-- gx_std_x6.vhd

-- Generated using ACDS version 15.1 185

library IEEE;
library gx_std_x6_altera_xcvr_native_a10_151;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity gx_std_x6 is
	port (
		reconfig_write          : in  std_logic_vector(0 downto 0)   := (others => '0'); --           reconfig_avmm.write
		reconfig_read           : in  std_logic_vector(0 downto 0)   := (others => '0'); --                        .read
		reconfig_address        : in  std_logic_vector(12 downto 0)  := (others => '0'); --                        .address
		reconfig_writedata      : in  std_logic_vector(31 downto 0)  := (others => '0'); --                        .writedata
		reconfig_readdata       : out std_logic_vector(31 downto 0);                     --                        .readdata
		reconfig_waitrequest    : out std_logic_vector(0 downto 0);                      --                        .waitrequest
		reconfig_clk            : in  std_logic_vector(0 downto 0)   := (others => '0'); --            reconfig_clk.clk
		reconfig_reset          : in  std_logic_vector(0 downto 0)   := (others => '0'); --          reconfig_reset.reset
		rx_analogreset          : in  std_logic_vector(5 downto 0)   := (others => '0'); --          rx_analogreset.rx_analogreset
		rx_cal_busy             : out std_logic_vector(5 downto 0);                      --             rx_cal_busy.rx_cal_busy
		rx_cdr_refclk0          : in  std_logic                      := '0';             --          rx_cdr_refclk0.clk
		rx_clkout               : out std_logic_vector(5 downto 0);                      --               rx_clkout.clk
		rx_coreclkin            : in  std_logic_vector(5 downto 0)   := (others => '0'); --            rx_coreclkin.clk
		rx_digitalreset         : in  std_logic_vector(5 downto 0)   := (others => '0'); --         rx_digitalreset.rx_digitalreset
		rx_is_lockedtodata      : out std_logic_vector(5 downto 0);                      --      rx_is_lockedtodata.rx_is_lockedtodata
		rx_is_lockedtoref       : out std_logic_vector(5 downto 0);                      --       rx_is_lockedtoref.rx_is_lockedtoref
		rx_parallel_data        : out std_logic_vector(119 downto 0);                    --        rx_parallel_data.rx_parallel_data
		rx_polinv               : in  std_logic_vector(5 downto 0)   := (others => '0'); --               rx_polinv.rx_polinv
		rx_serial_data          : in  std_logic_vector(5 downto 0)   := (others => '0'); --          rx_serial_data.rx_serial_data
		rx_seriallpbken         : in  std_logic_vector(5 downto 0)   := (others => '0'); --         rx_seriallpbken.rx_seriallpbken
		tx_analogreset          : in  std_logic_vector(5 downto 0)   := (others => '0'); --          tx_analogreset.tx_analogreset
		tx_bonding_clocks       : in  std_logic_vector(35 downto 0)  := (others => '0'); --       tx_bonding_clocks.clk
		tx_cal_busy             : out std_logic_vector(5 downto 0);                      --             tx_cal_busy.tx_cal_busy
		tx_clkout               : out std_logic_vector(5 downto 0);                      --               tx_clkout.clk
		tx_coreclkin            : in  std_logic_vector(5 downto 0)   := (others => '0'); --            tx_coreclkin.clk
		tx_digitalreset         : in  std_logic_vector(5 downto 0)   := (others => '0'); --         tx_digitalreset.tx_digitalreset
		tx_parallel_data        : in  std_logic_vector(119 downto 0) := (others => '0'); --        tx_parallel_data.tx_parallel_data
		tx_polinv               : in  std_logic_vector(5 downto 0)   := (others => '0'); --               tx_polinv.tx_polinv
		tx_serial_data          : out std_logic_vector(5 downto 0);                      --          tx_serial_data.tx_serial_data
		unused_rx_parallel_data : out std_logic_vector(647 downto 0);                    -- unused_rx_parallel_data.unused_rx_parallel_data
		unused_tx_parallel_data : in  std_logic_vector(647 downto 0) := (others => '0')  -- unused_tx_parallel_data.unused_tx_parallel_data
	);
end entity gx_std_x6;

architecture rtl of gx_std_x6 is
	component gx_std_x6_altera_xcvr_native_a10_151_eh2glbi is
		generic (
			device_revision                                                        : string  := "20nm5es";
			duplex_mode                                                            : string  := "duplex";
			channels                                                               : integer := 1;
			enable_calibration                                                     : integer := 0;
			enable_analog_resets                                                   : integer := 1;
			enable_reset_sequence                                                  : integer := 0;
			bonded_mode                                                            : string  := "not_bonded";
			pcs_bonding_master                                                     : integer := 0;
			plls                                                                   : integer := 1;
			number_physical_bonding_clocks                                         : integer := 1;
			cdr_refclk_cnt                                                         : integer := 1;
			enable_hip                                                             : integer := 0;
			hip_cal_en                                                             : string  := "disable";
			rcfg_enable                                                            : integer := 0;
			rcfg_shared                                                            : integer := 0;
			rcfg_jtag_enable                                                       : integer := 0;
			rcfg_separate_avmm_busy                                                : integer := 0;
			adme_prot_mode                                                         : string  := "basic_tx";
			adme_data_rate                                                         : string  := "5000000000";
			dbg_embedded_debug_enable                                              : integer := 0;
			dbg_capability_reg_enable                                              : integer := 0;
			dbg_user_identifier                                                    : integer := 0;
			dbg_stat_soft_logic_enable                                             : integer := 0;
			dbg_ctrl_soft_logic_enable                                             : integer := 0;
			dbg_prbs_soft_logic_enable                                             : integer := 0;
			dbg_odi_soft_logic_enable                                              : integer := 0;
			rcfg_emb_strm_enable                                                   : integer := 0;
			rcfg_profile_cnt                                                       : integer := 2;
			hssi_gen3_rx_pcs_block_sync                                            : string  := "enable_block_sync";
			hssi_gen3_rx_pcs_block_sync_sm                                         : string  := "enable_blk_sync_sm";
			hssi_gen3_rx_pcs_cdr_ctrl_force_unalgn                                 : string  := "enable";
			hssi_gen3_rx_pcs_lpbk_force                                            : string  := "lpbk_frce_dis";
			hssi_gen3_rx_pcs_mode                                                  : string  := "gen3_func";
			hssi_gen3_rx_pcs_rate_match_fifo                                       : string  := "enable_rm_fifo_600ppm";
			hssi_gen3_rx_pcs_rate_match_fifo_latency                               : string  := "regular_latency";
			hssi_gen3_rx_pcs_reverse_lpbk                                          : string  := "rev_lpbk_en";
			hssi_gen3_rx_pcs_rx_b4gb_par_lpbk                                      : string  := "b4gb_par_lpbk_dis";
			hssi_gen3_rx_pcs_rx_force_balign                                       : string  := "en_force_balign";
			hssi_gen3_rx_pcs_rx_ins_del_one_skip                                   : string  := "ins_del_one_skip_en";
			hssi_gen3_rx_pcs_rx_num_fixed_pat                                      : integer := 8;
			hssi_gen3_rx_pcs_rx_test_out_sel                                       : string  := "rx_test_out0";
			hssi_gen3_rx_pcs_sup_mode                                              : string  := "user_mode";
			hssi_gen3_tx_pcs_mode                                                  : string  := "gen3_func";
			hssi_gen3_tx_pcs_reverse_lpbk                                          : string  := "rev_lpbk_en";
			hssi_gen3_tx_pcs_sup_mode                                              : string  := "user_mode";
			hssi_gen3_tx_pcs_tx_bitslip                                            : integer := 0;
			hssi_gen3_tx_pcs_tx_gbox_byp                                           : string  := "bypass_gbox";
			hssi_krfec_rx_pcs_blksync_cor_en                                       : string  := "detect";
			hssi_krfec_rx_pcs_bypass_gb                                            : string  := "bypass_dis";
			hssi_krfec_rx_pcs_clr_ctrl                                             : string  := "both_enabled";
			hssi_krfec_rx_pcs_ctrl_bit_reverse                                     : string  := "ctrl_bit_reverse_dis";
			hssi_krfec_rx_pcs_data_bit_reverse                                     : string  := "data_bit_reverse_dis";
			hssi_krfec_rx_pcs_dv_start                                             : string  := "with_blklock";
			hssi_krfec_rx_pcs_err_mark_type                                        : string  := "err_mark_10g";
			hssi_krfec_rx_pcs_error_marking_en                                     : string  := "err_mark_dis";
			hssi_krfec_rx_pcs_low_latency_en                                       : string  := "disable";
			hssi_krfec_rx_pcs_lpbk_mode                                            : string  := "lpbk_dis";
			hssi_krfec_rx_pcs_parity_invalid_enum                                  : integer := 8;
			hssi_krfec_rx_pcs_parity_valid_num                                     : integer := 4;
			hssi_krfec_rx_pcs_pipeln_blksync                                       : string  := "enable";
			hssi_krfec_rx_pcs_pipeln_descrm                                        : string  := "enable";
			hssi_krfec_rx_pcs_pipeln_errcorrect                                    : string  := "enable";
			hssi_krfec_rx_pcs_pipeln_errtrap_ind                                   : string  := "enable";
			hssi_krfec_rx_pcs_pipeln_errtrap_lfsr                                  : string  := "enable";
			hssi_krfec_rx_pcs_pipeln_errtrap_loc                                   : string  := "enable";
			hssi_krfec_rx_pcs_pipeln_errtrap_pat                                   : string  := "enable";
			hssi_krfec_rx_pcs_pipeln_gearbox                                       : string  := "enable";
			hssi_krfec_rx_pcs_pipeln_syndrm                                        : string  := "enable";
			hssi_krfec_rx_pcs_pipeln_trans_dec                                     : string  := "enable";
			hssi_krfec_rx_pcs_prot_mode                                            : string  := "disable_mode";
			hssi_krfec_rx_pcs_receive_order                                        : string  := "receive_lsb";
			hssi_krfec_rx_pcs_rx_testbus_sel                                       : string  := "overall";
			hssi_krfec_rx_pcs_signal_ok_en                                         : string  := "sig_ok_dis";
			hssi_krfec_rx_pcs_sup_mode                                             : string  := "user_mode";
			hssi_krfec_tx_pcs_burst_err                                            : string  := "burst_err_dis";
			hssi_krfec_tx_pcs_burst_err_len                                        : string  := "burst_err_len1";
			hssi_krfec_tx_pcs_ctrl_bit_reverse                                     : string  := "ctrl_bit_reverse_dis";
			hssi_krfec_tx_pcs_data_bit_reverse                                     : string  := "data_bit_reverse_dis";
			hssi_krfec_tx_pcs_enc_frame_query                                      : string  := "enc_query_dis";
			hssi_krfec_tx_pcs_low_latency_en                                       : string  := "disable";
			hssi_krfec_tx_pcs_pipeln_encoder                                       : string  := "enable";
			hssi_krfec_tx_pcs_pipeln_scrambler                                     : string  := "enable";
			hssi_krfec_tx_pcs_prot_mode                                            : string  := "disable_mode";
			hssi_krfec_tx_pcs_sup_mode                                             : string  := "user_mode";
			hssi_krfec_tx_pcs_transcode_err                                        : string  := "trans_err_dis";
			hssi_krfec_tx_pcs_transmit_order                                       : string  := "transmit_lsb";
			hssi_krfec_tx_pcs_tx_testbus_sel                                       : string  := "overall";
			hssi_10g_rx_pcs_align_del                                              : string  := "align_del_en";
			hssi_10g_rx_pcs_ber_bit_err_total_cnt                                  : string  := "bit_err_total_cnt_10g";
			hssi_10g_rx_pcs_ber_clken                                              : string  := "ber_clk_dis";
			hssi_10g_rx_pcs_ber_xus_timer_window                                   : integer := 19530;
			hssi_10g_rx_pcs_bitslip_mode                                           : string  := "bitslip_dis";
			hssi_10g_rx_pcs_blksync_bitslip_type                                   : string  := "bitslip_comb";
			hssi_10g_rx_pcs_blksync_bitslip_wait_cnt                               : integer := 1;
			hssi_10g_rx_pcs_blksync_bitslip_wait_type                              : string  := "bitslip_match";
			hssi_10g_rx_pcs_blksync_bypass                                         : string  := "blksync_bypass_dis";
			hssi_10g_rx_pcs_blksync_clken                                          : string  := "blksync_clk_dis";
			hssi_10g_rx_pcs_blksync_enum_invalid_sh_cnt                            : string  := "enum_invalid_sh_cnt_10g";
			hssi_10g_rx_pcs_blksync_knum_sh_cnt_postlock                           : string  := "knum_sh_cnt_postlock_10g";
			hssi_10g_rx_pcs_blksync_knum_sh_cnt_prelock                            : string  := "knum_sh_cnt_prelock_10g";
			hssi_10g_rx_pcs_blksync_pipeln                                         : string  := "blksync_pipeln_dis";
			hssi_10g_rx_pcs_clr_errblk_cnt_en                                      : string  := "disable";
			hssi_10g_rx_pcs_control_del                                            : string  := "control_del_all";
			hssi_10g_rx_pcs_crcchk_bypass                                          : string  := "crcchk_bypass_dis";
			hssi_10g_rx_pcs_crcchk_clken                                           : string  := "crcchk_clk_dis";
			hssi_10g_rx_pcs_crcchk_inv                                             : string  := "crcchk_inv_dis";
			hssi_10g_rx_pcs_crcchk_pipeln                                          : string  := "crcchk_pipeln_dis";
			hssi_10g_rx_pcs_crcflag_pipeln                                         : string  := "crcflag_pipeln_dis";
			hssi_10g_rx_pcs_ctrl_bit_reverse                                       : string  := "ctrl_bit_reverse_dis";
			hssi_10g_rx_pcs_data_bit_reverse                                       : string  := "data_bit_reverse_dis";
			hssi_10g_rx_pcs_dec_64b66b_rxsm_bypass                                 : string  := "dec_64b66b_rxsm_bypass_dis";
			hssi_10g_rx_pcs_dec64b66b_clken                                        : string  := "dec64b66b_clk_dis";
			hssi_10g_rx_pcs_descrm_bypass                                          : string  := "descrm_bypass_en";
			hssi_10g_rx_pcs_descrm_clken                                           : string  := "descrm_clk_dis";
			hssi_10g_rx_pcs_descrm_mode                                            : string  := "async";
			hssi_10g_rx_pcs_descrm_pipeln                                          : string  := "enable";
			hssi_10g_rx_pcs_dft_clk_out_sel                                        : string  := "rx_master_clk";
			hssi_10g_rx_pcs_dis_signal_ok                                          : string  := "dis_signal_ok_dis";
			hssi_10g_rx_pcs_dispchk_bypass                                         : string  := "dispchk_bypass_dis";
			hssi_10g_rx_pcs_empty_flag_type                                        : string  := "empty_rd_side";
			hssi_10g_rx_pcs_fast_path                                              : string  := "fast_path_dis";
			hssi_10g_rx_pcs_fec_clken                                              : string  := "fec_clk_dis";
			hssi_10g_rx_pcs_fec_enable                                             : string  := "fec_dis";
			hssi_10g_rx_pcs_fifo_double_read                                       : string  := "fifo_double_read_dis";
			hssi_10g_rx_pcs_fifo_stop_rd                                           : string  := "n_rd_empty";
			hssi_10g_rx_pcs_fifo_stop_wr                                           : string  := "n_wr_full";
			hssi_10g_rx_pcs_force_align                                            : string  := "force_align_dis";
			hssi_10g_rx_pcs_frmsync_bypass                                         : string  := "frmsync_bypass_dis";
			hssi_10g_rx_pcs_frmsync_clken                                          : string  := "frmsync_clk_dis";
			hssi_10g_rx_pcs_frmsync_enum_scrm                                      : string  := "enum_scrm_default";
			hssi_10g_rx_pcs_frmsync_enum_sync                                      : string  := "enum_sync_default";
			hssi_10g_rx_pcs_frmsync_flag_type                                      : string  := "all_framing_words";
			hssi_10g_rx_pcs_frmsync_knum_sync                                      : string  := "knum_sync_default";
			hssi_10g_rx_pcs_frmsync_mfrm_length                                    : integer := 2048;
			hssi_10g_rx_pcs_frmsync_pipeln                                         : string  := "frmsync_pipeln_dis";
			hssi_10g_rx_pcs_full_flag_type                                         : string  := "full_wr_side";
			hssi_10g_rx_pcs_gb_rx_idwidth                                          : string  := "width_32";
			hssi_10g_rx_pcs_gb_rx_odwidth                                          : string  := "width_66";
			hssi_10g_rx_pcs_gbexp_clken                                            : string  := "gbexp_clk_dis";
			hssi_10g_rx_pcs_low_latency_en                                         : string  := "enable";
			hssi_10g_rx_pcs_lpbk_mode                                              : string  := "lpbk_dis";
			hssi_10g_rx_pcs_master_clk_sel                                         : string  := "master_rx_pma_clk";
			hssi_10g_rx_pcs_pempty_flag_type                                       : string  := "pempty_rd_side";
			hssi_10g_rx_pcs_pfull_flag_type                                        : string  := "pfull_wr_side";
			hssi_10g_rx_pcs_phcomp_rd_del                                          : string  := "phcomp_rd_del2";
			hssi_10g_rx_pcs_pld_if_type                                            : string  := "fifo";
			hssi_10g_rx_pcs_prot_mode                                              : string  := "disable_mode";
			hssi_10g_rx_pcs_rand_clken                                             : string  := "rand_clk_dis";
			hssi_10g_rx_pcs_rd_clk_sel                                             : string  := "rd_rx_pma_clk";
			hssi_10g_rx_pcs_rdfifo_clken                                           : string  := "rdfifo_clk_dis";
			hssi_10g_rx_pcs_rx_fifo_write_ctrl                                     : string  := "blklock_stops";
			hssi_10g_rx_pcs_rx_scrm_width                                          : string  := "bit64";
			hssi_10g_rx_pcs_rx_sh_location                                         : string  := "lsb";
			hssi_10g_rx_pcs_rx_signal_ok_sel                                       : string  := "synchronized_ver";
			hssi_10g_rx_pcs_rx_sm_bypass                                           : string  := "rx_sm_bypass_dis";
			hssi_10g_rx_pcs_rx_sm_hiber                                            : string  := "rx_sm_hiber_en";
			hssi_10g_rx_pcs_rx_sm_pipeln                                           : string  := "rx_sm_pipeln_dis";
			hssi_10g_rx_pcs_rx_testbus_sel                                         : string  := "rx_fifo_testbus1";
			hssi_10g_rx_pcs_rx_true_b2b                                            : string  := "b2b";
			hssi_10g_rx_pcs_rxfifo_empty                                           : string  := "empty_default";
			hssi_10g_rx_pcs_rxfifo_full                                            : string  := "full_default";
			hssi_10g_rx_pcs_rxfifo_mode                                            : string  := "phase_comp";
			hssi_10g_rx_pcs_rxfifo_pempty                                          : integer := 2;
			hssi_10g_rx_pcs_rxfifo_pfull                                           : integer := 23;
			hssi_10g_rx_pcs_stretch_num_stages                                     : string  := "zero_stage";
			hssi_10g_rx_pcs_sup_mode                                               : string  := "user_mode";
			hssi_10g_rx_pcs_test_mode                                              : string  := "test_off";
			hssi_10g_rx_pcs_wrfifo_clken                                           : string  := "wrfifo_clk_dis";
			hssi_10g_rx_pcs_advanced_user_mode                                     : string  := "disable";
			hssi_10g_tx_pcs_bitslip_en                                             : string  := "bitslip_dis";
			hssi_10g_tx_pcs_bonding_dft_en                                         : string  := "dft_dis";
			hssi_10g_tx_pcs_bonding_dft_val                                        : string  := "dft_0";
			hssi_10g_tx_pcs_crcgen_bypass                                          : string  := "crcgen_bypass_dis";
			hssi_10g_tx_pcs_crcgen_clken                                           : string  := "crcgen_clk_dis";
			hssi_10g_tx_pcs_crcgen_err                                             : string  := "crcgen_err_dis";
			hssi_10g_tx_pcs_crcgen_inv                                             : string  := "crcgen_inv_dis";
			hssi_10g_tx_pcs_ctrl_bit_reverse                                       : string  := "ctrl_bit_reverse_dis";
			hssi_10g_tx_pcs_data_bit_reverse                                       : string  := "data_bit_reverse_dis";
			hssi_10g_tx_pcs_dft_clk_out_sel                                        : string  := "tx_master_clk";
			hssi_10g_tx_pcs_dispgen_bypass                                         : string  := "dispgen_bypass_dis";
			hssi_10g_tx_pcs_dispgen_clken                                          : string  := "dispgen_clk_dis";
			hssi_10g_tx_pcs_dispgen_err                                            : string  := "dispgen_err_dis";
			hssi_10g_tx_pcs_dispgen_pipeln                                         : string  := "dispgen_pipeln_dis";
			hssi_10g_tx_pcs_empty_flag_type                                        : string  := "empty_rd_side";
			hssi_10g_tx_pcs_enc_64b66b_txsm_bypass                                 : string  := "enc_64b66b_txsm_bypass_dis";
			hssi_10g_tx_pcs_enc64b66b_txsm_clken                                   : string  := "enc64b66b_txsm_clk_dis";
			hssi_10g_tx_pcs_fastpath                                               : string  := "fastpath_dis";
			hssi_10g_tx_pcs_fec_clken                                              : string  := "fec_clk_dis";
			hssi_10g_tx_pcs_fec_enable                                             : string  := "fec_dis";
			hssi_10g_tx_pcs_fifo_double_write                                      : string  := "fifo_double_write_dis";
			hssi_10g_tx_pcs_fifo_reg_fast                                          : string  := "fifo_reg_fast_dis";
			hssi_10g_tx_pcs_fifo_stop_rd                                           : string  := "n_rd_empty";
			hssi_10g_tx_pcs_fifo_stop_wr                                           : string  := "n_wr_full";
			hssi_10g_tx_pcs_frmgen_burst                                           : string  := "frmgen_burst_dis";
			hssi_10g_tx_pcs_frmgen_bypass                                          : string  := "frmgen_bypass_dis";
			hssi_10g_tx_pcs_frmgen_clken                                           : string  := "frmgen_clk_dis";
			hssi_10g_tx_pcs_frmgen_mfrm_length                                     : integer := 2048;
			hssi_10g_tx_pcs_frmgen_pipeln                                          : string  := "frmgen_pipeln_dis";
			hssi_10g_tx_pcs_frmgen_pyld_ins                                        : string  := "frmgen_pyld_ins_dis";
			hssi_10g_tx_pcs_frmgen_wordslip                                        : string  := "frmgen_wordslip_dis";
			hssi_10g_tx_pcs_full_flag_type                                         : string  := "full_wr_side";
			hssi_10g_tx_pcs_gb_pipeln_bypass                                       : string  := "disable";
			hssi_10g_tx_pcs_gb_tx_idwidth                                          : string  := "width_50";
			hssi_10g_tx_pcs_gb_tx_odwidth                                          : string  := "width_32";
			hssi_10g_tx_pcs_gbred_clken                                            : string  := "gbred_clk_dis";
			hssi_10g_tx_pcs_low_latency_en                                         : string  := "enable";
			hssi_10g_tx_pcs_master_clk_sel                                         : string  := "master_tx_pma_clk";
			hssi_10g_tx_pcs_pempty_flag_type                                       : string  := "pempty_rd_side";
			hssi_10g_tx_pcs_pfull_flag_type                                        : string  := "pfull_wr_side";
			hssi_10g_tx_pcs_phcomp_rd_del                                          : string  := "phcomp_rd_del2";
			hssi_10g_tx_pcs_pld_if_type                                            : string  := "fifo";
			hssi_10g_tx_pcs_prot_mode                                              : string  := "disable_mode";
			hssi_10g_tx_pcs_pseudo_random                                          : string  := "all_0";
			hssi_10g_tx_pcs_pseudo_seed_a                                          : string  := "288230376151711743";
			hssi_10g_tx_pcs_pseudo_seed_b                                          : string  := "288230376151711743";
			hssi_10g_tx_pcs_random_disp                                            : string  := "disable";
			hssi_10g_tx_pcs_rdfifo_clken                                           : string  := "rdfifo_clk_dis";
			hssi_10g_tx_pcs_scrm_bypass                                            : string  := "scrm_bypass_dis";
			hssi_10g_tx_pcs_scrm_clken                                             : string  := "scrm_clk_dis";
			hssi_10g_tx_pcs_scrm_mode                                              : string  := "async";
			hssi_10g_tx_pcs_scrm_pipeln                                            : string  := "enable";
			hssi_10g_tx_pcs_sh_err                                                 : string  := "sh_err_dis";
			hssi_10g_tx_pcs_sop_mark                                               : string  := "sop_mark_dis";
			hssi_10g_tx_pcs_stretch_num_stages                                     : string  := "zero_stage";
			hssi_10g_tx_pcs_sup_mode                                               : string  := "user_mode";
			hssi_10g_tx_pcs_test_mode                                              : string  := "test_off";
			hssi_10g_tx_pcs_tx_scrm_err                                            : string  := "scrm_err_dis";
			hssi_10g_tx_pcs_tx_scrm_width                                          : string  := "bit64";
			hssi_10g_tx_pcs_tx_sh_location                                         : string  := "lsb";
			hssi_10g_tx_pcs_tx_sm_bypass                                           : string  := "tx_sm_bypass_dis";
			hssi_10g_tx_pcs_tx_sm_pipeln                                           : string  := "tx_sm_pipeln_dis";
			hssi_10g_tx_pcs_tx_testbus_sel                                         : string  := "tx_fifo_testbus1";
			hssi_10g_tx_pcs_txfifo_empty                                           : string  := "empty_default";
			hssi_10g_tx_pcs_txfifo_full                                            : string  := "full_default";
			hssi_10g_tx_pcs_txfifo_mode                                            : string  := "phase_comp";
			hssi_10g_tx_pcs_txfifo_pempty                                          : integer := 2;
			hssi_10g_tx_pcs_txfifo_pfull                                           : integer := 11;
			hssi_10g_tx_pcs_wr_clk_sel                                             : string  := "wr_tx_pma_clk";
			hssi_10g_tx_pcs_wrfifo_clken                                           : string  := "wrfifo_clk_dis";
			hssi_10g_tx_pcs_advanced_user_mode                                     : string  := "disable";
			hssi_8g_rx_pcs_auto_error_replacement                                  : string  := "dis_err_replace";
			hssi_8g_rx_pcs_bit_reversal                                            : string  := "dis_bit_reversal";
			hssi_8g_rx_pcs_bonding_dft_en                                          : string  := "dft_dis";
			hssi_8g_rx_pcs_bonding_dft_val                                         : string  := "dft_0";
			hssi_8g_rx_pcs_bypass_pipeline_reg                                     : string  := "dis_bypass_pipeline";
			hssi_8g_rx_pcs_byte_deserializer                                       : string  := "dis_bds";
			hssi_8g_rx_pcs_cdr_ctrl_rxvalid_mask                                   : string  := "dis_rxvalid_mask";
			hssi_8g_rx_pcs_clkcmp_pattern_n                                        : integer := 0;
			hssi_8g_rx_pcs_clkcmp_pattern_p                                        : integer := 0;
			hssi_8g_rx_pcs_clock_gate_bds_dec_asn                                  : string  := "dis_bds_dec_asn_clk_gating";
			hssi_8g_rx_pcs_clock_gate_cdr_eidle                                    : string  := "dis_cdr_eidle_clk_gating";
			hssi_8g_rx_pcs_clock_gate_dw_pc_wrclk                                  : string  := "dis_dw_pc_wrclk_gating";
			hssi_8g_rx_pcs_clock_gate_dw_rm_rd                                     : string  := "dis_dw_rm_rdclk_gating";
			hssi_8g_rx_pcs_clock_gate_dw_rm_wr                                     : string  := "dis_dw_rm_wrclk_gating";
			hssi_8g_rx_pcs_clock_gate_dw_wa                                        : string  := "dis_dw_wa_clk_gating";
			hssi_8g_rx_pcs_clock_gate_pc_rdclk                                     : string  := "dis_pc_rdclk_gating";
			hssi_8g_rx_pcs_clock_gate_sw_pc_wrclk                                  : string  := "dis_sw_pc_wrclk_gating";
			hssi_8g_rx_pcs_clock_gate_sw_rm_rd                                     : string  := "dis_sw_rm_rdclk_gating";
			hssi_8g_rx_pcs_clock_gate_sw_rm_wr                                     : string  := "dis_sw_rm_wrclk_gating";
			hssi_8g_rx_pcs_clock_gate_sw_wa                                        : string  := "dis_sw_wa_clk_gating";
			hssi_8g_rx_pcs_clock_observation_in_pld_core                           : string  := "internal_sw_wa_clk";
			hssi_8g_rx_pcs_eidle_entry_eios                                        : string  := "dis_eidle_eios";
			hssi_8g_rx_pcs_eidle_entry_iei                                         : string  := "dis_eidle_iei";
			hssi_8g_rx_pcs_eidle_entry_sd                                          : string  := "dis_eidle_sd";
			hssi_8g_rx_pcs_eightb_tenb_decoder                                     : string  := "dis_8b10b";
			hssi_8g_rx_pcs_err_flags_sel                                           : string  := "err_flags_wa";
			hssi_8g_rx_pcs_fixed_pat_det                                           : string  := "dis_fixed_patdet";
			hssi_8g_rx_pcs_fixed_pat_num                                           : integer := 15;
			hssi_8g_rx_pcs_force_signal_detect                                     : string  := "en_force_signal_detect";
			hssi_8g_rx_pcs_gen3_clk_en                                             : string  := "disable_clk";
			hssi_8g_rx_pcs_gen3_rx_clk_sel                                         : string  := "rcvd_clk";
			hssi_8g_rx_pcs_gen3_tx_clk_sel                                         : string  := "tx_pma_clk";
			hssi_8g_rx_pcs_hip_mode                                                : string  := "dis_hip";
			hssi_8g_rx_pcs_ibm_invalid_code                                        : string  := "dis_ibm_invalid_code";
			hssi_8g_rx_pcs_invalid_code_flag_only                                  : string  := "dis_invalid_code_only";
			hssi_8g_rx_pcs_pad_or_edb_error_replace                                : string  := "replace_edb";
			hssi_8g_rx_pcs_pcs_bypass                                              : string  := "dis_pcs_bypass";
			hssi_8g_rx_pcs_phase_comp_rdptr                                        : string  := "enable_rdptr";
			hssi_8g_rx_pcs_phase_compensation_fifo                                 : string  := "low_latency";
			hssi_8g_rx_pcs_pipe_if_enable                                          : string  := "dis_pipe_rx";
			hssi_8g_rx_pcs_pma_dw                                                  : string  := "eight_bit";
			hssi_8g_rx_pcs_polinv_8b10b_dec                                        : string  := "dis_polinv_8b10b_dec";
			hssi_8g_rx_pcs_prot_mode                                               : string  := "gige";
			hssi_8g_rx_pcs_rate_match                                              : string  := "dis_rm";
			hssi_8g_rx_pcs_rate_match_del_thres                                    : string  := "dis_rm_del_thres";
			hssi_8g_rx_pcs_rate_match_empty_thres                                  : string  := "dis_rm_empty_thres";
			hssi_8g_rx_pcs_rate_match_full_thres                                   : string  := "dis_rm_full_thres";
			hssi_8g_rx_pcs_rate_match_ins_thres                                    : string  := "dis_rm_ins_thres";
			hssi_8g_rx_pcs_rate_match_start_thres                                  : string  := "dis_rm_start_thres";
			hssi_8g_rx_pcs_rx_clk_free_running                                     : string  := "en_rx_clk_free_run";
			hssi_8g_rx_pcs_rx_clk2                                                 : string  := "rcvd_clk_clk2";
			hssi_8g_rx_pcs_rx_pcs_urst                                             : string  := "en_rx_pcs_urst";
			hssi_8g_rx_pcs_rx_rcvd_clk                                             : string  := "rcvd_clk_rcvd_clk";
			hssi_8g_rx_pcs_rx_rd_clk                                               : string  := "pld_rx_clk";
			hssi_8g_rx_pcs_rx_refclk                                               : string  := "dis_refclk_sel";
			hssi_8g_rx_pcs_rx_wr_clk                                               : string  := "rx_clk2_div_1_2_4";
			hssi_8g_rx_pcs_sup_mode                                                : string  := "user_mode";
			hssi_8g_rx_pcs_symbol_swap                                             : string  := "dis_symbol_swap";
			hssi_8g_rx_pcs_sync_sm_idle_eios                                       : string  := "dis_syncsm_idle";
			hssi_8g_rx_pcs_test_bus_sel                                            : string  := "tx_testbus";
			hssi_8g_rx_pcs_tx_rx_parallel_loopback                                 : string  := "dis_plpbk";
			hssi_8g_rx_pcs_wa_boundary_lock_ctrl                                   : string  := "bit_slip";
			hssi_8g_rx_pcs_wa_clk_slip_spacing                                     : integer := 16;
			hssi_8g_rx_pcs_wa_det_latency_sync_status_beh                          : string  := "dont_care_assert_sync";
			hssi_8g_rx_pcs_wa_disp_err_flag                                        : string  := "dis_disp_err_flag";
			hssi_8g_rx_pcs_wa_kchar                                                : string  := "dis_kchar";
			hssi_8g_rx_pcs_wa_pd                                                   : string  := "wa_pd_10";
			hssi_8g_rx_pcs_wa_pd_data                                              : string  := "0";
			hssi_8g_rx_pcs_wa_pd_polarity                                          : string  := "dis_pd_both_pol";
			hssi_8g_rx_pcs_wa_pld_controlled                                       : string  := "dis_pld_ctrl";
			hssi_8g_rx_pcs_wa_renumber_data                                        : integer := 0;
			hssi_8g_rx_pcs_wa_rgnumber_data                                        : integer := 0;
			hssi_8g_rx_pcs_wa_rknumber_data                                        : integer := 0;
			hssi_8g_rx_pcs_wa_rosnumber_data                                       : integer := 0;
			hssi_8g_rx_pcs_wa_rvnumber_data                                        : integer := 0;
			hssi_8g_rx_pcs_wa_sync_sm_ctrl                                         : string  := "gige_sync_sm";
			hssi_8g_rx_pcs_wait_cnt                                                : integer := 0;
			hssi_8g_tx_pcs_bit_reversal                                            : string  := "dis_bit_reversal";
			hssi_8g_tx_pcs_bonding_dft_en                                          : string  := "dft_dis";
			hssi_8g_tx_pcs_bonding_dft_val                                         : string  := "dft_0";
			hssi_8g_tx_pcs_bypass_pipeline_reg                                     : string  := "dis_bypass_pipeline";
			hssi_8g_tx_pcs_byte_serializer                                         : string  := "dis_bs";
			hssi_8g_tx_pcs_clock_gate_bs_enc                                       : string  := "dis_bs_enc_clk_gating";
			hssi_8g_tx_pcs_clock_gate_dw_fifowr                                    : string  := "dis_dw_fifowr_clk_gating";
			hssi_8g_tx_pcs_clock_gate_fiford                                       : string  := "dis_fiford_clk_gating";
			hssi_8g_tx_pcs_clock_gate_sw_fifowr                                    : string  := "dis_sw_fifowr_clk_gating";
			hssi_8g_tx_pcs_clock_observation_in_pld_core                           : string  := "internal_refclk_b";
			hssi_8g_tx_pcs_data_selection_8b10b_encoder_input                      : string  := "normal_data_path";
			hssi_8g_tx_pcs_dynamic_clk_switch                                      : string  := "dis_dyn_clk_switch";
			hssi_8g_tx_pcs_eightb_tenb_disp_ctrl                                   : string  := "dis_disp_ctrl";
			hssi_8g_tx_pcs_eightb_tenb_encoder                                     : string  := "dis_8b10b";
			hssi_8g_tx_pcs_force_echar                                             : string  := "dis_force_echar";
			hssi_8g_tx_pcs_force_kchar                                             : string  := "dis_force_kchar";
			hssi_8g_tx_pcs_gen3_tx_clk_sel                                         : string  := "tx_pma_clk";
			hssi_8g_tx_pcs_gen3_tx_pipe_clk_sel                                    : string  := "func_clk";
			hssi_8g_tx_pcs_hip_mode                                                : string  := "dis_hip";
			hssi_8g_tx_pcs_pcs_bypass                                              : string  := "dis_pcs_bypass";
			hssi_8g_tx_pcs_phase_comp_rdptr                                        : string  := "enable_rdptr";
			hssi_8g_tx_pcs_phase_compensation_fifo                                 : string  := "low_latency";
			hssi_8g_tx_pcs_phfifo_write_clk_sel                                    : string  := "pld_tx_clk";
			hssi_8g_tx_pcs_pma_dw                                                  : string  := "eight_bit";
			hssi_8g_tx_pcs_prot_mode                                               : string  := "basic";
			hssi_8g_tx_pcs_refclk_b_clk_sel                                        : string  := "tx_pma_clock";
			hssi_8g_tx_pcs_revloop_back_rm                                         : string  := "dis_rev_loopback_rx_rm";
			hssi_8g_tx_pcs_sup_mode                                                : string  := "user_mode";
			hssi_8g_tx_pcs_symbol_swap                                             : string  := "dis_symbol_swap";
			hssi_8g_tx_pcs_tx_bitslip                                              : string  := "dis_tx_bitslip";
			hssi_8g_tx_pcs_tx_compliance_controlled_disparity                      : string  := "dis_txcompliance";
			hssi_8g_tx_pcs_tx_fast_pld_reg                                         : string  := "dis_tx_fast_pld_reg";
			hssi_8g_tx_pcs_txclk_freerun                                           : string  := "dis_freerun_tx";
			hssi_8g_tx_pcs_txpcs_urst                                              : string  := "en_txpcs_urst";
			hssi_tx_pld_pcs_interface_hd_chnl_hip_en                               : string  := "disable";
			hssi_tx_pld_pcs_interface_hd_chnl_hrdrstctl_en                         : string  := "disable";
			hssi_tx_pld_pcs_interface_hd_chnl_prot_mode_tx                         : string  := "disabled_prot_mode_tx";
			hssi_tx_pld_pcs_interface_hd_chnl_ctrl_plane_bonding_tx                : string  := "individual_tx";
			hssi_tx_pld_pcs_interface_hd_chnl_pma_dw_tx                            : string  := "pma_8b_tx";
			hssi_tx_pld_pcs_interface_hd_chnl_pld_fifo_mode_tx                     : string  := "fifo_tx";
			hssi_tx_pld_pcs_interface_hd_chnl_shared_fifo_width_tx                 : string  := "single_tx";
			hssi_tx_pld_pcs_interface_hd_chnl_low_latency_en_tx                    : string  := "disable";
			hssi_tx_pld_pcs_interface_hd_chnl_func_mode                            : string  := "enable";
			hssi_tx_pld_pcs_interface_hd_chnl_channel_operation_mode               : string  := "tx_rx_pair_enabled";
			hssi_tx_pld_pcs_interface_hd_chnl_lpbk_en                              : string  := "disable";
			hssi_tx_pld_pcs_interface_hd_chnl_frequency_rules_en                   : string  := "enable";
			hssi_tx_pld_pcs_interface_hd_chnl_pma_tx_clk_hz                        : integer := 0;
			hssi_tx_pld_pcs_interface_hd_chnl_pld_tx_clk_hz                        : integer := 0;
			hssi_tx_pld_pcs_interface_hd_chnl_pld_uhsif_tx_clk_hz                  : integer := 0;
			hssi_tx_pld_pcs_interface_hd_fifo_channel_operation_mode               : string  := "tx_rx_pair_enabled";
			hssi_tx_pld_pcs_interface_hd_fifo_prot_mode_tx                         : string  := "teng_mode_tx";
			hssi_tx_pld_pcs_interface_hd_fifo_shared_fifo_width_tx                 : string  := "single_tx";
			hssi_tx_pld_pcs_interface_hd_10g_channel_operation_mode                : string  := "tx_rx_pair_enabled";
			hssi_tx_pld_pcs_interface_hd_10g_lpbk_en                               : string  := "disable";
			hssi_tx_pld_pcs_interface_hd_10g_advanced_user_mode_tx                 : string  := "disable";
			hssi_tx_pld_pcs_interface_hd_10g_pma_dw_tx                             : string  := "pma_64b_tx";
			hssi_tx_pld_pcs_interface_hd_10g_fifo_mode_tx                          : string  := "fifo_tx";
			hssi_tx_pld_pcs_interface_hd_10g_prot_mode_tx                          : string  := "disabled_prot_mode_tx";
			hssi_tx_pld_pcs_interface_hd_10g_low_latency_en_tx                     : string  := "enable";
			hssi_tx_pld_pcs_interface_hd_10g_shared_fifo_width_tx                  : string  := "single_tx";
			hssi_tx_pld_pcs_interface_hd_8g_channel_operation_mode                 : string  := "tx_rx_pair_enabled";
			hssi_tx_pld_pcs_interface_hd_8g_lpbk_en                                : string  := "disable";
			hssi_tx_pld_pcs_interface_hd_8g_prot_mode_tx                           : string  := "disabled_prot_mode_tx";
			hssi_tx_pld_pcs_interface_hd_8g_hip_mode                               : string  := "disable";
			hssi_tx_pld_pcs_interface_hd_8g_pma_dw_tx                              : string  := "pma_8b_tx";
			hssi_tx_pld_pcs_interface_hd_8g_fifo_mode_tx                           : string  := "fifo_tx";
			hssi_tx_pld_pcs_interface_hd_g3_prot_mode                              : string  := "disabled_prot_mode";
			hssi_tx_pld_pcs_interface_hd_krfec_channel_operation_mode              : string  := "tx_rx_pair_enabled";
			hssi_tx_pld_pcs_interface_hd_krfec_lpbk_en                             : string  := "disable";
			hssi_tx_pld_pcs_interface_hd_krfec_prot_mode_tx                        : string  := "disabled_prot_mode_tx";
			hssi_tx_pld_pcs_interface_hd_krfec_low_latency_en_tx                   : string  := "disable";
			hssi_tx_pld_pcs_interface_hd_pmaif_lpbk_en                             : string  := "disable";
			hssi_tx_pld_pcs_interface_hd_pmaif_channel_operation_mode              : string  := "tx_rx_pair_enabled";
			hssi_tx_pld_pcs_interface_hd_pmaif_sim_mode                            : string  := "disable";
			hssi_tx_pld_pcs_interface_hd_pmaif_prot_mode_tx                        : string  := "disabled_prot_mode_tx";
			hssi_tx_pld_pcs_interface_hd_pmaif_pma_dw_tx                           : string  := "pma_8b_tx";
			hssi_tx_pld_pcs_interface_hd_pldif_prot_mode_tx                        : string  := "disabled_prot_mode_tx";
			hssi_tx_pld_pcs_interface_hd_pldif_hrdrstctl_en                        : string  := "disable";
			hssi_tx_pld_pcs_interface_pcs_tx_clk_source                            : string  := "teng";
			hssi_tx_pld_pcs_interface_pcs_tx_data_source                           : string  := "hip_disable";
			hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_en                         : string  := "delay1_clk_disable";
			hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_sel                        : string  := "pld_tx_clk";
			hssi_tx_pld_pcs_interface_pcs_tx_delay1_ctrl                           : string  := "delay1_path0";
			hssi_tx_pld_pcs_interface_pcs_tx_delay1_data_sel                       : string  := "one_ff_delay";
			hssi_tx_pld_pcs_interface_pcs_tx_delay2_clk_en                         : string  := "delay2_clk_disable";
			hssi_tx_pld_pcs_interface_pcs_tx_delay2_ctrl                           : string  := "delay2_path0";
			hssi_tx_pld_pcs_interface_pcs_tx_output_sel                            : string  := "teng_output";
			hssi_tx_pld_pcs_interface_pcs_tx_clk_out_sel                           : string  := "teng_clk_out";
			hssi_rx_pld_pcs_interface_hd_chnl_hip_en                               : string  := "disable";
			hssi_rx_pld_pcs_interface_hd_chnl_transparent_pcs_rx                   : string  := "disable";
			hssi_rx_pld_pcs_interface_hd_chnl_hrdrstctl_en                         : string  := "disable";
			hssi_rx_pld_pcs_interface_hd_chnl_prot_mode_rx                         : string  := "disabled_prot_mode_rx";
			hssi_rx_pld_pcs_interface_hd_chnl_ctrl_plane_bonding_rx                : string  := "individual_rx";
			hssi_rx_pld_pcs_interface_hd_chnl_pma_dw_rx                            : string  := "pma_8b_rx";
			hssi_rx_pld_pcs_interface_hd_chnl_pld_fifo_mode_rx                     : string  := "fifo_rx";
			hssi_rx_pld_pcs_interface_hd_chnl_shared_fifo_width_rx                 : string  := "single_rx";
			hssi_rx_pld_pcs_interface_hd_chnl_low_latency_en_rx                    : string  := "disable";
			hssi_rx_pld_pcs_interface_hd_chnl_func_mode                            : string  := "enable";
			hssi_rx_pld_pcs_interface_hd_chnl_channel_operation_mode               : string  := "tx_rx_pair_enabled";
			hssi_rx_pld_pcs_interface_hd_chnl_lpbk_en                              : string  := "disable";
			hssi_rx_pld_pcs_interface_hd_10g_advanced_user_mode_rx                 : string  := "disable";
			hssi_rx_pld_pcs_interface_hd_chnl_frequency_rules_en                   : string  := "enable";
			hssi_rx_pld_pcs_interface_hd_chnl_pma_rx_clk_hz                        : integer := 0;
			hssi_rx_pld_pcs_interface_hd_chnl_pld_rx_clk_hz                        : integer := 0;
			hssi_rx_pld_pcs_interface_hd_chnl_fref_clk_hz                          : integer := 0;
			hssi_rx_pld_pcs_interface_hd_chnl_clklow_clk_hz                        : integer := 0;
			hssi_rx_pld_pcs_interface_hd_fifo_channel_operation_mode               : string  := "tx_rx_pair_enabled";
			hssi_rx_pld_pcs_interface_hd_fifo_prot_mode_rx                         : string  := "teng_mode_rx";
			hssi_rx_pld_pcs_interface_hd_fifo_shared_fifo_width_rx                 : string  := "single_rx";
			hssi_rx_pld_pcs_interface_hd_10g_channel_operation_mode                : string  := "tx_rx_pair_enabled";
			hssi_rx_pld_pcs_interface_hd_10g_lpbk_en                               : string  := "disable";
			hssi_rx_pld_pcs_interface_hd_10g_pma_dw_rx                             : string  := "pma_64b_rx";
			hssi_rx_pld_pcs_interface_hd_10g_fifo_mode_rx                          : string  := "fifo_rx";
			hssi_rx_pld_pcs_interface_hd_10g_prot_mode_rx                          : string  := "disabled_prot_mode_rx";
			hssi_rx_pld_pcs_interface_hd_10g_low_latency_en_rx                     : string  := "enable";
			hssi_rx_pld_pcs_interface_hd_10g_shared_fifo_width_rx                  : string  := "single_rx";
			hssi_rx_pld_pcs_interface_hd_10g_test_bus_mode                         : string  := "tx";
			hssi_rx_pld_pcs_interface_hd_8g_channel_operation_mode                 : string  := "tx_rx_pair_enabled";
			hssi_rx_pld_pcs_interface_hd_8g_lpbk_en                                : string  := "disable";
			hssi_rx_pld_pcs_interface_hd_8g_prot_mode_rx                           : string  := "disabled_prot_mode_rx";
			hssi_rx_pld_pcs_interface_hd_8g_hip_mode                               : string  := "disable";
			hssi_rx_pld_pcs_interface_hd_8g_pma_dw_rx                              : string  := "pma_8b_rx";
			hssi_rx_pld_pcs_interface_hd_8g_fifo_mode_rx                           : string  := "fifo_rx";
			hssi_rx_pld_pcs_interface_hd_g3_prot_mode                              : string  := "disabled_prot_mode";
			hssi_rx_pld_pcs_interface_hd_krfec_channel_operation_mode              : string  := "tx_rx_pair_enabled";
			hssi_rx_pld_pcs_interface_hd_krfec_lpbk_en                             : string  := "disable";
			hssi_rx_pld_pcs_interface_hd_krfec_prot_mode_rx                        : string  := "disabled_prot_mode_rx";
			hssi_rx_pld_pcs_interface_hd_krfec_low_latency_en_rx                   : string  := "disable";
			hssi_rx_pld_pcs_interface_hd_krfec_test_bus_mode                       : string  := "tx";
			hssi_rx_pld_pcs_interface_hd_pmaif_lpbk_en                             : string  := "disable";
			hssi_rx_pld_pcs_interface_hd_pmaif_channel_operation_mode              : string  := "tx_rx_pair_enabled";
			hssi_rx_pld_pcs_interface_hd_pmaif_sim_mode                            : string  := "disable";
			hssi_rx_pld_pcs_interface_hd_pmaif_prot_mode_rx                        : string  := "disabled_prot_mode_rx";
			hssi_rx_pld_pcs_interface_hd_pmaif_pma_dw_rx                           : string  := "pma_8b_rx";
			hssi_rx_pld_pcs_interface_hd_pldif_prot_mode_rx                        : string  := "disabled_prot_mode_rx";
			hssi_rx_pld_pcs_interface_hd_pldif_hrdrstctl_en                        : string  := "disable";
			hssi_rx_pld_pcs_interface_pcs_rx_block_sel                             : string  := "pcs_direct";
			hssi_rx_pld_pcs_interface_pcs_rx_clk_sel                               : string  := "pld_rx_clk";
			hssi_rx_pld_pcs_interface_pcs_rx_hip_clk_en                            : string  := "hip_rx_enable";
			hssi_rx_pld_pcs_interface_pcs_rx_output_sel                            : string  := "teng_output";
			hssi_rx_pld_pcs_interface_pcs_rx_clk_out_sel                           : string  := "teng_clk_out";
			hssi_common_pld_pcs_interface_dft_clk_out_en                           : string  := "dft_clk_out_disable";
			hssi_common_pld_pcs_interface_dft_clk_out_sel                          : string  := "teng_rx_dft_clk";
			hssi_common_pld_pcs_interface_hrdrstctrl_en                            : string  := "hrst_dis";
			hssi_common_pld_pcs_interface_pcs_testbus_block_sel                    : string  := "pma_if";
			hssi_rx_pcs_pma_interface_block_sel                                    : string  := "eight_g_pcs";
			hssi_rx_pcs_pma_interface_channel_operation_mode                       : string  := "tx_rx_pair_enabled";
			hssi_rx_pcs_pma_interface_clkslip_sel                                  : string  := "pld";
			hssi_rx_pcs_pma_interface_lpbk_en                                      : string  := "disable";
			hssi_rx_pcs_pma_interface_master_clk_sel                               : string  := "master_rx_pma_clk";
			hssi_rx_pcs_pma_interface_pldif_datawidth_mode                         : string  := "pldif_data_10bit";
			hssi_rx_pcs_pma_interface_pma_dw_rx                                    : string  := "pma_8b_rx";
			hssi_rx_pcs_pma_interface_pma_if_dft_en                                : string  := "dft_dis";
			hssi_rx_pcs_pma_interface_pma_if_dft_val                               : string  := "dft_0";
			hssi_rx_pcs_pma_interface_prbs_clken                                   : string  := "prbs_clk_dis";
			hssi_rx_pcs_pma_interface_prbs_ver                                     : string  := "prbs_off";
			hssi_rx_pcs_pma_interface_prbs9_dwidth                                 : string  := "prbs9_64b";
			hssi_rx_pcs_pma_interface_prot_mode_rx                                 : string  := "disabled_prot_mode_rx";
			hssi_rx_pcs_pma_interface_rx_dyn_polarity_inversion                    : string  := "rx_dyn_polinv_dis";
			hssi_rx_pcs_pma_interface_rx_lpbk_en                                   : string  := "lpbk_dis";
			hssi_rx_pcs_pma_interface_rx_prbs_force_signal_ok                      : string  := "unforce_sig_ok";
			hssi_rx_pcs_pma_interface_rx_prbs_mask                                 : string  := "prbsmask128";
			hssi_rx_pcs_pma_interface_rx_prbs_mode                                 : string  := "teng_mode";
			hssi_rx_pcs_pma_interface_rx_signalok_signaldet_sel                    : string  := "sel_sig_det";
			hssi_rx_pcs_pma_interface_rx_static_polarity_inversion                 : string  := "rx_stat_polinv_dis";
			hssi_rx_pcs_pma_interface_rx_uhsif_lpbk_en                             : string  := "uhsif_lpbk_dis";
			hssi_rx_pcs_pma_interface_sup_mode                                     : string  := "user_mode";
			hssi_tx_pcs_pma_interface_bypass_pma_txelecidle                        : string  := "false";
			hssi_tx_pcs_pma_interface_channel_operation_mode                       : string  := "tx_rx_pair_enabled";
			hssi_tx_pcs_pma_interface_lpbk_en                                      : string  := "disable";
			hssi_tx_pcs_pma_interface_master_clk_sel                               : string  := "master_tx_pma_clk";
			hssi_tx_pcs_pma_interface_pcie_sub_prot_mode_tx                        : string  := "other_prot_mode";
			hssi_tx_pcs_pma_interface_pldif_datawidth_mode                         : string  := "pldif_data_10bit";
			hssi_tx_pcs_pma_interface_pma_dw_tx                                    : string  := "pma_8b_tx";
			hssi_tx_pcs_pma_interface_pma_if_dft_en                                : string  := "dft_dis";
			hssi_tx_pcs_pma_interface_pmagate_en                                   : string  := "pmagate_dis";
			hssi_tx_pcs_pma_interface_prbs_clken                                   : string  := "prbs_clk_dis";
			hssi_tx_pcs_pma_interface_prbs_gen_pat                                 : string  := "prbs_gen_dis";
			hssi_tx_pcs_pma_interface_prbs9_dwidth                                 : string  := "prbs9_64b";
			hssi_tx_pcs_pma_interface_prot_mode_tx                                 : string  := "disabled_prot_mode_tx";
			hssi_tx_pcs_pma_interface_sq_wave_num                                  : string  := "sq_wave_4";
			hssi_tx_pcs_pma_interface_sqwgen_clken                                 : string  := "sqwgen_clk_dis";
			hssi_tx_pcs_pma_interface_sup_mode                                     : string  := "user_mode";
			hssi_tx_pcs_pma_interface_tx_dyn_polarity_inversion                    : string  := "tx_dyn_polinv_dis";
			hssi_tx_pcs_pma_interface_tx_pma_data_sel                              : string  := "pld_dir";
			hssi_tx_pcs_pma_interface_tx_static_polarity_inversion                 : string  := "tx_stat_polinv_dis";
			hssi_tx_pcs_pma_interface_uhsif_cnt_step_filt_before_lock              : string  := "uhsif_filt_stepsz_b4lock_4";
			hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_after_lock_value       : integer := 11;
			hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_before_lock            : string  := "uhsif_filt_cntthr_b4lock_16";
			hssi_tx_pcs_pma_interface_uhsif_dcn_test_update_period                 : string  := "uhsif_dcn_test_period_4";
			hssi_tx_pcs_pma_interface_uhsif_dcn_testmode_enable                    : string  := "uhsif_dcn_test_mode_disable";
			hssi_tx_pcs_pma_interface_uhsif_dead_zone_count_thresh                 : string  := "uhsif_dzt_cnt_thr_4";
			hssi_tx_pcs_pma_interface_uhsif_dead_zone_detection_enable             : string  := "uhsif_dzt_enable";
			hssi_tx_pcs_pma_interface_uhsif_dead_zone_obser_window                 : string  := "uhsif_dzt_obr_win_32";
			hssi_tx_pcs_pma_interface_uhsif_dead_zone_skip_size                    : string  := "uhsif_dzt_skipsz_8";
			hssi_tx_pcs_pma_interface_uhsif_delay_cell_index_sel                   : string  := "uhsif_index_internal";
			hssi_tx_pcs_pma_interface_uhsif_delay_cell_margin                      : string  := "uhsif_dcn_margin_4";
			hssi_tx_pcs_pma_interface_uhsif_delay_cell_static_index_value          : integer := 128;
			hssi_tx_pcs_pma_interface_uhsif_dft_dead_zone_control                  : string  := "uhsif_dft_dz_det_val_0";
			hssi_tx_pcs_pma_interface_uhsif_dft_up_filt_control                    : string  := "uhsif_dft_up_val_0";
			hssi_tx_pcs_pma_interface_uhsif_enable                                 : string  := "uhsif_disable";
			hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_after_lock              : string  := "uhsif_lkd_segsz_aflock_2048";
			hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_before_lock             : string  := "uhsif_lkd_segsz_b4lock_32";
			hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_after_lock_value   : integer := 8;
			hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_before_lock_value  : integer := 8;
			hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_after_lock_value  : integer := 3;
			hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_before_lock_value : integer := 3;
			hssi_common_pcs_pma_interface_asn_clk_enable                           : string  := "false";
			hssi_common_pcs_pma_interface_asn_enable                               : string  := "dis_asn";
			hssi_common_pcs_pma_interface_block_sel                                : string  := "eight_g_pcs";
			hssi_common_pcs_pma_interface_bypass_early_eios                        : string  := "false";
			hssi_common_pcs_pma_interface_bypass_pcie_switch                       : string  := "false";
			hssi_common_pcs_pma_interface_bypass_pma_ltr                           : string  := "false";
			hssi_common_pcs_pma_interface_bypass_pma_sw_done                       : string  := "false";
			hssi_common_pcs_pma_interface_bypass_ppm_lock                          : string  := "false";
			hssi_common_pcs_pma_interface_bypass_send_syncp_fbkp                   : string  := "false";
			hssi_common_pcs_pma_interface_bypass_txdetectrx                        : string  := "false";
			hssi_common_pcs_pma_interface_cdr_control                              : string  := "en_cdr_ctrl";
			hssi_common_pcs_pma_interface_cid_enable                               : string  := "en_cid_mode";
			hssi_common_pcs_pma_interface_data_mask_count                          : integer := 2500;
			hssi_common_pcs_pma_interface_data_mask_count_multi                    : integer := 1;
			hssi_common_pcs_pma_interface_dft_observation_clock_selection          : string  := "dft_clk_obsrv_tx0";
			hssi_common_pcs_pma_interface_early_eios_counter                       : integer := 50;
			hssi_common_pcs_pma_interface_force_freqdet                            : string  := "force_freqdet_dis";
			hssi_common_pcs_pma_interface_free_run_clk_enable                      : string  := "true";
			hssi_common_pcs_pma_interface_ignore_sigdet_g23                        : string  := "false";
			hssi_common_pcs_pma_interface_pc_en_counter                            : integer := 55;
			hssi_common_pcs_pma_interface_pc_rst_counter                           : integer := 23;
			hssi_common_pcs_pma_interface_pcie_hip_mode                            : string  := "hip_disable";
			hssi_common_pcs_pma_interface_ph_fifo_reg_mode                         : string  := "phfifo_reg_mode_dis";
			hssi_common_pcs_pma_interface_phfifo_flush_wait                        : integer := 36;
			hssi_common_pcs_pma_interface_pipe_if_g3pcs                            : string  := "pipe_if_8gpcs";
			hssi_common_pcs_pma_interface_pma_done_counter                         : integer := 175000;
			hssi_common_pcs_pma_interface_pma_if_dft_en                            : string  := "dft_dis";
			hssi_common_pcs_pma_interface_pma_if_dft_val                           : string  := "dft_0";
			hssi_common_pcs_pma_interface_ppm_cnt_rst                              : string  := "ppm_cnt_rst_dis";
			hssi_common_pcs_pma_interface_ppm_deassert_early                       : string  := "deassert_early_dis";
			hssi_common_pcs_pma_interface_ppm_gen1_2_cnt                           : string  := "cnt_32k";
			hssi_common_pcs_pma_interface_ppm_post_eidle_delay                     : string  := "cnt_200_cycles";
			hssi_common_pcs_pma_interface_ppmsel                                   : string  := "ppmsel_300";
			hssi_common_pcs_pma_interface_prot_mode                                : string  := "disable_prot_mode";
			hssi_common_pcs_pma_interface_rxvalid_mask                             : string  := "rxvalid_mask_en";
			hssi_common_pcs_pma_interface_sigdet_wait_counter                      : integer := 2500;
			hssi_common_pcs_pma_interface_sigdet_wait_counter_multi                : integer := 1;
			hssi_common_pcs_pma_interface_sim_mode                                 : string  := "disable";
			hssi_common_pcs_pma_interface_spd_chg_rst_wait_cnt_en                  : string  := "true";
			hssi_common_pcs_pma_interface_sup_mode                                 : string  := "user_mode";
			hssi_common_pcs_pma_interface_testout_sel                              : string  := "ppm_det_test";
			hssi_common_pcs_pma_interface_wait_clk_on_off_timer                    : integer := 4;
			hssi_common_pcs_pma_interface_wait_pipe_synchronizing                  : integer := 23;
			hssi_common_pcs_pma_interface_wait_send_syncp_fbkp                     : integer := 250;
			hssi_common_pcs_pma_interface_ppm_det_buckets                          : string  := "ppm_100_bucket";
			hssi_fifo_rx_pcs_double_read_mode                                      : string  := "double_read_dis";
			hssi_fifo_rx_pcs_prot_mode                                             : string  := "teng_mode";
			hssi_fifo_tx_pcs_double_write_mode                                     : string  := "double_write_dis";
			hssi_fifo_tx_pcs_prot_mode                                             : string  := "teng_mode";
			hssi_pipe_gen3_bypass_rx_detection_enable                              : string  := "false";
			hssi_pipe_gen3_bypass_rx_preset                                        : integer := 0;
			hssi_pipe_gen3_bypass_rx_preset_enable                                 : string  := "false";
			hssi_pipe_gen3_bypass_tx_coefficent                                    : integer := 0;
			hssi_pipe_gen3_bypass_tx_coefficent_enable                             : string  := "false";
			hssi_pipe_gen3_elecidle_delay_g3                                       : integer := 6;
			hssi_pipe_gen3_ind_error_reporting                                     : string  := "dis_ind_error_reporting";
			hssi_pipe_gen3_mode                                                    : string  := "pipe_g1";
			hssi_pipe_gen3_phy_status_delay_g12                                    : integer := 5;
			hssi_pipe_gen3_phy_status_delay_g3                                     : integer := 5;
			hssi_pipe_gen3_phystatus_rst_toggle_g12                                : string  := "dis_phystatus_rst_toggle";
			hssi_pipe_gen3_phystatus_rst_toggle_g3                                 : string  := "dis_phystatus_rst_toggle_g3";
			hssi_pipe_gen3_rate_match_pad_insertion                                : string  := "dis_rm_fifo_pad_ins";
			hssi_pipe_gen3_sup_mode                                                : string  := "user_mode";
			hssi_pipe_gen3_test_out_sel                                            : string  := "disable_test_out";
			hssi_pipe_gen1_2_elec_idle_delay_val                                   : integer := 0;
			hssi_pipe_gen1_2_error_replace_pad                                     : string  := "replace_edb";
			hssi_pipe_gen1_2_hip_mode                                              : string  := "dis_hip";
			hssi_pipe_gen1_2_ind_error_reporting                                   : string  := "dis_ind_error_reporting";
			hssi_pipe_gen1_2_phystatus_delay_val                                   : integer := 0;
			hssi_pipe_gen1_2_phystatus_rst_toggle                                  : string  := "dis_phystatus_rst_toggle";
			hssi_pipe_gen1_2_pipe_byte_de_serializer_en                            : string  := "dont_care_bds";
			hssi_pipe_gen1_2_prot_mode                                             : string  := "pipe_g1";
			hssi_pipe_gen1_2_rx_pipe_enable                                        : string  := "dis_pipe_rx";
			hssi_pipe_gen1_2_rxdetect_bypass                                       : string  := "dis_rxdetect_bypass";
			hssi_pipe_gen1_2_sup_mode                                              : string  := "user_mode";
			hssi_pipe_gen1_2_tx_pipe_enable                                        : string  := "dis_pipe_tx";
			hssi_pipe_gen1_2_txswing                                               : string  := "dis_txswing";
			pma_adapt_adp_1s_ctle_bypass                                           : string  := "radp_1s_ctle_bypass_0";
			pma_adapt_adp_4s_ctle_bypass                                           : string  := "radp_4s_ctle_bypass_0";
			pma_adapt_adp_ctle_en                                                  : string  := "radp_ctle_disable";
			pma_adapt_adp_dfe_fltap_bypass                                         : string  := "radp_dfe_fltap_bypass_0";
			pma_adapt_adp_dfe_fltap_en                                             : string  := "radp_dfe_fltap_disable";
			pma_adapt_adp_dfe_fxtap_bypass                                         : string  := "radp_dfe_fxtap_bypass_0";
			pma_adapt_adp_dfe_fxtap_en                                             : string  := "radp_dfe_fxtap_disable";
			pma_adapt_adp_dfe_fxtap_hold_en                                        : string  := "radp_dfe_fxtap_not_held";
			pma_adapt_adp_dfe_mode                                                 : string  := "radp_dfe_mode_0";
			pma_adapt_adp_vga_bypass                                               : string  := "radp_vga_bypass_0";
			pma_adapt_adp_vga_en                                                   : string  := "radp_vga_disable";
			pma_adapt_adp_vref_bypass                                              : string  := "radp_vref_bypass_0";
			pma_adapt_adp_vref_en                                                  : string  := "radp_vref_disable";
			pma_adapt_datarate                                                     : string  := "0 bps";
			pma_adapt_prot_mode                                                    : string  := "basic_rx";
			pma_adapt_sup_mode                                                     : string  := "user_mode";
			pma_adapt_adp_ctle_adapt_cycle_window                                  : string  := "radp_ctle_adapt_cycle_window_6";
			pma_adapt_odi_dfe_spec_en                                              : string  := "rodi_dfe_spec_en_0";
			pma_adapt_adapt_mode                                                   : string  := "dfe_vga";
			pma_adapt_adp_onetime_dfe                                              : string  := "radp_onetime_dfe_0";
			pma_adapt_adp_mode                                                     : string  := "radp_mode_0";
			pma_cdr_refclk_powerdown_mode                                          : string  := "powerup";
			pma_cdr_refclk_refclk_select                                           : string  := "ref_iqclk0";
			pma_cgb_bitslip_enable                                                 : string  := "enable_bitslip";
			pma_cgb_bonding_reset_enable                                           : string  := "disallow_bonding_reset";
			pma_cgb_datarate                                                       : string  := "0 bps";
			pma_cgb_pcie_gen3_bitwidth                                             : string  := "pciegen3_wide";
			pma_cgb_prot_mode                                                      : string  := "basic_tx";
			pma_cgb_ser_mode                                                       : string  := "eight_bit";
			pma_cgb_sup_mode                                                       : string  := "user_mode";
			pma_cgb_x1_div_m_sel                                                   : string  := "divbypass";
			pma_cgb_input_select_x1                                                : string  := "fpll_bot";
			pma_cgb_input_select_gen3                                              : string  := "unused";
			pma_cgb_input_select_xn                                                : string  := "unused";
			pma_cgb_tx_ucontrol_en                                                 : string  := "disable";
			pma_rx_dfe_datarate                                                    : string  := "0 bps";
			pma_rx_dfe_dft_en                                                      : string  := "dft_disable";
			pma_rx_dfe_pdb                                                         : string  := "dfe_enable";
			pma_rx_dfe_pdb_fixedtap                                                : string  := "fixtap_dfe_powerdown";
			pma_rx_dfe_pdb_floattap                                                : string  := "floattap_dfe_powerdown";
			pma_rx_dfe_pdb_fxtap4t7                                                : string  := "fxtap4t7_powerdown";
			pma_rx_dfe_sup_mode                                                    : string  := "user_mode";
			pma_rx_dfe_prot_mode                                                   : string  := "basic_rx";
			pma_rx_odi_datarate                                                    : string  := "0 bps";
			pma_rx_odi_sup_mode                                                    : string  := "user_mode";
			pma_rx_odi_step_ctrl_sel                                               : string  := "feedback_mode";
			pma_rx_odi_prot_mode                                                   : string  := "basic_rx";
			pma_rx_buf_bypass_eqz_stages_234                                       : string  := "bypass_off";
			pma_rx_buf_datarate                                                    : string  := "0 bps";
			pma_rx_buf_diag_lp_en                                                  : string  := "dlp_off";
			pma_rx_buf_prot_mode                                                   : string  := "basic_rx";
			pma_rx_buf_qpi_enable                                                  : string  := "non_qpi_mode";
			pma_rx_buf_rx_refclk_divider                                           : string  := "bypass_divider";
			pma_rx_buf_sup_mode                                                    : string  := "user_mode";
			pma_rx_buf_loopback_modes                                              : string  := "lpbk_disable";
			pma_rx_buf_refclk_en                                                   : string  := "enable";
			pma_rx_buf_pm_tx_rx_pcie_gen                                           : string  := "non_pcie";
			pma_rx_buf_pm_tx_rx_pcie_gen_bitwidth                                  : string  := "pcie_gen3_32b";
			pma_rx_buf_pm_tx_rx_cvp_mode                                           : string  := "cvp_off";
			pma_rx_buf_xrx_path_uc_cal_enable                                      : string  := "rx_cal_off";
			pma_rx_buf_xrx_path_sup_mode                                           : string  := "user_mode";
			pma_rx_buf_xrx_path_prot_mode                                          : string  := "unused";
			pma_rx_buf_xrx_path_datarate                                           : string  := "0 bps";
			pma_rx_buf_xrx_path_datawidth                                          : integer := 0;
			pma_rx_buf_xrx_path_pma_rx_divclk_hz                                   : string  := "0";
			pma_rx_sd_prot_mode                                                    : string  := "basic_rx";
			pma_rx_sd_sd_output_off                                                : integer := 1;
			pma_rx_sd_sd_output_on                                                 : integer := 1;
			pma_rx_sd_sd_pdb                                                       : string  := "sd_off";
			pma_rx_sd_sd_threshold                                                 : integer := 3;
			pma_rx_sd_sup_mode                                                     : string  := "user_mode";
			pma_tx_ser_ser_clk_divtx_user_sel                                      : string  := "divtx_user_33";
			pma_tx_ser_sup_mode                                                    : string  := "user_mode";
			pma_tx_ser_prot_mode                                                   : string  := "basic_tx";
			pma_tx_buf_datarate                                                    : string  := "0 bps";
			pma_tx_buf_prot_mode                                                   : string  := "basic_tx";
			pma_tx_buf_rx_det                                                      : string  := "mode_0";
			pma_tx_buf_rx_det_output_sel                                           : string  := "rx_det_pcie_out";
			pma_tx_buf_rx_det_pdb                                                  : string  := "rx_det_off";
			pma_tx_buf_sup_mode                                                    : string  := "user_mode";
			pma_tx_buf_user_fir_coeff_ctrl_sel                                     : string  := "ram_ctl";
			pma_tx_buf_xtx_path_prot_mode                                          : string  := "basic_tx";
			pma_tx_buf_xtx_path_datarate                                           : string  := "0 bps";
			pma_tx_buf_xtx_path_datawidth                                          : integer := 0;
			pma_tx_buf_xtx_path_clock_divider_ratio                                : integer := 0;
			pma_tx_buf_xtx_path_pma_tx_divclk_hz                                   : string  := "0";
			pma_tx_buf_xtx_path_tx_pll_clk_hz                                      : string  := "0 hz";
			pma_tx_buf_xtx_path_sup_mode                                           : string  := "user_mode";
			cdr_pll_pma_width                                                      : integer := 8;
			cdr_pll_cgb_div                                                        : integer := 1;
			cdr_pll_is_cascaded_pll                                                : string  := "false";
			cdr_pll_datarate                                                       : string  := "0 bps";
			cdr_pll_lpd_counter                                                    : integer := 1;
			cdr_pll_lpfd_counter                                                   : integer := 1;
			cdr_pll_n_counter_scratch                                              : integer := 1;
			cdr_pll_output_clock_frequency                                         : string  := "0 hz";
			cdr_pll_reference_clock_frequency                                      : string  := "0 hz";
			cdr_pll_set_cdr_vco_speed                                              : integer := 1;
			cdr_pll_set_cdr_vco_speed_fix                                          : integer := 0;
			cdr_pll_vco_freq                                                       : string  := "0 hz";
			cdr_pll_atb_select_control                                             : string  := "atb_off";
			cdr_pll_auto_reset_on                                                  : string  := "auto_reset_on";
			cdr_pll_bbpd_data_pattern_filter_select                                : string  := "bbpd_data_pat_off";
			cdr_pll_bw_sel                                                         : string  := "low";
			cdr_pll_cdr_odi_select                                                 : string  := "sel_cdr";
			cdr_pll_cdr_phaselock_mode                                             : string  := "no_ignore_lock";
			cdr_pll_cdr_powerdown_mode                                             : string  := "power_up";
			cdr_pll_chgpmp_current_pd                                              : string  := "cp_current_pd_setting0";
			cdr_pll_chgpmp_current_pfd                                             : string  := "cp_current_pfd_setting0";
			cdr_pll_chgpmp_replicate                                               : string  := "false";
			cdr_pll_chgpmp_testmode                                                : string  := "cp_test_disable";
			cdr_pll_clklow_mux_select                                              : string  := "clklow_mux_cdr_fbclk";
			cdr_pll_diag_loopback_enable                                           : string  := "false";
			cdr_pll_disable_up_dn                                                  : string  := "true";
			cdr_pll_fref_clklow_div                                                : integer := 1;
			cdr_pll_fref_mux_select                                                : string  := "fref_mux_cdr_refclk";
			cdr_pll_gpon_lck2ref_control                                           : string  := "gpon_lck2ref_off";
			cdr_pll_initial_settings                                               : string  := "true";
			cdr_pll_lck2ref_delay_control                                          : string  := "lck2ref_delay_off";
			cdr_pll_lf_resistor_pd                                                 : string  := "lf_pd_setting0";
			cdr_pll_lf_resistor_pfd                                                : string  := "lf_pfd_setting0";
			cdr_pll_lf_ripple_cap                                                  : string  := "lf_no_ripple";
			cdr_pll_loop_filter_bias_select                                        : string  := "lpflt_bias_off";
			cdr_pll_loopback_mode                                                  : string  := "loopback_disabled";
			cdr_pll_ltd_ltr_micro_controller_select                                : string  := "ltd_ltr_pcs";
			cdr_pll_m_counter                                                      : integer := 1;
			cdr_pll_n_counter                                                      : integer := 1;
			cdr_pll_pd_fastlock_mode                                               : string  := "false";
			cdr_pll_pd_l_counter                                                   : integer := 1;
			cdr_pll_pfd_l_counter                                                  : integer := 1;
			cdr_pll_primary_use                                                    : string  := "cdr";
			cdr_pll_prot_mode                                                      : string  := "unused";
			cdr_pll_reverse_serial_loopback                                        : string  := "no_loopback";
			cdr_pll_set_cdr_v2i_enable                                             : string  := "true";
			cdr_pll_set_cdr_vco_reset                                              : string  := "false";
			cdr_pll_set_cdr_vco_speed_pciegen3                                     : string  := "cdr_vco_max_speedbin_pciegen3";
			cdr_pll_sup_mode                                                       : string  := "user_mode";
			cdr_pll_tx_pll_prot_mode                                               : string  := "txpll_unused";
			cdr_pll_txpll_hclk_driver_enable                                       : string  := "false";
			cdr_pll_vco_overrange_voltage                                          : string  := "vco_overrange_off";
			cdr_pll_vco_underrange_voltage                                         : string  := "vco_underange_off";
			cdr_pll_fb_select                                                      : string  := "direct_fb";
			cdr_pll_uc_ro_cal                                                      : string  := "uc_ro_cal_off";
			cdr_pll_iqclk_mux_sel                                                  : string  := "power_down";
			cdr_pll_pcie_gen                                                       : string  := "non_pcie";
			cdr_pll_set_cdr_input_freq_range                                       : integer := 0;
			cdr_pll_chgpmp_current_dn_trim                                         : string  := "cp_current_trimming_dn_setting0";
			cdr_pll_chgpmp_up_pd_trim_double                                       : string  := "normal_up_trim_current";
			cdr_pll_chgpmp_current_up_pd                                           : string  := "cp_current_pd_up_setting0";
			cdr_pll_chgpmp_current_up_trim                                         : string  := "cp_current_trimming_up_setting0";
			cdr_pll_chgpmp_dn_pd_trim_double                                       : string  := "normal_dn_trim_current";
			cdr_pll_cal_vco_count_length                                           : string  := "sel_8b_count";
			cdr_pll_chgpmp_current_dn_pd                                           : string  := "cp_current_pd_dn_setting0";
			pma_rx_deser_clkdiv_source                                             : string  := "vco_bypass_normal";
			pma_rx_deser_clkdivrx_user_mode                                        : string  := "clkdivrx_user_disabled";
			pma_rx_deser_datarate                                                  : string  := "0 bps";
			pma_rx_deser_deser_factor                                              : integer := 8;
			pma_rx_deser_force_clkdiv_for_testing                                  : string  := "normal_clkdiv";
			pma_rx_deser_sdclk_enable                                              : string  := "false";
			pma_rx_deser_sup_mode                                                  : string  := "user_mode";
			pma_rx_deser_rst_n_adapt_odi                                           : string  := "no_rst_adapt_odi";
			pma_rx_deser_bitslip_bypass                                            : string  := "bs_bypass_no";
			pma_rx_deser_prot_mode                                                 : string  := "basic_rx";
			pma_rx_deser_pcie_gen                                                  : string  := "non_pcie";
			pma_rx_deser_pcie_gen_bitwidth                                         : string  := "pcie_gen3_32b"
		);
		port (
			tx_analogreset            : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- tx_analogreset
			tx_digitalreset           : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- tx_digitalreset
			rx_analogreset            : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- rx_analogreset
			rx_digitalreset           : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- rx_digitalreset
			tx_cal_busy               : out std_logic_vector(5 downto 0);                      -- tx_cal_busy
			rx_cal_busy               : out std_logic_vector(5 downto 0);                      -- rx_cal_busy
			tx_bonding_clocks         : in  std_logic_vector(35 downto 0)  := (others => 'X'); -- clk
			rx_cdr_refclk0            : in  std_logic                      := 'X';             -- clk
			tx_serial_data            : out std_logic_vector(5 downto 0);                      -- tx_serial_data
			rx_serial_data            : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- rx_serial_data
			rx_seriallpbken           : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- rx_seriallpbken
			rx_is_lockedtoref         : out std_logic_vector(5 downto 0);                      -- rx_is_lockedtoref
			rx_is_lockedtodata        : out std_logic_vector(5 downto 0);                      -- rx_is_lockedtodata
			tx_coreclkin              : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- clk
			rx_coreclkin              : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- clk
			tx_clkout                 : out std_logic_vector(5 downto 0);                      -- clk
			rx_clkout                 : out std_logic_vector(5 downto 0);                      -- clk
			tx_parallel_data          : in  std_logic_vector(767 downto 0) := (others => 'X'); -- unused_tx_parallel_data
			rx_parallel_data          : out std_logic_vector(767 downto 0);                    -- unused_rx_parallel_data
			tx_polinv                 : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- tx_polinv
			rx_polinv                 : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- rx_polinv
			reconfig_clk              : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- clk
			reconfig_reset            : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- reset
			reconfig_write            : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- write
			reconfig_read             : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- read
			reconfig_address          : in  std_logic_vector(12 downto 0)  := (others => 'X'); -- address
			reconfig_writedata        : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			reconfig_readdata         : out std_logic_vector(31 downto 0);                     -- readdata
			reconfig_waitrequest      : out std_logic_vector(0 downto 0);                      -- waitrequest
			tx_analogreset_ack        : out std_logic_vector(5 downto 0);                      -- tx_analogreset_ack
			rx_analogreset_ack        : out std_logic_vector(5 downto 0);                      -- rx_analogreset_ack
			tx_serial_clk0            : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- clk
			tx_serial_clk1            : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- clk
			tx_serial_clk2            : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- clk
			tx_serial_clk3            : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- clk
			tx_bonding_clocks1        : in  std_logic_vector(35 downto 0)  := (others => 'X'); -- clk
			tx_bonding_clocks2        : in  std_logic_vector(35 downto 0)  := (others => 'X'); -- clk
			tx_bonding_clocks3        : in  std_logic_vector(35 downto 0)  := (others => 'X'); -- clk
			rx_cdr_refclk1            : in  std_logic                      := 'X';             -- clk
			rx_cdr_refclk2            : in  std_logic                      := 'X';             -- clk
			rx_cdr_refclk3            : in  std_logic                      := 'X';             -- clk
			rx_cdr_refclk4            : in  std_logic                      := 'X';             -- clk
			rx_pma_clkslip            : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- rx_pma_clkslip
			rx_set_locktodata         : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- rx_set_locktodata
			rx_set_locktoref          : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- rx_set_locktoref
			rx_pma_qpipulldn          : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- rx_pma_qpipulldn
			tx_pma_qpipulldn          : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- tx_pma_qpipulldn
			tx_pma_qpipullup          : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- tx_pma_qpipullup
			tx_pma_txdetectrx         : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- tx_pma_txdetectrx
			tx_pma_elecidle           : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- tx_pma_elecidle
			tx_pma_rxfound            : out std_logic_vector(5 downto 0);                      -- tx_pma_rxfound
			rx_clklow                 : out std_logic_vector(5 downto 0);                      -- rx_clklow
			rx_fref                   : out std_logic_vector(5 downto 0);                      -- rx_fref
			tx_pma_clkout             : out std_logic_vector(5 downto 0);                      -- clk
			tx_pma_div_clkout         : out std_logic_vector(5 downto 0);                      -- clk
			tx_pma_iqtxrx_clkout      : out std_logic_vector(5 downto 0);                      -- clk
			rx_pma_clkout             : out std_logic_vector(5 downto 0);                      -- clk
			rx_pma_div_clkout         : out std_logic_vector(5 downto 0);                      -- clk
			rx_pma_iqtxrx_clkout      : out std_logic_vector(5 downto 0);                      -- clk
			tx_control                : in  std_logic_vector(107 downto 0) := (others => 'X'); -- tx_control
			rx_control                : out std_logic_vector(119 downto 0);                    -- rx_control
			rx_bitslip                : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- rx_bitslip
			rx_adapt_reset            : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- rx_adapt_reset
			rx_adapt_start            : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- rx_adapt_start
			rx_prbs_err_clr           : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- rx_prbs_err_clr
			rx_prbs_done              : out std_logic_vector(5 downto 0);                      -- rx_prbs_done
			rx_prbs_err               : out std_logic_vector(5 downto 0);                      -- rx_prbs_err
			tx_uhsif_clk              : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- clk
			tx_uhsif_clkout           : out std_logic_vector(5 downto 0);                      -- clk
			tx_uhsif_lock             : out std_logic_vector(5 downto 0);                      -- tx_uhsif_lock
			tx_std_pcfifo_full        : out std_logic_vector(5 downto 0);                      -- tx_std_pcfifo_full
			tx_std_pcfifo_empty       : out std_logic_vector(5 downto 0);                      -- tx_std_pcfifo_empty
			rx_std_pcfifo_full        : out std_logic_vector(5 downto 0);                      -- rx_std_pcfifo_full
			rx_std_pcfifo_empty       : out std_logic_vector(5 downto 0);                      -- rx_std_pcfifo_empty
			rx_std_bitrev_ena         : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- rx_std_bitrev_ena
			rx_std_byterev_ena        : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- rx_std_byterev_ena
			tx_std_bitslipboundarysel : in  std_logic_vector(29 downto 0)  := (others => 'X'); -- tx_std_bitslipboundarysel
			rx_std_bitslipboundarysel : out std_logic_vector(29 downto 0);                     -- rx_std_bitslipboundarysel
			rx_std_wa_patternalign    : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- rx_std_wa_patternalign
			rx_std_wa_a1a2size        : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- rx_std_wa_a1a2size
			rx_std_rmfifo_full        : out std_logic_vector(5 downto 0);                      -- rx_std_rmfifo_full
			rx_std_rmfifo_empty       : out std_logic_vector(5 downto 0);                      -- rx_std_rmfifo_empty
			rx_std_signaldetect       : out std_logic_vector(5 downto 0);                      -- rx_std_signaldetect
			tx_enh_data_valid         : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- tx_enh_data_valid
			tx_enh_fifo_full          : out std_logic_vector(5 downto 0);                      -- tx_enh_fifo_full
			tx_enh_fifo_pfull         : out std_logic_vector(5 downto 0);                      -- tx_enh_fifo_pfull
			tx_enh_fifo_empty         : out std_logic_vector(5 downto 0);                      -- tx_enh_fifo_empty
			tx_enh_fifo_pempty        : out std_logic_vector(5 downto 0);                      -- tx_enh_fifo_pempty
			tx_enh_fifo_cnt           : out std_logic_vector(23 downto 0);                     -- tx_enh_fifo_cnt
			rx_enh_fifo_rd_en         : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- rx_enh_fifo_rd_en
			rx_enh_data_valid         : out std_logic_vector(5 downto 0);                      -- rx_enh_data_valid
			rx_enh_fifo_full          : out std_logic_vector(5 downto 0);                      -- rx_enh_fifo_full
			rx_enh_fifo_pfull         : out std_logic_vector(5 downto 0);                      -- rx_enh_fifo_pfull
			rx_enh_fifo_empty         : out std_logic_vector(5 downto 0);                      -- rx_enh_fifo_empty
			rx_enh_fifo_pempty        : out std_logic_vector(5 downto 0);                      -- rx_enh_fifo_pempty
			rx_enh_fifo_del           : out std_logic_vector(5 downto 0);                      -- rx_enh_fifo_del
			rx_enh_fifo_insert        : out std_logic_vector(5 downto 0);                      -- rx_enh_fifo_insert
			rx_enh_fifo_cnt           : out std_logic_vector(29 downto 0);                     -- rx_enh_fifo_cnt
			rx_enh_fifo_align_val     : out std_logic_vector(5 downto 0);                      -- rx_enh_fifo_align_val
			rx_enh_fifo_align_clr     : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- rx_enh_fifo_align_clr
			tx_enh_frame              : out std_logic_vector(5 downto 0);                      -- tx_enh_frame
			tx_enh_frame_burst_en     : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- tx_enh_frame_burst_en
			tx_enh_frame_diag_status  : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- tx_enh_frame_diag_status
			rx_enh_frame              : out std_logic_vector(5 downto 0);                      -- rx_enh_frame
			rx_enh_frame_lock         : out std_logic_vector(5 downto 0);                      -- rx_enh_frame_lock
			rx_enh_frame_diag_status  : out std_logic_vector(11 downto 0);                     -- rx_enh_frame_diag_status
			rx_enh_crc32_err          : out std_logic_vector(5 downto 0);                      -- rx_enh_crc32err
			rx_enh_highber            : out std_logic_vector(5 downto 0);                      -- rx_enh_highber
			rx_enh_highber_clr_cnt    : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- rx_enh_highber_clr_cnt
			rx_enh_clr_errblk_count   : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- rx_enh_clr_errblk_count
			rx_enh_blk_lock           : out std_logic_vector(5 downto 0);                      -- rx_enh_blk_lock
			tx_enh_bitslip            : in  std_logic_vector(41 downto 0)  := (others => 'X'); -- tx_enh_bitslip
			tx_hip_data               : in  std_logic_vector(383 downto 0) := (others => 'X'); -- tx_hip_data
			rx_hip_data               : out std_logic_vector(305 downto 0);                    -- rx_hip_data
			hip_pipe_pclk             : out std_logic;                                         -- hip_pipe_pclk
			hip_fixedclk              : out std_logic;                                         -- hip_fixedclk
			hip_frefclk               : out std_logic_vector(5 downto 0);                      -- hip_frefclk
			hip_ctrl                  : out std_logic_vector(47 downto 0);                     -- hip_ctrl
			hip_cal_done              : out std_logic_vector(5 downto 0);                      -- hip_cal_done
			pipe_rate                 : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- pipe_rate
			pipe_sw_done              : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- pipe_sw_done
			pipe_sw                   : out std_logic_vector(1 downto 0);                      -- pipe_sw
			pipe_hclk_in              : in  std_logic                      := 'X';             -- clk
			pipe_hclk_out             : out std_logic;                                         -- clk
			pipe_g3_txdeemph          : in  std_logic_vector(107 downto 0) := (others => 'X'); -- pipe_g3_txdeemph
			pipe_g3_rxpresethint      : in  std_logic_vector(17 downto 0)  := (others => 'X'); -- pipe_g3_rxpresethint
			pipe_rx_eidleinfersel     : in  std_logic_vector(17 downto 0)  := (others => 'X'); -- pipe_rx_eidleinfersel
			pipe_rx_elecidle          : out std_logic_vector(5 downto 0);                      -- pipe_rx_elecidle
			pipe_rx_polarity          : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- pipe_rx_polarity
			avmm_busy                 : out std_logic_vector(5 downto 0)                       -- avmm_busy
		);
	end component gx_std_x6_altera_xcvr_native_a10_151_eh2glbi;

	signal xcvr_native_a10_0_rx_parallel_data : std_logic_vector(767 downto 0); -- port fragment

	for xcvr_native_a10_0 : gx_std_x6_altera_xcvr_native_a10_151_eh2glbi
		use entity gx_std_x6_altera_xcvr_native_a10_151.gx_std_x6_altera_xcvr_native_a10_151_eh2glbi;
begin

	xcvr_native_a10_0 : component gx_std_x6_altera_xcvr_native_a10_151_eh2glbi
		generic map (
			device_revision                                                        => "20nm5",
			duplex_mode                                                            => "duplex",
			channels                                                               => 6,
			enable_calibration                                                     => 1,
			enable_analog_resets                                                   => 1,
			enable_reset_sequence                                                  => 1,
			bonded_mode                                                            => "pma_pcs",
			pcs_bonding_master                                                     => 3,
			plls                                                                   => 1,
			number_physical_bonding_clocks                                         => 1,
			cdr_refclk_cnt                                                         => 1,
			enable_hip                                                             => 0,
			hip_cal_en                                                             => "disable",
			rcfg_enable                                                            => 1,
			rcfg_shared                                                            => 1,
			rcfg_jtag_enable                                                       => 1,
			rcfg_separate_avmm_busy                                                => 0,
			adme_prot_mode                                                         => "basic_std",
			adme_data_rate                                                         => "4800000000",
			dbg_embedded_debug_enable                                              => 1,
			dbg_capability_reg_enable                                              => 1,
			dbg_user_identifier                                                    => 0,
			dbg_stat_soft_logic_enable                                             => 1,
			dbg_ctrl_soft_logic_enable                                             => 1,
			dbg_prbs_soft_logic_enable                                             => 1,
			dbg_odi_soft_logic_enable                                              => 1,
			rcfg_emb_strm_enable                                                   => 0,
			rcfg_profile_cnt                                                       => 2,
			hssi_gen3_rx_pcs_block_sync                                            => "bypass_block_sync",
			hssi_gen3_rx_pcs_block_sync_sm                                         => "disable_blk_sync_sm",
			hssi_gen3_rx_pcs_cdr_ctrl_force_unalgn                                 => "disable",
			hssi_gen3_rx_pcs_lpbk_force                                            => "lpbk_frce_dis",
			hssi_gen3_rx_pcs_mode                                                  => "disable_pcs",
			hssi_gen3_rx_pcs_rate_match_fifo                                       => "bypass_rm_fifo",
			hssi_gen3_rx_pcs_rate_match_fifo_latency                               => "low_latency",
			hssi_gen3_rx_pcs_reverse_lpbk                                          => "rev_lpbk_dis",
			hssi_gen3_rx_pcs_rx_b4gb_par_lpbk                                      => "b4gb_par_lpbk_dis",
			hssi_gen3_rx_pcs_rx_force_balign                                       => "dis_force_balign",
			hssi_gen3_rx_pcs_rx_ins_del_one_skip                                   => "ins_del_one_skip_dis",
			hssi_gen3_rx_pcs_rx_num_fixed_pat                                      => 0,
			hssi_gen3_rx_pcs_rx_test_out_sel                                       => "rx_test_out0",
			hssi_gen3_rx_pcs_sup_mode                                              => "user_mode",
			hssi_gen3_tx_pcs_mode                                                  => "disable_pcs",
			hssi_gen3_tx_pcs_reverse_lpbk                                          => "rev_lpbk_dis",
			hssi_gen3_tx_pcs_sup_mode                                              => "user_mode",
			hssi_gen3_tx_pcs_tx_bitslip                                            => 0,
			hssi_gen3_tx_pcs_tx_gbox_byp                                           => "bypass_gbox",
			hssi_krfec_rx_pcs_blksync_cor_en                                       => "detect",
			hssi_krfec_rx_pcs_bypass_gb                                            => "bypass_dis",
			hssi_krfec_rx_pcs_clr_ctrl                                             => "both_enabled",
			hssi_krfec_rx_pcs_ctrl_bit_reverse                                     => "ctrl_bit_reverse_en",
			hssi_krfec_rx_pcs_data_bit_reverse                                     => "data_bit_reverse_dis",
			hssi_krfec_rx_pcs_dv_start                                             => "with_blklock",
			hssi_krfec_rx_pcs_err_mark_type                                        => "err_mark_10g",
			hssi_krfec_rx_pcs_error_marking_en                                     => "err_mark_dis",
			hssi_krfec_rx_pcs_low_latency_en                                       => "disable",
			hssi_krfec_rx_pcs_lpbk_mode                                            => "lpbk_dis",
			hssi_krfec_rx_pcs_parity_invalid_enum                                  => 8,
			hssi_krfec_rx_pcs_parity_valid_num                                     => 4,
			hssi_krfec_rx_pcs_pipeln_blksync                                       => "enable",
			hssi_krfec_rx_pcs_pipeln_descrm                                        => "disable",
			hssi_krfec_rx_pcs_pipeln_errcorrect                                    => "disable",
			hssi_krfec_rx_pcs_pipeln_errtrap_ind                                   => "enable",
			hssi_krfec_rx_pcs_pipeln_errtrap_lfsr                                  => "disable",
			hssi_krfec_rx_pcs_pipeln_errtrap_loc                                   => "disable",
			hssi_krfec_rx_pcs_pipeln_errtrap_pat                                   => "disable",
			hssi_krfec_rx_pcs_pipeln_gearbox                                       => "enable",
			hssi_krfec_rx_pcs_pipeln_syndrm                                        => "enable",
			hssi_krfec_rx_pcs_pipeln_trans_dec                                     => "disable",
			hssi_krfec_rx_pcs_prot_mode                                            => "disable_mode",
			hssi_krfec_rx_pcs_receive_order                                        => "receive_lsb",
			hssi_krfec_rx_pcs_rx_testbus_sel                                       => "overall",
			hssi_krfec_rx_pcs_signal_ok_en                                         => "sig_ok_en",
			hssi_krfec_rx_pcs_sup_mode                                             => "user_mode",
			hssi_krfec_tx_pcs_burst_err                                            => "burst_err_dis",
			hssi_krfec_tx_pcs_burst_err_len                                        => "burst_err_len1",
			hssi_krfec_tx_pcs_ctrl_bit_reverse                                     => "ctrl_bit_reverse_en",
			hssi_krfec_tx_pcs_data_bit_reverse                                     => "data_bit_reverse_dis",
			hssi_krfec_tx_pcs_enc_frame_query                                      => "enc_query_dis",
			hssi_krfec_tx_pcs_low_latency_en                                       => "disable",
			hssi_krfec_tx_pcs_pipeln_encoder                                       => "enable",
			hssi_krfec_tx_pcs_pipeln_scrambler                                     => "enable",
			hssi_krfec_tx_pcs_prot_mode                                            => "disable_mode",
			hssi_krfec_tx_pcs_sup_mode                                             => "user_mode",
			hssi_krfec_tx_pcs_transcode_err                                        => "trans_err_dis",
			hssi_krfec_tx_pcs_transmit_order                                       => "transmit_lsb",
			hssi_krfec_tx_pcs_tx_testbus_sel                                       => "overall",
			hssi_10g_rx_pcs_align_del                                              => "align_del_dis",
			hssi_10g_rx_pcs_ber_bit_err_total_cnt                                  => "bit_err_total_cnt_10g",
			hssi_10g_rx_pcs_ber_clken                                              => "ber_clk_dis",
			hssi_10g_rx_pcs_ber_xus_timer_window                                   => 19530,
			hssi_10g_rx_pcs_bitslip_mode                                           => "bitslip_dis",
			hssi_10g_rx_pcs_blksync_bitslip_type                                   => "bitslip_comb",
			hssi_10g_rx_pcs_blksync_bitslip_wait_cnt                               => 1,
			hssi_10g_rx_pcs_blksync_bitslip_wait_type                              => "bitslip_cnt",
			hssi_10g_rx_pcs_blksync_bypass                                         => "blksync_bypass_en",
			hssi_10g_rx_pcs_blksync_clken                                          => "blksync_clk_dis",
			hssi_10g_rx_pcs_blksync_enum_invalid_sh_cnt                            => "enum_invalid_sh_cnt_10g",
			hssi_10g_rx_pcs_blksync_knum_sh_cnt_postlock                           => "knum_sh_cnt_postlock_10g",
			hssi_10g_rx_pcs_blksync_knum_sh_cnt_prelock                            => "knum_sh_cnt_prelock_10g",
			hssi_10g_rx_pcs_blksync_pipeln                                         => "blksync_pipeln_dis",
			hssi_10g_rx_pcs_clr_errblk_cnt_en                                      => "disable",
			hssi_10g_rx_pcs_control_del                                            => "control_del_none",
			hssi_10g_rx_pcs_crcchk_bypass                                          => "crcchk_bypass_en",
			hssi_10g_rx_pcs_crcchk_clken                                           => "crcchk_clk_dis",
			hssi_10g_rx_pcs_crcchk_inv                                             => "crcchk_inv_en",
			hssi_10g_rx_pcs_crcchk_pipeln                                          => "crcchk_pipeln_en",
			hssi_10g_rx_pcs_crcflag_pipeln                                         => "crcflag_pipeln_en",
			hssi_10g_rx_pcs_ctrl_bit_reverse                                       => "ctrl_bit_reverse_dis",
			hssi_10g_rx_pcs_data_bit_reverse                                       => "data_bit_reverse_dis",
			hssi_10g_rx_pcs_dec_64b66b_rxsm_bypass                                 => "dec_64b66b_rxsm_bypass_en",
			hssi_10g_rx_pcs_dec64b66b_clken                                        => "dec64b66b_clk_dis",
			hssi_10g_rx_pcs_descrm_bypass                                          => "descrm_bypass_en",
			hssi_10g_rx_pcs_descrm_clken                                           => "descrm_clk_dis",
			hssi_10g_rx_pcs_descrm_mode                                            => "async",
			hssi_10g_rx_pcs_descrm_pipeln                                          => "enable",
			hssi_10g_rx_pcs_dft_clk_out_sel                                        => "rx_master_clk",
			hssi_10g_rx_pcs_dis_signal_ok                                          => "dis_signal_ok_en",
			hssi_10g_rx_pcs_dispchk_bypass                                         => "dispchk_bypass_en",
			hssi_10g_rx_pcs_empty_flag_type                                        => "empty_rd_side",
			hssi_10g_rx_pcs_fast_path                                              => "fast_path_en",
			hssi_10g_rx_pcs_fec_clken                                              => "fec_clk_dis",
			hssi_10g_rx_pcs_fec_enable                                             => "fec_dis",
			hssi_10g_rx_pcs_fifo_double_read                                       => "fifo_double_read_dis",
			hssi_10g_rx_pcs_fifo_stop_rd                                           => "n_rd_empty",
			hssi_10g_rx_pcs_fifo_stop_wr                                           => "n_wr_full",
			hssi_10g_rx_pcs_force_align                                            => "force_align_dis",
			hssi_10g_rx_pcs_frmsync_bypass                                         => "frmsync_bypass_en",
			hssi_10g_rx_pcs_frmsync_clken                                          => "frmsync_clk_dis",
			hssi_10g_rx_pcs_frmsync_enum_scrm                                      => "enum_scrm_default",
			hssi_10g_rx_pcs_frmsync_enum_sync                                      => "enum_sync_default",
			hssi_10g_rx_pcs_frmsync_flag_type                                      => "location_only",
			hssi_10g_rx_pcs_frmsync_knum_sync                                      => "knum_sync_default",
			hssi_10g_rx_pcs_frmsync_mfrm_length                                    => 2048,
			hssi_10g_rx_pcs_frmsync_pipeln                                         => "frmsync_pipeln_en",
			hssi_10g_rx_pcs_full_flag_type                                         => "full_wr_side",
			hssi_10g_rx_pcs_gb_rx_idwidth                                          => "width_64",
			hssi_10g_rx_pcs_gb_rx_odwidth                                          => "width_64",
			hssi_10g_rx_pcs_gbexp_clken                                            => "gbexp_clk_dis",
			hssi_10g_rx_pcs_low_latency_en                                         => "disable",
			hssi_10g_rx_pcs_lpbk_mode                                              => "lpbk_dis",
			hssi_10g_rx_pcs_master_clk_sel                                         => "master_rx_pma_clk",
			hssi_10g_rx_pcs_pempty_flag_type                                       => "pempty_rd_side",
			hssi_10g_rx_pcs_pfull_flag_type                                        => "pfull_wr_side",
			hssi_10g_rx_pcs_phcomp_rd_del                                          => "phcomp_rd_del2",
			hssi_10g_rx_pcs_pld_if_type                                            => "fifo",
			hssi_10g_rx_pcs_prot_mode                                              => "disable_mode",
			hssi_10g_rx_pcs_rand_clken                                             => "rand_clk_dis",
			hssi_10g_rx_pcs_rd_clk_sel                                             => "rd_rx_pld_clk",
			hssi_10g_rx_pcs_rdfifo_clken                                           => "rdfifo_clk_dis",
			hssi_10g_rx_pcs_rx_fifo_write_ctrl                                     => "blklock_stops",
			hssi_10g_rx_pcs_rx_scrm_width                                          => "bit64",
			hssi_10g_rx_pcs_rx_sh_location                                         => "msb",
			hssi_10g_rx_pcs_rx_signal_ok_sel                                       => "synchronized_ver",
			hssi_10g_rx_pcs_rx_sm_bypass                                           => "rx_sm_bypass_en",
			hssi_10g_rx_pcs_rx_sm_hiber                                            => "rx_sm_hiber_en",
			hssi_10g_rx_pcs_rx_sm_pipeln                                           => "rx_sm_pipeln_en",
			hssi_10g_rx_pcs_rx_testbus_sel                                         => "rx_fifo_testbus1",
			hssi_10g_rx_pcs_rx_true_b2b                                            => "b2b",
			hssi_10g_rx_pcs_rxfifo_empty                                           => "empty_default",
			hssi_10g_rx_pcs_rxfifo_full                                            => "full_default",
			hssi_10g_rx_pcs_rxfifo_mode                                            => "phase_comp",
			hssi_10g_rx_pcs_rxfifo_pempty                                          => 2,
			hssi_10g_rx_pcs_rxfifo_pfull                                           => 23,
			hssi_10g_rx_pcs_stretch_num_stages                                     => "zero_stage",
			hssi_10g_rx_pcs_sup_mode                                               => "user_mode",
			hssi_10g_rx_pcs_test_mode                                              => "test_off",
			hssi_10g_rx_pcs_wrfifo_clken                                           => "wrfifo_clk_dis",
			hssi_10g_rx_pcs_advanced_user_mode                                     => "disable",
			hssi_10g_tx_pcs_bitslip_en                                             => "bitslip_dis",
			hssi_10g_tx_pcs_bonding_dft_en                                         => "dft_dis",
			hssi_10g_tx_pcs_bonding_dft_val                                        => "dft_0",
			hssi_10g_tx_pcs_crcgen_bypass                                          => "crcgen_bypass_en",
			hssi_10g_tx_pcs_crcgen_clken                                           => "crcgen_clk_dis",
			hssi_10g_tx_pcs_crcgen_err                                             => "crcgen_err_dis",
			hssi_10g_tx_pcs_crcgen_inv                                             => "crcgen_inv_en",
			hssi_10g_tx_pcs_ctrl_bit_reverse                                       => "ctrl_bit_reverse_dis",
			hssi_10g_tx_pcs_data_bit_reverse                                       => "data_bit_reverse_dis",
			hssi_10g_tx_pcs_dft_clk_out_sel                                        => "tx_master_clk",
			hssi_10g_tx_pcs_dispgen_bypass                                         => "dispgen_bypass_en",
			hssi_10g_tx_pcs_dispgen_clken                                          => "dispgen_clk_dis",
			hssi_10g_tx_pcs_dispgen_err                                            => "dispgen_err_dis",
			hssi_10g_tx_pcs_dispgen_pipeln                                         => "dispgen_pipeln_dis",
			hssi_10g_tx_pcs_empty_flag_type                                        => "empty_rd_side",
			hssi_10g_tx_pcs_enc_64b66b_txsm_bypass                                 => "enc_64b66b_txsm_bypass_en",
			hssi_10g_tx_pcs_enc64b66b_txsm_clken                                   => "enc64b66b_txsm_clk_dis",
			hssi_10g_tx_pcs_fastpath                                               => "fastpath_en",
			hssi_10g_tx_pcs_fec_clken                                              => "fec_clk_dis",
			hssi_10g_tx_pcs_fec_enable                                             => "fec_dis",
			hssi_10g_tx_pcs_fifo_double_write                                      => "fifo_double_write_dis",
			hssi_10g_tx_pcs_fifo_reg_fast                                          => "fifo_reg_fast_dis",
			hssi_10g_tx_pcs_fifo_stop_rd                                           => "rd_empty",
			hssi_10g_tx_pcs_fifo_stop_wr                                           => "n_wr_full",
			hssi_10g_tx_pcs_frmgen_burst                                           => "frmgen_burst_dis",
			hssi_10g_tx_pcs_frmgen_bypass                                          => "frmgen_bypass_en",
			hssi_10g_tx_pcs_frmgen_clken                                           => "frmgen_clk_dis",
			hssi_10g_tx_pcs_frmgen_mfrm_length                                     => 2048,
			hssi_10g_tx_pcs_frmgen_pipeln                                          => "frmgen_pipeln_en",
			hssi_10g_tx_pcs_frmgen_pyld_ins                                        => "frmgen_pyld_ins_dis",
			hssi_10g_tx_pcs_frmgen_wordslip                                        => "frmgen_wordslip_dis",
			hssi_10g_tx_pcs_full_flag_type                                         => "full_wr_side",
			hssi_10g_tx_pcs_gb_pipeln_bypass                                       => "disable",
			hssi_10g_tx_pcs_gb_tx_idwidth                                          => "width_64",
			hssi_10g_tx_pcs_gb_tx_odwidth                                          => "width_64",
			hssi_10g_tx_pcs_gbred_clken                                            => "gbred_clk_dis",
			hssi_10g_tx_pcs_low_latency_en                                         => "disable",
			hssi_10g_tx_pcs_master_clk_sel                                         => "master_tx_pma_clk",
			hssi_10g_tx_pcs_pempty_flag_type                                       => "pempty_rd_side",
			hssi_10g_tx_pcs_pfull_flag_type                                        => "pfull_wr_side",
			hssi_10g_tx_pcs_phcomp_rd_del                                          => "phcomp_rd_del2",
			hssi_10g_tx_pcs_pld_if_type                                            => "fifo",
			hssi_10g_tx_pcs_prot_mode                                              => "disable_mode",
			hssi_10g_tx_pcs_pseudo_random                                          => "all_0",
			hssi_10g_tx_pcs_pseudo_seed_a                                          => "288230376151711743",
			hssi_10g_tx_pcs_pseudo_seed_b                                          => "288230376151711743",
			hssi_10g_tx_pcs_random_disp                                            => "disable",
			hssi_10g_tx_pcs_rdfifo_clken                                           => "rdfifo_clk_dis",
			hssi_10g_tx_pcs_scrm_bypass                                            => "scrm_bypass_en",
			hssi_10g_tx_pcs_scrm_clken                                             => "scrm_clk_dis",
			hssi_10g_tx_pcs_scrm_mode                                              => "async",
			hssi_10g_tx_pcs_scrm_pipeln                                            => "enable",
			hssi_10g_tx_pcs_sh_err                                                 => "sh_err_dis",
			hssi_10g_tx_pcs_sop_mark                                               => "sop_mark_dis",
			hssi_10g_tx_pcs_stretch_num_stages                                     => "zero_stage",
			hssi_10g_tx_pcs_sup_mode                                               => "user_mode",
			hssi_10g_tx_pcs_test_mode                                              => "test_off",
			hssi_10g_tx_pcs_tx_scrm_err                                            => "scrm_err_dis",
			hssi_10g_tx_pcs_tx_scrm_width                                          => "bit64",
			hssi_10g_tx_pcs_tx_sh_location                                         => "msb",
			hssi_10g_tx_pcs_tx_sm_bypass                                           => "tx_sm_bypass_en",
			hssi_10g_tx_pcs_tx_sm_pipeln                                           => "tx_sm_pipeln_en",
			hssi_10g_tx_pcs_tx_testbus_sel                                         => "tx_fifo_testbus1",
			hssi_10g_tx_pcs_txfifo_empty                                           => "empty_default",
			hssi_10g_tx_pcs_txfifo_full                                            => "full_default",
			hssi_10g_tx_pcs_txfifo_mode                                            => "phase_comp",
			hssi_10g_tx_pcs_txfifo_pempty                                          => 2,
			hssi_10g_tx_pcs_txfifo_pfull                                           => 11,
			hssi_10g_tx_pcs_wr_clk_sel                                             => "wr_tx_pld_clk",
			hssi_10g_tx_pcs_wrfifo_clken                                           => "wrfifo_clk_dis",
			hssi_10g_tx_pcs_advanced_user_mode                                     => "disable",
			hssi_8g_rx_pcs_auto_error_replacement                                  => "dis_err_replace",
			hssi_8g_rx_pcs_bit_reversal                                            => "dis_bit_reversal",
			hssi_8g_rx_pcs_bonding_dft_en                                          => "dft_dis",
			hssi_8g_rx_pcs_bonding_dft_val                                         => "dft_0",
			hssi_8g_rx_pcs_bypass_pipeline_reg                                     => "dis_bypass_pipeline",
			hssi_8g_rx_pcs_byte_deserializer                                       => "dis_bds",
			hssi_8g_rx_pcs_cdr_ctrl_rxvalid_mask                                   => "dis_rxvalid_mask",
			hssi_8g_rx_pcs_clkcmp_pattern_n                                        => 0,
			hssi_8g_rx_pcs_clkcmp_pattern_p                                        => 0,
			hssi_8g_rx_pcs_clock_gate_bds_dec_asn                                  => "dis_bds_dec_asn_clk_gating",
			hssi_8g_rx_pcs_clock_gate_cdr_eidle                                    => "en_cdr_eidle_clk_gating",
			hssi_8g_rx_pcs_clock_gate_dw_pc_wrclk                                  => "dis_dw_pc_wrclk_gating",
			hssi_8g_rx_pcs_clock_gate_dw_rm_rd                                     => "en_dw_rm_rdclk_gating",
			hssi_8g_rx_pcs_clock_gate_dw_rm_wr                                     => "en_dw_rm_wrclk_gating",
			hssi_8g_rx_pcs_clock_gate_dw_wa                                        => "dis_dw_wa_clk_gating",
			hssi_8g_rx_pcs_clock_gate_pc_rdclk                                     => "dis_pc_rdclk_gating",
			hssi_8g_rx_pcs_clock_gate_sw_pc_wrclk                                  => "dis_sw_pc_wrclk_gating",
			hssi_8g_rx_pcs_clock_gate_sw_rm_rd                                     => "en_sw_rm_rdclk_gating",
			hssi_8g_rx_pcs_clock_gate_sw_rm_wr                                     => "en_sw_rm_wrclk_gating",
			hssi_8g_rx_pcs_clock_gate_sw_wa                                        => "dis_sw_wa_clk_gating",
			hssi_8g_rx_pcs_clock_observation_in_pld_core                           => "internal_sw_wa_clk",
			hssi_8g_rx_pcs_eidle_entry_eios                                        => "dis_eidle_eios",
			hssi_8g_rx_pcs_eidle_entry_iei                                         => "dis_eidle_iei",
			hssi_8g_rx_pcs_eidle_entry_sd                                          => "dis_eidle_sd",
			hssi_8g_rx_pcs_eightb_tenb_decoder                                     => "dis_8b10b",
			hssi_8g_rx_pcs_err_flags_sel                                           => "err_flags_wa",
			hssi_8g_rx_pcs_fixed_pat_det                                           => "dis_fixed_patdet",
			hssi_8g_rx_pcs_fixed_pat_num                                           => 0,
			hssi_8g_rx_pcs_force_signal_detect                                     => "en_force_signal_detect",
			hssi_8g_rx_pcs_gen3_clk_en                                             => "disable_clk",
			hssi_8g_rx_pcs_gen3_rx_clk_sel                                         => "rcvd_clk",
			hssi_8g_rx_pcs_gen3_tx_clk_sel                                         => "tx_pma_clk",
			hssi_8g_rx_pcs_hip_mode                                                => "dis_hip",
			hssi_8g_rx_pcs_ibm_invalid_code                                        => "dis_ibm_invalid_code",
			hssi_8g_rx_pcs_invalid_code_flag_only                                  => "dis_invalid_code_only",
			hssi_8g_rx_pcs_pad_or_edb_error_replace                                => "replace_edb",
			hssi_8g_rx_pcs_pcs_bypass                                              => "dis_pcs_bypass",
			hssi_8g_rx_pcs_phase_comp_rdptr                                        => "enable_rdptr",
			hssi_8g_rx_pcs_phase_compensation_fifo                                 => "low_latency",
			hssi_8g_rx_pcs_pipe_if_enable                                          => "dis_pipe_rx",
			hssi_8g_rx_pcs_pma_dw                                                  => "twenty_bit",
			hssi_8g_rx_pcs_polinv_8b10b_dec                                        => "dis_polinv_8b10b_dec",
			hssi_8g_rx_pcs_prot_mode                                               => "basic_rm_disable",
			hssi_8g_rx_pcs_rate_match                                              => "dis_rm",
			hssi_8g_rx_pcs_rate_match_del_thres                                    => "dis_rm_del_thres",
			hssi_8g_rx_pcs_rate_match_empty_thres                                  => "dis_rm_empty_thres",
			hssi_8g_rx_pcs_rate_match_full_thres                                   => "dis_rm_full_thres",
			hssi_8g_rx_pcs_rate_match_ins_thres                                    => "dis_rm_ins_thres",
			hssi_8g_rx_pcs_rate_match_start_thres                                  => "dis_rm_start_thres",
			hssi_8g_rx_pcs_rx_clk_free_running                                     => "en_rx_clk_free_run",
			hssi_8g_rx_pcs_rx_clk2                                                 => "rcvd_clk_clk2",
			hssi_8g_rx_pcs_rx_pcs_urst                                             => "en_rx_pcs_urst",
			hssi_8g_rx_pcs_rx_rcvd_clk                                             => "rcvd_clk_rcvd_clk",
			hssi_8g_rx_pcs_rx_rd_clk                                               => "pld_rx_clk",
			hssi_8g_rx_pcs_rx_refclk                                               => "dis_refclk_sel",
			hssi_8g_rx_pcs_rx_wr_clk                                               => "rx_clk2_div_1_2_4",
			hssi_8g_rx_pcs_sup_mode                                                => "user_mode",
			hssi_8g_rx_pcs_symbol_swap                                             => "dis_symbol_swap",
			hssi_8g_rx_pcs_sync_sm_idle_eios                                       => "dis_syncsm_idle",
			hssi_8g_rx_pcs_test_bus_sel                                            => "tx_testbus",
			hssi_8g_rx_pcs_tx_rx_parallel_loopback                                 => "dis_plpbk",
			hssi_8g_rx_pcs_wa_boundary_lock_ctrl                                   => "bit_slip",
			hssi_8g_rx_pcs_wa_clk_slip_spacing                                     => 16,
			hssi_8g_rx_pcs_wa_det_latency_sync_status_beh                          => "dont_care_assert_sync",
			hssi_8g_rx_pcs_wa_disp_err_flag                                        => "dis_disp_err_flag",
			hssi_8g_rx_pcs_wa_kchar                                                => "dis_kchar",
			hssi_8g_rx_pcs_wa_pd                                                   => "wa_pd_7",
			hssi_8g_rx_pcs_wa_pd_data                                              => "0",
			hssi_8g_rx_pcs_wa_pd_polarity                                          => "en_pd_both_pol",
			hssi_8g_rx_pcs_wa_pld_controlled                                       => "rising_edge_sensitive_dw",
			hssi_8g_rx_pcs_wa_renumber_data                                        => 3,
			hssi_8g_rx_pcs_wa_rgnumber_data                                        => 3,
			hssi_8g_rx_pcs_wa_rknumber_data                                        => 3,
			hssi_8g_rx_pcs_wa_rosnumber_data                                       => 1,
			hssi_8g_rx_pcs_wa_rvnumber_data                                        => 0,
			hssi_8g_rx_pcs_wa_sync_sm_ctrl                                         => "gige_sync_sm",
			hssi_8g_rx_pcs_wait_cnt                                                => 0,
			hssi_8g_tx_pcs_bit_reversal                                            => "dis_bit_reversal",
			hssi_8g_tx_pcs_bonding_dft_en                                          => "dft_dis",
			hssi_8g_tx_pcs_bonding_dft_val                                         => "dft_0",
			hssi_8g_tx_pcs_bypass_pipeline_reg                                     => "dis_bypass_pipeline",
			hssi_8g_tx_pcs_byte_serializer                                         => "dis_bs",
			hssi_8g_tx_pcs_clock_gate_bs_enc                                       => "dis_bs_enc_clk_gating",
			hssi_8g_tx_pcs_clock_gate_dw_fifowr                                    => "dis_dw_fifowr_clk_gating",
			hssi_8g_tx_pcs_clock_gate_fiford                                       => "dis_fiford_clk_gating",
			hssi_8g_tx_pcs_clock_gate_sw_fifowr                                    => "dis_sw_fifowr_clk_gating",
			hssi_8g_tx_pcs_clock_observation_in_pld_core                           => "internal_refclk_b",
			hssi_8g_tx_pcs_data_selection_8b10b_encoder_input                      => "normal_data_path",
			hssi_8g_tx_pcs_dynamic_clk_switch                                      => "dis_dyn_clk_switch",
			hssi_8g_tx_pcs_eightb_tenb_disp_ctrl                                   => "dis_disp_ctrl",
			hssi_8g_tx_pcs_eightb_tenb_encoder                                     => "dis_8b10b",
			hssi_8g_tx_pcs_force_echar                                             => "dis_force_echar",
			hssi_8g_tx_pcs_force_kchar                                             => "dis_force_kchar",
			hssi_8g_tx_pcs_gen3_tx_clk_sel                                         => "dis_tx_clk",
			hssi_8g_tx_pcs_gen3_tx_pipe_clk_sel                                    => "dis_tx_pipe_clk",
			hssi_8g_tx_pcs_hip_mode                                                => "dis_hip",
			hssi_8g_tx_pcs_pcs_bypass                                              => "dis_pcs_bypass",
			hssi_8g_tx_pcs_phase_comp_rdptr                                        => "enable_rdptr",
			hssi_8g_tx_pcs_phase_compensation_fifo                                 => "low_latency",
			hssi_8g_tx_pcs_phfifo_write_clk_sel                                    => "pld_tx_clk",
			hssi_8g_tx_pcs_pma_dw                                                  => "twenty_bit",
			hssi_8g_tx_pcs_prot_mode                                               => "basic",
			hssi_8g_tx_pcs_refclk_b_clk_sel                                        => "tx_pma_clock",
			hssi_8g_tx_pcs_revloop_back_rm                                         => "dis_rev_loopback_rx_rm",
			hssi_8g_tx_pcs_sup_mode                                                => "user_mode",
			hssi_8g_tx_pcs_symbol_swap                                             => "dis_symbol_swap",
			hssi_8g_tx_pcs_tx_bitslip                                              => "dis_tx_bitslip",
			hssi_8g_tx_pcs_tx_compliance_controlled_disparity                      => "dis_txcompliance",
			hssi_8g_tx_pcs_tx_fast_pld_reg                                         => "dis_tx_fast_pld_reg",
			hssi_8g_tx_pcs_txclk_freerun                                           => "en_freerun_tx",
			hssi_8g_tx_pcs_txpcs_urst                                              => "en_txpcs_urst",
			hssi_tx_pld_pcs_interface_hd_chnl_hip_en                               => "disable",
			hssi_tx_pld_pcs_interface_hd_chnl_hrdrstctl_en                         => "disable",
			hssi_tx_pld_pcs_interface_hd_chnl_prot_mode_tx                         => "basic_8gpcs_tx",
			hssi_tx_pld_pcs_interface_hd_chnl_ctrl_plane_bonding_tx                => "ctrl_master_tx",
			hssi_tx_pld_pcs_interface_hd_chnl_pma_dw_tx                            => "pma_20b_tx",
			hssi_tx_pld_pcs_interface_hd_chnl_pld_fifo_mode_tx                     => "fifo_tx",
			hssi_tx_pld_pcs_interface_hd_chnl_shared_fifo_width_tx                 => "single_tx",
			hssi_tx_pld_pcs_interface_hd_chnl_low_latency_en_tx                    => "disable",
			hssi_tx_pld_pcs_interface_hd_chnl_func_mode                            => "enable",
			hssi_tx_pld_pcs_interface_hd_chnl_channel_operation_mode               => "tx_rx_pair_enabled",
			hssi_tx_pld_pcs_interface_hd_chnl_lpbk_en                              => "disable",
			hssi_tx_pld_pcs_interface_hd_chnl_frequency_rules_en                   => "enable",
			hssi_tx_pld_pcs_interface_hd_chnl_pma_tx_clk_hz                        => 240000000,
			hssi_tx_pld_pcs_interface_hd_chnl_pld_tx_clk_hz                        => 240000000,
			hssi_tx_pld_pcs_interface_hd_chnl_pld_uhsif_tx_clk_hz                  => 0,
			hssi_tx_pld_pcs_interface_hd_fifo_channel_operation_mode               => "tx_rx_pair_enabled",
			hssi_tx_pld_pcs_interface_hd_fifo_prot_mode_tx                         => "non_teng_mode_tx",
			hssi_tx_pld_pcs_interface_hd_fifo_shared_fifo_width_tx                 => "single_tx",
			hssi_tx_pld_pcs_interface_hd_10g_channel_operation_mode                => "tx_rx_pair_enabled",
			hssi_tx_pld_pcs_interface_hd_10g_lpbk_en                               => "disable",
			hssi_tx_pld_pcs_interface_hd_10g_advanced_user_mode_tx                 => "disable",
			hssi_tx_pld_pcs_interface_hd_10g_pma_dw_tx                             => "pma_64b_tx",
			hssi_tx_pld_pcs_interface_hd_10g_fifo_mode_tx                          => "fifo_tx",
			hssi_tx_pld_pcs_interface_hd_10g_prot_mode_tx                          => "disabled_prot_mode_tx",
			hssi_tx_pld_pcs_interface_hd_10g_low_latency_en_tx                     => "disable",
			hssi_tx_pld_pcs_interface_hd_10g_shared_fifo_width_tx                  => "single_tx",
			hssi_tx_pld_pcs_interface_hd_8g_channel_operation_mode                 => "tx_rx_pair_enabled",
			hssi_tx_pld_pcs_interface_hd_8g_lpbk_en                                => "disable",
			hssi_tx_pld_pcs_interface_hd_8g_prot_mode_tx                           => "basic_tx",
			hssi_tx_pld_pcs_interface_hd_8g_hip_mode                               => "disable",
			hssi_tx_pld_pcs_interface_hd_8g_pma_dw_tx                              => "pma_20b_tx",
			hssi_tx_pld_pcs_interface_hd_8g_fifo_mode_tx                           => "fifo_tx",
			hssi_tx_pld_pcs_interface_hd_g3_prot_mode                              => "disabled_prot_mode",
			hssi_tx_pld_pcs_interface_hd_krfec_channel_operation_mode              => "tx_rx_pair_enabled",
			hssi_tx_pld_pcs_interface_hd_krfec_lpbk_en                             => "disable",
			hssi_tx_pld_pcs_interface_hd_krfec_prot_mode_tx                        => "disabled_prot_mode_tx",
			hssi_tx_pld_pcs_interface_hd_krfec_low_latency_en_tx                   => "disable",
			hssi_tx_pld_pcs_interface_hd_pmaif_lpbk_en                             => "disable",
			hssi_tx_pld_pcs_interface_hd_pmaif_channel_operation_mode              => "tx_rx_pair_enabled",
			hssi_tx_pld_pcs_interface_hd_pmaif_sim_mode                            => "disable",
			hssi_tx_pld_pcs_interface_hd_pmaif_prot_mode_tx                        => "eightg_basic_mode_tx",
			hssi_tx_pld_pcs_interface_hd_pmaif_pma_dw_tx                           => "pma_20b_tx",
			hssi_tx_pld_pcs_interface_hd_pldif_prot_mode_tx                        => "eightg_and_g3_pld_fifo_mode_tx",
			hssi_tx_pld_pcs_interface_hd_pldif_hrdrstctl_en                        => "disable",
			hssi_tx_pld_pcs_interface_pcs_tx_clk_source                            => "eightg",
			hssi_tx_pld_pcs_interface_pcs_tx_data_source                           => "hip_disable",
			hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_en                         => "delay1_clk_disable",
			hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_sel                        => "pcs_tx_clk",
			hssi_tx_pld_pcs_interface_pcs_tx_delay1_ctrl                           => "delay1_path0",
			hssi_tx_pld_pcs_interface_pcs_tx_delay1_data_sel                       => "one_ff_delay",
			hssi_tx_pld_pcs_interface_pcs_tx_delay2_clk_en                         => "delay2_clk_disable",
			hssi_tx_pld_pcs_interface_pcs_tx_delay2_ctrl                           => "delay2_path0",
			hssi_tx_pld_pcs_interface_pcs_tx_output_sel                            => "teng_output",
			hssi_tx_pld_pcs_interface_pcs_tx_clk_out_sel                           => "eightg_clk_out",
			hssi_rx_pld_pcs_interface_hd_chnl_hip_en                               => "disable",
			hssi_rx_pld_pcs_interface_hd_chnl_transparent_pcs_rx                   => "disable",
			hssi_rx_pld_pcs_interface_hd_chnl_hrdrstctl_en                         => "disable",
			hssi_rx_pld_pcs_interface_hd_chnl_prot_mode_rx                         => "basic_8gpcs_rm_disable_rx",
			hssi_rx_pld_pcs_interface_hd_chnl_ctrl_plane_bonding_rx                => "individual_rx",
			hssi_rx_pld_pcs_interface_hd_chnl_pma_dw_rx                            => "pma_20b_rx",
			hssi_rx_pld_pcs_interface_hd_chnl_pld_fifo_mode_rx                     => "fifo_rx",
			hssi_rx_pld_pcs_interface_hd_chnl_shared_fifo_width_rx                 => "single_rx",
			hssi_rx_pld_pcs_interface_hd_chnl_low_latency_en_rx                    => "disable",
			hssi_rx_pld_pcs_interface_hd_chnl_func_mode                            => "enable",
			hssi_rx_pld_pcs_interface_hd_chnl_channel_operation_mode               => "tx_rx_pair_enabled",
			hssi_rx_pld_pcs_interface_hd_chnl_lpbk_en                              => "disable",
			hssi_rx_pld_pcs_interface_hd_10g_advanced_user_mode_rx                 => "disable",
			hssi_rx_pld_pcs_interface_hd_chnl_frequency_rules_en                   => "enable",
			hssi_rx_pld_pcs_interface_hd_chnl_pma_rx_clk_hz                        => 240000000,
			hssi_rx_pld_pcs_interface_hd_chnl_pld_rx_clk_hz                        => 240000000,
			hssi_rx_pld_pcs_interface_hd_chnl_fref_clk_hz                          => 240000000,
			hssi_rx_pld_pcs_interface_hd_chnl_clklow_clk_hz                        => 240000000,
			hssi_rx_pld_pcs_interface_hd_fifo_channel_operation_mode               => "tx_rx_pair_enabled",
			hssi_rx_pld_pcs_interface_hd_fifo_prot_mode_rx                         => "non_teng_mode_rx",
			hssi_rx_pld_pcs_interface_hd_fifo_shared_fifo_width_rx                 => "single_rx",
			hssi_rx_pld_pcs_interface_hd_10g_channel_operation_mode                => "tx_rx_pair_enabled",
			hssi_rx_pld_pcs_interface_hd_10g_lpbk_en                               => "disable",
			hssi_rx_pld_pcs_interface_hd_10g_pma_dw_rx                             => "pma_64b_rx",
			hssi_rx_pld_pcs_interface_hd_10g_fifo_mode_rx                          => "fifo_rx",
			hssi_rx_pld_pcs_interface_hd_10g_prot_mode_rx                          => "disabled_prot_mode_rx",
			hssi_rx_pld_pcs_interface_hd_10g_low_latency_en_rx                     => "disable",
			hssi_rx_pld_pcs_interface_hd_10g_shared_fifo_width_rx                  => "single_rx",
			hssi_rx_pld_pcs_interface_hd_10g_test_bus_mode                         => "rx",
			hssi_rx_pld_pcs_interface_hd_8g_channel_operation_mode                 => "tx_rx_pair_enabled",
			hssi_rx_pld_pcs_interface_hd_8g_lpbk_en                                => "disable",
			hssi_rx_pld_pcs_interface_hd_8g_prot_mode_rx                           => "basic_rm_disable_rx",
			hssi_rx_pld_pcs_interface_hd_8g_hip_mode                               => "disable",
			hssi_rx_pld_pcs_interface_hd_8g_pma_dw_rx                              => "pma_20b_rx",
			hssi_rx_pld_pcs_interface_hd_8g_fifo_mode_rx                           => "fifo_rx",
			hssi_rx_pld_pcs_interface_hd_g3_prot_mode                              => "disabled_prot_mode",
			hssi_rx_pld_pcs_interface_hd_krfec_channel_operation_mode              => "tx_rx_pair_enabled",
			hssi_rx_pld_pcs_interface_hd_krfec_lpbk_en                             => "disable",
			hssi_rx_pld_pcs_interface_hd_krfec_prot_mode_rx                        => "disabled_prot_mode_rx",
			hssi_rx_pld_pcs_interface_hd_krfec_low_latency_en_rx                   => "disable",
			hssi_rx_pld_pcs_interface_hd_krfec_test_bus_mode                       => "tx",
			hssi_rx_pld_pcs_interface_hd_pmaif_lpbk_en                             => "disable",
			hssi_rx_pld_pcs_interface_hd_pmaif_channel_operation_mode              => "tx_rx_pair_enabled",
			hssi_rx_pld_pcs_interface_hd_pmaif_sim_mode                            => "disable",
			hssi_rx_pld_pcs_interface_hd_pmaif_prot_mode_rx                        => "eightg_basic_mode_rx",
			hssi_rx_pld_pcs_interface_hd_pmaif_pma_dw_rx                           => "pma_20b_rx",
			hssi_rx_pld_pcs_interface_hd_pldif_prot_mode_rx                        => "eightg_and_g3_pld_fifo_mode_rx",
			hssi_rx_pld_pcs_interface_hd_pldif_hrdrstctl_en                        => "disable",
			hssi_rx_pld_pcs_interface_pcs_rx_block_sel                             => "eightg",
			hssi_rx_pld_pcs_interface_pcs_rx_clk_sel                               => "pld_rx_clk",
			hssi_rx_pld_pcs_interface_pcs_rx_hip_clk_en                            => "hip_rx_disable",
			hssi_rx_pld_pcs_interface_pcs_rx_output_sel                            => "teng_output",
			hssi_rx_pld_pcs_interface_pcs_rx_clk_out_sel                           => "eightg_clk_out",
			hssi_common_pld_pcs_interface_dft_clk_out_en                           => "dft_clk_out_disable",
			hssi_common_pld_pcs_interface_dft_clk_out_sel                          => "teng_rx_dft_clk",
			hssi_common_pld_pcs_interface_hrdrstctrl_en                            => "hrst_dis",
			hssi_common_pld_pcs_interface_pcs_testbus_block_sel                    => "pma_if",
			hssi_rx_pcs_pma_interface_block_sel                                    => "eight_g_pcs",
			hssi_rx_pcs_pma_interface_channel_operation_mode                       => "tx_rx_pair_enabled",
			hssi_rx_pcs_pma_interface_clkslip_sel                                  => "pld",
			hssi_rx_pcs_pma_interface_lpbk_en                                      => "disable",
			hssi_rx_pcs_pma_interface_master_clk_sel                               => "master_rx_pma_clk",
			hssi_rx_pcs_pma_interface_pldif_datawidth_mode                         => "pldif_data_10bit",
			hssi_rx_pcs_pma_interface_pma_dw_rx                                    => "pma_20b_rx",
			hssi_rx_pcs_pma_interface_pma_if_dft_en                                => "dft_dis",
			hssi_rx_pcs_pma_interface_pma_if_dft_val                               => "dft_0",
			hssi_rx_pcs_pma_interface_prbs_clken                                   => "prbs_clk_dis",
			hssi_rx_pcs_pma_interface_prbs_ver                                     => "prbs_off",
			hssi_rx_pcs_pma_interface_prbs9_dwidth                                 => "prbs9_64b",
			hssi_rx_pcs_pma_interface_prot_mode_rx                                 => "eightg_basic_mode_rx",
			hssi_rx_pcs_pma_interface_rx_dyn_polarity_inversion                    => "rx_dyn_polinv_en",
			hssi_rx_pcs_pma_interface_rx_lpbk_en                                   => "lpbk_dis",
			hssi_rx_pcs_pma_interface_rx_prbs_force_signal_ok                      => "force_sig_ok",
			hssi_rx_pcs_pma_interface_rx_prbs_mask                                 => "prbsmask128",
			hssi_rx_pcs_pma_interface_rx_prbs_mode                                 => "teng_mode",
			hssi_rx_pcs_pma_interface_rx_signalok_signaldet_sel                    => "sel_sig_det",
			hssi_rx_pcs_pma_interface_rx_static_polarity_inversion                 => "rx_stat_polinv_dis",
			hssi_rx_pcs_pma_interface_rx_uhsif_lpbk_en                             => "uhsif_lpbk_dis",
			hssi_rx_pcs_pma_interface_sup_mode                                     => "user_mode",
			hssi_tx_pcs_pma_interface_bypass_pma_txelecidle                        => "true",
			hssi_tx_pcs_pma_interface_channel_operation_mode                       => "tx_rx_pair_enabled",
			hssi_tx_pcs_pma_interface_lpbk_en                                      => "disable",
			hssi_tx_pcs_pma_interface_master_clk_sel                               => "master_tx_pma_clk",
			hssi_tx_pcs_pma_interface_pcie_sub_prot_mode_tx                        => "other_prot_mode",
			hssi_tx_pcs_pma_interface_pldif_datawidth_mode                         => "pldif_data_10bit",
			hssi_tx_pcs_pma_interface_pma_dw_tx                                    => "pma_20b_tx",
			hssi_tx_pcs_pma_interface_pma_if_dft_en                                => "dft_dis",
			hssi_tx_pcs_pma_interface_pmagate_en                                   => "pmagate_dis",
			hssi_tx_pcs_pma_interface_prbs_clken                                   => "prbs_clk_dis",
			hssi_tx_pcs_pma_interface_prbs_gen_pat                                 => "prbs_gen_dis",
			hssi_tx_pcs_pma_interface_prbs9_dwidth                                 => "prbs9_64b",
			hssi_tx_pcs_pma_interface_prot_mode_tx                                 => "eightg_basic_mode_tx",
			hssi_tx_pcs_pma_interface_sq_wave_num                                  => "sq_wave_default",
			hssi_tx_pcs_pma_interface_sqwgen_clken                                 => "sqwgen_clk_dis",
			hssi_tx_pcs_pma_interface_sup_mode                                     => "user_mode",
			hssi_tx_pcs_pma_interface_tx_dyn_polarity_inversion                    => "tx_dyn_polinv_en",
			hssi_tx_pcs_pma_interface_tx_pma_data_sel                              => "eight_g_pcs",
			hssi_tx_pcs_pma_interface_tx_static_polarity_inversion                 => "tx_stat_polinv_dis",
			hssi_tx_pcs_pma_interface_uhsif_cnt_step_filt_before_lock              => "uhsif_filt_stepsz_b4lock_2",
			hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_after_lock_value       => 0,
			hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_before_lock            => "uhsif_filt_cntthr_b4lock_8",
			hssi_tx_pcs_pma_interface_uhsif_dcn_test_update_period                 => "uhsif_dcn_test_period_4",
			hssi_tx_pcs_pma_interface_uhsif_dcn_testmode_enable                    => "uhsif_dcn_test_mode_disable",
			hssi_tx_pcs_pma_interface_uhsif_dead_zone_count_thresh                 => "uhsif_dzt_cnt_thr_2",
			hssi_tx_pcs_pma_interface_uhsif_dead_zone_detection_enable             => "uhsif_dzt_disable",
			hssi_tx_pcs_pma_interface_uhsif_dead_zone_obser_window                 => "uhsif_dzt_obr_win_16",
			hssi_tx_pcs_pma_interface_uhsif_dead_zone_skip_size                    => "uhsif_dzt_skipsz_4",
			hssi_tx_pcs_pma_interface_uhsif_delay_cell_index_sel                   => "uhsif_index_cram",
			hssi_tx_pcs_pma_interface_uhsif_delay_cell_margin                      => "uhsif_dcn_margin_2",
			hssi_tx_pcs_pma_interface_uhsif_delay_cell_static_index_value          => 0,
			hssi_tx_pcs_pma_interface_uhsif_dft_dead_zone_control                  => "uhsif_dft_dz_det_val_0",
			hssi_tx_pcs_pma_interface_uhsif_dft_up_filt_control                    => "uhsif_dft_up_val_0",
			hssi_tx_pcs_pma_interface_uhsif_enable                                 => "uhsif_disable",
			hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_after_lock              => "uhsif_lkd_segsz_aflock_512",
			hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_before_lock             => "uhsif_lkd_segsz_b4lock_16",
			hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_after_lock_value   => 0,
			hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_before_lock_value  => 0,
			hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_after_lock_value  => 0,
			hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_before_lock_value => 0,
			hssi_common_pcs_pma_interface_asn_clk_enable                           => "false",
			hssi_common_pcs_pma_interface_asn_enable                               => "dis_asn",
			hssi_common_pcs_pma_interface_block_sel                                => "eight_g_pcs",
			hssi_common_pcs_pma_interface_bypass_early_eios                        => "true",
			hssi_common_pcs_pma_interface_bypass_pcie_switch                       => "true",
			hssi_common_pcs_pma_interface_bypass_pma_ltr                           => "true",
			hssi_common_pcs_pma_interface_bypass_pma_sw_done                       => "false",
			hssi_common_pcs_pma_interface_bypass_ppm_lock                          => "false",
			hssi_common_pcs_pma_interface_bypass_send_syncp_fbkp                   => "true",
			hssi_common_pcs_pma_interface_bypass_txdetectrx                        => "true",
			hssi_common_pcs_pma_interface_cdr_control                              => "dis_cdr_ctrl",
			hssi_common_pcs_pma_interface_cid_enable                               => "dis_cid_mode",
			hssi_common_pcs_pma_interface_data_mask_count                          => 0,
			hssi_common_pcs_pma_interface_data_mask_count_multi                    => 0,
			hssi_common_pcs_pma_interface_dft_observation_clock_selection          => "dft_clk_obsrv_tx0",
			hssi_common_pcs_pma_interface_early_eios_counter                       => 0,
			hssi_common_pcs_pma_interface_force_freqdet                            => "force_freqdet_dis",
			hssi_common_pcs_pma_interface_free_run_clk_enable                      => "false",
			hssi_common_pcs_pma_interface_ignore_sigdet_g23                        => "false",
			hssi_common_pcs_pma_interface_pc_en_counter                            => 0,
			hssi_common_pcs_pma_interface_pc_rst_counter                           => 0,
			hssi_common_pcs_pma_interface_pcie_hip_mode                            => "hip_disable",
			hssi_common_pcs_pma_interface_ph_fifo_reg_mode                         => "phfifo_reg_mode_dis",
			hssi_common_pcs_pma_interface_phfifo_flush_wait                        => 0,
			hssi_common_pcs_pma_interface_pipe_if_g3pcs                            => "pipe_if_8gpcs",
			hssi_common_pcs_pma_interface_pma_done_counter                         => 0,
			hssi_common_pcs_pma_interface_pma_if_dft_en                            => "dft_dis",
			hssi_common_pcs_pma_interface_pma_if_dft_val                           => "dft_0",
			hssi_common_pcs_pma_interface_ppm_cnt_rst                              => "ppm_cnt_rst_dis",
			hssi_common_pcs_pma_interface_ppm_deassert_early                       => "deassert_early_dis",
			hssi_common_pcs_pma_interface_ppm_gen1_2_cnt                           => "cnt_32k",
			hssi_common_pcs_pma_interface_ppm_post_eidle_delay                     => "cnt_200_cycles",
			hssi_common_pcs_pma_interface_ppmsel                                   => "ppmsel_1000",
			hssi_common_pcs_pma_interface_prot_mode                                => "other_protocols",
			hssi_common_pcs_pma_interface_rxvalid_mask                             => "rxvalid_mask_dis",
			hssi_common_pcs_pma_interface_sigdet_wait_counter                      => 0,
			hssi_common_pcs_pma_interface_sigdet_wait_counter_multi                => 0,
			hssi_common_pcs_pma_interface_sim_mode                                 => "disable",
			hssi_common_pcs_pma_interface_spd_chg_rst_wait_cnt_en                  => "false",
			hssi_common_pcs_pma_interface_sup_mode                                 => "user_mode",
			hssi_common_pcs_pma_interface_testout_sel                              => "ppm_det_test",
			hssi_common_pcs_pma_interface_wait_clk_on_off_timer                    => 0,
			hssi_common_pcs_pma_interface_wait_pipe_synchronizing                  => 0,
			hssi_common_pcs_pma_interface_wait_send_syncp_fbkp                     => 0,
			hssi_common_pcs_pma_interface_ppm_det_buckets                          => "ppm_300_100_bucket",
			hssi_fifo_rx_pcs_double_read_mode                                      => "double_read_dis",
			hssi_fifo_rx_pcs_prot_mode                                             => "non_teng_mode",
			hssi_fifo_tx_pcs_double_write_mode                                     => "double_write_dis",
			hssi_fifo_tx_pcs_prot_mode                                             => "non_teng_mode",
			hssi_pipe_gen3_bypass_rx_detection_enable                              => "false",
			hssi_pipe_gen3_bypass_rx_preset                                        => 0,
			hssi_pipe_gen3_bypass_rx_preset_enable                                 => "false",
			hssi_pipe_gen3_bypass_tx_coefficent                                    => 0,
			hssi_pipe_gen3_bypass_tx_coefficent_enable                             => "false",
			hssi_pipe_gen3_elecidle_delay_g3                                       => 0,
			hssi_pipe_gen3_ind_error_reporting                                     => "dis_ind_error_reporting",
			hssi_pipe_gen3_mode                                                    => "disable_pcs",
			hssi_pipe_gen3_phy_status_delay_g12                                    => 0,
			hssi_pipe_gen3_phy_status_delay_g3                                     => 0,
			hssi_pipe_gen3_phystatus_rst_toggle_g12                                => "dis_phystatus_rst_toggle",
			hssi_pipe_gen3_phystatus_rst_toggle_g3                                 => "dis_phystatus_rst_toggle_g3",
			hssi_pipe_gen3_rate_match_pad_insertion                                => "dis_rm_fifo_pad_ins",
			hssi_pipe_gen3_sup_mode                                                => "user_mode",
			hssi_pipe_gen3_test_out_sel                                            => "disable_test_out",
			hssi_pipe_gen1_2_elec_idle_delay_val                                   => 0,
			hssi_pipe_gen1_2_error_replace_pad                                     => "replace_edb",
			hssi_pipe_gen1_2_hip_mode                                              => "dis_hip",
			hssi_pipe_gen1_2_ind_error_reporting                                   => "dis_ind_error_reporting",
			hssi_pipe_gen1_2_phystatus_delay_val                                   => 0,
			hssi_pipe_gen1_2_phystatus_rst_toggle                                  => "dis_phystatus_rst_toggle",
			hssi_pipe_gen1_2_pipe_byte_de_serializer_en                            => "dont_care_bds",
			hssi_pipe_gen1_2_prot_mode                                             => "basic",
			hssi_pipe_gen1_2_rx_pipe_enable                                        => "dis_pipe_rx",
			hssi_pipe_gen1_2_rxdetect_bypass                                       => "dis_rxdetect_bypass",
			hssi_pipe_gen1_2_sup_mode                                              => "user_mode",
			hssi_pipe_gen1_2_tx_pipe_enable                                        => "dis_pipe_tx",
			hssi_pipe_gen1_2_txswing                                               => "dis_txswing",
			pma_adapt_adp_1s_ctle_bypass                                           => "radp_1s_ctle_bypass_1",
			pma_adapt_adp_4s_ctle_bypass                                           => "radp_4s_ctle_bypass_1",
			pma_adapt_adp_ctle_en                                                  => "radp_ctle_disable",
			pma_adapt_adp_dfe_fltap_bypass                                         => "radp_dfe_fltap_bypass_1",
			pma_adapt_adp_dfe_fltap_en                                             => "radp_dfe_fltap_disable",
			pma_adapt_adp_dfe_fxtap_bypass                                         => "radp_dfe_fxtap_bypass_1",
			pma_adapt_adp_dfe_fxtap_en                                             => "radp_dfe_fxtap_disable",
			pma_adapt_adp_dfe_fxtap_hold_en                                        => "radp_dfe_fxtap_not_held",
			pma_adapt_adp_dfe_mode                                                 => "radp_dfe_mode_4",
			pma_adapt_adp_vga_bypass                                               => "radp_vga_bypass_1",
			pma_adapt_adp_vga_en                                                   => "radp_vga_disable",
			pma_adapt_adp_vref_bypass                                              => "radp_vref_bypass_1",
			pma_adapt_adp_vref_en                                                  => "radp_vref_disable",
			pma_adapt_datarate                                                     => "4800000000 bps",
			pma_adapt_prot_mode                                                    => "basic_rx",
			pma_adapt_sup_mode                                                     => "user_mode",
			pma_adapt_adp_ctle_adapt_cycle_window                                  => "radp_ctle_adapt_cycle_window_7",
			pma_adapt_odi_dfe_spec_en                                              => "rodi_dfe_spec_en_0",
			pma_adapt_adapt_mode                                                   => "manual",
			pma_adapt_adp_onetime_dfe                                              => "radp_onetime_dfe_0",
			pma_adapt_adp_mode                                                     => "radp_mode_8",
			pma_cdr_refclk_powerdown_mode                                          => "powerup",
			pma_cdr_refclk_refclk_select                                           => "ref_iqclk0",
			pma_cgb_bitslip_enable                                                 => "disable_bitslip",
			pma_cgb_bonding_reset_enable                                           => "disallow_bonding_reset",
			pma_cgb_datarate                                                       => "4800000000 bps",
			pma_cgb_pcie_gen3_bitwidth                                             => "pciegen3_wide",
			pma_cgb_prot_mode                                                      => "basic_tx",
			pma_cgb_ser_mode                                                       => "twenty_bit",
			pma_cgb_sup_mode                                                       => "user_mode",
			pma_cgb_x1_div_m_sel                                                   => "divbypass",
			pma_cgb_input_select_x1                                                => "unused",
			pma_cgb_input_select_gen3                                              => "unused",
			pma_cgb_input_select_xn                                                => "sel_x6_dn",
			pma_cgb_tx_ucontrol_en                                                 => "disable",
			pma_rx_dfe_datarate                                                    => "4800000000 bps",
			pma_rx_dfe_dft_en                                                      => "dft_disable",
			pma_rx_dfe_pdb                                                         => "dfe_enable",
			pma_rx_dfe_pdb_fixedtap                                                => "fixtap_dfe_powerdown",
			pma_rx_dfe_pdb_floattap                                                => "floattap_dfe_powerdown",
			pma_rx_dfe_pdb_fxtap4t7                                                => "fxtap4t7_powerdown",
			pma_rx_dfe_sup_mode                                                    => "user_mode",
			pma_rx_dfe_prot_mode                                                   => "basic_rx",
			pma_rx_odi_datarate                                                    => "4800000000 bps",
			pma_rx_odi_sup_mode                                                    => "user_mode",
			pma_rx_odi_step_ctrl_sel                                               => "dprio_mode",
			pma_rx_odi_prot_mode                                                   => "basic_rx",
			pma_rx_buf_bypass_eqz_stages_234                                       => "bypass_off",
			pma_rx_buf_datarate                                                    => "4800000000 bps",
			pma_rx_buf_diag_lp_en                                                  => "dlp_off",
			pma_rx_buf_prot_mode                                                   => "basic_rx",
			pma_rx_buf_qpi_enable                                                  => "non_qpi_mode",
			pma_rx_buf_rx_refclk_divider                                           => "bypass_divider",
			pma_rx_buf_sup_mode                                                    => "user_mode",
			pma_rx_buf_loopback_modes                                              => "lpbk_disable",
			pma_rx_buf_refclk_en                                                   => "disable",
			pma_rx_buf_pm_tx_rx_pcie_gen                                           => "non_pcie",
			pma_rx_buf_pm_tx_rx_pcie_gen_bitwidth                                  => "pcie_gen3_32b",
			pma_rx_buf_pm_tx_rx_cvp_mode                                           => "cvp_off",
			pma_rx_buf_xrx_path_uc_cal_enable                                      => "rx_cal_off",
			pma_rx_buf_xrx_path_sup_mode                                           => "user_mode",
			pma_rx_buf_xrx_path_prot_mode                                          => "basic_rx",
			pma_rx_buf_xrx_path_datarate                                           => "4800000000 bps",
			pma_rx_buf_xrx_path_datawidth                                          => 20,
			pma_rx_buf_xrx_path_pma_rx_divclk_hz                                   => "240000000",
			pma_rx_sd_prot_mode                                                    => "basic_rx",
			pma_rx_sd_sd_output_off                                                => 1,
			pma_rx_sd_sd_output_on                                                 => 15,
			pma_rx_sd_sd_pdb                                                       => "sd_off",
			pma_rx_sd_sd_threshold                                                 => 3,
			pma_rx_sd_sup_mode                                                     => "user_mode",
			pma_tx_ser_ser_clk_divtx_user_sel                                      => "divtx_user_off",
			pma_tx_ser_sup_mode                                                    => "user_mode",
			pma_tx_ser_prot_mode                                                   => "basic_tx",
			pma_tx_buf_datarate                                                    => "4800000000 bps",
			pma_tx_buf_prot_mode                                                   => "basic_tx",
			pma_tx_buf_rx_det                                                      => "mode_0",
			pma_tx_buf_rx_det_output_sel                                           => "rx_det_pcie_out",
			pma_tx_buf_rx_det_pdb                                                  => "rx_det_off",
			pma_tx_buf_sup_mode                                                    => "user_mode",
			pma_tx_buf_user_fir_coeff_ctrl_sel                                     => "ram_ctl",
			pma_tx_buf_xtx_path_prot_mode                                          => "basic_tx",
			pma_tx_buf_xtx_path_datarate                                           => "4800000000 bps",
			pma_tx_buf_xtx_path_datawidth                                          => 20,
			pma_tx_buf_xtx_path_clock_divider_ratio                                => 1,
			pma_tx_buf_xtx_path_pma_tx_divclk_hz                                   => "240000000",
			pma_tx_buf_xtx_path_tx_pll_clk_hz                                      => "2400000000",
			pma_tx_buf_xtx_path_sup_mode                                           => "user_mode",
			cdr_pll_pma_width                                                      => 20,
			cdr_pll_cgb_div                                                        => 1,
			cdr_pll_is_cascaded_pll                                                => "false",
			cdr_pll_datarate                                                       => "4800000000 bps",
			cdr_pll_lpd_counter                                                    => 4,
			cdr_pll_lpfd_counter                                                   => 2,
			cdr_pll_n_counter_scratch                                              => 1,
			cdr_pll_output_clock_frequency                                         => "2400000000 Hz",
			cdr_pll_reference_clock_frequency                                      => "240000000 hz",
			cdr_pll_set_cdr_vco_speed                                              => 2,
			cdr_pll_set_cdr_vco_speed_fix                                          => 117,
			cdr_pll_vco_freq                                                       => "9600000000 Hz",
			cdr_pll_atb_select_control                                             => "atb_off",
			cdr_pll_auto_reset_on                                                  => "auto_reset_off",
			cdr_pll_bbpd_data_pattern_filter_select                                => "bbpd_data_pat_off",
			cdr_pll_bw_sel                                                         => "medium",
			cdr_pll_cdr_odi_select                                                 => "sel_cdr",
			cdr_pll_cdr_phaselock_mode                                             => "no_ignore_lock",
			cdr_pll_cdr_powerdown_mode                                             => "power_up",
			cdr_pll_chgpmp_current_pd                                              => "cp_current_pd_setting0",
			cdr_pll_chgpmp_current_pfd                                             => "cp_current_pfd_setting2",
			cdr_pll_chgpmp_replicate                                               => "false",
			cdr_pll_chgpmp_testmode                                                => "cp_test_disable",
			cdr_pll_clklow_mux_select                                              => "clklow_mux_cdr_fbclk",
			cdr_pll_diag_loopback_enable                                           => "false",
			cdr_pll_disable_up_dn                                                  => "true",
			cdr_pll_fref_clklow_div                                                => 1,
			cdr_pll_fref_mux_select                                                => "fref_mux_cdr_refclk",
			cdr_pll_gpon_lck2ref_control                                           => "gpon_lck2ref_off",
			cdr_pll_initial_settings                                               => "true",
			cdr_pll_lck2ref_delay_control                                          => "lck2ref_delay_2",
			cdr_pll_lf_resistor_pd                                                 => "lf_pd_setting0",
			cdr_pll_lf_resistor_pfd                                                => "lf_pfd_setting2",
			cdr_pll_lf_ripple_cap                                                  => "lf_no_ripple",
			cdr_pll_loop_filter_bias_select                                        => "lpflt_bias_7",
			cdr_pll_loopback_mode                                                  => "loopback_disabled",
			cdr_pll_ltd_ltr_micro_controller_select                                => "ltd_ltr_pcs",
			cdr_pll_m_counter                                                      => 20,
			cdr_pll_n_counter                                                      => 1,
			cdr_pll_pd_fastlock_mode                                               => "false",
			cdr_pll_pd_l_counter                                                   => 4,
			cdr_pll_pfd_l_counter                                                  => 2,
			cdr_pll_primary_use                                                    => "cdr",
			cdr_pll_prot_mode                                                      => "basic_rx",
			cdr_pll_reverse_serial_loopback                                        => "no_loopback",
			cdr_pll_set_cdr_v2i_enable                                             => "true",
			cdr_pll_set_cdr_vco_reset                                              => "false",
			cdr_pll_set_cdr_vco_speed_pciegen3                                     => "cdr_vco_max_speedbin_pciegen3",
			cdr_pll_sup_mode                                                       => "user_mode",
			cdr_pll_tx_pll_prot_mode                                               => "txpll_unused",
			cdr_pll_txpll_hclk_driver_enable                                       => "false",
			cdr_pll_vco_overrange_voltage                                          => "vco_overrange_off",
			cdr_pll_vco_underrange_voltage                                         => "vco_underange_off",
			cdr_pll_fb_select                                                      => "direct_fb",
			cdr_pll_uc_ro_cal                                                      => "uc_ro_cal_on",
			cdr_pll_iqclk_mux_sel                                                  => "power_down",
			cdr_pll_pcie_gen                                                       => "non_pcie",
			cdr_pll_set_cdr_input_freq_range                                       => 0,
			cdr_pll_chgpmp_current_dn_trim                                         => "cp_current_trimming_dn_setting0",
			cdr_pll_chgpmp_up_pd_trim_double                                       => "normal_up_trim_current",
			cdr_pll_chgpmp_current_up_pd                                           => "cp_current_pd_up_setting4",
			cdr_pll_chgpmp_current_up_trim                                         => "cp_current_trimming_up_setting0",
			cdr_pll_chgpmp_dn_pd_trim_double                                       => "normal_dn_trim_current",
			cdr_pll_cal_vco_count_length                                           => "sel_8b_count",
			cdr_pll_chgpmp_current_dn_pd                                           => "cp_current_pd_dn_setting4",
			pma_rx_deser_clkdiv_source                                             => "vco_bypass_normal",
			pma_rx_deser_clkdivrx_user_mode                                        => "clkdivrx_user_disabled",
			pma_rx_deser_datarate                                                  => "4800000000 bps",
			pma_rx_deser_deser_factor                                              => 20,
			pma_rx_deser_force_clkdiv_for_testing                                  => "normal_clkdiv",
			pma_rx_deser_sdclk_enable                                              => "false",
			pma_rx_deser_sup_mode                                                  => "user_mode",
			pma_rx_deser_rst_n_adapt_odi                                           => "no_rst_adapt_odi",
			pma_rx_deser_bitslip_bypass                                            => "bs_bypass_yes",
			pma_rx_deser_prot_mode                                                 => "basic_rx",
			pma_rx_deser_pcie_gen                                                  => "non_pcie",
			pma_rx_deser_pcie_gen_bitwidth                                         => "pcie_gen3_32b"
		)
		port map (
			tx_analogreset                   => tx_analogreset,                                                                                                                                                                                                                                                                                                                                                                                     --     tx_analogreset.tx_analogreset
			tx_digitalreset                  => tx_digitalreset,                                                                                                                                                                                                                                                                                                                                                                                    --    tx_digitalreset.tx_digitalreset
			rx_analogreset                   => rx_analogreset,                                                                                                                                                                                                                                                                                                                                                                                     --     rx_analogreset.rx_analogreset
			rx_digitalreset                  => rx_digitalreset,                                                                                                                                                                                                                                                                                                                                                                                    --    rx_digitalreset.rx_digitalreset
			tx_cal_busy                      => tx_cal_busy,                                                                                                                                                                                                                                                                                                                                                                                        --        tx_cal_busy.tx_cal_busy
			rx_cal_busy                      => rx_cal_busy,                                                                                                                                                                                                                                                                                                                                                                                        --        rx_cal_busy.rx_cal_busy
			tx_bonding_clocks                => tx_bonding_clocks,                                                                                                                                                                                                                                                                                                                                                                                  --  tx_bonding_clocks.clk
			rx_cdr_refclk0                   => rx_cdr_refclk0,                                                                                                                                                                                                                                                                                                                                                                                     --     rx_cdr_refclk0.clk
			tx_serial_data                   => tx_serial_data,                                                                                                                                                                                                                                                                                                                                                                                     --     tx_serial_data.tx_serial_data
			rx_serial_data                   => rx_serial_data,                                                                                                                                                                                                                                                                                                                                                                                     --     rx_serial_data.rx_serial_data
			rx_seriallpbken                  => rx_seriallpbken,                                                                                                                                                                                                                                                                                                                                                                                    --    rx_seriallpbken.rx_seriallpbken
			rx_is_lockedtoref                => rx_is_lockedtoref,                                                                                                                                                                                                                                                                                                                                                                                  --  rx_is_lockedtoref.rx_is_lockedtoref
			rx_is_lockedtodata               => rx_is_lockedtodata,                                                                                                                                                                                                                                                                                                                                                                                 -- rx_is_lockedtodata.rx_is_lockedtodata
			tx_coreclkin                     => tx_coreclkin,                                                                                                                                                                                                                                                                                                                                                                                       --       tx_coreclkin.clk
			rx_coreclkin                     => rx_coreclkin,                                                                                                                                                                                                                                                                                                                                                                                       --       rx_coreclkin.clk
			tx_clkout                        => tx_clkout,                                                                                                                                                                                                                                                                                                                                                                                          --          tx_clkout.clk
			rx_clkout                        => rx_clkout,                                                                                                                                                                                                                                                                                                                                                                                          --          rx_clkout.clk
			tx_parallel_data(0 downto 0)     => tx_parallel_data(0 downto 0),                                                                                                                                                                                                                                                                                                                                                                       --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(1 downto 1)     => tx_parallel_data(1 downto 1),                                                                                                                                                                                                                                                                                                                                                                       --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(2 downto 2)     => tx_parallel_data(2 downto 2),                                                                                                                                                                                                                                                                                                                                                                       --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(3 downto 3)     => tx_parallel_data(3 downto 3),                                                                                                                                                                                                                                                                                                                                                                       --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(4 downto 4)     => tx_parallel_data(4 downto 4),                                                                                                                                                                                                                                                                                                                                                                       --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(5 downto 5)     => tx_parallel_data(5 downto 5),                                                                                                                                                                                                                                                                                                                                                                       --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(6 downto 6)     => tx_parallel_data(6 downto 6),                                                                                                                                                                                                                                                                                                                                                                       --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(7 downto 7)     => tx_parallel_data(7 downto 7),                                                                                                                                                                                                                                                                                                                                                                       --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(8 downto 8)     => tx_parallel_data(8 downto 8),                                                                                                                                                                                                                                                                                                                                                                       --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(9 downto 9)     => tx_parallel_data(9 downto 9),                                                                                                                                                                                                                                                                                                                                                                       --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(10 downto 10)   => unused_tx_parallel_data(0 downto 0),                                                                                                                                                                                                                                                                                                                                                                --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(11 downto 11)   => tx_parallel_data(10 downto 10),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(12 downto 12)   => tx_parallel_data(11 downto 11),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(13 downto 13)   => tx_parallel_data(12 downto 12),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(14 downto 14)   => tx_parallel_data(13 downto 13),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(15 downto 15)   => tx_parallel_data(14 downto 14),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(16 downto 16)   => tx_parallel_data(15 downto 15),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(17 downto 17)   => tx_parallel_data(16 downto 16),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(18 downto 18)   => tx_parallel_data(17 downto 17),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(19 downto 19)   => tx_parallel_data(18 downto 18),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(20 downto 20)   => tx_parallel_data(19 downto 19),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(21 downto 21)   => unused_tx_parallel_data(1 downto 1),                                                                                                                                                                                                                                                                                                                                                                --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(22 downto 22)   => unused_tx_parallel_data(2 downto 2),                                                                                                                                                                                                                                                                                                                                                                --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(23 downto 23)   => unused_tx_parallel_data(3 downto 3),                                                                                                                                                                                                                                                                                                                                                                --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(24 downto 24)   => unused_tx_parallel_data(4 downto 4),                                                                                                                                                                                                                                                                                                                                                                --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(25 downto 25)   => unused_tx_parallel_data(5 downto 5),                                                                                                                                                                                                                                                                                                                                                                --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(26 downto 26)   => unused_tx_parallel_data(6 downto 6),                                                                                                                                                                                                                                                                                                                                                                --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(27 downto 27)   => unused_tx_parallel_data(7 downto 7),                                                                                                                                                                                                                                                                                                                                                                --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(28 downto 28)   => unused_tx_parallel_data(8 downto 8),                                                                                                                                                                                                                                                                                                                                                                --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(29 downto 29)   => unused_tx_parallel_data(9 downto 9),                                                                                                                                                                                                                                                                                                                                                                --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(30 downto 30)   => unused_tx_parallel_data(10 downto 10),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(31 downto 31)   => unused_tx_parallel_data(11 downto 11),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(32 downto 32)   => unused_tx_parallel_data(12 downto 12),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(33 downto 33)   => unused_tx_parallel_data(13 downto 13),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(34 downto 34)   => unused_tx_parallel_data(14 downto 14),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(35 downto 35)   => unused_tx_parallel_data(15 downto 15),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(36 downto 36)   => unused_tx_parallel_data(16 downto 16),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(37 downto 37)   => unused_tx_parallel_data(17 downto 17),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(38 downto 38)   => unused_tx_parallel_data(18 downto 18),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(39 downto 39)   => unused_tx_parallel_data(19 downto 19),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(40 downto 40)   => unused_tx_parallel_data(20 downto 20),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(41 downto 41)   => unused_tx_parallel_data(21 downto 21),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(42 downto 42)   => unused_tx_parallel_data(22 downto 22),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(43 downto 43)   => unused_tx_parallel_data(23 downto 23),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(44 downto 44)   => unused_tx_parallel_data(24 downto 24),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(45 downto 45)   => unused_tx_parallel_data(25 downto 25),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(46 downto 46)   => unused_tx_parallel_data(26 downto 26),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(47 downto 47)   => unused_tx_parallel_data(27 downto 27),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(48 downto 48)   => unused_tx_parallel_data(28 downto 28),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(49 downto 49)   => unused_tx_parallel_data(29 downto 29),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(50 downto 50)   => unused_tx_parallel_data(30 downto 30),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(51 downto 51)   => unused_tx_parallel_data(31 downto 31),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(52 downto 52)   => unused_tx_parallel_data(32 downto 32),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(53 downto 53)   => unused_tx_parallel_data(33 downto 33),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(54 downto 54)   => unused_tx_parallel_data(34 downto 34),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(55 downto 55)   => unused_tx_parallel_data(35 downto 35),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(56 downto 56)   => unused_tx_parallel_data(36 downto 36),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(57 downto 57)   => unused_tx_parallel_data(37 downto 37),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(58 downto 58)   => unused_tx_parallel_data(38 downto 38),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(59 downto 59)   => unused_tx_parallel_data(39 downto 39),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(60 downto 60)   => unused_tx_parallel_data(40 downto 40),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(61 downto 61)   => unused_tx_parallel_data(41 downto 41),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(62 downto 62)   => unused_tx_parallel_data(42 downto 42),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(63 downto 63)   => unused_tx_parallel_data(43 downto 43),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(64 downto 64)   => unused_tx_parallel_data(44 downto 44),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(65 downto 65)   => unused_tx_parallel_data(45 downto 45),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(66 downto 66)   => unused_tx_parallel_data(46 downto 46),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(67 downto 67)   => unused_tx_parallel_data(47 downto 47),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(68 downto 68)   => unused_tx_parallel_data(48 downto 48),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(69 downto 69)   => unused_tx_parallel_data(49 downto 49),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(70 downto 70)   => unused_tx_parallel_data(50 downto 50),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(71 downto 71)   => unused_tx_parallel_data(51 downto 51),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(72 downto 72)   => unused_tx_parallel_data(52 downto 52),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(73 downto 73)   => unused_tx_parallel_data(53 downto 53),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(74 downto 74)   => unused_tx_parallel_data(54 downto 54),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(75 downto 75)   => unused_tx_parallel_data(55 downto 55),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(76 downto 76)   => unused_tx_parallel_data(56 downto 56),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(77 downto 77)   => unused_tx_parallel_data(57 downto 57),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(78 downto 78)   => unused_tx_parallel_data(58 downto 58),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(79 downto 79)   => unused_tx_parallel_data(59 downto 59),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(80 downto 80)   => unused_tx_parallel_data(60 downto 60),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(81 downto 81)   => unused_tx_parallel_data(61 downto 61),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(82 downto 82)   => unused_tx_parallel_data(62 downto 62),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(83 downto 83)   => unused_tx_parallel_data(63 downto 63),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(84 downto 84)   => unused_tx_parallel_data(64 downto 64),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(85 downto 85)   => unused_tx_parallel_data(65 downto 65),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(86 downto 86)   => unused_tx_parallel_data(66 downto 66),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(87 downto 87)   => unused_tx_parallel_data(67 downto 67),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(88 downto 88)   => unused_tx_parallel_data(68 downto 68),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(89 downto 89)   => unused_tx_parallel_data(69 downto 69),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(90 downto 90)   => unused_tx_parallel_data(70 downto 70),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(91 downto 91)   => unused_tx_parallel_data(71 downto 71),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(92 downto 92)   => unused_tx_parallel_data(72 downto 72),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(93 downto 93)   => unused_tx_parallel_data(73 downto 73),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(94 downto 94)   => unused_tx_parallel_data(74 downto 74),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(95 downto 95)   => unused_tx_parallel_data(75 downto 75),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(96 downto 96)   => unused_tx_parallel_data(76 downto 76),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(97 downto 97)   => unused_tx_parallel_data(77 downto 77),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(98 downto 98)   => unused_tx_parallel_data(78 downto 78),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(99 downto 99)   => unused_tx_parallel_data(79 downto 79),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(100 downto 100) => unused_tx_parallel_data(80 downto 80),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(101 downto 101) => unused_tx_parallel_data(81 downto 81),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(102 downto 102) => unused_tx_parallel_data(82 downto 82),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(103 downto 103) => unused_tx_parallel_data(83 downto 83),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(104 downto 104) => unused_tx_parallel_data(84 downto 84),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(105 downto 105) => unused_tx_parallel_data(85 downto 85),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(106 downto 106) => unused_tx_parallel_data(86 downto 86),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(107 downto 107) => unused_tx_parallel_data(87 downto 87),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(108 downto 108) => unused_tx_parallel_data(88 downto 88),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(109 downto 109) => unused_tx_parallel_data(89 downto 89),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(110 downto 110) => unused_tx_parallel_data(90 downto 90),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(111 downto 111) => unused_tx_parallel_data(91 downto 91),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(112 downto 112) => unused_tx_parallel_data(92 downto 92),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(113 downto 113) => unused_tx_parallel_data(93 downto 93),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(114 downto 114) => unused_tx_parallel_data(94 downto 94),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(115 downto 115) => unused_tx_parallel_data(95 downto 95),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(116 downto 116) => unused_tx_parallel_data(96 downto 96),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(117 downto 117) => unused_tx_parallel_data(97 downto 97),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(118 downto 118) => unused_tx_parallel_data(98 downto 98),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(119 downto 119) => unused_tx_parallel_data(99 downto 99),                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(120 downto 120) => unused_tx_parallel_data(100 downto 100),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(121 downto 121) => unused_tx_parallel_data(101 downto 101),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(122 downto 122) => unused_tx_parallel_data(102 downto 102),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(123 downto 123) => unused_tx_parallel_data(103 downto 103),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(124 downto 124) => unused_tx_parallel_data(104 downto 104),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(125 downto 125) => unused_tx_parallel_data(105 downto 105),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(126 downto 126) => unused_tx_parallel_data(106 downto 106),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(127 downto 127) => unused_tx_parallel_data(107 downto 107),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(128 downto 128) => tx_parallel_data(20 downto 20),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(129 downto 129) => tx_parallel_data(21 downto 21),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(130 downto 130) => tx_parallel_data(22 downto 22),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(131 downto 131) => tx_parallel_data(23 downto 23),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(132 downto 132) => tx_parallel_data(24 downto 24),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(133 downto 133) => tx_parallel_data(25 downto 25),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(134 downto 134) => tx_parallel_data(26 downto 26),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(135 downto 135) => tx_parallel_data(27 downto 27),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(136 downto 136) => tx_parallel_data(28 downto 28),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(137 downto 137) => tx_parallel_data(29 downto 29),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(138 downto 138) => unused_tx_parallel_data(108 downto 108),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(139 downto 139) => tx_parallel_data(30 downto 30),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(140 downto 140) => tx_parallel_data(31 downto 31),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(141 downto 141) => tx_parallel_data(32 downto 32),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(142 downto 142) => tx_parallel_data(33 downto 33),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(143 downto 143) => tx_parallel_data(34 downto 34),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(144 downto 144) => tx_parallel_data(35 downto 35),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(145 downto 145) => tx_parallel_data(36 downto 36),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(146 downto 146) => tx_parallel_data(37 downto 37),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(147 downto 147) => tx_parallel_data(38 downto 38),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(148 downto 148) => tx_parallel_data(39 downto 39),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(149 downto 149) => unused_tx_parallel_data(109 downto 109),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(150 downto 150) => unused_tx_parallel_data(110 downto 110),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(151 downto 151) => unused_tx_parallel_data(111 downto 111),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(152 downto 152) => unused_tx_parallel_data(112 downto 112),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(153 downto 153) => unused_tx_parallel_data(113 downto 113),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(154 downto 154) => unused_tx_parallel_data(114 downto 114),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(155 downto 155) => unused_tx_parallel_data(115 downto 115),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(156 downto 156) => unused_tx_parallel_data(116 downto 116),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(157 downto 157) => unused_tx_parallel_data(117 downto 117),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(158 downto 158) => unused_tx_parallel_data(118 downto 118),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(159 downto 159) => unused_tx_parallel_data(119 downto 119),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(160 downto 160) => unused_tx_parallel_data(120 downto 120),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(161 downto 161) => unused_tx_parallel_data(121 downto 121),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(162 downto 162) => unused_tx_parallel_data(122 downto 122),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(163 downto 163) => unused_tx_parallel_data(123 downto 123),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(164 downto 164) => unused_tx_parallel_data(124 downto 124),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(165 downto 165) => unused_tx_parallel_data(125 downto 125),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(166 downto 166) => unused_tx_parallel_data(126 downto 126),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(167 downto 167) => unused_tx_parallel_data(127 downto 127),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(168 downto 168) => unused_tx_parallel_data(128 downto 128),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(169 downto 169) => unused_tx_parallel_data(129 downto 129),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(170 downto 170) => unused_tx_parallel_data(130 downto 130),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(171 downto 171) => unused_tx_parallel_data(131 downto 131),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(172 downto 172) => unused_tx_parallel_data(132 downto 132),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(173 downto 173) => unused_tx_parallel_data(133 downto 133),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(174 downto 174) => unused_tx_parallel_data(134 downto 134),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(175 downto 175) => unused_tx_parallel_data(135 downto 135),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(176 downto 176) => unused_tx_parallel_data(136 downto 136),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(177 downto 177) => unused_tx_parallel_data(137 downto 137),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(178 downto 178) => unused_tx_parallel_data(138 downto 138),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(179 downto 179) => unused_tx_parallel_data(139 downto 139),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(180 downto 180) => unused_tx_parallel_data(140 downto 140),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(181 downto 181) => unused_tx_parallel_data(141 downto 141),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(182 downto 182) => unused_tx_parallel_data(142 downto 142),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(183 downto 183) => unused_tx_parallel_data(143 downto 143),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(184 downto 184) => unused_tx_parallel_data(144 downto 144),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(185 downto 185) => unused_tx_parallel_data(145 downto 145),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(186 downto 186) => unused_tx_parallel_data(146 downto 146),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(187 downto 187) => unused_tx_parallel_data(147 downto 147),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(188 downto 188) => unused_tx_parallel_data(148 downto 148),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(189 downto 189) => unused_tx_parallel_data(149 downto 149),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(190 downto 190) => unused_tx_parallel_data(150 downto 150),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(191 downto 191) => unused_tx_parallel_data(151 downto 151),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(192 downto 192) => unused_tx_parallel_data(152 downto 152),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(193 downto 193) => unused_tx_parallel_data(153 downto 153),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(194 downto 194) => unused_tx_parallel_data(154 downto 154),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(195 downto 195) => unused_tx_parallel_data(155 downto 155),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(196 downto 196) => unused_tx_parallel_data(156 downto 156),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(197 downto 197) => unused_tx_parallel_data(157 downto 157),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(198 downto 198) => unused_tx_parallel_data(158 downto 158),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(199 downto 199) => unused_tx_parallel_data(159 downto 159),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(200 downto 200) => unused_tx_parallel_data(160 downto 160),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(201 downto 201) => unused_tx_parallel_data(161 downto 161),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(202 downto 202) => unused_tx_parallel_data(162 downto 162),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(203 downto 203) => unused_tx_parallel_data(163 downto 163),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(204 downto 204) => unused_tx_parallel_data(164 downto 164),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(205 downto 205) => unused_tx_parallel_data(165 downto 165),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(206 downto 206) => unused_tx_parallel_data(166 downto 166),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(207 downto 207) => unused_tx_parallel_data(167 downto 167),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(208 downto 208) => unused_tx_parallel_data(168 downto 168),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(209 downto 209) => unused_tx_parallel_data(169 downto 169),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(210 downto 210) => unused_tx_parallel_data(170 downto 170),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(211 downto 211) => unused_tx_parallel_data(171 downto 171),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(212 downto 212) => unused_tx_parallel_data(172 downto 172),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(213 downto 213) => unused_tx_parallel_data(173 downto 173),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(214 downto 214) => unused_tx_parallel_data(174 downto 174),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(215 downto 215) => unused_tx_parallel_data(175 downto 175),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(216 downto 216) => unused_tx_parallel_data(176 downto 176),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(217 downto 217) => unused_tx_parallel_data(177 downto 177),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(218 downto 218) => unused_tx_parallel_data(178 downto 178),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(219 downto 219) => unused_tx_parallel_data(179 downto 179),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(220 downto 220) => unused_tx_parallel_data(180 downto 180),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(221 downto 221) => unused_tx_parallel_data(181 downto 181),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(222 downto 222) => unused_tx_parallel_data(182 downto 182),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(223 downto 223) => unused_tx_parallel_data(183 downto 183),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(224 downto 224) => unused_tx_parallel_data(184 downto 184),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(225 downto 225) => unused_tx_parallel_data(185 downto 185),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(226 downto 226) => unused_tx_parallel_data(186 downto 186),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(227 downto 227) => unused_tx_parallel_data(187 downto 187),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(228 downto 228) => unused_tx_parallel_data(188 downto 188),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(229 downto 229) => unused_tx_parallel_data(189 downto 189),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(230 downto 230) => unused_tx_parallel_data(190 downto 190),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(231 downto 231) => unused_tx_parallel_data(191 downto 191),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(232 downto 232) => unused_tx_parallel_data(192 downto 192),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(233 downto 233) => unused_tx_parallel_data(193 downto 193),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(234 downto 234) => unused_tx_parallel_data(194 downto 194),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(235 downto 235) => unused_tx_parallel_data(195 downto 195),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(236 downto 236) => unused_tx_parallel_data(196 downto 196),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(237 downto 237) => unused_tx_parallel_data(197 downto 197),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(238 downto 238) => unused_tx_parallel_data(198 downto 198),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(239 downto 239) => unused_tx_parallel_data(199 downto 199),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(240 downto 240) => unused_tx_parallel_data(200 downto 200),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(241 downto 241) => unused_tx_parallel_data(201 downto 201),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(242 downto 242) => unused_tx_parallel_data(202 downto 202),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(243 downto 243) => unused_tx_parallel_data(203 downto 203),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(244 downto 244) => unused_tx_parallel_data(204 downto 204),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(245 downto 245) => unused_tx_parallel_data(205 downto 205),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(246 downto 246) => unused_tx_parallel_data(206 downto 206),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(247 downto 247) => unused_tx_parallel_data(207 downto 207),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(248 downto 248) => unused_tx_parallel_data(208 downto 208),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(249 downto 249) => unused_tx_parallel_data(209 downto 209),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(250 downto 250) => unused_tx_parallel_data(210 downto 210),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(251 downto 251) => unused_tx_parallel_data(211 downto 211),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(252 downto 252) => unused_tx_parallel_data(212 downto 212),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(253 downto 253) => unused_tx_parallel_data(213 downto 213),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(254 downto 254) => unused_tx_parallel_data(214 downto 214),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(255 downto 255) => unused_tx_parallel_data(215 downto 215),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(256 downto 256) => tx_parallel_data(40 downto 40),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(257 downto 257) => tx_parallel_data(41 downto 41),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(258 downto 258) => tx_parallel_data(42 downto 42),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(259 downto 259) => tx_parallel_data(43 downto 43),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(260 downto 260) => tx_parallel_data(44 downto 44),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(261 downto 261) => tx_parallel_data(45 downto 45),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(262 downto 262) => tx_parallel_data(46 downto 46),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(263 downto 263) => tx_parallel_data(47 downto 47),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(264 downto 264) => tx_parallel_data(48 downto 48),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(265 downto 265) => tx_parallel_data(49 downto 49),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(266 downto 266) => unused_tx_parallel_data(216 downto 216),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(267 downto 267) => tx_parallel_data(50 downto 50),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(268 downto 268) => tx_parallel_data(51 downto 51),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(269 downto 269) => tx_parallel_data(52 downto 52),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(270 downto 270) => tx_parallel_data(53 downto 53),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(271 downto 271) => tx_parallel_data(54 downto 54),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(272 downto 272) => tx_parallel_data(55 downto 55),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(273 downto 273) => tx_parallel_data(56 downto 56),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(274 downto 274) => tx_parallel_data(57 downto 57),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(275 downto 275) => tx_parallel_data(58 downto 58),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(276 downto 276) => tx_parallel_data(59 downto 59),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(277 downto 277) => unused_tx_parallel_data(217 downto 217),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(278 downto 278) => unused_tx_parallel_data(218 downto 218),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(279 downto 279) => unused_tx_parallel_data(219 downto 219),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(280 downto 280) => unused_tx_parallel_data(220 downto 220),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(281 downto 281) => unused_tx_parallel_data(221 downto 221),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(282 downto 282) => unused_tx_parallel_data(222 downto 222),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(283 downto 283) => unused_tx_parallel_data(223 downto 223),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(284 downto 284) => unused_tx_parallel_data(224 downto 224),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(285 downto 285) => unused_tx_parallel_data(225 downto 225),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(286 downto 286) => unused_tx_parallel_data(226 downto 226),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(287 downto 287) => unused_tx_parallel_data(227 downto 227),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(288 downto 288) => unused_tx_parallel_data(228 downto 228),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(289 downto 289) => unused_tx_parallel_data(229 downto 229),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(290 downto 290) => unused_tx_parallel_data(230 downto 230),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(291 downto 291) => unused_tx_parallel_data(231 downto 231),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(292 downto 292) => unused_tx_parallel_data(232 downto 232),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(293 downto 293) => unused_tx_parallel_data(233 downto 233),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(294 downto 294) => unused_tx_parallel_data(234 downto 234),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(295 downto 295) => unused_tx_parallel_data(235 downto 235),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(296 downto 296) => unused_tx_parallel_data(236 downto 236),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(297 downto 297) => unused_tx_parallel_data(237 downto 237),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(298 downto 298) => unused_tx_parallel_data(238 downto 238),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(299 downto 299) => unused_tx_parallel_data(239 downto 239),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(300 downto 300) => unused_tx_parallel_data(240 downto 240),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(301 downto 301) => unused_tx_parallel_data(241 downto 241),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(302 downto 302) => unused_tx_parallel_data(242 downto 242),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(303 downto 303) => unused_tx_parallel_data(243 downto 243),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(304 downto 304) => unused_tx_parallel_data(244 downto 244),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(305 downto 305) => unused_tx_parallel_data(245 downto 245),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(306 downto 306) => unused_tx_parallel_data(246 downto 246),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(307 downto 307) => unused_tx_parallel_data(247 downto 247),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(308 downto 308) => unused_tx_parallel_data(248 downto 248),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(309 downto 309) => unused_tx_parallel_data(249 downto 249),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(310 downto 310) => unused_tx_parallel_data(250 downto 250),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(311 downto 311) => unused_tx_parallel_data(251 downto 251),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(312 downto 312) => unused_tx_parallel_data(252 downto 252),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(313 downto 313) => unused_tx_parallel_data(253 downto 253),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(314 downto 314) => unused_tx_parallel_data(254 downto 254),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(315 downto 315) => unused_tx_parallel_data(255 downto 255),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(316 downto 316) => unused_tx_parallel_data(256 downto 256),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(317 downto 317) => unused_tx_parallel_data(257 downto 257),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(318 downto 318) => unused_tx_parallel_data(258 downto 258),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(319 downto 319) => unused_tx_parallel_data(259 downto 259),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(320 downto 320) => unused_tx_parallel_data(260 downto 260),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(321 downto 321) => unused_tx_parallel_data(261 downto 261),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(322 downto 322) => unused_tx_parallel_data(262 downto 262),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(323 downto 323) => unused_tx_parallel_data(263 downto 263),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(324 downto 324) => unused_tx_parallel_data(264 downto 264),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(325 downto 325) => unused_tx_parallel_data(265 downto 265),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(326 downto 326) => unused_tx_parallel_data(266 downto 266),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(327 downto 327) => unused_tx_parallel_data(267 downto 267),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(328 downto 328) => unused_tx_parallel_data(268 downto 268),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(329 downto 329) => unused_tx_parallel_data(269 downto 269),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(330 downto 330) => unused_tx_parallel_data(270 downto 270),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(331 downto 331) => unused_tx_parallel_data(271 downto 271),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(332 downto 332) => unused_tx_parallel_data(272 downto 272),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(333 downto 333) => unused_tx_parallel_data(273 downto 273),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(334 downto 334) => unused_tx_parallel_data(274 downto 274),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(335 downto 335) => unused_tx_parallel_data(275 downto 275),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(336 downto 336) => unused_tx_parallel_data(276 downto 276),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(337 downto 337) => unused_tx_parallel_data(277 downto 277),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(338 downto 338) => unused_tx_parallel_data(278 downto 278),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(339 downto 339) => unused_tx_parallel_data(279 downto 279),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(340 downto 340) => unused_tx_parallel_data(280 downto 280),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(341 downto 341) => unused_tx_parallel_data(281 downto 281),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(342 downto 342) => unused_tx_parallel_data(282 downto 282),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(343 downto 343) => unused_tx_parallel_data(283 downto 283),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(344 downto 344) => unused_tx_parallel_data(284 downto 284),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(345 downto 345) => unused_tx_parallel_data(285 downto 285),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(346 downto 346) => unused_tx_parallel_data(286 downto 286),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(347 downto 347) => unused_tx_parallel_data(287 downto 287),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(348 downto 348) => unused_tx_parallel_data(288 downto 288),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(349 downto 349) => unused_tx_parallel_data(289 downto 289),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(350 downto 350) => unused_tx_parallel_data(290 downto 290),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(351 downto 351) => unused_tx_parallel_data(291 downto 291),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(352 downto 352) => unused_tx_parallel_data(292 downto 292),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(353 downto 353) => unused_tx_parallel_data(293 downto 293),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(354 downto 354) => unused_tx_parallel_data(294 downto 294),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(355 downto 355) => unused_tx_parallel_data(295 downto 295),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(356 downto 356) => unused_tx_parallel_data(296 downto 296),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(357 downto 357) => unused_tx_parallel_data(297 downto 297),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(358 downto 358) => unused_tx_parallel_data(298 downto 298),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(359 downto 359) => unused_tx_parallel_data(299 downto 299),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(360 downto 360) => unused_tx_parallel_data(300 downto 300),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(361 downto 361) => unused_tx_parallel_data(301 downto 301),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(362 downto 362) => unused_tx_parallel_data(302 downto 302),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(363 downto 363) => unused_tx_parallel_data(303 downto 303),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(364 downto 364) => unused_tx_parallel_data(304 downto 304),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(365 downto 365) => unused_tx_parallel_data(305 downto 305),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(366 downto 366) => unused_tx_parallel_data(306 downto 306),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(367 downto 367) => unused_tx_parallel_data(307 downto 307),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(368 downto 368) => unused_tx_parallel_data(308 downto 308),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(369 downto 369) => unused_tx_parallel_data(309 downto 309),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(370 downto 370) => unused_tx_parallel_data(310 downto 310),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(371 downto 371) => unused_tx_parallel_data(311 downto 311),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(372 downto 372) => unused_tx_parallel_data(312 downto 312),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(373 downto 373) => unused_tx_parallel_data(313 downto 313),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(374 downto 374) => unused_tx_parallel_data(314 downto 314),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(375 downto 375) => unused_tx_parallel_data(315 downto 315),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(376 downto 376) => unused_tx_parallel_data(316 downto 316),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(377 downto 377) => unused_tx_parallel_data(317 downto 317),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(378 downto 378) => unused_tx_parallel_data(318 downto 318),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(379 downto 379) => unused_tx_parallel_data(319 downto 319),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(380 downto 380) => unused_tx_parallel_data(320 downto 320),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(381 downto 381) => unused_tx_parallel_data(321 downto 321),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(382 downto 382) => unused_tx_parallel_data(322 downto 322),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(383 downto 383) => unused_tx_parallel_data(323 downto 323),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(384 downto 384) => tx_parallel_data(60 downto 60),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(385 downto 385) => tx_parallel_data(61 downto 61),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(386 downto 386) => tx_parallel_data(62 downto 62),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(387 downto 387) => tx_parallel_data(63 downto 63),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(388 downto 388) => tx_parallel_data(64 downto 64),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(389 downto 389) => tx_parallel_data(65 downto 65),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(390 downto 390) => tx_parallel_data(66 downto 66),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(391 downto 391) => tx_parallel_data(67 downto 67),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(392 downto 392) => tx_parallel_data(68 downto 68),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(393 downto 393) => tx_parallel_data(69 downto 69),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(394 downto 394) => unused_tx_parallel_data(324 downto 324),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(395 downto 395) => tx_parallel_data(70 downto 70),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(396 downto 396) => tx_parallel_data(71 downto 71),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(397 downto 397) => tx_parallel_data(72 downto 72),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(398 downto 398) => tx_parallel_data(73 downto 73),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(399 downto 399) => tx_parallel_data(74 downto 74),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(400 downto 400) => tx_parallel_data(75 downto 75),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(401 downto 401) => tx_parallel_data(76 downto 76),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(402 downto 402) => tx_parallel_data(77 downto 77),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(403 downto 403) => tx_parallel_data(78 downto 78),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(404 downto 404) => tx_parallel_data(79 downto 79),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(405 downto 405) => unused_tx_parallel_data(325 downto 325),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(406 downto 406) => unused_tx_parallel_data(326 downto 326),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(407 downto 407) => unused_tx_parallel_data(327 downto 327),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(408 downto 408) => unused_tx_parallel_data(328 downto 328),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(409 downto 409) => unused_tx_parallel_data(329 downto 329),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(410 downto 410) => unused_tx_parallel_data(330 downto 330),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(411 downto 411) => unused_tx_parallel_data(331 downto 331),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(412 downto 412) => unused_tx_parallel_data(332 downto 332),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(413 downto 413) => unused_tx_parallel_data(333 downto 333),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(414 downto 414) => unused_tx_parallel_data(334 downto 334),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(415 downto 415) => unused_tx_parallel_data(335 downto 335),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(416 downto 416) => unused_tx_parallel_data(336 downto 336),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(417 downto 417) => unused_tx_parallel_data(337 downto 337),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(418 downto 418) => unused_tx_parallel_data(338 downto 338),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(419 downto 419) => unused_tx_parallel_data(339 downto 339),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(420 downto 420) => unused_tx_parallel_data(340 downto 340),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(421 downto 421) => unused_tx_parallel_data(341 downto 341),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(422 downto 422) => unused_tx_parallel_data(342 downto 342),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(423 downto 423) => unused_tx_parallel_data(343 downto 343),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(424 downto 424) => unused_tx_parallel_data(344 downto 344),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(425 downto 425) => unused_tx_parallel_data(345 downto 345),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(426 downto 426) => unused_tx_parallel_data(346 downto 346),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(427 downto 427) => unused_tx_parallel_data(347 downto 347),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(428 downto 428) => unused_tx_parallel_data(348 downto 348),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(429 downto 429) => unused_tx_parallel_data(349 downto 349),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(430 downto 430) => unused_tx_parallel_data(350 downto 350),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(431 downto 431) => unused_tx_parallel_data(351 downto 351),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(432 downto 432) => unused_tx_parallel_data(352 downto 352),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(433 downto 433) => unused_tx_parallel_data(353 downto 353),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(434 downto 434) => unused_tx_parallel_data(354 downto 354),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(435 downto 435) => unused_tx_parallel_data(355 downto 355),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(436 downto 436) => unused_tx_parallel_data(356 downto 356),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(437 downto 437) => unused_tx_parallel_data(357 downto 357),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(438 downto 438) => unused_tx_parallel_data(358 downto 358),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(439 downto 439) => unused_tx_parallel_data(359 downto 359),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(440 downto 440) => unused_tx_parallel_data(360 downto 360),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(441 downto 441) => unused_tx_parallel_data(361 downto 361),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(442 downto 442) => unused_tx_parallel_data(362 downto 362),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(443 downto 443) => unused_tx_parallel_data(363 downto 363),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(444 downto 444) => unused_tx_parallel_data(364 downto 364),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(445 downto 445) => unused_tx_parallel_data(365 downto 365),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(446 downto 446) => unused_tx_parallel_data(366 downto 366),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(447 downto 447) => unused_tx_parallel_data(367 downto 367),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(448 downto 448) => unused_tx_parallel_data(368 downto 368),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(449 downto 449) => unused_tx_parallel_data(369 downto 369),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(450 downto 450) => unused_tx_parallel_data(370 downto 370),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(451 downto 451) => unused_tx_parallel_data(371 downto 371),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(452 downto 452) => unused_tx_parallel_data(372 downto 372),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(453 downto 453) => unused_tx_parallel_data(373 downto 373),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(454 downto 454) => unused_tx_parallel_data(374 downto 374),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(455 downto 455) => unused_tx_parallel_data(375 downto 375),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(456 downto 456) => unused_tx_parallel_data(376 downto 376),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(457 downto 457) => unused_tx_parallel_data(377 downto 377),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(458 downto 458) => unused_tx_parallel_data(378 downto 378),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(459 downto 459) => unused_tx_parallel_data(379 downto 379),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(460 downto 460) => unused_tx_parallel_data(380 downto 380),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(461 downto 461) => unused_tx_parallel_data(381 downto 381),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(462 downto 462) => unused_tx_parallel_data(382 downto 382),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(463 downto 463) => unused_tx_parallel_data(383 downto 383),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(464 downto 464) => unused_tx_parallel_data(384 downto 384),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(465 downto 465) => unused_tx_parallel_data(385 downto 385),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(466 downto 466) => unused_tx_parallel_data(386 downto 386),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(467 downto 467) => unused_tx_parallel_data(387 downto 387),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(468 downto 468) => unused_tx_parallel_data(388 downto 388),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(469 downto 469) => unused_tx_parallel_data(389 downto 389),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(470 downto 470) => unused_tx_parallel_data(390 downto 390),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(471 downto 471) => unused_tx_parallel_data(391 downto 391),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(472 downto 472) => unused_tx_parallel_data(392 downto 392),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(473 downto 473) => unused_tx_parallel_data(393 downto 393),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(474 downto 474) => unused_tx_parallel_data(394 downto 394),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(475 downto 475) => unused_tx_parallel_data(395 downto 395),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(476 downto 476) => unused_tx_parallel_data(396 downto 396),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(477 downto 477) => unused_tx_parallel_data(397 downto 397),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(478 downto 478) => unused_tx_parallel_data(398 downto 398),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(479 downto 479) => unused_tx_parallel_data(399 downto 399),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(480 downto 480) => unused_tx_parallel_data(400 downto 400),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(481 downto 481) => unused_tx_parallel_data(401 downto 401),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(482 downto 482) => unused_tx_parallel_data(402 downto 402),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(483 downto 483) => unused_tx_parallel_data(403 downto 403),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(484 downto 484) => unused_tx_parallel_data(404 downto 404),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(485 downto 485) => unused_tx_parallel_data(405 downto 405),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(486 downto 486) => unused_tx_parallel_data(406 downto 406),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(487 downto 487) => unused_tx_parallel_data(407 downto 407),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(488 downto 488) => unused_tx_parallel_data(408 downto 408),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(489 downto 489) => unused_tx_parallel_data(409 downto 409),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(490 downto 490) => unused_tx_parallel_data(410 downto 410),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(491 downto 491) => unused_tx_parallel_data(411 downto 411),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(492 downto 492) => unused_tx_parallel_data(412 downto 412),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(493 downto 493) => unused_tx_parallel_data(413 downto 413),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(494 downto 494) => unused_tx_parallel_data(414 downto 414),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(495 downto 495) => unused_tx_parallel_data(415 downto 415),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(496 downto 496) => unused_tx_parallel_data(416 downto 416),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(497 downto 497) => unused_tx_parallel_data(417 downto 417),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(498 downto 498) => unused_tx_parallel_data(418 downto 418),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(499 downto 499) => unused_tx_parallel_data(419 downto 419),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(500 downto 500) => unused_tx_parallel_data(420 downto 420),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(501 downto 501) => unused_tx_parallel_data(421 downto 421),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(502 downto 502) => unused_tx_parallel_data(422 downto 422),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(503 downto 503) => unused_tx_parallel_data(423 downto 423),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(504 downto 504) => unused_tx_parallel_data(424 downto 424),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(505 downto 505) => unused_tx_parallel_data(425 downto 425),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(506 downto 506) => unused_tx_parallel_data(426 downto 426),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(507 downto 507) => unused_tx_parallel_data(427 downto 427),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(508 downto 508) => unused_tx_parallel_data(428 downto 428),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(509 downto 509) => unused_tx_parallel_data(429 downto 429),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(510 downto 510) => unused_tx_parallel_data(430 downto 430),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(511 downto 511) => unused_tx_parallel_data(431 downto 431),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(512 downto 512) => tx_parallel_data(80 downto 80),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(513 downto 513) => tx_parallel_data(81 downto 81),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(514 downto 514) => tx_parallel_data(82 downto 82),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(515 downto 515) => tx_parallel_data(83 downto 83),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(516 downto 516) => tx_parallel_data(84 downto 84),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(517 downto 517) => tx_parallel_data(85 downto 85),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(518 downto 518) => tx_parallel_data(86 downto 86),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(519 downto 519) => tx_parallel_data(87 downto 87),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(520 downto 520) => tx_parallel_data(88 downto 88),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(521 downto 521) => tx_parallel_data(89 downto 89),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(522 downto 522) => unused_tx_parallel_data(432 downto 432),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(523 downto 523) => tx_parallel_data(90 downto 90),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(524 downto 524) => tx_parallel_data(91 downto 91),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(525 downto 525) => tx_parallel_data(92 downto 92),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(526 downto 526) => tx_parallel_data(93 downto 93),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(527 downto 527) => tx_parallel_data(94 downto 94),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(528 downto 528) => tx_parallel_data(95 downto 95),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(529 downto 529) => tx_parallel_data(96 downto 96),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(530 downto 530) => tx_parallel_data(97 downto 97),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(531 downto 531) => tx_parallel_data(98 downto 98),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(532 downto 532) => tx_parallel_data(99 downto 99),                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(533 downto 533) => unused_tx_parallel_data(433 downto 433),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(534 downto 534) => unused_tx_parallel_data(434 downto 434),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(535 downto 535) => unused_tx_parallel_data(435 downto 435),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(536 downto 536) => unused_tx_parallel_data(436 downto 436),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(537 downto 537) => unused_tx_parallel_data(437 downto 437),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(538 downto 538) => unused_tx_parallel_data(438 downto 438),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(539 downto 539) => unused_tx_parallel_data(439 downto 439),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(540 downto 540) => unused_tx_parallel_data(440 downto 440),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(541 downto 541) => unused_tx_parallel_data(441 downto 441),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(542 downto 542) => unused_tx_parallel_data(442 downto 442),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(543 downto 543) => unused_tx_parallel_data(443 downto 443),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(544 downto 544) => unused_tx_parallel_data(444 downto 444),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(545 downto 545) => unused_tx_parallel_data(445 downto 445),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(546 downto 546) => unused_tx_parallel_data(446 downto 446),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(547 downto 547) => unused_tx_parallel_data(447 downto 447),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(548 downto 548) => unused_tx_parallel_data(448 downto 448),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(549 downto 549) => unused_tx_parallel_data(449 downto 449),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(550 downto 550) => unused_tx_parallel_data(450 downto 450),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(551 downto 551) => unused_tx_parallel_data(451 downto 451),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(552 downto 552) => unused_tx_parallel_data(452 downto 452),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(553 downto 553) => unused_tx_parallel_data(453 downto 453),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(554 downto 554) => unused_tx_parallel_data(454 downto 454),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(555 downto 555) => unused_tx_parallel_data(455 downto 455),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(556 downto 556) => unused_tx_parallel_data(456 downto 456),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(557 downto 557) => unused_tx_parallel_data(457 downto 457),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(558 downto 558) => unused_tx_parallel_data(458 downto 458),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(559 downto 559) => unused_tx_parallel_data(459 downto 459),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(560 downto 560) => unused_tx_parallel_data(460 downto 460),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(561 downto 561) => unused_tx_parallel_data(461 downto 461),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(562 downto 562) => unused_tx_parallel_data(462 downto 462),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(563 downto 563) => unused_tx_parallel_data(463 downto 463),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(564 downto 564) => unused_tx_parallel_data(464 downto 464),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(565 downto 565) => unused_tx_parallel_data(465 downto 465),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(566 downto 566) => unused_tx_parallel_data(466 downto 466),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(567 downto 567) => unused_tx_parallel_data(467 downto 467),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(568 downto 568) => unused_tx_parallel_data(468 downto 468),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(569 downto 569) => unused_tx_parallel_data(469 downto 469),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(570 downto 570) => unused_tx_parallel_data(470 downto 470),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(571 downto 571) => unused_tx_parallel_data(471 downto 471),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(572 downto 572) => unused_tx_parallel_data(472 downto 472),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(573 downto 573) => unused_tx_parallel_data(473 downto 473),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(574 downto 574) => unused_tx_parallel_data(474 downto 474),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(575 downto 575) => unused_tx_parallel_data(475 downto 475),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(576 downto 576) => unused_tx_parallel_data(476 downto 476),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(577 downto 577) => unused_tx_parallel_data(477 downto 477),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(578 downto 578) => unused_tx_parallel_data(478 downto 478),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(579 downto 579) => unused_tx_parallel_data(479 downto 479),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(580 downto 580) => unused_tx_parallel_data(480 downto 480),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(581 downto 581) => unused_tx_parallel_data(481 downto 481),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(582 downto 582) => unused_tx_parallel_data(482 downto 482),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(583 downto 583) => unused_tx_parallel_data(483 downto 483),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(584 downto 584) => unused_tx_parallel_data(484 downto 484),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(585 downto 585) => unused_tx_parallel_data(485 downto 485),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(586 downto 586) => unused_tx_parallel_data(486 downto 486),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(587 downto 587) => unused_tx_parallel_data(487 downto 487),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(588 downto 588) => unused_tx_parallel_data(488 downto 488),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(589 downto 589) => unused_tx_parallel_data(489 downto 489),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(590 downto 590) => unused_tx_parallel_data(490 downto 490),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(591 downto 591) => unused_tx_parallel_data(491 downto 491),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(592 downto 592) => unused_tx_parallel_data(492 downto 492),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(593 downto 593) => unused_tx_parallel_data(493 downto 493),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(594 downto 594) => unused_tx_parallel_data(494 downto 494),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(595 downto 595) => unused_tx_parallel_data(495 downto 495),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(596 downto 596) => unused_tx_parallel_data(496 downto 496),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(597 downto 597) => unused_tx_parallel_data(497 downto 497),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(598 downto 598) => unused_tx_parallel_data(498 downto 498),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(599 downto 599) => unused_tx_parallel_data(499 downto 499),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(600 downto 600) => unused_tx_parallel_data(500 downto 500),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(601 downto 601) => unused_tx_parallel_data(501 downto 501),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(602 downto 602) => unused_tx_parallel_data(502 downto 502),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(603 downto 603) => unused_tx_parallel_data(503 downto 503),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(604 downto 604) => unused_tx_parallel_data(504 downto 504),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(605 downto 605) => unused_tx_parallel_data(505 downto 505),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(606 downto 606) => unused_tx_parallel_data(506 downto 506),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(607 downto 607) => unused_tx_parallel_data(507 downto 507),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(608 downto 608) => unused_tx_parallel_data(508 downto 508),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(609 downto 609) => unused_tx_parallel_data(509 downto 509),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(610 downto 610) => unused_tx_parallel_data(510 downto 510),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(611 downto 611) => unused_tx_parallel_data(511 downto 511),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(612 downto 612) => unused_tx_parallel_data(512 downto 512),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(613 downto 613) => unused_tx_parallel_data(513 downto 513),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(614 downto 614) => unused_tx_parallel_data(514 downto 514),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(615 downto 615) => unused_tx_parallel_data(515 downto 515),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(616 downto 616) => unused_tx_parallel_data(516 downto 516),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(617 downto 617) => unused_tx_parallel_data(517 downto 517),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(618 downto 618) => unused_tx_parallel_data(518 downto 518),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(619 downto 619) => unused_tx_parallel_data(519 downto 519),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(620 downto 620) => unused_tx_parallel_data(520 downto 520),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(621 downto 621) => unused_tx_parallel_data(521 downto 521),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(622 downto 622) => unused_tx_parallel_data(522 downto 522),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(623 downto 623) => unused_tx_parallel_data(523 downto 523),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(624 downto 624) => unused_tx_parallel_data(524 downto 524),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(625 downto 625) => unused_tx_parallel_data(525 downto 525),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(626 downto 626) => unused_tx_parallel_data(526 downto 526),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(627 downto 627) => unused_tx_parallel_data(527 downto 527),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(628 downto 628) => unused_tx_parallel_data(528 downto 528),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(629 downto 629) => unused_tx_parallel_data(529 downto 529),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(630 downto 630) => unused_tx_parallel_data(530 downto 530),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(631 downto 631) => unused_tx_parallel_data(531 downto 531),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(632 downto 632) => unused_tx_parallel_data(532 downto 532),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(633 downto 633) => unused_tx_parallel_data(533 downto 533),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(634 downto 634) => unused_tx_parallel_data(534 downto 534),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(635 downto 635) => unused_tx_parallel_data(535 downto 535),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(636 downto 636) => unused_tx_parallel_data(536 downto 536),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(637 downto 637) => unused_tx_parallel_data(537 downto 537),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(638 downto 638) => unused_tx_parallel_data(538 downto 538),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(639 downto 639) => unused_tx_parallel_data(539 downto 539),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(640 downto 640) => tx_parallel_data(100 downto 100),                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(641 downto 641) => tx_parallel_data(101 downto 101),                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(642 downto 642) => tx_parallel_data(102 downto 102),                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(643 downto 643) => tx_parallel_data(103 downto 103),                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(644 downto 644) => tx_parallel_data(104 downto 104),                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(645 downto 645) => tx_parallel_data(105 downto 105),                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(646 downto 646) => tx_parallel_data(106 downto 106),                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(647 downto 647) => tx_parallel_data(107 downto 107),                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(648 downto 648) => tx_parallel_data(108 downto 108),                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(649 downto 649) => tx_parallel_data(109 downto 109),                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(650 downto 650) => unused_tx_parallel_data(540 downto 540),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(651 downto 651) => tx_parallel_data(110 downto 110),                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(652 downto 652) => tx_parallel_data(111 downto 111),                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(653 downto 653) => tx_parallel_data(112 downto 112),                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(654 downto 654) => tx_parallel_data(113 downto 113),                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(655 downto 655) => tx_parallel_data(114 downto 114),                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(656 downto 656) => tx_parallel_data(115 downto 115),                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(657 downto 657) => tx_parallel_data(116 downto 116),                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(658 downto 658) => tx_parallel_data(117 downto 117),                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(659 downto 659) => tx_parallel_data(118 downto 118),                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(660 downto 660) => tx_parallel_data(119 downto 119),                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(661 downto 661) => unused_tx_parallel_data(541 downto 541),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(662 downto 662) => unused_tx_parallel_data(542 downto 542),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(663 downto 663) => unused_tx_parallel_data(543 downto 543),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(664 downto 664) => unused_tx_parallel_data(544 downto 544),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(665 downto 665) => unused_tx_parallel_data(545 downto 545),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(666 downto 666) => unused_tx_parallel_data(546 downto 546),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(667 downto 667) => unused_tx_parallel_data(547 downto 547),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(668 downto 668) => unused_tx_parallel_data(548 downto 548),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(669 downto 669) => unused_tx_parallel_data(549 downto 549),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(670 downto 670) => unused_tx_parallel_data(550 downto 550),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(671 downto 671) => unused_tx_parallel_data(551 downto 551),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(672 downto 672) => unused_tx_parallel_data(552 downto 552),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(673 downto 673) => unused_tx_parallel_data(553 downto 553),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(674 downto 674) => unused_tx_parallel_data(554 downto 554),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(675 downto 675) => unused_tx_parallel_data(555 downto 555),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(676 downto 676) => unused_tx_parallel_data(556 downto 556),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(677 downto 677) => unused_tx_parallel_data(557 downto 557),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(678 downto 678) => unused_tx_parallel_data(558 downto 558),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(679 downto 679) => unused_tx_parallel_data(559 downto 559),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(680 downto 680) => unused_tx_parallel_data(560 downto 560),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(681 downto 681) => unused_tx_parallel_data(561 downto 561),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(682 downto 682) => unused_tx_parallel_data(562 downto 562),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(683 downto 683) => unused_tx_parallel_data(563 downto 563),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(684 downto 684) => unused_tx_parallel_data(564 downto 564),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(685 downto 685) => unused_tx_parallel_data(565 downto 565),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(686 downto 686) => unused_tx_parallel_data(566 downto 566),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(687 downto 687) => unused_tx_parallel_data(567 downto 567),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(688 downto 688) => unused_tx_parallel_data(568 downto 568),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(689 downto 689) => unused_tx_parallel_data(569 downto 569),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(690 downto 690) => unused_tx_parallel_data(570 downto 570),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(691 downto 691) => unused_tx_parallel_data(571 downto 571),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(692 downto 692) => unused_tx_parallel_data(572 downto 572),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(693 downto 693) => unused_tx_parallel_data(573 downto 573),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(694 downto 694) => unused_tx_parallel_data(574 downto 574),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(695 downto 695) => unused_tx_parallel_data(575 downto 575),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(696 downto 696) => unused_tx_parallel_data(576 downto 576),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(697 downto 697) => unused_tx_parallel_data(577 downto 577),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(698 downto 698) => unused_tx_parallel_data(578 downto 578),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(699 downto 699) => unused_tx_parallel_data(579 downto 579),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(700 downto 700) => unused_tx_parallel_data(580 downto 580),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(701 downto 701) => unused_tx_parallel_data(581 downto 581),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(702 downto 702) => unused_tx_parallel_data(582 downto 582),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(703 downto 703) => unused_tx_parallel_data(583 downto 583),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(704 downto 704) => unused_tx_parallel_data(584 downto 584),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(705 downto 705) => unused_tx_parallel_data(585 downto 585),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(706 downto 706) => unused_tx_parallel_data(586 downto 586),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(707 downto 707) => unused_tx_parallel_data(587 downto 587),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(708 downto 708) => unused_tx_parallel_data(588 downto 588),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(709 downto 709) => unused_tx_parallel_data(589 downto 589),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(710 downto 710) => unused_tx_parallel_data(590 downto 590),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(711 downto 711) => unused_tx_parallel_data(591 downto 591),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(712 downto 712) => unused_tx_parallel_data(592 downto 592),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(713 downto 713) => unused_tx_parallel_data(593 downto 593),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(714 downto 714) => unused_tx_parallel_data(594 downto 594),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(715 downto 715) => unused_tx_parallel_data(595 downto 595),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(716 downto 716) => unused_tx_parallel_data(596 downto 596),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(717 downto 717) => unused_tx_parallel_data(597 downto 597),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(718 downto 718) => unused_tx_parallel_data(598 downto 598),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(719 downto 719) => unused_tx_parallel_data(599 downto 599),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(720 downto 720) => unused_tx_parallel_data(600 downto 600),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(721 downto 721) => unused_tx_parallel_data(601 downto 601),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(722 downto 722) => unused_tx_parallel_data(602 downto 602),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(723 downto 723) => unused_tx_parallel_data(603 downto 603),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(724 downto 724) => unused_tx_parallel_data(604 downto 604),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(725 downto 725) => unused_tx_parallel_data(605 downto 605),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(726 downto 726) => unused_tx_parallel_data(606 downto 606),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(727 downto 727) => unused_tx_parallel_data(607 downto 607),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(728 downto 728) => unused_tx_parallel_data(608 downto 608),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(729 downto 729) => unused_tx_parallel_data(609 downto 609),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(730 downto 730) => unused_tx_parallel_data(610 downto 610),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(731 downto 731) => unused_tx_parallel_data(611 downto 611),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(732 downto 732) => unused_tx_parallel_data(612 downto 612),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(733 downto 733) => unused_tx_parallel_data(613 downto 613),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(734 downto 734) => unused_tx_parallel_data(614 downto 614),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(735 downto 735) => unused_tx_parallel_data(615 downto 615),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(736 downto 736) => unused_tx_parallel_data(616 downto 616),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(737 downto 737) => unused_tx_parallel_data(617 downto 617),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(738 downto 738) => unused_tx_parallel_data(618 downto 618),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(739 downto 739) => unused_tx_parallel_data(619 downto 619),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(740 downto 740) => unused_tx_parallel_data(620 downto 620),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(741 downto 741) => unused_tx_parallel_data(621 downto 621),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(742 downto 742) => unused_tx_parallel_data(622 downto 622),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(743 downto 743) => unused_tx_parallel_data(623 downto 623),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(744 downto 744) => unused_tx_parallel_data(624 downto 624),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(745 downto 745) => unused_tx_parallel_data(625 downto 625),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(746 downto 746) => unused_tx_parallel_data(626 downto 626),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(747 downto 747) => unused_tx_parallel_data(627 downto 627),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(748 downto 748) => unused_tx_parallel_data(628 downto 628),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(749 downto 749) => unused_tx_parallel_data(629 downto 629),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(750 downto 750) => unused_tx_parallel_data(630 downto 630),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(751 downto 751) => unused_tx_parallel_data(631 downto 631),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(752 downto 752) => unused_tx_parallel_data(632 downto 632),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(753 downto 753) => unused_tx_parallel_data(633 downto 633),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(754 downto 754) => unused_tx_parallel_data(634 downto 634),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(755 downto 755) => unused_tx_parallel_data(635 downto 635),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(756 downto 756) => unused_tx_parallel_data(636 downto 636),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(757 downto 757) => unused_tx_parallel_data(637 downto 637),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(758 downto 758) => unused_tx_parallel_data(638 downto 638),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(759 downto 759) => unused_tx_parallel_data(639 downto 639),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(760 downto 760) => unused_tx_parallel_data(640 downto 640),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(761 downto 761) => unused_tx_parallel_data(641 downto 641),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(762 downto 762) => unused_tx_parallel_data(642 downto 642),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(763 downto 763) => unused_tx_parallel_data(643 downto 643),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(764 downto 764) => unused_tx_parallel_data(644 downto 644),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(765 downto 765) => unused_tx_parallel_data(645 downto 645),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(766 downto 766) => unused_tx_parallel_data(646 downto 646),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(767 downto 767) => unused_tx_parallel_data(647 downto 647),                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			rx_parallel_data                 => xcvr_native_a10_0_rx_parallel_data,                                                                                                                                                                                                                                                                                                                                                                 --   rx_parallel_data.rx_parallel_data
			tx_polinv                        => tx_polinv,                                                                                                                                                                                                                                                                                                                                                                                          --          tx_polinv.tx_polinv
			rx_polinv                        => rx_polinv,                                                                                                                                                                                                                                                                                                                                                                                          --          rx_polinv.rx_polinv
			reconfig_clk                     => reconfig_clk,                                                                                                                                                                                                                                                                                                                                                                                       --       reconfig_clk.clk
			reconfig_reset                   => reconfig_reset,                                                                                                                                                                                                                                                                                                                                                                                     --     reconfig_reset.reset
			reconfig_write                   => reconfig_write,                                                                                                                                                                                                                                                                                                                                                                                     --      reconfig_avmm.write
			reconfig_read                    => reconfig_read,                                                                                                                                                                                                                                                                                                                                                                                      --                   .read
			reconfig_address                 => reconfig_address,                                                                                                                                                                                                                                                                                                                                                                                   --                   .address
			reconfig_writedata               => reconfig_writedata,                                                                                                                                                                                                                                                                                                                                                                                 --                   .writedata
			reconfig_readdata                => reconfig_readdata,                                                                                                                                                                                                                                                                                                                                                                                  --                   .readdata
			reconfig_waitrequest             => reconfig_waitrequest,                                                                                                                                                                                                                                                                                                                                                                               --                   .waitrequest
			tx_analogreset_ack               => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_analogreset_ack               => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_serial_clk0                   => "000000",                                                                                                                                                                                                                                                                                                                                                                                           --        (terminated)
			tx_serial_clk1                   => "000000",                                                                                                                                                                                                                                                                                                                                                                                           --        (terminated)
			tx_serial_clk2                   => "000000",                                                                                                                                                                                                                                                                                                                                                                                           --        (terminated)
			tx_serial_clk3                   => "000000",                                                                                                                                                                                                                                                                                                                                                                                           --        (terminated)
			tx_bonding_clocks1               => "000000000000000000000000000000000000",                                                                                                                                                                                                                                                                                                                                                             --        (terminated)
			tx_bonding_clocks2               => "000000000000000000000000000000000000",                                                                                                                                                                                                                                                                                                                                                             --        (terminated)
			tx_bonding_clocks3               => "000000000000000000000000000000000000",                                                                                                                                                                                                                                                                                                                                                             --        (terminated)
			rx_cdr_refclk1                   => '0',                                                                                                                                                                                                                                                                                                                                                                                                --        (terminated)
			rx_cdr_refclk2                   => '0',                                                                                                                                                                                                                                                                                                                                                                                                --        (terminated)
			rx_cdr_refclk3                   => '0',                                                                                                                                                                                                                                                                                                                                                                                                --        (terminated)
			rx_cdr_refclk4                   => '0',                                                                                                                                                                                                                                                                                                                                                                                                --        (terminated)
			rx_pma_clkslip                   => "000000",                                                                                                                                                                                                                                                                                                                                                                                           --        (terminated)
			rx_set_locktodata                => "000000",                                                                                                                                                                                                                                                                                                                                                                                           --        (terminated)
			rx_set_locktoref                 => "000000",                                                                                                                                                                                                                                                                                                                                                                                           --        (terminated)
			rx_pma_qpipulldn                 => "000000",                                                                                                                                                                                                                                                                                                                                                                                           --        (terminated)
			tx_pma_qpipulldn                 => "000000",                                                                                                                                                                                                                                                                                                                                                                                           --        (terminated)
			tx_pma_qpipullup                 => "000000",                                                                                                                                                                                                                                                                                                                                                                                           --        (terminated)
			tx_pma_txdetectrx                => "000000",                                                                                                                                                                                                                                                                                                                                                                                           --        (terminated)
			tx_pma_elecidle                  => "000000",                                                                                                                                                                                                                                                                                                                                                                                           --        (terminated)
			tx_pma_rxfound                   => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_clklow                        => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_fref                          => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_pma_clkout                    => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_pma_div_clkout                => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_pma_iqtxrx_clkout             => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_pma_clkout                    => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_pma_div_clkout                => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_pma_iqtxrx_clkout             => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_control                       => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",                                                                                                                                                                                                                                                                                     --        (terminated)
			rx_control                       => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_bitslip                       => "000000",                                                                                                                                                                                                                                                                                                                                                                                           --        (terminated)
			rx_adapt_reset                   => "000000",                                                                                                                                                                                                                                                                                                                                                                                           --        (terminated)
			rx_adapt_start                   => "000000",                                                                                                                                                                                                                                                                                                                                                                                           --        (terminated)
			rx_prbs_err_clr                  => "000000",                                                                                                                                                                                                                                                                                                                                                                                           --        (terminated)
			rx_prbs_done                     => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_prbs_err                      => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_uhsif_clk                     => "000000",                                                                                                                                                                                                                                                                                                                                                                                           --        (terminated)
			tx_uhsif_clkout                  => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_uhsif_lock                    => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_std_pcfifo_full               => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_std_pcfifo_empty              => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_pcfifo_full               => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_pcfifo_empty              => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_bitrev_ena                => "000000",                                                                                                                                                                                                                                                                                                                                                                                           --        (terminated)
			rx_std_byterev_ena               => "000000",                                                                                                                                                                                                                                                                                                                                                                                           --        (terminated)
			tx_std_bitslipboundarysel        => "000000000000000000000000000000",                                                                                                                                                                                                                                                                                                                                                                   --        (terminated)
			rx_std_bitslipboundarysel        => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_wa_patternalign           => "000000",                                                                                                                                                                                                                                                                                                                                                                                           --        (terminated)
			rx_std_wa_a1a2size               => "000000",                                                                                                                                                                                                                                                                                                                                                                                           --        (terminated)
			rx_std_rmfifo_full               => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_rmfifo_empty              => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_signaldetect              => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_enh_data_valid                => "000000",                                                                                                                                                                                                                                                                                                                                                                                           --        (terminated)
			tx_enh_fifo_full                 => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_enh_fifo_pfull                => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_enh_fifo_empty                => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_enh_fifo_pempty               => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_enh_fifo_cnt                  => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_enh_fifo_rd_en                => "000000",                                                                                                                                                                                                                                                                                                                                                                                           --        (terminated)
			rx_enh_data_valid                => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_enh_fifo_full                 => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_enh_fifo_pfull                => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_enh_fifo_empty                => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_enh_fifo_pempty               => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_enh_fifo_del                  => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_enh_fifo_insert               => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_enh_fifo_cnt                  => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_enh_fifo_align_val            => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_enh_fifo_align_clr            => "000000",                                                                                                                                                                                                                                                                                                                                                                                           --        (terminated)
			tx_enh_frame                     => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_enh_frame_burst_en            => "000000",                                                                                                                                                                                                                                                                                                                                                                                           --        (terminated)
			tx_enh_frame_diag_status         => "000000000000",                                                                                                                                                                                                                                                                                                                                                                                     --        (terminated)
			rx_enh_frame                     => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_enh_frame_lock                => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_enh_frame_diag_status         => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_enh_crc32_err                 => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_enh_highber                   => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_enh_highber_clr_cnt           => "000000",                                                                                                                                                                                                                                                                                                                                                                                           --        (terminated)
			rx_enh_clr_errblk_count          => "000000",                                                                                                                                                                                                                                                                                                                                                                                           --        (terminated)
			rx_enh_blk_lock                  => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_enh_bitslip                   => "000000000000000000000000000000000000000000",                                                                                                                                                                                                                                                                                                                                                       --        (terminated)
			tx_hip_data                      => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", --        (terminated)
			rx_hip_data                      => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			hip_pipe_pclk                    => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			hip_fixedclk                     => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			hip_frefclk                      => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			hip_ctrl                         => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			hip_cal_done                     => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			pipe_rate                        => "00",                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			pipe_sw_done                     => "00",                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			pipe_sw                          => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			pipe_hclk_in                     => '0',                                                                                                                                                                                                                                                                                                                                                                                                --        (terminated)
			pipe_hclk_out                    => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			pipe_g3_txdeemph                 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",                                                                                                                                                                                                                                                                                     --        (terminated)
			pipe_g3_rxpresethint             => "000000000000000000",                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			pipe_rx_eidleinfersel            => "000000000000000000",                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			pipe_rx_elecidle                 => open,                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			pipe_rx_polarity                 => "000000",                                                                                                                                                                                                                                                                                                                                                                                           --        (terminated)
			avmm_busy                        => open                                                                                                                                                                                                                                                                                                                                                                                                --        (terminated)
		);

	rx_parallel_data <= xcvr_native_a10_0_rx_parallel_data(665 downto 665) & xcvr_native_a10_0_rx_parallel_data(664 downto 664) & xcvr_native_a10_0_rx_parallel_data(663 downto 663) & xcvr_native_a10_0_rx_parallel_data(662 downto 662) & xcvr_native_a10_0_rx_parallel_data(661 downto 661) & xcvr_native_a10_0_rx_parallel_data(660 downto 660) & xcvr_native_a10_0_rx_parallel_data(659 downto 659) & xcvr_native_a10_0_rx_parallel_data(658 downto 658) & xcvr_native_a10_0_rx_parallel_data(657 downto 657) & xcvr_native_a10_0_rx_parallel_data(656 downto 656) & xcvr_native_a10_0_rx_parallel_data(649 downto 649) & xcvr_native_a10_0_rx_parallel_data(648 downto 648) & xcvr_native_a10_0_rx_parallel_data(647 downto 647) & xcvr_native_a10_0_rx_parallel_data(646 downto 646) & xcvr_native_a10_0_rx_parallel_data(645 downto 645) & xcvr_native_a10_0_rx_parallel_data(644 downto 644) & xcvr_native_a10_0_rx_parallel_data(643 downto 643) & xcvr_native_a10_0_rx_parallel_data(642 downto 642) & xcvr_native_a10_0_rx_parallel_data(641 downto 641) & xcvr_native_a10_0_rx_parallel_data(640 downto 640) & xcvr_native_a10_0_rx_parallel_data(537 downto 537) & xcvr_native_a10_0_rx_parallel_data(536 downto 536) & xcvr_native_a10_0_rx_parallel_data(535 downto 535) & xcvr_native_a10_0_rx_parallel_data(534 downto 534) & xcvr_native_a10_0_rx_parallel_data(533 downto 533) & xcvr_native_a10_0_rx_parallel_data(532 downto 532) & xcvr_native_a10_0_rx_parallel_data(531 downto 531) & xcvr_native_a10_0_rx_parallel_data(530 downto 530) & xcvr_native_a10_0_rx_parallel_data(529 downto 529) & xcvr_native_a10_0_rx_parallel_data(528 downto 528) & xcvr_native_a10_0_rx_parallel_data(521 downto 521) & xcvr_native_a10_0_rx_parallel_data(520 downto 520) & xcvr_native_a10_0_rx_parallel_data(519 downto 519) & xcvr_native_a10_0_rx_parallel_data(518 downto 518) & xcvr_native_a10_0_rx_parallel_data(517 downto 517) & xcvr_native_a10_0_rx_parallel_data(516 downto 516) & xcvr_native_a10_0_rx_parallel_data(515 downto 515) & xcvr_native_a10_0_rx_parallel_data(514 downto 514) & xcvr_native_a10_0_rx_parallel_data(513 downto 513) & xcvr_native_a10_0_rx_parallel_data(512 downto 512) & xcvr_native_a10_0_rx_parallel_data(409 downto 409) & xcvr_native_a10_0_rx_parallel_data(408 downto 408) & xcvr_native_a10_0_rx_parallel_data(407 downto 407) & xcvr_native_a10_0_rx_parallel_data(406 downto 406) & xcvr_native_a10_0_rx_parallel_data(405 downto 405) & xcvr_native_a10_0_rx_parallel_data(404 downto 404) & xcvr_native_a10_0_rx_parallel_data(403 downto 403) & xcvr_native_a10_0_rx_parallel_data(402 downto 402) & xcvr_native_a10_0_rx_parallel_data(401 downto 401) & xcvr_native_a10_0_rx_parallel_data(400 downto 400) & xcvr_native_a10_0_rx_parallel_data(393 downto 393) & xcvr_native_a10_0_rx_parallel_data(392 downto 392) & xcvr_native_a10_0_rx_parallel_data(391 downto 391) & xcvr_native_a10_0_rx_parallel_data(390 downto 390) & xcvr_native_a10_0_rx_parallel_data(389 downto 389) & xcvr_native_a10_0_rx_parallel_data(388 downto 388) & xcvr_native_a10_0_rx_parallel_data(387 downto 387) & xcvr_native_a10_0_rx_parallel_data(386 downto 386) & xcvr_native_a10_0_rx_parallel_data(385 downto 385) & xcvr_native_a10_0_rx_parallel_data(384 downto 384) & xcvr_native_a10_0_rx_parallel_data(281 downto 281) & xcvr_native_a10_0_rx_parallel_data(280 downto 280) & xcvr_native_a10_0_rx_parallel_data(279 downto 279) & xcvr_native_a10_0_rx_parallel_data(278 downto 278) & xcvr_native_a10_0_rx_parallel_data(277 downto 277) & xcvr_native_a10_0_rx_parallel_data(276 downto 276) & xcvr_native_a10_0_rx_parallel_data(275 downto 275) & xcvr_native_a10_0_rx_parallel_data(274 downto 274) & xcvr_native_a10_0_rx_parallel_data(273 downto 273) & xcvr_native_a10_0_rx_parallel_data(272 downto 272) & xcvr_native_a10_0_rx_parallel_data(265 downto 265) & xcvr_native_a10_0_rx_parallel_data(264 downto 264) & xcvr_native_a10_0_rx_parallel_data(263 downto 263) & xcvr_native_a10_0_rx_parallel_data(262 downto 262) & xcvr_native_a10_0_rx_parallel_data(261 downto 261) & xcvr_native_a10_0_rx_parallel_data(260 downto 260) & xcvr_native_a10_0_rx_parallel_data(259 downto 259) & xcvr_native_a10_0_rx_parallel_data(258 downto 258) & xcvr_native_a10_0_rx_parallel_data(257 downto 257) & xcvr_native_a10_0_rx_parallel_data(256 downto 256) & xcvr_native_a10_0_rx_parallel_data(153 downto 153) & xcvr_native_a10_0_rx_parallel_data(152 downto 152) & xcvr_native_a10_0_rx_parallel_data(151 downto 151) & xcvr_native_a10_0_rx_parallel_data(150 downto 150) & xcvr_native_a10_0_rx_parallel_data(149 downto 149) & xcvr_native_a10_0_rx_parallel_data(148 downto 148) & xcvr_native_a10_0_rx_parallel_data(147 downto 147) & xcvr_native_a10_0_rx_parallel_data(146 downto 146) & xcvr_native_a10_0_rx_parallel_data(145 downto 145) & xcvr_native_a10_0_rx_parallel_data(144 downto 144) & xcvr_native_a10_0_rx_parallel_data(137 downto 137) & xcvr_native_a10_0_rx_parallel_data(136 downto 136) & xcvr_native_a10_0_rx_parallel_data(135 downto 135) & xcvr_native_a10_0_rx_parallel_data(134 downto 134) & xcvr_native_a10_0_rx_parallel_data(133 downto 133) & xcvr_native_a10_0_rx_parallel_data(132 downto 132) & xcvr_native_a10_0_rx_parallel_data(131 downto 131) & xcvr_native_a10_0_rx_parallel_data(130 downto 130) & xcvr_native_a10_0_rx_parallel_data(129 downto 129) & xcvr_native_a10_0_rx_parallel_data(128 downto 128) & xcvr_native_a10_0_rx_parallel_data(25 downto 25) & xcvr_native_a10_0_rx_parallel_data(24 downto 24) & xcvr_native_a10_0_rx_parallel_data(23 downto 23) & xcvr_native_a10_0_rx_parallel_data(22 downto 22) & xcvr_native_a10_0_rx_parallel_data(21 downto 21) & xcvr_native_a10_0_rx_parallel_data(20 downto 20) & xcvr_native_a10_0_rx_parallel_data(19 downto 19) & xcvr_native_a10_0_rx_parallel_data(18 downto 18) & xcvr_native_a10_0_rx_parallel_data(17 downto 17) & xcvr_native_a10_0_rx_parallel_data(16 downto 16) & xcvr_native_a10_0_rx_parallel_data(9 downto 9) & xcvr_native_a10_0_rx_parallel_data(8 downto 8) & xcvr_native_a10_0_rx_parallel_data(7 downto 7) & xcvr_native_a10_0_rx_parallel_data(6 downto 6) & xcvr_native_a10_0_rx_parallel_data(5 downto 5) & xcvr_native_a10_0_rx_parallel_data(4 downto 4) & xcvr_native_a10_0_rx_parallel_data(3 downto 3) & xcvr_native_a10_0_rx_parallel_data(2 downto 2) & xcvr_native_a10_0_rx_parallel_data(1 downto 1) & xcvr_native_a10_0_rx_parallel_data(0 downto 0);

	unused_rx_parallel_data <= xcvr_native_a10_0_rx_parallel_data(767 downto 767) & xcvr_native_a10_0_rx_parallel_data(766 downto 766) & xcvr_native_a10_0_rx_parallel_data(765 downto 765) & xcvr_native_a10_0_rx_parallel_data(764 downto 764) & xcvr_native_a10_0_rx_parallel_data(763 downto 763) & xcvr_native_a10_0_rx_parallel_data(762 downto 762) & xcvr_native_a10_0_rx_parallel_data(761 downto 761) & xcvr_native_a10_0_rx_parallel_data(760 downto 760) & xcvr_native_a10_0_rx_parallel_data(759 downto 759) & xcvr_native_a10_0_rx_parallel_data(758 downto 758) & xcvr_native_a10_0_rx_parallel_data(757 downto 757) & xcvr_native_a10_0_rx_parallel_data(756 downto 756) & xcvr_native_a10_0_rx_parallel_data(755 downto 755) & xcvr_native_a10_0_rx_parallel_data(754 downto 754) & xcvr_native_a10_0_rx_parallel_data(753 downto 753) & xcvr_native_a10_0_rx_parallel_data(752 downto 752) & xcvr_native_a10_0_rx_parallel_data(751 downto 751) & xcvr_native_a10_0_rx_parallel_data(750 downto 750) & xcvr_native_a10_0_rx_parallel_data(749 downto 749) & xcvr_native_a10_0_rx_parallel_data(748 downto 748) & xcvr_native_a10_0_rx_parallel_data(747 downto 747) & xcvr_native_a10_0_rx_parallel_data(746 downto 746) & xcvr_native_a10_0_rx_parallel_data(745 downto 745) & xcvr_native_a10_0_rx_parallel_data(744 downto 744) & xcvr_native_a10_0_rx_parallel_data(743 downto 743) & xcvr_native_a10_0_rx_parallel_data(742 downto 742) & xcvr_native_a10_0_rx_parallel_data(741 downto 741) & xcvr_native_a10_0_rx_parallel_data(740 downto 740) & xcvr_native_a10_0_rx_parallel_data(739 downto 739) & xcvr_native_a10_0_rx_parallel_data(738 downto 738) & xcvr_native_a10_0_rx_parallel_data(737 downto 737) & xcvr_native_a10_0_rx_parallel_data(736 downto 736) & xcvr_native_a10_0_rx_parallel_data(735 downto 735) & xcvr_native_a10_0_rx_parallel_data(734 downto 734) & xcvr_native_a10_0_rx_parallel_data(733 downto 733) & xcvr_native_a10_0_rx_parallel_data(732 downto 732) & xcvr_native_a10_0_rx_parallel_data(731 downto 731) & xcvr_native_a10_0_rx_parallel_data(730 downto 730) & xcvr_native_a10_0_rx_parallel_data(729 downto 729) & xcvr_native_a10_0_rx_parallel_data(728 downto 728) & xcvr_native_a10_0_rx_parallel_data(727 downto 727) & xcvr_native_a10_0_rx_parallel_data(726 downto 726) & xcvr_native_a10_0_rx_parallel_data(725 downto 725) & xcvr_native_a10_0_rx_parallel_data(724 downto 724) & xcvr_native_a10_0_rx_parallel_data(723 downto 723) & xcvr_native_a10_0_rx_parallel_data(722 downto 722) & xcvr_native_a10_0_rx_parallel_data(721 downto 721) & xcvr_native_a10_0_rx_parallel_data(720 downto 720) & xcvr_native_a10_0_rx_parallel_data(719 downto 719) & xcvr_native_a10_0_rx_parallel_data(718 downto 718) & xcvr_native_a10_0_rx_parallel_data(717 downto 717) & xcvr_native_a10_0_rx_parallel_data(716 downto 716) & xcvr_native_a10_0_rx_parallel_data(715 downto 715) & xcvr_native_a10_0_rx_parallel_data(714 downto 714) & xcvr_native_a10_0_rx_parallel_data(713 downto 713) & xcvr_native_a10_0_rx_parallel_data(712 downto 712) & xcvr_native_a10_0_rx_parallel_data(711 downto 711) & xcvr_native_a10_0_rx_parallel_data(710 downto 710) & xcvr_native_a10_0_rx_parallel_data(709 downto 709) & xcvr_native_a10_0_rx_parallel_data(708 downto 708) & xcvr_native_a10_0_rx_parallel_data(707 downto 707) & xcvr_native_a10_0_rx_parallel_data(706 downto 706) & xcvr_native_a10_0_rx_parallel_data(705 downto 705) & xcvr_native_a10_0_rx_parallel_data(704 downto 704) & xcvr_native_a10_0_rx_parallel_data(703 downto 703) & xcvr_native_a10_0_rx_parallel_data(702 downto 702) & xcvr_native_a10_0_rx_parallel_data(701 downto 701) & xcvr_native_a10_0_rx_parallel_data(700 downto 700) & xcvr_native_a10_0_rx_parallel_data(699 downto 699) & xcvr_native_a10_0_rx_parallel_data(698 downto 698) & xcvr_native_a10_0_rx_parallel_data(697 downto 697) & xcvr_native_a10_0_rx_parallel_data(696 downto 696) & xcvr_native_a10_0_rx_parallel_data(695 downto 695) & xcvr_native_a10_0_rx_parallel_data(694 downto 694) & xcvr_native_a10_0_rx_parallel_data(693 downto 693) & xcvr_native_a10_0_rx_parallel_data(692 downto 692) & xcvr_native_a10_0_rx_parallel_data(691 downto 691) & xcvr_native_a10_0_rx_parallel_data(690 downto 690) & xcvr_native_a10_0_rx_parallel_data(689 downto 689) & xcvr_native_a10_0_rx_parallel_data(688 downto 688) & xcvr_native_a10_0_rx_parallel_data(687 downto 687) & xcvr_native_a10_0_rx_parallel_data(686 downto 686) & xcvr_native_a10_0_rx_parallel_data(685 downto 685) & xcvr_native_a10_0_rx_parallel_data(684 downto 684) & xcvr_native_a10_0_rx_parallel_data(683 downto 683) & xcvr_native_a10_0_rx_parallel_data(682 downto 682) & xcvr_native_a10_0_rx_parallel_data(681 downto 681) & xcvr_native_a10_0_rx_parallel_data(680 downto 680) & xcvr_native_a10_0_rx_parallel_data(679 downto 679) & xcvr_native_a10_0_rx_parallel_data(678 downto 678) & xcvr_native_a10_0_rx_parallel_data(677 downto 677) & xcvr_native_a10_0_rx_parallel_data(676 downto 676) & xcvr_native_a10_0_rx_parallel_data(675 downto 675) & xcvr_native_a10_0_rx_parallel_data(674 downto 674) & xcvr_native_a10_0_rx_parallel_data(673 downto 673) & xcvr_native_a10_0_rx_parallel_data(672 downto 672) & xcvr_native_a10_0_rx_parallel_data(671 downto 671) & xcvr_native_a10_0_rx_parallel_data(670 downto 670) & xcvr_native_a10_0_rx_parallel_data(669 downto 669) & xcvr_native_a10_0_rx_parallel_data(668 downto 668) & xcvr_native_a10_0_rx_parallel_data(667 downto 667) & xcvr_native_a10_0_rx_parallel_data(666 downto 666) & xcvr_native_a10_0_rx_parallel_data(655 downto 655) & xcvr_native_a10_0_rx_parallel_data(654 downto 654) & xcvr_native_a10_0_rx_parallel_data(653 downto 653) & xcvr_native_a10_0_rx_parallel_data(652 downto 652) & xcvr_native_a10_0_rx_parallel_data(651 downto 651) & xcvr_native_a10_0_rx_parallel_data(650 downto 650) & xcvr_native_a10_0_rx_parallel_data(639 downto 639) & xcvr_native_a10_0_rx_parallel_data(638 downto 638) & xcvr_native_a10_0_rx_parallel_data(637 downto 637) & xcvr_native_a10_0_rx_parallel_data(636 downto 636) & xcvr_native_a10_0_rx_parallel_data(635 downto 635) & xcvr_native_a10_0_rx_parallel_data(634 downto 634) & xcvr_native_a10_0_rx_parallel_data(633 downto 633) & xcvr_native_a10_0_rx_parallel_data(632 downto 632) & xcvr_native_a10_0_rx_parallel_data(631 downto 631) & xcvr_native_a10_0_rx_parallel_data(630 downto 630) & xcvr_native_a10_0_rx_parallel_data(629 downto 629) & xcvr_native_a10_0_rx_parallel_data(628 downto 628) & xcvr_native_a10_0_rx_parallel_data(627 downto 627) & xcvr_native_a10_0_rx_parallel_data(626 downto 626) & xcvr_native_a10_0_rx_parallel_data(625 downto 625) & xcvr_native_a10_0_rx_parallel_data(624 downto 624) & xcvr_native_a10_0_rx_parallel_data(623 downto 623) & xcvr_native_a10_0_rx_parallel_data(622 downto 622) & xcvr_native_a10_0_rx_parallel_data(621 downto 621) & xcvr_native_a10_0_rx_parallel_data(620 downto 620) & xcvr_native_a10_0_rx_parallel_data(619 downto 619) & xcvr_native_a10_0_rx_parallel_data(618 downto 618) & xcvr_native_a10_0_rx_parallel_data(617 downto 617) & xcvr_native_a10_0_rx_parallel_data(616 downto 616) & xcvr_native_a10_0_rx_parallel_data(615 downto 615) & xcvr_native_a10_0_rx_parallel_data(614 downto 614) & xcvr_native_a10_0_rx_parallel_data(613 downto 613) & xcvr_native_a10_0_rx_parallel_data(612 downto 612) & xcvr_native_a10_0_rx_parallel_data(611 downto 611) & xcvr_native_a10_0_rx_parallel_data(610 downto 610) & xcvr_native_a10_0_rx_parallel_data(609 downto 609) & xcvr_native_a10_0_rx_parallel_data(608 downto 608) & xcvr_native_a10_0_rx_parallel_data(607 downto 607) & xcvr_native_a10_0_rx_parallel_data(606 downto 606) & xcvr_native_a10_0_rx_parallel_data(605 downto 605) & xcvr_native_a10_0_rx_parallel_data(604 downto 604) & xcvr_native_a10_0_rx_parallel_data(603 downto 603) & xcvr_native_a10_0_rx_parallel_data(602 downto 602) & xcvr_native_a10_0_rx_parallel_data(601 downto 601) & xcvr_native_a10_0_rx_parallel_data(600 downto 600) & xcvr_native_a10_0_rx_parallel_data(599 downto 599) & xcvr_native_a10_0_rx_parallel_data(598 downto 598) & xcvr_native_a10_0_rx_parallel_data(597 downto 597) & xcvr_native_a10_0_rx_parallel_data(596 downto 596) & xcvr_native_a10_0_rx_parallel_data(595 downto 595) & xcvr_native_a10_0_rx_parallel_data(594 downto 594) & xcvr_native_a10_0_rx_parallel_data(593 downto 593) & xcvr_native_a10_0_rx_parallel_data(592 downto 592) & xcvr_native_a10_0_rx_parallel_data(591 downto 591) & xcvr_native_a10_0_rx_parallel_data(590 downto 590) & xcvr_native_a10_0_rx_parallel_data(589 downto 589) & xcvr_native_a10_0_rx_parallel_data(588 downto 588) & xcvr_native_a10_0_rx_parallel_data(587 downto 587) & xcvr_native_a10_0_rx_parallel_data(586 downto 586) & xcvr_native_a10_0_rx_parallel_data(585 downto 585) & xcvr_native_a10_0_rx_parallel_data(584 downto 584) & xcvr_native_a10_0_rx_parallel_data(583 downto 583) & xcvr_native_a10_0_rx_parallel_data(582 downto 582) & xcvr_native_a10_0_rx_parallel_data(581 downto 581) & xcvr_native_a10_0_rx_parallel_data(580 downto 580) & xcvr_native_a10_0_rx_parallel_data(579 downto 579) & xcvr_native_a10_0_rx_parallel_data(578 downto 578) & xcvr_native_a10_0_rx_parallel_data(577 downto 577) & xcvr_native_a10_0_rx_parallel_data(576 downto 576) & xcvr_native_a10_0_rx_parallel_data(575 downto 575) & xcvr_native_a10_0_rx_parallel_data(574 downto 574) & xcvr_native_a10_0_rx_parallel_data(573 downto 573) & xcvr_native_a10_0_rx_parallel_data(572 downto 572) & xcvr_native_a10_0_rx_parallel_data(571 downto 571) & xcvr_native_a10_0_rx_parallel_data(570 downto 570) & xcvr_native_a10_0_rx_parallel_data(569 downto 569) & xcvr_native_a10_0_rx_parallel_data(568 downto 568) & xcvr_native_a10_0_rx_parallel_data(567 downto 567) & xcvr_native_a10_0_rx_parallel_data(566 downto 566) & xcvr_native_a10_0_rx_parallel_data(565 downto 565) & xcvr_native_a10_0_rx_parallel_data(564 downto 564) & xcvr_native_a10_0_rx_parallel_data(563 downto 563) & xcvr_native_a10_0_rx_parallel_data(562 downto 562) & xcvr_native_a10_0_rx_parallel_data(561 downto 561) & xcvr_native_a10_0_rx_parallel_data(560 downto 560) & xcvr_native_a10_0_rx_parallel_data(559 downto 559) & xcvr_native_a10_0_rx_parallel_data(558 downto 558) & xcvr_native_a10_0_rx_parallel_data(557 downto 557) & xcvr_native_a10_0_rx_parallel_data(556 downto 556) & xcvr_native_a10_0_rx_parallel_data(555 downto 555) & xcvr_native_a10_0_rx_parallel_data(554 downto 554) & xcvr_native_a10_0_rx_parallel_data(553 downto 553) & xcvr_native_a10_0_rx_parallel_data(552 downto 552) & xcvr_native_a10_0_rx_parallel_data(551 downto 551) & xcvr_native_a10_0_rx_parallel_data(550 downto 550) & xcvr_native_a10_0_rx_parallel_data(549 downto 549) & xcvr_native_a10_0_rx_parallel_data(548 downto 548) & xcvr_native_a10_0_rx_parallel_data(547 downto 547) & xcvr_native_a10_0_rx_parallel_data(546 downto 546) & xcvr_native_a10_0_rx_parallel_data(545 downto 545) & xcvr_native_a10_0_rx_parallel_data(544 downto 544) & xcvr_native_a10_0_rx_parallel_data(543 downto 543) & xcvr_native_a10_0_rx_parallel_data(542 downto 542) & xcvr_native_a10_0_rx_parallel_data(541 downto 541) & xcvr_native_a10_0_rx_parallel_data(540 downto 540) & xcvr_native_a10_0_rx_parallel_data(539 downto 539) & xcvr_native_a10_0_rx_parallel_data(538 downto 538) & xcvr_native_a10_0_rx_parallel_data(527 downto 527) & xcvr_native_a10_0_rx_parallel_data(526 downto 526) & xcvr_native_a10_0_rx_parallel_data(525 downto 525) & xcvr_native_a10_0_rx_parallel_data(524 downto 524) & xcvr_native_a10_0_rx_parallel_data(523 downto 523) & xcvr_native_a10_0_rx_parallel_data(522 downto 522) & xcvr_native_a10_0_rx_parallel_data(511 downto 511) & xcvr_native_a10_0_rx_parallel_data(510 downto 510) & xcvr_native_a10_0_rx_parallel_data(509 downto 509) & xcvr_native_a10_0_rx_parallel_data(508 downto 508) & xcvr_native_a10_0_rx_parallel_data(507 downto 507) & xcvr_native_a10_0_rx_parallel_data(506 downto 506) & xcvr_native_a10_0_rx_parallel_data(505 downto 505) & xcvr_native_a10_0_rx_parallel_data(504 downto 504) & xcvr_native_a10_0_rx_parallel_data(503 downto 503) & xcvr_native_a10_0_rx_parallel_data(502 downto 502) & xcvr_native_a10_0_rx_parallel_data(501 downto 501) & xcvr_native_a10_0_rx_parallel_data(500 downto 500) & xcvr_native_a10_0_rx_parallel_data(499 downto 499) & xcvr_native_a10_0_rx_parallel_data(498 downto 498) & xcvr_native_a10_0_rx_parallel_data(497 downto 497) & xcvr_native_a10_0_rx_parallel_data(496 downto 496) & xcvr_native_a10_0_rx_parallel_data(495 downto 495) & xcvr_native_a10_0_rx_parallel_data(494 downto 494) & xcvr_native_a10_0_rx_parallel_data(493 downto 493) & xcvr_native_a10_0_rx_parallel_data(492 downto 492) & xcvr_native_a10_0_rx_parallel_data(491 downto 491) & xcvr_native_a10_0_rx_parallel_data(490 downto 490) & xcvr_native_a10_0_rx_parallel_data(489 downto 489) & xcvr_native_a10_0_rx_parallel_data(488 downto 488) & xcvr_native_a10_0_rx_parallel_data(487 downto 487) & xcvr_native_a10_0_rx_parallel_data(486 downto 486) & xcvr_native_a10_0_rx_parallel_data(485 downto 485) & xcvr_native_a10_0_rx_parallel_data(484 downto 484) & xcvr_native_a10_0_rx_parallel_data(483 downto 483) & xcvr_native_a10_0_rx_parallel_data(482 downto 482) & xcvr_native_a10_0_rx_parallel_data(481 downto 481) & xcvr_native_a10_0_rx_parallel_data(480 downto 480) & xcvr_native_a10_0_rx_parallel_data(479 downto 479) & xcvr_native_a10_0_rx_parallel_data(478 downto 478) & xcvr_native_a10_0_rx_parallel_data(477 downto 477) & xcvr_native_a10_0_rx_parallel_data(476 downto 476) & xcvr_native_a10_0_rx_parallel_data(475 downto 475) & xcvr_native_a10_0_rx_parallel_data(474 downto 474) & xcvr_native_a10_0_rx_parallel_data(473 downto 473) & xcvr_native_a10_0_rx_parallel_data(472 downto 472) & xcvr_native_a10_0_rx_parallel_data(471 downto 471) & xcvr_native_a10_0_rx_parallel_data(470 downto 470) & xcvr_native_a10_0_rx_parallel_data(469 downto 469) & xcvr_native_a10_0_rx_parallel_data(468 downto 468) & xcvr_native_a10_0_rx_parallel_data(467 downto 467) & xcvr_native_a10_0_rx_parallel_data(466 downto 466) & xcvr_native_a10_0_rx_parallel_data(465 downto 465) & xcvr_native_a10_0_rx_parallel_data(464 downto 464) & xcvr_native_a10_0_rx_parallel_data(463 downto 463) & xcvr_native_a10_0_rx_parallel_data(462 downto 462) & xcvr_native_a10_0_rx_parallel_data(461 downto 461) & xcvr_native_a10_0_rx_parallel_data(460 downto 460) & xcvr_native_a10_0_rx_parallel_data(459 downto 459) & xcvr_native_a10_0_rx_parallel_data(458 downto 458) & xcvr_native_a10_0_rx_parallel_data(457 downto 457) & xcvr_native_a10_0_rx_parallel_data(456 downto 456) & xcvr_native_a10_0_rx_parallel_data(455 downto 455) & xcvr_native_a10_0_rx_parallel_data(454 downto 454) & xcvr_native_a10_0_rx_parallel_data(453 downto 453) & xcvr_native_a10_0_rx_parallel_data(452 downto 452) & xcvr_native_a10_0_rx_parallel_data(451 downto 451) & xcvr_native_a10_0_rx_parallel_data(450 downto 450) & xcvr_native_a10_0_rx_parallel_data(449 downto 449) & xcvr_native_a10_0_rx_parallel_data(448 downto 448) & xcvr_native_a10_0_rx_parallel_data(447 downto 447) & xcvr_native_a10_0_rx_parallel_data(446 downto 446) & xcvr_native_a10_0_rx_parallel_data(445 downto 445) & xcvr_native_a10_0_rx_parallel_data(444 downto 444) & xcvr_native_a10_0_rx_parallel_data(443 downto 443) & xcvr_native_a10_0_rx_parallel_data(442 downto 442) & xcvr_native_a10_0_rx_parallel_data(441 downto 441) & xcvr_native_a10_0_rx_parallel_data(440 downto 440) & xcvr_native_a10_0_rx_parallel_data(439 downto 439) & xcvr_native_a10_0_rx_parallel_data(438 downto 438) & xcvr_native_a10_0_rx_parallel_data(437 downto 437) & xcvr_native_a10_0_rx_parallel_data(436 downto 436) & xcvr_native_a10_0_rx_parallel_data(435 downto 435) & xcvr_native_a10_0_rx_parallel_data(434 downto 434) & xcvr_native_a10_0_rx_parallel_data(433 downto 433) & xcvr_native_a10_0_rx_parallel_data(432 downto 432) & xcvr_native_a10_0_rx_parallel_data(431 downto 431) & xcvr_native_a10_0_rx_parallel_data(430 downto 430) & xcvr_native_a10_0_rx_parallel_data(429 downto 429) & xcvr_native_a10_0_rx_parallel_data(428 downto 428) & xcvr_native_a10_0_rx_parallel_data(427 downto 427) & xcvr_native_a10_0_rx_parallel_data(426 downto 426) & xcvr_native_a10_0_rx_parallel_data(425 downto 425) & xcvr_native_a10_0_rx_parallel_data(424 downto 424) & xcvr_native_a10_0_rx_parallel_data(423 downto 423) & xcvr_native_a10_0_rx_parallel_data(422 downto 422) & xcvr_native_a10_0_rx_parallel_data(421 downto 421) & xcvr_native_a10_0_rx_parallel_data(420 downto 420) & xcvr_native_a10_0_rx_parallel_data(419 downto 419) & xcvr_native_a10_0_rx_parallel_data(418 downto 418) & xcvr_native_a10_0_rx_parallel_data(417 downto 417) & xcvr_native_a10_0_rx_parallel_data(416 downto 416) & xcvr_native_a10_0_rx_parallel_data(415 downto 415) & xcvr_native_a10_0_rx_parallel_data(414 downto 414) & xcvr_native_a10_0_rx_parallel_data(413 downto 413) & xcvr_native_a10_0_rx_parallel_data(412 downto 412) & xcvr_native_a10_0_rx_parallel_data(411 downto 411) & xcvr_native_a10_0_rx_parallel_data(410 downto 410) & xcvr_native_a10_0_rx_parallel_data(399 downto 399) & xcvr_native_a10_0_rx_parallel_data(398 downto 398) & xcvr_native_a10_0_rx_parallel_data(397 downto 397) & xcvr_native_a10_0_rx_parallel_data(396 downto 396) & xcvr_native_a10_0_rx_parallel_data(395 downto 395) & xcvr_native_a10_0_rx_parallel_data(394 downto 394) & xcvr_native_a10_0_rx_parallel_data(383 downto 383) & xcvr_native_a10_0_rx_parallel_data(382 downto 382) & xcvr_native_a10_0_rx_parallel_data(381 downto 381) & xcvr_native_a10_0_rx_parallel_data(380 downto 380) & xcvr_native_a10_0_rx_parallel_data(379 downto 379) & xcvr_native_a10_0_rx_parallel_data(378 downto 378) & xcvr_native_a10_0_rx_parallel_data(377 downto 377) & xcvr_native_a10_0_rx_parallel_data(376 downto 376) & xcvr_native_a10_0_rx_parallel_data(375 downto 375) & xcvr_native_a10_0_rx_parallel_data(374 downto 374) & xcvr_native_a10_0_rx_parallel_data(373 downto 373) & xcvr_native_a10_0_rx_parallel_data(372 downto 372) & xcvr_native_a10_0_rx_parallel_data(371 downto 371) & xcvr_native_a10_0_rx_parallel_data(370 downto 370) & xcvr_native_a10_0_rx_parallel_data(369 downto 369) & xcvr_native_a10_0_rx_parallel_data(368 downto 368) & xcvr_native_a10_0_rx_parallel_data(367 downto 367) & xcvr_native_a10_0_rx_parallel_data(366 downto 366) & xcvr_native_a10_0_rx_parallel_data(365 downto 365) & xcvr_native_a10_0_rx_parallel_data(364 downto 364) & xcvr_native_a10_0_rx_parallel_data(363 downto 363) & xcvr_native_a10_0_rx_parallel_data(362 downto 362) & xcvr_native_a10_0_rx_parallel_data(361 downto 361) & xcvr_native_a10_0_rx_parallel_data(360 downto 360) & xcvr_native_a10_0_rx_parallel_data(359 downto 359) & xcvr_native_a10_0_rx_parallel_data(358 downto 358) & xcvr_native_a10_0_rx_parallel_data(357 downto 357) & xcvr_native_a10_0_rx_parallel_data(356 downto 356) & xcvr_native_a10_0_rx_parallel_data(355 downto 355) & xcvr_native_a10_0_rx_parallel_data(354 downto 354) & xcvr_native_a10_0_rx_parallel_data(353 downto 353) & xcvr_native_a10_0_rx_parallel_data(352 downto 352) & xcvr_native_a10_0_rx_parallel_data(351 downto 351) & xcvr_native_a10_0_rx_parallel_data(350 downto 350) & xcvr_native_a10_0_rx_parallel_data(349 downto 349) & xcvr_native_a10_0_rx_parallel_data(348 downto 348) & xcvr_native_a10_0_rx_parallel_data(347 downto 347) & xcvr_native_a10_0_rx_parallel_data(346 downto 346) & xcvr_native_a10_0_rx_parallel_data(345 downto 345) & xcvr_native_a10_0_rx_parallel_data(344 downto 344) & xcvr_native_a10_0_rx_parallel_data(343 downto 343) & xcvr_native_a10_0_rx_parallel_data(342 downto 342) & xcvr_native_a10_0_rx_parallel_data(341 downto 341) & xcvr_native_a10_0_rx_parallel_data(340 downto 340) & xcvr_native_a10_0_rx_parallel_data(339 downto 339) & xcvr_native_a10_0_rx_parallel_data(338 downto 338) & xcvr_native_a10_0_rx_parallel_data(337 downto 337) & xcvr_native_a10_0_rx_parallel_data(336 downto 336) & xcvr_native_a10_0_rx_parallel_data(335 downto 335) & xcvr_native_a10_0_rx_parallel_data(334 downto 334) & xcvr_native_a10_0_rx_parallel_data(333 downto 333) & xcvr_native_a10_0_rx_parallel_data(332 downto 332) & xcvr_native_a10_0_rx_parallel_data(331 downto 331) & xcvr_native_a10_0_rx_parallel_data(330 downto 330) & xcvr_native_a10_0_rx_parallel_data(329 downto 329) & xcvr_native_a10_0_rx_parallel_data(328 downto 328) & xcvr_native_a10_0_rx_parallel_data(327 downto 327) & xcvr_native_a10_0_rx_parallel_data(326 downto 326) & xcvr_native_a10_0_rx_parallel_data(325 downto 325) & xcvr_native_a10_0_rx_parallel_data(324 downto 324) & xcvr_native_a10_0_rx_parallel_data(323 downto 323) & xcvr_native_a10_0_rx_parallel_data(322 downto 322) & xcvr_native_a10_0_rx_parallel_data(321 downto 321) & xcvr_native_a10_0_rx_parallel_data(320 downto 320) & xcvr_native_a10_0_rx_parallel_data(319 downto 319) & xcvr_native_a10_0_rx_parallel_data(318 downto 318) & xcvr_native_a10_0_rx_parallel_data(317 downto 317) & xcvr_native_a10_0_rx_parallel_data(316 downto 316) & xcvr_native_a10_0_rx_parallel_data(315 downto 315) & xcvr_native_a10_0_rx_parallel_data(314 downto 314) & xcvr_native_a10_0_rx_parallel_data(313 downto 313) & xcvr_native_a10_0_rx_parallel_data(312 downto 312) & xcvr_native_a10_0_rx_parallel_data(311 downto 311) & xcvr_native_a10_0_rx_parallel_data(310 downto 310) & xcvr_native_a10_0_rx_parallel_data(309 downto 309) & xcvr_native_a10_0_rx_parallel_data(308 downto 308) & xcvr_native_a10_0_rx_parallel_data(307 downto 307) & xcvr_native_a10_0_rx_parallel_data(306 downto 306) & xcvr_native_a10_0_rx_parallel_data(305 downto 305) & xcvr_native_a10_0_rx_parallel_data(304 downto 304) & xcvr_native_a10_0_rx_parallel_data(303 downto 303) & xcvr_native_a10_0_rx_parallel_data(302 downto 302) & xcvr_native_a10_0_rx_parallel_data(301 downto 301) & xcvr_native_a10_0_rx_parallel_data(300 downto 300) & xcvr_native_a10_0_rx_parallel_data(299 downto 299) & xcvr_native_a10_0_rx_parallel_data(298 downto 298) & xcvr_native_a10_0_rx_parallel_data(297 downto 297) & xcvr_native_a10_0_rx_parallel_data(296 downto 296) & xcvr_native_a10_0_rx_parallel_data(295 downto 295) & xcvr_native_a10_0_rx_parallel_data(294 downto 294) & xcvr_native_a10_0_rx_parallel_data(293 downto 293) & xcvr_native_a10_0_rx_parallel_data(292 downto 292) & xcvr_native_a10_0_rx_parallel_data(291 downto 291) & xcvr_native_a10_0_rx_parallel_data(290 downto 290) & xcvr_native_a10_0_rx_parallel_data(289 downto 289) & xcvr_native_a10_0_rx_parallel_data(288 downto 288) & xcvr_native_a10_0_rx_parallel_data(287 downto 287) & xcvr_native_a10_0_rx_parallel_data(286 downto 286) & xcvr_native_a10_0_rx_parallel_data(285 downto 285) & xcvr_native_a10_0_rx_parallel_data(284 downto 284) & xcvr_native_a10_0_rx_parallel_data(283 downto 283) & xcvr_native_a10_0_rx_parallel_data(282 downto 282) & xcvr_native_a10_0_rx_parallel_data(271 downto 271) & xcvr_native_a10_0_rx_parallel_data(270 downto 270) & xcvr_native_a10_0_rx_parallel_data(269 downto 269) & xcvr_native_a10_0_rx_parallel_data(268 downto 268) & xcvr_native_a10_0_rx_parallel_data(267 downto 267) & xcvr_native_a10_0_rx_parallel_data(266 downto 266) & xcvr_native_a10_0_rx_parallel_data(255 downto 255) & xcvr_native_a10_0_rx_parallel_data(254 downto 254) & xcvr_native_a10_0_rx_parallel_data(253 downto 253) & xcvr_native_a10_0_rx_parallel_data(252 downto 252) & xcvr_native_a10_0_rx_parallel_data(251 downto 251) & xcvr_native_a10_0_rx_parallel_data(250 downto 250) & xcvr_native_a10_0_rx_parallel_data(249 downto 249) & xcvr_native_a10_0_rx_parallel_data(248 downto 248) & xcvr_native_a10_0_rx_parallel_data(247 downto 247) & xcvr_native_a10_0_rx_parallel_data(246 downto 246) & xcvr_native_a10_0_rx_parallel_data(245 downto 245) & xcvr_native_a10_0_rx_parallel_data(244 downto 244) & xcvr_native_a10_0_rx_parallel_data(243 downto 243) & xcvr_native_a10_0_rx_parallel_data(242 downto 242) & xcvr_native_a10_0_rx_parallel_data(241 downto 241) & xcvr_native_a10_0_rx_parallel_data(240 downto 240) & xcvr_native_a10_0_rx_parallel_data(239 downto 239) & xcvr_native_a10_0_rx_parallel_data(238 downto 238) & xcvr_native_a10_0_rx_parallel_data(237 downto 237) & xcvr_native_a10_0_rx_parallel_data(236 downto 236) & xcvr_native_a10_0_rx_parallel_data(235 downto 235) & xcvr_native_a10_0_rx_parallel_data(234 downto 234) & xcvr_native_a10_0_rx_parallel_data(233 downto 233) & xcvr_native_a10_0_rx_parallel_data(232 downto 232) & xcvr_native_a10_0_rx_parallel_data(231 downto 231) & xcvr_native_a10_0_rx_parallel_data(230 downto 230) & xcvr_native_a10_0_rx_parallel_data(229 downto 229) & xcvr_native_a10_0_rx_parallel_data(228 downto 228) & xcvr_native_a10_0_rx_parallel_data(227 downto 227) & xcvr_native_a10_0_rx_parallel_data(226 downto 226) & xcvr_native_a10_0_rx_parallel_data(225 downto 225) & xcvr_native_a10_0_rx_parallel_data(224 downto 224) & xcvr_native_a10_0_rx_parallel_data(223 downto 223) & xcvr_native_a10_0_rx_parallel_data(222 downto 222) & xcvr_native_a10_0_rx_parallel_data(221 downto 221) & xcvr_native_a10_0_rx_parallel_data(220 downto 220) & xcvr_native_a10_0_rx_parallel_data(219 downto 219) & xcvr_native_a10_0_rx_parallel_data(218 downto 218) & xcvr_native_a10_0_rx_parallel_data(217 downto 217) & xcvr_native_a10_0_rx_parallel_data(216 downto 216) & xcvr_native_a10_0_rx_parallel_data(215 downto 215) & xcvr_native_a10_0_rx_parallel_data(214 downto 214) & xcvr_native_a10_0_rx_parallel_data(213 downto 213) & xcvr_native_a10_0_rx_parallel_data(212 downto 212) & xcvr_native_a10_0_rx_parallel_data(211 downto 211) & xcvr_native_a10_0_rx_parallel_data(210 downto 210) & xcvr_native_a10_0_rx_parallel_data(209 downto 209) & xcvr_native_a10_0_rx_parallel_data(208 downto 208) & xcvr_native_a10_0_rx_parallel_data(207 downto 207) & xcvr_native_a10_0_rx_parallel_data(206 downto 206) & xcvr_native_a10_0_rx_parallel_data(205 downto 205) & xcvr_native_a10_0_rx_parallel_data(204 downto 204) & xcvr_native_a10_0_rx_parallel_data(203 downto 203) & xcvr_native_a10_0_rx_parallel_data(202 downto 202) & xcvr_native_a10_0_rx_parallel_data(201 downto 201) & xcvr_native_a10_0_rx_parallel_data(200 downto 200) & xcvr_native_a10_0_rx_parallel_data(199 downto 199) & xcvr_native_a10_0_rx_parallel_data(198 downto 198) & xcvr_native_a10_0_rx_parallel_data(197 downto 197) & xcvr_native_a10_0_rx_parallel_data(196 downto 196) & xcvr_native_a10_0_rx_parallel_data(195 downto 195) & xcvr_native_a10_0_rx_parallel_data(194 downto 194) & xcvr_native_a10_0_rx_parallel_data(193 downto 193) & xcvr_native_a10_0_rx_parallel_data(192 downto 192) & xcvr_native_a10_0_rx_parallel_data(191 downto 191) & xcvr_native_a10_0_rx_parallel_data(190 downto 190) & xcvr_native_a10_0_rx_parallel_data(189 downto 189) & xcvr_native_a10_0_rx_parallel_data(188 downto 188) & xcvr_native_a10_0_rx_parallel_data(187 downto 187) & xcvr_native_a10_0_rx_parallel_data(186 downto 186) & xcvr_native_a10_0_rx_parallel_data(185 downto 185) & xcvr_native_a10_0_rx_parallel_data(184 downto 184) & xcvr_native_a10_0_rx_parallel_data(183 downto 183) & xcvr_native_a10_0_rx_parallel_data(182 downto 182) & xcvr_native_a10_0_rx_parallel_data(181 downto 181) & xcvr_native_a10_0_rx_parallel_data(180 downto 180) & xcvr_native_a10_0_rx_parallel_data(179 downto 179) & xcvr_native_a10_0_rx_parallel_data(178 downto 178) & xcvr_native_a10_0_rx_parallel_data(177 downto 177) & xcvr_native_a10_0_rx_parallel_data(176 downto 176) & xcvr_native_a10_0_rx_parallel_data(175 downto 175) & xcvr_native_a10_0_rx_parallel_data(174 downto 174) & xcvr_native_a10_0_rx_parallel_data(173 downto 173) & xcvr_native_a10_0_rx_parallel_data(172 downto 172) & xcvr_native_a10_0_rx_parallel_data(171 downto 171) & xcvr_native_a10_0_rx_parallel_data(170 downto 170) & xcvr_native_a10_0_rx_parallel_data(169 downto 169) & xcvr_native_a10_0_rx_parallel_data(168 downto 168) & xcvr_native_a10_0_rx_parallel_data(167 downto 167) & xcvr_native_a10_0_rx_parallel_data(166 downto 166) & xcvr_native_a10_0_rx_parallel_data(165 downto 165) & xcvr_native_a10_0_rx_parallel_data(164 downto 164) & xcvr_native_a10_0_rx_parallel_data(163 downto 163) & xcvr_native_a10_0_rx_parallel_data(162 downto 162) & xcvr_native_a10_0_rx_parallel_data(161 downto 161) & xcvr_native_a10_0_rx_parallel_data(160 downto 160) & xcvr_native_a10_0_rx_parallel_data(159 downto 159) & xcvr_native_a10_0_rx_parallel_data(158 downto 158) & xcvr_native_a10_0_rx_parallel_data(157 downto 157) & xcvr_native_a10_0_rx_parallel_data(156 downto 156) & xcvr_native_a10_0_rx_parallel_data(155 downto 155) & xcvr_native_a10_0_rx_parallel_data(154 downto 154) & xcvr_native_a10_0_rx_parallel_data(143 downto 143) & xcvr_native_a10_0_rx_parallel_data(142 downto 142) & xcvr_native_a10_0_rx_parallel_data(141 downto 141) & xcvr_native_a10_0_rx_parallel_data(140 downto 140) & xcvr_native_a10_0_rx_parallel_data(139 downto 139) & xcvr_native_a10_0_rx_parallel_data(138 downto 138) & xcvr_native_a10_0_rx_parallel_data(127 downto 127) & xcvr_native_a10_0_rx_parallel_data(126 downto 126) & xcvr_native_a10_0_rx_parallel_data(125 downto 125) & xcvr_native_a10_0_rx_parallel_data(124 downto 124) & xcvr_native_a10_0_rx_parallel_data(123 downto 123) & xcvr_native_a10_0_rx_parallel_data(122 downto 122) & xcvr_native_a10_0_rx_parallel_data(121 downto 121) & xcvr_native_a10_0_rx_parallel_data(120 downto 120) & xcvr_native_a10_0_rx_parallel_data(119 downto 119) & xcvr_native_a10_0_rx_parallel_data(118 downto 118) & xcvr_native_a10_0_rx_parallel_data(117 downto 117) & xcvr_native_a10_0_rx_parallel_data(116 downto 116) & xcvr_native_a10_0_rx_parallel_data(115 downto 115) & xcvr_native_a10_0_rx_parallel_data(114 downto 114) & xcvr_native_a10_0_rx_parallel_data(113 downto 113) & xcvr_native_a10_0_rx_parallel_data(112 downto 112) & xcvr_native_a10_0_rx_parallel_data(111 downto 111) & xcvr_native_a10_0_rx_parallel_data(110 downto 110) & xcvr_native_a10_0_rx_parallel_data(109 downto 109) & xcvr_native_a10_0_rx_parallel_data(108 downto 108) & xcvr_native_a10_0_rx_parallel_data(107 downto 107) & xcvr_native_a10_0_rx_parallel_data(106 downto 106) & xcvr_native_a10_0_rx_parallel_data(105 downto 105) & xcvr_native_a10_0_rx_parallel_data(104 downto 104) & xcvr_native_a10_0_rx_parallel_data(103 downto 103) & xcvr_native_a10_0_rx_parallel_data(102 downto 102) & xcvr_native_a10_0_rx_parallel_data(101 downto 101) & xcvr_native_a10_0_rx_parallel_data(100 downto 100) & xcvr_native_a10_0_rx_parallel_data(99 downto 99) & xcvr_native_a10_0_rx_parallel_data(98 downto 98) & xcvr_native_a10_0_rx_parallel_data(97 downto 97) & xcvr_native_a10_0_rx_parallel_data(96 downto 96) & xcvr_native_a10_0_rx_parallel_data(95 downto 95) & xcvr_native_a10_0_rx_parallel_data(94 downto 94) & xcvr_native_a10_0_rx_parallel_data(93 downto 93) & xcvr_native_a10_0_rx_parallel_data(92 downto 92) & xcvr_native_a10_0_rx_parallel_data(91 downto 91) & xcvr_native_a10_0_rx_parallel_data(90 downto 90) & xcvr_native_a10_0_rx_parallel_data(89 downto 89) & xcvr_native_a10_0_rx_parallel_data(88 downto 88) & xcvr_native_a10_0_rx_parallel_data(87 downto 87) & xcvr_native_a10_0_rx_parallel_data(86 downto 86) & xcvr_native_a10_0_rx_parallel_data(85 downto 85) & xcvr_native_a10_0_rx_parallel_data(84 downto 84) & xcvr_native_a10_0_rx_parallel_data(83 downto 83) & xcvr_native_a10_0_rx_parallel_data(82 downto 82) & xcvr_native_a10_0_rx_parallel_data(81 downto 81) & xcvr_native_a10_0_rx_parallel_data(80 downto 80) & xcvr_native_a10_0_rx_parallel_data(79 downto 79) & xcvr_native_a10_0_rx_parallel_data(78 downto 78) & xcvr_native_a10_0_rx_parallel_data(77 downto 77) & xcvr_native_a10_0_rx_parallel_data(76 downto 76) & xcvr_native_a10_0_rx_parallel_data(75 downto 75) & xcvr_native_a10_0_rx_parallel_data(74 downto 74) & xcvr_native_a10_0_rx_parallel_data(73 downto 73) & xcvr_native_a10_0_rx_parallel_data(72 downto 72) & xcvr_native_a10_0_rx_parallel_data(71 downto 71) & xcvr_native_a10_0_rx_parallel_data(70 downto 70) & xcvr_native_a10_0_rx_parallel_data(69 downto 69) & xcvr_native_a10_0_rx_parallel_data(68 downto 68) & xcvr_native_a10_0_rx_parallel_data(67 downto 67) & xcvr_native_a10_0_rx_parallel_data(66 downto 66) & xcvr_native_a10_0_rx_parallel_data(65 downto 65) & xcvr_native_a10_0_rx_parallel_data(64 downto 64) & xcvr_native_a10_0_rx_parallel_data(63 downto 63) & xcvr_native_a10_0_rx_parallel_data(62 downto 62) & xcvr_native_a10_0_rx_parallel_data(61 downto 61) & xcvr_native_a10_0_rx_parallel_data(60 downto 60) & xcvr_native_a10_0_rx_parallel_data(59 downto 59) & xcvr_native_a10_0_rx_parallel_data(58 downto 58) & xcvr_native_a10_0_rx_parallel_data(57 downto 57) & xcvr_native_a10_0_rx_parallel_data(56 downto 56) & xcvr_native_a10_0_rx_parallel_data(55 downto 55) & xcvr_native_a10_0_rx_parallel_data(54 downto 54) & xcvr_native_a10_0_rx_parallel_data(53 downto 53) & xcvr_native_a10_0_rx_parallel_data(52 downto 52) & xcvr_native_a10_0_rx_parallel_data(51 downto 51) & xcvr_native_a10_0_rx_parallel_data(50 downto 50) & xcvr_native_a10_0_rx_parallel_data(49 downto 49) & xcvr_native_a10_0_rx_parallel_data(48 downto 48) & xcvr_native_a10_0_rx_parallel_data(47 downto 47) & xcvr_native_a10_0_rx_parallel_data(46 downto 46) & xcvr_native_a10_0_rx_parallel_data(45 downto 45) & xcvr_native_a10_0_rx_parallel_data(44 downto 44) & xcvr_native_a10_0_rx_parallel_data(43 downto 43) & xcvr_native_a10_0_rx_parallel_data(42 downto 42) & xcvr_native_a10_0_rx_parallel_data(41 downto 41) & xcvr_native_a10_0_rx_parallel_data(40 downto 40) & xcvr_native_a10_0_rx_parallel_data(39 downto 39) & xcvr_native_a10_0_rx_parallel_data(38 downto 38) & xcvr_native_a10_0_rx_parallel_data(37 downto 37) & xcvr_native_a10_0_rx_parallel_data(36 downto 36) & xcvr_native_a10_0_rx_parallel_data(35 downto 35) & xcvr_native_a10_0_rx_parallel_data(34 downto 34) & xcvr_native_a10_0_rx_parallel_data(33 downto 33) & xcvr_native_a10_0_rx_parallel_data(32 downto 32) & xcvr_native_a10_0_rx_parallel_data(31 downto 31) & xcvr_native_a10_0_rx_parallel_data(30 downto 30) & xcvr_native_a10_0_rx_parallel_data(29 downto 29) & xcvr_native_a10_0_rx_parallel_data(28 downto 28) & xcvr_native_a10_0_rx_parallel_data(27 downto 27) & xcvr_native_a10_0_rx_parallel_data(26 downto 26) & xcvr_native_a10_0_rx_parallel_data(15 downto 15) & xcvr_native_a10_0_rx_parallel_data(14 downto 14) & xcvr_native_a10_0_rx_parallel_data(13 downto 13) & xcvr_native_a10_0_rx_parallel_data(12 downto 12) & xcvr_native_a10_0_rx_parallel_data(11 downto 11) & xcvr_native_a10_0_rx_parallel_data(10 downto 10);

end architecture rtl; -- of gx_std_x6
