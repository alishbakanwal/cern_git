// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:24 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bh6jTFBbhh8xI2/SybHJI9zKMJncKkde+B9IoZfRufaoHLVdknRWFrKPouSjdmHf
gkFyUG1ymKIN45ocWnuBbDN2qcyWJhfJpQbts+Xb0Vi+HdVqnnvq9bZn13zRsyct
8oGY3SE/MFNM0t2Q5/M2YYchiN+6Dh4lvcbjKtdP3/c=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3072)
xQ8eC+9KK/3+gCgbbTIY7yk3SrEoTmHwiFETf5H5BM6J590dfn0EOZOxD2s+JiLt
o7LYoIAemcqGNB5N0krdiqEHY/2eoYaCRKH/h62Qb5widkGV72W9SWFT7+BjkaPM
DhhVM7SewRcuCsP1Z+jj7NSfFyzed8xRG5Hn+O0EEd1XafMtb53hQ7fWLdsbOH5E
3tNbLp8709nPgj9zWx08DAVdYX6Ycwd8Mty9BWEICQlqE38T9yYokahP3lc8V8VH
cBxXksE6+GqXFD3FXfUfaAr0GKUw1iMuERSWZK2muNjGsCOXm/hNvRJls16ptsoq
/lsnutmA5NMj0qD/5OTeP31ghHGGRO0NLGGznWttW9hr9QbDgranJrIM6AVSnNU4
y/TlLOgFdl8BnxrHdD7yMKbkal9BeHatroQ/Btmbvy+YEmgIog3aii7/WvVKmAR+
GVZvhUFAQIk/Gt4Fxczw4Rwlgu9J5EwH8k5VSjfylVUfVXcSAYuAPwdSQHdytKQ9
GwoMRem3hy9mB6mDUS3ifhTwxRjzwk9NFpFcaFrNCrwhiR7MrUCcf+/eY+P8wSSu
dLQEypkYw8gjJjO3Hgt8Ex7pbE83hkYEKRbzrJ+udzHquGVmGJxnQNR2+5nUvOSm
F6EsGW1iMUys1cj5vButY9hUZ41aYbq7QKM0acP2WOkFY4exTLLvkRs8xN2WJo8c
/cK1oUEbBuNttLLAWeBaZCTHfW1XvG6gEiWXUizCiStILSLrOViSjgjQLeKxuqsL
N/XoYEZV9RaWoNq9gMTBgc2fLSq16rkuOOSkewSneXpp7ZTx6DcncPCicQ/nq7X8
mAW+0mpgq8BZ4ZPy8FH/KeLuFetqnJAKOtwlTJOgioeGlYlJo2q7Z+1usJhkJ5xt
orliOwMHYaEmbv7x5e0+BNbgsdztjHcJ5b8+krFTe3WeYo7Xc0un3AEToYxw71jc
UCVLDpTc3QEm7GrIrjSz2Gtd81/IE8Uum4qYxv9+58ZwoQ7DyI2pJBTTfim52qh+
XcMiyRxAp1DQny9CkfoXmbN4wDzW/lce2+cq9bblAoSGkNvYLyKVV5RJxaBeJ7UL
bbb7CrffYzMtHlJU6cweMnMO+LlzBCMc7hrmXfnwzaIqTFAuKgT3P+hlytRSnApB
j7SeT0O+L9Q/Yzlo7SNxeGZOHWgXk5z6+m0XBkClbRgZh481Z0kM8h9PaAZjCS2g
Hb/zYZ1HJm0o/Pp0CHkdJZzHh2uheglO1v52nzufS8vpsyEtDuJU1ZoBfXBS6olq
PqOBQZ0uyDEprKbhFrwseutn18Z8FQrH1P5kY9dxETIWKpWhepX0Nuk0Jm4u3QAI
ttC9rNhnPSilYqPnLxEUDHC4LrRBB2WSMeYGctZzmvg4riFMU/9BqHcRV5XjsV/5
s6LEIDvSCpFXobffPFl5eap8zIiiHJtKtHwHDMWQPOEfjxepsfopQ2huwlGatQ8t
ZNAYPhG/nq5zCoIDjz4qAo0w/ZX8rx9/t+sY9gvL0bxUQyWE46pVQZd5V/UbF1U8
mLXXdxmb04ASOK1UaFZtqySBOLCe7VuYj6/roxtht0tDCcW0GgNpl4XzgKiBMre9
ROFvcMeUwbgRRbS3RgLeui5HmVyLx9olnzdX0J5cJ6Y0v/WJHI51UKldM6U9dM4L
rBESd+434AjloEqwkR6BnLLBfVvRKYz82dzlksf+1NvJAN7KU8MdRORFoHodDlXI
hv+HGUz309KGCMZ3vRl0YQdnM+mkKxG1LnNm5Gmxeq4EoXQkp+OLPph8nll6h5UV
qyOBgeMxz60INmwS//p18NkukEPbxZ77qvmU4zjZuJNjdnWNscm2LYZFKUDE1yxx
etG50HzLVsYBm/FbyfS1UOjdbO92ijlSRcCa5KwlZaBQf3ADjEsUWfRuFrU6mssG
XTuuUQdElItJ4JdaemthBljk2VBq8IdZ/cQi/lXDWWTeSBUNHrgqiizgUfaLR/SP
YLjRvlpYvgZ+5VrNqRHqfoWiVHtEiznA+yGdF4qpFqC6L9r0hmkFaIlreiO3tlA7
c58ZRyKaG5RiDiQFBomB8IbMh6y9Tyi1FbPO5T0wHLGV6Xv3yjtUhM0NNxJYwVIs
/LrVQLhXJOw1Qbh2q5ZAF0WeppXj/ya/cMGg4A+a6U3u9aATIpDnl5OJvRKe4LYB
t/xnWUC+YlbZjTb8XARpJnjlf7kbH5a8k5CvgjSXL+tP35a8GmPI8AiPTStZbIae
zz9bxRvXiXKpNz7KS3CIGLipf31R4nDLPWOsTwmXDyXud+DkTmWs/dKp481671hV
Op6FyqKujrgBJqqjCjip53z35KScSszCyNZbQubvX76nneAGdFFxBRCEYOrU7WPA
XR7DfjmeKKZpcTtaskplkaKKYzBznWV4Kgi5yDqGjWRLU3wWWGK471jtj6qE40Gj
LQhF3ECbDCGBvaybJTwz7Qa9CYR2krVhDWXhSDq2zquUG37Q5BQZVsUtaQaBJ7Fc
NkgfPo7F/Cs55qZmBny03mzEZ7uWWgIk++JV4sbYMCmiwlNVPeslu4YB9Mla8jv6
6ZXomrBYaDDwf54Q82Da2Yi/FVQPVkhj1GIAPnQ1ZQvQlwte0h+OlWnS99Y8p9nS
yF5t61uTps/hIXW1UyriOiOtnfrnGOen0g03BYEfnbLAIrf08Bze/SeoRwn4E/F+
JPPIaNiGMOBfeU9diatQZYXGkx+Nrx5bteL47EpaVTC1Mxz55Qxfe+o0iZyWq4Xg
DcjCTrJb+wmWlrTBkztRz6QEUsrfVAspHE5YlLtGhCIemU6augfpPKU5jOiJG/LH
Fp5hDaj4bY0kp10QFj1lgRduHzwNrW7EzmKRoUgMDe/tAUM/g2muBjDDvnE5AjCu
+ui/SmqzLphaq83KW3ZyKqdOgMvLN3Kwk056/22hDca73VZDbtprBL65EqO/gpxk
BSSF94HKeo8KeKwZ4VGpa2GguUCmvh0vMMzolQGIa7t6btvjTAAeeZhTmA/tyW3e
GV7UUTuF28ymQQFcJPYuMqOH/FhzxhDBIGB/2Q6OENAxOmjaBffMfWm2SYIih6RG
+q5vsUBJmhOOQa/LMMDB8C5e/uGCMwzxd4eN4Hqw04ZJ2KZofZULE3CJl9PHrOQs
YT9/Z0c1uTWia2D8NoiEwdgrcLdPon3nM8oCpM7iG+unsyO1zt0b5RKz+lFMcaFM
2TSQ1s4OVSHLZT+lvosNKzQxxRtMxurQYte+HFF51QI4FJjENCh7B1+w4cf1U5vV
ma38tyW4UMVg2OGUXn7erOrzurRjaYSSzdLL6uHLoJExGElpnpJQ7hzuYhBDNtaD
7SC4C11kxOvHzh6ZHkPjDQ4z2tPLbsaccZD0Qfnm501DF32EI2vwUwBPVX80hs3n
AXwA46oS2s/lrHMQSiwDwKurfRtCLlPjZ5fF4/bhQt4h3pKcOu5WZPLnZL6UW8jv
eeD9WLWswr8bYPseGgBKqDLW/aodXokqzUr/yM0p38a77sr4im7LQuwyWLjrAn64
/iS8z+LbmpzcTO5m1Nq/kyhqSOqSFYX/xTfvM4dlEPcdqoZdWBzJI5gv+Y1nOdpk
iTJVwygrC1eee0mo3xh/Hi3qSf6xvleJiQWb+T2lRqpfk+en4Ym8VIxxNX2YRdSQ
7E8oVyvXpQN05g1Ssc26njdIypkjdnzYhdiQJ1BWnrI07A1w2oXV7eDiCDFhyeav
+uHPL8H+hBIQKnklrD9+39WHyZB0FEmyzCKyvA+slPGZADt6DCwvrnMIHeWNpiw3
2T0nfuQjPDfzXk8rTCAYL4If3LXBC+kZVmuPJlgu8guBUqtRERyzuOAiuzRshxQo
m+xVxyuV7MhHoNwAhXVLNv7NcUmhqQMsZyBtqUVThdn4jS9R5YrwJEqsK+Q8DH0p
Gd1MFJMMVgVFN5g7E+p8+Ee2bdrZ+DBC2oyxjY0wb7GGrJTm+NmyoLiVVZRHSLNd
WrslYqG7OF2oST9PSPNqp2FmfSOceakdQ1quKIDMs7oonWlpO4lyAwdm35r46q0S
PkGPwYI0/QTgmEoHaxsJFHa3TTqmvy2kPfDJ8bybMkjQIodKLULJXMI+bY0WOpCl
`pragma protect end_protected
