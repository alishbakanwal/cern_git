// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:16 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oJfYYinosP3ECIu+pl58hIn2FtTFvtVdLbPs6hrQ0zO10hsC0R9fOfhFeQp/QQa6
ocfjcW5aAUczHgD/834i2SeSuwKbjhGr0/S5q/dGjc0mBEZJ+ZQgGUlH4/vd7JU9
rqxcO7ujokaZIbgdmvVZxAODQtN2c9VKE/RkbX4bjBs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17968)
8JFGkE6HKpqnB8v5B3HlsTOdoqeAo/m5hfyGR/pKNjn8gq8zlVP3j9ZC12FmXvsa
aoHTbiDQ2EMvREeHS2hdNxnzjyIoDf6LhlGRcARJ8UXec90KFSz05frsukYRJqDn
LxWxe8orBoMGTBu7t2Tni4OfvgQHkh9MHQ2xklWq8KsqiJkAWD3SlkGcBfbn3NAI
hUkIFN8Kf3VF3v9dznbrY54L0pgLDyMAGwzrQYEP6+5TN+NHC5qfY8emCMSVlom3
jTz5gwPl8DgdcZaecaGu9ov6XyeQbNTMMP1MOFelnOwWtxrlSzpj+wUnSHiosy0i
H/alVUaZGE+LUz6elxTT+kOLj0yH8UEpqeuonf9of7iDfI2U7woUza7/cZsGInML
JXWHRoWumniQucTIdID2DxthfU+b+QQY58TqmEyVn1xMUDBft0ZaTXDnlOlr6Q/X
YqzoRF4PIYkk56BD9GL9G4q9RWaP8ARUrHLXrAiEN/Tbl4UKMPxR00y5eEx10jZF
u6tGvzbvhzSK6iDYz/LKXW9V2JoRoRzH5j/9GhO16gPY6bK+hQFZJ276JpkeDUD5
9O6s06h0OOh5y4I1vIW6b9ECKoeQVdThMCqsGfAFVLV+GDFfPk3u2B/J+2loe6uq
yFJeKIfn6XK8eL7yFrd5VzB46eqR6WdrB31wu0L3VkoGMWsjgJKETVhp67m4TA4s
L0NXtq8LFWJ/hJVmGcpnHhB/0Ox/ZXuo7FwR6o5S8IwINIfonFPaZT/rwQjpG74x
uvYyvpxyVF7SwhGAm7hVPskGsrnkCLNEeRQ0OZVFMYqnbOKcVX/1nbTOhq+6Dg7l
kYqQZ97bkHpKuee2fwGBCFC3MacBAp15Xiq1AJD+c5V0eRzDJpGCuS8BayoVACdn
OWxTfjuOHI/xWfN/Z63iDy5q3fa9LI4GNDYUza8YywuGxT+HOGTF7TLKskomfCQh
wJgaT4XkcFOMRBTllbCE51LCQOgeu4c0g3NDP5UtLFojfrsioBuu//SAJ17q85vI
t3/IAwFCUetUssyY/MWIOhK2ATVd0u/J8FbjqDZ0JdZo60AcL+QNaAUNyED5J5YG
dHObxwvLokMfP+k52oGqDJdwtpbjpjcvxNS3T3DrzaYuri/+ROnJYSZr0a2hw1vE
cNVKAkHKsqWdeuw8+02fD1oRl5t+wEb/GTXxfV8btouApW1r5FVFSVYm0MfGqd1l
dSFV4pun8RBSB9xVPWSU45nk544M4Kxk6SWFsyOGpC4rSQYbYdRbul3fc633zWX3
CM3QpD2rBzoSOzu3BLBDRrXR7dQWLEyhDVKfH4bQ2UwXkKm9r+yWh9SGscV2d8NS
9MO5ZWoSD8mXF8lcxzK8zAiaVUUIL0TlPDKHxc9p+1dGspxo0ibUI6HL1en55pau
pWDPnHVKfI/hmbdFaN1ThSWy11llHn6coch9SXFsooe5PJBLNLCModnWLOoA+aIN
47pqc59ZDhjpLBUeJKbNRxWpl4Ot1cLMh2xNpXaJEna4xuqhJ5v//u42UFxUc2D/
Jpx9UfhGPbCOjJq24JIXpLJ0ooM37mei+CS8HVIGJEGk4fd2XOAE7RiJ71MMpuGZ
+RuhWrg7r2ouE/vl5Nk1NMSsRNp31bTpdF6FzCp1A1p6Kh6CcUB0qzhuItfD1/Wl
HF+ZClypcCP1rICZm9hFz0JjSqSCkIp7w8QlOH1KCY4xnLQZI+psSzXqc2SNX1Pl
mtqEAK0tjU6dZGjuvYncwG1mBTTXDvRqevGBWH6oDplYEVFjJvC55/MxhR/am3JM
fkcHHDhQp7kudviHU5PHpV+3dW4+5QRp3j7T7IXfzlzNP2Hv1+Gnv5K237NoahWn
KEEKf8JmiXdb3KktkD/eMGWC/gHadbKqucSh6HWp0QDqU5Oq+aVwd5AtJV3U2bzL
UGlkb/CA2SyLWhKlPGXr5Bhhaewb3PYj7RrWFM95tQsGggwplxCA+uNA5QuHuv+6
RVRHQ2WJeZ5F7i48hHW0PwtfNZLzaaqiHqzKolhgeuNzZwpWlL3iUFVjsxZLdrGb
w+/XwsjLiaQj//0ndZCxN7vfmDd6/AJLBEgolsWlvJna9ibQ4syXE3F1zG0WLudW
Kl7tSNaeVay32/DWmsLLszN/BFnO+UpNYsRCkCOpeQopyfbAgXilK215sqsg2QHA
OGmRrptZTCyzAwf4a+W7pLZPSUtXFHJqvhJ7jmuYP1IkQrCAWJ/3u3xL19egVAyJ
7g6w8a+QR1kudv84iuRYWhUSvlMxOy9go9+d16T44HkFFYGPjr0Y6oGYsDoeftNF
sZkGzezw1YYJE13T3ZyuTn6dvFeKNCZ4lfyPfyAKLNO2f6BdcHFjcNP6y+IHtz1l
EnJ8L92Pff7VI9SIeLQcHXyUIFc0uREaEpC9jfXC+8t6JtbZLTlwq7zF5Sozkiy7
D2x7ps1mFhrNY94lCe6x2/6QCu6iPqby2uslEAHsnEbVi6AxjhrX/08JNB/wQ838
S+FkM+vn7SFKTlf54Hq2TzUN9wHiBa6+13JEZx9U7v01nT+Ab10aORAxuYxzPRKb
T9/ekmQi5ZVhBd5HJdqJyQxM6KiqGjfC7ILHFXxDR0tdOdlfM07J2khr44WRW+1R
zyVk9sgSE5AmkAPQGG5SOucmDLZlf510xTmyXDkVuYF6YQm03b26S/4FT3Xv8d55
RSM0ZmoZupVaF2+bpByTCHdnS/bnjLt0d0EK5brImivNsZ1yAU8uGkByNGKmHPyF
uNo8HdiXd9eCV+HOpntatMML7J5kodD5KtLvE+0tLX7VWqS5xze2Wt6fsamV8Dfs
Dy6L1r6Xs9gpAwDdu54Bk8pw9CKS016yJW4WPzl/aFHffjul4IuQ+/ubVquCq/7d
1i1pZZo2H9DgLBxw45E47XWYGmmKYpt4reL28UMRtu6liobrtkSGfnsSQ5VxQSfe
Q7m2XjqaaSZLtv57lUyct7OEG0s+YZnGQPqJnEOtTVZydMyrVbfdboSGTDV+F1ip
1cvrIaDFRngJWjOdAltH4YQ/xky/T2JtL2VdhqmdSBq4RXb2S+98tb/UD13nvJVj
jJ00QkW63kIp3hVSn6cAlQ9v1MYwWkugiLoYFYwEB5eCutBQ2B8q2a+RfiSVQNq8
sdEp3pI2OjhCn2zh//14OJOo47JfN1ZpCaRZlmaAh37sArdrOUmiy2VCChM2ItDq
6r7QQZ8t68ubLdFKlw+P3tUqCC1u0F6O0vIuazFKDRF9PfP/ntiLRw9Z4UvPjDxa
b+ATLAu8II4TSQOLif89uH/LeWp3n/7pCWEN9kQK2R1J511CYpxg0dhiMcTc8HGM
Hb6/vdVDYaA+F+e9kYaDT6+k8u8Uj3kS4R4gxsy+sox4lKTWBUXeNhW7bSCx9Twt
h64BC+dcDEdpeitGY89YxGnaQzJ74US8tF9VSurtDsfzttPLAfw+5FPTftdPLwi5
d+Zj9+jQf5IuxdqODH1V/S6JGto91Nr7shvk+Sysm+H8l4hSiI/c5i2oHKVytPQM
hr/fVstfup96P55IWQBkLomrxJKMrJT9TUJFigeWJtWQmYIGWrjlwex4iaLFUOOh
h6bqxcy6+W3sbR5NRRHDYr3OpXjtUQtKgiS9YcB7eAJ14UHK2+o9+PN1o6xFG3wz
jdsmBKRjd1acjBKb59W3hyT6JOhBLmCJ7qgs2mm4bfOafceNdUaJLjpeKHt7E1r/
jNlxgdFSnSZ3GXEaNjn562+CHQqlITCqRTmtbq/ftVtoeKsX6yquvX2G/6KMjXyV
5WUckCpR27QlGtmNeKwkfB5Nw7YTNh/QoUpPlMP4kT7T6KyEfunJTtNHw2yUyvLY
3CO+j2bC67w4Llji1U7xQiNJrJCyPqqPA11B9FE+BAAY4dzgIXBgv/LIEkOZ55SJ
JBAypBzUES6E+K46eyg8b1d00MResbxLiyTF8+PWEzWDwFwhgM+WneqtPD+bCkOy
6PTuuhpBeWLxL/VbSmuyYvfd6rHK8CsXDGNx+glzOdyWu+znm3T3U9g/3Dk+aknP
GpHNHdklc7hZIBS7nzGrwJJpTi3aalAczLXfi8qq5gQ4twuQyiSIofJd3GbOTYSQ
WbuO5x+T+qdw7ZWtX9RpWrccX69G1L1Ub5xsQkOqTbfkxrJi7+yW7G0qOVVUzlvb
//k09u8/odeq6B5/lmPyp+Js71ZnAznDiXtXbw/r8eekOa0CSB9knmWPdPpUt7l/
o/e8+03xDu4Ya7rFpDy2nEmX/092r+44y3nZm5SMK2IRo0lJnWmwmI97Jh2J9FCf
WpX00J5q27FlJdq93OAXmcaFMlTZ6Y1vxu/XlAH5A6rw+wrRAUNhVkhpqy4u4Gb7
sqH8eVM5+Ndf3tSEo8ZLrPs864rKF4kXln4tFHN3NMgv1IvgJQLeaklOJkp4q2Lk
y7N+xMymf8jTbK0lSEytK4hUeNoxoWosPg26RqQ2MKbytBSNZljZ7I5+7MqSdqBm
6RT+umaDCwsWhbRf1++Cg1+sSWOGeR6YxFtXJo4uB76j0s1YP51UiSZH38l7RarV
aN2QHenCXPyly/zaPieYFaMrTz3L8AXtUAXDZUwJ8TQG5go7qgarhns7JcWhIqKy
wzELMmnouZxeKPc8hiuIkZSVTNBl/HBCoYRL5lhR0dK5oClI+TF5Onq3ZAjSOcYy
g03Dl3ugof/cdHC2rtfVI+ULHsJxKN0G7shI7qEfRYbGVE16mVmNBBsIQXJiqOxD
QmvdXaBkcvFNERG2ZZsSPq3skT8r+wlwlgLUQEpldWOZaul5lkGlmhYtoAU7OclV
vRsj/itO+iTu3naPUD9maFhM5sGFRKR54Wq0gdwahsxtsDi3GrphbzY4LYcc68/Q
ORe3g+ytNcOg6AVcuMWchiQBUSznQfw1IlYsJKglZ/SupOBQAHrTS9aZN8cmHBlH
3WIP9Pu6Iuee2922terUXA38S8ueiLXm+3XThjIUTAWEukorZVDxUP4BybXAVHxY
5h5IrbDGHI6LXg08kReoQGw2bWnhKfZzbMx5Opd5yeuOt/gdG9qOihyMikgKF0bl
y/n8+ivuU5z+1J9gZq5v6uVGRhHapnxrAM8VtnJWO/e9CadoQswAOt9F0EvZYJer
dGf0OZ7vjfsq8WxEK0fdVuvcZlLGHNqhUSNZRsYrgFD5A3gLkXA0xXQNTZzbik21
WXae3sz4SnrY8FSFJo5c52HMeJwDpSN2eDynrslFxHYHT/B/lkt6HO0O59C4ZoqF
l7BZ+V/iQns1uTnpsFKI1jWWktBUyQzEsU+O2VHrlylOo+lc5MR4SCIUg/DbrtOr
IQxkPDrYw9Jz6PysZ7zTpOqCmK4AwUC9gyCkYBQ6byqEdr6Bd3x8VZ9va3I/9k8T
YXZimrtCksjsyCvkXCImjp7Q7u3jnxz/Qd9xt+SERm+Z32vOKzWf90om/4I6Fznj
gLv/TRN1fV1itMuJ8j39MlKR74QDruF9ShXLdRxyelwnk2mPwcNfhGKaAbWzDjLN
zYCbTUnsQCxkNa1H9PfxYBjm5wwKw6aTcJREHYFhJkei+T4EDmYaNuXqBP/+Rjav
KnGAw5Cfg8FAqesEeOelW68k5JYRfzigGfjepzO+8+NR4EErgNJ+NTlRbOZdSmaM
Rr7BJnH7+b5dqltaUba7yszFASukMn4zERvuoXbyoqgFopoo4WmK60oniJ5CPwpS
UorQ5MysGRF9e1+Y55GGuFI4fIh0CkHPyKLxArQHoKQTk6GGdGPjQeBHzifh98RG
kL+fQT4ViorKGPdtrzrgScgOf8HF2+YonpliAe3nqoyo+c+RBKKzjLZo2Wv4Z5ry
ffudrA1W7fql38liHr54UghnQmKbo5mLJfj4MU7eYcmOXqIPciixVz8De03fJeJD
dOpHg6C3urnXacGO9V0sDthF76bVUvtd3ihMHwSSX9P91kPObaQwxvSQsGg1hyqM
vaINh+0HPA4s+H1chOStbhKmUUkxCUBFbdJZQyd+dTB04AtvSQj+GSM/gmqWtqEC
PRtoyyAOm7WtTARp8J1RJQy99Ngtlhwq7KYJ53xWJmjPPPe4XKUL+OlhuAe7uelo
RnTsfQJvmUO7cPchWPuH9xUO9/3BezOEpHDwHFVVEC/BB18wmWBnrEJuJGW2eKrE
M4Ntgbn6eO2HTCNwvEkddY3MR0kj3akHU5uEo6pNId9B3i918WVnxqHO8d0EUHcs
Qoln+abeZk9nIJYRGmx3xQtfjKztJPAC1AEzuyL52ny0626erQyVfq4SjeRjtY7G
5UB6vn06Mm32SnSKOVuSrOVtz5JZ3GHwQUU98qaj8PaVxSZd2IwSjJpvfTtYDpFg
nOMytLQeuHTwSaobXaVxlpL1h9eI7w7Bcrfnq7Q2JT5CxskilnPmWf9uyXLrP29a
3CEto2yh+nR52TxyRDYlQ/Ncqzg0z0EfoDRMO0Mri/X2PjAnOR79gVljwYrbPERE
Tk5P141jXPB4JggSHiByLWJeL2Qqu0cjOIgBz9fsKNPd3Ot+pBRJgc/HvdvY+hu9
DF7YUOglCuPLhdU/m5Z9MWCFUBpTI+smi+Iwcafl2VIdsyUpe3Ce3V9lxTS7PAmo
bSQzgDsiq8fq84ZnnZX0HW3SIav9bVAENqqeLeqkFkxKU8l8IBqA/KsRwcCO6ic3
Uloo+p7ssUMPP8/fDykJTvu7kXFqMqPwctnlrYhB5hbjHC2ZSySNePom5b+7i4s+
Zb9MG2VU3Du1o466bEwI7Y9ThiQ/xhadsoQJev5NzxtWiUU9w3g44ZGaxjw2Q4jw
5WJXGlQsNl7B1JsLigr50W8fbDdti2GujjcBqawXRf8pDo75sELg7EYoeKUT1toN
kKJMbxDufE26tOzcFYBdDr/V4R6ixY1J6mD3gOJcnFWFK/lkPW6wRL57SHE6OhG6
FfIxPluy0+/HMtxVssKbIvhEBLZEXi3/4E0w1gNERmrAhsCR86d4lItRf+dVR9I1
HuFVFXUOSZghJovrmp+DwkANr1GZuBl7pTATY5JC5p5ge+0b3qPRdphBHznRA3X/
nDL1fCl8XgsKo7cruIkDPuAcjxjv5PECkjKOYCfDmlz0GMC8tEpIqWie6Gqn8J0n
XEpExPCmwmWEaTUQADJ/yY0njUo5vZk/5BqN/mOLqznxyliXRrL8vMxOVelOXJEE
4sm26Xz7n5KFNcrsQdsxubzxZlr+nDdMBH5TXfmTZF8TInfgX3Lu6mOrbDINlqqA
H7Db7Dlcsu2IR0xmUjhns29xkhZEAG7SfIx783z6LWeW0s5MmOq1yAFqc7xUcOmT
thNQUB0TDJLibaNfxU1b2HtTJ3aPKf18DDDccz3MyuMNHdw0fPF8CVeRvgZbqV0d
BRpvTS8+eAz+qcsnTDtl/au+t7JUSiVStVXGh3uRMDHk71JKGuxf4p1aogGAopqx
JM3mPK706WkNOJvZeQ2bZBS4uKqy0gpTrXC9j2BI3HWDLRPpyPn/d9MHObEZxU4q
tqUe/aNWz+IpN484WRusBFh0yLCzKDu0pvLM3GthG42c56ZXJx6hmS1PnxAqVKho
c5STdRkmkrT6qLZs+5zcFsVj2olOzSPkdt+Mc2GX330hq4Ov8zQLdfXilDou6oew
2cGNmlNsWbCHiar4er0mOdCFjJrsVMhu2vAktLklx/3uu2DZnDuPydmUygVrmu1/
vBBgpspVYcqnwxYR5YTA/BzXcDi9qBpUeKlyLolnLRITz92sK3F+QquI6h2Fb7ek
emU6LhfXBlUVaPSX2EYJfXvi1iU/lYcoAFdi9j/sz0Aw8FnHM7YHjy9P7OOplx9J
1/0rsDGe6EPz9HEa5Y7eqg1O5ddlKKFZQx5WuY/wzt5UCcgiH2qCN/iRsyQNSmqO
0s+IwiIqdv7/eBznJUcpGa3mzN2ETqyI6UJo3XrtKYtM+WOA//071cSvG7FNmvzW
y2hXJpzQCpQvao6Erxz0JlQ3mtcP8EBrE5UvlXtmWTHSWVaa5Wr3hYut4UctlckH
zBlDN4SYWbklfN86+diGLmmM2K5aO0NNuqvDBRaLsVp6YDZqNP7O8YAggLJMY7rO
9i4KtzIqi1s/7f1fTKcbgkZDsjGoGtmW5f1Uep4d7XCsfqXnxisvSHg131ILPFh0
DavIcjO6WOP1yq3VTNvrYYOdZyupdVr6WpRAXb+qJdrPLvWQscBA6VR5VkkMNibB
l7reb87gKxzQ127svwoKOqa0iC6yT5wfhQ8lHQ/0tiW7UnSOmKQdZ7aRytOUDXQk
TFFzLpnyTuupiCGgjErjs7j81X+OqxXgAMN7Xg7HrQ6svtlhCB+Q+yI1/vlEhaYO
xcNwQzAMflcDx3lCKlTRiBkVvloKqKXF5tcM5XuUzfRG2tyExm+OGlF6JDW35Qsl
U5y5o7g0j7fngx1ft+vGVYAH92DoVs/cL/NgMu0oFtM+zrT/+260vT/Qr2TLfNtS
ll2I5t/lfILY73fCn0VJ2XRy85xsnZJBcC32IWf1F+2cYIbmBO6aUyXmqwfMLmxk
TE9pc3c7gWkNgrVFUZ9tuKENre8+L6LDV+f/n5Qt3m6yL5F+ICvLXIZXP+b5e5/W
uu9UuTHNp19PokX44I9/4WdC3RqCEHFv/2sUzlDdd++4uMwK6EeoL1p17csOfyDL
wEkscQp5oTwgaWtaQrqZ/XTy2lPzaxwBwkk7vMarCVV53dxGBi0kCqCupYD08pFA
ticR7IvDngklA7c1+BNB2AwZj66hTecygSOu+nC3aBVSLxO8t8DkbeK/9mgCIB+o
1aoDcmoodm1mM1H3iYZki6H68dkZW5hNqrlQTJSaMrbuaV8BS509NeGV+6xNngt2
NIOdjhRHxOEyzlWvYU0D5m8bbPOwfBquebzji25azdxFHy/eLW7htrShdWPwR4UL
0I5g4CedEbb5P2aLvjqVzjvzMTQYSnq3YYrXihm24LwRaHWGhrT0yAQWaSBihLea
8DzuTad4iLmY9vqgj1PkM+24bfwu/obfBXGXfde/hWxR8Fzp4D/0C7O0Vow75e7b
/s81UWKNrjhGde0vScuta0G/1FBMD3imrCL2B7JaUSytrvd6jr13Gdq3ZFV9kVmb
ravIEReUBhe38mv2rchdAuynHakxeDjjontoouEBhA2akFbrn4W9K0l+Vy/aTAWt
8oiPt+QzSuBIwChAS2e2vzgh5xRvtxfd9mxd/u4d+EC7O+11xFNiaBTsDu1EXYOb
Spw4wKoUDGD+ahlV/8r6OO2HWU1XbEs12R2ys7UBznrDZZFbAkoMsgGxiZYbXEPI
sKucVEWSd/qZFUU1ZEsYRwveiu97jDYneCuzKIR4If1V2nxmBX3a7fFNnc8veFmS
/BbMzCnso5R569LzKAlwTdl7hFkyRRQfDTK7cCeEHtbpJF/G5s2WQE5je5CwJdR7
l949jYCqGlxOvRT3PuQ1tLkZk575ve4ifhVydiCPsWuYhITLqtpISWg1lE1jj3Dt
8ybFXR97VJGJQkEtyWkGHZxXIeGOyBOpyYXn690ZBAAAe0Chlt/ra8ajUDcXh2pV
+3C+FsTlZ5V4FeAFGbY1u0HceZyf0rO3wv70I87NPOJ4nnaXF/OHL/MKWV9EN/Jo
wQx+sjBFhPSb8mklRwbBTsB5hv+97jrvq7nlId4OwOgnwmACo7AEFl9Z++0jkott
/obB6nPV/hp39eBdCHqjhwgaTidJgy5N3KZ09vIClAa57a4n1+I5JBrfUWpfhYMy
CQhirchINxnEGK84iCMUL2iAkc2pM9NFTD4YwIcSlA8bKsPqklYfeTtYvUG2wcql
GzwqOc2TSYUuGaO+qaVAI6atWqKpR9OmC28JWFApHyg2IyADt+/gHliCi85ToT/x
FyQIgA17Can6ae2TGYpb2BAEOvpsMM3JC1cs7pze1DxOcxZn426o2/KeOZv1cwS5
UjWGTS9PO5o3crWBG4z4Fv7FC4R8CJePfghhLMrWe3T7TALJ8lTBXIzYFyDtbnPZ
zDnjC1FlAM4HJikjRE/KSJWco0BLctp6IWdaCYKsjmRm2DhPZqyX66DvGf02ld/h
ciJpQUDjJmHeYXj5V/GZa7rhoOYFE+/58whcaooc05AhaB5SXRxL2mrNo9C4WRbu
4mdEJTm/uOBjpWf0laaHCYGtJx4tiS7EvBAuRJZqG0yAtRE2ZX8S7Je5VIFg06Qk
o4OrmHXNSHBrP1Wf6hh7d/VzLovL7tkXYnEmNKMC7mA3l85+GyjPfvFNcPWBrleS
joWwq3aieuwc4IP6S2crm1cd8AhfYhPKxhTgHXnBf+i86KlFfFDVJ5gsUmZTxROE
LzCrc3zQI/+4A0nxPZaee/c/mqV5t+2VTAc7HDgPr5ik06HEuMfadisizWb1LG15
JHhJvCX55xtu1dOg9Bs6Z1cyEpIOnaJrK+cs9Wv6K086VcqNWAMr0KYqk9yKq4oh
3V9MDUTBUs1jLpaM/0u+uqOo35e0OyKrDNnMkmLIB2fKQtChjjRPUBqnkZt0aetI
Pl67ZAAWzvCuowuXtW87Aq1Z6UAFVKt8Yq5v2aTUIZyTrK2h65wauJsN2iLAFm0L
CNJ93fuRHKyudK5zyk5yPBXwWzPhY+mzdR8xrQDmYjvYsPpwPXiwJwpiFPF4h+1X
cPDA3zXSehz+W4EsB/UJzgm7IhENjJno1G8tACpNIEF5/El5xj86vzd7jzTciNkJ
1vZlBcEKHnfoLCDZsI6jAHnRF3kOZdChaWVuSK89fu21jkKUwDhd1GFjNKss7tSH
cg8KoX/r+AvH6ptN1yZTC55p99ikOC0YuViOUjqGE6Cphhc4hNDymLYPJlgo14od
ARbpOO3S41W7oexlKGcfwtNYa8NhsRFvehwh+XcbTQ+0AGVh5LKr/jFIZWjE7lLv
oJnOtNtcHqQ7b1FLuzgZQR30ALG/9WAKEgM2BBJGpS7TWy8Y1FihHjaASJ2vZcOm
okOBVlct5M6E32Fnxd4FZ71doNSIlG6OHvV1jM3t4myymEGFVKHgGssDEOyTl10G
y50gDUoJWay5xkjprQrovAulpQT+DuSLpiTZkM+8Josbju5qb4IJVmUu2O23xUJz
HesVoq2Z7WIvROE01MpbCuMBuuQzItUWDG7Tjdy+QJSlap1oTGM8hmJqRukaGYmH
xf1jIdEnhzd8Dsn2z50p/Vqg25skOX2Mp0Ii5AXTizgGH9em6tpvpK3mBGezgmos
sE1Ot4V6cO0nuRRux/C1+Xlp/1iVLTRA547QwqSk24E/SEqGgwhc6+SxVRVjMZgL
DJnOlS5JnkNaFkvYU/e8K8YXPpk2rsZWLrm/OLMnRVs0/HguH4uo9ajsfAJ5iEtN
onei53VzavxrajO0eSf5w/VDt2MHG7lJgi0+nSBG/I6DiqvGgXsdjHsupHfpwlqi
q2iuG0QJondkuVPfdEixptQ7Hmcbi6DwJSTGRF57OXz/pqg2ZhqgRY0Xq2f5L/lw
wg47+kTtHdVrusKk65NxXW3irqBlblWO0UqfIsvd093/4faaIx3gtYKRhoIRujs8
G+vyD5C/NiaaATwmhF9QyjJbauO+EKA8Fl84FXd0cKxBvq3EFPacVlNw/l2m8JIf
fKC0baNnLP82M82GG8vjrc+eSK6GWfHUtw3Go/qfyZHsmNJv+uZAvogQgcup8eNc
xKjlHJ4LYzfNEqoNm0B/3j8lKGV6ozzeu71achHWWsYZpRx2OknC3tOPyEe0hoKo
1zgx0XGVrwlE6sVsqj4QjCQqvNEeLo9FIS29nrEDQAIWRAk1gEpWisI3N4nqWzUz
i4YDZvujHOms8z2yITQTozqsZmgPGflj4pQHHAdq4299HFzCeNp9tGpK3DYncieR
mfSLgdT2/nmQ4I7a9XPnzQKffIBT4z3v5cy4g/QG8i4GB/T1fnzcU3wW3Ygox4Zf
o61FUz0tRHMJC2gJC8cSi4OCXYuHBhu7zRtsyqcmf4+RgKXzCRIChwuZcwa9VaJE
j8iead93RZCmQWf9KasDSFhhdAKVHCGmvfhTL49++bfl7Ea4wE4L4DlDgd9B7CGr
xUyrkZoISc77vyF7xP15NquqHGdrDZI5wtWAdR4VZg/ttijVTQcr4K+KEQ3b0CKq
WhOSrwWzZnwWt9wI3l/B/Ruq71tqCYuTNnDNGJg+/VhArsXoMjysPiIRh39+fwpH
7CCy1NT5ujgqxC2MxwchnKA3G3g+rDJSqJsvaF1ARAZiBVKaVVW11e18pasVjSil
D3/A+hPDpcMPZsrjcCwIWNB+QE2BrUZ+RlTMCpQuP5HX47w/0FysyHF7qOVtWwn/
leSUN1H2GbsGQseJDYTHO2gqJMYB3GT/ODiOr5qbAH7Ak0MQYuAtP2/jDjQg+sj3
44ckN+C7wAmCKODP6npIdf55EaHPgyNRBIg6yt8N4PU5X31oE0dgoUOYqEfffC1h
XFc9VLSYuwbPayMX7FbDnDnz7cgyG5YNEftPOh4PDcjvzu6pZvnxDnR3VxuwLvHN
zmo0LfQY+DSEJmqDJCF72WoZnootPUw1tf/iqeus4htk0ydrv/u6ZB0j1+eH1J54
DXZliXIJbjLeMOB8r32uxM0gNXq8RI3nK/LFM3vUA6s/4Tsl3Ht+OlZhd6Ct5eUi
4hi7QYx96D9nFGssFRuwSJTVDUwgMyuNBZu8eEIgrXFmcoZH4+HF8GPyDWeoitsn
VHqFR6ImY6TPwQpAi1m8yWcEfLBlY+EP0T7l2p01yoJCjLTA8sQocuXR/8VdpayS
fJKbxkp8cn9MIHO/MWlOoZMt12UlJ0JIkFfNvoyWXs+h1KyKnaLgwqQ3FEiLZj0w
BlQSE6j2dml6GtKGLpu8OIsuR0j2MaB+1g6+wXOCabLefExyCHAQs+CxRvSXjaqp
zhLwuAzzji0xdi3M4sMpSBUiID0haq3FUtkL4NmnQ6adfQHRwQwTfTO/jH5XogH0
ARZsuM2U6hPnAD6UBEltQU4WxfImdJr9RZ3yS/Ckheo0jzBIvXX4zS8xejrS3kD+
jZQ/9y0BsWGlI3pnRZFW667Ju5esMoq16U/qKl8LcSY4zpd0TxdIQnZml3FQjU9Y
jIlTl4p8nS/jyg5czL7XmE20Qb1Adm+KEQ7+5ygZQGX9opJmjEUdxbBFqoJcsANw
+FKH3+Zd16x1PmBoDi2t4mW/javUjYBG3v0s0og5kcDYFhS7QCK5+UimG77Y27On
F9WBDi36xGXkbUhwxxqus4kNlO41xjxU0Lsm6K/ViyCjxCRBhON6zRANKJkfhXvX
nDpCLm+IfDxaaS1uHF/l4o7Kzm8Tu7V/ZPTBftAIRBLJ73TQ6WPUBid5/yhn9LjG
UVKw+JdX/ymkF8Yiwif+4S82M4EmBsS1AbhdNIRaXGG+FVWaW2PELurzTrpqfA9c
iGD4wcMdhf9M3iSTc0Ek2P6NHd47Bk8FubRi9AwXAiibYbYcCulp2nwdHRZF/8VA
VkN+KV5QaBFqAgmvbAzCVmZNxzlmh/i41UpwBVQGnfi7eauzAYDPAK42wJcMK228
EGne8iwK/48+QNkXETctLKVySjLcZlG/N+3CUVSLnTuNLp3IYFureYQuo6r7qkfo
MW+heiZMcZv2pdoLjQ/5+XBQYNymdpGcuV5tNe9FZG5uZgqkIweI2HAWIDWf2a90
UdWStouSzyMUpdFlDauZVDgbuGzOi5mBh1cC26IjaCatgjZxeWF6hiOY5wazX+yo
ZmwdKuQTYwyUPeme3b+eud+iqU/3ATo9DHEhnVphFPSXGrbw02LHTnQ2kZwCEWKZ
IqNETV+6TByCXYkle3VjXPJ4SAFjH/sKU50ihEkjDcvy9q/AFCDsgHK3yyfzmMyx
+bB+q5wj/ABeXWHFX21Oh0tQq+z8eyzshlufGzDKoxRg4JGiUwgD1HHcieGroGpj
57B0VF9rrUTNhEsnzsR61UGrjic6AKvy79bOQnae9YxxXMITqNt+U7RSBoX7Z+KO
uP6mZja82vDFCGJBnOugxl3XmHoEGL3VJ6kwNMZxMPa7n0FenQDbmHvcm0jqxrJc
imyE9wHkeuJVCXARkucX/GP11RUayPhvb5oSxSXcNSJOcdNzOe/Y5vEp+re/MxG6
XUbfPPo9gfInYW9VgYTpzbtMbR5uwY9b7aVtvOFjdWqZT9ESFPSU+UlVlf6y0une
e8vSH1IFUuYm+khoFXIlOWOkB1cO2CW+wA1L4Af59/RTilnPbswbWxw0OkXgrED8
Qzy+AIKt0nVKhKUARDx2swkhTul3MSlrnETr9W3qFx7734gP3b0IuAlFcD42+UZf
y7MJK+TpLnQa2/Xn7R/IKbar569QrEiJ7GxDaGC1rJ7/xpp4V0IqWibnlKByRtEh
ivl5d5VSGkmYWjXRfCqK8A8lY/gtWHg5sgtlmiBfoqTIgpstom1xQhNVDVzwuxlg
hXZ+4cGXkqfWp5eW3ef/taAFCkNHogWL5VOXs9ZDVIpf6gEfoDLfdO+G2fLTs6u4
BdrUPz2G0J3ppRHJKumwP0+ePD1BWE4yGC1c0UcpuemsavQ2TaYlk1nvGb9GzRNO
RW9sb3mkJkfNhZctsF/cJwNCtgZvxlV7v2+/yTtlLYZ/+L/LnqxPZ9imglYQQ7PQ
lh4mVBcNfLH2dTk4+pgHrQnLYKTu6BOzUZyRsipQBPFzh4roKUdN07j3HbZhDgIM
GreTumbuP2F/mzHUan/b0YheI/JGWe87enKhg82IvOIb8x5ZiSk6XbE+Q5CW3Lbk
hfq8u6i1yfJH5ennVMUeRrbYP0kA4REsKr12AGG0okD9zjlBBNGUG0r0x8iK/NZp
miPXCJqaF39/dn13erAp/mUs3PhgkqGyzRgpFuASke3v3Fhe68r24MAqBq9VKq7c
ahhis7pSJlVojL5Ti5IR+t94hM+2uzj8t1wNRy6wI2LdWWdJhAfhCeD3y8iv83bf
2PeXsBmxeJU6/m2iRZIIsPUc9ngyFaKfKq6q3JKGM+Cmzlrtw9z3FLDe/3T0TM9D
C8mFdcpEf7e+VookMeLmQ40dc/QzKIqQYa9gBu0BzlVgUARyWnBeKLGY4VgTmgjf
DJSsu+CxlaeGjg08pSIj1ktROvyUzH9LRH/lIKminPy1jI+LOvXS+Im3YGcLEVQL
Ar7MmcXFIu+xTnxGcdlVVDiwHeHq2aqrvA7Q98xKyRSZWwsbEkWt0bVA1jVHwrPG
n90pd6/oqZ2eoIjFRO+gdLs2ZPiG+GAgKnzkY8i6zfdCX6qnwmWS1KwiRodM2+CM
88Wm33vZi7iQgHzU1le8Ufc0GhDO2/dVbe4B9MRVsZAzvZ67n9a0y9uxgzeULZcu
l1BULkUB+n62TGcyy8QFJk1AjzTtQvkHXMXRwtxMVys/VQ3JhiLr4TQ5uWeGd9Tj
WNbn5WLhvWCE3T/3Hc2w1nCBp10f3TRGVbwnA6yn42U69lLpPhNAJVWSQwm6caWm
u1Bydm9cF5XobQ5V4wqEQOVfgCTerbgmhuuO28U4Z3DCd3qSEekO5O8mA9LagCFb
pc9JVQZ73fvcytBwxuG5g0uyzzjYg/Xl94F7K2uj4gPQkh/0o6HmwwWNvkVTtGq0
MFpBn6R7P/6zZnWsWu+i6hWYqpaGVChX5cZLxXa1zc4IStnGz9pPetmc68uxSNZX
LTLzlcvvaUD35/0ohXNhIQVJy202Hl5An7qxJ7JPnBsSGj7mRPYMDFBGRDmCUyKR
QS9kQIALwjh3GHGqsIDV/NNCUjIv0oZ9k7ZDX1kN5cUY/iMWNpaWA50SSmm2o8TF
9ONkKWvmCbaUSo6erClG1CSQpY0y6p1RFuQdJA3RoKf3dbBj4mB9tWJ8qPZQJZYq
9FBXuysyPFv50R61o4s1AkvGyR+Weu990Z6v+cZ+WXxqzru2D9mtTba3xeOKVXQP
AE7TUz99+O2q92ZW8haQ6zQWyYxLd7+k3D5vh7U0/m+hT1JFUG3ZDBhmt5BkIFw+
Qu19V/WZihJP2RVpgSbgL69+46DXVeB/Aw2wfL34BPKmOtfmS6oKz886/H2ht+5L
xMFNuQ4Zm7x7o+t+l75NMoOcYGMBz1tZ2Iss55KhJjYC/SSCFqwEHEUyJYtehRXE
YoMr5QOp1BX34ecc/aNT0X1PikT565hCe4fdMxxEuQbI7JVhDE4+qOp7APQcDBgv
VvK2B9lbeCckwp5Et5QsSuhhic2B+mK5FloNYjg5yHHLhhVzzm+UbwQGdm/FODLO
9/2TE9rK3XH0ZCgpcFD00GcHLxhZhMJ42hEm5USBhNf7ejdkAdO+lGC3P2g8Dmp5
VDoyHY6qpUKc74LZW37mqfv6TbKmmVpQvqt19by9xRAyGWNnQf4aZCaQj9t2Djve
W3vBfVcIhZX6mUK65ohDyBYJt+Ff78q3HQvNyuLektDQL5oMEKCVG+yKY9B3Pcew
LV7x8IBxVfIzx7Szbr2zDXSPlBUPrcHfCLFuJBfICC45hFjjRzEjhrBWdOJaqBXn
py5/1MrIbXnhU5SOK1AE9fM9x9rT0EcDm1qdA5kOcHs7pCgfyN9ZEHGEa0e+2QZZ
ZAQ01BvYyeYLJl31cM2D3kB4veLBWZ5CZ5FoFlOxHq0QufnUPFSrfnjsCa3a2FVV
PfyD9psWfGic+RzrQpxs9+4XZ6WV3gd9eg5G9JBdVLQYIh0T+PQMeBK2o+SHKYjR
Iimga5a++uol76RjS+268VHPms0qxzYLfpLXs3OaRDEjkoIq9x7OSzVVlCb6OE1V
ni8HpDTxOjS5zqHRWNX3ReC3LWqf6DGjX3LeHLNp9J4whZUpS7GVsJIhdNAlJEAM
erSw4YH17Jqh5LWvOymIybEpHbaFpkGFj4Q1obWKk2r/8TJR4JwNtTFeKvDf2FnA
X+Jx+eDTRd+x0+llPo7xmoU4xhKz5K9tb6GYaLhFSzD1gsl8i9hpUHdxE9Nq2poj
xXUG0M7Wh7qjBW1CAwWeT9C2/kHN1CumcN6ZU/1X0FbWCLXSAG//qHBVEjwHiWSf
TMiuqFR+EerXLuyUyst1CR3zLQOVlpJhZVMnZfkQUUI4hWarSTAZtrP0bYRibXVG
YE4A7Ldx/naiILCSNSav3fZdR/2xjnjpNkibgJ88j8Znu5xS8KQI3Ru7ULS4r9k+
wHBsrgUvx1LfIV6jDjVRSZZ8riHIv29WxXiD2t3Ai2gBPMLbol9WN2Rxg0qsShhE
cXtSHoXZt2TnlL5WC7SWeUeZhwyvxKHoOfnZoPAKVXABzgWWiWofHxBEEoGjvof9
JU2h+RLyeff2Y5oU0W73DjxqWD3D2cPr+l6dRn43Pc7gZqGP+RUXvu3qLxQlZBNA
AQCySptEWI3kjOa8tuiLHtwy/nc6cn7UbCXh9RgC17+SJD/dMnPKfVebxr8kJN0H
FYj+eRoQAiLr+yB3KeF0ZBwxDhYWphSok3K2hcMN7VAhud5TqJFj58l3FHsTb868
iMoAxfdHzThBM/JTFryKXDoX7QzsPdPwO8IirG+qS0u0tg8gyDSB/QaKmz0ZJhsK
2IHa5vKZ9xaRqdBHVH/IjORqAkGGY4XgSL10lqc7gB8h+dDbtOBVH8TOvwkuQvyj
FJORpXngfO3MlETFa8eC+ayALKjmHabXI4oIxU8CpMmCZr/Wwa3e2EischSMK9PM
7eaeoUMJve7m/hn8aBe/Qgw4rYPilj+7L+1mE0iOKAOPTWAcAIPAbzo3bLwNdjiv
gkmPb3g2aJjMAJi2SwIqSXVpz08hDsqAvq4nKsLjKsCs8pFbcHidIKJs8LqzcFQE
6K12U8zmF5L0rj7D0fG0j42UA9pv4KgTROPN1YKCUgBcReK1u4TaNUH9sk2mLT4M
ho8X4ZrSqerjO9zKprUm6b6eDr2U01r3EnIKPcZzFMtRkDjbjEtJMVtZQNbPNqih
xwuaopmQoQXiArDh7/Myhp70jG6Z/ozrt3P5GPsq83kRzym7zvVcDEN6XUEqg2ZF
876zAEQW2UwIck/tUvXCQ3MzBlFUsrTUu+gYLHKTUYY1zIyzMEMRQaKzQAKwblS/
dzI/8dVdS7Xc2Pp+8ZBdmoACed6UTA9nBeDjPPJlD1H2FJZ7TbWygYtXKVwL8TPQ
fkbBEWceMXgszFFzgmBlGKuSi/PAT43l6Ma4LZT1tE/uHclUKsh76+3novHKv1Lk
uYN4ohv4+qx72LC/vsP03ogzHXQ/qbquwU6hUmrJF3hxSggYahqnjTVjFK5j1qJT
ZJlTvpBH3moXEW8jUv2bHkh2aooYyXFmTvSNo9jBruQ15j95NjU8gfwo9HZg36Dy
8AFG6RX53gL6AHF2hc216Hbmc+ZP78ipH5qaktCPlS/66cPSzZXG9VxNYyIqd/CQ
ZpP2IXkCjCS/J28VQoGPmTEDl/NfBunTH1y9xjVO1FSioVxSPlBuhglTHjfBrFSU
3e3NAv/4CjjzN9bkqsDch9IX4azixkazBJFN2uke7RJx+bnhIUpLYO21M2qr5Ttn
nTZBj7+kazi0rSpO0b9uIfk8w1Kur8xbxJgUjnJxpTLgngeeJvPWurtgn91Qq7JJ
yu5fwdcsL52WMSmIzNmTyladWRNUGpa7Kk+CIkeRMnsrvEM7mjqJsfY1uEHATw+h
ydiWUTEqTCxbNA61ZHyx63eB1ELV25bG+OhBGZzUiTNLBBQOHJqzGEjGn3yvF0f6
azzPpf8QlQuEEkxlxhM5J+i4wekAiz8on+T+mB5MZ0V46tqe/S1ngN8tqkzmxChF
Tn0TBTeltr4uFHIsn8fUD7jtM8Ogp/u7rLrFMmW0HYGwxVuP3Q6ohxoxfieQ7/TZ
yMrpdCOr3fcZFAFUnu1KvIs3BYPD3nMtaZkkUSw93ssg9trwVkw2kMwJYeD39HMr
izbQe1Bx3msedS665yyfJN9zG+udClvA9Sb7CqM7PfK9VBJqkdFtYA+qxxBknDKV
2qrwm6S/88Elp1jXgdHbcE9SI57vXl5BonWk+LOwP5Oul2j+IxyS5wbDUWe+8nvT
0n6m+tvxqSOfQ2XkffX0blRn5zLQiNzXEBSu9nhX99zL3+liu7yZZaXPOirNWzeU
MxvIF4VNrQWCknvJ7K8O/pHt67FoCAq4MEsTAtiTlmz/uunxtHBRQjxRdxmo+zlZ
5r2/Z+FfY/sS4JQtXAwDIdFArazNJXy09OqII9DGVLG94dg2ZpCcbiC7nzZax41O
pTo6+r8suekOuxdNhDzUYz5RAk5DF0xvn67ePxGtxTKlHkUuwjCKBUa4WQ/NbNHf
AFQQj9r/UYR1RjI8fC6UYaALiAdyT+Bcn2n+exd0thchpdZk/nuWm/m3GGha4mVB
Rs7sz9EB+E/HnyeXIYJvJoUQ0msxdBBl48ooX6BRJFSdxcrs/sGCbTqESVt3G0Dc
0VKn78m4bMVUHiIvoz1hH9qhk5mq6wtqrjyTZgvXhKx394Edy3xMqdtPXDMVKryr
jMWrlvOnwa8/jx+9n9Y/kxZh38xC0QiTRkiFowtOUMGrMW/BXvh/yNVmY8uz5u18
nOcdWT0pJfQ1jQSlhBRSJhqSRnx+jt+gBmvSnzh1g4KUMvznArKfFFCWun50y5WI
vLIFj2IzXkPfdRlbwcHc5x+nESnae+8CY7BkghmKLK654Z9zRlvfBb0onR1G3h08
wVCHtUWcFDoNRwjN+cQeKiO7EseDg3xZsm/6j/VzKw7HkONvT9s67bcHgapA5J7q
PSJXzqR3MK+mKF5788FFdeEWO50arGIMhyKNFOfPx3K7yWZErh2aSStcXa2pglWB
ffhYY0rWek/clgDrr6L7wBBUBSY//AMOCuJ88XK/zWK1I6Y6muaS7rcn13cO1p/p
Lt1bY+rHufE8P9AX+WCkSCw/e65bRYCpw1Kbh52VG59hwrrxGylZe45e9YZrHqk9
3a+8Xc3cSgYcfGzTDk/S/OsOeb/+kxBSHPBY62y7ZVoCqzc4gcYMhKne5Xifoo8D
+iUez/EN3mbJBBOSuElJIDMGquXqhnBczMbD6KAB+PlCLTB24naV6THI8v1RadcB
rtt51x6DyT2ZhJSNyuIV1lgkUdzcZArin5ZYgRnJQ70bXRXNmVnxBERS/X+R4J5J
UTcQcDPMzItk5itD/0bcSCelxmeuggXqAIRUI2ML60bD64SmAtO4XgTmx/sO/Umu
oWjO0tgyYAIByGhNWE3LGB4oXu5OF7B/RRCfPbk118n5wlxdd2DpfYe8NpJnJuo7
MT0aJPt2e6OhC9NkSvKzxADRHUvb+ddvsgbNM/NSTiKf9JhLBPvCvTcbGmGECvpR
E0Z9qc9gBPx3cXRDlU+teoH08nGb3M2CwNX+6LBXyEnCVoakytdZKcr2Zb+uReau
bw/L+qTPXSfR4WralhlVg9k1Lg0u9965RhIbiIQReCUt4ndmTP5QXJVfQv0btr9J
rX8nZtVlyhD2qr6d0qk7XE4RYxxuVNnDPIsDya00QA5QX0oG54T8X6UsHvbdeSm/
t22gP4jK+zWJ752GsffO6yVWcxv4WPnC4A5lqsUNxWXCPxDoYetxwCCMRZtLzK52
EmZiEhJ6D4dUuKQrYo/Xcmk81fALS+P2sBYu/u897O1jgHVZ2mbso4AlQtB7E2Ap
sQDJ9b9jQ4RkXxkPRoonE7jAU/tUfuIGC0fWiqunYPcnydpLUay1/SksuJT1nXPc
WYsPOyaWKxuToq/pVe3MoRNinm3NdvCB39IQinZMP9gzPjn3DT8N2l4Azjvqc+f5
S/jgxl8JhNVO6GoKczT2BaGmzfa504icfoZBkYW6AFuPPNrKViIQ9tCDpg6pblGe
JA2J9JsWbf6+3r3edYoxgmVEI0UCRVZuoa4GiZSxZUTpt9HcXjv09WHILF2//9qs
ej7yU8+npczFAwGI6X3VsikgI2nAPogPQK12IvO9JNLOOvqH5EfJtdfLr1qAoEJl
4MYNWmGCFX43lh0L1NwOW9P8TwcQchF7uR5C++QippSXwhexB1oFKFhLWdhc7/Ou
YyL2aM4xj0Nzz07hYAFFToaBaD+EQyZ6KTJD3IaDhCnBzmAkE81O0kPTv36R5jvY
4ufiQGBvnt1/Nd9yiydP8AyOG0bhuIpf7XjN0GNRTVMBLtYlubpK3ArYVlZrGWHA
qHORsFPsqNJnaUx5X1LqJ9UgYZcyha5BoZOvpfP19WUdw0LvyIJp/KNKdu0Fxy9S
amQISlx+C3+udJp+pJnK7uY3aOko4HAVoGr/wHfhiTshxoUgYf5ApIFCKfUpWu40
A92WS4VG5FjeYdi14NbWVq/O73iDfh6WYHjGKABUQyVKhLXSSeu8TTYYamZ48tiQ
dnHxDk3GKi/ovUA/e6SzUZ0oENBUj004fIxMCQB0AY+C7jTBE0IOa5yuk7TdgW1A
8lwG0imL6zOljyLYAp71rp0yJZVGP8MAewEJ10Vwr42WFK4UGINXtsT0GQ3FsnPk
sNzjcboSdRJ+jHOfMJiQ1qOOHxQjPloceLQCgMB3h10uiIyWQLG2KGw+5nF6DDOW
i+LNONw6oxbVnOaYpXRwideLoG2i5iM8f4Kf0pv6LNeME9zSSQfvIN82KWUNYkWL
qsfxeteqL0xt8UxIhhTqsJpxrIgQG1HD/hhRRJAulCJl5p4eXcim/xPErHb01hV9
XIxnK44TmhO9AAStIBs6yGx/WoM6NTaT9OqS1MJ1Ve8WVX8uQnAgGOjB8vqwRUId
/6SQeA6Cr+upHihdUrjtZ32p5Uauf8Bs8QvWUpxn69nOuqaRhKIGUK+qGjyC31gx
k4L8THUYGXxLwuv5Mk0QYJfFrPYRsO6sE0MZZrt2HT64/vLEMeC5j3IO6b2+P5AY
4zWChafu3P29hzTj1OBr3ruU5aNyxSsyS2DJhutr4QmDI8vDuu+pW+AyJApvM+Q6
qXXfIIBi3c10l5nLD97ie7lb+cJiFBsChe8rj/mmjjqTaI5FGLPZRQySF1YamlOc
5WAe48BcjFbbNMQmtI8VUAGcTHb6l0qdJLXRN5gZR0j50SFI1TIbxMMc89oJqWZx
auuq3ql4FIF5pBR2MG3h1NYdeBgK60Bn4lOxJITE4GUX6o40HObCns97AIk8fTUg
w3ee/S0Hsms+SmleZZruLwC8kpKEznX71KzyaFMNl2DSyx2VEgcMqom0hGwBMoSM
pEM0sIPqGFYjQokQ2w7XzHTwAddi9QrX4bQd3bgPb2oZnUVf0E5erbsNKcCYRzfB
WG7motjAdGO5OZ90SBr0mvE5FZK+i7K8vSbcT99/zR5ncS3ZE654rxHXhusJLE+N
ZK+0PkP7hylBJ34U0FgWCHXAg8mcGraal8VybKrloIzjiZ4WHdwmt2vMTp1KTbLG
nO9wlJ91icmebezG08/qMzYGeuUpnmi76AVr2mdd9upT9FFcvN7LLsQBCADRkCTJ
sgcmlHaCITHLcb63eLCf63MkD7lvv4GWN08WGEWGIE5+1S0rfOWUbyi0f3s7fsVf
LGX8D2JJZOxUG5rRf5x/DOTYh2NJff/wyfBqtjuFUitsuONDawElST8WiYwXwiPZ
PKkYiPgAz8fmC0h+DYYkvJwL+5P2p0ARy1qkLfYkGDKhkQ5WaAti2pnIVmjz72WF
xKzyfm2rTUkaeUPZK7NI4v8eAvsOVsOusR6IzEmLUVZvnF75e8LnvqtiqRMncsmU
EW2YThKmFSnB0Y1uLOWo7vkz9iuMS/L1zJme3g2cBrk1xdfhbmgVnY91pRfDuCkk
vDaUi9zVy9iBRHwEcv8CrNqEcWCzrothQDuKrBTGl4ykaXOJ2VzTrF7QL/MBNnl8
q8uprI84UQGj+f2dv9FTxjsrL2t1K/B4JTkQrzw76czslp13+2d5VMWUanCBPoVz
U7rE4KBg9wKnEt6nJupZsN7Wmnahh2WFfJPaJuH08RCZxpRWN+k+dcWDvNQTqceB
XrGnii5ZM0kdIz9X7tixpQZcZsFAbi/D8LSK1MX0vM2vE64zo3ZOfmcHdGBme2QU
8DZf3PpSMbSYaMbnyxGSHHbjY9lA7TuIvPWIm9ztyw2AR1dS2wQZl4jFNPrALdZu
YJtxS2mWB7urGd9sJW1ikJBHp0fGNI1RC55gYdsZ0rQaH+D64eDhSmTZ2tayINb5
wJBvHj1KmQY+/nJSSwLIFOZ6MNhIpVqoncdYLgMHfNOy1KNpxRWGXB/VfXLeW2Bi
jt8WsYa3NvrrV3eWiecfXPBm+1MJjyBkhGTGKRjqgTmL8Pv6hrSTKIp2WVGvU+ja
FOSWUKAk3Bb1Hw8714sSSxb68Sotnvh4MqpgiDF7Az6rigvvXHOJN3sH8LP2p0R/
9jkr4txRIN7mzhFq1WFA9cdos2XN3G51aeqijescBCFovTBjn7nB1lm2DtEaXRfv
2LwNeA5XnGbGCI1M8BkQ2k2mZFHEwxQcnMQCMEX+MB5udjZXrLd9Vco9VKINFxDC
oc+i8qHGLBNTuH/YhrXj4q6uHz6SKs8TGML5lCuCsV+j1/avhShz4Jd6YXO32OGl
CXPaXDahjePu4QapkwyOa8Pp3VpspCxbrZmW1l4k7N4hn8Pyqp3qrNLSkfZZ3cs5
H//iAfEV9bTH7K9ofDqjWrEtlDzoziUf1jSc9DMZDUIUTVeR+JJvj+6Y1XGgEeFE
ykIHbBKu285EwugOhYT0l0fNN+0OsJ1i2LcYl0mB2bEaNi/5r81oC75s9zMTnmeE
lGNodj2yhRi+tNZo/R2pEfnEjBilNRmU5pEJpq9N04DAtRVR3Q+e4o6R7EbFQ5Lg
UjxofX2glZJ6Dzr9QLIyQwAX2CeIU5+/hxDP1zhzOnWsWMetWzisi7Oqqq3IgJhY
UR8CwtbQGer/jDZxfVHh3XTsBGzayXK9389IO641YP/f9ud1sGL7tRgiJ7hrfPoV
BHLex6f9wKm0tBKChd2qvOcYuDHLLt9Zf0ip/Q8+Rslt4bYzWy/B8JdWXcwip1jI
t/EH9BpmFrlSkibE/sDqJGLGDz0XLyiKEhNdbYv9oM/H7KoOUYDifldJeeJGggu+
V5Dzs73TxFLNuyGaQg05rg==
`pragma protect end_protected
