// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:44 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lxacK4VcJka8Xz2ookwmbZb+uvVv1ZdWb2CSu89JT8qICWsGt3HLMHWrpnhv6kGa
LUOrUCAFZtIzIfsi9QbF+z6FNLcHeNxAn3TEw5vAUCgzs/8x6f14HI1si28lVPQI
uYjLYige1JlVj1CXHA2o947ecI13qQV4wZBiA/fGW1k=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7920)
/l3q+y8le84kLraZ1ZQxVY9vmMIciocyQcdpa6Rri04F3uTm5AcO9/jfy5QNI5Gy
npRZ8AMiPAwK9o3Rzz+RRAYfCZR2VPuKs/nSRTP9QeD6RLCQifM/5DIWFD+RsNFe
mo8L059rIW5kpQtKIbEcYJyySZS84HPDwBaeuz2VTWPvhSnhB07F0aFKRrerVLlT
9kfuL5gGIhABlNbt0QzOqgUlDtSu/M9ij5HmTeYEV1o0keh8vcFhpmPKGzAQobry
mC2W8KGrpaDiEffPHKoAiBh8VtkxIWnFClik/tSGCUlAdyRZj9PGDkGiKW3M8up3
Mq5DgxPCHrRaO+OwclQuGocRF4zSa6zhyX9u0r3U+YcvxBhBvPfBTZ6JCJvj+bSF
9MDrl2e58gxjOiQNScgR+9V1wIrt4/PatFQVI6wHPGfw/1QCnG3MnVueSj7RA1m2
s3EWn5Dtuizd+LDsKT3Lt1s7e9PGCWlfM3fUXW1ZKnXS/0DJQOSXYgMqqgjmGLQZ
JELvnQWqsBmsBAhrGwwcNmmPKhLVsjAVA1En0TCoi5A7JPEYCfr3M264zAwzCUsa
HLP24JoFB03yD69COsclvUvz23c4L1nEhP1qoyNHtHdfeOWy0s3p6L1vt24M+dcj
GNmpldy4zp9ZdrCpwApswXBbrhFReKtRcua+Jkb7+3e9OcAP2cRz/dXyPlHvLUbn
2LRtsHg6gtQ9u/gyuaYlh8YE5+6E6I9aJxrAWg0qhz7lcZrqR/Dy5xfQdG5KLznh
u2YRGrcgVAnKWey5JTmJe3O38IUP9nqPNgayFlc6HaT9ueQZ5lHXo7uHmNCVSUrk
Tz9qLEKxyijulDQfWcqCHGQQg+KdYc2rVPZKwooyguLQbPdXvfboQeFST7ayJRk/
PCqDiKwhKPlnL8h+JWy4NxHzD7k6T23ttUZlbwKG2yBlVO2S8Q8yOIo4avtn2Fkt
O1z8KAAvO/dFdeOKWW/1UYavxkqKE8QyRewajYTy8GOQ4on2FIkm7IZhr6QcCJxp
Wk7g/Ja/TEOBjDfoW6eqyNXZF0P4//ryxtVwjlng1WOCIZrLa7v/fMsP4ZdPlGxe
LVPU/AHTnDz1qNcEchWCTXtqyC/9hnJhzahPqgLf9Al5IEQc8PR74m3wIDxjaJHg
fPlEqqU19mmFG82zGMDgJGAioRHN3EZM3dtOCT5MBO6YCms5cEwBQXNdI9vPhfLa
chvEjMG/vyEy/EQ+4DLbKVY15/AV9IubH6DlaAs7cb9ocIw6hPbESeAH2qVhjKHl
JKwTZBTDJRQSHEdT4xXMdGT2VsmAY64Ps40xTGZJ1vkNZ7jNo1+ixPi/Qmly0dWh
S3n8QLrMn2fzTWrXss7yKbItmlrgeE34KvoeUqJCrMCzF0rOuT0xm41Q97dHnsli
ybsoMRmV5eAW8hUkd3JiJCtcNNorZUpbRsFX9fuMyTtthCDAE+Z5aURDHvHvXWfI
Yz7Xg0TYnJRAP7XX1oIBEK60fWQR3RKKygFAARaV0VAPZ8gYlHhahKenNlCFEQok
Ab1qA0ZwBoa6/IWZOwPWjH+2/lryQmYen23X1CUsM5bOzWlVDT0b9AhAvryAsMF6
9IXuMh2HrWReKoL2ddDZmYzDVwc5JLC3C+IeT8NptlYcohz6H1RZb3h/+QZKhTxW
3MOfA+6kPK11H5FSAy431GGNUn6vM19z1ESJa9fq9f649lhxkIyymohXHVeA1bbp
Q+a7FlOYtrNo5sgh2wMFnfvJzoud9OTj2riGv6ojTasd8IHCURU9PRwfNaiQcKno
an7O4CsNmDe0dzrlkLjvPCnEoKF1v8/EcAiJMH/FhH2/xejyf+Yiv1pvQ9UD9iRD
B/DxA1zCq0zZrwiQ6IDJIPy9Zq0okY0OCBpgRstrRfhwYWOKkeZhIwIbfr1qYo2s
/f2rw5kTRJxYcJrFPz47ZfhAPrSFXWJ/HAfAgOVAWny99mWvZEWUlgSiZ83RAAHs
2t39VEnU/kF15Cxi0kVv6Zj7Mq8NLK361PyIYwZ0FxxnyrnymvVJba2ejK1WqT5r
I2bQGlNHhN8h7FAzZAurZPjjNw6rTzPyC5BoppSrpYiHPwhJXXULJgmlBfm1WN1M
WlCevGx4RDe1v1uwzAtsC9vi7bWxT22Up4lk8vmzxVTgPIKMENsGseKFFlSqusc9
0rvl+LXyptS3PP3ArQy2gq0QGAtfMJ7KAGg9TCV3sN9k0TVJ9FuE/um/EDkuxCBu
PIEAOgeJb5zLgsNh7IAjetVQb15t0hykqWyO0vfBpkNxiwQ5R8XGSpoaV/Pu3FnI
6bhzko3oweHD2yxhH3gVMVJUJuOmYF7+LkBAw5f8CUuIK6hQyosziCYbJ755VKDM
HGYjr6UySEPssU2C1IMeQ+mhGNAXUFQa4fa/yioHlWW1AH5ttU4rTDUNYYsTkezk
gWXqTAg4S20NaHl0Ae/8+cGm1RDxsIpGji//yJRh1W8c1N2okpw3nHqVk+V7vGV5
rofwl+2id3ize9yOjdlJWD5HuSy/SBg5v8bHxiEKxGsF21LvY1XtViWRCa9uovL7
Wo7SMrSczf49bU86o2USFy0VXSaXrua8afWv/mzmycabKlGSTkDX9v07wewRh1Rj
jv1ymFEluNK4T0WMb6aED5A9Eyo2A2Bgs0s8fAGg1/pwWgXyVJDzar5zZxVKsyVB
KWzNIFXEMPVNyBydylW4wfiu88hN2oB+MiM6Fz0Yf87Yg9FOr103K5LVYqcbM+6A
sDhpdjqV3+EX75ryGDCF09huK9wn+S7/g/1zqhKWMvp5npTklyS0/CUkYZOlaFB1
fBeFqC6qNzrk02Y+z7NyAz25Dqv1gpVcPCWUGJi+IFtUimvn/iw2CCeI+7V7MJ59
PxajQP0t5qyhO7wh6GLjJs2iWfJDgHKKDVE+W55ChJ8Ps171ZoBUP4OuGiEyf/Xi
YUH7FNLsd59AD7SLQ7WbkkelduoKS5IpAd6yu/74ym8LiDyRvB/L/m9FfgRKqHES
KJKsdKbw+Gok6c9REZa+Tjjp6n638YBhcCpKhB4E+ouvJSuWf3ipSNEE4iu5q9j7
iX+7fFL9uWAxD7sLrmSVV8LAE3nHMnFnc7TbcGsjfbYG9Jf5vtCKIFr3FqPHLua9
/hIwWjD5WCDi5l4xfFrmqs6zcWK4ojD4pooC8iQhiRQgct3Y6oV2myAxeVs+ndjn
BpxoToLuWsVE0dQxG+tO+n4yYYi+AJWC1/2rg2dvRywT1k6z68TZdfqofxcav4E5
7UZx9UoikYMpyRXEUF6bkPAQo/ghuTRFobKv5sdhVMyBdQkz1rPG68swxPe5xpqv
VC/DZfQYzeGTLjHgztJWgQiBy1znVB4o+B9BaxwD8WfZxFXT2srgne/ZblnYPdNt
lwC7Y8vR4fshA2hd064QtnQgDW247ZrrMzMfe+VJTlJiL6JC4dPt3mjGAsspPeIm
DLgcn6pPtZNOKZg4Udp0H36y/jLZ9VbuJLEbZHAZB+e6kmOqhvvgb2B2W1FSUT+E
1VhuY7WmBFmdeGN6+1TqE2dkwvirOSBwgd56wOnOLCNSJZ5r/XbFUc63avYliFoC
vovSHgmdnVA94feYZB3StYVCgd/B0hbWWIopA62SGDaGl5+HUM6JLYDPWReXwR38
GoP3sTopvoEej92op57w+zjYIi0XOYC4KI8zS1EzyzzHwUy3hicdE8JKpU9t45nq
pcQPEfptxH0H3/5OaXPPay0cBXjpAHumGGRKVLRrUbzdFah3Z0NjwCkOrd3OjiPF
q/FToibj1Va9jHcrAeDjI0zcTMLp1Pg/gidWUbpfFVZc2sw2gBAbUt/MYIh6MI7T
51v1VgXrVUPBn4NjOY78wCGmDppXe9lZHPKKKY7PcUKESOnu22Rg0tP+d1jycPX1
ZCQWnSAGdvnHnNypseRDxIjZQYkVedGMwleRkl4x+X2OScpcRBo0cM++C4AwZrdM
8thQ28lz4yfRhXOkeB+j+sRAVEW9rKCVldkP2vc1vW85ufkw0rKZh1ZgnLq5zfHr
+jeY3XjqTUo5F1btR5Yix6OCZRds09/sBeH0iPI0Tcs2OIqIVuzp+/0EKjHO9ek0
PFH3/1lXz3WVO5CgXX45K3IojhG2sysBy2P+Tu/j/CC586RdNEEtyGF/ckn0UtZz
HFKgi4M3ZFR8c6DgSn1QCofMhuXr4Xn4BJJxJ7rRVJq5CArKrw5DpyoC3wnU57GZ
gsxiYlfUlt6zucMjK8a7LmXQEgh2xIL3ubQ9rFi8JcfKOUP0rZXWwtGvv/jsmG24
OsnAnYtNiZI82P+C/chc+yC4KYOfY9cp8L0Xu4K2v9pTtShO5DmTggmaTgkJYlGs
QIQ0cFVjeur+z1OK3nRDPUp97tjbEY93VsXpGBnxEWOZxyEEdO0EKdUAWzE6PoIp
X9ml6764stUTpIVTG0Xlevw1d8ugBz3UvuEc+OzWAwXz2rpqsigZbfg9qvemx+eb
H7xpwDuAw8rBPBkwQxxVP7icBgVu6quGwUohRsT+qd2EmxXk6/c0bGN0X2qI5i1V
ka0CODjHE3Lv/9LSEoZjgHTg8MNZtBPUxYe65dyKC2kjBGkkkwqD/25pr1IaiNae
TfW/UwjE2viOeU+hadoft2OB3cQjdbKTBHGN1CAP5NikpheWnkanw/6iaRmrDw04
tQL0Rxp2QGB4xABihGSrUnNLXYAEPhgl7W6gZZ4zLpn8B3iNTBF4/8+FdmE5oWI+
47vyaVY0i1g6PzaaDhipLGxUxyDYAldMr/WyBa01QKieHKlaMhzFA1KN0JV4/CDE
INcs12S6B2cn2Md+mk3IfZqwvStjTRsYS2g4MtNJOzVhGgCwakk6HBgfQKwa1Lly
wQUqnrVmMCBVbIDA7opsc5QxmMAWrzinvUZ336eCg62c74ELmC04Z/IZdtbuPNxO
U/FeDBV+3Mho1Mdg5GuaQ723oVkx0sLIcMm9BsTcLdhdA0WM6rKZY9uCnUgxB+Zc
554IJ2xRAh5wAP72g8/srbsb8wU6SjltDT9iMR2eEM5ca485HbakBohTZWxaab5O
ninUAJBEltHhmF8lt9ta5eHXi1vg8mgqwPKutqNDiZT+3fWbY6s4nklnhpEVdYAQ
RZpQdQHAPctiqXvuiJoDf7MOanhK+s44ROqcifZGDjJNKixi+8gmzQ9lHsm8dC+0
cnxKaadEp4pFGprFtIfmDRg6t2JVr8AI7ydfnWTljJOruHyVNmZYSyv/2f10+dKt
pjAVlQzxV6N74B2FK+XvzIoDQqKyfwWpN7bDYrrvn99FNSuwOVu3yKIBcfFyYA/z
TnD09Lpjss8VXqn1WLveOkqDkj5WENlZAHcZvZzODiviXUC/+aJdLOcmRC3EQsMU
VVNUMUN9Uvi+VWtIHm/IskbWg3I9N6q66ZBIqvPteT9SZkzBk5DGb2PdwdDAvJ9k
glW+2foJxAlhDXMkkmbgiQaKnMZvr8vBMjGgiuFeWXGvMRTUswrh0IDvJ6x0Gc7y
j0w8W/tOJU+ZDHacqVgciC0tDzWPzMkp8kU8K/ICWKCY/XWn88XynN05IB3+bZJV
8TrMbfd/upPl0HX8L0gMdtvCgpMlELVLeePTjf/NDBDcoDRXWe5neLTDLE0L2ho/
9dmoZYxWgjuV73jCqqHmsp/sujb0M6OG51m8PnfoM4fPEah+xUHEokf97NTHWbJE
khxeADPsB7KcK1JfZAbsYnXbbEVGd2sGMNhWKzDxerxRwMXdZZ5+sOJ+12rYycXP
nesnRibDErpgP7Vdb+QylIOmnlMSaBKemuNyigM6B/meiau0/kJDIh8cwlugShij
FHsKBBA7I2cP+QJGFcVYdmWORQHDT2M5CTQN8C0n7ZeAN0ehjW+lheJ+26GuYtD9
niZ48S5JBBelDEQveVbkTzexKLIjab4SgrHTZzcvdqOpHIOR1C7X80YHujAXGK2n
/A/PtoylyaLhiElknx0qXUY6S0aoHx8eEYRyqOdnQuLkc6lcajewsegeJLoST2WJ
7X5iKQL4S5+aRXWK94UL8KECLCpcRoN0IxCwhqi3hisIScuPQrrBS/yla7e5m1k6
JdmAv2Y0RMOlfxS9L4KiYNFtblY8m/zcd3HNmVoxJtWFU7+9WHPJ/e3BtJRUWBk2
gce2gmKk7qQRhqij9+m3wluRsUfvA4NS0/8C19y9nfPMIHJVR+2we1Hv24bMIGXj
pV1aoRefzPr2auM2CtwZ+VKaf+oqXis4KWNxVZzoGl4DmlkV8DOjAWgw7zjFS9j9
tuMunrtU8OtNDO2pL9eVKVQ9HNszd+JKLWKRWM4rSvdl+BATMApgaFdwG2QPzUsy
aWq/KhJI6c0gy67DxjqvyJ6Sn5arlrMjgo3u4nMpj8Rb3lcYBlHlD+1/dpSj9HdO
+jv6UOx7FWx9x3XGRXMRNuQIwZePlmJMEXM5CReeZgz1XMWnl7mmcmXR+c2/S510
jO8yW5F0WAiSEDH+4cnoIHE36RmpQRA99n5MArypOSJiwuEh0AhXQ3sOCBIvTyEi
J+vr7P16k2uzpsIaK/YARO0NhCYRDQWr4rabzIqc/8kp/xLf5gjhDiCvBI2imeTq
rG/MXt6vrg1D4q9T3qhHAtTTeXABo22o6syGtDWk5nknOl/8Y4ksqRWEVTFvG2BQ
w/UZX6oj0hJoON1UFCaZy1hUk1MRi1bIQNolxAY8zMMJ/dzfomTy9OpmDfReroLF
9Bc8tkz1f0z5E9A5WS7UTIR2sksulA4ld7b/hn+m7D/5zCSCEyxhXC/WQ0ESZ01I
4VvMYWEcLF+r6Pe1LahjYuyUGcOVgQUfh8bPyT8s/IWeCWI0pxlqZj1up7a0j5A2
Vn+nXlrgKVyMRNt1/2e+QuRNtOYKI7HFPnjFiYscYg4h/VYmPPZ+e/AGnNH7bvaK
+7UISKTg9H/aZaUvYfLkMh4SOIriY38p0k/Y1ojCvNKZVICr91bfIAd7z21xGcmu
hf1N3rAV/sFaB2+mba+zw7Sk4hiqT2KsBBdx6txhcxM3yScwyq9LS2b+oATuULPd
jhNRGODICHf6dm5yiog7/b6GKucHA233IgMP3mHDPTVa6oIWQ0PM48Lnf+QoV0n0
2egBV3Atyx6MqWxJk1TKgnicPB8yWbIf72SgI6l9QK7gwnU2Ds3slH8IpZhCfwcy
lJBmOKiy81rFTDEnZfMupU4gA+PXrzr26dvhJ13svONsxFJOzyP/bNBqg5Fgw4rN
XxjvAFgy2qYoT2nKkW5DQymwa0YpYen/w8lt2dYcxIpox/qR+KF5cEgk98Kd/FoN
JTDXZQ1riFsu9ftHI5/v7HJ/LDKE9/kYCXQpD02loYOKbnvj5ND/HIylhumLLrw4
gat4PWlJ1WElvS8sj3fbUERUdvlIkOwpNYTS28A71MlFfwZIMb1bmVZXtZID/mvI
riEfaMc5wXBeszYPVBedIicAHwvVWHvEJXpgJ1d/MpdDvf+p7fEQFFGgzOVQx375
7SGPpg5JDYOOx+JVB5M2ddabqgIVdI2F+8CSqO4gq/46y4VA2sTK7eLwcV6cOSo/
v6F5EEqUBtxmWn0XpLNqfjNmTEAdfGCkGWFnebhgmuV4BfaIqmYkJV4orhWgwM5S
MWwZFBVd4yIOSsiqoPst6D2IMjYYoRtajj9kkxs+dYSlCd5nOVDIa55nBaLw8QHI
yyHSi0DUvNw5bou5UJHktBP6P7yOvlzfjyxS8w/cwKZTZv2YeO5qJI9G99TUxtC/
X7r2mrOtC1BzvG9QocbKFfj1wt22nPLXA7rC/hPOLN8TyOKLvRnHIYNyeV1abQ8B
DqsFab290yfFj8fc24TFv93+BXVOgGZdq+he5nv5+mLF9K+Wmrb3r0vx9+ISBvGH
qlb1OQi1MHWgtOHYFW/5hyEDj0rlGD+MBeWH1OMoQQgf9Fm9f0bPept4E8nm2ADo
biw8pb41owLj3BTZouzYlTfDmSCTRsfM+Gbm4rzdz8o/Vq3Z151cMHTst1NifjqG
+Ha7iz5tkqSlkeO4bTxoa+iR7EoqE0q+ITDHBSvzwZPanMd4WUVRL7KEcoB+psz/
WpAV8PuNi2mRPiB9T0/z3h+GfjPjvUDlMhqMjMstRKrUOagimPrWjJLRL6tyhbBS
Tzd9Ba8u/ghIQ/qhX3VC6deYAQFVkl6WOeQacZaHCX76+3MfFgqxvxPgF4XQ5lQg
kCKbTAM/c4DI7EG1RDmlBlLfEuDzLuYNithQZ3pfeQGNzo+c/M2sGmr7zRcCjDEO
7R1YUrkxg+S+pGcZXVZja+mawKuo+RhYpo+DFHG/5zAjleORdjlvdJiiyxVeAYRG
PPzxCPxJtMk2q/RfEUlNHxRmOVWZUu8WwGgWCRDgI7o5VSKz1CkDGYc82gCDcWzP
kMSsiyli4PnkTjnreiASWKTQZ8fR4EzWtUWcaUfEeqvBdHoxKxhBgZSInSi/SC35
922zY+xhryzNyLK7k0iby7GzOadTPCri/Nv+vqusDBDcEwONkjYc6QIVWsixPQ8f
o6y9P/gTc0IG/Gg0pBOf0Mrm01V3uChCX4nEFa2603Vh8sYeUTKg0Xm3C+bTEXJ4
4wovPoWrd3sFhl8XOmTHnEp298fHns9Wl6+Mh2vNfV695WHNPY7KaH6oGRIV4ZtJ
wvocTtGWqD7WW/gQS4tqVEgqH5DNGaWWE1c8QO2XF46pHBVPdroifoHoiZSFt8YV
EndmvckoNaTV34iraexkBnP8uW37Lfd574Labk4FZbwkVImQ5WA62L1GS2g6RlC2
Pz95i6FOFWcxZpiFNsOsyK7NeptBgRGNKnMGUxqtWHTDMIkEEcwuuObK2xpOh+3h
704izd56U06hUbXV4IZdfiHASXtKC+RDljy7xkLWHNFzmX9gQpmZ7sIARnFzRdzn
NMmFDJGJN9P0L6p15O+xACIRNHg30fCeDbJRh2Gvs0XeA3tTcWv5rHH1C/Gq3mXo
HCrO6ZUeaZLneAbp/XPsrOeGTlK4CqN19EAl0d/TKTcpuYD40N9h2bNXf2BunpWg
mHA5V+d1eZFPOsYn9nIYuXi48YCCMltLIy6TlKut60tUcIPmYK/ADrkZbzLJyN1A
WAxdVG6l/Llqz9MM9tPWCN2MBNU77fcz4lhCxu8/ywvI9ic1XyqDxa/hNr7XNmhu
mUmxx/XS74COVEqq7n3qrGW+v4TW0AGEJ3WU7BgvmuxojQN2uDp5Jvq5ILWmPMbf
3rSfkQ9BT2HuTAZdDIF4ezdn2kTEhSP54E8d64OS4KYQfdPChh9XdRaHcpfRF01o
Ps39orjrmSOeXgbBIKRokSl0fYeej9JBxXHWDpdzxQvUp+AKoEFxhTZPQzBJM1+1
y2LNbq/tRn/CiVh7tqnjLtyK+MVKPZU+WbzsA7Xo5Ml7dqvZveYm0YlRCtbj5Uvs
bvGiWQKLN1CZGbZLmD7Kb0kF//8Doo5rpIXM7w2lgQOhQXrvDG20TpW/Xy2qvfh0
KeJqnS9ZBPc0kc2/wduypAKg8YM3cyJ0IAkWCKzGlgfhuuc2YesPP083WUNB+2Qk
GSgHOvUnG13wXFR+FXHn9M4da8QzLYnIJP/Y8YFtY8c5HbKLkPP513LFUW+d1h/E
tZtdSlVy32r38QXlSFvz4qhA53SaBrC2thXV79gBjykDxPyFABekp/CiqPA20GwX
W0w4IolBRyEVpwRgOYyzuxkC90sumDZ6XPu53t2iJ5xZw+uXGV2lCyltpezykyWN
UU1cVzo828xAY7DPSbNX2eBs8OSdOAeaFXk3Cvur0omVlqcgi0xJ4I89bsU6xYJA
cno20e4e+sDH+uUsCvT3zZ9z/aVv2kNkjU60DCBD5l8uhad5ZeKr4G4XDix+M+NH
ecqzhfUJAF3KxgVKiYNrtImJpDDIppxp5+GdnuK3XGAITV0UPnZy2VH46H8FstW+
tTgwleYyg/6FSU8dIMrIKXxWvGRKd5NcwKsa8xqYa3LNf0zIXrHQS3r9rePIboq5
Dnf83R4klnRAsVuN8TnATlqZfgSN83leDDp8sfWWPN4NyPfZL9GnlZWCj9YVbG4K
QiibwBDWFt8LjO6AihzWWS3BTw8NBhLp0YFxRH+YcpVRbJMEkpxU3LPLBQNcQgOJ
yUd9rSDFoq/EWvbcW9U/pnCGeA7xdIiRYCrOTV6t/jWVqJo6LHEkzD18zIwr2Q0w
v8oIUEgbZ2ZhIs7HgnO8TCgOYAdgxQtS8FcsujrP6dtdeBN6ap+7zlOZzQLfXRcN
L8UtZNJ6j03cDjzFOssFlqrx5SEhjuXb0pvr4x0sUnGRspNnY4mI3OOodzz5gvkC
INeIcimsYTY05ub7wRyEp6JTOncXx/3nXS0TFbyhg3Tzm2Qg0P2pqSRphdYM9TRk
Y9BxAdZc87z+BCJiiuISd+pVlleK4KogFQIV0ENQqiQKwOdhNG6bULVxxiPaF0qS
566e/hlmam3bxvjcszB/Ez89lFL795KMDiprP6sodx1UIY2fPu4qP7lZzfzArfOY
5zq6fynZ9Vvtlmg/UIslbnlmZEfbNK4WGL3el7Z3J1OhVCP9AqkyCcmYU7kjC8Ii
`pragma protect end_protected
