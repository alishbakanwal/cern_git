// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 13:57:49 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Dvdq1tiSEiKLw2AR/waUeyIK33Scs2ED6WXG1rW4XXdJjyrmUVGhX43u+saqUZoR
yRd+Xk4vMQuhpdBk45/sliKn+lI8K8aDIt9DiL4lvRCFMaJVXSSaMR7l89zy9Dgr
UE7EHE++ExFKckAxmbDBo0WGYNxKjX7glcn2aD+YIqU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9840)
xNdL2DBmD7rVsraQJgVNbUOFyOQRckJLUW5zNRfc9O3tAahxjox3fzWUZ/Yokwys
QKdRErA8zmj8YXWv0TQmc2uGIHouFlyhbUI5jw56L9DBPXqY1nlxKPbTMmN0Oaod
f2aTj9Krjru/oIfQ4/0FYhr4wWICUC5HKWlQmGu7cAoGagBUQg6ugZNfiJ+jD4kA
gaDHRbVhZS1QD1lwUyL5y7HO8zrECqe69J1/JS7NacxAbBIKT+DPYgtedpt6pAxd
rnC+qEhFaCcYQiDxVAxUCZRDWI1g8fd3rz46WnV4vBd/V56tskiWzApTASNayPoB
eVUt7ZTWHh5SsPy/KgTd+yMO0WWk7W9if4IReMHioxCsgaJsEhzGuoVrFdXUzwt5
7q+khb7WPnRqw1hpeYZpwcBnu6Iuz2j/eYtaJHk4ukDck98FTjOskHtE0LF5iCx7
gUljuP2LCSWevNXKIPlEQ2J8Hu33TUoTXZIbC7dUKKWIqLS+xmssFm7t3WqkjChU
dKdQDVI3PfAThdshM+DL7T/4sInQOswwGJb+qM/chwprdf9Hp1o/e0p4Yb3q/bvi
dqD4KwowidkjBAZqT7MuiAi44O6W0LKvc9jroYx/riAokZMSh2X3uEeY40e1psjf
heGBxbPGdZtzCjAxCLYreFYZXCSS9zaP2p6z5eAfxRcNKgLxwPJSNtzNEzkleBgU
tr92JwiHHc6RxahAfYyOcCU9ltaU8J605OI1TNJGlX9IjXGH0RIvc2d4wVTMZnLX
4yb3jxKaQxXPCakOKOupq1jik0YK/SbU2c+quJ14WfOQCWc3/9hvHsGMrzEyIpfx
bLpEqzpZUKzfuxSQAnNVwS87+8Einq96rJoKCH8+kU1SA6XQir9WsWkko38wbcoh
hBWNMjqJaclg30TyIHQgo2Rf9mzbNVrVuqOkhBm2aJhLBhNngqIabqV/OW6wz+BI
hYA4gK6amDJqE5rJKthiBjsuDGhvWx/JNeV/r770D4O4alV+I0lWtwVPgFrPDHjA
lk3RHfD892uAZu8fCv6Cf/F3XSB2VKHkOG9zqC6zQyCCN1S3NpDXx72CynT+/+DK
sqtnzpX+oXTcv2I9MQJbvBmrm1vVwda6V67VGGncvNRcawaVPgwnc7VL3LB35ikb
WvH/QetINdaksAaryVNSdf41xNYQaoY6QxgmjYzhWBne7lz2Iyd1RNDzLaq3wZf2
yKYhiqhTCTL1U8/Q5n3pQIXDunZZ50oXNwW2vkTEzIAlya+MEQntO8lWJyv2aU/W
w0XTGHfK4L9K7UFuA2MboYk8XIXcZ753GNIQA9OHwqL+0EAof1f+juEYdlLEEHHd
33l99zaJR3b+kcAKGULbqQR77BGhrDWLIpn84M28DaLmQnhX7b9wHJd2GPGwZde9
eZsjvxqT7MQBBPnLZtP4oaWJbAbDv85XHdxl0bS/bAlK7vCWUQ9+QpUCB7RMbTNP
84cFb205eGzp14H+6uvjdQmbVIF742sZSajlNR+9bN9DImZktGQ3sPNWu0VG3CBj
8HJGPQ+8eqZ8XKXzuL5+cqdzGa8rT3CZTw5j9L/O5U/k7fegMUaln21kVHigIxs2
u/jfg43he50Y9tpwsJkUeKKIihQWz/TTs2dCy0rdgLcPcDAHOpj8uCK24gmGPR7d
ul3VeFsz92F+FvmaaXK3exoQrBEU7dv++s2kUvSsOqyqdPmtGJC8wx73s1TT/T5z
BqqCkg1385BLU+sd3hNyLnEx+7LsHAatcENUwWLcuxAW+tmrG0Z6CFRMFrRtPEYB
5nuxBmMIR3j8j/MQ20ekf5KcYEwDitE7o9Ue4NsVtSbHvuRqybBFvxfjItLzKG1C
PvEpLCfBbD9eU75uVMHlwFeNCo9x2XSALp/C8hJrf4XE20XzIp7NsyMopCEOcfp6
QM0ivvyBx+yUn9ZIeJlb0ofkwV9ipwipjGILEX4lAdvGca8KNI+rwxh83OpGv8ZS
8SlQqCgF8wfCxNaWZpugajzlgcBr92s/ghP9DOa9dyW6aZnI9+VsY1Ttav4iA137
9pyo5K1EA3CjV/ClfSAQOZ2EA7xXfxsLSg3O7ByEgRf4gKY80aXkBAHWaW4+lRM+
TONkH+n0eGWe4NUpCcmIbwIUd2TWoxpfcjukwP9icBxQNfKp6FwYtX7h5fv4oVa8
j4Gf7yvegdQQsHQ9PemR6YslVPfzYgSn1UUoI3H3upRFbH6pO2svn6DyNjxiaaAC
LzeWi39xNJB4d185O7Bc0xjMXJEj37AeRbYrWXd820o4kr9SHxiDFXS5+fadBGVg
r7w6aAIGRYhpWTNGJBCeBJgyk47J8NML1DSBqS11WpSIsABTo1tV4VwgwgMsoj61
aEUteLb2EdEx1uLV8O6WC7JlG7rpxMR/ZkHm9uhmiIUSn/xW/EbnxwppLwbUva1N
115uiLFj0bvBQVPr6Osz4gke7tn2wI+2S8+UT7SDYi4aaKiF2Rt5WnLFA9V9XV49
R09oCtTTcfUI4i5/wlqHQ6eXXERPeZUit7zlM+g9/6vBdgsUqeWaL1x3neLRUUPh
Z7hlgOb79wnSsgzIFxoKF60XxUzpoIbZ/gA/kshwJq48nVKP7iLtOUCsfjAg3dzD
jqKvs8vpd8nlMbMsl+VS1FoKZFYqx2EmZ1MoN6dEM2yiU8lE42p13TD14+N1vt3Q
zzZS65LRHPhG/RiNc6gvN1h1UE0+emk5s/efS8+zsEgAKhJjfms61ByooG8dcxXf
u2jpZfs3cBN0Wcu2ZKYg4cHRT7rMdvMnzKCr+N6hUP68PMiIG/AJ8LjLxf16kpNV
7INdAt5YIQyAdQr7Z4YpFaNUsIMxYD1KiW2gBPExy+cFiJ8a6W18cb4tE4l5Tt7j
UaeLFVBYgteSxSs4wjQSKzT4fHKf4b2bXexmX9Ys4dPjHeUbxYlGuuKN05cGfSXP
KIoKd4b/oJjHLOWHKuqVamnyKUVS6ce1oheKHIZF5TIjYPL2wpN6R4c+vZ/vWQig
M8CK2dQusk62hWWAtbNdh2wEv/la4PX0l2EK8L3c+8cb+joaBRjUsU0+PbUPK4ky
1A5emdlE5yz2VlnaCbNlWXT38dwkZ/k1nzFgX1pw4G2E6YMYWhv8O9wSftCywHUM
zQNBbM48HupDB11GnH1BGFMRahAtQT6Mi9r1t+ZY7e5w6rAesFpsdHXJGC+9S/HS
X9UO7gX627eRUQLX+d1SnBaLXGdPc/ssNVUUnp+zs/k17xub0LXsGZiinNdKNOpo
6u2HnFqGYyoxA9Qz/w8WAkDrSgobVv2+uQJr63mCZCBh/DBPtHkV0jXmn2R9X9kt
AeAap/ffo+gNHKhM/CMNDS73nxpHZDJQ3tdfDepxFzfcrTo8OOjrZ1hgN2XqRJKS
2OVJs+qpET5C/03M3CerBiGAnyaAMtSfRqsyzLGZf5TDPBBT3Dp6I83Bt/lEkFXs
bmWmIfw3KV+Adhf7J9ICT0s6yPUbyKsO9h6eaDQt64dWQsq36KL8vjJvM5tTctl3
NHZQqniaUqGwxFmhHsQ5pbnaGtVS+A0Vdf0tfSVt9196loefLu8egB7xwKa3PH5R
Gc3Ate2GR7arDFjsHMRNLgoMkcuU+TLtPi3q8E6WTsFPbNo4301WhJpWyaZvkIxK
Ntjuea99VvAx4zdplKi/wTAIZgN84QuXX4FuSNl82LxIkN5f+Il+gr3ivfYnZ7p5
uMZrXIelPNWqJjKAmHg/CFuspFKyIh38IxDNXsGZ6P8mSafS/rBH0CzPRc33ysM/
QV6R6STY8Yh5bHUcV8K9CgU4gseLrUeczdsMynCjSDr7b1B/LmTOIt4OWO/ULkwA
TX3Q+fuLQyRSVFlH8kC4DGSp0O6IzMu/3fTFG8IJ3BUq9SxDB2nvvOCC5vnKzx7W
2POayHP02cyCuuj2FFVthuBvzeLhSUdIwQBrMXLhp0XcASKE3TMkuGDKbeSHWgWZ
DVTxykFOQIynFTKQAh/XLI2l0QatX6xjVltbXaq3TDAoebHKVnCq3dQvybyaVyZ0
b7GLYDSYkb6mwrpj0P8XdMf4I/YYnXKbiFzMJfCK/ZPrlIH5Cn3EO9tnPrr+KoiS
TK+rUHZJFBTn/3p1Rw+BPgSu7UOfuTA3Zb6AMPYR59Hmm3fnTVB3VH4o8lrUtLFS
xDN/aVqqgFiAvZfJNznBfR3YKgkq/BzptcFpRSVVdW+NYGsLc5qBxibW13jr/pwD
kPq4EdrF0PjzJIl8Y4Uv4OKo2s3pSl4xzFORyO0M8ulunr9HjIFF2lj0BbDpns+9
P5JabelwAncccwlXjdQLb5kkzgiA9wUzcB1mbWKeoKzkQf5k+S774+45K0w16VIV
0B9zgnE3udEGuzTnUv49y9JuP7VABPO6wiN0uL6GWxc9hYBad7s+xzyJFNt1pso3
gNLLzzq/iedQmkRCzoJDI2/2gAxRIH+dx6s6hOurBvOKtAU1vs9qqgr1AOUd5mea
Qh8Bl+8/HeOQz6cIqNqyj/7XjdFeOqlJXUjWn9j9oGkKvILFPnODSfC9WZSXPs+Q
WZaOB2pXEfa2ibaMszPTT3X4dHo7Lwy4hVaWnLro6nkN1muw78NUm8DFQWr1EwfI
3cTx8N+pnFEvovIIse3K/TMAkGOdFT0o9SIUTNi9mrjqwrbfo3tD2w9uBvRO2mMS
r3q7VoPwWKex4spxzNaFJBPFjATlCdZP8UmLjevIQNatC7UC77Ne0CqtR1hNWu/E
Ea2nRikdetjYwbMO04RYEGZRZtaQfETYKYzjbLRO5R2Kiyu6FIB/jfyBMzWjN1Da
1PU61iLzAs8EsIun7FwZyXZrEo2DWR5j7b1EF8wLBw4amWRgQTcW6yePEdyxGNh+
yfE8SUFvDOztl5CwQk65z1uG0cIbiCNh9OfwO+vUvg5JbvNkhHy8RHD1qk/KvGbr
LwAjPV2QTjLMgpcakTcdaiIJ2tyQoCd6c2ENqlgtEwNdRQZpClaWTWi56DM7pUOk
YAf9o+hA0SLPaz/TGTc+brAGdV3kUpMJyF6h5YdY+BAUrVbGgjf7sszYG1W0ZvRg
yUhigtaXczzpiXE7lH9BKlyhdlegSkCkP9v995RgzPmWnY3YsBKMSBSlfAzkLyWp
UJ2BltIkBJEFAFnY3eXZMiUTCp9NG0ttolfwCB5/Y5xorJxjQ87kAgyzbn3KeDiD
Sgf/OjPgg9rMSUbyR/4zY0iS6laAMJkysBJpoMMot4gX+G5L2Vxwy07qTT36cW5B
tkjwzjz9Qkrn5YTQel+dqoEZaBLL0z1X4D3G42UNvCbH3uYe1g8MOk2yX2VB0Xge
zD5rkM8YxKCmKPFLTgTsTioqvdmi1g2FqDxCq/QVQ+gsmSeAMzkvgRhR0bC4v/l4
7H0gGDwyy6hxDO7I9KeW1G2ocB1xpIvxMER12zznRly99DtxwqLu39kvIqGYjyVi
1jylJszZQjfKLq43sfva4U0cZ9o8gzswho9LpUMb12XeH80aujevM1pIDjUDvZ5e
RKGQjwimY6+ygoJ4lX2k8BiGzjeAxctr7+Tq9YGamTmjl2nNyyM6VyHG6kNrtaXu
Oro/mAOJo5aSOt1EMA4ryCYvsQraimQdTwPldOLaT+Foh4l0NhzcKlRpAyRVr8B8
PCg5Brh9xrdUYzAWGMx5Rr7EYFRe2SuxEhQSAzmk2pz8IFKn0hF7MzOjjRFMxjUj
K5/S1EFBht0VIoA039qcfQU1EFsy8f5Ma2I4x/ypUzXFJYtaYyuF1BEZECPYNfIb
6IX0eAW4vPBdmhGKtC7VqchJTturAMo0bAbv2NdDyqVptnmX6YyQClqbBkwMxWQ8
Wa9ltxVDKTrhznPXkWnww9LW+gI0exuVAyrtN5FkXxjTnq9hZHSJAvHFDuATTpFJ
/E18j3lRRlYH1EfMOCqoTas+fpzYPmGTlCduhhcdsi1s+hEudX0NA3ufiuGWZb8q
BkgFY/gIlJDgp9zDlTCgV0IVTJ3GjX99OS9i09SNgMToVPkb+pDUSJcypOdfO4qL
TCocX4/94tmJ1ae1KILZZRLyjeHZ9IzXOs5HtdNAq+ppGiPvJ5ay/NwFJg2voyDk
4Cu2vtbFIbwDG04UZ4s2psrZ0wHbPZqZUBMZogJeeZmtN1OaxebsgmMYdp9J0ifS
0FoGLNKtM3wTurK37qHjjIzedpuK9WGi8gHfwnJuNxccWE0eq55o0fj6pK3vHHak
VN5bzBLSunmcTv1pruAL12S0fImCtEVJSvZbPEIOu56bbFDME3PWJZ8ERgASRmBE
W7cBfrW4MIRob65DBuKx/uAzgAcR2zFLia6z79asZvQLb8CIZotMyuD0S3rauyYV
I9RXPgecWn2Cp2cHZP5K630gtvGTZRmk8WStHLQetIFFIZbmq8kFXv07QV6JK174
aMSHDZBpJs0xUWcLHrE/OvYUJKkVzqXFQFnLuRGgN3bQ3/Br3Oh8CuzN3QFtPjX+
xYHtaTmzUi+YOoWWCggA1Nyb73DSHopZ0RCKz58cCBi3WBlUHRMrs1BgHZgLL5vD
0pT8az+a+e+8oRiCt8t5VacdIdfSohR+AO1/3lPryUh9HL7ps4aigKUXdtp7/OyQ
KOg8IxXftkC31FboNTbbmC9RPjekm56zExdO/uvDVq5UTD+b5PHBAi7XzQDL9x4T
42bfZdAgYmqip/wdFe4CvlcZbtAOMdTtSpGTcGq+qsIgeo+XuPY+xMfRBCCcxvNZ
dxyANwO9kVKTVpyP3wOnc1I4s0nuF4CjrMTUJVjR2NFBK3cUczMGFGPMEkLVOzCA
YDIQmXo00oeEXbhVQ8WErflSu6bgpxyrLyJ8jHQarflvCXM8FRTERWjm/1KwnhBc
xOgYf1n7GIbGJQPv0PyHIUhfvJ8NAM0Auut7sz2iIn89ntnFg66l5xMk5GrwGmxH
kjWLyJljHLclZq7Tdihs7xUfBQAfs4LNR0Q6BXoLOAw3/LrXMKYpQtjdorhERomL
HIGI889OB2HDgmBcy+guNev/voJs0Xibs+yPqO16scn//URi/CU9kxTh8D75LXOz
n+RFReTDaCprNF01Es9bKgzgIY//hxySAMVekRsXPTkb1b09Z+VOGGTtNWxZrqF6
6gwkbWcQBhCemCVtwbgvzAnU0TWTHdRyuvMoJMNNAcvlChJaZk7wdoh1mGbJx6fm
40JC0TR9K8Lm8geFjwRtsNnIGLb4wdOatWzRDExcQ+9F6QNxlqefzoIliBXGens2
pgZK6O/8WiqcpHQPWzE3QSxH7PgwPARbG0IzZ9EH1D61Ch+Fb+NxVp8HOJheEsbR
ZP8Mvhf+p69gHzmNBoHxeQK5289j9d10tmNQiRdVumE1qGIWd2e2XXpf7xIWCeUG
COpABdZduIU9izrfmvwT6alVY2xfg2v8unTLg5VnQqcDji8vsjWNZ9Qir7nlcYti
11GiqMBG4N8FmPu65q/Y15HlxKZQ3yBlgO4U9b5gvgMuKfqM76lpXVFBBIZC9teB
x9BoONVHtSkQk89iRLC2kchSToVqZhYjgWmCF7TQIJpBhO7WnQjZUydffGuGPHmN
G+ZvaMtE+FK5IpkgYwY++6nrPGUxxQg9scv/KuC3YbHpGg4Mqv8AAhx3HlGwv2gV
31Pgl0cR46GoM5O+6GWbIUVirQLOmDqgHXiV+YqLQvEqOzwHHEbB96tvvpbEo0OL
2A6LilHEZsDFL8l65CQVm6YEuqB3/5yRjDiEOKRh7ftauSGrjQ5JFhGNnvmVLpEO
w7YHph2OFNmJbHaajgX440xychrBcoLDAn7uBwCp2kifVhrTUIcGR1lPCaftsAD8
uvFyodlg6ev/wwq9onnW7FC9EvV3YURRLBIb5ilc/VB0vvKhJyBox9TpARRms4oY
0E1qD+wxMIkZI0BOy6z243U7c2y4wEj2iqDd0LNor2+5G5eExaZMTB65nuJINZpv
+JI1uXhYk4hzkI9E8drnz+iVwrJA8II3eYvNUmyc6fDJXQXhXfbwXwodwa8Yovcw
5VAbcwiJ3prhH8iGlcIil0IIh3j74htdRnICKnZIaO0psotJKQqFGYJiYl/Q9h1M
0TgAnfyiJtCWTRlwIiuP33IzN4gyCe8znrW9o5kxbdz0951tCfq+uz99HejSfQee
hSf1eqrNL7MDU0SEnkLmmiDo8tjS92fHpi7L++1zmGa1vhdPGSYBan9pVrWVLPte
zlHe4ivtfm/HJJBeRI2yOIXfQltiVw5PMOpvq4M/VOvIwZM+4W9V4uAOsBoR7DTG
7PFJMuSIenBOylM/oCxYORANZnUcenVYjn/O6UqV7jUfbvUxhypqO1eZciA8+Wl5
QjhycDSuyOsi+hjodhk5uIpx/FdbbSF3Bd8HGnE+jbPOcZ8MzYpNR9iE7aaX+xag
SAETICqgJGWCu120D+WFB0sg+NzbByy91lqnQkqE4Zm/9nKPUYHGSE4OMdDpYD9K
aB267vH3yneNG9FsK0XVaJUdkrpsf53mC8FgpVaCfnZm7B4XDQ8ekIXzhEi6vj/8
BelpTMgzV+kSyA7yLrGmy8pemwK5U3CjJvMke8ui1mHK7b5zkhv+O4jI6ecnHlGa
t0pJGtLz12PPURWiHxS3Bf4XM+tk9hfZ0FfNtbD+1EjSsx4H5zxCAP44CR8cw+ju
6tKcXFDT7cW4IJCGADewLKmFjQMqKcSoX0g5h6nrpta/O4YOtwgic59Wya6BUCt3
tw2YORaiQtLrpWPhE0dbOk2EZJqckrbuRyh7s90VuVLFnH3cBcM9kMLL7VEvhjWB
7Jz2nAuIT8FQzLIZFGjjq/SSK7oy7oV28PU9F1fw2fm/+CimkDz3VAJwsptH8/QV
oLwv+ez0ZCq8TJnEnQCxYtQYgZrLE4XOxk0d1PLKrkdYd+AePy3a3scyHJUAmu3C
+uWF6Yq3md0W3VF2g+3sUay7S8/A0Ivu609+7AjzymQ9qW67Mq2WJKHCy1GIjKKq
NJjLbh46Dr5Gt2k8JCp7USnhb8OMHNYlaTBSRtYA3gc1Mm0MU9PDD1g6+Y6/Bv7X
I06iYGapIp2WKSdHQboStVy3Qpbrt0CDSmVq/tCCNEKIVToR38P/0hFuvl0pXBV5
St442I5S8JFlBBa/qLhk+0XsbkT4lQ079+kMKDiT1265g+TGobxCPy2oSz7d7Wjl
LQKlbgFRN0Z7Xt6+/vlRcY+ArS7jVXfcdcniywpr38dxxXAUpGippXTsBVcxH+WI
wxAf2KhRcEyDiCKtHYi204PjABYaRgDQN/g6Zw+HMXCYw3Oxb/Hp1iXiNyQxVs1X
c3SwYUolEQCCiKsYKVESoRgz7NDK+Oqd2/Q6qn8g5UB0NcPk+F4CnDsV/ktsoMXF
C3rU0QX2KhljJ7QB5xGOf4OU0Gi1jgVT+PCkrJKms4/zLZB9wNuwQO30peJSOdxQ
bDLo1Y/o0wlKR2VoK10hxK0P/AdNkvX8lbs/CeSOBfUn/SfdV1SlIGVwlcuyW10b
e009RUW2+w6Uvb8cdKz+7oS2EpdXifNGnK/730X+fuTf/AOzRiTMbJ7PxUKcvpN6
3RYlavgNnFNPWvqOV7xuI4NBI6qrjE5N+YTZikCsOC4poiQRcJLw3W+TuEBYORJ9
DgVH+OpjbqrpVpeKyXEtTA87smn8pQO5VO9+SuvCkj04T4IYx31Xw6TlFiCTvd+R
nIO/9QfcUf/31tCxhCxt32P5guwwy042Fuy4jJSw8QHymD+FkAWl7L+FUmQ/jO9o
yDcKEs9CoY1QO3Z51Tn6LK0z2CHJ6fr6nbnVgTjNCD7AFxhYb1Novp+jOBAcKmRT
LlOW10cMd0fQIJFEvCwAWlMZCRcpJzwXbxBdyBtLTZnvboWRlwStLLpCjgfM9fra
AlfjKLSDweuxi09jJi1BInibRWQMhEWPMbAU8OYALZljuQnz7I9s9LPCclHdt6fc
mSj4R3e97qbKG+QW3Kwyj6mbR5/v8mxXeDxipIWvkkjQFD6pmUFKfhk5g0ojWL9Y
NxTm9TZcl3rcdEC+6bIuGKQf1smX2Evfken9kHvn8CsX3BUkKUMnERA0qRiiczon
2dppZmBQ9hULxm4GV/Iz+dugl2znkjZjY5LSOs/6G2ToPt9tXc2d23b08uJedZLT
kzspKZy0rnoF0R9NiAwmm4dS+ywVwwaCTElGe0o9s9t7BGJRaH26IoB5ykcKy5D/
SDn3a55nuPRurB82MaPTLeETS7C/W0LfRFbnE2JJkgzSoLhb2UuK7Uq3a+tRrbI1
+Xlpgp55pw8+rp/dar5WEqxJGfOiu1FPK6RviLrWMRD2WL5HaQYpoKukNdNbKQfk
763jBKk4ihVwu2hVr7MEzVGEwlxd0lC2F3ymmf4Tca2RJejjZChMsXsHz2LZTTvc
7bsvbAh749m1ngOO1eNVqg67ZE2StUee4X9wi1ybfuPyhLbkdh1hPFe7cW/NGihL
d+G0MuAf7BiIcnI6dNZrvByZJbiBpkMt5+FLzQS1eo1yRycSowAZhd17+2Fv+MZJ
DagXNZ+aSgbKnkOIJ59Lait2jTidkVypqWTqYnIldqgXnuTS6EBd7TYB8blXmLah
XCqN1rdCe+3fRMl89E6Eo9y0xmtYr2d7F44ftHdZ6GdLmEP3Py35lqWif4m1MgOe
040aP5uF/buoXiTFFutwdMdhX2ljlhtG0ht5nQ46abiy1X/V1iLxZ45Rezys/BMx
x2q0ghmiatkts1vp2Paqhz2NlQeqcWLCEq/EK3n7ExVKrQkqkH3AtwNHuFvZeVIz
FC4NlN83N73AKcWKxkVFb2tbKm/xVxNhqtjNM8GJsPtUsUOg1TT/wpTjw9g49rG3
E0pEOwstGylaUFBZhoMaRur4nc8u0a5paG0N7Uisjo7kvcv54i31oBOUUgfsxUz7
5cf7JR7lUVLNTgrJ0O/6xzFLuL5OV/LsP2i5M1IhiY/NfkJz1M+DO6QMNgPjKmbU
oJdWrDvTk7eIDerAb/fVb49f2J1FmRDaosrmspWTtnx1cF0OLDGjxz+enGfk/ObC
3GbU58NGTVJ3Dxf2UjMsNoJoFKo+kuTF9FsTwVe4y27rU86Mp2VrJDNwkIyjF/jw
7kfocVmdMFjt1ykxEm9YrAn4TLWqbCkBbc8bO6In6iIdX+ulP1JNVbpBvM2xoWK/
ODF/A1z2cvvsWdfNnqB3npielxJWbrEy8Od2v8KUllXmh3iCbnMiEb7Ledr3dr46
E8JhusfoNJRv3agt7jAF+EYkJVtq6iE/7yTH9THUdjOfch6uDcZRfLjlIzIiR6G2
XBwcukjWuvNjfNnhcABky1drKSG4qtTDvShpJyv+vOabURDzPeSTJNEvbddMBtEx
uufZp3ko7Db6kF9r5pfPPLhTLYRiF7YsQapsdyCotUQVAt/RdVCx7ZHx+IQ914Fj
CPdcIDBaqahyZZxlM0+ZEutWmiKBP+c7oESKMaN1IXTueZZskqordYvaLCLDS2PF
oU6dZkV7Cn4FKt138QBg2AifNabhHOlN/M/Len+UeePzbRZtJnoTjcX6wdciXzb4
Kss8diMu+itruHHT3IChCdMVVVEDwuYnp3d5hqh56xDZN5xdNXyUC8r9Pyc2pot2
aYvgLQ6zaoz7k4xuOiUSczeqRroij7x/eLlDfr/44O0lK4sp3jKLFskyKuJA4gbB
O6bkSEq4mqgbzTmIfNVTXeQc75YWlM3t5mo+mTpnqrMZv3+9DRqAXqoYPOpolq25
bFkExHW9xvsSPZfXVr1407fJqPEVPeU38vK4lNzq9ZiEmbEeFVmQ01p1PwNPaNbG
9lfBTH/wHmitCYV2Xqno8B4k0P5EjjWe7+6x3RpsYvb33W3mxWbJnTG8URIq6NlL
sr1+XQiSya6FRlVkYkVkS6lWwjTVTJIYp6S06XLXW44AqBQ+1qh/9hcG8EJidSPy
WobgkZesSiOU5BVpa/qTWy61qnNhFXLPmmsB0Cv0ZKBIY+FPAINOWf4L4YlICkbr
4TdLck6yFLTC+BKpSdTlbxpjCRgtRTXAPEJmSTVE564TZHBDuEWBMT6RC1Y3KHGt
vpLHVMJCovIR21sP1aUd6S7PU5qBtRTtn6XJwwdtthhAbKg1abiFtBCn4MqVEP6T
2NKidT2Yh+ng7OOc5Mb3A8X0bqqFd2XZ6zlGkaclnitIG92/YxW9mgBLiyFV+kcc
k8o5KICk8u2TRi1XNRmHWvW4zFytmIj207nzwFhsw/uKfF5FpolEXOMwJwG5YMQP
ZySuAjF4aPWieeyP1TBAlwllJgS/xiglG1FH0oCncfgdjkoUDO4uFc+OUS9kB6qh
TGAdz88TlQwbNPRsX4bkzBtMTGYrtwDnbo8LZpfUqYHzTMcKdtTXvBASu8YhS5to
tilp0GyJvHuL7kI7pe3LvPhjlekgcJimen5kfgqp45CPtzDDntCg36QuTblgIgmP
mDnHislnoGwh0X6hUCocNei3Fbb8SpMoheVQy6AbDR12l6/DikPkw0MXkH3cDXJB
KQLZrYUtUmLU48dXblJxfVq6b4HTlMKn+gMggUu3dsDKg2RL6i8dbyUD1N/rsGFd
ap0Iv7YESrijmFVuyIfU0niUuLNgXiEDma2nM/l+WWMbFYo/fKqA0gnE4+zGsbrS
g9lEWa7MVwuhP0QkrwXNnu+8Lw+tNVrvuyNP7FyreF/5iU+9mmLjvim9OF/CB+M5
RnlgQQWc1Uq3vnIgjFvwG9dRIwqjyXMzk6hbx1+e/Y8prJ528lY4z6DyZneJCF1B
yc4FNwSu29wwjtzJw8tylbZywOl2EQ66XP0sZWzc0LUcNq3VSJ7lw+K+1LRNFiFK
EYT+MUrMzXNe/1KBHvb0YTkK8TVZVzwSlQZc3JTVrRbzbsnT9cdvOX0nWhhp9U5D
DIbR0iYNz0Uzy4+n9ucOLbvZn69lSKSTmkmjFyh3Aj9qWcOthjSByOVjJFXMVJLV
8mWrhtgxYn9lAfaksT4oTirTIr6yGsJojyYU0wRvsSDzc4JbpoAf0hAze53x8QSS
pKoOVmZV2f8ni/bhAuNJIsPhCAGG0zpMCxeFnaTMTg+qwyXPwdRVVmRsOzMFj+YB
oC7mwf3zR5dw37JAOL0u+u/hlFyHVUG6KSmpY0GYtb3pCqdg3Oo9trxnshm+om2R
`pragma protect end_protected
