-- megafunction wizard: %Stratix V Transceiver Native PHY v15.1%
-- GENERATION: XML
-- gx_std_x5.vhd

-- Generated using ACDS version 15.1 185

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity gx_std_x5 is
	port (
		pll_powerdown           : in  std_logic_vector(0 downto 0)   := (others => '0'); --           pll_powerdown.pll_powerdown
		tx_analogreset          : in  std_logic_vector(4 downto 0)   := (others => '0'); --          tx_analogreset.tx_analogreset
		tx_digitalreset         : in  std_logic_vector(4 downto 0)   := (others => '0'); --         tx_digitalreset.tx_digitalreset
		tx_serial_data          : out std_logic_vector(4 downto 0);                      --          tx_serial_data.tx_serial_data
		ext_pll_clk             : in  std_logic_vector(4 downto 0)   := (others => '0'); --             ext_pll_clk.ext_pll_clk
		rx_analogreset          : in  std_logic_vector(4 downto 0)   := (others => '0'); --          rx_analogreset.rx_analogreset
		rx_digitalreset         : in  std_logic_vector(4 downto 0)   := (others => '0'); --         rx_digitalreset.rx_digitalreset
		rx_cdr_refclk           : in  std_logic_vector(0 downto 0)   := (others => '0'); --           rx_cdr_refclk.rx_cdr_refclk
		rx_serial_data          : in  std_logic_vector(4 downto 0)   := (others => '0'); --          rx_serial_data.rx_serial_data
		rx_is_lockedtoref       : out std_logic_vector(4 downto 0);                      --       rx_is_lockedtoref.rx_is_lockedtoref
		rx_is_lockedtodata      : out std_logic_vector(4 downto 0);                      --      rx_is_lockedtodata.rx_is_lockedtodata
		rx_seriallpbken         : in  std_logic_vector(4 downto 0)   := (others => '0'); --         rx_seriallpbken.rx_seriallpbken
		tx_std_coreclkin        : in  std_logic_vector(4 downto 0)   := (others => '0'); --        tx_std_coreclkin.tx_std_coreclkin
		rx_std_coreclkin        : in  std_logic_vector(4 downto 0)   := (others => '0'); --        rx_std_coreclkin.rx_std_coreclkin
		tx_std_clkout           : out std_logic_vector(4 downto 0);                      --           tx_std_clkout.tx_std_clkout
		rx_std_clkout           : out std_logic_vector(4 downto 0);                      --           rx_std_clkout.rx_std_clkout
		tx_std_polinv           : in  std_logic_vector(4 downto 0)   := (others => '0'); --           tx_std_polinv.tx_std_polinv
		rx_std_polinv           : in  std_logic_vector(4 downto 0)   := (others => '0'); --           rx_std_polinv.rx_std_polinv
		tx_cal_busy             : out std_logic_vector(4 downto 0);                      --             tx_cal_busy.tx_cal_busy
		rx_cal_busy             : out std_logic_vector(4 downto 0);                      --             rx_cal_busy.rx_cal_busy
		reconfig_to_xcvr        : in  std_logic_vector(349 downto 0) := (others => '0'); --        reconfig_to_xcvr.reconfig_to_xcvr
		reconfig_from_xcvr      : out std_logic_vector(229 downto 0);                    --      reconfig_from_xcvr.reconfig_from_xcvr
		tx_parallel_data        : in  std_logic_vector(199 downto 0) := (others => '0'); --        tx_parallel_data.tx_parallel_data
		unused_tx_parallel_data : in  std_logic_vector(119 downto 0) := (others => '0'); -- unused_tx_parallel_data.unused_tx_parallel_data
		rx_parallel_data        : out std_logic_vector(199 downto 0);                    --        rx_parallel_data.rx_parallel_data
		unused_rx_parallel_data : out std_logic_vector(119 downto 0)                     -- unused_rx_parallel_data.unused_rx_parallel_data
	);
end entity gx_std_x5;

architecture rtl of gx_std_x5 is
	component altera_xcvr_native_sv is
		generic (
			tx_enable                       : integer := 1;
			rx_enable                       : integer := 1;
			enable_std                      : integer := 0;
			enable_teng                     : integer := 0;
			data_path_select                : string  := "pma_direct";
			channels                        : integer := 1;
			bonded_mode                     : string  := "non_bonded";
			data_rate                       : string  := "";
			pma_width                       : integer := 80;
			tx_pma_clk_div                  : integer := 1;
			tx_pma_txdetectrx_ctrl          : integer := 0;
			pll_reconfig_enable             : integer := 0;
			pll_external_enable             : integer := 0;
			pll_data_rate                   : string  := "0 Mbps";
			pll_type                        : string  := "CMU";
			pll_network_select              : string  := "x1";
			plls                            : integer := 1;
			pll_select                      : integer := 0;
			pll_refclk_cnt                  : integer := 1;
			pll_refclk_select               : string  := "0";
			pll_refclk_freq                 : string  := "125.0 MHz";
			pll_feedback_path               : string  := "internal";
			cdr_reconfig_enable             : integer := 0;
			cdr_refclk_cnt                  : integer := 1;
			cdr_refclk_select               : integer := 0;
			cdr_refclk_freq                 : string  := "";
			rx_ppm_detect_threshold         : string  := "1000";
			rx_clkslip_enable               : integer := 0;
			std_protocol_hint               : string  := "basic";
			std_pcs_pma_width               : integer := 10;
			std_low_latency_bypass_enable   : integer := 0;
			std_tx_pcfifo_mode              : string  := "low_latency";
			std_rx_pcfifo_mode              : string  := "low_latency";
			std_rx_byte_order_enable        : integer := 0;
			std_rx_byte_order_mode          : string  := "manual";
			std_rx_byte_order_width         : integer := 10;
			std_rx_byte_order_symbol_count  : integer := 1;
			std_rx_byte_order_pattern       : string  := "0";
			std_rx_byte_order_pad           : string  := "0";
			std_tx_byte_ser_enable          : integer := 0;
			std_rx_byte_deser_enable        : integer := 0;
			std_tx_8b10b_enable             : integer := 0;
			std_tx_8b10b_disp_ctrl_enable   : integer := 0;
			std_rx_8b10b_enable             : integer := 0;
			std_rx_rmfifo_enable            : integer := 0;
			std_rx_rmfifo_pattern_p         : string  := "00000";
			std_rx_rmfifo_pattern_n         : string  := "00000";
			std_tx_bitslip_enable           : integer := 0;
			std_rx_word_aligner_mode        : string  := "bit_slip";
			std_rx_word_aligner_pattern_len : integer := 7;
			std_rx_word_aligner_pattern     : string  := "0000000000";
			std_rx_word_aligner_rknumber    : integer := 3;
			std_rx_word_aligner_renumber    : integer := 3;
			std_rx_word_aligner_rgnumber    : integer := 3;
			std_rx_run_length_val           : integer := 31;
			std_tx_bitrev_enable            : integer := 0;
			std_rx_bitrev_enable            : integer := 0;
			std_tx_byterev_enable           : integer := 0;
			std_rx_byterev_enable           : integer := 0;
			std_tx_polinv_enable            : integer := 0;
			std_rx_polinv_enable            : integer := 0;
			teng_protocol_hint              : string  := "basic";
			teng_pcs_pma_width              : integer := 40;
			teng_pld_pcs_width              : integer := 40;
			teng_txfifo_mode                : string  := "phase_comp";
			teng_txfifo_full                : integer := 31;
			teng_txfifo_empty               : integer := 0;
			teng_txfifo_pfull               : integer := 23;
			teng_txfifo_pempty              : integer := 2;
			teng_rxfifo_mode                : string  := "phase_comp";
			teng_rxfifo_full                : integer := 31;
			teng_rxfifo_empty               : integer := 0;
			teng_rxfifo_pfull               : integer := 23;
			teng_rxfifo_pempty              : integer := 2;
			teng_rxfifo_align_del           : integer := 0;
			teng_rxfifo_control_del         : integer := 0;
			teng_tx_frmgen_enable           : integer := 0;
			teng_tx_frmgen_user_length      : integer := 2048;
			teng_tx_frmgen_burst_enable     : integer := 0;
			teng_rx_frmsync_enable          : integer := 0;
			teng_rx_frmsync_user_length     : integer := 2048;
			teng_frmgensync_diag_word       : string  := "6400000000000000";
			teng_frmgensync_scrm_word       : string  := "2800000000000000";
			teng_frmgensync_skip_word       : string  := "1e1e1e1e1e1e1e1e";
			teng_frmgensync_sync_word       : string  := "78f678f678f678f6";
			teng_tx_sh_err                  : integer := 0;
			teng_tx_crcgen_enable           : integer := 0;
			teng_rx_crcchk_enable           : integer := 0;
			teng_tx_64b66b_enable           : integer := 0;
			teng_rx_64b66b_enable           : integer := 0;
			teng_tx_scram_enable            : integer := 0;
			teng_tx_scram_user_seed         : string  := "000000000000000";
			teng_rx_descram_enable          : integer := 0;
			teng_tx_dispgen_enable          : integer := 0;
			teng_rx_dispchk_enable          : integer := 0;
			teng_rx_blksync_enable          : integer := 0;
			teng_tx_polinv_enable           : integer := 0;
			teng_tx_bitslip_enable          : integer := 0;
			teng_rx_polinv_enable           : integer := 0;
			teng_rx_bitslip_enable          : integer := 0
		);
		port (
			pll_powerdown             : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- pll_powerdown
			tx_analogreset            : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- tx_analogreset
			tx_digitalreset           : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- tx_digitalreset
			tx_serial_data            : out std_logic_vector(4 downto 0);                      -- tx_serial_data
			ext_pll_clk               : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- ext_pll_clk
			rx_analogreset            : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_analogreset
			rx_digitalreset           : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_digitalreset
			rx_cdr_refclk             : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- rx_cdr_refclk
			rx_serial_data            : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_serial_data
			rx_is_lockedtoref         : out std_logic_vector(4 downto 0);                      -- rx_is_lockedtoref
			rx_is_lockedtodata        : out std_logic_vector(4 downto 0);                      -- rx_is_lockedtodata
			rx_seriallpbken           : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_seriallpbken
			tx_std_coreclkin          : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- tx_std_coreclkin
			rx_std_coreclkin          : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_std_coreclkin
			tx_std_clkout             : out std_logic_vector(4 downto 0);                      -- tx_std_clkout
			rx_std_clkout             : out std_logic_vector(4 downto 0);                      -- rx_std_clkout
			tx_std_polinv             : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- tx_std_polinv
			rx_std_polinv             : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_std_polinv
			tx_cal_busy               : out std_logic_vector(4 downto 0);                      -- tx_cal_busy
			rx_cal_busy               : out std_logic_vector(4 downto 0);                      -- rx_cal_busy
			reconfig_to_xcvr          : in  std_logic_vector(349 downto 0) := (others => 'X'); -- reconfig_to_xcvr
			reconfig_from_xcvr        : out std_logic_vector(229 downto 0);                    -- reconfig_from_xcvr
			tx_parallel_data          : in  std_logic_vector(319 downto 0) := (others => 'X'); -- unused_tx_parallel_data
			rx_parallel_data          : out std_logic_vector(319 downto 0);                    -- unused_rx_parallel_data
			tx_pll_refclk             : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- tx_pll_refclk
			tx_pma_clkout             : out std_logic_vector(4 downto 0);                      -- tx_pma_clkout
			tx_pma_pclk               : out std_logic_vector(4 downto 0);                      -- tx_pma_pclk
			tx_pma_parallel_data      : in  std_logic_vector(399 downto 0) := (others => 'X'); -- tx_pma_parallel_data
			pll_locked                : out std_logic_vector(0 downto 0);                      -- pll_locked
			rx_pma_clkout             : out std_logic_vector(4 downto 0);                      -- rx_pma_clkout
			rx_pma_pclk               : out std_logic_vector(4 downto 0);                      -- rx_pma_pclk
			rx_pma_parallel_data      : out std_logic_vector(399 downto 0);                    -- rx_pma_parallel_data
			rx_clkslip                : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_clkslip
			rx_clklow                 : out std_logic_vector(4 downto 0);                      -- rx_clklow
			rx_fref                   : out std_logic_vector(4 downto 0);                      -- rx_fref
			rx_set_locktodata         : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_set_locktodata
			rx_set_locktoref          : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_set_locktoref
			rx_signaldetect           : out std_logic_vector(4 downto 0);                      -- rx_signaldetect
			rx_pma_qpipulldn          : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_pma_qpipulldn
			tx_pma_qpipullup          : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- tx_pma_qpipullup
			tx_pma_qpipulldn          : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- tx_pma_qpipulldn
			tx_pma_txdetectrx         : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- tx_pma_txdetectrx
			tx_pma_rxfound            : out std_logic_vector(4 downto 0);                      -- tx_pma_rxfound
			rx_std_prbs_done          : out std_logic_vector(4 downto 0);                      -- rx_std_prbs_done
			rx_std_prbs_err           : out std_logic_vector(4 downto 0);                      -- rx_std_prbs_err
			tx_std_pcfifo_full        : out std_logic_vector(4 downto 0);                      -- tx_std_pcfifo_full
			tx_std_pcfifo_empty       : out std_logic_vector(4 downto 0);                      -- tx_std_pcfifo_empty
			rx_std_pcfifo_full        : out std_logic_vector(4 downto 0);                      -- rx_std_pcfifo_full
			rx_std_pcfifo_empty       : out std_logic_vector(4 downto 0);                      -- rx_std_pcfifo_empty
			rx_std_byteorder_ena      : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_std_byteorder_ena
			rx_std_byteorder_flag     : out std_logic_vector(4 downto 0);                      -- rx_std_byteorder_flag
			rx_std_rmfifo_full        : out std_logic_vector(4 downto 0);                      -- rx_std_rmfifo_full
			rx_std_rmfifo_empty       : out std_logic_vector(4 downto 0);                      -- rx_std_rmfifo_empty
			rx_std_wa_patternalign    : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_std_wa_patternalign
			rx_std_wa_a1a2size        : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_std_wa_a1a2size
			tx_std_bitslipboundarysel : in  std_logic_vector(24 downto 0)  := (others => 'X'); -- tx_std_bitslipboundarysel
			rx_std_bitslipboundarysel : out std_logic_vector(24 downto 0);                     -- rx_std_bitslipboundarysel
			rx_std_bitslip            : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_std_bitslip
			rx_std_runlength_err      : out std_logic_vector(4 downto 0);                      -- rx_std_runlength_err
			rx_std_bitrev_ena         : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_std_bitrev_ena
			rx_std_byterev_ena        : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_std_byterev_ena
			tx_std_elecidle           : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- tx_std_elecidle
			rx_std_signaldetect       : out std_logic_vector(4 downto 0);                      -- rx_std_signaldetect
			tx_10g_coreclkin          : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- tx_10g_coreclkin
			rx_10g_coreclkin          : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_10g_coreclkin
			tx_10g_clkout             : out std_logic_vector(4 downto 0);                      -- tx_10g_clkout
			rx_10g_clkout             : out std_logic_vector(4 downto 0);                      -- rx_10g_clkout
			rx_10g_clk33out           : out std_logic_vector(4 downto 0);                      -- rx_10g_clk33out
			rx_10g_prbs_err_clr       : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_10g_prbs_err_clr
			rx_10g_prbs_done          : out std_logic_vector(4 downto 0);                      -- rx_10g_prbs_done
			rx_10g_prbs_err           : out std_logic_vector(4 downto 0);                      -- rx_10g_prbs_err
			tx_10g_control            : in  std_logic_vector(44 downto 0)  := (others => 'X'); -- tx_10g_control
			rx_10g_control            : out std_logic_vector(49 downto 0);                     -- rx_10g_control
			tx_10g_data_valid         : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- tx_10g_data_valid
			tx_10g_fifo_full          : out std_logic_vector(4 downto 0);                      -- tx_10g_fifo_full
			tx_10g_fifo_pfull         : out std_logic_vector(4 downto 0);                      -- tx_10g_fifo_pfull
			tx_10g_fifo_empty         : out std_logic_vector(4 downto 0);                      -- tx_10g_fifo_empty
			tx_10g_fifo_pempty        : out std_logic_vector(4 downto 0);                      -- tx_10g_fifo_pempty
			tx_10g_fifo_del           : out std_logic_vector(4 downto 0);                      -- tx_10g_fifo_del
			tx_10g_fifo_insert        : out std_logic_vector(4 downto 0);                      -- tx_10g_fifo_insert
			rx_10g_fifo_rd_en         : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_10g_fifo_rd_en
			rx_10g_data_valid         : out std_logic_vector(4 downto 0);                      -- rx_10g_data_valid
			rx_10g_fifo_full          : out std_logic_vector(4 downto 0);                      -- rx_10g_fifo_full
			rx_10g_fifo_pfull         : out std_logic_vector(4 downto 0);                      -- rx_10g_fifo_pfull
			rx_10g_fifo_empty         : out std_logic_vector(4 downto 0);                      -- rx_10g_fifo_empty
			rx_10g_fifo_pempty        : out std_logic_vector(4 downto 0);                      -- rx_10g_fifo_pempty
			rx_10g_fifo_del           : out std_logic_vector(4 downto 0);                      -- rx_10g_fifo_del
			rx_10g_fifo_insert        : out std_logic_vector(4 downto 0);                      -- rx_10g_fifo_insert
			rx_10g_fifo_align_val     : out std_logic_vector(4 downto 0);                      -- rx_10g_fifo_align_val
			rx_10g_fifo_align_clr     : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_10g_fifo_align_clr
			rx_10g_fifo_align_en      : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_10g_fifo_align_en
			tx_10g_frame              : out std_logic_vector(4 downto 0);                      -- tx_10g_frame
			tx_10g_frame_diag_status  : in  std_logic_vector(9 downto 0)   := (others => 'X'); -- tx_10g_frame_diag_status
			tx_10g_frame_burst_en     : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- tx_10g_frame_burst_en
			rx_10g_frame              : out std_logic_vector(4 downto 0);                      -- rx_10g_frame
			rx_10g_frame_lock         : out std_logic_vector(4 downto 0);                      -- rx_10g_frame_lock
			rx_10g_frame_mfrm_err     : out std_logic_vector(4 downto 0);                      -- rx_10g_frame_mfrm_err
			rx_10g_frame_sync_err     : out std_logic_vector(4 downto 0);                      -- rx_10g_frame_sync_err
			rx_10g_frame_skip_ins     : out std_logic_vector(4 downto 0);                      -- rx_10g_frame_skip_ins
			rx_10g_frame_pyld_ins     : out std_logic_vector(4 downto 0);                      -- rx_10g_frame_pyld_ins
			rx_10g_frame_skip_err     : out std_logic_vector(4 downto 0);                      -- rx_10g_frame_skip_err
			rx_10g_frame_diag_err     : out std_logic_vector(4 downto 0);                      -- rx_10g_frame_diag_err
			rx_10g_frame_diag_status  : out std_logic_vector(9 downto 0);                      -- rx_10g_frame_diag_status
			rx_10g_crc32_err          : out std_logic_vector(4 downto 0);                      -- rx_10g_crc32err
			rx_10g_descram_err        : out std_logic_vector(4 downto 0);                      -- rx_10g_descram_err
			rx_10g_blk_lock           : out std_logic_vector(4 downto 0);                      -- rx_10g_blk_lock
			rx_10g_blk_sh_err         : out std_logic_vector(4 downto 0);                      -- rx_10g_blk_sh_err
			tx_10g_bitslip            : in  std_logic_vector(34 downto 0)  := (others => 'X'); -- tx_10g_bitslip
			rx_10g_bitslip            : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_10g_bitslip
			rx_10g_highber            : out std_logic_vector(4 downto 0);                      -- rx_10g_highber
			rx_10g_highber_clr_cnt    : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_10g_highber_clr_cnt
			rx_10g_clr_errblk_count   : in  std_logic_vector(4 downto 0)   := (others => 'X')  -- rx_10g_clr_errblk_count
		);
	end component altera_xcvr_native_sv;

	signal gx_std_x5_inst_rx_parallel_data : std_logic_vector(319 downto 0); -- port fragment

begin

	gx_std_x5_inst : component altera_xcvr_native_sv
		generic map (
			tx_enable                       => 1,
			rx_enable                       => 1,
			enable_std                      => 1,
			enable_teng                     => 0,
			data_path_select                => "standard",
			channels                        => 5,
			bonded_mode                     => "xN",
			data_rate                       => "4800 Mbps",
			pma_width                       => 20,
			tx_pma_clk_div                  => 1,
			tx_pma_txdetectrx_ctrl          => 0,
			pll_reconfig_enable             => 0,
			pll_external_enable             => 1,
			pll_data_rate                   => "4800 Mbps",
			pll_type                        => "CMU",
			pll_network_select              => "x1",
			plls                            => 1,
			pll_select                      => 0,
			pll_refclk_cnt                  => 1,
			pll_refclk_select               => "0",
			pll_refclk_freq                 => "125.0 MHz",
			pll_feedback_path               => "internal",
			cdr_reconfig_enable             => 0,
			cdr_refclk_cnt                  => 1,
			cdr_refclk_select               => 0,
			cdr_refclk_freq                 => "120.0 MHz",
			rx_ppm_detect_threshold         => "1000",
			rx_clkslip_enable               => 0,
			std_protocol_hint               => "basic",
			std_pcs_pma_width               => 20,
			std_low_latency_bypass_enable   => 0,
			std_tx_pcfifo_mode              => "low_latency",
			std_rx_pcfifo_mode              => "low_latency",
			std_rx_byte_order_enable        => 0,
			std_rx_byte_order_mode          => "manual",
			std_rx_byte_order_width         => 10,
			std_rx_byte_order_symbol_count  => 1,
			std_rx_byte_order_pattern       => "0",
			std_rx_byte_order_pad           => "0",
			std_tx_byte_ser_enable          => 1,
			std_rx_byte_deser_enable        => 1,
			std_tx_8b10b_enable             => 0,
			std_tx_8b10b_disp_ctrl_enable   => 0,
			std_rx_8b10b_enable             => 0,
			std_rx_rmfifo_enable            => 0,
			std_rx_rmfifo_pattern_p         => "00000",
			std_rx_rmfifo_pattern_n         => "00000",
			std_tx_bitslip_enable           => 0,
			std_rx_word_aligner_mode        => "bit_slip",
			std_rx_word_aligner_pattern_len => 7,
			std_rx_word_aligner_pattern     => "0000000000",
			std_rx_word_aligner_rknumber    => 3,
			std_rx_word_aligner_renumber    => 3,
			std_rx_word_aligner_rgnumber    => 3,
			std_rx_run_length_val           => 31,
			std_tx_bitrev_enable            => 0,
			std_rx_bitrev_enable            => 0,
			std_tx_byterev_enable           => 0,
			std_rx_byterev_enable           => 0,
			std_tx_polinv_enable            => 1,
			std_rx_polinv_enable            => 1,
			teng_protocol_hint              => "basic",
			teng_pcs_pma_width              => 40,
			teng_pld_pcs_width              => 40,
			teng_txfifo_mode                => "phase_comp",
			teng_txfifo_full                => 31,
			teng_txfifo_empty               => 0,
			teng_txfifo_pfull               => 23,
			teng_txfifo_pempty              => 2,
			teng_rxfifo_mode                => "phase_comp",
			teng_rxfifo_full                => 31,
			teng_rxfifo_empty               => 0,
			teng_rxfifo_pfull               => 23,
			teng_rxfifo_pempty              => 2,
			teng_rxfifo_align_del           => 0,
			teng_rxfifo_control_del         => 0,
			teng_tx_frmgen_enable           => 0,
			teng_tx_frmgen_user_length      => 2048,
			teng_tx_frmgen_burst_enable     => 0,
			teng_rx_frmsync_enable          => 0,
			teng_rx_frmsync_user_length     => 2048,
			teng_frmgensync_diag_word       => "6400000000000000",
			teng_frmgensync_scrm_word       => "2800000000000000",
			teng_frmgensync_skip_word       => "1e1e1e1e1e1e1e1e",
			teng_frmgensync_sync_word       => "78f678f678f678f6",
			teng_tx_sh_err                  => 0,
			teng_tx_crcgen_enable           => 0,
			teng_rx_crcchk_enable           => 0,
			teng_tx_64b66b_enable           => 0,
			teng_rx_64b66b_enable           => 0,
			teng_tx_scram_enable            => 0,
			teng_tx_scram_user_seed         => "000000000000000",
			teng_rx_descram_enable          => 0,
			teng_tx_dispgen_enable          => 0,
			teng_rx_dispchk_enable          => 0,
			teng_rx_blksync_enable          => 0,
			teng_tx_polinv_enable           => 0,
			teng_tx_bitslip_enable          => 0,
			teng_rx_polinv_enable           => 0,
			teng_rx_bitslip_enable          => 0
		)
		port map (
			pll_powerdown                    => pll_powerdown,                                                                                                                                                                                                                                                                                                                                                                                                      --      pll_powerdown.pll_powerdown
			tx_analogreset                   => tx_analogreset,                                                                                                                                                                                                                                                                                                                                                                                                     --     tx_analogreset.tx_analogreset
			tx_digitalreset                  => tx_digitalreset,                                                                                                                                                                                                                                                                                                                                                                                                    --    tx_digitalreset.tx_digitalreset
			tx_serial_data                   => tx_serial_data,                                                                                                                                                                                                                                                                                                                                                                                                     --     tx_serial_data.tx_serial_data
			ext_pll_clk                      => ext_pll_clk,                                                                                                                                                                                                                                                                                                                                                                                                        --        ext_pll_clk.ext_pll_clk
			rx_analogreset                   => rx_analogreset,                                                                                                                                                                                                                                                                                                                                                                                                     --     rx_analogreset.rx_analogreset
			rx_digitalreset                  => rx_digitalreset,                                                                                                                                                                                                                                                                                                                                                                                                    --    rx_digitalreset.rx_digitalreset
			rx_cdr_refclk                    => rx_cdr_refclk,                                                                                                                                                                                                                                                                                                                                                                                                      --      rx_cdr_refclk.rx_cdr_refclk
			rx_serial_data                   => rx_serial_data,                                                                                                                                                                                                                                                                                                                                                                                                     --     rx_serial_data.rx_serial_data
			rx_is_lockedtoref                => rx_is_lockedtoref,                                                                                                                                                                                                                                                                                                                                                                                                  --  rx_is_lockedtoref.rx_is_lockedtoref
			rx_is_lockedtodata               => rx_is_lockedtodata,                                                                                                                                                                                                                                                                                                                                                                                                 -- rx_is_lockedtodata.rx_is_lockedtodata
			rx_seriallpbken                  => rx_seriallpbken,                                                                                                                                                                                                                                                                                                                                                                                                    --    rx_seriallpbken.rx_seriallpbken
			tx_std_coreclkin                 => tx_std_coreclkin,                                                                                                                                                                                                                                                                                                                                                                                                   --   tx_std_coreclkin.tx_std_coreclkin
			rx_std_coreclkin                 => rx_std_coreclkin,                                                                                                                                                                                                                                                                                                                                                                                                   --   rx_std_coreclkin.rx_std_coreclkin
			tx_std_clkout                    => tx_std_clkout,                                                                                                                                                                                                                                                                                                                                                                                                      --      tx_std_clkout.tx_std_clkout
			rx_std_clkout                    => rx_std_clkout,                                                                                                                                                                                                                                                                                                                                                                                                      --      rx_std_clkout.rx_std_clkout
			tx_std_polinv                    => tx_std_polinv,                                                                                                                                                                                                                                                                                                                                                                                                      --      tx_std_polinv.tx_std_polinv
			rx_std_polinv                    => rx_std_polinv,                                                                                                                                                                                                                                                                                                                                                                                                      --      rx_std_polinv.rx_std_polinv
			tx_cal_busy                      => tx_cal_busy,                                                                                                                                                                                                                                                                                                                                                                                                        --        tx_cal_busy.tx_cal_busy
			rx_cal_busy                      => rx_cal_busy,                                                                                                                                                                                                                                                                                                                                                                                                        --        rx_cal_busy.rx_cal_busy
			reconfig_to_xcvr                 => reconfig_to_xcvr,                                                                                                                                                                                                                                                                                                                                                                                                   --   reconfig_to_xcvr.reconfig_to_xcvr
			reconfig_from_xcvr               => reconfig_from_xcvr,                                                                                                                                                                                                                                                                                                                                                                                                 -- reconfig_from_xcvr.reconfig_from_xcvr
			tx_parallel_data(0 downto 0)     => tx_parallel_data(0 downto 0),                                                                                                                                                                                                                                                                                                                                                                                       --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(1 downto 1)     => tx_parallel_data(1 downto 1),                                                                                                                                                                                                                                                                                                                                                                                       --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(2 downto 2)     => tx_parallel_data(2 downto 2),                                                                                                                                                                                                                                                                                                                                                                                       --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(3 downto 3)     => tx_parallel_data(3 downto 3),                                                                                                                                                                                                                                                                                                                                                                                       --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(4 downto 4)     => tx_parallel_data(4 downto 4),                                                                                                                                                                                                                                                                                                                                                                                       --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(5 downto 5)     => tx_parallel_data(5 downto 5),                                                                                                                                                                                                                                                                                                                                                                                       --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(6 downto 6)     => tx_parallel_data(6 downto 6),                                                                                                                                                                                                                                                                                                                                                                                       --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(7 downto 7)     => tx_parallel_data(7 downto 7),                                                                                                                                                                                                                                                                                                                                                                                       --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(8 downto 8)     => tx_parallel_data(8 downto 8),                                                                                                                                                                                                                                                                                                                                                                                       --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(9 downto 9)     => tx_parallel_data(9 downto 9),                                                                                                                                                                                                                                                                                                                                                                                       --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(10 downto 10)   => unused_tx_parallel_data(0 downto 0),                                                                                                                                                                                                                                                                                                                                                                                --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(11 downto 11)   => tx_parallel_data(10 downto 10),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(12 downto 12)   => tx_parallel_data(11 downto 11),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(13 downto 13)   => tx_parallel_data(12 downto 12),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(14 downto 14)   => tx_parallel_data(13 downto 13),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(15 downto 15)   => tx_parallel_data(14 downto 14),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(16 downto 16)   => tx_parallel_data(15 downto 15),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(17 downto 17)   => tx_parallel_data(16 downto 16),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(18 downto 18)   => tx_parallel_data(17 downto 17),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(19 downto 19)   => tx_parallel_data(18 downto 18),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(20 downto 20)   => tx_parallel_data(19 downto 19),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(21 downto 21)   => unused_tx_parallel_data(1 downto 1),                                                                                                                                                                                                                                                                                                                                                                                --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(22 downto 22)   => tx_parallel_data(20 downto 20),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(23 downto 23)   => tx_parallel_data(21 downto 21),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(24 downto 24)   => tx_parallel_data(22 downto 22),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(25 downto 25)   => tx_parallel_data(23 downto 23),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(26 downto 26)   => tx_parallel_data(24 downto 24),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(27 downto 27)   => tx_parallel_data(25 downto 25),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(28 downto 28)   => tx_parallel_data(26 downto 26),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(29 downto 29)   => tx_parallel_data(27 downto 27),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(30 downto 30)   => tx_parallel_data(28 downto 28),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(31 downto 31)   => tx_parallel_data(29 downto 29),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(32 downto 32)   => unused_tx_parallel_data(2 downto 2),                                                                                                                                                                                                                                                                                                                                                                                --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(33 downto 33)   => tx_parallel_data(30 downto 30),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(34 downto 34)   => tx_parallel_data(31 downto 31),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(35 downto 35)   => tx_parallel_data(32 downto 32),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(36 downto 36)   => tx_parallel_data(33 downto 33),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(37 downto 37)   => tx_parallel_data(34 downto 34),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(38 downto 38)   => tx_parallel_data(35 downto 35),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(39 downto 39)   => tx_parallel_data(36 downto 36),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(40 downto 40)   => tx_parallel_data(37 downto 37),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(41 downto 41)   => tx_parallel_data(38 downto 38),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(42 downto 42)   => tx_parallel_data(39 downto 39),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(43 downto 43)   => unused_tx_parallel_data(3 downto 3),                                                                                                                                                                                                                                                                                                                                                                                --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(44 downto 44)   => unused_tx_parallel_data(4 downto 4),                                                                                                                                                                                                                                                                                                                                                                                --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(45 downto 45)   => unused_tx_parallel_data(5 downto 5),                                                                                                                                                                                                                                                                                                                                                                                --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(46 downto 46)   => unused_tx_parallel_data(6 downto 6),                                                                                                                                                                                                                                                                                                                                                                                --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(47 downto 47)   => unused_tx_parallel_data(7 downto 7),                                                                                                                                                                                                                                                                                                                                                                                --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(48 downto 48)   => unused_tx_parallel_data(8 downto 8),                                                                                                                                                                                                                                                                                                                                                                                --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(49 downto 49)   => unused_tx_parallel_data(9 downto 9),                                                                                                                                                                                                                                                                                                                                                                                --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(50 downto 50)   => unused_tx_parallel_data(10 downto 10),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(51 downto 51)   => unused_tx_parallel_data(11 downto 11),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(52 downto 52)   => unused_tx_parallel_data(12 downto 12),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(53 downto 53)   => unused_tx_parallel_data(13 downto 13),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(54 downto 54)   => unused_tx_parallel_data(14 downto 14),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(55 downto 55)   => unused_tx_parallel_data(15 downto 15),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(56 downto 56)   => unused_tx_parallel_data(16 downto 16),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(57 downto 57)   => unused_tx_parallel_data(17 downto 17),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(58 downto 58)   => unused_tx_parallel_data(18 downto 18),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(59 downto 59)   => unused_tx_parallel_data(19 downto 19),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(60 downto 60)   => unused_tx_parallel_data(20 downto 20),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(61 downto 61)   => unused_tx_parallel_data(21 downto 21),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(62 downto 62)   => unused_tx_parallel_data(22 downto 22),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(63 downto 63)   => unused_tx_parallel_data(23 downto 23),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(64 downto 64)   => tx_parallel_data(40 downto 40),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(65 downto 65)   => tx_parallel_data(41 downto 41),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(66 downto 66)   => tx_parallel_data(42 downto 42),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(67 downto 67)   => tx_parallel_data(43 downto 43),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(68 downto 68)   => tx_parallel_data(44 downto 44),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(69 downto 69)   => tx_parallel_data(45 downto 45),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(70 downto 70)   => tx_parallel_data(46 downto 46),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(71 downto 71)   => tx_parallel_data(47 downto 47),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(72 downto 72)   => tx_parallel_data(48 downto 48),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(73 downto 73)   => tx_parallel_data(49 downto 49),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(74 downto 74)   => unused_tx_parallel_data(24 downto 24),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(75 downto 75)   => tx_parallel_data(50 downto 50),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(76 downto 76)   => tx_parallel_data(51 downto 51),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(77 downto 77)   => tx_parallel_data(52 downto 52),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(78 downto 78)   => tx_parallel_data(53 downto 53),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(79 downto 79)   => tx_parallel_data(54 downto 54),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(80 downto 80)   => tx_parallel_data(55 downto 55),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(81 downto 81)   => tx_parallel_data(56 downto 56),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(82 downto 82)   => tx_parallel_data(57 downto 57),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(83 downto 83)   => tx_parallel_data(58 downto 58),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(84 downto 84)   => tx_parallel_data(59 downto 59),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(85 downto 85)   => unused_tx_parallel_data(25 downto 25),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(86 downto 86)   => tx_parallel_data(60 downto 60),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(87 downto 87)   => tx_parallel_data(61 downto 61),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(88 downto 88)   => tx_parallel_data(62 downto 62),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(89 downto 89)   => tx_parallel_data(63 downto 63),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(90 downto 90)   => tx_parallel_data(64 downto 64),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(91 downto 91)   => tx_parallel_data(65 downto 65),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(92 downto 92)   => tx_parallel_data(66 downto 66),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(93 downto 93)   => tx_parallel_data(67 downto 67),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(94 downto 94)   => tx_parallel_data(68 downto 68),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(95 downto 95)   => tx_parallel_data(69 downto 69),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(96 downto 96)   => unused_tx_parallel_data(26 downto 26),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(97 downto 97)   => tx_parallel_data(70 downto 70),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(98 downto 98)   => tx_parallel_data(71 downto 71),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(99 downto 99)   => tx_parallel_data(72 downto 72),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(100 downto 100) => tx_parallel_data(73 downto 73),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(101 downto 101) => tx_parallel_data(74 downto 74),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(102 downto 102) => tx_parallel_data(75 downto 75),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(103 downto 103) => tx_parallel_data(76 downto 76),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(104 downto 104) => tx_parallel_data(77 downto 77),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(105 downto 105) => tx_parallel_data(78 downto 78),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(106 downto 106) => tx_parallel_data(79 downto 79),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(107 downto 107) => unused_tx_parallel_data(27 downto 27),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(108 downto 108) => unused_tx_parallel_data(28 downto 28),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(109 downto 109) => unused_tx_parallel_data(29 downto 29),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(110 downto 110) => unused_tx_parallel_data(30 downto 30),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(111 downto 111) => unused_tx_parallel_data(31 downto 31),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(112 downto 112) => unused_tx_parallel_data(32 downto 32),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(113 downto 113) => unused_tx_parallel_data(33 downto 33),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(114 downto 114) => unused_tx_parallel_data(34 downto 34),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(115 downto 115) => unused_tx_parallel_data(35 downto 35),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(116 downto 116) => unused_tx_parallel_data(36 downto 36),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(117 downto 117) => unused_tx_parallel_data(37 downto 37),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(118 downto 118) => unused_tx_parallel_data(38 downto 38),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(119 downto 119) => unused_tx_parallel_data(39 downto 39),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(120 downto 120) => unused_tx_parallel_data(40 downto 40),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(121 downto 121) => unused_tx_parallel_data(41 downto 41),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(122 downto 122) => unused_tx_parallel_data(42 downto 42),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(123 downto 123) => unused_tx_parallel_data(43 downto 43),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(124 downto 124) => unused_tx_parallel_data(44 downto 44),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(125 downto 125) => unused_tx_parallel_data(45 downto 45),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(126 downto 126) => unused_tx_parallel_data(46 downto 46),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(127 downto 127) => unused_tx_parallel_data(47 downto 47),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(128 downto 128) => tx_parallel_data(80 downto 80),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(129 downto 129) => tx_parallel_data(81 downto 81),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(130 downto 130) => tx_parallel_data(82 downto 82),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(131 downto 131) => tx_parallel_data(83 downto 83),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(132 downto 132) => tx_parallel_data(84 downto 84),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(133 downto 133) => tx_parallel_data(85 downto 85),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(134 downto 134) => tx_parallel_data(86 downto 86),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(135 downto 135) => tx_parallel_data(87 downto 87),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(136 downto 136) => tx_parallel_data(88 downto 88),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(137 downto 137) => tx_parallel_data(89 downto 89),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(138 downto 138) => unused_tx_parallel_data(48 downto 48),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(139 downto 139) => tx_parallel_data(90 downto 90),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(140 downto 140) => tx_parallel_data(91 downto 91),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(141 downto 141) => tx_parallel_data(92 downto 92),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(142 downto 142) => tx_parallel_data(93 downto 93),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(143 downto 143) => tx_parallel_data(94 downto 94),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(144 downto 144) => tx_parallel_data(95 downto 95),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(145 downto 145) => tx_parallel_data(96 downto 96),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(146 downto 146) => tx_parallel_data(97 downto 97),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(147 downto 147) => tx_parallel_data(98 downto 98),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(148 downto 148) => tx_parallel_data(99 downto 99),                                                                                                                                                                                                                                                                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(149 downto 149) => unused_tx_parallel_data(49 downto 49),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(150 downto 150) => tx_parallel_data(100 downto 100),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(151 downto 151) => tx_parallel_data(101 downto 101),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(152 downto 152) => tx_parallel_data(102 downto 102),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(153 downto 153) => tx_parallel_data(103 downto 103),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(154 downto 154) => tx_parallel_data(104 downto 104),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(155 downto 155) => tx_parallel_data(105 downto 105),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(156 downto 156) => tx_parallel_data(106 downto 106),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(157 downto 157) => tx_parallel_data(107 downto 107),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(158 downto 158) => tx_parallel_data(108 downto 108),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(159 downto 159) => tx_parallel_data(109 downto 109),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(160 downto 160) => unused_tx_parallel_data(50 downto 50),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(161 downto 161) => tx_parallel_data(110 downto 110),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(162 downto 162) => tx_parallel_data(111 downto 111),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(163 downto 163) => tx_parallel_data(112 downto 112),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(164 downto 164) => tx_parallel_data(113 downto 113),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(165 downto 165) => tx_parallel_data(114 downto 114),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(166 downto 166) => tx_parallel_data(115 downto 115),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(167 downto 167) => tx_parallel_data(116 downto 116),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(168 downto 168) => tx_parallel_data(117 downto 117),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(169 downto 169) => tx_parallel_data(118 downto 118),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(170 downto 170) => tx_parallel_data(119 downto 119),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(171 downto 171) => unused_tx_parallel_data(51 downto 51),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(172 downto 172) => unused_tx_parallel_data(52 downto 52),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(173 downto 173) => unused_tx_parallel_data(53 downto 53),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(174 downto 174) => unused_tx_parallel_data(54 downto 54),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(175 downto 175) => unused_tx_parallel_data(55 downto 55),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(176 downto 176) => unused_tx_parallel_data(56 downto 56),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(177 downto 177) => unused_tx_parallel_data(57 downto 57),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(178 downto 178) => unused_tx_parallel_data(58 downto 58),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(179 downto 179) => unused_tx_parallel_data(59 downto 59),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(180 downto 180) => unused_tx_parallel_data(60 downto 60),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(181 downto 181) => unused_tx_parallel_data(61 downto 61),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(182 downto 182) => unused_tx_parallel_data(62 downto 62),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(183 downto 183) => unused_tx_parallel_data(63 downto 63),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(184 downto 184) => unused_tx_parallel_data(64 downto 64),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(185 downto 185) => unused_tx_parallel_data(65 downto 65),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(186 downto 186) => unused_tx_parallel_data(66 downto 66),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(187 downto 187) => unused_tx_parallel_data(67 downto 67),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(188 downto 188) => unused_tx_parallel_data(68 downto 68),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(189 downto 189) => unused_tx_parallel_data(69 downto 69),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(190 downto 190) => unused_tx_parallel_data(70 downto 70),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(191 downto 191) => unused_tx_parallel_data(71 downto 71),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(192 downto 192) => tx_parallel_data(120 downto 120),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(193 downto 193) => tx_parallel_data(121 downto 121),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(194 downto 194) => tx_parallel_data(122 downto 122),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(195 downto 195) => tx_parallel_data(123 downto 123),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(196 downto 196) => tx_parallel_data(124 downto 124),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(197 downto 197) => tx_parallel_data(125 downto 125),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(198 downto 198) => tx_parallel_data(126 downto 126),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(199 downto 199) => tx_parallel_data(127 downto 127),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(200 downto 200) => tx_parallel_data(128 downto 128),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(201 downto 201) => tx_parallel_data(129 downto 129),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(202 downto 202) => unused_tx_parallel_data(72 downto 72),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(203 downto 203) => tx_parallel_data(130 downto 130),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(204 downto 204) => tx_parallel_data(131 downto 131),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(205 downto 205) => tx_parallel_data(132 downto 132),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(206 downto 206) => tx_parallel_data(133 downto 133),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(207 downto 207) => tx_parallel_data(134 downto 134),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(208 downto 208) => tx_parallel_data(135 downto 135),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(209 downto 209) => tx_parallel_data(136 downto 136),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(210 downto 210) => tx_parallel_data(137 downto 137),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(211 downto 211) => tx_parallel_data(138 downto 138),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(212 downto 212) => tx_parallel_data(139 downto 139),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(213 downto 213) => unused_tx_parallel_data(73 downto 73),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(214 downto 214) => tx_parallel_data(140 downto 140),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(215 downto 215) => tx_parallel_data(141 downto 141),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(216 downto 216) => tx_parallel_data(142 downto 142),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(217 downto 217) => tx_parallel_data(143 downto 143),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(218 downto 218) => tx_parallel_data(144 downto 144),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(219 downto 219) => tx_parallel_data(145 downto 145),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(220 downto 220) => tx_parallel_data(146 downto 146),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(221 downto 221) => tx_parallel_data(147 downto 147),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(222 downto 222) => tx_parallel_data(148 downto 148),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(223 downto 223) => tx_parallel_data(149 downto 149),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(224 downto 224) => unused_tx_parallel_data(74 downto 74),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(225 downto 225) => tx_parallel_data(150 downto 150),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(226 downto 226) => tx_parallel_data(151 downto 151),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(227 downto 227) => tx_parallel_data(152 downto 152),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(228 downto 228) => tx_parallel_data(153 downto 153),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(229 downto 229) => tx_parallel_data(154 downto 154),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(230 downto 230) => tx_parallel_data(155 downto 155),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(231 downto 231) => tx_parallel_data(156 downto 156),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(232 downto 232) => tx_parallel_data(157 downto 157),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(233 downto 233) => tx_parallel_data(158 downto 158),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(234 downto 234) => tx_parallel_data(159 downto 159),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(235 downto 235) => unused_tx_parallel_data(75 downto 75),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(236 downto 236) => unused_tx_parallel_data(76 downto 76),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(237 downto 237) => unused_tx_parallel_data(77 downto 77),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(238 downto 238) => unused_tx_parallel_data(78 downto 78),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(239 downto 239) => unused_tx_parallel_data(79 downto 79),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(240 downto 240) => unused_tx_parallel_data(80 downto 80),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(241 downto 241) => unused_tx_parallel_data(81 downto 81),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(242 downto 242) => unused_tx_parallel_data(82 downto 82),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(243 downto 243) => unused_tx_parallel_data(83 downto 83),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(244 downto 244) => unused_tx_parallel_data(84 downto 84),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(245 downto 245) => unused_tx_parallel_data(85 downto 85),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(246 downto 246) => unused_tx_parallel_data(86 downto 86),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(247 downto 247) => unused_tx_parallel_data(87 downto 87),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(248 downto 248) => unused_tx_parallel_data(88 downto 88),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(249 downto 249) => unused_tx_parallel_data(89 downto 89),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(250 downto 250) => unused_tx_parallel_data(90 downto 90),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(251 downto 251) => unused_tx_parallel_data(91 downto 91),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(252 downto 252) => unused_tx_parallel_data(92 downto 92),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(253 downto 253) => unused_tx_parallel_data(93 downto 93),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(254 downto 254) => unused_tx_parallel_data(94 downto 94),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(255 downto 255) => unused_tx_parallel_data(95 downto 95),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(256 downto 256) => tx_parallel_data(160 downto 160),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(257 downto 257) => tx_parallel_data(161 downto 161),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(258 downto 258) => tx_parallel_data(162 downto 162),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(259 downto 259) => tx_parallel_data(163 downto 163),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(260 downto 260) => tx_parallel_data(164 downto 164),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(261 downto 261) => tx_parallel_data(165 downto 165),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(262 downto 262) => tx_parallel_data(166 downto 166),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(263 downto 263) => tx_parallel_data(167 downto 167),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(264 downto 264) => tx_parallel_data(168 downto 168),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(265 downto 265) => tx_parallel_data(169 downto 169),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(266 downto 266) => unused_tx_parallel_data(96 downto 96),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(267 downto 267) => tx_parallel_data(170 downto 170),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(268 downto 268) => tx_parallel_data(171 downto 171),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(269 downto 269) => tx_parallel_data(172 downto 172),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(270 downto 270) => tx_parallel_data(173 downto 173),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(271 downto 271) => tx_parallel_data(174 downto 174),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(272 downto 272) => tx_parallel_data(175 downto 175),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(273 downto 273) => tx_parallel_data(176 downto 176),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(274 downto 274) => tx_parallel_data(177 downto 177),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(275 downto 275) => tx_parallel_data(178 downto 178),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(276 downto 276) => tx_parallel_data(179 downto 179),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(277 downto 277) => unused_tx_parallel_data(97 downto 97),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(278 downto 278) => tx_parallel_data(180 downto 180),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(279 downto 279) => tx_parallel_data(181 downto 181),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(280 downto 280) => tx_parallel_data(182 downto 182),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(281 downto 281) => tx_parallel_data(183 downto 183),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(282 downto 282) => tx_parallel_data(184 downto 184),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(283 downto 283) => tx_parallel_data(185 downto 185),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(284 downto 284) => tx_parallel_data(186 downto 186),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(285 downto 285) => tx_parallel_data(187 downto 187),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(286 downto 286) => tx_parallel_data(188 downto 188),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(287 downto 287) => tx_parallel_data(189 downto 189),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(288 downto 288) => unused_tx_parallel_data(98 downto 98),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(289 downto 289) => tx_parallel_data(190 downto 190),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(290 downto 290) => tx_parallel_data(191 downto 191),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(291 downto 291) => tx_parallel_data(192 downto 192),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(292 downto 292) => tx_parallel_data(193 downto 193),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(293 downto 293) => tx_parallel_data(194 downto 194),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(294 downto 294) => tx_parallel_data(195 downto 195),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(295 downto 295) => tx_parallel_data(196 downto 196),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(296 downto 296) => tx_parallel_data(197 downto 197),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(297 downto 297) => tx_parallel_data(198 downto 198),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(298 downto 298) => tx_parallel_data(199 downto 199),                                                                                                                                                                                                                                                                                                                                                                                   --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(299 downto 299) => unused_tx_parallel_data(99 downto 99),                                                                                                                                                                                                                                                                                                                                                                              --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(300 downto 300) => unused_tx_parallel_data(100 downto 100),                                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(301 downto 301) => unused_tx_parallel_data(101 downto 101),                                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(302 downto 302) => unused_tx_parallel_data(102 downto 102),                                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(303 downto 303) => unused_tx_parallel_data(103 downto 103),                                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(304 downto 304) => unused_tx_parallel_data(104 downto 104),                                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(305 downto 305) => unused_tx_parallel_data(105 downto 105),                                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(306 downto 306) => unused_tx_parallel_data(106 downto 106),                                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(307 downto 307) => unused_tx_parallel_data(107 downto 107),                                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(308 downto 308) => unused_tx_parallel_data(108 downto 108),                                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(309 downto 309) => unused_tx_parallel_data(109 downto 109),                                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(310 downto 310) => unused_tx_parallel_data(110 downto 110),                                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(311 downto 311) => unused_tx_parallel_data(111 downto 111),                                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(312 downto 312) => unused_tx_parallel_data(112 downto 112),                                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(313 downto 313) => unused_tx_parallel_data(113 downto 113),                                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(314 downto 314) => unused_tx_parallel_data(114 downto 114),                                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(315 downto 315) => unused_tx_parallel_data(115 downto 115),                                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(316 downto 316) => unused_tx_parallel_data(116 downto 116),                                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(317 downto 317) => unused_tx_parallel_data(117 downto 117),                                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(318 downto 318) => unused_tx_parallel_data(118 downto 118),                                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(319 downto 319) => unused_tx_parallel_data(119 downto 119),                                                                                                                                                                                                                                                                                                                                                                            --   tx_parallel_data.tx_parallel_data
			rx_parallel_data                 => gx_std_x5_inst_rx_parallel_data,                                                                                                                                                                                                                                                                                                                                                                                    --   rx_parallel_data.rx_parallel_data
			tx_pll_refclk                    => "0",                                                                                                                                                                                                                                                                                                                                                                                                                --        (terminated)
			tx_pma_clkout                    => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_pma_pclk                      => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_pma_parallel_data             => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", --        (terminated)
			pll_locked                       => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_pma_clkout                    => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_pma_pclk                      => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_pma_parallel_data             => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_clkslip                       => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			rx_clklow                        => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_fref                          => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_set_locktodata                => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			rx_set_locktoref                 => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			rx_signaldetect                  => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_pma_qpipulldn                 => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			tx_pma_qpipullup                 => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			tx_pma_qpipulldn                 => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			tx_pma_txdetectrx                => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			tx_pma_rxfound                   => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_prbs_done                 => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_prbs_err                  => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_std_pcfifo_full               => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_std_pcfifo_empty              => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_pcfifo_full               => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_pcfifo_empty              => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_byteorder_ena             => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			rx_std_byteorder_flag            => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_rmfifo_full               => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_rmfifo_empty              => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_wa_patternalign           => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			rx_std_wa_a1a2size               => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			tx_std_bitslipboundarysel        => "0000000000000000000000000",                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			rx_std_bitslipboundarysel        => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_bitslip                   => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			rx_std_runlength_err             => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_bitrev_ena                => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			rx_std_byterev_ena               => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			tx_std_elecidle                  => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			rx_std_signaldetect              => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_10g_coreclkin                 => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			rx_10g_coreclkin                 => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			tx_10g_clkout                    => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_clkout                    => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_clk33out                  => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_prbs_err_clr              => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			rx_10g_prbs_done                 => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_prbs_err                  => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_10g_control                   => "000000000000000000000000000000000000000000000",                                                                                                                                                                                                                                                                                                                                                                    --        (terminated)
			rx_10g_control                   => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_10g_data_valid                => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			tx_10g_fifo_full                 => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_10g_fifo_pfull                => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_10g_fifo_empty                => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_10g_fifo_pempty               => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_10g_fifo_del                  => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_10g_fifo_insert               => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_fifo_rd_en                => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			rx_10g_data_valid                => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_fifo_full                 => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_fifo_pfull                => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_fifo_empty                => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_fifo_pempty               => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_fifo_del                  => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_fifo_insert               => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_fifo_align_val            => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_fifo_align_clr            => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			rx_10g_fifo_align_en             => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			tx_10g_frame                     => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_10g_frame_diag_status         => "0000000000",                                                                                                                                                                                                                                                                                                                                                                                                       --        (terminated)
			tx_10g_frame_burst_en            => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			rx_10g_frame                     => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_frame_lock                => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_frame_mfrm_err            => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_frame_sync_err            => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_frame_skip_ins            => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_frame_pyld_ins            => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_frame_skip_err            => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_frame_diag_err            => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_frame_diag_status         => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_crc32_err                 => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_descram_err               => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_blk_lock                  => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_blk_sh_err                => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_10g_bitslip                   => "00000000000000000000000000000000000",                                                                                                                                                                                                                                                                                                                                                                              --        (terminated)
			rx_10g_bitslip                   => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			rx_10g_highber                   => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_highber_clr_cnt           => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			rx_10g_clr_errblk_count          => "00000"                                                                                                                                                                                                                                                                                                                                                                                                             --        (terminated)
		);

	rx_parallel_data <= gx_std_x5_inst_rx_parallel_data(313 downto 313) & gx_std_x5_inst_rx_parallel_data(312 downto 312) & gx_std_x5_inst_rx_parallel_data(311 downto 311) & gx_std_x5_inst_rx_parallel_data(310 downto 310) & gx_std_x5_inst_rx_parallel_data(309 downto 309) & gx_std_x5_inst_rx_parallel_data(308 downto 308) & gx_std_x5_inst_rx_parallel_data(307 downto 307) & gx_std_x5_inst_rx_parallel_data(306 downto 306) & gx_std_x5_inst_rx_parallel_data(305 downto 305) & gx_std_x5_inst_rx_parallel_data(304 downto 304) & gx_std_x5_inst_rx_parallel_data(297 downto 297) & gx_std_x5_inst_rx_parallel_data(296 downto 296) & gx_std_x5_inst_rx_parallel_data(295 downto 295) & gx_std_x5_inst_rx_parallel_data(294 downto 294) & gx_std_x5_inst_rx_parallel_data(293 downto 293) & gx_std_x5_inst_rx_parallel_data(292 downto 292) & gx_std_x5_inst_rx_parallel_data(291 downto 291) & gx_std_x5_inst_rx_parallel_data(290 downto 290) & gx_std_x5_inst_rx_parallel_data(289 downto 289) & gx_std_x5_inst_rx_parallel_data(288 downto 288) & gx_std_x5_inst_rx_parallel_data(281 downto 281) & gx_std_x5_inst_rx_parallel_data(280 downto 280) & gx_std_x5_inst_rx_parallel_data(279 downto 279) & gx_std_x5_inst_rx_parallel_data(278 downto 278) & gx_std_x5_inst_rx_parallel_data(277 downto 277) & gx_std_x5_inst_rx_parallel_data(276 downto 276) & gx_std_x5_inst_rx_parallel_data(275 downto 275) & gx_std_x5_inst_rx_parallel_data(274 downto 274) & gx_std_x5_inst_rx_parallel_data(273 downto 273) & gx_std_x5_inst_rx_parallel_data(272 downto 272) & gx_std_x5_inst_rx_parallel_data(265 downto 265) & gx_std_x5_inst_rx_parallel_data(264 downto 264) & gx_std_x5_inst_rx_parallel_data(263 downto 263) & gx_std_x5_inst_rx_parallel_data(262 downto 262) & gx_std_x5_inst_rx_parallel_data(261 downto 261) & gx_std_x5_inst_rx_parallel_data(260 downto 260) & gx_std_x5_inst_rx_parallel_data(259 downto 259) & gx_std_x5_inst_rx_parallel_data(258 downto 258) & gx_std_x5_inst_rx_parallel_data(257 downto 257) & gx_std_x5_inst_rx_parallel_data(256 downto 256) & gx_std_x5_inst_rx_parallel_data(249 downto 249) & gx_std_x5_inst_rx_parallel_data(248 downto 248) & gx_std_x5_inst_rx_parallel_data(247 downto 247) & gx_std_x5_inst_rx_parallel_data(246 downto 246) & gx_std_x5_inst_rx_parallel_data(245 downto 245) & gx_std_x5_inst_rx_parallel_data(244 downto 244) & gx_std_x5_inst_rx_parallel_data(243 downto 243) & gx_std_x5_inst_rx_parallel_data(242 downto 242) & gx_std_x5_inst_rx_parallel_data(241 downto 241) & gx_std_x5_inst_rx_parallel_data(240 downto 240) & gx_std_x5_inst_rx_parallel_data(233 downto 233) & gx_std_x5_inst_rx_parallel_data(232 downto 232) & gx_std_x5_inst_rx_parallel_data(231 downto 231) & gx_std_x5_inst_rx_parallel_data(230 downto 230) & gx_std_x5_inst_rx_parallel_data(229 downto 229) & gx_std_x5_inst_rx_parallel_data(228 downto 228) & gx_std_x5_inst_rx_parallel_data(227 downto 227) & gx_std_x5_inst_rx_parallel_data(226 downto 226) & gx_std_x5_inst_rx_parallel_data(225 downto 225) & gx_std_x5_inst_rx_parallel_data(224 downto 224) & gx_std_x5_inst_rx_parallel_data(217 downto 217) & gx_std_x5_inst_rx_parallel_data(216 downto 216) & gx_std_x5_inst_rx_parallel_data(215 downto 215) & gx_std_x5_inst_rx_parallel_data(214 downto 214) & gx_std_x5_inst_rx_parallel_data(213 downto 213) & gx_std_x5_inst_rx_parallel_data(212 downto 212) & gx_std_x5_inst_rx_parallel_data(211 downto 211) & gx_std_x5_inst_rx_parallel_data(210 downto 210) & gx_std_x5_inst_rx_parallel_data(209 downto 209) & gx_std_x5_inst_rx_parallel_data(208 downto 208) & gx_std_x5_inst_rx_parallel_data(201 downto 201) & gx_std_x5_inst_rx_parallel_data(200 downto 200) & gx_std_x5_inst_rx_parallel_data(199 downto 199) & gx_std_x5_inst_rx_parallel_data(198 downto 198) & gx_std_x5_inst_rx_parallel_data(197 downto 197) & gx_std_x5_inst_rx_parallel_data(196 downto 196) & gx_std_x5_inst_rx_parallel_data(195 downto 195) & gx_std_x5_inst_rx_parallel_data(194 downto 194) & gx_std_x5_inst_rx_parallel_data(193 downto 193) & gx_std_x5_inst_rx_parallel_data(192 downto 192) & gx_std_x5_inst_rx_parallel_data(185 downto 185) & gx_std_x5_inst_rx_parallel_data(184 downto 184) & gx_std_x5_inst_rx_parallel_data(183 downto 183) & gx_std_x5_inst_rx_parallel_data(182 downto 182) & gx_std_x5_inst_rx_parallel_data(181 downto 181) & gx_std_x5_inst_rx_parallel_data(180 downto 180) & gx_std_x5_inst_rx_parallel_data(179 downto 179) & gx_std_x5_inst_rx_parallel_data(178 downto 178) & gx_std_x5_inst_rx_parallel_data(177 downto 177) & gx_std_x5_inst_rx_parallel_data(176 downto 176) & gx_std_x5_inst_rx_parallel_data(169 downto 169) & gx_std_x5_inst_rx_parallel_data(168 downto 168) & gx_std_x5_inst_rx_parallel_data(167 downto 167) & gx_std_x5_inst_rx_parallel_data(166 downto 166) & gx_std_x5_inst_rx_parallel_data(165 downto 165) & gx_std_x5_inst_rx_parallel_data(164 downto 164) & gx_std_x5_inst_rx_parallel_data(163 downto 163) & gx_std_x5_inst_rx_parallel_data(162 downto 162) & gx_std_x5_inst_rx_parallel_data(161 downto 161) & gx_std_x5_inst_rx_parallel_data(160 downto 160) & gx_std_x5_inst_rx_parallel_data(153 downto 153) & gx_std_x5_inst_rx_parallel_data(152 downto 152) & gx_std_x5_inst_rx_parallel_data(151 downto 151) & gx_std_x5_inst_rx_parallel_data(150 downto 150) & gx_std_x5_inst_rx_parallel_data(149 downto 149) & gx_std_x5_inst_rx_parallel_data(148 downto 148) & gx_std_x5_inst_rx_parallel_data(147 downto 147) & gx_std_x5_inst_rx_parallel_data(146 downto 146) & gx_std_x5_inst_rx_parallel_data(145 downto 145) & gx_std_x5_inst_rx_parallel_data(144 downto 144) & gx_std_x5_inst_rx_parallel_data(137 downto 137) & gx_std_x5_inst_rx_parallel_data(136 downto 136) & gx_std_x5_inst_rx_parallel_data(135 downto 135) & gx_std_x5_inst_rx_parallel_data(134 downto 134) & gx_std_x5_inst_rx_parallel_data(133 downto 133) & gx_std_x5_inst_rx_parallel_data(132 downto 132) & gx_std_x5_inst_rx_parallel_data(131 downto 131) & gx_std_x5_inst_rx_parallel_data(130 downto 130) & gx_std_x5_inst_rx_parallel_data(129 downto 129) & gx_std_x5_inst_rx_parallel_data(128 downto 128) & gx_std_x5_inst_rx_parallel_data(121 downto 121) & gx_std_x5_inst_rx_parallel_data(120 downto 120) & gx_std_x5_inst_rx_parallel_data(119 downto 119) & gx_std_x5_inst_rx_parallel_data(118 downto 118) & gx_std_x5_inst_rx_parallel_data(117 downto 117) & gx_std_x5_inst_rx_parallel_data(116 downto 116) & gx_std_x5_inst_rx_parallel_data(115 downto 115) & gx_std_x5_inst_rx_parallel_data(114 downto 114) & gx_std_x5_inst_rx_parallel_data(113 downto 113) & gx_std_x5_inst_rx_parallel_data(112 downto 112) & gx_std_x5_inst_rx_parallel_data(105 downto 105) & gx_std_x5_inst_rx_parallel_data(104 downto 104) & gx_std_x5_inst_rx_parallel_data(103 downto 103) & gx_std_x5_inst_rx_parallel_data(102 downto 102) & gx_std_x5_inst_rx_parallel_data(101 downto 101) & gx_std_x5_inst_rx_parallel_data(100 downto 100) & gx_std_x5_inst_rx_parallel_data(99 downto 99) & gx_std_x5_inst_rx_parallel_data(98 downto 98) & gx_std_x5_inst_rx_parallel_data(97 downto 97) & gx_std_x5_inst_rx_parallel_data(96 downto 96) & gx_std_x5_inst_rx_parallel_data(89 downto 89) & gx_std_x5_inst_rx_parallel_data(88 downto 88) & gx_std_x5_inst_rx_parallel_data(87 downto 87) & gx_std_x5_inst_rx_parallel_data(86 downto 86) & gx_std_x5_inst_rx_parallel_data(85 downto 85) & gx_std_x5_inst_rx_parallel_data(84 downto 84) & gx_std_x5_inst_rx_parallel_data(83 downto 83) & gx_std_x5_inst_rx_parallel_data(82 downto 82) & gx_std_x5_inst_rx_parallel_data(81 downto 81) & gx_std_x5_inst_rx_parallel_data(80 downto 80) & gx_std_x5_inst_rx_parallel_data(73 downto 73) & gx_std_x5_inst_rx_parallel_data(72 downto 72) & gx_std_x5_inst_rx_parallel_data(71 downto 71) & gx_std_x5_inst_rx_parallel_data(70 downto 70) & gx_std_x5_inst_rx_parallel_data(69 downto 69) & gx_std_x5_inst_rx_parallel_data(68 downto 68) & gx_std_x5_inst_rx_parallel_data(67 downto 67) & gx_std_x5_inst_rx_parallel_data(66 downto 66) & gx_std_x5_inst_rx_parallel_data(65 downto 65) & gx_std_x5_inst_rx_parallel_data(64 downto 64) & gx_std_x5_inst_rx_parallel_data(57 downto 57) & gx_std_x5_inst_rx_parallel_data(56 downto 56) & gx_std_x5_inst_rx_parallel_data(55 downto 55) & gx_std_x5_inst_rx_parallel_data(54 downto 54) & gx_std_x5_inst_rx_parallel_data(53 downto 53) & gx_std_x5_inst_rx_parallel_data(52 downto 52) & gx_std_x5_inst_rx_parallel_data(51 downto 51) & gx_std_x5_inst_rx_parallel_data(50 downto 50) & gx_std_x5_inst_rx_parallel_data(49 downto 49) & gx_std_x5_inst_rx_parallel_data(48 downto 48) & gx_std_x5_inst_rx_parallel_data(41 downto 41) & gx_std_x5_inst_rx_parallel_data(40 downto 40) & gx_std_x5_inst_rx_parallel_data(39 downto 39) & gx_std_x5_inst_rx_parallel_data(38 downto 38) & gx_std_x5_inst_rx_parallel_data(37 downto 37) & gx_std_x5_inst_rx_parallel_data(36 downto 36) & gx_std_x5_inst_rx_parallel_data(35 downto 35) & gx_std_x5_inst_rx_parallel_data(34 downto 34) & gx_std_x5_inst_rx_parallel_data(33 downto 33) & gx_std_x5_inst_rx_parallel_data(32 downto 32) & gx_std_x5_inst_rx_parallel_data(25 downto 25) & gx_std_x5_inst_rx_parallel_data(24 downto 24) & gx_std_x5_inst_rx_parallel_data(23 downto 23) & gx_std_x5_inst_rx_parallel_data(22 downto 22) & gx_std_x5_inst_rx_parallel_data(21 downto 21) & gx_std_x5_inst_rx_parallel_data(20 downto 20) & gx_std_x5_inst_rx_parallel_data(19 downto 19) & gx_std_x5_inst_rx_parallel_data(18 downto 18) & gx_std_x5_inst_rx_parallel_data(17 downto 17) & gx_std_x5_inst_rx_parallel_data(16 downto 16) & gx_std_x5_inst_rx_parallel_data(9 downto 9) & gx_std_x5_inst_rx_parallel_data(8 downto 8) & gx_std_x5_inst_rx_parallel_data(7 downto 7) & gx_std_x5_inst_rx_parallel_data(6 downto 6) & gx_std_x5_inst_rx_parallel_data(5 downto 5) & gx_std_x5_inst_rx_parallel_data(4 downto 4) & gx_std_x5_inst_rx_parallel_data(3 downto 3) & gx_std_x5_inst_rx_parallel_data(2 downto 2) & gx_std_x5_inst_rx_parallel_data(1 downto 1) & gx_std_x5_inst_rx_parallel_data(0 downto 0);

	unused_rx_parallel_data <= gx_std_x5_inst_rx_parallel_data(319 downto 319) & gx_std_x5_inst_rx_parallel_data(318 downto 318) & gx_std_x5_inst_rx_parallel_data(317 downto 317) & gx_std_x5_inst_rx_parallel_data(316 downto 316) & gx_std_x5_inst_rx_parallel_data(315 downto 315) & gx_std_x5_inst_rx_parallel_data(314 downto 314) & gx_std_x5_inst_rx_parallel_data(303 downto 303) & gx_std_x5_inst_rx_parallel_data(302 downto 302) & gx_std_x5_inst_rx_parallel_data(301 downto 301) & gx_std_x5_inst_rx_parallel_data(300 downto 300) & gx_std_x5_inst_rx_parallel_data(299 downto 299) & gx_std_x5_inst_rx_parallel_data(298 downto 298) & gx_std_x5_inst_rx_parallel_data(287 downto 287) & gx_std_x5_inst_rx_parallel_data(286 downto 286) & gx_std_x5_inst_rx_parallel_data(285 downto 285) & gx_std_x5_inst_rx_parallel_data(284 downto 284) & gx_std_x5_inst_rx_parallel_data(283 downto 283) & gx_std_x5_inst_rx_parallel_data(282 downto 282) & gx_std_x5_inst_rx_parallel_data(271 downto 271) & gx_std_x5_inst_rx_parallel_data(270 downto 270) & gx_std_x5_inst_rx_parallel_data(269 downto 269) & gx_std_x5_inst_rx_parallel_data(268 downto 268) & gx_std_x5_inst_rx_parallel_data(267 downto 267) & gx_std_x5_inst_rx_parallel_data(266 downto 266) & gx_std_x5_inst_rx_parallel_data(255 downto 255) & gx_std_x5_inst_rx_parallel_data(254 downto 254) & gx_std_x5_inst_rx_parallel_data(253 downto 253) & gx_std_x5_inst_rx_parallel_data(252 downto 252) & gx_std_x5_inst_rx_parallel_data(251 downto 251) & gx_std_x5_inst_rx_parallel_data(250 downto 250) & gx_std_x5_inst_rx_parallel_data(239 downto 239) & gx_std_x5_inst_rx_parallel_data(238 downto 238) & gx_std_x5_inst_rx_parallel_data(237 downto 237) & gx_std_x5_inst_rx_parallel_data(236 downto 236) & gx_std_x5_inst_rx_parallel_data(235 downto 235) & gx_std_x5_inst_rx_parallel_data(234 downto 234) & gx_std_x5_inst_rx_parallel_data(223 downto 223) & gx_std_x5_inst_rx_parallel_data(222 downto 222) & gx_std_x5_inst_rx_parallel_data(221 downto 221) & gx_std_x5_inst_rx_parallel_data(220 downto 220) & gx_std_x5_inst_rx_parallel_data(219 downto 219) & gx_std_x5_inst_rx_parallel_data(218 downto 218) & gx_std_x5_inst_rx_parallel_data(207 downto 207) & gx_std_x5_inst_rx_parallel_data(206 downto 206) & gx_std_x5_inst_rx_parallel_data(205 downto 205) & gx_std_x5_inst_rx_parallel_data(204 downto 204) & gx_std_x5_inst_rx_parallel_data(203 downto 203) & gx_std_x5_inst_rx_parallel_data(202 downto 202) & gx_std_x5_inst_rx_parallel_data(191 downto 191) & gx_std_x5_inst_rx_parallel_data(190 downto 190) & gx_std_x5_inst_rx_parallel_data(189 downto 189) & gx_std_x5_inst_rx_parallel_data(188 downto 188) & gx_std_x5_inst_rx_parallel_data(187 downto 187) & gx_std_x5_inst_rx_parallel_data(186 downto 186) & gx_std_x5_inst_rx_parallel_data(175 downto 175) & gx_std_x5_inst_rx_parallel_data(174 downto 174) & gx_std_x5_inst_rx_parallel_data(173 downto 173) & gx_std_x5_inst_rx_parallel_data(172 downto 172) & gx_std_x5_inst_rx_parallel_data(171 downto 171) & gx_std_x5_inst_rx_parallel_data(170 downto 170) & gx_std_x5_inst_rx_parallel_data(159 downto 159) & gx_std_x5_inst_rx_parallel_data(158 downto 158) & gx_std_x5_inst_rx_parallel_data(157 downto 157) & gx_std_x5_inst_rx_parallel_data(156 downto 156) & gx_std_x5_inst_rx_parallel_data(155 downto 155) & gx_std_x5_inst_rx_parallel_data(154 downto 154) & gx_std_x5_inst_rx_parallel_data(143 downto 143) & gx_std_x5_inst_rx_parallel_data(142 downto 142) & gx_std_x5_inst_rx_parallel_data(141 downto 141) & gx_std_x5_inst_rx_parallel_data(140 downto 140) & gx_std_x5_inst_rx_parallel_data(139 downto 139) & gx_std_x5_inst_rx_parallel_data(138 downto 138) & gx_std_x5_inst_rx_parallel_data(127 downto 127) & gx_std_x5_inst_rx_parallel_data(126 downto 126) & gx_std_x5_inst_rx_parallel_data(125 downto 125) & gx_std_x5_inst_rx_parallel_data(124 downto 124) & gx_std_x5_inst_rx_parallel_data(123 downto 123) & gx_std_x5_inst_rx_parallel_data(122 downto 122) & gx_std_x5_inst_rx_parallel_data(111 downto 111) & gx_std_x5_inst_rx_parallel_data(110 downto 110) & gx_std_x5_inst_rx_parallel_data(109 downto 109) & gx_std_x5_inst_rx_parallel_data(108 downto 108) & gx_std_x5_inst_rx_parallel_data(107 downto 107) & gx_std_x5_inst_rx_parallel_data(106 downto 106) & gx_std_x5_inst_rx_parallel_data(95 downto 95) & gx_std_x5_inst_rx_parallel_data(94 downto 94) & gx_std_x5_inst_rx_parallel_data(93 downto 93) & gx_std_x5_inst_rx_parallel_data(92 downto 92) & gx_std_x5_inst_rx_parallel_data(91 downto 91) & gx_std_x5_inst_rx_parallel_data(90 downto 90) & gx_std_x5_inst_rx_parallel_data(79 downto 79) & gx_std_x5_inst_rx_parallel_data(78 downto 78) & gx_std_x5_inst_rx_parallel_data(77 downto 77) & gx_std_x5_inst_rx_parallel_data(76 downto 76) & gx_std_x5_inst_rx_parallel_data(75 downto 75) & gx_std_x5_inst_rx_parallel_data(74 downto 74) & gx_std_x5_inst_rx_parallel_data(63 downto 63) & gx_std_x5_inst_rx_parallel_data(62 downto 62) & gx_std_x5_inst_rx_parallel_data(61 downto 61) & gx_std_x5_inst_rx_parallel_data(60 downto 60) & gx_std_x5_inst_rx_parallel_data(59 downto 59) & gx_std_x5_inst_rx_parallel_data(58 downto 58) & gx_std_x5_inst_rx_parallel_data(47 downto 47) & gx_std_x5_inst_rx_parallel_data(46 downto 46) & gx_std_x5_inst_rx_parallel_data(45 downto 45) & gx_std_x5_inst_rx_parallel_data(44 downto 44) & gx_std_x5_inst_rx_parallel_data(43 downto 43) & gx_std_x5_inst_rx_parallel_data(42 downto 42) & gx_std_x5_inst_rx_parallel_data(31 downto 31) & gx_std_x5_inst_rx_parallel_data(30 downto 30) & gx_std_x5_inst_rx_parallel_data(29 downto 29) & gx_std_x5_inst_rx_parallel_data(28 downto 28) & gx_std_x5_inst_rx_parallel_data(27 downto 27) & gx_std_x5_inst_rx_parallel_data(26 downto 26) & gx_std_x5_inst_rx_parallel_data(15 downto 15) & gx_std_x5_inst_rx_parallel_data(14 downto 14) & gx_std_x5_inst_rx_parallel_data(13 downto 13) & gx_std_x5_inst_rx_parallel_data(12 downto 12) & gx_std_x5_inst_rx_parallel_data(11 downto 11) & gx_std_x5_inst_rx_parallel_data(10 downto 10);

end architecture rtl; -- of gx_std_x5
-- Retrieval info: <?xml version="1.0"?>
--<!--
--	Generated by Altera MegaWizard Launcher Utility version 1.0
--	************************************************************
--	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--	************************************************************
--	Copyright (C) 1991-2016 Altera Corporation
--	Any megafunction design, and related net list (encrypted or decrypted),
--	support information, device programming or simulation file, and any other
--	associated documentation or information provided by Altera or a partner
--	under Altera's Megafunction Partnership Program may be used only to
--	program PLD devices (but not masked PLD devices) from Altera.  Any other
--	use of such megafunction design, net list, support information, device
--	programming or simulation file, or any other related documentation or
--	information is prohibited for any other purpose, including, but not
--	limited to modification, reverse engineering, de-compiling, or use with
--	any other silicon devices, unless such use is explicitly licensed under
--	a separate agreement with Altera or a megafunction partner.  Title to
--	the intellectual property, including patents, copyrights, trademarks,
--	trade secrets, or maskworks, embodied in any such megafunction design,
--	net list, support information, device programming or simulation file, or
--	any other related documentation or information provided by Altera or a
--	megafunction partner, remains with Altera, the megafunction partner, or
--	their respective licensors.  No other licenses, including any licenses
--	needed under any third party's intellectual property, are provided herein.
---->
-- Retrieval info: <instance entity-name="altera_xcvr_native_sv" version="15.1" >
-- Retrieval info: 	<generic name="device_family" value="Stratix V" />
-- Retrieval info: 	<generic name="show_advanced_features" value="0" />
-- Retrieval info: 	<generic name="device_speedgrade" value="fastest" />
-- Retrieval info: 	<generic name="message_level" value="error" />
-- Retrieval info: 	<generic name="tx_enable" value="1" />
-- Retrieval info: 	<generic name="rx_enable" value="1" />
-- Retrieval info: 	<generic name="enable_std" value="1" />
-- Retrieval info: 	<generic name="enable_teng" value="0" />
-- Retrieval info: 	<generic name="set_data_path_select" value="standard" />
-- Retrieval info: 	<generic name="channels" value="5" />
-- Retrieval info: 	<generic name="bonded_mode" value="xN" />
-- Retrieval info: 	<generic name="enable_simple_interface" value="1" />
-- Retrieval info: 	<generic name="set_data_rate" value="4800" />
-- Retrieval info: 	<generic name="pma_direct_width" value="80" />
-- Retrieval info: 	<generic name="tx_pma_clk_div" value="1" />
-- Retrieval info: 	<generic name="pll_reconfig_enable" value="0" />
-- Retrieval info: 	<generic name="pll_external_enable" value="1" />
-- Retrieval info: 	<generic name="plls" value="1" />
-- Retrieval info: 	<generic name="pll_select" value="0" />
-- Retrieval info: 	<generic name="pll_refclk_cnt" value="1" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll0_pll_type" value="CMU" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll1_pll_type" value="CMU" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll2_pll_type" value="CMU" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll3_pll_type" value="CMU" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll0_data_rate" value="1250 Mbps" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll1_data_rate" value="1250 Mbps" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll2_data_rate" value="1250 Mbps" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll3_data_rate" value="1250 Mbps" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll0_refclk_freq" value="125.0 MHz" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll1_refclk_freq" value="125.0 MHz" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll2_refclk_freq" value="125.0 MHz" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll3_refclk_freq" value="125.0 MHz" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll0_refclk_sel" value="0" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll1_refclk_sel" value="0" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll2_refclk_sel" value="0" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll3_refclk_sel" value="0" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll0_clk_network" value="x1" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll1_clk_network" value="x1" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll2_clk_network" value="x1" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll3_clk_network" value="x1" />
-- Retrieval info: 	<generic name="cdr_reconfig_enable" value="0" />
-- Retrieval info: 	<generic name="cdr_refclk_cnt" value="1" />
-- Retrieval info: 	<generic name="cdr_refclk_select" value="0" />
-- Retrieval info: 	<generic name="set_cdr_refclk_freq" value="120.0 MHz" />
-- Retrieval info: 	<generic name="rx_ppm_detect_threshold" value="1000" />
-- Retrieval info: 	<generic name="enable_port_tx_pma_qpipullup" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_pma_qpipulldn" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_pma_txdetectrx" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_pma_rxfound" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_pma_pclk" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_pma_qpipulldn" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_pma_clkout" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_pma_pclk" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_is_lockedtodata" value="1" />
-- Retrieval info: 	<generic name="enable_port_rx_is_lockedtoref" value="1" />
-- Retrieval info: 	<generic name="enable_ports_rx_manual_cdr_mode" value="0" />
-- Retrieval info: 	<generic name="rx_clkslip_enable" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_signaldetect" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_seriallpbken" value="1" />
-- Retrieval info: 	<generic name="std_protocol_hint" value="basic" />
-- Retrieval info: 	<generic name="std_pcs_pma_width" value="20" />
-- Retrieval info: 	<generic name="std_low_latency_bypass_enable" value="0" />
-- Retrieval info: 	<generic name="std_tx_pcfifo_mode" value="low_latency" />
-- Retrieval info: 	<generic name="std_rx_pcfifo_mode" value="low_latency" />
-- Retrieval info: 	<generic name="enable_port_tx_std_pcfifo_full" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_std_pcfifo_empty" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_pcfifo_full" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_pcfifo_empty" value="0" />
-- Retrieval info: 	<generic name="std_rx_byte_order_enable" value="0" />
-- Retrieval info: 	<generic name="std_rx_byte_order_mode" value="manual" />
-- Retrieval info: 	<generic name="std_rx_byte_order_symbol_count" value="1" />
-- Retrieval info: 	<generic name="std_rx_byte_order_pattern" value="0" />
-- Retrieval info: 	<generic name="std_rx_byte_order_pad" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_byteorder_ena" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_byteorder_flag" value="0" />
-- Retrieval info: 	<generic name="std_tx_byte_ser_enable" value="1" />
-- Retrieval info: 	<generic name="std_rx_byte_deser_enable" value="1" />
-- Retrieval info: 	<generic name="std_tx_8b10b_enable" value="0" />
-- Retrieval info: 	<generic name="std_tx_8b10b_disp_ctrl_enable" value="0" />
-- Retrieval info: 	<generic name="std_rx_8b10b_enable" value="0" />
-- Retrieval info: 	<generic name="std_rx_rmfifo_enable" value="0" />
-- Retrieval info: 	<generic name="std_rx_rmfifo_pattern_p" value="00000" />
-- Retrieval info: 	<generic name="std_rx_rmfifo_pattern_n" value="00000" />
-- Retrieval info: 	<generic name="enable_port_rx_std_rmfifo_full" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_rmfifo_empty" value="0" />
-- Retrieval info: 	<generic name="std_tx_bitslip_enable" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_std_bitslipboundarysel" value="0" />
-- Retrieval info: 	<generic name="std_rx_word_aligner_mode" value="bit_slip" />
-- Retrieval info: 	<generic name="std_rx_word_aligner_pattern_len" value="7" />
-- Retrieval info: 	<generic name="std_rx_word_aligner_pattern" value="0000000000" />
-- Retrieval info: 	<generic name="std_rx_word_aligner_rknumber" value="3" />
-- Retrieval info: 	<generic name="std_rx_word_aligner_renumber" value="3" />
-- Retrieval info: 	<generic name="std_rx_word_aligner_rgnumber" value="3" />
-- Retrieval info: 	<generic name="std_rx_run_length_val" value="31" />
-- Retrieval info: 	<generic name="enable_port_rx_std_wa_patternalign" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_wa_a1a2size" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_bitslipboundarysel" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_bitslip" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_runlength_err" value="0" />
-- Retrieval info: 	<generic name="std_tx_bitrev_enable" value="0" />
-- Retrieval info: 	<generic name="std_rx_bitrev_enable" value="0" />
-- Retrieval info: 	<generic name="std_tx_byterev_enable" value="0" />
-- Retrieval info: 	<generic name="std_rx_byterev_enable" value="0" />
-- Retrieval info: 	<generic name="std_tx_polinv_enable" value="1" />
-- Retrieval info: 	<generic name="std_rx_polinv_enable" value="1" />
-- Retrieval info: 	<generic name="enable_port_rx_std_bitrev_ena" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_byterev_ena" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_std_polinv" value="1" />
-- Retrieval info: 	<generic name="enable_port_rx_std_polinv" value="1" />
-- Retrieval info: 	<generic name="enable_port_tx_std_elecidle" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_signaldetect" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_prbs_status" value="0" />
-- Retrieval info: 	<generic name="teng_protocol_hint" value="basic" />
-- Retrieval info: 	<generic name="teng_pcs_pma_width" value="40" />
-- Retrieval info: 	<generic name="teng_pld_pcs_width" value="40" />
-- Retrieval info: 	<generic name="teng_txfifo_mode" value="phase_comp" />
-- Retrieval info: 	<generic name="teng_txfifo_full" value="31" />
-- Retrieval info: 	<generic name="teng_txfifo_empty" value="0" />
-- Retrieval info: 	<generic name="teng_txfifo_pfull" value="23" />
-- Retrieval info: 	<generic name="teng_txfifo_pempty" value="2" />
-- Retrieval info: 	<generic name="enable_port_tx_10g_fifo_full" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_10g_fifo_pfull" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_10g_fifo_empty" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_10g_fifo_pempty" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_10g_fifo_del" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_10g_fifo_insert" value="0" />
-- Retrieval info: 	<generic name="teng_rxfifo_mode" value="phase_comp" />
-- Retrieval info: 	<generic name="teng_rxfifo_full" value="31" />
-- Retrieval info: 	<generic name="teng_rxfifo_empty" value="0" />
-- Retrieval info: 	<generic name="teng_rxfifo_pfull" value="23" />
-- Retrieval info: 	<generic name="teng_rxfifo_pempty" value="2" />
-- Retrieval info: 	<generic name="teng_rxfifo_align_del" value="0" />
-- Retrieval info: 	<generic name="teng_rxfifo_control_del" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_data_valid" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_fifo_full" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_fifo_pfull" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_fifo_empty" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_fifo_pempty" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_fifo_del" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_fifo_insert" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_fifo_rd_en" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_fifo_align_val" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_fifo_align_clr" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_fifo_align_en" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_clk33out" value="0" />
-- Retrieval info: 	<generic name="teng_tx_frmgen_user_length" value="2048" />
-- Retrieval info: 	<generic name="teng_tx_frmgen_burst_enable" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_10g_frame" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_10g_frame_diag_status" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_10g_frame_burst_en" value="0" />
-- Retrieval info: 	<generic name="teng_rx_frmsync_user_length" value="2048" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_frame" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_frame_lock" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_frame_mfrm_err" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_frame_sync_err" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_frame_pyld_ins" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_frame_skip_ins" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_frame_skip_err" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_frame_diag_err" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_frame_diag_status" value="0" />
-- Retrieval info: 	<generic name="teng_tx_sh_err" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_crc32_err" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_highber" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_highber_clr_cnt" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_clr_errblk_count" value="0" />
-- Retrieval info: 	<generic name="teng_tx_scram_user_seed" value="000000000000000" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_descram_err" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_blk_lock" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_blk_sh_err" value="0" />
-- Retrieval info: 	<generic name="teng_tx_polinv_enable" value="0" />
-- Retrieval info: 	<generic name="teng_tx_bitslip_enable" value="0" />
-- Retrieval info: 	<generic name="teng_rx_polinv_enable" value="0" />
-- Retrieval info: 	<generic name="teng_rx_bitslip_enable" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_10g_bitslip" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_bitslip" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_teng_prbs_status" value="0" />
-- Retrieval info: </instance>
-- IPFS_FILES : gx_std_x5.vho
-- RELATED_FILES: gx_std_x5.vhd, altera_xcvr_functions.sv, sv_pcs.sv, sv_pcs_ch.sv, sv_pma.sv, sv_reconfig_bundle_to_xcvr.sv, sv_reconfig_bundle_to_ip.sv, sv_reconfig_bundle_merger.sv, sv_rx_pma.sv, sv_tx_pma.sv, sv_tx_pma_ch.sv, sv_xcvr_h.sv, sv_xcvr_avmm_csr.sv, sv_xcvr_avmm_dcd.sv, sv_xcvr_avmm.sv, sv_xcvr_data_adapter.sv, sv_xcvr_native.sv, sv_xcvr_plls.sv, alt_xcvr_resync.sv, sv_hssi_10g_rx_pcs_rbc.sv, sv_hssi_10g_tx_pcs_rbc.sv, sv_hssi_8g_rx_pcs_rbc.sv, sv_hssi_8g_tx_pcs_rbc.sv, sv_hssi_8g_pcs_aggregate_rbc.sv, sv_hssi_common_pcs_pma_interface_rbc.sv, sv_hssi_common_pld_pcs_interface_rbc.sv, sv_hssi_pipe_gen1_2_rbc.sv, sv_hssi_pipe_gen3_rbc.sv, sv_hssi_rx_pcs_pma_interface_rbc.sv, sv_hssi_rx_pld_pcs_interface_rbc.sv, sv_hssi_tx_pcs_pma_interface_rbc.sv, sv_hssi_tx_pld_pcs_interface_rbc.sv, altera_xcvr_native_sv_functions_h.sv, altera_xcvr_native_sv.sv
