// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:15 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UXKsC34nxzp2q+oPd93/EI46AMCB2hwnaU34S1x3Py94C50oLuIN+aAuVgBGr2x4
no7rnksVLgiqsR/pDaIr54qA8aviGS+8n81AqZz4zZZRZw2PH+gbhrHE+iGEZKON
cUiUwzl5PgW89guEeG/uAG82IcYYZlwyMuhNAHpXsfw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11856)
42/LNQssEOwstD6T3vbrBsHXgzbOCreUd85SOciSYqrNa+rG2wZDCuXpobMfs3mI
zdmrC0mQu8gRARPfLUTX3Y1rHpzb/7RgszWiiW3AKjnwUkYaJxPbzwfOX7OG1Q+5
II7nj8QckRwfpGn9sGM7exxV4ZRcJvnHqiXNd4n9gBn6kW8Sp/wLao2vA6V6Wa+C
vi9ZNf+OoBt9PoeK9fYDl8r1S7VMxk10TnIaj28R2ea462mJuaEFoLYZKQJjx544
YBUHby8hwtHFOntHiLGU5LgYNZnA5vHLDzsmNO+CEYbcJ1jckucMPDp2dx7FlKo3
7M87g3XOEvQ4y/muQtFafPfxyhKlTGfh1MSkv7syxH/ugCG8loYWhWI7FUV6XMwB
glg0ccnMTcNCmReRLswtN6iijAx+t6cbrAc7c3Nx3G/eSPvB6PnRC1VA1WeVbbWd
szYTRYs8wMC6CH0zAOT1ifOCm3xDNXfmAMaG6A/hKwOMpwZkNfmAZJPTMzhE5NeY
CSgUR/NAXMIhJhdH74kPp79v+WOSCQOHTVVTpE/kdb/RLp3vJRKbTkUXhwE/RKBK
VR9bN/pC9pBvAL0ZeacpZ91D5PQ1R+Liuu49V5d5KeakqngYRwMphFLCOAUu5hAF
JIfC0J/4LsHajPpfNMmLZ8IKfQiKMzNIxmnzDQMjQEFy5NMW6Q99FsIPAvIbQ0SR
mVi5oC1eLmqbZQe7bbfhaJw7PDdUaBmfnxLqtypHxD+MKqRz734vffjPO1/qqOA/
oNqjJHYXccDQJVq8c6BzklxSsV6cWgE2IPm1inBGLEY+sdsDzrLPatCR+IT+t/iD
bPDHeyTpunpICYZDMkgnM3ykVIDSegkYl41Yqgq7Q6mqoSr+ZJlxtLMmesaD8HdO
BR2LxKMyjQtQUdE9KroNPQSBwI3Frz5VULqHFZjWLaWogX+57xbJPEQd6YvqKCV/
bHflUebKpIjOdlwkkTCxxXG7vHbV7qBjMEcb58umI1iQoVoHjlvMYemrttZxy5Fc
+G7Xe2rACIOMVFmk280bfJCaeJg8p2LP0f33oNT473A8xFLUYgG6NERPyOxzikko
jvY3qtOPgsoqE8bOIEjh/8b7SkbD8rp52GrhYq2YJ8ZNkBpVj5nNpsfim04p02Ak
rHZiue7+RuwgPQjhcy07xIY0V39PT/ASqKE0pV8yHSEF13xx2HYzvWYP41Usd9Fu
MN+0kzJ+VWWFu4kOlcNuC3XM0IJ2lHw6ZrMm9LCctVF2V3j5hcA2F+gO3X44dNto
paGrEHORDE86ujLz8KPcKdk8tMNwIXF/pNy4+Xqj7ppMMmpSkXMEqcgJHwtDEIhf
SGVzB8kgCdxt4XPqYTj3MjcWwpFL9AdEVCREJELitgjFHHjx820Mn5fretV6g4kb
rzEg8RRTCh0wxlri/GIJU96VDnXboCtCpYFsZ5okpLuK+s0hR4OA5+Z8E5hkPIl7
SYfnQi42bRBKIdZGdhdz62J5uitGh7YNwEc3C18HglggFJ93ErT2iwwbSxMCXp5F
9D3erP1c4JkxxYIbXsMoHHXnmqoYZA+l/M7+3RenKFhXvXSCk1TR8zvkSj7BOu2U
WKnRO95LrdYglYV6Mxfc194fQm5mnCbjjGHBiSAYNBy31o4fjHuQbfJcHRo58Kiz
UwyKTsZF+iGZ6A3rVZ8zbwpVXxMrMBg6daR3Uj75uewUXK8bno/fH76/bZuybcMG
i1WNV9c/mEoh9qX4bcTJqAq3iEgzlwhVjViiMLYmaAatGO9zbLRLHVSEXoIV0BQg
/cQz6hW4Cs4SM2KVVNHaZxZKiZH1gkk8ELoyLZklbL5RlxCG1Tkzhqx2cPLJ9bm2
HxB9PdnpqRPF8z9zq5h84ek6DerAiD7Q+W8qKlhiv9TcOosZp/ticZMo2wB3d5Ce
DN1zB38xVX0M+EWT4Ac7X0sjO0jIrCiAQQFBwxFrJQzkPytTAiHQ9ePeLd4hQ+Nd
xV4Zuw4MbOrdpq6UddmuIxEHvJNNaGTVBNQqTcrD16GUPIgkFB72hXThT3IP8NxY
RuYQHMdC9Hsl0OhXu2GxlWaEA3LIlNvsEjrX4W9aV2xlpDDhSFE6vausd5arkOtp
NF8G7YIfxD15W8Kp7pVCNIg6r0fIm2vYtEGOXuJGGKvTjqDZI0crWBK1eQXiipG8
imXZylgKr03Xe2fTKPKi/RgNDbm5Y03PW2YFvYMriT37GmMZ6OvEA65ysxdxV95e
DqsH8otGGGk3kfTp8ukmRVhDl+40POk3DOBdu1A9hEttEeI4SMwGV+ij9cJKN7jI
++sD9+utQtICxTVBxEiN53LLn0jlEeEplrrbyKb2nQnww9vdOGZc0nhmNyvXfnAr
zKZkCMmm1AYD3o6fX5PDtEpR8oVtTFLjOhtPLThuKZk3f/BU9bL8+ngjJqTJg4sa
EEx9guwNglynGJ9EievMvMxzkVblWAg2nvmtY1FCRamUORbgxCBiVPSuonYt1A0V
BiCPAKH7e8RDF9RbDiyWAbEVRtY4XAq68GrJWKSzMQspNj/OVDypFWGYMJSZ+iYL
wo7a2DC4Df859I0rGpqXEjw0oKiURrX9dY0kRM9+PNyo650c4hzZB8FnyjwAjujP
WyGkQDLP6vIcOfgJKcLHl6Rab6naamw4O5wewP7RZ331QENMx+zJDnlh7sT34svs
smllpByVNhA8W1zsdCdGowWzwQ6uCF64pbebGeQJtvHYdCzzDWzSxUyv0NsuWv+u
7GNe3QmKxPTF0UGN3txbqyVUjeFMFhUysc66Dophh80W+aa6Osz1x0JbRSw1G2nM
BBpm641aQn2sqmvCI2SjZuPJyDYbj6/8LvYN2xWILaLaNtRhSCnR8UOEJVo7w0UW
2UN+sppX4U71EmglA6BK87Ri7w6MCd+79Ftdj0OSsJKavh1YJOxULDd43o/tmCY4
vM+4DUoWHZyVC721CSkhN0OeikuEp9vozxPXaHIeakVR7nl3av/ygKedZ6Z1P1VR
UxdtL6utvYfvfBJnpuDdfiLDVhO+AZidP1DaVpCG4jMsdeI5qG5mdxShUe4dJhCx
RBywbxS0eDKkqco2aJQdCx/6Jqq6uFZ7DtMdbjtFPIKilOJ/GPOn93ZXKuG2pAIA
iEzAzlH6aJYxBYOL1KF9AhA+iK68f/EO2aulRXzXAm/6HPF2iTQR5r2IZjgOD65o
WLxilPtgL3/ZCSN/P9ugRlJsn8JHvH+6p0LMn9LDQI55iM0RMKeOuSEJq63EOaAJ
cY+23h53gBZjk6k7m2vG+4YWawu/HFgJ2eu75Q/ggZUnZyrysj9Mm0mfSf0uFIvy
qHE48o/S/T8CszLBIJZKWnfVuikREji814MZLYep6K/oGGLgzoeiCvS/yXGMysFu
ynX5szCM6MTx1rMyTDTImd/aTmM7bTDY8b0VXPh4+isewO6Nhj94CdzA/un50Ueu
JlARe/u4hFJvT3AVMIzNckedMOdZubzcOyEFQfwqVjW2HWOw1BCiagklTuI6xw7v
+jYVcLbkOg8d0jIHmTcxiL7lEu1I4AzjT2ISXdDHpc8QGl+fsMt/pVwMfy05EgF2
Vx6/SRYn5HvltowFfldAvuoi/8RvJPA4w7OJSJgQw+rgWlQIJ7Bi0Kr1Dp1n/9tE
Yl9z84CxPzdp3GT4JqpV6JIthFnfjRR2C4TtbIVF3ajKC4mxVLWqL1NbGe8NTre/
W+yvDzI+Sa2uyaMI4yFTSo7iyfTQN2HQkIEHDcVk5de/GtqFaq2aHFniHHIbhC+r
pV0TuTy77iY5GQP4Q5upE+0PuXE8xg4rZWWGXfyoKV8eTQc5KfNPF19qky/Ts8RX
QOn/8OWj5UKG6XLVJ/H5vHXDdZ0ymKOvQRXJJCFGQrPqM2nMYRLS0j2Ny1SYC2zF
cIMNoqxBMum/nMsX6H9qfmqG3hQSu3xeFT/Bky0hUjG8pIr6Sm9Ih5HX5Dk9Cyvs
Fp44/Q5HQMTa2kqo9hdps8h2CMW3MT/ch4fAglAPi7jUYg8Mcac7ighFjoCltgtm
3dpu2L3whkPj9PHZPLOTHA/7PQdzdfTjGp2n806l0cosR6fA4sgpYJuqsAZKibdh
u5yqlsTby36WFQUJtiKjImtkt2YcS+CxmFdiokNGTDxhOKxJu5mUkdVN15HaNdYd
cHMaCe5dnsTSm6aYKq3ClmTpvoMehz7TEDdYoDzknqTEZeyAENu5wyWBV60eJAcG
L5iYMzxvUtiJ0Rn3ZfTX4LuR1NoTrbTi+delV303879OL+4P84J29j5EI2BEUZID
/ePMZViGkk34pu8zBJTgfNxR5OGUcOCbayo/twUaco9pV5HdTM+v9r/4C4b01Sv7
50FYKgCqDaHfMKwK46zJ5NJVudjsF4fR3QCSr5zQ0Q//ofAAW1Vhg7O1KLrYbhTb
vMAswgxZA7h2oF/4FRKSFjOUnAMlcUdeleVBxN47XOGEFaCwv6dca5Glqzr027if
NEbcDZLSl0ZeHMAbz4lX6VyHVsfUnC2JgI7DxTtbqau1vB85CRG+6xfVESYzCBxo
7UvFSZkvxEp4/69RKsk3gce2pkYcBEIHK0sYn8DoxKp6N/QtStaf3canENUBPhuO
XPQH7sCG8se2MEk733tUbKPtnCMXb/t/qH5L6jr4EET7L6OvvCUKUmX0X+hD+v5f
2XxAF5+s/TEDk+DDJ6FwMYpc780D8YI4CjYoxh0Uy0lqDmLwBK2iRAhyowJ4yzLO
5PF2L3J0TpdoxqE3Zr5G3LUF9AfOI0u49a7u7N4lYuMJZ/RkAsWHokZs69wJU1Fz
w5TEyApXBanUNY1cFOZjO+BNc1yrjtajMJKdO9S8SlAZFQ8nAiwsYX49EFwBstAi
iTe4XTPhcn6VYyctNzvrB2pkjyhe/q8mf6TI0pBa1AQsSA9Z2XLFfYGnny3igV5x
qQKPuV7tKdTaCQmV414uLu+KWfSy/S91scH3YnkLnhiAY0FupOv64Twvs2T0L+wC
7xhFNSgFGfJMVKSkBi44qLtO8kWtBPQpO8yzfZ0gb5AUZfZgTmLLaYyZPvlPk0+e
6pcU/RqwTmp0j65Dz37tAnkhBfSWHSi9oqLofQFzsT9hLXykpaufucDBZFuC8nO0
rDdQ8SAg2GuxG/ZvJfb3j/DfuR7b8NuVKlVrSZr07ZDM3DLZh4TGt6wgV67ixEUE
DTltMk8gxYEAD9jN3TPnIJED8F9AOdjuG1wVcgFWvEpMnEBhhde3uj1CWzX5wIsa
qU9GAX9GwlLF5oVabd6IZQ9XarPQlRVtuMhhQuSHL+QYq07LCHMiu6I2PWxiNQFf
+zQkXosghP4AdQvvZPQQT2q1tdYafTblKYCdm4imlcrcs+avdZS9QiC60wKiRSSm
mHM3ExdsY6VZGas+FgLsQBdmgp4vylLaYWz2c5+SIH9zt9PAyLeQqLMYpX/DkTPE
rXvThJZeHFgvpTXAcYQ1IER8Pf+fdlyAbnrVSggliwuQT2BWvCHPhfouaOjlknZJ
ngXZZgUFO+4tWaqbBzgI2sDch0otzDqQ4cR/GpcvCcxvXNUrj1jLvlIOT5dFrbT1
wGPYsXpWQJJ9Dj3UccPngd7KvtMdbmgH59N06sSPfTtJhqcORAa5794iqLY/Oz3s
gKtcGahX95lG9gtMKHTX6vYailjyHjoBcYx7+3QI5Jw0fTWQ2NeEXu4KqOsYgwnv
TgUtZin0eywcF61qB7rpSVBjM8h5yQ90MAjI7e+LzpJ9rl5QObx1yup696UCOhmS
74gqXjFSOaGFUxdfcx8rO1k8eRd+1Ub7UBgfBxXXnYAEzViRP3LRrRFICQCnxcyH
5pmMZPCchR+6pVxGOcXFNci7S3BRP8UrrSTTvERuRnGNAwj9QeK4tfTYt57ashSd
CI9fRrZ9vHQgKFppa7IvgWDPv78+AW1gZJYp8I+HLbAlW1D5eiLWksTAFDPa21sf
jcnoC7r3LLQpZH3QN8D3M8KA4CtN5sU/eadGtzU+FHcFMFh73xQrgGj6ZTOH70//
TQ7EcLhSSrUddnMJbyzg+zchWyAu2Nm9wKlb1oBugap1WeC1Fa4VQUPGlcqBrOHz
5Ed4th1oqOWeVDfdR3w+7qsZd48+FPU4pPlXv7sHREN7QnrfhFNsZhote6D4ruVU
7bJDJf/Y9Bqf6A7Hp6+W3zF3+Wpw+MpTZBERsCywCyrNT9GQdbDECqwbY5VaxNkO
0Lnr20aine6SLJIsajLXSH82IH2GeujlIBb4wF28GkAApNglchqPbstak8qX3+s5
aKPcGTF/H37Cvh+CPKzRyun6ph/iWVGKmU7vZMAgl3N2cpqXbSYoCMXaW4vrR0D7
8nAnJ5tfJzcx5BP7eQ89hfqKuaQdBprA1uKCvPuMbxsFXGlMd4PE74+GG78g2qhb
28bWHcOH+WWGP/QCqbhucMZfgHH9do7SjaphwErNNVWKjJfZgRrHAD9ntJK7PvJW
LObgl3jp3lI1uIOAat6O2wx0gDzDzwPb/y7KXxH0a80bbqyOX/g0mHqkvmTRC3o/
fFNBI39cXx9do75gqRz1iwZ8dGh7FzY4F1xt2CVaV9CXaCmmygKx+Odqshc31Ypm
QW2GuzHpnh2lq6sYLmXFvXXbET+GBrcHZu21GaGnMoybuGSrxLB/qDEq2HtPpliw
/BL60k815ELVBwBAElBY8w7uRb6lK+oVypxcVOgQBWrX3HrAa8Gcl15RkmCKC6V8
2N7She163pUtNaERH6YtQORXZdvZXfE0qJTC8F7dgnGhE77gPN/5CzbFJzIrO/UO
jXhcpY3qWDUTK4XBzofJAhPcoPAay5BNgTJq9cgs5sL8DEtZTGXxEZsGkAefriL4
p8xuBTajHS8rTLsEU1orI6NFPWbkp+Fl/ejZ5eRrNhUdtziw5+VCfyXeec0EgRSt
tnL7A0rHki5qD72vBDu5k7Ubn/jRldK7ZPJjUyfA6g52C1ZtaKOTmaXi3C1tT98C
zeLhnaW+wU64Ttkev4ZTkl3Tvc/5t1Ew2Qd9PIJH9pZMmhKLObJMI2O4ED/wMidB
E5S2tFqi/YwTmQmU6UEr7c7O8qAQt9bQeHTZpwx1njsKXCaMR2Wkyqec8z/txnXR
c3asxCdC/ci7qLeE3XDUAH7vm8FcRRiA5FaMcKKzj1Pm3pfhohhM+nb8znwyKOu9
Lct4ju/ZvjF3n+7JDgvIeHB+Tj41iSWH8MK4jpzNHcqXfusCVzY9wyTjr3dx02gF
XXGdhgWFddbEzRSICff5J03Wo8X1+Q9Rfiar3RLu+zFdA5JL2V0KrlxNc8qoGlsH
4Zsk2lNVxpdcwQkhH4awgHLymmb+BswVJEMzBRsSZKzH3XR53gSlbttRe04n5uXj
fSJ9bs3IpSntmUET0DstpMgH6uE/BWCel7UnxPPc03s6JC44hkvLg61OPZOYw2Kr
WJnCxJNm1JiuDzBvAaGOFLrKKGHXn5dTlsl7w9cDGsoqUg/oYG+MVqDbIanOFR/S
mdsZ8fYCbymsLl9c46vvx109dEV40jhs0DFIRaFBUn3WIdnwyEMPWACQufY4Nte7
ID3Tl0Z/OjVA/823n6UEfLU60MNT/sRGoXfgATeIOkvPwe8pF3IG3Ji6AF9ZK0JA
3dR8WyopYdimyiSGH/0qhrFVmnlN0/vjoh0eqFFM/sB4aVTH8F27K2VTJ31etATi
f8B0WEctVxKzm7T+p2g/nyqVQOzk6UI04qMMeSn9DVqCn7n3vxmrnO2QI75GWLhv
3uCmmg/yIW8YCmX4pGezFOodqiDA1QsarPWPvqJgwOWaVzefXSbq+jDuRbDWuJls
d1goSu5V8dxXQVSQvvnqaTG1E7eXKgqrltgz1O+mbu45IsD571Vdz7JLO+Q5nDoo
x+LBnf151d1toQZRK7h+xVaCfQA1R2fq8ZZHDXK7cFgKQ5Y0+9wCVjCBUe6srDB3
4l3Ufne7WX2HrYM6GL0cDDbeAB0WUIyOXtbmt1ef+ISmV+vEUi17nMIZsThvCJ5i
n1QH3aBSD3DQoeUQOBQ5tUKwS9Ry67KqU14CXp5OjSnr4kDkgILPmYiO1ZEQ3fd0
g7B/un3xEOV2imJt8HuTbLqWXD3pQ8OjYqZg9LXqD3alVfGbxCE5sExmVaOFr3DP
fB5a3l1Tch+ao3JrnnEae/L7ag43ltV9ZKjjPFgSS4I5PvuTJ9gK9KUWuax/W0ZC
VsDSYWtYPQRNENl1PyNcr1USDMY2ONN94cbV0QloZ4cYU+vap1naA4y96SCvJk2c
QWyEbdB1XnEt4AuQT1R7+79RG3hW4EnXE+xm38MfSdaJlqFTcUiwWERrrcdkwn93
E/vhy0libzAoOS9Cl4RT9x4jTj0N+xVhhrvzeScaOceRy7ZvWEk4yRzHE0YOLEVT
VmmGv7U0uxdJMNRm71vrOhps95LQoEKUhk2+KqBACgALWH9w8IhsMbhKtYcDebb6
eB32jC2L2hQorRoU3XQ9bC2tbqKrNrJev6uiDR1dBqK7ZZHZZUQnqVBNT9jSw5/X
jHbi2CmhxGYjFWa52u3GysF3oRdRKwCxM8iZAD3iVexPdKqmXwZqtscItU1zerqJ
jXG6eSC1sPznlon2HTZ17ubhBnaofNR163QcECvoeee+m8o6yNnUkxofCNTw6T9M
0UCFkT2eFbozcL+1xV7S0IQA1oaK6KuElWvolYHWgoS20NHifkO9SxcSUaE6sJDO
J+3qIKjNK/EtIFLNN7WZxmXzMIl5EmPIerZJIaed1/Acbzex5KbpdNWJ3VgmKb1x
fTz3Vn10tndR2GvjBwPGKzRrFbrCRNNUxfjIygQRg4L/y1hsSjKu+slhFsnHzI5b
oz3PgEM5IkWw42ENOoHxeetbCmUbfNpvctqlsqiVY0nUfPS218ZoYrUBiT3rrwWh
KxhNYkwvgprscCMp+kn/WxabZS0YRzK4+MtJRI3igdCz5d2OtgP81hWQ3XN6/uuv
fiaeYIKLljzvIvYj4HHLWmZQRDlAdMYXMo0cXDcgkLnseUT7rVk5prJSaC9Rrtio
Px8kOTGxavtvpYWS3aftYprrkRYnaOp+cvjYlLGcJGW0LNGRzzpDjwLXLkmaWSIt
eTMoDD0kszczw0TyuB9y7T68aJoElDkEh5BUZMLQ5KN8G8xYG99Kc0xWyRg8eceF
0qEGL8VSQMLAPbIVkETz/i6QuBiA6Hpwmm3BPlNyXXIli3U7Bxl130c4yrp2zTl/
PW+n+IDkmCnIsv8AD7lU0qhwbwGiYxEEWkQBjQU1Ezo7P4bLnBqYR6Ka8+d0bLq4
wXNxmNdbE3JZ27pGk1Ssb63F9+0DHZKm1hcm8wcbqGtPcJkdnRiw+IkiJMPwkyBY
uKiyiFJbWwKOzjOuN+UYVt8eWCBCvqB5q88SZwIcLG8SZQMQXXJPvgsvzCXnPP9F
/TKGBrG0sTT2ZJ8/vS9PgV8H4ei/WY8VolOptX+xXHCknBKfCoqVdYpzBHDGFY4l
LcUv8UTbkVPIduf3toJ1cwrlX9Bj1MAYzXMBOjNMeYVVa5Gk3lAblvpTqVyMVmvB
eJjliymX5U1LXTE9Nxt7BEM2yYiLOXPwq1qLwLzPI8ZWtnvbd3LMEMu8paJijvV5
pOyYMwM4FDh3NvpMIoevszAT+t8rTQah7I4MAUk/7uujwcmhnOry7ozbOloncStp
M0XRhHNxWlJs8x5Me/BgcjWj0GaQ4A9omauMl56j+cR5QeQnLKA6XtJdmxZ7OHvF
WOG1Aa/bbHF4T2wrontJ9l/caWvLd9+12VHp4r0WlMcSZyx5b7lyO1/gBE5CMRRX
DQE5Ku039qE9keSNJ2RKzJBLTytKfDLtelmRcSpdbkA0KeJ/Q1SJH5LmFGeeV6J5
/yCPRVgAvJryntmYUNo3o0KyKbP/4Hf7o5hpCHL5GP9KWFw1JcDq1mxEt776gI8j
A0WYLvb7e3eQ/gmIVxPh3OrvNNMDDIYuS+kJwnxmbZRS/bjgCyV0Co/ggu/frEVK
b+1meVDKNVWumeYWmW1VVFiJik6Hcq+uvpZFzRnLu3QqPj3GQUVWlYYIywvbA1cN
eZgxsmcfUglpfz9xIzONaauhnF9gKf9U1nsO7QpyBEBO1fSCnwZ265TTIUtGxrL+
6J6ueZ7H0kBKbB6w3NiZoHSAdvrCZ13NORz8GlPhnRBZVzMTiRWOyWAAOSqikAo/
fB7VU80aWoSJLYVNg1ICFP/lBPw/XfA7mZn74GFZ/fu6OmOPEIB4QwOEvUHMluGQ
XGljqPu+uJXQIMut3refGlkEfgOrnxmvMxGxwi8gKGix4mUXFewV9vL8tlE/Bhec
d8tWzTS+rToMLA4rGaK35D63acXzukuCVPZtGMej4XqEO1T0rfxMwOuFq9UAr2e+
+9UaBZYMMUS0+wO/T4a/x+ek7Rr7fl0bUjWhAc4CxDTz36Ohy7SkC/CG2AHodyK4
j/raASpQivNhFVtYtSKYpHAaUf1wsdKHJEHPgVapj11W/YPVR9nnco3r7wMeFP2j
lwiyCQOIbnGy0AFfIE8IaFxC2cheSGvnP2YWB2h00Wr8tOa453FMk8afjPXiMwcC
GS1yADeDi5FOfXp8dS5thozeSSvY85VbeXbBlqpfC1+MNtIwngFssFd3iXlJyKQq
fObI+J8xMeRGyNf7BdRBVnRl21z4VdMinQYzpKVJbiVb6OumZGwOaLES1VqpVDAy
z6GRhOG++1LOggfmaKc0jh2knMT1r32a4grPeXSgiG3RBGp5vdXuduEAJELv+N3E
NzdO3PnSgjil/GxuH4YcYLzb0fcp9/O9wCV3Rs4Ykt/Q0ju1NCshd6XYWyC9grpi
SLJrWReDrwxVTPaurRw0M+zWxE5fLA0gkzc8eyAjx2lymGtCQtG76qWm3/slloxA
l5YWjML4Ukz1O9kCYbDKOBDKJl2i383N38009+ms09rYxs0MtYkEOirkdVYw8iUh
g9L3RJoxs3wi9UEF/lTaKXd3RCNErHPNJ1Y+kkZkksHBH+DZQ0befiH6vlovInDJ
frXtf0eBQixvP2Dk90TV/zlLh2QDIhYnd4ZheT2le0diM0nCmt01hJcfecMOzE7c
Kdy0XEl4h3Y+aD+NLPKAqIigc3ia1aSHxf4SE9Vz2SzLBHCZ+KzpltUfSjgz251s
lAxpOunQvrhdhQOnUO3r221FbGZChvPC7JOuP7K6Rc0Fwhh0W1ggXpjMK1AcIbBb
6+gr3qvKtfYErxbGIDRZ8AR0m3cRnQvwv5e0PCoD1nYHAknpIGK8rq0T9tyh8d/1
bxa9674Wklh4KyFJfRGxBXkPZ3Srq1halJcJ8c/jnYR4A2k4saOWiU7LsLU96fWV
qhcqIM4Miva3YvYmRq+BKz5kde9YChavJW8vnL5b/biDUHCuo3EcbSMAkp/CL7+j
Ya7iGC4ODkbWGLuzik9W3FoljGM+QYFgjQjniAdR1VdR07CiajuBNkOIcFBO8HpY
dlLQaz9Zp+tiv7obcC5gawaQI5YsXySApfWb/yqSmnlMA6Bc9X8hlWJMUsWrTIb/
QGDJwIhgpAhkADPkO/BdvYqAIAgawa74HS9+whtI3OifwpDtihpNeAxUlHh4hxVg
oIcpCo3x2Ee+4UnexOiA1027QrYi0gm1wXAVmycx33+4O9pS5OHvSxFoHXoi1sN2
llyT9HM/Lvn0rtiyPLQPiwEDnsoxdlFT3hrnJ78GeUZjBV5Sp0bCgDHTv+aep6D/
2VFPUnNBAbpKCwxDn5Q1RnqFT1lUqePRsSlDb3rxzE4YrWfBBaMkk6rOCk28Jgpi
P1w1/7Sc+flPMiHV+PRz3y6GmG8d+ZQvSTltD8FLmsYj7jWio7IWoCV76LHNPJwY
QFxbOxGc5wCZTd71Ew9gdVxdz3DryQLN2VwoGnh/azMnIo0ifs8pJKcJeRbKMHSs
XniKR+ho8kRSqiqTLhZuAnXMCNf6ipyHTnx33zSFFQ1ziy2yceyEsTzV+or84UOB
TGePecJ1to99rEyVjhkhUfyJHtyuZC25zKD1WItpBA7lSbdR4klXf1pvauifq862
kmRvTWtygT72e3oxSksCbHshWL/6jNo3vgh7So8Sa76XSx3cewyhg7PrnPmoCuJN
vn8d8VkkYc/17wDr8aCschRoaq/mB8+SWY16LuEomi5Y3c6zknpRqoT4qrMXZDtb
1ZNtZL3cGEwKH5/TT3hdJj+WB5975CJFN6hAn44/XhZ4ccJHZ5bVzd5DtQPwpUA5
JqFRMuW1p4nZbjZ9jMq8wAtNbTKTcRa3pbdt6+gd23A77DXTUqzAnQlui1pSYu0S
/3FIMtTjjQf7gvuTZLZdDG6Cyy9Eqc2iJFGGazwhhnz2awoFGGMJLn5NNhEEFA5k
KFdhoLyL+LNOvDE/f5msfWnHaV0LfaHuHJopDF9i1Frq9Gk7YsBIWxYXJnUq1W5k
v42l5wahBWlIKM7J7JMJM58fhbaH1iMckwVs6C6h7xbab3FbRrYL/gTYTpFn+kEg
F+lVQRp3I70sM2J0vK63FU4cE197/idx1W+NWavfzVYAqnnLK/YaBGSsa31GnxGk
m+uzc10muGhFie+EFq7SCNS+0ZRUrqLjbmuDJVs3Xtd0KrDXgTUdUW3GU6hrsVyf
9nQ0IG4SZf538yIVJxC06ncmflNFuhsP6g+Mx1EG19pMgPo/DomSeavNavIOipKx
EMoAouKWpPQASLrXtedhcuqT2giUoqCC4kWoWZVb4MDIgkgS4oylGSXA3gPfS76C
wnMptGc9fkEXQ/Q70tQo+6T4twtJn/EXBRyEbmPcGiFc1HdvS1Uk59mee3Lr170H
oDAsy6oPWl7CX0r4KhH7cdKdrbBMwh50e6wuHcFCL8LqrJ7DpeV7bLDQ6UK49uGz
QyRZ+/7MYMkEP55G00sbvkinotLn1EhhlWGOAMuEz/+XkZSleSbYHlKQcjHe4SsO
CaYnzfmGncPtWyitfAJRj39uN1DuuSV7QPTDjiEojCBsTYIcO7MVR7EGVpB58N+T
9sE7oOJdDaAFK0nl96sKhVpFLcoMQ5YJY3D4/clel5JC23PvyFnqZG0348C65dc7
ohYi80AQrV4dhDpmboY9Ji1YoFglnNQNyofsNSLkC0oUvhxX6AOd9FbbR2qYbOW0
YkkkiiybWN+Y+lJEDK03YQbz8H+59tALU4nwbCT1Iy5cxw8SrT6HJnyxBYnzwdRj
B1TFBdsA3tSNV6QkGloJNYRtOklx/cXmz7lk3IAXzPpIG6p5V64qwEgvIqBf64DF
zPQ1/8+I3WEXNkpQfMrG0m841BmPH6QY6CGsTo1YSjfBp/mh+4MHe7nev28P1KJY
Nh5ywL1pZxxGz9LAgVSLegfOv0pKGNNp04rFgcSw2qbdAhxVu4ESZVwfZyVj8vml
52i0dp38BYi2KYVVEjmQgfLVQG/F8fCEhbQyeAhQw+aIwD1JeKfTxL5MOs5KEgMf
g3Y1d9IIGd6Xrmc71PWJcDjHVwFCNr5FcfrR83CLE39VoGO2iBDY2BS0ItuoZkOh
h295yqCrIjy4u/RrUY//iWMXRAewVHXe6ke6V8JrwDz/CA6+jlr16xaAyrv6LATF
3Koe1vaOgmdsNL9qOtIHsAG88ASXNzb6A1XXl5heUwo+m7BjBdv5Q0UjduVhRwUo
X51dhKi+sjaf+7H10CMn7zbpktpGQ8cwvpqyaopTkylEG7AbwrKb6cgHtcZoGRsQ
NZSfsobnA9W6kEN1nCRSuSSS9pQc5Ccnax9ab+Z4bqWTix7hJRIgBS6O241SDQEr
jTNmJIL5RX/7S+lFfeHzXdGFgw/56Tg6kypjW3mcb5D3R3jk9ySjS6l7sCleFypb
lsgJaZiPNi1RDjIDsBLzRNZ5vWRfN7rYj02hh4VWZi93s1ASgpvsgyCCkN9Mtq59
lh4PnVZXWMDOhsht35XXHOSKUZNsx2r8Qsy7xexgcRyxNkPeq8dFjCCCIIsnx1h/
Av8z1+0tY8cUvHLySPLuX+/GdriDlyM3+NBjAked0GI98TPXaMYeC77dYgq9jK9O
lV2aMmJxvM54x+BZYP+Mq7XIOInom4mucv2UbEUR1P3iJ3DuLAqxgLXVtKV3XAB3
T2Y3TRVcdgsSCOPOxuLaznmYYgKfwarhVxZrmkwuPrBuSIGDioIaUXIBG9GuHL0X
7z/t+9DgDMaZ/6vV0I983/zmLgyGvfMMyTiTt7bMm4hZIyBTJn2u1h/GExxBVFjv
Xnl5OnUwJ8Y2H/+9GpMsZ5TY/1ko4HC/cvpgfuuNDPIAphq/DpVFtPV16+NQsOoD
n+zzXhlCACJM5AYut7T9budJP+nD6e4pwcTGTYtlrV4H7sWdQb8LHQKLcrqaIDfD
L823jhuDYVgxUCVcK4vBe3wQa/GIUE+GZHFK9PoMZ3gpFz3DAanE+zfrj3K0zKGM
Jifdskt6n/4+cD+JCkSIvgG/xRp3chXjZWLqptC+dB+SQ1UwnIIfkQt8AZ9rfkYZ
yOAQOIBMmtNBb/SHtECRvNGeLiPQxEgjdpIl4XX4ki7L7o7I2pby5u3nqQMhwACG
CMQB+c5/mV/1X97D77/+29JmujohLMf09fanB8f8n/yK1ebfJ7XRA76rnGX6Hzi0
ntW6P0UQ675sks8PKViVYWSUHrZ1fqP7eXdL0Jz2wSZUL7tlGS5ugCY2TghmjtCm
d/LhpleBRs56Zf/NAhiWZp852K46ekcKr/QQ0vlYM3221nv6KHGLkUuJOM5kh6V8
JYPaGwjPzpW/hiOBweOaKVL/P8Hmykp/StZDVkOr56j/9xk3dqP/0qW6429sITdm
0gSbZ68jMa6qyZGvhXFpv3T3q0wGw4z0LC0CLyUrjGrWNQbvP3ZgY8jKl0BDT0oU
G+Y9Qmynic19IUk+OteFI85WF/QooElhBT9RD/w2gio9xRPCjoTiRskIzJ2iRDuN
+Nrd4NEeUwsblowLy3mICe7yPkucdDfkT/mauqnCqmggpm1EjQQ2fs3C2C/shgqF
1uOqGVRvhbfno2oAtq0pYxpekDpEOLcvCGquEsOuhp+YPRlq9EVS60BfjlH8woKm
+zULQTuf3Q7Z8wGbIN8zuOQqbt5D8g25RvtMmm/OHtK+TFU4SGSDbZhypBwz9NOc
ZJMk2L/QsbLaIh8Npjh13N1o4AgtL1RKQSRt9Ht8y1Je8K4HjkmxI76yM/JIR45K
fqhUUY9Q0O29y8SQ0zSOLT440L3wMEtXQCjTsnwxPsLa0/DYyyKSR2/Y52cxjZqq
Oi2AkjYVpTdHSKpB/OeNqkGEYyy+YwROtCgeqlgwEh0G+t7vu+z5hcJ7Zs5mJwZW
QZMv7P/u99YLXMEG3PWiCbKzWaEnFTd/Vl/JBoAu8LyjVvwpX4SbAeSh8WHV+EZa
1cMCITGb30NMfAB2FH55eE9CgAoaaXMXS+UPSPLkj6zu+ZnuE7x6zx38vjkNpqvi
fOcTPT3dsrpv4SwPM4r532mkSwah/VVSH9q5phTXMS8K3G4Wo/ZyYxqiT80VZ+e7
xSqgFazBH2K3OfIGMobfOuWPsWiFt2Vflf7fZ0vNxWUJAO3biopb+uC6GKSvdcrF
vUvmq2d2cACvo47uI7hUJs0AiX1hZVIyz6rpQRnBLe0wgKm6K7A+KV23S28Nxo7v
O7R0PUPRcL/A8b6YC5y8NMIdjEPXdGTXaHfZw64M2B0351jpyIX/eJTouIRNa501
Wza4qZkhCTiW+/xneoYPdhWThQEigK+AXwEdD6ax8mIzsr6eTeItopA9tDXCQ0TG
s3ozCtv5HLpwDqNxomizLmjhazZgJkx1YvmHPdb7CPrtiaXmi4zuMNvzP8l3R64V
`pragma protect end_protected
