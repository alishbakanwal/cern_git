// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:10 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VRewYMBbw9Whq/eCchDFVz3J4UCPc/N9f4+BYAY1dUjBIHv9mZ7PpIHY/A6GYim6
B5QegILvfzdigNpPDtnKHSD40G3iiIoUojJ3aPHkEd/B0rzB1RHPUi4yXCeTXENS
fCZAo1f46sGZQfz3fsPWVz1r3NRmyKEcQj7MdY7CfII=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 57760)
Cdsvz+gvJ9WqnCYhaKr28VBgyLg1/A5ersFyg5ZpPRF5JznH2FRYhUbyHvHmDUua
kgKY/X+ajfiTNLWVrjBLTZkLC2Bl5a+bmrXTvuKu5gDVw+0tepQUNvkah0a/GvDs
hterBFWff86DmJdZxu12Mp7D0wboN7Hcaj97h6/jyaUyb+qnVFQsYH3EPhJDiN5i
rKyWUsT7KE/V7bUtq+tiLtzlJFENs6oARCp/75uH9Z8jOKMLzTxLptJkLz8NEmUA
jyaaTGRlJCv4+eeKR0ELuuvnO9ab+jp+3LEUEgXuva8Wdwu1tLwvW6pe18SPZEg4
d+wOHGoo49UMgL5foIeOy8Dd8AQhZz3y5B26U+TbMP7KfWADnQiz7GMuXVS1JlxE
wNvP9BByYB9zPhpneczRR5/0fvAdO4FeuqbRo6MNfTDkuBmwhwjFw0olcRomijM7
0mX7C+KSW2Pr9VRWuhWz2wEtVt1SASYv+B1E7pUzvBbyuy4RqvSZPrZk8/JNXftU
wV3XS7lRswOPPgReQvozx9v3Q/WCxKRO8ywXhVXIFKKqIfug4zk0hcAc5Ye0wcc8
l5Qnvu58b0XRyAiigSbCt4LNlOaNzd3YzKVyZG1TkvUZLbsKW71+YJhyWhDfOpFr
HP/SbvI0pD0904DAn2/2W83agEWJVvLZn69QwGjCUxMWIqCKcacmC4xbv5aeKnlC
r5fsiRZACjY62VrPIb1v7Hv+bELVCQn75VSXS7qEgiIX4jAztiDvI7mPjJbJWn6b
GpnqdnGCpjJig+GZIxX6SK5Lnea/VDJghNp/T031p5PSPA61At3gt/sqn/57VuAp
CyLoC9nOmyVPUEhcafETnh5KT/KkGX7AqwbmSuhKc4jNFvuNuNCdZLKq8yAkuqDK
GhLS7STUJWDE+53tDetHf1PhWA8Pw+FjdIbNaRzB4CLtCRC5E5xsCuoK13VjlKcf
R2SRGYQt6T9QFvXGySyximdGQDr3LgYz/sQai43ip9iGgjqsKRneFtEQQKW640DW
MA1Isy8Ob662vDoq5ycrUJjow1atE3QKe1sBHpnZDsh3h70+219o+uoVX3Fch/Hu
ulsQ6LJAwUBcVappIOJI8hfWFFxs1Dci5fy7dt+wqPHry3xYxdLYRgALZ49StBXb
Sb41SPsY+BVBAd/dhF/uuCKehKUoWIyAJ3bRELpxJv5nXW4h2OoWFnjxh5XT1K5W
Zqi2anaINsVZj2+p/8YLFivgsNdb9WqR4MAEq1ipxlTw9IF7xAUa/EKwugkwBbEP
7vqVyorHT0+R7QnvPXXBg6oUtCE5ynkA7unsCYLQcICem7/26NIbUAX53WiyC5ad
hcMzq0DKZcUj9HdJ95KE/Q2MJX6v917AqQL8yMh5bJ/L5a4sXmhvqZc0l1uT8E87
QVf+CwOaclOYrQCL+hDAanAJy2QpAqsSvO5vReOe7B8HZTEIBeUdkzGGGdhGF5C7
KCQVuZJ3Aq41TEBvvILBpj/SGYjmVYQKEh6PLgzqyvwu23ZX+f4LRRNjnFaPkieZ
kstOdqBEzUg13P87Wkp6kqB8wKtgE6ls5jJcEYsTr9kDOiMh+b7wRtgma4V3iRp3
6bnFfCbNq7xujI4quwqJuE7jmqPcajGsFNySncUebWVkmSrn5I9ujIoDt1nRlzDq
iVB8UxhVxOuX0f22sy5v7Zlw16JYGJLdoQCFd8HmqT4VPxgdgeScsGfxhGW2N65F
8B2MKmfoD7yb4D/3mGOSbnYjC72MMS1nugcjPVGKkh58Ecck7HIZ6BqQ+SBpLGGz
UrnlnQGXSYGExRlUstf95QjW5XfmBuA1IjQXpsM9H6wIZ2Ag1dWQM2b2v0pWcJiN
t3bu+FtuutCUOEUNnt8FpgfviR8kAP4oLxaz5S6MD6LiNUcHpZtzEe1JYd+O6GOE
5vQmPYr7lThqAGAsmr8Y7HgqOXCwLAvQAW9+i0ZuD5cx1junK0WmPeDS8XWFj39T
0HwCB7Fo1kQWhAZVREx6Pn+oOVkbeIFSoHe6an3V5QgqmV1J8CxLO19kjJdDBIiO
yM+9VwJ+WYW/8xKU8QPPvNl7tiHtzMVrKp+qNkNMYKqZoCMdFmeo+oQPH2FMhToA
3IfZ5AxFmC+6A5WIExT4bTlmlET9hGQidoeH3LtCayJXoHTWY/Nz810sYWbRpDjY
xDm3ptzK0Iw3BGDoN9sWMBfICllHlWCOfeYPojHDnEOZ7v0gnG1fMmDYrvao56UF
vxycmv0XB/y1e6nwVX+Z6kTrGhrEHJ5RQoewYq844OGFWblHO3PMekMLgQbsWL8S
saH4LqzwaiGUx+jlXrJv7lujerFUtTu0hg8oA8o1VERP7W8sC3FmrbeGHz6ySBBa
5UgGSikuaV6wvE/lKUnQd8i4xKYiJQdEtqoaSNvNc18czDyf68221ENFY7J7ubFV
sF0rlez9u74StKUkTMZHY1EDjLXDDZHjwkYhR45u3IzSoYakUt+tlwBCyLXBjEOh
QAC/zmcK64mcbwyAPST635GezW3G64wYDHt961FePYM43xOerkNW30BYBUEB+NWC
ylbKEPRkPcBakU2sAX/IX6pI4jwIKHrQfR1/7AYLG0tcOCstIk4EP47Y4nBdQK0C
xJ0q2/zA7ZQaPZNkvym4XK2KebG9ljfq+0fmlWgsxf2CGArcwEHuzJC89V8BXgL9
zYPZ/8OjgCSWJ5mZY+j15DrA/xu+cy7NorUmhyTTyjYKIf4+0I5K/ZvhPOaeS5/z
s2s1X6bBYnP5rRb65jzVRw9PGBRHwuXsTw2cjCnZM+oTCYwSUx4z6JcQl0qJgxuJ
2B1aNELWpJCClkBxb4Pr6pKfhUBu4VL7APjs9LWs36Poqg9XwNuEuBANjemeAmgz
3wZQ9hxgUetXo1LszYOxmtg5YUJ8rCRT6AYlH0A+lU9G8eQfHX7qkaC66cI+cq6y
HFIHSh7QGzDjnO/5SVU3DUJ8wykR8RrE5YcdCeVUSFEueOkd/32EALTU+P/ReVuu
Z2l4lSnU2o++vrNZYY0TOWPVvZ+lobFC9Au1Mrr3YWjCWeVXqQTsb4h/0GUxmMJf
wGprBgiqPTxKc9nlhlYc94z2dlLbi5vhM04Ju+IFZR2ctgbHlmoDVyMvExjHXDNd
6CRZ+zlVCaiiblujteRNuqCYgTjnqbA4Gvnc9tnGQDLDh6lxiIMTp6++pps7EygD
ZtPo3TwVvslRP+TlVbMiQ6bULEfi7v5AZLlIYreG8sRPy7sys4F4CXl/8zE/allh
pQG091GCH3H6as5jDRGA6164eygqv0vQa0Rbrtjq07W3xExixsst0G7PtZSiSweY
B8kj83x1XofOZq8PbRN3aOo9HbSIW+Wo4f8nXMDXYFQwt6t/T4+hZWENgKERNRRV
4ZobPW7pUHPEjhGvStzlUVOZ1C11js7pQq1OSo60rghHeaNN487Z1ijGugyn/Sc+
p5MDVrTw/Vmj25702Ox/Lcn3olHFmKvqGzXqRJEsRzoeaIrttGMBIcNXXZLJhEN3
FfsujyRlVEWjVl41AWy4S1HpwO+i8pDm92bxmpsDLGYyx2NwQkZ1awi5s9GfAH6B
hKe19a/L2C/aXjOZztITuuXx+Hs3/5aWOq+pmRJf6erHYXsULmWC7M43GBClTe3r
MIdv9PeYBTeib/01gEIJXyDgg8B4r/hpezogHOVE4WWMgN5DmqBsRnXdxPZr6P9w
QoVCU4pYVNih3MkAOiKQy77TTdQirHASHhhriQIK0+ai7K4oAlgwtZtv5M24ITMG
+24mMxF9x2ixiRWRcwNqWu5QMDlC8ZXA8fTg8pgaAu7ZVsYdqD2RM5Qa4U94TMAq
w2C1Veb9rdFwgqfrNI5miuwvcrEgXGJpV4WbD/lwPaZN22BUHWQ1S4iSuKTxr87G
DRrrgHdDWNFnLwFN5/ION4VdoMePTKh/V6l7463GJ3UJh1CZgf3LKZ3yFeK/Ar3m
KziChbHGXt5MO1vQ0h2mzsPSDtAG533H9FjdU0QRM64D5W7kFzoYGmSg37d+jXx4
a6hu8nFu34Y2f2ZboVHVouL6xhi+9mI8BiQQz7v2tpNQnWPwhedcQCMVTvaPEcza
dwsQ6PoU3Toa1qbF2s9z9DDn0sCrMam/jLMF7ELNplhZm2u/RTjIQ20Va1LQCqEe
zCGB3dRK0JTafjS8T+M9LJys7O9e5ByiMGBXBzhUPEm6P3pmB2Ntbd9bT3l75Q6d
4cD//k/TSY1g1IHMJA+iw+D/qMllycsHYAaewt0GGjWrtDSPwdJy2EpH06n1YDav
kppPZPKQtW2JdpZmL66OT3C+p8Sb9OSnJ/jon2XopIJ38hnttz36Wyzm4CTpI7LN
wdSKm8r9jaxgqmE59TQefQLqxBQXJmtSIOwP7irTcKFS01ekHs1Y0X0lncfP8c9f
7d0DxPp53l8y0TgBYwsE7EwkiP+4ZnkadPRCxFW6St/CKQGHRVfQqk+ftuz/EFyF
+hur1Ld/Of98tEIjICRuObDLC5q6KIf0bikvmtDbFwtdujBG37wS150lZApSfAn1
OF3Z3VnEQVG6v+hOB6KcLy/LarWUvKAZwrA15b9B7eT0Hclsz+L1Y/I3TUY7XWyJ
715r7ylH6hoWNCWICx5zdRBCP12BS1aSsDiarkYE8OyEJGzktOPFwFE20aJYslTr
HWKRkWIoQo8FUQ8uFfItH71H1VJmbNbsBMY9NomCsoVFYF3G6bZnZQTOpEHgbf+C
ED65T7/cvbt5WfbYrCWSnk5TYyVIiMh5clJ2E6kVE3wy/UJIOBcgKVUxpBDfdEiT
HdKw7LmbcMcUmRW7OxLKwC+q8dyIjeUCZ/nzpQwSbQBtWpkp3KMob+iKg4rEbl0U
gY1oruU6jkfM7qJyzrdJiQ9Gszc3V8C53dCmV4M6wxsja6UM7v8/zhtTQL4kM5cT
1/4F8amLUCsNLSelGR9FdW6X5IIZ1ctJUGE84eZu3dDL+dX9RjNZUWxD6HxlTcql
zVIN7WNxG7nGf23Vc4MI6wVo8+jNWEWHfWcAd1RyZTOfleJqDmWCDC45pTwpO8o7
nNHvuI9zUtgedk8pslf9VhMIeAFeyzJpbNDh3xFea9L8XV/DKa6TQikh9J3yrlKH
guvVnJMpQRjjAe/fPVNdynro/FTh6DyG0ivmoyoxDwtHf4K0m0di9ZETpQ04dIAd
TpdCvMlp8vuC872+PWM76FSDyiOmcPqsZyUIB6UgODLUUpiDaVwczvQZXjKtRf68
9QpdmprDTqSDRjSakeFpWh3ovKmmTzY7E03dS/e8SttMO3wKRKejmtIKWRuY4ISD
KAQCDeIgv1S+fKOvbn+Qg4yzM2e9I5q05ovODuCgMKIPJYarJMw2GWwWQb9dvANv
2Jd8rxbJoVg5I78An+yw7xuZLkeJvx9mahLvHXw7tscdj1ZPOUx2akX5drcV0m/l
mWKacmjhi1IZ8+LAycDvmRcVK6S+GQ+Ljdxs2pRduyEi8fIlyxHJzUodmFaMgQRB
tRSJTR66owBl9Xg0yQDPbHaRe7fjiDoN/L1BB0n2Gys7r2HydVt9H4dX7V6QdiFr
LooZlYISzmXViMr9KloHkb2wMMQKYfy5z1lWog9wYBP9UDMTtOa7g7VcpR9TmgnS
wsiLcvw5udUqJIEfxy8Y3GZNZhhad1VSkOX3WqjACGd9gaX+BDhZxT6eyzcd43Jk
QaX0E4M12gmRXc7r+baFoFupxJ6pb/LouEJtYG2ZfxfDcICRiAnhV2D9QxhFEKyy
XSS9CONYibhVB/j4rOXUhjYeFpWbHhG1hmexMi6QTA8chEmrpjuDz4ekoCzp+MiI
Zg4TWTL5zwJDYC28hENXH51REFL9I0WnxWXUuElC/XHEH91IdMUpQOESOoaXN8Jj
pqia4IhMIzkTizzYpMXLIVp1kPqjnLRRzmPjJ3p/pvWfvSwBsJetntecYE4u0SID
HPiQTbb7z1hb62vxSs9sxdOJ0HSA/1uJDTDZCMClRpG7v8YQwIiGlBAaDZBJxO1n
SAL6ulVHXMq2QYeyl7EcOrlCphxWIoFcLEpjSxG1xGS6fdf9zJGxiMxxawTQ80A5
SQUFh3gutt5B71xu4SIdY6pq6Z/ytNlNWDs/VUkNB4zYfblnc5CtzhcqUcc/IkFZ
7T9DPN4eN3HMkJWIwOyr3e1aHqnHiU2MKvK2DYswM402n91vrRgt0pupODuXOkMw
k6353CcH4UGUOZk0GhAEAukdEDyz9JY60s+IU1dUXLbb+4nK2HIVBu6fvbmIQZuU
XBvLGa2riNwDu0sGUE/gyDN9DyapVWrbLM6fc8Wgoyw99pbw8esZCG7iVCOnh/Nh
5uhLRfI7OOR+MIaloX5+9uXG3soP9/oyMtPhUUqk7aCKZZBkNYTxp1Zozwh8JLIl
72xGfCe5uh1w4p6Wf1JQqV4s5KFjFNMrO+fu51pmUL3XZRuB+NIvEn3iEcjnEDKb
zlPeD73L6P3WhQ7EWV4vUtZHmT0QeaXmk+8o8S+VtXHJlAjpdBsTdd6wa/Rfb4ub
0j1cF5mJKy7h77qRid7xn0NbeM7uP5UsiNgqk5hL7jdT2d+p9hcfB51Z1BoK+YHO
vT76b/e5tas022oeAonzx06QgJTE8XxJpuksoBMcbdC+vOBJ8wXLnUPdMmV8Qf3E
MHPnNLi9c2uuMXdCrYyJt6p5xbBtghkNdD0OAnwSkUPn/hKlhOzOxQVMuQ/RvykP
MQARZiSLx7Zjb20gmht6fz41wOfPc52rke85CRLcfhQIaOmapAys5II3ZiJ9yLeJ
u2VC8VZFAyiXERK/AU8ZXMHCO7YkoBMb6iAnUFm//M/z9AlPrwd34QhFJIYfsGKj
0UZnTrux4nHRW+0sQ/Ptv6/1wH2vFMj2RnbW1F+LctSKdSUP+xqgGJCafRGblhYy
oihqncH3/uwuXI/OwAeAD+m0GU7JQZ34837wVX5exC1s+YyLao4XvWtMaWhyzN5T
xi0DAhS23oa5rVCb5S0ZTBGArKB0qjStf6ziqfdPAHMSMD110lPCzjuUSKaIKv4D
Z+WmRR+Dccc91lhDpfuVlQw9Cx0cIbBivR/MZP/+AlG7krIZw54UvJ8sTAolB5MT
VXqABZDJR7sxuiisfX4Fz9P3i3sh0rwe0pREuOBfBVDpGvJGY+YtwQVK7jRESM2l
APlep4gftKSbAaKJ50XemRrqw+JcIns60/CUY/60fXLy4ohXKL/PIxwHqslYZOss
rQqj8xnMharUfmPK/rui39D/Uz3Q+8FqR/aP6VyVdmsxzgmfeRbntVvIPw2/9nEL
5AuMu6FFVrjwZ0n1IYNXDKhF6+zrS3kfKGIW6pAPSbg0GQJRHuxYKGczQfPnkqb4
DznrGEI/zNwlV0VqEk/J2aTCsTeVNDaVKqzfLrAd+jjnyR6rrAo+5/kPNwFrxqct
TqkZEsaHWg6JGnCbShBbpBjH7dNNfuxFd1BkZ6QLoeCnbM96OKxxPBm7nrseFSfg
NCb4Xw+N9WN9MEGyVCS+z2JbcfFbsdPXZ/sgizplyzcLj//aocEFEWrPZqfWgUFM
odrI+iPPgzW/AuJuWHDVXLJbs2gEnTEyBe+13nSSCVjhYvK+Vh8H737JOwuLeB9t
JNx6Zd4AmBUuVjB2XKNGj3MI5TCHcCQRKAanz3cYIHhAMwz8YJ3RrMK2BXHbw7eJ
FMEvQ3SnlDVTEa286MMjc1eT187JniaDp4ZPb5L5uR113HGlcludwaHzAXtivEce
AM6hhECLATdnLv167bcf4ASASQXh8IG1MpM+z9YSsQ7WO5ZUM5axCVe1E06hQk72
G267690FzvlDDGD9risD4hrqQZIH20MjyjgL8dY/+bV9j22Q7jgnDPAIyo7eJDS5
Zf0RTTJ3xuxyuo35F7rGirM9b8/0tcC/3uJoRgZhgqC9UlHE4Lm9BMDocQG4b2cH
wOxAdPw4pD/ilF1W9WjIlaIl51zjn5T3kzHXPR4x7tIvflK7wkpNnqmKLpLXI82R
r4kQfBJpgL2cnlK2EBS1x4g/OGwm7HlEzYFD/LNHUD7nx6G9V3rfCJwD7U0b8pHy
TNZ3gum2v9IcsoBtew/1b33vKZ/wj+XlmJQPTXcimA/XlPzDUvSE7N1OHEnNfMzb
PafSo4hrHGfGtihAs7cHgykD4jNlDB6AFAimanulivovX8oN2auuaN9283GcniNl
1IQDLY1jlJipZmJYHJF8ffvg3DNAHw9tBWXSb/e/abJcIklxMShFzJF9lJeLosGV
wKJdQmDIA9pyYeOljHyI+Pwh93vVJVMvgtMp9t9+4CUHDoCDqb88VZcN7fUvNp3u
eUCkantH4Emx3mgnkiztaMPOoVCQv8mXp09gFnTO+sz76Pa1d2C/fwFIvBijj6Ze
NVN469v15oU0ZGCHyg8+xOpDL0nIVd/OQekAvY0MeUcxlY7ihN8TGpIYfGAm5EvQ
T4VPeu6CNpysbAYZplyd8pedGn8LJs3iSVTrEh+DKN1Hfzf28wHisJR+7LcOg24p
zNDMkD00eOnXXb4pzX3ebhVXqXgD8WuGKrkpS82u+PHjdejSSyzTeTsZNfF+uZ8B
K9O3bgzUwBy46rSxaAPCQymg42h1qzK0pUTA6OL75My+Fd8CRim2O82Vy03sbJMx
7ZZc4TGAEs7hPbY3QkqZz0xQqLwh8EceQGv36IDiZ6bT3OTeqJT+IeNlsg2jKBfB
4SLa39edx83bwVTiJAtf9izR/3vVYuAdieWPiU2Hi4/qP7WXDnvBMAvSqashMulm
z+Jl96n/uCHayNsudZLYptupTnzTlJ38ilKGF2VpS0O/cLmmPDz9+5KWF/v6zXaK
IVgkWprsdw24H7ZFntjwMVLkXXB+dynD4ZjygcxF4T/+JhtX9nC9ChtKDCTlFrA7
TA4bErxMKqe9hYxg3oiTkj+VMEfar0xBJ0okYR8t4VfLCVnxj/4BlhjuCA+gpX1o
Mtz1x4JFlX//qfCRTEHOdqr0corebYp4qDN1H/0XdokmCmIx6xAoa5pdHJvtB1Mp
4fLt6PBuojnXcYNxWSTsAk67o6QCNTnLsOhkGWSCbkGMutTAcmRNLH59W3Mzb57Y
1thXeQ1nKdAecJBR646xVYWosCiM6G8LHx+aIHQRe210i+SUpJ7OroRK0ROqcZy/
AWZPVGC1fn83ydiyA2tcu1E39mCG149QOI0qMjsRXmhGzz3fDUFpnfkggFUhTo2g
4tWb6qayK8mnHsADsUWejSv/XlBDGsU/7jJjIKVukGDwQFEoJi6vuaCyRhaP/EHZ
G4UXiVxw3o6kZqCbcxeqcRjouRIdPEhn6RpZ+iKeWEIpFZS1li6bB3ar0HV+c4jx
mH3wgRrYHOhZDwRxeKHZR6VQicyiC89+AQEt124TEByW7PYNjxV8JKGhICDlAODw
qvxBU+6bKsDyJLKTy9PHNDMRk9iL9ik/6NpMZnoiny9GIfgO26W3SGJerGnLgJ10
dPZATMNLzeCBucK7RY2Hp8xbU7sHJcaDXTQ9N82L4FfziBd/lxUrx+zgJohxqUv9
6pPIATQ0oGxlCSPfR+buQyC+N5+SW3rrKImm23eCw0rP2zRjfxx4uU1qFrtCd/x+
k/Wc5bSL8fbIxL9eoPY/ScyunSKrbuPsPTXKxCiBtS/4t4vxghW8EV5OTNV+MWn7
nw9hIWOoiT5Hf4YksQ4/EYo0EMw59B9Un8lev2Bg9b/+wp2rxAnz9KBj4a86ITDC
hU4vEzMHesd0CuFUIzxmr00mXX4jjijih0X8rz8Ouzm9hN2nOPoQ8e6UP7cHOWA2
c9hNexxfDen7ElhOQOXWRxi4QeuhEULL0KZl/c6vxe2wCmmy3ashliZYLB+8EUe6
XSyjWu+JI3POVwBZU9M5/5dYWSU62CYL1R1hKDUNrAg48YDIkjkSGcyhPsEpj5fU
VvXvGSe2p9fJV9B0HxF7IdM5qL8gsQ3ibkv8rY3+MBBzDmqBPy+C6zUxz909RsnJ
y1R6qY2Fx+cybIZaqZHfwbfrRHUKluxmul+M1GzFIfIKi1HBX4OL7d+3aZ/al2b6
UK/hyMiC+ph+BstWwmERRLw1d6H2rs8N3cEYpltwaAFgB1Qo+CP2jrCVpzJHQaZc
SykPCO7WXiAJPy2RMudEYWi0BFB3vsKluhVYyLpI/jYxtnN2HjnxFIb6daV7iiOD
rU9QsPnQELYvLc1rzBGIUDbl4b8ZVn6cce6MXQMK+e7Xemb1DjJPBT7/ZoXhiitd
6I7xm4qf6RipVsZ53Cwli8uKmWaB5SYg0I27JQe/4FpkYHFknI90aOre4TpDHDGY
qudquFkrCjwk9gAitULnli8sMz7aZUuey2pTSjQZnXbaFwlAZ8dRXrfByFusGIph
0A1UVJ4DSFH954Y5YuSfeM0gd/43alPU8bJrKtErRob9U46i7FkfUflz+140LWhS
zcVHIKlMQBnKDifLAMqRGd/I/CVUwclB4u232KInj/Bu5bAQT7psRjZwd8p0O55O
fn8qcoU1rrnZrANMyB/3CwRUCeYj6vEicLsOz6Yj271xt11wa1mOQSr6+jRwUdR5
95r6QtFqBR/V+RF3aq2hQjHv7hek1OQtw+O6Y7l2cjQAW+PsvVM/wzedYliMjo0p
tizFGURtXPWXpoGPFYK6WFLn7I7RVYUGEAR8VL5RzCb21R9j95FF+nwfeKfP0FvS
//+0Y7aDiC56EoMG1KKNQNYqXiEVRx/mMUqDvKb5U/YMC0Py49ZuEzZtK3CJg30S
kjVx6Zspp+TEf+iFGd3ewLuHVdjIFykaTIG8pvne95OiwDDWoOabCuaTLdj9NIE3
u4wd6f8jc3rmmMsjkUneF2J9l8jka7xlEL3cfeUjktUT7GIBanYQ/Jp2Le34ExGA
OFhFUUnFuCiHQB1nykq6WVUN1j78dNWA4IpeHDOVQp3uEP/m28RhTRCVJ63vxr9N
x4/srvvB0JvojElxfXLkF9b1h2LFUkHWTTZ3wXB/0ORgjc4fzeC8USkaNABCsQpx
eA0mQJA+Ut4lzYnQyW0DktbBv2iLee+G62mB15Hgo29IUZdOCCsDoFBszCtFKgLc
aO60MnziWqT7l+rQczqDI27pHUPxHiU7ugH77SdQ3w69BJqsUjfhM6bKfmUIX3Si
9mIddk3vBRIBNP9m9Ws9IDEtjJoaZ4WT7zQv+4utnA5NGoHsG1swFCQtbR1PmTCa
DiuHUDzWnzi7EDqjTnmuwVToHr6lXSSY0atlqaHEblleBM2FY9U65G7zdvkR2eXj
KGGT3TyJu0x2c2vQweMCka4RhGb19EQMfG2t/n7gLxfBbUzun8WtH/qQd/DReLeR
IkZBskVac+mmaJGDZsLxs/TKGiqIJjIox+tL/cIb053HOKI6v1GkRTHDkSD1eDWA
lbaDWSFEGda7Zjo9E3sRTfpeRoXWXL1GTTpQ+pXwGUroul0igpK7xASz4HKhaq7a
IgQbr4VX3YibH7SFYBdhuNJng2zn3KR9J311buQ5e8dqB4uQ2HBEcnm7n2h4dkYO
frTuTQ5eRHqv7UyHVCM9SgGiaJMgw75CsPX8lWIKppz+v6Bzcc6R17tKyRzztJYf
PHers6wsft1PxRiqz8DWZlvEmXqvsGvTpDTusobjeJ9zfkjL5ttt9vDHUQKdyjSl
ZPTySuHfZ/ITc63+taghvT229/ZNDdlXcq+9BffLByMJM9s2QwBxxA+rpeYxMEPH
dt+CVcZX2ze4SyS5P5IZkeMC83Rz6ybjs75ePqXeRgn0nHyfvXe17FCTi3CkLuzN
347njp6YXC735BsCcDwlOREVgoaliF3tBaQr0ynEYUEb04Gj/WqNKAzGMsGfVpb7
S8VpLTTOypMECBbuBln7ubqlzghf9TJZdxy2TAePJEvhc6nzDiztIvKVOHn4P7vj
IQYS6IzM3UC5+fCKzzjWQcv0lbJecgGQxpmqTmc0wvJpJmohSCyModCOdhOQvLBh
LDu92zUVZwTme2VVERywIXsvQYrhaCnlAZcqwJC5PNhH9y6soi0h4HDnUc9a9KyE
zbwIa+0J9L68e8iPf8MnItnD6m5STY/nMAR4iBSO/I7Efcuil++/yw/GZIS1OqjH
l5LHamoYbiBycL2H9sSyvrd0NFQJkQpaTBGY+gkiYroSqJJAE0WxQYSljbIn5lty
1euYCPDT6ULHa/YxnMsjqbARUlU5eCzRL6YwpYIF6JypI4h/FfewCVpVgLOhYvlH
18AUyswuo3m1Epf1ZfWpLHrvX+F0Mt2ghCZn2czPpVYytnRe2E3wVmQuBZc+cd5Z
EN3CH+9VYalZECuoaaKJVnh1kOq2ZymZ4vohI/7+yRWZoPW5pVfrwr/atk9D9YA0
DtI4BBGQXe1+ELzRl+xPCucmLXKqyQYmpYJ+fPbbAaIpxnZmoNryqfa8SJEByn5V
mBUEcWzl0KLsB/Cub2uBRHeFeu3RQYCaW6eBCRzpnEU5qhpu0GkzCZH+6dYLiQ0T
0gHQLvQ5Cja+yx4sdJyeW3PODOcVTi53OPDTu32iJoJq2RzNYd4TQSWwa+tVOpnW
627PpdaSdqKlMpDXOf0QjIo49Xz5RQJdyyMM9Z0LP/OJUhVCaBxtIDku1IMZXT0S
CmncswMJYDmLW1H0PyEBNlSiXAtqMp3IdNAJHqEywavc9ull2eG+6Q78nyWCiA0G
o80Nxj3fGEfyDAkY4IiIB0IJX3Ei99BSOBz4D9s0y4hWcVDi0BDuqxRP3oZ+lPp3
Fd8G2+yUUVw1ef30/8TBHU1DDwaGZ9l5i262wJTnev/iR4JwFy0i9WSaF7y8mLwD
/gROQTxoelHe3bFRo9xrvc/SibQh7wvvIElxa7FfDaGcA8Q5tSaEbKJkf0UIOW3w
uikvThlF5XBuyAmjdBg4IWfrVYhyfYBCYVzXI+V32tvfZT4EuIntJqF8MbRCMxWW
TdSTKnGtHjpffmJFSluDeVxCT1rFgjF89NtZVka6MzTXlLjKdGNlRAQefSpdw6qP
7byK3SPTHhH2xJMng5vkpQ/7fFnBAvDkRd79BsN+YQAzLr2njNifNI7rCG4rkzht
djqcgmZLhY8F6PuGQUK0qlpIn1tOZ0FEv1hThMqFprEcP5YIvo0EIxtlZiClXQkv
acA5X+qrSrO5jMQJ1oza7F0zMYTfrxkT9z9UeiCqfKxchCC6UX0NEZEx+MZDCLqH
pehvmx2yNiPGpkEe9yncLMQ7lR44xh6UEzBUbT9ea250OpVIOeHvSGBcjA7fFg3B
N/fFlFgiOssKEl4lsZcpMzQ4B0WSTedTLL2YRKxt5NcdAYDxeAIXS6e50od+iJQr
n8q3WqIvWd+BJODbolK6CW6nj8GHrOBJalu8mYhL8Wvgb61Nz11r2AjyoiuTu5Rd
bMdhC1NhuXcAbTux7IDikMAHV++2+ZHkrL1yPJeXE6H756I+FJq0PSXXKQe/X2jt
UsbPWVRZRpigptw576oBHTdqJniVaxmRwhSK1QSg2qvFcgT5LtkH5V3MkFEwwxRb
QORsAcwHlgdsKpt2Jd/E7yTqpNtPys3uOoVHk/Mf8RY8zQpb1o0+dea8aTsPVXar
TkRnrmC74f8bXNG2E8z5ihmY1YyIO3+NxnQpMToBV/z2zYzHycUN4I70xCu/LtEd
tpdV5lF6y+VuQ1tet1Y250HhZWDn9FvO0MDUxnhm85XctNF6JeP9xYUSkG0CxYOF
bRTz9Bcob9zgqp64Sv/yqH8RnEN6H33lkJjXsZLqcbyVu4dLbwA/IF7WJqqXFliQ
u6L15Lk9UEu/+j7sjHN6IzhGezpqptpC4ci7k9qdMDB/sISfLFAppbKz9l7iebar
ZL4KkiVVw5TrwmN61p34FkVBXB1cwBmPizZzvSqxat3YV9TzWJlPmU03N2zsjnby
u270X3aZrgrT4Y1IAbrv1nk817VYbW39D+PeUjuVMYI0k+hJ/vVL4MsOySpC/Q3J
oZ0/nHn+rsi8cseqVLPtsMSNZpzSoa5TpsQAgb9LYM/YJ30Cjm3Tb7uNRIJEXNQ3
PXDMEzWOSEMO+tCof8tuLIoIuMn0VRQoEfTB48k6O30zEgcgPOTet7AJd6y7r/6y
zezQHeD7VQmNB+hlMEDd9JcVMywQuKBGA0ByJZTPXFkQo0KU3OJs3TI3VfIiwPjr
l/OJVJnnF3i0moFv90NC2fjwZ1amplyQr5P/lSlUqfxqPMtSzUuw6YRiqCI6WHyv
FJ1tejy3VD4zORVEJEK440gYZXIM8CwIIqhcv7lbxmQpotXGb+Hyhef+/LmBXhG+
bGQqtZgmk0EMn4i0JkGMdc5RyV6VjtzLq+ud1nR5Ts75XIF2PTBy0jjTop1W4mFG
09v06ghvfqHMHtaNMfuuIow1PnAM2hdu5oQHZhvY9fpYv2csqbT7gog1m3b9bn3P
LrSsL5hFKKOxtw8+oML2KyeJYvMhfgGBvv3F0hYoAJwq9qoEKhgClNyiTrpM/nGA
4I4576/4IGSXJ2L9Rh5OM1Xlx9ZQ8v9qUCpzEIUTjA59ZBPcxw37jnucXjEsBZ1k
w3IPR75SnKZXIrs+bIGJlNea+Oo5YkwSnCQgsCy1jGeJ3xUHyl94GkOhB+JtZ1o7
Z6a6n5KHgDf+GQKP13AdWKfJyjUNJtyO2Vd8uTT+2ZDnaJ0rLicGQE9aTxk0TT4+
SuWukCKV43U69B2Y7L1S4uN69aKzZw+Dt9yrGtzpaYt7OScVkYsknsHRzQhjGSTU
FfHqclzivrHhehZrBcIcwXOmIA0jBlb4WPUz0Vg/laiNdPNuF8f7+XU30mi0qjgn
Lp3GlWwwIEcAX3H8YTiABr3xICyXkN9MYAw7XXIQ6sk5s+xe3udVzogmBCNYFThE
3NPF8A7FCpuEmtl/cz1pUlsGieU68nwN+5ZWO4Nt/ErhpvAHlN62J8riN8PNA0an
gvbRH0B6/nGQI/n7wC/JbTDj/jg4Ste7BYCsSFobGhakFdaESaHlJKimnEClrXd5
Bsa3r6RczJ0NoEPaUNSdDiI2IgcMAx7IY/62K/Jx/pS448nktb9ZroaBrKllAyLt
MtTvGhn6j51q+xS1C5XeMNZ2BAqMnBtF47NLpuJ0pnuH93QkVdgCa3Ify2xuAdok
EnkJUoiyqZG9N09MoktQpFih4iLCgRkCbOKLD43kYVZwUAnT8nGI9kXQwz+yXqpq
0HAevq9rujXZyV8bJYAQN7TJMhQPYjs2bsflCTwIzs0RITPE7WT6otH5XNNRepRA
nNt2X4SbaG/4JiY1RrdYLxblYLjwX1h/3xChje3aklELZhOHgQMuzNQxvb4zwgK+
0YYwKJ0f0Z/oV8cJkfBpb8Dg+B27Z6kiw92Dv5uRxrktKxh+suD92heorTfBj3Bz
xUGFwVQNGby91CWTvWBoAvTDIfeCyxFD8Ksf96NBslWNh8k9tFnp1VYxQIWKmu8J
zvvo4jAiB4/nJyMyFRhJKehh/T0rA0kzyWH5cY5s1jk3FnGme9Gq/ltQaBGsKLb0
TP2+lMorvtbBmvkVo6W6NfiGisOA2nt50qrIrYNHrQBZZy4D92WdNtsEX5q4paE1
Rtkzij3zIf5wCvkwsQ+MOKet76oVEa++MjMQvUONOTz/B/YNw/dX3ExA0i9WOdof
B7M6Uq6gNrG8IG/p5XYM93JVoe4nz39zm61CGj1wNvFVUiVR8fpu3m80K9hre8Wk
vGBxTJU9OJduVoRItkNwEAYZnxzd5BGlcKUeYO4Wmd8hkiC1bA1QL6BeIgKdApj4
aVRewhoMjLKxzEeeG+IJQig6JV4HE16C9peMrvMQgQnT6G2+oqeOxDsGEkdqHRWM
IFsKlu/6cZnlk3hJdJXc3kz4ddOmUq18MD0jR3FHYIkl233Hf5uzlZ+NAAmHoFkN
2BpD4+s1SjpknP4IyKCKFfc3/UZCt3zT/T+OSnWF08wWQZCjEv+4EHn5y/YyXJ/B
NbHa05tOho+uQqCw+nxgDC/YJKnuBZ16Glmg9FwmKdf3DZRb8/VVQ+8kSwSk3keu
DBaVVKTjlvYdWp6kBd6h2PgWv9nG4ag4Qu8TrKGsq5QFncrLul6K4iLertAECuGd
Aq6mfrDLf5YY7MGcKbq2oAHPYfyJJySUMAOP5xBYZGFh9qJ32YYb0VudNFXmLULY
EyrdeJL4Q/PZfmrQaElp6JZsFaKeU6aIvB9hQVjJAKBHAW6qLSu2Fy2B/XlGhE9R
Nsb94RJcYA2UM2klgC6Pc4/hpYXwt1y1AHS4IGAUP6PhkqprjUBPNZlr1i99UOJO
ZWiYjQCkMILFsQ9Hu5PUymeeDSFKWplRc2qcBuimRC33/rcEUJaFSX5iUywNAH6g
lPIq4qz90B9NduRsVO2oRJF5MLSmqa+R0k8dkwexBsi+KaT+G5RXTHC3CYUq9TUW
f0oxJl1HZPmsRInZ5yab1YsaYBeAkcVCN6f7fBMGhtfwZ02rYDW+c576pzBpxk6O
pod5i7Nrt/OkBl6yfws5+Pwva1n9li7Du/LQhKTKnRs3YuC6TaK3QPkfRGUngfC3
dkr4CwxjzBs5FsBXwZ2otJUCo2p8MMGHpLUG7f2fy/s97+/8JxfmfVxF5yEduzad
o3TgaW+8ehAHK4dxc0guSOhgkIKmJDmsRBLTK4zn10CifXCy021fIwKZ0Zm4Kg5M
7NH7phwMwbHBnWJNy4hsb1/ohSh7UQkvvXRDm0cac7d/HFro/H61acYHeOItw2Ur
L+GYWebo5VhyIPUx8tSqcinFP2zu/eU+XTcbeWLgMnLNFwJxttfq++cV41gapXeP
3jLG7+NofLdaj5uNIIiH1u7MxqcIY/Qth7xv6ocuY035vqEhKDuWm3tnSCcBYM+W
KZY/oMU3I3fUH7Px1Qm7HHaMYX3RU8Qivj86thTB7GLWGaLtbmRoKWPU8E+0bSGj
89RVFIdgiIPplxU496mIeJ5qZkoThWI5zcvwNSRoUhU/AIX+gritdChdnzwK24Bt
0/eQpfDQXR4awnx6TIMIvywf7DvqOyogoTH+8vC98a5KFzfIsIhVr+ZU4fmvyBNn
OWpu5PCD0wlAr+vm+Imc0ul6q2ikEmgg6sDV+Fk7ZFszFbSYGZuIAi2CHuIwcDsD
n06r6hAt7u5fSVm814+usyP8BJg61KqvOl9bzvt1qf715WsaKBmWh4fGeZB+gjuN
6n+DmrNOO+Tl0wo22WUDribHyuQRWKQLeVVqHx9/9Lld37gqix8PhaCmUvZVAwa2
+zD+RiNmt9tCozKCA071P4r//ko6yCEtvr6e/bZR6gp6KbQoIULBdEfmEKR1fTUi
Kok2FM11o4+4oHk/xnlXtKq54mov6C6JxEguJvOYV3LO68HQZkcj9kA8uhbQTInY
jCuS3He5AROczHYnMWSLt7Fcto/Eg0g2FsTmdM5vJdgYXPV3qU/vd41PkqZEJHOk
oqXs4nQ21X0DD9osw+Ihb2KjYWLIAgDe1L65mSwLKWD0xIGomAJJoe6N7jendT2Y
spiGoMaZOT7rGOBLl/OpL87JVUWqaJukdVtfziasgB+BZtQ/F/qYITPc7ue5bV2d
TVnBPleryPMVhzHHewOpdY+9J8njbjCDZE3kbhdWBCSKu3N2W4KL4yB8/Pp8WZhR
9UAvHho1bxNRX6ex9RlGsoX2nRcQpXu4lnmpqnM8GFj+MCBOAhhEUm2/GUhKRhPo
dddCsZI4zN9Pbl1+XG7KbW04vgX+dqmV0lxM/cAuI5Jl8PbWKAtc5M29/Pe17aKk
JqzDHuIsMK4a8gXIRBBjZNpJ2TzV4e8yY8rlLI8BDPHoIL/Fn8UugczlAryogjMa
g6dzOO/ku9TBbz2/x1c/u1llz8VgeXFXx3TgZD4ZJwYg4jxWGmNp8T8Vn79f2TGW
5glqp3hYF3Wqvt5FiqIUcw4ugyw7ap+BmqX2dX3NYHsy5TvnO4aHGISwVp+BJ3xj
mWBrEJ3fgjuBHwePIgqXxZYzk0mptSALVbyUsiRdVGBFAufLBhJOvSW5i0SU1Ysi
/qBH2/z22mWm0zFzjsMdfnwz/bxHCoFsO5pf6y+uZgpDedWpcabhk6fO7dDg8J7u
HDvi6/JHo+yNvVyTWXsns3nTq+XHXAC4fo++MlWB2iKC+vJQDWrN1LUUehgz+19h
pTnCg67rSZ4/XOr3Oz2fUkkiFuJHxN/jKMHx1rBUZQIOWFMRuGE7HI1qZNcjyne7
BgCqJrwaZBRD4M7FSCkBELQM6/9h1fwE5FnxDS67efLfV1l90kJ4FpRzxFTziVXQ
mYMYg0E5yQTOdgk35KMhEOxX894M7PElHIARdstmqg1+suCrozAms5h4XkTNPmUJ
eY0xN/KflWaWgZuEWq8xElKFsruafHSxE96Le0CpyyC8QbPhiQF2hYVgMGB2FBIR
hTD+SV9ykzSDJ/mYT5TgJ7j8V2upntbKyWjY5GdWH0XSpYtAJ7PyY8cj+pvkh1Cl
Gm/hAqX+DEVd4PO9lb2z7pkoKTbJOyYrXinsaGU3c39JFdbs85XWE3/or9oz37Od
UIomzWNae2wmCRuUV12gP5N2j9YWbCQrOcb//hvA8OQFuPlvS/dnzSsNvoSF1tf8
wX1vk1nPFz8KU1xj1CKOGouyZ3Fs4z2QL3+uWFUPOFIgDWmSeXIl7pGOHng1S1Vv
0XZ2sfD73jatfjXW9YNoL0MoYj7Pdafqv7bmglPG6NUn9pRPgUpf/YKEs8EhJPVu
NfCjLyzDZspEcLDhM8GjWpidCUx83PHzA3h6fNtAPlquk5Wne6smz/ShKGaJ32+E
Z5ouPvExLyGquPD7QhcY3StP7Lcmt7S22FWgKzD00mUqNjN3hQcYU5Yq80jQ2cib
Yq+Po1DitI0EfJ7HRlGCIXN5Jj5xlP92JZziY5vDjjrDvXDs8XKHCqz3t+/8/dWM
0mijE0pRlfY3f9TWWh96FAlVW3H6FKqAizC3KZ68I5QSJQVB+QoG0yOSQVqKQNyO
XOSQiDEz8pRzknPrkPb6z8P6zqxbPJbIV2u7bYPZ6QaKBjXYr3vIxcKL+mvdJOa/
vxglKx4DJ0ZE9r+n0+8L9OJLWo2t/CJOZqdTED2vxwpbGGg8GNMoD00RsT0EFvef
foJJbds07jxBa+VAyVBZX6E3MjMx+Hp9mpwQR0UmdgRhTPwcyg3AjJwmaaUgiBBD
//brZSLtrArtT6R9dW6jp9ChBbkJ60SSMjvjq0N3GIO6XqSsLpR1IWkERe7pPKPA
2bzAKGg/Y9QGC3uljXdSUPXnSfoABDtmxH+FBJMdt0IrnPS9loBgPti7mPJq33BU
V1vuE6sU/IgMGWAjKCKISNp8uTlkEU70aHZTFTCgsjZ6PRgzjci5EYe5UlXV15OZ
dUmACDAW0L5CMErEB/0t0rkJPhDBHL8p0XBjjdwRoJThbJb4cH4nlhSa247RSwCj
Vdjm4PoRRDRdq2zheTH6k64KU7TV+RpNBLcR/MBNOQLHJK3wcX1ed4KtxhrP5EzW
o+a4t6LeX+CGrVyehV3O6Lf5dIo4snEJ0Bm0LLZ3wjJ0rDInF8oU6D75b2MNdIBE
YrpJcf3+xDiC+HBJFr2Fdq/cX8PIzSI/OykuvU5CSehcHoZnlkLE3LZtqvmGZfrl
zCxYJwrycHhkkkb1SkJ/zAE3r/KgZ6ZXuXD2oPXbuNWdQ4XAg9TyaXd9n664I/je
WD+l+h2NaUvuJyBUTQFQJzdvEIX75o8fOBV+rtEnUCDmPMADGeWXpnIWHYNUCiNf
nBc4OzIoPHazTJefpGymXjtyeCfsTYP/z5Zdx0rLS0ubWvYodaS7LJ65FoUSyNJB
s9PczPgCFXl3PLZQWPL/ftm9mEwVR9BOGSKmSN/pgo8qnq5njz1B5NbT1nK/QL+F
j5gMfRmuV84Mj9R/lMF7qEzjucVaGsn60rmCweT4vlmGl1wk8goxfhbc8Ya5u9ob
Q1UFsr1sbkkIhKIiqXZINfxVfWpAoGDlBFRLkjldS5Sqd9a0o7xDNI2AjY5HbYME
PAwOsErlt5vG8wr4ZVASSukcrkhThdBhzh+MSfulsfOuOuzZo6g8l6kRstEsllJ+
J/pqpi+A2yLvCbvRvHb3mRKTWWDvAm6QbxbzJH0bsqa0tJM/R1Ht7n05a2qaKXPO
k828HmwerSIrDMkYiK8u3UGeXRoMgKlXDZBtvhyaLKoKiDQKnYCZzgeEgwrU51+2
Nwe3hfvInA3RpTfqYNm5VyLJwgYQXXyZxgLDDVTTlswwiHHYjdAlF32qO6U0vjiL
M/YGh5yZQ+pJPTyXjjxdWMgP2Jk6tJQekLFsXztQxxPo6BkgaO8laroyUQe2/enD
QV6UkBCC1kCxpkatTigrG9Y4Fdy6Sp+gYHd1/0wY3NA1E2vKkjRKOOMmO2sbsLKx
AV10zwWmPTICW9ywuaJ1G6UIoqbRG5tuBZZ+oyavipUyI/YqD86pHeSekUgHaXNo
WuCnAIKAt2mEN5x2TAos+uqO77CATWS7hMVngZYpdkuG5DqTqjVPfEUiomEXXUVc
w7kfjamWWXNAmyJQtu1UalqW+GnslgQQ6Mb6kViEKDTBwOlEOe3UOXHs60O9K0Mb
jNcuUPuD18hEewx0zpr3qNAznNX9gg2Kf1lMyePenMU4r16D21lWmXjNMgjU6k5k
chZ5YCr5P/2K5QLXX75y5Sj3g75o8TL95JZIzP+12/F+Rr34HjMiHOBGMFkW9OmW
CYdB8NlMClWFeUZJsxjYylOvX/iWs58n+jRNAL0q1ot/8Y4MgY3mKzgNwjNX4wPF
JEQKTzNdTD1iynqcyWxX9untjzx8g980kGVUFlt+WtXyR7JqqACnPsB7jYNKvBaH
nv73ICrviBPkNt3w+ox2ZVn5qzKi0FLO3IlvQGJEDLDS/quJ7ShfbIRY34k3TQ05
N+oSalf3b30Sqi1f0Ut4PnHkelVqHkC1bA4i7+XEGjbHNbat1vvAcN/C3P8d4MDW
QyOrqrRVG1a8vr2n9ENZOi+H5c5EhLwp1GaafpPPRtofxTQXxULpS1PGkbT4AgX4
Gbo+lm+C76YXgMtoId5AsqUby1/G5ET5DwUiRX6H+YxIjkEP0uRNbWTGn1okcbaQ
z5JTJW7chESzRfsrLkNbOtSCpnBVFv00vBwU1UjVz3bjIWGGR711JmHztAcMB7y5
HgllDb88hzzcWzN5ovead8v2mKh70mgQqYdWIkLlO0Kn1Sk5ptfGUc4dKz9kQ5Nv
i5QFeWjpORxnFmtverT6zM9Hj3+/wrPHA93T4giWKB1HfrVvrYu3yHSlldpGwdIG
2ERWi+7ROW1a34yy2kZh4bYjT6QvZWpmX9vwlBVXJtcXE6mJ11YJ0sLaDYWjJHk2
SU/rSNIuJZrnBZL6lve+nCPJxBP/ebbUlejPOX51xSOV/3EalLrTD6CXexZjK3qR
oEmGxNt74ded6T1p2PoqLWkClat/a5XwsMGuevVP3V2qDgofH6H2bIXCHEEyfIW2
/pxsQZ9Me9GVUmUPJzsK4/iHbjGX5OxF9awE3u2iD8J3BjngEJ+o8Z54Vsx7XOmD
PJEFKS3EPt/nhFGlxZtItNQIedQ032taCU3WCASfQM/jL0Ifipz8qj3ZyhX65prT
C4mXpJ/0w/NyuwzAdF/dalGJz8GrxS+y32VVsURN84sORyKTLpfUZ5PgeK/V4goZ
qpa3pBon5sZ9+Ygv6w8gA/re6BExy7+fKTKv6emqDEVPOfNFyQ1NIdn11x1VbLcK
rDL346bxdMb/EYk3R0+Xv4wNNJEFGQJhooMyeeNmPFO5tS33tP8VlQs2kIY0jrx2
coNaT0rTLzfUjyJKpa3VzXNolVK1iQY3xgJEMv0TUddxl1NWgPjwzk8zkq+3ee9B
7jr6DNWy4mYwDwqlfCPg40M85+eCoIRMhRYEvA2HQ+zq4xgpuNbQRfa0PZM8PBh0
4MJ21Bzp2dlzxXlsBREtiPWqKdTzoPpqQazCbIxSDdk7XdHwF91k2M3TkyJFH8uK
uP79RP4zpq28E85JabATxl6B0vfSL22xwho8siwFLVBDrHOxjHMfne1ZeGZ1PkAB
2RPSQ7m6D6BwzGVBARd6p2BbjUXUwQxV8lMxmiQEUC95YLl2dXCrNw0kIZR7yK79
MRTzGSs8zyczk+QULkYtR9kMm29SHh2xZtIdlV9qF/lzK0DWo3vHtD4nLEAvb5tp
UCooA6sOoysLMF7+AdKSIACW4NON6kJyUrty2ut/t1YswyUTQRdNbHLhpC9x6PIN
AQPxiI7mhR0hFjGDZ9WtAh5DF6OklO8S0mA4ZfrG8PPj+9y+ZBcPx7VWvlk2Ht0w
6ktTKRGM6HnIKwDfSRw/7xNLbGe51223/IiI54gkNP9PjRFZ11Sf3FHwvCYAuWS6
YkDLx7SL/EjI/lOCeSUmUFsNoanvkQ2lA1ElkVcL6rj5AjbaHaTsGuKbIgM7qNdK
ikV8MAjqOx4RCfRi5v5YcOLhnsjAWURQr9BKF8LHzuhyWaqe38zZTGNerCTOhWsd
gxICqn37iCrskPjq3Yqb4F6vQUPiK4yvKwGmUhQxOQp7v2792tMb+jXmz5dLoo8c
ijNZkcfFnZSqKKZmyosm8b+527e2gL6yRHSI7mCBUHSXlIcht3+bsWOkCXWNk6kA
U2MQ6KUyYfp8TMj1EQOb1WZJ0sGpbU5St9UF9uSbbJ8BFyYJakVgMAdO05APXEn1
CXOTbfakifJv70rJt7QfXWiq7Z/vmOEd/k3LytZiclwNEr9BWK/Hqud92fmkEWra
Fo154SdSoyn0vjCgfNwtgmSHXPHIAbvIX1SSsHrujnwwo9TVlUZ+ZRCo1rzf3UY3
IRowQJ1xpuCFLu88lBHSknN+n8F783aHhydTMfTRHVN+p9hENeppggDKOb3hzbPN
Lq6TCZXDxSbDn17xvYcu/IqHBfzYKvBmD468Z/ipDovTpyS1S2BqZEfy5hDQkUDc
5QW3bxwFB0jVPNGkIPEwa7Zg+vECLZhl9OTprZTdB8N8fI8KJSbl9z2HVujL0xr+
QYgQoIPqNcZIJfouMVvKeKgrM0Zso88fvKIgyi5kt0gotW/xNzWpKKWvBTj/aqXh
G6IPldnQ6EHKvoAwxH7ULHoyx3zvyDmYPufPYPnpeVvcnCrgsq5WDFYIcjbF3Hz5
/uElUgPSnNmbAlxfxYrUqYseezBsxnJreppB7TUT+iSQZdZpAL25emMJraujEMcs
Z72l6+eM2s1NdOfeQtRprqb4wHRIqMTJGeiR7Fyz8zKPC8iod3cILejRP2yGNj3t
sIazNfBSh0ZMfbIdMv/OxQnRoo86UxtYZeHc/vKBtovPgXAUB/jyr69Ao3fEgsaG
JTCygyS73T3AozPN/94F7Kue+HqHanZ/K1SUzARZNhU12k+OqkXfiXOMuKzXXVzz
bSSoCG+jqaS1fERptv+bj1EsXiPiqVS8V8N37lQJIdWY3C2d96saouLwiI3dwbFt
NYI/oraXcs6Drmz2EEGgWZpGNaVWUiVslj+dUlt15TH3f5v7m+apELPmBVHjmwOL
oNbFgALQF62ryl21yE2B1xubdiSPNLFpfsOGV9PGzZlImHqkZrP8G1LAbDTFf58r
eGsr5WkexYRamhcVewjSeE3iMcKjkUISD5J9JuCv4DpvXsVDs/R2VOqehmmGCqL0
IMUS7T11Twy+5jrU6/ZRlIpysMp/whqo3Q+dQhK3nSn51317Qlr7D+pSHTVjnzrf
oRJbftqJYWoxSMWP/jX5InRN2m1pL2uduZbuAcS/UM9R5KOVRzmt0gramFuEUKbX
wD1d/W9kN5wDnT1I+/myXYYx5Qm5Ci/YSSutCi28YnNmsjj+ET4L5qcDSn3Z4IDh
c1+xZ6XjLF40i1qrQhmoe0lXjP91YnjrzM4K0DHjaR3JZTSwKuRPsekGt0OML2z6
Z4KHk0RcZn8w0Pok3DkHlmQNq9yRz1XkPnNXeOh1QTnla319RCtycGSUMUej+iSH
ymjxVsa31b100tEtcWkxuhBn2kalpjAt/91SeFvszFMTNElOrqokg6vJpGwd5Dkj
+EG+bQbX86fuGSuy026X81fHJ3cdXToEjSgDWWNgLGS69Gm23qMb4acmJRrv9mjw
5KqS0yGMkewJxwgN5P4QP0aqssP8Iixl4qUDilCmu2D7FP/7+sjvjcE7fYKVV5DL
z3XpQBgdfIHaS/zl8vRFY7W2TMcrGHIll+xHXvLVDOqSDHvMnMlnNPP4STZUVX/F
Pcm2WkbK7t492lnD2ITdWhnVi76lV/DrWknKVivC1/gL4u07fGNPZ8x/c1CVQcL2
QOrySKU7ICMzx5RSUGB7lgXGlTDr37ARBlv7uvLBrq48BT17Mv/Qk9iIzQYT/2Ue
XdnrsNUv20QSZt5uNIc6/1P95jfm1Wsj0+ljsPASPdjLdC0m+ObdSxedRSDMQoWW
kT8s1AWbWOWccea0lWj1WOUQm0FaA/jTTto1mxnl3Dp8+AUW7kjp+JvfQCqzYoPI
bgbllaQz9lIEgpI9jB3Ko1iejpeRcEO2qhul7Ygm5CY9ZkDPGmhbS5fUIqeFGGxD
l2/i6Q+42SK4qF7qoT7m+DSn3KTB/Q/zrY/S6PRoWqMmxVT2BpdSzAwwwzI58Il5
av/3w24O+Aw/axAuzp+JQODZZdLJ/whMdMA9pFFzjn0FWuXiTj55/kY0s811HfY7
15YEkil8QYCPU2byZE4uf6ahuq6gjKXaMBVQVZVhXZ7imhZGIHs3LR6bUUS8WtDD
duBZBs9cj/HZCC0cZ1hlU9eDq/v46bAeT6stKe7y0XbozFhJPYw6Ybk5GmCBVyPY
4eL+I2bTmBxJNkE8xaC1eHL8ECQp9YIceaKr753khg+RrS846dtxFkZanINGiZ68
e8fydZ/trpEkTLQTocLZ54jVfzPC7pkJqxF1Wm/4DpIl+eqkyHE2G4UNkPCpFxVA
Zuzhi8B1BJTTvMTI7Rfi3cftErFGnrO5RkNr1eUs9gs6lyqA3UWSw5KS51HWzZ82
Jw5TgzMbQwGhh6NaH+yaqyHhHPNbA1hD34zytkJhFF0pS4hmF22p2CkhPi8YPSPJ
IPRI/C5Nr+PvSBgEHnRWsHfh5WAc0BoHQaOls/HbXcU8wriDPpqMriQeQ2ijKupB
FEO2srpdT5weTkCzDshXcYrssvHfLjI7Al7448ls5wa+4Oh/zCiiGdemlL29VSK2
+sFbZX5kf0XHzLikBrIXbzP75V2YowbcOWpcjg3IPdoOwirLI0GwmhREieLG8uk6
ReKtcfBr/QFezyN0IbXqX+wp6NWbHDR+al90CiUThE3dBWQtsPpox96LEdnoJbtf
xoKqH5u7OY1rS7QExynVzxQr1hXaLtxYx3BB29+EnhWLe4STrg7RLWQ2jR4d7TUk
lpzyCsS1phP502ondO7AwH3Lo8tVjwLkxx9RVda+m7dMegg7JQLCInF3jPcQaBYv
S8iTaJvxZy2cf+qh6uWekDgBCL8vgAl9ODakdmBznCMP+v9ODQ09qIKtBsKNtwFK
ijHHE2laylPpPBcsZnTgdVyJQT5uv/hEFcj0ERn4UFzqz/VjZvqLpIz6CNL+7hF6
WfLA7e5PBE8rgSsMvGq5lEk9Q+5JB0Gn1BrMiC/OfUHRzRKl0Z/6gFwBsnoEjm4Z
JSa4yIFUpnjdaH3/voBRjCnz1QWzy/Tp//tmJj8jpON5GK3OcoG26SGK6UY/Xx4L
qZM8IONWknnSVqE4qZgPGAnF7/OPMdg65K/rUFD6ucHzcN0zkFspi2NB3wnZksmv
Ume4ozWuCPN3DEveEKhODq1aOkVdvuoospul317ynEpKdpzNlYDV34ZUXNrLjhOb
uHJa8UzOmDonTgcdqVRIb3WU4PgP9nbG2oFZD0ukF3lWceOB7rg2i1XpHx25aMqI
z1WL9tORKCdivJN3jaIUGWnpPZDBbi4rGKhSAfABQsnsxKabDe4MI5VTBjUhoQFL
3ZrR3VjFi6BogSLfkWlA/6x2FQU+u1EZzMIn8pQM6+ly9ahvCwJeYvjCPnj0qrTx
x+esOyqBl9q3m+wXtzyF9tLlqLjwke+7O9oLzcvICHUumbRa2QUyAxEG2TFxUtU1
yiEzcJaJFgFfeun09aDkSddUv9nX08N3e6wnI/D5zEP9f5lV4sRuxoQg5Y4hZH37
yr4h1gQ0UZrXmTXCPoaRWkKWVE5CS8C5LIE4fqTvN92RiFiFC+/pzNjLjoN94I4K
1N2nCjhIQZw3BgsvN3cV2FeXEXW/Jn1tR0p3SHgcPv/AZoKodbmujfzjiwCGb2Tc
h8qI1B6R1FbGXt1TcWAfQA9PElk7aEjuh+rMtxaLpMu+TYkDUxqY1w0ttTU/Xs6a
+OplAKZCMtHq7/Yy7ZwuhfMTNaTJ4URaBVxNRKN7/Ie/lW54W4dkmx1YjORV+NJ9
NqbpJo2a+9t0LIF/oAKeckWX53LD5TGEZDbFTJ3tz2LBfuqm7i8Ukq36g4SMZXia
S8T1nx1Lac8RcEAmXITWyHObFwUcTdwaFfCJWIvqoDc5zgT1jvY+s7NZguG4td17
eTzT0EivJFdOxIC3HuGGhr9Ymuq4kuZJ3C4O8np0XyBZP6aVIRlfbyHIUu7Pyo3B
hwUA7JvBLofKlg9GQaJMst8PZRRUgRYsRPbVhshwXcrJC2iApMPwRO2ZvCLu2cv9
Np/zr2nQ6Hj+w9qJCQYtr3bz20UJqsqE93DTEQN0BLNHR41G8DQ1stpgA2Z8gF9u
CqVSwcokokn7M6t/EQSiROorAEzkmqQmAWRSZz8QaUxFSzmMb2dr0dQLwbIcChzG
IH26IN2A5nrTeJ+/54tlbo9sn9UjDZMZ8wDfW/QaXNgHRekga+H4+Ffje7fLi69N
JFnvrsOXD/R6U76xOVhv5WdT/tuz/37Q3Nth2JPwHwZAGKt0l8EdkpUsfKUeCACy
Ou5q5t7VoF0hoRdlU0MfljTBYtI/mZvZhYRPdcMjs/Clw4RZmVLM+MUhj6JZiaUQ
viSxZu3Ohq3apPxsz4igxTDx+ielasHJDNYNoOPGeAJuJJyuivpPfeQtidgSNtPD
xDmioKWwjL2XCLIAcsSw5S9TPN0AquEUCPUBimDvcHXCu7pQ8vOfm6XTrgmBVWWN
OIaDLhJyX0Nka7VzeDhVtSbpf+5UPKped/0brzJ03hzQSebjbHYLgoAL5QIzo6BX
kWpKsThZmBq/eLscFlrd/xkz43MmxqJagPj+3RleFvVVXLaKe+ZrcLozVtGfpDdB
4XiA+Rq28Y1ITnoo5bdsFneJc9zK3JHCqKFEiOF3/GIeVXNyrq8QDE8obpxaOduF
Q6MNo1E7ha4hfs+Isjl2LecMyfjN2eFBXqLGxCYzVEzoQXnF+Gfksyg/mEnXtojl
gsZzpSLRqycgatYtXPJZ1hiPZqFd1Qsao4cbwxVk1oaIeC2B8hNBe4xAoGSS0aPp
EI9Ik1fkDCrOZ81AQ8Z9KjAe/CLH2OU3FRr1+0JrIL7BOMcSo0BN/js3/w3NSiwb
MLf/7DCdyMgqqFrCwwX1W/MFJdLmvQ/Nb+2uX1xX0RvrpDbM/UK6s02tGQyCoSJb
IQQU3cionF8TE5S338jV7gdiGbpXJpnBVkBxI6TOCJayYYc8UgAI/unxa5iCI1rH
hJiNjXP8287uxvw4YxI2h4QBicXQSbUlxUZu/DVQPc1cQDImXIinieadPCHUjhOl
1OWTq1DNTvUHDHMuEk7ieloltJcUZtXqEUSRHhrHu+i8wa5lzNZ/yNz3bF2GqiBR
r6CTDiSayMtNnwWE77Qh1YYyQe7coR8z09J5decD4CiB0awgJ2/y+qaV994V607n
B2UQuEMlyEs/k3qZxf8Gkkk81e6XZ4D4MgVXwe9Fi6MApJ36/ylcKG4/OuL62POR
ti3J9XxnrMh8TuqvVEbHRIL+lK/IU/Trs44KXOxpZLrfWvgIdoVfK51U4N3p3n2v
KtNA6yL80Sf5tBmrBu8pf3uwQGZlTrpBcwZGrwTc8RCWg9X8UWNQlMc8A5KTK8lp
/EfWOzLllmdDPDIOEwndeRFGcH+18dMgULROA/0joaZlWWRGhJTvG3TvSq4XHw+S
QA/RV9Y7YWtdRX3zDF4DYsHWkBH79HRDlYKPeve2N5q25i2YgZGAT5stDDFmTpIH
4zfPf+/pQnUWyRKks5X1nSVBNbsfaDKbhTKBAVw9v2e+MBDmrYNxWk2Ws+nNvhxh
KsZKUUgOeZdJFOs3uNoENw1tIP2wmABLW1m7FbNM2uv+CV6ttdAITojzTVQ6x88+
803DCK/y9/s+SH+3PeC1vHc7Sii6gmKKx8soHaUwPgX48aRO+LhZwLkADUIL/ROd
biWl4Z9LsOKlRsb9K0tSXI4hv+rFItDDlMVxqMCFPVRXerArg3Pwj2FIKs6WFF5L
n/Aa6c0pw4USCejuXAtG1Sk5qfSjRVKCfJrx1L8FaTsHgZCF1wZm9ugxLyPw/EIs
XaFzYXm4ZV15vP7o9uYQgoMxnwKmRrEeg2AOHbpFStruPdQ+aKTq9f4o3e9+Hq1P
IBzsL9IHHPeAw15M2afPnYwJOxEDSwVVmmH2OFd0jlZ7zPTM1Ih65s8F2luug8RR
SazcSBvUary4iqaxWC21ZcVbpW0+HAUs4T8iq60TAzfMICC5N0AaDccVqBloO3nQ
/6uMyrEdAoit3CCtSGJ35XUbYJEemkz6u5wpCZem3Lnymk1j15HtX7Lr82JwSmWz
Kbk/Sv2it1i+5fotoaeYf2qn0AVLc0SW+Lz9jQ3Ujg3MS6G4BKl8ofTe8A3drKYI
E3gW5R/LPUZ/Wz4kmyRF1j31MjJCreHKw2rpJCi8hCllqoUhn1TZWxzqd3usAzR4
YNyKtMt77cUqPD7p1h60i29YMQ78i+1qae/ahvHLuV2o3Nvgey61gabZ6Kl3B2VA
bYbY3fsfKyqBrVGSPahp1m9O5BldPzV3Lx8HIGXXbuTYxZkBK1KT54p/HxcVsYKv
oGx2NdQXYk62P4d4EBKd/JZt0EcJuSqqBr9kpj120bQ3uJO94pbVfECozggOhqjK
VXKKgtINssRy34qZs+i0v8WekHJqaBuffrxXAqzT0rBkvzXTAI6Gr3x+2tMCOG/k
u6BlD29wT+dAeNpZY5v4MgzSfJgXw+81xJ+93S2Wwa6/pW6jNmhl1grDwKpZu8YX
RwSvtV0U+RXD8mO/ldCXKbUMBF5hE+vKNefpqL/AuPAmFKkY3+t+UtReU0kNus+Y
Pkg8nbvuCraqP2sWMh+BSCA+sdWMaHOlwq+N/exzi3bagqkd1aebz3IiGCnPl2fe
wiFaHpEbEq/1dNs7Knw6LnSmQzVUXieW1usbwFbVqvTMZhGLEejrGbZcb3n+/Bs/
4sisageXKOFNTaWkiR/ehq8JaLB66PQdG3OjQx0HMBs39zRKCdEPTt7e+ZbW/nVl
wXzYMEBwJQJS6MnKRBj0wRVXk0FCjhFt5iqnc8T9nfltzyz3osfOHmnauryad2S1
mDNF119+cJNIwNyubAc1ThX/aaQp7YXoI8pJLXzP6iiIU7qHBev+Bry4q/5LOE6z
6IUISGVxSNfmqjvGSbZ+7eN2k56gQZ7M9cvd5/PutN9VM7Oys211Pe8Tux1RIxAg
elpWTp6sFzFVdd6bh3P5n1HuPZ6zICvUDrVXpK9AQIan8D/UTp1H5irA8Mdz8ohh
O4OE2fScUQR2yz1IHrcULPUSAlj9aVldaR1XoL+T5ss6VVMxvwPMLmVyJR6XLmWb
r1pA/LVg+OG1aazrqrD+AizaLFTZKgz74Iavq8xD/tHvTkhDoCeEgLhr07gfBV6u
4Ym95VwTsutyhv1b8viTeqIkzTxsMa2IgProm1f/2fk5FYG0di4705IFZMvoev0p
/yJ3rLAXvOSHD+AoBpu5eBMynOoBpekw4XKlncFB4hNAwWAB7//2ygcQl1ED/jkY
sJ3stuFiNkRmZkDsdJSQX5hLVOb8Z5OCSuIDK9PT9B11g4QoU99PFAriiZY5G66Q
G9rRds4DiZUHeyPCrZW89nEdP6H2BcIlO++AyMgWCsIUsKZtxz/K0iJi7eg4Pdkm
edCipfQIMpo7MJxYX9aHewxsfdsrZIyaJGdmDgbeWWvJBNyIPkPHW/EVvVPqrO2X
ITP91RY5zJ2e+izm1KlMRvs+Nwa2eDcCetdP6RtHMRzsEXaAVX+Tr4cA8XqmD5W8
Vbzg347hcN/9VZM9bcYXeCWmR4cEIDxskeiL+eaiAR2oIlPnrfXOTwTFpoBg4vm3
/X7VYTKSA7t7/S0U5OGvIQ79+R2obb331nReyAOu3VucZlgaYM2NMXpKKWkGd18f
6JK/ozo2mxnMcQTY0+5GHHv7i69pdyz8Q+4JnjFkjC/373jj8ZdedkfTXBgf7Qp4
F6YHi/8JhuRV+8vwob64EHTsxzgs5H7jb+5ETPbb1ccNoDH6cdq4IZxj4SdbCxZE
fzwkDRXxk7kSFPTE6C2P11tfKRE2Yi9yFSifVVCrZSAbu+xVzG32LrNIdjxY+xM/
+Ez8JUZbjVso80NhEhBtngpPxq+SBhm64jjAKJdoTrIyG2QCz+qNRoI4oni3HzAe
Xafv7t+pvD03q37FqnavvRq/bPp8+KNqdRzM43i0cEJYkSpK4rLFDVwraQSiQ5tU
ea7g/QS56VVHuxxv8davgRSZmvz/3K6UZVvsxNZOi1ltJV+FZtZqKqzGipraFH1K
8n8U+PLHJbzwV1iDLzVY+/Bygi/qZDGvxLeRMep2rgi8MzSuufYUoBzEMTjkAa3d
lJY/pGJmdtXYPP/TkYRxcBa4jcRi983iZnAt5YuL5VAJN6cKPdKISFWsELDdaVX9
iAE3h6RETkB4Upkb3BbCskSnrv2iyvHCF6HWjNfKHI5xPRvPKtBmQRtwqJVLDk2q
TidkQNmBKvUfQfYiLswYiMm+rlUucLQrVf2vItFek3XZ6KcBiQ7EsK7OC8xwG/Kp
eZPV90HdtglJ7ezXj6e8p6SENJF/bdTzhwTqqKzRTiab6vwXPFRUz1NeGC9qD8hd
ceDSnleDX4pVKnDbh0TMrnUdmczTIZNmqUmKOG2nY+Biv0oAmKrkzQ22LjQQNEBU
gxEtVyVCP0EHFZn/8RZXtytva1eUycfuKzwLXTqU3R/fu9NCmzG9ZbqPPwJHjxSJ
hxBJJCGajdV/OaCpDXNNc8qmTzUqGUgz0Bh2aEKutA6bgh/u/EX+IGn8Qcwclll1
PLC18zlO/95O5gn0xOarnDlmyBtDUY/GLfuYkkeXySkAxJGEfLF5eKy2EUIcTitx
Nb+Af/D19teNwOk3g4n6DQ69nqZuux3RbuiObDcngqdHqbI9fBFNlOmh06FT46FJ
sLUTLkfRFLeN8ixykGr1RRTq9o63AMRrRmf1ZXrOHR+qaI7IIKilTDYppa9AjiLQ
zx6Ux3tx/zTUE5z7SH2SpNTzOMKmZj1sXb+AjxqhwrSm2QYtKqOfjE5gnS5qWCTM
HqgBcgKw0y7TL97bcfn+BEAa6LAGay4DW4Ts2lUXPNJOmBeMi9oql7pD9v9MPg5Q
fMS+g0Otd2ZN19uKnJLVpg0CrTVGXCET/wpUwf1vfheYY1Z1zRXZWKlVMqTnWXfs
3vkA0fQWQ0vgot/meXLKJONcc/nnk7rHv9umQQxx5BPCoLMPp6nDR7H7d0j/h3cb
Tn3AR/i9dngHRIeZqD8UvaIzvJWj/79X+7wV7fTUFrzE5h6rSXxpdj2y43vSN45j
6XHttackijA1WGX+AxICxH1WpsnwLsuwa08qVoq+wK28MAmitZXriAW1eN/UQnkk
4od3Mow81V08IS8DxPjcXcVIDTA2vZyVDPtj4RMqwuqg78cd4Jmvxbtmq/pY5NNR
U9jp0UJSpeuF5E3laWvFJ1xMFkKRXylxoGfYhSMwRCKkKmL6iliBlGEHEfgozTBS
CxgeYy9ycuHOxiuKp4BMqAMirgzeezKFW1G7Rwv41YpXVUa5K1vr0pgORg7b0pcP
wybac54TtsG14bgyDLJ9GVbvAyqXQUYPnDNqK3Za6GFQTQnXQu9M1gc4QWuCG0Qa
R26uBh0fnwu3ewkeI+qSNQf9b7TwBEcvosxnK704pwiI0slfhJz86cPrGzkC16XP
7uFvMKVz7Tr9WeVlCiRnW/eBQCeqMn2oAbEWWxPq17CQvBnfnoSqUH/KRGWilUzS
dXHZqyBD8+W3v8jDMntu4iCInWFACxR8z/wTElCGi3WHZ99quB1a7JHvalkiVOIj
9QKqlg0z/MBIpF+t6Q6BUgPMSklP1XXXPbd+yZ4YbzYe8ZMVQpCgnav4Pkbp0g88
ukNQn+TSKjuSruEc/VR+npr/z2FajRdX8fqFE5Fua8F4VR2VX7vvASu3vKBxGcSi
RVhbCBV8td9t2FZCeUyMx6bTTRxR7wxVxFz99xVNy2PYw7hqiog0iYm24uFdLRHx
p3F3dCNrEeFN1yIXsl9zf5yo1MjQZPs9Whf3KEyz2wa9rzncI5W5iFAXbbQ6Sb9z
IR79FvMRoJxzdEmFHke9V814gJW5YkfMEpoigJG3EgREQEIjempbewo5vQb8VQyx
ZDZF+iNYVZXjgJYsFFtJ6ETh+MrzOwfX6EYkkD5zQWNyujut+MIlTwbB3EJq6x5B
FOQxusV60tMnxCSNl6YupEg/q0pTUlReGVBBqd74Fxs5wOtE/8kQ5mXdkzQGLBt2
sW0e3MuKxmtorepSTGIAz4msbk2gciAqboeJsU9WW+aXwNFZA+Psiz3tZllxmMpw
vADbwStLv0l9MrEI3uAf9EXrlRtuP4Nu8nzqQur2wCWV81R5d/Rg6l4OiPNMiL3x
Y7iroKWiFC+15DEXarsYtXBLx+7VDlVm71ktCCCR2J0XANGmsw3UskrsyvLsPamR
QDD9oi71qlC6TaTPNVmdf93ftVKd2Uoj12Qy/71Wgr1Ezd06vbnCuyiwCaEr5chx
D7B0lwAPwsiKoMPaRta5bipE4Dm/SBV/iCkbrWOdZEK5N9Rnillc+G+eJRkUUvrQ
5m7+0HDYRBZ2Q2eqc9rGff+06+/Se9ZvTAsztUS/JjpR4n1chnPHDyD8vcHN5WIw
cAwO++2Ksi8jcLkAugOvHfAT9QLPIyYm+IZzAclN7rqm3RBegaMt1X41sBQmkjJ0
/a82ii75gt22zVTJ1mlbobY5tWzmldaPUoZ64bvtb7hwERwC3kJZXAoe0DEOOE01
ef+MoU9C6dFSIhk3QDGnJHDqfZLx4BGjjRQFRClZZWonRYFXpCjwSX3iM4xEQii1
02awxKmxEMp6/TZ3qlXMKUUVkga/11tykw//1tjRq3ihCV5MQnhTvszZFHb/jzc5
yWvtXBg/JJJDf2Oy1rgBSTO55QvQouasWQh8q4UQyRoN2x4B4arUfBfm8/7CJGax
BgrE3ToYz0Ckba4uYn45EXFKXk8mda0NgPsASnc+6JXEhXgNj/xK8KfXxrkdVIyu
5In5gqvFbMyvii/Kdq/jOUrPwY+z3l7gdlvqEra3KvLDcNcdMa7QwJrKOWYSevae
TD6/yTfldxsZ8EJgrIJIGAjM4DJC1GQTHmTUj7o4rLsTZ4DCanHtOUGAbYCpnMHm
0sGnTFjQMM2ePbmlx/PSU0lMYCGh5fjvWjX9NZFjZcBjHcL8O9bzEs1ymH3OazI7
bRch/bqmXC7ne28HjTA2IzvVrK4BlID+n6efALao3sa6eb5Gw8DKeJrm28hR+Mh8
TO05GxvmwbkYzycsE/Hjp/mb8hhd+J9QR6FFZkzQhcgqvnlxtRFLPyuhPz30RQYF
EctHqfk0u8mkVgi1K2rUGl8QmEUm/nAsJjHSKDLSNGGG6edDkmosvkCkSfpRFFTg
UycmNeHA+ph14zg0GB7bNL+sFzg0HcKlw3qaUBtO+YdhVwNr/f72EIwy1bIFqu4v
RCrJE65mJceQCFI5NJ4jdtkCIFHuki5pNTwOqumvgIAIqoVdmcnDDnhJ0487+yuA
T3hB0ds+WVRi681u4kQY7gqsijo+k4feV6tmUKSGW75Fz28PYKCMxgdCRZB36Yjg
V845+tCoOOs5kERdJlA0aKSBXOCn61BB5uH13zE2YJa4PAc5TJvxa1UsRLlbKMGh
qqr2XTVMPqejt+3GI/QgfadpJCEXf+wdfds83UI8780YPmma8W//47OTqOZnJlwz
EE7piyr4kEKXfP+resY1Nu6fuSaO7wPniMHP9EyPkGvkj4oVALNcIcr+igY1E8lD
DTtFBumVRWxvEx6mk3BHsBz741NBkm66y39ImK7KzvDORY633Di6/GGvJqqiUbHp
21M0sMq8oyTJngQpchjpBW2tTANkXoa8iJduV4l76JUQBdTru7qEUOdJQeqPc6Mb
OgRCugqCvkrwl09dagMSBC717ec2YxoiHNnXHvpQeUqvOnC0lCYd3n3e5LWN1b8b
bz2jHyvRe9HxgfWCOAkJdwaoHlA0vG80st+feE4fmOlhkUf3WGwHdq8npeOJEo/L
aZ3YHISE7Xmv6d88nIUQChGXcH6cMMofpvjFek1OQm6pJmo4ShzX5zJKXaqtvyg5
7EdLbX0GGYghZdisxnCeLJ4+tazfPlaOk0IAjvpSdDJPfhKoBn5CS/ja+fIFSzeF
iXYwZjm2csUESfHpSPcshECXLJS9YIBlpXy/r3MHUj6adZuJSZSz87I7EWnbgQYl
HpbtQQMbJICXQpLmFi0Jd2AS50eZJNFBR/R017fmOsUaYJ5JVeVmZTq28KB9l327
oI4/diW/8EHCN3eWnYFOE6Vq8gDNwM/GCq2Jd05qA6m7s29vPTGaZdOyQeUk3lE7
eg0FnKAQULUeKxrq1OPIHGBLjNDqviukijWMpRM+XJrheN8Ng+6bjYDAW8u1dw4W
h0v8yi/lhmbxTlzAFhn2+NBc6xbXZ6sefvyou88B/Z10C7uYk2ks8v2YALl9o/Nj
+xUumZC0LxFfK+NNFL+4ej3GFrM+Z3eByVK7ezhW+lluMK3yDvq0USl808vNTUU1
uNHPmOBAz5W60avZQwLnhcbYG2BbQi8MV5a2/lqZekY0UT1Shk4T9bwWtmsHKxjD
i0rHZT4rrylhiWC9aQlLufAG9QAliHBhXGZYM3hFpic95KqIPOmv/c88bIYAm/63
bA6h79zL0sx3mRPa3dHuMSMIvWj5VGVaRGA0bo2jKzp7axFg0RSlY5vLY5K8/1uq
kQdV1GBxZlA81S40+FOQwLWsPqge+WNGdjE5XQs7xMKTAqLGVKh1PpHGe2h1fAmb
4c7XfBWi/T0GCyZZuVz1MIlqNGhV7VAJ5gJv/CQAh66U/sUW92h6MGOawyC/C6Iv
UXmFM9kdozo8gbvOa433V9LSobQHUhNeu/IlE0kr2K+1Bn+982HUN5xFn4UFFPE0
LobCNn/HbXZZSrfCKsIcBhc+xvJj2vF3bEB/OAmb9Kglt1VMARR0LJQXln/0jdAE
y9qBcNerCLMKRPwq7FvuRcbkGahog0wHtoM6e30gbISFyrzzk9swEn/u3+1at7ng
I0m4Pk8j58ZZo7jiuBRjRoSMnjCNayA0AhCKx4TUo6RnoDrWr5+QGcMvUmW2Cy9s
960R4SN+uFnwqp0CI+M2rfI84ABZAACQUbZbMtzDhCKWrnZNN1r6sH+W78yJqyhe
ckJlknl4a4YOc/mHq4HSghVaDsJAFJ8za32ViXVKdgbvAIBkv3SM4w/w/j2EwHhR
VTwSCegztClP41i2IO2pnNFb4z9FtpHTc9ZCcEW6ZoDjhzX0bp8Ifmcy9kekD9Xd
tXXqsN4fmgHDkPfv/nm0JIePsLJ75DwwDvpistgfcEv/UOo/B1o0YK8/IXO2skxt
1aCPO0CnbrbCVcmwvQaPo73BP+lY4wE7Q8eBDEOx0amxiqGfuV8sFRaVw8PB42MD
QZ1m81toQqg0l0c9C3Dfaw+4BWb+5S1vf9P0Who8FGvdpg6YMjZsdA1bmj6bReTL
nX9aT6/Bgu9En/3iUXL75mgzJwPzuJey84JPugEdHpZcTW74lKNmgdF4F7grmUI9
SgGMBG3E0jOrnqpf/L0GdSIQ9nR4ypSUk3cfprsEmhQE43iaP4bInvhn0DgFUCMI
BiOtfzFZiGwXcnVi1yBglyBysP88Rti289SSNlozls/UjL2o/0RjT/gkYJQt1lPJ
McVPBowKhg4+d2aZJs4gFHm+CPSgTSNsxlGPGhHbkYDDCzoyezdLNoRci2JmXvjr
cKGwuDAAINU6q44SbEWi3Qocj0IZQMRbozDsApc87Obi/5b6opTql1qoPJCkhj9P
pe1CCAPS0ofclfn4hYwxEXNNjyTl4skuZ/HQfImhoeURxaK6Ni9Wft+xGedcyIFg
7j1QRiCPeAN/Iy9aI+mPMYRlhuVBQen2Px+vEou8e1DWd4KXTc09MWC9SXtOoq36
ggQxg1esOhfz5uIRr6mb57dy2MYqKp8oK5ZSZFV8tzK2cbeEu6DOQfogE8HAEPkf
nryMQoE8koZ9mSDNokktgdmtOHDrfkrtfmqlHL3TiNiV7hGI3gaYvYDp+XvW/A2v
Mzq5kq+Y+Er90T03AeFVVzHBiZizpb+5TH6PLhYBkd8W68O5j6RNO/mHg7saJOp8
3bJifXPIBeNH453/qoP/2+hhODEojJSCZrq1YGlknQMo0QKgMbjJv8rzge0Jp80H
FD/KIBb/nKHja+XLkElS4gdlQIjxjmOQxCczOzfoY84t78Ph7K/MU5wzcjsNqXKA
VZU89PLDgr0HbPyIu4DxHNWnXKfwGgCRLEVlnZq9OFZ50/AtMX058BGuC/zKhvV4
qAsNqpHm/1let+sTNzz++UHCi9YrHTiE880/t8FeK0ZgcbZiR043PPq5jOm4e+ll
xEjQQlBmV+p/FnZKS4pLAM/iau714HPBSKzSVS1leQptAVDcIe3dc8wivNQAwyWc
A2ABR4nf8kapAAVh/mSi6vCEMqbNfsSWH9WyZqq1zVYXI0ltZKubw4yeTbv9FEoI
bxyPAOH8lBfpATc6LAy/CBz5iidfpTBxgSV+QvK9PB1o4fb91kKgxpzQzcSn1lKg
tjGo+xTODCpmNSUWOM/b9pWz3a34P2AHiGIHFj1Uhbq9xLRvsOH9QRSGM53P55Ms
3ChIrLrkJswDMgtzGhFjyiY4jUbU2TTN5ND1fhtIj/92l8++VrNzXSSdIFTX0uBi
MwOn/B6sRZa+SVmfVEykEkxLq28x5UNYkY83rbv+laDvq/yT0Ou07+HHWAEfT8Cz
1UD1jj/sthrp6i1EPSD+5uf0cF+wupLoGfxGuwiGneYKkgDEpn0IfuIZURTAUT4j
RFrH/uvx2j0AjtsLVQ/2IPyjozzaTkaUV5veYxKZrzb5DuE9X6bVMjpcLroMILI2
jaj7xrjSs8dZEXPReB4Jkz7bDWSOgKrNSouqtCxlU/a0o5CGBj6PIaJexYcH2CC6
WQ4FLiiArc0QKaWAT9GG27JWVTjyg6bFaarTE64TiyCUe0MOjfkOYGC4IgBYR0za
9sfFusW1OdiGziRYk5a/oUcvogKFQQczEoeSn9iapPe/FjfV1wA7CwtSeUTvA7BM
J9lNnSSJIH2wKsWaXf+wixpovTHe7Uy9yuJrMz4kIkKQONkDF7F1+EXoaHZamqfZ
B/NiI0qf78k0x+5rTlrDxtLXhaCSOVtEJtjfpu+EiydP4HwSc6J0iWLQfzfyDglq
USvMG0UQ0LsRZmzaKanX2JAv0yVWHCjImkyUtjy2bi72b+NI47DUt8EksTcibw9l
TJZiEjh2t9UAMyroqD/ryBxByKROzITqVpR1Nb6JaUHpg/yR0bePaLdUErLU5Vny
sQFDGOxQC+eLYU0MI71UqC3lDA8OI9PYsJRquDuYxOztmU9tGv0cxTyplCP7HF3z
12fjtHhaT5OYJGMBxkcedFfmNaaOQ1gc8uJMmfxvZv57eyb0ldtLTbHwXFKbvDpO
G5BFNnlkUQ5hwGXG5D1y8m4klfXDYf9djtXFHUnyvnIFytoAXbJP93bT59gdykaD
DpSlM0mAhodPIHYoB3jmFjxkrP/wki+A6b5Q2JtYi6Na4RbM8M0c9INedmFyXOiz
6BGpZCG070LIq0lr5RHy9oYvPXo3IpzqUNQI8lFrdH2IwbydI3MQvr3IJHjRD6/D
MBVBi8DMkPddA/LCjQ0jfdZKrci0p2Wle3aTmDGf2vkkkNkcVrAO5YV/oFw3BrUF
tWAdfG58Ssit+z6wpXNxRL6cZNA8KaSkQzyiImkF5GvXDbmMmRy0ENPHNbhWa7dC
Wh51A+oWyk8gT5UCtN3t6y5khYZ+Tv/zN4Sk9K/GU6XEp+WaBSZLgfErtui15Zlt
S68hBgthGVaV4fa9TfDx+Ldd/Zxf0iVUBUh+0HlNhKje1jyxKQ10VJY62YXuDXam
pLVZsbTdjCOAfNWjebmKVhtivWrzTLuZdpMuISGFmVP8oRG4UkvcHPDyNkij45jY
qlcPgijwsv1Z7cvCqBUMbNaJhKaevQI4L2RG1B4zLQqk0gXZSHa2VUyOkeQA65dm
9ZIT8KX0UiKVJe44goLtIQRp6Cx59NOpDPhQ/LltX5Now2af667N1jdu0fpBgs+T
UhVp5dWG7iPSLPHdTCrj2etp1uVE9AfywLa9K0wf6pWV16U+lhSJTncNkkdaKTjD
nEx1VYPoOgLTQVK7KfDJTN0z6pzEzCgm8OYubAnpFAonXtd3lJp13FTeifTkNsB5
7Iei2g/1tKsPkTdMGEyHKR5nK12Te2TBaX+G/anERBOYZxkwhABXdTptGfamfHtP
4v9yuetDWL+uj+zlSrXEV1oI+in5eou5xMJ5xZx0laQCzn3GuH3WThI/MBd0mx6u
EUn2JD7cnf08lx8PzEsTwRlWMSCsTCn0JrnTd9i0LDj6AKwLlFbaL3WHYwST1Bky
F4h8Nw3y2gDET1qG4v+DdD6RPAWPBmGW3bQL98cDd90G1aotq3ai/HUT3Hx5V6cj
Wi9JZUalfUMGqhPF+GFUP0mUXRLMXhdHbp6/f5srLcVVYnRQxuB94L5CxApxm3PR
sE0Wi8kIaGc/z5X0V2G0gS0Wiiu1w6D3hBJpTAlqlBU/fxrER3MzC03vdxvZiiRz
9F++zTVTYX/TLbAVc1+Z9yGPAKNtDLZtt0BqT3wmahfvopt+sK4P3KvXsbrf9x3l
R++p+/Ntxd4Lb5Qv4jywbupFAMFbPfyd3WxmYG86AalXV5yU6uZ3zPKqkVieX65b
+grKcX7lasbT1CLAts1voEODVGBc4/VJ8DHSNxVwAftcpfjcBWHqqRnXibM5x7Fc
Tow/cDe6VMBUoHTeQF/6B4FYrt+CxC5TZGCanwh1ACSdL3gUnHo8BZTF45Is56j3
pItxOLbCGpAysk+MyzR5dCPDtOGPR/eGQkF6zlbUGjNPyqaCZKBLCuzOod7+ppY1
TIYL8TD6Kx5CFPWwClzbowpc5sW9EsS9fG9X+qDUX8QcWbquiSmRrxlQKojmbwZO
/clEtcxyDLTR87asVZZtirHTvDnMozvbRfe/B+jvSQwwYbbkrybXbg2eLplpg+Ms
C/PLOZoocmtfaJBWxUsHtOkq8cWCGWGTxoPW97Iqa9Vak9N2/LfDPpex76cMvW2x
5/rMo2l5Mkr80je9cSjuagFvGZuIsy7zLCx5ElpqJBgSgqVsWV9lmAwetuQMBNf+
xsB3cO6bbLQwlOrVUiJO7wLCb5Rm5C2ruZZbkhKIUUe5gSNC8rnVo/iBiuz3chpI
wHkWAba6PYcbHEXkgrNHma5ARqyXKKB4VRIgFpfVXbmliZiLXvwPkaVIr+xiV7H9
hJy9Qa7FGie2s4eOiRALYI5B4h2Jlg6j1nE+1fd2of/kRlZVJ3HiBw3rsM8pr9cs
dMgVN8yD0RKW3fI3FXHqhHInvLHp7Tyh1RmQSIVEhqpFLYCiZphdzq2+a2c5QEAr
UiF9PxL+V+XBv5A27jO5eafBIBWGvm/Qp5ECi8tNF5UvVmxzVHtDxr8x9g7JZjW5
I6LGu5a+P47FzKCaPhLi/e7PONay4I7ueJHOPzCNjXY1rXmbsdzvgVNKp+yUCTZG
eZ91ssPaOla9vsc/P08Uej9asaPgCQX8bA6AeCH4hlPaSN1gJaUPWlR1CNSLwpgj
nb7y1UhS7iodtern5KMJ9ALgQz8KcCy0oWibq1H5xrWRqBwZ2HRwnpMz2T3009iD
hAt63wFMWqCVl4nuCZJdvj/2KtmFr7s8AYTGbsBlsB+vLyAjDVeVaziCaV2r+EgE
DlbgZHhDEWHpn3cNZfjwU95DqS1ZcKUqX155g5PhS9OC2JfPfW5kgi8W+SpaC8gc
tdFdY1eMs10FY0S8E4Gw/98sbizQyil9LJcLfYdAdGMZzJSfuqyt9hCy6Hygjj5D
r7P3boDZfHWOroZ/oFdA0bw/Vx3JCTBZNVvOZ1hgG3kB+M4Bt+m7nitvbWKb5nN0
HPWUtNtqjP+lmWj3hMUtPqJdANWfT5y5/Ebu7ctMwB1WPA/3DCEssdz3zEKZ8M01
GPy9pcK7x7FySL/k2H1ShCxbiuv0p1E+mP40ji8EoND/uQsgzXRpxrwSRA3yL+QP
sHMAjc/6vn30Qyi/CREa2BBfCNFoMwVWt2ZA0cq6a9cxHdIRXTdCMPmeVob+CekL
TEXtrSYobbRy2mkMYtKx3LEMWy1qQBgKZkMugedVHHnp6t7MREFVPoMuCFGJBIMY
/7vY3W4T6k/mdEt6w60lxUA+xCm9neHrSiQyFi238vJGI4fynHNhxNJt3Ni4oDio
h6uoh5VKj3F9jIpcdBGU/8K6tQaJcBcVWwdUNn1rj3VcpusoGbNhGF4+8uf7IuRT
Lyq12U8n07qSxo947tjjHdTyeK9w7/0TVZxNj6xmNB4lKL3544s9zMDuX2COyH50
kpcyLOGs1wJwWKF4ghfGbvTKVJ/rtp1/k6//07nvfmp/R9/OK9nRqrYP+xwvdCBT
FNVUHw5l/pNadednT+Ga+8DQukQ754TQwCKTe60YPOhWccyduGCYajMjLLgDjKqA
r9lPngXuXW13Ijq2BlqANfPAkuHAhcWEGRZmH1tNOUtmtUIt7hu71y7+X012RETG
fY2qWSgXJcOoPxxuyhLmwI1MCWIpzYH4FtPH1uuZEjQ57O9HOTG0dgByEhdOHN0v
nKtKhf3G2kRR3z9lVqyJ26Jcn021gYis+wgxT79uI7Qz2Pxi2LxyAvMeNu3W+P0t
/6rZ+s0zxBzyF1glTYYTrTvIvQSSAUASjBgbAz/+fZEGCfLtW8g8XaI1tJ1SzfCj
JZYjItPEr7hAAgolkGQ6jFAuptvbY2RK1/6MD6ExXp0rdN3UhO6bPO5DjIN9mFj4
3oZCsm/SD23LbVuhb/29gU4/1XFmE3biCeT8McMfhTlth/D2yJvHYjPPGF5UZx18
wjI0DpvTB1pTRhvytKGGWSFBAvKokGavuembiusQ62hoSM6Np1MdC8CE933BXiRV
JdUi8rckVZQ/vU4LQFFMxzCETpTXNhUAdfDsB5CTdylxIcNGnFiavgi2hRxDWxLm
TsyEHHRuOsqr2pTxDYdu2heDoscT9jzkATnbtb8h3cjp+gb5KCsdre6HRcsXHMag
NfRybrQuH5fma5su+9bSQj/+7Gi8o0l+cqnGL8MjMMHpVcUYiVdSruKYZN/qEros
hATliR/raHqKCYI3STl0z3QtBluOw1alaNEShZzqF3U3Nsc/My0bibIvGQI4P+vS
5w3u8OqGnMW00ecaZ0wmyYBCgViuiDcTjRuu+n2hiawCOl5Sr88lyMHmXcZE1LVn
oB1UPSAAJnaMxnxVVQgC+i51dV2IalzjggEuRyxrPhIsdzq0wy+iF1Tw+fwXFc/4
llfG/agbij/o8lgtHlupu3bkdccYlmmt9JaTdI3QxU34LMzZhfY1vXzJdq92yjGB
HV7IS5XCAqpYceGbSacb7APG4c7YhQzoP1MIel+djUrzeourcbKeY4jNtREVAUxf
WV2EPlF8pprsEjyB7wHC+3cWnS5Good8s4QpWw2GTfKWwaVZn+aDh8TTloCXZtNX
nxg4GkZ/J4eO+ZX6bvJfu3+IV+XkIBlqMfVO1B9KbE9nXtGj0scTcsjFpFawnol9
G7lRlsZeduP6/OUlFQLxP+5KKckF7zbH2g9/effLMpql9SaghKp/Ou2mfplmAczz
xHyfigsY7GCdb7e6ue0hNF5r5bZP95/lVorlxAFdjsHayP6xRwAhPar1Pq1RT+pJ
e69GrPBYQJmkD87+vO2/fdwUglreLjkLm7tvdj2VCIYYEf2regSWvMhwiA1G3IdT
y84kzlNAz0w3qtmGb4nZ/160y32Epec2GIpWM/jpddBr42IvjRRktWzODqf20Utm
g2dvQXMUrP31MZjeHggSMt8QuZHPP2AIxf8bxUMKUiETnNJQaiivF7AvIlsA2tRe
u28uq24Y73NB8I3OT+/G14MMMjdnUK56OGWfrgw7olq55pKN6pnNsCVh57UE6suy
wkQtmeYeyNF0oZPCYyNd8GuYqZXvakmugQDZWThPLMNdSF3vsj6OEFumOOm9lVmx
uS4tV3hAvKH4SqChJVnFMU7GpwDfhFBeGngZ0CnafU0Ah0dNRsJpym0pb/bkkzKH
8borYWh/OgrTHB9tuZUumJDGqo10oF6ZC84HZcmL+80q7wDL/7tG33KZgoaH7f1T
hKzeCgRYYTK4Emt8V1C8bHsvGYiP0qGpRWf2QBnPnPtltXAc/zx/BWOIvkpsIOwi
WHrHpsRYUOulgh6s/ViS58P3h08BoBKLdEWkkI0DYufg3rR3CYdr/sBZQIWERe09
Q1NqFMaVFS6zP4xuujXv24IQxTZYKZmkf8jHUCCJ6FAX3WIGhJwGVdfa7jb4WmdT
BW3RIZjDED1tWTMfNA8EPqhkDK7xtnqbCzwaQ1K2QtvglDj/SkR0HGKPZI8JhLDl
fRESwYqTvv1qIZjOMSv+3iRGIrUxNwE6km7ngzYdZDdmvGSTdvdxtYOofvjSCCet
Zbg9x9oBMIohJmd3sJ3aGmfuU2nOU983AVEWIA8ivzjOrehSzy91J2yyZ0ws6Ttd
DzzMT2gHn1VDFh/BxdrQ40AJgeMei1Va740K5Jj7oF3B45G+chk+ENZnSkEUxywM
PmldcZ1zaeOLn/jD/IliFgZOlCbhas7imhE4MGPUJdIyEYoRH4OZRYX8KVWI+ITx
bypD+ODnJTgI3XUBh3Jqt31pBgzAiGTLTCdvAaby0fvIiHAWrY30dOFiedHKqIM8
fbj6JZZ8VSnPEbgDe6td30Z2Fo8CuaSelq8lj+cfAZlLZtdflf62oKzX4LAFJ11r
Rh2anOMWQKzDeLUr0bRFxloM42K260Hu5yHgqe8A9QfXWlakLiAmznzkN8vGEgLP
VD0qyB986KqWK0VZCbspEj4hseWnx0g0ka8HI3cJSJKI19JF+zuslkEotx0+IH0m
5k9A1UoSJ3d3RgI6gOhkZAzvFIA38jd1hVGvg/fJ880cj1snepEunzMQ9u17jf0C
EzoFSy9p2ArEmgMNOFcJSRWM68y6HmcP8F3hDmDGW3ver029mESeBhvzOTbp581t
qgsgZfbQRBfRiy3VtTyxnLJ7xIGZaIEGx1rxe9JCu8meAHsOFDs+cPBmWxVEaGby
A+NF70aN1QAoEBR52o7raOauvm8/g5hhtXIsx0vRpq+VbLd6WAHIXQtJ1JYoPkYw
EDH0/bXV+BtL2VrHvQ+nCNl8kNeOTme2TdlpNKMc5UbUQdlFn9ZFwjtAv6ARncVT
ItANTQI7RWLJS089eJlXT6+PNxwb1Vh9LzqWoKG00Q5/1SDCmkjKNNfKfxTmrbkw
U8cEeWCkRjs+qg1yMkp31eWhLEd75eBSX4XUwYXSWP+8jGbRnpTO3AR6NP6KNZ2a
+fB7v321Eq+HTIMnoERJIf/pduJlIXLj5GRbfXD3Ql8qmvdBAOCLOpKje2ZKlQot
+mh86GDrlO1/aW9uFfMz4NRiIIeaJtgSNo+gt12gysv37LE+ws2IaZs1dcN2qazy
f0gv7llu6i7b9bke1py3OX/Xus8M7DH0DvH5hy5lLd/3VJkBWEr7Al81z0PKZJ8/
Nrq1PffKatPPQbLa7maoOdeUuMMeuT1aH3TRLzYTLerBArWuWiQpiuZrrhHqMOid
wAm1fjd2tg08zxCM8k1jVVBm2qg21nMBGi3AKNuROmT09rf8i24yErevgeSzm9e1
FxVPF73pikXqpcEmb0rYwwxKSKMlPBu+gBZaCbqF6jqXWz2TuYK7pHPmMpDfVBNU
pWqczCHbkS1wP27TxnmWxGbpC0MtLMklMdvEtwfMuOlAUHdAXJ0KpZ4Fwt1JgEwa
s0ZAFt+V0tqtyyCxJN2CUu8UNUNLZQ2TbUSj3cC75KLkOkyF/u+gpLZYnbqHn52Q
bKeNKoozqPYpQslvXBl/XcBHoQ0ra8594lpIkXJHJgQ6pYGEK2NQOqtvjz/YkQVS
Ef1QVbiZYXsg3Cs5BYUjUu/tqi2jqiMG6CUMiTOUGaXtcimaYYfuAe89hUC6esbE
thWGoCEhPRBevDM3WPDPOuYSYt+F9n8LjWcfRxtuhLpcGyfsmOWXiyrBUQovYcQI
pGsp8HbNEEDInrmFAnGtT6acmTPTUSiIlzkjbdgKNEEHbOru6r0bIHIFtr8/+Y2F
OkXMC6wU3p5AsVi/JdNsdfcJEoDmp4V3LSPHp+QLL2E/l4S2Hi20uflGROi4jtbt
pigG/Z0b1HTA2aGlIpkdcB6T0m9yuwJB++AZC+a7h+bSMPvjmjD749jh3ua5ArCt
S6eznohXhJjBhkE6V4oFsS0dsKKhkb/wYEGfTrnD6crOVDZXBkPlW0HnBHOiQjw7
aHhNiclFo2OEREYOgZASohMyOUYEG4l+zC0MO8rc6td29jX01vkoOjSbjH/MzJEq
zMUFJblj/0zLrbj7J1+6bqycFlfQGfR3tD/dNB7Tt7MYi6JyS9kdYpsjKgYt38oh
gEiFbGqxmc25wb4w6U5LAL47atyiEStvSTVfniHfOXEx4VLkzlIQFByifbYLxeH5
VTHZFoWEyFODjuxFU411mBG7abqxaG7cjHpZ/uwMMyXt9t7yPNVQKVMaK7cSCalw
DjwFwiQq0EXVgmxYyH5Ox/6uNDXOoLtr6/DRy6H34AIoVLL6/xScs3BAnaj4+iFD
MA0tWhmvObJPwk8hm594Qd2OF/F1A8Q9fhg3uit5eB2rkBeZW2zd2/NI5O/PdMwU
SHjRBk+T1s8WlF8XtaV3QDfF14n+xx3dpum/FlmLlInSN1RcTnaXHET1lWGiviuh
O0DW12E4ljFISHA93FMib/YrZE62sMtRLrbXcAv0taXq8XNaOgeg6huL77A9J0iJ
SfpBENjdbc18QOWWkD3n7JtSfazLYuO6H1Cd1PAd1vcMgAUSm2WHo+U2EXmuNlHx
BIRwH9yoaadiM3lS1FgZ384yu7eoCesrQxI7nx/hJoHincZ6PRAGw+l3CWc6UpDQ
qvlH8QEUTSLre9tcJyzH6eW/HC87VVt24yW/mcw5tGbn0ock25w9zLNEhlbRJt+a
Vs0xrSLEPj0xI2U4DKOAUyeXPaTwjNHvOuSNq14SbyphDtCCXZg1gdUA9sahbbM6
RXviux1VrWZ1sw5N3yYNSBydaoo9Rztv066r0LaJIB9gjDsQRCSbz8ikBd5O9Ehr
JtEwB/4Vi6hkwBrHDt0kxSUX19o5Nua4cF6ecfUKGmBXvDkFCpKrtO9UV82kPqrs
iFTwetKcxQwDtBfg2dDLPxQK3dZwlyVv2OcXlXnh/2EEMDUaO54YrBt7DiSk+o6r
vma5xcbsdsexlN7eEKxN9tqzkec6Wiy1IIzDaD7jbuRSq4Vw26ukAfUMytyPWF0z
pAkEosory7rL2LCBho1SJdiNWUkRH9n4zPyI3N4ucTePARJlV1UJF3G0LAQkaj2S
vmgP2mcpYdZUUtBChLvpgBkA/PoRU5wR0f5jZIajsmVwGbvi6kRu9I59rVZ+rokb
0S1Eygs/JHjZ2vAgTQjiF8ohiRZ7NFeNV2DUFACgDJ/PhisYRhGoKUBjRLxrRYwd
N6ShIARO/JpYSL27dGyiazlkPK5/5f03p6pGN8kgWmO29p1oyrqaUfAWicWzAun0
RuattfT8tJwWLbBnGwJMCOPkVZ0+3/q6s7hZRPeFOmmYPYiRG10nKEs26KkoTgqA
PGUq0ue74qh4H4/prFTIi/IClI1+xVV26hzL5OOiEFjT0D/hz0JQbhRNfdpFy1ak
rXp6h2wgYOnmAeFaHgFKdG/jWOjQC+BGBtb6yiDomu2LZMnV8odB3xf88m9S3Z5I
vquYMBrwCErrxJUsHzXc9hxucaZ8F73KlcS8CC3krpsbcVCoMx31TYmgGN1LDK1S
haTvcNLcGeXVaNptmEEYyyFdIGP2UmlOpmCTKdhZZ9PBa0ZTwIkiVwWIbxQk/mzo
11NiLx4sAiOAyghoQdb5U4rwkFzcLLuNvUbEabgt8jFR634c1o5wbd1zh70f/y6W
mSGis0SLP5CsGPmnpyI76khC/u08/xJfGXTTD58ueHzZRGwOtHKAiaWvnVvGuIiD
6MllbUfaFr0c9VwhLOXrbHJOfhd3xjA9ibQ63hD+Rw+LMgFW/9kDZRXEOmcPIrAH
K7WvhzpiwNQMwwjOlNh125mk2yrDnBQhzeTO+M+dC2qTkQzF6/KnvstGd2o5RJ/H
Y4WI/kBiPLqIyyftyrhBQscvZmiCWwpv0ooJIFA8oO17t59YHVdf4+FsQNlS16oQ
+mDu2nKDRXxvuVHXbV8cgkuT5q0l90t6J3yeG2V8aE0BrBiB6d069aUTKvqn6vjV
PifB+ka2L5B/2FKT1hkmZQ6vGnBLmtXJOIe1zxLayd4iTtLgeCsbj7XwYmqHzFv+
mST7FZWcxgMA7+hx3P2RQ59rXxqNv2+geIHEC2ibPUayDPcBf/5U2wH25OJnw1s4
MviNQQitmXzZdLr2QwGC5d1RCx2xvRG5fessGQhs+pDIkzjJLIY+1HT8GkDOQm5A
56QDWa9Tao+f7wEpMXePdxeehelK77TusnTqEIqGsxjLPusKHGBmNlF3lgF9amqX
rTpZzubT7Rk/hsYdAQJ4ljUk4gw8iIvOLsUhV7U2iIllJ3yLDfnuXwZ9cA5wRlnh
LJFwQLTYcYWuHeQFVdDCI46JUWkBM5aowEoWdUy1d9tdPnHDPRibKrSiy9vF9Sps
4RpMvi4wsIKgJLK+5De69tnKVgbwLYIJmcDAT7JXDuyWb82ViOyXLj9I5IN1iiBc
fRTMd7/9noFvv1P8Rf/ewYiIvQgxeQs0j8fSo32oM2ghdnj6mj0fhaF5mQUrspKL
aciiDNzhec4NKtmssz/rG89temXRRu+s928WxO5ubTzNibwTPGapuZ77wizleO6K
aF8Y4NMsefwcmQhFe2S+H5whDvhkeO+tNd8QPciLbezTKDQw8/wfUFfQJHEScTjL
p2DdN7NNm6NU/NHhLk+QG/eV/OPKphifyqCNP4HolXqTm/IXivEFa8dNDlROdNr4
A94lWnYjJ/OKnASNouz4atsdtovDshInh7+gqEZzyhvqyEdosZCWA/GaYhb8JkRz
TldhYtxXU08Im9IcKylIQpQ3BzoV1ssqsChr7+p1/oiPImGD1O742PxPRqgGjxpJ
wvxy0jwdFYsjG5LYrmghqDmgzqBPDUfSPJlq1XXAiBkrQtl/ArE/tqAmU7ySnZn5
SCjoQxgL1Le3oykfstLhq7AFuBCqS909HQhfJfVj4OvR37PqsD10RF8JT2n3glco
6IqX5cn6lHiGxjJI6ytQjq5aBRdh+3W9vvxnida6Z5iJjwfMuJL0uqvkVrfMuvLt
2rl7Oc9DgGhVNAFsGieCRfFVfSp4q9vMaKKkJphvFZUgP42ttTSizfH+Qu6mT6Fu
gMI0AimDzqzSWgfuJGruQIo0yrGgv/c1BG1igEkn1yJnVAnkjY108N42jxwfV9RY
qgfZi3rkSdfdw/+JCoyY0TiDru7Bzcl99u4nfF9ZNMbyjm0sJJYKq2vya3md18yK
yecMjeEhFWBHV7KTOmucaKyH1KekSOdd6tyAgdPrpdhFwrOrujcGhE2NiPJ92q+i
yFMCJhc0wdfY0Z/I9SmwlCbCdajJBlem1MRWky6QcjNPmsCiSYuseSkGIPyrEx8t
JNG5iSQTKyK4RKrLdrsoK+qAHFKnYvihwJWH5gCpsvqmIcFeuBuhnXQsJJL7bsEx
zSlriBOvYjh3esr+mlb5TP/s+QoqbyuIP8lVGJon6UIiGSPiZK0d0dg/oeytdn2K
5dLP3kF1LP/Sjdfv4SY32iduRyPjOBo48SD2FcbQbNmF37WMywbbuGPI1veB2iox
7GXy8beu9OJmulXlZxFO4ucWQq+qDJxgY7eqeHDvUyzAwcqdAEcAsZ1gaS9KH4Sf
qF52ZEAhqb0pUPS6RIL0/QWk3NQMyAsivhh8o9gnjeSPI6D3VaMOF9UU+IL6xOyZ
lIvVxvakRZRxqU4QD+anadncf7Jh2QtsXV5XsN39LdfTOiPJ1FdEm78e8lceqxLD
Bh01lwpdEmMncrH5gebVObooAJxl66J6KGDYj5CFoTy2DKIIkinsocByfuZqbBI3
mcFJnGay8hZqlU2sL33QTP53Qoq1LykheqLzUJuCBCWff71v7O4Lnp4pBU9d79n6
7WnXkJcjsQ7DlrUCpRRLdVvSFBv5uwz6ny2g9lLV24YvrXEnWo1Cy2P8a8L4smTs
t8nONe/scYAGNh/Kbf2zTaPiob+IdJrVboI6epAxgQfMwsgi8v+ibXg7hLOpuf36
FiOVCFTpKWGwyvnMnfFL9YwaOkFKdWJmITIuLP3zTPOoJvg1cEnGaFvfsWqI+BxN
Tv/M7wn3H8oHQmFN+ImmLUoYoVLVe9OdC8HqKmTdxTbICBA7IS4opKSKew9bXhiV
cHK2Q9XtC2mZoej5V44DNIZhzPSagI/LIttB+F0Je/TfEkHBu04ATje8D7wXMXll
7Z0P1iicoTUOdeBWKuDlvwxaFRXx1ZmQaxUJW5z8hBHzWuNoqGFcFhkrctC9LMDR
za+jEaEog3MFF6D0Q1T+RrCIknl/rS7XxOCBrGNmE8gVN+6Y5YR6LuuvAGpioqXM
9mPpl4cnDBg1jON2+ySHy7THKTdIVk+AOtQ4SFzgOJiWcP67qPDmsxf+VFIKq9WU
XkaTPSI8xg1ZrEvObfRjJX8K1kRyIR2b/AVQPnV1fOHh+fM3BLtpVOi6fWHBun6a
pCr068w58v3PienTBi1CMog9RR+Vh3frvf81zrnGmR0Dy5W2rKF9DzYkmDuPcbpp
dxBLx6pgMbhuRfHaC77o45VQ2IQMR+ba/N64ezUKHXr9rsOJaowroUtVfY1qgXIv
WlrFZlayQjNDwTem/9S7q7DYimjkEQu20xGpdjloUzv3Zsi4Aa7SR1zPClEjBbXb
WAEnFbcfy+U+bOoGKu00G/4BWhWKwFIcQ/+8QfvtoUXRQ9d9ocl78M7LstQ9s140
kWfdBq3SKqjvBCyg9lFhunYSUCZJQnqOAmhuIgg6n40UXMzGpv4XPIjPh+MxbXHm
UXs/vcvKvIvl1C0gyZNUUaHP+mOphuAJi+mTjCWXRNxN1AlnnGz6F+/tnJ5jO3f9
GtlJUiIQdRbPHJVHHqy1b3MsuvKWZxs2yRG2NsZuxLXT9q+R0edTK2yovKD02OEO
A1QGmdbnyHFX4mt4FZQcskj+tgdMIe3EpRYhQKJzf+sA8T5GNH0PHNj8qP8mWLIn
PGST+953JZAIixtk0111sEvQAZEPb2V0r2GQSXhLV84embKqtMf2KaAyI3VOqo5R
XIVraPe5Dz6GCIkFw5xDEbL9774dx4wVmGanVB1bL8MrabDNRTJchoZRHRXhSVBQ
cMYwHiH2RaReGu8gSLCqelrkRioKS8jG4zLuszPMA6AhnnReN1RSTYJXEsWqEnYI
BLxvgHXWKDwQ53Oq+OwKAKe0icmF9OragYPX6I9il71j5UZWvXXgyt3y3MDG89tW
1aSeWz/IpBh6opi5kUkxFlt7PtYEL2ToPbaqZNDcxD/tWJk6X8j9SjQ6odyXGpIs
pMGqL7GaE1hV7RzK8u2DR51O/BrATF2W0RqDKu+k8uFi0tMSD0KitUrmUl6tDdym
29hBUNzI5kShyyMe8FS+rs2uFb/WoJyf2pwuFnmOgv0bYFw6bnFoeCbjfcdFEu/+
xovi8thBoU+96a/TbskT4Y2s4KDc4BszVm8ezBCarI8JV7ihUick3nv8OoR3SSmu
U9FgTJw5HHnMwMnQzx0ezGV4003hZh6cnOCmwOf1rJRkJpom1kqo71yUxD57hlHA
vF8SVyD0fwaTodPCWh3hCHkBaRv2bfG9zCsJZgk5wgzDifCmwlqJ0bZS9G8MkdHF
tmbb0y7EKJMiRVdwxmY9cYOCI2qu115P3MIPCxoaumCT6/aVcc1AaUciwxiH8teG
J//SlF1/MiA1ulgTwuIpQQsXg1pGb1U8myoqY5r28E5HTTDtZFYPE5/7Fc6MX+hR
KEcsAvGpsOjfRYZxIQMoif9hEcZqcSqXyy1Ls/wxartAXODNXo902IXqgQY+CxGG
2OmeuRjhS/77mjucUT7EAjqTHBTM+TmkdOcF+XxQKJ83i60ho5DI0XWxS/0bkZCW
k6EL1SbnQiM7XeloPkPNBhbArGJ0zhirl39w6TtqmC01tho0h9iBVLcIJsAu5+tx
P8inAUpBH/iDSF5iH/RLg/E2rZKr2V4k8Bnzs0+0iU/qz4ViA+vDe6wmHHPSqDyX
HR6FtKsuuRfRjk2cuaV0P077FDKDMY49p1ChqcacPFDoxxp3A5etB8A5Y8g2oaI/
9RnBOrj0uFTIJhhSchOblj4ljPJf2fPX45onsAGDA6mcLSpJUyZFzASrkLxkKZOm
b2WTsB+IbEfD4i9IDItUPmyejQ3OW+kncO5GbPqKJ4ZQjU4gY3A1ARe3QyL6f4Y4
KaIu1NSpWVbHlpuFLxv2OJOBtfdL+tg21QSxtqwz5hyrr1Yht6y3/r47mQTPF4tC
4sDq1S49WZVEryglmdTAS4lZjmGqAuqTlCkV5G7r+PJRLDb/3+FjHmB3cjYO9mb0
qccWKt5t6qwXkfw3Lfyb3T/89l+iP3Nr2YkXJYpar+cLVa/2+x6LkUDS97OQ9oB2
uW4aE75mUHpOK/wqT+lbi8OljtBiSwjDiSc4exxZQ2LmFg7RsTCq1X0TU3usKxSE
JYdcHhXbv/Tr3XG/bpUbzMpt4dZBHGB8ArRqzDgeNJSMFDCryOGw06PPo42xHb5p
1P3NfS5zJLFw/gEBww/7lJmkJk70fVj8oOk7lzFaOQepnlOvzsOr6gnZB1erGtOJ
JEPPrqRR+9WKOcQGjklyNRZawCatFK2APDkwopdYnuw14bfgwDZPNj7coFeqgANO
yKrEnobyFMkwH+teuzeFtyFFGv4+Vn1M50YCKJp16dHaRU2ThsGi7bKn5lJPH8Bc
9RGzJH/fiHKqNwuR30JPyH3ytl9s1qtoN9I0zeVyHbBS280Bbyut5Bji0dbKM2dU
OAmWmwq3w5urjitZL7WtvxKrJgoETePleyu6J0eL4BRjEp8Bew+Jq/FqN9kqBq5O
zfi4rARBdVRwCev8q8QMhC2OCdO5QqCDxhe7/LFcQNHlFX25/Txs5V5V0bTaNavv
2RDQitsMNS3fFrp839So7oO4aDbUlKX8j1yPL6m3LIPe/82VaGgASlfuUo2NyD+2
bi3KAI2wFzm1Do5pkAh0x86UV2PpxvQEvohlc+XHZA3dbbqLgwcf4kZWesJeLVQE
334A7U2GRwOJAOAdmTU0gKXop9F/PgD9DChMZ0+6aDjtkFuoUwFyH3AE/jklTOiH
IdFDwhjDgOMsYFCklCw1gyUiXScJd0U3KSafpiN3xBk/kXVL9UMEgIhBPrdEekEe
NBnP5r8smZHjpYcCyrkNb7FReSLcdMpcyXSquuvP2wuDdOl64ihs+F3/oTr71XX0
whdAbPxJTgiPQb35rEn1/EP5uHK0GmYLRGDTFyu6WLdO6vAHodUmd30zq3srC6zr
9M4gG5z2lqqDNDT/rucmEkDEymm6hyZK5mnLRToQAbRiBKybnqEaB7NSqIbekO1I
nS7itKcyQsMpLrtVcyQ96Bdo0bs35et7D5thILQhOcrbQ0Q7xEb5XfOyntpxG25M
6rGnV/NCgYtr8ZVq63o28usFuczjK/3X1M/XQtM6yybrdF4y5YSKr/bDPRjlYCjZ
XhX1M2cjiE9FiMicliJF99dB0vagw11WObLxU90cyeaF5F8HIlOMgHTdVJNlJq/w
Auh/+9jvQuorQHu84kCXvLthQYzA+cVQg+HhYsA/UXgCqtbFyaJ+UDnkBLyHy9D1
H3pFbUF0QEDVbfyb9M3SFVQOnHlgpCLeZnRTbUYNJ0yntt+47+3E6q+DogxcICoP
Mf+kA0KfE2Pz87E9yrIbq8+VfQNztzcniK1eX11S4s7qQV6OUCdw7qbDUim1+XwJ
NfxGwZubB6wJUfsOajSoGNa5VlSrg0Z5upMoGXgC/upuJ6J/9+Jn7B8PeF78XqT5
XsrLPwe6lZtZLM2l6thDrGFtpC65zmy7Sh0LEVSZKCL221MYzIahx57J4fJAPkRQ
hCTQdgb7Bo0oATmywIy29pdF5cYgPHKNZy8ns7N9Fz7hVOSvPmd/6DXCDb+Mf5ND
nE6jNOtOlqY1AWnd7/zjjkxY017i7UfpaFl7xoJwbVSQxh5BjBSPyQAfRyjhxlNZ
PQDnQBvP1P2gvOkYvLZLh2MKiO2CJ/bz+APgNLe1vYyNVVrUv48dDFgTFneKTtwX
yXKe92U1o6l1gS7rf2Z4cl8KVh+dvGjw7L8xSaKj2EVO+8x16h2YZkbciJ0vUOJf
mPZ7nysWP71gF6eq8W13caSqwrJQ3rzq9ALxBkGOT89YM2QDeeCUe9MLmuJjN0ow
vJeHK227oS3ZOB5WO7Zk+F+DEQIBPhsLhHe7x+oVO7s+6luBx0/zrraptP2FB+3/
V79Lytl5sCEBcyTUtSyi0KCsPM1Yva/9nohDgvLvJjxx+65+qmM+5oSQWOZFdmFB
NTgTwG4j4kX9QTwYYtYcEcEaez5Ovp+1qmsEIbjG/Hw6OxswaX+WBvE/D+inSMWM
uHMiKO+UXgqdEPT6cTYS7z522CQWNEgvny2zvptnQEjCwVI82aGtVYz/CEa39Gpm
GOGEbY0GnWVSaEAOIhCamBPiTbR1MXPKm+jZW/80nMJcNGb5UKyv0p8hy4duaiZX
8D6JED68B18iAMBRd97h1jFmn0Lqq/7TXYIHZN2ZXpagmXEc9/sKAOW9nIYW1H1a
7VwdiPewxi/MYU0dZ/lC/brO/rg0z6dL2cVaawu98y3bPvG6x+zqqEyfbf5jUF+U
KEeWxAFBs9nG71lLuyHOqT8cIisxKcMJeAdf2KnBLNXMJAEJRrIKVHVhS6oqtiDa
fs44Z8/md3dLcCNt5T+gAnZobq/eTusL2LtTpJq3Dz+Wa2SgFpSxuE+Mt/D/WAsR
DTHhDJIb0QuH+IfpjOWc8yEp++PY8fqKQ9cl+5HSScwrEHy8S8Wbhd2L9IBzwh/E
7fYro+zLfjOrnwaLLB3QDxpNOMB0akr7C0U7UWP+0MtOgq5MlaXLfZXuTb7TKwgA
Mv4W+nr/q5pqV5Qy3MhIdh1DAjqcEXVjvvyfWTMGvKl9Ujj03TDX9LghO/TDS9T+
GYO9TAMa0/pqiLEjFurazPGNyUPQPBOphHsWyYIgO/0r6rN6WhS4cesa2GuUj797
OaGZCB3sln5AwuzxJXdHINeBJe249DMFahfgJNFLEcjzSI8sNTIV14rX4PSBMi5r
yoAL6txyvE0o7tCj0GBWL1UTsamEvIK090tN5+pzxPOr3SJqyHkxPficQc8ypdlF
Jk5zGhPYD4h9ltCk5aB67tLByuZI6wvB1tMbk8BSHSoLzCB0YlewcG28AK56cJY/
fjfhdaxjdWsnzfBKOfllAzdyEPfe/QXI+udF1KU5sA99XMLb7Z33bLZbj6SQix2p
HcHJ2QKDWOQrUMjNcUt5GoLrjHNzaCG7IVOGItYPzpAGajEa6b6uXVk1ftdyn5bz
Wxyuz7bnrrXjEQkpeOnje0MiR5uqo5Ax0JytWWZ1M6K+Te/dTGR4PZ4/sEHslzBK
UePV11FqD8qrKWQuc86PB9QRJPs2eQTQUNKA6gmj852xaRFLI7v6w7UxjSQC5mB8
DtdS8DNISXKXt5Ik400w+u1ywdrLl9BPQU3LbLjwjpR2nd+3GIXSqssi7MZmoATb
eD4JQ0TJ7y5sbUYb2rZG0erNEy8y4ylom7wDesG3dO5lYem/Wgw+qAXiyrxJDEMF
CX2GOvK9yI5t/+UMZJfNjA3sfJyu5xNnSHtLOmoRrjlMRywspOdeOnwdzFMLCYIN
n8G6wDv5++of8FyjNuIC8XFrZkXlWz2W50aKES4qXR5jbiPcCow5qNHYESJaW6vD
+0YUrFi1gD+sCOeWmbKJ1KzSfJ4JjaOR+awEWpCNdQcUMjpKSdbpEPRRxAw72t6a
79EmD1vpWelaWNbqq5QRHb7nBtlJcpeyl6RLRW/1w6ANQmqa0bDLOJaSipxTTaU2
sQ9olDVvQGqo+/kfB5jw2hGw6YwbBd2s5IjAv0d3Pm5CHECwuZZ410rOg5q+w7Xo
lt04G95I1m/6XpEBeizlYxXZRPbdAKVANB+TfjVy9mgJ2CM7cu28JotrQzmcR0Z9
LmkQ0GUq5QZ8LQfS6n+id/wXObhVZCivqaaTFgbcZbPXrOOWGcFMP6aUpWzjvVY8
w+3JCJMabUBW3RllgTvnpjJPUQBO5AuMC7gamCMoSUtFzcjGpUk5qdnCFWaG6HY/
+Us/3Po5EihUJOUvvmValg0aDW2bJuup25QNYRLTR9x4LqhJVr9ugxex5/ejNMgI
s7Dkzq2j2Z4n+sStTjseVw0vJA3JAPstMmnBRkp94sc3K9Ew7Rly8o3PSGbCvbNh
L4Y/P8rmAWQ6zE2lrnggY2AaQf1k82sUoy6FEPr7aCvTAYBW+ehaAaIvi6cXaoP1
wCAjQEIr2VZT6fn9TnnOnnqNNySoua3Dx6Z5dTXZhJ81OvjpXf+IsB09KcnZYuHp
tOwanXgB7FOHEQo3i68zv/CtMhz9zoBkAlpp2WiwSK8SB/PFQ2BO89Zo0czlTE1u
cTxrQlV7opB5s6XrPNgLtZbUl7iAkQ1tMRoCNib5l0fzEKbxBcEtRpJOt2YZTuCk
CF4S6Q3EoV7ZkideLi6nlxEOWxexcir5INtV/oHK128/IZf3REYzrYpYBh3/E4xO
uPrGmB0aLXlcxvrN0u3jzWGWLS8e1K3q9S1p8KjMe+Y8ExRH+lkY8+SEOmtYnrQL
lq2k8bfsNEvTfSmstBTJcx/9dzJbQahogSmFj08bWMxUMO/C7qmQgmzNpZtiBTH9
KxZydpq4mwD/EPSqykwm7+vYz9U2rAj3yP3h8SDPGT0+vyQEZ2BywlQCwnqEBga+
YE3PLuymfN9NSpJGV/BK1iWpgkpkTrheix+jLfcItkqvHdqhEFJncBbWa4EBEH4+
TbIWjZzhrd9rQ3EVQ8vSjHeDGiJXEKiAnMV83zijBFoA0z2PS+LMZB94FwKLf6qQ
eP0T+4OorlSaacU9129rPkz2v9K5YY7LjTWwZEoWKx0rL9sYPgXpDU3ocLaJKn/z
C7FzauyVWeiJ3JwmZRt6MlndjRrYjOcvP71lMsAdXyHC2o0f1T70Z7Icw/tpa5R6
2zKXA3Qq8h9l/NlfEv1zEW5KFBg4ZwN7plsPtsd+OF5cF6Vt56QAnHHKLxtM4vCb
xJ3mIyRP4qCortrQwIAccciBsw0XDiw/8aCZKVFYFhnNRCcYqGafW7/1FjS3KG8I
QIpeZTiUt0LL1hg+s4HouNsfrVvsOf9TrSMm69f41gESJw63aVWua5Wa+smecZGQ
FDlmhOXWSMkdO1isW/hvKjtlUal6VKskGBvZ3DugFuxJSNlXOF1S++LrJQJwaO1h
Pls4+nEfceiPLc7e6qwMespUFhZZ/2gw/ZmamFvWsMu6WQHN1dv7DG8XPPl87Abg
ux25lM5/w57s39zrocn7T6mzX28QLoeA6Gi4OU69V1+YSO8xnKiI5W8TkR+eDe9f
zqjw1WnBDR7hQtB76ZY07nvagBkxSLL1cCLkoR0w3cVmhEmogXC0hOV6ow5BJGTz
cPiTNU9r4aHStvF0R2AWFvPTtNsKO1Ms3u3u6d8pNOXs7+kqMw6V8ZQRSKSRSCzv
6/UtKu6HdojDwbMEiWE+yR0VRADN4Ix3fqU4qAhoyV9pGPfyXzvxWXHNzPsW/nxP
cuQkASXysxv6YRIeNBMLdiames8stfrxrb6GUBHma5YiSean7RJZ60q3SIgbmsGp
CMT78Qv9gvO4I9ep7/cyKMFyTiV+ntDc21J7IXxXkhcAuB6o8YVmjAmFO9/UVsJJ
DhdTFULtrzqmc1WlKI2dDQVE9ly+XlYC3cqrO2pDg04OjrJLdlSB2d2xVbD4jLyF
G5FLNclb7jb7WuqMrI/adHHqD4+DYXg0M6K9wwebEFbmR7+oFB5V+QUr6+VMXt9a
4EgG9esoJ3SX77A5AQEDRVR19pCaU2gluKsK1NCgfgcy4OgeOAzVHrA0JoNpRexb
bpcY8Ibwirekjoj8zUUzGSTPu2ugFJ/G8j0J0HBi0lBJgYH1aDKffO6MIQIJcE3V
DYH62C4jqX46LldEhWOJKx+lwc3vNzVQ9ZZow+osVucdSK3SnGUKzxG8tgkl2XXv
4i0cdHEpLdi9XyOEwf+oETkyB+127ptXzsp9k1vUjJi32FL0zCTQW10VW97FAQs7
gIXjmPthccLtfelOksQ8kEAagC2Eus1QG/ZZyba2s5bxlp9wXEqNO3h5JJkc/CR0
TEafxUcm2eiLy7uU0UmPK2tgc0xDA23XAj3z9Yv+qTy8GJlurNhy1UR1g+6oB2K2
+URf0Zd9YkTt7b5VIbYIO7pmDFD6eIeC6KpGDUaBtfXK+frN1okZuITno3wHSFuQ
g2qb6fQW/DC8lBB00WRj2uWbVXK63bv+dFfghIexprUhCfzzfUIDFF2rcuqBbxWj
2JgA9rs8t6Jr3b/gRk4xIiOg2Td/wA97Uke4qFbg4YjgZr0rjSrxOGupUPLl5vRE
c7Z9fw9Yb7H12hC9ic6RJmCLaSTO9q2QG3CQ6WplibRmewmV52FsbAgB4EMYWf+U
PWde0MN9xjP3LGJ9vYcEhYl5tRUgyKzlia6riCyYrsF3x0AmyZNxG/fHZ3G5H32L
RooL1FQD5ypjqZulgyoJ9mGpyA4NDvZKZ7FYxfieGZ3Lo9E0Ir2WCakVSsJ1iZ9j
0IPu5NHDIQTJtFzmf75IhpvQL+KnZMqj4OJ+tjrLAIWeChNghc3kFIrPmuq1+p6C
QMGOr5bPPF0HWqBKqraUQODRecrV/ZvLF6k0bABT/4pCcGJ9HClgpOSysyV+RrJt
tUOTPVmSNYwgGVRin9B/OHO97dV37gj2baRvUhlzligXfE471CTvGwUsVy+BHyey
5IEpYT3uW0Shl8K1Yk0r9boDb5Ew40GaPGhNnHyvAJh8wHZCo8mnlqg16FhuhprO
Fg3EL2bwE+yPQiyDjLwGiqnxu+Wr+zOZ09gS+VsEkJSwT4GHlyHeCAdbicbteYOp
d7qAx5x+iR4F9RTHkx9p6ggkBQS0Lz3bbPsESiMSLPoXm74f9Sll7O26biae2Mix
iafF5N8HcK4hLJdGHFUDypDTvLnDVkPnVsqq14uMOhARKybTJJCcsH1xHppN6riR
2zaaQ1izIcO+NsGWKmpsRWxCM3JlyzaCExSgkGYqzY2B6T+AbzMJuDElj6RI/h+3
uu7+c/dPoJpqqw+PJzUxuGBY0njk9Q1gRkjBiLTylP10rXfq0pStJ1NFtE8G+egd
wxkK4/SR3/4slkmup275yvDmlMhqK67rNiK5VxyE04wUjdgsRu6D5MBuORWya2tF
MAYRq9Y6cfxXojmwJlCAt5j4VHTwI94M6LTpvi/ae413KGmFmX3rKL01bL1fwp4M
uzcoz9h+ju1S7iWDIMTlICcYzkOo3h/W8qYUc2toF0+uWIRrkxW0dmfF/ESxV9Cz
R80eUhVDwcbRxlbgoIuLRYV8pfvGf5cPHb05OCERUMymD9NM+QwnBKvK4YJb3CdL
m5MsGmPV7QS3q27LgysZkCKELg5cyHUHX5NQJfkGEYVxm5LoPJsXT/dIi23eNUel
eClsZzo+ZQMgvEsFHL8XOPiSDDdL+1BPbzxT3ZFBQb4HHwJvtF0Apy3PliOYoDCu
iOhW80sCXe8I5W3Sse1DmexljG9L7PGn5EWBJ+0Y4B1TN1ba8U+Y7UYsfcpcS0Lf
KfO2cqsZqA6P4L/ooW+hDyo0gBdyP/r4f3utGrav476CFgFQnZ5+5C/Q3BpzYX23
jHn0ZfZn2+ZU+mTMKGHnlIyso6k/8nHKu8DIk50m6whUqyANXGdVTc1QczIj/daT
ceCviR0CmsN3x4xbtH1+tDavid2L+Kc9k/WjqHao7PpA/wAU1V9RXqTaIreVPNnY
UFjWPoLI5ivrEd4K3k+eF25OwIzRsojKf/HuiwxtdV6svmOOWDdMZY66yPoBawlw
WYVaLLCuQzeHoXLbldjmknypXOOM7aYcLeWQjf1joCw1zlnsiuo6eXgBSez/aHtV
cMy0rPXgGzcsWgdUHqIKnMOXIegrjJwOFeNkbedzK7ItzI3lDdFQm2n2Dc14BYwp
DHvoiD03FSxBCGEznXjuXTOQy73g43PKc8GM36Q1iSl7AC49JLKa2AqO1rFk/s/u
CGc9PSLyFepgHVh5llJWY3Iu79u03IGr3pssDThNQmFBlJUy6ZaXK2ZOIrrvUuEs
Dc6dyyzfVxBVRF4B/apC+dHoeDZ2oPGsaGpR3zrX3Ui0BMvJ80vxRyHzodAdod9a
1ic29iwOHoSJvAQb9db1PIK9CZGRLfOSy6rgnnaL/5HvFQOySohMSV5/ChL+uiZg
NwSRoJKhDndTxVoNH98TsUuKvSVeoILep1L2tvO7xStWydenyzJoNk6lfzTgIgtT
VT/pC9hVaAWbAee4WyhIGADSfQ+Lf6MCbI1uR9Oc1U7pZJKt5Q5SpRgZNNGGbmnH
XcIG5QrrmJZ8hj1oEAzFkA3Pk4T3cjgvAVSgeAtaqjeeJc7o+iAJuhAqGE2u54jO
l+ErgKAY2ymRc1KuiTm5uIsfxJhAWwToa3pErIqpyyZMGkO63VICUBO9Bo6dzkCp
PYRK4Df3aREnzGeqEmG7XAZasufyy5wJjsyT1DP8sZqz5EHocfg3Cth336Iat1Xd
DHN0fuA9I+UkpfUE7q269sC9muZt/8Js31+SAftCadRx3YaCiS0slmzWLyGTAUTM
bQiwocalwUuMC+CMhTXELlz1odKBq+yGvQedjP9iuoIpCG0ujNLrEsoZfFsInmRa
sVv1/aUW6lgozijdKR6LbDLKfrqln+Jkc6iZv9SSYtAyRS02YexErW1+fxLxhy3w
bGp2vzlzpD3piAgAV9WZrQMN+yZ05GT6/8vEEHCfGLwszbXTS2XvCCJQEaeh9xhG
Ic0sHosihiy1PynSTDGKG10EGQpbJ4bdZwb3AREpxBqeQEEX4XeF61ekSgWPcIdH
pGE6HZQtU3Lm+kmNx5bd7bikVCLkkTKwTj1oAIPiEHxk6epwvKIjflf3DDkTZPQX
Cyn7B+w74b3IETvxJcmiDP/NDrF/J0W51N/5YxTtI2FWnCzsslPgZ2HQNLdV3MyX
AFgNUK6KCwcEK+0MCcwzabnFkmyv3WBGnxqqLx7hGRvhtDmC3luAbQ/HBVSynY8N
oKYzqHX8V8c5GAsMdosa+cwg39YjOcZIo1AJKQwj/Tafp3uudl4WKBFsF3EsYek5
XUhQ/Vvq02nLi9TUIrds3tb4GAINEOAfF3TtHHnJcFBT7xqEUdy3UqiSrbZe5Jex
EgVVkAupcCvd7JR/BrCSJ8SW2AcpRWnpT4c3syLp6jgRlRyyA7yeCgK3EG1Dts9u
JwfVSF17J/p3zw5MlykWnqsJjJLCO2lHxTzyrg23Wpu/lHBnSKb+bryh21S/7JqY
Ud9OHi/OQKlCFsnD0KpisJcIjlD2A40cwSR0IpQJ7FljyVcyZOaPdRAH2OOfRkNe
pKHW7jXSb3MYjwoe7wLYCYF4N8ryUPIxP0GqKfPhlt6fmM4hUs0qfSmCRbxUwjuU
RlIk4quxn87PVncTV3DEbvV3jrlpcbhIn7UqtbHvdVsc1v3tVdpHdyEkxIFW0zRE
1FdHaCNCxYYwtiHYjaheDcwFh7s46R1v0qJqGSZK1T8FOhO4mxmandDaEPV4bea0
uMmzngVpdAZR+kqAk7DyI726W0DKJrJyw6L+goFed9+1XzH47hdT71P8nRxodlDP
sJ7ZEyETOlh6QXeyaaj5AljNRQcM5eoVtfMe8dqGA/Nqrb1tA8jfoVQMnoCqFMj/
x4CfQd8uAsDatYaaxgo7rZkRvsv4lbvVzURGCLGJpTKJpE8tXyEA8eGbdJgF7G2o
EOzHBAsVr9n9DPmklJ/RpinLHyhSnbVb3p5L5ji7Rngbz/hV+ShStP3uxXHP7nXi
dgTiT5gEdLLZiv95URled5CES1EA9mNGLPgMckUp/x2qRGXbALDArlq+153omQjA
Pr9k7fs2yP5kvRGVWtM3TJDQVVratKNJXm1WTgAHM5Ku0soW8LXRYAu4dX/E4rpP
GQcIQ+VASZQVtdzOjnpROBhD3XYx0gKhxE5tq6WAeQ3+iPfgCpepT9vit9eGwSXS
FptNvp06xuvJAJqJ+J5B/CAwxlq6mMGW4z7fTB765UeTYjH1jdAqKDusxhtvr97h
cYZZl28ZwQlb0EsxEEqBfmEWMi5glGezLgreQbBPiOlzvykV5PFa4XXLupVCGtlv
dPMX9omtbaBxIHX9nIODWPkAOkmZYyTEoKrwZsPGzoTj00sOSZ1BGD2w2uauvVeW
sOQ5c6mYE52ZtbZnn4nfVhsemqtfPoOAfbC3DzZVFa2qNKbbOE2cFjsbRfKUIEm7
idX+iP8G23z6CHmDKjrJD+f2FUCbBZj5cFW6SPGuwKAddrgSygnjCIPTKR02gV6e
o7hYnvKzQ5HhZbBQB6edf2+ByEmGwGdK67UuhVnOmM7Bc4wXmnt97bvXNlZswE42
Q9RaRKAavpoJqJ//aMQ1loRYFKxXC9N72kAYLBBCJMg854uNcH4awhwhOcj7nXZk
Y8lRtK3zdWrpwoLo4OoxjFqadxE+xLR8OozyVAE1rvBtFHodIybez2LV9qn7I0eD
BbycCD0+Lss+9OCx3d8lTtrdRIn+BofbpHF1Y0NnxT7HCiDh+TxUwQ2asEXcA5vX
wwbFaF3TGdJv7zKMXSGszmMlkOri0o9UHuNT3ARpdZAZIAQCqhOYukk4wJw/H4Sy
ghYAZJOh208rZv+CD/j4O3DUDIiuPEiaptkx9pJBJYXHzKEktlSN5rIInXXBd8YJ
WQAjD3crSv9NgngP4NpxlapnAL70V96SXAh70cQfvDt0ojBGzs1uaH5Y/6tznHqY
Y1sLrlzyMHrf5jpeN7TOQ5C4R0dK2Zu2od+IBFtGOLYWZvlEbnh+ZyyliJEye97Q
VT2vskJE+kYzxBherGIhCec+s4ibA9vMHKXt12WDqh9w92XfpZ3TwdGh5UvUgQFd
N6WNryK5tzVOPBTG32g7XN7Hu8zij80ilet+NWvkggiHlyC+JmBjQ+LcRDJRLiIZ
00hH1I4rpw6me23OQ/i221YgxuWVtWbKFHyE9XZECXKLQFYAAgzwHrXz277kH2e6
9+EadJ0wqXLD/pfWSiSn8hgUNCSuPdcP6hdtEoi9e9/6yrC2vQDrI6QYOy/CAjCN
gQl04U82dm+3qKnC/H/m48nT67j+nQ5l9CEif01YaMaSN2dJetH4mv4J3IUpQxUg
mJa9E5ogCEXsc5cNrROjhNjP80fvg+rnLhfceRPStzolWhxRP0MBNbGPXMOqajAE
OAOU+faRvmbULTC+Mpw9PbeH+oPrQ03zQRqj0guTf1JuLSC6N7lPrUAH4I8tEJbK
5W9GWdAQhcrXW00WrdZJ0b1rNXU6JCMQGeWCB4WKMIALmyI1WUu/kV+63N7aA/7+
7MZbR1SkgH+8c17d0KJRB/JxdtHKEcE0QICtbRw43/FAWk/0ZfgotDTk/Sn0nfwI
SGRncdKczFCC6EU9tft36Za+E3rQjHT+R0erunMQ3aFpHF86DJv/9Je3KcqqQOpP
LWvkCDfufgt/rEi11KefbyOtJsXM2Cn/zfAlvf1ESMQBXT+KK7w4J20RdbQZ0whV
aV1GHqT/52eeAO9wDGd2mLHO5ighz3jxDW4vSaDSpjDJ+zzG0U1mZKrI8CUhTABF
vlY+jZtb8pDwOGADlxTV8Vo8GklKA6hR4apRP6xCXKu/DoR7vpgZDYIYSen+XL4y
svCTsSMVPtW295uJ9L68RlHpSaex22b97DKuxJPmzy1qxz35+Gdgea7ihWOSXLpb
hkwc7QyevaCom72f2Om2v+KnpXalPOpLBvsvje/2jrnnvyFSBXqImNcv2GsKpMAj
TafDiWS3px7/BLBcsmRfxXXW7rWMpaQaRUorunMOQE5oTzKh10Wkyu+4ejVgHnGX
VvFsNmrUbNKzpGkkKyxzqLiN7Uzp5OWQ5pdvpMS5nVxJB0RZ/2gnWwYQ0qTE9Xt0
cvxpwEklm4OiLV47R5MamqyhenY/U3dk0GY89dQRsv3RXLIsDx2sxaeNcRHFidR1
G9cJJVvANEOnkbC4hBFSHbaDGVHzWwX0SPvRDTek0ZXfABW2p2ln4X0nMKMpNZec
7Z3lX7YbguGNiAK3m+QUPGOYFeBzOnDdqrxQbwrTzuZ4GdSHKF4aQhc8wgx3Tlj+
9W8MQfS8rOm/t3l8txNkSmuqN2NnXn3pUW4RjsSnBeSPvLOUZEELSb0CSuqDZgxk
VNxFuZmToYFMpwIpxp1ok6NTXqIM54J2c4EHgqlOXw9+tM6tF5kaLiYMzUpF2oVt
BYB3lA8dJ8hrGSo6G5GiKFdC03OdzQUTwTIXEfGRFlqeXFRmLU4nVCKKLdAUrONO
pjbbKwIqlViZlKDysEthcogwcgV9mZ09G3GDJU9s3biN63mFOclMnkaPXLmbcksD
RunyFpNd+2RF2k6JrBKH3zW8KpQ6YtX74OZpJgxBFIFA7p+A4SV8WJFwsQS7Mquw
1eMPXJOXUn7QYXK2snRoXo+Mw94VRA3hU4+c5B4o5A+REMBQdVXqQlukVbka2BFf
8KJM9yfbbcbkYXFgnfF3zQ7rXHOhMOC/Wfkxhcjn07pMDBG4WSLhkgo7RdXphDSA
gFmNDMtqOwCUXUw+OWe9S0vB8h5WPGj6xqsoFM1FglV2OfH/VVydghHikStmpBup
RM1RMHCJFSnTD2GRd+AXUBafT1e/NMxWo+EhalS4OwqMeq9eT9AdFRKCiVlTBE8y
vtLHAwbeBdsUTYaEtulEhIMqS78gTkHU1QiFkeMS9ju9EtS0N4fFi7KcNvDReTXd
6hv5f058CUygB6prqwlbGLo0tn71rOXa80xu2/i0+bmzfkG6M6Tyb1klnwm30ygq
d6X3uUf1Rp13pB4HmZjnN+0hxjeO1yDv3gTGDl9hDmMw0nEDJ6KP+gYU5KxDxGpt
MUiUGS5pVxgYEo4gjFnFU6/N9SiKyup5WXfUYrAJTsbTn51zix9xomwY4VRsvu8V
p4Ef0DVipRMehOuNwRrnWBRDJB27oA/rb+pVizfJiXaUtvKJ0gW7c1aAC7WnqzZO
86y/v714i0jwmmyqAX+7mrMHW+buHW1RaUQQ7BLRV20dMalG9vtI+HFSRjNWrJ4G
KvvJgbMTs8C/0kvULUKmUIm9MwOHY37tVyOFjno2oeHiMhnN6lxtcrBwZYo+9iCI
PNgjB6/XvwGURekaCWMcU0fD65iJONJwkUC1XB+ceXEOq64HWeSunwvEFodgWMuV
xbkIiMUotvnKuHVC/gkrR35Ra0+8iN6EAxSIASaFZY4ypptZQAhWZojnOQIIM3zi
TLjvdqpcZHrEEtmYSEtHgTBp92RmHihS1H9pXHwtZaCRnCa5PJzP3nS5sCgTCAR9
pUppRjFxsBRo3k6rMlRTPCMA3hM/8RR/DZcX9MkTOeFsSx4mJGEcAKLDraZbKhVL
Ta2nD+1Mpzqs7CYIfvH72+3CbnObIvuk/m6WiM/CJOMJQti2kTbm0C1EV3jV4Mt/
a7XjH9e038yZVsnfx13YptAZHBKuyygcZXkedoteSj6+ktExfRhDXkm1isosW6si
wPTUDTRasa2HFOKEd1E2PKNNHYblSf0yQaBgE5+fc2A8haZ/R2EsPR7RTXyRjUEx
BSew+RzVY012ZZGz4Oeia7cLvlTpmEvQdz3HCaPTxiM8x1xumu2mI2Zmrx7dFqiY
YnIUBhrQpjvYROwleeRf49y9lwmR2DiJS7RRxuFGVmZun7sZiMacF7EI1ScOGgY/
Xk6XW9XwcSssu+l93nPT3mYyZgRRGKK4KWcy/knmla7+19yByMx1Y2S8b+2CoNXe
LaeIehbpsnPogndOwQushWYnz4TYqA9oXGCotA1965rZI7MefIn17OAdyugFLZ7Z
rJVfOVyYDd8sRAZ8wZ2IwU6zhIi7KRM/ig1zdvoEPQQWedQ4VekZWv0awimYYtUs
qe5NrNdUlq8hiOupF2lWurS8b8Tq2o+HPSEZX9mxiSv+hI8O+uNbcObcDtGIITRA
d7fJ+aOW78UQzydjLAceLB/ytTdTfjQ17CvXGBJJLgwpwv1HNA23R/JmweMOJkmP
JDUlLI9J1bwSDrQj+rwCfr/0emo0MNB5dAAreiEVg46mDVF/7XTveeW6liT8V3oT
VCyg/o9Y7265TJu2ik89EeO2M/rEbXyoM1sYETEpOjnDvf1d3qtv1X6XAkDZHYVO
S2ahoBPxpo3kb4X48612rNViUm6ouxG8sU9Kb8eWI52zGWb2T6BtD7LikRhehPIP
t7Xxlo5ryEUuAWNYbdYaMjBv2bNMtQRJcHFMZbTwYSb4kA4+O2EcuM1IPzPV4gpQ
P6uMdUGr+HTyUZewiTsbvgeK3P4gXLjSQmNzoXacbMHfeRQEExasCRlcsxwK8NDt
EmQC+qDEq83Wj08HsH2QA8V/AISOZ/yR2LnSZyLIWulBemmgIikWLNNssfVQ9kM+
HFPvUjTMsp0uTqjt5hS54N9E7tNyZOl3JGpIWNqP8ANgLhh1DdqSd2XkJ3gj1UWk
J94DsfBpsJDjWilUdIm9AWlECAu9exccdLBaN0AMxtvVk7NjGtCNScCXWGllnqTx
/iitGiDRpZHfFiuLNKSYy445+Z6gG2Jvas19GHXV/hnDIJ3QOti1L4aFv9n55Y0M
5zkW1b32JTC5OLdXIcBXSOTAdwjonhOkYMBYHB5NQRUrk9rzmEYBOxaLg95EF7T9
1OT1uwqpe1Nwv+I5nSTARk+fmA9asV7mbUX9SdofjfskkVnLVzidXzOU9b7Zkg9P
oPmrFBnXdNtOWBLu4Nt9h8TMfyO6usS2xe5+11EKLlk3UsPbzm12HKKJgUbvHlCz
6fIUNYdQAo06Lpb0djLElP9WHk4dRPTCOL+aVn4rlkewGPKqE/QSDwWvDi6UU82b
N4MfUew/qIKt6MDOmAaJt7OjfOll8XfY+2u3OFX5bYWfLW+G+nIco78dL3r8QKSb
NyVfDEr5ZVxxmQKhWfoMr6P8p5Y3cCZV0XD7KF2AO62bg3AEAIFzjRsXZ4x3oQIm
7F8BFXewm1CmGNZ4eSSv9mGega48ggRiFZkZzDmwsDBkcM/osytHuMOC6XZsnR1F
sW1XcbblpWxpNvYv/+bptrtXLj5LZuN6TO7088Eb7WmbWPhZCOMmAdwithmbadTZ
R17IwmAP6eAo+LYMWjN9zNKi8DIz610byPDdg1ctCloJAGoPDKxH1ZGj7rpfHn+r
GCpCXHeHmBwLE/JqzlMs/M/XHT1Dse1e7ha1PWTNXJaadoeOZALEgJO2qppV64Mf
njqpJApoJJY4xb2NidKgB4o4wMPCGnrukMwaeYfm+eZozCLbF52JiyN9UaeNNJKo
4BJceJeoAb3vxBVxP+h4I3hxF0+iq7yWW976waPy/hVrHt1pZJocbDDs2231kJAk
jvLiisFVnWo+d2NaBFAXuIZZpaHiWKd6OrX+JmOVFDId6wv6n8OAzoHn3dITFaLL
P1IypoQcIzVzqDsMMKm1/bahuuQMxl8AqE5Ei57Khac4CU3CLVEEqmElI1ce66vX
TH9+2vhLZ/nKsbvjtS6NhJ39NQgcZs7E4LCu2PI4mG+NFfjH3JvTMx7h/JVCDXUh
TLXXswbIJixri+PN8sCYvVkHvY15o5He+afZkD6WyawbI0J17Fk/GnfvPFaEsLPR
S9RdUR9RWEn+1dA8zD9fkAQAS9WFu0zjj+QdBI4jvUoTwDcvJGG0R+HTmQsdEAe/
wRutIAL4OC+oO1dh2FwUyg9+/tq8u5p8msG5jKz/aUU1IXYUq3jjRwV7Fgw3YgAM
odhdTpz9Acw436HoiN6ZdB1vaF6QGyJbnxQj/xWIU5EUD5Zi5+atJ32JSYGIRaTs
Pb5QWlT5WJXyQ6q6s8Vd3jSfniPYwY8sHpakQlL9pFS/bmuyilY49++WobR0ePOV
EjkEHvHn4Ng+YBwT0X9xojCBlLBWmstMEXuiclFgyh0IVGaQgi2gfdhdAevrKvnR
dsiMlNVP/SYRgavQB5hKRmE1TjwpvHE7r4xFXxbqFD7524YkgrY8mkzZqwIu7Y80
VBckU9nx8HIsgcUmM33FGytVxyz5hwyMxF3eQFGXqNDNCIpfvUvi28kmkupao/dQ
md0CPpOJ8aiCKSGobo/AjRx9WwTlvB4I7SRQS8hX9ZqiOagOSHjRfX100KGPlB7T
NI6dex1sSUNdh3HNK9gOSC13szzBbe2ETgEVdYI47hcR1JYfE9Tr5VI6g0/mQN/G
MyQkkTFSst1ep3/Bi14/UcWCdp4W5G2is/PiBSr+CoNVVDig6CS2rvV5O3iREPfX
S3vd2AeCNoX3r9Db1iXNyL8VC3DDHVfBQzidxFic7d3HfpIp7jbvUzHXl+ft8avD
k7lmMsJrhi4l29zgXKLFYnn9tG08FDIFW+oiSre9es+m+7/eBWksjXC+h3S+O2E8
WsEbtHeJXVXvMMIQF/Fe4EddnF7TC2RlO2rNYchoA2Qf0kmBPFa02JEc8q/dc34w
XJu7nbMNsQq7VxCbgeaDu5nxJoHoXo7rce/eRpDx2qVud48xBRqS4NLDjjFF7C/5
l1/gS8lgsdhCYhcnyNI30xyN2Myr1XkHjjMWLFQk1WkGr1eG/h5T5b6K9DGTqewt
upMHleuj1E2PTp57u3E5zLKjT59UFqRE0LOm90f6hwdhiuC/P7AS8j6gG4EF2lEf
xlr99btHdVGeBecT/r1dPMxBy+6nFXtweY8LiH5y+g+d0ea80rd1nxM6A36hXfIr
geTXgMmXe+e7IPg11hAPYtRVR/RGA30ZDwVU53lG+DoPkkBcbzckvVWwGwcfgPsv
j7v9fVCu6lpgPCyQdVztoHygifyHC3ie7JITOsKmF6bm8pNVzZaCqVBhWSVQErRF
XHQxmrgjTeTw8UX4eCWXRjvvSb/SbIeZ0JuwANVDtFzsNgC8Am1L6VrqM1Zq/HLF
7yI30HG82mb3npCwdiBDy9DzmD7zqobULl4QdlI9lvAK+CinzdmPAYHH6HmgWkR/
9tVITZ318DLqD7HGNNrlBX0fRlVw/j6KRVtzG66ci+96aCnqasuZgYAT/X2guDu2
XIGVV0ldLboN+6F/ZwFhajzfW92z4nMeGji6c6h7DYPA7rZuLN8/Jy19+MUIcvvk
9mxakdPjdabTkA9t9eBJ4jaZFSPoI6wfRZtkJ32GCYHeupfs1xOOqncHNUNq2cnF
/Iluyz4t00S6kPGXQfTaYvIFpZFcbp3RPoyJNsIyI7lH5RBwQTnwzEziFrXP2TVJ
HG2tYKx82nXG8rYqyMzBrLHWYuzm2Vh/G8291dKlfe/FfrJVoAR56p+CB2BHHZZ2
Mb7dqyX8f3/pJZPmWmolh0po/uS1iDqdwSDjZChJS70OP7KPF+YCQxwdGmB8+/og
IpOJMlXoIvZdISIcAgMr68OjErr9Q4UX05+zk8hZedCBDn/QYcYaVPX0ZBIWy3Q4
x5ezzvg+YvF0HTBWQlRasKJk2s2P785OMxs2fqQYl3U/3QESyt6vKI7V6d9gYgxC
Fln7asQzLD9P2iDjDGRWXfNKguBaOLvzVaTDLekrpX61hRpmuYwHRdvwuwqfmkp+
bSrsG7QriJX/jUi87mf7A1mAGEz03saj3sut3TELpidMi+/kQQ3iAuT2DM0Kj6IY
EtoPFVGGPOAMA7/nD4Px03Zn3//81nhSz8Eu6gzio2AZH2KZ9hYAwv29Kn98CZvK
s5dFJLZ8Yf2ww08BB750s1qB/eunSCzwEhOXE4M95oNBaDjW2tFlqhYYBolfOjeV
zzYrKjWLakDK6js0HW5eURUMCn80zuZX6vKFMBYbluxRmQYQ9akJL2zEqNRDojsv
bPHYS8Gm/G1TBq/0IGIhfOTBQsuox6pvXjbIv20UDqFmRVIBoD3ZYJeSC3u735FU
IeqxXmoGkGUd3Wym3+pwmSmvXSiPrcrLyGrkmUJ0kTOv1/UN3211mFweElzNrSt8
m/EkeA1BL86FvTB/EbwsTrDPJmMrlnC7/dxrZ830HRu1z1bd5La9k9zsd6ffARY5
Qnm1BRA4nwv926tUlV5QMYBcaHEVsVUEpQoJGdcoQihmFRSY3qKImYOFTXTAFWxu
oxU/cc6HZQpjjCzH2jb/N6IaOy3kG3WKSYHQC+a/4+L+NuOsoLditwVzMAxskgpp
KB0eoxTtYqtRU7541GBQoAMqMCtyE05IGDYk3XasiNB/peKbimu3f3OQAnfCrQdJ
wbtjfUf60oysOpB2A8Y2HSqSxWzX605kPP7v39xMcOmhAr9HWwrIs4w4lR87330H
EFnUC0UBfcNua20D0rS689t/rSbdMlsVay5UR5eE1jZUSV6/7Rkaqth2rcFq+++M
7fRiZoVokys6gYBY4LhPTuzQ+aNfBxOFEhgDB6VWSyYsZXrdcOn6O4AwKweIkh83
a1+z+1syf3qtQ6QO+AUQ6gJ0Qmw25o+ABfd7HHliLdF7l9eLfs0xPw9DhSg9P95D
mjo6sQmUmjPiHZ8Y7hOgYZMddLK87BkXsnj0BbnI8rtmESiMdkfMA3YC3iPNbDjf
uifOwXECOR2CGrX9OkD1PH5yR+6cNaKAwbz2HCw1jb7ngu9l36r6Uk8OzMMHscLJ
Buse6hAzpvWhBUH9HmjsKUFLXFTukOgh9pVD0OSMIJR8hQyqXuSy40Dsq9VivjQR
ymoKvSq0vlKmUTVpDcZ9re1jyX3lx20oipM4Oig322U1QEylc+VJqim7nBjkwAdt
TKcUXZZZ3Yq6pf36vQoDVgwQi9d2I0L1Ko7fF9QixvYnQ6qjZaHH0TznJjeDEbY8
w6CTwkkaspP92ifpwg81bSp+JHzhT0lXPbqfop9nWiTEEzuj5tMZhRknGyGIVXws
JnNd+zFW563JVdZG/Tio35qiNBr+Cs2Z8dSEJZxpkAQ9qtWsF6hXpAZTgn0txarO
lIA02BuBZh0L1RQJwQaRz+dXzPIPrRZMC7i9ntFapT3B07+EPYdps4StQbpF0lWD
CPmRD+GYTcu8WZ90h8WQYf8wO/l51sCMSebJ/koNcGxpBBvTAX1EpwEUl+oXbwFz
mzzGxlx1j1PAy/jpfhEYyPVRQfZmw4GRoZSsvl2TbnOtb2/a+HZ2ceDJsnblY+kq
l+X1MLL0w6phpZpuP6j1FuglvzT4lFlPRH5OXZXLgRpjgjn4qeAY87R1VuBuIAzd
ZgXP/HYQlanD1CWFuvX8VKpCmiv1Y1abVV5S9OJfTke6Yt7y6OJvZ/X5IeIYsxcC
9FIPLDK3olKFLeSY2wnnGs5AJJBd15PSEPuq7ZYXjbObuwrWbK8LdDtM15z8CpBH
ZSyOC0esnBizVLiTXFHTZLbyyD9xOakP6ZcOURL/dXJzOaOZAlnuxd+4OTq4iv0x
H99QUWJ67f/f2pksPlkZAQ8t2rhaiP1aJ6jRA352Mi2Nx7DIWUXdY1z7umKeEDRn
+gr45nf2aFxW5i4xdhR6tqpoal/4oURa1QXJsV6FQqicdZkIxYHSFWWTOJbisB/J
ek8kifyWiFuyF1svqIVA3+0Q7xdQOjFzV66U3E5xQjyo6GanSa+RxlXpvrJ6/3F3
zKwN/oJyLWcBhSfbmsCIogbE7VI3kB13iuhFhAK3KY9vCYli1/5Kn6MF0z/r0R3M
uOEaRsKjSUR+ykjK0WWsVip1bbhx0NUnlY64NWqH0ULzVltcZPChrKeW9xzkiQ/d
j1o29SnFuFEkmp7bUTf/mSgY/AxNRWld2UcTObGFYy4YDJ1uUgyNPsHvt8T4gDNx
83Isx3eVVuW3pvsRZKYQ2B3FCnZmROVK/Mynoj6K7fFsk54who4rGxBdKnDjRj34
7sO/O13PxewuhecsCmWxiDPlUnG8mUY8ultd6f4Wp/Nn8ynRQ7gX2eznqiQd8JCb
SobXTUZbI9S0ytue6GSEU5VvbBdRi7VdKMdluAM+1PQS7NnVfsACq0A4MrIbEtj+
al8QIY3FFd4I/SuLjrlJwmrf5wdo0IndxzTM3hJHE7ZoK6W2z/dxShE3gZacIBYG
PjN+m3nSBMgQiWpgU+HRMxAKb7FlZKp04TuTfkUrVRBgayX/kebwCZ8ZRJwJ+n44
KceQGj+vD7yZCaekhhB/RieQa/81YE4pPhH+E48wi6HWUUSHfe0LKMbcPj4NMl3Z
szLGVqlvn/WwSmG0I+g48YwVoC5X/tqh5NicHDmsJQYYsnPfs8qh3JLIgH1eVvvN
+4YUx3MEgiFqX+rf1F0ZtWGStnQkjbgMDUPo0cQDbiYYEjOXRt2ILzsCeJLSP7Jv
CmLoTswWUSPO0arfGsydFVcgSqN4XT2w0WiEg/BHDlJkcWKd8zRbiUIoU5PzaJP9
3HgfI6JsbuQxihuKDLq/wn3+9WwlMEKY5rXAp2qBtuJokGpaLrwPkLJB64XlldcY
rPDx5vIP/69dwC8py7I+P75SctrsxzSLoPFfdgX+lhyXE1SuzG2vWaXkDjnXynxw
GfeVrXAkTYmHg1oHBzdiRflecbichxGZlB1C3ADu7TK1V3XtNWE9v9pRpS2aiChg
ZuHa3MGZvPNAaRHGXvK9NRcBx59psoLiyHHK4MNugkMxkQHsNYi4jhsX7gJn30qh
E5/QFTUMbWSNqTeOmcCyXwLXW9z8MQUR6+fz6WBbdrzb9s9h9kBPMg1zQGtfbfNF
vm2yKvfeWBB/ZZs/DEqMrUM1ZQDBVVfA1JQJi8VumhyKQYsOFeG65OJ6Efm0xbvJ
1TfnVCaTenPs7DhrkYG0+TYOo4iT3DsjvyYan+bRDuPyfKq2GjfMK0a3w3NGt0ee
0YGkonZ+/lBNWsCrmfQl4Gkp8hfPi5sDxqUFi3wHGYqOiplmxmjIvnW/cFYzeDKW
i/F8ALPAPqD8FXXuxXpCwB3gI5P1gLszNmVR+EOPrN1UR8nlNNi+65oJfNXdqXlj
E6b988P1hKhxcbK/7GOXOfqJjux+BWALbravNTm2ukVd64rW7fofeXRzc2LrHJWq
M3lXHVDQ8NTiqp7/XtRf15Miv+ApUYDz10YY6sFoFDYFFnuUnXVdaH2in36h+MzV
KcKZd6a3gN/XEzRQTKPFPUZPmrU4gB107b8YikRbU8uE+FHOCeTTbfN1TGEKVZQs
2M1ZwGdOSMHmNjA5/14vc0hXYxmptlqHKkiyzjpMw8/6EA2qXkoHd8TPn8hMV5cT
iRgFxYI70vigukkSX1cscWrJUTjPvDo8EsXeoG+tiRBu8r4pVTD7py+wZ3S2yH63
Dj/+TCV/h5Vz3hGwGtgiw5kqZBRZIY2LsyeHC3XqrYs7A/hhr/gBWUP31JI1V5yj
0RS7PM/0nXg7MMxBtMNQDGDESUxx/b/V6DcTP2PJANG/CUCBKWYP0OHKa5AIXpSw
JumdKlE6JnaC6ZKxOZQhaU018AJmi2pQ7LkiBy4D0r8lAf46w2GXP0hXpsFmkEEn
cWfR+40qzZ/lQAppQh7jcEl9ubqWuevlMz1RvXFuMcqJdeEio/tUy28IwoLg0JDc
Y2fyWP5CNXmsq+oJk+wlYR2X4QD+bpFljk3oMFivqD1+hQxvpZXc5a76L8UV79/S
h23PrU9Gyi3+arPQJbZvw1DGUenQd8kL3G4uVA73iCmM0dguSmxSr0SzOHNfM3bz
949yDemf8UmGNU7/m1NB2Yevzu9MJ8mBKte46bciTFYPl52nWLXCNmDe+C0qIX0n
k2PHQV8t2SSTIGfSG36uV+oVA7P1YAZiYmDYA4EQGEi1b3esSH67/9MJhuS8d8Hh
ddpvgIInmwkKAP5cUQd8jVVZDvuoPr2F/gvN1JZJPlKyXrGcrtS7A/EAV0jbijVb
ntdNvZKQVUQW9bcIYFY+hek5cnQPQEw5nqinNmnos5wp7i5FjcoR1wYxgD4hfhDP
4ml5qxHZFwzn5ztiRu+jV196RsZb5fKhFNVqPly346R2RV8OR3X2vc14/aEWBKrE
Pw/8lf50vSo0edZZaYVyHGVGqVXJVO4YgmdGmtH9jUB28BtM4wj8bhJOIVTXA9aS
mDUkrwz79Lfb0QzUTbJNfPhjzApGzPKiIS3YiXTUpvgV0agTxCvLgjHLjkO/zI4v
3esArDlL18YJCLuvRLuwU7rJKGqiriNFsbTq9/jy8atZzRq7W+QvCMXXmszofRWJ
66uno0hu4JrXohw40YBxIWoZ/R3g+LXM6N3qZvZxRZpmTJ6AkXZZH6IPvsYM4Dpw
asAkB1GGZG+wzjiuaCysdsnfB1zLED5ct0RUaSg0jSokf3GdzSVQoD9AGgCrKci3
x7yphwM4rUtWJGLY9uwyHTF2OoAd3xbu66G9M06jOm6WZy8sf62arlv9Z0hWCpu1
ZWpOICtHgWunK5kQTPi/D9IIcNoualc8OuoWMJbumocYxsaOOmWW7+3xieOLpFY9
bgTCp/YbP9uYqWDVafO8iWN3OOugkdPs9IueVGXEHmDYXyGSPHd7PJDNXbjnMoxH
7iAPW6bP3459ReB5DDvd6jo/3tkJG4dcjxHeWwOxNYx05Ax8TDzu7i7WjsNMORie
vHzfQJLzwlJQrbigNlQzERHG90/JtJcJvYjeuczKIDFNezXwJwUQWSVuj1ZaXSd8
nnXWDMc2iVLmWCWMregmW2mecfBleRLPe+CPXdisE+fgnVqSSvduST7t8WSCwDuD
4ol4cuV1pg9wNISlczFiyZP5RrZvcYqm414e7eci/e3QDSdH+MLNQsrF5S8sI+tL
yV9K/83VpVGEoN9djWgQwSXVzGoJbXRIu0SBbsGVnzri8y1INOkcFY1O6HqPTGqo
PgZoWN3FrqZ5lNCAgrHsx/qScGr6F5bewb3efxI3ZTLn34gtdd6tz6PfmvpdBBgB
uxiMpBGgix2f40BStpt9jSg9jQEU1G16bRPEoS43q1bDZZaruw7ZtjS9nIA0aqZN
LDakNUE/wj/VpHXxJrgKm+Yp5GkGBsOHmif2oypJX05dZT8DReudWphufbjSXpI0
WIWD4vDkTMPJsVXbsk1omF2lCxvyKAKjlLxvVHGD1HpAQj4PLufg7JBk2YBXfDKf
cFhDa24wQwk9ay+mlJqbEcylbFbDARJeA7ViGV2vichPesxVVwCo537t4r8Yzczg
jfZMOMOyC92EnhUrLwLG16pGtaesDoT6zquo5Q/zChMSLF6Hw+gctNK0XRIKgRnl
vHUvA2LZG45oe6dWdevJ2p5Y91EP9Rj2mg1Ctw0ayn0XcVJRMJNwJsj7KrhrlTUV
un5mQr7TpqeXtvO5r9J16WFLJMkx68f1f4cASvPrHqMnO6JaobOAxmumrnid/118
XeUDy9bjHx/aces4fW0EvteZtboecuLmWVfT+nU6Pf3NSHlaNTrr2coludSPkSIs
Ka5zTHGp6E/LHNyq2SfENzW5gwlCXHYOpjY7gja4PWUYS9t0gBdjvPwXDSfSRc3g
xCC8WePGPfy/DYGRK401FHZnOaz9NlhirkhSkcafksNO5oKj3hIdG378Jc99tl7r
zIZMG0nNyI4EnL/fL4sJGtSBCoIBsIau0yGXznQVPZDX/2cgIJcapCNyUB2cNs+N
s0uwQgCeKbV2N5qphO2FhaA7Fz8oLrjbT6qFdn0+K/5izGgvRIlVJ0EOiQy4XXDp
E230i6mlo+J40HobnjKE89wQPIEXt41eEFWIhwUQeIUwRzZ9WwOM/CUmDdJ5kLI5
172PanSk4A3h3qwzqIZLCPkhwpPyvKOzbyReBoXlZLfdHnvuYJwxIJwvzupp1E1s
0nI6oTk4pgqNGN6Tg+Ib5R4mTocOo57F7J9uA/diS0vb/vk295xXCBjkSqXxMUQh
/pUkhMkSXAFyzihV9aokxIu5s9uLX/vPQsk7K+Ja9yrqDLKOsa6sZ3Qwbvm/ZYRQ
IQ2YJXMXTs7tujLpVhusd2D8ijT41E+khCOVdKozANPTGqUCK1HcHwg/AoHWhDb2
Gka0dhvsRuwQy5U2uLUxrroGhzFekh8BAmC1j01j5FrwYA3bXDWv0iSJtmffBWKm
b29DkWS+iygI+aFxTLg6vtbCdxfxkla2sPWUpo5jU2EGCsChTtNrC/I8m0cz3Bya
XaYiQWfKH8fnKl2lnwzyKeQp5S6BM1Z5tNVENUzAAdVWvHNs5E6tQRcxbITJidrC
ILOUSn3abpq8YIe/dbwf0rMO/v2YxdG+Eth1cTP47KxcVKHVZ8JBv/a0khkdwtsi
yKSqazMnUXrK5ZMwFjoQER6JJhTY2TexFjANNtumEICUlbc29YcKola1jhtt0ahp
wfBIBdjUtf5Afd64n+ScKzDA3JNAjE8hFLRJmvDAFXuxHW3uQTnQjkgRgbwAsMJe
EFvdIqDF2bVKUKFK6besPPuZj00pf4UXM/dPd8ICXz8IiHX7KLgoWb4FdvzY47JD
dIdDJEp8Af+ycJfe3ct0nL8J9qnuYNZYEqqBryF51P9/+Uci+ynzFiagyKnwpERp
uc+1ZP8m+Fh6MCxdH8tnb22EbLU1GJLHYvcC9V1S64fk1w1my8D5ytZf/uBGAGUW
BRxqCnIKDCIW0W1HMBgmDNdykKJoF+wk9pKjzQptJ6fowGeeybZhMqj9n4sxA+3L
9eng6pw4zv86PPdZTXBK0faI3G0pphzmJg0bQoaKZKlT+hbwRSVdv0DPIzQXHvpN
X5qfjbEe9tJ7AMyQNMnuLtFUX1ZMmcVRiNls/KwWQREWXigmi321ILcMXgEsUXVm
LVJ+dVNCLZgrYOq3zkvzH8/qKxDT5dwyGe8uwN9ZnIihimu/Z/sXgMnNptf6uzkW
zCWh5dERyKlh64Zm8FQWE/yVkOdCqaYGNsd2l41gCpFsFq+ERGv6nKvbb4hKPbUs
TksNnRpGiIn5pCWsExpycbaYWPnCA2/ALFlsxoHpnU8BxuT8KicDjXT5UUfqn00u
nqB/dzzt6tYKSoHomUDeTgAZ25LkNTkLqy7tX1YlqtQdPTWo6by/gtUhnjGr/dJU
PMfuGNgh6751tz6GcXy6LGDWGkGDuM0km4xYwUKGlTR8zllKCuUqmNERaGBeBLJH
7NWujZzQLhx3JIFlM9Vj0ZsfHsJyfeDbfAT6DLaKKX5WicD6ZoYTH1YxtPGbNedg
gbBhYiO5VAms342VFKBS3lTG2bS7V1iroxC+g1R0sweTrzpn6ij1b3/EAsGzfZnR
KMk/oTthpD8OyY53hTWvMW2WaIQgoZYrVq9ketYKxa16NpS/TM7WdKw68RB0kVP+
YFAxx52gQDsTBn9sPaOhpMWOxJPCvpXRw1rnMWDOx0Ta10QnbG1CZR4RAkJmToBA
NnkVhGFbDsGFxueyi58M1q+/OQfyVC3S/SGiBzLHztJR1mN+PrmqejFA+/BbO+l4
jPRWxQGc4KeRtAR/nhA4fkH36kOQw1ushJoZRrJaUWO3XgzcTWS2l10uNSPu37nE
CeBn2SApYuw6eRU1koBT+4Skxh4WSDFhEnFu9Ip8lZWE2jt+bw+Pk//IoZ4WZFC+
Pxe7JvXYRGDDZJviZAYE4pGiPlpuegmCZQCGSdwqxhExi3clnRJ1VrPsYsS3yP2v
f4Pr9Krgv2wd6nL+rhsRVL8kCFcsCGbc5FRynQfk2Rt2lLIDhL//mFXAHsOWPq7x
qdJUtqF3HqTv1Rrd/GPgyjmHZVdQ7wkAj9X8+B1sMpbQkubcz80D2nu6/bs91vaS
1JW/hO9RDnNWpRVpKWlA+ZpltL++5I33RQp4fS6bwEjV8StRHEgkoA9LSLpGGtxW
9hm2lrUw76qs7PPic8Fm1Y3zJD0XlRY/O08WKiDYMbCJKPT2rdOiOFoRB3JZHIyc
Y4Z3s0caqraAQ7IFlRCaqTtXdovsH2Ze9rNkPh/EGYiBheipSG8PXt9mANJ0DV+J
lVxz2ssMSyxZbeWHEK5W7/qyDHYMTBrr0TsySaJ3thp2mtyi+ML5aPm5EdHhrdtW
axO9frsb4ghVmvBQpcDcbWUu6FAaATZ/k6wOgVT4mDZMKeS/r0+meFb7WOrYATUu
xfX0gUfb2xzth7meLhjnp4iswYMPlR1WnEs4F5pUjUE0UpIxwz+3sLa0ikjQa+It
vvkCAGookTIKQETfHsHvwcLnS4d6SWtBOPdFBd+Kv5H5LDejmrwCeOCHMqNR/HRh
WowGuoHfNTKOjq43Su+lk/D2lIeeQhsDVuqwsHdxO/l53rWox+avTOeNedR+fi3f
tAGgQKWRBAPdBu76VVDucGeOYUAFfJwn51u1ElkbsueWfBB1L76WYkpsl5f1GHfZ
VXPAMU3q53Zu5eCFLhX7xw==
`pragma protect end_protected
