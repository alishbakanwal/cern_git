// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:41 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oN/6sQZDiJJ4aweaV7IGJHn5nsa8pqKm++VjUk5zN29XvDMhSeZTDkcIs5n61AAd
bakumWJUVvbAZLVp/hNkHAXY462Ku/4GopiytDsc0IIE1Dw7WI2440/pdLpyh6Vi
H+KpadkSgtfULC2Td5uckVAmg63x2cMEmqslUAzJNoQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28624)
CURSsxpTX0eW4DQ1+IYZUkBEwss52RMtL/+9scfU/3nn5vOYT3t5Y9sLm/676QNR
PgqMDlOseMDg4uQcehjtQZtEYxdFSXktPGSBuQuvpBiPcfrte6mhBHvjcgO3YkyN
w2HR9PuF3vdvDw93eAmMAYwiwT7Y5R1aIcEyUBeD64hZQpR41kWiDRN4ZqzuIJdU
KpknAPJrnJV/qitdQHvlrcKSg/h5FiWEfVT6LgbsBYKsR7JZIlSTun6Ng0wo6CZY
q/vdyRu+wGLgjfl7qoGBePxuRcpAkz47rmW9HcCKL2app7PXQn6KccfjEf7ZkTwj
qauziZCNpmuwsPwZPS4DISaGunpUcFQW3376iUx0FzqVskGu3coJ/P7OKUnYxAtL
52Vokoma5y4R7dXpYMnqm2XGlkPfO6SrxYRZGSd/pUvgya2IuvbvL3E2JQMCG4Ky
IEkbXD+7ODbHKCWvjhGaNiMOe/QLxM5qxg/wy86JdmQJspGY7ldmJH/hLsVHaXYl
DOreyRIbhcuYws3guGm2wu1thx+Hued6Z5JwNUic/OS3ME6oyGFMC73Trgllenso
qgWVc+UWRT4k6/Wjl5XzqEJOw7Lb6D4O/wux8BTn2dsdy0r55SW90IK958YGnfzc
WrSHFSR6C9iAAu/FHK100UuPCDtUcIMpwY+zauCSvmS8ViPugFlasS8P/c5LYMyp
WrezHXTBVw6kVNG3O2tSrsVoEWLjhq3G8fbGWEtATv01Y2lhJdHjEycvrcG1ISYE
VYbZ3Jx3QV/puIkeCMZtIw86jx/IFvHzO2WqZi0Uwm/r8jooRYqasDYBBU3wK1Mu
TMrE5CmGr8qFYmWO3yJbG+DNBwQuR+fr3Ud/q5d5K/133A3Tep0Yp8vkxgsg7aBs
DavRhdMiXwM9eP9jTIhxUkRAklZoZhxMCO8BsWXDpy7J0kz9cAPeFUs0CUrWFFCN
Xmb8uBEo+GGy68U/8u1HiJs5ueDirfffJmX9gYni/QT5xF7XMKnVX2YtTt5i6KbE
pbl7w6FLEEb8mZdxrICsB2HjmqNBqEoidHDAExLAXgmQyK79VH+0nhqF0OFZ3HqA
VKVyqkWl1KPE38Ngh5MSgUKV10QIrIZhu2fADVY4koxcWGn5hSJ3k7ptuihfMnRx
cMZGjW+DrlV87UM2RZ37iDzI7OpzrBPkFS0tHqnfBBYbPvThjFLHi1Wv0NfEsZfF
VYIoxSuz0fxymLLG97XZ+TdoTjFnXpYjsTxmXdiEnit0pl0ImvGx3T4P46UvBcth
wEJfBjD60ORfkT41OdWsi6AcvDa/RepDs7kHXjrymOuGmHlx4gP9TjR0zDY8JHpu
jNzbeSN0js6V/Y4y/S1JEIICiuIMzHMg06NsuwaVA/DhljA2s5esRp0Bi0B1L6y9
bMwbNfyZZwqtFrWSikTpbVVKycrwjx5ZmrR6HUxqOMWUl2GZYVCm2etqnrm9J0H8
/MMtgrRrjmn/RkUtNahqUDxKIonucprnVZ8+jyM99/CEhkfpDAuDJFRmeFxbDDlk
Asb1KY9ltOjZ4Piix1gUz43sXB77LEzen+sdMJ0AQluv+i7OTQT82CJYQqp/aSfo
qCWjKDX5r8fmRAstC0cMOizeKP3BTLdpGcxyjLNL9qZmkgdCPb1VSkXbxXwMqOYY
N0LTC1/Kx63KeYY2vabJEm2+3kFWtUo2NyW9qgynDMe3Tbo1KEm9wOXGSQknj0ts
vhxlzKA+K9DI9Q3dKoyHdSqx71oM/rhnYMewDC/fxNyDZH4SXxDJF1cOi2MsPFJj
D68ylRQN2WnjpAG3PSV+aDpsCtH9M2Q7pelHKlvvzoZOb0O7PkofKUoD8zeSVNH9
CrtDD/of0/AACz+3cfeAaOZAqQy9KL4b5X3etJY0AnnB07VvaFE5Am76ffxfTzjy
MhfhSx2xuMdMTt8SY1QStpdV1E04CsUe01IzFU4x6faJ9523SFvdpJm2FvLJId2D
h0IrsbZwRFZIQwXPr8OC03QFIAsZrHqjVGlNPcjUdKQFli3c4YcGogsByoPQ2XWr
jSgdsr6/1ZbiclBPXMT33kQ8FF5CcKkG/nuvLRO2+MPIw2LwESyUL8jp/RPTPBFG
dPXbqiILW1ru6atXC8lGIE0dhX5QTIjujgG9qnzGX3kRfVibxEFu7GM1/QZbdv6h
OzH5XmO2TgMFBwcmAJhWRvQGbUaRn0/5TLamv4RVYWD7xCbgFjI62qFxP0DtEJFG
wDG90LetwVZnKmmqHGgCKq7I4ncTBkRE3ExahZWEvuhR1cZws14+Uz2rt7FmeObf
nlt06xg2h1GNbSjvKMMD3paLCsxHr9PeXxDrPFeVhcYsjdPzqLQlffg9w0Lj8FI4
KPrh/1KQ+rGPJYUFWz0Q68SAI8pNbpdDxrCgMFJrD9fAzjKlckOQQJrBF9tPVt3t
WBXDrnm9FWZHI22CLY+n850OMrn9qrGJX4h6zLjLBIT+nhVNTS/0cEnfWu19Jeeq
+rTDjsQ3qqZ9thmk2vyGNdkwC4apHCJudOzc39TAcXdYPOUtxgaqS/iyUp4wN7sY
ka8X/LK62d9b82ih7Xu0gLjG1mUWi6By0S6mVN7dSKS2qbzx/EmI58DeeQa8zpSq
y6XqKYdRMhIasmeEUHmVn7v4wzn8F63pRmr4yxYMKu8IqOyty/X3bKCwlBZ/s2hz
4ETDOqroAo5LZwe7rV8lrrWSmEwTYKia+x4GFEa9nLDPVgcNEQyoNRHLwN+dS/pM
AarM6p4rFhW0zajZzvZTAY67c3buTc5S/e2ydANi+2c8GVjCdGaXAz1HRQVuc85i
20D3DlBA185/41aRNXCZmhH7BGuIW80WvTWk+Oe/Y3QDLXU+TrpjY5pORv7Jxz3V
4QULYpBGevXW0DnNNWQza1CCvMeGgYgzzI2P4C4JxQCdYsudpcDlEMSwcT/3T4aR
mWRyJ7obuZmrDKc5DXD4oq6333/FRyWAOXG0gsosRfja/MdK28WE2+WTDb6fZxRp
jzCoQKVhRyuIWqECOB2AbmnwYmu4ovlV+n60acg1Yv2FmLt1bpbSKhy4EkT9aIPj
6iMPT2O9HgQo/TriRlhf9OGKNWEryUadZ9jbvAvb1Uela3kXIW6m+bD3I6BgV/1F
5CPmcN89+ewwsRsSsmEi/dNFqzv6BUqOyJDDy0BOl1YkRkDtgMplSfkYu0CnSkK9
GY2bLoKk6L54nwl4a0ukyLia4nlAZedrAVhNGAhu3UKcDZ5eS4iIr2dTgiSQneey
VjXFPQbJgnGapPmCWjvSJWV1gJrB8TxPZZ5etTYZFo9Vr44LSIK4gFk9fT7o8ku3
dvnxnCbONeNFCcuhJtGBfI0tfpQGWmEXsuJPs4wvIMjlB8AUDBZv/CXjZD23fnEh
FAQbEv3/NCfrAmyNKicPc5kvIXEZ7QPnx6GUcf+vnwaafxUR1CjiyrZfe8b2FOA9
VmlEeTzjRpTmt+6fdZfkrY4LjN38RknG2epY1eB13aWI/RXzwSFnJc7Yo5AAIRMd
wAnogrhtmEr9Fvy9Get2DyWzMVFoYcEaf0zoYfSMwyKFPT4hLAPM+jXTbCAPoFRm
U5jMoCYxjuj8AnGG00oI0p0QYu5Y2TR18CVtsP1iH3isbC4XBBQFC2M9idpuqfnU
kxglCO9EQ4PqdbR+SSmWNkXdcrXknU2cif0/KdkzRaxjZ4qpzq/6YIkSFrcqf6Js
sSdZm5zQf1eX75bsXxPBEnXRjvm2GDB1gREeX0eFCGroxe5gg126HXCovjSBtgsZ
h7sbThV3poUne5DjvlAtwg9niXif+ahTE1UGqwbycFkbxbhrjxv9j62laKkA2XZ7
DoP/p7j5y6NwW+P4ANgoSaV8HOrcWoPHp0YXABikhWEiTRJv7rT8riblfyi32c8J
hoeFlbD5B89OUAJt/vL0GjheqqfhDPdR5xbRap+N7boSJP6VG1fqYK26PuBLQx5L
a42KfRXMbPD3rW3RI43c+529WWLCIaRJZuadFp8IU11CCNvg33ZR9+svb7uVGxqA
aE/rkMtkSyazcdjl1OGWX3WjEI6E0m4FRCpf+1JxTfwrmIfoe9wtDh0kw5QOaVFB
X5HMlCR4sPlAWzq9rvSN+UrbYNKtL+yD84t6GTqDktRbshxJfPVXLnCYI10ZOFby
KZ0CeA5Ei0vfWe3PFd100e4ZKFUMb3JpjaJ6LNGxkkcWKUSSr52HNjTP4asun+8I
nC16mwjQug+Xp4ZSSjWsQItNF96s9rzvtaUq0sYsLm6Iu+GC+HP4iMbRIOWeMTBo
cUnSD4xwYA7Mkha9fEZZTwydLeqYTpbbQpqC6zIMi6NN93BW1be2iTvMI4MdB+VN
3tWmsePJDumCiHeLaJoo9R4BcfOUdhbKNLcsceTJoNobOyVAK4B0OA/dSMnJd+Ty
n7Y+v/hznWwlwzk7nfwzgnLGV1S/mDqdVjseYOVLYCo86uEXP/mKjp3XcLVQXwaq
rkMDno++B6OJxLLN2Uj2WevR7T6DVjKaLVvR8kzqv+AjOJ8MLBVbazG042+JogXt
IPMMeg9tKyMOyKNOLpF4A7FXwHccpqsGzDWZe5wQ60HNKk0Hug66QNq9jVezaWJ0
kWY6l0rk6ieNNuGE7UdnUuyNsze5wdYy65Y3qG6UtpZs0bLVNxeb/H+kanRkpeTf
iWUZ+SAHFJAV0yH+XNzNf2tTHBzif6hwgsLBG8kCJIqkqInuTlu01Dd69cFft1Sr
7W91DwR/Yz4Fl3WgdEXaFEZLviRCMupeXoXSvKhUcuUkUQViwcRRTmWNMl7kcqDV
dFnGy6KWWFvtI4MRvdg/xb+GF5s/4sCJGaI1yto3ITd8d78MvSU8A1fBMdjVBQVU
5wAFJftr1BPK1xqP2gh583ACRcf2KxR0pCDKSPjituX86LPPGvx3T1HW+F9+jgdr
J3nmbhfQvbgkkmY3+0Xbq8IFhND2BuEiUpvjac4xzJN0oEyUsIsUdHCI4ihAYI1d
vY5R7c+jxeRyXMBfwf6Sn3FsdYrGXBDatG74yveZZ/T3qHDXxqIbn22Yo4QSuWxA
i1H1xmsC/XDT8rp6WAMD7q/WfNs1AkH2i5mLaCDjRfshy+IKhuLeuGsZKaJDFTwm
q41XnEuuBHljQODJ3D1DWDxMsYlEnH+c7AfyX0NewBh2CnLEaHAw/SIHI52Me5ok
GPPA9RsCx3bu6urJXlJ5nwTxSBCjOra1N9SBt62+b0BeOH9pnj0+o0hIlomQKJwO
RyP8uUMqwcuEOV9de0idUokRsWK/VcgFUw4Fz7oGomj2ZDywmu7WiEyyBzX4Pavc
rK6PidODg5AL+ZqXHd12KIHJ4cZmAsvlMXKV5sQzMylqZLvFyt9OYXuaBeUzAIqc
3NuQlFymoFaIH4zZmQKrIst1xJAychRR+8kGxDIC75ReKytmVrjUr+sgMbm0jOp2
r32ZGEKqfCILsEJCU7V6+MJIKbz/l+ZIw1+3kbbWAughdEY0AcW+lxfl1m+6eHbC
DMZCGR5mF5dnpbtkgSamZiX5AoYYqVklPUPwMmtNlRJz4jGMcjwk+BwctnzunDWd
/LWk1cgU87iz61757HxXZyxo/XfSxunYMkrcO1c42tsy2D0OlDXaDy0+E6VY4AtR
dqx5Ir1uQ4BioYI0xJd7TaHV989RstgrjVtukxhWVAHp1VYCtanflLlZVTq8/yYe
LfiTkh7159VFu3heYfhTx+NbQ/EaGZSICPb6fU32djBnzL/HnTUiyxNxII/ICaHe
xRtek9zPk9B/ulyrb+XTnWcfzdYBpuVZJ17yQ7mt4ldZlm7iXIfaPNU1+w/Qv/4S
HGxtfZbeS3pVG24W4fmsedmIeWh5/Eaz2zB93ZfmEet4cDv2PKBXNZdYbM9WxZsI
e4ANTqzyPRbXbnIWQIVwYXyQTBb6bYpQSzH2MjGamtKcCvhF7n8lOi5XCUprkoRZ
23p59fTcDnnlheQHPHmimMY9bXYSrmxdQqwNNaUMCIMgmVpy9Olr/WcA26wpL7e7
qqFay5gv06fqQtQX6+mVYnZWjChHIvd94j+BLIEJbr2z2HEb04Nnk+tx4agnJVRF
g1bm2kO+l6bXvi2O4vq2hx78tVMuneBocFbzZ3tUU7yjpodKDp3F5hX8h1tbJJri
hGys8Uly+Xbt34/r9HBm8S7nOpJqLbhMc/Lln07oLmueZsdRDKUoPVWd2qbOo023
fRgLlRlN+8iWJE6Zv1vdRav3xGuB8mssBlbrkQqcSx9cNUMAA7dk7RAcx4pyJR2e
00DVi9IThWqBPu8uK6BY77OLwe50tjkfRSQ53L2uJw8HJJcza4A1xcTTEcegosbh
8hHUQfTfw1M2iWH5MrdqWjqYltbk1HSv/wHR7e0ZGCMPhIEcjYD/TEXQoKhwKLNY
hUrS4UrhlLXCtiOitX1xQgHAS7wD8tKyTE2WnpRaKNgZ402itMnDwqtGIUi4Yksc
6qbJnRd0DQ4pcjlVPZBDLqlDhRAHAmnYdExzfBrahgz1RRlnb3V5yl6HOLCN9FsN
9zHOBklKi/TrsKgkIi9+MF18lCU/GuSDeRPVdhaYMeew6YBHYjhGsYPAqMoxIoA7
hCwuYBPhTMEmttlihX4mrgfzFPb85ycvWzskQ2j543E3WtASzrvJ4HpZahfal5nx
Xn5+SL1wWAOw0yyhX+b0z/6fI06waT3uv4muibMaB66P1SQPEuZAISlrxzxqvpK/
Wt8845uGa5i4pwrafNfoLttYoDBaaRP2jEMgZqKRknyS+wSvGCQ7ulm7La4VOeVn
JQ7OWx2YrhoP7p32x9wotMfK+JaRR8HnwMg1Ujna93BWOXLLJ8syXQtdXBRldacm
m3RgCahObRsxnsbwfTpvUSimOduQODgX9pEOsxs4AiRhPUQ69h0WidEsWQ9VLYbd
0dIqO6ATwYJK4IWAJLKM1NhsXO6cpVzvz0pVCswvbuelqYefm2tg+9F0MEk5zPLA
U2TG7hyiZnfd9bwo5fPquhqff86TleFNscbsWFbCfzeQqB8CzfpJZYapPAbTx0ct
ZAuYayJYwXTPT/qMkYxSBCJ7OOb6HvxRXGbAyXd+pFNzwYiU9gh8T5qL4I0uUg1o
SCoTwtK/UcagGhLcR83rVIanTcu/jupHBYM3RIFCrqqvzfoChQiLqmfG6KNP6jow
HIn0nuBsBJfXispt4MfmE79mel6WbYyY+mEuEd+1vap4vNzNuCQbgMlN2Z7t6yAK
gZLbG6r7mj7ywVgjVpljxniFPQICm1yH+hqAbMwpDsYFW72aFEJN9WfoQHBGe9yS
2eP7KaGtfu2BrA6EewEMngqoCwKyT9NXwq15wIEMSK/P+HvjInPo7DiQHHOTOK84
0N6yV2/FUqwmZcGR5HuWjVouJSnexS49lufG6kWkW2jbQi6WvD+fg1/E47rk4D0H
ZpcLw7A9655eeTjduZFtpmt4KLCq96AWQnnJEcXYo+fakhAHNaV5Ux1q8rLw+n5S
JzY3TWFQhpqD4cVQADctZXA2xX87wzZMCZmp/KW7LgWk4JzKTT/sLzDJ2Ojx1nOh
V0nUVJiUxVQ51MJ0Ngkj54iqD9jlAY5KHyI69wJSFaIRuiDSVg09HobB5v+1keEJ
tNCnDe9ynSDkdRjr2XawLzriwM5E/27BHdz1Tjt7vBu2sSQGZZrEsiexrBC7F1vm
3LbSJB7CQErZ1U/wGPN166jJjWaguET0kBZWEBiZtjam5v8/qd1VcHs6HRfYrmT0
eRvkWYC1Rjdjec0Sc+O5Ez+hEwseii/LXM7D/qQqNOYvsCRGNj0OdUd2FykG6m1j
s/WQcJa7mdcEfYgoYlOgg7Gn8HeoqiKpnfCTDYQYoiUSPxeLBY0lDO6GK6zM9L46
xtNnxnDEwz2ZVGi8HuXoP59TThcykuCnMMaGvjaEOK3OQtTzMjALp0mzlCHu/f4D
RFIaYgrpPwAM/Ldw3Vb7JE2WLZeHf884fWw6oGjvvcoSzqf0ber/CnNunk+ii/IR
LyL1YKpFdACW+3EjmXo3eCzgeC3BcPpyoXJaU8ETVjCGnKkDlkC7/GAPdVy/Rys2
F+JufafvHDQYU+lFxO3kfg2RqXlXNeCvwb+A4dENB9OaXd26xSnmvUAzlsO4nJvZ
OENcIm6K1zGaUC4ApTExRg1LQCs7EVAyV95WMmipeuORu46WhI4PoaVUgU13ILYG
eRFcmS6XxGzSDbCg89vRcYc70Eui69e38PjE8Nq0O+rIATBsb/My9S+9jYhYo/Ya
uDnvLRr/OfZ7OlX1YDyXbhumdqPmWyXFGxy7X6SLpRTCgDKybnKAXhzqlh5Nuy3L
6DWOe8TvARpCya7hxp6JFqahzc9Vy6vZwGgQ4VaM5wAKEI4GwjvZOHCpkx/hzUFR
rfK9wrUuGOIzIIJ5PQFpU9/l0TqwOpj6FoDLfrpPZeP3wLFx6uYQnN2mzVaTpO92
TfyBQVwt74S8djlxMwN6ywu/E1Ug/n5n9X6ioj137BEcpWYl2lYSBiWRyGrLo+ja
+g88jsqwrmfoV4xp4xdKj3JZ48yWebU1QeC7CCyU+5f0G5eYDefi52g/th+teEtj
e87Jz0E1bvAEhc5nhZMFumvWPmlAmdXNoncwwfZhFmNfxvCbY2H+gpXYcOD8y7Gn
aYKrPOOqTUeVfiHUuVpqi8gD8Lo82UCzCQzie82yZV+Av8O4GiemlIjHKD0tpFbp
EN/1vTIxhmYpqHjrcMi06Dty/vFeJVJbn2Z0sJVqQo1tv5RHhLlDiKfXWg5r/nNR
fhuQD3JSL9I0QGHqdmJ856MVzmypS8nnND69t3/CaANhq76Qmye8Prbmf+WLeARZ
pS38jAGfpGOLOJiKgK6la+0IziDUyfnSiC3Srp23FYyOu+qvcJCNoM9FHhlmfAHi
GGowgZ5kH6i0XOJovOg3/hyPb2PneL0cVjhdWsC1bwL3Eaqfevv3ci2Z1KRWX2Cz
uiGW9lnHEuxf4D8cHm13jMwjBq6KUlEyDRtmNqUj0wE5DJ0dQKkz1ajCnHC0gwBn
BQOa5baKebknZHOgSBToEgqXzRL92xRDgpCPs0olI5MiROSRCQUUtsXCMR0qchal
Ch/xBM7AoB9s9mAfJ1tUcElqDCJKljWgHzsxeoqH5D2cZwm/FYhMq3y/lX9K4Swu
i73+A91PyoNEdfLFPx0ITJvlScqIKf79duognPq6skYR/qWJMamXBDqNp4SxG2PK
Ge8XXLV5GBxxFkXPY4/Shc3I28XQ8T20T1p1a6uB2Zhoy9I7dr6h1ssWmOT7EWzF
T9oAm7S8hfNMmyTQKeWN5jt5D98t3Qt82YAZQ03GgZtLo7ljYYe/reYBXAjFjEyv
rOSsKf2ST8RegOyki6fMfIPMiFBkp8vHhMe40yK3xWN2wSezS99HonbVXaP5nafP
h+iKG2zNDgUSqxXeiCItKf+Ly0SR7zXdYo8caidKc4+sZPaBzxQdyrS3VzL45TeR
3oBEL5oaIuH+rmngFFwn45Us9HK9X9TkYkzyXMRCzCEuVoKj+uG6iMb0cJSMJUJT
O2QVNH3FCSYFGS3N/bSxOlWsdsBaats2afWX/CP3cIlr/Z1OX1/D/Ft4QLZxiExs
Tw6NO0jOWDoifPZX1UzxXZvRAPt3jeQYdF4aMVW570N2vDR4OZxa+5PxGZH8ze0t
+W8x+JeCJQyZDgz2ebcs7L7hZtMaPLeeuQuOPCYp14r23jNtcWyTr624aPjZ9rFa
Rv+HfgxBcAJN9lAZuW+Bp2FXzauaf5FhLEnpAJbT9jNm2jf8iO2dhOh0S8Gcuimz
WoecnVf3ncHZIRs3JS9b8i7GkR01If2bETSJLrULCqGw5ULSwlmFlhV30035tEA6
uabn8048yDfXFXDaLVS5N3SSr8R57B8cBzJsroyo5KIEKVnol2hmJTTb72ZNTmjD
hl+puET/t+Azou7t3cwswGYRszPKX6RWPSfuyh2NSiGZ28EpMFp2BWpy08CQmfY0
V6Im5YLHUTktBHGfVplkOwSlOchAqK98Qnk538HXevhtVg//9eD+h0VkblHcrjBE
PvyMxQm0k1QK3a1S4pyzP6I0EEOIi6cQ/JjSk1XSXNUgv9o/VKBP4fDfOq10YlQ0
v/yHzDvgO8P3gn1dfzrI7ETNlfdS0kdaogIvYp5b+mG8Zc743bIt07LIv4u0T0/x
V/hBhU/mo5xX1LrDNb26MYOfWge5mnRa2MB/oU2DuawIITMzPI29iiVIDVeWYjbI
jWUK6b86CFo3RGl0Hohnkn0mumT4CYz5e8Fb3+mV6x2VaDIImGOL0plg1M2X6+DW
4C0MP/oN2wFmQwP7JvGF27sOHptgl0v9EJXsWewJ9OLzsOPsSNJ1TCObKsK4MHr/
eK+qXK+qfNBZFf4MV9OrNbyU82YXYW45cg9uaZVIseTLyCvfaPAu1as3qOiC2D5P
t3vrIurLOC2LwLNlMvO/5xCuRaBsIMsak4nN9joBbz5U63KFNGacJqaAOFppU9GI
YsnzaOXVUQ1jFUbA7+LK0rndfbSFXYsJtrz/ygzIsoRe9q86l5h7UnjE3VpE3i/W
ZE2t4OtiH37lgdU4K0vNFI4uE/AvQkmbYoGN59YKnmQmj/CcxL3lxedrAbb/MW7h
XA2QCsWJhHgoTCKPsKHtUnFBmn+ipYT4VhbvBYy+0Nh2A0gFkg68yBH+JposQPrW
ZG9FQqedWByPIQcdqduOLeAqvT5wBUNB4u5uKkty6wQced24kPSBJq42uEV3VNoE
HZK+TmsXpzrNEmEC9lhPpzac1RxVl2aVT/0eEK9hNmd7QXDFbVRycL4avvVXBN67
0lQCb+81TYeGTvjgZTImBaxSysPAy7RRyNFzMKLZcW40J8PiyNRHXGtkg/rBi64P
72T5ndJX4EJUcHTniQCAVeSqUY6RxjYybLPysTDGLV9AzVBBqW9R4YH5TTLCEY4u
IJjpfnrXgGNPVzvULle8MXiuzu1PjMkiDVBqFpdOzgYbZyKSna5VV8536XWiEqKn
B8yS/zJ/bRYfegi1KoNgRJnTVYhUP/jHJ2FGmym4AMhOvURjg/avRm7vIZ04iWzX
oXDNoqwXjefnNOuFYoZ6NacBmqquIzByBWyAVLCT0edj8MZeh7sG9EgXzYkGfjva
tvhtnTpMI0+rND3vttqHZKxJthtQFd9BQ7tpXb0qCtFqSbylidEj2W2vAw66O7fb
Zdk+pZoU5god5ozBVLQ+RK2BhW+QQ/V5lwoee7+41lHZh2xdWNFmUiim+7AXaMtN
Dzgqf66SdcUgGFtIgACo22y6FPlq9edLjqyhakWjPLEB5KqESL8mxKbkvOc3n5tb
8aKwWPEcIYPtTS5YCGMAYwuNSk2P/9xnmPoF0P5FXXkg/wTesTiDsxV9iO2UW/LM
eIDvHk3M+BTop/ps0cdvQnBTqkoQnBPkbgI0Ay8cDSXU2SifMeCCT4uSH8nSu7Gm
C+BdR6YaGsLGE62iOOZGYK6bEHc3uAFvdVsZ2X+eb/ArCQ/F0HFK9UTQpZtSjnkm
gbY8Klys4qQytPiDD+AsQbZg2m/N5EgY24/D/Itj5/nwS3eOVzBDcrZQrmn7VtFi
rPArUea2hfyQN65+F9SjWyXN3LCfZrnZDkbxodu7pPXFf3fb/Fyh8gRkjFbP326H
IwIyl+ov475i+GtpXTNTRb3YEyUB9DVdCH3CTU2QAt/1o24fXMk0mqTK1vShgqLm
sVK6LyktP3YwBZqkj4BzbgSXkJw9JGQzXOOEdXWz97ZmK72tm8GfRL/hZJ/cvLEJ
ar0I1kExieeIqLiL/+FdIO1aBWxqeyEsAuuypIFAMM/tSHprdK/e+J5Fa04cABIg
qpYpzuGXYMqZN9gdAM0MGvXB0c2ouZP+gii8KDRjrg04/jDQC4ZdE6AhGEflLEFB
6ZQgglw9Vjmck4t7FeLiJW61m1ld119z7jE7fXprqqsKb1m43+IhD0o3Ee1zy3tv
VkP4dNOAK8rDwyYHfaI6q0d5g6v8sI4EAhNSAmMzkJPLYSgUxOyBks9UM4zWq5R5
Ap0kL0wtOI0Fo8DaTug8+wp2OjXGezNCssKtGrF/GsMJjmSza5Y5Bhc9QdbamUg6
/lnlih/33Vr+b6Y/aTUdoVPETFB58gFx1PfDK64Q/01Ba4iXFE4hxrKu7GT1jlBV
W7OJAI+SHYOpw2S5/hnt15/tIcA5HVaC/g9NqEMCNcsy9vkv3mRxztIbc8J5gipV
Gn8tMTBszBQDlTqgG7jugk6OEBu1wcaHWDWEi/fB+ieRfVc5OkyptHK3MvYQwy3V
oZK0ktYUJ8sBNz/FtS+2i8TWEy8i59dj0KePhBjEdfPIzuuVPPZgSwrz1OmfYBJY
oAA4K5DBiE7GIsLsBQeMUF6C76OO2ei2EBVLR5wO8xNLmo1aI6APe86kBFi7Jhdv
qoOGxlIxRiWtIm4Etr8RqxZV+CKnH6UCUTtBUtanTpIToAc7twOvpWXShCqhXHG5
QiAqTBDwXRf2P5ULLhTfgy8p7GqSWwlXWNSyQShGRh5NnFqja+hLw6Qmc6Uo0X5Z
FfLUYbiPIPenP1bIQCQ9lchW0Uz9jZfLhI8e80qOhkgt5PkmllSXYVwDWlaX96uc
SIkNF9356chMQJBhx84ANtnz+6VDCF4Rv/+T5rxkLMD+WEvw+1BMzqoheeHjxkqH
/clK9W462Tc7vWe2z6JJ8PonEqoMrjOfW6Osx9WZJvFcofs+lGkizNG6wCVjS7/A
zV921cf3KYcgvDUVIkAiLnJQu9hjw909MNdYHHjEmQu/dzGxFASd1Ehq68GYzwcB
ylUljam7DDRpT8nJ55K2LpFxPXOCxRWBQURrDOt9oMMoh0/obOFYyecNmZq7pBY5
ZbH5nCfARY3QiADNKyMXCopQF8/d5CX+JLL72fBid1sFSY6o8sul61Mxe3fx8qSS
1MnB13rmPszERpBk4DH4Pn+j+Ub86SnHrMgUNK+Z+euMW2KaQkalbQii7kWVhGQn
q2WjVyyfP1UvkVj3XWB0dwsA6uylt9g7g7mA/WOn5StY254en69gxR5MOti67gt2
649vJzjOYxAtz8nAN7TXkSPHCijyIBmAbT0g8fZCJxl0i1H0YlKIywlN9TYioRGq
p9MFPkkLU2z1QYoMrh+rFmXbnes53ymbk80WNDvPlOO3Ldw23CzxBC1WjDb/QUXI
DFk+C88SC6WbT3rGMG+AmD0laQM1eXEZ6JdOrrcGnUPgi+JekLtBENfJ7iVTvIPF
wTUWjWBbUrdB7qqADDkmMGXWr7e4ncVXUnEr8qmi2pf0mEmNCcEkZMAsYXKPZSGD
nLOap5tdAUkT8pVjN/5LHM5MrvSv2giAbcTwD7dU1D4Xfp0v5wW4oxMDMFubRbeA
nX+HfLtm9Y/5q5SqEbSrczw21RM/Ifm/k7jTg3It3kiGNIMH7hYiFp+xE2D3pCMb
2QRL3Hv9+QZ5CVqt4ot1rNhHcyE6qNVM7AotHO0cP+A4zAazoF8YOJLqkf9ZD1yR
OckYGT/cmdT5rnPQFynPFovTkqbVEVNbrEWMBXfR86CRBkYH7fbZy5WSzsbGLthP
/CbRaNuBmSUTL1fqPorUpXFYhXNYe0b0yL7AQQB1KdCbEz9NqPfBOVksNa6rGgD7
7771kSxf2lvM/ZfmWOliO9TbqsW+yCfoqvb2MXYWHTk3CIOO3k8SEM6+tCLzmnQW
IB1sIpXA5cd+kXQKmCfTrZdytfMUarTgT8aDV3HIeSFcqt5Iw9zagSjqw3pRgUwB
W6kYJzD2HEnBOfcq37hLNPBN8H5Nvj/yahLi8WiM7DvAe113Sa7c5BQAazgo6JIF
m+sueLIwfsw5km2iTWJVmztAbPS0x/jB61b6wI1JP0M359hsyesQapGmMK44RQqw
rsmSAeCNzOT2xH7fXimzM4FbbxrTZQj4TCI22MQeblWDjehE/aYuP4s4O0M0Slwp
ZPIfymjV9Mp8zwb0vx7pSeMBi5yCgBCdygzNWiYY+Z7BgdbF8LrHUfRlnMP+HySr
Bo8oaw2Y9bvZ4SuDSfPGCjJnP5NThQfISdDl6n0hyrEuhsw/YLmJ+KXHWgODuNrV
8/ACLV++weVwcfof+hYwfHuhze80KNbSlSnx2NS4jktNJASLCQ5mLmfcX5Gi5oaD
gn6NALFMrXOCkh1nJYcC8jFDUpo9K8VFMXALf4ku70L72dEOyLxrltxJTovi0Km+
nsMj3r88QGBDZRzlo4J6lQlPAcBmxmShq//r/Hf//Fz+4eKeCBINU/66eOaKWjG/
hn51Q+5Jj82ubx03T+orZA8nNv+3wwo9CLEHIKYNBUyV0bNeEXkKOPQceKtOn1VR
ccWt+Djk8EKo/afFaWzz2VGnzt/3G1GwiDNQiZYTb5Yg1kj4ZLZUZAp5O2aBgGMv
ORYhYQejNDHqfiNMs/DXT9kNynBbJtK4q1s/XUcqoot5K7jg9owN7DbeD/FJ3UCc
ZtUfnN53Si1+tZ/b5e+qxcAxr6SNm9HhZICRhfiQGXksI01XN+IWHFDa4R+jIyCr
qiuOUiO8SDArkvp4YThUf++Aji53mtbj+fOEu8nHAgs7NqWt0KQstoQa7+fKCfHS
4yAZmHxaY0EhFsDWVQxS1sP+YeKoGzhmk7qgly2+8B+2FNYdVnWm+dA8RCaAH3Qf
FdyvNa1XMKBO6LxAz1l2GWB3pCE0ih95KKNkyJOQ4A3BtjHp4QMMaJFnsHQvkR7G
kC404cjZ16bisJ/lFI0CrgI8AfaNP8nuXoOnRqZmjFLn6WAKrsFI1Kr3rBsjDUUr
GIkGufSavLY3mJ6QR6SP7iCIaXOoUgz5wq3pK9/9td3ceBWPD9cy3mneRhW+te6E
Kn6tfP8fqiGJb7RiTdaXJKjpLRjN6jNtYnRZ3na0dF6iL2xJp9k2cwxeF0R2bN6X
FtQedb2haV6g/hVdkkD6AbGl5DvfGjf1kkRucX/L+P8N0EstGlSG0RW5kfpi1O9l
ngocKvtV4hMBEusfhcBCHT7r13GVZDflDt4Li7vvTINvhvlzBd70eZHHsYoeygLH
bOCM6IDVhc3mW7r0c+GGlDn8xfbHPc5C1w/MVoJGxVquDW5fqqQ8So6+111bXRa0
fJfKIGPhGScL8sVvQp7TXuMbkZ7auF4ptW2C3ywzQgrmSBY8SwUUyMxkF99zGEBh
WbWHenbRlEVF3X4yD8CanMO7tiTLKKDeSzxJMorUerS8IHHcRvWuvIoGkxeYWLUU
0y1p/pod0NCPKZUQ2ucHWpiq0gbeA+10zrZU2sdCjjbtiAvChoTNndTuhkWXRkZ+
dbVZYmYtwytxoNSIlR+i7N43aQ+JOAskTBG+iETUvOR8Hi2r/ovX/C6AESyk/D5v
Us8nrT/Why8YGv7xFR/9PE8I4odtiEeyC1TlaNJhTnljpoBK/J4k6Vg6X/6L0aBg
pmRz0OL89ySg9Cf5USWGjl/kGLW6xrtLCjfhPsK5UYOFm7Y5TRrz5BV1zBxqAuc6
iYk7YrxEXq3Elp+SoXAu1ASq//kxrNrhN44e6gB2svsrhYNacGLUNozB+HDiv6Vk
+OT1UKZpwTRCqkpXGOtVC6pwt8U9e3pJeZ3GWM0yd4Re45XYrxxa7Vmh8H+7ustm
0I8C7xV8U5ooY0uOZ0wxcd7o3XmgpGnqdA+joulwzHc70dNrx8wyNPGDq/L/Eqvj
fqso1u8/1tfnAS37+SFeY7wJ1Ppx7cw4ZQmj11PoDDs76kWAMPeNLL+GvQVbPQRS
5CUimzvFgIDvl/HOj2Oi4fSUGHN895kzsfMddKg8zYMFkXnh52AwouI7/UF+cI/X
xBoSE+/dyRwOwhU+NupdXyQxJQBi4/t2SMHAosJOSfNZ2O4K6+Eswg39R2NuuAj1
xChAvxZZmKb6BsOs3tGqbkSormAKk+F69vP1zM1kV1N5tljVXv4B6uFJdB7OumQf
gaMQZkLhEB8E7u70nstHN4u/pTxbVvK587aajhJXsZb8KaKn9EXls5ryWtM3qbNe
pzT5hvKlwnWZIgZuDBP5TiYILw/q2ByaDPKMTjujHCioOXwxOr2A42qm/jrjFJej
bmQcLN3G/nDLJm0N8nYzmLNkbEAuFjF0Pms6+h6lEV9qEkA6QDI0q87i5jke9ErU
RTHJbdpZj4FNizbj0Ew3xXXYna8FYxjlroHK+Q/9pRge3we5hxnwJDr6tHhbsFAQ
2/kt6Sd1J4BHYm7jbIG5xGpSww3kyH5jPPqhk5Qmf+8UYzFlPrJ5lS57OgZ2f6F9
fW7pONGLJd9blQeh9KbkzOSuTWuquIQ+zKHonVVNcNU7/I1bfNNm1lUtm1KodN+K
uW64YHJ3RH3ULpPhJzz1syCrwmXZV/P2YGW1cCP4L1nKj4Ldjv2LlBYhPdLz9ers
peRGb2C9tX2LcQAk/r6UEcUtYc0KX22GmBD5Nnx+oG9ldwekDU4Bd9VoHT1htPh7
qRFxPExkoLbGaAa50V4yCsx6E+/09dJX67WfhQ8xmX55rryo36r6ySBXHT9jD5vp
UYR8+MEqyeoDKZPJvZ+3jgO3FZ9LPKBMYewoWpynDSKJmCGTfVrHkbU0hLFhnVqD
HxSRX2lUGT/mrWO6XQIUFZvYOvDN/JKiDSftmMszcQDig+KK1RfeuaKfesZ4ue39
taAtB9v+4IZhiaUocpEoWcve29fUZJ0BFi0WgzdA4IuVbPEp+qee+8qjxcgrw2++
wL1VisOvqAGzho/1RVgEnlRTDulNKjp/efn0unnopwm27EpbCjADaWEuiNPrGAaT
44PVcXsPHt5cUQtvNw+I1WO9Splnn1fid50o/rwjhaKxlsB3qslxl/LNea1slCSN
2fncMmymyLWsIt+gnCLVbMIOqPhnqjVq0EybU8jDnoRtdF7QU6ppfV0Awt+hZXFo
eWgktFjZiuiVg0JGQ88dNuehLzr6b4EHO6jrcIVq0WFdXJps6ciLKjYkjN7ee41p
QoGiVK74G/eIpumsi+kWewiFD/Cus4rc5WnFm9C6fPrVjhrBYp4W83P6yZqSWCZ0
H965B4jWj/fL8qg7b10MRP5t8URubFBShrDltEhYmsKyWNoZFRS0Xif83lXokc+A
Co7mK8ZNiP1kk9cntw5W/Cnld7PKACHeLPoxdhGn3PzJscjrkOHSFNTq/sB9XAly
DfmZGTa39yX2omdXuZLG5ORW1eDRjnHxtj4yoJlvPXJ4UWPJmfE+b8CHiXoAPZBl
AnW+C/GEQVNPwANz4QJeqQNnWOsGbl6GrMCV9tM/nDgA1LqqfTksqHE4lpJl/3cu
rYk741KArh5dXZcXyjGt6JU5tK90+GWXFPq6aqMeuMQbL6yHlvk/lgVFK3iDG8Zr
xKzsru8L9VktPTL+gNUIdv18L+6G62u2DmKW3fGSmnu6+8ejUpWM82NJk7Wj+3jZ
I3ZCy73vKsjO3mFH0+moBzaHYFBdwbp/ysu1wW4bdWq3ViC4W9XmWD+H/v9UFIPb
ukzEQB5rKz2RA9Q3jTGg2Vf90fJJMGFNew9UaVyEOUlQBJ45T1xRVPbjaK79ohR4
h0kDtsjWJY9glajynX/i/PgFzZAHzOnq+PKyQkujmrmPHA0NQgrdOgYIqH2yGOId
WQKrVsImL0bJ/BQCKmhv5L9uaX+et64uZ7WI8NOIyM/TcvHD+Zma1kmrT0o7OpJP
Aq5gSl8szhMftyRbxZoLY9ZAxjrhqVtBJ0yGkq9RijC317QE5DKrQ7ehBCTBdhRz
UWeAW2AIuMSnzvR4E4O7QIjUgSMXhBM7OPhUZ/MrBVRClE/fOcY6SPqcPjaaoKTj
5P29G+tQ1dmgYqqjnBvNTnNsjtDotdaqk5g1LNfWJy4MarSFnnMwE0QFzMgaZsZF
qK/ZOs73dJ1p4OQiFmqg9x02tsZ6pbqMyNGOR3L5SMEgUVschmE3glQUFObdG1q4
1BifeU6e5x57boswOtAF85b3n+/DLuR+aP5BC5YYioGuT+M/u4uZYgFR8pzn7khh
Pv5jwcGp9Ip+60sNz1iL+EJ7O+U5xl7/17jETCcDDiEDdc9nAypvAWvEsabQAUHG
ut1q5otExtYIsYL7YTaSfUD6r0EvHvvPFrdj/yUvdL1NfySo7ULemenRk2kmCgKl
6jG9JDEmIYN1YPBBDZlKOd962/fhvFBThVGhl3QsUKym7znRRBxWp/vsR+K4PL1d
dy3SZ80dmRcjSGb/RpSfLtRQSCtW7r95zjyDHFIn1A+OMNQfOXiJ7WtdtrK+orL0
r5S7S6/899xheHk4hcESxmR9pPIt9z5mEwJcz/I03fLz0pblY7aCmM8WmcTPDZho
WrDwCsFdI8TLkXU3eEGv39cnpugTDenpJg3IdPMBnBqj4jkmzIuo6934zb5Gz2O2
IUPbQej7KLjQmXtougEiSpkVSQxt+XzKE8iUDPCk8JsJKKRM71/TWAm0fcoDgcJp
ajlGrkAkuAbIoxt46MKxuLvLPrghYXQzJWPR84d3oWKO8eorB9J7OAnskKWjjV2j
k4FT4UrbyYKU0HEc5qN9bAK64O/olqq5ywaZHk2F/02/XFj+RvBl3DEwSOKgynsp
bxmCXK99LWLP3gdnHVJkPu06pofIN1TaThFnzC/DIXyO1vPcDlkXSbOwAnc+nnRu
hOT2hYvFpkrHuR6WqFgKLgAuYoEiL+36o+gqw3lerqZEOg1De5Mzuhiof8FBTGDB
Bm5pkHzc1ES8x28W1o4MyCTG0+qPUgyp6l88F3TiDSIOjkASk+Xlei4yMu5QMTLi
NSZCfuww+p78t2VRNztyPPxYatY5PWvMAq3kn0OBKeokMEpEC2NVvucFPp3+kgHH
gP263EDnzXLH9nqQWzMbIM7+8yp9S8inIQtlbkYAqFpui5u9OSfnPesg2sOwPYAG
dEhX92aXEg+yWCwyPIbiHWteg/QXxPLWEex8Py4FoQpgKQht/WhuEfI1Ax/XYCnf
gKMewQW59VSBSjhVmzqlWIhw3cHc1UoGrRkIGcnqcH8lPpKwXHDIqHRHAAwzZnbn
2/n7XhILWnRlWugqs5ZvP5/nq9Ib8T9cgLQdz2/K07Spe9/mnykkNfkDERTzLWDq
T6Bte4NDJIyF2rtzaW8u7p5XqV/YpdYxZrvrkKOmNkZlbGuTvHQ17trVvYng9nff
6h7zPdQ2GA8UghivfbomnZ3uKK/32ES9djgvuJvIp8wFOCOVPKL2pz4rvq4ugaba
WxsgZKgCkjsoH5WE1CtKQOPcYyxU/lrTbaEewneWWtgmeRZFB3ZaMaVW9EZzaJ25
RRUlq7JvKD9ek66kNPiND7ysMcxuYizQLfgovBRBMXXbDziTkmv3zyqKdTbdHUr+
wkoNXY1SD5sZd63ej7qHZaq8OXNdqKGAYx/VQBbGinXQS9cgCWhYrnGADQubWmPz
jGdAfSjw2lPmhoUkeFNyDwIicXOPRkq4t3b84X5CPzH0sGA+NyO5FI+bFKr/RA4C
4XtCm90zxgiDp95uXbXdayRoE8z6e/Gs7Bp59VCEgL6Fwdn12F1ZzXmMLTkD/+T/
mrf+lPcQqCX7Fbc2jVkCHprFUkbOgCHpd1U2b13QXgQldBZHahs71Q7Bj463lF3T
XqXWkWAlUdIF+8d3YVJwSTDDug+fblGBy73krclbr7RakV4lnOsWZHUP1aNw7j+S
CdJRiPgL9vaAKSRrs6h3QLepKGs6ViQucIsIxlf733SASLgo9CYBMo0rPEdOV7m+
/lxTHdHk6JKKuCn+KVprDZx0B1Fla7RrqUlhfGgtehY9JZsmT5mZog1l1lTeDTDi
LtRXsPpuubJies88/EXWmQTiMKsoDZ/etX1vmtb8D8crxnDesurHHcAuQe1bzp/Q
VGPNd5YO/NWjFCL/zq8fqwGT09ODV1HO+nJ8+LLtI1zXYn4pOtlWFSLNUc9lY7cv
KZelyVWQUFsz3o//xcVGA7qQkgXf3FDDJeLzYJAkgvWAbNVvzMaUJHbN2TyMkkub
dZCztap9kzqt5BsFzixiG6K9VBYJFYI0fT5Wg3L0GQSHWYZ+gIBT8uO9OZGpjHRl
Z7ra1ZQ9qlM0wL4hEDnWO2DemdDFoXkhHAUmRfofol3qZikRqpQthC7wuhgwNyfb
Ere3EAHsFY1It45k8sJ/aXVmcJMkf2cvY8S3PUnFvbSrGxc1RG2vhmgc+PjGcXHf
4Ec4QNcU7TEW6UNBIMRSWnhgAfVEqsqoO7HuwiApHRmqXhy5ATm+/r2lWXCRAVZo
tYftMCOnQLv6/wJqVMLuL/YlClLkOZjDy/EzlE0zGiCgqOTWdSRomGmQGr8RqiBM
MyiXhN3ZMa19IgNWmo9sac0rbe6G28TQyWgYow574wYw9hThE4OJYQEsYmcWwSBZ
ogoBWa0id5Zuu2qJyspqv76safv+6VEDLA0rAvVIVGNR4poaFnwbL8ZkXUDYHUSN
zIJ4okYypTCExZmL/g58+uguMenefViHUgWZ7A8hZAKsHQEqNLI5xbDwqP/cE3Qq
qUfFoKL18mtcABQwsPddRr+GtyY9tIW3MdEZT14/BcvdtrGZlTuMW2rhWYjlDoRa
xCyg8RYdcX82i1Ae9jurpQirw4v2v+bHV2W5dH1LLeu7DnG0blwGMmY0u+10Mm58
IpY5sDN2ndjSJa6669ms2ogln8Fqp/juu28xO4GRvVaI47m238lQSmXw6320boFc
u0dv7Zb6dgKPgDpF0M0m/LaV3fiqG++3CRS2u7KBYBsg/aM9j8zwnJ2Xp4mQXF3H
2kAcVLCxKtU9x9m8gOdm/S6xFvyHTgOHBA5XdMrUYFzqv9033BUMxCW2NprFhpGZ
FdzKVFWe5B6zYQtsOio2jl5182LOUUJ152fJyCtbC3kzGgyMux3bUxnl+34ilcje
CXZzoAZz1RiKHK8eTwta0w3IrwUM067XX1RJKI6IXE5ZU77FtamR7LjvU7AkWmkb
Sj5WPSklnVtJFi3labf7w7P2LM+14UheBp8SC5FMmPhCm8pNsiUcKt8oHYYv/ESl
7TRcZ+4DSYQVSkyddtAmlItYPkfXqFEfhTANaqgCyz9FbdeYiDdEJz/KOOrKaZ8g
qM+8u+9lVVX1jCkjApi9JXHJXEyW96uovvmLm5GStNDhwU5F1tgtuWY626we9Xj8
afENMONvU0fDUOXhxxQs11eK3ByzvRPv2t8shK9+JG2desF5eh0t6gfjC+PoxmtI
EvzcSrtxi1LgJXNCKDXwtYSWfXgly+O/Yv6PQgmrw+LrsBKXDus6RQSY7uTq6a5a
9BOAzeiWg9JI4q4cVHAcvFMy29m3R+HRewQ8Z1p9p9jK4e1WGHEaPO/CP5nJf7Lj
E4iuVGL3KPbZDLav4tU/c4loTSk0gv4jA+vznCNIlByLHTB9wCouJzcHHjpXTkk8
85VV6gchjlOOwwnOzhCj9CYa3vyE0Ro8rAZLTOvRmGJhQ4ETQo9HF2LVlT8lRfE9
HOIT3k0it9BEIKYaPwWmvv7r5mJfawZ+s5guEZGfqbOqKh7pwwe8+46mr0d9B9hJ
z3G64EIVd9WC3JDHc6TBx/7hOGETLGunt2PyXo83ZbL8Nc/+ZTb8JxffQX7PHXuB
GbCPirAPa5Lj2RA1QSbNXcpAeRUCtIFcr1MFnnmDBurN45gZzG22TK1wRfBkGlGC
AvTF9fqyIGyfPkIhf0WVutMugu3U1A1cOsVJehn2Dw6QnqfLlIrr3OV9Svmr+DXP
jOntrXkjLSSQs2V+U8HDfxdlFveKX9tFo1jP+6F3dtjJI0O+nNLXkgvDac5O7IY/
1TkK/ex7baYKmAUX0Ux5tIev5aVHbn3XznSE/j/E3fxehpJRTlSHHN0CSP4xQPvw
bcbhFYTarh6ESNGmAoSm6xUZOluWEc+jRvR08tBKzMbwGrIBlGesB95EJl+PVuGW
AP9E2039yPYrhuXpw1gxNtxGTZf+8BRRHEIlqm3tQiGPM9diSD14w+XMOAIFmWKu
Tu9kAaMOh+hrnEh0+k+85UiRYAANZQA3/6wo1cTXkz+8NAjaFN+D8M1nTmC+C0Pj
vi7HhXvFBi2s4AU5ksbZB3FzpaqLo7XvRr9QQVMZd417mFpik/xG3Wc5JUSwYrYN
kOat+k8Gf9ydbkzMEsR+4U/KziyARnav/Vc64NfSiSRfC10gguwfl8gX5gALxpXH
eNAm7iAd/PJsetVK/GH7TWf5DEp+4ayLeM9CoU21NNJFs4bWyP/F0vudOA87tFvi
WkF4IZBULaPUjaUHZF+Q4ZJu7ZvCgHcQd/HeB96w1l+xG5x7UjmQaPJLMElS5841
B4qAYzEZw/Jsfcx5f1JhlM6qORseFVs66qPUez/7kZ9EsN1V79yLbjkN8UpfV1re
ZrAWyqMDcOZezkOVn6/IkIDCDxl1L13rGhpFbhnZNoWltodra0TdL7p/HDH0AdXe
b9V1nsSL7eRNlkcFdyQ7RBM2lQcXoaAO6AWp0JvznZcckIHH7NmE7ggBYHJAvgZx
T5Z3HIasKTrit1fDGdFwrVbxrXjsrp7jQYXcLK7AwlcokuIQJ8oZ0L67/7Y90dYH
bqBzJYm2bUk24EE/CsOT+esRMDtporkuC1aC7WZ6sq4sSwOBfkxIrCync38NvJtQ
fiz2ItFy6jSRGIDAz+qObIxiRysfAqS7mBnSqM5CvvYW35aBnRs/W1ERv2e+FSAH
2B5P2EqANZhS4ge4OzJF6tIXaMc5dY29jGsEzDVhLn3aZFRxcZ/d2cj7n6yc5CmQ
X5CWKqTVBg9XJi0CqC9VVTJCliynJz0KG0UvICwPHeFeZxpcPUdpRevdHYrP8Asa
7RMAOPIC8Uv5hr6Hj9JLfxHZwCpXyCycasL4Ae9Z45LyjkBte+W9YcdNtuF5F/1X
yf76Q6Po8odHJ8UYFM1GpKi+QJ3PR1DoiqD8FVxvLNweYBFRdsbo6sEKX6+rhMen
4+LhmgJVzSCX92WvfHFCA657DwBwN+i9aLW38lPj6CvY5a8Rv3U6IxCXNQ2Ooi/S
pORFYLuyxsZi5gD2L4VU3TLpGSdoFmuNhm8xmU+4dHW1GVnBSSLllDdYgm8ev40q
1VV3UhHKx/g3GRiqr/eMQCYJYBQP6ewtkTBSncQI9aCVfqElSEgl66KdCQV94Tbj
2Lo7UykQqOZLBQVmpn5VgH54JrtJCCEeneBzyXuhn7xPHoEbJtTWBFqhdrOIlHHe
a8fY24OR2aWc5uX0zAJT8OaEIqUGwD2p+PBrVKJQ2Oe96+SdN0t6E3igEesSlw5I
4j50fVVW+tsBixjmQWDcneNHpBUnEfKyQ7NRLDUMchv1hLiPXRj7dU6NxsvGsCG9
67ik2SeOESwbPlsJaoWDpCygCdamXkAOxo69AMgFYaw80fWjhCDS9JTHMaGuoZXM
iqKXUUxeTaj0YHKcuqqOgyNHm+TE+S5u9h1t3tie1+cYpXZtO9CT2Q8fONLU3Ft8
Gtq+FU83pO9MOVp/FNRyJkoNdKjGA1nPgofMWAm6d/lX6Aa+qgnFOnKwVE6FA9rZ
qCbtvO5Sg0ym+CaHvAOiB2c/gtxgA6YeXSoURYT8OP4INzlei1gg1tKjkHJHAYiZ
Usl/LnXk5ujJaMixOBaOnrcl6ptE/E24f5DW2HXKBURLdQ16D4AmkTjh9Ktf9g1p
Ou6C+4NV3TSvJNVtjyqrFtWoJoOHkhzjOOjij6Ip+YmXra1yD5U9BryxMpu/RXYS
yJYEOYouvpIt8Y2Z+rSlRQSGy7vFIuV6u9zVzyH/7vhDqcnxgjHtnwblB1nn5jnl
O29k8zsGyETnb8Gcbj8rvZDUYtPywQLuWkwy1897uqWXL6UrhkHm3OV7HGNpAypM
4gJ7JElrLVIrNXTUlfjigVwwoBogxFQSj0DjR/M/nNKjISdfXW/Hz5+nCKa+9rEe
0hXOTaa1LuCCD1IS3xxmBJSFf/YSgCA/Jinvk8O7Cd0/rYExXk4IMf96PBhUjVyX
0+5drYj1J5uzIWk1qmPKNIH40ZIu46eZpTHVCkxbD4aJ29kBNCH0DSdGV97PMFMG
+uBavgZx6cSoEXX6S3RPXl0MsanbsW30kjrGUpFRqooz3M2fBB1cQOQS8UwuPv33
vAzzzuTSR4uKMaG36tYB0OdcjA8Nk3qUKa543HUo1vpFW6F+trEq+HWFS/wyJ7lq
YGmMCRJFTjMhgGrog2dLvsne9HeWsdFGNQhtL2fw75E5zXqEjGoI9kr+aMLjm6wL
T9ElWYiEmKdn+jY3cgXQpo5LmVlwyCFYVPOY5QBGtcwsooJ814X3XSLxsFZHEyXA
Ofn4WOAUYlmvSrcSmuQLyjqWLsqv68sinoXqDeZCZuHvt5UVTR/a6+tu4bzR4i9D
Ekl+Fvm9d5HDcZPqing/JxOaAdrfj/asD//qlG9rpDhvCeGYNOd3gSEqrCFhowD6
PoxaIBOm+KXl74fN9NW3vtLXywgYLKpQhKBLugUzN1i9eOtnxu2y9X9nM+YvAq4I
f4Z5xLfONampvv4VqB5trH+bDuBRfOJO5xQspcuNGlILtGjE3PdGlg/cdWp7I8iY
IDbO4rTA3cbWnzm94RNLL4t3OnfJ4mCBwXZnOl/o3F6rx/9244n3N9y0bIXpHO6Z
HENrIjq2cM4uFdJtS35qd1eC0x2eaeKC36MdBsQw94y4TCkWmAXIYXezMJD3aW+R
Xvr42oKVke5j8pw2FS1Pvf2vyZL46jMoFqCCBV+7pSpl1XhvEfa7WoSt6ZTc765B
INH2fa/87teL7zZHQukHrCfEm3OgXZQwQ5eG5lPuGNOtRYkNz7gojnKik/z/rW0W
NNgNy+IIJCB7WhCs+etewgTcX0XptXIqxCTAtMjNtdxqKEU8Y9/30GKAKhqEvchX
1k9oeeYjiLtTVUNN02kas6Yb3wUCCdu3P/O5BAlNb23OEMi2fMwsJt7/sSDpPKxy
ztz/kVuFCBDVGCBxzH8VZs0jOLTXLxVNcc2HIoMyL1XjnMQv6fjITqj44JxBoe7S
ujMR+LZCidxApwjXxQR/IGngXoEE79zzZxPn5jzQiIdlZVYpYA7bT61vGMK8DFHX
taSRLTUxmTEgEgnqm8HBhD8+Sj0y5hj2duC96s3iWSHa4CGG0F+3i85OWkuCMZSN
d/tUbH7nlGYKsiezsbfII79qjkQkR9Y4OMe1daG37VptfhmdJrDBd39OyrLdQHhU
vsB7Tk4wne/6G7Hj1SkeyaVSCWiXQAdrvwePSopDuSMkwfUCnansTuHIedgFMI8W
NPBXJiyHygS0mKUCKy9sZHaon4slAER+e6vcNLwZzJoHVYwiaA/m5dMCkCmFn18F
Wd717obxYalRbUEO/RvcXY3PQX1vKnRkHns79sC9qhvJ+HlQcybEPkfVGVZJGNNa
znvKMgJTVvg9cJf34FfRL/KeB8TFvwkkU2kZ/kd86rg48EyNbAtzQKFNol8Pzhft
C9GEN8H2wWDytYy48XffIIsfK4PTDgqHZwrkCYD9h0+tdH/CnW4L80M1GGGIKi2v
Ug+RLbwxNH1Yohd25AU2ZPs7fHRgIbq9lqHEYtZnAY+/+XJsnjw0elAY3JwYE7wt
tPGmS8oVZJRYxAz/oXy4PUEu8+NlQ51VhKldAEkJUQ1192vuhdVvQ92MkGq6PMfN
MKh9bKkddYPCC7jyDms7Nwd3svvEdP0V8CsjnY9QoJhtV5y8+ci3vrRe4ZODQjOT
wp9vJ5KQlee36mVLkuxFNy95y4Gse/rt1nCmKLLG6d6mw5glXQ/CFnKs9Ag7zZTA
rEr6q35cTy0iEkINKuwIVCLxzIGNErQGlrCd7wQfSx51s9sZIPN5qWsGq1irzTxf
0c9NH/J6vlpQLAyrN8gT6qDtiaYFNMc/YvSYvFnIzuUllcCP1IjmZruAddD9jjHV
QJKEXP90SMi3Cm0xzOn5z1XMBawfsRxYZtgWGOSDkzRUWSDxLCVLGKmd8ZtvU3es
Q+7ISvUd2CSgWpUgDA674ahzLJ8gY+hYNGZGDFxuYgZFhfJEPFTZ3cPTQOx9hCh9
/W0VvTgc3R2GEvwKB1uI5nyZKH809o9DwzkSNKVftm9d5nQHG8rdSTjMt9ooytfy
30lgPaEiB/jSGpmdO/Ni0Z9ivYcA6QDJphe1OH6VPZukbxpKpkIlIxBKmE/z08Dt
9Zafvg7PuTB7lxO2iQAtTKH3WU8OPBi8y1WDFwfr7q9Ejxk0DfXLgp/TNG8FuYwr
vlcxo7AdxvHT4uPF7DLGpfkIpMlwsSaj5K8dEznHR+1LYQZ/dL/VZcGIW5BpZAh4
EjrVn9rYNKSuQgzyouR2ISc/Z7u0krUW1sN0eKSU+WuuBMSDggkf6z4pZ9kNqVv3
Mm4nIltb0Cvu73p2zYFqNwWwzXMBVZAOXIMlgRfWAIgftqeQxnIMcdBciRN/gkFC
lJKK1oc07/4V+nNysc3F44RmTT17A8IhJzCSmraGDyRynQq+7OTcE5Vm23Sot2gY
ejssH0ZfBzeBq/iN9ABQ/uO+Sn5rOjgnbftcWzAZfwj8N7V92qzSLwwci2OZuoFX
qpO927w1iy7h3TLs02wKvmi76WiGELREW7wjNJJjqcwd+QJdjRqjS6EECVCS2Miv
we69r1ceRdFiQUmJBcrxnNLmMm+djb+l+Z5mzWrFvKymB5WjHLgrgAoryxFO5Wdl
KcJ0b0yYedhlDAZ39K1+//pnhRT+KT6P6PjalhK60dtwrdk/aHUjJB8xy2ZmDXLA
VGwAenQjC8sZshfjkSpw22H6zDo06Di22TpA5o13/g0b7ZVtlohGN3wqAfxBwbHg
QJxap33z/SPQ5WFlFo7K2HbNETQv0PlQYOGaxsF/IBBmN3gPphWG6I/Behkz/CAW
mCXH7HAB6MHbPZLID2PpsNyv8/GU6dKCbhKoSeoIJop+0JwiDnWQDjbqbdzGYJG8
BxjNmb+LdPm99kXtz/d89clJZch+Eohy+mQkCceDHKdsKZZ2oEvay7a4QkgaINFv
+z8imruP/3GLQFWOCBVKVWIVP5zcaoVRPME/X7btt1IVpp8DQqQON/hyy0JWA+/F
YWLkE62c2I4Frx9o8dJ63cCza1Q7oOgm6BwIEsipZXE6RizRX5K3U9A20n21ms3k
/qN1DzvxerobCdqRF62SN3NFSimMOk4HlRAM6WiljzwkzxtFEXdRhFwBv78OE/j6
rltePYV/Rq5gcc1hCmGu4y5ETuJJav/4f1W7YUMBmhWj2I11nt0zBPFdbJSq87pV
zsCGJCn7TuL1gZ4PLYF5rUoctT5tc8CU/FZ2ZTYrI8W8c8C3hGDkK3XRlKZK+1Ij
wHPMSWyFxWOe8kMeGYgz6dTvTJiIzl+SvS237k4IBVQV215lQ6mDP2idkxo5gTKT
V4XZclrCwDrutnITGVJs5EMcXrziyWyilnKN7Z6XOlIUQarJxD1e0u+tEpXwuT/B
XhRHgf6DZwzT4M88Pamj2x5+pYxfU4kApJci3M/GHzW6rUnfKankiJRAb0L9JP9m
+rCLGelUoejSe2GfDdKJwTE+pcKYcMdY1/iPOPRZ2+eRkE711Y9YpgkMQzn7vAqy
+eNFZl51k1IDUZvKZhYkBHkXdTCM0hofButOShfKEZJaz2Yj2rwJ1ikCM++Pr5xc
WaFAKYBgptkXRDs7axN1h9B4b65cwgpej8OCkVLdYsqwJUD2yJazVLfhYZQJ0SzQ
6k/rb8DwHAvIOw1F4qRyY8r0c8oJPtGM7c8+7MdG4b67q9/mu9ZDmPyChBsNaJCZ
tRzfQkH6cvvGZacd8bJ0zSEDn1WJ3DHKmlfLznq/3Ry7s558QheP2IXBJBf6CvAV
zQL72CFnnlOsCrj6xoNTrSr4Fe0PUKU8JxaTPb5wOe07GRn7aL0Lvv8CPOoN6Cr5
H7fb9aNttggpRatTW8vJhD7qqlDRVUnugY9jeo+shXpdq2EVLEAeNfwHrcHKh+yb
K6+kvby2ivnZ9t/a/cPlO+Uat39YIVKL9uXhgjj7/rwBhCdOzT43SUOcTcZ18kJS
7yDYFWV3vhPLA+xzy2T2TgVjn3U0DjeJN+bRp42KBVMm3cCyf76ai9l4U2cwkak8
n/T9aiONuzLtQZh7lzv8LzacrRCI6jn/45Qc4qZdnUjPBPocBeOmXsrMMKUzBSOA
3abv+i18ua12MeoZEae2ew1TekxofglANdAa1d5nfA2drhUnYaUmWEpXRg9dIX+1
4rlnmk+VR84napxMvRF92mssfhYkN3IaCQ4OHnokcpvuXkcJAjlO8WlNfghv/8Gp
MFdhoEWeciXtu62KRBxr/i2VcryFIZ44UrcxoxQ9SWif2yPK0TmOiQG+2wgKolDr
TTO1zi0DHFSNSLl/ZUEClHe6k0lr+4GQ9JcTlmJJLVjfkNDcvWnfxq4htD1phQur
CAmMQl/VSARK2qjGTZLqD2GNJ8Biu4To1/nKkEYsqjy35lpVTMKnzpq4hZckBsMk
FuCVOyotCJXZ6N1J/4yH5ZWD+Ft9twDMSH+M0rgMg8DbTXHN2fYK0rQVbpdwHsn8
46yWUUhNu7XUUIbF03drvhGTUr0xqS47MVedJpAgLcf7ca4teDqqw7Z+oKa0FBVG
Ov18BxOXKRx/uxJmPGfE9KEpkHYEHlYnFZHNFl6ZWia2U09llN6W2UaHpdTo0pre
P9nLMLey1iBLI0i095kaSwVpuevzWGA1nC2/JH3l9XHmRwoe+BACNu5p8rL3bMIt
qpbk1SOQNJZQZgeCpH2aTW2i6w3mYrHzlZmi5wzg87eteNAXqATS4NRMSGbrLlpW
t6Dz0nfkjjTckSfJfW6xKd8y4pOhTlPR2zGuYD82RdAY2zt15iCoTZdwpNeNOYHo
+REkPf3iqUD5MePN0ijcXxNxMOdF5rHrGbGqXjDAe/pt23aaXoGzuvJeLHJoSFjp
J4S6vY8N5BtJ298tmVcYz78deP9oLtlNX/UFC7J9w+Xuljy+UJuyqaJSlk/iMZ3F
Y1yzHOd7D295yDsMr2g0eIuODqohu9Q/vSVv2qit9XWstUR0srhC5cbDILFt99pd
egltUInaQzgIhamDNIZLd2T0ltCqay04iVGHbjUJXVkRa7jJ+2zj7hJqLJd6zN0Z
ZFcBCHgtWOuhGudCKL/Oh+Ik8PccR1GOXGKT6IVA2ESDtMnB0FukGk7X+ueiu1D4
Wobw8WGDeQRI51gqwXx/ZvU6XOtoWyW5fUsGH7L0hDnUFy8U5GIgAgHu8NvKfUqa
tkQsuorwRj0ZRqKpog+kemrqehhJk5TigBfQN7LTwUU0inFoPfmns2xrheO4s0CM
GhUGKQbjKYyW+hoKGwCwv2lR6c/GK8kA2DVQlqVpawYlk96LVydPhEnalhGrAqkz
fhRCAqfEVQUvimTKbpCkNEDlXQWwUPFzhZtDPEqTFSIr1LsPOb+56q6IMe/27w7V
pYSF3FTcKztNpobkRzw0HtgaXDB8l2gs77f+lBTxyq/Y+cDOX9ilp3uWwss2KsMy
h+nWuzXGHpJEiL2MVbBWEAKDslWOshvuY6zXTcXhy2i6ylZMba17Wq3ZPlgFcMq1
tqW3zeGmVmNXnlxRcDe0G5PM5/XRlyCO7OzTogzoD4viwuWahLOfp3qKs7YQKY/v
1oPT3hQ8aZ3HML4SBWV+ZlIxTT4/wEQUPJx+K6W9BB7wrlZ44h4aGQ2t941EYIqy
H3QQ3JJ/u68Gcy3xLii4vR+mPu671c43lPksdPXtOi/k6Tsjc56oY7KHQTwvZr/5
KdmlDQpzX3GSwWxKieWsjSMiWjPBhqBZeCA65d5p+HC4pnhLfoWASru06sQITpkM
anQwyszN38f1xoheFKosJj2mMBZv1LVE0bvhbnu4yRNBp0LxkEFugXoU6F0HCSUx
ZGEb4hBfc1etv6YKu1Fd/zMtKy/hQivQVJ2DScHZcPjn1t/6FLXIyRuFpm5ju8/0
QK9YBFz8hoSiwDLFNi+OnTVgJJVbGfeITVyNRmdVhGWgLOVxruA9sS2lAw6QZxwP
ySUwW4liMNA7dJdt6uFdhNnlQlQFMawdC6n88m6yWGnRHzI9wvH/WzADJTHw94Px
9ghxWAsZ3gv/yzzSR8p8ByZcs/WB4V2rMwSgQffsnljFrHGjKXjGkADZHQdiKKZI
9Cu+mbOXq3aEpj7DSvGle5PY5MKjkMmlxCVz9iAF6KM9GOqywKnHvbXD0OfZO9Gg
SiQUvnA4Vy1+oHwzLBFuK+Dy9aRPeISTzoONUvGrh2NrMK0UTuv5IMLjURe0SdSG
6Y1Y9SpFN9KwilDo2k4icRzks/LD6Ak+DgtE+3lmj8UdIamNxpvAnGji13CrFt9T
duY+PN3Eqkl0gZf4smwt22bs/u7RHTVeV5MQuxKvpTU1Btx2CqpQO53dCkJYrRZo
i6LSwqi56vDT/t/na5/t/tkj2h4EljMQglO90nDmBP8nnIQKJjtH7eaJPqUZIcsi
q1NJVjyZD4yKD4sG+8Pnz/Y/pma/7uk4+0a3o88W30B09kklqu8WXZ/cz4V5I2fW
8agAqME4ArcV3Vi3IQnBqVo1Haion0myrFZBgv2h0JnDiPthb3VFm3QGUCqh03gN
TvTG8HZ4OOje58HL0cqj8zzJq0n29DnMP6zMJThv1ShZdaAgD4pG0ZCIZjhvC1xl
ZQMFRFmS5Iaea1pdFGt1DXteicovzO5AMYdnLlvjiT8pj+W3b+x0oOLjXqZRkpYg
YP0tu4jNorimFjP2EjXYgiuT1jd+L7W57NWftbbpa5wVAXGfVqmQmq91syahPHH+
eyQqz0uP95t6VRasD3HbdoPcD6tiMgiPH7cMFKQFrDC958MZfIGy0TuI6PKNhCs/
Qdp8NDEQfqaFHH3uKBjwmVs2p41NR3Znr6rpyRXlwwa+57Ke3lOEwsH79o9RI98e
3YQwqKLIgaLKFigt0mukNslmddi1RXJspcqFoST6gswo2zXRPXp17t+624mKEkKC
ZUnBbJjSANwGcO6GVdzEsH3uQ1Wfm7hYTuf2WXnSSw593g6qvtC4/X9DdTpYH8ox
WD1ZvYy2YJsD+5lfj8kZD4v4FmjdERqOHId6QG9rYZwqKBCr1v5CwhBqnEhzi0Iz
FetvC9NgmgjvOtj9SJvbk9ICo2G6xcbQQs0mprGGmiGbSVWCKTpliC6qqXFx38ZC
phLQ9jj73S7070QYxgKOc4yM7xkjsCevrke8k9yDti6naANT9t2exvw/y8AuJBHm
8ibeWIYEVn4R1FPQO3T0M4c8Cd9torWL5Pb9CnGSjiyvmhyJRkWbI4caTD7CygPS
7HnjKAP3Z7QaCK5f2yFG5qhfIMMmE/noPivn2y7O7K9FCbeerpQQyxGp7FtTqMGy
tCQqFunyJZl8pEr4waHmw5HpZPcdBZW+JM5KCXyU1f6AIMiBv6Erc0BX0uRZDqPN
JznZtPcj2bvvrk57qdbg5S6ApiUvDsHBhOOFiPz54mOpBcIMNfttUbhKEhMiln+O
5npYMgt5dcTaOTLBXB/J6yP/3iWmqg9tw+FSkDjC+U2qwwXp+3SHf5XJAEXI5NW3
F9Z4k75fs3jQWH/FzWShaz04PnCDciC8bk8YnyZv0/8E8fT35F1mO3hPfCKRwHn8
jJcPFdPjZ3EeFmSLAzJLvPGvrEIGNyNyrY1+O6owcZ+AcN0mmyocadH8y0XK/Gku
+suQwgiyQREO5WA/JjV7+bROMCxJ+SzyqaVQ0fMylgP/RKEzz9DQCHhsqcxClMc0
VQXoYNk/XOpcPRy95tKlQMJCIH8v1TS+4YgT3BAWd64A9LOZwLge4qwp4+weWBMk
+B3qf8JayQfRh2/yIIIlnB9IjW7++Yp3zxkrlZGOo12KgKVEx27a880W2A4Zy0CT
KK7wQ/+MruE3+O3KTx3euaTEhTNxmPuiYjF6ysG98/ck70UDGMBvs8gl8SwWH7Aq
GgVlxM4bg1EgCl3J2V3ple0EnVijs1bJPzZIF6/wkFvAWEnoW3zBmRCOVsy3RZ0s
/rokLRajTSEX7PFqaJlmLXyCtEJ2o0SSamSI1U3ZuQ68cadvmpQcG8d1rMkkBOYq
PHrwEKJWMzgiUDEr84FDMcsxM791F5amJyP7yFvVcSGjIOE2kauE7vsfDTtAB2Fu
UcbgLGD1oOnsrIM0e4XA2ZYh/D0txpaNOp1ap/EeHgbpHL+4n3JB/KccXAud0i3B
FAPO4+K1kiXWVeRjvnyjPTMVjxSlmrfUDDqIschpvl4MMDMWgryNl4pqXDCVC1Fn
fmejt9NzlqCOhZUTLyaggQ9yd3wnZNrIBOq67GsJmlkAGeccCnDv7IXHjXhGoe6F
3fM9XGaDO+xLI2IR79/B9l6pDsxFF0CTRlUtP7qEeHuf9HjoBVg/3fosdecj1YMH
KpQGWNGwzk5sq9A9BdFRvVWlHaWjbfREjdYotGvdauc/4qr8Eydl+T6xJmecYyub
/XyWKLL0JHxYrGknb4ZT1fRCR/w0LkyH3k5ccXr3OrN0MGn2CHSpQQkt8n6ke3XN
0f3jWPWkxvzMSNjrOY89jrmapgjmqrPSZB5MVf+CTOB6PnOi/9OAFz0cL0RhHhJe
GqkGqSB/ZqvRYvsguY/iCjp8Dn7xmIC5k8QWDAb+QzstQ4rnUlhbRv+ODdTVHraD
o/FeJ/ouEkC3AocGvH1ZShYeBwrEH19w/qGGI+dqX32hMCEdgTaeeV6yRYqlfhFq
05KAQePNivUPAxXUikiU1Xw2miiu/sBxZsZQmmYHhU4Pmw4DjhJy0vKJEBNkU8tG
wte+6mqvTCbd9eBhOZotzuyy9D7x3YMQd1srsQRGWr17Wo1pjW4SsUz9wHMkAuRM
oLcy8k3A75v9O1Hn1XCeP1FMzFcZ6Mcm+aoZCGKzdcYNb4BMi9nPHzPMO1suCK2I
GNqzIF3Vr7ZRdta0qjFk7qTyTDhFCPYTSFFYR6PFQqEaonCUvgBs7GYNeZL5qBia
wINVNUkAL8OfUdF//b0cwa9I1/JEXu8QQtJ7DlduOsQUmoI0wY4heAOLvpkGVVD1
gn2LBj4iGJ4VnuZOUrOMeTSXDNPbnxfcx16hndhGjVXo4ABoW/fc/yjT4HWlRDZP
clZu6p5bjIABaPAMv0kJArgnksjNWmhgOv3BCdoyofxcrrutl7yVUMdfyFY/+Oj/
G5LX/rUTnTb1ZU+lnkIyYViwOrJw6Fp4n8Y4/rTRHYI/Ow2TpyzN2yq1IwCw7Zlr
37XD+ugvrKuIN0/iWp71HyN13n/h8O9Q62CAovuWcY1tUhjt3nzrp2zncNm/Dz17
JAh6SM/HQlNeWgOeSu+Emc3DrIvUYzN4sSohgcra51A3ISNjUjdUURvQG9jj72Kv
Ea2g1XBhmXKZokSjMrBZAGEVCAYgUIzgHhtR6HlgXECp+PDQvifJEo9/NJOwc0S1
IpbL1oLCi9Y5XRW9+yu8mKFtnJUPMj46iEPoa9I+hSoVvD+TCjqE2pcFY+dQgCq3
hdmAREP5ZqNo/JvtUQM6TDR5YrlGX28ib/7nJocZhmftjC5/jcELzu/UTiGssZVr
0GM2wUBvvB0eR2cmbA5GYm8IzBLTmHCxLT0DuJGitTb1TgRxZj8FeB4yiBZZ5Wc5
2uDDDSGzpcqbsFOXEzkGrKIJRZQgHWiSwHWU4fgW+GoNpRiEtWCe7djw0RhPPmCY
tZPc1asve5e+hizAxgaTIwlutLWIk/0UbtGMMOTTigG8Z3HMpoJdpD7DAx/Gjy9Y
3TVEfhmLnHDCXrvTUf0zPDiRNe2upGKgfV9frQE5W7VRHcpSLi3NmJcRuj/lZedH
m0cVWL41dY60uSej9ijqb3jpDaINJvRzWQ/zPSQjVQLHSGMDj+tGLL6HtMImEgc+
9HuqiDhkAFqQlb3Z4Raf8orGWziVuLwWNtynNookYe9/XPbs1sb+0B5IhABg8xhl
414/usFKy6dKhlI3fqiKhfrOw4UaOCXX/aaAkouvD2aJ3Ryv84f0XxUTcHY8gA/7
jp7StFfGz4Cw6mgb/qcRpksxpBxZR6VrSzMSyV1oNT2xRdJu/Jck1imy1bZPwBSW
n8/qvJFwVYYYuIh9feAGeoHQlqllf91EWkQ464zzWYljP0LW33jMRkhW+TRaOjR4
Lp8OP6YuOb88a2uLI/ZO1T1+FGlq/h4SOxFDfSLLcGifBUaEYYDWp7Xj/PSKtKmw
49Trd0YGkf+BjU/B7/8YqG5rVsxsrTN7i91s7A1UinXXEJo+mLRGmhiU5CxO3vJn
W0JvvZKMK4/gyRiCTO7wWCHontRbDZjdUU+qpP/cSRy3DRxoLJKq29dTFw4BOk0o
b+i++JGXtNjaoiAjK903X2qLGjttDggjPvbfWe8VL0oGpMU4p0ByZaAvCdCGvYSy
cGbZGnpcbL6ZnG27XivxZChl00SeZ5mExBeSwOMOcLgtP32GkcfT3Nb8zwJzvQe6
icxextqAF3BlmfVSZUjSlikmNDQv2onZiWwbfjZvmhxayFCqUsMv/wx2g8WlxqKo
mvy+VgorPyxOPFcUC/F8/Q7sXkD3wNsA4sQaV2ARYnbH6ptovUcEIRhhx15Od+n3
TYREMppwKP21T10Jqj0jktBuT9qG5tcJWyuifWmx2NOLifeD9A6QjF684WpIStH5
dbHciWUgLvwQLDW/F01vSBEobyShOdQiuKdb0oQ5TZ25UZwxX4ERh9+Pc6Z3XNOL
AYzcKd+L1sZ57wEEwPMyV+qB8RzGXb+1EGM/Y9iVRYCrRDOm3ChLw9wh8sjnXl3U
6vGYALMMjWInWyAgmUvYQtRNe6M9n1Cir39mbdY6lV7iRo2QRNPmrbIP/czzPhq7
N4sDTmQQVTlOI1azYo6Sk0RNoNV171SZOGH3CYzkEuvdClTDYjE787DGLb3koiYH
8aZQQ5UFQd58c9rfB7+uHOJFy1IiA1yhCukG5QvN4D7llbXWnmxIrpCWqXRCK0DL
w+TNoBHfbJs52q+5CUSmIgcFZiw8uyB2CdIXO509olZSZBJYJlfYvRLquD3yGv72
7keULOQ1c9b+YpiMs9N/vwNA2lPRpbhqePT9c4iCQVxfBteYBoz0AywQcp8trZLG
LutKL2M7hKQD3wLVYy6b0X76PLmdoluX4JwYrXM638qY48KtIZZK+Q1HOo8tDQ1w
KogUqkO1Hvc9mEQ8ZUbcqdAxvVg8sQw/+g1Qc8pfkzj0G197qLSrMd31PGRAYAnd
of2mJ8+YtbDH0tbC3vjaQ3P6cxCzrTYq2gTpwYPTq+2L5eac36/DdVjVXIn/l9dG
I06KIooK+Q/UAGAAIcuXZ6gX21t78B0TCT4/QzpWFLiBJgCVDxfX4g0VeSoJUDxe
76KJOXuWPf1PgCaFGitU6nymycB1DIKq2b2SVfemb/3X7BZB67q2k5pgvncSYtYZ
TIWo4x3vqbjdZKI9RUUrH5ZZAiuoJJNybTCWAewqOtbIYH5wQJT3zUiVkj7a59/i
GKeLtzpMBIECXz9vtFAbwlUqhHaIpVaNjvkmUrXT9rPa36KbfkOTVd/X4UkcUqUq
m3VfJHQ2apAKlEEAXE1oh2yDC/DLvowE4tSMCA+FjEaQp3uRrtFfs7qrBSZsIWkS
3mStqthsK6WOzGwRX8+t7VQa1VYARYEUK+uJkzRKBWWZZtbnZbE5ylvwPRpa8yfW
9D4UBHUCBoNZbAIbe4KfnP2FnjvxzQnBNiBjOzZrLTB155jpQV+q8i5RCfvEmMLt
75Uzxv7gzK37Es98e39ZD0ZaTP5aJ/Y8299rcAIBF7O0AAjbVEjpXFY3vaodOKoF
vfnCeneEveRcH6VId1M/kx54b76jxSck8UJfCSkVwwQptE82c2Ne1jp97vBwp008
H2eRTkY9FODT3iZtP22yr2ObeCcO5Rv/Z76hS8WrZkB+scoHrM2HgvzBriZtQds4
JI1hs5GeCwfPGFiHjDSHTzi6QM8L+UKf6v+A/WX6FpW3H9Dq7Y1JOKMWsHjz12qT
nY1VV2EOiIbW0bDkPF6T5EO9y22xZYOyA8+w6hUyNlsBw/eGZEynaLOBo4T5nUiW
PqUnzaFRyS1mYfmzAv29R98QTd/aI8A+o2D+BHBg99fttuwkoMcd0OkSy/VP90Vs
EsTXirlTGN0li/0QiDXUVu2ghML79UyiiTUvuxxwCe5YExLwOLQvtJPRWAwGa3rM
ZrLuDdJBcdFeL3iUgjNgQhAIi98SJuPYp52pZut0D8+7QKR7sc2yCJqzgeTNe8fS
GDv2gotk7HLBZIYl8OOIObVHFleqEPplwqCTsOd9FUObAOnTe2rOP8jdbzsgYajy
T9qrNUrG/jpUODdqIP27xGaYPNiWu8t5YPUyZ88f+an6Q9nBXEMB02mj/f5Qom8E
C6PfiR+8EyRdR0Nq7RYw0l6wmd0IJ+DxT2qNI4oZIk3nLPOSI2Sx30Ke+81aF6dj
n++TBjw+/7mmFq4rcenB5r7uqCW27X1vKKUjL8F8BKbF1q4Hl+r8abE9K+y2e8Ah
9tG4MhsxRAui3L74Y5bV9W2AERuGtHSJ3095QH5NnLVH0MKXNwFrW9DsVozHIYhQ
xyPj9qAlx7ES+STqs5W/xodyvpoDV3kHQ7Z2mqPhYCgfxAoCY/dOo6msLUhFtJFJ
6Y6WLu868RP8/HP8M3YpTVgyKqXxNg6j/e0LTda23c2BTf8cfzJ0MSqxfJBmt+QB
FsIV1m8OTX9SqF0xzdJ9+85tfJiyjruA3WvcEgvCTvAs+1MLhXd5xjfv3uWZrCYQ
DK4Y4kK/pDZKnoOw9mC6C1rk7UJ5fk+ZC5xthMLkIQs3Ns4fPO6nq3PZyn0GE2hQ
fJNmgPgtuVGj54H16haw4sKc59IxzaDxal+RxfX20zoAzgkGGt4ZckswtgOb1B8P
x/bfAZV7TK4pfQ9KR05hTR2b/Yf5yZfAxHiLcqqk4yA6H9lKOjl/YXzA1jJU0OMb
/an0Yio6FWtwHz1koSQxbhDy7byhX8JdNgZq44TV/GH+YHDFJTp4/oUoRh0u5jVW
t2Fiporo5YqlXb8px85vb1tn2b7/GpSvMGgQdc3fX3c7+2miZR5wGYFcdNYVR6dE
VLfuqooeyrTx6ZMEyk7xRs41MeBr7z+Vx4nE+v/qFXuo/MZDDC/e+8vESpmdxKIx
TzYp/16BWuEl+A1ap3re5r01lR5VbRBv4mqOl55XlTxTu5W6ySeaav8SkcpCytP2
7U4edHAB/obNAB0htsf05LrWRL8izkLXmncYuNF8MzEAha8rk1hFRlNbhOc2uZaM
svTWkS71G971cOP8/1eDTw8NYwyNw1hSRZu5VBkWF4dNFI2wvIpFtuXxGJ3x0Qwq
hGm1sNNgDY+EKv2wmKyrCgdDVMosWyDeTgHQSUtXzZVPO1OeueTOoCzRex/hBYSv
19sY7ltIjiITiyTjB3YWMgRxWqcXr81sQODpeLha1QEe4IggIFkJbOlePAWm2zRq
ZsKwNJxzF/LH/eYgsXyjiTl59kY/KzcqbkwS1GV+j6CD1hMfTuzTNL2MxpZ5Kq0i
Q3Jwegx/A5/idLvGT7xSjZex4BO/zGQDMeS7s3ioZXHfMHMmQEvVjenC6j601DMS
KyuD1wjOfvlpuTpMKfoK/eLB80AOHE+XmBoQU38CRtjKXRjE/deU5dYeiOwlJ+7Z
7KND0cENM8Ts3z85Ed8/MlkTFsNwqDwfjR1BWPHHl8izgobUgPy9YsIiMMkGCo2u
iLxqqgBhBD9/kUTkQeu990pDUkrqsGqo7aILDczqCCHArI9r/BEOMxmK9wCbRys6
axzdoRwtvYVSGPN9X2bM4NeQwwt0KeRANyNFl7cBAa3ir1rIY3LwRMNvfPqfPLxy
CcbRGfvlQXHXxf+ujmgz3xdgF8L5y3kHkTLMKajdzC+vTy2gnrc9G/ou21eBprnS
ooNhQOmKBxIf129vSQ2Imyfb665n08v31H0LyndVunXtoiSTW+8DnlWCeUUixh2w
z7uU9QxU99CSeyfA4jVP3AlEWdK6Zq0ZtmAWHkhcF0x/rNf+i59w8ajIwGgfQSa2
KhfWJVxZ0/5JhTBuCCYHhBir1kJwmq+SBvOiIcYKN5JOLcNV0tCN6WYPWLrXHqWU
0mQ+7BnuaFdJi5tnL+fMBBBHyFaFGZaXURuC6BgxTz4ZOKU+j0Oui0bMsVNMWMgB
Q5krhJUDAOCoA2Prb6J67QaNMAwG+Y0+WQJVG1JEpcWAauPyjyl4BGvsHR6PontS
nTujTCGg9SEPxgbK0M0RMw==
`pragma protect end_protected
