// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:33 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
X7pgaW6vibw0XbMc4Z3489LiUQbv0QirYN7oV5fai49YDxBJQRVRqXXyBIrl9a2T
d5esfyKixGdi6D0R7Ri20iuu1hDH6ryJ19qFlfY0I9FzrIMFgob/SzFVmW+mLTQN
egWe3Gpp72mMDvEk0EuCXyssNm28LEaWrIdTxC7mqDA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 93024)
BupyXogJna90JBd1NnlRctE3MBTcPrJ9eJmP/W9P6UcXOxPbfdEWPGOBTcsUBSLs
UHK0I4tljf7yDOzyS69UmwfClh+F37Np7Rbzt1U9FWOFmGZ68IBJGerYgzmMftfr
XPnPa52Bei9sCo4jDgbGOoGAO2XEqUz2aPeJL9jPeK6+QodP+8r4Yj75RSsyAbCP
a0esOYjPsjy6dMs9gTWmqlJVtscHBRFvlme8J2V+L6JeHvhVpzCu9zYL+hZUAXmn
ldObJLV43kTMPIjLFux0EEC1Y8TD1hdWxJjEJ23FkHz1tY6dTSxyybU0OwlcI1In
yNfru3uQhJg5skqIv2zckn9qoW8ThK8bOM1qO0gGm+9pU50IxdY6PebAHnqFPd4U
+ugHgmFt374FXtCwsOoxKpzxwFCDu0k5fLgV3X3X+ZFvtP0QsyaG/Lkwxhcy0ETI
j9M/zA5Cb/kSgULZgHvWYlJyYGPQdktvDR6vbQS540naLcrxfS4k6CA6K5K/Y7SS
uM0fwCgxeY0N1eGtjLrJnNRFSOvAXxby/QyDB6IRuI7ctUF06QHUtgRXj14k6d4/
LL1dbngAVVrp466rwiTV06wCxz63zhOLKB0U+nc2SdkIrQdX5iJXcJfLSbs+luvn
0IcSXPoP3F7lxxucF+dJphh9AGqUIhnbqURSYYIzhHcQBoIHZ9noNFNjJtGu0XVo
vNyYjaDY4SJCzutyTZN2QnDczHHz9x+1s3k6EQ+QwDMPIymgGxcBNSP00ypTDxl2
WRt6fshGkDgi6M7NKdAv4jwc2AOpkiQ6GOdUc1vNgkOu8bEd6krLUH2Fj09WUkja
RhTATW37rC4haqQFSxbmUVLoRv/kioaOEXe8ow/rjzSX60ps8yidaxjW4ah2S8/k
yWUxisx9KjOTLqbtS3UA6+bAyvh//Arm2s1yISM4S/hf8quh2KRots9kmYQrakR2
WLwb03fVGZTornB8kKOvvXOwauWBg5h087V4tIeja0c291NBbXglYT/9UlyY8z0X
kjKj/H2KXcotLpqCi5liJtxFWhlc+TcWts5k/c4GEnzlzG4po3UkRQ6eC3rKrKKM
gbm6RaHXZWzuqbAOzqil9lW3ramF//zZ0Aqi+JGqR2v7X1Fag/QloJxzYmqfusVi
+AnwvN/oSqKlQn4AsIpK0ZWU6fKowVqBLtxjuN0jBZXzQPrkrBpJDHl0T+IkZn3b
v6Ep9D5z8nHvXIakadKEHAhYIP8gToVgT4ZpRom50gqSpj3JPN6uL72StUosBvnm
urxRjJcuU4mvO+O6c2KJ+EdubktPVH2h8nmx0MfOt8Boq9X1OFRBTqbZNdGm/m88
YbJUSs2mzmDev606eQvTX6u97biYvLRS1bBqJZ2ASH4qoOa8UaTvSzELcrBEo6Ep
7ayTTOJBidcCGVtWSUYqua7GkIT42PKL/os5ZncdPT8/FQ+2YajEjGWRUcpOQrlV
NpVob6TG7d0kYCs73YroiwCrKibSVm2Js2BDzchi3u00V6a1KRi26l6+B+sXVBq8
cNiJ8/5cYn8mwZ2v5c8dsDw9VYY0mm0Q9QPUzEo3+ENadMHoYMIHV41BxMDzdzvb
n91f7rgGngIyxxRYpaLwQT7jadbdmqWCN96IMq26bskrUXPxHw4oZVrzYgxxNY+j
OiS5nbdOyQKdDStKE9LXSS9Ay11eTMc96FVoztM9cIfogLPI/10qJOtTsbyDp7cw
RoVLRe2A5eCbLJZnQZ0W4cTWBvdM2SZaZajwxIsGggheseLPyOezmPgrnbK/7I0r
taR6XjvWCagZ25dnA4iUH5pOIRC7XKJC0C7vuAHV/uIL2CLFGYRLCsMgOD7mKVqz
+5h5dY7HewWxL+T5/kQ049nDs/cmhfZnyM6oE+m7O6TCauxPIVrjA4AXoXwyUNg/
E7Jdu7sgPH94BCHPW9d/nbFXQzRWpMorrFToCK0/NpuV+kJjJBPT5hBeABQnWWnM
D/3ggW4u0WcFHgOYmDlTkEb5Ubiz4EgmWSatZpfB8F2TzJ8BjWfpNHFoKkPXT5tT
fpCHipkpto14Ke/e3oduKGjPpZFGO4Mu4FTXLtf/pzDUbOCJ2/9/BjCJan4IDOUt
tDvLua10mLzFm1ft2NUc2uQxraERLFhZpwuclq49/sfegJwC0+ZxmrONW1uUAvKZ
IX/r0EHYHX2m5ndsEIvj5vodHmw8KTap9BogmBkks9yrlmkEatxdk2wufywG0TbA
3omO4/EpeQuMUIBhUjjNUez+j3OGpIArbnTUQ+a21f+WLVf5Z+wlfKdvmjONGNlt
KnM+1R2hNgC7/fWqa2D1rhdVGeu4vaSUcVlIUfNtAh1u32o433xD7LlEMKoTmK3S
ir6s84zc6JqqE7kcVn6Q5u4quLdZFv7Foryu9ps9YvJStBXrJY2lHp/t+LdNQggM
lp7Zetpg1/G6J+Y9TyijrHiY5Yue0WdJI+25ymgKXHPt3nCJWqnwGjdq04IWaYu9
NgiGig2WCqfoQd0xpD9OPmaINBSkxyRs4YCdS0V8bNOZOMEQYBilNVz8N16y0AQx
bpsALnEZBZhYmrRQbNOuAgZlsegMCigbWkj6f+RtkiDegBaYKSHLTPYqv36qBG1N
2bTBoRrBhqGvnWqZ8HCSRONzW9B8ZLGQhUjeLVSr0d200+mUFrRvI0BXIBizyC7+
UeIL96pPWVxsUNhLzTbmcZTMEqlHoLFh34gGaQ+AvAHPc705SHVgdPhMS0yLA4i7
m/94khxRpaRi5bAlJdfK8lTGGGtfpi1TRZizuUw3FTuvyErkiZeO7YJMk6o5DYRb
fqBYnHKgANjzFMUs+h/T8IaT8m/JB1cyyW40lRat0eFjQXel4pKNPANiXyruWZFL
tTZGR9UhGe//6PyMK+RmBtlEDg/zmcDb2XsBxJo+XHHB9Sbk4Blh4VdhZ2R5znHG
b5dtOJTV/Sy+Le+IcByFM5bQKNvtRG1bL9K33zHhbmZPzEhWtxdT9Jch06j4OkmU
+3AnblefzlE1sSJ6FkZBusd0hz5HkXEUNpJVDIbAROY3PmSZVGn1lpcnySMJERPZ
r/laiVEueJpdVeA8RO8Mli56pxXeuO9TVg82ThTEsYbk3T6YAhiC/iBYRTBFnmEy
ovmSTHCtywYmC4ksg519bGhYnAI8f7FDj/8LN1LCErFxN6g8tNAnRnBG0BU8gBXm
gxoe8403eFxxjyykkMy6BJBLFN8YXBhlrFCguS6T78oCAlM86vA/VN/PXcMBRnXP
fnzX6hwvfrYgN00u0rn5OTSau5Ot+PavUjs1zua6VULUYKEZAOBf/z6B/DBXCkOh
iz+amygu/rQIFaiAMb6ZP4tyJCrsBwNZANbrgsGLuatBw4HFASxC/wt0c14zb+t6
SWLNBBQHAMZwy08UBkKYDDrEPCw/8/XbS2Uf5oRss1sDiM9TNHxC2HJCZQ1IMi3G
jNlV0pm0RZFHFDJeNnABdba/asC8S0n+31sTlijKZt/g8n2MxXpIsdWr3HoehekW
GAoWD/W3WDaDu6c04tDTKSaBmHG4EMNtix2sPQv/3vxpin2FYBYCUdWoYKGT48I4
my+d5zm2ml72yFkPrbUgGbu49HY//ozWwXL29f5LxyLEMpf51noGg7qFxj1F4bjV
tc30oTTIU8tL2TE8UIAnp1+Shf/w4/aC9d18utLOFBg4kCYQKCOl9iyBcXDliKDD
JZwlJmC9r2eYop0hMnZjlfaOosiANP2HOCWoX5/1bOWH5iAzacqFIGf41wR5c/R5
JTPfUevdtwkY9uAw1upI38WF5wzMxD4dkY3z+TeTJghQuKmSDfvmxR5ZdNzslY3e
N+Ykb8x1PG/1ZfIv9fmNvFB1mXVmOYoS8mK+ISiD17LFWgJDlpfE6IVQRJ8YS92d
cruqKao4V/JEqRppmLgC9HJfG2GgjY5xWoCzE8DL+Nw+reOkb5A/BA6MqCO3bDkR
b2AfYNmpCc8GECZcwiOe5hcUeCGo7lC9/wBChI5LOcQYJKWvBzdLAhZAujbR+iCQ
wE78WfNvOD61Noairx8FrMutLE1fcM3MVMIbEl6K4ukUvyoh4ShIdoRpVdjQw+eE
TiJd0bBmYQxM3kxDYu11zjMTEoBn+eAI/fPHKdx3ZwSuJgqX2zstLUeB+hxkaISv
wv3odN3BSB38XkfOuSm+CeYyP8OK3shF70ciFn0PcIefjHMxVJ/gqvPkutwlUfnI
x3gBt361YBK0RuF5EdgsSGeA2dDPSUPG5yLRm4aEDFTihSFM0qFkELWqABJLgPFE
+3SoYymvbTJ4yxSAUY/U8FiAUl3f2OMTVZfyTuCHRXMOMAZEY+zUDcnrdv2scLNJ
Kp/SKqEFll7t6bvy1zu7orn3ioHT9+V2AY5jaAY4m4WMfiQcyO3QDOFz1HlmpmFQ
X2mCw9PelZMF/dJxoNom3ArZI+5jcbuuaIWxWBQb+yHIsw5ZnaeqXD49HZ8o+gko
q7rEVtRU20gp1Kx/brKeXtIMJOFZLBeY2iYcRRjGAi7bJOpsGxwkn9S3qGZ61X/f
UPjwOjT3pIN7cIPIBoGgsXVoqqsT/nGZRLwovtL0l2Ynfj6PJ7wxjHml+D96Yl1o
J1juS50jknFOgAH2Txi01m4rp67sxvvZLs7uXLXZ216s7SAc5XNIJt6jBvxtUzqU
HgHIIRca8GKZpaFA0GVT/gNskYOfxb8ZGKVKi8pZ/pv7h0M2W1sNs+LCy145ANdD
2AAdWzzd7JusYFtBgBHGZNdknkZmLdyXSqAyFx2JVltQK4ltoZbr53lojPt90tBT
bNcOrkZPrKXDQoerFfxPgCLhHAUNUUSMXJ2Yt7AAAdSoFhmjyi+Er2qgH32xmJa+
VLD0+/p4eYa+PUL73tBUyqxdEwkx9MAKkrMynFglf3Y3VaFoKQe7nFk6br5c/3OC
+huoP+OL7DqCiTgu6Pg6hm4sw871d0EI99nLZu38YasvRmlWIZ+r0ad4zSPl9WhQ
WOBnS4R34CpV77tEe/S0Z8nXYLX9q2BlCTHEo/TWiTRPrUz6bZET6T2bU8lJri2O
k9HtVXsHGW4rGv4+bm9jTzZsEs3vekTJRZ9tXAz1UC7KnAUwDEtAIe7UI9PNwoc6
zIaSBI3/DOnhW4+6Au3nj2O4nTg76K5ZFyx9zWlAlbqrcozF1h9WMP6K3z1DeB4Y
yei5Y3HuP33DRRpPEZ9+wsws+9T8cwHUXc/Fa5q0SW/tczpF6+7kfclH4XDiwrWf
UtFs+Ee49rWGVF8hoM0S8ABNFP8v4ZjP8UPWBFlNb96xDfTchl0IacqftDKG0o/4
RpVQNaVw2lK3KkSYIwiMsBb1lPd8L0wbDd7VlpXgNlNC9zL2g91+7AUdA6bfWtG/
mDNZ0T4tUDNfYp+Fv3GSzFMEp8U8XbgExl+855PhRlgeQS3GwfnVVmvC1uoN73Ip
hg55GBfCx8Gt/eQ0u4qeOpnTuEUoW6rmrp5dTg6UjO8+rlXJEet+NAZFHuRS0xSa
u4PCn80rFRrOhRD/1hNgE+eVlxt33wbt+nA2Cc1w/xhg0A9lAxQw1kevT/x3P7/P
/VJ3Hed94Dgb+lWhcDfRk7/uNbD2IR0+06vPDA+6Oxn+ODbWkQVLri35cKKi9HG0
BQO40OA/vlVXtLie/mnHUl5kqjRwFinolHRpmYbiI9SqtNV/RgeaLm+cNCAiWT5U
r9cMYsXrvCuhHZjjBPUX/i13w6pYVfHanBetIq+/BY4UJqNqvsM27s7PhTSUFSqV
NKu0X7FrZZn9UewBgaOqZFQrIBDc0TK9pzhIqWRd8vb7adHTo4pS56eTljTQQDmC
HhGHDmJdETPDdhA6qbpZuwKnbN45WjqW/C+kwlW9ccCK6ooXtWsF/IomDmq+P3y7
xCORV7CYjutjNBHbHaKJj/+uFcZHXK5RhglRzE805AEw+Jxgw8NNh2mEVb4qAQnU
zU3zq17SLQW/yQ/IGOdcHz5NjZl+fJsC4mUwqpbfx1MTOpdg9G0+8CHKRr3EKRAR
cU6oADeQJXGuSij6JCCE+mwrhBr4opC5o/R5DiGZEg06O4EFgw2SheUaRnM3nrtP
J+Rc9zhAFr8wXQyXaVeXS3Nt0R9IrvSlTQdP2Y1tSXZ/gUME7Az/XY85XzdYKyxv
syIW2JMsKvqpjAUAFyvIhv4DaV0kzmAmu/BJj5Z4zzX1OoJL1rrONb9Z3YnV3xhA
YCSY7rYLcwiTWnBB5f5D+4Z0BrBjqPYzWZHjFW+A2IqNYgWIrGJ8uS9Eh2ZqLJbx
Txx2Y+jOYdITjCev3e0flqqfskp+h0TG+wTHV21ua5WQ1I8zc4HMMRx3Jcu+ywbs
sBkVfEmcQkW0/hxHAp8HEM1IKmLC4fltv200l4Q3z29PyOxzFtKi8F7LSME0Eb4+
5c6JkWtA59NuqdD7VRhlyoOUi7jLGDMLYihHRE/UjZgyhsyWODs8xcGpnVbCpKd5
NOun/ZIknZ0vQeUJewgKqlhbUo9PeLYOwxvv5xfYRkgYpcwfWLcp7TfQWeiIxLo0
RNq/iNx+4UPXorWNYbGkejZHRULs2nlqr8bEVu7Np6n1kwqHncT6jKYlgMpV7ped
im2ftzFw5s73LxmlUEI/2iAKg/kV/xiDmp5xNXbvMO9lru6SmqWfMMsy3xijZWBm
nfzUCDtjoroy2KAvkgruap+aLYooC41u9yvGfbkWp9Xd8pjgFwZvpSDPutqOXPJp
dxRmP4pMNiGg9it5JG4D+ucrX1tLMcofv4k4SU0JoVUyxEnU9huosQiHIEDFkHiX
89+ghnBFbJgHmqUhTGmMTAODGL0qB4+V4x2lD/yP+vDIamMRGTO9cLwwtFmFbY9y
B3fKCVQsEZfh9Z0T2DPRXGAoloIhk8Cn4lPNZkYHpKg2mC0qdjk5nBUC2rkqFVCd
tEPVmiXecIqZnh2d64BLA0ew88pA45IjpB3jnGVoPFxEMZfQk+1R82Jw11KuHjs4
XXldO0pwnMMyEqYg7IVfuInvUaEjF6s0CTXwa3+1T8dWWcJTa3BMpgox1qkW2HuA
eiCvbjTgr/ySaG9xOCrAqSXs89pSMYET6pSfSDyEMofKjejAe0EETqGb4vDIHCGM
PjMXM2qD8d+HQ945eibpZLZD3Ct7NKueULBI/IrZDLQaDKC25NvAjkxsaZfzEJ0F
sthAE8sJVHHTcgW59xXYVfDLoxMKnsEtNTJwHuQXhD80H0ioybtlhZMf2E8pMcFT
o9C12TEpUgpG9bzv3SuhuQ3fkK77TzzhHsu0YViLudK8uGk4v5Zwf5RkvDY6lCTd
//Cx9kbwMGtensVPOva0O/sO9sEd0PbDvPSAYHtF9pG7kOa9wQXawV+CF5ipsY4V
gv9Cc0QZewOOqATiMlP8GDk7J8DCp38tumMm7SOu7ZfGF84HNpMglxZ2dVCeUJy0
DBMXGcroi2CCs4Z2pcMGEuvW14eM80/RA3oItGN0Bh2UbsXkTGhQPvbQiHUg5NQd
7FsmrfpSrvaO23+rEb6tv0WYbkZfF/CoDqDfpKm4pRN7ERn1dH1AGzHjuILbmHKJ
ENqklBhfjm6X1vOHw4X1mSJcdfgj3ruVKIyMqSlhZV3pNhjoiT1pkrAJFKoQJWRb
llX5U/VGSsTvJ5uxrgKNrnYj/sCMICtyh6MkEefU2jNB5RhxRkEVPVTGREhycQNq
YTtKRy8I37vLnvWigcHm+dujspdVS98SoFscOfuVCo4/ABxm6i8eCU3VZk7ATIzS
zyrm2cp/ozWoHH4ZndU61s61nlAngfNbe9vAKzmA7sePk37SyG1c7K4J3QMUBnHc
VRmuQjL9UCHQqm9gjp2w79skTixVCxyMEJlMTESPJW3chVVpyLHVYjwwDszMacsb
23xaDF/WGZMccxFvys7XCM6dWcurPCtlx76ItobJl0m7SWKxkTYEveXeMpsgAsd8
u2VZQFzdssYuwp7dMa1GrpQ96be0CqL8I10mLWsehpte3MdFHVWnc7Ku1i8tLzIn
y+r0WxQMpG7KoCQ1tFceYnyh4Fq+EsxhPPSUc+40Tr62o+L/OdIVhsFBMCAAFpBK
tlt0Cs/wWvgEK/q1vrIUsdIj2O1ydjlBvXbuuLq217KDDSm79Q7d0whCuFkjyRoa
ndYXynVpGWFJdFbKx8saScU6jNRSRdNKeRYPNKATbo/O8HnFlhqRddi5YDmfZtNk
+XL+shP7xn2JFePyq8UGWh+S7zg+NVN3DZ6Q9QJ2I53eMFIzcyRpyHpyRR431b+2
QUUbpLMpZ5+sBhM+p69BM3A9tmEFtwPhS5ID7y9dVUz+bj+HwjFqJBnVI6z7AEnI
fBfU9qte5/bDT8QvRFYo2j38QkHcvFzJSrqygFikWjdWYZPlqjWQ4xNodNS9kOwS
x1Wj/JhprGpk+fg0rjvXAowCLfF5BvkQRRHnFoO13Uzceq7t25EgMvgwx+hQCByU
KIOZbXlcLViKxqlM/kjKBIJW5+eqD33Q6a4oMfa+ogNWb5iA1mV0AsDXd32UexeW
OkdcO0Vc5IVI/HTfJN3xJ+kfexJil4RznqcyrrQXz2Ry0vBDq/kE1yzRvA4CRPAB
KaO0l4JfP3iZM2ENSpwhJkfnGFP0OQgeznc9v5KsSvXx2KXy7fu+yXY4pS1krjA9
/5bz8QKzUfnsOJyxs3wm4gDi0HOPLD3OJB4HA0DLkNx/106ac1wUT5moz8x9lWwq
IKxAS1acQDk4xWb9x5QMxBMXHvSaXLEKGpNrRkFz93w0h/0HnPKOrh+hxFZ61alV
uDuJiPSL2Xei+2HK55RpfINqd4X82Js9o2ONQtfakKWvEChl/7eTxMFKFbTH+NIF
Kim3mP/pO72eO353YtnSoZHVVka3GxizHsY66fQnl2Wwl0EDPYlWK5PtVr6EUUMF
yeimH+tYDlhPHSAEb0j00pSXTKfmbZhrzaDwUe/xg/vpJfAO+3ka8Y4N9ebHVAnc
9qn08dPTd5xPLUS9VPaorXzO82Dj3xFpzYP2x8FkMvyECe4BHZ5eR0vRO+HC9qZO
A6z+nULznKnbJh6OsJYujLxsjN3+fsljmPHODCXOKStvoJzEzOTbKM9dT5ylsYEW
NZZ9lxymsteSQ19ny1etANPvXwGA7dUr0opkDGfQaVCqtyCtudEsvwblzdU82TD9
U36Ef8OvU/NCA/y41YBfu3yD5eZ8vP3ZEOLkGmSatZ/fTpimziakzaJdklh3MU62
zt+9UZuMMgaTvoRouKMJ61KZcA60+0Dhk6o1Zyn6UlqLWfmrEvVFTUh6B57h3otj
s3f1oKloahN8gaEiV0Ppl0kLm7fQuvKNd1q/3K2H0EaYh5TItmnv2ZhSNeueVLTs
17H/mR7XcXvTyJafkx4kiV9zBc760Enf8Qt3ON5S0Ya2LLRqCec3hoREpKU4Qvyx
mXvoLcawpVtFJo+iTmjC2v9eCkJ38AWChDmFqov36GupZffvK5fasYUxlkhg3H/Z
jTXjSVGNQ47+ZUGHtJ499w8xuNwew9iWkgr7xPWddOYJlIc9L/xpeM7EMLOuFzSd
JTbfl/Djtsw8vyddBqOmhlThSk8FkFGjiRz3jOgk8O7CYnWQ8t7eBn0eyBQYmGZ0
zADAqoBO5xt9W9YoVUgm1TW9uXbXeU7ayje2BlCAGNyQtmn0A9RkOp1aYgS8w0Jv
yFTr0bCXseIO61rK3kn3lxZ/P8euDiw8fO8nn7NEeYcAkhlu7Cjz794cWnVecEfb
o8HIhHI/ktwaylklmZlhUGMUc17ERoorQWiCQfkfx1Qrbc4Ca/j1zfccG4fL4tBS
pWavVijfCOPbkjeMMpzF0wW744jyR+q+xJy05tvFHWVGI6kH43pue3fkBy/L2Dac
foCAb2rKHmKNx5DX8We7AzRg1kl8wcsMwxU4EsirWM1Hzh32vEmn6RZ9W/RnSSU2
bqrREeISqFXe15llZEzPCH/kwiyo4f/LTXbIZWCYoBjs5i/v5ki0KxQCu6UjT6J4
vjWSmjExbO0QQG3YzfxSzlQxiyehACmFyddqA30KgyMMktJubfX3Duuv+wWQ+sJt
6xp3N3ronME3FP8lTlvYwCLrZAvsySTuDE+bXIdQYMoGV0cKZzj/NszdSzENLOU0
/FoG/ZqoQIBAnMqTZZJ29LEiuOGb4CC9bw0zgMRcB6xYs6s8E+fAbOCHv54DHgWZ
doIjm1ATOjW1umT1IGOR639iZHOOWj6YC9Pv6FzBdJg252h2SNDQNNmUeYe6PuIe
2rUGEWAQDpJEdhcVmKqOsDcI0DibUaQ51RGZEZdMDTo7Y9ybO6v7l3L98t0YbrnG
2+Wh8Bku8Pg0Bf0QbYl/D0l1DAuN4eZWB6ATD4jl/bEFgQ/POPlgJuc8e462qhW9
IrB6qbrM2h8VlAzB/97k1HB0CW83XtwmnPQyYUBgYxNdK70se7FoR48D8CQwsFw8
UTlSvrC2jQE34wEfztsmSDafOP790Hf6melKF93tB/HSqwpEQYWrvAJrTtA22Eoi
FnhySNVBofuXYX3lTr9hWnN1fi1GuBeLxjZWHtC6BwQ5975Q3TbTKtQKG2Xxopeq
Iv3MnKFNAr8AjbiOjIBd/KscSCV0BsC3ozBsk7+l0oa/F1lhBGY+i2yPVVRkupQH
3Jq58DjKRMx0LDxS1kwCtkShiTeQsGhY/nKpMLl4Q2yAGTCUOcKXeP9dezMxXDWv
ldbYb/3ZAQFhVLE2XmycTFztnV181Glvdo1FLUUKIZ47VihmR/kgkMeOwAkOgYhv
rh4q27Aeusy5dGK6tC4+X6gIQwKIdOBF6dDURo/vZBX6b6rq2sbviZnBreEp2OsZ
I+nX1BWK81/qMh/3uXsmFTD8q7pDoZQAhWYcIPUq6OwoMJmsbVf9GgsHsIt15GSq
X/H55vYkfIjRAg45bGO2d69sTi5Ud63KmT3jwemGCvNyvEW4+iMIUxN+toYtTqG1
5UJpNzB91rGMmvQ5MVtHo236VjaRxawGvfK/y9W/TI2NFzqCTLURx/jfKyrApiHj
d11QSQ9N+cDfABnFjRjtyzc2xbwFtZlqFlKibn+srWBaUYItIuKDyOqkZ7rlSJ3c
iinnTRqcKTKjY4JllKMSUBBxzwBTVbOcwAN1KFnuIgZJqoqovondW/xzP33OtCYw
mvdE8MEosPm2WjNDrL1O3ng0TL81eIMEFedECYkwGGaBudL01nNBqRx3J3NK0rER
wutScNyXbrr5o1QHcQ4B8nuBAfFYR3hvgUR8MaN2I77RuX/Sh6kn9ZVQFNYHO98V
QFjdK6P5NabZkxB90ojpJoFcxt4Upj5V0bFqIcvCfGpPAlhrqBsmQitUHdJRqboW
eH5Ks8eVjDv6zessH07xWIPt7mWndoChJnt+vHSlKqUWcL+HP6EGUGEbE+WPRuUt
+W0/KDYy9PiDAMWEvLAoPjmPVWC+e3ihNvdYXcQs06hxajXsJ+LtWcslW+8IhuP/
0FzHKBCCVsr4Gw/NG4mC02tU1nIwK6Ls2kq+0D+yodkWd3yG7Iwrm5i/+SokqoLE
o7P1YBWUnT87ZOLA8d3JbNvVOWELiRWKLMwnDwIlnads9R8BjTNyX5aeV0pJ7xKy
efBed2ROeiXc3P+E1/RhxuqctJ787LdCwv+68Xjr8rZqnYh2TgkhWVYcVW2SQMYO
W0JYTHpGaq+PK3mJJN1i1443AXjiLYa8K4GN9CFyC7xQ2uRQfqxdUYrnw6IJBTb3
yQJ1s8YqaWSwpfUMpmw2lQngP+V3mxUodtD39RsY+S0Qumu88sIcAeDvQyzRGvqV
AAOXl58fKd1nAAH1TwmUmT5JVkWualjlJAzVDzEUasFA/Y9Y8PBPY0fC0dGZvSsb
e2yofeWXoJyleWQppcJEiO8SSPz76HRVAMaYNC4YLuRoUbTB1S+4ZoFtIGkSr8hK
AkBqzvbxHOfStQzFczjlZpdU6Upq3X950gBjAcnBiIrS5TtVNaSDY0ldANKtEm9g
Vwf2/cdL1FVrdMpx0Hk10ee5lNxkAIXQGgq+sG+pRwrM8sEylVWC+pEj/dBXtjVW
brcUjcXQkUFAIoKwaLLmFg4Jy2sYEB4MNqwOtdWUyip8dgGUKtR7YtW/na1Ej778
eTlYS7aS5CzdZM2bTZDcSrIwwOnr/I2bxVOHV3nAxLy1GIjFgApPApqE2dp8k6sC
wV7vrz/IXAKr7HLwXePG7JVQ1EZO8WQWWoZyzaSejH0k3i7VkeboAcg2jKfTPMQv
AvoapJeMErXI61DGjeU8q5zJ5AJUB/LKRe7Khv7jp9nAh9A5L5ouB/w+Ns9VPMm6
duTHyt14CJCB1+fVNQeSsXDTnxBfv4XxYW81exg2c666w7nBvfJhiiIxp3k9CgHU
Ckqo6PrNxWajCT9rqNsIuE5OVOi2heV//MCOp2D5AcZKGN/JGysNNeT3MrBFB+ZF
NfjULDf99/65bDh7BPjMbcYYQpq4gJwOxiQLpjqC2txjVDUlLZGLYkK3JdOExYdG
b7j0sOPOcWG8RCJ3ctSd3PfGW3l0hJqrbTPsgju1DbClIeCMU84GQFhYXW0J6XM2
NyQJtAIPTFCvywNysw4U+/OmLDYnCMv+9LlwQJrjE7uaL2bhTVc7H3Vp8TPz20UJ
qLFhZ7D1t1HVuU6Zl6efdjx/Mfr7CZrNOdoITiAwCCWNp2Emof3siZN5ftHJUXgx
pzMSGJ7CZpmrtnXM5vtBs0g328T8cWPFq64nJPt7xGVmoT4K4VyykGh5bu5k9QFQ
SgNgswYwlbOkJ+D9QVsPwODUL4V+dk7XT0Gt0U7e6NoHFegmEm5RErvVIfdaeI4B
cnMO7OUI5Qqdc3RffjyEz+pmksY0tSGKg1Z0/M0g2MIUMznRxTHHdd37INIMeETG
OPCCn3oW7zE37dZj5yp4rBBhR7tL4QH4n28jzLPnBa4iLikf05ZSbl//xASFnjkj
kriWFXPhtHpFySnYI7koaASuTAT0jsq5gh+AemM2bIFCz0paqiGEuFaNXjewJGK2
Q3aFXrMcxUsC6H5aUaqqUkqrHwmZ81VxnObA1NQ8ZUZZlJWuX71vvcsvb45h/dVB
B+VsZCt2OI3Th9ZA0/YKf+qJ3T4Fhs+bfz0KnU6xYp8t2nZtgpPo/n8arHMk7UVv
7J+MYTCAE7KrJr+W1mQHPMDQZm+O/f3VSr1e9QDPs4VlQivppnWBTgS1Ef7IpxBF
ojeUmzf/QMngA032AKt00q4ij2ZyEJjDc4Xuzr0LgNfLBUwJpcjyLENkA1mEq+LI
jMLQQ0dtvUObMB0DwIumKQB0/crxal/ssNjBdOtH8GkGibFPprtxrjHtDQDWRPaK
0y0qkgkVkk1efsJKc58wg6oatkzyZ1pIpOvsy0LLf14/et2tVY6nNYwLq/BK2GZf
XEVJSTu/gW1Yl9d0+AcT92/61HUM7IuACTZF2sJyWAkLUwYqJMTtn7F1iQ0kf0x/
JdFYAaU/PcKCQFAWOMgkQKBuBqKvsijWYbrfIQ4LDgOzQDFgHZai+bb4AlQPo0iu
7QqiWQzG8o+ipyz8Myi1fqekW7JwYJJyT/vwOiehgWyFytUmP92JWrFvbt4v6YVe
MdbZZ697WtVTHG1bwIVRSDo8JfD5E7yYXsYYyjTbLgM+cwMN2m/Lmc7CpeqU4wAi
CK/R39MEG6V/b3nON4oZxcZKihUbHKmDFC4iSS/aqVpympXWP+SclL5NHaQZjR/b
yi2JzXn5aOuh3POGg+TyTw/Oe8fIT75XTRLyOJbAm0GfgErIb6VYC077cuGOpP34
QKto9J3D+lCVrCSzlPVVeWViKjvbA9inPS30+iN66KZEDeemPPDL7wFoIHvGm79Z
5qvdj2TcEzN0RPdGuVN7GOSNpvHW0/rNOB9mJOBFbvYDjWojA8SJ7FvFOPFzdrzH
rTrUChArgxXZKe+tQ7HVvTFNUdYjlC9Kvwv6HWCnqUYS5Z/YIe6I3LNZJWwm3T+T
8pxCvxphrzVOIteOhA1oLFAlf1x0Jlj2YEOaPayyDn9J4DIliynS5F0jSXFjT+qA
tDyKHwSaK3WJfJzVKiX/HWKOlxpSrg0lYs+oZmHUKslJaU49H9iZiZt6GeKxYHts
Tj7LgmSmp3r1End2VV/cc//fgkuo3Dk9eJ+0/LJKiqTlgRXBy4WEF6ZCVQflLJUC
3GjTeAfajZsH2JN/5ENEPGwX8/D3p7pZifeyl6Hzf6eI9zTp/zoJNfx+rUgNSkI4
k9lNf0XiIJufPKDdB431inL2hgUcuN01I1esnMfSXr4zCmo0NHeLIYtgKIje2Hkp
umuDvSzwM5/EM1eoAOSsJ6o7+Sb5KYSyQS/I3C7pL6/1eiOh8ch6qaKR6bftgqPe
pi+Z7+n6NYXNO+A9AhnfKnC4/5+q6mi130By/B7yFFeZYoZfv5UdODSUhsrqwN17
M+nnOfn69oTnLYBfBxKIotjXVUYLxhiRnt/0crgzXLgBe+oE2o9s1tid371xojSs
lfRvIeT+qYOvoIKvgOMfl1JZi/1+35JWnMe3/6nx2aDtV33XRokL+B1WuuRTJZAj
EcfiyMHkA565aawXOu6vS4XjIrGKj9eQVVEIRWOPOEgjsXpzyTfjV5n3dWzhR5kr
9RKCn2GUvT5q/ObDnvAY8d1801JF/bSzb7o1KZrbmMsxoQWjhsRQdUdJJ2AH3/Kz
QHR/jUqi5tU6A2StKUPkmnMSVkxveMLg3HNQWWThW75s7eeXj+UiNhH875S5Lb0Y
m/uP4vX8ADLHgv3W9i7r/O58A48fKsUlWy3vbCJC0rrd6JqFldpKzqZvqsvMZ9Fu
kdxzNfcuKjYqXa5y/Vd/6cdIPDaSL7WZTAdv9+kbSAwQg5u70Hc9PDgAzgQYFzQE
GcsD8KFW1JCS1WStsCGgXFlSIKUV3ZZsDng1Ik0rbOsDmlwDU9nG8Tr86ufC9mhv
DYxBDL23BkvLYPEOzje1Otkh4IwtUmcUlOqVbxUz2xpXqccxHZZP4qzqq9647f5Y
Nf4cQ1Q9bkQ524d9MsxAJPSs5jKNa+4Wuq0KPW5oQao1knk9yCUR86gfBZty8FAs
AbEzKz1xJ8rn9imF39+xDRx+BXBDuIGusMfCznnlhyiRpLe3x+HKVL8j7AFDX7t/
fpjM16eyi81SamVoAujbbIzCP+O+F+1ELKyW+7XeJHGa79y8vavuLEvJitxlbxqf
cYiXdBGfsiPdiIvdOh4sfGEhODgU5AAbhW0o8DbnknMWVMZclLM3KWP6gcpscLYB
TfTcg1jl/gsMhrk3eTZ1MpitbdmoRAnnwDBSNQSS5nWmDSoa4zjV6WPU9IiZUjXt
660lf7uHhmKBjFLx0jZI1CY4rHy1vI0dPWZaOzMNP6FhxW9N4kyd8HLeL5lMRapi
hSCi3nNa/tx7Y7RtXsf2HG1ItSSIr/n0icnGdozOD/8HYLn00DpesVipMLZBVc/B
F+XoqzL/T4zRv8sSarucDvaL4fC9YL7hR2HF6b+EyIY/sBj/bUMt1Aif7xUFTp4S
sPDXV2u6TrMiW3ePg7iPfJ7fKZiPPZLbijSXsow76AijR6XVSHd08Annfl0JyFj1
cSMdsFywfbiN57OCZnuipSXoxu/N1kLfkuP5VE5IQLJ3WS+k+dT2dJVuDppO03E9
+hqAFUJB4G4LsZ8y8PlfJl9OzbbscxRbkf2dlkxWI6p42gKCF1X3Z2wocOk/VzVK
cuwWZPtvGIfZVrdJD3bQmq/dtRN6ZjdfAZk8yrmd1MXTD8HFdG5b3QHBN8MGHYvr
dphlTZlvXhqV5SUWZWqTrRf100bLsi8WpJKplvMKBzRRhTxXtxz/sTdFMSD8W1pW
qD9Zb/sRi80M6H2cyGA+0TH6j902XCf98iFd4cW+xqrEg9kmNBHa4cUqxFyyJpja
ABox25SyjqZUP9AqnjAxIw9msbN9n/Ep+AUD/QraVCS5jDdsZ3NogqPl5C7mfqUI
x+OArPkDIScE5XIYqVZp2mQLSP1Y3BjxZNnUKiNe6hj7P8KlIptjaznJn7vJXysD
RBk0rCzDegBJtS/NLdBHz2sYObIA1lLxw16rD4vAyqApH7Fi87guSosfA59D0gPv
aLir+dl3UXO1OgJnJElifduG11rufgbnKAThvO6triiXKdodDUAgGuWKfqxcN4OC
Q8v27LftvBxFBMrOFb4W/gYWZmPkxJDXlIjKS6bHUFbVlckpdWN5nLQWWJgXwWh1
2kUEPMmKU6ncLsEHcVHrpHx6q42jA5P9zRkYBJCOGV+xUXbdRRRPqEBAQR/QNe8w
zNfnjr/wVA/1KpIJcYBm6yM6afGf6DCkAwwUNvnEtlCFu04KA/TOgnBV+5diO99H
/Aw3pp0n5oMIMdA0gptp6topJ8HiUb2BHfCuEjTfmUK/0CdM9dWWP++c3yb76smb
JTcKXwq20no3M8nNFQkfbVwYQHcReTtw9oJaFsTrpzemDm8tYuEn3EaegY6fwMqz
8Lk7u7CjMpVQbtm8zc5lXIGE9zC8H3UtxlnpzBW8gxYSvWjydxc1aI23U1k8yIH9
eBI7uiNKl/eFwAB0zBGf3XIBDPYI4JQHF1k1jNXYfwLZnt5fqi2KVyGyQMxSWsWN
5o1ZBtU+C37cnP01bRCMeBbWfqSmNYef/YrHvHGHpofj1HIWAbHUHnjf3g0Db0lR
k6Xqdb+p80JCFifPiFYIfcGWHjhK6oRuZFLAuYX3Khd6J592wvcgtmUyRzUJbSwn
R5K3ZhGnPZA2yLwww5hopWVxj1PkWpCX79kmnCb4SVbasRKKpaOxEhs0vdsbrYZ4
gsITlWkZ/31yMcnuGJhkKXZmRqyKeaW3B3HG4/RM/cvPD2/p8HDVrPO7wKKfIPKw
cMjg6gVS4AGYgzw4v8s1P/8YHbsGuP2Cp6Teh6iC9EmdKW5LDBUWM7nirif7M7PK
ioSc/Q7KpejfuYthCxwskp6DaKQo0jXdpShenzwa9n5QVkveBrQ4/zW++KlQBKfG
J2tXuJssRwZICjD/MvxZwkyZRUFEPOcpwqEB7XL8XuygeQ1aVjFAIqHtvfSRdO/k
UPgctsR09iomvOHluZVxtq9wKZgu6SHQ33YmzBN3anTWLH6CCjHT/un4WVN9pNbH
KO40kpn2tdK+At3koVY9HvwJgpbRK89NfTaanubTluU/T3LopRkyPjNom3br55GG
8PEnYBm0ApFJEHFTfvI6rIJgKnx9tBKMfqL5mfPxiG+JHtDK37gAbPeoYHa4fs1U
DuYl/BeDNGByO/Sv/IxZh1tP12oWU4azuqWTGZBrECP115sHAz81hJta/NYw+b3E
pc7nJRDf3befXRMsedd8VHA+BMR4wd9JfjJpgzTkdbx/Ph51bVrNuROSM+2/UrK9
3uk8FffvB0D2ObLwD8/r3Yj0wPHKmsei0QSe9/ENF9EDkIVLISFsySFeOFznGxvF
dX5zbQaQMpDsm8elJwQ8E38goE4SUPIt8ad2ePmytn6cGc2lehhN3Q3/1D0danWt
vImjzzOohaw6Qi0O4dPlcOF+eDnP/vyQd2wfKoE/NHLkej3Bgvl+XI5V9nLj56XH
JSZQPB/dqkXYBaIOlU1RUYQythu1BJxFPPRSfH/n8FyK8qrINd8FBdZeNIxbGpk1
9ResAmh4lJw7BkZGk/ziphEDxTej8ZVAanca3xb0ieNQ+WkFUnvr7uFYyZx6/qn+
kzevwbXmMDFgK4x7JfaQVsCbu+GtrOdACBokcQb2R+xH5ljDGlYXL96j+OoLBawe
+9hgs32hV8FUzjCcagVeFlcdo32NeG86Ws2rLYFXcit5jpWfemhW+RSzBzDHiW4m
ISR/C+NrspU1I2gzQUn7d1e5/yjjhbxGjzH8H69flLlefBuctgy8/yENzxgINEMR
gupCnkYaeDQuTJ65xyCTZkQIbuLaJVOvNjhBqVjJxiggROcSfcvWV0Hi8CMyj9DK
Z47+kVUlE7zlaxv337HHCmeqir8ds+5XO5SQUIyNZjLZaiwYsZSDmMWQO+3RrXDp
mcE/vm9QWSUuE0bKAykw6YuxjRceu5MddI+46n5GWK/7DfNPknMww+PK2BVW6Xp0
O4WaMhWEaHSSdJxYcG35FVTR1HlGRFY0mBxYI7vPwE/KwGegFwjJi2zRQsrMKHmc
cNLX8q9prgoftyuygoQqFqrNkmvROUn7LM2oqtfgaCK25cgPnwIlCrJXxojyhevO
zTcLess8nwqXivons5p+zDExE4xWPre//T9rPAAs5mLS9NHpRxoLV0xPZQHCQAu7
oAJ7jHMu4E+rTqAKBFc3cTN8WKLkWeVGkjo7+mQUdnTc6tp0cnpHVOy16PEqmuCN
3cNZqxHQRu6TMkp7+4nBRwSjmOzp3HRQ/KdSnahFo0rJnTYKmGmUQOwdrfrTgKmG
N7VdSkdqVnR5KYZGAFRJLxMFkHQcw3AhfDXMHf7Evt/9nRz1SAFGucz6rEWWyLxk
u1pOGcsyNW2YuXYUZNr5SPXO5TFkC+98CVaGq50HyF+quuaHxp8CDmBgd67Xjguu
w1xV3PQCaAyW0Qpd8udVRtRTyPZXSZR6109UtBLa+7vSwpC1Yncwccaf4KqMPW+X
OJunuJbm14CYvMIo+nkYovEiqR48BguN5/m06qt29t++kipwO6SKUa5ucrwSEv67
OurAXzYdxU0gREe4Vqxv42kY7fN2Zm15zIqIYnlR6QvcHu9UrBUTruRMwvuTe8kL
1bOBuiQmzkcOTuxQDfzlE6Zpa5TeTK+up41IdS2VUJb2F9ullJFefln21ny/U/R1
5F6p5TErCn5racN3rvgF28H2h/ONtrMhub+Db7g6sTYRxCmuLsyxKS+Qwv6vww70
RQTDTjok88PJjYbcQ8BR1ZAEHMDfYmZqq/gFy1Jd//L5yQ841+UWklOngZ2f7s1o
boUnkfLDmYH8SxczwDJXEMUYMvPGHsgzdRC4eoxF4viRO/T7Eh0zf6Oileavzvnp
5qesZ7fvJz8nkJfvf5gzudF0SX6eyO7Ij8amNHpwuZ7WZ+UDixbsg/NYgw8EaHvS
u2zu8iTxPVPUuTo0trePIso7FKYWFh029yXox2GPcmtv4yIWRpZDAKP/iIMG9xdY
DbVN9hqDXQfxX3iz25cmMPEi3CuaSbzUcRx03Ncrkvzd+s/NOCIplz+v4Fo/d//2
ZaHBqhMhc6iiwcZMRnYoS3fIL0glWbeMqrFl1fbDkhyxugidvRC/KBlq89vNBLu0
xtjQnOQvHA4s+RJ/78E6gM+3uc1mH+uuJX+4LYmOucd6UHWrcup20lnjHIsCJ4Nd
4R4SmJymKs5gYCzWsfm2bB5vDucrE1A4hAPHXcSbT9U5Ymf9i/lj6PtbyO/I4+xN
IfLWyEh7Z06SuQOuwwR2n9h5P/qmGLklu5PuT2usXEf6xFguTEyQvl7JrrkD05ab
lOehVEUfJZehVHnJDIw8pAsqObcq+DcPiN1u08plvbsCIawV8cXeCBIVCr70ZGf4
YjMLsbraPIVIOUxnmh43Lkb4LWu27D6PpRYz7wgcvVZ3s3efiUStevf25eFsms+z
mhVVj3eWwq6zM+e9jUwyK4cY69D7okM0NP0D3ddKbZ+QczKqr3v0Thw1Ve+VXzNU
r5viAEI4KRUr2CubBmSkWS4hQ0+/299QDc3MLsbP6Zc3uO2NZ1tIO6FqhAjJUWOZ
3bPK8nA3Y7MItyWlcCPzIFQ7mvJrOZNjJy1x6O1AI1/nszIiGFKxitI6JZb8JoYt
sfgXhyHD93RwOqaJARnGGDii61PwU/49IvYm6etoAZHruQFLqV4U3BYm3u3oCRJt
LdoJlcUJl+qlJ05XyYLENKNWhtXjlMSXj4jv5p73QcsTEitIE0L7nXg7U8yPSB8t
2s0GL0rjS1jmrgDRHBRgINlmqbQD9RsW+Qd6o2a9rVxpweBM8gOHzq8f/1rvTqrG
TSjh0IQs3dr0qvk94YSanBs/SAy+/RsY1r99ofexgrdhD9sSuPiPgn9tlWOftZxA
BThygMqdlACwfax/ODxD8ZIHoXqc3+BQVajWkT9CNFz3hXiMqAytKkfhCyZXVfLO
fei7SgPpYIQZzZhU9V6W7FzQtWLcmJobTYIqDNmnxTPZGNbO/UJVkTjET3pYKjA+
Oh9bRtfFNuc2L4MV74mOYkPyN4LS9+XHCfuBMDasv0JRUptzwfvAiwvXX+YwMh+6
3KqdA2dS33dAY4iMgjxKQ5W6tqSLqu1cMA/LOlJHn0UIfeQBf5V8F48/npLJ9wEw
gLM54nvFCOqglbWOYDOFSJ4wHz1Nf5bolti2QURGmZNFTYj3pfHW2INhOIhSQDSM
OygQiHu6poTS8ioBe4V/VUydUg3NBfMBHfWP2ZOaMvWOxUyr2ylGspX3dcQOiAOB
0hJJd5A3XwFcFZqp7cmqkm8QlQ5K4s4b5nls6zgv8nmBjtM95glwks8tihxJZ29j
kCC45BmMsWTzgpxIj0SUMbaqPnrRGCvP6mEFZyqBhvUW/WNBPQA6ySHkp+IKuOYz
yxXRNVdDYhzaJpu6O4dYCxUFVe9o2Exm9chulMRh4tL5bnQJT4h3FUU+sPD70hKj
9JXJZU3JmAi17m92UeKPQ+hFjZnnisAaZg2uHl7K/xL8GCNyOWvGZl0IImyxxr74
yL6ZmRH4/4euizva6qXt2shJLvRQ3NR38jwec7/6/4LPTNi0vWDwf44UGkBNiEZf
7ICUsL4p+pyHM0K6R0m4YhpPtOy1ZTf3FfYY4UE/k98/vEbWG5KEGlIPZix39bLa
DnLw47qTcEhPxM2JRojLXvZldfGsW8DbeWBMSl5CyBKr52DgjD4M1u1Qns0V1ack
gzjW4E8yQs3/fMNo4n0G8Xdfu9QIp07YiVOrKYutubnkOlPf5cm4J8dywPRaefXw
qBALymFtfRg6lybM2puyBCFJ8wdynG4fo4f/vVXHoBelf2VMBA8j3PvupBxCzQkg
eeyjwAPykWV9eK5NNJdeKqR+7mVMSzf283ef4WqGEO55ZaRrq5IJYe+XBrtKgo6U
8yuYiMWfKaE+u0e0ZTaTmnPUu7p2JtaMOG9shKY/31CmYIxvl7Iu8FEhDBUD0QPf
5aG1Z4vfLvCzhdFJ89FLbrnLwzn1CUZAnjbtN82jgGUGdn9rKkV0LE20AQf/sWiE
EiqEDNIy41sZxVxHMuaj96kZSttBSGA/stHy6gQxXDhNlTOLb5ODQG+0NPV81B87
fnIxmTdXqCbIAVJzDIUCozl04tH2ODm9AS43VKW/xbJFhcJ+jF+K6ihPFKNXhQvX
WOKVOtvwZ68ElN5Gmei/FRVCVshxdUkfMCu4nLONZg0WDLxCBX+yP2hNfhBMElwM
O+B63ZhC2pGCu+oOL8QddiUJbcryR0MLk7yaEHQLavJozFVwGl65kZftC6ItDeKF
gjf2i1k/DQrVxu+el41rftUk/7SPzzOSUmK5LpJxVOeCiONw0l/rYZneeXp0QvZi
WoNHsP6NlytXcoRLdOA0pkHIGgIJnMNP5TTWpOYNy4a56pN4Gp4jYB2G9GVznjnM
af0YAGXd2gkuAaiKThghfWAJgoC2K570WdQ72SDWNVL/lRGGFBN9d2f/SGZkjo9y
OPwmQz1/9meyRcP8qPqRsE3QpEjjmaR9npTY+gTnuxnbv7tS7JM/2XJxju9zfedF
vZMQzPbRUrmpwXSTl0+N+KupMShm10ks2mfK79TwEpFK/SMuyWAskMGvgYahivI+
9TSrPyWKkK5hrpXyrcvTt+ScuXh/u6uClE1WuiwT78xmitFG2LxsNO7ZcCCl17AM
fRHK4DEiVsS+UMrOJrxlCXlwSnSZP8RGce0DbIGHEKOknIrUc9+1jXH4yurha0HO
UFO3cXE0xN/0RUMSWGsrowd4tQknh24prwOSqkhOghcvxhJrDxBmHbv8EFyMxKtN
YtEKtJxmRr4TFsre/ILxSfZNppXNZrvlkWZpwSLUcZSmE/m0Xc5VX4E48LCYOipC
FSc3d/+js5UvDE8BGXbKeSIzwMEfQtsE//q5jeHTPBVtBuRIVUz+ZlFyVHQu1+T1
DybTUJxQ5Fm0TDnfm8OXEAGNkHM9wib3elI2H5FacWxJLtx2zi08DPEKT6uE6KRN
m2FYC+JO3AN2Dt37KD3qiLS6t04KRLjv8MOi0XYxL+VIQhP6RmWBBj7cX1XRWNPG
/kZrxeBbZMZuxbsW7x2zxsq7SneXuSbnKRn1Wl6ETFl/4RHjDW37LYoXT82xaUNO
DatKxsfENtiparN6S42ai8042t2ub0QBymxb/f0Njn4JkYQ6wF1o0BtsPAzW4BHO
dSoiw9AZmVGCWE1QAGGkpyZERpYU2wCLovCQox9U6KH4qTfbVN1BpqI4lrGJRs/m
8ju5JOnnInGP8S1+s0gOlbHQ7fvzg63vIfN7ep4VNUH2cLyl0ECLlVYBnaUrb8uS
2bwfA3xzyqfk5QJawdP+8hSP5OsB2Cx/TXg/uOeD24/qd+G69PJyrEns3TDEfhH1
1k5hD6ArIXP8H68Jfa5MRA+JEwt5PsiwZhZCxr/FHTY4UbzkxHcZ/wzo76thpEb1
VB2O0OSeG2xOhSp7SGF7CK3hn6R15hTtpVqmFtuhhDivOec7sSMguiG4dyRjX6cT
pcRx+rmBwBedJFspt6dC8Ofc+wgm307xGHgq6DnmpdBc+c+0n+7c8dqTWGMVCO3p
Y9Rc5exE77+Xq1jpU+CuWfGz5VoFFIzab7pfsA74rTX4/CEBU5gL95/XAvrTpXU4
SoFSHad/375z3Q295ReuydWc6CGmCxt5XyrrdYglHMj+UoeVtrCAB3407sr2tdRk
zY9PyZaycsYlwJsooJXOpsQdyrgxB2pWE8UCUMWEU6qHLucRIcAaanRNMspVVJCb
/Wjy3nHDl59Y1yjxlVINSAvzSxzVimpUyLmyoKJeEHxB6N1Eyw/MBmlEtc63tBXZ
xGRt/1Ir89F/+O2wxboZJsEksCLJAlKcNf2amQdtVjNViXpiyQTck24rgKIXc0hZ
We+jG5es94e/WzSxr82Mj3NcXP6zJ4tpuI69E7fZb9x7a/RTiJlEA9lky9I1iNyv
MD7hVMDFGi2ukv3iKqMarGfZpxkIRIThIWhZO5kWd8PUqn9MMKn0Uvmaw0w3RMdL
uE4trPtFLHLlAeiNhC6xAOZKq6e88ZlEOE/XuGPL750UPkMvBfJFgzci/+q8PyTm
RBe1tSbQLNDzo9Zts6ewroQtAbADOQkDnguWXFKklW2O31JsrR/bTiD71WdfL1mH
YuFDT3tx0SY/HNGzjoH6/EHafy2iZjARzQoFHmfvhVvrSd+kn5tCgxNxQG6nJvMW
8KwQ7/ZQvwFgP8XeaMrj6YZ2gcK880ds5s3KWQA+MSACfhlGMWVNo21WKxfPWGg2
8ixjLuZhCgXRNKviHDobalrWZfWDCDR2FOoca10vImJsRi044gRvSCDGCAh9tXjP
gQhQUITNHRqJ3syo5QC7La866gLCAIw0pkrXVFokjr0MFH/pTdaJgwYaafaBAmbw
mm3KVQZ7EPfpaf0fYWUKMjIOhXJlUjKDfc9eK6wlKFQB3Z53uDRufLQHpxjRA+Eo
0rhsQKO+7ykyeCHy5BHL387r5D3XWx8v6160jUrJo5Pfi7kQ7iCIrXniivqxkakv
MRqUDhn3L4fSHApV+QDEfWolLA6m2hctf0LVLwsdCG1zVNHDENGAXFU0cdu0WUH8
VzYWgPnOs31iLc0dpmKWvt1+lC72B6dcfKEExNZvkg6mdZxy3mbmzzP/clPFzlz9
jCUUovTyshlOoV/YB7MTemiLV5iy38TEsrd+QrTCo9yszakiwJsYXXtELfEBQkHy
JsbThS0Em2C5S9qwgQk61x+uLv+Ux+FkxNBR1RjzOMUbartQitmCTgAYoH7tZEIw
Npe0APJd4H1ZjTjCvHJOU45Of0rLrk7aoqxee0Z3TkH95SebWVqKMCoL6qEySfNs
7TvX8pLF2oR/weUJkN6aPfditR88uOrP6mnJ3z1ADDYNFvNikmtZMDK5r2/2KOyP
mLfV6S6sxa9TXoGY05C/CqiQXsuh01h62AI+6THJrZQeb7s0VtbfX3xFhQ3b3sMw
61PP+UCaryf7q3gmeKS4Y+VnoGVafoIf5biho1Gzmfwmok0RxuNaYPVBXryxzMhF
dDrQrS2ILXMK1QYgwbq7hJ7bs5vf59mew+1ZusHe+3+aKEYYuLGWoj26zKOicVOc
jD0Gm6j33glHYwODvmEzRCw+OAe1TQXVQl4ZMtRSpUIL1nVUxcsAq/GxqPAPVfDv
5LfukR4/NTYDLUVhznyCPE2GsRpT26Uto412arlhGhJVaGM1HKHY8J6BgUY70VEr
hRiDG8QSP99TgF5y1DK44ftUI2D5mhs4eagp4Ys2E6c3LyTwou7kAM8H6us6v38z
KdsTz728nw3bUwg48DZ/frYjje9yZ4CPCMEHJVNTNIXZE+LLsm/fCfD/WIMLk6q5
tnV85hOs76CcSFIoNdn/nq6NvWTX0DXmoZJUVNcd7pRq8U6+pEXgrDJBJDsMz8v+
Ma/qgHtRQCZsaCvExvGuIwQ40srvKQEcOY4QBVc13OPh9vi/jqkSpCh9wYou5EA1
DskK/egSdJUKeiNUU//JT+ectEef2wnI3VIhBr/oUM4ydbsjR2CaTAufNaDdOkCe
gZaadAHrqN6wEshRtWxPdmLqpJbC2OxA//KTUYWwnndxpg5TPECPUNguIY++K0SC
gkm9gsvefqcKvhfbO4sEA7f65AJ1gYZs9gOXBqJpufxZEP6SYxSihyJbljTzsZLm
0+i7oqcNOZZyywUVCMCm1eXAgTL7UZ2Tgtwt0ZPVv9LSgQUlH3KWW7DJ9NL4Dyyl
lFbWNjJrvIfGm8tmkWOFVmFivaUC6z8YqUFUzQSw00YC+dLGjp7XI9+XQf87jQFq
ZHIYZumDHK2AvMaGmGQiJzn+/fBYpoNF0NpUYVRbYKuI3Q/7kUX54QI/g76DQBha
3CLLYrtt1psaJhZ/P4jQMl9RL62YCcJwuyBB8PujZDSrQK4mTUYS1qvbelKy+VNE
ZcKqgZTHFKMxWDmN9pUPlQI1B/pjxBCPQJ7yP3mOHjG6AcPrfOfgtl5P8Y4Dz4QU
hVkg2wvn/jCp9R9/xr6wprmPV7rQSlF4bHX7R6355w6a8s5hahr1EIxbVaEXTxuq
oKJpAAcfmHkr96Tf+/+gZ+gf4KnJvRqwhEjoGg8gyAi6Awp/+LL8lXmr5iqImrSj
wqlujpWjQL5J0BkA5xz1YLzBsTFTcaZN0TgTUkrJUfUG4afUxBb9sXEG9hMPXEYI
usavA48nXBV0mFr45k/Mtp1KWzCh3dmxwL2Uwc4oEwx+YzHe0h9LDENSPVRfxoZH
XFsc50VlSOtlv6Nxijm+cMnT+3fOR54f1RvEc8aaloKc1CeADWSrA5t1UtECw4ku
ngL3oTunKelWkZGbkseUPlTGKeOixLmj4wnBbI6rLRe6JQstbYJKOybVwbAtfF5O
BXyRa/bWN4AJuX3uyjZWV6E+k5HGchqGdRg7idM3SVW9t7e6za1EEdinGR5L3EHF
EWtLcE8woZQkGPg1NgAi8VlrMIkfB7Ib+CrqVBMy+gZrhlBEGYcJQMz4ZnASy3JU
6E9UezOcAQrT4O2iWRX2xXkUO4lBk+1pbxp0gaHWs/gqwcwYy/cqoWwD3ekPDvdi
3IIFwp4xNCcLNtxO2/Sy+3X5hk6nJPr8JXtPN2OPh9KoJOacrFpnN40gnDp2ESeJ
MAMY7PK0I2QDfWwmArJfgo0JkbCqIwEBCD0hrJMhAg/UqUwWkY1TcoGc+Pu74y5q
cEOZm2Ud/Egovc1I4/ygv71mfROL750Zp3c7oBkVb/DSUsG+1XelmrdIQKkKyK6/
SKYmn1HPMpe1ur6Q5oOHdr4yIQc5A1DKeUt8MX3eBp5PGVrimF8oLVm6Xzfcn77/
6YiZb/Oa14Ux/2R/lpVmw1tkcicmFt6ypmbl47G/yfwlPJEDLhLkhKQD5x4fMa0O
Qw9v9m9hk8IzVNjrksnsORG+MIENKXy+11mWKTbXWihWfAlr5Qu0x9hLwzjbEOE5
Szk3newGSm4CbNUhe11HigRYweqAJLbtcBuyz/SrKDWKNBoqHKLf3cylpDQZjZeE
0fKOK/UrWoUHLuRYdXQw4cQYLIoCvTh6qhZr/fwRVCWTtUL+9ZbrSLIRk4cfHVgK
i8JLkL8s40eysr2lNagD47R8NmbAUuCcbZa9s99A51Zc0efJZ5G6GW/MMWQ9DxGG
fCfcvqeIg0TloVUHStESS2/TXiBlg7C93ubd2TW4JmYdeCNVMet0r+m63oTBuJMT
MNeXDIYT1HarxcLpgT/vh27E7KCkxEvNXkhj+lWxMuck36l42RXP3E7hAkTFLLvh
Y5gDsyfV5/QK1A87M6iSaMBOQSVrc9mYJCqxmndC+zsXXjUCKfkV37S8zmGQOyRx
6+SlH0dZLke8QsnED/57eAYNUhQeUqtnZFYKQQBAktlO5qUXvd93wz75vEp1EV48
AOFlZpsfHmusTISPjjEQ66WSEAQA08BtsMgdcl8MqnbQDwnHoEPs/AcT1/FD5Hh8
9bzlRmPc5nfQNC3r5hN+KlIH4T3AITF4oqLht1Xb2icchbjjD9Ie+KD1hu8evCRz
CmD1LD3FF0oWOTPTm48qye9ZOg2v943Hk0uyP7ne1HVvqZ3oOr3XGPlhXNQOKqbD
cd/l+M5mqyxHLRpvtzkzZ/KWPUw1rCidX8hzRDuzvF2+CSeueHDp7orUO/ygtDhu
N0dBtCcxYNlfXPbqYAUU1dCH/4QRd0u+JleLCC7tbiSGks4xI/YGjnIleTh9+kb7
d7Jl4iHNES52ARI5okmjum/7jh8wciSr55/GxG+DE/HGphNMfPXpzY/mYi/Jxf76
GQfSc1+w1D6WEou2MeVfK4y1907OR1A7nrLIVtYRCL8bNiqTc4tyXIpmSeNONnaW
zxoJNmS5mF2F7bzVcnidAATDH4beokEo6VngmLI7qQyeHrOfCchIDpY0y7MvPsKV
OHV+AuCvvXe7cdSlxF/2xAdqioVidPdecSnDh0Bko77ZeKCh60ksMuvqXb8azLOR
VDhUbcYYkphjL+a/DOg6WDniJ+l9fnfs5CJFOG5LvaisrQov7jmEidhuJF/C6i2f
0IcFeqVDIIOON64pagoDKC8AF/27zh7WddnoMQoQUCThSiD/GML1R/PKckiRxaj3
Tuz0RKHDWjLqL2OUDs4Ic5Tmb892mC/KBpD4vB2qrs8m8GmVCgyJRNH0Z8s40Z5D
wph6zVQTRhH3wbRqT0qfsDGNWsVUHZJCDVyEnv4g4EcL8bi43tKmhy7b2wq6UgKa
lsEKK4kMvNcpWpM4JqCi7bW+M9/HAW7FHxX5UjWncKzojzb4mN2SRYvdJCNtpPCT
aUh+mD95yXkonA/aeP03R5oGXJ4gtOJd+DLKeQaCI9sIVIZHxEbRp5Wi7ran4QLx
hJpkOPUdC1G1zVYyvnZw/wO++phgrzYROsUigeNmwme2sEkh4LmSyCMap/IZbpIe
NdPYm35CdGWJEwyzxwgf+pv9vW/f4gjHVl1KYrkGly7tmMejmTzA/hOQdTQ3XUD9
YA6TYsH62R+zjDhRzQqAUBH5k96GhEH4a7Q/t5RY5+k4QMmzQhikvmlMf+YZF1QZ
eOH2mFGwIxu0ibCmyNVyIl91yHit/MGCf/WolZiXBdyFOR2x0+xqSpsOR705agkv
BzHxc+4412U+z5Kn0IsQzrpyiqwMY5JGTxz4DH/SkAP/vRrHATdwIN+t8lK/87tX
I9ZINgHWTXN/+PIBLDLqpE0DrUh66T4gbuzxYCdW8FNCeS2lhJBh6+fI9TwjLgK0
uCDfNwQwIsaZXSWrcE1Kzr7HG+tQMU3ZnIEDeKqbTiMIqpGeF69kQUSGW/3tXqCW
XRa6WIlLES87OaAezmv9iWPeua1E5Z988k9WuNBhE3ufLwRbAksa/MNZKwLcbkFd
KQ1wNIv+Tai71sH4Zz0gQyHmDx+3qydGjdOTb5KuOtSOm5hnpB1soiPKuffZ32vP
IvKWR3/FKo1i8ntiaolLoSd9SDEorA//oVvI4qpqAfoN93Cd4tlJu/Qc+I3/8qzw
4LBNeevW2eLjJ2YOqiAktUempdA0fmpsoN1rmbSBvdl5CM+6nUUFYhGCC6eGWkdS
TI2ZPAMXZtxYgajbFjgFwFPgZSNzZaehmV9ipLuug9Drbkv9u5mLEjLFXKl8qYK1
9mV3E3ToPSNkdmnkBWednJE+cdc6s4gTNzwm0J9B+JhzkdqzR8AL2qZATc+QxkT7
Dm6pxpRyeUK8446KcPr1tsRh+Nl95HHXdBZTjzdkT9XhT3hZvpQ96z4m2N+6JZax
JNoJjmVnJnH0qCnL9PqrlCH97T/KfkD2FHdlEAwDycLsNb9MUQsnT6XDWYJPFZ3Y
iqf83WNn3RS0p632ka7bKOnp5Ko+OpKDgJVBirDuyeihwWPg4SAm1utiSnpe1pYy
k5hAhNVlMXzkLlJgf4ztmEX8MHmcq09t1BGu0eZxmH8Its18C9eZF13BJGAt/Pb0
KemG08oWY7PQdIlESbEtcpm58trv4NejFT+m2kCPxeki7+YpkA8HRvw1/xsdKcSK
Bx4YNAailb2sYGuGV9aptdl3cfRGQ7Ze2Oi5QTe8Vh/DPrvGzJ3hVT/5fioDYGON
e3/vfifTQTown8xt6jEzNvKZlUUL0y13XiOtP9fPwwPphorHwiu5bfc/Q0h9nW/h
FVj5/SvfHXV3w1wli8wFcB37yn1s6Lkiqq+2ht3enIdeiFVb3015pMDLyAvqiWie
OyhUc+XjQfcQA+J3JLZ/wUFcgEE4FRWxGl9o6/NSRKP1OqvtOUTLMy5aNryhZtIV
3Ve9E2BhY1a/Jj1BMQECrFZU6MxlF+O3VV9CKv0JcWPEmP5SeIqUfrNjxPQ+/chq
Jg7dZS6IHFjKmgHM6LsDogmsKLa5G5uoPmnwQl5/AuK1cspev02Olqp/xWcHKm7c
6oM0uDmOwrwGMgd9ABOm1C9HW7SbFu/S3fElhy8sl8mPzJulDuF//g9kwFahGUCx
p46GEu8dWfnVzEkYwOEDtRRC8I1y6dzkr7TN80XjMlfYgUX4APrItA5sCrnnSIKq
Kv9S5FdWBQDXpCF7MapUImrXQdrP3w+h4rRJojDbeDPp1Jno8vnBlOm8KCOSxp1I
qfRts7CvyDNBwsSKiVLnHfPphYlYK1qRpM6Kijl5ozlt8z5KnbJOrZ5m+9egoDXd
t80dMy/+S6POaPkszI2FD/Q0kDoGLeGwJTZhPImqcJ6xYITheBACYWEd4dXAbc88
GG+hBoijgJ1If+87Pbse0PfBeSjG2Rg5srIGt4Xm5bB1xEKKt6caOVjRQH0RLlX0
Z4jGQniWwRjmh1tV3KlsbJip4qaW1iWyI2sE+hEWELdNl/N5FJxo/o89wtF/Q2Fz
wJVyyjiK3m2AD7LBLxd2mcHZuZTi5oeOrRbPCSjtibFP4IQKbmpxRJc1Qh2iGMHq
At/00OFDstK/rvBhJtDgLtzAKvTAG3Qb04FWgGIGM4fpKzSy/+PAOX0WYr+qazWo
3McOVPAbwl4uFKwccrslyi3LvkXVRCVCd3kO+dIyTGHRx5JaHy9k56SwhKVQIOal
yZSc8bzhC+rcqLg6I6L3yu+9iIqo7SIK/aZqUmL5ucDitt8d4yoziat8PaXGplZU
TcDRGOrCzwXTQEu3OClfddvNCrRFdAh5+knP1UBS5GO1iBk0yO5F/MjTbGemPtgN
EFL2ifwS/zoD2EP8FCNs0ypLv5zSMpcq7DYBpcWxGCkrjl+MZvRQX1NpRCpbXEl1
DXcFPIdOTr7JOHvYkCNxpscW+/ML5mr258JcaUWBkFTKgrkyMpGKv5m+IXOQZzOo
xqLv5eJKQhncjASa7zc85NJBwYCDSoUSJqohmGMm1wxoxLVmBXyoDnULJeH9vLLZ
1pzMPiafJ+xjW5Hur5rVTvkarvPEEVYflx/gKbVHziizGbyRk9RKuYBdNEE8FVSc
hczPSZlwUzU5rkOHJ3FoV4b7eZ7MpU82BsMSxSLtoRPzVggoTQS6b2u/iwvk97UO
nOAirMGsGtU8MKdK1vpBfYUIdKcRQZisvTjWh/rmd2GvW4tVQWEUXOuXbR2XyIDq
iONqBshJjfRAAuPPpSYatYNoMBXm6ksTYxFHXqMJS05As5Dm5ipU5gywAOhh1DZ+
gd0difLNHRG5W93xPv+gOvvPdFLUiM8v9BeiGmJAwpY6+sSrnSuBs3F3BAzQcqi6
uq4MayImCKA2Ap0rAIhAvGq+sCrhriQ0mBRj3yJt48CqZEy/1Pbv0asu47elFaC6
ObX3Veo4j5h90z+S+Zog0665FZvSBBvj6PgtAhj9A0rqm90HM7VbvmZ/InXIu6Uu
RDORmUW3Erg1pvwvv+jlavqvIcbZd2u+l8PrrdXaZQwFZ86SM9ONJZSqjWwNyH5m
m7HT2mHcFGiME6o0vO/q6JDlCq+hLhbEBMkjJ7u5FUKY8pMJjRXvArasxbhCJNV6
B8Lu/2jDwOQQIERd/qfS6iGvcTkzILP4YR3JbVYRegAU+RP4Ihb7DrPlESH+N04a
FckKVOVeISztRJDcq97ZZM2a3jmb5uz0/A/zjFaVGR/51ABYzT2iHI22G6YGJ+fg
kvsTc9dZrDdQkL72+ZZEjKFizYVB77XTQVYiSPsRG+T8ITzfr4pBdVPFmKgfpac1
VYh1slTzwvQl9MUIIIv0GuHJtKMH5oxt+Kg/c3ItY+JgugMO4o1RzCqKQNjQ2c1Q
qa9vUpz31YAtIVAI34VE6GQkQtbbkq9vH4SuCVOYQqzDg1a8Nue7Y8hqBpznrHfu
wsL8oFRYANoqrZqf/ETIAwjsHY7+z2yEPWM7fGqanZDAGdLwEKtco5NTRQrsT/SF
xBHoiTemiHjknIOBu/R+Y/ZsrynCfqRLKfO25xUFQHvtk+NYJzdSPEu6m9EObYMo
Rd/1WP7d7ZinQ+qa48qgDvTCQsE4ZWFMr1lD+tHmu0YH/kjj8TwXLknJXLuJIXGS
wW3xK1OoBkegLCfWrNb9kZcpwmPgKP3esKgsc/TKX7cqkKfWdkDdEzuRlU72/13L
HQN8oven1fmaf5xyCUYNJ5gqx7xdwHnyYbZ13s4anpl9CqucnLeaS0fssEPTwFdp
I9bjn0hAi/1IbPd4UZZFvcVjY5YKbUDEf+bajFiHVN3DjrhWynZ+65KRelnzO9EE
MZJOFDlIdEtGRAM+E/UJWq6joonuSbW9OVpBcKsra5xLoWQBEM0gVvfS7leZ44/i
ReLusJ/wDpP+BvO7UCGi1JwlwzhO5A5bLF+BJnxw4uMMdyqau7kq4d3Id0EJnH00
YPKvxJSiVQjFk4pvFotNQTSnfTJvMZGOslo3JVOnlmqCVPaYvOhJJ8HPsLhLexnP
AwMzgVEpPWHv0o/e8r/MH1l6d5jrxmGkyKlPX08X/Ru16URherMel/cSgRUj1UDY
eBQ3y47K3oGfTla+f/C6Fy0N5iTYuBks6y4AS7rZfCar6SD+JV6tdRdKj3WTcamX
ePg582hdlf6ewXw95EcSJjtIqP7WF6dBjMhiczWMi0EiPC0oS7zJ4i+LhseAh17r
h5Unj91/WVULB9vCHn+kS2qLrsow5nH8Rs/ZlJd0LObo6KsUPi/A7osSdRjEFdCH
0O55fGjYlQoMd4p0FYbWC3IhR0UfTHVeK+ERiAv18Hs8XSqzI8i31fzhAGDr412k
ePVVP//z05i+LW4/2FxEyWwUyW9wuCICltT2j5N/ByzW5vfaDtu7v0B6DooAMHeH
lxJGOXddz8zSweH1yXVOiFr6Obg9X1G2gyNAlXyHiTLgwCoN40asnaPnrfOIOE4p
mJ1/pDjz3o15os5544KOElJ+Q2nNj+QOUkfJNyRViWmsgIJzOnRt7TsTcGkM6cUf
cDCIZ2iApzwLVrYxv5iiUy3MPvBhK9W9svZN/Vxp27kTQbNGixb9wL+HFIFdw+0J
d86jlPpr2i+8NbAbcjV+5WQ+ENT2v14KWY17zYILBWOrWzrWizXAr1JcfXX0hbqf
gl9EiVeAh+PdupI5AKTPMsdnLLb2HgcLfTZ3kg89H9XdVto/lv5VSMZWc3k/SQ62
S6ItYI15XQ89ofVHD7pqh6F4pvCvo300SiOw+y4FzVXFXlnDfGtY47Vu8IUwl4f8
Tqk6R2nM9086J17rbVyS4v0ME2Cji3nEMUfVuBqST+SFkyh6MGZ5ztxh5SMJSmav
NPxPXcUslF7GOyBgnkUhauB6Z0pmdwuRIVU+/jHMm+q10eXwtaa5gStRIeFdwAUv
fOY9t/OWau3S98jxbAsBcvXC64mwku/Qbkp8+ekX+5AyaX9wF9EctRMq7kNJzDA8
LRmNAPpMdBBePX2rJpTaNm3+xOTEiyo5XpsekKKZ7h0kat79kMo+BJcWM3jmI8f9
kBKMot6AbYcbiQpqX8whQwC0PQ5hcrFbw0fbLe8d18exe25gGEiELmmv2NpDvx4L
HXZg2O+EMlFx7/2uuRmaneT79JsaGm9E+iEbKSXGO4hpq/qW2hOHVT7B+WemhN4a
sJ+p7FtyM9d2IJ1vuID93IX8cw9X30v/lpyj0Gim1qJKoL3df2U597kN2xaAftkT
UCtOXfxzYmn5QiaRxrRg2HbQ6CQIA6K/KRYTuscDE78x5mv/+KnQOTrQuQgiJUaQ
tQeXmBshxcZB2fdby8hGjpRLMONmhR6UQVwMoqzGOEAJ4PMkidxeaVQzfiHUJxpV
3zEw6/xPP7rnMHIql8vI/4eK237itCa+mspMICzC63IeLiuUQbZqNbfK0q100zTv
IuxMzMJzDast9NFUvzdFypSX3S7UTS5yRRRQVjtFJq9GFfqmlTsbPT02qvi9NYr6
/DXql0RLoHSG9zR+vLqFjPVwjtKFDwLi91yE5ldnS4X0rlpbdUisvej/HxLXRdqO
lWYbpB87gzvzz7e8apwXDjLu/qMXfUVaWzj4vVzjNXC0dOE1JzeUxVX1FZgPHHEg
bkmi06qVYaQ6uJwfxA9E1nTCKW4P7itGralzq/FifJ7hqv4sLyfGDbIXD3rnsukq
F0pFCDaF5asgV7S6rQ7PXXHwiYH3McDsC11OyZ0xBGHCPz8OadejQnibZs0BTBUr
9Q9jG6GQdjxMuPN6yJEwfjPmmkR/rULF92hjjkg0F/mk5XM0vfScca4QBx3/oZMY
Qzzli91weA6KWnZO/Ps8MKPP7JZssqIQWBSwa8LlOIUj7reKgCjA5HKFx9XpAMcY
O3qBAUz7xkQ3gDPu9U1w/HLbvL9HmU0p8/fCFR8JAGHgydnR02/ZRYTHNqMVu7Sc
28IjBJ4KC6ADnW2XemV/1Hegnv0epCjHVYSTaEXzbRyfpTbM4SEa0qMUbOPSNvfL
BWGad1nLz6vKW3z+sAjyUzKqdJyJJDIeDc2wojAUl8LS3QJX/nv1s1c3WJP3xGya
0gpdiUzkmG7swCaFw0LVDgoKqFCxEEpgJeQ6UniWhgMmR/XbtRNQ3MTxL13cZPve
K+ceaEMig82ckg1OG5waJ0xLK8potK3jMJsuxWBN7R0+a+3RsJ7YK8DQSbwa4Ofk
Kt6cNsJrx4J0k3f38iYOZJ9oVYgSHf7LqJZlJw3n0JPITa0e8uWaOTuKyc3UCgB/
k4S/rndr6XaL4nfgl3sWJrfbeGWiy6srl/yFdx4UwFsZfESFipNkr194gXGi3PDt
oRc+OKz+KZ8KRvqS+ezB7SJlL9sDSVIHpcpfWN4YcCliteogvAfkrOfYYx3Detna
iM2atTOJqiEzzQErsmBcYs/U8FTWTZZWfoakWjLev/IrjpjQhWYVAjuq7U9N0Nd4
MTF4QRqCWUL4d1GgY4tPGEbxkpbXWMmzdj4Gjch/uaRl4QcvwqdGugKLd/+nw0N0
z/OEasxZzBkeqoXEYm9Xu8l+HyM0H4L/2HM0tt276HMIOxs2IuAhhlggBdgS/ARF
CAOMauFhwRzRxePQ53PjotzhMbDroAK7K3Q2wkr0YrRkb0a455Dd3dEC6VJ0yneh
ZPvQZ3zl5+mi/bVRGbdLroD6O8hJO2fLXjjG+TRzz5mHD9fI5KU0zHZ+dKkuxehX
kB9GhM17wunAii//H2byTxO1wOw1CMH+BAbXfyDPynCTQrOvwaaGgoICBlESn4ao
bxNWzq1LOQpnL1GPxXjF4mITpXw5vKz7vXviHxd5YnNK2l2C9GJfqoqjmZQDjEkm
kIBSdZ8A6FYsPasXumT+AxXtFSNq1qaCYniEKSVfIx2nLk37gFKlNr9EAQ0HeRZP
JBva3Kq6LZdwzw5G0wjvCHaAjPpRHDLItroL9piU7+lQZurhWLYwqSXDc9Iy0CcQ
6jyKHQr+4WfMh2K7sYKTEaHNZwi6LpMEzn44dAxPSCGBjy047GycBd1w+5KxoI9O
2XZs4NxQeqBicxMtTKixXq+DofI336g9NVtn7eGbluD9sV5ipe+t7QSrZER3OMvc
tqCjsjk7X4FjDdZn4xt4fuce32OdxpljTcCtd6cLG0VZl5ozXyor7DeIhDnIy29u
1OMNmQ9WLt31ENyI5l1wyveWo4TgujVt+fZrSbUuK8MaeaFzPtH1clL4cMUmMMyY
OHKzpsnaboYilgnJOqtwZX6PNl8GBG3BBPat4Jd3mpq6z00nkHH7My2tlCraVsvj
oDSs9TziRFZSOjUJRxgfHs4jQGitL6a6p2IezheMAlRVf/FT4xSD5Tm6jACi301e
2LKwYXD+z8iMVOcJzfxCCWMQ8Xt6Cy8eA+7JDWXPJe4VPNSpMs1U6AEjuqQDNzoE
PBcVJFvcPweB9qBtcfzJEdm8HEDkjXEunEoF0Zd0IPr2TttZXVQxTzwqKgHf2/Sz
6UqRBp6xdfm3EojT9ac8ME0uOAmMmdB+aD/mCozijau0ldXZqGfISi2vaEZDCTAh
XCtit4yDZC59hHZ0U/2SVOz83LFWCapQpqIf2Koy3hxR0lWy2WRMKRWhAU4lW4uw
9hzGsBKTD66f2BWrkOGVacvLpVnPSWVaBydzrGdta7S5QUjTWcw4p6SG2lF0y2ux
1cchWzJQg0lKF5ZCOUnX+9yV9DA80MsAyGlIiGPPZ5p+FVDgeBEYdQ0yUkpzKsuf
rXLEJFitg/4F5Eozo8XJd2nJTskGEhMypG01BzZ+a4oWu3pR3/0A9fdiSha7tV85
lzy1rNFsLK98o0WevRo4/KI5PIddGRdzwLIafIp+07auiuQLTyQ84gINcIZBWKoq
s2tbrhKFnIcmJxD3fR5gW4NKDsmFeSy/oVNl2CiBgqvWiDlLuvWE+3bdfDRXkw/e
8zWjgslC8rp+fZwU1meQUhtijVYhRLHL7u06ATJSgg6tG8/4f+BfxLK3x//CcwWb
We+ZiCVVdu3nChRxmVdWtJHYVeqizwIS6Fs35acYSqkuY/PvOhIru7ByPiTPZ+ZW
bi7P9FChJ5DYJQyX1JVCbxhBYbRYMCnGGnl2BuJdAOrJgnhfgOG54Uksjn2Ml2f+
pysqsaTAR6RXhnzZAoSvO5Q/cxnhbYi/KTsxuULK5z3HIJLStoXFT0wz84sEKG//
xD9W8+crmWb48NNOdhDP4Udxew1AH3lmQX7tMfE6wPcvyJjvl12CxXMpEFtp8AnP
McrMGhmDbZkGm2ahQpf9evNQLtrjO1/lvlLs/QEuzaot0fiaaznBq8RfcQimv/Uw
HtDGoAn+VY6q/lXovuggPqXuPZTHX3cDsjR7x+r51jTYdOLjZRgrFjBc1W5so99J
XAPvq4Ei2q5qSTJj0c1OeBGPCLnGf8kh4mqPlULrBbanLbACzNxXOWwkXD782icJ
NakPheUF0+GDsaRHa83BfSXbb2oI/xi8E0f8JKZI3xeOyal4WLCJ9hPsFhVorta/
PJfTBh9AyfWZQJ5H+q8TzYlWcZg3XKrSn/Cbb/TMQAWm6EalaPNr5nUFnEoRYTHz
3Ptd6NLzWcrca7E7M3vN+AeN9/59PqO6nNaWUqOL/hPVBhKeuTnwbL3MwnPWZO4L
SbeX8mphhkzTOgxBYX3jahGP6bK7ax41jytN0IY8Gek26koo0GBipdzyLe/DD7E9
3soxV9bNfHqB+LawVi7H/OoZATBqZ8PzeizwlHJp+SHdlIQ/Jqa+7Gl7AtiXrCew
EOJVFlc40eZueUgpM6668c7yxNf1J8HyhCS6jKsGUiNIq3Qxw9H+6TOAMtMIVOYK
tXICLNmSPXF5OZuHkkWzA9oJi6s4juATfhRYTIHJ2Kl998IF5hIhVc6LUAsHl7DE
ZiZI/PAjClz+2q9+tYO72WIVoCKUnsSTomK6dELU+6Igx/mIh3O5lEmRzfkrmtfv
wDhfIFAMVjKpb1SyFMp3TLD71qvkrRKPY3M0uNXZxkk3EJd+pPNj5mp9jHcQPI+P
70NocyATEtDafvoxzT+iMnAXZuGXvI/965RykItRE+7JOfTv7eaaabIzB68XRzcd
z+mnHGJ+DWGtz3FQ5gCw8SMHAletM+p45Yp+3xPWA24OluqGX1M3KaumMLPPHEo3
OgI0eu8MiZtuKWS/1K9FSNqUclNHRLX9bWZBGVHd5vImq93U72VNf/OIm5w9snFC
XoxmZA9YQuJlite3qIlehFzrbJbvAv53dxmydhFEzwpQF2pSzFnrRRRswpS7HOXw
OqpF9d3qWmIbhuX4iH6oMDCvIOCpdAXkWTlJmgLWxhgO//folieeD9cTamEJ71mA
lr6tC/KNjvjTpEQx9kexjdRvv0kuyUzlsXumjYV7g0HbSvu9k6HbK4OsuMweYQH2
NBrsnuD2EGbg7sbaytz6S+tOfmFFJWOcedc/gD2RwfoJKVUtLV4IlAMk6+sh/Ibo
8kBMGBpVHHOpRFPuFsBQ30VvjOry3OiziVlee1iSsB2Z1+iWF8auga+s1psGjEv3
de7z2jJBS2ylP9/CXIrAD93ivkjwb1HyW0zPuNvbH4JltZWCqFCr75JJ/aCZrs5x
xDRKMBY4RnhMcj4rImUkyPh9xt/cXWV4Rpo0L/xoZKO5AF32AeccZp0IC5/pd6lX
CLEMYuFPwWlJoAMQuE1yiJiXmu0BLO3uNZjdxLcGXaL8q/4wDgs77GAw1IhJ4rbd
sQjKwwU5TgzntT5XG6+a2CuU+e2ObmATVsYWyHUwp2ExjTE31qM0Eh5Z6G99hxOB
8RrbjGq+yVeaEo1eLQflwKnLTiU7+5svUn9Ehd8LBs0FWRcF6kNHZ5bZReAfoe5t
RGj4Exdirp/on9ez065fOcjYOhfhBCgukBa6vW0Kl+AaifGrJgGD/Xx2lz8wQP7m
viPfXJl7Ct0kQpz5feMhVLSI0Ec9D3h3kSn4PxGmCm9XsNi+l7VaEoqOGIBI6G+p
b/9PtRyAkyrV3/MUUW1gftRDZUfHS2sglZ08iY7jpwqpYCF11REuQH7K1CkaZYzu
p3ub23PkJtqEoc0BnuuAB5rs6sJ9qfUM5RKlgzWntgwtzOQ9g6VUXc/dPk35Iism
zTgmaENA2Uss2KWQhVCDLggzzmJB+7krRFlt73O3S6tJ0GhDaiczcKpLbdIy4v4P
0iNybv7vbnU5Afr16q17dw+gW9A9ps87sa0BV17oEL8JSUzaEOoTOk6c/QNpsKRw
QQ910a1lsvs2Fxvw4kDCWZ/IlYwuthTgMpTjIL6ljGrMigWooRWK7lNnVk+qdO0A
yza2nKyeGXcoBD7XSrwJH8+gnp2Fvcjsa6wiYtG/UevnpLzOAcCMczPPYgXsHwkK
oQUDl5tVjcEfx9tQdx/TUTbF7C1j64vlFPiCUHymZPL9tQ43hXGkHHERWRJZS6hy
JrCvc1bBG9ozf8k4SLaVpcouBf+y+MZCMHJZoA/6Tf+fBLvoko/tjTE4TAnOGXGX
JAicS3p5l55dLjcK8Q0o2fKWtl3fRb/roz8YZ+eXawEJ8YaBGVyDS1x3l4yn08qY
ZwMCaVkC6PQzj28fcMM9T5DJYsB32kkHYrN2sz04lBGJIQUpM37n8MtoSHhf7SIW
G09TJlHjDvJVQ3iJI2ZShfqXwyunhTeJew0XDatUtoKrSfTV0jitPF835CdOPmJN
OrFdsDiDed0DKP///jIUvXJ4dBbbTaBn6rpe2ruwrHquzlkHOFC9/z+SF4UDT0wN
h1viLdVlYthFfC8xlZOlIiN2Qz5jZlkIGPO//oUSkmjxIMSSUsoaYKS3FXdaaUUB
GE9ErUHqbFLFWUdm+OZWDEtx8FnRVMfKv2/F3Rp53eZMqVRrSPjuCQobTny6N7hF
4IU1hH/49Uny7PYriRrp6pC5/Pl6px5WFMegt+MGogc2vR60CluKS6puax9VpjdK
7YZb+0HNsu4uabz3KhzM85ZktTbLRmOF/eWT6/4UvQjC3V9OIKJhE58r7+uPOjry
w5g1iBqIpxSNje56h5zf3E8Cg3L2bOkrkYzMFERoRU+HL0T1E+I0flfiWDUeX+ju
mm1YRv6N8df++ZMNEuSI5SglNMcMFVoRZlPg96X+Lfh6NFwffAlR8GkbPvze5DFN
hKWvnhvxrgXK9D3mazoIq7wbXkmVOeMmZJSek9KB8x40dX1yMQuEdby2UlzG/maA
oVlS919H71KSW0lmZcE4b9so7Z05QVIYYwQRfSciAm9q9VKK5QDh0VzBvztvqmTW
ZTkEM6UpJh50RXIO3tdmQFYVo78Q9G71dDuylIsNr/EFXfliZwSOrocWZIEGlV1V
FO19xLi2V+poLeq32n8T9CLzLhkeKhXCUq1dGW5HN0YSVKQ4hhMksFjqLZe6/dht
GIHcaY8vbFbzE+dKvsYPWg2P6oaB/SGBE+Hkz1r+UKPWL+mSTKr3MpicPAntzZJu
7FYx1RmeID07CdgYgsmPlSxFYgtW9mf7AR/9MsKvVzyABTDEuViROn/iagpMZJam
6UBVf6LDab9MKQYEiYYyqiE3QIP/atinaYA3Xcupv7qht9MHncD8NXt1uE2zowEc
elpaxkUVInkddtsev7esMHG4uH1CMEiBZ5U/EjSvt3/sW49YNH42TT5jjbXqzvp9
1Owf2Ef5YeXl4zsSls05Vq3JVgLFYzLx9ULodN6K+UoJXMZOLPUwJWE7Uc3p9JYW
zesawLpKVa+B3Vdy7WUfGe2jAPjjnmS41XVPFmbCX31sDUSsZfxfxrRglrkog6/D
VDY7dR9Z0o03guG757iqg0NdFXLik4H8PW7F8UxQLqBe6eJX/LFXIVJjMsealRjI
J6U6VJ62EJ6iD24qWxf7Ff7gDl4lNzGiwcxn9RSFFZLyJPORO6Fw1JyzNPk1KNKI
DsaW5AsV4qg+lnmWlYbpoML7NzUZSO+b/7MPmmpw8U4FyFfzHnm6MmCNyQNq1LW2
CLG2SZlF3Zi8bktcBtF5fy9FHlWFAcPNYXqUKRDtnIXlcZxq6eI8ehOMuucHaFTB
1k9xK+mb189MqxMWvq4QimfIghGx3gh0onK3rD4uK9Ysba1azXJIeNKbMUyU9gvF
nZ4NejxJInxq7yNkuIpaeFH7KFbezFTkYUKhTfM8zhD4blPp74keNaoYw721gV8/
4Aw5xU5A2OceadP1WI5XRp5vD83VLTgwfpaXX0hDbvuq7J+lZUDx+9jKxE2eTldK
PqE7uQWmhY2PVxlNItzEq/19eDkaJFekM8El3fLvSAf8Eq6DSJU/w5drK1xSaqx3
N4ZtdEKWO+N0klMJFwMHFgeFD1OWsbf/NAjUVRdvXk98TcuerSex5Gz3Pl4Ev7sp
Jzrh18vFIUodpz9RIAQpOa7dwmUZ2eqdAXhbldB2dh5Gr9CRgxXaTmAS0ouOJKbO
gWdxY4W//ZE1Pcd5uGq65XaB8fHtx4i84NVfm0WJIilIjAnmDmJvwsUvAO2MZy+D
GOgA8KRpOnTZ1vE6MI6cRFACrkrftmIa9UN9FGXAqTm6FSPCS7vObiEg6kJ74mck
+2603NiQkSBxnb+tcEStr0hOQmbbR3ZDu5xBLJPf4L1lzhaqyfiMIUBnpD2NFNFN
brRs793QiDn8E7CYjyuILkbpBP58QZai/klE7c3LuRWCmBaYqSX3SzNPxXVFhQVd
hbcbWitBR8exB6C0IXOxDKBH1YltoWZWX3Jwfg7OfCluma2P6z0ATtptZMMJdmQg
lxwZl2iv4MEgioP2v/6qAh3aeSTjGr5aqU7jqStrgtpLyQdIuVGemlD307p4gUgl
92Qe7vT8cxw+lF7heSFAC1FT6Nm8yTEnlmFYH+weH7faj8lrj8c/oMJKekyZwLQi
MpfIeJeiLKJ2IMI9m95vUIsa/W0PV+ujUMfuhfAgwlyQk+kUs8xyn5++5XJU1JKj
w/xJcDRE8JTbVADgGsUWp0Y0GQjew8ns937wjXIg3HnmdWTAT83jty45TREVtAWt
2j8ekloA6LTN9nJ5Fg1rlJX6BURQlO2xmSFnEC+g1uaTbG7sQuYmHsKGLFVuxG9U
ANNvbaXNtkfZ5KoGEBEoqp3RT1yJW3YaUtBGScia4StMnJKRIIxnB8gN4bOgJmeB
c38Xsm+yrW0wqlz6yak1Dg9cbXrIoJRn3RYmn+ONSVhRDgE6Wpb2RbyP2vsT/xtd
0T2n0FLAH2UzNx2qJv6JyuqDdzynXjKVtBtoXncffT59kSY3P01HslRuqYGg9a+o
1U1xeFn5QpZXIiq8ILlGgCLSxL283UybpfP63L4dSBTqXTwr0UuNiQuP8ehcBr91
2wlV3mIKRM4XR6C+N9jPaH+xXisBLyaFBsRovycnPFpKZPAoDzntjRO+GcOC1YaF
vtzK+MxzNbyxS0vLnMYOns/+gleBjS9kDlgUVK3tVVluvPhxBOHY+JiK/NSj6laD
a+9TN2RwGGIkXU5w9tTu9y47ROoTAzXJgOA57DqYY4QWUmx78YjNDgBXMd+FGaiO
agONkzLHYDPkWSD8pRE+9UFIcS4YByjb/8fZ4s6huYRKV7IHgDqo93x6CMiYyOWB
jehgSZqP59JgKZ0qqLMFRGzg7iTjEAJS8/UgZ8O0r3Sst97oKSiqtN8Xsi4+8aZ6
llRxjmYE/f5S57ZxPsvmPm60bjGdcbWi0l5V+9FK+qVp91SQ9q/flDaVRgCrirm1
9+9kMXYrU8vqG/zk2XaQ1dFkv5ziU2b8/Q6EQZG3HXIv8QHjfqkhsRsjdTLEV30b
Vf4LIMkA0NLhCYoftFr3W2ecITi7Uk1XoWsw1RydMJcOTg19KhW0W5h/L6FieS3L
Tvo9Xylsr2HRWyyyh9i380rzzbbc/5US6qroHs49qsiJIsIozutXi1ONHA7iU/rK
k45zqs/F041YzNgW9UVyQAuiZDubC679rb5RXv4UUo48SRYU7F01CmUEIhypfoU7
woqG423EMpAwUbqKC+GWGwRWlXFrh0UVIBHCfH7CJPeEL2GT7GKxzzYrGmYT0mkr
lAmQ7/XNb9aSibLV/28etHi78bu+vDgE14ZzelaMSd8fc537hseCmjlBQskvHcyb
ayDe4cqjwWX0vHlKxpFQcNXg0496RUAfNt8xpSdOzLkdBKUXBBZF3snuCyE1rAGr
pJEVLM2g7O7eyesCVCNbrIrOvZl4JOW10aSwfBzsvAkURVwQ9WdS5bkmNSh/ryIH
7I5zN098qMnL93z/HAoMgolPS9PbaOcB9Zl6X1VbTX0BPBoh0oQUCR4jJQi4nX4z
rV5OeSn4mk5poFmv2Dl4w10wGxcce/lM+t4TjgA9O5pXs8YAe4kINSNcd2ZlCs9P
vOaX/FpvUmARaYBs4CQ2zUV/H7Tlkq6kk+3XEa/aobQFl1SbIaA9yDCUpB8OfilX
es4HwUyspzEw8JPPezrwwCKkZ4fRfiY1SAGbAhXGLZhu8rzMt8jAcQ/R1md9Uqvq
3U5kIE38WyXm+JJjewrydpZj+zw6r8REDKvTRGEFedbBhnwkeVKxGDSi4aK04y0g
lOoobKGUqNpMEKJwwjtaWU/iChRu3Hx1URp9iVUSusHEXSdbcKcFA56O0NiKNsNR
Uyl7017AVgKKKeS80YKCx9VyScnEhnEIr2YcrQlfy/werUmxk+fnpbWWRfXpt3kC
3Dtn/PQ8NoT/XFTWw1P9nLtzhk4IwP0bXuzUjG7NNxkxvbvLjcNeslzox/61/T0v
l/vg2wyBkiv9+0h1RPcfRN6C+PpFK18INohpQ+9U8y+mbU13D7r/cwBOz5+M5Mhv
dRB5k0SCequgPu8oVEhXBMpLfpnPEFY64Pvgm7Z0kR2T4jJxexpI9TfJ8MHhArFa
47kk4fHga2WwBUAb1XT0saBJH1/wqreyipH7TQPNQBNC7ckY/XBOgzEVznDIOQOl
9Uw5v99Caf5qwfNf7Q2W31pnxCzwB+rHzfrfF5UacUIgrYEyK/wVlnEc+l63KkEG
Jkbq+15ooXpHNPBW3erbI3QPrnNf3j2UeQrcwTB5H17nLYkHZwAhLUNWtsGadjRZ
R/qv2j3URXoNwSaxeP6GIYuMr9QhYl4Z+tzf7Na+s+oRTuDD1G390DVxZB6ld4NO
GrRK/jlltLcUkCpyQHGZmynv3OJx8aou5WIpbmaun6N6CnXAhYVD9CwqXPNtVOkM
6d4dYK3Qqq5eP9WfAzXn/rA3tWv5z1uD81mKIlzT3BoswR9qTfwbwH5LIwqtflXV
QOOJn1CV5ZtA409LwyxODaxEibXkY7JU5wcyTBlBSoQaiy5wjHN73+j/dLBNDHi2
1WeWVjLVFs3r1a/ggV1W6VjLqMHcP61OZY4tYV60OjozIxTLOEA30Fx8L6nsDCR/
RVh4Suw3l0AgyDDygZteUz+67Gi9ldMt/BG5PLz4Dbh/HTy9zrXPAvT9hDZoJjnp
F0oKl6+UKW4Q76j/lwoAKKT2wXWIx23rQNYVPBKn2SCg6P6NrXEPqHaYqrE2BIIu
BbR1mAEQGkV2ycLdTfCdw2tluQ4QBp7QQdoDTcGRT54yAwNbP2AZNkJOoW40dgeC
1PWTCYU1GIVSDviyPdJnSPsBC6GHymsEzxKzXFaJJW8KxKWkDCEo7XxUGoTUNkvG
HV3QpZKasCkF+V8vm7V+dN3H+YHDnOwcvug6eM3eV7tv5wXG4DjpjBFysTi+Bjo3
t5z+T3prTYyr0OKbsq+nWpyos9Jqtli+EKaJ0FAcGCdeSe2QvMigMX86WvK4jQzY
20RZeYVn14h4UD8EdLZ9xIrVuardcGleFBoqAVqsYVnTZbZsOL79ZWm8EabtZUO5
GpViEXLZurGIDuLpHjHoZioInkeFeu8rvLj3gOxruzZypZTFhlEZxw5PQvGwE+8e
CRcseM/vJsaiZVQH9PUVwHLkScfS2jSKlZKXyGEhK9rwSxvxlJ+yXL43ACuzZrw4
vURC267FqyBWfYcuM9GAw9N+y/5+Wyh06ppzuJPUxUVjSJiaV8CBGGmOG6INsv9F
TAXhEXpbxv4eDaYEBW8xo2JWmyKPQJwl2K6CFlCtY/UrVn5ZBozH0zK0mGx4Tgrs
G3RbYKJCUaZPbijgnc9AW+MeHxIbCZI8T2xefYkFFA5iSF2vVzqFj+eGg9sv6Xxh
utdIc0F4HTeIay3Er+rhYWG5zj+NLmH4j2onmE9oZSuzVsYi1Qvo6Fqakxr82MOE
/0HTpsJlc4v91zdGu/jrpL6RUT06XrWFcuk3ro0RpKnBDrbSLkFxG727lNGA+89B
FOPdx4hiXXR9c7pUUCmiXk5crIusb+ZygNYSRimEL8p3flnytYz20lwsZrX0WFoP
07VUpAsygm2S9fDAK6W7iX0L7qGHAH91j3scbnMoFAM2hpEfZNRX77twsD4BocuP
nGehGp5beqaCSNkLhFlxQqX06yf8D3SMw54keZOEUIS3u+K+sFrm4E8q8KXEGM7O
26Y3Kq6tAE66IkaeB8V7A5zfdxp84OCnTgPSybf2rSPjRIzTR6LL5EnlZd5PXgZk
CIrJKvpbcQ4EqeMXZbK4XnlU3h4VbTvz23CWQtFpWifLkHwKY9dHuX46CpSG741q
KirRc8V2RrVAr58wx3ZPKg1n4nyIwJi+rgRnMR5BopYHajpS8l83+x2chsS9O7PJ
EeaScq+8IB1kQ8xbAnYcqZDqVM+GX8bsd5u+xAD+WFig5N+gIphIKA3W/9UR+tAy
JOTMzS6qlg3gpGP3rqLCyA1IrnXqKiWE1hwDk73cjVy5jLuScCDjQL3yrvi10FSM
vgqZl5V6WllN883OB2F/8QJuJUZMEqgq038ViFvmDfU2z/BnXZE5CXtoFHU+Pema
0olLjkjbGBKSvXCHweKXintNms7pDY+df3JeHCkBs4Gcm+wQrZ2TVMCIum7SVehI
ttxs84WULpVvlrWNQYwVk7q6CYjRNdnF17j4aGpl0pIPSZ5ySDaAyrkNJMyCHttE
b0O3GD8FhTcUTW0JltYJfhwFUouiTQ2SgvOzyKLVWFO5gnLYaW0XPLwAgMqazZEr
Qic547FgJlN+QRckps3J8fo4QcCNrO1Z0qwHFdXuRBtuE37YL4WKfUjPHXyFWZtS
uhiz6VJSxKTqe3yDUiJdjsZZPbu/C2/lCWnqKq+9gdEXZUKSAi3P/K+jXK7aUJ3v
wwlKbQ1CWas3uaAdvf7b9FIzqPeDRea771Rxh60S2GopnJyWln8Tk/7sJNMIqQ0J
xb/4eIkW222sjaVn/K/VjPf5YTqE8yDcre7rm67UfOcUZztaIKKuKIhz4MApirBk
trGgFNvSBAKRnC4nZTuekwKB0IQMkm9ZQcuP0J3AUUSuMBWHW5bYs5Z7XWSxMFjv
/EMf+TPlukQG2PuBmAkpG061nygxTrp8yHETVHs4Gnf5BOP94faCBPRaDm+CbFfI
tYcxV+4+iByYdINe0OT3nDvEjwdZwIxIiMDRtLpkFDxh3QNhW/Mwfh8czzDO2EuL
Jxb0dfRQH7nlz1BjrMqQw56r6Gqk0jdxxwmam/0AcnKnO0bc63kyqD2/nmEyID0V
mZTfI8dXDZq+vq6gmiAzDYFcodf48yz1sz/dF5ETXSqzL75gjpaYqqWVRNPyTfwh
a/WRlTDiizB69gm8cuQxcNnx5lutPGZ0azeL38yJLtR5fV4MP5hj++MTicO+ZIph
nSB4Pab6U71B3sYGeDkpYCHE7vp647Am4Txe0z+Z54Yh8HPncvHUXYDL7Zu8gttM
H1IhxVaNds9Uc6R+lOVgqz5SWM7nUwVtOEMGKexJ7641tFalw70lFlvkO/9lY9YC
QWmDGkSTRN9xMKQg+3fBfSAzSRSgNb69d5p/R/rOgh6zENrgqK8s9YAUlIeUS9eW
qgP+Fb8GO3V+jvl/gzD23oo1SxulJlhEuYmNu1jH+YoaYQrkvgsLNBIpnN9cAtqn
o4EjuloxZNVpAWUhI9TdBlcykDc3C/LeZ6STC99YyUIrBzgsQv632EI2Lmv9vdLH
ta2MxjXVOuP0KwJrIuQOKIoH4xtg8y9yFWiLL+0DNydZDRYYrhZLd37+bcgO4lqz
nlZtu9GpnuKh4wZ19kQ8PoQTmSftTI9pP7BznQbC9gVtqFsIF9ZCzUMnyMfiIENa
ErLBL590pn4cBz1ORV9CUWu3GveTNCgiAL0Xc+x43sVQaVt3cIitx+epHZooAVRi
TXsvRuu03wJcU7QnZOtSe/jKFGV5u5tvouP8LLKqYRSjOGtAFsnQIzEJq6GfVwfH
k8wyfqgq5rEoU+sBtqifuaFBTxgeQw2a9dQ8RYjNoOG2Iba9ghH7EESnaLEUwrM9
3pyBD/djosvm4M6H1z01gH6UxjgZIzKmvcO+W9V5quTKr2EtIo9YEuBrCErZWT5s
tveLfDFUf9Nku6GxAeiOkT0hRoa+tyTgCu89iZSLS8tGR1ZYwNs2chZf12CSkIOQ
HPlQVoI4NpdmMGhxr1D9eiEvoyy7sTtLxohR8GLhDRK/MXOH6fqHdYDrd0kf5ooO
JE/LrbvZ8PwErJBzPtTkPgqVvzfKsM1uzF3tRcq0ei6AWm/vHsZY6gtYKZWeMRCN
tfsGuF0yB9ap7pz3ZsYr6SQexcV5ggxECMgupyKWi5WjrHhKAJmv2JPYVfSe42jp
/fNmypaLa0gKv3gWVq9OqAxI4DV6O3zBEAz5HX9cHx06wuJ2a6PSprfJSQvOvkkt
qRGf3aTlaJMu6oQK2FPH0jQDkA8QqZfkzj1wfKFpqPEADjKBz0DE64dTsK7Dx1b4
0qNL0yf6NlMYv11HMQvC01SQRwrqUn77+d2zBqaWcBdXHozTxZK3q2NM0Zy5LiJk
y+6z8ojlxTcYfIc6OkmJlgHvSVp6BwFoLWvKys0pJYoskzYTtZuh2FwbN98uZuAW
oC+9grlkwm1DgWXkn5a0hsY6mpzDsgrXaPrV6SAR2DLWf4aNFv21dEnRDtBH7xbS
zpm3ZvUEz+7Fz4hjYop6IgzEwj/+reYXMmWqtY/BXfeVfKr7KuBIAMW4MIDJHOYu
Wl3g1URTs+LzsVFwe5RUAIhLafHh3/f0AK3RbALaDFoUAGvTgzX7efnmdQas+YWx
3sW4e8NQ2s+VOWoqByjoXp+r4LsOgwo37AJCy/2AnqBft7+WWqUxeyp2pGZ0bYhH
GRJZDbQC5H9/2IvXzFIZe2nbHr0mrYF2aKqgy1iUIaU3mGrvIKNjh2M/a/pvkBko
SffnsbHsx897XP1LBO2DJ/KbIQT0QfMrRULn/ZN7/QVnJx1EflhsupMXRTOC6aFW
Acasy2+ANz7vNDThwCcCvfWZgEHJ2zE8P6CGz+AfqUHlj2YA945X1baqyABVX/0m
WYVaN0XtH65CX9Dj7tqy24Y+r7V+XJEUGo8+HOLvXoBzidYKYLhRLP1Kz1iCKuIl
eFZAnjxzTHM3PqlDSEwgRfYvDdcw5DvHHFEgSa3CuQmlssShILHt1v/6hZeWGK+v
awUvOK4/FL1ygSaU9QNHhWV2XWd7CcrDSdp7igj0tid8glTWrUFLvXhf4A2ggKe2
ms1YafUhacTyEPMHak9uL56u2lmPC/dzC2aSvmqrS6egzrwxkp46/yy3AjaEvaqD
E+rthM8IcAC4LcxWXu3YDSefhydT93kOy5yM1rgnyqx0a1fM1xIQzf/ivRSwYmnN
Kf7Vx38iHhve1q72r9eCf3ejZ54iVssgKmOdle19oET9ZyWj9kLxI8+KeiH4k5m9
mnDZ+1v7c6ptqANx/R0C6F+oSLDln0lZCIHIAcXkhVtodgpLBg2UiGkoyqdMs0Jd
Vl6DOTOK05fLBNDLmnFkvwa6fS4K9kDBIQ1n0l7T5/B1GIKMHS8U/yi8o32Gz3ut
gO/tzgiDQA6wzMpx5f4DoJHk8KeeztgyKanJFC6W3Z+6iKBSdFWww0ycgQk4mjsh
OnxwmfWQ397jLjU00qGgCCyrDMI+ucdauKTd01EpcTtMitvz6BnDn4IjRCEP9Jgn
EZFWFVYM2O1F2ZKUclPfl1k9mQ7PUgK26OABLvUf/DFbae7DWaVRGmAz4A1zq6EG
a19jaAwE7lNZOf/N7UBZfY4v60VNsqRineC+JqNXWWWNEoiGOZ3XoGZGcBqeh4ZT
TvKudbrL1wUdp0sIr2FrFblH32mhAtS8nT7g9jOamooe3NSo/tvOxubZnPxn2sZ5
8ZSTkzOhAs8BNQYulNBzpJapwhWUWxgWWFEepF8SrBQzdKO6CseiArNANjyKbifG
lXtQx59jV0nnHzbFXIujqBQ8ZwOAhvwY6q345p467XkWAQSJzRv8dTByNmPSZMmW
ZEqboyUtUTrh3G6+jjMO5vgjf36bK6aCPCRpRy3v6bpuLbFXMnT3/F5MlBBwXusK
tNlCzTzKyhesonWC4GP6Cvb7/Hn7bLr9yICLJah+Ylmpi+hcAYYdW5SOpMIVBW7H
CjPZNm2UXFQMdzMPJXeqeDaq9yWY1Z4gk23rLFyta/HxCs4cXIS7KAbPXdlIycp1
Pm3GUqjYzGvhXC0EMU8mTE2qMLHzkv5p+Rf0YmWHioSRr5RgxBfE+u+yszlBa46a
VNcW79Un5A3hY/jVqzYVCBgCbTcSpvGnRS1u+C8sK/t1um1RX96qx6yrb6IjwCAG
nov7rJcZfErmCZDeMTuwCMRTZucOGnWxu3kq7NbEwEUR7sE30iphQ5nedV9Rtfx6
vR/KdMxIVTW0tJAIxXdngjowi2G5KQsl9f4GkPeKnEcGDUAG/UM6qwZUQ6rHApi/
w0oO9bNWjekZ/foiltAc19L6pOFHc7WmG/UiMJdor5/Nj7JK4S9iaJhY0WUIMDCG
hEI5Qu4OG5BcKnPmvHCeNGW/PF/kli7JViAoWW0naccYG3TNaRnUv6Xuv6yEcds2
ZXgG1FOyJhhkRBAgAOZ/snO7XryKlyw+w3OysKugYGF208QEG26MNOJsfp6zKv0E
Y+lop+E2eWuDHHmHY+x8IijwtxeAfQZODx+Rin1rpvv2mZJSr4YdlBz2n+FO3dwc
Y+9ua5NByTUn3cnlZeAbRSGhJTKw6IkQ+YAo4t5Il6sX8V6gtssUU+tNn/Y4rHlC
+ejS5268IKdtJ7tEKomPQ6AVPSOuhpETAD/3qmHFzO2XtpaUEad8PclLTjY2lWb3
T6hQmViCTjBwBClHD0gYOOe7aZPaDl+YdmbVOTiLU/NZCxWSdUlX2Wp1+5UeXruT
0SZUZ+5oBZdr2UvK1q+eVRR95pe6GN+RvM4PZ9R2dEFdxcEiGyFUKxxq3YNewrov
v77wA1eyxnNbmdrswRu5wibXXRbyoskRdHSuE1d1l/TsXERsRjbAnq83asQos3Rl
86pW6ELT0XsAS/MJf7gCbZ2oYqfWny+lllFMCgUyLqYQ5TGGtsoZVx/d3+VGPiLG
m80wTg4bemZKPSmccmPtW0croV8u3dmgD8zbfjc4xBwBpzeIz6iuvjFHGLUxweOa
J81sSlPDkQa06XjYfmJ5QYWvLnePwfBUMT56/ZlW8wgrmsEEO6f2zcnMrBc8aP5A
Y++fGquwNhY69T8g66B3bdbKUmRRyzo/bqQJIopq1WMz/tXZiahL/3RQoYB1YiTJ
HMlCgofHyCmkHvbs8JSo1eS6ZqM2OewJbksKbQHkjXguxftsPryWChW+lq4kFtjb
72t1vOsVf/gL32hy4A+6URoEaqLqKb6rlq+Jf9HIRJwgOFzhFU7SVfpZIorMTXBT
5dYCMjlYf2IaLfCu00od6pP6jMr3dyeiwnKNSfXiUPsdWxXGcRQLm2GyxEhjQHc5
85Ipytq4e6fC3ESRAn9YBDedGTne89bjRl6QS+fhM5MRDVaynzDmoCfW15sS+qNB
Ex1LVUsjc08luZMoWPSxZz/IJlrK4et1P+IGraFnBxAohzsz6ZErKUrn4EqSeuk9
b5IXRJUacoP3QNfCYseeV6G6qQw9gTysQ40eAYD7jmtRtQ5mLHC5Bv+LZ3jsBC8P
YTe7oKiIikyWJG2/Amsw11qRFDfwF42U5366xh1IvDvXksGRmbvhRuIJ+35DGohT
N+o4Ub+P81OrVZVWxI2rxd0CNuI66pA8btqAW7WzEwW6ytYTq+ZjXaD/1CNTcS+9
dveZAezrXVoktPSpuv+LZ/62Wz+kjoy/AHfSdnSFnOMpMd3HdPCWVotXEAKYHXtj
WTlOmlIo6X1W6ublRgNpe1v+0St4/MV8PXbYFFQg2hbYQXQ03mADN0KEwxWOXRcp
ZGyOPZohT9Jr5w/eOrmbQNX1gTufDNKeMunAQiKgwyd3+Rzowc6wd8vHsJigT4cU
ttGSU2yHI3IJbpRd0yayfnu0lBc/CoH98wmHYzIczYhMzhQjwiRcl2m52jwtlOhh
2JVZesNkEUa5ZHCCBVL6oHukez7huRMNmiSFetyMnOP3McrUwcDeY46q09lObPA4
C/6BHLyMKYBeRYEWQHZKkv/Go9BR8TBKsADpHLY3qcMQysC+MLTmEo6MgYacnPiB
EE02QD2Sh17ptgRTzNHaTXJPBR9O/Fws7/2HHKsl2SeHD9/QfMG5DTFNhBtZdTqV
1Klmf3y69rFAb0JB1zqWEO/n3ApMlFYV2M2TtCY/WsQRRYJZkTkyNjkyt6oncxnF
7hllyYZ7frY+9qEEM1ODTW/nrxR3lXEx+OG113o91vHRrwXIa4CMAHFDmUhEK9yo
Q9smaM1b1+ZeEKveOh0C0edXltXbpH7Hb7lWRdgCX14kQjbLTnHKwzgQz2Pgtw72
QMEU9WvTR9FJoWclnlMcjoj1GDfijlR4IO0tKc7/oT5lOtc+K9TBDG6d7T3Gh7W5
utCPdzlWzYkobm9qZvy3C9MvOnkv8ehfwJqBFFEhbIfHu1nKsjujhysrdtlEZ7/x
e9KLbN+xtdPkshUZtA9WW/fVXIIh8Y2VGgh8y93iyQUM5x6dwHfn0sOiIsDCOHhs
ooVfU33wIqDaZwAHna/7PbuK1ieqc2/vzBxl/qNBYicSJU/c+zDFGg1Tn9qwjdH9
X8yXDT4PoCAAsUqLPEjvC5f/FbSD7W2NwMppnxVD7qzJhdIsTfYuBrHEr4UONfL1
GqQFP9z413XsrAK4SECwddTsEnO8WP/BtD9mxojDf0KDRXY2DL5Kbb4Sl2hNXXaX
DmoeqPQX6iD64EOge10dgDQs2/4hM9Kt2xF9dQEOLIb3Sh1OFFQNgx+EnBRvmwT+
d9WUJ5cLUlIlBlXKsXdsMikP3hY2/N9HtdEPLvoazd5rCT7PvEtjY8Q1DH4aPkL6
ldzNNjBdhwR7AbVS7vIhfrFgRrdgM84aNS+YDHPA3r44rr8yw4mvVMv1LUGu2K7S
zTEMeHr5XZ8WNm5M+kJa4mbg3gCIIlZY+Bk4zziIeEX8Vreaz5qN1qWpxc4GFzrE
NuOjlmyzjZ3GH/sktSJdOPFW25zJr985pQce3k+jKSlHKbq2pEoyLF5pqc/lq7GO
Y0iRc9yE8VRxhdjCnSlEEPewOlJXEDYGfpePj8VOVDQ4fn50Fuxcf92RzhsWtkH8
Dxs7kTMyhqQbGRh11rcvvTn24ZTM238dnXUwrUMcqUypaXlsf/BYBuhTjIb60s70
44O2UOvTxVgzOrUVt+XvWHfOpS9kewB78EHdcsHdde2G49hCXzA4aXlx4/szELyh
rSrwfavJLhzlpntCVa/GNfY+ksOmoqVuub2v25KeZ8TkPa7C2PYHmU/MBjLU7DyI
m0/7Ulr+ceUV0WUyH0y8ta3Xlkjk0MqgPx+bqkaiY3pPZSRqa5TacxInTHA64BRE
NR9f8XtbxoRc1+kxkQjKXTA6bo/HlkSk81hF2jMQ1O742zRaWaSI5Fneglfp+XB+
N0ukU95Gy150LLlXGXaRgacqWtt/DRQJ9sCLeiHQk/iTp8Jm8m1crZCDuogaoyd0
OGnIWH9Wjn2KYeqDy3TGqTwtBVwYU74M1AFtrWKiDQZ/n480OuJuYyns5J+Bgtt7
Z26RelHCeIk+U0eUorG6OcV3r97MHVVmIUu9j9Jnxj7LoVYaIEUpCC3qa2MigUpq
rPaOCae2DtxvvOogAtXAPfg0zviRQ3L36jPlkKLJbpiWQolADVr2+mQTJsMTSeJ6
wwLufEABW1JBo8wlOUywfN29LUTQIK5DZ9WeSQ7k+c+rzBiVXr0OCGxcRV65tH3z
uD8yvOyD3yxliipB5Jiuqkp+p67cqhAyWtWWzEOddnDo6OLcWfwvP8haNfd7vzSg
/+XtaVlYHUI8OFlzHFUCrYlS2A/OKEU1bfiIcxmqr5Q5wL9VpPgF6CEGzZwWQ+8X
N3MXMz/NuVRBGiJvGpdiMvlGSRpAnGxHt0z+ihjVea48hLGAIW3AFIxYRqJhbseO
gduT6BknLhMoPFkZn4NpMvJVYlvAWHYWSL2GOe5myk0pgpRE9bZ7d6bWaR9f5yBS
mCiWob5u/IXz0eunZWBth/udv3ZS8TtA8KpGbqWXzDV/1wYFQoDdAxPf02em4F4i
Gki/J4uTK5oKfTJtgSSZpKhoq+lbQ1Rr0EYn5m3RzZqElqTqZNYXrtDsAmVnpif5
di18pfHVv1yyM3GsIlSEX4sHMyn+3oSFtiUfhRUuh8UlFHb84b0Q1um2exCMk3IC
CPdhflRqxXqeNo6l4BYl063NkDggDuYkLotHYlki7+kjFd8qZ7yHUs0i+MYSqVhr
SRsYn9waokmgLCg5CvDGtoVqQtLN221xmSCeKWqZBjbFNpdgt+sH4eET7n26nwOi
34n9Z0l4pTFxRWshy8rCxDhxBntDynh8ILe33awNfIpSrRYD3QUEFnK7+9nTwg/6
9lAQj167rm8CDScdeB8+EeVjmcOJqh9kx/tK7c5xd72L5efJgaCCXkkbfc+6IaaD
vWFyGEnMCgwWIyhgS267nS9su7eUSTA7I4BORTSlcCZlxDdRxOe23R0FiUh+I8ix
f/j1kwPW57VEo7ryK+s3SpfJwo9SMXKqiDTRAEABxPkyaWgaTzPXOh+yJKquHYT4
MQyHAQGaJmGkbaqYqaEIKxgaF48MbiNx4VtDeqTkDXUriRxAUmf3lePBNEtnwLfH
SLM0YGj6j+8025HSO0YyH1SquwdPQFNEo/y5Zbmo7sm7Oyd4crsObrtfxvX5h6uP
22zxOuM90YajoHbtpXKx/BiDPXWtb+K+2wZ8q8rZ2tmGzGix0J8mXHzsFLSgYpsW
fLxkoip+NwLdzffenlFdmURSlSU6N4c7wHeHP/Os92zZTkt/cnor259QW5EofXI3
ahqTiYqKojLz+h/VBdj6xmu/wDIt2/R7qJXrQzzvwY9DmGaMsYJnUPpMia/tGR/+
5IqthAIauHyjvCYCa8Zx7hjRAfMkJEh+1XhLRbONpjz07EfpM5UNDap1GwsPm1HT
TuSb1StmyHvYnxvLVflKS+co7Y1pQ6+QkgMGj98drobtfxu7Rs7qya5k5hgP1zs+
4ofRQjgkOB8gbZkMSZlx7BuUvufSElqlfzxVry4fHoBBVZYD9sAN7xbbjPUpa/Cv
XRrtks7dd04UfD74A2Mr6nvNylLxiYLxcwzRG437w/w8a9u/1UjUReMAIuwfRHBT
6Ed5oa757A5PkP9+sn7x8yOOfXEmeYJ2SA93gwSoqEbA/lyekWIzWdrJupKr8kDZ
ZA9Wgd9D/JJqahqxguLq27ZbjUO4oNV9CVDmmbhV1w85IbCEy1nJ9pMgu06yCWJh
k4tzjYRxJTlMAOEOtIIGiYMgpOCYJP1BcnWken++tPJW1XU8A85BiRUZ9t7N/EzU
LIOeef1Qvj1sc00VJUQpOijWrnCzwYMlGius89Fr+j+5VhVTJHjW1dB7PCJ2sZjs
cm/2Ag/1QMUAC/NPRx3XnFrUdF2LaATBPqDxKX+vYkzVnN2MHfv9a3Id3WW6efri
3h+b79VspUXy7G800eaW1XRTAbWW/fIL5U95x2frvpYUAoGCU1cZ+nJIe2kuruJy
Vn7OH8jZs1UkmPXi38rDva5jv5gTQeNr/t4DI45lir+FGQjbmjDSStCNW1FiG2Cc
3g/crVu0i4Q1orKN8FOUtU17LB+mfBg0gFgn/Kdjt7bXMjbZgROt5zrsK7ZpL+JU
ZoBmAFqyALNd0W3IGE9RXHWxl5rhbAsnLvsUvaY37jqcOvzNrMQ7SwWuleRY/zjG
YapvNSEWIDfJ6vl4XTUuRk0Zl0RLHhKEIVmlbJKoOitEIZgjCegEuVOGF2aaemc3
eXaJp6NOt0+3AA1fjMyQ6BN38Emff2Kqh4RvgNmXFmSgJDTuxsJ1LhcAs/+bWg8P
sV/13kkWP4wl1nBG1DWR2XFuqBnda7Z2Z/hoobpXhVKqtpYJ5LYDMMgkekyYodPf
8+zAwhAsaV2HrYzEVtFfkEq2EzcXBZI6hUnJ9Jgqf18UlZQDOQrqNLP0XMjK5bAG
MdkCK3ueA8Dq5Q+3LTAYPQUL+DIfB/7S1DJh6DT9mK2M6xpBkpZhb3Zfh519ubBf
kJPoJaQRE2ZnPDHUxJIWrwYUshZenMmJPjzurkITAezQvxSbn48V/iZS9jyYz//D
d8aUJ6w7T06YgYFJDVIoyfZytryr+nrQRSvb4z8LjM+g2NLklyvHMvs80T/h6HA0
AByBjurl5/J+UkqhIR++ETy0iZvgP4HvXmcGhBs/WfsNnzMnlHmu1DosY2wRaRZ+
YC44zCW+p0Ux1GujFowiSAQIdbNdiDJqy2Q+6C/FxV7X2LhvLw1PovRcj3a8a8yx
Q/4tLUF8lc8IdrrvUtz0nNRMXRGBCZkM4Hu3QXSPiN7QxCDgtc1IIFVlVhKxdOFw
xD0pu3TAQqfLGZhWN688H6wPPVkTZLCyVggELIiMYxMwac8UaDblkk4xC6jpL20l
p24v9wQTZerPq0X3kHb26brFqt7VB+YhvsQSHuJlt5GSIvDz/vbCSpZufQqlCb1Z
bEZqBg4Ze+r3KUppQT2Y6h2Vd0NtdH4/0w6xGosCxCBewce6bO0qc7chz/Jd0OH4
O1aCobryKIIL5I4ZHV62CIc1w65XBVfsQ1OR2F31+GoLzu5wEgVlGNMKKDVKnI/j
LSj+ClVpbwrldxYRXWDLL27WAGD8mgtgbrn95TBHcgDIZebWTwu3LJAg+7/S28d7
tUlqWen9bU6iJYeIAXBL5br/0XlLSZGTTJ6teHFulu7jf/1eWBo0UbGiV1Rytfnq
1p4YpLOjbCfL4TPUTRN5YyW03fNxdvm0BcqOTRmVI5ddv6tNivfHLV4lAoFqlX6H
6FUxaX3e72E8QsdQxi6icxXnNNrmIWaZaeOabyfTMlcuaZPaiGdv0TQ4WEZPkRXh
0OAGoTDyv06pC0UuVJ9dzS0nOKZlGfc5q2B+mY8lTUTs5G7r8h/Gn+SbEbk+xiLy
0uN3sqTThHphN2K9DYvkL6bfvWVJTEBFz/7YDqBVg5Hic3Ex1+Ktvv9Ox0nLlcN9
ionzb/J2JzPn7i9jn53R2dydrvGzPmqAUoae32TTSgIurjuQns0XXuXhf2+UPNMh
lSrO/zUVL2dF8Aj3Beo+Zcy7kmGEka8TctCOiq5u488nCia4xtCrOMjOBNUclpUh
3yF4qCd3s78I7/H71XjyRQZZtcqmd+7cvDmA3dLZhJUjtyE1db0QoefHFZmvqdeZ
okR+Ian8HAY+c982o5tbhSsZ6hL+H3DB7OWsuyx2mXzxpJpEg00Z+ptoPn+HXibg
CLFGGtUjg/uTlh05DxKSLpktRSNjnf2SzQiDbOqWezF34005vyfnoFpLGCYbo/3p
A6bo+1+lo6oN2CQMg4uc8ezjHnL7EeDuKNT3LzNEFvuHofDtViU6rJ3UZwB6j68k
5AgeCvNP8VjNualTiOa000ljGIC9JYvI8hE1Ys12ZEoZF1P3D4deEPbaUTQiL0+9
1kA/PDqKJRmcCkjcHNSIFLTIEtrktwpQhN1DsJ/OO4zcmK97RLu7/7wtscPUdDY7
YUdSezpVBtxs/zsSb5IpADzaOfpSTBCgfezvxZzuzE8x43+9koAPirI0baVsYL1A
Sr1DRqSK4Mi14IVuOnRnioZUfT9i2PrBxpQlx2N97+NVkb92XPXGMOWM5j34wZaM
WSWv9EnuOjnpci5PnkZ3Q3o1KZuH/1HXa7YzagsZuBm8gWnGpzGZb0WUm+AYdBUU
Fvm9EwJARQORlrBiqimgitWhlGhmbDUZ461Fkqg75ZgRIGgHh2HUfG4b6t7+2zSK
ntL4U2+b4/ZMIxjlCMYC+n+ORW+rry2W99L0sLN/fPyohLAxdTHH1cT2Fi7q750q
I2PUd5kCGiuwrl00G117FBtfYvLxlFdMRL5/FxMNwEIAU/uLCQbWMozpuAaOnBC4
g/vuF60sNf7KV0ejOUCptBB07l3cbjgaP8egmWA9429dg6uU+kOgP8qhTyppZjR+
ZmuUMyGCKSw8rm52DMcn3zqzLJEHsFbYVBohvTDRmPtvmyaM7Gm6HTjNFfOGRd+Y
DZt0Xa2IeleICT3IR8BfylU9gZnivg2bxdpZGUiF7f5o9I/dNBXRI643TDcZSeiy
p/PlW9cZ2b4wKk1hF0wySr9yCdY/76J5FsZWDhtolW7Y0MxV+6dCU5gIKUm2v+oI
zz9NyklutL19dpesh0jbH6EhPmkH2IT9obYmleMZ+0mP51UcpEtc6+nwPHAMWjPe
aTcFDduTHFh/2GJWfQxiAIJjLlssvVqsv0nkgry4adHV1L2JXxP2udPOzhgQ5Dbc
KqZ5IsipKaRG+0/Zd8sS45cqtkJ97nZQ+fp2znhhSpMxMxwpIPjUMTf4C6A9mBEa
gwRHw+l7Xxvb1E38wQQ5Z5BHtlZ6oWRI/qsWS0ItEGNhKEAL4Xp3MKUMV9BI9vsZ
vmleCOa46wDh8B7Ch9mSkPn+p17ChMI8uTluQ6IYGy8HKYbNu8u3SaDKNcYsiDER
ZvtygAPToD+F2wi1jbttSPOs7+7nBLjAvZfgdfg2LgP67zxFo5Ypm1F7nCmLx6IA
ReGSS60kpASIBytnWisUN692AtaDZVLkG9jj+hyMzTw09/wNczZvDqjFzgNP928E
0wG2fYbPHDK4jrmDL6o+QO0nBu9gIk8btpIGWtIzdvdpXH2MUZpNgASZDquy5xLK
1d0M793+Nr/tO7KUEHMCW1ya+u0fBkCLQ/6elSBr5yucyv+37YMDY21pkMyRp9tJ
7BTbIIUqWV7UuHQP/w+98K/8HT6A+1lVYwzuaF4ydhQKel45INVVEVtgbk8Vcowi
A9BYORTNTYz8m1KVKu/pOJVTqUTVjoPErz6a04XgTZ4DgpAMj6pX3SZMEyi3+5DS
9dhE85N6DG5pACa00uXbSFZ7bVamM1o8a5IpGbXgcQUAPR/4kgE+Mg3wFp3TGXW/
j/lKZdmyN80SQoA16vErgdTYI2uyMYUGC2oBVWPo5wa9RZoPweHsjzseqh19VZ6F
Mwmn7sBt7WvcRBGsXpgWUsmGJmLZBSW+mN2OAPzT0IoG/zaji4z9++V4jbeoaLue
ewHUi4M1X7KkneOoK9E562KjS3zfCswg2qy5fcobowDlKj/Perjf4uymA+2x4QKB
C82ULR9UxLjuxXmfYvbksdToysMvwWFwv8xeAnm6S+mBlFAnwVCBPImg0OXk5HXo
viQcDe8U7wWbOS2RoRIUrJivexzMw1ZoGUZRIq7AEh3BTb+r2mGsPZgiTe6jV0vr
w+fIGazMyN0NpPKYR6F6sdA0iXtX11X0enZVBA+Obpm1UsGUT3RDsCx/8dkWAHnX
DABUYj0a/KPFvxN7SoZZkaUmrHcgNA4W93zh6ukNp6EWG4qFXwVP8EC8XsCecAP9
KRIVagZHy6UxdHxWPF5IRK74kyGwPIT6kk0o5CvhKBkJ+MxDZIpEwNHr0K1UOmen
xIeAwq5EnJKweZNrCSRfgW85TBwPHJl5/I7Ix0ngjQDDaL6MUKpRM9+jXzJRvlbv
acKWMM3f+zgY/3j2/OHL4ROuXvnMhRip9ji89Aqt3A0RyuVOAm5XcDDTzXaZJPpK
XpQvUDZKKnInJ2zUdPF9dlIGT0Mk+O/ZVLRTFZUgATgWIJXbT/GjxzOb7WNE0YfF
HXiuH19rPW1ROQ03qd/ZGRN810fr3G2Ckwh73oOX3+xPZptpP1BQutWnozHS8EbR
wTZBiFiac7prf1IcNg730Fk0OPlImIjy3fTmfNYC5VdSNPLQNrdpDmgcansPma2V
mrvah8vZSXJ/3pFsWIAQYXu/LS/P8ZAcy4I6pcLxTyYIBEHzw5YiNdWmg176qFSD
WTRbJ1Pc1gVMTm+nFWVred7l0oVAa3pQzDf4eiJ8G0kiw9ZoRuDjxrgn3g2zKs2K
k+ABbiWpNxWXlDE4nq8rYf1x81NWibkA9ilWSCupKBic3TiOTEZcmvpzNo7LcMWz
ANLKMZYreiCYXWn1CZZUn2jmbXS+kdousQBMX6K/RAN7A59bO4XuuWWjzb//Py8N
Dxga3IhSsLi1VTdeFFY48KkFGJmnFkpCCaY/vPowIYeCuVnhttw4dvnDebDSgBud
hVeUrshEsP8AwN6mkS1aTxjJm1BIIyDkpxG/yYpfg4XEOxAtWDYNNmF37R0ojT/M
jXDGpXxIYGDH+Y5PYS5U1FDp+dWs3fo2h2RqSSbkx05G8O7s8OI9s2uzKgFyeyU2
YHO4CyyrWqRLaOymVLJbPo0SW1aB44LZGP3kQLY41p+fvfCweY/RgDKA2hI4d7oq
wtnSIeZJ/kRGT0ADfyC/inhagcTy7v0h2Vs1dkfIvYjqfV2+q1RON+DgRra/mJFh
EmkIEgNmCcxLrkVg+dd2QjybaB7Qn1gqbQXaMXLpdeFudRrSaCKUB2ky8B+i8lXs
7Iq2V8bkyUpyW3zcpDylNFk3XIFAZS5h/uVaqlkznwWpCRCnGULeDlNTI2sg7bgk
4uPhze4AHDKNgLl2rnqZoj5pmDeopTSIXms34fLlgOz3X27ni3tAZrNs5sPXBH5S
GVpBMJJLvxVTcUEO7jRkBpg33b7HGJPQB5Oc5yL4U+WcOvU4mxy3V3EzqOiTBT+Y
8bkRHNddMHsfOmIRnmFau9cTc7SpbAbEvqUrpX0V/82e66GVeUw2YVebozAXkXaO
ulvOy7FpwVPWeYNBASYpWoXf1FLG/Aurvm5UlGPweF5QDUkMLU8gQWv3Z6OjI8p8
U/xDs83laGbFmVzwTMMvqrBkuNjfocaBNhvCB53qGaO7tlKsysvtbJiP7zbxqlb1
WdgF38reVLeeR0iIxBpW//fVJM8Wm3EcogxulxkJZ4SFOff5E4/uaekYbWLzXdNC
OQHY4HJdG0i1QSyvcDg6qklfE4phJmkiLPPO2j2EZ+EP+yra6L+JupeUgTZmaCak
TjsDoEVhHwBVQUuRAYa6i0/nn4K12HqXLBMLRBoVtb60TLgLOcsZWJrd77OCIPk0
6idtgE6I0mWPHXx9gTu/R6+3GJwEZBhy4jxX/MH4e8nzQm/qCpb5kBGjY3bn1R5p
7AztP62bVLtC9OXuQAeiy+lz8nDxmj6ZcF8kMIm94F9wGYGBXkAgO94C+pblSY64
uvLQAA9UBdsgkSzuAGSzjx+fVR7gql2Xobn8QcGRbkNehm3MmJ7y05rwBfn0LelI
E1GIdSWv2Lh5p9PteKADKkjEW5gp0TOHEWoUzJEHdYoA2YSTG5BetKH8LQJo/nY7
C+E2mWohoLv6vrQQMchJBEz832Oz6Qg7BIkp909bYQ3/227IN3qnHTW+shmJ9ZC9
gPr5s36FAqAHrcqNY8/Igx73e7z9splYzh3MU9nR4W0v+hT/m0U84nxzWVmW1N0T
FWPxWSWk5KxSYiPH2fnzpH6zNi4Dq5fOPLR/dWih8y0uEnWn74kR0zaa3cYE7QU6
4qBCizkkfvPAp+HzgzTNMHz8igEJQLXlKKs4XuAZv+Zm9eCWkEt2iOjS8DiBQ+aY
Jl4+qi0KD1zL+xevCAC1dCJwow5jGS5gSHUo0VM4Tfxtfo6WI0/vKlNES0vRrbcl
VqE5Y+jYD54b8n25BpYADk1ugwPXJJ+NQiDoIw36kyuKNP3Lqd2q6Z9Wh+/d+klF
GjjYven60hQFkDi74+umvge9onFoSEt58SCbQ18Nf3gVi0pCHONvUszJtjjcLwpX
UwMZH7xFXgg7ssehDo3UxgDCgODoI8ZHN8Wm7wj4e9nvB6JWZwJoK7xT9uGtp+Ri
+66hlz0MK/B87FkjQNkNzw19HzSnBm6nTXL+bQl7/eK1461vR4Q29q8ICM2y/66a
04tVTH8fe4mkgRCFm0EmnrhNW+T2Pic05fz81D1+/W6DkSMWmAAd1JNiSvnw/Yos
1fK8YOG/TRyXwEwXC5bAlu1ZJTfbWwVg9jM+WxWaez4Itq95BDTyJneHkyNjRR0u
0Ur45nZLv/MLs/YEbhbYTp56nEur62Ee73BibsroIc0Og+OYtiNOAimvBXsBq5ba
yaBShkGoEMuuLltd6K9yp9NBQ8Vbum+n9Zm/I/NZ5GFKM3Iq96xspWCUJg7gib7n
HOSNszlBYsFEMlJZvKVJ+shCqOAa0Gf5HHhVH8+k1YE9OmH9mnUsFMgiP3A9jUHj
gW+QmfXfxExIWcDQJRzYhj1CE8oy7sRbXjX8TUR42RkfDHHEfVv+e/IMaJm9nGyB
S2k8SvHbmFfT8T5tLuWvPK83/TCqqdeqQurEgME9WrTJ6eOZNUD3f13yk+1TEfsg
6RcuaOh8N/4jGOUiCaGMIa8jNiG834KF43ZYzIprEyRgSDI169rlyi1wT3z3pHd0
F/tXx7ADkCwlP78dDQBoixVJhl7Ft0FneLv39TSDDDwGGl7jBAodJz8LyfMQnQHu
VKt2ZCA6zvD3V5lVasSBJ7wrT1omDwNqZ0ykW6cR5FtBmzhYNEdF7rk7qZa+x6A+
ep2ygg1kZCFh40SQ1+G9Q4FwNYEEBuy+mO0aQwDUNp6oCSQdlLidAfPiy12xTSxn
zEO6gmce6dO9q9STNgngli6ln3fA7cWR7gyzFBNH6sR3HkSEIJqUSFQ0uRU38+Wp
Qq4/JYtI67rqSYGGWpAjuPa5PBhVnk4BBZ1J0ZladdCqT0cIkzsbrVj0gH6/LA8A
XuTe4hD9bWUd59FPdqxIvSZdq9/87O8VCF+59KFM3ofaYN0ANaW1QdXNjSD/TO9L
/prFGEm0tUW61CdCOWSth26680M5DZw7OwdZWbMTmWeXYFBsNkON1D91mE8TnLlE
yPHBkCVKtq1cSjZHtEGKVHYmULPnVlIzocPQDOofgDGBPMu+CVrwER9kiY2BDzp8
p6okHcl3pYOEC+9b58tI5i6R+Vr+yH5xackTOsmLNM7BRHDCWzwoMmsargS/Jlrk
w2ijJZlHW4G9WHD98zMeIq4WUL+vuwhJULAvf/BRkH8trqcXd909l+mcYX0ShEsm
yVIyRSIgYNh480+Gh98Lb3ou0LlQKl0T6ErZoyaWHaAZhah3O+QYXHnlkeBAmgRe
W4J3Dv4ttsUDPL1JYXr7sTruB3c9DSPFJE+Eqy8rsAoouO27H92y8mZEu40PzLP2
cL/Wd/sIU+L0y6W3B3LwZPwZzkFElZs1J9TpKe+m1Mn/Rx98NjHzwPioT4lhh8sm
UTC1RtiIAC3MmNRKXMfALY48WcwcSMkdqEKpcuWB55O41LPADieIG4n0ejzirvPo
lzWV1v5lrlCzfuApky66RwvxSnes3q+Z+6iIKpPF/+5KFcfMOCUxJWeKKQeSYeND
yRcBvoX+cNxQXr+GiWXLWL/H4ChALv/FFMHM4y+6QFHi7xH6RgV4Q2uNwIt7PpNr
rqAJoDBM9BWGmkQijAs3N2Y9J1v7eiuIOjEjLgBTE9ABS7r00IgHR9ImMxJU8OED
ys261Hbewt7Z4dB0YhnZyLJqUOBL0zuCrypFGNSbXPZy4HxI0ffQF7RCLNixZQ2u
+qVTwkSH2twaB2YAvmy5tZXKIiDqf9BFcGBPEXSXKtHvrYkFIaW3Cc9AC+BJsqa4
iJLyGGIDj2zxNbZRavw3KPjKSRK8aRtKKuoBY+uJATKWf8s9EtIrrjQpkt2nDhIP
JI3M+WOVqDnnTCtFFepJwmesABdCeK0IIJ1osWEQcrYTht/anUujZH++c3zsu89w
Gb1pNFvnXwJFhaV1EbLPaukO34+ouY7ao9W38IN7jTNAfLXoq+8r5HJaCcW7l1JT
cs8qLiyFYkuAqEuHYYs9N0u/H46sHBSsSToP3S/GCsMBOMIRIbT12D90vi/n8n6K
viys13qDzU+qyRZeVn+oETUBVixWQfUedIL//aiQTMfnwz0A3iIcFkei5iF3bZAL
WNzVstiSQNQ99c/Ew+51gxJVxaKWeZEyZAQYikRKHMh0A/FrgsF4KZtXo788Z76m
0vSTwo0+5YwHCORbyLQDXUsE7nBt4N2nXHmLkrQIap1ZxAAihPhUv7g8HXOqabsN
+iN2AGzW4HRIv34RQAYa6GB6q/FbgMWUewTd2QHXIX4/bku/JGJ7i/ANiuA4WJfV
O6HsHW6BHuXwcCNLj4BBc8XnPacxC4QiW3hwy7b/3XgnBaeuhcwZ/cIXGbH1kVJ2
lshm0+LtK/saKWokoRSx+AL+7LoY/pk5RSlMh07ZwrgICTXKk3eqJFOzvIx+wzf2
WsjGm0nvrdgciuSX0BqvspgyvpsDISHMPAqjcIR1RknA66z+f0ubqodBEfuFneFG
2v6h0h2FTSceDu1CbJsgDhW34ZgCv+2pHtTtZP7+ROMnVusf2aqK+1x6lOgWwqME
Tx1GINbF4PaIL6BX3ZOh2zF/YUJBODAU8hzVIKQJfoj81Omip491A14vnasItBJC
h1t9zLY5GsXnwHnV8ewYoCgwc+SoUz58CILsXIsUq2JsG5L0uo5ZWhDe3ocNuthp
gMKnIJO8OQtZKry/A5WwzZAFCREcGNEYVXj68kObwOcoPXQl8Nj67Tjg4WZPVu6k
m351baAeb4UNxhN+cCkH69xR2+faX0rLUUqCZapI+BQ51b0OPGhJGiC70kwY96SB
tpH/M7vS2ONZAzLRAS8buOWkjRUHZXJ2vX0VEfcrzZYmQbsh6AwZZYDXjaN506GI
xh4+ivdQOV23p1xR1vCRPACgacIf9bGDpIhBkx4y5DvoKDH9gIEYSU7V5gwCvjMF
YePyK4EeN9Y+Z/EE+S2eYHqgYxzH4zfQdJFCgGFxp0WAFHeNgHrHiP89ZtqHQSyT
hy8NevMpkh2gqRmY1pDq/PkvQ9BiHYGuZc1K//UDGGQmQhQumAka56VIn7GoG/fI
ZvfQc4nKttE1n1LScHxGPszR1FsdqcaVybkuvIJyO3Lww/4Ca/a6OsWQmx3JgovF
rS2aSXdQD3rjMVfz829BLvl3TCNMqBwOOn8Feu9PQSixQ3669nS8HyZvtxPtR8n4
8I9DHOdqIJwrb6EW5VTugRtWg16xzTImjBtBAR5vsDAuhZWrw5A9uRG0Rdte7tzJ
qOH5h4vguDnOe047B1QDSaivm68gJjzmYRw8ZdFccCTe0ptMYEpTUoOQbhWWttHk
h5xCtotIEpSa3nRTSv+Y7pxetGdKSd/gQdYGiccOxSYxGYB9WvP6cJu22pE6AQJ9
2AmwnArCQutF43P1+iPC4wpH3aYnzZVIe3opkqC/pG9E8w/tiRNEduGZm9pcMZqX
9Eun0qYNY6sMc2hezIErRt1/7nNncUFqZkT1aG+cqATwHUFSPm02QWEEKZQynYKx
i7UA5yTKXq+C/kydzuD3z+v6kab1vcWEKs78tD5zPSBFQRI2ZrEIKYgrLs0gNC2i
O1zvMzzagbbfkIVQ+JILWTj8k1RVN5YNLwtPWYJQ9sZV+qK1ObvYtpRtT2B6raWY
mwS7kQ9HH83j4UH7R71HlWs9+VljgawG/wZvsV5eneANMtep0ygSc1Fnf7a5x/bJ
2XnAqpIEiY6ji2Zk2og5b1sAl+tP1IYOhKrOgXvti4aN5KfHQOBC/oGesVIm6NWN
4VkHd4uNQKNuDfQHXcyGUx1wxgWtco44rUWpanqpLo1abR7el83Q8ZVJE55kR+Fc
osncAs6SLmMGMcDhQtUpddGqzacZHoHUrBpwlu4IWV55wzyZBwpLI/6iEqjaq5Jc
S6bDJjPtWZQhssmEmLPTmRK0O+sIJC7D1bcahrTWpo7cUdRtzxjkuAXSQvOhCLbP
XS5vqyaeYwfjsc4mAJAtLs49MNr+UbgXEXVQHNa3qDEVyp8T7Hvw/KW7r5qIxFpJ
pbDL7s6aMTHkt+l0GNRujsaFy3vyeO7E1ibuS2aERVO/KFOICh6MDQ74qkaP+2R2
zGL+paoJHwLkLFAzlwpfU7jogHWr9xwO5Lbyz2a412EMWmTkh9EKnw/sbjyABCLB
bm1mXZR47aG7x4xHs+CotcnBHVPJzbx9098Iyq9zpInRO3/dZUn3D+Epzza8vxqb
fDWeV7QCA27xPWswCe1mYCYjQK+khgRFLgiasW8p3hxoKBslzL0yWhGgSYN6mtMC
QcCOG6N6XfD4DqYR6mO0eM8MIo94LDHtnljakKXg6mkuMD4T/1w1j9C96rJdllv+
500kAm99A0uJTQWUtK7Zp642WVo3yhNt5iW/bEGRaPV9xbFspZ+P8JYOlc8CcuDw
mDLDlKZPknZ2152xHS2JWFGwUeEdaKo9SCdPQtsYS/dJU+yOiFJfP2NThj5KbITG
Z1bbruuJ1lYitVLEJeydMap80S3xr2qX0UAieI1JcnOyHLZp/sT/ENNhgNQdeGUc
AaVdLiTgWP6HXZtMQ8rCGvEKemYT7Muaxi9NxuBXHzeC9oo8pf2NeHm2/+M4CGD/
scas9SbHH0Z8+pUuMhQ4y10zBJm+MLRV1C/uBuAQV1mDflMytpN/qEQKlqGyMVnh
G6aHOdYOmZi4hFUuIhjA4AcVhbRh8+qdiUA+0mQ7rK0nOuQm0Qfq8Z7zn+IDraTF
xs4AbmFUkJRqQFKLEOsr2Eaefh/Fw4uNU1AQJcPdEwDH7dK7ZZoNmvT2RVT3GbSv
hQRFrDGTsZY4Ysv/LkirFN1W8tURtjFh8fi4Y/IUhVwhPE48tli7O8BFRztplOmR
yboiysfnV7w5a5Jy+hZcbnPfMEp/0YSJxbYQPW47dNWmbB71z1xef7x9II+7Qt/8
WPc97GCopZxATNEo1aw2Onnq4GxT/TJjSxjwp7GfC2Xm10eTa5ZxTfn1Dde7edfB
+uHisSoDL3YpDABuGJzhdyW/6S54zz35BlbfRHg7JVDdD4nX0nhwYCjDo8+08qyh
4G4dPwS/7fDqsI0/A0qppajPp5oY6iS9dMN0kvvhJnqFEqzn58rPmOegMZDfDpyJ
NOKuVQvWeIIDxsUPd3+DzoYxYVLgl26xxVI2C/BkZMtPxWRMWvsTfnnH1HC5LIAd
kqNQDTl2cQKrsOrHGVx2OqS4oPKDJ8x796nbuGO9TXo4xioAOSNnwZz2A+l8TSq1
8AHxZcmAV21VQ3NXAG2X9h2BFcjOpuTaJFqSTp06V6IiJnLO96cCstaQJH7smfZY
wCd0GTxEUyFAH339yY7gzeHVf/NlAq8kjk3cB50ZOrKw9tIu1YHpMG3x3tq+BDnh
upxs/Zm1WIDnYc7/oCxgYOgYIcYI1h5kLxjJr45I+v8Vam6ZorLk+P3RT4OViqQa
6id2+cKk3h3glJ83PG450MP+NxiaSve7thz+MmN+8fR+qxqC2R2jOzHHqKl2OhwL
mIX6vmyemw1Fu9MI6ix4sB3pavXcDp+n4WpSuPTgoKAGMRGT270yErdQM6PXTb9R
+57EdNChprTn0cpLEDzpeXxQ1YG7GKLGI8DDrVOKhBXDvKgRSulV4h5Q+tdvfJB1
+WBlX7pb5EGRGSuoZTc3AwzlW3K7yiqc4tjTctUSZRzqeLZRJsMmHX0F+F99hYco
wZJ1AysiKOLdcxpGu0gbOYBYt49iaJz+ggoktQDASccQ7X6Arfd+wwxo9/HazTDw
eygJ5eUrTYsjy6HOyJs03fW24xrV0LM0oJcO3gahR+U3Igz1h0HOca//4d7NVz3m
rgaLmRQ/63COnoBhHJm/yOs5wk9rDLrtO4GTCR3PJ/M0bzjV7cUCE4djB050CaFn
rvBk65EujgDe+Z4m8fvNN8/22Gxt3K2V58B4JRt/TrmZhVUh1zXkAdRNI9dh0RhP
o3VXl41HGItNEcTvwO+jyJdIsZWiJUdV/cdo9E48I/+3kkyXeGOXkLqVkzGeDME/
Ex7rgHcFzLf+rDNo9sIR+nilJYQP7VY7LBbvdpJWvcKToJIlJ375SJiko4e3WluM
K0uUP+r17wv437Y7ozQWe99vX67EeC1Sh3zNkuqGLMTmK3gje3ExD1bdf71kXmEN
k6CnuqtaoOo7v7O4hctx7lRkHuDEXD1/kd4s6JYnoody5h9SncsA6aFDSqo8BuqZ
L/+lGPCzwe495zdk793dNIBIMf0BnqctAg09HTAUxJkuXDAkiWZnphMUsNcwb72C
QUiJoyHMZ+YQzX4FoPOX3o4dbvKewPhbeNguVWabOuh2UW88TpYio6c23xQhRa79
rO1D/AGZTd+SyUfQ8mlWZ5CM7rAd6xfLKVi9m0HuWs1TP122hyL6o/ESwsm/xkZA
s0FlPvh02hCWOhiQQu9PHS12d6zux3558lbj0ApsrM03PYPhgnJWw46r4pDYVcn6
hUfe7HLDJjopsDrHzZHgemQ5iUCfHrHVsNixI7ma+uEEKJ/oWFcTqMBucQco+vhR
d5XzafAF8ecZLa3bF8pdkPcxZebR3HL0pbrJuEAJjkgBER2og+jMYlbS26D9HiK0
2/TE5BZWG+77wvdlWcJYHLkiknzPU3eiuVY/BQKnB6fTlfuS2fbie8Wmr3HT30gr
2ReMWsHEDyd9zsnrUqwwoFWHgN4mSxyaq7h4lxttI8V8UnuvOWl+HFlrmJ454Y5N
iLFm6B5Lhi6AAo2Qglu6YLo6hsIoAIkUsxJUe+80kv5Mj6loA7bOdYrCyf17gSHb
mFIJXD/WJL9uqElEe23FfRTuj6bz+eGH5Z/XvvKI2ZUaEiQVlRN4k5Pi8uNuaMtD
aAmHbgmTh7JlsYWbx1m3x1Tt8j0UcAUjvRddlFr13h+mYTVyYpDyGwxi8fq/Ra+8
v9j1dK/VXU2/tESDWLuZsCfXkVJ08vsVA3SDc98IFkBiJ1kGc2kyVFTVZEzVIfsL
OjJIuBTLfvwFGaCaJC7GzRoH2plSThjn5f0nwHqp7yFAqxOB6fdEjMsz1eS06M12
4Juxv2Vhs57tWbeW5B1SlQYzF9X1bfNhnQW+60O0I3bW7WxDXBYGb3tfzu2u5Hl/
XxDmi0l580SFzcqYO/ljDoR1Sy7J2luS/jmKcrseCwkMqX9cPSlEFn1HFJdKgIgn
x8w4UkZNznkhRgd8NQ8xdeREGOc0iLtTddq9tw4gvQxe2wriIFDnBpU0r/kAWcKs
onmaix4H2ujO7BHqrnebsfDKLjeR6jlIFba6PzrtK4XTe6JMmTTuiWo5CyEHqKrI
fkwWbECHTUv37jCPP1ABlzKdn5RymTB3X3ZvC7Ge7nrGVXwQYuHt3GWMflBfbT8q
hb+YnSSfR/Yk3gqgwE73j2emgakpXfx51PDMuCnv0GUwgvmB5nxfdZclynSyJXJV
vQm+7rCNerm3gzBrukv1IjrbT60uvfP1qrydegVwB5qOf93mOp9GJRBOruaVfjf2
fk013ZxYQCCNowwamHeLpZ385EtstvkDlf9kiarb3qUAMHX1iP6HUSqtn5/ECLlg
Zx1BqlxQ6kfBsu4Hq6MVTDYki5YTNPjjZzZWcWUgGWXtlcUFAHxzkMFXha5N4xUt
QLWZ3mGzGwr1jjnO9xBN6K6aiVISdHeWxp03L/HOG2pLbPMZEuCEOKOye8iQIXGY
TCLSVGSa9PcDwpHJ2PxavCtsVUrLNanmXlYXP7oBYR84/i97MnvpMcB3TAxLIXBO
FqMV9xCQEUEtWQugdhkQZpOUxfUdJbGaJroH4tFtJBu2PMeVQkdkM9JCJcSoPmOT
2X67/AlY/my92Hp0sHqI9TYO9JgEDPakB5iRHN1HJqbkjAqdXLN+DcG7RJVSvXYR
9KBmu5dZ6qrPC92XGWPypiZlr/P0EbZC3xIZZ0UHgSnSzY1AQw8cpKMv+Ws28JCc
GrE5bmi2RKfKCDeQoaH1Rz2yk8zIOtGYYbomFx0y4zWbzUR8tKHjKWYsejNCZmrU
ETeXai0qlOkBscxnKFhJO462bhzcnwOflNkBAKnApdmcOgB3RlrsxDg3J/E02zMr
JqApnmbXi2+yue/rGvF6qa3SCuYac+PhG4aLUnT8T+NxtgG4e+3NhBAFdCh7qKoH
3eUI7WXfoqtvW0GrdrK2KXQfbjW3vWYAuot3t+6Kc7xJlGKQJx7m6eCS/jFcixwu
RP5yB8/zOHNxIxXU3XUWFgD9XHpshKir8l3TH0IQYXLRIVh9TvRi33dpAJvWuz3h
yYKeXSqvC9ByUjK7DsJazC0vJJeCHouIP0DLB/n1ghJU7ZhW0cque3/wzqGVdhMD
fZUGdGFkIfoX5UUtWwRLv9caXjzXLLwFNPcQedSOP91tNZ557pHHjEiASnIuQ38u
MEXy+ncv1QCVflxN2HZrFBckqtEEQt1lGbDZuAjPwsYIhHHaJUp/rX/bDh+K6RPa
EvJdoB478x5dFNARXG1Fbv9b9aw4Qj9YhOwFwEGKnjH7G/9PfSSbL1BRegJ/qGMT
daeXw+sDR9Dvxfj8xAZLYCKj4mbq2l0e0InQtevaUVwEQ1+WmzhLxfSvtTh1Uj+5
zlZ+NxXSTBLJEnbAZG7ae4uktbMUapuN0J1ziZ5brzLgWSphN+Y2rcYycobjMk4Y
+Jl3cOKVSjP0cV3CBX/iTFC+vnrA6RcGm50+AXRs8SakgfivTzEzkjRhA1W5t9rT
f//ysbD9pbDwlpa0vNoaCQ9wFiEOz4kPmXda9pOqG+IViPKsFt29dhVxdIw9WuvP
7CDjpA6BP/AsTW+NXOd2ZIEnJ1jMuCEDzEW92dULGPjFN7JTi+vvaEpt1HwrYII+
YEf8A8Q8ExPmmaPMdSKos9t2ovkK6RKkYv0sos8Wjg4+cAFGNMPAlEFWYpS3g8lH
XtH1ADSwaPEzWkEH5gklrAYZF6iVmecx5ba8KhaPd/6I0CuNenP0wCYV328LSt2S
DSl9ECT9tAlSvIu6vpEGGcfWrt2qFmCJncqhVZ4x/+RBYVblLpHTVSSqp73Jx16R
Nue1vExDYP6E5E6QrKuiCnqZU6vVg0qPqOJhay6KyWiHWrOOPnkCkLXXYZ/CS91i
M2Xc1HqZcWlJy7O1Kwq14dPaemmlHkbHlc0ZQBGPvFRWQYhgkArowV58u6cm9Klc
coHRkEba+7yI84zgVHE9Xfjq6FBRxfWuifOhGh9Z7/Dc82o0zntETq984D22+4J/
BeFXUsjvisLyf+HfHKvfxjvSCGJP1jWVPtDmyoP91Z1DTDrL3IMCzswYcRYG0vDu
+fnTUU5L+cO7o14u7D7uIYfb29b/OB+P2eEVn3J4DdxVx1nuhWjdPeKEv8vpUmCo
AvdiH+ZyJ1d8ZLOUqMgJiKGi5WK7TolE8qvP8JtCO8udRMbv+DecGlEci/MqMhAg
/kjsPnl5/1NBZY5bJUxvQnrrmhvQ6TfgjEqvzVnFUHLP/R4zYBlkOxec7PFW1CiS
DrJ8vzQWHdUPPzSbudSoRDbFeNOAIhoQFTql9koJS7rE/nGivw9O0jxm0eN4CgHl
9IVn50fK7Ql67oiZVNASTl+2n7mcxijJ1pFOLcYRXXGYCESFWSVGq2bA0E4DLrNC
agXl1f+wXNAowkBx9sn+WGNBAfsfC+f7R/H44Tcs3vn+7OW7McYINXAflrdCtJx6
tZ/z8C7ZVI0cRVdujG3D+EIVjGye7DAb2EcRp4JXKXnhEv1nHYBY/Thnr7aeH1zs
xm4HSeNFtcGVkTKsySXPBTVgZEOPZVkJMBu+SpKW7bvZccWzIJxreOMR2prKgDsH
6g17UuO/wrPt8E4MP83i8tIkZh23HfOotLeg38r4CjwdyTSFlkvKILmzCv0bwYvn
/JdjWVmB6XApRhy8zu0VzdxjGW7paRRkFYStRLFq3ovRMMca2yF2LIGi8PTshVlo
m9FmjIwpM+lukjJQr1n8nBnfhWMYLLMtJynsibJR069hsUCHQB7hnIdKqsnHBtcf
I+nEeyH3tGb4+I1O1gv02JboeoQ55qWrA0CKmT/cl9d9XCOX8CGBt46NyIQRWAHH
zvZdG8Hl5wnG3Y9ihi6NcSDIqck2ewlaREnxjN/dBQLcO9GwvRMMqYw1W9BeLpOH
v9Un6phPTqsNXdYxeR1d6YUHDqbKteZvvciBHYqYS7G4231K5CS6JTQHT+bef0bC
9rcEdu8gHWtCyOmgt66RqAkz9f30j4GQ2Q7qWKp5N9PxJpMUmIRICXuiWcw5PE5y
IB5Vr80Z2Km5VT/HJfbpK0L8hTaw9rwjQ3V6KpwuQ0CHJZeQ6RWea7khCJRvJyh5
zHDA+kLz8b8f3jpboo5/SHK+NvAddS0Tp0k53rY6yY5t2BroIQa+Avg2SMo5WAjO
Mm6cWyS6rZEgKpy+5ZDQcUia91oshla5qVk1CD14r4WokTko1kZZuaO8F3tLLAZ+
XH+qd+ubHkOZbclJgxBu5HFSy9Pgf5ETQM81EiMFwSMZH3XWud1KMWuEB5nRqQ4I
bL7lOKtbX5h6Z1erqHMF42UIfk0Mcq/OoqIRTuqgcKfzBowXCxhUGBimKbTfqCMs
XoTU0UgtcBb3q1cveaxF3SgK/Gw+U4H5IGgOfpiZktE/9ooT66PesZ8QpCCtB/fC
ilm53N/g0UvsJBjUdr7pWqREm/pvWeICJ2YUf2uWlse69B13a1b9aW0EzmL0Es6r
j/q39lLQlnuufKXTISIyYZ3S1R3qiRDPe6Kdafho+Mv46bsXiOkt+wDMzy5OqA5v
a27MUqacsFBaxK1wsqvrVTkUqtkWpI7wgOHAKwlZB4jOHAXoAx2dD58Kg4o9b+K5
AclUvq4ZK767aK2/JZAVaT6Q7ApNz1e8vYanpl1dRfsLIYRZKjkvt9fe4AgPbuzC
cExAAooT+N0O8mi/Ex7keolu77WdMDjUlM0S2P5aYqJWEX7GdjWpNqMqMOf7+UZ9
07XfaTYDhBE9FHwqyVL4ldS4m3fUeb84JiJMvXAEGCT6ZkqNHBQnBpBIyuumKiwk
XsCnXecDeSICgOSU09jOkKSHJ9tm59CztoBiVuMq9Ag5sSHZcxgt+knrCmCsBK7M
cPak7lFqGvti8kZS2fpAPB1axn6yZGhEwHnUXrcqdRmuVKZ3AUM6xGjERTBuXrq1
HCNH/+kRgZGeOBkPERfLRj13rgjS9dDT5jpikMj/s/q8uaeB6YUEN/RnMX1ciRlP
aPdW1bdaDbcavmp+drDAJp7HWVEDEbfCX5/LKPhzU4smIaJncQRdyCcM+4aax3zO
g9nlhZzCGHNdtZEi8GjFZem9nzS8QbJ8mhos9wwwaBb3HoAJiwB+4bPezXMAZtIT
04MslZHS6Utf0+fb3EAU/HMI5tlIdqSiWdrA8EOZhrJnQ2RNZEieWmpu1ecXBQGi
16U3qb8HcpLspQ2APbRvtv0qI5bhNdj+rV49LhL4L+0IOzDS0pHaWWZ6eAJZzfP5
4U3gQCPIz8jA4hQcAXA4SvCV0Fcpmm6tA2Z5A7mIM9xgse5qzyQHt2/qCBArVMxi
fwVMFduxL2TwF5YwZ15evAU39y6pecuJRe8E8r8UCAg/JxSgu3gZqyvuqKc8BDqI
cpLKwZBGvYrXyfpcPHkvtSuaov/JOc1Vk7Eu929LP899rgnrCs+1zRL/4ATqH+og
VdtV3+hKk/uFaP1ApUDlWr9dfiDyMlnhAhQlD5TJ3Sn1uU5H0Ga3D0zwDeZ04sk1
005c/izLp2BcyEL9xNmDH01LGUz6YujKEuIqerXDKozUpuxqCkZ1Fdojs4V8KLft
90FyoTQqaBNuJZm5offGQ3pQMhPuHIOT/IwWKkBQpfz4jwns3h8HZUjXssr4Vu/g
gTDO7OxLkrnrfos0aBo60x5enjl/VSuitqjjJfbXz77RGG9YkiD19pkJrIxyJ+eB
8NmKpe0YM+K+dy6PVAaaas/b4tFCZzknGEWQUT9ESwB3vi7kFt3SD+DxBTUa7ava
/PzrDMBFN/AQ3aJdZJHRaYeZmWrFh9AuV/v6m2C4i2w/B/sIHzjqbQoY8+/cgzmR
Bxwxe3ws4o3mzuph+/XX3DGWo4u4ThyKQupi5M2qHS4bYK19VsNF94n0ytsb+64E
PNmU3AkoIcHlhz2GPN24Yyowya6M3n1dKity1TfX9+KIRq7hdxEYj5WbCPoTzhtA
NOiPVfyp6WmTmk43ArN9qDoJ/nCoM7zkvwxqH7iAH0QJj4F+8lmvdSRheH9yIouB
G+2io2TDIaik67aoQEGxDI6jMZFKQaf/bg4e2GD1cdkcJYIvnzTU0YDhrh3MgMtV
FlEG+zQbYkPZWB9nLKF18SHlF8oK00G0cfG6jsDBVzquO8o1zmwdcbMBE6nax1Q4
ADJrLsKygH7mqlNTBqSSmiZzAbNvx24vByHReQBn4Ka7MFjoVValKjofsf8EAsFU
Js1Bful3p9+MwHP+3XEzzmKDhNINYyqiMqIeLtvPXmlQ1Y5pPSpHkk7q3yQYLIn3
cPt7Q7GxvMi+ew5i3dThpQMLdLZCtApNAPibBDIF6Y7ja2RulUJSjREX7nxLAvaY
C8B85bowXneaUtNKpt26CNxt7C1UpZUwFn1AKWGKl9MaO/eSs7hvJQ/4UUfXKJhP
luC3DtUTzuxQs2vKKP5HRt/76xT69urHK96XM9gz0YvGwRRgqJE9QFn1Pk48PHdo
6WVoWq6gCBfdzgnfP/nBQVvPD7hMpNv7OaAxYEao9lkfWcLq5cyQ9eFgLRv2t1R6
0KsZLoja9awIrtVrTXco81Lv/cEoGTGPyCpXE4+OD+Bh0WpUoBya/CSw8AAXK0QC
wnsshATTplBtxBDswbEgwKT35EJbQ/tEq0ZuvVBsSxQ+BnfBf+PvTOYNYIxPhjOE
JoF98FeNY8OnsMrj7wOPTTsJO7cz53LqFHPGjePTZ1SOIBxHF3g9T6K0U6pLLhcA
sfPHNK9n5YwmeSWashtxYWM5gzM14Okx08WTvc/hCDTsyLtNhL6/dOvtdvR6cYND
aEGAyJfoWIFzbrKTB54idsoSM+L+Um68+o1mjjYDIX1pQiNZQdCoUJAHFm8kRpF4
Hm4rvx1CSiikJpNjZNip8rE959P9AC9FclV9axziihd3vEfHDIGSZKBPXtdGKoyB
Y7bgWQocg4L7/nGrJa0TUwwDPpuCzDGdas5WCljxEibDi1x9jXfuYGCkgowAM8lV
2ytSvcUAx00ScJTr0JFLdtep7Z8WE9+tZEBweauXhmr2Z8lYIpkhgcp3oBetyQJE
BqNL8J9BKUV/ZbfKrCs9frQTjCK+nymhTzWQWpDoQWtQmeWHWSHnj8gdKDzZjNPA
2iAusaz5BlSL0dPbggFCtqByPhrFy4kUG/mTWFwbMSfSXQbIAJXbCi3uj22rWyai
WUcBantrcHWTJ/1acsuViBUdI/Ya3u9QSQtqWKCKSvLsyhDLSpfYIIYu21Jj9Zay
xrDZCzeSAAVEVqBMUdC53wSThKiAf01IaEyVTq9eFBY5YOcr5Kgm6hiSlZNrguu7
L74YIlzUYI9+naVx8qX4pR6oEvT17ryXCgfmq05hV6ubAOWkdW/VNCWCmb8V4Ldm
XYGweyyZ8w9zPe7gJEsPHOOJxSvz0xtzGwpHEKOIQgJNx8I+P+luzs3TtmCj9/Ir
Jf1AdfO08o8QDUGSh5QFk7IoNOV/H9V4PPEziIxb2u7M/vZGd7M/YMWpFQl1AyD8
1G8o4l2uLLnSS8KJ6IxfcPFxI8ZwHUF97tpGqjfid3/z7zJ4xRgLadDM5P2rqmNI
oDI5QVGrQGSxf+CUMNplvQTMIOejLe6wj8FSfm8a2d1AVCdvTEyoDukBw4nUlxv8
ovlT6YK8U3y1Og+9oFTcoe2g+rml8+F5HyGTiu7Pxbu52muIM1LFoXcn9nbHCcvS
IGiibJT3eynEqSlKhIjlpulZ5k0ugWLQOIlmpEyAmzwo6vgKvdWtPwiw3fBhZWIg
tYm8cxMJj/aZKaVPHRzhhWkmtiswUVTVMWVfk8/lYFpz82G2xSGGTP6zfNY62K0p
GnNAChEls47Ppe05iS+vPZuIjuc6KVtLbBuMWHXIzDc9LdVCliXahg+6FmDSv6xj
TxZQoU8nqk2uZqTn9WZWS98R4fAO4k1Ug1OWoqBwyXAE1ZC+9Fxk25UHDuvcKwiT
fkpe8127RWT+dE87Ui7kftaS4TSLRvSZJ3qQw3BO/VDg8mvotU2BMpGHap2DMLCa
31LWoBkRoSKO+s9VVla2xqOvbMCfWRXsoQ/RY4S4M479p+gFhOcI9n12TtDVVgmB
xABr9+zPlKex4azel6g0YG0ffm6mCyZpvZlC/mpBiNB9aEiAr24xarHer1d9XZAJ
oAuTHlUzzlxQ5wcbiMMratd9tE8fnxM6uYrHFONQB8PPrFNPmFJb+tf0LQEGDaFB
tFt+0inStou7l1UBxfuJXr/b6mLb0NMZFvakD/nfcdwfY1JXWFqL7SrRpeHB0Ief
77P0MEa96DAR9aiav83XQr71EODnyIEKzq6JmMHU0S/FXQ3eoZAgp8NlPNShkwUN
ZlEhpLfeDaQc/DEec+U20lY9/sU/PmiMUoshm4FdyUK+PwN3p67gpt+ko2o5wJOx
UgnERNLU5VjXpXMUBr3xn3y8yuNAwzV7rihi2gS7klg2HW0h0aX8H0Tt+gADZz6K
kTlPIzeYd7OYrOit8DOvKnFt0R7DEtw/V3gD+EWx8cZP7swVGqTYgiALibI//LpA
fp1u1uYMsMd5CDyOPGTqif9OuH/oDj+MSPpUIguuJBd78deTba93x53lTeryGgMh
smsvxcQex96lCQAx4CZNwy4cbJE2O7PfVSX6t5aDfQ3fEQ8xL5j6S0tdC9uwwlvn
ZLGlMsV2A7WKHEDIgpQ2b7iR2Qhsf0tChckNUhDV3MvvI94wcsgFET38/DnSNEZS
oQ3GTmH5pGYoTK/FUOII05T7repfOHJq5uZ6dcUg3+/MVZ5veb4mxYCz+LTtg0iJ
K/xj6bYh2GFyj8u+sIjd4UIIYkdctxj/FgaY3Xpo5K9RLdO7Zq35kpWifzIlEg5Y
XqJmiX10IevSoIY08qMvxmjbNpToOoZHc3azbfJzeGj35/I+3LHNsUSNr/q9ypA/
6coq0jBGa3BA0gIWpu8RD4SB53ibX45j6PX2trYCYPsDkAuecxRTLVHxPSPJGmR1
WWGUPyERUU55382DxPcIbpIfQmBYEn7U80KP9UwK0echcNmwIBiDgjvCV5fzAmoE
s5kdfTdf5kmzwkdkdeMWFl6hw0uhDLRFdXtigwvjdYcOa8mxpCwAg7n27TzqoqjR
LctS2P4akhhw4RXTYYEQC3NQ7xgAr/r2To/jb6YypNajKTL+VJr69BfgzOKpr+7I
btDbkpAXKQjAdQHGj0QXYKtPHX3cSFYW4+TVLLVTYn6aWsdC7q1oq26oHnR1QhZN
5uzBg1Sfh9WaUxjxow+GeBF7gM/Doy4RVGPtgh7M3swJnPEii/9kyw5Cp0fifEN8
wzzvukc3n0veeJwD/aDhAwXra1VDf+tR44as9EkP4EnjU5fgID1rtppZ/345dpPM
VyVaVA1bhI3Gt5MJ7+yX5yCHLPcg0Gvh832C6GGz221t+FgEoZtDfNGhTNWtdgsW
LpZzqLmbiTwulpTZy6FXtq62Z8UitkCQvuzWlK1F17OgR+0vTmY0fgsjCXno4nLO
1ss5RGxLjrt87MzsO6vOypcoG/OA4Wlh0N+KwtsARgAQxxEFIK2WjBDFVO2Vpx6A
T4WF49mQM2B6ffedsdnBLq5cu9vJBVfjcYb9F6YknR+w7EMoQIEu27kYPXCBu5mP
vLzSNz9HSbasXYtevPhkrr95zNg61DOUfTNO8ccqDnJiOjbNNpX3BCLPrCM24/Jd
+gCnG/qRz8VZdQevlzlK7mqXIrSAA9CHK1h4vMiNebolfFPePYYC/+HluctaaD1n
loIGbsFFafSTogTwPb8IhXBlrwluXG3lLbfD//ZKjXmyzyCqr3pJkU1Sa5qzm0s8
/FdDDW0vwgst3CtwUsRAogboGHb8I/sX5Yw1JbCKFGNNnBkyElZcCEVulvltWM9u
80dz1CnxjZtYau3y4KQv4G55bO8D1Pk/DgQ15PfypnewKfbzG+l+HKLtzzc0fmgi
M72ACaVHCFC1q83EqG9pdiaZ/QvDzYM6cm7MvhXCfIYroOAczCiukc6CsZFFIplK
WTCT9nQNObp9UtPPt0CiqOU0TRnv0CiCXnmre2Z15aPSLDax2ZFpkzdit/c/ENm5
WuRUqcF84NcTnqclNcoQaIIT5Ue1ZIw8POb6Kq3BMvj6cfRqnRmJjkTzcPVACJys
HXH1RWM62l/PItKE8npd7B+xMope0/WsLp41T2QGGMJZTw7tt4A6NXv26mlNqCS1
TWalP8QdEehBuT5+7OSYlFsEOZnXGTsfqhKPxjR0lLJ3EcmYoGVTVV1egsqqYWew
zGgz6y2X4v1aqdx476e1zhJPSAUdSw43vTaIJRYpAqs36FGFqp9xXxRh3PDJLMke
Z+JbUVltS3KuDPTG3tdpV+F8msnOKFWa85KCAtCIGWGRV1f2/LWwdyoN85s3Hzr5
6k9Wu+ZGMiwkEjrdxgpDoIkk5Q0ftZ43n1wg+9lU3wq6n07nYxjyo6i6z7aarMIx
L/UCkR0mjZnmKQQfO9hGzBE666zKfaq3cA2NK7O/T3ewU+Ni+LlQInU/48CgTCxv
eIiUR0+WZ7fmK4qXUJDbWiEaxvg/Wgw0JsHQTtVEciHdYpjRJXi5Jbt6FfJHRIHS
4z44+/xl8XQxKkZRlJXd+7noW1UfeU8jZtx2zQTErO3J0XM1KWqLz035q0TFyGIC
IEGGkyzjxQnxW7G8w+a2idxIJ8G+68sH+nlTM9wdrPHQjADFbwHwASXwqybSokhx
kPaATlR5Y0dTM9jS7f7VkHgpassY1hew8YNP9WPvBjpWrKx9ALDHSZ0TfVp8dWqm
JzmeqEMq7Ur5IkzZwp8ZuTJHGG+fDoIGCuDS2Rn30rh6aqMXkIiYP5PJ7w04e3KO
jqu44NQHZljnZMahabr+/Fkd9+BONUBmdBpjQHBJN7Q5hd3XdXPp1RgyXvqqpdFm
ldeRaRhWyaIKLoCpgZesVSlC0uEj7esJCJSS8jleQmzFG2tHiVYXypnbcoRnYMg4
C1SIGs1lY+HzVJ4NVsVZiGc6LMhC9asdSwGUkg+OgvUEGd3Sy7vJblPKbb4WMdQq
zK7wPV2PGKvn2WGt14RNbLxZ5fR2N23n26bug2ubtC4srI4QXNEdW0vbSlylte2w
rMMbzY/03oBwpVy4qlPR6tKnIINRdmHUx5muU5RQxCNNhrWDxCmVLCUexxzRGhv7
9xWSZeNBhVelACQLszlJB43WF8gG+gmfy4o8AaBbgvJmE7T3QVF8I8us50QOa/8J
GKqBVrhM7PPvUBLtRydX2jIvDoPXIjA3tedZZXWyFPT/TeWzvVhhCNiFArz2PZoE
TiukC6lKMPjIfpzEZ90ldgDmNwRohcB1+R3P4QLSI2OKUcGxI5MOlRmX30Nx80to
H6rho+y+9opiJM0pkktDMYhqbQUFKl7N/hNGRwXeVFKMg7G98rLDEhoje9GEjO6x
shIWNb7PJpygBTcZd2gXUUv9aWBg99kY8D3jedmql8oPici9cVqyIlhKtgDNV//D
P4rxGcRpZ8kXOJLqJJkbGddQ41/vxq0KovIJ5u/ffR3nZczZIcz2WwELSxFvHYLj
VoRS7PKVYkY0a8vYMq6+iO5X9NSAtEzOMVGMp6yvXvR35Pgo2KG/h2pgf6M2WA0g
f6aIJshjz5IiguwbXaLzsrc4Ftep2TnVYjOS9frUGE30HFFXkeXem/ZAwjCgl4UI
Y8sgyOFyOgIffV1V5xcLt1tF0jo2rCJGEoCuplFzJ8Z5OUmN6/tcG6jtjaT2ySex
uDg0yqMOtwC/lHe2fHPeWyZscTKEe+45GIEm/FGIKGXFEedis3Bk3KueUrSxT1+/
NmL9pK2y8WfJnJ2nq+A4VCeSEFQAjVfJOJQpd0VO6FMvQUvIKFqkZTUEmfHaLKf+
hshWO168St3f33yuSUG/QFoeAkU7u7xdGegGsMhzcN3PKHoJTsOu66BarPtc02xm
zZb6vp37qpQSpMdO1kuA+CeAjJl74huImXQXVNlrFyMoX1Ry1vuCE5Zds1pck0D/
bdwlP8zlqPvuccYi1nWd2RD7ZzoqoekbQObDRenFXZhOqLyrJkYb356J+ksCdQtE
Eo+h59alWKlF7IxGRjv98d/r2KkgBExCx77m4LMfkEcnle+YhPZVsb7QxQWE4Cr2
jpOFg207gCGF8sAucAH56uRsqSxyYDVuszQbePJog83nsAXC+xxQCUKqqmAYPktw
P5yCD8wcn9ejl4Bxty8aJQUfQPH7jVDv8fEUbKax48P4vwJByg18dsvMypFlG+x4
udGDlOSv2MoCpl+0iyhdPR8FJ1OCQhIdXw6z2YUsaEt7iHeeAjddZnVVFpTMMEe4
oGrL+LxyWR8TvQ1L3nU6/vAfQiY1+WP5g64upQ/f9IJ3j6xixL/EV6GnUcW0tJ60
7h3dCSYQT+uXgsbsc0svpng+twV60uv5bXEFiERH5klZXtWTZOmgqeTIbKcKSatT
ktArW+NZJa9vI+kuLbAgWIASBIJzNt7jJq7fw7uzGk5j5UE+SLKD/TIH7ufkZ0F3
t4VUUQqFaQeu1rY6EBDLHKneuDTM8mBkHgz984cZcIZPPqnAhWFpAKPwhwx0V+dO
X4BbfGuLb0wWRkb3DtoM4OpokqnyY2qsGg86/Tp9waGNg8KtyXmmadVJD2cgOw7I
xcexOdj3TZekGPOr0lDnVjxoYmhvXH7sxxi+wiMKBNhZgucK6CX+ySB1eJxeQjND
ixxe7k6PtqLjCkk4IK2PPqsAyksIcbzlmKUgjmrJUfWcFP1TSyQJjIEfOM50OW0L
p2Ehf2L66mX6c+B3crGyopfA6XoIpdc4lc8jSceyzHOIHirdY6UCZYCRhJ4ccZWi
EzBVqlX+RBblKafEQIHBoNXBZGyHRLwBKHx0t/3JP/Y3xCCUQm0kr5s/SrVGszox
b8S0E05Hg2pNnC7f3oH8rNhJ2pPZN17jyguP6FgC38BWC8jw0/ACcxOY70XiD2X4
rGsuIn0WYRzoppjukjymICs67iq2rIiT+oP+sRx9nE0CLFh+SblaYrAd7MDklr5q
9WIbAVWlxaVT3uG2Trz2DFeaOgnsWiwIk7ve/C0pGRBm+sdWpU54cu6O5EVo4PE0
6DERH1kukYfITMcjw3QZLVBQtNMf8Oz5b7a75IitYirAl3JfFTZ/lDqZeG/qSMBl
ECVoQ+DJsPYsymfBMLyP/uWMN+8xTHywYkAPDVUTgptURAYsShYX/dY5fJzGsPFp
Jn+L0dov7GbfQ1zsmeJyJE9IeNiIyh6PS4OAqXlg4HFmctDIFffIASx47NLV1L33
Lax8JU/hY5m2wwmyqINYLd1JbzaeRJS9ZhpW9Bo8Nmz2CDYzuSG9N9BCfxrA4jsR
mI4Q1VL2EPZgkvM9rDJy2vP/COszpqe++RmWpFRNvVpZ5lqqDD2vp5mt1Yty8uxB
RFHBdBpTN94w3FHApACTufvsT362CJQv01q5KKwr/qqX2qgSg8RpfhmNarA5LIQg
0+4yCDdYtTrAFBmPd5mm17tl3Jy7lkdTi2LouPVMwdx4Dqye6pmh88X1JllFt1fg
TGPgcC9bzXk4cYvnfAAoj1Vhx+aeRld1zPsFEqfx0RVsPaYHC30JHSiwH35cPhir
IFseVT0YSciXz+m5Qaoxurkocwv7FoArB5Iv5Um3GTLM3ncfDnxVCRpDfXDHfPr3
3OnXndFaFQ+Y2h/g6BbtG5wbeN6YJEUtkJ6lDk9e2hoBN1r3pbjWeGQNZ9yY8kOY
NNG333Td58e/FsE8AAxqiZ89f5z/ZQlbu4gBi0Qtya4uy8cA8Pfez4mf4QrJHnwC
Ivioy4PhjyZwq2IQAvcg8F8jqCRLEjjDBgDlWlls0uQFgWKyERWfVCukTQ+1vK59
8hSScd8i5TiW90JVTL9zILcKhFXXCliSirb6TBSPJDjAPkTvasTPUfz98H/dMgAX
Q7JykF0XYyUWKVRdLxK31SJvcH4h0r5Vj9SConFW8vwnzkZYa6l9tuarsBXhSeMt
jeHVlsqpjJl1G2fcPRmDtM3QMBJ/guQovJaafGJ/2rrLY65233odRETeB4jk8sIP
BGbbJZ9K6pOTr68AlG6m2xmdwK6aOxWO4K4MShrrdHF1ZYCmGjhPPyIZx7Wd4r2e
39qB3Fj+WiAy7wqvsP7heg/VX1BefmlRpENimOQ0NS35NuJiBQJH0hDQB/bG08EN
wsbjYxFZiYFVe3DmfkhELqJq+zEHtixHusORoFOT6dG7/E7Pv3xwqzECeL52IgEC
ttMED9oxRKBM1B62hYlqCxqI54gF/NqgN6BSL1cI++PeRZ/HR3bt16olO2oGuay5
OFQL9kHztAcxwDegc+Z7ureUXM/8TplC2KRkPwCjjNJ9BEEr+EGZbfJICteW1yGL
0u33bYnSEE5QtjVliAiyGKWU/7NuZJltTKB2BrQ4TomtpoVbzfSLNQLkyBuUFgh6
t08IcbmZJiVREkHJuFM/w5jS30WhYGWb21q5Ib9S74RrxHDVqOvmmbjLFIgmnQ6/
ibzlbui25HaVDSFsTMEHc7aynLZpCQ77AVb5zZ4UL160JZ+OegXwDnULnhhxuWwR
FJHId7WuU7Wk2yKLRztoxOtQ1vpObpsjHtTZMgoeT3PCTctt5s8vtaXGqtcpR2lh
L/94A0KFVQDbnVYjHdAn1C8sSK2gH5UaaZGHDLq80CEhWIbbarZq5oIQA6CJw99d
Zgd1JjgrBMqw9mTtXB9DnQUfE+cm/PFU0BB0LlA0nut9+3Dsm7/ybWlPiqAeF8pQ
cTI5I6T12faj5ZucTayZfNxHl8x56x0eKv8nEEQCNFuubLRKArpbm0u4sjJZPbt8
0/daSRAFnjlSBtrdOQkTosyu8dyNqHLY0vXRCQdATbKALEGJEJJiIHuQCr+hGvNM
fYKpQt4JSvWtYs3culBE1dvislGVaRpJcvvzfGAjCZ96jqANoaSuiNQ+NyOU2Osr
rLbuOFqMvMJ7b1Qd7R05qytAHm6zpFBl+0xKU0uxEJw2EGXsCl5lQ/aYMK1Cor+6
+7+/rAboVD+Tydv8o2OqD7r/o5slDP9nhR0yyKGsLcIacimHwM3nBETjEK72ynit
wj2GDEkmoQ5HqPhvmGiZ3Pqe7EKB7vNgviYOoc6SEhYVrLQhlPyq9ToDZfzVfX0y
KtPEw6BT6hshgGY7tU/LZ2mE63QXKREkojH6o/N00bXjS4oUNcUu/DKiNaP7U4l0
ZbV5UPNtgArP9fyLcZz0dTVdPwNzJ0ra+dF/mhxKH0zm7JRgUPV6C7xjeD/qlbg7
7tF4sGZsnK+IgU+a5xP4GZq4oMF3bhcWSI4BqtX87RqaQ7nBJVCi8COTMpJZJ79o
J8WOe0K7AXTEQXyZ9XSQi1xRXu1H7bgLan4EqLLJ5nCHvXT7TG5FjfAd7aGVAOoa
EHzrun2F9zWbomgRB8x4M+1EqSMBwtxjjTZnI56O5NdviTNp2+m0+lUVEQadL7wR
XqH6CzbVnz2jjbUz129aWzDt8Cbe5X0k2TwA+sU+LtRcOJzLODpo9MPE5VEof/vB
OeB+MQ5u6IVa3S2VjPKuu5P0qMwQgslxSrMc49fOFTEdtIcaFlcwQeJsBF3y8ky0
df3+4ayFufpilEjUdlLsOCdPs30DUUEBGHzIFemZKbTlWw8LSHQrqbmoCU2u9CaB
vBLA/3ZrcuyNrmUPxlMkxQM2vEQYex7ODQHNBXSF4L0ReiiFBjZpd7wrnLkVDK5L
+E0CkzevTaUNP8kFe+70IpqTW+KvL1MU3/xiUxK352fPK20eNQYGzjBagwzVQFRw
4hNkYFJu3v8o8bxw1+G6kgvN3X4XmkaxlMCAysf7pO/CY0OP8i2KW4Kkoud+F+HH
MoRuX9shZ+iK8F5w74plPxE/gkwIj8daULpawm/17H7rctHiAI1dbkANCJ5GnpRF
YNcoQH/9wwEWUjUuOyZ+iN0cmAu9YHsVEZVZrxq3BIcKGaeSw2SiREiEYK2H1Cwz
NSsa8pwJrSsfDB3e5xwa9IahF8wYf1p02/HlYx8tYVTaUCSAQRTuwBkqbc8bMkNA
zTkv5kVhjMkgMtV02IgrStYnRuhUipxpZbTpXOLRcojpsq2hqJ98WmHMUZY+10L+
rMxxKIKYw5c3/ud4E3nQBuUDw6I42Kyf/gCS8QvlGblp6LARLuXMYeMxvVYcuYQP
188OrVKUBgfc0vJriTuwRN6PNcNeOqYVH+G98GR2eJtpOkRx9CYksx8z05Mritbw
M2ryKCN0jry5h1k9yY1mT2BAce61P30L1jcxmj1XJoL7DZv6VUkL+7SwO5ZyaTqZ
jT3B+zsgWwCGbuGSGfmIPtt9zsjyn7gnwdHCHDbgX3JhRrfeh0Jssz4+aMAlOhrz
UblvksI1SHUcJ+gzyCeLEf+HWRNHsITtpLcdEQL3Uzs1guro6UEuyqvUsjFGlNfV
vgxoZ5/n3Da+OYnQld7RQDeeT1l2CFpPrZRa9oKw1osKbj7KUrT9pfeM1mN+wgRP
8y2dTVt7k7OjoUPOpPYTYvcg9NLpyKbldmHf2sS2E+t/VtH3QUviUSE8AGRLHdjD
dKUb7BQ1c1bEEKluaWqnesdbPO1fG7+tZGo7pwiMY0cAcdNwPxS2BVa6BdYnae8w
jTgfpafr0CfuTOGZA/bzCniRn52p0qLanAfK0vzT2oQx+dQ6xs0rICFM+tJEaSCh
Pf9PejudfOQ9OdKwuExay21IvqbayHZIZTpx1D2tK9biSDENTZ4Fs9aINwjw57s/
oc2tRmdowtpVpMIUxTM2vYOv6OMb0/a3TKqn1Ow8kEXvuYupMVn0q2B8dLXhqKOc
tvVr2rxHvxJAd2GrFfbB1aDre2C4SsOTYuDgT8g6UzsAo22VrcUUsXS8PDkBQ0n/
hSv06H90utlLqvQ4lAAVm1XwWKn0VieVgcksDHAcm9acyFgRo5QcWCm2m8MLBM/3
lXkEzuseGMUXSJq2c4mXOVcoxhh8CElrVJxamhCA8MhaVCIPYrN29IQVwK3/UPcy
91NLcl0PrGTqXmA3G3Bkly7qlSfWCTaak496Gh4LFZ3J5i+FRJHFzg7pAFYlemT+
PMOzaeqor2kusmqTNpFdam2o7/hzs6q351sQhC4vMBknkWpbKu22c5CDIb76J5kT
7w+VfR2w0/+srZird77eaT4xoLyvsMqyVCsAoXf3MbBXpiSRoHvhb5bySzms3EkU
+MdIS2uhbOQVwBKH0GsDtnDBpA2eJ/ZnpsVdBYhhgsY8PP7xzJ3gUzZNKHlQ/lUF
tpUau8HBkipJU6mQ4dUhgjF7Yn1Zshp0LhtdsFGeYqqF/AXWyaT5f5R2jliZy4WU
98C9s8QP+CIdL+zivYK++Lv9X2R5S2KmrAAbXJk/uHBkl7KbM3qxetzkObibrw4i
HgmSx4p0+CdrLwnjaxopUZ5//pGCfgmviMX+OAnRjSNvdI6v7KKg0TJSNucKyi/9
PPTpvoNLd92w/k9+mTa+IlaGMbGar3HbczSHnHl4A/kOAzjYOSHCLC3mVGXocFXg
NyLauceGWLGBTXrWPX5qVmT+ppnrQl+vwM5xvunmn4X6VoBSCuhJDnhq49wqL2BX
4Wx30iQuFvJy09Aw/XhXqjKaG6zIaSdJOMWpq433JYxvod47EvFZ9kNdPyh2aPLw
/OXmCwhIA9zxyEl6Ix3HtVTN0Sbhq2VBPFjhlwLNKCtJ+JIKI9UgGyl+gMI8jBYU
NJkyLLOQTKr8XriidmlSzRm3sejySkp7k8pKNh4PJXYozlwpqLFqIyQUUWv63jWR
V51KLfrprvDwtagIxV1NGuL/ct4n1K+beBhaUXpn1gt0lF5VKtjJj0wZYSlPvRHL
fFrFC+8qwsc0bsFkwtWHVl6Jqabs/vWCcF0ItnmCj4y1uJjmjmTTJ7uU67F00KF2
+J0oNo8U9sBUskix+puNzxQ/hPcRHzboZa9sCHxyX3WKqPwI5NacPPplviODJMgL
rCIwyzBYDOVbjePLG+QcXJCcHAfia+8Z4Gty5KsoPqdmp3gzfjZlcMRI+Y1A0CIT
xCXD6WwN5sxUoTJqh/AaT4/9oLI2y3YpVJEF8khx5yW5XH8geT7IPhfb1FG2kBGD
t2Q0aDUWY7hCrlnFayahCUi3qYHY7kcIGm1WqO4OdB7TDoJ5bBWwNm8JY8vTH9lo
kgG4SV8tyle4Z096rlISQcHLMf76mhQRSg2f9gTUSn+nHnC5rBEsvFY5i1+IB5FK
GlRYTo8M7L+MveTRHfIMTQW5FwdZzsapQCcJ4wQENLJjz+LABLJu79W6rJFw4t1o
alMqfcAzTH9Q9yyurBG2W9fRIypiO7ziZc1O82sghk3r/26UslxrJhECJtt9D3+o
3AHseQwY3VX7ETINq7x3b564u/zkpgokCpCjfPWusPdv3qUPTy3Pqt05j2B43Krb
amtgLQGifWu9z/8cUH4A8lc8IR5xlqS802//51rib8MJiUOd28OemCsj+ww0IZOh
UgBIau7lsEjkJK5icjXbbPtGAb8kDR86g402JazSIW+go06R7QXO0ByS5JtKka6M
RipHOnUEGmpsChnCBfMbCIk9s/Mid9aWioOCTX6ymgeZHYmJaaX0o+svcIhtK05+
vzZk9chNc1U5zYCIHoaogL7nROmfNPYFb5mOxOOC/MLE7DnR5XsIUg2MrQuwPzbh
TE8f3JVnY26OjQmdcsW/QbMNhWKSVKomsylfi0BCNvMWG5Jjz4X7OeCq44GVBASK
4cqDJcq9jjVDFCwUNCPPGsWJ5TwWgZw5zJFcSNlHaHik3kw6PixQuyjHjpoFzsVe
Dp3H0dtjWFTEbfnmgNJxIwkK6YrRTb/HqzDPTKyBiCAi6RdX1pBJTIEXDKkr+bfG
Zh3ZWU8WIA/AEKTfmyGb/FGZ8hBOcDyN4Mf0yQpBy3NeTLTiNk9t3wiqrPKcpckT
/SdRHOeWoyGGrtUfpsasUyfo1p6Rjpmte6ihKBCMqlnaBk/WCbJ0O0AGmwSUY4NB
sYAX6SeGqWwmlEbq65jAXETWwj11w7DcwyNxSxG2ap0VNDrW0t2R7VOyS0EX1KFw
Ioq8S3lJNTtTEfdTnZwYZNgKHtLVlIb7lOm9oQv6oJb3VQlTlHHazFqXRcc5dBYU
oMQSepa9g1sjSYkLhf05LdiBfZij7BqgVnhe8M+1j7K6bR2fbspX6vvSbN/buMDc
dVEUX/6Qe6CER5GHsHqHOYFI+/PNIDZi/zVHtJBcMNWukWKQ7Rntgp8j2sXxdDpI
4tjADgGf82mOAl1jy4L1DoXdNF2w9jyDJvjI3454DHa3lb+Y4RVvw5kuNlJXM9PI
A9SU/rOhvOUmR8hEjJJNGyZDYyRgKEO2X3W6l8b78Gkdlm9GJs0M3MBDYx30aTC/
LdjheporNohqcm1w6gRY9Gt5dnFdwvgi6rFLx+18hphhirBdEVolbhLI74k2OcPh
Lcd3v99bnikgKcg+KOetJV9Z8F+HP/02UpjxSkvwmec0RK/X4Ckifd52bBcRO0I5
DtYMiRa9mpH7bwg9EJdkgVt8Qtik4NqcotXvpiwLU9uu1/jp8vWl28VJW519I2HH
irpCTH75lZ0vKPDJWDtHQL9JtwO+XWLm55sblktuCzTJxkfa7VkB4DrT2WbuPtPi
C5UL8O204SdaKCK6iH/JSYU3Z4FYmhZn5VuNc1z3eyNC+fWORULWoyR59OK8Ra9P
k0re1g5T26JcnuQsOeNjO7gtGc8Fyq3iGq0PzdQPfPXLYHwsux5bp8lgavBsF/TM
0BpjuGyukhiFXvd10uMBV+U4r+Yx953S5ZAMZ1oqvvDNYDIQLZRw+Kl8pNThRyv5
h25JVdt3epLmkSHPBkB7BJXP1Sd2wVMzh6/+y2MmYDG7QRoPCXl/RcbLPbJLPoxF
B+GFA0lnE/g77cbZ339ADRAGV/0uwatbyuNvbxRDKYq3LRzqpfkQctGE9k+07ogn
VihXxM3Cmwp1Hc0Km4QmWq9dSZvirL38LZWQfuB0CNcuIa196hB3V1r7oL9sxxeZ
uZw/HQ668w2FEbPthaSO8Vi6DsenHsqeDq9Umyu5eoYQzS00ro5W3Obm4N39/1p7
g0r1EA1ONCcWZwCePQIci6Lzz+tw175s8w68032iMBC1xCd8xH1AqT969VemO3Do
oc5TQvHiV/m9+nGofBDd6I4HbkR9lcODoxVdWHhTrfVtu9wtRjq4gDDR6toChNTu
gNhC0ErGXSC3tsXAuNloeclEF/kbHhhh/XxqEUPwEHDrfzMmKqHbFoLHP/GUqKU+
4T+YWo7e3R2v9vIbXuYh/FSEGBfhCpKueO4wTBo4+/36hAmfCiu8sU+rdRI4U/oU
b5vhqi+x/bf8ChAJFA5CXngNJBVFlymuD0pMtlHCTeTtEVoYzmbmVQBu/iqdHZZ7
6yuWUfsaBlSJru7aoInrOQ4rnuGPtIR94CNKhxf1ER5JN+kaCZg578OCzA+BJh7Q
d2tNzuRDVnPXgmbuf3hHdkEk3djiak8tcAxbnF/m++GtBMdHWGeTcNKdojpaxJJJ
EUVbDIbmlW9CeKYhoPreTzzM5yDbEqS6gPFlwASlPxTpPhvXsqxxnOh7I3CiVg8s
6RINhi5sdgT7WXqk74lbiEslpROqH2ylbOU5k49RYxjm1fyqtChiRaqKTbV9S/x/
TyMoJaiR9VAxUMY7UgzkdqSMQ4AOGeym0L8oOoivh5ORgN7Mt3bDJIGkA2wjHnag
Y67tDlkTKbndDmCFVDNoOOwmLgYOjf79PGbMn4hXPoWqor7QbDbdWjaALs52xGIs
5837MU0fyWc9BOSrZBKL/bl+HxmKfR+IMsnT6ekBe+eKMyT+CUyL03iOpRe46JIm
axcMbO9pnhDn42NzUEMyetMf+HwZoVsjmBUadgFMMv1z2lt+pWZxTcBm9E+h+Ed3
vqPPfJOm2LEZIYkNpGJJa7FJtK0T7omanH16VH1EdhbO+nZZRDpv17MODYHbzAMt
rpr/DUzY7cpqBvy9akajf0osbDA+jPKYKqwz7jjjR1N39jgZmB35UeCQRwjW/Lvt
d8o4Od1LZXmgpAaMIA83QdvVfrY/7BrId78Ulf1wkrZRt4LGBkjh+walmbz/NUUB
k0VcRAidGOonTnhjpESuUfvT3sJMxhuiP6Mvc4Ci3ORz9eJVTIx5umwMyr9c7PAV
0TzeRsfI28Rk2d394JYoiwO63CKwEQCOVYLzXj6cxD95X2VumhT+Si1tL1s6+FS9
yNngvEAJ1JvIi4wg98362HAaRCF1EGNvIo6Isg4ZCkKgXI2+KWD/KpjKsQioGveK
GRu015Nzcf4EuLxLMoUN6yCBRJzTXi1wx4Yc4gYRDKxecxMJkDTf7SqopsZSl9YU
Ld6rdm/uCHsV2oH9XGVU/GCSTE9cTzH1MzmTe/ObHD2vLi26+7pzRcvV/sMxRQyJ
iLJZ+C3l8yTYBjRS6HRWdkDJDTOz3HMM2yP/PF4RU7Sa7Cq6/BOX/E2eq4UvLfJf
SDdpTPVjZz6dS7vV8JkZLUdT4XOqqZsAiu4bFIIxJEtz9SDokJFwSB66BUblF7pd
M25Gl+lYblaAUpGOl8F7gtBGLKHjrUOeKUP0Dog9zczSgKmsLDKNYNfsKkmGSVXO
NBV8kA61ExjpdtFib9e5OPCytFTu/OQHYFO9P+gRt1mO7BT1WJ9fVrX1bfsKIiHN
L+0CqSl61Tj0IxLpbLl4CKjjZhAcBlJSnWZy7RHrSoZmxKM/tM3nyHEdtmIFQiiV
TenrmAFV0zl+S/n0v2ntnWS1qE5vkBTrBl7dN1rFEuQic0wxU4tVb5oKEYUoVLbF
3Q+3kWYsOiSdbIQh42cFDxrtNySNVVtHI7jyuvJgs3+PhQGHqTQzqxF8XC4fb8S9
UYiiX1TUx9vCdESrvzets4/1UUYfTEJ7Y8AvXvpP2/FOIyV0wQscISohoKygsmiQ
pJn6WgunP2n4HWBEEWNMbEJ6VikYybPPFN2XdwZzGXQ3+oDZLpdSJmuAYXzdZsTR
wtF2eXCXfSNp1Wo38SkvheRX7WF7QOjV6RbaPMw7Y9fAOudnx+rVW6/HfYCTShDu
VaQutSO5A7+aAzCF5qX3z8t+8amKTJ9g0zKLk+pfjf5vpaE52PvLAq5E2MUU79X6
SWiC/KjAYqz3vbr5L1OhE9FaWI6gvg6fZS7TEDP7xJ3omLl9nDYimcHgLeNuHDyn
wabL9jvsWgWVJ6dBHCVCzj7IfZQQ+/RxW0FsiR9APbYD8Ywy8h082vcqAs5s2NS5
dHOirtkmohpEewNhwUVjQXw6II1DcRkX4KOiON73DDyn/tHQc45uxD29c0NVHm6G
KVbPHHS18g3fSad/gPnobNFB/JrUtWaaVYYKhDz95fTQaStVxhne2IzMnUFEkJHr
q3AsuEsrTRi2DZStnX/wD1I6kk0YNtu/6HOUOShDtBCFoCJ5gkJpUNUDRQreBiLS
xNRWaaGNwLIdNSPYSYvYHQtouLfXzHtw2R/GtNs/Tzzcy20QUeQw9wimAP9YKjnJ
T0QLUXuuXeLtNCq5qW9ICErRQgg2bp/EUVoee6REQN3BiRY2MfoteYKKvICSFnhX
8ZGhXzUhzQGukVhyRkkXfG/jDkK2FgrTRDBtVgsZ/CHtOvweo0bIy5st68iZeNjY
qlUrwDTPJIeI089OosdafloXHqUDmH9SviFxYziuuXv1BHS+5Qq/fBBcOLSMyS+R
yG4Qev3iktRJj/Oea7Uk95jTVDvBYBwpf1ORnhmh5aOTP2Ahqd/f1hWdO6qnf/Jy
l37tjUvpJtvzdCsBlFzoIKbydSXg1VZ/LkpXJ0LyBug6hSxO6Dv5h+ybKyp7EQ7L
mP5CQXpeuf8i3ptbDyztqHYIkzLjHkY7cKqtIzGhc2iv2JPx6hWO93IkSFApFTKl
7c749G1w6YQFYZGrKi44WhA3rBe9yqZ95uvOe2DOYTmHHsDjrUbGDzW6GN2/VfRh
BDuEzQEKMAtPO3VIl8LV7P72UwgCuthx0nu+a1XUwcyh6hgH9nfG7RY5K3FAw09v
fz0SuDFv/wkFHvIJ4cB0Jeh5+5by91AAx9bO22ogIqEviOg43M3lDLkXw9Dgroll
sDFbUuzGFsPdKO6ksavSE63RbwaJDA/4Gm3MWsyTB5G40NgndzmGeY3aDbuIMsnH
fCEAWCM7+psg8Kp4a1dqoBlWtcQdkQcjVkqlz7BQOlpGEfbUnB/j4cLES2+e9TKQ
cGf8lwViD0p/kPNQsZzU/4mmqDNzhqlfhbWAdcj3WonxlFwu/Oj7LMmsS213yUfQ
XnPnf3FsYM36AyDaCbtJokgVe0P5QLQVT1yZeq+gLGU4SHkXS5/FWyF5yE/9oGce
Cl0mfhiXux1dYBmdmy9UvsD+ew9Z+QcdaX4ejv98jFFy2Nie7YH8/qeQwXyekjdJ
quin0YWq+uBH9fp0K4riH8ydTs8Z7dDLTXwOQBX0oSlSxzTnJLG9eDZVTg0vMH3f
uVIhl3aY45o6BmnVuYghu0ikLpeiFusBVGfEWLrSGFrUDU9sDP2HVNbwgY2XDfMK
nXJvbVAADd5gIt1rToQMbKKp7y2aKVCJ+dvLnigtZpqwhp46vgot0rDPAa07Df7R
rSgm0zOa5mhIVy7LYnkk7KWPLGqcTZJwEamqel500B4PZ1y5jyqNeI9HGDyAgibq
H8yiA/wZBgSTVuwYQMQu+tNY+l+QRULaj33hLDLTn6tGh0l8v6O1eIPmI8Bu9zpi
1Fb/k8EEB9pyQHu4LmnzkkUgDzOFuN33f3gIk6qws7y3hUOOWRQ4i2KSoMCg5UPV
nUBNmi8eLWG/Tw5+M/BxOuXo5jqGA7wtKYTBFWdHI/EaHJYl1dbDxvjKPu8Zv86x
stxXBZYloXbFKm4V11yFoeVvgQVO6sYXTG2+gwkoN8b275BxZSjlNHfD3yxcHxOx
B6BXmGO81apQ2iJNatKi0hgNzg5e0pKaWmvuK1hrCJL1jaFgBQYj7peGgLkLWspn
3CnevT192DDW1gEc6dgaDbR8VDKg0W50YEY1M8WXQSeg6ZVRb/1YVGmh0f8E5bUx
3Tql8i3dRVvL7iTp/zfh4H3lAI1cxjZW+yU5cYrtW6XbVrSzhe441M2k09pdavQB
kteS0ssfJzzFN0KwO9PkEGpgkF6eZ/J69OcMbNxjCN1x8U0XW9ymlatozg40Cog+
1zHTyQS+Rrh2PY9e1EZxI17Zb+2yNNnyZ+DDl/1OfEpvIf1hOiXhCS254UmLSeVc
YeWsQMI3hlJdbcUvs/ZpeF8MxquVmgUXPrGYzjuLGIPcQ8D3cQPWaR5LoT0krYvV
d2ztkIELPAxoImw43YHfaYf3Hwf/aryzwiv19EjlROj2bU9Q3GZeC/yhu/NMgyWw
zcoSRaybWdffk5BaSxxzncsRp6EfbKQqwqBRchwNNsw9oBq/D/fAa2rUqSUucf/j
eGzaXKNL9mCQoNfRR2blkXLfJIoH4FuFUh+M1Mh5grQY5Uqa9yPpWuRDkIeYT8EH
OZ3K9M5CvvO051jsR82MzYUqeYwZE5pRZ58GpFYrhvMfO8ynwvlRn9K+UDAxlYVO
nELV5eTBvzumrVlr391YLzRiIBV0mPn8MqpW1dfKOOnI/4n/aTqDfI8k+iyd01pW
s6X0ycZfRYeySrpGTfhxwCAhW3SmJtyZoeGPoKH4w+D4vLgSPsoHX7UrsmI/NFiH
X1nNaxYvC3taVgEdKWiipMRAqK0sHaXJvySLJEZbkvLKYVzVpbIsyxVYU75Vfjgy
aaGlYARlnnNmcWATy+ZIRsWjCdPSCqBvV36/aXUNch+pukrAZRiNorlw+zrxPHx2
o+Klk2HXcmi019Lj2pMTfYfJrR7yeTi+YPw09gLRWUaUT9hLBs8QR9B15guD4Elf
lFUvHOIgMpAl2kfcHP7/LEfTtAtMM7oyDzdMolyMniGxGJ2GTiYs0WP1sTR/a5db
v9T0BTuSbaS71g1gGrivbFZ1WdVltVgXImeTkoDORFO/DzB4b7mbf8yVo9RaqEO7
qB7/cxN+eOanwrMvH9ERt5fF7J0TNqvJceS3ac5gwuf1Iu1dteWQlQLvYTdMdrTv
5ImV4ohu1N42SzFJdhzUNrtykIrOBnL7WoqZzIsO6N1WpkcDngjcaA38/5EXSmlz
Xj0Mh9bcgca8sIQfEVERQ2IyoV5MPlFg7jKDn7gZmy2oCWYi+5gd/Mh2vcwNen/Y
eU+SaRGpX7XwfViqIWflSea9rnoTKKN0CZjkq2auN3UaOjT4bj4p1z+Gh73NZG+X
DBUqwDfiFIszRbB2gkeSEpDoDGKdBiZnesup7g/eiGTRmlfSBUfPnhu2sHuU0kSn
a9WkfH/kiEaQ9cXZuZmODTttty9dtEfCScLY7dPfgKuI0ijhl1y/Dr4rApMyfSNu
yAsjciOxDdan5OnAxh5MJqV5Qx3kTprN3QL5R3g1YYt9DauOdNjnpRPBy2so877p
L25haJue1XRz5dLwTaaHEU5m9ThI2NyHaLfXUyHOm1TKfmlqOlOuQSE03OdOAqxM
klvlYtz7yXg7h5s2H3c2rAz2eDlw5rLv+D5Slrw5FkYREa7zGYmeG6nK7b1JJSJi
Q4KsPaWnIxRqfzt6aFzT3ruEVMqx7wnB+Q1sLMGJEygnoYGao+bAG9+wWfcf97Jc
+b8BL6CZjSYeWawG/RmKQ5ltzGVEqY3H2Z218ypdmb2Jxx0G6xRivW0jESC3KfNb
j0ag2z61+NiBlxEQ8Piyw/AKquHR1nqiI4x/fWVaz8ZSHiEJ9V7PHmoDl/c7sQtt
s9TZscFCbJuP3W+Y4+XAUOvDKl7G95C7x9WiZfkhABmpMYAd3rydj5IZLvygytaw
SWSCp0iWJNPokj64HHfs01UAQT75IAOqnEDrlWt7tnFpaThCith36GmFZd9W1QZO
V5x0RnO2DH2UyYsnB9qpabixmRc9+yoWaSFWxBlnBuHpRQjPGohidT3k4YdQ7waG
87umG2HzoCms591fEZGmXaQO7+OSfrJcrf1Ftq2o77pCWXdVD4BfMW4vy2jqLTBF
Fov7CMweqDa7V+Q9Ynp5cIJ1r7vOnUpP11RcATN3nZzSyxN19GB7vuupMhxxShKd
f3bGn+Q2fIuw+NtcwHDC+ijNp5aGEjQP5+RYC3MmZhmr1q2glhMi0h1+Prr9jtfu
PYDX8TjG7AwFXYyG8YrIIzJfnPogm6tcuOI7xehtsVvZy1171vv5j+ffaWsgQmjv
K4JEjDAo3cbzhWRUnaRhGYR+aemtgWAtZCjOWTs5Awp9mCtbFo+hg4LperHl9WZ/
KVzfd+vCRkiyvNDhPPXeKxZX9dZeSYXWYC+N8nIVxnA40T4au8OlhC8BYrBIkkcA
CcQXeEn2Q/6PNBSJk7fK/Yq0IAv/rpt+4HW8Ey7IDoBQKD4o/PRn1CfJpVS2lbiZ
yIS9/I27WsjUlK27it1n4HP4hmdOaD3knRyu5hAaAtuG+foVYgpymcZIgcIQ9UPz
S6poREeaNlBpeYoyhmW26ME35h5rdU2vjm2Ltcd+Cditwpd4bzeRhFIoCF6DMHrp
MlwcEKvowNRn/d5OVjRIZLdajVZuYbZCm1ddoADLNA2palvtIqT1HrT6Mnl5QLdw
6g5LvY7yfzDN3+euO6E9Scy24O2B2jcT61E7RtqSwskzr2rYtpAMQfkje+oYb1GL
16M72leYNQTVQa03BWPseePmszdHwsHEHg94PHimh/e4naDcBs8YSAivgldS1Bm7
hfeCtihCrIxiNQvJYKr3Ob06MvsnIjdzap/zkWtSBEIpbVALosyWC6jPEoWG7JQM
5wO8nJ1bNZqd6PTARNQPJ+mI1JVTTlBLganIoC4gvPSAW2HH/BZ3En1IY+6w3O1N
hpXq64igoHuL46OGnRj4GG1cWUmISiE6ILrZ5+mqHU663NN8OfbE3BRj8q2UwejZ
eh7OXWc3hJsAMPM9Gxpw0pspPVCwO9F6QjiE1/KsF1jw/mY6g6lbJd08ffC4OnXZ
+6apRsTrth9OKFDAbCdevX7C2UQDQhVUxkIGJZ4kZmKgLym1rjSDfvlyJ4LqLNa7
J0NMsuoizdUkyuvvwvBMY2pf/Jso7szfw+tq9dWg/0B9O1sdozPNv/Zud9bDs2cF
IfMWnTCyjdDQmq8FbK1mMR3G/z+fbLaBY9DPJlkdLTpskr7R2wjJas6jpLYWRvg1
O1Un242ybHRUnFEoaUMUenn2vsaQXJMZuV1FhJHXNGbt0aN4niyHDG9IgqJI1ads
U496YEdz6vracYrRByuQlcQyZkQ9f9TnLH59bOPI7EZbYZqU/c6z+3JRfI7FrmZa
utPIGR/8wHXfx188W1onF43CxU1BdkY+wt1DVvG5l3zLVbHjPoi/oJJbeOY+OGuO
9hU8EOkGJbVys8RxrdiM2+8G7sBU28uLIlCgLwbm/WFTxzWVJxkQ1n+JgyJycSki
w17KwX1PkciSmfCxJxick1eoG5dKfsePqjh36NmgIV/x/uaNjgwEi6/eEJwitUkN
No3CbJTe5wlTYbDB42gfljGu5NtYfMr7sJq5yGoLlKh82gueD61i5XpLX1/uSU3q
TNP6QCbJTpeN9SB790s6PA3jH0oNFV1tZlJ74lvhx3uSNU91fZd4hOCKajaS8zus
seVOqJc8jyw3JHG+q0IN5fZAQ4ANEjs0bIYSbrhtyErtPisrloC0/o+phe5R1wWY
GROtwgpnKPm/G8gyLOLxnHqDhAgtbV2yhB3/V2NeAhFlawUSX1P2sOjJQoYMsZvN
3UdyJPNZl4/ehC4dC9X0NHMQXzimgP4+ALVZGBfWhLM/61UyKQN45s0kkpQFAJZI
+x6reob+N/PBwomFLFyn0aSr+L68rtDkc8FlFMo5PwJ50OneOPBmnj8hO7eqd7iS
s5FeK4bwWBW+tuUi4V4K0KaNjSsFQ3iRGyl6I8UwZYWVQuQIuhQl5pPmS6y7Nojs
GysttACv6oFqe5ZzkcEH6KwqvQ4xY4vULF2LwEgLZrL7XF4SkEgpfiUIfeg73dvZ
GCDlbHP612U0t6v05LdCwCMkyckrPHSDyWAZ5hIgiDaWDk6Vg6ux2FrYLXAiW2gD
AebcS+Xk1dzbg0iRApYgYCxKmcpgrmZAWwg9+mLQDTZr9g/mU+2DcZn5hbO795L5
tEXHrQkimzJ4jv7uKBWyG46FPAw9hAZEhNUu5WuUzBiDDtpcCX04OBvCJCW4Q2FM
L1YxA+mMXIxbVPYU7ZQT3pPP7NdxNhIYWoornk42yh6wBRizjz/ppLPUYOptVRsk
fR8oUrpycWGC+oNB5IEUpGj4FHYurqBG+DlzOlzzusY4fpzJSBmeVJdLiSN5pOTW
rtuG9Rf/vomNyasqDBzt5qkQfLBNGZd3Hyijo7PePQ9/84aPYHpNsksKtKetTr1z
kemcpc7dD67gcBEAW5+DaJ4bQRmuMcrYrTi8yhkZ+zXrje8aGzRUXIkyoGoN3OJC
+WObJUD7js+1zlpRQ34/4r2u62V7MNOI/u6Bovk2B9oIHE0p37vWOX/Rm8vJEE4h
BWQE9vRDtSnyrRIHq473RYZMOYIfbRaRzgx7/GF3M5bxcFS3tQ0LV0qVwWzcvGlG
BFNL6xHg0bjo5ov/FKYGFVOBPtaLe69NnQcJdW5atK9knTIK68KRY0kbOTAC8Sb/
QzWMB81dy6NqA5DxmxsGk0cUudi+N4csRBG/0CKKjvFqrwubvEJUnnHKDzuiF/d6
dFB+eGR5GM0Qzi/KVpRPPE/m9P+2qdAqQZAOY3Kp1bBneJDEWyNY1q4COZ4OuX6l
ybY6hlvsbD9B6n8fNu06bV3psgj9PXzR4oGL7wcTBTMig4ImWqpl9iDQzWm6S0IT
FknA9+e9JubbxtY39TAj75m8k9/hxVYUlRjvM63vLcqTD8XK5mwvt9ko4JGZ9hGL
Sh6PNKBxDPfl57r+oNSb9Uj1R3OyMupRhwOWqKhN/AketbYwFekrlpH6eujr0z7Y
3OfTZZuq8cruAuya2600ANoV8WiUFm3fztOd5YlePy8a882u+gXTgRulDvnch6UE
q18eW36fMS2dmDJna1embjcJNciqxBdkuFYckqS0mgljF3Bd094hwTHGbbIiwvam
DtvP0MCujwemDcikJCBU7m2QQQTc+LGhR0IKEj8GEI5c2T5bwR91J4/WlNreAD+3
lwQs77QIi8D+k9PyGUxznlsjfvOa8DdIXWMPgvG8imQ5N+PohTTxN0cH6qBpoysj
v1DsTKU4o0rdkUgdzTlvnxgQCElIBtU56b51QQYXv7xq+TWN48/jS29ne+NjIAkB
tKpxHu4lNLDvVBAr/CU/aIbT2P06/KpbaeHLtzxScPFSccg5RPYpdFt5aSM1t1O3
XNBmZEDMN7ijklwkcsEC8lrOEUT9p37UmvrESZwk4rru7wUUrXMXKXvys5bCTByD
exLeSOA6bAoIfIW7EZxnai0lOWYsWkUAT7M+2saGwh0JpSXWCfEw4uJmdsTjhhsD
yI+OkQ3aGGuYjL0RmKv1eAYJ5JAbaFMEPCNcfyOYLI+nVFuxmc4ImHLjDNSsP8ll
m0KZKyQgSXhb2oqU/cYkFJBs67URPtVnTlawMhbSjGtDGzVQci6CrVkyMk/37FwU
Gu/YM7xnrPFm+QxLzqosxMRW/FWeTIzgMvf9QAo6L64rk3UrHTyAWibopIWxewIH
IAl/5REPM1v6mslzYuuDcx60QE6NNfcvtqsMeFyxG4Aha+Kz3PxUFSqSTpSYxIM4
Ns+DRYB3Vring7Tv01/KnNfKWXk+P5dnzqEPPv3okl1bAXOCAnsO38D07yXaOzle
fP8TmZLHkcj0/Se3MmTWsXSWCuY9OSysmfIFec7EJmz9omA+6/MgubuJnCR1X1dJ
Pzw+DzU35TS388ELbEysdgeLITxtQimmlp0IU2czN0Y6l7SsQr+UEHtBro3lraeT
XTNF+TojQPP3sYxXj8d4KL47rOS6uIJVsxEjzhNJC6q2Q5EBvDZc4EaS8ccAn+2e
1OozoyoI1ZcGKLQUlOrd7wIFuf2up4f4SXhxBjTrCWByo28+d+bUnOymSfh+45Z1
adTXZWG+opIbSauE1h7vtndu2Zoy6dQx2ZmVkH4+BGC7TmbNE8fnWbhtddBXr9eZ
/yqL6WnRPtv8Y2GhROqn9UyLigqhrJfp9Ga0o66s46SWwVwZqlXDSIMgnlm/+dux
3jIs1KiAp+o3DatKlPbKrRhlRM7LIu8TaWRTCh1FDGseCkEWgjqf8jsbmDTDhMNT
0h9U7QpNxp0x65GMMP/IWnCl49JFyozqZP/62kGMRxETdqjqWiVl2e/xEUirE+CV
t3HvOHGflhwfV9whe+1hyl04w5I6d3hI8VLwVs8+yyUmHOzOpLoh5uEuNz/iSmR0
Qy+DLFSoWizg9kZba3UqGVRhINXQUDexIz7w6vhUyU257MH+4isRYITc8eauE7lg
DG83YbIm6RYA/U7RC7AUCv65WAt0CC1BRlXK03ytCdnvA4sZ0GiWZMVUXPpIp3V3
K+/4S2tbDWoyJ1MpNJ69+q/XtGJ91QjrOLvjkq714juFsdM2TK/50APNTMlw6QFh
u0AtMNqc1JpIOLypDPsQdLLDRgml1804atQmeADM1z4fQMuRU9G/aoCuHeuJ3SsN
C5O3K2J98LIQsF8Z2Hh4+nziLH/Tmp0D9OkizuJseYRmdtf3yh00694K+TcsWqXQ
tB5+cbuaKLxVqscriwVKz6kTmWI5F0JYpNOQbMOo9HtNoovjUFDSEFTlwZlU9xCZ
hyiSKp/hhYlwM58DXp8/SLcBEuhJehuR9Zsh6AS4RVtzBnBM8VMuJLJEEjCjssEZ
umcRFJOAhdE3DyVXqox0CcFBpXoKljQsceanfs7P8nLpT/Pi3mxWhvTtcCpllxCF
PNEzPKErViF1S8LVXzp4Rk01U2kkR4DCISVxwf3wsC8zwCpyhwV0KTJpMhKsKEDF
cqMzmEUounjqwCOLanpPRQlf8SBn+aw+OzjE5KR7OcE/OzKWtrrfoUjABwmZHUW4
9+70shhbP/hF2EEMJG/VXzwPzQ1izTL6x1rBpWHsnWA40XsEecETlg8yL3hGFjVF
0lQS5O2xMDV3O9N8ZStzwYpAROWXRJg5svXmdRASGXWzO1olHDq1bbpVfNM9RAVf
WxCbiDyE4KLuMK+lAHEoWXgo4canILaC6ERbMQX+lzsmBHk6h29fZy4zUqQBTNuo
tlLAOT6sISke1Yx5YQadQXy9kJffROjQDwKvfB9nSHVUDH1LQaJalr9b+OEo0MPF
fW0Tz+UhwOrT7FzNGPWJYUDUT0otS8l9vM4a86UdJRKj8Me+sj6A0sLQeF+xJyYL
zSPs8K3nsbVd7r+LcUbPjVKnj64SVe6OVihi7LmkPLPTFnthOeFVwmD+DBA61JNs
ujQWJuxtwLf6DM2n3S3Vc+AhDZnhy2NebDiQn7qllYN1l86do/6O80eHPdVLKVh6
rtGjEeWe/12zAW6yIi2cgWEUr/ZeB18CwXopNVjRTxoNcVVgPiy6Wyd2DqkvkAns
kVrNS8BRbIQwcKhmCHz08mplBsQQtkd8fhKOBCsmeospZDFHyJucvSK/bLIhiSOS
Kb+ARYFCI8PJHMPI7GL+p12xo8OrbZgY4N3L6P6l3JUY7lEVrURL7Njnzhk9aJxA
iTzgU5EcvRLkRdjfbUnfuYq7p1KPWqRVnjvRigJ0Z4InDgA9iOvlsQi2XIktVG6F
kap4UpAbJ2QC3t+yUu1nEon2lWvlJTEvIMrjx6pu5LHK11+gttXv+8L3mQoPlUnz
LfORv7b/J9a3EC/d/mTiClb/J2DJqbYu560GuusiLDoggqdOKO3lJpL4lQqHALER
2ILB9E5jNTIeajo960Gtw7Fl7FNbmMDA6qAak3jsCPvSzSJL2pzyRw7HggBCP5uf
16COTHNg7UkCCMYQFcbr4/nZe8vTiEkMvHvYcSUasGgHpS7EXbzgVonZd8Q4LJHb
EhxIbWKO+etUK4Oj4ZF1SfhqcHDfsKK4X3uafeyVkVRJ/YetLQnAatzDQubPhwq3
47VvIFk6U91Umu0M2mutEfR5lx6fh/RNz3GtadSfEKRdN02z9sN8EUa6IFXAbJaF
Pga+E81vGt2o96fuKQAnIEfUaWXvKLrzoISy6gf8yA5vcIurPfqaMNqluSyyVUT5
RP9nJLO2RQ7G1A/begVRtd27uO9XoAnv91mm5tX+YRd/8lfh4ufg5qr6gfamEXCT
uGCZQpTWYwj+MlluCI4XAQMF2GfpCCBoDD/6SMDK2bUZ5eu/WPAKqKOkdSLj3xF4
9M3BrYMcIa7ZyRr8/gj55biRmMtOF5gCIJJ94PQNooe/Pg4tmXb0FJnH5qLWHwpi
DTEjidEp0fs5ECdDIZH/A0LmjS12FOlHLYDtnJJgyuip0RG+2+AVQvSkyKfExRo/
ik4KKRYlYWOXw0/NmMQSuSP1nTHLkuj1Nhp3niz2PSfGuBH46KOvrShXYbHE0nit
S4ylVcBbDD9iC5uxqn/n4j+D+pu1aZbR5kxc+ROVdZdFixCY9RYgWDEi/de9LBMR
IWYMg8IyFOCu+7k93JXdSlu+teRzwFB2FMb79V+xxfeomGIW5WG2XkjGEhaOThpf
/lIUdW1rrS/9c8aqwqG8H96YhCLl8P8QD5PgGeBed6r+4uFFlNxeuaBQGrrZnLUU
A3cnFr0WH0dNhnOXH7xHP7MaE95slUQei+tUWnUOaw47HJV9jizB0ozE7stxsycq
CTKBC9sZAtL7EgeF0JNeLMHATdr7PkFJ7tAy7YSc+PZIsiof8zmHWf1+MZvsT98l
y/IHLOAXI7OnNVA84zBsxwvLwZbZodKCfjJOpGdJ41hakkRGJl0bRevOv4Da/55Z
n9XDMkg4wvs8zFNnBSfsz2/8f5hE3KOWrVH9zq5OMWHuoMwY7hxy8bV+XyEVTwdU
YpNvktPTQkRr5A7VzNtpXmfZ1Ac2dvdCT1/2u3FUTxzwVJdBjSwWS0Z2Nuddfl80
JfbnLeM6RBK8TR4lnlAHkwjQy2Au6J1FWaqZ0TpT+P/KBsrc6FVG9eNoYUu5GecL
cMPgEhB3vsusiAqsc8Srdb208LZpXZbQnr/5KK4r9SZ5h2duB416W4d/pRENLH44
atEIcTUGT2IeeyP+AnzV3o/L/ENAObDWXscnXaG5BS5ASE1RKiMGhfUXXprQrqPM
7yG3VzBZtMfpJ4OvaauD3P+OFBe7duP2WP5H8r9sid7XuE/lN1E+XgPuwWBpnO1o
zNSEJu9aLJBTxm+7KZRXU7eASNLza0Bu75fzluPfnFYJL+u8nFybDvs8pGB/S/CA
65Er/qVquhusay0zFW2EF6RRRv9e6HM/52b2P8kDbjNIbcysh4RzFqWVRz23bLQe
ZM+x78DNVNWxok/GjXPq27WP6ROycLsuMYVoN3PE3+AT69FqAArhnzrj0TLuQg5B
/1u2r9IEoFjq5OXr8anj8WI5mjwy6uGhOANa6XBAe9WyRc0O7iNasii2XHDaa2FZ
luX1Lu3L1qT7pCXklQekF4prE4YiI0yxr7UM6xLT9XL3n5nejUI5y3evZThtDT6u
ejvamXjZ5lXpEm9hTMUa5iTMBlrhFEHxTl3SG2IxelTAPa6V/MRsr0IvCufAj3p7
v5ha6UKwZRFAge83J0YN9Pw067CUcdq3BqIYNwfKgggWHXgVg5SW+K7Lj4fbaa24
NpngQniT1B34vGlzXK7bqKbJVVtm1Vn1gKoDEdPb8SQYXWBsRdfBc+hrhpOZhhZo
U69OzwoShAnWIp5EAJosPGLHjHEwPGj/Y/QP2LieYu4BeY8LbI8FST7z5FD36tzn
VkUP4Y2JDZj9jsoLpu2GlZ/5QhfFh6cLYhWZlH3XazGcyh3iMuOXN8w03Mk1DYFv
UezaszgVy/qxX0ohYcs3A3ZwmIpAk6G7OvQyS1s4NNILnM++nhJVL+5LHpLpk/81
vJK5ruuIuuU68qUzhBv+HEzQgQM0QSUeakOx9UloQRIwDtAE3lEkJjVTPJjTJYob
TyhpSKrqqlW4e0jHEBru/WzFLSWeiIlZSLIgk4kZVI0ReUNZ50OZTxMNBjHq8Qwi
9+YmekeAHfUiBCSLrDgOf0oR+NylYb95/z00tf7gLsg9Mpon/L2AeenEMgXpoBGd
EoZag2/NV5334bioS+4LiD674xGiqeVDcvY0yysb6d4htF0j+zSuoMOnGzQCrKLq
cFDXvPX1gN4SWWJU28Al0ScLeSXhelFapLryM7ADUw28R7ClP6NMWyVV5Ra3LEzE
MUmn/XMc6pFfMXSaxtYKiG/A3urye7pbtGMm1lcQOPoer9V+ikwCLb756ygs1FJZ
j32GzO/uKJcOtTRUe0I2LjND7l49q550jMZaYtz7UObrEhBHUWkwy9HCmeG4OJOy
c9YUXg74VG+9A2ekGTKBtDvvEgvXN5uiEkcFd9iT8HJJ6aOSykvAbHv9fXqvTqZ1
y3PIr/1h4C0aFCNoPdA5LEr1N/AeqLn2GVYhqP2nhuM8r3izeIIuA8tMs7akiQTN
twkfkvXv+momSOFK8DeiVbOso3/gmd1M5w7PCNPlWWlSSfR6yGWUWRdfuunuLLBO
GyNnvTBqlyNklyKI3hZE6szuK5Jct76n/gV1wPq4/7gbUrD0iiEhVrghOc2pM/Ov
QFPqpYtjQ2NJy5tpgnzp51Cw4U8efATdzdq9fzyBKzc526s/VZKCltsdBGzssO6Q
aFNIAtEKgpEIl1PLYdczMrz7UTLYevaQ/zB15wwCbJ0T6kuhMCA4LkmUfxKgZlht
JvW1+f6L7kQTiyXEUhDrpCNfqN7tY0jHiSkooWjGw7khmJkBYoryank/F0q6Jw+Q
GRc59gIqCl/uLQbC9ERh+NM9BcmuxHJwEmkQUnm5+ZMkaLKh9sVuFvgZHh9BX0sT
lXlz9s0vAS7SUTVUqY1XgIRGkAJRUFeyMGQ/+M7MHceTtqhnQaPdVcidh9tGhDC6
7bDeAVckH1CPDK2jhWlbjh954cja65UNrpLs2SvXAqfVXrJzcxJtr2TwltuwwLmZ
NMYeuOlFC3tqd0TLiq1Pn/mDTgqa2CWEtNmfcSMb9xNB8VrfpSOMtrdUvnUWZriF
cQQ3ksgcExg3ZuHB/P6FXzUwYOjOGepq+atolKiePI2bZlsyRAHnNwDWNAt4YLHV
nc6lGc8CCqNfGvckik0d31GMKUk4cRqQvy1EzNo5n8j6F+PKB7Cbz6f4AvI85AMq
kDVV6YCX1q6ESoESpVtdQjf5PvpCDI7iY48b+B/1nI9ylTGKCcC0ehhzK/8dl7tQ
0K8aXUPDdMU77kLaZIs/Sq+E85lpYSMz8VJpB6/VTo8pesDLYKNjHCg1IQsAC4KT
yUi9xfsJoVO2oM4BZufiLOofig6t1UDd7zigEqPU1xU5V9QfCxHyp96xWoF9ZfDu
CHnOIKaN0l/oxaztBsC1tOiZQ8SskfHSkVVZJP575Pn8n25W4Z5CqafkzwkAKote
Ax+Spm0OdLVBxpQ1/pnaA6+Tmi1pHNhvQjRe/ZbqfYozTN6HxvYbfG4xyaFvS9gX
MqdxGAeYC84hC/t+qMdjV6mB70m9sTLcMOpLWYewWat4ZEByF1YA1nHlqCYJPU3v
xGch+YMnsso3p5iAfz/m7VTo7SiTOYllauFv0fobGyo5DHCQsJ4rK1tnF6HhcIdX
9jHQ4G06/YEkMiq456neZnLh+GyYaw/MQRMqu45u8CLfXohOe6groZkU5yak0jzB
uKzcwl6u02ZmZ5tjNAJl7zEWqdqbCp8FGwxSA0465gkFyVD9hKLDsUbADaRmuC4b
Dvm+PPyYed/kMmtXlK82brt5/dfTj/PjdLyJZL2vroypCU3BWptKRDG2tgFvD1TA
MVNCo0MVQmOp6lsKsnjoUs1df0bPF1cuFmCUNXRoh4Of8DoekdDsSbJ8g/LkxM7N
5QLkOLKeKnBPXjdDGw541Rf4Yv4Nk6h3tEbAZDxDFR8FJQgoNftPWeH0tVP2EPmy
cgrwG3kyIPKyRQYSZNMztP1fIUrJTuVpqJh+DDs3nv/50hX9+jNYvCnOMg3fOIa1
k/OMpXlmqohNkz84FerQk3X9Eo3XJ8bpXGF1P41JSBtm68YO53wb5KShkY4SX401
cWCWlX0SLM9hbpm35jcdqRCYR4ExYO/2I9/RUswF5fD1M/KQR7beBqulIBQGnLnf
NU7fyJdsoBHFQAoM4561H4Q06KGC9YGG/HEFjgYVibONvweqqHlqvQQR9qhdryGH
akR4xcUGsJCUNwu6SAbOqe5EzHLpEQptwX5BUzcE4zDPrG9Gc4owRTO2J7jCGJrt
JIYERJTyoWSinGPTU0KVzgzPZ8+yNZuFOdVCfsPblEmh2kLjQ7qTaUjVQbjat+Yr
YiAR0jz78/wbXiGNRO1pwXT0/9oqeSmVNrAxE5dKzEfoa3m/R3i1PBZALBDCC6GE
Kph02cF11fP+6fDYB/Lg5isg2EPqegTzdBcesP47yh+qPgw2pcp4mA+KFwaXm7bA
YkmE2TMHE7RzPS+m5IOLWHXSigYmQaFb77r9GJydIc/8NSJVlci+QRq+N8xgZzq2
cTYA+cvJDIdhYi/+m6F0rSv40NmZaU3GR2Q0sriMAqzuSRu7NFd4qpz14D8kdWNT
ecgX0z0kvCPUcEQOMX2D9h9Ne0y/UApjRt/lCVY9xY/t1iD3DeDkFpRh3ZobSc0r
5vKd63/buzGQ+C6RuVvvoHlHMEDaJJ4b5HENTfzlMwBF0KPhD1czwFhlOQKtisrK
/bZZqAngvYF7JKcck31G+1QovEZUQXvOv3xWNxylHdPlnCt4Vb4jvbyQlOkhezdu
U74gSwFpZsqs4OoyXQQ7BnRW4++iiQuxOM4V24aHJGhfx7gn3ZibaKXzfsuOrKer
nGlujz4sdsUzw7dslc4naxxRhxfytwIg9GTcCwszv4QUOSSPIL2U0uV/Lkvv/Ddk
thYFM7Nc6JSUai/pLOhVBL6CvmuSgmKFBmJa7kI542ibcMeQO7Y3YZPZ0gB8SpXT
OL5Q8KVf6CPM/Z7kJNhoP7ER/GpsoU5CW6dQv94ccu2xJEUOl/ak2w1JY0WXFKoy
hp8WlOSkoiE3LK4jOBgSGukkc1SagbYDDzbn8/toagZjqgSmj6OLwr43N2Ph/wuC
mIp8WLwqUikjbXoS902PWFhBobWwP2OlBTLAPB2/PubMWPlB3fw2cLFhJDO/UKrh
IxOmbfOgYQcnCLcF/XnpeiLJTc/lG/j8BO+ya2lwM/YpiPXzldV1AK1nHNWh7nUG
794+ybF72VOw0Co7LwfBN5RFArryLbi6xSk/NjPvuLb3nS6oab2I/TSBoBOLX6Fo
x+ZsyWBWCxMcSLQdYr0WGoU+IDH5FuOzty2LutF8ML9r23Dq4QUcVxdjlvaVUTP9
ydoKj2IbrgBUwR2yXY2CP/oKkzpPxP15Go0auwlt8uSX2rQ11qv4LuTSwctWZhxV
IuDEBWsUQ08AMetv3c066YvdU+6E1QNiJD+k/FVg2oenK7fYbjm8LSBsB436uptx
8OmktpZTKEUFm/HTSI0PN7kkIqa/1giGeB9Qp7ZcAI6jpAv67yrfGGdexQ9y+owd
JjB9ldUyau4mBCQ15ZCHFlK7SepJxZPdFYalbqFdmPOkEAw+6nG+RHQsu3uTJN2r
63IH8NhYYM8pBM0hGjI0RLjsR/6M7YMIsZgzxKaGz3jImmogJBRp1gLvAokFocjH
CUkI0wvJ89JdASByKGiA4Ky7/Or8pxjFbIJZMcXaJC/cRkoBy6h3ZLNE6BIGGT6X
rAPAZErGVlgHiS1WrrP5y+91tGxe61AXi2Gt6E/PHmb6L3d8yMtwn42YTm/JdWAr
Yg+QolUWt9qmk3Dh+C40th2JWVPVEm0/gyq6zk2jJFzQcUgjDxx/u2y2nMmiTGrs
f26WYHdi+WFZddtya1VlA4TIE4eUL/0TYnxh06uKr/+5rZ4BrenlG1VplGElxIaQ
XNLrgiKMhkPUoDzsUY0L0Sh/2bUzLM+91qVgkz6sQXQrTSn00fj/kOwHnOR7Lc+2
P1ZdQNc+0CyUGfeug91Erj7P64dg6mc7/TxKNi58yOuS2AYQ/QUonzvmkd+/MaZm
CO4f2xw0g630dvIfUVE6I/m35GhSZUgNjVxhM0dNSRrLmwPqyCv6HVE/Iq4n4apH
Z9ixpGtKrf62w8VVtkh6elYcZKD2xRTjh5IyxE4pYVYWzHI1+mUeJxq2HY8KpjFp
tevfyTraq7MByJtQEQIovTmgR6lh9tXwSx8NU8MsC88sHPkw7fZRbf75IBSOngH0
VPiNrT/O1Zwl8sIBGgGVHm1nbwq1eg5m9WgTyoxJe1hF3NVyedbtn5AiwE589Au9
iIP1uKxEVGdwe8Aqu1nQMFBaa0m/9FGsYG2XAvA+F3xqRWqDYg4ABmbUeSXlDovE
+w7npT/Gbth7vDpIA6QPiB7yds6Hkc9zaoztwLriADac9cF1jiEU68SOGAgdtkSu
ehENwUACp8j6C/PAoZ4YXQVeiOv7CXo2Jmk/TehezTpxfiHM9Rt5aNrfV1IJEGlT
RkWAsu1rMnV8td7wTku6qMgEbpjpo9wVtxiwz6AFbgTKBs3dg++4bLmHyXchvLxx
PcaCXG4IcnZKl2xxyhwKpJ3z9nacr7YIQII7lHuoo50HXUR7rEJeNnQpuFLK778X
4wxakFurkCU68yUaOrnBBjiKoXnQQdeK7VlHRRz5feSLXdGPK5/mxxUW6VkWuh3I
cBeMrh02ZRH1GmUUF6CEPhgXddQ5/leU95ordEZT2GlrfBFNGL6SMP4xTceiVabM
0UGAnP2zIasKroSS2Nxrh2ifq4rZC9qqOmy4ebHDEpWNEh+69JlH3mUvz+9kqiEf
aUI7gVt+Y9FbACVWyWVjmeut33Y4po/AwEtM4akLrhFdSiNNbvdtvpU5uOCjptlJ
NrNKNherHgJ8ac3EPA2WEfapjQPHBvcesR8Ip/1o7mOdZppFAxpQYKw9cXQY3dRY
MgZKMyhK/41kxiKHHDk1vTg4W0SlxetZ2vT8SOsu/OhiJgy3SRq2Jib7mzp4cp5v
WiBYTptdNuZglLIfniqAYoOtytLBl5cIaXQ6RGy1tmqntnMzNOXCnLJ530/RcMam
NfWfYsnJ1d3WcXL8lWhV5nKOokkRvSSyZAfFKfewwFuwn3vMWU0vU+bxptWGno5F
YqGlpUaXCQ/1rodsPgJIweVG/SKlDzFZhWqSeojU/tsUskT7L4UUCUA5CZVaOTgE
A2xFH7emA1ynjRkuQTG2Q4oBNp+ZR434ueii2q0LWpPEf8PtZ06+4DSDv6yscmsG
3Tou0UgrY7FK/me2qhh5KFApPRUemr77m1zQZh8gpwJTBYlKDAiqOyUPrMd4gGi6
09Uo1S4gxf/fFaCVPnOlBn1fAbDu0JEz/zpTohB7SXgCSWj3RTpZgUQx3NBMtKpP
CayLMilwKIuWyQgXpT70xseREc023ls96xNul3Z+1vFi8hOO3myncyd1oW8vFFEY
1u30skGE5rPsZ9kQHnf0ua0NY7vHjIKiea0n5T2DBqadw+7axs67s5UumxSHl6v0
6BecflO+iF7B1eyz2aDyp751ztOaRn/dcy1fEk7hDDKKlc+LSPACBQmupujX84Yz
zRX+j8d0pClk1YeMJivZGNDLVQNd3BAWd0Ilsvst0Vq0cBIqgWykjpMHhVd0vTyh
n+St/G857anHekNTVlLhLGIjawhL0yM1IvEMelaN0iryztRV5MNr/takO2iu646/
q0PBzeyiFBiO3zI2yefDLIwwkDmZ+A1ObpMI4vi1sjediUnm3P3W/dZMx7M8Mzvm
TkTaw45tfg+XQ6cqCBOo8M9wycvQYL6EETEtIUkiSMexhOWB2kWGz3/0LmvyROsb
Q05n30y/NgOmFSRxa2rXUnpChgzEae1lZGZp+SIM9+rq+NFWy4kUIXXVtrpsSwcm
qXtcUxHdvaYfET+Pdxy2vVQJNAEXWWnrTroTThMurotkYZQRm+fIyXHqfsHsGiD1
7pooMHdGN8bzeKxH3R6jyrXPPcv+XVEgZxCsKGme9SocLz1lTnYF+IqXoGDmGLo1
1w8PRkDbz5rvc0oc2v5PUhFrP5YfvVzkSAYJ/O5y35lnZN60OHsA86yJ68ZSs3lA
lPRRpKri/53IM5Nv855LoABRJrrfIvjtMkRkwEs8Bz0kUBaXfC+STK85r0H2FXF6
EW4PGy9Jrg1V6L1Fggl229rTWLCk2YWPvZ3qXncKfQQR2M7wZV0KB9qXq/pWx+AQ
cNkHOkPAVLVgmeTUYdB510a25P9+GNYgw5DBmf0Msfr98h0CcYXIf5MBZvLPmOOQ
fb/etAqyvSMdapkwnfJDh1UmJZvkIMoxJils4B8/Xcq81k0MKdDiNbrK248BdZ0S
+O4S3p5hY1NTV2hlvSVOcgFdbYkdy2wgS/yZGVJn+/l5+6FRf5gW4407uZCQtRNB
6MIrL6y1w/yeHDn7KMSUqTBwC/HbrVKaqzgwT+raZlOCKdum4cdZlD5xAqhfx8Pk
kKlQfoz/kokwU4DNldSKTep2eg8oJI/VOIxhtRvLla00iIcGw9pzE4megRonxpGy
0Sf5UMfVgm+KJZ6bz3jR/grA09GuAWo2LlsEJUBj8p7V02f3fKMPKDB4Boyw/DX/
k0eNAGBGTcy+tKierO3hjoEpiPsEOAqfoyd0DBYkyixX0x/RXXxKdiPtr0OZj+IU
jvFKiP+VfZYKyHvwzkvJIf4Cwr6KHp6jr6USaaB6bo4L4EQuHMnvPpNlAySOz5D1
1PEUCylRuws1s2uEWamX+J4rhYsLppxWuZWXiTiCDdBVCth7f7TJYTENTxcCJ4LN
AGf2nufCMv7T0EcoSnPTRCzxL7FkAy74AX9KZ3qBvOttnqxdAg9Gr9Ggjz4zqeyn
FIvRcgspo9r8XoJFo1vKjvrhFIqLdFfpj4C/t40tfeT9/dn6bBEEBIFMaLUrlbqc
SlryLU6hoQ4AhOnDr7bBnsyOIjVw0f/EpV2pQP6M6TOG5oQ1gok4GcX2klgVuSZ5
dQxCYGj6c2PC2xqcL+Vhii6gBNZ71l9pGd6m+E/s9lBHPw5S6nYORfPuprgG7EIH
moQs5Kkrx7sxZCxH8HINWq4ExXamLOmw2WUT+GjRCjI3SvB8s6EbftieOMdbFivd
qi4Mz4aBWS2Z9VWRGHLg5UdmTt5sWi2yoRKy39/zXHrPE/0d7VfbeBuCnrZgcgcC
d9pnoBFzHO6IrqNp9RT/E7Ntr4L2mX4mh4t3rgWgNjZ40kKCX/kcxNpQsWYit0QM
hpdXPq7+y1d2CkM13xsBy5DgWPwCI8TEzBRyF0aG/tuUNuf/sulVIH0aRlXgWBLz
6WIRcLhlQyaU6IeaSZBhYUzVyAFLwDhOKDWgKo6Ri54c4ww/Mha6/sOSFnW+8BYD
IxV+ACValICl+X/u/gZRaxI1nxYoq09zJZUcpA7kxvkr938stiCK7o+pTdbxFct0
oYn6OQ77YeixXK05Y/PVrDAcckqvqHRXa9n8pp+f1iqHbR57J3BthkWfy6qjsEvk
+FdYURXQdDBaJLItB0NV7nnKMLj/k3CvSir7peXByLgJyvSWCynOb4NzaRCzDOfd
AFxtAeeOogatGOB89O8y9Rts8om6HaSZQC/Og5fFggnBehl97ITRYFAwGO4shKHo
GBnoBMh8w/6cOfqqFcfip92MYRynqydhV3RQQVTSkyhZnF6CfphTr7u+gAHAuXhC
5qoxKRr+s4MPoxZ/KVJvwImaYLXeneE8eIKM0hgCkWdiJhDRl8n3x7wUMtrkfMvH
TdDymRLscVTx+qAJXKr3yiOX9p5Zu+0UqItCXplJ9U7MNfXZatdf8tB9S8XFhu9S
t5Wi/4wnYiz15g9rT17NUxelAtnC8SxYapykJRWzq8IWfHdUXVjNzXmXB3G8jNFq
dwW8Nj9ORj9e/NdDJ0gSsVOoI5pBthpWrnc9rCtUKPXJxtIJGlF8Jm76/xG6rYXM
I5xK9a6XGOf6QDJv1fIImQacLtuDT1+wUMVe60ZKjpluGVADMIkSoq7oitOAW54O
IZhleztXhVaJS/vp61W1PFW3DQdTr2SOflbt0/hw8LXB0BeUP4yUWeZJjYIZMA5I
kcdWbL93bLeoLPXwJEWPL1pLByXiyFNn1hqJ/6QQ6R0C1MqSW5l5tyTQhXVsygk4
FXpEjthtSAx06t8h9P4q1K+VAYyTJaKDk32kmohu/R95CNExB86AI216EjgFUrir
3D8D5SkuMWXBfu75bs0iziN30bDmsPkhbCzZcoLfppt3yODCmN8y6T0KrZPjM61b
RrJbb6KDABo0pJYfTl5lj1odYYir8kedF8Xuu0DJr4ZCgksAZ8uXZruaA3o+LyQc
GBWpAzJegX1spKfwTu/T6BgN4CzPP/wGqalm3FQls75UkWp+Gj74TODPMyw/mH80
m0cLu/G5Phd7GsAjPZOsKVSY3Roy7FMTWA/FB5b4Q+l422ytCoWGfI5kvxsogXIi
bLkfncCPbRjKqYzpL1fYSo/+cLipcMgw+qnzRyxOfzUiiSSDp/p0AQhb6McOMqGj
TK08SWzmzWUVZo98Bv3Y9fNFXbsdq7euezQ16NTSwJhtLpGz+DObv1XPUzgLC0dV
dm4bv8MXHun/MohRZU0t8wkafvHhROK/uf7bUue8P+o277WXqS5SA602qlVVfvix
KoAoji117tkICeQOWlB1axvlaZwx5ALpWxsgAwFrAD8QgNLtUTEqGuKDpVFwgM4N
Qkt5lXe9pJQtaI673iZbRy4MCuVYcp7D1ZCMLonk1eD/eoH1wB1sMvLrXh8lq9F3
Ku8uxUXkBkHIENZjt40dsyxJ5077rgxShs1BfoDd2rJ3QpeA33Gd5eaPfC7xk9W+
4QxO0ekymAleo+y2UJIuydeQXGz887iEqSWnVEvKTn4AGu8BCRqOlhwMKYmCcIYv
on5GRn01Ap16v52HAgJTmaBkyqEyI1V2+AdZCkqQRy7Aoup8kl1CGSL6G/gmfzNj
9c7/Ky3iNarsfsBahjqC5unlFB8bKCmANPXTFUtstN0LiAEK2APLrjk02i65Xu6H
UcfWaPPwauXxyV3wMxAHH+bhMeSIwIjLuQHBfaGcszFRsLBT1dxKDMPyMv0ottwd
eugV7ntQ+HXDMQKw+6ZpdaxN/f1JUkrv/v4vSRYYasqKhNZXLjv6KZY+ZlXvUpVB
x0luTUlqUOiDwt/mzSfwJ9RAgqN6CM1Ne1UHdniQqfm3f2uDMEy5P6ohMI3RDpW8
UsTgkHEgPrJXJfBhWDfYl6nx8/lMA0INrezswzF/8vn+dZvkxBOgtYjCNx5sZZGA
lBamd2xJNQRrbXN+ErPFpxtKOwBnIKDX3Qlim+GPJ1neyORT98YKQiZ1b8eounbp
yCjvM4FrnULHU6RGAxH+NYhZJ2lajXhfH2KOhNbfAYLQQGHHTJmH3II8AbGLCpJ/
n17tlcQkgTTp/i0GgxIpJIQmsnzlFd25JVfs/GegYOtBwmyorADfEPhRGRjSNlAl
00OkI8TVyWqQdAL97ZVjv7+N7sp5w58bglcCYBfDwYqpKUK30wcZAWqBbol4SHZy
w3kobN8A2Wck+4MIcvoaEKGx/4urgHRDkjJc8coRq2E6jXH1xePYMZhY5c184/Bp
0a9+aB2cVwbbaIrfp7c2ofDUescVZnhq49kfc5u6fBFdZx2VV4+9JN05Z4Digg1L
H72PVy3ADdbKrFyq3KxQb3v01GExJ+KteqSAQZ2fwtB64e0yTblQ8z74wKmTRDaO
vO78fAYKIt3HAvxAFBkcF3OpMsizMH2ElgdHsnEySsuVl2CpvHjl7UmQIHLSa9Gm
9EdzbUdEFANGFEpApDPpYchGkpTIGsr4Z9QC2xf3GTA7VC2ei9OzBdarpTzqDnk2
EhKvEd4yDFs0B0zCaxZrzlOxtjjOuvTmylR8AiToJCIzvSMewHnhMnqmVU0skHsj
7LszJG2pHsgPaELii2Fgz/NOsmY61d++k/CJuPCVQBzH0pZUgo7vH2vjjnT0nGVm
Ezg/fYLvaYq9VtFRO3sZQmTyppvTjDVWCWAt64cbEOCON224jSL2BUb89mJM3RAg
lB6xmCl2UeNb8Ie4AAlPE4kUwL9WiIXn4F7VKAKdFWaqxisQh8JwxrLkCY4jVuBd
rfrAAUYgM7m9j8ziODdvAbDwXjLDMT56TylXXwKUhM2+USOmtpsU1eLL5E7etV3+
d0mQSe6MjNpoKtzdZHtS9WGSEFjXrtnmAWPVtIugKfMdEumY542/jiUf58MgcQVa
9EX2EWV+MNHZSAxBEW9kOKNNppdJhWrmPjE0P8rZlSJGBOp5scSanAj79X+ngHpR
p5CwN1KtBjEMAVY7ixlVziFN3kZMpEvCoZNR4Lnfz77HYLK521iV89Cs7/YTpeTg
P3Ms6+rJbMv/Au+I9RZNuQUcBM7S30832UTIQP3foRUBn84wrcAKmRCQ0SP/40mP
QjXaRZ3k81yMccZkoakIS+vfRcBsptOENrS8UDGxBmf//u7pKeZJbB9YRct/dBod
eZbbaxafbFJ2KG1LCqRgKXHB+tLN8XbLpfCIeLnKKbDz7ffOuUx3QPviACildyBq
LIqCRCs7x6AVM8+XwTCWz4pX16VmKtNp7bieZZTsG7Iehc0whmZ6f+P0SXv3UZsl
wZRdXam58Tbnn+HJAPVvsDQb+ecuLF+vyYaaiAWcVWXbQKN9+cqgOyBa+uOCdHed
AdrvfNxJt7y+egkgSg8rKh2qX7Og6qX54orn32SzEg1zsfNrHE2RSFulTkjbwwFE
mHFuOTyQeXlhERRTi92lSryNMBKNCmi8Eka84pykyvSAZDGlw1oXpO/nyKdnP44Z
Xl6UQS0HwJ6FkRq/sTyPzLhlWM1hwJZrILRm1Pfv4tNrNQtzMNpzYOulPGz0i8rm
4zYCPrLZFt7JbIOV2H16i/hCTboDGYs1IIWvuZRoGWZOrp65Wo42RSVeBhDLxsGa
WIF2W8/dhB6kadlXDju8Ks9Wo+Ut/LwQs+7f+Nx7pUy/9VPJZgfg4XTzF9Il8RaB
i01pe1noWBJhV6bBBVXPh1b9fvLnxm3MSGEMhljz+E7Ff4wfVxqbN1a1x2P/LLdB
IM/2neOCq1LMOkqmQTzeSDKi288G5JmqKmnInf7r8YP5Pwcp604o0SYdM4qQHmvM
QBDO2aGh8nTP68Kd19ev3jlgPKTPOjTPHZ4t6iMQ8tO+45j+NYcl7M+vUaggyWLj
7hdP7zIGjDhmewsjSp/jBGU+GeqS3EUrAwItk3+FNrFAcL+rtOpDOgMabR6LtIh3
wA49NI4xMlEv+e4lEQfgHtx6tP5rbpMg3n5LX3/45w/kE7KBKacAeeKTe1IoOtL7
/9JwIezvesNIcILRKNTDqN1GMTkZ25PH7Rg/KrvfXZ9ioyL4bJJ4NIkfY/1yQGra
0+IFMitMcNBd78gvaLQy+eYzRK/yzK2qzEzpJZNfNDPAIe/6VV0eUv7YxLx5rcur
XNQAeHBEoMuAagKlKla4ZQcxSoxDNA4VC3d/8vO8yHtdZwO3A6LSi9Q3r2a/+bOK
jhBDxGQND8A+qUyI6ubg8gOcTxolzy9W7npxH5JAJwn3vgzd3zHY2WC7g5/lCppA
zseRfmrFt+2NFw+xLKnIzzw2EzGgp8NSbzOY3EkL3aQ2xt2OSbDdcCkHTRL/RZTE
6N2JE+tBWt/Ov/n78mOTp1a/5OjNYrw4aZyaAYlFAXZ9LQUoga9ERKqVFZQ+6V2D
YohznhHzu0xdgR+yfIwXWUhUe7BX2oWaAaZ06Zw55mP+wYhQvhNDArO0pBXMgvGc
c/9m6fGq9SXpA+MGvcAMcmcIqdW5gyv6DhhF3bgDkghrTLmKwaqS3kEiuGBQifLN
63hgb+UM1HX+Z4NOrywEBUSHji0ISaqQEMzFzwOKJGRA4PaFzMDWMxCpzTchPB9M
z2CrJ2019jSWWTJt/LnIwHaAnSqzued5yfPvMVngryu6+vvAzbi0rIGSb1rgNERJ
8ayarkxu1NgCGVl2mqA7c/PjCXaArijQbxxkVXVpNLNZc6g8pmkpCUycn0O1BofT
atEl45/zZtBEENXZjmMqzQ8xjaN4eiSvP+zBaiHMseAR3fAlIwY7NTmOCNO5sfbK
dvxpy4pRePWNC1xKd7Ja+jKSc7bEb/2OxG4r0MNmLUGHrGZOM4qDO/J5ttXt5EOj
q3OA1lr93PRGnRf168XYGun4/Pu+isDZ7fAkCs1YMOiPthgrnFpB2Qw2xS1oc9Zz
tDAhs4MmODQ8O6/ha3NIOpahWitpCZ7E8flbo6EL/yE3yCwQcIi9xuAYY9FLOSij
eQB1cw6d8mnCwwDnEmN9tEmz0rNlo6pmtorH9JACy5E3i7TiVamoFrOPMKXCZLYH
Ke0ZYq1yeOMtM0//eEnPgp7xl3kf8n8Eer9DXZDHYgAEmT5M0YDVy87Yosgf82bn
e2GW4XyLIOQHMhYAXbZI17vetqJ+wvEmnZQh5FuKoHaBnF9d4eGSsLMiDowx0tLn
gXsgYK4PvhytN7t1VjBNyAsAypdgPkZRrO00nPubiMQ3ipkSSPbIyO1k9pMt/2g8
sSFmuLZ/dvf0yhnI5LW0YKqRVfhsTEHmd1TO3wLu1cThLc4wQc6O8YyN7ENdO8wC
ZSkIIHtyuVnsZ1jfUCNOAPuotK4EdLTLhP/ZN/O0uIwf289TQyc6396ueFJ5m2jD
cIq0+fNAlNTOnMW9NQY6cZpY/WOXBOi94OGfupsA+MK60vsTmiFojinr4y+ZEqfQ
9mAwKMwONhhIgDXIKA3mqawUPY2Kcw5dsDVZNv7aAmpI+NIEYlfeNmlcYbul6IHj
oINa0USWA7L+nST8qlaLEmYO4ZLurE1VVKyGwRuD1XcnD7MyDgo0AZfqk/eeFbNm
GlgMdZlDbhrVUsUTmarfLRbp/eLzK2ODdXOkfhd40M9H24UiI7D1aWNGTb3l5Y65
1EHJnr3mFC0uB1jyk8gypBjFEkcV4sJ+na8y3B7FDMOgWLupW6zdslBHpmXwvyz8
0rtZLJz0KdzJf5sEQRYE+z1lxe+v8qitWqZAj29+ZVRYxmF2kbnTLXZthyqKnnub
i5NOpyY5QTVGBwM2OyoybjdDZrmNyanroDnjsZbXwWLtIcPPFaIVTZV2eng7lZDW
Nn/TOZqQPghTMSgJ4AkmtCM+oJTGKsNtLpSpGZ2knkJwFLce04bi0TqKQB9eMCtN
DtVcyRt1EyvWNIrz4jvFaqu1S2Gbn1uR3Q7w2dY5B7hM5CjplcVfsIp1uTKXl5QS
UnDNs05v7fQ6FUaQYydFbfYtNSbCXhcsXQBxil5/h1feLi21LRS+/RomP+O2azYw
N2CdQgmdX85kQTsqS9MeXCSNGgFbTwRajpNBce1CtJUpofWqtvj1u4LrmVV6L4/Q
Kx1jWlTguFWj381EqLmywNic96X2S8HkczI5IiW7qpPp1R0c9sHTQ9H58lQEipym
7Mv/8IfT8ri9zXmko6JCyYnt6HKL/beLlmwbzqnbopqTskKuHxHNPQGFBgmF1Z5F
BeSlwV/VngktYY4v0n0+J7IvugsW9piHPfe9isqfEAwIsoSR8V2JaTbKcm5Vyt0v
oGeom8bz83CtPZJYGW4UlbxHzQ9brqgCigwmoNczIQrfIJoa0QBspIZYU1t75d2j
Z5y5lcbE7AftAs/s734gp8b1pKzzjfumH3VXn0SoA2AJshXGPyEMnv3KvV77Cde/
Sk24JSesse5zFAvIRC+xMuHxvIy49PHCa2vk8yEOwLDR49Wiov4DloquwWcafYs2
9Ow58pm2ihSCtcMxB/L98AYCI8bpas8+tQXczHCpMgDDDSBEbYeyosuTgRcs0E+P
rvzJDXXb1wEGANPdw02bt9kQfsI14Qyk7SkL4YfkTO2G13pjhEzjLw5NzNqo1D9O
xuN8g3FAySCSu6HNfhRWavQjUmPLnmr2VtFYqB0TOt2jIBsIa2gNxprjcIzObd76
KlhXGQcCVCI9VCDs8oZ+dBe2DaPVZrYztcEGjSQZBQ7EjIFsz4LwkeYbEs8Zbbd7
3Q/iVtyemPcXEkPinD2MW5My2EM4WlGLHwgGvBJxkcBt8DaMnwnRvqNL87dHhF8R
GPqXQlLXcbYWUx40TQs17qiGThkTr0Pld/Ko/6ANGhWmYU3jxxPAKUweUvLLgaFi
0dl3zBh+frbceTavdP0LHipWgS0jQBmaO2j+9MzRcz70+/x0BmAYUestbvMAqAiQ
GQglgvWgQ27ozL3NU9lbZ1Lla1rMKlNCYrkm5xCZ664QBPK5bpuC6wnaUUM5XaIS
ZxNEXJLKkpqFcFDCGWQ2lKcQU6rI+teglfougemdEH1Ag6wDF3b0IiEKDKdcxdaf
UnWN/cDIev/oWDwwwmpL0HG39HQ/gVQPP6beNewgYV1GYo3qM0KFN5dO/zx9YhyO
H624aI/BdUdPIZyaJQrEquiO6jpZt6KkNL/yjIf7R537CQaeLChjSzGNIKOpiWkW
Ns59ryCC/pGccs/+J0vLC9w3Qe6M6ukg8P5OWT08nF2vyjTJD5686tuDRM4GRfZ3
3OFRnG66IgNVNkGiDrPqZborYbQYpc4MoDO+9IhPL9dayRB3pk5xLCfpuTLOuuM4
faWtO5gSgZZnvT3nUWb/tk3jODdJGM5KJoC58aCwhNHn6XlEmadeByG0mV+PmTBd
olnL3vBtP9o3Z/mXXh3VX7MDu2d83q4G/WJvNWyStbtwMVoPcmwwy3kdbqVMrcS1
Z2rHU5e+1ejUe+Fcsqf3a1x3fVoDff/StiLslyDcZbr2/IP7Gr+PwfHrEX8xpRhd
xuD0ZCNDm4mP4+XmKk5LuDnkgDBfqdHJrqkYrQjo00Z4kkSve6WZr4GK2N+zEZx/
Hk2Ue0ZgmrWbTleLT/RMnvlvVD3cwbBJgincX1Rj2P0w4eMXEY998Au90yM0N56y
Xih/vF3k4qEXJNwr/x/4JQ2HYumyOyfl6gC4Sx0LDKNjJU1XVOm4+uX1wmPKUEES
C+CFAEr5wcoEv/wk3EPersWoAElws7UKgeHEGdBrst/M6Og+/zizfY1Ll6PrHWCd
L7yXwlAJn+RDiFBPHl4jH8tWBYYFJp+KEFvesu1eCmDd/Xe39EN4vAvVxcecQhZ9
g3gS/toZO6jaL+eRGpAZx+a3WxLN/VtA3nFPihsbw2ROVPVr5Z0em8PmeBP+0dhw
qibCB8HoncXC55aOF4e4/x95y7TN357wvVM9PSbxWG7l6t6ebjTYdZnV7h3YoJWw
DHhVvDlEUEWfwc8K/99+vP0DGCQyx42p0m/aVMqmTmoyG7ygcWtLywQq9COfVRMH
K7C6eof1sSQPnWHe83q1cM4PsJT4V+GnHXonsxHsRo1EwU5maFe5GXPmhrq7XREE
I1uZaYXpB2EwvgVzFsN/mmfD3uPvrbd9x6VWk7vCn+3K3DIQD5eV0ks+X2aqC+tK
UGzeMHN+yag/YCVVPjj9z8Kcsg3wwA/WXG7RKdhFvUYr4U/ofJGhzMpQjn+cUbl0
X9lyedS4uuz4J67Ls9lZxEZqEFrVklNslJj6baLcJ3azANu7faPXkUsVhlZS+sWn
EvhjFRpa4gHW+q4qTBzQLFBWik9UEE4Q/BhtyyeTd9YpQvllWv67fqEeUTwoF/nR
ta8KXo1OG1+TVr7cNSwl3zBRFnVzjli6z4dyYyX1YNpb6E6TPXqheNx5ul/ekeDG
Epi3msJhJdIJJeL3S1FhWCOEbRDtZ/h0VE3ADbSqrtFld4Eu2EpF5RZTt0YeTzqy
AVMq7VDifY9rapoM/0BwKeSdfvyH6GiD28QLbMsXwn5yhSICnBSDImHP6Z5npihu
towpWe5/leLnX/sW8TVs5FzMXhvtDLG7aIc8bv4IF4oCJq95fzw27dL8N56v1xCq
/TEboXxOZUCO1cP+khjZ4hl3e19pvrihKVIS7+8HCzTxyKjuFYO9vwevnwJy0jdo
tjH9b7/t9dJxlamBz0b4DdD2At0yy2inATlMzWyyPvCHVzAh6/tr4JrGG42S25Ce
d2oCrlNswQPe8pEkMkSPuTU0W4OoPcPk4V3onLJfBQHxXGQsJHmTC5ksKPv/l/E7
ZQN/RhBYd8Qf8b3rCMCsVisxXJN3ga2zlX01CZDzJ2djNDsEUnys/aE3OyXBOEzv
TiudnDJb3vJfabw2lMQj6CWJAT/viKtQAXbS5Wbxrpk4tQh/V4xDRyuyZOBYUEkh
zdDNlWUBlMyfw/pjEPuxV0iAbaQ6CHU1k43+1RljMVbb1Kx1mcaqowITAB6GBmbB
Nnhn7gbeq58sQLoBk34tFBUoLZEzRgQgEsn9Z/Xc6UOkP+eCqfXXB4qRQIzVApsN
F6A2YpfHzTkR9wcvLzVER439BwNIV/l8P5ZOSTgSBVOAjx42mLTQ3BsxSbySu4ze
TehS6Gl8TecIlxOgYr0zUL7gB2dv39x9ddTzTanjVbEA9t345r28gfpa35N8KLgt
zATfEamw+WWQa/nH+0GFxlWalSpncUu601FrLRFtocG4JZcH+jsvq89Q3PY63QgN
dJUsLnDh7P2Nc64VAl3z3JIuEwUiSED5TinQlKv90qWlFKrvfC6DIROyjHQx3O+E
bfr+5ELqh1VoCFEsI8pTDTOBdq3CWo+VMBLhqme1ympag+0oz/ffE4y8ffeoKyJn
hSESdxqPAMa/FOFvejfDVzRgF7SaUQ3NncPEUm26/oDdemGNYoVWGgKSlqB94uz3
037yScJZk052YSx7zWo0uLvdT4yNOnZfBZdJQoO8GhGhekt4BNr+MYAbX0Dtcu3B
wij5JF5PA5o81SlXx8Ik1Ucb344K+4X8X6wqTleKeEvpK7DV28yALzvI9nr3x+Br
3Aw1MTRJvdP3N4giuxh6oEXsBG96L1wbrAzKIMRLswsuqhG7fo2r9m+NkhcW9W3T
g+D65sVrE2F9BcD4z8V/Jn0cTKOoA3/vQbDyccyKJdKQhYbT/ITbksiGMrhMMVYq
1dJ3N1u2rz35chlQUzUanEQGhLZbdxGJA28pbAxy2KTlLobfeRplxDKRb+/eyPqe
ke7KDMr7BJQ1SiYOGhllpiqENLKfs3ytJ4PDTnTqNKBaNyE/xxV5dnP8FyM9MvYE
xuxoHSpvOVnivV1I7aP/tKt3/7naLaHyX+n1HN6iGyHEp9AhcwSg4qjaWiBfQ4bd
PH6OMGCtSnMbVw4oYFSQyi7wBpy5ba7OD3yk2SnZRqaS32Pp4NebK+L50RE4Kh1g
qG/FJOUFJIrdlDWT2YdHIHdwpQIK3AcqAxseJvK61EpZhLQrzgi4lhztyGD3umDE
zjqUbOfq+QWctX4jkO8jsBm5qLhIhqXbDDh611T2kMtYPsajqO+o5HxH1khs2OGw
yiy16IA9hbXZ9TUDyPhUYQbBj/W2vBFr6Xsv9Z0QXk1Tu5Y0kvBv3YYXnxT4p8Yj
mzWzuxlgFRkA5QzCiN3EgHB/atfpIz92YrtfW0PUTjOAf/Kwsq00LOGvwqayMnPz
wR9s5RFdWQ72abLLaQ0ylaomW7hHq3jMekn4fyi7r2yks0yfU3xbWAP6NnQPAs9D
H7cbNcKC8Um348+xAleVxaG//fnb+SWSBYAqNxBY/cEjhi+8+g6DQ2uFkeviUYkC
PZ30/Y6ukDgqYfOt4+oZRWIohDSz75XrpdQoc++WHnu0IM4ojWHrupLXRt+rxUF0
8T2B/CxFKiibHCiwoXWROUWHS1Bp8ZT+hRT2XAdO0CU9M0nfDArulLmLKViCUGqW
/B+ThardrNhjCaRw1naEr9k6dbOzYJqT2RBytDJ513Ntp//unrtPftzKRGgQEBoU
6oiquHHOZ6T1um7t901CZ4xfkRVGVp8wX5rxEP/IFgE2y+iGXEsV28P5ZkxwjvnM
1xPqLGsLt4Mdv+H/scD2NopItGT5yfySHjNtaAmWr+ozQExbA71lzLSTwOo04FM9
DiPjZsW/AUw2g5e7R5v6/fEsz9z6RjkaSbHXd0TWcxq70FOv1hGCvO3HK5s3nNiG
Db0aXh6g5PoGMNEblNgGCIz6/rIBTTaKxhlfQIB3I6lFYJ+FJ05ukbbP/tDa+2p6
2eb1xmFT8Tls5HHWXYZs5L91/ZmVj3Ot2bjB7Ix5x6Lw7HnrXzHPGJS18eLo2kqK
jwEX9ae4sqP0esfqCY5Z5J3qfdiUOm4l0VUB7l2r0B7XvGuEHSxEFY2CzhM4PI7z
XAssbDGNgK5CiJGLxsM/0cxmi+e0IEIz7vj35fWsg5K3pRZ3UH3oVq2gRJX07AvH
jHQ74SgOwRN80zE3JKkSiXvk5vP+MnIwTpOc/+vhIRnwkikckPWwF+RSlvA6MfX1
jT+jFrKfVLiLS1pCvA1YmpGSec4uJxXbWucrXICRCZZdIZTk2mINnm6bGJ0bgLRD
hfPsbfO4DRlTAYJaug6mG3s5gOulhMHGMgFZNc7ZB9n7I7Ii7VV7RzJeyHflV8BE
dvO1D4DAgQOKWg/Qmgwc9ymATJo4CAXyZvea3KznEWJcLE9lUmR59P0AFhwI2do6
YOhzM4cbF9mJPULbwLsBcid2EHPMluSGtxD35MUhE+LP79j+BkzJ059XRtNinbkT
Y5Vmht3gbbFR+w7YZGndTHTdrG0JDGEArZz5lh/URGkQf1scsBxm3RZxiNp2Yezl
Vm4MvgAAaNRwX6gBfcJk5e9KSFEikHYsCiryPfUfhlaC0gYb1PfKj+SmVwGJEcTA
NYrRyT+8cfg5nC+QIA7ccGUi6SXgsmmLHo/eOW/AOc38EIHMgh/5ivJhsuP69KHm
QCPBVxK+1x+jTvcu4F3GCmhDPMY1VKvBeyEV7UBU05xH6LwDvUfKgJ0Skah7Xswj
6a4m4m1ZgGbCrnDNAUMIGun+bUf+cy8XmXU+Ic+C0KO7S9Tcl55oTvckJmfxKRQK
y12yZ0LH6Pf2T9XTIcpC/Wo6Bm2BllK7Zg+flBLNkPl3eHzbSGR4Lvk002+1S9GM
ijl20PEgEXi8B2gW9tzYGtSoinfU8AT1P8Z2bCxrUji7i+ds9v3/QFWc/omEXfm8
qUBcO1a89tAY0PPOr+7NdZgGHiWEKh6o5bEvbVFavenAqKFaR2sag58iEACBgKdV
eJtYlyDnwax+aUQsv/y6GgU5tIRQzpO+b+UHZFcmhbEgQyjhPCNTH1a9NklVR1z3
JLycjNGPpsa6Tol1MY4mS3hbT1QBQujyYNW5/pMSg87HymFI/K8RpUzh63zM8KAq
NtlmOeqsuT9E/vJfgPPQWnKBWWhhpEkMwIGkYEtrmnrIqpadjPmz6OcNAdG7/epv
MyGPOg8w5WjVaQ13+yoiAlPSUSRBjTVtxwQPlULyZ7xp8WmrXyOswemXxqIM7dct
6ALmL1TAhDiACgNazBkJz4cFRwGfsMMKkkZl/Dlt7WCityPZfPNA09L2HXeS7hHl
cXNpXV11g8qjhB4PFLP/0rAxBgbZKUa7LwVUQF4OiY3iQrvtwCNk/h+9SBgzS17f
Y+46Xi0dCqQX9QvrNH9EF+2ifFJOxPAKskkLOhWFjQvYtLWFkharcDwDSdcuRayV
SIIkDTn1rBJuOhVvL/kNM8rk9ESeNvJc5m39kQ+9W/Pn1vrApc07G2jtO1hVXvRR
tCyPejGKo9Z2USNFqn17bohYaMT5RZp1oRM8Se2FEY32Gi+ircgOOfw3ljsSleA5
gDLZ80IAYOcVq2izI0/GKN1UbxPROIJq3JJhnwlDJ2mLhcb9TR9qVIFhj7q0Ajp/
bILJz5piGr+PCJn0EQ81SLtSLapyFLHgLQ1BrHtFt48UQjbBL8Cyy0AnEiCuqR1O
mzOAGZSUV6Ww4jvoD3FrtH9qwA3rtOe1aycqeQ78DLAZ2vkZ2NZGMyzfZwN0U26I
FobsBFduSIIxrEhbn7XwT2VfRMO1LgUDyaQql/I3HL2uYxOAFDOaY0Rz/mE3WMEu
N73pTGvYNm5U9vi90t4uEqQ8qjM+6kvF9CpoRfXihNlgZsBhuCjfESGJNIU2lPiF
FI5yyh1UoyKWxXv3dcet1BWZYkA6dXZmtSM6r5oPTsNU1IRJZklzrBB4MSHTKLhu
rhGRRTG9ui2C+Fxx7Lkl7Iw0WweOEYyUOqUT/PqEnLN5o492bWpYAIl80+tA3IUC
hfB3Er60xiZnLxbLwQIH87HFr6cPQCro+aS39GrdSBajXKTLRtQH6Pd+ORm+wl8c
MUMtYKBdB1bVLPBaG00hXRW2zEVA6OnqaSp/ueGjwLxDTeQlgH7Gj4/WH+YwNltN
grfiQsGf7rLOcUMCYMAIquuSkCjevPtMwngxljx+OpI0YOBKnWJ4qViR+0uzzyE9
7DZNt+YcfCHnPIIjlTkmBW6f8KCIozdm7zTOuvFT5EvRZJwcpBemrYgu6n3pgOXN
HQHaJRfzrsZ7DHGXP6ZUWRUAMcx8LnWXNJmqIbWbuaDKMdx17tu/nz/jWkN4UWVN
K4wC6BhuvkhD+qe/lSeLbxqpLBoQAgZCT4uruheIPFfVr+eAKnnYDcr6Zbw9az+8
AOyMNftkDJdbnGo7UtcepxkJdel+uS81SFBIUa93/5gaW70wHgM6n3JWzKUkYAwM
GN9G3xGd3qtZ2GAmVvzj4PzClW0vp9xI864rYX4c9ucssU3H8iNQ19pFQ66lFcVj
9O/NIQKpO3Y/dcXNkGwiY8JgbvCh3PVPIH7tSl5kSkEcmc80wYjRBixYDBtIEUc0
tACEI7wEUlmTMiJZ83Dz8zVGJtJ+EMN2B+jviIJzTTtXYoFwzBuYPVtirrHm4lzf
XHTzekB+19/Gl+DHWvx9PdbVidtjruK/at0t+3lPGaHWmDBW20PnJ1wr+L9OPiR7
PUsIhNCc9pvtDTBlFxdehotJk43K8EBAJSl7fXf4sqUdX7Pw4uRcWh/tRkdNyOLw
WXbjdbxnoaY1oXWtBfsXNGiBwZ13Ej1SPRpaPkJlVFeU38UCAI4KXhzUIkUDpIbu
M5hLNC62J1bPTBJy7wE7wC3hg4oWPw0WzA4nrsRQImlsVe6bxpy1zrkyWdQnt/ja
dtGpIXo/vRIvoAcXy2rNKf5mvQMh8YlhssrsLnDvQe7G9DosknbELDUqQrXLmrY8
+gnQjvxpkrqS1KtCZgzXgfDJSbZJgUFSLxfRSz2gWLLvgf6JnBM66TmHJZRcjmWv
+jFiqSfWqGVTrlpNHaKISEF6thUE8/VBDFjwg3LFGIvcpV35ChtXWCXsI0Q7NX+4
wX1pi9hBFwJNfbmdCybFdefH5DAox4LxjWtFt/hyqr2hendnmPXO9uEbVxhkGZYn
6czx6bCE2QO56y9slXVSL4pzDYGtSLEmJ8OXbvXxeaDpnqWUw7mfjp44nuwSNBnv
DQKyi8vn3+46xeuxwsn+irmqRYMAazWlrHb1GceGEvLWYMYvYmPECKy6RGDoFfB7
HgI5PGZOP64FRHwGq9+dZZRHO8qEu8GnRX4kZt2tOenKrryhLPUlR34WVf6UseHa
jsm6Av9t40PWSzuqWx0hLZIMa/DNll+8peMzWcFNSbHnUYJ7q6L8s8UjwOqKakN0
NXmAO8gZK4bm7BpiBDpWLTGVsdJWKlWxaftza5rghgqrvS6RPnvJMNOWAojIMPtI
NawRe/pLo5mvMiLYCHicL95oFB9u4ZD4YSERUoPjlI/CIpaWoI75fJCgrNWjTM74
ZUytqVDo8dgCmCi+GImuJ3WFEbeJflKfvv9f2RPFbuZGLqpQZ4mBBDNZJNDy5RWS
+201hvD/Xf43XS7MShICWJe0YwpHBYMzQ9RcNttWJ27ykaMRFDKCYLOj5uCJ2RWt
Q1M4N1IWNFyUBtTwd677K7Gv1spToS+nah5w0QFm1/1wASVWbfQZGnpmMKZWyWmZ
+DyWrSHQ52FYXtNPAmr73PLcnni0bkMLpkB3RVItMPfgiVPDTfCTNkC978GFlaj3
hZeotWG0RxLXaGp9CoP3r4L8MWeTTW7+8Q37jLw7S2Sclz7TTpTw58njduMvtmFB
mXUvIU1CKomAfaRXrlY+7ij4VBrUCz0SUQydzETdNdr9bpk/Bf+LTyNgriYJOn3i
2+6hyII8h/i2SKcTsxZv+bXI3u1ewqIHuqgPdseKR3r92h6k7WN51lkSk1SQcAPY
Zfxp49TGJCC4l3ORVyTWMUkz2+9FmjRCDO0DDAues+qO5SzyQoKkCUfhMlU+SUWM
AJ+khTEQmUDnIIAAi6dKQ+Zeh0liCMOKzrH+Pu6YfgQ7TG9CivtAwsDLwtVZUZyQ
JUm9PCZpkvCgQrDrDp+kciu1Kisn1b6BgAAXEcUdvD0rcPSILuMACHc0rLJe4ghd
7f96B2ll5rp0ZnGY6HI9yWFBThxbyjuq71YfPb0CpXEgIa9px2mgKIXFUfU813jd
IjUA5Jz46s5fUHEopBpSqFfmxsjixsHOR97nzs9lUcc0sv8e6asNlX6xlAhSrZny
T0uZkDzz4SCQXAA0OWYH218z1FN/HQuDMAciIzFjEbEk4mBD6huUH2Dh5j08Iz81
IPz2MLu8BEjnKLWXa3DHG9bA3/+mNQd/21HPtBvn8lzfjE2vi9AHNUXYygiMbZug
5DLvplAFl3lL/9ZV5DQKZmD8He9uDA7chjCgVdk/uyStpSb7Jj8gN5fCh7QWPewX
AOt/DuZgcKRyQhtp0J4nSflo57nBpOO8TF0whztr14hZce2tOP/buohofjA9Tqob
A76KBmlhfWpZWWHu0YJaKGK99xxWvXejKcwpPexTv0SnCQ8y403HxEaFBR+tRU8n
hJFRAWfnlCXfp3YrWiosxmuz9mvNCN3lhNsaUqkeaoO65AcfEjEQ0oTTvo73Ma//
gyliRrVaZi7BrXw8TlH9MXQo37a2M2rMciUHka4UcuKzdP7IWc1ryPqWJWSmHzbU
169fQj7np+Q5EGZ0cS5nZe0LDXqS8NMKEg6OX8MB619Mx/UpCI4C5mEOBNjTxmah
mgxStmbNUG17NjZWdq9jGNGIETo8+VPMRFJFAyUcNooSsC77q9Ih3qSfbOD8zPlD
AC5RNnRz21BOK8P6addalJ4hC/G2CTLMsfHDGh81ZOLN6e4eDulRlkoJzCY+Fbfq
pikIQFnlm275nEo54fNzbDpHIBUbiS3lotEs61dFaE6twj8B7XhzBLG4XgnfLXbX
8FbRfcO8lsrJdl67Xjhmv2JXCqsKo4qqwfGLOjL/2J3rW1KWeKgkh29xYurmXMHb
rWGEcd0vpLodD1lAlcpqjA1K2rOrWFA22E53EcRUOXw5F6Uo3Y6I2aOxddx6Acky
YH2kKwTRzUjDgvtAUoQAXj9ES8xnNJnyGI66fRY6cpwvEO086PpBTaKWraMu3n19
SZTjS1vovBwkRRyLgwQueEnKPH9R+2WQWVquDo+1sLVTM6SLcVKok32LLp691vFM
px6cWAD3XkgCdH72edxIr3GY2M6NMX4pk6qNsY6Ri4QbGpp7R7dp3QZVcFcBunXF
Q2dmUpR+zPLVPMx6Y15qjTCul2jUxUFxuHwgp77oftcbG3ctNuFZwx+q3Wz5Sy/Q
djd000rVQz/H6aAdzniHo3RJj89fHtK7LCA2oWxQdJ05MUL+8rT+l2c868TxgPSg
zbE93ZC3dxpUQ+bLWmILo98ePNiA03SscGQq7X2mApa+CIOEi9dbwqrGjo1C7xAP
flZ/QblaSvC9oxQ4xau38ySa/UTCwVM2PT7duZQBPpFmNAowQhOS/o/kXNfZpW6v
C3IxG9lSi4eu8kL+CcrxN/gu/a/Tv+bOzRzFJuU53Piv1K0XNt71ejXpH9RXNy4f
OYgyEwLlCPGvQ6OmVYVwqlW9nM2byBB9XpBQz80HTZhzdUeYVDFPdOV2Pnzb6g/Z
38mlyYzJM40E/0Peqj5n8CR572b9bwNQy3MJtOw0tGPVHB+xttEvsK/QMOouoAbt
BscxRSkxcdentRbRCohu9k4qtLMUtg9EPs/YWk7nB0v7N6Z97yZbIxpXZuemgLud
sdgiuqJeKDhjiOOklEKMzRPjpbFvrq+lFHMgmXd3WvGtsKMCYlgtw90HUlAef/EH
uuQgL9f5WTC02EgGk0CHAy7gGHDbkK+i2lRFgoNRrLGVqqKKbimAGNu41rblnjEW
y6KGkJkQKcdlqoF/TBMD1Q0Ex3WsOCoISHvc8eDrzz8tTvnAuL1dk5DRu3cLH8a/
34g7tZHSlqp3U2+GCYtSru2StM1lueXsmzRfEGSvOEuksqKfWwuu4+XFjAYOK5ih
WWOBUT5a8/oLc9smPKlkUzZJuTlpxWJ0iWm+hJHrqOwgd6W1D0r8GCW8fktV5LLf
`pragma protect end_protected
