// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 13:57:46 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
B6oNvB5HBKpxEcHoQEL6XLgqPVl/Sv7gr/d8mcwO7JBA0J92O8e3KavBc1p3fJNc
1Ie4b33X0LU+gopYP5pBKVk+3zm6b1F7dm7+WMBOWvEkT/Yg+N3+ufU6tpdOvnCi
gOgRcEl440sempFkAiomK0KZClmzuUDyZGGujOe3wUg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5744)
+vd7O2u9Edhwm8rTuALvjvX4rh+gr+lEwslObGZO+PvlKP279sRYP6Y/lCnDhRLO
RwC82GQNSl0nflONF9h3aBAWsZBCLhLQmxqy4r8vlgEMHlTBQURIu1dolrDH+LQG
3QR+EQm20JLrgVRtcS0lgAti/7IJnnCbuj9dEQgVcjFuBkhh5bEWdkasr2nmmEpz
5iEvsrlvh93dOp5pPrDQd7sG14rF0SqJwAlZr98OKE/A0sw9rYTXtlq/4yGjK0u2
ZEFHuidWhDreoYvL6rKcAEjiJ3Wkk58sJ9BeMyopRGMgP249JCWaX+0xlEXKAXpt
ZbKBwqs89hl2kzWI2LLSenIfJH3ZtqTvLxEHn5kLceP6ZAYOFVMR/tnv5fMGHu61
0DitYIGOIe5XnkUH6Do4h9goKElh5xtftDK7m9y2apri1pu+Fs7f2PaVYiaHWfG3
fVB5KLZC3sN6tiDXBHaHJAvDG5R0O+rX4nWIIfxbffcheNMDnkkQ3X0fjwYxMMCU
H7lj80E54WSM+IB4tGQ17Qi2vlgpoCLEGCxalnNXR5M0VEySWa1OlVn1ugyQhEo4
w360eq4A/d/2HQurUYSggDf7pITTN9O4jLOK+ptS17RisudtWFKuwBMUuCbZ3XIj
fL6eQbMQf9W47rIi8QtDvHtQZSUqnFi/N/hOkrLfUMuVrFZDJqG1rWbbPRz5scSQ
tNaleeSDbk8uuI80Ctvkj7UqqWvUf+ygMPK1spxwr2dxpZpvezYH+awrKTmkIKxD
BJArR49Yn2b+mMpn5UAxagMxThbk/5fcKK4yLLTjd8iReMmAFFI0PD6CrmmGrcPc
r0nGPVq3UjeibFb6ZRnauHJJL4WcjkG8/LYrWlSuJwKPK7wTpRQmphtOeDVAvG0r
BuV3YlzakR45eMp2wwhkQlRW0CtfBTa3xvbeyiAH8fWIc48D9jYXHVUldp5TO12h
J5Z/Kjf/qYLtnPvuLX8HXd5ZCopkcquW6aeaUCXJiAU9NnfQNUD/05ojcs4/Ohga
AFrt1Zmh/DfsPmN+AchcNYBuIeBh9c0YF2JBm6mBMixrJeiR3Tdy82qr7uW1Tnr6
9s5KPQJ0zHgZKAGKv7+aZ9HEfuexZVNELZ7wxXCQZLwGkd+0J0UrG2s9v+gtE5dD
Ny9SVdSL0heSKsQ6JucQdB4gWimf40POsehr1ANGOO5Pkb9vE7z5unh43exso7cW
9mZiXsO23/LOsbhQuM3nMfvMC0Mb3boIP3McfO9ee4pIqCsPJRGSXMrP9ZPc3kgI
g8DYw7m4rQwgVNQPKiLbkJff49kaXSlPUWa4Q7YYS3BX1QJyI5f5P4BeC9lfSygA
YmdtQybe0MFnx6NsPkb8jRe3caDIC7gvw7lqkmr+uTwPs4csRUYFIbKDi5zqtTC3
D+iDOXvRQyus+eb6GprA9pUzTH6tVwPOM0SJUm9OoOi5GScBK77PHhYNubsduxw2
N9Gq0iAhziR3b3bk3h7uFEOaz7MLqrE+DjeEnm8k23sk0Jd1e9APyNZ5qqBPHGaM
1m+LD29LVcNU7WVDerExoYWYQQ9eFxpnkJ7r0FkTEWcT27kuwkg/Pz4caA4MuNLl
8sut8jf1UeWXWpi54ZcHHvmJHmolNawjbQUt2jx+LEaJ6wUz7ozaEWMNP1Z5WpBJ
DvjH797DkGpSjv093N+RzsBIi/Ob8+iVLDPkTyfZXxg2AMSYEssFyso6FZoFTEUN
BOqtw/zxVgUQU9leQviI6iyq4MemvV6b1VHlIML/DE48LOKXtkwUIdDQUlmIJ5oR
ahOGZhqsFrvqcpZH1seyNEGkAN4mvOehGV19G3iC4yBIrLPwDEbqVMhtXcwqabs5
QeaPnEn2M58P/UhhFMTLmH0eYeyUFY8jtFBQIh3RlBTnV8H7eemCAo6IUhpBvAze
9zdDptUYYqouKJ6Kxkk0eaZO+hWgeAbE+tPzC3fO4zJ5U6Z/pQrLbXxVSWytFZeE
YUxo/0Azl4+uDILiMyUpJVwDm5wTcj5QQzLELkRIlEpLaJr5tpn5ZruzZVB0k5lC
zfEGELxTAzfzoGCA0Pv1To12edNKfmoaJMXAz8j/KgXRAjB72KPEHr/5rDf98blo
QhEmg3liSyPT9xAsPOv0EhtX06lghcI9JUf9Y88MzZ1cq6+pPL9d1xSy1tRU8UBl
uuY22nsgGRJw3rA4/AOpOvIiaOCkEPJ/HhIcoUeOdYfJFtZ/jZKNxEgP7nsK5LvH
M/abu/zEbg0+VGtMxQg0Q2ic72AGoiK6OScVVL9rX+sLMOhy9uql0YbJH2ViLjlX
80qF/3F9ygx7sfoqNg4Kq4cUoCZg2NKc/0wouxYnJwUO99w4g6ewFLFwRHXf7bP6
uFqpMbxHMiR3NuXvcaKxKQYYJSEmheC8CTCCRah03MIUjF2hibjoSHNdPuHQgNFu
4e35F+opqn126spHypRr5XAeccTryc6WC2YSOnRR69WpDvVJMpA0ZzVQ4LcOOxW4
MrTy+GNZyqRsdrTta9FJcrKgCh92hs/NmXm60SvwHCaroCjE0IQlw3UVDrlGEULu
BRMhpAaGhKWY3M/GPijWllFK6L7NuwR+yKv11ZCC91fuJNa/Hc8E1hF/60xVIQFG
hT9EGgROXzTLV2hQYxNAEJDBJTNqztJdmfSEz0NmiKKmsZj1jPCH5OFw+YS6WTAB
XMqNv5IaM8XGkH2iWU3kieN3SKZSsxukE0GcxqUcL0ywFw+EIm5xAdb3PTvkqw+b
rH9V6PCPg2q39FRPIAdQYFve5Py9xD/HfWXRagq7ghMkJK8DaoviEEobvWgFZGz0
vrkF0DcaxFk1qY8xT1tHBOTFysifmE6LZDh5awUxFERtzc+N+HepiRiq48Zsl98z
KWPv1iHDOD/TIYDsYqtKoJPvMuwOHy6C9PnP2KQQdkR0X8I9EXk6QGLYT7x3TvLj
ioOqMLFnmDzA/qoVpBWp2tzI6a9f+q01nEAU8gI7s33aB5T2s9BXLWtxB5t2CzE6
ALTpcCNmy2QVWMCsbNHavcrV8Y/mUb9toAZSi7FDYFLkcB7k4kpgMF5q7xgSwbCR
2tI8o7Pr/n/a/BF+er4jfETpQ5wqf0KY9EOGHmOitYpEXyH8NdonLGr3UUMfKvGg
NLLRcjHBQxw1D1dINtl0CZIq8yjCTcDd+m7h+eAv0AEMexWyZWtjfydzUvQ1hTiw
pban4+4b3cRxbIpkR1Cpg+3aP5IX7Lp30h2FQTsUmLaybBXc4uSZAOJR19fYqIZm
UxosbEWklOoTx0ykdI6VFj9ao225p/VlRJiW2K1q+sUUsjxF6YJepu9EZ+pqEbHD
zQJrzaHdgRJColrTNG2fhg+/IDbz9QAT3Zzu192aX2uEXNHiB3E+4ARMDTaTnVSO
tT2BTXro6uBsrNLDpMyFHVNJuQ2lCzekUBo+Hy8TWSO+LrzS9RXByLzTwOiPAAF8
mYs42G1m2wKipLuLZ1B142Ro4vkr09T/muAmn7WNSZmj/JHUb2KRSfRDta866G9q
d5JtOuz1wpv93pLY638nLPru528kD4mFNKqvwlCRR5wzbgAE86l9xOPLcBQSaGEt
S3eHlOTmBPq4HYcYJYebGjIle8a7tQGakR0PcJsyGwgxJ0aWJUvAkdJFOn5gi8Jz
DjhctM56CciLrp3/NjUuR6KI84TgBxNrEKtXeOiFRjIDutqKjl4eJj4OXaj9ooa/
HFYMAzY1FjVEUY0XEFq594Uev3prQFGOfDBUWWDW6huo7kFbkMuCjwpEybTJkNgk
0LK3V57m50qcNDtz5xTiRnDlTM1+c5VjP84E0eElBpHShSxz+GZIFITJyJHoMP11
sP016IufZiG9Ct1WGhA/QQnVfyIXuW95sZ9T7Z+8iPUwySvhzHyKT8UAZUvUk0T6
4nnHiu5fnkxb+k0RHx1Zml32jHL3+FjYjlCVT5NBer2VnzNm38dbermvJRoVM0RX
DlGa4zfZHtr0n6uK+hV4X98cwKT8IpRxrR4ssbu1OxSeWMLbIRWqxIaOKO+tBnrF
kv7zWVVj9gnl98bRXtSEcLsBmBt7tswiWI41lYf6L3J9ivqy9Kg4tI2h4NFr3qSe
qustZnDxdAYo4AhEYSYnwJySzIsUjzJiOL8bV32aQ0laKhcRO37lMxPPYzP6+ZOb
PISwMQncT9gCdJFv52YGqBuqwoFUnZLzQwbcZS2Dfk3XgF7cGobuNDroZvbUy5fS
z+wZy7pDsWNKyPJuhrW7ddABoZMMugRM6kNWrIXuoia+WRsLbYxkdObqZegMl5gr
9Wk25T65HIzRPZFOUORKbADkBtQbPD7lSXuT+7E3cJwsVR9G6N/Bgcmm1/j9MLYQ
a8LcWFqhXxiysyND+elUn5nlWjKdEK/K5UGn+kHjoPg7YFxNMI644TM9dVcaBgey
5rc/dXJikgHe2jQFe5s3gvK4jeYBseAizc9kUB2UVAy0VevR7RYiEYxYbCkceG/h
NsgymgjMhDbcAVXHPUmlMScs09r5lEtiqtqP3OYS2wAXOXwnS934mcJcB0MDVtQF
+MMcfkhhY48PKmrOEG/zCZ5oHfpL85gvi+YU2PpCSvkrRZeaF65Eo75wyPQp5cXg
dOTuL+4T0kcjT9qGSvOxDz+56OqHlWUWOjUAOGliOJEhcvA3abKKfD1cNEU9lqUK
u9NM+WONhN/0cE2HFDE4Mh7X01aN/dq7gay7bXSIHh1W6LerctDoedvNp5JE+Ywl
86qhkilI75QnpMltJ8zvBVZQ9KU3wS/6tRefok4LZhQacDTaZ0P2cjWlNHT6hOOE
wPa5x4jePkhx/Z9aDpJWqoL6F8tM5LWn20Cm6SPzAq3XCastXcHFJ1O5IKu5cHVo
U7alntv5F1GqjvmudohIPe/x0CpDawUQiRlRq8aL/4Tocv4VgUun25DyJud+XKDO
loJMBAsMA3o1fZgZPLQuYIh/wrWH7dJDfjvwg4iqOrxqAjjOJPg/S3HE2fH8I7+p
UdGuo8pMKMNLVPE+Cijf//iPaG9VYAUMMY0OydWH6pu3zlp4I58IWHdd2w5PSFjN
RcHO/8FvDN4jNjKI5W3VeEjfVFnpj0T9CZ1he/IdMMqKv/q5rRlG/ztT7a9AYgkk
OTsQMNvoo4sTSIXJN7wDPhaVI+8zn0wzFu+FH9P4WsoNSUslNMbl4eXXLDo7nMVL
qe4XxsQ8Xr7x1qYdMoqQqjVYGJiHkXNojH8cFyTXpoLgcnTYpKwOllUZK3oUvmDc
Nosv9ZcfyF4rq78lEkCFVKXkkXrFxYwelGP7aQUzj3Jk8V3A4EYc7mST408H+rEA
mLIVKyajw+0W491vQDvKuzJJpUnbMJloN60N4TmmqAa4Hny+vMWkLrlSHr9DB1cv
qLlSB0Wn8Nfa+g2J/uoNEmVUPdRrMTEFkcjrqO+IHe012FY4QAtiX1P/70nZuJoz
TAloOshGsqSojSkzxMbhAtiIRhzdd7zygmiJbhyMRylc+KcDrL4gOgENOK39DMtv
23j7SNVSdU/jQaBqwJXMRlXkEJtecdXzb1Yj2io3oiIQwZCj09Hw95Spor2OYRar
ec4g+p5PGDmrRstnErblKZ+ruhyyMNqOJFSxXZ2yPQwCXltIRjb18f4EGecqj7qh
OLX0OTHDCYoC4k81aXd0agToKIXJMFDqynA+QiQhmR03GHpA1b5LDH0SBJm/+eNU
N6inY9UQdeLK2POLa3662Fc8ZfpNXlt//nlU4fPkRB8svUTUljvhAFd8jSozy6CN
FayELFj9zoIgaJQbZpD6gSXPt3JAsb50LyIGmXmjRadVJYx9bubthMr1YqixqwKR
Y+mIU1P19GXlV7WOpPx9ourXhIU076RHwEnEKYfDBA0qqld9OlVzy0jikH/qwf1j
sdXi1Ke7N0M3eAN7biJ02LmmDM21rFKQWpWnz0VNQm4/BpOxdAyS05JKOTf0UFFA
F6nbTGkgbVajis3rooopIYWYxjVIfo7cUJ7bR5Wal2+os+FYrkujXdBv+Tl7ciOh
hMkcuROIsGi+dWgvE71TZ0eJdZtEiqQy8Ug/lVj5uKCCYL+PuYNRtygQWYKlvolf
jYop9AHUdY/AKYwsigMQxLUK+BgPiSpqB4BQVqBmD/JTMSVAi1AaUlOUFbU4jq7i
HBR9nI9nglsw/aQ3+qrP+LV0EzJeGf4rBbKlz6AkfaxgZmK3JFejEEDduIC+iOjM
26xWa2W86TuSGXJllz9IPoe3/ic8z3/MKLZZ8MZYVTiFCmDtF/siOPUC/L1oHkvw
wgmZDMglTlkn8t0lkHxz2q5HlwwofYX312rYeouzQq2EOxngTe0jRHYcP3Kf1pn3
k9l3WYdbRaSS1B02ruJuC3XtekGIxczzVKFG8gWTvewgX90dUls4o/RWSes9TJFH
5YuwgGq/Q2+tbHqjZKfTgbhz79Y+zeUy4T0qjI1UoMFbU0XW7O3pXjt3tP3hjnwm
mStkBMcGfNrpDQ78kmdeQysjx5hcoIqMymldujIuYARyK5EqwK0s3UZFOa6gBUpD
ToYMIHq8omxFVgdN4JiO26akftj5At0jTyYGINh4Fiif+nRYd+VwiI0VeQkvyiT9
shuJ4oCLPeKLq20lttrlCFcJjSaqKWxMP7GEJ///9RPggg9LRfMKRwBTe5HHbvo7
MNWLPyEuyZUB6TeBPwC8SJw5JWZHRvDg9P1vDcx+nLxC36QCNyGNwO8tbLrdBiNH
zx8czHFsNjJiZ6CoYHrdXj+dtIdffFs3zMAscIHy9NfvlUC+3UCs0ftrEN8Lu/fy
iQ+Dbi0yKcs+bw7/raP1xK15JvGOZ9bVQJd78tVsJFjf5IhOF6fsc89GJPoJlZrf
bUa6Vo15TpjO4SfU2KAO9L7jajfMP4bnYeQsfdWOOckLAfMpWflEpt7jNgz1KR4P
SEkC9PV1MenWbK8UFL05PoCubQ3oR4aazAD9NGlZ4lehIxNTwDq95wNlHZLuvnUX
GBvXW6pzbNRLx/n5t/9yuUFFKe4p5EAc8qBlW+sCcvwj+RxSRQPBYMfoj/ovZjrw
oOR5kdinRow6jvEVaKuA9ralaF/JpdIUrMSPXXjLk08yWpousz5RfHd3UeDbHqzc
qxZGsioeI+Mlq6lSax2WJLIH8LglrfrOFQTX1TQR8ktzwUP6LE6gEdPVAhElz2p7
s7NY2Ci70Zh5gfmsg6vCw2c6JJzoF/eVp5i3QyQH8MAbtoEGT7SOw/GYXwqMVSFj
wVTDC/8JIXFw8eBGoBWTQ8MqFb2azrNzFPQKO1Ihbl9KTjk0Y1J5xbkElB9T0kxx
hhzhN1/z3pXeYlk5KYcAX3RVktsqsFofHox8SDggB/KMbbhNX0CIqfl8jk6KA++U
VbAQoGdbS5NmiVB42LvEi4gtBOlHOtZrWda4iORwqb0yRBuN4wKOgagG9keYXaNT
0y1DTvnDl1FRNObwF1vZI1YuOwCfYhgyX/vzStG1/nHuSJ/0tRZXn/iQ4ojUEBeT
T6/mlS8IbVSXOKzo9T8qXqjrH6WT1HziKiYsyaM0JP586i+IioGYrK56F1BoUspz
3cSIBJojyj67aHUcV4pqUlhO57oMXHWawh+KPcQZdPe2r2cF08Q6iIswJ9rceTk2
zFCMNX2+D9+hBoyLLEt17f6o1xA852liZ6cKjsG/I7s=
`pragma protect end_protected
