// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:41 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sPhn9hQqg3+I2mVlo1qzDfqzMkyOTrFkcsn8iuc/TQgp96Uo+FPLJfR2qzfU/7FG
y/fYdLmMnpd4peUjELJjGVgJVgZPcihaTxcINkHOnd7SXt0pi+600Uvm49NPI05D
vM6bc27UQOLMhI5EPDunpxGjx484whSAtXrQMMnJ0RE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7168)
JlmhGC9jelkfaoO1GifDskaKpuBLx1MKWQ3wOkLLnAm/qtOqGvctx+8wKSf6O70x
oQi6V1LSBpaqwfI3cTPtcN4guH73FVaCyZuIU4TVC6nsOpv6J4lfGCLZMNOP57YF
bPJgxumR1qieRbldX0aECcIxo0kJfc9TJgLWUaY/DCioAJ7AYdZIAFoT5/y9P9Sh
eKtu+ZD69jC50/C8lowq4sByd+gUqtQHGnaFi2AQJVo/8yNcNfALLf/Ij+pJ2NQH
/RJ+qpAJFL0jZrGslIreF1sM3nD25wvH7N0MqSr9BojI+J5M65kDTNxgI+hQpVFm
wW1rkuMhANOYUuI+ZfV1fpYjbpqGcOJHgpbJjbLg2sEDj+1WQDyJL6G8pZrtB2oV
uy6/T+KppD/x6tedSGTzrTXj64tL1rkKJ+cLaDlQKK8LO1PLvONgjXjrz+BYpqX1
dqrmJL7zt/atkOsVOcDxCQzLT+a/bSpdqvFdmRg6s84Fis14KOC33YEX0eoLAkwY
egJnhqqwxiSuBvd30YNcjIk0VXA85sSdCdpqANsJzTn+XaR1mAQfTe2MjtCWEnr4
L41fZdEo23aVwps+9G5cyfvEQL5svmTef98qc4imKr21lQTY2rhgcGMPEmG0SNlh
3LBMccwpwFw1apfFhaMGK2HJ+77/HgDq+OjXXFDjup78XSQ7Hj52W9UJXuPc+h27
kWD9xRbUoBg2o31RnS5aY8aAA4yZHPt8p9H7I/A/P6VkcW1EKlrpiXyQ0isdwHtc
E3feSAOXhRI3innhYMcBLljt21QrgqkgeD+rKdGek5k26796HpY19Rv7I9m4RnoQ
b4oCUL5g6kKEa54ZLoh/Nu9kYf4rl02VrW0ek8dRtrBZGf0sBRcICY1i10hmwX7P
D+9b+dT4qHqdwQawobHeU3BosBgp000MruKltUO0mTjW+VOUkdN77fr+5swjG6XM
PlTNvq7VuU2qbIrwHkgcCdVR1qG5NQ99KY6AXIS+mr+O9OZf4JcKFZmYvjFE2yPd
PeM1eR20zyzzutXc259ezttPwXQcthu00omrZWagqtV8Sl9nisy7fvbjE+i+a4Jd
O5iB4ZnspkA9JLiCaVWu8Py10SpfJLe93yGGoMeUSwWe9GTWZ8LXEPLlNi+EM2TQ
v7E+nMiUQT1fsGb/YRcVkPA90M4xhU0Xfeo0GrQiJ3KbfBk5myenh5KahwEFQ+3j
L4TFOKsF/u/03pJgZixHnL1h/mevkxpMMBPGvUIgZ1zfQSXy/OjmzfuoTW/qbtrp
8WgctckR2ORDz29QLe5pPvqugBkqoDOq3zBCg3GM/YF9uc8BUEFEOd0DUIilZ5sZ
tIgxYLWq1em4YsN1uwbSAJ4Ma+WrxA0Znve44yGIIaNlKdHJOxE8OZFzoBEO6/VQ
qJjPrd1OfEmpWqfWoOxpfiNzJlPM2yNX69W/+YcY1p/Kssj5T52gSoy/I8OoZGgz
VIEbaQkFYljB9z88X5emgJ9vhv5Kq9h5i1oH9qhuTFFj50CDHXsRq7vK/pwhnObj
iN619k75lW9vRQLog/zFb2lr8xU9AoAGsby1nV1xCe5mapSuyiI0bY04IoTaIy46
8G/pdlMksomKvm7PTGuSlt8suKxPxUAPBuYBKQRMJC7akIf3APihie5zj62VODBA
BcP6kQxM/3DFFeb7mChSOW1WHQ5UsU6qBfsrQaJyn9y2GGLY5wYQiGed3MgoUYzz
fyzb+9BvrwluGBBKw+XUUY5KaOat76N99t5kkIXXO+ZbRTDVwBpt2nt1NAmfAQlF
G8YFWUQnPW9eY1rNO9CMfl6wzilKab8n+QJ2sqSEWJwkQ/KH6XPv75CPk8Nk8LEM
qbwSb+h1Un2utsQUn0w5MNzf/bOdT8sDM2juAssGGT1BKOjCva7rFcIkF74/ZRYS
xUHJfQJtZLF3d3RIdp+8glU8mhgxKYrw6vY3ScB8CkIGEjqjL0O5Wj4OE8jyWaDC
A5E3jY6RP4n1snefanoZKpdMCQNJ8SxCAkEAuUX8wHcRxHOYFrX3DuNuXMhiLxD8
2VZGNysv+SkbC7z4QYBYpspoF4L64eWoWcKtulhU3QLccdpShX7LUvIJWJT3EFMn
QX1oDwE6X4C5zsuEnO0HkGYjXIQCkW9oxzadxWt0iQf6KxmU5sPxCg+vrYXVmwI8
+U2Y0Kj2xxmYsruTvLXAfP6R/FYvdIJQbh33W68wCoDfL/kLC2Bki6mZasb2AEyD
cJKE2yZrka432KeG3EJjJ11ZL0sVL/3aY/z4cmg+3ga2OcyZES+wFQpNGaLC8z1r
S4dDLkr+9YQQyN8vqZp6B5tWv1ThPOPI33P/asDasG1JIuQ+5kOIUx+1kfe6Bi8S
N/H5yMlVi54zQ8g5UUlrE7ixN9BAqqWOigikfS4d94gxu2fd6HAA327IIi+h24QR
JXIklmLOMPCgxajd3geJFiVpWm0D1SdDngLfn88FgIcoyauD+7qNMhKcQKv+PZ/H
EPN+5U8+BXEdeP5rJCQj4ynNAIq4/1+0GfdmVKaDRgczf2XvadlPA0izTX7G53Gv
N9CBaDAb/wwR5Y5sWkTAMQ0agydiJNeq7fJpSWHAUfLOFowGmebmdfrekIVWQIjx
WWjZGh2qjNQ0wMorjOLkgQQ+AVXyd9v4uAIOl1Uqkq0pzRtzaXcNLQ78/+EJX48t
CMlFqGnhFT6rSGlAus+1kjvG8sE+PwmjjxUTTkTu2de7EVqkN54vluLy4XVTCP12
nG/eWvd13NWiGcX145SdzEjDg423TWIcubrv+Er5FzEVsd+Ghe56ZxORkCbiQ+Kl
8oHiwIiMkf1G69WY1E7n8EIbeMtBKORAaqm6hQfN1oL1DOmJGYEmVMTZnCS8NMYa
uXL1dpB4Ty4L5mjl2adNsWx+mqUtu4WkweY+4/JuSFJpgJRY/4fnO8/5Zi9CbNZv
NvuewScIk0fYqnM9u6unPxHhl2vJ881Ha3Rd0/C8WxbfHenF3tcU3hDozdy39csF
M3IBXff7Uq5M6A8b1QaD5TX8jw2kKC3O+QjyxwUvF/i5Me7w7sxWzg9dN9cVN3VB
b0JYOyhV3NMhkrPFKH4kmq19SEGV/du1LVGTxfyeyYSP6wTIZad1iq3NMdQoiy+d
H7vr2da06UHfK8vGFf7peIG+y0PlURX3HeADOMtY73v8x9bi147nWzfd1ye3B61k
73iOpD9AgOzRchhxfTgg1bo5+42BuQ9OROmtdxMtLdfxlASSQrllX3bcbb6EovJE
W1t4qBuBnmirnxvD/caRQ0ZVPIz0/9eZ/QmMvQODdTuptpkijID3JBkFexMIe6/x
C39c/ktVZGzoMUi1Xy2UrPMEu2zeTip7atdxdDJwfbvnwHPWQGoLWP9NykVnk9FE
KekbHpW72SCsJIeIc4omUeoZYpMzHZfGZILq52PwJkbqBH+RKAAHsKTsVIQ4Rc/w
d1sRQNRfs8D6KdMcOonIqXmdFvdNM63vgrqdNg0PYafIX0ooXiy5I0PuUKe1kwXC
eyGWuaKy8OQ1jBadPzRryPzS3uwDBodRRiZFoJ5qujiVIlpVo2SJRe6u5K/U6M6b
67Tm/g+bZegu3l/IRTjfBdDCftMdyChkSDd7fdsfMXHfYRDbniJugB4CCK2CjByR
AiY2NbaxiReFMmslIwcGRZXuAsrKDybLVipV50vxm/xbdF8GW5lkoPGRjBTFRcNA
F0LURAk4qxcdTKRi6gZER0ETlq9OIAMZ1f4Ucg/4WrtY2SjK9oJgJWaSbNeH7jJX
hpj/oRe+DlDm86YtpmjSmqUCf9+FpJjez6j7/OA7CZYhwvwgMGP5cs/n+jcdOSNN
1l8yNnB+TYpi6Xvx180yyJL2C9YKEXLTyKh3X5sSsu9oItPHcZZpc2J1vmANeCgT
HadGJr7ZxwA2xmYXKoJrxnGl18SYROYL4DEE6JlSelUbpIMxwGAvPmhI3k0AcLxM
Fsy/69aHMLmOBNJz72X9a/2r/giksqss89N1JrAnOp6hFdGWEaJnVVSXJbh4RvCS
8Crxdhjl7jKFhLSnJRR+9Sb4xOJeXFsG8NE237lQnaNZkya8POBDhY3uodX2gziQ
pn3NJRHwMeUQ0BALm3ZY6Ux1Gk+Y6Xtu1ei6Ry85zFhWfibzvOoNP0SikW3k6jmE
rPmyDgcw+pHFRztDGDEiZ611UbgjiKhkjOSsH1hvF6IcgHBGX1KiF0anjeuBWExU
SZW/y/f36NMO7M/3BqifB8FyOk2XhUPkOpG/FOiAEiG43ypGgiCMaDaL3jQyGQOJ
LVLvrsHEc8WEt2Oxd0q5fRR9eY+mDje3PIPMS0tstTwKR8X3RjrrLAEu7wLSfqSx
ASezxM888DKXwRzMGyVoRYXIayw5kAOgr/eBdTjFLh7et21poNA7vLN7+pZfcNg8
rxYICBQWQgOpSJ8xvjIOLhz20hcX3Ba3uXrUoswZKDIHFi2t+BEYdElfkDXjYLdU
Und8FrxzXcJXrmeS804GQpgI9dZ2oHQQ9MOIw05ZVnUQDkXLqnCHPoWLfv9E0rgp
i3c4oNjqHoXQKlQOYtKQdVT9ODpEebXkRDFs9WBascyUJATRGqEYsWXS440ET7UQ
7eWr9Fk4yjn4nAGg1GzLMCjP2UR2ohBZ+K9aNkSoHaCtL9T1j0wwsZWaUD6z/h+4
Ypq+ZPCMmwvq7qwwJyz5ITwuPyPqsHBD341KNTBjmKvZq4ZdbrdzYtwvLzo9OZLZ
Enq5u/nvyZA+XP8yNBjEBLVWNIsfHnYNKp7+MO6KRoEkZdeU8R8TfPl/Eskf90ji
wQ5+4jp4z/ya0P0TsfZoPa5535dOkXT+jnV1KJx+eMJ4s62zGTvdFCWXUhOw4PnV
k+IQB7BCkFYYE2hlm2XMcA3GGzTbn+Rn73U7qMt4MKF1x6+bzejNp32evtUMKObX
QSWMHsrrdtd4h5YoWiJCJu609a15l/A/HogzFsQlra6eF6yETrQ8FrQWkizdLQ6b
6NxUCqrY7lyFPR1yge/8HfHC6DbNjYPQQ0WLTTut2dhQ1xHH75NvR4n92kP5K4SP
NeQLqZr8nGifJefDk2rNiK6dCgeOxD1wNxjc70TdR36l+LWuMrlAT+lPHNKNQ5gR
rn7N2ylBT7xnOFls0Nv081NMarwhRRKG0iS2M8Ijk4lVULBlDzj9ezvkDIi2lVdF
UEAAUX4h3tXnsxssISSfNYGsAVHdFDEUiBxU7cggYIvXO3wQI4DCUGbFp39+V2pP
laguxlvMgguiFw48KJIfxd9Us5zXhCWtDuP2W8vGYlj1OzK4c382uzjomoOmi7OQ
kZ/YECdeMeMZ28IoplvAceJZf2zUvCmYH944RV8rikdAeQNv0hT5qIt0qP8EmitP
CtoZmvrMnMxmE+gqagBSxwnxLVLQpQukqUI7CfEKh4J5DweJjyctbL03mBGbNew5
1dzQt0b0DScvL3vkWsITnO6W1pJJMzvQmnmh5Io3/20Div1p8PrCyWHrFfKY8nrb
fIGDoFkU0YyJK757/DwecvtEnhz9+O6KD/5ki3nny3dm/kqp8gNJ/kOII8ms4XSI
HIMLpCMiQERUencPwxh5xpKg9CPz3g33fL9AU1NNFjcrNuh+K2J0rz9EoqOeroI0
Uy4LI50L2FtIM8pyUlXlO28h9mUSiwHLqeJWpW6ezJzuLIbbd8d7k+WKsMm71IE+
2b9z4ybzs65rYYip4qmttPb9psL/Ooa+2CxX87Gf69HRE83Y3F1YY+34VlH9Hw0q
SpdIxno+1ayCu7jzXYSbF11FBc+6IFouam+MzEHAkKKrt5BHVZWlEB6ayYkAWz+L
aqdo7+vZ24t+OY77ZcP8eaUK8nuhpqqhdDwd0IY4i9vQLU+shSUO3UiHk6AZAm+K
oAz9NHmBqk4Q3A6f9c0jYSs5eznCY6L7Q4v4PCaZjGuX8HNnhnRZkaTuc6vsCqKh
zL9XkNX8TVU7WV7Wvs/C20VPdXQ2L3XW5G743vzdxXQhqOAZByfvg/vUUQL/SzTh
cBsq49WTw/fDXZoLA2Ry7lg1BiJMBgPX/5hESqDJL3uLWiW26RzjnXo9P/0EaR+F
9ZEgMvjXjnr9eaw/tG/fh05G5t/B/J/wuP/3EErWhgwR/H3csNIyyec7UvcdZ5bI
Nwiw2BV+2RGDUZArkpfZMIZVHIX9F6k2I6MpB253DTTxPURTWdK7xwmlXnNhuENe
Tzf1qeB0z6oB8AFOn6YxhKT/yTbMMIEdjEe3o2SLdBqmdBQ3PAJHrwnxKVX91DFD
SljzHarhLMktRLCbNdMJW22PMbQEswhKRB9F0nogvTQmc7gviZEQObCJuSKo2Edr
EUFnME3yihLwR8FWNS7DBWfhP7BoJoMzes3EYQtkg8/epmZjww/xyWeGj5RkSU+S
OIPe/lj3nO3E/1PDqPy+dj3rSPFJC8QgRNEuBxGA5R2ZxBsf2S4wckZngfgc03HP
vQ6MJtLoo9pjzbsXwVDwcvqEEoehFySv3eh9GY+/btf6jBfFURM0xE7RtoGkY8Sb
xn8V2gECcybq09h+36JVD56YWgh9lZPJd9U2G/jjP7SrFjzI2m8Hp4W7ehD+xi8K
TUyvVFapAu1cHwtkPPEdeVxLT83q8w7bWgDGoJ0TntaknkdtFHpKQ+su3TdSWbaA
dUHMbaKixtQ/YJfM5JIf1n7beTQYhd+2krN1MP2xguVKuFG6y8EiMfmcqTwsOwuc
+O9OkeOde/j2iItAqKeSSo2y38kJytM1Mpv2VJKRYbR+k4i+G2P+0jWV9Y+VHfRa
E1lJeAbXu96Jd2DCBZLxGRvZjVJiEvhW18nFfO2Q/Pj9RwAy/YIHZUN31vsI2aMk
Bv/bbsaCM0DW3CZnu1MXLn4vqB8rmK/AHLpm4NPlf65NvBsXdL4mm2cnBnQMwsQx
O29CqS7bQS3GvdzdM5FTJBKWjrjyjvsoQg6W9y6xhc60+jWs74q30Ock+3sq0fRE
KmQzGLokgmjh1HZQG0GDx0rsDKCP9814jZkuHWz1OBM3G18PnVF7X9At36MeZGRc
SHuU1vlnSaoI0+XKsbrZ5zjW9S7z7xWJRkp0+K0Mr808Cob08T9KVSGZrJMDT6aJ
BtJAWdarN0MmaiPksLOH0JQl5Za94mfMUzX3zKjDu6T5fK6nWjy0xfMBWRGSRhhI
ehTzIAUFRqS8U3dGdIQhDferS76DXnM/4tfZz1sCD3N7RXK3jMY2cOEQA382AuDR
OQiD6daVZWtOjWERUGEPNnPl71ccvtEJNYBR0cQ7rT37ZrHNJvY7AEf8xPpRZOZB
cIXlpeqOJv9Dt8VBlQk7vqphehCDdS8WXgkfx/IBZ1Xhiuhg7gH5MWh6skecmRLf
fOgbyX9cuTyD99Q/e9VtFSnjPiTchlvZrm0FZUrshCF7SOp8M3DMsW8J9jkw3oJW
nlQbpvHOTjx18tZMOOG/LNX/TWVGBh4H4SROoc2I8NMPaF9fu8UyAvGWJ9G4aHX/
KyuBuKbfz+58CpmdFQ5ugspOALbAkCOPRU2SrlJ7qLkl/2YnIUs+BAQvoyhbo2Lv
S1qTRF96NeBJlMUmXWONUKjgdjrFM0dhHSQ2qtl41jubIpryJ4ssapj702x+ukBQ
uiA8DANGbk08mw+nwaG72VGnONeYdEjjtjy+RkE93pN0r8uZAbkQu7lXBPpOITID
pYLSSQGF8JUuQQgc/j1gsdIkjeDcGNr1Qn59A2/jVVs1hJ0OsWAGeUrQtNsUIJ/i
qqL5e8gnu17odmAdlbq+3jo6DXOcZPAb8cpQlMX8l1aVlKMyGvJpmjR3dqoPQE9+
eGZ77tGLq5aX1y7c64MsD0qHH5SLq4J8HBJvPIICnrvN4fQRcxy9cCBEVJBvgGqx
q9JppHzMErcjlniIyqPX6wnO8B4Aa06IiugKfpEhJcL8YyGLF2iwbxQJTFJciklI
Km9b3a2dTAMnNOHKnIeNtytGV3oEfLVWAXePN/tvQkDTov0l0LcRrFSceFMuDWEK
3oItVFAQ9h6Kf7xmh0JoEz/9nZo15XBWvOtqE/LC0NqMhwNsMFPzeKrXBV96Fj3Q
ksCf022uuowX5HGZ71p7TM9g75r3ghPA0HDHapZAQq1pa1h8TcM6N2a17y/x84BL
hd+m5cqB8owNf7EQV3LimNtyQf1qwhvc69rrmXi1MGNn3wx2SQ0jaPm1XsoqEcjG
ffuWm79O+eeK8eHnMPtsURt+xMGMxlp3RVwEeGW/+DbAnMK6PJ3WCazVj6qAeEeJ
mHs+Cxw6e4g17tUELHjoAQ1UPiV/QNsWy6UlM0u2UERG9nyq6Uf1rVZRJIDzZhwz
pws5j71u0Ne8b8mUzCr8MeXUHfWtlQb+bA0JF4H4fnMus1g5By9cW69lVKg8SwS9
goTM6YrCCaKfXHMBvhI5Cgf2b+SMuV7K6tpNaBUuV4THUKw1sPjXe+UQ1ju99SyP
VXR9w6/UVuTyZcuK87piXBVDkVXx1Hv7B6dwKDdvhmDPvvBa+/24l/xWe8oH3TEf
U8eX9p92czt2RtsGQTSRsA4TQWaBtDQi3y/XLjXgknBQYWxvXQsrds83/YKKDQYj
cJnDoYyErCsccknjRXf8n2xNrd7vc5/jVgRxF0u9cQMcYTE3lBqlniZt/34oP4I+
mZSdZOA71A0uj69bm/dgQrhlYTSB1Tyl2oNPY9hX5Enz4Fh0HVKNPJRJqChWNmHb
fj4G0neq1OpuxAhdxfOw4W0MnkcXD5rs277KxDhsV3Oy5Mju4K3tsQ8B1T3j+iGZ
UbvM9GbZcAEgUWPH5be4TKEYsse8allW6Ts1P3bdeAEWS7Mwxqw/dRZcxGl40BIH
IiXUNnEcgXNd3mYxsKqXJyZzG2gHFipVU52HADQzegGrtT3JJn7b3w/kTgoDMuNy
8kPmRnTYE1pGl4jk+uYhXCG0HM+NG+S3SJ6dG6m1msJHSF/NQLjBCTtfs7si3aQb
DijdB0LyeqcaoI1HoGW28xwD3u58QNSNeFSqgSg/9mr90GD1O9NOx0FdLAS6wdvH
b82o+ItY33KMZ8K14GS0sORHV4M2p24kgtKnrhd/dUleb6Ac5fp9l9gTH5j1c72h
groAU8Ofc5UJLoI7VSNhFpV8JmxZuAbOaayIbNSRCnPD6R+h9WStsGuYQVPk5aGp
IGolvnb4bIC5V55rUgVR9MPuNSkGeQVJu1VsWQdwXiSjS/odXnoJVPYqjMGpqOdL
8zOfJQs1bvXBWRus28HSTi0OBNCgObhKIcZuOo4JRAEioIhFQhrobzCWZDkHyZzq
whBQ/SFNUgLi1m/gGtRWpnTMt3T/iWiKdy3CmEruAWOtDtbY43I1+ylF3bEU9N5a
E8fimL89ADGcQGnaPL3hFkh1dhXjataeGePHuqAxSQya5Qagfwhrq8Buni65CKfj
gb0lmulYN0oiC2DkrTTW5qeFgmAoDZ6xmclE6UGBkiZ9HtOlcC3qxlLZKXbFByBa
ltzAr6vKFGK6KvXeXae9sr52DzinT0C06yA7t21sTOJDE5lwbSH53bF4qKJChzlg
dbz93ZR/PPxDm6ngD5s5Zw==
`pragma protect end_protected
