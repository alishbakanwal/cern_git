
module ax_data_issp (
	source,
	probe);	

	output	[202:0]	source;
	input	[200:0]	probe;
endmodule
