// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:34 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
R66zfOnaZwQlpScqk9Q4dvDTXYLZqlH1fOzDrlujf6kg/0Q92v5V0bLSmdqlUcHj
qvheUHN6n7wV3NZ9FKeEOGcKckkaF5Ccm3n74Gnnm6iH7fC+4hjZkrjfruD4L8Hq
fn6/ljHUOWrRfG9hEqFTcG4eMN0BS/U1ZgsEsnABVKE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9184)
qxJ6VzVH3HrdXUsS0eXl4mvdag0MwwbwvkOzUybXdTNpM2Sa1NqjFXOoDDy+zGsi
J0uvi+gnTKVKgF2bBUGvxVxKgOVVUB83pCozFZveimnFG+F2REY9X0bRNOyz+Ze2
TPuSFvbQ9Du/90oUdFIKzPLXg2x6lVpm/i/wwlktElR+fOopvV+tbi8SvVeZTS8k
bELdjkaYSLPZKc8XFeJZCqRHc/I00CRwWqE/fSJgWFfPzEvRIpUkAM9i1sNMmDOq
1BaoIV7QaWSycvA0LgJocAn7Y3r3mAAViSbQUmRIeZO1df8rhx9fsCm3trxEz453
vuMrzQhVnut2BGr3jENiBg/GGgkcvesBwgVS8XTmY6jYxUjTPF7gaxttlDYqehcu
/y0OgM4pNTO3Dq3i+KK8rZps2tBl481WPGRvcePG+hqOgDISWZyF48ghxYpSmD69
vuIjFW4mO2pnwzk9dEOWNS4XUPLKd0UIZbyoLpvk1BEPJq15q1YF+qjmUtlBCvSo
NYCtB5hWWYApLLCvGphHwQirdZ9GLgWiA93H4BagKolBnSIWNNQBZfGm+kd+wM71
ojrbQlYRKDkL9+sivKTkhWFVFxzPseIjL+OXN2d+AjzF0NkaMBH20F/w/tdPaouN
eWa7AmdKV1w2z5oQNqmlP3Dv0XRTtmfv4fIdysTwcUciMTlSKujfHEeOESCXe99Y
rFlsP8fhT7/B3SXNrTpZWMLliXlZ5c0LdzXHhrE6wwVGS8/c8bTlu2pBd8AGsaLd
Bz3Ybf4SAzl1mfAyBhLXY8JGTKIWB5X/FEsAtR/scXJ/ZL6AhYE1GyT55eDyYVtk
5/UWpBowUMWwy2+8T5084U/51C07rJQcAb9bjeByhb4u7xu2OiUZtO34oKe3eeUw
fX90mRlRx9V4UsJOqxILakz5Wqe90wsgNoSWSjlkX1lrY0t0U/JJFm4Wq2WVJuW/
UkicMmBVGXAgmCg1MVIwAX9S7PCKEkKWLNnrPwVeAqiOVVgvdUses9uliiBZIxkr
DmJ1uKnoscv4jMASy6Xdk5haEGEbJpg0PeI+tMAfnUOmERSWWBUhSrfWPRu4xSrc
o7ke6G1bcMamgQhKEOC40u1U6BHbk9kZEeSc2I5ontHGYt0a2Qe5ezU0lBDuWY9H
zAG0oNF2lNdz530J6EBDuAkk4lxQ0Yk1SBhKdLq7feyhLX2+mWJUS1KMak+x2xbP
PZt7aAFb60eAme2R7U9iU8BL72DpmsmWbYo92zeP8MVtJir93Anwjl+Fmdrk2a0I
EHnnQFYd7CpjrErFCETd30bN2AF9TpQHqxKjSXe6Me9gvN9TirR/Z8ThtQJFiTcg
k3eZs4zofoRp1jfmERwiFnMwcbfPrJjeNDphYhNF+TwAc3PB8zihtLLxdY3JWy++
8qKUrAmbhoZdNiQrlwhZa2u70YswfY4ERKP2rWSlgk6xhAHY5XiunqKsL6+aRro8
ZpKx2Z/yqhRgtA5S06us6feiZtzLAAXLcKy7yoI6C6s+pt8ywn8xlDeOpdHj1jMt
HEXbtPVDYy0VO7FlQe8fwmlVnM704afzt8jySz+afjgulVhqdsW6m1Cu+nPIrnwD
dwwjpg2jSQuDlai/2q4zyPtZh4QHSuX/iQ40om4zPhXDG3U+LJEgImqiDD0+PXd7
gyZFVTVZvSuPdlk1eLALZJlpbag2GMEQvT95yMeieMTLF3MRfA51OrsJuM8+PnF/
SRt1kPuUBdfS4Ft7ttxcpsgmzVPaHUXdJO7FI4TBq8rIczPxbRD6NhuD4qMkQx2M
F6/Qb/9m3rFRsmdUhwlWBQ4kzpFFXYK8y5yfD9YPk9Rcm7S1A/3OCVjLyezKgp+m
xg/ng/BIzROfGWSHYN3+qpvoTAQm2HrYS40H/o+Z62dDB2pLwo8rPUoaI7QuVarC
B5ZDkhEYOB5UGNWyxvT+u6Oor7sGBOxESS4fYayzhPNgMWgNv1NFYmYuKP9mWQ3x
p24BbwKXvnuXBnkkph+Vs5Tw3wy8tBZ5wb8I1ikjhcC3xg7v2DTnGusKkFVW7WE6
8YjmrFHm224tyX0LeRljPgvMzMIvct09rZX97+dC11cbko01XH2Ki494jDn1tncu
+lE0XbKRCznblb1msj/9wPBg/E/ezdi6AUYHg1KzgGWXJbC4rUchJz7Eo53BflEn
zDkNzlWh9iTvYbl62HkPJBAL0tNhoF9aRoabcD/vnihZ6lo1dB6rtIhWH1rcPC0T
eeR0aQ6Kc3gHhYJKoakvuG9bOohDIXydWCoYtjiJFJA1IAs4kXW+TXayL2dwxYzc
O/e/aEgUexzxQVwPeLvIDdWJJX6LGDyet13c6uP9n509Jjo45R0KpyOhJubqmaJf
7j8cWJ8IPCDIFbzAZb5ZC6r65NgqTySfTcAac5KYhublq0D7KmDUAecC1SphWEkO
gyK5x0M6jtG9FRP9+EEzvnlompDzTa45WQiNcvNvE1VjLvSEyh8Oa5P+XjiwOeE8
vV+AJFU7WEtfJODbJ8oQS6VYc6sl0Swew5Vw6uMChQBzhS2qRPAy18wh1atX1PCA
+ZCZBj2f4WqmQ6QrO+vb72h8jgZ7GpiosSBOZPf5Ckp0frSRE3EEVSwD3wUGBf5w
JQKf49n2RY7pR9xeBqNzs8/icz7DUYEC5GAwXvYSpDautn9I4uiZaKkkkWJ5/Qm1
lte+LSbN0lbLUuyYjhgZY78uckkVd9JqkKEt43qOeih0ICDKL3UX4w2H8lGZ7D4L
mIsovqW1gkHlDWkQUDadHWimi8C0dm+tC41B7ss+qOa8kRAfZjaRJG9shpqtkdtq
gdrSByn+tbAWPAXkDsIXpIistDkjHT2CDQwB6XVACnmTv07JnkmT7+N+RWrK0lBF
TTy59VRM58nqKIOgCQQBdJMat/a2RMG3IFBlbE/5VcaC37+5cbPocbKFvnnJXRaa
ecAkHqQ+dUooIzO71Ps3Q1pl3TedEn1DqS/IbqKUPpBw5nPpbWw6KD6UFgETKkdc
WiD/g0Ew8oC/2BhkdWZG9vN7uv10pd25Jvy6EjLjAteVDeVH63rsz2a9ObogHZzm
QmaVZnjpt+E3HAkm5+rptnWVZu3uRPmGnZmKAc/THqS6m13Kz2g1MOLuBqqB0l2H
ji9BCjOo22HqrY12ZmYMQVpYJ72G0G6PQRsVgQ2e9/SqVOGKyasjFbeND87NcqQq
2lOy3MB+vFEmRXyOgdX8RqVMqjKkGs/b7sTT5FRETiMtEIjnd//0QT0V/22L7GcF
GjpjhFbSObkCZKrmbUoqfgPEkSL5imqPoom7QFEngysZDyC/DIM9zAl1PxFrSSdY
pPCVWzsIM0NK1+EK5gnfTCKliHARp6UKhWSbdKSk+8ZcCIYgSCWB2KtfwqjRAgQ9
T02+y6NpOYKe26i8E3b5JRxIMgu9Srd/gZyUJVcdkUvldEhwI4zLQpkibFCA3SNa
MDgRmPkDfIwlnukaeXBPYdiutii+5URjqD/7qAQjdlzR93CGmBciKRQamchZE2Pq
PqmQfUz7uR9of/mOBqo3pQLRj2t1+3Kc5R+WKwHMc442czYd/F0QzYqlZ40OkD2B
NHUkf3xevbmgfVUnOBk+hPTjRDAbKkCOjmtP0qWpHpH2M5QhQayqTMzSknJ7vd/H
fr8FQmIdsAGJb1qszr2eD4EXiS0hctwFveUX+oMMUVkTzdJNQEfNWmxD7L/zMrSt
lDgVfVQJcDYJimX5JM53yTP7Lr7NsPHMlHHqsn7YNanZuwvYPmL/rUG45zH7z+J9
iLf3G9llWZl2OOUJFqbRUdRjq9lve8nehjkY4CV5Nu5RU5r341DxVVuZDkr19fjE
XPB/IT+5mXnaJG6IyBiVHs+BqPnhBv09+sEV0h0/xMH5bVJURGxXpfXetqWYnqnD
2d/pSgOAhg78lruZjMSI4F2nNqK2uEaO0xO5a87QUyuFAzN52MFcXNFnmND76NBM
b2U/SV76rWCxUmY69BRYnkD0Ha3k/Q7Bw+VGSJyBIQWzEZv12pzIxrAI71adLWyW
WKvX39x2ni9Gqji2sg6IW5KOCqysOpzJLIihXo0F/TlX2UCSPKXMbd99PO4SzP6B
nIuglk0HztyhL3k9wL1Vaqy6/xT9gSq7UbaNeHAT0EByS0a3hRD0QTCoFWJ6WXEc
aOoHJuplVB4h9Q/p3CTYRWnWUU5nmDd29JI7oLcyqQ2hbHk1sGVuH4rVF1n0cUtG
CoRWd/rp+ItqnieJPREMlWkzqo9mU01RCn0638WRShH9DqNtrR5Ug0nyP6kxGMp+
wUBkl7eFLD4Jx35001ls6aQnnVsfuH5QLDYtZAcKPDkrDSbfKlP7gfkmXaPHH6fW
IwDlmlymi5bDj519v2GWJM/jH9w4v5WKOjW4/YHWxx5G4l0dWSXy/DOYYmANjV9h
NX+OlGh+ehqELuDlMW7v3bLx1+Fx1mCSjMUyLnJirjnsXTxkQN9RBQUn/RE5GuDv
c8/7VopHsB6TsRFI4dBDYJ1Zba+tzJOKjm5lO0sm8ylsTSiukFG9dY4T2961Wdmk
DkLUITvYP2BGlUG8E8asHkMjvhv5XWJvDBxbQvXBpD73jMvMyDkJ0vNpeSP25gxk
CWjZ2VonvuoVbD/JVMoqQTuRFF73HyqeYNFHnECXqZ8zmmpz+OfAt/xshunGfEqA
NFL20cGBXT+kEvdAv82YUBhC5lZxWz4UDOF9jnxVRMA2A6WNiqrhjN7v4pBST2L8
fVXzXuFd9pAefAARLDJEgL0yqEzda65aamZ43cR0YTd4Abx5Zjgr4jO1MbiUH+tM
hUeTXQKUPOoeTRH5d/MYl/TPmnQ2hMtP13nMIMJbz4ESkoJzmKUAWMXkRvP2KEdN
8ktTCcYxoVb4y5nZL2t8PdAYHeccuE9WJbHp90RLPkGr70PWrSyHBBqKaX47s/3y
9as4HJN/HuAuH2er2q3XbGcPFtwdPQGWiDCHwJ3JmlHTDRI6lJS7xEn9WwlQ5+Xp
MfqY0+TKsRyJFcbDZcD05vJVSE3b7CupsoJJz2Bzh79BFxmJ6NJQ02ZtQS5oM8fW
K6sAiUTEmKlZLREPAAqIs+TUsEzPDzf99q+XnBjgOxT0sNF9/9LPDE/wFVenVOu9
rRq4fogekljpwbYX0NmT+VeZXhv/JawyKkCBngPaGY4Kg2O2gKdcr040+9snUVhG
Kcs3zE2JGmAvpzcdycSKkC0sVmpw0H5UIKcauOfiQu/2N7S4ei5w3w/1oT3Jo0sX
BkrXKq1l4JbMQopjm9VMuW+ZPug6yJLUsnm1TVLhIeZNzD3R2zrzbsAB5NgTHAwj
UPayUdFgs0uiqQe1Wd1LkiW3klCcxkXt+3MY4Cs0Eto+3QHMLXaicKyAxTAU51o0
ExkObmDp5E/hr6ooayoXFhlOIlkmVzNmMQC+kUbs25+msCI1sV5AkBAGRNL+I2/3
l3JxPt6RyKnp1TwNH3Uux1xzvbWQs/vLjSAwuiQlnKLPpqlCodY1shXV9ESM5hTz
e7peyFI2r5sckkr8Nu03jv2QBZTCe8EqQiOKXShL4pdCLCZNaV4c2ul1+oHkLQ77
oaC0PupoNgLQlzOmY0GeDJiOnMZX5PhVnFgb8hvP6YpVTH2FP0iTuP2D3brXNyzS
1xFG8M8dVeaB8pfZryO6YxMv/jfE2YKzmeFEg+SoF2imQAmxQ6wKlP1A+ilC/zF/
SPnLvkTRaOAR9pJMM+5NEVs4e5RYT4exMZzj4SdnHnLNoYB0WBo6cTbdDxuTTUiq
Mhs2ZIaZHQepGmVAnhY7gF92iIOGSjCKP6rcmoZ7T62MQNcrG8OF+46a9lRqPC9k
2+3jSxopcZO2PEqvurYv+awnnjx7kF1zr4Z1rKEfDmc0+zmrWQghI7XRdAbvFYDw
4OG4jsW4JD87ZxLeUuxlzdFfIqNbrbH1qbooo3gS2s/gpqgGW5oE6pl2lJVjUxvI
d4+ieZgaCoBF9qr99qMJKV2KKypeIUzjzT0o/Gw+n+o46s2Dry9dOhckE/oJGnSt
ECvVMPR1tESGqqnAGWa9fwYHjr0RgmbdGwFvq3vwPOjdsv1CZJ7t/lpd5YzItWz0
t+9a+5jgvpHqckqU8Qb5vrcIL7VN8gnPZFJ+qJVNAtLZbhniJyXpw2rm78btUKBt
mrLJEHA77z7hsKehQ9HSwaEr1FhEdAQ30a+M2Nkhv+gjIm9Y1DENdFOg4B4/zh8G
PrVWws5TwByiGwGqxgHgMBsDERsZFC2imxFywpCuFxJtU5JWSbSjp3zHxIXrHnfG
tzRoAboWpp97/91byDItPccaW6sCSxnmZO6HzvOyw2Z6we3jVH06Y/nnuOH8El/v
FOVIsNhP4HXk5NgmT86MYhcLNw0EvugEALksSILuUmB7e6PR3IFKjNGG1YY2x50R
hA/PgM7KrTGFc1DEvaqFobAYU+QKHmV078KfwCNHTIQrkHyPD4H6WV7BKEtYVSgq
yJARv2XceuUxANiMjAFw9EuXhDyL6B8D2QENr6MFwWPyF65i8CsTUxvBLiEMRPrt
ls8fqrHiqeK8GOJGNI+pJxCZL42v8pMxGepeX01sUz4EapP9ChIZcb+o0ab2JBZm
3vxNZtL2PZ1au1Qq5PPsHuiByeHUt9W6NkU7A5hEnDMOsUlanNmybjSOqhYK1L6Q
26MtBJsNXOhh1y4kGdduVBuaqHl6+xiANIBK+5rSgCAyGm/R0CCgD7LhktSwJyqA
YpRUGizM86qKy3mOWvk0pSD7zILq1Fm028gIjD1cbT3aHbzOkFbllLksMzBUaQ5D
YKRy5iSmSo7LW1gV0SAptp8x+X80yOharviDQHdqkK6qTISM3mD09qYH72kUQnvX
h2GXsa+7o6W+KQcv8idx+UQjP3P/b8VgwTIDwhBy+3uTUa0e/FSE/AWs/lMzfLBA
Da4wF5Sas3r2oWv14hNuEO7JIaZsqutU/nUpMubNKUsif0sqk1RYnZre4BJY0bRB
ZejXHRUmFquoCEGJeT4Q5FWGUgcHq2jMKl6zHct4u1+Qm5234qg0O16DKvrPlR84
zoVCv2RtPmE9iq8t54lYV8nXdmXcnZJRkDRY1XXgu5lRGP62zpBQvVshr0yK7h0B
LKCm+NfRYCD9x9BB4/+2SxH1V1jkx07vWYD2ySlMTsmaf72TV5Y6MAap/RmuMp3S
tElxnXwwWYfTgvu6wGnbHKEM7h8nxfxO6SW6kIGA3l4atMhB45+id6XS8/UYTaMU
swP3Yd+6FkGzmWtl6AejZurOvpc2+5teOiDC8YHIKgAXNy1q3OgO1cUGFZQkLYTF
EixFhstOxN4oj5t6tyYRL1IRVP/lWc1kzsBJOk1gE8lUQJnInAvZik+EmKh5tTYd
F+1CKX4j6vaHdFTqYkCm1UoUEgpu8jd98aFfwHBF/w2v8ZP/z2HEuiwMqo5j4tcl
eHMR896L8L1szxVl06VIHZS5ngDmaf8oaASxb1vtOzCOA0wfr1NeX9/qNu3B4p4v
9GnyQHhNva3pJRWfy0HM8CVBwL6EhJRcPLfmeSL//cZkqoY4stMR2fdNCZXpMDs8
SI68+1dEm3DoPbnqjtcOqL7LIz8Unb4ES59jwHgaY6+sPRwkg9vMBtSJpy/yAv3U
+iAGA7a6lAosUVAPVAwYT66YuzTS6h5HO2I6h3hTNacLf9xQI0EVjKGQ64TAxHka
4ceW8w4mQjvnd8iaz3DyClLI17B+6GQ/2NlNocwd5KBQbQAcLfjcWzkfyJ9jXsLt
wtpA4om9NQViAiUkPrbuIT8ZhjVz5TqbIl6hd/IKYet8oi9IOFk1OTxubFFLEyBC
vUsG8Xdqea5LkK39uxC1J4k+lRKWb9AMoFTYWuRSs9dijdD1gAa2VuwzvJBXx4gC
mYx+F+d1CJijrmjt8xY1waUUIkwu79KzAjSIUeH1VsinRbJx4D4IutP9cRXGSumy
HwVIA0Sq58cnpLONntF+vzhTe+xGiCSRfW5vpL4f0BkQ0nHlY2YzYkdrZio9MhvG
EoFkohvnYdTqSfY85isdjLac66o8Exsm1S7dqMkC3aufGGz4Q+f14FfO/3IcsBwE
ltEMwJhlvUq4XWL2HVLQTgMXMRZydsu260GoQg0mOvifIisS1fcOBVwT7hxoa6Tx
LyOHmXiEVxRKRjbCF4YgHj1NiP0Po1k+iPnQhHnMqhKnmGOmUKqGoGUozG84P4a+
oAS7LooNgfIauxTeceb2CkcFooAZGWGxk/h04hk2ojQGh2cksNq+cbzqQZ+Gz/l0
tKVINYIRozlkwaIui3yLH5tzl0aWRqrMQHUwQeqcVuremA1SZxLYCB5RAok26uCr
1GBGOUavJd0nm6NhuhYfV5Ntr8McZyKY/F/pUYO5n+dm4S0wxHuCdzvw7xDZlH8S
JCGtcg6CH2U61H89P+7Wfvs1FV34YeOzVDRmu/gQSZxK45i/ylHpHcu8kSBbsvb5
oSjURaxOz8Mzw4bW9f845+8NFyYreKmLAo5rlTzbmYdrb9fhdhiwRXhfWGdpHBZw
kyYZqHgCYyuFlny54aPYqe9jCdW0/ldeMjtHV5f9LB4wW9POckbHrwPOtkgNJi+a
dp/xsCI/nADjH5WB3ew7wqNkVl8XhBqNT0C4PidOsIQjETWSQvufLWf2DDIRVUIJ
OHHCC2WInBDC5JtIry3xaLuweIXBMB2hIS5AJ1bFRq2TyGpY3GIEL9g6/s9z7joT
rBP6MF+DJeXGUfoE8rWPmnfigmfi/1ZX6/LkIFI4gkEJJ2qtcMBVwcRcWkSPLY+O
2kvHcnEImlPTIVBF5zBh8g+nWv9rsD14vC2aacGxeeCaHernrTGcMDc5BpkFq81w
47uPpoMh0vyF6IEWGhZxyvSP1MEQ1JRw7cry97ReyNhNvmIoXHCAzDYqiq7VgsLa
R2JZ9Ca98J2v8IPePEC6KDaLd58Unwl3LmKgqVekgFFR3wgZFA4RU6K1sNKhau6/
72WIFxOp8+tEa97BRCWC5wa49ENrZVAsjsglqRWEbvK8luoUdTyRqZOYBknGUbyA
9VYDlWSrDJat6lFDGrrh/oRi2M8fUaTTvP+mXkSg+oxmgWedkVYBMiD81CrP5fbi
6oCVnUbZT5DwPl4PFn7Aof8CqzpYYxxm1LVKljo6v3wdZkpby4w5QsvV/IEii4oT
UMEbDYM9yjO3hlzAuDyXBvi7hRmZbcy/BMmTsUrSqXHGe1MRqduEXszqZ+L7wP/T
UAPFOAv5KbAz6DwML4j4tId9Hf3isChub9DLJeERnCbgTIiIVgPiq+c8qgT2koCh
EhGSYXY9gwwf8jEPUKqWiuQrc3P0FiAq9G46maW0+y+JlKCnE0pWcbmlBSqivSRg
OMg4slC0G2wePjVVX3pFNROyOhKVdPU2j3Yjieuxb+cev990VGsvCJmLshu0flyD
zMwF/XXIKIoIDDqG2YzDpNysPmYvXSglKQvzi0nxAZsPZFYrvu1y1xl1o3D2ZLBG
1bsGov7e98IkW+n50rPS+blua0aoUZSNyq7QNspYE1TEf5MDpm9sL3LeT6iVy08z
4qNOn9O71pLX7Mz9k/z6MCdYTbZUvLySyHm8PFqzT2jtH2KnLuE31cSFEkSwRkGS
hYCUISI5kGwwRXAdLwwf/Xuoa/dqQQnLG2PxjKHKdsZfWFF8ucAR091YVYil85BR
QJoOOua/cuZp6HB4QwZj/wtMuoNILCn1a3bwZ4no5igLwweX85UEtgV+5FJBbyhY
uvB46BbQ4yxaoXgQo4me14ZsoDBPHXVtuD8PcRngjEPqVso6zgPBWQw+3dOTXSIX
cyKhRTkSMQXN+zM0MsadVpVEogJyxvghQG1Gswxaexgy90UFVMPHaxxHmyojnhI/
bdQnHVmcwpC5V09KbNBYR2Kg3DUv1Xt+igw6EITVoiwT8im2NazRhLDdJNPDVYsi
4TFhvZH7UUt7hfJf2tHzta8sItH49crojGYaW1aoj+DfGuJprmW3ru+bX4NlyA9S
oWbYWpwaUKjL/syYnx97p0v/XG3y8OpkO3OEQMmMfyjSqVUzvsyDbenvnwsEutQo
bGYYR8o/blW6ovSA+03EDO6mhODN/3s0JQAwnDI99CDH+NVMZkURNaHf9Ytld+HT
ZiyqtI8Bw7LQXIU1W1Ry6ZBQA7ztq6RYc79CIiy7hbm45rAlyJ1ywmrJt2y8pHi8
+Buqbft99y8ZPCYcobhVf+TVSr0/AUVDJr3NMylAZvAbznPKiKY3rucWOInf8SLU
K3NSUse2JEPYX4dysnMP7PgIMy6pTZzTFa1BjPoLYU7+Wp+1o1AVfz6mJDexts+b
Rkon2wG6/Cqn2xKe5MbmxUWsP4zfYnkBFloQZdxN3B2PGHo3L2QnGiRlGKNR4C6A
3Xfg3i/cLOiXWGfFuM11eb9XYKJHqQngtM3SBrggv/15RgIHejnY2Zysqh5iBp5I
UR8rYxrLvG0jLR/YRMs5zOL8PfgpAOH7ytL4p7JAGSuSmCKUryYUw9dR0xEyLS6d
rtT+66fKEbL8qAdcbVTbjnHEPdruzp9iERPdS4MiVtnROFVJdac69wZoh1hEkEJq
FYzu3ZLfvohEkCibjHxWXAZ7u7KT1/Mvh0OMrCvq+7MF0Pubapamuh7ZVJtndwGy
Z66F69RkesbT7FXgO95VoZEUQq+ZWMFtZjYaGfHIRW2xPPk+k6tYM//HW7NOkTHG
1Ry/iUJKR/bamhfjfH9Ddy8tDpQ2Ijclfx1kk6uN2RVeg1Y276yant2/mblNe2Up
E8k3wfXcZ4EG/a6YAKFo8zLwXau2sjJJTVWa7cnmdykiXnlHqrUhE4zOo/VOCgY+
NgsIVuVuuMTmgP+RhI2jUo+IgENaiT757eNXvkdPpbMphSREoXqQfAnU2H4jx8Kn
5Rs6GkXBDG9wTnx5SBjMsGRsk2iHdOXu9hkC0oDsZ+XV1MkSYZmAPBQNzei+detq
GNOwHQXrDNf01sY/QT9TSkAGhF3ksE4pXi9bzvaK/Txqebks7G4SEzxQX3/CuyT1
ggBS7NjP/d52/EBdHNYHb2dBmVN0DXC18qhNUOaL1cLCrSevMK1ZQa+VYVTWnJqJ
42fBzAxuK2zKBGpSpQTPKCCTfVbgFDqTLQEkpS8BiULpqYebfVWMXJpiuLKtWNOu
29a0M1prvTMS5y0ae1I1cfj8ig0pXSh+0RETfql0tZeWizwFk+Q3gifQ1UVJ6q4L
O5l8GhZRkqyjCbRKft0Xz0AKmzyacn6nybHjZJf/990lUoURp85U7wRIgAoSMIk9
hAeCSm7OjoZYIOiTrB5JLD8fqJWWRAZlTk0yoUB5RZhE19qNHYSzLDlrNJdweHZO
EGoAuGvSFayJvcV+PBC6+V2fGpWFJI4c0n5Qes9o6xdtA+HnAC+ju6Jair3BJFIy
G9xEaKnoLD6quoC5E9yhfMMua5Ni2o/h4EtazOkn6SYJq5cW0TateGQhIu/waiq1
+l8Up1UNQOtXTBGu5LqTcQRUL27w6KRLwUFjfvqdsfKSWYio2uFPZLF8GlWkE4Yf
F4KKoOGGDpnvrNXO9NoZKkcq344qyLmdim6ud+hFGOTiQIcZdhBwRkhF51OpMZB5
Inuh4Lke2STzfVoLpKQQ+Upmi9DmAkdHNTL/e0fhi/FItY5h4AmRp/BhR5WDVXeK
uuw3zeP6RCZH9vMxKp7C47lpqffpoW6ECTYR+kOQBpBFbvJkOhueExcqisg+zIJy
m8V0Yi+TRP87uoGMFCi6w/T6cmFerqf0n7zCqnaRkKjc6MduD0RYiMwTVmTMN5Oc
2Ov19POAzXzxcZyueI3tP5QTGdPsrHFygOb/kL6f0qQ3b28t7kLMLEEO7MbkZAMB
TVHSquXA6pjXxsEwKUOPfbrXWeKRMlgOKzn2SCksqwZILOudj+OFhZJn13w1HFkF
qnSmJXt8X10A1rNeqSSj+aKz8kwkwl8Z4aFg67J0gpzRkiafyXt7DAPK5iakofJp
AQoeb4n2YXVb4NxOggsj9S4TTvJsR+A70vKAnuNyVupJB2gkWVz1XwTzji9niP5z
AlZRsMPpd/Oar6ckRkhkpNE3SbQFgpxh+vn6H0vXODNcK3sVsDQiJiKP9iLatQhr
mkosc5/15lpTv+SO1iYmQcHbuE2mG08halWGhWSTLRA/339673KT1ayuiNZkp5At
mZFDQnbEdoVycNgh8d3mRxAyzfWjFrfMvdEfG8w74FJMDtQlkupPQuo8JNJBid3u
wihKIRPL/OTX2ceZ/LL/fA==
`pragma protect end_protected
