// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:10 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gquJLdv+NiSjx4nmT6KF9AAaaWbv9FYlS2HYRcDDo6i9LYjzBpg7gG8Aos/TP6g0
MKRNUlLr+gqKcwNZspKlO/W6rTNA7cGsDSsPXVN6fHH6xdgIep4sspH/eK/MY6uf
DLBb/JULNUc2JVncDF2/h2hhZ2Qojq/Hslu/ni1IKfE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28032)
wdeYigecEEuYal6g8h6dFyBOtlvzMIu5mKCDiXLVzRamEeu1M3C+MuPvc9wRE2eT
CMM2a22prbqkquOakHp0OGvlfQ/HGgQ7OM0w/1Kp0n6+Uj9b5fjAE1/wVqJo2aQq
9pRtTIIAfwINdnU+rsAsd8+vJUDLkIXtnY11OKkY6iZsW7FfrtPb3mRouvBCc3kx
2EREhWnoQwlc7GcwJrx277b2PhwRuLw+w463OM8/sxAiBErCnDW3SSwSOaHLZNN6
ieMcGNtcGQMpi256sEfXV7vRJKfkc/iuL1XXudV1WaPb4siNb4J5VMomxbz9V2b+
eBUuOWk/6HG2gsUeieScAcpFudnt26UUo0gG9IK81cB50CHKW2UBkCwe0CYnjiy8
B4wMYzKh40UGZM7BGGlUTbf5WJjNslXugwipV35Bd167bMVOqzcpt+DGCRYNTygz
WeqqyXmpFhPb3VEuGcYwO65mC68GdXzakLHWjfGTHD1R2rMDudDcs1/EZxjUTpEu
KKht6IhjVNIDH3VrnRWUBYIy89i/0ZpHiJ1+R7JcA1Vnow9ujTc65o5swKR/JEiW
hzbzH6s055mIXSqfzmmTL7kLP3b4lPvPwqwYBQ20+cXU8DvtjEd9TRFgdTD5lndu
Ib0N8cjyAqtNjKCpr4g9L8dCuDzerLER6deko/CUCd9YSmO5n9qBH1cuIRSylHS+
5eBprpngNeKSNiIrMThr8fPqH5X2msBpvpBGM/4QNjidjEP8aYti3ulfegwaSxKP
ix+RNvaq9Vj7E4BADUjzMkc4G9aeCcfGN+c2IzuGu43yUcDg+VIbU7j1GAyVfMcD
496kYD4xfhoCgKzCpbwv8IRF0Voxxc+7JFG9arFxTNyBgrS6bWQHkJwSpy5GEOwz
c5lT+sEF0wW1QCkUOIIzFlzi9brxlQtLHcCRZhLKweZxoyCsuh2xOdLdxTNALgUV
kCxjmO32mlt/V5MryzwYkv4YcdN427tr5BUIcH17aNNl7kSKA9bRuqmriY0SUclF
+aXZgUVo09FY07gynOyU8FIlqOh6maw4lLPV5vcjns6Db1U5A7FG//lj1TFXIIFN
NHpB12vmPV+Kz1I8vaF04c6KuIT0s26thhhUfyE669pwgZwhH5r+Y2vJNkaTBIEA
7+9Hrf0zHMrv6hZ/gqaggJQHmbTVyAkpmY55ArdjuHfJMwguv1FodnsPuhiJ0Mu3
U9litAGjmxsQa0iFK7mY8hmuI+HhTIlBZcazK5MQkqVGuVJmrQMu83p3Od8sd9z0
o8rq4Irn3wP5N2qUGwdsPXddfnBcF9htyMIHB5MbdqGzd7jTFFlmwTQViIjkedhh
kjtjp51ixvQsAC2fNP5K9wiI60E0FBxVRXqrPRM0d/M7X6soHrn2GskT6UK//bqx
FGNcxDs2vyb9ryF5xJEyW2hop+OgGL9vNW2kAixrrdtA52Hw4Zk5gSFoCBKgga6i
zvGuEp+LS93j9g3Rw17916eszdIQnTTJrpfGITrZK9/L9lY0z/cCbr5D7WqbTl6m
t7rWiJ6WTTdN+YDJwDY9rS2ummbf8KS3d1/ZAkNLb5x2zPFmyWnqCFyoVnfN4l5U
W9ols6JaUf7srnuQouAvLkM172ODeFTrHjAwyMz9CLnOZ4pnsA3oBVeRDW2On5nR
fsLyQGQDxIYkaglir95yk//pQxKBo2x+mpEU+S37L226UOP00gImlQztyyI5dY9h
gd8xqzQ9E3WgLZSBy9AFKMJmYBiJz+1R5aWBQ5fNTNTtNureQACr+fjbMmuLj0vv
CkW+IE7dI8ilgYVGNLCL+P7SzNOsU1j840ORMoOB82nn/z9Fm+KDCX3iQ25sfx08
cCOQr59NFYYZETY3kXPPThexx5EhXJcazBv7EP38ew1JKPE5Xra/XbYL3pKALE1s
jP8aCfZUMxDDazU8rCl4crr8gk+A7Lr7xwAUmlsdtBbHIZyOxmu7twAik/4oexPc
zMwcZwjigO+zahLXGOSXodewdKBTdiggWVF33ILttUJoEFtWjKf5+6WGVlNxRHAa
/xN2E2ZplN9TwBGyV4EjNIkdVAHZxOY3fX7IMjhZi7/BmSir5d51m2F7/fpSIvDo
VsbsZj8bmle99J/xG0zDKdSRfA3ISAK0vJHzcyohY5xduvQbtp6F4ezTeLwNxKza
x9wUQgWYFkXMxxcX1pddba9cAcGBdgU+S7Y9AUcd7cxcbrsT++lYo5yh1RucE72L
OSYO1qfa7a+GQURxvWC1IVpi6ducQYo/Wq9x/Pub2ozxExJh7A//FfSe7tAc/UgQ
K2Fev4ngpvXqCpWy6HNRWj/0hEuRineGPn6jR6S79QRgKRu/GN9sAybWlWmnw1gf
6LNKrVAQscDn5ZKlskl5MFc7G4groNk2G9kZz0JrEEYosZBvW2bS6VFlujHnoo5r
5hS+PY8LfBywhIYAjXCsU6dOmwuplz0CDuQOaJLCwS/0d0vSXUP+lC0cRob3qiVw
U+Yt6Q0nO60fhbG4r8IWH4KdA/CWXxlQwOJ8S39SaOrHF+Ejr/2gkjJ4anxZufGz
HbNDNgycrmC8u3IYoSSrD30ovwcTB7oXpW3tOQctWeGQ1GC8mSVNpDNzZ4tsyGjt
lqdgedgFKW00EuJ6qqiOjLJkTYSKDWcEMZopq8A/Fe2JkCdmjPa7Ov0GJJGx90P2
5/TS9TM8g2focbzoEFLV0u0aDE3O08VLjW+iFDDyCuYZrYRALdM9+baJoKWd+oRu
REn34at+qNRyWE0OwfFLfCPpCKsYuQgy+xITt0h/XlRvB9GXvmkv01hAk+EQeaTG
qnufgHkNeyb9ERINRFJSPBxnTzA1ap0OFdPf4eALKR8K0Cw6eoilbBmExE5H9WcE
Wsxz99UbNxz7McHOUe/0eBIMrlcCJT2XZZp1wP4mL/ZPzitjQ2r325D5zonFBqBs
WsduQwFYPLxTobgtK2jdDxybUx6LfqqC4GgCqrr7cvuStnehtaDnOa/xj2LeO/X2
H8U/ncIkZ5EXetnPN+xXE2rtSVF6PQM3P9NbmAxJ4mnHQfCBVoJ+OzcWJvo+BtBZ
kB6qs9wnUGfRdwSlIGA5SCSvMnp5/1L4RpYVB83my6ndIfjTbhVeEW7BBDkXjIAm
y6U3yf+/loMkztIUknRNzWHrOZyOAdADwI/bQU+uF1JcItNE3DmAey+x8qoLqsmb
971oE5E2r9jazwc7dVsv5a0sGp5sl71RqiTljTSMcUXoSuDfdDJRaNtKxvjV/Q1l
2anMVdq74tz6cCYpBR5Upvk7I7GKi1fTcQqB4ek6drTZOwAwCWMuTTJA20EZvztr
YIshiQqDRWMdtXyqHS8x1QHIp8FdhhbAIH8GSCKvjoq/AZXuq3I1FcIigILcd3o8
sE+fKqDKb3y1ZPL31kPWgh7NoBVAEIiVYtLwjcU6pHyEFAN3XygthvqcktvEDkCv
Z2EbivNjDSa0fYWXcSDA9rTAryjlQouT9iS2tdKJr+Blu4ihO+CSHeK6YqQ1v1OD
jNlYJDzj5RCWL+AvSKGZpRjdqAZLLcC4aZ0W3WCCl1l7RPU6tkR9UbcuPZHWeCUb
HD/7aKsuUGEbQKK8rD288eP7QaNAKiCHGrM+DWTiOcVqdNLG27iQ1ujit8pMBESB
DxS3y3qhbjzvpgKbBcuhwFEPUXGOIxo8wdLAObdKEcz49gDMNZJQ9HoV16twEqFQ
2j9uyWf/toju6d4SNAelnfuisarVnWCFVRHLxn4yUItOS/zbp0BN9KdW3BFg7+gF
3EW56ofrjLgceSspJnqrXH9Y+L7d3Tlfslkxa5qOJRF3FWMd7+IDKG7gqus1cskq
1dC3GdsK7P7edIXJVxY04tfwAJJ/WPY48mvgyL0dSoQPaupD6ekrTm19naqgXsXp
CCj1kHqSod4TO0JVL/Y5zCywFkxPJTQ5iNAwZkT7qsx+qwsJTZhjFc4ScNMI9L4y
n1tY5kWaHNfatzzfSreQ4rLn/MZawfvWufGbwGrlG1k3bHR61BOmOTo18ac6XR8A
kF7ggC9r4Nnh5JKj/9A1HcSxMPZ5ZVr0k92nfwa5HbQ/qROVKEYci9W7tf9QqN69
Q19udPg8TUQTnera3zNgYRSZjqCHirFF7igEcqBwlslFsmhIPG7sM3lEQAWoJVZg
eQhN95lHuzVC9xZ4EXBGfUb0bk70LAUU12ty3pN8eYG2t0WmH0MmBam/CrBxacaP
ndQKPmYr0+9IkAu+vhekARbaDO5Nrt95Q+r5H31Ft2FQJOjPxd6GRAIZFrBGgWj8
xdMgqtI5Ln0tUGviXRgvpQz2DOaWA9ujbDz1q4+nr388D66v485Amn+yAVNoWXp1
PIaTKY8tce2TLaix2Uk9fr/+xg61gprGAl5Sp24dncGo+xebOeL/qjSgsqh8PcaH
UJd1fW4qHqENcJYS4/YuSYCqT2UdfCknhz2+4gUoHaxNNiswS2MtCnaKPFj/7cwC
nMLlOuQyn/TK8Jza5xHFaK3kWw7w5eGEEZWhiSQOv5gVmJHA0xZsVe74sRa57qIl
qi0MknFYk7j8qiqy6ufxIWFYA8NCX+dvEoDJJIsfqIj8Hf8I3wH5e8/5qBXlXii1
/ONnCWp1hlXpHuFlwD2wx5KZawf9Sf6SWDdz3UAg9S2JoipdkP023wt1cZmHSExo
QWcIk4EJD4XtppOP/huqLvFMaf+j6XWhaWqz07TDruh13kmXGvH2u2ggNYXQo7oU
YruwYYSK6TmPPXz81GQNbE5IC2Yf4B/tFuYtra6Tc5nvPtDWziScR4l3k2A9R/oL
k8odjXej+RlK42qusZxtTq67IgK00JmiBsoshjd3HXWJglCkbZb+aLCbuooujaL+
g8Pll1EtQKsxbKAjuHlovPsmY63S9DWMsXcUXr+uMOQJeHpqRg+8OP/eTHoXZfCJ
4Gvuw6pOfQ2KguSMC6P/mDt4WW5xlbnkFHnjWIdTXIH9bd285eUT5oHMm2rBtLjC
7OoHKiQQPJYOld1RRg34fshIvy+qvMGAmLsPRHeS/aV9mYAK4UDRyimt7Ydqkt13
3GEA35xp777CxatvHj0vsw9Z2cxceWkjchfiOA4HTdcHy86ZFFt5hjUqWddtgLnE
tce6Fq5yCXBBEPa/zShWVmiU7mtobHi3D9JIby4R7XAajRejWpCSQw0jrnzuOC3O
IOsi5EGww25gws5/imJLz3rHN1d88mUm9DXh4QvWu8Vj5wN7iI7wkP/vasifv1zj
q8XmKFx2Zwm8moR8J6sH/RJVDg10LgJ8rJCxKpouvB/2n+6cHuuOP4zZWb/dzXjT
IJnoCa6Qj36lYyYR+Jq6jhf31zJtFy49RalD+eex1BiRQc9KpKHDyfj59QppjD4y
wIsRyOjXGO9c2h78nh7y5XGfXc68GqZFL8o6uKciKEDKnPy02v1PJpCc/Ozq+KDD
7eC9/Ts+usd9Xyu0e6skJx0LbmFBvde9dDsNCtG/PvyiZNW7KNyxI6/Ih+J0ZwNe
tstWVqWfSocUyRwebLElBsEU80zsSUdvCgS+QNHX5xrcd5bR16AFHjfr0VmV0vc+
53ONd6xojV/LozE/5EGcvr6paM4H+KQScYN/7p4V6HFp/uWGBuwkzdxVBzF6Scw+
PM7fEdPFRPcgP11O4+TkYgWfgedTPyvwBxWK8SGnmWlkGysdMG/hR3lXf72nGwx/
ydnGx9BqA+uslh7JJcE6hacHZrK8TDkHaB+JkHFx3paAkWq/0kzEUmgwHCFLlEiB
Q88Tp9Z5NKwSwbP1B2EZvkAvQL65zUbSarEFvLP6/GBh/QkOgVpA31tFb3C1w9Di
51SU+WGQ+AwtLiNwiM+7Onf+VL8s7Cz+mve2BLMPvfZ4rr9NvOjwXI5MLcXsOAZU
HzH7YR1EFaidLWfEWj8MyoGkQvg6fGdzJebzLFRKdMe7/4dvEdFy5wHwOvTsDGuG
mqnB5g5+Oq+h2cu+tTQwxuLQt9Ao1Fm0RjeMetIGXi8Z5uR37nN/nstHbN3cZgYS
MFXeosFSYycDPzNmwdrAeguBLV7n8k502hY7Qg2JjqIHPkVvjfHfhp5Rk9OgVZoR
007f8Ch7ahHZyQErGpOjIBD9sqbA6TwriDrdLrp+zlKpYfR43YHhrDZ+9TCN3fQT
JQy9891r5+k2sF6IkSzaOxEg/ZnTqjemqlBr/R3nDNYColrQdTruO7ZQNAbCUAGx
gzXCINBXGqQ0Wqe+4+MfQuPavfEKnWcE90Z2ygSWaBL+yPouLriW8Azut+hUo1Iu
Ej+8P8x9XLC7eh3cM4ZrfPDc39cC25ttvoSOrr1tpP+Fao50RH2K6FiAR44FpTYE
w9Gw2ztcEqEkA//kL6ufMXZJQsTMY/CIEGjwNMWVoVYVHjbu0B7wUiEAoH9t385W
YyIXhJwh1ApCSCTgoUMhrOULanVq5W6MVkKOCbvUbDrhwI+gZMVdGPNE7QsARAc2
UmOjjLBH9xzEZWCUIdGZ+YXNFopHvowdG804ILGPArRAf5Jsm9c4pSprAYq0uFIo
DWTJImk3Q/SRGOo9YRvpvxP6zqcW2BFpPIUcBs9SvzTxlzBNZ1K4Eo0gqxjP6MET
UpT054+yp1wMqQgEkPkp3G8NB+xMqobSB0/wpQN9JZg1SkQ4cCsjjudhb9GPmjfa
r1jrAlvApSCNgGHIwLE1Zj7LZp2xP62+pKLYn2eHvW3pAt0sn6IW5jcxQHAUqixU
iRwV/+MJ5ZHjeSuEtHWmlyeBS7mEzgfMvPqGCM5+7s9bUGc9oxO22RV+Mc5oBqYQ
fHZ30O7/J5eXIBJWWUUK3rBYWqHJN/hlSkhFwmDGozlcOVe1xdjMFAg7krID4X+/
bbM8eSpux5phzMafspbDWZvCBFNkBGXwRu8oGyWm5mImb5uTVazZJbnwpt7oGVqY
1ECinTFHWY52glxHvXvdlCZFWfuOUdQbYqMIj8LtCi9lg64mqascjcpF53WFFlVN
9czkFKQcafO9oAJs3q+Ar7pPgMQr0SltNyOdETkYcA132W8qefgudMt1UYWcEv+v
yd9oGHS79x8NZuoaXp8W/Sbv34ggqt0Mfk2+R09Vm9Ur0a8xZfnsdJ0FBmkSKVBH
JesEt4o3RD3zGQqxT0KA3I7Pq7oe7T351+2Ch2zM33rzs+DA7EnUyIxdoB2QSRfa
6c7J/EApk4aAGY9Lb2+2IDd0H49nFoxjX5k38GXAEwPJFdCQFPk4qHfm72duo7lv
MDOYyYbVIARNCKSRmbTQ883c4XLc1YCbdnxciDU25et4vV2Ex9X14vG26A2HEKdx
7vACPz62rTfhBCA/TrPmdG4iuXmDeleA98AetiPPrLYqseCDnfFq1D9Cu/tyISni
z0uFquJx3JUoHP5rIyVfSRf9IB90WTFlmgziZUnmF6fZWK9VcFud13klp4aeFseJ
r1M0f5tzmaq8XSH/LdtwtkUKWPYJyJC2zqx/TH99rYQync8XnJDZu6/8TcAaCSQc
vHxWKtaH5CoePdnWf1+QKV+0Osr9O8xBCntphtytquPq687tJsN6GwQ0aEmrG2j3
V/c2zsz8oomFetbrP821euuGy+yL8ZlOoF84Gs7HqtFn3k1RWVMlRjhJd87w0GBJ
kmDUWTzUYPPNffcYWGrj/5bTq1tzuM34qI/UqjFJLq7oV0FtMh6ih/NnRBVRuZI6
cHnoRj3VvYWtEHAH88uZ1cF7vsrgsq2h2PO3PH7p8QHUMrB/qgykfI6tjJki05rG
4XgRboETFDYs21sY+EeZVkzLWjR/aiGRFyKusouBWKRzow2RQtTfFzjG8s4XTUg1
fAYePtTjZpex4mKbKLHXiXPIqZMo/0hhkTZvWDCO6vy0Du6gkGxof92HeFPewJ8S
dNSx19kz4oK2V/zpVSoq6XqtjsYZFWt7pFwBWPIf79Y2iCju23/UnT5ec0sS2y+P
/BTGjV7fGvIIlN4dfTsN2//heZly2FIhLLJyxc3dadLQ1cFd3zu3hR/r2wFwu8f5
RscG23iBEOC6M2IGVvc5EAbVgLBSryXr0nGTwfAB3KFfvuxpFAJwDj7/TvEtiHvY
hi4YGpHU15/xgSfGkG4OvsEFtR49b1m8KzgxPMgLQdVvn+YoCdJGfnD0tu7ZUpTC
D58PFmx84CbGtpQtBEsGO6aTrNNLzcLqYHHhyf/RL3zstaacoBDNCryoDz36Zo2y
PYmWJGWl8yiumRsJDgYmjTd/kviylNHfkBBfBVqbAZsDfCvkDIgFeHxgiMEGpdXo
W3RwBYAa4Ka4CiaG8URND4Y81yHUhOVR9ZebT7axkQ5oqTo7elnJwP1vIJB7maRX
1u+CgWQ1pxynDD5JmvKea0rVS+049VuU9oc3yjyC5hbW18nvbPsj8J7ENnKU45QV
km4NXzp+qZ0cJpW9ryEWWQXrDSUtqhs4OjPIhYe9MB6thFHdRqKV/QaqQmEeNB+Q
rvgErBz7bIAXthse9ubTk8MiekanqAoymP7S8y8qSMBv/HaYhq+HBWDsUVUdp+wq
/ZhlzaPTQp/pj4buWZkRTSH/XFe5+hOmtLvXitM70Y/HXvFXLyhcJyQd2mfyM41o
DCPmpDnw/47/cId1gwdrzhWwNZau50mN6/E1uubHiYbFqkGUgkrynY0BplGtt3Sf
JzhMUMK/LSiURCVFQbvKDV+dfmEgxHPIvwOK9OiOCeF8Z6FH3JXOTMNmI/a9uCYE
MRSoGgNTl6xI5wZfk6csBrpLcagzquHAGQvIA77CFMFpQcnJyBxKcNAWeaA5fpfj
p2GA87QFjDS5QEk3lJAK1N7WZOPUrFDdHjy8y4Pr6nMkOdlFHpWVSDBTOyZOAEdK
BR/ENoUPs3CLWKuSZF4LduLXxgcZdsuN0j2VABG3KiWz9Z0GPBdrl+Pkq/uF/SvN
UI5ZJeK5xfDtfS+XQOmNfbculHYzol8oT/ZNViM69wDakhXXzbQ/0l5OsZB7by1g
FO1MLZ1TPenBuAEbJsFxRB5umE5haxyrizvL0A7J+Meq4PxaZWjciELK4aSi9WvT
Zx74likmOuHUoS8Cs7rfobsCRTzpfme78pARjFovH71IVWM9hRdrK7Q/OOh55+0V
nrq7ToX93kA3r/754vToNsrMzjowROqNIjm85Gt9CzmFVz7G7Hjpxv/ZFFMjGSui
Yq4L1Ax3p1dRbjhtPbSN6AMgDIyHnufe+lEAmyupydQPed2DX42O/lTVTMPmHb8M
/oKX4Zv9bSym3HTBOf59b6EBDkUPhg29Udaz0QkAI2NXAYoz+PeMv5T3TO5pB5Dq
VurUyz5QaCBgUtmZB8KbQV6cvYTdUlS57SDRIDelCs7CgEULdXZOyH59bwrdB8jd
ibrx8ADtnaYF4Dwu787Ld2CxCj0MTOEvjYR9lIPTH8U3WKd1EOcDS0Ed+hFqVo1u
TegBXBnTxcRUYrdOR5MbAZbGq/G7Gqw47obckxQj629ZdrXDS998aEFJN6S/pC88
ON3j6ydX8U148yMocSqWFVZH3YH5KI0M07CNQ6q0oqPRp8T+hhgGP77OElHC11Er
Su/Xg+Cbj8kLUYDXuz/oUp2z3tENLyraqUgopgLTthN1JtCWgRsSXfRYQ2vPmovF
NHniDE1ijncYbYtSIjlxazlDv8e50H5aIMCNw0+gkJUtU1SnLE5D50v0rzYNhVdr
txqO8P7XOqjfTx0CtQae2ahcZkQpWZU9qf9Cj/7gTkhFc+zoHme689yLIsN2Qz0u
gN6fywtqxjE/OSArAAMS1RUnFjHwkblmygUOqsw63YS8njIUOllCcgtzb0cSAlMP
mSJhdxMst2JUUYtsnCEm7NL4vdFCKn/+svelfSklMgDmohiA8XBZWLsiLWQ7MyKW
t40hVN3gO/XY/ymvi1CnR91PMewza+SC0nBshhQGTtnZydJ6iSIMMLZ90KdPLrxE
JkPpD5dhmIJylaOV6eDmmRF0nUAxkInrrCj78mThHqlRxVrE9TpP0C4tOTO7XCHt
SQEk0tuL4855vjZjbWuxecbZl6n6hbclecDXpNpc6BlivjFXCRHlnCyHaBMqthPQ
KeCociuibQ3QF/VQtc+QIoLLkJn6/9q8uw22GYanufMiDkOOSgGKlD38GIOLxaf6
oeGzvmo+VVPSs1vScGBREchfIboSxVQsTSS/r7+FLoRsgDMBK3BcODk0egQ+ynDJ
8eP5+2wERlCMiIfA7SVGyMbf1Sc4iaTijL4X+V1N1ucNmqj9v2V0deaky/+Oecr3
Rc+lP6LBTenyF6ZKPNSbYbwrp62TkaOPYqycW11LSAwT86fLZyXufaTsPTCgjP1s
lrjUUTYOHr51FczBrmqfWQoA3fsymyfYrzzp3fauYeWfh6wdCiiwR7I8nVenLcG5
hSsu5vR1OHoJoZRRq0Dz3sM67KeuirbcGVXfog9iAFeDY3hxoWhWw0teN5MlKW01
/EVTLkA6LFLOVS+XrBsDQqv4giPXC6rrNy6UIJW2bGbsh7YwBNqg6gkhVULLbwF8
e7Kxx5BMzSm5waPjJdzsKYGilYD7w/cDR9l2xCqhD7FbHeGo2sAMZovBJmrJs5FV
zbi4GdfrKP5sW62dCDWk1qnSt5vs1UelWF+49LhMpHSnp6xgw553g1qjB+Fxln/R
hyA98Mtv4XW5nxelikR6ZrZtMq8QzqkekWmRC1qD9s7wxY7Q7G+ze9xPdLFwtuLP
85nP/iXyXrwXZkYQJNFgBPqoBcGwz8BzgSEOytz2f/9lvz1/CgXqTLbAajtpkBCB
tKjoUAhtpce61XsWzDnzdpPnIyvHjVc0M+gEACn2EpumEMz/zWxRL3s1Y4E5Jlio
cylZS4Ce8/NgNdU6+WL4nr1C04WWH27hLtaJUAhYnTXnK3KU2Wy7sd14ifV38Pck
lkao8BcqAPQ/1zxMtu8GjU/QZP7M5UIhUuaBI7/yJsoEbSMVs4ChlrdHrnDVFIrQ
TAJDBfydYqKvTgQptTA6l5U9NZ79ySUAQb0Vxn+PUf3B65a8A+yw0lJr1WoWLL6M
L8tBTsFXMuFc0MZCRB2IIyZMP6EBWNhZapF5XCSsP2tUsShOjnAgYfjlmFmIj3Nx
OdwZKWvxhWRXSE/ynzu/iOSaoiuqBTRaLzc2YsfldDAAZEMiFVsCQsLYs39nCCql
mx+F/IIVPjtGok2gxiWBxiPXTxiLr9nXl6R6ijGnjw47GaL8c9ivmvoovA3fRVpI
gS7T2fjUYBMa3wDSQdQ7EGeMURKjq3e/4JqABgyz5fFjVDsyiLAAApgtCUjB7ZK1
pac0KjTu/fYp8n7d3Fc3R2H76l3/TYu6KNu3KPOS3F5Jh6uwKceHzTdImAJFYul/
z/L2iiyk6vjdHSkMKCigKlWaZA11FvtbauauqM4CL/kX7fIq82VAaLJ8/trAg41c
UsqfJmLPYBP08dCBD3OUYApjY+LirRHO2EmUfxd6atDwx4ijCyllpRBcKDEAQzh3
EoNXlZb6ZYKBkcCqxdWMCHbu2NXtIknkYtMKIHgjSzk1iSA69/ifNkvz8+z/z0yN
amik4qP3QZrbNxeN19ts0ko7ViGXcnR4uLfi7QZg9BqNs6T8I2D9+IUEQVomqXnV
iZOeQoywc96seko5k7TWIlW8EG3PRDw1ZL2dNVWTQc7v+ovx9AxZkyNkD4hqglC7
FkWGb2uYwjtEHYSdlX7JtWziviQZ/hTaeFkQuAF7FNwlee8vDlv76ONdGcVSWsmm
G9c2oDvH83tlnzQtYurmvg8cMqN9jHfQUaxd7JGMiKUtPLedLMoHs2mJ3Dy5/zTd
1mxgYzMtC8zMqbrpMGv0ypYaWIpxPyvp5Cl+VWXCQusp8ukY4npLDsdgkT9woBnb
7ByNoYkqOllKjNI8yShzSZ8FR7DiapcOzoDx1VsL1ewbdmEE+tGIsx7pUamYgAoF
bGldIwpFSwXj/0rHIVFW/lJH0pb44vPgatqxZT2MCkIwdHFi1K/QnpxH/ecSEXh+
/pI98DQ+MxP3O0Onr2qWuxI/059syEHyXGcSM990+LOPg6/OXwfzMEfUc8x0F+ZN
plcHcIlnule0vWe97gGHEZuu9kqK/XZjo/AMkPtPIYxGrMZSVM9K2MiT1a8QeeiS
nDyVM65o8VLi0vHCjjcixQ2zgcDVS8mJyffp+NqipcjoDw7+8TJfQOGhsLlyx2c6
BvANiMgzwulNmQP1jSLmr741IVa2kEOLKYvjey7nJ0em9h8JjUQrvKTCflbcWq7U
0A6uQxKDuPSeBgGtDuff53HYqZLyNF73zb/D4DLAPA3mxt2HOQH6+PJb7fR8BclQ
c0N6RD25J9VXtWW6MTUHFJyWAM/CXjkGpj7yt1cP9nEO/XuBo1R4AzpRco6RpIx1
zQsmRq+gX3PDO2OkZSbFIYDfoGbf1iYB+fYOUszO6G7hhkaatfMAOAUtZyskCcZM
+wT/mqtD6CZ9SP5+by+MiXtxVTEkUIn3kYrBjDakF22d8nYCY927zs9mVUHYvUCH
67QkrhEwhE2ucwLWvEVmm6ClycUEHWky//WxuhZbvtFOhpNGS0p8y+ODJBvbsM48
nUc8nfeQqoermbqezhqXxT6mStGA2SS0zS2cKGn5bRxHRqaPVuHjNJVIYn9Rlu6U
ldJ4BRi2CsX333GLetqIv57MOTrDxTui4asCPSWE7yzuiXdujY47bT4aOpTgr/2B
7JbsxXMla25K2a8Sa0nHc3eeaUlMB975agvFadagTd4VZDM5epm68KjCOHHfDljz
5JlBg95awCqC48DJDOMUZG7TeNNj+TiL0mdmzQSfL/5OuJuhYeXjhVkF6s1Hk9fN
GJq7CWQmw46Jfuscuvf7EaRbQJpAr7dWlwQVQJimBCBqIV74d3EOURnymSeYyz6l
wLatL7ROpzAKQdy+deeVPJ8M9u07cGLGTPDnsRKjE1izZdHx82BZPlQyg17tCDCx
jmzUNRkTcV+hz+7kTS/LqdbM/ROETZWyjQ+pqUWOCaJBIQEFKPdECESSck39ogP/
hdo5/Gor/X9Tn6t721k9D97MoqEmTSX+c+8rq8/J2YZ95gKceJqmNXn0sE4TrYHH
B48DhtMoyN87PDxFwwt7I0bxl3qkpbF3ppWy+ly8U+UpoBXBbhWYoKXHAuRpXMPA
sbTxOHS8ZjPCd/ail1G8Z6rf31ysjPeWvXsF6ijcvIaaHwWDzuhpBbGO6CUApdPu
C5AEZSRkmkqpinkRjZYnIWjkBF02KPfOVeiyCrUL4UCP9KecHKFRwjTSAuU3Hk1J
Orw4LKZQLgTAQPDJWlaSfynaZXWVfAf8HEjNwe93Eb12VN5LL/B7Ba7ueDKdB5Ym
skdQkCv8OpzefY97Tdn+2RdxbGfuw2TjDMKBcgm96n2CU/QDvJGOQYiglPYw4vrG
VAb7O/9sUzy6XQgZOaZ0N5OEDDzUcdpcd1Q/Mo+/p3vYFSrIQYVSTunNEOViym1P
bzxq+r6u7APEHZUiSnOgucZaM1BYJRDtfci4v4Mf68jBiYPGT48A554tzo522wha
LO+8nhxHtWEBojnFro96OxBbOEXS0UzRdV0/ygKwEbcCD7zuK4A+WXt3e2F3dWlg
3MraXYk8GVlcfemV8Mclrt1WXH00e5JQ2FbK+GChQtU/k/TsTNuTtQAx0t2mX+4r
mJH6ZSBYzxmkE0J4FNZ3zhKeg1NJoFvu5rEC7PSU7w5oOBAV8TQ5TmZkS0cTfHd3
iFmkd2jdLjT1qfr2/jLjvowa/ATdjbdA+oDn/6WBHz80mbqW8th8My0a8EZE5gaW
CfrEq60jhIXo9+gyGZI/PEuwM1u4mkreI7qOZ/f9LWFNnTjJW1nSkBespiiNbvDX
1x/b0Oj4j5hQcB80vL3sTJ/4LqlxqGg48ke0gfExTJn87nbFG4yvU1TLKLSuB/Ur
3S3XUMn6MYHbG35OK+AY7alhUICVeCl464kSojsHu78Vcok5PjQzHafivT1sTXBR
biSEG89ACzQtGxxETLJuP1EHKqKwD9Pw7bahkoxzEZiB8kKTdbihKKr3MUvrsh8H
zGz/TLfrGkKnRYRadqUkNZNxE5y9vbqkS0Nm9T4oFi4avxmEZ9mgHe4Cmk2kfxAR
OenE1hZwWm1dvQ8llEO/x140DBiuSwSAU/VedIpNXW25sLK58uIF63sJv5gwK1V6
I5m1E3wTXhgqizIq041lNy9cWPca5ZLyCtiiWPIssCEfmx/bN3jq20aimPgYMGuw
upCHhgFzQmkRTtZG3SgJSJwkdgDYnwweQS594fa2kkG5rTgK/orJTFcxdeewhGgx
JSVXaj+Za1tH9SPyzIbvADd2O1bx0G1Kp6YNEpS2ok2FdMaWomxtX+JRzbo4G4xc
ojbgtOY2yFnEeVtOE8nK8R3orusaohImzt4v/Kvz0ymZIopFim9qW5m7zuvytlMB
x1Vs/i2a7k+8060czjOcsVi4tYN/akdh5mX3XruCQNCO5OZ3uRwIKn97RuRnsZty
Jot/5GMQjCQJGR2guk+gY+zf2mpg6yIPKHCwVdONPYD8wFSD0GXxyn0VxVcnvXp9
psXqVx9RAZ4q85nHRFyJtlMLvw5Dn/rcCgHgCDHDLe3X2pKjetYXLoXKyhjk8KO8
u64+fFeRKj5BJ17dvKAe7Gdi/WO7G+8BBZZnkg/fGFLXpW/mpfXWhJoo6YH7kEVj
GCDc+yLd7KxV0lP0kD2IWF1SG08+JdPP6NIZyv9iauHAbpyxTNqzwEDfwez7Hs+M
QvWht3xTtd7P0cqszin3bizRU+5YcyIEvhQnkw9Cr81yMj7P9NXdEjum9n9iBVuK
G8P5WHEa2K//7r6G/TDM4nFOfhpE6HR1E3+S3tpbc3a1SrRV2h1tNW71UZxD+yJj
tidMzyGMQsrf35m9jsN2YICyYmsd5sV4dabnvftdzRvOYroHC/bjrc+DWJFoJ+ad
0TtChsGKAHLVoGa1pR2fWQXbZIQi2+Ose8zB8hDcMKsenXgLWmCWEIuFsaVTv6X3
MrQpdW/8HLKe3cIxHCxEwng7/94hgGz9kZ2GBdAtHAXrqLvjS2u0klXH4Vtp+zYD
f7Iiqa/lp6B3tcv7/jQ6hFtqsUrmqKwwyT3mRkS+5Qg6ViF2VzwtN9md/yUPcpit
R7f68QMorFvJRhuVmYZgzs13h5esKuI/fHAOQWXbmgiZE38YMtC8Z1nBVoKTBMtg
3ud7dZjWRZlV4Gc1idqxG4K2ZjVU74Yt15HqcF/zurwX13r66yVImHnBFpO0Nmb8
yPBkcCu1qqT/a79kn4TLfNIjGsM34RiVknTYQ6bx7xg4Sxiep8okuV6VBYlq+eEw
Mz+ElGI9wzuag5OZS4Mb5RcyL8ydZXAPZQogVR0nKfkuZH0tr34WkYT2oZmXHTKF
/6PoxLr5nmsjilYiWtWHJVfGzAL56bs/QkbEMRbpMSDuiYOrWfq5uHaDtoN9TQl+
OvqaeLy4w66sTsEMBpQbZzMgv/Sp+1Re7BrNAaGQ+60Qy1kI5Na7fRPw6B7FO+BR
ZSvI6k3uKXEA5HKGv/J5oNBNfuUt8Kp8c/PigkZDyHFVpQPSkxkH+i+LG9MRLHp8
iUu+bi8Hx+4dI2HA0gxYc1b62yqAIyNt7CecXtBjF7j+cKLSuzXmfJLzDpmAq/sh
fuyE4dX9IKVnam5mYgAStLCkZM+eNhYzjQRE7TiOE+28LqXWzM/dEvzUbc5JTB9O
UWhgmH8KPR9YWtuZdGHhsGgb0+Mx38p7c8K3FZc5Zc4GEDq2srI9g7Q+DzyalGAD
xAmAQ7FAPDzY4+BHs64nZLTl3JvE1yDj4zZCylkmmeuDp7R9dOUH3S6zcfl2A4Eg
DLJ8JEmqU6teiqdrEXitCP8aE5Y7LTx+GKsQjCo7kvMFHul6vrs5Bc98354SO/XZ
pP8GlHtL73ZldWngq5YU7+wQpTrH8vbdW65P/200GMQD9jkGWbFIfO/mWBDNweNh
+/r924vZsEOpwMuxou2/tTUcqGultzxcpUb9ytcZ7wXKWe0E1++gNvQ9XjpetoJs
BJgbAhokAgpgMDqyV3T8c4j0/vg8MBPUDzF4Zm8vNfP9WpF8bX6Y3t4CMaQGEyxZ
ts+AK18F+f6RbomThhreYVLEf/ZMRJV+zJORO0V2qaHE6CsCps+kkh55iMAxHaia
myNsN7eXopo5nDfOvIrKn1slhRlMTCoXLmsRaKfYSdYWMHcHJOIXbQO8Kph//LRX
u+7CoYOqpo1VxQLyrvwrWXDANn4XOZSbCtN4P8/41+bLDM1RR+hkqrEhqk7vTskG
AXzvyo3+xdYM7DsK+oEEwVJkMZrXrlsGq7RqoyrONeOdAacyL56RZ/5YUNLaM1nl
ZaFglDDE2JJvKksJV3amY0t7JxzYXIpvSnIL0dhloLeTqJqBGBZLPP30F7QsSppI
zEQYusb+Tovj8FmMUJyvJTaCAUX+nGJcxcn8JAVA3Mw2fdsG83jrcHhuUt75kc1t
62dIaDjryKRis+We5xXtdeEeIvn9dtMhxf2ekvi0+0P6RcOv3fjHtZgmYPsLl8xi
/ZpPD2NZI3wZ+oUn54M8L2ZCe6Un0033Aq6BwsdlvpmENyN+SGNwVfDDz+KCflq0
XET2qBoK1BtSTeOix0UJXtq51i5ZoirvOoCiHgqs/b8CCVBOe5+pUmNf4fEonRTx
WXVYcU6J9KmNswa/QJqsqJZYcrrsiZO1E9kBYh8aSoR60AnwhFD/GhGry02gpjb+
h2EntIzYKjjvmJx7d3lDNuw6tHEwJ5EPQ4AvI/abvIbjT/jwO0ITD3kQm0iqCTpu
gkd3e/OTfGRXB8pgduu8DQWA/t5O5bUCeeZt29CVPpXq8M6PG5mT9vIS6bfLsgZi
laEzkQEsca6WKlSwSiSIbfeOg6BoFtpxNVTAABKs5RsBfVOLMwSVhBpe9IcczcKn
qN4x1tDE4N75BwBxHHhtN6LKApm8blWpYULudzuzAygAIohu2X8P6iWc1CbmQWBk
q7TBtSv6M4ZDZO7KbgIvNyoSzK9EeutrVlW15JeY5btUjz2RDaANE/5L8zc0wH26
KpsLrX68i3TWtU4u/M6bncKOaRQUUSdL8X80b+D4MPiFDWktSR8eu1Ui/L56LKiF
c/e+4c1h+GmOp3KYNcDDRUfJq22yVa4A76AYpHz5BuYrlrb+MLqCjb+g/MCklZhO
t3OIwfsqXODYnOVxWpkqMPndcOEw5svPUf2Yw9iHnQTdRla/CiUlI5ICm18tQlyl
Sb8FodOO/V43H7fxNAAnsPWqvrgNPp9nfQk2O+VHsMg7506tKgHRlOFWuKt8ac5g
JmbxEpF2pOVpzyrlW6o7ZHDRDWYCdpXELzGPuGoBg8phF3SzWw8Cqib10cM9kBtY
JyjaaNylLrz0ZvHvGeqiDZSoiw6EADGqMRU39H+WjjXYW694M2ikWhkMKZaw9yKI
VZPspSD3PWmMeqzSfLAarvAnzOZ8chXKRpaJxl+rPYAPAS972l8D1LslZ4IGPN1N
/Adx6mS1FQmW7hCXbh5fAa90O2w8PFtZeqQjgyu7wPK7L8Xe8UTVGphgy4iEOKaL
VXZ2li5Ek5n1GXMUJdW8oYvSkABbYgyDFSl1i+u6SADPnG+62BYRU/LemcxrcE2I
8PebxhUHFZVZ/nM5hCtykBlz40mJwixpGS2B2IX+Lqmq+7k1qO8YB1O48jz/qpnZ
qfs4Im3njuMKyYaOEhrsQ2B1NOlZq03LzvmaMzE8yVuLRJyy2Mlcz2GwpFIMY/8e
kYlHBCRMq1alosAQBjW/YfBzIbs9nEyj2LfYYjhNVpKYzKktxAQWx4saUUu7PoIc
hnIce5kUwV9wlspsa1vqVyCfrrf2lj5rEGbeamCZmR1GNCyJzyE8/+zCIwpKjPgz
m/FVElUtKQS6PwDqIYLI95ne6rN/TQ4Emmfs9PJdqT9t6bH0D0cj1mSyofsakoq4
udF6fgkBVbkfvKg7LMmzNHef+FbUibZpE3+QxzZoZQDUsB/HUv6fLKQRavmDmZiK
lNPkRnpkE31p0g1LbndsKXke6QlvKXM1WsBUpzy1LHIH4Ia3AnHBXGPwBjC0SLlQ
9tyknnOCI8CIe6/TrFH/emOqGxQYRW5/z+7duRtleLo+qfbw7LwtKuLipqkA4uA4
sP3rgAacS6vzRJBqvzTBh+vqBUhrn5Dn+HAogF2PQYDfHd8aTETVPg+0G/96grEU
mhhYAVqzMtdVzvEHAZBAly/brdGL/g+JLvhayt0pbkdaD3mwv9goUGd7+0CTzRVY
UDU6GHSvHN0hKCvquWTuH5yAZzlLOB2HIcYtb4pmIWlDTKz3KFcqAmZiQW6crmI6
ai7sH3DnQNXDSkwxa7PLrIBkNvt+Zxfbq0zRhpKiMMBxq5Pv0xktBLeuygutG4R7
Ve+LzNyX5/4h3rz902HH4Yb22qLXkiQg+1d3wr7oa15fjDP+IJCkuw6dgaprKN7/
2K1/bzOxk9vRtTDf7KEdia16wckQ+Nie0VjabTYcxrLsp/9gXIilNd741YyKg0qf
MLAc1K92RF3OokUMwxmQhUJwWvs8gEUiJvKSOduLp4g0X0eCXXWFcZXpTYCDUgn/
M5SRYCTNBiFceRixGanvh1DYO/YD+BsI3CqqOkjqPY9FR/xRkhj54a6WpehzwV2I
9csenJjw6jCTDakjFid3XpZBjmf2q5U/OD2RHjBUpL250vpA9hJJ1+Ys+Ti2lCRo
cWSDBHWU4+Gn4KyHDcNDiimQruqIeJQxE1SYDt7HdQ/1LTHZneTURMAymRPwjeuT
H3rlqo61TNvkGThi9iOIMwSXyaSdF5OBPiSMDLn3oOgn4gYtp6E2dRIzYO9nOzwC
VeLNQwK6kRs92XecaZMPLKoHPebs09UcQUGK4CpBmkhZR4zEZ1+CFDQd3rlEC6Mv
AqOgo2kGBb/yuppWfGYwbuMwrC0HUmiRxqqDoqmqImxb9qwnjqu8/Wsfbmz6RUg9
6y/v/L+gPt4RKCKlvvV+RpJY1j4/YoPZC4kuqEEkJX+dIlHGMKaTbSRb9rLZfNOZ
uw/TD1cJ8L0A3S3Q1PnP14XnWlQmCC2NQZQt65YPitJdg0ALiC8HjAwknFxk/OfE
w5VDE2tuNRl1I4MxnYPGVrSoUFULoGcE5wbkB5rgqJaXsvZHJqmYjbKYy0he3uhg
WCapAwersurcMNOKpOVij8xBWSZ4KebkPUWjkIG3SWLruwk9M+6ZQe0H8aG7jxmc
iay93e317ejEYs+MFLY0RlcIxsoUDv9rfcYmIkaKAIomCNpTNDGiut/rJfy8Wk5c
ULoj7fZvB0gbc2Ot2QytR4p7V30iJXFmlpfLRrpRZCNtgDsjCYmRAAEr/VwCLRNv
Y3W2/+jJrppgpREVQsi31HZCDPFRtPF2U+9UtJ1zolRWlD8T3dVQXBWWJ+1JK1Jm
0GbHWZ+UBaHm4OkCDRCUCT38C8Eli4xyE1Gv6hjbPpdVO9ZNgAHnd4QGRH69su7u
bNOzS2rq8eq1pNxVu644iFWijCLZaehzYj9AzbGQjP4eQzApT5F4YNCC3/sgUIHV
UzP14ttYAN7367S/rOEO4ZypvJfFr8Edry42nnnagC+WYT9AfWcJXxUzZLO1zfRf
4U9lz8F6dpv5p1O9QDiV0SkIR8GF8jjwOe68p636Q/FhYEd0ozTJYTd6unExb0Ri
sbh4RgauqEP3yQ/VJjW3Wnrr4zCSLH9mXsJSCMfoUE+uxxKwmspWR7zoLh3rCb+5
xtdtra2hLfDRJ2MTOvN+0HWyMoNJBbpKnyyGFWcl7UGFdxFerwWHwj9Bfbnf+pVB
+jSN2QRPA4xNG0tKtO+Ua7bF9MNV0AESHM57zt/go+b2RzDb3BqVM2AykQwPolox
cTSJ6Ezgjsf7B/oZwEzBQcZrfnOEPbW40qclEh14VOzuccaNESLkoLWosiGtqB5z
MIemF5POc0tUzRL44Qts4vkPjRTClAYqDYGV11y/YbgB6gaxqWYnzHpgkffU36yI
W91dE51XcULOeObPsjQHhr6/RuFcpN5sSNaZZ5qSqUnGxNbDvuXdC2Swbmaw7zWT
ag8N4alW6d61r60N5LC4mHnTjoZJqSApeNOFtbU8EVbUXJvzGXLXjAAsbGvD2Ynu
v8MvdEVPi+yYQPftfRpfZ0KIGkTeFtgAaDySDIDblFCeM9uA7/u7DHzz2hWb+iHG
irffm4PPpdbqbhHcZ0jaLP3Dz9Sya/GAzV5qtZG5/Hh4s45BN3nwHurOIYy+8rMZ
jA2Eawjr3kJ5f/h1JSsfCYPUoUEyxdZJGrfjESPfaGkuEph3y2X08u8hDB+6c4r1
mN6i+N0tKXi4sCBve9ypAd8CyjEFW09zT1HzzR8KI1AHf9Z5Mcr6AUIweLFhIdVc
QfrqtmvYt2kI4D8k/A3myEjCOojRHxrRlNPdPWY+TsH9jrmBgsQe/ksLc+7vheiR
el0kmTPBtwhOtqAudEzGVvDyR2D05yYT6iGEoD4/4Vr8Nd9Lj7RhxaaSjNoAeHPT
wigyz7u+BnnfLZqIarYo15W/xpQONL/TdVnREoc/h/vBieU/0Ru1JjgOZqMvOn4s
Y0M221erqyIbgTp+WQT5/mKoyhbAt2xP68J4Oo4ipLuG/pnB2JWmX4TurZ8cgMRy
Kj7zirkk0vfA9+s4Vbb8wFR4pCbC2zZy+PaJy9rDpRMuKapGaDWl0DO9tT1BveJ3
nrkm4HoxoIiooo5RIoLyM+3b75mfm/V9TnXeNFiNVVjecnii8MVWr5ipCea9cDY1
7iIYZN8ocRB5FDvqIKPUE83+Q0qNQ267irJH7H3RPMrfNmhDdPjDTA9stTkVbEbX
eTjZlDV8b0RLgdX7KeLw2PpqeHKeyDzTm+izuiQNxFES4+MjfDirPyrybNdAuKzZ
NL/1hEnzGqVE4Q8T7Qi9wSGaBv6n/SaRNT2ys8evI1f6V8Hp+TscWQtpXoNFSDuj
wEjLzUfU+NLZIEal4/diMCK2BcAISM/X0oJZc79QpD1Q33Zr7/goJndlKoPvx+dV
5jOSwEPbPXIRbbheRgd++H/PCEovm5JHOr1YF2NRod2/YT1OVp5yOWoAzIcPzisL
RwgI7qHnxHgPJ3noTj2wUus70IgFOH4Ui0SeZdjptPZOD8yL7T+Q5+hvzq5UV4te
wFBwRWafTqjHzxtTBgH3XAXjm/TIwVkS7hlGGXMGqDlJaG9CmhicSnoo3tSJd05F
am+VS1XcOVEz9DuBfnhSTUJItCQZ4X15NojNA1HoNLHl3prdTUJsEBZjm3bS79hE
QStj+HY1usjvdD/+jQS2FCYcAvPKBuizPHAVtdoXabKAfsWS0MbMFxxaSTnBrarX
oUZAwNMVtFB15Dh2gFiginYhXJL3oELllLmYPyC6oLRVAXWX/AXom7SGpWI2OIdE
J4tQDbD4y0nhNbR6QXpcz+edU4GBYoro6RJstJVhygnkpMN3/DjCNjSrgQQWedZP
3pDFdDPl7BYOlcElbi+DDqzQZG418MVDPJDARwRugRCDFV3gx9upKTfDwOblotyW
ykNgXMraE2D2EszBy4DP4MdskVgO9WS/DlAL7re8H5rs5GWSFf5pmEiyIo+tL57a
ZQLHodxLC5jc0W8UkJzZeuZAGkm2NzFcLXV4/TK1cpAKg5YckFYDCg/IkM/vcBlb
xPFEbCC7CN5KTRJTRSNj+CSY+lS4LxBQ9WcHI5sEsq0fGhKE6O+Ihv89pNI1pcVF
Q6GJ0Pew3RmwCfZo4cdcILxryUZED/JXt9yGsWPWYEd8zxj/ytvjUp1Lrt1wCbWI
15fZWUl8V9FCx0+Il9iDMlI934PqSdiL4UeaTIyvAwkJ3NtNSRqx/84t3Sa1BrFH
1mKGnfquR6SfVsNC+vht4WylAH+8P5G1P9YwfJD4TWodGetG5di/2ExxTGRaW/T4
KRqle4DdNyMmh9ghlmjl4NkL1hF2QX8AgymYANjnMq9pixChOlfXvx6qBeRIzBwb
k5IchmyTfulECY3C6HLNRuKjel+1qmWk29mhgF/+JPhRq+5Ws7KV+qmcak001BQK
/TafVMhfZ1BC+a40Nw3Q4/Eg51wA7C/DJ13Q8IQD/sBMna/sWKECQ4OdpEeIrR+H
vhciUig7zUINiK+Oi8z84M3nQdX2wat3MhmbJuWAhWKBgY2c4gsGtH5msVdgkHH2
SDWlwkNGNGfrq5sK4oapCojSG2NlzU5xcA3Cx0vC1SrgVB4PQ+UjBDzLnzxOyR3V
P8uqLbFEj3pkKScay5FvcaB0Juczx1fRaV67Ciz66UGdUdwGdh3y+spW8RABKzeu
TWUxtgS6eKv8LcuC+fzsc4tlHKwvA9YZIAtHJ4Z8KLH6s7fpfKgzNUTPxY2Mi4eT
d3KO0XqMmHauE5Twmk3CZti61b8eT6TKcYeEKNkWeBkJRBgax9rFaT1K7unBm+vX
G07ij5jRQLXAndNwC8UWnRfuJhOD+HX+GVTw0ELpg+d71KYtA6V2OkpCpFXjkeMo
0rA4LKrrRMqiT3eQGmUCgXHZsQ7bv/2ft39V5DX8CCPiI3sb4+GjOgUNdKSAdw0q
chCqSuccKJB0/CVyd1xdoMlczj8djE5oqUMS4BO6Zm3IPqJgMJm+bvZUSeHe20FM
oCuBGWvPbiKm3KbWBjuUmfLTzVcVxMPWCPVFQbJjQS1vv0sYt7ZSJHhZRIAYoeSx
zX6JwUQOT+CdgX/Q0efRL5Cmd64SCQfV9GO5gF6gCGorpyhP9Nu21NTSjHGPmSpU
FiOktuaaCCY/xhViUMJyYzhRj99x7xOdiAzgm3eq5ZbW80nKmyZOb9W9hTaO5a72
YS1/lY234a2mmGbnnhWZbi/IdcmaLEiiNKvvp5O3od61InIVO9vZAN9pW985/uTl
OEhMg7ixCfY1p44e5/JmGH+NNuUJ7anf6tKexCYCSqWYnpb8YCDKjgObIAhf08J1
SfOIaDleJvvu+JZVX+EyOyBSV5hhrIpS6dmby4GNp+rDYwD/y8tpXlohwYohpmFW
aEui2y+ay6BX1WUls4Pk17HXjHhZCzmosn0G6xcRIEhYN0J6VLM60GzENF1AhDue
XTbVoJD0A6nK/CcRsrPr+2AAmOa2xlINSYxHVZXkokzPUfLDW6PtCSPoLHPaeinD
YR8jUtDGlEElXmcK6QYVrHkqSAxqXFaGz8wGFcU5Y2RsqjdL5qeTUyjRNth4BT1U
RhASmR89gmCoik6ZuPMWCYeITaN6zqCxsevxC3i074lKIRYTSnuTBtlE4upJAE2s
NTOkBbD6G5prOJ3B+GCEhLiuX+GulQiALrC2iYXCMUhDbAPmToD4ijYw9JsVtm1c
BzzhJPvVSFftxkyzuWcxx1zQBAyk8FCdNw3KWNsGyEu+iTi7X6fyD6t2OmDbJkxz
0eOdn8VWOpfUkRspBa+hBYt5c1iy+cPgoS/wHfbkYVsuIDswTOo61d8nHNAUOuQ6
aLedlSsMROV3aakyE4n4uBDm5lU51nmq5j3PgtwKblcAs91YSv78TcZuRCF6rOGV
crwNUIL+nO3PmRrKB0MFw7FxT+rIet+le3UvNVFssoGcgvbceyFnSQNZVJGgDvmS
tNE0LTaYY+1ET5I1Cra9JOXB09+c4qdxkq0P+7j3qkWOlyFwMo+GJd/aL1R/QDgn
NRmlWkUQ1s5W3bzLCM5A0DkZpZpw7dGHz9FDpNxVVhI/6XhrvX+gCdFDffNrt4RA
5UUzaGzo6iRd+QcHACPOQhX00PRFaWWLWTP7SphcmDgFfZKAin9CW/XuS18J8vgx
v/TNFynqawZxAXh2BTwnRR0hAvZWEZKjSP8ECQptveJKMHooOmfWwyG5IFv5eXWP
xu8adLcJ93Hnf2aDSscIFGBfM5y4FHpKvV/erECuPBHLRwMuNT0Lq+yJhs9y2nPP
nHx4n6gzeShi15YLsFoHqaPu0JlRlr2BILFRYzRHaIK78ZDcwhdI/en4T1evRxKT
hDVOKIOHrFH+zLm7zyCpJhtdx5HT7AkvOCsIkaM+gCeFzBa9RxXGR4NmeNewC2zv
XNgsDUmh2m3hGWb/1OeUZLzGFFflNrG7vBKPsAOjHZUHNyp4fSRXyrVR95Qa/gHm
Vc+DzHGWuGwsbzZVOi0NhGxfS3UPvdevhREgC3ON6hMJ/h1v09HSAy/pylA3Ssn/
LhB/baGAc59Ce5i6q6Ju+yCtytgZdd5d7SHHmyhgBUBX7fntIRtTMy3KSEcmewqk
y9dpjdKK+GthW8LLjQ9Tx17qLS5DSHrEQ09rw38M7gXu54JtQtdY/aHPjmLcgwOM
aIK2NkfpUM7jV2Q1BwMHvD/08FNY6nWnc1rv/NE/qdXSEIeiC4eVnZWaYWIrBEK6
BFSXE2FdKyzCMHMAkvU28lZ1EGj+SYDJMN2FkQlqmIXFK1jXl2hC2q0xtB2oYNgo
Ep838pkW1ZqkYAqKBBOKd9kLNdzlJernVWLBEVJfWx+FP63RSyeFovyO6TlXUUWt
1BOYUCxz6juxSpjEiAVtjbBustqjUWkyiLMGe8Uud2aI5mc1dw9J2vhJK/r1QLRL
+NsC1jZvIaRVHFaLF7WT1vrFHu1Pz1z4CWr/m8DT/48QDKnfPqCiQIfR+jmeSwk5
gaJFIbcamwvfZ/Q5eaQ3SLkMhEHKzPt2bolJbTkdKBguN1qMe0IvBC91bwsmJfz+
SnYdxgWylYhS+f6Aj8KBN2bJW80rXPQozKQkJwospWhcg1SXELU4ks6nnb8rt/pJ
wF4A9cTBxa7YW11rTBiZYYhViorQyKP1RZYtUH9piNL8kmfNoEFHwwmPQvnmqufW
skPL5RBxcaauY7uYuI0hSWDcK0OIWWqNB3SfbbfRwjMtJ5PfBdFCfr9okhr8JdG0
4scWs1hkMJ/TBblC38H7smIZGkKGGaIUC9LQvGLC4MyNtSeHmO04r685ZhEfk/6d
9nbcvJ/bBUWcW+wJnW/NL/KspH0OPa2fBOJbMOJUg4j+v43Qv27xE7UV1IFC8b9W
qy0A7TY/HVg8E7oqs3/YgTQC1VmDvbYFY+jzYcM0VPlp3f2davApgll/hPB6M6Y0
FizX5705d0F5TeAPn2uQjPiY9zM/ckZ5eoXwTh9CqUAbU60m4X/7nYR4ozwu74do
LfXTbbM1YoIanzm8g8NUgnPZhDDGno7rBxhpgxRioDJcIVCdBGgvuZ3pubdhQRNf
mDf9bihN8oOJKKr3h8K5lsYWSp8Q3LcOjBk9aE9ADoGdOK1+dbHyGTbCQxAhsesY
MPfftVLRj9KsTYKXBH0Qq4RLSsVy2uWsO0XUyxJrBuyptzVm1NNfryR/blb0xX/q
hE5s2Qg/jTdBVN6cuQCdgs4cl6AA2tB7EDy1IBl0kidMRR1Jn40WDILAlMXZjASr
7d7fHbHOS4RZ8Oorn22kDC+uBA087mnz660aMqhsB3UxiVz1yXeBIJliyFdJFuLd
PoTKCkm8X/0Th+JyCK9snjXF/SDG8gB1EPodu5JB3lFEZFXJB+sSGp1wqIkTXChB
xHOBdcEKMTmmoLSWDsizeq4dgAJ7hOEpecb40/otkKJ3pb9Z8Op+8GlUbrSf4z/R
e7U9QzBnVUuiLI+JVAD+7tTwcn1NzfWKkqVMhT6fw9BCd2pguafmFZd6ZO93JuuJ
y5fLHIZmGqsRJzfjTF+BAd5ITBtXtq7JEFSDgA1wwY/4BTedR/dtFr4UKnMjsX9q
98zvtyyRI/Rs5/DXtAuyJkldCDNgyM3N1T/deGWSa8EjypY6tUTEw6bTNSiZST7P
evu7LSY1GtUBzu8OcbTfwbwCOeqc2pOGuSZPy2fCBTDl3lae+uwbU5Ms0kESZutj
8aeSnKTAOgguTJjfle+732zltPbJTBm00ZrbR3vAFTa61hnBggn0OgtwiFPD7izJ
jgzXBauzs09ZYS5kj4wIzuHVmFRYg8ug98IzLW2sqW5FBaWmtMJHb6BSKQEaTF8c
kEDmnUts5lH0Sq7BzzqjnrkNB0FKQdLiipwlOfLI2lrPG5Rk2TKL+5vq7lZZZs4i
0csHaW7jNOS9KkNuMwBgve2epGl4Q3no72RGTMfK82ZkcNT7cCmaTmlClousTMGW
meLw4ija3kG12ZhfGIhK6f0nELgO2AHysvJOxenz6Jf74hxquYjOPkVqcqCqqIZ1
pjlmRm8kvWLw/sxyX63roUrANex1KFVRB5pZIVNXTWB4/0fUC5Potr0mKa8hyKCL
m7dOO+Sqn3bvS+g6x0+YNkHOewz414X+Yod2gy3KpLXdc+jVW5D5NkFdM0ihVssU
WZ/80+iUl+ELMLNQerezxYQJcDq5QBxLxlbf1ejKDBr9k2g4GRaurdbWbvB7J6ig
mxPJ8W0NHaKMAQpHAgUjb1mjQy5bPjbQ+kida35HNH1EXKPen3PwSjqE39F6nHRB
TpsLhy23JJ95LepB7Nf4dDwrhbwMHXFXxsAbkRVdf5KvK6uQl7sqbjH+7kycoh0X
Le5pc7kS2nRL6ftTDpvVG3PvDJS6O8cAnEKrRoF4v9hNJDV5GgdZZIuIKS1fAjif
xvYg+9JN+F0/Q2bg14+r/doTOONrgkIBDpY2bKBbTucsuOjqEiRThtcv7m4Qw4D/
lCFWh0pdINPF+cPaT8UQd/En6rd0Ugs8WpgUnRaGeMcwkrhAhC68GoGMHwZarm8k
xbR3B8JyggMc2rUnN+tZPEjwHU97jf7HO7W/Fno8jsSDmYFyCYs2uwTYfTCyvgao
NjxyWzFymNJ1wqgVMWQCfKcBYGunQszmFVGaK6mBc9V1ghSrzhgCYHf2nqGLpXQ1
JzF7E2J/B3w1Ywv5SxE7roT0rbkgdBtCa47WtsU03/Z/dbNNE1dGaQQVSBV2m1je
ga51o6lEKAiLUbfNr3qgnsMUErxOHuRg9zUMig+7ioVCjrqqPCkz8Qm5GQpfJdDO
Sw5jE7IrtYYLZX+nwagMtmLSax3uLoutz2y+QJl2g0Z5MLrkkgYO59ma8q/8U9fN
cfhPYoI8zCcAlPZAKxTQAtl15wZIMjw8z9js6yp8pbLWBeJj22hqwEOz0AEoFPMa
jRzJILWs/09f2HeUKep4XgIFEDaud5tGf/RBdac+r8ZwZG1Zi2Xs738ed6/yMGaG
+uZgepoOdrECTMl5A2TrfaaV+HiWnBLT2WteF6jJQMF3xWbuZn8ocOTGTrv1xMbY
XUz0WgazrcbNLGgnHl211nJnct7f/0yELPVQAUha22V6ES+Vls22SvMX2J0GMnhs
XVE9dPgTuD8h2cDs7sptJntUdyYq/K+9Pq1DTCwFw6WUiq5TtvmNzU3JaigKzOl2
PiuEvzvCmhXzQbeBSOuwgK7k+dbbmgh24R72OysDirMRRA+bMkxwVdanVrPrExrB
FA++W0mtCtG9JPMpAPGYS+RQrtzIkSVu/1eHFyy72nplK4JRx/Qxp0tCbI1JYwAf
vWbCYkxy54wGmu1VYTiy4bOOisz5tqAH8D0peCBR+i1BkyDj1z51x/kmMYO1VadY
dG0ey4WZGeAnKK24CAw9IXvXfQGa4vC3oxJzG7onYKSkIbEPMUg8dW0HQZzMVDaB
fiJCari2RE4RsypsP2xnZ8TajFINRvDkjIUdKzTs5Zmo0UkkFIh6U7a+vuz5bN1s
rPU82Q8V/56R39tz/OdtexANjno15xO4JMV8ojWAuy4lQgXzXyp70gWa1/LS227o
uXhIB61OmVsoYmSaNl/o3mCVFVfnP2S0xFr+dLimNEfQ+rUsXI7fJuMXJpAH1qQO
KzA99mTAPOOf+o4xTZnqdo8GlO3/JeD/lH6KsST04NrSLbnbcs9xkD0E7Fvr+nTb
nDIc1yhrP7Mm9objo9N5ZiFP1RCOk8rffoLZYVH/pUuhgQaoJ33Tdn/o7R0OhVAR
ST4wKUk7GC6DpwoQGV25a98LFRDhX7X8qEuyuXC+825sZ+FGvgJuFp6gFIeE2M5/
iJPNzeaGscSWn6fE2cXBkMFMLc5kpqsOH3sr4NCwk7d5ZiznDvLtjMRXYzx+hweS
hhnsLUP79vZlVmk6jxSkIMJ4kB01VA+vOKIevyDIKHC8wbfm8fmO4JDISkM2js1y
8jF7rQfQL1KIdnRo2fUTyypU2NZ6N+Awg1hxTWhZzguMvROYaY5cw+LkUkf/IeeL
KAsY5KxSuHgIqsxnDJWwUdI/auR9jNT1V5Lmb12I4R9Mfz/TLyNhWYVilnhL+RPp
wmunX815b+mtSCdlky8IugD0b/1V9b8Qa/+tgS5q+MX/EZHdpdZO/ltvjI0JT9BO
zq9R12kOTG7o8DXnRloiEk6lkkipcjML+WerQT/e0R6X8xZtUg59q/fdBJ58ZTOc
TeVgb5+ImCYBYGABzdpdqccee0p4rilG/BrzWxt+P44Tyy12ZX0FX87+9jF4k8LM
NZ6SVxpVJLffqDLBXRn1tbM3h67PWVI6zItNMrceeUpwAa0tvj0n3BncG88HSr/7
ObjwtjW55BR349y5KdUJzzWZZnIaZvM+VIsoxa2kwVKAduZ/nDdNtRTu1M2cNwfE
JzkWJ9wSkEj1RZkaH2aojcHE3mjYyw+zK9EuDSKywZhwwSKv1hpEmXds2F4o+orZ
WHdklcLL4+FonjeLDXirzcBi0iikPQSE6M1/+ZFddwXpbqsNsSJfpBQorpu+6VL2
jPHxLPbFIQi6lszTMRfKQOhnBBes4ppvxPHJf6lf+iqYk1xSK1BWK/gJ6uO4CEVb
Yg0MLWov+ZnaL9nuPGaC4XT5zAqV8xG37wrWqtGbjna7hBr1eRJuAACyP46ieouD
T/u7s5NwYgjIxrtCT02zrBi3TIu167GrSoRyeFsO4AmW2crXhmrBQDMjDOULRgyz
ug58WPNj/7A9QnIjr8MtLn2ILdoHWNnCq0iQXEHRuAsvVv391e8EL9YyefStRplu
r7oEvZokOHnk36LfiHxpAgtmDC0jh7o3KLhr2wHCckIcChln1tg/3du8WZ1WWRDi
ORHPOv3Bo4HbdOl1L4VBRRudftuAZB7iGZ8yieU5wzuypJ2yptVfchFBTAU/5Oie
vtQ8+QzYWnUCTJ+s+PZMpPnJLXQ6/vFZLAheSFcBd0rbVhHQRgnlecpwwF+m8pjl
Bi//I5YhIJrw0sVa+OfxcHiym0HBaWPEiAZX9ILnZDwDHeeyVlUeTBviE5MUMHnZ
C2epkMwMMI6Q+eAJiDQy+X5tHGmxU17VDaDwiOdP0gBzOgzw+J0XhosMGxlEDp6S
Ux6ON2gKAPYxZEytqVWmAB2w6uIi6nYFutblLhrApQoJ3dkCSY2wF/TWjUMgkIwC
B96IUU7UzNG+Cuiqj2exRgYAHkpU4orDC0aDsYPX6QiNdzpLnIb6fHgn8hvsrQao
u40QMkRebiygqUOOWxeqUk90sIKVrhGSlnBHLUT+ClfmO6/nyGzG1IJWzU6l9TzW
lenZGx23yAJi2SZmQ1z2PcwX4wvGfeNQob0fs65c//kPRhwokAq1aQGmYJulpygf
msCNuK2iTbgEMHLfgMQIxsW3O6n8aDaKZYtHr6NM0vX2M8qOvj3anSYBuNu9Petu
zU7y7qEflDA24TnrJkSLIkZiUCgSSZf3tAIbjZyH0tgay0tJVq2gd2SjHvaEJqqM
sld5Ig67w80CV4WZMaCskQtCaI+M8q8eSlf/BmKjoBuB/ZZtIz4iNJ0khaxIdjZv
5ar54FDsnXUYirodaEBuQ9eXBrfVvl5uOd7H6TGw8OKYADvRLDy45wGkgM+lK0Ga
fCzcHxwBvykfvVOCG+ZYAYv7ddtonKnuuOxAzIAJ0W3aXo/THyOI0/g8nwVPNu2R
adjRyWM8bnYsNa9CQ0zmELIh7ija5SpRwKGJrXEp+38l4A97E0L9g0oQLCAj+1mo
4fjSUut8IfArzJj9kpATuTy67keImulVi4VqMitgEYUAEZ9qhf82qUp3VDCJ071Z
sSHzoEWYNnxqoh/FO8k4oDjYqU6KtvAl0tgRiph0/JKLAlwdCedlvaSNjFFZ93w5
R4gsZ2LZm2j3GeaoWjF2x0mUb1SWDCcXzr/TXP55ffQuXMdjo+uKNOdFqMq8ms91
Li/pH1PEEGIQMpBGH9NfXHasUaj7OhvnHKZTozp9tyduNt5E0GkEoXv7kyKAOYZi
U9vnLEPZAPJHmOTzws3D9b1sOrXFQVqeSo+oLS94A67z0wA+uugwg+OwJGXLMarh
2J6sAnfW7qDfhxCY1utjjLv3IErNu5OY/pJTyj9QSqbhExj7DzcOEld8c29OnL82
wLTUQWI9rBIXefTU5+vzKyUe6oabAtgBzT187im4zXTKA2ugljSrVMd2FdH9+SZj
0F5Iwzj9Ysik9OdZmWdTTfV5GREfnhAD1/un5Rsc3kElusIlWG+JLUlQJpjOzlY4
T/nNFoPs3zUzQ6B0JyBMa0jXVxVd51XkiGgmV7evmy9CVDzncR9JbqlPLYuv29S8
tubO3YXPMIGdP6CXGXAZu3mLTSH3LmV3fc+Wa2wCxNomgFUQ3x4xJjx8bp9gfupi
J+zjmeeBsHXxBC9mqg74K4w/eq7kXzPqe4z6KK+ev/WvhjLFl2VMuSf6C3ijfDy2
sD2047MLTfwZXPApYiqRkyKJVPIWBmVAJ97j0+TTLVgDbXoZMrL5Bc3Mm9M3nozV
5P8P1xPRySThReJ9aQDEmLzz3cdyqdqNDGqbAbqfBaIOEO6cJcN335C4bf6WZDrL
YKudvcmXVnm2PBKMgjAJDmzLURpK0Yoo6tKhgQ+E+S9rKpBCubiOs+2MVShksS/I
0eGeov8Ki+ZBMPtjTt/EDLopLGxnb3ZmdJJxAQdr/qJi7zEuJV7kdyg/dfsDws6A
IxUSNkpSwD+UqCuKg+EQ7I58w9aEKia1aFm5jtIO0+0bCAQTmVuvbqDSQratHpkf
k2t3rzXN46KtmGaH/5KmIbFSTc1n7Wfdp2H29QpLluezFI9VNoRVetQPKK9aVFN1
ZRXoFRHTgVGQonlWR2swgWIvZlpIKLsbVouJmpFzbrCIVQJAYn0j4xiujeVgTi1V
3M+CG670226B40sJfkgymeLiRTTa7huE7k0MshPaSR8jo+C1gyMQkzt6JIb5VB1n
L1mC0DIB5qDfPYT3c3xCM2Ubl3lTLV95nh+x1N5vW9xjRhkp28Eu+KLBopEQjwAz
ayeMQeaTThTvmyf4e9P9FAKVW41hDOFdKZRJkGtXFXQzv/xHTUg2xTlF0U7z4qcQ
J7mg2cpQ7BQgapBrfusuUbGoIxGaBcMqR6sVjuIlTTXwUrY1k2w7Y7b0Dk51kbw1
j+/wgndiTw8SJ60PtBvG1C5ShNz/o5HJhbfAHAOEmtIpgi2KzHO1Hlzfgm2t3I/Z
QE11F3CS9+1EwScd8hDWyxtDvL57iCk77D84a5pUun8+p0SENur/KFz5oYR44J2p
19z/5v5tssvhNxqvh5DBJWUFcfFmwX5I3l1Tasqfa8nsfB4BBp63Op1nLbnJYUhx
Z1cq3SCBwBwgpQWL5i2pLKQm2kXbuWpCYMEiDhtFxEH6fg/ECJY1/IIJ9iHvaIQJ
ENd8XFLM/S74F9MZ7v+YGumq70YdfcofQo9ngxyOn4pqZ3ZAnU6knCbFfY5b5edq
xxxrbLt0tsSrwsDqfeFgCKtalpUeJkW6XbSVJHywAJeL9bRnfuS10gFvCMjwSptu
s/jcHqgFLpJtchGyGGDS29I3+PUTXdIUj8FaMksvqOTaI0ONRM18v1HQjc4PJGNw
MCc9ovkZlVjFlm/8Mt6GkDddQcSkfTyqw5+6y1ZqFk7olHopz/HgBT/QvW7K2mSz
hWmY0Cu5GFEUka8TBHiEyUiviOJ2oH96YjNZtwduWpTDUncu7IeFt3PAb5VkAvZi
IoxVVCiabEOFhqcr4JnS7Z26ALcUkcAGCRcweziAeNUFR7SoIy9GFYjSmSe6qi6O
GjbV3PupTX7KPptRP/p5BjpWu8fSnOFId9QW1USAXtfPCzYQH24YW/P6Gv0svGcM
UXAIKu7G+hWfog9oBuvBOnCXNeEVlTul4G36ladeU7vj0TgUvBj3xmYlbx1eYdlU
Yrw00ySKRkglkjLt3fJdsJbDpUQ6IzzLLsduxHXpvHiwOvUbLWpelBkZu1yJ6E0e
9OoGlgOwjrFBGph+Rrqa3WPwhog2Y8HOE2r5mBoMsJmlVI0W22uEtqmKYFf/jkPC
lbBFLxfjkgnmXraRgZLyJ5JMVLrNbkqq8IHsNdZUXxrU12YYnaPTKghLmTmq6Kue
rik8j8lWoKUH03mmxoC0aPYlohxDY/reKW72/FmUIj6z5p/gLaZSSZRKRYPFd/Tn
zQ8yWD9OO2PE0ABKW2rTBHyXmmXlNbTSjU8R154+/aR6hc3sJwUMDTHeB/c+0q6y
ppxf2cAGkgfTbqN9njaKM9PdOPfBFUktAPmPDopNt20+5BVSTUAMMUS3HGZeuUP0
gI2GLRPdHtVUzdPVa8aywvYMCLP1ty+Bo7hGFDuO1ZD8z76UMNPr7KzEtCYY4poi
vJHS66AnWtshZkq9mSylrGB9aJAPcV2ZSh3pN3RfvAlYVqX+RahcAIhsgjZnPNfJ
/2VbbceD5uzVWjAxdZZb5gC1OL6vwvZ8+Iky78Tc/uKTEQZqFlbWzhG4BYv7ZVQR
v9jCd2jyJYbiM1lU77pgmuYcSyeTz9NcUSzBF4tdWewqi/dvpY0WTyf7GScbuRf3
EKeik51OzhM9Shgq+yYgBAPQM1j5tkYuRibBWiK2shWKRJocX6UTBx4dd3awf4RE
k4gkO52XH5BkuofBxqSKFM6bEuuOxW1jwR2sMrl6NzQTzvF2dZbe/5fFAIUjDQVv
uCNV2Z0dxAMxLh5qceOJAe197fcY6+69jpN1ssjmqbHqQFzgHK4e+EzcEe3Jpr8w
MrP5P3/wFfgrchM+uXWH9nAx9EylRWUaIJ4j8Lsmd+CEs0I55CxTJKFQfTaTg2Ee
tMq/zRfc1FaJtXjccNSLYesnXCJ7m02g/SWKCVX2ypE3hTdK0ELeYWZMm5tQae56
AXANBYQdST+GmwiKkNi4gStV5ieL9n423DD10nXTY8uOSsHE0idFzgcerSn/YD4O
r72MlqBPZhULuZPRrvUr9PZmLacc53R7CHtObwXlfl0cMw0XhHdg3Qee9BHrGKg3
xgJ/c2xWQUdPwEfpOtOfl0PVpzaFxihpTbSG1by5Mc6zzzs0V9kIKKLAAhGAkZJS
7wvmM+E1xcvDif9tDtgQW3Z2NAmCZGfcZbyUB71vQRUrE1z3pMF8nXzyJgMwdhYw
man1btbZ0shv0zLRqoRY27TYHzQryEQkdBDlSECG6+Ct0Oad9C30h1SGMjwkB5cv
jbcO73HHBisfuid348gvDZc6taFkUp5MAq16q16682++ouM2tU88Nv7dKezcjake
BNdeMd1x+rNiY+N2M/9G6FDcijbSoJm07vIHbGtPkVWIc7jVGNSsc3PwKxu99Jyf
hmXP4s1rR3fBjZ2xp/xM1wrHj6BV4lrFM4SCmuQFtfEpprwkiRwHznqxAIzLsA9x
urLehLnEcxivpc5CJENkERHx4ggmG5/2ATlbjcrjtp9U7mSMZahfGSEU1ulM7GYk
gJ0K55wNxKRVuFKHRrHuWaDG5IuiXEtLZdo262qEN8QMEKHF+SjhbDclR8sG9s4K
OGllWG3E89FOaWMgN6TMrEv0xCJxQznNPnpgp/bcT+0fkQ67vK+ZaOK1ktTeOtS3
1xMLKx6zoYgO5pY9DP0QQRgoB0iBr7SxR03kLiQTJ4gJcEPyWB6QLjSc0YAaU5E7
jFP72hW0h9ZYag7RZsU9QpnWiLZ8GEAb4PM9zCtH7ZSMDppQYkJnCjtXbBI5bZuy
in0OssRCSD2zGLncWdC6xu4K7gN4MPwisKiZWozLNziOABqCySJK5oy4Yl2mEWLM
uV0VPBMlC0x7NZVWKYKRYvslrBkJ748bgD+13ZtJsKp6ecPk7l16fpnKv6EIxc1l
y3frEb6Lx1iT8fQpdD/x/GT/+jLTgbrTU4jJbl+dnRaY7ZKRA074EWfNopCH7TuY
ZIQswOpMU2WFB/4LQb+mKNKRI8HPimKvK0Va3pOyDCKJ142dRK8ih59VKhxbG1Mf
8Q/xhQEN2SbbIOZKm4b2j7+jlA06CQpG9HLBk35fO1RtLwmbfzurrRD0xv3hfauC
NItux6mWsWa+hyX1HXHKxGqweD+5XsPbBY8ZZqpnEVMkv90DA83kgCoJ+sn91QDf
4nocrwktbjzIsHdQJVRKOYcCv70hLhw5u4l3UeCjHaU+OGRDFqeqBBM6lhYQ4o9V
5ckgiM6POCAU3xE3xRHVJpleg88piTBAmgG+z6XRCfO810YN5octnTnoyzNTd5ww
cuVnrU2mRc96vBxRjL5fezFaroZlg6TPEPL9O21ZF2KmzwvlLHGhEVXiUpff5Bif
qDMnPmzQo7Kjw4oWGmH4AWgkRfWQ6hv3SWOKd3JjBk3SGlZ2/r544Ox7OcqkFm3g
GQOdmxDEiXAs3W95QlHv7PnhCOAf95EDxry0ok3zKlqE85U4LhcGhvGRDfqoOXv5
kz2ZVCiEy71FkTIeo5y7Aidybi3sf0k1S9eFM+j88i7QPBThN3QGmA/9H5xn43kJ
thekVimXV6yP46wbXuJ81Ik2IgeUh/LFNSJfTQJ3D6dwX/BObfYPhXzCekK7/g/Y
BARGm5rdF6XJwQgI0PqqtB0xDD5aJwQQSOnPMqk8wP43O1gM/uEXaMWzkgp40NSA
QzZXdfJOmCDalC7GGuZrEv3NmGfB/rCv01GWJa+e05KPoDcXXzSrl11i9F+tpjPW
ysl9BhaRBwlkIoed91fxSvCQPHwewsv6s2FDXn3ArxpOYVafvvQ3dReeEn6LGR8H
0r3+Js7MhBShVUtR0NTF1zpBhbCXCZWDqgoDf6xQlg0vb9dGfD7tjDIvRjjNcxbY
5vc/yqgmtWgzbdnK42dk8etg0CUK1SMDcK4YONyN4rvQSFpWnbFGpQTQjnDRpwUb
P4FQyPFppjfGzbSAhL9zFte7ckkGDIQaj+PyZmi195h0KuefSkoI98IXPVORLame
W0NddNv1dD/TnDQSYlZ+foE4Ft9kuHqasZhZmYaLP8dL1OHHJP4CE4EwMGgEf7fy
iMFcJEux1eALVs8TCP54gpiSII9hfTDqS7kBmVUbsOdswuFi5qzbWLcdhSZ2Dx8P
9M1XF8mAtJ+gwK1g2KOLL+MZwvFe0mIc86ihBoTTfBzPiF4gwt/ccbXfbAGQfrbp
mqqV9CjNzeqL384kvDEUTcWPRQy3gXbJ7fePXWWjVS18CalskaPyqTXbxF4dAlk+
toRJeF/90oQJGOUBl8/tjKGo54nNZqzp57+zPbdS8ZNlIz1ePTm4zPjseAkelHhj
Llc5QvskIhSFREoc45xyfFSEAwVz+/jtl0PASgkqgSwRs5K0jeyOnB0IPib8lGz5
6JC06f1LlReAB89LFbewgHvcjLP6h7eq2iA0bW436h5uNCKBDPsR6oJpBRnvEdSa
fvBniL78zWenOHHAE8aDzUVQUXzkRMTJfADlHDC9SBvr2NDBEC3+jgQEcySqp0bn
NAb+RhgwV410q6AoAnSyxibM0Ex1Hz604UtlDmP2cWeEEVyX9heW4f5RSyssqdOG
PhWp01TMXhiEKwFSRs8Qei1BLBjqoHZmWEcTzLpRLKGY0MgQskVdyzPPksz6lKue
5hbm+W+cY9FuExnF7cxbDRcublDaFPxnp24OiRk3Rsywb0rNayD8GRylNhte+e0W
rmtfvI2JSQMTay9Qs7yegCDL6PU7A/ekHFDbmM4A+7MfSyrtpajQDMoMBXR8qUwp
EnU9DRFTauNWHvfOx5FmXqhNbCwiwtRrzCuG/XiuBoBb+u9041AinBzzYkizMlZc
nokAB6b/0hUvJ48YihbKS2y+mQir3+ni381jivuWuUqzc04Awqy1haYHZNdBQZiY
9+3taY2ueGk267phqLeJlSXZaBN3hAMMg9q7o3linpDXDUYklefW108E7fJ4gSS0
8DhbbtIPC/r73iANAyq8XkpB92VZyrBkKaxTukdJRHQKgKekjGQnRWTF3vb3qMO1
/atP7pDg/RV7od1xKw8VFz8AHgxn3CHzBDOxVVxWe0BsbzFxVQWvEssSaeRxHrU0
rIaVNRd/LutvrfSxPpU482tKreGn7Iyb9ycWKnqLVaDeT/xcpV5204Rc7Tv8EhYs
DM7a22FDSuqZVkL64Qeixx/Eeiuug80GYffW1UraLWqIWSf99QTKpxjIXhdVex9p
joZc5bi1U/CAbfS7lbesDOS3RFCYvWyoI/E/673wb7+8er1etL9FXeUCE1l3TFcr
he5M49m6aIp7ylKnsH0ioQrUork432yTrq+n4y+0QQcqhciPg+dDW7EC5lD6HRdj
JzXidZE+BE2wliqgu7ff1vJkHpdnm9GGVaL7uABrjmnWM2CoVzqm5ZHhUdjiyeM7
kgh/S+krZNoOiBAthDCaBpPjhOBABB4LA1foLBQ7pkv8r5u1aJzNE6oqSr9JLbBR
Ci/PdxwpFCAc4fsRSkWZit3JOamE4wq2XZXKNf48KQhP4N8IxM5rs4r13T+K7wYZ
9jTJnqJypCRo3nu4RbqbQ1a0ZBNKp4UXsBMiNaPngF2gigSAJb+61DVqdRFXQiVT
i7b6Aw3D/yAj6bRSR/qIxX3qU6mYcZtAv8avhBJMLvY0wwcapKbJQXSWzgHkmUBg
jtPVC8H5Bh/3mgO9OIHA0MTYbakkKOtdXw/4Y0lepZMdUotvyET21EtKEQVDQC8I
L4mNqZoQn3euisPZuCeS95zpONjtGR5xQTo/cr1Owb0WRRajOH9nCnEkauWZfE6V
y5AwZLQvwQvchS4OjLm8CinxTlsoym6+ilTSdsg3z0NXzEd7nJRaogBu/0wq5hc/
lPxg4VwPXcTbELDWraZBdrEIGIFFNqIAWGasY0hqWhfryzzs0o2WkL1okqx2P8P+
SC0wiOjnZutwK2Xwhirw7JT/ozxKp2kg3C2dkgkg1ATIwq+F2uY3WpcfX2Ee54Ng
1zQpjQHR639yCgL8o8M+ThTvTJfQFO6wtaCqpkuYnaCLudntFJvGPjWn5xfmlk0I
Lw8UWKxHF5eXksdNewwQyfTbKM4wln7kNZoVanEUAIRNW5tRhUU17HQk+/WUpmmz
/SsQKasNn41oZnm7D9vHZI4kcyBTuU85pntYjGvxJ33LWl78CgesgbBXvZAdqjDU
HzmkvExpxQjAKrohLnPD7p7jSb4ErRJBSYq6CLMKfhk4+K+6GgwqYJIhviz6YxIl
4X1qJzG8KjzoNaCdVR5aPmSeCNUwohulsjEGdljOrJ3s7bwFZvHwhHlhIKJb1IqW
q2og+ZBj9RHFXl6aYP6hUXFChsOUrUAaev4sidmtyyRdcpTh5EcrCKINNjQlcO1b
`pragma protect end_protected
