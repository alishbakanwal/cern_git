// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:16 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
iD0/z4c7fDPXt6+jbGTOa1DwjWMMUosz710/WPQCD6/OWTIH31D876yBvLqzt9hG
WMwthMRZybiYbDv6eqsnebxcNNf+l2RFHS8AF0Z7sTQiDbxWvUbqT4xJ3eqRiApP
MncdvpqjkXJ1rcDqb3dBsd8fR1H1WyaO45AqTHmaLUY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8592)
M8auqihLwYYvspiqVYWrpGQ4j8HHc42RD98ZGg5zXCOk9tUSBoSgU/awSO8ONjbX
Tqq4h0sysjhH07Ous2a8fK+h6UxE8ohrXo5NZBYhKrwuJGLeZttTmB/V63pZOR8Q
Rg4m9Bmqzx1Ib4T4m9DmxBauGJ+OTj89NrB+wQVZa/pDuE63OnJeZu4CFumSaWyh
aB49Vs/QN7egh5NfUHGYiAgtn4/EhlW1PkpN3prrw64YozNSS9Y9ROHJRNmbfkIW
E2FIRzeBIrydbOzDoiKJOR87XYPUDqtFUF67kwjFR0wOBEAuTSVVEXo5+sCLly5R
kglXHTdgbAPUkBxeKbSKAvkKOryMfaZ6lfOCYflG2dK9c3fQQhmktLRruZDspAgk
lbpgdv6V9H8U7UpydoUEt8TjSEmUu4807sJu4NOHcPSI11a4n42dq8NbKZ0upTUk
OK4VCb9n5sQ0TTUkNKwtPXaFGmxyEJTssObbjruVDK5Yq5S9aeO1h6As5lpqbKs4
IR4sgysEyR8/34BJBcFCTIjIT8OepcSEYa5bF71y+HCkGozx5MaCgGjBqVMcMseo
1jCrg7NFo2VIDOkvgZyKcWo7FBjBWiqhVUBlqQN7QCjEjoBPXCfFPPFQUfBrXGM2
Czhz1BImWhS0in/c8EhQmA+iRpdYBl45JL9nBHFnrBQrlUeGnwpJ1t8H4z9GhNgC
ieT8T4QuHlEw1MZzTiqvMun/a2VzrTK7gI1nKNmymOkoKJeuk64jSXxpvGl3BjzA
FE9ETHdGKspb2zO2FHy0hDBlu9+xlJskh+LwWF2Ywe2sc9OtVkQT8YXMsLlxiK68
feG+QIeNg410HBLrWv6XJoIbcj44lHD/VU16fi3Uo9ZAiy/khFPkUhpxs7+JLSGx
v/XiwBRp3iSzhACUloqhPy4TCmRsNZwxDNDBF1hI4hLWAPUR4Rx0tZVtJaiSFwAO
BarUvCfMAW3ES732SYwVG4eirAb4KCFszV/iutG7EiBImF2fD2eMFTpGrCL+73ot
hc1aCul4P71lZLlKWD7aY9clmWEXOTIVvJno0zy3r8hjMzc74Ha1D7RUAiab5uE0
5UUcQUxQKxkRlW9nViAK+j2Rr/So6iQ/FGVuPZM8P5O2tFLM+sLK4mUPR0Ddz8pP
5o+3UOws0l4xVWg1q7XqAnbUexwsVtnTQqG06iu08OPO14emOx9YouwYp0bzJ3LL
SDG/qtSQKWxzlkfwMCx5MPbO0ea3y3ZH77GNMBzQyjcCLjIo5hz/L9KCwuWVaRNq
JxQJx+rSybi+QRhtbEMSM6UuGYyeNzb/OdfxKXI5Hz7HI72PyxE0+3xpfq2xA73y
oDyHpHcxeCRIMwma2uDqOFdMnhtS3RHycpRp5LZBwvAIXQlhZRBCY3HdRty1K7aQ
wGGnRADBBmCRJdIjsWbbu/8hW314n96IA+jZ2pU86uPhpZManjafXA0D/rWpMkPd
AMXu3FziYt3axUCTrrr4wVUrRN3XONGtJTEZymZknkSuNzc7aTFq8CZfmRiBIdWW
zKMG0oGk0r9Lmv7y4D0WeQR4nHbxV42Ngjx+SDigxzGsKuTi/kT5UfZdD66BFNIm
9w2fhvYTAsHJWrJLzUPZ8cwzM60Mdx+aGNSEKBvQDftJU2XFeB7hJ7rtQdG3UoTS
WdFOH9SlibsDeZjSN0ViV9uaT+mXgS5x3ngMLNK9rMXGwsl5hCBhK6FFnbsUELMU
P91MuqHpZPEPs6hcO+MAgKCE8i4v/L7FIs4WzPf5wNZTIDuGEKFfyyiRJaTQ+8pO
7kywuzfB9gH1GsKHY7swKy52VKFs/tKMtJ/Bcde6IhryVNuJ0YO5iVpG91CDiI1G
TwUPcOy0mmy+o/Q48xR+c+eK0tgwJ6vrkbwp7bn05jBG9soRjc+7/35MBrrhpi+m
4lPM0RiLIGbW57Haj/WImf15SG2/7f1oCMzZxjTjX+8K3NUrvpdVbMsUkX5dLANL
5Teur7CCz8qezLLUEuJUunpcMjWwurvfwE7qgbx2w921GsyBSQwWMDrX6IxDbz/r
FB1+xO9+lHwD3eueP65eXU2CmbvGCGvEaG1RdOjDDHlXVKE6Khw0um1hW8+4Vl3l
zBXlTvQUlkkLzLMUINDS6rC3n5OBFyxzMtwKErHlsLc5VKervVQ+8OMCVKVS4xjf
rvpQBtS5rxvz0F9IsOZdoDzih9LdKsqe3zuyo8VEY6+F1Q0Iv3bAXIL+gy7+vkKx
2FCyG9n3bXncSFgqpbQoMze2Vb39noZVWy5tKs6G/oTbEHQj7ELnLG7Mnf4HUDSt
T0RB5HhN0CSh7WfEPBlYfvrHH5kUcEsXiy8hIwgnBx07TRSveQe2gm33smWwFYTI
9DVSvjL5qIHXkeZr7zUNk5pUxFS5+Au4UpfW9zFBbEl4K1CAkOWFCV4u4HOa/0Vn
mpnc9EZIwwWYxl1h/nbGxVtxMa8lB3LzjxbAnMf2BTl4LnxK9GHudTsXguzpooN2
jvALOTIzNq+hCvwgJy8qLQL6PuXcHKpwApBbUp/qR0fHZl9uauN642V2gcAIvn+b
u2fivUl90Wh58MHomKM6bAReoXm7XVa2JTJ1dlJRpEIrQA3sQCcqp9iP7uWr6Fk7
5FKV2Wxz757Dxhs88vXCd8oqP8aZ+mbFmxq+5M91wkyNhgphKLt/8UPP8jrdAsDm
UoCb97Q3xMlIcaABroAsBclImjVdLCOkB+11V3xW9T0xyZm2zajAx6v5rHJP0Hdt
OcJWZZxUfbHIcDAVt0LT3MvvnP5tX+j8NeRufKtw378jIauF+EM5cwRXKV9ppu6+
KEYmRFFdrjzCVXq4yG7IQQI1yGeNME8nrO19ohurFSVWiKmZAnZ9aZQBd75LszUp
NpgWB1cxUnfJZbWafBDaCn1v78VTwSxTYNnkDG/mO3V5AhkNDwX9Cy3wQ7tBDU8k
4DevF3N4VHiJD0H0Wg6FLNtgejotsQ4hJtvFgWa0ULSiCBqGVnz0SpE8sEBsApIV
EMIcNgAouMILEfpvEgzB1TWmZyQ2aWY0JSffWbJdxQdY9vR3XGDkbV3FWAjDAUvr
dr5ahDp4l7YoUaf9Xj9rO4/cIL2rGO1tLfe9FZWjgkCQa3w7K3VqcIt0KfuZLN7D
J/ylx2dhGjMZAwuy4UivVucgscW0Y3s4O2FeyrlbVfXnb1HKxPguJkCud9B3r324
9SF66CpCGCgEfOma1jWqqwHPM4wmRLqt4ie/uNyYhnaGnxr9wHqLtQY3l11l5YZF
Z7PibZiRf82s/fD9hZql1OY+J78SfM+6e73hkkdjFJ78V7rg7lAs/nb6AbCci7L/
8nEc4aP5H3r8Ka2tPTY9dKGAXc7AiHPBWlnW3xwKkHONq9qXpqdyvbnsQ0mRUhj3
pZoDhxpTQj29Zgspd4yZcBmNHCdqicX1c71ze8N/LCtLTN2db67fvJZBfTK9TlYv
jEcKBa+yRuOV/dGLsIL748STx4vOlcxf2O0isTXJemictbiZ/V5cFifoHBY3pM9d
+/VLKMs4XtkMOwxrSOKeapbUJaKpoA5FHEl42AydfoPJ71/Y4EGBj7D6Zsl/dv0f
TaAKX3lwtS3QOjzso7/83xSNCtGv8+nyOOMFnbc38qbSXVXW7EDtgLBTl4DKZLA+
Al8SQNf1+cJfYJsoaT1WYkafgpjlQc961Hs4IVU7N7nDkBpXzgG1sdffL4pcBxU6
jgnVRUUAF0/1OTr/8RC4/xUhAIAmNXMZyelq2lpb1uUUxOJGqyE9FRSWY4Vr9Chh
fz344cwqRuYjjJFl0Ty+JwuePjQBan773x+QUjxRkuZG316I7N9SBQeApN7PxA6g
0N9W4zmUK5IbXpDfDOrdf328UhQSWiqImlQ5b6CS/fhUluSj8m8O5KZrpG+sjtA/
oF3ODEMm9DfEobpDaeJnNAn0SIz23lUK7Qc2OU1UUFrlKDmYzNpVp29/GJvKq7i1
TZJauBCCp1uN0tIfK/YuGUBX4/fsy+R92/9pwSb3Arwi4AYIbMUfPMVrfiBeLJZZ
4+M4xKeIhV2M+HNBHRe/ustNWB1Jsuzuz9R66E8dfKgaKSSv9sVJOcxAjhhoPApy
qHP7QZOsBvVWvvDZhfSKdAOxU3by2NNzlTj7lCz8dWbtZhQj/oaJOPxvkIDkHql2
fgWnc19UxErjW5wtzc/0MMFEvcgdN9IS4oXrTh8Se3HCzvk3pQgs+vh1gYFC+fvo
UMkijLfGKSv1cViZvhfXv6oyA9X0Io/tj1pcjf2aN1KVC81e8ONvztAd1Xul+5Ri
QzZUIMgOWIhqnPHzK1jnX6tugLZR+IpOqHINTOdVyBDi0KlwCxpAO9lZIBNKePWt
m6obFuQzPnr/lmuhodHJZEBloWUOiddyLnWMQ0o87HZYIEzZ/ftC6z9iwelhPb9p
Q8XgfZtyqQtgukY6t+eNTgfjP5mLN0nii3nFH9nGCX7bIGnnzUTLNgKk1epahKkE
qBk/vRHEM9MZcY50783Zl7t6De1xDbE2ONQOVl9aE4pF6JnkvOgQRdFqEF8gygMC
G+ZnXY9JxERA+H967Rs6L8CAjR1DsQKFiDIS/j9T40VXAM5f0cNKcpMM4UdoFF9z
FgemAlV1dEpg4vzE8UVlknTeIuQcJ4uMxOrovVx3TDXwAJCr5HdtFJ1kGE4dD+78
ZI1b+0h6I9V1wg3Xxk9GdZjY8ehMRjGTd2whYjUu8oIwT33dKQnZKI+k2a2IzcMX
5fiBN865c2HGi3RWiX/zjAkRCY6UpyKZlqrAtYqjCb99q0MT3hWw6kz2KLWnAtdt
kicngP3BMCnDjWTBFD0yNtmB8v/OZ5voWlsG5V6fJJhkKkTkXW0/VwyE+BR3S5Hl
qV1Ovrcbv5sn32UhMj2zAu+k54/2h33BQhbGIf2T4gPw+yDJRMDnx4TkMWSfAjC6
cz8PoBRWUudjN0euQaWGevMPW+zo3hMfQKeemnFGw0ZEUkrzDgSilffhZVD5sdhb
f/8C2CkptPUcPqITcvsEhy6FeQVqU5h7f1h+EFL60yDO4CLYuiUGAqTnjnIx6QGX
K/SxHZzb2sHsZOdcjh7T6zzjDC1cJt92uHrybKlkwIp5DPmUnPJrvrvnbgPgXM9W
uuflyaF9avYs1gJ7AVTe36cSR4siQxk1b5eX1is1Djw7zHyZVIhLaPX2lTdgKGDs
a2Gq6ciVlaTOF/pcJc43OjIeQh6SPzXYIwLnMQhJC6a/jGpaP0XVM3uh6HjF+RLJ
il5DsCRW6iVC0Ni2vBvzzAEq2nr0WhO+IUU95mZbcljiT6oLOJuYYzFkHsQOzVbb
k0Ryg9jEr/4QoWS9h7fX6JPGHt85yg5bD5Xmjs/ZWXn5u1a6yLer41AzAdoyoat3
n6GHU8/b9dJiUBYY4cQ8f6lNMw2ERC2f1WsXl7DuWcjis4GQTLADrfwq4ap93o6V
oacKGPvcySvNspHwL+hXuccrQecXCK1Kjm+xMD1py+UyxW8esfQCo8Oo2xY3OpfX
l+nT9YEfXTAnIKHqYKT7zM7fTdycOKIdKMsyfqHIV+DJgD0aWv7F1FVhmzXVNvNz
s89+Eko15DHdJ19eUrFWRIyctZ74Eo1YxbhcZYyN3ifBc9+Hw+N6/iafiPvFSXfs
3DtUK7HsPLYkjeWP9WFMO8vkxUDBMMefd8r5cg0KjrkE0E7hqfbeex3H2zzq+8gR
nFAGahLxcWnuJzl9FlFEFSwSrodRoCQe5GK5CHUcZqliquS78rY2QHT2m8xP/Ygq
zsFS+SHRGcfWqEKLzWfA9+OiuRBo1VupJZYc07/kBk9jas38Aswp9GKj9Ogd63bc
+kYXL7DzMn26TuStExdoOQd63E7QVi/Q/b5Xm1dBOrN0lCSkWOip9G7m+qcGtE56
nDkeMFVINYwEa+1usBjwplnQs7qx5bT4VxGVfc5BQbSdI7Xkoh22iWZt63CE9e4h
RH0kE238wXVs5uRMbH1neUNG5PSeY0RvJKaA594NHcZr18N0kkGy7xk1vr5Na3dw
ZPJDgz2JXWHr8sUeLN9+LaL6pQQJoKJKnJGw/D8IIRblWUl6n3IsSDKWzd0+hmxt
c3pEzF6d9MRyR32d7ekzz40jXyOYUBOfZ8OuCWn9SPgwROlgkGiB4mfh+BIytzTt
+Ch7iJKQf4DAk+/s5YSBwgsos9PEx0bhdhuGKfipoLIEXbujFoncmCu5Isvc9Ief
v1o43ohpAIzt/9fphJWuEOCp3/qmtWJlEU5vkjLt2zvb7JYz6Smv3O+iz0L/HDm3
AQ+jBfph4xYSAg98Om7p9He1ECwyPthIJRhoWukwFHXzwna0FUZ3ZMa04wE0Y9Ge
ysxjfYdu48S23kjZKYfMQmGaqsvDqMYmUezBq19NmP7nCbgyzkptTv48ZHERZtVL
qR8yGxPzieQsKrMv9iL0MMdMYjq2oXXzZMiw21tB71SkXQmwG/dhVAst6+3jsAJo
zEC9ftOj4EDLq1pQdZYqHpwHKVjRnMY9gnKc1eYuDGUosgQUtRY2AWFptN06O5+W
iT6Jvov9474Kn50WnzzViyPIPPwe+S6XZLodL+dQa3vlK8WC/Rnb68P1GCWvuLOI
Cc63ex7eBPUZfmERs3Ar7bXSsHTUGJ1osTilwo+CUCeV5D7hr5AjYghqMwTN90z0
YBbED6hePlEcNlojxEeKRWBH/NZbKsRLIp+Pc4uQ7GN31xvsj4nna/Z1ofOYYwQp
5q1BuMFywyccbmPc0OV7pzS4J9wJUPeoA5gvU4nK1/1/neCfqVaxA1w7j9BpkRdE
knd7TmFbn9aqpdVNd1uo8s8uoNVo3TkR92EKwzNr+tPCukpEBcukg/XdoCKnS5Vv
EDGFsfZsnwNZntln+rKdquexshuuVcBx5FwTmy3pZD4j3KbFfIZ0jyArM2Dgvq74
coiZKOjffaw+Faftm32+C9crJeaJSABuk91cH8LlPEsUed+SPcRbgLIrv/0SLeFL
rb0RiktVWwkPTiJsyahkjGqzuCixeH2w7zICQZgpKcSa2RCRpV7pAw0Ugs6gwiVz
iebqyBBrJxALu6o16gPLQMwCM9/xh3xF9tjw/tYxYTWU5X3x4D51NlpAdtaCaVK7
mKgOPziOp5xxUXPC842ylP2YahnVVZbbjUuHVatBvlRJDj6zjA7lS0y1YV2xI0XP
G2m21XKX+BmmdIJ3KFdYccj8oIiJeZV5fNAX1p0YMWpUtumP+EpvVfWgpX2L6plj
cV5VgqcDzhB+FPXxhhSmq0xmrz5N81o5OgEQEZ3iJT2E97aUmC1JqY848tuulKNR
stWucIJmDXB4WFK3WYNIo1DCmeWrO1vKN1PKBwbS2x6zPYqFL9aQ9tOEZhCX+4OV
Wxo3Q7CjbM9wmDwDVa2E/cB0nt4Uc0CNifXWxtNSIcyW7ad8V3HuuQw1QUTrVpA+
uKfeEi9VqfdiQ1SreWpAdI1/tvgvWYWeH9AkENG5c6AyDpDNA+t+oqQ386b//AyC
wUm6kAMEBxBMggcJTM3tlPw0KOyS4cKhu+sDSnVi08Et05OB1uvHIvTxuOqBHBaV
rMUepcqPea6+Ju7tPgbdtRf5QWEsb6eqL3J9oa1EYbbgj91obKD753V3aKjzpynM
HwVpFlqDefS3XIpqgIBX3Wvu9D6Guf+QJK8STadTwyoR0ZlAGXoorZjNt1ZKTURO
Wp87THM/WIrxvStoLnC8eYvOG9cIsZV293KFDkqGJojJfCLE5gG+tQd0hsqtyNL9
c1lPTpII+tmLfkLDFn4pVTx88+7hNVdYN2DkRCMlfZBIvM31RlH1N8v7Me7x7KMe
7rOk+VL5NjLkpvNCSp6d99S4fSjX+tbLcE96W9SyAiS6IDlXzOvXzD50tGCkmsz+
KYS1hRxKF9EjJpBfqfLXm9LVdpbnCcg/VGL5zgKMzIEho9TPGlVal+2hzY4BDCw5
dVXuM2NUzYIUYlgL9dfAicyxnMrABXMTsO32CV4frVET6SEPcmMctfxCgy47Wc2n
WagUwZc3Dekg7l3wFbgEkV0msMvNwdWkwkixcNlCVhm6Dlt2G34M0fJ333m5uClH
aCuSvoo/ig//yU3Gi+uvjW9ZYbwHv0I7F//itVOfkVHPTYPOadg0l2h8cri/Jb43
meG+/gXCSFzoDAERUU+bzAM6/y4coufPTbPvImhijuhradmGQaEhaC3/b6BK3D4p
KZn81Zs0CvFttJR1CGh+WMtWJWthky+Qcx1o/thHRegtrF1z7HYFsMwG3kM3ofCb
hWwWuXLWb6HMaLmXXKqhOJI/pfHJHJ+HwmxAYw0nPAaniz/iAyqjvrPDyPtmUd/I
1b7TOFyXIi8f76Ks2K/V2EaY8eoqXHqXCDJsSKcWFthaB/81WNv7N+DgBT5Lz/o8
rB1d2NalXG1uv/RFJUNWWo+WlXjLx7uI3r5kdNzKCQ8AUSgqi1Df8OblElzbATNT
UXKEF1Am1/geQJ/j2avjKzbqYRK/cTlD3ocddh8aWLeJAgpRCU186Qf+fAu5nWVE
eYFyxee2fKaVDwKL9tsyQ/tu7BsYiBWyLEtCcV4JvCzSzpvnnW+Rp7r+xeXOB8yY
+uEG+qAvdNPyQg5HEbNWNmgg/ltfHlFd+CPvJ61ixs529WgMuAuOeZ3/kCy5HP20
eyWVGCpk4snAcdevnWWjuh+mLMuH+Rxti3ybsWf0TUB3waUUNczopEHaNE8xN+RS
5uJvI9v/iokkNKhxFRGwwxX2pDEMtfQM6u17FkeL4pXdLSV3IAJ+CKJWW7NbMF86
wFrAiFXKJXigyf5kzxogC3bn5kYL0mmpCW+ml4eYHmtNwQgw/UP90O7lv82kXv/o
2j44ygWLiLqXczs7SshqyZoZkVUha3sVajt4Yme41BoriowazQsfGBNwSOonaqc3
zzrc8JkZGw0+CiZ7OB4v0V+utKVQ2Mv+DphV5FV78NK6DvLnzF/EipcAZvQtoxct
1o8GnTJfSjoUWeoocvgWQGf4+lcFl9A5Iw3Zcd1ISc7AuPbo8QaZswI7EvK4ixlf
lRr2BT2X08XjGcN8fXaUF9l6ZoZFqFqeSPexPvcpK2m0Zxt+rYnfHK8XLCnd1IqR
QJHoK9ZN6oPncLxwcIf3t95rM0T/VIX2hk9ptHsL3bYihQv0rbZlbx+sK8BmchYC
1gpXJqKoTE4k2Vxvh5XSLChO55cRQ42ehUocLxXnP0blBHJIgC1psxgKWMQHQaQ9
Bi1eQc9UthrLs0pDgNYhsaQcapCCk2722cOtrlMT3PL2wkwsUyNX1SHyXTWedCkf
DU45LEhcJMxq/HPJkiqBtm/sHeKuyqL1/CMGaE2Wi9wEF1AVl/aw7FWjBWiT+irq
Tk1gmN96jTT2DlpgA+p5nyca/Yx+2Fbctm7733JMmhyv/wYA7879kGf7paJcSBpJ
8BWQT5AYiwSRPuA1rQVJ8dfWprsTCqjtoys5JvneNxNdcxp0cqi2Pnw798U50Aog
kAE3pUa2Qsd4p8W1Fa1ASea+edMMJfaxjABp/6v7sRsSJZckdOWGS4apKsDRzS8+
UX9E27wqIwVryaIVBtHpMW7s3OrQYn0qe4QSlttKuHbFDsbTDNF2g+Gw1zz9FLSx
xBzoWHheSeidFfc0BOgOnJsNu7qh0GZSytNyqJMuxF2EchUIpd6MzbQIibfBbo2p
8XCQY+AnVUbgY2XMts3nNBwVKt8QXZ5hnEKVfXFkj1lP16LsYRo5/T2PYPO/YHUB
tx7Vg4XfYfh8Gu63vz1DId+HlXYPjgUIDwwFsSCdQMgIesE2BXYWwjRkQvzIQwkx
oXuDgGJjUAB6qn7i36S5UeI45LrCX6PvqK0Z3VztYeHYMtaq4HiXfDmWqVOLEPTL
aEWkvuIkmNhTj34jyx6M7Xvj4QbzyWp0fGaF7Pbu9ukrSNFTwSiI+7ho31LtRJ9x
a070Wd0vGgb6/E+AdLLnVB8slUNmJ907Bd06dC30pEHeWkrjefPCRfZFcLARvTz0
YeQVQLfB8nNrBcvBdJuQkZ2jzg2fpV6po1G2A8hVZGhvJn6HJC9NFPky/Rq/iVJV
BUyOGheDAmea0DA+m/5cdpotN787Xd5RqGZhhDH73DCYDc5rE/VySmi+VuTtE7b6
LcQKkdu1uiL7GjrkuqvkZErbu5C8n3DbzzgmeEK/kVfdebuWV+1fH/nbfkNkqnzZ
p4ZcppGXp+xlSjkYFgCtpLgS4BMhH/IOAVCTqa1K/fAkcz8ru8XFGNeHRxTfPBxa
FtELZT6mmyWDH87vdAdv252Hde2VprPHzZevmuKsF59b46D83TUrAWBNhMwjfnjI
+Mx2wUPcHlv9mRn5dw1JeUoCL21G07WEJw757ezJeEdUvsg6BFJC35uQ1dArinyk
JIK8VKsxV1CdBPo00jQIcDK5vOV8ZeZYmGEvWK5Uy+oeYRGaXBLgmoc5M67fwFqn
K2jm8bankShp9FRrBvCeuZJe3QP0XjFjWmw2ZcC+qmkeBnJ1uSqeGiJz3M91zroK
BmF8m9Mvot8s6AFZPvUInkKpoLszWBOynI3unqkdlGNEM9YPjLDp4ubSMAIZK8kd
p+fNIuKChcVjXYOMceLgHnSVU6GbK41kGjoQwpFR3VRGMW+YxmS6ezUvZmKh7iCN
fdmfgXeCMcI78rbjRIxqTnFQa/iF13v53AU2b5HSHSKbsXNNosUyxfd20PnedWS8
BFZILc1ixZ84P0ScSWCLCruVDZuVDYCxoPiwf28cwhW+qPuzlsi2tBd1N+jjN1WB
N/WBvFUAso2jy7AKDeFfb0xo49IF/9CT9QFhIm5Rdgz6qG+pb8DeKMT5Q9BOAhaK
+eRz2DF/A38Rr4783Zc8E+iZ3u5Q4gl8kNpY7MXste+LNb257nCcxnyDcO3sxMnt
Gx2aMPExAPmzpzfxDWlmmYrk4DUNZy19b6R8fFRySXCT4Z/xNEx4hBMltFOpLsyJ
6NPloNqGQMQEfmuD10ihQc8xiI81IgUGvVx+bs85UJj+yQNVmTSAle6q7kx0DV3h
sfmlXHEv368jdok8XPjKOfmXhR7qqApKmZpEWEm8NonUTPt8Gpoupv8zg2YSwP2h
wugodJtOVP7FXrb7S+0dVEDp1SkMl8QizRHlo5yZqA+QfMz7bjSWizOAKugP2NFM
9KF7gmhFz/egF9+r8BltatvXByCyOO33ei/rIz+JrZvv+sylATnwMXtGAmG7Dr0K
vqe7P3qJUlUm4rOWMFsIhCLsjdAT0s+s82ECWd6fEEWouzwP6AbKJ7APGm8LB3gJ
VwkC6GlmRl+eYIEDmm5mkPDBVN9HksyV0uIyGPiLfLjnqRwKd68W4JFpCPVVJ2vr
tSh7BLtx9hS4U4cBvnUHM+QvB2i4DM0QG3GfzZ8rx+ZcDLj+KadzmEeFdpIlj9AC
Qourt6BZDfidMyG5g1J7EyZ5GbHWwl5NQflaTDEI+s1puzXSCbo98Y+OhcgqwzAH
`pragma protect end_protected
