// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:28 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QWTXT/ffnn0U08x/5fSFLOQ9e4HiAsfUE5viHu/8FHFh/3W3yMD6ufu8UdlOqGB4
7v0q/TLK380ZGjyjQlx7YHwu8z1tOEN4m9SZwnPwZhZVf7nij15JPFbXlGtZhuUe
bG2rMZbPFFQtWNp+IbxPPOY6E/Np25/VK0Rn0lDGiNg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 75232)
ojfhnHND03ZTEF60Sg2mygP3VJB3IkTMDNdKOlnbIgHJ7v73LE8Kg56yZr2yoGKb
1U9BM+fhmdzMfONKuWTx4q6NnkMmW9TB7ooeFh+jwJutmHcY/QGkrJAQSf4vWxvr
JjWQyiV/Bls3nlkVgs++fy18IUXbdYEE08n/cP/ql37rASnUp2JscLO8Ke52vuue
vXM9jELmYK4xKY1/4bus4EzY7lPZWZ2D4qJ45ZwiNzJeNM5udXYMtXIfTR33W7aV
qy5uqjd5KHxnQIRyoeH5pmcpka8lyjuG6azYpCmDUQaSF/YHS+C5Hi7a0X29aOFi
1qh9SWC81KoO2C50LcD6Q7372IWhlGFTU8qMZ3mKgQzE5B5454KWVDo4LS/sWbOw
yGbCie/i+hKPdxIkqE0jf8pb62FbVWZSpyhvnDFtX1S9K5X+/mIBn1TWS5C+o8Jm
lqiPBMumptEeDAjuUp630I2w80MblYZEthPGfhjf5T/+yzb4tmuDzg17s2BaCdxi
9WnZluuAy3tL6zAr5mGMvPKutpGkJ2I254gyuXAMcnjrWfJME7/GsTXQBJ3/uM+v
syl+tdemBKyxOjDvioL6VR2uWpIhRu3GHYuYjZMA7j72qvaplhLCsP0q//ZqIlZg
eBvaGz2UOSblFWLDmjlW8t+a4Up+S75BV/yx1O/l3ckT4LaYq0yKvpu23IaXNI2T
5ENgr/plzlQM/pXEKJCDv6bJ2Nma9RjB4h57+Tx70Epqhu7DDpqqSeoSpVBbs7AX
kUQ89vdKuT9hGPIyXjmVl+SrQ0DYTW0INTwZY2TpIM8reBFlUk+mapcVaOq9v2xU
BU/Zz3YZgvD2ZkROxR4UsIfh6fX4apaedrfXPEi8fL7IfaUIqJ5Qc5H02GfqZtjM
ZtqTfutYOd8qPGvp4nq/E4UpLPkdDI9Zz3K1pF1304Top4dhIc463jjDr7MPecvG
Q6xxtgE1BVH3dBZZUUX/w9MigB36BI48SKHVhjRQsBEXTm+if06Qwji/KdlJKckz
1bCQjx0YkNtuWU1DieM9VyT+GJdPeJj6jeoVKiEM7xqWilvBqoTZoWhWUtbkxU12
w/k7yJlw7Fo/eP0WXFytomOzsGu2tgV3QLA/Hklwa0g2gO2tAl2x+SJbQmbr9XF5
Srkc05U0XwUuchl1T+XsZZCGcqxvYSIiYLu5YKA0LGU00/EB3QtjcaNzZ1LmfrPr
oXavxhyy1ITa4mq36KzxEwc1Sw1wpu5xJNBt9m57HCEZSzuSAKAzeryDlAOJOHA/
9ouwbSpogBaGxv2pcqL6yPSmVkiqeT1hMALn+/w/nLQCt2ieCIjpiPvbdzB3L9ne
ac4qH5P4/BS5+sJ7M4fds4vh/WSe5iTK1B8PQrFxlQN1Rg+Ar4sqCh68GpO9HhR8
mL9LLu5PtlErur/MQttknwAOqovFp6DCDGThDsiWGL+n3FzJ22l2n/5bZH3ZUy4m
OnoIV9OPp1TTUVXDWieqzEG7KA/E9Tnmr432uBfzkFbVEHuv6VJVlr+uu5/UgRmo
IUgreFX6xQNalojS6icIRDIWulb6URti3jOa8nAxBBWRs2l2d2q0jVWdZKZBuszE
W1FrP22aou13ZxrUxc5BpuN7Yn8m+zRBFZ/edUg3AoaPBBmsGUElEQKseLtmfsJU
W/ZneHngKcI6P8Avf+Vxe9+nL0z2pxRHmmZoSMK3RY2cbuFvOUjpZ1a2MFEffYdv
tsS19dRW5qHjX5ruqmxOtmshtPkuEaydnwQ/5BVmwhZtKkMH3QEd53k4tWN101X/
EpF9iOtIDOAoFRfLl0lxKFz9MytEIuibFgR7RD8cEERlu8gW4nk4CDDXgLqnq2eK
fNzatmJcQuI+FGFaeAR5ByveT52fiH0vGUSxZOpNRMtLOQI/FQ7eCZjnXaTzXQAb
JdQ25cL99DBMZyUgdXFnFZdNTT31IvPO8RkJPectn8RwpV2O+FLc1ZQ1M4N5EYoa
efaoJof4pe04Wu0DPw/1N+Zbt4fBSCKaAYsZQ1sLSZtaW0z3bRhYGYI0fib58+hd
RmmMnzbgST3vAcwzUs9js8ans7dkQ76KUp5HiPzr/vv//x80pROojj+Bco6YwAbv
d4ULGArbl/yDqkhAO7Za/fGXcmQ30TkRhBdk/vqx1a5vuT26QkmrTWV4bTif0fwQ
zX8IeQYoO9axmH1e6OiA5ztFfokDU92z6R889QUq9uYnZQ1vlYqT/QuMdHNorT3T
WgUzrKyAofPu9VlP7SsF9GjU50+trrtmZkpHANc7XUeBh4Gk007kiTFerOm3U47m
U1vBBp3rN+vWsk5E740SS5wLHUbbPvVGYWhi0IpdBpZBEGvmf6p4UD8BRE6OF1kU
QE0HryoG5JwZD5YCL3FqHFa5GIjiaT2xuQIQzq2w5eHb7MFWbNxaWTl8ZMk3PUvT
BssLu0I6ECU4j2cTxrVUTWZaLIzXXICmjfRpaWO33Ouyw726oyQNg+c/wwQ5WIVx
Mc0thOzM1qfyE8t3vBqyDYblxAIdMUu2pmidMa+TonPRNLjy636asfCnaTh1y57b
MPx4cJQZFzs4CDvW0tWQKsR6JEU0iRIr83Xz4o1E5kKbPTiXFtS2QXONh0mULdwz
IeKz/0+oytG9oqiNhHXyknq0KN54AnsGXUr9JHpouGu5/oS9jAiPOnfSO3eI9/QB
uUdORXG7B7FQx5nmniH7pL72D/ACGqzhvt/LYABUOuU7lJpIfrslT/pH6JfyemR5
2N/zkV7Ioh5Ak05N75zU7kEOS8GeTm0L1SayeAYPHrIXn6E5dDtUt8ecxE3TW4N7
r6iqRH22ORcMd0NiOm6rqO4UyY97WJdPQq8eVAHxNV5mHbvaB00ZanFDWRUEWjGN
P7dcl+KwrZSyN+93k65JAOWSbI06dbPT/Bqph87NnYzGQCQwgdP8pypZdfKvdKcL
ccn2fdxr5GOf3lgzDS1jaGjoTFjX3Bcac6Mf9axqgPHFCgUyqFoifF7ZfH1HnIgr
7dx1CUg3AQljpf4xMAo8RB1fr7lVOZWHnbBV9MBvzkbZRW4CqFGOIzBnHcZPZmTl
F5qeeVp9zcC24XuDAILHZgCDgIPBIA+54uPOW/CjGiuBfNTNmOxQQF/66cTVF2ab
iGWdmQQqoR+b50sB2MhbLTExKsJVekHnzuVutrltQibVEPYgDBxsc97zH7UnD+/I
8eHdpGnPLlvk82xdiPg0qjEFBrPQZE+46Uh7otaVF79d8A5OqIIMUgBLBPxuVW0m
Zi7DaM3BH8tA2WnopaGLEA5VYieDpaJ2YU8ELrVsAr5FY3MIpLpvIsNljzvFwzzu
LC/IjIOvs8YDU5YYSN1AMKRMDdkoVVE27JOXrYkeFPiY16F+15HFeSMW4XuNeQGI
x/ocgc1fDzWYkua2wBzjg3IMUtct7C76XySWGFpANGkiVgp34GgUqsrFZtaHGNpD
l4c7fvehcCAzAz1yHa32NM21cDjw57Uy6IVJofHMSDqX/NrxcB7H6YIx0hNmrFF2
QzYvNv3wyq6v1lUtMuZyrLIBJSuTqDXH9X7ieRvKjry62hIT44UYmIYtm8OYry7k
1IrV6/jCZJgxHRFBskWMOz62Zh7mLRPvsK9wHmajcJqBUic0yCRemHWiaVOXlQuP
UjcsLxm8mzLz7h8zDEzcOU0gJm0hCFm/CibILV/ry0+godr6mV+7izChFg1D0/64
beSD/3mPqGhr5+wsjGi/tDPf6LWNNTfQUwllttvSODzp4018FuaaF8zsLiOxgukN
yD4NZ6PQL0TzwkV3jzKOtu8nUC0YFIbIvKL2xX08iypc0XMXbuLTUKxOd2Cq9CMN
1glc2+OQ7VzdSqoD1Kezmf1Qsuo75Qi9oy/bC0YvjZWCYzDlWqgFgPsdWq9NoBHp
vGwyuNYUZrdxLvSZ10OcUz1iMpDOdtSvEk7qp266/e72FwaG4yZ4TddMS4rPRZrG
3TshiswYlnPk5sdov9ZgOJaNnomz+MlvghFqE40XcciTw9nT+nT3sK8eOCzM+mHp
ozpBMiMbgkaskM5P8HWh6xHLbWXyaCC7mrX0OC/h4tEAkKz97kScSaCRMan68tfI
nwhKaIcYYqO15p38q7nePBHpwmONBVmAk7j3csdvGR9KdZ7qzNGO4xesRVss3x8E
fuHb2eEacm/G+SMjrSh//VrgaPXlnYPwCJLmLCj1a8MnXEkN5l0yOH0i6fpSEAjO
D6ESAYwcS8deyzPCxwN1QrvmtrG4aIuo+b9BSh5vjsMyA9WFp3sYKVMrnQZXJZ1t
XRqlWxBcCMe0NEjpkXy3gPiH1+VHvZ6vzzonzGcSqc1qtMS510G6dQvemOlT230t
uz/SOnXxGjMUkyvYG3iRFjpA5zweV4F9E5FdqhjkwoYh2YTwV/de26zivcBQy5DZ
n/DZAAWbQFspunsweh/JTCFU+JY2a0idlQz9R86RjEyMbyrcjrVYVpVWXb3+H2B6
aA9wEeOGI4Xv7ZZqwqxom2dV5M55BjrHVdK0g1JrYuoMR1gMSv5/jjdfjwSgWyRF
gFXR2ionpQTUM2mjAXwHWUWnKuNUPt4rb7gFKOQ43jiCc3GH08vb8D0UlclR8QB/
17FWtLQkJBRz7z0Wx2JGjQOtW5zZHTVl3t4G+QNvlmnMTc88Kcqc7+R+ceuYf72M
/DTy1Qlclxl5Y2OT6mbojIw58YIopzx2KRdE9TqhrXBqmU8JeGLA07Nwg6mJZP8z
HvnexNaA5NAeJim58Uznux0S5Whc3m6fLbdPSiNoRtKASL+Nwg9DiMuDIFg1dmDJ
EK8YSK/V6gSx+W+Pwa1KyzwCOkl8l2mVyfBhkaN5JZVuyQXLHPEiTAMbVveN/wY8
oCJ6dJFDl+PoYtgVI1GuDbNpyy5dUdrSan2wBbDPKElDWisvJNEyyjSee7iN89fr
mn+voQh+huhlPLvYbyGZcqnEysMPB9JGIGMJmkPh1Wk/uR+/+F0KI2X/9zw+B4lB
loL7hUtpqBVYa94cZv9sMp/PVGCOMGCK0aJFw5ogWlWBjLDakRh2ZT9xtn5P+s66
r1oeEy9o7/F7HgqDBJkueby3C8sqx0Bk1lXI6HyGMWZl+XGJ34VxsZg5XrR1QMqb
ZMCiGqX+9bkJvxI/3wX8ZwCtbw5fYm+sQdhYcQnqV+l3JJTESv1XAw4zDLrJr45A
OzohhSODRtZGnhJOZQGjpZeLBi5X+A5qz2e8EEk2K3/bkNylfrGfcPngULRQyXjp
esUC1r09vlsXtdw0a6zlmL/nt5mki5ZhrRAUsU3DeWA+GQ/2Ee2t0VJ74lKNSTbw
cy5UXwtb9Sk2oAtwhmAOij4Cv7j78CZKPIBtzLUsSNxnB0/KIcNGNhUucqo6aJiw
LIXL5GuvLQMul2PlJ0lOV6IsRRCd7+3/a/CBVjHDYcK9VH7qY9EgU79UwqjRJXtX
dsPLm5SkrZeumEInBFUcobfBkKdVyWAiiFmF4ZZ4PIzTtysZFU0Ddv9UFwzoC2aJ
NyWRilsGa5W9xOLQGUfpryZU9xO+VhQQhsZ+hbZ5GVQoFIfp/5cO01/RubW5SC+B
lUhkmeu1yWNC+c3fnbVdfDz/rKnMQojVsfnBuHEki6urE1n7aAYT99j/aTFNzzQy
mIGnG1bDzK0ICi2K3Vhol84Na8ZTkeR9+KlP1l6dr0u8YLxb4VzLBR9tR62RKyyF
OKxoqqfyGsgxBaGbJFgyPgHzqTZVbEq1yL2oDQl97FKnxhq6qdN9U/o5DwJ5E9Tr
o4+mJ0LCi8tPk0b4hY6/k+KuRb1vdVOw2LaQxaCqtk39BF9CcHnz8oBBAj12HLN/
gfHkFxTcrapi+Jo8+RLVD6TB7PjaGTdL7AETV2cik1QrUF9ry08xxddNbnNQo5hC
vIa6JkPQm+ZLPl1ESdvH2YHfdF41EcQXusYVCarz+Kidg0YD9jWMbeluUddbUVec
AMQBG2fsxK1iJSFmQqG4sXEjTQ04OpGaPeawaRxVbFkOzOEe58HI7mfDVW32XDAe
0nSL6QFKuJgNQRo8c/Xtreo278BxpTyW4J6kPKMqTnneonPIXoPjrahF9jlZUwuC
gzEhQljhBhlgG0qxZJ9XSDS+b/GLvb0P+2q/VTujq3L/DFVD/HAfkxb2WZZUdeei
bkG5oplROpcmpwvgXwXFRKhcIXkxYSKB6WE5hEisi8Tb8ggXodB/T0gmycnU6x6l
QjSuM2dCVKUbdVVWvtm/QJE1+hRXzaFFba8e1ZfHoHgeaH5ovg3nzhuII6ApmK5Z
K9mSomoUg9nlIbrQ1nMA4F4PnE/fcUI84jb7u0Wt6wVu/Dj2XoIYLG66q1sr3Y0/
zlsiqAsDJFZnlCdbuTbYv/vE6N9EhRclLo24bexWT4t9/scM2qnLAF/8Du2NAAF9
fhy39UcIyhZ0CDc2Jv9CyH12zGHT+3BchSekU+WLpP91KTb5Tn01EVuMBtC/ywSi
nLlQwf3WyYZm0dn8alqQJQUIRMbB632Gfo7XsUAdMYkIyk+u4yI33BcPyvVX9OEj
uUlX1a4bTGcO+lMs/u7Ap7M4+M7nSUF8qXMAcVCZ7DcyPZENKRrcHW8ZfOZaeJhK
/KyRFJ0CCXGp3bQb/BcRBY1lRK5dfqq1Z8LpDSSvdlrg+8M71xZwnB/Zg9v+F1jL
MOTITqbubTwXvu2UGiaY/UHg+GKPX+UL5rWkwJmAxLKhoBfJBQWAtjEHoYpLWya/
xLPDnrBbwtooJ3TFeaAqU8NQWvGda3CAPF1zS6uoFJuFIIFngPdNiWpIFM560bg4
nRuHFx1TQ97odEtQMmYITaMrNISkGPig93/54OdpD4TVOmKFKvRSrLj0NtaL6HRI
5LYq/GEVr2/STAgPNT7D4i8UTavT1fgH7dGoDUoGuNmwdTfSPa5BV9vU4b3scYud
qSWT/bZmb007FMDRZLOubqPsTymnOYN01uJ5aYfLFWod50rLVVMGQOQoltigZ1y/
OaikwvzCs5/EcGYk+L84ZB6Nt1FpVvHPu/37yQQbE+aYmQr1/GFj27yfWOoOfQfC
19DyRT1lstfsq1PSxcIgaTUa/6YRsirlsuVKBkqFtv5qFWl+xIUEriiuwaLl7eT/
q2LL5oFaY/OBIv57DBCWPHXVFCGWcj0/aSLx5TNkcti8EirMd6uMk2lL0dwjrjF8
5dIMFP4fAVyJY8gaplbizIaM9v7SI5qoQlXpNGooIhIzT9Ry34t6MqxURhS2Snnb
+1aZ6NVXtdZUY+wHJS9h0Z6fWcuB0s01bq2ljEZu/Tez32pRemK6AFzx5WbUT5XH
pNJvb8ve1z5BgQoliGJ9jbSEUbrFW1/q50K6nw7zWw4ZaQeDvHObUy879NxrcktN
kl8d0tPYH/w25NhY9p7Ao6K83qPbHrNzH+iyqVOx7ulpM/FBX3V9t3HtMPdBgUXg
sk+epJ3f+hywa9RecqWxa/2lbJUjTbb44BozUIMfaVpGjQQlZZ14H0yisi9SVot5
ebBLjvHeCznZNsd6fMgBzbjoQt2Rnk94yLO5U0BjhSt3RTnBUuKnm6t5lkPrpu3a
Or7zgiccRgkhyOoC0L5siAt+Cc1T6XbMcLfSre0xSApWukkca/ASYQ1LdH+U24xf
+sU6/dJmpYLhl360h0fDBRhxWd8VN5lz/qAWNR/FMy9s8g0aDMF+iV9ufkfIz+dr
Z9kuzAZYVKyUitXZg66MdAWl9seQy3YkFejpH6LnXn3q8XvunSv/JloTJBKCWM1m
YgkOrKl+LdTpwCtSBqh2CN0j+Zi5WoRm/6tFk1tZOGY3pSGd/ynVQUiMvCkadoAX
GcDQmFuFFHqdBjpm6/x1SYED61dEt6rDkjkqp1B687zBN5o0/7WXwloW8WSHQlRT
nZ6TXAFVDHDKfvUaR1N9fH6u90aCAsSMWTr2VNK/TAXsDxIupobtXSPWGvgQq7el
NK5MRuffEKG6KOVVW9lQGjnhYHUgsgycJdGiG2ops+vy2AaA4xNZJm2pbk9x7CHA
PUxHt0IOzi2LhM70u5x3StD+q18hyJd8jmxstPLQn/yS1FCJLVzqaB0RPUTXNZUd
RGvpX/MzQWMo0du+FM6o5TZ/6dDSgx44AvFpCkJMUyhZ6oIKc5uJI/C8Zk0xHE0b
dvZpL1nyB+bdJfMNSdeC9Aey4DD+Nw2gbCFrgfSlgCxPBDoup51YTgzRLU7NXgtH
R9eOqeN6Gg5kl4ijhHaFS7WYU9y2llxaF2g44H60d2l0dX5ojWTPv98T2mJMvUV9
rdDUkmcyspLvOVU/MN5op/+/hQgojBIPjdjKuQkY2Ix5bN5PsZEbN4SnRkE6tPqk
bHcC7CPOw0nyiKz58Z5TK4d/XPUJGzzX328oqxZ4pD3fnQ5QzqFscM5ncSnofmM2
q/B0L4vfCEPSZ9qFlNCBOOXapdRi+HjNwRPo83J508jfMDCkpo73pcMLFJofdMsC
F36qGAXh0IDdpTwaCCM0rAdfllgm7q0+iy4swSZ+eJseg2pOHU9QgzgiWBaC6Ilt
pqYTUDQDRk4F2R7fZD/ikvhOsovwa4PTgWpZsFo072VmjuHgRZNPTh8AdumHyHDf
VpMeMYPpJU8/ubtz3k9yMPPTqkbRc+OwSobqRdWhdXwAbltexVTVbbsiu2VhVqD6
f9owqwt6cLceUZrzoefZb6K5aeISYRpX5yqp7Ea4sM/B+SZ+5pCQoqF/aK5zgTQp
vL5nfpkK05xWhfmM5b2fxa3ElfONN3V+grvC8yMgwgNWYVW7EhOTnGFWANo1fEEh
mcGIMYmBQyouxyhrtvY5260JaFdv5Y+vP1tmDbOF09AwEOUr8efx/6dyZD98VHeR
Anw2aguYOydqpV6MRaTAr+QBDw6C0uIsO1wUe9DTxhzHJ5zXfCK5meiCE5kQ+Xaz
TZcCqDHeMyvu+ZEO3NX1ExgYmmPQ2k+rk8PgEBfn4D+lwrSVwetvnaal8105O38y
Q5TDGJV4Z0F9rxRC5aUesG99Nmg3Bo7hC+Rn5bAQ1vtUB25LujT8MY+bT9VsyF4T
W+VPM1/2TAbEwa5NVvPV3tOoYxt9U8wM402Emf67N3bjsbYRVOXG12Rjqcs4w7eR
YG43ALcLru/T0Apx85iywe6K0aHm8y6pJFvlB9QYawHVFfFYcNknFIS8Xk9Tb4oq
1v3cjesEBTiosRKvlJS/IbGyWEOECm5gdhuUxqYO/Q856XqbD5e5VstGIKIqgKNf
vG04DH5npRVEWWjCnhmPZgBPjS4HUfGcYCfz4R17M4e/u2ClYBOzmGW8LH+GJXog
IF1jaw80vTv55h4keIwAvnfFLZo8CwNqVUB55VjauKWRpG+N2+El6DshFIkOuMFT
JdO83PoM5NQtACq+0fkOPVHgNmbmtcmGo0uCvLB8XnuSRv19iBimoX/ztzDWZyyb
544rWx22GVcwAZWvjAJY4TaM+rxnhzdAckb2fw624RK6la5YCDKS01Xt5tHHZ7ZK
Rto8zW5iXqKJv19sKsavGX/XF/iSLI/VXmoIYIEvDII1l5Fss8wpw4JVckoxAbIA
IB0VE+UauloOxLTuj7Oi6Xrcq0ud4208QaDpM+4nv6qsCwPZyC3+I3wgyyDHZWYw
iEkWOU3mWL4z4pLLL0d6f0uU9NjhRyEy09hDIsqCcOF0P6UzghWq23aw8nL+WIGa
tB5wjDtG4IesJIGM5Wvt64A5yu+KjecO7ITU20TjuRl+OMj4zwhcASuAosM8E0ea
oJVd/KrX+6iYyCTCyuIXBdW7BHYv0QYXoVTTzyNJFmtA2tvbHrQqpcDtmop8VgrI
UUVDNCtSyBmvO8raZDaTivVsoRIOWJHqZQ2fIVz+sgwXxO26ye1pw29rRUcMW6CS
Lcy8WlNmbaYiHVd+6t4i5yHUZvVkNgcomrzlKQjIFgXeYF0Wp3dyIyu03IC+itB5
6pHNBrLDNftIwafgDYhZvdjDP/UWmCmfYmBemnCg/I5XZZFuRPa2TM0EdgE75/qE
+ZSsFaHE6c3l2Y+aZZuNZE2oF4x9xA4fFAlviOtI8E7TYCQA3+R9hKDfPGtkJS4k
JjU0JM+MCa1iNHDJKZQaGpRuT50W3kc5UH2NBgM/+Wqrg34UQBtiGPGz/qTpjiJe
yvwEcAcJOABSjuE/tVmwoQ2wTP0UMo6TEsTJk4S94JklBtZLjGlghqi3ChDK+R3g
a25eFqpfoU6X8JNflJCswSm2GJJ4MesaYM0PsqbmeyNBr0gHhaoFlWCqFKWcgEAK
IdTJO1/AVxnOn7LqaLo31kG0/BDqJTQdlemeUs0E8Z7YXdlog6VUuw1E/jXHJMaC
Sru+sciVJ6iyJ84XqlpF0Cdm18XiU4nTwnhL1m43/6lLey9StpJe9JL6u9k+y7ON
eesoa7eNnS6Rj+Sb1r4orRgtTPg+RAqtMQV3KgCJPKtqpeadNvZbz/xlCxk4X+Pm
bwUwnQbG6kjpX0Lis5z/u2heH5l0afLfaXR5ByNP26eAHsebf/cPNoFnYMPP7qG2
UUWUKosWalGXy9AkWQ1y8p1YKSbVro0udPjohJAXMfuJCmcU7ifSe1hrVOURJzyr
XlyZr/rQW/96nkamNdKMY9Wfn5K8QXrapKAu9J5KI7diBmq9Y+6giMDmeSC9W9NT
gVMtGWIHqRxN0gMJuGuBBOuT0c0aSSZ2rYeG4aSxh4NCXdBeJz9lTzhdCjCN6JJT
EmS+Dg2UrbxArZzRGm0s/V/Q2jIpsmiEO55KnTOMXeU023x4BFCa6O6AKVF4IZui
JYPF6929z8YzLUJIcA+cJsWejyozgfyKQb8j7443jn0uciDXMNE+ZVXIfS4qGPlf
udg53zS2ySWj8LUcgwTOcpCdBfsoGACRW4B/0/kTHg/L4/y1KXZ/5h7nbhE8aO3i
yhhUoBXvJhL2aP3SkcQuKHFP0ujuS7Ag9ajSwelqJY//pIuzIZz6DHK1v8Y4CxUV
ELARWujs7+VPXRq4MksYE9byzJGwoHkoFmZT+hdgCVLpOaRxH9d0+sX/K/PZ+Pk2
GEAmm0VCW82hzx/WetRCHXmGBwGqwkHMPZkm5UuCtuBfWTfg1xSl8miFU0GHtpsm
tAKUi1I1ukJr1gttgpMNYfrNMc8XIdoPfsj1/63eJBBauFeqFB/dYZmOQ3aHnzKM
tiJ4j8fWc64bNM+n/okWa22bsLTVmrjp6dzaZHI+rURanCTpuTgDeebg9AVjdZ7F
r1qYNi44/Sce/ovileZQXXa5UadLQImTQJ305tiKrmwYq86u37nR4kN1mT3uEDJC
a+AY8vaq+5Ohgq/CdysxO7TPfsq5BGOpT9NdQ8ukWk6dyQds/2vRQlNDKOBLHBcG
5S6etZEB+/mp3Fdl37W/TW0COq31UlFe/nlMSbnxEoGXWV2zlEHLs4JsRDMOvwR/
bjzlLvfoCyktVAUrdZepMK3r4aA/DwFvEcbJQtQTTtnNP07sUJEVXt+hvrB4a958
Sx73VNneLa0lDDL4rnJjeXZZZ6/KrbSU7inPHdMUM6HMEriMx60o/aZ8o6s+trRW
cgw2wUkUn12nzsvKG/U6pS/oFaJBsIZEGE01FxYxUKoS4QLHJJza7oPUCUDS71Cb
lq945PITrCXDl6IeD3HVpEAGe3Ez83/AAjQYhCX/SFCIwN5nJEIhnWkq86T4ecTm
wjEJZLhuzLgAfSCM7UFr/c2I11J8xqFb7iYAmjPDPp3fU41lhfgJC1DTFAwm3swZ
d5Ci8AMAVageZ8yNb4zvO9sELqYy7f4JZofaw9cIBAQ2WLoTHIiujOBvBnjfuzwI
MKYgaPHZjdou4jWznOaQD/icg7xh6N1SVffDKJmvnfvT5kl2hM7r6Q9sy7o0k/5k
A1I3CHvS8N5IDJnPpF+QQLwzU5Q3Hj+zO7V0NQLimduBAXTugbt/UhhzemWN0f1y
77BQmMNYYVjqwPSBgzRZXuPwigwO2js7IBriqJaKBDbWt42btmHDGJiLfA17m4je
oHknAGJPRp0b/nalMFuedjJaxz8k+Sk7Ne5IDdwPnKtLu0ml4V3awVl/j4k0l3PI
KXqTEAI2VoUm57bPSlkT/0SzCtARPuKDTSkeCtv92XuaXkq+yPyCvL67MFO93h9G
Ne6UFk5mr5hF0yDQZ7N3OPbhuh4qq+mnDmzMbwIehNlBaeCZOR5z1P+52JWK3Php
89l9ZXrUdUiBhZZBKDcalpPckvPukrYTLVTNdAnkKyhyvOZIjAPTf7ieS9+T1WiF
VM5QAntZVt4O6J2Qv5pM5fgqzIoxlhCdSAv4WesfWFqfu/sxRzF1jY4LGqqupoEW
+uCbKDSL9aDdvf4pIFbno+FA+7O9VivXaH7LUXC9ftZ9XmD55+q0JH6JkOIyiAeE
STAVI0CDmNSpHGXJCzXe6xedLq9z1wtL6TKDJ45irDmgoSc70T//vGh0EUDkov4x
o+/tSCroaTBpbK47e6sca51aaFnr8+t6whJ2NshEdrqTsLULAToHHyWlBmQTGZFK
R5ZFI3kH750gsd5Op2XMDm+qkAQ1fY9T+NYwC7PVTL3JLOfaQz1vvxO5LdJTLq1W
/xGSpdvxVUfGGqkLSMZj70XoxvMo3JhOCFcW9dOwISbwxrFBg55i2/mAuNnZvfhn
HIRiRZ0XOrVPCb87mVcdiU6U+44thFIfXkfKFz3OJh+j3z45N7CjhAQjoBR/LN1e
S4Dwbz60SWJi8zvAJYK7E4c2s5MJgFvkcv1CJDACWpitl68TL1aNqP7RVIg8pSHd
T+DM2J3bKVN7Ep+85kvkZknSIsG+qKG15uly/HFWqdzouavU4M9uLGPXz0TWmcQK
nKsI2H3EU4EwhCkJzHUNXYxGrhd8uriK1979VmZCibKKPiA0zUKh0x3lcxOzU06k
4aRCF6pcyBZr3deRlJOlNnCbgiG8AOE+RacBKpz16nf8xcPvnfiDkR1k6j7MmjAu
quhdwTRAnRklaXYK6a6AtJ1zjtw5s4tp6R/snSooeLn+MjSLww15EB0kM4b0UPB4
Ogel2gxElNQ7AQr/+bgEV+SQ52/9pmJpO59b+KNYW1AUrwd4/NyoE+mRZUdlhq4u
qoN4nlkJHbmLx04ix/7hpTGLutxML/N2Nfh2d1rq3mfQNWhRt7JnRLxH+OZ2cVuZ
k7sG4PcumuAVT9D+oBn4Ai2ZJOpvC89KDcxLg+PFOPgWLDZFvjsJGnhk4/zjWSu7
nYOc/MckCejA1ANOlPRm6UuT2iDwqcM0M/NMPswwsNiyjwXmqGYVBnSjLjHnACYQ
U4RVQ/J2cakWOUT8PqaJAVa3KgA3ah/JoRqQQRgEo/26Xem2hmoCdjd68rIIvxf0
AIYh9va6DCE4wSfIGSquQf/US2CwjI2NmSVXL3l3WvmmfoDnslzx2TukyHSRAq1N
cf5x+WiD+drBs7uNT7ASohcfUuwAirn7rmtnJKqg13bkprBd5HpEgMJYK5y5CLeL
Pe2u6H0mUdN2AW1psgMgomUAk4wwEzlqipHL36XI98E6xOA3e9KbwVWKoMPQn0mO
hH+YEsLByPDYxKeq7LUcMhiwtceIlYivTTxUPCqzRtLUhGYF6VFTnVLpZRSghA1D
R3TFjEblqnjVUMHD0idBizAR38u0OQs0PESzLI2EP2Gtm6aEzwvsdQC+7lxoj6RX
Z/H663H5qJGguCeTey/DCVXOTUnLEw/opdmKvq3utmZHwKzA4w11ofndDYjr34f3
QMBRaZoIm4fAhAqrRXA37JLy/JeX0AZxJ5uvXb92CT9YJrAM4dgL7sxfl311S3wL
5wrCg4ZxwwzUByf7eR8hy0T1rYl74kQiEv/OjVk5MM98YbEo85Zt66IP08+Ll09P
Zb/pK6yXCJj2NcIZYTK9Hj47yeP0d0WEUvw/4i5CoDQ3O0JLrdNIGyM3Qh7koHfF
mlFxqk1ARc/Uwnf1lw/dT16aAidW4NTRw0n8ZHIfH9BqcrI1YZ0PZ0dY09amDqxd
I6qlo1jrUrhYKReTD1wMROIz3lnFXlcTJ7bz35Z09wcODhIDnnV8mOZxa/cF9zl8
fkELa/+7orm4bGDHn94S6AH1oW+G/XctZauaHQyq6Gm8A1ULROuhTubqgEA6CN1n
fhYARzdLAxWRD+us8Ofqks4w2lYVhgfVI/KZ7/a1Rjf4tPlqsy/n+BB9//J20Vbg
Hx298V1yLQa9gWW0BEUq+7Xcewv+5fflvyhT6l/SC0Wb+pwpiiZgZP6Mi/Jg2QCV
tYWlFbi78X07csbZmSYsRXuDHKW3WU4p0eu8c3tz7Ycs17Dcvj7pyl5bMiJ83542
ETE5jCzXUdC4rwX3fQQkVlLu56Bgfnby1a0ghXJEUe8eIFgEgi5szqJqLA7cOSbi
DhlomjRTq8LlgQZLuySExNAHNHRqhIfeTD9cyjykmB6CAdnCDP25lXU3VYddL6Q5
b5/H8VOrm/+KIwx9Wnv4g5aON+eRx429/mzUxFUSow7UP8GfCBDR1VjH0nNO2enA
4H7XTeAwQc4KlXq30ywd7DNVAyLs0tL/cYjwzrVFAg/5isjXYlocsxnATReUuXFB
IXRD/bzRDnnLLgfyI3rHr7sTbx4Eargy8jr7ko8TLJuEQMUd3KM7Zd0MCflXYiqq
6vuSYtGbMq0o5J1roixkTQTu6KXmqbauMbPYBd23va7CHZIzn32wqRBCwJ/Hk52g
mfpSu+6UbknuWM1AqlQmpxMumlD/IfwLlMcLJzUVHL//AM1zYR0UZo8BCxveadGF
xO9gWXux6H0Kh70t9LRofbX71Rzvp/xaJwbui/oRpP/TMNp7tswcVyfMb1eIY5z6
oxVIN9LV/wiHc0pF4zhmM+OoR8OI3WGUY6d41TtqLmEh265A0j2oh3OBaBDcBXcV
5lFcAJ1mM4ZRK9/+GHBpQG1+6Tc5V3LPQUvJa49lwucji6/zb8neyo8lbHpjouC9
xTUMSatwv8Ih9tAJVYiwVTz1Y6H9FsOBz7220UXVez/aPdEaw61LEODpuKcUoWAN
jB4VoTAjT4GTeS7dWLx+V2IeC5Gb2AiwSAatw3J/qT6DPlYO44s/SE6KZ42UIPmi
GKLzggET8TC8ErPm+yKQdEtFDVkVPP1RIu3gDK+NWa7gRa/ljM+Ggvu/JJSy9Pj7
5jHFJDRsZlGF932o/EX+Qaw3x37dXHaUnZmR1wnY6GOZigk/TgUgGCLC+fDQ/HKH
llO5iV9fCep+KMAEF/9jauD0mK62DXXP7RGFH9wxeukxepUxrj7jgBrMpMh10KmG
FaixcCXaKuZ8yyA9n3RpATP1avJilubegY2Cy7OgcuBiMCsPZeZO0zQ+v0QyKEr1
8qRIyK2dc6iTBna5TblACwNyI5lUR3CTimJHLf5lbVI0LzRIDVYeaU5jyHRK3zOq
SRZSfL/Dx7bH2WfyjlLUiT60lOqM+m+zLUkzJYMUj/uAtY6j/ejkhCZmmk98q6Fp
htfjqTcm+I5EWP4My9F6B2gxUvydRTtZjPRpgbxPSmfMaolHbAm99V54k+EsEpih
LeVkBpkh9yFpFUH1eClsGIud7vmfpfHsAY2D27WmjqJ06PjQeoBmZMHitWcobLsi
gbOv3HClI6uKWbvzeorQzeeuvxXkAQsTkrSzZV+vBdgx0jQRmTzzmjfsaCt4FVgC
7RkDfCNv7i5CQ19TwA1xsxag59B0UUhwnyU36N9CiCi6jnHmWTpE3RKT+MLURhcJ
efeUBgQp6J2+yVjqTZp5xIEPuuaoP3mfL2GHw+az+hYbkTc744d+sdhJ+MNxhaOv
NijKSTREQZ6dsUgXVwgLiYjnXcuYBNiicauP2B5VcgPwgMd1o+k+xj1tTTqihCVR
r4Q69nM5qKiQmpqwT3IOi+CfhmfvvSfjKpYqbbxeMDR8XN+W6Zw8UI2tee5kN66w
84twfNkBhYEw1sde0r3YoArZHLtS3hMgg6/SImDjdcT7YsSB4vlBuaSBqXAgocR3
MXLXKqKrLlD5PyuXOOJrA5oV90jrTNU4RBRinSGKVWQoWD056Johppzu5OMTu5PY
1IFkubqUEt0vSwDpgBLgPTatQJSN8SIfGAejb+9DQnIek8ibdJJ57QejMB7nbsaD
TOeJraecdQ62Jq63wRfLVc8aUbl9qkY4ScQbSLP5j+TFahUgqRauqj9wbULoZ+BS
w2M0BIy5G6yhamW/a7zogPKi2HNfUO/eVfvPpZPwO7EW1ZOzzfLeoHbzeNSLWn+g
IGOBNimZOftoaptK8D6M1IVFvjcdZX/5Si3YEAusSurpCGeCI8WKZE7eqwHZFyPe
d85KGKksBNvsG2qgeGhMCbuEF8l1F0iK/90V6awwL2f16aDzPHeXMPOQk1fM4eA4
h3XR039q1iBDAonxrVCs356nt4H8YMXgInC3fCq3eErHAUsMnzoxzHxwAb2rDXgJ
3KvNTLdN6kavqoqOFxrSnNPp6H2zLSyl4KTC5FM92YmjD/E2v3NdvthIVlOq8NQZ
bhbLhkMkOAKCdsxxrvjl3/GWgsjsB+QOiSf0m6wV9ljJeMZYLqWzF5oDuj1FujvC
p6kcDwFGwGsK8hhhLhAL+6HdaWfGwV6rRVGmwj/pBHSXs4dXQsksq1y3EPeaz+Zn
YfyunDDIQKkbDh1WQNeJSYLU9M4hZmZzgd1GB1+RAGbXXAyJc0iyBu19JneXQi2n
ZxT/42+/diDXjePZ+8qhNkV18ADav7QL4LzFW8lWzels/q/yss0LtvZC3eaoYP7P
AkZbB8O7tFBZrj3eaYMRErK6U8D5MafI4ZLAf20VlX7FC1eiHu3BPd25UEJ7osST
oSgTxVWt6tiqS0H6ce9NW7odk33L214CX5/m4u6pl441G5Xi1k8/Y2Q6UPPIsxTu
Pc6IiNrccqDz3DvlAnz91U+nJn851yvsXwidQfZABZ8tfLCsBhnaKJn7bxdY0ljl
9Ns6I3iKHejWcClnQHApSrj6HDQ/ldTPFfkYLGS68wYUac+KNvEeEGfYPHfIsgSm
b6XYYj2CEIrNgIrUkwcHkdIiLy0VQLGyAFmTO3P98BgJ4w4B5s83ygb5gWcCfbdY
TECtq60WFZPKUOhMc5FhSG0I1XzSPW03ixnkQvJfDL1Xqw75wmuNidGzy+MDYU/n
gAKxmu38/gizyFqlquVpdGXbU7AY9QgOlx0D+5c+qEpP7olcOc80HhUb1hOtsL6o
Vhk6P9u0/kLJc5vQMePOF9xb+bB9HE391hPb81Jg6iGyBntoR4Ki2NgWyGuZP2Xn
7rve6EYe7MfcZWffa1CBLSEDwXQiJQbfd5Gu5Vf96JfOlI9tafmAeBHtuNo0Zsgv
hZoDiuOhDn8HKCM0vRLbUMmYDHe7w6gkWFS9fJI7Z5g8tfhQsYeEA6DeREyPKgp3
ox5JVqyHTaRhB3bb1XzRjyrrAWyOGIt9IM9v97+OI1krBqLCgkqkXUPdeaRCFbfu
RpOVQ1TOvbllpaTD691N/cgty0sRD1zjwQJX0tTv7RLGn3vDMXnC2G+yv98/8w0f
D3b6U8LeMcfMYLXWGO2/LmwehXfn5wP+8oTRHsoYNRqAdPZr7aGyrvIoEoOuPQV0
mCMZT4dWgAxNMwAl2MYaLRTBGpEYeitoxVa2RMxy5cgKvg2rOBOkV+fJFLkY37zS
bqeLQTHP0F0K9lRmEto+PdPPjSxfflZPx+ZrGRhOc4QtuCtCz6La3v0CKtCPYXdY
Tfs+gYODNuCFCN6es/hntvtVOa/TjPuZ/KDOzZqI97kISrMO9NPzpHldj5hc72g8
5bAmvfgvQcmuznvgYHSdosUzovKyLorB8Ouwsh5KfJBPsijZou2osHn621lg2YiL
1EKMMSAZ92SlpKv9SZ9WGWRo6FmxY+DpU4aYkAetx+cmPygFkI0KAZFw26CnIjzB
tnqJn4cn60EPSqK9DL8zxaG3hfP70fHaHZm3ENbmmiouqswfxgIp9CrI2IdTBfVR
JJLEfb8T2FLaX9LoJq1l5katt/jQyZsR1zvc012wbgoUXJ4eKSO/X8oGBYADHVgy
CiG/vgvxadOHCaMhnxPigvHmNMvrekUAaqFd/sKKO8/fPqEQywsY9oNh8HYcrfjX
/zoW2n1ve7CUS+L8mXp8A9s5i9/EPwa5/fbPYcfspvusA1SPiVpuL7hcpYfQHE4O
C/CBnBFtt6LeLG3/+sXhHXTDcPN8UaO3/Ni0cjVpDjofiO9svD3y1Zn8A+rIYQOV
uWAmYGaNHvaCr6YKubNNkTmoiP/vgGJDwLUK5KQs81q456FqRlIZTR78doWt/4da
ECmmGuW5ovihnLPQ97QVkvNIYe4DUgtSNBj+HzHKxCSMrJabooVD5LUrZzS+QzB7
Rd5A9KY76z00FmeeDTpuqd4yx6b6yLyNh/KoZQ2MU6VDdW6FnlHGPaJsUrCIB9vW
t/hNVn4JdllAynZPAcbkT4bROBbTpIJfafH8f/q2zMSkVuQaZdzIGM1RTio93ir1
ptVo+/XgYTHFw7vfIzsQFLo7D8JuvnMTkou+rwWlnI6LFQiBURsN0nXYRnYC6BBa
2YG5YlFIgxIV5swnp/4OikAkG4HnXLgwPfPLOKB0BxHx5jyE5uZLTw4i9iZ5c7eD
35TsEWP0CfEHlj5usf085ni4BEDyOUpUwxY8spzDXoO4DQrWIR4ASZUAB95K6sKJ
5rbZFcem/W1QR9wCmZlBDH2mlR/PMyhrUemA23QNALHTvNV/CDluuBXPOkHSHIF7
ciLmd3tymHKARcxblQIarCLUfu21pTlW22dI7wusVi3EqYegHd70l3BYSfmjoOmW
Y++YKSIgtYfH6swznd1AP6+FrzUiVlLJr6B0oZhLLnAtDMEieHiOtVnmHAP+vZju
jVVTfzWjbY5koiG+JmJa3jH0ifMZgWig93FXVetDBGzLXXZmSKMBkLXnlVDrOIIi
VTeNWv0f1RwImX09yhuWDlCYqTS4StixNNNBiILgvyFYHzzMHq8koHcbCn7lon0k
5lVjzkUq/1swdV/WAqykBHjaRgXpb46DsGrLtfC04x0spudKzFRuZl5NztXmitAL
ts6MKNnHnJD5W5xHfH1DgSU1xAAiS4JXtaeVhFZgrcF23D/bO0dhsyAAOSHtmuV1
wmUP7IMWhF2eNA5BC3kIpOF7v4qPZupcTBMhc55LUmLTO2Kid98VAmh6HYErGM0P
zqng3ly19krjVBdia0iBAOThVdYBL4e6XeKxKMV8RQiNopghTcpMRch1w+4ufQil
TeUR+pacik+i3G1SgKQW6uJHEWBO2mvgbEwKYbpqFaFQznCwZYmgP0AuxUMcXKnl
ZcgESZGQQatcDLvrEC3I8rpY82VxkfOICf8rbdU/4F4TunTSIc56lxmfBxUpiIMf
bdbjv56nmsjIcUNuHuTgNgZn7JJTjTZa8V8Fjqaz0VYRevPixEzhoBwBqGrfzABm
WeJNdILwxX+gJiSM/7u9mRo4rHm4VuWNMpaYdI9WLXunOzEFJc8mVDah206mROeC
Q1H68425YKW88h0TO/mSi31oDYo2fYKQcNP8UoBb6F/KOzHNV25GYIY4NE2VuDQu
+3drzh81Gn/QNxn/26u30932f1RFC37n2IPYh5F0Kt8HQHojtYE1OYyLsE4cEz/E
h+ZGcrsGDQ6+gXGHcCaqTnTOmdnV6IgNj9oVUvELao65na/TGz4TYk6VV/cNdRaP
bTaU4AQ5omEytOQVtzQuzJFtLcxOfH14r/2JkWwGgnNGbV1VhdvG/054+hGKl6sy
25ruxN1wrV84uI8SzlaAwmp4B1IhGVNghcl74nsel8bmLc+56iu50YHGp8khRq+8
nqjF3lfozCovhUDtfL6DxSFv707b2nfhC8kAz9p9Hd1w/GtM0pxmMCHMuyLjz+WE
Qdcg3mQPsV7tB4bvTFYUiIreF+6Oj9yLMA/jLTktD9LqaguLul9zHejuaIRQGtxs
lw3+KJkrpYJAcWuTtNSRla1dGept4AsHJ67oaS5etWfUFe15yqBw3PVq4WkZFBCK
ZewPAbGXiHrOVZlJtII07cc0qKgmXEcHL4AFqd8SgN23VZbPhyWrWJtTrb8UOhVe
t+Yy+AOLT9DcEg/DwRWzhj1hstLe2qhs1Kd4l8i+K7O8kpyo6gpraO2At13ZchP3
SHGTeSnTqjJL7gWb0jcRspcXYxEI5rA+/2j/jH/vv9m2SDqVJgBzCTcsdoh/mfjz
zWxwQJaqdOx3xbmNueBxFxMUwbF+e2EIRQIFrPkQ4jQcwcNiG1uRpsi8DOJQCc5n
UHZ7IBEKpHTyRzmt+s77yh/kNYWI1yl7Q9mwQN1ccVJw38DWCB6GM6fO9Bv8IIu8
Cgn5tInnl1g67WYPCHpM5KdPFDNRe6+T1Ra9JRFIEoXtTViEpuSVRqP981sr5UoN
63OUnpbqNcW7Oiu9cPI0yKnHwLtto04PN6Ti9qYVKS8huCwrrHxLPztmKTMM45NT
6XR86E67nvrYNrlXEGvokMp4vlpJGn/86fqtn/PWg33+5QW//guDuBusAlBvoJvp
0CgYreajjwM8wlDQvobvMnzZdIKXSkmq9aQBP0sWkdNmZJRJYdLaYno2Q/Pdm7ss
qXJ2K7fExpH4JTZZKb1DROqkgIKANI/os1bo9qiR15xCEYAglbekJptJb9gQlZPO
pP5mi0PkZLxiS2b4bUQiSucDwg8f9+nOYTQfpzPQJSOotRLs4ogP22mRwN2Iiict
25A5hYb+rTmE18zABMcVBNUATdXH/4vuUMmeUVi2nKCVb6bKzwy2KyAc4kcBcxDW
pEKU4sJwQNHtIBZcVunNfVVIOpkFLmb5A76A1BDOcPVaiB7a5HVQTcgiVxDPpazS
emJg5Qk030QjlUbcPZ9YQv2bvKKhOLKMcf2gejbwgyW6gjUo7DyZrTTL/xfW1GjC
FAyoiItCQK2ABG0E1l2JEslw+ThrspNbFLwd8A79djtXtF+KW7L/SWhtgwZeXxm2
yM6GS6RfOpIEeoXeGSjDzw3BZbYOgEh0eGlp0L63EzTN1Wsqzfg6QYVOp4USTNzB
XKHKNjsIoT4R3mNbYbIY2/W2drxI1GFnuYpHhYBvvXJfm+0SMK4GkFh/U1fzIq1N
vdntotqMv+eT5qVmm4tLaOFehKaD3njrU3OrUooSF1cJeXQB+zX1zhLgsDJjx33n
U+TlHAasD2sj7vgUhNxVMVYcweVq4XhHucS3widEfNl5EVdb64Rc/xFVn8HgMTSZ
q1hIwnuvnrayPxNEulzgl2p7SSfubq4ljKiyObTBlv7mAef51oYsVsj70JgwmSkO
f7dmiZtoUKs0JfVJT0aK1Cy31ewhrVea+Ywk/0zUNXblga6w3o9vSwjZhzTsXdtk
GJ3azCEUq1+LDpYsdwd9b42STXmCukGh8O3I9bHXEO8DmNVhVYFxnTd2B1BcPge1
GZBxSqs6CRmWVkV40YM5lqj39n6D6UQCo4DO7urCq0qKtTUZGq5p0150iwgjZo+U
Md4EcZypgBIhZv29tcfQAZF5Z4P43/IJ4189zqKtgOhuwqK8ss9NchidxlCKi5kS
SfZAyxXlC5k1GubGAQYkl9CxHAaZTnlOwxNARGM8BBi07++9wTwSwr6wIt2wuI0t
HnaTE2h7QLxcI8CzZDnayUnp19EVq0HnE/Vny0hFLJ3G2OWOklTDT0BhDTl32Owg
yVvoU4BlvfhkXsSNcijTykkrS44jDf0fqKzT2y+KNxnB+oDCtWvmYM/z3QnPU9Th
SSUL8wm8lQ+odok9V41cCUM6p0KRHRJOxzFk5i2WjTcuu/VxZssMsu05D1BbDMzV
F/u/a7OEpC0ADjvqcGPVTQuWAtHFbmjL6zubQBtVhUVpvviLjkqaZ06lSVe+PVmP
hdi/oWB1WBvIHBJN0a91R+V4uEZctIlIudg+eb1JQoYNaEsS4Cjj5PxBBotvbbmp
e3qms86R1xGkIijSJsmoHj5za6DKSVBQrl5Bz0LhdNm9lAcwJ3h3/0Cu9KuVpdXS
81RmNOOIT3rCtlbbW+aoXpKLhoos6FADtOtjeubOiCmyQvDeTu8Z4MdzS99awXjr
aG0pL52Bc3HoSXNkZZPOMLRJonxedQa0nYL3etztunuW0w6EWAhceVLW1d0FSWbj
2RtWg9Qx8l77o6dPLmuH4BVsl563NrjYn/7xsRlPCDKt8s0yOnYFzVnRLNWwT3Jf
K6zu1+X4qlfs3ZmHXDMvV+FvXSniHaJkSH8SUrqcSv5bm+Rt/6dqm3jrtn8ADS6G
NNO8r8l4eqnoy6nnpWfjFhEJF8dMBIUg/v4a4YI7cyPHRpzSHZoxtX/qoE1+T3DL
t0H75VPWxcAz2dhnpCMwnmcCt2QzArfd4cN81MTCcA11tJuc4fwKBBtf+91y5xp8
mrhzcI0KOhN/1eJpP6/eFvcjAGF69oXw5bybOavNdBWVbrLDlhgGvijqjDiDuvw5
6EdPCDKTMZB371YO/pyfb0cS1aVEJI6OLBzWw4EL22oGXZe9zQLQ0n2PhBK7WaNA
8kETFUp+mb0sQzn5tQXaYsX7hBndoYhELQ8+/Ci8UIOKjVg2qOV6MahfgUHyVWhu
xDf9NY7k74KPt60WJFcAaOOt7/iF5f4y/4DLF1BnqU5/hs8ocKeo7x1AjU1O2mDn
2sqwGagftrK4rlxd9gWDblE5iI8z6IxiJyfmskW8D9d2JEiUCBCbu8Tthu0k3l3a
U0D4zXtf2T+n0lkRjLhQCMQLXcnDFERUWdQt8dZPmIbpLO6b8DcOl7/GXuP2WHif
m43oWfHlBexzwuZHjEwLEOgdaet/iB6oYTJAeTdMDSh40s4Aw1xiR/i3z6zkEgAv
kduFLRcP7bsi6YSC/0ylPFfpurPHRFb+qmpmsTcXzu5Tle4ufZcXWE/gRq6JABwh
wW2GJLfn5Osd/2B6s9oqpFqK0i4PdMT77WzUxwSYaq2ErEfubMVS2h1e8C3rbBbT
N5UKjF1IMUoPGVdUf6/Msd+Ek/MiwdTpOCYqV75u1DbFtcJnrWJIiR0cfbCjLOJA
mYqfjEQthpTolXKF8zg/QOANUNAcGQRnH2scxAr1zZITRWBgiwgz8/hRC/qI3lPe
BoE06GPyFrGHtaCWoLV8c+NEmJJW7Di1ePijhPIFC+AxNepkCvjn1SIdiYuhy+qU
Du/KEvibg+gkLSnmhveoqFr4zpvkKndQ/ME82cgWU7EFGsAF9fj76Nl/5OEPWywn
bQr4eIHh0GXagvhYBvlDEJQMCy3pzIpHUEcIlTu+8Ni+RIK1XjrrbEFDsPnx2heL
57bIvlrz0L0hZfCNfbqrvBKO0sVszsPkf/JpYTZ6IYb5VnICxTVTOduvqMoeC12S
/VXg60cEEJpw5tdO7wiQFFQ8Z1m2xyt5KpHrWajWKG29LqrttEnVuedQ6uAzLPN4
EHuXVmUuitg7zlSEAgr4k+cp0gyiUqZOTpEnjolpDT02ByxWIx3yNN5iT8H5EPTj
QVEFKZA61ZYgZyE81yaDvKhca9+sCdLXNOTnflunoxOr8Jc9mzOmw4yAalco+foI
xvrtirDWs5DRDTLhgig3qXLNMGy8nAamya6/kxOAyyZffzAf2h9WA5JY4fAZQVJ4
YVX53Q7ZlSixZGrla9EV6Bb8WXUmzCAVeYVuUd2HHbE24OER/YcOZbvlAK2peK5c
yFwZe1boCYrcVYUEA5pN14xq+TBKXXHmXR+OrvSHssJ8u7dgUMDGEBKg3Hlmb8dm
1LIExjQBL9A8gejkyXLLP7H1rJKvpi7pa1/MTLuEqCwTjxa0lya4AToVmzfGNbuW
OaFdu7sCZSxQSHHS5o/NSUz9ebKD8GVUwDO+2qfi2eGWZSf+p1t5hWue47ksuXsq
bBuC/XLTrizN7GX/64CN3yNtelG0Pw6lw6MZ9HRd3iKi3WMud3H9nooLK+DlSfCw
chp9apkv296v2MsypbHAAJvUc8iKD5R8EScG+Oa8KEZk2rmJlbun/619XL5+4a9G
TFTlRV6/fRYdKH7yCICDg+LGJr3St4LkdX7sHubpf5XCY4dPol3WKIakX4ugOz+u
CwDuAQnwEOoMnMOZ8xVcP0QELzDzyWIYBjaY33E4T97aOlL+NvRRBxIrbufHQAEx
6OGEcOwjjHKDln1WpIRBYXYRZbNuh036ArL24xskaFfDIK2iRhdWRsC4LqUt1uNn
py2oVyZh74i/wFRtLFgpQ9ZTXzGHcxIaNup4JmPEVjJpgjfJ+XYNY4o0+urJJGFH
Swf7f83UMxq1U4gg8Lc+pi+++U4KiN3Yia3qnJ/TyuyoTUmC3MOAQF06dR18SCGb
JNnwOzW8Z+FRCX0DsHkSVfUZZ0HQ0pKnKFL5cJJBoTWV+a0ZcqKgKO5ORYxc1lT4
n6DsMhrR+DySu5e4P8NJCVI7efo+RJW6dDXSMq/xFGNUmmt/WFPXq4ozBIDMaio3
X5vp8FKsNwf441kbQ882jO7mSQCQSyML3ZyXbosuDxSKjUXxDUstaF9bB+C4hAKM
ZoO7a9UmiJFlTPV0MZuhHa/8mWfm6KrvoBm4kA+WF4SMe3vaRd6QvynkD0+kkecz
S50eYuRZYQQH4y+iAJAxSUt56eyY1fHzfhhWUplLpYSvfIsGvrgRxKK+8502BWFP
NhYaxWldLUywYGabKmAuCq/e2qFzja5sp6gkvvs/B7pT6vJiBT4jDhN87QgSCOAZ
3jBhknaQ4cyHywOK8jqGxK1tN4PrjQMK5X2CzVY9u4VqUaJ0a3FIjZqlsczW/CPH
rocR6NgAn1wazBBoSSOgZ9DfdL+D4NU4O7R4rN4hq+EjBvtS3uZOfOTkyJ1jBWYD
faLNS5TCfJl1V1AvWjlfQKHtvbrglvEcZxIf4mFVxbkqd+F/BSYxF3PeD3KEXD2g
x/pu6Wn0Ij97VU0PMaUZwXdBBfufodagFf3eENuZUIsqd6EL0LmX6HgdMULfKHwy
yUgaFlFoY/28t/dWV+YJTPru8KMyc1WKnl0/GENx6eaRAWM6RoKJiIDhvdkXOj3E
ZMerWpy77PI5JXxVD9TSmd0hVgtSdRv8xyvUYULho5t7VZBQyqC020NmrywWYSoM
BPAy9/60RC7vT2Wb5wnKq4epFxmBl53gasdBLQOjNmU0kjbbeXXDi5AJh8iP29BV
VkWCfwYPNYCKy9rlOZ7WrODJ4cFercxvb0+o8wBMgrmMlXgLv/B2IueA54wNUv5O
8oA4CZkO7X/jucZMSnpacRjErIEBp55TXwGmTNHQyxWEWAZoKEoLrk3Vx0puHY0Y
Vp7G7+Gag0t85L6L+PLA/gPV9uB2U2fw2JFguTTGOB+zZlD7a4meVj7Aedcx5KHF
YC3/PD5WglwSPV4uCvwnQYaL8qBWGIEU3d1YCXekFfM/9+rIYcv6ihmQzsy3Ffpp
f+gAfMZksyqzJEITeJRNmAQUM/tTyqtZZdY8GWeZTNTfmI7bZvtd3CPrnTW2CTuZ
COtqtZisnLkiNA3yPsUUB4VQKqDOGovocdBt7QJ8U4I0JOCYwmIVFiWTyJitk/tn
D9Tblp9hExkg60ECwxX5FfsU+3Yf++r99LcX7TSn8wDnaPEPnjBrzcXCb416BRWY
NdEzNiOrSID1/8kYNQVuuqOSlSb9gDEhUaXrTTsRaXSAwqjrwGNsMmiBltnhUFH7
fiLCuNH+jmeCNwJL9Gw5sWHMDZCNtmThVyibV4hfmk4hSTCvpMiwivh8qyRktZvj
JOh+v800w63aSG5r0wUqNC4WCU+wxDweHzTLne4BgUK01YbrfrqXRavr8dMXvl4o
bT0TNyW7OoCdGXP0hbnIIyYL36TbiAVECAoj5PB//voD3G1F1wu6J+qKLOtlMRJu
Ff2cHJM8bkDy1MJB81q3qHZaHImJDkLONFb6pjpFtjf3VzYpNKkGIxR5WZQN/Flk
gKq9IWEdMk7mGuF2EvftCFHHpBhjIcxOheXka5CWSxieyt4+hWwN5stp1AnFLz8N
rb1xOGsK4iRyfH3OUYNBkL2sfVUfvwbzhCnVVSXxNmmEhaW6hx6UNUjYBbGWt3ny
wXX04WPTvsRMUfF0kCs6El8R9X1JKC+S8C/mUa6nRMJ1Qu2RLVuvAPe+oc1dBDFI
vaM1uq389/xDUcdAYWkYbYMdhVI15pP4wWergrqbwcjboux8eLGPca/bSlb6MX0W
9+N9u+ovGpCGyNX1ugkfIG+FXUSPeUPx6CXIJaP2LIwTi+yAEwCPvtlVYnbmNhlK
YvfQ3cvKZgVC2yhiqTJ+UD2eHm7PrgbIEkFBvryPXPh+l52auSnX+atRbLjgVwHG
s5k1imJFIrpZ6yan0YnTil7Dk6i5SNFu58aIEyzfbGpwYXAk7feEQic17TmZWK+i
9ZkOZLELWdu0lGZkzNVWwqVityxWpmQSIXNdDg6JSPiEjcHBppnTLmV3bOXczgqM
iXhRE4juQnho8QzA7hWWDd2l+i2i4mr2L8QRAjSt4H58DEShAhRtNfS+dboMpkDc
mkbivtbot9ZClxad8nGdrZRjFxDauulRvUO1CSqkHgzzAX6+XRHVtQSj75t8leDV
EnPURia02dlc0/wmvJAm0Tsk1zR8UbMB5UDu11BEdIoFweK9+PI2b3kY2GjKbdON
YKsR8ZFuWkBHKQMmJWJ7sF38+a8GHFmSrqeNhveCIIOnQy873dVmNYIokhy34Dvg
1msVtK8ofotB9+GCrFsbE2n16fJCBL9qzsGwZsE/I0ovSOxG/BWYb1yFKclOVAwl
u0wvOv1Q4CixrQAoYC/Fo6XjQFMhf8JVvXOyB38LaImQNrNR1BD7fLua/cN4RFHY
gST7eY+2gg1Ua/zYYCaKiQrDQ/q9+w5vy6elIxYYCEIcRoFU0KHsRgEJvKRi/cg5
qDvXgj4QkVx+NjKLmtwkEa3fFEGeRSjkfCgD+vjs0ZQ+D+cTzfS3kN6CuOO0QQOo
8FJsDZEt/HMrT1h4xlpJQgdjiJZL/EuD+V1oGqCmGMak30kN84726zLzgxE79vK/
3gra52Zp5nuED3ybj8Ug6k9zyYtx38VRZimZ7FppTjqOmHMCIIMeeZfh6chhBssS
M+mskhHurINN6K/CH7bsbgqv4HQAar6PqA6J4eg8uiDDbmZpcH4nxsxmVtIVrSss
o2I+fpdwGYjA8v0TvH/3anjsTAOpKFvKzIx92Cl5l21qRXh5wHCRdPVD9o42bsD5
aN9zrEJXgeh8IBSqTuX5Dk7iYB7LRXBeKlNQMI2+XmEw4NtXF9r+/6UuTVjAtWzt
eU8h7dpghXo85JOjqH2UnZqlYBqcg9R09mC+DlTR6oHCG5/kL3ydLnPU4jSyzyM5
/wZRAQ5T68koXmRv73esQr0Cc737CGAXATqiYIzAlyLVxRS0mk/l1aM9rwLP4nm+
u3hLI2mhunPE1irPGTbj6IElTFjUE3290uYkrcnh2ocDOoWN5k30rJ1GU8JGkHnS
y6/PSBrHJxYvyFoGf2ONED875N8iJaJxyI10avxUls68/W1/OsjK+5hm7VeOr5I4
nfWOyWw1N3AqRS7yBIdPQqXHQG5DnzQ75cdifwWOomxMMKGnyZWxz/yTrgUdZBFO
+bt1j9UbpL2JmWqkvUwTFOqQnr1uOTaHl5DkYoIS9rE6kXwODHx0G3RgjUdgjqEU
S16AnizcsQ81kuR35EVxDHdoQfhbOayj/PCprUHJYaEOZOjuzo4UI9WItzZl/vUt
MTtgF4mnOw+FKFWSYb1Ee8gXFBDRDsuWAWNnwVZR8V4IEQfYVA54LoaklGYEa+EO
8pQghApkkC19UDXtyL3sCVAWBkinWNLineKFPBdHLlQcft5ievlDxPxVAQDfUEvv
XEzEc/O0F+IDmzxkz+yTeBdEC68YEBhAqf4Z/RVL4i35YLIKR85rIRAN9UHRSsjX
FpshNNvveBtSPf0Nttg4ltMPKj/RB3bh4wbTgrjAvONe6DksoYJN7jNbI/GL7Pke
7deEMliCzXVtqNPvRARAuyt9IvET8f60k+nAoxyjMrgD9PDavkQhPLlLpNoHv2Gv
PXS5HHNclAKoKbssmfPLzWCMeeCWFmRIMuvsJes3s4df+ghLY2YAarH0iXwLafk1
Ou5d0WSgD3RFGuLKENV6YCXSiAbRAdsUaXYA9KSIElPb4iX7XJGs40Hi0AmcRZPr
mIEEb4m0zEJDYXAhhOgG91NuEZPC1aZII6ZoOPn/N8BY/vdHvDbOd+4GKvYVgxU4
SU6dqVrKDb1X8e/q/f8sZ8cUiOUyjxAe34EvCGq0niuBxqpBorrC4e1g3RMoldXU
k3yXueu8Ut667mwMI8SWwkDtBC5mxu7UEqhLTUPhj1mDka9+0C6czGwWE/0UpzHi
yVaGR7qkI3PtScIqtMs7JwEkLjoQPTS8BR2ZIktDHbZMirNQyVYLRBpVN+gJaukN
RowZyeX+7wd3w7dNfHVqX/QHVRXlygcC/IEaFONV5I4io/UyV+/V7vcUPGBT1cAV
feAnIq22JDEfRN/muyLjMSE1ktZZZ8H65qpaDzVb1PcjR2RMXPE3b2tc3dAyEwfV
15OKFkSgQ6jYUHJoLg3EVcvUcicH7cYgUc/zCQSePZ5JyQvCxbf8LN1Yt/Zedo9M
SZPo3/M8ZWlKbqMQPDT8s0iQmrBILmTVytGX766uAyocdRnCz0Vf8GRxa3pW+xBl
IvnrWm9p/Idq2HnheSzS6NryxqX5NJQH6/GcDr1WA7KW7DDPlqTdm7RSu4iRa1vU
4s1Y/ISgXOhcn3p0yylP+JM0zImp3zcF55c6jF1Ma6DVGzKS2gOaCySShG5fMmKJ
7VckvwAW2O5rg9m7JKKFI9YVsJ1X9Cg+9+DLA5qO3X//beou0OSf3BHcN4O3tTB0
PwljLlhTj46p1UrMMq47G85bkzZyjUh9Nfo7WY1LVUXgZKj1wJ4phvF+RjvnFIEC
jfvHOAhilOCaG/4OL8zXXq9WCnEl57ZT5FHzl3mBweal+xKXJmPMybc9Q0cAcQhW
G7ahfrZJupYI3ugU3chhjAQgM/sRkkNONgDVDKg7xbE184605hGcEaHuphyTijdH
/De26wdMPSNR5UKHJujzNQb2B4HUtFYJ2yAGmV48CtAM36sG9PhGuwz+KaOHqX0l
NlJ04vLlZcqovlwKtH0fJznN+7ZpKcC5tgnm07C9akOfeBamMP+lg8IrcNRhu+cW
ZXfaiUo/36muDQ9rQNC2qWRsUuCqw2Kr6vDnpiI990T8MNyFYiS7SY5/cYyJirpJ
qXBV8FzmI43F+1wjZ+Gtz21fJuHH9FNy0g/NG9/iqt5T2Cz+2SoA6wk38F0tTi+b
2efe4U3Lcjh7nJQnoAszixzQNk1xm1ZXoWjar4ZCtE4SoTrGGY6UdQL+WpkaSCnr
BoTfoe/ZGZt9rCiILc07YIQgPxuHC6yWtb3BtX/h02vhBtXV8sHcGQZfNDCUs2ir
SksZA67oZrxHSYMGSR93q6HxkajZQ89GhMxIPMbFytXJ9MORgnBU33WH9EO2DduW
rjxQt16cPSdFCdI/dRUuxrug3PBDGOTFyznwq2Pyk733OnhchZBQ4hAYftV/b3l7
GKY05ivGL0AQnEfmP3H+WbX1sVsF+1vTgx2mlWMmJAvSIUuLR3f+/pLun9ii6dIx
fmU1/y5yXKiEG/5N+WpYASpVOif7ife7blnK38nRn6Ap2Rxqoxgr9K9t0UGeOCNb
N34sMs4irj6doG6eDKWxQzIihqxvjm9OGwbx98hnu8FL9iMbAPnyCPhDjs45hL1F
r8h33dF7NjCd8HrgUt3snCzYcNt5au6hvX7Auy23Bp7E0wF7J7lPvbuTLDmMzODJ
bFd+GtAt/EpOxXU3IFN5N+HD7ERWYyolvuxNswQ+g+5hI64Bgrio9qWykFS1Uwyj
9GUjZdqAuPLlhFy/16usDJ6ER3GB0PlLs4qH8l10ClruUtYYtiKT/7hE7puGPm+Z
C2WDnsNmxnstpEWiz+l0prTmv1N5x89yrJaoIh1j77GvwkI9cdCo+ZYby7XgKxtG
jMaxnCn1O0EOMMIR2RrUWrutmrh2HEeM9OUCfqjPErUMURwIOjyO7o4wSdkF5VZH
TLQsYedAIqpc3ByR2NOllwX9JMSOHQHnvGIDvVd7zXJ7V43xMg0P6/3jiDFnRaTx
MHIq0k9IQ/gRWOd8qtKaihFNtvXm9OjegRvowQUfT5T7kQHGRyOMk97/GRYDpeep
i0cTOxUeQM8hsql9Jz28GN4Rcewmyykc5CKO8yHV6XXYD4zrH5mxS0w+3f1myqxq
zlzMJyZUfNDgKCeI/AlvU1rx1cAnH+ag2ZyFuVJjglq2hQ2GTAKB42fQQ6g58ImR
argaOkut9JqPewthhuf2L6F/MNCXC6P2NNeWOJeyFG/B2/00sSYj3lFVpzIskoTA
ZejyHB/JJfV5Q3acKlQuT+GnxswdFChCHgwsl/8ppRYZVstD8HZKzqxk679en4X1
uZwvYPTPagt+lrTY0IoN1kTz2bHMh83iWLxBtjjDThk0P+C2Rs8iB5lux+dccHA7
+vx7VtyYH+TF89nSNvsYXIjYYo3yb17vkzqxLzNzTcfNoMLXNZWiVLlCYx3UNKgT
324HVPLgKenlVCMYrd9KCFWgH/QG1RLWLloUSip/i8dA88BvC5Hyuk1D1TZyAlqJ
rs4paYAzlYPZCYwN3x3qP3wp89d1wtqQi0RSuNoSFZ/99ymIkqYoC+yNutVdKfja
wewxt3NgEJbs8KzXbQixFgocGVnQ+kt8wOfmf4aRnpQBSAKW5UuEjRqU1zeh5XTa
0lFXIA2DLyAbBZyZpgztcZGE2EDK7N1xBIbkYcGMPmgEkS4mHX6m5IKABVEe+H9Y
xycnJ3B2yerIUf+ehdtstEEMh34rmVge0RRY0lXeis47joxhzutHmh1RsRmvn2c0
Tr091FkndcX9/CLssWD1zMcqVP5aKkan6lGCE6xyyxDw1aXJDM3XjzWDxSzEMKq0
7BbIevmjblvv1Vd7VYscCUV9G+IO9VIv/HreYmHaPFKnzgsgiXXS3EBbtlI63lyM
TZd0Ugl17V4jmBVqb5GyTI9u6u9Q07R0kXv/0sETVHmtvCp9SUdkgUX00jgjyINb
oWIJViy7NVVoQQ2GAAJGOUSCCCJHSkLOSo2Reyqbh5dxWV7QrbwoJZjBKuZ/tv3j
F75MZfuq6UAjuXxGt67TKuATWPQna90zUrrIjfB2EwxmWB8A09yHxZHk+kkas01P
qpdSNdioqbuHDQrqN3JvtIDRKL0YGjlT64m+CRtuWJ830zetT6zfpPAnS609Yonn
E7eTvjy6uUIQlOO0PMvpxHwIufpIsIrBNN78IteB60X1GzF7KoqVhppseQ2QunEz
rxQv7chgtPRtp160pWdAcaiCJdX2dhsaJ1QRtg1bq8PAJwP/H5+eHyC6Ez0jysb+
nEK+KbtaXki0Yamw4s7xiXTnQc33eO5dB/Kt4s90+fEZ5Uvac70yZ7tc/iBh/Cjb
Zb4z/Ek8qTRrhhIRV6fTsLrOywkxHha8TdfLX1Ngf8ck4c62dwhetuRhc9qFQ+7J
B4Regmg6u6O23rSMboyBpyzB1loclTeh/GyDyYKOHNqH/55Ubzg6s5KEYwO95wLx
QyxRyRvHLNbVzghcynrDRazWBoXRjLLBRICOMz/m8Z8V54toRCQf2zDATWmZEvI7
clc4bTuvk8fmhYTaD2X6KxvhuEWyh1F6Lkrb9EB8fmwJNOyV38Hw2eBCb+zt//l6
te8IE8eyjgxONHw3qd54aAPmzFgrSKc3wrZnYaBQ4+lBCtOoPKq8LPJAFmvbLTlp
phl/sigBIxxAO+hSB9QRIuPHjZ40+ocg+OH1P8zVa9uVAcHmZD+2IrQzhZn9oky+
ROHzKYvEt383ESMo+0eOjkjcufKUQc9PIqGMZnrJ4bM37idqqNCqsLkDkaZFCgP+
pmFMZ5f04H1rOez6LdJDzaVFXBHYcdcuYCUYXNeBMJm9ZF1TlKYMd+Lue9gX2aQl
0Z2x6ad6Ay62y2kz4YgG37A0PWHOirPyA5sDkRR1dJh3MHipbko7faWgiryJ4Mf3
PsCiW9lUAA6K1Tysv+3/XeP4AShML7N/zddgqNoISBVW1ki4MBD7XQppEWweJi2+
attC10woWn/K+PIfLboiA0RHq+3082GtjB1Pz7rJn6hN5L0EpU5mEBCbsIrWnHML
Z05gACyPx3hj/6/FCXd+MSkI4ChDGWZbCokFRtuUEWcE1V2vW17kzRD8bNFmiL5Q
XtiRCVGC3Ulwafu2I3rLQzHLsda5gTgWksyBSRcFNuznnlWTenwrdx/CbhIdeaY7
VoXnFKM0yAI5W0TFyiDX5w2i7UOi0cocReIw4NUIm+g238MhKNs3wGrxSdLV2Fwm
goqagaVWsk+Tus1jTdRMyfNagyoMXlZyfVWiriD2rDiFpQpgyQb90jHYXiCi0u7u
DkLvj/Y1nB5bWr4rWTTll3XQWXFoQQsGwF7yOHm/5/NjgmwoMSOqY92OmARafCAT
D4xNwAW7rsOR9+ocsJ8bcyC0/DKSx38JR2A+MOh3i84rk8LrNVxiXo4bnl60S9RU
9gyX6O/7CHNIaWb8p06D62Us76NPYq9W5JyJ7OEMn0pZmyBIGRT2NTsLlHtSqxJ7
1nuY33xejZBv9Z1ImXJyyZJ068GKa8v5t6fiJf72Nx9rVeLgOMdFtGM8dG9X2vuB
NiSKIBKWLtou2uxF4sUHH4hkEZRSYopQWiAzZEPYCioHu6fHQMNr67htXrEBLtye
x4z9qV63DkyMzFLeil9RCCuwi+liUo86DcGbPlViScywSsX+U+YA96b4+G6xugS9
7CcxPWC0xqY494njvBTlUXYOkdzPZ+PBy9ETgOCisJFTJthkxWVMXUeUIkmz6NLq
GQc/fRd/ajpjLvyiqnh1hbuvmR4jYR6niRqtZxOYZbFDtb/lrfQx9k6wy9lQ1Ehp
3iso3sM+AS2cXXz+t43UTcCK9esNkq6nRfJQHvH0nWOhbMnHN5RvR9B6tEO5ci3J
aUg7l6IwHKQu/FSbBZHUktPQyLz2vtEFrn0BC+tMvfdkmdZMvtSG7e9sglFVCsdL
7CLxcSSaSQVwDMtu+0ZE8MUk2WUTlssRiQ9H5Ecd0PJlz7UIw/09O+3U8QtGZGpa
i+AXN2aCTKxLYpSUx1eGHxhWeFHm1p71rRG3RvSsmRYXSD3/lPP65NEMu5eKF88/
NLSHtiJk1vxqJxyJh2rjhLzHGlcppavJSb6deSeTBBziPb9bt4kC2XnNqFXEhE6H
Yp347HUud4ouQwq5i3BYAAhUW6mexsjS/QhxRZDqaWJeqFkrPUornABkxsl0xJzx
l8godY2llfuYxRbAkmv25Ln8bjGAWyQpuDJjJVu9AYrs686JFb5FoirBWFKz/BUK
FA3p7RlONYsj+neVxccHgUSm8KymRH771FLMVJSIEySJFUs1aTb654BITlZ6Oth9
AMifSzjWoBCIJCO6PABMx6zwDV0agArn5RXWY0yBkJQkhPqZamtYcepjJrQRMEZ9
uyFjWOhhWU11MI+nAGWNZPFQbOph4bWweKxgsjNJQxwGUAukJMFoHGtYWmraF9iL
hKaSrVYThM4NRB4+97DSFqY0VaXktxsfP9Gm5bZrQuF1VjMC8sgGFHylN6NR8A7o
z959yNjwWb3arSe2xHcjIuoP6b7AB/VlqQ9gxWyOSWSaMlQX5P+abtAksh0DMtdB
dIYI4SoDjpWwHNg8x8Ojh1tVx2HIGYk1kpgGUY2CosNmSdCSN4w1UBgt5I3ZK5s5
kmknbOLNoXN2a1Cfm0k380h7l+TI0MRvYZ1+2fI9e/oX/upTiLQvt3GkrxB0DVsa
lkT0stsVEwuUPoipR2Tzv35zsi22Ytc3YMff+wcrRplh9kNcEVw1GVjkF3NVMQiU
EDVyseKsGvLWQrWIOwoHhBj2NA8sgEo9qg8EezBqiJGKi6EXbwsoCSRJtry7ZowW
MyUUvSfYuZZaB359dI3RvP2sxnYP6GXZVaxOFnkWNKo0MCYEq0A3KbZE88xKWl3/
5Iy6NTLC8CqxbKPJ0H3n9GoJ5C0cD3okQ4XlAE5mGI16kBj8D2FlDh1dQhxmNzr9
Iq4VD4mWT9S/Rm7GTKohNkfeZSiVfZVOF8h1Z2qu2LWTFXA3sufn0qjRQ6kuJYig
1sAQ2QN/GSmir6ALboH9Jj97a2Ow9+mmW0KCcMWxcHHrU0vPm9dBKiegtP7FopVZ
cEmv9+0NsvrYAkWTZCt77YNT2DVHRnrMLZohCZibjxuMK+sET5Wy4KGmBS2QO2RM
nKL3VPi7vHeRk87J8fAl0MzrDenPqABdvpH9BanoiKx5ARLxAy+2WOudM24R1QwM
fJO3Es+SE08h2CCUBJCbKcl18JlezXZHhDl82ldG5HIHBvEI3nxPGTwfP9y3EiHL
tWzyiBve/bz6SRjO7R4otuBw7RU/W32RKpQuV9xcCaKmDFDtZYQzetJZ/bkOwW5+
8Aw3Oxi9mF3nwbW0d/iDSUuM6RP1E+GzblFOs57p12p/VnuNhhCpuN/rJ+89KHJ3
ezgWjCKfa8I9vNa11GNZYhCdm42mSldiJ3S7y0PpaHYoWkmLnrQOKz8RaVPo8eLR
0ynjekCIAXLXJ9WDyX/Fhe5hEDBQw9yfvc0ODoktAsdQNkMb4Km3JUtdaH1IOuuQ
fBWRdTFhiWIqza5bCd+nHA6r4XQnj6/Mi5iPR1DsaUlc2nK3JXkfuDtKUHpwZ6AX
GsHDhXnaZjbCL5vweyfa46N+HsOp7/MeFXSmmT62mhFA03XJ3VLcQ+4hr8XksFU2
Q1ZEiGVnyfpsfo73PEisq9rxCRLJElkNJh/fbGjUQpqJwuSS+rwFG9OZ38O299bb
1SVHfsKHXqVf6BcCFF5r+55MGziBOgGaInV2YI8+cEiF7kRjFOpQsnMf9+rL2yeY
bMLtmWWZ/KDPoEYI8Esjl9u4bhDlbVKaPKNPhMSviFiflhkAe/qLN8m7nuLFEdt2
teicUaFid7QdO16ZjoLhIvsTuAwhwPycOrQJ/Dd2zfIkvANyvzMGoO2VEHuLpr1W
rOMQZLNmRRcege0Cf+Pkr6Y6uolAByNzHWJqF06HoAMlr6MynFNX2LvAAeRlh959
eWwVI7d0TdsyQHus3WHDZuXpEihW1iisZj37limdnznPy3tucma6u6gBplo4I7tJ
tivujLmyoAEp6UPkibv4ZNWlxxhl3HzSUjjnqEorSXmRjdMoqEB+Y+qpA0y3TK5u
QN1UQLC4XsZ7Ym6o+Q5GXtfzELMnJoNtFk3cUQrPZmeTYxMg6CIMVO81HHCysN34
UzBHxVY2dkTL13Md+uBbS44/hSje+4RQfF5pcgt5chrqXYI3Eb1uTfFxPYDv4lNS
uzolw5ST4nu2dLDRSQOH2NmKwkRX1s4f8iPS1KBXjSsnPim7QWRzkgDupRba46W1
rLyqP+ecX7zASSYXLqAr2L6FxN2ybdJdhDwwSYsuC4kbTZbNSru2nhKtQJmNHSIP
0UUsR3ZWdErnEYxQa36iF3Rg8TFICvPjhRgajff3UnQ1He9Hcxhv0au9UdGteaP0
Xt5d4Fgqqn7b/RttFgVDumnurqWcsbSkf/hx7MHwS8eQ6SHbiIf7ZCZS4DDreieG
z07IZiQGwMiCjJZffl6PmRuqoOO2QOkeFDBsM7lQlIgM4Lr+B/kvfLq2UuoX7qY5
K6YEMsxplhFmdfSGCPbWPRP+/MF4VIK1ZfclWfjIGPiDX3uyIcOMAdlFpglU1RCr
e4BqNDawUwcdvRTEMZa3zgJ0EtkGjY4TqXBxlpH9tBeHWlhjnzoFVjhXuyfP4wLg
35BgtSLtkMqtE/4U9EyCfary7jf5Qw6i8JoLnpKS8KvgSAVBMbwKPB5y1zZ7zR5V
q871rKZew29l2vvBrOb3ziZbdmcYeeaFJDV4NqphqoqganL7h+gaRNEXAOShiI1Q
eqqbTRjxk5SyX5pYkjZhvRZxWfmvg2zfjYaN13FOlPbtfM9UUZopKXT/F5OmfFzm
AGsU5WOKk+axHPDxL+0fzlsA48/QWfv7oliKmkTrNGs5yOasc9h7U2BV7L4X+U1Z
5v8U2/QWYiZNNYnpUoJOgmSgEga2aZ67DozuBWWH5qIn8L6p+8VJHWCp7Te9HdyS
+I2jqdLKmHGjtDN33/GLUvv5oAsHVemDsGEeQuM2HKwkWNQzQlIv5J7VhVUaL0o6
sLZvO4Odr3rkAF++tZL+sHrsnttVRvx2+haNsJqprHPEU4WLJy3i6GDhP6ChlreU
Ym13t9PLGGmLBsXfiAnvTf/zyFFsswqO+LKSiXgf5pEDjRujv/6JVBT2my26ioYk
UVQIYhN5ZiI3DBb7BKz+s4SN2rG5en+r2Iap5Xuf4joxdL5e/OVj58xi+KK0K2h+
V7wn+6Zr376KuGdqe6dQ29uc6dSu6p4exWYSI8G8M8JxRLIdYwmFPqg/pljo8f3+
iok9ueNEVaLfC87U/1+X8+oOWD9MnMUmzsq2tc+QbT0SmuK4tVDnbnV3mRW7+tc9
VjlsrYnAL1/KiEpC4s6+8tBhozOn7k9wUMowG5tpb5hf4iCpFj4IQpRPZ3+Vj8B+
uXH+ffkHFJQeIPQy1nUZIaYQwhoj/MnPwfQNf7pRzd/zuh6eUY3QGlINoDsiHUUp
o14+h4z0XH40EWL920+azzrEzrdPiCrFqmCP3GVSxU0jS/UQEeFuejeGewyAKgL8
wA9tRpK6NGA8AucgvdJDvVhqDnFRYeSZhODE4+6aWxZGN4pB92bYcMiUTkiuDALq
ACXlO+b2QJXOqBVNEHpGRWv0vwmtTDm2Ewze/gbW3B6rbftC0Y/BuhxlElHVdYnJ
08KuzJZ6ZFsoobU+MnQqtuU2VmFf9Md6Kr5+IY4n3qObXDyuNjG+Bg+fekRrbAQU
RYLSfBrNcVMShY3EXv78Qo9SZMY1GZgNEDvF+D+pcWUjw7hPpXZqmC0Cuh8Lk6cK
vabgZxkkh/meSMBggBC4NqGlkgfj/PET79tj9yTbazAcPiqPOgfmCueOedge0FGz
UbU31opB07NNMJ+6f3HwoRX9ADF37baQiX4NSi5w9ILUFbnxSSEN5iGD5TJTvuMm
HKogfTZ8YKFNJ+5e+3NTnZh0vIdpq42MEa1MqB2dzITfRDpugvtD9zSFzhIutRC8
HMOW8O9jErWydg99lCPmmrIaxFQM2UN3zIRMsu0RXCNeNv68mB8qJvQ922Ne/fsY
dQ3/SDIfFae9iynpicLb4fHbRIAGrp7b9gUBUZtaUnBbjnL2U2D5q+Q6OkyyJtCU
iPU4EOUM44EUVkTadhA7Uin9tmL036hD3cDHANgveIJOMifrsphESpXJC6YdqGLL
5ImKacHmZyKpcVkz1+gh+9LYDYe/gt6hCSIp5AslxfAp64jNj6THXUGlkWj/kQHV
vIfIBaWSccPG957kKvmNrRi4zlYblHS4o1/V2OChsEb0FvpQKpW35zUHi/hV30QY
gV0Eap6DuDLpU0YTy4/xcq/kz9VtZma1RXK0BaApz0Cj5Q4bv+zWm+d1b58DJcvf
Gpzcy5tuq8aTjJs6D7XAtMtop2hhbiXXpItYxkFwRCHBmxexDodqa64OKCL8qPoE
djUFkITVNj+oMAR+PKVFwsQ9NG/V8S/4NOA5NwFnkgqEsdWqemRJGyS2s3Wy2ETP
LiIbBGQhH9n68/+Lqo5iVqxRFcquN4Quq6WHyxzgEPI/KYtTAnnWpsXUTKiK+UQU
vf4/RdrgXtDzS0SS6QoRfXSZsfDewcqDOezjTnf+VIyoOXgdCX1RRNtsc0Fi46/l
HmKSRcmTOXjKK52NQ7g4VJNnk6kUs2dHVRqYBHv+8gn8vyw639IOdtSBZPRDVopJ
qPrIUfx3IHlr2h4X3MRDIYKE166pJOcvD/qn00x9S64SA7suCHSNcDERE0MPDKZT
+L8XtAwd6ytUcaDgAAc98yrhVcPEP89KRqvuYNsVDz3Fk+wLt4Bj0wAEsdHbOCun
X8kGht1HOFYIwB7HtmFUFeTcrsQiM3ZgoCi9uPh+LLJrdz4YyawgV8pkN4w8Wf7p
w5ka6jQ+todw4Jf7yQnTqA7ixmuh/7DBQvKEc4GoUZRoCcOXIYiHQ6fIs60yBUJp
fZLgafytkyJhWNPKELx7Aq7+vrD836C7y4PH5+zZ87ifpX7b/J/Zmh+4vilExsqD
VwbMWQQfDYT8Ng5cQtbNWMq6v8iKIc4taqnWeTnZy4G7yQreJv0H7C3tX4/IBqC9
UwE7IQ7OrDoau54bsostC7JWJfKX+ch3lwzQlp2O4v8/RDSH5FyxocR9CwJTW1At
5+7gtsPrc4WuDHbsS3l+bPS9wRrCg3D3higU35SKTZGkMIX6D25oYjDObHsAMJZm
NnvHix/nX+V/PHlXSkecVOWuJa8R4jrxwwKr+gybN05oEVCXPpJbXa2R1dpycf5L
+Besa9LWR9zCnccpMGVF4vSqEhZ70GdRW41vW9EoWGk5ChF425p1enHmiOynR52k
ERG4LM820JSuu0hiYezdSQ/4x9WjDaQ+eJtVUYPyYQKf/tnmxIJ1uOg6UwuofGq/
a03JQ04L+H4SMV35lbN5MvW6iWEx0JIOJNCgIyuZyFmUvd1SKKQiphDrlBZNpP1K
PSXKch4oEF8ajHKGhI5Z94EXucKoHv3It6DrayDQEkRqTf+pKRENIP1qYLmEqzdv
Pi4oriPhsnJaepBwZ2LP3I7k4ludrV/82mP8clPnwHIB+OoYiMQktDvSqZoexnBk
isw8uY7L7W4basGFor0CMc0cy41yTWg+9udy+rQ08WhEasZJG0hhi0PMwYSPl80y
F4cz+f+ftENP/6074w+QPT3RidzajBs2SmMy84pVdj4ci5cNnzSpfUpYYU7ERq+U
spyATj0HSfOFpLqEpvl+vpkMwhgpkLb8pnTeLVrN/oU7ZsXcSeL6lTVd8s54JKwH
OYkxEPzk03+AZLmZd9osRHOhd1CiMpnOOJbH6nsQ3hcvLW5jxsDgNByW/rYhdm+/
4lpjFmXqwgLicnDqbkPjZe5BuFSk2xNAVxUtwWyGisBpdfye05o+qO3LxqpG0ELb
IMpQ9j1kK+W4Uv7Ybf8m431KTxgrc1q24hdwEOrYzj8OJ2kKuc6TFpGzPqk3XTjH
xE6OclPcKYDw9hVNtBGz0CR6LQNsWEyUtN2uZb2NbYfYv4FRe/i/QYc5RzZIgBOv
9JiE1cOLdcz6iCpUUoyzfADRPVmDkpcTE/wZqpR174R2wgdAhQxM1z6PJJVe0ySq
B6HHQFu2qjmET03R95bQcSCul4vFPB5/AvgYrIIztt9iE/xqZXPOQgW46WbH+z8m
iIcI7ox/CaKXmtVELzcH+tOIVmBMo/rOdY8XLB3tjOfA8pE2CrXJBLBFH3m/tzw1
8addd9M2m+OXcn6YLh78rEd3nQ+S+Gsq+ndqq2KJmVkllVfLPvDJDw5ds3Ee8RcQ
Cmjwnj3Y/DCkHNLN0iorF+a6E+b4VX09AX00UUk2vr94AedWGlWZyUZyCaJVFQxP
Ylcq6v3ewAXpNbGiq2VGroyJJHl1bFAINgyolEijSGuEju1LEAR+1pRXLbqK7xSV
3yrr2ivHKwGcd7YN4ZZeOjnFdtmCo/i6gfZ456y1+yqc0d2BcOI9qg/9Da9ooBTe
gz4rZmqzx6YiX+FIlVZ3PtbvUYeBAq5BLkxjNNBKb/ypdqaAmotH2vjcPWS/kcMC
Z7ZIkbt2uTxp8fC9FVCS8ExeHm17ax45Dp809OZbC0s4npYWVyMUNJxCFYYhOcF5
NGqo0YoTWLePK9OswWqAFO4LwYovcqggyhFflCg259aUTcKjLZWfSrqjyyLO1EcG
xOZHIAuj7HL9p/jl3loqW/52hRVVnhD/aBPxsRI/TI+w+mKOuOzFzrZxaR3M5pcA
V9MAcmCIeV6XyfuxDq+LiwosRJ7NDZn4t1pcdsVEqpdpLr9sZb19JM9yMA5z/uPi
tlAeMQb4ikku7i4tcnkswJCSuD/wVRvqlcv8iIOoV1x/JO7L/jTRrt+FbnRo+/yN
/y8yO5E6z1pIsFRIGkJBOqx5k6yVRh0sEJSxALEoV0PGyJ7mutcmbmEK1MPVwWot
QXW3MwX5TSKJAb7zxf8DtRYXokMGtIiMT2wlyaTPTzHnvuZbdaX05TMVO7Poy6bm
qNh2mlk7ot4ow7kTrYeThr6AhUFSV33ir2gAI/qVs+daEqt0lsZ7F1dLQyhQBq2K
h0N2+h1PiSagwIR8M1Wimrkm6AYjaaKq6aagnuYOqmGQdQSN51ai/28oycQFtfCF
jRZuH/C4eOBYDQ1Pdc0zhZSOKjbw/BoJKFOO1KgaxL8PxQCLQx3FB7vriiUtHvCn
qaGARrQGJIk7FCm8WlygUewOWxjzkY9xB54CIVgDpT3SgL4naVCS/L9j0cQZ/28E
qMPfsCa1qPLrca2cJm3+EyrjWglnPKGsBj7tfB8tjbPewNCH4eXFlRwBzlAG4BPS
z4f9pCi4bvQw4ueW04ddw2J2B+vL2Elz1P13J77Yq7gc/Hhs8RcGonWPHbe8NYDX
amVbFcoCjFxXUMLV9wgyu9zR9pptoWqzZUqfK780eEl+fRYz2601XePs9ea0R8vE
CdwnkOvkId1r7vk1LrMb2GbVm2A7VtNixSUvGsHW4ZKC9dfmzinyp8SCt6asdFmH
HT17uvRJIWH5Wmh/jaT98wKgItB9/lkw7xPuc1/WVFalvU2WbGqAXPqy8fTbpbqX
p3Rl+SL/iuyug1wzZIA8+ADwpuoqI6G2hU5dRs5nPQmO0c3tiZRBOXSmKUupBMAc
34hskWTJUf63BO+6et5TJCTTdpDjX0nvI6ekuAbGuFEo8tmQzpmrkVjeHOABVaqP
bCX+YGB9VCJ2E9KyxRmLU4iLUEy5KzZzZoqnXljQqqrpdFAX/zoMkjmiJeq2VX0q
6IiwEi1tsyJq52SSvykAdyeg38XN0DBl9GNtPsZeQL4PWmZCNRMCj9DsiIpzvt1q
37Jf970ptlniyDd4W4B7rmdJMsfHngQTNlzfSUB0kURMRb+EYG7pGtn+xz3cSukv
JwADLw8klr6WObALNQ7TH/oizHs0tBnwhor1Ndl4peZarVqENdAhV0izEw+1Cc8U
I3ERG3mR461XqkHdUbLA8v/g+GMvPCaaYp46boJBAGpy8rTaq1Q6pZFt5Sq27iWz
WamAbfo5/Iy9vnIxs1ezuNVTDkTtCMFykiWRt8iijTAFCkMDmoE779EQUolIE3Vh
TpuUHGjt1wMKZA87H0A+YP06qRHxB5NSmZPxPw1QQmEq0uv2YOuTHObFBzwk2WpX
S2XbadAXt7oia53zl5pypKp62eQYq3Csh1gT78n73h5cgtyZRYRAvUhqIJmiUiYz
Y6392BP9fOIW/1p5I/0WkUcxLZLiqYqbWw8trtI7EESIoPR3/zShlkvBmywPX8Au
xvL8CrV9N49M99t40MIQT5+aV8AUCh8ejJVTudrW5r6WSBu+3lNsBn4v1uSRhntW
F13zOznJM2iZwfZio2RiMZcrnihFBZZa2vmoYwML/CLKejWfg6pC5CzBFCaEW2tW
+CAvTcOP121uDasjp5f0xsUoMEsYRfXIPWo6BRlQ2jo4uyLtSaCOPQ24Z+X3UOr0
xRLb2gJCKMq+otdnnBLZ561kd/rAxsVGuP+rqK90sHQGrWehJkRVYznP6Et3+CBF
wMzClCzEUbdaLjn6z18R2B2CiAK7pC4eyA9Lwcl/RX20bptfr3FAI8Zap9dHnkNU
K62FYeuqy4dobMMgwTY5J3PdMOcE/2soPUFYNfbdfPnqffRiOdMSew/2FBFjFbZ1
aJXHKShuMGIp2KTdSq8K0HybW8AND5ydqPSrqYe38x8l5CPSWfaMfJFFlaCjTCCK
pClFdRY9P8VImVBskK5Cz57V2AjTE4kU7ol5ZjeuGhKwlg+wp4tgGHi5V0b2ZgMg
4fAYXpCWYUUax6n2Ea4hzvXAGZB4Mp5vtgx8eUZrNwlCPoH2KYAsoDJ8pTYV3wub
u3QASO8h98jAz2vzsNHZZCpHbtzRNqBczobD1WWxn6m3aevxKXwS5pUKAqLpA2Nk
Jg3u8lHlr9/MqJGdJD7JlUPuJO1trSmObZj2s22ZpoFFKHQrkkVzqmzmXByCxlQf
4Q4/lyZDvvHk2U6hT9Ig1qZYrdI2mXQjEZjDv+nAuo9OUukXa6pdrJTyTukOk8Zk
1QKWuk8HyTKaaO0ncSCjxe26JpB1gVXpQbL3fqKjf5XkNEN4PGlAWFTNhoeauiGu
kMbHPtOtxRzzJjmJT53aEYQ5sUVdB5/7okU6NLpEJAQ/EXkpghyrn1+wllrvVcFH
oRikoTLy9SGRFVqocdWeR7xZ0dyd0GP10GGfizLNKUfqHJc/U+Ube6epfN58Yy01
hDp/y95vzjo0R2uoCX9QBebmyD3DCC6MmAaohdIvZPT64THxxa25lSU4sG1I0+D1
OVrcsnH52cQrrZWxEOGZph7wxczb7cFQagsjHEvWpTHE4goDEyRDCI4YCjm6S/ft
92dN1MOm/s4/cUUVn8Rqot9VGavIFDtBioKLU2UgL38FuDIuUh0taXYwPWSt2HXC
plt+E8Ae3kADpt6gd0A7Zwlpb5i9UslG2uYjTQlvv3E+pHZrkGT/rZ73T/PD0mvH
YOHvewwlQ8JhfV27pzwBlAOp7ua1woq8DPTMMVdtTCdt8+BDXMqRnccdimhcF4AI
MaijUeIigWmnE/fJEk0dUVc2lu1/PRjNVUzglnpJZ5biquyNil0GPN4QiA8jXEic
Yl5OD1k3b7xoSlg1FDFRvRVfa73VTy4JC8x7CqflNhKKQ0pxAo+wge7yTiGrix0m
djvQcEwI1J51icJkh5yRCDhADzmL+sZbWXqGDMAJNxbooRMmii0EsLz3OJFwPRR1
VBrKlpS8imhFwy9tAbXwjZ24fjBK4IUQ7oCS4Eszkbj+N+GqSqQ73xVWSo45buJr
hdP09HGwXpnqZm5oHyeODuJHG6vJDPngk2zLzYiP/rwlbY2E7V5/vc9XzRzuRMlo
u/AEeZYmmThA+pHkLEztLu4dEVfbF21KGwxhinhS9GOUpLtbYq6uyE0O3J2NunxC
A52bN9NMbf3BeH4IZGDR1QBwOGzBWxXObD7N3QT8eu1bXSVC8E5AgIcprYPr0KX3
y6gV4BPbkCvzxjZY2A0RNEtbRH86qdZsVBd9IfiYqokyfv8gJONfOO1aHEsq+aoY
g98yyuui2y5c4xB3yi98dCwVCN3/Kdh2PvCF+/9EGUAEy1MHGTsRGrlviArSHm70
vdg+cibuAnSjeH8o++prV5zn5RKjkrIORJNMSi13w0/X3C2qWkWx23WlLO28iweG
8sSOODVlRabHizsRwKO/pZIvnq4zbjAOj7Tyqd956X+Rghzk+/iWmEReSzT/EIKU
9hAJtro1/WWGxwpLlvS95g9YVgNQSYlYHeqjilCyK1c6IpB4xMt7NL10FazTLFMY
M0/cp4f8e80NEyRQTzOTgGxGc0QwMEZEayXnVv28BBSWCsrBrX4oOZFV7Ma2QCam
9pv157zGA47p1z6jFkg47mGJfunec089A5lvrHNlbg3GQ2VjwBdklmDM9+k6jNFO
jGSNEvOKoZu5+zX4iYjjcvJ1biGDAViozCpitUz3jvUg7A28FLebL/36K4coiXy9
o6sf5BiJr0kZhtAMtuZCidZzrwIqPMc9PIbfKWtEdSLD8RlPeyVJn9MO6Q/sizqS
nNCnoTse3tw+MBe6+osN2qdtw7ESZAI38cIg08mwv5woqZ8hWc9rvf5VaazEqgmQ
+XP/Sf+3lDywWB2XXD8dTdWC9VsGLZmtM1DMMEOBVTUEg/u7bzMBx6z9090QZSvr
OZx6c9MeZyVkUsNUhflPcggUf6FbalPqf+qANjFpNf/VDmQRJPkFJE1rsaH7vokJ
q56f541QEUoSurSAUjLJE9iGvvQz8GFJP4KJApmqM3Tzdl5i32tJqzfA+Pcap/rO
zkMTHJiP2OCy2FynzhFQdYLjXwMrMGyUnuspHCK2ZhwI9ExbSI4L0gvOwc6HzGWH
H5fuChwWe0K3aFCyOkE/Ff8E/hbJ3T22tdPXCwpIGeKrgusz2YCHLxFDbA7qgeIc
B/096SzYX0JQ72+sfAV1wuaQPt1Guw2YVef5mlmvnW+rq/iPtfY33zafDmAdwRmy
7tdD+eu2gKmQCOX3Hk5w+G0Ey7U42uj9I+5debsFIN86RkB/Fx8n5AUrqo/QDErN
ABQPR1e6MAQAKh/vDzAc0mfX1Eurd7Pxzaj96dMnqq0OfuN8TtwOdBdkz4SP+vCo
5hZoUz11Kl85ql4V4MpeAMV3J3TTdQcZbwhhP45R6JQ4C4oDL7qWRuy21dJnk02a
mQeJOzpLGOnf9PFIGiIeLNXpE6IpaTsMuZUdRXv8WN23EuHQQwzvNmgctzNrsU2S
9QAQuvO6JDTmLLbzCKzZh+883pW8KMK3bmTgw41ESGuSW9xEeTQGBH8YSgZKbhwu
/rxTUZ+8AbXrBO5OGwQv0uzmkqMzFwGW4cZvWFF45VMlWRpd/yw/cujSPz6sBvU3
80UMiuXYXX5zPQuC7/+cQKNuFH7eCc/AgWhVbZRB2eiQU8IWhGUc6AeSWddSqDIL
bfK+DjNIyulCFnPiLSHN+7iqrSFVN9hkjx8fpcnAjzH2KcLpacWHYraO9kWBsxkF
oGq4/DJje3rNRvAxVf33cVtYSAk7qV97FxZofIcPpuYOvCMp/oOxL1eRNylsGEcA
jHgNpQIDm3h7YbLVDZmcEoMI0aQtpSy99s2FNAU1UKhJc/F+dL4juimh+K8Lka7x
VWZLDls4i3taly1UcMYMm7KybrAUc2vG+tYPULwYhYjmHQy0bp0MGFoQfW71eAQF
HrvX0tCVUMUMZuhAu6n3IiDo409RfYEFGUi4OjMMStFVbG8wbnzyEe57SUGuwofS
SnKo6e3YlMUrvwcaianWNVWGx0wPzq9WMX705GNhmaxYFPzcIG+tZk8Th1wuD3jG
NY6/0rYyoKXDVuYwoYgP4U4DckCwOqUTQbaJM69WekYYdGuvpois9H4wjQea+Zh5
yFXJohnMjy04nobbC44GxlDCyRlIWt8wKV+yQyxw4jRWREIHotmDuwRg8InDM6j9
CTo4B2bp7650R2V7ox9ivMnP2YQiE7Nb8tRP+mfgJ0ZWFzVT/eD3/pnV1dixFnoI
7ig6dLyKX+5e6qGyWnwoMoBzp+1CCc+XYT+UfkNlQ2tZs2XZ6jSUfXUojhwb81OK
RQez3x1OUL15jZbQtcD4H2+NgA7fh7HA/O6jrBWQUuq0XRDOvn7ObRLJiwtti4ba
SZuStdvhcfNrhUHUlobFBHVwHhG4rBtoNvYItnWZTsLR+UxXeLECM7AWBOO7m2JZ
HIlqTXazjEJX2iFaqsXDZ/P3O+NZ8W8jMAqZi/tv4c8LCEQVUwZq05a3w2OBJ4Oi
8O1gtLmiIadXqe5obj0qNmngbqr/2Eh59R3SA+OZRnfbicXufOjZApqLsw/0a727
Gdo1oNBruK5Ka3KOXMlgiwbY6m7Ym382ta4yqpOVRZKe8mjA7jOAOyPp3qn+kmMQ
3a3QCrbyHdk3bt6Ux9jF5zpUrD4CD5S0XKQsTNdbngB379CtScnAOYlvgQFXF/CG
x6BbSgnP3TA7rGNuwAc0WWTXMGF/marI3lRwb/xjBk6IP6e6qalVdhvIRJ2iOKx7
cklvQ5irJvygjFv64zJ5wKlC26W0RxMY5pFOgsLnIrNlQMzfCe0K5BZGizQKNIM5
pesPA1UjyGe1R0l4bAk9vjEKFm2OXwH7j85bOES+ydtvd4k8XyYMYeL9BFsq/x4B
QD8cmpsjFG2OpSCwYOjWpdt0WGKfDnVX34sjmlLEfCFF9ycFL9heu5RWy9htmM0y
MW1CjLXR6wocuOPnXuHCZVZl+zeIQ5UBdSb5C3hnQ+LOh3iqLGV0D8GHA0W8CNbI
/yqIKKMgP615oyJPR0GAFt4yHg6ZWEOPJojy77jsXQPZQU2t8GepAilmowbbFsj6
oyruafr8JoByshmaqIZvUmMCzj+eJxRaof9WGjo7GEwGMad4Svp3YmX0x6fiT0g6
qxISEveR1uZlMVBlJJeV7t1AcX2sqijZRaf/2DsPXz0lAalhTO6hqYhMVI72YVvJ
tp2LF3QrisYpnfJPyLiebSvsRSDAStDu1YQ/0/8HAoakV6uibie2yBHBFjGDw73F
locvtMIAH1se9fq5WqrCdEglkIRMEvV1npFHwRLjoe6J3mT4EJwgtmfhqrulbJtG
UWGECAIK4EMHZmFJgGePBS0CjJ3093oV+V6iyRniwWJfGkhEEuzuBP/raaqgGjt9
UbqUoiNuoPV1HypCNDP6NXP8ZBHgcr0wksoH6GCAQ10o6Zs+BmuufzUwsG0SOOPt
eg8kNgLXWXCuHHxIpOkurFVhOxqZkUBDTqLonvLvQ/IufYize4/aLgIw/lHznpWM
J8DkmUBLYoZfJAhrBUSlb5fk4GtA/8o53KqLIze3FfPjrVdlFiNjtTunUicGaogs
lkBsvA+SLP8BdrBIKLz7mwhVIb7mxoYIkMD2AodAaEMrKIGnRHhdKSxjT796QW2g
JXkFr7yMHwnPHmbfnnd1R6qzxahISFaHskNaMFWeXJ2B6aoX54wRX0nSyat5xM4S
uq3IZBGR7imQizIplv66ftIcIwoJTpPIithtBzB0vXN9ReYdsCzFR4ohM/moAaAU
QkojQsKBedCVY56o3Z90CaMunFqyyIZPAFBf65NfAVuFmSFqshiCqGljilRe1gfE
iiESKBDvj193omLQ2LIkb3PV9voAcuFoW772+QiAbSTt/VtgnVmyaPX2vNCtbyn5
yZd674QMOt32J9Lr01W0whngeq3GbnxEnzV9ZkIFR5im1e8SYokuyg4bK2mokywv
y5iu+2VVLEaugmSSJfGX7kqFOu/yYD76iR3HAkqBQDec9D3LZDwSEPaTNLwt9Ohz
ZqFAa0G6YdbuaQMYw57eEu2Vzw4LJRchhTwQhwgEwOukMPjB8bLHj9z9j+x7VX5O
JEKc7aiS3SmW1OcOTTrmvEig8eqk1fyYnjc6iEOijVgUKtEilY3bWO3i9vrO5jpI
yC2wnxdYrGm+PxGBf15bSRrOb/5HurDeWSkhssF9Vsmf5w5gz/dJoEe4XFTjc/mF
OgchGXcAoJq1Yi1aiZbr8vHWrlroF9sjsRCpguV8UIte29Yp7d5/Glv0L8dXh2KP
eLQlUqQOe4H0m/dRcwngTeDWb2RVfaeJWm8Dz/U8PjqJKpsjsY9NGXkBW5Xq1lmK
PMNUOcFJh+rbqLubrDNw1HyC1U+YD+xhsq5BwauB52JVmhpahevqWj+txylGuTty
sLYUflwfFcWewb2RD3wpt0VBS+0rtUNBqMNaJslhK6LsUjAz8xfrwoWB2wPAjL6l
57cBeJGCadje+pwLJy4U2DuRBQdNFuydCRjVBPvy2wlz+PMl73PYpkJU7+7VhrFF
PGdQHd/S4QJaMegB4BQOVBYAFczT3fYBP7Dn7NjxSIxJxVAmgJ8ClTW5R0EAg2sa
q/OqvwZ+AMv1PGoxncOMQhfKbiZFt2uFd2wCH6Otihws1Py9aAyUM3ETWC38LBpR
zznl8ln6hDo1DcQs4/agzM+gnIz0iRRQdPVhJhkC/N8Le0Vb/F6l5nimBCH4dhnI
CybT/oZl8jxHqMV3rSkBfBdskCud732KbtOVgUzR38KL/Q4KCbN8Ygi6CYFERepZ
SkE6eOzhzgsNqs941Vst6QWKfmB56WIDK2iQt0GBjS1wnAy8MhlIAlk0DfgAUFVd
rbuFYWt4Q15IYWBrW+qVjgT2v30iUMviGVqYTP0w+XQfOfLON8Hh9xntZB1GWU47
HvsuksvdPYsbFl7o3G9vtlUwJy/yPmAc/UznNFuI9d7sCuABnj1aWZP6EykT10x5
7vaa8y/VBl5vWjuBu9lETXOItdQk6UydzSZtv6D1TNQcYHkAOlmVYiM36ayopDyC
MGTz0oKYnN8/CYKtEf6PrMn6VKhpVljbY1560IlgtqOtNJ83aSVQipabrNxR/wPR
eN4WQjoveLHcyPhw91x36PLjjsAAh2UfZtoZQz9bHTfzI5+m1NsLdGhyMNuVYGm0
22+ykX5iXKbxYnSbj1OSEQ2oJnCQKbd/XyMD8Kv8SCUTAI0/3+4w1PVp9nTJCjId
9ejFEKU5WFJbVjlT2q3qWBQofZvP/qgszSK6KZ8r/1I0NlD/+nWV3H+XCZFobqKe
f2cCYlPUrN4LWee1/jgl+kckZDmbN/CFx6Mnu9SccBb42iVwYwn1Y3Xqn0BhPrH9
1mJrBkj449XYuOec+H0hYAIMrFjw3vO2gSqiYMghtjFsUWV09Q9o/gwStU1sx398
xklYDvGUCP9L4F0ST5ziCmIyfK61CM8Lu7xR06LnVx7m+3FQXMRUfDm2aiNXq1s6
6A6xi1LjEfGOdrMqB0JLUbrk7oVlTqyJh1Kz5a8pCfi1I626V7k9SEKZ5ozEfZx6
EWHnbM933/EKUzb2ZAQgQSV4BhQQ9hUwh2X+qluskIoYfx0X4XMu/8ipm0NxQsdd
S1t0f0yzwLVcn1LXjbWpkoNA+348FThhCr2+bwjcc2UbL3QWojsuaSt8BUi9G8V8
dFEnu8AJ80ijk0f5J+2BPc05dbPwlEunjUTPq0OK9LkDlej/FmmpfU67bgBcWbP2
6rO83d9Mi+3ierroUzWGysAGErb6JTEffyEPGB1q1WAT1CEOFzdlGhQreDdXhdk6
wV7sFA8xD73zo1JA/n7rqrnM80JmSH5QjFuvoAUQMpUureJsdktZccO+YFjdYjLg
kMRE2wiWPvB94asPwonk6v2TgdCFHUQsyLBdS8EdrbeTIVt80J4H3z+fnzywEFwb
umbB1cQ0YpJrYoPW+0SfPJrMR7q+1ZR73Nyq70o7eEVw+cbltB/cOlDQU2YZQDpV
usGmQnHZ74luraZ/pNCAGIYBXmSWjbr0cOILf3kEwTYOh6AyeCJl4QenSIHptR4S
zfXW4psoR1pnf3pzFik2JkIWlnpp6uAzhqU62gNZqTeRYl1rg90g3dB55wyCms6z
HoakNJ+V7rTu2u2A+5PPwsPzkcuuu5rrxmPlzo72QsC0DsKnrqnMplbkblYcqkxl
l5G4YUoEWEEzWJ1yXA/hrobsSjG8cFyDsvhqBhYfNyj65a5geyejLwT7Rmz+5J7Z
vCzluAmzBYtwP7ct4lKXIUP0khzh3mClX0qttkaTp1s0eMRDyk8eJQP7Z5HG7DS7
1IoH9qqSer0+pgqKfNmVkWo7xWRGsTmw26ET2rlvM3Ne5KpWadnaZm9ZLrMKTzGQ
oNt4RlMlpH0JtrwuOX2aNGHXGWCOv/iWQXVkpCuQzWG48Kfijq8BaqLR4WyBc2ZW
l9QgnNyU2faa2OGc/zJsmpRNQsNa4obxRf6+D3PVCeW0+ab3fbBLkgzRhzfVjtj5
GmZXEH5cjz3fKGR611Q3MFJMB5B7vPOC4D7IcgbBNP20Z8852RxiqC5w5hlm8rSU
SrMO9Y9v8KeBuw1DSAwtlHgJVmblSNbT8Fug8ZnQvl43+N68iayj1lRCub6eTEx6
wMaLeUOwusqXiy8J2+JF1FecftW1YT3J4UM2/2miJNjPK7povQxT6qB+DOo95xkl
gSzVHQXMyA2sX5IfjtWSTDA50eyk+XkD3O+O/13YTle+DXHfavgS8WMd/JOeGQ2s
OS5sOGTBx683OyV8GTsP6uqLo8HSzco9GsKIewcmuQ1YoVM/QnsVm5vY5nThZHyJ
V4q2HH23EwoLyk2iMxxVhFYmbUycGbH/r893Kv7ISB1m3DN7yUhk6vbTn4qjcNj+
OEm2dPeksda2cvnv1c1ozNjYCk7hNPzeBpFUXantRrkIjkIFo4oOq8bAWBG1ugle
h0FLh0/YqE0qkmN3YdI+Eq8hSG7vO3tPO8JvF2kCPtQR63oet4fJfUOMvvzuVd/z
+0YMAf4PpBjZDJ4n4pxn62s3PAlBux5nP+ENevIcWIdBKnlM7XbOG9vxiznGlj7Y
F5sMFTjTJb+/56QnNr45nlKHTr6Wi7anH5N6uL/Hbs0nPPt81oG4Abv12DiwYWn3
R6EBx5skR8Qx71Q3v4x2egNPgR46SYWewIPSZZ97YuBvn1KnGmEmV69MY0nkqYOE
lFlcq+07zbaW7HJXbYmeo9iIfdPF3y7IFDhxLCxV+runzISIqoNGriFN+PUoVmfE
jgtRtp4PJMRhab9268cNkwTrU6QVDAuoGO6hdRsUEvI/cy9B/oEfixxAy103+rbf
DDJnNRBaA49nNe34mxE+pe/5XBiJJiRiEhTQW1bQqZeCV7QsHClO/Ctah3sBGH3z
qLAMVgxt5XwIOhpDqvAD5TFTW9Jnviv+GN8ayBZsUGEhoukSusf058d0JgwU+VmN
f90JFLjhSyg6YaWiTsU6UWLWxj6eG26hv9O5etWtm2pZ3SAWKuDk+iEqvhYK0esl
Kgg3YRZN5fNMZCtccO7Y9CO7dlNL0Yren2GQrTJdDOanHF99g0ENJirYeGwn2DVL
wctLReZNGG33mNYlIdRNjTis1bKlz7juqBvAE8OUT5ng+E8QzB4Z+9kyOQVzO6xh
1bGpJGa9V4DzOu37dPI7TNRUiZXxohnXZQizuSRkR9VzkIoaB1pRTGAV/l0AX3yu
3k3TgbP+FK6AQ75+4RPFXb/HYGRLFCLUJu9tlyJQa55wW3TYc8D82qnxYHzd6g8+
FHysJ7BpGmdiERL/wrOB4UYuQRmhAgWgmL1K81Zyfxf1KZtP9SkjUgiteK2qDxrF
UdU1vZ41Lc/knBzfEYHVeudaO59d1ciUrW8eVoSUR/lwjfJodSlEiMiZ9AtHMr01
f2mPc8xhvx3GqpMpjdThKKKr6RfVZLusIrLaIubDFzz7q4C3uwRQN/3SyRyonptp
/M/3oqkaYYqwtqX/tRjTojTPx/gYsbPQ/niTHzPfc1ThLGkzJhyLL6FV1U4xnsOr
okGMmJEybX1da2qMO6KUQOLkLiO5G6ByJKgUWfy3wGw3SXmoGLfLvRatEbGMeH+N
xvnbdrq0mSNklSH0EaYaorPTWTIlI4U7YKBy07p4EnRHuvV6hBOpFGUc8kwo0rWQ
NjerFP6MhZesIYb/CIn8OgKe0tYzNbvviUX3ZJkmRpSo7IDYPnIE64xspqR0PRQH
ere/J1v+2SNpxDCnlvVumeQdcggRd/wHclYcS8frxcAL9e/UhWyCN3uq08sSn2CN
7LbSrxxXF02vBRxc/JO4wqJ6M3GPQgfGP+Ln069KNWyO21uSx2mgK7KFEbIWSpzx
eRvTSilaJNTD1Jp5tQZR/r0yYDpTI+N4NMiE3pXjJFI/ym/2tdH4kqhiT6be+R3N
MjyeJOKRdo1imynkOheMk7BZ+uFdtl+LxPBfIvzasGm1q7f/YpCgkN6RJCZPuCpy
PU7xCS/BeIh3K5c48jdr8qy+VmA8ZM6yQ9vNZO+njzj7xykgWXNWGxbcNySygkgD
9M7lefxeDTS5aTf3XMQjPXYJkJAcPfUwgrT2pOlSeJYAaLLaotZ/Zu2gSF/RDGys
CIKNEy//3alD25v7lzOj7HFzGdjQo2433pkCR/irH3RxtsTB/PhEhhMhozv94IuK
CjwTX3pfMNk4ho7aqf4kbRfP6uU3kqXpqbb7I9b0eijS91C2I7kipn6RVf8gHFCi
eBjRz7ZOeLI/GIPkUu9zpKXK5uVScg14s6Ix0KU9pF50OZcNhiZhlIBmJU10NjPD
NejnxC3WNulVfyW9n0we1Nr9yvo7tKYjPso7wANaXY2CM+gB1JAAJSH5uzCdEhCU
ANwtj/H0QCUXj0T0RfwvPR3HiGKvHRfJbyxfds8l6ijgAck4pVk6C5f88doNQnE+
Oggc5RlNJeSAZ/emfI6tngNuQHfvGaTDMGWoJb+l23XInohbyyXgWtnJkQxHM4Jr
SG5griNGdU4Fng4CrboRXbeYLIwVU2X/XPKzA/kblRNw9swh0l6UP3yNXa3neMDJ
YJXmz61Jb8odQRKfUbxNfVqM5bVEtV7qjSQwMKwjj3qPzbiPTmUjYkWa+OcmTQiJ
oPS70BgKrWUTkdZ7Nu1cVgINRknfNtBt4hSppEieY8Rwiu/jEKlB3F9srjTSSDNn
lTOJWtBsf8yfkot/ziISE7TRriAv1wR+FuBDKkq+u+vIqYz/QxX8xluRp8TLBR4a
cNajxgCQrhXZ82/RTYMDGIepSjSoY6Yl7WhvvLbwsAWy6Sp5PmXBuO1kWmYX5rlw
tNezeUXwKeA/rEfeFsVtC7tn3aorzdl4PPXCEEBkXrCbdB8I4zvLHsgSQOVA9m9P
jeE45wOn1m1Y6gX6xFTNIctlxWH0ux/LHbSzEk/qVp35yNAIYvCuDAUEvL3/IloH
/ElD6jz6fOoUVkcNOnf1b4wgnMSnaX7eNj6WGesFOHucGv/1G0PoOaX6kivmo5tT
3v6gWKMe4DdgyrWueXsqOiQfdd+e7a5z9KJVpq1nAJxNHVqJyI4n5RbutNU9NuMp
vRv2iAmnSVw9PSQzFEnkNTTEQjWqnUbc+WxmRJzxHEWAWanMlbfLQfG6ywNqQKCM
6HILm2kfQTwCFdXoysLW+jkxpJ5xG/TtzCegQP+9kiBi6wExZ6ShdhFwHDRONh9s
NuTmdwWcsXwG+l3YkPDBYhLNvhqtCO92y0jqIX94HsV+aBH801oIPk1XjuwXEEHN
M4tB5lK3FP7CF3KJZsoxNyOC+JzQjOvUDjmGf3WRz9F1B7Zm3USnVdAdZFNIyN99
90AMqSd0FrY4qWEgHZHryAdfUv9yf1pijCtnsP2Ax4UbWBwgzJeuTDZdmyDKazrU
xgNlryvB+UKq8zjNN1/hHITpdXfyqrzLlAntdMNcEL5gkCKrcdrNCX8c7ajZmFUX
sKwu1PvY+bEEZ9B2EdITBPODYmH+UNp+99YzthPx16QusL38DOTUUIoRU9yjK46T
ve2+UEEyqy7rtczQDI0/epPUIJZeJyYJnfVeA7qqDhoQI/JDxTD+XEsazW+u2mXi
+WV8i6QwT1lRniMGdysQcXxfjIEvKhwRvLyDGH2XCyocol1aEim9P9jyVTrLG1Tx
A+gJX9L26G6ZJT8/Y/RLXC/VJryj3KDuhUZu04jUF53JE2hUEYnpEt5hYnCRRBr1
Gqdo05JqWspJe/9LnmmiIT7WN6BPutPsJscxlysQS4lOko2UdvtxK9sPZ7y0Z166
Rn9rBRXCllO4sq7763n8VJtcb81hwXyDdi2JzzRhlBMtSgEznYgPiPlZsV3qgWdc
v0IEVBAIIMgip9y+YzvGQaG7AZyIWWef4C57ZPjd+X7bqFl2oi+3yrgGMV/OEVdx
H5Mc/Q8RdVq7FsINQb5THU0XKoSooIqtf4/F63Qb2N/SpGwAqe4NxEnd9jUO6XQb
lri6+hMYAIz04H1ybevwBDJkNXVvS8mKstuomFesQ0XrC8ccHlMnXwmMog7oQWRL
7CAxIaJwRm3iZ4s6lZA+AsjJsFNOcSqUQBrU/Ko3ho6pUo+2a5cO37W8w1xULHH4
ThF0rV8H0NBupk0rLbXHR8WRnsv1ZKz1EIlgk468nS8NTMdqehwGHx6c/oPD1UtJ
+RCDWU5tdMTC9w+J/eA76jdblFQ8254VYnu/MDRU8tgB3QKgc1kGwRzQjpsjWDrt
A41be96XjrgxXTmdHnRJwg1ICCbG5pDCYg13i6ktkxyIKGBrVhTQKFLGH/IKMTSS
PikuRlFl9Cj2K6M3w87ie2Hyhf3DiJwS+yH8wbyNU1wUkBoVV8Jz+oC5K9GgtyJj
x3t/9RSqrj6r/+tt1iSAuuiAAn8MJ9JUN1Vi+llzxCyqWbsGxdAlpdF4SsIQoDgR
bDRJ8q81qvdu+jFSzz//QMHigkmdGkWpRIMbPhibCXEtb700xv9XrO+kB/oxPYnj
urQeMfAe3GrPxR27R2gloRDpUvlHjwlGivOYTHVQj8yD+0CWIrp0MQwHCy+FVWT2
PUgrFJnOAnRoFIJMKRUYyS2CmHcmPAW+2KqwgDMRVBhz9doNIlBp4TTkanL36upF
7vmGMTHM6U9Y8JCxIKVGrlSWDaFZacWEQQRRRGdOX5kZF67IoOQQ84B+n7/UB6tw
UD+ei/4gu1PLB79NHckoqSgzX7j5Q4n6d2lfpKxwPrwZW7LjiZydPRcKTMDtXZXS
4l87TUAuHTPrws3frSss+WtURzdTOKL5NLgWAp2lrYX69Wk6gsVgUgUUbP4Zp4zp
3ejZAn62OzPjoor7/vDsQT9awsxeJL9eUqeOlWOIsukrlioC7ayYzWubu3mnilum
ljhf2AZZVyiMBmA/6qKN1O0cjBgbnXso2LUsVXdKS5bnT72GWNYLC1Tv71HOlP3d
i5x5GQHqWX/FTe/UYUdmM7iCrLrVtRxNFj0eOqW7/Ru27avTrozL8bog1ZXfafik
Av/4KV49BWd84p/keOIiJnu28ZYqxVngdj3g1iG8dLR9xyjHfy7W6a/zMUr4AOSI
XRGjB0viGUmQy3Fi6ZyXyRtG79TPj9WGO6LgG279go1QFAr1ueDR3n9j3MwL2omC
BP+xFLur7jDLT6AlEpMS8hS7NNQf1zuztXt+m51TK/L6wCUVrSqsR6sXx5jGbj4J
CtdCVnhGAQsCXqXF+z7pnRE2DQplb33ORXtzysgvyIrGOG8Wh2J/eecv3hSui9rb
KQMss26ZnWJ7bf1ql8wsaDqo9HbaOKTRWpucL/r7YaGaBcfgKish4mB7tgob+kVE
AiOuQG86pfN7fn/xaduFJzlrGLjWHn5YU91830l1GhwkeoLYqmZn3L2silY1HRdQ
lRSog621iTxF72NGTyJygZsftmE3CHcXu01DeZ/UarCgUvfle0AqalWRrkBxWLhx
mfACvF7CAEQOle9s+IbFR4bk9A1zf+bVj0NJMG8DHwmTCVye4sKqQTdItrnsxDPE
Thw/doroUu4EAc85TpD+5TmYf930UxtqJnowrmhKeu2mUVFot9cGGzzkmDg0pyIQ
/xuCKCvSglpEuQAYwFnZKGp1EXsN/Uqt+ULbitznHj8qtT0KhhZBQ8dt3vYIz8NH
8iRXSu5Z8xwa7OlK/x6uvZs10OGnagwMnpCkpcvBCrVgwR+MZ9SXVcRRZmG6CcBy
L6SDZ6/Q0e/4Vs1uvv0fzCYKiNJmRonAG4uK2+86y5223nthWM/SXbs1NBSbmrt+
j71iz2JC3bEI8KoT47IyWKfe5Ojwm5spaVaC55xV8ad4Kf0oW5TjT15BYSimNC6t
mHopjDVMt5lrea7+kEWC9VRsqnBhQF+YP7tlSB5OuvejE8WcUCnkryHD3gfWLOnH
/s4uNZYDF72wsOHa2mhtP2IyaEH8fC1o4R/ICkfiYEi+czdG7TSBzpEUSnFSt5rl
7KlFh+lxEhq4sjlEbEhzbeNv/SacUon44YPM5NJanJRWUqfX+ZoG9Eh3CyO3XnVN
h4xAgKTLH2219VJWsauSRu7OloPWj+TaxC7vE5uiGCqa5P2dboelNvDxnR8QHl1H
qh9vZoHLJnoYXbE06VU7yUoIfxguVp0mGG58NTfK8uxLcuH882wBvz+RrFyF3ZdZ
cKUmDCn4vckKsuV/gudzbxuZUb2Bjgf827pWtFPAv2PZGUE46z8WkmscgKkgdvLl
QwzOqcK/v0xZi4Uh66asmBbq91auDuBH5k7oyVl/RtJDnReK9tIj0mVtKpSEPTjv
0nLsfxnAKD5bhV/ZuSaTNY3cz05DSWu7Tl/NM7kBj/Xn8A08J9rie+Z7wuIykQzw
cVDI8P6yJW4GswKWsg0h4kbp2mhCOyqh2DBao1LSXt3rD8MaAKYDmcAoDPApduQK
aBF8/U5zAONnzBwjcOqs6oJTiVTYbzdLj/NgyDrxHurwmMPmlITW8bhPCLxiOYy7
1ld/WWmWVHZWItcSRy7Jd5+ggdkKT6hc1k1xCopM/5DoQztRCEc7edvLV97JWF6L
jR0cTpdgXBKcNb+bWs4OxHwLQMh2VNlE/9cHea7b3u6Zd7qivWAvMvXSs54IpNDs
n7H1TdKC9NSaY/QCHt1HKYgVI7I8U4C6wgI+A58Q0VeX8FwHKSTNdZk6j4ohclug
Zj51Csvr+cie4/awzVUTkQa9/3MYJi59i24vxC862bkRf5AIEUtrzjF6nnavGVZp
lpoTxMZyjr+acNMd8yIvK40FBDkx8Cp6gi1a8wkSg5uwGhBPfSfK5L1IAE8b6vx4
EZBk4BEjcrNIvSKVo4pwpRfFbDtq+8Nz35Bj2Q7pBxbIN8WRuuZfJ5dFj9hcgLwI
bpoEl55apWRS8k6gqyn95hyL/vEJi+N7jrLbbHF1Vu75irsYu9Hipi+Y7CpESwmJ
Ojzj5fo2G0TdZJQisoMLfP96YGBa1KMl7M57MRQqoGHDcoVuLIyIht5qLU6bTBUi
eec47H8GFtbbL1JWkx+3/exo4fGfwrI5g43wCiXChlrwtYIyhRFz0cBK4LKg9QrA
b1rko57KW2c/bKc6CjrtbyNllzCDbIvMFCs+BmwzIl6cJwV640cSXNQxWw3qYzSP
Ae415fr1uH09bNYzfeCHSVnCLfLVNHJbR7cT/gjhjKkdqMWXE+uDc6csRya2AXCq
wBbbWU4bwhzAuYQZa/n62CsiGjog38Dd9ohdtN0+Sv1Y1d6Hn9PjN8feYwxOkIzH
jalspJKTartcbbMdEJnE8ri4ZSodXqpbVdiLHCEebZ+jbrIyhr33sRhXQaIFC0Xr
0XhvB35NR2tKDxDQ5SPeJXSELIOvAP4U2j559pbjSYCQs4jaXjfeuD/IK3npELzA
ePq/zVlVkai4VaVxjMoNckkf15qLHKTuc67qtRl9Ifexg5BOXzkfYQHXR+l04BkJ
G428b7pmdjB120OOzqNyl+UuTKrvxZBMoOMraryZXvwpO5FNO6dySvL+mAsdAqsF
oJp55enNDVGRVQ3BeKMbMIn/hARivRZqv7uWMe9/fzoHD51uQAoUUTdJlhlNilRm
VOMs4yW6HfXkQDgFMyi5ToTe+nYxghnWQ904XxDKy0yv4o4CuZTiDfns3TlGg+ur
UXwnnvxrMTX//3/y2pyvvleQ+t9EoXBSTP8WSdZtnOUOZr4w+PBoME+wlN19oMek
XroAmW1zkzjmGLVXW52IUnQoGggcbEtxxGHcmAcyBS9DfMExisTDnzevGCxiGkXR
qwSOlNbCc22FtSYNu5Lqjx9HW0kIMCrbzyYk00JZqvaOglf1YJNqIQ1eAy7+X5PJ
XLR701cDG8EzJjreIyOFlW4Hm8HFF+f5flkbX/Pr+/d5f/0oS+uhSTzX7D5tEGt1
GHFxYdJWQc+83PQPpZiAhzwfbq42d/y+t1IcYEfYY8xU33O/FGFJgr6FYAPoqRGs
59nYGk3KvEjqO3krbb8YH3j5Q+xrAiy3+fdX/w6Jrh1j687Lgk6pQHVlQSAdlJjw
QLUzSrGaQKFzTVJcZ38f5ymZ7xxThGmHA1cYa4WDulDVUbZB746ybYk7BWC/1ksM
PSFA1QoNMnAAdJ4PtbkKrHV7s8Jo0iWb4W2m0xDcfkfYWNYwqoqOhXmn2feKFyam
dZ5HMviYcHpx9UVUt6Ox4K5IAUchRd2mxwIXzJFr52w7r22I3zw0qNpc3Q5i0PfI
dGijEqWEVmNDL2sct65L1C2k6iN0fa2Vbu1Yszv8zUo64Jnz1+nAR2e8ZuzkbGI7
NQw1s2vdGSTsv8bfyvhpaqo5kPlYAR2BT3CTnZpG9mkLzKjmROlroMqCr8KdeB9w
DqXCKshkR3+kRUuO9fK3TF4aAKUrHlh/AaNh8tApembZszV61eyNnVvjejz597zl
qit8vw4FgJ30IPpXrYAZTE+ohWMFSEkOc3WDRkB+HIGlsesXE/uS0ZYGhKWuVlru
izCOO9icFT5tq36y04Q5Sa0nJ6YM+8GlfV1XkWJfwl2hobJ4HYrjejovmB+RkmdW
6HvmM+a/LZu4mBAkVZOHwJM7p6sFphSwTtR06Fq2NgpEUj2EFD8hch6V5BUyii7Q
UzF+Dr1XuAW4wdteIvl625PD1S4iwR5e0udO7kLtyNyFtbUkZITxwV59h+1I36aF
W6vlEfXVpaV4HbGZ0W+WXkIOtqQz7jUJQ1AJHpKCeXnYs+ZJ8AnfcTpSV4ZB8gm/
NKUfm3fItcKjLkBOWKLc5uhMvjw8jkN87JzlIm/CO75SKTIXCz30ItkdA2PjBA3/
1AnAw9xbPe0CAXLq5GxPjiVhklgC1IRatJ7vHwrv1In5ZDxpCSQvdOXMqp8iawGX
7xyQijw/N5GEu+2OJbDkIgHL7sDSKDn4noQPxZJmlGmfe2cC9BlhlECrAdvjzx/d
kacOGsXfjDCYkurYLRgMp9+YVkHVf+e+0LszRbL6QYhF/EC0YguttnUGhXGw56mW
Rxj46SGtcB4R6fue15wtMP2AnWCjYyejgztNeK8v+TpqokCmE2mhcispIN4o0xvR
EVKvPoK00walwE2tELxWB+/aStwQWcfXp7gzUIdoxuJ9ic0kIatxpocnOjt3xg39
LGSr0YtoaYeLzc/HddVBWrVhU/ZCllMBY8jSrzLiY0TRLgNgbiW5OvbVnw0VTbak
m49BwueKZpN4/oJQZYM37goafBZJAzAEkTNMDsBOOd4QA8q94vr0IQ0vdi9Feskm
Mqjx5C9IT4v8AuBVJxN2ZcZGZ91GgbJ8YDQ1suQo4UOFO/KXO2573OMFEdl5A0NR
1YJwwkSdxatmJX4MTg7X0umLTnALost+Oc4m3LydtOCm9ZsL4+nC1nBAE1121zsp
Gvi5OZ6OErSPdsMfvHumYHHNJmVLUPKGRPwKosmEZEd5diobQZsSyEIrqlrrfhxo
u1yi5Mt68Eo1OfHOgxs+CjVmnWLGQq0FwzUVFKV6JM5gPvo6U7GlNdoSjh8qDO3I
6hHeHVec70w3HDBarE029Bmyd/yYPs4cK5cFMky2r23Yyt6H2YKhSA6ORaZ1jqh1
k5NPUTXkyz7glrarmHUQmKc+B6adR33K2OW3cgaCvMcdDh9Fs1o5a40hfNkCMHEG
6PgvfKsOPCnY+oFcUJfC3CVnS2foQ5z8Rp7LZWsP45dF9FHUpAq6fsZZyIvgQzKn
b1ZdUsJULRbV5atd/sm/z6vUvza8xzLCwS4GWubBGKPxe6w6O5Gc8Bw20Zj55UOM
/UbvI969RjS17TALoVZ3s/z7E66lH2fxr+kpjYDig8RdnXaRQAObUlfUhxbOlL+w
+jTqXOa8fnUJz0ctH1YiMVLfuzwEefiP+Rei6ETnx2yTeNAxCcn95w7lPdkU9pQB
n3bqbbyWI1gjsR00ihL04G6JmYMQSF61vl8YFmEX7kYzHs1YJ6Tb+cS6FcE4FCKl
Nc7CpcrjF0UCrwVWtcA+oqbqFwb64k9Fwhr84w8LkYlnU+hpwCREV9QRDrlx8HU9
VwF+L+RAPtXJJI124ejlsATrVJYJ13J/XnR/wKzNjwH1tBJByx3T354Wq8bHKg0o
5NacZrVHnWvCh1rTqchBKgMhdynSi1YsH1ubnGLkD4e+sTU+0sPoGlM9bJZrzyEd
u2gKvTPKaXGaERlnZkAJSgOfKZmsQtAXxLzZ9vpYnxf+lpCyD4CB6LpcwBtXgk5T
Mk3znCqrDxTtcwDin7+aWUgXUPFXwk57jdHcWgzW81efYcs0KP0s+hTJsTIQ5IGU
tWxfhtjRLQ3N8+3p4zGI0AVslexZfGkuXb7/eSt4pdn+1iAVxktUEJw5QP4eLlIT
98HyvR6DOQsCu86P3dk1fSboY+Epu0yF5ihH0fqNecAyGOZYqHoR+SwSCh7RPdHs
dBzm7Aj/s9ZSTgLQPrZ9sm62MkRuDO1jppGsXTOMv24y71hH3So8lutSf/GN2nJQ
Orv8CJgpCO+Ycm/RIvzCs+xy/l+1zVV5redVNPI8lXub0LCH1XxwTnJ4pfrkxdpq
bSu9PYk6lK7+TXtV1yYr5wWaeMy5/GRBDGkxrKTVJHgKG1yzNjWM5ECgUa0lv0K2
4jjk1VLkHLl//3U+Gv7Z/CcxnG3l/QQylCJdeYH1+uGFHPliWQFBvK7vj/o4Zyty
atBX2qOxgXFnyRvFOlJtwlEb5Kdaz9h9mTz3GOVvh9XOnHtdrlXYP1IT2qgSd/wb
Xhl9hOJUSAj5c4gcZTGKEOxg9UAqa5pmXB1ZkX2raLkEGEyKdFRgL5N6jBe7sZOG
hfNZtOdhfCgtDZYhe5j05N13foLpAqmshzHXHK3sZsama04UAxMF5Nhv5g2KPKtu
SEYiVbwrQvYCGTxiCO/TyWxiNwG1CylR/ZuJvokFWsVdRYZWBXvkGJ15QnUYfdAt
8BU+i7pagKfsLcjL2KUcEjmmqHs9fSNZvAL1hWqkFQMAQh49NVYdIxibP0KdL33l
jILPnmkXiKOWUxCGWNRIZeuWwVQZr4/A6Cp2yyzNFf1YbEqeQ0i/rraWb9Jud2mS
SfVlky/Z4iRaZGDKwua0rya8n2rR88vGEinlky7JectjNgg2uxAprpLYS4BiqCGO
kya3vxC2dUq5ixFyAgVQkYOEvbshmnQEMKSVQl7An5fnfyskflOONB2Ew03zLAQq
q5EyCfGi7/+fzlg+0ZuqFsaQnOEePhZDNcGCuG9BKxVCfXNTEVZxh2gMLK+bkXCK
iushcU/C+9GB6JiV1m3NMIqdex7yr3IyN12EEj0IMSs+gYRRAbWQ/87Onx3wENuq
cnTN6NazDLFPIruaKRr+s9nd3GK8ZovcpmpCRtUhtaYvBg4MMzFn3RNi6RDU0CQv
+jE6nzYW/B3rpdbtdy6K2Dbra+X8llvoVhUgE0vLxHqbvA9gCqs3k+AkqoOlvNji
FGW++8b3UvcHLZXVYnv58gsrjX4l2bhJ3d1Z0xhGOCUSKRJp/h0pILUSzBFMbeZ2
uBKdA9eD7krsicb3pl5yJ+dxbegHCO6KwPNtoUxuPyMzS+sK57Lm9wA20SJtr6dg
pganG0DgcAyy7DOKl0L5yJldlC9Z+V8ixMcfcoB1B5jvywUB0d5CeS7Ld/tE0bOY
LJMiI/Ay8D2EkqrlULIuFc2BmuGtbgrCA4xZKV/WinMAUYwho++BpLcNS3tE25aa
aSFfPC1pJIF2i12D1bh3FcjET5ljJ6MpP1FpiXW09SV+3ZiFIfLhXqXgcRFHLB/8
CU4Ah/vv2AtoF9Kzyecu1zOh2osVDQSM5jE9GPvk/ktDVHmCIr1b8/TlUbb9x+EF
yDCknW2+ibsdd8wV2PtGOrUfJHUhwgPzi9B6aHVfv/5JKNRR4RMCFpypXWTV8UkI
PGF5oPvSGrOmqvv5u7qmGawgrGlofRRO5xNoXegEmYgGUdiDAnRQhgojHXgauXYT
xr5xegUFzroOzXSzCuzgGWlrxSIVOhHfkex/kmSpinF9umpLiltec0sznQ1RprLs
m44pc1HZu1cOKZ6FDm01PSRUTr2RHtGh1DlRyiytwNZMrt+zD39GwoTPvxhA/NvV
DuXl/XjS95SZ73uDXFzkcNlGsVvWxLZ7JGvsBpl7kyK56oR+HYbstlwSs7EeXkKd
MHYd7YVxqim0YGk3mivcOJb3B4uGeZweUSSMMzFUcgaqYvqr/q2uhxtVSTKTKGhr
zP+dzMCO5++/th7qq9UR2voS/5NIw7xp0ytxv9jWXTpVgowoc/aCA8S5iLiG8a7g
3Lfa+d6EG7pQVMkAHR/wQ3WjTMGHGTQy7zsrXxkXWRqqNQx9OBAQxjl/c8ag3MWa
edPLS1jInQ1RpNp+SPAEHtAxQPrJ4yynwXe+DUhq4IlE0MBDDnwvX6mdMgAhRT1x
pfQBtMZDYyUK5MBsQRTH9E+ouYB1GuEwQ0VM25S+zFndNDYucJnxnVWHUfLueZPl
G0ji1SgpHPmSpuFu+43fZBZy0oklvep6iaIuOVTuskr6tz2VVtSI5bkdSqhm9jlJ
Tj+kFvf3utj08guFPscWY0cgOleK9lHAZd4Jqt35hficU12MCP100SwnDBA/AXxf
60iggfjUzlK0/9I8C7Xrlzm+AdUh5XaXU1tjrJuIBpzzkHJ8EEubXcc8sGsZJF1V
4Fr7LQ8xwz8y9CSzYnuUVRTa4cflDunpwYjQ+6VKz3ItfG3pjpQVJxHyTNdMWa6Y
CdoczFO/234APzMgVmCoyOq06/uOaLR4WitUUfCMndKWJEShIM3YrGcNBAA6jwDW
3uNZFQTf1CPAcIo9uTCMikxtOddxQpafoFxs1Cokm0Q4wKWyz5hZhyc9GtiTYKXp
UFAvlqsneuTteeDhhKJ3ZXRS2Hns98frDeGAKT/L8Oztje4gfshPeHRafPJe5E7z
wJ2z+TfJzIDelJ26Z9jHP8STIan/uUp2FmudZxvpNRbCCMq1xkI00WXqwmAWlmod
7NVmHKNyJOlsJyRunIf/8rixP3xSAExPoJIX/lnas4WWxQOOyMLPzsdOak3sQYaC
t7iD02DCDUpYYPZZ33TFhM7AaIInOdmH4vy4u5alpuQerlniD/hB/jb7mpZ1HG7Q
TmGOQABYVDKwClQjiy/4tqtfZwlT5pKyYvqx7bG1+mH0TNpQL/1gQMYAgCIRTqM0
ZGJFvBfQ46oxidksU+t27mZyQso04XjaGLqMwG4qjRmpkqa1EJtA+JyGbX95+8yX
rgJQz81wf+GPER/PEXtonuc9V0Jg6Y0PF7yrNLHQIesD4E24/ssppxaKZ3BexMTK
HnFDbYcJcgCryq52xfdAPnK8wZt2ZKZSmpaVOcgM+p9VHWNZnE1ZC7vu6Wjs28ZX
sOnsHmdkLNnz3UQxbcd1kiaSkgPSaMs/+/7MDmg5HN89KR2qWxSgZ56Zanco5I43
TdNyIotNv4zuE041eSSl6qybtUveA3zZXYaVA4bUIAAepGKzBCWMuL6k7b4ksU1b
7fxkLV58W61nd/UMf+RkEaCKuASxLILbux6XkJMf17NvqstA45gAtfvYyNlC32vD
VZevm/E7/AOOdjPnvVALuLl2ereHFizc2+bMAgJsFxpYrL5EdlTbxicEcVfq7/Kp
zjAVF4mSPCVlJkFkyHZppHug06pMbYaXyhSqvmyGFFbCsx6/eYtr1j6GXuORpfpH
HB3gb2GfO2o7w7TY9aK5u7ND6rUWSFplycztzo43hy8UNbuui94NFS8czLVy/8nf
TitKdF5cEeH9eDz886jkqm538K7R9RVnuD5olssh6bScCKifMDYy3eFnLMiDHnoN
9KfrGnr7K98Qw7vqkE8viQ0mLllnqUBBikeZA5NOLNfqV3o8qlCBByW6BfpvWfrW
lOevgh6inZsZShGl6s8NI6r5og9H19vKQ940TCEW9LBvt8UXL1Iz0sn1EP+qPSaJ
IOEJO7WsVAdYeyjfS0XBGie40OKpisVYgv5v8eDOjTdkBjgpvr2XVxwGgiQLWAsE
GlwsYyHH+nOEqZon1SNAvOgDofLOS0/2AuqcoKCJH/6imLOX+qUgWBk+cXE8CvEh
47SYmR57BY4ksKeiyzR06vIUtM3gefFqOTT216DwyirhPfUWe0fMrNVERYLGzSHc
08J0Uf3x9DmijBOumTA9me7QwptXYZ2/x6FkdtseG0aEY21IiMshyn03MYNZ2Gyq
Jgq3PVeKe1cyXL/FrVIddgmsyWjzsquYCJQhKuAQeFKGgUe6vp7hUd6PjGyo/1eR
UNPZX3X9gg89+BUC1MMaYtPYXj4QQyavQKhu0b+LrDZU+gtkK55/Uq+bN9gvX0/n
DUz0o9+saVt7HzMhyUPgLr5Bw91nqNHSdr8LiaJFLLNa0pYeG5m8+YX3bwBLKTed
dqc/z22ZvooliIe/YAiHIJr0luHqHgT9baTHZVdDtQAyRizPIeNgjnk3mQpGp8a8
kAdoUUJxy7Dq0N6/0UhJnE5EVbY4kFhX0kiQaCQKBTeITvNEQPIKHEqLieznYKZm
zI7cXCIQD351m3rQxSeJJC8rgwLKe/YGSpEWpz02CacuXen0bUxy2IoUKdEJz1D0
AsXOToLQNqgFVm/089hRS7WIO6bYWRJ1fhcQxb8IHMqe5CSBLTr4q2XPO+d10gcE
jFQ01QI+wtD1Cncv3c8l6a78qltzcDUZ6cR9O6/NsWsoxqtUQdJ44bNKgY/texUD
MRLiEn3FqK7A8BC1dXk6w9IZi8e1veTHOSXKro44PVHeAm/JsibDKWY/0u8xs0F4
JEy4XlBUn6B1u+u7YxQ8Ge1UcNaF0DHk+48jXHzB3DndOslA9VztkbWRnctyvfBt
qwFiGG5gcQ3XRwAIncwCdhWSaptxH1pqqvSPUdq8vgwkkbDyauLxxOg0WG5tstqW
E2cd4jpHXU+uI9M1X0c0itgVlM+fz1a+LUGtKT2vks6lf8iXxDEB7fIMNWEOryUE
uGMoMs6M7Dc3q5yca0eUyiNqYdudUqGj/+CDzJ4sumTIaYQYWBfM+9pHXt8VTgRj
Md4aTVB51VN9CSGVDNRiUe6kob+d3l1ClQGqXHotCPSdsv8c5ezJtXEjV85Nnh3d
WjwYjO2k9r9yOx503717BVtCIR9wuTIba1bfJw8Kn/zcsR/rKU59Z39wZnSmlba2
jnswatk12aJ6zMIGQNRhb3TVzvHBtnI3fJh6g7s82N9Dthmua/2ObuP2uE8ddbVY
DfIhjdIMHAvIRl5d+IUPNP+64uC6/KiOboeg/y8+rH1oVJudaDbq3WZScXZg5p6I
oZeYSiEAaXvHVbTdwEM5HiO/jcfEmdK6hGIBrxvOWmmuBCYwGe29rKhoK6iZZ5+c
fAaOHU2T9nYRNvACTZBtvST5AYY6fVHTLKEmK2x3Za7Ui/nX/h1AgfzINns75qiP
mGE8fSh1Sq3RJ6xhurNbVIVmGALiWtI5rfqnVP91UCcffv1vah3X5NrwX9UbAQhI
2IOb00Iz64Xbe/aCYEmTMwQqyZD1FoSisa74YZuYHkJ71TdKfybNQB4Ih51hA3oK
lZuK0nUUbMvDnwgoaexJDF/3XKNwqaNkFZxpoQAkAHS0gCvY0plX0o7X17+BpKkU
A65MxexGIzsxkUmkEHjGcCvwx+2lJU63z5GuslJlXl07qNp4ngKQn1JpLnGshK8L
i40UrJV1r/TRENgDnbNLwILxvMIo4+Ex0njd7/ZedfJbl0tckbaCMa+PI1z+PQ8n
DCPQIasGxGQ4yU2oXra2lKe86Y61mtyvN+Y2EzgFbEJRTf7bgurxCytW/Ek1EAbE
e7mttaC6SGlKnpmBSHVQda5aMikzcCqLPyjniDN1yNpcH+PUsLze6aa3olIyvBPS
e8ZCnXKKq9zicFeIKpeuNi0qVMVjnqPvSx33hcDke4Ekc72S4Ov5Ugzpvtb3+hWI
Mx0ZICcQ8xEAZo/3JE3/nSSd4pZXNAlC/2L68BeaTrIDGx+Df05Hi2XmaXM8nULR
0LnE4top08DC3wCFn+kx/WEb2CI32V1ebTDzdcY0ic24Ft88RvKhJkUh+KJWTW0X
RARfBnIXYDdcWFumYAcy2sRhRsy3OawG2tjGCHhT3wbbXzzbu/EYNa4cR6LyU9l9
pkr9nhp87IN2mFQzqrr7fp+fFuV0vO1oRi2WoJbXtmhdZhSCxFLJKXzRRF2VQVgE
I6EvRUrmorpYWdMHXvfNUtZLKqY5ahG/x40f1FqPkwrusx8f1PiVuBC0NnDxlZ3/
W+mX64ldrenn14uGifwdUwxAAEdcFzUoZ/IVb1wV8adxffkHhIBLi2Mg6kXSfk5M
rKmBe6Tl+V1NBsYDvCvjDtkg/xadIGd3tIExUhgsm2anuwPrePW5WHHWkCwFSDvK
a1Cy7ur9zB385/r5NUS7qJ1H8Bh1+tDk0smDn9B0oOUF2CCZd3hH5kVFfH5jBxzu
3wn/fAMCshafZI1UIq5dQiU0kG/hrnG88cKl/6hWOywBAR3SlDRfvOv/heg949z5
+2D/pyrc8jdVl5OouAxLUKQVPYglu6e+fzul09BEx5xW+rp0THKsZUKhsIGogDnB
TOyiQvOAxIkM1yckTnGiBRv0p8+mmDJOGG49fo1neTWsloZegtSDMiOeghqbQGkN
QUJ/BzU/Qpr19VUzUG1H0ggt8c2FHQ21+0q1qXMOxCixSXlkkVxfNPY/yn3rgUUR
bp+SZqFpGRTEbpvTytJU9CZty/BIVGGDhnJwvPWxgEYJZjz++xnR8kprsdQFoZRl
7aEGWhbpnqYiAN/rccrg+wZ4pGQoC6hOQVhMJtXBwe42vmOPMHQKgo7UvlGqPq74
2VODXZDely7zanVH5nTikhc+J6Wk2zQ1Y/q3NYlj+NnOeGxBd4U4AZgnqHwL3tUI
9HU1Plm7eN/gMoyCzO+vf0nK588UrawNYo3J0mYl9dFDd4tcrXBEFJZRvRiSNuTq
q3pyG8OGd6o1W6dHdatTj9ueecjyCUGaTK0Q32KpnYoSUAsH9DRo08AMmMHV0kjZ
TLiXKRChac2j4sa7CmjY28dL8GJZAtElcpI1fdChwpDy/TNiVJa4skbAtyfQVuoI
rL74svLssLxnJJpDiRSIPLEPUMpv3Pl2kaoskfryUGxZX996a3WeCIPqA45ijAFb
Eu572gVbwWOtoOm6EPGLqcP1tlmMEi2bHm20RFZ6LUAfsDjgnIiORrrAsmutktj4
tryWIHsjLwlaghqfor5BTxETHSgPnDKyRuPFkLMKPva1GMcSdDXMoYvPfesokBph
f9PuyHhusgQBM1LYYUE1Y0LId2PQGJlBCEh3URsmTuYTjdbgu6EFtYZlLe3aKNwQ
OkyXWD/U0fE4m3amSdC18r7bU4bVHnqlmuZ8G6FNMmSY3tP4211l4GG83fMASmgF
OUMBN3WNRwHRMkly+tOMXdds/4NuVOoA5mAeUFAZzYOrxRVMjMJO4ZwH2TAnrxh5
kifn1aoNXPvIn4aLdUCkRaowohcyAKczsCAUevXsJpRdF6S65aeIHIQMY5X/Dr1C
jp3GL1SKmDAw1Hm96KScidVkFCQKPDbIDJx4uk/ond0bkihGVg/4cb60UApmSQ3g
dTzU0HTvBlzm1wC/kAk8zAdjZakYwc0ewJCiMYz8zNC4xL3KsR7051+uaHkF1u45
f6Z44ZEx8ey/ZJr6+VcQLbGCVdRGA2m3pHaUPhOoXWOwFYR8QAPB4k3nquK3bpXt
LLxFhjTD63vISm6iRBxdqazh0wH8pFwVDpTlcQFcMW2GHo9VTBR8aXl+ayB3lNgk
SQhr88nJbmJNGCpOQ6IGeD4KugyoUWWrkg08Z2xf4sNfdMLhvxd8xF2/ZW+eAQ4V
YnCxSuAMybmi7cLQgY70TrlQIHWf+lVnZLczbCXtsL0zb7/PBCs1Ys8EFtX+N8U1
JXPEDgcvyw732MPkJKVZvg5scySrqLer2Dg/JAdGEDcpmV9St4PRvscTYLcErp5Q
AzhifOoQyY3UEYxfPhNqGDIMPkCMopJiMQf6XxSCrbpyY297xilX4w8uGGINmN3D
VJhcjk6bIlSGfv03x0ztr6gritEXRMFT0waxBu+NpKMqn/9gmL/wFtuhwiOmKD3V
HE2MJKgAgQrGtCeyvWftAJihUK3yJ3TKwgqWH7Zmrdb9RfLsIOUHZgQ5smzFMW+B
1mefKgxu15IT+osrxmnEEZuYr47PhjFkGZY2jCfhKRDXTKhgt29T//Nzg2+A4zgi
c/0C98JvwqEtCxZheqRYLXokEL6GDLrSL08LlzCTQy9w9GBOZsgOVVEyPrgU1bDH
kEhL2d5nVVS1d/FfFigHbp2UBJx+IuYKM+xEDjJ96cvDS9BKZpnYYShkCPyNL4mH
utTqJstSRJE1+jrczsNp5WVbV6NtvIBRWu6xPKOMHCuY4OSmsIZmDDTt5fDoRPVx
nsQFudFR4RsonqJeEEu7cHTFIdnQ/xJrolIF3w9tUUtO6y6XRg2pLwVxJfAYFLxL
Pqn5t37BYln1IBo88VI+HPj+EuAW+Gjec+fZ3XSgIsrXoRkB0sIeUxtar7tGGEpt
M5dviX9jps1T4347F23PK8u7GK2sA3+PM0gOCYUHt39RqRgaWrtzyfeOru40vOLb
/KtRPzaI1QeKv3y8VESMNm+IHO9QSx5u9SND7LwaWZX8Nus3JF3QxrVs8/XjrbZk
H43WZ8UqBRvPQUXcAjq3S6iBVopvi9eu8qpFfSPD9G0AWU0EP7KtV+sQY9SMNv9Q
BuM3CKfkvqs+WGD6dzRAdKrwLQzhMvrBkI1hI3wyUZ7KkvnS9g3mDVh07NOB0r85
2mOFP3sGTeOkeTIUUMFHKFh3djc3+ppm6cq2AazO845+GIY9mz/sTK+4UA3QCWco
aGH8wjoGBe8YGOPeavR5VJXZTS1eXAYiI/HV6Qmx+FYJPJBTGY9DC7xLSH43uJ05
6QyQfiM1fnXimVJMRUK2912Z8x/mgYVwhhT8gpDR67CXTQC67A+iFCuiF0Q8AYpE
YFK7ayEqmTF5SVi5y2/X1gFK7LfubE2oOZKeVDw3aHpqz0DuGZ17Lj0HkYKtXxZi
z2kkETYanQmDvAXuYDYoGSHE/cFe36ZyzX3tlaNvxeMtcKvn0zlrEQwo3UhtXFa/
OSF9SZQcx8CutYwk3XsetwFsF9gox/3z8GjDtaC+SXzGU8YrIcDwX0cK4eNUbCQT
UYq++K9COhYMhg+7jSLGOA22e9ufR8oOTzduNAKzF6X+Z9Wxau6blzjZbLOcPCUq
6MJlxLZiFiItCTchpqNf/HNnzqgOhuN0NuJBKWwusAejweIk+nQK9Pt/PhWkir8u
lchZneIYZXnFNNnGwg4mNyAXTZ5f935OSnprj7bFv4qgah6ke42HmNTiiospSUbc
WhrMEwNu9O+I6C/ejJAa/UU25022urGaKC0IxmOpDn+npmBY3uZ2B1df7xhRzYKK
uxOIhwlTMhu0fZ2ZXLaWprc6cPR+wG1XqGdd8y7OC0DwqLuwNpxXQ5lET9weTWRF
NEggi8QD34bz58tCTMoxbO1Q47xtEzaeo+YA3qvLmRWOl7jEGFBCctig8XBVgzdt
/UY+EicH9Sk0yT2UmJkSHCp9n07P+2TR1a5o5giLkitHtlvuj8bXXHMDdPaNXKcJ
tgTi9dqmDjHwHNFEGChuuTtZRfZdOiR1I+2a2ZUdwvqYG515b9BS0SkqHkBU2UDf
zqI6tW/NxTgf+NDw0lJI6Ia10f0XLFyUhMwnDKj+0KRVXUMTp5EL5MkGNL3Kir8+
YvIZCHAfzwniYE04TJbl5fp/cs+V4L/ab/R3mdww5u2YU7TgycxbBdI42FRaveuc
KG+2EpCLAhj9TNQEBWXV8kNt6Tn+SD7OUf8eqWc5/g5cUJTCcn3hhQqKK27qbUmo
u6rMRCWKgeAsqUlebB5XKnB3oTCu00qYCqEUKR94DC4XoKzJM1QUmxBDIDsd1EKm
S2spxN1BeXiy+dsjs7QesIj1AudlvVIk7B22YiKrDx/whVWojjQXWieADg0YQ83Q
1odGvK7CrCIFcjJrhdDLyaM1KRzsh5QzrJd4jX6ta6MHBtvwwUZ9JS5pQ1Ip0tTa
gtx/x/4Ucyhov/v4U8MAFTxu192mcDHdtVeMyC0k7+n4d232FTkcxbdKdG3zNOtE
jPs5DaygbIbfFRBYEfr7kdy5Nxsm01aJBPoTWiVkACPOls/qPTk/LBSqMRgC0eCK
R/WRIYWOGMeBF6K27ZUBQQsJugV6ZHvBRcrdSZmt+bXg1+KVCCnqJ8i6bkN7CAoO
f0TugOqQmJnJpp7tyBayxKFE1pQq+pBZPt8rKGdg+A8BRsO3lTPC/SyH4i/wHhtE
Trh7x5ufANNXctVM2Z1VsRR9ZT/OWSMOIUPJ3E8ourxF1dAMmVMsgzYKQhFaGWuO
z2//t6GEDW0pi2/WzGne2NiitM9YgCHB/hLru/9umvVqMDaBPC44p+6KrPSmsckq
mwPoaR7jJfTPO9R3121tNTTtDw6ykYnR1L7Mkou5SfpcAabO/VDVH2yC7yfgVZHj
4jeGUq5zkLvVU1PK72cQTkWGA7yy6+TQeF+c8FipNw0D42M9mIfghY4ft1pYaoiz
TqoinRGd11HEWy/GZ2xpAff4vv8/XyE63tljXFlnpoVN8+kGWqN4X6L7K1sWx+Uj
gMj0RuXp3IWoeH5mCTnodKzZpNgrwqSTt1Lvq3lnH+ML4j7Aiogpc+CeZh+fszCM
FZ89ypzEpgyb/1w+bjm9IXnGc7/qbbCcnlCUQMC1qI+fmLrURusZFvX4ob23ZzUK
cT0vrW8SiK9q07Kp1a4kuFJrpOUuL5qC8P8UrP0QL2CmLGtpUSJQ/JCX//uWxgV9
PQNOy9WXwr4rrL7msTu4GCcxTkTg+ISlHNHkPFTn3bKnjzDH2YogWMb2jY6Yyyed
iT+utTAIx8iiZ1AEKsGdJ95T4qRnPcz9gAmb0uep3K87dHxe47KoxYJYbzE9Rt6y
Q4gZ+y6AAspo2w5lBxsoyV5NbR0YEJih9A7l5LusRW+q026/rLGwumrRRc766zr5
UD7cOWj/miVZlXgDKJTN6wSoH2sDhyjrqP9UWztfv7kGW9Pqtc0q/LLmFyEFAIW4
/ILXfR2fMKoZFMm2t+Kaz+gnf1p069r7nfxjWSGtxUptv/itlw9plyZJG88peORm
bJKkopSAYK3y3K8hsLq7rLqD6ANQ7lOxytw/E9on11R+SIqCx3JBjXxqc+R+8kiR
YFcI55EV3p8y6wUrSK/UR/IN0LmNEWkxsO1DxvLJJIDytNY/CiNNnOnczs46RBx+
xK94RMWhDWyasKwr60MupnjjBWsvNRQwx7R8Lw9tvDE8KQAU22LXwU4W/fT3AiMm
M7aU9vrV8iEnV8w8lgEgpNywZE6ZfWAwX2+UwnKFQrEXrD/ltztnV2u9HC0ORSXC
Havq6ERVsCv0Xf90Q0BQ0NbZHgFXmgjXCHGgXE13yD+0/lmxYEL7pxtJOme0KUYQ
WJXJCbKT6kUYD2cOF50C1+t9T8XpxCllrWJ6d856mJrSr8Yr65ugOBGEdo2b1te0
xU0e2yuxw1XRb4CmlroueOeeD6eP0xShUqW8SF63DtcqfWy4UZt65NtQYP6Nrxzt
qnit+tAe54vYp4sXmDL6T2FzWkVag+McHgKVZXqWHZW4Fl2y/NWpafOJA4CI/W32
uqr3xnFMJeE/V+/mA6Glj2YMW5aqk4Hbdmjg8A56+6ecRhDLTTOaXYzZjTTyx0zx
WllEpX9uYUikGhka/tO/GMEREwr1b64/GyFguZeLNbMENFbzi2sfDOzsNisJPMHZ
pt1fx0A6IfNloaCZZa+mFbYM6A7RtnqnTcN7vkIQu6ALe4L3BWmxQnmlLuEnrkRt
gQ6kLp5YuzwqP5UGTkIO52Vq4tIOerCgJ2k/i9MNb3qYGPapwWrHbpFvImEk9Bey
c5/SaTm2VbeUw3bmOHK2N7M15NnLD6brp2725k7ls2gBYA/VcYfgC04CQ8fzMfwb
X7qmi+a10bdsFbhvlWBSvTahORQ53SGc/ZTuXSiQu7odYBxIIQ25VxKJzNLJtayI
radPNPNvkmNXerKc6d55uZt1MFpIWveoD1h2i9sC1a9/nHm8Ru1g30SeUDIocDTS
lf0+1aTTrlk8k2bmOjZpyCEExIVr+qSCAlk5dayStoGcj/gqXxmsfQgGFprmRFZa
JL18ilosMum7q/O0fHfhzySqQGR0QnEEbfl4e6QSx9id7X/VnotAhqscoHxLNOz5
xEAk7TYNfc8xRMrvujcRYbTtvwFPuQ34UuvKu1lUeDfPe9bhkiQMl7/w6bD2yBnR
zSic3XAWC/cpM5n1Mb4l8KUEDfWQ2Jll2SzgH3zeNeFU9sBYm+gyMtzaxdKwC7PM
2Gk8j0AiAlhie5a1i6E2KbGtO1Mjo57mX23lg/BitUVnoy/strbHqRICBDUD0gAT
BqNLoDUyeKZcUZDkR2ozW64FFhZy/LoDz2w1DvXXBBn3KpC+oYMOqGYXwnFU3F9C
dBlfh0IfDbM6z9LE3/6wlzUrrj2XYZxUDctshNvNQAKCMts2bEF+Nkjm8IdWCdsX
kI6bthQmg78mpF57VTZ1aJBlH1F+Y/9uWbwBcwe06M2ucXwaf0272S6JJQExa3G4
PqdL2omIDPmDV/UQjckEUCRxS4auYAexvqFW1twmzVtxVVUkOn2+oGkCYhAOeXsx
Lm7o0X0/cxpVt7ZPge760Of6xwIxJ/MGJOKx5gsST1p8uri3jrcsZGNIiaFrFh3R
UAnbXe0sqcdMkcm+o2T+Y1kcSECd34mXId/gXj/DevVFXM4WemluAg+bs1KG67EP
I5Iv4hq3YxP6mgAjXI4lcGKlsNL26phiVoNqs2YS0RelmfP/FWAn7N9iKp2W1uJO
HtkXdNtax8aghfDZTgRG4W2v2f5Db3vOP4ZsCDLn6x7m66NbrXcXYp5uErgSh67D
kL27g3wkyI7GVEuO7lD/gr2LDkbabQxCdvNLzd5+uux/0ldQS4ifRe12owfAVNiD
3kOTO2ZNpxYnVzWoQ7F0+rojn7mVl9Lpw7ruymVLtBUGSoqVGw3Uf3XbMo8s9yKq
CLiSQcq97RVSZ0WlYoauIdZQUnsoMrpn+FXFYL8IlKo6OvOlxmAuMXL4g01pBjh7
KH0kwnzmW01lIXwJE346of2g2KvmyUsJ/disOac2hVsqSw/YPSbXdD7KKnjKaqaC
sXyz4bzVjZs2iu3Y3kLNtN5X9tQkIHi3gOLPS7jUoO+WsPfZB5VMunoPo8WkK2tD
nMxKOb2IIh75uL+FcUc9GkvfDUt8n5HkJUr5FnjfQA8uVr8NX5/9ThZdtae3J3jC
vmIZVauxFBWNTqzVaBhOvCTVbjlSUjTh1ZhSvP7bLeZV4b1nVgiJWGzO84ZTpzDN
l9lGtmK1inrS2zXqenJCiEivPO5J1lrbwx0Ls0/WFweBUbnWfet+MBCk0AyhrqaJ
r78EInf+hnhD1Q7cL4CPxgHcR9hwl8jaMT93n986nzCnFxcymFV7NqBXEyE0A/Oh
KrwgvY6x3FhkiR4adLYWhyzY/oGfAAPdPotc9WUu6UdlDGbfVbopgo45LHDKtMPc
u94RASlnZ+V5R5lE0TB1mPF0H8HJaMYWUZbuWIgrB7LMBNhjZGiG2BpdhI4lxiZW
jG823W1aN9fN4eYiBOkdDfM0PXuIjkytOmSbO5PtzwJD+1te+UesrtB9LRpk4Sqb
1XPDAniAhqzjxt7yBbEbbOmVHwm4ZoXlPKypikPCBjAgF64OfFhZDsJkqSSfP0lB
ADbebNHLlMdbfBhQ4NyMAxougLIOxcQQhswx/TrChTNx0UG9wvbmZtdyuarFOVqe
0nsusQGynjz0mKE70dLaomyFDtgilYMO/trYJ9txYH+O9ADZbhlh3bcRDNFvuKpZ
s3VdkGk7EEn0k6kYwUhAQNBUfGqJCeZRpSU2UiFOwPuZS1LpHSDRAEj0x4Fd5Da0
S2FfwfefP0ZjyDVGobUvGtyq7pyWkTGIihH+YxgvtRsRkQn2ta0sRRuMJ0m7jEhd
TsjMrLcN4peEBjjlZkFA9DMqVUViBj5rx1fFvw8QqRgmEYzU7nKhV65APeUnMu40
IaxBj2elksd8P7ik1U4GCCmwNyordNzpViwNhyehj/SMlWBNKEGphB9M2BX3+5lt
eDTwPLOewEyfsYGRKz/E1LIQtX9s+wDXtI/px3X5yu9vCS8JOnHSoZw+zDvdZNTb
YxNRgAd52DO+V6eBFPdLEKQhQ+wKxvaZpjG+sZyIFxGOC4gPRGxpcpI2YJTuOQDj
xPyzEnOsAtCcZMDYne2GrNPKkC3Ju3qjIlWvZ6aHNR233x6+5YKCSPkM00JC5ouM
VB3kpDAe510/lM5WCgfnKjf3VYNRBf17OCS/VV90vfCz5OngDqkWObOR4lXs454u
+zXeJhtLU6qqGkSZLGDahPtSB0NSQyok8cn5drt50dbbdXfxYpRbec6rxP6FdUJ5
1cCt5DMJAMa0JzOLxyDnDrLSqVnTZ8APDLbqYgHS25iie21ij9Nk98vUD49Ut6LN
16h5fZzRuoUOzV30VHFbh7QhajLFhzURRW4KhHo1WrEU+r75R2pa6/UxDd+/y+mp
HRKV+qFDuQDqoOF5SNtVd7lMvHzq4l0R26ZIzD9FGrk7WJUz+DiBy77zB86/vw2K
TNqHd+Kxl3trnWLu0V61kZuhRWGOcrpAy/BWZt2cTMx5cBLwPsvu/QUMTp2wZQ51
V3W+LWemFV9pX+5BnwCoFKhytKyETJQDpJPnSxpCcm0bb+LZRZ7ITDi1van+i/56
G/hNPTXhm5CPgZntNS3WygHe3co51wrCXPyNavDgF0fIytuWoLS1k1ahOW3a7sRy
JucaB/osGqZaQvz5NgJ/tEGBUXlaqB1g2r63VnOkmVnXpf273mtBdqW98CsjYbt4
5wrIzfrGk3+B1mv6bQcpOcksgwBLQvm8Bxz3vVgJPm3JYU/ExpMGTNJKdn2/4nQl
cauDbdxh68v8x2dM5sx6BDhEvFYTeX97WnJKISdpXw8QMXFclIwCwcuMHgIper6a
oO1iF1Q0RaCi0GdBvD8ZIM1vXuGEJ9syrfiVuEdB3nvYCFwCeFZsQOBnUDouzdFu
aPeCnZdgP+5VbZDq8uv8uxsooHLWdPBw37qhnaRzKAkM0g3W5V+iFDllhPN9qpJm
/mg/T2rTkHc+Dn2EgcPtxFydjmXbZ3uDoCUFDWoyHYYF0V1qvpYUwQRtpl4YfWrd
0/dYFty5dzI0+Gchx21p4eoDonRlKK2ucNjGeypCjOLWgx3cSYG4Wrtmwi0RgSrv
xlDrUHPRU7dhjYGGKJVpkQsuX/2u7sO6TlvThOiELMlF0aM1nURyT8fJ6ZkCcAhO
kRyyFMHkB2YqTFa2FUmARGg7U1tmwC4MIaRx7tHcXZELjJOWNDupitoJgHXGMi69
ftq0FkjI4g23mWKtGPDxsSbJFJOFuVJF3avruxWf90R+Y4r8ksAC+nDYJAXvXXvG
r5ecPcS/KSmItyXtSq7+iCBh4vCuWsO0dGO7pkhW6ntuwDacpTOAUYxSXv9dxQd+
CDbcIgJjnUQyZx0WdCBihl2jYk8xa8a8Fhl6qTUBzqktyznrT/XUOoydl665lrqy
+wi2CtjRtLNku2GJJ6UewzlRbBmoCfAdGTrDCR8s1UOqJQujlCza8cJ5StAlV46P
zBn2psFssyf/EpBnsErzFpJYy6oqvSBdvPtNi6O2ql20m6n8X+JwFHvDnJD3X3mX
CSRPcesJ12RmjF1F7+r1DgBVK5yGeNJwvtF8eE/Z1AP5OuAoVZ9MDmWKH7mNtWkl
k9y3cnzsUoioosI/qmzyfjjAvlVeOeYaAe4kjM3MrpKlpo9MuJAa/9JkduIEV4zF
smUieHsz6iSmYvAzIdmLqyXghCHjsOc8RuKLXB6EObGKjGJ5GtqkYVcQAV3qjdEc
piaxed8jw6Cv3iHT7EKnlQWRC4oK7GeallxHzMEXxnYWMlVffkHs1G8xWudcrXnv
RAHbjNPZmGkKFrUf4pfZ6bzrGux5MSK8NyxzI1zmpGxaG0iVP8k03TM/aLqBDGmw
UgYfF36BJIriCsRUQmf5h9Ow0OnecB00jbAtGfP7YFDQ0SvBCVda3qGFdhHzPtT1
d8jAhbRteej7UWyMZZIx49gX3Nen04riW+A8dMFVrF1JWxUzkF7q7cnpJA/KpIvS
VCATpx4SAYXBk3r4xVUdEJUKXMiAvQXjZ2biUP73sxa62wntCYf9wfzu+l74eQAj
gYK94A9apVbU7r6sUIj4kM/k7Gag9Vw3siQDN7m1wejzsF5OZUiECtnzAu/JavNk
6LUSRVVGxZaQ6JZPou43rCMcILjb60FXQ0tXTEui00Ex8KuDOI/SyqyM7LLc/Gwj
hkEfHrJ8drt7nC6nlmLwx4pKnzuUZgNKcicAcNsNO7R1ZBrYfUBySJ2sRq3gjm31
xnfh4NgBWIsTLaB5FW2uTsZ4G29qZ4uvRDv51twwgKpKL0BGzjbxytXMo+3UnEa/
SmYcpwdJHBlsLImFwniJwgFqztSmJsERmssIKPxZMt9shbXctKPrw2MxubQTGHQn
28OLw/im2eLoretG8glH6qs6IMUaqgvvoigbe52BZzZAw+naEK58GK/Yvw1ciEgI
o/UdGtonTxa+vpUoZ2LIz4M2ylloLaOHvr6pxD/7R4OdKSQiLkV9dMpoK+6o+eob
BNZ7CVv8htwkvcFRgJgWyfI3Z5STlDyVq+wu4ZcYY6hNSqmmRaLaH8bG3IdTacit
WFETD1XRAWMLYeSyd0J0wdLgsDZjQBt9H+62QTVZn6IFQjeV/v6JVFkueYAD8bhP
0EXkmq6iEtdVV0XLY9LMU72NsCvx8qxBtsp8JLRqKLTSjtUoxrcQHNrSE2LHpALF
Sv2ao7TKa24ur+jJ3hPVU6FHTGuKu/a0559/S8tIWV7eg6/chZyw9z7ryBZRDtrS
VmsJBRt7MU4d1AQKbrZU2Sqd7hJxh4WSq3Ubn1BJDMb3wjFdc3usdwAu5uDns3Cw
mKLlIVYY70Ne7Gx0GCf1GHurnU5ZcotesnBsBgvM8TxnTgdZNNGh7sx0YyAWFjtN
mUWWuMvRZKEY7bHmF01ed922/rbyunGHOwHrxHw0aS14CllhR4U5Y8DE7+2EsS2N
od2LTcR8fgL3aMMGqhExD1EL55te9ozhZw8/xe+FIUImMkFik0mmNZpYZylEl+rK
HEkiRQGbLXmTJK4yykbNC29c3qe2avsavdgjWOWIyTJ5HIdyoeiVHDl9ACvO9rev
dNd3Eg4Fk0y7hreKzwbbVq1J6BW6xWwa7QRNPLRLYH1wWY0lfeB1KMCKFQ/ZIy+L
x1SmX03kCIt4LFmWrZBScshBT79HMFfbUmJ5iyczbwPBQCDPhdYiR1vnMjBt4kY8
I0Zu+rLHPrSKAdIaFAeP7fap8EAjlkVwCp7gGpHr8qQJzfVB++FXSXd6Lav3CX1c
iuexg8pjzFWZazG/HnKTW7fhaVbnUy3QEH+3+1DDqU/eQcXJGpGdRcPN3QW0GrB5
4gZQVHzleWZPvEgd90mm2Qk/8HlrUDY3R9MiHLKqCVD/7yLPNYesV8Idlvoymo+a
t5a9RqF11xw5VByaP8gixkx2hyXm2W/1H3QfMaRUvGBxNCJGVO9kDakw6QeVoa1l
pPUWf0Vn56KVnA87zsUlk5+3ik0N+QxPQoUJc4mhF9rykEAXIQujthVeKbuDdbJY
30SHm+gIfRZ7PcutWzFxoyfZhZ++2uOHc5pCiZGS6mITIWqYXIz5aKMviEKE/mRI
jYCXFiH78fIuhkNEvutGs4UqqlUd+XS+lfyFUEY7tjHCNKkgAooEW6F+hXu+L1QY
c4pUUchHS91fBlb5YWt44FzI3GkoVg2YJ5pJiakiOpUTZhFcs1HAnwsGcBLjHMAm
vHu0mMeMKq2XflC95DJNKHA7gN4JFFf19gLN37d/BfyZ4a4/5wkkRWp+kqeJC8vV
3nhk/wwDfQvOw3JBV0iV5vXI1PnUbobdfhRt0IF3W5BZyoWHk5TZqaL2DJZuhrNA
kFXwjmFYVBgUiC6V2Ggx+hBd7ynYNP+OhF2vxtIcudzM2HcO8oFFUvIXTbVUfVT1
VmjbCIuFacz8cmzm2OuxULjKMYBXLO47DvaNa1aVHiVxZBcJO9cByDy+M/MUPmgr
4IrZt7sPbJuKiaclrip+I4vzE1wE/KzdfWKd3Ers6emCALPeOoI2U3JiTgRJhnlr
6udSvHxXOnqvn17eI4tC2nQYMIeXNGuhyIvk70NNE3a5OQvGpvcoRVYkEHhCLpIs
VvpsAJ2qwvKiqQ3nf1l+09hbwrMI0QExaLlSb6wk2ZFWmHMtZoEA1/dN0GQ4779Q
nGewxH/spiudr67hm9Sw91moN2Mp3od15FHPKLBufpddhsdwpnVMJvqUXnYQ2+IR
0/AIzPxeHVkpnPVXfWraQRu85OH1pEQDFO08KNMGn6kjbRO27amyshcIcNGUOmy/
qt1G7OU4h93uFJvyl2IvGISRFyLtMkoTS+8NC4eGsVHLQUYVejDDmaQp7YodU4Cd
5PnYfRT9Y6oT3vH1zaJTFLkfGYMDt5V8RCM3aedJeKBSVNy0WFUHcIWKYzKQtgHQ
FX4FpF4LlzouDoeoBlgdmtKxTPYmJwxMUfMWgGTskhfz1i2nUEX/QYbyRRmceAPo
TDPicrCC/JMVag8yDSsDDAH42Pnc37J5H00bkaQGs/VyXMH2x95K0CTBvdLHzcNV
zU+lLO4juvzCn6eAg2Rv5/WuKdc76crOPgsInis5oD/AbNPXbxKy08M+ZFHvLSdJ
n1FBgV0KErpNP7UENcqF0kpaUfNCoWOlG75+GtpRYfFkY7FNHWF1c2BrUWkYdVfz
X8w52u3uwBlJisI08NpXgzj8LDzi7zVr2CLcN/4lnOfiivMq0Vbhfp7jnJ+qf7O3
orza/7+p2XSofE3eCpg/h/bgAoKa+u3Q5+Y6FKhw/FShZ2NUuxVWbMG41IGjBRlZ
RDJJYyFvTtDBEueCy4TK+ZSqMA/gqeMC4lceg8257Vc65Xo8kk+VDtlvjdsD4jTy
6pjZydFwNBiNHUDTOa9XO7+1RQmnqYn3V324okrug4tExeA/XaR7GDwzTWMKPP9N
LcansOIbg0JU+vP3dHe7/V2VjRDqyJYLCk7wXf1Zwkp3lmeEp8QxDE1KUWKmHd6D
cwElVDLcxPA3eQx2501vtLO/Ffb3Q8g8UwtEWcsrN69WsG7iJ/zg+gkaW2zGXmtd
Tn6gw+io+8lMEesbyy9EVaMQjMlQ+Ehx8ar8LYkRIDCJhp9jvQckIersp9ZzTcjq
yU8kQJoPw8VHgmhVJP45nLHwVd08FztZTQo060L5EDJ+hm/9mDDrsdsjy2If7uNV
buUO1sf5ELlBIOmcDBLchOJtbM+oeWMvyrWmwI//UmDvCyw/4grx+Syc+SoeSuUV
OTd8Mco1H51cIlGr8qzzOHZLJ3VkM/LYHqht/rSA0WxuqTHMR1gHO6R8dZLCPFt2
ZgXD6GlV9E6gVfFpIUd7AkYmQRr9j5pdSWQjZGNptTFbrkakxkY3pTMK/0mDX87X
VeKauO9jFUPLHHsgOuNoSX8G4DO0g1nsqcmMEAiD84FBq8NCheR9+/TDWevWOCBX
IaCQWNuSigUK2mPWUGjQo/zqYep15lw7vZvp+XUEM/j98U7Iwyj47tt+Tq3Hq7G9
GdyXTrpvM2RXbKQwFDus3nzxxc6mThKUr8/5d/XPcOFnlB7WcwgU+jynyJ0HwA9e
+UjRzL4Hcx/B3WyQyv7H73dwjIsecG/4DbWtWeVMziiXnP4GdEI5UTp07kq2zzF6
IloohkiyEq9kDseIfm5e3O1xCd22sU6GFC8Wo9S1O7BwE1nWXufDOoAyLbusP/H/
u1LQEPoff5GLasl2fBZ65pptHNJLlG4nMk1BJU/yOzxZbMeo28q9dxvXsXVh9kbV
H/ad+LSFsxucsWSXRWpNQs6JTzspqfzk42d5b1HCHlg3P7+cSx4qTfK+JIgnYVQO
4t14I1yv2h0UAFnm2MnhAgVqxBjcAy6E8twsrnZnz7JYjg/sxYZ6sRX85xBDTjZ4
G64vOoOYQrDhmDHTFFGaK2CLnBk0/CWdgw7LsAom3VxnmF8Bg4yxXyPDWETqwZOK
gBsF3EjAtD0Ncj7u/xMFs271ccA+Df7mj4/kusBd48VhndOTudAhW5e6jWQVV/GI
GymYH8D+Z9ZBL3Qyfqk3yKWs+lCAk6KwH3g7TU+kKzZ/hMxsJQkBl0QXa/VSuwQC
4NgqnoTBHMCjeJUTV1GSRKkEQ/HwKs/UmrzRNwzaFqym3y/H3rSBxtfszy6uNOMT
h+auukLEUH/QC1+E3LSz6Dp4F+f5s4dT6LIqztyeQgRGyHa8OQs9LZ6cqe+4ea7C
9I2L5vCdoxK9z0V4ZVMfgDuAVprF1XPxXF8RSzy253vj73iaNamRtR+/U9X7FjAc
CVN79gZL+2u9oiXTs+vbWKX4Mn9rtaY+3EsCDaAr6uHpKni8IiwrnrtDOoYxfmRa
KvvOeGpwFF5hjJjhHncg5Pf9KM58tRlMBz6pUNre4Zx1E2IEvz47CpJyLBVxAxar
4FiDrs0OKCl+i0liCK8SBQbo/CQ7qjlHAxChIsbNSQfTkBjS+Jg/ThA3xO/Ze02g
Nj3AXymc2V6y8anVZc1qhfs/FjjNCqQcnZDrq5iW7iCg3pD/OCORMnSA3LL94MW7
PoKXcbaNlEBuCIGq7WB0eQKUUuY3gEkO1pMFidHSIRy3TVT8dJF7kqY5q0qHhvIY
q5KUlHECHgncG8qwpA8Li9UnZVgR05WRpe7PwB2OYfMG7rG57z6/YYl3rIP41A4P
XoYxY5UQ/X+wgIEwWM9uTXKinS02VmfF+TVjDNGY9vEZcGRXXs8ZRsWl4yledfMo
IZ6uKhRU3rRioqUhb3xWQOuw/Otbd6TLENwWDS+YW/37d/4da0IwSNITGuPM81sY
ajTeHifvGb8MBTlq5tMPoRV4X2q+ssDg5A8bdK7p0e1Xhly/QP8HZhipRpHivPJL
W5yMZVGOukdFYdOGLhGsAVjdkNUF16aMWS4ZVIddMmwaB6nWxLZwYWyz5HXP9hef
NAulJ939kKbMdnYfjpzZoPk7St17k3Qf3l93XiS2Spc96k6f7TXutVUraRN98TPb
Hc9AlPNDTzieBVzjJm3LhJVTKK/eDFE1iJC6qKXm8Umot4aNum6wvmmuBh+HInnF
rVP6rU0STYN0KwrmsyuEv0M4UYAPlLpueaVWdGJF2JJ6Nj+Mz/lcf/nzEB6cG5oh
JCalhoiYoRTTNBIIDCqitgFCPaKvNLxXavnq37jG60M3GM/7H4DSA6/e9NdLH0uo
mId6IHwphXt0n782EWV96fmDDRVSKmAygX7wcZ0xsVVAmy6C40N9rgThx1o42kG1
N7wi0LJKV5NDbUDyCHkJmT3qhnElOzIBxkikFJC4uA6W7El7DXVBaJSCZbdMIfyn
KzWkXvznc4GxgxuDi8ipieFMC7v6aZvfQUxeyDWdjGKVBfakVDfLAj/w+Zdh5XnS
IATrvJZwYwvevH7YOfO7D7682IfucKu1hx+7+7K3bjNj3dPIsy15/rhzCNkXGfzW
jrLHwEP1bDNSC1Co4CNyTza6nOvcDlVWp5y/g2eLn0Qu2OiZ6PiKBk3YhASX1aIp
a/aoBmhO8aIB4lU02yrzMrE8Xd+PhiSAUh2oBJqnZtg592HXzk3QqtT8PYTFgUY9
vgJYSZZTSoVml67PRUZ7HmygbZkc38F5dSG8Yc3JAI5wEWYpp9fQNREQfNAVbAIa
Rt8dPhZeok+Vl8IOPGuQCmp38GFPcZl1JvPR5I6p0VkHE/3s9VVwti/1g9lC1Jbd
aQH6wqeQ0Qwabjg4QMw4H2vJmAcRPNWUc9AXrabpyvZRIQv4LE9gLLPL/DsKW5C5
3FO2QC5ZQKntdoMTc5oVGrt/6H1ntunpgg+R+OD3pg47598k02zM0lwUHFpSZWWk
0uHvgrVFcicqB3mrh0kJGUNQQ+iXqoOnyrr6+t46qU/dRPOUYqUgCcUl7YogtOud
IcklhJNmN9TDq9CJkVTOERB/0Uw5F59ibQbeEd99kRrtBbopCAyrdPb7ubjG6gxb
Z+EObdPEFM2e+hKghisw+Ex0UkfmqKi+z/pBgjJsRImMptzTi/KuKnZROGe4Heky
Gspk3k8ZfDyQA5aO6oVCfU5mdjT2Foy6OP3bGO6+0HE41r09tnuRNV2aYZerL6zg
ovx+ZuD/swH3+PIoF3syzxI3rg1xBvmkVqtmSFiUd401AmVwPwitc6SOhDV5WG9V
HFJYRU5bmi80KKJQSIldARWycemupqAuTnKSw495PHaSyo5ftq5nzUp47cQCHUWE
cpdSeNmSa0N+oguatd7emRd2jrZo+Zzf43NBrRPBHo0XR+UaD4PbW0/V9imoyr7H
5v3NouikNyG5Hk4Cg73xekunQ+a327qwAUTIIej7ef4+2n/iZpfsjCNb24x7sx95
rVL2OZOWbIFbv58JTK/YcMskRniZqb3bAqOW5FWYYULqdhAUUofnVfnNuDaAb7R8
qhQYUXUGuXIUfNYmCHopg/kk08p3Nw5TM5eEfPCX++/qK8FuzcvU232xdVmuz3Xy
WrTBms2G8FwSIhOUuBdoWlqbS0yOYnUDRcZHVjIBAIAEFBAOlZzvQWOxbpGwQH7S
rwtq2JwiYhi68hZJPYPbZUX06LUlr7nmxK+8rDB08I1V7viAbeN93+ON8pV5UyeU
pgDZ0DcI2OdK/+uZ+9YBTIcQeMB8SVm5dPdBaPVimNRICvvLxOtiT05HF6Jqog8Y
dc9vHlv/VvxbfbOQzQP9jelXpScrYCsFgXziqzzSetD1rZIgIejtJsnX4y5zlTul
soh4xYAUQK6EkJ29N6Fgkqt9qhUbMmLo9zihBZNsSPUTepIPJ4xKt+KoY23fkW4M
CvFpKFU/t36ef0vKaerlsgE/vUnDj1hzwG23CFzzKkQPCoRHmeaIGhhYAoFRRIi8
qKmcqn3AvCA569N+hMY2eTzwswI8L0PptbcnLh4YvyAM6xpCjd4AIglGOcNRZfRV
Mvut2rK7TXsGJXPAZv28Ytv3xxH9gp2GiDmByhjDB6pRVpNLzIMo0kOXJ+I6H4nu
2nc+okcFKh1blNXSQ5XGFcbEP07q6kVQItgFfZ0lYbBh7GmTI/PoxJvtnVZlT1So
G48TlQJJIgDXSrdXzpWWqa196pDYvAGnXhG2q/TJojOyq3nufnBC16zRJi9Au02c
nWXvw1VvKes+uPSKyJ8HwSzolWrnWNWdSe8S0l4Ak+h4UE2aL0Fat1x+YONWwSN5
CrfMKDo0gg/XmZ92ElpZFz6OpuFuliHF7t9wdLnFZMtbOLu8ff56bxwV47J1hrMO
j/ywsSUdD24d28IU9XyrNCQwpYZK0wEzgBqbi7UBbQdk2FFDisGqCrOBnRmPNT91
bi5id16UFKs45DWaO3HMqSzUJ2dr04q+4wOct6GFIi6Q9vskMsXVNK/V8G6WGgjc
oxus4dThPkajWHn7Olbi0iXwQMOeO6JRscTQVfmqL6tvqlwp9h54hxshH+3k8Og9
JsPAA7sjZxX5YZuQrPfv6obVLfbCGby93EY+5c29S7NCXV8DtdMse01jj9MNxBZF
C2aFnuWo+N82OPkLNyS16ybsS8o3uY9prPyVRZA0p2ZQWeIz4EIp0Nwj5+ZML2mj
77BbnR0xmzMnNQDkkUADWlXTNdhTyVbrHq3YAA+tzRHqYYV5G0DgRgkdoDV8MKsb
8UzLgMs8gqtJLiG38Ez3ZC35TQKGp01nXPXwhwIXX+y0EYnzm413nIh45jQhUIj+
8UK3pz7z+b4S2m3p3JbLeIrmXTdngiIYDfEEqWvpF0L6dlPI2knDwWfgmm8VTcpJ
DmkG7zpOi86Mlz9cWpYOkySMgrrguqkOt8eRxyDXVXRgBs9NXtq41MEVIX+aj0M4
fOSTUL4k+QANsHyR1rg9/xNqnSMEYdl8LfzxD44if8fr+JFriCdxwsp9z+JQtPCb
sXeya5058ovs+g+K/79UscoUxDqsbH84Zpf/UyUQ2geOTpyDumpuCIDyJcZMJeS/
fLK9vW2uatpD96kVEaXbIAuvaFGth5g2zgbV3/1CMpxDzYpbPf0Ga3tpuoFofTPy
SPor3o5KMFEcrPNsI+KSD+BltQ8UaN4rhWjW/0RLpl8mym6AAvgFQeLC+t/cGKib
kEkM4YwOElleC57JRQVb9GfkKF4MpZ/1nCNZdUcKh33DFf+Iicwt4uJFOv/mZ+8e
CXNoYTOafPFY4iIwtEcRSdySaObcYzEPzDIDJpCeGFr6Vxndpohvryy6W44FqJ9x
YEwkN9qAzT2VC9KOofmST1bgYI9GwWALEzZ9Hbsej7R7OgZzniZC1ok6wyXHNLdC
txk6HfaB3pkxVMOLDAWYA81Oy1rTH97X9R5zqeYRpIiA7fVmsJ4VbXsIUV5hONzW
pN1yJkIdsZMs6EY3oDPV09/1dhGGwEQ9PHZfUeLjvwkGcPrj/orILa3Ss29IyLLL
6y8fvVFZ0HzVxlvTtkdJWXJ6P2MMYipl5gzIrypqXNkgZvQrNxlfsVeQ9vitESEr
ORuZbgDvOUe1kHRRdMimSmXSOc4uQtxryTKoSwKSbIZUIjWgdjzB0HuoEU7qO8i+
Qi2dNO9igWZhX6cw2eBC/+7q/CIyZw1E3AtS2c2y7+T7WXcmT0r0bNm41tVzRqv/
DDOP21gzWvRT9jRcnjEI7+ibQGO5PXo7/rQl9TBNXChrP2AR6gtWqDBmz6aj110P
lWhTImTY7K3thDb6YXnMYJcwETXoyiB07AYR/exAvlnNyUa9vLfwpQXpNJJIJsF5
OpYd6WjchVn+SCcldNaVcrovFZ8YqAjbFJBbZcjsXkCShzLBhCsGLgK3gT/LetfU
GNZ0FFZDlIeTsXWS/DFwNEVXbjaN3LC0aCoFX2Kk/nVyIo/HIs8IB20sL4Acp0fK
xpUxNJv8i4b4a0LbnNOgP5JuJbB7F7l8/X1inC6+BMKi4xeRrhJoF/WxBXY+gZSI
/yMVaujcwaEKcEVYh/gKmhwlhFm2uO3Al4PicrpKusvR1JYcqaa0YnO3jGyGjtSr
rJUD9/BNDLkHfQskNEICLL5iunycye0ySarYUilCyzVTXStft/AC94g0CuTMTevr
MsBCctTSUwS5BLQg+qInLbjIyNGNU9ONZ5x80D5ov9fp18h0UPp552zQ7ZDtUFWn
D7jnUrGEkwiu3CL0Bv/Vo6utu5ssV7Er9bdoP7EzaCvAfCcNcF7rM9OFYMmWI865
FXpD6SoUTNjFUjNvvw6Q5/ztQrAF5GHugvRaWyV+/pQ86cmj1RptgEjeDuy/VVaX
pM8cDsuIpFiqkm9UBlSatpeI5g1W92BIPKNmYtI93EB8Stxyi4oFixHNch2JUdvf
V1Zd+C+ubOXNStceoVeFgXZgyykkC/0DljP6FJE9zq7Wu3RsKTOjU5vJK3Um2pMt
tIAM+zEZH0KmqD2M/VKXkpXwI3NF3PgsQcOvxS6IaqXgD+je/OKXAS3shjqj2reJ
uuTdVtrrzP3wXzSz6UofOjKfrm3kawOtgHMdhzMMQZ9DghSjI70/kY0mfjdsEpWf
mIJkVJa8k7J6nTtb64XEg6z51fdxTLX+1c7dbENQ/+Qud+jcLkatnAgSqSljOdDN
MMPsthjO7O8K2QaeIa1Z6b11KHl3d8OtHFdkPY2jJmyB8cYGzYAmEEJRdAu4OP+Q
3BZJY8DmW8xp4w1grLCpJ/Qikl7tcjRUWSiA71FxGwTF1vdmyDTwflgft31knGYS
U4ctsZomlhjAhw1HJqWe5CHmyB9vGYB3Y2Bdo47zKsIlpl2rVxTOMHef9bB+j1R9
PlcUvwKsvK9P/Vl+B3/m8OBsp0eLTHSebARTeiaQwYeFQvTK8VrWcT9gfTfzgEsD
R2UMRgTYXwBtDLyUGtmW1jZDF22WO1xHIOXKCc8PK+bD42+cN93KkWnvhAPlg+44
4qo8EGFgASKVuM8/XlDutnosLS8eA/Yf6ugyjmIJ9o9bzd5itdCag4rgjLwPcd2Z
Ybmg/ZmJbNYN3S6LaSPCoQHbmZL2AfKj6UY0/rdKWdNxPATazkku+4gkHIm6Tr4q
RhCt2JUSvrRbZq/C+MLxlq1TzS0JAokECZiLHh2Hldz2pBdavj7QiW0b5w2ybK7z
ATm8MryCWGhn7ul7J+jILlV4NxUwQkPw9gz68YNIbHKEMc9u5hZ7snAku+hZH76l
ozIpA0R/5h+7uVnROaO6bybBNv2MVRuLOO3aRf6/bEX/4lmEa7jSaRrCuRHw3YyU
i0jpXKtoRAcNbti//Qmooa2v4T6Kw4vf3wDaRhRk4ssGg4EIo1RuuBgwkVMQOSz1
nbPCiqh/axB8CTnFBVbqtaBUvhHqIqj9XzUoCvSSdbaEMWPfl9baMzk/r2jMvvd/
ixJEbfPQv3c8kuFuYP/TJExQGQaBw90r/Knu1VDAm1O6yrE41zSTuYuU1+sm8BKM
ycYLHWTVjhWIzkguytpl8sQQVN/wPW2KVOO+n+B05gCuD3j9GXNgtsQXiCgeoxsm
H3m87+f7jPHilpNVdnqnhex94WZY4TYNVAKddAcWVoPGelpRCgpezUdWmKWGv9Ba
Y4CJWTruF1aKDdGg5CD7WiP8KE+Xj/XDDlbSV2aXQHIU2PlHhnmqWAZWnYSWA3zh
8UDXupT7ju//ShrrWqe2BF/pD3MtGA807eup8zGDi/nWKh2eQEPpfbx/1r65FooS
Di61j1LgbyGVz3knagL9PcE+SXD8NKi06d/SteI+WRLdSrfha/7vqGS8OqQQ0rS3
qip4WFPjF1D7DcQPeb6V+sTXgGTyyIUbkZ5dCj0U9buAWk35TAC1AHG15qIT1q1v
r/IrXBlnjh0p0OLrfHLQJPfK7rAZd9OpClv66T8ULCq0SQbLfW5kCgz+ntFNfQYu
6YDIPkBgFgGVpyWmoZnhRTmGs/MFDu1L77A2mpqiAmLdrSGaoK/NwMPpWdu36Qsm
MYHB4uqO6EtCXYSfogxbV3cheZv774lOhwB2IqY+dLA+Ak4CsrMNxj5mNqRP3uvd
Q2ON5uJtqG4TXJah7z8gQZ7mgY07nvsltldLSPKo3gccXVq9phktc8c1MCoBHdNp
Qxi2z7EzIOp5YZLcTciPcs+Wo3E+piwjZsdhC55qbM57UrzcDWVFwyOf2Lsgt9Ze
OVWtTi9v3BCb6BuORaal2Vi1c+9DD/dp3+J7lcvrxS7c4Glv7cm5uJf4P8tBZEQS
4EKFk8p6pDQCNPSxX8Ok5h7yQ17cFbnxX5Iqm7jM0U5Y5uKriRYOqNN6eRihtsul
Taif9J3O5IclxuD9TXaIo3CiZLKLpLgQuCZ6PnX9nom8ny60zOajSwLDbo9mRnFP
sCcg0U1pk2PTrgaPFwyC673HIV5YmKxhr8THksQUr40GYXTF+fztseQQvs06Lx3v
my1M8dG3irRCMI5/vK2JwgQbIXX69UH4v86eoByfbauzTVIrN1LisXhU07jOk9DR
GYcskILYv+yTV4sdQHfxSiR3LmQnFmd59ceoO5SlmTgiSvY6i6kJ8/IONv3wboZa
Or1fQet8vYvbilArnYQcVRUgR0tnHAm1PrQxsS7rRTGNk8iJcWVc4GRFT6nu8wv+
Lk5jwFDgT5+ncn7viQ+/k6E10UkGtqYU9RzOkLdwhpEKqklaN0FufOrDn84ikV3Y
jZu7vY0xom1S9oL41gYObSOBjL/9FlOg3TPRrut6tu70MVam5MMpyDckSw3zyEge
hiJ2CJK6UQf8PBKrf3m6xggjfT+MANUBSoytBrY6J4KoB9qBu4RfTkkEvLt1x2PI
rVPwXR8O3d61BsK+COOs3ikB375tWmIhjhi0yugEIHtxl0AUDZnnCWY9M1/y4IBd
Wxqux/fS2lXS8dad2QoTHpguyx7sf6a5mKiERUmY48Fk8MV9iqqyIPqUTbN2uOUe
2DkYlDL/CpAp03d/CtKxhaGcZiigdmhxUgMSTb4LAAGjnisiqejUFHaMS23ybFRV
O7E1ZeemLcuT7cgr9KBQZdjd09P8cI2UkIV5xQg51d+M0nzaLDHT6KOYrOuKNrYU
QIbi1/wEx4lLacxa5gK9MxFJK6RBCvo2PwTIOwl3PdFEqkXuqJ7bfQRXaz/9kV2D
RIa/X63eInvTku2zQJKOArGRHROUr8Zy07JTBmTlJ+conCfJO1Xvtzk8tiFLviNf
sdVBt7Y1m983TEEGP97h2iu5lQW2/g+Op+xDQH32GKWilBVlpCqH5fIFLD+Q2HGC
EcjuQOz/gtI06hk5mYSntfKSq2f42WreqJCqYUlsyJ5n7va+CDMBBpamy3o807HF
h4VzxpzaAQat+Jw7DJwQAmhO/pVw1M9x+TnWfmaOVO3VlzGpc/FVJP75V97edJOE
Hf+GEF54Ao4jaNmomPGJfF3VLCCuT6rne6nRNsdTw5x05pNVY5u/6cGsBJEdgkMO
k642h0qvNtQMbOJqKLbDZrADuUH2WJSxKyalPkcno1aaBLogKVnR6X5fmc3aoOdr
s7cWwsEp1vC+jxO/yunbq5wa9NJDZuNthQ6ZSs4zaH2vCogiWvZ7GTF/agHGISZG
TWOaP31uofxcncq0CjVGwdR6F5m/0hnSKsi7kOeTYjjl9QG8CXhI351dN3y7WB6x
Qki9ZISTxH4i9J2NkDvX9TElr0MpViMULobw7oEBxgsUAdFyM+V3cKtpicp54fuL
itty5r3D5OO7ydWl41RbDM3d48CER/9Gl4RpabbrbU2NNYVIN56lpv+zoqQqkaOd
P2ZhpKNXCHK7nGjIJiwbIqIk7XnQKfQz7o8bz+X0mRlQNw1I8c85J9Dt1bvHQP81
E+TumedNxid85H0d4wM/CaMXqJv40gphpRNhW8S3duu/HdKF4ZuhC3M0STCEJ5dJ
M/LmQn2O8iFyHx2jA4vLTG+79M6e9iPD2cSPhTdTGdSmml+hiaP7l1jy8mr0nhwD
SlRCIJcww8DySLzKWQqV6JXSNYDAFaFAVvkso/mJ74nY+XXzFA6s/vhhAmZk5YCY
mQXQ5uMoKBAcsEENxrr867P1fvXC747Xv1+USzTXxRwLQAL37THDtLLYv4N1hYK5
K1PF+DA2SSYl4+l4RiIk3R4YCDJeMFFZkyjJYNm7ZFJYFv34NVOSKBmNeHIY/Ik/
OjENpJuc3gkpElbvbprH4NT49HZ/xfrFdTrZWpCeQmG9ETdJlnLcrxy+yAqtntun
poGbsl24ZXSFwqdQJ7ACdWByVB9suNmjW2uTbX6NAa6n0rutY2UBJ+KIK4zUOs0+
XBsjaXMIHXgFuS6tPnENLqAeSzYPO+Jgk2a5vFKPOIIYFLzfIzD1kylR/XZiRVRn
+u57ILrLnr3LFoGzJ+y06tmfHANgQvpRiwW4XPu3khVJ5jo8aWm4NRXpaX3vWiHd
hkWpeppYWHQBfknoZ6oC6u0woyrKyEjX9uajGZ3tntoJZ8l4CF1wPLMe/Zr3jqiP
mxpA4xlIAMh32bPPWQVdLu+n9Hk0AU6VnLQnMsxffXbtggA2ZMVzJo6nYB/pMjmR
M10mZcXsJiDoO9u76Xi5CzOXal8tE7y6INDGfa5zKYHXje6t+NyxC7N3E116DgEq
r2NgBkrxAhzwTMSicabrfQ+metEHjSl7EIIClMG7XzeyAyPfX5+KlrZ8YrQrMKku
qQYTuLO8WDcfWuLIgXFRLzBabvVzreCoLA/3PS0I7DLOzQgLzj/2RxwlX0gFBpvl
B7g/oXuSgAdJAAaR3NOvX6u8mIyxlO5R0G8NL0dX83fqSrCvTzyQoqyJANnPwCNO
vOj5uMEOGXU2glioIYY0dZCtDKto9FI9DEK0GJiGhfdhtwWsVYRPWcPjTlNJmX/M
6R/EAJZOnFoAw5bGyXbGWwlurhtsTZ1NAGUdf7l12jol+h7FLjDr9wDZvkgApS4T
+kbNLXzNeJDoXiJLl9TJzKfzPD5aGJe2nlmxDX10YB6dodN5JBjG6i1RdabXc1SS
g01ajjLXTZf4iF+4fAml7ne3YquTb6AandjzWJXTJYyCq6eufEo8SjxCeF5pYQ7x
Dy4Ggbq0uIAc253lx46dPTYH6i0X5mbgSQlnF3eHNtjKN8OFrCa5PjPX/uNTWDdS
kLkp1MmSOyJkMEt+lp0dbFs7VskyYibTQZsR6YljhO1eok2HHFc2H+9n4pLUDB45
+zs28yLVHtHEpb6fnB3kiK2H+pNM1eL1eJy6RCpzzrVu8ihVHTllyXLpkvXMqj4a
faZm3WzzV5ecwkwecjglwZn6bNd8eSHqFuPM6vjRMRjFnm0o3TrYmJqLbzH5Kw4F
yIsUrtcML4Dqk4jDDGpTH6ft1vmlzBkeIdOOXw+lg/AKcU9I4mgy+GxZLuOl3Ucj
3oLIKJZNtESNTVbFUtr5jKhEWymMaYLRS7VBBRItT2j7izNB07RwDn2MW1xXvRRh
tosy37Pzebzvorov9qVCkvjb/NFbKDgAD0sb2UW8DQNWjnltcpGMZnmjFVxBwtqm
t6xSMvLxLta5SVevabrHaOM2Q90HTfr5xS0AIbtbE+lnKslM3/NjMq2GxTYRpj5/
meuBLMdBVt0PVmYmDUjsrINqtm+HHzMbOMNWY9rlcHyTEuKO+536zPgL4jRz4klj
l6vP7c44y789fIu3KREPbd6kB8g9GTrBE0tnLHYBWcQThG1GC7/97rAhPCvUz+dq
JWsDdiIOIXha0BoMNDm98Tr/p1X8n7ATFPEEwH0RFKlZ9I8vJkJgSz8tPHZaNze5
6xBN1un049nkhc4GBqDFcJU1j1krb9931RX3HXTBRdKl5nM07OBhvSXTEeG/Rw92
ZefH7QrPfaIKN8pnLbpsvePSjDJPtFwTbqWaB1OSModSbn0X4mqCUOscFxVuKlmA
Sp9LljGBvtjk4sGP3IggLBn61whDzOWJRZJZfEMqaxHhvBfylApWCY5yG09/u2Ev
bEiTv3IjAXrTKF235FiynHYYUGasIqcLbmR3AkzVvZa+RDNKMt7djoZur0RVmMrU
4oKIY19Ei0seK13eMQHGiHbuZwn3cZo61QJKucXwQh7SIVfAwCSNz6O2H1G2QAbS
Usw/7Hyd5+a0IKabGhIz0kIlTiSkPY4o21J2B4Lnibmoc60fN5Vn9gD8IacR/QX2
I2Hx+MdB5JMBd5V/TkYF4olWttrALxzdtgSGHcs2EUbpqpSa8bj1USBZmCv4XVZQ
JkMRuvffkmeX+w5hln6qIPq/oNx07fbVimB5i17xSLpqXdhHdlca6QCsw2MuKUUo
dcVyQK4lEKTEEFenOG64suY5HDvFvqxWz6DpcEzOiMAGCK5tyJsbNfjqZAJg+ECk
mjNLhRcudauQ3B+uKwiLntDtSoZkPndAuXizKLFNXSonvIFOJjD1IjeCeP3fC1E1
da3EuYwdSKXMX8+lzjUhoDvNOcGmxFxNR+J+GISeW6H1WmXnsih0BRgkxWybQtSp
W/t/Q6ryg2/9JQ8RVvq2g2iFRoWy8ccLW3mX5KI2CvZqRxwo8y8/euKyL+PFq4ki
3bReuWNJIzoT9ab3XGJ3PqgifQqVLoXKyUcvFn6QH0bjysNbaZbQBOlTYNe5H+dZ
R3WHtOk5tYQTVRodfS+0PzgwJLVX8EHmldsVe76LQdCHAF/jgOu98MIPJGyyFbv/
Cf14jpx85SI6H9oi6+PKas7Avzg/VBGRbH28NOdkg1Z/y8KDprGlmHblyYSpxD2U
wZeYT/5pAr/ci98awGR6k8IpuN/hLZsXnZrt6x4rkqqT+qvmEkfVPva/7u8/RjyT
DN5pg2mGg6mMrwPTY25AQGGiPaP+wMrOkoJhn7vFjWv3tdlV3sHBx/hVzl3ZQmai
o4wQBWT6BW5Okw99PIlSx2G8PyOZoibV2QJn6g02XqBAYTj7XPSw1Vn+umZPrKbl
8VW4/Dz4cyBw50raux/RqS5k8tUbSNfe/qxWn+nzdvehhMGYgrKskIb2IqIMPFib
FaAifLy0RO8WhROBmDW8LCUPu4DeS7ILdyXJrOaqc8OY7QdV8Kc0XJe5XKAzYbIw
olcwahF8yNpE/3p34DMaMpcTCYaJUDcmu58o9GyvrqPHirXHdXQgSBOGrx1RKbrJ
Ck92h2X+OuSYBfvgRyYiGgfhhOQZ22BXURZvcZfsDt+hPetZ2ilac0SiHnlNmU/m
ilSio3KxBduK+/orvBnYlJPKLuCIoBvo83w95RlQHr/qdJVvF0Q2ooq5D+bhVqsb
3TQ+A5piKv5s3KQ9qDnmtrZE9SaeCrx9CA4v3pe+jNLQWQbC465AHtfkpiXVJpPt
bAAqICK+EtQ3h+jru9GnU3H063S0k6GwQCv3JX6sbcz15FaZbNdgJFF4G+8fENoJ
uUVgRNnl94sZ/nu8QuWtPiPXrSlO6hkR8nzzcMvgCjANnjoxi0auNMTwIdPQ+HXZ
T+s9RvY6KgnF1QqFecr6SGg6rKsQL6vsFqXvTTWxind0w+9vT8jTxcButuxdCUXW
36Lc0mwhmUMu3QGheuAHpluh5gBoyvFhcTXT2sFVn27NBluhj38hvsnqZW0MZMif
msCYulwLI6OKyZDmfFDiJ9FJECL0eb0FQMvejduacraBvVVKS26r+UPBg4HLX3Ym
qz37YjR1CTSs/kaRpTkt1p6Nt/PA1v5VGkTdG9duj4Cbfpue3uXmqjm8SXLmz9tA
lVMsNogHfD5PvfxSsoxCelkOHTbWB/WpqBE/SilG8tHmUsk2JkqOKC4dWWZIZd5W
Zw75vnIfyrZYVtKzx5Tt88HiBHf33wbUi4m28SEtthW2QRYK9IyHak8viJ3vz6wo
h6sFSR2kO215kEqerwaKXhTYZDS5rV57iYdHSOz+9NrSfy+Nco5//rMCVtNB82Xc
iWo7BPDL4jVAWDzWBPcPB05pZPMcJgINdqHHCtbYmbC+/e/TrvYJ0Ur73Jkd+k9O
is9CHDI7fD1fRtx/SE/IF8Ih5hHwWndBRtruUf+0fO0Y9ci/TqiPjnLNRTIkXtlU
v/66yA4juEYZTlyI8yvK6Q/dIuVdj7KOPuP6Ebk8cgHuQmMt9Yzaj2RDrmqI14E8
IbzsdKFEMA82mEwaQK7V2/8/OovF/uJ+T5K54xVNzRxXbtnh4SAA9elksiE/sdnT
P7Ui75YQ6gm0YQc1n6bDscmQXgJaLe/U2JF+9kKhkbRLGhhdW6zZgWNjXjIUbDCy
q916EsSKTi5f2e0ItOIKy09XxnP/xQ0tgQ/fXOS6USqH7js7qAL3kewHNuZC8dXW
b72LjP4//4PfSNVQgrXDNEMkdnlsQSTwTK2VTDUY635r+9pwLwCjFpgXqi1D26ZT
kPNr1Vxt/2I4wlJDhew0medRTbXpi2APLl7xjoPqkjBC+8wx00zj9Ge9G/yXZyBo
TdcMB+dd4S19GPNk2+1QNuiCiFtoBmIZfIidQPfX3qudMBIXimWnGw7DUwXIx7g2
HnKm5Befb7m9JrpQXRsoXA/Fp3nWVG79K+Rop8oMbX6VPLUYzn+/fMxsVIKHj4u9
nZ3sA/RKmiVFsWzh4hJN39ikL5ooYjoGoRJlw0ezEyBZLlX0U9xzmvxKzKiIx1y4
Q1fRBtnnsECXUE8DgedkSQFm6VIJb20XSXal2COTBNtiP3YfR51Py8io2F6iZnD9
IWCx4f/PKETka7NlXscw8PWw9gp0qp/jB6pmDl7anryqzwbq3Vb+eGW2ZGUZzvof
nz33KWbp4Y8ncD6aiT+QuxLfYcC4kYQXt6016UKit5Q4a9rAce7xd8lrawFF5kzF
ew7cpanujsIZjnc4PgX/EhpS7uKFsN1r8Sy4wSofwzuOWeAxfar97pXn1QdwxK5P
B9RQA9e5rME4DCwOCY3ZkD2tQW6tM02AD7S52BocUASvv7v+MQxWNp1VOzUsRX9F
CZcZv6D8wZKNZO9uDc1vmkrLq27geH5Z8cWmLa8d3PmmJ+4qVZa3UWEiBcthAO5r
sK4bD09rrFVpd2ea/hZHHbeGBQKUo7wK0jX1LWucsh55CFk5Nu+UjCLQL4HjFWcq
7ShD6R1fMjM7lqeyYNJjxGiHwLD6K1QwTrWPhMK2lk1bjR/wcGmhjxu4DaD4s4Gc
aPifaojbZ/hnPijqmNxXIQHsIVHaPPhlKnQwsl7/x/P+panOVV40KBO5UQ2ivgKa
c8pXNkzaw0m4xzvxVxKf/pZYtukAQ4a+R+lwqnSZX37qvUdWf8jlXqCd5dygmRfD
Vr7Lb6+V6OnFyUR2QtltGUddiIOClZRRU7VkKtVYehN/k169TfK6mQxjst10ti2u
iXGddr8NeJgWplkLgYu2aGEUq1GkWVXKP7aDf5XEMs/DhG9tliaXHzCDiahiV769
tEV0baOvOL/KWhkXkT5OggxwhvvGWcKDKCPvpj5q1IdXEap1TaRSCFXTiZRjpxem
Ba+6xpZoYYCT23ZMELjdXQQAprcLrFjqaQ3Bhoi1q/Ro0/D4mUv+PmYQWPNp/sUt
LZEpCBzyzf2T8RajbVX/WR2k3KQdLegoqflSUUtMzNpkUC8n7cCXPOB3JTpcdz55
LlDRfJOY2BBqAc5RwfPPc0cyUAQVtj5dWo3yba5xir9yU0z39dtGpHY+Fqy/8Vjo
TMbdnYAyoFdsN61F57H/phVXfQiqcDvRLFkBI90yS/oW/5mhHIAHsjeQ0PmdNw9D
UG1EdZUlmdcczFFZj8h7xWAdEN/uReyVCn2VN1VRGznpsG8ZVBu3cj+yXLuHPtcH
BVlEnM9QMul42GGlp6VUAp6kIX6IgdTQG2bVYp/0F/wdfdv0ZkN6JxR1G2dScoZ4
fBpRN9VL53fmj4NOjzhwZMdilI/7LRd4cJC2Db5c+NG0Dmv+eG7ufPmADAOsHB3o
R8KVN0NG2fWycohjTO8YzLtHDBu+TuEf+eoDIaGYbA+2QTJQcPRouHb1OG0p0Xiz
a1bkyf4Rk7zxWy8bp8TVORuzcH1K9dzLzzaTYagwdSB5zraExxGkd0MM4V7iZoxo
z3hekh8lbhz8mobz6VHBwrXIxDak/NSRSJ/HOpurZXkSCJqy0utO5hmhiJtSMvgq
h0Wdhw80sBm+wv4RbyEsntjO6qO8HieUMKd4MKfm/YwrujqLHlZ8QLwcidP2zcgf
8+PEIVDp1eN/ZYQuYntIWdKSb4FtAaaxVxAt9iXxYTWq5SP1Rujq8Q9F3Yiweq8l
4xmDfOcJxGV2ElNdhk3LgEUg+JcTHdyrEwQ56VyGXeAAc5sCV7U8YH60gOL1CsiI
0MaJztXtNY4x1b5fNl4+7d9GfSzOFX2wnUVmVb6qkEJbmLfllP005jO9iauv4jVs
QSiR3IgjeO6eoqcfiQbgJS+dR39iJRkfbhALNeCWJCiLwjPnw82eVsdKxD16k387
RbLX1tHem/6DkxQGFnN/pPwXS8PyETGF86I8kr7zUxgCCqbs2K/JJvgJmIKMBtBD
bwOjG/lwyedk9utz63DnzBx4AiDzvnnnrgQuG/BpWsTYIuWUeKab6BYtasNNa0UD
WRELiiLMwyfC7y7YfUjf53OuH78GAT5RtpRRvgIf4CuZXZkGujKnWMGx1xQrcB7/
sskp3/unLLk2ag5QI2Lc134tVgFdAOefEE+YFTVD8N1bYa3c4AsiE6Sb5pXw2MUC
eF+8zT1i3ICFomr3P/3p2GqseYZsYNqPr1n5cdRTMI5XRYwWRDZcjOCPNIYoBwQB
V9b/qIGo+XwZzfpYEeEPKja3OPx7gtd3+wqCMbLZbFimba9aMHQwjeJ4NArTXiUe
aM5jpxl9liTkF8gsinMlidvjB1UOFgj/h26K5SZkId25pDv1GBe+RQo6VWeNbJLC
0WXf3FCTrfW0wXIP6WaJNjq9PlHTqta/q9DXrQEGb+xYP5akaYEIuflOuQR6dUXG
3m/mP2YlQmxxsubLyYjLPYS+ZLAek1vlITli4yoEPSVlZGQu0T8uYxl+qiNmwiWT
uDN2LvclckR9UMmbxcHS1YsdX6IV/ntb7IBl/WVI+tNqkH6qJwc4gRrHniU74Emn
oJYhZ9w7YDH1hN5nall0j6uj7LMHz0arqfZS+r2lVWCQ3hTdw8hmWOY4RqpAf/vS
KdRfvjhQl4dgc7ww3viOI9Sqyx29IGi4shjhsHttpQL/93wvQebvieytvRclaDLw
j8GC/Y7xkOVxTyf+ZxLRjuSaIdxQM0JHr7wePBddZnNXNJDxjMKaBiidCRhyxKN4
mSW8o/afqiQzI7h1HK7m6d8OJvHVp1C6jBuumH4Fl4Xn92FDuC8y9HfMHi4uUHva
zjf8XJFteeJEtKWH3up4fi7q2uRIuzaMAPcaAO1KEePbFe0oKsmsiBLRn01YVO1k
XnVnK+JXvB92WkTWHW4Lgeel/oshrG79hs3sbMbeKCKZdzdeO5ajwfSjFH/hcu3M
vknwQ+XiGWCdIvmXcRp4USrH+xbvJXo+R6bsOD6I6cZn8dhUH/XkQdid4xF76kt+
tSqzy2VECR+1+5Lqww5RA/l/6RgVwTr7fg25jh2xLrSagp2HtwEOpgViKxTDC77n
m1VzbzcKoG8dAVVI0Tjb1528IYH2pkgQUHBw47SceTp8rUCWCf/Pm3pMbdwoSXaV
OgBn3J6V5FItbl1yFBQ8yRYEikGcTpxS9PQIBuGpBevbJSX41j3J0gfr+XeyoEyk
Vj4U8gi1fi3nrq52hm/OQLqpo50g5A3x+kANXKCCCFgPlYIcAZntdRA5fbSVugZl
eqifDN4RoEpLGrezXqJGWswR/kC73vMV9bfLiEg9S/liznEBrWVK0b80cGV4KMPN
qy7tWQD0VgSeIBCMseCspNh8ZBRSiADBZPEYMBSYiSi/GV0i1Zk9JR8zOimmdwLT
zy60DPcfgwTPRrXCPxVYG1KR3loiyEZpjpKDalYOpqOElABKXyHqrVH3zpAl4Fwd
Af+WZrXKBCNr/IVTnTDHYdd2935Z2hPjbjkvoolxFYnga0wq1DKUp6HoAkXBELM0
Fy9hIy4z5GskUEXfJveOAlDN/GrYb8UbuG3yk3i6f1Z+3ninCIOlS350CuCXNxfu
0qzYwvlfHBkqs6R9MNDGGbGgf6xQLxUAZGlAWuTwnyO3tDT+7q5GoiUdUzZ6XfbB
QTuluffUPXpWauv5ga7HFtbiTcx2mKPKqC1u34VvPn+ugMZAO/8w6aGMN5gA7kw9
QP9lwUL71IfD7wgk29kWs4Dxgplnp7i+PsO6lFsdLKfE56YIQ2kPXGqdn+ST2xpD
5lYYHTOeo9+fTi+UeQNyGIJxByBfQHsFjcdJPM3p/rJYgfXdPDee/HZ3mpn/oIPU
hJWWiSiQkZQZUtkFrQ425fZuIdBd51DJBTNBwCXSn6GtNyppGlOoqD14T5m4CO1L
q0p6kNDHY1CseqxWXGAXY+uWzUc8fGFEF87PViQBm/xInhm09hNRfC8SHFNJ+O2I
AT18cIdJ35HT1w5MeggAbmINNfXjMSUMA0+L99xfT54ygpswirdfsKRSd8+tqJ76
32MvQM52xkwH9XjLnMNWBbiVxVOKH5quG7zTQLudV8opsXsS8RIHcK9qgNeQvBKe
yZNZH9q+jFe6OthvSlpx7aWyz5iq6jfpUSyIpXqetN9uiyEZ3PNN47z7Xl+wPFj3
3z7k6TflPG3GOdqKt8+8od9mTHdxdyjTCPd1hVYmr1d83R0Vu9svuqC3DVecrIML
GGJXrZsb5vdjQPj8SdkslXmzfPw0xPu9iX+kZbsr+n7vojf50K2zdL1QcRUnnFbv
gW/P4afaY/m4ZPQHQWOI4WU+ewaK2TQ61vAZ/s0fuMYqUUZezNBsMkORhVlIgEzA
62oDYbkR2mEXolBnt1cyF9tQWH+NtkXt+ravLiB9GXzPky9rJVUyJ0CruH43yMtF
l3qENeDde1LeOnER60MkXFG9IyUT1L4wmIT/n9D1uiULpbfGtirxH6LOL8qPX+tX
AFYbq5SmKojZAfDRj13oJRmyu4uLVbkAK2T/vJ4Say6rkuep82Ddj+OMNd1vRiOM
KZBxo+LkArpDu6YO5ePj4EbSRJU5uOvJVlcTjbEPSUZZ35SQP9YnnXamWEKx8Hqh
NdXcducr4jiVj8Hu9Hm596QBuzH/p1s73mBZMD9tKPha1rgFFQqhPlx3OgCEr2MK
ADxSjenTc48zCvf2Soe1M+TdOwRz389ROadefF4vloFB+WX2G62xzXPr2T6ZV6/3
ouV0PArsLXNrSo1CWmz8tJl7uMswrpL/SyllBhAw+BhcpaFTN1+e+0dLUUYbLZPB
4Dd60pNGsO4izzeIO5ZKR/mg8n0GKbB4I7R1OKsP91Z13zAWHs1Mmmbh7j6I3MIj
FJY93Yb/8cs9tqdlkxCui8t39HRLEBc87/WJfMEyy3LYnWDhLDV1KudnXQs6TNVq
VYhnvoigKdDcVtC7MjEGvWMcCsREEUKUhnHRs6FMVqzvvL24OJpvN8YX6+spEmjE
kf1uAdtxwyFKtsQKOir6dzrtumkyz8FHHjFC98XGglzI8pmPhl+wqtdgLN7kn3E4
HRySH3mbqf5dW1hWFx+jWr8syIFFpHIqtDb3QBJRefon5S8hMgyW/3I3EaeFoSOw
uAxxD4qR3Aqcn29z5hH4YitoIEzvxeCAAQlDaoWcYn/khzVlNx7tqiEs1Mf52fvU
RVUC2MS/1i6qlAcyn6N4MI4DJuM8y+P4/niBKZOwaonnPeia2XPB8fPTUFCC+pCa
HA87iJ5QRPBis7VJXFLZtkXftWVb8UrAjdJ+S6eSPeIMA9PO144MdD20YnDoeeti
1/KLiXkJnvWm1sBbFM2Z7V37Mf7xZ7ly+qwgAQj8pa2xksE/ukds407l4cZHr62M
lug+OAc5VQ5AVKrGqZPJRAOX8j5VLO8s8iD5QY8yRZW0yi5/LwbNgIzgQRa9F/As
R9EX0rW2jzUe4S/bOPhJwLNOIZav0pCVxlSiNr1IeCEyrwFafIG12YfOoIu2gWlw
c1ALT2pUhbnh1qq3Zqz55l4Ca2V8TMOJbXmtgWc+89oP3Rh5s/tYyYp1+LA5CQ17
SkCtUgf6JBUBkKJixXFKJ7bOxGSFvJ8kiabSH6LH9TZ22IAuTnLL1itnJEBN3G4n
t6VDQULWtxGMndFEesY8gjl/9uXOLSJpnsum6VS80O/+B9DTyWzgCZf2sRtCaJyx
Ycka5/ddLGgUdz65C8ZPYHr081RvuhZTQV00RzarSmPadq9X6Toyn0jTCjF/hOJw
5Y1/d7gLuJ5fKNI3KGuXQAsgH/70dMg4cPX7GOYu7OtC1iwCgUmLIa/G5oNjUIBp
6Y6+HVqUC/e/uZqUKc9qGp998ZQn2+CzdCM8J+JQin2Tk/rLnt+hK1p9yXw8lbRr
kxIE8uqZLJ3y4wJyxgSLSRZUhdyUaDaF+AX6RPh+pVU5sE8ynk6OLC6oRg3tJPo4
gh6TH2ZSozU9aynTAA+uf8ebrdyMjLV03r9BKZckeL7Rc13mXIF4ATR9p0XV2b6u
KaKtR1i2IAjcWXhR+qpje4v1j/1MqExShJ/FWorx2Xzx00bFXgjlwXYXbY3LHJgg
KRAZaewRiNHO+xuW6/XStxHmOwhJ0s3PEKMNZl9wUzWWWOw1WT2+Oyj9RNbuo5Pe
8BdmLW6qk/epFRWaQ62wBPP4ncu1DG7Nyq2fUFsFzXOLrSIaeqeRa9+pie4Fgqfe
gpcJrtwhYp5FpsPZxGuNhUn9Unmzq/RsihlSbuThLsm3EmDcFANuLoSyC9dY5nau
w+YPNhOljdEFIBwlj9fuR+oiZcSPkiHFGEHDXW+GWBINzVr1x9TmgrYYqhASYC++
FDOfC/Rhbh4PHRxIxQl5fIQ8b1uBhdG/6c61UAWyVFhVWzRCg+t0VJzhjZIt2mVP
LtaGKB6mA1RrbxMD5sSZWNfKhqFwtKpJncMJWr7Zy9II8w7lyFUCIq/Jh8Xjz1oe
wQdI2ukbiDq9Q1zXbDM/tTAH8FDWpiP9ypKHSYP6dw6feecrUOTY6CCpfE8spqC4
DjoGb/cMBxyPK6QUTu1BKbXZ9aldFRf4s+UpOcUGaoSkO2iNYUO772qm8YJ8VDPh
OiJ16jm8GpiDvro/RBfKVOHRHHS9ZQ2LMg5pPwhAXoo9ndl9vwLeq/27INNgm0qe
Ac411uUg5ri4+PNX2pI81WEmJSvhWdxBzT7/0Te2Nxt5QUWv/ypS+8EcNYQKnHlK
jSB8n7RRVQiNnDWWp6WBHAtSM/nNN4A/jGgkPa8RgrhgQttddn7YPNoFO864Lu5o
QvzBs2iiYnpns3s+7E2aICqd1vZP+QVfa/moZBks+p+nZzk8HA/MA9dQE+FkOlmK
UIgQeyUFQcPksg7+WgP/AC5euN207+0TuJ8nXuHQKBo3eV91dCloMxoogSw4C/Nw
BT8QIQ5d3/gJAf5DUGioeRc+BH6B5JdRkyd3F9YBepQy+ro5aOr4pbDqfD4sooPk
c9gb/vJZtEcy2R6d3jdZk6T5iskb1opk1pVc2vZ9Yiw5UfAC1bcrda/M8sDNPTzb
CqRjsj7O+/2VtxdvUpNzSxe6sSBNO8kqoaIiBxXwvZEkMRO1tymihS/TgdHhPoo1
RTY+fJUp/kBYI0Z3+Xkr0YARl8kMxJU96o6G23SC6bggCvrDWyHWURMkigj7IciQ
PhBXt0Q203011J/1IHivw7MNpr4p4JLp4k/OUsH9PVUBouCUfy0dH5RXGBtc6wbG
OW1AJ7OMQoQP8H3o5wF88UmFyCq//apt8m6cf5T2vbqHilvWL7C2rKEBcS+8/IVG
PY0aw+17tu/Bj2X8nZRLyg==
`pragma protect end_protected
