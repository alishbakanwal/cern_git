// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:09 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SyGsZdlv8IdSVQPcbzkhXz78uMS8MQeWWofYJAvooiYaKwgOTFX327D95V8PbcnN
LL1dUw9vHOCLS0bcKTtbyHFg5kr1oxltXuL58MhDEo6M37LJV14Tr5+qcG9FWRWX
PMVyE0sCjLsAo+oZktnLyF9lgWe0XQQwIdQTAFXSWgk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30848)
S4lw/4YRqD7OLeAomVA+CmfwY6TBRhUv0EI1RuVNKDvB/ftJFmUGZ3kYLnlA8KC3
R76HowE4nsOQvUjnUpumTZQo2OlgTXn8tfCBbwGmpxKlTGbhdhM1We8kRgWpvn4T
5LSVZ02RlwCPtSpJq3uP/Ah97N8eFgBURhRxi/95MN2zpxrpMQEvSUQcayDxIwTe
LVpWxlJfjsAJIu4Lju3XWVXe8h2bivP94hVukJRM16675cuEOnNTsFpMVqcUqK1q
WnmDnmgWffSnjM9LxcfYyRyDc5QhsaMYzMLl1Fot4y6ZwO6lwaXBR5w1d+Y7bgc5
tl7feB37GDTW+mhJBktAHHH3oXw5QlgsgG0SekVRCuymcocgdeomHj/vQcKc80jp
vODQ6nLcj9ztR2ueUcZTsdAMQZqb5skhoPzfpnph/kfcNrcoD/KP3TI76t4HLE63
dqdw+jbpnIks5pHn17t8J2LojrIba4IJBweIP6qpvCKFw3hyFFMhLX9c0PdjtZTP
hxGD+XyxkNQJc53kBhWS0JuFAFq20JfYE2CX3gNT1G7dmQfW51bSlUKUhCjneFLn
Lnnes723IMUFMEUNVClL1+hrEWvWTtA0ekKPYIUY1OPrFb2MM45vwctRuEMEzdmT
Lg4ZplGMz/O8mlRls7Hvz1M9R/u8hT5dx6+QQEwZqrLDInO7r3v8VVvC8UIJjquM
CClZJa5ZUV2iZPdRP/iyxZ9TaTeIijd1AbplSmZZQxR4MdzCSlQh4s20QsmMhQfh
AnA2mY3QXV4jYeI2jHy65Lzde5ZzXs3uT3T6uQUMarRZ4/sIauP5v7doHIcMU+Uu
Xi/2sompYtjFu4Ez0IOLa2/VrtRD0wRcV07l2o1Zi84QsBOFTCdQ/xD2+XpLplO0
Os6hhObTYxjT0KuMdnI2H//sGh7UnbC7cq+58gwYdy5BiCxivan3CPm6qn1iTsNz
4z53lNdNkz8rG7zXnr+EPhdllKJ1yHn6kMsEYD/jsN8yoZHClL5nBcyMuFNJF9wI
0tQFWhtMplMEf2LVWpu8vxIAcRTwXczo3VXiQQFJokpawQbFnFCpm2SF0JB5MWrQ
WX67EICHlmtSnztjB4rOnydNPMTPsjbBLeG94in73EeKcRAdzd9zbF1BdIGMoNii
KtT9cHzlQHeosw1aql6rmYg5PdlrFLJI+3MqsAI0iojpaRGD87YpqbaaM+9STqsy
LcCv7Andbxj4A6tCDGiv1zcDCe5fGTrwOR2PmYjTjYidzNPpMQNA2vh1cd+UMyOR
EuMvLINUohbcXe7rVoUHGT1ZAs8km1OxfKkbALWRqRTeLhGiQ7mRKpi4ua3yysms
QlHMexFMw+kNrEERXyiX4pPwaoQog5CPFWUPdFRhrutet/aHKMAdQbqT8o7FIn6x
y1hFxsRJRHxEI/rYjmKZlHxdbp/aPnvE2CD9chDZO6nX/mZ8YSkkyJg0QApVHCiS
ZUUpadd7rHxc74Ol0PCM1Ts8u7qaMfSRga0zb96n83tO5XhQVlqTxDQ+l+dzyzOX
7k7cQIpA4+EyOyhYMLw2H4i1kQU1y1AKkBs0IhDcDCPaFHeAUsRaBgyWluHs8E3M
Jy62/8/5xK5MQ021/rplbtC1G/V7KAHNCn66RmelBKYYt/z6QH86i4cqkX+aUKeJ
Gf0ATz7MZKW2cqbpvJAJe0F/q20a0NW29ltWN1gCSWH4VFAKPzOyYaBpxYdCyBzr
68JUMGSbj4quIiRQbH9MoedEdTeXsECk4EUIt84A/gqx0p3QBwUwOeOI0PYSVzxs
3cCu+SmJHxw99Q6E/nm5Q1rfodsFaUW9JqDMFBRbW8+FZ5XwpF4peSwf2UheeFrD
oq4A8G/h7cbUKAVnIDyhA5YB8aFzq0sp7N6Hg8WpwfPDMs7xMSd6VL/R8gyq+d51
0KYQ4PAXPMX4D2GsPmhgHyKdHbxY0xETzf3pmb/dGny0BM48UwNWesWx1HkaRP9V
HK7psSVuIew3is0qjnpLVGMidzSsZXAdZCsLhK1tACnnCdjpaqost4OR0Jybcu7P
V0oxhApOtpH2a5fDf9mcoHGrTEoKoV4zagqLrGGUzq080ALCBvNRiKBY2jcWDyF0
tW1xFrmYk1CNaDRoWEDCC2igHXuwi8xvtNAUSGjLT0FjB1yUWn1QWqnhG/tRMPbV
FFaWjB3kXGeP0KGEYY2GCGeFiIR5U4fmC3LRqbLPhoqdUgHRKCieS6LrQqUfGU8+
IIPemN3NgnNEXtTZHjCkV9wft3oFIpJjM2IGvQsgWaqAQL1Vy2QsntU48rbQ7vES
Vr9zNmJ6jISvZKPiiqkl5XCkCDAIRHRToieuFJpfQRFCGWFKGq7hBYfhYjsa+8BG
KZFIQrdtb+D7MhxMKlYth6aKs8BDc2OiI8sbqDkIRXRh24IMwoOh7SdMYX1VyrJo
74tAL9mvBjWJ5RDxntgJ/H7zOYxARAOfGDYQXMWh9MyMt5BWPlsgHMeMvNtg5gtc
ys0SgvkFMUMEKCxQFDjforf2ujjCExFqocmqVW+9owb7fb6Ebn7YLF9cbSOfeCLQ
f/UJmS95fEpy/BRgaUgtfqv9X9eIX/b37zKiaDKWAW1UpfjdTMqafBSu34B7dPWc
KDbTnTc/arm6e9GHMi+RA0fgqDCJmcKNDD9fYkm3uuA+oNmSzR/U3oZU+dIguZit
CiWzYlrV60KdX0QOquMn1V8u6PUdUpAkYSZfnRLOzo8orpaRuwLYCrdsPhZDSy08
V4pzq1LASKmuJ4YeJhxL6dWTI7sNTzyLS33g63cL0naLqTS0Fu7KIueGR8jFrDxl
CtH5Ta/UZtRjd5gP//52YJGskAJibLrXfzsd8nIP1Y8nV9vOdUfLkcaTy+eOLOLY
MF9mMunftmDBw3HVSXDrcc4a+jvUvia4DiC8I5LrGuUvgWfe8GW4qexgv33hyoA5
2WWiBDASoL/603Ns5NkYHspm1l+uyhM6DxpE3mGaEzznPTOBgB+r4W0fDT7JOHKu
7SYr7O0OH9fB3RNNEoQpFlZy3XDTEn+6cagOStBw5/qAWL9am1aMvzmc7Pmzv+na
rkqDw9tzX8oSyLTstGkOdjIsMN/fkH1UNLN4RzpYJ1iG903kq90+SWKsmJkWYQiT
VpFN4CGSjUNwA3qcZacLyYYtxIaBd88/HSaf6N8MHH06f62evBBOIYt5pBmf/tuI
Cs8+t4N7nb5JWdfWJ4KkN7Yzm3A078FeVCfICjUPCPedYUf36mmigjcCF7sadcNU
3IdxuF1MVol8v8vDj2/0t+en38X/qVDjS644TQDylFel/IcZImLDXKo26heraFxT
L3X/cRat4nkZnGrNjGKj+CslwLqRA/3Q3V7jqZl+klo+6DwelWtPiQgc/opUi+V/
5G+lqbNSMTEC3ryP0+pfPQsG4lkWw2Fxv0Y9WdyZ50lisGeirSsyMnZp4NFTAXph
6N1d4VcU9B5h9sVTAy2eyKNz22+DjqOWkAqD9izNzS43XObwebbBzg/q3p2JuMX3
I6tWrTp3nSiD9uBsctr/ZZoA1xqhn6zVt1u8OHBTKjkxSmj6PKivjEntJZIZKxZ2
P/E2j44ADDuwCPQT8ukDETc2t+kx17gc6kwDgsWPO+wy4+HkhE5nmhM2tKzAQoLP
o81DnITLr+zDxS4zw1Jcgu1nCS5pBolxbG6lWv+5gkOoMaRV1Eas5MiOMqrUik1I
o2rjUY5D9pGh8D/r1ax9svpHPdliNbYV+8sZl2xCSFBJSNjR1eh3h7O0XBJgqZgR
EVjJqnxd20oHn/M9GH4afJYDi7ZK3hujzXRYYfO1oDmW3Yq+p5LL75usH/ehYLF1
qUa3lUDWMyfzuw5kqOfdtrkdMQtl8Zy7NtDm66NUJkEybYx43K9AZaVRyIYS9KlH
Vvv2c+u89pNreqRZ5eAzUESkpx4f3DfGlspP8SV/3VAYOOKhYsu09tO/rkqwK350
QqLUS6yWuTB0QGUa91nkniys9ualBG1PgUkPhJ9ZjA5VFRoOGRoKRDdKYA830KAf
bVF4+Ux0FPjEIYchFdOPFC7mA2zRgq4ERUIW4WapRoTPb7YOsUOV6h5dGlsmyu73
WSiJC14DaDJ2GZODc1IQOtsMggKNqki18+cGd5pRDI2ewd8vB9pvSIYR1EIqJs9a
38DcYQUV6v3nuQFaMu9OmpYCobruU6Fu+pVUCwa3iU5Alz9h18I1zxbwh5oC5W7T
RYoTzeRshhI7j1L6v2Zz5uxHl5OTsRfYd0LQbbqTfIRj7GPEyWScUHFd0srLZEIy
8chQT/oYMRcOFSuGBotS5w9/XIPtWKvpRBkNDgWEu30AmuFVLvCI1/tS2L6Uqwyj
n4Pk6LthJllEC59lcuo9xhj29RndlDnwRfxlSadMVyGJ+W0qSAB4V0jdRKenW7ru
UYrClT5zwS1aT7VYF+EBdiawodPloBTKfd3vZERNGnRHDeBMasG4BpWuehqAHBaU
uNUbCh5Fpg3YyNmEfCPB2F+1rrP8Y8q5hyrpbdf77qnuhecYbetMAPGHgIrLZypk
mPlXJtj8SwrOK/A4yE+CqUcM2Nb8z4HDmHwrfQq+lTvWV3J1ZovzjdfCYeUMrgOq
k4KpX+nXHL2Ke1BbifnSELI6gs73TzgtRFw5J3OD0g3Ycl8Z7TjHu54PRx1YOgpj
UnakVk60IxzKDOaxWUBg46xpfKA4L7DIxeHYy1bWRokFzt0y34j+Owdu1qYrHGIm
z8i/HUnqhkzB88JF4njd8++yd2tKuwj3t037whHdazh7tMbXjqVKzfE0CIt3/+Gd
2RI2kDbLJ3j+TktmmQ5TUShdPXsgLKrdG2An/DBOhplb5FdrSRYxeQLG2O6K8qi4
rn53fSR3JbmcgJa3gXHjXzntXA8WghRLTJ82O1OvspLpdw61gUmUG6ho/HCwAA9e
X/jCkLIu9ARTdi3wLwup4kYwKpc00UPBDrNG2rAwTlJO+OGnb1SvJsZP43gNegRa
m/eiuzRvRSD/79juu0G2Qvo+DG2+fgNcjIrER3EXs47Qcz8RsV7hSxEMeymd73Tv
tNujlzmo6dB74BeBhilKYmjTpyR9k4M4p51wKQPDDBUrWAT2/+j/7ihULLsT1T9F
oskCG067icuBVh5T5cMv07qWNqT7wsuHRq837hEmm5cLTpYeDvW9FRMyca/BjmW4
7nxWXlwF0aq8M5UOkKbzdwj3sH0OkXpKgQSy9MHEr7P3gcJCJfVDv9La/7kS3Z3z
P6aZnYogJrpVbWq5JZVQgqdhxUHw7sOMYjW0FeF+Gc8yeXYNzSp3rITCxkOy8s3S
9rzTEEfw2S6vA0JzUAhm9bX/80KUpihfpkAQwzThN8pzMgqfb+swnUXH8zIO9L9L
wDG5MKsVx7YCbRa5jVF6FFiNJJ8GaIhlvVYy+dtz+Xze3FqWOqs6Thv2b9LmC+oS
/W6mFX+x58foc1ln+7ynOVuUaH8NZJaKssfJqlhGlAeV3krbMlVAZ+7WVaA6lG5I
eXSU/H/zjS1YSISv7GNPi4G4tlbwAyXnpXYTXliXJn+XScOqYuNjunpOxeLLnDmp
CkTAGgHYzK+EKWsAIUqnBIKoyxNjV/9dJy/nw9zrMKDgjno2e9OJ/ckKDKvGNqEr
h59D2jlpnR836bi39mwSNJ3UXOjrajfC5XQ8v2nVQVHzjDeXsOb5od3w7md6/Z36
EeY/v92QnV5/KFLEgLntC3krx8TTOiCH6ZCDvCNLAt+TdQNwEA2x4ukTBdXmty20
zOds22rs1QBSnfjAa5CwOs5SJvVsejWkVBLOMfncVFVKCZzaqZ2MEUd4yCe6dRtA
rR4mMK4IQL437/rgpAlVlLefLQw4akduzBlQlZEvEkddRG07Wrt+5VsbILElxq28
LJu5/0eSUx8m6iSiTg/ETdoYKM4iKgUuCdU8aXD1LVWloY51uWC06mk4iKZuxYxb
aBrFZurQxpKBhRXeumvMRsECSGBNhXBDAikGKIXftAZF/DwngiXljo8SqCf+Kq2N
U8U44a+v1bowIqi4WbR5ZiAvN4Frn/+he268+SuEpcE/OSyqhIt8qgFmOW1uhJuG
bLVfy11gGbCF/hTKaLVakcirr8GVAVnr5Q6cgb+D+2X1jwhf7bf2+k87OZdzcYEl
9OHkAXv/3qVyS3XS/ceVrqXyxYlEncl0Jq6GWkrlcYd2aBwhquQvyV4rgjWMZg7C
8qoP8JtsFF5RcmY0KtmsslV62wWypRflkXRHwKgGw+87nwDyX4H0aUrheK0QXe8g
uxppBAPJfdDkj0AyEwbYhzDUSSeYzwE5+ib9hBOmZloAJ8R9K2o7KhP4Lf3FWeyZ
MKundj4BSFwHL39w7P6DfzXQTcbbaG4dzMY+in78mLSiFA5v453EivCCqq6Ikpq5
wZsVEQ3430GsIhTo5DSzeMISAIjA+1FElGagqsxYJAtQlBi19Ma3fgt18REFE+Xy
z9Qkzy/SN9w7TJouUKHf17DUQ9N6btzDzmSHxQxrQw3Ie5HpD+VZpmCDYEdQeGaN
KC0O9aL7S6nLbz1GdrXbPI802x8oEhGDhWmtjiEpV2Us5Qqg4jtaReB72uZSJ0pJ
MqyaYpxbZU9f0rcYw2DnDlPIk9/AWaVOPtnxiCZDB8TnuM1fmzpOSY/kmdN4LaVo
l9cQH7v4DPmJFxNatvmCMva3O9S7uSQfIXn9aQhmOTAOsugFd880RpWbrqKC3yKU
AFjjw/a4KfYxxRADD+ptrP7wL4z78AwZhSH3geQ+i5UVH8h1kDQJ2II+UiDObzLt
+IIR3dqQHhFZe3YZBHtym5ry0YQ6IFjYT3zEZibePrOWC6upoE/JfRzCOAsxO/ek
Cq5Fi/bLkbI9i6l0jA/ukrnUDbcxj85ju76PvEZKkgY2yTCXMZPxuWTsPkjMQoKS
sBpBVXc392rsmvbwAb0hkZuqVF0e0O/cDZKC8YTkJ3n3V6WAijTrEbk60B4SQl0y
Sm5A8j9Uab2wCtmYV9Rqn0zow6KqPuW5q+i7Oq/x73eK9xJolWYof6AsA9ppeXYL
BEG8+wB5hAdASoA45fWVMQZMiahxYGjloBMudaFDIpWZReMRJviUgJM/YnAX7Rbm
r7Pai9ahsa/p2m3CDLc8mjOqeMXnhgHabF4DJEcPqT4xShMLBwbBV1JnGVSMZeo0
45bvK8asdEKSBDNENUJtE/wrZN+zUS5gtCm5NxLLZfyNFw3HZErG5EiqaMSMqOAD
RfpJGHf6T/kJP4oZO58DiHGeeoyxvy7FS0ijBlbsaVZa2wv5PVwarfwN2kccYUMf
9mfh+F+4seV0gNwmxFZbu3HtKJyoUs8S0FeBIi/OaIs6GDpXwHTUTufHRpvzEBFB
jXH8iMQ+Ce91zmeuLeysFjuuZOI9z2lsjPGDQiXGFNgapEy7PTjp07F/BFoQ3tf+
mkJE6TgZJpzElQhns0krGs9SxoeOkVUU5N3g0w8aBcaycgO+vGUTb7jVo+ldeCnv
dabeuZ/4QqLYjjPxVtVf5EvjrdB51sOo/BYpze/1MyzacL2raP2+jNkbN6Wf90EE
VbMiQLwF3rLnRpqgxp3UpNdd1C/OKAe5l1ARlglFJwjpdrpKclF88lTPANRaqYlK
6aCyB7V0TwBt/v3BkZiZC95TyjRzBqmsxcvA0aqztQwI4XnQyL0Hn53XGgC8rZNC
Xwn5G/4ZLnIzlF299Un0VaHz/7nOZqKM4n3lY+B3g5dne1FWplHy0E+DUxiA2hHs
P1RZlVrUSBykyhcKC9xcuniO0HmGFvhltCT5rWC/5JEiEVrxmwK/AODCPXXvnkJC
KrgwtZvhuct0gC6UxuV/qZmRfJvsmXEGmgOdc2CAM2LhsQ4IOai2vxXGhOAFaTOb
ub58UXvOUj1fhVnbBnK2M/+G7cSydGCLkeL8xgDrHE8d2rlMvlu6bxqHdVvbOstZ
OHzA/j15t/OYJ1dqPl8YVhN2ZIDTKz457jhh6r1Utj4E2Rl4bdiS437KK4rN7X0N
18SjoiviERHTRciuWcfr4d2Wj1lpwv9N7Quu3Jqbvyj6bRUMD6qDzXinGdLVjA7I
umnFpJNSLU+DtgYjWNjAP1LZ+7jQk0hktXAsCT4xaQnItet/hFbAa2kyjFAX4Qnf
pqqva3jiLZd8dCSGI0LEKu6XWQGiURR3ITCCp1/HbG+MVEXG/Pp/N3VEOpv1w9FB
Pr8icmCINuVWSjKdG4z9N7YcJhmyWA9xw5vSPULBy67wUTokM7oOxtrZTexmlL5f
BeIuVBdf3u8hVWxWWCx2A2tM2B+yeX5P69eq3v9kjHGjDWNWqdteeDbl30eFbX61
5OBqBpBAfypoy1Yvkvauan8835/giAavyqfXISBlzGweZ/EOMuH+5cVvvwk1boK6
JgaDausCZOkRao+OnGTC91s5vz+dSYVoZykNT+APKvsN//GuG97wsbudwXldGbe9
2KOe6uIdog7TDFXDyVMZbSDhnz8CNCxFm06duDKfE1/vFrrn+8mFmzZ0RNazZGvP
Y1CGSln05N6p82vgVPrkqMXNoOnccY3xWIIwcp4/C1Evz2ZpLyVrAByiWhQgZ1c3
Zk5HFucYyze+gXsxZ3TdnDu+ltro+FB2Vwbc/7oRsUh6tEl+Ln/PuVnUFOxweimW
FNBwufeGUdzwZ987Sk85Zgzup9O0OPivaDaK9OOkkOSRD3pfMm/ngkTbTuK504wF
CO5RY2LslWEUljLyxbUnDcfm7Q0UVUFSONGyYv1BzPbV6prX0ZSFFPgiXviw0WJc
VUZjz0T/tg+wB5Dw/H3GlD8sP/MG8X+ugXCkaxvuD/oDDSPmH/xJqEp7NkGNW6Sc
vufU0ax+oGiVF6CFxmRwj4sdpMiEp6/8SZUe0CSq99TNSlwBbODlXCkhz8j2pxJ0
bO7LMRucwcsYQT9Mbbo+0MxPDNbvAoHREtrBIE7YU2prCv2OAiyf4d5ZO4brTPKX
CFzp+7sCs2wsT323pL62MhfkTEYQggA1m2PXaDC4Hzi4Fy9SXR6X0t/P0kUDNvWW
43HcYB76mto1fNK6goM9eKztcQkPtVosRBg7yvVq2MLyxNg5XGtOFAXP9JHfN97J
2alRPIfrWSa6MNTQHn4FEbhBZ9KZ6dDazZlPNPF0CXWVkRix/cfeKChTxxVWHquG
w6EzH+nCztr/71a9+RJEwbSHVuxwRHPznhpHKPf06le8ghfS0Ac0SulhU0A1XXD8
v5RiUEMIo9+jdgXQn/Xx7V40soEFmy+TSLQiw+0qaZqHS03hGQiufTQVloncavee
aOnfRsPR/LeUmZeX4kNYZbAd45vRGOqY5l+fA1UkLdxuLnyPZEgF9qrZd3EFVGvS
Zt+//+CKG5fVKdP/GJBk/sneUUuNBOQ2s4ualCR89rPXIOGn5BWpljdBmuvh4oel
m4WAHOvs+W3YPR/u8y/LL7PbmbnKCT/zvcRtwCs+CXxc1AVLafUohuydX75k4T+I
xIIodgT/oMAnkMCbyQ3wxYMhkZYQBheqBBHGsjGGSHFi4g6K9JmSdi98Q2EgkKFg
bhvUPPo4dmcVXwvBDS+9ONRKYbOHOANDIPJjGR6AktO4aZyasizRQ5UGIJkwRQ9u
ZzNGSLyA0En+KIdRKtl29eBtOIkgje6qe4Nm/ulqbFPowE87VI3anCXKSZD7pioH
0lp8X7r80Bd6b6HA+JMULsosnFOXSDydypG858UjTSrLjezXAfwzfjMkEdRklgCg
scw3ONRKWLnPCN3nlh7y1GHpb0VugwwSq/PSN9+sxEbaSy2nT0hqLmpDg9DPah5u
sT3VvmOZ0s8q5ZxjeOAalDwYQreDZ/7bsyy+7fQFKyZWQEaXZbhG0bLGIl5o2yn5
DF+ozbhJuc5xLY9exGRFmznyH9fRrk/eiSYJMzawD94Rb4uTrEIMTG+gNRI0ltiD
LpAsJBZyPjMKeeGPblyjEy0jBLCYkPUGIUEwSJAzSYzXdZJVMA22QH78pyhE97NA
1VN8M8ZoSm17x9Nd+Q6gQvWxjZ3j+RnAYVztiA6D9As3W3JxcViUnxFJhRVoDT//
EJRkQqu0RGrD4BbDk6e10E1vCVz9RYovItFHDxyv8hiW553pINp2FExJjhg2KEYj
EBObX9cCbesbHWuRILey/ad+bb5B8wyYdUNpG/kJ9en+ydarI4R88NonGY5gCbSj
WnxGJLK+TIX7bPif7B2iVIqV+STVkmTEvJP6N77KTLux0wtUAQ8sJ4KQNBKVwBbS
z/4gi48iAfb64uEUyDuNNDn/m+zrmViZlLKzoSWpksuaWCHHBbBoTWSM7DiBBOKb
DW7Ic+BqKqY25K4kdUa+jrZFu67ez+jeDVhgdeadHLCwiypUA0anbvaeKoR5EdeD
WWQhyAQtG5Mav1RAW5/8ciD5eM5Dtn8HtOrbKVWeKb/SRWb1LaEOCW93FXnIEc6c
eKCx6FnccNxwTGhWBU1vvpwKq9c8hDLBiFUXFKfGH3/TX9bhBSjJ/Fn6kvAkJKp0
jE27JM+fDnnQgqGF0+3bD0bbtzhTKtN1SRWS/5UoSaN1zNYdJoK360zX3Y/h1n+R
ZiDMzx6Ow/79CbJxTzeS8rXMaTzcjJQ+xWABbRLIOpbleRUDgrUf8vHV1BaBgqJ0
TUOLp317jjSVxI6cSfxg6CyuQ1gAR3BAwQ++QtUH9gzxqTJNIeBOcg3U9+4ZM5Fr
mGIV/EanN3xU7jC3X8lgKqpNkLvf5fQ+SDOraa1rNQP7EjPfIz+g3ALAyL7Pb/i+
mM256ajwPoRAPECe6GbHRR+pwGmhAiakxxHMs85MPeM9MwG9UMlgwnvQ70th6uvX
/bqf4kPydAW536LiHbZ7LKf6xQqrNG3Nq8E9+euAxjprbGU9iFFlYxII/Np84mzl
F192GcoM3JJmavihLqsuVHpWG5Lxk6tLfzGOxJ8r7TblDzrZrbJPI4lnbjcW6PNB
8rnH/fyxXJmp5L3pEEP434tw2oDFLBvZO7R9X+Ox5jg9REYgJi0lUb0bb0/grq/o
zxlajyGDuBJBEaxqZyPqUUxsR5G8UV2SIvXzeldhU9gtpjho1Ds1b0nrS4XynOw0
Dy2KeeV4jhIcKExNHzQy5AvrLUr5Gb8JXJDnaQ3m3FHkWslna58u6DnceFUCYGQW
U+BlVRJ8cXa4m5f166FgLEi0eHj+jR2fzFFFz2qE/GKerFbsDaxnUDHEdQet9KlQ
Gmc35mBLw/zVCGk3MnIC9pNKx2xg4JfO+KjA+kxqsDEhqnJbzvy6CZZBW/qTWlEw
aimBR7eavwtdtLYBH2V4oIRlj6urw6gWTbk4KPks0RcvUp0UxfWYDOMC+YpmB1Ie
RNjTlqkRAHSiMAFX33Kedjr1ddGZHIiapBQCNSex8tbp4Zeur5DQdfm5zMc/mdPO
tfXeEM1ow0o4utawdnpQEEfi9qsdej/dHhwfbm9LFR+ZADK21FBQ2mGqJoxhKmJP
23T+seWQHTXnPbwxScB809KDpL5wf+lvgziIw0EszRgA/UD5H7A6f3k1YrgC0wFR
04uBl80AVJOF+VnEzQNvemAH9kg00xoOfJKiyYmpCnkj4t5CCgjaXltaaqZzBsel
67W9xtwga+gWeLAPCcT+VMnT0skeLC99J4OO6AQnFnkFwl7VzE57YOK/5lpXn+Cn
ahqmWeOc6SSS+XwqZRer2Sck2LIJJ1Unf52iGFneWer6x3lX3D1EF48q6+sJqTAL
psKJpS6vhTsF7HBuouwT2GmcD/cV2oztbP3vYo/yEvzswpSEIxpWxpN6SKEoHdwA
aERrUHYZcUB+DhMldbz/q3SwJPP8yMhKcfj6YWO0/POwXlP5iFT8DSJORJ6QRZqJ
ddIA+WnmcNo3/OFA7bwTYAUrAZzoXEv5ywao3djN85Ini2sfj6v4wjsMt+2rIBv8
WWK7Rb2qVTo/rfvXon+kEJ1Kxoo9reGGsS+/7ldRMZ3apBfgk1CG5lznp3L7FcAI
ieTid4Y39X74GM9Rxa0mZnCEiJv38XNxdl47LCBrK5C/7sUuxPPBJsnsDFHWErEw
GlQXdYUTXNRZmpo6P7joC006x3vfeJRai5N7tgbNSpp620sWcPo5+WlpWG23Rsji
NCE6NOX6f6NqiLSasg/CZnRlIS1QYq2GjCVnPI0IrLrQo3O8Pt1BNARYQ0IiNYjN
b2GnGLdN0ZZFz8mo30ICyYDp71347Y723INnm2t3eFMn4Hf4Hh69UPGYERU0uJ9u
HuOILPAhiS90YYnNmFkQDdywx1m3CqB7WTPCAyYGsITIo65xkDNUBZHUm3uvTHg+
e3lOo+xltViuU8/U7rnNfKtq1fy8ee5L+7Ab1gstrsXwJ95WF7wC0TLj+bsEFhFo
ldgCA9w9UYquWwDT/8R3MJmhQQSkGJE688hqntmvBzVK0ydkFb3WrBGDBsCPakVG
ytw7TlWKLD5QO9BxnHAwyzwgJaKtS1+YHHi53WeHlLlTkBezP+hOQzApuqeIJFFK
sbquA5cceMXMAy13iK0O5lIWQASyrUnAihJfHaIsnoYu0jkAs6S7Me5cYjultAXP
snOrav3sc2iSThPiUQV1KalUPhS67PGaqIWhMnjwNtTCT0UKB8znhPXOb6PsxuyO
dFnpfuhNSNHIVsgOjLxEUXVSZHVwFHTzSkgc61Acc8l/AJg1gBk4nkKqTwna8vvr
rr9enKMN9+DvK6dUbH3ycwDT+vu5UX+2czkk4w9vaiHQ4E/bsDP7i5OwAqvhJeDY
fhDOC5PRxTz7as12w+Hvlea/rxGVw6DvXpFBcSMO6iEBq5mVbLKDe/E2hgDS58t/
WeV4DaXZCbiAMvf+ieak97RtzmZgOSfbLRs8NQnWoJf/FCCXNLGbrsFCwT9uWs6B
yBchV5ZofQ313rQTCMfbBmfVi2MRx9BaPl+DmwA54FGiUk5KojYImbJJHN8VZS3p
7IvBWwQSCJnIgEl4bDRu/jwSoGnbvu5lxQ/iaoEirqVuMWg/Fp3QEOw1VKeF7AQh
jhzNoxvXGYFqGNi46IqWwuueI6VQ1u/NxJPhcMFEF0QRssYN476MQN2M1IzPEmor
zUAfrVia28UjUjX25MUlM1hk+CY3JgRQII7TKP8KbN0N+y76GbHj9mZ27X8Cwh+D
Ed6CAL6lKcvqy+5EjSeJBDTnSCCf9/TERh2m4dljxgsubcezb0Mp8mBOCLIrCq7b
Kfk1XIXKSqqPnCDsdBPsWlQDDOFjDuLYIBuacoo0BoMNfgq50Em8U3eJ2sT4orzN
y0KVKmva5f11+INKyq9W5GuMexII2J8yTDgeI0e0+rfRSH09MBj4oEURtytJNZUL
MTBmmacmEeNFY8714Zh61try2LS3XQf4Nv+b+iPNMOfDsHshSEOrhMosmEi3ur5K
jJA7iJccNgDUoE4ZQN6OgNjTH4/kaBEvXzYJGIW1USHSEgUPJbqAU3afi5YOxTLH
h2pp8y8tkpX4kmzgnCcBRNjC4SELw1+QeFgwZv0CxUUW9rcb4Zt0JdPHtjRFXyYP
DvIz3dpKbEyvluvbZVh4JOCDIWTzn+OLznidQStFlQ1278hpCaN4tc1bz9umVXqG
SkS07yMLEfcllMuiOw2pXefFg3DM5xOspklwKr99okeABTVnOmDMxH7pZOiu72vg
bmAcbJ3hkjyZ3cozrbKTwZGoevfeYHMk2+2DkAVXC0gq8PQzytg2cnFtnSKcNM4g
5DSO+Vva15Uefyr+qooEpXkMSp/XSSADYq85klJnNsh23EHqeSizfr0SGvWptCtK
20fqkjD1jHMwj9QcJSQ3M8rEH/So6w3xIFn7bZuQHcw192HjzpIqNtZoZj04JxuU
I5L5p7HJH1Ammi8KFuavaiJdN/KmFNE/GIcOuHqdp3aAeMS3ylAL2mF40VFX7fWM
lYaHAzSf57LWrkYaBm598XECeFX6LNv0AyulPotvw75pk7RoGeyCrVKSiwCvz0bS
sdVsN/pX727n2NafCh0YusDJM6usOzgf1misT21XF4hIYUPLFFW/ilgQksj4LvDV
1CukQbeoKLxm2+uaNj/z4J7rAzmRu7XtOaPNiypMWroGGVTKhyy/ooHHurkb0bak
S+1lNzF6diJFQI6lNraGEAUJDLACW284ZxBeAQd9P44jBIU7uXaEhl6zbbazMMsK
pB+zfvHCXh1eHHzm8UjL5HKmndvk8iK+IMG8GuvjDnsKae0mlFhWLwWyAM7ye+vN
NRUChMYbCS1fs0jgo+F2cj7VBDrMa6ayNNR+CIB5T+QLEmjQ0G/ecq8mbf/5LWdO
0qeABvKp5XJ49ySaayqE1DR+M4nyLejXRNSEFI5tkDtaPsHHb2mExTIidwvMtiNM
90GCBFAV7DbsNdhH5ZKqFgthQ9YVhwc47McjZ/ywQlfgEJPa+bHuAftNfxwq9p/l
Qz9Oa2fhRnS+hOhVLjfw928JG6zLUlEsiACTUrIhn40iccs1cpr8j+QmfR55jzO2
ekE9+ZYDrUoLVBvVPV0T5e6X5C8SQJ5N9UDoPWRue7cNZIksUObTOair8uIdNGk7
Y4CcDH9bVv5vF0f25OMfrjCmqOuWmUCXT0DyxHZ0H1y/oU+KPdxVS257I/DVprue
gT209ji/qPmdGLcGKbFZE0g4T1KFULtpflraWTd6/xeAmIANpR0T/ViRZXaJc0C6
mbDajsuqTozr+sGsBv7EGS+ubfKLqYZonNKE9oQTrY6+MjfoBXA8v+8bgnj72FYm
dYQC5r9XM9KAPRRINaitrHvFE7QjglOO9iSi0avX8C9lVet8+QUGh3HqkVAC4SOu
yD+/S6sNf9xjrMYv6Nmbj093Y3Ov6dEbeRlR88Ovxc1h0FtYOSF1n6sptJihMz7b
9UucxLhyN6i/3SerCOOQuefVZwibvw/AIDGqAXITEoa250uE8lbKRjRtyL5m9Xl4
U5R8+FjIPAgy2TJ1La645S4EVOeIBpln3sAfwykuE6QeKe/RVNspCeL7FEggzmuh
cBtYKHxZdZ5v+DvLuO0U/xY7aesXfkrjR53hdj8rhd6SEFKaIqjZ1GtqXaUflfn4
EzrYUtfW275cqZReERLId1ZrV1JF8NBeUhJsdAhAsthNQXZzMyj6fxbt92Cnot3E
L9eX/s2nZuiJ2XR1aZQ9iNWE4gLozmbPwhwLBDdj4C6Cjj3ZRo3ns5wky1Jc7Qpy
SqW06R9lxtm6CS93vP7eqL2BX1lDdUu75gAAE+IcheVaH8jS9jaAYeO9axHbFrb9
t5eHZCBWngb4uJdxh6Jb65lJS1RJ650v3kRWx0/mvDbFF5C9xG9FQpvb+UgadSDO
5HuV0gDWCB4dWJYHFBV65EOciFpyfdPR65xCPgK95SoEWcMRkcXDo+Mk3UbfhsHu
WGtRoXM2N0BG8IT4WA/rWkjQ1uhR7GrNaPII2f6CTGi+WzSZMxb06vzvZaJoeyB/
Q5lWVvMZEQBdu6W29qFjI0vzCzTSkxpfbdpEpC4HNT8V8v1Xul0CfeeQ1wMcuaG0
V7rxo/Itm7yo3V2BK1gDDYS2zPNkMrGYCI1B+xQN/gHenN1z3+TOALYLxYHsblQt
B2Js2eMy6ywPdSUIOl3cSAnmTlzC+0OvVPg0hEQOHLFGjm1t2uOHWAa/NbM/kRnC
felWoWJbFY2n1ffqCbHWkBXY5RmZZ5X/zze4WYg+w8BsJJX5Udkm3A8A1clCqjv/
seHIZ5D4vVwjo3zJTnO08urccIXxS528SywAqfj4qGDS7cyUnIuRCSkC2/3fBf/o
cWIB9EIaGJ0vGjwtlnnl3IvxeSFnAViQtAZeI252VtefxgZPLOx/AWBB15CpjtuQ
FAdJ0+PthH9ekk+1KPZmDt3Sb2eZkGrWglxAQVHJkTvXwhxw87U2B8YZomtDlMCM
ofv5j8gI+CBrMtNOEfUBJEVi8obS4e6tLmYpDNGxcUOqK0K9FguPGIpMlP3HKwDH
uhcYGvK/qEVUu4FvR4xTwkmbbKtlEYuRSa9momqV6I+tgyrpZYsxwNujOU/M6DHq
xr/J3B1gluaMpp1NY3SDBWhdRjzsnIRexaz9+Qj2IRghn7HeZAAqL2w1njhmYVKU
f/9WOTNK6PPfpxQl3enKEKbywZtyz7QLjWEv4LcYj/i8yx65/aTuZCwm5E0p1e+g
s3tLg606JXGAXNubvTMxt+T0FACtjV3v8ox9ipjJV7RTHM3uL51zb9DeRF1bQ8Bf
HfBUXicGPmJNgOyGZ7UjaXF7EkvYGFYKqQtQcZKCoUT8ySvJXfGsghD6MGKdecGz
D+kHTtgIxPfjyXNKJ8S3/kyJV4oYdxRukZ8v7UfH5gM6CNjv19ifHULOCbzHR3sm
Pv0/PLdn+9rdr2Zzb/UeVpBYL40JH5rbxzIaTqGQGUjfPvxNn1nQpZp697xjVKAs
3Ocv5uNg4H33J/ebDScvWF7P8pK+9Ht6dFs6+Y9OmTAGjtO+Km5NEZGrCYtKywty
09OKBmji0TldjFXEQRZpg9CUdzQgu9PBlzV25EZIuivw2rJIvzhVB6RChPe+J4bZ
nTCNf/ZdXKpuumEUM9nuUrCaxu13YLLEMjgEE532KWa1OsHZyAXOlywFoybCMkPy
qM9dS4JLBHoNlFZ7ytl2HGtqdMpo4so3aFVGmxfEXkqoEcInAmD6BDRYjt9dLfHf
316WG2Qr3VZn8eDEPO+H9i+t965+iPWmTsbXXb79kQ+CkilABh6jn6cf/CnmBpPG
pw6+mVcIS4XAACMjeUXDykuu30iwDXXIlo138c9OfxzevMEfBpzMQC8EOwwWzhF7
Jku3m5mSloGlk0VArlHYzZQdg/Y7yWi3siHfbLQwsSVM5xNYpCfq7gE9DaEn09E7
oGZEO8t5ebdZmRPhqI5QG6vCC05WaLqviYEo/VvKdvpiINI2wC87o+QVGZeq8akI
/qmLaPBHi+MYWUOU1CGJ4q6dvPXpCWzvs+pukyjBI4814uBA2b7q3uQPVUfgeJDL
hsf09kijMwRDgsH9ze6jDAysdP3MOScceChKnOzlYHpXBLUr6IKTCecckYYOccvC
HN89yIgry703KjVHV19B/+nzXDnPsZS/GAQwHRC841/+47D0Hoczz7UKcz/4owR+
bJFd8sY1mxB1slUYs4hygff+bpsqkMISzgJPNnWgcUvCKkInoVX/4swLE2fZyEk8
YcTzK5NpaxrG1LFetCraIyofroMbO+dNq50noOmD9C1+k7JEeD/rs1SUUbjhd/0O
9341kaGVQJ+Svb584oj3/433rcGJXBEwn/l1CG8Siy2LhFIR6BcKqikCUH49tsPy
nIlP0pk02tBBdLHHj2ihe31BPu/5LwVP4iMVLUBg68GWFsVkB04Ws44+5CKemY+H
kd89l1OtsueXvSDH1vAoNSvL1JeRbNBKa9Mr1U+r2ZvIqtR85k/gtwso4yEAgl28
SOZuNBP6JhDLvqLVhpe6MgwCO1jutg16L6JKPmek6YintqocxSyjW03i+RybOohH
LGtTzwwWkWOy0KQy1Cbr2Z5LBnutKFf9GdguSHNNd0YilKh25FlITVqLRGctPlTb
ohTL20ZhorPbCKxYGYPZ7mFPqQReNRv8Z+K5ufn2JNfy7eCJWASmeTaLVXr3BFhC
uFrJnK80yztD/dbRjJ2zxdrQRHAeHA0lo6QPPzEzhKwhm+izFWNT0tkCgFjyL+IU
5mwCv/D87h2DzUEFUpoxASdF5WkwYKs/zPeVt6FwT6vVyQJEE8vJJkVc10+O6jV6
zZ65pe6G9L+mEYlL4ALtgcKrGds0CN+Pc+7ADIgGKYnnel55SSorw7DJes7ogPsD
24mujzzK/d+te6UEVvMBHDjJ4Oj0b2zEBaPXZbVGjLfw0+aU2ftxw9AUetWUUcUX
+pJTTRRrMMMreEKK6otioEGQWHLU85fix+QbvXxlDL2vdp4HOhaGbFmsxk8lYr7I
sVlyMolJhTET4whp2TTyyzkPEuNGXvnJQA01fOTXUsJHIDX0EfCedxOd3RvoNrfX
nLhGciAEftDiQAuc5sxP1UIQ1xCUkgiZdBfng0uLS6MorTdf8IxaLzMpOJ4DoA4G
v8CR7MLenxK0CVGL3tXZmgVplW6rxbdyzMXzZUpFZO5IuHejoNWeaM6GCBW0B4vi
wVigbtOkMwlGIFWShJ5aLQ/l6+fCC/MnBMCB2xi58ukPy/WVSv0cfoB1HbPlwZYU
9RB2oLhhetvea51PQu65226Q9aHiTrO14/+q9JCHQH3C2I2tXq9SCg2P6LosVfJZ
PsIMOvaCCXAR1OnQr+mXt39G/guJut+oE89k6Ov0RdKqmxt6U4b18gOvVDIlzi6M
ojlQHk7/JLxggikBohSB4P9LXlDQlCbGiTOC35FaruRrt1VHdH7SbjOpLrs2vcY6
JbKYv/xX80JQOX1V+0UVP4hlXxe/vEd73UtZQRIGcvq2uhUj0zUK9msR0p7wqSXf
yrUQIuVsW1uE6DDemZfGzktRxRJ1JFCXLjoq4FB1F/4ppynRNDQCNN2FldG+4BNw
h7vtu/8Abzu5q/UQsIkuLP6gBNlT+5sierCR7S3X93VJDnJgl8/YxaqrkUcJOZKX
7OqlowccMosG80cl5e8npVkg+FHmTAotkCwO/iWn4kaNcNl/GtV3m5kI+9aY9IKz
GEA7LrGwftHwLJJJVnIoKMo4prEqqUwVwbldsRD9h7BzUJGx/DUzDg87mqBhR0ME
EVoBsJ7/py27XOgxfbsw8h9McsleFA5ALz4+UQk/EhDSjVKsJlueNYEaNsK4YwDB
eLKVEFLoVUKTAmaZCruPXfe/0JloDplKJK0jW+07PozJ4o1vQ2oydeWt4Fw/wTpP
HoU4Kd8EOYrpcqih70xmgEn30AoiGyo4jtIY+w/UkVEJBEpMamZQ4cYUjbpf9l8t
o2qLLA2Rxzh8ikXVdlBU1uQHgv9qrSiMQE1e8T1VOC8AIKZKF3jdHTns6Ggw37QG
b9//uDO+xUcsXpN9EnnyjJ8Es5u/tmpiguXVDbrqCz3BUW2u9025fNxYQB2QSqjr
DyjgXoyS3LdKnw0cY0UOQ4DwtIj/QMEW54wDO0vVLZFKryl7EKkU1FAaC7B9miHv
UCWrJcahLeYfmZdafO99qJpUv8EMiNZo37WkQx1NArFBx0FhxoTVajzWnJC1BCdj
3JrlCgK1JA1UswfZ8/kk9jQNgnIJu2UbkQ+qz6h9fuHr0cieVkIxdkaLJOQxzbKf
w3Xs/77nCGtbPrDsmYSromca81Kym+Uan5XrkFVNQMR8RkyobJIr08eSBMYuVg6C
Y3Ta1SC8IKju1fzkfwdM6ctKhzxSDdl9hcJqG5nHkue1dA29XCeoPmG//vXPIXAy
2l/yPb+a82Uj4kF+FlbrnpXOrYRZCzk/N1jE4z6iglyh1wknVMcQlFG7ZOQdwm7q
wIqhewBDTtH69gWNQX7GYYdZyNJyHg2uepRcX4KbbcowteSD/WPDqpMVcizq5b2N
Mn+FGMmz9U7yHBqFzUJODHMZRQ+6l7sICcTxUC1Z79VR0U1Uqp2fpx0iTYb+RUKy
CQu7OfH07FP10b40m4d4MGfqyL52SK1/6+VCMA7Rz+Y0Qtc4c3mwY938jtuy6KCq
ECqRxz9JZWNJC+IZGOrQMW4J8B444N4la9FQyVpIumVFAND/hlG44J/cEmL50vuy
kJUxtdA6OK7A3XLNInOAcB10FZLIVCFizzCLRqH5o0ElvoH4Nac30xaRVGxjEEFI
rM4cu0EXEMP8zpzpaFqin7FGrUtIt2DGxWH2LJ4oR5MiM91w/uWhAvUKyS7ClwBU
6rt3BnPjdjObMeeSZCFnCIHXNrOjULM8uW4YspIaIFJCcCaw174QebtHOP5MBecw
O6dGfhImURk8yTHOCVzs5e7W4xzIGe8nHkpSfBBSwo54UQ5/m1kEFYC6xsojiVdi
HGv3N8GhVsr58lREB5M4CpuKzjwHvyxUPdK+pzL4JIULmBSbIi6RHezR3a1JrQmy
JGvJLRcQ//cjtnQ89ZCbWAqhOzNQsG2JRkDy9SFLCfH8lMdPzPqt6s1oiMyfkXjz
uOCtgifm3otZG+WadlL+TfmJnkfXPQnmFIMRqdwCqR7Q6gBk/hP+drdMu/K6dFsQ
33S6xbrHU+6rEaWIDmXuHnNFDvUjt4aDQ+3rz/5jlkJKcB7EWkPyL1xDwBRrUMYS
5niVA8Ku25cRmSv/gW1/+vKla0Is+pOyWVoER3mkjEiCa6cwvo26b0nNXMhC5IGJ
YPmcZJWG53ueZsx88Y+o90AHHlcI0EPh92w50XokIrk0k8Tmnc2qA9kua70H83PL
s5OZ10JCQzcrgI3arI+fw7Yl3YGJN9LCp0iLSwlCEvhI7sQ7fwBmIkzxoS/ZLzc9
MJcmlflGRmqO9K6o6+JQhdq9PpBhjifYLaMv/yN2YFvGAfQqUnRMdx4gloq48ieA
XL6LXJ+qCB4+RvKqyJCZ/5bl68phULq8olge51EurYdWI7QWPZZKeSa9uqQ+3qGp
iCAJ/bfxkCZhHWAsjd0UJlEEW2e8EMIWp6V36PUZWfC9g4pT8utU1qwi3m9yLPO2
6Uazwr5XBEnG6B77/C5LtP2t+bzr7cSc1g+NbPoLjVpJPThPTzfbipBZ733vYKy9
uSW9VnBUPiAfo8azBgR7uMsFwGAGfK+m3u1+EQssDvuj93kzEI/detrfm246rScA
EWdHWyMPunTDNL7TwwjrNoxzdlqRDbe4jABxoAWkJxNBOxsvqsSns4J3cyjaUfBS
8ykQ8Bq2Thxq/koKcjKH5tzQ0DLh5VoynIEr0ZlzGIpfzuhFqnIpgfeCTJxfZr05
I3yN4LCNRVK/7B31jR4FiroiOF8ePBpoem8KNN3WwuJ5UAa1vOa6iFe6O6VPU6cb
1INr9e+EOv7dW98BuAU1H5aFEWYJrbn6DLGChuLvX3ujLf1YZazho1fngnZ4Prdu
u7GMc2WyjQdAUGxe5xd4JtK9UJc9/jMuN2rx11l+vJ0xpbZIKuYbzhrJzUuL0Rie
zPstqEWEgNm0o1bFEuD541MBXFs8kDKeq7OQs/F8LJLG98hFH7I4KWhD8Y+vXNi6
5jEvEuoCBTrABCkJzTvekHy5xFpxsRPCUAnDifEeaSMvDSUclgEwtN2Pizgq/PAT
cxT6+wrL9uENlgIwVgTP3fAKMO0LSBvfvRPP343w699Aly5mHzLUsJqPOIJ6EDM6
pCsg0tve5J5o9zcaB7pmaQrAT2eQ2dtEMRHajY/DEewjKJDej0+27F0sMSNkoJeO
fVSSQYTz2MjNNh++nLoRnxqgRlRJronlvfVWTbibXichDJoP8hm2R5TVr/gSUbby
0+YDqBnoW15FvwzDsUEoWWBxJyb6MEIHW5HXL93272u9aHo4+ru6zt1Tb+ntgqBN
2YTQoHTRS+RV6SnfoEiHMVGR28aIVciFZoicEkFZ4a1EzNZqE9Zps2KJZXXz95rv
05RYy821RuQ6CblBGy2TemUf0UAsdBVptMpJu2dQbTZ03jw+1Y2aKo6Mr2xVMZxN
7jsLEo2apZ8RBVjjNcOrmpXe6HFjjb9pMY8jAqSIGUs9rcVVX3Jumjq3GwU/gI09
djyUOmacc8pyE9nZ6zvC5eWZ/h5IwpzQukbVY4+4ZpzYLTRmDPLuZ7h9HcdCVgBe
8hrnWaCr6pXv5NKqMv/4xdb55igZfaA/mZski22FVW8c/0vRsP4uq0Hx3/NtAFLF
8pTcDgItUVyWOySKEgmpHsscwt//KTGv2dQwzinZ1SksTw7/wnFaFxSj59EcIjuG
HWr+2OpfxG04t0ny5UQ2jC8xn17dj+HvvQ4SEI9C6WCyCfONZGc4Kcz2ujwzqk56
qSGmi8if0AM7TZAPub8L6baDcp1QjdGySoXLg5uWG+XV3fYejs9kA7W4PlURwPHY
WvpFPLBarfo4zZRpZRXbWO0+l1J4SA3uoLPhlEdmrDi0lBjA+/9iI0T9evCqmcM1
RePN2IILM0eCJqNBNdoWl7G9X9KRo0/lGlN7doeKna+qeqE3GJLO23OMMaK1ZbA3
PXKpM7nSq4mpmFFygRrNqhR/549vVWZgzNWMcn1M48uPybO5YSN8SGLNfnkrSahW
ukF12H2hFwc7QcLVblX534ZYwVHb9FAs5hTis9Fl6Z+Lo/nLGOMDHJw4Fmo47Nyc
SmwQDADyA0HgDErw+uoLnfsAvY06RtxThkPJTm+XgWyjInE+Qd0j7IGd7QlAUoUW
t36Kl8UOAKAMZg8T9NdvzqANPjm1qsl17X0jl0cXFgZQK1HLEr+mCaXEiLMG6L4u
Gkm9KpppgXI7wQGTSWSi1XGJwqT/yvCBWuc1cpdfcvx8yKsPhPKDeUg25VjXJUmb
wUDI0Z8yDA0UMWkjXp9huX56vJpWdmY22OfI3AAcgRxTc0AgkxqgASt+XxmX+4dM
pFN96Mb1/6eoP8fCgtiLrEaflMWa2juvG+CFWlGMEIaOlSwM4VISkNc9wMmEmc3k
ZPplogRUHt87BolUc2ziZr+/Q6aLQOH/hf8y1vzEdhQ6umVEgBEzkQJoVolRa687
sk8RMKvXbSggTmoLYXxqO9TzuZ/eDO4Pg2yn+JI+WztzqXYa5CzbRlJK/JIcUM/m
JCpK2ZHHruLG1zo0npu1aX4InGkPQT3NVeAgzR/68AhvTNxdEjLpw3EGJFb7BUMM
iZ1jbuFU0iC5MEJwk9MTz95j40NbU3RgmrZNl/d3yhYmvkv5kS8Pl6Vhlv/TC+/p
olkILmRdggjYf5Bfd0yqYu4uWchrPHm548VLlQrHmFUH1LgFOfUkDM7esiQYUaBS
wh3IKRW6uBxftBDyG30OW/Nn0ycQsW+gtuTLojRe8azBwJNJ0/ARJYdhdkPiJQrC
1A3414SsUZ2hcWSzbw9d+kVG5nj5DOvHyaac5y8I7E+JYbfvPBTweWc39F7QOLnP
z0meBcV50XqH6m+3iFTRTBWijMwk1+hVnpmUOkDfjPNntewqc3XVS6NwHFIANqjC
d0FQtnwam0Whyf3VkS2YNCGNkda1w3xxdT7OzbNuoglhJm13dK5PJUck+F/gm8Yq
xqdO0E4Wo8oExbJ0IByBkhEXbgVQmAmIyERPVmhWvSBqW2L4uKPfbEq+1itQo5oG
TxybX3yQiOT/6Y07fSB32mfXD1QaJwt8PpMIeilY+i1k0dYCpU5AM88WjrX3bI5L
Y+rlyaBWC4v4Fq2A3hFQ6iWhO6PyqEanuTaZzWz7Cjq0W2P3tZX3+6MxnAno639o
BbI8pWeUG16fsjC/qcZ9ENNmCubNPLkJTGZqirgfb+tRQ6JEFjGrYUgsKeNwQmx6
ZJYVNW++VQjLfKsjVDb1AnHu9tlUKMdM72okeuKrD6zTlaN3nC+y906XY6oXrokQ
Sv2m6ymGpZUraPSkj0hofGW0YbVNv9TZhpiKCu7ddt74kYOTzWU2e9assqgaoa0T
AGp8XnEGqba9scj1A/qKP28X6T8h1pS/Tjg8jgnqzOI9YWWWQKyGZAopLYwXVhBL
zdqoIGmLVuU257kfmnXG/q8HRdCNRq8wVALV0PZXvPbzVqL7KbcoEiXTnrjfL+SH
UdYvPdyHtetO5OcIfAZVEWe9Ot+7kFDvHp0fdlThudq3VHxz/+nlPeyD1e9rF2ru
2tCAbZHT96sJaIAx0faRtu28Sxsv8fOaf44ISj3Pbdrin4hFbj56gMhK3MlHcFkD
kjLaUb+cIKSfPOEhkN5YRV8oyCUhBaYTXcWoXa2cvpw7gmr+pnGkceajRLs6Hd9t
fCmscIDrx35WqSw0By32q1h7gFNVwDRzHJkA4TMn5YeHYTQ2TTes/OFbxYyv2wFu
n78OG+8z41SssUacrsACC5spIkmjbKuIha6mi4QyYZPy8KM8lSopUfZC9ppMei0f
QeWCww6IYoJ0hnggaoop1mGG/1dR6Gqc+9dmvgtMxHcCHOfWcYtkU7zO5dtlusot
OWq0OV4auuUGxi4eDR78BkhNiMQv4JCtMkGosT3zOHLJ04zDcXYljV11TTALSgqy
8XOCWS4AHVyA3Bv4sAjoIOSPdqYxCU8pVPdMP+02DWXgWet3gagSw7vdubXAmFLN
5tqN0itHehByZ1KXTcJ9vKNQ+YsVCYXAM91g++XpDoud/W8sWJ2AJA/rGXg/Bejm
tlG1w91vonBqtqZg15gZMX+t5155mJunJ9Jq9KVQo6181VZb7DmLjsysOWh5rsZp
nVaONPtsI7y8yze/RzQXhVhWzKfEegZ+X3LqeaFqi31woq10Npp97QWPg0JeecpH
iiFFzvq4vvTboT/7CqtacvfpQ2B977LL0zoVk1S3wW+ZzSWDYAJ6d6Ps6Y2qKCi4
N8gzI6EUYAJaeHyC9Nbm/sVVZ+21q/1xXbz3DP1Gqli4WBGVVdZsonNto69riEGT
6A2v/htzRz9m+eyMm/rU7BoJc26Wfx1mt8Ipo6TfuNlNeNeo6Owdz4hiRjF89qMF
aCg6HN65IXhLIbPGbqU0rdHDZF40qcPSlbCwWZZo1rVNDF6tvTbG6+Cz8Lp7k9Gc
8zEgzGuKBX/iGrwo1SYJtbH1QaIUpCuPb3MDUM5OJ2ZzfgZoGq45S59n4dIGUWj/
Es/GlHgbpEko+kl0YSo6pt3U7nbURgNkbNlEf2YloQJZ6WtOopGat5R9SHwgnP3k
UxAqCofC9wC6iQKw0DIBNX8jjMoDCDq78ZlvqsRsPB+0gBkMGOF/qzDA5A8U38x6
mxYggB1EOLjnZZlKV1x0Q2/AA5Zej7FKqN/gw27MhMqU0TAPuvL9z1q1sN2zclum
retuiJ7GwuBH0z/Ix17lrN3Vt4SwFkeUJcA/IpnohMWG48oJ4bWZW4s977qgfqKT
PEPIlPSHVk8JzYb8jXlQ5Pa5egqNYp93Vfngis+OBtCJbTwkLRH1Od4UPBZaG6CN
zyTN9HNTZTAtHqa1TPXBF5U4x5qDX5V0xO/48wzPXJ5k7w0Aei8Q4icPDz1l4lau
0pEjGUMa108mTgbe6OwYgT/CxTXmsRqhuRdISXd/H9x76htqhLWsNiK4ZOFhwt6G
pdlH/cGRff4zhgHIYfsaYBFpja42hvgOJBQWG5AYgdowNC1RIus+AG3RUKJeBRb0
7DX+GLCrGDiHVqlFKZ4wn7X+oyNW2nwe3Sf3Kcq/VVRf+yRvFy3FcuI0IH3JOite
WVH6Thy0fmxRCoebejgBZIkUJ7JSDowldwjPyfiGdPkH+QoJ7S7NLrVNsPTekQ3y
ZpwtJQUTlXVS0POscse+5TRDh2o+rkRnYL+DvURRqMTukHThWycsAX1y4XARtPLW
Hp1msM32daz2OvLKqm4AeNMoLQBMI15PO4emOYWOsZxKZ6rFxzTy2yYtdXwpqZJV
OKKQ7sUJUszIAs4iWZRVQXPhUBwxbnzTzqRT3fuEMEe7Tn/tK5t3/wB7odQWCHyF
lhnSHHBKhaH30r3atoXzutVG5U1qwa/MJvBUmX8VxLSs4Hn2NDNX26Ri4NANwOnF
x3ItqwD8YByzusCe5avxgqbHe7Z7Cqo5DF6koDREz5rIcRcW2MOja5+i8h+nh6qO
pyOabRlGjkfUj7g1gtuVNFnBtkCbND4zlr775L2NuUAL7ozIz3/pBtq1nhiRfdPQ
dXiFI4/o/2WSAdeXbHjDUmmW10jWJyZStxwp0p77KEx5WwW9O+pJ2JEYD6UISvx2
6fYqfln+P1tg61skFOe9kfP5oEQuMIpOEM7TRe5YbOE0GzQv6J+41Em4/4UGFH1O
A1RC34Bw/T9jzETH4DqinaADXjGSIRuXWkV4BU3D3V2CCAZWsEvC0BXhHs0WLUhR
HWtZ7XwtJGdsw66i1OG0oDuZ4v09lD7pvhAtv52Gd/Fa0cHHNdHsOSLrt6h3TnVJ
iXcCxEB8ZjjxG0fpv/198fSFGu8J4qzMD6sDjaLSTlZKpyF83D2FmzFp0wsuUkvG
zEXf54Qz6mHnG+B0ViBya7yO1XQEgdBqyqCwct24HC7/YZJkAbYZdoNL9xpepXQw
9BGmE4qX/HylM9BFrztgrqL9X0pT33nxaExiYqu6rLPNGeOVqj18B0xdmCnUMycN
JzlWzxEGlZdz4LXM0BiPLblJ7mztCBMCJIcBgLcLTBOT1IFj7G+gm/Wt7mirMr+r
/PH7sJhaX36lgPcs5gGzxPZLQmdclszeMScwFYmgWrFZp0QwAU/OymozEu6D0ulu
fJ+GCOhKKDa3/j9XhdNnqZXBuGqdVzM5YicK/oggjn+8AWQXIcLwLjrJyZeydgzc
oyqPcIVZeGiwr3DoiFQbflxE9WZgbBbAkrTFrfBUGaFa6iTdqYKLCep1hQBBGos0
FGB8L+Tvt8L6oGhZtOgGNxhjLgqcBSMmluInn+/RRaFajD3w0S7YKHUj1emOmdml
H3uwJHXaDzvtUgESKVaA5exW/BC0PX8vksxQlK2sPlRd9udQTEIJ9oU1fuNIa2u3
2Dfd/IU4MvRgplHeSi45v+/APrlvYdH22jIIGXlfvSXm6uFUYMZ1jqMjllVgS/cH
4G/tN1ZWDcXGZinhGC+6Q+oc8nkUFd22ibPS0LV7J3lfy33duaSJ8suT/c3hTA/G
eXP/DH6mf2H2eVqE5LL5gPz3RcRb3rtfvDCc94OVtIjIc01z6YjfnJG9QfoJonc+
/NiGFRG0WkIMHKOF5r3PuT+eiYdbLu7TuKkL3t4KnVZhGUKGqwlKAWNQKyAHdOFD
3kyluqSnn/v3YXs6s9ytZFdpAXRBCnxYThMb6Y4jlGlKD1jn/kEstYKqPzITAbW1
KN2DtSel34rjm7JS8vKGLplG+qcoP7UFvhGE4ZoTklTexYCSl1JBZR+1Z7k6aL79
ypshM6RHvQeEkV5zF5dIv200LUs7lh4jf4d2VFnVJIu8kkyfZQG70w5nU1u0gNSu
MxSi03QZV0j/tQUsOysflcbrPRff42iOahXn6iYwn0KDPvT0RiY+1X6zCYFeUxSd
ZTNVMVGPWaOApRW4uZZMj0H1ndWHK9EHG3cWc4bOxEErN7TGCm7DF1TDEyqZvvAH
xuDnGqsfL4JfHaczNpEaw09NjxEuCR94scNi+SLNx1R4L8MDNYy9JuMg3RATkfBK
wxjJL1kq9i9qCZ8lVZNMygG6IiOQUx7XPLlSzmXzcfA8NQMGkkYumwxQtbOg7itg
eZCbL7Dd1Mi5bjDsdr9znYknvqTB/VUyr36LXg9/BHGg51HCowjrMmGAXUp2Bvk9
FqW8y0HZnfe6qtLg4CkIfNr+SRWrbFukp8APhWyozLECiJt4eitE4WUkh5T4Xdde
cFtXk+x/R6AWZI97lHi8IdkFX3zBFrASiSW6j5Ya2tdKrDjJaYQv4hZwqayQHJXw
9HhKeFS1JTs5J0aSa4NFdgH9BPiSMMC7ty02UaKbH324h0F1usUYxSpVKlyz+mRe
8Ojn1tphirKUz8RW4T0I+3fLa2YCaIJO8uSvI3sgpfvYdGOp+knuGDiRab+gx2Rv
vRXROFFXmFukhQV6x+PQE7cR2NSvx6jyzpgtQkmHDN0IFcdk3IOxJZ6U0sMdCLav
X+31+YRjRNHkuedr2AYVpSN5CmbnLgppAdHzyxwA13sj7VFANBYalgAj65+l64VQ
YLB/dMnyS863BnaWwwzwzV5/+N3d0XbLsAL1EZm/RnVUBIVtD2ciPPzVaYGdfblk
bHUPSDErRB+SsA3ftiqEi3j5SVJDE7x9g4eIrp+yScWhdZjmF9bDkpKl9h3ypgnc
vOrzPY5lfrXEexcyWTSAzwn0czwo/vVSBPa5mNiu8DrDpI5DubofQZZlo+Ja7QZW
NVWnCTN1Bqq8N1HXe2xlYbx2R+8DtgudP+9OrzDZeOl4xP/3q4aWuQWSdptfLcMp
c7B/pYpbyrfolijF4KgWKt7TCh4J5Q15XccOpzgt90iIHBW3r6UEc/2Wjzr+2ESG
tfckLsOQoC8sqxFjqqpzpVY8QKfFa+hzMuR3djAI7JL5I2WRjuuY8/0Iit1LfdqS
yI6I8QyNyTUcncJzq/ERuIl9Y+p3gEEwaV8Zil1QZHofwj0vtECjAQjwr20N7aup
h6N09nQUflWVDft8PHmXMckgbQDbsyknLEXlMxV3+WfPDydtWgHi5AomhNqgsYUG
sO8SvHEqkzcQdCqJwLYR+6m0RylMPpj8xMzMxQ/sjJMc9nltPctqxD+uto1TnKcZ
cvdfAO13SC6hcWVj6r/8QFBvAZ/oAHob4b0VnH7hZalVTHTWKxCkhzBS9AoWwqcV
97tMDpSMjM9Qodl4/AsfYRDWM1rj0mX+DX3NzM9Pn0hamjIru5jUNzrGTkIBrhGT
WvNHfXWYie7ggcXBniXaaYSnlyUFS+JtfgYZ+b2m67EoLoS2dheTpCOOtGpCoXC5
Jp4x8w/OEuJXVpTQPPFarMndKzgD9pjbso3aWjiRX7QTYKNiWauA/+eMYIRCpAp5
uCMkzAmtpCCGG8XEld3p+8yLm0dV/MB6bu1/epq+jnDTAX/kif2++DKJTvajicq7
SVgRD+A+0OhhdHapnOfBcNxAYbO/v5Wy34/RH4+JJb0h3LEcmG0CyUY4KrS1+Dh/
ebjalaUYRp8wfZJIzFaYmPcNMj+7ZZC+lFdxrJfRiz/gcAuiRAfX2ZMb6bMx7KM+
vh6k6zRiFtMDcaFJkfwDkuFOXTKT3wY6Sue2jB22w6iiUcvG9J+AoRIAvolPStz+
QymnkbWSMqolwOtii+LWkV5JnNcNQGo2xfSuFFNKSGFDL57pQ0yIBxoUV1lewQ/n
8cQ3k7TLHUpoKjh07n1XpKzyz7nwlgc3ACTBRfc7dJCcrGt0+RRGWPte99KpteiQ
nDawol+tujXqpVh97fjPq9JqOlqKxgzwF9pYQlksStzY0W1CigNxZq8NubunMvt8
D256nacXpQnKj5soFEt4t2ACkO7BKzOH5HnkZT6t0y0EV26bOH2B1u849Ty5OcTm
b3NrYTkkC7i1mfNzJnpBBUDBaV86WId26JvMCyeEjacY35XHG8T+JVtIes/3oJrN
t00dAA5cPOK2NYbmIkKN9x8yl454VSqKReKOz7HcmmPLxYo/QQQul9BnW4im0qwB
hXRm9PbdqEmozrMFAwhN+sjsQD+fyOgT+01GnvrPuHIbFdTbRli/baJuRk6STady
yXVwNtUV0aCm8Y9RAjFZ56LA1D5tMJUcY10T6f4xTGgnHW/J3UngaMRspjqoJMIL
3gCfCWYm+A4d+tSzqZEu5wKB0I5yxBWam2ZhX+7r+2M9Mj/JG51NZiOjxw43qtfw
AUcVqO6C8WtYrC1XeQ7kTxKjw/Qs0VMh0htlHM0uSThJOVTKq9Q/egHc1UO61j52
sQAUgb4w/O7vq4PdT9h8dvbnC3590tybaunFO3hdj0V1x+Wl2GrcZoaGd6+9OdzL
+dxBtCIMGar9VeDhqluU6xjN87RUCEtUyZaOGlXsd9rYNiFUa8MMDqyZCdhurB2I
prEPzJyZuWQOvUeGX4O004rKBecryIqf9KRtkCY03UGMRU9kbirYB4PHMq/2gVfO
LYho08pHhNgyKiKjeLYE37Tz3JYOOvaqXsleLFNbN0fPrLPX97JjMvCfP4QibRYl
c5yT1k+//P0PAowdSZPRbl1/Xl3Jv43C17BuVQLhRtq0PD/OGaHa4XJflYJQ0n2/
tdQfiPLE/6QsIpRhZKBFP0END806aoQSfN2mcpg352956r2a9RPmWTT5RqT4LEbD
H8CvPBm28f60GsB8w0uJSNu0mOf4zf9DvJ28A2M9zSE2vXMflEtsgRFNpjePnW/q
CjxUtVfstbaGfBmZ2fKwrajE1azPcV8KUbZSXMdCc7I6F/+K77HWPy7ofY8puTbI
4njp2JTGNRJ9VkeuSL5bmjPHgIqh6jzMEcaU88K4EEQC33ma4EKMVi0usPq0UWCp
xdKYqfRlyXrs/XPmP8sXvxB/i8BvlyHoWJiEfTsVOZ4bWqI3nzeWZdnY9uS1dDPw
fxAq4QIVRhbzgBzjqDLYiTAtBLbLVHKVuVpLSD1Y0v2QHOFMvR1PCu/ReYEk449m
DELSLnTEosz9+zZoaAUzC22rVJJ3sfqRu/LfIlUl8Gt+Jkwtk3rL4g6czUOeOcFu
TP0yY6cjIo2fG2/tmD03RVlXP0IX9qHYFl6NlSQSKgaCeWStbKjY3ewxRMJKbF65
vugShfMY+LRStUhBRt7WtpWbbZ39ukBkcklmjHbDiEl3R3S0OhcPyqwpr6C6V/Jo
/xGzOwPpvfa+WC/qEJxSyVM5tC5mnpaUC07LjlvAY30rqcagw/P8+ULMliqPwvd8
/yIDoyf0v8a7v/cImtj2ulatWDybMrU8taP3kivR+N47RaqvBAOGsyL0CxIlWpQh
4SvD6AtVgdO0IIxj3i47nvYl45YiKdg+vCltS5a4LKSgiNnd1cQwvWys9/KIuUBa
EPKOddLfWqF1yfJEZ1inWYMIlhNAPFfzXwIVR4yAykbFR7SVs6I/KrGUA50WOgJh
sEQ6Gl9djc2+Cb4DwE9Aj9JewY9eZ576U836FAHKMH4YFK1ULObpa+Bxa1vuU494
CopgNphc+H0YqAVsmK4UGryhta8uJhOB4jka/7QZLvy0W2Xn/6asmaGvj6I9fng+
IsRZ8Dpmid5w4iS6TCiCZUfbHoMjpHX0ds/4f7ar2aWd04asfJFyl2R8x2ZESjjA
q1nmEqzRvMJq9mbZpMxKQIGHzV4YvVFyyoCXJHQwLyI8eId5XRsjFiH8p74fCMDC
vglr03whyx0nlMOI/b1m5z+UsOULXiCuOJEEC4Eqv0LqRneIBwZCQltRwJdu7/t7
bfgwJQes79JD2JWGu1XpkNGss3xKKSgT1tFo5nVs+GJDok7JlQVmq1WVAEHdinVD
uGZ/ebX7cJMBm+xD/aksyGB0SkysZCBTwhDDfucIzCtiw9J7wHHcVd1mVTsaggIw
4I5vmu2BrbZcwN/KPw6dSfxeLwal+jpEHg+bXqxPmQLTzUFFsT1XzuGOh6eeEQLL
bfXr7jkyDlM9+HljxkTGzs9ipnzOxott+XtZ2ak7BoJnaHFpGbx7dVADmyuWdoh5
t++qUk0NXx1wFfXun6Bo5PwCF6Zm2htlJrMhlXmjhvKlWsGauirJekAJ/xwsbmnU
1Jo6dNeJHei1pcauLf5JPgLSLElpgpJmymcWHZaaVebJXVnZSh6ilX1kL+zMvnR6
75S9eSPkXjhQdpejkEmKEC+LYky7o4vU67aF0UvMkxiK58zUSUqgJb9zBn2b/9/S
IHAdCIX3uxy0ESeIl2Iu3KSqYnvRFAA5KOfcJhH96vH65hhyg0vP4Q4suiqHHNHM
cqxkrse1h0Lr0rjmX3pLBbw/1l62HicxaGlIRDhXn15K0GZWhZtlPVxqHteDB+id
7/mk7VbjwX/scBg7F+iGn/WwUF6035/9sZvOo8HZpCbywxi76b/oJQ/c++OY5aEb
b/bYmhKuTBOhaMaM9RLeO2J2fyYXF1do5Rm7iZv7s3rE7MDy76GmgfJjn5jaUUrU
ePOLGaCzmCjxb6+zmFUw9tZUcf0vfDude8AiHtIdRhS1o8KKR9QGtIy6i44JqlGa
mLRDSLSCRFKVUVf7p+zIb+Ofto4urSOfnPbBWGzZUKTKGuJCKmXjMITmXqSkYK3O
Nh51yXlVbiKStjntA/UMWwDNU+w6wtXNMg6NgFiFMwhNEWChnPuHxOLEnPrdxRMc
ehYDgzKQDhi2Uz6/QDnsg4uajfJI9vjNg80wOApaJH1vHCCwA5SlolVEfWlss9OG
0ys75quvs2C/fyzMA6YCVrtCLrby7xwxUN/38EuEkiwPU7KZCTSJGGRpTVJI0XWK
xSz8+SlQpIZgVOM+hdazrz67mCXLkYZUprFPfJlxpx2l+wV/V9kuMqHQ6OOOi2mW
x+TCwgXLoZ34VkIGryj5vyRqzaHVct4HmGmRYOpB+TxoN4nQ/ShuutpLcjzDRk6p
BcEc3IW7zr/5aar/3rQJUgXA+SWfV0I2f0m1bFgWcBoFKPvn+2CayK0pDTGHhVzb
fPJxBZjGRAry+Cv6IpI5DA+9jFRXaGSBQcalDzTHocbn+vNdu1/Y0dLXhRTpY+rE
wX02RnNvc9WnHEVDd0EBUlQL3vae2L8V8yKuajcGcB407LaveRBooT48kjobQgsI
9misFG+GGmoq+RMgS6dGineMpizqncr6CnoHWIykLtGk3nJqDdpyH9SxvlO7DKdy
5XFoqJgqq2DHRClocPEOfMlK3dDdA3ztV4VrWmAv4hTkxXLrkMovz+hZJj5Injkc
OI7UYfqPic1RYEUMg/Dn4fsQM7U+maCHtcq3v6qTD2URCmdBXH4ustM984TzaTle
MH5dxAidEuwpKL5bS02BUsD6DmS69Q1mjBq8UYdOE3/UzifMmIZEWKlfiEcaA/zm
GB7ta/Sfi45o/wJCrtSIDUB00PecNiU3lU+JdONIhwEtoUlDxnz2sCt/wrh2Q94q
xpPRxqatIUqRlwlwDVXTdTOM+KMpggFxiMLlpcyOVcK0F2roj6FuTILYJnkshFEn
i469HRwsDfTG2+Er1rTj4VeUr2G2U+h+/+rRNk+Ok+0+45Jo4XYadWNHmrvaZfoj
BGLcEKOIXsONVItVvobwPNmBHBvcXHrrXM0oGm6eM3Uxull/fNugx4evUcQZZb9I
1hYb0EQyyGUYkjllrizZDNmkD1NTEEXxkzslxWM8XnTxpvBleRMMw1Kn06abNhd7
3hEEA53nDXlEladx9Y/ttuubny9EmhzIpo9N6GfROvaPXz5L8qRX/acikHROFeYT
LTlB0lpTvAc0Bugv5jQPOWkArOkLYTIbf9+MxTuKv+4WI1035Vl7eikiknegKtpn
tiAKAZb2WQ8TeoG2dB1Amx9a9f3G+HQbc6jtTN4MImNK5T6khsjJMKNNg7yEhoyR
bCVyj9Rg394IJ7o87yx4J7bPiZNhSbUShR7jFmQH7Ha8jmNKDfqEuKF3YBCwUekB
AB7ncc71f5y/1ssnnrxPo2PlVGJSXMQRZsct6QtiyJn/vt+879qwGy7tcLnjKIhG
eLZwBZ+vKsUsQyI2PWxMKN966MdBI9r6Sd0Ig/BLc5zLCXr5ZbgT4gbom68ZUYI1
NiJU4YqWBf9IwvMp8d/PEWBwMYtTo84LVt0TO6vPuJWF5Fu0hl3vWxsrT+CSVuYh
M9AFR1oFJ8cMnDeAZ21+llwHn6GnZGDE/MDhRmp8U6wB4L2diB6jXRC3Jr7P5lUb
fVcnver/zGLQHLQkxHFO0C1WQE+jTFSNmLZsFID4MJH+mjyg+pqVeweqduRNl7Cg
ENUdYXY/SkXhGSb7DcBbbdVDdpQB5PLX94e4CfoXE+5Ysd+Du8h+M65cnZfrSGiQ
RGr7BylkU5UVACpVfo5OLeoePndKa2IpHwgyibZmOb9D3uqwYnQOcfxjiYSK5CU7
7Jdv0zb+7XXjX60bfRdVCm3TxBT/nnTBwbtN+EUMAN8KM6nE9HnkN8UFMI9EiAiV
0NfyiOBQJrA563NRrkPFdTThajQRYeFY2gbcp5xQThH5Ly8pKPnrDXeYSfeFlKD4
BAjDDDh44a3TpgbSbgTw4fwUzHzT7KUBI8ZkYeDOYJvgpokePPrTnO/rdspB7lX0
9RpGvEwhLhTbqR5aaLkQLl1FfBYyL7H8pQql42aCoawbHTIvOEZGS3hjr1xJCtzP
xiqgvINXd5ldM4J40Z28QzdCU8/xs5eTP/3JCWIFrX2Q41ceB8gI9/XXsV+oavLF
SKZbRM91DcEddQt1wxmgbJhTY8L3iE3nJC80Pb56oloO0FvDFACUiTuQ9UWSi1K3
+gbyTKxXtDh4xFo6OOrWXUWU18BGuMk7B07tr4Ye8Z5YnSUR1XR1FUUq0luixllO
dA7gY6QclivVt75R1shUkjhLE4dmMeAMAqXDqKFyCQi1X+I11s3oKs5ADu+jei0y
c7l8H1thW+hZ2h7zN2+qIJrojwxK0fG9jPxJp0VTSRevS0OJSNBF4e86ie0PAZqw
iTBRrnWj29yEODEz2JLcRVMX0LoWYsMwB5AobvgPe8p6hGb1SSVrwEWefCvhBkv5
v9K+LiZ5zSl1RWpkHRBw0okMcuRVZUb7LwKK+gUsfNrNC4GpbaryK19WjvMn1oGD
YG271ewbGnyE51SaL+RM4VKjIQkLAqaxD+Fma5luamzXSdWRwzjWhP6yQbEwxE/3
hxIQLg0e4tKJL8wcxfmdxwedvi9i1r6I/IyhpBxjcwaN4c5dB9UZS0/GSS74C/hJ
WlOrHyPLTAqLe14Z6IuPElY1VhUQjXeTU2YKsRVAanKFKKd+Ntz8A6AdlagCRhJ1
jB41OIce4gsmFRZ1WNyxu4Sa2OAcb8EFZWxilLStpbXk4XjIw04adAUqacyT9C16
RItioFMIRWaureaaY5S03GhGzEk3nLxUCFSHAUNgfvfpMT1quEtVGe4ZKVsdp8Eh
1vlyMC+VJ74zQXI7JpCR0H1sGTzmXgPFa3j7IrIgqR3Ner2PrizcUvc46eUbeKSl
j9ZjqzTXi+S2wFE0KkE2X9V8bMAhz7B5+evx0Fu4fuJP1zEiCZ852aw4soQxUOl2
OpRtTg0ZJ73smFVlTaAofs8cRRxPvxdIBdGHYQsLgtyMourgbAdc4TuO695ZD302
LuncyT6bytd4RqHsAuXqww/tJJWczwOqYStqUcY4dJIjqTT+H8naplWi+Mw1S5qv
YYoYjUHIYCqOHOT2d4O1v7AeH9ZVa4ruH7fGsEkkQlriJS87VORyV1z5VcisdjT8
vD6GSffJprLXHddqbaVLufFCwo+G8FXEkSwiXP6lwbKeyl6gG3Fv01dQ9STIhSZp
lBzwusqjLeA3x3iCgGUZ5BxcnWpdQnp5tyaYNlewNdGA2GWnS3kPFUPRoVSX+b3K
ZxoRwsPqfq9qV+L5BOtg7PPqRDtFOcnphEthY1GWp1a8rDRxqJIc0+tzjP3IrzT0
cJK8S///3huIh2W68Yp2T4VAawFCtqgHFx1ZwkdUKkOp93Zbh+WxQdpjZ8Yx6Y0y
15tsvNHWew4YfDHYRnjSMzK7K8/KCsGl00uw41XDIGM8mEoso67n73TS9B5YyHmi
ZJQO3vPxa6L440xZ3Awz1qTMZTXOljAO87Ip0f4WLuBUbL2BBVA1BUtw84H5pTcx
7d7gIOxXncSvuoANA9t/DhP0exYUQVJFamrX/JNXfSjSmNSU2Qe4YrWJ8zXGY/wF
Llo5CGQMKVJR6HZKp51sNWeMc2f+Y1+Xxy8t8W0ae0AP0CqmVSjuIjDc1S20Qn+g
lWct44qa4YK3nSXqpMQw2s4o1fCrM7ysj5+ajund8uUTIMAg9W0MIxFuMcAy6+KS
npXDUCPFBmcTCBQXWhh930gSds0G6gh7ECMq7c3ZRB0jHHvKaHjGsy8CbyOZrnC/
jmOvWySzd93QOykzay4PnaCy5jV8Lp5QVu2baoYLZn4I7hLOXZ0Tup4XGwrYO+hG
vwNTyjs0a0W8IZP8GPlMTE0az3/3B6or7VHWJUPbWHBDxagYET6S3Qj6zdh598Jy
36at9l1QSOe5GncmD8/GoPzgwUykYqC/lcsCHCD/P1XCdCxzRSmzQWJmUDcvUJIG
zg95cyQev0FumSYbO3g3qOivp17d+kzPZlqgvLUxBkqm6f2Frl/9Z9/LdgAkbBcW
5MYCbNcAjX65ETPi2T5z5mP4uRBJo15w8/oqbA1PnKkAGc0kKGlY4p0ZcersBTJX
Bpo8kUsZIn5JfdDfk/eli54t/S+5/8LO5C25V2pAzichPU7TpB8WJaX948JZGb/q
xDZj0hWpsCfLIZugkN2cSrnOzihkohLMv/Rmhxhygkgh4+FZrXOn+APzOMVO47ag
+7UVah1qGnS/Ak+FEUF9+lmnsEiT5h03J+kXUSow/i4Rh3faqzz0yhJi7VQ4OodC
kwVL0STB+y2dPuP9NKmTI+Bh1W9x6gFZu/woCK2Mi1Y/u9wU7Ky4OeGfE9Vr8+E6
UXrcKU4bMTVqW4bs0gH689JOgEZFqeUFDVcX/f5Y/RqFjRQk12B8DdiDoFaXaofh
iQPiyRzSL7yftVnGWevAsLkSrcFHSUJZz9AOk8CpW6lK0pjz3QvrrG0lYpWtqLTI
i+b9vnCtWtFEFtWsS1tNyECTvfnGwFby35o46qcH4zuvZR/S0LomIoyZ8lFcxojg
hPdjiUCb+4srhB+l+y5UcXZ+A8qrc7/Nam+vTkAksVdBIHnsW4hU6IA+dCY4gFcL
4n0orHnfQlhOFsEOg8F0Lhl9gutCm6BJvhyKDMpYItBi9nKo3YNV1Sd8dUcVAN/z
/84TNFMie6zA6Gs+2mydXRLLygb7/NOX8/zUgd9ZnXr8Dg/e7NWrzHhb2OnJNKkN
Iai7ndKaoDiQAMkiQPSRyWY6yVzMu3vSkl5jzrR7bmsNNfYV3SIPbUNuKsMgqME0
yd5DmtcAIuoO4/GS8x56xBT4IOT4Aq7qcBnoqZTY/EJzFYmBIeKy/H2OFTRacat5
Xd1jEdUbQfJWbK7e2FZHcPWMFp+/6LBUd820/mkafMOdnLF2VPnxUYvX/mvFm1/b
T1dCwBqBhnFWWRpYbtIq4KKwFEfF5rIrIVZBBlVNtvi9M8YazTI7mvME6o1lBlnq
UDvfjg9nPmh/ayIODmBc3VXanwBIUNIIJYpG+28qTamj2Jf07KpUkNDKuLI90mHt
xTzDGjL06d82L7YQwBa9ZWg8AYjf8SBMp62bDD/wsgUrFuZAlgyOOPoWM2wroSB+
ZaS4gXbE5kqVC0mB5/xyW9x9dQvwxy1HiBJCJxaR2zIQjj0wwHmc9e6+Lwlxe/+L
GV6TlStzNe5+6JsIDSiu87nXkCWNjpHcNTjFKAIKBNY+TOaZF6bhpIjyTP4l9IW+
JURCT7LP+8HrndeiCCHXy225E7jYo8bMoiAhHvn68N5aP6Hygj7bv2bgSWloN6Os
3gxC8reY8bE9ZgDhWhkQ8DHYqZ2cFSNPMl4uukMX9/Ad+F/z6t/Xl7nkmSZIoKUU
w9gZL4yFajk1sw2upXIhAOuagQX//+1wmqt38/aB66yqwkt1x0g7+pDtwFj8z/Qb
ygMmA8PuBywiTek9+UD5vvtlafh2hYoa2pH4+VGFgBVRsvsBSgdYnbPf9R6eEyCf
6qnfwHnEOMWTv+3M+4HM3xVSnsFfOjtrlGMBJ8G8jsRPfzQ3JPHkayIpJbDMcyLH
yYjfIISsVypl5r4rionj07CJg7KUBmD7eWATAT4nvdmZJon43r+Zng6LoLeXAOGJ
LawOGa82eq6lsCthi/VgjCnuuoLb9+OXx55DIMw/2aNFpLOog9KFkxENK+0uFWP4
TW6+suam082TaI/jxrzZTBmL12yKCAaFSpfSy5T9zQe0m3CWH+9CgxXfURlsJzLH
inaRxyWpGFpvlMDFoagCvYe2YyibiSSmJtjabaUVkvLTKfxEAhoBTIuUdLC72P74
mnrIZch6uEtA/N+0bZly0RA8bmzvodrE49xZaCBoVjA+zdqpkekFi/OkCJjs3jZy
UpwrUfd5MYn4/46CHG/8rseUVAexR3madNHRWPd6D0D4QJpzcswas7ekPAFnwV+Y
R0yEgX3ZwF9uxlDg3ysnF/ql3jriRUVdJkgaOEW8jyk3vtmaJbn1h3F1pXYz/+gm
xjF3Oe4dvSr1hGUBfWqHxHQGfp0b03SB+P6W70RXSCl0FdnweyDTD7GJvzJQXyRf
d+Iu4copyPkMKjI7qndi4znXjoxi1EcbTrfC1oyW20enXYIeD1IyazbXrmBH/cIN
371jEgad2t2Z+Ap9ADpFuSbAW7oC+e3pJ3dmC5Xm9sUEWiy9OMqZURV5+yNnkeJC
QK4QktdRmUGv2Vk0SLC/E+SUozCBa1tNWwqzO2bQyr2OqAkxNsAjvUPO3LSAU5fL
wHDZasoQ9Dj+Cjm0LbDbk75pPSZKLxJ7z4wll4zph0tAPtJ5uqYazgFsghrMATcw
4bjKMJkn2GOgc8JgxKRWzMYgyVNWvVmJX26SH9UGPmhN5ZImddimzhJkk8r3gDej
8YeXuqsHeCJ12cEmXNaTHL4eOVDskjO3pG/IJSqjswVJ1flnpbQMYJacVMmDDivV
puJxDEDxAQxMmsgmZKP7nz1UAkcA8zoDXcK60R/pT+kuFRMQhfCWMJRxkXLTK1K4
rfocQA4HpfHzAEZ+xpWwfUq6gRWc01SQ7wKUY2TIwRQgpOHg0l7o1Sfr/iNP1oAE
aY39tRekFBHVpqZZNTDg486xa9BRDAGWeTfnYjcv3lXkcxrz/BnBIYp02Ci6j6kw
FhxoZd5B5xZGZxWETIifgaKyYzqGrON2JmgeseZferKc93oNeyzNlYUUUBN5YLjU
u/THHPXuDxLXCqdY6nfGemK95/Q2QzKolnK8eBkpulPzunTeVegdN75vZVlJXfIk
EK74lg/pb9Bx0aNGxMSPUz2dZJwzPQk5rg7vi2vSj4tzQzTIyK+dP8NTZFdnJ/vh
/bndRU/rtqTp1RWf0mpJ+AXGeyS9fdAeCnkktI07rIBIfjaaKY1Le0egG4MC2mJ8
5gutEdU+wxF7UOfZx5TcPqKztoHOn/qPA1ORgUF5ddtxX2W/AErziIIfz2DabfpJ
dOVvw45ea+LmvuXqmN6/lm2dx5f5g6CMiRiRVQoqTUI318bLjr/8De1o2yYp0ZMM
SjtcNLwhJT6SalmXVJJiGmVKwzg/3zhWt7vu62s9Y5DgRXcQ9U6+g0aDo6oZUWZL
CXyZ2Xx3Q/VFdfWrVnE94PMtrxsID/fdtiobMPWyjit5roAmRnahY3w3HA7mR468
2whAEKK4Oj3wXioPiRCkZS2lqhFbeeNWG3bsTFd1wGsXHGe/FF76cHHvtA7MB/Rc
MRrerh11lhgQCJipS8z/l+/thSoIMh3NChmKHDK0xYsgOcZoUctw23Tq5VGdKWNz
dxmHTI+/zRQopgd5zOOps4wT6OhDNVpIFWH4LGCDFwUax/TN4tFSkRkRa3ITkFnF
7AY7bcCgaOxK2OoCn6ptyYsx/RqeZ1di6xH+kw5xjDS6Tdra+5U/jxnUVkCjybnT
VcliSZT6MJJOF3fF75juBl+nLzJRSM7ZblJk0yEY+4910Wx1vg9Ynak7LctaU655
CcznikmU/6TEfS8rIz5cwfBJzQU5AGNDP7rm3dqwL2/Uu7306hHAn3W8KhvAf4Xl
ceOMC5Lx8+DmzPlZYt98WdRgiSaHa7IDWbLWfhmNmgJAfsS+EFB5lL4poMeWn9fY
6s5IUip8P8Wb9bqRdu1n+R9wmOaHffYB9d1mACLQcAXzJ6vyXOvTDq02j3KarwMl
sEo6hCutp/nIiODhT12eCBSuoZaX4lQf5QdKMQ1UdH29RhK7xk4mt5hkwwC6iI6/
uV/opNtik2A0kqGHmNpfjHsaXLaUTopz+BzeN/lMdDZtXADCjFq9dtqcKqx8X3lm
/+u0GOye/2g6eQbqQSjtSF5RWGYGJUkfDnuDRilAAriXmxllJHEUO3Arb0c5op4Y
MeCHc1FD5wFJP5ahdIAHp/MJLdUhwhgUTMOGutKP4r1MFcro46OBfEfdHGpPtdN1
sxklx6ldLtTKyz4nIZGv4xh5Pz6/nmr65+Pspqx44J1jI9LvMdeMJNgn7p2pGDUi
2I1IJ16QbtzYqrIqm+RHvDRjgVCe4E9+VhboMawnmC7FNzu+XZ73auaAYhYDVOEJ
bcEqnL0ra9eYr5+GC5ogfNQ12ji88vOAhhQ1qby8xMP00DmCcIplCQ916iJ08R9e
mxBHlGqacToKlytjD3Xx78VDO3ZiQWDpBbWbxf4ynP/cQ5iNFNR1QFNnXEFhCxFn
3QWvtYDcSUoi2EafgHcFGM4U31axno03l6pERill1E60WI941BojJ8Cj9UQKxLJp
ZTscLmko4+tSKEyV939rYqR/zf3vLgZ80L3g3nIx/MbI7qnazQ/94/Gz2st4vLkY
lW+FnRIu4dN6MGz6bZGNDBxLIDZoPNQTK1q8dzJRFKQxQOVgjT8eCw3me5vUbwaD
sRCIfvEkda0K8wAVq7MYIkBRMUcSbVHsSYop3Q2XElCEvqv9hiXYcfLcIXWargJp
RmMlMK5xiYcZhXXcKhV4udCMLvnZDiwgPyms0UHqPo+kqCAZ2BmBVBUkmQdJOyQt
LVwqWVNa+SMG1L/Jkb/fcahfba2j6Mngi3fSZDJme8+cN871HXap4ZOxAAN7WO/a
VfEMbSxbcwXhkvnjoMOO65SWMi7CGCegWbsjOpwuGCHFsJ6b9o3hmNx/ZFPO7V21
6lXJpJf9p3YwmPHOBqKIp6wTrkebsPVAyesqwgYsxZ7UsgQPrVLJsF76Hgahj/90
9LMCnn97c1ww+N98EuFfVO01QSii14lv9j99jl/C8ZrRxdacGCFX1wMGxlwIRuC+
xmyyn1HYpw22q2y6v7KKIme/yb5QHyy5ju6X10JLXfD/vyk3YhydE8TSXZaVdPcO
r9ZRT9MeAGCZlEWsNBHkdlD3DFczUHmt7qIS05T7o4z9Szggw+jeTGStDIkw0nE/
kzRX+WcjY+dZe5amZhp2ZyiD6F64iNpLshJ8jMAmSgn+Fj4jnyQ8jfONtJix7LpI
rP4Ztu0qfHdCAG424XXfsAkbFc2ANY1Arr2s5JO00ORCONO3U6hqFHzw5ID4BOlY
Ow6ubFr7lNZm0WPrvSYtuoDMuGLCe0ChEiz5QcJD+kMIvBD1jXtYmPZUr+8NK/ZQ
HBXCTZD101GAS2Za5sFTapByb+qfxyx5E8MTN1MFQfby8sFODqTWTqwJmVYFGKoi
xVSeJ9a2lhuhNk8iUsaBgeMtb6YjpEfuDWch2enLUGJqZg4BA+dOI2NdmLlIncc8
HJPTp6oHdRQQ4fCMqI0Xjneqh/gfOaHo3fVFeSJhRZzXXdBbb5vCIrWpad0Ncgdy
Xy/vkuP+la1zyCavmmz+RxUdw5QGSEuhJDt12+jOu/37mYXhTpdi1SmKgWWx1aSz
MbNP0ZfDwtq+DNVXvuA4pBwFadfNMQ/92KGiqXtOL7mRP2qWuqJz8OhO8BXYtjYd
672FbFBTtzqkMhVm56cOg6JbSLO0haaMSbNeXVxuEbPmJSF89JjmwT/jOPuW7hlo
3ZWhwQPYU3YwytJA24jNpO6GGfO314xUeQsfsdwNIUk=
`pragma protect end_protected
