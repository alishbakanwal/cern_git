// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:30 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jsE/Keg2UR1n+ChC2YCbbBnSLdWZb8JWBtgIwZpBVh2uCuORirKmQlQYO4KnHB1y
dUz0jK2EfKgWjYwTsxMldgrDbCdmB0of9OesNNnQfvWBSujMfqv2rimji3NbXkw7
wNub97ThJuLk5aiGqmydUxAhf0xLeTnsyki63e4hcvI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21920)
e08DQVZlTTaGmU0+X9++YarCUFEOVE+jCCMzo4tb3QGhPknHs20eKXkSzOcCaU8d
bZN8akYNMvPrKDxXAzT8cVCP7Umib9duQ7CktPxdrL3HUafWgWYHSCSnnoWcpIJi
T3LyTKVlivU6h+SeEmygZ5MB43iOzXmVW+wY5IH03suWeuwUJvuxfd38j+1INw+Y
TSN7rYl9WmR5puXcK1NzwkJNsMXDWHgabQTCUSJbKoThlxfPEVLFqj4cOWSvgsrS
grE79SSwkPsabN5WAvACCyA7Wpm2nphQ6WbOfoOq7SNoboPo9S3uYG5bL+TKwpcu
s5j1Nw5J4w7WqtR5GdTkCCMCVNNtBzQM6byEVqXxGqDiaMsuG0JWG2LiGFYMFaiw
+Y2bApf/iBX1++xE1CM1bDj9fi6jMxufMBxOYpuXXRBgeFKICf6XVok4wxltmh/v
8zDhLUifK4guCZGm9PVeIav9ynO0QG81+pI6b+6yKiDcKO1TkKdy0GRHZgpJye/d
5czq/1iRcEIB4wHNSIJx5K50m7PCyPLRLjPk8v6EO89AY4u5uWgTVycZVdOq++IN
Jmn/piNmrnvedCMVX4ZdwaZlepJEu4atd/A1eYy2jL2FqNe6GLypHg2x2TGTcWOe
W8Fgb5wKHHhYHBBap9Ked5Lrtuzx2V3lB4531jSPmuQbA/4Vo7HnSoCaKKgU+ZTp
0bF/XUbh3wXmYCA/3U65jp3KXhUctTqJ0T9a/zcV0o4WbxoO1gPy7pnB4lXUYPa2
EsWwu8JpRlzUZotlvnoz4bx0GeKQ/NFocmG6f5pMmlc6Tyfw3oSIDZ6cgpv0VGym
uFRcoQxoyC/ErRMwU70Jf80/k9nqZuAA9ilBipRyaoPQqvAnbLtrPLy8zx2bzNri
qMw5F/WYTq5Jr/HYoQkDq26dUsK5IqTrI1SBHL7bonuiR49LwpCTAtLz4nBuKwqV
n5KvQqSvfkTnJlB2PUE/Q5EPjgbX0SG7xHIX3ullPDg3gSpP74Gzs6U6AFt8vmE4
RvUCim+H+CSCczgocMcOLgXwf1Ti/r7fB5LWESIyMh8fdzKbNMCLHoDw/rpDlG4S
FsP4CgzGIC7iTOg2Xl3eQD73pE8xQpNIme8xbTCZC8+yv3yQ5Q8WFwTlnkeuIYI/
c6yktgeMhfgtPPHbJyelZY//bz5m8aMXdHpngJHOHtUdxPU6VO3oDc9xJOUTMEaU
QIUf2Xbc0zybdoUbcXlPz4nSCgxRAE8LOHlb+n4W/kvJ9z2Z5lOzJtMJ6Nj0a69O
OvRzflPimRLlqVwbkSZ+i0uFYTXVG/VtIqj2hN+zAbHQWgt2OLVm3269+bSiQbGS
nf/uGDrtPKfAuLio4Lu0YDFIGV5BVPfrPJPikBHGvfqsxul4ORI33YobjCQidQxw
HBFs0XIZ4dX/Mp8etiuMe4lGV4abvBDPEFYVp31TjIi8mPzzYsztAJ4PTymwZ8Qt
TrpzRk5Dfaj7zNJgcyh9JRc3lv/+VnbHPJR3ZtFq3aS20h5IkhQey8wr1fCktkq7
WMLtnvaHbIEaJZsTCe6BXZ2OUYRrQfE2+suoAn0KpJGJ52mFHQilgXJ17o71n/Sl
xelwVDf5kZt3tpJzraXJOwMGJpCg5lUEWZdnDRaVSrxfbqU7bIOCxu4DRZ/XFLDH
yckUdJD72ghboVMqcSCdqPQg8Rsb9nrM1Zv0aKfQ8qpnyz45dJbrEmGmRsllaJvB
umqP1FrSCrenYchy8O/T5p4NmT4R9NzMqhIQLnTxgXIsAboJg4wqNe9luvFgAu4M
HVy97TRr/rmGxRlLfNpVV0zfx7NP6EeOg5f4y+jKO3QBMetz6TZt2t6SmZi68yZ8
v4r9lxgoCzul8ubse+5Vc3EaeYcmMs+bdFRVSTVUXb+5XuYwNORVdkY8ZZ01oovN
66CRnhSk8XAgIFWL+8g0sswiJ5SRHHPzPRXX7JCfT/Ljmqx6ryQApH7fOJx8PKcs
fbAxrfVIxaCCwIimexoI5/Qh2S2KJ9sD8ntMwY/z1c7yleE18HvpjjXbYCq9TYJ5
9tznv3eNALIEhyf5lHuBVta9DE0+/zi+j6MFGSyiVZ/k1hhZXCUENa7jvrF0nABE
7Ylio7EKNDlVmogHUSgdtXnJPiF/K1G2hpEvVwJC7AOR6U+V7puIAQwco6CHTOVg
AAFkId9y8F7B5c2UVRlW4qab/STMzwfwyQgCsoKrbvWsx76GgRpH5sJm3lCwyDrN
MV4IPyDyxchLaUCrX47T7AGCCe+Bm5C4KYY2KKCSkUgp90YsYqyxQTBa5Bbksy5r
zLEMCHgQ54cfstaRjh5mXjXbSZhdebpjbEYkQkGkUDfsheL+hqN0rQhYTOyaZMG2
Wj4HWzs8HKwKARjRkxIdgJmgMpseQlDr3GRV+t6hL+NZMw640iMEgf/BxtSq7FwA
t9BZE4meVP8vRTqenHHcTdypfTHbjNbtcjmGr44ZDME2I4/OKM6k2tCYhYE6ikog
wUASi3POKdoJabAZ0BKUAR/Mlexk3Y1j2dvhxA6qWEdsaLHa+iiKBI6s6fQWjIeC
FY2/C9Opawft827kNrypZ2X3hWcrTwi+n3iRRTVcffZe4fWaMJNRAfnH5BPMRLEB
I0aVL5LYnKOzdWfgmf+yekQPVCOcBwjtu09mVVmfc4eLNFr0OYqil+iZcDJaZezy
nXXs0Yft96S5Dil6I7hH0CuexfOuWE+XbLexkys8cJFHRGkqO5V/hmYak01ZCobX
Ypfev93+G+u9csh03vkh/EN9F00XxEJK2XF648HHtfK85XviCAVp/ceZ3jZS76UU
7tiscF6uhaxRrPmsB6kIVR0/31pQ0iMF0bDpcbxsdszsHx65fl9QXZIs9vQz7d8W
e9sGw6D4y0vm2eHoUlvRP9xFhwimeiiYd0NVnQof3D8bJbGUxwoZ2R60vAd/TMZQ
zUFfqbckNKmpOoGwqfA2QoK4vJx3J8efpTRZjzFaok0sFeF5bqAN6jy19gUxeX/M
KhvoCrxDdfMjCvgPRGjGoKUF6Z0XZ2ISnT0hHuIHJWuw/v0AZVP363bC6Wwhh2dM
+/APV1nFKgicyS20/xXjrKFGV80aICNPzXGEQQlNql4vBLHufrYnSauI+okL5cbr
AUThKsgg3SrMLEBTGrfVAHcutTAupORgK+KAdWdaYjsSh62PHWvNOHon2rm/BlQj
Zqt19WA7PfMjXlyX7Z2S5GX38a5TP9UQVmpwvqm/sx9pzTxgZWFc2ib/8v/JQdEo
+SDZfGL5+k1Lxlp8EDrfCrSF2dVUWlOP7ekaalM06r3osk8xCEXi/6o6Ew1b7YNL
d6BLnocTTc0tiEQsA1/CA1uFuVteic/bxJY0DEaNlaXpH78tyvbLI3JPXj503MKl
ZYyzlaSCooq7gLPGpbml2autgswvTCWSu7FWyyNtJ4e026LQ21h6wp7m733if83X
EF2cYDe/numJV/m8clFIrmn+R/5Ok4CNbWnDpkrQzDXbv/XQltYvFKAeB/cLtUeB
isLdaM0dF15tvz9hZn3TWzvQKun7zjRGaDE7uN7DRt9p9vGh0y3tTXtI4ddrTgaS
sWmCTSJgq0Sne47G5hf4hyJqNs0CTwVDUKk7weQ9iSo42Qs5yGkJXywEBBua1Zdu
sQXJh9RIAor+2xjbXPkNQ1Y0GtxAiVBKksZxZwn5lqvnEuEgkV86tgTG9+jeV4oy
ik9J7f4u03UddW2gpf3C5dZXYIe9kOWadlKZ42O7sTa6kb72X3Z9mBVRR1FJKIEx
fRaJwSGKfBKGA3YczA+4qbmH3SgP5QJ/9qHbDkCejMFPH7p5s1wc8y2PiLdr6Phj
oc+flLcL324/i1sS3T4oReuEXIvTBd//OM1G8PQOV7abacAZcAGRs4HvExnAzQWV
z6pIH3DcNuZDYPuvRLqaILjtar3C6rwz/qQUM+nHt8pdUcswuW10KqjuNqPdmFei
pOAszXRb52ySTpZ81W6IoEEvKN7gzEsX/4/qX6OG7EcGH3KylIyIZaWUU6rUNHf8
zBMa57dM35fzrTn++i28xI1X1pGGt3Ku/8miZIMnqdujoHboKhV3nsQCihwUeWJE
mPvTkzqP9uTT516a6vY3+y6lVuqgSgR30zynTy/vg+dwtrAYk2Xomov3Lok5j8gX
3QqtHTL/uc9PyCPzBzmDGS3PsfeD7hojp0z0wxvKh3SzIAmG6pBSKB+7r/n21sfq
MXU2xWV77lUk9XYz62UwH2NT8c4mwkPZtvV+vV8y7bcCu54ImF/kDQg9P9EHsobv
mL+/25RLUntMaq2nLCrdAaaYoWzitNFqEaViEEm83KYNQqX8S0SfMCZ7mdKBc+wQ
dtoAiTsouHzBGgt+dhb4AGHHjD5oI+TVqCqS2KhlkrIhqVzK7TSqkmHN3yJLqCU6
gP+tjQqzxDPPcsjSaUQIqM9OBxnDMtT0TrpEe9VWxh+sHxUPI+odUB41pFnyWt8U
wbiDxFd3/CkIz08Yni+ZuMPDDERE97vFV6R7jSipFuUWpobtOZVQBbrRkNeGEFJp
RUBcUtO/ZVZt5huRDbYv4j9fa688V7Chq8BhAxwh+cQMCzdomz6ZQbpaujACc2Do
ODqdDa30L2wMRCsv+AyGp5ZvWbPSgKxh3GwXLYCaR2yPGVwowIjf+2W0EGYEbKBK
rSFFTZjWqOTrdzf1aR06lBCZ2TwQ7TxoKU/rrhggqk2Zc2A/oQBmuXYip+52amOj
+6lpOsiRK2u2JWHZxiXzsAyFVBlKb6HT56ZYi/JezBB7KEa2dn1Y9+2ZCFbfPBso
dafNPWrH6mKVee06XdGEtZ4pTatt6rbh/n/bdelz4JBn7zeYY0+ZkvX4LxfpqJiQ
S7WZVm0afJ/301i9OZ/LBDslgbut0CPgQ4vlUpSZXbKQBxMnGvtF3BKuBYl0SECP
AX/t20r7GelOSucjKa2+2piNtr1xtAh7hOgM2COHw8doiS8f7DMAyF00cJn9Q+/x
VTeaNdyXIqJkUQhW2STRLXFyYeI/bzs7LUqjBgLPE69i5QQftEsSowOYryGqtoFC
3XC219+DjvCTuVbFpHEN7kRqIYmZRt6BVpUHtvCgFPpf+Ahkm0Fc/mWAUmg5BQKF
/a9gf8Y1Av9iLiB4nJu4+xOiiEVBLO40HgA9cXwuYO2XpIVVkLyAVR94ts1FsuEH
3TxFPM7J+aeXdOz2XN9OUigHWSVFqacYeUzgEITkNvAhn032fBIzn2eSDgqrLEV4
34fDFkOLozW89TD+ulRdeXntfZZxkIwVnoRMyhw+vP7jQ3dsVdn3yvhJ/wojlzYp
DOAjQ4xKcJU9x7+t7s14QiM2p5QfCoj0KnKREK/8WO1MnM8LiPhYHyWR3kpxE12t
VyqotUvJNIFge9gJkszY6J3TQxvSUzXinJ4a/xKYzLdHJSR3cWOTnxRTlqGelIJt
tJPYG8rSaiizk87gVGKiBBt/5b4JaPe6JWZ5xpUy0679Midr5tgVFQ6tI7g+p4+N
EUdb3+rpR1jGkMMnSFkIxtguX71wmUfNkdyYeex2wbTX3I3PBYZ0lWvvSkACR2pK
3w8GjZXpmZ1Uu3kV7MZrCGBGqrB6RNcORbW1pXOOiSLKGaP/coU+gHSEQKw2Fjuq
PUkVmDrQnRxa5mwA8dasEtkE36mCI0KJlXctinpyF6/OeW6Q7aYYWClPJjePLII0
hs6Ib1BCotcBqTW15+7auMzeZCVJ5oGQ9x5rlW7EVodEpabKZlIMDyHM6xNB2YiX
40hgUi/JbJWkFZU5IGUJAieG3Xs2LxhdO3P9aPzHRkcZHSksgdx3yl8GZtjT8l+r
lIFMnC5l42r/YjGAbTSy76WgKQnLN9glU/OfejzaP2CAykBxeLnrdztS1sqp5e6G
QMf2hSFeWEdP97u6T4il7d955I7mxZYeBAVzws4F6c0oOzpmtTfFYW8pc7TK7qF7
k8V8NrZv/6DevA+xd6elsozEzzDaZAxOgyLlYOLatXuO04zsU2vZwmsT0HcyNd6O
ai9xOAsMuu0j6lsxAK7nzhhPwFxpGiaqNTgJiQSA63KI3ys991C0VggkcuJgobnx
Vm/jz0AMgSJKHnhhBfiMk3bpWocZqeUPwZjk8OEANSv4r9xhncYgfasd8DvMv7M7
za97frkoK1ZpfyVGgBfwLnfiD7UhoAo9NFFwHYO/EliSDGz7IXrke6M7dD0dbIH4
TAhyHV9IJ+RGDYvPgkVoG2DF+QLf4+hihFikS+l3QDEBWUoUbS6QL2Jac/Dz7Y+A
BgWWosZQ2bzhFBDGTrmQPEOhNjb6ZcqOZXRdkQFyhhvrmcm4sKPehiScD+NAYvxu
oYFd7JLurJmypWrwWL9AdTXTiBuQ7H/wynq+BcCX8rjmwbvpfe0thZzn3gnWzqpl
wJuryudQgp85Cy3V/T1YtEYhh5Z7wzuPSypWUbx+BE/1RX59KtJ11X8I/BVHtzer
EaE5ApGw/AKf7IrO6DEvQi/oq7ShfW06IG8oE0q267Z/n7g5vc3/GUWNniXscBdM
q0k8CDl2tc68QSYqHHL4dMDlhlk2iJ46uwE6MBJeQvxzYeX7T/NbP4SAy0nQupxL
bB/cgeGRmNRxxCQQbD4v1uRM6BCkDnWCqqy64HGuj8UshiEc3sQeklG3bqOAHQe6
1Kdln5oqLvB6psiw0c216ZGwbW2W2ZtY0180ZHBpTwI2r4BpCr3QLoOBj6jl0jX8
z9vmNN0+LFYlLHfix00LkuWjG7/q4OoV8hC7Vd1ufXXoN8qyTjTZnyBRBzqMPiJW
eBKcGpoBKKePHJmdjrxcgHRgp2j7nJHOBVIUykNcRMCJx4tWO9OhGsLLjL1JLh4J
awPn8PlzOjtqoa5L3lpQiTBGRoorvvLQ7f6LqsmKuRIQ3shqajAoq60okfgoezsX
9cIKsLZ8LNufX6UCFOnM3dV6jgJX7QPC9sUYDX+zdOk1yrdMScCSwWiN+zCHAU0y
B6Zy4iWVbTA8Iue5EX7lBAbmfTVVxyUIV1pwcCel158hohAZSebB1q+drVHbFAcz
nybttPZ0ACKtn8laYtBFTSylg1nUose/HKrZOC4xSPaJhFtuMeXsdDiUBDkp/Fv/
dW6yGMp5aBgukLnwBUfsLz64jP9j/qGH7Jf4RWPQ2fj7CfN7wVEqiBaXFPQpysWk
0DMVqN1m+SdCI+V44vCcP5aZg6GKDuitmYeaOeiHBE6SutIjpYWspDPwjCW6duAU
GKhp71i4FF9T6W5ynUEtXV3qAA78wqYTy4EZPOGg6NKhL7/FZtzNUwZS2MkuCY5D
qkkXs0h3afbV2iqnqSi/O+WpeKNiCYBUUGTJKQPehkwbsDwEbNi88QV5+JcIn9b3
55XJFDpJK8sAAZDAYBylS1phadZwbiNYOrpqfzCoK8Vx9hO06tLXh+L8UIWm7Z/I
PPVTXRqsv/CiYmiT4zhQpnHVILf26RvZh1+D7kdRLXNyqlk0EtW3uJEQ7PW4F+kA
7Zhf+k5ecTpq7hdeLHnIzZ6VwyLCAzTGnBYzPI6plaNuU53Nfe5ehfo+jVHdWy83
0CreMsJ4PEfoilRUzrjfKdrXOnkHmxSiyI2p4FdhVtALY/NDmIBC6W5hqEt1j+Vb
j9JvKK3YOCrvA2bz3Z5rLCzgelhYialdMTbZA9yOYw7sOx5nYS9SPJR8vKqyuakt
uX1IxyHypxxYdzNxgC1csDmUaRprHdn/Qb+arRjMi1dFcGzjVouUbyyui8RwQ3hG
SxcS7Tu0ZSAEGj2Fr/i3k0h91bC2ses3hWNNG4DmZh1gSjPfmQ3XSjykfCu0xdjv
iL4ORbigDXZzG7gwO+hKU/mluA1kiUmQOw+Spq/ITuMR0Lr3eDTe9bCI3ERR7JPF
Zp8VL2qCAyk/NAAJzq3yIdubeRgjckfGog6L80TTz9L0SzJbXRgS9kIqIUklZYE2
fe9fiHQvF3wjvJBYv8WDBT+sgmyWMUaZsvArE3mPPKkTanfPCilhHYHyD6eMeBjn
0EirHAIKtjfGTtyuUbS0kdcKdlmiHZ5E49GF0ARGtc8ffS55eZSAbsVAI/YwkniZ
11VME6SWpCI954CxIvxAp5sgdmDzeLBgi2iTpl40QU5CqXqBoihuEjdBoe17WjbR
Hk2/hbymzFjaq3rZLZ5KA/uj1iX7xchkbP1ltVgwxT5YG2UA0FpkjheyCCg3KcXy
QqYoUof3TkxOG/WDlqx6Y4jGev14UGJJ6/zR6OfLTWkdv2KuhGxSaIbS7SboP7w9
EiYnttbvzRx2woodp0QAuQ9E2f0T3KyA/Ot9fwE59hJuuvG5YJGSOrz5xF/35SGD
1EsmSkkaFFFoF9rbWKfIric1qxDQLEg7pMqxT94eLuWuqCX6JuVdFmPogZ+OnqMK
mMRS6UPhRoRlbrFQ56XtJEfaBf5MGJW/joPXP6IZ00DpAoSm+KB/LtyQE7d4yrFC
6NBKhPtPTJiQ1gEc4rzA9d+aOHAJwTAeHgBrMWDkma/d+FE7YKu78NYDTOCRO8rZ
4HOV8aI9k+qYvssCEVW4BiDrO6Wjaso69fgTFAsVZ5X2UkbiRAr1+BWxJIVGtve/
7CvJutRo400ZtnMisWtuCXyWh3jBYA4ZZh5ozP/Ff8NNmHd00Uo2F4eLP02ibXy0
P5rqwAfUW3K7BYjQeI4qNXa+7sIPj5fIfwqoWyEQc1fEQ7WAxza7qThdwh/TUVqB
rcq+jZhtYlAN8XXtyiEgyXfRiA0tWldBhLpILNUEA/jb9LG891PkB/9X0KHEfeZT
LiIB0Y30E74N559vLZuT08OVJUf7NskxzQxZFnjBTOjvTpb2FznhOBd6SaHbYan8
viE5oIE1PkHFihJ/YenAdWjTP5DdpPNtMcgyVdJ+28dJNjxeOVz9++WgYYFCRP0v
iuGyzadtql6fN/gH1MxL615+LGYgHRj2/0AGEkFwvoRzu2XBJfd7SLeGEc7ERVDp
IgDYjvZCIQ7U9e027Fk6IufelEPVYAzyPt/CXkEOYTKivUy1Azpu4Z9IW1K5MUo4
SS2kzIJECaO5CezrKf8yr8XUti0+/3R9O69Ttv2rj1XKjVnlggZjscsjctWSFNCq
5ZIVSfk/2gHh7S3LYp/LSpHuvLoY7lNv0lGVOzCuEQeJBexWSm/f/POzA6ISu+Pg
Snt1xLgJnKliXehGRAKXcEM67DhWU/LBrL38+bYxq1Z8gZx3QJz/LadStcRlVr2C
+E/Ybuw+M/sJ2IfSVVsmvb6t9DQ/8h/KvSVM+38pSA20L2mtOYDnrB93D2kjhdtL
nGnRPMpT5u/UIRy9oTIuc52/aJXLWtt1888pMZy+m0NJw/M42GOwwrQWPumPaCU6
LQ8KWDbb9oo6fGJviXU92BJt2QD9Bzc13JeW0ePs5iQFJgn5nkEEf8lgaufnGn52
45+bIXZJI7Wzof2Udj9yDyVO1DOFnPtapa7pUFtd56q/t6E+70ZmDIKNxrXc5P3C
7DBWyVWasLZe+Rxx2GQvPAzLT/TNF0TaFSF5B3c7+npojBeNEKK8BT7rbCXRe8ZW
JifWSa44K4epzy0NU87r9BH4JqqnqIVWPkTkbXSgrvjYbU74jIk71Ao7e7J1SiTQ
KW5KRxw9i/bxbHu6UqNBONjvSgNDO1MgeVpEThHluuiXs9G7KhRJ9DGIuD4Ry1sw
JSnsbdbQYTeKlaL9Rdw9p7jjnnQrldtQxCxtKLzQ0hr2s6Oao/YHup1FBu1GWfN+
/anwZeUgfODT+5ODL+8WrUWyAUZH26ByIzTclJjift3rNsx/UgD/qh8N1jnsXj2H
Ai1PWF0zEtONotzaFv7B09RTaDo1Yl+u8V71H5dXMv/dEAqI4J1GG9Ygozo8PrkH
U1IzqdxemIBVyEg+apOS3TS61I+97ggBo0Gbycu0asKKAEgoGx3QoCdgXp52Qr/e
KdA01+EWj0RyUQoeGDV4jAJ9ZcCKhJUB2/t5mx/D+U8pAUYovTpx2HotgZc4YifL
BrnAlFMeBeEsaWyGveewfbraZ4Gta97w/uSmFPbzAzF3jEpoDqG/Z/5BJRF9rVWW
8AgUwEPpswJYEMppK30Vh6kckrx7tpKWH3aRPIpXyoR2kQl5VDc3nWruLhfn/usR
aJFf0zMbR4jo3rbVMKUMH6RMNnbU6FosHwhgJzScBu6rWyr7cNldBHKNjCIA+s8j
b2Jn5YK8ykKUJ7UwqClw85fSjlSsn75J7P/vcrVKuQlQIppa/yzCo21oJedF0SF9
VBL0toHCZDNAurNf4kIF/gn2gH1g5Bm5wFjTCnJPtvMUg+UmxfpLT0s2Gk7LW530
aPyRQszZb9IOgO56ReEgYXm5BPQHW8JNvqd8lrqtp0S1u+GqzBLlCgb2LGnsAcRe
rm0g0bijTVZFHoNEZulB/RvR4VNPQvEtciQpnvC2AIPmK08M/KjGYeP1dqziipGx
N+i30bLWNhvZQAAc2JF7H04xMslRzue4LyWqnklmU7ONLxRS+lUOdeLDYMPQLJyn
tRY/DnirqEPJVvXbVv9MVNAxcItc3TmnxqrLwgq2p5GJJCwck4woelGjU7AfBNge
0goLTSJI+14U1K+oLfzQmSIUdSSE+t6dMVPtAc0Evv70a25aTSDVm8323Xey0POe
XfljwBztFfi8wx+vhwDqOWAPAZ6UNKKISEoorhCJpPu/nQfrM1yAZkiAFrdq4km2
LsrI8Edfc+AWfM+T/ZUM5TAgQ/vUkSfXA+UQGDxc6wDiEamX0zfK7sWIhFpkKkDA
tP0wyLEUkbxIpjArzFB8ydFWICuC8WR929ke8isJAc++giM++B5khEyjN9GvbRuv
7HM6FLgQCQkhpPCIg2j/Kc/g0UHRkN40FT2oJhe55SDS8Rw0IiMiR3KrP88umXZM
Tb1o/b1tOpt6G8EXqLas0z2W61w7n8o5XPyRPWW7BmsqJQ43AYDEGZ4PHN4K4323
pPlOda97zAJT6cBabcj7g7CvMGmtl88RBHxziypJRLcbWeF9QjsDld6YUuKbc1pN
wif1i4pPgNgmulPFWGjXCOCzf8iOMaKfgnPxf7svar5qlp2hGUcg0GGMWgzwT1Gd
iNeeYBNHjOgaIMrxWwW5T98T0wOKpixQQAkvgzI8ds2cghz/UVzcVZjwyhOPU6UY
xeQ2jAg5AcXYCF6N7sjJbeoWBRJdkY4tGfgjcG4P1rX+fkhBhmYKD3cf2eJOG0JC
n5mbuftXd05z2zqdNmZCi8krxVIG8tT2P7cSpPsGdSsfO9b7u5zkzt6S39XPlhXI
8/l+RLBUne9hRXSWzFjpBeX6uw3Za9NuV0BwcjTCiHTScOgYMP5fRhy0qwq6GEKg
WvVbDjs8PNoB2DqD2P2wGjFVW1RPH/XdFj/3lTwJjHnjeNg9zifEPmeeFbN0hffo
5sVw5E7t+N0DwmOOfrsLmc/3RqTiflIMO7DCh94b8pmiXvckOY6jszAfwk+enPcr
O18Hy1KWohtyGEeet2HAPXMXTa8KI2fye2HuxqwRoJjNjZekShUs0lBJR2u3OLsZ
mOtDW5fZM47I09TN5HjXzeRESbfNdqnUYl+SpyY1RjlFdUfIPuqdJVvW7kFU5D1a
45pVWIzp+wcjFGJ1u7V0R3AAlLdJwUH3KhEbzDEnOstVRYpp0JSRm0+mVOrGxKeR
V12OuFES6vkt4GyCFB/gqXL6pxoAeC/8VdYxdm8/adxX+k8cMjUq+Qtk8D9sXsJO
/vxUP48y1hUKuptInfFY6IXB2jd9Acx9ZPZfhxaR7uvHSScsjmXLEZPHSjBrag1v
epEkCz+E4i55hNVqqpwcHu8yoBHBSbFzwfixp8VREO4jo28ZhNgEhTt6+smT9hZ9
yZ/wyQCsR1Q4LmTbY99q+NYDvpJ37igqMTQSHzotyqMiXNymYd78U6RvbwF7YDdp
kC6/jV5LGZxiDU2VSpJxqbbtJf6apN0nvrJwDHxTODpkp7np2IjCTGpFL3DrWYio
r0SMgET4vIBZ+69KFS8katVKF2T6W/y8X5SH9JHfEu6j1DlMt8mfV4K/VqWLmgU9
ToMMGp0tUB2ZeY6GQ1mWpQldv2Hmvsz1o5XuaFJfzEKHoy1kl9ulNL/q2CKc7ajA
0ylskTqIFb2KNAJDO2r4tKPUDfQ9MGjGI8K/n7QbbsE6FAanxpz+f1knjY+o1+Sb
9aaxGZPU0DagXWemxf6zuIs00utaVYAamMwPO0DIXYHBDrc1ADnUwh4kEH0OAtx9
F7u9yaemPnhjUXany6f0xNaB7BJ5Hkf/H9sAri5WjLFi3VRQHhyVJOQ6ec9wn6SI
8lQfkZceeiOub6oJMtkdQHxuuaMgzmDPVPRNs7r+LswwD+pjn8VgI6+50UIhp7BQ
oy1kOgQGlwsLhVdVzfrCI8CFoecQf9LjRalQ793llTUv9ubIkyvdQi1fTxHxJK34
BqCF2rkgwOMwTcDziVVe+03bGYFTT50EmwPJ7kVTIwr5ukie9O6RnWdZ5Q2stoJP
F1dYdJo1ot+VsB2CAaR0dytloswcGUx+mhfaYQ4OhmZh4T3O46ggCaZRQyn0uME1
UpsWpN+cbj+D2bE73Wqrpv/8gf9ow+UBHpGF9QpPzbzgqc634w4Znqbn1+J+F3Iq
IVc9TA98kkbg8SSWLup4ujC2tuN9anD510lG1ZUj3D4Di2djQEgKW0/MWKkz2NH8
9jwMZlvUSLh8CWbgr6gYfOzHWYpvRtfZ9/Y0m6pd/ZAN8SH+jcY2H99qx4MqLvsw
zok04Yb8izeGBwVRGTJ615OJdXiX2omWVCL7xnQSNO/a4/UPBdcrFs/QduGnYJWj
5+/8ochBN5SVv8jBi9HN6p09YnJA1f7bGxqfS3ImYmacJdGx1EuLSzQZb8aFLU1p
mCvmifHQnXz7ay3OM/Xx/PNlClWDv6Pa+eYG09BuY9qEoIztKd7zuKdnqOeZRq1x
x2awiirNFZQHyxHVbLtYKMLceYD/foup/Z/gtVWwmfZy2QclZkr6FAsvzgz6YgoC
TBfyHmZodR50cmSWa0H9ducR/M5gxelPYgUNLqCyLNYHLxwV3jNpFtgg/YqfA9e8
pbl24Ut3tQjgu7Hj+ASc37Xv9rLpmDCGHKfuyhB/W1ANXdhcpXLl2IMBwCbS1evW
Ep4T36MhACjTEMjzEMqQ7LXA3BxEiIAzOdB0E+LpZI4WeoLVDrAjh4nDGUR1xxcm
OG+387VHT9JtrzXU+08J65EFodFyBXjOJMMnfnSo65oXRHc5q99c8VEi2ryj4uru
9ibtrxwcWjfaZiD9RtvoPiPc0z/egtrH6qJJS1Rz7coJATRiq7IgHjA8L0d4XKSn
+GKTD+5bDGf1jNcNnSGZwv5mfi1sAGwj7qjoAhJ+rIFuKb1YNhvAC2qLkxlw+GmA
APU7NQRvlqe7XY7Vq9Ray5MnlyfhsLS1dYIalEbU+u3avw8t9SEHm6t+lgCNoNVd
fagaTIDjOF/WaodnqW99WDc+k3qd9b/XSsLIWc2QVxIktutIbi8KjVjixAAErkPF
hpl2FRAKkVRAD3zRjr6asE1cxMF5MhE6aoyk5W2CnywdmFi14l6oNk4V9P3JzWBO
x6zqOkJoP83ny2knV+3PiPqny8bQceZkvqbSDEpGijqTTYUibm7n9nopKMjhhcFt
fwLgTDSTrhVwk0w+SMcBotRnt402OwNUt94/HxCYh6/cen6bWMk8w0bzUEaVQbOJ
k6Y8TkBGl92caQp+zhAn/1QyJqDagn7qMJwS+eVgspTh8Tud1jkYKs84YX2Wsi9b
KiLLr43Ihp6yuui8oWjRZkNVPtNpUFJNcPbiwmwzy4NBa2t3ICWgNRvPbUnMYxoi
LB9pvGawmll5SEGaXhVpJVG0fReRXvnWXYsU7ByT5GvGGl/n771Fx5ha4N7KeMnZ
baLGxPaByMchUXm6REKUEhCIktTjBoGBVrI2hnIgByhqC674dI/jE4I92a/l9BpI
4EoPIGl6te5ANcZmQHMpis7+jcKQ8bR8guv0gL9ZwQ4urgT7laRiy1xG4Br7RE6h
FY6t57+pIn1ssWVaupl82h1omUoowQYXJSJ0UBFdIUk0Qz1msFgmttUwnz8l+2NT
hmiz9XLoH0ZKPH9fUUEVwRhaemxd+24p0C4QSj1JL5fRmcnYXALR7xIx9d+VGcpn
RZNMB5RIZfASN9g1xifYc3d7K9q0mo224gyldvd/ibyQPM8079P5NPOvBRpx2QjT
+BVUWnw/spUOpTf55xIrHOKVmhsq7+F9ECLGKWAyGPmwq90FXAcgkAw1488vpTMI
2e0d4D4xqxWj8oTLuazVvN1QzmGi4W3l1DOBbNqzrA3e66RNgF0cJ6NrPhfVgl6D
Etvz8pDGrdFQHyz72ANUYcMTx+q9aMRT6QirfMW9UO1iEuWnWX6ubcULjxM3q7aj
F8f+FoYFyiK0DFAKUXw7e4YHddK+WDkE9cY8t7mQJFyVM7KWaovkZJF0ettfZLHZ
Esm1FbqBXmm/0zgnapZYD+rk9ucfMuxr2lVQBgV9oX7vmE8HrhOMyj2hKGk9ru77
OYhq9en+wiqv8gixlUlikXHZZ+NsxneOX22fD1mpu+41229m8wda65ktIuAIdtFU
MEGSG61tJDm+38NC9NqJ6f3JOmsJcCoE1lQQ2rjJ1At4Fv6XjcFk3XCeDi2ttNQb
pzdPKcMX7RzhP5k5f4V9PVGXxYOQy+A9VdY1oJZ4GfL9keGZ+6ImH58NCF1LGS0+
giCEbQr0pqpQxLlsY3C7GcL4jTI98PKxvJkkuidcBkpkhbcwnO43VENCJ6D076d+
JuRzgdQHmL+MErPBdDscQsj9YWXTMMR0kDmib8mOrvFbvcZjOvvTREQ8WllKbdYv
oh3jji7FH0fDxBilX4ke1DD15hC2/OrWv1mZrmnnLJ0g8pUmDTDc9h9y+20jjkrk
Wf/kcydT3jDRUL4B7VhYMQT98v7At21ZvkqeipIUrojXeh4fhzLxNBYJIxRvbnrC
R4L8uYE5kqVIZk+Ysfiwo7bKdKiHUV/wcNXiCTk/KS15LAJ752Pb6vj6WrAXSuhR
4rzDsKOHJvxffnQxIuR4Yvi1YgfB3ewAMOaAAml70HQkqrj4++jwaEu+qukHHBa0
MaPjJmj6HMcwxQ7H1/9dO8yU/JfrWx7quckw5iViduvopzH9vykvr2gRn/4+vDq8
Joj7FPmpQ6CtVOL0uw4jIA2/rPT0p8MQuxDEbzkzc3W1hzfm59gm32qagMlQ3v5I
rE0oEWWezi/eV7A89pPgK9w4Crd5MA6veRYM7nnYSC8IRvneOt+CJk/5o1Boi0WT
Gjqugcpo+rc37VdNOGYNAejo6mvazK3pVQ9Kowih8HTsGsPIm3OHyXOVpUM55aFV
HerhjkgEpcL1mQFaT+uZ1kzlwLdN880tw+eRna2qqyw5mXjz3OY96c9Chqe8zw7h
7lVLpLRW3LZxmMvOR3F/QalB8VnNGZ3JbaI4jL3yViyp2+gtbq+HXy6PLBoglVxJ
rPQ2+jPo24UgpoFhIrWqRsdJy1OBx3rkGNyU03/6YfxTt3Ed3RE4mj1cy+y/5R11
WvRGLLByVZ6rWLEJKElGLTQJjstkfT9ate2Ouww8C0sxO48r2IlAj2Q3Y9AubVrE
5/Yaj8NqzSEtirMWk4A1LZh/hXdPFIJpJYNMe7FvqZGNGZC9g/TT421eyRQRYlHP
RBR3KrJupTPDxEEkyPfYQULVbH1xfc5fDbNIwQ3Tz8qfFMfZyoqzzkDiMiA2lT86
WvuD2hIum+OAC3cOrPFCciHKxek3oWX+8304BnbL9hjr37/EtaISkm43GALvZy5S
VcRSMI5YjvAWc/Q7ZbTPHK9a/CHtwKKIz5qw4ptUp7YqmnMevBlNUPGydy2P3Eri
2YoP6Sc78dqhJvry/IxYGxYWLi39rMX/b3+5mPsrYnLyRI0VzsAfa9/PyFiVd+4+
F5Or6Y2m8kmFxnIgd/75PAVSh5yfqlnLL7V1hdqJHYO/01V7cE9J/iO8QyUNqE7S
AMZeJ9q27alI8D5EBsBn2lAdcIHKdxf8Swqw10CBzeO2BXxeSWt3kQWZvUWao7kP
fzl/rcWzFySjUViMLVkokK8YWsAI0OWct7q37nQQktDa5rZgoIR491h6IdLHz6lA
NCLDzciWZOkUGgCYohxZKh0m79gzYunjWBq2Gvwp1LsSZlDVI1EzyIhJVMhPjMXC
UmXPVVJLWKWv5zCvgIlhimx9dT4wq5lnRLEaJdE5Ulmktu5szRp8T0veTsL8MDmc
u7MQrG0LdfnRPIVfj31s7QKtozhK62bZ2tyhYv2Xpg+ldYgfiCUqkGyLS6TnuzHm
Td7+BlL6uPMYqdllQwP6gZR53iggalvlwB5AeYTY7kDGC3ecdJHK8zmsRm4srmfk
tT63H7IBtZZoXnTEz6wqcf4SfQozOnRXXPN8pChmTASs8ACDgNmMXay/S0XMgTcp
XAp8pnfZIBZ6pL95Ph80JKcooTA3r+GLzGJUTqh6qMQx+VYycTdJTP/sVk/vcy40
CGUhVAO9kN8yCvFBgozVNYVB3rk6cMbTJjlILAq+kid0K5/J//pSU9jOhkirQ/WR
4ja0zgDTToQQFbG/O7ei7BnPxRaK/hm7KK2U+JKJetWhl9XwdDqtSy73wNqUiNnw
mZzlWgTjo7FiDs2rhl6+1HE7GllzvWB5spDt1X8oj5waG4Sw0gvY1jX7cqZn0MvJ
zzwhfnj0nM3eZ1N0Qb1nDvhGWQNhpVRfYr9ULIZzdkXF0hjnewH7+mJ3FKDCysMi
BpH94/+kcL7mhUaN8wyhBkAc1vHlQy0quloXJOnGjyP8P2oF95lUo9WGPXyVWptg
352BBvaoA7SCLv09lzFaACS3Yq3BaAKi8t65m4j9qXgq3OToCAgDk/PwaC0bE18/
NbAdY4YacCvskQnYxS/+q9sM3b/43tf5FEme7g0pxFhaxmuUx8ElRqk2yC02c/sR
AgOpLvM/3K9/d3TI3ruHaXePNcTKt+MpB01r8nKvJb9aKm+dHpv6qlCyiVi6X87g
xnmhVieLAEmPzeSpQdj3ibrZ98Sr9Rg4UF+OyAJGDGsJnkSWdH0RqvZZqj5I3Jmo
TkRq/Ljhn/DobePO3Iw/Jtk00393eRmjIpXX/CHBDFpcsGVD9FmxxOccx7lJZ3+p
Z3wXeIeB8L/k/489Y2daU/fgh89h6+9Hqrpd+fOZa87aQm7F+YmE2e9qXlrHmhvz
b49a7HYDUycHso4FnuvjJjUftH9AOxynLvO1/UZu5ram5VwBuHVweb349OhtkBuK
iigkZukYIveiJvo84OV58vPPeMGteIosOZ1o3YgWpmFEUHR65apsCQ+Dfz1kFdKo
ZCQ0LcBtDD8v6ZJ2fbyOZVRmReadOjru3obAObafeNtIhetxY2RZYYwxIjBRslHb
88mT79cwVy1A9PvoTQ+qazUjOOqPm6zJKNknNPvqaBClizPjlgj46o68akTXBYAa
ThVx3VHlA6UDj2NynQgd/ZRIPMbNRxckMcfbfPV7JY9Nvlbg6pgXQAN+39lmmtNi
0l5FVb1wMfum7k1n7ZKT4gtQMdImhFNkMnY2jJHq48BmUoQrYIl7+vbSNdLDc4om
wY+9X+/saWpLlVb5zwv0r0nVHgG701IGUezUSFAKyt0TKoXaJ1TLWHLoMpsww8c4
CrfAAiGbXIQmLubiTNRRbs890kAr9RGR+b+B81PnYvrDWqsn12qWAAS34s3d7FoQ
TP9LQeTKrfBpSWk5sSmDHJuOrD2TuQaWIek/0KR3CBceKNxE45AOf8fQyGyOF9CG
Lyb5I4Ms4/cLEfJcWP9IspTUtPJXdRjPjNxFfMQAZMv+X+inn746J2Yx2P6Eljno
Py3X0Zm8IfjUe4fhCytW75nuqFBB2BuigbvAcGd6UMIZii/nCzYInxWTnl5A3oRc
HhedjzSf2mgQRu2w/HFOnkNFzB1hU/3Q+koMHYk+fhCedJfRADgHYTYH54A8sBpQ
yyiyBIUFA21MyLC4UC6lXA8tSeTgnkSFrNw13hKYB8f5uLP0dyXCmt371eDQyUs9
+Vibu/O1hLNEYn5WKSbBkZ/6huxhdYEwFod6ZCIpkxnOvQyXKHgVZyyghNi5moOQ
tvoa6TcYnD3mlg2tyfpAdl8YPTW6WU2+UT4uyH5rfM/Kapsp/wf2zoUpEW4iOrN6
LBh/hcEr5fsAZPzcnR+FGpMd+AaFO7Oz3ZDle+KLQRVc9XyEuMMtOg3ad/6eBX7Z
/9rlsTATcwO/mKu8y/5UOeE3F7BU7Ix9p2w+iFO/QABO92bQwIcjbH0odI1A3vI9
gGFOqNiAbjfarQzjWqlZ/hHMKdJhhU5yLdgb633Iw9A9bn8IBeF/ujirqpSVPQwS
llizqElbfj0dXIIWeN6QfV+o6rx62dcb7QuHQlgT8lqF4FHQfT9utizEvQ5GhWSv
4aPyE8O+cRvhF4ojoDwtXK1rbt/NdkObHJUBpGy5Dm8Q3b94GkkB1EP42d939c36
CjHd/MKYAfr9wIKYE3iHskkHbLRNXP13wf3IvzDHfdrTnY070z/lqncIgmR/VCPw
cRcNR3X7k9qXBMn6tBM+zAEQKVaC6lYy+RdLpi7hnWLe6p2Oa89MTslrpMOhwoE1
5lBcQTc+Ze2LVhM7dDul1XnhAcj8RT83UMcBMV8mD/cUu0aOsODWOS5rb+qe4B5p
JPIbIfzdkG5rYLCtnkp4eUxhEHp/maW+HQGG7mg7L8/Ze6qTM6CilAmM5qUxK/TO
FaFJkBs52f4iifQN3uyyxdlgng5AmUPSphm8/ykTraQX1miIlhIZM6uSnm8M+JNz
8VBU7NOW9o0bSTQOD7/Be9KOHB6mUxCFT7CrgetJUbX6viGlc1ivbCF8p5zy642A
nq2jtRThybeqtnUIstf/W7QDHvCzk8sWR5qYNAPPlV4jehTDnrU2LGSoIW6Zu/3f
k71saFJCINu/vpXdca3sqOy6e19xkb/6NNzILNziY0cjMpsdOV/lUAWy3OrL5hAd
K6BLM3lmciYCOxbIzg0XA/MhbQPfs9NbJvvhSh6GMM+rLjhLEt0s6lItIOYSIUxl
uM5mMdp+0sTtL8eHkq7RpgZg7rH2OiDz2wT3lnCwLgGzdU0Cz53tqNw5p6leu5dr
UFM5J0Sg741ebSG8anJsSvJPsnMtopqiWyeaIJ4hI1qXcZ7fzRpMGD/MMZ3Fncr+
rfAdC6awtWQmbjqGpZRHQCUgQtvXiAK0q4RmGOXPbmvTtVM/bLqwn3yoZdU1CS6J
EG9p/dWNNL1CsH3e2F0a+qChUjcsjpPwvAnHjKKZW8vLyMx0vbZEByce5D+apoE9
yg32/bjCJ/uLp2lGogAz86rJ+dzaUuJfInfx7iOnZ3JZwycq6m8sGs+AWi+vuIaC
dKtQKyXIu9LZdodjFNIbFn/14EdzPqR5os/tDiRKjeowNQngsVebQvhcFSeFT2Ei
lxNrS9jGNQxH6dl4O6yQyby6EGwMIGFAaNgeomocnm9iUw3x2+3FYEPC09oM7NtV
BLm6fKt6M3xF1vp1J6tjEwqOxtVS+S5qmAqbq5218JTK5OSsfMBAUbXeD3GS2X54
wDzmYqz7lJTSdXvMjza4lDnFxY9uInM+8oepDH1c+eGraXunHMaqEnmF7FjP1Q1H
BXLeWIn1piDB7w6WrZ3PDtv9cOyw+jnzzodsiWTYq+1jYZd03BmbWq+/Sn64wzE4
iZeeXL72oHRBgWxQYRP/GUc+8BlgcCPNtNmwhdmFTw+oDdTnMoinHJ0AC6yypLzC
g4wgONpRVtufc+nZrK8zmgaE6XbV3znvj72F/f+sv07Uw94Yp7tkMgsp10bRO3xj
dd9WD13kW206MlrNT0LvY6UzW5/mKEDVH3M52siubDOwLGhGnjhjvVAXu/COJPi3
mIDJHJunuSuFePrLcqBz1ZMwvyEY+9sQ7P6KSwl6Z4Lcp8IJR6nJYfEUNJ2QrbV8
ZRk4G+tcNjJ5Ff1xWwv7n+K3B0f0AH1Cpoe6AtdjbauxU3xfg9XJyNJG1F/MRyXX
Pb2lKJKLkCiKay5iyorpy/Q8DlVcGZCCQZqs4+Uom8I5WYEjfP5/oqky/IfXFgtY
J2sWrihZwbrj3fkUzXkluns4xdXhh2H2LmboPqK7YBx+sYrHz6N8Yxq79YoAbPMS
IN1pHJ7XQurj3IVulrO1+goLJ5IoqshLsKlPO/yLzisgk0wcZKxGKgaOAbqFnErY
Uc+mhudyBUzmHlWOFqgumVPWyd6NnG+6+2NYIAtjFG/nm+z6JoulwA0KaTOK+nRv
vIuiBLvOxlThTVGQA85ZibdsQXMILRggXlYJMJOb4DLBFBHRsGkTAWHRTPm2zFL+
ncUYhQ4mrS8rS5cIBgJZ+vmOFfYSUrqLPTjg2jEFvebUr6DCycffvr8hb+NY3iR7
yQT2H/lLMBirahX/58S0khVeddmXMztVcQ3z9HDaom6iUNzNCE/j4FVaC0XOTV1G
gFHa0RA6R0WcuVcZtNVdcnioOngNKSU3PMiYbmLJ0dtdZkTi8cZ4SoL+NfLKLMnS
t7539cfqZPCLpW3LsNq0Y5fKGybmDfjjG+lbJmQS/5i/YiNcneTk2SbxNtOQT2BC
3cYNUbDHSWFllOGMhALIf8h5fZMiHzdI/Jr8w+K9xIX0ij0u63C8D+rtjv82u/Lp
eyfINNZv3GSp7FMQjDhYLbdScvOJbu7fxpn4Mab8m9SZ1snnALs7Fw8z5sctnswV
4vwGfFcv/njIBE460Vx6WCBLZyeU8Tihdpgo8j+K1q0Vog0MPRZACdPHF1/D6605
9Z5eTH9RdklccW2eBHM0eNHZsSFOy5oN40U0/2B8EHl2PagDsNtmNX9AaAz7MYNN
Q5v3Y81fLhVhCy/CVKXsaSprhsQUDA3s9DnQ86NEq1JXpkJrGOyf7LbZRThtNRCz
dmUwMo57KmvrGQVJ5rNl2i3rR79TFkbkuc8u8WMxfFv/hyDPcDjPSallq4hrQuWc
xk+Ojf9JUNx2xrzgYn4Mx8pToRghwxiYo9u8JdKedr0wLKLBr+nCe+zLQ+196w36
9cl16E585rGBosqvLGedY+VhTq87kEY9lj8HNJjUcYdlYhobzge7FoCjrJ9u52ed
8RqhT0efFIlwSsmzBv7Kz7S6TzVOlca3Emxk1Y4QVtHY3YTqdVB6P0lDmKxRamxI
57qc6VDoXPbOatk3fq2923/4+Q2nVwHwz0J+rItTWYxfTBptOBl60jbYVR/CrXuD
bPFg7CYQv6k+k1xqoBe+31kytjHT8SWhc7IH9TkMzYwiyJEoTnaf58bSmNXSAOzO
BkliqQUqsexvBlZOcLlscPaaclLMWURxD+YDxuueKn2sS556TCw9nU5xWHYF/unE
mWJ57/6FydO4/ZrQ/PigqhhxreD5IMcXQ7v56ixlZU/23OJc6pH9Mby5KPvFHfoD
VTOD25+icLwfXfyvdsV8OOSl0tDM00vm/q8pYNvHq5fFQ0jLs6O+DXKNK8Rf9+zW
vCYcb555M1+rTGj9QYZfpXIUyUyyHcIvpzakm28x7L5SsDKC8YvfdtVix/I4NMXY
qSQoO3+YtVAKAnPqbhyMRVP/gOE0SNqrb1lqb69X/jyjonwlv73s2oRlaOtrv4yX
40EWwGwlALyEyHQXQYJpB7lXcl6mOASnKBp7+pX3H8bFq2rLrlj7bZlctIDWi4vR
1vYq3h6FzAdU4JGjzWBk1l3SYwpaLvLzQQDGWXKkNCJ7iUP1xkhIvIYAowTT66Zj
vvWurC2yoTp4hT28/RueMPtSzvFiJ6rpKzkM5YdxcKwCkvahFwU83nb4mThNDP+X
AuP10QcaAxbUFS5oiGfXUNlpjLeuPyaD9EXnJ/p1siVmN8R0DBnfrh57PjBBxgum
R4C6pF3BlIoXtUnnQINgYeVjjjoj4bWSTFkzxREGRun7Gr6ZVnG5l9nDs17xajfe
crmU+wQwPVzAiLC5NqRUdWlB/4oyjbebOFI2p+HfbEiOIsFYfHQLTFNDB+ZwSSDk
NH8ZQswctn2SQHOyYlL2s87L7r75zlovj3jzTAWRbRl0/RognxU0bJ1oBt8+p8Ku
KCLbg6YTwUfZ2Ol2IZIpJtboraUUh5+kHL7CvT3K48qLCyIttdXQOTNaZ0AwhgW/
LYPvBVhYiyJRqV7w3ejqdDUAEYYy/NFQAfFDwjumXlq3kkDvTCix9x1O9YddZ3az
kdQnEgwvnv/IuQcaDYLpqflD4Wjk7YykAHHlf3tAPEl0+RK7LRgbhCRl4/ygmH+o
Ovx1s4zHBXae6F82x+DUErA0dV00zngIR1nm+Vefc2fdikV/7jeQIImBodQjFMiE
6OOuVJZfaTPwwjJg8ob8r6RkoEdTY/NkJVH/iE+ewO5Z1vSRSkhJSD4eslE64a9p
GCAYVWYpbNEbb+7FynGaOh6lUh6W0XQ8bKywu79pQyj4lUAlxK6n3LKmr7+x66Fj
t9s3CqUG23FLEGNPvlQeClfAlMSFczyTtkDYU5f0o1KVfClXtzotbw2VOzqtiSGO
Sq1O+m0vDWGyZ/qxFkR3QxZmN4sgc9NVTKgWhq3rlvooO0Y3XHEBa7SbwKbPMXvf
XwiMcWg+YshYOQnW90GYLy9luKkIcNteEIYEiPuA9op2XnbUY5f0VrukMzNRL7p0
2cY2vEXP9ax/irUBDkxB3WN8RnW/+wci8cPxQDA75IXCKWuH2S/1QhZwfuq/Gm7l
1mV7VrIdN95QPw9rdFeTgqLNy4Jw7/o0xRiZjnIZ30NH/Af92tHXP/cI2LGwrCpq
M8gVWU615+WDFmIWMKlFo3Mcp9Znf5vnxsLHNnpwGG0Tj7mSjdLk2bLBWD6SQ2JI
PojoZyS8TTgUYY/Kp4/o61O98d4nEN0smNUTa4v1DDoInF1/5huMH5STH+B29axr
Ff5OzmLzRDmaAkfhTbOpo9OYdZ5Ks44+A5mN/OdbMwG30HTXAwaELnmbhbg2ArqJ
+RtTyOJTeeYfaL5yPE6K9JTFlvGBadvZdPhTDprGgYUKGIi+/rGIhpNpQ8d3IFSo
J5M8oH3/FXcfS0GopyntU7h1qdC8xFAEhz+x81rDyOaGl4GGJza0Vgmaqbg9bl+8
BSwyUMU1Ogx8+FTVZxU31vpt0wsymC/U8XJ4+WWdmYaOn0gw4mco4RnbV37Yy+i1
CUUTI1yd0NzOgcgPQORS6VrRNy5uJU7L/O1ijnK+YIu1VKGDsbDUefE/B8Vt9lrW
3qyHb7HMX81hsKrcBDAafl4Tp9AwSYDwVvd5poHMHuJyWI5tmPB+3ELCRNToJn9o
TXoRCL6gfeZ+i546mNby9S6DM9MtLprxcdJl/qxPBrsrGxjH7Vl46U0ma+ubpl6t
lHbGIMv+vdNA2gDXEufgPMtnrMCGz7j3VAUgaOB4TraVmHDEk/KEXqygM0tPTb7m
/UWAPiLVIKeDCeOXaQB7MnOXg2nNh7ydOEZa8gIrJ8rcdeuEzdk4I9FrTxSAQkws
mPZ9LQ+5BPpDefzMbGUtP6DCKP+uT0hgk9dBKrgfW2F7X01PPjwgM7hH5UAf1HPl
sGbXMJLmEhFhUojayBTQFBfIyxaWgygbZDL4uA9DbXxO3SuWbHEf1j6AVBPRN9JR
UD3FNWapEZzRjhHx/hd2D/PMjNsUgSrmCR2952DWYjYYDN3bwiFyEeONgDELir4m
agE7hkVcaKSml7TbYTQotI6IBX8Luo2Hjg0kqthEQkK2+xGnHcedj2ZpLVD7VUlW
XCtEczaqhu4NGfKZNvf6zeJRYEkfVboSlf9/EX8Hn32LfMBEINNSAmP9A1vI25Pw
LFuKZUEAj0Fb+tmlXZCeu5spviLdFREkBwWusk+AGzmx4cMkI58YAUdzMV+P9Gzg
dYePjq9kmVWy/bl6gdzREEC4ZepG1WGut+KM3jEOULc0+jib4laHHdOcKTSVKhbd
ujv8G+3dkI1Dkj+L1JTrK1AR/R8E4Tii1xMkE+axT/5xpcLGUhwTsD1D7EufxXZG
Tt8jO7a+V1ui1+pXcadzb9aJB/SL3wRQf+9AgBq5+5WvhxlLuodwFLuAQp6bCN+y
XVlp9CU3kMv/+WVaIfmxcGdwSgure0dTibfqzToRt+PF4Od+Bfpjh4VHp/wsuHWD
4vyU7hiSwul5sIPSdZRM5sNBAi8HVn6y2ClNgkjSigILSiik/KbRlzPmxt0bwp/e
Mhn/a8p7kL6hTgdVUOHS8FGbb5aN4pQZxD5Mm9Wb79vQFG/XSC96xfJLQJth6lDJ
oSiZSKa8fr2vVe0poLZkzRXZWOV1x9RZJigfOq2hpDgSwZzeUFTAefZzNAIyhL18
J7KmMZtFyHilYiC4I1SWEe+tsfnsOE5Z0puO+70rhzn382t8uu0HznUPkslMhcVl
A+kCJ1P02iKR+noom5UEjjvsUiX2ZLVcmHeYsT1LeglOnXqaLUbBnh1ej5qUsZa9
mCiCfbcMiOaULAaOJ5V7dfeHWf7SsjDhdfM/t2/TaFUYYyhqACiygWT0njkV+Z66
dIUmHqIKbWTPIssxo/ivE4LHq38nFhmtEAoLCE/SmfOLmCWFBB/F6l1QVkwH0raq
gEmuYAexRnLssZ0WLCWXpfsZAgjvuHZaR7X1yGKGrwBq8a6C7IwKmCZOV0R2evxp
RigyQKMX4owc7j7j5wQZ11/kVQKEEN7EhwH/uIG1FAaXABA1Fl7nZ1zRDwVn39/M
r9fsUUND1t4WncT3Aam3qDeRK4KinsmHZGNM/bNcMN6ICnXtn5iX7cWTDtH5OvRW
bnrZgYaMVialpAmBGqhODTcp/twTsEHnPEWi2xRaQZup7Dhoeza4V/SSCS4l3aKI
38PNUFXS8ONpdrRePkJOAoRmKTY0bD9928Kvfiamdu7O9iQoRQ2/no4un9WA5/hU
JFErD79pVLTR8IHfpm5JBpGFXV+xcTOA2IrHtMtCn2Uw6SwXrKfOj99sKNnCztOT
D4SoiF6ddYCBIv7CPUQkJitQG4fOmkrpSCUPv/664P/5KSM4Ip+UkSyk6U+6KsiA
03yrMYifcgBA+2SVowoJtpQRw+kmJF5RHQW6VIb6cgrGxvlgSJqwbj5CVsJ+BSGu
EXh9Ta9pv5ny9K4uKrRM++zN9CkNgCLwRBcTutujHwtb6omK8jYr4TnOR594xHSx
lsYQg91P7UBwX06NkGxSK8ejj0innqj7yRI25rtx+yG0JudeAmRFQXgRiw1OEdaR
NMjyu8ZF7DHh/M3cxBPZ6gJYo49us+RrpkkWeSQ+M7F0zPbDaJF9AiA84wq58laB
YguUfNZTT8GyCJkm2UXEJTnSiEhrEF++GZLbnIB96REZYq3Xp22LMJM/9aMq7bXe
oFMXf2SoiTjeQ5hSVf0VtdDqq8oED30bYVdutBg3OFwUjTTixMOrt29CVXWkKjMs
OXE7W5o6LXjl6PKtVPHSCyZkR2VkqPQ51iZj5IGFJS83pp0Z00fE2kOVcvfZoaO6
5mLPsWDWp14ARFAlhjRZ3FZm8XicVCEdC0S/8/fvl+3fZso7Xf6aqqWdDDV1SoXG
pGFlgbbUxRXLjOxn+NY7VQpU1LiL0+bqmOErKXK+0qHvMBR9UNU1L//CAI2Q/aPt
gSpriy7YcDtR3grR3O/o0KM/i8cCafxWm4A6Ux6/jOjg12sMCpdEknJqftWb64rk
g4f2JqbPvmy0d2jOeFHtsuFjEgEQPwSwqkMKFAMXSBzmCj+TMWMcm24iXSS0IUSl
RatBwjn+DyLT8dSDzT4aAzaU3urNDWm2bBqWhxFjFwCS024/0WCgazAAUh/o+Ofj
kH/X2LKpgzjVAzlhAkWFmd9Z77bA9VzRNBGbqQ5vGphM20lQm4of3m2nWsOU7hfe
dv8I0JWCbQRN2DTUMN583Skm1Fbt+L1zXByWpmQM2ZmlRzScMwt1e0eiKNjJOmfN
Fn7h6KhyTi5CLSskuRi7BkQNowBZ13Ud4H+o3zhK8Un+GMq53++GyhMcggoVah41
nSzR4eblkQv0mvtmHK8HWq1ByncSxNKS/xV58KhU1wndMAX3m4tkOur92oVZlj1f
zrwho8dKznG2BX0BHzORr0eqYTE41X6fyqMnVgjFBUwqhiQfcmjU+NUbYtQRguuy
YdI2ZkCO6d8BjYjw7MZ5r2103Q8QsuavtzFMKANDuEPbdJWgD5oJzxFkvHoGY95n
ecwZjAYG987zL9RIdSu397myJ/oKF8jigGXsPdl6Pa00nyR0RZckmayaMsrWIB+7
sbYpi/9u4OXXjce1ZxfGurQ0ffMtIK6ySP1tP9rkQjGIEnIQWxvVwzd/TgpZymaO
VBn4PuGjrCMMOlly/6gk/cke0v5iMNakk7qgwCognpyKV3hUvzyLRrSIX5q9HeNM
7Oybhx2po1tCDMKNoUKR3C3AIjNp2XItxv6AvVRiMx9DfdAOM1TaFb7jCRZJRVjl
R3TIx3gAbfkOLOXsrak392QCGNMM9S5YHe7qalySK6WntJ09/khtTxR4V4BndP4o
z0suQMN7B5TxrtFggPeO1utPwIPG9rljOfkwgEnJzsr9ASbf46OqgNXu5jydTMRi
YU9kYUqDBpCUAG5pkWbwU3bC0RxGyuDQDJyU1uU99aIIkDMymbWSbqCOKvaAN/Ym
sMPMPeOyAhOPuO+D+D3yHqWWuy43U4YVy6iOJ/j2oZOwdLpcuyE+ER8734DnXcR2
BUu2Hx3Sh1Qxttp1gtHr4besYbaGMTz6QvUTaFYX0vRAJJ+tJcz6n+9e1wm6VreI
n8NqZSPC5aDZu8PqIA9FfmkPdQEdo9ow3A3NNS8OLFX8j2PYK9Kss72DpUGr/GJv
l8gp6r9addHsg7YgETU8oy6iAlY4QDdvfEmA4M0829YMLt5EKV2cs6v1D1JNV53s
Y6hnjkt3haSD41S+QFVsSBqxF0jL7AiOSLiQUOYhkDJi6MLjIlh7NEUcwh8DVUfh
rMsnrRhg0BRNd/ZkkS4+9jr3Jux35HBO8UiVWjvYT/Rb+6azQtVeN2AKg+qok6a2
Q7sPSOL9tZ5A6Rl4osVoqSJ2xUfQvhISICgdnVL2mRblKZtS3Ud8GXsHKgMZO8jS
ZNDTrsBUA8Et027rkyFdLB6dSghbarHzPKEGWN1vZRddnmL7IZYNOm2FclED/EZr
yfudufb7BQSaiK680s02gAbL9XgdTilq6tDwmVCC6EXM58SOVYEr+KlFOXRiauAl
WHDdIt2GxoWRP+ydlr2fpqIqwvo+7BFS7qd/kSlo/CKBmu6Dziel/DUk/Tvb8GoA
YGtyW+lzgYDiR2SX4bV6TYtGy22v8vV1yh1zKnCgK/bMM72xBrkPruDXyxPvc31D
8UZtpnfvoteJcReWza6QOqRVCVKvGx9NO2D70Oxzqs2zgwWd1tmrB4Jf0ueLUWIc
EvxtRLYD4cRhylFXP6YxvOC0i/2z6GrwP3cLaOi2+QBhqdDrJIeR9TGRbewAd6z8
BQIPDaQExQyNwh49MXbKI0BKOKMZHwcdD74iekDuD0ah+ENz2pD9xSP3keV+BRWm
rq/dsXqgiuGTtO4IoyJbQRLRObY768g0q/tA4KDq2wxn4UBXPDdmEVuC00KAxoyU
EyNKcoZ6EuXnWJO2mlZ0OMYj9Vnfvlsfkm6e82olBzD/PZQI4r0aWuQu5+sSZKsB
hfiQxBHfgHKFvHThRpL4CqB9NtAsMofZo5lG1OeAW71SlfMIgEyATYg1Y+w9tgWD
4i3e4ea4JyPyBlBZOT1ilXw9hqddFbOkeJALuT8cab98bjiWPtP+GSiyCu96r8ev
S/aCnCGOblptRpMcLujbYWTohFCWF909n2qCbBG5Bv86GNCOaWd0re7u6Xz08uoH
m15+PtpYeqWuw9XtIoHZRKJq2nEYdJOPf1Cut77EoexaXnRgc6DK7vGTZfQ555Yp
3kdLuOdQIUuMuWic2aGndhZbpNuZgnlPBNeMQcFsxKMwoyTZLXVnRebHmsgRBb8A
7JlFsX7q7aCI0dtvCrfLG4QIjeo/voqFbplSsxFpxilzPzJOqxiQhhIvqUPCGsq9
NQ2vq4Ml4RWRvadTyMFZV5Txa0mgF7ooeEIBC494AggY4X5MAW7XjLW2lOjfyEG/
1WzAHGXon7DgoqRVVwN+CgWvhfNLfs1qko/SxgI1hSF4ftDAXfFw87tMyHOBNKUC
cLuSX5MRYYWIl/sJ0bgJm61uASovXUyJt/UzaU8tca8QEMUBqz6qp9hs4XOFAl8u
hKWzUGsvf1FzcqScHWKLCLBYlhgrmPwy2GEyjXjPzTakAC12NTSiHxga0EWa/A+y
VwqZcOZHf7TKy5+vj+IAzV5qs2tHoHlNUC4KX558FDQua5/B80Vd9Kkoxr28WPfE
4j1rpZvGtVXrI5P4pPBpdfDfPO4wJc9hESpo6Xo/AHKtGL7NlKUNIuEInA+oS+n8
G2/l+fmUNDuMOtQ4EpldLENun2MADhUFp5m02jDCHfPCsetp94/HA2kyMIlfuIKl
KOAQBl8f/niQPdYV4jboiJpLKqaY9RtacbOjMWhPM8bkIF38BFk+8nY+LEOZGEKY
hIibOO/o9de8vIa5GRqKKUaf/ZOj5hG50NfGkuYhhObT0EOHX4ZCdXKPGP2I45C/
FoEn7zcl0Uj/63auzNQR+3UOl5LCJISgJ7r9kjJC4ye7hD1haH1Qe2tCkMgJcji5
gpgGlConI7v3PCBK9Oo32o60FUKkGiSQ/0+Goho7lKhlbphTunF0FQkanu3uQmVE
VAIPsTKEJHRRPkmCn3fPQX2ZOC5au76Hf7qt4VQW07Y6JfrunHNOV4bGgMNQ0vBv
T8a1HC19M5ZvuxIKuVwK5ADswnGGS2humAlpsDyLObMSvABa91NX5cGXG+YOemCv
lDcw2XyuFeHHPy3+qJj7Gk447v994eNj6B5E1EIvuKDwuUVkrCjOcaZOiP1P6ppd
NCNPYjDG8zlDE4rDxU5vxMthGsTQley9rddegpjpKm/ZRdfJHozBSp3y3aOV9V6T
OavIBlxnin1TnTuHpeQhA2jw4hk8KcjKFYCkOjExxzlukDYr6hrYFypp+vEXVtAL
E7Moa36bxsWK9dUR0eczocJN79FVoLoNAIQ6vCL6YZvAwB+FefLzyhp8ZTUnfZSe
ya5urIwFn8IlC8y2wHiAFJ1cWgv24RRmiEknJ+nXcrG2s8HA85CSvST/nTge/Aqi
NRktrS22wQ7nQ6jgXEsIkIxxJyeN9zEE3DdY4XN7xIc=
`pragma protect end_protected
