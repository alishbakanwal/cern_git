// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TwOuGbyVYszXX+EGB8oqJ/PRfE/2uqLGWo0miToEkAZ0dKeZSOr3obMH8Y1baVDa
81Vo//jMNvK7LSV3/qKxgQdb7wYpdVowJo79h5dTBtzf4AbgRwly85s9G8q5PjaE
mrQjSzEXb2bJg3rFODydDPrW5a7HqJqWF04xOrIsP2Y=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8352)
1aGhKxNRmiJ/VQU42GmHcigoVQeRO1SyGeYp9WUFO2gj8XqpUWaOnWfxNl3G8lfS
j/e4Yumci11HUj7az7kykKguan07XLvHV3BGSJUujTLJMAnem9YIDBl0mivfv0DZ
btijIEXuI4tVzC0F+hPZCcYxhwf3kPB5iBKNDMsexEs7mc2ma4BPCWH9L+K9zyo8
At4t3DXzYIdCCK4JlwThhrwl/4k9L237vRrl+yAg/DL/D7BJf0qaqIo1jMrDpf2o
KMzAhTO3UhA6WPXSvWVzBahiMsmPphC388YJfE82wWcZrwNJNl/n4hw7a8ItzUqn
7eE6Jxj4vV9whj6/jR5OJ3AFQFzSu8dEDWCyeCfhlrVT0ezZlcTsHbASr3MWhiOz
+67Z6oNqgoyj/qLRvTxVJFsNBRrAdN/IpR8VQRIRA0oANrglqgIianitWTPlhB2p
PAk29ctdVTSVsQ0tsHHggcMgi2wVT5UDi9K4WG7+Vis6iBPVzO96L3+dtukIQAsW
kfPQuGdOGwMfhpAWispt2UXUIA83nzRxUVCifNn0tm0TlfHieVEhZoMeyhfh+T48
XDbkPmuqEsvapolBKPKhJN7hvd1kYjzH4UPKtCsh9/6n2mH03mXtln0k0ADVce6D
qh66nDzfNjSq+A4NXGYdXLd2y2bype2ndWfXxz7/hDT53hyt155DTWu5VbnOiVrf
SzEk+eo8xIYckHQUupw7eTWl1ykIJ1Dxyfkuj2LQ/zJufJf2/robaLidKPSrZ6hy
+U/tdIbeQoU9OmCE2/UAxjS7Z+Hj8EJlJKURgMoEtgZQ569trVBbTLczuTsEtJGz
TKWJ8jxGp+MYdpLpQmuv+6bUgygIcP3w4zyMMsm2kP/Ia/Q9qhWU9X9BVxXKXa1s
ZjxDSunknRkzkjjgrXE76RvB1Gz7ZLsT0XSLBg1Uk/O0fEfvRIbvdRgzd6VbdNDx
ilZEXQG0w/ZzrCkA/4tV0JquOKSOrYbwEQ8JYIAzvx8xHweu/0SJsdVfx35GsqG7
51Q5xNXfn4i21Pb7hfQOjxm0Wp/UXrzGoLwJ0e3NXTEcgIjl5WMwNMdbdJIT0XwB
URPZR2cpqrmZN/IWYHqTpILFAcFmPOOp5uOfPQFzrBUuFFePnOk3RZIpFaiSW19h
F9hFdyMo1wOSzcMTyzgnS8lbrH8CIurxwU5L8EJajwTCRGwemLxKvIuLnmEdQYmO
vy5oKUrANgpwNt5/m2y+VV8XXOWk97vcenZxo8+LilfM6YJ0HoAI9iyUvTfOdc09
xRfdBzwT3XLxZVEyDLI8mizZM6GOJIVWfuDOQ9JgDfBamjmb/S9EPzqlAuAyrH9x
oaKAHIkpUJuohrfhcJukUA8a+9RFb+PXVED1a+ZRJ10ZhlGFiMHxrW64PgAUMluh
oVyLqje48s0wJVvk/QiGisxdpSXPecZj3boAnHuHtvie7IPNI7dWuwXv1844pzqf
Z1YyrO8qL7+D7Vm3Xk+nOBlVAd52Bdmi+JXBxZs1RC47D8s8R58WdeQcLPDTQiqh
UTDBrNEfvXFE4U362DYByEBIflGXHsklipxFiaPVFiMW6GCNRVCPj906m4T0F6WF
cPfxIR41hBzyaS7Y8ZN7QQxLMn0dlB72pYeUsWeo1M7BSUZPVBm7LwOOA22ycI9S
XJX7VaedUE1Cg6J/1qnAZCs0B3uLnVRjQkemULniH7AMTo8xuVQAD0L4IsVIOoG3
8H+EF4EO1gaFTCz7cYIEBsLvaoh+KKzU5LaPWdLiwmn7VO/lBAcedvArN+ylW9k7
R/2S34Z8wZIRQ3Xz7TKcZfVm2JZrHTsPdZrurhmNjvNih+zk9QkpUiQf/Qph0PHn
IXFPlqTEeBjpP4j/m3DeiwlYA1QiRGMnFstdbA8xXKPuwLpGlH3QNs7rQadrvA8+
UYgP3yYmxVtoZxF9f5sIXV4sSmcjlbByPDXkP3b9U+GNcKWCpirRNiM/iguMJfrW
AHLEYikPq7W20Qbpf4vYEx4dFrD5ROrrpSt01s3119aOZMfJDl6rElFY7BJycEtx
tnjymsdsFkH7SwcVfUMzdurvKBV6XkM79NTc0pDe/QTQnty04XHgwX+o66bOy+Ec
Fll+1EDcvkPlDPrD5DeuKKqcvI9pj7JLFz85C331kQ9sKIuO4z3WU8OYRIP6tLFr
EcNdFOKoPbNkr/3TscTK4+RiW8laaRWZY2I57E72LnQnRCo8iygRWHH9NFgbAkF4
Pr9HzXxiwNAF1S8fSJ5qwI1mLdYWatP+8XiCYcAviqREO19ZmnEXW06BP3jWO58Z
EGeVLJk5P+xAOCAgaifoX9mFwL2ozh/KnBEEwaTLan9x0GJ3l9PJSy408WnbeZzM
iduBsZaCFlWHWw98lAQh5L9DqU+WfC+ewSKvtUkyjPvduBC5pnyf4HasXwImtpT5
YoT72VRBCScD8ryZUa8ZOyHP+fTvcx5DdzeZMgL2/qha3daGCFAo62vR6RntsJ2L
34kFeV6bppUJZ2hAV8DdXGUp/KXq3oARs5l9vGuOLx5OYu2RYaKwpPFrtfFHi+Nt
ZK+nR0m8XTqQpndYl/YedlBJVJuMX4sFpTaw5dg0aDrvJN8FGCzlaLnb4Ncf92+9
Tfh+CLe+h2MKU7TdjQd5oFqtHWhdTOCOM6xhYBl6FVFg0HDuScqSsW+MmIDdk/Ws
DPGDowZi72EwKsU/evIMVuU4ZHBmUKuBLjzWKsIli4XrLh9pCc/GpKnoLw2CsYpJ
XtEa/TQoZhxEF74wtNBIMXv6w2xzi84Zz3v0EM//SHSRF61RvPpNNTxj5TtPOPif
Sbn4EekM2uJgDPRnqQn3lPndUWdhRAVhHEN7eZcr/SJY6eJR13+VMlh80AqG5jdt
F5iGcSNLOhOtAZ/Kxh3iOnKkJENiB6rECb6R9gwkpfedPuo/qfbaSB1Zpjf6noqb
4Z0BJwkgjL60iE4K9+iD0F1MfA2ew7Hzg18x9NHLNebLSKHzDO9tXqkRM+IRmCeC
RlSRJvj9vFTiHAYh7rIq8ZdwFKNlqbGi0YtsMsaUK1orph1u25RNr6Tud4eq46NM
ma6cOEGRLzwYjerIzJ44NAPLlefQ7J8sUry0PVxA7KUEKfC8rQ90q3RRKz9uitNz
0wwax0UkiYmX+JAsv+JVjbzZUtZzHQsAHmHH8OVLQ1pzSbEAp2ShncjIGAL0h7vq
WKPpvphbrzQxHKF3LcwbMUgXQAlE/vc4khb4KzzvkWDHYIMT07/e7kxlG1b8hS6J
R1pBqpNGt7uzTEWqVQtxBehqeY87bpca6wYNH2b2H//4O8L+Ui05m9yxjp7JgKFG
DGf5gCfznhE4dvTkZs1VFWl+eccN69UjPUmQC+k53T5SjVPgq4vcX6A5CcKKOV9C
p6jqvQbZsStbgCG+nsM1CtGMcFkaB1Vx0lk4jqm7vEENrTEVc4/XTMc2wXScQRQA
76RjgZeoExErAwExNsLnSCTTK+/1kN0bGCLJpyf8/DweYnBoIz2mclrZMMdkFRZl
ED4s+mjc+oKbEcE5tmwbUzDUGKu2/KhjeVAqXIvBDlYGO9+FM5xYSpBTcfGiIUzz
Cj4kdJl9fV7lv7KBApRPOf8KHMkq1Pfe6AeP7MNoIcpe8uJUV5P0zCP9HIpKhHii
fwl6VlN4VnGDktGreSJTkPCxKPp4bJNJjcfYrRoXASML70GorhfCSamkHS3OV106
F1fGEczjESAmrqpKWFjtiq44K4/xT+qPGVfkH/TEgEhy9yV9UGTSekUwdlVMbcfT
jYzVheiJxxZN2aoLx6nVuXYZykKx8Z1fAS74bnmHimpAA1g3ABkmMSlZkJnk0r4T
7NFiI+A8jyuGN4cREsP8OurV7SMcwAA7DgTBnQ5XZPOEvqBkFvh95mUCQaS74VdO
vP9k1h8Ysszx1nYS52dpWOMLtqpurITMOj2QxmysG2LZ5Ud7pG3auudcuI5ZiWf+
LcyPkoUfXO/eq+xvJke5ScB4qpCBT0qP30LpShsvUccfDCMknu+u5k643tRATBI+
OKYZRDweZLfUp/1qLqJXKoKChiKkE5K4ubJ/oh7AhpynI/IIBc0otXdpKglOJaec
2R/SzIx7kE76uqgzEFlAe2vJqqQFu+NfvpbkuFkY0Q+UhSpI30Gr3jsaSPh6Z8iR
R/dLgRGRdjve6F86gYmsPv9/787vYew6aHhhyTXmyIj7+80ui1ydbQ9jw5ZIkTJ6
s2MiLN9JSToCJckKbUR9pqDBU2SceLaIfACccwests5Lr/cgzOhv7/THuMnWSe1D
btQnConqNO+rgBOWXqDrLKXdDnYSGsWB0PEp7ZensqZrOxNFA4N0zB+V9IYxl8PC
v/22y8AzgQA+bB3iSpC3h1CeoL7wtb2y99Tlz8u0GLxUhm8la8fs3ui5wVLILNTZ
0x2z1tRM0gBzVfvrdEwMJoCRA7WrgEFofrMwXKGoB3hbHC3A+f5RFQY9TJkHVgdR
MWtH+llvUPO8hMjyIYqELFEfRTsQabMipnI1G/+4EPWo6aj7O1oG1sGWrS1wFmiH
JBYUm+KTChfYb8oGC5YK57TcIuNT9UWXUGO5+bTTJgZdMHMJa9uNdqPUDae+j6Sr
H98l4x5qvuT+V0sGA9tKC836Hc3Tta2SWVyhW2MI+Y+RpPQapZ5GLJU3KtNjmscg
WxVa1rplTmSbjjsArrJ2EBBmzqA+IVvlm9yrnecR39HqgN3EbEEGdlExJs31T2pi
CCxayDxLLm0JQlYahT+yJf2abfw4htL0ynCGgvTcMVy163gVcs7T6Y2JYLgKyya2
lzlPrm8kZpNdKuyn95pMi8Huv2C2DRcA9s0TlGE6Rv9TCf4LXkE1vJuXc0Bx8q8H
yKT4AwyC8dOYNp8PxytbIdTy+9YiIPpzZXGTFjGra9CwQ8DzFBUjEoYXlbsQ/6Ss
28Hyffrkcm9bf4HWg/oxII4G+KGExKTWq2Iqq+FX218tWEoTVGe+ZgyB/wBiDHKy
47vpt8f4ZS+Gyw24SJJtR0tAy7y2u5k4pY28PKslwtIPsC3/pyNVH0lwqPJicckX
pvqFdciTKYSKjMX/1nfzRQ/u70gkKiF4MqeouQ9B2VdjPa/kBZLntuRgo15XAP6c
TAdtZXNAeH29dS0GymEupUGTWhC00cIyfCQ12ZJkSU7OblAhxCWeEZpM8hxuLEai
4pfEhrtFvh7Ua0/Sesy+U/GU7PD5ZHDyq2LKsEvmyZAxenuyG0fMNA6SpB08WPZK
YD4n4EvTfjxnnwjkSC8DfInI2xRSAFrDEM6kh4kLnwzFZQOrD8JSvQKvinoa+cV5
lctaT/g7XdNL2EQA/sRzF/ocqWSrBLCf8Qy4ZjuKL9iGtYN3fnYQSgqYvCflmcOL
6OYB7CJU0k22dHyvA4YO/WB8chw1QuNHRhK2jYQmGapDcOPvOoQcjsOsvQl8trIN
G4NeYWzEtPqbsZCMeIuKwKfoIumXcT6CkO4i0N6PvMAmNQ6HIVSPd6aLrMg/YZix
LhWL4gooUTTXGd3bxcVfVY7n1v23+UaVFrJi2+/vnX94gkxlOtWDYDlJWl4TqirO
YmDJJdlOKB1I9mTl3uhOtS3ah1eNcOT+B50jW38ofB6r7fglUMhtu2SwkoBoaDdj
/43ouBj75bcVZLLzxuWewNXaHGQJQJYSIywM0zj5qRL5EG+ScrjqdO+iR9JN80Xy
5XCz2Wb7eBBax2W2sIOW+LeyLvR4hrGHMlaNBxQuOmr28+OJmPaGUDlUMNkz/5uS
SaHYaUM4xIAGw0RJq3q1zfOAJTifUNEriE2++1NSkozEspLt4lpOsq5KemJT26cH
6igJ36/thgJKk9ZI3ptPUAfe0vi8xDu18462tfNZVSgYyAIZJKJWfylWhJ7kC/Kc
neazyk2PEElGDv9DHRWTGAvk1NsVMe7u1h3AOhosrsRJHiv0g2pjbUfzO4pIXmWw
c68KQgY0ueaOBurfqRhBtAdr4l3eiZVXoOmQ/+xPf+U+zzZbSFKVDBWzrHiB/UcD
Bk+iLZVhj0DP/5apoV2Z6ro7gokKMh/1SZfhdU5maZ+OBgu5I3Jws1Ign4jcAF2P
f2XtyGgmgWc0nGtlAxObA7EoALAtdhlDq18bpPONYuo0KNeoI8k1tH4fVQy++ep4
6x6n4cDEzFaFbJqCotUKVTz9QS+dPb/TUQb2vbzVc0AfxuQ4/pfar3Kh+IK6kPD/
aPKWqXZyxjH3QuVJJ0KW0GuNCyu+WVa/dUay3xJTQX7UkkdUjvAj+gbo0iERoGCf
E/T3hjiTukgFeqXUXxs1MZwGE25g0tDjCcT9l7dvQOq4+m2zp4WVan+ULVB5/CzJ
TVSLrb4Ud39+r5/Ald2C1/Rr4F3Nv2MT5fW2ffahYgqLVjecQBKQEvn/nekxC8ez
qxDIf7eS0+lcMseymBGtae/zEXKRPragB9x/fOTfxopbtLx5aXDkDEwVR7JxAUrt
3CoKICCVY9c40yEJZEBzwWkiL9b4uQKT3S/Ej1Rh9BdMhpUdfQU4Cm/MJvzWxLVr
cmlBg6UW5K/nJtNSM5nYsr+C7xwW7NlDMwU0ovEpZNva9gSgrn6Mqx8J2wRYSdgx
/p+ij+T3vttKW4FzsF1Q4fI1/BH17Nu2Bd9WyT80e4Hb+EvcrpFzMfqjnJsZ34uy
A+OQOmpSKXtsxmlsqGzCWIJhFqrU/arwikj/26YRccydqdWh7d47MOJpTnztlzQX
wV8XHjvyltsf8PNRsy/zb7c11XJRCGq+vYTCoRzbRlMP7oAglKQYBzz/Yzs8GWLY
T0OEdLq3chSm6+up/hW5iWQS+q3y2876TRbKJ/eLsDNOVD6FsZCB4xdJWj7Fl1Te
ME8IHFlQLoPehcgxNpGHkS/sJLx97tXKCKbPqNx5XAWBak0pVj/RrXgNfsFTRxEQ
vvQHQS2K9t2SWcoMXHF/tGUywOAv32wL+GlQNQhN5Ab5z8XtfAP61GygblCyNYRC
z19lINlR8qnZ2MCVJON5h6wjyy5q8KWkSeiNmxREhY4NULGzbjb4vH0JjduMmbcs
3RG+2CFAqAz94rSYYOkNj6p9+O3/QOnGQmqSs1inHHg5Lc0K5+k0qiQrB7EcvTX+
8MWw/sbWuNYrhD9LFEfLb2IJ7C42DNEbyu9wKOsCJIR4MWMLg0o0IhQtcjOTV9pz
fkOB2nJf7bZjD/F1MjH1CwqX5ByvBrIk78NBzAA+L7boQKhlH7OajbBH9RyHuY8R
bZewAUFjlAnuNwsfYSDdk9JAKjB3BddXVCxI84omb08+Lq0MueVIEVifo4PXC8Sm
QRxO3h6MkkFynsEOWnaoGVONxRM5AYeqiSiC6fRBc1gO9Gfr7u8dZWawm90GqUZ5
sY5Ty430EWRQ9XNpUafvfzcrsaOKLhkbJ9Qt3zlfy6QXsZZkhg4WQqXp8XY/JbaA
lTBjH8P0n/AsBTpS3TL3fvxbX6JR2QnSMpjqX+jhi5hyvI4vhhIheKJ96dpIZL37
7WyUc8nxuimw5RvM94ZqlandcXVvMOw29EP0oCagoMaD5FaY1wEvL2Ctewh3S7YG
cQw0UNSncMFcGWPe+6Zn00YvtW3NYhArXQeEoYkiC81H8al24D55EJvZ4ogXZjtv
Nxt8epoQs5sKf2hGrLOFpGhyHMVwjBQOsCRIoGb59TvrPa34OWR5OPhd0MMCy1XV
9QCg1/xOKw4Q6RKVa866Qxk/EBY59KA+gGWPj0db/d7NvNsVX1TryTB0PqCbC8dt
2h0wFIuynYXiEJYqnb5YHWnGBmiaD1ZYmz9Zln+uzcsKq4Si+yM17avBkHfYB5rR
isjC0sJ0x7qHdH5wQeDckEkNvaV6anUnf7nKoyeAGq2f5hp765Uuhr/rZJmeEk4B
3KsxJZIW93N5ieTHjSs/B0kfSR1NOufKqPlAUT44DDXnqP4lqYr7zJ2ORE114vxq
4RwaLcv6Ig2LJKodHovyvvwGb9KoPpAxMd03006llFA0hhjUdQKZpJX4eVptAbc/
2WgcJdcqKJ0GtIkOVuDXlZxykJbyYhsWzJCqsop9JG7JtmQv68KUX6KlG56jGRD1
62Wq4/HPxz7wRY5INKMk/YzHAUYPG5C50NUSe/ibk7en0Q+NS7uHohb9HmVcWDTZ
Y5yj6DT2bom3XYIKsBcXg0rrl5EC3Jm8p195wra5ZDAlStEx48liImLa8p5ng9z2
mMwkDBWN865Y4DyLB4OILojiD9BW6LHBHbFqlEUOz/d56Lf752a8r8mkIZEQU5eJ
cYO/NAa149+4YiAhhwHd5VqTvyYxmO3qErI4n+fL/YlSH68PGhl67gzYWJKmCVss
6ISAKBaJ9pR8phARepXRDOHBfIPMVs3FjX7MhzaPRmyLvExIWxOCJ8qlfsm3dVhR
5sklgRtFIeB3YvXoVg5TdgiYNZRRr1EwWacqVTUY049KsCEtwv47bUdx/fQKLAxw
IEBA2o6N/6GPPLEC4REZfPLRroSDql3Fzl0JSesT+A18cNcVYrSOmtyjdJL35yPi
9Qy0/l0b+O1TxhQe5pOQLO0OgOA/bJ6PtAqCZbzY/WdyE8KYETHTzMtfVxHqj9Zi
nCWIJkw3QKM0vMKD3iFPtN6L7ZIn1JtZF/o519QAaL6X5IwieXDdgo0TSNW3ig1Y
8BUr0VaicIxEtojmGjM043bV5CGae1KAW+53uFDp+Od9X//5GHVmhxlMt8vNWC1k
KwVk2qT5DcBN9PCSJv3hrrQ0J8HKhrvdiWcBJ72LGL2CRB6sSo7/+Rtr0YmHvHx1
OPiGVJzIqEKt3Cyw/3Sq3lK2O2QUOD/xLsOcb3kZyXs0YgVohXbSuc3kgKGp/MtI
0FKOqCR19zrIOE1Byn5v0uSQkEnVPA2EPT7+aoYvw1bC612zIaQZi5uuYu0RigE3
7I0ud7B0O0L1YQeeOaZ0/eKAcjdTTYNKpnQIQLOQ3xEugMtrbTEhmmIMXhx8iTR2
eCiYfo804hK5oz+C2KJRG13t1eJlX4Ga/Y+uFy7OXC4e8CYaa7IldIGcdWYfot+j
3KbJscCPMgMP3lz9QmEdsRU/DHHwVbeLp4zUbCrk0SwmIkDfcnyjdoERm0tahXES
1batpyU4AWTptXz735utt9BmWfuz28IRMfqdWb9qWRxA41RPX4lk+7bt0GgbVbTg
bhYD6gi0pXf1A+qoo1xV3adUqSYCPfgMOOh4h20MyECCAaAspqYn3b4pI7sOzNX5
Eyqj2Ath0LKd28uT2j/LygoV0+QqQCLh5h852PpEzESXtpu+wMRsB/yaIY2OQVfR
ddTCwl8atB47pbj/+iVVSV9Nza+tGlDxG2iJGN++Df03d7l2PBLg5iKphzmUzd7c
GelK1asnXJeJgTiJ4EGg/H82iAtWPQz38fjxb5ARFvD41Yeus7PNd5kzXNV9Si66
Hjq822yqlWTd6LhAv2sboL7QXlydQPcpARcx+s/gHdPwp3eYDoHKTiN4wWk+qz8+
CA+z+UozJtHmmjVrgVcatkHVuEEHjFerwbITHWB4hOzzH9h9nI2aqpG84XFqVMcD
D1sIqqkrDshUOrSXJIO+WyE7R1WORTq1tbb2c2CFWlcv0GiQiPjj4TE1Hdx5Xzsc
A8ZQv8ktQtEvfIB2WqNIbUnW1S2UF81btRfNNjy+XwPOSyOXpGZQECvZ2vHpJAlj
J0FKiywF3yaR0pLZp1weBVp533kIuxPJyZMHKNoggO38lLDKHoBnjrrUijSCuFrb
QTe0aGqWTjmlQsUvMbB+TxlNVfAXCPviRvX1bzpDfCcg+buDbpWw4JR+4cWX8Tqe
RmpiKx4Vq4H3h0M0SFbjsVLPw4nWThO0Q14K4RwdHNZ+xL71Lv3/zMt7FNVe3yuq
kSvFJAzh00JtAdqA4mRck+/rLZJVlP8pQVrpwyDtM3TDNXEosZQOWLt6itG4HX/j
bGd0c9TIBYrHAMg/Nf6NmFhewdNhS/wQY4dh/p8GGRKk6669OHnzgUH52Dl8wSkS
1A3X9R0Rb7PoMxH92fMCBWiTclLYBrNM94oEOA9m8FYmzHGQf0P/ZVT8XFNAp3y1
ycqFdBSPd5KijIBVRrOhOtJ6l8LWsMxAzH8wtz9SPDLATr7OTb7h04Nw6xjcE5yn
/K09yXMy78KnlIqPzpfyM9HtuLzixTKYuoC2GrebSkFLgPkk/2vfy9iFByeyeutG
oIKUGIHfu9zHa00r9iZHW1BeDyH62sxz6riaI4DG0qAa9QY8Hv/k07L5qyGxMAOE
AWShRsxOMDtaQ1Bq/d7JbKBnuUet9JnRfvFPESJd9DEOnDM2MSH9Qgi2ID5+/Otd
49EMv29k2flCk140Sa7tkhgzVVk/TRjFMdKPlbaYxYZFDNZVVr/dprDz2a63pStH
fGU3Tu6lCOB0Tep+hdQ45x3tTAt4wY3Vz5VB8qWzi5yFWERaG43fE8YlrkltVAkW
LPdqPyUAJdsjg3nlYGxKUypy7Ii7aGEpLa07+jMgDDJz12gtQ5sbIL6GtStQwsTQ
1L7F0sv84cbdfEtxIE+hu0nvyQDBVFOEluNrZ0wyVAYv5GJW6x343LzPf8hdMGri
Ca08jgXZUOJ/bH5ti9E4uS+rg7XKTwIy6f9EMXz1clHERIpJwkq4IEJe/i+3vWi+
vn94RGe/a3mBkjFfgpurz9ILF8x0rtFN4eNcg4qMWhDuAMc/Ottu3iuCHF/4q0r+
sdhM0DFav66nq7Tv9mbAhnYxiU2CnzB8mZJ0juPLawdl/hrpbaOoNVOGyMScN9Rp
nzAQNvTOjjmFeULF2M0ZOS4z9CSLCN1J5Y7g/xTUZS6T9kvEmIdmvCY/iR1w/CPw
GtPGtTErrDp2JOMQ1RdXzdfcaUW63oqSSiBWBpRxa1tbLnSPieKSfsWNnGbRsTMB
FQPTWkBT0G3/TtMJCfiSVcc0FzffJdFUTFwRJJRyoaOjqjyQOTB77aqCSJEyIdgi
ORolLYSeP2npaUk7KsSMjaFBcHWCRk3zGHc8Lt0HMXx2UmYJJIMxVOUGJXqIn/0m
f4TkH43pETVqnIuunCV2f+NGfMuj5RQTHjipPvEv16HvK/AZIv0XgX5h0mNVnP6b
jlM8gyBsSjmy/geKuTwKtabh1cIFOhzLIQO72hB4bSg2F6XbVbuwnG+fCW6OIofD
`pragma protect end_protected
