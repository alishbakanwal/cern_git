
module ax_data_issp (
	probe,
	source);	

	input	[200:0]	probe;
	output	[202:0]	source;
endmodule
