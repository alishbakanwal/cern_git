// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:33 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oZeL2VVXMf/0HFLYygObFo5yCP4N82Cvh28HFIkGyKZCPYkgwpXqGYX9D+N1SJVr
FKNDwQlXjTJCj7gucWCgcs9yv/plHB5DPibe2ALmFO3flivTY1rFS1nbPofw2flO
f+V/VLfQ9iQwie+DK1Bvp1ORflUJwWG+NUomnzg1LPI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5568)
oQgAGO+TpMspGZieoG6EGdNDDZscUWsBksymkMNOoJZy/lj5QdkFSdwS0MncySOv
LkiP6jguDneBF6ogiLPI2zkU7vYzR1mrsComBVRJ0pVWt7ljKi4Baf1vNvLvuC8m
3u9CEAxKPYlqqeaJN/5T/ICsJjDXzCNaMuTH3MQ4dmj5M+clzxxvEgVQ8oQ7H9jI
LRJbXdlrMkPQt/9Jwd8f0KfJn8XvOqq8mFydJmzWPk73bTfx+8jNwlV60MGhK7EW
F0FAy0CVvK0Y8L5os+G4ndo/IHTA5Jp/0vUS0IG/x1qU9Re51wu6zsfTx9/q3vwW
5789U2glBdYFAs3mbcepYgchRzBp3QaanFy6YN4yOeDLZKfpnQjS4f620NWW/NuV
GlmOKjP7xr+yyrrDGZKUR4S+8+QCuQLSO8mzKLRzKOvWqtSOH3Szn0QzYdAarCsS
XCcIgqPQkipc7maz9+QVBwEmIDUNwn/rPGAJ+Aca/5QhS3tO8z5f8kG5vSZzm9PZ
Z19t1Qshr0q0A/47O66bQMg1JCr41MEi+qXMpKkK4kATvSz8pjmF3BGBAJX0E2EK
eZ3Er80+mwZh8DYsdYAGun7mnkRIeeU6EsV61Q+w6g5pe5P4PH1VH8Bmk2eivlxv
XGbXKBxHhPqeGVm4apbwtk+R9ob6E38oPeidj0fBqHRZxcv3JmQpWhNyxTTwWFQJ
NTww2EFrEvHm6o3cLwLgcaAn3cXzF3f9yT5TLUSmE3cAFwyiHqBfajFpue28/51v
gh4dqAjmkIoFvl69y3khGj6DDv7rrP7ICMfsnx8ULV2jmQCiW9NhPXwS2eNWhTU6
RqVeyOBWzo/zlFLmKfI0A71km9hcJwU5AqnTF0O97c041lf5uj52H7+53MlSWCsf
YxrQHzdt4lvsrLz6QS0onQeqtnEJaEVhggdydDKpszeUx65OC+QFCKapo8Kn1VIF
FxrS5CmGwcUHoc1+UUqZNsQTUyivhJl5k++msneR6QEHOv94SguE8ExD1IHvwTQo
2sRYf6Z9sfoi0IvZggMu+LdkidqrmBlphm9wTMRA/GJWM2LHxN1LN3hBaYzvbAAh
u6r6CoiBRAvnjIYbqXPqAhxh5ZBDaM0fKnRr5G+YHIq8qYyF9sXvYWhzdh3+8NdF
X7URYN0duvT9F1L/rxwe9v9NJbPHZMM0Hz5Ua2Cd/4mhqlroabsR8XVLmxDeig+Y
8iEW3GchHesHaq5bj1KEjs2BUpqTxo7DOLOplw2q0nAjZAnff30oef5utiBhnueC
jBrO/vZcA3qFYDiaaDSeILoh3YkpVmS6J4qh1Bvua83i9O+lZj9bbHYDI4NSB+7k
X9XbzKXXpkyB1aSCPxBjH14N4F5P+IdgRHHkUQxW5LecCH+4OS42epO9vLGVIojS
2NUjxOF+HTJAUiL/X8qxiTbUGpP5LkEJ/NXDGfdYGfJg6q4OxCVuNkzg0NFDkzNG
Cr9ANEuXn83xoq2CYjvw+0AWmxYHOacZwcw2ig4UFyqZF53YUT1RWEXz6rI88fMP
4yJVNOZTCb7Eis5fW4LKpe3cPX9T7Le9xg3kAlHN/yge6D7uGbxeFhAaEbisM6ur
UvTQDmAjHDjjJGjUkfemcvK553InRs/4FNM98L+4HSvVwdhOAJoeure7XqiuAMQU
2R1RO2bzeKYgLtBHZkvytiW4CiveCovebayA9cneD0IGGuvKHS8ZBMa98FK+Jati
C1iVnuZRam0ud7kJaSp2socghtdJ7gv6BwByNuW/cPOXk2uI5mcEOVX3s+a2Wchu
qmeEh7MFH7VajqZKXWE3akAVO8OZY+jx/CXTo8mZqNRjhn3tjCE292j7cK/M9L9O
uSfWgL07eQ/UQIJadLp0RgqVUO94QMGJuSRrzw8a26Yj9d+ZpzMuE19nK4N5cU07
M2P8x8YkZFkXkMwiu0E+kBJS1Eo8iii+yVus4nfMrjCjcZnjB2hTFkf1nA35pQsi
rrbX/OY0LlOR84IQJDGANHuMlOnJEk/Gun57ARMt4SghtyM+fEWvMyV07bTfUrH7
z3Jw1EnK2p+l3qSL+BvnJjeVj5S8MJ79Tn5H/2QL4DSx97mEZiB8FKSX36xrI+Me
jEjuNL0lCGwASDUsPuHqkTfnjIc1wavox4vxLTx47IBBk3RUaA1GBGjDDgXUEyRX
WBwkWU/IgAHlfHpN+9mTZMNRgLXXDGFj5V6ljEqR/YUWlj4KXP+ifpR+cIsB+OYG
kUd94/S8ulJZPoh1lAzS12a9woPIEDyPf0Y3IUwqhhq0Z7907kOpYpEvmqa7iuDI
VSiFL9C8gLIb5CRLV77JXNjsN2MHoCGAGEhjsFrRBrcrivqTGxD/jUT9gtKz4AuW
oKQadKOD1vFHBEPqTBsHwhGjZj8iFvjR0k/ZarDYYabZq+M8xBONQIuETFGLOMjO
ppr54i1ZqpqCONAWOh9t3R1SoRmEbh4R/c7CABE2GH4s+9qjTT4IquLF6WlA4/zL
1Jd1lpiPHsuwAk+Db9dldqu0zSgv/zZXYJCFtr6TQnfZp8PKzoVurTdNecpROLiW
qgEhl0rZ/rxXbYWkqPx7N99iG7w1dHHojCVG2Z+NF6baj6PZPupPv7ePQg/tCMgC
sDNMFTGcYzLVO1cx42kYfUlA7x5qGAemG7cyg+/AAGdIMWfqVk8t1o+AsCIAyKLk
n8bcQ32Fb5OH/y0b5yvhMCl7forY+T7SMtedThsFT5qfx8qtpEKFeexmVBXgVAnS
1Xdb3qxmaBiQm2GkOhgBraa4t0LzS5Dumn+IqpWHdr6IzfuRziS1CnDNzQO10bJa
ZhbEasnGY71Io9D8kYZm2xHvJ5MS0879+NAXp64mTBZNJoHPz/pKX0r8ybQ9vd/O
na/vSIK7fABMyj1WL11CnxqoalSGov5JnzWIdDJaTDJ0vAp8V2vl/0jXYdstXzMY
wNTbJo6fzytcteu/UQ9EenWonF/AhEzE2jofcwDQVnzu9iG+avYJsoijwsr0QXV0
wNEcF7Fx3U+4iU+PSqqw4EntOKFoFySRMRBq39pVfGrqWm1CxUtcdxehwnylR8ft
7Aq/0HsXHv+VChwxhTVDzxxcD2G8fiuT0THr24zWzUfxSC/Jt32Lz35mvY+ZoXjQ
xK4blPFZpY2WvxVJfaInnzOgsgAcp8qlYFJOSEmS4bC1gyiuZqCueu0CO1f9mRLf
yvENiGqgCo5lS4kRWYU03Us/Z8Bcps506knIcMvqiMUF9kVRz+3g2Q6j5ZlII8gF
BkXDJrQLSUUchMjyDurF0618x+8IzcsLKrhkfXGC4D/nuCrBw0hBLmIPnutp4wkK
qnomUaQRVLN+KchG9NnHIeIi0xrA+gBMqBw3p/z/BqQ3lqBgJ1ToMWSlvYTP2Jov
GAIaco6bn/mZfRN5WtZ7mBRPNbKcJbJzOhMpYW0jNSUQVE6X9rhRE+J/yROmH5T2
QGm7Rw5CwT25DOGVsNv+9iuYvVsVgbbZvoAtoyDSBdWmygQzBZwQT6jKPMMOtddz
UJmt/XMKZKJkz4T2teENHG1XnLHJ+2PLk90W1zWKOspTOeqcd2MVnhXvUDYRammk
wH9e6uFT/z+SuWPemRHLYlgbGwlFh8r9Xhob+La6xNDhVgqar7m201fhrTeQM/cE
ndCz9OUkxhreYhW6s40Tl9TveJjccDMYvRPbKcR4MAXQSdN7+8o2q0oQZfrS65ri
Rl4dcqnW+UPOecsezAS42Q60pRHWW7gEdgbTcR82ZekMs0/fEC7mecKgpGPKpM9q
97pRbGhQPRJMpHB574W/7T2OhzdVuEMBOuh0g5O+mEX8JKz9zWZc/5i3cnSoFvU1
EIWnkM1TqRjCp7jJ/6cqAXa/oLith89AhpR8enuylr/H8wQeQgTqxUYGznUnbYso
rQhOYvYqqFZ6+brTyLax5iXYfAvJU2ne3VWm610VoCKMWqI6QxEjecLwqR2oG0ml
TXKw80BaByEK5EbvpBwHKP8iPUt3miUrslWd8Oc96RRT/frUFW7sb3gQt8P6Vuli
cQ9EJFX8HiUshJ81ly+GKfkQqmRiIn+4Q8oeOwzU+DkRmC8QFU6ux1la/jdxR7hU
Nd/iky0UIroVkfG7/oJIqJsvm2WJvgFfSRWA/NZOgl28fWhfd/hJoqA+OB3PVFe4
dqcgzHxB6+67ymhLQKsHbnXLZyoWSDJDidhtxPQoEAb8KH1/+aoVtH+jgPOJbeAR
OqGzMn5DIqkhVRq6bzunlSplinV9NoKz8owTScSoPDxBarGb625/OmFyxlfy50bA
+1COFM7vQK7GiQSPoY0JfdgtL84pxmR2MVtXhZpZimAPTTAndJ2K/b8sCwxA7tLL
JPEuOMGh1deRw/dK4zFJUTRK7mVEgsu4InjHNlW6R/w9yoNV9yk13byWoVG58q9i
vIWpocJHr7eyq9Lx60HjT7f/KFi9wpIXjLMO6L15nwtGUL2UXZhbZWRwIHHHu9kk
aHONnpOKL/JMNqeuHjBryVLmbwUlcEnMHDvsYun47Dk5vdUckS9E/d1R5FP19L/m
q8xJ+/iz1Opz+9MzVuYyGYnOcm4lc49/uwtN1HBjGv+ji1UK4NwOAAowmmYJrjd9
AgUVTxZPSpLDdpPLEKurfcqwq8bu8q2sJ9gWMv/OmKaE1c2b4Kl7YM7b1+nLMxRz
xaBlEkROUg4DPDKffmQOaQsosKh2KpPHurfpqsfnVJ0kZmygs4gxg4b/kj2zWdkJ
etAqKx4C2P4aDbqkc3UmBazgK3qXgVfbtDwQRb9nS64pDGmgxtYS+UniCvrG9nTs
cN9axVzWJ6YIkAAcB3l3J9UjkGEdlXcqvexIO+/NkuyIHkpPTSeWz+FH/O8mUY+c
VMfvImKgAqvPCAdKQVdP13Ezd6ZJQQxdlnC6qAwiBXtBS0yBXwu5ysbuL/IoJSBO
YgIctxVydtZMS7Ozw1QCk5G+EW5oix95R3ee6LziK/bkYLNwlFs4Di/tWq9lyKYQ
nd9j4XxuhbF2olDWN6Um1H+RbfdSZ1bUruZ10La7o9yM91mrct2lNqaU5wES5YLp
vKENKgQCBOAUUM2QF6SDpl4HxKLFMSqxMLdo+SeaPKtRTIBc8ZEj50N2ABObRQZl
BfSUWKK272rqotg9JC/CWXm6F8nKRzwZzWAku8hZ21lYSOvyiPdCUTIDUgOx/DX9
FNa19bA1OJaBEmYnj9HcYeVIaC0k33RrGRmLv/zcuyhx6R+K8T09ISk6gFkHCFg3
fgf6cVBiXJxzSFIOJhtwzQGlStqM3UAumYKHnbP3uZzysnCjtcJg9ASKoC2fQoe2
yEVlA026i88Mu/Y/hs/GYDlPL3GkNhLSLcz/72YqeD61IMkAeew445eHeSVyEgZb
KlJXST2o2n7NFys7a4ypsP0tYksq97KjvmjrmYULVPz7JZ7Vz58HSoUJVKAMx5Jt
wHQcgOY3G1mSBN+EbDvXG1zEr5vS/nBWeXV30xiy/SuBK3/EpHlqj/A0/ga4087e
uG3pvBrb9LdVMQ9At7fVwAAzIQC1pC+ohOD7Ovc34kfxRgvGLKlJTbCnEKc8WAqn
1gsuQq9hP15COFTEicZYbQCmEmZGYHbFxnTrjHcGRfGRQIgKk+BkZHiP7L8kzmWT
hayXk/0qWAK6KhNrPKQyRjiphfbZUsFk+wo9i/WjsmMynn+7oQ22x3k3i7H+/YTk
1j/vs4iuOxsR6tlOGtUQiMrFxJ+tarUAoS7zUFo47mgz5S2PiD6AYZDtzywm+QOm
1UmE6DfkKJcH/tfAHxqMKuEHuda0I45cY4/59BJlbXJzBdrgEevc5+o9BLZKkVeB
f/eM3KOS4VKsNGhJbxZQ6WL4X0EN4sMFeoTtWVtbYL/1wBkZa/3dXk9m4ymFeBsV
D1RsEPJnKctKKOL63cfLp/0NDt7Lo4HN8dyxx54J6b4DDY6sDVv3RT633LBiN+wM
sAVPeKO69ez6f8Bvh1lLCPeWVqkEgsoklpjrqOgur8pg5NPP7h05zMIDRbHuLvB+
RNwaHnM4rLHDrpXZKZDtaD3XayXWovb7L1JLLPUBdRZ/eJr3gqVjwwLrEhAobddg
sMjKnxSEmg+W0NDSzpov5qGyqL9jYqsSNWybZ8RQ3lZmUbW3zk63k9n1AXTpgYJo
HLYLrUGe++EvVywR/xulZX3bF9GtcbyCp+Z1/BlalEREkocjrJwP9lalFWmCGC5i
x+GxVRVuwrLv8viKkpojcg7ZqlkrHSoqY/MZ6kDpp7WJ/c/RyWcX1tSpVdXdWSkd
8rgfHvmSplUSE3vNoXR2Gt5DhWQl0sm7UstedvWUkLSkh6zvGogUlt8DB60dSk0s
+A7n+0m1wg0ZuRJC7meVv2AljDiDdmqknJt2bFBiCI7t/YJsivSs7MwmpW3vOxZD
55CvXpu+20o7wSI8iV6AWBMRQYAbqfS4B/2FkS32NH9eOOSrEmp+5Yda8yIswadU
6QUg/6SIP+PFYouguktskkQNX2etbQOqD4S6gLj04i8Z+rPpNg2dBXMI86+oGC3z
qS2wmOFJHeVEZfx69bqK1yd2yVtV4Xwdbum4MzgW5iXqMoWmbshv2z0cGVGGwM/D
kkiGHMkJEXNwd3Gnsq2wtkCgOww5XPSZ4WrKYZxfgtH7o+GTaHcCbfM0YnvcSGOP
uGk4ALatIaw6giSpfTjta/Mu4AVO9bncVZZpLm2kr47sZZyI0P4tLDoW6mHRFLx5
yLJGyeqI2hjt5VH43uT04tdAtRplZBaTyJIO6pPri1u0cyYq3DPDtzwqPvO0+0Et
a4NUzy5jOU0By0r6v/cBucUSgRNug9rxTjjZ9bM7kke32c6wHqPuwoteBdXp8bG0
mvcb0TmJHc5BEhHpr8H7N51wVJq9SZzku7FQad99JK3Sjufz+AOBHLLv4fUi6osP
t+3uaqahV7ufbCZ393iWe0SfYrbvkoPriDrrf/+S40+QNSxi5STDgV77I6Z/mDQ2
Wx23xdE5icDowuWA/FJ9Q3ABYRU9ZohmrBmM0YDrTjOIf/5Wm3fbg8t8ruhLx9tK
GLNhdgY8WhywYgjfL/UexgHLxc7sbKOTAJC9Z1/x7Wo7lxn6I2qC19ZcnpiLry87
wH6c8ieiEKnTmHZ79kMN3iT4P0DM6T+N0G2UZnSIeMxmSfV7fpb2LomETyjINWFx
EJ1sM8lYKZUk0Z2ttHaMAtKGEVSsogN+zIbVB+PhpQSJUYHD1GfQQCoY6mfMEr6j
Ac2mwvmTun2GGF04t3pJEg5PgBMyhwMOIXbpNCKhckydNUvajVXZjOzTWLcCNt1p
H8kd0vzQAeJwXO4eQXMz4u16mZkuL70VD+7SCdBEPMPTVgLhvKn6yprichwX2ufX
mlRNcewrCoZl0leBhWEP/fpQiaWBrc8jtlEvakg3/eyXudgQwT0h4P6B+TPEnPI3
`pragma protect end_protected
