// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:31 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Zt8aRBfb1LClBCBojp2xt5luZi5e1SQ4Xfh+cqiOkR//EmJxVSpFHFXgrDiP+7ch
nw1JENL/2Fa3S7XBEOVvrK1Zn8J+OhruzkV5ozjeJeCzzHOi0w34IpjzxDzEcGDP
qt7V0j7upM9WKHotqHfkSu82zoHakSVUVMPkHFP9ZoA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11328)
uwwbaAr7h1p02ViEH1p6b68G42z6ZzFzxREoPZC7lniYjAHgxeVeOo2pHSUMLBPX
sNqOV2FjW24lnBxdADQBSDf6JRSoS5p1mUVqO2lLB+9T3k469YJeD30BCJADJs4M
ksnMmBCj03P/5aoG1IJxAg/FajBEvBenmLoNrwOXn0LFX92GFrs6AmLGuKEMhkJH
UZkd/IL6FgEoguHCQmhE0oUAuThnLe490O/Uy/kHcgmZJg9H8J5S0O3h1dzHeXzD
9B+rvLUUPv7zCHJqriZsATknfAA21uvH7qtzEvF0ritGEnMZ70BpkC2NnWw64yCr
HmnUj/jpqqZIlTUF04CMifQ/pxPEKMXl0jwkJglNT4yPuiNBEsOn/+hwsJdlpJqj
cSJr/oVsSjdX4AZdw3lqv/f1J+ZF6q5hFquF6VeIehaZFZXqZWQG/4y3Ulrd6MVw
gox3/5bFtLoQ2Fw5XPbAcrVecDCe0dh5KMkC4vPXK6LvmhmCl3uaI1gsBmlKdUli
ULTLEJZgPpuVlvzgDkSazd4+neho+h2aOq0qw6MJtXrofgNBjQQnYOe9nK28nwC5
3DtQOVLsvEHYpZhy8M2ASBlsu0pght0m05YLUq+mpixa/LhCUhXJNj95x353+TDz
YSmeNu5X0ujB7cEGEDkbzsNIymLZF1GcmpZ88cup4/vYWQ/AKgd6OWM5KqfghFVV
Lo8f+h7wkGatzOAmGjAmyg6zQRR6WXzh52YsyhbUwwRcIWCKV6kzSn5h7SSmI210
/ZmSu8IpA29aYz0O7+yha2x4b8qTS86URtrCqCmWop6y0vTvQKns05G2T0ZbJTrP
Sdptp0o1lUldw9LkgPtviOb0plhHxeM84azm9jRDjebDJTh6LIP00+ojnpi1mwae
PpzoEvluMxgehKF/+5FqXieklBHBVxUnsyTQ2/cwIsNoF8POGQOzTfJozgUhMco/
KV3QX+pmlabSEXNABHtUEPXy7fgTPFgMxPq2OwtEkIXZmXMwlpV1uqGZZZ3DHaAH
rS/ZjmTg6I+8yl4X25wbmw9wMPhk/wa8c3+sYXV//UfANBBSnuICRS7fiKP/lj9M
KJi/ZZRLSAa0QcGSt6Jwl4dF2Gve1UzxzfVd/uFY6XGJ5qTmhu8TAEo5to0kDXDj
GMsA/vkOc5YkJ/6GYNwFgkO4hx6gquYewFWMPODymsj2szzC7b0O5GAEKPiY7IUe
MkRX4UxZPqHzjCS5EzOTixK9RCSEQl5KYtzKrvLirYAVoLqd0R6MVxsluXk5TyDP
049VljQhw42fEtt0sPwS7ZfmkMHznwPMKoONO4In5DKMFmOEuShtYjB2JG0EvZEe
iOhfg399rZwba2iYw04nw8wm5iMTsBqo1TsG/l43YR+xSuXecomsj/dghF92Tyxe
0mcWP94zrl4V/k5GvWJGdjGXimZS9DF2nVKjx90YlZqJHST7lOGTtqnEw8NdUIv5
qMOY1eWgcYl1b0vt0K1Jr2LQZ9uxdTuqBw3Z/bsm5kga12yZt+KoS5yAAhwCki/G
3dpPr3Qg3cwht16LRJpZxPMExWJ2SAKPisp/jOHjGypGaEokcAKe7OfBvSpwyzBc
AM+Fj69I+dk6NDwLWduAsehBAkXrEULZy/sVLyBXuQRGXGpsd5XXrwnU1gkap2/1
dlG6dSqzA/QBYZQFLsguyO0yPdSm2TxqY3I8kSOHUDPKIfHpPYatL+ufEOtW9KNp
IDmLydYvXx2BKBzoG3kwKAkJ3PmJvuLa1uhHDV+V45c7kV7KxUpTDzLsPRfms9gn
gVPAcpPyvxSIYe6+FKCz8HZjFCRe4oouMSjDrkXh53RydtrVXyEVO6TAT6D9royn
kxgPDQCBgkV8397b1M3qL3TDb3QUry+N3DoEs3EVkdu2E+kM92uuxoESsXaNdhOL
nfRPOowLscbmFWuyUJwJ25M9THFpiG/2zFEXP41PKby0gvvOrG7AejWytY9iu5y4
3VuX27vr8qEcfFeATwI22cN5ATIVge1l6oZitZqDCbWJXJ0Un+NWL97Dccoy2OCj
EnxlGefmUtlsOJ0Pmt9VLAoAdIu2ZkNixNyEODIKaizgtimWkYHVRUyAVKHB+c25
BEBQvzxb+UqOmHq62XcE6C7vxNTWSgZE7OmvdvgO5MPBVLEt8ln0SzIwXmDTMV10
xd/79hSS9MBwxDOElFZ3BtMK5FXm4oHpOZt1jOFkLTjpo56gO0GpGpaU7xioE6nO
htfxamsi6AzQo5Y+npPUrVnZxFVam2POmGmDA1K1xu4XOfrpjThLs8uLHlGZHleu
QVrbZ1c8FHq2mB7xgGvkq/WRoypg1j9MKD7xlRi8OsyJK267sqnNF0nt7z7vSr0k
kLEYIg4pRbOBbJirindyjC1mdXd+mN9rYn7kG4BboCrM6UApChpLMtIDaICrp+gM
7wIo9aGq8y4azxQXjPLPh9cOes62FNJREaCNUnXmlYLufmVMMghby0xXgDH8ChSa
rwrec3F87bxsG53inSAhTohpbMVhEAPlKFHNZV2y+Uz7v9LCltjL+bhOhwC0yCdS
OwjiGFGU72xACr5n0bZaJZVE5Z4rBTzhblvY9S/E4LDr5FDeQaLgjV+57MwaPeou
BF0Um4eyKiv+XGVldd9QLWuXTUWtRlTcsRUL3PytDlBMDxsR8hLgi+htbrmSPgBi
qev0tJ8I1OQmX/QLxysuXaF919ZXjn1EBu5MMOOVyfY2XRAzjv+Awc8VbemX2SgW
tTZclc7+7BGegRkMvhQ/pjgEdwHDOSkrzKyazcZtsYta3R2Zs2lt5yOZJ3qHLzbW
gShmz0bgUoIMOa1bCgbKVN3zbVhOGl7DqbIsST8WCzQXrhHZzJzzb3h8aXTnWCJW
GGCrEEcAFWfn/U64fGmOMCfg5G5uxQPS5W5scgvLPGLc1z21jPjMPsjG9UmvRXem
OFa/4rpWT0Orua3tKPb3eaqA7yKRAlLI3bciOt218dT5nx28T9hvtQr9fiS8o0Zu
yHcAni8Inbxje6uSeAxpw1HA1sBVBd0U1/qF2AULLgxyZcFj8zGS4+sB2WBSTQNI
AErelrhiPhA0Pw1ejHCJnMOMOCmkVI1rzNKcBdkK7QMV6uiciP++sdh/13qXPPPw
qXlRyeFFYLidC6ZH1pypMKS/XdD4uN8aCI5UtooSOqYrKuU9So64tho5t/v/rLpP
dO7P6exXO+2tnE0VPpk4bqIfGuic/VqDRyw0E0VSaa2Qu9P4uW3n0Z9p7+bwxnuT
+BAWEbNy/gz2MaQQ9RQdhCIQy4mdqGT3kgldQpZHBW/JjbAkrjfR8fSIJEJr/zx3
Xe9/wP3/7njtHkdG03c3rwuyk0g4oJR+Exd5gXzG1ItJVCfchlI4UWyKF0wQ7uI5
AtEGLnk0rr8UKPblUpDzMNaTVSAE/spPpWGTDzZLIZOvs3grt6NBhDeBMCkZmvje
FsUvcgggd6CUQab8iManO9Mju1/4MJKWlcmLeLqC+E3Dp+ZyttkhuLtxbs4IzSf+
gbuqtjmf/4kWlnRibUI+JYntBQdrNdgZVGbT1JlbV6pDM4mp2Fizoukk4/bHJzVv
P+IbObHZga0ccvgowa5+3TWCSkJx2TRynaxhOIlPzcBdDI1+FWp1fTFuKHnHbQBs
rNcyOXOUk8//UAEQZwqQszmwYNLJxHToIjqH55RbPFsFTYig1+w/QePBm8VwhE7e
vxqOyjNkWw99B0O3JXzhCnEoSdXDsQ5HuJ2ZL8M5fX4uQAmTxpPj1PUkouJd81Ib
DJFA0z7KHYfe/4XzZfPxRktapl7tiLGmPXiXcE+mcjyxqFBdP2AqYQgAeNWwLWiH
vep2bWKga/CT/wkp0Qy2VDYyuE+19ved81fNCjBtabA0hMBZmeYGpef/LB4IZm7t
4Rw12qBtNNKJhkoLk2nyEs5U/AADtrd8bW2jrOut4mOo+gm1tOuLfRVrvVNDoZVZ
PJBx79LnGqBomUOW5E+EXw1j3puH7hfiffwCkpCHuOBE4/SkJeVrxdEDn3y+szFj
KJjoIVLEFVJX2hmwcwMhEnsHOE7tDE7Q8Dp+kyH8GTq5J1sX1jiH7Sj81VgmuC4B
YUkO2+8d6wPl9J1DVVVJoEQfAb6uktIqcfS9RyvvJ6WovvRBGvoyDzw9rt2/5tU4
7AGL18RaL0nsbc4IqNBWyF+dN6qacUr2zh3cnAYaMp6np5qqdPWHVNiJxf0iZicC
pEtKC2SDfFXTe/xF8OMJM2FUscNL/KrinnMQap2XzZPq3Qy3wD1vfEku8Y78novf
UL9HVV2Vo2q0LlS8MNT06mz9w+TlwviqUsoPwjh3a+Xh3YTs1zNNVFHsTEV5yvXv
dq879ciybh4AJq/2E6y71VpFETX/PqsWcxoatSUIy6oAcnN18jlV4a0PmLSwkWsI
mvwL85bCRplJ3vAotjJOsDIh2swwWtUt1T30G6EPRYekj3l2TP/S2IqzKVpskSI2
xDBMOvCt9SeVdwnh7kifUWT/IVAYLB9+Xpjv1bY5y4okwMGH4qAJ36/TEtsFCK4R
3L/SvsKh+vKvsKC6tBFkKthP4nOm5rUdk519D3sxRCZg/VBhywtrHJFYg0n3pUYT
G19bpfhzXui6GNhxnyXkfpUAfS/KGrA/MN2JaWNvcC8bx+fFvpDPJMlatMRHamVB
tH2Tiuq2X+Snc1VsYI9tCINHujYzdjokL9KZjyFAGb/E7jr7q+H3/NuiM+YI6+n3
Gpe634GPQZrIFXibfdNgOAII8I6nJ2CtGctxMm3AFULb/iKWQzRVwBlp+u563l3o
ArhS0PmBTlzjiwlF2RSZFpJlkqmDPrXwtZ9zFskf0JadaSKUR5R4O0PkKcM0W335
1P7FSD6kqqatHC9/iK4Q0ocm2jNKh+OD9bCcQjntMGSVi2GOUR3mV9C2NgSFm9B8
hcAWbsDLgt7XRmNKPBxgY6237eBg7wcZBCjcT01RIvAPtSTDM7pCpkZ0BlXAqGJN
yw8tncEnjbbdW2ZyYOTotTAzl0qqg7kpiEIhQh6UrC4uKKJDlo64D4Kj2d4PtCzG
W64dqHOwIu8ojandZ/FmJJNOa3/Ln2zrX+jPuIlE0Y/StBmdQryn4mwOK+3VMGtw
tJCiV/G+aOlTEyggpNRXyPakCQWK1bmCD8uhdmCUWcmJgXtvjL4nU71Hy+Hrfq9G
6sXGsSeOABjv84KGxXEd5Kp+ei4XyHy4RfvfBqLZ2AO8hvAKtMvotyJN5PHryqoU
QDKQ/wbtxoR1j2EcEL0uUzaSc0+2ihcQdLClGZpP47dDnHhPsHENTt8p0vir61jL
L1DYnClp2hmygw+FGI36KK5/JKn2jZCFUs1nPo4RkqJeXFqW34WOOVGpVvSgE7So
V5Z6KQo9R+WqSuPQA4I5n56EOWPT4wQOYbkOaUKWcSCmv7m5Vb6GBnnA7V19naZM
tGBZMOKlfdDdgp7B2hceAl3b9Osm81X1cJFR3S3A456lIefJxi+eQx6hiXAV7D7x
CAkiyRwkMcOzG577W0ZJ6fBrbVrGSx/r22Yg8K0zupUCpUFkWdU/hvf/qDbdhMo7
YyOirf+SpMc7+dCcLcGhVn7YXky+wTzyo82TNV4H8MzeOtkhPGxKTRzk2WfgwYra
xYy0A82zpbhRjrThBAwrO+UUQQnuQcq5EVNv0lUHr9JV5OBNxXYzUPaS70EkIAB0
JGnAX6ewBCZXoJD+Hnq3zpAJAm+MIo8QrF51OoWh3hTuq+wGZ+AQ+9zNTMEIE+6/
3VMLK5jT+S57RUc+E4YDz4lm3YdJSN1vSDay7dDtwBtcKHJBaDOdafN+CokAgy+i
QrqRUcJtJq6uG4P6vyHSHQfPUL+0O/w7UTBFcc8xop4BwTiJo9MtzUCNBa2df4Vl
JhPkNOntJ/lWBjGqcsjivppyauqeVBs+epl/VBooH6tdw77ZrK+fYz/hZkq1NOoz
nh+mTvfQbsD1Hz2Q/B4WUIyfqZx8KSZi2amSi//AAXLbPw7OAM/YrLKwK5/bzEAr
Fvxdn+5hNtzloqSobY2LrODsgRAI4s79l6VBb2ZiLJKNoeug3uzNU11nEgCgXVbA
aez/K2E3+Mk7Eyg/YzI2M1anvwo3o38MBeYRCIT/A4iw2R91rKeavn2vicGYyxjR
Pt7Ufqmsd5hBx0mqVI7a8SF0YyzYrIe5j4a8COAuPjsAnfE8nK/UTy3Dbfaqpqp0
KGl/6x06MjPloSqukYrW7KUbUaNJ4EpwGspKoxeRZjYTJvNZFcqegRriAoojRAWX
sqJdkdtmhDSdslkA99G9R1byB5fxel9DDA3j8qsvdilaYZPsDxjLHfzG7gt5s3eG
tvgjOhAc49pgCutGgZ6YQWJ7Z5hVDLGMccmeM9mms1uMWW6F2GupeMtZcgsISxOX
M6DnjZMMRUKF+Rc8/oAlgx/zxomelLRGpbMqVAqY7LSpLWOwUYDDDKgxQPd5o/eU
7SoVlgXvi1VFC1Vj8+gWq+X4mzGox4VOEiaM8vdK4zUGjwJFbpvjauAdz+uXceLa
gl/iJhbnHpmhtBS47yxhUPKlUZZZdyq8PT5CuoTQPARrR02vJ5bmXvuVODW1c7U4
9EPuOHuiPPkvt1LMznZI7NT15hJblZSRPgAPTslW8h0PKugwQ3caEaTcXSLzoUfU
bOQyLGOxjOCF1vGKJUZArbFvqq6/1nnm9ZXu0RblkJQR6qCZwqsJqawYYbWKv3jR
qKqcGh8WMFUfzjEZle1VY1DTso+dbRl6i0c4hmHbsMilegMUgdVu7zLv7EG588to
v8W/kS873D+FX0c1hmY2Awe3nu40+LTDGqdlVWWahVaL+Oaw9UtAd5qAioRWHuwN
dHWy9RUlICoYZUBLSZYKWPTxyRvlkQIMskS+yleWu13FrErqZ3VsqXeRtDVW9fKv
iw+vC3bKFuqJDpp+mG9HMO8/VVtJ1iAiaD8gBt34RTjQoE8u6EbJWthVMo/e+Fwn
Tl9avphRvIvNiowWXBF45RYNoVm8zYdV7C0kXEw5SXWSEvcdXzHYKtN1Y3o3Va5L
zZMvUcWYm9Km9uy7xJavFDjnY18r/sCCLX8+frl+yc5PHkk3smjAxSIB/yCwDUc1
H43RulQQ62zRarvswtyR71FhaXXAuzAFOehfFlXMV4763hNnbinOlTPQH7g3gK2M
gnh8iTzP+fqEFfS2rcTph7JF18b3BapvHZT0oIV+ByOfOPv6vL6L6uC5Itmr4J4A
x3uJbeafU1Gl1uF7GILiZgqEOqRNvtGzZE3RFDG3fGYaxOOdMSSOycVsNPDS83GS
M7ku8JjT6ER10wAOydE7vGRrjZ221GF5D0LKlqezalPnO5gVCrpzYt3a1EMIFX0H
a4+Mll1Di8LybWDPrh6OjxYqjtamCS3KieSk65S+XMJ7gqOwCTebOie4mzpkRw+Y
l/L5/VJZn6WFv3Z5GU3rOgr6ySTjxCzNNhUtWQyQ9t2e3iHHjQY3YQJqCfnKcycj
II8ZmK7PXAAck0x8wllKux60VAbP93a6xkWOePtsN7+TPOKhX6d/3LYzaUsbpfCK
AUUXTL5z9XR74ZtZ9Bm8u48qkYdR517dyq6bCB1n0cxBWJG1DGZTkecEqyD4mmnB
IQbuWzRUcVid9sBsob7ESwNnSYokT3w2hgl8XrgsjyMEozB1w88uLEWaRNQwY7eJ
sG17xXl4cT19hZz4Bsc9iYywfGlX6s01zS+XoinN5V/JJUzn1XBg0O5Hb4JcTjK9
m7eQ7h/cfiM+7MgJ7OAlYXS4FuPErvyoLRR7AvxX2ESKMYUjEP4lQpHiNWW1zJFn
gT3lUlhFk97J1ETyzJJhUYYwyM+ow42MJZk46XiZuHOlxYQzaMOrq0I4SZZGkmNc
zyFc1Ptu6iHVp+N8OVGDA9gJRzoc3rIfFfTWcKn/H4o9cOtB7FJfvy/m7qpyzF6c
Won7U5z4QcJeoy2aMcAl188g+hTar6f+9jBTVQ8ftGdqM/Gt7llkjXoJY2L4g9W4
5vY0XJdQERhLvjKm1aNl305vw3uZZht6CMu/90DVXuWBq3bExgitip3JBNHb12J0
57zgOSyKXpCc0KuSp27lRNiN9FB8M/KJ1sX+X2ZoeKGOMZVd2e2GzZdvS683Zf4k
h4S8n2dUPn3zrEtU2gx5KicGaN10yN3Ugrwg9yw4ukyYnLB+NqznA3OFuS8qIKwW
rUY35QH1pR0hPtmWNuwMLgeIsJJc1o5HydBRz+ln7Jv/LAbjns9kdpkdLDzX/ylu
Zxy5BCO4k4Qr8Xy/RfMyT1pjdA2u5R+iO/tcqKzL3Or2gMMV04UzH3nQJSlqm4ne
IMKz/jZNr0e9E77V823xtQU4aKMt0YvIJ3MG8mO6Ra7lKpwoH64EE54ktTIXIPkH
T8mf8c3bKPt2lPqRPAtC5d6WZfvmXfTd/x7eRrJmzA/fHlApHkoUFrCdYei/0kIp
b6lntTE4GbS4jdFJ36i9lekf+yUmQ9mLwufo0J95IvY7tLlAu65Dhw8baAHxp4bL
P4YDdRmXQeWdiX7I4XRBUWcws9MQNF6OTLArYPHFQQ+wbZDD66n1yB2gF6CeIiuO
f2QxGuoXvMxatH5AGp7mTTcgGJOAUlwiJWgR2EA066oQUIhDxsHj5wW92pr9mayx
yIdYZ+zWxkhPXiwoZ/IQ0z/Ggv8WXSr54s6ACbRT5vfeWXREjkBE1QbSAKhaDePU
ZYRWc7iwrQ7cCzzWTB0b/3Wv0CnRsMUdTn2mrGb3jFm91+DZaKTeNMP/WL2MD9wG
F3LVC0GNzNIgWltcW/3rt8VZXpDKYCGtChxobBlivXfU8002/OZapsgJWB+zTMro
a4qHVsT4zsA3hWL4c0YVi6wiqTEA1MdbQolnEYRJ2idGuaUCy2nRsduVJoJifz9t
GnvskJqOFNOtDpO4iXWpD8kmPVtfhR4R9VJUk9uNBzG6lgplDdYUSwuG9C9zp8+h
h4uQjBMKxYCgCAhr6scMblFFCoit8iqbBo4kGHEx7ldWlyRg6LwzSqm2Q8LPKpMa
tl5HfuOu6BuBQttR2189D5CdOd5ddDkyuIzi6xyYbM/gmQe+95RuM9oXbT0/hWtS
eOWM1l4IQYH7Dsl7ardkFTg7Tv8vcnFnhe+XxAYlQdmi5OTVH/ObLiwMQR9E1fAe
jjO/h+FFExnXZ/PGH2qXM9drE6JWVR25MbTQFIlRGUgivclTR5cBHoaEIdGNkAb8
ZggXZPIbUqbjeshvH5gsG8b4U/fk8Q+T5T5qCl28GbQ/iNvfjrsR0H4vJyIg/FWG
sJe7U4jIqzyHB6GGWJr0x49K/ev+/Mq9lyUZ/EGUynC97I8ylw4OSGxRCz8YIfOe
YosHj983H4q50MEz6AhOh3ODT5pKl9YvGVc1GqsQ4LHwegFrgF9+S7y9GPF2dxXB
3my5yu6mictKNgXoRIAxH+7zDx7CKiqYkA7z9gQtAdvuOy9D+2HVzf6c0tU+p4EB
lE99T7CXB6KY3B5bPqL8A2tBsa4qgl+26x9v5ryTkmMxzx7QPUbgNL82z/C83a+6
LhqRGFQ2eMjig1wcVVCklPpZMkSTp8vYNs91SYmNc/r38x+PWlD8QpTyFzaNukkg
z7xItemmu6IFVqBm1ZIGtiYPVQAsNZ+QMDCSgDBnadIOCkRQM9vmYT4Bl5qoJH+9
2tCW7rI4maCvMkS4Yix3/3xXkybDqTEUPJDPqfymFeALsN+SEV1yXebx5x2GXbZB
Z3TzknmJ2GXXDIROITrZwpWIyZXwx8AnIfiZUl3jPw8EMsldl1QcAgQtq2ipqhBh
3579rfPZtTSFXKKlu2sKAUqcHWPvuK066ke1vCta8hgwHPtSEfvmEyqZogMLoWAj
61MOpLwY2l3QD8yxPa+OW2/NxY7rjRBLNL6v87sGdqq9DanvsIQcJEnLYvorM1jS
jXbBB9pRYfL5YRrtfs7NQcp/9zFv4fH7FDVhZ1eNcPYG1WzLtDtHbGwdIZdeUMxx
SbnjD2GcA2eEx1jdmOjga7K50RXUn9LWPnApBVuP/yFQWyHYi+dLV67jq6A0myPO
pGnLu9Rb+SFOVYLz4snII9+NZrro/w+5Kx2aUyTvVsHFawkd6dQTuWPzLnO1TOMB
DsZDC/qKUfGapAUzdYMEKAJEQw9SYU51bqlQOOTpgD4pu0iZEaY/TkG4yKT29sMt
Anjf8iF5lZ7H3a72y5EFttxaXCRKEJhWtOUBMKa2a8tmNhFdEM6skfRAyYxAw6UC
b4WnvnZ25IhduHOKvUrSn5qVo7zTtJJHs/Clz6Se7lepCAloXig6adHqFfS4pgox
3fdnfsC6mg180q/6t+wkjX4rf+8PHE//m3S6SxYjWQp2pLcZzcAuDCfEUklkEoMH
OnzaLRWnNwrzgLSmbswqgRyYArcOiLTipFot6os77Hh3E/OZkKGIfIFcFa5Grpj7
POgc5y7+mey2c4Rm+9eCIGZuvM6wc5+kNVEJQMD9vy2037BHkOywIEAz85jYSSKK
YDXCI7SBsvDSHr0DFmo6Tyx694SniStn33zP8PDzUfBsva6a9vrj8PwfeoX6HDDC
h27PtYooxtiEeBWLBsc5OXyh08rQRNenh2+lIUIenGH2Ms6rPL4gZUqRaJGbCi9p
ScTBL1hALwANrDIUgAmrzKA+AYhcy1Z584dRSHCmSoMzfuDw97uXkBeIlME0e8LJ
c9a3JREZoCqEPjTVc7Rh8X8zrdk18+Pde9z3jmQ/BUDiRLS+y2jO1K/3YeK+YVCM
32C/7jIGa3ebZYhR2aubfHOoYnf3ALmSwGCM+nhDxYMKsnaxlfJj4Q/R8J4AydB4
E3akaPpxb9qbPCGBU2S45Fiet+J7NybzBE2lsABx9gzuuI49+Vd1sZZCXXU6Bbmy
2MoaMWlx6vRWhO0GPEZhM8oENrl5u4KnGdH/g0PzQPbZUpQ8llui9SY9LMoQAhRS
0WsLh7Gr9HZqxxj93eLCzXicAX6wGNuloDBujBCjGZbenKmFIE+NP4cczTR7h1W3
Y6iQEmhMuDM27OonKuBXNQcy32eRDCb2SRaivLeO2lkwy2hg9/Y28zdnXdBof3yV
uCGMkpJ3LpCWvIaMIvtP0OeTN5C+mqxUFTDahFXV0NWaPfUSv7NG54+1JLGeHVS2
/+hwl9Q3/VxYJ9GlT1FHj+vlbSxjyseN41638YR9Xmxk0gs5773eloQWZyUrC9an
RMR+Hbcp6NxtH81gLOKbAdBAhFW4quShcoF/yHr+3bDYGPmukvT9AkwgXj37a4+f
CUe86hE9YbEUaCKStMK2r1KqW3UAo7e+0GO01VzpEVauBrJG7xc53RSp25xyHJOe
WIsau0sy5kPcvYDk3nTVk7lGu0F7/WtMDpXIIF18HAfySPmb/mOdAJ+ZnSl8fsij
WNYNRJZo4dHihrymtHALY46yYUa5evolh2pRsZMtNLJMhJMkjK+hckMpd7AJ8sCC
cKheRmHUKxmArHArjrFNXoIjQTfeFILL/sHCBMjTsWMVNRnLWgOsjwcWsJemhnYl
ViL9IXTSNaqWabAS0dko49hg/1qsSqeH5wSOIlQWzUCTAeWi4JtBRbXt44AxH8Ub
IMMaOLXe6whq1uDDtrUXBIXL35XATN0Onj04a/BdUm0Vm+vlJkaaTJkJqWFCXRLe
GtOD2oF22jPNIpYuJoRGQpY8uWxB+DYXB4p3fQtFAHKAoItpm4hSEB7659iciqVm
MMWagXZTqnpaGallSip9CuyXweYozve9ufxblZTWCZAB508lGwb4h9fDmDA0Ew5F
y7xGgQn8ZBUbzQq+bJhUj7NNIyX6BjRD/I/UaqeTDrQHwn5wNL1Z441JEelZZxQO
AxidNUnTrxTmP0pPms8SV32WyJcQ3uiIRzT8dtFwN1kLLUz2IHxiUZRVVXC6NaZe
BhzCnzs8eJJtwQD4ZGgAu1MXYRs0RD2JswCREYgLcfJpMIEO43VBKH/pQIHaNTlN
127CUbrzYPnMfTFHhT9I+fdpQ2P9kZq/0fb7BCwfayBxmaHH1kaw0AM4JWzWhJ9n
mbs3Hr92yElGdr0P17szORJSGhpbh3btq5mECpJIa2VsD1EfsVtAMFciyZ/u9qRi
8oasTn2XB9gQeyhaQopnMv6Bu/038llJ6xHgtQwAbTnlrL6/bAbLqkXJMU5X5KwW
NRm4plGD/jwCYH/A3VKXeUuAP4sJysAiZfX5+SQfYEoYNQSBX8crv8NTMrJLnU2Y
223BgkHuiYx9jpaGx67qmXdSLqAbVoa7C6g+dMjhzSWLMTrmlxWWgPngfn4g0BfO
74lwVmHnIiEdjS+aS2a/xXBiviCGOwX8C4luONcit+XdCW3plKKOVZUdSYA2+E+s
GsQ6lDxeq8uO6uiJXJF6pJ3rgfSeb+FHal9Q+ijxPMiFnEISUZoDgwPQPwGj2rWz
3VOWDwXtRaFPa0KaJQEOxr33P4pLI2g/oFSWtlVAacycwKup/m9raw5B4n9lyQVG
9664Gmo2OrbP/cfj2GqoYBIY/6paPwx2zZ+XwggJZaowKNCiwR7XokCt6FMYyke0
ZJyc2zTMgLa3v9mZva6A/6+jOqFCkDA5GUMr3a+sob/JLqF0J5cAfNUSdLNzetJY
FHgVLwuoIo0lkR8Vtsdaw4cBsUgLdlpjubdrt+RzEvR8+ILAE/FVoKWt6Z2ErcAJ
vw6MckhSU+Xsd5jjWkIRVgOVLKbKdh/IvnZW+kYCUqynJnt6SGf2CIft/mrcj+Sh
9rEw3qjzJYUJsViqMghAzEjubnk4l3JPwt/XBSxmXJdJ+wR/U69+bUgYkKI1nffT
LeW0tbqYdF+LW66h/zO4SCGc4+uZocWyWT0JCWx3luP64e1Yv4olzR1bjiCHgMCG
tjH/uZiXzxV6BX0TUvAbs+AsAb3Z/BH5LQgPhBqjOpeW7LThJEsWfsAT6B1hwScx
l79LbBfhyCXkXD2M10eFT49boamvLrfDqaeOzebSg4wlkTvQgd8n5hJJrMSTQHSa
6cCoKRCvpes/AbiT7rqf3UEkBMaNDQEC6Oh0hJnTqLi+NaoLWAiQCRFkepNB9/oo
8t233qmt+Tm5lj8mHnzcLc7F1n8FpxnWqGalFKwKZABCz/CDuIgoBClY6/8KuLvc
fi1GrIuhVZQrh+kl6ZIAN8aqQsnmLpa+3gMUPmNIPDTUWcXAuzQgToCOtnO1RogD
w2xzE0V5qkhlJXdPKkMdWJ7F8m8WBP3M9tM+butAEVDodCOGXBHjsdJhFg2jWutt
2TRcYK3n8NHjvWsyqtLTghDMFGnqOMgcBXUl0OMlw+V/GA9gg7SeSQm1fPVXyUsf
a04PmlvMw/HxSJH+fzWUSb30ZpgU5bBrNOXxCy31NuAmZIR6QFnDdSj49rGG8fxy
iKQ9TZpFeilpIztnwhXYFUxiQx0+FpVnELL3oJlYt0ogiQulTDqO+V+FCFDX9oAM
LXFHmfpbSurEorAM5iAqA63MuM7Ju6RijzmLroUEpeIMEDUzNQ8tyMmH/BaKWMxO
5+44rfKoy7Pv1gy3gUPHC322C5WuX6dp0jOfyEBtCPCN2E/p74x5vTkjUyLFbXIH
hNJ7n9EaYD/DGOjGSw6NuS4/EqX8zTdR6nttIq2bDuMMKbWLKE4sGc2DEhXOTf8T
k6Q5ulsumwZz5AqX9CdldjPDTzDKfTMLI92kddoiG4HIzOPu6c5lCLE3rukRrO8X
FARsBeY980DdTyrh0TN91Vu4acnOawG+vnxjIj9kd84hp6BRhsg9TvpW1B5IB5HB
8QIU6MD4+jn3OE6p1tQXlKAEXLdAX6j+PxzcfVSyCsGuYr/2GW4DL3JSA1a2JmIn
VIVggNXRjnJaIQ7a9A5ryeG4Pu9eZaK4Ve45aQ6OdtIhbHj2AAgIsVIeG5Vf3HxS
WOoED68AqxKZIUPo7euUXBr1MiszjwCCJq1R62jIKrO/SMDZ8navyVvM9cjKFeuF
sau3g9MbUEEvo3L6hfXekdUli202o/rSA9OMcmlEnibc5bmpqPIcoGfJhtCA1/P7
sYj+C0B+6SllHdXzfc7WgG7LDjq6b4YbKRwO6gzErqJtjps3jg5UmxX+evtB/KrU
ksbN8eyuBIEG9o2VQiCRsratQsc7Om7seXGr14BkUL9mI+XRoG5/p8Ontw7cp+Xc
37hN3EqmplaMLP8VxCexh+3EtRf2aDdUkV0GK8MruVCeBM8/jZSQy3R7hZXdfISG
bFDJfTUxdVj6Y3WZdlymgTeF70jaL2p73t6klxAK4jMUKLuGOPnZeFg8z701gLcK
IHlvhg0GeedyDgFyxeD9DQ5HcM56b5w92UPxUrw8OGM0sLBZjx8cy5MkMgNNfrHh
HuPT4WEqSvaNcrlpTa/ug5acpO7Gf8AtklAAHFJhbSrc2AZ4oUFRxfFFwgoIMOpg
IcmGzicy7DMAgXHeSgK0nHMpUdisdhaRXl4OEL+ddD2gvQa+D6mM5XazgB6Du+Y3
RSysG+smrbpb2e+LccRpZl5n/g40FNx0va/3F/hgbG/YJMg2jtRoU1Rxl2hwLISK
/BM4c6T3hVSTyR1EpOajyM16nXujcY8r2fAYh0Fk5MT5Oh578lru6sBh3vvp7OBJ
jyppfklj8935nRLTk1IQV2g2sXtfzXhCfYVl1zFII1ch4eM4zZjJ/m3nIV72oeOI
IldAfkipHaR/kCSVyGHybeLh7tX/2LtKTgFCnn/pdwIxa83u6ji8LU1Cz5p1i4L0
tldEYy9MqQf2GUWO3TJvrcwaL3IYMhmjLFreeFQx90ebpG6K+MKTX0IaKWiluDpm
nzpeX/f505mwQKpjLxcOMJkn7x7NU5UlOA5N5GyTj/BoCWKrXsunKNXN5ZlwEL51
w70IsxhHUb85TcZHFbf9qbH97vqfnWqKsENFmVSKNz7jwsC1Scl+ANcsNZ4biVWO
aa0DXrZkI3fI0pl1Ch45s8yEiSTWkIjX33i80x36Kpi23xQ06A4NDzlXlUJ75nhc
dhE3eae8Ian6MqH+71MjhTBMKU7sMUSr4vnAnVs40UmJkYlaiSxfRTzR/AX9nHOB
JOTsQDV59eHZW12R2iPyz8GUxKLjBOQYy5xGSiJwd8d68F+iFOOTURwtwl9j5lAd
`pragma protect end_protected
