// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:38 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
c920bZRRlMJy2GF+TaRjv7L07WZ5CPl2FZ2hPVLej/KCxsD/QgAY/PaAOibhEm+C
hqjXVm6Tm2xVlkdiITrFtkq1i82AeXJ66B0XjmhArBMwQYyAR1PexS/Wqaq9HO69
6t6ySS+DLtwGRQRjbaqzcgLi7FIKUgFlcthOolurQmw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16320)
T/wDeBxNHVt2Cbk0sTICYoAG55pY2mbLhVC8UAfP6Yaq2sojf3I8YdiAkXT05K3o
oVJCoqBcWKkO6k2WnBFMDT736KQ7tVm8tCQiQsbuYOkKN8rFgOebD0Au6hWH+uoa
qOTsEF2hO+bmYs3V1jAu0/FZu8WxmsjY23+RHSbOMNp64OzRw2Odt+DniHpvPNvV
k36nH719f3S3HADhJ7TcFIf4CJd6nic2ps0b45CugJBXTXJBrpq2ugp5NexXXEZB
zO17txm8h17C5/a7QwXcvB6aIGdM/pXxN3Jz5TwGujYOu0bOuEwpTJUf7LUNnMdb
N88aQo49uejSXJfoGzctK+mgp/e5j2L+OCeq8vYq6z1ychHYzIHtjTuoStfGnAVS
tMsToxYlYex3iVneIDo4xp+oN5u6sshRvepy5YdvhH7EcH8uLcPflcaNyopABWDl
fnKL3PWs9uM/yJ3CZ26brdTOJfT7r3JvQQJ+U/YgJpD5az/uvZbkfVOyBjjavHt2
lCW3IyhjPJnBqPOMSuNXhC0ujDXHczH6VO0JWfNsruVmrnse7tRV73j99RlqegiT
TbwBnbk8HSO9CHmJjRfaZ90SCXdVS5aTwv/blw7RoStQpqQS5Y4EQH5HGb+Azu/+
veIx5BIWQyCnK5+gC9e3gbBMsvo9A0NYB6nEKJK8udmRTjGWAgYnWTYX8bHxctgE
GL9Yj8kYKA5QVcicxyExf4DfvtnFDE8iNlc2kXgUuwSQfTGG63s3yBF2+Hzh/Ob+
ml5PyCutz4ZGwoxYlSTah/KRzFsqrxlvwBTU6U+DKA/OFXgpAukAqU2lQOXBFHMw
POibguB1p32d9pxADKFp28r6hyvf1JFZeeNk5soe42K0dxdQbOtD3bmWX89SzWCL
0jX0dk3yhzHigri/P6O/juI5z0lLTnlUu9jYvJfgH+0JFqdPA2NKND5JwZF+hs5s
p71pShrWIoyfowrsln3y83iqxFLfKZlRpu+lRBX5qCrV5A/gfPtg+B6SfrZIzp1h
LYtfFMmRC5stVaAQdulkiOdE9rHZ5onHlnFel/AGLjI3qmXjtyyaPySsgjW30Qk8
7mRA1istoLPhQETDgMfiAWKzlSesmP3EKksUufXFvZa7MSe/hLZ7wIAaushwP/oS
JW794fOjLvGbHrtSl5BGp+3+YQ59oRpSo+WAhG3OJJlvPaZlU6x/K48JsQBADlCr
/L072GdCneKvmqyW/nBNfh7H4PkkMsCkSpSiu6QgsI8+xngJPwArH9OasYw7ATVl
vZ/z5aq7dOCUPtDr+EZbc6ZUDbLlMg8/M1Wb2xDPW6aL+ncYHS4uUa6wz9Aswb4/
hA6dDGnu9nRtODwNlKNiqdtpUKZ9jcBeqHWZRZRn6AEoDNuJeP4B0d0095uYZahc
mzQKHVDnUK8PczmD5qlWGkSAJRCT2acvY9Q/IG8Mw5nzINHbCSAdpm+4ypV2QQHs
yy+560r+i0JqDN8QnEMkrR9QLnwRYCfx+CIXpqHl4uWdWOVYa+bn6+aqHdSuCxMu
NxAXMlwLSpSX6sl5hBat1PCpfHP9ZureixGjpSWTRbkYkpR0fwxUblqS3WgquAwv
/fLTS7mR3Vy8MQObAo1eJTz8yeT0whww5sl2sF82zHrjlajHNT/lP5L4TPv9TXwC
zVi2bWIWbC4WcobLuTxhzUuX0BDE/bNxn+aBeHzJAKx/W8Qm/9U/UOhekHeq7Al9
ikwJRtFsWvqOIILGIHSYPHR6kSwnbk35U+T+GdpiNb3N4UFvlDT3gPWMfhLbk+PL
VOO+oVaYDSyIxoDXZoMfLNP1YCQhZhEoX3tH9/DYFvpJLdxgfypjTnIfyZW8peWq
oryCGWXBfnfT5+O2F1jrtMMGVPs5GnYF20hlAYI+SQ1t5PhFNQw3amwtNixlds7d
sXJsulNRnhsSHvr072LEENMwn8Qeq+HWrfcQ3DQARWw5PRB1fTLGw+1Qfj0a9KJO
wtUnL6ZJs1eFwcOjg4JbwKGfoC5HfL5R/QqhYunz9Ep/rqWjzv0wQ65gFyV+LW8T
c6NUuj+Zycj7pycn3OgEJI09hl/jEdqz9ON6qaHyBFYH1vcgZAEiB4svDDilX3cK
i0cKMIATFbmaW3nMvJO5rz/i+yjhTmwVixPP8v1H8GkHHB0gb9+XRxF9Ot5VW/8c
BrfOC5ycZakHQOlxeGgEJspPUYr6gjvNEpvC+DcYTpSp664Z8Uu7XlYVp2lZltgY
qj1aufndBkv6YHemRr0JfK1cPdokdyYTDBYyXWtxvx9HHq3Wd0G8Xn2ZA1cKa+Kj
lEh/V1Jx1TmhN3X47i+LIQGZIYBbHZOvOKTOpayAug5RPDB7KUaDZp2O/1RtRg7Z
/VkedDHFdumPsb7ll2lBGjD4phFBeBNgNz7HDuhzESwoKmkq53E7oqmpFFKU1m+D
ts0XWMV3kIhELUf3C32oM0Okzn54+QAqbLmvWOg/EThUBB/5Cf2ahdGCzu7PBIHZ
W7qz9I4AsFL9623CdSFRJ840gpaexvMgmzGACx0Bes7hZULQc12YpQGk+gdwLHhM
rHIMIgDKzVbMYSEo7oEJpSeshsoS/o2Lzzqk+9EbHXt6P8P+dSeNIJXdNpMFyq3D
y2TcIMMqI/1FmqMe9dZHbqGcRL3siYb0zsYk2bvNt0ZOtyJwj5MHOV7PjAO9XjDn
k/GkHjntuUgm0uPxnvhVsrJiMbYbrFRe5xsk51DxlGlliaKnvYB6xsiQK3Mcg6nc
ZDHSIPuJ9Xs56wb8MwDsLgIjsz7YjtwF3EGX/eqW8v4MBaZAZFdpHEN5wfNM/AM5
5L60+GAez/vq2rd8nhRpcoxm++uQKRJ0WhlI9nyOcSSz/r6mgZdAsD/zFDsV9lNj
U9uuBJBnItbOuLwojIyKfAvSGi6dEQa/KP1HL7TZq9GMlPI2rf/u3V+Hoy8O88PU
A+VaAY4LYHem28rZtHsKg3JS4UdH5noDGquAoeMvdiCdzLCIiNhh9gidQ2wnTXDu
U7JJSK5ECDy3dRZ18Typ2WyyfXE55ukoeG9FPfMHdrUiyHWhNcM4bUHsitTGb8LV
MwUGcVkPEDwlNncKNc6f5IPfyuAZErDTrJNWsCQqgYgX/P/YXAtOLTaEnx/h69/c
iD4T44JVI9sQjn2iWooxfdE0o3CLLaIGlcjKfz549zjSAL99l6SAhwxufuTZHErR
VvOB8DL39ISZMK24Ui2U5hnEz//PkRPXR0705zgMJKH0H7LQiRk21fcGiWXaMq0u
B2M/PkFAmzMYuELbU7h8a2mvM+iDxQ5x3rmDjMkKKuOyskHWj/K/QQ2lziiGessA
gkNCHOp9dQUNJ1d8l7wqXCQWbYo19Rv47mXpoZZviBhR1MaUFYejDTllGCUxOLpT
dG0XL5arzuAx4nVRLYRj6fUluMG8BBhuaVcBbbCoU8ypgfuWVVO50Bk1ogHlPDU/
h7WmQXXO+Q8Y15yRHcfgV76ZgHUMjW/I/y42fte9kSKu215cnpGW10d/FujIfnhr
/RPFyjYT9YzVkWZ9QfKOv5SL1idysaJRz1hnUlAHAskKyCU8M3cux5Td2uflvA5C
hZPUAamFCJEPc4sfoLqeQ5gN/+GnPJknriNKADEWTn2zIbZxlhROrB66oGGbN0UA
HW45gYKxK0w1wYM8O7OZKTwmuZuR1y6TXTQv6qPpFTKRzEHsOucJfMNe+TuzToVS
LngnIqAh31+vr896+bG+ju3QpEf260ByBnvOGscQ9QyBfDJ9LqEAk26qUSZunoYY
yH25/A66DzNggqcfNZpqcZpQmloYha40u3v3rCicGR3GqNJ8gspqbxQcBC7GpZsn
w8tvyIw3bVvIwdGLnmmGNCVI6WLteapua/HG9+957TAjc+eLGWPlAYYJXEmTk5BT
hcik7Qam25JFEwtmT/ZczozhVBa4LwtRlHE3BB+lqLHecJcGN038BYDMtR/7ZR12
3w66tMCEHwvhEhZGA1S95hhcSnrEtkXmPD4Mn9RVs9xe0LQajt8TBAd9oS0WDUkT
rHjUfnMBP7q136U/DG37pUP8lA3+J5Zm6F4WTnrz6kpScu1GuIqYW3g3JIGp5qKq
OsEshF2223rYgyZkzEgyjRRvQNdlz/AiNLVzTmbh4vibWVBAtHYqiSJstrlwoxsi
Zzkf6Rk0FKUF9H9FsWM86M1/EelEQ/ZNzC+eJnD1ARVmEgQwBoKhqtocQhScFiM3
bk28NJXT5UA4HRnpiO8fBfVM2KufeJdgVTC7OlWsQ+/pnR/luuxbqaietQYkw7zU
QJf/z+TynjojD+54b08i7qhJgqb6hRX6ksj8P8QD27Aouwfl6LXDA8SyOY5UgI9M
PP4MY3cl1MP4muKV8ssT9r/zGfjfia/fEIRrY+jjRG4Fl/ImAu6JETEiDoafXMIz
mORAIhq3OqD7LyGxr5B6O5hC4gQ67QzVUnko1rRcf3xh4Ya5X/4eDSi7LX2R/mMq
JcWV3wqRrR/P8e1CEiA4byOjo06QIlEgzjFJBLXHDFkc8tFzCPQtpdGtNUeP0VIT
qyaQ5hSrSODc0YUwEv4YhV/7+Jl2th4AZPuqfTwBnMN6TjJumyDYFI/WaUQCe/aW
dYIqtTyn1j1vHV5E3td56P2zTk/OgR5Jv7OUoNU0BzFh7E2TXA1TTMlnos7Ozp7W
FyRmfKP5AexVgR1twl4bqYI+XUGgvVkr8TN3SGrMemYGTZGosoIFF3nucMCvAApj
ibZw1EmvNV+LFGWuHZQLciXu3BRcpfqlgaAy56fQ2J3EQ3AKxTuwjgiTHBMbunyR
Gszz14VFFQj66++NaDbZGgkloKaNmRpbRWgBsoAC3E98tbTX9M1SydJIO8xGcu/f
7FUoDESL6nj501TxSUL0kLVARDW/6S85x/oAZ4sa9TJYpGkOo7NGw6wVBb7+7fzC
LM7MjjY6PE5DXc/YBVRNeUaFSgevKWVr3ylqZIYTgiyq+EyQyVjW2Zm/GFlHy0tY
XmZ52lUfaPz1g6Rmcl9WXVVEWuSSb7mKv6NVXRWGO/l0q5iBXgVZisekC4oELA24
yxSjyvaaOrMkOmR5g3RQQs/cZReNseAWL7H4nUoe3dMxglfqxWXXs1jztSteqbr/
akUP43pEkyllflnTqu52r8IDtC0yhOn6wS6TJey0q9Qn0fylQYfqYiymyuSG//Yr
MAxuocgge1uIwxcnN3PDLqUqYLg6CSMr+qqp4yeJ/NiuOM7qQr1Qr5QMiWc9lI8K
RmVYx4aL3fE0IDCDmk5eGsnfeW+OJsVouRD6x+m/sPX1E0rdVEB/bPblahYcte0z
hTfo1o1N3cCSYh7Ly8p+8HlBkP/NOV1NgDs4A2lKYuotg+LhKBrx84OfUjVBs3N2
4FNlQjBQREvmQblEEuBrXbSMOdNnxiX80yXrw+dr6bHmVXKa983Of+/jg74/p7Pj
BkpiKc1VNXDf0uO9xPt8ZOaOw+/5J5sSH+7MENNBiwGO6WvlyuOtK+rEZrnilxbb
8ocTcpaLcgTHuSSOdpoVnT6PFrdAV2a/lgDi0IIIZFAlJkm5HUPXbT1JEKxAh3kz
I1tRvpR608siwaGTZr8xRUgVEEEvAs2ec9GuPUrTUtC7bDmfxfmz0kb89yfuT2DL
eDCdjmf1DaqgPlUYg1dZavg2TXs0t+8cMoM5JJ6d8G7kafhIRGXT7NeBiVmDthUd
jlEcdnu76yp3QuwKQJr0sOoPG14TG3QyQoGnbNagk3KfqFsc7ab3TFOiLLDS7iyD
YHr1N9/qk6LQojXwLrtfcYSJ2irOZz6XzIOAPW7KCKLz9HD9x63EOlCtMcQyIi5W
rWyaxIYGmio9sPO4Qb7B9KZae91ZpBCbFOVzYcPRaJwJY7bNDmH/rHJFIEA4L4/s
xNaxz1vAhigNAhn4Hb4ObhEVipvD5U2Sp8CHf2z0S890Gfdn9ExKnUVI8uE+8pii
FTB4bIW40MlQag3DAYcAVYzRk/sr60Ts5tgAXJtsUGRddtHJQmy0uFA1SIFpWbMe
dYsL/9duzwY7mHTRMcTJ/fh8KWJMrlbBi3mJXnbBVsNflLR/DS5e9WVxFgyDQQYZ
dShw0JkygJL4JNB6YqjL6zCfkx9I0OcRLXD61nNz3HFjbAgYH0zYLTVkN3rNLbeq
tL51UC5pKIxW5RtOYQGjjzf0kydRjhipoHfwtV1rGs54NZwrIv6uWmqlkP5ws6Ub
LMW/t7yJx10JDYcY74VXc0UvALuYDTSTsOLTd7an0AhnbU4xbbSRQQq9E6nANscq
bxyr+FvRJxw/w8o9nnufGJKK16ooN0YvFUMtac9oYa863Lhxg6VscAMQgw9rTJn5
CxMaacDTbvGYwwVlW9RgyzjO7PKjqqrABF3zNkibXeVJ13siuLcsYxWeXNSEdIpM
3CWqM1uBA6Zr7q71Pph5JU11neZcpa6wm5GlfHtp8sBkKM/92S5AwHzxG0AGUqZ6
b3d9ZUow8CJ7u9Bf99fff820IrjABgDNoLevhHjWDHWiD7pLB3g9VBQM4Jq6G8od
Yx5xgrLAjekcdU5jdxk3oXbjUUAACIbJWxx5UwKfKLW3VKwrrLpm0S7ZRL5+4o/z
pQ9xSLc2Ga6sEQLUXR8DeuSv3yMKhQDoZV+X2Sjd7GU0AeeV39fZ+0SK2ZhaP1+m
PqEpJoihjChLWaQZyo3QYs8pmf3qkJhycVKSooQQ1PFON/NxbYZUViDhxwlkVTJ0
x3a9F1Tit26RRbYx9+WTQCX4QhM1vhgDScznnX8KRDSz6KQSgzK8NDvqIm2GjsLZ
PTNs9jHlmOFM+kjA9QJfqxLyMuFoCzag0RZCAdK39+0Qhjz+VgeekWcdZtlsiNzL
g0jYOWm1f7YhK2C0wLNboDzwd2klZg0tW6qyVOrYSSba3fUVyeX730hMEt2ZYv2z
ZUrVkLjIaH/WnSelq9pJjl2zJ2lLSuc6Gw5Pt7o/RsgPvwTeCabE1WQJu9DmKE4J
Wy/GN0ifj7BNCn/2Rzy4SN7j5E0UZzRB9mpWGlvm361pbIp8gr8GNZDTxRahWQhO
8CqQCoMdw+dXYZ3d4yBZDNM7PsFyotm+c0RspCWbAcVYjh5JffqnJ31nDiqYp5pX
vqzsGT2GrtbyASpnc+67d4o8bpl1ojt04OBAc5bBdauU0l4xt30Yy35FUK0iMLhz
VmXsZ6uIF2syGGv4LKKL+Bnc5K1LHeVzsbHzpPmoHwU0TuUTm58wrlHHaG4j1vzK
k0QR681vakMmMUEZpX+gQs0Nw28j8S1WOis9YX0pUDofQwAxHzZ1HS7ga7oEhhN1
qPd+HX+Z3sDk/AkShJAOutaZ+s1jCANcqaUFcZ9EEai6ZwCZPXcSPsswhn4ceg9/
9lS3V/bYvAP6NbvwrHi8rJCF7amKBHvHQoHXSM2oR9o0gRM9tyHtOiRsX1jL51ii
3kX/eiQqcQdWEzxafczC5LuuX6Gzv2XwilT48kK/YIM1t2MpfZJyhS6PEOV9gUUK
5bbaPByOM4Lp1Tiy0FDB9K3mVgKMexoM6ybtgBs4IaktdVOsOqCi51bq5kmxpRd9
dMwxXG5Iw4c1H6grNEPk3iOmBSAwUgoU78iVKdQP9KcmWqz4L5dDhWQM6vh+myiQ
tjUuEdb2YqKRBHTIo71+QlsWGeu5ENWso0Mf0T1URFo4e0rt8C7j51QV8MX9rnmo
y562PH9ifFft0+4W4ctjkMrmETxYiesALfs9/kZB5v7/lc36Bc+UtZZ6NTlbOrKj
pAXZx3a56J1T32espZMoFqIwkFXq9d20ID1EuYUHfVI1MpVv4CRSSHwweGgd8PpE
i4gQwFg5yCLpVMbMf0+coMsW9Xyd29JcG6UTjN95jJkwuejwjhdUdcqklhuh5Dpk
ZFd6cKyoHtkgDh7YpgvU+cpMUx2Lq9vrRhNmpVdW5aKF/wFt0XfPom7XJIu5J6j2
JZ6sdu3rqgMYlqgs+lekADtS0Dc4aa1DqtQebyo8OmrxKNSfkCGk6UJizh7R3jrY
u74JyB6zwD9rhty+6odSW25k6Rzp7pcKWXotQIW7moomnhAO+M/1vyYGgzMbR83t
CfRQ6vzZrgidpHCadNm6BziWHnTlMRiEnBV6nCvoJ0Ej0w6xZ4HSB+fBpQ072T0z
fh33VasOWYS8ixvOBduPFUMxLkwGXeZUWHuLSQX6jKfeH7IQTsGiq4P3QSCMAjRP
Vvj8AVG6mxF6Cbu3WkZW6mPcVGwvr0qU7GK0NiJNvsQdmV/x4yOr+HHiA8QhynGA
0P2f2G4YEhrt5+aW4LTa1ljiacv/BHGISZmT0OzcND7+/3m8tNXuGuEsGhHnBhDt
gwFzvZCQqNMUGw1UF+Gl+yfbt1jHZN5I94pi0uOYmKrf1OgffAsRrRBSkb3UuGpy
qjptGB1rofCpizbsKfUXhmKu8qKCfRniyrF8KCiOBwHnLOFGHkt0F8k0UJ9u+179
HkR0yfvXyEbyCrS93PKv7fbVCP8sd9p2O70KvahsuPLBynCQKDcYjay4SD50Uss8
wi7IpUvQTN39wvXPQ1KgOZQJohZP/g1CqEZDNZ8SAnKhBjLw+hy1hNldpJdkotFW
I9oN2Ivh5HPy6RqGJhyBG+odYTQEUsJvNeasctqr9YI+jTNKTsb6yEdDTAk2i8ev
/MdQ//iD1rmBlxNzP17Cywi9eXcsUQCt+BuU8Shy4ur/4nK6JpNTtznPObL5wR5t
eltUM3NJwzk4+1e+z3H+7E1VE0XappWHhLcAUYDXys0DQgaMk4yFuaoUiQzZkxHi
Jioi9V5vOJD/S7mb9bd6cE0H0CNYH2ifXXojjF9qqtSfj7O9nqIqBCOvVjShS7ay
UgIJAcJi3NBzY5A20q2xqBnJUTLQfgJry4L+CpJlsf+5vb5wncPcWi75Tqg6EAX4
0d3vVuOL8nNvBm2Uyb3wo0pIz3tqxtRm2jTK8+FdaV0bwbQ5s89zOE4pj+C+b6X+
/1CnsIQS9FLrAP7lvTIYqqV1ORUhhpZyn8cGAvAONA9lfwH5tC5tpdmFr5oAiw2H
DTByR+yVSaKUfQ9qUc58axco5mBA/M1PD8N2YvJahVxjhBgx1UB1K/33lm7vd5U3
Nic8xuwU8YkIBWBQzNy/ha0HK4ZolF8KdqrIKep9KwLBI1oBYF3SbrIBjnNhFgmo
TARvUyQanJkOBYq6R/idGo5ZK3PmE1NVOzl5dATn6HpcyKdO7yj08fssQ9mOHpk9
iRMcH8485CZQAYUTdj8bw5l+qUSqS/NJP65emJwE/jMz15Y5MUm29VaV4HS6Clk/
5qKs7qmu25j63jDVIT+/1eyIFeSgEX/8Bxg+twq/wpPQOSnPAJYP2QNsLvtxzzwb
4Bf9wMbW75VVzFYRZhBR+3nlWy7hVC2c5pvRSRucIhS4JZ+3YSr2KmexGE0aROAU
ykxFkanqqwTf7kx0I0XUcY0vD0ZyRpH7oSbyIZTloKRL0XUvat+BOJ3MSqi8m+vL
LZfRoENJiZpVg0Xt220AahUXzbMDCOfe+BGSA8xJfOQjzStmw7pAEMGlqEvNd5+l
/bo667qkJctag6QPSba0F45B/GB0LvBIt2xSr7uf017yYn1BsRGHD7lGv46KTtUx
Y2IANHS3AbVmHRW16toulrpafWGa5+dAbfYiSI+r2uWb3ogGwLHGX0V0QgBHTUuq
AvNOwMBWALhIFBJ+/gQkwyJZotzR7w6hj7tdqfl9Dx4IpqU2ZIxnAVAj/MZ7xTFS
mymswHnNrAxtWnSo4hkqNXQQPJI601iPduWqzIfor686yq1/fZ2ZOUYIWHwy+cFX
7ic+B5qHfA+J7zJm4hO9LuRd9dWpkHex/WQTiLo2i9FHUtcFK5Dfhl6QAV6gjHke
rpdf15MXMRECCXbpg0FRCNyPwMPloVOg3geWXRChxjYfHfnCQuKCZvgeI/hL/Lg3
8jqi+yeSRm6pjtbdfcZPekdG3qcKyJmT4WDAcdjLFMWcR4FTeWs4kds4YQczYASx
ecJu48UXUsgZ2mAGFSMDxRKEPLKW7DO65BSAfN+n8GOBZFrz+G9hj6rukDagLcNE
wY2qgq1xmHwYFcjmuqtSfoTXyd4dPnqIybDcdDJ1PNTOVjtnZptAX0WzXa1ECuHi
QQtHOxF8PzJrwc7+FAKH5A4reTQm/EJ4f2/G6ovgH2t1C1dJdp8ABRUyDMNegr8F
mhqu3nHhn7VcWzL5d8ViEqEHcy0sN/QRS9/dwcfaF2MQBBHZut38yhgyJBHJAZmD
K+yKg7C9TKy1saCAJeTad1jdygUZwbqSMbxDl7oraW5hHhjG7UFlTaVSRYHhOSTm
iJcvBMGb4vL6XFtcn/TC2EaRuHalM1lURRjHX+2bJ0CJREIXAqdDnXRTRYNbaKox
ULvdHusYQHAG+A8Q1wd7Lk2a+VaxtLtIyVvzQJ2aEVN5iT6rhVdqXWWeNKospKpo
BRQzFFVomeGeBkoWHiH1fH/wzkrlIOxtVv+8zS2a3Dtu3ZhLprRbTdcElBWCPZ2V
zrKHuUCiS2hyNT6pTBKtIVftBwjIlKnqiYqDnXvMo8hB/3J98DUvvrF6xMl6Z3sZ
qq9Uk8lbu077QwkXiaWuagIAT6C7MF6HeElijrdnyEWEBCQRHU2u7j4Fz7W4wxWC
/RZY1T2VvSQt2Oa1EwB6H2AA7lDMN3sd5RoJNTMcV9YLsXvBlqye9ClSxhbuXmU5
4bZfguxN18ha7IDsXFPLE0WOrcdMcHCHCDeDWJ/T9hKiSj0OO3wlIHEbwCRR197Z
2FtdVR7GTj3hwaH67FKeftbJkxTQBN52eVWbHZwaB0bdcqqMCn3i/NccWMmmGh0M
OCVM4ux++QyGGO7pn4MDVEOhlFXUdOzrhpTciTonPMco1Sjb036MwQtJSUVYU3Tl
bDpVZWTId4DUvKEwSwC3sIH+xnudR9nIv7gH0zwhI15pq2ym4IJXLi+S5m7py+cA
HzSdx4sY6tcJumXAcDVGnsqxjgBn2TgOhHNx/gv+BqD7cugyThA8iU9s2QNzUGnU
gsjmrEER/T9H0D1kYXwNav6QD08c7kIKrnSMHLc0DSC/JI2uB5RUYGl35WyeKi3B
FXiKXiyHTuwN5Cme/YJPyHK3mwkTW+oAqU0QaEY0wfE07kqilYgjqnR5o+q27CE6
hCg74UYqV/ohRk9wt35bNr7ryX9ooMsCnm3PgOlKtdqO+hwInc05W7BEB7poCnRF
AxtbNjEB2UqewbGZMt5WFiOi+AWDB3uKERJVHCeNva/zH6ITMbMCPi/0LGAyBNKG
VeITY1dcsR43NLkEP3WvSEzgg40XGiFTT6UtVGbJ0+SWqNlPqQ9zG57cLE5iI3jL
pPgtvQtMIAtJ0NW3I05Sw4WAniTXMmT5vscvqxHOhTcD6dkEY57d4EAY2vGyaZMf
jGOHFK1rxrNVm9WtzRsdugyTNlL1MsPj/AgpPAFM6DdWKdCFP46ZcfSyvL+pSFfy
7r+B1Wc/gHUKiUzGY54SfoKZkAaMViBJegIJbt80VhzgfA9+Id1Y8G06i1mK+KYk
RaD7pcpWX4W9LuQX0YT0njmfpBratLusy/6beIQfVujiIxL9eYt7FfewHjnl5ePS
gFx+qlRx/MvBAYkACZ5KcPt744AdAAqs2oQwuHO0nJCBjuuz7qnIX/qhN/S9pn7f
umaR5yxNKLSiF2uTEHVyHPuxVujObyPO5BQEENuzKRjJBfD7vgr0liJnrQy3JjNq
pOPA37HxFoljnZZmejMdIpX29v5ZDesa+9ed5FaukBR6RWJSCqaIui+cOa+YNTHL
UOZ89jyFTLaSczwWnw4rKWHkO0lkZ0XnyKSIX7FwS5Z9v/CUysYr9SyxHugQ8+uN
M1UWTy3sp2kl6O3A7UqxrXOQTnjkcGeC+N4EH4HzDDRwNxBhAzj3EOMRR/ux7CUu
nFzJh+SM+Oy2wxt3upTG2KsZ/HcXSrb4f/1O4x/0eU1xhssP9MT8r1YcnaoGtMOw
2CeZzBvGBZGtHFdaQaFUMrBI0DGU7YAZZiTZg7Ygep+sHWV3tTsg3t5pKKJJcIQz
f9xvRCnuVrB+FbUnpcj9jqk/1eLES3DiNxiRLQBW2dRwq/uMW7S8aPhC2lYM8RPp
E6y2VQYr+OY8hmHA9eD3PGr5uTZpfvvYmFzpzmz7KZ4KzqTewpTc0bE0p9SHo5I0
mCCnoDtXaqor0bok2W8Tw5jijRJSMNgfnvql/wm+1xv150gnJQKv6EB4wnIgwYKi
13aDD/Yk7eREgRQ9KUWejQdQGMCa/TyiE3AyCxc7MkRqFM3cLUxc93X1rc5+gggt
zXHNO6gpflyzRtajWP7eHoSq3FNNTWAELYgq/Vcp/VnJzSi6ozG4qOm0ueVWwpTZ
GABVtss1/iyQ0y/zxRwe27PCPVnGkkKzM6INYXiWEsSjW+aS0KFZQRqfFwgO2eHx
JtQyn1kfu2zp3D/E5Opk6IID5EUkPWFRa5ddEActCOzvynyKzkyqMVboS5urNzuw
hxuKsoc9jc99XHtXZxyZf7TdIMU63QLi9frwed3Cu9QYAXkkKnAsrFW1dTx5h6U4
Gw7emJ+T7ncKB4cXro/n+KogcsMKTW0+rm31751ou8BUpYlo/n3Am5oeoi/JAR5K
/nf1aZNEVQONvrkuKAazH7xtGoqQKeKCRaPcJXlZp9uxyzyS071Q71sfV7wyarIW
dB/2m21CG1uVhel5Pi6OLBlcxMkNmtj5RnuFOqvhHtttZEEgJoQVc3Jdzi/NPOYF
H2jd5CHD3lKFb6TwH0NkjdwFuW9zlkXdSroLgcYoKcJf+eX/d9Oi7spNwQ2oelsl
1ApR1ErjPVpVT9DIaMqVkZ7ZEdYy6HTU9gBYKmF9w/U26xPLqyyQj6zeP5FTgZpD
5lMgpr34m/e+Pq/DysPKC5hDYZoV03WxtbxVIUgohK/hvrTYp6N+0jp+uTbVBXLj
jxwV+J7C4pZydkSN5Q103Mhux+z13jch9MYdBddXStYh2DxWyy5MU/1PtTK6lHWh
1r4nCiZCnGlLCj+puTZTuUxpyCRIxvJm+5uc57kn3yRqh90jYOMIoLdd731Bey43
nJoIfRAcZDyj3+tSiQCDsJU5pYU+hsgmEXLdVxed5SBOeKB+4k9pRDsnZmbKrOOH
bBQS9RzyJ1P5p2zYQObwDPKuXtN+pRAnd4XdCBHy+OYQcoSJ0FZy+336nyPeMLSV
TQ9YBSNteTluDSFpp0XmJHK+o1ocpRg7wZpyzHaSrU9CeDHtAe3YrOzwjjigxjKa
KW6Is4t5CopW3n9FN7g78Kl3JcB68kACe9g8SPHz4Cw843+TDNWuM/L+S8PhNKdk
jvThyyASDrmyf3jcc48drkRbD0AmYwAT91Re5gQFs4pH9xrCMClGhfFuMEtnl3Ff
VdwJXuYzA9DCqs1k/J/hDHUBoU6aQu5NpzII3U9DVF3Cm5m6f+rq1um4I75YMiO5
tgVgfrjYsOK2lmB7I4i/GydRlIZcJ9P80CDKfUYXTUBQZTeuSEhYCOA/fuxJ6KJ/
8loDYb5zvg36xUKWyivxQf4qZY5gj1I5SNdCItf9kitHg9s5sUUFyZWBldPVBMqy
hKGVnVmZWw9Pavec9XKp9iWOaw4SZR0W6fAOz1zkQfLNlKBnRozYdQBWxzY+8hyt
VDQDvlhrnhaWksfqyVz1e2eDjgTLhcay4zAikURsLH8qmw14b9CuuxSJ1hoqdg04
uQQChslbYerlgy2Izohtqzdg1xf8fKfxTvhVpgCeNIRlLk8b4M4Q5tTN8kF1Tovb
ObUEsFzZdqoAzvG9a7tqEhi5xEJd+pgzwOrZPzpE72w8uIXMlh+OkYLT4af3rGqU
XOJAmodkb+U48oou6PBJl7GOwYfldIAlOrUbql7sVE0dsjbVv9wic78jxDOJguxG
POzNtSTYCyQR8JzVOKtcGO7X7dMCI13e6+b9ZRBsrAM7JL1VN63qjOHfcLytWhk4
jocwWIqbBvkWQqQMMEyGmUUhaFe3CIlgxNB2dl6IvL9DkaUjtJGrxBXqb1QKzPLg
tUc5511AMUgnWLhM593xGJIywzH2AFV6TBpJoH1cbXo4mMjwAq3EJ0BX4fgO3qpI
fxvhMUvBZCDaQ4mscBo3PN+gNQKGdgXEZlgrRm6M9Iss+t7hU5fti1JCLTxVj2KF
2VrqRWg9jEBBcUVuwrAgcdbdkKFnu0RvpNFw16Zvtnwmh8iiUjCSPQK8zQ3qS9tX
9arrWEYKcIRJRM6ZocCVWOk+PXJ7NPzI19RVJ0EwwzoCBzRD9skQkVGlhHTYCGXA
dUYYS3+gfzDUuIxatKfEhXNlSK3zOmeLQ617WdeN1fvtCd3SImPuyrdsKr7eI17B
PJVYXIslEgUi4QYyAkO+I8tb3ewdIckVIpqR/7ei71cdeHW5k5Ju/eQRku5i5Ss9
lU2po4UN92WBPelDpEHE9Mmij5tlIf279SzW0qj92hr2zfZbEG8/hpEiEbKFfhZE
WOQEdrGqGQmLNGDsL8PmsOZHi8k+v1cYrSKb2BBiS2+Kqscb3ECJlymJUnZxmbuH
Jp+ZeoemYNrxXyVoobO7duhH0XsckLUg3uP7VbuVm+BK4M9/9veLLtNOe1a6MUBy
57at2TOAgsFlbKKnu+cwBZ/W4FIUnIKAaND+FEuUG/D0iulICZyVR/fdtegMPsdZ
QFbfdDW5L1IR6QGGlnyzNcO49F5ZT3SC2Vm7vdbhxJ9ARU5zqUsThnNEAx62AVgn
YqkeS5PnYGiNG2JbISY3n8E5TSQEv2mIBNkvTUVkFWFd8qwpeMDnTrSoEdaFu8eS
hJ2Wn0sbWj51oSY/HYqwHiN1jXzAPWYE1Fe9ocZ5ww2N0Iw9D5AHetpB/BgBN9Nm
nA2cvFZawC/0Ayh6YTRskPIYEZukMHMW5ZLAiY++8yb1B3gY9UQ4Jo8IQkdH+3vD
uZFg10c/Kw7Osfzu6pwX1/1CBw5sIokbRq8H6T9Rvect28AitvYinlkezEvEAzTd
NJeVBHcxr1QnYivQgKiDuOMCdV3rdm4qHAZ5BMZzEhj2iTvYwXmfZmU/5/Hzaa/M
exCKv3Y28cwJQQ2hC6hTyUPnUdn9t95O9w1WQDKNeQXsmYufjv7/dL+x0E6raWGL
2fLqsM6rOeKWGOliY5hTwatljhksLQZF9Jp+VS7gWrroL+9T133+TH14hrUrrUIr
jc4wQWrlEU7zneMZPf08Y/iuOkFzpgN02EABSeRGkP1I5cE58EWu3Hewfl+rJ5ZS
UcRuALcLI2p38XhQOHPJnbae6XLu04qtepa1PQfSvPrVvJNcdA+llLVAWPm5hW+p
aei5dgxb3uQfNy4D87ggtRNu2K7pg3Je0Q1/hBjXw6G6IXpurMA7CjBe2GDzlvHk
U7vzW5C/fe/XlhYWtXlUP0U64JrIA4SnpwOn6/o0ZCWjQzqDu5OuVKtAUq/7gwew
VpNV09fbp7uA99No+RIjgSVUOw59hAcBrL8F3fj9mJJWMYRiWzAUjmHlgXM9X+JC
riEYybTZatLtV6ktXTlpslqLVzTTY6zgkiwXxHm8fyervPgdlWRzo1ZdePA8/B9N
4GNjGmuv6mgkrUVi95q3Yqiz16rqv45frAGoLixz44SXxNOneG0n0NIuKK3R6J2P
GbfFAmjphgcnJLXc8vmbzVEv8EAylNTEx+Emlj6c+gn9h6jFxoB3vk8fK5+ouWAg
S6MvJgIkkFcFzwyLpnt5SOlE0SM2y6iTUW+LZdEE0N55pq7Ze7fAXZHOi+ZJLikZ
E4h6C7yXKa3g02zmwwfQYwynk/tRao/dtEOWmcKmLTcuNxiPS/ne7f2Wh6iC7qIU
of0kuefHa6Pcs4GdC8PWoGN2qbaS74sbcwbBRNfRSRk+YatWU5WERLGR/z/3Zmig
LcWth9XvCdsWkzU3v/6P8LUDNC22kns20xZLh2z0atnG9KMCMPAgpQvxLFrxjNce
k2S+7LuB43SsEXI9PFHJdw5FAsf9ndmiPg3bixl9yPYrIRD1i+s5sM26xaR0LYG9
VhxuH5ibT8MQdwgwkTPApnrhsCMuIKXg2rftPqOfiLEmYhnjkx5NUmywipdShIeI
ria6D6sw4jSpb8yS1pGG7GRsXqbSJOFEtxkeH5OdfQS+lMFy8fuZqHdz6L6InZZh
HtqiU5RJI6suOsGygkaRMZL9hesjW7WGYLvNptXkyaEw6LfxOf1+n21NbluOKEhp
cVD1LTxM3HBtaCIuBSxbdcsoXuDs4gq8Q98KFi4tRWLj9S7KhkykrbiQFdCRrdSU
ssr595wS0fQpmdz6xtbnHOErVAXIrg0+A2uqvkKSyGuscpI6MXbN2JynIqSFiQGO
li1n8OaCQpwXPBv5Mu/gbVgZhJeMgdtl4UtN5oYWbSknjsfMk9ocxMyC+TSv3V0D
E8c5wNC057A+Ds5CttgwmrCsAqpPXC8o1KyIXO+TrbFzDOw5IK6/xF8JGvqpOaFh
mUKCvD1rK+uFY1sQqcE5TFO1ESz62tSEi/NqXw/fWINrIUdIEBVYYtPdLgNQkRzS
JbiMKgdhAfJs+f6xUJ9ust1gqC/qQ9VY8lQhVf7RqNQnntBKFRUoEoYIvViH6fhk
GMGPznjjMR85XjWRbenwUly74woCTFLI/DUrHm7xOkbXIm/t/HF96unx7zFy4nA7
+84d/3xKcRRZ2APXFyVGAuFMKME2S8FcbXguNUdEpsC1NRjtJ+U+Jg1nXVwi2ZvN
9hkGSS2Xsy6L0p44SAzpQfPmpZJ6K+T1oBDPGnOHmlPB696tKL4f9l04pPQwy7pl
rUFJ/KCjuIycSmwdG+3DxQ0dFTkn7XrWMGEIlfY9JXTPMQvGy+f74F0TfCq04gxJ
i3Yh1AXPsajeMefmmOUou7naiV+Ymvt/Bi+G3BPndYSIreabLHsJBRzWoalt81/4
CJPxsHqLzpa7SePy0rvtlVcv2xOp00S/KXeBl5cHbKKUBZ+Yo8kWSUfrqV0nxQwZ
0VCRJJkggyrIK/9GB148qUlGw9uC1R9280drys4q7TOV8bKbzubfv4a9eYNW+AzO
6CXu49zgvOJnmxqk7mVqwo2xVSMd90xlb9Y7vlmzIDr9f4m0i4GRVTQzhQPKlGBh
g4JY/42Y3Gb7ETGJVu8dBTKoDYF++dxIeJC0YWNeOsB5pCJ58yda0Zc9K+2guxTN
3thJN/jVRBaqPY0nvNgHtJJkNwzI6HthSHnj5nY3IPEzLOOAIuY+/68EBznsYTmG
d2KPU403uk4kU1OH58iKUc8cRSMgQDAxNAWKuMyj/IPWBKvr/Sa49o40RYpEL/CG
0/A+DFL5WNnQ57JGnoA3Tk+4xST17TQZGcLuzzF9orZCci75K2T+a9MGNzuRfVXo
gCJCLgDftQIEd2+YzPCQhQxddLPIbBZLD8ldbrHGznTobbtz9C0kXX3tcVp/BNlw
QozGEXhXJpGcoIf4dMCGUX7k59zgHqT63vZtW2YxBDmy1HvXkZWpA6RXpbETSFi2
vONWsiJWSyXrZWtxvtO0OzkQnaRy/VDr19gMtxLraOblodC6tpID1mRM7jpOGMh7
CNOVeTdHPoxXlm1yqBdsGpow+clAoSWFP+33V+4E3HcvlQhAr39yeh67sQEr9QVh
ZbnerbnXheSgHx4XJL44cvg2lUB2aRzh++jOqTQgj2eVlTYt8DZiEXakny2Z3D7J
NvGK3FLkyzbvx8IdqjAIuVXyUXss+QxlbRf4gSX2o241bHWnVmL+9M8oJ2lUNILG
mlbGXAKCEN+M6BMyWfFiG+jZCGMy6EDa7KOADRnf1LccQQRiJyf9sX0Dwr41pHoy
5OLvvAjwZPKwlskaIJLpGvzB5T68kf/cuVRCpBAQxU0OynKU2G3l/NZbrD9C6Hkz
8NqALe+x2+lDU02klq8kfZFOLtPVHuV0llY1wmPOOpJ0xTBteP/Zqnupk+GSNrTI
3YiQnSvGHHt9XqR4t/Sox249PJ3Ok/ipnURlsZxGl6hFsd4YIu4MkruJmX3M1Jug
28lvcdAq0Bm1mTFFiS2XnTRq2yPoP2FMUa4egeU9ULTM4O39Pv+UmsCY7BgcO5xz
iaMrcYZwQCzKXMAxFaLVK/GnLPqhPuR1NHL4eKirwEk+ojy7gpfpf4lDonca71ZB
byNb38A3I+FNCBDXUjwPUJbH+YC/WHQNCfT8Ge3KM0/24S8cfmKmQUrrvdF18YE0
+Xd+jeyV4jK+bLUCPsTfkV+6kf5OFIwWZxiUWQ8M9/FZWcDyO+o2G6yYJVSSLtUU
H7cfm4L4iSL0C5IG2pGL1J7B7y1T6WBX6Z7GPKEsJgDDIefllNmki5BFUgo+2W7p
mTS9JuzlpA1mXWdjBC5IqwQHo2YbI681gzfb/gXuIa1hwOeFtX6xnCBSQBow5Kyx
OicgATOfJtNLqe/BrwdhJMO7CDqwMpof0rn9h0NXK62cxU52orJHD2h25CWsTqDH
0OGVYLNnyA1OEmBK2aUIrObnnJqSbk3AMGNYFnSonlZEL2xPgC5GujUcAG5erGjW
zgBEBDFaVfTiRVPdL+jvrHmTrp2cPcNIrjOq/G0+QGpHLqUMEgqL0wC8DLyiAgfB
izhvQYtQF+AK7Qgonh2XdXW5+n7sCnVeotfuDAZrf57gz4H24BSv3VKS0vh9Xy/q
As35fjNBUwXsInXUR8zeFGsWtxDKkRSUTKdDrUCWScA71yxmoFSauDSRj1vfIVMg
U5djq17iLyogy26KQ2goL7/DPMENKvKYVFh4ahxKWUR+Y3ScJKlA1GxsWhEeJHPY
eKEmpcoeZM/i5kRNt0Pz5flzKgbqu0EFhb508M8nDEflDCw6nfkjepDPUE/MBVR5
L84rIF+Cwy++IF5QFPsqbXYTRcxcLbhWq2M8wlaaUmG6tH3oJJzv4Gf2Y8lv0IBc
AsrO6F8ac1Tf7cDK6O/2gh187Gftbuv46fK60ycBdf0vWOY1Roa0ReLhsv+DDyiB
yC/CY+rYLbjP7pkGbPh6vYmAAJt53c3BIrJDeB18NaameDquSKfEw83y9AESdnfB
oXB/09wcmnKQjRRYeQATiWuOTmdzM0NRGvBngGcyp70h5tuu8BEfrGl/O85/9V7x
pTu1+ytszkZUcNLj+Pc7gdNtyn3HaBFuq8a1xZRRwf7OsuFBTXd1a/spG41VA1p3
kPy4rIZ1TmOsb7jQy8CGHqi6TUCbeI1lC9Q/7jZzBH04uOso+sbBqjXEnQU4Flat
JW1UfX5mJ1hh6ynbXVN8W7fjXxR/4oHf1xFyp2Od4k6OO2eRxNHa3Sc93F1cR0+A
zfK5KLeoyKADnr8LXcPnG0t2ureLzZWxRalhIY2XlESuzX0eEDGdUBrBiUp1LbrR
SGhk9Zc2MQiU+qYo34rJMMQSCkS+rNGTEMJ4g1ojmqT+XPAsHlYSpQDsJIwEV0La
p/7+qoaGDWxMDKxA24sugBrzqUkRjHLzlrSBY6+XYxTjS+Yq5dGvRF4UtYVEA9qm
0siXQ0R2AIYyGz4BmguEPJKfcMXZ2ALTp6jjbYdGkHhdppy/UD/fPWAtYYcOe2pQ
2GK5H5xqT0dW1lkOgKDMDFvFpfWBzmh9jORa54KRSerkey71zbjmVm3GLxj7pyY7
SUrmzVko6CVzDfQT0ldg2XYoJtE8k+Jk1i+VLjD6F4xDBFEIRpRMx6zfiEalaEMP
zAwf3RH/LHk7X5tjNcREhGXXa8EeRxhu2Ud5BOk7AXMPMKTZa7EXZmYoAnig5YOr
4m2qzCnEVI7wV00RLIg/Vz5UpZ20N5tb124Bj9aq0XRPWpwLJY8gJ5LOYfe7jp2e
mBO7RqEjAgp5LRcIPT3mHsh61KaCcZnLGpVR8X7W2Mf8sjG4/B+z7lRMCoBdabw7
BlEEDS9qvdR9j+rSMSUtLI1nUHbC14AwMMnFv+81u6VSTMIpR/ykzO+3NMJQKWvZ
CP+prTe5hAXXFNQWt6r7/sHrJQlgbf3y52wVsBMrOI4BsT8jskmV7P1NX3TMIAum
oVmptRL/fPBUBczso84At8MbiGBx7f4jp6ZxPVeSOKw3uGFSU+r+RVqJ8gjh5Pyk
mm8JqoYgeN3WYa+gOrtM+jEqWFxbtwGMX4lL26BS+nqacLvq4lpWnBbAprpgYJKw
LNn2bP1z+Zz6B6Faholy5Gq8fG1LeRk/ilZ7ZQ3BWh21z1dbcaTXbj6JaUQ+utor
7pH3j1ekO3q0YyiPJM26/OFQkkKE6eiyfHAOT9V+HAbL+3oO8il6RDSxc1PNTVn1
mtvL0cm9O8ON/rvCt4OHxbQlwnXgPU9VW25v0KW1JflxFSbUQK6hGUiLkVy703r8
XpWyyQiPxtmDaNAmG/cLH+Q/9v0rtAeEISzF4tPWn//wdt90uEE4VK0uKr2XPb1i
8lPCDf+5qsTcOPhS3Kl/C1JSHwUDpB251eoRUqsu9Tk3NJEazBGHJPv+7h2Bp9wA
4JeccnqoWOt8aPHE9LjhUIIUb8iiyzFGx6Fco6qOLfnTXBX+GaZgILwhaAGFTgZV
KjZEa0asUoV2l1ErTNK4Tv/F6ZDdR0Kww8ySWDoFcHrMhvgLr+03frbCIx7RZYcS
XcebDUxwUdVvxeFb1Z4f728hdwrWx8xh2qy1zihVfibVXkvUr6PTglcCqDgvnALm
bRJ8UxLkRTprpkM5eEyDKXM+9PS59oPDN1WGlKoOR6gO8HACj6m0o431EN3CyeMR
lvs5XJRJr4zvqXsLQLXQ4/YhI7wLDmkzuLsWVJFOyRNz95+Wd75RRcJuzXkSHkkL
IgZMIvRRv/CXUgC0k59hqAM/wJBhkEgMI9pLC4KPY9pAhXNl7t2gSH+nm6od8BP4
XOPz0jFnAeuuHJpq1HGZdSTlSNOSjric4tRZ5xSRT+YSO/amZ5NdUUHwOAOy1Yon
pbKdE1u8EHlidgCMrz9Qp2E5WKvpiYidN0M0rnqpGYXXhBL7hJhkmB8mbpEAeuE8
ySgjnr2zFNXmjKTkqniskYjwcpLf9EFVwQiTkmTtnQSYk3GNrY1JBzWlNM5Cu9ar
Tu7dzs5r/5FLJOPslepTPSvP+2Jcm9ypVi3g8qyVi1Sje/fVdc7MQx6civ2L4PEQ
RdjGfyK5Jgmh6zFR11i0ivjmBlu17peUi6R6e9gZnYumKzgSQBmGHIMBXOqR+/r+
O714LggLTMAu71q6Hiqwo+MI95oqPmuOM6s2W0fr6RRc62jY/SZo8zoTJP9M2QMs
GWo/nuu8Hcuwjk+aUyK6sWYw81hTMWnsPol9O/iix2GIOc7pY7V2MVT+ritk2Bj2
HA/Oal1g+kpVuSer+QQGRSgA5EyakC0ggm5gU1IKkfSXR+W+DRz2Zvt+34nUatb6
jajN2zKvcuSfo8MgO4JmEl+Setl95ty5sA9cBxgQr3IZuY1shjD0pVeHzjr1ndX4
YeUY9pFwCqgrAF+NNpK/TQwffq3Wv+ZKbBgAyo8de8a8prOGVpks3MwLSd2P/Ix1
NIudbGn99L7Bh/SMQ/aApqmk0B8WgrkkuuRjBTMpGx1iok3MzmZwi9ESGAPYV1HP
sI2dCJ8QMxfR6TnlaAMM+YQwn2Gb4ef6PimluiHxhkU28WetUcUN2LTDTNo5xsOb
wpqYTVlnPq0ZTpepE4lre8QgDhd9mCNTlAqsaNmXylCSWXJi6WhKRiNn370zcbTV
xpgoBOwVpGLWXVTO2g2Q8EIqY3ZQsRHa/2WIM5dfIuLL7xV1w8zttmyOsqnbT11c
2jQJh6NHtX3Cwr3sJQtrBTt2fwXoC9bSz6+3it/JmezPclXaTNXvnM6+d6t9cwyF
`pragma protect end_protected
