// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:15 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
CVRTP+9tCvnzeMetqxzOmRaVEM6vi36Gygp9zEdcXVk68jH6RUyP9wEsYrijFRp0
tHuk8VFfNeENcavfC7g0N29BL5Pkw1TlHKhDapyHpaVPl1sl3iviP6fuCUaO8Jls
jOV0CV4psSaLaf36Vn6Kby0PPDScGRTrSpxMsh9UcH0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 23760)
esOUUdPu928ejhW0qt5Gw4qfQ8TT/tcLrutNqp2YNnQd3ivlCgF8gSpVbwXZ4PtJ
h0YQGt5lO89rlCfK9qT+DvUyj+dpexWDJRbm7tGWohxLMHYMSWoFRpKxAAnf9jaU
yb4R4qBRJ+Tbq8tdWcBJ9+cYYTFVkamznQpOsRj7a9KJjecjKUuEN0QZPVx8BE5J
4ld+at8BZ7sZ2ERDd1JhK34KqhvGQW9Oj85LVdizuftcTESg/1YJaGAYDc8R0jxR
6se2OommgubrykvCRMo7wwzxTBEQojvIJ8b6UzGRS3ozM9wl2IZZtQiPMVOQI+w0
Ad1adbGfPnoUm1c06qabfgLqCnKnE3XLav99VbUDhI8tUd/tGwXSN5eEn1/ZaGdL
hRUbPrf6zzLawCP1qnnYeFcFckhjYwrtf0l9rp0BmlBEwA6qHN0gU12GQ+YVGqyL
G27sc+605ZvtiBTNDEfly86sPfmv8twiuR0TziCpL7BgmgmXBU0/OjdPs0JUmhfX
V64gQ15b5HFrjZjIiBOSCagjvHb5agylvGhKxjt1ke7REowUP02C2wrxXUoMrJ7F
VF3xYBuiAWsSAt63Juxy5SNccMl7Q0BsUgLFm4dDqJVxJ3zL1GxTXrM7iJB2R7tp
nwFqHaqaFnn57NsH8jzAM2YYddMBDhL8yuCpf4FOyF4QmUKnLKOcuHCVZwo37AZm
Q45PsTvDWj64lgoB6EhQwi6eV1ROoiIrlajhnl2g+7HmNIxhT6NoOhIG1WMT+d1g
IlJlrhwWR7kIPF1nYcKH+mXuW2YNejz6V5925n0kDQY3BXhT+uFe7r9awW/eGW33
7QyHhj+idTgBRexD+wQDikltiJI/dL+Ei/XERM388ZdwhqN2D9Pf9j6+BTfq7YkK
qFQVbDmHr9u3H/d4mc1Ij13O8EPsJJ6bsnjriGaM/ZzHElEGEYgdywihRCjbvW88
tR4TMt7LUnYNKRISaAw7wQO3+9KWWV2aCdtnnkY8YtPX7/1F3hQi6Sf1/+G3Q21N
tS5+hq6cpwQXIvpi4LeiC4C0g4p+jc+ZLFjJMBEen83WGjlmEjBXqjcewnvGrqnb
VmB4hVFZwePdN7/sGWo5/MztSqaF3cyMWloTi4jWvjsHn96BIdC7fk7rPM9qTR0k
bghqjvoQzEON4cIYZ34JYdL+lxEQ8vFoE69bhhIMw56MCCKiQUYvlRimhonIpVBy
GOeCQ1wKJSYJrquAjMmIIKtGOU6pdGkvUXDb4orr3cRhQNqcp0DvF2qU9096UDRy
+Su8xjG2VpRc0nysv89cli0c/cccr+5KZAHx6uVyaWgDmC29E6cxBb5XYzlROMyW
7UaoGIQmtI1W423eOIzmbUF2fkvu80QwsKh2nFrPsHE+CNx3cF3w34AYP3CCxTm2
97TGltftca1cOcFsw4ram23co7MA05VNeA4DP5JjQ75XOZeRUdIyv717cp47s+Bc
tQgceMBgnlX0O0s38yLx4tzOrhVCNjqyP9gpHIbqNDEcvEykP9Xrrp/F5D0zAom0
/I47d13Fb1DrvZtFZusPbvRVqBlgwVea48YQAWoBIH8BdxMlwpQHDbp741rmdbhm
ep/C36S5KR9AiP2IYkyNJMiglAqnJLXdWMXFnY4cMu9CPkP9qWiJn+8U+uV4G0/i
+6l31ZjGvOjIp9B4unkLxOFYZG4s0Ezp5D7JJmFgqMQzSiQt6nmOHmExuAbKxAx2
GPVIBFmLndPXBwVc2bzNziEBex1Xs6Yd3eTyCAWy0Bcy8f2IBkys8GTXPcZdhHTT
bB8vTt9oqLBIURf5ek8IDNQUfaXNY8Ea9gPuL6GEvWr73FhM5ohVs4gxCpwaJWGX
uj1gjeY/InDhkBqlG2J3Op6bJFLVh3CBC2B2eLWtcroNjjDs02z44eFudEvoKzHF
onajxMhkoc4DTq2yYkNm8KOZc4EgzXVPwv0nStHDqb9c0yGD8L4RMpqLOuXM8tBN
4OIp9/shK7kRVA/TVCBdYCZnWiBQkgZpgHxrxtbrkbzEEDiZGQ4CX5qPsCeTvM+J
F1Hgc392n1mbxhKccZ5F6UxojmFl+oTOIS6zpoWAex0GcblWQnt6Y1mRIvhwqZar
eEOQ2kbuuUzUCbJhbSgSWADk3KhwNEDzpW8C2FZVSTsN+D8ld7OR57XrdRR2ZfDd
0AttkT5j+81GbhjDhQ7vV6YXuwJ2YbHfhKGJzx3s0LtxocrLHnfyLq+UGCj6dRB4
iHuuP3xGlMBuTIjHxAz7rfW//vrvFV2kk34aE/K0LNPnVTXg5ZaCFrANjNlw6ZGg
t9Z2jQP+OrhEWsqfNghtIAYUXEAdI8tBI0pISWpsNvk/emwHHaHlletJgGsP4sqk
goAMKtg3lpQwq8X5fK8cePIWIkR8ij/ua18bPDY04PQr6YUix/N3jiWrEDNlSi5v
jfMEEKBx0G4uCAfTISPOYJNEWA02Jb17ieoimjC1UQxq6hXEqWOYXoW6V6Jsqfg3
CxvDlTa2XttbOls4L7pzm4Y49UiQGWpb7IIWcZMvAgsYxg70hjvMdMLi27uVIIlJ
nSMrFGUyv5y/Op77JmSfFsUpDX+Grq5/dndY2yVmJ6gXGjgBtwXstL/mmyvcerqH
qye6FuxBV51rPJwa9k5aXe+r4i/1j6jGDjtSWMd3pDFWAHHCkIS4S+cMRczC5Xh1
Shg3TJyRFWRI/qOrBF6Gc1XjBTRdHvh+d3WkTGn3ZQePlYiHcpEUDHtq/Ee7eakS
/4TJZOXB/r+5CZYR70/N/DMZOhh+fTksjSdXhzAM4I1RKpDjS/Ifq6+7qEBBPu2H
egxJ2lGLRWsZShYF08dgvucA7Be8+ssZk+bVxtgX0/uNcBiGRgH2JmFOV2iiwyfp
RSwoNW2upeERJvJJpdar1cIIDdV6BPQkkHjYBbMFWbOS2zwTnldIp563hCcBnluh
J7h/dUSjInRMjElQdAW4VWrO79wLIwuqdhYEKkSY1SermbrkNh2XceKcL2a7hmyf
8AvbHYocB5+PKGjo/u/BKJAb5NIByuVK6MCQjxOVgi8swt70EcNyGxppqGl1x0NN
3dHTq+RbaRjsnGfGaYdaEZz57SUDOQfXed59x5nzVQ+ZpLpA3gfxsZ2r9hn/BS/z
Ds7xUvUankF4B0wbTGGaUjk+QMFWfx2OhGGx++qwfGvZW5so/p1KDO8GNJudQPVr
NoaIQ6FsltnCKlKVGhfEwK0xbYAsDREiXIn+zVAX+hd4u7O8wSoZ3OBrCdlqwReB
722RRwexba2wdSjdvkdMKcP1VaDv1D1gty5WTDMOVKhaKYxC18K7J5dqfqn0pt3j
E5Wr4mXHxlMiVOjA1RYiCAks+6sBy5ekN4d3C/03FhC7kNCH7ZuuqBPfHFClOIsu
uX1cOX1BC3jSI8cfZ2io4Z4oyuULsjEY/fhXyjCbdncfyBl3drT2OpGrdnY6p4fl
mNF8A6IGb6wUpMUDZQUnFuH642nkYL9xM4EzSWo5WpBalzaexDlJy6HKDhYqRtdP
lldSkWAD8bpZwrr9rcGHUQLV0o4vK0lYwKbu/rEozACKc+KGXZt9jtrzxztMuWU6
Dd1MPGUdQuq1hRIcElK2LMX/bNkTECLLmBOY3It+lsDAkCDrbsztxRKneEJ7LuI/
apxqGyNsnXdJrC3iUDiC1gsCJ62LgMxUVJz8EIaCvZYYVqkPbGx3C+MZ6R6Dcx/G
UnucOfsEr59jMLDca49GwKgndsHD+w8dWOYce9zHJi47gpUCs9Inw55AyUL2LIyc
aIfQyjFOxhEQm3EgPTGK7yvnAkUDS2+Su/fOLFQ/DFoq+S74ardarGLCB95OiuQq
2lK819Exvh5cp8tF6wjMFz0NnyT0fRaX8ufd2o6x+sUtbhSbLwVBnJbrUBAQk+kl
L1jD2650dxsQpA/ItuTa8C9GHcIF5Rwx1Dsy5Vs+LDgITGC24cDcTz8rvhWRCt2B
0HOideyaCF6NRKj7C9LXV9VPou+prsY7Eq/B/AbeZQ3JhTTTH1QK2aIs9YL4PkAA
ioHblzurIn5Ans7tEqgz4NQGUPBSi/9PIwJXg8i9QQfCsZvKAlr87mlGQnJGT6op
8SqQMrdRqENy3jHZdpJN+RQwexwTa++jTIb0IcFDGP6Ouas9KyU/U/pUUxQ2yrA8
0vN5lHNs1gMJ1QpBUy28a9rEdKbbW4yR71Tyo5B8OT7wvmdBNp7kGQiur5gR+Mcv
Ar7yf1vQaiJDHCcc0c87vynuED9wNW/+JcO1JELcXyNjV+HpzF2JiqMvSekKGZTK
hxA1vBOM8ZFflIiBUe4wKnbrbfPzLnH8ngZUxMnXMM/GQQF8IWSnTEVWVUZoYxk0
D+xPk7U/VYw1M/IyJr9+n/cUJLJkqczSPQIyftP1jYNyX8IAB3XkxoD3rY5M7oRx
QBNiRvC1mYN5u/PESz+RakE/xOojXBSv/sVhLuxrJu019ZgiTgsU4jzbhQtDsre3
CYCWVb1eDZjPD32/+4qijf2QVp6EDi03UgBB0jXI1fd6ThKSFGFTFURsD2ft4qLr
Eom1eCb/rL0EcSejS1TW+TErfoX5emu/TL/L4JVDaLqx0JtkLceMhkGDP7P5rtVv
I5j7EP+3SIBIabkv4UCAj7X6clgpYngqKWvblirxRAwuiPclazgYCRA41EueAU9u
xsXn/RiZW0eUOqYAIfsbeSiznMvsPbCz3lJwzWBKBIXtRO2+ORiic8LmzUrWr9DN
7+/io7BiPoRCJH2ldL/9hzTPs9xlwejl2bWN7RnVlCZgmqozh80u5MJVdAbnVQw0
+qx/dtpR+t6uEasIp10oKymX2voQrzcvzgE4qYM6DWP/YTP1zVz4EpVFMH/msNFs
/PN4QpcQcEYUUbdZw2D6ASc1T8es0Su+gtoc8DpSSpx17+fTNdZj1IxteRXOAidY
DW0an0z2nadHgCXsbAz/Tn8Gogpt54FHM5aG+1J8PUFAjL72Wwu3WRJJATlCnK5Z
tWE/ydHzxfmtV7i4HONLuympLQe2jKhyxZtHiRqClnk6Tw8SA0D4JfXC7CCqN//K
nTut8rfPehfCdspHII3ZfSDF1OwO9oJLpeT0Rb3kP0mTtQwVnYwo5Aw4oEh01D1m
pduMMXDVfNu2aOARF8/UT45M1KwqiRx1Ggd4r+8ABKtdw5SbtWpevKOjr7IXEMB4
fDxzKF8yFiPMVfAMO5IgqUnN/dfEl/8WY2CFWzuqGpHX9ca14r5N7pvvY4i9jvIl
KqQljmtIe074y9oyb/nlm6Xlki1NS+2ECZ0J0SiWq1Us5uPtxzLyeybZaYN0VJin
rzv9XJytl5bnv8gxCjv9CYeHrLs570YAfoMLAiwEnPbEgqxGiSx2WdOlqEY89HQN
/VVzDPlQ//+QynzLcrMsuyfH2hArfR8aInpA/waBh0RcNNRQf+DkpBbvUfYMtKdM
IeBL/pGzWge2eh3UMBS3sXUPMLbTeuGHt7TJi3CjutJztW3Xyn3bJSS1uctCO7M/
tWu27MF58EtdtLLooiXPTiT9C41ZZTWu+7fwitgHlhS0SS5Qyh4o7T4gnhIp3K1I
EhGwogBjz5CUzzNw8Wh2u4/YD/iMKF2/cQbTQJoYTueRoCqT4dg7A/4cNfUpQPBd
j1o2uOTCiduVea1Ia7gQoAw7QbX66PiAkj+HwDnABetshoYUTpFnrkiUA8VhBqZt
3aJToMJfGygkuCfTC3z9wyBOerxPdFcSbh6IW4yWfPKurpLzUu9qub5UI7RiQWHR
V1IEqiAYI6VWU3kM7XxIZetspdBxeSrvVnA0W6OuwU6XRxuVbYF/K2ofAFREMHic
YDVM6pmIWhgAPEAj6OshfnW0DEMz9pz3R++uoU2GkB48VuX+GCrkWMN3Wfu8yQQ9
GENBoOa/gd7m4slQwzcN5NELkFAoo5JdokLRZy5MoxG9IxT8s9hnMm/vGajHeHhh
7I/Zz9R+D4UPSXxlUYcSyGGeisrxbxKYAe/nIH1lsdkQImHqfs+ZkvxkhFne1L/h
0AvdOJOrL3+ATNRNrXdUrW517vy6VfokgFNPzlyUvB1t+Bbb+CCTfy57K1tv8/fj
vgC5UYUj3O8Q7QRZWS8ToTGAaSKsUvJq/GEqqny876vMLsdCYyz9g3B/H40CNEAQ
ruAoEkgRU96g7sTsoiNly5e6FUNN7NNaRuglFVismtoKq0Qk57ikdvCa4RCRF/Dd
oeBm4D0SaamMxamcP5CsjNok9i8L923qFLni4+2PdZtg5CGq+qGkUXYH8oD5U/GK
VsuCB95Y2Id6gzLlxIAGcMd9bRDYRkicNxX3JJs+BlMjMhvvCvmrU4iTX4DGObIH
h2EU0cQzU6wxz0hgWFn6Q3fPVtWRN1n4rYXEmql22KI3ZMebBqzEEfiPZf6gMARJ
wSkX87/14anWBPJPz7gISFyDjVsJkheTKrribVziXkR9q9XJnxcyRq+NtGkDXElq
2U3iRzVAH3Y6R1oYfoyHuR2pJGpSdldqNtUFXgFhAnhSmUL9ax3Z0r2sbzQpBrFY
MlRMa5cJN00A/k8egKH2MPK9Ttedq5SBjSGuR8ysz5+KBbvbS9TQt6qLh25K+xu1
UbXXhuH5CXr9aFhvq4ZoNNBdJnBa0/neTbuiyi8wbi+liUuAzjVq4M6jkXXjTDCG
MRsNtXOx2Zr0F4KIb1tA5XXhsrKRfec3SDEyirXES7x4+NUtweIapKu/8Sj7cb8L
z4iTc8PGnz/jkyzu4SYtXLd9M0NtAuCGYU9G3koHxGKJnuvUpH33M/ytFdJNDSXj
JW3k2dKNrdzQIQyxnHiXxcv7ypU04BNxvnRhm68XqOKqTCO48+CMylxKbKry4dc1
nuVSmDNxAJHyzWd3oa+aEox6C93HQ9DXzEsD/g8CPsaXyryozNvd+f8XJmHRFGRq
YIw/JJSIzsbhdODGRq3PIV4xX9C3Y56lqPvbHW/As7zLllAzr6kmRMGNnTAYzENs
TTqt/t3kTBwShGtu+jVezbCxiMfiACokkSR/7Oy2qjuTmC39D1Yd31pMqgCVceiI
hdBCZvF0aW68WdcCilCeZ6UxQgeMaYesIaS6ounJnIZ9++2r0ajPgSrO0SYeN37E
wQZmw9a2CvYAHV0N5NpuYfvSwaTUxO+yKADfQm9N5aawO4lRN38O4Ib4qH67xli0
eEOwb/E24PnDHaD0Tv5+WMb5Z/6kzQaJX/je0DGTOQ+m5HdEt+7tjlmtnyRVcmMo
4xC2fBSY0B3iTXKvDCtY9kYkfEXqedOWq6vob7ZgtJ1Kz648Athesn74g62zguIg
l3fdFttw1N/0sZNeikmY0mKHYkBjp8ULAoN7le7Tnc+rXfA5O5Fl9RIklGL5re/e
2SM+nQG5xA3/NwMTxUJI31fBut18MAvySlYi5GOS0bs61Z225KCQFAyH071f8fXt
iF5gByZ4dm8ihnd20bddhoWKGUmzLCqSksNzeeFVe7tkyVcCGrFbArhqZHnbCNHj
wlM80i/JYQnNUkU6YiZidn2Vx96UuOStJ2F8UzZh47qpn/Z9jJrWoFklG1shNpHj
tVeOF+lj9pGigkjfdRxBVJsjAE+xIF1GNFX6+kPF//ViVc6Jgy99Jm4vcPHWWlXg
9vTu/VPOllktHX5g9zgEEcFm8drpVCt6S6+RPPCeaI/y+upzbnHNdXOMMiREqx8E
NKdEXc+KSmE1XEw0YtGZC6o5/jwT2mT9GSZArTx/ucTozbv2A85L/8nHA8wqn9a0
mtoAFWjEnR3rbjIttkIgGzV6sfXKRkpjvjMlLsva9u5vrZpmgQSKA4ph25nzuZcc
xfO88YXDPnZddQ1qtnxD7aYb3Ub1u2BPgq3yUiuJ0756PiqhYXH9iLmVT9d+rqXO
bERIJhk2Er7aeCVyTHZo8Iido5V6lpY3tXP2dAfOYg3X0rKxtq48kxvxx5Eph6Ia
AvBAaS+VGjbbMN0CFzvs9/EjoSKiTsixhxapMVPkGQAvl1SIkIBoR/up2gwbCpb/
6CQ999TUQ+wiAp1wAtQN94mMqca25iWD0xqdX2delCSaHyn9gwf1rfRvdnZ9FEtB
3I+Q4DiznuIE+j5SeoS9AR53gC6y53Mf7nCyWuVGUSipZ+vGmHzV14WnkmCBktB6
rChpA7Q8f0+qYHNx2yKa76ktPnVWHR6rzOaiDVom/lRe/11E3Di9Qp/2yvwgsvYI
vLpW9Hnhv0twB36INgiL0XUtduAm09Ku+Jr+28lharyMZ7+wMvs02ccLC2lcnRh7
Ntr2IrAtkwHpJ8t7EGUw9n8GsO/GxO4bic+UKmo9WpFdKJirrE5SsdV4AZJYoJbc
TSOFljVPEOgPIIxO1QwxVvTbaLLzwSjZ5O2Uehq7yQh0dCL0dgB/paq1bRLTbP2W
+WEsCLTK4NaatcwOd2uQnucAAqzcPcvdrn+su2BCW0Te+bxFnC67RNW/x2bk8OdQ
grE9hxdrmyPriCE/ucyxfTvHCaaP/x0Z9oLijuINByqaqvSHSZ/UIlgB8dRxfM2N
ffI7Fx7K78CQmu+reFnSum3k3YK9QE3OWyrhS54UuuNWGlV6k3sMVEefPxFJ+ozD
tOzCFlE0QdVUsd16X6+nNp3kQpgykfj8Q9SpDUDKfg+ABbeYBRR17QJjParlFdea
tlpvGeLFn4tlpce7Eqdq6ywLzzdBEPAFONxx5cG+VA86jIYwaiQOjAMGhGtfrWDb
aHIzrulY5JgJ6ILCF5+5h0tjT9CbFaYIR0w5NbfR4r6ySONLMPOKop3pEtp/Wr83
eJhaNx+w01OSETQ4dlPv/NUaTPB1yp1h7E1H3nCpZqflrfJMKJMuBe/vlMUMjdgV
SJEMNiE7D447PYb4PLRkr3cfl5nJUcr+HJTxJTax/z4SzBYV0vGJGu+iFjoEBc8Y
IlZ6vFHRMNYQRWHE96ndfE1M1EXqOOUaljZwUCUwHsxcy8c4v0GyazOMen4EtnJC
w1TwQ/old96lnYGS903OLnYYyw6GXNS5mfAgPP4xAuhwz/8sb8XnyE3MHDhZqFyz
go08szfMT25xzTiBH2wJ2j6TbLA7kq3un5+chMUriIAQc3VI+trZGCOrocHbO5g3
P/iTz38oLjNnkSgpbjO+6P4PA8CbLd5fHDJiJtLbkVo+pGMQHlM3VyVJAMta8AOJ
v+63AG0EJBfYdXYvy0zdzz6fZ1H536eH41/uddzVnKQbCg6wgLREdcJvBWbL71Pb
PQ8/fkzOpzjytwAXcZxDmZe5eyemxml885BkOkDK6yS2B0dS6dv1e/RTb8GKYbwG
Vc2rqoS9+u5mVsHQS7T76kt7JekxclESu3F7V9Ymsrb/Ln+60g1PPBT7iWER9GzM
6LLG4n9UM5YXUGJV3TBpLP8bb6fFSxTg3xIfs88HwQTdAapXuHPFKh5zmcOWFZBp
5zG6r3z51Q4g1bN5EuqQCZ922yB/nBXGMlKF7QRwe86SuzNf+tvuXeeBfb7q2HOM
FKDj8qqFh3w41XsgQ5E+6GvzLIA3t7kFJ/Q6E7eT+xszvp3tYeTEq8yCVextvl9t
lKCxBYFWn34avL2WsHWByCsfr1IxMLzeoxiMED4FBSEVaX4bS9o9GSu8J4Hy81wS
1IvRxgT8549MZgRe/xSaQUZvaGZ/waEIwosMMJCJYgxU5JM2IB3Tsuz7vM8xBdO7
Xs8Kn++i4cNQsnKnzi+61KsB8INwHORvuh/Jgwrn02DFih1RquLb3jrxp7mTM8Yy
3YcroDRzpvVK98lyYj5PR6bFUK8gflfTWZ+ECh059O+w5FsWtCIRYjA5lEhos0TM
Ghpddo3GyvNc87VTYGs+3MQneGbo/Hjim/ID6AmrjbKFdlUX/Ede+VvG1+PGlHz+
CyrxrJb/1ydwJbJMXYNFUt4eSgLQGjXbQwqH8t4wJamuYnP3lBzKQEY+H5xXiNaF
1HkUjgaenAxv9SbcbvwmwLZDuzQzhUGitwFw4VOB8pAv5iceLy6d0oD5qnDf4XCZ
roq+nVJ2GNfjF4jkcyFfxQFBP32lOTGSbBmzOWdNHoHti8eofgEZ1vN2MGbPLmSf
ZyMZsuRLqNCyCnpu75ZF7iNYLj4PUrctXm4KmnvYNUAuoBlj6h0PFt8Ri57UHwtC
RbjdTvBOUbTnmkDboeB3HEcWpFt/HsQHlCuB4n2KuVE4CdwAJXVUKx6iY9kG0lHY
6O9Ucsk9cJKuasy6cgdOAcNZioW0Y3Itjb4Ll5w4Cd2BtJGKI+U19hypYciFKL1Q
5bzV/6No9UeOoB5y8+cOLDBQE9kdDpF+z/xsIWFqUuzyz5+z/b8CJv1na43QlsF4
qrooHMfHNLqzfFyOb9ss0wxnzo+qbvVndsL/C3BcZ9DfdcOidDAid9ypPz+uoUVF
3mi1U6dC0phX8HzIkqZMRqhWl1BqIEeMYPc5oiY+LptRA1Nc/0og9/dwXxz4E5tG
wWIx8v00EpfKvAY8hBEu6PZDI08IEXOgCDDZxKTc/DxbeAm80xYRCN76lxqmnY0S
pgHDx0KJMNKFXGfvHoPKRltA4RBScan5vyHYMM42IpN2aj2OLkLicwS1ZTJhR0Dv
b0wBpD/m93q9ALZMWRu54NlWgln6PcAXbzzB2FOPJhfYKNMJdqRFUlZHSCtZBeKO
SL6JO0eoK2p4TZRhQxfgu4kiCOupWIsJzcBwhhJTcHuD2yxtZGj7SbI2M6s4xFHM
c/SQ/AxcpsroPjvDvyiNrKYve7K4lf3F+F+CQK5WJHt/+BYBbBa2opYxMcwfbfqL
Y5Cu1eoxCWm93kicwspsRKm41nuiPdy/7zFLTnaJjAMTGcr1cyhUZIcjkFNDhD78
if2i6P9STsOItDswcowsbkFzQuIEGc8KRzuKY9vltqpTyJaWTJX1CmvY/HA7xOop
V4JIdE2gqxiJxD192GP5hqUDytRk+73OJ0fnczzldbqCmvG7f83KG/NgqskSh7aT
P0AeyFERF6SSwzAKBJp2vS5wu8Ih5o8FoVE8OXpwcWFCGzW78S7mnTZpGkV8955r
SVf38KTFQUONfr6aU0Bu4kvHM1lWGwUkzp2nM8n1fCZmQtwKSZcxIgDmK4wh8nw2
TTVjbRjDNNI5i3VS+aUPuuxFPyaxNjGT6FJevKJlWBUrXnIgsOKPnN5Fd2uSaP8+
Gk8aZyaUA/1WoQzJKIv7Z61PJxVbtKB0R/LFo0mhN4lD3gCF2dEQAtOXVurHirlP
fc0qy5sdWWSFjIrMy/EA8xtluOLlxFMevCOyH//WEQkH54u/WH3HyZLhJZKBBBco
Y9XTYfICfzmZxDMzcltqAX0hbOZenaO0WmLbkVqveW61ndLyZEHfZft6AxQijmhZ
NI4qQByZc7qXxf27teQsDBo7/M6eeINLPpJZork/8zUOd5yO5HU/HGTa92iQtMhb
X2QWm9MukrAZhPZVrtx4w8z/k+s3fFa6kXem8ovuo4Db1pO4IMkasF9BW1IREwnU
Lmi04GVbiWMy3/BQ0siXB/tx1x/r+G0HOvN2YZ9nIMrgxAO2jQfb1Vob6VOXzWw3
gLaC3PzC25jUBogmuug+OL/QgYPBDt0do/QgMzJozkkVXWi9kGR4AvJWeycghMrN
7j87/CGJ/pW7pZ2dH5cb1b//uPdyktuPaDEMxWK1qA9Bm24VJ3Ebhq+cGJzNlLSh
+nZMQn13pJ6VbGWp17tMMZ2gS/hsj1MkTujwYi0dkFPEgc6+0WnVolJKP3A9TpVb
UOZNo/KgQh9JmgcFGf8ROJkuzbsMB3KUu9mfoD3mVcPhhirdRb3QHYNlJICYWyrz
iRsmFlRMbTymyWueR5OnH6RzA2tm2OBogO0+qJpyUCK2m18KnRNNYLb3+nYnUieh
JFMa9YM25mNwXWp0GSF076UzEWxnS6cJRZ8FwxZIw+hBlluJYbbReLPY7MCRKOWh
hUj1eMT+/AcoTKlWBm4WSOq5hqaQVydmDfTZP5SSOYZbCXdzWtFgqi5nkZMGF5W9
VsmdJPZn5s7ywZ6WvPliVrPXa2+IJnczwL/SYCnZmWGvynqCbuyygVUqrjX8QQU4
1tg1+BS6f790av2jA9WMeqhyBEo55TB+MByi56CLYduJHHjFM3WHgY4PjSdjDFJ+
IOiT+cyx1OfGgbJFzurJMqETZp8Y4WcY/A6MskCc17bxLI64pIZRMRrLuHGkNa/9
YeiGPWfRtsHQ8w2lVrS0tUlQKogsmjHd9r7s7n9VSyrU68VBDJRmPOA1rfkB6r1O
4ZJCXHOP+faIgVJmGblkEAPKolirYl3UZJnNf4d8lT+vczNwlO/q+RG0S6LHoNnj
DPessGq9P4zHh1cIqVKsBzrKeja5NgzCZrE1EpnuvHCrO2/OUOGaNVIs3Vulhe/h
uVMQtbx+6OxgAXjsjn7nNM1w9P8LOi7i+4AIPCvKdZ7KS2xEENAT4TUGYMb9e7KA
RbQE+qfSxDGxHk2MqeD1kgXy3mxZ119AHfDN2+uv07fsxtxMUiIp3D693m5LbYov
xMVb5mJoLZ98VOXGEIIpxGfH84cKXt+18mMjmRcjh6FUM0rs+DqbEO1+OUYTH8Aw
UmMsfPu9b76nGIh8bZOmviXkkHeVDQhnjLsV4+9lcW2sTyPYFF5QBNUl1YSVP1y0
pqBi/f7S1NBSx39GsVRqklpMA3DoUjmI9er6nahZAdOAOL74cLHTHW50S10vn1+b
vBjkyhJdGyWaKRuuJrM8eKrDdDm8OFOPisUfmNKxjMCHlCUPjrwv7GnCb8ElH1ix
CwWx646xKzBKXVzaaSUJhXRpTHk3Cor5BmbCmhX7WZFNqig0/Ng0LshO65bwTp5I
xmyOE7FleVtPHUdhucxUfRwaPaedYsings5o/RzT+MJ4DX6D9zpq3VqpI+HkjGL4
RxgEJEsFBYqhK4Ec+yVD4Il0s9BP2Mq6lC3/qe4Gv+DibMdhc8/uqRna0WWRbz1H
8vv0g22M7PeN+RiPL+sazBufoeLKj8dgxhamCgAhu8XPTtQKOFxueJGvJBNhlTiS
qkwoesYr4yxvisRDutnI4AEfE3TNPLBEkKJdma+J+EDN1MbK367Gk6NqBf+3xHic
7FQbYi7GgdPN5uSiPehjS3GPiDAQMCX5zBfAqalUdYjcX+p5mjmsj1pGmPp5eZCI
C9n5YJE8CNCx2sqyIpbOAnb4i8eD96OM2BPzoEmdjnyTYMNSWgBpbivVI6L8CoIi
kAWEYzL7ZLZA+1DoGB/RdvwvMwF7ChaWV+eKmXvBehIb60appd5Byx7ObNLzbXfa
mkCO3Vf6w56GLI9cpvKVIpBePsmo4gZ0+qvAyQI2v6wZbtTS49npqsnydyEVkVaX
sG0W1VuUj+wXzY8WfzfMVW/NE2CNuWM0PMeGyl5k5H0ecQWoZH2fFF5TaN6vbDOW
PmHjmMveBBincVFeMgSz4o76ncW4kQp4W2N/DNSY7wz8KSCrYRHqtkUphvR4l80D
PsKhcMgp2dqU+o7NntSfjmqTPft+PEyzxlcu0dt5n6Cs4KIkd1GXhLhL2zXLSI2o
QwmMD2o5FbGyhMDBoPBBXqZu8+TNoyvKcP0cZHRKvynb/ErIls022fHTzJLIjTvT
Tg8WeziFJlbzZZ7Qx1TemLgzhenqt7+xXOGlJSOB/wnGlRjWApIkzyXribsob5fv
r09i/woIdlsJFuk5gzn1DZwFUb4LAkeTkV3+EQcheFTAmXBZKJtLPCPXGy2+LxyC
S2m878teCT/yN9frARVh3h2YMHI9KwGLFTJuvO9aih9nYbkajV60CbCQ36vSIXEu
b7OdEPni/dJR70egQwke37Oy/uTR7eknc179pR+RBonmBT8tGKPDQNvmvAAJbk0G
jGLtL6edYL3BZ4pPT9MSfYfkq6FjHEYBFMPkfU/kfYcjCAKiz/0Cj4nEkrH+QF9/
ZO2xqyu5Qt3Erf9Uy/bk/BtmNw8VPFwfK3Ka3hHUtuQJCd3Ek/5DdU2hFZxXx/d6
iaZ5JNhUNONRFwvcI2YeN5GlL5Fupu4fAdJb7bm6hHcYhHu9y7xX5e/5zH3RTWH5
z8bVj8NA42ietIvQSwKSDRZPdNRz0cEbKQVjqaxbc6Jf29FX4ldgEtoBam3jrleN
FDxG3nFwq5TD+4ynsGb3BEfEVclYEQSKAjD0YAZf55XKeHaUwVeqZWvVlainpwFE
5ibuvNAC6/Hi3OVoCtimKq/nGik+JoGsBEg42E2WJkOzwLGUpRGfgvakDVTBRPhh
GR6/UveEt9ITRehZyrFbdxovPUJupub6wCYHyxIZBJqRqhveyM2kZGZ63wCriIAv
9NuAsEXI7l51vH1TSQ/qt+8tZ992b2pbq7Hz1wX9mht/pa9mDltW1qmcp1CCnTyx
VDu+Ux81Tqf79TLhYuLGQdGWmMh7mh2ueBC0OuCfDOQauFqClfezJE3pB/78a3fK
XzpAm8AlXhPMStKAgSve9g+X6SoLzfwvB+svBdLpnDcv/kCTj7M2SXSkjCxfWrY0
osMGsw4JgbYavx/d52hclok1DejllJ664GD82Yze54WxXz2exHkTVA3fKv/aBc8a
NQzDY+JG6rOrWo45U2FU5P1RXWtaQpIIZ0d42qbzUwFGVpKqBV+KwXGKbrFwZr4G
0OPoFRVUgMIkttg79p5NcTW2m1+dqYMYFXyjTkhVp8XrFcZ5noLvYmI4RI9SfDQE
uGz9lJL8FljLWuytPkp26p/haw8JcT/vAFqWvkTebJT9+VxRxyvH5vmIZSnfn1S/
vP8qO59klNtXjfMnPYbaqkmmmpiGEoZie8/Ozfj9tZPWKo+1Gx/xiuQNB9pHboNa
bxXBiJL0d5mgA1DaMQqvpeJRgXNqhaX3n3Q+fdj9WMb+q9ejjvPK3IV3CwpZdsdn
tm2gd6PVW6knahQihrXS87ZMj1mjy3P1b9BfCHk9YvJE0RV8aAvS3XAOy4mgqIdb
U1AoyDERErZVA6hLuSv1nsCSNPtp3m0YQ1U4S1ZkS/iC/iUwNvIPVxp4ZuUZIcQO
TJIzf9vH1ZJ/LHcVvGj3iwp3uvEADFZ5MBHmn+YkAJmEJN9VIi608LUvzcifIRYO
mYPaMYa/oDIHZzwIPamU1LuVdU5eihJNgQjzIpe0n9IR/j6pqddRbJ8OebtufVg4
jSEhiOi0mU+85KJLjE9YeRlzG5MkCvi6jlxGUz+K9nNHj4xiIes5UF1rlVULaCpb
HzaSt0ZHrW4UcbvXTXhv6LmsNbSTa4qFwBu5jzY58I3WyHAjIqvxCxesgv2Qg7Oa
RtXSF5ryTJTG+oZyH3xvjFtOmsI44QxFP3qNvgCpRLYHR51OkZkpT3Q3riMx76Kf
6Csn/UZBwgqh5En+kbdaviuyF1Wp5qU0xGv4g2eTaeQlvOHNYLMKvHkCvh7k9lts
/aFno1x8m3bIEderHxYlaXODTa77GlCu2aSYZADhe8DkXteERJwHQ6DfZu/Lhuss
4u+jiGKPGXLHD4ZS+R/uWyAdPaIYYdnQuKLM+g1zffX9LVLwMmfjezKRmyeL7Fbc
5Kfrt09//IQwxSqtc5ka1tg15kWKzUOYrGIzLEAPhOhrzrF4BcuKsuOv0fJfBPZM
lBPkAnxJ93HaLhYHNBh6wErEAaVPiP7sRfA49jF2bB0DA09ZX3lVdlQ0jKm8kX9F
k0I5uA/3u+CsbyrDSSTBp0CJK6VMNTC6kxawzDNr7AsP3pBbkYgPZWV/E2QsXVX7
nusd7JZU7zunwVhO1sXqY4+1JGEPrTh4cOFoTiW6pSp4pnaw6c8ZEcHl8rj6RIBK
5IyxUpO58o/MnSMGPrA0xHQDuPfk23ry8122jx6WWszjWklhyucMCEJpcLYs+uld
/slCmGtHLzxwxwfYNdZ69jXbmJmsOQVNnqQ/a1J4lFnWb2B8OQc15iag6Dpx2trA
lT2fC+rL/EQQr5K8D/UQYqeaEZaUWoEtKR/VHItioD9eQRwLShsIDkQTGQ+N/hLG
nzM22UX2uao0NgMqzjl/W63KsU1G+0JmT0AoxI6TBOHRN13jNyT+OqqeIdSQY52p
XJMSqGjJZiPFwT8KkWrtQF4RcL/6/CBT8v4qYNb8Kv9u0fEUbAfRXizgADjM8lWo
5DqsODnoNsmG9wYco110BsOH6uEWSjzyxLbA5UTQxOFkhT+tnjeYc12fXAxV92ey
OjVf1VVlCAjmW/9VQPWK9Ky+mCkgBNkkauzF3ch/btFHvW98aC1TTEoQdo537WRT
hM+XxdkukKuJrajmh0acte4VOtqsYkVkwFBLPkEPWgVkA7fWxvDB+sovoRsDzBEn
wYVFQZcUZOSP8nL9EnqltbrfJqhmb9JR8UtJQaz7LYLi/lJXyDffUwKjm0uL3HVW
YuEMbVgrNjocYpHMjsPU0WfAAestzFF2poa8Q8eA5LSTNqiAFXHbbzXdNYsagxEZ
QiRUujr5w6S0i7s9srZHuhVONp5uFOvHa7ju/0WFf0QaHal3FfoJtp7gu8KIlomI
4ZD+Us9c7xY7do7qyXeNGplhQ8w5hqtA7z88vnf4MRexXHySi8l+KrWhlDgt+iPl
7k6cI+zslGLlzuj3mwZNvxMNOZKg/QoIQjnx4VybpyXJxd62kfmIyGxSeYcZid4g
IAiSsSwy4szrQrKGMudsMxAqBlCEapvEOiIY6XfOTl6ZmBNtZL6Rch2oTkVvjHou
At3ybpKyOWCnHsTebxf6Hycno+acGsiUV0c356mDeqf3tMmri6M5b3+/D6Zx1bvV
ttGa2vhQ/+qCaPGbp9UCiCyf4V/b9F4a0H0COiPF5cUV6y+wqgCr6jn+FSP2ImxH
0wpFkKf54OM0EubUedIIaTQw0zsw5AoNePOViHeW4Uuk0t+HYxbUKV0gJuENIeeg
XOb+WRz/Ga5lTovcksV3+Qsyrvj4EbANrBJEFQuj4m99p7GxtSydNq4J5s8lnEw8
E/53MUrXHgpwfV2NUma9qtI+Q+kv9di2HgNzA42cwM0zrn+PFXdCc/iYt6IlIYgK
r0YPjAd9IAksmtL9FDrbd8BR4uB0agWXBaQn2D7wvfRdeRnwiCnieGbQcVftVtOK
FjaEMe6DyLuVIe8nc/4rVqS6IbwfOJ6PNd+gbtflTKzeXdtEmauh5PbZo9qyflJi
AT1iFnPXr6ZzNrEMuZUjhVoHrbhsNGF38hhmjADl57hOUTaITNPX/jcTVAd9Kwnt
k0x20QLsoRnWbDPE8KdZe4hwqTaQt404+sQjJlME8/3JEeGtqozhVD9lMzkm9kaz
Nr7M8rScm3JBqzCRwNVPuFiXCYhmk6ax+tvPiSZr/2SRJzao4wf3soEge++GW+If
cAT/j9sj7/V4q8BSikF+0pj1g5YQD2PzudtFuRdA+i9FColSwlX3ndhyBLiAw04a
LqSZA6SHIcu3yS222PEaG4e+UE7mIwlJAr5FelMh0+1xfOQA975f1qUONoPpikZ0
pGZ9t0VmoxcQP3pbMRNLSFwvjOBv5gHQY2QeRyeTUUVtH9cpTiS/fvUiG0hugAxN
AJm+fhyAdaM3t85vmqRG3tW+5BkkC/TTEpsuKinshRHMiFqj3l0JFii2SbmJjOnl
Weg1M6R/1hCbCO9vPTM3Gu8f7cV6GAjms7sc0aB+n/mVAwr/yExFkajcfX6biPCD
rqYrGcyiyx8J4LIoS6l0ZkxBKZyt6FuW91H0Yr/pr9J3HShVND5Ay5A8wVaDL/48
egrOjLPRs+9/AQmqnVzaOay156kufExi0GT71tjoDHPOkEjRWWh6TG0cVIu1pB5n
6yXjrf0uRqz9B6J0CTSuVwUuSdXGzzLvr7h3zS6+MVi49tcLOgkOE9l0JYa4UAmd
1k36kLYmYK1gMHyhMdMZH+bf/6coonOksyMD+az3Z/Rt9TGeyeCLNDFLtpqXHAjS
MZDMUFWLrHa1HqAuElCgqq8J8vN3HPN2707umlMzt7EVh/ITzQSf12iCjAnb3RIS
jrnGNJxZuTo4cA9u6HUNwKNJ+tdXkEv7txqxKKae3erM0BwGXi/z02qjxFK9idqx
56/h8nyRdN9BQ38hVsySVq+M2RFbc0gXwkj66/g/3FP6Qhs/HlJ3QB4TpJw7TGiU
DdB4Wct9wEe5wheL3/k+5lhpq29OPxnGICfvQrbsg84x+VnV8NWt2Zcwzez4gpen
AlJ/Pso2KTMfY8rveuGa8SdkL+x0cnOGu/7EBipzx7fvJ7PMzXX8xbz/w6hgCkHQ
PGpQnJm72etfffeazMcwXpAxuvo06vpxJFk3QqG1TDi8UX5F7mFJ0b/DiYBsRxiT
zq60OtTkV2vm0N+/1P7uw7w6P2bvU08Yfd5M9PPMSHgSdODhe4VfBzRrxrTVQvvv
8B0GXT5La3WREcq0ai3RgbxuwiYV0RMV6FLHqHLABSHzEQ5zN6ZXdoQ+ibq7q/Bs
SPTtR1QrlCSiVo2scJaTiqYXOoyOsdqt3blKT+fclu9Xa27RGwmks0JvOyhVpmIr
1rAdvoS7OsXCyjjAttQWBfmzgFqK4X7nfnZ5vmy2MR7t8i2NW55qbnPhcgIHP67O
FfRmWQRGYUeaH2cJmmjA19tV22+97ywXVb+i/VyXK+hz49e3/Kj/QrxAgYpeFcp6
7w0GYK/KJ8lQZ6CX9CXvGBoTO4YYCbvSugRZRqNB4oZQgPoVJf5donrzfXMdatgh
JcP9k4DFBPiFBHAgm6cVMRigKYLvY2Cl9NlpMuPJORIzLrSmdIyKg9zJbQfW3OYS
i33xu3uL8a9Wamk7T0HZGjwAhubKTbvWiONdTW8M1ndCOkEFxXX4gaPNhGkhcU0o
b3339nZ+001+OpH2ZcRCV0JB+oM4osqaGmXtnTjS9B0ZA7yH5VeV4NZT5amQwtZh
a8SfIx8o2ZEDABIHWABCgQSbKjninFcvEP4Ww52ErnGftTKwlAJaH63C/2eN8nGj
WcitjyAzrn1nvqQ/wK6x8cQdG+RppJv6FHXyet56Tw4/68hoghohgotr64FrJKUv
8OUFFFCzMSFkTE9MQ6z8i8WXYYBpGrCzZYQzvLtIIbZeB6FhvVYCUKJVq0xbaGfL
Ql1WJCeCkISks2HR+Z64Gh/hdASPb6pDJLLIBtnSiOOh8wcLLgsuK3djbnW10ucL
J/TWM4gNqIWlmmAQeESutUgNzmZNfdDIgfl4tiIZU+58h8dom0zQVObuygzl/nvA
TqF3i+u4ML5/og/tLOKH5jkOiZzj6suTl7Bp5zkBE+HYOGAaXxQ9Q6xwhgAIEhFA
F2vmB0OyYTB6ehavud3H1vFpDs7+XcEGlZ+C9cdS2uzwOxK3xmHB/2BJrFqrIWgD
rRUfWcBA19ocTZpsOTKPKy4NTRekGgSpBWJ0kZ6l6GdoAnz5HNxZUnDg++Ax64Xs
8Lp57FtV73uTzmzTn+OxZ3y4MrSyyKNiaV/wsNOQ3xlpu4QmucHd40IbSTGPGTPr
lSur1qqHvAfmhsVrEz9XhLVPA0XP6k7hZ6OZo+hN3cpCWA7aKGc9Xmu9EVq9l7ZS
sWjh0fZ7NtMtAIWnxr1xwVM9NgekoHzpy0pNbI1gSkzIGqGwF1c2p0WiiuROqDBM
7t2V/Y/tfQnKuOCw1SoMuE8mgmSauVWpxHUgOuGMRrevVvuJb88RirF+cbohkb3p
Yl5KWsdWFtAIJ+X5f6rjHq5kvBH/LNRzpdKPVXowoOcjhC1Mn7fq8XXXrbt9co8O
QYz+iJw0s1zSrVpEyIApmPCbPxGcWHkw1rYbySr9GqVeO4FOo7y+unUe3sfIw2eR
VnGAfFlS3GORFBxQlpSm3RDzNjU0ZEDRtmLQYF4lyUzreR+DAQZkj29uKSoyHi15
Ne7MTSuj0jXE35fTYZ6cqKywbB+s4lEvvnMmds7BDm1uaz9XEqh+mtsVPEkeLC5X
uchg6irrfToa8z07lcEIdw5cpMliLkUjUFCqUbwkNZxFQNkdQH8TinUFm/CF+Gud
Js8PhXsWM4V5UOeeKMHCnyOHrNfsLqWIHZNgt/dxzrA7HFtTD0o95NKAsdNGZseb
e6pONw/ec+OqzBIU1e0dXmSUBsKQ14YaK1ANeKwTeYgZZ57+zLKVG65TywbL98vN
RBmZyYOjv429J6Qggxdbe50CN1CZvP5kfAiRpuRNLyPkwQwjka3daky3Lq40Dyfz
4t2hB6dqlx/ebzLHvAP+Bkdm+9F4TW5IO7uix+MYpdGvMukluv+ww/wqiuBd2Zv9
7l/zQy+wijSNN6PatHUaMhDn42rcx8fRduTQRqAOJt+A3LmyP90m1x59mlZ9tGaj
X21LGyNACk+NfiRQo/W3mV0gEc6MOge1fq7UztfTxvlVQBf9MOg42Z1wAy2cmmSH
Ct54jh5RGUem5S4IdIJVSbD2Insx05V/YRo17D8iG2wBjvOywID6P/cAv2VcQ+B5
j30dn165Vq37Txko7VzuHF4M6fpUwcU0LFwtuPfxrRP+bcPs8PdYzJxAqmEAxP0k
ZaUlyjYGH3a+2xFuksqgrnTHbhNP0vbVaMXp7XSuQ6GRr9aybDX3OFJdhIgjZF6y
42a2b779uqiJ1Dzj53g6Xd0lj6Z+B5AGFkJymSGSF5+zrmMf68a15JMg/kc3Xw94
LVomGnShfDyWRsuWlMe/tYT02Na+TBggSIgMQSJC8ynExayPJaZbR7PAFEXE6OIY
lCfEQu/EsnINATds2+iQWk7L3LIW2ydGElPlqY8it/e7t/XY7oojegeuC/xPIJdY
AbyN9JOLNMIu2HMnIwgTBy5FYd3Nb//06rdlA3U3VGOp3AbOcYlt0+c1VZyFyEl0
JdBlax7Q9KijGYje/DfoKG6yfwAnbDkR5AIH1a7IUFND/5rJeyC/+RbB4wsxNYu3
BFxznmkAj+eGTnL5rQVhh61WbDktkznGnOwOUMGPq3+FEM3b6aol6ZRqtflkGmxq
7dS1tHgiwlU3B8Zbo6AZNJcPqOQyVl/5uWXZeSKNaSdE66C1VAUbX3iy41rSD8Wc
2B7xsYhxC4DoTX1DzYBsXqsmg1WgM/7tfSK7NeY5J2u2pUIUPlncReCS7vv1Ahe7
Kjj6ZtjFno/i87eP/J6EVQfsveRfvUXK1bmAQ+BvfY6d+0pylEYvxW4nQ8N8Rov2
LhbX21/nru9x6iDKGONK6tCcToPENpNDBR3Gpt8svCBlHFf3aPmiZkTrhiQtckkl
kXS90eKKzBnjMOffefpun+WpDX2SYhuBQ2IrDLf848JSZuPAhBsNxKbU5v116iKi
3bASnotiF8iL+s8+ykD4kmLePgtiUONptjJrgqS/RqPi0ZSyshW0dEJejoV2yeE0
x4gzxDNMP+5QwRLbUhzQaF+y03Ax36WPn6twhhbRl8FLjT/yIUTySUSuaJoaBChu
IJzzAr9FweF2F10ZVgqVkZQoYR7BXXVd+GShN3/XVOBMkco0yERzQVb6LvdUqFbY
BBcq8t+i+1sqP8OSejguLosFyt959JiQi2pokha5FsUFe20JYIeDOqe5qfrwJsZo
grAYIdiRf9LIxSmRUGqzLmpX4Z9j5UqtmYUUb8h0uRBdwtmAlhqsb3ESXB4pku+K
hxmjcT7RjjoS1ZrNSiTT/dH87ZjMSp68/Q9GGbd9uoKW5GYJFuVPRtY4BJgbJB85
edWZJ+kpatJTKxBEseab8rShkxSN8GgdRo7EXoPkpnGcG2Du55fpEfVhk5n6kren
CqEOBc/UyMGDFzayw+HTdY3SxiSb2WOFTsvXjxg6QaAKMfRfbfUHTv+C6Yn8Mp/h
YZ09CLLF7jtyWl5/v48NPStfGaHBIGMjCJgCOKnVG1C9RaZC40uqaJvxPOY/ULRO
ckgaTLeel5ENJbC9tgtHQRDjZBTzFFbFxjMcEWXMb1T0S4IFZp1eOt0fIeVLp285
3I5fKx8tH4cvVHOGD622uGrL06of8ZWaJYj9ubjJNhZm2LfI/uXPEmdxY8hgmF8u
oyMQY5og8V/oSM3t4eNBLxAra8WezObzUqOQFqZU9xdomR1trtNJ9kl854aUsJvx
jcYMMZIZBgMKAw5UYgV7buTgYglgTqNKowzSyILEFjJor/TN8ByMMN2sNJVlS2Zq
5i8rgsGqgUQPb3SjXOmd1caF8fJ8v84BRou2q0LCFJR1fuUR0OLAzL5ntFrzgURr
HnrtUe6K2MoTT89hj79O0OzoeAlGWyVB4Jmpa2sJUnk5Gfnfr7ad66ch7rPAOiuV
BI280ucs1XHwRxb7MfrBJMoE2iWMzYRPuslRXff680p097lOOsDUyBdLC8E7d+sL
CVNh6HpYiCZeD9NS3BMbs7AtJWCecjg0JAarU4H8T5chKPSHQqeFdao681CgQtTA
danXDIPU3+ErUPurfJz2e7hg22BUmNe5CE6HSjFS4gcctX43+1+ORCR+PO7K9hvJ
BXFG/5oH3xas1w+ky+uLxtgQYf25DI5hQ8syPDkeFg13jtULqsvIZcqYPz6A+iEn
e3CtJjNUfqkpZfPE8sA344mnM9aNFVUDsoWutEt5hD/uoBP4EdeX+5LgSQC3mXOz
Px6YzsV56BvclItBqVXaC1ywuFWibCeSy53MYad0uA4aFlO/fY6aBSj9B984IfLQ
bF3M1oyWaPRlBzZi+oWO+8TDZ8cKTfizG4SeLU9gLIUXkWHYW578hWaPikKgJEcT
t26D5y5ijsDyn4RbCzRJ4kYztQuLrNVJK/zjZEHusXHKKuzKecJx24lmseEBvvQV
ovoraQnjMtu/cMAVzMP7LKb5nl/Qb3U78ooS1xaz3AGzbEVPZL72j9DamKmLq/1u
InFSzGLh7WJS/mzbJngjOnkYSQnTscFle+7OU/Cw+gUPrFqIWZ2sQsy4zwbFqeNa
S1cLASPWDl8I/yCmxzAhrpi2NDB8KFqjfT+k/YFpHeFIp9LKtIxUG4e3sHVo1x2a
ssM+giiRCdswViPCH4j5gA9PPj7pZnpwglOR45NnnUBLozI3Kf1AKCwiEJ2vJZbJ
VWAvtA624/9KbA1rxf2YFWM/jQoGN01DkZfUgfTD/zZkGGfSpH/0knUpS/XzikgF
Z5f8KJeQc+jVyZcqsJQdbDXwP1iVteY7d5B32M5/phA8VxXItQ4KsJg8kd4o/8+1
Yb3oCIhrgC177WausktVZQsUpEHyHydUFrLT1FXFp420Z5DA2J9GMJFshS8Qj4Mw
ltE0saXQInKkXuKxPwedMl5iLyCEJ8aXgcyEJoVPuR2kKxlu0pJTWDikOndzI/hl
kCl1QZ7tJJhWkLM0g93QVy1sNWqkI74LzSSfBgktdwnuxwWRomI8BplSGWpGIUEZ
aml+SAMUJ09wL1KXnetUG49q/wwUGjljPJX91D5pshxSAgBEwcbSl4mIf0bAB5+G
aRXPyRs9a2VXDEfflvccMQJK8m4vVcwAISIkdSxcbogzyFxzd27lDDDi0VOCUAQW
QipYPVWIuA2+QnSB1yxAG9d9bFAIeKlAmz4EjXu5ZuEFbaTodspdyMd/EvYu7NG9
rofKJPwOFTxrOT1liZgIHwa3sjj0EIlV0Y6PE0ZP/T3vFJ4gwSp5zO1TrmHFuveY
vsY2fSYIuCiwZWPjAnhgY0W+dfNqU+fEDTgihpfOO7PzPwqWGv35lhtgCj+s4LMN
MSDqyPSXi+WcgGd111MhKTkGP0dunc7TfzNdz9AYgeGDqQ7x6+/5Q67EymTGyJw0
1XpPTjcHb6vCDiUN9P7ip6XiXLgYPB33cc2IG/H5OWAnkvFAfGSSj3Ih6vSBPZWR
aWFyDrg/7OpYRNtytzjFs2qJ0dWWE52xQ48x9YwP3UWrVGvpDqb/p8ywYkagqMSV
tD+nDj44Uhtyhi2QMVhICwLB5H5UgPWEX4c/Vs4ulXla7AacncHNX4Y/6ozBoFp6
NCFkC4BR4m8HHpRGBgc2rIE5k/RYKjtvKiIlngf6+a6WhPETUyLszR9Fpbd+uU6Q
IEseY1cWmVZkWamEzJu3lFYHw89lEiu2IXMb1vfghx7gDGLOXg7KVHSxf1/5jqLm
F6H0UTPiOxc3ElIG0lB1B22rg1+xLzLnRHWVvq9SBVOi47+8vg2+xvygwAeizXF+
SD5ybSJXfohEdhszLcFy78NK2sxlyhk3Y2ZoWElsIUxNqALL/76VF1LWKc3sD8kJ
mqG7UCPmnovFfjSJqvHeaIWfe+8wvtBgyCiEmnclnIcrJZv9JTt0WnGmEYT2o86o
HkeQM/7Zh7mIlm+pfm1r+Yi6cI4opOxx7ROmzJ1bQUty+S2EIH3yytRJqHLkqZ6V
FGgw+W5py/dg4ZvzYM9AO20zbq+oKL+Z02DNzU6hdkwGqgUTmDpa70CVAf4SbJdi
8B6FCHVlJV7jkP/mKCt3JdSvvWK8/DYVQY/fcdwGmVQc5JWBWN4B3Lbd+VXV3l5+
vFC5lwzT+UGq+0Ok3uLsWfcKhQ0i5kBihwWkeamwCK0VFUNMV1jkxOPQozLkqYtx
ljiHOHiNZGGIW3ioIoYiO02gXCywPG9eE+DhRIkTgp9mYl70u6+CPw22MLbvakYj
ITag4fQ8fqX0802UdxhGmA6YrvSO9XpzYPnhnvGiApzHqvmuRlt+vi1wWajNlOL/
Kc3bKMPHKOn6zeXv0jLcPyq9ptBwEdAA3K6ZDdG6s1hSYjxX31OtxXNzU4G3b4Ci
JYLz/r8opte74uFXwPmYi0mYXLsNlL6EqCgCzyXpdRn5GgxMkFdIm+JU26IcwRlh
s4Dnib7GguXmlhwcWQeVWHcpE1RrQsFSF+Um8a8P6JaIhZOOcvgF6ajGDbQNV2q4
Mw2Xc6xDNtDz9RvfsAdjtstVrf5lX07/bHB/sKNM2F9UXit+PJc1JFM1Jy4XIM/V
oRC++LV+jPRjUWwRGInNULefhWw5qtupAFqhtXaluzt5aTdkocxsfZ8t/eTbEIJY
5/gb29yN2WZZub7bCT0LJN+vJ0bmOpbC0dCoHzYjHmhUI6/GwS5OO/ITJxEut8Q+
oEupu3s87Y1kr7sbQA7hHx440GxKqApvjmgdeHDc0HmH4+/HH9lkvpr3hYnnBwfR
FfFNU6w4XMeqRuyr59ho7wZXRCq/zkb1qdNe9F8/G/sL+Y1JHLku1zyAATGR5Q1l
ICZPtxI0jWlK3F7MW+c+VIm1L0m24WS70/7k6LhTuva8h8Qd8mZcuqLZwSv60u/7
8eFAo5rOXPKF9Rl9TcfK0NM232GzK8snpZNY0kjfGjYmikMstBFJvg6AXaC1iQrQ
xEtS9fD0vXHBHKRVDy/V4SOGvoOq9gJuUj5qPJHaab3CuyZh8cWha/X3rAMONVoH
oV+1TLq70Y23IX33wAlqbOyeUCscWrfk8/hUIalHOnsSj6uqOGkUW/peMpnDs6aZ
O2KXbh/nqI7RYDUa/i0pFZCzcfPvpEXehKSgKLEFZ3G4N9UX59mmL1gKt7rkAX0N
X8uO3MlqRiPq5hdBeglQPL+UUOwZqq2+9VJ6FTucqiP/Zrds2ENDMoWu074x2rmS
HNgnFRra1Hv385lvZlKGKLaFY2wlEXgM+JkzacMIFqUQdf4L7sCIUHHL/lSVrgov
IrMkbSBZ4XHEuQxXy8eOpo/UpdzKqFp0FiBgjjDOtf3OrcS5tXtaALBaJEZzXvvO
wif2z9YcXs25yQ1ZpakhaVdPRXTKFN23L07aAQCti35VpGQTZfw2OAg6M4okoqZa
BUq4sIMULntB7ZYlVu7fhhX0RVBOWXdNwPBac8CGLF8SOREp4gGHfuI1lYFSNBzg
m1xeOq55Be6P82XDgiQr1UsB6caROF3vnbQG9/EZuMzoIAjCjfrKaSBvyqqI33iW
hc/cdqINDTpDAfj6mq9rCOLU0e79iliwPlg4EMQFPesAIVJcOuRv63iVLBZ7bPw5
yZZacfVGKXPu7d0T4CgGGhsEppq1C2F5U82qXQOghBK1PmKpbDxA3o2zuu3KGegY
7p7XukgC3Q1EclPZxMQbcLUge7rk+Gz2sjKM4wMBaKijeH+kfl70RPztcJ2Uc7Ca
NGSKXIX4LLUu0jSBi4Ooykbebd0iWv+j9R0aNEaKAt/tA4P5Z123t3XxrQkxr3Bh
CtWiPOLDC7nv0OEUVJ5u6UrpFTzgxDRmHKXwHGD8AL1XR0bnmZvP8ILRNFu2lo0Z
nsTLVDCGFmlBUYXkO7qcSmd6ODnEoH2bf1nHxlfhru6UhHyYIZlG5RwAz3fzUGw4
uDI/kPyQmlZqaI7+6q0M+lG8M4vWsfStuOcQvLadtsxAR7mTk5W9vD7Ou/tlMTlO
n7KZiZrvr52NI0xA8uJ2mrlpsSwqsi/NVUPW4nPuG+qHB4UI7W7GJAtaMNDaeIMw
Eh213ByfV09dKFiuiT16ziS9tR8DlWn9dAHE0lHSe+W9wiiLGduKOj4i18U6HfnR
uFa5h71cl8yk3T8ehkY0bDdn/6sEWpz2528X9ThYBNux2vwUoYNdebl16uxRyzi9
MdOadDMrKuuRpXOFZfDxyKDtynr4Q+6Bp4lknFJqxlxjQ4BXBBzjCdeNH8K0DDWD
zlaTkZFFOuKJCYPoFPH0KynBBR1+TLmEXzzGVpAq8MxcgYVyqHZpfseFzj85L4UP
63uuE3CMYbGjS+bbFz6NYpf6IUorf7Es+Xu/31e1jdfa6pGUKOIA4n0qRI4c0GP2
ddlkg8l5aPPYxaRybUZkJHgmhGZoZ7Z0oXoqjZbtQSS/lmLw1KegYtezrEw8JyLZ
U19j5Ctn4aAeuo9nEgDI0P8CpLYa6ESZaXZhsL9hkUgizm16OTUBcKwiWOxPvIjO
iLd7czh7FkzVOedsp67sbFnpn/y5n67Uga7QZ1mM/WpFdY3tXa7CxMLkgtBjjWn2
ks7wJY/WN/Tlt926dYPsoSNelAduewcnmiX5TiKLQKHowT0Z1tccXJm+nHTLWflF
oIHE/UzHe6VORy4Na06SIcrte3ZhDNqx0OkZN9wOmUAWQlyrNIoW8MolbMTKoq/b
eKrgqb6OqTPOS5zY4Gmn6pYT/In5NquSAA2YD2H/typ1JIuqpfooLi3C9eStVBIY
zuLAZv3LKJZosvq+LyKbm8BpWclQVOIHO4aDFU2FDS9c7G/SJoJ1yXF0DQwzYlwd
DvjKnxNBjAgtEXmalk+Az9G49rlbm04ZxWv25UJaoPwytn1ZSbHcuUYpyHFDDWrh
5SY3x0iOTtI8Pdw1jaleRIICLEea5ZsLsUYqRvz8FVAdYMSQfyP9ey7dIIfkg2iV
Ffi35pGWsTrnD/BDdMavopZ4ht5bB9pGEjIZ7ZWPpyKYXtxaadzJq70yvSUcUd74
TJU/lo0+Fm/koHkLmzB/uK7dAXiPNPy8wpqNEdp8FYha5nzSNFpi4va5018XW11i
Cls6/35sQ6dpAYVwTAmaMpJ0YUP7zmcWkC+5HgAsES+SWczTZumv1J4JzYzRAk23
Ug/YpzRXUNzGr76N5FPTJe5GnLbALGpZjbiDYy0zsnZ7V9zEeY1CXzCowEv2Cpi9
Eowsec8rD8orZjAzKghpGon+5keim5NUnn3oYyjBy72UzpzYnKgf4YPgfybPE82E
yqbTSsfaJrqsv/oBhsD5kPPmtarGG2KUMj9Cc++v/1o2mEOuapLd1Clu5Gn0X+jP
k1apILDMJKKUdI/0HfM+M2r+NTyWBnnmvB9m1Szfhcz9q7sOzm4fs0YYTcGUm/D6
DvbcFuToyRXqVMWiknSB/yIZF2rCPi5F+RBJFA+6POA0mZGJ0YWzQBpIk7eyqi9c
l4qXL2kr0zu5XNiIsxMD0SeG/BhE80p2fA+yQfOIMcX8uzsI2o5BgXSCN2m/dCzA
StLZJJbQL0IFtKKbI7k2bSH/xqJkqW9bQmdpicyj1GKAE6gY7XKkjY18Qm6ZngnO
1YKlsBjeAJeob9qZHGJONapu7pmFn+P0FRbvUdlBwLtKS3B9/jJ0FURVUz+hM3FU
SscNicpEoQw4O74GwXgkBVT2dBiY4/0Is6igv4HZWY1AkIyworNY+hjovSZD6vga
dYNpjqqdWE2AbOFzlt0nDbjVX+9YoYVbzJQAlXLu1Bjc7giVmubp+W0rzMAwxM+t
CdTvD5dUDqqBOtmXYNjUJvmkWrjfQhIlvff4y913JTaien2/MJ3+yVOjmd45UW1z
cKx286DP//UgT4P6aJEREXy9zvMF3nGK4pUNPd76E9XsJlVpsp+j6z25FOJQKn5a
cVZ6siEpFfmNtpcU9By9xXytySO0j/zRxy5aWR2tfJ/I4Mk2R399xIvjQqRyPX1C
miD+PdmoPvXrI2z28cFMrI/I0VhA/mvwoRleQ9Z5DIo4P9qQng9xHCFeJG9LLxM8
7Xf8bPL/+uuMyUwpm1bQQ6WqrhBRDoJdtihgLsrp89WzxNMeYXect7HmxStA2jcS
UBDd38bm2s1CEOjpClcShmA3+xyBeCdCSnbyeLLoch3HMaOkWuS8t4gyB7icgnjI
8Z4aDKhpdTmBzyTfFRcMlTJ7TmQOlgrgsu3JMCYQpM27/4MgplAznfFouE8BCikO
R+PeYy84pdc7GP54+IvcsMRahEoCK8nL7n4KuLFULnMwoR9BzUqFMUZe451RsYcq
qd87RH4Ah6Pn3Lwz5m7Pk7Sgt26jDQTdAJrjP1ZiOlBYiEoVI3xDIFz85t5F1Tbz
J3SA9uSKpojKMDcZWJR2zAmAjPkAtqHaKUAUUvzcoXP8oBWBW1lIlwAVrtJFfUXm
X0aQe+NPdNZ/GL2EPbITTDLes3CXo1Kl3sXCVtt/sho98Ay9EYr5Ex/bTcVdkaTM
YPW7AxUN2qPqcczNcUcI1uT5x52F//MewlwaJwS0iArAqBoqwvbLAE5XOGCNActL
oBzvSTo0n1N47EWKGsW+8fz7WsSVs7wWP/PrJsTTaHVPY/gww3n/RCQJfYwMX8/9
ATWZoKpE/Yt/eU21v8A5Kyhq+NNxw54TSbRLOxOf32JtNt8p6VgBBZPVzD9euAqZ
QG8mhMSyezToKjg/gltgMnI2dRqO2Mo2eCf7xTK/uI/kD9MS0EHfdv4aGQ3h6NyR
HeDZALTn0o1NcLaGV0stbijR+yPNud8ML473+VO5Tzc4Fy9bHBNQv/WmhEQ0qcG9
VHPa+w7ULJmmMeyU+ZNgNwqnn5ykSDx7ZTSjrlt3fk3HAFAtHj7tcmNw1QXLh0BL
jbJP6+BX6eJrQOuBuTw72UUf0SUl/YzTZtXPv3Ru7C4b+5wBWAi9yhPkbo1aighg
dt13I7mGtPZRMIlXrBqUK6z41t/LmTs9cyQNS9f0PJnob4m5xjwRqAl8zGXfrPRf
0saPirJFqXCA197SJPtjDQL3GbQq7T3IcT1wbLv61865pbm1veAlPcFWssxsKFOM
UFSkF10GhEvnDkAoj7tUvEvatm6MaOczU7BBwupRcl2YvgC0aYrykPEH5Q2LKZ2W
Tzkczc/woLvPQxHbd8l4x87FIV/EAeNxa4S5JAVtzteI0KdGZupx+IgSQiWaG+vA
FvoJg1Nmn1UKC1jNKWLPmrOauDg+wPlnSduHQa/+8YvVM7IPQA7XXUnldWR5D/eh
YOMw8DY4Nbl7Em6v8Kyj5XmpA3b+WWd9ni2mizFsO3RPASg89tHXFsovMNHjXMtQ
jbGktoOC0zQSSl8SeWpkkqb5oAX/jWPHqutkGgb2+KZVmJYriEm+BbObP51F9G5K
SDY5qvkhgGbDqA8/EXElIQQABTbF1hFZvr3byAubbVjnREKEwbFTbK7EI95VUIhg
PN0ciS8lULwnC1nWeHyVaqcXKY57a4P3OvmgWSYFgPIskYNHKPJFT1+kWgTwrFDg
Y40avjkkR3MhgOgeHQJ+WoKg5Mr/qvxoX2izhJcfRniijWCkhqA+O8hODjbsY9E2
3TnWc6+3QseHL8qDwErCqfVxOTIgwmHvyhWRVu3vxq+uYlo1Rz+9sVaTmUW9vQyJ
TJiYeXMN1CZiZcoiR90nhiIibcy2rNlG/BFjBBwszwcWGqfJIjTln5NIkM2AmfiO
MyuVCowX9qN3GXQ6jfXfxm58eJN2opzLANinY5ylnp1xwd349f0IQhCG0nhjlqNG
6JLJQE8aJNp212D9/pAi1lJjmoslEQymFASxSFpRQIldm76pGVHt7NbzrVHkfCBO
GX8uW/t3OMUtyhVBCyN+N3p5RV/+8eVIIRed8CwlbQx6BtgL78RiqOGkteprL0Xr
VXvvjdGR0nd4fk9911V/sTX4nAEH8JsuXxI8wYpBSjXhJ9lxQs8fCCV2nLgs09Ir
368e0I4pRA2JD6PoCSIekp8F8zsqsoY/8xAqAAz+atoOAglmqWzv5yJURM0HvjZj
lNmh+id0VXpYgJxLicRxAi1KE5Z8radOfE/aqyT3sGH+aAb5RZKS1XVu/uPhCI/e
SZ7/byo1oTpsb3JvG2x8iF5bIbzaFclV5n787QcDf7IVSfTLoMGNGdMmsppRtrOg
kr4Qi8NlC6qbosjaLaaSdX0OH3R8vpOdhLhE3KLZeVmziDPqUmIKp/VmfFBGGKdy
uwhTAHcWw9aknR7z2cREHfAVZjzqxcfxESft/AJIiN1ZIcFDqcwR8uNPGMtLLqpc
cwzNHZpCTnxoiB793RB+U7PpKtstoBtJqC6XHNg6v/OHL1ZH3lUbpvrNtEUORAwg
CDgZMIqD98aaEuWS6yPQ5CYLspnOckezckogCZzUth4uqIEitQ2af3bpv5N1+GTh
y+x2HhtBR4XRp/vEYHT+oB4j2lEEF1gKwEGnq5MaDgVMoTooimJTqYhz+QYFbXoP
8VIH2mSq29zbN9JiDnSTljEdC2Z+mXpHbnOX6NEJVrqjCL9/NaZK9+4GZ3uiF4XC
zPcSKmQMoGYqB6p/SzN1vIyOdNT5kb7KJMXbv4AjYJQmB9LTowYkyLRSTaFzjQlb
g1hsrqyGoDmynY55g0SM7cqNEbb63WkP00x6AePk19BYWLhS27ttNVeIG2ER962u
c5MhvUOmSLfieqnJGsCxErB9j9Q85l02m9DDuZfyk7DtWw2SVYEckm0PCO2hL6je
iGEpxNMU4XtZWmjiF1xD7cJ/f55cMbej8Da5O1AvlKuSm+bn2ZYfjrGKP3GhoFKd
C06go3U9b/OaXCFyls9xUCgIekeGLhO6YamAS3mZ9hgnbLBYt/Nzxy+WtkHwBdpn
OJvNq78233qyRTXzVE2lmJ13DSA32j+IT2U4BMK9USkfhODJs2Oa5s7qmJMGZuVW
XcR6M2p/mtmHlR+ldjsbKQIsDFvxFJmcYWTKOkh/8PXjn1KUdYcVfZnAsyIm/vLg
E2Xc6LHeIYdjVh4hPzYCdP1y1Ntj3ERlXg8iF2dKYn+V7v3JOwoaiCDHh92lAFIT
v1eGz+DLGI5H7meI8lDkDFYhOZQTbmyNAlPH21qs/KDkXpfaEfk26HT0GdPAtxqc
5lHmRfch+sXSSzLq5wybI/yCragsU0ey0iimhNzCikRn7jn7ZsuYOh86gMh172vp
oqDMyyrCU7LTZDUwbdzqiuvQUNQ56+pvnjg26ReuQTO+XH/24vABBWRNje9G06Sf
9YK4vC9nuXeEwXoQYWvakFpgv7mv4OIuikeaAoAlXwrisfBI0DXboGUlnPf0vl3K
pcfOmNaWKnEWiAT2DR5RUKHlGuCep6lBXeKy9pSS0m7Q3VlHwiCnsiMzyg/anBqi
i2+M5p6zkrA6NbSmH6y6JVN48gCax3K98HNw3/KVSgRquTb4RELfmpHdMx6b7X4g
Q4diVbehHDD7GW+VIfir+jOcBEbMl/34H0FGf3wIHryS0uyvA9CyctO3aVs2FYdy
`pragma protect end_protected
