// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:42 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
q8PWVl3CcaJhCUzD9qgRYdRKo28TlnikkQeOyN1tocWpqkR+/Q+QS1ELAQwAiWUo
b33+fqU2cLTygmN0ZNEzLbVib9Lp0IR+mGWFg/83cdVPlEBqlrAYnlUMHPcQVGQL
XGSsPd88IDVyHxF2vJx4m+cd6jcMtGjE0hb1fV2pZ5c=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21760)
Y+UpcZ8wvNrLhFAus1ufmDoIhon6GRItWB/z0anpfeLjv2hC3EjySFpM/mFn5cy8
IOagzuUjxPhDyX9nIY8OHrNwNCi2jZJWH6LhPjiTnJT7lgkNE/CZdwT+OJUE5qXc
TDmkWCFkonNEUvsP+BA1IzfAV28THh5TCKSDCVPr9/pTEgIJln+paGrMzjK6ey/m
JPAZyy7e+dkkZu8C8HlCYa7A8/Lte7tSVt/iW1RAoBhtj1KRWmDqGD3AgTh2BL+h
nRZXpMVgVUzd98ydH8c5fVQjMklnDrs79BgcRbxIX98q8j4T0E9h7s7eQdCHKxQC
OxmhL4g4KAwRfN7dyXeNoNjiqOQz6cESlrmHPYSRmbmJBzqrlkQ64rQLxC5i3me5
El5Ly73HcY/ZTu0yzDSvrx/156TbXpK5KkVd7yyxLdO1jtWkcKxQOHsYM97+I/SB
n/x+y+CdLczPTNbJKjJk2KbPAD422PZ3p/60ywP5MQ64FNSHOlzOzFBMnuo5rSaE
blVGNJR0S2Y0Cu/ISru6DLRM8EJNmtM7RsHErPvD5bl8WbT9s7NPrKbXq/RLgymp
N7ByipeG4oBA3pEJsmAXnTmjNY2V/OU7Eyh5MCvWHeXZxtlVG7vb90ZqdBS8uHGJ
OMwcoOA1kRbi+sQRmohiwqhWUm+YxAp+HH2R5Xdxa9uV153IryncEx4Pcy7eqN1z
lj5w7/u4315FgrMU0iTDaVHIMeOAiz1qJkzIni/nHM3z4HJ64sBk2yNEnicgofYk
PY04ieJnWPfSXP14rVwzsYfp289whxgBqdFZnOwpMaFQe9H5OlWLW1vHI/iJtoEd
oMSv6Tim6vcaHQSdNGASwo1KAeapOQjfKJdkANkLxutu6Zqj12KB/VJK13uwyruw
KT4uwUoG3m6k54cs5qauLtoFpBof4Y4E/KaRNRMqUi5lFHiUT1L6PQd3z9kyFPsE
J1oSD4C7y5CLV+odI63UiuQyrGet2Bx4OE5jLMjAV4C1cP4II/ML2RxPniPcp2w+
Wdzy4fqtTE2kmfE8rk9HVGVC+p0m3PypkgYsQa04d/FwRdi1R6u0IA5YTKq5oS9C
zKDBCevx7e8zRXZuaodlUCp2Qjj94ilL0K3IrE2/rnjHCAJJrupka1f2T2MOgQdz
/uoMbqFK9N9gxpngVLD7VNibF16uE26agQZ3MJ5VcxqyshErFB9s3Cl78BoKiMo1
L1DJ1xQo5yrrmB9Y3me+a3Z1A2okCABP0OrGd47QkRfLrldMP/x/Uozk5iHz1HlQ
tqGd5Sjc9+Sr+uaRHIEW8Z9TxEPxmJzADq7fmwizphfSct0Yk/Os2MxW9gY7VtKc
dtrHoXb9Qo/Psmfht46nOw9Gab2KELSGrrmmPiKzquiS8LEvz1mHv7McOBVW9/TY
Hmr7/GA7pzMsnTmlilLQ5mKrceLAzlmbgMhP/KLbq2fJ0tPthMWQyblI0OpBLMFd
jKZme4S66SzfOsTdQiM8ZAv7GQqFFb/Ks/15vPZXH0ZSrBox8RCTbm/nZs+jHKt6
KcaMMCfwB1SaxooQbb1sCQydUViqocxsjE2dETMAvKJNtZQbQaMlEJBy7C+xypeU
C6lTj+svuL8OdmHXLR819rx/1shl2Kl/awgWqDb2hqKa5zn/Dd8YxT/XbdTA0i2V
NyObjpDg2fbXa+600MZBe/zAXFiobIuY2yOFQ8opy9EBrbBpYjMx17nxzdQLkg5N
3PGwlIZb1Wkk+tY6fBaeKM/3cp0A8+sU6fltdu+2iV6yDSuJ2yJAcgnovFvJNW9Z
WbAReCb6B07g//GDp5vhDyOhJqsG3xfDMsYQTPd5uSMdufWlADYXQE75R8Z2nFzh
LUN+R45lMTqrZsZ9isKkHd1JBj3nyvb0wP9ioDwaqWTNuaxLbd0YWc9tlTynO8oK
Mpb+HnWgjR0dfNXDKFOcqR8TC3B5N7tt4lIVb/haRhWbpGZYdjmgrr5omtguX5lZ
9XBViWSX4jPLWr0Qoryu6LKi+S7CuceWzd0EE4uOvA0OUR4mwIzf0hLXIJcEjTiR
oOQqK1LiK3hY19Pxtj6cJkWpLobZvLUgZj/eEcZFI3tUL3dKEPF51vPW1e8M/tlC
HAhaFoD2lrVdgGZjfYrFutI66rYX/VQgF+tXiAD2ENHl1FjkqaFN82RDeK8XuE6D
iUIYDE08chU33va622nowve6y78Bz7ZjUqY+GvE/gtQ+l2bQFP9E3kS8OXsKBHdh
6JshZVC9jgpWqCiqeW1LnME+Dx++p86vjTV7zALojC+p30B5b9hS7LmD9ljxC1du
xnZnfFgTx6nzUpt98duuivelwHUdiar5Stj5tpg2L74JjQpfP2tzfmlroFzF9fEp
TbEPUWvzK7h1auiM8ZyOnSabo1dhW59ZTZbPJd+Yfu/78PCUhRs+RSmr9Q26e51Y
R2dVccrqGN3uY7b1ttTY/x85rK+lK0KA0PH80Y0lcMGCDu+4jeeIFkfGWY1EVZO/
oiVR4u1gO+ybU/ZHmfpxIq/0iC2Lxr0dXbVN7mFNxQjdd1+24j3y4q97ASNFaAIT
Xpwu2esG+5KFn6Ua8/T2C+xxPIWsy1WVj9dwMUdtgZOTNaxPVHaTTy87FGY3roPK
C3a5rQlcYizR/7W6VdoOATBvGunsW6OAENJLMXPFcrYnYPz4HSpwaZ90V8ZR3t8P
luet707eFWmuXXg47B9/vYesgDBhysIBrRxCbs7/cAaIQ4c4LWwWgo9am3omWhnl
xTHKChHWyZSUeZSLiC6UkM9KzqGMkpUR1PS+g/wAG/8ARwodoJlDnMftq33F5NMn
nv6sy/yjnQ7nKRRTeb9Yj8PEqD36UZzTeaLa+JJ3f9EyCElF1c+Jay7ONEgYdBXC
HtdcARhc/99I7mcN6pL4o6QZUqrAUp/X4XlZrPg2HgJFMwrD8Pjmf/KNPy9a5kpa
Q041XJZge64ZaZMJA58IDn5OQgwhI9RO9ppF6tM4FDiU5vykqA11MlLnoJt1KoeS
kM7MeYYK2LNSItYr258YKAV51EqbUjQZ9Lzo27RaNuLqnhMfeam9L3dMXiAuUOC9
pDPjaa31EgYXSiOEeDLcc6ZDCTsLjJuf1MSokffuxOL+IrFy2LySpY0gOoa/gNAA
SAMZn8jqhSP0j0BDn8ZBR9OGdgy4cKJK6Xt/OHYHnhJptvyezt4DxvBIEOvvZlA9
rlqQDhWuDiGG/w4oT0YdtNInoo/SAaD1jm4y/RLKoB5ehweV+HME9EKOV2cXdPGj
/+G0iu2aCVdgXElVCiY9jdC3lh0HeUGxlwkWWe9p1wec1db6Kl/t39i07IZKNbJ0
7MXuMYGtqyGG5+sZD6N0BcoYeKuim2bMEhOZhAB7Dnux5Z1hOdKcP0ie4uJX6rKA
48LKyTzKQDb3wW8xXoyRka6XRpuQkrRn6NsPV7FJR6UZfvl3FQ6eOaQWTcq/s19z
3NS8Iyvm2CGn/EkEkNIIydGvldI7+CXFqpSro10/8cyiekDcmi8x026uSYkLJH+N
jtzKQowkS6NjQk7Qv6YsHdykKYyEnpIz5/MAOF82kVcG5BLthze9ciytX+nP076w
2g4tUakAwzx0Uc675L5LDPAOVkckxPykav3QRz1KdaNVQT/wPuvLi0+kKzAOoHqu
8rY4FD9Ce+TyaNnqeWGyJP0ZtGRPWiMsrb+qPtkg6jjEfKiF0eElAyLtQntDzvHh
sU7iLPMVq7c52PpK3MIhppPjv/rvPmLqV8nSeg1OCzlHnBdeQv+BzZAAG8B90gZY
qVqiP42RDu0X4ZI3iSwrJvDA9rexpM6JAtpfdZl9JREV7eMgzos/ppyyybJMrYwX
WoSoORaOjWBzK09Aj6RbU/p+32bBUj000lbDHEnv+SaUCBLLEREOPMiznbug3QEe
yoRZh47kBglp5m9ImP8ptqQIi0Yinq/up/0l8L27WQmdZRy0ECK2IwDA1KB+SoYt
DIlrPdMJJCUDitdBkT+b9FOo9Xb20I39tPi8I5JyDJcolivcZ0EemSWD34fXdBHK
mICVCGoWhZ8s0Yu9zgF/zc/gl3tWgLiwRXHQSyV3tTBr/DSR4w0J6ERonLvbQoaX
Buuji4/iX6uWJmxOkqDnZ+bsdA3FJCq/9Y84ZdHcQVgvUx3oWIOVoF3br+LzQaSI
R9FlMEcudqqe3ECyNzipIMUKqdURwe5FRpB63yO/oQhwvhzd5Wblrb5e134h8DSC
1MEHIX5S1DPFaA5u2YK4wlY/1c0q7ObWMpI5U7jRtVCJkbSlkK8u7V0WjNyBIeN8
wodtppQ97xMiZ1Vmh7IXBycX1QOEmkqzxwsDNz/dcZRClKYoerBrQBABZLETEbHy
YaWfHNk3Nfv0whW3PNGjVEwsZZ4wOwZSKRUHtCfjc+ecyy5wdtjpWT17py2fGn9P
Oz5LiWud2PrAl37SKKX3CKzqhJAw2wBuQxQWVxgEhVWSWSUDkXpZ0YT9P8IwkD83
dWX3zlogu3TdsRKnIw2FViPnn0em4bnIiFbPbt3Wl3jq2jwHI/zNdGwRk2hgDx3l
8pTGn0z41aYocYbhTpvYTZ5TRUJpNMG8YtM0JJPHS/wa7GLIf0Oh4MHUyNqzqVM9
O3TsgpNzDlQ/LA1XnbsKr/ODVayxiwWFAogR5HxAL2ToSnfQ/c+mm/clNwGtaIOP
0UG8yKZeNevdMg8QBlprbWgv0yRhq8z8bVRZ2z0mozii0A6Y7DPgnZkE/WCmsgup
TDjR8znTgL85FDU/Id7PgHli0AqlIiwrcbpHLLRg/saIntvElBhCpHUkjlRA97Fs
C1FXl7D+wysqt3B36k5NpX1z81HTL7NikyTnRoOBq56btKdLStwP8o/tzQ9ySGjQ
y/k2eIkm9LHOAiFvY6QqdftkL3Ul4JCl6OmWypWaQ12Es+Rd3iG2Ini4Obi3DNSk
f54i4iyahBfYcxLB32XrJCnGCZznBScWY33RRi+pmQ690iVIwA+DNT2/S/t4vD1T
wxD2SK7Qvv07yeTzgU1OooMdiN7VDXHQoANUYn4YuUBgmueQip0cfOWcliqWmI6A
UwnIs0yrbKRi9jdStmvDQkLgsvPuL8tc26FBtPxSLdB4AVj6OkZCyPUnnsjs7Cup
I0KkpPkCPvC8MAz7mh7HaJTcv2tZZZYXXff4IgP8gK5vUIJRmcibwwCQNjKjl3dF
/+zEfe95LVqAkA5+nMuE7L2SiLSD65LWQ59BSck0KqfvqsGbrTBYqSVPsMB/JGFX
bboAm1dA5t0FWSYcIpgvqpevwYD2cFveMb0PnmZxMMUjblGtuOfnaCynpklVXytH
d1T/kIBsALPQKmOB7rPHRkEfe5xpZxR+d6WcHEBdVyQ3ye6A43TKkNV4AC1NOGau
31ZzTucHAZ4N4riajR3nLkXazV4vmWaa+iDxRdeTybZeaXU2KAjtlU3tni5Ob5o+
HnQ9u9PmQd4kEYAOFvEwCpQ/tjoVpceMYuc2NvO/FsSVhYHmzVRGdD/D0hXzJ2Lf
NIRz367ol1MoJ4g09EaH4opi9Bo0JaeeRho43WOMGl/XBt1Yp2D4kAW8Kz4Ud4g+
V6r2QfsaaWywQnEBzMZNlyZVnik4F6TNCdjZck4YdQGYX9G5aN+ZABnYj0CCIzsN
q4vR/SFf2j/ii1fmQTablau8uhi1+5G14bFI/shSyGbtK9vTuvsvLoKzyalN/C9z
jBCzTI8kiGp3dp0X3eFhHbP8PUa0H7QZxmmI57rq3PwZh/qEz4C32VKTJHpDjnY7
+HfR07JfnH+oNGXIsqNYLA9fRdldI7LHpe584lFxX2rvSBuWRFwOK26xdeOYDYwM
BUZhiP3ouuxCvtNLBB4OokcveulCLg9rT6Vnp7zK45nSc86A8DJPIvPScd4uwMiU
dvlv1OpvqUy7VCxP0gVswDSaHOW4dIAZ40JMANW1wZarxG+OoxMv370j4xoc6eC7
XJUKY9e7MambV8JjfU3djiou+aIreUng8BCZIrbp1Ysty3Ayy7RFMX4XGkMckipk
4vkb5ANYASkIRhe611TPRoUXti+sfaxlLya3xf23ZzesB4LQX3BYnAYLFO5DqvQr
lLfA7YUCXq06Hjvd2jXIvwGw3ZMLxQSiz/sPXJCWGNB8TaPuWwbAO1lZRoXkutGF
GyBygN1mPNzAFG6wLa1tNjrhs1HcrPWBKPnBslLrXvHDMYJt7tVLAbBFdGMkbtru
FSkAuq4+qjm77E4fyVsWl3SRECgI7HUVbqK4sJ2yFJ13IzMbpHLVRq63SN8V/a37
eHx5WHpbhvSfkP5F9kHmlng1ac89sKKGsyJZ8zucetXBYSprQJiN1EutkFPtKpxk
EfmPGF5qCs49DwtJA2083oRjVdJAgYK34jAQZkPoiW0cqKplzug5gbgDx2aGLk6d
yr2zlAMjCqWSf8YD8fj6gLSBdCmEL1hdaLcGyzmNkAfSlEOnVDy3gvQbfEY7vtQK
bWc1MWyJHhwk1wIrttulkwlqXfBAFxbJcZc8i0pK7q0XBWljARKLqJsi+MbM/pkM
qWpkPQVHnmsPHmVuIMxN8cMR2kJ9CWfE6JoAp4unLW2ioLiIDfDCqe15szHFkI0K
uXKGgtkPdFMDzihAeV8e1o5rVoatItUanAy3PJn2osaGRQXeeFJ/NKN4j8bjiXUX
3mhWVVdpfowPzHwmUd1IBDIXAWeRF/BpH3AL+I2WY9TiF3yzAZsNhEEpJE8fmigf
Sa0BuCZlG/KLYrjywpfn5lEPojS/d+taVS9pi7Aypl2M3md60wjY+hRD/OUcmqO1
omkgwa3HMcVujEbuLdN//wBFtzS0goGyovwEHXR+E8mOE9HVAHAX4gyArQ+A/n0u
wpEp2DZLJwUouDoI4dG03Ded6TyyFSCeA5vks7SZ3uTrmdhM3AaFlXNgTQop+Yvi
EUVH+DbDvaAWrz/an1uUwv0pP1vu/jgo5QHFs/yG1SXzz8+g5PrmoZMNbh0qKqlh
lUUllQUEsRwXXI+2oxkFvesMjMTCTP+UHeJ/THNhZK6MAbH4joz9EX15BqGF6661
gKghtrUbQtulJ1EnqEsWNxk48SeYYYWU6TKkcvLep9Mxtq9Jd45/LWUv2MggdpDg
pcJ9Wl39AcbXyyMN5HVaul3+QzVASG3boRw4cSeSj5x7sGosotQZNFMYel7y9zmA
ECJLep+auKzvC/SBbbm7d+TTmUshhx+7oZ/gxED96mwq8jp4I5o7MzlDS0klnbcA
1vTQ7FIHjQJQI7EOQzIQd32sz80hmzxamA0fReK2kH34egNj/24qZgoXISh93Vct
c9zyWRadFD42BSnyvTWvLyjJ9PAVASna14RNXKRR2tHarDZ5z6CFnubAVR2k038m
bGVa1no+W4E8lXj4GZuGTs27H7vmCQLuloaZyLm0eTqGF5C49/s2ZQItckZSvgtL
2jvJ2xcLpLErc5NXNjhOYysK33FclN5vomz84RSDujh6HYLK64oChXnPSbHGz2N7
nhVyr7XqNmkBSYPxY/nwCRORHdHxokvSyTxB59KDoD2EfAjqdmOrFidpYxtV5dG7
s/mfSPq9nl7ptOaQkVG2KDUQph3l2odOOuHULCCrQfMMh7wM89wV/BR7ZMEq3ToE
fENGwDHGTHNqrAmN6/CY7Kwb2rymEhIcIB86JttRPm1zPZjv6etr0ucu1lIZVFQd
KXNm9+Hc/Y6MLBYBiiLan0QsJ9x0SSPI3t25xNUk64KEgVZZXSqqWIAwH4p2m2Cl
maSTKw0ogwBg+7n4TzNPW2F8B2cquW+A5xrj8LzZRSaACntbyL24in1pOyW+wyLv
Wz9WVVqaMNCLqGGsyYKAgyT/rdQH/O+UXWjjj4xQWKY2sXkv+ehHW1lKmYKW62Po
wYfAIjW06zIjaI8/afRqKaor3wByG5kxsHipFfuILoGHcT3TykYjTu98jdjfbBWv
em2fdlI9j0sxBOXNmOS/JNBz6wxvBvq0qL3axs1XQu1Tb6EJUSyDrfQKvuAdPjmt
sqp88JanikWnxcDYzztCBgs248aYB0Gw+LdmOw9Ohb9gwrl8WsYK9k9JbZ2dERuU
EaT2TEN1i2VSnknlA/woN04YxqIJA1rmKCfMubxSaTzCGq2TIH22dfCXKoDgkdaN
MnWaCuNgyHNRkkrKHT/iL+PPwV2KZFxuJr26wqJpZ1RlFFBx4ZH/Z+sm68A/ikN4
uKTUhkHqa7RbLfqZPd6ojdBMLb4AoNPV/lOaKRGn1AaAnfNvO4V7zr2NTgvCkDWF
7S3T3x+JmDId3Sm3XdLOPRIBfwcOk14J/+k/SF5F3Dt7NniHTuP6VvKgVkdjhPGW
+yWsEJFB7X2H3JmEfp78bRob+iNYV4dmoPSZAMj5T/NPT+8RVX5Zk7crcr343XX4
9eNGQvwos0H1OaqwPxHSoVqRNq95UpgT/yS3qzos6HyQbRdJyGOyK0vSpEc2P+kc
af1Wwgp7FhH6lznvKPg9IkNoR2yGYyhY2oBr4razisUHaBhwb2JaXHICgr3Hp4qZ
Q+5jZJRYb3Qyk8AoKFP2l+I2KkCcl8OrU4lfcVXo3G7ol7ZNtO8TuJTf5uezlprg
KVH+kjHsAF8nGTv1sRIqk9D9wLGCrBrPgsDbFZAhQAU/sTcg4EeojjxIiRY1sHZ3
VVHIPM4SG2L/6PzJTHEWZiPvXPaM3y1mMFsg5Y7DtM12536fxMrc7StUFSJRSsce
Blr/6IukJ/gX++W5Pze0HfJaGnVIWr/d4/QuYci/kzIYmTK8yTvhIX0a1LaSVQWb
pNjhweEsxPJWCbl9E3v+LSCQkBiTMhoqcGnuiC6sz/xcrP+fzKDU8/os4ZqGwpLU
6eOOXZ7ecf8QOosAsS0zE4m8RErUUsEZcc/YRPVdObz1lHXaehUqgxnIHBxswSIb
vqyQ3gQF60wnBygecQTARIu71bZTDTrYcPR0BbZI9wbJU6GURraCEtKS6C30wFYu
OYbXKF1oHw6FJPHZR7gZ9Tb1DtlliMDmt9TXnApK8He958LzVRdDS8Oi/tY0cwsO
R97THUggrePzwT+PJnJZ37QgusnxkR+PjlXgETSfHeAlZXkiFcxVTi4HU28TZw8m
E9ez5zQ6JN8oceEPXn8ODWL4zNmftJLXZhitnWIimaXN9eVVN8FQjAyP/hhjE3ZK
EZ9RduKRCWc5NY+l/Z7fGLU2Z3hLCrotBGR3amjdKDdyuLuHjMp3qaRMrbcsYP6K
5AGF0M58G5T+UHhioSI2qk7DraQISQR5IBakPitvdVx34j6DRtX8FO+rhLLKIYSI
XjjgSJk2d4XeYR30yYIXrcNkvccob94jBVOLUPCVV7B3iRLzQPPX3M0SGBnq9D4h
bXdFdaNUuXmY3B5Ju84qpNyYnQpzPMl98xO/sC34IIlgOiUIeFTjnzPCLstr7jg2
tCOVg0HNMfd6u3g+GbrkL0prXes/0Z0uVLYEDERjov0PXU9fhgg76RMzGgTofHq2
P2hVlHRI+d65uu3A0MGH4hLPrC60UYtgFi4EBoZYE2StKa9/44MXPVTS/ia2bWCB
QK0tIV02/M1vg849TxHKfAhHcKVhV1Y85TzTWvvWUQqJHGX4j6u03c0GInwudS+6
MhkI4p0YuheWbhR1G/OX7Ged4Wc0/w0UmJbBDYp0FcsVXqoZgji+5MQ7tJLPesDN
GYJr7X+g6+vWIDzfFPrUEJApRgPKBqDVUVIwlLzYSf5b3jnJ0zefVUsMp5A71lpz
3OvGZHQQjgIuPQ2ei4vzrcKRz7IlvPmq+ENNENjz7ZDyU6jF3tTK1P6sljed6oit
XDjqyGIdqYV38ck10nIBMuo3xIewz8QS1/3URvqN60RnJK7wNcCxYKVoz1rgb4By
1p1xjrbKz2mcPew7dTfXjViPtVf/aVwi7wTjnJU4aRSn2JSPqCO2HytrDnWD9+AC
LIqm/2to9LvN9HerV++gBBKPY6J3v2f9FfLaB3lg8Ade1RwmHXFoBqFnk6WIS6wi
RmqsfHdoVXW1nG5ZU8YXAQ7Zcq9wDwn7lLVLGIMsx35lOq/uSZcJfyvVV9KJD5iV
MM7VpoOxad2cnCqjQefbL2pUcYj+t3Kpa4jIgzxBnJMVuFFqIJCg+Da9ov1P5S0C
kvAmTYH/zwtQm+wUX9+UwQLRuCBprT/Yw0jy5gcUE3J4Ejn0l/qm2nYx0auL6aNl
ifvDoKOnzbuCuVumMBrhBTsDNtBqdH7goUqRyqqIZOO4LZCAMwoJ0kdahvVohAX+
Y9ALttZ4+oi05LTFk+cxRytxyk0+p1qqTt2S5p2unCqPm20PAtTDlBts3zlVopBC
48WACcBvQbnpWxULdZyokDkILM7jrLdaUaOS90XSUsJDwPunlp/bHdJEcoGHnMxY
HSwHmuLKtx4xw9ik6ZAKxb4cxTgDUvyOcXpQWSa2ga8rpy8unOucst+8iFAuNMg8
nYxT7GFc875s1o1EuUCTBl5ZumhKkZsKuSkA/sl37ZrVkd+h/Z8GjiGobnBpA417
6adEQuMs6N+myqMLAsH3VyXPHIywFN84O5Jo4OVJnpGQP9zbH1EhwMXuaJ/7vhfU
0nzYeW+mzknXBtt0njOhEs55tUoyZYGYxwFdSwY9TRXllwS5eVlRPts9D3kcu/rz
wPzY6deTc/ULfNTJockJkxCLmskjBycP+qMcJTgxaDdTAZdisSCmkQpeDZVFWx8T
79XfW4W4UkCDL9nNs085zAHMWXYOEfgwfI19qu9IZhAD1lbBh28OzR6ks7Wk/Cqw
FYUo2epW1m1iz0b7rH0X0IZnb+5XZpLEtNAw/uOaWBNxJdBhDjH/y4T9nH6n42Aj
ytzKZ0KUePUuvOuAT255qNI6qRShUas3AIVIIQwXDkXQrulwiNL4o9MJ2uvC4nTf
r64BYFPsT0Ax80EzMm4jVU8CDep8k3rl2EQgCxAU0n8h6qRDfq2WGTLxCQiCWCS4
u57FOz9cgbc7+ycGF+hO/ysQjqNbk/bBVJEC0N+xLgNajWbtdJP35ekTVRjpa8b0
sZP1HOxDWh/Igy2mqtRK1QqqNMnmdSlLq8nRIRZ0YUYFTg5nKIwRd5WTRdxdObYB
6au0C2fAMiYXydk7V9btkfYx3BpA6aC4r8RoUA8JoIPG0tJkVq4eUv/rWFFuK0mC
SF01+Py8CiyiRXu/F7fZJsSufJf032f5qFikXtM/I6WjX4R+PQiQsXFWvDjmnGXh
jD+MwjhECbFxf7w03EzA593L3qgFQZzKbJ4KuXW1nXu8jUORDTZeXSzmmkAwOpfo
1/G9BSmtU1y9y8sVXfEKRGgGyS5puIkG11yAvX3+748UkL3C2n0t1D1lADQf07Hk
dE++XjpCk5sD4Qp0p7Iq7YKDx1mjp5XemykDWGzUgdxebDxmRWN46O6zZZjsTVKe
LPOmZzvMwJ9CDpP6o2p+phF6CE/LO5kF8lPImsPzzXYZj7DNmpw9w7RYMQ8z80Pq
5ZuZhZ3evBobxtHLsSfa6e3kLkmZVtrStjtTz2m3N5LJ74LYKP+YrkRkJP5lBD7k
wBfOrYlu02TJpGu8hU22fiCE+hIAxWF6VY++8yIKE/ImJVEgHs5bESkAbHmwnH3w
lbdgweFlEjkZ1HSu7NmJ0AzNnYYIJriNKbQXDUkrDaS1lpz7PrV+1taH1Fv0xjPP
n9e2BZQUw2Sp5n9s6esY9YMKCqKwPCE3qbEgqZjI8RdzQFAG+N5Gz6Ma0xqMBAAN
Z+TKv3BzuhCH4MWr4CB3KMaYWdZEOgm7+hWDkD1eJr8MeDqppfFFHnOHeEMeSNoC
ukpUrfjEb4hJLTbl6ga3g+ATaqIyQAzsb6k552uLanlCcTQfNI1neEcUn53zm7kq
YjJD1QgrTdgdNEWjHuMWx9Nwg+9RPSCcFymotrVjEW+s9gKJUJ9sI/Q5tkRgrTp8
wAVTAT05fZ+AwUcHpNWusOmQ+3JbbUO0+IYxzQurjgRGTT+U2IH0DAHXV32+uzWm
FKE9KVlh6Q1SIykzFfqf6NrgDaDmPbgdn6BjiXJTNGIIjXW3RlVOGZ7OXa/VQ3or
8msWtyfKzAK0/XBwXAu9ji6/6QBAabLpuusbPY4hpnj1V693/3wLd3NPl7zdtKQ5
7cBD+WNp7gzhL/leuqpNCG0e7UpkVU8x8C53NgrIpdwOGJIqD1LtHNoq8tYh6+56
Cedcrq02Ju2b6+udba3su1lXVqFlX8RzK10IMn+Xp35OrxjI5fZvuMxR99cmugQZ
RFZrHkxaLwAh5G5Be0WFPEH1gpRpUE8PdPl/RTf9TTiCtC4pRuY8CqGLdlv7GCDx
EdqSb4IBrmjrl2l4Zk4rQX5c4AjvwHwQPX5AmteACZ0DEw7RGQbAmu9HghuuDMXZ
HTurtF37A5ixrHy9fDsx2/VfwyyYQLo3zW79rnApWkSkXHJQ3AFg35e94PhhdfKV
dPz1AVgPJwqMn4/YA3IWHIh50oMhWsMTQ8ROL907o44VQLWMAkI8JAluM+DYrPU3
1Xh7LZkK067dKi8LFckrMkps5B6r6t/ZdclVHeQ0Fpj0/3Kic4F8KN39QPxDdSI+
56fWBuMLFmaDdtVl/27hbwv6jedRfwLdMGgPCtosuoV006AUb3WmdLF89IVzWIpq
kx5OxGupTZs+wEsZqCOQdjYxIdbLAaBy4GTrLaseR7Gm/bTX/m0EOON7ykfAaT2t
7cvktK32bsWclH3YKN0g0kRXmWF4V6ar+5w8IVSxYMkjATAjBrJ2T0FqVzFRyvyC
C45y/GnRE3wkEH7462j/xguA+M6yP5Ee96K6anePEzXIlSRVmVqXnn2giU/USbTr
7BbpoXI8MViXVZb+bAL7iaiU0EA4f+BvFNoeHPRBDV/UTt4exfb1zQgvSyxCYCep
fboJ2SDlNvvL4PcddfiUeiCYpkfgLbbreWFkppAEDi3A50q8e3M9P9tWpUNwujKG
LGDVuVbpaEl9EoS704fbahtcKzurCYZtqtsclpB4jiTEeshpkhajkf+7OFPo/9vY
RMc7xYQy4ppnC3qPbGYA1l9QqbczaaFX2ZTgeM5blIzRUmEJSOqtt8rzX6heP9tz
o5yG1Bjl4/CwMQO8WjDX32vhet/45zI6wgJjED3+DpWYLc1hOsmSrCeK4T74EE7A
d2j3PJrmktQd+oSwLDSo/S2IcvDFlV9aKfuKziC2eVbXO3szUPbsMLi6T/cxwUmp
QD6orEBJyqursKlDh6v5PfjE4qAZlAblGLCS5K9lFXm5q4JeFhMoS6M7vDDcS1qc
zDjxEhqeb9737tfVynLccfWupwe08lmgSUd6fzEvSmTNmVOSzVAN9hdcZMtvi3Hs
qpotKhMqsGI4bRxro9Nopg89r3lBq3ZKp+W/udoyTd8P2MMDu/9JL+/vRd/HNZiV
S91VT4v0qDwhpfQQ8Jdz8PfoEdv1oDcum7wzGlg/09r7IqGc6+QMplhJJbvoNYsP
y45MgOTUoKwKUD/nDfCQ+ZJworc2ewWGe56OFjv8cQkugmohRROH7emnw5V6Isne
deY5S6iQaiYF+UnJvYHK2tccE15EOLxWeMzjKSnjrp0pr9anmWevrsMqfFEFprNu
ZiJiy3bmKAQENFy1s3KidbSZmijb+1jss3fcmiC6cxIqVRYPE5QgL+B3I7PyroQB
40o50i5SrRHZY4iZC18J2LRTeO4yEV8U9sMyAytwU4C4gxBx5GRSC3Oa1WW/UYCa
Qx8eOJm3xec5S3g2Uz/Pt6hrPCZGrOAsQ/3q9Kzs04OeN2RJJyhdJvh9TJ3DzDCT
jYsn/wRBEjMjXbIhBjUHWRZaccAXFUxLa/D4v8iVoC/hBdsScE4mYaE2Lk56AduV
GIMRj0vuEFfPjf3V1Sxtvn5LrUyfGgsDe2YWHI0nYK2w3LEyCjUyhq2RkOVC4DTD
VDfGABeisA3vsKtTzqQAnQdY8WyvgUQSwHgywgjxosGr3g8CJwyXEhd5AroNTnfP
45drOkY81Ifq1BhAgongjaplsRzjACumbgKGGDPV5N6oS1Mvs/YIntrZKAX1kJuh
3Dn0nCjp4sLaIahzt4++j71bm++3BTVyW7PkOrgl7FBb1WK/bps2c+z78QD8kWBO
irZCDU1yyZON5sxxy4IcMRbKOhK/NeVpuMGbr58qwU+G+HT7HapNRig5hP379re7
1LCv8LrfP7zc/uvGeAY5/IUf6EQj+Fc324Uaz2jDujp0gihBgWDUSc78qxdccJPe
4UvSXP6Aju4yWUvyB/cHKbFCM1Ee6q/4kFLNSlm6Abm0QE74Wio6eHGK5aBbyawp
ZO0k4TZtN9hxLqyuiRgXMu1OnDqOItIF9VldEs86GbFh8PIuM9QehwQVuj54ZCKj
el1jAQ0RQxU2976g2lF/vZuT91Qy78BDJykA6+nmvtJIg4UgUR9bKfWVVbP+CM9t
qhIjHvI9C65UzRGiI0/iuQFsUY+M2kz7daX4kIOcsghC3DN+CGpGCmY3sNe9kvQC
KjImBTTZvpSYPwr9o0zTEGDWpDy0vLQp+Up+lKJCFCaxxXD9/f6JiKFR7EIVfHAZ
iFvsR0WdiiRS2olhaI/eXL6Mr+Xld2gncgewBMUfwKJUNsoHSietMTaLmMCHJazn
B6VKRbaaH4qeRekFu3qDGzT2MFFbt/Fsabira7troe4woKR4M/t45PGcK+G/cPo1
reVOK3xlUZrRcFy88G6YyZJ3/RkyXV8rNfmXbsfoTPd/pswSp2Gtl/xHeMBiQHNV
zfqVCVBEN2AuwqQUmV3aW9WuZc1r586B5KcCB04UbrzDfd5Av+8Xdiy15taQgqzT
TLgT2lT5fGB1YO7QJjKSxORl6Cw9zKx6BUcyj3hYHrrCHFSjfRwHbmCdLo7PsTVS
Sj9Uu4gAfG1+7P5SSFV6Y14PfpHaNYLcNuHDgmHDAp1vopMMdWmQNgYMgkPxSYH5
f1CH8JUDc2UfOmVuTlbA2h0b2l6eiuCyFkbh7VAN/GpFmS0jzv8nQlrDIJmL1JH1
7jDTR6pOJHTJZFcoY0+TNdSBY3wPCTAf3D/wJlF/uKkPtg6VKCUkpjSxvN6rTEvr
QkR241OQxtOXrp+oBGKtIMi6Coj+u6tJXfYcWSM97ANOxgXZ+g5uRPRQCCeAlDs+
/KU0BHw1HA3tCtbKGqf3JMF9IE96W8VxzPC+nL85fbGQyBWrV8ka+LM89KmXztuw
LAhHfQZS4TVXVNLwwfXVfpwnimTxxmb3WZpoLo0+fyfH7KSNKfFy4ZDH5Miir2x/
MUAK2CqrIK5S3ohwbiADiVZErzQ0+q8Ixopx3ubrDnKboerSGlM2UU0ICmH1uTB/
NyKAjqj2/f+myzNAsNxeENwtyVoEXBJhWefQNPx5C3vB1yghSM9ZeEDgzUIqPU09
9lSCJ7J/+lf7idBhHyUDbupW4bPKXNsAheIB660Tcvhkq8pGb/Z37KTRyKwQYBgP
Xmy6ODAEOzGhza+ih5JLK00in0S/63WUFlw1I5pVpC2PtgIpiShvHBGPleK+zKmo
4QVNLxWKgFuG+dLG1kMKWYQT8QXtmoMSCEx7mQj+bQcsbwrmziHpVOrlguNXflSz
LnYr1QexRTLpa6Wzta15NiEvqfGG3DBRqazIJzSjJmqU3Z9qnz8cF33vdruEybwx
Qg5gQegjXCNAv5TwNMluj+ur+ZJqzICv3e5xvt+jJZ78FkjXCCxr9dmn0vNphFPp
penT2ZOaXhRqMnnPi+7lmvwvHT1rhX0Sm1BbK2UEPNfj7Ziz5cIixN5bqJWbpXg6
gnP13fNYqLr3tekh9Cl4Ps1A2SCFnKU2+KYjJHK99T3WSk2GttHRQkJfieF9VS7o
t/Hmuq4oFXWnGMMIsTSKL5wh+A9hSxhOk9cwpfnNQqINnKWA6UKJ+cxRzCJ8mb9u
LI6fbELDNyMAIpkKwhA9mdZWoeiiIrSKUJKenRuevNHhUfvRLHxruCKbre7jdWTA
1Fq6RDiUBFMEowXGnB2TRrmga4Ly2x2Y8ZCXHqydPC/ye9vx5VqYN2xzmGzAsW+E
x77A4REe4S2h2IuUCnnVn99J8tjoaVjeWdy9BYNWbBsXG+jyM3IQzZPXYE5vmbkX
xW36pjtiHhwrZrQmIiZX/+jyWPrrHGHsyupL1qM74LexWbp9xCKurKDNsC/WMSSz
SwO1jpPNURi49VycC/OvdkOciAVAtOs7/nwh/ZMbItqTyhh7mYYOCu+96mSYPi7F
NSShJ0uzrd2X2z/uGSfHmFh+zyRf63NILy0JIryRXj8f4jORDKRSsAlJZS1Fd4DY
DF/+kdLTFq46b06uNFfdZCmOD1DBF7BQAWfaji0UPgR+1KJOV34vLsSuImaujVEk
ee33rdA/qL6LRtV/qvM+76FF+o7De4nLqtDMQLKW8Ratg0UWfbut6LVNlE3pPYpS
2McYZKgt9wIu9ngwJEYsKzSUHsJN0WB2MWwYVNQmAC2AEXbPBOMX4EdC/7JC1XZ5
4aHgn+mz3OeaiQZe28Srk2/9O9kxa80gYZZJWweUTcqGZtSzGunoVJcHypb7ievK
HbGY/Ud5HII4nV/UTjxTHV4Bgw3JhRjULL57+H7ac8rV+deBbi4nYLmBSzfho/Y3
ExSF/S6ysvUmAFruAo+K5jAgqmUbufKyiM5shTcbrGcLtxVdYpzNrMPYW5wzBA4W
rnDiCJEN9YwEGJKBbNgGFgJut96FpmtU0ZrZ18pKuWlrX9nSj/uBPywdS4t1ZZ8M
9x7guKhxa/OJyzYvK1ESDgANwi5YYjIExNcaK3wAqlQfXUvOi6QFaMRdYRRr4nDg
EBw/ZpM0Guxa662AR0gcwTulZS0rz1hm+ThRmZkBRrxyOT5Gsxpg4GpS41l25tMm
oJtC0169T/+VCG66JcRORGMOo1xSCD3AALAFnuFU5ffF6hLSHxoJ3hd6UnbeSbLD
t0bWlqAGK6D34SXSDtHO2GSCb+GUUpBPFW+p2x5f4KDCEMh0vU5Sb9eaOecFPnzS
KxV/BoaQboeNOli2RSBzeZ5lzvkK51mQCzb5i4I76otBuiGqy6R1QczfQxqKhg9P
ybmomR2Ef2gZeCd6bJvFZX6IWgoqoGLmITRCdsbxVVvbk4me3PaCRnDU7jahnAjb
i8jRZKFbnzW4R1u2/k2bUqHqwZXHRm8RjXFBb4mqG3Pdd/fqUSItXO3+vyysBuIB
mP2UzGFIQDXlxevp8rY20WE0C2Gljt5WuuJi3crWqbTmW6QaRWClWxfD/bbkLOgM
fUuH8kJrmJJij4kZWaYErKjT9Yk78bHfBNxFUyIOIbW09dkOnKCtyLFKD1LCfsLF
6gTs0ICZIT/BCbb+myVpVRCiD49RegCOTCuwuXwptRNeeEP3EeArNAAI5nqTZJJc
lBKUmzNoyN6aDJ9JvO7bZfBWi3t2LNWnELshnjrszAH2en7KKatFiZH1hFDShLjX
H4CkIc+UJXbDgvJns0k7TMDhMqkz4zPf/U/o915O+S01iFxCRraiEa/gaZVLYGYP
8K8vUmBaLY5hRwtlMhepTeOqi5k0tiW8mwXc/AGgs9beWCsmrMFOEGxzs6wFVOaB
tqHLg6Z7R9fACnxuL0kihqu6K8g8Vuu/TWw8expRByLTMFbLiBlExUTSxWoeriGU
T8imjvhBLZcjZ866t7krcCJ9XKDJkgNQWt5bbfYocwEs4k3ex1mrvmhOnBsmUtfd
R8UJ4cvEBOlkksYKsCNAP4dcRzqvlPszU+Y/nnjR3wKzmwN8yQy6st12caX9bBr1
qMLXmnNt8xc1MzucKrBuj3rVX1rwlLwZzIVzQAgpx++laj3dlptrjpE4M7vK6uhW
zxt7+g0qFMohOM5r4vL5qjmnuwpaMZwmghTOJceZZKTjortSfVsiGw0I83cNWfyn
QmhImKxf0K9L4cymBH3DmW03paLpz0JOQZLj6d/i9XeRXM27SI47XTt1FPHmx+Bx
CbiSQrrUyW75bmgZOA8HI/dAuKSXssUqlQfuQ3q2piZPhRngR7KwHOPGi3gdAMwz
5d4MKkyY3XXBjGqgAtARZ6GhAB08mcdYBbzfNie2k40HrdxKe9QhUHbaAe/xMywz
9v+ck19tqKxrelMhS8CFlli1K/zBPdYoiHTAqKT83fGKvoUFQpy6nzOobDS5W4Bt
gfUtZi+dHM9eej6/VrZ2GTE8m79w8dH9priJoQB5tto4BQ+oO0gU9zxwAO0dmenv
t/iyWEX8dwMKRI6w4qaj1Dn04yjYUh+L5iRuPSAUSBTGPZlByaRJda57EYMvEcLn
o2me7xti8g0eqGxhrQHDAELjruM6yPN5BGREW3jXHU8UjXLN/EfKVjsBjSjHP5Jr
rnAdDZoi5flTa3XrKWAERNnPx8+MOOeZoj0YvSHK6FRRuU8NnmbqWpa+bAVXAwF/
oypLFNR5w33yJFHyJvm73xqw6YI9G3gW2dbzp3clQOIuJJXm+1BXPo/dkxruYExl
/gF+55vXvg9a+tzSXwOg1VqXmr6vxEqSHoUnuc0Tg86nSD2kGbJUwQc0BnohVG7X
fJepdlQMaElB2KGiPNFIOOqQs6laSIVf97NjBt342DWXAUzvSYUhqVkbncvVf5Cy
6a4YzE8QY486AgNadDzctcvyQPcYB890K83d02efvSuCXV0IbuWDwCGPXl9yTyej
zKMmptSpPC62RVlQlyl0dNZ9qEEAF86RdPMQ+F7uSbdMT6Wft9Mdt6hoHTtw8jv5
3FlehTvUADRE7vQfHwNfYCx+6gEKqB01gmisaiaeoY48Tu7Gv0r8+ptrdWBhA+gN
Nn8k5QXgpcqOZ+Q8mSmispseNaJ+4C4cfSKSNpokxhpLhXxLiudYVQ4OMZmIfAVr
sikk2bCt/PlwoP2MLIQQcL8SA8P9Vp8pwXUrttuQfoSKxbS3JyZ3gLpA2H55Vgvg
Qes4mLn5+aswgM7QcK/yFMy4GHbAqfSLi/p+6p8EhaLCk7ATJV77nclSuyV1JiAY
hh/tqz6mLpeaY7wkgrz1w+pItg352o9aswl4HYV4chPnRKV0LEgG57wDa3fZ9JRw
fKd94z1cq2MgDpT0ido7ze5k/RzLvVpNQ7ft+Z1fRATrGvNm1o4lxoW5MNEQjEXm
v2TNDFJS9Nv2iu7niKxPOwkVpaQBwIkxkNPLG6UIlgWoHwxfuUkERxlzNg0hDlpy
Cny0UI3LYAZUcuUwWB2p+GNL+7tKGuHgNzEUQzp+O/otV5x98DCdqKr3QD7R091T
LkPqaehHiuEX7slqea5ZsN44oK588CgOM6UVI9Mc/msXYJvdBaoknsI/QlKKrEvy
KZV0g7C1xr2FHSVOfUcAQyLvbuIJxSFmDpNhmwLdu6QzNE+OAJ8WXpGyVnoEXTIQ
f07HBufoGuBkt/n4HftIH5IxaCxKHfXo/WdnXFKiFUcDokSWoE8FgJ/lqibEcBIA
pid+RXX2CrGsX3pLlv2SS05gI44VfoUEdH06A7z2WdB0WPlOREUuxJ1Jro4go5I9
LMQLGWGlwRUI8i9qqBD/nrj70zAC2f5sDSPOb4WA7PbXpOpkIynv6AzZlJt5fXVG
TQ8dWWhzPqIIYPEWfdnWDMBXaRY7Z4uZZyUs4R6ctebJxzcAC5Wfka3jJWnxWI44
1ucO5HSIXITVlLktI9q+NHB0/PaiUgET8GKY7gkGAyCraYjBsNptfEYFxMVDuZ7M
UiLUeAiBMZG8UGE1glVzFelxpsHNelEnDrMe1r8R1xBG4q8JHYpdR+V6z18DSBLU
o/tsHGSaAnotzQwAOhhd1HMyMhoxJzUvCZSEdbbhHsqRea2B3wDOwXb7soCdCbBQ
57HLHD3/00Cfc93vnceWK2roPopP3vSVZv7tK3U3fMDOs6TvsYwP7p+yYHSWl4wH
weWtkOUFtGU7NgfEAXFnI/hAwtLhygyxXGupi3EBkbXfaoNLxTxhjXYYGp1lqIcF
Nt5ZU85gST7/neTgfumSfyDgMPX6dIpk0dB1Xd4bJfZDQPI5vOqzhI2BdWnH/ROU
EcTzC5f+wjmGruaU66BnutM3pcOYgv9jrLuDkqKo8FdKANuKWpsXUFnlcviENkxB
hnPAlAZKVgfTE/+ckpkDoYuVfL/Sy6a2VzMH9SUY11HlChHG96t7GMM43Vnf6tUO
ajmYUsHf82nZmqbQ7cUSoswu/hyt01EXBCvHPVRZX34/ocEpjm4JqumXhgRRGpb4
j2UeeyIatKD5JJEXDbMSFVwipASH7ZvaDwx5KnnDQvWRIWwhyd3Uo1qM6LFMxbdw
kOxypKCUahUuXJy9C47L6TP4gVv/DLVqPZVe3NTLJ2dC6vylN/nI9/pwRxSY0PWC
9dZNMobUVMxPkjVwDC3FDrTNIo9z5n5ZfBCwmlbmzOWnWx/TXU0yd0ocLMpHTfKQ
HVRVCo0sEjWHZJRAEclBlS9zXNk336hMmgHPNHlxn5UEd9sVVyjuJcyxG/M1B5WF
eul66DDTbEFf/UX5s35djnhPH/SiJ8nIUYEtcNMB2wRtepgsomPL6g21LKNcMK1P
fadmgQfk9KgYzUjHs6hsUVMaqQDWAbFJl+J7bDCJG4RBwIHsrZDOSBy3hvC+IQTu
yTOZlw4mHAHLHpNVxGQKGo+8ERKqTK5jlr5QU/w2U94gete4wDCCBfUln4kb6D/q
p8oLAYV0HfZl80tO317wDBuNrP7JDDJN0j2EQ4onCFWgPzz5b7iMtPavtoGIq7I0
Em6wofHkVib65ssdrpKl8GU8RyIEAPpARVCTDZ6jyA7ZRBNxKmaPE7b+hVG+kNUH
KkqXWPDHAVgRTn/AeyLyL/H/0S1gE3GOc1Y9/h60ae74KGPgxjz3exyjRdMY3SnW
+gZrVTDAihR29lp7RG7CCK2IBpSWUbdzrjzB5rLiu1WsBLTuFOAA+4uGCYgPQMVa
Lu85cDkrWQqzT4BK6K4WXNWYscvu085sgEnrQ515Yg8LyIwhY0oqkkQUXftyQ6yd
zqUD66lMIPQCWSxvt2v0iQAMzlKFPzDTDWOPDuegFVvUQgV2qk4YaWygp+5BGBDB
zVHeOTqjYrIsJaXHe76eyjJSdd7ZsvfivNg3ds5nLdaQlJ9ZlYXHprtaARmgc5Ez
o2K/aoGJeYRe3sU6+VdCbDIpfPz0PNESxw3YMMVbm/iSFDANl/btnS6l69aPq4wn
Zbx1agmZCfBNbnBMHYK7O/v0tmOotmntzyYEwwH8In+zZ0gbV/KqP9Z+7ITFdS7S
w0sxbG+VX2hYlr0EGbzjonMK6ur4CqBuBfN7cpoMN/tqgBNMqRmfnjwXt3ffh0X6
kuDavCJRsPZEihwS9crYqngxtxb99tryukWh+QveAKTuieT5mH832y90NdjeptSx
9oQBVTFXbXv4Gd+9XLRhSplwDMKO4nfQJEnu4fU213lLxrFOuUHCqg3QfAvQ7W7h
7TBRqJcJSnupTMqr2sijxh7eT9izJsWizsTeKrEYywJp9vT9h3bpfXJwc7wtYeRD
4MD9I7Jki6ta37vL6J3VbxwN5mkfAZFjS8XcjkEES/TdX1g2Q7ZvsGfApf6BoeGB
nAFjWfOOGTdSQrxGkDuL21GdTSGB1V7xRVmirwuS9IFNr2XaQFrQt1d/Cj7t1xly
qt0dHohIBvc2m8K/GS1HSLVnvI0AfFrcP9nfgXoL1hDnQlODBF+hqKh6YRa4L/5b
uV/AEs1zKSu9VizyFyM8wQj86antqAaeYGFU9pSPs70EaU4JuKl+0ywtDp7iaSwM
cRPpArCEJAvcifgZRliuNeEkAKypGSYkTts0tW+SfsRkUsgilpPnfoxIRirAHXgt
Dd30nanIyuZbrMupYJSIl/0nx4fw8G2Xn5V4UmTb5nBrvHPGVlOc+IFqdo9FUBMx
70OR7er3SxBYlGJyzJMJ2q/j1h6B9Uv50+xzMyN0Po6+q9qtfpred2pLEGT6ndUv
r0K1SGEh/afLiw3YSS1uy2Ce2dIKTlu+NXcFlWs47fhlbo9k3/i0u42tosZKBZHZ
T2wxD7HO9fkO9fq13DMxw6+opB2QAiFfC/0J0wQjtwNCyi+Xyy+jdevGOgzLkjTD
HLre9niU3TOoJK7JbwuwT0T5HykVfLBBdj4FB8m0fQTbQZwBgMwQL1VIlCr0F2zv
IdeSBXh206WTHMU8Wf4sR5KUVD85NZJ9D3Fgxy7Fq1/cp7f7zGsCfkxw3l0WjScA
FhxoANiLp5gCbxKbPaOYMRsck6oyN8d+V6OlJAalTTiigJzpbD2SwDyr6uGqX6L1
5tmJm1iYqm/g0v8nQvYfgBIMxaKuDsq9BfDhb0e5DceX8FhHwAUyK7fSzhwbPjZa
syNR0Ca/RbguSEqf3TooQt7eF6VrLJ7mvJhO/M7awbTnbZ9HQWTjTH33zuxS423t
Eql3QxDpF8U66zpOKM8Y+ZcU/fXQi7arWqNOd0wWIAcvr1t30AZpV9X57nUW7b21
PQKdu1mVLIL1aSo6+NpjfQYfdGaqCcySqlmmX4nFdKPeY1v2sKmTzrwJXIRmytsp
1clOIeEeXrD7wgKdnwEy2vsuyACWCZPZOrTBziwuDEmByg++PtcBKuBpvuuXUuJq
uIdn2v3JfymUu12GPdsqqfXaEWIpXltiITj3gQjvA6WwXZq7cMyBWjF+dcrGmI5V
Nb/Z4so0QfCBrAHaGmrOGhioVT3ehqwxW9QhbSLHtVCMfrkGSLYTMm9fL5bTC/RD
p4crrHHfj8/+c4XJVg2F2bfLTyYGSVYLttY8PZYdTSrROcTEOLQtz2yaC3hQzZkl
CrtN/CxRMqDNYvt2P8DdhxnddyjiCmBun9hSsNtF/vef/b6tzwcwtBoPwk4+ms+p
bPsGQN2jzPJ8LneNgo+Fl/yMcEmT44N87/M+JckujZ7yeQW3QRQwmutiFmNw3jz9
T4MrnHHhNnrjQWkX/Yh+eWduj7UYZ93Hqmrs9Vwmyo2m5e6wvXX2MyLxFkc0Gs0J
Eq70e153HNMED34sV6IWtYHU5ViWabeFbRd8rvwV1TvqUOQ6KBQ94XwIBUUslEmb
gF9zKT8uZOqP+G+02ssyo2qTT0IAZ0AXQEj2QBrplS+hQG63bt7ExNx1LDWX+isG
00Sj3AW+UVyGksjEZLbx8mo23N+l+oOJFQT+uQ209DzBQ2D0phcwY+SKqrB7YNv/
gBAHl6jncw/uMUe0TYBnOe7Wyu8RsrjXF0MGWy9Pm2FcCzulCpjRBIxieS+Dh6O3
KOZvNgAtgQEgpSQhLPsfQdAI+lSJmdG6ac2VtrrBuHK+3Lm1WloyvVaUjsRV6AQd
Wqstzofhx3x/0wawzdc69w9xdtRxwRFMap20D6Q82xjdTBiYWMbaoH+b19ROqpE9
PicFAt99sZFTEkGnzTyoywrkBxUI0aE88w6FG8Egm6WK00wH/D5Hi264QGua3Y9m
U4Sj+mw1lhSGjgv9RZ97Bw4ujJvyeqtVt4jRapQ1fja1cPCM9dnsIUXY5r0v7FLa
Z8TM0GDJQe0Y9hfCw1M7o6QeQu2gZcaK6mwXahm0TvGGTirQ973+DcaSf1EN2w5e
BOWiJXXZj55R1xZZIqOVesq78Wpg2qiHY3MSnZTYqwQ6BIhTL+9nQQU0ytmSaI/h
SXUe9ZrDhuuS4KxSi+Sh37J1HxAhkTbaFnFCFeAg8ZPXWwt0lrehi++aH4FfY88u
TktOukWPWLJs5kftGhpU1dZ6KZGbEX+pJb8GDt3gsLNqYwobExSzsTnFE6jEcdGS
8uQpnUkXGBixkOhKWWRDkZHnV7TxI+RSkgGlczikGgifoEb9CkAEks8/zY1dAQcQ
CHTfjsa/PEu19LESHn0pdOwZWcYmhKTPkHHmklcI2Yn/2MWIKW3eNy4BHwUaefWx
+C9r8He+ks7Cwu6RQzWJYJ79WskvNh+vZ0v2H6k90B5oxuS6fydsEdycb13uLcLa
vxVYoAM7jGqhjEr3Zgt8a4DHvZ5QoiAeTPsPlsb8s9MdiiYDBEbuzX1UBIp6PA+J
Y1soUloDuW+u6OM7QIiAkEgXBOw1yiyPnx47/XVoorovm6flNn3zsNZf0nI7WOMB
dOAwBHw0L5+smPj6pxsEz+EMzbCA5cjdpP4P8nWIwElRgBbE1eAZ63gV/v5T82cg
4geAurNDTcrRllz2Dk4Qms4hcCv2Wx5xD7ovdDTXwgVqBqwltXUX7Nc/77YnliDA
FKlpAWcLA0Z9IHQ0WwoBuT5nDwvFfVDIw0lKyy5i384/K3XkblT74KSSodQ/BFdc
LEwUIfkKNdDSnR+n1PYgl8KKwO3WBnD4X3cDbJ2leZbYsgbUkOuqBvuM5wt+jwwj
YADyJ21z+JG4ybLHbTQ2KWBrVQMddPdgthUmfu55QT9MV3//JKm80Ml7EwCCeFOY
+wlPD/pJruuzo3N6KxSvA+nOJd/HGhHjUzQQAyzHLQxeySFS9rZYHh1K1myVKfAL
K6mntncVY9cZ3r74UAG6HlztQoSZEG5DlDUP+Vzw882y47Pf3dFhg1NGVHIGPQsq
p5+ZmM1Njd/Jy4lKWYfWD015z+EJcebWiCEyPWDpc1af5W1fGP7i8sUnrc31AfBR
tCaEk1xWcvOa+ZfSqkwnlrZ7s1rHPFoPzbByDIM+lCVOtkg0b4PZxmIZ6Bkc1DDH
tw0ZPhe+5bnO72uF8mAfDD3HehK1ueiEn+cmETBrYMC4xhDj+fZdqKzT8E8BPkdq
8ALSVYnNxdBK2v74iyD5hGN6h+eaQM7XfykexLy2MBglrsvsbRcrOM8OVG52imw7
Ob06P3Qxa3D4bLdKEyqvK1Bh6VLTGd1hIu4XVzxAGgbktBqVqnAPDpQXkbK3EnxX
EAEhvErjfsvTSuBLfN2XkuHVnRwK30gRclIzcfNx5N/1GBbGgv3l1OkRP6vScBtn
GVKmBrO0eO8ZJnkJi3XShKd73ij3o5MFH14qA0bCvpYPXBEdEkZTHLFkONBcPfT7
7TYg7R5BtUZfAt6lmDPf1pIwZGeJmElKDMnfana4xMirM74ILO/gVtu0adRKAUmQ
ha3n9Ne77ZgkIccc1g7Do2sRjucXMus3HzooVIMCNmhZj4fMv41B93qVkFwb+FnE
TopkMyUp8unTS1OyMhhYHdGKIoEWQd/qgBDkJQ29vPORx9xLoyjLha0t67oVuBM4
qVPnNceQslK2ygv90CHVQAHKD4Az6G/yx4l2oIBppHtXLzSv65IqsjhcgZJdxMeo
P+G1qWYuujALFjUauRQpRzTHTxpTydQEA6FA/MVdwSF0+JkiBgDbkUsGEZ1Jxusr
+D0RzrBUBSKxYZ8YRLlR1wWj2/scyPo/qNYp4ECwoWkGggXqzz6zDJU7/3B0G3i3
R880YaSrqDQEU4rUEddL2Yw4FzYAHQe25vlJS6dSvMZJRGQMKHiqZnDZLcFFxVaD
oeohXt1cRCkPEFEs0KOIkNKX1NK/Fbv3DwmKkY7MrKjXOhJNeqj3i834AjhpdMGj
rCrbXqdVy2WuhyCJKTTo3Srj4VOKVlWLiOyx137lOAAK0XPrNzgunGSAsvpgMM14
EoIdDjrgxx8FEfYNSruksoA8o7rTV1ZKpxDPtLNyTyYkIWzvpxyyM6CpQ5bFWTTI
wH3FFwOHsqIHjoaxKo1ITJ0vHDbN/9+6gUY+n8yp9TQZ9aDo464JAeaxnr/azrDw
F0Fnxh668FKK9A/tpZ78u2skIEjVv8KZTOokPLGhtsclQ7LHFVTOq0s0neXPfd3v
Sp2+XYKqMqDTZst5rp0ShVdeRuCZGOqbFDaQFcNndcxKHCKaSWJK7ttbJurK8gH5
a0UBKkfdledOJPY6TBYxF3EQIRt0CZ3B6B631ZhiaPgk6AF5rQnR5gcsdZAl1yRB
zAv5HUTanGZ14x1/ZQJDIMye2Uv93DkHDenSLipGEQYzDHv5EwVGV88SI8MrIZ9n
D9PwVc6VUY1g5VsRyg0oR1FTpMXWMrl1JkK0jRy5rhI3+ar0gt+J1HFjBIN2eQug
wJTQN8JRPn5804042StxY+IUCiZ9rc4WVuIt5ebFnIflc5M+BwGxEQYe7IBUV0wF
EvKRXMBvkrr034fJEYOGQqduhTLRa87iIMo3weUSBXgU/VpCKLnc1MIgsD5oDnyo
VCjM1UAzud3N8l5kFnrZ6MWc3yfnrR6lOxiOp+GF+l0mcJcCo0InzeNdzjBngkh2
utt/6/FT0ABN5eXKYdz/ttFjr4j0b99dSWEs8ZnEXgDs4WhFeCaTOg4vIGeUi2E0
o1Q4qJC+n6Idyxarq8WJZbCymzA5TfnGeGmZsOjS8VONlHo66jxWPscOVjhh3pXM
J0Bl16d8cnlNxvpUu8iMizOeFmzdPq2Yr+Nno3yE6nywrYejXq3o897TybciUX6j
52OHz32lZtqiPug4NF4z62ba6xXqtsaM5yxoKZdfUvwF8zamhTRhQmUzCXEqQvLg
mWwen1+diLPg8D/G2cpMmYySKmYghvAsnyY4spP++Y1qKQJRy1mDRauYD8oGmeaU
+mSud+GbtdGCm5c+SQqeoa9GGA+LBspvE+48EXhH3oP1E5ZD5Ouw1MY8oGSripYN
e2Nsb7uPTSPdo1D3Qoa8XWjNcZkB37x782yf0uiMYKso4m440p+WuG2wU6OEIVj8
3EzDR5TPVoI+AObmvydU4/X/KaOPVShaTVjIM/mb4egnUHoEiLX3x0PTsqtu+/rM
nUXVgRDz7lJRLBKDevvY+DnkluD7kFQc33GnDX8hySulOD3qGNPzMiHlJmykZwkX
te8mUbUDBiZpDBNZbVcd6X1ZEXe7QgWkhN1TOYqqJfOBK+/zXBpDbBOQW/gL8yU7
hOnlWNQnDqKSCdZiJBKNRTUF2lVTdY/wntmv4xII+1YAAn8+Ha/tVIxPgX9Ln9sr
6Ha3phpaP6BY2fRCcUbPpztnD0VfCFCd8nGwcdKFDVrnDP/7/qs9j7ZPDuUMevaj
O1rVzd0g4Xnx2H4cSMr2HLdflxffjPNCaOo0cjeE7qalsgiuqIm4qtDmo02Ge+SG
OrkI67N6evgJV3bbXskIjvgWBy+T8aqwItmdzBo5sR7tbexcd/8mslYzFWJTEfTZ
OZazCMx595uCMnW9gck/2cw3APTmLXisG5NKtAnOGML3EQRv+YyTSMxbHzHEXAsI
d3sD988oRcRMXTEYHJB8zsYD5L2eURUXRaHOM/GFYQsInBXZbvjW/ax4xhw4O+b6
rpTOcCfcliK8EDtaoBGVuCserjYiaHsqY2xrTxnzwmc4mbBsLtpOs6dIKImulSf/
FY/pFfBA9GxxXvixmhfhApcfFwNTCnI3i/XjktLBM4pFcj7dQUGzgUH6zjz+ust7
drruQ/1AfSaaJ10rPpiaot6O4WVvoNOzsYpu9uFNZRNS3rLZ6y6vtsd2DDz4T4K8
bq1ZnCHwA8g958lyWl2cu0HkrMyDmnzZoh29NWm4y6oKYUB+3WAXxQoaaVIIgW1T
1oRll/xuUHKusVemApFNOGR5ABbiCV0sg+oW2kK0ucr6CSM0dlRWN7kN3MxZt/8e
MykXFM9WJ9o3HOU3gnVkaSemVWbin2gMJ/vgc0AmtbKDtBJLey2BLuKuZt6jm5Wf
Pkddb7t+2hc04FRSzDDVez+z1qljb0vIDaerHPJ71v0VIA1qRiPdRxy9uoE6+9wO
DD6akFWAlJ1+p4dRRg1kDlDytzAb7K8XcFQGgfGDQg5Dfo+xKMzOE9zoleXYtS55
DbgE0rW4qZzt586JtiUIOkjNNlU5bMI6Z72HTlWPA9w6S53VvWOj4KFfWaUkIGTx
DIfv1aPdWGY8cQUY4ITxCg24tZVPASc1upFaMu+VvebyAMv+oZp4O/yTqpWDJyI7
Ew3MnRqxuTccWT1aHtN4jntc17uqD3J18rJ6225K1Zec7fFHz+04nuTa1a55jhEG
Dr+HNXhr6uCFqEAT5+SS9UrNSkcs9N2xf8XxMpoVAtbdUmlCUpneVQ4XBYdJGJ7q
NSB86V3f4qh5/kBh1SuKTv5s8/y5stM9VZLUQRhv4b8KtL/N1cmSwIpAiq8CjeDA
AJLD674KBafudYQ+pEWNmbWc3B5zqp+3vM8rw3Dqh3lJC77PppxBPRHAG2it0Aw9
vG4WLbS0/21g0sLXmzoTG4WUmIWM99VlZxyzawoUQzhLGl48fpGpBAJNIY7kHWM0
3jY8C+5sPPr7LSGWdTbuKaBh8C6rYhHd1/jf+b4gqndfSxvLp9GHhe3rxJBsEN0j
AoWw6aKyu1/ySW5C3VXgijk4KDEXlxuaSEC/Fb3Y8qzk0pHM+kYG3JGW4M8SipFN
+osQ9s++2DYiIHLruywBnYY6iF4cHIfKWjbI17bxYCHh8FiSQliRq2uYDAup+PST
aD2VOSgTgoIFNyX5Bo9+WDWBzXtLmeCZF/hU1YTY3sLrKQ/r7ZS2sR1lpliryIgY
88u56mhwIA3eQnuK0bjQUDcBi8JzZvghLEdDKHwpveifCdP+GA60LRl9M5SbfnFy
ZcD1paf10xrLADz7NMUybG+eScvbwV1uVvtuJk2WDE2j1nPV2K4tp56uEZWOewkG
ZCAl2DdkswH9zWMXiLg7ymXbygRUEWxaMAVAigX49JdPkvmqVChm1cg62IaJfkxP
1JBK7mXpRolDjKNem7HkhSDejuy3Gup4lQxNRRLHBd8D4cwVkb4yVkfcUOqo7E9b
B+cN8F8Arrk8MTXp9iuiPleijdq8PMeDsdtRrs+FXwCSTsH4Kdx5xaaG6cqhzu88
qBe3lvCxNsWr4kr9jkrIJfzq4/ctqn267WN1+QJoMdXJpvL2i/hpRjiR0SRm2cxx
QxvsY+zlKa61fizNwzzyqdlVZwd3PiYEZxAnGnOvpViqbBBYlpz/gt9Q+s+evYJd
T2JCYCzI564uKfcEuR9PTdkVxqOBlStXDgUdFIebbiK05OJGvz9CZTsDAnkHdroZ
hB9wqBgXMm+A/kAW6Cz59NUq/dLidC43YRFfKlOsVCgjsxef8tqXeDAvL/QRa7WV
te2qvRCJtAkvwiCUMMQ3xiCQHO1lucsAbOEhUUIa6x91X7naDwl9bVgkBCBoUCqk
pPvtgu7KWUiLUflprlTomg==
`pragma protect end_protected
