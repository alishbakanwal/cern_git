// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:09 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
p++Xbwk2EX87r5bhhxUEN+JRbKCaTaSe4hdjq3MlnxR7w8gRH8uS/DJXQyZoi7Bd
X7EUfdt+yxhwzPl3QYsaLh51qb5Ow9UkysG2sXE6rkM6TXMXv7FbOxYTj+UZaK6u
VhLiGbIxkMPLSGpMGTVgd6sJYAPaN9L1a9QOi6EvUnU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18384)
OCdTI2uednxpaWccF+J4zR1vgNG0yieL2kbs14g7jlv8jukA6b1lUCjbluWMDPLg
Aa1sDfwBWiFagNEz0eNDGhk5zxRVCRIKplJ1+7POlV51otpFtWy9GR5nJJxhUpZX
rjVaVdIXZzzUX76M1pG6YQhjgH7jfvqLS2nA1h+zaDh7d9rcMv6X0elwmC3rKyXU
OZ4xRoWoO4qIfVZeP6+Q68vGm6JxXpT3aGwIPLubkYkED0Ce08soOFqLXmIuNEMB
EfmxYsgYfuoa0vtAIZATd/DUU6/I4PiWj+Fv8VOrO7S/dIeH+mHDqQlfmA3+oxaz
lkgbD15YZTFSl73DP8v5Hh+rDkOzGPItNiIAKYpWGdUoaW17t7mlgrVO0Cpnh8X4
cxw9S79s0o+fhbZMUC6ALKYtVDWhZafRPFdbjVMS1OO3uUYTO+V6EQPj/dzuziM0
obL2S25uZxQMkqMX1Wv7mET42LxIWUN4bsl9DmNku5EmdtQKasRDETCZUzcIRMkl
dQFzVAzKztzh0PohkI6xVGETKrgC5QKxtYIuica53Ip/ADoTlk1BIVr7Gur6BBTP
sLpa55fyJ2KvBonZDUcsIzZRbPYH3r8/Rp1Cqh2RQ3PlUAcixze+7Wdp8Umms53K
nd8ghhHSuuEUee7n1wzbXiR8S/LKIuS57gdH5FlXCecRpZetUI1vcGjHjEahh2DA
eizCcRGIsT5vLh1cxQJ2TAYko+fewtvk2phG5GGhijXJqJ7A9a4rZUdGze2v9MFj
K0k0FXuVTRjfOWtKinRTK9VSt/HHQ0nw9Q0aW1froLW2LfbZYPqVYkjOo5dBAPJe
E1C1MmN5a/ENuU4q6Td0fMsDRTOwTDa0HyjXryleA3qQ+YzAmuO33/7tLFHSPgK1
gBvANblSU5s3upIhjswIGlcPEqNS+FC7H0wo+6rSNkUinphlrxeXPJEnK5UXxtVv
/JQ1UjLYpA+Z0XRFHWh1t6ghqadh6H5Xtx7zuTIgHMGp+FBkPMp6RtZKV0RKJ4xI
AcMNywbyNjaEnrZS/bB0AsHlSldw8EncMvn7LAZhpAzRwwYId8KHsFdM9FJouXpD
g352sKy/cM43kznMFTcTRznoi+yS2hFLWH3+7m+sruPadGxpcMlRo0u2jMwvz+Od
cAt1Of3Vl8C/PvmWaf8yTgqvo3ZzQ4AE4atmMnORiyYu4ZnZGeqyiX7t24L4WmyG
9IZLS1ofZ444ePaTatligT18N7sEw1Mlg+7UlL1qf8QmtquINLcVLtvRRzpNX4a1
4asBtrSYchUNjvMF7a6rwgSjQ97x4NWBVvz9/5DGYJ8XJxusC+eKtBdVskIJjA9C
tt8s+PSQqFyyN74zskSjks0jJMUYNXx8U//EcoklJ7K+3TJPf2TktWV8naeJf8rJ
To/J2sPVl9HBIKav1li6Z/2VJmejc47alWZZrE8Jf68hpeKxS6nzYTRLfQ81BfU5
NlUeQ740SE9POBbAhZLnRnq1nRmnc+AfFSOaQLzMVDBIoVrPMwYsCLg3UrAMZi4D
YGdhhg723ORfgcp5i/pY5vUq9Z4qAFBizV+lNNdFmvQnv6HxOpjW7XJCaKvqVES/
Ue6IWjxPDa4V2K7AkeJXaO+XB9qc8UvwfdA9096jNR6RPaNJZ8VOtmxBN5sNA/Uf
iLwiMSVvlNP0xl0FAk6N8yte/aof2zCJZriv/Y8HW+g7wkj+9WyNoof/PblSNZWh
5NyF9jTFe2bFjK/ee0qNKxOm3EApL9ci4Hl7bZQT4t30mV0g7MdOXeHL54EJ8a3F
INs5lUsmfpxbFjspLiJ7EeStXWuBUwPyCYdsRf6ALvrRKVCaNv+UBawtrFmRZnVe
cgxDotPUk6ZQC3ZOYfgxdFvtrKAFshm8DMIPKcNUMpS68c9zFwnzErlZK6kJ+CSl
OiWy8LcRUfOgTZqjnNHOPjeUV4BiF5FdKSRTzosFa9nriILVWiWOWeWfcvQUV1pU
m42PaOQcJewCVI67zCQxM4XleNb+lEre5Zz+eYJ3mITop0Q5GHR7uh4gSmrHjtW3
F+Yi/Cc1whnv/j6JP8EjBp4RY0mQRNSUD500g2or3p9rMXOxDSFn7tsJ9/6RBqDw
ox9cww+Gai101cKcBXUbNVa0DuCNORWfzB5wEBUc2UD53r67mJXGTJEqF73ix8GP
XC/lFKx7iQk70xIIt/vWXc43fUvkNcpHnVEelHIzaPR6zgKw3eyIrEKT5oyqZ5tB
FJNZwPLPSGsIoP9rxIDV0puMg0fNFF4YmxsQPkNe7kNZrzZVztuq14dzwrwTPuZj
wr9Sf52zvMAj6PGweljzhqjoYaRWi1R0Cbw2VHdtBO9pDBKkniyQ0GdlPNVCucvp
+9+N7HGCv1b1l27JG+Jy/NlNsxBoglcr+8/7+CfQNDlk3k/n4mtM/WbE405OAFkm
mWvdW2Rh5udkvW/8S3P9IJfNceYMCtDbqGVOxQ2lRwPWRrtjJw+dKVUlK48GzsQy
eRwwat0NywSTRrZRXT77audWVFpBvVuyFlanZr4Ug11XW9tWgYzBo1c3OhXpYj8g
ZWF1FZIYFOg7reihewbDokiU7sZBytAqQ55wQVDJyBUrqhyoHBpCcVfIlnovjW+E
gCCcDuzaFdOSsYREZC2/K8Qc9ZIlTu6RbGvpaeVnxNmqSkfpUFpa/BgkmrlIJ3I/
V2hXFiQh04an07pPLExg4UhecSwCzxmhBg+bJtO13WUNmSE1B40xkk57rwFmMGIl
THSLhLENutpmLSLmI86c0gATjgcpWiGpcPqIR1PKT7LQpr2kFwpqqA5FhWQJ9CH1
UIZKDhhY77y7JVQgvQ1o6DyIyHI2pZVsGbcoyA7rCDxlwlgRLRJDIEMvdJWp3Pla
j6J6fGOKQlL/6WAZt+mPrqzvCaqzCs44Ug6wHbv24mBCocRYact0IU0KfaV5KAzv
Q4ETRihiY9+drerRHO+0hgRHFgZLJrejM53gB05uJe18D9Pjj92OxFkhQfIUiY8Z
5FI8RnLtWx/q5RHuxq9lb5Jg/MzLeqrMuy2BX0cGP8DriOLek/aG0ngibL2yp8kw
RZKpvkDTSip/e+wUdiragckqhz4QnFo0u1SFXxXw79vNl2jrqwm2sdRQFyADO7ff
bQ9EPPtywDsXfiHNZkmKLhbxe3zFNYQKVrP8UmZ42oQHK21ZdYTv70NNpnWS2hDa
0xfs3VFpl+uBWGAi45HmKB5mUcx/KHNp6jZ6qB2TAd1Lw03k6lgBHMw9wgalOZ1Q
p+lVPe2kxuTgI0xeej3b2syXwASXhT6Z2FFygiiP3+AWkv8luYSj1bb+hX81C5eU
C6pMAoVJNNhHVGXzyjQEVt+JTTsdpeXvBJYBgzfPyQsS36M9LVhElel0a/NempTJ
ikgjA2ShFKkuYhsapelWRJtrYl0rhaNrJSqh3iCP1+DcL4y85KWaThcWZMIWmnnl
Kfo0a8P6kS1xtonK3LZ1rQUzoStppK2znSPdiqImSLDk0jH6a6B6/9xVcNid2bK0
IE2hIktoPGDDUVa4YmBUhxTGjPCJkupCdeDFF3jtRNi8yZk7icp9PPPntllGf/re
ZOP6KtxZiUZPt58PSh+2gzoJFPEIw3AC1WEUP0ZmqrM0NcmJ/QPtv4XxYK7Cvegu
Gthhu1rdYaNg5kb4rk/7YBK89bqDV0dWz91QZELa3kvQDqapgCNUBL0o/5WjgjXv
85iMC0zkh0GzPMnCn/9H5gjWPVw7BLjCMJ1fjdrwgFLDvFHbk1TfaCKyN29w7W2K
8FVIhTl63P/edc6671ofsSGs+73WmU17HAmSS7uf2/VnTmTXic7hUP7W3LYc1fVa
0M3YOUqURUi7z4fz9Nxbome26klzS+j4v1cLjFQfw8Gyhyy1+vHVLOIIzpQeMISR
r5ZRHd2Dxqi26MtUmu7gcT32a2KT0D705ghkmbGmFUxiHR6MVC9B07qihzr4p3d5
9el7x3TTFAr7U+BeP8Mb7HDc5v9V6wmWPXLcGhK+hYGFpUog0y3iXy+Jh19jTlZX
5IEyQ5aiAATF5NDTZi4EFI/Pr+kv1YesL03AT5tE0fiVWxAU3Kc9j2zIA2vjEqRb
o9+whZRnnkQCckK+iZ1qt4v4/kN818zLxXHiWlgxkVlj12fQI7lygU8W3GeKJDS0
2aoKKvFr4BKHlXEITiN5Nrk3Ij1O+3ronCQTh9tpgTxz8BsllTOmW8nM+M8+kCWn
pcqAKnc+11HAxz/bu3PZuJXoLmz94dtDE6BarT24YQYw+6B4D7XTGWcUOIc2/QeW
jrXfQNe7wROTbw5jimZ6cTsRXJg2MQhJPwjglsISCahrt5qswHp00uHmTHHxmjXw
Niso79eGh0YGif/k5WiZgXTrXGexfM7FOMnxQg2o9Nk+hYGObwm7q8fEmjrtK5jp
rsMuQ2+GiI7yHIZPlFRbVzVVKp221q4oQuwZK/G8v7psJyB15NfNHt1dim6n9cYT
X0S/qOONPneQSUrvZuxDxIG0ePL7EkUZexj7i8CyaOqoQhHgqEqu22LT7fWgWvhm
8Lvs5Ad7Hx4zY9h+/ezGZQqBfKwiwm6exKdW0RjUjWDA0D9A3f0cDcL7QTyjCzKt
qi/coawa7RPCnINiMZqauZESmEn+AWRP69dbyAOSwbdTLW3rkqLwlV16pG01WsfJ
z+lGNpy5OsWcrr/qYQVTOUY17j3Cr1DtEiACd72wQtFgNyii6TAk2qC43+Nqu0mF
ZisuK44pgj6eiSoJdJHH375kKMKE9tb6kPxDg8evjC8P162ffTlqbrhpBEmeslLb
Qz9acgDkJ4AkHBiWXIYMXXi8YNmrV4Blih0V6qwzgaRYtWIQeuqkFaNGcAL92Dcp
/Nhg8hC7mlnqkmTgQ1LgN4iWtRWrp0yYsK+2mWPK9SHrPCNgNkp4pgi4Q9UAL9Ls
/SJGSgwWO9Oq0poVaPjMnc0QLCoqSq5GJFXToGyusXhlTe4zr5uJ3uDTFtPJhjdP
FaGG9+EeJaE6qg+PA2MMds+XmvIulm1HzY1+YTprUG76PeolqYlvWwZLqtWLGnXM
OKuPM/k+xxR/Gph3qgEQy0HC0GiSJXFJbif0hM5eX51Jr0dSCa7i23aJJt86uFGo
pzk/me8yutSeHB3DcnT7WJ8UeJVumXiwl+QvCJZVwE+9wTzTSnhRNWG4uuxj+xZO
+ppr4CRI5gLVoZ5dLnfBmdYDh+vylYBkjkC77f3875MkzN/I1FwUEompr4NDe80a
NwBQV6DUWTM1cWyTT533S6mv1vQ7KF1TxDlunAWYg5yBIhHZ+M/mWBKB6Rx09rM5
Kymdr4/Y/HObkCGLUcxXGocNYqiJQC3R62HGPR8gqeA562hbYo7HzAbxssOVqrL+
zvTptNnPfp35lRY7opAEPVXMmLYsr5tb7gMyCUTZHVuS3YZUVLVN0LK1jU2tB+i7
qYWhtuTA6LJqCIv2lnFERYhgXScQhu/ACsNuNE7TJSHWPuqrm+3Kvab0/cSWACMf
hVCmkiQ4BywTJpGG+j28eF2IGYug5h6PyN+qLNBW+hTI71BhMd2im9FCy7kYZb8z
iifu82vIN4kkzIe0e+yD3/9l7e0MKvdW4hwKeqYGFsqWl6x5dhX+BkHd5VswYpdu
knQVAkE1yO5BMNaP17lPKCcAr80y/dFxhpqdpQopUBSPke3XRw3Aca/c/1hwjJyG
KZ+flhdtZNdWTpUTvHodOcTrl5NsJDwBtDVTaqmiQl6ChvvWuq0NN58u6cWWXQkC
rpgByIMCHpDmOyr/wNjNXlXsv/7LtaZjMnqrFUz2+QzRmWDc56Ma6gPQk9TydD1L
AgrfoX/A4D+b1yAllgfBZ7ggFcYkKYtzv35vYWhIKogmqj+Cp6S8/mrroed3s+Xc
Ms2TXFIKwBPkAQb94YLmVYdhSNwSKhq7ZGE3RDpfaGNE+jioplxM6pdax8oIU86N
jLHHU6dnGodNRMgO0WmjYStHEtIsr6VGlCh5RZAYwi9z/H6+fEPhrnuGUi7qNr32
/dPo7uTRO1gmuRr3Mhe5Z95u2nkegmXjMO9xIJR1kEBZLS8TII8+4/rDprOcAWY3
TNA/yLwQbPPhM0HqFbyXvHqCIpTCk7F1TvPSPZFzBcNEfeep41/1WlB6IjUqfV5s
j4k5TGVL8bH4XDaIyNwHznJ14dgUSOn3xGSFV9RMerG2dLKxZYczjY9njlRHZlYi
p5KD4IZSzFT8DEJDO2Xpyn1KCocHDhPcM/bs+LWVtN8OrEksIJKuPTEJYEZIuu9U
fCUHrYl872ZcRUaSy96YutCbdM9lsQjLScFyyYYPKTuRS5fGwu0rn0EnkrdDowhG
bkwhG6O3u3avN0MJQTbIX2uiZ2k1IUn+yNwTJdeS5lHDGRBPVBin0TIea1s+TnIO
qvdVB/N7u0cy6JcIS8sfjwar1kmAk23kppj1VW8tZxziK9VEmBLf6mQOKHfGn2TL
crQh4o2qhMKRb8c5HogubEku0L2GtGxWg86Twqeibqxt2L+DPfoDmQbpHCfFAOM6
0Kz/+7zljzOtE0kOyOZrBEpVc7cRaE5hiE/WkrjZ/M0eX0ADfYRSFyoKF80N0/BH
wU96cp+UPoT5oy9HP1Q6p6/7tp1L8LeGiYcLDKOIxk3Xb3vhusDgDERtZX8uBW9x
nRMK9bGUpqBy+pIkHk75kJNU6/aTuOOM1hPAQj3lVALQCg5Az0VaVKUB29BQBlZf
JATAkuan/ywFV+5zNU7Qu/Mts32AVLK4JvuJJoH6ftJMFfMkNE8rgktN3IiQLepG
WINeBFNGmNfuz2YsJVkPw48svrxFBKu7IeQSC1pzWzJ23fDEd2rlwB4SueiAmK5X
0XsGATPeYW0qfmIB32ZjYM0LVzaT85Gt/f4WQ/qJdoEeo+JsLIQiYEXOASZFDnko
QUqgl/0rbajPfbURWuyg1VRs6wckPol3BUW8YJygcvTh4fYw9wM4kboqSg9BhZB9
UHPX1AXZaQDlHgGodoDgaqnnXtVANXDM/thS19ijGI5Zs/U82ZdHuC2o0XhNmksP
N2k4sxCf3XwLzx0bqWs93PLINO46S6NTTzfYkXI3qToQ3lMhIFH6Bdumv02EfsS0
4DCnq7uc7u4+Al7hJLOAhSOOyYvpVqSOrVtqEdZJFYb6Uj6mgCvLwzhG4io9Nf8S
CH+0Pb3E9Ia9Je+ObXXMcggUQUVJn1t9YsY/RL9nWQNZYiRVfR8WvtW0nlzuBldx
YkEpdYAY74+5PLN+mWGCtE+qXPMKPtZjtSek8gcavp6ajGpSeOUEDxMKLqA4EcTz
1yoW2HtsESD/oOKa2NkcEThfiQtGy/vSMdkve3ha8OS7dvDSyeA5ZPTFb3RhQa+b
TIMJTfHhvcy3ydCoPNV8T1Osmn6HThSi5mgT3uFIdGve2tlULJAJPKUn9E+tLMoM
JQRY5Rhk+WfBbxzTsV3RUBTZyw/QjljpVW97BGlib3ewzJuA3xb7s/3NW9IWHCgL
iRhC/Y1ATwmXWtExCzkOqUwt0TzlhcqhfvfcrnD1DJosfjNuqVW9vc/0qntpDPJt
iB9OowbHtNCNZE1h5HtgNqRG9ftnmv/7w4TO0sitYJq1w9RtheFkW1DQMVcuHpSk
iGlU0zBKdmuTjpilIva1GeLUBXv6wMeqn4WHtH7KUYvRMy6MwVnT7SJFl/4ujh6R
qp1ZfC5P3bEetSzR0+JxKzamCZ0uOZXvo/CsvfW2nrJtSceCgg0vxMyPrEYIiQH6
0BRNRzydEEouO4/D7mW2BSbporFWGVu+KTUkdmoGc+blQxpU3tX03CXZBhpVdQU6
supr2DJBGP5vFYamlIPVEoot6Vt1bAw6M9B1gIuqr/x8ZCyIWSsIJjcJi1DPHdri
v0fL5EvH0NyOxuMdNGg37bQ6dht5WvWlIxu7pOBFr+p9kBJKBfhTAN5JIsLuAjuF
1Sx+BOQ6qpKzUfJXMd78AskkEeMZdGJJj89peOlj/F4gdC7AZUmA4qk0VJy5vGL/
FA08GXDYxhuLAJqJZR4A9uky6Q4VXJ84BeKWWROKTB2vExQpoqubnSCGWa4WaiY1
V31cBrd3uV1GkPg4/VR/Lgx7/hfRKGeouDqUQKmHNcFfjt3Rpyd0MOCXSPBBtzOp
xZ48qKaqWgNyF9ZvZM6/ahdCLHPJzspd2KPtpgQHW8WmlmO6gwVFtmu3gs4nqGtA
s5gK7bK1SrOVxsK6IkpsgKXNkLZGJpJshi26IhdTj01FY6lONfh8IwQOcP3UizRL
jXsecEjN35U6+Q7uNN5dmBCClqpXgYhhthIkUVKZEBD0L01auCcmeeHfWWPTsKsF
96uMZtzrUnNSddTcW9/UCiYRUD0BTSaBT6MjqvSsN1RZWvxns9fdmbmjthq3fQOC
F33qY7vqxwOKW4v7EaSlbZjkwkovPMAtDkPrDBEJfve8AbdZDcd7Qiu9yXifDOh/
5/6pccR14ax4RsMrhjBbSEVIMcMhzQ/uHMAx09oWGrAfukupbxHVchvLf9IWjDbE
ZGKXcq9bG7nFOFv1wJ4LSIvj216FmFKSRosYAMSieBFmbv8I+2+gPYUMEVgI/Irv
ZHUBZE+HwMPMR6gNwJH2vupa/YErjVyT1WbwmVJKzyvwKT5hwdMLZ18dQvJQkHcB
JVx8euhCDVSTCiJKcKCg7Ww3EE8ZkyWH4Hl5LiUVfFl3oQSo88AU0q5jiGKE+sn+
xP+/Pdj6n8Vx8w+hHeElEiHtz6UYDIFTYhM3Jv1p0UODgNKoLHVwDnnKR1E6VuKG
Vxg4kUpcb1qyzkMZBiYK/Bp2N6yw0Lf+oiFxqNYtZYBLAFdzcdsGVUU/pSl4IJKt
yuMm7Q1IA1qs7EcbOgONbqVBpX4vj1MAmgwYJbCR52W+FerGy3CsHj58fuTL/l61
2vsndFzC80u7JiO5DQMw3jH4s/JkWSjSIQfCkNbWjilqLHOrx4+4SQg3yEZ2lGOG
vhGHsHePlRgKwterxxZ3oWlrgscf8vnpnM8FmiQVJl8HHceQtwiD6Bl0ktq9fTYA
0jFocJ9cOH6IgPbKrtcoQ8NO0Ko7/9+vaMoYnmHn7ewH3Xh8Sxwrwlk9cwCv7bF2
Hq1C3F9O33Z9kKRlhbJazaeqAbRsOrQ+0W2v3RmSeMgBVBSlEy8g+3KMA9USHsJK
KWSV/Xlt/1lkB1m3qcpg23KC2OVmVjA1OKuuOG4zzqJAWgX3uRZAptObFJdg9fR4
MpUDytTNNSaXo26UOSYYSpvJ2EQm9fHVhDN6ak2+2zZe9Wa5IkT6bKAeKeR2DQAm
wQus4fY23q13xA9LQVdggeAUskf/jex4mjkJ+fgAjIZ9xXMjoTjXjCGCMWuP9OEn
u4yMKj6eTk8KJ38IGMXP2ktqZ0sn3yXmEhzk/H2c9nmgguDiLXnAY8lrErBhQANW
00OiJWLPRwxSpt2yy+bBfrpahhsEN7s9vvcnVr1qZU9R90PvHb66j+IT3WY2UNdj
I1CMfAsUd12S1oYNwJtAjsrePajUR3WAAJKXDqBiL1wTzCwHT7ndQPAsi09a3sje
64DofmG9MTHhDFzooSa3R2lHYKdbAtmlpxJvRz4LVwkfThBJw6X6xyLfQUmAY0vR
SevnCxt5LLNwYt4nBymQajiwAhVIN1kwjgBGsoNTtAsCSoxs40uRYzTm+wsoHPvB
5TYorF2/3XZQLhsLq0tLAOiIoBWnzubUMe1d5DXaNGbOBvTdpgku04VHQF5RMehR
IiBAolVX5PfrVPO/6scUIaj8+fRetU94MJI/DBU4N46UZ1OcbdV4RgsJaVKg9hHV
eVYYG8hh/C9jvBrJ+vhhacEKMnOcvQnyKZMLDMBUHpVlP+d2XeGxPOiNUX3AHs2M
RObm80XC6P66NDkX0a0khLqYmz577hVSez21ZiIWEx89LgRyx9nGB8ICRXbClmHy
+w/Vjg4153XxnAFXk7qi+0IhyzeemC44ugOXgAjOPjyy2U2I5aRDM60z9A7YLlAU
FEuyh9jXJVLN9sXpKyQBPxLGZ2cXiJ/dz7PyWnAaxjqLhODR+NHS2/XAjRx4ZZNU
82s12o9QaBulE8m6zLrME7evMEBV6SpNXGpKjHOSmL9rJaAOBt/2AeUL/44+mDDV
RT8vQj5K6z2s7HV3gy/fFmbvq3glBUefhO34cxsfzhBUtuAX88qu11AxFSozqFHG
y7Md7k+G2fbfm6JFoaaTWySaqoyFmye3VZ1TowTx5LXl14LPDS0+IwnZNBufoUWE
NapgT+rrts4pis4ink80HYn0foikmzDMWfjETLXKlwU60GHEvzQOYi6canO+Frpp
nxV1af2BaGuz0JFEJAQRHstuk2yvoqYQWMPeFb01E9jGgz3IlpI7O0KQkemREaZ4
wyQJNs2KBtIWoWY+mL6hRL0TjMfEEYdkF2cY/+PMRJYjxn20EXKjljVfBFJeBEY7
hpoSY24hwlN1iwexMxzRpdb0+zBFKcq4C+1RyCCX+whgM67Y4qZOORpym36coSLT
sgI51po6iLhD8npb4YD9UjehQLMlk5pBL2DebOQXit9uBWermvmzKzP74i+l5eAT
xo4WEXi1sNRld1lM2f9ApUcdeYSiRXcqvGWzkdm67ExwCU3xgiUOsQfjyPuN3pB+
8krmSE0C4/cILvnycQc4Nm7Na1huR6Dh1ffgtN+Wq4bLpjw/LPCjoBZvAJhIEflU
RkyXsQwqfn9Cd0EjN0fiWGWS+6x39cHwYE29u0SIPX5wJYkx5OKAJicEZp9FQyVR
5oAOymnohHxUeaXFRK8ZAG+8zgTCIS/z9R5r/zEOEOL5BU152VGwRbV1ixC3ICnV
V/ROfZzTIA9rxAkPEpz0Eg5Mq0xIHmM4aNUz8NnlOxUyphOTCUtdpIotnokUKAHp
uDCCW+ezv+bLWJXbMf+5k32ybLBQ6dnwtTIChEjhZVoYk4OwrDc/FS7AhQJGoi7a
dBnevILZxzgXZLqq+FL781q8beKftaFa3GWEkf/n2I4IPMTGvaXrvlE7nnLv8D3u
fDJ+dgOXesn5CqrnIpOILz4KUVUXqR/ee3EOjmtvIJQ2CHX8uJ9KAVBSKZybD93t
FS0YlNHv73V/TQu0gfuzqUuoRiiVJO49aY5vZhdrVaFiL8PE5km4ir77mjCtikB3
tFFiPUHi0R1I7oAD7X7rnqdTH+m6OVamEFXHtJmhuh7x3LZ8Lnkp+B2h9Qs13BXN
5ydrGi6w86JyIChxslgYJM1kxLR62L8vB4utwKh1qm1jIPpVX3pVcWEBr9snVppB
mT36WSSQ/3tOlZ/9IYq1SnoCzmHpRo8MTC9AHYnx+00EVVLwvecXIShGmdl/ol+I
em3uE949ndzZfpdDFsPSqakGTOQhpf5Ve0KakQJ03sWETiyqbCnFxC1SDu05lg4s
w2jPRrBpVN4x/r2EUe+BKwjJajaBsYvZXT+T+rvgMTdv2ZxMMBLsUFbb6ulIZU74
KjIapN9Y3ikLn3UmpNfZChgGSHt68abmj/mjhwRzLyvL+qtJ8VrA1E0Uo2ltXQlM
CoxgJfGrL7IUwP8i/AYufOSSoNTjX0ucqq3yXGNGAJ81EaoexboMwI6fLZ7f0CeR
DsY/YgndTyA6eh+RvezGRqjtZFHaNiwdO9EF2+JfTBPtiJ3L6rFuPne905ylPG0H
l8YrxM0p03u8PqktQ0Rp0e4NaLXUCyyC3i4IhoRnsT1qgsXIeuAlF1XrbYVldPmm
OHWSfJH47rtkdKWkFO27HLbfO7+lHk3l3rrqvj+4cMvFJJmahPXliEn3BF2s6l9I
bbOyKlNTUp8R9JrYcDrf1K88miLDgoBGV9mXrojljO+MpE8yRQRu2YIQcyVc3Tue
pqUMTykBFW0GhgwtHgZTqR3OzRXMSUqLtfXapakic5y6+yOSz8h/mbV9PsrL50M6
fj4xaf9PyM7fH1IQGlhExrnNbkFbJRGh7GM05WANPiAyB0i+IH4Hy5swkQwnd5K+
07I7zbphPW39U2OUaV2zm+ZDiNn9uvuF4HgPtU6CHfZdQeOYyYVk6jNwc49+SeIv
9aCzo9hOSLnHU5+LrAVLAbuRMrroAoVUyi34rMvk1/4D5QPJtJl0rYFwSBUBP5Ev
x/5lG+yF+euDNL6VoLZHBuGGK5F83X/B04wyDW+XHg4iyxTygYw/JAylH+VviAKz
Ep91FVJW18OhZ2z9GTcwP941lOrrGJWxTnf4pFUyWyzFGg1j6IssBCwChkr+VtCF
U4Iq+yhopS9ieDqZJaeY3r67g0cjdXV2/wT9Rb2f7TK6szIo6benV7Z07xvpwGEb
Vt7dNj5CQ/Xl6U0k2U/WJo/oal4sCQVcMR979qIf0UkkQG7AzMHr6VrSHfNsKHFQ
zrETV2UfXvAWXBd5Czy9heat3oA9I84UlrMwQqAe+aj51Rfk5EWU5uoAVYifYcQr
KO5eeKr4vr4J4LOmSdZm9cMbGgUgs5hLeKxPOoFN83IRjIVIQJoET1CYs84COL+R
bhEYbBZ5q0vkVpCqs1kE/C9FhT7/QQ1iw0t7G68QlX8zwR6CZ+KTPNnjCRWTBdi9
44287TO/Rb8QdVLlNScp90lNHTju5xKcJhZISqS6ll6GQD3mbPwKJj5puH9dgdil
QOHD+IIytHXNJG9wSWO+lsJKASlp2CFGN94bA9vnh+PrqtzhrdvzbNWvgWOeHXhO
8ldZ7FFkvi/ACheRvR5cqSZmMzJGbFmJ/shPk77Ox1Fo3qSxMryUbx3V3QSYslin
2K4mU4ksn21r+RcvOxs2Rl8OapAUHYLcJ2gnZk+6YWLKJyosDOQNGg+97RC7WIqZ
qOOTEf54RF8X5NOYdIjRdZIPgkvllucOJCZkMw9SjpTMJwPJhyXiD9FJphh7AmGt
uX1IsAMssOA/rp1F7kR9IFcRbWmz+FwBXJ0Q3ft50djSEt9mZ7fGM0UJ0slBUPI9
bxWUoD8mvVwk5iJj12EnkMCtUuiLYSXI4XZuYXTqdz/5dogeMRJeTigHaTON1zQj
5jBLOblSrv6zRegLoHo7AU7DSumI53h+hzP1BtEi/O413ozZUwowGosDikuoiOA1
DAj/ikD06Mm08XQnsk08ef921COZrVwjntkcUM4dA1afJP2yXUnTtBie/v+46oTG
1YwilDLW6ZYuAlb3gzlebN9uYZVD6zEvBoGYPXJ5vy+EhGblQCsV6b49thrMcljM
ZsahaMxGmLbAM9iMx6ahrZXeQlevM7Hxa410jExY/iUaEUxuesLJ4SCznTjbdQVn
Q1nG1VW+5tSCkllB9k3MeUVnLFqas8Gj7zB0ZkW8rc4wYwRuRUkPnL6lz1UHiAIN
c20mJR6SF/IGi5jpeYX3kdAWnCpFwsGHS2bHlu+QOLbNX4Nuoymut2WyXKvLhZ1H
mvO8K+Jx8qxdLQ6rkmR8CXv14ZHJhPeSMV/D5gFa3QdaDZAVDA8VuGeZG+it/nRE
cSoaJwJ7GQE2IBP5TMX9HgNBJkocyw+/n6lOVqrYRkIVtuaZXUgE5vZXr5oqOnMQ
2W+UDFQ3VCOpA09zMnWReaDwveDuPRkMq2LLDY4KTkqchRLpMNtc7vrprHE9PIkO
TLcMbDBjC7JnW77VvtgJZDqAR6eHDr2kBKFNwpYPl5mQA3ZadS1NU3M2db5Pc1Fg
hn3TDxnz8Zw8Ifj8oyPkutlcTj4Mypir9v5DJgyczqmql7AbMkWcLZhB2zJJsZre
WCEVxSb36msa81VdBkZF5D02u3gEtxMTfGuPRNmA/oItfcSg24XflFo8fSPIQJQk
Ca1K8uvKIaXb2yL+s61iKi1hQg2cdzyCGgHVe88sIPebvxdNElgJ3LzmeQ1gWHAm
T/YnE5rzFFmSMZOaTMfYgX09bksiL4LhsmT81VbdPW8OhmkE5NUoJ0CrjuLNxABD
rVt7ZCmgfWIzrd+ts7y5XgDhNCNFSxC3rWhxN7YL+QzgYZadlzAuZiPTMhowAR1T
5PjfqVwSD/YVocokgTijfan/Gh+1Uv65ryGYDQCwPXI8D8U8ImEzQ9XogRBj1NFj
j3gZhxddXy59MH1aDAbv91/mSIuAVhvHWvWS3T3QcIq6A3s3TgVY593Vg1ATCn5A
vnF8keJZy+ex7hU7yLGEpZDD45GTBPrvO/XjpYmJ8WuhcOdaoKwVAXjsaooEumNb
ki7yPezAV5N73mHiVi64FsUcQcAGV8W1/WovvHq4V01cMPBpR9oCYxfYPua6URhA
tgqeoYBkZgqSx9+h6d3sDMVcWW5fk0pt6cjt9j52QjasdoVpdXx0fT8I6AL3DC4+
oOlrHP3ko42C3wfdU+SZdxc10GqjVnNPH4fi0y3GocAh/CmqzcP6Ysca6/1S45Ku
ADzMEbULkNLdbkty3AAPT7F719saCIPP8hi8j3jZjibnj4sLGXvj7cwcYW9ZhRum
kI9aiHP1LrynZpDQJhEzIuHG8+tsN2MZ9lNKcg+VwCjQMg49YQnjOFnSGjZOXAiH
qX5ei062Vamm4O4rYfwNq6+vatvQAl8i3WEDXIUsZDYT5TdrZblJr3XlsanRpJaS
23Au6P2DIg+A7G2RlPYJQ+q8YN77dHOIccR3O3AFZ1CpfCN/M1iobwbaFLQ8TP9m
uvv0WaFsy6zVDHtdqjAK6Qk5KOdc4z8MhwiOWzVgvhEc55RP8I6o3AaI3rfAQyIl
Fkn2uELSVq7+qHAyWv/SHdJ/+vciY2dxohTvQ3G0mtkJlckfcZqkGESN6xg+ECV5
WOu8KPIgC6MXY9WMd8PKx5sGKBfUSjVn3wFM2Oi6c+lnKlmOdhjFY+JDIeCPFVUX
7Wqp2E3g5UeZss+TMRhIKhiRSylaJVxfHBaiLAYCkfU8C5Oy0QTw1P5Ub1UfkP6/
Sk8XgG+GKDlqelP8J1ukxVxvb9UoiB9kh1ore/zYzI0RJwBJP4OFuQGOh3JxQUp1
lFW8iEC4LjM2UNPPi9zauorO7vGjFxmpfXRQah0DvTSytjd1GyoaTpvTFbzx2nBR
KShfvqHdj9noZ72ir8v4Hj65PF11tS6QoyqYGGZgpscjy3h/4S19it/1BES05JyE
hVS8LizC+YKgQ62v7o7Iwr0UhS++8B4es9FUSgS5bKAD5q4Gpxl3su2y0TpjnvHx
QM8a1QMIH36UtIHUIy8t5H9ARu0WBb9ueJjhL8KfTszdqemvhIZW4OMi49PHMD1m
YCtB9MeJX828cuL3kK/8hlPmUWLd1tpoujtZXF2dVtrQRU4i9NzDVXyrTZYvd7bo
3dzNA8o8qYaO+S0a3oNaHx6bKYeF7waRwSs3IbWdB7wXT0QXxlTkkxItLC4slnnl
//lxcPCA3F1OztdPQgCEKpUQPz2tliqJV6F+GopJ4UrOLHFKRlVgumcdKEp+XbXU
jWtoerrpBnGfi+Wr6kw7PdNzQqAaPkYvfVCsXxlbyuZYtJnEYaxjeVGIqfeHmxJA
E2wRv2mcSeGAdQmB2IUZbrYIjKkFJjPnv6F9Ior020+tGxKOuz0PL/BlpZV5tOoT
I1f1A+8p7fhmz7Up6KI0dYydcqq1o3HvQWrkQB2bvUrxLcsAXxPBgWBX3ZmY0hFS
FhOSYIMzrdjXQKB3SuLDofxXLgVOfTlvq/rwHJUPqBw9d+qQaBDDT97pyoqEwlLr
wM//YTFBBQgNuJD8mkxnboCEb44jYyEU6ID2x8TmHDIgAkoQgyn/T7sdoiipKrB5
6mtjetOG+v4JzfvJDGwlE8l25BC1ZwkuIlvBQvowAg5dBv6vO7fa2a1/kx7P0TQK
CRYWi4zvDSKSv0NlwAtjan96igUSSEr7Dba42MK8MVz6Ut9xUk+KfWnxv+6TE38a
J0QogIbwspbiJU3P+zoJMauMLy2P3Mhj+CYFkvqCSg4dUxhIoR3Zd1asUG3gtFRA
s6K31lnCPG51Wxp8f9topAI4E6PAw4baeecrtcfWkV+G8CXHBd9umjqtO4htIqvd
+YfdFWTQsbFcUeVqL83vyCp2KjCjKA19LmWuOkOc9D1lxR0VRR0IL/2vIqccMZOb
BoLA2DXEF3W8H8xsg5Kv6+ZmnuTqcZz5BStt0Z9NLKOffdxl9mrtn3biJGwPqvIC
mehUHu6Uqfh9YU2ThudV2HxbJjl9roIVAFRBHSWxGroxDjAub3e4xt2zi7+W4a2D
ihqTgAMoFC4f2teYVmxDlmxKOpSyro+RtP3JTTPjJx3cmJZPpdr4WwEBcwCTRkE9
XMMGWAvw/hWZJYGJGV+BF7KcrTbLocx9WcOnBYha/GtI2ffcVmgPvorK+SwG2K/a
USr77pAb0FcFet3MI0VDC5R1KF+Td4qc75DUCOov9GVOEJ8kdMCSCXJMd2lfmHht
RHYLB9Az4n7QGxB+ePjmlbBepdBNUgzNmmSC6hcwkuNP2tMmEWBhaYs86svCsUUM
WgTDYJ7QiWXu90leGb06lE14opXtJCY88CNSH8g0T54C2PQmdtE6wAB6nI8YaUjM
FwHrYBnOx51ugi2MjDmM5BhEWlAZvv32MZ1O9DrWkV8N8wROOFbPi5OjITJq4wQk
5G2oLEN5wKrDXu9F09D9yE360D3BY6hJruU5OBUSgWqQ+gblIcuWGUbVET+iybSd
TP6Fl4HbBD8ef+es2t3C11hrOBst7Nfsq0Ap81DRR2p9oMVekZxC3AIQjFHnL1wX
XrFZlizDTfgPd9H4vaorN0aA+WltVXdBTmnQ632p9NmSr4kEJuXEiG6C/8cBL7RW
N6REKvBmt3C89HtFm/Opc/ihxutKHtrzq9ylmliyTQ3X3XkWKU7Xx0TIJ20OlilF
soi7yrkcJblo3TujS1pLqv6mPehvn7IL3TJrKbLzi+0XmW+0NSWARh9a9qlFlsPl
ZGwyWtSUmAkXjyXCmfiLsM1/L3ocr7o8EFrZQc0k4mADQI72oRVoSx4bKTIcm+N9
wirNoN1vOxHzNMMFHCGtcIJciAD0f2d5QB3+ZeIl+8clCPm19uPPEgbcnYzfvQLk
XcfsiGt68xEWW1T3c5IQL23f1mgIPgfcFimDaLwyArxphJ8O+MmZlmy+zUIh4rfe
+J8Gs3HKA4V3QA/Z2vPpWiYIK9eoS2hEANh9QmJ5gfAevN8SNV6fzzcSLddYCjJp
tSPW5hWrBsO4F7qQ7zO8lp9KN08kveThdYfCtSV6lSvuhUl6G6W+mk4Jwi64exr9
6s4g1cRk83wvzRN/d7MOO8zvhjwh1JhgnTTWkkzIB6KemqcSDuCJKBqA0SzYmKK1
cVCP96T/Z1T9ScevJ/Un5OBX3eFV6nyD5j4dVk7Mo1Reguv55BoaCS5DNdg7PecY
2n91lmW5z6InXSx3iuh+BT1TVnWbXelwkO5hAyCkKoLRf0o1hRh+S8w3raEOG7Qi
v6mXkReK5J6YcuUTqSjX2S7bEN4Q4w0OHHuXaFaHaqbMAcbjja9iTvzuvvDyeFCx
UQBZHgPejcbw5ufzZ9ovwqOzoN/6w7xq9I9hYqPRLoWKVY8gH/lMUEIRNYfauUFf
ji60fdU2BQVhO0p+GtJyI5DH6mHS3K2X3F85FzaDg1u+kZEcUIDf1W/FohAqAXnp
B982y2w+W5ZJHc645GsoQh+m+DbA/0COaFugqkLnALgDUawzwJ0JnP3KMDNFg+aV
FzVV53ipqIpZOb1hHefoueMYBTfQM+YONpiwWhXQvD+P84CC0FdvJ4MHszXm4cY+
ywBtY+pC9hkrQ58WmS2arKKwM0YbPsN891c9Ndjt3jtepjXDuU1LAEEJ0QdU/5ua
0obGxiytfrS0b5Qf1mxWqLGzgmGlGvb8NBPgjqWFIVmT200va3Fw6PttB0I+OCrC
y+bFVETN5PZIsTofsxSeWbwb1e/tVOiQYoTQUQI7NmZTBvhc8zgOzi472w9HUxqp
aPbyj9A7Vx/GdL4/OIKOorLgi5VE5JkZ1LJBYFO/DDm4Uyt1Vau+VP6wf1tApYYk
U1r7MNci2yKQiPKeBV/eya37lw3c6AIh9n8Vszp8pWWAKli8ZYJR9iMjLt/IxgGX
rue0Kp+S/yFKzqujCx6m5IbFewDu7hFjB263nQk3Z6IkAUJIXbD56/rtdSt9Xu4I
wgVHs30Q5rmiGnOJGXHhR2TveavvgkglRZb9ubhsrBHw2S4tR1/xxIDDhTSbu8i6
bXpNaG85x6QzMz++IMqTBVNA40jL26AnDd1c29jTOE/RJl7bVy+pyd7KgkKIPJWh
iLwGuX5y9JlaaZhrrMLaea7wsxVdFK/lo4LzvPjFm9okoMD0Bwgjm07hBQpspUc5
FTkNxdzQtBXKZa0tbz1sip7qbKNgz/osdplb/KEhrdimHdfbMUWrWOVQKD+QxLFP
dNhpktYuvXenakp7D9J9T0S9a1/tsoxKFB9Lwsz2fjELN3ALOwAtd4M6y6At0WHU
ExcB/C1D0bPhLbzinOcBYJWEY00+oRwgzmZEpPwKScCjmepjl4ayrfr4fSeVBYEy
IQ/JY1/fyPLbdPSn6p+h2Yy5pQ06TJ205zyFnqdkothykP1fVC5rSg/XJLcD5Qhw
wZOIzj2f5VZNoJuE1bc5r8ou7lx8kSeCjDKvxTfX3KOwRqSu6nWbRKShm+dOx/f0
VswGbtOJXq62UpIdDLtV9tBNkiFHbVNd08vXVjH4itSPAlQDXXOIvFa5FLwaGNAY
TlUDuni/1NI3Rugqe+IClNCBr1D+4JHHfMk0K6lldCbQYslWn6oYxL38doN1Pi5S
7OIyr2IluuPyJffoBlZiOUsD8FAYu7fhsPlPSxG45Jqi9wBuDPQ7MMOQ+yresHi+
rb6eefi/dQwUlJhU8QW39LDy4llUc+emzzNDfcGr7cqf6Kv7DaH4+o4rdym/C2ZY
Mg/HtUX9FIAewdu35zGJn9Aw/FEVDt/q6VcpHFoG+ZWfwJV0Pi1rAm6aB1GBDCON
Z69a8EBOIejoozvv0NxYUHZpY71rccRTCtc80yo2eMt/Q5+80SzNTvSiIH2RYHv8
cK5X/sobGOPjSIMaSlwBkiaHTcujgx3WDWZWx3e6gQnnBEypmG0XzLWBE0Evzq7k
HWIEH9nhrV3KRhQif/zojZgNU2MmcWxdtwqHYC4cEwkL3v55mxMbK/MVx0nwOzCW
B3LMfvZ0Wvp9KMM2l+SHAjjX+pidUudx6FqnSaDGsSlGjfEdYEW1kWQPXuv5OQqV
Ge0MGDqMnf2ntLdhUeGtvuxztFfklTbUSjPe8PzGyCTzChCqbpLqMGXmcwxlKpHl
rcwoUCrm1M3QLEkixPB5rRyW1mdqjKb53gBfxe9xtBqI0++Vy5cPWkTAttr8PZ41
AsA2H26SwvlCHZ9Rz25GRKMYvwp9pYWtgLbpp/l0Ijgzr8ndLk3duCjl8O3ycDrS
5C4OQl/gij5aPxuE/EWe81077KmOFfsVBB/RP9hrp3bWPGb1TAqvqIfsu2VZvTXd
vEUziYOCIR/z8iteGdcyJtaPQ0Ylau7b58pKk4HvxJjSstnCcrAmls3oBhQdgHS9
/5zNdmasYOaeWj1XXoXMwe/GOZ7lakycbYG0FjRVRmypnJrcoP072myEz6SL9xCb
dz9eTPBevD0RBelOSdU0jsJP6fqaG+B5cR9JwgixPUc4/JWqKJgPujQz+qjR0SP9
XWTSPpCxNjk4gjf2CO2ufaQsLg1H4s6diFcEdSyIrNSu4a2W9oBSlt7aQ/XHrztC
yCYvp7ufl623+cdHrGx106aUPUFra8VSY2SN0BAAXx/oNfpStOkul2l02/GhAt2Y
srMPqREfe6q5Qq+F6T74t0btFpEkL/OUd+cJ7mL3F81PHyjXrZZYtiid1/Z1Wb3y
LPMK29m0B7k20ZMUzP2cBiv5M1RAoMjnl7yxY2ZLTjH+qDhaNAkYhwz4RXHS98Tr
upvO8DiNai+3ZnzS33hPiwqS1K0LoE5lvgy2wMYkLgzYjyXx5iobHnzpIR5Il68c
4bQ22F/G9S+EDpg+UAMZNABt84VW0PeMb6CWA1F046V2nbMlnJa/w0XnTp75QbuH
XLM3EAqUmXEjksZjROYr4psdTD0FTVJgPXYX1Hco7vV+Z3+sVm/JOOn7FR7+KSF5
4HVfUh2Wv21BUH1sXzwyP2Ov8RHRzRwQU5yfnMeoVdLN6lyqLoOxIpou08TinWib
oK9H//2/mzzxI92rZsS6ejDz57s+fQ1Igl45qNWn8X55O9EA2ioZYsM0ukqb/8nS
B4BKdE0zQexpp45zopOqxiNmgtw0AwUU/k5Sb3LiMqQ97ydjQbUmO+5pHBlqgtRt
NmV7N/8X3EYFFRY6zeJIBidWw0TtxSLUkRcSlp9rVR7KOP8A/iTdRmaUJi12fYwb
G6qENcTn+rgzFsrJbg8xo8pd+qB/AXuzAicYwT4qGqKr0yR90OdI1ChYwXv0OA+J
TSLSxQZIEyyBnSus53Si4+i8gXzHadpz9HPJGRxse23ilCsDfefqNQQ3oGsdF/A1
EQ5YBXnBjCtdyOK7f+xD+AEC/+18nQwGX7iTOHnMZdd4w+6BtEDz8MctDqHMcJL9
+w9Kgo+I2KwBpHvimhM8VLKk8HPRPHArde9//i78OVw1GK/FtUfL+e9Dv1FpqN2C
F24GB/PSXnUlzVsQJ03t/LIWoOavb0hllBhO2dOGb2ThSrL9btdx7VlQTvy/2fny
oGTRBkZgM2Cx60uDuj3SOS8Zvaycr4KeEtplLZ4nCjZKrhGl4f/YOAWrIezH+Fqu
2QUKDNpp9xkyPcbQsAlyIeWDipWZpFbfqDaiccjGQ9RXTcWiZHhksFCKQcf83tlJ
t6uONsHE/yB2Ajj1i1A4/KsyDJJx/ge2PjgEYpMDj57CyvOzZ4SdSi90JzQv2Ntx
9Bep+Mt7Ug8mvuU8mfHP5sz+38iRUU4zj069HDwT/AywJ04ewusK2lSMXBNU8Cdg
6RuwRASBHU5jfWqQPnlEDRGi6hUml9Hi5H6m/F7NgQFO4yq56/2pPOeffbK0HNCl
5NvQ5k0gLMSRQxEFtbuVDM+O1X3jDxk8/qk/7cnd8sc0Kr0iYJbEKh/kC4FfDWdy
r+bJYuOY08G6tYVscOh7XHqicUFFUFHBH4aRE8ZOALXl23JC4g/SekFrt52HsRlg
4oUjy/LydB5VHF2KG1XZlkjjy4Ld7jqQZm4uX7GmzyZRl24Ro6Qj9MbKAOkrBSVm
GQsHg29Tm4wH2yKUhKnO8GCdLD8AIrpcxgRMKn+VdgRTcCp1RSJmQvH/aEW8lDrb
BE//yrJBexIONi37MwfgAcd0wxdLZF/lMGDUR76Inyzj6Wv+cBhspjNxlOPwHfdt
usr+lU/6urn//JvU/4+ub9v+MdxXoV545auojUrtcaq3qwodJ5TRdHO19u5aEKtv
k8ocGaFad5QQx8Zr5N64mBPagkcBDk7ibOUxXosRwLjTG4Uzqvxf4pryqu9tELoc
3oIuSMTNaTvL0Ku8np+bla7952tMh7QEyBxxXc5jiwoqrltk8QaZx0QXLXCFn7CZ
lhQictoQO2wWU/X4X4FcpPG3J/UlY3Osq97+FZBjdmkEqpaOW38kFEOUszJLAxdp
QVyQrCreBANDo8omDqYStcFQT3BYZ3VhoDuigH/8HFAZYPDdTVNM7uIg14KosFhH
ADAbX+VXJoV1JgY12pzd8sz8u/xz+enzWwlWSgl27xRR//DuaZCgsDr8vjW3AwKv
lYeRkAwFIeQmKEWBS2UHTMi1BUkytMD1o3Nol6qUUHvPxYT7ydyOvYHZ7d9gJPrV
JVnlxV5RRmRNKh3N8FyN4q0nDViWf8ZsVwfbNCvRzlRMMyDzT3CnWYzMeWbpA8cL
+y9Pe0OqqfYFvr8IDWJFajjEyMg2llbaRqgqHvSAVTv46JGd4Mv6Y/+aZEPz/lbu
KWA6PiMroLwH1xvg+8AOtGeMv67mV31fXZ6MoRq9S7AVDiicn8EpFv+wAFofpMTh
DrZNef8HhW35tU1UVw8WU8+RPh8m3/7Hv5RAuoMyXn0F0Bd5dNBmaURbMoQjrQQb
GVzu0HU22De98q8R2cMetuowpzzqdHZYlPC8SliUtOshjidzkNpGtBihUkNoxrO1
GiWB92C3us4qkGLmsuKvPzjq088TYrMMubnA2GniR/mRGU1fxCN48Xd8cgBnCm0r
iA3rjBHktjPV7yIk0T+J4ieqNRQk7Iqg4Z7GetzyJNfvzX+WSTTuAVY5N6Yifz2M
71El2zJyrAiIoNkinmkNlF0fTLOo/viNmSYkow30As++cqLrjVU4jFqK99rDSjMk
bH51aV9WYAm5+USVaVrhA7HforMMUIhkCSuOw9x9kR5a/G2h7XxLRemzKOHZL2Lk
UwjtiDUWuCbIDKQQHjHSWlc4QbmXjINWGxbs8gZNidT+R1UTppQ9U4eXjLaz3nP0
5Tjvc3aV2UZWj2FKKa3+QjtjwU0EkrahqADwHtlTs9O1F7SP+eKk1Zv6SQjwwtwg
6aHyWN4mxL1f/gLJqzsMR7irYKir+K4QhThN1dIjTKAAoaDfYoJ9+dawBVufN6Oe
kMvQbYTqzBV0DPa/SJhg9FuBVXuKX1c6oohkHGUaxxPTDK4Rqxo2omCurfEas0Eb
l8sl37W+wfHITtRb1GdaCudaSO8K5GESJU8DxvYR6T1+qTsEN9TW/AhB40CVQId+
jCWA8/7nUWfI86NmfYlbLMPWrhqDi5l85l0zrkKDK4XVjxMzw2YUfR7W8RNs9D4z
4ewEs+X/O8ltDunw10dRnFhxbVEgV+yNrPo6mNuDXRkY8XFpFlnEa5eS5hiJFBL1
tIYjJ9mO1bvrbS6F1URhELuvi9TgyxH6EkeE5sK7PmYuCe2/zOtnAe70USSypRwX
zzkP0prd3D535y+IvCDy6M6d5NhdCYmgIM3kOlc5gvX+/nz6rofrZbqpBPYx1SnZ
tgeYA4u3abNtfLXX+AvlF4r1j/odhMmIVZk0m44rA7RSmvEdJXwg/JoPoLkAjQJF
SaCSoFiVFS+WUInGIrYIv6a+UFDVyAwBYerENcjDDJ6QAuHNmmzxDF2Fp8MiiOZ/
wlEZCZFAVB0V/HjQ5djzf4OVngiyvSv6heQ3Io+Lh7TyR3gP4UTWA5inW9PSBdtZ
7l/CpIwWxIQVPuMfSvKtQYtcxvhBag4wfUDPAmrCqTpV/8ANeBOzuMPskihgRIWS
iVlgBuS3lOAlNZQ24KQZ20QTFMxH6m1GmyMm9wJPWtNivGjnUb5BrjlVNDypIiuS
w4qzb51E84EHrszcQcCnzvSeN899IKGG1UZbRrFFWSxR5zVkKz9Z+bKBhv0vUOv0
vz50L3BlWgXMkxtslGOn7b3nRMVrggOfxPMxc8OJ48xAZoDD0SCcnu5KAy12FjUK
WGqV/HPuOuIHtv6Kzes12UNqosGMWuLqrc61WJ5YLnxwbQnJfthWkK4YnklG5jag
ty+DqEF8+tmjk/vhBO2zk7qgOVtz7c4ItSHAYYSa82lm/3E1tXRVDqVtS7hTgQAG
u+kfyqcxiNBNeVU5KfjEtjlc0rkWNH04DVMiuwrPtvf6YT805zpeGaESqWHkk5j2
/bU4bINDNpVgUbEF2G2rCjbkt70vphelrbdnXdIP8O/4PqK8RJfOvVz0ZkKWlI6U
1CdSCfpkJYd41p37P+tRckbNGiyLXeswnD6NdpPMUwp6d9ZNud7bx2HyMBMihRP3
HMdDrh6qucI1ZIp8w4qiKLEU3APzR/L4Dhqd0dQyocgHL7WagDPJ7Nv3I6qcTJYp
X9P/L/I1mRop+qU2MguTzjuxBSSk8IoGjfKTvx02rzP6fHgVBPTCPGO1p4zVSwv7
pqTPCp4qDbXjBQJ2FselACg1tNjmwqqb30fynIfJg0c4XiRuRdxgITej8x8AGiDk
XgQTyDwtsNPLNnyO+NLs/BfP+4rachWrJdx1QO+O9xBvGlWz5m8mU8BwlI2WTago
y6M78s64L7U5qw7a80M0ktxbSnabBXiocA0WmTjJwl9kwh9RjpTqjd3aEQGITrul
KuUHJUIb/z2juimYVjwhfBVbM7MQI5CSI9qilse1MbwNIjq2uMMjIH03UiJ+1spZ
EuFaD1G478JcJbwj+nVtzDyFvGHPymW4edxOAkqg7v4qZZnBoYon+9k1MKxF+9jT
yA7P4Lg5nHy5RTfSOi7HHkSOfWRW38OOCZu5k5LWa5IQhRuWQ5M7lUm/Qo8aeGxO
JQxc3FPpmacCRIA1OyTQL3Ki1ZEGu/0tpLvecpxC2ZLX9YltqJR5Ge1P0QzSVP7W
vG47iNjZHbeY1lpYKmIKiNSLzrggZapToZBHjeSLl4hKavmQIVZ8E7Vfqba8ALRy
nJ54o+CZNYHYZ7FlzztY66ClDQA5I2vDXX1el3k+HiMzYj54vS3ig1TbYyczzgF5
/BEq40toABGnVHZIe7aRVDN6UjGky7YjSRTKAWvj4Y+5iyNXxiMV1l1fipmPl/n/
ppAEYzfgHBK6PI1++ZH7r3rIU2Zrf1un7JzTVK8QS59qxTRYZ2z3i9IMWBbDITVC
2nrhYtnsYwMGzswz2ezbVQxy9nEbmB5r2p8PxiKL8YdL/Z9H1xKl4IqV2ws4qv/5
`pragma protect end_protected
