// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 13:57:53 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Jr4/E/oWGwXjrDmIPl8/QiVpLZOypL5v51vk2nZf29fvTgYtNxL+FNKyYHFcqQFI
pPKbURHD+2pdzwK39TrhlHhkA+AMWMTt8eESw7CxD6ZMRLcfLf13laiBs/AXYi3B
BUb5+EpQ7+6tbbMefbSs/MtGrTxIRkNRew0n2PF2yfE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3040)
IRE9dMNWhqsyok3QchMXD7JHomZb55Jy5Fd85WYH5E40J9Gr/URLj2P5Npr7ftIn
twaefSrexxa+vCOnc+viSFcSAJ+WHJx68Jz630auEZ8qChip9tU61fI94DFtKwbQ
2vr5EqToorI04kqZ7Ut2uGXM6t4gO3CW3YOPRkNMNKAA9rvV4BoPoAGzfnAQnjVp
CfSmI6E89njG/Yoon30rv67b0zj5bQi78G2koEjKkQad3eDdfsL7reUv834p9cso
C16LSEBkXKvm4CR1rK2+H1fAnUQUSvobWrJBxSlP1p+UkiLtz8BA+dzMjff5Qzk/
47rJrOir6dn3oKhrLiw1FomSksTtkQWl+JA6ediX5Q8Ll7li0KiGWVKGTQ3zbF9B
FzuuMNmDyETg9AA2xH2sNthtxsX5HXFLdhikqpsVd7/RzYvqKy2tOJtbcLFUHNDB
zxuQOxyG1aqXZp/3Yiuf/CZrhBF/RejAFmT7EOfnMY+eAIUjmDVag6xpwR2wvmpm
hWlzyElseHhenTQ8DZ2HXtzV//4uUMldFBdAWhhAt+Gw/+YCpdy28Y59zVaSb9rp
wpvpF1nua4dyLGZaAMsphlRejywPw/cy0c4dDkTHCHY/JnDJtElDjb9LSRLnyPMY
nP5kFEmJsH6LCMb2jzLk3TKVZjGUy8oi6lhb3wkz5xTwjNBC+LDBQp70U2VKyjZz
gsYSaBQo3saeB/C55uHXLcPnbGZpWscz5eIQ3HEFxOz8r/s4bdWYb/+u9HKbmZz3
yadlDksOO/1YlzgH1lj1wbc20tO73y3NQNMmvK1kdPf7Gl7E0sbA8bQEGXSWmWqn
kA6SRAyL3kpCFQlSrWh1a5WUYei9yLCfb/gtrU/1VxtOGseSr/VuUewRaEY/3UPx
fU8j7AdCnHKZHHdGMZynLQNcPwoz0995YpCLxtR5DtoNb4yMbUNll0/pyJwhZ9u6
x+lxZnqfCzEVPMvQbHS9SVQkDYpVb3ipGm/V5JGjyZTze2tTF3P/I3HymzaOSj57
O3TVWpv/iJvVLE6LbgtkJvxBbMcO4JCV7up0gk12cJiZne0nmD7h70b51l68Ogbr
69ZPFwiY2O590r1JxmD/HI1em81qJ606bSS2lt3ynSEd+6N/KUOtO8hAygRTML1X
HLlHsdEQqFGfBFT3idIr/ZTx6vKGRbRzzToBXtDF9w/wsDmUbk29M2jpjegEPaFu
UHglFVLOManyL44rUT4l+aTtXJwdX/jTc/J305AWbig4HAPo1TJH0zbiq5MkLwH/
MA6S5PXggoLLXAq35qjjOsAsbvpGeH3u5AHzpEl5PAMKbNHlIUxbvcO82Vw7A1Cv
g9GQS+fXPAU9l6x0zrJ//O/rhAnEhWzcvSJ958a0FgISQAQmikm49pfU4XwDli42
YYdtg5bt0BcIbvd7ao5pOktlnPqPxneaC8pl0vc764mHMTdNBnWBsCK233UL0SDy
yQAHVjZu+TtuD/qceOh74qqIslGz32Nv7DEop2qDbMum9H12AiLzv0CUHiWUqF4P
SV8lg/9CPKxYiq+r5IMXQW+ju1ju8N7u7IInGGZWahqOS/ZA9NuACtPWb0Pwxf4N
bIeP4Phwl+NgOx6rdhhpmPh5QA/y7xBUC4phhbt8i+kzzEm+L23QrZdKjP60p/sS
xcsVtR/UyJge1eEilcz5ym6wyirWF2IciDc+qvKaQpTYdk1ZS059kjUipa9wilyw
Ng/SwG8qU/IWK2pHXQL2gbFjsHQvgAbWZsaQt0DGvODYxF8LFCdVxKKK0ESSdIYB
1EsDFkf3JvD7SJdJhfMz2qbitti7jr01cPZL+1q8Rxnh5esIBR0smWRG+77coD9K
HvXhVkYLOGvWVSu6K7UVLqyYDdIfmkimGwHNueIVl0dFaFCm8zflx/c6KMKBHsFm
290/RPFQ6GtICVFdRvGOffNn2mjhhHfzYKaw0iP3g6A5dg5fR49priEUSfiHmOb4
eAHH/nUxVIzSfh+MLjlyNMaYuiZJltc1fULYnT0le9Of//IKIZdhcULjPgfMNgVi
7iFqXV21626I4u1vs+/5rpMDdugexL272WcJZKqGfG+4aNDOpJI2zMLdg7/iM29v
ym1JW3rS+skvDveVBgbmzOQikXFyNEwh3/LCEwsCXad/4cfe0QZkK4krn/vWEGFG
3+PGG56mwDEc/BHvFNaY1zGBbWTH1URlhGpHTCogsE2tYu2u0dts1l58zpdvKS6B
LGPGZ8/SFSQP1Dsf0QrjLn6E6GU92lK03bAk/cVhnWh454AklXk1eHdKinSlNfJR
mqrUb2sw4fu2CESio/l2MNm1W8YOOPSyyCPFP6yp15Ds39XBdiIcM7Jryc8ez84V
ihENfg4Ukn6rKgGIrXJGIY48n9aFakV2nyy/pJzzbJ8MXx/KDs2OUPeCs1OAFwb1
EDIEzn5tgkk855vIRrUB4JEUXv57Fm0U2wid3e0juaSR7YuVL97mGfoI4bxhAJPI
M5fcAEOvLpAtsKpSJJ4zkkwjql6+ExNbMrgWAJm1prs5VY9/g0qMcoWtPHD1Buo8
I8uNnhFlwhOdFSeGPZAaQ6VC9tVuoGC9AW/qscuMoNZBVv92ouLqsXvd1V0DRPK4
PmZLdO66rkZ7G2N5g5KfxDIMtq7RTA0hgPB9cR1dTKZiCcesoBJMS1rXFYfHOVY6
BT3F9BjwLNqitr6AQHzbj+nXU/k0Idjygt/cyiKazkJZFaVVkngKBbkeAYSYW4hB
fez0ULdn1v9jgcpI3yE6FkVvqvUUX51Rzwxh4bDBCLirQg9ra93tP9x0BKSW1mCI
se+au6YkPwU/9abpw60qZ3o+B5UIuXYaTz0xQ9+5AQUCb0k67xsfmh3Q0LJqgKRj
zd+0+DXR3+nRb6rFGjiFnXbaxy0R9XLu3x1RqzgmDmq6/sGV80td3MWmuvMdI5xL
y1JqwRo9/maZ+rv/x/IScmbJz659CIlUbCSXnevfJtwWmiqeyHV4sppaOHK2Flr6
BMrqvfZmK7mKiXTdjC7dLvwRW6vn/oo34aYKQ3v0wpuTguc687l9Bqvl411WXcva
e85c0zMAbUdDunID0OJ83IoxDL3sSRBBmuYQEGkjbhSxxKEPtylk/2fndSqVnxaz
A/QY6+3EXCRm8Ki4QNf38miFLjN7n16mfJTrPeS22l/0e3du0QEHb1OodNwwFfqy
UZD7KFtA4Xc1ofPLErPrGB1QQyuVULet1hJCVSoJIRiZPj0kwCFCKtxbTasCSxrP
9j7POLrb9gjbm46qjOBLXtDcFnAGKWRjppmVrVraHrwy7+eyJw1bzq6P/ULNTqG9
rNQdcUlNeMHvmAu1R3mdRpMiFdY0msaChWiW107Zj9AkcwSwIR38f91U0bnoid8p
f4NuYt4S2dl5Sf34wt1eddgdbTW9CfreKvdp846nLnRAvMCTdF5BlyINtAuWyDB/
rbpA5qkUoysAQt8i5CekezgGv7u5yVTk/rUfbtO+9PuMhXIQUsJxSvNSDMikE9U3
QoAthhS13xNNXKHHEhFuqLzD08mR3lZTzPzuseECF/zPtnkF6ZP6wSMJ3hCJxV2a
eMueKbOaLC4LvaoPVk8Mq9d6GG1i9tF5BUnawY9emwACFNXTt7Do5pzSwfcsekxk
s0XOqqsR+yWDNjJNykjXm5ZK6NTvD8gWu74MzI9spUOF4Q0TM3ExTnx5gES2Wr0D
zsiMYKTrFZWfsFh9ta99V4IbHZBkUnfsq0cIfHoju3y6Q7Xk5GHQBjNAULtVfUi7
78+lfGDXiOlYjEmUSk1UAliUzufaMq2JGGTQaDo8omYgNA8q4TJ1EOtIaslZasm5
e+vIu1IjAYTk7JeB0vT20EaDlF6zi0dXjTBY8h6ogzUbd5MgYk0iGZMroMejbnu6
tMJGOsuCtwLa+6ZwYklzI/mLShMwDu5pQZyiWfdq2h620Otibh0DF+UhoXuaR1MI
qbR9NiVWqeYqg9y7eahSNtieS0XImrpHUUsmDDDsZqFo0r+Hd7sspALUKJug5o0V
iDbrWNcyZlRjJ+3pMblYig==
`pragma protect end_protected
