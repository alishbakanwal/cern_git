// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:29 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
n6HM6gS1PCNRsm2dPfOGm3kiRwCsTDvfXnulztcTfu1vtu2Sd69nEEDTAP++w98s
0kXfABzy2Zjjd2yY8v5RK7dXEKwtgwU0poT722bNAV3shiRBfQF45ntrSJDDf/VZ
UdMB+ja2aslzAVfmEOqbAdefiu/AnAQOUnKtrtlfbb4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6544)
hLjFykHKPVNIz31P0Wx82wkwzUdY8AeyIxvR5nPJeVlulAFMgbnUrl8EfFc+0w88
f6PrQ/Xy14jJ5hvKF6GcsShBuRLU8bL1zij7Rej94KzOyRuIdclzGlHOV1Uc42k0
xJ0tNTPPR01wQAhBXxDXyFhOGl36/SQMbmOFDs+hbamp/yTfTIEKUVcLq4o9Qikr
iPUrAIcmj07foLpxQQH+nC8/mcPHZY1njq0qfeZZmLvnRnWx35vVW/Q/WXjfpgEM
merSzjf6wc7ZIHhmNTWRWLDwpQOVX6ayRDuHmbLPoGn9u4Zmg4KwSU8BsqfQcF57
+fW++Qjva/uChgk7FBkjnkhJxJQch835o3Qu0RcZr/UaWu7uAZIcfUOLRd+fKRro
7MWr//6yxO6zJSUTH0m71vjhk/Iv7IeDBk3f7kHujS9HrYdMz9XldabDciQKW+44
kq7lx3VMUlwd+BQXl9e1UGS3fh2STCBSWoBT6nYAaJUxvEjPkNAO9r1qZmUCOHfK
h+lOIsdS9C+jwCl4Y5guGkxfj7Evaem+/3kBDUd8nf+uiB1RUmRQwCCwrEB4z++i
N71YTvsB4TKpCvVwOiGiacFd47wlJATzOBkgpxUKBZ63PTRbqzAsTIpN2qNLg+LW
FAxZnm5+TdfhcFt7uewzcJpzvaQRNHOxudYnQ45jeVWKyN3LKeM5PV3jlb7ZTlXq
MfsCzNqoUkHQwXvQI419IzfFnGZk0nVyPNMomBwuycaxxtv3Un386k30qJyfYQAU
XWXezJwexNYjMMn14IM+zh2M7ZYeurisVCBQhfV3mfF8Mt7dVnmnwwex2oJrPX/I
7aReL4zmWcaIb2vVnA31BX2S1xk9JaXa/T/mJgqcRNvkp4YG8EXv73ZANXpkJUVg
GHKRpMHl3gKqykCxDensh3YycUi+Ftx/BUhGDZ2K8bOiFsEC+mAeWT4A2DYeMjif
zTPPEqejGDwvE3ry/8uqNRmUIuLiOxBu5uCQchM9zZ1WBRWg+rS3SmX13Tvjd0Ys
c41M1DqclJ7z77sKp/LEQkrVfSjtNtrlnl+P1X59yg4IGY/OSi0YD1SQxjQescDm
aHywN9ZmgX+2jFHHSj4QgNa02UMrsd02PyIClpXwZ/TyWs9ynFYVta8ujgLpvsEd
Pgzq7BlQUBiXQkOpQmJaJt7P0aAgVtYcjW8VKbCNlDnJNwgaCk2glN+OjhmFCHbv
053sfU1OIn2KH9OpJkC6gfMt0eWAw4/gVOO2yMNg4WNGBX8c+tvcG/Bfg8xA+aKq
sjqLIA2rj1D9ugjji3xo5bR8sbwIzmibIw/qAFjeJWn/P18fpG5FGfjVPK+Tcr4K
A5/j7+Zz5KB76euIsU+h6iKiYs8rO7GaOMGLlRijX+k+xFxLrFrHWTk4aP0JjoTG
r2af03Ycmkp33pZrmi+0lxovV/zcTZzAoBweYX814wpjHq/dHl2ihtxWb1O3fu4l
R5YtuJTs1YrAj8nyxRMvX21NY1kdznUK8VsvHOxCdYAcC5DxVBX6M2AF0/hyWnI7
QgDYq73hNgRSfKFqSJvr8u0XFzB+JNO1WWjsG44fBZrpBZKIT0W4sst5VeE87tqV
60B4wFpC6mVMBGaioJP5VW8FkhQwDxtECkRz3X2KMWEKHhsHYNLzIutuIffXUCRk
Ga6DW0iQJfcQgYShEUB46wpARoReDUirgcv1W3LQGFZs+yVCKzTZrMU9p07ZIV3M
/lCJDChUuU+F4tKEN6KEfCaCgA1+Fs1CNt9JW+kzeQzag9NMcR20ajNO6q813HtE
hmUotYN/kI/HBBlDGTlycJKiQ4/zMDWjrfweI9QsXnT6IBJSEZUt4UHX2Aj3RedH
YSdR7IIKMYK9nk8DuwyU3pQUH9fPrAMmYxenWGWRUaMw5ZjHOn4gdjbW++6XaDt3
XI4ChD40D8fn7o6u6/dv0XMw9AizLUGQlSogEE1NoDdMk9KoblGEJh7R0fQJaFFE
hemnU6HMPsivBe+DVJZ9DBtVIL9B+dgI9SlYszxoZGbcjhYgifKoPS+h/SX1noCv
ZcT+WWOAeOtqXkg6/c0LVt8L/JI4RVfUG6SHevjiMPxZJ4cdNMEV3jPjn4s5ayW6
qcDGUG/pI0+w4GfOYqBB+k099E1RHtj2WkTfL5CDK6QLhrx+lbCgx+ROw108GVws
bvNXOch1MZRRcthlmGz9UZLGUkzogmuX6TGwMDj3xh6DUGXbPfoEwyZEqmm8ZCa6
8T+CzKEuoA2dVMvxmZRRDfGptKZnZe+yyFpyW7aUaDy5IkNWO3lWpunwh33Y6/HO
tCOo814e/Qsy882Dd1Ssvb+BxtlKQo2+bGpqvV1WYjvCEBAV1ojKDijRzc+pjMCP
DzqoRxXOpU24s4+LBqtESD1Na8VqnFjViGxgUFanmp2pcbQ6lSsQ50hcvqkO7ZZ8
vxXsvG4d+owep5eiiSCbv2p7lhaHIUxTbevsF+ogFvMa0yxWsTsNuTw0dNeZ1A+u
Cqx9TYIEngHQXvZT5qhncdnQb+yYaQozVM5vN08ATyO7865d15iaJ9rFq74jUG1X
pJX6ZSqz2s88gI/i+TuWVgWqiJtl8et25Dz8utbk8+l2hQHtZWPmzSjmmnOByK/w
prPLol21vxV0iE8Q2LLKIWIJeoE7Ro/FUpnTYikUQGMUIM67ZhtcYn4Le0HRT9QB
Dy2OuveXiVxbyzbaW1ikbqjv+HPxntBDk83NxbAA4DaqMHle4P7BFm06UMCbmYq/
EqW6CSZb0OCMOI4yjW6CKOcIHnvGS9lwkZHgOG+ExE5vqMRo2ZfQSrN6kxJPxvGl
mOsloB8YjopEhYYiZCy6Kp/zjFyQ66El2gsksu68atnSLkVThcvcB2VF5X7f90nd
NyiFsSGjvzhzAh0bIBjk0eISlZHKBMMAE6QBQ3MQ3z8byK70h2h4xX0QcNt8cYBb
jH1Yy65DCiJ23D9dPJMMatwGYRhUbNyIjrd+uv0WhE00Emv+t5LKT+8/yGKIInHY
d5tZ1zJ8cpuvYGJ4R+syfRyaA13z52o0r3zHo2x7lXxBn24rsrTsCmwt7pgg5hrB
exCGrWhQs2ybY9noXjW+7ZynO/wshoZRYkNKlYidUWC2zvkVbRrbyy8J4HD/WDK6
KYs+wYA3umKeMIGC4CvxP9vSP6zNM4hhGjmH9U7qYORMbOXhaDGEuIuYO+3t4dxf
H54joXhaVGQ5aSZLPewB9WUcq/NXUOuac1cfVURMVf6HCin8pTvrdUGMzOZcN0zq
oi7RA0/NihYw/gLXRU0qPnpDaOZHaV+5G8pDs/bWm/gJTQoOITy0HE3I1AZIKdeH
WXp4dmIjov9p+wsOS92qs3mpqhUN6/FXpVQrbciGeyHXxTx5GOyErH1HC9Ej+TI6
PEIvmJPpwcu0UujjtmLNA31C8rqqMx/mNyLNHxoUZQpajRGavmq4LphensPuyLe5
sIssHXZUOTx9IVNqcD0ugSS1Gvy/a2qINK4gKmUoHC78v6cMWBVTNe4ViCxFYscf
e6hw+AvoyABx5Tppy2xMX+ZoK6odoxhIPAcPrEyPuE08U79XBPZV9eCVN+MalAcG
oGfvOsH18mnH/4qCfbp0nIIp/r6RyrCEgjKxZ5edXfCRrsPNJWCsxFerzDDsUgMd
h65TbnPf3xZy+g2Jg2sdV9h9eOmdNGc7n+dAONbupLf4upGpVtf4N9QBu44YxRs1
VL27JyZ4jx+4oT0tItD2udQQGxhfqd11SdVTpjR+biVc4OFeRh4z54iF70ILv/4Q
k5nBaOgvmFoFsc1gMm2G89h6MGy1eQ5HPavBUqiLtfeZ4FLt7fz+fA8ItkvMvCxj
dMRGcFyJDaUWk9upj612BzZyUmgMONF88R52AajyvwKAGTWxu5jB+wGa2pCPliRb
nSH7W+kN7hr23NfzE9aI8xRh991IUNGJaU9kSdpq67+oQUZC+Z2RLYTLZ4wN/E3+
rXy9nRHw1Eec52JWmLP2SQOI1s4y+KNUa6ZAbQqHoVHXH516AJ1ros9zbYAO7cik
VGZw9Fu41D1Lba4cfjrbeT79NWF6dmsPtT5i4Dl1L5/b9BWEgJz2abqDKcrQXlF+
gY2O3G5DKNiXpOhVgmpZOhv+WNSsJ5nHNkw78ko94y3ZLe91UmonjgHDuxD+2GBZ
xuj+ueNMPo3D0mfOrc3i2n0DrNfszv15Fi/it3R3vwyHnAkD7OAMYmpKS3SpR7qp
Ze85jg0hev1fkG0R/nE69LLiDTnQrNB02ZI7Gz4brGBfFooJ9e3ST713YA6b76BB
l7HyrPw2eSk95xKaa5ots2brlDr3EC5iZPnWU6xLME9R+FspqLljJhV66NVUz6vU
zNB7Af8SHz9xc1e1FofuuCH8+nmNh1CEbz3eYgobGAym3gVbCEwyYeQkSj/SNwBO
qTuO6r97siNd/OvkGmzpmoM8+nYRzxUPFckkIcWJBXLB01mEF1D+naki/fWRb7CM
LatsMPIDESaHsaPY4MPCdey0PtQV/KOQtHxM+QT8Tm/teqD5pbBSsNisovMbUZD9
d2sEgRK1jdpk9jVbcZKNbX8o8THLWlsDzSfZX+qclA5+chd3mXQjDRBcXFZZ3w5X
BKgoNJ8yCz3RqhkVIlDhOlq+fE6YVVV/M2bbPcDUCVW221B1pz4zQsQCL3M/8+o8
ZSE0YmkfmhO+JOLalf31bdHsIej3raBgHj3Jv7iFbwvtTz1jVK+Oto+pTcp6BI+R
bWCM3BGcrvyQlMs6qO6NIbyCRuyYFHisqHbpO1DXXRQbM44BINRLW9YZO1vNVIlX
jr5H2ECf2u8IfOeDm6Hr6rxzk89yfIrqWtynD3SRVUrKLu8KZyeD1uHT9MMwE//u
o7VGCqwJZOZtkEkLTUbjhVJkjnGhc/PP03r/BAvNV4XI59Wojfe3+LCW94Y3nqd6
yEsChWCyoUB9+O4KBm/3tK2nDQ6yZbp0psoe6buUh6W1RxUBXztoqLkUbc0Aq2FG
RKhvPjpKAloLUoJmKdC29zJxCVdodeCECVyYsMkDb7HQRWS/N7NbECyR8toLu+tv
aJGPVS/CAWGcj8VFP44RIhuWZZRHr8KMdsEa2wlJLm6VPa45LnVMqsHLq5HquvSy
Dw9RKhWWNFy0LhpBX63reWv6IeYw+Fq8EI4fDoy7deqGZWGs9u2Man0Z9qGgH+Jw
89voiMWwiqnoQqCvSk2zkjK+3XCcUzAvwVCSdeSZsE/M6jC0DpX6OICzxaVndWTm
/I/tny2quJrs5kYJCSh+h02y61S+KjtKmjiWlx6tuNBJEY4TG/fXhfyT8bWHnq2/
fKqAXFbP62N+yvUKSRrL+SshhymUcvYq9Qkc0z/buz896BjJaIE40+Zbt5yL+QJd
SPA0C4zphUtlMngKhYNGhIhs6P3oWkZe2pqoD3kmF2Qvy0bUMBUSicuihsDrRfd0
FUwMewSS5rHih4m+xi8gCR9b/RAXyOpK/hVPiP6YBiFRDV7szQqD874rRBwqhYbV
llfrYLa3MOSSkhUrL/PF9NFb4m/qB5iwC21CbE70VcAAd+Tjpo365JfdtMVdVZFu
JWOOD9ptmtvlfUIip4WEaHAHIhS83+kC6PMgy34tHU/gTAhfn91GqG/ZaIuhGnWZ
zF1s8epfmx0cAxfgFKtjK1xucSy0dH+tbw3NBn+E4sA9VRpQMmNqj8U7/eiHjpyP
cSQ0GUbCXB1Xij3T8fz9xt48+s6DWQ2TKdnvHV7CUsBAQhFxVU61pyyzYEawqsSU
4AYROZ+z3+mddkwe66FmeM/3ScxtQt+MaRy42bA5SaLPiYlWGYaqjgzP3Pbvmpo4
HgWMuSq7EYEjppk57+Yp2nh6ziwAhLvhMSOG5bVYN3AKIC6kg7s3dk+NRin7Lmoi
LYOfLgg4s7/AFso+HndpsWY3eE6Y+dOMAulgmXy5D7ay+AjrAXDldR8dt1MqDPdv
cldHp8S2flvcYK+WqX/aBNgbv1qALV709jm5Mh6/1TgIemuYGQ+EzeyRfMtNe8Ss
ojR99Z2C6Ac5RGMh3qvo9B49BhFM3o9KvbSL5c0wCwPJKJ+Nh0KzjyUi3xw2xnt7
s3QK3znAJ3qSpofrpxIlDOIECnox9GYrx3SWVXF/L0vzsVXZncLFmItCyoQGlTQf
LGecC+qJxd/DI70O87BLwaSB4W++Fi6U387kNd0IHFvSzZd9mgwJYDhYST+4JxMZ
itrFjzEO+1/u3dd3EpOj/55FO7KNAnXhITUBQuphM/KaY1+Mo2SQNYzLrTs0vDDd
Xr+k2dVgQokXL4h9EYZvOKvkly0w8hysn0msCuPAaTP8tLxvB/nfU8bXP60DYHF2
SDNTweOEiki3pov5F5KXjhneU6NQRP0y9f9caMgFhmLK2cWV4LFhBnm0EgdWMqXp
I55esTjIc1nk7MjJikAp6lidcbA+JMNxj7iq43v3d6oDHpL26HzY2saIZUykgEPa
GlhnonMZJgqru1z8k4VHdxnhB4zFg/vy3GpKPtiIbctzcNqbWuPMHa9YyjXhrDuR
7HkY1xtbecJbanjspi6Kspooa6smbmkhLgK50MqOjy+jbO67irYQlhFqxykIuvCf
fsTFuqr1TsyJu0nHfWMfMVm4lvX1LCPV27iJ1a2+L/8ZtST4dyB2Uxq0E3/5mbPj
BBiS4U02uYf5ZOkhvG71c2qfah24NRffRaa+k4aKbKFrm4e1vd0XDqSvWW+xMai6
3RbIHdjN9BSiVqQ50Ewm+C/3qFeLY5pwbwrSpYvx6t5FNraLP9VAW7qtqIRd+Ev4
q2gda9wl/4Hu8YeHjaSkdGwCSlXSA8ONiZbRMtNNSoqOthg48ByvR6aGp7942SoL
A2sHSzofLMfXsPMuBd4UJ5Ow5zIXu6cXVQtvgdl1ZPTwW2RT/KwTyBtECtSuXQzh
jHU9wgMxYtkIHrzRJ3xXPXgbZshU6/NBouHY1ysZtdem4un9o0E8VYwC9w5YXoiC
WSrz2btEEhz4buRclfZiPEXqsv3RRjfDNTmpZjinS0lelW3biNXwLwVh6c4dO7X6
jZMZkX4sru2VgrP1Agfz9AXirldbkMZLU1fWMUNGTdtXVy3eklmEWNv+zKSdSlM1
eg0Ft6z/Bvky+2x7sTMKPa4I8RIJcU3I/FbcZzUPh1G1hk5WH0o7syCAj9BdpBe7
evTPyQWDO1OJV6nXKWJ73mkEHzUJzre5vRFtSLgNIxGUa8LW5h1LS0EwJsnNQ0ZE
PKyVFPpeoVmnq3B+CmW/5zK2Ep0iFD6kB+NIDn2rwd7smvDknnlYmnI4/ZoEQnac
uN0CQr7zXw1GeS22F9cgYvgx6zN2XUXuyJHiVLANnw2Tle7T4hcEH7HvdRjPzy5S
khEjKf3JW0jmFqR16meqFt7qWt1xNzwmoSOByeyJgymcoUY6f7xU3NUisgrtid44
hSvrf51pUrSkoX/sTirPc5xhTATm8HxlDYX+eOQcVebwZS8FC8SoWHn69bNuVfqZ
pMJMipV4I70/3Uk4UHpM9kOb7svb+5bSu8+yfXTL5ZGRZS8gxzqsryDcnJN1dslz
CSReRjaXo3rCHtyZE3V8m2jtqCKx6KQOTKX2UeKZr8xzHDhZNAQe1J1tD6Zb8cxh
q8su7kAKFw+1wMOwReSb/AS2BM/gsf7SHzpG9z66FWxpa2WHnmOQqQqLTcnxFoWb
TJP1WC1Tjdagzooqc0LGxp87EQhlkMXa/slR4RgwrDuLw1yX+ZXfKEOa8EdMLzwh
0I9V48Cs01ReR2XXrDhyhNvaeO/MLnhg4TiBuyWVIJ5P2oxMLxqiA7T+V3PCXiVc
iFNxUEUkkVhT4aHXa+np3PqJ/G2PeOskpNoVJbhK7bwAL21P91v3H8kMtziupEpL
/THz+3rBRs3k5zxP2b/cYAhGy/553OWI/8gFRIPUH1DfJmmhHknZogVeoENr2QYA
NgbUrv926BnA6+XSsi9bNuPr1iRuV8MGCVdpRtko/oIm7WBMm2g5l52rHzvy0DnW
5mb9lSc8I0LubA4Obln/7oC8lJmVIRojhtEjjSPaYRmv1sdW0vc8HcY4HJlPjdqT
SGvQKbaH/QWc+4VKbJxliqFq4nfHthvbhQLzgrylP/XeOr5Zg9MTAnXBHwhqS4rr
ubpaX4Q3lYgnk9TawRrWusQjqA0FYdJiPvZbNZzPZ17uVrPMu1Us5IJ5f42njI2Q
jNtF7lNBmQlfxvSCccUjV6bqkaxzC/SVEsHsr5zPqCEp0efIgNdYhVh+cR245F8s
usVnvKklFA3Jz4bhL5zDA8Fu16ALXI3sbBkQFt1MnGsX8hFs2UYBw9efz2EAVIHF
i4N8a4HYZ9NSn3hN49ubtlu9qHZksUdAFzLnUqmm34MLvkNC4nZ2Yu2EOD0RRS7f
JoD1M27A29EOFpno/EXTedZqwhtjv6g0kJBxPiQjhfiDsnGWUPOSReTaQZmuXPMe
0u7Q35bo/hli42dEyWznjKKcvv5hWWToJ+N0OuS+I3JwMpYzL6GWk+jt7OHUxdP4
hdM9GM2DHZ1Pt6ycPDENuov+BombGelBGqcDSST857/zXAxj06CSCaeyaMqs/M/Z
v8mKLgonHZke2rRtiGhYgfep8RlUlpOrnN2/tkUw7JsYsI9ggMbSVxoi0IRyRt8c
R32BM4U9lwMvE4nf2LOQ89T8UsgzCCX5tTxYOc4bvH/KFzhdBjQX2/3T//rfWKvC
0W69pG7suA/n9B/Ffv1ayA==
`pragma protect end_protected
