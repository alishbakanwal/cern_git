// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 13:57:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Sp30udYmW5jUZC+NuC2ZFXgKW+RiAmraZx989pgZeQfqFo/yL0sS2UrABds+NWUu
cnSDajZM1fnDvwklAIKpSygp1Dc/4A9n8CB0CmY2o0TxJzEstS5w6hnJJNv3EATA
rliLsFbmRzsm5jL90/Gq7pSA57mLGWg1zW0OqxGMPXA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28224)
4EvSY+hNSyqTeWX9ibzeYaB2oBF0YjXkrH843yTtjk6+zzmV/XkRvgiJI0kxn0pS
vIfRecDMHydlBuqiXr7psd4cNuLZpwodDfwyUb9j0CM595oGw6aQZEGTEjCD01Jc
5F5tGIOCy1vm3tLrMI1KQYB7JlEhpWnPZb83cT5PSB32/6FabmebhLaQGf6T5aff
KBEH68XIRIYf0g7jW//+tsDG1D4FZNU2tsX+libZDvHh1WBG1gnbwe65JlL0UIl8
t8DRNLJZCIFZYDFSxqpGNQ3j0JaOG5boDBo01CHZ/yADEjNad4LvYgb3L07cKEp8
PExQpbVMjHiUzKZstcVFZC0M3E/sLDyhNXb/gM/yiMBO9ZkXyCeNQgtX6Mz3XG6Q
puhTbE8XDI5Bxh7Sy+a6tI3JyY3owgeTCdBcD0x5CMhPSkox5Ki/T9wU3ilR/cGt
bUBHeXRroW0lp4IL4z7pPTn6ZRG31+/p+ExJpk9yy483+B6OjKcyqKM8wj/0kJJi
pvNLm99lz7RzbiDWg5Bcx204l4bG5J3SHbz1lvGCSByktNUilM2E9wk6oVlmcoTy
lRK/L6drHVObMt285TEVO05mFjkamFQxR3AcpmYAXHqNlYhxUlVzYXGfyJ9pOR1R
iIzePjbHy0WP0iGQjeoVZ+HegKYpeQIZ0rO9lPvtQFTXXVgpZgalKlSVYuVFb5xf
modCGZo86YJUdNNYxeESUc2DU0lE6oyBCJpGITn4h4MG7CY22AOXerKYZ3VwFCEj
NQYaqm+gXrk6Js87CGAR3di91EPswVuN55Upv7WkD/1YSaGgAdpjEOg+L5ZaBjM+
KDHxO5Zb2ynSW2N+qyG0Q49/GyENnlbh0ZnRsFU+AZr5h6ge9O00CcLQsdIJih3I
E+3wABcpDGLfGp2jvQsXw7zzbGZXhnBRkIm1pk/kDD2aKBOU+UDTfNmqPNbpY3dL
DI0K+z8wJ+80y5toX0tIIHXyV84g/LpfaCUOIy8iLyZbfiD4nZP0CUWLeFKhX02K
qsN0tPweG1mgWepAcawDnb3jMWRKIqvuBa4GSyB1Bc+Noc+YU8xtW8AMsLndttIf
5BOYgXe7oSoOL2rFxe+q30bndYCvncqLeiJW1LLHNYCjn4xO7va2VUYtheZJHuS1
oW6iNNHMMyDWVtNYhRWs8Nx0wO9t9wcVoZDOLqMh0AWrJthWTyvJVCb9otho81oi
fW/ERSjk2VhDFT4xdYtS63mcHo4KtPSv90100gTFWKvlKhzLVlImS1cSm6iIQo7K
ih4L7Kd+Pt/y8ttV8FlIw0eAB+5JBTcn5NR+IGiVY0Su35UI8WDiXE47p87ttQyD
qSsko7nug16GcvzUGexBAgftEV9wryBtTo1JQzXRAIYCAmmnjn4BPANimDWe5rau
jmR7D7Fiwh/2p+FxRQUOgO8lcEXRPxcwglBTia6UMCxBhdtzUDkxMoULVM7hIx5W
WXG3zQHJ5dhky6MLwnqHKR8VkUHwy+y9FGLdPobnkOmW8UjLUd4BZ0OSMG/MmyUc
o62xIcEO/41Hd4Ai1/oFWsBqPfo47V+D4E5R5tAwI/owSdg0NbscfdaT87ZADQOJ
EazQn2RbcU7NSMZ5hyrB8G7tSa8I/7PGYAyTiJOR/S18daRLF5Inm9kPe5FbN//S
Zdrxxz9pH5ao9Ej/eV49bvM71WISh/HZ9xme9r2r9yP2AWgJucKoqxqh+S/clyP4
Ts0ACRbxpTt7rNRyJKJwBPNREpL6iwwKB8H45x60tKhl96GkOJizIkZbaBGwlmW4
mL6rT7i3+chVcFKc4kCVqLKWFE1eqTY8eTyug/qUz7j3nS0ScMai5fU9AQmdkxPb
C0HvcbYVsq9Gy8ohtyU0Th64yUaKFnNie/ie7ysRN/oi3enhXjF3948TTiZgh59W
zd42xzq5OArtwJtZGk7ujg5dq/pBYH9ThdoPn6UHy2jGcbgsiO1OE5IbvIPfuWKn
UT095ynyh9pJ1lF8NiILqfcI8Go2yQfZeQV+TkBXBgpl0hr8UfXqeeKFEfJUXKHG
1z2sIZBX5wVLuj5U+jX7OeyfaonMJszDvzqopqcYpWv8L/HbmgsTrwsiXAMorE3O
qRz9xFqyeI4nykU3mmaNzqJTBAFscqy7pmP6MPFYzl1Nv7pbajTq58sNiFrJfMp9
6GVY5b0lJ+Cql5Go4pvm+zXmoUqX4wjXFb+oYk2zacFrwmQ5TV1kksHa0ntQ66uH
GsBZ5LNI6lR4eXHcylVwOIL+SQXglh5h2ierZg3Sfuq9vv1dPWRcSoDUI/S26tel
sfo7ODwx71WfSoz5ueHT2pPpoVO35xAjzvtCRJr8BsfmjwuXY5xuVZ/VJiFY4s8U
bqUNdLqp32rgTsqO0f61cbo26HfIXTwY/EX/qtb7nrhPNjhMv4FB9T+DJa7qbbtI
1M4IUDpfyXSTfxifKq83w7zeR8BEjyxpnJHDAG+r93P8mHsYFzuzfi53pEwoAxTf
aEfhXJQ52vsvsILok2U/qPBciLC11cs5PP2xb8b/WbPr3eejiK7ZI6JPGzRsFjzT
8+hPPxdz77f4VbRfhyNzsfPdQwsjd761RwsJGibrZzOgnp9UgtpGKF1M/xib+eZ0
qeT7xgD9gSoTAMunm/rzE19k+3acke5kMTxPw3B2wQjSNpokHnOzuooZVlPOaTi+
hJV8Gm78erxDheDnzsq5Jte83vhy0ND5ttNf65f+6oeIg5Z3loRdXahqYlB9DyLo
J31rK6fIjAng9fL7DfV2/6VqKuzrj9A3ImQ/ub6KL762o7GfKa/otdydFp8lIy8U
uUgvDVwTgNS1As1Y6eCnYpQDlgBLXOcIo7ubGDar0JFpDnmlnPK+MsvXbGp0yzI1
nV+SjomjDaUNFKW6Ta3lEEY7KWnwTgGmxQDXUqHaNRCQEJytiioMfbicUxABAqUv
zdf54JteVYTGODo7agkJfPpq1RfzLAxQlmp6grjMITe8sPo+8nQcHTGMgypHdX18
pHiBZC9GyFcSEFJghdBc44pwHJ/5iBUK3SRwf0N8QpRf2YPKEYMBXzDpFdp7j1zx
I/OWVfhPHb1MrMX3OWXU0SHDd4aIuO0hHj+0HCpmKtWiHKHDzMM5sB4n2NYbESLm
IFPxBbYoc/CzU/0H2rtCxf6kBkW8k/AptajZas6K/RRs+/WQm5u+LuJBqY+RexeB
78YzZJDesGvDENeBPVFDEXnq8z5dkbpv84xvv4Bwa5TNR2wL1RlTCL7OYGk2Hz3c
0ihUgl/UbkUl0Zc/0S4AQ/8BVbTWdBZlMcwhOxEuktEEWCZf53uCmg6xYS3H0C5s
+kJDnI4oAZ85WOXJSKE0k1yEUqqMOg/KbzXeepT8PMFvyhMUTUPqL6SLkEhiWwaL
FyFXhGcvOcvtGmuuGVHjC9eJTLRlHUyrtcVZFu6Zfam9XaSprYM5wfOiJ3zAosry
1s3Onl11dfL8bp/MZsmzWa2nM9E/+ebjO1w6APlPJl99Uum2TBS450oQpDvQ1VXc
ctKp/FEKRJY6IIPj2YzJ9Xmm3CdkBJ6bxV6K+MzDIShyrWNa8koQU2WET4Sw5F8y
3wUHzdy39Jc7CYYE89N+XzpzO82dbGrh2BZOsBIMuzLGaTfpy5vnLsedaH95ZmgT
PTuNcuo4zu9HEj+HcC3g650wN/Ah5IewM9+jx/6LV0jtY5d+vgicFjv35q8k0gOX
XcdXSvQPc/moWFpkFLGCGqXNnk67mQtWLG5ltLyy1v1SXux41O+zGUktq9vpUZMp
IGihdCq1dyV3EFknAPKRvXm4RVUlk2VBz2Z+MYzRxHtGhAzUk/Lv65nKGOk6Pj0S
zWklclunQYPSVR9poRl0IH3Kz23IiSXwwcChc87EOPUqGn78L4GkMdy0LgVkpvCz
v6+ADqqNUnXse/p5+5CpV9GIk4xfzQ50jgKRZbfRff3xtS+q3alcICDDMnP+GIA2
r1HCHrVqDsujLijjysjJrwqCSUhhXb960GODXpj4f+tjByD4ZVkENmGzgYYXR4kE
hVf5cafrpLcg+osfea0SuBoRw/u7mOjRXB3GGcfyyWbTVeJ66h5bdsbUf3a6jep1
J+pPnuFbi+LIU2dFn209Y8BIMNYRPCq5QuuaxwfAj0+euQn8K9tDdEk0GiJvz3wJ
YMZkTzzM0VXRYKksVfuLqm+jvRZ5hqtiTXBzE2mE7EqEmMGmISmhwpT2vcgRSz5p
l7IXfkScXb6ApP7Yeb9vXD3nfRqni/uyD/42M3Z/5/bW2pI5JBiJLAL6cGayzc6+
ZmOelFAKkLDuHn9UyUkP+b/F5sNaoYJzdqj8W1dz9AG60VivrrRozD2Ajl/ZXZv9
3uCJAonXbTr4MXN7moUBn+NrGMXnyhh+Aowl7Fz1zxJBM3D/xMIGquSlg849FdhG
gvpAv2gkJOpTsS3dVHj+nHXj6JCoZo+lwdSXxTlqmaBkwyxqXRMxnC2kYJd1YZ+0
B94hQ05BAQxuvVbXNDxKMfpP/DDssS/sEVnniRY8AT/7OAqeMadmph+5Uf5FJ6/y
NAcOmk4nY3jnZXlaJ2ypzP2dOMXGCwOYV6kJ9Fu9U4sIi+MJglMwhgOPWDqO5e8Z
wg3tr4A60J7MguWFxeZvzBCcQGcErv1ACFiLTVn+fIWSivF4o+b+ps9jCESsAk2h
xWWy5X2aO2HQ5GE51eAZwqVGQc87R58OWwpnkQAbIOPIxFeYuIunaTgiD61PsZUx
ZKzQzR2oQjbRjAHRByHhEDywJTRMwv5tvGllJiP7RO5qELlC+2VaSrJqF7kNN8Lf
swHbEcxmSPeCjcwOohlT/eP2o30J6aGQmqRGUg+teh4KSXfTRG0H8+RqWFkFIVuD
cl4DJrn9LOhomVpYHCsGhJmx1a7WG2AfjiW5SAc4giOBK3p1AnMfhkZmROpkM29U
C+Tpl1gi4GiRqGaIV5Cu2jNDcvVbnhl5IYqEkKfwfk9/vzAk91bVHkmWrkSsAiDa
H62jmD9XRTpecI6LUyN5MufGHAlVmsv5vLorBjHMFMRPyvUvM6+kXuQNPd6xKCBC
tgtXJtDDZwe+gRzXxiF8NmvBZkOIRW2K/rDqMReVPvS15KIPw0XblfXmsmMaNXtT
YjeBWSHKBMSlvcwlujv70EQnSUuoJovXqrkyFFuLJ66V453vUETqa52p2aIDbGjy
p+ZryUEEwrC4eRGk+BD/sqhIISO15oaI5aJ+DSEjN8TFc/Okk5l+q3uDos9K8q63
W2v3i2wWYDlPQE+/ePYgzyu7g6mfqfytEE8j3ok2aXxOZ6HStxMjBjoEYevcdjRW
h8sAvBUVk5MRuLbEw9f9Xyec03GGQ2wVOy8oYiR7zYKHDYDqtZBP0lmIWvViBgNl
mtRDi2XhpYNS6gt46hAR0Hy6TKzb9qBCUZeiAESTyz4cgKc3UTm1k0pvjurSORP9
qPjzzLFbHYh7DN9vtrQdjCQ8wivedRRl56IwRCC10kVQjcauLmiVFYxxNm6hAi6M
jqF9t20UjCnKSo1aEzvV3MbJBizz0qBPO756LFN2h1tbQoV3r2+mX0aD3RvqtfIn
4Qjyt/8W2M5EkWamrcRk+09mPZorG4KTAz1LWTFO3Atsi61FsFtbpi0H4cag4OU6
/nHxzSq2GKEt8d3kzYQuNlpMYshkR+rhJYMFr9T0NAg3BCsq4kUlIJpAzB2fSFxV
5gW0+gLys4WKd5n8H3TPvi8GwpfqV2XBBTa5B80LBU/VQscIF6KxHyQQHWCEQZta
yQBCZPoRQy9r4qrsuFDYeajP0ZJ4iDOE/zJHvTRrXA+zx5O7lujfQSe+ocKmWOx8
PS9V8iVkWasEz2oupNo1VPb/b8Lu/aq+2T3jCZXtgLT4k0Aw5LuNLLTWVYu3d6vY
G820bfli/VL810De/rCkkdfLMusUj445bmNKbBx8fw9vju7/sbCmfFCccTDRlKp/
hmVxo9z+I5AVkoNwlRrJZQq0XXVMCBaihkgNT9PSIhOTaP64HP3Uokx6f6cBq19U
qdzxaiLaRKb8hOjAVq6bK6AfVGC1Z7jl/rv7lwFCJ4MfJ52WvN+//24/Zf/81X/j
gRffQEK06s3Sq/2pnEDjL3Fg5oZ+Blo2gQh7ix8UnzthJL0JWUy+dzWJ9Y9XHR3+
n+dk0R+SIPMtxcBeHxA/KVZh1DM2Z+jogYOZtUW3gZL8qcW+0F0ZojrM7GN+VhgA
EY3wBIb+ixhEFddX0UODqVr339B6ixenkdKVAvoM521RACeKNE+VHtEKRnm889pb
xwg7qtKhgJjKcPPi9MtYgQtCPPMco1WeDQlfZN1Hc+90btt6mFqunHhWwv1GyHRj
blUOBAxceVUJjJqmz8EV9XxOc7vRorjJaW3hlqtJZABotG1dreGwYjsZEzYB+Fss
K7huNFW2h/PAdBhAZp6wfNhZVsKrUyOHhk+KDX/8BiANGRtT4MbpdCPqriiFACio
rqQ9wWU2OdXdGz8h1DcnWFdLXFmWbNMydV0UhQsMKoJcevRhAgNo/aBE6FlhXXmW
hjvEV/JidVkIzWPfUw2vwg7k7ihORLGjbc5ZcicnPGo8/rgU0SYxMPQ1V4/PgRCe
dVr0+eU6akwYa18/h16zwGCZ5lAl4OywdqHUakRm0KM3i7uZTXMbY1WLWqmMgNUL
CXN4ZyWOE2ex0FbLtMkH0HfbLgpONkFf7BczwA/957Vrrh/YMccHh3ask2oj5N6l
BI639KPAlJGtXeljbnbKEwlSX8GUl4Q6WAjhW7qrLgii7txpU+qofHzlkc8SSc8d
mGjnUh+nlGOyaNUDo+cRat8WqxduwNaa+PuzBtZi7fX6BzBiBAK53rhUQ3jR/n7r
6GzWox7yzhnzShOLDNKVMupNja710lpO0oiS7dArf2MMx6lrwhrFU9xGRVK44afL
//Kp+QrM2Pkomf4Tt+pbMBdMt9dEczfZQxskxNWzGNAkjZ8ijstWbM9d2aUkKfvH
TR61lQ3iWbCp5r6DpHugT7bUcy6p4Y+Ib+uZmVxx0JWkd0IguKcpXufMsQ5UMilv
HnX+5vRNC+CmwwHNtE/D+ZtADEog778wCQ7fKFtQN1FWZBwIIK2NEVTOy0C9mA1j
RJkTL5u57Y5+PyUb1Vob8z5tMF4eUzKRl8WKDZAo0Kih0mVnXb7gR1oSszp/x0f1
NMvWHf4uOP9lQYbzPPCqKZNwNkGC/BCcFQDHa6QbLqoIgC5S+oZEgk82UdMzfdTp
RmTfUJmCjNsqPxSqH7IXVhsmGMVyHQDlVNgbqfKgTAK5MHcjJHOmmYWw499ql3T/
bVfX6WLfHdGVQoqalLQnoVgVuZUYK/EkHzlHLTIKnvx08YnGm3lt+XvCoAVUXMgt
b9tbc8/tSCqZYKd11/hdC5H2s0KzmoZcA1tmZli7aCgq1bs0FEelXMB7Sxfp5gn5
yklF+bC+jVCZRHOhG6CdOVuzMLQeGORFp3NdOHN5ln3hnJqNC/wsLIXPjiMfCVME
VShTqP0c3/1VU3F5dS+dsMaaKqiIB6KpV0Opqx8UXL73yJxG/p2kbaA93T/yA86i
v9yCDc7DMVIo9Y5JACReS0+HJagYpYWVLDVrv4Cl/qScUvZbpIMFMXrNiIDPlx8f
xTTE3dFiRR2lPyOUTHo9iGx09dFvItnmRYIlhkyEMBIKoNx2dAAPwsA8d2jsCCej
Nrt2a5+0khtJF3o/Zi4ZflR9IYqvidajMY5kzavJWJh7hIGH83cSjrajj/ST6JtV
X3MkVPE0iFjE2DDpN8JgEiyS80j/mGtulAInl7vc43q4hFR00vEWnlcvRy0LUbSI
yUnI1FsFi9Y2Byl+WwPMBgQyjkfb0uJZsAhCH0ma35LCbUREOEX8nPhYWTPGbRjk
rkygJBUDxwC1GHszkTQcEM70zRfcwEwQJ5RB8PgvHxeDxK6eeC9wWgBQEM2OgfDF
SVQOGYYaTTSlNp3a//HWB8IF9fi1n8GwQoQ4qtbD0JTTa86jCg2ppwAVyfiE+Dsx
cnefEZXcoigN3t2x07HtLinFPpKyn0zVSEflrhQEHiFcEVPzprxsDc1R/kxV3q48
NEW4Gp5nbI9Tt5nQ3NW5O4alFv+vc3/dnqQuO8jdge/mBB4zdbc2kM7nl9m56ZaY
IDehTCK5TPugjXucQ6uI+a+bvDJUSfhI4l4jrOWzV3/iOFxnoC9jDlvWk5EGEbU9
oAVmN5dEpoih7LasECDQehkXTZv0ce0+qWFdJczimGOG40YCDNML3L+5tcl4Yh6N
fjR7L4jAhby/de0/Dp0Bm8MFv9VJBXJfwcwWzVD9uHvVO2ZVTXRV/GsOIZCPadxP
kWr6KRs9/i9LBdfPXRsnHAXRQFMNlNbUxTdOCEHJY9rHGO+AsiQkAfb3a7aNh5oO
DZ6VJKa/06mjukKswm9dUBOLBYhpCDIzQViYRh7IxD113LM8o8k849ToI3THPKxs
R4ZOatJtTLae60AoJX5qFqyxdCS6/tTryxw1IuBKVrz//q9iw7ZeFvSL1OLvB0mc
DB9kag1D5j44iwyZP4FF8r+qXiCSClrMs8iHru3ybcKe58/9Wh20HyQUDzVpFW1r
6x03mBns3/kLcirFtAIieipYijGadeAPWO+CxIihrmuXtHwV6EmQw2ckuEJtADpf
mU59I3ivUOdP47FINJLaRgc2Z32/u+XX15Tkyh7ytCAGM0rp6wMKQTNiRutkLICS
8+npt/W0ebtqbmumCzkZbep0GBSdmG+DS0MJlIAvPjRpUOFZZrLQ2rEfkMdv8dRS
Im8pWynIciHlwzf0MIoi9JIkt8zR7wOaMG7j2UQvCCMECl1vhKYR0kF7lYgP7ZU4
imydaKL2bbxIQlu8mICLieUgjdTNyvbgDJAPwmd7PUQPfoC74DzjdbEgNU1ofENT
rbPbRSnoArZdZZEwptWSAv5eF6xeqcYBPelZ+grD9wJjhnrx7+soGl7ugqh4ie+o
scr3CE4jDFRPL1tDNzAi1lfgeTEIzRX1K/ts0Wq3OF5rOpKUPEywv9MJfh8jFost
bNFaZZWrNQmmavlHwYzA7soE1t6wIJbMTky8YxGnPsuStQvMDafuLMCuePSH1d+H
fvA5zSEzdSmvCat/Ia/hCzOMFozBL1lTEoRcK38IbkdkMg8JpVBSynTcLvBmRGs3
HS+K/QLSXm93bV2ZO6rl73iWVnbUYHgCDQ1L3N5C0DyVteKLQQ4WVqppIiYSmI6u
vR6/EiulRbTddMe0Nbw3oB9eaQSCTlKxqoskIFydmNXqT7gdcJWrlXGo+SKrPPZS
q4g28HsA8FF3g0sPRvrPUSaIpjac2HbaFWzJ0xwC9Rfdr1VPPC3zYQ9X/vD7HdNY
D954F2KF7hOOKxzI6NzESs38/J1cLmyEb4h4BJNeeKyqLKRqRD9EmPhhctscCpwh
nqx493RQiq0PHX475wwPBhzW55LstZPsrRBlWTYs/Pfi5py14bpg6q3JYpmJ7FoW
ZqglvpvCIwVolKxXvmTK9GmmDPlxMvcWOWU2RtCMQX0dwHKvvar1ZSf6+rhnrnVb
9S4YLAlUWZIQwWfCizA6j8ouefGeisfOc5DqetLnk1MxJgWOTLlWyAhxgp/KIYXJ
bh9NXSJRPI2CxNeNkrIhsu+YMIuhQJ3QrA3joOiOnX8T7N0X5I8kbgAsxILAAnSm
TKfvdJ8k0o+dIDdgZ93oJz5wXxZul6rXEU3dy//01K3iXew6oh+FomghHEcwIKDN
6hcllAPqJ34aLaz+3QqdOtCa5+7kuLTP0SWGm0WrR5rXf+Ol//yGNb+5pjFdYSZD
n2O7YIb/Pc63xqd8jHZgOfD257Cyfuy0aSQX79aDx1TsRJ6+sHMzJcviI+QsN7gG
AW3Wy9g2WznFdFYLaMloSK1+YeyzJqZgxZfHUGZUemjJIHT+IX+vnUSgoqsfDmBS
DEQToQjNSo4CZXIa58ljoYWuoxoym6fO+lUqLtjMmj6HFG4qLcHDtSQkYh7esxzW
NGVx0dnzZNZBusHYmAMQw0K8gSd30i5bHUWII8DeaJTRt9M5XAVttq+IPN+5f5IL
Eo66Q/0vZ1tfnk2lUpdCygWkpqYXxeZjDdlOl5Abcxmv0sYV8KkVIoSDQGkK1k+h
KSsPxsLjeg6XPj3q8APo1J8Kj7VyojcX3uz6JYFUj14VYgHueTnLrlv6zeZ8fcqe
7j5tL4oohR3WVUKOdpmQODgfICuE7kGetYEijeZVmBWHzQOI5VN7PXbgpkSbTHMU
dDBXv9h6avtkvxH7xccLBqQdLhvqGieV0izDCdPdiPl2Cd3oykP0aGoYXkajJGV9
pPeHo32f9nN2ZP5Hc37wdESM7iLMBOgLxnf74mzk8WXot+ruRr+gF3mbUK3zEuPY
GQovM2ujgMfSZ31m4RAO3VK5hVGkEYXqpZeUWeSVanT0UParMVzIiNcKRyy367f6
3SW/wamxVsajhkjl2yF2ksugNltZ7YIx8Ud7UY7ukoxTjpV5XGZjzyFJqdWS9HD6
iHjFT2GxPF987ZBMMF+d8myzFpJDSI57ZoQs+6PNoHVjD53YgubGxLgVYvzjQclg
yjgM7BaX84fT5YF0tRIRxI3dwQjBuqPTWB5vnsgkkdvldPnOOOYzSgQ5jmNh2uSN
xRmvozRJ+QsLbTtCh/EM1B7SeK2IgL++IoDcoqvguuJwkRyPYCSKubughDsNl41/
omNeJW0cznLcBSNnAqctIo1+64M0xsYTIwDUd73x/PfGnLDj9U4dAJgkCjFOyZ7V
+jldALpkbYuGQ7OimB8oWsqKNQVLvDzN4zsciUnZN57k9R+SwZUYiGCRZj6PEIeE
iNYvaqTtGCGpfAP6xa8xLMmXeHJmz8WeeqRyxPsJ9SRBTA24RCMF0vHKD25zGYf7
M0CREFTkoX8zSMf/LQRGzzTfv8GhpzJJ5bjQnUAzwcZkJJp/C9wI01Kl0Fzd4MM3
XdzR3/4ooPxbD/fKPtpLRrzzMXwrAN4Js2cal4g7FPtvmL7GbG5wR3OuBghbOspk
Nt4unI8dl/EjsWSt14/gQXc2aP4DYzY3lgUSBybjgGJWALftGJ6cDKh2U+FA5dVL
JZkF0BnW2SQVZMAEsNTnDEvflYtOLgNxUxrT+Q93WGxMuITTUFCeREyfZ21wkdbO
wDoEoEtdvgl5SHRrx0DWsAZSjrV+31H8Sw2u2Q6S98N2Gcs9uMByQyAzNrhFC/OS
a58VR0gTlwB1wGTfEAaZnBdxubU4r54fNYU7WPgha0q2UFuCwOaq4AxmsSSC41Ty
3hKUwnLf3KAfTMCBRsEnrm/7hhdxYm6JDEyi29GaQ46UGrxH94KhACgS0kOd/IZG
+Jx6mZokeNizy9gAxtftlAJtHCGbWCigKb/PlfBkI1t6LXveNTlmM7Hq2c2hP9qH
6rm/7On3Q/G2MDYovUtQBYIfi9bxsu4b6RabBIhspeVR/10iMFphJceUbUh0aQ0p
p87R48+KsaYH4/N4AHlSTlSwzqEFQplVhOWSbTHKwOfSJ0yZVi0nF7jZYXj5rUOp
tuGUxY4yLPBzzQLMTydoDYaYUwVZq0bn7DYp2JetOqoz+zE8Aw+TRtu/ZlQlg6f/
xuEpSiwyJENEcmU2hXwXbT8PR2v2ePvb4dZoUVVpngpSgec5c5DsbxowTyL1g8tf
7RpHIXKTlcRQbKBxM9sq9B4W6bYrChUIDMLlwYDo+cphVyIEArDCoLgr+ly4F/1j
SAS5QiFe3Exn8eWdGrp/Cdlf00Tm8j9drU5+fTB7R3L0k5+190QFbsZ0khMhi7FQ
w8SMbudTnln27GsiMneSBBBg2eqTW4xr3G/6RmOp2+59FyanR0pXk73/3MySE8TB
yNeLjoZ/eULWiYrD0WMBjk9rk0bOgDoNUtWaV7+/lpj6cwzV9NxpPoCR92XQ/QyT
Wd8WnpKSTVM2b3lIm+drfSoRjt02zkGY6i1fOTPc0wDEagB5FaCBeHqzvp9PPK9K
6qqiMizL6e2EXHCHprVO44GBD7hAU+RklQqrAK+rZxBksUlliZdFRc6WWzfCfA34
upbVQiGNyaQZRL4ZM+OaBVSNq8T17/swudRbHmZo9EzLfajtybPrYpDtgnPVCSV1
Ufl1aUAQG/oK9NdHGuvcV5cd6WG2UIuv0RJUnmWId4mmf55xfXwwYd1T2/UAZ1w8
YzmMvm+UPjGGXoOkg5HIIq/106ATdeZkqUYT9i8RaLEsWD7TrlzxuvjPhSXyk6QW
lnuqYbQTPdr0JwZRTLvw6hYa6HDil9o1zE4282GBebmljGpT2Jvpd3K3KQQjQ4qh
QxZuNd0XmkzoamTaL9oCA3lSTjLOgjMQ3i+DFshIGCE/No6M75IoAARcCUtS53cw
brfYWUmPtoZN//FTL6tutgH1Lzv13POpAWqG1IxgSMCHjPVKdjSj9XYLipY0SdFb
eU/xfTvym+e+yuxwYUHXYvtGo8ijcGfH+/q7Hh4Idq+PmfhXUO2Q3eHXoI08yJ1G
hprssdp0MksT/rjk2x9QSC3M88R8a18Rh3t1m7X1DmzPoO614RSca0cTvBZTyli2
eWbKV7am0K3t40hCEZIgKBIuQNgz5eECIdFh5m7D250RwJ2TJiOnHBNbZZ5BiLp8
tSzd9MwJmxLhZm5JoXhJ3fQUiY0gbqIYtiAVlDXxi9eTrFMJFe0bXIR/nsYLa243
QaLCrRQaKFFjfuXpIA+qSVaFYkxtDzs3y6niCED33R4lg9PBw3B0K1a/apVbj9UK
P0T0PYSYqbBTFDzckQ+6EjGUP/G2X7/lYgvtdMklhskrxkoh9LQ4eqlP8Zm/u4K4
X1KHwhLNNrrMS4AP/kW9FhOqak0Do+h/MjPdWQ1RivccHfZNm7o6kcY/ZNd/xG6u
aF3YbGDhm2SzBJlf9kM4IGWMzxwXc8XXWq5vZB4w1cy1hSEki4UV1BkXqacVItBy
u/35DNBD6PV1gugwN0veJlwEVmhSUYQGWmExW8JpTUOavDcGM/i2Ron5Yps87CYh
gnnClFPCyoEd2aXQoVrw351qLWsh7weNmFBDT1xf0NuaKaekYhotEyy6vn1w0Io8
3jhhKl417NASC/O4jqbKrZwvooeV7BGQ0FiUwumJvklz5CX19jJlcGsSKch9jEGJ
vJGeB7WDomRhFyc1w5uoKkQwnySw2wHzuKHJE9X8XALgP/eWzcDkMR7RFJJNE9Kg
rlFgEMZBTzfVb5zSEaTALLjh+s2ZNSCjDKXkXIjz4vDeyK6CQlJ3bf3pnX0h7wI2
G4E6u3rIW/FH7puVkXMU+dgqjlg6cIeZOoHcCKJGCj7zkJuCJnna/jLnqJatb6HM
E6PXSDF5Bz3NbqdyZvbc4LwJaOinmuOsH1z7ayLBZCam/qCqA7h2JQR3I9pYqCSU
4KWvpk6O6mTJzuQtKCyFRFsgzDjCktGuURD/bEGY76TItJwep3SVaW310OI5U8Tq
x9fT44dCWPkE8XbL9nNKvbs7RPi16ZDSwXiukjgCJ+6Jb6iSaYETDKCblTHIhVwA
B+Nhaxe3J4yiRt+K2AL+1Ad6ogxe/dhIruVHHoUtBlNc6LxUDBQ5VgaVQaCSUr4v
ob87fU3MdA4zKAyqTVws6BBRh+5TbJ4+UlgjXS+kThR6EnABIhnTDNskU6x39ACw
VhEj5MMEYvMB5eDD1Sc3L7DmdYA11ue8sy3Su1GvYWr1lDHo/VlmVGFHg+ly4cZ0
zXDbqAcCBpXqYYQBnTQUKGqML7l0hrXDJTCGP0YoooFvqepZsgJ/MmLgxguCyRvL
00balWz8y3tCohi5ALYkczBLIrYbJzU7/wOt9f3vAMlLKS4UR+DukhEZTs3qe7Wq
OmLeabqEay+ZlvxJbLPHih25wjEajhxypVSUjBfJ05uE/TpBa7g44JNxE0xMgGqb
yMo7Yh+55ct3AOMz/GNAkJiVnrRp3dtdMlVLGhA+mXvsVBkMVS/lYnJH7nQ2ryM2
5vOvTGQsixujA06+7SQVx+cHaTG/9V1F+VW92GY9uvjIRu0SRisSw9jon/npNs/W
figY9kQd+aspkDvVXKFiNhPFlt4eB1tsvVepqpfiUePiJomax4nnQpIKQsiEZ656
iUG8Zo/UB4OnaQDWMNhx8tcVdmcnbGoP0+7UcJ8IdhWhlep7f1c4dlKGHaRywLPY
/ktTBFMZKT8oTMYYQooUjuiQduDoJAS2QhTt3u+qJE+RR+WHGJyJ9EtvpWteImuf
hMk3wyT2X0Ji9rigAtAgIuDQoycgyQ8Oo5v6V8Ap/SGFQ7tZdYmrXAVJ63H6ddX7
m8ZU7FnI6BqneGStbdqDAhQwI79KJ2cdQJsYrGVjPGQL+Mji5ZgmAnU741V4xSlH
MjbZEtAgxjI1fge+WETdeoRJKQjj9Uus/ZdjwVo3a8zByqs3awY306w6URHJOlu3
T/BcNcJ9+9M6LAE4/9rBAOAfUZm2GxqLKuYB2Rs3p9EWiFYPUvIFlpwNPzj5EjQc
6R1q8o4flviqv4b8TRKl+i101S0hoo0jfxMd5auD08ubZISJPDwX40zOC8fQDcBY
LJ+ub6ciKujFw/UM3qRG+kUkjV+wLS3k2zMGZ11CH+5t7Nk51yH056mCisE55jbA
owWmZP6uYWhFQbpp9E9cZyqPKyhkGg6bKdYK9LB0OokXXPX4slfJHT9J4ZxeilHW
uGmvxrNTjUBzwXbXDrnVti78Br3WjyTg2z6/Ut5RFA2ECwPFsazcmTv3o+kwCKkO
rUun93RPQTj/24Q/wk9swUm/TnPbzGI13lOTdKscm6UNxzI4gel8zGFRYdjTU/h1
Ht2HdYkjoTYnwTQafahrodpIn9URB1yVPHhuL3yM6Yq5t+tVMZnAiRA4ziSukAKZ
/27XeWmVL6zSveW9uEEfFqEdXOZsVyY0HDwiFrVHuAAnQT8tj3RY90S3FJGg8/bA
/aTD4oFa8nQqUwuskox4vgtKqjju7AviGw4pG8iedjANcUYeDkMhO+KSjBlQquX9
ynQk77O0sBrqreYY6sx0rzxa3JFT9LQwaW/nFefQvaak41+lOxpBdnUPSJnACjyX
Vfph3j0kCK1agXVJk+glTFKYb7224JOD6YXvUDMXcBThVJ3NT49K6Z3740eeZlSR
FECQ8qyOoOA/hnZyw1Wf8DiMVbWAv/LM1vv98ErkNc7We8lHr0RGJ0dGodv7Eaf8
VeU0+BcRA2TniHp5QLq/VjNpPyjmtvi0I+i3ZjF4Brb358KM3XmRJ3CskgOkZqD+
x/WwGSjqueWZ3bvXTW/EBu3um5RjeO/Si8kn3nYzAXMyd8kHN2PJ/+K4Fl23I0uI
gUCv5Pke5vDOoCT1thshSOcgVLRZyhTWnoN4O/emflRUnscD7ZwZp4ehnvdSWtsP
4CFXJMN4PF5j10kU85t4p/VxfMj0hRWxHx7f1sH9dT8rPk/4MJvMEiwyT8uIIp9S
1+7LXcVrBhCEgguaB3TIh7t/kuGowNx57gEZmUjweIG8s4Esrd3zrWFJibm/EEIQ
fj5RsXdr+u+3fwSuNULVpqglZ1vC3MxUORjHf7mnWttqFEwhC8rI3RphrRMhtslw
S8bH4wp1Ef326z4PU8UNiweA0lpyE2Z2IYBFNoNozVQae6QKYZIeiv3L51ATkrrY
FuLA1Vk90rhAuuzhqB+jhB4F0fN0C8yaXw1SDjoCKpgFV1m7J5tdebmVk5izpTMY
TwzkNgUotRlv2HmJJD2TxxDyTjoMcZJBtoIW870b4t8gk59dQ2boFJPKj9lFYvmw
QfdVeGTBchW+S6cQCsaalPvsnKRSk5dUXhccgTQAILn3hXD3283HSVm56IwOytkA
FXYDpFDxHaKhsSBPFwbyTdLZtgD7e6QDU1woB4Sb0/YsaszsrLacG/KcjTJLnkJE
ihlohNHA5lv8qig65hdG/5rQNyuHV0RmFm2Kd2XUm5Hl3GUrWXqzKC0sbV1YH3BX
/Q3zGUrj3ahXc7k46dYp6eB9gOxv+xCNTgqXl7P0ORAoVTmUeIpH6m6hFlgok/Gk
2I9nLz9BvUGcEcQiVOvXys9CVs7tc2AR3zGx+n4t3GYgLvgCQQ9MPxxVyytGEMO5
J32eKRS2xnxMs13QCXE3/GV7CiYtxqarDrWNEAXpPIwuyq/9KY4Lw3qJB361EvCz
zjSMkNmRsoEYfFOfuVdP1tg5NPFuhU34wb9M/kS2LFISj3bVCKCljpeuycSVUujG
wRy2JFtphSpaM0sbGtJEY7l/EsB399ZWUwVi1vXTrM4dnWp4+R7Nh/YhpVy21258
vKdFg7JGB9yVBzQ8Ud1JmT7pzqGr12uCiOB1XmQHrBEAhxlSRyyR4Rx6429ESixN
t8vjsL4MMumoKZrLhrkm3L+YoDUrtSklaPnFU3L0zMj5NSL5453aC2GeafvPiV3/
Qhj46tQLS31eYI90E8I/J4w7VDZiQiNe/Z4JtZMLCoCFOEe8yZeVwM/PNaPpeLLR
ReCMuFJ8TWsnrbMakkgl8gIbKiOowANjT8ypTUeqMEo1jWi+jzVa0bCvtxGBFCYv
7rNPgG0qritLjytQ2mYcEy9k/vBPhwGH9y2w0uXbCrJ45WLnomJLPwdc4uR11gVp
jRvWiIrNBUIQcaR9ybZTIC2J8GVtM165oEqt9jai4HsR/Pt6fzR4cyQV2dtyT+Y2
+jm+OnoULDO4pXz/0cQWexhwOlvrP9FsRg7p41c/yRNc73E0sDJuxDvR6mtnoh2A
dvnBOtRZr/+50eRxHUbFFrBb6qhqoNGeNOXaLk2jYQQ7LjmI2N4KXKXCKoLROPkM
xTyBWoHheQ+iAodQ0bpXQIz5hOyzw5cY5rx1OIf5ETBKM4hoDG7VAdA8QiTYdY8Y
Xbmv9BLq1YLdtN8BcSafEmRSWpFoZZlDo7TNOaMLdZFoqmKCNR3UaldeJJpYhlxa
Ao7LCwbF3F83Yb3mwnPwB000ALvQRqMlOaeaiXb+1oRn4eHPcN/ca6VGIp/LDkBg
s6NfFbQbqzYfyiAKJUunC0Rzpp3B3nC9faQdWP2fBMmMcxzfiNAoyhgLn1+NAK93
UV/Ke2gYmWppny5KuOJOb8g+TBCZblwhyy/jXeltZ7T3kKdEzxcLBfLCQ7ma1ius
NxP2wVCmcV9FCGuXoNuuLE2JsCigolyNxBNOA61BEsQZwwm2KUAsKQ5VoOH8SdzC
iu0F/YfMK/m2v9R0drTJMoLfu1zSehz1I7yVi4Lu/kMGpqNHeNofwL7IrFbbc2Ja
RjkkMDqGP4KcYWkLxs9sx3wRf/7O4EAA5MgZmauEPNKmWXcBgrvuP1rGOKpmJ1yY
qEuA/KWpg9TR0S14ZEV8bKLMWhNtnaXztLx0nhpb9LFe38Pxrr8BGnH89leFtEOR
fraLDc3Fg2PiPt+AbLS5M/HePKlnO6RKD628w3b3i9ZIRmvC/o5vAkZffkKaJDCw
B/9Iewny807arOo9WfjOKQmiuzbWM8pEqz3H7C8UnkuSLlXzsA1h9tksjMpkd3kq
M6dy/7TZlpHE/s0G2JlLZgNmLS0/0FSPdeeqX3X46NiMwf3UyIyrYuuLjb/5AmD3
so2IiZZR2DZaWnLOGeSqdMf9okXAY3frwlOGaNJHcAVUVj7mdwoc3CWwWKwOzgIM
nkaKTTfPnXBv9VYyCxga8XQhJvZatI0jcXTrZQclBWgARCqtGHLwWfPgl483Zcdp
wbfvzynyj2RB4ENUylo0sOFuck2ur+sxdSWqg/Sv1UlZS90h+yzSGjrJ0NzJkEvm
VAWxhifAjoMKpeU3ANluce6KhYI3SPPioDqA8QD5XSWvNbe6ycRJRYN9cwwmVAru
FKCHY0opZO0wqVioXew5BHJL7rTmV+wTpkFh0Lu8RWN2Lb3ylQIq9LL2W2qCs0j9
hCw1eXXHe+96z2gUEAOvEN64U468RnrQsClis+8LKfGVbqrxBgcsl6cfVwH85jWp
aulELSdgThPeax5OaOiOlxRvMMn/37InSpxoNyiGsCACrYKfikOF8kUJmmFSl5B5
i58mDmnVr2DfoYJwh8oh+Yhq0EKHshIH/o7Kj64lheiAwRQm+dBOLwD7PeaOj97E
d8yaU9H9eSIwZbCsrRRAg+ZmgWVePQwBs1iLuEx0KDQllPizgpSfCfVMTAt5F+Sn
S+/AEUH8xZ9GdnxRoqzUpCPL4W0485Rfv3IRksEWLwVMzhRr8au+VJ4U8/LCBt/7
C/RAyxIJT7tIqTL4kBy/ywJRnLXkYJydm7q9F01CGHXCw9QLfhgfqtUjfkv9hyMF
fxFZGdYpQnANtMwEdVoYchhgRDVZrj3LunLQNXr8Do38aDhS7lIHxq4qmx23cVYq
rUYz+gwpQlZ1yku2VmX4rFEType70D3O08MzlTbXjsIUFVHglfe3kAld9a/JJA1F
hw0ZkdLnnKQYMI3i6csInNPzZXF3mEkt7kSktbWIqvWLoCDM/JaWys3oLgygs4LG
LrmizcIKKd2epU3FaMMYPDApZiD5UJtnRUjQAAkUAzEW0e4XGtv9Z57C45+zd0ml
SQM2qbe//cAc86PEBOAd4ty8Kd+yhnbvbf3gjIaG8yXynTLf9fZfad9pbhprHNmB
ywL1q6RohL2TWIxck48U5zGZY8OZjC8kP4S4EH5UAGsO4q4yQQ7Cdss40YQBMN91
xE+3b7mcCY7vYJlZs3yaaa1V8Me/jrRNenBf+VTU24fHth9QKmlfGhzcLFSSD90U
OVICtjRaN6Oe9TRBh/VWq6k0F/YFVjb2O8QWvftShDvqND5B+ymbRxnWgkQXYSiJ
bIBVIr+L/6vIQBzrPNBM8NAFk0h/i1XmIeyQjsbq+zzgnklSzQVxQjkUDme6Uipv
v1V66e5UEUxeUT9a3KHg+SdM7RnleUuhcEN/+n9hK2b3mDHquj96gpMomPEjeJjD
WIpDo5t9jDI/kMpDe2a/eM8Kih4aJR+UQ8iQafjwRgy+u/Jbs1sd7VMCecnfE1A2
VY27jasOVYxj/ZM8AIl2hkgkxFQ0pPGIwJRHUb76TKZ5EzRV7hdsltu/c9mROhuc
pzW0LjtKIPjPaYlPLwIRZpVH2tlouy/bQW8jVJM1+nego+zpMHULaW6Lvf6UjSoL
Pvvt1uEaykD1qIsBECJqz69ltzDXbVvP9A8MEzvN5ipJ/UwzthquY1bTAnPQE23G
jdphmakeo77rcUdeegrO85XrMnSpyp6h0UUL/J+G4DvZE1pBJ/7mFGCzz0rDJPCj
PlLphJ9HbB1FjoHlX04FxErK7vMBQ6itVNGos50QWWDbwxBCUkCufxcCjx1Pk78u
55e5sp9qxu5Rk1fA0TnUrWA1+ssvrUOi1s+BddMiuDdzDsh15KODsEvUKUR3Czs9
OvU4EqDKMfw9Ddqs+tpBqkk8UYtmzVmph3zn0nz/5uwtNH+sUIVBZHJUAep0wE4R
6CRYSOOOT2NUJlDy0lRGLyoaqU3mXmyev3R1v5+y7RIM+Mvlqifo+OUu3J1Pnd3A
W50FI9FiQM2HgO+CkVZo24ld/5j+pydxkF6FBu+LoKAGAqZ1QtEEjn2eOZ8NCD89
iXZ/LXQq9zuC1PQ9GssvtHWtMcL5En/hjxD2bY4OjezkMUUTlci9Vwreccd42K3M
QDxOj6iikIjvajc1c7rHtTnY4vo84U1Ma7WgwPWWVzXd6tA9znhsn8yTnohqswn1
3j1RIgvqyCgxG9tokIMRAYTcq8QSTCG0WR3qfJebqxNWe3LpcUdORr9CR/SRTdsr
9iksDbzoWZj1rAiHk62cBYzKhHeK3dnYiYSvUwwRwzs/aig+t6PG1mXQld4yb6ED
ESGG5cemnwySvsccz0s0tkTcM1k/syTMA0TEQmXk10SKl1no63mEcSeKOJIx7Ny5
wtxF5VClLdsJZH36XtwswbssCIKb+33/BRLFKwioHN+L6vAoA2pdxdpbHSp7qImP
vvUOrcQqwFRisvHhL1f4Rrrwt5J7gCb/TIu65bvExqd2QTO5MkC90IY8PkFYDCIx
tNnYVLRGOUZFBh2HWCCBymSWJ0PS8LiExQOyJSMjnR04DvfdEmp45As35FHhAJyH
UOtmjxfBDEZRDvvnm3pHCBKxAM6iBwdFTjhCdu9yJs3OGJkNA9piGPuuy2m7uxUi
8r6oQqVdzeWT+Ap8d79UTKAwmpgWnTpjiZoB/KlPqttl8NRrA4HPvlYe/B8UCiiB
d4MlpS6moFSNAIzDIns/hIqNmIckTYBffK3VDQxK8BSYtB0n7ZNMDOjV2+CfPUH3
Ebuvd3U17fQeEvbYyf/n6S4ZnC/ivPEZZ/SOW69ADw+b4cvGbIXsccWfm8gPbUF7
AM3zTn+i5NG5ml72Hds8Iqonk1IgMqa4G+sz1ogBDuNZlpG1rK1l1HlCiHtJC86+
sKDacCj/Me2zFGCMoaDWUPNJVgPnrxJgLAZ00k2XxasbaJcyaF+BLvfsGwPvZllU
xrNtg4fzKJ1H9U8JB8ttwJrMwnLi1WPd752I/K5Ioh+LJJELbQsA3VE9f/l6oeY4
dCzkUQEIE5cueTO+eLZEYegzZJkGQiFkq90BR1QsCy2C1adHZ2lGDdOxaWga4DaS
HfnMa7ERR51HuXg95HRuzwtnj1uyEW6wTIRMLB0GJsElEJhQ1UBBsEa0df1Absyp
pnkTxVKnr/RTDwMKGLO/Ne+108EY/fV5Tj/CXRwsOgiOf5LvuXk1+mqibzQvn2xz
IUqbonpu9IOM0TNtrBKJeKxuq8jS4vqsMaJzL+A42BOcyrhtDim58J31iBOIU3nr
bwcIsZHMoaC2M0pmNfLgi0n3K/m4gp0wfNmZnbzPN7GSyGVcB0ARQSGugHyitaYz
oIImjULC1nxTAFerbNcqrJTdLwfKiuBdyD87JzWoYs/b8c8EFer5B5IJds896hnm
ST7O0x70ZjTsPlrEZjocmGoFPuXVXhudrF7c73b5VHIjb840jo/w1Qcg76I9TGyi
rKhlYb2w4UvjmhBDqTu604BQg33FGUeyWhj6dmbydeKc76v5aDo6PTr+KQjmQEzs
CkhEAhw1nI8J5KQ5BeCdvLbxQnWLR/gZB4hJRgcOdL+MU2nkxQyiswqw71wmpKG4
V9F9/+VU/ge1aOzxOtpaBPO2vtxE3/D/4bEkbQNh0tGGlC51Uj5PfXksnwar068C
cYLHSIIXcu7O+FhjF/OoozVL/m4z+FolK+WUAHBOpgXxGUpfzibyoxhGe5gXlhEy
qxmUq3Kr/hIRQ7qDEIfdYuXq8VHrDg/S8tGfwIE/hkSZNOVIZS+aoYGAanpOASJB
QkkSSwbNujcrksmNEfBJswaiCy/cj7scWm8ccjqkLL7Uzz6Wasm5EOakTmPx7Hha
Q5aY1rO76Hwpbu+K0srdNZ5ZpInMNywJBUU7QoQZ3We1btKY8UqbhxDo17eW8Uvx
vtdfNMBjLHpKwFnjX6G4364pa2ebIR48Vwnp4OpEpxWgF0Pb7B1h0a0r4sXQycb4
rebu+VVQ+bTBUW6SDlinbhFID0P2GJfaU/Urxk7hdAywW8nlxfaveDweZMshyQaE
WLPwpDC9HZaGkWnEVtrkN3naF91bKQFbrhdXILRDRI4pEw8/c8WNy0Z8FQuodtDP
yFNu4rcenKCPr9TWai8t3yzOjHHUuvK69oDPvfsh7sgiB4wH/rEQLEOzHfiIdyHr
uTgP8kRPtRepHrT5cf9YTtNQBJ4ySgStD3KaTNeddNOevMg54HWEviOOoY+jroZN
XYa99ufNr2BdfqdSvzdiHQ2JEhl4Byyf5MIOvSgQKiO3jylhgeSQe0OtIKsMSeT2
bUhwv4uQQ5jdcZTxHFeQV6W4xK9PDOfPkMqNXJSYrfNogyjVhJnzM6Bjfl+6s+sE
opLYnVik9Gb84DQDNWNazrjna6MrqoMX7f+sA2grvJ0ZPivdFa9Z3jlKg1YebPr6
zSd64oHyBVbszeAmL03XP7i+6O3+K50kL97r+yiFB3tNz0Hoj72hLq5HRBYQPtwz
0Qs1rJz/V45xVpYpL7b7wUd4tVdpt1no0C8QasUpxnVbcnG+YOmTOBwTcYdPfFmn
5n6UaM/DVQAWYmKlxs6njFqpTPUOMnpEB9pcFqRGiqKAaF8ZEwJRyCA44VGSAvgx
2QU0JLVy61sQsnsa3ZppYV+1qMvSVXk/Dbehw5Cn4pFkqbLMTcjpEV26Ln6xaVgg
HK+NhTFOlVXtewvHibr/N7vE/zBdjp15qgt5YyT72Wd7OLm0TbOwO67VD41BZEry
c5G8NEIBo7Q8XQS1vwfIfqNJlbWWQzF77XkyfPFOcOE4w9ash4h3Zh3FquQ4iiw6
9cbKCZK2chPg9LasF2Ao4foF1yuXNd2HFOq9YvnCPbGs6O0N0nWgpAE8Bn4Y8Dp4
KdNBXGSGgfPBWLTckBX0hd5i5yM0nsSt4N51dApbfsyYbDn0LX7XmDB1lamrvE9g
tRtbB8xNe5ZOtZwU0gMuvUtgYsdWHYq89qE54PXOir2Inw/0vIMIxB3BKJFXjrZr
+BYGXRldnU6irQHMyEQVCloHbyngrz26dlkSePJM31514HLqBEYNPZXIxRiXVHAx
DKWppZBhDgQj4p8jrK/RwbpRkXt10pKTbcDQJQVy/8L+BWD4+3EIRKOibQsHCskC
yaJY+Y3mP6KfDjfMpW7kXhph4KE53z9rwcevZ/pr0FkWRWDzmxT40q50LXIEUE0b
R4ZKTkAcH2m8F+EwkKBCuNiePGKrcAoep4H1LGVHfaWMEMZoYFXj77Ko0E+N/vw0
pd2FSCaG6EE5m/LKhdhFSDOmkKInv2Dw9atB1QInEJkhxWbUyQeXt/7KYYkIGxfi
7nJx3qpTAoYt/i1vh49O420Pd73ei2X5EVeGURU21XqSfVM+sbYIYFRdfmSog08W
KCelMB1zkp5AVUmeV+hCPpOAnnqGG5BAIY0VC17ETWF6v5WMP9PgcBWXabmh73KS
Zc8W0ZOCAitxAURtS9Ik6/27NDeAaoKblcSZGI2wmo8RRJDMa32zWDAhoKvpZP6e
y+SB9SusGuqiGLgEqPl6E0d1gIq02JnmnJwsbEd7e7Umdrw/PoUfSXzqhBuhn+ns
L/VrbFWzKkj8H9+2KyXZquk52DHY1oe6BW0w6whSzNRCq1Dypxp7z4ciDCK4E1SZ
ILbQJT+ViXDJ/vtxAq0NVFqwWPu7rTYMMEuK9XaRkoIaxU6wJsx87FVIMJaBR4IX
e8gRKzh1fYZh140YuddpcplpUdJu6sl/n9IYAq6Xks6RHF/hqkua0HE8HTjzXcZy
QmRfWGj1NTdfrWhRBc6yF8RFQ4GYnnFMw68/Cv7eTQhG+GNdhHiBjgVWJVVGA08F
8xb71KGE08LxCEqcBjvOH+A2vs8EmL4fuJGxrugGyq7w9guuC+YS+RITwRnLM8yX
qKy/k3UvZ6S29eOGGukwNixlBs32RciQvAL7YxEzKriA8+EwVzZhj6dh8w+rkWe5
SfVOsaQPr31UCiCBg3/56fPB9dz9WQYy5wW+iU3H3Z3QL9j1Ih1n6Z/B86cDx71A
dGskOJxE12Azi68kVaNX2Ejk3LjOFDiqBY2TmEe2P/CO6x7XW/6x5nOSB+YCyrim
lPabbvJw5EcOhrIO3ftJg2xDL1UvGZTMEkaTOPAiOt+fSq/5JrZHR7ilBazkuh4m
sxkDDjmmeA7NO9Ib7/sME2s4L8K7MwQUvHD71MUjDuia7pRR602KFEvdnZrpP2gi
RzTKbwS+OS4pFIBw/xWzdCMwHHR5dexGFKpORXMwOTTp1+0w7elTXUMl9UblL/zn
R9trPahgMRq/0F2p84grtUNt+DDCmwKiQ6iwpcB3bj0S4xpsAi5MvN+e0HOIcFoD
q9gxtR56+gRE5ZxejFvEQylhv25p4HR6vB9vXAER1jL68iJ56ok3u67en4Y95n5P
BUhWUsbiD/lJeSWHOPKwY2CkKgVi+NZ56BjntPJBQ9oRt8DyDZGT5KYmFO56s7we
kFRzMJEH0FZggGbU/vMk6H+GaOqdMo8Hjqr5ij3pbUUmtRGWa7vUm9lSM22C41Ep
l7/jxN9XETf7aaaQdH2nrYSeGfR1mpXQ+fTCxH0iqV9djLnCkfSZrzNbHadcICXY
puAi7gCwDNEzzAb8Bm4ejuMEIFkLMAMS/TfLhwkOhaMI+NQgKbbtEVp+xOgYFGCH
ETDLLHCXzlN4EcK6uSf+K9VKNA+rJkN5W2MF5pS4I64X+4TCfwBHqN5OpVzrWHEu
qc+GF2WtKb8NPC6PzJDwZ4GCpIyNy0qGyYZ1tbIKHsN4rgbEUMhbh86fArkepFkU
1TSsMSFtM0x9jsTj3R0B8oqyEX5vEamxQ7nEqLnWEephyHu5LN1YFnKR8sAcf4qS
3DQb4bwxYakJjC6zb7vEdipENmT655H/Ve0s+nZqEecqn/E4XkNcDny8C+xiGCrH
9ZtKM8CgjSzUSN5+v5vWuUr4akh64fVdlh1rHuVgi+JIV+rEpav/tws/3kBMUgM2
dkgGPMPcyupmYfPT/BnmjsrSRx/d63UWIgyQqeB23Yz/e37i6k0rWI28wdK8+TeD
OiYlcevwMcG1wrm6+vSfDTUdA6eLoZyrubX875QjwJMeCYb7+m5jJBe5K3L+FvV1
DaVIJIS6MfCEgMSijIrY4LZgXNzS39JlCLbImJ9e+r/7sFEX2fEyNcb1S5BGLCrD
eY3R/Ld6mmbyZXsTm5mqFQkN1pGyDLZ+u9yxmoi7mQ+a8ahT8kR9pZE99kQHklAi
XoFPc842qYe+geyzPXBdEE/29mcyxkryO6lULWk+dgWPpk9oXokp0GwdUMKRaLI9
VUQZRiXEQrSm/qpMeF+wUGsN2eEVXRtYBgDEBVCcKeK8boBVSNx+BZ62lgT9XTGZ
4eY7lVp8I9YCiwnjy++c9ShHwDE+Bh6e1X6ee0ULIh9kt/EHcYlDbmi3Ndq6pN7H
D0GBrnc3drI/bjhCj8NDrZCo3jCmngt5d5KBFXPL0RAs8xEKUeU7BsDQ7gFXZRR5
Giyhy3opO0Fx/JJqZCAemEfk+mvlmZNDPgXj/guS2JWZ6nC1eEaBiajv66eWs+bF
eIkpr4EJDTlcuzpOWSFevdPA2hpgAFACfvwuxur6EnIz3FoRRVNk6oF4gV2nS6E2
E8SVL3amfiUBMlL2xriQp+kguc4Nv9JbY2so6syB5kRXOPxEbxzZRxzIsvSzeTZj
DZ0f+C6sahvmoBf3yvS3dnYVY/Uvl2z1Y9hSzO2/mHR1uKIUW0ugFpe1Apzm9hYe
DMcwWsvlHGQFc2J3HLr6NoeS2gVNjWrBWXFsYO772holWGlDglXo3H9ZAWtUWJu0
qfJ0rU1UQw3R5fdIxKNCkpdFvvkvfnGTshxNov/UQUBRtoHevFZoucHBcr6QPmtA
0mXsWIfMfOkCXCqJEng128myrykCJGovOPbX2pGlEzdkAlXpkc/wdYko4kMD5TqE
aNHswOcpMOdbwYAsWeHCB76cIwxkmTTyTJn+yqXTCRxznSNNTQZ0zUNQMVy9B6c3
MyUtlhQ37oeNujQC6JUsYslAZXwRTaPZI0xh8YqBgRsDJMyJPdyxIul3xXVk15Bw
KAUdf7qXgpQxGolLbFllSrOh44qQtlx1+UxrwHqvNfCXeHqHz3LFL2mI/KQIgWmg
4oE6+oz7jtQNMu7QEoDYix3SrZO+rAppCqZuWvXCcDArgTVHoObXl+eLqCVF4qY8
O1rtIzvzwyjCOVbhuDxnTjmRZa9sWwGyt/QDJz0m8AfBi+r5vHV2E2WX5ysdsay5
lvQTqpRCwn9Sb0SvDmhpxMs8En30OO29H+mPYKe3ZXRhltCYdHRAah8IEyGGNyXb
HDRclZ3/QUxSnbmuhqrQi/AtdQ2oZKXUaWSJQbM+l+FN4zJNn9MydEmqCrDcPIaK
ms9aKG0yvkJks817XDmy1wc0WdD8SDEJLsGjHAdMjXiggPtglrEfi5Qo6CH3E8Xw
nKWMeGifH40JfnfZdqhX4kde5FYN1ToeMYcLkRhHnDc7j67p87F3OInxu1nOfzfZ
f6clVvG1jPd0MXjuSq9edvYYm2Q1UA+tT4V0i7bNKT3oj8lYYSDwL6dZGZLv4Qmh
Z459sEMteM23Z0fp9zibdi1vPjjhizZ0qRhXJW+oEFm+38pV4Om0W581qd6q/bZZ
bc0GXuwpnV87omqaflgBAqSCK1541+lQyg1VcCuvnizWxuNeE8wI8wXl6zySBPLM
ewgfICGnTM2vrTyRXnlqygsZjpP27yan58qewXNFL+Zd5x3aOfpPaZol+dqbZt2j
PtC38aS+qDcl2kpFtiIMv8oQlIy/vRKiKsMm8O+R+AXChWz1FNHqfA/9bOdEyFT3
ZaNk5ycdF4WUXXQahe9hKhlIu5OO8BJiGqDAjvOtMyk+wof/0B0/9TJ7g/mOo87J
p1H5cJsSbi8fX9mA4ICydgMz8rvVletnOrsOB/CFMqiZb2/0YdhyLNlQhQgHXjRk
shXEJCyDMl3z2mHj2QXFCfZpxeMv3rQ2tg8wuTOr6D+wOvqpNAI5rMX+0SrsNnm8
O0wA57JdYgPVyYK/bLQx8zuRkYXOMyb+b7fuR67YIxlylHD4kVP+7gGIyGpdB/IY
8YCTLSpP5lRDTT1kaWCzDqMQIYfA1PRp/00wR1gnwYce/BkflQXYRS9Ho8VdGAXO
aR5q9q8j4ZfYTn5XrMNUA/Y6HBCIp7UNmx6RsRGAjX4PC6AqMOWxAIATlqP9hoT7
+C/xmQtxPmkWKP8LUK/FcIjxJqo7ivsxaVqnpRzZfLG+R0i9K2ZslFDXhFCsCgo8
2JsYVhGi8OGta9AYxdS84JDVLon4bLvj1v2SixZV+S9nxF8LKa5EZ5YhZrhgNrFi
gJsnIL6lGRCVisrAmFNLeXyUr/h0kw6vlpV/9tIWpsNUf8HLYEyDNeINaFXxNURc
ouvw9OgeBDi8zJRKZ89DDbN8jcOoumk9S1KBcuUpKTFXyRQLnvu57yjC+ZBhxekc
tr0x/LUfKoo5SihMDIndG1KmdjzsRgS4c/9lNMNAkUZtUXnqRCTnuq4sD1rXb5I0
Ex28E9ww0IuVkndkvskbXDOBmMgcYO5bSwUnU/c5jrLneEzeO86fkG82SA1kzm3E
bRarvdembP1MmL6i+KoLIkNki4KY6g3ZXGBYUSeImMb3Yw/H7vMS7xuGWUPqN9gI
wAaL08jkabq5VqiQGfJcGonQRpkqJzlEcbNjSHX16VxPXpYsOb1tPyXlnDVDtSPJ
znw/OixrwOOoPs/wQUmRDQU8LMAVq58ao0HK77knO7nG1b3JC6UQC7Y/zeDEy7yl
zjRq3jEF6dPJjYpIVcfMBoygoRf9oevvKkXhNcx0IS/0ypJ04wTjCFpDecKp+Mfa
qbR3mccxt9J7nkOlTZIkd9osuZn0bTiXJUx+D29yhXxpyDl1G+f7dr1Ed3+YsQzD
T/5Dhu6KePHpu816N+h8pw9O1ai6JA6Cycyf+EKHWvflNn5rSN/i9+Ge4NI/CeZO
tE56W0r5wOocc0zs9DLCBIPphw7AlJrwp/5wh7cMHJHw66lDQAi8r1jOWSkzDzW1
/94sPIBFOs4NrtHhrFGla1nKRRGzFLfKb9N9eAH6dTLjBabF65PoTA1k9c8N/gXo
yz/A/Hos3x+neCFcS3umgwbrURH4aF48ppdZVCkRlFbGtpNtsd4l66HtRJRGJp4a
hjz/obvu1OFpTeVWlJ7eciNQyKlxGvJA4Gce+3qFEnjhPHGp7HeGv7kDFKsYaHFV
DQlzYVbtDJdqwe1k5sTfxtzJ2zmdVbJGD9OomKturXL4Vo5lg7+4hpThRo/Jqv7K
TO90Fj0El0R1acDfnYeKKDXKI5fmLCFRteOZigk9QearH2oK2cXcsgebf1531dxZ
LKsjoijKEKcDl2600r3QsYZmIoqJNsUfN/SRX8WBj12+nogwa7Oh9Yb2dJ1bNyR9
g3Al5YT9VKVny2NP5nTctC9w+vLSZ4ZrSmzNcsP4N/Y3x7ee6xHJPvjn19qd26kR
JwOsq6zAkp5iDFT3/qScJWQX2KqFYT6unvIoqWLMbLPOVtVYTY/3MZS240RhGE/q
gtWwmVoR4D5MW4AHGOP6ZRQ//k1KhYZ15fHFx2pbMnqnnuaqn1jzQzNNN8jZ+GlS
RkX0COF2zWdjzRg4YixtMSzXHAP3yVlupKcjrkGqR1642TtbCu/PNdSgn/S4mQco
7GqPDqvL2TkqBaLUgQ+mqyE4Gk7xlxZawJLl9Tjv4uCthKY0GnU2tvFKL1vhZ5TC
lNVB6z8xYDS9/teimjOshwyFRIOUER/vamEq74mTCkGXeLSGuS3EfmMnIwnp70Y1
G/wpwpKTngl/9hjp8eMp2hBYLHI6QmCbTf3dCzacSTS+ccmqc/JGMcsJ5YWvBP3u
rCSIALrxog2lFL1ohfhgWtGijlDiNAJtDgr+xbjsswDjnou5dpPz0UmE6ul26abO
E8v1dbiMrL3WsCOmi/a5KbyWDAIumQ79Xm85E75ybLLWp3MtIibqkIewJMVdqtu0
ZQqKFXK/AdxqwKOykILj1xYQU64+lYrxI5hIsHHjJC5NwdIDldPmtOgB9hPPH6do
A+1jkpXB/v2+6H38gMOwpA8reX5YDMQbkua2xrXDMjnQbTmIQg36JsBzcehzSsL3
n2K0UZirVSNcGABGUxtehflYVXK9emKNwOo4oHCVvGdf4i7xnRELyk+qdYbxHkoE
5RsFl1a7adQG+FH6MQtyxb+o5ngkw4gGe8ynJu8/p/A5DBYo/rJhU/s+A3NowLw3
hFpsDo1mLzSa7sUucTRA42iyzlQ2iXtYXrljtWN9utPvl9Eq8Sk0RvCB7sIJym8R
FA5626eiJXoj1J2fe3YtLVdJF0Z01pnCEoEs6MszNpd1ghA6F8IBHhLLDCblgX3H
18VL+Xmb+cyyFVyBiDn6NlbZv2MRtxpsz/id4uI7Bu5YImwYDgRBoz3pQ1XYoOOY
dB9r7ukxP+7iLOBXuksvyM5wJveGFIx45htGTloD2Amj2PlxpdMRtmvc3QiUfeFO
Xpzg4bJV5RezI9b703GitsGjH5mcxV6Fw2SjqDQ0PS7MZBmxOBsC+CSo+wpYwVim
IeFWDl1jz8IgwErM4xeswiUnCvk57qkyvlhI+ge6Vtbz4cJkuDDDjHBMyiYGFix+
Kabk7iCoFcbKdK80AH0ZG9BhLHVsTgDsIUeQlo8jDPhQKCq101pIw2tmbAhEHcwI
mj16qe4e0Hyep7to2JDjaK7seQCEGqXOmH/Bi3xAWGulM8ugMDTETRO95VTadkiL
+qc5mHfKLlwvy02+UAh3AIkjqOZzi2JQzFhXHStzBY71YXcc89XU7ytUF31NcDcm
Z++V/AEqodbA3tkpKUHlROED+18XLeQyVIEloK05OoiOdS7gAGAmAK1/VPI9QoKE
HDJ0A+k76rhogp6ePf4x6rpu/dOUrWZyEJzmEGHWNqbRgLItaIRbn1LNYZ2eJdSm
aGOtRvbFIOnG4e6bE8ew4Bn6Ri7uSmE0JtoPABjpd8uoeKi/CKhvuY/xR/STBDzL
vj+2goJcUzja2jwc1sPdRj7OPfRcEwCE+HM7Ky/4PXfsfZ8b1pzdkFag+sZ8xdEg
xu9IZdkuzwZ+GkhaZXzPFv9JSk4rzmF5qS1XXxyDbDQoqPm+s/nWCubr0kML5MGa
rUHVMYsY7Dcmn4A4ecKMkoAcpBDdTggMayLsgF/Cxn0Sfaz8X066eaO2/1W+HRzZ
hp6ay0guk9yP9cDOO6NJ1JqqaOE8xa/Q7b1W4GwwO7wIFDikRfNhEaHPphLwDd/q
ZpYmLPL8BGlTaQ9n31xLKDjD+RzmWFPQUMEMparvMfAArL3roXK/EIyiz2I78vk/
26s7+z/AAE6iWLqlA0n//WWk1vXb3g/YfpYW5DpvlRXXCP2xFohTTW4NOLI6PfAF
hH9Cj3tQ8b/uW5ye5Ae3QaNkUfr7XM0AFwG44pUGdlXh0eiKz8nPHlleG8Fqi34S
6AxY9Tyr8VTdJ8KOXCRUBUNcRO1uIVXbXoghE1oRDYhDZq5SI5DcIbYUG+ST4Ai6
4lM1Oc048/5cHPL9OBmW/wtQbzOGoEouKCVi8UlKJY+4LeNtUlrNFjpcJXsZUQgC
LBz588brNT7YeGLcyMbP6aympxhKQGrsqRHksJMOdqCpQ2i/J+NE8IYAm7TNRkIS
I9tbj17Qzb4EeiC2FW9grrpb45xomHokUb9M7UwYFeWyPgqG6hfgAILQBHPcHLJX
cRkR6YGh7cjxo39Gq/w91W53Gj/qm0nMuPOu3QGBPZGgAtLExiNWZVx/4EvtTnSE
dVCpCV+wo0BcAx9SJtLnr6LM3UPh3/CdrxEw0l6wwOLHmnL6qJ0Z05e20mATno1o
O/koL56xulN07FsOfElFrvB4m32g2Zupgb1si+1XfU3THBqPqnKzbIz8WOehtwZ9
siv3/d+hgp/hpcLKLaENaa9MCpHfE/TEzG7OVTE9PXPi80ldTAv3Y4rFGtYCnL0T
4aEKfuOg5BxGaAJyvo0uqzLMJY7aBNH5byZh5onPODgEgITuSzKEaqrnVt5HDXM2
ZnwmMUE0kCis1ZjYPmgjbA6T0nrj3mj7U639bJIXXJP0HNfTMr2gtbsS7P7XNEHp
MbphY+IoYfoBdh7QAdzgIBC9sGirPtGrsGtYfdqaYkdxpCDCMF/D5R6PjJdsdSOg
WhkWzwfqo6LI4lnrzpGqXA9pNePALWlAsbJggjtdDzLUNVb3/kyt+fQCGPshcU1N
SQiu7OlQLlyEB+UNVmpSr3O78jZ4ZYGbPB7l4Mcnk1SqgFjUwHA8UnDVZrdDT37e
Rgspazmt+p1VtBWS1SssEzsveHKPY3oWMwgV9aKLKe8IDfef9C8OwIwtXWVtG/fw
9hsiqnqAb1x8Xcj/hOR47XkbcA/YKZ4CrH9MZ9nwC1Rm81dZtW+vcwzBikjvKB+7
DvfQN4NOYozjlF1oIqs1XogW4DnHT14Y+zpNGCo8pkd4kH4mShjNM7LlmzkK6fFz
dI+7TRKPwJOrT/9TUVFFuX0q8qZ2MFCDd4GV/394Av1H9OMsZGJ8Wskmrsyo2m05
bqdlPSP5YazCEaUbeu9/rbnYeBbOEvUMu5/+ZtqPkecudWSzF8lZeZnIAzqoYdtC
zgAfaTnJ+F4UhymmHVJNGu3rckY9H48ZSn9LIbQjdVPuDNuwiUj7oCM61P+BbZBr
VI3chpQCviYfEqVj0n1wARN6HiV5mjgfFyIkCgzPq+oFXjif2AODEWd14qrshz41
5Toz/eOR3UvUrlex4zs5U6/o4ERnXoUk5B5di7WPMyFnESTLaog5CbPjiSBB733f
t3pnb7bihJTR6OWDx1l7AcN9KpmCIv3yJ5n7C8t0bJlEzlbBurr1E5pQ6iePPqZB
SrvV/Vve3afnXyLRih3ucmYYAd7U7m1td9mQ8NSd+xOEDSmuzibOHYl1bmTIwrW6
F/m1G8h8rYbSr6tO96DtEn05kH0gCZzHi4lGegmPLj5wtSwaEIBnP6FTGkCR8ucz
3bCyui1isVkKpKxBy+/dwg//ZJhI5fvGyE1xa2ExbE8HkhuxQ8ZiPSps5ya4Tmz3
RJ2x6F2M6vb9UT6sul4xvaO4ATHAn/1g2jcB6PsmmpriZKnlZft/qJwOqxBXzH1U
b7T5A4vgtVswsgYo6jtVMN/2eCm0em+OorSi/69bT05rs9cS6K0J+PR1ggwn09N/
oOzKlP4//WxMFoZ1Yu9xl6Xsw5w1XEeKXHFbKt32XFex/snqehKCk8UEziQCKzZt
WgZE/WW4mwwEnCwxEdA0GnXDxi6iGcyT57NTazwKjg2Ue+utojQRajfNwFfUhKVn
TVZeMNALOz0sPyH9kG4oHH+C3wTf7WvVfHisZwUMnWUHAxK1Ql68iepHJOUqqowl
qGtsxo3WxWqEFLMUJPknmlwHWkci/yb9htMRSVyemC0I+h9TOd06T0Bqg7nySziH
IKLyWQQ9W5mHTn1KSVTll6YYBSEHxarKhCyF7kswmc3UlsTcitPrEMh53Kj9giyx
NHHuJWivNapmSKt8sUmIXj+w0ge19+oaGZKw/nitIFAByMUsbs8G3Dq33jZkbd/X
vhsjZFgTCSZeWLqjx5h+raWavMe/KuzgaTzshSoy5IWOuZGv5w0TQhJtD0UXktzv
R8XKbxxR8gNde3scvqzKCYA4VnvXcl6kiQV0J1xYoxCqUfThOISd1MDlIYpZfoMD
jnb5xNkVPBvayqIUVbnL2K9sxwh5nnviIlvb5Lh43dOM4gbi2JDyJTQ1lB1C887n
dLvd4wr/PMEVClfjoIC1dthMSB8iRg/Lbb/55caIUr2eP9BlyJIagzcf0nqffEkr
aoELLh5rrAAONC4ieKofDgyl8hjRwJqqZw2y/bcXKukjP0fGBqSmPcxkhC4Nh8/f
fxEIiExL0PrtNSseWQFvs4rjlt7y/waqOLFSuge8ufR1bxd53TAwvsIkeQk51Fp3
+pKDmBT5kdx5tac7ABnYWJhESLTXfAB5VE+zhrRyNe6YI/puucGshBEzV6Q5b3mi
zDQk76/A7hO/X1XzxwklRuc9gBAEU2G+jZ8MAbuL08sw4F9kWKs5EQpg38J585YU
t16epntDX2FRJtaAggS7wF9cz4p6TwYzu94U6GOkOa5IhacLIkOMti4Ov8riaOL6
DNqn4gpJ10AYPvkycDMfENrsexZX+3gY9RK3xZucIBUc4aHBu9wY23LX4yiv6gJy
vfr0nnnTYXSm9newExA82oCsRqlK9HsgUamzrE4GU5ZtLyjEfGk/3gwU3KRlyVdL
Y0rD2bU0VkewC+prVgsVPBCqjs0x39k1TvYtfpkJz2bMd/C8gkXGdprsfwFVQMgZ
ADPlHDJNqMEo7VTHuykDUDTQQrBEWQeE+cl6E7ZZtWsxrqS6okgJ8KzB0wJQMGdZ
SgX+3yVUboxDO3qkeoVYUEjF60OZnO9smfSPUIfy+RNovsS7LxRv6EvfuzjswTlz
R9OI9hnFfmLDdMDMkzAkp4JSC5xUVWBacCnSwLBbavHsvjWkzN4S7alvFKg2IThe
AgR/raYiMicfyFjOr0n87UXBS9eMELm72ltK6htdbYG49yYjaHCMeKH8rFy7TTck
PTP5jFeyNUIZ/iKQi3NG+8SW51x0+R5AIBkFHn1Q6Xk1eOpXcOeDqdRUDnzEw9qS
55IOBbLZ4AP2KWYbJeoepd4DDT3YrAvQmYocINDOpc+FJHp33xk0RBE7bYqtI7yY
BPc9c6NTv0x8MsIjEGShIcMDW0VfxRq0+nileVZyn5o4tqTJkbmHsAXugdXzgnlO
8wM2GzhD51rXVM56+xQB8cvGyug0GeEu3RFrPnQSprItkuk9n8cuL83Vp8LeRwTs
RxgWo+L2BS/H5HxNIY/geo+WrtlqVNyKLJ5TvTHgBNmWWs2XN4ihgi8pKt7ccpe/
Y+kFa0IMfIVZ3CEdykv+4QXQ/bPLe4auGiXTZHgZCqwECTv8sF3Od+h6emg3IQGF
uznw4oXLj7sV5uVf9Wi5Jd941ODHGD4eJafnv8JahxfKeF2sz13ZycRlWqAwzTud
6YXAhynqg5X91Bmpq2Mh0JXR62PuBM3WijGUa9Yyn/HcQyxHCeqJt9ZwOdYOvzIf
OCKsYx4K5ya/NMGrAlDDjmHAGLVTh0KiBeDTk0dSwza1Py9dzIBm4xa3YyWcp2OC
fiGA95B6kUmVHxViWGFnbZdnWIJ6BMEUPdKbFstPUEbwFMgmvcV34Pph9/Lqi76n
dJRboi7bwry/KSz3NaoU1zUV1L9veg1rdkn8JjEwdZX8OSkmhvXH+LICREVy9V1i
DLvPlVTz3tgz/+jr6c2KPGYXn4sF6rnuB+EKQNMGrUoDLDa4MAgOGv8HXWjxYPuj
gklZlb0Wl5wjANVQtz0Icf2KBSbCFLDOi9YQkwqT3VpnOcf+SdO/T9Da/VyslXRI
7MS3EpA3BqfV8DM0hA3mM4/erL+mOj9J73HLhTQKRRNa4cYkJuhFMP+BokJM5W/j
/mjUYfc6QMe3cS7TMUoqDMQT5Y2DdR3gXKxhlrAs6r4GRrsGVoh5ciiO5b4bVUKn
wWurUTx/v7WawO+cAN/GR0Q1sTaNfhCjE3GmV7DU/IG0J2G3eznHBJOddQe7Wi3t
DdhvCqfZ6s3amrYsXjPWGjVR9IXD8ROKpsTPKsWgtBjQP+KpM6Krwio7geURI7k4
aX6868zOIkNLpfttSplg7OoLxL6abir4uYLRb2MJ3tBjw5OFvNZZfa0FbRbp0/DL
VDItRLnbHwyNApHBQpqmCSEh6S1OOfXzY5xGRsvF/CD03Hin5Gpjl4416kAe/SME
PtjChU5qdo7a9y7kZlDC1xDaKs4cTFERgeQMnfa/IdlkFNl2CpTG+eojXnFLLhxx
/yl8k2jvobq3Itup/Qa168vyVKtGAyvH3fqaCz+gCnsMDro6tTXEY7lt+uJNTMUQ
N1TSBwnyt1jGmpJCcjzM1AmikzjnO+AEMsAZK4g0s7Hd2/zJF3WCXJSwsHNFGow1
zAKC/wVXWXmIbDdlk74a9nGF0A/z2eP+4iiCj4bfVqLnTtEf8uXJPe2QCNYq3hRV
leH47fGNtD6jHkSB5XQru9vbo1973QUVAKZS5bo/LYmJyoMxRh/UANYX3K71FOqh
SXuV2WAM1A9KYa4h69ukT2XbzL9CUuddPIawYL9350dHVNKxyx5OYX8DqZunTaiX
WyRT7PnL3bNDSsVZ2qE6JcHB7VDDLo+kMigP42xTVqqT6/4Bw19cEEbwzvIPHMKw
/mNqdq7S60AxKhiI1RXLtQapGUfpZv6i75FKO8W9TuvNjPMrEeGdhWn0pH9WfZZN
lFNVFsOFMD1uRSL1xmMgvCP29m9XriS+ebBCMW4q5JxBAKYHs+vP+vLVniJrsj08
l+jJm/voq27YCWf9UQrSp3IoeV3CppfCE6WfK5Czjre1HPulvH01epaQXILJ2LW0
LRa0inu83svxUtPoA+Oa8QewXc5m4Aq5FgxudJGuJwwVqa7AbAG6MAcpu19IUBNX
OHn8zaooFoID6X/Yo2d8tyqqgXdmdrlRcrHVIh2OatSdOcYNO+fvhMSjRTc4Ser+
Ja/uV9StomCRvAQcVl+Bbq1yu8ekhlLLVm61StAp/zv/6/4gMaJxSGjpDqkvhaa5
j60piMML6Lw2v1cRXvN98NcZWeDyfUBxZK4El8BYblXAuiRxGZgwbWXqjLxYl7Wd
fBJnvAu+0zGUuM3ZNDGBKQ/uArkxRwK0yHRu5mlDpyDBRoRyAB1zV99e7AQWRGNe
+eNQ1hTOdFvbJNs/vlOONTh9KRXOCO8U4pJAmwHA9GWI+MvfL9QRJqAZveeVw+2c
TVdWYr5t37gXm+E17aUqCSgZCwfLcLEz6mkw8rhMc9qtQHGJEc3KXWqsOFEjB63M
PmfvsYAyYJQV2CtpIWbQQCUzWCSO5tRBJIX8LhBGw9kJeQw/kpkZazw13Pe96Jpt
BvjnJ1wshFWNoPhUZPUV6c6O4cj4hE0wTcYdDdXYZyFoOMzCq5vMRLQtiT93IXk/
BtKtDnTY3Y0xh5gIH48CnQekfgHFMngfDC3uPNeqGWn8nd732vCjIhbFZbzrnL2q
dfKG21f/Orn1fjMiS2mVgbRk/l1tNSJodjFcNWGfBqRl/16Rz2r7PAXB3bCwAJcf
BDd6fy4ovJ7RDZEa+hzSgxkpGewkaGhyaeeNAPzfxPOzWss3FDdrRRlhwavsAxAD
EnfpxBQ/veGAQsIDqas+4LD2PyfwiaO0U0nQxl1BrjbRmY2gtxWgqRn0JNk2V63a
voyaquQL+FouarjIzAeOFw3lWk808Ia2wKj0e3pBN78fiP5OhXZoMnSoXF6zE0Ww
+IDKQz0ufIlioDH8AXVMJUrxKeiUIfJ4p6SzpwiJbWUD4ZmL2eUQNVf86HxzVZcZ
tZsWyN5DlrXLzF1RvCErDgflIwJjicXllnWzXDXgaTYkiyrft6ajaoL1ZZYt0f37
o4uEW6eqsIp+UCEpTXaZAKCn9vXfHqB8yjrv3SWO/CGsGLdHv7Snf6oJ4j1gv88S
1iFvmsAtbraDe7BDq18c0xRQ+uYyXCeVWhj5Vd5bX21w++5nYNPF7JF4/qm009HX
p+14jcj1Cu6eSWNBH3mNCTHz7z1NUQbxK/9QR20oQ1KcDrsjbzRPT4zkm9n+TJSg
VsGJ69AAtCDqnK2d1caRAADubqvUHM0sL14Pq9ZN0KEL7DfclXL8+h9RIgP0eGnO
JyFgsnJ11OrftZ6XbZ5Xf2KpsNywou84XwU28+Nw2t9yjQBq93DkBJZSL7u0TNv/
bTHZILVPFblHoCNRC6y8butAPoeXKxsbGZpZNF9P048NSDk1oN/WN90OBhGNMbmC
YVtZ9bVueH6Zt0R9iQ23YFzradSdVSRC/Eo+8KD8xjVy8gW0p6Gkoe3cg2TCJmeW
bcI1I3vL0VW2znMIqKjW9laakbI2p2utFfXpxw37jmp9FX9BofTGoB9beuVJHTs3
Sj0Y2mUdy7UB1iTfRyi9MTC1uHwdnd3hzjjDT+wVBbX7t1xtJ+E1vN4XR6bivGG6
dvwdnaji/LhFs5HvKMl1/ZG7n6peN9iz4nCQzXAxN03uAGzrU52mCySpwdB5uAbd
gEZI1F2e7pFw3m66L/llaG630AvhcSthY5HXMHrA0R2x3tqwcGjKhHM6NC1cSOkg
15qFBZsF9dRx5T1QX3QHOLtyuiBsq2Up+Ilp6vrUkIbGKIcizb3YaejHABZI+UKF
HlXL9k4qY1/Fhl6Tv+JTnsXnH38wRHlKVwT9gGFl+DJRDRxIF47IG9T3kr8GH4WP
pqIakXo+/jjmaIaW/Q0dRAgFhSQUhuot9mY66mqgvezrZK0ATECRzwOtN7JdgG/O
BQ/toWhUKnmGMsvynJRneo962xlvxdlzYygKjRa0O91P1vvzEKrnKkaTP9qMXB5r
KAjPHi8xabQFUfJYWA5cUlmWDrd6EmPG146t3z74VScLHPaiwH78SJLRJNAvH31D
w7eunfVVwCoKaheXTdz1xGMzhXDRHLPcvI7Kq+2Rxq/TzpdaeXRd8CeAMsoy8dI4
lnvHgrfHQqLovXZjM5uL1lXuEz+x/uXihFqChxAtPF9VYOlXJipteRaSiwycDhi0
cYuXCnag/ONXmF0u4EwhatAuzlqn44MgIHPnh5a7oC+avAE9Gig6bXE8vl+NduXK
9NzBOrRDMyykN16DYI/LzADoJ2DzqdheDTX4EHljs5OtQ1bvstbJIgjOthzgRJ4Q
tISdcCsv0McfNZHHvSHdgN5zlavPcaX1HrVWi3aVnUJZ+jCwhVd2QWAK3OcwR9YM
pv1I05IVTmqPjtVE0PY7LGDNa9oUyru0EmdmJmExEq0TxJDpP4OLIFgXnenehnbR
tEJR3NMwE6jcqDbvxi7XO4yzTKSz6LjlRfZ0F1zoNDPqMPyLKs0sTLvTZ6ULAyZ7
72LLzN3G4wkSRPr2QKzC1t5l3uXt5ueP4h5ScrNNTGGBdKns37FzEFJFdXZon0kD
JUprmKVLNvUa6LaX6KbZ27J04hF3DiFZrjuGmuXHuiJiyhGy6WDgqAXUM+Aac9nm
LVrLwHMUn2R/ZKtFhfQvBq0IqsXvjjyMLDIlzFjKC1kr4NXdbyU2RWo1vrw7zltH
`pragma protect end_protected
