// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:41 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rrMngXCTxePgc5QsEGDLdPSfdY6eJ744OAeJ7O+e1CYizlHTiSslxX1vKhKNRRB3
U7SqC91br5Iv0zqHMQoMqYXWGOFgrGfRrFrLRV+VDWzpwCTGvHtPqzMIw5FJvfBX
BciWE4AEKVlWlHHcui9wroUWYbs4FltUZHxWSwZ3XJE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5600)
5hiatwSanB3TIwXPQ8QPn941Olsj3Us7CbeQoTDC4SxIiOUaEJWfuj00n6T5tCV1
FD+DOF/0tTFGt52a9QSMgnIvuoHF7j1i1reWfi27RqE9DQUj7U1Fao0ebKwCdVIN
iWgBxeuztD59m1JX+6I3iBHTgp2FeclX5H/9tw9XWHFxrZlpgtElwCeRTJiumfSE
WEK6b7C1WOSXeISoSDmqoIIc3BsVPx9UOW9QNef+zv1PL057EKH7cWRY4f8wEdTr
+9a5VL8oxX7z0GmtJiumLQHyrOWTg/ftHtWCWel9w0IrwvXsb5+EzPdvRAyBPEQv
vBGSykbmta2jVwtsa9H/upfZFiJZU1hICiExDwG1ez5TLkfBn26WNqNUYzIOOBCc
P8Tk4GXPnXVon4QI4PIMaBAa5XXDtNqtEuIZRd8sKdxMbwsEYRyeWIMLva5nRYJg
brozAPXefS4CqsmN7RQc65Q13kyTqqRwXSkUuytB4bU/NW+3f4xUelLIZ2pytqdC
drnHPs6I4qSQ7DlZFWM4phNTEIFhh41sdLB47rdFXPexbjbJf9CTIvxylB/3nEgn
99cJCeU51CzJ6r3iTRcN/kxLsI6HAWuyaxacgRM/S71yOrlpLRI12c0WWfs/WRUy
m4ccfnwlukTBHaPKvopRHk3o0pqPK6ew6n49mgt5tTNgbRCZhCiFjs1/djwuVqmm
dMGMclZ48xRdhxc7aS+MZTeaC8LxuIOXtjP/LkQs/OJncJ9EOrok8D+ydQ1yvPHg
lcbiqzo19L+PPv7EFDMtqL/IM/fprOX5fu6CKKk2vDrDd+He5zlch7l4t/mdFpXC
FqSJREHqcp0d//jjKUQv/niVSsPSR8hMWSzWnla30bq8Ud6PgPSObP0N4lZDG0eI
Oy7DMF5HI+MSc7BtxtAqYFxRLQxdSrZHcASKKqMFtnpFtkbTt1awrxR23wyF3/Zh
AN/IfdhM6gfclOHVRo8PdRIYuBwkELGkd3zhOQiQ6ourqNOpI+PUGaC3DhFqZQkA
L1bF8fUVfXiQxVtet2op5fzAYMms3WsGOCMVRVvaJ883sinJQKPJSUxn/Jy+Dj+V
ctEmeSWpwd8Punkbz1vkva3+YvzKZW8LoBM1RI64CzY0yuYiYlVpbG/F0jO0F0p0
FKUTSakSN90ubstt+SV7JNOWxdJKUq1gHsEqcCyiIQxSKDn9T+4WDZzaZ0ys0nKN
ni+gJdkTRIJPDlhCJ25y2OgpYvw+rNXk9QgcjYunkQ1yKddrfgZcFnoIngMZM2mJ
a0dzCXphyB0Ix8jH275MjMUtUCeYDaKcXepnof+/cRjhCCWH9bgO8vzYvtjGe6d9
fw+8gFMVz+AfW1FiO4VQ4CVgOtCION6yj1GuX287DnvCZwBc4IwLH0Kg1ZaBBoNR
7Os1WHrE6+7Y8vKwPUTmdL73OGrI1Zy4uOpQ5GZeuycyFFTHwlU7ZVnMrD9ep4Ft
jm78aS0qNQmxotjXeKH8e9TqFHY+HhabqC+Y9tyfHZX/Q4jtqj1v8boLtSz5wHSQ
dxnwyZYlgHU+RlJ0ZDXpru6XwYg8Jz8UY2hxmQu4Y89SQzZ3iomBzPoK4000QP3I
nWETcRc+Kc4kOP0X+aK+IzWB2IPyzPZK9PKBVZhtzFJly5LPrBjR+BePS4/SjSDh
djwRE0lZHm1U7fZaOcNKs46kaTmGL8xyXD0++D1x8S5XOeLbtnR820HQ94lHG3f6
Ctka+sfjkcZe70it0YTwZ1AfWPE6LUlc73HPKqfNImek0YFK7YWbeknBVZttkN/R
n+TqvYa76HTYifrvQmWHNpa1G872K7AaYXcNjrdCyQacAV3aBeyKusL5QYHTzNrU
AIAhtdZ5LMSrmk2sgp8GTBbF8BLCUUFQ2NdcnG4Yh1AIC/YjDBgnfDDzaF1+HaJl
JhQevVeX0csnO7Q2Uzw+8i6tQBMTePsD3NsrcyLrGGQRSd6xfi4ZGFa14HEbC13q
LPP7hXMj5ZE5zIePLd+C9/83P75aoiv6s/pG7LuZnc6c4MOK4u4NeF6WY4k3OiGr
i7aDWkNsL89T8nD2twoGJFKvhhCZaLUnJX2CE5owfKzBQMPZqxF39zgj3ariZiGE
nMsZr6Th9HRTXSq5FPtfeT+lN35kO2vXt+YuGGDceBjGsXwJUhScbBQy8A8uCAZv
3CgOqHmesrNQ7kvyExKrrkpuh2f0/9IXOcC56zh1rzYI7KtDeZ3cl0q/z8b+RaHf
p9HgbqbJCLinLT5DkHPM9nVFeE+1yGaxXwrrGuhoLUye3zHj9PSrShIzLB++AnfF
3IZ3vrcTzFqRAkFITFZXH8lJX9rP+8qRlc8fI36fsHUVU3a0liuL94Wg1msdx45W
0AJJVogkWoW0eN+NSLghSdPEtsyOXzBAbmMw5d8sPKW9b9ZkXI3tjZwKm9Wpi7KJ
WE89MUXbSSK7hoGGDVL0hav9YQAKeo/aAf/BqsiYWvumcZKI1p7XUO492eksDO4r
v/YbvewAOgStohypDgRXsvcdzd9KQTlKC4msun6qm8az7D7Ygsb8xDYVFT87Rkyh
bnbWjMtuTrQ61Ni+QjPFaCneUGmv4/bOxLsutZ8A6ctNpI4SPtJyK/YXIltYa6D+
Y0369h4aI5QrXjsqd0whvvVq7HgWezB285uz8KPwtrd9VnhxKoBbvyqPUdRTDaV1
PlVgcOqYsPtBrGSHT+xijyrBOcLHEONp0lSXsHsYDujwaQqKNKX0FXy5b9QbGtUz
Sqt6G4e+I3XbZmBgImcDTRtj0f5L5TEpi0irFiBl9zinqI86FXSrvi1VWdPlzLAF
7ovU6L9qQYr1LTLRZgG0H9M/mWBtjoRo89dLK8nDm1jHevTKfbWnJJPcu2xbsjbO
GJzxoYmB2Wy/vHGyIoQvkF/4aHUvi3oY8vnem3slFA1IvAmkAbNcWQ/F6VIbfrr9
0DPj2i6yPMikzDnUtMC3oedLKTnCyRL6by7FbX9kjPNV4IEGhx6XrD0LO22Fe3KT
gkIxQN7FIrO6w7QVs7WsI5C1DRHh+9QSy1H9kMYDmmJ7+xIat8yCJV52ci0HmdVh
MBxIFm3o6iavE5zmHgEIznatOjkDW0pnGRMTgdZt8CjgGaJyA3QLPj2lXjDB24aN
yUnJyxUC9iBkJOqLyalFVGsz5MQtiKHVuumJQ7z+XnZWLdXgCwMxOVnPsQse7N+d
Efn/G9CXf28L/YcVXHlaH43dHPhyB6SziABfdoHE37rSxoUrSQYzU5M4VjgsvM4t
lHSQI+tQp2Gc5Df2p0RHapB4igVUr55LwV2UHOiJnrLaRdVYw3wiYllsbMN/kTHb
JUpAo0nnONQBQb9eqJgJouR34UcIEsSGKMT59avMKjKeBPBwuVH4FWfvj0Xe0ig3
nVJ7EtVNEQnOmNonS6gr0OcW/ZUZNOAXjWoNG1SIZ/W6HJ0hzLNksqcOvWx/loIg
TPFWGZ8dALEYdMXCUbNWgw9zfXAk3h0t574GafOg00+CWuj8W2WrUJ8Kll6QXW9/
V2tE843BQiloS31EOQbtGX3GyEfblxiizAckeRw0GwQ9sBnjIA50XpahgKhBYuBK
XC5gYUuzoyy/P36wP3OVeq1zwW2UVKr9927kVWrNcYAIi7XpSfska237Qn8r8ppo
fN7S7NC1fd33uUvSwVEPur1Wdh0j/9EOJh22Qrt+i8LhJh8gUUzvxU6tgSppczqd
MGGV1JLai1KM+9eygi1oS4Y/vVzFnVNf0JEoyqlc5oFxg8ShAr3dtVReuY+nKAck
ybK7/T98uy3gYZLeAPecIix9q1APJIqY8iroJcJLKum5pLZZ2atnfA1g1bKqvtki
/Y2ZOd5DYMoKrtxrjVxjmOoXckid/bqmJ4MRXAtiDEAsZuYeQ5ZNRPPxXDRIcty9
lgkcrHDhSo6EwjNh80UOyFeF6VOtI4ZvzmYYYdBP5g10m4g4tREGO7ZGIMJqX0bV
BZNhDu57pe9X2ODv6VkDdes6YD3oNjo7+Hs942pJzM5EqLxyDAh5s6K76wnZNuaO
jFTQtG6vBznpN98ZnSFM6Dy+BqT8pWpU1WAwkBTeyc6eOoDatQRA9msEsVv7bF2U
7BtyjjRsBKZLMfALRry9S9l59iaWL6UsUOkXATn0GBcN9ytUaDf4Sfr+tG9r3RV9
4unAUNUWoLI3rzgoFbWBSCA4+ZyArMphknyPcN0aYj+Rve4gZVoaZsXWvQdzuolr
hgAsEcfN8ANvOBsMMZB+DwDJnGLgyUZmOW1Qtftmbke+YOELX90CvdkcfVpm3LAG
jcFQb1dVFRoJWjfxyy6WwCGoybaM01QEoNLZ3sz1hJ3gUVvUtd5qGrZ4oDpGh08E
ieCz9ExC5ouJ2T0Ct9BKbz/IvgREBm4+2Op0LBnB96GBjl6D2MPRD1F1IOnC5cfL
1U26LvbX4UmhMyqsr64nL9OEdS9LDkRJ5rZndwwrMcJAhy7F4oP4oXyb08gMjH1y
gj7GCfOCntMotscmSMhS6UPdlIYEgESK0RLlGeHIkbrAEaq8wEaQNtE53z014fc0
MtlhwIo/oxiXiT4AvvU70+RhG69lQ12d/76HMl8TL+FXLm40N/ndqJibLpEhPGRD
ikS7ODbgV1y5RFXYEO4vLilF+O+QB+AdTN2asMQapnXb0sKNr0sqHePJfDrj5nhu
Rp/TSccggbu4X56TjreFMk8mjULKZ76GVCpAYff+YaEJNJDCyfZstGdC0Z4BPerz
5laTIFwo3HpB7Pt8ElzZ5GHXiWvp0OuNzSLjCx3X05PBegmh7wEJs+a8B6uRkFtM
flgFN7iiY+f4no+9gbAxAk9oS2Y8ealql1JXrBZms8DEfM+cx6Kfz3BqeGKlJkMG
MdV7ZxOGU2Ip1E7dFN8MwI5iRsCTS3NuUe5oRLVhR6BxfJca9pCY1KPpNvuyYL9b
vBEOKKr/Vt6veMKqeKAfxc5XONyKYu58Ua4oIgFDT0Zg4cZhO8ZNFGkANbG9DJkx
C153zRMImioGGIBu3fYk7Ug0GkwnPk8qu6t6Ob6EkpssRh/8jEPNb1WS04gp5H5G
lD5hEhTaL8tiCkG2AvdZTsP5I/qktXNlyqJyhSsz5p1uht14woWJLvDQix9yPH8i
DBiYBtHQEDbFA6wBW8FLfEC3UGu2Jkl1pjzYnYmaUkEbUKrMk1EGEJ1IN7L0OTqo
3uDT9tfNoo4wFIjC9Yey16EivTUowhA8wemcPNGfh96hkiEXu0POFWN9o2JVtNmY
YWdJu+5MW9AeTih03QXSVvg8n9IOwL4w0PgpK/nqY+rbJFQo/QQ8v9fzcviCgGrp
WmSwLyLs9YRyJl0XSL6hFG/KeFvcS9E3zSDao7LSKe5s1F9QF/MdPlYq41/afzYK
ieZmBIlBPLs/AISMEeIwm8P8OVxcQZEml9O7U23+FpNagDPMp5uGLKha5Q56+u+e
A793MnNuEvbU79jRQYlDE/UM1zZd5KIMR8Or3jefDDQGBS4dBthadvaTuGBToo7T
Nbj6Z1HcbirjP2b03tCVwS+SMG76EWKsOJ8oI2NNUuGwT/H+bkrjDWVuy4mBgBAM
mXlSYw/StwpIIRRt1Jh8AMfy3yYcOr20RKjOg3p4FvMT0RjVZYODj/+hRyGvfrMY
SUx1zlPrOOQgJG2FFYYBmC1UwN8DDlYEj2SyRvmYIVJQqwJ4rzU2T1d1dHmsJp2T
IfPI/K7qMxudWGb+Sagwgb47ijQ4M+XouvX1eYyD5MuRCJQYQ1v+iBMsoU7x4d/X
owGGj05YgQ+LpF9mh1TNW4lFK230PnDdylzhOdcauEEfTgc8DgQ+HgKTmOhXwy7V
l1qnbWi7DIiNH/xMuebaNj9KlWe/hegoSxRm0pPeO4yQvN7AxHIbdTKpNqbKpqDe
6HVcmWAEyH0onDW8Vwsqwec4OtzoTSFAIAyY7fJQyBG1f4yNUGJVsa645FdwBnNq
nt6vXFzstchQtLsTvwSwpBbggVJjp+7Oi3q0twm37rIiltxyo9ujsnjmDFWVRcTa
5+afEY/TB5eHjQdkhbrif1nqqqdLtCBdaHXEIbQDdNlMv7mhVPyP4VSzaJtJAL1I
GDoLvpKT3W+5iRD2XO7dFkWeqZg/MIKq6wwZwQqmI8B8UFd4M/bBl7yuBfYpZkBK
2o3NOSmMz6aMqDmthkI4qC2q57SCbgZmiQn0mtc/PZWF2ukszzE2Zitz5EltuyUh
3gYaBBZIAbNeRa6Q883iI89wjJ/LbdKRSmWb4Vlv73DXnw+M6f3beG635gTpBB/6
B8PbiEGW+m+V8O8VNF6GQn3ugBNKcrKsTrf9xwaxxkKavRYdU8knxFhfUA2Evgml
/WYQqqwnpdMPNxSltT3Roy7rwJ1v9VUulUtQ02QO2B7V/y06IFwGvg9g2KDL/zQv
4ojanK6F7R9GqmrQr9osk95eJOXaSIoa44PUsd8U5vzUAG5+PH2u6Haa0J4biAMg
AEM8BKDjsMoRZaVsqDn19dNA76JkNGPUwgEAO1a5SEZYk3JlPKQFOtFWY67JNz/4
PeX5uuBrWH0XDdrVCZ+PTonTFYVIa9jIirV/AJvmKu2Zjt++wsRbsACJaS6GLnVs
WDENHOobhiPwEpQgDvELLDKK8afL3IPHkl2uDNm+Dv1Cfv2R3Miikl3YvgOeDie3
ApZTPabKWebf3azme8T1ehirzf8+cARaJgUxRBXYe/aqwVEeb+P45t9/+0Yzmpnl
cZGCfAaTi3R7M/epjF6utJ+2G9yrxfXOCRO9BCpuRfwAxrDZuLVfr5M4kAj2aTcO
KI5VB5wF5xPKPKtO9fLg1Sf0f8I973oUiaksRwGbeB4uAUcpe+K6Kd/XzuI6OVic
Dt+/oxoRtT56ZyJ6e6iRgj4bTwqQ6t0iyVtu719AqUEQrF7ZEwKw1MwUao7y6Sp6
WkZPJSqW51uE+X8L5vL2rYJusilwzSt4mwSkwUvKVeaivBcwg/Yqx/yl4aiQtDx9
h4hwyS3x1AfzL1MSnim6rzoV0g4u2NGcqkVKRl2O0G+yHyc1UCDHChoPymJL/AtE
nqXJins82b8wPqb4h485syg93LK2mayo++aqACKXSfdGLKBFFa6YyW4xp9/I0Tp+
o+U8dIQNzsk4wo9EYIB3Dvg7k+4Drxi8/L4oVymwDHew+eIaBYUkykz9XYnF29Oo
xjU/C9XGp54HWCEnRttP0abb/MOcb9VPjQ3vkYchGczZJDJRc5/zt3GVp1itd08N
B9I/VYtRA4USAEnInHawDkXrEnjO57iKkn3MBxQMJYI+NSjy+M+CO5HdLaKXAL6S
pXIb21IBW7H85vJINefeJP7PSycGCLfa1PtcVGeV5OY0H1AJMT6mU+F7h7PqeyPj
OcwSOHjuTPPmWTbwIOYcGNj9iY+joq58dKNLKGBqKFovM8Q0/qwUN+WORpe7IyxI
XzRyC5YodscwQWqfgzlp2H0yhqgqyMh3RPnWglKJkBY=
`pragma protect end_protected
