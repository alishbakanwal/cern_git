// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:36 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
prW1+1QC0TcWn5V4uh4ehn+0959fcOtGnk5P9+xSQ9noNsl6Cfuuzwxix9foWoM+
1zmJWg6gdcIU/oWEZp0LUcYmLbH0nmUAzzvPtPmPwmIGwdhiFuiAXVDLnk5/zRdC
D4Zohx5s/o2iUM/P1yypiTYLCUvsOW5qX2JBn2amZ7s=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7232)
7BKfsnd76l/HdZ4dzkJUz1ZAFMGKRf9zKQt2a5CmcQr5mSsJCtlyOGOgjOJau6YN
zhr50YkWyyRGQ8tyCEzXczOaCZEnK7OF3WLxCtSkFIZJLcWw/tqBM59vT6ugNDrk
lv4HNXEtWr3wP9koi8MC4FgAq57Ss6Gg3UYBbCaLSt6bWdQPA+ltpNXdIvrkhJnz
fj66H4IJOGuStuD6SCEXLMAHYEOehghazzqOaA/E5R15Jg488D2vHA2FA0g2GVmz
1ySWgfdrBY644q434t5YhDp94IpaChcEDnkd07nzm5ThdBg17/uZXNtncwNPVGyk
1SEiDiCXBSVBpcCMWLDWyS4R8atm/aF2dt28oBhiX1N4QoK9opGQhpYzZdgpXH6Z
sp0hoSYxIq4K/w7+QxQdoBb73yniqukwp+OyRWbaa03B0LnBTNln6z3yqphEODiy
gl2D6gZGX5ghOUKaa/vz1kSXIwr07WqejbhAQD/5QBRg8RE76N5HH7tCL5UIQugz
q9JFU6J8H582k1n0c350K5m61zv3VPVYw6DldIJKUPJ+Mx4nwZeT2CqQzV+oLKf7
JWpXSiP468b8hEyRyCF+OpgQJ85lYvMZYpbnMIDS9cVsL9shCmK3Lio4VT+l9tC5
Zm3AOlGQgua0X9zMTxnfKBTdsTRsRlQwoOtwb0UA5S8eii4y2KfCzVLVKXk/qMVp
WadPOwUd/9H86c/GqnknT2+v64/ROX++IWJT45ZZvWXlV7Ezh2hUjDurmfHyq7L2
NFNHjcnE7jk7jcRR9OmnXKIzc39cLu+HH8m4F2uFlL8EgGaamA4U+nCWOsiRT8w2
/Ds003U8Y/R+c7n+Hkl2CWzkUDLkzu6yyJvGNsrAIIMOkntJ1eS510VbOOZ196Fl
zgy+KxuR1XkPkcrFaM5limFiEDsHX/7cd48N9Kx+o3SVBKJpGq5pcsKNfQqADrsr
p5gfNRIZDP4zQHijddA3Mj5+blhSw6x3wQw6jnYlkUzeTtPFZJVmmtnVmh0BBCSj
gfH1I2BpNgtTiA5UhSv+Ca5nEnZ0tckD1g46sTiu+UPjvMbHNPAEFBdztPWNTQux
v5c02RQEzjNp7mlem5+UUtRjj+zco1LL7uUFWq1V+yheaWTn6/xEjF2xbQhwG2Eu
a9HzF55XwqOyI1wAKhBPanJIT/pDHl2JweoJOfzlpgYtSxTPrUezFxyUr9SRxd7t
f6b/jKPbX8nYOVLyA0n7YRz66K4cnCY+PXrU4WJonwqCU5Ak2Q+bzIwB+nCSWyJo
8BEDFyoUfN0wrRBUJ/EqvkQk3C2HBP3CBp20cTiD8uW6ndkga9Yy54rLAJC/f/jQ
5QySMKZhc/xr4iYmJHM0RD4Wuns2oidHGl5s/tfZWepyfFdSnvufYaKm/xlY3nzz
Nq7U8q02imYA8YhJCAPQ4T1xd+YPcITkRzzCItXqVgSRIjVeTfXqWRAE27Zmf9uC
/JmR99um1sz3VQNSCF2Y/Xsxzzl8tsRpOWIgrny27VR1lmgGpbsHvFmlMzw/J+mM
WSU3XRUNyY0ErQWml+0hhh1fBemYgdvOgu0IMqGO6qvHklmhMecNe1P4fBUMsWoL
RTwvVeL5vcZeeAQR/DhDr2+dkT8Fbc6ef0iy+7SrDuMTVlcBroUj4WhrMvmy+91F
dMqDngapgWm+cDjh242l/l7vyP24DI8DbU/+I0pjFRdPKhMimjWnNEXlpdcedAn+
QC9UUceSHhoxRijfxzxVnKPA8PsEFNOBC5cSIuXKfXin7fy8C3jCSj1QMtLlSugf
1n2TYpC3Oj6rSvCIFoH7WJbYxwZGYGiUeq4wlK4XUEeGu3itRFk0noeySZpugf6O
mDSyEr9bfXcuqVFzF7lUATHnqhNTU7hInZe0Z+HBUygu9mfLzjPXnz/LTNsLu94D
rD7uUycKqNaIS11j1PmckshMNpYkG+MvNvUR0cyj2SdnZoR+pZgedeZPiTexu6Af
cjVDSp44dm1e+6hJmQXMcn4vkgmvfHsomWOxXHlML8mqPbCzsMY46wT3K382ZUGN
wW56ooo0on6X7THZXOjtyDl8L3020W4OnnpM5EBGyVZ0XZcgApx6/8Y7JzEuCJm3
5WEQf18cbND1XxR8yILKEhvcPik2ynssxFG5JvS3yVpfMmGR63e3D4Ls9Pbr7P5/
ZIlg4lnwDVw2+gSONT+HK2r3IUqtRUW5X6jlwD7sIEGIdFMLonNhdjW6DRT7k0Vg
sCz/2fuVIeO5ucbdTfLsxdDPF4VYaUrgy5vaC3BYM+pbFPJ2/ZU6v656wV9+OrRW
ykhyV0+DvIrFApI6ijvDuJwRJ4ig0nbUpRMZnU52R9K2Vz0CeSXDh/N2RAMsEkl4
0wAG0wQg5imXxpJCp/jHoAqOziccTo+31DIFyRzjhYsQnP7unzmfv6N0tBJUFkhP
4N5KN9LH+nf+J4KH6ZdVY4nuIwxO2xiVGeOgqh9i4UbOGlcK+j2F23p2arG3l3vt
rho8fDxFeXKuqeXtj4tUDgNWrvySxyhKl/S5lexoYVMRgYfuI/pMKD0ZVhKdJI0n
6zbKNR9cAAZ54iQfW4nW5PDpiDi1AkekBcqqkP382oJuN677w6azSkmpvBxgvTFi
8mqFBUtE7x5Ac2ew+rlooVdxu/p4sNvU/v1V/s/260OlYUbro1heZYEnrwMj2NFa
ogZAnx0nzPLYyWij3EDLPifggz8mxb0bX3wDuOXl2Dbt3nxgtO1fE44So0kFGvTX
HKRAM4V/lUVhi64vKbpfekwsSqsQqfFJ131Dc9qeppj8IHzHgOu4zupTc5Mr96l0
bVDIht0HJHIl0KBgfhssvxhfzhtXtcvn7EGhTmFYC7eW5JbVa/mPhBA2SDYPvNZS
iVm46E57kH0Z5jYmHkGTwUsH7AUbm1wLaun8gyiLGL1I8Hu2aGWDtQZClF6URAkm
Lzngdxm5CWtljBo4mpGOksOGAd/6EQYPz9/vJqvmvuPqxpd6NUo7ItgSgnF27eKx
L1pZH9ymYi2+H9YM64niwIOuICoOqn1C7Rqdu3kLUxDs+Qo4uB+TgnYd2L+74IUg
Hj1QcOS3ZJ46ehx/4et2eK87zVte8FQ+97ZK5u3o/1RQdDpqjbJyMAci9xR1RpAF
bfz7hlgCmOICmt3CNgKB82o9z2QGS75x2zrBsX+5GaSKPxGgpzzMGfWrIir74ZLD
hq/vxFPZE/fzzR46lBU3s7KeJYQJcGv1WslrqDEIdOog5QQJmMaVruMvFkuJgPGg
lmJB5FWxVLYwfLQNk4F+1dHQolOA3SRjEVr+8b1GFV2l01kV6vfkKviGfFOcQumL
rhb/ohKApJbRfc+WVqby8uNIK5SnHGEEeg99+4w6xCBFk0qy1KEyd+5VZGg2Bp1a
jGzjQ4FUoBpo15qPL5nCVCBsONevQjSmOqA/4jJFaCkHZUD4hyazMd482NegD8z2
jceXEg9s2F1xfdzZ3/9L2rFUJmK5O27uq9x4RJMgIVLwZUEeC1m+D+9+XO3PXe2L
LyBsy0xagrJI0/+x/P/RLp31ta4oLLrUt10MaxjMrg/c75qxU+3bxFsCOFwfI/eg
Qi2mpIPza7Q/NJpo+BM+cEAZUAPdmU+iSuU6RyEHQ9qHHpnLVGJXcqiBbshW3/nj
DaSmnmNsc91rpHIRKKnfkpmRuWuUzEZFXm6SeTivgYyCHkzziqCLyHdQLw8pt2fT
SiKqAASr2VcsccrTM1DBC1taOCoPwHZRHJ//fWWrJjMPkMHr+Bq/S07ummxstKTW
gvvw/KJdmng2xwhf84oBQe3s6myWWRJ/grO4q9QHqroSi7QY9XwsFKrHRv9Qp7jK
qCMkhsiNl/wGIByuWi56QiW8MbUcnFR67SuRqBYvIPucXVD9DhKNZm2Sz9vMkcp3
BOYmByp5gWp2vQfuUwwGu94Jzia4xrU328FOcAuXG4/dtlq23scBmoyWJSMmMPx+
x8kQOJPBBOL70DdqEwQtL61RQa5z0OkuKoTnfd3VpHk55DWT/75dzFBm6LmfNKI5
qFufbARTHlEnDDsprcjVNAZ2POjz4dWSykfFaf9raSIaflSbxuDD2Fr5NVubiWIr
B8aK1AP5BeB4Bnc0nNDQbvxvbQnIHwvTTTwzCXRFUE3li3yKS7Ze/cMRjP1BNZc+
fFm1iP4DWbJ9v19a0fUM3lYcYwByAAyOmKUuUnhYs9LUPP9P3U9lhjMBv979bCNH
PYO8YyoYm/MTM4DYQi9QHf4XEI4mL/nWYLsDMQueRX0oSRKI+VmoBpVk0lsWxdE8
EkAQuCEfO757TUxx59S+gRHWVUmXc0VbmyaqjjfYjRHUiT4vsh0Tj0zAkX3EttHX
962noeoRd2Pp9xrDfUW1jewli12Ib0sB0ZzlF+1WDQg+B3zOqSUSZrT0jxLAyB7Y
u20ev91J+XwtXY00prPRYsvBjw2TQ1K4cICYNhYBTkEyhWELgbkUjRfCx2KUHeWz
DT/gLHzCtfD+HzgkYJ4kktCCHr1BXtRaivF0vaaV2M09OD7L+3LRlmRR3LTjOP7e
lSwEHwf9XEhw4up5Qw7n0EzH9UYOKwe9TORJ6SdWg/Q9zlEU0ZtFsMhpsbYD0Nwr
AVsLmFREmD76Jvb6prDibNg3qi4Tm37kKixEPb7JqaCnWTTLePtzp9N78HDbNK9X
VtgNwGdbOFndo9g+bHx8Bgtnrffp+VtDlaL7FiVu7SvHKYor8fHHLxBUf7hIwbL2
1VwVRjr+4eM105/BE35vktAe+ZPx8qOXhk/wlrZLj+o6M9ACJvAK47AfD1QAzmtm
PeGxHYxKGD+8oh3f8nf1QbRtzHujYn3kgbBmrb0C+7sWeexALqfaVk2NDfuq1/s3
4UtdTOfoPSJHuULlYKAtSJuom8QNLGs3e+e/2OxsW6iLjPhtjXY4iBvsXERQeo3S
fYnKxp6txwdJMFMOcCyjgmZFJus1n49RQJy3xp2kkkKfTj8Fxg3slIOIYLPgKx1f
fqA+cNVJV4yKwtdWLuri5QTJemrwdqC/p3vYQgOOapw3D+hBwkZoFndG7E8VCQtN
E2X+EPjSl1Sq1vjc/9JslrKG4DbH8g5gn8KKRfHfmS/gi5RC5738mUip7P/LRJEw
H0/LWhKgR1+pfrSrwfNRgROBnnOanKC4yR9aiNBlEtvsYuTOK4TeyL/j/aup5EhA
mXnLc8XiBmnz6LDvEuUAKmbd6ApXhWTq7PnOt4lRJoPDNWY4eKr3ggewEb0Fu+9i
t7lDGZ1x4/4A0rcplQIZevEX3JK09AwzEc/F7VGo7fsHJhRrT9fuJoFoDuLv2fC6
YpFP26jaJeRHgvvw8UDYRI2eMoNWo6r4YgOTzPq4RQCXCHYEn+P81EMP08qWOeVF
qtDzuklNLDsvuf1pnWd2amSQ9joyciFJKZcCnIv7Nu3BQYDCDIG2SU7ofPIz6T2q
bVLsL7TH1YT6nj5g5lnJe6mXG8+oWprV3Bx7f7kblKQl0FeHhT+oxQm6p8ny4IJe
udlKDkfLfUkWDs9yGO6APyD9UK35CJqIxZYGSheAqAcasnHofDp5e/63Vg4glZLZ
VJ3J6Y8bf/SDPWI65nJsRv9ZnrCGJcDlLTmMD81q6JJGB4fs6Pu0GIv/pxWjr2b8
AdQ0foHA3b8NvJDV/wniuP0TeYNeWP7pTVaVwX75isCiqSS+E0tECYtl0nJiTIO9
DJR1D6SYbyu8goIzzCGjVEK3pDLUEJYHSWxViXn6k66CW/ZuB/m518dNsPL33D5z
ifg0YQ7HPgUx2VEHaCSJgWen5fsEmW+6z0tFlXkY8kW2+/Q2JCvy9NZ68uDmo7q7
Hl7P3F1MD9eWD5Zfi/Da9Yk4Y1X/KEYdymKC+W30zWT/++h56quDSJvzyeeJQ+vG
FewIfLagOgCLtVcIXKN+BJ8UuXgEFKqXvQpBxsR2QWtIylH8mks7sBoYJUAqz/qh
M4WDvoc/Y010EdnrXQf9an4+AvSZMo60Z/LP1me7BjUr/Dk/MsjLTTgOdkf7wSYR
vELi/kb3PhLZvj8KXvFgYsVxaWNc7j8J6100sHZwwrp4Z3zP6lt7o+fp4XW7PfIq
IxUfjVl7xNpF04jdPXNPYcD5F8iMgcmVqJkiXilYY8aHR+6pa8YhX0g8gXgA2/eS
mxC1kPLeTciMfbiEoLhQealaOFpKfKie69iuxFlFnHgO3OMgX1tjRU7cJELjFDQD
wGfIB5cX0rXmRVaIrdzZNy2nEgG2o/ufNIe6pY54EzQaVWgsmITzFwOHhKIjzbpY
UGZwRbkmJAD8ZmB4FI+1OH47cL1ocnZalGgAqgdq57M1lXawo6SkweShouDvBo6V
KT8l0FSOBVFOt29+0ZJ9gMiZp1CgCV4OPvn0nY4VnREO5Ja2RucbKIwUaOuEp/gD
YtNnFEzWM3RhGmjE6/RCBI7e4te3W77W/bcEUFveLB/euw+TKmmqp+eDWOG4ldGh
/sBjJShQkPvx1CX1wTHzM7RfX0Goj8e8SNDGxh9uKO2NEWq42I+Ksh1TEOyv4Cb5
zG17+9xLqAX04VCL0uDpUm3wqfbD9T3Sn496G76Y+77o3JNJs40BldmyVuU5ISe7
/Mnn+IdQAo8W5a6RTdRKgSTV1efMHOCzC4z90aSavoE2XRt8Nq8qJ4aWt6+T1wfV
IpA2E/d2XVn7FOm538T0zGOApgtSI5rfEte/MdE7FaF8pnRf4Jt9xKOL+vmMlT92
Q/13xM8HCaZG+f9k6hairN7i+Y75YPBU3lnDcOogNDOanJFHV+Z9j5+d+YbU5/5q
fehJfqRp+7j+W9U/zy3y5rqEljcgJ+yaYa2Iw6Op68gpOmQZT05AbVFTodN7MKq8
6D7251KOCpXW5DTxproLU1BS0W9/d2c7JBiEZIGrt8QRRF0HwevK4rJOaK4xiWoG
KH0QVVL96KRcEY0DPEJ/GuYsekxTfO7j03eJpV+MCpOyY4W8l6r6usIt3oSzpJ3o
bpzW4aABGPhLHG0OpgPq9OqC27rOqdeQsVO5sPAFqz2bpDRbXETRS0c1Yx7f7SMf
LYfUftELrRA41KXQ+wdrb5PdEnwi3GLQ+0uvOoHFeBO9hfec//mha/bGrRLAwqqt
WfP1AeqkjsuEy7cHomfvYem6xiXbQPWhcLDddyDUa0nK1+smExNX9fELHBZfBIim
ifom7noa88rPVfPYUvm3JiR4tlCNhm3y17KvLU+ySBsZw+bFy44pCyyMD2JdsXB+
hsYVniJF5/BTlecMwVeOSqWFyFimsUuuOnqKCYj3I1/vanpcnNfuJkS/hBeF6I9X
JufFRoDrAJG6yaPqKkgrAnbtk7dKfCBoDYqhW9LeGiu7n3OIbI4Qt7Eq9UAORedT
rA3GRAQxIjayPxqYz2GqKshekypgPzbIQtBAEAmeJ1N9GbnJSTVcBaO66bxumj/+
qYEdYjBuA7FED9mVeD0ZHe7GHuKOcJSssGo43ZJxOvOPQ9dTc+P+xLqTmXe1cTiL
4hnYzoeK7NJ34vUVe0Jbj4iTgZ8kxcLImM6nidPrj3kRNFUvrMe/r4cXSQQLkCxQ
/vAb4vHlT180eS9prN7Z71VdYa2LFBb4HMt6gLI8hqGjmiwfsdALVAZW+If7VeZK
LSxBRMC2vcMrk7vkU5QuVlZEKZl8CmD5wfRs6LzT3jVStO3LuvTQXE7djTBVIpMj
HnfsdXBLHk1Bpe3Rs7tz7QcvatLx8QJWCa1jBMBlGPNtQ22knMO3IVNYb5ve4ji3
oqKdd6RuHEXeQ4yl0n/qXulVqXciA3pCjIKZqlhxhkSD5bZwhSDFKKQB74pAbUf8
9d9ibgUxMpiP3zU/EAKYpaqHymUCN2bjWb8NkxEOZ2Z3sRLiYzL4+e0X9SHmPbVS
OnN3jT+BkkrTvZ103ydGo5PHlwhRm+4WeXPdJJBQlbmdgVCP5nbhu3L9u1m6hQow
VS4Ks1jS/uXKmOm5rhBey3jlmzVbK0cFwc+zAnlu0zs4gk+V+SCIB/2anYQ9yYOr
DFld/iwbHXgBj+WHUROJpT/YUJEnKQeplzkMQK0Uue7r82wabwDnf3P/QiT/8Xdd
oQpy+Zhx09kT7kKuCYlKl6RyZT2v1y1lNBMVAeoZhygLj+1IldfaNsdy8F50nG9h
FsPVeGw/YjRkXqlXYw9jwlNtqXeoEYhtmex+bcviRI3UzBF+ZXA92u0Oasf+wf4S
UEQry75wmIs5hG6Ot1dIuaiMYvQuHakCRnZeMT/Qo0Bqpos2HlCCj+6aTrYRrCOn
Qi+BY+kAZHnx0eouSmIVjiOp0zmZFw5GdI4bT1q402mK18Vu0cKH9lyZo3xMBW7o
IxO58b/+AsWmli6UYa1T8qY0VL16FdvlB5iYf5nHN6waPmwT4/Eu0iKDu6MNYVBr
3bBEP0twf4vqrV/K23CGSrcxDgkAKOX4MP8DHTQCLmShzrMw8QDA/vXaJZB+KLnu
WmXQ0TOXgo6VBPUWLdIHt0RmbmMtrvqVyxm+fPyaZ8ZCtYDYJOMm0ENvmB9Hr1yR
VOMfwq2qu5KfqTm4a9Xp7j7+Nao6A9J0KvlMlotgiVPH7apwzlcrd+b2KbJMN4YR
8aA4U6atg+OR2vlVapV8FiTV/hvs7r+Fm83CDwjXkD2pM3a7j2wjmjQbpiouL1pp
vhEaQHyy44rwezxvHIVQxmuz0HBXcFDrLhZtO/PRqKoI6ifApurpg0L0mHs3aeey
s1wY34fixv6NxgJDQ1Zk0CrH64fz4y5SVscdwui7y6LVwTVFu/UtqYE3MEQYKSdn
Fm18jfwUDd2iHIglI5GWxEXERbdIsAlzJgpzsXHtFkZ0FbSENWHpULNbo9fVLW69
jiEbTGQBmRicTu4ggJ3ngPHSQq6I8NeQUgESe9X7ZevK+5PYbKF6VY6bfWr0iO5y
lQ2xraKEC/QqPH+Y5GEWiN4j1aZu4D7czuO8d/whXYisUuCt1OptqsdAy27ag8Z/
dRN2qHmGlXs0HhYek9t68cyxmiUN4FEUoLjyYFPzIzG8ECNi6IqmXxxeteGJ7vJm
OUf++Uoh/i/9pPi0OLcfTqdbXj/0YmQgUdts+db8c2zfnmvrD76YA6tmJ/Mt/iMh
Y0LY2IMY9oQ/pRH1s6xJvWC1yUH9GuJmVLNF7kzTsotGc6kf6XGEurZJ4jJUkrIJ
15bal+xSSebVaiYkK7OC5bFMWr7B6S+y7jKO88N1zJ1U0bnP6k93yBICLEQsnqbX
HNxf3GjjanQcsedAu5rFvJXQV+jgvjdVeg4dgtj4AmX+tweHt0+h9TbYXpm6ulOu
/gp51pCGEJcQE85/H7+bOasu789BhZz5/x4hU8YgW0lKpVrVIFZzrOXmvcv4yzvv
Mi5fZlcqrYCO9L2V/YY9UgpaIJIjXcKWMdc7xmuOvlTCNwnJ7VsYJKkWg1HvK5t8
d+gd/zz2jSeFHpGTShHVKbNwmYw9owuhFqQc7JeH5n6wq4lXlRye3AMHkZOsPmlb
Fduh9mYgPjJRbZnoDITjT8NG2+6NPzJaeIRd5/VG5R/Tpzqi7hmveIb7UdiAfIOx
JT0q70FNjGAo6cDOkQyWrJimsoUT76iS1vlGj2fSWRA1daWMhu5M/gVopgBdZh3P
7/WYA7lQ7r2VIgZsbjXFD8nyJ4ZzRwwFP+P/23TYhc8=
`pragma protect end_protected
