// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:44 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ek8mP6dCX9KY4UGd6dF/os63sD6eJNSv+iu0QulLSHzYKkse42l3fLby5KPOQD8D
rOGxrU2LMcBLgpGkzlu0/Dlz0Ah2uQnC7HnD3UNAXJzCCLY4KnarQbSFSIsUVtsI
6QTOe0CqLxSoQ3Ga+0KFWpVz9MiPdqjLvFZYXAWCxq0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7824)
CYGvz3AX6Rl2QWnp5riJrUOQCHL79KzsJe4PUIKhhOZCJm6fh3e8P0/eKq7ExdKP
ciKZic8nd4WhBWheQYMwHpqnLdk6BgNcqtwrzoUpmaon7jR1at/e4LbzKIMu6ub5
q4tytbsxII4IJY07qkj+VJ/q6YliVWVBWUTC+L4dppaCD9iFg+KPpzitoHC6TFvY
ucFPVSCqVlFfrrnrpizdd1LihrqgjL1gRlAuyGEJ2H38gVJ3S/YPUpiS/w5zTj2R
OaBcqXoh5HIdV+3XoHE9qV4wIbVj1hIOLC0ovVGx8glgrSh0gs6BLX7zEU9Tq2No
4xaSqFZJa1mxwpwnWP+CgnrAI32lnz70mqEUu0fGlK9m0nFq055LivCtXkgjCK/b
CMxsyekaX2cBYJQumocHtxLrKKwMV+jkWFoF9ZyHyOVs6zATk42t92GSjzxH796U
ZsBirjJWCcpQK/Dbk9bGAYzFTOmL8rNfDYdV4omsC6b2K6T2Dx8Cmr5WMll+PQBF
vkyq+KL0FU6s+OX+F/sMtkwcToa7DpuV8AxPxFtXCTJOC/Ofpol4qw1T+sQW6Aj9
z3N4Xy8HUe9y4I1Wh1T27oBhfMxJOfX7aLDJo4tiFDjc9EXRGvbfB94teVHgiV1S
BE0sHr2P8BcmRJmqzexo0jcZzUcedreDGXIgJaLYYvIsOqguDthH0l95v3gukthA
ivKHr2IdGIzxUFaQjiilC/do2OecP/0O8ujK9g9gtLYNDqW00JPzW3WRXgsa98Mo
oFiEscYPDt9hr2xn7T8KFDrDqyE/vjjrXJek3qp8Zw9+Z4hmOW9OLAfjUu8e2kiv
oAju8Bhm6ylvF8Lu4adRYi0VGl95KNoJfofHaaRc7ysDfTvUnuP05V3YxQpwvShQ
aQZ8N3aOae4pcYRcP77WTSzCPDRjM7VFl6Ty+5Sv29DGEiiE1g3JfDmU/QuSydUl
fPCnSTarcFQSvpc51p0tpRIL15e1MAcE1oh/SGRGKl7ir/PVcyAczjSiCXz0pFfV
8MK8DDpL/4sqYm6LtzxRKM0krJJiF3NX2q+1DJGoy2PgU92Ih0SH+6kfjMM8wTqc
g4g3mTT25kDY6IhyfvKJRtd6crgu43Cb9s+yv+97lrAN1ex2vWILt3cWLsqOq6v/
zaUBL7WNOdOrlB3UFd2/Awbgwvtwrqgl80toorA4cVA0nVD3q7tg/rpKB7tMRF3l
su+Ktrnn0D6kDPZiwu43Pl6ZBikkTN9J2zVLzx8wmAUgnr0urN/LhEsyR1+ss2sN
5vUdmjzll7J2S5iR/NQw+qJvoHKu0mJp4XvkK/M5moe/VdWY5qlDcRH0dMFLNUJf
Mk97W+DSZ7GVhsTGRjzxUxCjkMyL8PZmje+ph40l/tZobe0UfZM+OIOL0toPnMwB
gRaymrEmge1J8+s3JQqHqEsHDrUI5kYD8Mqd3Qx6aynCS7+U1V+ipKxzjGiyHPIr
nAUr7/C95041I2q7xjm8puLbmmBVUUlVngpIzvao0Uo1Z3NDm+wqg13hDZ7wI4PZ
tSdsmD0PEb1+ASu2S+mtF3OErqmLcwR9iSiRz5C0UCxgqwuyrFnOIRGOrWWvPyF6
cBcSUSHK3U2XaTgMky7+gmLUceY00t/Dx3dQ+wxX+V3EHqmbHCLUDILxUIzOT12r
no4Xp9S+MF4bo5vyNBnKfNpVdPL2xFP9qxoQwQi8sAd5CUT7U9R1cIBgNvSTf07A
kkV6Yqi//za3OMa1cm8sX2R0XqN7rFJNq3DlnVXSauKnwL7QogX0ZeVeDB5ELW3M
xlG0zBIog7hSsnBVHs2FL7SPZ2+4BE/sC0L3iKRyQIMuYfmloX9ThZOva7BvEGIp
2WCsP4V4MUVRcBCYNyhNqVpn+QwxSMRE74bhcvvpalXCKBv1TXXQb8apTSV1p4ej
US2Su6XWl/RjVvqY7vz2Egu0ZxvqeCFrjWknDn/s4qoCYlqQMswZTSqCIhm1FOgh
21941xsPoiJefFAYWRGp59LNntoU7fsPzsvuxGW/P/0BSTiocRWtDB24yF120SRC
5O7XbKcpAdM/MBuUnVaeq/F46FfygGBzFT1izokNOvkb+48aJ9UHX9kWO2aBxSne
CF5ctjd/YMh+i3iZZJq8pkdr/x+9r4V8iOgn3c/G0dnWs1FgtqjSyUn8iUBMJEgi
wXLlT6qzb74DoXWxjVh1pkMJNy2+eXpBNrO5a4PPVTV+4LlmPQa6/HqGZMfhNR+k
gdk5Q7iyuhBattwoK5ue9uHWrh1L8jDCKMZjsotB45D8bNB71lJliYRCZdx02j0R
VNwiUC4gKKra4XefKHrJlrwsQyBmf8dcwfsjjJ8gKfJUfrsuTeu68KQMOOOLuacg
bxxiDNuL1o4vBGIaS19YuH1lg7EoA0HPHno/FEShIHBGOlKu+4PF/MOiGHx+tyl6
eIwsXHTnXeWDrZeQF6uLTkD/qxtUxm6GIt4rQGRG3O9j2OM3asmdZqPODNouCKye
i2byJJRocBrT06paL3y+Ab/d8lXooMkhaId7WF5xRkWpvVVIkPA9maUzKo+3lV5f
CEitKTYBY1w8FwA8FGcO5KwjlKjsEioiULgmOBBB2RVzcXKtDMVRMiRgdHcoYj/m
mmGF6Q0YqOLFDlS8jnd0JzStjRYSQy2ZqNlFoXNRQ0h0h30CBRQvnnPd6SAvPtG5
+J4zDvGLOfJrcrr3A9BWK0tjSwuBieh1BXlS3dggYf7mdbf2WkmL46kUPdIhGmf1
XmxM6vhuqxQnV5E96eOs6TMaJAJjhTA0ELuDuQkH9Pt2Igd1Amvwh3xZQfwbOE+U
cCXxgiFGgAERN7HQspT0oBt1lyBxpl3A9XUEnu6SwR78qfAu4tbPprxBnBRTVQ0D
SLuiInJjkrTZOWQeDAUoED5VU3OfI7TRlu3cStVbKlt9lksLZbpxEheLoY+P0Hgj
d9M5DOrPDZnMo1M18CvRajEWXbCjt9uddNY6OY5GbgKi3nMn1PrpIjJppCgQo5PR
d2v3zP6UfGbkmHN14V/4dbjYE7GvNudCubbnin1KuXMQTnr0cEpXM9sl20Vb+JJ2
jc7/gqzPPha+1z50zSapxeD6H2iEnb+bIulU/EqRcf2e/ZlhsHt8DpegX83WFZzm
ixD1mJevKJFev1qNFzyqqInSR0PwgzX+W/0mTR3zGRXSzz9SSwQyAUH1Z2TldqIp
xaKN/bGXYS5mAyWwjSRB/tQziVaQwXIGMNtK2tc81Z43rPB9MKFK5G9XP0lOkfuX
iy1eo/EGHqQJ6B/UvUwwzdYo4/K06pDCAI0w45CYXPwW6xGxZlsbO4wftmv0ZzBh
N/6HoxGSs4wOn4LdIaomYpjuY7kC++zUrDBzdBZmFFzszB+ggkFr17lMzJmNNcl7
mWc4NOhmc4qYs76n1fFd0M4bCJVUbDrrlqANlF9YceEQN+luoDKnw6jkOW3Z2s6P
tH3TYIsx+GCKsMk5V4UHgaBJA2yFreOXp6U2pzhvjA7oGan9a7ieiALhKw0Wplty
Oj1feqkIxtb97QZVhkjWekYVlBAoqOauKlAlKnFRtxDddQ6YcNizNwXTh+BCEOCS
S+KS3yDnjOmEi6f3adlwAYAAmahGHb/O9YrC+tYDMcbIo7ryN9DSgL8Jf+uIljnc
Nr0iaWycMBc61rjY3wwPWmRZb5TUxclwOqxZ3dY4Rcl6McmA8/Y7QzDkErhMmuD/
9Ssf6PRs+3o9btGQT0eBCFQxtZE0U4s3tsgpA2ekwbbEX4UUWU7A6YENU858vJQc
9CTtDvYT221SGvcLNGmSSRK8u7dRR293E2TyrIl2U2DrMTzDoF0+cxsgycm+NH+l
I06tqvBkzmiuO/X0WSRLqyonPA4uuG9cYkSlchmRO+JoEg/MFLasI54xSpZ0eju3
dfzSV8VtvJAkKjip+j8CKiEGjUTM4kfSTB1MN6hS7bdFAktOfOIuCG+YrxzykSHL
m4v5fPRtI5YT/PdmZZBg2s/eyDsIP9udDHUiYcB9kKTsHmvTCYPvtdjI4Y4BVtQv
+6yPTE1+/gACylqvLUV0w9kEq1mdBQdW/CAOQT4nUCK3enrYDr9ruWAbVPK6Al2Y
e0WNJCipitZO9l/STP41RxZpM0eYfdv5412Tgv5TSlu9asFtnVEOyG/d8U5bJR20
MaKmz+eB7OpjvYjx/slSDg3aUGTBxplHM3RWePCXRI0dJY1enQLBq5o8CVvjsMiG
2AjQ0EltATdeeE4zS8gGtY/X9oNERZGrrDcZGEBaAREChULClPpKcCYORv/ULUGL
WEg0E1c6sYjLWR30VtM5873JQK8McLs/fqMTHGFWeJiU6izBsNEv6TXkD4ghKbFq
6FW6/6Sbjwrhofw0KnNOnqMkPfXCwruphpjvcqv/1tS7yMobVYO5OTeWMBBbHbkE
TegBCyJ8rcmyC9WLdTYgOhGqMfa3b99gUaHIuYm8u+W3VAN4WlOeZJveNFK4M3g6
nPAoieB3t02C61KseCa2QjwpXgZC4EwYpPHjDBGHb9/LWTUpDIy5jV+502I66NAO
niC0foceC1jOB876yHXSzjW5NnA9o0+4vdXHhqStCeBKNoeUducm/RGv+a1Lznv1
4XJV1d2B2IQ4uPRW3awM2wODwaapg6gQ+zA9WEhWnTlNeGg3wBSzT+BCleF0+afY
H7Ydqd4ZXxNK7Lv2Mgpsk/cHIH1Vm/8N83VQF33jCiPjlTk0evE+zie3D+HqJJB6
Fo5cxwevwFDaJc1QPT86T+X6oK3XVYgdIaGrIezTvGm7sTlP1+1CP84mQrmMUu6W
oGE/zbtbwFUHj7xjpalUFEC/Zk4IOg4QbVZqxs2SjfcsNZuuorips+ZaKbLSMpHV
8GnaT1BNyVwJBovfuRrSPNJ8p2truLw5sazVQAxQB8JsuFczjLfk2TLDcrbjswg2
Jrjk2KK/+8EHJt8o0WPBwaLFpBonl1NBP9meyh8y5Q/WPhphhRFDxM/fJ4u4YzQy
K1L6Wx4RVShumz7ec/xaR1m+Xxmr53FXN/cAHdhxZ++NAQ+FvNvi5wWiw2a5UOw+
L94QoA6HzG5dutCTVBnL2fsQ+ZwaJgmFw+1liZZlQmnSlTA10k2NgFPIeCyx9fKS
0S7S0AQ6zjZqMl7fajSf/tAHi8DchZH2/O6tR2dKTMj3PD11bDe6ypVseNgFuTXE
8zK9fBVSQ0gEQf/UGNWD2jM9ooLj1hY01aKUqydyFbdThSXfCx+pkRcAhNUgQetz
ejPWV8fY4wV1TrZungxN4GVKYqmU8gRGGYJvFm1QOiyM18ymp5rlD7FbUru2MVJX
1PR+L9LH4nVMd4GKCsbP94hVt0ygcNuLmgUyYBOAWyWdgydsAd45Q/ECYlkbh0zX
fVUDRBb1ljzKxCegM4GL48vmv3jpCwigwFCJJcbFZTQOtuyCr+ZFce5Z+slbijP6
qzYFqwGb47SEuI+LCBaBPY78EGteKthQCSJ7WQdnlyIm+q/phq6aUapss7FQ4617
O78w1I5BSN65TnmhwqZIB84BUuZlfNpwJgo1QAhuXEGwiaEvebELScJcYvuWxYds
Wk95k2KbguIUVrQ1qDzFTXCifaL+rqkYaWN3wbz+e0SYawsrDBUkaEucVDMNk++d
TBLVckz7RSOtz+6TJi+2/ihOF6d5GYBB6154Dg9m2faG0wWCLYR9wO/GTy7YVJ5E
kDpm29x4MPCnYLoUAdk/FR79DBQfU/m/NcJ25Rt4SWpS3Dss8PDvMFB689YSekDc
LMGQ0IeX2WXZDS8mVUPzlyBqsiGSRni69RuAyQI84j5kNXDIfoyGL7kkhkZbl14l
SRZyejDQmn0S+GWdIwELH5kC0GkXzQfxhFWRXBmtQFd598WTqaQMTAfvm8BjNviq
oY8DY4cGc1uqgYOfLgUFa3J7sND5mpjvsvkv0Et+X/DcF9IyHs8McFuU+7er0LO+
7XEmU5KqshmHkGOCjV1mJrIEjH3TH0wQN3UouXvTpnIbbU8FKO/fD45aIOuKMAK1
mpylU0+lL6UbWe4fQVtoe9CWWz0PvQe1BPTbdKTtFH3ZzpnW8bM33UILdOd1x4Ow
qwV57pOt0mifeqqitHoBnfMkjf3aEm+8EKIBXVOeTKdkoVubZ56kH7Wp7RKhRCtX
HWy0seSKmqcQErqLY8w4c/uAk4AxvnkplqPhqTFOyccNlFQLmkr+Bzxk6gCHqBr/
jbZkFLt518EvyeW5Il96X+9/DRwnj2vpRu9JM/pstZjqOFzG+kLSa3ZiGFUcMt/7
zg0jIscZ2o8gGraP44WVG9gqlVw7Cv1kRm7S3qlYUQIXeSzgBDoDOTyYi8GO7x2I
bjMJmdLs2TZYeThrsDnNSoy4jN5e5XN7N/VJeEg1jTzsWZjNfhNer3Oln/6RO3BW
xsjSPsQDNmAmEx2yNDSLrx0adC36wbT4PIHIP+2V7FCzZXdsSc+AndSk/ddvE32p
v3uG54U6qPDdcq8ehR+nbTX5v6rp9cyE5OzOv3ouvxxi7eYih7eYWKcOQeggknPt
JMkqjT5nYqmVFzo980qRqRK4w31oTeJJNIJy2V5W2W/vYeIGDQ86LML5ixFgrF2G
lq3pPIMROkyGojk4wfFJbFgn51g6wEMrpenzBjRQ26f7asD6q7qOBjyJn03vzXp6
IWsWKG6coSzsBQ9KL2uPldxpyYvh0iR61+9EPOWwDDocAO48CsE+YbE6Cu+Ti9fj
ylzIEnVDK3898oAlyxm3Wtw9w4kXJa7zsSqIUvv+LW+KHSJP3VMd/kRmJ81RZDkj
N0+Xxo1iac+KwQUEehNozsabtD0SDZK9kX9pnwcHe2V3INFbkORA8nRnEYMm9oaT
dl+UShTJZEBIEB+4+D6Vs8clIUVhvB1UIipdFtBmq3mwGoESyjPxZz+Ns2eE1Ul2
rcZsn4/CGjwAvzo92rBK33hKiYbeSNgy0/HsgF26BA7nCYQSUThV9zbnAez1QG06
4e2A1vd+6Xp9uKVeGfI3Z0EN+lXckXnWI/RjVEvTFf5UrdpvPQdEZhFUt4N+p+jX
C52uvyxVxZfxxcf7k9PzDM2SNhJGB/op7MUBbkTRAVtGV9kV7fb1MxlioJU3wIjq
qo+JHUMV4Qq1mNgOLyDNluH6kJivvSVAaj23oMX2/kC8RDsYNnXEWWOmcN7KNTui
a6Ao2lAGM1+BA1xrmkeLEtIkqu1jZy6qspjE3JdYNmlanZ/keMaDWGRRl52lYWLM
3DlXIvkgVHWt8cr3umY0+CNqvJbBo8PpvlnY1Nwo2AKVIYMykOSjYHKD/T/7XktO
1E24Zx2tMrphNsxkSfQTM0IYpQVhiKHGf6UrQxbm96HvKWo0eJQ/rPlTILI+8y3t
0/A5MnjvgjT15uDedXtaUS62cAMi000LbBhDVVZTB2T4yYmcUc/HKD7FT6UKj/nU
E6c8xRARjf7uojJ+USNflnFTkbuiTiWyjM9x26jV6AlsNjdXyhjQBbb+wwYFjDoO
3T7T3vhtu5bG1BPSafKpRnqH6sC7uA5O/LXDWHwgP98dwvp39OVUpRyzqxjJ5Vol
gmM7udY/yOIkGxyPWfvTIMjuh8IwWhbj+eqIZIagVN8WiUKW+Cl2AXv4bhBLvNIb
lXrJrqg3U+Uan70e2ZobtjItuSXQMndKXm4CEyDN5LzRwFkZb0R05Z341lLy2/FW
7aNN3PLwZrGRqEHCzWSWfXVNU8O0zLIz/vkxBfNeACquRXPwAbVJCFQGxzgVW5Vx
JfYyf93aMgoVfQTf8SWejqieiM6Ie+6QF3XxhZgdlk7lfwNHYL8044OWsMuK3MTt
Z5Vaw/IGOypg1m9vndeIlNo+rZR1VCnYY+LjbFzQadHPtgH+WRxP9nxlKwcAwCwm
G8M8Qbn1wOY2znzZih6QqgyUP8ZY5e3pCjtgpcNCN6QuSSnF/cBL6I9jKb0JUoHy
kZ5NSqQ5oyekDcBy1uoGAbnia4sbF5sTP4QhObfA6BWL2MLfBh07LcoZQ7m/Cttj
3dMJ48zA3QRpq7asNrFeUNWyLczwJFLewP0Q9AyAWqRgmr5busCKdK3tilK5y0Dg
hQQ0hS4lrlcYS+io/fz3V3OuoYo8CEayuaq2OJ8ECeZ0Hu2koCM+ksy4Tp7Km7x2
pAGOt5KbFevcU4dw2A5ln2q8fFVFPVrBWUrIk0m/l/2/ImKAWS3R9r2iJ9PWQyAd
X5iOBkVzkpkFbfUMBQuuO0FZQTbZcWIrBQsSeLSZTz5p+XM0HGGkmZOA07JvyaYg
LxX9e1h0E7m/A9Er0cCpb21PU+8bP9SczYmE2f4YacRDp2IbRBTua53vpS+52EMd
WStK63L5xL1XJNn7GsitD76OOUf0Yi6icNnIZ/Kr3ttDvg7PaMMenIk7JYbgQ1MO
ZI2Z1ytizRzf95+1PqucTV2JUgAw20vQZdf9ScrImPO4/9emwLnjYcr3ZdmF1Izg
S9erXEvPxDZxPhHQfTgoAYUhSYdEmhyVGMk36ZePFCsIcxw79jbCQrPGDMhhiCzt
YXHZzoNs2wovDY4PX2tlchdCyxfkNkr4SzXZUYX6Nn1n/Qbwdfwut2lq5gh1ga5S
S5S8togn3IPaiFjY4FSQfzmUc6JwWQ5JTklrCXLooDECYug7G6lJYQ75K5E8oEFy
ElWxaEIeeCtAdMJWHL/IildCVidLEDzvmpZVg/FeCWrb6AppxylUI5u4tTCBenAB
ym+eSTQ4QcD5743RVWcupxbL9irIwzSxQ9qvbYjE+ZB3v669vx1cE3jChiyurGTa
rdNg5n3oB1t6iHrQMpr2yrJY3uDUPhpzRor64RcGx7P5SgPEkjUZnmakwG7+7UDn
ZsoFKursV26fGhz0LtorE6Gj3KbaGkZvOejWLdWI0GH1UXqJuSKnYRj45EngzkRv
gzj8HEbEsXzj/ruYZDEkHfoSAUFNBbnxUxrLfWUVPstia6pQWzOw8+pdGuljoKy2
KmouJbPCIXALZpBmqRpY7oYI/qIV8Ar5y2z18dVo3/M6NXVXP8av8D6VEWbKtORl
koJ9dUGJY7+QSi9Sbd3brhpB29fazR6yBYAnxe9bRhp3+pc7OAksNnWwX1zZGezz
1kGLcSvZADT41bRpllrgKYWMfQPSlK+srkDIZCYmtqq2wXCbES7+xbL+JIYejqTD
FVAa5iZeY0dJkvMjaRDrIGmty19dIlYnGNXGI3c0OzZkoUDMDO2RUasay1649Jlf
xkrYB7UwoBB0Ss8J9ON+5VDLaGQeExwcAC2X1tXVmUCCbM5g4vPdiHsuwEv+4HDu
XMc6JTDeTW2C5PTYuetfxcpheIx37gYRfvmqdLLMj8TBJI+6tQKPA0BRtLPnEJfm
AagBK9y8kiR6MQhk0iSMUZ9uOJD8uEAgRNyzJP7vorh0QoehaSpMfrPd2FB1DaHZ
SLxZtsnHi32A9m+J2DZSP1ODd+0y1+4Uiq1y5ouMS4B2O0M/CGnbIwXU3C05CCcF
8jxPpfrKhJfPgbX6Sez6z+2jK2fyJRnluEE3FD/63cp8GR1iocIKqMHj7Dmz2weQ
IKH14B0HnRFvsZ28LjXduvl8UdHTod5JEaEWhv6L9uOH+X9NFBwVin7EPH7rqNRQ
34BkhASEGYRrUJY3ASv0LsFLtgeIEuWhgUzx/num4ZHVQjmPbnNe3tuh2nCwH6Mt
CQLQD2oT9Q+Th2EyTv9Nc5wfHiyOKpu7q2J1/tQ/GkotUAAFIgRXdbIrsRSmblmB
X6F7+wPZdZTwBWF3FuwUlhJraWud2JVFM/9r+wgCzmSWJixsGZvy6HCbOmnoVImt
kKrT5zuTYnbjWVJJboLF2LRXfF7PvO27MXAVRUfe4OMSfZb1Qvf5ikGjSTSAVdxe
YDG6mTqwPvqjmEB82GP4ZHkZkvONjzpyR+ZNfauoXjc6pFYx+snPkz6prK1jGFbi
qybNgEx+nVC6L+BmD9kSUlow6JMWtq7fLgdKMZgPxg8QNusPMXiDbrgqV8s8UoEJ
SGavuW8stzJMQNqdkvuxJgmVd4CUsKoE71aIYkJCy0cFJXVczeEhNyPAIa9LFCzH
qfVWj4Pj2yYKkLrDrkjqYI+5yrRuWbBy3wIbA1h/5udqrAU6vYhgo2hiGipooLGJ
qR6hWX2hoR7qWoE2FpSQNggAPZOMQPfuV4yY97ssX+0jyQzffa9fhyM7aSw4vNX7
hdIp4xFv/bUTRUb7WdCKEEcwCwLMjeHBl5rc4IB/gMC2/dDcXe3qIhwnAoWpWP6K
cTqYFOLAl8bV30w+5x/x79hfwtEO9WsAp3bO+anHMmEPGYSCy5Q7twmEtifp7kwt
HYYuJjxt7sg+CKjnygG9LlszVnkNWv9AEisjHDOr1bbD219hCKG1dPjp9oTCaeM8
E38ek6wSHRkYXCz/FY3q20Am4g4I7TtFaoR+mIQUeUUBqYyV1B68YE6OuS3wuaQb
`pragma protect end_protected
