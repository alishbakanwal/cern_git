// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 13:57:46 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HCV53/Pjupqq8LFh/3tG7p0ynd5h6vo3p2u646E3WVS1U5YqeCVVbwmEQ5L5/uVM
1KMGF7RCIQOOVv11XtSnk3haAbJhCrGDHNOZIDNog6LZ2CF3M5mczgAoIOjP3+1L
q22z9XB+qKv7mQoXrnMSUzF8HO0P4G8qvyVm0Pj+BrY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12352)
rApTHMVHvTG4autldzGOQb/pv/JNny9H7kKmtbfrH6ePG9Af8MrM7oL/jDjMvJ1x
GBTqol4joJKgSAmdFkQl5Jvn0Zzn79oygOHAJJn+VOQO8fgAKyvdf0mY4CVXNqul
qqHpTuZJF0Nd39crjZhJAxnXyoG5YzisZf2gent1o3javLzpEtQVJgpUU3IFhwdh
JcDB4cMf7FsLE4lBdKCq5DI0XodBL01H34kJCYkx/D5IM3c+WfrCmI/g4Qys0QoT
lGGlxPs3lqV/rBac44qxIoR5fJ5SzECRqZHYLnBeZa8tzurrKQGTJrtZfiGayDLJ
xw4Tecr7Ugh4XN0nTKarNyuJkJxpjB2jRJWyzdAeUtG1Rt1l/B9UYp/Re33Vjsly
5HjfE9nS1f4IXUQnI2VGTvR++RcX0cW0+QtoMjrK4c+dSbsmnSy0RhISm8kXrVSd
aPZ67T8zprNPDdMZRSO9YWrNpe+081YfBgTyFeQlOJaH/fUYdYydUM9iFmTPaeoG
o/Y15gJxGTN+m/KwjyySeUHyDm8bK4b1BrCjDJNjO73Doy383Gva/sXozhLp+a2X
yAyxwvfASWb0VfM032R+tfJOgAhEIzEZmUm4OBy9TPYymN3CZGZsYcIPN7zD5GP9
tcYncKEER3n6uOZLiRWr9eudhxKFQOw0h2e77q0j8yB+25rqZR4ibKDmxxbDRrYM
TCFAz6j2U8eVLGuj+qEe5uaIuFAM+hZTz2lgGwGHozj+XZDkqCuibL66DhVdXufV
aGrG6sl9kLSBc3pjWjGJ/yp/N9mVIiO/jcxbasOh57SAA1JZioDeWQdnfztRTmYp
ljb24s46OlRM9fRt+XPoQ9kjllu01g/DxUQ3Spmehh9NxKn66MzQYhCwXRgMLeeB
sMPzFji3DmdWEs8LP2KW1nqIb23aF07vss48oSuqie9Woz5T37WuX2xcOcDxLDiE
DEJLwDvfDjO6ltKobKXSO5iVz0qJPNEWg+lddIDp2hXM/dmCRDIUABPHK8OFb4+P
+NIsZE1g1eoTg+h3pwnHeZ4hm58868VISaXBr8A6Itemt3U51+s7wxp+fV3TITm9
JgGo6OK6iywg2QX8fKEveLDNkbO55MvattHTHUgBG4XTDcqP5I+utsxHBoSCsVaI
6QjKdguybN8v0o9+NGnBOwTgEKCCPW9EpW7WROQ185r8AMaI+jXsMl+Xns2p3Aik
0KrWHpjmTIDR+DFt3Qzo/2eDEl1LCTMF+wANSew5GJQPCCm5enrHwg2i0A5W6eo8
mnoj3/hnQEiiDC7kE7MwWPc9gCEZhdr3TN8iSw/KiMOl4gur5AnUeEKf//VwQpYA
A8Vu9j/F7iLZSiKLejqA9ndSsJAL8X0hMcyEfm8UZXwA2yrUjAlmOpEUFIcMVP3+
+seLovhS0Ff1UiQkEKWK4Iqj4wXjZeIVT1qO9BwhkRrgghIuAVNHwgArM9YTfHib
LXX5lZyZJN6hDl7gxp1JXJvNZhbp4qMCBt45QWXHv2YE+YlSyfp763YQ6JEfZ9rE
Q+iSl8Ww7RbYe58/ZoLjzv+jjn6zljhbC8P49nq+Y5Fli8zoBlbxBZXLwcZees0A
nvzO1RCt14Fu+QHQp6Om6VB0gDRc/Gnn4UtgXIoDiETKzfwArCXCD+MxJNzUfxYq
XNF89eE1eK1r+ADFHwAYwXowhHJSYgJnwOvY9RJBEhsBvMuX4zuphitzQAQi/F3w
ZjwceEHnW0i0L3PSLYKXTqKrhII9z1K2yDjRzSvf/f9Tzt4BU1ubRvnczc8jQDup
ZPkNHagrTBw0ji3BsIWap7YiStAWpuSvbKfePv2I9O8nZwFBL7w6A8O38kcwY/l+
EeKck5DQJN3X3I18ncVJwg0ekwMXMzG56/efEy6dKzo9T+r973MXYs0zGtSFgFhd
NiBzj6tFdnwGuz6baId9M3YoOGG62iMw6Z9fejKGtOsEdBrs51hUBESAJP3KQt5+
ybyrzgDbwniO98dsiZ3Qhnu0o+cVUdz7HG1EUIG+0rt9OAqs6+pqeT3x1pYPWuSb
7v1o2DWj4mEAH49dGG+/uH3+cMtLNArSp+GdwfyDYq0f4MvH7pEjnFL+t6zN+bnm
bm0Uw1irReFE6JY/yF2RGOikFI7viA9I+eBpzocOcPR7ZNryBedmwD3XgG7L6OpU
NUgHTp8j4/hEOrZgKiVqCtq4mcJ0FQliDJiJEu6aJmUtoq9KB41kKq4/2ueTkYob
hlKBicOjiuG3h+3/f6S7pIWRniU1BGDFVNaVNhFpJRwLpxyitnDfTr6slzxrSVvn
s3tzNAfvZABLIe77RHThoo8oKXa6MYsRdth7piaDxXA3TkcvTyOiZhZB0OaQEyee
JdEtTNPyW2kp7geTZpBTVoLRO6SlL+rybIvtvL7P8Jwg6aHLKPjZDuiGh5GG8kYv
aZ2d1jaqsIq4rhd5MY5TnQSShkPc1/8SEAXyNkPEh5FPL70n4OJA7158eXe+2nfD
Qv1UwX7waqSqor7p6xhB+5vURxQW+kcgH2cLd3UxufbcSRbv6MyYK2dRhJfA8B8p
GzM9x+rCMLEkpCOjrSoG1TVl06fgOBk9hAgXa+da644PZwYrh4JOc+P9u947ALyC
KRe915H6qoNyi7i6d/BMJaMyGopNrtnWhxbl1TzGoaJJCmfEP8GPlXkZhDYgZbcm
0/YoyfnF9A8/1vnc6wq+CRwXZCvMTW4kkbibm11/tZENSrhW2f8T6PPVGQWNCz+7
6WmWuTtQK7+jpXUIEUDyD+mdN9SX/2CvqrnzSKnwqzlpjsa+txkZ3NhBexk7ydkx
F9J4YBWe+S3RpMIeJpFFrn3FbCO9Myw+qe914i3Ej2tzYlZ+JkRjThubghnDKWHv
Vo9mdpbiCF2icey19COEXrOYiqV333mlKKP7mliNbvVQmuh7OsIA+qkAm/uzAGt8
rJWT/aPrL1d6RMWwuTXXQIFNmOeSGZ4tTt72e1GOcP9IIlj0cUVlv1+swaullD3u
WjxQUAjaBzu2UaZhDALw0YCDX7weMlLQgYvTwboSaxKzZykBNWJRGr//Jhho7Xo3
xgNpTsZNRENBRtuQ+x/jWbHyop/60jyZDGfA6hK1Vo+UJtO0DtrKcDS32oOlS9xk
8SRW4Yg0BOrvw1Ar/Qjtg7LI58nBIWMD0OVrPw4k/P4f2twBr7l7YB/6IQpviuD4
fH30x6fpWmla8z4rGHVyTwePj52aqzWj9BQTKGE+wNxY4AoK/BY/Zv1x6rhnyd/D
M9/uNq1aJ22w1Ynemh9Ipc5Dqb9SIdKUkT4E07R/GmvYzBm3sSjK3+Sac+noypK6
4dBYQ088kT9rPgcwQmfcZdcqibheuEYF/ntuzAQC4exE6v6nxFNvwVmDGYfO+yay
+OAQNhwlMKCuacUW/bly9n2F4IR3QiEqRfgveBeVZJ7Cc1rYqUz29bMFiGpMPuoO
DjD9ojDXovKZ7CIarN2aFAJ69U/8fbIdq1K7QEnanT5R6yRduVTJbhF+HjX5GBI+
Ig2j31DhMD6F9Aj4f9t2/K1PFCdzeOK2iNBPAlywMaPjAwQVcDPoYN1+6NoQ9tX7
CGIl12YQoXUFw2UCqK881/7BVmGaZ7O+ma0NafI+Fuob1jHiqXzwuwS+D52QJiDz
VZOMe9C5RY/V3Alzpfq2OeXltovYibCALmFE+vyQij/UG3AGJYcxWzUCcw5Qwftf
u7ODrGDbG1ywn9rNXjHh+O6IA0ehpo3mxDgiD5JknAjeOXs/+1xN1IeJSeKLlFOp
HefEv/6Vjtb0QL2suIeRQzTfDOh5KMBz4E3z8ZLmyNlhIISKVddEJK41FCSNE3mf
GwuTcBdIdxzB2MUR11C1DTPJsalCt5Xl4v0v2L9PCB873mm4wS92h2hakVvpyF3q
1xKUizDnuVouSwOrya1SwgJl7YKSGcIqP7uKShR2quFt0NWnhAVbg2aaPwhVI/Jj
Q1TcDtCMrSOCARRVGd3wVxvqbqxWG6jZlwjPpBQAZDMhMEqvovN0XMflgoE2poJ8
y7+FfEFRXyQQSUIO8GC8e17jDNpmDvFEtG8PQGnTUZ8teapATWzlNV9FeWKTLPE5
Pzi6IR+ro7Un6u3gadqbRqreefhMylXS1Ayz1IT6ealJ2ES+l/epBdFlRqOhKf0V
IOzyeSMLS0zSs8SvUn3DOvNeiTz7ztTumZMkd7pAFkIPCsRj4H2KhmNvmSZ0iTMG
mV9V8+ulqoB7ryjc/pBPcqRkKB1sJRRTJI15N+VE4GtV/fSeA8wfSe6MnoU1v6Ai
OVhj2mg1a49VfrPSEP2XW1cSBv5iw6SI2JFh6BafMSn+t7kaiLUUNksebPCgHwL2
T87QoBo79IOBvsKzoAnhrINZjBNqZbqJKZEs29Y/7Ri+kDPkSbef5/0oSBIxPg3Q
/u10FKgTu7i47nIDma65pR25yAevRaYZaBzlzq2e2ganDIGQ03Ok/JzcHYkD1Omm
oI36Azn4A1n2OSXcw+wps2WQlQLmbF7FljgXuXVsrpivyud8UjRtTwjdndqYe19C
aAfsPJTgdKh116Buc1ugm1aoOpnL5enUqWnme3IPsSuBOoj1xW2kdYy4A7AfZfGQ
Mz8h/53SBgHK2Tt/cRDO9HOIXlbqhGYlXWbAwo/kMHMebF+KeWjdT0PdaoNxvO6/
+xQ//THdfaHmZPXo3rE+dn4nbZjmXDOxuGBnEY2wGvLYR9934s6QZinXPk+3vs9m
VOfzW3GnQDW5HY0Y0RpV6t22Mo85jUiG58BQNmH0sPWvOhrH6X/+X5X1U5US1Mqf
pY/HKH4Skjh5Kv5X1M8Bod3LrZjKaT8bzIsjXNvcWQbJyXK237T1dC1ECuxO0U71
nlpXMcHNZD/1k74omqNw3Jmo/GFkU1diln9JwZ2txyoySyDvH51SHTkhd2EspNTb
bvzgKSOiCkOVL8XxUSFPlxFwaFizw85YV8hGfdOwasJWLOgAZRSG1mPUWCrbVRTJ
RoxbZsnb5nzvyfN9Nkmo3X4exx26sLjO0riP3DVvgBkGUYmiR0w3DKLdvNZ0QXDY
a1T2Xxid8/YUTxI86vb72bDyaqO44Usz234i79W9VEL15foOC5U0tCpvWUALcU8L
kvaOT2yCNnE98jpztL9z+MLX+Y1qvSGJ83qCBYvuH5Vdm1X9XC/SFHB/v2XWac9S
ZvgFCFKUujQ7lmlRYUDDrJ5BH1PW82XCB7FBWpoJ0JbiUtLeLmNVt31y6IPlOZJA
igBfM9j9ivNIgeohgCyk43Gzm2e+7ASUuk107SMn8mBKH5DJVrc8YB23EvtLmwUK
PcCy1npUCYUQonxCPezXDQNT4dx0D/14YoeKDsPxa1FyUChyf/FP6cjDLxo4s7rP
Xw4ATWZgLyYaRr1mR6H6IQXRzHleji7mQr7Bx2XctMr/E7EvdL6gOdgWn351yfyO
vkBvTqtlLHwyJqKBpC4twapLzKAovtV2O0SAK5UUmdPdiUpET83oS6NQerIx6mJs
/so8qVHPTmhG2OjwDnSUuQLbHusoAhMpuFiU+D6NcoicxHxwY+s1mug92B1ouSHF
+bLerpksmNatrGjUK2Kb8NJ2OtUGIv2NDQWwaSkbhfmvRJ7y7DivUnKOXTUvKx2+
SU8mChzbH6eatISrUD1bZwNB1h+WaLjSGK8MdVl4NRC5iKxVeq0q8CsAXclr6FfQ
niHk9MHlQN9OTYKwnEA6mcXOL5ozpYqOqtqZO5L3V24yBU1x1ftyYokzlumOGggs
LRCg97KNYg//87ot6QdkjpzWmM56RGEtSvwqrPjIZ4PeFmn/S8YVgHvKICOPViw8
uDYZMlw4BCbiMjegSeAkLeQ0XnLEN8MF172Hgf287C30QimJRQrjVT4iDMbzobwY
Zu2hjP5Pl/P6Fa9slWKevb1nQjBExHFKxpF4alr2pfXwzg0S5QRvVjlvOAiRs3Z5
76ApceJZYkSuew39jYIvrqQvNiNRuqM6UF2V2e7R284at82+1r021noVS9DJMv9i
1oi8uGVKiR9A04GJvH+kvD6pTWsf5GB9R49yvVtQzbSjIBffOZcr+gzFvf7l/NbY
+WvrpI6aWzHWZ5OUwKfjuzmOF4BKRIMW/3fk9ryH5OUu5LXBBKRakW0u7CeO853g
sXk5/oRk1Ty4M7bKNRZa0KZjS4aLEnum11duowVwmOYVK4cKr1Yxt2fD2eTmy6E9
ycbpHjLkW3GzE2ESdNl6iIHFlhZvIdVg9HKIJfXRSAcMQoAvU8DMJKJHZ7YFoCoh
eVCbIT4F3loAxlNF7xxGbzD51RUE6435VYFUOZlsYHWDo3m/XDusCYpkuOEZOlOr
Fo5lkByyiuQWMc3mX4dq/9Tiucg/Hc5hMCUGaWkL7/MYil6BzOfaAScH381lZKvl
e3uUUFGOn4fY9PLf9DqUve63XcDRS1erD15ihnQZOXaaLCRsTZ2RrDSboqu+aQts
XH1YT8qSH09bYidi8PIDmpCTVP1xUkjH5hgZhzkKeAIztSS4rAs5T/+mj9PX3HVV
NVaElcOLtfKg8JyoLBL2xz7YxuaA8D1tAM29kTkGbzLfVNoYXnPgvkYseTq0uk9y
m3Fj9pS06K08usAPZ4iI/tp0wVZc2Mj3cjhWZL672YQ2UBtvJ7hVwMlno6rUWo1K
e74GGQKafSCLcNKv70+6S2xHd8eMRTQKV3vOeQgm7g7lCLLyeYCeeELcc3Lc5IM9
HhDvV64mVjB12KVChi0dwjuu2PeYXQFhXWP38T2dGuynJmPKBcQlSRHS16PObAKQ
PugFOkd5mNB5NeTnEOXOgDmPCVcG02LgjEHQwXD5bwXLPFWu3bCspG8FazHopRfT
iV5beZAu0LL0f+u0LVY8hJrVH3Doh/GfpzMy9uMu2UtMTsM6ZTX3mS4Ri1oWbYKn
gAfqaif7m/Yicw8NgL98t62giCoB0I0UbZ7W3Yo1tFw1PuHLkDFtTU3tUObcVib/
ze56mxUZDF3Ga9JrOHBmfBNpRP2i6kjtEBQyBL5Wo9kjLD2r1QEzUJDh6m0xe+VX
iakyynu1laClaFcMaD3Vg9plS+6YQkxQiXjpIBSWQn6FzS5lo43T1RTXQroZjiKs
d0rbQxowkGu2lqrw+mKljLh3GlFBEL8nA0SPh6rdKjnM/l2siXhSZXgExDmCnE2B
12ihp4LnGy8tHS6bdQpKD8JBJn156uJTmihwnxIe68vLm7ox0uV3RxhPd/1gXn7W
VwMPZkY7Gh9vkTYo4LrMOJ5UiJ21A6F7hQfbDor2fAl9RHu5JsunJio/zQk1iOFR
BVTRANowAJobDlWlHzh2L1QtvQ72ORb1znreyWpMzj95q4gz5hQTz61viRwbsiK4
vVIybNuj1GvY1Yt1kLY4xHAs+IQCtyGn9ZLo7p50Y2WxKjStkAy4gtQ1byQvHqmF
2Vvy4p7z3oZMiYGS9y/lJka3lf7g9CIyc97v46cvOUGtkuuJ9e9HXasU02Poi8Rf
Cl/pYm/2EYeppacyavkV79OjI29iR9UgdVgD6MTQVq6Sk0V9CzFV5DpRsUdwZdAe
DTeT3OBC541UQazCyUVS7TVGyl2fq3kmCekSxYPNeDQaUH7Hu9kdSb8oTsVQ8x0q
nW1mjSmYTMtt/Aj+ngWRuC+xdI8Z91/Le7UFvMqQhbZUxzFl1BN97j7UsU77NxUX
wBEHiK5I4kJ0PglOeV5Ic4Pe/VezmBbVforl2lL49LUTnEp3mH05JwRXxRioHx6x
Twk3oI70JA2b9va9IwovIPDD4Ktt0cfT6cWeGF0qk8J0lt0qEOf19CqPEGK7sB1L
iDrGWpGzQNft2IllTybPsZapytE7UUPdacZCzAFH4in2oAdUqguKBpE+eGTBMFb7
iB1woEhqs0lPC78gNwfFszwii0IOswvtoLxBBIEPqRRnGbmLi1WFo0X+znUSkOjR
00Cc5e/lLxD6rvSkEtviAbrrYkGvwYgzsMRcZDNIT1LV/LQNV8BCxUy17P9ddmqq
ZnZtRwqmICkgoSHDEuJm0nWzuYp2Gq7Om8sizuA4XaU20QQ2Bz0vVY4t+It/e7j0
gev8AgXLOcYmKHIAEqu/6PcZGQUYj/tEPrM4W16b8oeIKBn3lqKB2sZ2SK9Q3Ok0
plIiXKMEeSft1WwconzFgkE6zAxJCWttXl+3mGh30HJMmtn15nFFUFfqSKd88SCq
X4xw1ThmrDEuYamr8tx/bGBWr0a0rvWQKGvvtnh1rc7ZSCuoLkznXPWLhmKa6mFL
VnKKN5LrA6T9oz7K0WuTjAhPyVlkSma7od4wK+L8fgGBJA+yxLo64/cyBLuDNdf6
RYzFBwC7YwMBRIplMFLgmqyPZ9Sd4MMOBTEz1q8nG8cNNV8UbWYZxEIcQrArD3gL
/NlBlAoeGJH0fC5upFQGyar8cTHqQiJE5xVWW4qO1qbCk+Qhw5Xjcj7qR/8p7BE/
mF9tnYUrOpRzHyvhqMIq0Rj+n03tWWYBzhxFDqp5zZ/215KPZTCB96TKzGMtRou9
sfJDqDxqtD7UYqXk1v7meQ7T023jviLj8ZE8VTxjkNIVYhwyg+CUFGi/jCHuW+2O
FhlRhyCZDfVpjMN9tigazk4vQuchFSeuvA4xa76Pe+jpwTUdl+xsPS8XXS2Y4Gbl
s+yE2dCyGvReXHO4XhcHBYTKnU170NKU2ZHomqTZvRoaAkw0HdZIi42enC95KqT3
c73NjBiyWTzGqQy75Ai8obj/CpVylyVlQk2bY/tU0crx7CPeRwEX6Bc1WLV0G5kP
Yq2DC3leaXbGlSBw5Ylj5AtvwkWmgBbrfRiuL9dc8eUWucsuJ+3KVQcYIoTdkosQ
SG0f6deitWke/eZgWbZ888m32I5PR7WQUQedZ2CyYSFpd6AoRw+ED2TrCOqXNfxM
1JDM7B/ccLfzx7eCFcTWn7iWexDqV8zpzemhkE/wMr9J6vZBKaQwQkC7Iusv0ASJ
S6TYt5F3O9hlM0Qhgz3v/j71HjkMXPjs0k1MkjxbBGSmHlvjjFH/TNwGh3ZfJHn/
mLVNlaO3vpsnRkxBb9n9a1Fvhgk0vuIj70oVNMP9gqePtU+5k3h0YJpPjbxOB0qd
TIt1n4YEzaTRU8t5DXWdQA6XYBiVUMcnUKakW3L0NHQBoBLc6Lu7WOBkPeySwXhr
ov7GKmISLVyfI77bTtVOgqFxd6JOtdkwfyogO06l3WFVVEbRrOXSlR8yxKg9criZ
U16oN37xybjJo3IQR/J1KY0HZFa/HauMW4Ze4JQX6X4txA2g4Q9iLYs564b9wLJU
3U6LPNuwI6lxVr7xMKMTouhvOSObMn661SBDnJ3NQ+bS/pnawsZ4Hg6O7/H+wOwY
H8qKdWlcpb86HZB3YdQ96f2JPEs+GRu8W4Cd/Bv8eQ9sZVe+ifKIhjbZr7jl3g0r
H+jCsX92EnZYw0sKebUy6e48b/EJGzdxNPgvfRXeumF2HbxDKxQei0KC8NygeTsv
ZHBe/K2p++8BrO9Wwad/z+8oEUIgy69RybsDRGRE+trLJsrSDrbfu6AeBbcEi+sd
IheIi4dcrk1EmnnfAESiWzS2S1qkJKqy8cy/lwEqUQSvxQ8IsqbM4EcrP7Xl8y63
cDjZ82Gu/YTTgefmaK73DlkIfxN9FoeET7BiIfAT8n2zU3okR/TMKSQGfl5drBfv
WYuR38GrECTkXV/GtUnTjSBngpOmlx/9f/WICN1pJfB+C5qP9KUv843nUMlzX3S/
eCKMrL4JAeBh4fvi3kQIivjiqVUPHD6TeF4TDBQ1VWqFzeyf2W2h0V7L6N3tnenM
WCHVW5majXYQokz5XdzNGY/VZJ8gBnTgjYPtfD072hCxgMbd9VlDqpUumzhSqFqR
2VUih2qvFG4mHnzrRg5EN0FaWIkiMcpiXgsbGcUdEf9aZ6opOI4OWDBerbGiGBn8
cDQHxN2FJHNe3cU6pWjHJ3mBqCOipLR6Oh19JtKXzGGJ8d+HwGnBfcNzW0dSFNTx
Zi2kDkAN3zXNeCWSR0d9s3Nn2Pblrw36T+QrzEQSoBJJprmbEscFNs67R96kE4xF
7CWiDhAhQ7sQMT32uU9rhPXkyKztsYlqzAs7vmq2fNgmLLOm3ZXtt5b4aNtlqNgl
aexDIzenyVR8KDQGO5tfH8nESptjJfKe8bK5YYspx/C+BmSR5aW35VDVToOE7pJR
zQ4VxqIe1LZzIhd2UiFV6AZyLtDDJ32E3mJ00UQh+HgVyJYvNMfusSRjPCawTez1
9OgBX34zmSnKzjngWFCWpp4c2/DqVbywP198OdxjZRJnbMA4OO/sRC5lFioDLQ8A
yvOYVsZnitCqWlVBWovNGMbWqMzy1+YtbQTc1vzy6t4sN0K7o+hyJTz55wSAOB/5
nWpGC0DbtuVYzRb1oIADI/QxpYxshWpHKItlHnUaHtLqbCN93PDyifAeKPw0MMQE
/QWDPftA9VaAvAGaKnpT1clSqV0T9ch6zsZGVxhX7Oqmt3YCsuo0D5G6xaR6bGMt
CvZxOYHsREE6QCZJTRSiliDUs+/NTqGRydu+tYZlhL/sSWEW83T3BBx/9B6dWjIP
0ql7+1+vVFTvl7YDSouLNnr5IAIP/JBdZyod+83XQRBmIsgL7biIqiz3VVEBzwgJ
JbN/lN7Fq1ZyOil1Pq0EedazhgoX0wz1+gVDqdcx4fVfOMoncORmD2Mk5CjFGMiO
Z1HS+1yEPS6PHSL5tcEJeDZ1qDPDlQwLiNTNJErR9F6IzpO9moVYuwOBx4mPCt9z
V/0N+7PHHaFd1zHznBQ4w/vqIuXMsbIw/c85Q75DYRN7cgYX1sagoFf2inKOU3BO
Ib2lLVba6iaHwG/dF1YvgQaPl6sPPKmyDwSr8ouNANsjpyrUHyH5xN0hHBdMaH5H
8hbqE0PAm/Wx9JDkvSlE+94rYy16j49jyEnG/jghvpuv9CVOxGwZ3QTY1Nym73AB
/yIhoRQIXZQhhhp53umiAZwWGoCscLw2yCmukh0ztC8h9jAcchtTsdKvlA0SRqwp
m5G7YfaK+8I2ZdkJBWpjhNBqk3tTFYamRutM84rWSPET5WRIR1VVjPew+PV8jgRz
00wPGWvWLJCoprMtBPTJsW+PVKJ+wFUCc6l6iHAjJKpGqYXp/EaDyK+dUShhHTOC
KEQ/OcwdSWv1IAC8+Gr0rZfrgW2WFAS//0KXGhRmOsWUd1hziZS0P9s8YkFAEO4J
lcel8e1okm+CPruat/ynOHg/tN6pgot/oqTkhIFN+vaWIsc5BOW31qoigre8TiUG
vdjES/iEgWOzqQ/f1HnGT9rIJFWVVzOwnA3ihZHtXvpVJ6/I6jgGtSl8ve82j4tT
1L2QUEwTeK96WRnWzst4JO/Bs8nxUvFhaOkbVPQhA+NZzSuxuZpfMFTgWL3lbW28
suvWI9U1F0TiiWVKVct8cIyThSOVmn72WcU4ouSEOmUPQqDf37H4EyTUsFDtFMpI
ptLxL19oMMTaSCXGUGIPHKXmnKUdqVwT2YRtuEbVAHZsJKzijZUfiBYqEFf8184g
OU9VLKJo7XLcC0GK8YjyF4UPlBtT8oCpH65btwBvTNcZQVopxDCNqZyYpPev5gcH
MZ2UOaKkwGkUQ+WlZXLGyJ+zVy8wzITFskfU7AzPBR0AyXYuNxeV9Aw3DvdSLr8+
zXY9LzzOoRasdB8lO7DpNh0amPimVwAqkuPiGIAJeZW0+F0HSeP+UwhZPEWpuupS
BhHZRjZa5JnYoZVIWUoXImi2vW0waIIEirsxwzwrZ88XUx3a1cQVp8S977UK1L4f
bafQcIDk17nX/6CClYeLKzgVqegkeeqr6sh9XB7WyLO5LplLrX948SNnfEV5FVxV
tUWWAwQ3uwnANh07mekJHuhce1+zlJ/r6Atje+3iYBkKQwWgnZNjxUZnvzGE/ArH
j4/RWj6Hg3bNWqVsXPo6now2r7SlR+AVUadHkdSrzWVGQa31MVMjVMpQPVCD4UrU
lswH/df+r+AyYbvLwOreWTlsDw7l3XuAMrBTxi94ZnA36ejWiR2txvjvcDY3zEj2
Us4CHvpi6wSb5TPZnp5d+ZJtALtrO9Ez1KxnmBi8V6UXrVZ1xB73UeWskIt03pDx
YHnpz5q4SXc8d0a4OZ80wifZDgz/rGV4+C6aE2IdLe8rrL4D+UVIQd3X5S+45XNx
cBO/wfl9qhkChT6Fq9VSTi5US6Lu4Hi9EuTZmSbQ+Y/SNT/2zODWSm3SjwhTQznf
NzaDyVFGhGvVvYeGqlVtQl2JrObPSpWpEXVT+NGXtE7xu2B7b18DgcMtc97+wX/d
G5JcGj7NhAdIG/NYNSF1qwO0MnxV4UiRnEarz8+Wnt2xzHIBmnnb9yRYUKkJWGOZ
Gf/MfR1np9F2Dz4GeZ+3IcWpi+x9UiFvrG/8r90D3eTe+Q0G0bZFa+hNXWdMESdS
6bd+6H8u1Q6WzS5l+y9eW/f5PVdl6MuN2aEfbOzRzRdRuuciZtLh6sDkp71s4cjr
E7DRKszAVFwrKyTfYQTsQ3gA2jEJJ2RMg3qJ3HQV9R3lU0xoSv+nbB0CmXFPMmMM
nsntol8TbSaZrKfaRHJtp03Vf+OOqLqrdqRtHVyJ0LYho//jFgdVclCva8qJ5IxC
xy3zIfRfRwX+OCxTxsYjuVfxZFecwoKWFRxmhsoK02jWfwG3yIPBvQeYhKGRjR/u
/+XVknsQWDA/a6ztJA7btcHIb/EgmwNj9iThUiwYEZV2Sw5JpjrfTod+NNF8WMVh
D055Sfzkw3LnygCYlnx8Fo3pQ0172sdtPb3kUmPd77+508twDzqc78uz2HSIo4jv
MdRC73CYtCkgIWDKNXoe2uxw1rY4pOXHObEuNCKj6rcXYcilipQMTxe5Czrx3f0D
LfX6xBYEjuDH5n/7AaN8XZEOYoQUtaMs1TgNON67KHpuGOY6EKD3gjmdFI0i2WCB
H7Sh7rJxD480tipx2t5NkMzf48vssCevv9Cs+u6saoJnGspai9UVS1jKk1P+OZaY
hiHv/Zo/XTILAMkUaEHqTPa9LhbL0YcdhdTz4jefCDoYwzGjR7h8c65YxWXOdyOl
lTSGGGZfEwoRrEjp/YobtYAnEs2m/Ir3igCrE1mjiJ6JNEKpRuUfQCZESZK3FiDa
YruHzerSdo/GWXi310V2oiqOf9fE0vAS62Q3ZWjsw0p7J6OLp1wTDDUm3dEvqmu6
k5wJHA3A9eeDDgr8KcyEykRTRj0UVzBSZsxJS+X6Fhtyp8ukF/OXvanUGIDNBz1V
fe0eaPXFV4quI1cltonHrTO0cj9dYJsBWFf9/GM6mIf5fU5GwBh549hdExiG2HpW
4IoHifArdjjhDqFeM65RX9AfNcwEXMln8gCoct5jLgO0GVP9rmgm2jn6ivQk4Nd7
Esxw97Ofu7RdJ2CEE/LGLKTGmVHf3u/emu0jZHCPvKF/F3XYCnfzn3VIjGOFUTCT
WCajBk6tmD2amyetZ4JITdTXMiyY34SGwIeBTP5nBpDi7IjAIv95J+Aj5h153DQm
Eu2ub16zsei/BhT1m9axuKJk+QeFDYm2L6UxedgAj3WJlvaY8sz34UvTrj1R9fai
ckYaD0L8OvU8snpvUumKcF28AqSiCt/guPY4iUTIkEeqLBgXHkqq0/ehGAo/R299
ZAWeW1ynJlqtyyhTyGyFeyNbfyxNAQhBJd+QDVWpkJiJbUVoyIASK48YrNRYTkp7
SEeV+MbcEZzqhkIqD/FVdvSpw9qPunTSbdgFrES3a/L5mLeUWcvfrzilBQLA2j13
p96hBP7N8Ugon+bCOsFaIm1gaiwhMAkm9ftWdq8l/khHeOdnhbsB0qcZuOyXpyJQ
08BadtOt7v85HcqYGJ9jjZb8szGKn7aEHjd+uMYJZFknDvrS+4RWBov/J516yLdG
zNigVkEdd+4tyFCpfvRdtjn1yG5CS8tPvbPP/IW5d8hjuPL56fGNDOcvP8x/wKs/
wWC8mmBiZIfMRNRTa5lPsMEQOpk2bSHCAd8Zxzu40VXFyOgKPppa63GrAqCdZ7gE
XMGBafVHfqGnCiwha8G5iHlIkTltzM49jUtFZ8ubws3o6oSgcuVtU5AEaRpODdQy
hWRF+azy5dfOmTHHngGcOsjN4R0UeHthn1rBdlvEyzvl4jzzbDbGj6TCQ8zKAgqd
t5HgTZFaVVs8CBPjpOE6FeIdFNeeHePDkYoVZVFER1dqw/15JZhIqWyFqKjclEzM
Jr90qpM47wMVyEmYsDanvPmN6u2vDGuHvtin63zwV/1nK57EqqDjbHvgjRlXPkGS
tF+/+7yAF+QAmAj8x3ixizIBy25kgWA98MtSttRiTMIIm4fBrIMGQOnTo/1sh7pR
SbATFAAQJgBY84fDhA403oZVRPNqc7adVdiIa5onWOqafcupGETO45XKNM/9P+0G
Sac+s6umyrmAyabTiVPyMVO1Lv0RB/d8NuMSg1iUxHF9n3IXIL4Ba4V4zBAmTdLE
0+4KqiO9EiWFkp00VFbvuVd1GAl6AeIOO3iGITiClZ3eY4El9PQzc/I30DGwaaik
K306RN0k9JClRwmhOfnIP1Du160oz3upDyHFSIoRY6G6eatKUTVxIJTctqgss3Li
OaeIrsoFSpX8x+6bi9ipssCe0yRt1UPsYYDlQ1pkhbytbjv91rRGuMBwMNy7E3rI
SajWiDhDwwlykePWZEbyrmoIsAtO+bo0VBey4vN4ufC07QVZmzzpWFQL/F1QniYg
93kNCcPxUdXLGaAJ9zLI7IiwChCJILyOILc3Jc17Jyo/0bCwUfpItdWgcOnU2IGE
PsuuWoY7k3wIm/Fhl8z1jzo6l3OCQroa2/xcwrJPLmxIXrtA+s88ZL3Van4C+wtO
NwmQxYSysefJ/HVD2GSo8AiwGMFoLu6YFZEw+0pCeN9X7r3Ol4AEl9CAePo40ZUP
lmNs6DwjXJvPU/eoOkaZjPqQWHSKvs8fMz1zAl+eZoD4Zr2ZcI7KXy2JpBSCb9A9
DLbqfb412hIVUG33xta1160W+TNMi5Wvi9G58TIgwjF0BiFg8KATsrw+hdxttd4S
WliZJS7WEPAzLwLI/zCNlywQgP6qyctJYyG9BzYj0VS/QO+SKDIkdUX8xtiaiHlC
jhayvEjek32hzYOwYUbFCOKvKBJKtnyyNjF3paXvCNt9bOBHnJV4VwVSSSWrdULJ
61DFMIMLg7xzrgmnQFPsf26tuqwQ+Kk16msSKSH/Qxw34OEK1k/snsK47E5anXVp
d9dDPBEyqFqg6uAXtuBHwnDTg1N4vPImMxFL/PAPFiHoClTlVO0VvSvDXvCI2Feh
CcoeWUeLG3EiRH/OqoLr4HRrFRPR8LjQBHNSKS8OM2RvE8ka9lifTbUSdBdL2GEo
18I1Y8IHzZkP9Wvwym3+jGuzoPoE/5xSZa5/Xi2v4qoD0V+1xxoY5R5IhYS7zwAw
w3yu6nyZC/i0yDyWpmvQ4WB791kLTf9UMwX4lqlmATFFFk9F1IL9dLIdzX2OtosH
YfuGD5YcLQBuwQmNVixxQIUAAORGTtbXwM9ANqsXQT+GpEiB4p86mo1y6OyKTgKS
ZvWIwvoLbDoqovndVNml0EEjkzKJuw2Aoa3wNHJeOER62qITApp5Q187ezL8J26F
hEV/3aaN3O9w/fNuu+4UVaISwg1BD9a7uCza5ksJWpEqkEtbOER102iBd2Zad4t3
Tw6AlSKLOTLA0lF75KjDkJUPswWZmtvKgwZfchh9Vbtt2mxM3pSa6JLLCwQRqjwW
mJlV+CascIthgA5hINFOHhczmtfZTQoNWIGfU8mEKTBWsxewTO9PoY0Dt0bxW5rz
nNNeryNrUTkL3NzEpa8Wifl2J2VL2/9BkvOhE3hH8IeNa6yqSMWiEsT6QrL9LRl+
pyf5wRqsL69Uh51cSIUxryE8kc0lLykwiPEBBaBvzg8vNrs/ZwDW1N1ZFzcjb1hM
JzKJZFnedZ1UdPB1CqhbQEfyAx/hJvRXf2kujN3w7gSf3yKkJx0NhTomHLjd9B/3
84m6Yw+DRF3oG1VQ8WwAqbeKMT2PzM4r9qnqYdUlget5dNC6uUW2YmzoCSgxbqzX
2yXPWpkmZjbLWj2xu2g5ddgq0A/pgB5ijdvcMnnYGiUQXQDb0QDwpQN9aTCgHWvB
g8+Ki+EQOrZtV1a70g6sRHn0s4hVh7+vCgtfmfmoaArpr2hkSWWjk8TurKX+P/Xn
iV+9MLBKRyauz2fZMmQ411+lkUTUPKrDEVacqeBSBusItXlKowbQ61E236nBztHq
PYKtMrNcYf4xbUFxa7ZK0AoynjjNujXqpZ0WPColaS8ufxOyHJx74ZogPIYyTXz0
i1+svI6L84itgbkki4mxTV0hUwWldrJDp2uDQC5ZLlTt2BMyy6e4nwPH0mZivA4Q
6yhP4aNq0G0ZQS7qNHUVckc0oac/pAqoj96sekUcWnIS/PTRCvWXmwXwMl6TL9ft
5u6zuJA/L+wheRsrVtKI4g==
`pragma protect end_protected
