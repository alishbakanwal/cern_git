-- alt_cv_gt_std_x3.vhd

-- Generated using ACDS version 16.0 211

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity alt_cv_gt_std_x3 is
	port (
		pll_powerdown           : in  std_logic_vector(0 downto 0)   := (others => '0'); --           pll_powerdown.pll_powerdown
		tx_analogreset          : in  std_logic_vector(2 downto 0)   := (others => '0'); --          tx_analogreset.tx_analogreset
		tx_digitalreset         : in  std_logic_vector(2 downto 0)   := (others => '0'); --         tx_digitalreset.tx_digitalreset
		tx_serial_data          : out std_logic_vector(2 downto 0);                      --          tx_serial_data.tx_serial_data
		ext_pll_clk             : in  std_logic_vector(2 downto 0)   := (others => '0'); --             ext_pll_clk.ext_pll_clk
		rx_analogreset          : in  std_logic_vector(2 downto 0)   := (others => '0'); --          rx_analogreset.rx_analogreset
		rx_digitalreset         : in  std_logic_vector(2 downto 0)   := (others => '0'); --         rx_digitalreset.rx_digitalreset
		rx_cdr_refclk           : in  std_logic_vector(0 downto 0)   := (others => '0'); --           rx_cdr_refclk.rx_cdr_refclk
		rx_serial_data          : in  std_logic_vector(2 downto 0)   := (others => '0'); --          rx_serial_data.rx_serial_data
		rx_is_lockedtoref       : out std_logic_vector(2 downto 0);                      --       rx_is_lockedtoref.rx_is_lockedtoref
		rx_is_lockedtodata      : out std_logic_vector(2 downto 0);                      --      rx_is_lockedtodata.rx_is_lockedtodata
		rx_seriallpbken         : in  std_logic_vector(2 downto 0)   := (others => '0'); --         rx_seriallpbken.rx_seriallpbken
		tx_std_coreclkin        : in  std_logic_vector(2 downto 0)   := (others => '0'); --        tx_std_coreclkin.tx_std_coreclkin
		rx_std_coreclkin        : in  std_logic_vector(2 downto 0)   := (others => '0'); --        rx_std_coreclkin.rx_std_coreclkin
		tx_std_clkout           : out std_logic_vector(2 downto 0);                      --           tx_std_clkout.tx_std_clkout
		rx_std_clkout           : out std_logic_vector(2 downto 0);                      --           rx_std_clkout.rx_std_clkout
		tx_std_polinv           : in  std_logic_vector(2 downto 0)   := (others => '0'); --           tx_std_polinv.tx_std_polinv
		rx_std_polinv           : in  std_logic_vector(2 downto 0)   := (others => '0'); --           rx_std_polinv.rx_std_polinv
		tx_cal_busy             : out std_logic_vector(2 downto 0);                      --             tx_cal_busy.tx_cal_busy
		rx_cal_busy             : out std_logic_vector(2 downto 0);                      --             rx_cal_busy.rx_cal_busy
		reconfig_to_xcvr        : in  std_logic_vector(209 downto 0) := (others => '0'); --        reconfig_to_xcvr.reconfig_to_xcvr
		reconfig_from_xcvr      : out std_logic_vector(137 downto 0);                    --      reconfig_from_xcvr.reconfig_from_xcvr
		tx_parallel_data        : in  std_logic_vector(119 downto 0) := (others => '0'); --        tx_parallel_data.tx_parallel_data
		unused_tx_parallel_data : in  std_logic_vector(11 downto 0)  := (others => '0'); -- unused_tx_parallel_data.unused_tx_parallel_data
		rx_parallel_data        : out std_logic_vector(119 downto 0);                    --        rx_parallel_data.rx_parallel_data
		unused_rx_parallel_data : out std_logic_vector(71 downto 0)                      -- unused_rx_parallel_data.unused_rx_parallel_data
	);
end entity alt_cv_gt_std_x3;

architecture rtl of alt_cv_gt_std_x3 is
	component altera_xcvr_native_av is
		generic (
			tx_enable                       : integer := 1;
			rx_enable                       : integer := 1;
			enable_std                      : integer := 1;
			data_path_select                : string  := "standard";
			channels                        : integer := 1;
			bonded_mode                     : string  := "non_bonded";
			data_rate                       : string  := "";
			pma_width                       : integer := 10;
			tx_pma_clk_div                  : integer := 1;
			pll_reconfig_enable             : integer := 0;
			pll_external_enable             : integer := 0;
			pll_data_rate                   : string  := "0 Mbps";
			pll_type                        : string  := "CMU";
			pma_bonding_mode                : string  := "x1";
			plls                            : integer := 1;
			pll_select                      : integer := 0;
			pll_refclk_cnt                  : integer := 1;
			pll_refclk_select               : string  := "0";
			pll_refclk_freq                 : string  := "125.0 MHz";
			pll_feedback_path               : string  := "internal";
			cdr_reconfig_enable             : integer := 0;
			cdr_refclk_cnt                  : integer := 1;
			cdr_refclk_select               : integer := 0;
			cdr_refclk_freq                 : string  := "";
			rx_ppm_detect_threshold         : string  := "1000";
			rx_clkslip_enable               : integer := 0;
			std_protocol_hint               : string  := "basic";
			std_pcs_pma_width               : integer := 10;
			std_low_latency_bypass_enable   : integer := 0;
			std_tx_pcfifo_mode              : string  := "low_latency";
			std_rx_pcfifo_mode              : string  := "low_latency";
			std_rx_byte_order_enable        : integer := 0;
			std_rx_byte_order_mode          : string  := "manual";
			std_rx_byte_order_width         : integer := 10;
			std_rx_byte_order_symbol_count  : integer := 1;
			std_rx_byte_order_pattern       : string  := "0";
			std_rx_byte_order_pad           : string  := "0";
			std_tx_byte_ser_enable          : integer := 0;
			std_rx_byte_deser_enable        : integer := 0;
			std_tx_8b10b_enable             : integer := 0;
			std_tx_8b10b_disp_ctrl_enable   : integer := 0;
			std_rx_8b10b_enable             : integer := 0;
			std_rx_rmfifo_enable            : integer := 0;
			std_rx_rmfifo_pattern_p         : string  := "00000";
			std_rx_rmfifo_pattern_n         : string  := "00000";
			std_tx_bitslip_enable           : integer := 0;
			std_rx_word_aligner_mode        : string  := "bit_slip";
			std_rx_word_aligner_pattern_len : integer := 7;
			std_rx_word_aligner_pattern     : string  := "0000000000";
			std_rx_word_aligner_rknumber    : integer := 3;
			std_rx_word_aligner_renumber    : integer := 3;
			std_rx_word_aligner_rgnumber    : integer := 3;
			std_rx_run_length_val           : integer := 31;
			std_tx_bitrev_enable            : integer := 0;
			std_rx_bitrev_enable            : integer := 0;
			std_tx_byterev_enable           : integer := 0;
			std_rx_byterev_enable           : integer := 0;
			std_tx_polinv_enable            : integer := 0;
			std_rx_polinv_enable            : integer := 0
		);
		port (
			pll_powerdown             : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- pll_powerdown
			tx_analogreset            : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- tx_analogreset
			tx_digitalreset           : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- tx_digitalreset
			tx_serial_data            : out std_logic_vector(2 downto 0);                      -- tx_serial_data
			ext_pll_clk               : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- ext_pll_clk
			rx_analogreset            : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_analogreset
			rx_digitalreset           : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_digitalreset
			rx_cdr_refclk             : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- rx_cdr_refclk
			rx_serial_data            : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_serial_data
			rx_is_lockedtoref         : out std_logic_vector(2 downto 0);                      -- rx_is_lockedtoref
			rx_is_lockedtodata        : out std_logic_vector(2 downto 0);                      -- rx_is_lockedtodata
			rx_seriallpbken           : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_seriallpbken
			tx_std_coreclkin          : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- tx_std_coreclkin
			rx_std_coreclkin          : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_std_coreclkin
			tx_std_clkout             : out std_logic_vector(2 downto 0);                      -- tx_std_clkout
			rx_std_clkout             : out std_logic_vector(2 downto 0);                      -- rx_std_clkout
			tx_std_polinv             : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- tx_std_polinv
			rx_std_polinv             : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_std_polinv
			tx_cal_busy               : out std_logic_vector(2 downto 0);                      -- tx_cal_busy
			rx_cal_busy               : out std_logic_vector(2 downto 0);                      -- rx_cal_busy
			reconfig_to_xcvr          : in  std_logic_vector(209 downto 0) := (others => 'X'); -- reconfig_to_xcvr
			reconfig_from_xcvr        : out std_logic_vector(137 downto 0);                    -- reconfig_from_xcvr
			tx_parallel_data          : in  std_logic_vector(131 downto 0) := (others => 'X'); -- unused_tx_parallel_data
			rx_parallel_data          : out std_logic_vector(191 downto 0);                    -- unused_rx_parallel_data
			tx_pll_refclk             : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- tx_pll_refclk
			tx_pma_clkout             : out std_logic_vector(2 downto 0);                      -- tx_pma_clkout
			tx_pma_parallel_data      : in  std_logic_vector(239 downto 0) := (others => 'X'); -- tx_pma_parallel_data
			pll_locked                : out std_logic_vector(0 downto 0);                      -- pll_locked
			rx_pma_clkout             : out std_logic_vector(2 downto 0);                      -- rx_pma_clkout
			rx_pma_parallel_data      : out std_logic_vector(239 downto 0);                    -- rx_pma_parallel_data
			rx_clkslip                : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_clkslip
			rx_clklow                 : out std_logic_vector(2 downto 0);                      -- rx_clklow
			rx_fref                   : out std_logic_vector(2 downto 0);                      -- rx_fref
			rx_set_locktodata         : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_set_locktodata
			rx_set_locktoref          : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_set_locktoref
			rx_signaldetect           : out std_logic_vector(2 downto 0);                      -- rx_signaldetect
			rx_std_prbs_done          : out std_logic_vector(2 downto 0);                      -- rx_std_prbs_done
			rx_std_prbs_err           : out std_logic_vector(2 downto 0);                      -- rx_std_prbs_err
			tx_std_pcfifo_full        : out std_logic_vector(2 downto 0);                      -- tx_std_pcfifo_full
			tx_std_pcfifo_empty       : out std_logic_vector(2 downto 0);                      -- tx_std_pcfifo_empty
			rx_std_pcfifo_full        : out std_logic_vector(2 downto 0);                      -- rx_std_pcfifo_full
			rx_std_pcfifo_empty       : out std_logic_vector(2 downto 0);                      -- rx_std_pcfifo_empty
			rx_std_byteorder_ena      : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_std_byteorder_ena
			rx_std_byteorder_flag     : out std_logic_vector(2 downto 0);                      -- rx_std_byteorder_flag
			rx_std_rmfifo_full        : out std_logic_vector(2 downto 0);                      -- rx_std_rmfifo_full
			rx_std_rmfifo_empty       : out std_logic_vector(2 downto 0);                      -- rx_std_rmfifo_empty
			rx_std_wa_patternalign    : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_std_wa_patternalign
			rx_std_wa_a1a2size        : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_std_wa_a1a2size
			tx_std_bitslipboundarysel : in  std_logic_vector(14 downto 0)  := (others => 'X'); -- tx_std_bitslipboundarysel
			rx_std_bitslipboundarysel : out std_logic_vector(14 downto 0);                     -- rx_std_bitslipboundarysel
			rx_std_bitslip            : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_std_bitslip
			rx_std_runlength_err      : out std_logic_vector(2 downto 0);                      -- rx_std_runlength_err
			rx_std_bitrev_ena         : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_std_bitrev_ena
			rx_std_byterev_ena        : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_std_byterev_ena
			tx_std_elecidle           : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- tx_std_elecidle
			rx_std_signaldetect       : out std_logic_vector(2 downto 0)                       -- rx_std_signaldetect
		);
	end component altera_xcvr_native_av;

	signal alt_cv_gt_std_x3_inst_rx_parallel_data : std_logic_vector(191 downto 0); -- port fragment

begin

	alt_cv_gt_std_x3_inst : component altera_xcvr_native_av
		generic map (
			tx_enable                       => 1,
			rx_enable                       => 1,
			enable_std                      => 1,
			data_path_select                => "standard",
			channels                        => 3,
			bonded_mode                     => "xN",
			data_rate                       => "4800 Mbps",
			pma_width                       => 20,
			tx_pma_clk_div                  => 1,
			pll_reconfig_enable             => 0,
			pll_external_enable             => 1,
			pll_data_rate                   => "4800 Mbps",
			pll_type                        => "CMU",
			pma_bonding_mode                => "xN",
			plls                            => 1,
			pll_select                      => 0,
			pll_refclk_cnt                  => 1,
			pll_refclk_select               => "0",
			pll_refclk_freq                 => "125.0 MHz",
			pll_feedback_path               => "internal",
			cdr_reconfig_enable             => 0,
			cdr_refclk_cnt                  => 1,
			cdr_refclk_select               => 0,
			cdr_refclk_freq                 => "120.0 MHz",
			rx_ppm_detect_threshold         => "1000",
			rx_clkslip_enable               => 0,
			std_protocol_hint               => "basic",
			std_pcs_pma_width               => 20,
			std_low_latency_bypass_enable   => 0,
			std_tx_pcfifo_mode              => "low_latency",
			std_rx_pcfifo_mode              => "low_latency",
			std_rx_byte_order_enable        => 0,
			std_rx_byte_order_mode          => "manual",
			std_rx_byte_order_width         => 10,
			std_rx_byte_order_symbol_count  => 1,
			std_rx_byte_order_pattern       => "0",
			std_rx_byte_order_pad           => "0",
			std_tx_byte_ser_enable          => 1,
			std_rx_byte_deser_enable        => 1,
			std_tx_8b10b_enable             => 0,
			std_tx_8b10b_disp_ctrl_enable   => 0,
			std_rx_8b10b_enable             => 0,
			std_rx_rmfifo_enable            => 0,
			std_rx_rmfifo_pattern_p         => "00000",
			std_rx_rmfifo_pattern_n         => "00000",
			std_tx_bitslip_enable           => 0,
			std_rx_word_aligner_mode        => "bit_slip",
			std_rx_word_aligner_pattern_len => 7,
			std_rx_word_aligner_pattern     => "0000000000",
			std_rx_word_aligner_rknumber    => 3,
			std_rx_word_aligner_renumber    => 3,
			std_rx_word_aligner_rgnumber    => 3,
			std_rx_run_length_val           => 31,
			std_tx_bitrev_enable            => 0,
			std_rx_bitrev_enable            => 0,
			std_tx_byterev_enable           => 0,
			std_rx_byterev_enable           => 0,
			std_tx_polinv_enable            => 1,
			std_rx_polinv_enable            => 1
		)
		port map (
			pll_powerdown             => pll_powerdown,                                                                                                                                                                                                                                      --      pll_powerdown.pll_powerdown
			tx_analogreset            => tx_analogreset,                                                                                                                                                                                                                                     --     tx_analogreset.tx_analogreset
			tx_digitalreset           => tx_digitalreset,                                                                                                                                                                                                                                    --    tx_digitalreset.tx_digitalreset
			tx_serial_data            => tx_serial_data,                                                                                                                                                                                                                                     --     tx_serial_data.tx_serial_data
			ext_pll_clk               => ext_pll_clk,                                                                                                                                                                                                                                        --        ext_pll_clk.ext_pll_clk
			rx_analogreset            => rx_analogreset,                                                                                                                                                                                                                                     --     rx_analogreset.rx_analogreset
			rx_digitalreset           => rx_digitalreset,                                                                                                                                                                                                                                    --    rx_digitalreset.rx_digitalreset
			rx_cdr_refclk             => rx_cdr_refclk,                                                                                                                                                                                                                                      --      rx_cdr_refclk.rx_cdr_refclk
			rx_serial_data            => rx_serial_data,                                                                                                                                                                                                                                     --     rx_serial_data.rx_serial_data
			rx_is_lockedtoref         => rx_is_lockedtoref,                                                                                                                                                                                                                                  --  rx_is_lockedtoref.rx_is_lockedtoref
			rx_is_lockedtodata        => rx_is_lockedtodata,                                                                                                                                                                                                                                 -- rx_is_lockedtodata.rx_is_lockedtodata
			rx_seriallpbken           => rx_seriallpbken,                                                                                                                                                                                                                                    --    rx_seriallpbken.rx_seriallpbken
			tx_std_coreclkin          => tx_std_coreclkin,                                                                                                                                                                                                                                   --   tx_std_coreclkin.tx_std_coreclkin
			rx_std_coreclkin          => rx_std_coreclkin,                                                                                                                                                                                                                                   --   rx_std_coreclkin.rx_std_coreclkin
			tx_std_clkout             => tx_std_clkout,                                                                                                                                                                                                                                      --      tx_std_clkout.tx_std_clkout
			rx_std_clkout             => rx_std_clkout,                                                                                                                                                                                                                                      --      rx_std_clkout.rx_std_clkout
			tx_std_polinv             => tx_std_polinv,                                                                                                                                                                                                                                      --      tx_std_polinv.tx_std_polinv
			rx_std_polinv             => rx_std_polinv,                                                                                                                                                                                                                                      --      rx_std_polinv.rx_std_polinv
			tx_cal_busy               => tx_cal_busy,                                                                                                                                                                                                                                        --        tx_cal_busy.tx_cal_busy
			rx_cal_busy               => rx_cal_busy,                                                                                                                                                                                                                                        --        rx_cal_busy.rx_cal_busy
			reconfig_to_xcvr          => reconfig_to_xcvr,                                                                                                                                                                                                                                   --   reconfig_to_xcvr.reconfig_to_xcvr
			reconfig_from_xcvr        => reconfig_from_xcvr,                                                                                                                                                                                                                                 -- reconfig_from_xcvr.reconfig_from_xcvr
			tx_parallel_data(0)       => tx_parallel_data(0),                                                                                                                                                                                                                                --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(1)       => tx_parallel_data(1),                                                                                                                                                                                                                                --                   .tx_parallel_data
			tx_parallel_data(2)       => tx_parallel_data(2),                                                                                                                                                                                                                                --                   .tx_parallel_data
			tx_parallel_data(3)       => tx_parallel_data(3),                                                                                                                                                                                                                                --                   .tx_parallel_data
			tx_parallel_data(4)       => tx_parallel_data(4),                                                                                                                                                                                                                                --                   .tx_parallel_data
			tx_parallel_data(5)       => tx_parallel_data(5),                                                                                                                                                                                                                                --                   .tx_parallel_data
			tx_parallel_data(6)       => tx_parallel_data(6),                                                                                                                                                                                                                                --                   .tx_parallel_data
			tx_parallel_data(7)       => tx_parallel_data(7),                                                                                                                                                                                                                                --                   .tx_parallel_data
			tx_parallel_data(8)       => tx_parallel_data(8),                                                                                                                                                                                                                                --                   .tx_parallel_data
			tx_parallel_data(9)       => tx_parallel_data(9),                                                                                                                                                                                                                                --                   .tx_parallel_data
			tx_parallel_data(10)      => unused_tx_parallel_data(0),                                                                                                                                                                                                                         --                   .tx_parallel_data
			tx_parallel_data(11)      => tx_parallel_data(10),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(12)      => tx_parallel_data(11),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(13)      => tx_parallel_data(12),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(14)      => tx_parallel_data(13),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(15)      => tx_parallel_data(14),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(16)      => tx_parallel_data(15),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(17)      => tx_parallel_data(16),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(18)      => tx_parallel_data(17),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(19)      => tx_parallel_data(18),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(20)      => tx_parallel_data(19),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(21)      => unused_tx_parallel_data(1),                                                                                                                                                                                                                         --                   .tx_parallel_data
			tx_parallel_data(22)      => tx_parallel_data(20),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(23)      => tx_parallel_data(21),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(24)      => tx_parallel_data(22),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(25)      => tx_parallel_data(23),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(26)      => tx_parallel_data(24),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(27)      => tx_parallel_data(25),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(28)      => tx_parallel_data(26),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(29)      => tx_parallel_data(27),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(30)      => tx_parallel_data(28),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(31)      => tx_parallel_data(29),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(32)      => unused_tx_parallel_data(2),                                                                                                                                                                                                                         --                   .tx_parallel_data
			tx_parallel_data(33)      => tx_parallel_data(30),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(34)      => tx_parallel_data(31),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(35)      => tx_parallel_data(32),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(36)      => tx_parallel_data(33),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(37)      => tx_parallel_data(34),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(38)      => tx_parallel_data(35),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(39)      => tx_parallel_data(36),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(40)      => tx_parallel_data(37),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(41)      => tx_parallel_data(38),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(42)      => tx_parallel_data(39),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(43)      => unused_tx_parallel_data(3),                                                                                                                                                                                                                         --                   .tx_parallel_data
			tx_parallel_data(44)      => tx_parallel_data(40),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(45)      => tx_parallel_data(41),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(46)      => tx_parallel_data(42),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(47)      => tx_parallel_data(43),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(48)      => tx_parallel_data(44),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(49)      => tx_parallel_data(45),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(50)      => tx_parallel_data(46),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(51)      => tx_parallel_data(47),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(52)      => tx_parallel_data(48),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(53)      => tx_parallel_data(49),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(54)      => unused_tx_parallel_data(4),                                                                                                                                                                                                                         --                   .tx_parallel_data
			tx_parallel_data(55)      => tx_parallel_data(50),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(56)      => tx_parallel_data(51),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(57)      => tx_parallel_data(52),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(58)      => tx_parallel_data(53),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(59)      => tx_parallel_data(54),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(60)      => tx_parallel_data(55),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(61)      => tx_parallel_data(56),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(62)      => tx_parallel_data(57),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(63)      => tx_parallel_data(58),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(64)      => tx_parallel_data(59),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(65)      => unused_tx_parallel_data(5),                                                                                                                                                                                                                         --                   .tx_parallel_data
			tx_parallel_data(66)      => tx_parallel_data(60),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(67)      => tx_parallel_data(61),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(68)      => tx_parallel_data(62),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(69)      => tx_parallel_data(63),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(70)      => tx_parallel_data(64),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(71)      => tx_parallel_data(65),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(72)      => tx_parallel_data(66),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(73)      => tx_parallel_data(67),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(74)      => tx_parallel_data(68),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(75)      => tx_parallel_data(69),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(76)      => unused_tx_parallel_data(6),                                                                                                                                                                                                                         --                   .tx_parallel_data
			tx_parallel_data(77)      => tx_parallel_data(70),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(78)      => tx_parallel_data(71),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(79)      => tx_parallel_data(72),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(80)      => tx_parallel_data(73),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(81)      => tx_parallel_data(74),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(82)      => tx_parallel_data(75),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(83)      => tx_parallel_data(76),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(84)      => tx_parallel_data(77),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(85)      => tx_parallel_data(78),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(86)      => tx_parallel_data(79),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(87)      => unused_tx_parallel_data(7),                                                                                                                                                                                                                         --                   .tx_parallel_data
			tx_parallel_data(88)      => tx_parallel_data(80),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(89)      => tx_parallel_data(81),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(90)      => tx_parallel_data(82),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(91)      => tx_parallel_data(83),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(92)      => tx_parallel_data(84),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(93)      => tx_parallel_data(85),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(94)      => tx_parallel_data(86),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(95)      => tx_parallel_data(87),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(96)      => tx_parallel_data(88),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(97)      => tx_parallel_data(89),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(98)      => unused_tx_parallel_data(8),                                                                                                                                                                                                                         --                   .tx_parallel_data
			tx_parallel_data(99)      => tx_parallel_data(90),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(100)     => tx_parallel_data(91),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(101)     => tx_parallel_data(92),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(102)     => tx_parallel_data(93),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(103)     => tx_parallel_data(94),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(104)     => tx_parallel_data(95),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(105)     => tx_parallel_data(96),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(106)     => tx_parallel_data(97),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(107)     => tx_parallel_data(98),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(108)     => tx_parallel_data(99),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(109)     => unused_tx_parallel_data(9),                                                                                                                                                                                                                         --                   .tx_parallel_data
			tx_parallel_data(110)     => tx_parallel_data(100),                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(111)     => tx_parallel_data(101),                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(112)     => tx_parallel_data(102),                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(113)     => tx_parallel_data(103),                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(114)     => tx_parallel_data(104),                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(115)     => tx_parallel_data(105),                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(116)     => tx_parallel_data(106),                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(117)     => tx_parallel_data(107),                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(118)     => tx_parallel_data(108),                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(119)     => tx_parallel_data(109),                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(120)     => unused_tx_parallel_data(10),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(121)     => tx_parallel_data(110),                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(122)     => tx_parallel_data(111),                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(123)     => tx_parallel_data(112),                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(124)     => tx_parallel_data(113),                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(125)     => tx_parallel_data(114),                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(126)     => tx_parallel_data(115),                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(127)     => tx_parallel_data(116),                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(128)     => tx_parallel_data(117),                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(129)     => tx_parallel_data(118),                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(130)     => tx_parallel_data(119),                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(131)     => unused_tx_parallel_data(11),                                                                                                                                                                                                                        --                   .tx_parallel_data
			rx_parallel_data(0)       => alt_cv_gt_std_x3_inst_rx_parallel_data(0),                                                                                                                                                                                                          --   rx_parallel_data.rx_parallel_data
			rx_parallel_data(1)       => alt_cv_gt_std_x3_inst_rx_parallel_data(1),                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(2)       => alt_cv_gt_std_x3_inst_rx_parallel_data(2),                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(3)       => alt_cv_gt_std_x3_inst_rx_parallel_data(3),                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(4)       => alt_cv_gt_std_x3_inst_rx_parallel_data(4),                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(5)       => alt_cv_gt_std_x3_inst_rx_parallel_data(5),                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(6)       => alt_cv_gt_std_x3_inst_rx_parallel_data(6),                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(7)       => alt_cv_gt_std_x3_inst_rx_parallel_data(7),                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(8)       => alt_cv_gt_std_x3_inst_rx_parallel_data(8),                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(9)       => alt_cv_gt_std_x3_inst_rx_parallel_data(9),                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(10)      => alt_cv_gt_std_x3_inst_rx_parallel_data(10),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(11)      => alt_cv_gt_std_x3_inst_rx_parallel_data(11),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(12)      => alt_cv_gt_std_x3_inst_rx_parallel_data(12),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(13)      => alt_cv_gt_std_x3_inst_rx_parallel_data(13),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(14)      => alt_cv_gt_std_x3_inst_rx_parallel_data(14),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(15)      => alt_cv_gt_std_x3_inst_rx_parallel_data(15),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(16)      => alt_cv_gt_std_x3_inst_rx_parallel_data(16),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(17)      => alt_cv_gt_std_x3_inst_rx_parallel_data(17),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(18)      => alt_cv_gt_std_x3_inst_rx_parallel_data(18),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(19)      => alt_cv_gt_std_x3_inst_rx_parallel_data(19),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(20)      => alt_cv_gt_std_x3_inst_rx_parallel_data(20),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(21)      => alt_cv_gt_std_x3_inst_rx_parallel_data(21),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(22)      => alt_cv_gt_std_x3_inst_rx_parallel_data(22),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(23)      => alt_cv_gt_std_x3_inst_rx_parallel_data(23),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(24)      => alt_cv_gt_std_x3_inst_rx_parallel_data(24),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(25)      => alt_cv_gt_std_x3_inst_rx_parallel_data(25),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(26)      => alt_cv_gt_std_x3_inst_rx_parallel_data(26),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(27)      => alt_cv_gt_std_x3_inst_rx_parallel_data(27),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(28)      => alt_cv_gt_std_x3_inst_rx_parallel_data(28),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(29)      => alt_cv_gt_std_x3_inst_rx_parallel_data(29),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(30)      => alt_cv_gt_std_x3_inst_rx_parallel_data(30),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(31)      => alt_cv_gt_std_x3_inst_rx_parallel_data(31),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(32)      => alt_cv_gt_std_x3_inst_rx_parallel_data(32),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(33)      => alt_cv_gt_std_x3_inst_rx_parallel_data(33),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(34)      => alt_cv_gt_std_x3_inst_rx_parallel_data(34),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(35)      => alt_cv_gt_std_x3_inst_rx_parallel_data(35),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(36)      => alt_cv_gt_std_x3_inst_rx_parallel_data(36),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(37)      => alt_cv_gt_std_x3_inst_rx_parallel_data(37),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(38)      => alt_cv_gt_std_x3_inst_rx_parallel_data(38),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(39)      => alt_cv_gt_std_x3_inst_rx_parallel_data(39),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(40)      => alt_cv_gt_std_x3_inst_rx_parallel_data(40),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(41)      => alt_cv_gt_std_x3_inst_rx_parallel_data(41),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(42)      => alt_cv_gt_std_x3_inst_rx_parallel_data(42),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(43)      => alt_cv_gt_std_x3_inst_rx_parallel_data(43),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(44)      => alt_cv_gt_std_x3_inst_rx_parallel_data(44),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(45)      => alt_cv_gt_std_x3_inst_rx_parallel_data(45),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(46)      => alt_cv_gt_std_x3_inst_rx_parallel_data(46),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(47)      => alt_cv_gt_std_x3_inst_rx_parallel_data(47),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(48)      => alt_cv_gt_std_x3_inst_rx_parallel_data(48),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(49)      => alt_cv_gt_std_x3_inst_rx_parallel_data(49),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(50)      => alt_cv_gt_std_x3_inst_rx_parallel_data(50),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(51)      => alt_cv_gt_std_x3_inst_rx_parallel_data(51),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(52)      => alt_cv_gt_std_x3_inst_rx_parallel_data(52),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(53)      => alt_cv_gt_std_x3_inst_rx_parallel_data(53),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(54)      => alt_cv_gt_std_x3_inst_rx_parallel_data(54),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(55)      => alt_cv_gt_std_x3_inst_rx_parallel_data(55),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(56)      => alt_cv_gt_std_x3_inst_rx_parallel_data(56),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(57)      => alt_cv_gt_std_x3_inst_rx_parallel_data(57),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(58)      => alt_cv_gt_std_x3_inst_rx_parallel_data(58),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(59)      => alt_cv_gt_std_x3_inst_rx_parallel_data(59),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(60)      => alt_cv_gt_std_x3_inst_rx_parallel_data(60),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(61)      => alt_cv_gt_std_x3_inst_rx_parallel_data(61),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(62)      => alt_cv_gt_std_x3_inst_rx_parallel_data(62),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(63)      => alt_cv_gt_std_x3_inst_rx_parallel_data(63),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(64)      => alt_cv_gt_std_x3_inst_rx_parallel_data(64),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(65)      => alt_cv_gt_std_x3_inst_rx_parallel_data(65),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(66)      => alt_cv_gt_std_x3_inst_rx_parallel_data(66),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(67)      => alt_cv_gt_std_x3_inst_rx_parallel_data(67),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(68)      => alt_cv_gt_std_x3_inst_rx_parallel_data(68),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(69)      => alt_cv_gt_std_x3_inst_rx_parallel_data(69),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(70)      => alt_cv_gt_std_x3_inst_rx_parallel_data(70),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(71)      => alt_cv_gt_std_x3_inst_rx_parallel_data(71),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(72)      => alt_cv_gt_std_x3_inst_rx_parallel_data(72),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(73)      => alt_cv_gt_std_x3_inst_rx_parallel_data(73),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(74)      => alt_cv_gt_std_x3_inst_rx_parallel_data(74),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(75)      => alt_cv_gt_std_x3_inst_rx_parallel_data(75),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(76)      => alt_cv_gt_std_x3_inst_rx_parallel_data(76),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(77)      => alt_cv_gt_std_x3_inst_rx_parallel_data(77),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(78)      => alt_cv_gt_std_x3_inst_rx_parallel_data(78),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(79)      => alt_cv_gt_std_x3_inst_rx_parallel_data(79),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(80)      => alt_cv_gt_std_x3_inst_rx_parallel_data(80),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(81)      => alt_cv_gt_std_x3_inst_rx_parallel_data(81),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(82)      => alt_cv_gt_std_x3_inst_rx_parallel_data(82),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(83)      => alt_cv_gt_std_x3_inst_rx_parallel_data(83),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(84)      => alt_cv_gt_std_x3_inst_rx_parallel_data(84),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(85)      => alt_cv_gt_std_x3_inst_rx_parallel_data(85),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(86)      => alt_cv_gt_std_x3_inst_rx_parallel_data(86),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(87)      => alt_cv_gt_std_x3_inst_rx_parallel_data(87),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(88)      => alt_cv_gt_std_x3_inst_rx_parallel_data(88),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(89)      => alt_cv_gt_std_x3_inst_rx_parallel_data(89),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(90)      => alt_cv_gt_std_x3_inst_rx_parallel_data(90),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(91)      => alt_cv_gt_std_x3_inst_rx_parallel_data(91),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(92)      => alt_cv_gt_std_x3_inst_rx_parallel_data(92),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(93)      => alt_cv_gt_std_x3_inst_rx_parallel_data(93),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(94)      => alt_cv_gt_std_x3_inst_rx_parallel_data(94),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(95)      => alt_cv_gt_std_x3_inst_rx_parallel_data(95),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(96)      => alt_cv_gt_std_x3_inst_rx_parallel_data(96),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(97)      => alt_cv_gt_std_x3_inst_rx_parallel_data(97),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(98)      => alt_cv_gt_std_x3_inst_rx_parallel_data(98),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(99)      => alt_cv_gt_std_x3_inst_rx_parallel_data(99),                                                                                                                                                                                                         --                   .rx_parallel_data
			rx_parallel_data(100)     => alt_cv_gt_std_x3_inst_rx_parallel_data(100),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(101)     => alt_cv_gt_std_x3_inst_rx_parallel_data(101),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(102)     => alt_cv_gt_std_x3_inst_rx_parallel_data(102),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(103)     => alt_cv_gt_std_x3_inst_rx_parallel_data(103),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(104)     => alt_cv_gt_std_x3_inst_rx_parallel_data(104),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(105)     => alt_cv_gt_std_x3_inst_rx_parallel_data(105),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(106)     => alt_cv_gt_std_x3_inst_rx_parallel_data(106),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(107)     => alt_cv_gt_std_x3_inst_rx_parallel_data(107),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(108)     => alt_cv_gt_std_x3_inst_rx_parallel_data(108),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(109)     => alt_cv_gt_std_x3_inst_rx_parallel_data(109),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(110)     => alt_cv_gt_std_x3_inst_rx_parallel_data(110),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(111)     => alt_cv_gt_std_x3_inst_rx_parallel_data(111),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(112)     => alt_cv_gt_std_x3_inst_rx_parallel_data(112),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(113)     => alt_cv_gt_std_x3_inst_rx_parallel_data(113),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(114)     => alt_cv_gt_std_x3_inst_rx_parallel_data(114),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(115)     => alt_cv_gt_std_x3_inst_rx_parallel_data(115),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(116)     => alt_cv_gt_std_x3_inst_rx_parallel_data(116),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(117)     => alt_cv_gt_std_x3_inst_rx_parallel_data(117),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(118)     => alt_cv_gt_std_x3_inst_rx_parallel_data(118),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(119)     => alt_cv_gt_std_x3_inst_rx_parallel_data(119),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(120)     => alt_cv_gt_std_x3_inst_rx_parallel_data(120),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(121)     => alt_cv_gt_std_x3_inst_rx_parallel_data(121),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(122)     => alt_cv_gt_std_x3_inst_rx_parallel_data(122),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(123)     => alt_cv_gt_std_x3_inst_rx_parallel_data(123),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(124)     => alt_cv_gt_std_x3_inst_rx_parallel_data(124),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(125)     => alt_cv_gt_std_x3_inst_rx_parallel_data(125),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(126)     => alt_cv_gt_std_x3_inst_rx_parallel_data(126),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(127)     => alt_cv_gt_std_x3_inst_rx_parallel_data(127),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(128)     => alt_cv_gt_std_x3_inst_rx_parallel_data(128),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(129)     => alt_cv_gt_std_x3_inst_rx_parallel_data(129),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(130)     => alt_cv_gt_std_x3_inst_rx_parallel_data(130),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(131)     => alt_cv_gt_std_x3_inst_rx_parallel_data(131),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(132)     => alt_cv_gt_std_x3_inst_rx_parallel_data(132),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(133)     => alt_cv_gt_std_x3_inst_rx_parallel_data(133),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(134)     => alt_cv_gt_std_x3_inst_rx_parallel_data(134),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(135)     => alt_cv_gt_std_x3_inst_rx_parallel_data(135),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(136)     => alt_cv_gt_std_x3_inst_rx_parallel_data(136),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(137)     => alt_cv_gt_std_x3_inst_rx_parallel_data(137),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(138)     => alt_cv_gt_std_x3_inst_rx_parallel_data(138),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(139)     => alt_cv_gt_std_x3_inst_rx_parallel_data(139),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(140)     => alt_cv_gt_std_x3_inst_rx_parallel_data(140),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(141)     => alt_cv_gt_std_x3_inst_rx_parallel_data(141),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(142)     => alt_cv_gt_std_x3_inst_rx_parallel_data(142),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(143)     => alt_cv_gt_std_x3_inst_rx_parallel_data(143),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(144)     => alt_cv_gt_std_x3_inst_rx_parallel_data(144),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(145)     => alt_cv_gt_std_x3_inst_rx_parallel_data(145),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(146)     => alt_cv_gt_std_x3_inst_rx_parallel_data(146),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(147)     => alt_cv_gt_std_x3_inst_rx_parallel_data(147),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(148)     => alt_cv_gt_std_x3_inst_rx_parallel_data(148),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(149)     => alt_cv_gt_std_x3_inst_rx_parallel_data(149),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(150)     => alt_cv_gt_std_x3_inst_rx_parallel_data(150),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(151)     => alt_cv_gt_std_x3_inst_rx_parallel_data(151),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(152)     => alt_cv_gt_std_x3_inst_rx_parallel_data(152),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(153)     => alt_cv_gt_std_x3_inst_rx_parallel_data(153),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(154)     => alt_cv_gt_std_x3_inst_rx_parallel_data(154),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(155)     => alt_cv_gt_std_x3_inst_rx_parallel_data(155),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(156)     => alt_cv_gt_std_x3_inst_rx_parallel_data(156),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(157)     => alt_cv_gt_std_x3_inst_rx_parallel_data(157),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(158)     => alt_cv_gt_std_x3_inst_rx_parallel_data(158),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(159)     => alt_cv_gt_std_x3_inst_rx_parallel_data(159),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(160)     => alt_cv_gt_std_x3_inst_rx_parallel_data(160),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(161)     => alt_cv_gt_std_x3_inst_rx_parallel_data(161),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(162)     => alt_cv_gt_std_x3_inst_rx_parallel_data(162),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(163)     => alt_cv_gt_std_x3_inst_rx_parallel_data(163),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(164)     => alt_cv_gt_std_x3_inst_rx_parallel_data(164),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(165)     => alt_cv_gt_std_x3_inst_rx_parallel_data(165),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(166)     => alt_cv_gt_std_x3_inst_rx_parallel_data(166),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(167)     => alt_cv_gt_std_x3_inst_rx_parallel_data(167),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(168)     => alt_cv_gt_std_x3_inst_rx_parallel_data(168),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(169)     => alt_cv_gt_std_x3_inst_rx_parallel_data(169),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(170)     => alt_cv_gt_std_x3_inst_rx_parallel_data(170),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(171)     => alt_cv_gt_std_x3_inst_rx_parallel_data(171),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(172)     => alt_cv_gt_std_x3_inst_rx_parallel_data(172),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(173)     => alt_cv_gt_std_x3_inst_rx_parallel_data(173),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(174)     => alt_cv_gt_std_x3_inst_rx_parallel_data(174),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(175)     => alt_cv_gt_std_x3_inst_rx_parallel_data(175),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(176)     => alt_cv_gt_std_x3_inst_rx_parallel_data(176),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(177)     => alt_cv_gt_std_x3_inst_rx_parallel_data(177),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(178)     => alt_cv_gt_std_x3_inst_rx_parallel_data(178),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(179)     => alt_cv_gt_std_x3_inst_rx_parallel_data(179),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(180)     => alt_cv_gt_std_x3_inst_rx_parallel_data(180),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(181)     => alt_cv_gt_std_x3_inst_rx_parallel_data(181),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(182)     => alt_cv_gt_std_x3_inst_rx_parallel_data(182),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(183)     => alt_cv_gt_std_x3_inst_rx_parallel_data(183),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(184)     => alt_cv_gt_std_x3_inst_rx_parallel_data(184),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(185)     => alt_cv_gt_std_x3_inst_rx_parallel_data(185),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(186)     => alt_cv_gt_std_x3_inst_rx_parallel_data(186),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(187)     => alt_cv_gt_std_x3_inst_rx_parallel_data(187),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(188)     => alt_cv_gt_std_x3_inst_rx_parallel_data(188),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(189)     => alt_cv_gt_std_x3_inst_rx_parallel_data(189),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(190)     => alt_cv_gt_std_x3_inst_rx_parallel_data(190),                                                                                                                                                                                                        --                   .rx_parallel_data
			rx_parallel_data(191)     => alt_cv_gt_std_x3_inst_rx_parallel_data(191),                                                                                                                                                                                                        --                   .rx_parallel_data
			tx_pll_refclk             => "0",                                                                                                                                                                                                                                                --        (terminated)
			tx_pma_clkout             => open,                                                                                                                                                                                                                                               --        (terminated)
			tx_pma_parallel_data      => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", --        (terminated)
			pll_locked                => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_pma_clkout             => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_pma_parallel_data      => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_clkslip                => "000",                                                                                                                                                                                                                                              --        (terminated)
			rx_clklow                 => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_fref                   => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_set_locktodata         => "000",                                                                                                                                                                                                                                              --        (terminated)
			rx_set_locktoref          => "000",                                                                                                                                                                                                                                              --        (terminated)
			rx_signaldetect           => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_std_prbs_done          => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_std_prbs_err           => open,                                                                                                                                                                                                                                               --        (terminated)
			tx_std_pcfifo_full        => open,                                                                                                                                                                                                                                               --        (terminated)
			tx_std_pcfifo_empty       => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_std_pcfifo_full        => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_std_pcfifo_empty       => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_std_byteorder_ena      => "000",                                                                                                                                                                                                                                              --        (terminated)
			rx_std_byteorder_flag     => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_std_rmfifo_full        => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_std_rmfifo_empty       => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_std_wa_patternalign    => "000",                                                                                                                                                                                                                                              --        (terminated)
			rx_std_wa_a1a2size        => "000",                                                                                                                                                                                                                                              --        (terminated)
			tx_std_bitslipboundarysel => "000000000000000",                                                                                                                                                                                                                                  --        (terminated)
			rx_std_bitslipboundarysel => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_std_bitslip            => "000",                                                                                                                                                                                                                                              --        (terminated)
			rx_std_runlength_err      => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_std_bitrev_ena         => "000",                                                                                                                                                                                                                                              --        (terminated)
			rx_std_byterev_ena        => "000",                                                                                                                                                                                                                                              --        (terminated)
			tx_std_elecidle           => "000",                                                                                                                                                                                                                                              --        (terminated)
			rx_std_signaldetect       => open                                                                                                                                                                                                                                                --        (terminated)
		);

	rx_parallel_data <= alt_cv_gt_std_x3_inst_rx_parallel_data(185) & alt_cv_gt_std_x3_inst_rx_parallel_data(184) & alt_cv_gt_std_x3_inst_rx_parallel_data(183) & alt_cv_gt_std_x3_inst_rx_parallel_data(182) & alt_cv_gt_std_x3_inst_rx_parallel_data(181) & alt_cv_gt_std_x3_inst_rx_parallel_data(180) & alt_cv_gt_std_x3_inst_rx_parallel_data(179) & alt_cv_gt_std_x3_inst_rx_parallel_data(178) & alt_cv_gt_std_x3_inst_rx_parallel_data(177) & alt_cv_gt_std_x3_inst_rx_parallel_data(176) & alt_cv_gt_std_x3_inst_rx_parallel_data(169) & alt_cv_gt_std_x3_inst_rx_parallel_data(168) & alt_cv_gt_std_x3_inst_rx_parallel_data(167) & alt_cv_gt_std_x3_inst_rx_parallel_data(166) & alt_cv_gt_std_x3_inst_rx_parallel_data(165) & alt_cv_gt_std_x3_inst_rx_parallel_data(164) & alt_cv_gt_std_x3_inst_rx_parallel_data(163) & alt_cv_gt_std_x3_inst_rx_parallel_data(162) & alt_cv_gt_std_x3_inst_rx_parallel_data(161) & alt_cv_gt_std_x3_inst_rx_parallel_data(160) & alt_cv_gt_std_x3_inst_rx_parallel_data(153) & alt_cv_gt_std_x3_inst_rx_parallel_data(152) & alt_cv_gt_std_x3_inst_rx_parallel_data(151) & alt_cv_gt_std_x3_inst_rx_parallel_data(150) & alt_cv_gt_std_x3_inst_rx_parallel_data(149) & alt_cv_gt_std_x3_inst_rx_parallel_data(148) & alt_cv_gt_std_x3_inst_rx_parallel_data(147) & alt_cv_gt_std_x3_inst_rx_parallel_data(146) & alt_cv_gt_std_x3_inst_rx_parallel_data(145) & alt_cv_gt_std_x3_inst_rx_parallel_data(144) & alt_cv_gt_std_x3_inst_rx_parallel_data(137) & alt_cv_gt_std_x3_inst_rx_parallel_data(136) & alt_cv_gt_std_x3_inst_rx_parallel_data(135) & alt_cv_gt_std_x3_inst_rx_parallel_data(134) & alt_cv_gt_std_x3_inst_rx_parallel_data(133) & alt_cv_gt_std_x3_inst_rx_parallel_data(132) & alt_cv_gt_std_x3_inst_rx_parallel_data(131) & alt_cv_gt_std_x3_inst_rx_parallel_data(130) & alt_cv_gt_std_x3_inst_rx_parallel_data(129) & alt_cv_gt_std_x3_inst_rx_parallel_data(128) & alt_cv_gt_std_x3_inst_rx_parallel_data(121) & alt_cv_gt_std_x3_inst_rx_parallel_data(120) & alt_cv_gt_std_x3_inst_rx_parallel_data(119) & alt_cv_gt_std_x3_inst_rx_parallel_data(118) & alt_cv_gt_std_x3_inst_rx_parallel_data(117) & alt_cv_gt_std_x3_inst_rx_parallel_data(116) & alt_cv_gt_std_x3_inst_rx_parallel_data(115) & alt_cv_gt_std_x3_inst_rx_parallel_data(114) & alt_cv_gt_std_x3_inst_rx_parallel_data(113) & alt_cv_gt_std_x3_inst_rx_parallel_data(112) & alt_cv_gt_std_x3_inst_rx_parallel_data(105) & alt_cv_gt_std_x3_inst_rx_parallel_data(104) & alt_cv_gt_std_x3_inst_rx_parallel_data(103) & alt_cv_gt_std_x3_inst_rx_parallel_data(102) & alt_cv_gt_std_x3_inst_rx_parallel_data(101) & alt_cv_gt_std_x3_inst_rx_parallel_data(100) & alt_cv_gt_std_x3_inst_rx_parallel_data(99) & alt_cv_gt_std_x3_inst_rx_parallel_data(98) & alt_cv_gt_std_x3_inst_rx_parallel_data(97) & alt_cv_gt_std_x3_inst_rx_parallel_data(96) & alt_cv_gt_std_x3_inst_rx_parallel_data(89) & alt_cv_gt_std_x3_inst_rx_parallel_data(88) & alt_cv_gt_std_x3_inst_rx_parallel_data(87) & alt_cv_gt_std_x3_inst_rx_parallel_data(86) & alt_cv_gt_std_x3_inst_rx_parallel_data(85) & alt_cv_gt_std_x3_inst_rx_parallel_data(84) & alt_cv_gt_std_x3_inst_rx_parallel_data(83) & alt_cv_gt_std_x3_inst_rx_parallel_data(82) & alt_cv_gt_std_x3_inst_rx_parallel_data(81) & alt_cv_gt_std_x3_inst_rx_parallel_data(80) & alt_cv_gt_std_x3_inst_rx_parallel_data(73) & alt_cv_gt_std_x3_inst_rx_parallel_data(72) & alt_cv_gt_std_x3_inst_rx_parallel_data(71) & alt_cv_gt_std_x3_inst_rx_parallel_data(70) & alt_cv_gt_std_x3_inst_rx_parallel_data(69) & alt_cv_gt_std_x3_inst_rx_parallel_data(68) & alt_cv_gt_std_x3_inst_rx_parallel_data(67) & alt_cv_gt_std_x3_inst_rx_parallel_data(66) & alt_cv_gt_std_x3_inst_rx_parallel_data(65) & alt_cv_gt_std_x3_inst_rx_parallel_data(64) & alt_cv_gt_std_x3_inst_rx_parallel_data(57) & alt_cv_gt_std_x3_inst_rx_parallel_data(56) & alt_cv_gt_std_x3_inst_rx_parallel_data(55) & alt_cv_gt_std_x3_inst_rx_parallel_data(54) & alt_cv_gt_std_x3_inst_rx_parallel_data(53) & alt_cv_gt_std_x3_inst_rx_parallel_data(52) & alt_cv_gt_std_x3_inst_rx_parallel_data(51) & alt_cv_gt_std_x3_inst_rx_parallel_data(50) & alt_cv_gt_std_x3_inst_rx_parallel_data(49) & alt_cv_gt_std_x3_inst_rx_parallel_data(48) & alt_cv_gt_std_x3_inst_rx_parallel_data(41) & alt_cv_gt_std_x3_inst_rx_parallel_data(40) & alt_cv_gt_std_x3_inst_rx_parallel_data(39) & alt_cv_gt_std_x3_inst_rx_parallel_data(38) & alt_cv_gt_std_x3_inst_rx_parallel_data(37) & alt_cv_gt_std_x3_inst_rx_parallel_data(36) & alt_cv_gt_std_x3_inst_rx_parallel_data(35) & alt_cv_gt_std_x3_inst_rx_parallel_data(34) & alt_cv_gt_std_x3_inst_rx_parallel_data(33) & alt_cv_gt_std_x3_inst_rx_parallel_data(32) & alt_cv_gt_std_x3_inst_rx_parallel_data(25) & alt_cv_gt_std_x3_inst_rx_parallel_data(24) & alt_cv_gt_std_x3_inst_rx_parallel_data(23) & alt_cv_gt_std_x3_inst_rx_parallel_data(22) & alt_cv_gt_std_x3_inst_rx_parallel_data(21) & alt_cv_gt_std_x3_inst_rx_parallel_data(20) & alt_cv_gt_std_x3_inst_rx_parallel_data(19) & alt_cv_gt_std_x3_inst_rx_parallel_data(18) & alt_cv_gt_std_x3_inst_rx_parallel_data(17) & alt_cv_gt_std_x3_inst_rx_parallel_data(16) & alt_cv_gt_std_x3_inst_rx_parallel_data(9) & alt_cv_gt_std_x3_inst_rx_parallel_data(8) & alt_cv_gt_std_x3_inst_rx_parallel_data(7) & alt_cv_gt_std_x3_inst_rx_parallel_data(6) & alt_cv_gt_std_x3_inst_rx_parallel_data(5) & alt_cv_gt_std_x3_inst_rx_parallel_data(4) & alt_cv_gt_std_x3_inst_rx_parallel_data(3) & alt_cv_gt_std_x3_inst_rx_parallel_data(2) & alt_cv_gt_std_x3_inst_rx_parallel_data(1) & alt_cv_gt_std_x3_inst_rx_parallel_data(0);

	unused_rx_parallel_data <= alt_cv_gt_std_x3_inst_rx_parallel_data(191) & alt_cv_gt_std_x3_inst_rx_parallel_data(190) & alt_cv_gt_std_x3_inst_rx_parallel_data(189) & alt_cv_gt_std_x3_inst_rx_parallel_data(188) & alt_cv_gt_std_x3_inst_rx_parallel_data(187) & alt_cv_gt_std_x3_inst_rx_parallel_data(186) & alt_cv_gt_std_x3_inst_rx_parallel_data(175) & alt_cv_gt_std_x3_inst_rx_parallel_data(174) & alt_cv_gt_std_x3_inst_rx_parallel_data(173) & alt_cv_gt_std_x3_inst_rx_parallel_data(172) & alt_cv_gt_std_x3_inst_rx_parallel_data(171) & alt_cv_gt_std_x3_inst_rx_parallel_data(170) & alt_cv_gt_std_x3_inst_rx_parallel_data(159) & alt_cv_gt_std_x3_inst_rx_parallel_data(158) & alt_cv_gt_std_x3_inst_rx_parallel_data(157) & alt_cv_gt_std_x3_inst_rx_parallel_data(156) & alt_cv_gt_std_x3_inst_rx_parallel_data(155) & alt_cv_gt_std_x3_inst_rx_parallel_data(154) & alt_cv_gt_std_x3_inst_rx_parallel_data(143) & alt_cv_gt_std_x3_inst_rx_parallel_data(142) & alt_cv_gt_std_x3_inst_rx_parallel_data(141) & alt_cv_gt_std_x3_inst_rx_parallel_data(140) & alt_cv_gt_std_x3_inst_rx_parallel_data(139) & alt_cv_gt_std_x3_inst_rx_parallel_data(138) & alt_cv_gt_std_x3_inst_rx_parallel_data(127) & alt_cv_gt_std_x3_inst_rx_parallel_data(126) & alt_cv_gt_std_x3_inst_rx_parallel_data(125) & alt_cv_gt_std_x3_inst_rx_parallel_data(124) & alt_cv_gt_std_x3_inst_rx_parallel_data(123) & alt_cv_gt_std_x3_inst_rx_parallel_data(122) & alt_cv_gt_std_x3_inst_rx_parallel_data(111) & alt_cv_gt_std_x3_inst_rx_parallel_data(110) & alt_cv_gt_std_x3_inst_rx_parallel_data(109) & alt_cv_gt_std_x3_inst_rx_parallel_data(108) & alt_cv_gt_std_x3_inst_rx_parallel_data(107) & alt_cv_gt_std_x3_inst_rx_parallel_data(106) & alt_cv_gt_std_x3_inst_rx_parallel_data(95) & alt_cv_gt_std_x3_inst_rx_parallel_data(94) & alt_cv_gt_std_x3_inst_rx_parallel_data(93) & alt_cv_gt_std_x3_inst_rx_parallel_data(92) & alt_cv_gt_std_x3_inst_rx_parallel_data(91) & alt_cv_gt_std_x3_inst_rx_parallel_data(90) & alt_cv_gt_std_x3_inst_rx_parallel_data(79) & alt_cv_gt_std_x3_inst_rx_parallel_data(78) & alt_cv_gt_std_x3_inst_rx_parallel_data(77) & alt_cv_gt_std_x3_inst_rx_parallel_data(76) & alt_cv_gt_std_x3_inst_rx_parallel_data(75) & alt_cv_gt_std_x3_inst_rx_parallel_data(74) & alt_cv_gt_std_x3_inst_rx_parallel_data(63) & alt_cv_gt_std_x3_inst_rx_parallel_data(62) & alt_cv_gt_std_x3_inst_rx_parallel_data(61) & alt_cv_gt_std_x3_inst_rx_parallel_data(60) & alt_cv_gt_std_x3_inst_rx_parallel_data(59) & alt_cv_gt_std_x3_inst_rx_parallel_data(58) & alt_cv_gt_std_x3_inst_rx_parallel_data(47) & alt_cv_gt_std_x3_inst_rx_parallel_data(46) & alt_cv_gt_std_x3_inst_rx_parallel_data(45) & alt_cv_gt_std_x3_inst_rx_parallel_data(44) & alt_cv_gt_std_x3_inst_rx_parallel_data(43) & alt_cv_gt_std_x3_inst_rx_parallel_data(42) & alt_cv_gt_std_x3_inst_rx_parallel_data(31) & alt_cv_gt_std_x3_inst_rx_parallel_data(30) & alt_cv_gt_std_x3_inst_rx_parallel_data(29) & alt_cv_gt_std_x3_inst_rx_parallel_data(28) & alt_cv_gt_std_x3_inst_rx_parallel_data(27) & alt_cv_gt_std_x3_inst_rx_parallel_data(26) & alt_cv_gt_std_x3_inst_rx_parallel_data(15) & alt_cv_gt_std_x3_inst_rx_parallel_data(14) & alt_cv_gt_std_x3_inst_rx_parallel_data(13) & alt_cv_gt_std_x3_inst_rx_parallel_data(12) & alt_cv_gt_std_x3_inst_rx_parallel_data(11) & alt_cv_gt_std_x3_inst_rx_parallel_data(10);

end architecture rtl; -- of alt_cv_gt_std_x3
