// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:10 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nDM8yY8qPp1EhXuT+jRJCSuC3w2kB3EUndXDRHQ/u7L2CKCDtr5rtWk5yVHYotCM
SjL4JvCZRCvlFI4CKK3FLlsGnji15vWmaYBqexM8Z2ENP3jK6a1a5EPs/iB5Vomh
NKW1SOzqY8IAPABhtGULzauK+fYt2pMw1KpkZuGiiB0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 125472)
7G3w5Jbti6tBeO6p/trvGpNBaDPSEU2n64c1rK3gEledaBMD8vAvH6tCMj2YSz0u
scjQo2j+s0Vo8Ap3FXk5Tg28Rpw3KypXm/7WjQNkUT3dswstGPOuFUOsgpyHmcPa
MzRvoZQidmpjbnlV7U3NTesBKjdow/XhbZyrO4/POMdjH722HZOLGc0sxHWlYm8+
KELVLFsjedjAdtVbuk14Us6Mbiq4tqoF1ZG9GTVvYi9q8oQ+kXYExxI58+WzppV4
3VDat3p18NydFfo6UsoBKuYGNWrCkhFCQRoErYox2Ep1Ekbk9aAX+kLcm4vhcRth
o376WpOjVYUC2LFVjYGGx9MDaLBqs+VdaYmu/MRPGVr0W+LDTkAdeN7QCUfNiN7T
uoLwCzL7UaagdK5fxy24INOyC0MUyL8adTTqi/Y6KXkmgImLtEfh1/ZNjj4h4xh2
PYdfPgplF6mEWIHRColngx+xhYvo79L0OValvZeF3yvm4mn1nWS6LcwOQSJKY7Re
rlO0mFxMIMtE2HnwrfJh5zLEcvCf97WYYGOtXB9WVSYruhhGP5gDF0R9s6U9EwcQ
3sx5Q2IIcAj3t0cIfF1uSNnBCM0Zwci81wo7b+5rm3TVphtCg5x6onHoZo5DGeLg
GA13bpG+7Ylf0OLfaSU8Hd5XHXTwhW4TMOGjQxlj2f+b9MJ+++Q19XU79aBlze8R
10telUu02qAdIkm9k/ri7JNR8PSP/5J/QAae8sna/1GTNpP/pzv49YcTZ6j1JTUu
PzcMHlzfTm5jQ8Hn+0fBoyq3LNNbjy8v7douQbPa4BixYCxqcZ5uDBcDPEVRqECe
/Y5xmdTKHdryur8EZS0+chlxWtS9vFgFpat19Z2i5BvMLtfWYN8lDQa6bVX1UTc2
xbQSUInmPao/QODvBIu8QityHb8UlwgTLwZMaD94tDKVnNh5hieE1kJ6dUPOLxBo
HSlvy+strK9jZ66ewYuE3l/IOg26OVcbnw53K2O/pAJ0ufIkomtcJeEa9vG4wSU5
G/JgEpVYjoRUdlvUnh8O5E74KRujImm6CYLl+knW6Jb5HJTgB4t3f9Cf83ZeD+tc
PBYVDzwgtd1CY70a5rVT4xVwwiooEk4kmDH6xxmnU4hMJ78orwnAoyrZId93nPgX
hQMVEsPd5PQpvz2jO9WTXiejvDnHZGWMlCCQ7q30vTOc+10q2yqmK8M3mhnD2PXc
ECi8HHbyrING6PfK5Vke7UroKxgoIQ6DBZGA9ru8bV9FWxxkYm0XyPOHyxOk90lM
YIdBKMvA7i2FnmhhC+Jlxstp/dNEs7nXAhI/jpndGwBRgmhE3+t7esHDEuGxMJRs
Vr92WSexUICeuvyBW8fNgGdtm+5CbM60baVNXlFosMjLK1D4N8RO/rUuXi0dqlGj
H9oTw1cIDQawktFuHvrngGqwPoEb4CthU0x25+87365tkywnlAO+OvtOPmpx/IDg
HI7OTHsjqh72RSvwQkrhbkiwCSp/dksB4NBgAg4QimwCUyG7ZTrImT+Cm18elH/Z
Fhnu+VjyYJbgsYCDRVgdVC+pCjha3wkjG9KUmlZU34t1TMLXVEikEhIPYYh/oESr
q6lfLBKfWijwIeifRYaDXXNn7GMCnTAEsCPKvIoK8akyWkQcra9ZnR2g89DSPAH8
sWjkUOEGbqS1qkdaYEdjg2w/fWSoVASpCEqOhKL+uSNOulqeVHxTNjWyhW9YjpYF
Q2IwbPkp4JosboweIRd9lGg9pnpNMFqkKryb50Bu/UWbaiZcMKJmie6ccrfaaVWA
YCcc8wJ8UMpnpS06wVnjaNUmwF0Y/bYJx0xwTzmzfUAzRVqaDBvqfvFX4Su+PkSH
RbcLxOe2s1BgilBgVuJlfVFuy2Jpls6J7a35QcA8GxWBUY/Pz/HNPRRVYEomeBSx
3Jb5aJK7AjkMS5v0sCfzK/ZctvnzmcOanK1UcLKkNCZCFWpgqfvxc2FTMLortR1m
JwrWShxkha5MFQWH9u98DUIrWBTTygsoDAbUamPd1bQ7aEx4VFKzMLOQJC+HQrJE
e/3Buo45n1MxNsqK8wx/dITsnkkXhDLWE0/HsdUxHhSV7Bg1pZ53tewDFf489AlF
/qV1GGLrZUfSnvoKcypqFsVbzpCvZstF8H/wUSy+nGYY1WCDlE0blP4PRqVWTlxz
z0rCPTRRq7Nq7SV7B89jat0CFSTsJze67ZLdZJglOg0U4xr50HgMFMt29/9IWe4H
/6jBdYzEWzyANProX3YQBAmlPFrYMr5v8wBJJ2+9jJ/JUwFuICwAQ2/Ykyhm8WVj
OvpetCD+4iIXo1pD62+qmbZtJywKz9X3bphmBNmCrXaVknKM4hQXnqGduspq4LB6
JdUPHhUl9LZv0eED3vMoYhPrGw54YnuomroBh7WiHpiewZ1BDKi6nttKh+QLlu+j
UJFxNKv8zIbvLWxCrzNRGnNRIfBhu/bObLoY0qNsrycMYOlHAOGRQXKTCWIQOnXf
b+TzLadd68uD3zTdGt+vZuuanbDVNVyudvxJ6xKNwbbTFxpcRoEw5KHfI69KT53w
+zpFOzra/9Lh0luaHKkK6vTE+5V1auYqFh6RnAi0CStdVgez0GnfrOEauhceOKCs
ajaMYAisaqNViY8xNGIcmT+UIBvg6Mra4dmGK5bK5A9/uxXUx0EY/kO0CiAy7QIe
R/rlvAY57zyQHJRWIOUj8FXtoSYZLY0O7HDIMfIbGmorq9RBaMkzBU+AHMITpvAD
ZA4++2+SJ1cHEDofDC4pWPA8YrMx5rtH9mqfnzTdXMijtNb6MN784gOnBmBpB0E2
kc/B/9li5bJLVY8TGqB5Tw7LQ5k/UbFx8niqkhmGTTHy4EqEAfaIV8mu3oIKmznK
bPdGwVoR95X4XmuHRXz/+jP3NhwWT3O6VB8OwIaqfr74G1iZoTPvL7hK/50ZHYG0
YMHbInAHM97v7GYVR4TY2StX0UdF817vK4dVIrSnTfQ+DRSUwyeApAHOXqGGjTgc
fSn292RYG+nZbZWd5/0h1SfUpXn4fMq0HZA/btpdoDYwICwD6ZtKKcIMnFKGrxGd
X29T1MJMV3l5uihpSvKVCnRp/5z4pBzilW2oYUOm0MlSChPUEl4CsSr/OUqi5c7/
wj2hPhiNLaOHL8LaFGidJmCiyfMxiVI/5yJVwTnitiNUj1sKZL92kUWX90aVwHzg
VmMLzwPEIxMuBaKJFb7NrOVIbwFM0A6L2UBvDLVLZuLWWbCnUTop5/n/yK2fHuKi
ajIvTSDvuW8G/5Ui5fuK0QbVjdi6kKL7EJtpPH7XhyMQ1X/PXdD2G8IkxjNtBGjM
Qn2f2RUpPF7gFL8PQ+1FZ2rwPpOQUQuzcRRauNxjwt2nLnvjsnkR00MJpaytT5pI
6tBQ8KxeS2X9qBwnxAKEaUnzOKkGHugGz8VN6qd1HIihkD39a7TeMBE5F1z5i8Xf
T82C0FUzzMf7NHvmqgHFAdueUsF4M4gce0l/1huUeWkxfYMM/r1de+IUM5vesI8F
t6m8qKYZFd6KG7dAShQsEM6fpRtklMjT1VlHTWUSqjOR9RDfiN5puEDcNyYIizhw
8bqY6kaov8ARzdHYwB5GecmtmkLKYSiXRFijYjGEzvkJ8qKdT164QcU0ysaxXipq
fOJDjuSUeVg/vIr31gIXNa/N0W/SLs8cFrgnIh90tJ9sX+ozmB/+A6sCyGHcCgPY
kjBSA3y/qkbJo4iQYOkpmzTvigtsq3QgFSUpuggvWaCPtt1G3CLsGyvWknCJnHiK
bH3P4yQRM00svt5QMk+YkqkUQYFSEnekG/CGwA1ZltBat5O56j84O+/a/Vw1qyAp
JHzGWGWrMEXBT7w4xT72T7Cy7U0pehEJLCCTUO4MtX7K8dmEaGWs4eOYDkwjVPvh
Seqvnmd/4MnC92iHOEbEP5CYY75VNA6RrubyyiGFp1aqG9sB90jjzS985guHjOGb
z2nc9oFSjlhMQSTHZNzkwQbSkK6mq6gS8lnb+0Wov1EvwcSLc4MvLjXQSxmfQzei
BTU77A3qPqgg/1iI76idbS3dlgKn7m+F7KGvWuFMP+vhWdbKWd+2e+dlx6sZmgzC
UpNUPNb+9mWTrc9gwzHlv977YFCptcfR77H4aSO6BT7kxs0w63stPF2Rr2b2Euw/
vmyZ1Q3xueKdIf/5plouc8uj9RTrs5eGeC+0qtGjSqsVZ6NGuJjmjCSQRZ2IAdci
zBif5tKOyN6NbOmtQiPFWpIarqS4HmxCHGl//tzCSEGnrDzlt8bvc/iIl89LOGoD
RC+GBzaKrDv4FPhtoyGCqyHN8htINSoXCJnPgEixCC/5waecKQkTX2aIkbugCt+W
uBaY/NITsgxMD9x2iLbPgqNeoNoGPVgfFIWNRJQv4g1tXhOxDDJng6hgKuuRG9j8
wtAtiHd5IT+t7f//1SYNJY3ysFVrtoP/ZBSe2ns3DWNcjHgCHyMPmFZ02o3IFXl4
TdC2WVNOZzUP9sRQi7Y0bwlU2j7lPwZifA/uwMKmIn9TFgRRxN8C86vbTQG+54Uf
4bMna917BJH4n5dFWxe08nYkyfakT7HqKS5UaDGC2QCj5NQMDf+N6etVulj8NH8d
obiKljso3TYL3UA9qwruTItEn0kLTqXKVD5HAhzamvsKrEx0v2U+Nu8b/tl3Mtxh
F/ta99Z5iGgn86c9Eg46VVRbP7xZKfGtwutpmYSyW2M13J9eRY73eYc/Rfh/Lymu
niAm3Y3TuGCMkNOgGOWKSVe/8kHQodAqnX8J6pcL/r164VvbgLxLAyy0z5+qapOB
HDsFitLO8nPEZlGS0Vixbx9OP5lWDaB+hoUofNGaIoDvYRAWFNkxAjPYjJWvqWhy
vKoeQxdv0itqah2NAFpp49rT/nwVWBY7SUL5T9qZciDEbFvJ9KdfxdDT1QCm527o
e6aeq/MjOpKjgJvK5vVehtBv1rqYGHeBuXAAumFhjvoQTVUg1RiM7r3xxGpPC5ou
gfa3CZj/W5WS2YBN+ngZGcWgyeWabdo+fQcl6B2TULKrUy8ysGCrwOGk3IuCNEWM
gHtM21ov/r8YhX0ptqzj/eQGVCeUli8oGtg1n2GmgjHuD2eDVoEjVneFwhoobpX4
/i10Sz4Be/Sm03DkUZXBBWpg9i/LELwAdqTxZ3P8gaOPa0MHJ9r7gNKSzX+U8vvD
RD2aCnl3rfwaKaK2zLVZNDCirdaT1RVw90IBUtBt2nTgpyWQk/jr9kMFiVgCXG1w
al7oyKVtFZc/Z3hLcpmfVe8XhzvJdUWXoZy0/Amc39fWpqF6UaY64oD7c679Duon
9veBfOcgbX4XLgtFYKRyxouB10KuoX2r011FGjiPxiT8LFkvaSUtarsAAc6Y6d14
cBs3+2bsJ+f5WdsHPrD/wcsTP/HJFPh2RXqmA+D/tdZ387IvZXYSxtWk15OWXbd6
APDlL9ggistkMsk64uCmMxGGr8Ppi79ejBLpcolE2vp1GD8ppqt05MFeCA50yzb3
HLix7X8pq+gMjdvdDWNLDdrPoqDSi/JBU8SqkOMfWxFzRfSOXlzfTXz2N6HgRImz
v/kZzh1BqG4a+Kk7SdCAKRD0etyIfWy62v5eSILqt8JEjcrFPZaV3Ik8qfgn0Dr5
sxOuscHWvPF0gPbqLcZEdblbMog/CtWj4LsG0+bcZ1xFsvX+zhs8fzUBKUZxD7hR
pyuSiXLqqzIejqBooEAZKmlE1Vzfgf8IwxFz1Aw/Aj3g4/wrNJatwK/R31QENhmF
nolRpmK2p21Zjn4OqV26sU5vliBRvfmsNB5jY0iIAvyx9cjA6b1e7M8NY0rHgDQz
3z8mIhG+z9W4vrP5US/1gpKAP7+b+I7+W7KMrDBhtokk4YEBVQmFVIV2FlTScQn7
EUYQ2Cy/1PI7A/ib4xn9WeVO15Qm1mSDmJH76MdkTNY2NSnSVikV8Tcj9sR6Rnn9
7H5tlodbJFRGCip1MbwXcFDFPlQzXYdRtd/SPrzmu3pOrgaTosgeS9kIPPReSwjq
/DPVTd+GBRGGCplC5YIOd2ynJKpRmJzF29rArKhh3c9nkE+xkVDN6NGGR6K2eQsb
Uz6jCZTUav6lkgZjBz/tw/kti+YqHW8sfWj5znUMeG55FOT3APEd2XfszJB575ye
/WQw5UsprAMl434x6Z1pUg4evJjXQW0YSaC7Z+rLjU58mDARR95GC5S3Wn4HZjVp
KUqB9Wgn1Tbu6N7tBrybJUyxGf2i/rvj9JOAZCJ/Z98NcCig5/ImW7AXmDc1Co0i
zV16bNXK3OFbKF17nC4NqIsrfFq+yp5BUijODVX06PRKoRD6tnYmnjzgHHuO8PNK
ouQrpGDcwmYB0T+vPq3UrdnN2b4jEb9sWe3E7FMgxf4VCcw/9TDJfKSgqHYD/IIQ
Ms2C+pz/bEeNHYLf9+2dO2lnS2OALAewi/Dthp5LX2tRITMytNMfh3nTwN8ck6og
TI51FhPXCVlzYBBFlFZld0AJwbsXyG3bSU2ti1oh/ljmjYOUJH6qf4fBD6Lux0U0
PtjbrvI+dbP0sMK3cYWgVW8sZrgjI56l3Y8R9KC6fC8jkAVLOSlCWp+kEibkiVPr
Dcjai3F91dAeI0PZyQpKIZsBKrzyEuynJYxzuigQ4c+DkksdMHGovkw1YZgFwvdk
M6TA+BrzTdOI5wump1die4uXhwSId2KBO+bocQ7mLcGXUtu8eozR+4OPMXcpPQFL
sE9ZpxBI9ZCbBNKZSiykh/JpJ5WnuAyTVkc4hE/idAH7RaVgfJtqCmkMlbj4iV/f
/oiL1eM0QTdgEZesEUDiUgXSVZ0Js0kJPktymtglpT0XVtuqX0uhoYJS3hCDZ/ML
fk/lFOf2421hpXvb3W5Nn7lceunovNFAq4YAeHF40BxknyoqSksPnXARuTZ4pGGh
waOny2JCaDumIViqatwIQbEucdAJFUlxWaltsL/+SEBSTGt1Rq84Zje3fLAH77cF
xFr2/mGTPX3J0iKAts5HMpA9kDa/OE+7+L2axXBwQWb29lOJP/RHHWOq7m6HeKbV
7jG537TbBy1qJU4ndeBKaepq7+ba5DMCcmTM1TGX5yM6rGGUrULVK13y289hKTp3
bdsHzxGjrPLNjr/euabmMgoqxu79OOgJMB+YXBlBRVcA+3vovDp+7WCY3nhgfaJ4
TfNe+mfEhppP5TXx2V54gzjOv1chLaCnrGc4/sGM8+iJWZFxpJhoMSR3BemuEQZ0
erO2ON6pBsFF9RdLihqUwGzpVB/FxSlCJXKIfUDGgASbnyfjzkPdT4ng2+O+GjT/
Gn05qyPqLAOoeE1qw1DxvRWu+lA95zC5MNv/jM7Ih7e6SwpUEnxM9XGjrhmt3gAD
kvyC91jZW4KfESH37VWkv27zws86i7UdfasCuo24uR7iI39yH7f8TIA5XT2ieBKA
9nLvGpXrzwwDXFL5sTIcCeuh2QiV/LxVeTnmsot6LdX+pyeurfShQlDGHZdbxuFC
VeqcPN1URxvdBOOYVAvjwh3NwFjkjUuCl7spEXSxk5oTQ+/Sd0ittxqaLTqzHtSU
duFJEWqWT2RXpErWYiVjOc5XteFBGCm5KNk4wo9n0ceTNdZ/leTdm+FHO46zg5Tl
j8VUpoJIdMAF9hKs90GQ55VJh9246H1uZnM+BG/M9Tq7ozygQ6xp/Ug8rRaU3iOO
4SYJWhNTkM8P+iWy9RzV/HiHAG/+mBfM3Sg6gIyK9TpK/LrK/o/dLJjv3Pv53hac
CZdZOOBuvUePSrjJ4GxniI07W0rhtwVnEMONwtKdI3WGNJmRPHKN06Lwc2/loHf7
h0tbbiOUSdCGFxrKUX8i7wKF0h/B97VTx35X3Bm0fMbSn2yk2xj4XuBASRxC7pGL
5BZnP0JUFkVGfCHfz9X3XnqcnRQY7TSuh4XJ2O6BHIajr9qFCdf6p/TwNhCbsjUW
ybKAsOMbB4NMtnSVc4p0oZ1K7qNKHQwfwf282AhF+5AV1z0n+ok/J7KXQSUqFvfb
bZR+SniOHvYZTK3MWF8xcX3hkkp/XzmsNyBzivWh87v4s1rDrJk2++NnBlAcdpck
MR8fEyD5c9HzzueI5YiZfkeDclWhs01ZCpywODQ/KbJ92ZOu2d9k1PMi87RXHSyG
WmyJg/Ca82CS0aLJ6c0OM4zSxRf0kgvVQIyCz8qdU8Srq3xUSShvre6A2mYs26L3
hGT0VuHZZcX89TMB8gmt+pm0VZAYK9PzxRJqmdc42SAyfGbQESyAYfmyao3HdMue
5r9HF56K2MThB3X2vJupU4wiQUozI5by9mIh8gSmwqt0QE1fUHbOgDEP3g0Vvwu9
yzkcxKFiiamOU5Pqz39RUOVB/zFOguPB6wPpFOyQv4v1fYMLHb6aWWCJsRwixW1b
wRIfcyHQB0Vj4X1/45eZR4JQu9x0PDr+4VlzdR5WygqFAsm7DyGprq+mXtdKNbIF
Hr0JDfhzz1xlYL7SoxWUVhLnWQJdAZDfJA527UXa8fK32ldkebA0ZEdt50buBzeU
aJ3YmY7ETLhj9EkE8MSFGWUYKm83jT8zK+lQBeEirPkDWUBhkvfSBvugz2gRGBiN
DZNkVntFonphAre7vyfRCHRb1upY1nTt5RiV2cXLAywJJKbx+h1n7JrXZp9Rf1BO
M5LWGcmZp6KdW16pM9G2QcmBdXmkG2iWjHy8K1CfKGuqKKw1vdBSMnzU3H7EhBrO
KCZG3tbTtTy2BYC0X4ITDUHglnZocH1izhjbcPUWcsTl7enhJCEGESZ8Z43pejgw
6wB+2jJi5tWPYojUJW99zVmg0MhOuCQnczpxSCKGd91Mgi2Zi2cmpsC8KhgPliqS
tbA8GzppxW+NlgheXq7aeKvevZNYKC5OUDmwRo8LR/QHgBpjmuAUffaLnh8nzY4M
30FZqYX2vp5kIbY1eMKKnJ8eWRC0s9vldwN4/OX17nVf5wc52sFh2VjwQaCMkkKv
y1cMRI+/BwXkhNGcSSUn1DnBCM2qBL1VMLMRqxOA3aK/PQ8g00T8QfJJy6dyQtLc
MxucUakoWzxaRdEmqv6mBsGPVavKY68EcOuVCUOoUeMeKo3slqd9e55iA7GFxTAQ
QzMQf0WWhjB6RUN3qE+N3ZgFxhL1Y0pc0A1v6Kjg8gEontHCqW5Q8TovdezIAxtP
0Qolhy1IK4REUQPmrtoUW87/N7r9YYUDH3oRqTYMvvlGJi+8o4/cwyDd4/jX9T7W
NPqpv/wYxocDh9jXsyReOGf2CMKfZiOjUBi3QsksvEAsE+4yTZG9BFWJQVvH11Qv
Y4fEmsm6xNJYmgcchHQiNfoD2ZDio3awRo09w8VXIvpDOwT9Pgom7PSIQfMqe8nr
jbUBn3gLkealaUdmXHsRV+fVodXBbpJltydgAKvUTkfrleAgZwSLdip0JrmC1pNq
p0kad+n2y43ORw24UUvLYXR4zq5Kz1Y7Lh1FnQfrmu0RO6QbG4paxIfN9cL5IS5Y
jVEE0uZ507W656xMCZrmGZifXzSJKEIbItHdYA3bnmF9mINzDqcsq2ML75vjyVMI
1bwB6vb0oLlIPYNN6bob+wIUgxfE1er3vslI2W2oDk//J+oPiK6wBqzrbvOFQcNo
iEd+vykDOgx0G4Kk35reBduD2kxDxIAoV5LUUKq6CBsKd21keEfNlaOA6vOgwHyB
24XoyP+J2B1qXBAPbRTmXRbaY+NmU872VMq/qNQFy6zlUViffGeVtZMEjoKOEKyk
xNCdu1ZOj1v+M2saoAT8EeDIk8Pa3pom0kdOwM/Q2LVdVSm8TIeE4/etzRBWE/6b
APDcxtitnAfHRpRC6RgLtsXjO/JW9IqD/J1ckWJE3B3sQcQowZv1sMiwxvaC/lhI
4Bb75wF9MzIpQq7iDkH6NoITLNNntQwvbQFRJueslQU6ERvje6Z2AYsfJ/l/apYN
xOZT0ZUaq9jwbWgizJKOtR3/zEOHt8CoRVf6ZdQFWbiZ3NwhRXEw3p8J/mIxjdsH
js8c1mxtVSEpOzQQlcIAjaC7Bz9oQROkUrZX2CAXcuGZpbHVB1HKKNwW/tZhCCvJ
VF1s6F/YG9mYh68CvEg/l3wmY7QKDEUUJT3PgO4Ym2M6VELHhWF8+q5O4/M9gwML
rShXKBXqxOVOVxKk6hn3M4PTDTjkK5P+PiwnWsEwOX6aka4qfJxszbJiY84nGhd6
POMGpnokDOUheZDTGxAXwlLLMrI5g4mS3RGO1i757i4jTO01LmtiKWruwmCVdzML
qSfU5g70zMkBfB8Qznnc911PEUXsRoqM/QShCZgQ031cus/6nlGfaJYerfx11lVd
mRP8hWPkAZstYODjniqCATT9GMPNpkmBT4kW0QYdKrEUcN9RgWwc2lojvQpdBEFU
AgNL56wGaDVh6q06E5kwSCfLFYQDKfmUc0d2ioqGgPw0neMQseu5fuwwPoSYdQ11
2mfloJ/2G0vMOP79dBxiYrDbrJ9nJQR+vlZTVwAOY0j2wwT8FM7XlXS+llQcQv8s
jhFx7DN3WQgQJWHn8Ri8tScIT4r9RxfS0x1dnEBP4rOIJN5ndqMr/QXC3g+uI6WK
YMxYL0I/VmnmKRvLaJTqM7jiLx2CZeF2b3BHya94IYd2vMzDR/IAuIVXXYH+UaQk
VHZXOwNCBSMuGsgznmZ/de6Lhu13FE1GO6HquvkGZ+vioyCn1qdVeugODcZRVJH+
kt2veeK99UlIZo1gNp14qZm2s1WZk73C2J9lkccS06iK5WPkIWmryEl9RkSrn4im
ooJWqUDmnm/AvdlyWiGvrX7m2MoZ5JOYQNuCd/gRaF3RaDOOwByFbDcUI9X+emtA
GQeN9tpFJwOU5Iribh0CNWfqBxq+1tNuyyiNvy2ELjMlHNdtWe9/7HnNjJrVY2ht
foBru4IfHEjY79I28ZXoyV3alDWlhgi1BjIXcx0hnObCxVR/YghdUm7eLlHGxOnN
8TPBeNkk8FA5MhfE3tbNW0R1YFo7WghsWlQB1DHUPKBUQm0fcVYQ8UBbzRK3lown
lpJsw6FVIjOpL6RCxKEBAMgV1R3kD6cyA/ANFXLOAlEN7TFXHthnHJT0mVCvoJzP
nF9h6iSebMWE9eNjQ7GLirrlPbqCT1FHx3e3HnUxb2BGGIs0tNugqpggjS3eGULT
i4BXXifcCp3bw6fNTex11NiAVb5tmsJIWhKiYhXaI6QWDNC8L4FsFYGlMes4ucaP
+gDu4fBKlI1wMWG0Gi6ljbKLdUV+SlJTsj5vhb6Yu4ra+hk+MjGVtbzkkbKYmLdJ
2M7EE4XLvAiJeRhO5/Dhrzjfac5TJ7UzfPo8XR20gqqbkfTNw8u1b/zV2IP//2Kc
lQP1mdKtSBLdHVv7RkNvtuRFgRMGZqNyOd1HeUuYpOlXafOhKorRY9Z9BnnWpSF8
9UEgUgpFoieBN9QySoogxc1tOVzdCqMtbce0WWT9vW9+7+aWGLHJlRX8m0aP2SC6
diXQa7uG26rgxGl3qyZ7TLUwxZOUWbfEeFELLZDG6IqmYOTj9Gu/mRbhYGnV4YgW
apyTinC6D4mt6eJ93VHWVG15Qf/TKFs/EVThlQzbhmnQFCwbXZ9T84ELjafWoGpn
qrUX6XOGCKAKCyPlpkUkR7lMrhxnzXKJ/BrhXpyHyWOXOkzsW69VGfqErKdqKQHQ
Ao/L9oYrL7D7hi2F4MoZSEKxmFdsE9g5fPKsv/NQP+orSm+w2UDNqVsEqRaFH3nC
KNbZG5B5QwobXlTUymVxa+IYFWE+vHczdn7xtkjURU9yqaC2GcF9V9ekA+48qCXc
dUcg1H8VglIh+U0OwHcRpHs3lMNNKNWUMyPZIAAZWuuvvBOqg7yK66Nuvu46r5YV
/rLq2cJ7p6AXo25F9TSDFml5o35VCGxfK3Ehf76VYBVJj36VB4eyVNah6GJqllWl
IhKoggNImltwvwq7IWdSm2AYfj/koFPz7gtH5YUCR88NPsXsX0F7il9qygjYTIUc
BwsT05i+y6ySMNv9nAVxexuAmkIOs5hlEvate5VkrU50eFZgznx3Ggt5aFuiLOjy
S8jiuHJAp5B70q/QRTwVebqI4ok5QMNolhDiwU4IQEzDKDg3nIZesef41/FrLLyD
vkFh8qULIjvBZFVw7hxOTmBqgCJ9XJIqf4wVAilhZzHTB3Ul5sHB6/FDqPw9ny4G
7khABmO5gue8bxoWIbm2uW1sqS2qbkVt95IwrSSjC2Bx2zaekWgz8Bcz9PKSOm/N
eV52cNy89NSTqr0t32U+ltb/4aW2W+aLEt7KFC/LOJEmcqRsbWdszLNkLNENKsdu
a942yww1f5y27YF1ZPd6PN/DqsEhD5gxwV6BwhLCfnjT6rtaD/144h5nofhRnRoA
n5UgWzwr2cdpFbT/af3q+/pHz1VpOgyP3+NjoaaLh3eKSX9/3bFV+Of/oJo19QWd
o+VpCDlN7as/TC6zqqOK+0yZvlhBGGjn81YT9GeLqi4mJxZONRv6JHkFcjJ299qW
QrqOnj83Ch2eUQR8XA7jGWDq3kKfqXDckzKgKQuXE9ieIQBy8ZdzIe5c3YbuJlKk
mN066eQiZVa0JfNMVtTfq2gdj7upJGPdUc9VFbKXxrUh0HN4euyRCWwbv5LbP0+d
Owzziddj4YCMvXFxjB2nFNVgHTnS2Pb19zrMxy0Qz4g8Be8snkjFToOyy4qns1QB
yb6OQCgf+aLyof6TXnI0BKLOWWMrQWKPOhvgMRlBVg/rqhBB2lY+T4wbLt39FN74
lt4jOvsLBO8sO7moiCCylzfUOgWsjRT56YuExh1J4kFWV+PEryBjCm0C3Naz2GcA
mPKQzQ8lRSqu21/GXsXBics2GJxU4FiAOoS8QAHHOgPJQQUYXXDmrAocGBdoLVRO
m6WBPQOJW/fCREvn18KENtvVYczikaf86XiMZliAH3ZmBgyXDD7HvljoCriNdOX5
lHdPdJU6sjJ/nqNvHYHZH8Aoe7QggU/jtSOd5fgZd6EBpf0afRj3Dh/t0hiY64AF
dx/g2eh1fy4vbck30AOlQIREP67x/D8NkgtjPSD2NF6VzFDSOTVJunrE2NVTNqz2
TqidT29Sb8DK8FBjovJ9ykHd40amPJDDaggLON7VTw5/UjmlxGK+edoKSCXIZ7Vb
DIF06/JsUUL4JDOhzyTcyPNB8/ghHQgZhTqlYghV8Feg4mVMAddujTE865XFg98I
LOJ5t4ZovjT8vW+vgAgkvD0D9v1C7Przum9ZyIy7VCYJ3/c9fHahiLpu6LgJ6tr/
rSPNquJ6GVZH0s4kG5saceMMLcU9H2FZ+730vip6XOR5ImoXyEj5knzMbaViKWpF
doZZ4YpUXIk81C+yz7JZMyotDiXKnyjD3a/87kSyFfCcpySMnILuR2Eop6QtDSgf
aCbE8fKy2oBzP8gC3r3x5oA6sl4oe+Se2XHzpcemKP0TRb4iTTcy+BbEyPQp4+7n
VoBZ/MHyUM0daAm6A9QvlbwQdaqrwAIJaFPjfLZL8oLv1bx0yTq+joYHkUalgMF1
qLxj0L+j+HwFjYqFbqzuv57A07U0Iv2BXpcjfuunHv0zyJjg3WZ72ZkpCnofrJ8k
5AvoEW9MqFs7rvUjjYhjO7gNFy6eEafokfXqMa+NREgsUoYQKREDalKbEsxKLR9O
EOI3j4q9XHq4lagN8dsnHQPi/6/s04w72QV7eEn3O3jXBLT5Dpr+9/JJNB1OEWeP
1fUIaq3DyumVSAGduWPlhdKaw3lfqrgsGXoa8qSH7WdchgH7YahLs4pJpDT4l/hd
YpuCEpjTeXOqToB8Ep+xOZuuYgAMX5948dNIVcbopls/F1NTqoCb1wiItjb+R43A
aRgWhibQJ06OVgE3oZqI7e237CotXAX/QlKbWlbRyiJ44z6vYRTj3kfQ4SAJE7k4
kD6YNVI7o/I8nSn9Gc/mJEYmIypr7yp1AY2/8axzZLFUIAx8vl5ufgRDEAtgEYjs
YpRpoE8Rx7sTh7Y16h9NHp3NyNM66QoiwO6Dte2s8uh3ToNExZBVYkkXuqBSgkiY
0DZHamI/vBUD82cyAZMqALVEUYD01JGdzG0OiKIrowkS+j4wsH254qSUTLsEt/zG
gXQRS3uklVWUARfZ0cTYKCd3Xb+/45ugw5lQZMiMR3JRi2FgaR7mvkdI7w4wk/W0
4eKkS+vxKdyzxH7gzefeOV5N08FgShtMRZ8+pKGVToV8gAbJxOSG5ReLhZGSTYc4
9gblGbMvhb07ZGG6GhdSlfp/XWvuM0rGm+dSm1gP1agb2bdzMH5iZz6bTw9G4J52
n9k0sAHfn0o6BDvmEUhJP2C8Gr4WHHG9YDV90fOWtAbBhYUR+OLHwVgkxoQwzU4U
izpS3EVFkt5szzBvJ60hX1/Wz8G7CMN4hexPkfcfwjSZ33xj+0/h5jDosqJdN5L8
za5/oVyGRno53KAY+6M2rS370KO7S1Q7iLMg9FYSDxeMMJ/G9pr/eD5IGuXNZ4g2
8Yw1M0O8Z5drC+ukr5eTJ978sI9k/z/KQo80PujW7h/HOpNQF/oLDhZjFrNQd4WY
0A6xtVM4HKXggTSgNoioOdemv+O7f3ZUf4GgEMnSVZXTrYKRRO/CYx2Jp9vWwp/H
ydvpFHijWkVNr/O4XpXkoOOQlZNMhnBIW1N7+6Y4jNvMJQpQVKfsipPyapkq1Nsa
bK+P80ft+yEn8pedVBPXVyoaqrSfhISxmanBlEPC65+S9c+ma02a9ilSar8Jb1C1
k1Rq7qIroJe4cEaA/Dc8gsLAGjifDzm9+4O9QEHiOdQY0eHQZzBZYAVQTG3S9ZZ9
NAXdEmWxp2v5fLtQRwSZDBOFlg6LPNFuqvHRCrkFayA5feXtzXVTmGmi2WIpfwH8
LfCYj1aDHRSqhnr0DiDDtV6+uwTJMT6f2RIxVVyhSEk5mmCRtjPMArDzbeo3hxpS
ROZluq9R0g3K/zNdV/5N4pOffzc8QHLxfFIn9fwajPmicaifqcF+qW8TXIfQikou
j6Am0ziEMD1pYoupkAPh4AIZNy22pFmUekQEzHRUKd9vGJdZhlaAyBUAtADKLwL9
iVrRIFQabJIR6TDMCNSVZa1DNhGtbC+xDeXfip4RXmdZQygdURVlD+zxpVf6ICJ5
WOdLlgFY4W0gKhYaul/m6N/5RDhHdLHIKPYLePH1xKasx6jVB7l0ymFb76ZklJ4e
Gqkw5OC29OMmDfVgnAFNAThR8mV4wPVASJ0yLL8kI6kGGt4AgklTPvs2IikrUc32
KcPbDD0R+955HsgqS0UwMWBiuFZ0FBrANTP1/rn4MkQIyyJ7huosAiGGyzmPTCIg
YBp5Oo/79ELSCV0DuJGJ1332hHIeDjTK9uDTu27a6eanoO3GUFQrh8FVi6Knf3N1
pJG9rW5OBIUwLpwWBXh1zUOxtEgwRmjE92FUxcIRanRtBh1nmHZtT0EdXkVN8cin
qM0dOL4tWcO1oVTQQ9NwTMmPQlkSwKdT1lvtr9UdQEtZs9s/GbrIe68ByHRmhvtB
hK2mtUQDhXd7nnTucuNxhQ2wSOMw422ibK3kfPJUfD0LdYf9idCTnT1e7+NTzUie
u55MdWB/4F/GkYzNI4zLIfQeFd9JWQq72EoOizfFBtVghJoytsTWj4/d9HM8beL3
APrLMyvpza4LlMndnlbzTEt4ke46qD53Pd7CRiP/ViSI8vbBgkD8YixzzIA3pSu1
oM0ENIhOD9gLAhVgkG8d+xeAKZUkJuW39nXmM3Za29B8HkNUyPpVLLcfx6Oo15uZ
OXi8LPJnBg4RUJ6uowv6W+JRsM1K4KNzlEcjl2fdwj9d/y3U+m4YLYL3xh7XRCkA
B11P6wwBVe97Pv/pjTBzOqNP4hcDiAi/vu1Z70esQHeBFtUGQ1K47CwsCQajfb/0
+6ViVBvzs4+fCDTAq4Jz9T1hC0l19CrL8PCAVU8xBrnidT4eRsF/8K2mptJUMvl/
NbDvTTJJM/WX/ielUGSKFEn3F5+eljxC7S6ILTqRjkh8EnXKYmmiSKrk+bYvA+H3
+6gBRZSpJaCoXlPlww62i0ZLcnjnDLbyUCTIylo3zaFhMrAwwTsh+jo+iDWYURYW
MBwKS+C5rAayiBAFxolVvdYTNHf1GaGg4VzyykgymTwtYN7BR5dGDKhFf8Fjx+n9
bhdnY/itj3RMA0GBswny5weFfAGlFfqbQVNYHcI6Z2NtgMqvovUvzThxlNPWjhKP
e/tt8tSxKpnrYPqKv/fYiBntg8tg4wVDobYY+4+/KURwrCRhbxw9L01TPEsd1kfP
QOHMuYAXq1keB3vebmX+u/3y+MzfcWhdEa8oNf6OfDlgzrbmPkYVOaIz08ftB14I
MwC5XpMNcC5/4iTfemttogKo06xHwhIwgx+LCROqaRgK6Mz0KOGLirJTjBPSm+K3
siHztgRtdb7F/IQXh9fBLdZeMI/XNPCYGPs1Abvi5qfft3QqzCku+Gp689h170B+
WzRHetoNnD0i3F4nP3emBg8EojEWIjTJOTVVaSQQq1N099Ly6WL/ZW7T3AqS058j
BX/gnFxemEqiLmo0cBihSnBZfdyatARJVOdYHcRYE64cUJRpLtKfJsxj/Weyxvo5
yjL6AGFr3CYorDI6Fg1amUOt0TMrb3kXan36DmpP042XB3jG+QUyY0zy22yxsAhr
wFuBenbVGoZQMPbJSGBvNdelYG+QosjPBAwje29B9p3iVijvJOgBfIwhvFiuOvhL
p841R9FTttI+oOUwlKJ/yTI+p5rBZeoKyLSzW+N/q1p54Nrf6233UimomazwEhFC
Y9apRXIW9ZINZB3SHbvs3tmScIscGreQZ65yyDM8Vtl3rrpNBlW/ge4Pw8WUr8Kf
L7WlxpcMfMrKqXNz+PEd6nonoEcXZsAWTEUb2Zuo2H272yUn7eZehPGMxrI50/Nx
/daewq8ze7vU+NBgvSNvMbF+rfNyn0On1K2A+FfRDxEIzHpbNfkMPATZ7WVvPEBR
Xcw8juz66bgtV47OfS1iVlCE90NgFhQBq6LB0EgwpswqYTQ0ph8ozoEiE9tDeHQv
OdqAnnAs0C3XJMnzEw2yVGh6yps81ulnGSNmO/DTmJu4Ci3voarVRYkdZyyi7Tsz
Zi5WjORDdpnsuqARIxTjCtw8zkwtVJtaUEic7jJu0Ga35nbsBOjPtO1oDJXUTtZE
NpYO4+WoufbbPwDeP1ubsqaiqjq+jYCgLsUut3OcbifS9iyBZIv1SISya+xGe8Kc
flV2/vF0ug/JXOXfXi7GQsuJe3S9JXjDxG+97EJuK7zJ0E4/Y+R5vtJVdc0SJsCF
O4GaLibSo/GpJNmEk1oRblmlzcSxd7+pZP7TvGbkyg4fvQLwefHfQP6N1BPUQxiL
Dyg+jvmYfGR5BFyn58EdAfrJvy0uRPLPk3lwpjq12ffQahSae/WdQ2jII2PVF90h
lYxThSqVoW2qm2AI+4HROOp/wu1kboZq97S9BNzlU634BzcJ8zeavcknP+kx+OQP
tJJFD+Jh5wz2Jh/Subvu9lXJDOD6USmRgl58PWTtKeNn8Ah2T/TaT2N+08wvmX+v
U1MpO4tbDRnFM3xv5ZxRbV8kG3cTOqKemyIbYTJpowtpMTMFk/YifRWv7k1UbY4E
5iJ5eRVseE1gAUMoZSUbGbgG8/i+o/K6sXE5TeDm0PwejwzJJ0a8FcNqyFiDTrwF
6qi8f3UI/f0b3twNLdQrRAMfzhTs2jozvNnBNsO4oQ0DI21J+se6znDbJ1id/mHw
NpdhAk5ai6Hm9EG88dhkkpKTsES9GOP3Stg+9UdaVIm8nXtjF9TLMMyrttrPfPrC
1S7MpLMat6+VGqXl5ptTkNPAdycHkBNPx35MQxoXw6sVkJIxhIHzB5kTmpNi2bb6
ldZ5opw3mnr47fAK4o8n2mhg9buRTJi/Q+cy6pQGgIbmRTOxT9bP7EW+oK+hnqJ2
SQ69UUm2G5CI7rqluJbfW9Z5JK/0ChjJlQ9GQ+AcZkGiypRXu/0EBkuJA/nFUmEI
1kVSCAnObH8YLnIm/T19T5t/G0B7pLqFfcjBzRuI0+dz896oCG12gFD/ldCAzNCr
Yf5dE0MMt4pHsUAc37UnnmncSlpkglxOXc3GNI3PoBJMIuLYLRUhybGqCO4UhUGo
eu+OZUGpoIa/sxFIuIIr2IRoRnWr/UPLtLRpkvFRREX09uZhxIA0VaQ41w3GkNta
3Sf56mCIYfXMZVnJ3VUEGX2AapYibYreEEKMg8sU5FzNiAwQFlAZ0PDyglG9Bexh
Xb+ossL/xiorotnbWWqYDglq3CxjJngQB1tyE+7+oYdzpHzq4RYZmjo1yAoyLTKP
1RxrdDPYXZn741WQiGOHTu6tADhdaCLjYuf1k7eRiNfZZrllCEKXRsbXCinqY3S/
mAulZSMoTMn5EQwFotSmKAOvdHvQ0PLkwdYJ/CfMDgFLnD6dC/PHvSVAsW2Fo0jc
l42ZTIRty9WASXXT/xj5lr9+ux2OLMfef+qcLqMUaWzKC/o+DCQswGlaNYXwYHj5
5QcGS/dwX0zH7BTiWnPr+eQkY3L4H/pCKhUm+5dOHEVvIiuPZFySdpesUL0SiQg+
KB+n0K4ZzY+Be6Ffx1QqiIChAYui3BGJJlwq10NtD6OUJNHUhQLs498mPyaJptxI
Af0IA7Zczl9jkJFGtCkvk6w9vTLGJGjbvYZRIIXDdU+m5UrMaOJ8CIj2CSMRRX8P
natJ5TaG2vPmLGy0KbmdGQ7TfFftiEzCCjXnD0zXGDzXDBtNMChxifDxUJGEPcHp
j5VBdfwVhAFvttxEI8PABm5lIoqjZZizYlJyOnpUldO9TZyASxjsYUN6LmaHLeij
YuyaJeE0hv7htJ9EEIjZPwtCHGHTc2vWfp7J+8xf3xPZE+w3pDw77NuJ3mdv92Gs
wpupolNDf+qXcGmbzXExgK3zmCAHa+uMbF1sK7O/As6vr9t+UJOQzp+OxeEMUMRk
yEjdGOR/ZpKApvwJmdsPz05pbk0btzN0y8mj78THv4Ihr33vRxltw8w0Lo5mesMX
PA0bsd41e4YipqguR9j2gSOl2jLcvS40MoN6wP8KlBUPLcDWkeEdx53PPpWh1zoS
FStZgROo5Gqhg2K9uYRPoIvWC1hBLZnigKcN0HuPK8aoNd1DdIpp8y6rJif2Dam/
6UyYSByUTvt7oXkLiR4nP6WaFSgRvRoMvt5Jse4q9IoTlGm6lp16BdnThuUnGkin
9BXccyYh3nM2j+pCG8g+9qvrQwdgu/atMSNBRQnUBuVopNs/HjT6Z3kRaDvyb028
QpfFpbrBaKCnWp+ptEdrJS0FuTCdN/Ug/ZV8ecGtc6rASLdIoqGBFMwcCXCAZ3Pi
Grk0QQ+2ZsgVfXDsYeRcKkNI0pWjfD6UO7sCdXYCc4c6ICVQ/gD5y7VfC4niFp5B
xB4lqe5he5RFCAVs1QX+VVG5UWXO/g3qXtWBOTQv0nVmQ9SmJT7LoufVWGkhWdrf
dkaGn5Rb3EtsZS8v769GjuYolcfe5lqrHmhViIZbF8ZXOLNSFWJH7L8pmLRV1m9e
Z4EJE9DwDNmkU34jTHfCqJfnzlMtaLKMvyhTlEKhyBUwbM/burj0IHxLgR5hEe1J
jg2z9xUYGb7A6PL0zy2lXA8vRP8Ev/74bubbsFEwP33UPTptAxTBqaj4Iuex/G0d
JGOchCZmCAszdVbcu5rzPtO5C3792w1AnyXMnuH5IMNJG1hZxHxx49crXhmz7l/t
nHb6dV/zzuc3+wNvZVluAjARGFFWDRtfA9o+teijAz49sdMctPp6ozhVtveZj9kN
rwhIGqZVADYrBirIq3Q9pxGIWqsvIntXDLBShVmOtKCwuPETiPDN/oyggkWPqqlq
pFt6w/FBJjlfkKL9wsMUzcDGNspj8NGbgWqKxIno0xGpdYN3CiT7u+fUB16GoTkL
bct5iPgV6eleE6DwQZCyBP7mwt2ysOibVN5eGU79dYlYVgWM1kR+I7pkIZw7o+Jd
svAmZTojeT/gOyDkLVWiHx0OExrNV0GLPdagiF4vRxURWUm8rlZ9VraOthUxxRsI
ZqVJDBHQHwaFig2aV1wQOQ+C2I2gIlLCu3kbyyL+cB3IUHj7/CMUxwiiIBQpukvh
aWFQ6I//2EZpK5ec6gnoYTcsMSiv8gIDUeXeg2BWYi1BT/F8Fdhv9PNBsle96HIm
or1zjjC9qXove+Qbf9kdiLF0M8UwtImawNasHc7nu6QtpUoOLRJ7OYrQveDzhOT6
IgjqqXXXw2tgEdI7gcopV5ogq/qMGA/fUFII5puxYj6+V4PLYjA32KQgMFeYZ3aY
MDwiwKM0TsxXHJAtF/83GQY//OfHP8Fhkkw5XW4B3XLLB/KgR8+0VrYfF2p2N9Rv
KbucCkDPJqxv21+VV72lWA5WEqy6NwQNK+yBRg+EpLILLmUANfLiT1aqWfy49TC2
fcNZrhLBTY7Po8lU4ep927D3XPT3IpMZd0AABxWBBlXsVEVg4yUg9QdbraWPHzRv
bvivHOfbQxtTjgldka6miI90rzTP/WTUGb1ZL0BDSqthPAuJWGrDnK72hXiG5cH5
Xtuc9CFuxNyIapDEtu+XlysFT/5h+L5+fZS19cjvJkqV5M9mGyGvPnRAdFexN61l
urrntruq4DOSjdLsIjnGdocuGFWBn8qsu50sV72H3ik2Jusnb8OSVO4Y84pGcdF5
xAMkDUsfEeSkQZAX93gFmQWq6ocXMtne/DHBT9jkXGHUE+cJ8KJhIVpoNQ0yiwSR
8hE+Ya0d6IkdrqKJqiebmAJaV7ubv+XxVCa2wcqTUT6qQ0n5Mnrp01SIViZfi7qC
m07wv0brVxgKmcnYjJbQ+bQja02YSfn+51WmqHp6UalxHeMxsUzBYhVpmi65foYt
wqGIeenYr9EHMfBEkkeTqIa7MOeftY6AjQlMHxGu7xz+mwH75yisbBq5is7AECia
GCEYcqrZIl+cgfNzR0llF2YL1MZm9SP9XlzBYCSxtAvHbWGpgxgcCy8VqVBIQAcX
+4uJq2FDBdvSWxZCmOCeBGViG23G6RLTANqeRbUO7xMHDmHZ4D5XzZOpq66kuutQ
jv/2IFgCM78X8QCSDR63zVkJx6FtBlNAyNE2LSmjqoazlWEY2qPVC5afpTZHBzku
7pyHg+ygRXmySlGbwu3AkVfy35RGOKuL7624z4tF39zyftbuLbehRLdhENSs3OAx
iV8MmlJaHliVKXZcYOuoM1446Blz1N5WMz+AG7Jlg/aSrETi/lmFjjubwutHys2Q
R3vx5jPXylDi3pF7WqlU9z70Ku58E0ocfuJKNkjAdfNromTLW7sbJjZuQxCw7XXz
ABYdoCl9EOpqKKmzLO2KbDxC67V/YUL0pK4SP5LTcjnBVErxK6HZeTp8t0hBmFyJ
/VBFo0P+bFtfbs2GnRR5DAiOwvDHuDN0S/EDIAiC/bCpqAM3+BlhJyg6vZJ+JwLq
emgDJY+5ykWFMOj1fsCAQ59spRY7qTsyLyisy5d7bJUYafzAkVJ8oRkbfVMn++57
fjbvEqUC6tqHMl+tiH0gzbvPhTzNJcYuV4oAmd7gOJdoq2PAPxyAdUtsFRyPSR3M
5gDgXqRBQpKcfM3nDW0NOaW7wsPwHlH+nXAVoKqS1jULrjK4GakZZ9B7mZmXpRZF
fx7HEIA0MdrGNRIog/KhT6P+MLzszB3sBUkwnmj24G+/x8NQ8Ul76TJSzESvrZ69
TKA0XRb3vCswZVHedLnQY6pFChUpefizc84cUes591XVS2aAoz//meGIeUc5/N58
y1cll7hYmEUjgyxUNk8vsMQLygeWzfXZNKi97cKSkVyULS4DMjxgEdSAPWFtgJ+U
hYwIG9co51Ruusfp26K8cJ0IdWCnF4OSwJNRhGv0d+PWHroho0/EtsTbXulFd3Al
uoIkbOsnm8Eq5VFtZIsjo5zcZqj1vV85VmdpWYakoHVtfzsGqpknzPY14KbE0TLi
3iK18RLT9h/U35E1Anf3W8mQxpehNN63Ij65TM73QYL+mF0KdWac+ClnADlMGL32
unRiGVBJ1JX2REzHDAbkvQ49+bbnLdtqAHXtlcGClFUE6fbNDI/7LOAthLbTZKeQ
uf4pPHNGLy5T3dmevDnpAXhLnvfcB5+b9qayWm8vbVazzJrvpc8XXUlSIGw+YnuV
I9EPn/uXQk1nQ2u33FQ9az2dCiiZV4aTPi00vwlwKstFDvPXq0l1vKKSHFveqJCA
emKJ3F5juTYCJEz+GbmfIr78HCtosrt7jGx0st8V3uKLBYCezsTkaDb2rECHunMU
5aEqC9D37Cqz2Pf4sb/78hLk5EwdTBrP71eS6/JRpsCJqnkkvS7UcaaCBZ3RkQ4I
lOGqwELNKgDSoet1z+tpGuV0VjcaqJ/Xd4ysNM5KYmch1bEQbe7RjiM1eeqp6eHg
R0hTvQbEbwSINkaVcr6fAb4kNs6WuBR9nbxa7b8vqbHDSuBAdmSlXfwWVUZhHtnR
6P8+6KQvtNOKXoDAOL4vBGGwwqZU+Eu3T4y1wx6D3t3efFSFSXN+i5X/QmP5jYb/
oB3Q7dnqbge1/+puByfKq+WmzJUQ3GvI/5fY/YjSWABi3odKhcYJBpmGhT1a+mKI
Iuc1haYUv1gXKxCYZc9vcfXOh10YIeK9fYzPV6HiosEQ59YYehxIUTqIXSt0SY6/
/ZAevu+HYG+7TsELu16I5XTT3QJt3K8EwUj0aHlM2E1769oe/q+YSTzF9FbEF/qx
y8YEE9GFU/TmJNvWv5fsUOkNdZSZ4rnQes9b8a3/r4HOXuZSfyMAPfDj5tHnsYup
TaeX/iKt1aXAK8WMM9ZdvRFxMEAxITQtoEJp7OX/f7oJujRBlvWR4b71e0iRHpO8
e8jVSxLPp06seZuKZDhH9dywQHLwabmopl3WCl5/E9S1n7luRA+R/Zzl8rrv+nj0
PMnej/dDbAVLo+q7M50nog9KpFh0GYH7+QrgA1TJn1nar4ryAQiwlXHkICySRDdb
YR4MDOYkLivIaxfMwkWx5zuZNNvrQBcPP5vf7+zwQq83TrKeUnmr9jMdUCa7+BW6
VFYgFOgZSRWHGc3fC1Fk52nnNoDqqq1O4KCNAFhzR8OwbQVZTtimt6tvyZ5GOuGs
p6s+fMVVMnZIsk2SOU6uPfLFRgOyNLDQkz+qXzDgX+w71Gc1CiW4sXrZ3R8ep7Qe
lH6hgS1V9Rka5WBtrqwVuwjbza58VjZSxOCw91j2hJ4cQROgNO8IzmV5hQRviauY
KuK1oszVf90k/m9Yeo8yf7weyqbWypG6+gABagPDjsnNWoQVC+pHi1hKHnCrqbZI
gOvryU4xZFz+YPum3IqM4GvvPQeWtnF/7XvZjbMHkiN2FVQXX/XS8ze2ff/jsXmA
kZTCHfWr/yCzqocq9pwJHndtHfy3JKkiOQztJiT7BO/F+Aa86QEFNkcEXrDdvpAj
eshQvYTx23yvjfF3mAcNhJlCpjDmTBY0WlSzyh9P1BkiKyNomSIq8qPXHMKC4FU3
ZNGk0jkrlbBVqkwO7lJGd6e5LPC7lc3+drMMnLTeBmuZZyOdcuRKLfb/By5ACVIC
TEuT8BPGo8JZ5XISeqrYjeUGhk0KOQQF8R/7lReQ3GH6mAkPWAECTPrFin7A9Cgd
zupthg751JJArWmRyb0grWC+G3MVavtXejkm7ZVdX4rg700b9zPHt2fIR/zZDKXi
CsMRM1UAIgSAvRxbhqMuoyJtxpVxPnldf3KJ+YleXBJDdV35rQyig7E8sISntkl3
Q0iM1FbqHJyR1DL4Vos89aL1uRKj1iZrGF4O1T5w0exsWh56V31QDzql3r4/oD4m
8IiqFb7nt05nd6QGeDOFA/Pr/lfyULOU0zdFrAzSkF36h6XMXS7wKJJEB8D8I1TZ
t7Deynn6FKJleM9/e6WU1qckrtjtLEmHosr1bbggp8JBjMPz6JjbKzHqZR176RPx
p55CEoRUT8APFvLa8KoNGPfFW0y8c64uBJNZSQrtkzQZ1evnOBoeXFkfzpi7Q/I0
7Pi0kNIWmzxgBA5p6278uOW8phykmQ4jwOlqUy0B61vSzuvVBHmikzByRzsWkhrF
mQa/0v/2szCEw02OvCvD5hmN+sV07y3FLmO67NHguv5ViT1+hRr3Vmpa74gErI1b
N5lC3ozfl6vsHOwCIMaS926bLKxnku2RhjT5E/RlV09gNiKph/AfNQv91ofBjj1l
TXrZLPVYlYjhYFbHGz0Ig+NA50IZjaYhwMHSdkDgPDsLz69cSSD42ovPkSFxbg7l
gP9Lvl+TSOEE6AjeC3J5/f3LRrdGULPUoS9QzQ7KMpkX2Zp4j0U2z5+HCF5XLIeh
DJk0qSHGPtSgxOEiogXHyZp5KOssShlwyTPKNEo3Uy2W+8FMuFqLJ0i/N54PYP5L
wOV69bBzRPy/8Hi5hEnnVrr44f2rS13nzVa8z+jFBz9+MNUyKL5DJ2Rxfww2HvfV
dfkCItHrJs5PP87xZZdXa9O3sSpYqnFCi4enpOd5CoiDweqbzJiGV3J2BdHXBTCR
gfFa6JXXlfNcS7irRsFx3DweclgbNC5J+ykZYUXppNdIdmW/UXK5NVAvITyVuGgL
S5ATCt6Y2u0gZhyoBS37YPNlna32pIGjUwLm053mNhmUOmx9mcrrFTyep5zBMjaI
7T2qW1qsF1yeNwpZNRvGKndhbj1TPkgXWUhUJX0wtZJCchjv7J3/82YbrFeNZ1jk
6NjLa1N1FaRrmpAe39ZhUzW7AI0L0H9e5jelujAv46INOsOAE5PbIYfs6YGp6/mi
Y5auppmva+O820nCANxAR5rlSNjO2LnN8YQAGrFfQZZJMakFVC2ERCb3aPL59M5R
gf0NGd+CXRAX/Unt3htwE5kbfbiDBEniOm9rjIRaZzOb2GSin5WdNw1e3MnuvhLO
zZbLL9alhzm50pn8vQpKk6j4Hc8cxMvFmhAhfXrxbwyiYsCx2m01sb5qSUXJ+O2N
fxHzsA0LJf9ZMCGIwA88TYv/U9LPtNHsDYJ+FMj+4uqxnuYGTtQLlBMWp6pY7SuR
phuTWx/XfRDR7ry0KGhh3/uv3vpLy2YZcCWWJgvhjKJXREdmdHryNEE780qfRRJp
5PigkAOHR6FdI1ot1EpYKi1+JwEzzWG/h08TWgah/251+d0cyIbGKWYjkz1iENhL
szB65MRlH2zwYk6jggIem3c7A9NsASviwXT0rizEB/vna0Wr8ObYHT0YsNb1/Jk+
NWEpT4dsAUE589/abkE9+FHLYegyOW2nSK0sfDrPpyVZeyTArTm/UWQZa4YVu+3F
BXyVuC0CXreh+rIqOA0npVCLBq+pkqJpPcY4BKVnxRuSIm2kubqKDBZ2RdG9VS+m
ARs4TfEWbHRapykizlYfazUkQghWnCLJF7UeQQSzCwaYd++Kwm/Cy8UfKJzH5CHi
Chs5AcVsU4jGjY+7IEdE0ruR47HSgEsu5l0Fpgtr0Avoo/c+CHlWo9uL2jZY9TXb
DBiNLXhPobEoPfmbYHK9cU6uhB14zAKgNlv1XTfUlo7JayimrS6Hp6l6qjqX00DH
b7UVlxRe1XD8MK+jJKg7PK23kZj0ID2aPCGM1VnDzCHxp8MVS1MytTKJhewAIKJf
sM/vXHt/5vmM9IVy6gnnCvQKEmNQX5X9gMntg/Fr9jGx/LfulaHkUV9c9d9J06rU
Lcanrzr9rIqpP/Isw2qa/85JtQW3+8FBJHnWIlRPAYX0FdVVw2Wz4rBf6UCjA10V
DgLtya+SRhStkFtInAdUAML/k+Ey9F2NY4TEH/Drp5N1qOJULM61Q/0mUWc7+rNA
zN+z750+Jdhy5wSWHQtu1tDgmsIdQfgKxLyYyjT3pLup2UpE1fDJZ3SPs2CJOWe8
IgKPAwvFlGX6Q6ZxYI/C4jL/JdviCHsdI0Au59NKrz7YtbfZM7sGaWgvbL/PC+1W
Ty4uoKR7JveDYAuBnQCHo+N7GheIR5nw/d/ajMO6ET1TupypQbBKKCpdzL0UmP1I
gURcObXZpe2Ii3ZCDPsImLmSW1rBS4o6scT7vSl6PVWyQfDByEaZje8XH2JTcGdw
+oc+JwB1OIOWC6sEeyjD8FWIn8OBn1tkCd6auXB73Qo6LOao0d0LdRS9rJKM8qXa
+PfhJtIfP9KrCx4QKvdiG7Tq7khd3La6yCQigE+FPv9v/p7ZFQlscAwravOydKr/
uD6qglq+BMv3T2g0XdF/GzbQ679DfFsl3S9O8fmfl2VY9DTY/bGjXcpSYsLSfA8t
ykTJM8eEJlQ+2i2AjgPUijPG09gUcHg8SSfHD9dgrQ53n9mI5bJNm+dVPZCxtWPz
rGpo6u8v6KaLH6P0rRiiigdxMb7giDPNlIGd2klfonB0YId9fmb7nS4zkDo2kPlp
kte8IF8w6r0DUj2X3r7i7jkku9apx1PEmZaJLj+F3rPFIa6VACY1iwWeNtdctPe/
dv0tA8vq9RlPXUYcKWyXJ8RqsDdVPkletiyIcfbquHIRNHwZgTIzQ57/rprRzt14
b8BcMB8CTXjx4necxaoEWfeHwQ1qTjn86rTV0/37uWz19Viy/3JrH97syTMuwrjG
+nv96TXvkQWGV5UGJX2cZJd1/3MH07T4qJHEvlxL24JNbY98F8nNvsoYEv6GULEP
BSG21ksp2VULMjnAazypfODPzTEoO5iwHuLOilfK3yO9jhL71RJOJclRD0Grgc8r
N7K1G4LABXsDywRQcbYH4sNuYs6wqNdn7EfwP0NDsFJjuAfhqfOyN84x1xluv9RL
YNrcQhBK1S3XgQE7WkHMbUiFNOxaQK7Djqqemfbp0yE1GV6mK2lPFW23Z2wxqxTC
oLX3TBJlGNVIFASErE2xccpDiqs9h5IuiOKC1AXmM7hK7O/UQ7feBWIECjoRVw+9
b6zAZxpwphfMbm9DqUjufcfKSez4lxh2igRSLvrReH5Obx+p6odsC/cBl5bSAzYC
JdgieNrDEqpVThq8U2u+upXP703iWpDBKxJlngXRXbpKYWp++MnWTpxRZXB2OQax
jGeejder5uVGBk4vlh5Li1H8nJWH3S2zmeRhWS1AWaTzJyHAIOp4hSq76II7cZwN
bhyGzY/kzS3Tp07avLopyih0mj1FGlsT/buZAR10WP/VnKvnzuMaEHiGznRs9kta
2xbGySdbKcnqhUvOEG8sITvEyjHT/SNZFqHVNzEOpn2ZEp/3ue9917upV1mx3wMp
gFH0NPfzNoVHrO/Ep/7E4Cg/gRcN9e6CFUNKtPKz5p6a0OEuVfFDj5F5MysW+LLq
JZgvJPeymdREtU8SYTJSlSERFbQQkF2Xe5Uc2C/Yvq+PldJX56CmCWppYHZ3QiKu
b7hBNDvnb7XKjFlf3kX9uPpRKqc2WMXLy/6v4gxr2E0eme26Hx9x4tgAOqAZ5Zy9
VrLoiE+tMHScMOv7E3lg0wwe9y4KEBdaQKs0sZtmlVhjVhJHEWTq/vc21l9pW2AG
JwlbKzDr1YX7rkwDgVNsx+TKp3ukexmYyV3gBOpRuZ6lxRIPsTfEMjsSmAR5WtCk
m7sq8sTr0dYc9dHs+tY9knanZs7bjELilizcIPkBHYgl7QR6i16ylwS/+b+nip8w
s5tY9k5v7I7fkNH5bv6ZSHrnaOYp5g90GSIo2YkmtdQpBzCfKHFqVfFOo9Q6t+5f
A1lbuBc2fZdk2A8a1EhmhsYa13QieoVEnmQpktF7yQdyNLsfWsKTbZOvBeYpdhPs
uT4dTgrUpwVW/61O9ZTsbyBviAkIi8+gOxMAROvsnyJrmcRhQs//ZewM3rwZAy32
qTHGn/pLrg/B+S+b3uljV/N91xoslnVKSK31RJrxlQri3GgU7ZJg74XB2pgL06BH
1kdWUs+SVyX3QNZKL+hqSwY02yZw6KYvbjArEb/L4Bcx5ER70oVQxxoNJC91pHeQ
NReRvVWhnXW1kmPLLZkEEG2rZiARmam/m8AP1JuxAPeXQj8hG6qLAcMePQy8LhxB
RON4Y5KXknsqpMuAENrnbQNNZIVTyRcKYAqcQNuJuT0n7gr3LB5If3UO7e38c2KN
X9ZZV7FDn6DOJlbKnKrhhPAmmhix79tsg5pqulGG0ATp50maWYwcmqdqYh0O1re6
aVeoAT5CdV+OZRnJ6sjadc0gO/voKiMW8vZNCkNkGMaiMtMIlGY2P0gMfPcuCbey
mxqvjtHC03k4Rpz7wvi0EwPpt3Sqx/Ts4eoQzmtSeJR05EcberehiQMsnQxH4/Pd
cyZySGaY8cr6Eia26cjfaOmJXZHx4KTvPPSF3OSw9UFCqkpgs3WyrZFGmjZzY0OM
Bs5u4X93uO1KBxZaj2B3zriDm0SCjWx1FAFJ51jaj0Acr3ts84USu7QI1di/o8IA
VEzRuem7suHitMcSPJXRgYaQkru8NFHe/uNNYS7p6haObOnftoQT+HK8g0qKkXM6
2sBa91ZQdUY7mvd96v1+ZvAalY+6XxVl206ndtgey6nMyJxQ6/BPSC97WotgEzO/
d5eK9e5k9UeAGY6dAQuUVORrd2Zp/r6wg/mTcTsidimoBkKHFGdHccBUsZtAWJ/M
kmlae399w7g3hSmkcaG9pU11KgYWGVcGRX6tDpNrraL1cRa2ciSwOS1BSDTEwggj
2BzFt26CDohO+GkHt3MN4q0w6tMGpad6CBNB4ltG2PMdIFuBZLBfQG82nMJEXpCk
Hh4zCXnPR55awJyd4Kjmx4lLUa70pB2jspi3k5bVNJy5g/09Kjv3UHChSb7daVEe
CTtUlukTOh5BwI0yKx6UhqwWSK0nerAGedN/Xi5TW65Tg9fMcyBnRL8LVaABEYVj
9E4pXIxXS0q0NHOb4F1db8VLWYJ5iw6gPZ4Of8QK0X7yKLMbgJZsYkP8uSCRqQx0
xDQ4Jh2BrzaC+mqyVEsDfUdkesmdRKEcWHQadc/ifFaJJKWrdWiVa8rhp/D3DqTR
sOlQRHpsL+HfdgVIJcEeMEzE9pQD0r4ocyYNqD/uFUu64G40ajMNPHwxsZohEM+9
4CVRvrRP1+Ci+qe4Yi0f5oQwa0N22JihRr/37N/9zlUDnKwsSPoypFgHvN7jDMre
Jq9xFYx3qWBRig6v8PNkYiQ006iP2/ZeYh6BaM/yeIukN5ucl9XHd7Cid2DSFR5B
1VqiYTvw8MlsRxqrzd7WkTeUTdJrFEmsi9RBu8fmxtlQYpGDVf373oTAxi94dPwh
JUqmuMDh79VCjNtUlzxkHeJznD2wgvTUC/mi9Oca+74WRGXI5jxuDl+khUIM8wHp
apJf3gzM1cnuJWVKMpFVQJ8tLguysWmkuN+yEjpBi5B8HY8H30FON12Qz5M4LxrX
TwQV7UXNu5mcmfMuqVKKRuSnRQaWkRqDl4BDcG69WElfQEKC51YfJS66qPQB0j+L
2BsOugqyO1pg08Li57qRssZQUTraOzAPe90aQ7mlykLn30HeHNJCrwTNEJwJYpYH
Vb2zkKW+1lx6ftFLB3MTB6xC0/aEcq0G1wjS6DsbEqBUZ4tZ00IvS7M7eN4+DvVC
/5PhfiDrOkN1EMMYMCdRkq3ZaQcQK2lNXKUrFaaFKBBTPIbW6INvzS1qeJ+qT1Go
jK7QHLbG2p/Jwsdm0WgSkc00B1BufdrtCHhCTldUawikpU8tnjW/XmR1+y/O1kcC
axVS4g6+sZ56oipV5rY+29Cekm4nEIpa1Erz2thhUFPSTbSw7xnIDdhHdQ7A1tH/
Wtrj15SBU3tjqsRdbeB/RX6U7Nu6FiCMIpEo//3lpTazZUfu2kagLUtJIrTwMJtN
tnwTiYXrmhvCWIuSQrkz2Vog61UiHzcKLXSRZGFql12r3+4CiXqg+wS6y5YRLb1x
8LYvyocT6N/wheKh8b2dNzGNEDwvMVcA7TUWPyHeajZLescYP21ktb55dBMNnAYB
silnkFLizLwGA6yi4CNZGih3PxDoJYcaiHX7zNPPJexzSndmneKvMzSmg1cmxMxq
uUJ3O7bajT4QiieCJd1t9lCoBYJO2hY4rRZWXpXWhj9nHCXQaQrKXzGMMRdvC+/6
Pg53eWhOnouBxIDK191nRLpMFNrmvqFHO+kmUDJ8wBoNyzoBiVJph+LZMNpFufAq
RMbPH/5UldvQG8zFJJp37ZJGYTx90XQ+3VLqUuZrAEeGA/62C+SVvi2DzeyUl9js
xLmPVH/jLxCtg18CdqSo7GcJA93ixp+PvO2QM30EaKo4ehgK81ZS4QecIO6Gr000
RS4XrbdFZTNNGV4QjnZXaLPC9KiJiN662X8mzIMEoWY/PAr8KwUApHK1IEmcKZ28
lj/nWkORu+8onGtaTQFvAFPAStO1HiLyapnjuwqwzY/AUjfCpWc5QCix572OXFVg
JUPAWiO/0SbgNUqibZdVbhVihoO/qrIq2f4WLWGC7NuFLC/4BWNdByGKCWYIxnQv
NP+KKitwn1VPV3wwI+Vgt41ZZlX6y3QZ1rCIPMy9UOv3/SqKqGAiTzVsxjeia+xP
xg6mJiWAk5k9Drpp9Av2l7la0/5J4IgRD5IuP4p701a2pU02tM6ca3ujF8BXSXKM
P9wmTT9DDvMYmKgJiH48VXvC12962wb6HApcqffHpUeu62RYSmiRmbuwCUFp7toS
BIyL1bUcYxmwlIUhiZBDEsC/GgJ7muS3h0CfJ8ZJ1nlLVWLyDb5Fk1b2cMRrFUyM
g7jiTwAXGBzUDJpFTs7BwdcIemmOyzzLxjKy9D+BbD6jMmgeS87Fkc0g3TWw5N5u
qFNUH82XZmLMeFzcb9LwR+vhwloIicswK4+CXNFnQPM4ELoM7oZGl+DWqnGwUZ7m
2yG60OU6JfBp2dgq25qj/TrarMQZebyrzMreR8RLk92+AH1qdbdmHR55FbSRuGgM
Q9yWlHXr4FPOLjHLuhFeyHNe+oEjqiiPA+0YPV6ruBmSaV7oX1GGtJNToSnGsF2I
LgMHQrWdfY3oXqVaN/HVvNHH+5nTKZMHJzcb0Yt/7Dtqa26EAnIThFHgsoEIsPs3
ak9av4kyk7+xEVnY3nnGq023uEWsL0XF5Brrcq8cNz3rk6EL2C+5opCjkKXcrEkJ
a0JQL4ZhOttHgT4FHNHPtvVwT7y4HNUouqZM19H6cBJJI4L1qf7hg0GxEAUR2G/R
+6pPx7JfNPMD2d1RXjjRyF3NFJYBOywCY2NjlzWE1o/IwPIQS5lSH/JZDuZ1dzmU
NR/oNoJBikbKN/0ga3LN+z5T3DdHPXdCYjnT94OmIFx/c6n9faAyCotX/IhZPykS
BDDV/2w1Vjnkgi5h2EBkuO13cADuksRyN125V5cxXxAWryjCM2yoM66V+5dDbdAC
gWk+xBYt0nwb8f1la3D/RQ4f6BrgUh/4RlSuB806GnpCVa6xZw0BISDumSMUOiNt
uJAZ1XJSzpD87A3mzFXRLxO2gaCEaSqH8tHbHwzn2dv5KHoyBjw32AmX4k0P4/9S
P3lZJnkZUVsPIao2hcBs2b4ivnxJNp5jHYVhbqVxcUF7qSgJMo9Ifh6Dm8+vGnIX
S0u2X+4E7pAIKIJ1Ma2U+CuazKfU7DW9fjBHSTDjYGETE6PvFImCm7NfLG6qiKKI
hz99bRO3Ktfk2E4qQS7n/ATUvtLakicVd+QycRhjzljFwyUg3KmDTCpZRaFkTax0
QqynvmfAE6oZu94W8KQC0sDu2BcZ5R/uHo3KGo1p+F/7npaUYRYZDdvP2uFZQ0dr
+JIJIrTVzLOjFfP40p3k8o7PiG1Ec9VqxVSamkuSUvoO6xGhs0ZUep9/3JLy0ZIa
YPR6NSv1G65fnuXpP9/M8I5F3U7rpBitIlcCDBhKoTjcuN4KsIWQ6JZ1JZ/a5aZq
r1cPCnptdj6BOHPmFBoIeLQf0NlRAJs8LPKl1Ip9qozIef1hxY4qeeRPnF7Lk5PF
sIkhVIOzjYw1DkHzVgMc4sAAvrnKGrHiEXVYA8QELUNt/T85Wxy3c2dwCX4cN9AC
tq7SaJ1c8B0OYWNKPbhbRVTUSIy0bqE2kqhvF4JpfK+HGbeAR52SsUGM/gra1Vca
dtZoagNpmZc77FVSPtmwU3x+GiNmLcltiTacR/NgpQtBhMx75/EHVBhDnb/GvxUR
0ox7+bY8o3TZsiX5McyGdoEIv2JaEcMPleSj3JV42T5+qnrKjpHcKqTknV0PBkHj
AyCRFl1O5zTP67XyhgCkAbDd9lia5+c4Xl5hCuJnjRpP+/G3xRJD2ThHHfMMvuDg
Xu5td6Cwfq9Mo1d/MTL9xHLeGI9zT35DvuCvEmUOsR5/yI5Wz5sKWbU6bKXL4wxQ
YzwEYQZK9fiIz1fvJ5RQZmEtSa3Tc77VWz01XdPqzPt1yVTl6WLqWNV1sn6tP7z+
KQJbzN3zV/r97P7sj6riI29hDxpHsdZX+Q0si1mW08ML3qFctSr13xyfxN61sMUS
HiXegY+QZRgiAJB59A+j8gbMw3VHQEZCty7CqRaTb9eClADemnURU1yJ4mhCbCju
aN9Uih+uFbwiuAAGJ/8yRufXTIAirro3HGPEpZAH8Qp7e8BEWRIFCxGbYRkF/gRY
cRdfawbnL7YxYx9YEYTZBj5QdGso9BNkFuaB30twRfyMrOpzsCMR9dYpamRZ1AcM
cxDd1rXt3Q1RpjFLw2xXaHr4GZbXd5iWwerimU0Qh7ZXTSSr0SeQsaAGAKWhP48U
FlGu2VwSgg9jx0cj+FefBO1ctgMP9KiFuR32o9iWRZtDvffgGBlvFfqpx0FyLNjH
XGLRMainB1ZiWah4CUqG8YKECw/SMumsJ0C0yqQtu/9Nfne93b+1JMacKxnCHaDP
jsS9DNu1Z6jdX4QWcc0e5fP/3gxFYBDQ9dNzQV7TkXFz1nPPwJl2C23/kwvxC/Ym
Xa5d8WNVyrlDt9kvox34gw2zl2q8LOl9R7JxPz4XTbS8GejWyxmYl0uXNvQrc2d+
+y3TCfMn7lJVSkrtrqW4uTAMICncvQRq3nZ6b4xP0WdXufEsR4G3AqWREykNnKfb
NRsk+rL03pCe6FaRRP5BlafzZ0WoQ9mQ1QToXJHSxiBQu0bllBSIYaYMogX9U5lf
rauKooBjkHHma46gPKvwKx13LM7IrgC0Ge+RQ6LflRLjG3Ny2z0lx0wpOMXa/tzX
JP7B1cU2aXk7Mns2kFK2BlCGS2JRIIfFDjaRDHfFfS7Af2hOkTvroyO0IQOdiUHN
GdPS08+dCb/Ues9nbKK+ifucnuIq1EwOkxqOxxMLP0PQhJkmQI6k5/k+wna6Htsa
dAMCNXLJSihyjG0M9XszHlGkcDFqV3baMi8yAmA52c0jTay6Qa+JXyFCM3H4HgMW
o767n1MvRl6i4pQSzG2yot2V/xvqPHFukLMtfmVE/VtMwFpQ2azEDFMygd8dy6ov
o9nTSIcCUWpTURlnmEOCfPYR2VZqbDF5CX8XkXD9bJfFI98eWaQpLfJLcMmo2TzE
s+b05uQmiy9Iq71i8tIFlPm1yHqY+EpaNlxYm9GHkTSPePruOlClkyHOEmv0RTks
LzHMQVs9qOXMGDjyEqDTQhzwCU13CUh9AY+udT1ATqHJn70XuYEa7uhWu7WOgQZu
2T+EYZghzAPvzQ/0jKOJWolDbonWUgQk0UrMKyGRoZooKxCVSHcqZcu4o8aRhA3+
kq6SEgkCfxgT4lb+pDy0J4OZnR+O/q6aWsParJ8Eur2wtiwtBUu7Zz7WZrCeTVVV
luA+pqquxcxQjnzRXv2wJP6TyP43VRyQutGNbyYkzGy4ZrpshET8mPJr0VaDWFGw
Nu6DvRn4W2PfzyDaoGc5C/1Hud+xXZxx6agZAI3/FgOp6Nin9HzKjMSatrqUTVGV
oE272StvLaYzfAn9PSL6yicEziYcU9MJtuCa4+o8WirZfIAiMSU7hdS5rMtNuLT6
7I79JviHgE9sa5SYz0QohE9crBt4//qGDlEZMXfevycrBfmI1uGOspGSUOlnVTeg
UJl5snFqlHX2Viw9zJQWHfv3bSCoY6tp3zcZ2jHuhbyD/Qba1ADigMj7ruMbOIIw
nMX0LHvqOypYH+AdPv3lKUlQcTmx0Z3W9WiV8bC0aF7VOVgN1T0wV/HQ82eZObI/
wZXrQaH9//mw0SgVAEwQ3aRwuNkQ+HzzPQrybXApN7crhkQP2xt/5lFmH90C7rdh
MURMIECag6ZIpeSXZ3SW8n2sgfjfQQGlx86ApICnoj1Z3L9VVL9LE/9sTETdrmMZ
39DOMS87eTgoTyzZNlUIBBHqPjjc0k1CtI43nTUhXY8o6up+m7L3eBGxEa02kbkN
GmDvmninq0VhXs7z2SqOIyRBPw8V79jyKeUngYxs0LMuDFeeg7Jz0wtdb1Y5CY+u
y3VOOSXzVKJYlcPk8nteFVtw24X4kRyXKODXDqFA3u88xu6tdgsWj5BwFBqz73On
iKKkKPeyQJoOvJR6/SfWe5JEdSBYSHCYIna/OK0H7i7SKVCG2RS4FdAforYddZI2
4leTbW+Rp3ixrSg7tKTE8jDnShKMmWc4wR+sfVk6P2ml6tJSc5fvLIcAy9jYOFfo
pwfth+cuauI0/YOF/pdeIIumeqjofx5jtwjry/FHOFvc8YTP8ECv3qnK+vJxdi9A
G3OXU3UGkAAsNQ59oY8xst1TBn4323cTFjHZHuY3DhQuz3BHh4Htylt1MOYPJlqf
0q+Cfpq1V4RiWobPCZVDd4bOjngMTvRetRUCEqSfH3aRvfNkeCWgcWW3qRSZ9y1G
LAq2FC+eINmpPH3UIZUFJvwj4cdIqpqK5u4f7O3uMDabgou71akP/C58bs+I4Gr2
WGOvjvFzPh2/UdOjPtiTWOe/mtwGZROU1EWJa1sY4SXk9PUJPvTk4sdMcmutwhQu
iLyM29m/DBs+jzNPUbbA0tcFeKuNEErUbV1OCfQ/mSpNTfidH7EANRCdzoqXC0bt
PTQpL8BD/zUXru/w/xBSi4Jci+RSObPTw0vZYLQWXNWVpKQ7nOHRG6rJYEr/VHNS
OgN/tg6eXSr11Nl/MLOthVyQN6TljouU7oFN0PkczqaRlFHFL9Bu/DprBJB0ztP2
zBwwwDCeE0FrbfbOjQu/75MDvgcR1GBChM/OlMhaNWL37YKcEjwFAsoOW6lqyAg8
QPb6eSQ7MTJ6QY1k0whNED/xMOf4D6VkSNlCGEPFe0d/UqX5943gtZfG4NThJBqX
emuQ+N4ao1E++bWG9PCSAcyBQfvOYGiWMnfZ/NJgFh2hfjH8TIJans1OGdTMIicZ
nNy3Rq7OqSFFqFAi8q+KLEKtr40MdTrm2WJG31vkWE4utZp0TO/ZYgG6lDUSlrql
Ai9hJckeoTuE3Fq07JPBvEcAYRjKKdzViF59YMmr3BAyiMFBPdMdy31Oslk+nF9S
Hpq5W1YyRIkbFK09+T/XMWrCWvKlJw51D6md/55c66JkSVW8Cu7Ks4atLqyLuksS
KEajwcG+5K7qfgxcgh8M3g15Plt+ZLJ+wDSNiIoFdHqHXyW81x9bGqqn8u/RCQLh
kjjrM3XWSfEw0SLGb6KeqjW0wkE2zlE609o7tOnzduD8tej50zR7CKIc4DWhePLY
ZGg58/FRs9lQ1gU5MQCOObXG0vHxZ/jUVikIMTMNayzCdDR8ANpEYwHQLcUfddTR
80NoePWK7Edwj7JW9uX+DTi0oo9WYkprmjQJ44joQuBsA+P2oCY6DizUZMyLmC0n
2JSRRXx5/WB0XADwd5XKXem7khdUhy0VMobtZBdR16/VcBO97ITaPmEus2iXTXkM
QpaEHzIi7l4BxUhIdVV5BHFMd19LHmyWZC2Vj6hjYDqR1pK4mtcBCIMgd5ULRBJf
zb8mgaPkyIfD2szxc4M1nHSYTQfiohnfyl/t46UgVONEX2yu5Hzz2AybghHpSQj4
qemMl1aoPiHdh10QM6BVSk0/3P7cxJdPj378ISDzHbjt7LN8xS7d75kuxZCuv6GV
mvhjN5QmCjq8pchfeYYfHsN4u9hfoSKunAV9v5HWs7FrkyPr7dYIy/+fdXjlVSSj
Ncy7YbWfOpishAjHxyyzK3XXw/n4knwI5j+UDaNxhOJ5FsAS/PptO3TZMutiwz1i
EjDynT+F4BLBllgutkwqNrprJTdUlbjbIJ0+bN54E1wv4aM8cXKzYOeIh2LO1JnH
uSvvW8VrM8LTPD7gs384Em6G9SnX6WKf1vvjUJux6oo7Us9B74twbWDp+pPK6JaV
kOOiiIHLlnYEn8M7WYQc4qN3VYMfZpnjV6n6BaYO5YMe0ezkP8QUSgjtGON8xCC4
xfXUSAC/YqGmtZ6eGTPZoyeUr/QNxjNK/SxyKcTcwr0BBccw5MQmle4E+P5G9rda
Gxpr2zOqvu85mjqxbAyt8IOVhVW9oXUdQdIQ25kBUN5nd8vkZDrtKrRFNBc5xdhj
3gZ30vc+Hz2NxseIOn1u/zXO7SaAi647Bx06BN/DEE+F+M4TxqJVO7Tdk2DbxAn8
WTIHZFMdyG4Y5RSbad07innhlUtWACXw+9eYd8EgeYdim1HT7y8/A9PWBH8i/aHE
rHgFiceISyvfPmnHvDTRX3E1MQz6RbbW3XKTokHNio0sjhf2hqVjxAC/DSetVwNE
udTejfAcsnvIqUEI5ECJ0OY075SEbDlJnv/HnQpKH3eds6qgv5LglgXl0lxyII7p
vAa/CXBz/nLsI4JmqsPZUJ3+2jj5FCDJ2KPGz3E53KH2dU54Fk3GEOx7dQvG7N2b
ToIinkHfNdHHVNoRS70LkAph4y7dhjqLR79gJCBN9SMAkwDS3T2DY6TkFtN9GGHS
8Z871aUSO6MR6/1i7nPmrTnnRkoSaXD/seNdNcrxkdmLpJeUsCiUK9vtuL3tJHN3
PcEmI0Tzi5CQiswnsmAfZvo9jSHpjJkPfvdEDYaTvRAVitmT+cmtUFnxzCwUv0rA
4xO8qJTB4eto13JA9mHbE4AT6GXjAp91n7pVP4qttANCALZxK57R1Qysc9BmfRtE
a0UGmZTR/9OVXjkUlXfiREwRAe24TmPFplu/ckQ7vXOWUi9byHlg6AXCxqLFstmK
UW/W5PCjsTHKemKpXd/XByd7VjtV4lbM3EOtCsc7tOTyDoULeMfuzwwAf+5fTIfW
v6gHbIsu5vPIN96jLIIe2qHgQkrEJDJKf8mp7V7YCdESK/L/Yo+UHDQOVUfBdb9M
LMc1BMz0UefgeSMOVzOzFXb8m3y5AkXv/NkZK+inMMQQlNuIkV5tM1M3NhQTA0l6
t0BwheydOTZVw5TZn2MoVkXbGafeUlucX/QGvMex2rAAGQM7c4aWpUbrzynaqmsv
0PS+CWIbYgRfA6kC2uwc5+P5EfKXp2YEvllOGgEFlPLtwLEtkVo4J/MOs6eQwueJ
KLo9Qx9KzlY8uULr4JcxQHA6Hz6s8V0m2N4SEHMWGmdbbpyphOtdgko7mz30wpLY
jUgtoIdDd14oawghyWsdbb0XKivAn/kVjMli/3OEWE+SiNXKHe0SSGIcE8ItG6Ht
x4I9SOMN9q6bbdDRC/zQo5XpyNs8MGedGF65R9sseLXtb4nBG86pH73XkKAx2cmt
5O0YJ0JwBbW8aH8RjxYEC0AP5hRLM41j0NYV3NLRvkuhcq56wV+WUUL1gVag7LtJ
jb6NuvDORojqBXU+H6ujWHW2jNGjgmftNQpChUnNyX0LrPAm6QK32MbLATjYwOBw
L/5JUvUv/xOYmYrOarN5JpOLJY8Cma2ws6wRYUiYPUMpodRebr8QMq9pxyM2BPqh
okiT+c9IudMbWM8At5ZxrmTrIC31mjm8mFiNYEUJsutQEnEu8zjFGIAk9aox0o3/
mavIIRRH6p/q4r6ovSe9VhlvpR5comFsBE/exKWUj3rcXwSQATHTOjx+tIfNoJ1C
yRpqGIX9Jxzdxq0yISsh9cUJWQiv4vBqco9oJJie2B5+FuXRGwjXMIMxXUX6unwQ
xrhH+3lVLtAPdiNzVB87hbHY+KRMAuiMp6bcP9FMNYcpZ9vkKD1ZLhBUcqX7DSKo
FfXDMQ8L8t2Pd/XeQj+WZLy0CO2W87zxoDdcT857VRzRfChAnwW9saNZ3cextDt1
GTb7JYKLIHUEZeZ90haYdHW32d6bSMk+GUgI2IgV8VgTGDdBtmOYD/7hnXlvP2cV
ksMSpyxBgghGDcnUHiZ39JLQrAiuM4nBv4bkKOjMB6jTF0gQbx+WI+frWzI93jzh
xxEiYf7Y7OMygsijc90y+lmJS+1uhp6ghH89xZhQhFic0vDXbRXaxgZibvLH7taJ
+lZqBLlCsXdgTTLdvPfBt57DCIPaCIaZOgTNCjg291tjWi0rdzvi0BkzvxyylaaG
jkvZXlkjf7wFAXj/+uhdkWhMrWDJRzxqBJbHr5p0wjwZJSryt6aND+Iw8p4z2A00
QDYcQONMT7Xlq79+BagPGTg7Ah/Ubmg4uSqafPF5u8aBHqHz+1wbtEMGMWQTPPK5
71wp7jAyc5OOghd/x1tsWAKPioTpDnublZaWy00djzxLdxaLLbPJJtdogpPig4Dj
RgHAm/wz28HThO1fGrTORRD48qMZxPINWVZkNuGBj6C93Vqmi/gUdzkgnjVv0BEI
HXef+GdiPyDrY3tMx1j0n8pQguSKP9bFXmkrOTn9T74oj7Z7kgLkg1eib54bW3hH
+nbI81m28lLrA3I6rrYLIiFngVmsbOEB29x/7i0qwUAdUUUaG162Hq/AfUAEkKpe
t1ohoPGX5Ox9c+XYJ5+LOWD8frdAi3kws+hfSo1xYe9cOtOO0oqIdoo6Jr3QBEvl
pun5AkfkiAW3o5Kh6Q4Smr+tFn8pUz9//zkMi8GpTFKPX1hVV7Gn9vJmQOLDUrer
wKLmLCODGrIv8LCnJtA5VXXt0H/Z9Sf2Utb2BHnUKNaoS+/S063a9kyyqBt8ao8P
jW+ZMea1CIdkAPi1fo4CpF65nTpu9klsl0ZJsNfaYypgWkIckjqBz2ewgYS58aBA
Dh+2R8179bie9WYhrhYirSLT4XDbnB1L3ZEKesSeguVNlmYOZLxTJytZmWU5CKKm
SLGYBA6K2Fno/9nQKLHR6tjyS8un5+eRTP0PS7dAkzNVDvzuSEOSZ/FbIFkslAhx
bDmSfuVNjOuX6uCH4mPzMzEVxFon9Zz5opfVQH9/MMBf1+dXxZjGaNsJ9GsXubr/
G6F1BMK0BPp83ywZ5eRL9Ny0Trh6k2Ml7K85HlLM6P6XDb5QRzYFDDNzLsT+sTE+
6sLk8Ni7aLvoL9G722hMu/b42qRW4ee8HFZbY3cWSBLVy02Je1740cUZCXJuztPt
J4bVlaLWps9SxBg5PHBpcT9zwsDa20RgbWBDYFk0yMtwj/wQVC4kfBLP/i9oFTxk
QS2lCVmTRsVkJKJcnBgWFTPfO1skTg4MAJn/LQsCVff8t0dtW+pDKbAup8CuI/iI
j9FVM0NuDPYV0Q0jKyl2l+FCV2nfbNkknXx/UnWPTYSnJYU2iADe7F3By9V3d9Vi
pztxmxkxD/uvlopddSXS1+LZnuVViAPbStT0NlKWwMPf78eIrQMtPE/Z30QS5sXz
6ppuMksmSyi9P0kvu6+lnGxGGRP7468y/VGc0XgaTJHT9b4YTu/zrrUNUwYYjXHj
FcupoKs3v5yrtTAodAvSR95sK/WHtB5Ihp6T2TgsgDdmp+Nr+HWmStQTyJ3PrIFB
h1rx87j/cJevRAHq9pvTXjGd0+mt6and/ekj0jOdU4H+D994xyNjakFDcRGSkg9c
NILRdIFcAx4kSpBxYQucjzBdj+Pqv2eyFepHcT5qfkUxJm7QG/sEZ30yI40gXIUX
hgIbNVc8FCpbsV3vhhZzus4WyUDoCkJFdweh4JJgu5V7YN2C5KzFEo1vxnESkwx6
TouKW9a0XTzrz6MPWvl+CpRcCq8LSFyW/qYvq6qUV01jJd++NxxpmeAMpoJom3SS
NV5Nb4fh0EMqyttn07MU49z3K079dUHWtDZ26FYz0jUktrMYXLaibcH60OdVDCBU
bUd7FfVfIuey6C2OED1NptHXbWa5wiqiuVgP45QRxzBNi5u72OxTDpRA7ezIoIjv
TcE9uaNNt5omDUPXZ+bbF9XeXQW06E3bm+kAspZJO4F/z60+lKTGg98HBvHLNZMK
4VTOZO5/GI9elnV3Mok+joD6/qb89sVWFT8PcbH0Y+5YI9MYrtLQFaa/9a7b1H+e
mGtuYfyKoMZ4eJac5O4e4VXBKAEpOdiQZ6kwtbBSTzClfStQQ78omRyExwSo4Enh
8+O+g0PY8HxaPzvxYlzz20aecY3+biiUW+YCZfbrGLJufxA6vRVkUXe+JtyUHW35
owEGi0+Cyl8hHS7dWRpN8XjS6W8gBE7gzJDbqmM9vA5BCbk3UM4Jh9uHXSA9FPik
48KORnjpAPED9FtZF4bcmWRy8AlDrPtMTWbHkwl8fa3byBECm0anSFLnTiAIESyD
I1AASuNMNt/TL45UmeqnYlCA8zMqUeYKklPXno7KZvQ9wQlEcJh6eiAw/ruLn81P
WPN6nv7eeKtM8nUgaeU59mwVBj7cJ54dRskn2ZehqqGqFxytvwtPJWeMbvxlZMxJ
ZRZykiwoXeuzkBQhXR21pxcuGP7rOhyvN8p9dZsq1uzYLySY+newG5dPvCcSzzvQ
FkZOAKN+ijDUZVrR7pMHW0dwzC/dCCOHoHj5APsEjcV1ftcMhZoDj4ssM7iNTlQ6
jAcrVLnEj7T3eqcWE2qKjGt1tKEY1G3j2RnZR3eVm+PuNdFL71y61IOifxIFi3mH
5YGgbSEeo8tN0KGLnsZKTvQ09FyGSmnQSDQfI/haqiwmsjpHPS+M65WdhTJdeJPK
CeHtwAasO1W941wxX4EUkDcGZGAhm+DcI2b1pbBx6Kt6f8Q068rZDWvBTk34Fm+v
htGtvW1/YCUPHJqT42KMEEfSz7qDlBqd1xguVzlM/YkxyMCEXKlPbkJgiihEoZL9
MPiR3+zu7JiSfuBz4/7I0EdfwQJmjU8cE9XOyCL4SnYhdwZw3e8+cPhqhuYgZvo5
6CHekNcJzyId3V11VaWp53sdXtEpJgXVG6ASwf2uT9hLvUGOFSKGUR2l4htJubxf
8NVxMkAx51fA+i831VpB/RBPMJ2NN5R1OQ0K3AdPx9qnHYkQDmq95NbvM7SNL8in
8Mu/3u/g16kLVXIB2DMWX1tmMCx8BpkLRrU+5DBrQuQPyisPprFALUd6YFFZweVX
nYdR4OyGwpPJemR5NKDXfl2LCURbGljha2v3U63KJcMShF4ShCj3vDoGgOHwNvsQ
1EpSG+Yj8JkIi2I1YaPpdcWj5/hg2n79SrEDauRIT2uA6/idmrUb33JMdjen3Dpy
iNDvinnAhTRIO3xzuv/c+h23V10ppiHicCgWkvjumD6icgyzjEi197Zq4Svy88Z9
WHzu+S40Gs23a5c75LuWKsM2By8fM1WUKapUtKAy0NuPjYyHkmCjY98mQnaNFx2j
9zW2AgvR8HxLq1ch8vjsBDRjRjF7X4fq8/7ex7AjsSh2p4/cA+ddmonFVEyl0Nmd
2ziDQo+bs9cqfMoUpWeitSgRa8n1ofrTSa44DluoZwpAUDwt5L3ovHvH2pv27WDu
tNWSPaplWIDoGOi/P8LlbMn2UQNGJRG0kKCYPpkRWV0NkAaFEiDj5nAJH/Z9TJFJ
MHHSp/B3lz3W044j4rYX7oEe3CdYpox3QaBCU6QCyLzkD3egWovi1TryWoIYTErA
5Q4xtaPYXY3ionhGwFAU5+TkIWzMVz6BxbN9z6DxJd8IVqF3GmSfZpNvR/OwQ5kW
P+IgUbI9FZ4QCU1/J1sVGtXjpJNxFhyg1w5I8WraScgCr88cQ642a8NLlIow4Rre
Px61fshHrKloaBRHKtEuuDaA/wUBafnq1V3SLH/S+uYNkS4H11ZlFRwi73vAixpF
EIcVdNki0dIHzsIAl7gm+ENAzkbCIPjkHResvDm5gGjIr4mPaCRzZ4ppbZxd6WJz
E2KMThkvZQTwOCTTEzwPAg4pWLxyXm/bfh9W/zYvbsqtZmsGkm5BdmpsT+2fOxGE
dgTqB/UghRSB/QiY2Z8qHrY1tH1FXFv9boaWrR7Y95iJai6QrpE31FuFis5x/qLm
iRdUPqz8IYjNPyblt/wcR8lGhrnL8n8rolYEG4HS+TW1vfMKHDc4n0/pBlPzT8lU
cvmcazqNCbKDBBwlTf3JBkKTBW/mVlLWkeWHIxF0tSIsAAtzYgMcnA8XUed7eSfQ
QRfvj/zfhOd3/A6yCDi6FYnEWpGLt5gfyC+6pyH0xWZ8tfsUfQu3KK8H87Aiq6Cd
oYsJFk8mmF7CdIOrQr7rFpYjHg0hsc2OrKTPQQ1hC6PFcUROfh6USFjjJyGe1KJi
P2+iiNt3z3U/P832CnCTAfI0MlS2TfiKzPje6oVmrXD81ZDCxA/gFU545SGElGnS
pN1qotafmB2R330sn7rbUI1kRtZYjDjJz2BWbJcV/Vcjg7C2Nt0Bfk1sYAsip8QV
6QR9/z1P8clwEBXO2GGN6V7lfEdwc+ZlUTBEFNelX5mu4eJjsO/wRct3kfdF2BDR
UP/G3Kvvph/rwr5qrUMSwWo+Eo/wv5ymtq0SwC2jg7RpYVT1aZioQ0oKNXcF6zjg
o+g/6l3JwMPHJFRCgTgC1QfM5drrpLtmfIBMjZgk8Xxf/InFZlM8h3sj3ZLJmZjK
BxzB5/rzZmRTfb94ochpzp9sOvYjW0sJSNcHElYNJTOUtnSvt+f3D/oYBfwBcZXj
hvojW/zD7WRlhfGPs7lKMaOcFdeiyJkV0Nxs8haKISvV0tEuL3/h82pr4hofJo1g
/I0dLpUY5vjtH3x1AjfowY/dSXnUOlbt0HJBiJxtGAfZwfkgMLi88r+t0r84brIl
yJJgN6ksRVH3EviiHHbqDN7Rj/wJEkdSozvDi3t/jtogxmE+eebBsom97CySz+k1
Psr2QX/XWr5Q0I/gUg3E1AI/Dy4u/yRtRByW7wZyB3n8MMnOdm8qLzKfJqz8FStj
G3QXiVWpcLgMf1OSIQksygbDDXPu6gWAep75shlL7mmN0NSkB6NK53KsIstbERrZ
eZvCk8ToTc+OkUBHric2xQeJPQyGgx6t/QsqSUTPitsn1ky2drSZteZYeB7h7Shr
Jr6ZoldC9sFmpdUyIKpinoHyOu/tYgAezkzmF07AEKPpQd1+O6lUoeqW+mVhEBcr
uUFnyVv4MAK1kU/yo3ECQEJ/g5iaZ2Et53dJjLXfiZmqvpSqYcYtnefc6wY7jpeQ
38gZeA65K2w0+OLoWdwlmIhBekhXMl4tULLsUPaayH/a3zOJ2tWwrIXdX6gzpp/E
ZdrN4nzJT+jx9JHbKHRm7mWd2QD2Fu2Jbvj1VtwEZaE+Q2P7SaSPkusNBFGoZmA9
sM3C45eSCxkJpA1EF5F8UVF7sRAbsOIkKjpG1Q7Wgfxzj5VFQ6suYY8BrhGK4x6D
Aal2fNlnoNhC8B9V0Li9xYM8fAihepmXF1iXeDxrn+5tc0M8Zeej3qIXUcnK3Jhh
kTfgeOeH71KE+Eb9bAn0yrbIp4uYrUzQsJRcrHyOtfJMOJQxe99S0dl3YvWFitLN
8sFyUCp6h6T0wX4ng1C1cr/Y6ppGwU9MCqxQh35AnrW33D3eFNulK1VMZ1xzfVwM
tDpH2YBlnUZXGQcR6F7vgNiuje9msSOzZBtSYT/FXMYvEzEQxiv0RVtdjVwfXOg0
hD/b6NKGMv/q55Kdjywqy/o5gTiuCr6ecvQfJT82Ai7i9NbCa3Y+t8A1uqFpFVgq
ggxTII1aU5aPD6pEI9b0VxK171sBBUvGedlaZ6y9sF5Lzy/WmoySb946fdpbo5bN
W0d5f2pDDCNBZ/4Z0TcnwVAEj7MyIRhUdt8QkMIo00H9HfF5+OVhQJE8UiEMafHw
Fe/D+7/GMBRigg6w+mNovr9U30pG2cBzOpuW5g5628AyNKXgn4YsiW2R1l2g1SNA
TsqzlWCUE/YI1Jat32i3nULlYbPZZ5KGyNw4PW3OVIPEP2MFcVelsLRGG1+99eDm
YauBNCTn7Z77xCH5wbFQ90bNs3+5hlCdE+kygCCAPlbUEVWJIvE0+x7su5Zzs275
7BpEztm9JfkBOVc+WjMMMbJv/jzrjjH7l7lysG1ImWCRtSASdJOK2H5UaHsP2f/W
HkZMDPQ6qyzLtp1RO7i3us0+mUJwqtHqMdIujc9aSgf5mdYt4kRQ6utVZIgySPhi
wBxwStTgatn/4v7bxYhZJVkKvDmvafCfEExVYMDWK7ynPmOX6bEnBbxMHE8MB7OK
h8fXHLPQd4egmCtSR91QejZw2idSoKvMvUnjSisx4hIGUPFslz8oLvJMthV7rK9k
6/sCCsrxz2cSbLfJQrgqTow821vVQs1uoPUfeR4MT5nNJnguSvyaqXhyqUNNH2l2
7hUBbghybcJilgeJEUej82Nz7cuVhySZRB1XfmWZFgGuenyuRhNXbiu16CHFDVLa
0azLT7ohpU37TuhOY6PM7qnfeRHPPM4mhyDK17V29TT86KYJMupcEcrKqtzxbotv
y5laEqtsierSfK3ET4Twmw7p0hBRnZbZSKD0xXdEtJBkUbBOJFpII+Jju+RhDLTj
U+W7Up+hdlJQyBtoomYtw5Ga0+DRMFcZKGoC6zqGzb3WyUP/3s6Mb6VXhAg3F2pU
eRKVxi/+kyfy3sRRP2wgIri7it04PiAQo7gsFgT/U0lifnsp3nvfNmsem03PwpKA
15U4zhEiPzlum08tMBlUiOmpu+xmWrb9oCx8l0eY+o5FfdZd5ydkjAoNI67XBt7T
rSy1mppLJkrp5pFIoZJ1O2Q93rbagaOBLACp2S/umIDQGQz4yPqd8UtKlnhxIwPM
3W3fx1iCJhXzDAN+jPGJnEe0AaxqhPsyWlMBb1mZummfdmjKFDHy3799HvJROYZV
FUJN2Axxxt4O8inX+SWahESlcbuWzU4sshrlCN6DhOoWwVpac19nWnG9d7br0JzH
pyIUwZrXbgSG+U4oEDLfU0RVkVPWEaRkHP6qMeMNYTQE2n6710n40YU71I+r85H6
mRZnybLo9M0WYMnUuiBArMm3xpGD7ukm+Kwm5UGSWAf1iuCouYgzfOMLHCGNpDFw
5Z0sIQY4dMGxBGOpRQcYqDCxkZT6DKRnMAtSM+mp/UezTICl1mB5drBCII68VXRy
hJoFNiJ+2Xy8/k55Ta35xe5EGSUFzQCZfWTCPjW3Oq6MqyzPO9QbFxDFQKPwI8es
N5Wx0OBNzhMU8rOGUS3OHXfHviHxWtZ0j8iHq1ij6+JFfWtr9gvHEDGseAO0i8UE
msPbBpv0A0bKBAiwwLK44tV7gqLdnTtVcfu8GE7CjM4XDeg+NbIDMdxXe+muQZCA
kQPHsaf2bK2xBPQbwZFrmNe0z7N4YT2Li3JU6dG26dW4zke6oynTzhCIFKBkIbAc
KcbhAOP22yaoaFJYn2vn5Mi2P2UuF9AJe+nQRM/z1logQ8kexoWSWd5ydrgdrf92
kE3zrdU1B1aM/YKuAf+HLmJmQ96cFcKKNFkYUYLnprwCNHaYh5Q3vyWaUhXcPLIT
qOBL5n8F1SGUBoqthhkBM173rXPEtq2bldkMzuemGb9C1aHpDOAk5a9GRDOJS/mE
xpz2K1BTErGPb8JmVLNz5m0TjijdJspMIkRWGndevFnQTxmoPZIQuQgzMqTDTcBv
8imE37uet8s95lq28R3hnZeY2lYTzxd3eI1JtPto7p2S00QQIfpmJE95RMAIURc2
bJHfFPMW8eyOzkyl6iCQ00t2eNcpvMGcYQWBCLyHFjbFc9ECvlST72+mPbzuZbB/
ylMX0EW4sSSgjvP0yY5/OFUSWNtiSw8F9hNmImg5Xm4UGMV7iyUX6r2vmsoymB8p
OvE+CFUqTqTfhkLm+IrPSD63WJuSHQeks6X8hAbzsQ/ckW7Vt0cbdwHxA8rt2XLD
tpLg0ZyEq4JitLstHm7bMVm/cooAtv+b6j9DSxm8TbobhLQFt8Yf5ol37tQRNJPN
O3CqF/EneuK947atalwMaoMtXkmM1reoZZtTo7J6BT1XnMArrYexVcJv7lfSs2fU
C/Qt1PZ4YHWcjmXztY3qarjJn5gZQDvseIaNEd/Qjshwo5d7+91MBTxM1OIEHQpt
Mgbg6+sTet5bbsl9tfhj2LgGNeN3Maw+tC9O8Ydteb/K0oO0PFvQL0npP5OLkByI
DvZk2BD0SzHQpaQSw/TFVfF82kL7Ly068MC48s+8UnnnnVlhSpFBQwEigZk1c+et
DBrZpANyr3dz4kwkOQMTeT3m6WIoxv+SGNvDeHrNKABmBH3Fut7UlQBJOtAGxex5
UIGo1AANq3RxubyAyZtOmaibOXYeLdfp2Z/dh+RxazFh+naZoQ4Wh2ydfSeLjpyr
iw0roNOCjbNJv7hRnDu7kXmuSEgwS0TpJDIZzF2x7+SKSvaUbScrr1qxrzNCmf+c
bzk70rIZtDUTv7IlMc+PZiwnl8VxB6UTetwlXqH/E3vcgu4TUj6edJ3jw5mZvpYn
zcv+EezaB3YCppfd6qc5dSnIpJUWMQWOyi3NPcfGnqbLQTPujJb6DsIfIX6dP+4J
wKkeATVdqV8ucqMQ21nSplbR8Sl7RJsdlJ+eWQtUkaq+tjYsG3F9wKwq+c2KDarH
/7TJiiOkoqEWA/g9oYIgazYruXkP+TZgFqWWK3s4fsMFIBFRxwPy3fxsH+jR6US9
UJazEDYmB24aeoa4G4MDoHWuHGglm2WbxUmVp3v7GkrIw8LI7464JqrMIen0fNwy
Y2ChuvI0xQ99BiKpSib5lMiu3B23F0MBgauLZrlB9DXVnNh/FahqwJZG6MnQu1Jk
QIXj3mrYxDpoQYcfMiZFlAg8H/oSAV1Bq1CCixBMuDJfNeV8QHLOyox9vUXHDY3S
82CuWY5Hu3BqYPR4Bq8X7hTo4AZYbAwdQEa2pHsgmekI0LC5+rQEmA74eE+YlUBY
10llrUGEQSQ6Zb35EterYKH0cKYnf22hXS5mRYPgb+tRMuGt8ujBLZ5S4SmL0VXS
6lW0Q3ItZzJOV/eVJV2916kKxMABM3uwWwDUxQ/efX/a4qYvPRhA26efbT421Umh
rMg1HpMZTH0ltEFPconRaVEffCkQbBgOhO3do6TtY5AK8mKvYUyvmbDDjQaPOFeT
tWrIkNso3aG+BYKsZ5zpDEfu+Vx241oeC9pljoQ2s4dSl3bviAi6aouQvno4j4hf
lrZXiGI74PgGcVcKeH6X3Vk7v1xbbrFN2ecO/JxYUxQTxQd5mWEoZP/gnvIvoK3Y
IYUyujXS1n98xtk/Qz4LiXQeNN+gFeE+OcLXtg9c1xyZpPM87jmtie3wMYJLpBdg
hI5tIVlcFKicFUHwaFRSFKTVljl8NkjeKkvdD39mYw7IGF0kJ12eXBQxUbYa2Avm
nKpNvhzzt2wFKXjsvIA/r5RSmKZ0eoxfhVrfIanOJ/TdGY4AXpVOxOszFHRQcVWH
0N7+Q78lKePOU1/1Coc0BTsFQ+L2TKmv9VHBWHdYn6NjoHPkfs6abm26TI1LwV4/
w+jqoOyj2el5JjIyM+w4sgs8uN9M52bQGBG2n/s7xUcd8XyG4Cm42E2G8nnq6cUi
12ROVW4YEDs1TnqTbDa1pEoqHR5j6M86Idn5cyl4zjkJlUsXYhNecf1uY7VpfwV8
NwKqqGHEiBbd+/Hc8xHcipkiPpxcbdCd3Pcj5aJLXr1EXebRcyA0r+iuzgdx4NJL
X6eINyoeGtaucwYdDs4jyBP4Cda1VcGXpDnBfRD7Y3p3ME5UpBHKbkaTJeaN1VsS
sfITQIyKGrpiuzzAYU5gUxjSHubNxNXgJC1tS8cw6+DjP3c7nCfj8DyBk1H0X5CA
C8UZaseVaO0p0Zsq1z0x5BkEgAeq7CGfMoSAC343uUlMRqrmeBHUgDYvxcLPP4Fw
UHqMlXava9b9O4t8/ocwzgzKb1vTrJPJGYNHg7kyd3J3hMlHTLgRUVcmFUxx+73L
LgLAUC5El2P9zdwKiLBD1OJNG7a37tqHfU2Z8L8ZVELjCmIk/d6JDXibujvTMFRm
35r6goIEY+a1eoXCWkkZoz3kXcEwpEvAfIm3PnaZdPuNsnHLRSUfmCHzGhSOUAHX
L+roCE+dVPR0IJ3VoDwyV5IcuKQAdY/xVRD1+oQT4//X49mc5QPyLotRFveEvWaW
/PKp7VqiSYc46b59NM7KTu18lqlZ9t20O7xNaYicgmPAyKRvO2zUukTQ/vY9BW4p
+o1I0k+xviuwfT79pjpiEIFH1mMTr1reeIMtlEVOSkLNL0/CSBWeGD+3yp1ktLRN
oNAuGcOtrhh3LjQosgdgL/g8qpbXEN9C3DEkEhVe9/6RpYHNWAhAnZyUzN7AQSs5
AOh15nJZnsZMqrrLJn0mn9xxtOEECWmnZd/kW0UPgAXhHU37boNqrCtvpWDwKyva
VhYzDd6rQV0FXTmlovSHxWQuNdliA3PliU8/OpW2HDzvx1kdg9J2xmgc9+YQsSPB
09ER9Zx6QwaniREV9yw+6mxwhp63xbigXqgQTmsyCL4hkQ8OA+Ywzc2pej5GL8Zq
yx+BC1GvbaqMV97brwwWc0u9qUhxlcqGWkd2aDTQJjFuiqLbsXoZEU7GnWM1smFz
I8jKdHjf+otCcjMaJ5AmsA+at7ESs2KVqBgF7hL8ROq5/MKoXqKa5TjKL6SPvoBs
gqwWg6v5HrOsg8pj/eMCcbG0z+NdAuHttsKp9edFdtJt9uU103ww6cQ06yYw7/ea
mrGXOmFvafaaVuoKsJsq9B40kP9+GGxyk+5AA5pbDsFoHiaHB50/AI4sQtdeI0ZP
/k+d1YMuLbg/IJanKGokJSm37VwfpgUdxxxC1lwN4yWHEhrSUAz1/Qj2NV3DgKMn
ZFR+ltCe2UjzpmS602ro89CY6yOL8U71poqusGXvdXb6NOjGtSwY/EESP3kaDwvE
55Trfhleay3pSca8ysKwP/EN8MO1De1ePmL566BUurcZ6TIqcJ0MdZ+ZbDYt99TV
xrT3iY1e/mzvuyQkFuVZGMJMO38l++SuvEUPItiYwBzh8j7/Y+SjOUzEp6d9uX/Y
8bamAF2ShYHocaXpaVefvlJe/7DrgQjHZGEbKxi7m45D0TFToVMR/0D+cbQh+7rk
9AdsAN+xpWiMzLELoS3WJ6KRY0j8N30kpdlDl72ZWvFNowPe72LTMIspZuhS/bcJ
lCJV9vN+IHl69FZCIbRT69jCai9Xsd4EhhgBP25eAkn1Pp5GKqAau0l7Io7cBZAq
5WiPyD8BOKAxp2rgD5lo+U7GnzkBh+qurxCXgBK8Y9e3c//OTrUyZMQXXTYSGLZ2
LuMjunFxjcsYw0fukaM6FdI1Tz+IIPMBkdbQiXVoQhgU7YWGnfAWIB1VljSLOrDX
c9C6Clp4tPB1/FEmz/qlHNWbosuQnsrBu4PHS+KDVQ+dfMz82TQ1vjJpgI3b8T52
V0eTMpMQO3ghAaYoQFMk6IHUnlSsoAV+YfBkWJWnVU50KFHhu8mZvJFfywIuoANw
oud9U2Ud4uYHTkugTuszpPiHgPPsHSQitKXXUMEdjFbFo+PU6hKf9LidWPVAkzRF
V6aQgGtNbkZ8h6XM6DaS11QHBVYwE+PCJJ4ToW6fQRVOsfea1g1ZjwPne068Z/y1
Qb+3xdaKO4/Csmxdqr51nP3QRDID0xz85L+tP8NmxGYjRL1iIz4cux26r3/PaydO
mN9QAI4pKsgEl/vBgkPP6QUHsQBXGuLOV/p7A90mE+LvhEgsSeKd+JLj6Np07DTP
WZCsG6TmV8V5BrqOb5fr9cfmCeWA+CN9TqY/iLzystms8i6In29QcLaIzkG6yVth
qLtsx6tZgdetUotNjlqqWG9VXdO1oU+WgcH/J981eJfPmPSW+onnIfZFrKz+huBb
ODVgxOEtlyHAyhtx7nrMd+/epEuummWUak4B+IxNohPmhDCN17qDg1LFLgtexRX3
fd+Gbev4TQU4uEVTE3q5AZzmfRQizNJQ5qCwwnLf13FKNyrKXyq31zYUyV59Thve
NwMQsP8jEL8id2nxvccPaHCV1BBzoe062cp5AWF4meWI/VmUafoCjENqvI8k47qZ
qnH0oxVmVRnNrfrEHrEppNBbmg11+GPFtByTos1LPo1/QAXm0bD/6cUZrEBvHvtZ
xUjvABv28vcbkmq3g3F3Lz+zwYeXjCjj5slT+Jh4UzpE6JLFGduhc2LDR7s0zUac
leIzUR3qYax2KLYpH9brLM2NxybMhTE807XdFup6T+PiXS4ROftg2LQKIE1Xkl7K
LG3L12jjrDab7ndiqR0q3dgsdtangJefx7R0M7PiqfhNvwU7OiIiQsSUe6mHvvW7
j1i1eJCjs52zlo3wQTEc+lS8BBsQUMH42e0MG1YFTOiTS6Sy+36HSQOhxlY0fXqj
nb7ir6VRIuKMmHHyjhoGd0ICLhJs7Klrq2RxzPsfee2pdtJ9x1B4EbIwhb7K2jSm
ejFhQR2zziy0z3zRIPZlawKP4mdZIzhkv6N4IbhFUdgiGs/JQpK6pNa0SCQdMZdH
zlKh3UhE2d4KZHOdDn9EmXDd84mEQ4S43hvbNxgHhgHf6NmNZvK9SicaP4AMRM9l
NHH3ETLHYmcRu3yHhTT+aPkoEuD9/BpzPf0hWb8UXK+U5bVB32WL2SUCbM7pl3Kv
XIVW9bDRcIGUBluaAw4moHIHFjIgPPphOyaEKtxv7w0x9N9vwfDbC75BvbNMlp8F
/5LqHiVdDvf3a25+beBGuWUg5VE6XL0xXpP89SQIZSkufZmO9FFWdKs0/MD+LJu7
sEZDUi/goJOJrePKWpu2lQXyOpWftTBGl2yCrvhTo3a25L1pxnJyeb22ozWYxXh0
qwYbN1Ip4YPkiP80PW17LmYj1zH5c4p9Z72Ck0MPBZpZODfLPYQZlD3PGZ7I0Wk+
OmWlEMBHoO4E26T9Oi3rlDjmXQ3hdrrqAQzcKfYOznKZeJuqWm0iYeXQtLkRRkHM
AnBA6FAfAbJNfNdrIReSTi0/xxTYMRQA+mnD8rLJsFtQfHkkpdCs5kO9poIcyQwe
7kDUnqV5InVB7HSJPEQLHNHnEnxZNjfvAJissRhFimeu4nngqqQY4LMGOsYiAeGy
BZbYHT3upC9yYwJV5wp/aImTgrLnLgza4HXWT52D18aATrVAWA5ClWbMK3hkjukT
1PopfBa9o6rY5EriMtLnB2cLt5RPDL/va6gfQroFBMS7ZWxjVuFtf7w+M5baDdWq
Brn5+XN8dMjq0MPKEJXeaWLllxTXyV4AtPgNe9Xd9VgBOn9wNmfL0o1vz9SYcrgH
sDfdiIDJpnIfIVlgb9ga5VZpKtw1iGp4NJwiP1bMpqAIREwSYe4ZPcyIIxCyUhfb
wVQA0C5MU/4jVA8wUQgJdzAE27gDE+okpoi0p64wHxBBzv69lKPQF1gLDXycLQVD
nFEkv/gWYNadws6FzMNjNwjkX0Ul11eMmfqGjo8jm6f+hdOyxpEnTERqOmGXUjHT
nr4zYp2e8PRmkbZlxIJGSddL0v0MSX6SGU1JKurOJ2IdYI0lv87TXTnjJp8UjiDg
ocy9bm8Pj0AzYzfcO/wUVQYeruq8iLfmxHFZ+HZopWvTsOe+2Nv8ZfNc/gh1/2L6
IpURvOavyJdVGfofhzxfN4My2uB0OpMD+Q9KB2dZbL7r0NHv2CTnPkuG1WYGOp1x
Gpv7/v0jaxZiWEkntUPrKzUb9n+olpAUo72ryTC3VJyMDOxiyJLDbfFDodY+PNrJ
ML0XVlMVM8nkEk1iYIC1nB7F7qhRl8pw613LH8y9NBWaJqaF3978XiZj0UxgtOlR
KjPvENH8FYHRsJ/6J0wuqiIJzHebjLuTHYftrUoiPuF710pjcdRIuXc7EwEH7b8L
x28VMjbnnkBP4uUB3vtowgb4ahS01ThMaAkyNQ01ualD8s7WyltTXhwnW3l6YdA0
BKih9cAcXLx6x7IooY4k+70+jaeR1T9AERTbmHXpt+U0DZYfYcVtw3gg2jql5aBU
Tu3SVIq10gtjHDwGue//Ib/SpYjBT7S8AvV5Jc4KCVck/gs1+F6IKEHIiJoUX6yH
MigR5FvyiZNUyfTe8I9v6Hpv3aW9LbKq+Y9dCThZA9WL0vDXPIDriNOND1wiCepB
piM2lDVQbB4rr5k1QZ8vlxzpzcSUDTF+kIZd+T/oaPut5KXC/Rls3PDBp8pOajkQ
fZ7IN8CqF1rSYpQBo8Mur92V6y1GJNht1KYGMPMQ7B7JrmMJXGl+0bSat+U55XHu
xzltdkG2b2AH1cSDJmfGTmC5k5FsEjSJQNlrKirxcF4733V8rUxgE+NT4efF3Xsl
N9Y2UVKC7zJM/CAfXLOXBRYz3O4rZGVfPUJgD3F6ar3W3hFKEBs6yWfoCglc9Dum
UmS23kh0XAQVEn1Zv2fzStJCED02kE2ISLdGeNSXZAc32NGtmvzIpTkTbo/fsqtF
IhHID9Rqbgl2ZSoi8GkW9RkAUCr9fqVJLE9p/NlJksvyBALHpt9cDuddxANp4fiW
cKe4P3XUzp61G/0Fprs5QQ/MOZpMiWYbckm/4YNQiLBocb5SbSmajl6c44+CmKKK
vOItAmXT4QQT1iVDftN63i+BKkZCY0fXeD6IeZF8Bg6uAs8yDxLCtr6V9dOo/KY4
v34IGpIdBD9LJ2r/kD8fiZaII99ivlu1lfyBdYiHZ+3/DudWTNkTj36XFZz6Gs7e
0qYV/+aDvRpuVkE6gbjWxpU8shYvkrj8G2veZ1sRfDVm4pROyyZqGtFTeH0tp+8h
cOhihxCZrI2T2JnzmAvBIP8lnHUqEiiNlvZhlCCnwCam6ETz+XCzN8Uuuzv7dZty
Pnp3E75CS4A2bKJC/5k8ciKSONY7Wav8Gs1bjNJNZbuHS+XVHoG8CPJkoa6BTKNu
ly5tkXjPzB+OFf27WexZtophddwwy/60g6AvWRyZ15lqD14z7TzpNlPBW3Yl4xK/
DCkR+C/1LcjiV5lgpVgrF8oc79iIcaJilsjWyid8RkELHCMizpNnhmP49KIQ777y
XoDxJ1tieqM/al2jplORSsxt7dLiEidAr8mOVhmPBpr8V2OU2rY2DLk7v9s5v9/w
Y9ILJULiEe6ri04OhcyFq7BhTFaD2pN3aeHOE5woFZ4FhAZf/EzHJ5lHcNg4VBRd
nSgo3ihL7zkjOER1ShX6KfVgW0YA8zwb5S7o2hQ9MN3NJb2DCwJ/Ww3E9ECDHNVp
JeO7InHxYJPEEJGpcnc/lB3GEkOUq/I3OjYB1a4Zn/uThI+1knyq1X5GJPJ1K7T5
D3cGSbUgxXBZC8G+LHZYRtGnrMY/HXUZRcra4ndZeb/0gnbHZB5BamChS4OQ4Bui
gg+QzougfKF7ORdcZJhhObC9vn7ZsI3kkHeKcDkX4w250Di2PHMa5JU3vWq5BFEf
Cf5fsbAe7p/OeyP1xP54WsNppOwyM+J/NqneH5uCSF/1UOQzGlawMQbaCeZGssvB
+qZ+r8z+oYu6lY+X63BCFAcxlH/K6SvkyeM8vWqhyFYgR++V9qSJmEjICVgXF76G
GQfnCzrfP6BOkCGgbyydhSz8IBa49aLOHmJBMeDtx8OsATp1QiIFnUEo3BZl6O15
C6SedJStrn0z91+iDtt1bTXRAji9Xvj9jmFHUraO8lRrBk3MiDCP00YHiu/YH8zg
4nDYrUvwX7fJQ+qPEaUhgWBLgrt3z/ykcab4XyTEhnwSATYd2gLXT+Y1UCDGW5ae
r+j0S1eSmHA6J/m9bbGuSPrptpMwqWOCcXJmKybzYOiWDRaQkvhMz+sV5eP7hHEo
rd3GO+fRfTtfa+CCTA8e+NBHZrEAwvqFjthU9GxmI1KLk5iBghGw6T4f8LhSg+BZ
U8uOC9P6sJP+Mu61BgQiw7GJm0SW1YR+vFxNPEPKOMbRdqBzODcmdIkW/B4oVDQP
DzhBG+CvYDD7EABuTx0ZCK0AXWCzGJ8cSOza2AiVNShyG3burqyVX8fTIA9lHwCV
I+ZStVPEFCFY6+C/qnDK/RNjYIwy/pAQJULnKbbRQsUEYj3ZI23bQ2Q1Hy9tb6Y8
bSLiIBqhizNJkRxyUJAF0pYYGNpIDTWcMChZlykLA3yo6JH3MP6fM3SDAvL7Q4r8
GaoRawsvsBV8ZXcuwZkEC4eWq8jVnaNGxAW0jlFhzPdMuzimN/ELlf+9NnJn+u5u
YeaUNY/O+BPj4gxZw+QCF1wW44dl67Nb4w2DqAY8LgZO3s73BG7n8gc7L5VuFQAk
sVXl/AO6oHCm/S9mqkxLOQSoVPdrwX+lAmJ5/e8vKcMOPXCnV96lcI2NNpVlOjgS
hz6V1UL5jW6TFRiajt4eXtmJZOQ0IQvm5aFixdzvdCHbtVGM5juzYJfKFEGy7Ewj
h0G4kIsdXOdX0Xw5DGrhJCY2PmrzXBbVyboLMLCrJS3pkrScQ1DcSfnD4+YZvj61
8lBixQrQX83UntBnlObMi0L84sT+Ig+HlwyV0noGESVqsYauglIXt5qWbJ5ZadrP
CtG5mK9wDES4VBTHhdnAqZg9qkppMDxjJY9B0QTw+73wio6tKfSxk1St0BcgwXS/
PlSlDaP61TAN4NLiw5rsWaAhV99+gip3Ab5GeTcaBlptZe1UJljCJThHLdQbR/4h
iSdKtfkB1ajvgt3qqCueWUjTCKu2Tcu2W+7GJ2ONnAnm/L29sRLuVw/RJ1I4NxAj
u3peMGWexATxNAQbgYasGa3X5YAeXngT/OAZTAA++v4lAnBfwwINmTobERrCZhuS
c9vUWV8LKpcvSiRR6VviRWeTw0IlAX/7oUry+1BsRhPWmX0raudFmFzmbRTk0TEi
NewH4Hwv3ut6mTjrnl4ZEXnNqDZd2csV6UWseMx5zgVs9OuCT8ObIhsjguQguMtT
rI2+4LVvg/aMmnNs+RM/lBXsVm5xOww6QzRXxUo2fvZC9a4Nqy68y0uxxPM6/Kre
RtCNNxjFXO03M69+MhN4kNXrw+ckcC85IYZsMEUe6usBFQo3uftxtuUZa3uyXDxQ
2ziZLzsHfgApPkTVhFQEGGlhmLQ9JgcDzMWHEmAWhqEUd+mlgXpqmQJhq6+0ydIW
btDZHJF/XGgHeUC5+PgwQy/Rz/t0FCIkg67mYro/D8OLQ/xVSrEeuTn8BfiDtCqc
F6ym5pQVtEVvdL6fy5Mt6gsj6cjhAG+YeAprqT3qWx0u543l+8ffDKFQGH51fZQ9
5n6szrlXlgx9la6V/kJMuG09Vn1xOSwPi3biA2PKvra/fLTs6mzrtrdSrzQgjAPl
IOcBqbq8R4vR93BPbpNjU04L6hjaqndJJS0k4+pYCD2LUm2RjXZi5NR/xVrpeJyX
wW/v/9R0Cc67A2R+5rbSvGhlUgyfSM8DnYWwsfDt4MPxv9v3ZV3Ry7hQX5Yx1igb
doLDP+8P5qpFdr5sT2E5kK+HPvV/0pXrwm0G1j46jNAJSMr1jT1YOuXLdsX6tmvK
PWEL5e5JFrl9FNzCWXVRfFPD6kRCuOYhcmF/5JnVVuomQsREBg+OrjUfBl2pwwJV
SlRyvnX4mhcGfYFOyp9qxcgVLLhZO37l9JEPHtunkLlDMiYKS1gt6CrtDgVxfc9d
XGpZIGlVQeTrEueaWeNLIi/T1m7RvzC20bKWWbbaxHpTo5oMc/77uCYW7tRcRkyF
3ZGf/ncchia9NnA/b6UTASOxblpfvTl/VLViCCYV8CfVPNp69ShuDJ1neYkd2Fhy
5NDkPtMarUUCNjY6KCh+Z2Bh9C+gxMsHzPeixSe60MYZ5gxKbulUIZv0NqA/NhhE
yC+MJ67VzS5d7au0ctK77KeAoPnhgirsX3aqt6wnEWS59cL1Ld9rryR2SqOgDFQi
Qg6YBgUuHGExNxcf6PvMTjuH9U9XMVGkAILMdvNR+ixl09bUEDh+V6kXqaVEg5CA
WdsQ5xS6VFYfPXpJbK6rFsxCnkoekX9gOPw/X50tXKwKfw8G9Xjz+OJyPp+tjLG+
QGoNe4g8C+Kww5YTvwRFq51qjI7e7VQ5KCQrTnNBXsPmZfAOHsUNCWufvRmrJQug
Eu6Gvf6RTNv9eZ2nuMwy7M8l8dhzWWUYxJGkobOBQg+TRE4IgXskv/QScTHCWGII
sprzTVng9Q7cItBcksEZc2KkwHh9neyM9DKpu7QVCmJo/+QVZa/Kqzp/Ee97UP+W
lmZLAFybzNYWbw2ekyBZBaKi1gygIxGCmYzQTXY3uW1I+AFPLcK2sKIS5mmZTrTO
3MKUTpX9naXZQxB6pQ64Ab5br5+ihXO6gBx2yl9uA8evkJmdQ1Wcbnao5jk+wEgy
aQZIfREyY3tnIewO7pretYqfaHYSJyG7fURaov3bNp76cq+nhZwU+AbbPqAoZxO+
YRp8tjI0XyYc5pJBLEjeRBLFXt9Q9ioIHJmUxLKZD03NTb/TVsgbtkIwlxT3xOA/
2tjxqnq6AIjKTocGN9otydJ0X/eCO/BJK7FunEYCaoUY7Ijcz124hUWFvDX/8eFT
C4UP45XgXGoftrnU6k/yCfariIf7UET43xmXvy6hjGPFRunwPbpto7qI2Tuhqqni
Qx8s9mk7E5oy13AbzV7SyfhJZHBPn6oR+EpbAF7xBEuyQ6IYkALXI2nGkmqGLMtC
LVhRFbV3UfIbOAN8Bb0D7oic8cl7s0bXHo10EgYkysFoHovkQdHnNg5/CsuCOj3E
UmYwcoD2f3Snliqaib/JLTr5bNCYLXhtQ9Bb1NbhSwQaiqsev4Il0Lsbc/ZB95j7
Aj6DzYV9p69FlHEfY0M2KRJwATU4Dg9lcqkS94yXIBUrFA1ATWBFZ/ZqqnRzAEEE
qCXEHE1ObK6yuQUHPCCYIJ4hDcNCNXkdg4qfzgyBVy2hqXHDCeiiR6SSFsekh4b/
E4DRHhJbPk5c+JARrqUxcwiJVQ4Oqc7pRRan0V4ZG3fyj746SSwhnYnrLo7k9QOT
skKlwI+Hz1U3n34FWTJtVuZpWSJ7C9tGXXfcBe8SG+0ZnxVSt1c/4V6EQa0YJfWW
iEkqohwQfYhpIb1KEdEPYfGqb3rfatCgxDXe+No2kcZyD3wd/DzeDPuof5or+z/M
pNsPP3bY+2kaE88lHsYW2s5mptC28N1E9tdwLlUdas48ueK5SnnfkSS3xOWR8gFx
ihUMTnlUcvBvqHlzhGTdZlE3vadcw+FLdKYJAZPJxMuzQt63TKLKJHuHHFzo078A
5f0sc0NXx9/a8RDu5adHwdB0gD7rgrZdLiOcVGfjLJVg2bjHQjdjcyeO/ynQYkwe
znUgKnHMVjohAcHfefTYXyVuelh/KBE8iA05lvsg0oT/7De3lyNJM9OYHAeEjvBk
UM1q6qmeCeVm+BAnsClhb7A3izw6d0HJ+mZr9eaSG6SZnbBe4ZLsuzv4Ha5nIl/9
AaM6PQrdr9oVKE5o4HasXIOxKlm7v65DcGiap/HSVN1QOvUdE2h2tqzwMyItzl11
GRjfjuOJ2EQ39eExbg3LeeLKvFdiq+VTRLhIXl/VQa0UG9BE5XOkUD+Y8hQN72Au
dlPuUx25mzM/j3u5O2m7w/oPJaJgwU5+gwj4MyyyPxipSTWQab6WQiMuuxgWgjgm
E2D1ZhL0CdxuJxB+SYwyeXU8i7v2J7/vUkJ2WDPUkXeidMgHPCtnjLW6fFCEF6CV
LAwh0aUXdIv4yQDDIzCZ+9KsQ+B/h2NxsUKKepcceY/ArXOXybPrFHI6d8KUqkpk
fS7kJlL8ROuc+yr+SYaclEb58q4FIlnf3BLA1SNI5qbn4XRVVytd0PJFns7DscGp
adn58WNdGldBZSmxzeQORCmL2q1vLaEnpfzv7tqS7ht3Z6PPss/tMaHoSNDmcSMf
nq8+cW2C0MTTAu5UoxkEWnQy5+QkYL7MKklkxq+7SQHA28zkRySVryMFr5WOHIo8
PWBK/pFc+d/mH6PQeQ3qO3AIu8X6GwRncVsz494aH0jW4w1aVZrmPv6PbrDDb5Wc
qvk3ZqRFFwJ68DUjeBy/y59kLecpA2Zdn0o3N1mKjgbqgbNpWShhsbCAvYHaU+Le
DYE22vM+hFJwOZdUocCpcHBoDCBQcd//cESVdInkcA9HsSuIblLXW1mnMMTt5r1C
yZ8Wtyvqpo+6uahoAIB56jJR9jYKnmkpSnBHQNyzUnYcNQoPY9LlF+1QE1ngr7w4
paoVo431G0fegCEclLitM9R+T8BGNmexR8gLGZQ6cpTfuxAlnH2feFUnUt1N2Zpw
YBH1y0h//GE2Caey/iGx4qIgvq43p5TepsTNgBO/B3z3RPNfoupCiHzU+SpWsfWJ
GQZIQmYM7uc2+UOUEaW91EvTeiplru2AJgzlCRs6iIeaCHXA8YkIuhdRalbZxvCG
rj9BtuJv5k+HNMIn7xColt1twWfGpzj84qIUy5fy9NOvRfo921KKqYadMIBObxzA
8yDYZFOtfQiBU8vX0Ij6k25lJ6PU6PQgp8FextMlWEW609GfqMAcAFj37SIU2IqU
D0bop2BATtqq2mbrUN0vpIgXLs11TMN0USFUWbAoAhOebVc7tokSKMDJtfRwQfPM
inx9WDu7V6gWNR1OK2enkyx4pJ+uuUhBJx2cAvgooWkerAKF65v8To+M0xMWbkPr
V3BUvwOOMs13JV7zkXTP07KbOmLRXQAkh1wz2THbTCC4m/oSHPNOgvR4GeG7hz3w
MXw9zFXfRNfrQAir/eDHfgiuQJ4QEFRPWSAT7OCas6SbZU4HHXy/F0qf3cUjbXIA
So1pJ9PhMYHPOJW5iPwzYqoZgEnrLka8lOPDQNtzt/8bkoIWaeDnvelZ2DTVU7NF
goZIPHWsGQntowd06Xu3ap2Jz2SKSH2fbdmpVjS+/oIdpzGb3e5yNgwJRoXs4ctZ
EJv1Q+6m6+SiXIRpiAdj3YnVbKFs0Oo5VS3jL+NAd+P5sk9rBPj8Dynd+8cvAoR7
c8DdcvTg1GVmmeEzf5ubhsg2jexkeCjBxEL1jLV0ZRLXmC33kpF9IHNiyX9C4JmS
NB5e33G7Bw65pdc12GCOlgMW1EKjz6/CSasvGEW4xiEnZJ0m4WX3dDRPKjE0V5Ja
+JZH+dP/AyQTYHbk2sFPueWAIYFmAABgaYZP8w4anvKkHYc1dImX7VBcG/A8TvdM
QUwnM2htVHCUlD2Q0N82rRVQcTwgH9DqzLnX5hrNnoCsOb1WUeUBcjdw01GKI09Q
wGTKGQ1XqFfEu16j0fqOsUsEuVnDF9TUd/Vazy4zVJ9FMtB4lLmUO+YAcsm8hQCI
7yr0pSHRGOgNEGzh76hm5lBlxmkoF8B+vlTYYE4mr+ySIVuehQO3urGIMk0wYbHO
KJLkGInENzIlhiDKrw60+uZ77TicaZvgfnakHXGWIf7VD6DMXO4qDVaXteoqrEvq
k6QqTnty/KpdxFGzf+fwmw5ewqUDYB7RAnIf0xvAQwPQIoRNXRlj3P7nCZbbP2/d
+Zr0MyS8MCrTjYencBwFks5T/L331i+Z05Bs4wtAXrCncL2Yz6mpoJb4YinqzWFb
TQyzG8r067itk2iPSBqjCYK3/CTiRDQSlQwIy9wwKm7SP3UKi+Xb7YZDcmhvSImF
xuwldx1UI1NPxrBAZC4db9V5XpNFjJDRyFBp8z/g5RWydHIyVP37i2cFWObUTdyF
N8Kh9cZUOHzS/VVHBnXxZDGFAuKC6NwaJPCB52rUNhCTdhELm7yD5sCKtfqMu86p
M0Nffuaj8LQJNThzgjFfTVn1brL9rMHCenlOserDYdEzbqF+SZfpsrHKHBimM3s6
UNwU6/RbUkgi0akn2YaeuAD7mdsBrSxefUj6UfsjQCkTn6/hhBkIyF4XKV9VBZBy
IGn6LLOiYlEe7NPOEbjunBGsrVdI/VDU/NaGCX84Pj82QHtOjobm6y9lY0Gmf3td
5plPl8UNSfkkG388YpVBSq7vqRposlc0mqIeJ4rw7S+WIoOGxW2RNtTNcxVEDJpU
5/tSuuzccBZ7jel0XEDCQEFqwOa8++u2POx6R5QIcDDCsiCAuiLQSALT4dNwFVei
jvnLcDGQO5wUy0iuOpBRTB5IMB04AG738LWOlHaaeoZ3m2GRk5dcB/awLg/d4FMe
U/+2g7X8f5gp/ry6DZmxsZZCjkOkQTrh69HRqgJIR3CwYM53z4529lv4ic4De5Lh
nRsWaLp5jDQvoIB4C4FXftBLFPKBAygxawN2AhHfHZF3Wz1mSbsO/2byCba+bNLp
vNlL4bHxNbPNM1LKuSJ4gSRdfmCE2+Q3OTUOrJEXrEyjqvUiOs4cq2pgTXtLMVUQ
z2oi4J6Ghvh9CGTO2CxP7qH2rvwvXEggtKFmkpUfjNNp5SRxMyTbsA+ZrTI3SWUV
kAJiX41wFQ2+46wAHqocVxqlsPs9kOUPaZoSW2nVgcmkGI/JIOoHLEoYZufbP8lY
l1pgmYXiu3XaH+SO0mAk5yepU8EHXJ6NJG21Uzao7wJTFWiUgx2VsB0Eq3raOLOv
ijesvsYrShEFFkRj16TfltcMCdpj5IsTOoXxzzWq/BRLlJj/zAVpUXbAk1yV5w4Z
ep4gnknqyt6UHyIJsZHPx6kPt15tV3t1286UrjcZV96uJ3Zqn6HeSjt9t3qqUVIn
b4MU97KZGmpwlFyuw3vmDXAHIbyvAvFhx44n7cmrRoWQg7dbGBxZ4eImB8/m2lKL
ML+z68KuIpky+ahWGCoLwr6o/51oC0r04isnuIiu0ai/ZVkgURv73c2eGLQCIutJ
SE0Uf0cxOxRmfn00+u5gHszsTwugZf8DDLKUHl0+SaWVx4iFnhV1YSoPKYtcnQRU
MEL1NdTxFYG464YbUZ41UQ2tvljxMkDVXPKqOf6W5zkj2g/pw9n7/R/DACcVlZ2I
J/2B/9P9Lt0zh9UyKkdrtEh4piuPaZfrQtF8VaazEMrOgmLpUSCsGmveqSHvAemn
z749nb8btUipbGTjho96iL4b6Y/ruzDjBW9w0M5xUrcp79XrKpjSUGFJRr2IyBB7
S7x2+7J50jqZXuS4p4K/IjmNXDwQQhReivM8UyB6pLHG34vog6rZFQzfDtin48hC
eW/NqjX95eHyc8Gl3vIpvXkqBAtLIuKr0dV0jeLs9VemvLNcfCD4fc8TGZLY0z0e
nul7yhjcnMsWmbYuyKEeSScDerwUmBbftBAm6moa7Hn4VZ9DNwA0xDQrchsM4+qM
8/k5ptTrHUaEFCP2g3pOAmP0RlpKhoQKzdsZXXhCsLSco3I0B2jS4pS918YZME6F
KtHBGbkKaD8KiKnsFe1ybWsL3LEegFO/gu/pivsTdex9on0FLzJGCFSEagR31n5B
7UNSX4JBbN+t0HGmI4xO/DNbb3Qet4TkOxCpfzzB7H6IOqj4oPllLoxEuE+ZU+jS
HUbXpEIwf2W/ugFOMNsS0L77grDTRp3nnKIyrzb0ETpz6dD4L1hilrulHELVPZvt
/6whoj6JFUfuLOR3u8RQRSYChd+BgJ3eFGKtpxEpETOTwtcuBnoDcaFE0V/kBqPe
828wXaakbenO7FkfreL1QCoUj6nvtQav6nojuuAMGsbfjlD/bnpAhDxtwWyLw8pq
K5L3GgZsKOpwARbEiI7yioQGAHp8fi6X2qy+zBl4jSRZwMblzI6zzRMB0jd34b7p
FNfUUQYP4fLuzHHfmXm1ckfWme3XAoAOeUhpOLIm5GHgomOVm2/dUNTDqhaNX5v1
14JbO4BdTxr1hXXiZItkWeL16ktc5J0jWzNsJueGh8dqG1mDiJfryKrgJjc3o5Ou
LmiyWRPjtSoOCoXylbEMxthpxuNvwtxpCkmUkW3Ow7cVG2FY7pA/5cQntJxfcxrM
hwM5sL42hXF9IlfJDZVUh/D2VPmxRTo6fVIB27ADWgl9o1BtWezABDBH2TPgFbTU
C1k/O00y8HvA5JlGrhJBSuSAChgk5RdsTAKzjpXRVciR5HZdLJ7+tuF+ZsgBhMat
vRFq6n2vo4FFe/AWtIM+Fd3mBtEzXmBIu6fyYBeF0DPl4Ok/Fs7gMJralO9TZrAx
1bPKZisQM+MwrUMGBJSt3cfMU1Bf0bfZ5c5hI3slLeiNx0legyBXNMDQ9cFXq12M
SceVIOa5lEzFq8zsLrWYBQ3FGDR26ePFh+3QI0fhxe9TltgDw4KM0JHiSjH8Zxcp
3Q/Ktq2qescfeXjl/IqrB3sRsmHk4AFROrm1badNTB5FibwKQSucdUbY360AHsm5
fXAiZ6GlRFdmyIqAOAHZ87n2GhJwuwdegFmL2GpfQhqZxKUJvIvphYr0UOVcNjXS
qzd0R06IbnJB5mFJOIgKVJH0YRTBd7Tiff4DoQbEP6BNDT3iJs7DMpsRXi5w7xfB
Q1KJ6J3+W9X9qf9MTAMvTFrz1xpEk1FJGOEv5xld3cE+bfu+WyRtb//H7OYbclPF
Bla+mi2KRdUzspI15oWkBM9JCoXZyZJy0U9ADlDHfQ3kUOH02/zsMajIsE5YddNX
KINctqiVpTGoqwPEwVgiQ7//O74E2SkPQ9RxfsJ18PxxIYyJyVJ4S9ZYHpS5kwbW
uf+D9gKkLZgocR46TMRgNtwmbFdULBagBvl7XAXpGwTRggh2K03eidxfncZJP91/
MO9e5mm8fD0Ytgudy6/Tiw5sdtuii1Jo+biH5eqpbGzBsP6oNa66fzGuVrPIObqE
gYN+O6KIum9Tpy3JcdhMD/YO6+P8lKv5pLCoZxqp67yT1BJDuNVuhaB3Nl9PTgjA
JE3WbMoZ3ATZZanWq1230TtmeZzerGN46QxctX30W2lxln1XoDdbhqtPuEAFM7Ht
S/XhlV9LsaSZi/0oqzsMfHaJ9JnrkCZ5jMC4EimU4yIp3PTZd5neupA1v4xb8hsT
/X9nnsSeskohrlsuBGet3GNGc8c1nZyvEEjlrSLoyNliywRfLpcgs3GXVORP18rF
UqRz6JHH+1N+WrPSNhxoPZoAqqfc3wK44xxJ2DMw6OYCjwSJbiJ25GJWWbpbxDI5
qSX689N1+iTVAODF9TIaCw3ys88R7niaTFRoKtcS39y9WdllysAI6A0iY6iOJWnl
5s8Fj3Tc6MCn6+m0X6btYFfj6wCAY7qyYKQhsqPCaGKRfcoMDv4SaDQlhzKcSv3d
vXh5LCYUeAqV5XCtuYBYMZ3tsGx8+TvYe/OQUMVpWMY/PmYLBbTVV3H1ML/yTS4I
XaiDf9kTlIgPVnu8WXDyDlpNRZuwO36W2FL6yNAPRJkEIHC2bkZcszcGVLUGJy+r
UHDD1akS8HorZ6wb1Renl4zZPbIuK+LoIuMjRCH3QOU4OTy1/w1WvMqh3eC8GAFu
jighSDJ3jRlou50LH8DrKI2ZhP4N/mgakb3d4C7008aT1WLH1fKzAgRpJkH3Ms2B
LZS+UZAKUo3Ycq+URMtgdci9RiGIqyg/IFVmobzBg4C7lPS2MgQBbayW1RUGmefJ
rn9jsDHkV5yqwSzkE3IRa11KkxLaw239P4QuuQEpntIdcqI+53jXmpYdstlJRrQg
Hmw8yvY0u2KlVY+IkFEob3Um/i0s7NZPVYy9V7VNDafM2iWOYhNrdFq9u54RvsMP
XsJY46lqq8p7lOySohqi07m5exEDH/Wm4Zvwq2xfQEl9pGVi6mf10JMXHKiTSSNW
P8djyhckNCTMp+kFgSZq8MiivuiTxX0/5m8bNSlT6qcR8rs65Vadfp3WMEyYnETG
w/xJHa/fWQcb491SjFIPsJoBPdrYyKQuFP2LdXoCoqeOUvyEjbE9NiY+riJfE4kC
lbFwoYq83Ut6sD9Hc+ZDNdf1fUaU9iebOt2/Ac51nDNH9a9LI4lAfiGRWy9LXNkh
Qv4Fbu+RcVWp4sJ4VzP2gxvNyLw3sNLabKcR49lxsLU62lB6G2niQlRb6NgZ9jiw
/FXv9gbW22JTtp9intpRJcwzkT4eEGv2txesd7/+f4OIe7tgQrE+k+9oVE40K7O2
wAt7vLaGlG98N0P/n6xcVPegaYk5ikqgxJwfYJZLzua8CbDCA4Bm/9fQVJditR5l
FDf/SiNjJduh7UFaSrH5csGb2h4QgRDz+QAOXLw44SR+suiTeADxteTBzT/0I3t0
M1LZDyzrKcTsf4oDj3leNA/EQL9feQql06AxA7duMaEtv9HDVO7a4ebiBlo+a8mH
OsO7Aw559KbIhMox8uSxgt8b71FAApLhUyOgzWR1dsoNIuNhEYorDub+4Z5uuAaW
7veq2UMRZIBwN5Kn6FFLZclQVPEDCM4Z8VQzNb0BMDOt0u23W/DcXYEWbxaF5D6R
vjMh8oT9CVnkAw7c61GvVFaQxAX6JCkdedgdwdyPDUyYtHncs7dEL7pqw3deSv7V
n6icvFXzCr38fGop1I17Kyeaj/pVlx9T1klGxDXxKysPnZnI6IXmeG+b8Bmctr5X
g7Y51OsaEHbUTXzgeV1O+KZdRjtGzv4d1nVus/mbRG+zcN0o7ktq/hocj5RPoVI3
iHX1N0p9U5go7r5gzzetKiovNo+OPQ8Z+BIiJ3tFIITAQHg4tno7XU4DaMG/28GY
I5CsnwiMqnrUzc4htJh462IveOPHJJC0SvhjZwEz8nM3LR2IDzk/1caR4KAP56SL
XcHvhLBVQY8AG7QsX1n/uXhujk887+bmZwI+1cofhzhGKKEvJQ4Cy7XvrD17/jZT
d8AQExvTV6azSNfL+DqKXb8P3B9KyRa70w+JpnP2AONvrjzH/qgG7OhqwUKU2JKg
puhy20qRyz9sq62Zb1u3VJd6034I8X7+rqVb84DEXtNXv/3RW13fgoiGb8aIgHtC
bo0Nwu0Gliuiit8WnNTtYtL68J1p7N8TUG8qhyKP6x8GFTcPWeZ1qRcqHNoHfQv9
53dKMwjmabfa4YyQkI9VwmVbg8hInQSrKSeZ7wDAmTzaxjj8DVE3yo95oTlcvlug
kU5gRdorNCyGZ+sBRhI0zjbRtSbY0N+Vkfe70nmb20Y2IG/Cff3aaycRgt1/Im/a
ruVX07k3abZSgNuWhYCBo4eHGsyedRLJhsYe2z6PyhrYhe3PZ7UciaPgX9Msir83
JoKrnNv/IIScWg7MLAJqJkDZ/ItZ3Pn+yFnGjR0f4VySg1uoKMtoCcULoXrpQZxN
NsYmK1zyDPn0v4ztRPCh3VTqkT7NpVpr8MHZINHpKqEsq9eJPNp4+kreQ8WhTpc+
P877EQc3WmK2F8EUacbp+8zFdEW8o1bZKRsT2H6M0MKwfP3DhSB9Kr23mJFMdrXC
JuUx/ossGfbN/C6gvyEwdxtFEOXly6/ihtv/bSlE181AYMKoe/yrCKgwnWis5Lg3
eHLvfJvrLse7yyV9LTx5TE+7tVNYo8gAqXf7VDs7iu1RPuddPjYFQOzb7cuUzNHI
txMax/nk2KepE61wrI8YLxHEMi6cz7tp8314k9x1DbtCceI+k/iHfYv55TsW/MOg
geMh+gFH0/HjjqFVxILpoVBvCieXXPHmPe8qV4vj9iDVB4a/WPpjIwpRB0SoEfNv
N4jgEjr91pxhzrndkONwgi22u0NVRioKTyfOjX1oXl7TekndSyoavMIMedO7Sxiw
ZtDaJFeGl4g9wg55YYgDwIbugyqs94A9V4Eb05GyAG/4Ho5b9KWl7x2G+ErVtswK
ooDfRplaVX+c+nOwQPV1CUWNIOP43z1+kee0QzuQIVN1bz3fD7vAD3FxIwxBJz7Z
Cvas1Pq49lMqQHWphAYL4jIsJ9GPw5BdpfNuLRio0INqWy90QoiefLCJDkbxHDtd
AZGC0T6wFrob1TVXUrJ3Z5Rg7vE+kqSj5/TpMmH0DNssqIifwzXaDvK0irpfVSCu
nENw/n/RQXgweyr4vm8LLulh3imm1IDVSHRl+GSIvQo+AmPKA7sPvwPHQ2XcbFSf
83+4HaNLRjfRnd+UL3WOerNpA1Ct161XmKYwMieRiSkskPBcvpp9D4TBTqgCp2dc
uuuJKq2rIZF+U8tJ7COt8270ya0CrZrJcUtBxkORTjlnNVca4xUaUfwiZEV7/1tv
x66cpngVk0aMKNKLMog80sQeGlgDd6tmlFMMjjaEEfoksga1bnZ6oMsbCbl3dV/N
vlkB5LcYG4Hb/W2ucHTLl0jBulzqY04bguQgzKCkiBAsTJTLRaatDb/62oYsASKz
hUD459pRtdcKcDu7nXeSwy7T7Bh3TsOq3URIbpG9AD3Pf7Duo67+/0mm0126fALf
mStfmz68aevp3qqJlmOyIGPAyHG4cVEDesYFtG63PZmqko8loB52iwbZElco2JoH
9mzzqOJuGsQARGmsVMHic20nCTdFv8DdK84N5kMocVFg4NMyJFfbd5ACbejcrI+d
+c/KZLthb3F3k1vfqpkUfIdE+A5PAYn9NBpNLjxdUFsmXmHWwWKsOHf99h1oSU1e
kkSaALnDpobi8BSuHbf1cG/+yycavtL3oKqKd3rCs7mDXUnx/waXz+DlmVOMVu7w
LJZtwGp7R0UoZX84bEEiKEsgvbNuo6poKOVEArazr7lSgGERkOyQAKOplZtygH1C
510st0qUAQFwP7/Io/sd0QOvXMBoKPm1liD2yEdtdqfrtZxPnuxJLSAaRFT5aOH0
fZkxAJ9IoPDiuv/qvs9SNWKNjKQt2XHmcqSRlRP6dBr97E0cD22+4EDySKVBSfEw
DyyBOND8G3LIkCwxseOK3zn4SEl/gsUVUtveGFEuWuMwOeeQaXellgmo6yUgBRFF
Wb+IkmgvLVYNDm8x0hU71HlQx9jo/kLqjNDHKO2yWE8uAhncJtAhGn91ETA6jin1
VTbLwCZQvfmf+AYVuCqMW9rn+IeTIxIB2Y8Z8e3i5rkNnTmpVREaPovfEVK8Isf7
XkLIgPzBjtC+1p4Qy94K2Y++UIf4HAXEdbwVQG6AyS0PuDNBLHMTkLntoULpCIMb
CVab/hbARjED3Ku7t5JX136YjdEnJKkA6Kv5aEnfWM4fmDNRF5eORWcp3Fd2+t1w
OepT6i8MrO7i/dm0U6NeD85kI+LgHIGSvVZsDE8SrsA3gat0xuzoty4RCJPECeQb
SJqV+s5kjXdmu0CCgEVe0uKlz7/CYCswOmz+buxAkhR0r3ShMUeRinsodw8LeCo8
+6wT0cWOCTgdsyGbl2kJi9y0Rx71iPMFns+CO961J+eW1eiPBpQs3S37Vqsa/sj4
3tLxftyvyIORjErLsAUMCs/xc1DxDFPSZiODWXPhHdLKldxxHmdw9KrWPFPKtwob
E5s7cao+Q9ERijoLncrzhq0ME5tH5zyx79qDhkRSCr+Otn5GMmGIJPL98HWhWp+V
1j/DtGQCmkDUrp3VongfdnI7PbGQsUKQK3ncBcsjD/BWjtZ2pzg+TBaQUjmHNwfu
BinIt6vMKS2VpzjeCbJXOta96JlGiIZYedQWEcrGyIp/oeord2qSqzxoGTveTxn7
zLa4OaImDWU95GAz4APJHnEDNYIHNPuBKnr7qvbPlM2EQ/mXNFI5dfMzm6GxEaGc
4JgmtKJA95RBP3ezT9+J6mbKpcOoXSh44FtQBt4Jxjs1+wvDP70nOoeVox1Y0mdD
YmC//ghGp025D92QAlsIt5Kjjk0Pu+jEz1cPXorC2D9ZvLVTQT5zxThMuL2Gyhri
CnDCk8KG+RhlQQwczxLca4mtKjDhGWFTP+PRFupwjsE+1sc6rQH9n+w5NfGchdUU
Bti1fqWJvxCDMQqQJtU1P+01SszKOSg9owe2EneC7D/TI/theqi58HFJK/HlDW93
CVe3hXY3CrB8/hJA6xrc2XlqAvLOZjEliUo29xCAV/+OSkExmQzlRcUkVMnI2xfj
GEhluZb0876rx96yUJlgPix+YgagM2c5r17zFRLqsBX82J4+prekwEW/GvocOkK2
bayzBOv15GMw3QK6ZxzRTJ55M2nclbtSonOhK8AGgfRd6GV2xaFSHT1ycFQeZTtN
kxZbYQxrR4n+aiSSBTsNcXJ5Fv7IOl6sxvXsZecpx0wQwxJ5KhIbzNDpXDnGn4Ql
easDOFD8RchPSEnHfZJHb20pvtX6amAa00h+BqzUwtNogpqVkgx+mQYto0yhQQKM
BbwMbfGpvNmIEZtCLBy4YXawemwyNVcqtoow0eTK8fcD8TKgVoyZ+PwJU+BU7DPD
QBIwCuPBwpRmzO+He2unSGZl4rc750YotyYeNTPgUCWGjjdF7ZWoNSyYJ4lBx2J8
7VlvOEJjuF5EpBVfWjmWLiH0QlKMcx2vR4jO20qEJwbL6w9gLVpOl7KZWzYJI1fw
C/+r/PYKVDZaM8c1OAU0OJd5t7mnTI2N+r4bKr4QMgMJ2tGrinzytl6HfXQeQPff
yD3PiwP8sl6ZYKbd3o564EAciJgrLjxC6g994a5x4FCeaOb/ExCwFXsJpjtO/I6i
0HsjupMXloPWT08DblBq8eLcd89cD6sUbRCuUeh/1vQEc1U54AmzDjGtLLoxMutI
maFgAsgLHb1tokMYrAbQoj/cX8E7ohThXqF2gI8uLXypiJe/ern3CmtcnYMj09RC
td3XSC5CsT8p0hOo+abJB8yFp51fW/RlUGMM+sff/DjaiSdGgy342VZlmMrm/DPv
Bjxnpmt4YN41dgNs9UM+dTbpmBAkwY0/aqkq+5Z8DU1VlyuhNy5g52XcFrAmZ9Fb
hsq0E/stuyrxIr4W94hZ9wBQPprLzdWOQce+tTJdmDbbxgOp9gJNPR6+FhhvHVyS
0bzn8nXhxsvEd6Dr+YgzoASdUw1dxDRKcWEtZEftMYBvbX5r1RfNIuM7bPv7i92V
AfbBWUB8QmZHAZi9Nyu5UcYJMlAlaKmzk80d0CXN+lPsfqtu5zP4sQ6u8ZofGwyl
+502IIrNxDzsT8Zzdf6IfV2numyro1kX4x3j/EeTscVc8Z3BxyqVJ65Ix6E+oDSz
NnH0CCtIBaaDevcmyXk2iK4PdhaitPCpXe+G8lJ4lMPthpd2X5BsRek6fV0wzEvW
jDhFg/VHFxN6xAAS5aYUHE9TAXDHpLdp52SFVLil8Er5Tl4ueHrDkexubIE35AGH
FJaC+YBM3Biv8Mncrrvq4G3DafmoSMn6rLUzwVgzHIc6nRS0EBnz3AgZdge20AiU
Klb7LW3slCOVDnoZ38T/IAq627qiAgGqvJMSryeqX4tAnOXf6bKjgSq4epeKMsqd
M+WDH6fgSrd18erSNGOmumKxhwStvdB+8AQ8mdNpnh/H/L+jvWmHDRZjaz48btZh
+9n36kvbYAUdFpdeZp1gbH0yPZq6mnGK4jg6kfSJ5+kbdc5A6Y9HDtkRi3Qx62iS
e/SWNov3XQC/5iOaDlXfCi67WyAtJ5rWPM+45FSIIdcj7CTRzIHLBbvYdGT1+3se
xfFUgMLtyT1eNkg61f8HVb4u51j8K4Csm/1neYAJU7z/HXb+r9m4nTwHjnOaqhQt
x/xJyeoyG2aleamQmG6jnGHeTV72e39OOoE8dPtSnvM83RGK/WH0jzM5jZOEiGGN
4b9MfsVw5zQQiFXLAKZjzurvRMwlFFy2RVcx/y6NbxwFR1RRkhI8NBGb+souGC/N
Lhq6ljKW/nmINFbpxpPQmVcaCNmSow7X0we6xg/cA3QFoJ4Tyh8dPYjFCJAxDQsR
hOpVaDr8OeFhQwyAVgqGy9q/iG05Z9KZHi2Ia1g5MExHJleNW7H6R21T9ZYZMtW/
rh6/zh1FC25dvKO24xyZnCe7eRHRQQ4Mgy/UanbVnIZaZyPFL0s4EZk+Ta1FZzlI
OcJW5wYjvMtb0ICGbCdp/FPUsvnLMND7pComNGpegPee5V9kIxT8Hvr2E3yQf6+T
bWsUChvvpxgq9ip0wDMiHqW/ykzxIrgZpY7Pwcwo5leJn0JMgB/FQm9Fyf3/Tu8O
WOPdVtNbXcgMS4//3SjqJ1lf65nQSnEZpwtjaCEiz6/kKqvKN+wt+0vy3MIhXkQw
8Gtt+lmzfHZFbaX0POEWEsWXhAjshDTMl08HFjC2VqjiMt1DEqA/yjjy/GULPhKh
KL/YPjo5OXlKm7lK163BJ5C8mqDxwB/Hnr39JMYvXQ+0hmRGUBN11YKFKuMjvV4i
KwhLrb/ufnzdQ9se8+V020QNxucHkfP+htkGwbhvqBseo0rLRpQjKG5Rx+69PNdj
9t795e2xeFcBUYgtRt5JjjW01LBZQm6DyjBz+WugNHx/QnJdoTBEVPGyDPA9lUAc
8lA2ea0BDKUUsPUDYiyeI7ZFwrKOqjR7bKDO7sWw1jIj8TZoWrLarjgK8xewTB/U
b5GkMqiv58X075YHCOjhZNbsTJpqkWEJm6Ia0xXufq5XXX2OjB/Fx19yGnuGF8hX
TsqBWFq62Cd8esZmPVN93RQJizwzUguQ9ELcoraO/Qw2YOBZ0Mxr82INPLiuAp21
3Gb8sWKxCXaClF/E2HzX6i29t0fDss1zKpvxZ4mtUennYqxVxcw8mclmohZytRuY
3nKrFdyiNzo8SytxSqxcdnY6enG8wCS3cwy7kjSvMMC2KZF3SM+NMCJMPknAeQY9
H9HjGHutRnYomiYPCrfRl6uf0YEVOAgVoS2cx9ykbj0ipooaSqsRn0YQjrY3ukgK
3YVTPvHxuGQWWaD/pPAjFEPp7QSMNLje9DFAXNBITXRv0BeDEkoivOcAer/bM7p5
7DrqO2m0qeCmf5axNAZcw3TeEbYqFaRBMSdwSaq/b9w7uFxrufvXB298D1HvLHqD
5kVM8FrjRquAozrOxPbpJPuiLWwH/AL2lzRwxe93nZpziEvVlZ0HOk/o7FfXwCxs
SAmoA+CDjbRxqOJsRF+nDJU+2/uDVS8kYGFsOXcOiFZUSRovM7y32kv/Fm+Ke7RR
GpomuTfYSp3VRqxU0Qit16W6iB2SntCPQZXWJm1C0C+MGrBW72Xae8cxVC/HtDv4
txdPQ3dL81CU9BXMZi8Rn6d1ZxxAiz0191804tx+beXQvYeeebD+0gU3AZSVKwAU
cKi7Q9R3GreN8oWfGafFgGhtqO7XUUNGnxYUgo5rsrwV6Qn/Q9ST84dH/U1YCJRx
p6S9DjCIMTzaO2fvTxAezY2liva4FTpEpBPNFkrEMcR7qHdsKAbp0mr+WfB8A+vv
5/QrKb1QIUzFS/TWDd4YX1eENkPjRZZJXAdol4mhr4FZS0UIuQP0DsXvYpLOM0Iu
fiyP91G96IutKRAMrSb19mFaIscnHJqB+buBOUS9vPwpTS4mrxnlN1bLI2TqPE3O
yPnbWOafNL3O4PSChGTqVA3Y9MXDxJWppmWSBEIvvNb+7W6zbgmusPbeXWca+5mo
FlQIbdnkBSO0jhfTnUZMEkoEFw3HEd9SN8OglksWfBh+SPPaXMmRBL9bvv16Fl0J
fmfmhM1By8M3+i5aw0ubvJHUkBrM2S4N+Bi28kRZNbDyehFDaNOg40rEaoKkmz8D
jWUB3a9AotYvDrpp0muhQ02Hh9O0PMu63a2CODicprsA7SSXdWUbhP26R/t9h2BN
3dYUNqpcXrvRUieSb/0X8MM0NhY7JIHmlDs9D6ClD7UjRdCi8ppFZXOAydiqWTfg
bMfyhEkIMbKKIBsOnF2ftFpDo7L00LlAoOhS/yVmQmB29+ymzUzn7e3bKd34Kipl
BzaOQwnvOI3+J+wWPYDlGGZ9VwXJMfKmoo1aphi6AUP9YSOO1gDaDTRFPkwbIawr
2tHXCVu738IuHk1+6W5VdBYvW04QT2p5YSLKLp0702aVKHZanjxY1ST6GCq0QSGU
Awz/ZNoJrkmV9UorHKM5XnMMhl5BPe/CPdKk6av8nLIvzxSRM4ZK/idFitXgflKM
3YVYB5VOGQcM5URs225FISlc2Az/94ogqYX0iVu2UG9docgOulEwNSuRYglLEfe3
HPMaru9rYVHmjjLtGcYS4IuPjMgXWDbX6q4eb+STswFFLuEcrRTSid6bfO7+76qt
ng+OIIccLv81hYHc7zaYTcWvdBEivFkfGk/xGtYrUOC///fLA94AiN4aajul8W3/
cvjFG6YqRtWnKCqOk0JdE/5dXj00R3RUlL1I2uYeDhNsVcC2+7cEqBYWiTuKZKkl
bxoYIQTKz6lfPrzFknbykV6wRGscmRPXOE8BR6zahDNZwd6PPNcQYh6Gtswp02u3
SFZskr+CTGZm8K4ztWf8A9qXsGwvCQGsXyL0nMCxinzflQw8C/V0HCjld2KkxJjh
M8bqH16v1wR0mD1YkfmgULOS5CPP4YEico3KnRi7ocI/Ed1qVtv/j4/EBhq9aVe9
VxHJ1d0iHNByWTvIzN7FoT+LfDGrc2UTFEJn5Rmi/KEa5GNpsAb+eBOmQo2nJS6+
Yhcig59diKFsFLgW1hfxMJXJVhbNPbheTA8S9seryaIyy1drNj2OXu03RgmrLT2x
86/bZ15QGA0epeRJBE1wgdTN64XUByOF6d9lU6PXl21COr2urnzxpGoVjWEuyaIG
UiPSXmZCgEqo6QLg47faYteml6HMhtjayCHIyfKYZuISffhIvTpud83Ewxt4T9h9
zBfaKXphqBnyWZf+ZOLRkXsVJTU33FzR0wHiP6O3ZcAqHFMNJohWToYesqnGJc6K
gRF1/GZc5yY8WA0cfYx5oXt6+HQx8UijuewcIpcL3fhlI/nx4MCMoj5cBaA1fP6R
osFxJ+6rWdYWCfBbFU/jnbgQu0j7OW2e/Hukr3hrnqkhyi4GJ8HWz8HV0uAMpvk7
ttBNuUyGi0Oxg/2UumD3SMC76PMt9gJwqpmtGXjT+EGg2myVrcTW8mJ3RTCBCHPK
KOFaap+JKD3kDLG5Zp1knt27tEqL8D45EFIp/uGxmTMvNogBaKchT7BdrmqaAPSl
9MEyizjCkFJTh8h9aMhRtl/7dqZNbzauDd1y32scN+pfRI4TX1FnC5NOQup3TJ5z
QoZe0RO8QQOAQT5JWSLZg5qk1MEtY/uN1I0vXFcuJvoD1XCtXeFJvaKG12vPa6gt
EM7TIX6pKz/x+dMVDusQQlfDScvcCV7JVF911rs1ElO0C+WvzalC+4S6v/aoQ31l
UvYGFe6ANb/xb/MfowZQnj5XFKjtxz7sod2W2jfM1WjgL5rtBZTRmccYZr4WnD1s
ZLvh6ULJpieXsyBUYXolUiQewXSP0csJEJksM3qRfd19QyTvokZJJp9X2AU7Cl/Z
Q/Ph1MHS7Vr5VOt2vVUU1GlMXqpt/kpIZQfvDBM+BfZ90w3jdmDk5Y2SKOReVM9v
3DBbLrYPUZgwKvkGd8LS8Oyi6DTx8iHhy2y/lmx6najuS8q+aLmd2O9dSH7S3LgG
Z1aKzZo7cpcLSqes/Dryp36ZYt3SzyCTUoG+apG8qKu3lClP4OffVBNRrV2gTfZO
Y8al9l3RLLk5Ci11I0WAZQ/q7XrsYVCUza+8m4fS46Df3K74DM+NDO/V051leHrD
HPxmZYo7uMipcIcY2c61WW+gM+4ndhDrTPhr1PBAhklhduiETMEVhleCTsr3vMvF
I3VXZYFW6Kr/5wMf42z4vq7NppO2ESMatb/hXYtfIOjSGWluX14NEckvxUQBrvqp
UE8bSOsV9cMwIPEkXUyAekTsmpP9/PZpmSFjRmZT2eozf73sMXsY8pm1PHv4yD+q
y4SiKCdLcz6rh834VyREr2W5uN4rZ68PeLLxsQUQb3xKxZXixM/imnMjvzcWx7tf
30tasPVDzTAv3bfVOmmzXkpVztfJXURlLtlbDZ8WV4oWZwBD+G6dIuySrH7/S+gX
1KRus20aOHB6A1oas4nDXHq+0E3Bj5oY4qP0CzTpXPDpKxkzUgzZzlIW3pQbzP28
g2RnbSQKdaxjklsGVgVDWO/3qHysVXn95rOltDr89sKmUyiSfKb6BHc4jcE55+Vv
L8OkBx3v7GKgkV+P9UVrFkPxLyHTOr63ZxNo3ZgE5E5dtqTVhWpT7CbyVv078Tsn
WFNe/JEsUQiGnase6J5EJesdmazHtei/RmB/FFJ67sdVQgBVuR66VnbLeUIo5yKM
eCDGwD4ThKRC1q+VAumiyBaIo9JzbQcEHGpSH9AeJ3l3v5bl4iK/RGimxQq/RMRn
nwyBaKj29jhN5l9cu/Fu841gOZQW1gE4kENBH6dl184ITWtfp96zxDGiHTaARBlI
AtrHBCtq7Gmcn+qnq4/u73wvoQqAVC1OSRAqvDAe/AiTbZbDFnLG83XwBUO9NY+d
LYmRNaIn/ONF78ICTAO6vOmHfN6337hv70TJAB3nJmlzxI2kPgcZpXIFvozsnALz
hfXeMbbKZH2qa943Yd/XNb8ez0u9sEOmUVPIX7MRl8hwRcLm5Ya7+Iob6vmPmN17
1qClCviO4F5HuJRASvFqClXaRn5Nl6kCxusOmEtXvTCYF2QyZPj9yUjVJ3R1djxV
JFGvVcDCLTRSZdzjYuQt94xIZzzxKhNvMVRPzUuKdRuHBeK6tG+9B2zlf11BhKeT
GYN+IXR70169Owo50Z5mqCx/j04/ojzIUvINe1ZLWYmSUT28b0jMXxNfCBtAq2vP
4vWbN+st0WL1LlixkTkP6xjrlO8nxg40t88iBwvSHgq+2aIh0QMedRKCG/ol7Ux5
nL9yZPc34VsBSQ8sveYOD3+njQfmMe6Bqzfyy+DsiKo8n0KAa6ALn4dDj0Oj/lKG
n0yJCBMElTT3miR6SQBVvmu6hY4u97OUwedAAGiyVMycAeVrgaztE+FaeI2Y2bzG
7vWVsP7kgkP5Tt8T365E5QTyFEt262bDSwFA9pUyxZ74t102ABtzdcwxUDJzQcmR
al8QtIu67AWzQ+HLT99/vOpYvvwJochcEPmSV0BtVJVMAlHUQj16AT32TMzHOkLS
Isd2ebgC6u8LieYZlHFkGSSFW/Atle19NkPG+hBd4jtIb6GZlMkexBjjcMqVJgLI
xaNy4C8NuZFUCWfehu/Edw5nL8vTwn52QX6LMloslviZDsXVbuQ5qWPCEDOv253Y
eXTTp/BLEeOsPNW2Kb/zCCIbOAoDF5phKF046FTnKwzcznzGhMjAE4NNQalyuzGK
bfy/bkVUeVyzdZZwcdJ7MhXhYeRCKqHzS+Q2ZHwud67hMwuScq4Pb1SrvPRuVULX
Xl9O8gedjWMdvdK327NrsZcnLBzZOxi19FbTM56so8IUACORAq/hdV+zCVDhTgCE
ovT4NGuT/6ODO3sABiQpdinPae+7uP4NDuOBNmcbs2TMBvMTQB+s/lJKJKdg1ZQV
pBvOegIWUq0Z+OMK5UxnuqFpbifVljYwkXtvA57GBSm2MEXQszliqsQespAHX17M
VGIqQlH56L0vPCGsJycnKEAJB1BW72P2ZNhnceRvbGV3CaZz8No5fGvXzpe6dfJZ
NRC5E8QvFyGxAgOLVHXhBqRbk4ZOrNIbFQTfcYFwifDnt892F5dALVBT6GPdtHt4
J/98qg7a4i8nl8FcWn51BiKwoIbw5UbgatdjjDge9R4bbJboilGA+35jc2pAfqPN
lKTtO+lZhwdg1tMmFATanvNyR2vRyzGneVqGFFiRCKuQL5sN/6iRjgubiJEvNRRC
VNoepLSg2q3RnO8vuY38VEl9qWkTOlultzBbbf+Z4qADY+76vZUNJnshJHz8ABza
5JJQ4XleN7fcFYyFd3tZPchvSgwPZSkaGER0dITrXWO8Tdjv212g5NORuAmhrYZ7
Pug0VQTpmaFr5BvJXm4jEIN5R9LlBL+Ien6uL/bVqskNwsLFdvekVI8RspEY2ku5
QgEQr/xOWv7vlUSEGhu1hoC06l+v4/4wpxZetdy+lGD2S27OvqhamGrb3wqRIQpb
rukzDDZDhSYJz0AkaQ/RARxC+vPca8brabORgdicuUB6ohyKekH8HIEmGa9r68AC
kmUZoPeDeMEeedH5HNhoSsmMSnsAtvG3PuHkUqmm2z6/nlG4Pb6Pp1foCxv4X52M
jFswjpukyTPzYmLmPdDyACPb6FlVGUofTcA2HV0a41BvfxhsGfnq+EpI8cCdBa6O
6r4qzF/KuF6cMQ3npWc9hHtFSWgRWTR41cHTc4yxw8xaQuHqUY+utRqnYx15oGON
uZa8b1uyLoHkEj83GQbC9ZpsXSVOFcG19IsJj8TNyC+84cQ2/bb9bGJx+MQK4+An
YDK16FJzeN4McKx3PNOz2XqFk6/h9BnMv6ltvcwhuoOZZKoVCm5X1MC0HIujdpPn
6DBIGQo2FHpWi4HXkyaBb8xuc8XhUKQt3Kmc7ev/GEBno9c4ypLI1oryqmLYHcUK
sGzxuAS411ysFS9y1JU1teCm80Ek79sbT0hatu7G0FeAWUoFnR3Rav6BuqpphAIf
Kq+Iq+9w0aJFk8ANDHwLQtmnob/tqUk3o8SYnbi88VxluD32M6RNKGM9+EDvt2Wk
yKyJNHNLesgjqWFWfJzCtU7qFwtbY/XhS19xs2Qhs45XbE6ZdEhizGczJYGoQyDA
qFnxb5SkUMoluQff7Hwk0Cu6Ic51BZ/cREtSh+vMA861SgomwVUu+u6NM98h77Yc
FX3RMNp41qVRv0U2E7zsdgxW5US2EzZWy61M2NiSp0gvrBExcgyOqQb6sP6GOJDe
HswWScggsg0tZgYVPcMTM9AIjeIlB1OFYx6i6K7563ZX1IDrfITGus34cLscUzEU
iNB3WhKY0iMSKVXw98eKXEsAhX8/tRPyHwEQu3AKoaWD24F2CXVfTzODQhBKMrrb
MdT2gMrqj7u+KZhHnNtm6xL1eva+coBl8nLZa0g4NjYCKOyQYwCY2hJXTl6IAyfg
ZdFsVK/T9bKZGtmazAUQLFQy+8m4JDnShJetXahkobmAb5sNP3bqCAe+jofyHzTK
EuraSdJvP2yZ1edn3sXGIgL5e4whZAHwc9Jrq977esIFPf/ScdEqixMMsFUv6ACM
tl2xwZxhkC5jnGskvGy+7+dk0I7TWafG30tjib+k9p284XS1+35/H7lxb8htEoLw
H2n/QwqH3TV5K14GlkwKteSAoMP3ubDc3x6gETLRGkSgNyfc9GxUB7Ni2QqTTpPs
59bt8xtY9vJXqggFd2EsBJD1XidHz6DFV8RZ90W5h9X2dTo5IuVC8vhwZJOIm/1O
UGCahn8PWCXisDej82hoKznXtzM0A2yPcBLrJKfyz+U3dcTgh6+9Ep1wDlybgYab
THgrB7oxEwkLFxq0p/9tmxS/QPn3jml/m9bY8B8rsQtlBpqE3ZFQUHSOvGKmBp+m
3KSSZgJzBl2hDCK8ft8InaXBXJOn9k78HvLftDbenL//0Er0LoSThUrbJ2xFlVZw
HpsNhuopPQK0DRbHsxROM7wPdHg+3hqzk2Mxa1glUif/zouyTlogv1Iixbvvwts4
CHffPWeM8ILkYPId9wthpBBVu4qoVyh2dGyckcPxNPSjJewcvlHzJJdCyN+IBhJA
rmfs9vBQWa+DU2/tzW/qmK7pK8kTXAGTL8imLNcU3e1HM5A7QJb7eu15MemuCRwW
YoSEA3JEiucPlvwCPLDVF79I36EEZH58CPc7HkU6nlztIOZvZm4dbzaWeWytNByw
HpagFdtVvzIj6m4Y38l+X5MEtGMTP7Yujp1tdjDR72APiNFdiVSb0TBz8sZBv28h
C9RGKXkyPSuzWISUGEd4ffCH/lT/rsjILjslAnYuaiFjMCKJhaRoEX7aO9ZfXDnD
TENy25/P5MO/J/+SelHSHYj6611c0RIrFWm8eFRtbYb8QuUEJndN0S22fDgiRzeA
8HPpzUNZ+2hL8BSkZKpOm0LP0mnZQSwMJrd/b3b3w1XokH1g5C82yDePmqGFJ/Qi
NNRvfYGxGW3nu6uU61ydYH2OW3MYsm21wqAn68xgNJev7jQUzCBSzdCQrOn6krWY
MUjvC3Js5caX8YhylRmbQh4ohbrML1cRf6h3mxUpWrg5b0qX44sWwbh2ygFF9IUn
hhOCCJnqMgqb+el05T5OWb3yRcMmDazgwl1tBFFjfptStv3wTqQDuEkSQRrNQMmk
oi0qaK9He7dacmmH2S88EHY0rBLPh03rbG5E0vbjr7KYTxhVMqMRKaiJt0N4BPsP
RwZta7VRPnAFITxcs65Xvb/yYPb2j5SdWMadw57FGP+duykgnrPVOGsEOX+whaRw
NytWSLKbarPr/uxzxnlR9Iwqs/5q124K9K5iFADQ8YGOq6QKw77XT80urPcqLgJY
oAscRib8KUfHuzg3fLpuQsgvp2XbLzVYyb/U6jpIkCAfGNu8dvm7DIHFZZjPZfDN
n3u7CV3XFgxdjuY9sihMvZLvKwNM+m3F15CWas2/owvPUgOOdhTkWKT1i5nPLE3Z
7DYVBBZLa4cWzvOfw8kasOBpSEv9XCIjee8fjwiuCV192dCDZjm/VyJuUtxnUSxA
EP0w11i/mXRS6dU7i+CFGTHkj1hCX6R+PHwOf77wM5YESPC30ejeqJmzxRlXiQY+
f2EVjsO0lEbspcPOTLTylrdp43qWwIlz/nd7j4SwFBIPNQCY6c+krd3G5RG2dWOb
UcrB1HZFbq5S9a6wgCsB4smmROQc3VNlxINVqYsOxI7nHy3eL3cl+l/V1K9ogCDG
bQKT6pTVAtt2HRchSIGKiNQCMjMZgWfNWpP7YIbpUmmNKa+k9H1W0tZ3tOJLcch/
PdSrAt2CVqbj36x42JSA35WGNKHlmBxmhCUJ7b3yedvfFvwHSGHKnchYOmyfBsaw
jUQUr1+hBrwwQ12pwC6ITMVSAOH81t4kqv8psWFnEeJE+79BOMQsIRXILeIHBU+p
DIIhqRTA6hFk6APhXdXnxDg4Nzg/Hf0mSOB/qO7XxBlud+kl8YxRqMAjPMrZcDVL
m0l8DTNkaJt+BRLwImtLHB0kpWgHG5gxqkSoCbfeydCn8XOJiozdNFKQTnWlXAs1
jaMBT0S1hbpyHI8ab7AvrmV/Mvha0YjQ1yScYE//m10T7mPGAni6RuVmeMvNWA5u
e9jQUrW7KlaeFYSarlUu9eEX2b7/xZz4Jh/0eE6H3NGiRQDcUSe75BKYletscmla
FL0ZecxALuY7zx1KAAT+oO2ipvnlyxu9cRJ+FEp2pWQuQRZynLtGAoU6QB1Jj2xL
XLC0lIsBmDbpJ4kbhJxz6FzvPU5Ds4i9bOEzz5IcQu9yAw3UxTg8LLPDzIs+Ld6s
SfIbehXtzoaPCYFxESwVDLfUB0FKBEuI/mmejf/Zkif1Wvunj6I+wTgdbIt4PtNL
PaA8qsbk79cm8iClZoqwRi3DmPHUca42dJyGgoj3wVwwwgkIzY8KznhXZ7L31+qK
Gtydk7IVYShegsDobe3uzfkBNwAsrpfD344K7mtebi6LW7AF6wSIirwyuJjYKr3k
qsQaRBEAQPSS+6GhgYZPyuMOh2BcReoXuPYCfR87ayOf4cEbbY5rnTtX1iDlslXX
JBZGaGa+GG+47t98ID/fSRxthyaVNy7uWyD4v9NEm7RUx1SEuWv6EvHvjBJgNMRu
Duk4yb/r9I1VbFO2Mp/nWJK0ILdb8RjdyEZBAeZd7VkiI4I2YrKw2ueNqVuWVZ+t
UKTBx8b0/NYk6JtXkjK5K1IQzedLJKQJib0os06S1E3oRlxirBUhRS6xPVK03hXo
9bUHEoyOVr7VHB4/ybPg2J+/0fJCISRHbuT8+eKK0hFFcI/Ddiom9CqN1c7kw3WA
tr76gwwI1JFWWbPJZsLXB72Z0XPsLVV59Dw9BzUU3swFruDTc9dbhjo9q+VOlpza
EGFgt97e3mPzx3g0bWXmp+OvPtusM6hHc6GoTulxyxjvnX9CfdvcnpHAhoNhhf1L
2/4IR6HUZRoG0/9VRc3B6wJ6jQjXmL7VEJ61TcsPuyOKbO8DlC/rBuHz6ngxaSBj
OlHHOBzW2UNC6KPQJG7aXJJc9TXvyiYRt3K8gwAMSX0MtKopBVj2fSJxdYy1F7m2
E7XjpOXR9SBVtAbMhgfZkSs9fjCjded6bFXm0VB0fTL7T/t3Q7tjP1tRryXs2w19
XFSkWDO6RgD5wVYyFn7b07A/EyPHKqg3s+cNvnjyQTah3IU8HdrybVrEkznQGIhr
7kCtVora0rStSDtWeEd115UAsbGvcvlck/v7CWhGSJPiEopyiuT5+wPKy4m/b49i
ZO6GaKjURETBPkFcYyJlUaK1up80MgPvIsage7fAUHOKxtXdsMiwOTpQQT98TSAP
r6QKO7NufVyZeaSgD2ao/IK73rA/M62ZbxStPu6ErAzx5eqzixEaRtlzl6lj+Er1
27AJwbLBMNsNKY8qUrK5AGtCMsqby5YBc/ZG2/YMR0I/FWSi5LDtuG0wpDEMdpXp
Ny9+CrJbME608AOx83wCYoZbBtKIIOz9/T/2OWxAcobTr+eYzIFXVKMSKnBQqIQB
xuiv21SSYIUFQt5NSIs3tLCLDYTvwMyn89NcjpXqAKlT15aETu47d2JwKvciAR6O
hPoG/ryXua50Rn3oaaAsI47uYeqqxZOl34kpjVPRtDIvEqVnIQyfdDysSCYHQf38
gMPQ5VWycMjGN/RTULugh/uj2EYkWb7jn+K9fav1b/I3Iq2lCiEc7E8/d211JhYj
l3MpilLufkP5GS6vS5TMuz390ZVrrb2I1LLT8lPvJqSM4TLvCJcZWb0IQfgiG0Jg
LFUiKayYVAakv+Pd5qIN0u4l2VxWNS9LE6Wh6tCEb+Gter3b+97vai2ZGx8+iJ9f
x2wJRnAHQwzTKQbjNo2XoPfZ0DVLm9plkLJOGey2eFDibylEBNyoOg/NSp9EJhrE
xwljh+fV9jI0Vvb8cFRtf0t0dVxBboczfdoRuVitTiug9Nfvhsc8HQ1U/gGXYWvv
JQUqhdP68R0vgskMX/PeA5sNgU5g/iB6YWBLS+YK6PKhYcq8nmHh/+n1D8yyTlzA
byso8aB+Gcz18ilxZ9dJILTcORXKrIb+lUC7aIRe5jwPA5sg09WlveJOdyCk+s+5
3C1rLUPWonT93D9+KL33AvvhFlIRSaYJCqWUJ24ykjeNP08Ap1uZ2woyrhKLg0p7
w4D8Dhsjv80Is7s8Wf4uYEns0xOc0l7rhXHxJd3jh0tOhu3ErVzm5W2hU9Cx6Inm
T6y5eJnBsOIFFdCoFIWHZO002FV8B0nDQKzTkaOKr7imQrFhU0BVly5JiJJA0AwM
6FFUx2b9nXYe+BlCPYpuiAuwRju1ptVEApJgYItpsyxL7MvrslXaoqzWy+T43aYm
0HhKAucsxoppFISkCXHAXD3fUmjUoCWo9AVhpKsZOX0EsO0ub/S/l6HkMCPZ/DLN
zRFBsriwP7Mq4Q1EHEgFEPzPZwEuZSPRK5bFhcTDKSgeeWUehiQYqdVYXgG3rxeQ
/MSryQYDfwJhnNz8UZjJYEstwh/RbV4i4j3bJm3nlE0qkuhuy4+2PSVGwSAG71SU
EMUdCXVkijJOfTvpfQCYztpdgoHveWXMZioELWPHc0jK2iROopoChFgmQNXwUADM
A341oEbGiE2wcMHlx/14ZEk0wwP4XxRcg+TEzeXf/covUTQncK5Ht5nsG5j9JkOz
rv3qoEQcSFegJ/H4hb90l2KLsegfn4xu7v7ltaIJTgboiJidHx72AuyISJJBm1H3
f60nYhLACXBLBF5A+gTlQbR3ZZDUD+QxKx7r4rtnN/rBM13PATHTBZ6q0rCmvxfj
D/W/Fjl6mW57nSemxSfrU1V4ZcSXASIhNv5+PQfEJ1eJB/Us9Hy9HEND3RdvQxOX
Y2YG/ZuDq2mc1s/rQTWm1KHXoGrnWHlKeaBUxmaY8T8Bx8cPx6uVL0C1inCp/7eY
zfUOVA/n750BYYfKAUIYQFFNYOgOY0ERRyeg5rASF4TS5HinqHU1r+bd75MA4mwe
RvZt/bGe99v6j51vy967FjawPQfucBUVtq8jR4mAmUAolLG+OmiI4LzCmtjuyDge
dZx2WfuYGa9C16pEKorSo3uKosMVUwCcJtj+YN45cKoB9yGq0IhUP4bG3s8mRi11
wQYkNe5kz5eLmMBq79wUaWi9qtBVSaoc5MlBo+nuQZUMIVKrJg/+SfK7mwOFNTYY
pYZ3WcNDcKHTTLpGG58LvUxXzFZ323RHDYvLQ/hMARgux/VC292to+3wxuQzbCZ/
D9BW7/kVGHgYcCnSwJ0GHY0MGkkBhIW0/5iKwlMc7wZaVwKhCihZt6ux8IYb/FC7
6dVYlbwpA7eK6U71lVvEz7bHD7QhjnKMNADC2ztvZC+ozrHaaCiEZP40tOTamxdc
lQda1n9GxiP8afK0UGBc5ZmpUqy2LQf2ZSVbDddamOiPD0Ez1xq9smDZCN8jpJFM
bjJsvGy6QprJGKUjszLdgaTm19n2yuXfd6o2ZUmuu9dx0z7TqAtl8WB/cCp6CNut
s1HrQkg/eXRAZ6iYNaWVnKyakxhwcl8Jh4T/uHJNdgCJU8lzTgsQguKAnc7Kp1yN
EPw7SwtNxO4+SYeZvLh6/7HuUuRP5SNsccLf5Rg5xDH7itjpUF1Azar58mjh9W3S
ym5lqfAWTLo+OeLeRrMLIT1Hx6PMWh2uXEIBScmKlk3EJ5y80MDR0XzOBfZapYup
WQLsHuVrS7MLSctJXp1cwen6b8b+JHY6mBkHJbXpHwCaQimEe+fzh6uS94numuii
pZBX+ZInOvYEg3qOIg/BStGWkVWjP1DzkBRaNk0+fgI49qNbJKsgxNmNXV3XKeGW
bK+L1RiySf5kRVGsdTt2tmEVbcmxrHDoIl+5Pp9FEkx3ETC6fGUlCpF1L8Tx//U1
eVuuh1IeulUWJBiLLoQDg6oREOS17Fg00UEEVtr7Rv0GcurRsMBDiQUQKwpT7h/j
U2CcSBwnieZJ6rGSHSmzY+NotH9Ga7NI1Cmy15SEiuoYwFTONoI5xrVsVcUpafup
353GuIkGZED/9jWbPWaUvht4+2lQB2AsGdwfmuZ/iAd0Vk0DLFaejSKteDFm3m0W
varEbpD4O3Tvunr2NDeGNHCFnwjuGAqydW8jP3gX588ZHNzlVfQa3zSwdVgWMy3B
pjEspxbw0v1piL5TJA8mbLaEpe4hfkzyrBDp5weC3t4hTyTnO4OZ1IpnmwtkcpKS
jOWahW9XLYe05fFCTiHkRmsH+B8uzmKeqSTbjOn75IgnZafqEeWKbx7PVEDnBVjm
LBLJhygkQwy8afAoZuPDWn6Mt3Lzm+V0QYuBG8jwodH3Kvb8u3gsegWnXRzdQArp
77ZTu9UIiUj/ohSlsf+DRSBkRk3nfpB5M/PjEuLhsIciUz0cdYjTbECA+DCl8uyq
wJsLAQGdwwrcFIq/blkW8p+QCntYgKDJRvGCZ9sTDxa7Sa22/T0hEIy49H06y+Z0
rl7uNDdO+Z/AeIbHOpADaoXt9nZymCum/oQTJVFNUykebyBJzaXdNY93198O4CCS
QEJnt1kd87cwpnwqaBeeYRuc3p2MQUovIXFLaAbbZsy27bbhVG6U9qj9GPml9vXk
lkunOrOm5vlpcYO0HPNoMw40zkTOhcbLYgypi3jjD35AVIE2bArwt+wtwsia4u3Q
dBs5VGlcgWQTr84gEB6CgOf/bFKUTF49I7vMB79U1sFpNiRz4dIvsRd4HcVH/ztU
yGkHqp0DVM+6UeBYNu7TrECK0MjNjO/vHwmULT3zncTikDow6xvnJT2yUpPsGEg1
PCKvWXGBASEMVE69iejfPcbbzZDOTrDE5vWCbBgpEmLNxZDN50GyE+0O3W8m5OBq
uGPDHp7bWqGs2ZKAfSeWXjog2l2Na0sncYGyDuQzO0Gu9wkigFvpf9VJ7VLEjpLr
r7Ou1z2nOa4kwaMMGKkbx/7dTtR9uhKdUruQHz4M9XkZFLDLWLCPDaegLwkqc5IX
JN+f3NHKK2+u3QZvZkL/GHBAvcS9eKtgZm4bidiM8Tb+LeQjSz0uM1v1Kya25ybx
zGc/UKfsQnquDvP3IT5I7bXANiw6uTOSIZrqUFrRYOIc3L82uStBhCjZUs1vkocL
c8ekJzAN5xsluyOyQsm09pmpwxRdu/K5xyyQZRiVHpPxNT/5up2IoYiO4ivR6xfh
A8sG/tzlA7qjD1Mq5yWOpXJVLm2KWVxuJ3GgX6YRNC1dYrY8RtIqUl9tDleT7JN+
Usp+DYDOUQfvQ3u3v71p/n8sKJrljzH//OQylFn727alAAxQM583HmL7U5A+rofq
MSgftsKxQCS7N4Y406V6UZaf46PzOkR+KW/E8oChnzslKP9Zf2z9YkW9eWgFm4Fq
kxBmdEXVKS107HQkvOnw6lu4ylGHU825o7xeRBYGi3O5v9fXD2NhMH7n7Wzh0DIq
ICa1FF9J8+pjCwrbJXyF13boHtEK1qBmrLI92ft6XlPMZgClq6O5RzA+D/BrfdFT
bOwVfMEKnuFSew8Meoou4P0GDx0ijswR7XQvxq8Kiuq3p+G3F3eSRXwpSuRsRkif
H0zKJFYzeDh9IW6bxCpjVR8nm8x+jhm5KC+sAwoghC48kGHJQxk6X80QMiSACEUN
fYKRMcabzZSaJcAxGj+dIVOqjfj/XWfGI0DOnX9koYpSvjbVIoiKzUKRdOcUYSy/
A2qeg/5mIVT44WHa8RHRghKRfaD93AN4pQukk4SO4WyTjjivjPKWGp+ucfbuOG9J
G9X3/diHWqdkKXvQwMShe7w3RMwtjldnEoJnR5XHZaiFPS269eb1y8KUDpPZ3Utw
FbvLgvvYR6fD7jnPpC1Z0MrLzbv60+grr1D6KKKpVxZp/cn6pFJhu4Rnd1rsfO1G
iXGhz66m9fedqV3bXDJOA1LlBteukdISGSDpWbXCaJv4kOmK9lYajPfFDh9kbT3L
uA4F9BOpud72Kpuj8qjLSoDxKms+t1idwXb6BGMRTVuHsr03bFfO00oRF7ow7mNz
jVrsPwBJy617/lYsGKZeQxGelQCt1BRjQ9sppMtMC0sTTR7q2CNaRDPbyZG1HC+P
wOxwFX/NHJWxD4rg4K4Vi27y3ZtVaDEg0XPxnvA1eBqw79Ibko2O/8oJfG1LlnA6
e+rr27KmsfetxqJF055N4PBdkBVieLpAW90h4SGoyL3JSn8cd6pcvX5/ibHsi3Kq
wCS7649byUcDHNdWBIZcSGwxrW9SHvgt0NlxncGmQ5NM+nx2mT0jn51Mu6Bw9gfS
fRht/qCjP9GweigoA2iwSqDgOnSxOiJUmZ+7z3xiMhXALO6BvCUBESJJo15omHr0
h3ErUqSbEnQVcyAXmKABi3uWhyDL+3c/SrwBPXYWRiT5mB7+G7Xv4z7fysIoMZE7
6DybJK1MXNKp/GWwzdTNmUmNmhfIVnBvWgKS2kSAisfvqGw+ae4eO7y3TYXznpIZ
QyQ7gVB0lxk1s2i+E8iVERkkuRqh3F6934sGw4cmxSaX93seF1CfMNhkrTme0JtB
GIJbDS7Obm9yLC4dokq/ktPfu0zhb5GKCmc2snNsuy58nt+EaewQjKWY0+ZvrgKM
uRPqD3AYozQHlemPFFOGFnMbHj1+jBBGrfSw9a9Jk7/jJvLMri4seywfsb86BQ94
/gSA8+esdKX+5Ag1C6ihb5igKM/5is6uXEvuuUU/NY0YQoMLaxBteDV3UQhxwHfn
MPeLyWUYiUUye4K28MIk88Dn5wXT+s8Z4qwlGY1G92C6VvFod9hwy6CcIDp+1J1p
qKP6f3pKgP/JluPkWiWfwh5CBbupoAUd0PdJ2VqMl6Y3csa81bPu3rqxQ//EfxGn
3pFaGN3reaas7nlyJr5a5S6EeP8RPjk585cKA3ROHjkfUpeSpqb+sCbdsHQOKSEy
pwb15wLPcHy4+1V0ge6S9foCllwNfR23V6Qw2i6EEn4iACZXbx9PhGnSgvACsxdA
oQQj1Nr8r6uhGRcnvTLwge7LtIdBDKennoyFFkBT6mt1XfppJYHbg74s5n6lQgvh
nk73A9ypsTSReEyyL6iTWkt4NRdueycE1apP17Nh2LLCab/CbfQquSckz4jyRMsz
jyqgFc6R7QZ4GzkzQD7jI5MPBfdBJhK/n1lX98gN7/gN4gypkTUuGUwKzWPVbMsZ
HCEsqEqTBOpoj2P3M5thjArGtywBy+UCRTaxUkY0iXqBNkMDIQz19KCe6Gtz8ty3
1CyPmcVZZ40ZvYMLpUch4ZWQ9j/DCls21uRu61zNmVIJ0uv0X16vcYKyXigJP0X5
tTaQyBteiq7+jBN52lorE29hTX/7Tgytn0PNpXsfAE22glQqjN8lO+z5Sc+qlRCY
ECKUh95Ag1WoWtB4kKwheiugnkozNJmSrz0NkvwfA2o96hGJhNZreM4oZVlKhqYb
h2kwAw/PbXdurWNOX4NpCWb62iFBwxn3lJEjKYxKRTlkeLpvr8lVLneRi5FV8xU/
NGyCV+CH620/n0S/FZO3OGTUrH6MeZ6A5uIGgvozQ/NegX7IbP0BrbOtzy33vot2
m5huGjyTxYFZIxV7gCkYOtm7PlpXz6a88mxtqDRS7/tFA5TD7xO9RyC3qhF2oMwg
DAa7VyJ447qNl0b69c5q88DrjmsZNeQ3bny2moN79iXzpKD8GC2+dUwYCar3l4jF
ykjFbUF7WceDbd9BVVR7GwYAlhfL/sXwYtZocUimBCkc1BQnvQxjrHTxMhRu4hR8
p/7d+GBRE1SJzPzBL4w8rCc6bJPkHBkTEAv1wiRBLriJ0AtOeBSuupXvQElwBvL2
cVL6fJmDARXg3Uxj2WGnaPxwybWsSt5/d/eJU3Gm1lAQjiaMpANgVSy/UlxnQ5KX
KcI3Z6M35qAI2SUBSPrx7xplfNo+ikxOvdcThBx6GdtWmXUgHs5wM4ahRuwE2m4A
NDl+X8ATgnbjDWASwKxv0bPPnTA7/Nb/8IOoKEXXAhZgBaEPcZk0vIQcDp2kkPxY
hamOZVYlHQPSQEnFG1ywCmKv02t9jWnrZ6fnSy4ySnuHTebpp17s4ZuBp41c6V88
rTUdrmr/U9UgWfHnac/gcTzYX2nKn183/nBpKqOJ4s7xyjowMOn3HLLJP4i4qnqE
fBA2Alu4pbjRPwLpCTcl/OqKv7m00fBJP1HG12CcTr4OSw/ic/lBJ2o/2bpmCjcL
6Ma6tGiewCofk45tNMq3ySOX7WXuoV1l6jbg+WzMi78ExLpA+PZGqu4cZDQcaDdb
GEnz/bwwrh7va/Ltyfiv93hRoExAyZp1En/Df3qORb0kV47z6V+1TGr9ckID55Jj
fbLrgevUbbZ1gBHcaSg5RmAFLcwnka9qbwJvTEwuKupY+npmKNbPS0EhEGDOmOts
d9UjX8KtnqRhFxoKEMDFTxsu+H2qigLCXcL615udBr8LODQjknmdoqVdBYPlpU2J
JcdvAz2cQ6qVAJgjf8YZBoYqxz5p+uWasNwh/dEIZPB/pf2L21gcg5gnXzhC+FP7
WaLy1cdZAfNIoHSLM65nDMOmNn76BeaG25rx3matRoQ1w7G85h+RTZNtdOJ7NVNt
2tMq8EasXTIsTDgR5Tv2IKWzNQ6dqEmjPxmT+VahC7OsBd8d7kx9SiRmRFzj+2xp
UF7dfWMdFPvRpsGldWDZHmfm/+tZ7lU8GUDM25d9jq2yWGOOtsY12pLl0x9s1c5Y
JubrJBPjWilI7kqnbOHKfE+mYEhlat+EHt4wq2O0DWAPNnAM0LGQfpbyIYQ+Cqz9
5gQXnmk/Ob6qx0iAXtKCzRMAc/BccL163Mip9bJVndHEmHkfSn6vkQlUq0GvHqZq
9B7U0nRJ76K2AZ7M3DFF0u/pOd4nl8GTJkx23qaWbdfNsmcOt0XjPrSkR6coPHZ+
byUE60qlvj+G7NSo0eXoy26XF37fQxNSlzSGzzmbOWaZUq1yTrLFV8wa9a1wZnWo
CZDywBDs1uJxir1oyfj8787FWdMNkSXubdXr8z6pB45asIjpBevwpKf6oyOBfqgM
PEIwFpO+bj1NpUcJoS6sB6wfsZbnHDDJWQIGtZMyDpw7vOTWgmssboNaKXmS4g2E
NjolgVYuPh6FwIfMR6HGSc6SgPq/jVf409u8ziXqsQTGKZsgSUH713XwgCVyysyM
nPTmr8ZmtDKntwlBXiyK0Q0qCnaY6zZTcK4a7WxAYzawzoocIOKhE9NhPk1BMUkO
2Grpp/SrhIGp9O8G4jI4EGXAa6wsYkGQMyNwmIgFJAeydLmerxRKcIwVDo7/9l0X
Egdj5+zFp7FI+IUA8vW/xY+zgtfbwZuve3Jld5bcHKKBR8A6RtxEvPfhiMIb+I0y
FUm6Oa8r8HU8DUeJJ42jr091ASJXPqVklMWckDWoQYgYwBaif+qMhiZdCMLQTxoo
+sdAm2RR9nvOi1Hua8Erx7KNXxXoOhgeZEI8C5lmZ/jLP1r1jkF7PmM5cfNet2pH
MTSx28j5vCO5FliyNR9xg9a2yZy6MNJvFEEHnIly3Z+dk9DGVkLO10NIrsysmH9J
TML2cLiaEQpQa+YKzkSoOFkvB13m5WjhyrMSTGRWF6KCI1B+a6Bo7WW/5ho0AFr3
eqhLv6ZJqTv3anIRQu3DFpSffeck9m9OLC1Keb+8AfWF0+FHfISL4sTO9y/kY5LS
1wqfqlBVMUsiGBaJ07VmMU0gHXHrVlHnal7xnZjdEoHM8Kghikd54VJeUIs37P+M
73gH9+PT60C0rP9WCDmWM5XYM8gAl4u552/z6Hw61XK4dft6Otztac2WYd27BSeq
9Dwh03PcaKcVuapIsXC6Z8beFdoKzL53zfi47mFY1i0ZLKkrp16+1IE2nF8sLJLr
gVV+uIo3OkSr7XImsg5XLUcqQPtgf4lml1E6zp5+McfH/DK8CUfHnOis5PGM5eaq
9SyuHecAwzxjGjGoEtv9CQHa69iuzc9ctI1Yl/1BgyRfhlaHNWntV9RcgvIJPR96
OsRiygSu4USm1eEY/x1VjxPeXvv+Tn2k0SCdszowqsnK468I7y/IXhgG2UBIq2GB
D7T179ducIth8fB6HwQxlhZRqAIophUYiYiQ8JQQpP79QMF3pMEs3uUE26Ujr56S
Hy2Nh+xJg3YL1TP8DtpjIDhgjHvO/hWyk4tSEY6bGBkXd73ib3gyF0vond2arb1f
5A2+rkIv84Un6nTMLmPCHoK5pZa8nQwZJOqiX4eiiMlTIXXM5fFhb8/rK7NQS3QH
IEYHvpMoMDEsxPGP9gmz3e0muCXO6admcbsb2tSbsZ1ldCi0DlDDSZrK22R0nOlY
MZ3YxgnQZNOAXoxsG7xHBwySvO44AkShGfbxvrtI3QW1D1dOLQnYFbeHhFv/mPIo
U/1KyTFLfvK8zHXnA32N5l4CkWNBMpi8Qa9ymKF390e+cvhUoKD3CQ9LBcyLqTvM
IB9wcC0SlHCY983XR8iU5RKuNyaqpA1jiKBHd0fO19NUOW35/8UlJF4ai8nX7j0d
J3p0EXUQdldncgNbIkogrotiAAkAzE8mFMIzXRsqf+NjGiNm0lByidPf5sh1ICyt
JvDtZZ5YDFWwnxVLzXhmroI3ZC4KGR3jJBp8XW7Zgj19oIbvxLl0uvef4DzCD94E
GQKvn98+lPc9oZUUs7SLGK2WO6gzRpduU+7t3YM0LzDzLB0nBBmEpmNPxAzWupHL
SsHQQwC0aNZ5Mvym7IOGgtGFuf9FWZIXsoW0UMxfFBu5AZS+cdmq3a3AW9ctLOzm
RrB3gt8Qew3C8CktW7aOU8CR6vFALcZeEFkfdw+lhuvyREKbkxvtqVLY2sUOSI9F
mw8B8z/2w4x2bcK6xzhxKENFwpFV/juND2oTXXTqwsoviJG+O/JD6JrFxFFc4VCX
R3ritRBsUJ6nssHhx0j1x40r4KIMeA85UV5fpUSgA3Gr2RhPRMyeAl1OwBnjFXAK
DY1EN7rijLSWvF8bqA2804ea77S3S7z99Wd9+UkrDlPnEC3TuZ7mrOWAvI0lCNoh
HbAaFBL/KIhISrg/nmON0KjqMdC3KxFO7uNNX0wPb3t0t5wbeySQFy9OUdBAHk5m
Dh8sjrnwBWopFsBRSIZgB1+ebs1aXlD2Ab0uJxNyAmvVAXq6llL+IsszoxgkIfLY
tEsYJgwvC5WjJE6tqMu+AaGCNSI0cSD0bnNTalSMIzo92vgOlVsNWWbqorYLvFXL
+M+VykiSDJ6kqDb7TuLM3s9gjKKo8G2pZgSEJO4mFDAg58CKbHvdHAJH/xiwrCSA
GwtmJ4UH214m6vCBvqnFr49/0BVbJ6a0oL8A39/OMaOnshDzv7sKfBRpIvc8P0qc
5e/Ti7CZQhojYaaY349rbcQaDnEqdtw0Or+gxS809x+R1EcIT7ub8EkDYl8fJKE7
JQU4lR5Rh4Gk5c9ZMn+XUJIb7D0hILWSM8pL/7jygGz2kSftm8M+OE9S7q0+7abC
BP8yVJ1/PMOmmWGIdhi7n2kmAMMd1FRXcZvMDtp8Fm7UXmmanCWks3sJ1WqRwaFK
JRlfZ48KWOONR5eezoLyZXAeW+Drpn6GPZuJ3hc1y0hVr0JNqQ+GCHAMddXT5Y4b
xuAttbZ+NHUNGCOvHWVSPKXJ64x0DOCMkSkjXmk6+727VJ8nEstkQn1sh4b0fFEr
vgrp3Zbyw1guRy3kQBpBD4hmIDkZIoMPpQovKNf+xEkgx+YSoywBXYF9HtclK6Yt
OOgaYlXhlHg8KWO5mmIkoS1QzM4wrN6esJXc3d65n9HvtsFjy0cdeauAz+2opW8X
qq78v7JjDQHmuhaZPcL8g3sVwrzWoNpTXm69lXfekdHi91ojRezFnU/Ao4Uq3Jrs
MVE24spFgzjqBdytMG4Ecph+WmjbZkBoO+riOGHmt2ABPMB3cGDZWp+hUgo58YVm
xKgiAmitg0gTVZuIOfwKE+qFjvAt0TcwiUZP5jXuvpmkaxXovN94PCl8R3vNqY3w
O9x8kA5Mi0nR8mkaKjPBp+a5kZGDVJV5szruQJKqdnVkgPFNjcCJBjFLjqYRh7qf
ctNI9ugd6mhO05Fng9gCjR8+vFBynItVl8qRXe9lHJpXBCMl65KWDGl/WADk+S3r
pYcF6n6Nq7kIgpQBYwah8/LonTZIK6YagWbHjnPZVcavUo0qwJJ40KmoIPw1C9i+
ynJomLTkqoYPgBfHB/yhijFo3YKSbZSpMpoviiE2yLzO6fRWGetnx57R5Rlj8Zux
Tef8jIu5rVZjxnJjQha6Iojg4OdjC4VgasySRXJRq1D0j1Ct5eBcnLBETSf1zfOQ
1cehNtmzB6LMkF+RYizYUyAWTqVB7bGNdYPdjyDAZLcwHRzs2ZUumTyRtLCwCluA
EFhnaru3aCkxcaNERZogw0vrrTuXQ6pB/ym5UZqi1a5dxj4CRTc1CN95yTtXLbn2
w1zaElC4gQrpGdt3mlMNVKaX1zThGFWxmCbN6sgLAjuvn2BCkyWshTDt7+O4dIWa
GKD8ElqDZfVvWTHhnE4LoBvAxrvUESszHEYVR+jaX5HyvEoyS93Hz4UAsP8hOiai
XI3ReZuHXOkiaIwYxrekaaCqW6mbKPufNCopbTljLPUuVnVG5W4/EnKtum59MW/Y
ADcxK2UfBG1d0MhXJiV5DeStODhW3A7ob41iMZnK/7oiBvp06TnTJsMsvcVe2PPO
Tu0kgslgdQ538OS8CoHblp498WiN90Zy+6W0A0K65liIixdZ1HnqvPxYM7TlwJAy
ugGH61kPjCfVoi/9VrIYyhBJ3ihqOD5dvqi1Fx4sM8wPfxcAX+eSvQpmRcxARGlX
HzDGORykoWzT4ly1RON1UF9jSmpDqJbf4yS2J8bi+Dm6kIn4pAc9h6uWHJNiW+bK
Uv8Jjigl4NVzgF2ZrqMIcqNGdJjeaEPTo1mwLrSqcfhybJxwm+KwJuSjvWhwqoBZ
Vz87M2f7H/Oc48fEVq0Grtq2VYkqtrqUjZ5EtzzvaKKSyUJmwoXHxaRBWG/En9B9
CfVSIQnAlfTRUKy7hGmRr3SM8/7/BJgB+OXOV6A3DtCc7s6DeavO/vYR0sq7sFzm
Pk+b3YldTHLuEFHG/WSpVPXyPDBCAYcyPSZyWsdYRSxxTylDc1vB92K94okbcd+o
bfux6XXrNxuzg3ZH2tJvFYraxik0ylMSPlzTWpgUHQ65ZDRZhNy7E/0wHzkoPW4X
wUm73pUedJxhTEoigSJA7l7rHo3K/VQlTSC/q+rcFgPU4Yrkmfi1P2yqIIumtTDm
ccqQWd92vLDMkBtawWsUk3LLkcUbgoEnPvftiR6gvtVBDh1gdDkaOEiiyRD2ooiS
vfXHtUWdCBPO2AAb+RQJm0LpRuHfFNra0km2XAJQ9k8qcbR3l8DUS11xZsUBhPI4
HbcNGtRiZNDEikau3z0YiYkeg6rgn8qhZV1y+ZLBqS6B5gHgdPG+OlCgr7Po9XRE
vTllp6Y/mjcfVnkN1bORM4ru1RKdcYRhb1+bQscPn6IXi8jS7QAc8WeBKV7AZJLD
hibyKzK7eb5JvVFfhjBNqcHeZgaYyUag52tD6pPH9vsd/jvAgEQ5mupVUPCnqI2q
8e1CzdLB7m5TFNUrGI2G/OJ4+7I6FbJ5HPWqyOexB1GRSU9whi9E405Enwcobksu
yMAUbVOeFlts40PE3gwCbcJjRgCxOx+f/XHrAKTTHyn5gwBpa1Bnxxoq1YbWrqkF
6y97z31w4bXzbdfX73ZL4SWY1bxdJRrWPzoXq5B0Kw9p5FTcDm1NSODjRygQUjCD
b5ZJ3vUlbENyaeThbv0UAXfb8zQ38uBh2k12mMyGQ1l/L/TB3rdShh1CHE9o3+qL
l0Z7Nec4KaiHalF8ItfJd650z75MKb+rOEbYJnjHS7XmbiYhJzTBpAT+FpPrp6YU
8vB8k2yBz3RVr4Ts12PYlq7rjOZLfQlrd7+rJuhkinjzhN78vvcnEfvZYgAj1Lrc
UfMiDaTwhXNjpxHGdoD4aRClK8QZvG2FNGgS2yzprDuvNA98lbKrPMdyAQdcNHOO
0HLIPaP8wMXPFXXdKhMAoWZ4D1HdcpHqw5hjV0hdpw/BkEagRHPAxHhkqiVJ505H
DYvW7l96rbJ/Y2xseiECYh0ou8sTv/B7N5Mb8N679Ux7HDnx1fW+BEFz96Q+Mv8a
+7kBy/rIa3fpp+BwmzLl2Dx2O4l+Ohc7UjADcBedcqtZpXLVJeQ9v7iduGUABt+5
3StigsnMMH5I6BdUJPwMa9tGNk13GozRS+6a8nWJP2/Cwl128KqAs+o7ZUw21Z1q
sEL8gk1Pyx9pACs62CEqLB4JUdWfWgRW0666QdhKtWsvo4S3DPvfobZSO9y2lPQq
KIafot5N6cdGS8ryZfBaDk4hd7QWaxYuJ0Mw/IILd6GAf+rTM0g5Dfe7hxqa7dbB
lMvOPWDZ3tDDBTnFTDGFKfXMcY4uGjYbgpBwNX4W67apB7w3gTii0xGGB5lGKLkS
TpBH5nKkBh1Rejqgrc/bZ4mqB3Zcb1QjjAXDI5s3QHlbLSdrKupmYvF6NT0s+uY2
AjLBl9o5qDJ29KWghK80zVqi+hShgRHfctaCB71wPpW2vxMRBVFlLx6fcmH1plGu
3bWAuf8S5WPzUOr6/Bh4J9oFqVHlARkKDqaESxEbNyK/5d4G0l87sO8w3ydMWugx
dyd+FyRidxFSldBPmWUh33kW9mqDcpRx9iqujeemqcT5SHP4JsrWcHJCVA5RrShT
eWvNJCMOWw1mhWEeZRdxbspljzzSt/i5Luby/Vp5R3js+qTqL841wwxYoHftbfDT
2JbmndnBMf4CfuKIN0VXkSgz+rgD1A0IZBftyK+uxCCBcTPP6nu4vL+wl7YAMNrZ
SEL9I/HN8Ck6F5KjVTQtlMsqElXmgvGbeATS+RhTQX/Vj3//oniKQSL8c8HZWl6c
Go9A9JHEa3gCEKmiZODrvQNvgDBY9HOvMxVWgpc/M4WDsEi14UiUgDiMj5hNp8ow
xn8emqa6ffbArbxXkk0M9h3Uz7vz7dvF/nlzS5d3dnu1pa6UQRFhqlEA3QBCxFSp
tYXWmbfJKfK5yK/JeLKBrwbPDJQ7px5Rs+xSraM81MOurKZ8jjJ4e/vnLqzHSCaW
EI8IeCribaawEQ3M8OthkxC+yk9X9zVwEC3r238/2MS6BPiVEX4W6qTdlamdxAvB
c7mTI7kv1CxrYvp6Q9V290x8XrS6KnBedgDI5eGx7nOBC48OkOJoA9w/kmJFioQY
m4QM1uJdrTtbjOZ9hvqp9aH/g2zw64Si1cuqegcTcpw76OKAtVrIWbn1UItORANL
kqwxlX4WjpheUZdODUnYlTLqFV8CXk6KtlcXLNVxrUXrjfRJxXJ6C/Up15k1Q7Sr
dMn0v8yE6UbZP9uUTQfQxC3/FhF8NJNmwENO6d9XYfJTcUwHZJj1iHLqdfHmK75N
x7SqpRJKuSaYlnXB0QSq9oxzIL8VY/ZQCGEcS91tG929Z7g+duLIM87i2+qS9kZt
h3mltZZ7YJhjfeJxw0qhz0D3XKLMl9pRwkcd0DguFVJwTxcnQDITZVZSSPPBv2Ud
MujxcLwZVLv1/M8XWeKPfTH8g7VGwT6rthn1Dsl1rSgBgV3/w3Rk0UgR5HzhFVk6
HQVpntVXKzwVm6u8495+3bHjioWl87x5JsJv1pZqAJlfFBsrhvsZsr0JwV7Aul71
Rk9oPz6MZV776RrpsR9MA17lh4cpiwGtDAt6S/vxer9d4Nqr+uBlTxmQXS7xEw/G
l3KskdC/RQg9dxP15PlFBmOK+MUOCaJhwi+SVdSiUQBYBBkCqe+f+jadTdNTaVHJ
yZ4hZrZsrDaDtC1Kj/Uh+FDfHqD0pYwXsfMOrFCZS3ZsWQ9Cm+SWGAaBKINhxJBi
Ui9LDbb50jG3rt0sAKRXq9cIzSNzPx92/KpO+TVhlkObk4P4tFgoc7TCzDkXRTrj
xbxtPb/Q2d61DBg+cbzO1fF91XEgJ54iu/VfmuCwxGIKYLoIcWt4Wk+wbAdC2PBr
Zj4unCC4T5rrdtUTGqc9/0y7VNeNZ5lYZ4m2ZBkzflC4EqwZGxnervfdsIk8AOyI
wu2aGupJ7AluxycvSHn/+pEBoT7gaUk3lVyr8KS3LA3C9UaR7AbBwnnipmOIuZgy
5ev3HAZ7i/ZACMJEYk903yA3Qq+kVGYzEJIspjhTp/wbwnDNaIO7oJtFXaFjfpPB
4FnB9N0YQanZ6ds8KCZSQoO8kkEcD270Z9jGwdkmcWpPAjA5+PxKiLfcluKA7CXJ
V/IiTUEjwPLCWzq46/InV+VMtnSUuOnVfluNg9O3PbgIiwjI1QkSbN/51/HxEPmP
zyRu5VkQJu3Z5C46F5kEic8TCtB/TAwq9ipo2zBNCml8bXJ9uPjCQLtMSEpUm8Zg
pc1gSqoZ032Fmf9WrC6cC3b75m3t2ACbz4vULriwdTDNRHK5elI3xSf0INIWVab3
UJqAfVemX4jmL+gHSIlA4xWRPHO3iSFUTNxLSDr2jxcX5cGlHSXlnP6Nsqsb7Dag
/PQZIyiQJL5gMxS0rM+XPdFYWDwWfoaq/J5f7PPi1W9YzfLoB0AbtiyPpWBXEeLz
kO83TDjosRUanCsr0u9CjxSTLa08ilBIwZ7G6ZgoYuNo0UNxsfkgqSC3dSs35xnW
5qLoVX8wDCHgKv/+BiMAigVc7+Hbljz5hcUNDLmVpvFKRAyACUwnxFP2XrRodD+8
VtVCr7tVGKxHv7P6c7Gpy/OvXqqgSQXd7TILPGsUkDO7H1LsiuuRr4+fb7FG8oBG
t1Lwm5luC0pSGETLQ9BAMhTtIWogqe0u2Y9djJsD3LGm46U4+uk4EhWN+N2tV7Qe
E0GPYnQ2JabwF2su2bhfJjiSCcDzPFZCmKBq/lVSb9dAZESsUu3Z21fC9MJUkrqq
XUNEl/Kw78k0DcugjoQV7B0GJz7QQ5zR7lJLtUalxDMjymFZHNb7N7WG+TdV2ksa
6AIt/NlQzF1wIkytrXzGnnf9FbcIul79qPEPbZXRR/haAIZu+9yezkPh0IGQ74Ac
s/+SAaypwA/IRidLr7JP9vw12Vvjich0gHzzXof9O2jTgC/Qs8qVZWFskEcmiLrb
rGaTZa+HV5awURRhE0jT4+ZrWQxZSFbxxYU4DbmtP3CVsHF+TBcuYuz4Law+Yc+X
syk41wrp6nYoU+AOpDrFdanWmMKaIQS4P/msNJKGu1Ef/giAr0dIcw+WjTeef4oY
QFdS1VQs8A1nxXYK+oqihu0nkeirxnxxSj1EYZB3UVs5d++96CjQSKNskO7CPJAA
2R0v0PRbUoJ8jWKIr+3IfAdfB3uY666Qm+drnV+s3Hw/DY/R1UzDkYtCN//MqepJ
3LvTiwQdEUaSnVB+nbRepN1LXL18+4k62i808VxXqqXbWddmNAkRYadTk3L+U5I3
uJcrOoEJ8WLBcrsvLYOc1iLJ3E2HoX8X/okGjzLyD5Uh9c2LB0GnU+P1Rvjs2eWX
Edep9iuEpiRBgChVcith/VKMC+a9WuCIdCBUPBktwZBDAW2gzgn8XYBfTE6qU7lJ
Bfo0RJiedkgRSAQOZTU+3r5GIs/m0r0/6H/2jJ94bsUe+wIOSA3GfQyHmC2a1Llc
lJTnFIBJiboAKc45IgXXd8gbQAgruaHlZwxtLLp8JXV/f7zlDPkI9tbcbmPQr6r6
J/ZszkThnj7vAddalCnlGaDT3kLhbMyC/6FPEbZKkBdEm08WQbTfogLAC3mO9KmG
h6IJHIdSS8M3+qmhWLGjXDo/bxLUkGic8H2OHXOeXG2r/K9ZfXi/fgRlUITVYKRL
ymI9gZJlV2tSgsRh9QCcrs8ftUl4GFS7Hu7l/Mp/dJ6emuR8+9XTV2wybbjlMWbb
wptivFdJXi5c+woV4qwlCDvmdTQZWw5Bxzzxj1yebPi90RtdKywMz0gwW0zRidZa
jGSiAzlzEnULfnJM7hO3BpaeOZjIeNgkAZczK2gAlCWjyndl4uYWEB7hveb4tjg3
C9EJKSodZGxJpr2hLWzfid98xozJmClQuHYXWqPPAnpG0hMgfw17YFuN6a6WkxM/
CQu/2ws2Hb68bzrJlkpZDD9jKSnAEnulRvpeT9MVGPVVWgVVhkRDTTFkp2Rmoi+g
v0Fu41wBneURgRQyxXP0mhDzGPbhGLgBFKgwv/ywK0rF5dag/cbs4iEtppImeJd2
83vFTGPnCRd3YW4EppXn2XmEQugD61OPzNsi5sWZiIVBDzkWZMQzMiGCyuVBER6P
Xorg3ywYiL65b+XsG34F1DpVHycsatpfeYe3XNfOR+yHSoRokKIdZWS0XZr4uLft
EEqtHIR8Nc6i+0a/dZU+Kg8pKB5Wyxx5wappS1a+aknQcn/Xc+/TMXUuefxMkeAv
LGcReDntz0fvHKesvf2+VvjLTVWZuHQeY3DJFpcHpxQz4GEbdGPZtUQClCddbAWP
UssFOOq7POJvg6NQbHkUzPl5qk8BSO6gjdJKY2k/EO04cNglhfloVSyAmVQ2biom
MmLiuQ4+uLJRFrkZEVCLvsvZeMD13GSXED0GMwLXDKpw9Hme/EkqXN0QjtGgIQmi
yciem0t+iMjt0zsLLR9kNEmexNqI+6glqwD60RClPIv5RGrLi/GZIgreilnjYyeY
TfkOT5eZx7l7wRNudHQF/V+tuGICMFzUcWktpPXHcsK7sjWES9CwVjTMdjtwkltt
eb5deRJEidVKE7PqhQSEqBD8SnAePhiuRPqJX0BzQLn53wkJKNSGY/gSAt6qjmM2
93ykavap8BYG79ESHpySqc/wRDpYXG+no82x4H8fL9qI9y6SRBIOULD0895G3P3s
hDZlJGPHXMdBijf8QVrt+bXsAUmj930PV4wwn+yfodwPbST70L1QESXJ/pA0hO/z
4bXgWyieLzZlB0eHBomwBHg1aNDiPInZzUf7ueyvRmdL6BPWMFllpdvWoZRgFiMU
vC/i9qPSIG+3sX5r6RRSmC5kLKeFEbSluB/BMIuhQRO4CkAPZ+acf8DgIUB2ZiZ9
bZ1xG+4UA5UV0lWSS7J00iZ/saFLJubHfjKA8dbYoqFFR9gIDCWtOMvAtL8i8dpt
nJu/AEvv6Xs7OsekSQRKhsZYjV6WxtGq1GGBlJu+ylGB4aL666p04ePzaFqSx/hN
spm2f0XT0rN9Rv1GVn3yQnjZek3wZqFWyu8CvaEsMAIKrgyjA+My/UoThv+7athV
ZS6swKkGDpHKwixuUC5q6MOfElroaRkLhx5DsXsGDODAECMdpsRIbBS9GhIzeT9G
nBbh4ig6QuIq+BakKVOMr79Mh6JXizRT06w+8tWiSyo5X7w1oSbCq+CHpbBnsbzn
yitWQw9o8HJmwtbO/L/3xYuRkbIVjc21kKHETXIQYozyU+SnSyeHT4x9KNdbdw5+
r8vVPoLumOgzPkQNDl8LnS0d8HPMXisZL0PWq1SexnPGyOwpqu0IiHv3zQ7PjTrJ
T62qV9Ui14xhxmMhrXYBE1bOLcQaiHXsi+YBjtAkmUzwKv1XaLz3YYHmgb+gnDnB
ZizWv5d9iI/mMXohOTjNyeeg5E8U8q8auEE3jDRT0km3spuk+NEiw0nr6Ct/fd2a
IycqoLXAW5fOomyDjJuKp/WOnzh+xhdRzwKW0Jy+nTodIL9xBbMMCVUFN6yQVL5+
lLybPbNft6Zu7uP57I7Hpi9bpgkyNuG3gL6qJZQDYETYwHSjM+oBp+yi44YEW17r
tZLSuZanXZ390TWwM/3xF4xYvltiOW2HbhrH17TxuQ1grVNIb6ldO5ktvHeAanCZ
3okZmCztNRKNA5Nmv2UBoh1fl6lomoDD8iMhJIzCVf771uH+Vhph/eu1LKRUO1gv
/LrZ3seUnbOfD4rzpN9G9+bTrInJ580Wh6fdUveW8D+5CRAUsTSHMFlStP/fbZGB
qxAg4N87aMCm16/UxUBAvbYkfbHJ/T4adS7Gp/ih0og315uX47jRWz2FvCGDZ7ET
Gi/quxIBrUrnrCVpHBDf3556bG7oXwvcX4h1bGI/r/6vDXyu1MxA2LwYAKFhD3RY
zCHPAUM6xfL/doT3MbTFieDYzAiMeWgfZ3Gm9COfyXMO51Uo6ZZSb5DYyausLZe5
FejzcEGYR6nkPJuiiL7GO/jfD3b9dmZFvYiVzQWZX5UAXBcAB1URkDYKtLoPpHZA
J7jGOmlrpzZhpmJTU40LMxXbi0MYfCo3wwfPaWGZEdLnjKI972my1V5dst+2Vh9J
DtvZih7L45vG6Q1+x9iO5rsF7mFAN64Ai5Yk99TqOxqy84ryH7qwU1JBeSFewC8D
mFWMpzFvmcHWFpZiXaT8L7ffQnOtJPn9E7GCD427z0ONt8smzeJ50oICExqGV+d2
XzhlFlL38yUel6/RkN3X/R07hF8gZ4UTyMtmAEPsqTSLnqkRsNx4bt2Y68ARg3Ad
0sSnsA8642zT+hA5RaQRhK32Ch8kOyQAx9Zjc8C6e46/nvU5zCnUwDF/dNn1WXvc
DmTySugwrXwKF/LpcGWXfoNgKa8TfI3/B7OJrV3rAOCj1IN1pR0Ybxic7XVTOiPW
JSLBylIrRv6cl3tR3lT4qmZS1aNj+5FMHPwdqVcWo0gL4Cima3/k2V2lj5rdgl5h
aof6RfoIqbKxoXSIwfWVWQJS/aeo01ZIfwqiAy+aWF3RrsrmYEB5uzrrgWVTkgDq
mJ8LTqqiI2Lf10L4zMtRAphOsF4OEzqIsyHDKST1cBNIjvQ3aBMTIUaukwhpSK3/
fTo+X8kaWekc7RlyAgEeRxMN5OBDh0/NsmcvwSZE7NDXt5rIjr0pdoBW+Tba9+UU
rw+kmaJLWftrINi2vSIryakDta7Vm3l8WdWsiCi12SUJkrfunzbACoPH+GCr8ZgB
p2SGOvjaN1XCdoF4x0cZbehuyhK/8Uk/hZ4PQW048KnBhh4ZV7uqMVqvjirs4XQB
3IYfMPLDSp59+fbxFlrh2fKnyQ8kaY1SSZhPQruml7V+39B5M70xnS+TzLpv11Ml
HgS55WCAHs+NVUfm4E1fv6cyeDR4NPjKm6qLsfzCsxsOtiPl8KDFDDzwOn8uw7z6
3I6ZYT2VicRs4nkn/88ITVRGsR1s7kbVHRn7sJRDvOQ4/k6vsQ4+1yEfc9+QQxUn
SHtBwVvuNVDlGdJweXU4qA7HFDQPWqQuputA+x5yR6twJVbOGh0D/YllX3sKX29P
ggZcXQWedhPdMsLdj+QpHeMrEPKW8DYG9p3sOYoIYp0ONxt8nm1gTeQFkDkJJMKE
cajLQcXm0iIIibwgLonBDmEq/Stj4Sm5reAZ4fcEWJeR5jh3vxxQRYoo8afk1LY5
WAdqknVBdfoJLLG9JHqTRJ4pcGsCa5zPhVDHEFwRen5XuDh2SIV4Rlr/w/dc9Pql
FRXtzJy4MuwoAkXtdLyvMrBIynYJw1s9XfiJ492Mm4dqP4h039JfzC35b0AeyfPa
JTsZfQL+6RJAxsS92lW8jPjYki8xrbIHl8/DzsZh1n2awXhgEIu4yT4EcPyzGXHe
5WKiu1rHZyRZQxxpfALFJtvw4sTsF5skTLisVdcRhtMih45Z/osuPLSrTVamU/lt
zizIzZwRJCpezxKKuyX89XsEahP26xaukgVQxz99CaCYHvx3D1Ajd0T7iJqv34ns
YExUdmJ6YVnIqufiNTmAgV3Wvbk0FsNPcb9rIoBlfPts/76v3qXOhHP1fexrmoQM
umCr77dFSBcfWqA0ib9Ia/wtSAwiQqI2Ayumo0xEpISwWdQpJA5u2OSCrAMJy7qS
/uRvx9CyUcN2PRRHKo8nHN7PaGv62Sz8wfYtK99ryxMQ31Tog3hP3yyz2H/miuHB
XKuPVI2QBzRelKpAnXNj7uJeMAOPZ24aOZDJemrwiktOQPmTUp4697kYZWh6hPDY
1+6gRSJm0YDU8NYn4YIBJFtKd4HjK3RL3zhDtym+nd1G2FQa1Nu1Hz37L2A1z85m
F5hpw7Yjg4CRxDj0MTUQBK6/m36tmkQ4tt03+mDnzyiSWsBz2sGMttEql3er3vUn
vgXZiZpVK5S7hgKV062t0HeQYLzi3dDTXXI5dxIIb2ycFkNvfIusSpjnJfQuW3DJ
z7BxxAUdnsbm5zLY8LnQOCz3oIjitqp4ut9QwAczufvi9FqdgURGK44zJ7VGPga7
Sc2qyIrNJjqAdzl0EjSJUUOF4dty6g3PNj09k7Gdn51m01WHPxZIrqG7I2Yp/akj
R6KPFmc26ev5RnblZRMj3cgvbU19H3HGtyAbyJ5FnflqLClds6OmQ5/7nlahrIQJ
kgNN0ahglH6Un9rYDOaHac5xdZyNiVYRabb3CXDO1wcjBEFFTxGAWjW+WpyKgKTU
5x+M/d/DHh8KZeHZ0pN3iRCHK/pwutWKpMhgUu2JcbJ5h0Ifoo3UzdqyZIJPuI3q
rIJemRZxsq29T6O8i21t2r6mFT6cmricf7Oo9tgjyRtyTAfx/o21HKwRM+lZIvlo
Y3Aa6vqbhQgTSh8/GvBeZrYUADf92Faj3ro7rFXho8nZoYGxg54Bk7KG56ypZMde
3vaMmSQShkkI/1hstd9Vxbr8NAkLfYREsEp/PIiN9sjHAGDjstFApAdJIXvHdD+E
YDC84WostspO6WdENOjeAnEdptqJWd8gGuOs+Y6EMBr3aPUG7VUySNpdxbj/MnkA
D+7g24UimSBqEXlp7NnRsBzbDdDEiEOV82lm92dHo8IqSLHkuJbbgpfR6oINOf/j
Eg1ZoAR6z307xfNmOet+ZpG4PG3cwZ1Zh6CqwrY0Ffb1IgbBWef+LNKvzRtJfxXT
79HS3bfQK5D+ofM67IIzbm5Bo/6D8IXuL/FVZrCtzYDaPFx3QLkoJmruSg39eLTH
50N9Wk8OXNSiB5ZjuxJ4PRFRZUHLV5AhqRf2ATwJu4Hi8GfG9eC56R8IuJX+H4Sp
h97ulX2IkuG4F2gfMbSt3v+Du/mvNVbZy9WCE9HBE/a61GvC4wffFbT26oQRDi+p
8QCEmvQS0qNb9Pzvond+2cFb6/jgOZt7Yi5K9hvMJ2+bvUEAKZHp/+AoMGYGqg25
NXFpd73wUcdG6wwga9QUdRgaWVTPjdwtbK6HAJ2+Wfqqh1EeCfnu0G7NEx2T47r/
B5haM0HNvI1+KaF+CFYc/BHY+5HrXxnbISCjelRo5MRUMkUS3CeQdQnDArXpsDlk
sCOFyVZ3NCYhmrMpObpq7cOguxqEhJGgjkWYtwA/4KaVuSToHxJtUtudwpaRJ0mK
aPpDe9OLcAGH2V8Y20Ij4cf834E5H7vBpCliokUBKAN1g7F4oI0XqtEAaNK6jCpJ
T+j1H7YbhKXh5vYvdJ0qmpwipVlRQoL6mYqXW1yXJqLOajDkBAoH1H7yWu+h6BSh
eedvwd6oSxZKv/i/j0rIeXRGxvaVREAdXqcxZmjkc8ash1x7mQdxtS4bfT30XH7o
5oACmPamGIyE+0pCnLiT4RTBACLIPqSfpPIdIbkBhqmI6Cvdp1VdWVzoHk5v8SDR
VgkQ7Ckm4YlSe1rVQlr/Pccg4BSjhJBQVoq46zHXa5aC7wuPOYt0Q+Nwkc8Uoe72
kHzD2ntBcH8WSh0Tpa5pFzvblqpiw3fjUN5BmaGxL3VmGhVbaf5MH0gODZX1WQdj
RqCsMh+ep+HT2/eqkJZIrGKxOsE3Q2LYLQK8hMRrQb6BNaupfHe9fsZtM3LiGSWi
j/ws80owpUHmRvycCe7n1ojpfWnQftoaSnxsn3bZKvfVFG1D6i3wIHSigqrNWC/9
jmyNN9VxxnEKc7TfaB5x0uc+5TCGloAi1k+YvjrH9QprmHxNZzLfiJsoZR/By/GS
/yh9l23zI96mCuL+0qs5eSA2fWz+d4cMATK9SycLvknZBCSjosr1lE/9VduYR1Tp
SMOW+6r8RrzUt7X2tkSlDpLchEAzlAX37dAT3OSCYymnNIlGzFK9duB4y0yjqmsX
gtIBnMuMon4FigdUB2ZS2W9hT37bdlfcieMDsYkSbSDYKuqlMTIsFC9z7FCIiQkO
Gtb4Mf/hiKNsjnDBj3iAbL4unVIZ4dqVetIbBYKGADChum3vdvVL6qviI+5qJwWZ
kxg2Ig+A9kogk9muC7JNyLeP0htMTiFum3bRXRsgx/r0sRO/sNYNWoanUjEN95lb
6o8ej1TsgcWJE34MZ/j0/MtwPMREtpyqJuX/K0vQmfNYkAs9GAe7TlGC0SP+uACN
eESAhGys+vHv1LoYuoN7P3iWTHi1XOvW77TwkOTnPI+E9TAHol6TElup4jnuR6Mn
h7ftgXFEQUK8UxqxtxsfkhfyBcG7SoqGczfmd+QzuJM7NqYgxibMySKbMfM73h5/
p7747HS01bbkk1b0s0m0tV8SQQk9l9g+UV0K3z+7jgQbErUUo8XvWrag2UhIeiEb
GmqtpWZvhOXO+sWPSfwsrCB7fjxKb3M3iU1VUHLo0LMp4ZrJ4xv8qu49TGqAdnJB
dV7GI0NEmcsVjdz1Indct6wxe56UD1DxaSDiE8dvpogTrddaHv5I1TmKFjhyAryO
wrHnII7TY9M4MNoEmaXBbB2cwFIxPNgv7iiCAC7uD8ohPpNw1Gd1Zi23hBWFfgEw
Xi+l7vZyYCh51QmLr+ACrAVS6avLFASKkgOq4+QYaJq5i6QEfw1bGct8Vo1Fwi3t
wc0WUNi6dJKNbbwqPAlvT07G+jmOVO3VMZGNsPQXARyYGcAJfO23Md7dJqJPGhPp
KMjGHAfdZzg17zCDdzWu1L+FwF5jbGg/Mq6IN4mrY+a+KCTjMjHHALWQs2LfO5g0
fDM1kvpMB+/4IDa6FU/yj6L1ccv1ARbSCScEYPk3xY51NriZFsoJVB86FIDjNE7+
NB4Nf+NbwyQkX0QCpeFfqokJsREfMq//yj4RUFTabWmwoEznfewUcV9fu9skzDUH
1gN9ZtuAKFGNPOUHsj0/+mynWSZ5rXqhEZCpfXOKpgYL6pEfp+yOUNGBCVfYvqL5
xy+fzx/fvch1302aE+XfyhmG/Ak4yeRGta61+oeCS7srAU00EECslkVZYWsxk2bk
njrs7lz5dcExvZLcSWa9PkLL+7iam1Lmtdb0ioq8z6OczLvEKUDEm/GfvbMpLb47
Xi2Bkms4NAGjqTVMCyKDXrAy1zGGz7nqE7K5nN94qeO5/2BZcWQ1LGnYFY/zgoZp
VPGzMKT7B7IyzFl1ML3aJYp0GVGmqIdyFrkd/9CqPtdmrA8KOqGJUZN4lE+6TWLS
AN3IGzf1BlRUjyON1kIH/ZxA7bHGfyXztKqPejZnETHnscTBE+WoS+54juNyVp/b
vbqqGOHekIhWdpTX2kFozXFYD/5GeJ0w1LuveuSqx0Bvl74KP6RSy2QVhc20zy+R
673yLoWBXvXirqXV6X94dGUX7Fu16X1W8z3slASXvuz+gyvGejEyVzz9npNVJcEz
SXX6QInpKurXHnhN6RedEr3c44lf4BFeFs1yomK5Dsf4SZyIburFBxzmLnPCSPDv
jtjVrqzZDPJHig0TUpbqbRPAh+Q4INcuoxVFyfIvOD4PZC/X1zZtVRNDDAZkQnoT
myyLyCKKPQlYYCJs/JA52Mzzf0HUBQGUoxF0lEGas/PikMnNbIxunXK/YG4TunCe
00CcB7b6OzdwAPfAccqwNvv+wgGR0WAIM4ys3J2BRIiulM61wOcmhjbAKj6r9ya3
txIDeToxmjUOZr78PtuK1OniP5doK+ZkNi8i2U48NmId1h1ZOGFVKQqWpCRvTL6u
gXZDWTV7gtL2OZpgI6I0E2HBzCMCRCIhJN0E63IwoflkgI0rIXXzQ9b++ObS0xYu
cVKSU1+OwjykA9Pe/qIrqI6mghQeZDQUyvOLxAFwrMnJVRbpWIUWPzpeCrxQY4BN
5sLxpXhI28kzHWF2LFHP2cXN0Hjo1CYuf0Wgg8YtP9cXa3m2pbaJ5kF0XTzoWgjq
b2cSjXc/hc+vMgUhyG6uBLCAEmv48+xAXO4GEcsNJDiDVVr+h8ib4ZHjlEcPW50x
2J7LQfsfxr/QI/si/qvTbfPC6ZnLrIDcfB3vDEU5ITftgTQIFRGvDJyRTgQW/1A6
48nsaY35rizmeiCEgRkMaHOZE71eXFwaPjyk44h1ddbFFL2EvU+lw8b4VAMP0jrw
36R/CYwd3WkE258RZwq8Lk0lLpRaIqwyPQ7vYdN2XOnyqJZS4a7+w6R47w9NEFGl
44mMjtRQLPmK5F0AFzjISxkic7HaapwV3ILKl45OA0U4py+H23YWzg0jWyrP27Uo
NZpT8oqrwcOdWJprp9hc9ki5h3xqRvtJKkuOTSGkXfpRr4sAcs9jNVJH8KM2OMmI
0ss2fmfreDDXsjJ89WJ/a+HVXeQTu8MnS5jw1HEorhgKA19vAe0RBkFqsV2lMEhd
SRLRrHFWGiKSjf3BQ6PsDzaq1fbwW5K2xOaQgclzatlc43mT4Cxv9hkZztsByiLg
7AbaW5BHinzu5ZPZfofnAHRxw4DxZwT4iRWbJH71sX6P1EVzQdezfLt8cK51lEyB
IMOWTqqUXGEP3kLBmclErgxaemPCAg3XIa0lgo5VRd44Ki8nh9DZfLVpZ5I6Xzar
K0Q0BwMN/hSkcuUUuIpSYEYbg8qeBTn+Yhva3EwngAzFJ70GwlavrEA6QDlaUBcW
jFtrT5v8VVQlSNfh/uSwuBkfPGGvXwKQzANjQlS+pjYs1/0yS76JAkr+r9nUdSIn
OkXT3d4UxG1OPIzAnQrTyB2KntwlEHOH3Uqet53pgxFqsCyQSpIzdvgCY3WxTHTj
qars199VMzvgzziin8diw7Go+6tSVx+eR7ql5xh5XkVY3KT6KdNJUoY2BD5LUd1D
rfoIVAabp/cMKJTyacv3ipBcnqAeRdGDdGHxbS8hZNykdrayURT11Wlssa7ffPBV
YfJdIbOGGUo0OTLDPZjnb+S7aqwCDXaDJzEQB21v6fYzQXILwENotwBZY95xX1s8
7ztgLHmfxKriepyhTrIJYBfCIiFyW70JgZC/zji6IQD8BRGAQL1r3yD7ARpHdOVT
i5VNZHUFc55w/79bFRGxFvYAwO8VlSAOA7aSPuEvD25ArThQYjvSOuBRYE6jqToY
+mDVzt0ZFglCkqv+RGIAdNU1mg49nwyWriwKil1JCjZBzP6HN2q765tYFfVqT5gQ
glwMtAqBScRUIbStsIDrDWUSQld1Da3ndcfqzSw7t43s+4c2TKn647V+1z7pyM/x
y8RGlojGoLhyq/XKS2WHZGkCq2lBXBrWZawfusH8Apc2DBay/hvQP2nwtICgV8LQ
pScuWiA8TxmgjRzKgEXWvqecit7U8mEbmHhsA/I9yi+iGEceXYV7mU2oqd8EQgV6
kOe4IhOPQT29Pp2jUE/nmkaI2IlzcOTnS3cgPVBwTBXpgZXQVcB4G6oT4sUjh+B6
bRvw3tKzryCYT7gSPhI7hjioS1Pka+gfSsvALx0ONESeaKfpvCT69+d7Ta0b3D15
Mw+EvpEr5Tk3L2XkPj3k44y9oJjgxEI9XocSYurhdMbOQmxvb4YOEhvNl9eVu2sn
rsX34R4RZ0gZc7pj/Q4KEAkHsi4550GOa4q9q1dL2cc6ZSM5Tu5GibaECKJiZVlW
KYAr4bhf1lo1t8gFZOEgg3wpJllHm1ebemkfapMBZPq/AEqUOrDg6zt1aCBuyyXq
jjg9hIAx/Et4u6qwzEEXRDoG3waITuwb9Aj9O6F1DzAUeYmVwAAyagS4ATECJYKF
PpsTGC/shZTEyP8IuWbQoYJlGzbCZJEzjTQrZ+w2/0dUFWLC9cXHcs269QYy5xNB
1srCM+ByyvWScdTHu8TLAgYs3jI32opgqDo+9qox7OoUmWIP8KfSTPJQquOMhxk0
FG4L8V7IHzT3/UTRddVtjrIBLM2KkuikwEzQ1BzWOYDK+HEKEaiDl/F7TGi44vtR
GmednrAUZQDi7tztwAbp/m19t71SYrkDpT9bJCzUyV9K0YmhpCUb/yaGwJjt0XIr
QIl4M6VubUj86VcitKC7bFbP2Rg+sicvkSP/ELhkask2xY4J+qR456wKbUF5kEK4
503oEaY/FT2mXYTZ+x479rV1lLWry5XJc6C/vyO8OS0xo5kvidvy3tpuj15tjjpI
0N59TuDGUIqJe76zBH2mjQrq4TCncanmF9Hr29ehDfBp8DbrlAs/17FTetZBa/xe
D5/BmIrKQQyEDhBauD4bnfybpOwRPtCYNgaOPQikgBKUUb4G+pIIYYc14G0HnXR3
SqpIQdYXu4F3MaO8+E1POHmPVYIeM2jremsicjfNA1OZLO+qNRg3SikWM0bXn+C3
tGkIyVxc1++IUVm6lPSms7+eEeMUn8Q7be/IJhYj0ykGiqehuYw2VDA789Znf1Sk
4lvCQIOHUopH+fI9ppQvYm1fDHDhu1GSUeqr9E85r1bxtJ6D8TOCCls6/fEEg2nR
cmEoXa12lVR1/PFpvweKgvCMoS6+5WI5Sfd36kqYamiqU01ArAEk3/hN48L9BiVh
MpiYTyQFWpaPMOgg8rzprmkgt1z7urmgyZJLyLkNpFWmOLaLoD64uNfEB1Vnumfa
+TOiDrlbU1vBGkUqZmpZhPOZ1UtSZ5oPwJKJzwzC2RuhIx96Fd/qZtxwpPTeAHD0
/gxMvlrNI9slSkQ2D7LKg9GGURu9EaYHFY670Sqisbogib6YBGOS5I7PfOlHWPc/
mKkILrK0HHuimquZd9zN9yeSHR82JU+IXTmk+4tsM9uoFrk2LIK0OZ9sujCZcvh7
zDAAY5Q65lTJyMTikLC1jIZPExgw7sxd0m1ATLfjgPBaSTCTQKFSAn4X6yLn/1Qk
kK1AupxH7+3M+a66LMUnFYu2q30TrpCUUEVJjxzHipqxW3JveWfa89q51Q7lqQWA
U1LGAksEvoExuklIRRTiYPA6FvIpuaABrO3a/6/rtghmZHQeMexssaBJQL3Z4xnS
yeD636F9+b5vN6HR7Wz9jGdI537ozw22IZSXG88uVljVS7/7hazXpq6ubSn4riQb
zEN1bWv6i6p5dxjpU5Nje0Too9X3wfapM9SgztI/Pt6upCxDhBEm1P1dkLtSpYTU
cJdzvuGwXGkyvDImk+kmbwc6g9TtcGst/4K9BtmmVvb7/WDX0zWoTce/4cH885RX
F5ryXTB5CHRAmCavHRr3Jsd3APS0+CwBgVK75zYMEWxt9cpwlsNfoIjBgDJr0GNA
NsK3ZWGDyASz31U3x1RuO5C6s1GIi04uteK0xe1uFh1iJZHVNyKC9E2vrc9w/8uI
/WzTJHfYnSfa/n4amZ+vtgk/oGO++oxSAAGw65sPKyf70ImuozCza+cBiyEJqKA4
WPtgIFSmZqxZpLvR998Q2Mf43lzPdErPSpWYtB8Rw4a8OubpKMoXwbIJTrTab0ga
ruTtzLnPwdSuyaoYTsIEw8kDnruF4OkpCw+fos0DvYIaKrMvjC/fHJGDbroE7+Xf
Zp7KtdAJ4lr8CWp1BqqPwNZy3RPDziDxxzeIkMjsznviq2PRIlKqiS8MWamukVii
zw83VXGKDWLwjfEIIcVpn3RbJkhRa+9nedvN+hsHF3TOqbqXLN4EkPkO/+Nn0f+1
LpmPYENZjEZMyTsppZhs/nkKVg0PeijPnoIO6beeUP35/BwUoPOdC+zHMObQ6gBn
KnmQvZlU8reryrJS0aZWzEpf/GGFFcD5FK5gy+xpGShemjj2IrW4Fu7uzmLweaKX
SIAEC9HhBeoQ3M+LeGewBygLPhVm2sss/9Q5uzkW9GPSmq+Ng+PwuoZTHx7fx9tl
/+QaDO9DciMjG3HLy7njPSC+exazQcbKlJR9K+BU6hlAwmhGmBkhwwVxXB95OMEa
3HQv2BrqS26f+E320g2iVKzaQ3yuCbEGEFcPbvnR2Du4tgd7LZJhbSpAToSO3V7T
HOEmTWOTqg/L/rQkrIGDGCkVkvqM3A5bbIU8UDGBSXvUN4imctsLVuUT56bPn5gM
6bXFrM1K7syDvLcJnzOWgYMDtg85jLSv9Hc+qOPae5xrLnMV2suIRCgbCdGRbpNP
j5J92hgvNGkC8WvlayPj7GNArQHXI/e7u85QNzgALkABdyB2bVu3yHmlynu15CFE
7I1mMTG45SCiEhcdI1RmcOyv7NDwTVgqpGlbYEZOLddUTb0OU5O5S4O4iMTCiy0o
FSZpFcMMzExTlF8m7fhHAeNqm+6pFVvE3q8PxdfG34P5yZDcvqKmyScuUlC2twk6
8H5bL+jc6aolQvvieCv3MglISLSWMDO97mqyk2u/ufWXz4BjmDkBtiFU/9kXeiky
5kCwwawv1s8POz22/WxNauih8oysadOzxyuNrNhCl83a+aEKOIqfymLM0gYDbyB7
zcOhT+k6KTOBkYu02m4xLuCfuM8KLYHNQtUzszW9qCubLtGSQYBTEYTI46slDsmI
lDLc05fZO9GiubM5F//0Oc+kXnDWsq6UwlUQmpiMLjOU3y9LCcRn6wAPkVo8ZIh9
Y1c7KK4TZUi3S+aeT9F66BRMsUa3thOnfl0ouOBSqUBO7cZrVFRjMXevdTMg1NSC
DZV8hJZ9QHsxO36Ye4g/bUwhf60CaUKpTK1hQ/9JAJqOfQM8tvcK57y3/DO6BVHU
XMpWe7uvlh/JFWBxQ7F1hCRh5/C5c9ymWMwSOSlWihPjftm/FhVDwxDcrK/Mcbwe
J1CKsScSQr56YrAVV9KnyV85nnJL94fuKcq7kObtkbk3ZPQt8xfgH0E1H/L3qwed
uyBdUdJQZzEmuLYkYOzHBs+vIgK3r4lHd67hO7rSQ5twLr2Y9eSdHw//3LHkXbY3
cXtNOHzJGdJ3JPS/z358s6OU/JTu6wpRxTnfo8ZKi5Kfsieo48wgBLsSlEK5WZvs
7Nkcf9X3V1J1EZC8MhBq2vm2AXkS4qdH+cP97gecifa6nG005yxdi4vK90Kq6IAa
XxQPEcQ1GO6Z5oGBmtmgoq/DQ/XrIejFxgPK+RYRe5TP367fK74fGk7O6CFsZRjM
ykkVX9cKhrClNNqwV+pwslvB2YJW2Gr3Nx0e1zqeB9wf0+c0WPDwIuSTblNfNwCO
Vj98pQ9hqbu4NTtbIOtwYY5TI0xGe+gvqoPbZs2S0742G2u5uXv9We4uSN9wlb2S
GVyGxjH2WapEXZOtTtNL1B3VADBhgj+KB0tFN+hp5ZXm3G7B9DbeM9GlxDYDi9A5
sZvoDGTTfKUgpTb68O9RqCxw+ZnpIikhIEfWNth+fE8S+/RfNmfOiOonfCljENg4
d37XD4zhGBldv7J0Z9Ojb6Ll5zx4S5cVNLQ4xvBed4rqgfPYxBLOlS0e+JYeRWgz
PPvgB1PIlf+SLKdJeVWV+bgEVGO4bBVbleSDKklFD+mx1KSU5zGHPMZCihF20qeC
ZHBAW44yFl4R/5444mofnlX29kqycLVPVfzl2i3xn7VtKLRabWkuEqejrtQktuTz
8X5LBHErjN+D+ZVi9sWKQNNkxQWw6XrO7lc4BAUOQxO/CDJPqau6yL4HX6sansvr
JbDSLnD53+H2PQAdX2jdKZnMTjE6I/XttwWzHYPbOE2xUevaU2rGFAGkWbGUs7ZW
bJ97daCCK0N7zQLNpjhsYdeS8SWedPez8nyVBxLjnB3wWy40hCsQZYYq2/90s+eX
tFMr3hcaEgnh2v5r6ht4tuWZgpJH3Q0GXuuaehjzobnW9fikrBsX4/Pb69AT156W
APw+XWChAJXO+w1HL4h/EdpUou0qTpJiD9rrKomkcwtv9REFg7p6/l475uyRI/a3
ME4ZKWh1OglLQr5G3FP/GXyMSEqkmMc5WG/D/3//Sbfuqy7WRS3jdQoZbjCeewWJ
bo6+iGSGWeO61r7+QKu6CTDa8sd9a5RDy4laJvWCgD3xs76iGxlLlWin6OxlgKD/
SANIxi8aJdDW691j9w5hofBwUJKfRmfCp1Ao1onFKXXjUktBVjPoVmS/kiHX9iK4
/TF51cRwP0X0cFzr8YMX/PPRqjA1lt7GhJW0/mfAeqW0Hxet3hWXFSGnTF+QoArn
CbnXFxPWz/MT36JseUgrO8eZF/7QSLCl4EgMGDVStkzzP9dhY/bPvKk9Uxd2mGzm
ZJquWhaL1/0aIxNzCLFQskKb4/GanBhokdbBUJ/U9nXx6aOGEGUVe+25hsTXe5e+
rgGtGY7FtDGIRQRcAGlVOXtA+KT3VUp3Lw11gVkKaE7JGuysmKn4YRZCf1VvSn6Z
2qsiJwS7TiXKzbFEMOqmu/imvfSzRyJFhw/uIAbQxZpc3Cnom7dWZ3j8Yxm0vXK4
TwXTCJC2JWCC+famwYP8nU0Gz9e2fIkzx8ThLL4urW7aIQim9ahi2V6Hmt67cxvb
x1FyYCMvGJthsa15AG7nasNPlpnEjgvqw94LhFuQ/PBRzSMLcO5igXoZP4lsK8aB
RojzuFkvnwrINksJvHWhZjfjhSV46bwcxKp5bgyZllMkjS3lF6ZXS2qQfBJ5tDEw
ur6vevskKvOTGMb/Z3g7Y0Tqk91ltIV8geKOdODEBB8kEt31Ko/pHjxCdXUExeUL
3V0hy6Xs4IyhTuMzlvKhoHTFDCCc0M0PotFhelRDn5Ok/Dovq/WCFCKtsxH5u/63
ku6b1sTCBA8Uh3+wz+A0VgPjiIvGseg8JITf8g/xHbXvE0oS7Ayzi9pKaeyp2P2l
+gnOTcR2/EoMxqiZwI+laPnL/ANEb535V+qGkG6Hi8TiT9pkcEPh6aHotvHxVgNi
lOjvdhMbaPXuL8qB/d/zWWrb/bCM5LhB8mzSc2NB3QAsmF5gIsnx4ogXJmGkJyUL
5pckJM2DrImMekUtPA4BPmUbxwlMqqs7XcdN2C/MH3s4GHkYBTHbULXIK9oplySl
w1sgWEdE77iyMv5uDrpxSwmn6/QN2FblFTbZRJY9+XUO845beOl8OK3bkfurjmxy
VwPZUVSS1R7myJIdH6kq8MPpcACocqdcALwCJ3NKmHkdkomDxeeKZgojMD2/X+ig
MbvVxfQY4/WO3cXeD4aHQs5BnUjHlZri6XbHH3zTwJC1J0wEVvFK3blWm3ESJ86Y
SQz+4YvaGYk4IHRdyjBW/AU89fxg5QzkWfAzcd7q2rpFdI7FaGk939K8KEv4yIJ6
5tCYTw+Ydalzp6hBmrsCXqEPFjQ2cPP4O8uLA4dthPDJqpbL5hXFSSOY5xvfHilF
dVUrZvNg6TLeFYl6XIdvMnShy2AFbhh0vefItnxArXDD0hHAwe0NR08AhlL27zUh
dpg0q/sXJDS9lxrdpr8DpUJ2QhgjXOXAxMkmKsLvB13Q5M/nUOnAYDQpfcQcmlqh
eKKG9ytK5iFC20jd/vE4yj+hp/7lCGcVE/gi6/yVao//b/OrsJ0CoWMxC/s8tnbx
fUpVrrP0k0x12BL5PQxBy6srWABg6mUPWb16p8aL1LnyNyhzFcxdWAxPjBrWJf+a
j5CrL5ZncTMi53I9f4aaBjwDA7LDLriAeX6209RaoKOUW1n9z+Rt4yBGNc0/TBv3
HC/AiX2xNceazMl4JxXO2Y1ZNqKQ12ZAD/rBirz5Ho9P7Va/7usR7YfWZ4RzP8td
YjgZwQcgnr74NLq1XSWfWDZT7kHuY7fOY9V5ecR+PIfpvefu24Jgg5UArVySBPtx
mXu1qQp4B/RmxXYA/bpdfYDCl9+N7RrzYYSOj/eTpyJwFcxA+qdbKreVdedD22X1
Vr5uqEySlhPhv3m9rJcsO0CbOwFWZlg0RnSELiXO+NkSXyFLCn0YIk2iS2ocRyvT
4YnRKZWSqGoWBNU7DAUway1XOqDU1g+oEbIeWpig3gKxP8YJutCPGP+NK2FpC3Rm
ZfUYRfHVslI0SLEo4JXXesugrmM0F6eNUgfzoXa83JLIX+1ppZpeI5ahVvmc08cc
jAYXFuRJpj9oGPsuBAsEveCq212VOEgywIGVA9iH0ZemCHGbFag/ZfnZM6vOPtEA
rJrbcyMFppE42WCiTILA5MdIf3uMg5mk134xGV++2dlmTLwJVIaz648VsDUlnhAo
qFqgRBZnxVZhqlSpdIkxy2ZnS6+7NTH7gyVd7/fQhN4is8rcbtJ9/UJ+SZbBPC2G
NDZ1j9StqVswMypcKHQeARtWzRLwrogJwp1j5Ct3AWwLeEdN6RCqvG+JLFFJN0Tq
szC8dm9BulqJlisP5LsM2VFZSr0C5KT1uzi8Bhcbl+WKdHToN7q1xiAvmuAta1fk
+OJu9P3q6wUFd6lf6b+iDYRtjfvkig/T5xaoFtEUmNWDV7FfrWBgKAKTMDlcqHr7
ByEEoSTBpU76M/jGUE8HG2I6fef2WJDE7T07OqYbXQrALvoTc9mGmBG9CYrmrsDt
Bj5Lf0pVhKHMysWN6ASNoYBKLRhl2wYVyOl/04z02f4x890KuxqnC5QD7mIsnms6
yMoMC/djDdzjb+5QpZq59wkdGEMOhMjRlwqvNtMTQXYCACum8VQpOlbYt1PIum0t
bVShC5qgwwwqMjJjjSgu3p1c/xbVGScYI2G/nsVJyZuFSvk4g5N/B+3lz48FmadT
ES8AiGeMNpBfY8tCvI5U6s9kEtUqMqRrM9qy1Yu27YbUl91ULzwEqbYarxfhtQbC
fG89fbXUv/EK/j9zyMGKDmaOta3yGffHGIkEta+FHbISCFZP1eli57avXL4WLPjY
zyeZ21557X5IhPxOSgxW/5NG9UdC5AnyWPU61zEtygZmPW5AtM65Mf8JciqC7iUD
B3huG/0zVvr7uetvwsKihk3Mz7JsjVaTthsEfEUhDBIEnGaZW0XbELWnpKPOIHYf
39i7/lblDY/tdztK4PR4mTNiJIWF8o74Mu6qpUZeVaJUSm+OtvGBiyB/KJzzyswe
QZNA4KtdR3ZeCS7EwQO1IzF0lJvebZYFj6dqFu04/NNEb3do0RQypt7jJtZCHSe+
/oom6V6SnK2zzouHLqwSAuYfwoVqVwmUBmXVS5y1t4p6g+8+RWavEMq/UcuKePHB
Fdvr21z1Qb9vqF4vaWliCo4Q1Lxiy7gMvxOlOKY8bayqlnnwmbMQjBAMeYol6Q3H
p/OBWvUyPJjiviW0o5CrsiWJBxfzp3RrVgZFCMM1g0mZyTzT6ggPD6HKFg4x69Q5
fIny6ETg0CQwOfkqfd8mpQKYI98NY5hUay4+j69OSbtvrbdeC8lxZfzyC28px5mF
87XH/BdvFHA5ixV+XJtpWuCSkWl4WezjLoqcAhqtI2IfKIPHYvdZglDh+UgRwtE+
Ej+EpShEcLTzVqU2ZIhaQU+J6KZ2W5lZonQoneypxuo1MWgqjiYGi0aEcwFqPlkk
RnGUxYNCyN8sTXi0oQKqb9R6NAu3WdfwPOUJKdllmKF3VzlNEuMUrtUEwEu5G8qR
TQJOcfriKuBG/8HR9E3HaZGh7N5gzf83bQkdC55SbPgD5oH2bM6qaylnHblXf88q
mMDMHVvSDAhNxS53zLmLPj6lgjA3Mx1nMu1tT2RkmXnEX0wZRqDqDH0nqWfuLShu
kjEAYPwWTwrbFHodWUYia5vBr3pzYZW+xXnEyW2JiI3v3bu9bn3gnNu1vsXVgkkJ
haYTZDvmRVp5WKoQXREEALSGN4rK1GOMQUExdsm4JpwHgPwXMVy5FAQZ9sxnQ9+b
LqZ4iQdIMH1PMEd47Wg4eLGbIKAvhCRusohu8gCGoeYynWTT14Ts5vN35R+MRvx0
oc4yxcM7t/wNdWmfLzfAYV+GZoVpVEblG1F+yvEKkTiVQKXAYhLxdbFs0wjXhabH
zyfU0B7w1HUjvqQX2Dp1H6c8nNL+BPbRvO0KMvkJPoPStIGSOicYsliSQMzu8Vgl
J5RbIrxm3rEmrhzqA8X3cdOtLFEQfkV3uziOoi0DaZuFE6QpPdFcIYk1ujR27NjO
O1r8ZqsMYk1oXGg0bvSDezaNIHznCy8pk69oBtOrFIb/beTB2eepHdE/vCy+aImC
JUwHoch0Wk1v9XITJpAWj0EnKblrJgO2HzboYzAIzJgLia4rOmV/XXvoiBXoDv57
bZ+SMUPel3Nbth0WtUmwY2t6Ia2UKVwTTqutczUNuTsFrpztcMfK1TwcITTiuM/w
hy5urNdI9gep2fP5tVTpeRI3DIviPzJaE2sCu/IyS+1V6MEAY4uHzbY3DkRjFKgq
N4geIQepTGFn+HyME1gzDSkadTFKJ/nPCIVsIc+JMTaNI3VZp3KEiZ49x0JhPrpD
KgdwwRTE19n6RUSUONzax0gbxpS+tKu0RW5cR2noezjm1lSy6qb13QrCbnK0Fazw
2XavzS6Pf1bzPvVoARJub8frbBAM686+hSaIDCvVbACx71geeQztlysjKo9sIUKH
uwEDEBzAycrOYCOT//8xt9OUK/w4mfsK2MLrqREuqIEhkRLM5www9Gucwlp7ygnh
c7/TKPrXwmyK4T7clH9/Benw50dmAXU6eTNFAKRT/EbUGdlevuAvKHC3qKQfh3ER
JFJN7rw4+YMxFxaBIDkPm8Sz8kDmcWbUEepoXjuZCXx/ZFlB83op+KTVvknTNEeq
TMYbELZvkk3GeXSbuul23ThQJa3mUc5Zn0UQf7c/y8U6+LrVIwzShyXaD+xP905x
TTIlkiDkvv2YlC+NAAjBM7Hig+Hgly1zzck3FPqP5FOZzapxXnCOtCF1z48IRSwD
f62EGjWFJ7/sIYWpm6kYe7eVyRWkjy8uG8pcOw+0/mIC+w/WeusaF7B92JQmllg/
WoB/+MeWnD7AoiOoR6aPWHMcTUKz1BX2du4TTEIFxWb9OsR/Q2J0RHXUa+Hcql4p
eKP/NrKDbjCr24KfRdc3xbxuyPpwZXqSQDkl49EDZu9UYHNmDnKgZqF8oWbjWGsT
kSdUauV/mgUblBEcuRN2Ww/ENSS664+z8EimE+5mk5pvQgqoCg+4S367+FejrwaZ
g1qhEqjPAVNew5H2ulyqlXeJUl5To/baC81KyEC5P3uzER9+NvLtWW8Hkp+cWdD8
APgK00Di0GX7almOQQVzkbrn35gGPmeyvoJTgzg8NSAP3/qKLTDmD7S0x9fWLIuU
8q7HPS3o+3t5su3rUFE9K30sPNwU7bQxYnvh6WwAxREOrnAos5nr1tM+C5fT81uL
aLuO/IXX0wIoV7QIxG9yQU5tO+p9SPW/GjLKV249lRD1dcg3Oe+PeKwEmDWslbNC
2SjKVKJpTRYljAostkZpVfu107SzSbM2iYmZlYvTkBr0Y+0M3DtygCVlJiERucGd
EnNjhZGzrGrP+HfFHhqHELG4GkG+mw6PUXtVy65EcSSWwJ045c+2ONpzmby8CFLe
AHlSsawkFPvWFmGWFQKON6FpIDQSu/jgA9Vc8MYte4QzK6JD6+zG9ii3iZUmnWQD
yJh/HQOGnr1xE0zFiCAd5o221dlu1OgTlpg33YrcCNGHftHZFVRWKdeXs8aFsq62
7Bl+/3bbbdItvdqCEzJJSwSu4eGmjGyDR39+khZWJMmwdbyNMLrNfvM0qIcHo9XM
H8pZFcGUtfmrolMvaIGlqIQnKmV/jgE5ZiCR0HAPk/rg5jyx0xZ7i8Ji5UwIjTL/
9Xygg+8lu38rdFqst/zFSlLpS7VvUx/eFIyaLnl8NeECCjYiytaOETRpt68R2iS2
JLC5wep10CSWLkXQsmmw/YAq5S2jcMwkgeNAx+/PuXwxvVDqfRLxGuJr2iv3tlVo
8ElOF5lzVHxw/roNlMjHATtL1RIJpXOT/b62jV14TsZKaXM2ApsoVmi8huEiYnjM
IOO+K/1tlW3ao7DOvnat7SOSvWTaz37Pe4Q/Lq2FABQTp/4h+KKl9TA0IDAyO3nG
PnudC9IvgaGSmDikvY2i6kcynLyF9V5JSkOjvlQZcMWMuX+KpBKyt1bvihKvaTJa
L436EY2BEWObAqR1WOCMoDpKfJKHX56f6cEzHLcNMIfbxkanumsWRxcyePcVZX0n
pF3UjTnxLOY48bfTPcLOb8iwPPdz5feKTma17dNfC+pKLOVsqiZ5DikRBv0wsBH2
DTSLp66z8UivRQFUa82iGVziQ/I8t35eQl9MOG+iT+U45MVuebple5hzifpOFyAM
Z/NsBsksjnGC3RXXGJfBHYkXfAUnqVWjeNxbqVkRf7/W7rWDdj9+kgjLMdbkzczL
ZM6Y+NFjbZUKZsMKjFRg4DVkeD5sRebf8vgyVgkS9G9GhcBv53wuD6P7d6Y4u3vW
ruIGTPQp67yfCDFXM7LYV77DZoEZFscGS65+ymJRr8ZHuJT3C3ndvOas0/+sLTck
Ch0Ob2CTt+sCO4Xl9n6wF9qfZWWCRU0NdAjLGytF+Eck5VK8WzBU5HFUvgOiJAQz
nAm+mn1T/QFyv3YGwr87CwWcTcQzXc27Npjvqp1h8zf+ZUzozkddLZ8LSPV2IVwy
CLTQPk92UIw6X+IjW7IzBdprceIWnu/Y2FBWu1UdwSfVe7PpakXr4YqKUoHrUXM6
farcm5hqFHtKQqr0xO+/JmEmUrVITkG88UQ7Fe7wZcDmwBhY+VdmnFoNVjg2VZmo
YUuyuV3IkS5ZEHqxUJftDj4UHi3pzveC+q31iTiFKoEd3p1k3oQaawhLAbYXFj8E
Ug09Zw0Kbfpq9UpOCxp4TAcrNdPWlu8bZ+tzCnbumD4CrVlz+R9TuJU46qkbzGJF
WUKj7oet5mPsQNVCr5yR0cSDWMKX7l7bTlz+RoRZ3u1cwr3/JiFZc2MTXpkNRLPj
vOiTdYiGTneJMc7ugOUFOVLPp5kZhVtWzDu+NRLdjOIhfWFCcJvEE+fydb5wgIkU
/I+61Q1TQpkUKtD44L5lWFKriGEV6uLbGhd42yX3Wz8nGpQkXzeUtDRlEFUcR+BE
V9SMQ+zE7R27CVeX+V+jtBV567cGiGCVSmex+4aK1jMD4r14B7mvxso7dMpIdXBI
VlRGrWJLGskS1VfP4DY7c1VFDQossZViFlcka4CcjTxPNwpetDo6tNIe+ZIHAN+w
zC84tL+ZjBqfd23tTVXRFVfxd/cm0c2m+LL9X54bkRCm8wxVH65DRUH+eBFanM6s
O4AmpxUEYF+wL77PngjncqfV/uFAJzSHC2K5+wsvN6ZdIUGecCkc+QHvfDIvVhOW
zdXsxrQ2YIsxSO0DBJRx0emiIE1n2CfmeAzHSg9HENuei79itJS+tdcXTI4+iabz
sQsuyCnz+kAOtKdFoG3Zciw/puRP2hCtWqNE1PgwZ5S1nam7zv3GbjJcxpK2+gsg
hjgtrjwBsp8KaR5nBIQfiRC6x9Tf0msAlGMc4sM5r9fnHq4AJ02cnh9nr+5+NLJ8
3JGZroYXEH9K3gwJapQEoGKsXqsSx/jq3Tv436TpXctZUtaJRAfxjyXcehsafdHN
ewP1rspwRyczpnTA/je6wWH5xgbW9PwRxE5TTItSaSPkYK5VzL5UfS+F1IarMQqO
6arIyfWJhzsplQamZF9sylfzjjV5iomayNxvBz8Sb7t20VEEEbmUrDR9iEf4q+En
LDLXP4SR3GByAkJloOhcsJdkZmPpj2ox6vYbKAhiPTUShuIeIawmG2sYcZ6+Qy05
Zbwkxzxf/4+5BfunQ3LP539lSSdI6DhNwQ/N/Zgrp1yi+KwGHM2spC3VCGC+3dPs
P+ULDCfXyzbYAx6zDFCU6khOxwHq2MFFVzYv/+nnzX6Phm3ZXC7a3mip3SzjXCZz
+c9vS8tXwNVMAwiHjZQdvP47fY7UV3J4lERW0WcXhMvQbQGGKAByOlAr8UOwTCgB
GCkRsYGTJlxC7pkhUOqew+chDhZ7H/ynVngU84eJWQz80U+t535wahM/FR5wEWI9
QRyMRSJffant3flyoNve1SfepVwgb7VxYNuw0gdYMdWjm1lAyCEzJdgWAHelFso2
Lg2MdbB3yzL6QyXeEAQs+IxJYw48FrJYdvLhpoXb+jik5Ml4DlzrMJD28lOVMHgU
aynUaSvk09ea2yJ+QQ8p1O5PfFVTxXYkjKRWB6nbvL+fPq3phP+7cgtPQ4cc3XpU
FEF9dq7ZxnWmMsAz5JFfBd94VwW0DJThGrEx3JmGKSL5ioZN9Fplk2zTlgy6Ax1E
O11/8B4ElyKw0RJBDS7rnRG1gP3Zz3bzEFW4ZoOFZh4GGw/jlhebZ3Qpf0zw+GGC
/WJjgPV/ZQKslFtBLrxUK/6/DgzSjc41KLy9zLTHIaw4CokATOwUg8Sb0QNEjNYy
NWhV85/XPTyKr4HerZTQgn86I5B01hIyJrn8TguOJwpTWNcfaojzYN4w2PFQ4tho
YT128yD7bO3LcKnN9gpdMM/BQBly7hoC7BXpC/XDL27Z8CjFX1dBGlWcL1hI1xqo
H8fp1xsKqHSTfI70UZvT3GHQ0GRNm7erifVU97rZ5A6yxhEYFXiHqX58kl7NyK4o
FFXs8m0MxJ1hwMwu0bQbaepn+ETgTxE3WhmldYUKFPyBZGOU+xm69NE7ADX6UMNc
2lkJ7xYLd7ZKZugXWUTgSxCBYdvnmN9Sg42/u1UNaZz2mFVEkwcS15T9HQiwgg9u
AUEVB8g5suTvcpGx8Zwu0Kp4Gih19wWmKeX5G25ZHO8egwekgyepsz4LOmlR/epC
ytofQa8PC4ZmC6ZGO7ifesVCOJXqDyyd1HuwXfjVXyFC18oTeETBJO5FYlpBB1s3
H1k40w/j9PHkMbBNpM1eUz59pSSjl65dp+1yKMHnHBdMB8f8MLZCkdZ8TvmAomCu
p49VnUrdWow5dr/0pmu4Lhmqf0Z2aH7Ma7m+IGxQVJ3Xzgzdzp/TfVDc3674HPUV
pM/IRR6MnZM0V+qB7KgkDQ0aClpc0nf1Ppr2jhyAZmlp/og0YSachK9jycm4Zwvi
QjV/eBzyWLpiRs2BadKAy4AoS0NJ1gy7RCV5AU3BddDmNr+mQqlZjSVB7OOFE7EC
JJDYCIfTVZS5F06iL9yeXhAL6rYn7FZ4MC1akny0pE5bIkImOGIKPBNadi5+66ar
MxSHLvyZ15fHL2y/ln8wbhQ9ep45z0jRbTgCcVhpqyyjtSr0dYu+WgNveheLH/Hk
inYcvguGsIiWY1D8/g+VNpLGQbhdxYC/4nS3JcQzvhT0mwQLUdADP07NLK+PLSUn
oPprROIiL2F8ZZGcyjX8tieLJwAM5HNAtGQ8PAr/9JfxBJUe3MnaLXLFb78STQD2
+6FqgQEvV4E6DPk/AxYZ986elJWmY3SXkH8NlsjeiZGVTWOAe1+RALeCHQvt0mdo
7qi1zyRvmNaF9UTWDmLaH2Q792qMbS/CY9Pw8dsNOVlGjfbhPOvAZYNPxwuYnIAv
kJtUoCy4N/9kjHfhp4fYcfHLo2Vl5lZxW6cOEMWiWHQgcVbB4pJQz8+DIDh7CWBO
fZ9dSURJ1ZxP/meqpJVqAnVRReOgdaWs/NR6CTA8cmNWCD4JKBYIIlBB0FuIY6hc
hU2M1k9+TpoefjvVKoskDafJE9Qvdy/sZMBZVD84I1b7bzRtVahuOdo+DOEkE0TF
H2EXAFHOX0EA7q2K4MPacq9vPWguIKP9aREdVpEuwNfVqlgccIYP0LZ6iSnl8M3E
PMTVryDmPWn0smZRzQjANbG8WqlsmXQUYIOHFNTUdoOguSLzMjVLFJfZVDYcQZ+i
ED+gxqH4GghF12s5ePwHL410GsfAumys9jg/wGtMp7V1utbEVrYmG2qEH5AV4dNX
oTIrZavFF6pFgxwFljtaIoA6AhBFZ/mtk94YjqCP+ph6wqjkrLupkaIMYrg1Otw0
fe/xBF5qjltZsKgtI72KK+f7TeVT6DEGvoBAWkK10bJkKr74KsG1eKVds7Ebf+UF
9x8xT8/ZlvqDxaN9+u0aIUNPAhIJXuBM+S1VAHT0tJrCHaiu0pK8M+MMwJ/f65G8
+3P2BJrVbDIQE5mkKuUqSTS6QycWlzE8q+hu0FHOFL08o0vnK/MupEvqGUFlIMb0
Gc6IhnbmpO4Sz3HpjJJk4y2H+lmzrnJtcT9AxMb3DuXVC/wqbA3bz++7nD9aes+u
WF30hKTNnAQybxjkF+ZJ4ZYxPotKoGx8No1rHYJ4G/UaEpclvERmeRjXJRqW8JWu
7cHC6+45yKxk1v8cRUfo9H5WbMBRD9Wskc5tw+i50f8idEOzSMTuP5hJlI1ZQ+B9
WLM9Oc761LZJcVVrRbHn9jkwmN8R8Kds9h5pyWrfnk/hjJp88ylNBkGXUjcReHLr
Cfg/ZqRuMf+FF1NYkrCy/s6bVaPyZ/BIDAeLiILJ0kqblgSwgEbCq9oRHK1snCMA
6m23CMxgcyEYrhwT45yoSjJgreXzbXfcricLn0Au2cUCck2HkHQPcdPy8wHg1zIJ
eenY+TTNVIp33mAHFJfMNz8EQ4lCW1F8iJAd/fRYhchiC3gpo0zn7QLR3DFtV42W
MpBKhqGkLskh+R/mQuoCOR7LDn9iFcd/qiwY75y6VwG68oOQKbDQ0NSLcF4ZnJjY
1ZIA8X8X2j30ZKVAwiccpy9w++ZjCvsp4SsqNnoftQfEv1SeJwwE3e4wOmKSKv4B
h/SkihY1vJDBHp5lAqFdeQSq0wf0RtTHvsSXt3IVH/DAvzQsst770HdzSky/zHnr
S6Ftk1H5TYRQESUgFW/Hr0lqa3TKKh6DKei3pbvUuCcSCj8Qe7dIbNVvIBglqrXg
ICNLA8iK5T9d11rulZqNMApe+JO0r9vi2ElKQAN9h9pETqqpRZzKFpQoQ+q03gox
O7GKbKASNsIg07DaoCOmLWpJ+bKnwmI03pytPJCjmEidxYakpSFE297p1c6TABaf
H5DYAhMWaYOZ7m7lP+Hw1gZsffSVuHTZw/gLOwBSxMiemxV007NdBtmy3yqg0c2P
mXjTfNi+hsYUP8T7uFNhgYQW8asnFXaCzVlmROTmWwFuGK7g9O71fbZhCoY6tkim
2TKsV0rmNZakW0zMIK4aTDJq0O+53i0LgojK5yALsqyepzYNE3JOmwjKSk76tiKG
1qiUYbMu418xe35qkKSANWil6em9saFe4QiUJO+/orXAvNy3w06X0ujQsWOHIurN
KFpKac9igm533qPwviYoZW5k+xHb2V2X8uJF9CaJjrL/NPBuhrQUGM69nC/sOWmH
SAGWA0PEZTMXFxlzvXulPon2xmMhsEJEgmvuL6oBdHFZ8Q44i8ZAO5xM9078PkNi
UsU+9+Txx2pjGTp34wcQS0rHFPAHR4wXz30W7oOgyJeYEttcgSq6bI1Rj/2gPomL
aG67M/eDhVbPcBBTg0t8Gs052CT3N7kspSP2/WX/aJdFP3rPHa3lpf5KB6BSRegX
p/Tw3xkbPoQT3xuSK0U+HDIxPPicSwDjYiHB/4WyLLcaKnDnl6bBu2RTuxOqN+mH
dHaAysdR+gUirT0Y7cmZ69brJqJtlkFa2x8FceHNa1qH/kSghLTkw64fwYxzfKMf
bgTG5DndNXKM4sXje3zUbO7xpDOYG2NGz6mwrjUcHNTHwlJ2OV8j/os3Y6DS5HY9
bbVs9EfjRt58u7iucAHITtYhpqDzbUrFzSfCqRWT/ImDZeBlEdDQDpW7zycYMV3D
Ku52BrWka1ROm3Bz/aMXLs4kcmKj03lFzTfyE8bGBxrdSG8lgUB19k3ncrkOz/SN
zO9aVuxplpwOLjBCtNgg63cwWzNomfgcnoru0roShC6fihIhBAaEl5p561QceqyC
EVF7H+Tir7/S+Ua2ZiZK0dOIBKsiKGUA7f7PUeOJbQf4KHvKHOGrFiWAGQutZ8hW
zAiNeRmNbqj4+XuuoQWo7hbdFH8ntV4YnVYFlqRVBwfyP/7GELUZfcngaOziRGyN
jT/Ly5GV71c2T9H0zzQrNrxcaEtECVV0oZrqWDTEWRCUxT99O0ev/6z/LMWOcJSU
69G5CaJS75dsKsKmn7HTHCt++Tw8t/l8c+6H1mSF2jTbgjhnjWgTPZTHVw+h3hhP
WojPe2Ks5ais1+OsBZ8fm6yiqBOTcUGzuTMZjmXWNJms1LgY6GHL5uuDPc96f4LB
rD6/xYHhw9/KxKy6j/QLepmpoi+pXw74jUAlkchjFFz1hodOvF+FVXeQO7w+85LU
sEbn0H4t5nl5pC2Bj/8LsHSG4D56w9/kCltPT92pwjK1p7QTHgx/BHrf/vtZ7Ve2
3dqnCdh+budotShuazDBDPYxHPFBwRq+zyrRMpAqrPManWRuD+/hz64vRzUpqqo5
8XoP5x/+8eZimbne0GTBO1TmZhL0zXlT1luRSzxdwTcll/+5oYhh8+73xv8aZnxH
RKXpJr5rZL65Tbe6goDorUhzO53dWtBfKxaOgw9axnGlETD9z570CUpIIiWKE+qr
N7sNTzLNoPdUCyKS8T4OjTssKr57p0+rsrdZLlMy72CWDbLRPbVaASHNR0zEGCTk
BELIzR7YQIgfQ9Soayn4uunHB6zf6LeKS+qWB2tn+oVsi6zvtqGFbya5FL2ixvqP
xuqwuY7WXwK5BOklyT3eZFOH/R3Ylhd97CxhddjP187vEfnl8wsO/1aldSHEs9pm
u7FDKWjL41TndXXCjcXC+YNMmn0HpTMxf2T5McS4GcquL44wgNwhwSMulIe46Phy
83+I52rNcBy+iETOwfT9tykTZBEjNRfFdR9FTcwd4y6zFVm/hqUVI0eQLBSzRbz8
0XQsZt6UwAr2/Yqzmokxku198LmTr9/WBYyBLGR8+8KqVI2+zyx1VXgOtEBFCulY
yYfoL0nqDIRxMiqb2L2RPQQTpGpEdlRUDp0ZT14qQ1q8o4LviViuVYVCMa/c88rS
og8uB5g3VXrvQY7L+Vb2L1CFz2G95ikFKvtuWeA/AdYUqbFHxFFIPjLva8H4Sfn/
Nvp5664jWtsOsz9B66e04Zg/LAFc/YKJXh8YWSe8E8hh34Cbyifc4CSHeas8lZgm
B9xNWSXNFw/YpsTcAa+LMYHusulqK7ulmmznisor4pzPVAJHHXgEA6KL3ph6hxva
Q08F5mQoGwwo/UBHPY3LhHNGOUxu02zY9tjiiBtNRxOaPXhRUe11IKARCGn+i7Rb
Dp53vk5dTBOFn1aqIOekQhlgWkPDc+pelSy8wbPOSkoOOUQpwlU6+JzpyjrT8LBM
1ouvREsao7n2KJ2lI2A5uvfUoGS+jcV4Zpp/i/9S7y2TFxuF+VrfhmVuWSt57t8S
m1SS4c+j05sfYj4wMJJtzOL5RWy01r52+SsWVG/OW64UvJWhsYzCZsGmb2YxpKTv
O9nVBFfpKX3QWC0f/9PE+3AfnQhRiDvy8/4cjRdstwm0xvSkTDowQMxAJvXhf1bu
biK/qMhiuGT2LkN/wbfwVMEn7YnDTnD4dCad+8rOGFjUv6eF3IXoZSTdQc2mo6g2
ZYiQMDFNaq6OyXalpntTaLob4jX8TOLUKZOaVsMGe6CwCOiZCd73V8sIfnga7rW7
TBXItvUHmBnVnkKmSJ3CcUl+NAgI6nODrepTP6d96UEozRDRY07U3G6JErdBXtIf
n+eg2Y8/QZG1UNIcJqMeHdDRRSMnSLj1787/JBjLhhVXzp3Heq5gnBNdPMqORSMh
/z15WhF7y/b9kmTV4Js+pB0qsRtD18jsM1Q4NxnGmSvmSqKU6UtGfSSBx/ihf5Ro
3WTqNwvU09nSWO2NfpQQjS70l08zEjowsovBtTOYD+MPWui7ErnAecPCXoyO5A1z
lwJyi6d0MFbJXUer6E699ft5PIfKMUphQfi7t6xTFwDSLmImFcHEeGk896XU5V0s
LV0AClaJKyc0tzj9b3YXTJVA1+SvI/SpfejQOAwHyvmfDnB6M1fCeRPrUBL+sXAD
Qe0FXiKhUbtCkZ79YdzqkgHJ6sQ3gUEk8QhUyMUEG0dr693XZxIgabipAe49PWmg
h7qqWwwkffA9LKT42uXnG7cWdDoNo9MdWJEwyJeMmx+YxK3BGBrhnRcpkC6KoH1W
Uf01nl1/G+V1fHphiDQcfwz11G99tywNocmbQwrTS5gB6d+lMjpUhwgL0utsNEKD
Lqi2wGa5zMFK3hCvTn7E/XrFi9fyfrXddY6SRaPgNvE7vQ73cxWSva7klnRoH/jO
bXIFKy7IPcKEIA9yMoLBckiax4jUs/Fm0z3o/pjNxTMRBojZho4suo02gX8njISP
r8DAWpbcFTMkw+fPr5bbDWuQPePeHRmc+mKfoXlouI13hT4t4xOAIInzAQiwok45
rPGfXoskalpY0wK/5xCDjkulEB383jN8V16xifyVRU5YTRsKWy+m80u8KJDtkfLE
GMSvDM9kdJaxKBmzQSUQ5LSBkOs94Ds8ZlKEWK5RuMoE12FSinecIAnowYSaTAKc
aUsmqGlyOgRSq4sTFCmFmuhVzhgnFcTUO7DyI3CYxfen1QBYu/Uck076GQlMwdKJ
qN+qCfI5rx9uF1qymMND3uPtVI9e+LROp3MrUBfMB5teGk2JnC+nuEDbYKvi9C7q
6Lz6lPbnIQTTrjyxXnHEUrSkoydtcu10rrHXa8x51E7H5Z1DSTJDZYz4SAoHevDA
xTbjrTxWTuYusU0BWyRObj3ABeVIrbuqoHo8r6/GiORgjBJmvdD7M5A+2AjC47tk
5iMFeSHuuJ3py8mowgAyJbpj4RtvqyazJzsv2SSedtVrGdMKwnhG66Lo5Eq5wmtU
MWVbFbPD1LUDBeNH1JXnGJ6iqdBPZtUWlLOMJXseBeWfoEuiu606DVqu5dMTCsOv
QyFPYqipJpcTTSjzTJ3RWkigBJXGELcBnXPHwthtDumNsq41MSf86B/EcYUMZpXf
93HgMp9QKftr6L+NS4iBkeWMLZ0ggc3S/O1Z/rVGo+U7ttk9kkoOMVo0csV/t+9v
AWPkZC33rGCIEO+iEjCcgLs3LRuCP5KPxTPTclglL84KkZ6dmADlsB89ZnX9Z7sT
snG+PQbBBEa7sKIIUl4fdnpTvu/ZzdHZuNQ6K1qhS6HGgxlOLQEAeFtbWZ6sJpoa
HjMckEH3++434XYwUVIv05Ghn19GbpgWcfM1fX0IpUNmK1SnIKDnglDngh6eNF4j
dOps0KISjg6Md9ZQ5ZgckBLPvcgxdZ4qoPHcvoGN6iguGMy9J+J8/sWbydmfuPmN
lLKhV9cpYvhrWRZ18XwdE2j8bJVGOc4fM3aQGzbIxTl2CX8WODsSt6E7IEaY4IpX
HgtF3szU6lx6gQR72jdEny+1oUC6okQ8/n45WMgtEfgRO1sdTIb86XTLUxKhmWku
qIAs1vOM93kHaqnwK8VmBIjAi5/HqiJe1xiqoMWMsnan6/9l71PpbTLIkZlhbMy9
eRdDh0ZsQHM30pWcieEL23VwtollrPbxKz64kW0/c94jfHErSujtziREaZFkSbsM
frwUKLxqECd1KhQumELKPvIVM/NqO4xMfEaab8959FBcIYfVvszwW6Qjw9n73J37
VZxbmz+Ds/LxnXraZ8Mkl1jer26AFC8GHoXpoxfALQOjBlM81x8SjyoG9ivJEfbx
is0PbVva5TgpMb23SnyxiC9gYI5sDrBrH+uXbZ4A9UYbGRw6NQA5YAHOWAsEbVcu
M4YLq1M1xIKeHsnWUFwtoIdBAwPFs6I19MP7OJsOoV3LdipCQIooer58DKQax6u/
W/ectMfVnKPmA81f6Ke88Jw4erx3/MYafgnKyJdtnpcZl5nWZS1oEE28KF9VOQSa
6mbdMWfFR2HvZ1HbfypFGk9B64uvSgqlXvFTTsPfvOgn/npNLkrArDin99t/kV4L
N7/nYNbXzspfAXW6NWjlgVjR6asRsTo+mA92LW8sG/0GljqAzILixOh0YnVIVqZF
G+n6pagGmQx1fqEVWaHdW6ShitXtACTVyTlsL5UpKOekApaP/hSJB5v0ICXQOcdW
KdAnN2/lFaIAxF5lR7pGe7MqikKHuTcosnBF0LnadU77Q88IDXKvifkWlMckdmji
GBGZIX6/vaTiVVglnK0zs8x9ZPl3u2sw852PkKVlAmg4kSvGGBegPEqRyNDdr7j/
9nA42tduCeQtAWipdp+3X/cT/alR4YeDXJfKDEaGQmF7ofKNCFIVXW0vep7Bo8l4
P02rAhAJaI2QuZGubHoBu/q70PLHKA4KK7Gg6jhbZX/9PR8Jmavv0YiR2t7+R+2e
1KFjsOdGq2Ca3N0L9xjoiXU/67PykniqF3ykx7M3KkwUUGImtXTjvvqZ4RPz3Jcw
jy+pKauBF16NI0Vk5aYFktgN2hghCjbHO9XOrP6bfyMEv8kMYll6gqx1qZrRZHgm
T0WM6o/SjNLrdlx8FtWmwqutmlGJneWUJZPVhgE9VfVc1J/qZ22D/poJGRErC3f4
QpGg/P1v7Pb4XyrswTqkRI9paEDtYOkRrrDf86EqudKKOqXIO30vb7CuJCUVBcri
8UhKU3sOpYSZ1EF/0IgxClfJ0OuEvve/4YsfGJdeRbpRVSs5ecp5M8Oeu0z6Zmui
raXvtYESkhJFL0Qu7n6poz98eqcxM+34i8GR/3EzOZ1aQU2CtYctCZYQvbf/ax2R
3lN/VsV56e1fK8TY4a+tmA880Nzci5J/XrB5PScVTw4jvoMco8KffjYZ9drRRkdR
ANsqkzqqOb1coBEqtgBOYmEbDcEEq5GcZVOa+REvqf5Ok/UdkrBIyQW4XHiRJE5c
qhRLwbWQo8z1lyXYAELl7qLJmgZA7wMF/Un6SQLXMcgqSE6dpRbbnd9RGyU0c7xS
0h4u5TkNI1KtgpFu2DL5QFnRunSWzwJtniU0gJ10ahEjN+SLZxAnHnmb5biybFbn
FzGodGd8k8KTtOv0AqXJoL9x4lMlbP6ZM2Evtcsqno+bMXH0A3cURaPFnEOtbKrF
7TmJe4A1qvK6Zrw6ouFUpU4GJ51GiH8yFT0FTftsQyn7mq8T7L61cRUXxa5YV7NU
g36gre6zAugOjI6fHTGohWpMJ/XcvWQ2EXfswgJtEAKhyuai3HCGXZXyblIXCyOy
VEqTrpt/cJjnjm1G3u8KFm+On0x9SrG4ayBLMmHqReZN9H6I6v7Wr8Uq6FDSw8MO
thP/4W0vy4z13eFhGvymkBRgPtR9qhASudkN7BxDsMAt15SEsMYeOYo8U63X5AJo
XVv+1hyEjJ4aLI6CwdvOcL9fmM6BuXNiqr4GugB+FBHvMGiuYX8anDg4yke8DK6I
7FATnzQoxgwoKnRB0ExWXjF0ED5V4t6jsDBBrSzkmEpyM+dVeET1xM1mLEPFvzVa
BuMCmYmY6K8d4rhbL09REdvPServMAeqUw+T766s8r6ehHO2PlFpTnKQQWjrlC0x
SoP6JbyPXGnYvmB27uhbDNGTeJQTnQrrteuAvpDw88JNQZIRGgqOERnLC7PYLzwu
cwjslAcCF7Iu+H7c0CfP0nERD1VAqttdAZm4iDPXOp/xzDbkfanpdly9KzRacdiu
BUTtlT16PzZkVXx2CXCsTa9fXtK5N7lBvY1qRfeu4Avw4LjLTqolm3ZQeNcM5XI5
FtbDDG2K4GdgC2hJ2hRhC818c1D7BlQnuY3IFnEYf0E292Q8EfxYA2hCZRqFa4Z/
qO5kN1JfNWcaHxtg4gEooVVMPjTn4ixQUvx+IVj/Gqt2O693vcjd8k9/P1C39+Lx
lXz4a/NSzEJvlNeZCuNRcwLrE3+3aHXVQd1n4qQyAg9pOOg3cuS0rLAUktpy3zNH
svUMJ2qWJD5jTfNM0LFNKXAYyze7wqEcVuiRG6UvDcx+HpBbVOBWVGlAV2Olu7v8
x0yQoBDXEiygyzTFoaPCNDEm+qRrcO/DvwiPBBPsrv9Imh8QE4KJGTceoPBJfQVX
BUf4BDbVuEnFQd1o577uWYBh2yEzVnHVTzFcYeTc3WnWtr4t49y2x+cFgp+K03/k
f0TI40trJDNFsKzHPs1bsX0yn++zM5c4aW7ETde+w4rwAMV7ZBMTIwMTq/hhO1zr
En8S+qslrDe/+HG2RuO56tj7A0yVEpU6isPqz2iPoRUdbhqX91TzNQLXjVI5pEgm
5m82I8Ce+9neTjocnUi3a+rA5dSyhk4A4gaAjj9xT3yrpmfCcaGox4MDvh8oiokh
ckG56hL+IbuedYdcqxM435nTiAp1bWmXV5vXz3cOAwle8YlXsfWmc8bq7xZMJfbY
WShIO+NCSdU/ggK7ZGH+Wq0GmsXZM56UrHNkEihRc+oyJQUqbAOn5HnHBDZdYVYD
2mpDFj7t7SnKZKzjJxO6eDOwbDIuPtPONdjHJDLpN7J5qGlp3DISCa76Wt26M3mV
yZJ6AkCXKHqPY6DiXIwAKuNx4Aa4YcVZfDV2SKAB19ayWtVFkjpCH18iGy/l8jP3
pm7fCg8KyZj0uFqv2so7sjQstRM/logliEu7XUPY0FLUW2QQD1zi7T8ybiF8l+0w
RXGpxneINci5ur6mo04r/y9AgqEbhVQTc3o40z8ghYCYiLX/+g/Y5kKYUjM//2Tz
tv4pVyuaL1ouoHZdypJvzxayS250d5GTmtOHWwsESECnUqhjQaqVo4JcsOrwcE4d
aIWRNMtWm6jKwe9neOOq1/HHIgM7BS2BCdL1MqXm3/pwOte29U9pVIsxl78jTxtR
FGipvNmx5P7ZcZMmsdKEYc2x8KAIuZ2ZX3bRRDoOD7TPW1pz9tI3Y44gn+xiY66r
O6so92mB5omhQqlis/YJ2Mawo2CE5BcGwPGwCBQ+yTLXz3nd0myniPJQfbWP6vdN
CXvbMOUa8wIbZkfSvs2bG3iUN/Y5ybWhUs6DCRF5CL5tBLSs/vvsnZAaUrwUu1l+
fttcep263EVlsnoKwz9knCzzQOscAHVVQ/6SeTk+YJqA/eXnwMNm208b4HKO2qry
ZpsTYbGOAK1+1C6PQBITENforZaWWw+2BOEgUDaadnAPhjt3iL4w+DFg1NMygCko
3qAmVZoLLdcsotau5CTMX0x59M7HVR4CNoYleN30hHu9/YClHc6kYnUhfyr0T+wa
kTRRpN8/b0lUnLyC5SN+dEax1jKmLtlCwr1YfOxI3NXgbVz4vB+OpyGDemCCq1JP
zmbVIyf+872ew5FbYH+fEfLrrgXATDoFjt5BmHPH49+C7lwoitxEwmJGFfdTotzQ
fwQZDt5vs1Ih1x342hnUPTqvLUNjiEwp1R82ovLEZm4KUZJgNPpFAIU6rzb4/3a1
FuS1ZO/VxFVSTF8omrzxB4CMZ5W+sba0eKe0XsdehkTteMNUokCxPXqo8sVB1E8u
ZG7pjmKTqs68pGQcll62lcGaS7mkOb/k5wuj2dR2U8+IhAznr4S5qXfbVVFp5xs0
gavbEAqBUcpLEhZnhYZbC/B8pMzOGUZbE8kMDfDFd/9MdbvZ3Up8ryA9g+b+CuwG
X8nTq2B5sty3l1ufN0bkd7X6Tak+kHM5FA9Q271Awq6SVLfs4miloNQ/vyvh5aIY
nMScCEYcHt6XxUYv735IWmQQi5/qei1aPSclyALY+97ARyrFAfWhZa3yN53xcYA/
VPGGStQ/haD5snpKD9dCMoY+2oLCbvN5Ced4FbrU218FZ9fI/zI6ZU+9I7pDNPS4
63wzwyQEohG9hAMXSuWCIWKv4JTolonvu4MTE2pcz9kHq1dDYjAaNAlZLbXBbrLs
woVId28HlhndjK8shRyf1tQqRg4KF+nylGS1RjyDBrolSawcQer2aIKWm6qEQjIc
3HVGftlOXG+eFAC4U//vU0NfTTwBDVTvZdHQunjjajDUcpb5pA7tTMFR/krgZLBL
kgZeqlie9l1NKbYIJ3NbGo3Smg4a2fMUZTxgxlZbOXxP3at50YKh8R2Ut3u6S2RR
ESuLk5N8SgCwEFARtDlwz+7KgYQZRtyVCZnj5T5UL5/rF0j8luw5Ec1srZRKHprr
ANrXsZO07dIS+iefWji8BAqM4H2B6HSImARmaanZYUZG903f/ie98YGOMuw0Mbp/
DaEZLIEhF6M91ryQBKs0FsbFdEhmTZHO18+JxSG8toeKGYR7sSSl71QfWDG/q3P/
SRSsEyV8KJeJBiDmlPvcEMWh0H9Srnq9TEzZ8cafEDaY2xFEBQNF3S1HGj0kxISQ
fCvJ6Q4pU9tyKMGRnCDi/gz4RFlP1hEpqeYY3GhOAvnZmfhD4TH8j1F8hGkWM1yY
o2w0Pf2YFiMOcCJ7mr1BdD11V2i5c+Nwho1lKoLM5n4Q1vbfuWkENLNCOumt1lpy
kt36CSczQPMOueiV0V9Is1j7lFAgUlga3UQbXoXIEqS6Pi7748uvheYIBcAvlHGx
PP9JXnoIumEejForSdiLZlhp2OSphf9tzvnrLuqxt9rPt+R4J3TyX8mOq1+PW/O0
XNLnyxn+YE7lYwiH07TINX35mUOXk+OXe8eUovLkyKinfvN3IZz5JnwCGf7pA882
7VMbtR6gG2Q7Oeat3k2ZOTKPeKmsK7+6PZAQ9qzo0OO1hGYvRZ78J51ffQ85T3hc
y4Q+GGsWwlfVbdswlet5+6kl0XmDSQ4Ahr7EvXyw4tkpTsLoIa4Zktd55ufpFX3/
wDCZK2Qq44sJoxRlaBxtcq2q+Lw/hrYVmFma3jjB5HYZap8Zjm+BR4zlmqUZdiXF
6UptC7Gdod5hEKeCRIQdJEtmbPovGfDH5Eh5tqjg2ZbOIqsU0azyltGYMWFjR6jq
xoZU0umcSFrKMcwxx2nSxsmp51gFEYACfoz5Fb5bQLdH5arM9sRAUjGsiSL4fYzc
5Ft99AgzvrpPdhhWsF+lLr3h78UOrqgir+DZLQCN8p/PtbmczPVPp1stMyRatnDI
RAZXd8Qoh3iKbaX8QD40koir6JIPQLPC5OnS32Zu2KQtEdU3wwBQGmZicHF7v+qs
vXQdksAFa7t4E3K/+5AAuX6/ggE13xGR90JhbQnOk0ioocWM8WKatqOOocdc09RF
kzB/e8ZigPsoISu2beUYABvVzPxj/+RqAJvAv2z3Ys6JXiLYCLwGDMjWu2i0Bs86
tebwGAltE6tS0dWiqLwEp7G9YvJs+4NjiGe+lqiGKG7Hod5lA5wmxPWIUBUo8C0S
VVvpaKxxM0RledUfWQyN5DKPQCG5tdYq/FO6Mbsb/OCEC3vrM/dO3guP2Y6D5rVX
h8O+3lXuH4cn7yOJFP6q7I+u1f4sW15YDIxVWqPnuBMUmXguVmJbhOfeQFlxHPnd
2tF5dZgCEJwk2INWnm2oeBmw82sAz3zdJ/P9dLQPYxXkDO/S6YB0s7vB3gyOUFuv
Ni+r+2OxsieKX1Dpr8RTDWw5d2pBTsAmcqBCGxf0pRfHrSJOSyE1mFcwUBFIY55r
LybYqZF1bRywPm/qozip0rdh8v5ujXrFwGGHLPzAC855laHrRB73y1+ttHyb6IHP
5TskPfYmL0nJHfrcqcTsUgb/S1tjT+HQ41eFldwYOWmVlGzhwmoMux1XAfVeuTmR
12aLq+Ju9A8S5YvIFpKr36iQOI4HGRSKnABCBy1rCsnHLhFd8X6HBIY1X0SOc2SP
048Os46upZTIJln+tcCdXPJmhuTCKauMEyJlMYCteJTpqKJdnR7/m5nBMSe2+bSR
Ehi8kkfubc0y4CigJMXkyf5auN+g6ISlbv8gR8v4t+QWQ+rg9Te8QwvF5XiNSLMQ
HUI9/4BlJ7qeocn2OHXE4Ss4zHMInrE7wLoYz6abzQbiDcawtF8fKwZG8dKn/sSg
xIBOYCgZ7LOCjJmwvrgsqWBNKJ3c7rwW5LIkrmGqzrT0e5LJOr5O0+mBJZep6g9v
9lLHaCm15YjrAkih1AM6Jo1BkxO6ue5WZKJO5ZW4a1QWV++OxyycSpd9nmw9aVsV
pll+FAYeSP8V2uJ8unnTrVVOH9c3xCeDG9oG7aiaAd9FWI45gpIhzwnTaJAASIc4
Un68vWYL+pUVMotQWm4CcjpNI9QQisg/s/u72NBKXlaKy0/Gj/Md3DQtHzejg9o/
pep2W6adVewSrwH12kY72rO+oi+teh325zJQDc0WMq3gqj0jUCgBxRKTalHpDOy4
VKVV4wjfg8YLj2NwAzwaIYxKvhhsQlmYM4S58Z3LD1qOu0qr7bx8Uy4KyqRkWuX7
4S09VNvxv3daAy9Jvzs76fb0lPZLMIAK12Z1KMyQN6PxID7ZSdanOZdwwyxVOgWK
fkeoQD5D36j+RCsnY5FXxgMrHeUuSXxRm5RmOgHIjwZ2z74lBsinNCkHjAW54LFM
PJGo/j7LO3253f8wt6hOPnhtbqqbs4KZHMtOwHKp2cptvSkYtbuPRwIdM7LgxS28
CIAKePM6UTHnL98JSCoOXYFAiIUFMYpuhyEDsutFjIexBYQv9hkVPDCT5JUqWc6L
yBIqgEhhOx+gaQ8tnAxfC+pDQjb7WECAgUkU2Iuw348Xf0MqUU4iITvHl7zXLwiy
Yf822r9MnawLe8qHRkigGJPVazdH1pnJrU1bg4KElsAMpgHEKvoiEENEOBjxtENx
jVYhRc/Vc5PCHqueGMRT5N1OqQuIVUnpxsG/C9CMvO+Y/zLuejQ4ljSkPAbbCM37
zKDUhC03on6A/N5OY+QZdj6fN9d9wtNFaDqjcevQko4PkIm96tdlBKltW89xzjRi
WdnHDfb2+OrbaiA0fJBTAE0BEMj4cPgascUyFImV4k2WSFqN7dCf+8EEbqHR6Qna
ybbcizN14zZvaM7bJjQwBLJ7K9tLF9CSr2GMlRypXQZDD0h8rMPeOkXLGbVRlpIJ
ir2ciCNEZgy++w7rQwgDwI2F6vfmBaguLzE6IeaG4aj06bEDA/8OallSRdJfS8lI
ndG9g7qSu7DSKepVJ+9gp9pBPtW8xjlN5BqHfnYshhZKdfJSnjEK+H8AcICYRlNG
Ltwr3+BjBBwF5E4lf+uIooPfT+RlwOvziMkpbTBAytjPp9N2gccz0S+DezrjsWjP
5bdOi24i/ezrw1m8d2GavQSQ2Ugvk6rEmAHobt7/lEf8pa+7Y3zCB9Ssb1D7MsTz
KGLEK8NUnTQ9r2xgZXPH/XxEwGXQ4m26Mdk8Z7LKGX2VwJVWG09jg6O/FgqwLnkG
ISeLUKBETeHx2cu5HFRScqFB9Hl6KaHAFobUp3iJ+YVSJLh10D1PMM3lD/gMmr8e
OcKY28ae5j7OjYlMpjKzlsG6dnIVVaemaH7BhFfyWgzaZ8xjJZ8tQHkgLy1/1kI3
/8MDW15JHQ8HKX8fMdsntYzCtfB4BzmxyKC2LEW1Q/3nvGFvJByYIXSAWyLj7NBp
Ccu0Rvcnykj5Ks6NxqPq1td/Q7e8rtXF12izZeoLa5/7n3R2Ul4EOibY7XmlGnSA
y2RKGdFFNNt8K4jMz/AhaV9kkQ5fh9WM+ZVg9QoFlCaKmJcoahLVxfP7mtcRKvbD
2hRS6qkbBnjieIK0pCy8kNd+xKhVTXVAQOeCHpV4bvRzAkMe71NNZ2BDIkGTEsdQ
v76GojkqAedhbC7NF9Bz3giGsAsgzmD5iNeNVxv3N9R5vjVZ7wQ06wlEAjITcQNY
L3um6UyquFzOI2R3aFaoZEXurt9GeXV+u9obna1znBnakR1TTOk2il5T+hO1+Mvm
RRkBoRavGjdVVO/laix2/9QciCaIHscQbvo73EG408Ybv2AjogC/3oUvtxuvVF8Y
FKKgFsHhuJDZ5NvtfLibVcsj0NhrkuFw6blKQUFn2J2yobdI55p/EJ6DmQKGHJdL
Gb4M/fneIzixZDaNUz+CtDQddMnLguKSzQvwrtqLNFel8RVHZnVvBvwYLDGHUv07
KwSmb21qREKf0fqYJmm7tcoEQsm0f9cF7Ta8BTKnm8b7EM/teWctL1XfJk2K02GI
Gsm0s6SIKhNAh0Ph5RPq6hAtDEickFfvMYrVju6/jlgcGkE6stkRY42KLW5EZ3X8
mzNp4YeKvWlQJrZRQ8i7ZLB6tpUNbUNU8CBt0o3spckSgI9//HSaVhQuoZ/zBHV+
7y9bApVdXXBHo+rdDy1Q1Z6wDGTY9+hjHppo8hRfgL/Ea3lfBNEtTVg7SacOj+NR
xcZCrTBrnczoO6JV6uwvwcb7yljqupn31akdcrEUVXXDBmSNfWMOsQWtAYKRuhqB
vSaAvmwBY5/NfNXTrIBWnioYY22NdAuxd17LG6De3fibhzTkjBJUyCOt/ceF4EDL
HCY3JG0osfzuNDInm8BUQO9BJdFoKV2sWXoaTO5IAjPPpHcMfHxnsezq1TNYna60
B2VLUXAT5plDcnmaJb29PUJbY1en3I2lIHwBY1/aISBWv7rWsvIqgJFpufNZwi2i
F+9Rwu9FAJ/OdaOhuVv3W3Y/lxanCMIZuQhtKZcYeuAegWLGn1BRPQQtpTGzlvxe
AigUdgNnIJ6DrN5XC8I2Fh9k9z7WSHcaFCOze1IogyEtTSMPyA0nwEhWnLiu4Ko9
AXihiaSLpcSBMT72I2rm43oTvRvK3/KhA8VAWxtGL3Dxlu8lOtw3IrKyekh74DoW
2U/sACZVEt2lqeUYsXvaO6SXfEfnVZN9FBInwJS5r4z2I3onkfJGWsng8BYahT6m
Wqf/MhX/gibRTpbpAKDbafHrPH1d/MZb28X3Ojurhsbuxrap4SsYBwnvtG7+lijW
4St+hHNmiC86ajoXXoGTpV5l+PvNlrZqP+ZsBMnNxa+9CFKfeIRNgKOOYlkJTU4y
dCOzUj8IauJm9PRa2g168sJ0lIPqllz9H1ocYZGAZCVzMi95irZtw11c8ShUofKw
KHIiXaTTjigOn1/6kNGeIFuPDhW6lhOt6YTQf5LnCiPU9Ub3bhcYU9iMTqV4hkBd
ck4Qql1UhhLCxaFoj8fWsTfXTV6MR8Rpr30+PJfaBz3QI3DWwfjpTkjL8Q9Q7JI0
Q6kOZZz6Nh4tqSqesbpKSVGKTFyJPghz8IP4ckSek+hoI7byNu10to84xykUbejt
srMCQXJDXdTcsxEzM0GVqRuXdRw+AdFKQBKh9xFOi3Mf6Jnn0tsWbLWsgybLOIly
I3IvgwYu/CoeCsVjEpPnz+HJ8AviPJi2WGRqOMOeSeAyWF56L1/t/eQnfe+3UoZ9
aUXTJxfk2+zXW7W6bplfjN2chPF3HaBCUefKUBjfRHsAYt22B78EKAQ/CYhqIGyQ
Wdnra0G4bTHOD7dtaE7c1Esst05g1xVPTEQW0fEuUieZBJn0sUc3W8TG68hszb1c
mQDhNhaOO+C1vdiiZkDwnx0wZ5BaorVrQce2Y93xqLCn/cGAP0QGFiCdQLMqyk0W
AOw30b0v3AdtKv+ukhvBurU+g/86mazjPLJEDry3qxSRKRv6zPqJd5XDGR2PZumU
AZ4yzTTYsXQ9byde+WVmTCA9yfliOT4gYviQYTw64boIYy6o+FHr87EMFkf9gk2u
sZSOO/WEw1VTAyOsvROtSqFW4DYLVW+V03q+DhrrZceYX5uvz5U1PZN5+Da3FxYK
3yqBSD6cZ2o/X3b/AxMq/8MI/ZDXA8xRjQvLOFcd7PXcj+JLgK2LabeLxDng29f8
/k27KY6sLFtcEJsmdyjuHQnpE8e5VgjDihqbz7R+F4h78UZO9GzEq2+wVy5BS2AA
QnJP1z/beLZNx7YEq1V4B6iyAijJj2Mn5AojBecPOmuvudfEpXge5L36tSS9X9Sp
iEO/pWzp6uvN2tIFagY9suiQutDTIw2Gf/kQx6AeGoKJGaJknVoKjobsCaqccwGh
boUOzkqim6+Am9wvTQMJA/NKrdAHo1teZLMWCL/iXWRcMHFwJlfQy9vjC1B8+Kzr
DCvQjNKxfnlVbXeleEUGdilR+cfJlHvV+sWht+LnHjMh4lWfTAc/GUnrZoaHaSgu
o5/udtHRRObn6jicQz9e79QDlIe67HLSD6gC+ORjkkDWXn+OerYXNyV6c2athbR1
yZmn6BmfgyHOXPJTBTlI+QvyG/STDEkw+KwdzNCVDzUbyL+tCGzn3YliQ5Ctg91X
rl3WADf9VCJFk0MJyzZX7lGzsSM8z5WU5Ad+Fa9L7po4TbsJYMDmZ4guY3on3eqF
MQu6qfHgRZWIr5oKkcekuILIRJQj/l7QCcBTbKUxObBJ0VQPdH14Udi9kveQX7Nu
m2G03U3sh+1GEdspk5CekSd3dmEdO8Z8qgtjEYDmPbfnIV1TLoS5Jk4MQU5V0nmB
DBFowG9lkla8o1bwZW4i2wf8OmEgM5bzHwLz1wKSGot2mnR0oGe2VIy/4sCg9HXg
RkdXfeXviYrc0ffIATWJa4srz8rzBii7ViDewTPidJUMzw3H2uZNwXUrGxqJzomW
oygitF4t5G6oOARE8/zK1VJB6K3gQgKBv9fvDD1W1C03lm4HOaK6uyC/+jj5IfH4
WrGL4vUKPVpufUXLpDTqsBQTMa2ASdDxJ5oe03l7iS8+ZhugAzwqt063AC6MXiIX
KjhOrAPY0TipxfNQk90vcm+ktVRg/Ysg66Pqo0CYdEK1kDw3c1ETws0Z/KnAgEq2
Vec+o0dFHj0lHQvWTzTim2F1op6SoqSSQC+OLv1oBh/CbzKDzVvwQHFWThFUBDDO
kBhku5DL2NMRXQela4PuYXSWW48MLM0Fboe8Ti3cxr+kXycQ/ZeT3C2vHHGJ7m1+
0Qlb53mVNVenFGdeqgrOk777Uzm6N6N7HJ3kn36kfVOxDXObFHQCVRElS0+4AFUu
aIMQdHMpHj2YEq950LLwZvaEgjDi4+TUzsAufIfTv+AXNJjDtPyU3OR8LE7+Iz4Z
XesiKWLetWIGZp+m2MDXSJsMSn9hhq+cbdOE+BJR0PdlGLpDaLJLtG3S+1pPXb5V
xdkrwbjUnhovgnffZKXHor+ytaqcjp3MUa5AoTVjwHpxow63BMJrrR+09yhxN+51
5GN/PJO2v6QTazDGHxUQ/q0OX3Ud02qupHI1BaBUCUZ9qDY/S4AcGlzv6xos5QL8
OrV8IFPLbkbAJpVIuPnLd/btyh3I2YPO0KiqLRIiEWYXkudDURH5HSaqs9TGrBCE
165VnfQMhqNfHc9+OvMtahoa/K7H1c2NerdyTv3GNBQsiCOUpZqalw5TWGl/+MVw
wOKUjLPMF3Aiv110p3L1mKse9ds5ckJ6vD/YdBYLe+UWzqFHc4PLIsMymeLhgCEa
bb1cFn/Exn7Lm6cEXSiZC6VIU8iW0WQzGU3M8Y+s+9D4ubmrgHA2Z5vgH6rEJXwa
42U/6A272P6Mf7nTu1qaBDtV33LSNDufIK2/+Hv5EMxiuqT/UVqeA4VpTQ05I7P7
XOFGcSNPH15qz7CBkAyCp2/CoBUbFkgqaFL4hVM3uACecOHwjrLHD7szKeNfUWAd
BXT5GHfsPve3nKOOhgNLPGYr6Gge/w1NtAN0xkMfhroZuTtMjtPKH0GWWMJGK1pG
z3SJfxPdUMorlkAw8EFEmmiOkUPgjwaXKpdy6zAgPinl31n4lj1tixhTp1UB/ZE7
3H94mVtMErZnvI0swDlEkZeFvTtSQhu9fNOuZlL5tBZCbg/IkqYrKWh5xUhrhOyH
yH3Urtqg69JVTZUZZIWstWj+kHV/aiwWDaqjG7IaKUJ3HSawbMDAKbB9jsqgjglr
xCA5XKW2+Ohw3IcoFC0PYJBAlHpq+jTkL0BrwJChQ/sa1PhBu+3/I/jv5CSDvqfm
ucAZILxBEp3gwlK332HhnIgrJv8l7SgOq216T7ubzKRfKwrshhrdhSj0xNdJDkB/
bpeIZZbueuer7PVqtbPGyjgu/VGNFUB7t4WN7rTFA3mKZT58zU0D3o8eHPTZeoH9
9i3NtIjgpeem28+Q5TVD4S/NrabcxAK7ebOl6uHqMKNPIdy9cnGWGmXpbEmnTvDK
hSkITXqSzuCi051c+IkIeNJz5+wE8d88AWLpYw59pjUPyzRwbTbOrcGlDAtpzlH8
eGhl2DgRWDkM1gTm5c+8qFuEMYS86Tz+SrjvUQ9GFavR8b+z8w+HKDVzaHV3ltRX
WhQZfbyfYEUwGOowcdWVRmfHntUqhUldj6tbH229CWRy5WkKRpJuPsLwBGz8+UIs
0QNVP3/pjg4k4s/TIPgaNVoEDHDYXmrwhurC27ZMSZrhOaro+7BeH9immsLdR4qV
VcNYURqvdexdMenRAKQ+UddJeqNvizNeJM5xGOkq/jA0w8oWiNO23vQSpd/5o5Gs
mAr/D9GdAvcFawZeu78NyiITljK0xqf4+XAXyaQWfexq5qZPb17aTScsTvXnmhZI
lUDYiAFghn2xi7eFGGvhB0w4TXAbsmPkau53l9ZrhwLPtHDyPshVoA16SHGSWdBR
mb94kLaH61oJJKNgxxOYyb7LJtFdtK/kVDbKcVbcfBHE0N09p2+Rog51qMSI9ze8
33Qmxcm0E/H+L2F6tdbRiBURJUAxrlip19McT5SkwXNNXqZr1rbxjtI7W/1WK2KK
lTQTsFoTaXb0w6MBLB7GoIfbmJtJ57Bv3dMWWmQMzSJKm68M86Dxw62Rxrb15QZC
nQ0bRGtqowaRAK3hGwZmgyhidfNCzyFqF2OCzVlA+atfOJ75i8c7C+k4aR9J4IbW
lQ+V56YaL0aMuCxeq9oXvdT0kCn7J28gyMMDkNbbyLA2owKrKW37FWFDaCIEGJdu
ITZUc/VHLkOd3g6JUERKv5pfl5W5OTTQnQzL0Y0/wXUnuLyeLRgHUPbvEQ8PwLgg
THsh0DlOCF/XoGP3JP3SbMO89KdWuIAig55Rmq0u7MLHSAk7gDyVqabdJjt2Dx3l
a8yw5zxvp+IsypUDD7zZ3cx7afU4yq91hORUuMLLXcmitdowFt6YX9uoFNwryEGC
Gt2U86oRwflniUwTI0tUsv1BFo39e802jHrhNjwR29AOIJBtftBClBjhe3aV5pdG
0VmQ2nermGeViD2+vQbU6L+Ll0cboqH8T23Q2FEZ/mzsvlOQnhuiwxPXqAfUcXAP
XjgkDwAVWviQwSJ1zA52uVG9F4VXWYYVh1OeN4WVV70q0Eg8zeRy6dKi57EUKviE
V/nEK+vLyx+F/TTI49KD6rRubbcKGAFSjRjCHJgCjII5ekPQBlgNVHAMAoouCWSK
KP4XgZUr3Bm6de6pup6thFNflD5iYxx/61TyZPXgTrp4crt9YAiYfGszmmgo6GzT
/YzluWweoAtnoSPyIN+JJn69lHCNiHsr6PY24A3xVJGDplZnhvNNPjHLJ9bW6Sop
9M9DhFdXbBklUK9mXK5JAlZ5m5l4wLUUfndtag7jwGoVUrqiaE/89Wttj8GeX+j9
S7w6SaeVg0ezhoKo/j5+4KKXpi/zSWy5w+hkpQWRScQ7fGG6guxEDiEjj1guv7uM
Slzc9UWEK8NHn8gNA30hQfjQWFzmrpy1pG/TXbgbfwoawLFnB/VMKa5bQslsonjw
W7ZIoC/SqYfATBoc+5o/s7y8N9A9SGVXx8eaLmY1BmdtX3BaHw/JwGvwv67CJxs3
1lMwQs9Z7SCjfsWfzYxb5adYfyoDNwwzaTJahP+l7LOrq8uSabZwYRT/U64TVVOL
Tc7EWwuzJy3D324CR2XpUiQTRt3f8JzfZsgbWflZiUsnEbJXsBDjuVntI2gxAnk5
hCwtqGCnw7XtWrGYUZxjWmVx2Zti5zHUgg/MvVc18J80D6ziTt4DVoXD0rKM0ewF
Duqo5Bm5Wr2IT6jC4/RZ0xevKeFV+YZrAL/FTkSBzC4ydkAOdUMcMqE6JH6nWyD7
pPDsDv//lzcXqX14Cg5HDEBmnt/kzmsSHczPostcARK+oJ0tlZ13vSUZWfm7Q2g7
6mhchTFGB3YuON9SF2a8zg14E5V/daCx6qcxNssPUdA5pLHumCIxvoOfOtO7h9xr
1lw5MLQ6dBuI2VSL0zpdJrL7VrL2wgbsGmZ2ropJ7xoIkNFVp/BQ15Y2Y54VHqSo
KfXGhQylhfl6TIGCL50SPPgboZXURRpwR9liR6XNYzDGazNZLvQgKKWwQJLTq04Q
bNtmr6BiEIetYNnZ94Nm/6hGFWhHQf/sqos+fPU4KnNualOWaar6dKus3rW5e0mH
y0Yzu0vBQIF6ML3kFLx+NC0Amg1aE9h7bQy8Wo5Vx16g1BZbOKJaQ0BiYGG+2X/J
gdImlIFDM1SobCwtOlZ4kWkyksmnZSyGOJRFShB2JVaCl/NSH9xuH4r08ZWSH/yn
7ELpzsrJmdQW4CU5womvVCHbrNkGLfSzHy1N6K4kOi8UdZkD27whzrjB1oJpV0Te
pff3oPEAE2C2GBn4dMGVZ84ydndLNsVqO90cXsIR6W1DrAny+YjNdS5BEFMMS+WI
T2bvORHXus+N7ieztu1IjIXoN+b3Fs0wbV8A6sCGX9c9UI8rmAtEoXXHo9GVx2ym
DDPPnxBo+WtiU2Vb1xlV2xsg4EaCyldGEjUsWA7uVuWbaeMxZy9CHt7FjIbk2OSf
vL8+gxg2jtsAQtApVyz+9Inj7aqAtD/MMGKf6TvnTezIXT+5dvHrbZQgpyKtvDVD
s4IXpatoTd+A/2EuaRJgQ25HudoIRFRH7Q1C2KdIyHNZBy70AXoAbEt++28uiMnR
Il+HvzUybttmx5LPNlj+lNeLUsx3C9yZnwIA7zfWVUp8qOICcQ/gqZJvySfNem3/
kiYOyrGzZ0ijiZr2FMioCi/IX9qR33pbcxiWEVVuax2rYgKmtJJexJz4gG+/Y/lq
Jap03NIXgIGR9pKS6ThuamZPR00vEL047Vy+5mksIj5n9x/kEKcN3Yx7R3nyxjMg
BwDQFzgA+t5tbuq4FwHGfZWWrCKWAjRIaBPytsgGSzqyje66nWcZgEgnfgouKJyY
1IG1kxtSi18FD6r76GDb8f5TPLjn67/MKgi6kNbZjFTfE8mOWcSmFNrwrXOAONOv
g11TtfYXtgevgLjiP2scOF2CQjiXlbFEbdo1e3+Uasds5xEAh0iwVNFxRNRL6c+E
0PbKo/LoCBgm85r3MllcasI+vh06hYwtf898kL+CeJbky4F9bSJ2LtqhSRYlLBj9
6Zo0phvg7dFy5yIE7kMvUh1peG1ur/wHNVI6udaSGlFaTJT9ORwUZ0lxwWRog1yK
JG+QCCXKo1LBQFOmXkkO7zGFrFupDP6BMwJdNn3QS4BnJA+/2nWayOrA3ABnMeGX
xTYVfdImBITsND7qRrGDLzqjqBXS6LAZ3Bz/aVdVzQ183LuPhPnfH0QOgoyLDZ4t
eflkXKCEbrGUUvHCfnz/9dBAZapthib631KPQ1/ohDg9fz4OlcFoy843wbMoSu5O
nU1lMDl2WVez5zysAALMHSGFEhoiX7c3uYBdYrKIo2KsvdFJltR5N5TiWMQj1Ptx
tKvAXm0XPiRANN9ypnvThezNu5iPzg969mWQakBQJGMzYeMMAhr9nF21CI8453Qj
Dz9D5lF0soyMta9yrs+FZnNKvbsodEMYc/kIhLKLI14cy1rhOy3h1yRKM7VY8mEb
mHTi7ngZVn3K2QvLbXAIBQz5l4LIhKKnkLG+a9ypoXDYuUl9ndOBQ3ByrvKNhGb9
w9cTfkEv1pNjb2UO4v6aigcKgdBfOBoMEbZSDSNkYMLgvgqAwbfKCC+KgnC4GZFX
E0cpclMfKs5eyVfZKaObMK30qObINFGdMCeBDcRlbrPhu+c+TTz/krycgZQGayIi
PhuPxGof5I7J/Hap8l7C40sMxGSu0BOaCz79ujavNk2Hgab64l4HkPETCukS1flZ
A5lnk7gnzmujb2OGv2l5Oe+qj/Tl5715eSZv1HvOsYgVAzU8t4XkVTrUGQ4p241x
2dAdtkgDrx+wi17dmvohXD78Aw0scQKbk/v6ZOzcuYlPWA83EwCtaUYVOnXkPBXP
NEVEmYy6esxpbq4lgIIwJS0o2fkw0c4KS86yqHy/KFklJm+nHbVXSyGQa94nm3VM
CDOPnlBtGN3l5eoDM6CUMCWW6DdL1AtXKZUdRjDRaRy9Nmu7j1xPu55Ll++4UU9C
ZTuGCEbvzuLMGmcdS/+mYgKi49illyiwvI/vIt7fVmPuI8RWYFkzmvk271/xtucZ
0Ecvjl7F3eesYH8zaFxgaIRIZI/YY0pts5gWH4iv0ZwWvWTIhhqfyzk7vivRVdAJ
BvpK6ACR7MYtI4esNaBTAmKu4akkPMyrx6ZuL9b7CiXt3XDEEAeumcPQXzKEulSD
ZZRi+SNgViCcFqEr1dkqezUdnesLXXykZ2My8s8jRpZ5+xniudf0mC6Ear4nmN7x
YfkT5DDFc81vYdCqbQCj9puQnotsWVNP/tFDoOHZdrHe86YKR83QKRbNx9rF0ql7
5OYfNmIhEi8e7ut0215pIywIK/78CFGhpcN78j5AiTF1Qcbh+QrY49dsuNJbjrLp
dYU7f5Fc+THM31LuW/JAcsDPxiDcZbHaydqC8Xes5hi0QoinwFSKr27OKxgJNdXz
e9dFiKE6CrL7BT0nITyJVPOqvE/xiiYNjgJydaVjIlgLUbJYRYgkDZBHzdYicTZ8
oegqRNRINYtz94Oiq0JrsoWfjFhB+N7C37CrfCUtnhLC1sQod9aWB3Icmh/2p1Y2
d5BRG0w+dsZL+fxpdJJKok0zABPOT5GvhiaV0kn9zeX9Vo9xPxWOaLNvoeQMOsVv
GxpOoaxTOzkvKp/WuLD8L3MyGxgtpAJ7QiSvMNWFw8uTuaaXeeAYZi3eib3l1b6D
L6nc/eutquA2oUt6FCuXJ5OGBV6YUOKAKxgPQ8ldQb/Wyonwn7Y5xX0iN6+934CG
igd3zDpFiXOGD56+tK6n44RT53oDX6jOtzcdbzOVxTWUuq8uD61EdeoJ6w6W9plq
JdQsiwV9onZmBti08gtJzbh14BifLUgNfqeZkMLzmy7Sp8rdy8Zioj6QrsKnWdL4
O/1ROgY4OJRf0bcLV6b0pNJIB3rDySeeOMy6Jn8hssqGTKV/uo4NhAM8ZX44l/od
by08Vqb0y8TIrvJ/083r+KlnOjLwEjcUj95Tq3HNxqgmN9rM3K5onwUexyuU2Dec
JLIkbn+JP5zB0lR0IXFsBZvKt0IOwNP16jhmm8wauBSHB01mBGuQU50HgTEapYOJ
ko0Avol9ZfFsmLDw4h5Fe3/BCTC/7qLVOgThWpMtcfnUYCKrT2+7LqGa5GXYZD5R
hhejgUIIbubyvODNyyd2BaFfnjlQByP195FqPIqgDx+HCaKvkixK2pymV8kA1aBJ
p7cqhUyGt8MnQ1hCNRNZZ8GeC9vMVbgY21mfONbuq3mmdIMMOP0pCRVGiv/DTMKk
o8IqAK8yt+FzymQHGHBCZuY9Mz2AEDhpSIqw0GqxHmGzfEws4psk54ziZrfEga1+
el6OUeit72qI/yE9kdHzkENQw1oERJ3C3l+luDLjzg7IJ0kcngi9ImDfeG4jqM3Y
BjabUdF4i7E4ULxxkLYEtKDNEkfVOZ9s7Kj/YrhVxlJgu+wu17rkIB95GSYdAi5D
XS8MLD3c/JfISV/+civbZwTfXEv0OEqKxVMVKsKaFB6QMZXvWZxHo17ibcZh9ZIQ
5W1EGDwlbQtbEAG3cvx/b8hO8SLqflHPl6gfGaAGeF0IVuhwveiVimRfmG2J9+ND
gYwm8Eg7lrMPiKLjuevddUQjuRBn9xbyga0A5l2Ur9T68Jj7SWwnNf4O74OfBcBN
FcvMyQwQV+qN+Y6Q57sf3Z6EvNXAMAA4axWVC+YJhl4XZyKFoizsePHA06EYFyM6
KHHFUmLLRNtfyi4qKI0V4zLMccayRT/Nu7JKPp4XGgwQkbBvzf28lxWmO6xbCcoH
ki0PtK1qr9dRp0W54KOFiS0uAivbktzvZGDZOU7IHHxkBFoTH8L0kzx/aC6HvzT/
XB5BkmvEVteH6DTj5D0jpT0+F9ZZsIAV12it9pR9LD2avtrLgy7Y+/xiZeNgroYE
iIy3yRjCKjIqC/GUYnwSVqfLZlBxT8lO1s22T5L/v6lOfK9FdCPITRp+5N0crXb6
vaMlYlPAnprML1YLWqEfVaAHNu65iNkE4Cj6Ugby1KZ+lSGbaOQ1ClxHpxQLwN4i
uAM+qsFAvYbde77OwtlTlCNj0L0CDYQXM/5bl0RO0Ha6dh/ofEZuMutP7GZ7bACG
077KjqvqejmBrKqP/+BOzdYB4ABJReh93P71shZ0EAMMAKuHI+S3EB4TrgbPbd5f
mYOO+m3RLesc1G40HMUOwTCsuRqm/unyOkoN6vtSHHuBnMS9uHGQGra31sjCednI
jlMdFtP0/DozjZ9ibjiBTUdN+mlgl2AfsyWHaoTDco+ROdh81snxFJOMnvm1VYHV
ZYlQxY5qQV7FV2vcqb2h+b7fx3JnoQG1QbqA1MvSzQzOA9QW9MmtduNSuljD7QP5
DW9CiWO2ntkk2xvkUMxMwBPBul8iUXnNahGqaZZLw4GzL46lHbo5q6iYeDYswjv3
vQ3a2+rmnJjSAdSf5LVzigyBJgMrMeSQlAZ/xrRUSpxHYPbYBogUUTrnYEs12zcM
qrv2d0JtaYTeZviLvd3tZEY6iuZmVqLC79P38T8yZfrGHYmnMWrRnZKwbBfRJwnq
2zTp2mdeEMlAli21Sw0GZ33o7rvhIZQkRW7BQ/fJ8H7x50BDxnl9UgAiukJkadTY
VuSeRB2VspIcV9dbfI15aVepNkIsAvo3YwMtvK1MbQWMc/H5hLOsT1hsuN6tYGHL
gJZjlVVTngSTxC+z4nkU2b4LGkTcoowyoJkekxY6hYRXUBgN+TNzRIck/ZFM7CX9
7pipbsJ/bTSiamDfeisnHkTM0Hj1tZjozYG1Wmf7JlzJa2N7fFuqLvV4Xwi0SHlb
HmykE7OhsRyGQss8qeX2ZlBQvPyB9DScEDv96NhhWkiuNOFnmSE6MPBtgDYgmMPF
EAcXCLAgyGgGQOAAXw66v5eQcnJJMxt2b2ysV9BExoL5XfZhd7eA6CKvp2Ur32BZ
oHiBiUQErtB7FD50fCNdwBpG1DJPgwd5OLiosV7Ud/gkC0oc+LAFVM2Ri4hdhTs/
ZVU6GTdWUQWnt/KujPZk4oRb5U5Ebig10DKNyBohlyyuxF+4vCDv9iwoduliN2TR
DKdeKS75llSFA1rIDlfo34PXnjrMr0p/rTa8leqgJw+yByluGgjWA2IrfvCZ/24E
nVlSpk+VDt1unwM8nASw1QThRN4ycYXPZKOMIz138v7rshLbzZQ5gvUZJ1hNxn7Y
xMmS2tIt8H4796mvNhvuqY6Hvby35qe3nk/iQMqYlqy9eod9sOCW03nyAEqOVXaU
mHFLPpbLFbFjKY/WAkUh3ElD6Y8jpnsYslQlqqpZqJ4mNGT2nFP1F7lFXDQjM5DL
qne88WiowVTooyLEjfcsBq10kYXSQ58etTWlm7KEYG7fpRg5PNSP6Vbtgthw9S3L
Ws735jXuN2MHloA4+415j45ErFTX9Zdh/4SQwDLJMkRLFyKUPB8kBMw29Ro4OExC
TPEts7PJtUwiG9Nt6Zm25fz8kXG//Eqlgn+JT05UDHmsUKbLYhCRCtD1A9Q3bW0+
E9tsL/GcksbRHiU4snnQWWnDL/aETEWe3+V5Rxuz8mCS+S6lziG1bIZflKEl1JRy
aimBHnJ2U9xXqhnvAIYgQQM8jCGCISo03OiXBcGhvkyzcf/1Csh4C+xmV0dc+axO
PRW+5WiVZ52LaplxgmX8jGcGZ0BQYcc3iQY4ZT60mZ9MJwfekXaVdX2GVY4GXRy/
TyX17n6GoqLJQi5BmFU3CrAX8zrqKwTxqvrE1Zfd2OjtjCiMgebqZh9qS7Y5jdvk
Umy0FM8i3Qas0ptq1P94PqU6qPS8GuEf3EIqy13jp645EkI494DXcZLPC342HDlB
gchEDQsAMAU7k4z/JPfTzWGd8cNLUXoyROWyiu9HoIh7U2SnHXcRKzE0CDCEGBZB
X3icBTttknYtdKZkzMguxG1xdh4KGkIfFkiJB3VIckknnLUiKOW5Qb/XzttWPTR1
DqKblI2ak+LABukxYudqSEmIjpE/1hCwWS5dVVQry/jjiRYe87ZTpF6nCAI0znqT
LHQ44vItlAY3IluHKHJe7hhL1hDZ7nJTJ2OjIz4+bEVXn+DdK20qeWMxjXrO5imK
Gt4HzNN6TcNifJzQF2mb0/RKuco3WRt8A8njt+Z5K9YGARVIL2q1F5fN+ukzERVM
TLohawCyvNUdqIcTLaNJs4FFuylvkrZrW5iwDgu05/shZQnumAYe7kmfoo6bEI+g
hd3SVEVGUNaIk9yaBeymiE8xrNwlZqlCZnRbrPJjEQEhhm1ZvwpZbMtflXfR42va
uyedUEEvBh6e1q7Y9d4LhmuZKKE0PvUlWE3AHPIY9U8XNb6Qq7I5JqNaGo7dMEbT
pu7pYnHxn82eAxRz7Qs1XwLP9zkPRdVDRnPJOuUW65UBzyD6J22bVGNIWOgQY5mf
nvuSF7dz0DY0LFLzLGF55qRrz9pGdQmztZqdkzIbGFvl3iSRoB4Gv6Zm4oCpP5Zw
N/L264s5DjgUJ9Ok1AD3mWea7hPmpKjuUxi2v4OWL7PT5KitVN+x73C9cRhmmxX3
Ws+e7ATWJI3V4+zQtUsfVnNSDu9fU8OTI6a9URjpKOIzTYxR314qxsqNuUlG7gwq
+li8t6I3b+0EDd/pbitkjBNL8o3TM+Rk3yLZrtpSDnh61NesAlivUw/I66QDymko
9TJ0OUgQPBlFWf8kR0KTc9XsrGpEE8sd/ZJYIyTDYPmOJN8TVcqPR1Zhmpfwk2cm
oUoGreP+4kTgHCXB3KUB9K4oUNmNiMSFVU6SDqlnfLej6nr8JzYy9+WysWG7MifI
zl0HEbQjf1JJX7tELMZsOkIItYf/5XDv5ihSKASrwq9BDaByy+KggTDxjksjkKHT
B7OI7OPS0E93D0cclm0Ugo7K90X4gpB/H2x/Q+e9laY9MJjSn5dTucz0REyjmHr0
pK7IiIo7+W6uaueUJpzUgfX4LOE3ygvenQ6g0qiiB2Fvz+nK/9ZlT28beELnrBh7
0pbquoysuEXyigRWMHe3w5OS+TDC6jFzlvOqQrJiLxyol/YAse+4gCeudhw053jS
hO+5Nrcj4kReAERCR4nrzna/LnLqAmCTDgmMXQGOHGfkUBT70VsIpqHwdnJx3zCl
L3nkHWCeGXRCYniNkNMyum+tiKTq4aOEGMU3hm+2SPvRDYjALkx7cX1pC+z0swBQ
/ek6xV9g46deUUNj89T41+iPznA4XQJ/S7CyZF1upP+08YWA+c/grwBCaI7DswlN
PYu5NbeDDEsZHeFIPm300bDq9lWyz+wBbh+xmEA37yEqjEaCn3b2e7VdYg7O02EM
yEf3HNgvx8E09hgsrtkUj2zgSRIUSLR/uMg3syV6jbYH2nXceH765kL9esAjNqyX
cz5YONfSfY7PGrCZIterISqlyfW2TeS/cB8WzGkWlaqPlDLPvO6qoIUZ2pSYFUzj
CFXUNJV4BQoJQwW7ZBQQ+HxIeLLZLFBknhlGassM7f7SvqFgVaQGbXpBHaem1JuK
6UBkRzIRPIr8ryIj7LsZ66muEN7dZp58TvvBGhzfcpDGQJka/NbitwXFxTRylany
5MRaPcJ9iEHc8NhkK6Iu/y/oKFyZA6YoQXdx4X1k9dmYjBDOE8t/CFI69J2hbpPp
v2DUCN6SiZv+I8VLXssHClJXaa/0f/s8UzvyJmm+xaBzPVbZRWlm8BoW+3jvCbDM
srd29/YA/kVjnhX4ElMwQCKhbTz90HM0d5d/BREuQ9XHd7uzo5B9umlnQBy6Z8db
ff6YmAduDsY6JNxn2UAcSJrawRVo6RlnUjsOgpU6bmfqgN/JBz27YC2cq/fHpApR
qC+a60Noi/Bz4VliKlXGOk9VyOHrMeU71ofHbmwSOw9d+kNpSKKk/UaHRhmBcVGh
aon5iajeH+8earw2hXlFYxh6f3wXx9/wULn41YI1j+VWm4DaYP8/PII2gmA0rGPJ
Y0BFekKgxsltUWndWmQhHNq7RdKSGtvxYxrbHaw2wHeBqam3UECEGtF4cpXj+h7g
/7hhvrsWKNmEDP6LZ3/hiYe30LAZs6I8G77sze0k1yeEx+vC483wq8ZnE/NHt8N+
tgT3vAa8Jq/D2aE2tK0FTJx6Ton+KZHjndJMD8ahlzPYY0IBL+InfXguwHXNxkO1
hfkRnf7MTxhRYUSD5sMYfEwhTy0J0ka6c8/Jjajdrjlx56E9EraEwQ7s75X6IMed
y/h/m/DmwdSKyMQE9YpuSiUscyKFGos+vIJghCPCWTyoIKIeZnAP9Br6bjz42FEv
M2rJYX6M7yJWPbib2odO+sJpQXmhMoXPC8V1FaT5Pr2eYTA5wyXTcQ27tDHaSbac
SEjmJ4zt7DnEVNTAICt5AC+lpIQiOKeyTySzfu/cAYcUdI6shKITAD0RCN61HJ0M
9f7wV+BBlpQMCjVCa2BIwUPEv/gtk4gkrM279EICrXY6P6Op/dPxXmGOszcqPMQR
NihWB+v5+YpTPIRmCFrb5fh7zKAxonwruAz+Ii2gl+YXKhY0rtkprw0F8UnJ/b+1
DujUPt7rV3FUqn2BK+d4GTjdbNKsl7p1WF44ywcEVnh3BRqZd09k6fgK/geY8yvr
/hgMt3bO0YU/eisj9PwipHG252lYhuEBXJHOcQEyzkY0cjgtuqHekenSlWWR6IPI
CdLaUeDGz2iqUwNKg1kn+Yoj40r74wKycOGYnxmEjvY9gjt++8quGv6uqAHJQn/A
ZvRBCt76ZaIsHi3jNEwR1kKDefQCU90/JW5qaTHEHE5VS0OHJnZwY65kkuSWBHxB
f/mngTg6pB0jSFAhF5QEmmD5E1GEDcGtRW1BbH8BC8hxmT0ZpvUhnvv7pPGBVXyX
JexY+ol01eN1QdfeGPf2yl4z5JrltstYOoWiF8Jp/AzChnm0gp3dGmc8CDtiVOyO
st1dftyEqr+EoLZGI2Xmu1iL5mVggaFWIHiRQczjUUyjujuRF8DWIJ5Sgf4kx4Ht
cE6af5vructMfAFgWyTpEQf+rmxXH8fwKezfEDRp4wvZ5Yi6DkdIydCyXtQlsdG1
0nu02+mj6hhz1NUIXXsYvG0DmGmmSqeQwiR0u3xXfzJ3nrXJ+thiZF2GH8dIwq5e
gmVE65tor2IcZlJ1Y3otgZRfcu5It5wQONERSatBZ9rNl/5g0cTuniwOEOpvJbLN
69sw4grmY1qpGC0cc6HCF1J5wkk6CZw0tu0YSweRv9dr45STCYq+7luBT+OxOF4c
Yr4gGas5qbOtyWwg4CH4ToTEo7LpZ+c3oNheYl5KKbLM9mcD8dr1HGxiol5BJiU9
6gE36x0QgtaBwe87Hpucj61fOwfUm2nxUu7loeHoz1Kp7xQlVUUJdb9AkIekk4n4
ItUpUxADEYpX3rFWZlL1NUreEFQRdyradQFOJNGFhSJsFpDJkX2tgZKSI6ki2500
8akh2qSYmVz+qzQM5bC8WKgknF6zSXk3gF6u3WRYOjcmFXmJgqX3RWFUwsKEd3C5
JGnEG2QuAxJ6TNFade2T4I8oWR1Icx7PnxyFNFSknQu+Z4jZTsLLEEI7oBpzszLk
195u8pr5mmDPgFg53yMI36yicJDtwIV18BUlzmIxv2UGwH5SwTeYli0QM6r6Of0T
FVefqNnbSAYXw2QgvuOls3G3raSm1j4L+sBcKdePRFVbgJLNS1X6x6UaTpNEzPxC
ptTv4sRff9BzIiud1iMUWjvXwmMRNWGaXAQCtS81HVYlXKrSAteh4zRa4knaef7N
lJ664XAQCXpkxec+3rMw331kUMN1iHrD9gvrKxN+tzhiTwvVG+GQV1p5tLD1CKqT
CBLqDNISdTDhFwwJXoNVilxgk8C7B+7fAE19aE+h4dE4Ymb4bHcYRqWpOjKBRRk2
nh34/2v3HA3AIA0F8lOEGwoAtpmt+MtD1xwFLWfzx7t8uqOtu1hvbVxPHxkcaLTG
XuPJvCJfo8QWiyhtNbkYKBS/SUjMOfE167UOq6SukopYoudS4xW3Aw69bVKZeXP7
rVRDddWNkxlV3+CylRDjtIsAaTgMH77OYPc6HTyEIrnm9GWTewOeNdx0S1udEkX1
s5W2oMZmH6sNPlIZwPoXZhdksNqkPfOukdD0qxg6i7LGlkcnyHAo8+ycYuLRLa33
DhIUwyEE9B4X+PWf70r+IWiysCL+XNtedG3ateE0Sv/iwR7Uld/4qaG5t8s4RJzH
Kbaboa9dGWSiHLbd1i2Y6n3skREShRf9nyfa4dtkfXtAV4jEOPatU1YuVpdckdQC
8/Jhjv1hXVA/P3uG7zwE9XKK4Qs24wBNl38JpPlh4W5Ofd9o7AYYpBEjzwuonQ1J
hbHhKJPiLbJontO9P+9uCZMAleultZS+OPT2V7prcBdO7mNzlPBiqBeTUZBZI5E5
ioRwE5orbi8PNR7L0IqJxBG4Rgr9orlwccUtt3zeWZ03gl+WWUZl/YgNV3eWjzBq
nUxCd6WMA/U4fKOfty4ULM5i40IEl8QJ1JkN+xhyz5e5tks1L4c/PYzTyfWTKZ1u
iLQ7huxso5glqu65AqYrYZyWiPYqYKkgwZrEDhrlZkSFiVUHZFPhnHyzYGw0xrwS
XPOuF/OBnAN+3boNzXU25sVboc8Uu+LNj/e5xuQcxw7IhDeeCy5apNkHe0gOCwyK
BxtzYjjnwH7YiugVDXzUiqpkbbNT5K1o0rq7C1GOIZIBUjcWjsecoTsSZK1F/v9a
Vq/vPbReJltTbEIq/1BW818qUStyp75CZcfHiRTD2AOUqdssbNj+F0kHZIRsM3gf
sk4sEriJAzM2eBtk5l7mX9WHzSzFX4jYinK4a5lcituLahO8wE6KMH0B6Mg/p0Qe
2ikE/U+gyshZeWE/Ydj+7Xixdm1hqUtGdpgb+B4yyqB1JDY5ooGUuUxBiHaFsa7F
vd8a3SclDgQ64utpXI4mlakSDT4qrG2NXkt1l6kTdsR1Z+6DurTuLQdbb9Cn/bs7
JwJWJdnfZ29YHxHIvfjgztEegqOmePwuwnIsh3qmKPKD+UT8IWHblzu09GN9K8si
QEnfwePZIEemT3GHQWGpDlZV1XKPQzbRGp01LGfwiAfP7m55D9ZvHrMKbq59joFi
gOaKaPyMvOlHYfRoUIiTQvXq0rLzVxRZiWElxGvGeZB8PXnNThmgTdoUpMPGqf91
dCOxY7f8w49xgQmrWwO/LYbp/+JsaAyVqRbTCk9Hs6i/KgHzx6XNKdCOvKuM4sYZ
yBsQYE35lz5HJ8/ANIIRG0VGHakWHnU3cSuynCkzIX8+yfewwpq0NFEw6PX4NPtr
6GQoAiORc27EeqdNteLacB5TfUHSZFCz1n2Sak47JErs6Ro5YfVdZBfsAmMjmHJY
J1M0NnGTEcJqChXeR+mUugeXZastz6+AOFWkOCe6nnMx78zSz7GQDkPH4GOaVIAj
sqerTacIVGx+VJYgF+w5jich+90WTvpS7XjyRlddP7oc9xpW5bIk2AAcdEMPvb+x
3WYeEHw1HgrNOu3D2ccyA4t8FF71ASOo0lM6JRqmONHNXdc0ZtEuYTGTvQYr7OWR
nRKTnqZkbneLwlhpn2/YvNph0+s1I7EOW2Gyyvt+tECuaGqHAPnYskMbymvvTSwF
XU1eDguFJ+acul7xtDEjxyKkai3X54vwT5LqSpuh6VOCuGvIP9SlH5GV9i8mwuc1
jQxFrewmYPubeUKv/oGJVtW2uwn1l2ZUD/DiZwhf6x35pN8f0g6QER1oOPARCM8x
7y/tN6r5PXPDbUSBUuHia6xz3lWvyTykmSz/vkdn3Twc1wNEAO20NRRey6Ikex61
6c/3ZCcoRQrxCmzHwHKwfVEOCWqJxs9ciHDEtu4Un5D6L2Y06AsygpxUk0FESONM
8bYXYUfiouweiBCdtr0xe/P6IJLsp9of3V6JQTMxaTqXwpcWBrmKikvUMfa8aBTJ
mMn+OA51yF0hFOy/Wer/uR78sQHlsnuOhTl7IN3k9uGtXyqydgO3+hloEbn1Ljo1
z0voGdwbf/tTSq+7xxZ4To6qolTXU/BE/U5yZiVBOvLycadkPyf4Vd3SMx6K77kj
A8aZDIbNVoEmD5TG1oCD71IkltGuXVsfEHNFq9OVSS/TmGG9BSe4Nm/TrcJ2mTrF
5gZU1BAp0k74ybyb/ULRGPe8Hf7YW6Poo+wd17RTYMqo18B3nXuVwVGGBS7wR+VV
W23m9KruXl4Xbw06qU3HDxgOS0ASz7WwkfYAdGX121BSpknkKjgolp0IcxPoCszh
fQCGuqXLJoHnY+5yXpk9hx33Ub6aOOFDPL9EMSvGwL3F22niArMsyKm0IbVIIlf6
Q5hh0tqJ0F5VcRBguSDd0CzamCw+y2NU2BLrYoe0PayZEpCNb0xqC11yCMwYr7nG
2/fJc5x+i9ajaJNgQxOC6wBIfPRY/rWm0MjZ2xDWb1Jvr4JSZ7G6mRof7JzKgVEa
E6fGCbavDGleMv03ITqSm9v+nxxwIk/a2UbpcuPHSskozWep+fLjQ0Jleun7OvaX
XhRRgMN4O4spX4ysPFJs2oxwpivt4fBFr1LPJwsB7kZo2cBelEDapkD78csE9Uo4
4cRuZqekyDhn/UAcQRZRZa2TIDvPLj6mWvo1WQ/665awi8mk0p0ousRZFs6g+M7D
2gjTmLHfS0jPmOdGfOmLS8r/bUy8fI1Ma3BcHW2ona7gTLQ5ukc9M7dBOhA9oHi5
AuqrPfwh1hogE831I4E6hgcCgHThpNheWG7BvAgk09iJElGrwAhg00dFOTBX7oMW
oYFwx2tlLL87Vd/fvpCcGjFNokvG/RT+7MUb4eGjoyGZxep5Lf8BViu7qZRl5c+T
P5HFzHJAbVjCry3uCAtrV8aCRpo85RNUJeXWQynBaIHdQgo+dvy5UiPWaR2/fHDN
4PPWDwJtQ9n3XDgEgbN2fV4cWCpKjCLefuR6a43XBnRFg1NndzFHY3AstSknULst
ci83yjR77hVbzIHWidRfk+kuORcAGsH100MBIEriUP7dyeH+dvcOT3Zo2NftZVPk
0129MDr6lFByes9jQUC0ysh2I828NxAvSGPtJi5htw+0UiMNNIBQnBY8HX6dD+Cq
E6I8dYW739h58hEKR3AiNewRhkfmNxscgS1bK2FW9jRT1ZYLfuivMY35ihozt+/E
mXwSVvGVbQYVJ+PW7k6Tql2LXTwTXXh7bvLTG5PPCPdcOOxv999L7/l6X9j7ago1
2/TPQ89jgezxT5rsWh7PtPXRfvtEKhiIJ/CPEB6+qeIYt+hatUoXUFPYziL9x1XC
erdcRnD23q4Dotj2a/rfxHHI3gg/rjUL8tN3CENlyJsBcSDg+b9hmXbUP6BxNz/M
YJ6HY6umpmtuel3oiCPd5PN5ChuHSoLjvEVQe35ugyUfNcYobXVh2e3/w0A22MhE
nr2hmcScq5RR09YwgWAve5uj496rxQyli+LCgL0MrLY2aOywSGDjsxfWegOASvmd
k1VnSpEsiFDsC4p4INq6lkHZYBl98XFdAMj3gAv/EG5wnXoa78V5X0MPu4SoK2KX
kIL0snqxGKe+og9jbULpjGQjFcReySpbe8Cy840eUjZSi6/B9YkE+vbJY9lVICO3
uHkiJfeZH/OPlmbMvkxVhVha61fUWYkUNyWrZBF+JvUuRhX3j8vQOPK3lYWv3A2/
mEU6olXx2rR8RgRncVxqoSGoKmd/swCSe2lzlABu33vxoj0RVsJNeRnpayBNPJqk
kFHzFIWXBna98WfyriMehqYb0y8S+BOhU6FGAd19sgZ+t3NFRQJGEEIrPgYUEFO2
FW92yry713IhlrGNHnw876FJs2Z2k75XC7umjE7GRmsV9ocHY1kGR9B5+9v+7eMs
P/qqXxMakt8aU3c4wqloR+ZvfUz8PC7SUrasxWsoN0B1Mfq6O0+bEI/aerYhCkwB
vPNAbFJS0RMa6iTyR/ORP5biwrsc7ku7U0mJdszgOq6BstkzK3mFezQDZzB/BI1a
uN1QFUZs6eTbzzuWAfPppyzwFGjYvsLsuQFquSTmeabnY5Yu8x5gDOHwFSeKIj0/
IfpH5OfNKwrWQ8XpiQOt/uBnXIPucjDywA+/HQadZ2aoenXo5vPjPfHSk4DMqEke
/miOO5Wmy3dkayWbVbnST3KvcH0eVFVN8vrJHA/TFuaLftGOH+oD+yWzr6O7+RZA
ZOEXcn20/odJ6zZ3iMQS367UzFLKuNl1sZf4AAMQdRm6lZpVKtI5dzaFw8TWKaWn
NO57v0ZRKIz8b+JoTSx/ywo/5MatgfrA9fQlauv2mJrwOExUgvE0r8UfC7N+h5V+
MD254nilKPrXl4tH1qbsvFv6a7+m7SKKTwPJ+HJWkPKDCjYpUVY3GmgFmEhsYND2
wpkp7N1q5wye6gVD5uXk0tlbsLCJ0xWCp2SMisIR9yk/quI7SYKO+YYqDdoWBPx2
x9cPi0Mj/IQSxEyr066YlZRO+qU/LySAYaZ2wMTtKdWyWp/ovzcUShXWmq/g45g/
unCB3Jl98rdVtRTHCaBBDQ0laV8fZzfWRynd8E8X/dItgWuKkQdyyUTsNrPnh03Z
K1MgBK5G349T7LgtmViBphnGrQnVIF7a8nNIw1EkruyM9Iag6goxLNp1VYSR/tSZ
ZKhBL/NZHOkmUt/M3eBWFvi2jBI50aDC4Scyp70s/J6mOelpupSqmMq0jh5JNCps
JgVlVIEva9Cj42rQevKwJRBY9RHApPKo+CtYBHUvFot13Qpz5KXt1Id/MeBubILG
XNc9pE9MtH7XAPdm+fM6bVbd8Z3rFwNhh1y4BM1KjYj+ngynZ7NucXp2idjlzYFJ
M69Ptyno2gefsO2FGLElYJLJciIHHMUreK0U11gT9FxcbSgRT0l7dYb1fQi1wU66
ozw7y95SkJwU7N9EIOf3alXN/ECRmDi4L7ulS7WeabTD6Ujh/HZ8hkLcacWXx6Ki
wDHqb4bPurlxLXzQwHXeaP5w1Gn0Qqgf4mprqhyGXYIPI7e4HSx7CjJHHV3+8lWb
n8VxVn98CfI0yYRPaDI50MYGqGXKCXOYlBZBx5O1Lhsx3SDmGQnHws3jZ7rPNclV
6NJLHX1lWQdZ+1bnl2SW8RU60SM/U3JmeFfqIPo2rvLgEkNI30JLUo6uMq+0fRHr
KZx/df+rUZMbEONOTZyo/IRI1ez/z17xIh8y6c9LmEfLki+0LVeBFOrCZO0ApCsi
U3yFE1dKQWVG8A/1yVggra9l8hOagyrM9zyW5JPY15OdPI3/S/eWKUt48QjUwvbz
lKHyHG+ZhUYG+4l2wDAsCO3QEgmB/8HjZPniiyQovw+DV9kxeUvGCJ0+yRNz8rTa
dk6X7QTfkVK1KXgoi19I3M+9OcT9WGWaXjaLFYODf/LQ8yL83Sex285dE93uAazd
lAUYqT0RelcUzJtJWkoZKJJKl69ti+kEKXiyXuAvE6HRVlReN6b8C478GHpBTUzh
9aH9lYGkbEZ2k8o4Z5uE/UUFw0iIT1QDWfmy+5PIu1S6KqfdY5tJGGswIPnp732E
BuJG3ENXofyea5jgYV47P/tRH+NIVdrtPI3aBGvEecVzEFcHIdmNhW8uelKGWg+h
wnS6Fj4qG57jINfG1AMncurEZna0S7rWUZm0oNdqF7CDyXjGMN79YFGy3cYZ/cbk
x+7Kqk+A8O+3LFTLhgUnaAZhA1BBnWJkuHIBxr1SPFdZgW768F7pnCySp7EEO4PO
4mTkjhLqzQDRRls35GegVzBhXvKtis5lwIOim5rTQaVCAhRodQXreeG0sTh+bIDu
aUnPsDS3ujULpL7rJPtQg1HBI4TTxmKlIrifZ/xY7qAbswGjl1RkZE6Zr8qXkM3p
CZ2KZSj12Kd+76IpPZSfIxnayX+7sjw6GmR7qladKx86uPmrVRwwetCO4z/SpZ3W
d/ZXJOWa4K9WCl5IKZsp+kJ7QwqgVhYb/X/iSy5J1En5Xo4Vuetg4VgFKYy3tABI
midD3zTffHqDWQPjLtpEsVQA2UMYtN2GWMbOCuT6Wh92snqdmxnRGPURkHyljD6b
Un4G9G87cLUe066vAitesr6HIrWfyPJAzz+pNbpnErG8lh5+DQSbmtxaFAGGZiyJ
JU+zvFRRlUY1JQ62utZUp5AF8AXjLPDqLdJqTkwZqQobSUIsh/dCRgQsv5JImazI
W9WT4zPzrJAe8H1VQXqQaULFzOlGBbbzjxKGIm8oS/H/PulfpsTfhHnFac8ZHqkE
43OM2SmCbZ1ZGb7cJVoBAhtIyHBXz2GEo+n52xCp2Y4Q0+mtNOSNgaOOJU7nGhsN
ZBFci70QtLLqsQ8vqpfYqKTyKoOnDzEJkVfrXoMQqNwVPUfLQi794/vqokzDUsrO
G/huBA1i+/FQo1xvBm9Pto8Y0bP0t67ApWsfAw3Ey4nJzWHYq2zA1kf7fkRtgVdD
4EiCNzB1n6AZUC3AxjJapJZh6cHiQw6W7l8nYxYIjLZLz/uTqGbj5O5YTMQpgvKS
CjQBrbRlB4ElLAydur8IQOQTdq7LkfDImSPjpN8EyJoxOnYMFzeu4CyvwpM1VWfa
1x3cvU3la9BV+io83fYvpfCAMBYJ7XPC4IVD9IVgMfTtCng//QGVvsRI0mv24QyQ
VbvlC9oIssJIhfwyP3+Sz1lqQQLWNtF0IChXRFYSsABeD+bgjr6MUAGyJLixOeuU
FXb/6VAhCuR5s0n5hAxtYHK2Ovq/t5Ej6A8AjoDBsfoE0mv2nES+zC6NWZ6pQpfa
hO7DIzL/eDyVE6GZSUix2tyeXBID6LIzTqh3Qkjc56rISaRJhpoZLhCSAU3qHaXC
NVZjz7dcyhrX5KdXK/voB1vECDEkzNced8/Olgi7Qu9n8oK4o7R2K7NhTVyQQSWT
B663PJpVSGMhhghtur3nUZl7JDP8J/EOicVdsnIgvHFObbQ4q9EOtdbg5Ohj4Lqe
eAr43z0eQVDMMrK8Q6Y6LtqStS5daoRLLanWXyw9IYYYYRBQr7fGtMeE+1ob6L6G
etcSu+ZwhgSQpDcYOKHdJOT98uW6eKSzCUjVjYbS6aUlfdqrGrfDh6QUpy9Qj8oH
cb6iC/4Xes00Ihemb84NRkdue7N7cbNIT8Qmv2piI2wI6XSGsGI9zFF5VSmU9eDP
WLlm17ZK71xJLSrrqEmedbFtigBCpXgF+N/mqa8cSn+guv4UVobcXaYu6nrRZKEB
1oJ/h9n8F1h1cLrEspV9HDDOS+x8DYaY13kFO/ObJVOnrmyFYYQXLOY1TNpPckc2
j2ynSJhUkDGScOv3rMqXvtF/fGor1xuvY2pfdgjRIx2VGYJ2O5OltQygHWqRlQDS
Xv+dzB5Edf6V6orCpB9JMdVgiKnLqGOCl1s08m7q0VVxgpiXbmRmn5dNHtPMAgDw
rXKS+H/YDl4XPbOY7TSrfLVt7yqokePlwcs2l4Y4b2WGeSOZMBlUqg92SKpiG9ky
x9luwWkfHK4M5Q0gr/kAj54Bf6uN3w7fSImYkmJuRAlkG7pSWXPhK3NHPGOgP5ah
SpqAZR2DVMY/0bpM5gCineOD0++vJYU9lisJiGbrKUEHQL/mVfBOcUviDsBLEHpk
MMyYSP8YgEZck3KTft46IhBEKzyJOvGRePqCpttxXu1U814bIes4zYnlIPGyR1Q/
+EquVSe25yACd4cEkm3JKwEgp8Tg0ZjTqMJEo1C9nALEwYTo+C1ubswig9p+z1Xc
AgPJnkXNzq404in4l4AyiVdMOnxr6Ti7DzcmV2t5I5WbCXHXLPR6VLY79yde+JlH
gGJ9Ml1ErhMWzDHFN+LNCAwuKumYEct4O3yJSCjKYhwV+SfwuI8vMCYLtoPm+aac
0a1WdZFGg6K8r+hIV06osgvo5HtfQbxj/rrKRc1B6ysCa3O/eAiWVXbNL/UU0lvR
Wt4ixGPFJ0qj7HZC3BYH4qI9viDAjvg0kCAGyTG2tgF3G9/A67yeq1p4JsUgwCpY
1FOD5N7xa+MxizZOvbqc9sU7BAnZZjLZp+/72dO3y4w8NraCxPG7AoAisRvdRLVN
lCk8oJ+m9NkT9oIeXj4AQxgcOUbbM18SVH95krMO6rj57RNJTRG8T/zVBI6oVAUm
9/fjtbJ0NwspZ5LpTJcY0BF9+EpdA8Pg5QvMP7S8Eimb+rugMdqA1ozikf+QJdO7
NzQ2rvJrOdOXPF3eKBAk5BfKfVT8LcyKhw/OjYBAT3xTEcC6Cpv4chBvnQz4S45v
IxMmp8ZXVgVEEnteJaDFSKTqat+TbXlOt7O7rA/3TzJFcnPNuaAfVp9UKZUVNa72
bLJIMC4bQIhhjyRYLE5VjRHIinoW6UXshxqR+DVndRcId74dylvTSku1O+ws7uOj
MAmMz5ymOsoAwBVM77CfdJXXXYVt9TaabaVeajGbIK90ckSh123Nnn2wR+kOChwG
js2Xe08Nqm1S8Jj9NgPACDl9RVF84Zcd2zHMuCHp5V4mI68ZYUROWtYKbBA7I4GQ
QsbT35hxkggLXMwuG+ZWSFac0tQbhJWTHGC2jtQlLyDTqyr4I5E45pxyw8RsiCoG
dmeT2LxUk6LdGD9YayA02QkaZ6potfskNTdkWEKOnhl/MhMCB7VSMfWFYmiO4Zmt
e+sxobhy23EK4+y1PiUo/JrV1DflWXqiARx2BLHrxKpDbKQtZx5d9vpPOSq7dl8t
adV7K0jyd1a2VSVey8xlsUfXgHZErViGs6lVD+jtwiRlhvoBOowbZSuljA3wbIVr
sRt6BlIXvaFPX9pUF7vBo5PSI5LJ3woX7rRU87nor+TQD89wUMG1tuE54YWTShm7
hzbOD3eiwpCIy+xW42vq4Ncy7Jw0mzymWknraRDQNrRfs7KUtAc51RMOHiFEWPO/
vSrVgsPU0qdfjx9qUqghyXiaHZEQ1go2d5R7YlAqK7u+9BCtLFTM/mLBxoD2x+z+
LYVa4Q6ZQsOQi6xdh+IvGefIj1PUAldsdeY14gWfDQriupp8WreIFdDBiWEGApxS
fVhdDIpGF312a0cc8YYwU9qQTn6OCjtOTXlDwrT5k8af/o3qiAUeySh7YD2kfdkt
pJkEkDRbeagGvi1/peQ5Od8Wv0JQkpI0yo3cctO0byqTcNwdspHR/HVX++H2UKKk
rDWilbhL+o5GRAJ1l+ctm2w8GKUwpBV7YgDOCbFou7In7FPWtblrNuYi6NdfryId
XxxDTefLj1kBiolbNpKNa6DJVJzRbIbCa4D50ezOff0ViiHBX5OQM9s6yuDXMHbp
f66BmcvifY62/9q0asn/BWFPyaweYmy4kI6pPfMGsDhuGErdd7gPQgzMObo15Flv
Ej7Qk8l05Rm7msDa5RUAqpkiLwG4mYxxeyLZUu4eqAwFd+PtdUfOfulGWz8igMYo
SNz/Bbajv8iuid9ZNc/W2eztGBpAZUaBqPNeJ8gGTGKwQB35ZMDWqmOfO4ImD8Ga
igy0E9OgZUV7rKCvgGnY7OH3bxccWEMNK5bnqiqy1obCYwy2JagbqhNhu9LstNt0
nrObALNR1pIkRQA/vfHc5dEiG8C0WXUfS6Rgkj7W4pycQRZawcBuoYmbklTc/Y8K
yJssdvSgPozZEeaOKns1jZ6mj5/EZgezOU3Z8982BFsYmFZilkQqqZkOSSiSmnZX
EUnkzJIsYx57Cmu/IzJr6wDPUwfkrv0cJMEldY98F9sXIyBpJS9mE8C8rISi5TWV
V2TTt4GTl00/Brdn8mjqWJJOHcVBuU0QPt3sz5IhwnSJy7Yff20GG4qco8rO+8Lg
KgO9oR0uaXWidq45vTli9pRD551mpNzN88eHWShzdV4Pmy9/qIXT9svcvrJTnfyn
o59nJAOzRZFDYtiPYiuQDSkuijc2o7yav3DHmWmbrNIur6VcE+K1Txng8j7Iqr2B
Y+WRLcpsjiwCNzbj5Kpc1tEJzgKsWg5O43CfFv1xQ6d3CXvWWy/UGeSKQ4LOrKrI
fr4yiJgY8r0Bht4dJkaVhqZ5LeuEuaQzci0e/geVJ4tOcV2sOEI9vNnhvwPdX0GN
gpyzsbqDenf+Z74XQuLjzCTnEe9o8Mee/VTCC/GlD4308J7wWP8ZXSucJR0X8T9U
JE1R8WAZC8KDC0hnTs/vbf4ANzfRzZuQvq2fXDj9cbWZWMc6W4GqsB1RDEcgzkxU
zse42iPdBorfEwH3zDgcPVr5BfLJgdtVJjYHCgfPKi0CfP9Qov0cSlnSn19jPJ/2
DgM6arlDfZROToqSfl3U2c4Iyl4DYuWppWCb9FmlcMMH6yf1ChEhVBJo5ivAyTR5
qqBfxf8gyJgtva+kP5F4dNLd4A2CMZjRk7p+8S8TYoY9P6IwVFF82s/aKOExlQFS
aj3qoKhAsii02cIPHsqP5kx9Bx5i+Xnreade+lm4PFHBAbeUxS2hqDxuQgEL/Jfm
jELmEngnpbeSmtoYItAsnh7otwM3KaxMafT9wYPaVgqtHA/aiEy1Ev/0/iSP7p8q
fQrQjEq2/tr4CHrplJcJZ+zQIaI05SyzEgPQsPYlN2lH/8+rXI/wgNHwQBnJBumK
cZtGhvEOj8LDzkrTesDNiQT662EtsOoKboQxv/sY7k39gFYWh+GUDVF3FwPwwS5U
yzgm4FE9y2TdhCWK+efeQsk31rd6SFUkf4I0fftB1E7bOKgiVJ4w+IE01deeLECH
7wVSBtnTGnz18rCJZEw8qqlW0uzojfzY1NvK2I6iy8nN1e3cPlTcKaQHnOHde21w
9u/fc2J7p0Sb28tA9vyagXR0QW+VCnXnZYChG1fpuIaZgpLP5mzE7oloaPv9osla
G02sDyrlHXPi64qT5/noXnzY3YKmUpVUdWPlmEcdZtv1r41F92p45eUk0G9lrmwv
FKhXFfwH2K6aDkavpasQeRC9tcVpy1PLv0bakeWpALoerJXsJnE9dkdnp+3Wy4TU
MvReMgRAc5HSIomjkRSeDahOfGtvFPP1V6F/JAT7Yb7s33Wrta3kWtEvoKZR892X
JSZrzi61SoaIZNpyDhmZOL7tQukAkz9VPqEbuZAR9O18OxWicXy6unfC01Kdt8hh
CJbfDsNCcYXcHevR4dLNIxbMUKvYY2coiFjsM+jtX0jKkHLg/rj3ZQwohnxaUEfA
YipbqtwOR9ZniDIPYFcZRDgpYYK4uL0JU5foH8heki6RO53RXnjQpewJ1kGbJ5dZ
gd3ur3Lnbrwyu+65T0w7U70F/oRhF1pITsHw+wXv7O2zPPsPWP9LjjeqsjBYiEOP
B3CcY17lb8NP5ihhCHk2GGypKcHJIh3Pc+1dbvvdi1uUbUXyVvGJrmn+z1urLCZH
DQd9MFbMasZNmQ2o83L/SS4OlqK155BrVuiXHYB+winR34dh/9PvmLmEYs2tvz6G
KQUE9VGvg6k2t8CdR1C8ozJSaWUkYnc0faFm4IW2ZpdkY6IiM+AsrOMwrv9vISP2
jytuJCzvz342fHyoCFvZUAglegAGdxX6ML/7H2xFr3ufjTdSWZT8ArDKJo8zcQcI
IFHecG9R7cyxDKMuvF+IOP9QeOqDshcGhBuX4B8MlhIEE/AVWmX70pO9ju/+iBl7
Q7gr7jq0KA7i1y+Jg6PjRtWWiI/VU8VhJOkcPtE2WnJuZiSkwjQNB2z78ZTcgUn0
s8wdybty+OaWWk4fTcml/QPadAcSTWaOaTqc0RFWlxhhpvOJC8b4aNE80CI1u5Bc
YAyLIWD5f1Z1VElE6ISqH7Doef4qgapmcG/ZFEU3CfD11hC16sqfdsb1e5D3vuT3
XlJqTXzrqdjt4QCqAOBns849S9ssfqdHpEQzu6sAeVHAVMSaXkLTrZ6ihC/I2R74
3v8lIFt6jXKrhd8EAx0N/+YKjfQ/m205Itso83P+guCd6UiSoA/rkcK03qt7EF2J
E5ZwzrVJGkOvWWboGYBXy0vSPqJXntxCTTgjARvX53fMrPxQYNAHsUImaS7h8FWp
m6BNknxCiMBgWa6QxSy+S6++4wsjIzm11YL9B2krRTQQHVVZYTdXcn3xb+gat016
N3bUG5+ZBLUfwCeCes6XzmsWBSLIT7ZvdeqLokwIFkygyLNAVxYWigMCxG4UDX6v
FNYTDQE6zaFAZbUIl63/dWFM7il4aoiZrcBslmsEPzPeVIr1WU+jCcqyQNKJEYI0
zMN+P1vuj3QyBhqqUkrERlgQxHTPqLFZ6nol8WsC04TKcDmMJ4UFd72fpLNZaTwh
npiXqQipObtK1WvaM+1+QHvm8JcHp94iXHufY+jvnD7L2c6NVz6PlvLvS+44TyRo
tdn/zKqHjXSVu8KRZxHZLZKfrdA0qLjNlKAkvcgsJ9JwPvM+RGoVJ4OUC76JjdTj
zR9JjAQjZfpx8NHnyGvvTz5oJyErnj2+PIkAOYwtV8rIODM17gfnOoErejxHP8tH
n54fZSqsuv1dxJYmjYTQ9druqzDlNUyWY/aQkZc7Kl8msBLUR90ES+iVFqF4pOyc
lzKbZYRXliUy1Gs08tS0lRWGngmqc3OGUoNmKx4rPRWAEt5hOvkrq1HjdtvGuPNN
g1Wkyds/n3YSj+tleV9MKDqbC2t91KoUits3omrjwwwe8A4kSxRAi7V6NvWI6wz/
yrZmSpDae1YxQe+YqwL2iqrzpfi6S3f8i6q/yaikoL034fHlLr8iSfrceJMkoG/U
dfaNgxrF/NY7mRlL7vg569WDCMexIjzY60EPVMhoIF5nmtqe9TC22CUj9vGhvGy6
PCkJC5H7v9Cf9vUYmfgV2RlYS12wtOE5fb/zxicVRwRpRwhfcgxWKAV54kGWaA/3
5K2IIAbhTzmCFhsLvPuwulMF3WFflGphv9EKyvkZ4xWjgUehMZ+a5+VMGPqAysEW
mgTLQD3JgmrebDc9nRMl5lXbNfaN37Uin9lqzkQg+oF7XIUOLGbNA888Ufpq4fyW
cN/BvKczcWas9XEPYrnCuXdb27WBsxJ5R3r8sddqqL1AhBjWC2JoEu86Fpmrxj3H
2SYmG9sC+BrVmUPuifWmzOgYoExwWfuOwgGLKqqDKTNQMeocdfUHkaWCYXUokF8Z
QXPaQnG7iMjPZjNXILCw580rGt/u7pBCb8wiRnB2DYMlyGhjRw6Qs8aWim4A0+f7
77eiLZoxUUmwuTq0jwU6eFrmChM7aIt8OGr0EPwcsU7kb3a2dw3W3s7Gf2zj4k1r
65igMRFP8VC0f+bdJimk3hFP2wkq5AhfeZ0A/3H8FlDxYgxyyZJUBlHhpoXr9eY6
IBP/UlDDdKisDFOBVetkjJnyKfyHYYsxgkUjT8b6gMyP+qLf8Td8kHhfC1udBQju
gJr3S7CKR5dvcuqBiuWyl0XCmoCRABO2iA8B/ipVvc4EO7hBtrdY3l0FNpF4rfSJ
UwsHDpMW+OkJXRY3DYpfOkYkDEoEV61bOaKdXfYbsL6zRGx8Rz9OXLrQoAJ2815V
ADjbesuVFD+fyBTqqWoKcXKWccFZKKWJiSLwe7CvNsN85Tn2Ub72z2gd5V7Uk5Sm
5i+5x96mKLthtKAujUdbMHi9bG1DfOGRmVAZA+s1EwXju0MWIkIQDgt4vDkm6dRh
Xl2CvT6/l31GotTwwt7+tBNui+pzVsYWbUfxJm2at2H/tgoax+7DMTrxYmUUaNIV
xuYzHKCOutEaw+lb9bx75FTmfwGAFeqCv63rLjyItq/NiSY6n/LAGP1J3aO9hM5K
sXWx1HzOOPRsk9HDK+cAB1ASoFe5N/fYC1za/9/zOEM9fWIXL+6v657u741BeeZr
t8fJcPy5siEa46ofRaj0EFIJP2phHhXIZcujmRbmIK18RRl6C2BMqGMwcFmk9FAb
h5p0KHBLG2daDqsrvm6YeVj0ipAMpH8p6VBpgntaJuufpydqAmeNCnrYo5eCcUoc
oQO/8un90W0HeKCtk70F6L9kj2RSxUuqvgey9o4rKbQ8mpNxR86H/xz8MAWkF01Q
qNPYk9lq3KI8qZdhgMzfzd361IVG9ZRfOY8C16rPa0KDl9JcJNtgo8gDm4nHtb5m
mYp7KPU4mOY69N4zJkwxrN/aI/Sr69jUQFFzc1Zg7+5DLTilCSWnmaCfzXWUiG7l
PvVqJbN5t5xwVh7ponHW+TCAQn3RZwp/8msJiKimk1N7tBCoGFkzVlwFh1QUNtym
ptep2xzKCKoDDl7RD9y81k4i1evmFSTX1QMsjR3IkKw/F0ChfRIcxrnzAWX5wroe
ChE0nMRBMUViUCKBZbI1ihKaL4f2gXY8TPoDcc7mKwnvk0MAjyMDY2639k0HLmfI
4kYiriyGOltFor44UpdwvSuaj7JruhRn3RjoyWTV7mT2HnOu/5CzRfiefMBYD8BI
5SYW+msXdvMzSEVynuIp2uQE1DJwWO3F3mvsPeRwianjozTapULRJVNeKdnt7zRg
yPNEUVw5rANFWFQYLqgRS7OMCYK7gNqlUE73mFdDWtAqxxLTnZD+pdM7EDOLFEAT
xQzM0Vn5yX+SkJADMbO7l+rUceSE3+dtu/+9LzoqZqh/Nw3BZsIS3CiJWdzj0Fp1
81rqVI70eCQsPUppORLIfTvcuheK6DHMNXJ0R4BsShGbvQhvzh3H+pfb7i2sH7UA
+ToF4Cw0sXi+bTt41bvXd5+IXCOmJ4u2gWaVKa620m9R97JHS42UGLSH/xP1TCSv
yS8JdUzvMRiNtQk2dZ3T5zQU6aB3dw+fFgqRwGIJr0Qkmjzovq/eMigXZC5QXMXX
U62LBGGIjbHC1RqyBWJih5hsxSMWVHvt682VLtJCCxhuYi5QhPtTvNKL2VtG3eLI
cgmKppYeyDet1i4SykqPNzSVJHUHcQqILGA4e46vTgP1GGMziJa57fVLqB09nQu7
oYdGDGTVQnaY/k2P/HBLnxEC7h12YOVqygvHnq+J5QWHb3ynZHyuN5RJ5XcNu2CL
lNrasH5btSc3qe98S8Hr1pUAxfbnwtokq/ZXUMtDeNDfzGfcDArGsI7bs8NJ8eeS
QGrUEdp1a0r3h3tDirsFklmfLbX1M5OCKEXOyF3QDyiucy4WEXpv6ljr0ZWOWcKK
F2RGElCppCJReV1TQqkJKh7q8npOqbUOjwmNAOrSiVEUE3qiO+L5Ow/PXuAQGe5M
hGoG3FL72Zq4pMalkfeG1ahFbE+evZiOkqtLkegHugs0LqiyRJTkgc5sqKqb8mgZ
JfRuL5aRXOVRpEvsQk1ew0bGKDd0XGwWB+31hp+zFmgcmZnLFn4b8HZSo8HnmYaL
AB+QZH7PSlHjs1w8kkwhpi32RSXoWEg/alxhqDH0wzZ+3ofkY34GYKXUy/3vPGS/
8gtMruRNwnoiP+wSOrw/Vlfizukc/mpu/o7pobB5TVaRrPvcFRECLvBrRY71LLbR
kBcvZcdhVKKgQGjJ+lImrSoeIOdzb/NCFG1hTsS6rq1F0nAsDyyXuHIjF2PqoVEY
N50en6EperngzbCOajmQPviJs+IDPvBlLQPvqNnHTV2S3wGDB+Ys7aPpa0O0R/TW
RrMlc76m4TtgRU4Zf8A4lWMgu5zNIDEbpLbivbj8RE4hq7SU8aiQeJT4qgOOZ8It
R0GrRRJPg3enFA+UWCnbDVGafBOyo2TID0O3zwNqmWGFVOIjjYyqbQQuggVnZMa0
bD7IvpbasahCx7d4ol6coUJqnDNAI4bOJyxYQp6bNe3qtb8AxstU7KdAGySaEWQn
MrEms7qaJbNWl3sekb52z5qWX4/wC4nUUz77w2LXeQSHCNo7w3lrAM8eBjmUrBCY
VPvqWY2vq+D4ZceTloFuADXI4MoZ7t7HCX+nLglruguuyZDGUj0rRjq7rtwHJoK+
Q3XRKdOjuNg2yK5MJQ4S/ypEmJKWgIPcO1kxux85grsapK8Ln1t7LOgl4mEs1Q50
Clv146WvLpTHA5IN589y+ikhu8xEiS+ZHRkVFEeB2RgeA3tMDxP4AKo6Bj6a9gBc
GeTsDj66onGgNX8nBw2b02236sDlDBa8yfkLhFq4kfBPosNhsFyZr0EZfnp+q4aM
Q4RkI0+goukyCdirESyGm3oKYczv4f9LtDUuoT8FuN//ORSXSPfAsc+PtwrhS3+h
/+MYS8S6MFMG9GXM/L5Uc/XOYH/JNNSAyNps8yIh53OMfdp/haV+iH+Yy/i3UI3Z
LMMGPssVE+2H6tWEKfyOcohFaSUSU4WvShGo6/TKAakbUcx+2ygBF7wWDKbyTSQk
Q9o/3xsxk11qoQ5ADsb6+YMdsGaJMtgVyknTp0yB3axw/93mQkoY1BbbzYR/OorX
Hq5gJTzZEAImy+cDt5feQ1uTAUOxplZknGYIgPSyvB1DDSenzEVU4j2iWrVDCC+F
62FbtF92G/QGp4vubS01l84pVbRUr629E6vudBBn30nlp04Mf717tFjgD33L98ER
MMiaah5GmW2mUANcfooZcf9Iiwl00BBAJwPq8o1E5NglqK4nGlzvOYuVZuYCAK20
aLQmaj60F8uinNB4DpDGUOwQSYCLiXUHX2TegPLSsjXtgNOU+++F7Uk4PSsq0l6G
f/hRObWRSMJ/WFaaiG0RUcKwAGF41lL792VI2UtBFX5cDaotg0GlkE/4D5EUYmRv
8hgBu7STKNyTS346bJCtkXERbp9KS3Y2/fEPRXijYW+PTT/aNp8XCDLcKHuFaYiR
ug6M3xvzNZRYLZWdY5EzGX3d5yzbTjjgNa6fgD3BQGcpnK5fM+ZMihC0sVz3j0Xe
XtwmcYjd9mXP1th/aoTxlGgxjjo/VWFl2LfPy0fk/M1fFebSqESAQXrrV7nBZEFC
IwXV/tIaAzANKYpLTGBjMRAhcN+ohiXYRCvR53IMorQ78GyJbdLjSv2uv4S3+7LR
3LO/lczwaPjTfQzvQZPUJCm3sE4oBDjRcn/xQtslHPDnIxS3attHgFyuyeHcGjwh
po4HovIkLRDnXFN38zqRoc3Au84oSuUYDYmnRuzmRxuQR+gaTWN3Radn5Cnswoge
DmGzKTlS+9NUPdRZHgipfx7cyypUIc6tUDTXppB7MLE5wDRMUQXGiMP3tsQfRxSc
`pragma protect end_protected
