// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:32 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VrVHjVbKp6BOqr56ihJtGS9LLVAP8NkShugxwak7FqGy+1cfmDrFe7HWXPNJ3gKT
1VElShBCH29PTbCS2BZf5KtiAdRibKfcYkwvh5qxlq3cTpgKPV5zHM0zlQV41Ove
DRrGsV7sbCJ1Hb52tJ+nZznXVAQFi2aJNW/F6D5otS0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5664)
wsK3CTD//seG+d1mpet5XsGoi4A7pDXGBAYIiKCwXDkTk2L4K4hZXUVzZ/IXVkl2
TMXYZm2Ogz8ixnA+rc5F3Ufr5rXPiz4VFyybxzQGrE2lWDnARTJ0AQHc2py76qpD
ES6LEzAJoP+MwQWhiWinKBVoRgJrXy7cHvivT/Glsq4N6e/5W+dDmBJh9jLZO4H1
17VUbJvzfeQlCZqdBqtbn6knpz3K/42QNDwXMyLfM0V+HSvuFmoubuiHNWzZGamw
xJ1hCmVG5Mo+gULouHi1OPd5yWMq2QhT+0+xdJdgepyJJVsVpZfwC/y3b87XULTC
ktHmDdykeQeAMkXvsf+YPlAoq1DzNkWIsSkkEhMYtlJg5Ap0ldjsIgFzR8sMspub
98aQbYSULKhl5zlGbwloQT23CWUSEERXwMJQnOx58u+Ic+8uX58pN/+KZiKAI766
KuFKaWUebT9/zodRXfZXcJJVV+e9r3HUVQxq9gJFFIdXE9vvHuDxNeL9sawK1u1I
bK0BwYCdZCtWC+ypqK6c48E/xhvR0AUl8oAh5w/7x68QqyeB2Vjut6qNfAsiR7QD
XvUupANrGDKCfTAST9QOWQ2h+aXPWYP7Rhtcwt901f7/Bd4ZvZhulB/BX53m5CMb
/JoYFfEQfg7Hd8LKHpR0nv++cYXHKP/ROWyQB/HI9lwNyUVIvBjFqewKd4IMv0vk
r+sYnfF7db1tLe6Q8SVOmYi+KBgGmm4/Jw2mPK7fsFyhCmmrTet+0YcyibvtWufe
jdTm2IRB7sVfX8+4Hdk9jhXNjkcF9FeXC4RZYFw1LoZ0ATfmaDto7eBtaNjbBjyP
qYxp7QDqHcIZ+O3pglzks01dcmVanBIqdA/hsbrbTyLpR//KzCS35P8P8lIdJiNO
NiByVPAEhTvmZN/+poT38uQGBQLYrVAsQjpdsFuXeDMkHFSIYdf0FLV5GRYRoBGt
8/ayZQiTbZf/CRxygWxlcLCY+ivsL1864alj2eZVFRx6k1fQ/ove0yi3NHFVYs2r
hdJjc8e56WWtGm/O66OpMzL5vwtPg69qk1yGKSkug6GGsrAYrPEICYkfci8Y5emo
ZmzT1kquNHvbPQXkdU+JSljS+vgjuqqwQxD6O+cGaQBDHv9H0IEyNMF3S7I4P530
kgKmnZjNsbUBF+/aC6pF01rP+93RXTo6iEUo0DuQ1ypmQV579jv7GJVw0CUu+xoI
nOAbY/CIvec8UV5xNFnHnIX4/1AJkI86E2VR8FVOg/3BxtGBK5lyaAS3RxB+BqwZ
Dylpi+UhzcCq2fgIk6+W6W4Y7oZm5A99NsC3HQOsVrY+ynL9vbYbLrcvphJmV4dL
3mEgpf0ZLMt5SetjSC6+ZgvI/h4COFOT6V6eBYYjgYxXXodJLIxjOxsZumcx/05x
WApBmQKZPRZZCJOQBf/QILdiNAsW7VqgHVNmYb/jPmCJWkaH5WRJZiKK5lwQa9sz
K3XEdUaVqdauKMsoXZDUyRTYhvoHtDq/Gvr0EJG6pwx7pQBhhGVTWLN+iqTHia8H
YnqmV59vEyoLDSwsBP2PhdhCVFxr03DQa4PeXjFNMgdsyfdlk0OVAZYWgu7iNVtX
iYIvheBPVNhgcpgeU+06A9Rzx069fvmh1Go79b6eRZnY6A0MlgK7JyGe7O7r4KLy
FN6qlvD9EcoYiIEi/Z4NBgzxowd8W65+Ecd4jEkq+UrgV9wZlbWcA6zloO6tTP9r
jNHSxnRpUBA64Qwpgblg8dfzptUDP8ieDM+slwH6XMyJHhqBd/geKgFJATMEdn3u
vdUjAtwmk37s44YtPA7MvjDM4ztlrdr4eupdy0QEwLH9crf2iXkbyMhDdEo8Ma50
ryPzGTEcPPx5QTPoh3nU8liU/3TeW2mjTd+XWg8o+eXxZ8Uj5zlrxr15qBQTntxI
XJGvbnum2y9wRyuxiPxjFBM693iy+5YjGxvDohlwNniJkZnT9ZWmB9Kq3sqo+4BX
tQB0heJLShASVxcEQ0lC1Qf5vW9cTkXd+LGgXoz7Mhi7DtNT42dBOTpqcNoUXqbI
Dyo5kmnnWXSFR12PnR0UG9B5wsHa9wYlTizJA1qvpdkcftunYU90mEges4NqrjGx
6B0QSm4G+zzJ51tqMZReiDW0NbqpIn3kE93EpBAn1OIVT/bljbKC5G6rkCCq/iZS
elLN6sNeJlXBxUl7eKb3mM00z2Ol+yFYHNHkg0a0EPiGac7EXy5oB/1c9KS5bW5X
qNT0aaaXSm/mwjYyxQmoR2tkjFiqgWNhMKXrUyfyZ4EQU+qMk1J1YaZKbg2SWPkJ
xn/6ODS8eb3ayhEmjbLkXSRT1UQBRY1inuKOVeXGboMBe1zO9aXKzqEaqdYYo+3F
J7PnDKm4MlVYHD+3Z+d3cvWQXHftpDVsec15KWkWfARksJitJQg/KTGECE3jBk1x
Zz1Y8Z4b0V3g/mcRFWQBT/DcpDScYCL9LqOTNBXxzxfJ0V8aQE4NHHWsOSS0rHje
9ylygYxqLwYG2Bmt77ucdUjmrGzZctBmp/2VIcbGXAW6E/vKMZUmtRX+ejSfFJgF
BO3nkPeFHSOLlrGEaeHES1MP/fYVu9pCTdFiZS5iSxwdu+Qayeiw3LNxvfWlC+FE
0Be0MufUimeqYjKXkaP+3Tatm3KHwd3K7T3vH+m9cJLG1NJ8T9Id2HtMWnYtRJnj
H1YtMme9+6ZL4gRv0U/+i+mVYUZeMnjriOSoe7PEKw+8HfX6K196ou01cFNxTYOc
vOickNQZbEeBahVsUv4ax3n4pK35HBVHHVJarSFpcBJDVytAdt0tlxT6q+MiaRSu
bJLrSK2qkc1QKJOmx86HBk5GnjcSdm2ovvvfXNuLayDeyuFiYkqK+r+BJpdB9Yh+
/8fBPSYs1vZn2Yby+pLX4eW+W0zGZD/6QKBrv203uceOOwkKmlxFYE/Ura+1ADSL
DDjZHl9vR//TGVqdMZMnh++76zeQtEe226eV+4vNn/xeluPQxv9gcWyYgXBKrd0m
Xkau6XRVIJr792WRTgRReDIPNRalpgAypuyRDB5bH+skZeKJ8Als4MRwOSnclfIV
wbsB5fDLX2rHoLw8tp6EZZDaJ6fZ2FCqR4v7Png6RYHD6gCFtmZfxKqPy91wDSQH
WRYwKXZw3ZTyDqpUN/TWtP5vnbwQDkCrLXpPE1xnZNTkHch5hZYLc8xbNypjqP1U
cwrxeHHY7SN70TTN8tNaWqcuqReRSGIWBy51LbUgl2au8VwNDvCUsfuliiWSyB+Z
m4+rS8KRDa73Pyc0CbAHBUfdACnS0YpUvjTabeAXs3KC/et4v8kd1+4KirQpSsL2
9rAEzEF9hPODHpL765cQoTsiPZtd72NR1FxN7WCVp2kBkChms/kZ6b7M9vHX5q0x
eAoXt0s1g6YeRMfhigSB0lPHM7jQ49KPdSrjg0ASIgwQDON6tXdAiF7xGFvoPeYw
8qG+/5PL3guxsY20wkAdNF0YgsXMPqxB1IS/AOY0/dxAf4bfxxisjHe7fbcZzo4r
VXB3gDuBLmgStuKjz44WUu0MtpXfCy6+SpuK3dsY22nJ/MnlpOMoeqNHnvRVT6Ds
n+hoEwO8hkywB604wTewR7CM7Dsy8bzqGQrecNNrPt2J0HZQRdRadupeqtR6PGqt
Hi03P9DKhT1i785ya+zOK9SzBAq5Wpzsq+ZU/uYtflQiyj0TPTAUTktCR/bzyKL4
ypr1CnLIXfozFwdOi7+5usuD1Op8HmkTpBQTV4krDXM57dCDJGu6CgAUkLemNkb2
8aBKDw3fTq+ZLYuLxT1cPsi4CwyBYUlL8upZxpgJiAT+Rmy4UhvVYKhNHxhGCSh2
6p/Vz51EdeoTP7VHg4O5iximavI0Um6UotNxspCw0a6zXx2GNAk+HvD9ncPM8Ng7
B8poDc10LEDtI0QdqGtoPwMVKkDpAX65bzMzxy1DBCnazNEPLXanvcmap6vrvt8v
dRU3HOwdsvCSaOSI2k4BzBCPdNQCR1Cxkopfcqiz6jAzH4ldpfRyyyaRqnjpQbqY
5ByJ2DBpbXVd6cTOjtbZbm1vCTy1Ew/uoN3DxTKVdqTw+mdhuv9jeubJTaMOzG7V
71FKLVO7sCsogVcdTVzD+ru3FuZL9HwwTl6/YaqPpZdVnTks/BeKCv89wa0kdIti
+rHAK2wBUgNWd6OoQKX2Fu5DZAzQoWQBBGOX812kyBEkFAPcrgpLwZ9cvV8RlsFt
TTo4pFiCePm41aBBTZciRbWJWDErmSmmM8dZBqs8wyBBFxWhLsFJLRK7xRoryaZ6
79wJQorIewsFeDaIRCQKPycJrOrw64+Tc+m5ikVTTrRfGLt7KzPk9VHvZUFTu3C/
f+JAARhOrwKjSbMlhZaPyF/bo6uP3VoPjE7KZhlBLFvY7gvQBVqpAWEIi2a7zCoX
rsXNP2gcA7JwPEaqNzw8viUazM/f2o7ZrTMzzLO2jc3MxsSqXrH5qL6zyXG/Dap3
AtVwPMmwIZbosialLuDl+Jb7KevSPqgWQSLAwU23+eo9g8TCwVplolMLLwzAKbSG
Q7JvrAliCjQapqIPSBegoJBN5RNzcx82y7SlA+a4URRq+flklOhd82LjKFbCiNmm
SWV2bX13N+fshds3DgmAeYNjLOHEruD01tmoZbCk+4hkmi+aORl3T13d+OBZxypF
L7ZR5ciJTY0nlu9ckUgizuDANCCznUZnWSdN8fHPVow7WeOQgm1affhkLPUjBS0l
mPJl8Q5VHuxTha1XZgj76kXD0GpLcrmHrj2jWVqpirMCm4dwbBAEv2coPfRTOvlV
ziFmrz0QShbJB1h7/VcPQHJ4clmQT/B8X8PUDOusYJ6ngIj2FjBe4JbJ2tbx+C4j
a7Az9N5Oz6P9+dZ/yX/DW7+TZ+ocAgUAx4pkOMyJ3FbBcPtf5sLE1unrnatHQzb6
X6BPrPbFpEagVrZnw8qisNuuR/DZp+WU0zzRQGes5LfBGyE+VCLA4shOJwp/meKq
8w1UlmDGn0jJxS7KomDbSaLzzc+4zlUvrMb8YXhKgMo2Dj6o8uTMiCcwygixqwtQ
OTWv4knN1aRMKlh/qEoeSqU7dsJe9CBvKac8gozJsfUGAGo69xuQd5s5I1RIa+LV
aLNi3YaoWaBT4o3EkEFOoK4lu/y270Tu6fRLRuKICkiic5uvXWD3rY3VpJC5Fz0G
hioxcUKNrn/8qNJdCkPbKU16BWb4UdGE2LtBKnuwkEHN3hP2rfjcEKpq5x11KY5j
lk8t9CnPmUeoz9LN92MCzfTDw1M+lUahWVLXfxTYibQ1wb+Sdt0PWOlvhpT23WYh
N94Xt1WWWJNHHs0vRG3j9/72QA978ky8TDzxWlUl+SpbaD28hltp0aZ8xIxlFMWf
Q6lg2yZ1FGvZ6p1n28Pt96itB1tKlx0LrPKrXNbasO3vcy4ilhdCb2B2NJ2N0v6q
nREj88HDY4nvK7OO7WfFfBM0fYPV8X8TWA0nz2RsM4E5xF94z7vjdgQ4lDyeKg9v
NtlDNYPJ/odsxpfwBCSKBG+MPso4yFX83IyxbUPmD+prNWi/mdk687dEGV61zQYl
SZhyMFTXvnCkz9q6vgqoSI4LEke7oLmfHwxCdxjJligUT386Ny/LtVzhjJqGeDQS
pZSFn3bdjddd3luA0J1WEvWlgUGWEsjMgOioNtBSD5PgudI7y/gRxZwnKS2KFmUg
Ho4Lw65jC/FIQHmIfF9AECM/a2cTfUUIOC2qGapvDLOpCtTmJnhVsyXxlSQAHY6N
CV3maM1ViJ2jR9dx5+wcQWBeXafVQkG3ClhzO3o4cul1Qx2zOUo+JJchSI4AvbTe
Zye+Q7henMOadZm7ptLW/MCLaogmaeIj0y3tp+SKyOk/uNdwzOKGupQd0qW8kywa
qVwimjIhESoOnlZ+14kfdJap7e5KaUHgvnT2aqpBJlLkpr2QKhJE1GsFhsNeYUtf
xCFWZKlaCFVy1R6k6TME3/+XDRw80UDqPDqiC2hhWYxjkce2Oz2+Bss8pA2vdh9i
Zq0IKUOcsB0SNZeOH09+pm78oc/KEpxU0qbBlYZYteRAoYB3DQb1q3v+rAlkkZ98
zlybjlkqRokClewWy3q3V06YIZbA3o83u3v3aByVLkxCocEV1xAZ+GP2FmdGiGO9
d77GqwxIE4Phmxz2UXjcu+d+uZEZcR2WswKnmSLFV0XludQehDK6jpNaXMk9/Y9G
TwpWvQaeZ6I3zl21WovsABLclMzZ4cMvLa0drEp5d3YVMwpHBbTuE38RgtJkUT9K
nfu1wn2dniZSrq5EPVPQkif6V6/T89cl+ckbTONxOg28WUj69SduP3qWkD3GmYB3
p3NY7xd5zjfY83qWS2mPoB2uWfFc1aYeMKKH/2PkDGDQqLi+1z43NHqEqE8iex/V
0H7/4RToojzz6ZEZTF4VRm2bgb0r2ooO1ZGOpn/DvujcHGGgI4BZtHWsGZjHoALq
wg4yXflWmdGSnbdja321Jt3FwTsBBgacxcTqEENeO2qtiqTKPq8MPzjWeGcvQmG8
Tl7lGlDjKcNIhqmKeCYl+3V7PszM43fgTgpTIttyFR408PBHr7vREFc/rb38yqos
bXivBxn97wklR8VGaQXpu9uY8/WBTGR9gKWf962XnShxKGt6KQ1NnEqTxjyab2/V
1Zc5TbMx6GrEcwnZHLz0FQix0ltR8SGIzGQ/x/uUYKrPNvsxptV0F24Kdr+USQXg
GOFVaOk2yhTuQ5uIY31Y/lHeZbiz+Q8Q0MhSaz30eykvDtsmZQVq3diOeU2hJ72j
3fTcw94YyHUfM8wZacNmuaYeKII1vM4Ov1LeBwqKZMpqrxpTUs2ZKitOKEjkiT3U
fv4vfSKkmQOc38wRN98t3qb5H9rq7lLlxM2IOuFjQj+jWANmEFIhbVBTYUZ3ADyK
DO0iMmiHfHcImY/rl+HZF8f41T7USd+79g27TngPcJF5B5DGevrqthkKzeVcgq+W
e8f7m6oGtH8yM0+b1fu6laqIbMH4AyKb/D1zji0zC56fqq3jp5DnCvLonq+6woeJ
NXLW7DDRphDwOLejhsZCezUCZ+o35Ol38SZkOJjdEP11/Uvj8sP9ViYeKC4EZ07y
AVYsspXYedw8CfFABWVyMfySE8LSNagQqYX4IXA5QWAT8Fm0+42cM7RThaoi81+t
0IiFYCMQFpc3+m/K7fkllRor6Y49zvLvt/PMf+wgFPvEX0DWPwBcRCPdpuuHhV5N
u8hNRHH6AxVvJiSojeAr31gGi+asGoYCxTasWrRsQzbt+UQTHZ/gIzmwohFbZyan
MsPy+Us+rHQolC3S/cc2kR0rBYWu6yl5SAK6bRCXGiEVNFo64/U3GBCSNS0+qnO3
Z6ws4+LijWScdYcoKrMk7SrS7hB5zL4piEXcrYkJZapAVpO31622YHoUpr8I2UKX
KQAs9842x0mgnZjekpr4DPMqjZnvKgLEsCZoI3JCrp4BsfdeFjY/WrCPuwDmFq/5
LGcFcvl9SWkvGE/Gdegg9HxnUSKELZg7rStqkZMmURFQi8sEC27oNs8/17qHY0Tq
`pragma protect end_protected
