// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:39 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
aV9TsMD9tJEr9z1OTL4VpTEIxRBVZJeTuRSbmUIEvNGgUoxFDhNeyf7qgzfsC4B/
7PFLlWcWkP41HDWB9I0PlZKZJEoVkYo+sZIYp1kpf8otre37oMKUZHxqy0VC04Po
YhydTXpYiU/vdI6HWwuqy/Z6XR2WZdxPAzsKuobFBwo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8320)
n3yQSD5Q2/6OpvGo5TZVc77+hZTEerOzuDy1lfzehJts71hlxSOZgmHOFz22+wgQ
xZjRNWzUtUADveWZOzrjiv25MP+MuxaRRuieytMHxpLd4LNzgjFBD2wQ/2+lL+sd
UwoQYwW6k2lH0dEvy8WnzBeajkMGm2Jvu43V3wV36K6UxX9UZZXBUavO+ko0NsFq
2rEov5eFtfwZPM2oQEvz62NidwbE1+glAzyx4AsFBvkSEMbL0vn11vCOfpX59D7h
DeJHTZqtN+Fu6O+P0epqyEy10o46MRneUAaNdO+/zhp520+2NWY8Aj7rA6F0Bdoq
OnahoPikipQd3I1mJVc06RQuvciOXeJ1m9NWii5SyJldMGhfnuFDUWu7JSnCMAv6
fHQRgD2LJJtc6jNeeG0uBES+x0fxwlWkLvNcbr04o8kG2ZQ9KQNytDDF0k+Mss9L
3x/Amb4X5ApeSnPVzUsjvKiEKfmukUMP9cbTGbqRJWt7rduw8t9v3ZRfMmQz9jcu
vJylQtfos8tyZBtV9+QgdC5mBYWlUXhz3Zgr4sKhXsUIIB1oVuApN2J8q2kpkswh
1IyZviNqEOXerdftCCmOxCtbslO0AG1rivvX8/qKPh5N9YGQ2M/U7tF20zEErgyB
BUy6vIM4NCevORvsFAYERxJ8Gwi3o8Tt1WEM0T4NHZ8xBXfmNng+MmTuaGCN0vEb
mkQ9JKiaQnWE2aVej33c+m/Q55zm13Tti+mWRx6dTlj5ZJGo1T+kKYwSR1mbBQMy
UkJyScAJnEr/LN1o5NQb+c5DSwKDUsNXaCeg8Z0hvLljU08gPCt8ZKQyvU0xSt/R
D483j9DpWMtasPYJ3nSGydN0UHVURnrPJYK0xjmX5w4eDeG/0jK9dR0R2dDMucKI
NQps047S2b1CVI2xFnAQShlqrJk8r0Sxz4acFnxWdRxI+zm4DpLDLcsIbA0/4ps3
KoLdCLh96oNwTsp8/fgSBgc+10oAV3sNyFhuLRKV8/Hg11B+pkFr6LSMEWZKXb4w
Y9qHrg7fKqta8idZxBTFeDffcNveFqa9JxFiYAWlKXwjQOsKxYxxuhYYOxkAZ8AC
gkI4m2JN9qhVT2HDnofwbW+ysXx3GDGSgnerMtIOIP9GKFHIfhW0ftWyH+pVOPrP
ZjI4bOEEgfz/CzHM9HTO2pwx65Xhdx4mX1TbOvyMVczX+5obVG1/k8z1ZPJFF3L/
cF9jyKma09SyxWmNzbZeFLCxC0RCcq/7F4ydnq3kv4sqIWs/z5WdQnUAcEHjqKN4
mWEorTz7fCbJbQ8jx9EZtRY4PETRi698+HgQwrf9T5Ajhs3IHqj2TuAA7A+K1b3H
nWJF0eUAeDZkCgryar+4RtUCfnM2RUvr7xnhlG2ja5HWXYrdkzA8Zz6lI9rssSNF
PJ1hZnHGaoEYK5hHHzduGX0C1cBCXFtbKKjPVAK1y3UNU+y7Nx6/sW8a8W2lwxxb
INWMOBWs+mqhaBZcpKuzwjG/3QjO0roeICg8CQ4FyX/mjGhpmoMCRR4Hx9xrVWrb
wC1/L4e5czQ1y9LXgcXf+IoJggIMyri8kfqlLqCPWRXup72Z2weZp3R3aavskG18
EzAdEqLn5XSE3ziTjessm78k0UVVGDzu6098p2nexNMbfKTvvgB85QetBkoUibB7
9yVbL8o0aVX5QJO0jqkF8G5kMcRK24TnH+tF9ycGdc01Cz36PDYpcDyT124DhiS3
iSRkO9z2y24ylkaS0FuxN0cusY1b3i6WemPXYfVezPQuT5mR2F3qEclQJjrNko4G
0bC47pgBqPbqPlGbbU+ij9r0RrSTYDjjrPzrJhDVsd7dfA0ylmtYiHSf+SzhAxOC
A2o4lemq2HT+79za3nJc7iNmkb/3JWaTZLBJHt2nneJkwNmqyDEyTIpGd6SGuhcv
UYSd5vw7R3MheMPaT+rH0jX/4t6CCRKLaVVRDVIyBtzrehndEAUXzVkswDGbpUyz
9gNjnVHr7fwkM71C9jjKdUpwX70kGjkVYlboHUkRBeRjUR6Ok5vZmR7euuxB8yPX
ISFWVJzf5iFgy+vY/5qsKqCsbKh56UgWIpcXCSZdmwpfRj5PEkbAFSugNDS58++S
LUCt453xP7S0QRdWLOT4H0o+T+MrdtMfZj0/k5mkifhkDb/P4RzqDPr2IUksfrnQ
okzUFKyouFfuz6856fNQYVjoozBSuu4gpy36D/NCeBcPnqa0VSKIeoOr2TiZArhO
VE/S7X6a/CNfDGD6vMlugVm1igDhCJlxl43nC/5iuN0j2R/Z7HYgLAO58PuPTs1r
3Jp5zZQoC+PEgT5A2NaU9g8K6Xnu1H7LhlOhT0qG6VA2VJttEkGDxB5DEg8ek0cl
3eid3zxabwqw2G3p5kx2nvL8KgN+GfKNvYzFX17UFFkrd8C1FifciFKK/9BDyVdm
n4ALlDbuVXpv51jfIzQ232XsZHDF/cvxMtU9tvryImlzIIphACasauxvFoIJsNi5
K/62fnQ58eWypQwT/sdzv1G4ZN1SmfY5z7weBHjoxweE53AJWNa7/ZV6q314trl1
RPAISt011c+Rndy4EfFQRt79ojMoZzo0n/NUR3s1f9VYizcDcehNH9HDrTB30Kga
Od9mgVmGUI1U+k0c8e4YHrhBdwe1dQg6q+PyV5fDAaEwGo6wwaAmbxd90UhvOQse
VHQOMLs54FMoLr3LX4r+13sIsE6rNh5WZxxKt4oSfZPOlotIPJdWOG0MsapMs+jV
CoXUKW5KX3vG/tSzhogAx4spYal7TC1focwiXWRLs9Gc9oygvbJVuNNmMDCks8ub
GM9IwJ6axxy5/L7ZRPgCr3Va47sP2l++PtLQdMCyqAfDMLvOSXI01rlvQ68BU8ec
J/YBguHmiRSIKNVge8AjWIlsMxL7PlK+Ka/8M5aVuMR+XkV0QU6ktq8j9R3qa/Yo
U5nR3VVK9OCGTwsMwWTmJ4kwzrngqThknBY5Gy6P1Nm3R06HQxR6bHg1FDIit74p
sUp+aaVRXAQ713F8sg7xJNtPhzAS7d9BEX+6MHrgTWEwyFwYRdQBBYPRWAvCOsIz
hVIuqIwu4QsxIvdSzes3sh9mneW1XRmQ4DWfHsxXjMj0W6uOeUpAbDTHkBA4mmNa
g9mDElsvy7uz/4QQZHWZwY4ZIL+SSjsLHvEF/IagGFkFRNfYA7k3p8qPSlDDiJQq
+cSelHOWSy4NxqrYHYq98mKE13DNZ3dPOiSgSqHG59EJeMA+E/bPW7+eqZHPzXwi
jBQuUxTPDH+pHyyszpA19KCIObnVa65m29pjvIFrSWo2o/GTlph6RVb16x8z7niV
C3ERxo+GZYAFz4N3N6Z4v9XS48H5DyhVmoCAm184EozT7bhvyOE2mIR8cjlle2sP
hfWEdjzNW07PxfiiCa3wuL7EuN1cTxmYkJoHd1yOhzBQsVOte2KRpW1BZFfhEipG
nPjcjPSE40VMljMUieKpTejT4w9zlsexV6SrsJXCbjNwlxEuRg25NpB0ClbQd0SZ
+5to7iTqFqGmF7FVEIe5FOvOOYe7925SzwJbquv+xwyePfpBoPD0h+6IXYacuTRK
jbWWeUNLi9bThDHD8ffysBq+Nm8dpD/ovOfj60/Mp3lzaOuBGE1ywnJuQ52RzquJ
sy05nBqM/1iUiTHf7bw87bbI7ynqTKXrM3GxnUM113hYhqe+mez+KyMMjaYEwEOY
9k3L07YoDrC3Tv6l3PT4cdG+2LVn3g4YCloLedFftLEAjcsj2o4dnMNG3KH9twHY
bjzyD80mfRwiK74/WmMQjdww5f9qu/C1K/WZDDR2EPUjKUaA7r6Zh+vAr1K5ME64
9LgYJxCUH1Gky8y9lKk1QQKH2IsSoz1lOhU0k5wfJmYtdtM04rQfVemstW7T7OOo
1yUTowXfGR+QOSVZ69TIl637b+xyslcici2xq+Z8GXa33XUJ1KR15hYQfyv6fkcO
g+Bf/DA6gCU5ODI/+nk7W8hp5yE8PbkFUYMZMJkHg21u8BGjrZHG64BzcqiuwJ9z
sND1j82zyLJFTLVRmI6TPob0kt1FhPiBXogIjRiHdI6OGCIdzWvxEtOWfdtGJ+ZA
/LLicI0dei65RBRFTGDZ9QBopsgU2cakt756YYNop6M1nKNg35qJJ/n6JPVeaX++
PAK7PaA1m67qRkGxGYPk2d02XbTFqlcXZPoE9sDJ/RUhdq+s8IBo7Hjzsxq9K0G1
JLFERKCdwOSir16uwwZ5Bm8ctVi9UyIkzaX+IBs5HWo+TRQWcU7D0uJUaWBttnBT
GCvhOKK8Yw98TYN2NozrTy/g9sLUGf2+E4phTviqBi1K8kUEeSy4iBIVGBeFbovp
+9qYfffDG9UpA0q+nypJS3AnRHMqK840vt7aOZoBgajd4LX+Fs/PjKV028Gx4xsf
VvGBnLBffW/S5hKPMYFyt+6xgy0zKfTsQq3uXhVlqwtvA1u2NqqhDrws7H52CwT7
6L96mIzNXUyfMmZGzMFAYGHqGREi3ZLihBcN9ohg9NzQYFKZF2Q8ygOvbtBuebNb
CDA71NhQJ/k9f6ow3PcDJh79COP60Hzh1fZVzhAIe8cDUeMjBIq/bXmhr34LJqcy
jSqoJqIwGeUYhyzyWMqapx9aFCTIdMlGEcm1KHPySwdM/OtsG/Yd9SCFfCGvIOx3
YUVpc0aUeNOHX/d1NAR6GOCRSl5DlBMqbWwgENSt8vPvfSObTNiIGjEPHDwlMFq0
GZE9hJQCt+ccBqT/hD+BxMQnvjirNGHKDDToD+DErgYTef7/gJKV37HQ3KXFBZ3H
f8upa+qgTl4caZCkF0thLhhjT5DGVQVQiNpaeuApuBKwlpKJTt4yTrKHfviTGIAw
LQh1Ge7NSHgQJ1oIuKETbBnbNT1TVeIs5NXzpfvo8heQZ8NJqTR+/k1PF/e3ZHdi
0sHaVY5kQZNLp+gRAYVaUyfOAox5QVMSTKsEAYnUMUsv1ulWs3FZqADklSQWs5+A
QmDZjdtAY4yQI6cEnGNtrOuaj+ErBw2t7KxQx+pvixiw+xVSS0A3Aky9y60Eryd8
Of6HsOpAFsSOCUBX9ED2JxH0/63So/zvZjHlPUKZzduvL91CqmSVHOs7gyGSHEfT
RlC9sf67JqJ7tCVVENUTJ2xccD2vUE7lMhyIxzhlQhfijpp01imkYRCFOUH3rkw5
nyQElY3rvf8U40oubVEF+SMzlackH76UlomDw3L3/U6ur4GZV4vwkZAHosaubZqU
VrXIlAOFRDZcBH96CqGoubxT7oeUBITfhZ2Sdw6BoNrNkCkju8ASjesnl08SeI30
M7mxym4bzDWSsIiMsFU8d3TBecoPgKdoCtzp4gcnhJgIGYzHlwlOfF9xQ3pg9Pa/
JyLdEzOxb/OAJ3AVdx4qnOGfijt7UUSOuapHTbktMmkhmLqGV8cELcdcx2yzHnc9
B/ZMbPTDlrsjaQiDjwMYaTj3NxbsECKgdQGPRiJTsIWrj2LDw6zGCR7B8AN+blhy
8xK8HCgyA4cuoYHDZNfJPZAeM0RCfJXNwpdc3LGyjvO5ttlZuYY+Tccsw6njHZ6W
3qMBm0sbhKOCE3ueMmmpJuoEck5S6n2YDeFcgeFLSQ42opbBOF2xTKgneAvwFBXX
Kz+ojTKav9kNtWbzyGQ2aPhDgvTfJao3w649jFfgRAibgil6TsSNttv6lk6Qzjdg
RDei7hj/cXYjvsioO9++Kn/kABBsINZvdP7GmM1jBatLYXm/fzbTBa5hhyVDMtbf
Tt3/+kFz8q/HlfeEHxRF5DANnq1GmyMaT8dtsJpWNynwMNIaI8ns2xhYB7yAf6tQ
Uzch/sYKl5BeCrwYVM3wE4uKc4ojlwkfzInSM66/LPlNoIhDhKRLjq/ZCy2ft8Eo
R5XqCCwZAD9SSjXEL2hRCPIhYU52Lh/Jbzze+PufC8tTmBLzYBZt8Fa2+OvdY5eT
4QL2+t5v3TRs8LCddlptrF9lkYvELHCQm9Xx0Yk8OLSBYQVo218eG45T1hdgs+aO
VFUwU7pMyR3CbaoZntXarpVa7sfnQ+5XAg8zPQv3sZv1Qm7fRrHcMmOX73pRO/AV
r6kbbw/YpG5yhZv06sgQen8RAQDS5tOAf1uVsF2dPZdM/Iajyv9wO7m+EMuqn3KH
vh68nMFMdNC+aIdhOP9EodrS5IO5zvdC3T4DFJOUM807ab+e5f/8NJdmxxe7xoPN
x4Krl5YtrVkoyZX87MZwI1cM328QQdWJsCZga5ReSGQ97UlmuA767nMORY8CwhrJ
Ug9EXokJo+2XuAczBVOBCW8fKfyj8v/rdh6zQGOOjhopSXqLSIv+zwFm5O0eX1d8
MROua8q1rGNAjMah56+jzPMHgqMR1pS87y17gGBYptGI4+IqSGoutsQFJqyWDHuC
Jg34WeQzndY1qvJiL6A1bGim5aJHHU64zGSEc/5POJQxd4GQL+c/rZWHb5I3Uwa3
T0iJ+6DItAQSBxugKUVxAbWhHpp/St18aoreOxMBFNvnrDpFDIqAiN3kUIDQrHcT
QdUcpiI0PbFe4yQfajM6sVxKMJCsyXqxlNtqNFHHn23VvoIP575qM6Ju8kMJZbJz
kD5oU4ppVHe8M2pwl2JukxZBUsamMJGBHbJjPq3+CNbRRoMXJK04QNH/B1WcoAMf
TeTSkhbBsi/bNTFl2qGghK7JSe2Dp5o9MsxVDRLPn/mOroMzeZbsQF2KlHcs9H+m
Guv7XgiRjRUGOWvAqnObUGFc2QpWLivgMqHBGsjz/zrXGOdBk5Y3Y2gDe+p4npo5
5+XhU702VgxH7Oi/kKO8cVdymPD7xc3KYmQcXOkP8EezoQQRIwRVGqKMMPhNb5Zz
XVyTJCPfjZmc8dhpDnlr3G/F5r3QXEni16yMYqdVz9DulmtOvPBXgXyc5ByPG/h+
lGUTFRzcYGpdyhvJeoHE4h9dWHfuL6iTloRQK82rxcirM5n06KQgr1P/IU+W0q8P
TqoAXQfZWFn7HykqZ1kg+r3lDpYEUNPL8TXoYf3epQBEzcYi3waxKXl6CtCAjjGf
cGjvhm/lAkRFgGB1VCaomk+qHOSdrhNj6TFvYos6E64AzUTOIbswL0GnhN6auQxE
0RN026PVaPNhV+7kFouheyBgodpJqvb44mu12OWwt6/Kzd4URhOBHlG6R65FJvZE
eccIleg88WKklh0IvlVyHlWSZOD2RtXrjfrIDQ8xd+x7e7dnWFWkbpzDfSTwzqsl
uVZzz6cmhPQ5uN4HUFECw/XVRfUQO+ZOrzEmuRGLj17gErL+3jCyUD9Fqjb6pE00
9RGq/YykamWMR9M8URIYrnFnv4EYI7RJ3k5ToklfGqlncc2Bb05bjDV+CRrREWSf
9pKKM43KvXfaoLAMPrPqayunqDViS3ybrkpuIsD7WbnbJAxUwttORZ248TH6koyq
NYNLmW1iL209ziVaWH6fws9/avw/IEdewf24GT0CC8WWBS0LPDlaKDtP8nGm6yDR
WO7LR5PRF3RrpIwdJ/51+2UdaENPNoh7+gpQArHPKpBfp0TbmQwaBDVlBV3aVPWK
3H8Bx4KzXeLOnQFJGcj8ldsChJB+dANa17XSqQ6Het4DVPqKQQgdDrRMxUh+zd7q
w3ajJYqos/AIZniwUs6Ltio246N2/xxn5q025Y1L4m1rIc9pXsYqbV635lcwau+e
4UprjI5kFzeCNoAykRuRLfzDe45HFh1FcFJiz/C5Pij/MokkWWhZvt4AbDw0W/j5
TWr3tOQiq6by65cckJriKrJXRp9AK7icRTKuxo1c2ICfi+QMmn5rFqhuOmGwhCQB
315M3MblmtdsJR+W7Mx9mfZrnye1dIXQmNJKomyobr1pHcx4YwEkaS4Da2jS6efP
omHhlGcVZ0wQYyajZcSVJc/Fxs1L0PetGT4AGlu1/ome2lcx4ICHlCuaaA1QWt8J
UOHeZmPy5UMe8R+dJfj+219yIVmvN+FyLoQy9bDSqr4V3Rm74a2OUZgI4hCIHjsf
VOkjNJaov9JximBtugsJLB1K8OICUljdPue9P0S4MsKrjoy0JGaLsRFX5u5BrfCH
A8gZDVBAJBNGISW9OObDXIf5+naQRYSEsKnrYO/PdV/grSESo/xSD8Lq9GrHfm6Y
Hlcmviu/CzuKteWj0VjeCm4Cj9GzwY4g63/Fz5HzVFUWcuE5+Jh9Phe54GlFeXDK
8pRlKahVEbAucRY8ntPMfL+fqLu9o42MfXFuyFCiVPvk3q4D2F9KFEdy/5Ij9X0x
vAT9waUmGiVOy4JFu7FDES8jCoY4/OZ5qSgxfbBaG3LXvjL19lQCBsD76s9JBVGb
dyC2rpAw7xTT789beM6niGpqInXOElZXgXaV6BORBpJyMXbC8eNA0ck3Jagl9nyw
QbOHzpcPk9Dtv832dPEBFiT6XFp74qJRK8VmRwuP9OXXJLUSV56DBdM7DMlKgRhY
HYY5jMd8iN1Bv2/BpP2miTtfAtcT/rfxD/M/pqjWtq/wYV9fb85mR5R9e9Turp5I
0LXCfk93ppmjzZPQd8Y6bzWnbk9RojjCrcQHAM8iiyV7n2/k6s3cievFVhtnBn2n
ae28sc2B/Zc++kK1XJ2dTtj8yKsBAFGxj7wRZrW3RxdV2WCh4f45DG3XixyhHREc
O2fe3as2BqOkI+g0uHjIP/n0CLjAr5BG2yVEw2eMqwxAtq34dMi3Re1peL8XWLod
CAWcn4vs1mzAVpJlkHRPgCI0GjoBAOXsSRewZsKSTbngkq/q7uPucyWYjusZP8RS
rUOmOvikh2cKvCZuNRL/Osf00+2g4Pydugk3+xid5hz8vvpelEbCCLtPiQ+YTQv7
4fIZCmiFvtZfJUeHb2Xq8Ie8rK9xe6UuYurJUZlVWodmkNeFYHwrEhkT5MNLEsZb
/afFU9GfOZPUY5eWCK2uGtRiaOdaGh7EohLhraJAiir/qIKxQl92T2EMxyL46/Lj
TI2SKFhv4npqZ4powu0dKWkrTGLJ8OYXIoR7QGONPaLSa0kBVbsSq+vkIbHgHBtN
JUr4WNnPnkbPn4KeCoOSVhg/VQbxzmJNVltN8o9y2fVY0HqXySLPop6TA4i98HUh
ILI1LeR3+7GbYXw8pCL/b5ji9fm3ACfq6WWnC1fWV7XNncTRW4hEDCuPxOo67XhN
mbVhgOJjiPWZIsd6hisyhWvlZ/rJxd29mvcIy6sa7xGOrw49AED4opfmkQZSof2k
0LFSpBcBpVUYpK1AKqmpiWq78CfK3+MSUloq38B2tVS9I0PIfVWhJRrng2mBKc/4
eILAL9polUkddf9/fNSff6vXV+04hmi6F9rReri6B+1ZER8e4o83OqNThKXZeQoe
NnZbwZSxLb81GFOIJ209a9lEnDvI1VqQQ88bKlS7bPwt9d+zNsX/5df+NeecSTuQ
AxtSx/jvsi8Gd9iVozyyPty28kKylCfs21zA5l7pY1ZHdZA537dNW4B004hYFFlV
rghkhaqABu5HiTxUxhAuLrckcE+rz/G2KriCo1WSOOes+YBYFqJhfImUBzy8VBeQ
3Fvdoptkr3XXvg2OkCdP141rGeo0YVk+IhusT7Zilp5jw56N9U41X0CMTFnW/f+C
soBYfqpzW1dd/hNibHNqhy2WGx8UkhVjkYgFXEkmRJVgM2WN6cgOvaTG/VR/fxd1
C90R/cXX4nt4qkihAv8S5eop2tFZ/JVTtRH2Wlh3jFpxga7Vf5RR+qmsrnNoS1w5
pu1CQZNAoXaL1Hez0ErHNrvgbidwPJng+lRUkqJ3pHmfiS+uPw+4wSs6f35n6fZ/
PdGIyQ99TtCP2Uq75v3335zAU4ZRmVo+BxM9jLq4O/6BSp36pNUvkIDT30tMn7HE
k9s7rLwJMwFzZ/amjFJaKdvXc+2vpBKYVR3seYZs/DYrrB1d1wEzAVTePs+rxMDd
NSd34qSB2a7RS2wzBcAYMp/cxKlhhD0SH7YjPH7SMIWoBvxKIpPw5Ca7l0JGxFxk
b8PrcMHouVqVbVhawJUKiFFpet0BUIT4Fj1zbeOu6s6FVPYHRXPNXkpaQ9CXaDYl
6Uh0US976UnxYtORayBD/cdMbAtgNx9IMqZMtYRnMQpr3+Rlx1+B2zDMowfQlIB3
QLBuaXNirs95H3plIT1HZH65AheHeeKS/ctAoKcsmuDGKR9cQWKdW5F5gkB7fsMm
8NPkbeQ/A8PNyPaBAyY14zTfWXSZr2qotnzFNjgJ9PoBIOki9N1SSFEZRTDrIDYG
GSltcg9dE9W82lFDe9h+u4/JtuTMGP2FPiFvTIThIsEjnDXjn1NZBsmw3gP2Cv+a
DzzQ1dedaReW96rislDls4+c3kPFlIG33fdOK7DCk+XuxfbZca39lBoBF5DxLehU
bGW1LswLtThXhsxaoiwLPmDhcgwVMQJ4GPSUHpImqCxJooNK9oXSzCW9iB4FHVoQ
mMt2EN32dhZKyJy2MbTiDNdan5C7o3af1WHe4+aFycyVH8LNw+P5hcNmSjQxVjfn
lbQQ7Sh95VbnDOdTQxnM0hWACgBXaiDrXQeDKp7gbcKmUBXw3cJUSYv8OsKkKa6s
awcTxuzULu0fHJi7M1zZJIt4rfY+5EzKlTK01y0IaUYQbvSKtLEwBjs/xqfnZgt2
OB0Dj7bVg3uo3k5hibiEHndj+Bpgkm5GQ9Kg+sjdcxCEDTj4uxDT+8h7BZNXNykO
SLUw93Dz5nLtHZESm7OuAGxK/hN6v8aYOcgA3Xngt5WalRxcxuMen485dl5i6EWF
Y5VYLL9+EDknnEEk7vasyZtqBypg1QqYOFwyVnCq+9jqlzu5iJRp4WioBi8lT5O/
nJLAvjJbQMK2b3ew0j/3Ms3BDqWmCs7+W2L9j9B1BZY5GA9JCgWAE1Jd5YmsFWE5
3/MsqUvVsKuJQcMOt7+pl8cX+jJH38s8TYzbiCoF6FyKvH3hOxTppyUlJR1Cf0Ax
k1kOBxWMijKw3ehitEENibOorJxjBv+onMx0XeMENvJEPPwJSPLPuA/+c2Y4DE1P
mYL1rfR+SynzmZqAPb9DQ/uzn8LroPf23huGo6qS3RyIMDetEN/2LtQ92Rq2n3K+
/hmvzcyjMJTO1pPCqDIRpw==
`pragma protect end_protected
