// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:40 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
r3tQ6z357p+r8scHTTYnlCv1D7GcywG+oz7j74oOtHRJmBKQsEMyOH3RNfb2KnHN
mevc2GkNZkoxkP+zbYWd2JIxQj0OJcr6OO9wXVgdmP7nmN1yMkBMoXhqaJ1s4wmS
+eWSH7tjlmHGhiq6qBhdzoiNILIT82lR89Qm88rqwUI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9472)
JX+sCuHuAiH24RIM+7E6t7deCtmjxaP9GbM/3fRATsyd+fxHf3EbDOMkl55nLGU2
O9Wyde7IIU6FB0fXCP7d9FVGEW1XhBZ0n8b3uz0PMngC6mMZ2JzEN1t4ExvEs4zT
mzw3l/+UU0Oohc+ZxjvzSaNdW7VPgnVyxmWSMtAGWGi4eAWKq/r3C28e+wLb+uwP
v9A0D9GN7dKgJiRwjqhottCHLkkowO0kANB9Fts3q7fKoLweVZZsn1vNBEHcZUMB
esURRPuJh77iTgbl0URbXjEJbyaRLvmT3Zvw/AhLPJCFefUJt3EMYwVzAv/F56NF
4VGxWic1oh30s744S61/GqK4ymlCXKDiYjGmRCBCRn7GhZVjQxcQ6MNhRV28aF3e
YoDenEAAvqzuTTgic449y7tbn8+1khHFr2M0otkEfcSnVW1bADRJdXADvTHFsVPp
hgz8LUIpO/rqLIHDbCiPJ9eIH/BgQOF2PmsgELBU7wtm1OwnDhl0APNwgBso9hfB
wnoxRHavmnlk8BhLA7upOSzik+3A0be2bWt3iXRmXx+Hbu/BnBLwzAf0ZgiDjh+I
5e/IxT5p9QXECIhglqdzBJYvTfQvIYNpZQR7MmQc5BxL46HD8IudTl5B3sxk5Y65
E5JtR9SNFLKOhX7ZTmRd2lUT3PvrkDuE3o2J3WY+i9qkOjmUX/uTW1yOO5RMIJl4
nVaKldyYC0F666CX/HJN4vo4Za6V8YY7wTNVMQV+mrFgmPjuCP9tyr6PRwTG8l3y
ldxd0q0DhX7YREuPhGd3401uS7P6AWnx/V0GYv1RK0CcAvCMyVUZKSttXwWa4Xq2
irStgPBPFlQrFI5GmcJ09btm6EcYc5UbWBn+YAgMs8n7eq3tFzo/2xSPw5/uGVBP
EtZfZSmVM3+Go0l8IU7X29fomhAYfowrFWBFoDavq1eSV65yYAbMEEZNdxHo8caC
0nuR3mjCpowhcnMmkiOEHd0MhtGmy8tbI/QtIb2NG0WzFG+bkUqS19PhPPXp2zEB
AGB0Clg0zw2lz6z0W4EwCI9u8lycu/tGWegL73zgrLixxD0Da6mvnAacAozP4K/3
xVKr+fluGkFKMjdTHeGfZiRTw0XaRyOY39MRfG03QGODB6QJOifGMhFQxcMeG6IP
smajnbRjkBVof12dRs7ndN+tuZpzW6X3D1VhVoJscgXjeTt3tYR0eW/WSyU24t4q
xNPxDH2JlKDYFlla9XzFByuloi8TfQ00Pm6cIsE1z6SU3rJrtz5ZZLdaPHvdTZVW
ZyzEcMjodl7W7Lkj+pb9H5FhI33ora1R3kjoXlPz7yEcIOsKd+dP4TlniRzklSwr
c0Pz9RfyEnG1R+xOcc6sJEE1bWTnepKlDXEjx2xlyjWE7G7n3uX5pvqvaxcS5g17
iAqV+RtRcW2k2dDFbF0JEmnzb9bAR58yPbbUro5zNRNDpwvwkKKOW9lk9SFiYXnp
WmSfdEHtvAuCqLU1rTUFlTb5wz53AqE/Euh10nFfDrESFu5N4Q598sjQwZHCf7ZZ
oo1w7GtlTHbze9utj4CF5seKyEuUOK87hDPAYwEpz8R90CAIURH8iLKxQukWED70
WhlDjR3FCMTq7k+I6irAT28EWqTlgKufV6BVnCaVuSo0qjJFyUVmSILKVL8ptgFs
IHME4VaKEXNOyFbwK5VU71q619evDQR+jJ1RdOas+FtTTAUOP4UzymjsAyw4kXFS
SALps0LQPz3KlVDCS+pDMCeSprzl+VdkafPSOKdjxt0aZc1MiL2VexrHV/TjRwtt
wpnDzv5LGCej/BLYUK7yijDvwlGHdCtVpC/SYiFOrdGQ8AvpHT77cIrJ4R4dKcEG
7lvZSxYF/7UStKqQ8dkSxVgijYnUXbpiGlbWE5iTm8DzYMx32bbhqLS+NbX3WSec
T6wSNOqUxONp35nYBY7ZC5H4acwmudPuhabmIaKzOjVGI4NLoCoMceq6adxIsh+/
jyg+9Lf4TA6ZgABzfTtw+//NKsA0HQyVZb6OYW2fDt22wD+gmNGLibv/+Akq6pxz
Jar7h30lI+bu4OYL8gF6Ch6PwHIlWaC/XY8vcGdGt27QTnvmnfoRJ/8vdrzS9SvR
hIvVKqCPfJMBRmMZVdh+5W2mplv8NDS2dmJdDy/dirE78bb0r2ywrw3Vu/IdepBu
yt1RGLaB2KWT1aUcLAdoKFaV7B5rrFnLw9xJNNtl2RVKD5vEGsEMsuwuqkY07AtD
DH2GVDvnB824q/Fon4F3/TuXQxiTKwjmdzJmwwjcU8u0clarXGYGcybew7oTPapb
vx2aq3AAfJ46qrPHnZzzA3gQKBuyreY8d8+kMa1kcxrd9UBy7eROYQZ70bagUmF+
tEIxXc6TTpeo5WDVuPjmOEiglsZO4ncdtcTJFQyyq4F0sTHmvBok9+VNuK43LQOi
ZeAAnOfFQukoAb3H5OshjwmsLsfrVjiLIupwuANIdWVKlffbjghQ2tBh9deeKOvQ
pZdWSKINnSuAXqWh5iqJay6tq0aRwr5By4KvG92gLjfXJoIhVFSLnhbVEzt6PIiG
D/oPjRKTB3hzWfwtlbUj3PIKoUZZOS9jTElxgCic1Y3SsZuSDJkOIvSs05NN9gtj
YcRCtwHsvRAPuPWXD3JDHZsdS60kIQosg0PLy9XL4SJHlCzZp0GgRqR2YW5EqwsN
8307tXMrDrj8+fYxi02CwEc3nJEj2866oimlFEV2h6fpSulUXJgtJ8W/21kTfxET
6r+cd2mJKjSDaOXgKEjgWsWSU1FvbU0i8IL6Xld/LsyISbO77c4VNflxLcXCQq37
BTOZvzIcGRVeQAYZ7YCy6Wuk6l4JyTetJeCV4HUD9vMfylygWLuepm/smIj6dWMx
H/ZWhWk6pm8TsAv5whDFVBJ9xW3oNN7SAhqC5Tfsy0wWyNkZSmGb/9DLtC8zC763
ZtiiY26Q2HcqSV0RM/VzsMM/jjNIbrYRqN31767W0r8fP/V1iGycN5Q3oBpGH4ir
WgJGNv285i5PUvBi56sUZghj2nFSlc8Bscq68wzCYMgyIz9QA4IcUF3ylCAO3aKU
1ix5FhKTq3ZQ7CPD2J0rPZLzjwm/TWjXyWDFrzeKnsvHyNTJBb7XI6EO9x9YXwdq
WsxpOq4jS3COFtgELq/Z9qZwgUnh0pijayxSJRi7i33N8irlxCDzIZ75yupH/tY/
NfSW7b8ZspDx6+lTdIe7QRA6xzA6Tow+ujkncAHbtNzOU7+sgNIPwQvVoXggIQ1j
45ZbKTRoQj5bF2dxC3NM/2obk2r5QAguQW/7/Ec6e4yVZAS8ihDCJ4bd/IDumDnX
A5mcdsEm4BrowdaFnFI0PrUmhl7L+C60Idk4KtZXj9AfUC+Ib9BOpQcq1TUGgnKw
Q9PBGoGW3RLlgHPdg+Mi+bhfDSZop3i7KM9GRR8Z7sAABzKh/VjfR1zV6XkaRPkS
C8zDD1QMok5sbWz935sjzFI7fapcEmuJ4kVyoPpdNK9QCuM3LdBB5dr4+fXiUznL
PCL/8ftX4rPMX5qWi6stbAa1CLQM3tfBt1DTZYuo2JS1g0j6Ixf3OX5mrqBZmbHJ
E6vWsTz+KFuAN7YEfJpuXRCNgWsHbqIid0cUj9uljueY/aiY8govNaOC9MpHrwRr
I1mF14xGtc2xDDRFx5BpLwh16b4SR1Zq1Dw8rpluZ/YGZH0WL/ZG6FN+s0OWBsDY
6SltAA6pfvwnZn0qWS2FUbXHJPHrdFpx33ZObF1hVK0EQ15dj5sa19ewMukLo2KG
OHqVvVaD6tenymCVNTtVWad/TpYHyEl5CLpCaLAxvkwifAlb/CfM2psQJXul6fxo
noaZC9yqB4Qk4FOYp7GdYyXACfcD0HZoZqjCIagyWe9EgAEPiWyjk15l7Wgc7QIx
3+PNTOTufHbIGGquQWcpIxs9BmFQmu7LqE1rAfU6i7q67ys+UezkNw6Q8D9U855m
dh/T2Smb6fFh4zmVJ0+3+U9IntyUJlKZYQhNtiLNtS8nIDVRpVPwcoinmI+mPsPJ
YHPRRYIQ1jQeT4Ox7FIgh0mEC+2DY26o9+75lWMivNrCPp6H7vZSEmWVKhocBSwm
IypY2bri10/Jb3lS61mgyZCBT5/gb6FcHXyXgrtM+ncMANUhBfz78MA/FDXFycOc
ERqmq60W+2ecaaxqiXa3uvG+ZuLxsPf2MTbQccMqUCJNFB3ssJ/7WJdPIs+qg0Ai
OgMr3nnM3iClJaoEIfXKpt/mGNdyyNbfa1Ej3UoER191di2dyjYkiJaZGZqOi6fM
abtCf5Z7UZQsC3imuhEq9A/eb0h2Bc55tI4IJVGB93r5EzwPtdWciYy7tTC9BVLP
0qfi9D9WB+kyjcqIXt7gLhEmvolO3HnoaQn6k+XUpquD5eqfcniJkVBnO0yqLENu
7zF20pI+tfUeGJA1GDFX3m3ZmSDMazk2DHV36kCjnUjo6v4TreDpNsgOsVvE4Wd6
l1cgP2otWd1kFdJq8NkYXVVvwOy+Ujppcg0z2wZCNg5FuAaQ2FeEsmDrmi33IURC
YELkGJQkiwUSqs1tolxTqg6DEKu/qIzASm2kAAbomyK3fGdhSWLYe27FZ4qmrfdS
EXY1QT9zRYHtQzbUYwjm7W1TuiVBZ2t2YdO58HUlbQBC+zo5+NXqlxKX5py9wqXw
5pv0w7VfMGsAndTX2d3dzUFnUCLfKQcWWBMsIUwK4NamNhEeKHjJv66QuhBAtAJA
BcDAj5uvj9q9CYE3qX2RioMd3PvhDhccXBAl/45rbYrHR/lRyAF3Fr+heeYffhnK
MbeGHIwjm+ZmY73AuQigywDfG/32zo303RzbRKGK0syeHxyPOhBFlW0s3STqnJbz
CFUP2LOAumKWSu+XxjkUfmNK1G0VtRW6B/dWTKdYezytoEd303lWZG68Ptj3h+xV
vYRclAlfcK15eYF7po2X73rNMZWdpKrqH6iy54rlOqeoj7I6/Y6dUvJtleNE8xnb
1YqT9GFpOjRlXN9m7NitePzC10SvucGbldGKbprz7QsGXcRru6choAc72Afthq98
g9VMsCCAzZBeWvupjWUjDUBhlv3Xxe0lHrnD574yDR2zpWW/6WUmWlkBzAHL6PY0
D6sqZ9rMS2AcyRXmLNYPqRRKGzSmzqsdjUocr7PXLE3j4X9hgiLtFuT55vuMa3eM
b/vZXJFY6VWfNDcQjtltzNh8tmoc+vXZYRrhf+ZtLDoJiM+GzukyzN0Me4BFnAaw
nWADPhg9sfbYYUTlnzUkc0Y1nprL/ihyQxYGURVTArOaZJ4u2dvMSFxZvshyHGVH
sMWeopNwClcevpPj1e/o+stCyYUXkPNBUw0Ys4YZVSFjCVNlZCRZz5H8ryWpkgKT
Uttl247wyPKF3WXJoe2hS63jVZvFrNhxTA7+F5u1baOiQAQu90V6rCX05e3M6vvw
pjn8kJ5lyqO/YVQDjUDC2u+V43G07ppQyW2xg4UNpGm+bzEzVrw6qIUQ6Snv1wQr
WKXgL4QPXymHxS2wZqR5WDow2w/+yxb9iAIZHVTz9xlJijGGCgBTQ8Rlh4tZTgzn
4Ug6JLl5mEaCSeAFS7OMtOrt9nDZRy1PxQIrT96DdDdL2bQiG7kYjqoZItkRyShG
phh3G7bjPYBT8Kc2UAWsSmGF7YR9y7bOtcz0s461A7vguYrytS9PzhcDosX0Fz6a
PBRbMLfMVvyjKsfCr+vcFhQdcKbsDqgBptRhfLkXLaEg5D5rRr4AdVTK5EhcpqR8
AsMFZ0YoMENGMMNd4I9BfBwPDhTok5KTSzPqslw93p3nrx93lUYUg+6avjn64GMy
5W7muDUpGULMPxiSVY+5lHlEFdT+9r/eoSGutzvop8LbAWkN0/+c84gCBXq+q2hv
wegFfIcbe2CsDVsm+85ALRzKub/1a+yZKAiRq9P/MDphUODhjLlOtpkTEVo4/vZL
zrKvhZSR7c+72udiAvdq4SddGdL8PjflVV93RQ0vO1lxhcEOLJYarwqkslLigDxw
LoQK8ZfL+SKojbnjTWUpUZg8OblhHQ0J7Zgm1IxMMnNa8oC8jun/4W8LaoeyOOy6
/Yv0VJRPRoFykK0v9SRsmVzAR9Op9tqWpmj6wrVpIOF+346nd91PLXHPWBQE7DWF
x4WENxHOm/ThJGVP7iDb0gzkZ1fTYnYC5DbMKRUTdAFIeVJxzXK7DEy+PJ4xdCkq
0g6iB5YLXZTlTCsyjauRAlhhRUXxjXKNJo1mWHNZtNvQIcc6tTEGrLvbmHt7M1GH
KyYHRARzZKhpvYMkIlwGOohkdt77c/YSE9mg/tbVMpM78LdRwpP3J3RI+KiSu6ZO
TBLnZGj7zPvpmQ7ReUA7UpiSVhXFjgDhcUxgBq6Kq6Osg3TJUJEJc/eJ8Vsk2YvP
/4KZbkOEOqT1r63oED3OxuYAzrPUck71BBygOmf7zpNRBpoSg8Yl1LL2fYR0wFjk
pqZSQq3WrSny+jH/2x7Sf+w8N4wIT2trvFHwh9ZKWwaloXOoHfqnX7V7r3S4L0wo
f6tGgCJ3DjFXGtjbcfWR5424riKkuhIajRAtdbSVfz3FMbyKwuNdQzGaZW0IA7Xp
e8BrlabSlTsn8+/XV282kU2uZfBSVYz8sDV7694PmtkchBqwRQwIh/1TSgTauOqM
3DHct4WTewxeudcAGnUc7xIJA74W28WK+Fs/DTXHq5B9lS3r21YgUbipcGlXHwcQ
y+s2fPp/1yQzn7nTJLvPc1U680tfIQ1OIPJ13SQBAnq54tyW8j2ILcaK9kXhAVGm
44IE9F0kGZe3rPc5h+ZESf0ygUH9y/EhNqPKI1/SPG5as8xroJ77w1gGbPgGw3VV
A2Ixw/BrmFUqL5cr8W2NiAm0ZD96V2VLnwt6E2cNP/ft3krXzPXvYxG63zEqbLfI
a+5FcEwaS8crfSgFqI+eAC+IN60Psy6aB+fziL7Zmpe5EZeN8w5j7RuRorbZ8UMz
kK33JAOCPDWb0qcn2j/PQ7Q21tnJZhqeRjuNAOT8j/Pehs636BC8B1yFe78TkHE0
qBcy92gHtIfunQ+c5z4NEfaBrHln3futNNn38Psl8PrdFw7YtyRICaAWi/8OlpNU
VxD+rWAkCUiTLv8/NgnzIrRWXYdRalC/SbgsxexfkjFTw0XNg8XzAlSbNexL/l+U
GQ9pHPNOtwk4+jROZxnvkDS9UhilUlrsv0diC0z9wQEkFkFsBixYJtnbLO7kq1Jq
cMiUgQ5ksQmR2P+lU7tnCv1jDUo7u2Yrt5q+lC3G7iYdVAO0eUWOPwpJelaK1IHU
hJPvi4Xinw7aTUicQwqVifDajS6+EBMKvLrfH2WIC7Pl4CweoyNeW81oQMvqIb0Y
r+wBdZpZ5WmYJYlLV7pjg5Spug+VhZEPKQ5V6IHnMi8+qzugbWzww0d/0GWtvnQ6
Ao33nT4sgPhgomg3YiIzpWgoWgak0KiPJwxI8OPyyg8uWnhzu3fQtNPVtEsmIblK
eyjy83GfjWutL5p8InX2c1qf4LvyuVQ5EiCwWwEdI9aptKYip7/YBFVXRkeF/LD/
oD6wgOyWOM4MXXcBhPcV4003K/eWwK179WcNN26Rf21VyZjm5MRm3O1nrTXjHfsk
wTiwIUSpeswtMSO5cfPZbAtmoZnUVhow3MHqmnEr06tMG5CbLsEDeeAR7x11BKTS
23FI0xv9n7bF3oG1zQSRkV0gHNfl+p2vSf86nH1z4cSgQYXkvm+HBra+26Z+Dyqk
9z/fqPqlKGvVuhXWd1L8vkT3yZI6jvygq97z8HvujClaXRSodcuravquB+/7av3W
+5odwAkR9s/JwnLxvrqwak05a9sTXB0Y+MKwsx7xD44ymkvT7yX3IW/BwoflSPLH
Eg7NqMHH/S0WTcmY2CQt1OEj0J9ah+n+M7FABToKDGGu/mWF43H6l+2TkiaEoUO9
zlBIy5YntUcoq00Z38gDSP9kYENYI5mCTFGAZ1DHnsLGKtNI8dFL6Qi5iHc874yO
IJCksl3f7aJfLQKmedLwmWtvnMch8FmGkXG7w9WmDNVS60WcK0wHUyMQjyB9NnsV
MWMGAbU4L8VgHutVTvLUJAYSrbGEMoDwbwC7fOCWDMoyxI2WJshtMOgVrTPWiX16
wbFzYYpDHpAa8lTgqlqHssvN283rgRJYBtX9++5/S3F4dBMWeiX4bPbjNEIwbcnR
zlaBPzWbumAImAD/cAcVkgkIQzdpAI4a2ezZGiki+v3k70ki9cLrJ4POwIz0ReUQ
mL3vKYgSpymWrjq4QftLzYyqY7mb/t7jui/wLOAUHn/B6SHOnG1AEPbL3ISw4UUH
o3dZBMijD9CEcyIwzYdgLcM4OZAZIiwiCZnaOvElQSl3J4R5fuh7yzJeGCspc0H1
xO1w+kf7Ly5wv88Pjn8btGUDshwpqJ291McQsrbzrrUGQxH8pPsTuW5MqspJ8pGI
+Ix6Qp1wf6mGadKV2KWXFWTlJ4h0JkVu/vb7dcQc9zbXfX5O1/2p4nzwRsO4bxwp
hZKMcQmPego0t3pjtFquhq3GYpyczqSU52c9vOrwxJ/UemAwuUlgfF9AzqXxj6fG
aMA4MBBz7AvM6u1oKwmvx7jI1mtX1CLfxdH9YyogF6tuBPnIRfGi+wPxkiuF9F6h
SAUKvd06neyAOj2paMDijjPMP5r+xsUj4e3mrFUX5anYy7mASoSC5UyntKKLhzTv
Pz6wB9lidXWsm84gWbI6F55h0IgX1TBgFxOpCSh2Kt8QZU5iv8fqaY19kJLSTCcj
lNSSdSxDF/BLfeMnLOuMIQsVgasca59LTJG53V+AVDGtBUZUUC0+hNk5kO//Fas7
60YziIr2eKUUxhBkef7N5jL3soRulV1T/at0StQCDZzX6FgdZ5aBBBWgMaSyulQW
/uK8aq2zAFrejp1h+tbRGifPf/UxRj87ACz7/BnUG6AAOwbEM8yG6v6FkmdqPB9N
4StFeKdKMf7jb9ewDn5Ln25hWhnXCp+ad0Mn7PtwIdS7wBlSRm1o5f52C4TtuJ9U
y3RgCQS+gzRNf+S5GjvS5LDdbol6NktrSk7lEOqZ9Ia72T+XyhrdG0OzzZFm5DDC
+MOR52MS+GGjNGc9JxG1gEH3npyszmM6nEMZd7Yh1BQTV4j5rfgrgoL2DiGuxyj/
XrMQ/8v0HyK6iaa6sx9+DlAc/vVxPFfFeccOufC24OUkDWSAi1kPp5zGTg8+rvlJ
UTK4/GLo/IqtlbUadCi+IPSp/jQUjMqw5rrpya9IGfi7/EKtRgRlt/u52stjYPIg
v9y+gpPZNAUTPR38spEnjFJh4ODphFtn6Uo7ErkGWD3ifvIEN/VCzChdneAAF9yB
/r80DgXij6v1kQM3XVzOvxsozTRxPzZUVmD/Ket3ai0T+sXOKUmye9WVH0qJCpfv
3kgCxNEPfbEIs+HhYGf0A+QQG2/sOYBN/Ry2hB6Li8BEC8AY5cmlmzwB/Y3QZo3Z
K0OBKWqchZMmA+kibx5czDGnQzcHItI1SaXUD1yhwXrrtSTnYiLXTMDoJivjIviS
F+WBkCYrK9IkKFcEdP2qeYDj+FqvmIs8YaVd+D8f5NM3TpCdh8HTExn7FN0XEvuU
erT5ebzEVHcnlF2tiMih9XglWfFhSSSWLB+ounQ2tLB3kn6WCLl/pOPjh7ESjCch
NuH17sXDTxKQSh1sTU6lDbh0ezro8hkbLgf9Ev19VDGoDiqC7hQ7MVD6wNh2VCN1
ASkuWUA5pv3Ap680rqP/yjIpXtrPXruNNEXZWOS3aUGLYsyzYhMxXi05KH3o45lw
BZVw0vTGIz24BLWvj4faNdmVYD+asCHdboyxuVKIxRn4LigrJiQToEQyaH2BL2Iu
ahOrJFr5uLhu5MfHGzjKEXPztNsAHQfS2YN8sxjB+WgkXoF/DHVPNP/psajznldP
8lAvDnvvgzFqU7z1V7AzMDdbPRMHiRzfn8JzEdI9aJKEZ+tdNJd+xVoRnGrh87oo
S14UnVMTin171VdjjMI6yoBjYZFQIJ+XZzKgUaSsddWJ3+G29Ms3xPMH8QcfSIif
09hACNZVY3iyyaBEPNcqFbMuutDWvRQzkEqmX+gg6U9A0i3Nsu50L7sicGgKnVuS
hAobTB2hkIOAboXLkpX8+n3bGSe2lRLJf8q24WC9MLbCGGKFyzlUFzgfWuADjXH4
e0CENP+EL1mRvAfQR7/9+N0/b/291GCRkQkCzlF61AwvzUZ1uJ48BvZsnxROKwPZ
C5X70+BS5UhF3CgGT882dbnfRvpyVcANXMZlR70ktncSCN29xM01N0BnH5htZ4a2
c6InPj3+W0RygDid4wRNIO+av37JquXQJPcPSgVrq4PeFjK76Bc0vinrlrfw+7lP
KszQE68QiyF6pDjsLYMj/JR0wPEp1P13Kf4x/2TWuiGjGQMmnFLDOTI3yEfAJGR1
Xz5qzjW3EqYx64O2/yIF4rr+4iq/y87Inki/MCl1xd9tHzldeVWc+3u2WbXZOWgl
YHB7Vr0uZfXo9B4GPpU6C/Sg7okCeK0zL77mYpwmhrzg+T7WMImFRghZvpOG45fn
qkC245hejHs+xUwMpHzcdbuHF6FNOiXZX55JvD/YG0nGf57yn2BOOcgxCvvZpFQ4
20Lv2pWOK3sqv4Ry4Bjf7fCrwboM41FIh3aebKehxNSoH+PtIfErB9y84N5J4lFW
BHUkz2ayxaNPJatROfroQsV5NN+yRTLcRumzFjdlQRtrUq5P5e6YQEB4JJxmG7/1
LwLmXz7hZPIbrUoR7YbsU5ednNU4g02j8Cf57qm0Nj6wlWpQz9Q3gpwL6wEE/L7i
+xeyo5wf1r0kilu8N0l7w/rqXDn1tVKNBuAMMB2B9PYwsyZym1rQhF2o/Dko3UAq
MYywMuezwc6lmyLrSaU/2Mk3bTQV/ER8onRrsMAyeojE65vYISI3KcWUJ+GFaM32
XVxM8vglZH5R1qyIBCNYi5kNsSow99aW3ZTPlj85hKks6DT6VNxsGoE7igmLwDa9
VoptwY5XFyUDvKjOaqXeVgNTFUaP56v4ziqtpZdpPkOvQyAKMEAEZcPisHYGq/js
sLRUpnEV/vXXiSUOXvqEg+nTNviEdoNwuWa1z2KTBa9ju7OcuYyDwS9tOXpRa3ub
nExjW/Y0i/Hoy31Fcu0BNXnrGNY0yAmRdvUG1opKGNba1AE1HWRUtMj0eg9xXjC4
LrTOqSavqwPQJBIQlBMKL6WB5rxznSRSesi4QJ2Id7CPcRgl4ta2oL9shbjDo1Sq
xY53c9RvqI2KzIslyPAm75Fi+tQyzud+KHdWOnJACi77qNGhzu5arLsLw8mkYEOo
X+uTPtOSEidO5bezH/qjlKrD3hsoASh+oQAoIoWYRqa5r8sknBNJrHbqtrDV20V7
DNnoym312IzjQTqwGRyoNmRQlhqZXl7eb6141mWyJR+Clo3pledFT3jqNNzvuSax
FfeUoRA3jXXYC6A8iyyT48zc8kRpUj5Ml8q2WavMN2CTKKIg5a8QqJFKkME8lI+X
nXpQ77vbHZUWUU6PQVOvNKpyPaid8IVQVkI2os+0tAvERNVispjDXAIK3y10Wdmp
N+V+i1Fd82eGUWpbpq+MYN0bDcVH5ZHDklZpTZ3E+oQcGqke5mtsVx8EQe7mZSXE
PSkufHP2aa4hN5pHkIrM8kTOAqCc2hr155dvd7JxlDJmCQAQWLyu1xM9mFGB9UGC
Rpyub9BkoGSBl4T00V6TWUcmnsO8y+y1upX0wTl7mA4R/GNj8ZC9k65egpNWugzZ
nIztqUBuV8oPFiGQUhX4ek+FXUjGX/cx/T6Aq+V33swLGezOll5CVpoidjWxFa9W
falXUryTIXL2JwT1WzfqbLrlVD0IKxvdHHIoAtajyrRgfXC8LqFdJ7PwfjVMHbeF
Jvpr++Wz3XIdbTAexcCqdmt9XI6gajzZik5+tm4F4EsVFUgzdYtnQZs9LrudxAzk
X/q3mvJzM9Zcq7EpXwrJSv17ZX2Al3OxM95IPjyoXawV5w49pByH4nw7xPkyCiQS
clS+Q24IoSkHTvN7v3TcQQHkQcPLyofkIfYl2WiLuHTrhA7LTqBbF/BSR3Z69pKG
jtDNitziiVu0UuwDfpDu09pibQfBHRa3fcYoREhdxVF/I3BQKY8nVgg6L4gqJ9Gj
YYJwRWbUba6b67WXcdtGFF0rDmoCh5Vv/a8Qt6efnGtFs5pcpChGH0Y+49Isl0AX
sC9oyptWqZ25G1MSb7AdwT/67qnyBbLk5VDCop6ERk+Uba5DhHsDFIFBmpz+9m55
FJ1M5fPekrt8l4ZF3HKkwpT2J0kRJvLnV/Vy3DVqySCJb06CU/6DSNalKMfccahh
w4pEaCjMRVtswFAxQJTSaFyfxR1CpaUSDfu23V2nA3Dbm6iyYlHY/HhD7R6ysyaN
d+j0VG/Fil2294aYKo/BcQLwqSSWRE6MDRPNIQaJ/HPfHhhtHs0MLEZNnOhFFaTJ
wsBqdtatWPLZSlKlLl9bg0C+JrqzON55TxJ2xgSMvbQbuKdHfL0RvdvzoKUB5P0e
688LvlCfg0LDQrGSRJ2HSZ5V5aiWSmJpypVRIgm6SA9QL7SuuCdf/SULKkoAUPAz
IYoRjbTqooNX5ofsci98FQ==
`pragma protect end_protected
