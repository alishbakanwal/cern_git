// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:27 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nXAGqzTtkR2Cmz4TrXk2xFAVn6PRC8lsbIzqEPJK/Av0jMCFzfOekiXFTBjHNFfr
NNmQLSHulzrmcKKOeXeUGT48cR6Pkm8zpFJQ9QTeqjkNgEkqD15Mk4pj1B+WMlt3
DtD3CKB02XocIWwyDlnP6LM+cP/x+lu0mbz6A047wBI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 49328)
zXaKRWqH7QUrZHDtNRbLIQrFD8+nuipmD1pQq15MR91VGi9GJT683/HOXSBfwJcl
q2e1cf+sONkIJ+fiK9Hr5F5AfampXuRT+IxUII2kuyw5UvuNB8hMycKN6PAhlXZE
lyc8S62h8I434XuPrSnK8ikmvAiD29FPufVt9WniUxeBXYvtiPA4BC/mPLcZ3EOa
YVQxWozpzQSPyUPBcYQyH5Mymi+Oehwk7yoza13djM9r0OHTXwEfsO+vUNleypDp
qdgmNE+1ZfzVnVMe56D7AwrWOlxUf8vJnqlrolgR5CMLTjVXto4T1h4z18DYi3BL
JbPdLBJXHQTeX84BceNJ3yWD/TYav/+1DD0PbgBsvZnw8VyXbYV82WaBb2WD2xoN
D4fX9gyJSVV8a3XXEDdejPsX3xHEVEqS9GyLn9goqMLwLiaC3PVNuXJzJtlxY/tl
2j7KCJE6eXqNfCVJA83CLQkhU3YtNCPVhAlpaBeVKVbY/L42EbFVPxHmvs65nGNc
bCIhRrKPyupLEB3cPxxmaQrO/q7JLGK8hPHOmDesD1fl9Ba7E18dkX46Sx4QUiDJ
QpqBxHF7NjjngOHl79916scKDSh5c0F84i95VfT8Jmp3jYQMqUGgoAjeD40AdRhH
Y246p8Rt0QS5/1HbksqfBwi9hnatininTfdlrqYZeMwd3DAMg6+nIOQNR4NnP60L
FFgYNwiMIlImkvMCm6eY0LWCOAxB/GckKWykRKRMJyFXq4k+rd37oryBVMDf3H/0
zfBAc1W2MBdvvZTFE9assrUL09EsWyFCggAwbQjrSDM5LjFuqyzetJ7zVeHw9dac
7EQusQHsdnQj6iG3GZXCeWMNbgf09SWioe2FvcfJGVr0Xd9QGY+dWS89jPTHSeD7
WI98pV4xLVIBxV3tMj7M1AG/309FyeUrGm8mIueu4hGt3gkW66g7r5Coavke2V5V
2sgSy7uI117/GCDq2eTi6lxDfwSV+F/JGRpix+ftNRfse+6/xldstGaTN4nKq6aC
fkTZWYf67wYbNIkGTd5So5cUnGuz6RvTJ0Sak9m7Fzx1aW140tIyVhWjM+ya109W
K4p1ZMyXWfkxtuFMfOefEZcJ2FoBuGTB+GJDkZfkn1171Qac0F7Lq4vwMYoZviLh
7z7ytBH5IqYPX8JL7n7nfPZvSz2LoQ0K7mn6OuiMHJffQO6YGSLqXH9PFFM7mVCJ
Yz3tCrGj2MwTJEA3sm4cb5sW6zgrc6lz34aJrKZpTtVAeYJuDqGe3lbWA0RiC7Rt
7o/Nb6fSVbsMfDSdwX+YiEZKW/b4VectVsAz0sjkCFyrejoYnSOHIdiyZhymeEuZ
Gzlr/g/LWY3qWC8GeNpbZTaH5Aij8Gmmv084HAm52aWytiLqcvfyL9xVU/RnqdIV
P34Dq8sWEh6ZxYmWDOgGvQ9+gWGL0p5GVs1mo/KEYHvoM0Suuuef9ibdHJV6/I4/
8lVqAvpDBS2B6rnGvaM/iwQHKZ+lnpUaKLp23aqDulDYpxak5roxOiyBvo7z2mU3
rSxUQ93W0+BdTDKVAGQ2O8jJi7BXvXCGM5YI+/Bk2WeQjPnW9ZEOyi4ugKbI1Hbp
8RVmuXkRSG9Qn60yzqP4o6zW5YG9XTBiPzKQQyuaC4jevqw/MJkunPW2bDCg3XmN
uD4i58WaAedug+fO3v8DNJxOKWudtcsY6iCl8l0NGZJywpvHAECmI6mbC/cGjSNk
Q5SvZTn8Ii4U7Dvj1IKYRlbEYj2c+BcXUFORHTXXYkU+K5GaIbvoPeJ5uElzywVk
ApKOrL3ZSFhKojeKjAuM57xX4o2VlHgAUPAMV1+otrOPoMG7vmF9kDT3lqwVmP77
E4NrSIEBj6KtYTRsRVza6JsNITG21Xhgu61BZXSNLWUUKGMdmbhHlQVA2SBsK0I+
cg0JQsOL9gm6u01ecRd6DU3umgcg2Ye+Qvr6Hi9/MAlXc2tgbyks+5Dqmjb0zEbs
wZfvjVno7Ec/myzG3ukA34+eePVEUnYS5xrP1zLSZ9Lg99M3xDIx4XjqjJqi6CmP
ETgbgBzSoOWYxxoYzoWNXfE3WCjqGO7FyL6VoOgOcz4kqQTXXGg4yzgJwW4kz6mX
IYHtZIjSObdWijSsbMiE/u/hzYzbNTXKUBG9Jy6PQFyFzh4V5HO/rw65WfCQrFaA
eF0WWmKPp2WG6SrO6FNy7tMuqax1RUlvnDXCuXI2aiOuta9nLt6xTLDesWxWZmcR
b+63lsrhzlzDhyj9QLg4EX4RJGHTvvvFEZncRnNs7jmKDaZ3YmOvIeb7Gem7rtwr
iZfYBmTgttYcwJE0toE5xbTKHFd1q0Kr5EifCoyuJR/bXg4no51Ml9Z93yfe1AFo
foOjgbOlWedxyGIDh3drujZZdvXmjwE0KxluqdjrTI+UqWQnHqV0Bg0FakwVpOhF
2YjdGJ8BImKtAGkr+2MKVPPnDjkz2mnF0iL0rP7bX7RxT6Tl8eevS50e0RlSV/VJ
/1+FhSozu0MS/qYlLh9Pkhp97QgQsIwVkMlil/iBnAth65NEIBcD80LWGws4E3vI
O1KBcU2eGIoc6pH+ho3XxO0jxDJIlmYT4GdRLhM31aWlLO6xMiTX4C1BJF3Ymwvf
TpQz7X7IFaSGsmaMQy7NIf5uRxeRHC5MvXcjAlwxC6OHM1LR9LKheBat+hm/6L1+
jgyXOPoMG3SrLwXbpxgikaLYBCu1yPKH35GDXk7dHwkuGDZv9RcF6aD3DI6nWU7b
RwDCpOTPYNxfXO9AmdjLQm3g/LwBJ1vH/rsjNk/0nHQu5oNhgYl2S/SFH283SkVd
EdJ5QT30FvHAoboAKlKQDjsahPng0OxXPd9SqcQiSWdQYHORNdA4eInPD1wQ/liR
Y7IO8Z6JtA8IlS6Lu5Ai40vll7qpEo60wyJVEeX6khhGoIYmVzP7r+sbCMbq05g0
DLhDxB6CbK03Q/s+Mxd6N1smbIzBJ9y6LsWNeLgdMROkFpt6kPufgyLim6M82cAM
kh0/G+DdQ/Bzlfx7qDo5nb67ZPuR4jMA8mvQ30CbWgSLK/uwUrV82f0bMp8uQooP
tC4KGDoJa3xDXUu3GXDigFqh1RncVnjz6ILEJYm79GkpsQDMyJHP7k0Lp7OZWQaE
8B3uSnKmIqQA19+mHMtN+uSRV0S3m7M5VwARNnG+tBkoPra6KPWbx5Ps6rL8xEN3
VAkA9axhl3KmpZGi1pS8ssjhUscBP0jFwg14noUw/EYDCGuJlVC90wH4Vfl3aR3a
BpSg5e5HUBziswJ3Yn7Om84wYRwBDJ662Kc2dzOOjW7+vPeehH0oHKwQBPQVHs+I
FQvggt6niFYptteGzYhYdGkUWNPdVl8o5ouy3yWjy60y1/rO7fHkzYjW76df/Udy
4T0hCNwsFO9DlywPmGXTiCk7nBAaQ3PjkRfx1rCyBAW312opGFKs2pQkOZFbNd83
A3GHJj4lhCIneNRwnqEuroRoYech6WwxsPuuQ1mQCUULVOsefCvKK6IDZurPiHe6
7qiXxB+198w+mq71sqF6vFRfywVF2BYR4SX7yDNArJmcYJ+KYtHmjAt1Vnlce1IG
OSbP6IO5RmB9X59bjGG7B9FG94xOlXvIGfZYPoJf9yhh1QYsP+LlyPuj6xPV2WY3
gSTLiw8ZkZSYKTVC+oH5SaD4sPbxYfrnjTTLoT9z2pL7K6Ef+BnDFBVr8G6WLa35
PlRjpLBH5P0imr7IEgRojLcPhYEfkUoIz8qhAophJfskN0O0laJGuKnaCwJcAco5
TIDBYp+RYpBo+XHRv9Jd5/Sc17VqOrFCVJssBiW9lsfp4l02H6ZPqT3CErNIM+6a
FZToCCKIJnAFXahPf8FwBzvG0xUZdC1nKrA6giasktyhXftZOkfpeGVKTsGlvmlQ
s8nSENMhDNuTQSpSbkIhpXOVUifweilKT2s9Ij6c8HDV4N3Gal6tS0I8DVKR4WJw
g3TJjho7ZAKbmIIfBngWT5UmU+zkaUm+09JQipePHyI39/IrRD92ZvG+LNSUMBUS
3TFTX51JBdb/bnftRTyY1WK/ZwggCfxWLDtE5J4Zp5ThfmLrvw/oiiPMaOMuMlZD
hNWvMCdLF5/KsT5CsqZmpzDbNgeWV3xYW2nAZCPperYsoeo101LwJtSR8gX3TL4x
3yg2j1lWjFl1cqk2Ejd4e/GLt/LbDxkQUbHoBfaPuEStUR3zboJDfHFIDnQQ327R
0tEwRYnhSVxaRXQaRh97FjgLPgtDMuwow4EfTFF0aSvEnkyOnNCd/4eMChBAS/Hs
l8Umh5knKR2Ppfp3g8WuADCpFMUAuGvS/ZgT3XQrVaPIYVnN/TfxpnIh0YfOzO+6
zqOzVAQbWA2U5mWjwzDFJ+m9K+1FNuixSdN3EF/x8UOnLCUYtG0UqpPBYF/gLhNf
5aOBt0Ib3q5ocroaZJh/1CauVSVhWN3VlIAKGynR7YvzM3uCLjNM1EROWGoeye+9
7DGeblG7wObM3NIBwM2OZJWNJkgU1imduoBs4vvAih+5OIqmTR9DBqtqiB5dPetA
P6j1EMl/y9qEE/sRZpli6uj9XHDGC2cnztmIYrxrmAFfZtBIkwRuus086WBUloiP
vKuyluA3OLfYiRGOwp9CxjirgSDUak2U0HShrvZMxBjfD07K3UDCritWLOvK6/rj
wRjmDSqv2zrfYSwD59N1zXhkKbVPu59UopraGBsirUE88suaGoxfActo7DdDAq8h
yrZbK7weBcbEjrDOB3OvGEagJUxwOvMpDbkklGZ1N5HZdi1oMgM1zu+WO+BLjZBn
E6d+upQcA7so0PVbP330vIZJDz97deBYNff+3QSq4RWaaPXaBjvCXEXZh6Zw2odi
XAYzgTfuaWsGrHHdkHZJozACWZ+408Zg5XjIPwLfwZrilK9ZQhH9hN6tojVIPhLW
u7h8ywVTsZkBgtPZ+xFZ538j0gYovYAqm3T56+FliV9K2QuaIBdY9LDUqJVNxmkx
fSpE6+SdBaVqhK3WEZOqa8dw+zNhizVJHiczzz76XVtsiSneTbjc/828nKW7HOpH
DUjslKiEmMjFmSZ6v+ipNcDY2HaOfFqxoWGOTWjcl9/hKOwFAnVVaUsLA52G1qg7
udCZspXKax17W+C2fbcLBFNF0Y4WUBCD3GcNBHo9zAiZyW3nAqU19/Zg5IELYmfV
EI6Urxq+NtC3z7ebiAku2oN91gSU1frWb9yFGjyhVbyElxAHQBB/fUS7JPqFgQWl
oaTARg+1/t0fBuK0G2M1Z0KhAO6LI/FzC7U0CcZ3gR/glw09mV7cBXuPDVtuj9nu
/01BGDLs12J/Ighho09gb5Wx3TfCKisnOFbZTWJN2lVr8v93a+Eic7Ijh5hB2Ty9
tozDrEMRrWE60nBPLawuDjpWyQ556I2dAsOjDMo2h0+KMu2MdvMj4UdG4Enk+P5n
7cGDKMLgiriKYe7qqdJJjY4RWJ/NXZnjaTSQ+6b8VWQWxPZQQZlB4w7GVOlm7+bp
QL4g0nXeKdbsxfp4MlvbGCBH9mnGWkrlY2XF7YS3HEvp+KuZbHZ0Jx4G6udddCcF
Y+Ef16sdJKQFuyxdUCdyB8Jz5Li8TXKf1IO0Uxa9PFWfkOlJd1B+e1s6kAVeeu4b
WNOEasHhpVEufAb/cZeynyzn2/nphPSKchOjnZzHwBjE+j3BTZVHyLu3ZwB7a5mU
/V06kiAVzgL6hEI0ACkpwhrorJnOpEkLaQE6neBhj3j14YV7DOAbAi4GbYQoTuE0
mMHR87emAq9Q1GLJg70wIjodwg6HDmAASsddCTIsSQa+XjR+vPevETmCCsVSCSJR
AriNAmSNCxhza1K1ZxPZezSnHl+quPw0bAmzCbnLKx4db9wCTLisi03HDJMcg7m3
eCMAnHmInqAmOJKRn/eJcl/dcBaLByO48yaLseLtn+Sn7W3fBeIbOVIhlaImhvuZ
KPT7thsQN68VXvUvhfO7qK6Uzyf/WAuNQfsjWNBtzdQo/fNQr/qBjpgMIJ1ZcU/N
WNKrpnUgETZJhxdhakuYVvZKIfUZZw25akD1/dsDUeCnuZ3QI5muMHzHwcWItzZH
qlE7821AWVx2E6VPrVsr45t2rqiFYeJrLMsah29LhhnI/U/TMXCKve+Or0P418Ai
zOKFFtcw8i/4cQ0mpfTLAcPNq7LGlwfMLvY5XfJu7hXattVuEH/7RjCOLaUyX2F5
5rMpyzeIMhmbfY/vPmUKAmLRVsDxdOQwR2TYARcr+mvlR9+DlUNzULqhsnDrIJOb
QTOyZ4vgXv6Tjp2aoVJjvZ+YUJK9uHtvzvv5TyMUcpAxbdIyxS+q4DdjUEGUZqmr
LFEzRT1wJ4sVGoaZBU/onz8IZ8E5HwnEjxLBGzFXnyhB2xo/BxaBTtnvs1HkGDRM
vwOj3iQaRB50vUIr/l0FIolVoiO5b3fgGYWxE/rIWEuXZiD4ADCA8tuzBEz3rybO
T+u8aD43vaXf9etioj+YQIWC+5sztF1G31Ntdzed/FHDKeujrsvTy2aB2b3K2wh+
UIkWxtSU4J8hYEgDac4lpAoDP3tb/hMvcX2Q+vJ44t4Te33M9iNkB/O8wAtpp07i
oYbYVrzFsy8MWA5sBxW4P5KGWpJmK6uI5I4ojEz8iYlUkXdNhg/R4wVkJaMDpkvM
kpO5AAxFNIHrLr/cDAHA9wfeCuu8faWEyFRmdJ6fxa+bgDrINVu4jFFtUUoPNUHk
CXvzSg1+sGC6EUajyo25fcsDdw0WAbTuqXUKeiNZT2YX6D05xZ2MdRZN8oPHVAk+
CVKmHk2KL24Y46VLbBUrZUC5ly+01S8kxZ9yefPLdcOBP0G7JiSk2Fs4huvtg1L/
fasD+SlLYpgBZYXDLaXlRnX3q11/iI3hv0pKyCjiOL+6+2PhdJvKseG5BAXaTfzK
PRFXieL7nCuZzlZHA6u1nQMYJwNHgTCGqN8KbI79os/SHx2kdIG1RI32TyMJ8dBp
mIAVdPnW/JI8PNWjk/RduKQace/uk0JbzkYmjWOJVLYc7Z4F5iQirW3tXzy5lKbP
Z9ifuBGboVPMNRksJ/F1R2t+2tZr/RUpBGL4W+gOHUpieZYHfx4B0eWRuG0wGh1u
RlQtjd7HMFgbbBxWSS45U5TWREn6/bf92QGAWmeQBhxQk6uC1aMjPkEWMNYwF71Q
mehHQiNjzs5h1yrWUMaFb4U0r7qOUkFCogUbm0xsCNsFtlkE4KW72qA3EO78Z5gK
Ujrv7s9BwvPxAIRFH/oM/7ZKyA0Ra5VNlAUs2DbzgbimktqmCZhvmet+7duG3g9P
3SYtKK1Y7ivop6AdHhUn1wvNQWKSWlxJ7h4oUOTYgrzOtytoIhm07DX+R2+S3Fd9
7KAmX+4J2zQulhzB63o9elRpxbyQDkMg4vnQWBoxN3HisH/M0BVosQvJbHeaMlGH
mKmUroFT9dmj9ONxeUzoECdglOkRyV9HiCmRrsq8AKdOl/B2DhS5slCtlDU8U7+M
CvmsLyMY1/TWKXB+a3JY3hTg0Mxq2wAYGw+MrMRlLY+SWcewbrbWiXH/kQ5PAdLy
j+upqMq4gPlKwqE5dQViJmYMB3gwPlDse9x+KsojdfNO2QudG+GOFD/mA+tMepDS
5GsUdw/H0n6MMNjINoA5TjlOSzy5z3JQPpJH/lwrTwvOCPm4rBYvTWwPSNaV412h
3NcbULiGyYUYLoOHtlYm9aY2fpfou7L3pownjgWotTVVdcnS+IwnkETGfqk6UcSm
Iu+1djzlxp2NWc0t0s1VmesJtKEQcMXN1nsikXF8Yxo3ejHUPsMZ6x9zvKGfrShD
/07iNcIqk31QFjl/JfbZSg5MrzGFVDcbpQIcH/0r8O8ay+7TbPR+h5uBlO2YTuYu
4NxJ9XHIXlCt6QPeY8hnVlNIncbRSF/LyMDGjZnPJ1YZZlezvtUbBia2COpR4S5m
3gZTHS4XZpbGKNqMxMhX2ogD1ew0jUROh5hUkEWkC5tx7svuZiIKdQBIu4EaIFcM
TzWhAr4FQaHfgIwiGG8n1FEDMnPSic3u7orBGrUzcuOi8DvT2Kic2vQbzDeHEk4U
2VzHKI8RQheXHjsUyWcfazhv5YE1DM8ZeuIFIKSh+7NNfgPm9WfMvtxxMOYVbxQp
5rc/pEYRzHdfjPKWmacb0QYrRFtIVGpySP4lmUpSQ9od2SnkKC+5p1uSRMeq4WH3
24PFfJ59o4Ns5gLAh6A7datQdiaFDItGXzWergFkdQdpGwHfAiN2daWJXFAzNXGy
V9e0W5X2TLdvvSPQDrKwDlrKfAJp0sN+yeh72s1FcDW1AmNhn1CIWPjgFjbsQuIw
+587M6SPcmJJ62LTytyI09R8gWoE7cZvoaxHdlimVho+d+IUw/CB3DJ4pT0rYN0p
ABowl96vPGlyEPMbTYPE1BzAq793XrIkT6+FAGT7QOJqeS5xkrLcHycXxzKE9R5G
sNP/zQ+FRB9fNZU4FT6Q5n0a3YacT7LRPkUUDiJ0U7vIwkOLNldpHI6IH1eW87cG
Fcu+g/WBTRlZ0mF1Bqlyvue7qQmh52NFfUz4VccGZdODeR6mW4tH1Yr+jLBqQqRG
8wOcLBhafkwZ+TCbHx21CWHW7oyPow7SitY3MS+E/jvqYv+bNHWVFBZPcJea/VoD
oKRUGIF69sx7qG1uYV0RyeATOgyfxYXWO+JfK2zZRn0xXp9ZLrHdpxQs/rn0HbKN
olAqq7cLr41MDMbcYfRrGx+zKIUjGgsGzKwFNlvNahxJjRZNyf5c8elwS83XRz/3
uKFGdajHI7JwYy5ufsvBW2s/RY7BTR7oHIRdb8OlYn/KpcGWcOp+Mjba1OhKnGdO
C6/LwHrJnh47ahY4iVDdlu2lr60QILWm4OWyyb9QzREeXrFYDt+MQui+gkrpjZcf
8+M0ap+IAATPDha1KeyTwTN7SkCxDqzYh+dRhM+8HezEWWP+Td0YwpUkJAMXHmVe
unJFJz2SCcLqMpj1CIJ8Bsmcv/wOo4TIVMJ2iuJY1ijhr1fvUuDGz/NVdBPb7Wq7
Yk3FtNohPGckrn8ejVy14EsN0AOj/Q1L6JmIQdrJcKnrVA7EqgFws4jvxN4AqDyT
BEtpZ6AVyIypWt364Zz4wztsql/ChbcccF6nDjLQSZPoz2Cn6If14H0wu4EfaJDL
ga6QzpULkA8HTF7RCB6iIDDErATMHqPF2T2T6snDlcdjmmMLnVKaybgpVzZPnWHt
/wfRk16wGffTmfWPgQz1W5c3gfIuZztNlvwN3Bxm/0sv1stlJ57Fq7NHs8fKg5td
SKMmxEOfz0JhGwBZukKtEWSPoWbDwfhIF9Tko3Rr8QWLPtbosStnMmRr4XIwVscA
M+Gt8snLEb/n3a68NTGUD7JIGrgBDFzy0dco0wWBH1DKVJt5VDjMt0PK3JvtQOmR
iUFvv8TDFWGbqvPbYVBUnBOBChydJmuUukylefnPluyamMmjXM7UxQKqIU6JW2AR
vZG8ggnK9sHKolyQv7x9bktREnHRrMzY4Xo5twy11ZddqxBu4OtKz/Up00hPNhGj
Cv9TBvUqK7qtzAvttWGKT9cK4D6wv5vjufuHxDKOOu+d1te3VW5dCT5DKnGOHMX1
QnEIKu3ZSsgeu4OvEgeoYqkHSROvIuKfJ/UyCK+uKdR7cWDLgsAmHBIXcOllei43
3eiU5U4KXLunVY5fPJj6LkAh+2eGcYja+KBBnBuiArQKrrpPZvyJCNZGqz7uSGLw
nkdM8UR7MbC8dn4eMp4N1OUcTnqDtBBJN45Nlj8MvqPAgbqJLR0gXzQkcAkR5s55
najCJ2cbYZjnt3sYOJH33toM8JbZ5B1jInJvnawruy1Yw4RH8g/uwZIKH9shXE/M
gopq2WQFljnFGPuv1KH022JSX2B4yYQ8G2WP6GBz4lJfpnZCKjwpAC9s3ri1yZ4g
rW8nqxPu30kODzfyyGnylB1uRRGXHxbQIn0X1Eb2P2YlXVDSRIvJJi7vokiatfES
QzT68dtfQnZ1i4mbFvVV7qD47oJq5r96cmmAVMqahKrJVK/KPOloFmtHgg9wuK3s
9D+ULHxuw7pHnQDWEwShpbG43uE4gPu8W+lHrU4BCCgvcpocL/xbQBeGKU4JdZeH
E20SuQtDoH8v3PHHs9qT7ra3GQLHp/kbatYNoG5/HW4RK3DJRJKwGMrsSUBh6Ixh
SGtp7EnQmCYmeYjFWIv2hVSvraIgbun9KVaQowFWjslxWNBl5w2Yrh6DlPDtxJ5q
KCDuPsKCU6uk+TkihptMZl3dccwUClbmvEuL96yicN9xUAXyddYY9HdITh/IHqF5
wF/ozR3Yc/OP/QkTb4712pkHoyUc/wP1/NEYkjbFfjiHm4701C5eIPlb5ULQJFcF
WwvDF5awzVV1D16ZJ5SHZ5QEpl0Ozo0Wh+BTyO2qYkQbfUB5Dj/xAQQlzY1yv+PO
lwFxCLp40QErbV+y9RO1gicz4MXq51VOgIZ423V8+boIuPeUQ6yIAjlX1echQR4q
HvFUT5a92DVrnvctF3k2cbtB6Z7tFA9Eo5wZgVYquMLIr0545d5RfmYmgn22fJgh
zwU2ASQshErU+HEaXMozmS9aotSydWTibuSVtXL81URLcyDqLggffnVVEgYooMKX
e2/e5RcynuiYu8xYtf3ac6eh2bPBk0aNtIisMdxDlOHMQqI0eGOto2LFf3sT/2lh
pO8WuErtF5qEneNJQDXeHFP4H53xGpHEs4QR7EhvAjniuUXV7LAErtAW7stL4u+y
MlHne2AUF1la86wIQWUCF1R3fKVpwOpq+QQpflsGFkd4aHqVQ/AtA+pzmMf7duiz
XL7KzLuVWnDS3WGkAYWBa8+MgDSEaHHjykTQhHdGKd5eU2dIck1kLyzMFLIbqHPS
ZK9ta5jpLLukpwVXOzcFfbXQnJyabJJ+yIzpdpPl8FkZf2T5U1DpVf3YpYiEUlrr
/yLn87Y832nVR0sZL0+q3GWVezmKGFN/Hy0Zr+cyehguPZK+i9V5pOAljAEgXbsz
cuC1WZuvtpzU/iff6XUzX4ozfcaD/usLsPs9gn42pfya0r/fRJ1+2pJW2sPOTMFR
s7rU+ytMLL8CUcYKIOP4xcZWxIJcnmFKP8RTHho1Mj22MZm+VhJUyYhPnoziN7JG
B/5CK5b0e6gO5CuUXzX3aYlhjpiYr8XYLGuk53GOXvs3ZYU1lb8WM5UErDu9tK6O
IChu/bE0Pp7fbrVnwmrBgJ9riSBNL4oKFUSrtB64LN70IuUGxTNs3tnFpu3ywFLj
i4S/72kAsaTpfjvYntW0Hq6shL8AOI7uXHJ8Ix4w1DxP1UCGz2gbOw3JS45fiQgd
xLVE2SLZ7/s0JozGQEDMmuExyCFyJ5eFiTYPOHeoU0JKaPFNdGtq0Ap/71jfhnxh
BZ/UZxOMpV6Kvsi+4osIrW6tKdFeaaQSw8rIerVA6p0F0yENTHwOxuoHMxTDlTLA
E7K1xSeJBkZXu6YLPkaGi25LaNNgZCy+rYLqfWIW2yEkUTg0ZpdesiR0hYyTAkUs
knbgqPjvOx8rdyVgFDwY1ns8lhXsWSjZohjBUbYqLvjl/7H50WCpXQQP6inujDlC
xqP+PzO9qV0Zrqu2qCSS0cxv/Y3b61SOeygj+PWg1Hg43U7D02ye7k5iRX2zQmlz
CyMg5ZDEKEFOJmzXRFXcJorDw9O+ZIKPCuz+33TAgLhNEcLPzH4KgujxvJ59hmeN
5uB1uOan/4ZaS3YNjeAfYTV4T6/q5GSl4vrrO2U7hFZpb8uYfmuLc5t6CFb3zqgk
QG4GoxgvwFLdZALH//xmYpUsTnF1fnvU2n2WvF5vhd9U5+YGMW70zXqKj7XSmWD6
BtoOglXDfKKfBhE9yF9wNGFMUHyg3ZJaWS4F+FHgOiYFkJNfbe11YNd5VA6ZiKVm
7dVuRKcswMLlJw7ogefWVhJE9i2If0/kBYt7nGs60b+oaO0AjIExWgqxld0rVAct
YIkfzfMUXN1ugLeFATr+a6A3szbarswnKL8dQvgLGHdxpQAfeqZTgmwWKOC0R3Hh
9c3Fl6geQU4XZaUPEm0DuOl/7nvzawJ4+RXvE9Vbd3Rp5RR7z1ooqivAgDYnP2Rr
MRBADV88Ixb0Grk/kR1grIivbkd4m9wE9f/KimsfgSGV5s8TbLvGnO418sAUtfM7
on0ZtxmcEHgxabuQktG70dUyZDOXty0oee+bmvUqOkr0KNbYa4/lsKeiJy1AXgAn
TpfH17utNEm3YmCD4zWnCPeTge6hZs0z0N9g/mbFk1ABBOW4Ph0j6UQZ4SK3YeBK
gjDMN0vu5Jy+edlE4lX9TRa/gmo8akq+kUzSU+cFvSRqEQetUeKpeGao+ZnEc+Sn
NIyjjwOg78RPW4P+VbRXWqHJA9MeAQzth07SRlUkFuc4C7iYgfeIK1t5Z/CgbIsL
YmjXtBjJhA/H1R0YRPGXm5gqhhyAHTLOcI1YoZDgvDRh5FEegpKH6Sw0oZSqclXB
7EZf1quJRt1xod+Qeh54FHGy/K3p5yWN+ioKTM+KYV1Q0ET33ZyEzzBtpxqJSoKb
Q2DPAj5sgiU9jcgPI7yPWCruH2VRubuV3pDqILFVRvNnnaXJfOajWS661DWhrbKE
nYlXbMT1AAALJXfzhE+qiWlufeMlIpaNJW2wmyiHqOAvyMQ21rjGk5A0NS8Z2lss
1dAOBuBPKw6RAEPfk6fD9unzT7NkFTpetpRg1qLswXAr34akwJOszxaftUfejoej
TLQQO6P6NCxXcNpPg/0b0vyt/biJEhB5Cd8v3COviGuwiwygyNN8/4X30VlbnHcy
p3p/66TLnKPmmEX6hqK/IrIqRb3HID5DtYgkilez9uJ6vMSmGLqRq4aulV+yWE/S
2RFbxjS6FEuGPpdbWoYQ+hd9tpLyA5zOAaaPd9HRYfrfE/fCYp/f22c1vzmj7EVh
f+9tHBOZnRgX5tnABteVe0YIldYN5ivH8KG8NHZYZRXQoHSJyAWj4pNAqBqMjPxx
4032eZFLA9cO+ZosTkEIrPu0PjNVj9+5Bhw8CJGxJh4BcPN7vMHN0eMZiHbqQFmA
PFh4FaJDQ3XfHmLyH4+K7Ut1V+1l0lBqzD7qiPu9ze/xlxHYSz+QSXfAJMjbWE9M
k8S60vicQrdJl1U1ODcnlpfenKcj+Giv3ka52Ukmx9SafBWY+ze/IrQ7AqrBxpbV
CK0nFkjyL539qNduwGN9q09hYW5tgl3NwA8V0yaM8Fc2dh6yJRzuMkgwsfGP6Aik
DA6iYUrVUIhpTayrwL5u1vxRRWRRK9aO2ggiqjDPZah/bga0TLhZGlgJimJLxtH5
NroLVyIq2A7/Y7i6/RAoyr4mjzaTa8UtfFBt8ys6Tp7tAsHVHp0rpw0NDTT8QqwS
rw8w73hKRZ65N/wdYMvlTBm41vQNzNEt6XJQV4/o5ExKvKUh02iJap30Aq4YZKmX
onIhV0T7g6Jm8CjndYjw0gHyASXsH8xxCw7i5NgzH/UyLnZIymjtopczRI411OhY
uTd5sq1/WGNkuIQKvTM8WQU5dJc+0VKCLWFlrdlfgi1RH7tZ12/PtSA36ajObe6q
wfDTuEGZuReYzyCTyYADscpMg9EbyFRk3VQbmj7WeIoxC5M17eyncvOVIhw8HbM/
OxZ4/CdYo9P6in+hfDiG5LH/4TCj3AEW6Jq+t5UqFhGArrPQMsugMY1UcRhoHWIt
8QW2IdBMIoWQqUbg9RhoiZqGkea+0K+gUc05/BPeQ77VW8gSiCkwfXx3GpgItBjO
tPywAx5tUQclYaBcflJmmXXobG8+OsfYgGwjdNlSlMhHqCgXpniQDtH8PVmzqGDN
UhcZs5bVf7hzh4rpK7d0sP+l4O6HzNPvsSSK/l6X6219gYjMC8/eH+InR5owQwgU
PQ9bHP26uw7s38mietkHRTkfMfgPS3AMq4CBMTTvdd/xW6RfUiKCfqAK/XSZt5ZB
ffjm3s5rYmRoISISEiDF23j0YlU6dLDqdJrJsKKX8UfO58ImTvL0yXyT9/yTycAo
IaA7wJBV4MqHf/fTMNMztxbox3nPRqRSV3/awSmUZ/CTvOyQWNuH70VVM3e/SCr9
y/mhM7IZF6Avf8via5djGM7K2+/dBU9cvxXaBBjmy9lxXoeo8DDns0qckxFSNVpA
2W8BMWGPq6WPaVU594/+D6KZX0J7jE59o29uozuDGJMXIH9RvXkcXMStOwkMYJYe
P0Hy72e9bKjC72ZUab2XRjHW6lVPTHyHOCw34JTl6YGDOotxLS2zk8fMFh/PkT7F
CUu64+WleCFEhDM3bNh4sM9CREbHq6gCbwm6dDMj18O/Y6phkt8HkMlOATjy1nxR
xgEd2fKlOO/8JI/fgBOHgseHyoH0hfIoHfE/j9n5Y8ukm3cAXNmo+9PD8cn1TNdx
TfoexUUgBg9sR5wjRdHeBXxKBW/KfLlKFfGn5GcDb3B79FoNUMzTYsUUFl6IZOvO
hN4Fldj8+4RvpmxoQTmn5pDte9q+L9j6KpeL/Hi78YEW+JJ48yCMRYZHmkwAXoG9
4pG0sBtDOWpt7fmnp7DHbcYWLm4qE4v/2k742I0E6apAH3UuFto1rN04MfZmputN
QpNRD3vh/pd1Q3NcAYfZHXdLBC6ilkhAbGTHcUbPJoRpeR03i/U2awrw8ogCz3Ti
Nz0et0vpkRN7ODbebtHIRtWhVCtlgdj/3IDpXUEm3Vp3nlR3Hzecs/6zQAqk8410
pUnorin2Jcwzpgj89pnK6vLYOdqZeMe8fPN7SO3VCvdegX/dJrIrfRR4F2nI8uQx
hP/hC1sSaMoXV8ld3YTF8HTkNGaVwaQuYBZ6aDiZ2wndfmg3e2dKFOo261+yPG/6
KhfG7aRM/lGVM+1EnMLu9AdnzqgC454vcwFSNyO7x/NZ8bsuyfns0EyR6OH0CyLu
69XRU2MiMsh54NNecKy19T33hYaCRI9HlVFYrJjh6/hCX87XkiHn+3lJZT17abpw
gRFPYuf7ePU2MBIhIll/BNzgyu0CBVyapHXlPdcv7L/t4T1vOoL3idZtnwZQDtQy
qrakRugKob9NhjiLC9iiKKddX1zapQUPGvGmpalD1tOTMWz7zZUOyNszIvjI0Jhc
U4hOJodilbzureM4fZXFhg4U2l1OKK4wzey1A8gBQXKd0wf8EOZ9g8CgI1EADn9L
r/Asfm9LYKTUSH5P+Swpg8tWqnIvK6b58qiPsRS3Oszhv6/pNn054jyADvFNWRN5
Vjnnmux1oinl9xa1+4QW5z7GOqYRrrYhaHzvizP4GdeJEm51cuboYT3pqceRd9c5
ONgh0aEOaWf3seoXfQxH6PS7twQfEAGgiMzu5b0PuwotGyrIowVPq/rZ6pKMiA/e
cm1aKUdhyxLztEbM6CpWMBl157jFdlz4SThYpT0Xmb0RL6OOmc742ArTvlJnTLfw
5OonLID9eNcfnHLYjH1TFRMNk2TJ4ZqiJoazMemqPAdbpl9nxdyN6pwPkOYu+G6g
Wvp8Tk9qCogqLru8xMajvRJljg26HBgRmVZL52IlXv9pdhOSUHyjBmWFfepqrRC4
ugGVnFKHTWQEr5+qq8+0AjA74e7m++XiTQ8dvN9QAgpK++phG9XltO4aakh6jBr7
CRiEYX54igouerNgMKGvEnZL4GACMvxi+JtcUHL9wSN8u+6bk5tWj30QPxc3ck8f
7Gf1vjaA+a1+jHm4hj/OnTsm31ARFsUne3cZqq4Gel2bNSrlG0DJTvZ8xFbVPTMt
7NNF1OGE3D9F61941ZfnrQ9qDLLQO6fV8imawOuMrH5L1SYbnnmY/ANEOkI6Iej6
2G+b6ylBP9A1Rl6HzJ9vu+J/M4ZW5Epj1JDYSQ7rA85R0Ba8vXiop4/l8ksT/Fm+
5unZqnDqdR7GK67CrLDcuPPviwUp7RjuUIHEDvsbKwRrVrXju2bN6Gj/tW0YLf8i
KS+s9zEhjG2dhGc1j8Qmgk3y8bpis7cjM9/LCP6Lo3GUX4NJ7sVu77ww0Zow4qJo
y/K1UB219kUMRycTVnewpj6VlBu3mG7iKo2diEGI8E0yFoY+wnYlyikJMW28fV49
Le5a8jICP6JHdENuOBJpXjWre2IXZGPfJFaiCvrcDI4BjiOcSrg0MTFN37yYv/h6
Zj4PKY0cugs2mHoRWH+6bORbjXAm3qfGEjEpY9s2szfTVN8PXxg9XqlVBGClKTnR
5tLKbmZS+4ab9O39Ayd+qUVMNdokoxIkcbhWwNJ5fSGNBaTl1zL6OQVNrTm2+iJo
JU9ELmzFWkbh5hzuARQOsCDM8Z/NUCqdKvyt9C2tuvYjTQ8aUrIdcdk0rOoiDK1s
uApJl5MLN6JiUhEWOl4VlUNjceqNrHyY7L74SY57fkwGjBmAFTkHuvrN10M8/skg
RiMloJJZ7FEfq5Wjhrz98LyRm8UihmBXc6tjojww4WmFwnBnw2653W2cDItFf8KQ
Fltfv5MmSlGh6rbVMI97HHnpN5DH8EHJwc22sfB7Hu+2nhPMq8cs+feOZZxYUlei
xDrWvETCw4An/yM6CI3ITWchJbF4YFUk0joE6KSI3VzqIGvc9ZGDsj1tNq3/GnBZ
j9fqx3ycETg7akzvIolj4ybZCcS5fy3rx6B+1XnlTLHAkMKzebulyXN87btpjaJS
Vn5SmJwxYw5QZxq1Q9j5NaPBuYHmBRI0xWBRJIjcXMtI1ZqW7z6Vm2DigSUKSC/q
9qpidpZHSjF8pUy5ozk8kGAGO19eZHcnp/YhdK0KwLuuLOVTDV38/O3m9fVVKHcq
S1syk6e2oaAbrtWm3c/PPOZUF9UZUjeV2kM3Kavo6gRxgSpwWWWdquE9u1fwzsj9
GcbtqCYWtL1BNGmiNBAkSxGQliWbMCXoLypgo/MdXvI0re712t+R1J7NVkrSwxSB
0CSJ+EHIwxbfrrRBa2ABQgUE/+/34ClyVbaY5iztjF9cUKppjOD/A3IFOmyQ4PLw
ro9k1s2W1Fzzchcw+GhSb14t2/59e5/8gaPG/B0OMYZinHXAlJvzg7QBuj10Jnbe
QileCbSHhklBC/yTQLXVnayz79mS6VhwhJRqzrD7ZZTOZNJ/2+X1ZqTSY5kXHhKY
c50FRu+RRlYNvq+Ey8ZH3PDsZq4R5WcJODJ5QhS36u7MxVlPSe7LBGsN0JNteEPw
XIBlLeyR6aRumGe3O7eLLfFRuYB49L1tEJrIPNldI57ttF+3cBntj2f4uykYYxc8
w1+QS9NjaWq6NIcSDNHiJwAcUUarI2jJyQSAIuhavFr1t0Wnhl9M+W8UvFYmmlgK
yHNzl1QpL9yFaT6ARr6kkahK5sMX1GoGwiFPot8X0NNRcUxMpKs5fp5ck8kUDDIs
vDS7cjBrG5bHyMrwZICoGs0RdemY36XzVh+kIdd+NdydTGKykapLN/cTRJYMVyoP
RNZbQRnh6pBqcdhWlSg4fg7h8ni5QaI9bVIyrfo1SAUfDtUMRfBQURP+r9t8j+94
KgJLeuzP1ZqRxSiNEELCgyrrwYsINDVOUIDUKJT6BZGjDqRh5YGDFyXscwIUArqa
ljA6C7eUEQ6U+2DRfwwuBPIpcW5jc3GuJoO1DmvfSZe9SlpUdRc5QkzQi30Pjz0K
cURSajMAVGx7ix8ATkNyVhJ8m+wRtab4Z0aIKdWS6Ylbww49ui66a6TnoQJxU5NW
GSupXizHXO2gJkEmOHtqopycrPFpnKCRzY1Ky12XM5+PsG0Jp6btE9BGXlxMvK6f
LzWg04VeG/4P29TF0Xm8qDO4Sn6WD7hZbt5vxpJ9FwdFBBdrMSnSyJGvqX7m2lge
NZ+daOCj/5/17TlvawMVBOOwA2t2l3DGxlv63L/dQZC+YIdW3bKFGRzvElNiNeRl
6nJSVw42UTm+B3yb0qF+IqU4ZjcepsKoL4+YR6cubae+HLX099T1wkZvpVdTOc0A
gkK21H4WF1Kvi5jC0btKSY91OGefDFIZS5jUM2+Vsb84OckmC03d4sb1np5nQEIJ
MPRT36kwNmK9k4+LvzLy4TOF3Jc6ZQj34ZGk1PMHjsH64kwnWRghq623HYaJA6Rp
itGYduQI5iW+P47EqQvhsuGykCSb8sGWn54EYYxyEdkFiKhauIVNmypGoiZNlVf/
BDygakQkkEjX5dDn9MVAoT5CsKhCIzDKgreab+TQPXpOUbgGrzNWIwHohAZKj71D
7uRK9l3UwLnpJqdHyckfAXedmIKMkuXKb1WlERu1tHp9ZHFimXwnbU77VxQZX5Ix
vDDOh7CV4omM77cj41OI22VH753GW4HtWm/MDl98p3XKGZTT4X1cBsk8JVCDO5tD
+NfxvAvmPAx37wNyBhQu7Z3GMQoxLNB3ce1pgLYATfwl9xA8tH3NjBljyNrTmP8c
0dnfnFXzGzttw5GoUv9b0ALZhJZbVkXFCSHkWa8hidPWTS1Dmv/sR5UaluRcAWr4
05n3NX1ILZSEusJ1uXwqfrmtpb2gOIewFHUaO/3Mn+OA4tJnpl354b4Up47p9BY7
zynVZ8NG/Nqb/DR1RWS39J4RW1l1tkgl5PlF2elXZ8DD/zJlPt7cg4InCXCqjF/e
rnQ4GSJ5CJZbVWMRxnRA8qtg45+v0fwH5XT0uPnECfmfV2678RlcHcnkT4tN8hQY
ExuVCPIpwzz98nPFFG1UQahgP0E45taxgJ1zk4wrUqqOk9Tl7AHjN+/YknvwqpfA
FrjH38sSso6fQb4wqBEkqsANbGJldf8FS9cZQXnUXHSQWTy1wZZHySRk7rn/3yyA
YCAXJg0qGoreCn+4UsbZ4Nm6S6Zx3vMuZRnGoO7rtz2youGgbzFx+pxyJnzfkPml
xhYouubPxk44NMN5ERKKUJr3ENK6wFGyCXCVmMtpIciX079z6KSkIf2GZykXFek9
Bsv3HmRtN7bfIl/K2fYmoMQhosPwnSV1gyf7S0eaQG2Ol3cxI5TOqhfvohDi6UXR
LtvoD9jw+K/FgOQ3gWCjZ23iEAFvsCrlZ19spMuXOHxnVhMxTabxNzElaNoExf/T
6o70Jflhc/PvncqKKe0oKi4u9jVaGDbmnIrgc2t9K/53+j7nXQx7+gRniVUrM1Cv
HtkCn1vwxag/sLLPzLMSPP9XLMuEiZHk9AXOKb4Nd1MjAGy2q4AGbqeQi6va/EBZ
5CB8qkDXqGTB/CCr7WRLiNvjrBnv14Tp9YcziBP3CoGui1VBdYZrMxil+pbAQgsb
CU3A4DbX6/Ti+xv2zleqCgBHbqQBwjbhE6OVOMmV87bH6GWYeZzxIoskTHw4+bSm
enZ9oTA3p3sTY+sWo3RklpVIgZsFp1Cat8vwJPl0B7HjSwu6QTV1fZXmQCyHvg9R
FXybwzsoySjvim9W6QAGfy6BQm/CoRS3sfZvrll68pPzLO20FbshvnyWbckhSJiv
9J3JO9pMX6iCKVCOk40IuXQwURqkl2iXtwIGXMgiNp7nSPcsivAnX94N1ZydtLlC
Vdf4RiViluo1hE/lHbnf3LodsxrCF+mcQ6VmXnuhn42kwJPP3uiB0vCw9Ypu2JDM
yL0WF7cTtT7Ks/eYqx/iVcOsjBuszi0pGO2gz+sN9hwjUPX07wMBdBYreBeF211E
UJrNf+x74I3l16YFJfEkRcl/+gJn2rmb+izgIKFGifAybW3tdUEQK/nwQiRbL7Tu
FKVzUv4/TfQAC9X2J+aMtN04jMMVkdD+9VoS/qtwhlh+CM5eu1MBTlDhutgvRkI2
AgQM+FzLIw1DsD4G6stJ+TlI0yldPHhwj4l9J4H4IBURnDfMwQirhFXWMS3HmC4r
02nVk/ksaAwAj2QAKXmQtt9NKquhEZQ5xl2ftg01pqe0oaMyzbK4sY3z1WWmrLs+
iJlmR13mIVdy4fluvg+N3bujWBBbqG2cdsQYACW8cH298xWcU7HQ1cXw4ogfdYHM
zG7VBhZQYv7wRpHPKVRqCUZod28S4ukb/u3zXIl7Hured1O1/1u3ROxSGjWIAMF8
QrTcROkAHEaU1IOTSmpxy/BQAqFrz4NOwfyngNp/OMOCD8ejNmSqkL7WKP8cZ9s8
bylHtUQlJjyD2hbtLmbTIGtH1wN4FB3mK/OFeiYZcF8pkck2etS12zU0Ip6pCj7m
6B6VdKB4SGh+hRHQ4Vw2NUy1C8uID1Hve/Mld6EeMqwlFTWtvcXoudQYex49uxLa
G8qgggTd1qVoMLKkpOSdQU5tBNmbAKW3KzVUeEn4LNqc3/7/WIgFX4EIR3zHuHuN
c1Yc2DvXxyqX0TnkWcdAjVljjSjq+/HYDJmomw6MBxNUcVNtlaIK0X5SzoUYxKNO
CWq1JI3VcmLxHvDccSccQGtjkul0DUP1eajbdU9dwQuRKt6d9c5Ulhk4kqk2u/yq
ZSZug3QjLfdqUSMA7O5QM5IhZC81DeYFoqaDgONiv1gzMKRe9aotbujDC5Foz6dx
mEXoJ4KL61flaZ6U/vKGABp+P8fMQQH4daTzSXPLj+yAABfVZkcqTccBaaEErCVU
OrI8qXzzVoQ4+Sw0q2CUqU54ZZIvmyToB/kWAGfS0wJj+InIbgfwozK6BrNwl3Aw
gJjswuuWwoimQCPY6051NVdYk9OqcF7jhY8F6dEvHE2rQ336gy4cBZzVesio/eR/
3XbRTDBH/0z8IQ6nN9KVfpLTdxdOI27+sP/rPtI+Hse6ZVvcpYJaCWPzaYWvGgkJ
/F3n/42/izYHGFE5lD41FUP3ANaErdmVK9sGFkPdeSrM+SLjuJhcJIlNJY2i4B85
i4KJ9byXDEJenukroew2meT2scU/oEysVbo7ltFfguHKStlCR2nQgu76vTcwihNN
0t4NYd/dtqhS8nztgb3XaieZzYjnNYQVqmKcmXVmrOm+DCZYeqIASPc4LUxIeVq6
skO7VRdPn8XYSsOGwWylljH65/FvLB1SdJEpSF/ML7GH0mlXoCjupgtv6BocXTNB
z3Fn8zHrnt2M2j3mq7GOkmHf3EzxHF17WroFGiRy5Hqq99LzngpvGBTXKLhfz87O
vDFN7vdK4rdtfQqR96U35it5AAHELJxpTN7sKRcCaS6QYzeM42oXBBTSOfkF5Hc5
iKFU3F8vhTNcREjaepKwMOZjhtBT4/aCUDZZH2sGVyO0p0tWR0DnDhJpa/AcDoIb
8ndKHc1Q3QtY+w8JMSvBAPxha7gt7U8QU2u2/w/2ssiL8cZMVFgBjwEc3+o5sNoI
Z0ML3nodlKsAiY5G0r4wQ4EdO90vRm3RAcbLqvLd0nS2mwRHM9hWdIhNDD7G4/wp
oWPPRBKAFQN0lBjs3hyObENzsZTo81uDdLsQuspVEtWa47k82MrK6VTNhxEEoLcj
tp0DxFX5TlJzoLdyi8L6Mi2kLWAJE+y4mk5CcV8YV/oLN7Y40Wc8lqLxq5UmOK4f
P1g/QfO8xlUQufNW8JLjrpEMkjJ2z+smC+xw13r+Y531HQsjiYZmPKxvLomRga+h
4L9M7bXebnRGXtFV0UcwZ3/hfHi+2rQ4e3A7F7SMq00mUjr0sW5nhf4upDrQYxzi
aea27NwJpx3rJltpclp0EfjeuCTaPorTAZMKBpaMd2chYdIVSVBk7+YSzwnqf0pD
lmSTLRTKftF3DA8qlcf4GmSKjHd2UNyJ1o7ecTjRjTYqXUpsXu7ck+EBWtxEvEbl
OMX3t+KXjJIHBIaJMhk1NeRu45oEU/VEok4O6qWy2fn86cWUk779pLmy08VnDXsi
ipQrMMd300kd798cFY8mlNJsUJnwkzLr80xs/dBu4cc5jDdlYzWH30tI0veWvPBb
p8hTMz1eJ/Mh8Y2SZfAjkEjbCGh9xbOzfs3Oc7TmiXWwgCnQ/R9+el7r3VxOo/ei
u6nZc9nZP002BafP5jt1v7IbhRpjsuCrR+Bp8LvY0iKNFTdpYMHrHEpj8MYv/F2v
oMCMO3ze4KMa9aNkg1CGbjnXzfetckkdf27e3nRu9G7usizXjn+nNfEWU1lHjh/s
w4QPQUrO2nzsBj+CtDiduuovSFLUOdM2nosK/YiIoNKrtAy6YnvnVDBBWsndvjQh
1GW60yBctErDUec1EfmK7mBPEd/4BWLn30WMh/yoRvzFcdub9ZIB/fH5HGaggfga
kGN+ICJh3SSne1ESMO8f5ee+Ne0UNijlkwjezTTjum8bNArwvf4/4ukFxm7WObOe
gFjOliL3qfTS+SZXXnSti9925aYnsdeelhBBM9YH6wyvmgdBoAQFMKE+pef4Wa75
70m17vHNGFzA4xp8xhkkkr+Lv8NR8vYhps1Xj2etuqvEISXjQu2eNcUBo8seXIUJ
TBKRpUCMAKC8/7vR96LHmLtggQtRMwQw5FedO4gvz+fMFgdJx/AXDFuMJuOf9UCt
PLdhqX9uz6B5lHKCxNgmRXZLI/2D2oIwGYyX3tyov8TBlwmW60Xu4cUxX3BfHyig
lo0ZWDQ/EQEsuvZfl96nadGsJecfKQB5Rdy7o/j3DN95pie/hq3XA4BoiEf/63jK
RzlvS+SkUVX6Oa+JQqXIlZ5+EhiBVH3ociizbGRn5MHMlAByuZoiPVIqXLHXDFWc
GK68mtJMbmxDhlJRSAdZNC8KZgJtmPqL63CMLKQ9TJ3rlqYbpoIdNOreQk6Jab4+
53maVvce/tR5zHu1rc7G+88ei+9lKfDRh0tSzi/r/48ahPTuB0L+IY7jUZ3aHQQT
722EIB2sADhNFHiwEobPw1R5yKY2UMBtAhf961s/yxIfkgj5rWjgkdTTZw9HoBv7
LpoojDymarHyR2tLvGPCVP1a1KIFQSvjxN9F0cX8tnXfzQBNL9QMjzu1k/npZde8
SA1tMHtF6l8KvsQcihcAeDHfplyxx/5EZoBwZcRx82BBj+Q3lk2mkJFKpYZG7BTp
+67tC3Sn4Eg9MRau4YM4o4R9CbTat9c0nqph7QelkcOU2GHWv06XWaluq0N4quyo
RWcW6zHPGnJOCQoisz/yRmKTt0K3SsnB0ODs8zR7oP6dU0YEPgAUV6XQ4t7n/wif
4/X3xOCtq7wzfwtX8c1L3vpxnUhtT6qza3xNaIdqC1ElME45o1OOKJBF8r4v6ytL
bcubeV0EIAEnAz+D8/H8ijq70r2jJrZZq7P5gJOfyvfKC1PQHcAcm5HKk/j/+PR8
spyUpXt8KzowWwhj6Q1baAi4/8MyBsH5MbqI50u3nJ30lBHgyPqyx+Z8759q3VHi
O55kI4vJz4IpoqNv+hG8OoVPAyKLOFV34aQ4YArKd4WOYg0RAZv+Hmwbd5MC0VJZ
OrbS/SrB2c4tnbWkDNmTMxOGwambbe24UgGjmRKbowP/W5n9ukP3YiEUOhgwBAc5
IFeMIM1sOTIUcI/yxnQC+fnOyTjfY7HHkX+ua5YSZVWiFpO0z3NgJVuog2GpMXd5
ExO2YAsozBbfK6jisjOj6XTYYOwpHcMzn7sTpGrfaggANcuBO2FUhf68VFTRjQcT
kb71udI7Wbwuakd17LuBe929atJI6gTCxOfnKvPR10pqLi93jKUKmVhdAiXzK4WU
5fZ+WRibXoPXD8dukoz3AF19WYHPROJk6g52XQB4+Qy6AH3APGNAp4kGCZKJKP+o
ZmLRlRiH5Y3BzB2h7JBUGMXJ9ADyuG8MBSqP3cgSZPiz/acJeIt0txH6U4b/SNQh
SRa6hCJIMI7rAoLKguSCyM7Pp75YtXD1KWD3UNBa3CelUvrz48B+HNxcInEC0RQb
cyhrNQ+kATpbwWGjTHsWwEPoU1R54cnGeNhzgJlItWTHM52OuXmhwLjKttwTvSpX
VHPWmRADZv1mzIhi0ES9J0lI2ycqNKGHJianUETzNtS5S8jw0voieMIdlt2QZABA
nKpY2dldRbPLBXCZQZtd1DyMZbPqQBOWuHggGPN2zTZ6KsO7kto8SrqVigjy9LOv
CzGL1m2DJJtzmRx5nXc6Z4+LsZOpdrQAHbdy2rCBMg5WMqSKmmZdngNcfZRhd+jy
myn1fgOLElpibmaJTfMUrMHgBeJhNSQS/24N10BPDHjslf9fZw+O4Iut85xR7OD7
mSKej2BObSc5dk4rBgFzrP010q7ZSvXK84Q43B/kUnj5duIfR/v4pvzbs7p6/PVL
6qNYWadj2u4sUA1LtgGPeY5iAHAVBnoyRgdNRIL27KhmKBrHFl9Z2hSAhwNC25Sm
Iv6BjEO35DoSX0UWUxHkwH97fTs14vM3PYR9SPfoPWFluZYN+IovDAeh1eOQIkkn
hompRVy2TGeXPIHKW0Sm2PsBEY8tZWgxP3NTscfsP6FGduONOTecAuWKx4uPwRgS
FLDfTT09w4NlpHE59rhkME4Qv4JYnWeP1aYt3HkVO4sehviX+YVX7JiPKTdZLCMv
jCblv29aiZAoMZvk7AJq93FOHndFf+YOw0+FWpPFpNyoauE/nTm/qfB/0mG2lmO9
fCB1/QvJu1XkoukHn4DfQBWeNnHCSViB7ZWB0zEH/nApK3c4UScGU+l7bidFJPqn
5FeV8jSD7OPz28wnicnX5LdXUBeJ7litXHo+wat0Fn+acA+0l8IYDmbyv5U0SSkV
8IWU5B+p+YxG3bLpzIGucGwtwYnCkgGXGcVtja7GF0Zw67beq4qU0NURLLuDsJ5/
1Iu3GqYBYtDpEmbPv5aDwdAsDilZFbJCxgWs0Q21/7xn/ngw3Kvv2WYWjGePG1w1
hGxeHw7wsJgtQc9J+AxfKyyg6sh1uS8GCmLPuoAGfk16Mne0NAGbQLkyqOX4lem/
s8pEv6FHcus0B+f1z3/rgNg/pTVA0n7xpIN6w0+8utQ6zmgvPPT7jRStMtmGP4/J
o8GNazW+tTi7H2EZesPEPhfLK5unRPvave2ZwPPUu3xVP3D4PR044g1xZ3H952Yd
LcsvtU7DXzddEhpfTkln0iyHWhNsUbmw3Sq26quzANNi4c4tbHFzxlrY1KVXhD1d
vKYMrpVcOAGMc7X2nrc9QbplgAJiTlQT4X9i7Mr0njPpOnZLC6xb+pzYmPEla3X7
HJWFA/t4vBbCbuDFyWOGG4LAX9Rb5y4J+l+6nSwC2XA2jHZoeTpilWaMSQ/Rs5qx
amoCF8sWnrP44pga4RxBHmuuD6xQ5IOIfJC6MdpXppKRStyA7tP2Fk5WK5lLjzHV
tQNhxkbLnUa0SjvNY0sZHIQJZfsJC1huhUbSWOGWUv/PHntG2tH6RuroGFOZeSTF
5XxtebEkCaYY/nAsnfxNr5PYcKJs7h6yEl9vJi6fmDvgMUPKs87W9tkP6kklZnsH
OTMM1m/h/JeL85jS6PcQ5ZTi9pODzudDGJwd2hE++d0SgzBwCrsuwm+34FmIlrt/
r5450s715NuuOCkiEddCFbdwTcReAyJXfqlVtcUSgM2mqHvpl7EJb5u08uYIH755
0BU/DsD0dY1fD1TyM6lv1P9sg/xJcOv7RpNas6jbOMGnrLbOrK57nIhU5N3fBDYw
6/PjqS8g1ntDHZzynty1szFv3Gegdx1wAeegojzdqXC3wt6xFuOvjdWkHX0zWJyb
67l51iIqaeC6UkEt9gj8hhNUnQjM5tyiHNOLrDlc9Lvd9QtWSu7f3f29MeGWhLla
b5zLwjLeDlKzxtHAZm63Td9aV3g7BOcYjh90daiPIeGG6W4zce1RUV2ObiXl7uZm
qD9KiCGuH1hNeHKKyj8E2Po0DxTU2glZXDEQl36bqFu0+c6j8Vc/RaVq10CeqF9V
nXDlbSrt4N0BUYCDCLL5I9aV3BmxD7yab8vzMQ0Vouj+WoPqGrpmRb1+hrjxOG9a
HrpnBs2M5+s6Gb6tzxuFIDeWbxl0sHjSJa6LmTMmF3uVlYsdsNFa2BT0oBIr58HF
X06C96zt6i/VzuzbmJ5tbDrxxq/BnV+Q4UUtzIdIssknIRLrIM1Zv7oxj1QNT910
S+te6tIVi7BaBav98Iru4aeKAaUYLb0OuUV/2ggsuOAEh5FwE7Fl5P7beerkuk6f
HDXbKtn09G7UVMHkUF2+PdpqpNqmIQemCiWBD4fm8o9aqTgZwjMw4eF3Suu40iIo
lBcUPyhZ/VEkJl+UZ8oz2FRwB5Y6SuHXmCsAzl02ew8QipXJA4P1saPEBP1myZ6H
tTimuEqF+VA5WM9UBwRtsYKehk7Xc9r4BVS2IGcwKPsIuNXSwWNK2YzcvXv6LIXE
yPhdEvmV86k10Oes2rIM8EM2gibKwTCZ08Q0+NuKKbcnRczX3BdRP+hm9ay0Yt2M
E8uZYwFMVU2mPC8gApY/rYpL/0ZFvz3HNhuhLvUlh3RTHz9ThwXPH0VL38O8K05s
SY5PQIHFncUuLj51lw2OwJ5s25U7y928U9jGpija9VQibJo9aIFBCEmfxqDqtMqT
5VVZGnhH6P0pqJBED9ILJj0Uxng5/CbxsCu/FnyHj422OEkJiK58boU2rfzBmR/a
p9NPI7EXBhfx+x8a6IDOdfbuEhkTR/EHL3Rg3QmSMLVU2MUYSZnD/XCZUlmzBypz
K6vIYHpga9DMtu7S7o//byPHBkd6286RE/ri1xJaG2mZfnTl4kNzw+88MXev5rbr
cMc/SmAhqlOecZmQpMJmy7aMz3XjN2DIGlgIc3MGpfPhKp5eHEoka8BzeoAd9xqP
8rVKy36KyU/xOw71LHlJd5w2utXTTxexyWOdvEK42EcqDph35UM5XRl5Q6uysCJt
dt+olUKg3aQCBqrHtqfIPr+GNJ+foApHgeIeZuX5baphxdj3UVdy4sif13G6IsSy
PvcWBI5MaH0QGfDYHp/qjZ1QM7JR6BhckBReSJogoUKc9jT5M/dLMQI7Zf3Xxdn1
nC8AFCh+luM5Lg/C/rYWJZnrvt9OvGmZ539s6phDYK4b3wLQhZXBf2h1RXr8IjzY
QPtNjEg+OZoVaQOSKRV/MnOivXEOkF0jvDSsjz9vQMRd71w7/T4GDiX3TF98kBQ7
Qfn+Z8IsQgr9bk+T1sWzUr9SRvB3o6FCbfW2wVciXaJ+YWLLs2cYAVglLlAWNWL5
Tqtt0Sd5bUVch8z3VlOL9JkO9OmmFThzuP8LXSe7ZScISzA7h+jeHIErQbLCd26F
90N3qJZ+FaqqIxiD8nnjm+drmyIAgvmhYW82zbj3F5/u5GFeXFNXVtsJzff6xhiH
deOTyzVohNqUASDa3g0/RsuVPTmxA8B4pav+2qRLKyJcEMnXxOZUagv/BqFvd92I
2UdmiIK2+eDr6kaf2yAMssvJ5Bak+aYcsvuZ48rSWkmVFDXHk+9YdXWxeC7A8gCf
WE6WazV9/sZ16GftSmTDxvFACYIs4/OKAU6HNzlsgGl9akakcaLLmzis5ClPaJ9r
6X6D5z+25Pyj/cwvx7sjg87mXJJ8B228ZRHBES2FDsQ4YtWOnIvcelbdtkUj1rNV
92D1Ozj7hyS/fcCwq1mX/3wFQqpQN6AHyhuUgG1/Yk7hoTPAF0T3EakRQNxJX85l
n8aFWNQ5Y9J1uojArdynBJE4/g3OKW7v/VrPpFhVi2MfMPajyFNopCG2Jgq3m4JH
aTKDCekq0JTVHsNXpMxKY6kpC/70aj4aAtlNGbMaKzACJNer2jQ7OnIgWzua1Ra6
y6p5v6HAyeo4zQBK2ZK8sSnHNye7KrDw+YqtUBkAuLxQ7W6UyxWOUNNa97fodSCn
TYvv4SG+NsvfBnZfgj49po7JQTzwUqciXxOLwGP8CuGCFlABwudKR/udqm4xEili
H4tSkskSwnfRFaEH2DRPUDky5FBXb8LfJ51MowlxlDXwTrYKtqdxn3OYtXixsc25
1vQwSmS2ApwbPWAbVGjS32fxxbI1OC6ZY1ugQWgVgZxhoc5MdKgjaDMnCAiY2ipu
rBZw6cPl7B+Kw+UJF+ySXbBcdl8AQqWMVlGAX2j3pZubsKulgkNM0ISSYCNMSFtV
Yhz1gw65agfz+hg6IVz5m6xlYO0ZScU1zX5pM04ygmevEpY08w5/H+/HQqRtWHWm
Bvu0/qS1UTirUpQ82w1fCof3I8KX9K6kuNNJNwz1lMUQJQOBjED3M/C+dsh4B+pg
FsnQS9MbhbzgrtjRzRN4XCfv3tIzXmIUGpVZxhsYj9aXNnaZzuazhYHbWEM3JZYX
VN0Y0bLFCLfHg8XbGXFM2S+DebqykUItO9gMIsZ/Ol3+qjYaD2Sc2H+wGY5/9Ax7
1i8rZBSuuW5EHMJ4BZ3tt0LywJgld+dV9wfTqQ5myNr13oDdqPtAobqJv0J0ni2D
pd7XXx/r+Zi937F2GBnoardsouwyu8sxXCHB15tw/Jzdf/M0jp6Pv6qmasV5d0ta
HId8G5j/Tu8OKKQpvPYNwTEWmt4GGxzHRPY/QqAchBfa1YYJPzX1t6+KgOuwss8V
fWBJVRl2XmaB7d6KVxZTVFPU2Oq2z3JsEwSRjipFPyqfQnX1cm2ZOsVUKAgQ+O1s
tlfOpTC9gdpUbtm6AvJLiVHc6dGKkG6Xr/Pr7X8Aiz3mIMQirxU1ddIueUgyb5qQ
Bn3+l8QiRPEvIpvtI/PDGxWzdwhZNkzfqLbyJ19Jyfos5M74R75y6sGi13L6kKiJ
k3q0CxZxE6vfwbi8Q8iggNghYLtj7SsLmzFZsEOTWJPmAn3RZt2GzAktGDd8MHK6
UudGRNDS+ae0ielu1tZ8P6JsOku5/UEapsMfgvHT/cNtb4JH32a7qCrWOdWbnHJa
XuAkbYq62uXUgGBE0G1/OjnQYkSgXF3q94QHyUxPtGEKp+ljUjQtfY1iXq/KZE1A
r/2iahiiGM49GP9zSUXxgDEAxwQDIeCZMbXHHDAU3IAlnMFjJb/ZBPFwZj1Xc7Qs
ppl9aITjCCQ7BUvcCmqWt4qcM77+HJQ7B3bFplvLXseuAJLz/dwRSH8BPkzRbYU1
9plGfJLvhrfvlGIYUUvx9+zqVlq/WBqynJM16M58436/V1hjJmhLBM7IyLHrnh4z
EPwGiZfxLtmAr5EMyTxjpUMPjx5Sk+y1ceJEZgnM4g1O6GutoAvnI4mN4XgVJZ4w
edr4TiLEaQB6zGjGabEZjKMLQax64Yu3Kp2epoH/Cyf/O3hCy31GKxsl8pcqr/KG
OwudyrC996gk6/q8djOx/kNkitcgP47LITWe/Zd5SecxQS7E7ir3c4MKjxGHFO7A
Hr9JpcwcjiIddUiQTFLeA83I7+D35pElbAsVX3WRBqcNP3ElAu+ORjeO8zH64Vkf
Do80QNql22R1yUPLr2q9O61WVF//c6lh7eQTphXiNUX3a8P9PLntDjYPnZaPf0JF
+u0fSyZI0EyjsoCwOxVDqyCjhz+aVhoJ1J2wxJG/MAhKeEoGOXh8yFEkcvCPCtzA
TDWQfTjuNCQukRJr+yZudFo9it7pYTprh5w3Q+V8bT7ZmDI+kMB+PgcA5nm/tFEh
3C+CSLDOOJG+B4ioghAHlk6Afj8ZQBj1bah/ETmLT/EU5Iq9zHcExM9DLUucr+Uc
zIwbEt2WLSoMKNGlT6LKRHSvo7spKc1VZZHDYlhZe3MtklXkqAzleSKxYKeT4wcb
4YWu0aWBSNSSGRGMKWIDkaHQr0LlncCDBfcBzCdSGJ37RVjepKIZOyNuLbwNumIJ
8qTZMWkkD9iLV4PihqQ1Ghm7bo+vsGAXHskHscQT0DajxzJPCY4x0Txf9E/Sy/Qk
8QjfNCfi+FMiEfUcRxgP3rJGtkzPrnQGbPMu51nnGTjU0oa6ThmVuKqbfNMWrgBO
cRgxWQ8pqy0W7y6hebWfrtrHCyRF9ijEM/tiT371Ph7aWsakl75ahAwGVXX9NwIB
wciV9Meofdu2RTqkNHHR30AzUNnElelxpInPQTy6whz7BMRcvmeoHfZRvYg41HQ7
mkzs66ckODaWSAwt4+9qWMXZMgUj2afoHr9FEiIFYeRJgfk5ybf+pG4BFO2lpIYV
V1GgwlSmBwhShty+sjOes3GwP+LjpGQFiry5+ZZJSL/oYnp8unA0uwqjQAYmJESe
yufvdA2OEK1AnwJNOFmYjWflvn54rHpMzrSoVNUuZkRpwEzwRZlorrnEHBqMtLO9
rOdMNGXM4udJCMTb170Ps6pT9IqLvupZStaykw1uuSL2HY3s3e84RYIYJmx996jO
pBXOrs3oSP9VJuXnulKZ7te/nU4+tmL0nQ+Z9Gp8w/362S+lMjxICv5NfFJR/jky
DBTkxZqZP9W4ONowdZk7IXkjAVB/udnrG2IdZ6QdNPsE5lB3Oc07DgNxvMWUXEha
Ox1TlhYtSR2azNtfzCywxRK3uqBlcW4eaUmXuesDujagrdpaxo9AUhtvUDex/aE2
9x3UGW66a9dATU9ZME53kWPDYz4ST/EIELhscsUlvi4sqB6EnTSwev8RrE7JKKu8
sKtjaCK/4KDAmljLp9zsT7rd80rYRsQCeJJg9s/VN/N2zKxXh+vweB6EoVme//m/
B96Ezu7usJx/p0l+n+1MCYSfKUTILX2gXPq8fqsbcUWHBgWyyMglP0H4nYLxhuX1
0ejUmykNl/uAbFWC9umR4giaEb4T48VNp0o4KT4q6rF/li/rH7v7Yl2SpkYi4MCu
07WDiofKxxLQ4rQkZ3txYKCQO85BPZ2zW0alzOQlCQbtzbUJzem2X6xDcYk/SWuf
kt4sCR54VTYR4lfJXx3erQck2MnY+iCp6IFNI4QwXVtYjnmaxrbALo0hW/4Vb/5s
W5dA98EPpLfE45uea6Qp7WoVhRAgxnc2YnnCT0SOuY91W3r336Adk1FOT8c5/o0a
7Z7HouW+MbSNazkE1Jy2hd5Pt4gLSqtK40kgKCHH26vPB23qMlFwuZb8i38xQJPP
GH99hzGWdTj8PmHln++JpHFnFcTz9GGBIwOfQ6NaU1bhVfxRCeSbAcEp2H3fd7Vc
35dJ+SeKUgJGFVnPP28NNEUdWejXgs8ARTuJ5bF7Td1fkxjMBe/GNa/vZrHKvyy5
lSRecRpW+a+lQhDskNKqOy8EkY9+ilHYglmPJeRpM17dwcjIa8NJg1I/Iy/gb46I
pBmNbfrmbpQT784ivg8NMsax5xHOCp04Er9D2O86Dy8B21r5VSF0qb9v3bUWpKWs
zlzxZYNMzns39FDNSkj4ynRXKane78D7om3y+rmSZ/iKiDBCVx1e7IR7UZrg9Cxt
1JeffmYTRQIZM2PzU7HUkV9gkBAb/ETsfNK8WExy3gOF/ARBZ7DgWW6Ok5YWqxV2
B9MKqGDl2B4dgnFxQNK9RAG5nuVla/A9R5uylA25/d9MVrD9AwdeU5XTx2I80uLo
xwXNI8J66aKzig51PhBTZ6NAsrjggaNt7e7qnMof1p5fA5esShtA9IkrJVPQxZ0B
xwxCdX1ps57zeOvr8zsrsvmO9+MLm455GoJpezfZURarkWbhRHO2m8joMx4xHwU/
HqBPil3Wv6kkoPntkxbH2G8Zq0JFT4w8QK4WDn4fz5PEdrM/Iu8Iewe1+ZM7cCUs
g/2yVpcRqNlxLWgomjb8DIYXJbLaPnmc1ClCo9KSqAiXkHwYSuOHdGX+Hubs3ssb
aJI5EC3uqywwQyQ2XrCZ61iHgeNyXq3IIWpExBqPeY5hvlvNZAkIrOvil6tUeDuz
gwt6mE13wXojgZK4JNYOVubvxe+GQgl6yXsWYXYFs18Pd6eV9pJjW+xrCtEXi95c
Jc5YbQ52n3sZ/tk64wQNKvMHHPC9nbLXgcpZJq207T+qhqO1I4Ri+Xe4s1MVyZL5
eEppD2C4hbySbwSC7zjTs/cB9CJ0SkD5aA7yr+BRF1KN8jB76PMUSDKSDO2BjJN9
cKUg0bnwCnVr6iA3JmTBS6hGc/96Q9YMmToyXlwTiIgL8iZsh3dyqCC9xe7a9ZGl
AoCPEVK4Jd7vcbQy8gUMcye6k/6ttYXv9DMalxVxxKxAyYn5rcOJjPNqJZBulp9j
v+GumOhKdvxLazMyVAAc6NAX0KdlAQ+DjIz9D2rfuMnAyHGiCjpCHDFagpne5PmJ
O3qUKZhUbmHi/YaQT+XqH1BejDljDaeDCcOASmaHCoGBIQHYXNctM/FmpAiCZmRB
36nuKz+z1kTvKIZiTW/9eeZvQ74coIxo9ud+ODzatTkH0T42L8/MfkvIh2QMdYyP
M+t8vjH+ZIKU+JGXjvfmiCBiqhCBOCq1WaaCNp8L+ZLTCbAPTgBjNWb5vV/I86TG
bwd5kcBo3ixIsAE85WoJmQx8qeb3OmZtW2hTWvNgfmZ869ZkGdT+wD4/vqq5vexX
DKNoq5NWVpJrexgvGsjgiI2Rpm3f7rgJzoAf7+a2druU1OBjORtVA3g46B2vUccP
A2djuryNvPGIRhEy9UHF0z/rSbYXkvpUICA6sLR3Zer2n1mC0DgAB/zudKPbb82+
YPu9LcOvRxKsv79W034Pnwk4hWf9bJxCINRsqkvG7lePOI6HVzzfDDlmDpEYeraK
XzH9QgXHVotb02MyIlBAd8J+GYtylq2n8p8q0JD7MoxNJDMviO1TZqMo7p+6pFVt
A1J1F1JDf3ReN628uZ54g06HC/0O8KL/ZjZ4wapYQdKaxeli2mhcBMDwECbiz076
Y9KgRLZsMniRX3Fy29swNl98aR3EhSoGKFZHLC+Xe9LpgMh+WTy6125TEtdKWvJ7
dWve3QUSFzmCZD0OVLjTr/MFwr4XkaRaa69zo3sLFcgMrkjHRT62Q1FpNRfSovmL
cuCNIzDozeSzqzu0tRpvrjyKNx2vFyTLWdC/ulD6Nnt27R/dst3ESQnui1QQO2Z3
bDWlPBg72zRKJaaS9i8ujMJIH1a+2XosjzTnyywH32VSIbXVRr4Ss2hT41IiHzlg
zAcM6Jpco2IvG7YSKMn5Ex1tnvzdBmUxlA+yrSzrgU/YS8JJ6ZR4xnsROvEwG6/Q
E5zow0toQVOYoxGhYC1/0UIMS3aKMXeGlX1rLYSsx2+FAIdCowgNIwkNvzzK6RZv
YmvJ16jJyLfpNh8JUn5EQ3/NcI0uyoDChTRT6xixOeljNreEE5HquHdV5TIWENw+
u/hG10BL9Aj+3zcCUxchjBNl97nFpAv3kBptfMqGsk6s3svVlyYWTd9FxXlhcfOx
QATTHk1IJxPJKuOgfG42PJB9B4ugfk1TbEngI/Q+IBiYtzZCx8H6CCdgts7EEto7
4nbWbuksXFpza7m1MrELw5NdNOAbMmgm+p4rnwuYg+BvEJG6k5dZBOUKGf1xI8va
H2JKytB1SNYHWVf75SPieZv2cIUfzGCQ7RLE/JfP+NxkNzZ/nyC03o1Ul2+32DR9
WDIy1h/9i460RWuk76+rzLWy7lyh114Ho6TzFtniNHIY/EYfg1S8tiD2vw5zPAHf
XwV2rLwhh1u4HljGC8dWbU+Mo+YtmgHrywTGzBURusBQkbFBc8n7VJ+kgw73uD13
Y6DrdiSveGJJi9zOQiaFRfd8EUbIfVIv5L2tnLk4HXPRTszF44SYaBUtMGriPehO
C7+5D8Slh/pe0jOGQ/7TTVxTXQ0cA7HE9y1+KkvTK4wy+Hl5eE8q11Y+XyefoVNN
BimYH2ejZBDszC6sSRBJOZyfDkTre9oWM1WVJY8kkyRbju6AnkCas0nWxD68tdJB
0y8ic50aCzz7gFkIrojlE1JDHJE7qkUMzg4R5F1CeDCK8QcdnHhIEVLQEaa0ZZHD
WHXF+5U+W3Ox76L9AGwpxashexC99thOGcR6BS8p2iSYRgzPZuMJT4P+NtizI+lt
0rpBBu2TgC292GNBYGsJnwQUt9EPud7ezuvYzwGS99RdcTaCfEKXZ+M42YJjxvGP
5TI4Ostab0fkx2LWukKv2v/bPAn41CFhS27og1nHB9AjhL+z/7XGUUVXBcKQvkyy
TwAFlnS5zQ0sl1T3pvfIQ+OvHvBmL0foyEBpjMMSr2mJLmGnfBMF9FS7YjCwaKOM
xDw5kqOzwPQOt0CHDKYNg64phf1+tN6wYwszrvzyX6mPcKIcAcHVqcQQ1JHq9Sr5
vX2+rsxIIYtSwyj1IcRw2MHsutGKQDfcLvWFYCzgfzgRm9CnOcSSnPSdxz6A8jeY
RZWbrVqvSbEoluctZ52bWKIrW8YD2KpqE96jZ7SWztzMQZFxKBT6K1EGNVK2GBWH
ClFaKt+RNFw2el6BB7Fvpu2IlQUdinx07xBDCQBAQ/BW0+Cf4pJJ8wNDUwcFPjkp
6hEUxRZKaYdrFcq+nRHDPapd4T1aSbS06dKO8XvHSrYlOQLjHsEyTqyyIV+6NvS0
Frq/VqC9hYn291cvhqx8rjC3q/Lz7XKhY3DMF3RLrWAW5av4x9KEAKNtSpk3v5Cl
1XK9JWbgVi7AFjw0JKO0B94iuJifBFDAxKf7cWc3i1ht7GOAAXKG4tip59tW9yLv
dTbimnMd6UQkoIyPSnfVSJrYxePc6BUQcmdjYtyVem4QzGHgPZ4TWtcCFBEfxR0m
2s3TVTfjsmt1uXsUAYoqNYctDqXZXUZGdsjnqV98EsSRvqWiInMigjWA7QHbOkuT
c72C4DbZzhaCcO/lVjIr8dYFzx1sLZBMA1bqIU96SLHtHdmB4l54yaomAQPeVADn
a9ba/QCDINjGTLmFUaXfpPPJYk8Wxmqexq2reBz4/EWi6Sqo17RedpqZ79xssSW+
E6jmQpSjxsf/CAiEbJiGW38Y1pCLOtqBrAM5if9afH91ImDd2ZbtTQ0cOhZYPejB
nWujcortOo7EA6YbEFvqNwMdT0d9L3g/AMNw5O1mS6Skb6twyu3FUJgGh7SHP4WD
/BwxIQ5L91SDTY4DQN63Zd5sZTVLTA+cYg+oB6fYEjXwsCI1uR/sny2iFo6coKZ6
JHt4gn6BP600CGPlvaIS8hLNpwucNzdw9wiyNEPnhCMJ3VdlOSbI1/SZF6GLat2f
dQ7AMNFWtprcwR9dRH2fVR3rtpqreNjnamcP/BHrSsUjmqU4uU9Le+995pH5v1bX
iWXzgXwo6cSOi3dotomgsKtQ8t9tZXTMkrXnDH9HefJrOPiJr03a2tgZxosF8j98
vdNWwJFa7YhVCjEkJPWgxWdLrLp1/9INyWRRU5f1fnOKC2U4yjeJlMQOXeN2DdW+
X7NEnJEx2SuPUS14cDyiUoAy7G0AFzVCcVkeLWstpuufdh85rlDLaK66rrFj2NtY
tcOva7m4JWYjrisnWM4IbwENAfNRuJpRzTr5y4rNDRDdw8CEcJh+dWm3hnuTE2t5
vZBusoqlSyS1o4PX6XR7I4flWic6WusLDvw87tKu99vA7UQfSM+QiKbG1z5vpb/2
R5nFMmz1G6kq/ZAdiiftUZogAj7f6EIdHgybTsl71FYIRjP9VOKNkS9hv1hm3viB
8Hj8ng+Z119LpU9SUiC4L+5G6vLSkplJ66hW3AxICrxBDQvQYomnkc4r0D9V25gf
zOJYnraWvNnjgYE6rEdrvZgrgarDR8mkJkk2zNp/VcSZ6np+a+2QWn2DQbfwhioh
3Uy7suTsxTic/22J42IACP0rGf5xXCUA3YzJ7Bq6+fyUeTUKThUYD8Wl2JujMDvF
YjbXbpnNL6Q5KVrrtv+7v8zzHYi3KlkLhwh0UnhRgO7xkN5Pac/lXyM1Qjb5OLI5
0e2zOJCP88d55UjN9C9vjRdcnQF3Fcc4t8tcPZga94pGSqEUIfxFgHHxenOd11yo
R1WboHOTpEnuPRhqY8jaQhAxS9TAKbmOWgsARPcHgSP6bEMPyrMFXuPqEZRKw6w6
M5BS+ObEq89y+TZGBUjr2uGWh/bsqRG75Sf2ccdGRtcrBJioKkx5sP6dDDGW+IOC
bMmpj7oGLD7oCNGend6Xvp4nBp7qabJvxJeh6myXdkG15p5pokL93wmBRILJI9dH
jiidZ5+97uRF8N9QwIM0SUGcrRU4GBwwOb8dZfjeOjYiHE/0V5Krs7PXLCMO+Ihd
BEuXpkVSQ2UahzDA6DHHCb88+V9w3F6ihHRiIuHhds4tAnX+3finw8NxBgBiNQUP
wU7V4yD7ckgJ6rgyukUR9EpQdqDe11UfH+3pE/RdXgvXjiEW5FPOzFM/ONVJmQ8f
zbjtGdqVxOAEtsos+ujIzKokk3HWDlzR1OBujFGcA5Ih3Pp/TTvz/gOJ+nfK+to7
glXJyuKGtY5dOwuWpe7x4/z8ZTRK4losdaCCGryEMEUBaaDm8HVOLppH3HMmzcXN
5017byKLk9XtXCbCyGvltkdg8pAdST4sM9wD4yOntZ9XWc5TJvKh4GeNjqLYFB75
WkOds2owEfIv8YXFz/1HLjqjF/t0HR1YL2AJs4gSrj6Q2ozTMn8otTL5B2M2ijSf
PeqH4GwJYQuU5omGC6sb+ctPdp3acMFNoeqHNa7hxezB7fL4iG9BElWxy/iOziXv
TDOO4U4Ei/jVcYb3ReH9FUViXRgkgk9XeoOw45VP0d2SUKfEzJrWDh83y/Tg31SW
pGYJ7DMigiUH16HBZugR2wMtClCWY3qrfW1+F2hzWxCIzm9FR3ja3QIo+qFulayo
xtMDx7sHIPfSozfyw1TRr7uM9HoNecmuAtmLjJVKIdn00ZJE6Z8M8/82Px+L3lUG
AY2LF3r1QWUhpeL9Fx9szuiDIbZbJFeJ+oIhrGWttTQNWetXl309nqwLY2r1hZMA
0AZRLW2vdcRd69BHNuYUQptUIqyfIo1BA7OJaB2l1nG2aoaavGhS/t1QADEGOC1n
i02P75Gc7Dt/cgMnUSeZELKJPxXHHtKPZNDyR4N3akjq6klH2urYUP5/gECOeaRY
r6L7mF6vba782ZfYQ4oRYcCtdiU0e86V2Bv4TiiLzsBe3M4QQEQaCSZXgzR+dBf/
BUljqvJXCKyVzWFG6W5evtb9x6iaDd0uQUIiBR0nSTvbzQ/Ob1FBnyV4a1m9TzZq
e6/arF/Scpe+1o3rO/u2KvJgcFV1cqihTPTCQr1Vj5yFwQ+NfPrqW7PITsEU3wBr
QkXxNu0JFRXLjRSJoev+HnAWuaN6QANRsb/I889weeOUoUUBxuQZBsd1gQD+/v0T
CMVWQgmLLwQctVfSmm9wUX4V12SDQlfm1IFf/FcSHbRP/dvssuCfZ7mZQMKo+ef3
XwbkdJsLoHIttFld5d4JgRpyEIJw0z7aEL6fCUw00OWfCPGPBKWm5nsSD5+EajQC
2SIlWlUweWciodnYEZvHPT2SEeTcInfSRq29Gn+2JkPJD76sPTLDVTiDJxpLEjxY
2r49Ge17xOr10pYE1u7lnSQxldg30VTUIgN7SiumXGBwDRUm4HAadWcwU2XM0n/n
GTqEaaP2c1h8g7iWjFN6AVAN96fUgTwUk4kn8w7JFYfFS6T29JCpt80lOGdHaQQR
E8eeBFuZHLV0tI5WhpRHI+ChvhR1nx9E2BbP6jKDIOGrHQf1G7XJa3VQNpUUsZHg
H7UIS3XSeC0GudXR+WIEQeZKhQ8SKRZENOlBjEXEYEy7cIyJ5zeDbNNt/3IOrNnR
V0au/HMy0CfWm1pfH4Eh8dNDWpMk4HHvm8/bAuwpk32cIZnroqKIU0/hCXoKpGa/
PRHqvulUDYIUJVv1dfrU4MPcVKdq04FtuVbU+0aFbYvUt1oGq90J12T/6DNcGFL6
I2TXVTI/rTcLJNpNHTINc+B0+8buFhr/DBuw+a/G5R7o8VjwSmlcogwopye6B8zM
UIiidiW605YhlMTJbdX8Ly+vVt38MDJPkdQ91Ot5Bx+clE7TQbWZjXWtGYa6nIAB
olWt/mdIg/VK7FTfnOWLTJUapBAuqTQaq3qq+i/gl3YVgsiJvIdor8elIqP/Nq8o
vO8idRrB5AeRru0pCrqRLWMExYJiV0n1oQ6645fkLinZgiq2T2IgVSw1xtdxgwA0
jTX9WpLRhMnpZmt9O2G4AQkePDz5HGzgiMKrVHwXGwqIffNPKJgV2gPF4t54A/vc
pc7X/Y8OBFOJ5OkPPxVXQX7/QF2jSntHcfs+0EBsYi4UDX//bn+zofahsGgqxYrA
4Md8SkqCjR+Ofun0XHGJAUQGeszL1QV8HDrcA571HcAp5Tw06xJbJ0B5bWzCSVXN
7DXFzCTXmvfMzJZ+C3yiWu653ArLbdl2mnmPWleDeNpPng5AXnoikszFpLX87qCm
TylkzvyoJ5iSwGHNM/nvWEefv9TXwFwB5Tx6PsbRAVN4N3YoyUCkleOeOjVeaJD7
WW8t05UGaRiYp9qzSUM7WhWpWHnk2jieGMmmW3fI48oiPU+au3Hk8x2r0QSz5I1G
htwIuE7f6iNNmwm/2LpYgveOusmWcLefah+SF9B7ui8vGTufe4/wCR/YtYmn02N0
KBGY31OnlmPCtuOWZODvyheNDpKeNIYdcuXkRAmO0WYjMuVz4OsravG3C7E14SgY
FmkclDaLMSlNsBonHrWr5aDgXjDsUYhTGoVViL2FtEpd3O5rGvRc7Rj1M8YfxmYi
9IEW8Y+OQQYfmuTnvr3mA3V4UFOOL9hTYAuHsZO5upbR7D+r7erZ9Ao2cXKm76Zu
MmyGXBRxluNK7+qZyCRt0g5GqoBA5wam5bTK4hT71xvQl1kxjVYREOYo2QdQL+ly
o+BJzjqnrQ/QEJzYKoT81VDFJAZj1SZfQ+YZmC5tmkoSjEx3uSkHHBEmkT2GUsn/
aGu0mHSvLmTgaeyl0iRKg3WxD1wjCkMCDL5pOfCi7JIjKg709DMteq4F0WnRbF5H
USXbBSOVZGT6cIvzalcFjMIpY5SMwzrDLWq7Zj8f12rBw+HNZCviQ5/HpfUUnOi+
XGXHeiXiqcDYS1cd2c+hRnivoV1Rnx3OxWwoaU++2br+65/iQu+Dro1/Cu5+DcQo
/Rp7BI3q0QX7SDISKb1JulfYLGx0B9XyX6oPgX4X7nrCKDBLOPXB38q8vsomDVOD
6CpAsmMmVDusyhaW3rBt7ugu1cq/1P0VOyfvH0INWfp1Ugre+DPTySFnuu3V6J2d
ePCBlI1e0BTw0/vVrVYBpW8xqzrjSu+AD9OUs3i+UWEzz+gowBMnIGqpEOlVpGuv
tHZZNTNPGks8jqbMIJjbFMK605TcptAT8gnn+OqKF/a/4dfmoSh4fwpf1gTjWa2l
cGiKlBBRIJrD2ZfdWkN+9QXz8cgTCcLPSMWQEnfOPNWRtkAuuqvwri1El8DvKW4z
ni/y+GY50bhMXYadIGevIYFnn2m4oAU9/5RljVicHQlUGMFbwwOYHT0HNBuTzeSa
Cyw8yP9G4dw7Jg86WEXBrQfMmzK/Acz9Flz5FavAeUUzEN5H3VPTNg36l2jOGXrf
J0uWXsztyEzQRU0pUcLgh/tYuAE1DZZqCoieAHY0ZKADS6FhEeQzud0wLQ9J4KVa
dZETk/c8Ha399umLOGcFPiU9CxHMmPOJb2KDwxAkFX3T3pout6KFstG7Tr00xOG0
eb+SP+kYLoSOd2T36JgWDPbtpadQlvcmUrvjYs8O/4pJoJBr4C+dwKYpmrTBrqZ+
XuaXUEAPz01W0F7n+zuDCTjpqEchR0KaDUBt3xpSESQmqEK0NQjRmym1Vdi4o2L2
RSe7p961HUW439dapublvDGvAUehDVxUbNCAzPxUprOysQ66UvkSYVgg4YX99evc
H18/YWIAUQnVBg/eIkc5kfJmhvG6NAlh8lNTnF+przifiAdIDiwIaXLL8CTrLTEo
FeetFkRzrvx1z3sh8suZiy49C1q5KgKcLQJHa/yWkH3G9BUjqDj1oxs9JHtOlqSz
LE/iYODh1gVVVffvJ1TO63iDstZTPy+v3CzTqq0Ym36AzbaGHlhBGuUyzu4AmepC
NVjMm52xgCtCKwIaCr3tWGjLmr+70THBovjgUcn3s6FmQBflyYVwPpu4ORGBt1Tr
zU4l0Sk/SnJAqPxGU2vR3v2ymrK8Vi5oJhosvKsQoBnSd/i4U1gB3ONDgKmkveyo
Zn6eJzLqGYvBZ3Yr5ir+x8ARQHk+H+oEfb8/JQvljH6kPpvP9ItSosOqTEL+ed2C
YSIc92lzsZ8/vkzF2ekenri8XE+ixjwOuzgYCM2VbGw2v/3TWyHfQuJ1pUYMtM8/
d8RZRk4j8LTI/GTa7BehP0XlyCI9h6FYflbJDpyAiOEROQnIbD6heL3qTtdwDTMK
wXSzWdaNEsLz0Vk0YJLmRF3cYs34SvdLnIUIUrB+TFCUeadVoUWqwsggBYozR0XH
84pmVGIxFdTIP8szdAEYuq6Dxdio4iJB2cRWXP0+tT529rjqE8ShGP1tgP3qdurY
SIi63/EJYKNcnFHBOI40/Z/IDEbWc+MjC8bqQOQbVbEyoXw0nFs7N8dZtng3tImp
t/qHz4ADr480eOCHL31bnVbUU2tqp9YJYmXfvZyHsiHe0YIhELHW6+Y4yFnUl76W
vlp62UtCpL1sGld1V5FrRZki4sjRUUEFeQGv7FJloi79mzhl4vaDMwEM7W21SwwR
7xwe6weVGp7KHAd+8wBgAidLzEzfjDACKJsTEtGkRYZ9Ln5316lnBbVsyooco5xw
lPanvh6iytR6yDrR+RqCNCtdKgXDyYspQNVjlQv19oDxHKs7jagOFyh0zVWnpVL3
o3BDTSW1rfqC6Wzg0JJg+b3k2/lrQJR5GPw374NU0C5AJy3EUz2N6RpCXIOb1m6m
Xy+DHAQNLGE2sKeCxsrYz4IDP7NCYbVHF8QhjCV2pxbt+Ny3+Ke4FguPOUe4ZaR7
GPylLgR8PHQlxYOR7ohUYqDXmWrgTHDsI/ZEIJpT2H0NQFXINmXgdfkBUnOzc2Yt
0VuShWnj7xhYs1VPCrRY20EwYtHvetwtcqpjgTQl6l1Eg6Ce/YF7rEM0aKdwnURG
Vs2bqgoeNIQE8vSX4jAQfEKwwxo23bb1mtBv4lTrFFyONSXS7onNK50Ggm6yUeTA
7N0DF9/CzivIzSRIB1iQ99dBVmsfR+I/x7Itm1SMPz1pN1cnawk9ZMI3lOBRuVVZ
xDXfj+iydVWkeHu/YudlNh94d8tBahjhO/GqV3rN8AdVL6f8Hz77Nmr9cxF5r3Q8
bdMY6po3m/QeDjA84m2JcGaIV5QVW7Hqd0V4K4QkDmHc2I+HraGKF9NUihz41pLC
GCx9JpdN+ufMJi/T+TuRWxxqLoeUXXdIp7eJ7wP1VW4lib708wmV3xvb31fXykbo
E48tL9JuXvYNE5Wza956bZ9Rp/Ejnauru4YgkLnAwqelIbXoeVdkhGwSlzNxQGxV
Tpf3cvKxDoMvsOa1oYIVySvwiUUWEYSmiilnes3e1n/9DPtCX6UrX0P39BW/41d0
zmoF0+7RnpfDNI2jLt/p3ZuaQfAB1iWeSDv6C4l5Z0K4PkeuZOrFVMi4yLZYGwwp
AZFpGNcrj25CBuPcvCJlkAgGZpgVK5saCJoOuRUT1NMQ4+PRmCQTjTbbkE3eq6pI
vyyPL8FC9Op0c14v1zhMGdrLJ1hdSvqpzH9qAPiwX1zM8vZ/qttc/9ViLfAXPTjB
QG8NvcMltax0dTZ6mlcF7TJyD9S/r/KLUbxwv4/D5D8Yh4WR4Hp+Luj0N7BTGwon
dU5QjZhdoP7STzCSxE7pk9Sx3853SfVLdGwJ3wAxhSjvKIOWcmAV+cUj3eUAv5lz
GEIhpvHchzFMBp/63ysj03OhHy+nJN7Fub6Xbele2fzYuNW6QwMK0TAtUFYLR+6/
UYKAYhZPRfbhYk6SUMsmkycsJmVwhiJgmuhDLHzYgpnyDnVb0lNXjv7PE7djia3J
rTcx8kdAoyORzwXdvRe3VzzWJ6uREoYc1Hth1IV0DgynNZuLhznGQpOG1biaAddV
01SSvO7NSX+rbTRTTMoJEczYIUh5fUuFwvm8zzxGToozBJhWUh2geW2M7yxpVCuy
ZWQfvWiqRJLPBDr++l0BmUBQQofLvTHsmHh8jWaeyoxb+uMgG/sJ/q8FgGR+J8jQ
YhPoTE4wD+ktPDMZxrad1SHC1Ky2EbjsX84qzPR1Ywmq07SxC+CqMRtxFn3I18K/
r8v7RDwZYa4/mH5TLIy6x7tAEi/lBF9Kg9mhSVBGFoQJPnmIKxi72otoGZQAjxqF
XNcdnYRln0oi23hHViyrzaVkEhJbhix53fZLn5Usvu3ePBbfg9ZVssQLqB2mgHGy
FDXFSoKM4zXgWWzfZ5KvLot6dZ2cnD9A6A0+6igaUXLCUU08OMox/MM3bwPFDKND
tY40N3sht9e8CTBXxWbkvm3/T3/4bmd0F7SGNqps/rlPOYPo8+2R0uu2gn3DrclU
l+ilk/wNAfZwPLga5QsTaofp3Za4MI3+H7vOKb982oVSh/UICaPpEiFxQmL9n2u/
wTgUpPKZ/cscz5onGgLnFBV4T2JYJvcxX3S1PePH3C656X0TRuKswAZUIBvL29sY
M8DGmB+ntuk0YbrJP4jDWZqexGCm9nVvvYco9flqbjm+4Q99g/2E9rk+ttBKLSUD
9oW2AhH/JL7gTWnBSFsy6wuGwgG89QuwqRUznI7iWoAv/ucWR5BYqfyFeX54DdbM
9fvjb+3B3xbrs48ITSk9q4DSmZwnx11RMHZfe5rvNBXAd+00RWVkEIDiRnFb7Roo
NKkMHm0cjlPQRmpQqOpkDJrbzVIzD6pRL0Rm/DMKkN+ebG5ZVq8JLlsqc3zxSuaL
+F8BAgzRwYzj39IPqqClykX9avMuPkblW1MmLlILRT4oiXxk7JlI3TEg/B6HOPpV
PVCdpZKl6Hr3Y1I9wi6hiLeRwwIlaSo/cEG83rE4aTAAxCWoOgn2DTq+OyDNggVA
ahM+ZlIDxAEX/eNXF27OeMEKI5uluA12dO2z5K9H4NUN9QJzipoA2Y+CaHLmEREA
KtvY1s3ldhDf3IvrNXx67CFkWz66kdRqihzy1sW9kSSmCA+WwkhCdPe19erz9j2x
YwyuNh2OCn041DdNhFM4erlkGn0XX6jKfHTio+QtEBQ8BiEUikk8U7rRAk8h1DKk
r6A7EaeO1XA9+s0JoxTOp4mLGKEyF6E1Ql8+OTHH5HQGS8iG/1Xy2AsiwGwwRWnJ
m8aBebQoYYl2cQa0nk0fKVInBciHOOIpoqSny6C9v/WUijzzAEdV5iQsNa5rgMik
DuP4K9S4xjcjmuUzoW2wEzbeX/t6p7EkkueFq2g4iq6wJqg4UOG25PLtsaoGWcNI
Eiw7aWJy5jUfNjq0L+wKjnUOpKlCBtTwhcXRgjoi38ZFFuQSGRFvQtoXYhO0+gce
fzYKyRUCgsEI7d6L/ZJrqGfNxy2mnnJS8LxLtpaN1VRt3Xjb6STSV9Yd2pvwsjl4
r07PNWHtOxt3d8OYR2tWLxuZZcI0xjXrbuGMgQ+EKJqW4oCaonNeR8DhUdutODCF
5VFzPbLq0wulUbywWDYhjO74CwTJ+vCzuGT/Rj3teOcANzPYQ7wIlhifEC4iTOKP
UYB6uCEZKpXDI0JbAcpDvpAVBCPBJepMah+XU7urqMfuhfxM5zWZZ+qoOWU7EYI3
Zfa4crzD9gVOlNnK2nM1jSovp1OczT8YY8nTmtxBqkKzuhkDWWw3tl1HMRl0Zf9V
IeEIgAIbHX9qoQjQW3avQcrCeUsujXjZMEnyF31JyR2KNiRXh+ARu1aphoTiD8pL
MfeP3C2AEUzHkYJPFW9SQmF8qQO7YE9PBowBdCu9kb4AmHAQEWytuj0kCh5tPzsU
nEihOGu87qpdycfuzEy60OYwbj/W+Nd/hJnibWpvyk0V8qdYtSNcSZ+GnePudv7k
ecfUkJtutKymlC1DTlJyABROk6Tc3W4BF9Bbq/bVVZxkPxwZCeznnwy/cLLacbdu
QYxZwHYnFphse36xFvWYF2zQ+IB6K64HbdMGFTWUKAZ8uwEQYzQalYPG/wxLBdPk
bxL8hDoLiirZklm5/9bRXVmy9qTeMuwPgP1GcuKlKerZgAfDUd7wtDJ19GqexDYR
w8AVWV0quWQpZJPbp47YRtqhA3v81r5VzIIUqi5QTwqLz90SP+YA2nUpd0Ais2FA
tU0h2rq4FsvjpTOoPfTK+oY5mnPaDn/gH26jBkqYJ8HR30i7dyvPClZVzjwXyryy
xLR7O2mqyXDRMsH6TLD7X2RLxKdSlH5+Rbfojx3XDH5kuF2gcHBrbnSsuj7up/eK
LeUCbq8h39dCj3BjZSkX1GVldypATPRQvrOyK1Gl3muBITOUK00CTDeojRZcXMMp
/hpKuGWeb7h4+EdcWx102yc1xEb0wJj2fwjB4L2g5yghAPZz9T/mpeISEvGFCz+u
QNSPM2vPqqQtsyK5eCwCLegDd91WTOGG0RPLfFWOHtJQ67xWpmV5hHgVOlRN8lnF
fjfQ0dNKEuN1gHMpnnIMm0N6V/h0vVCfXqXQ+Dk8aFflk/XYalbE42jEOJP2VEt3
bNK7K46A657ftu/hHT0rgWgTB9bRQIhEdIctl+UtyJ9cNb7VE4fq/fLmEht5s1Vz
+8kOkdThC9+0Bs7dCso61siIBygteRgSCxZQgVIRuXZQ2UnPrVRO6XjWFSggfx13
NaX5zij5Wd6Uh58sNT+7+1+sWESmVzEZ1vvCjARvv1QJ74w+s3ruqViZWJ1ScCIW
kPBq+JZxpy1sYlXOVuuvK82QWXIFKArsP8f0ggyPOMA91H0qZoQalBNrRi90PCej
uw9D9ZmhUmtYMJSOT+3wwmfoP6wRWD/xdeMa0d7YHuQL6H/w1aVEsvH6FpEoAi/G
ycurdVin0TlSGSd+Q5ao57ttG+0rEQ0FIPkhLGgrcqn5s7MCeg0hOfXUBBvBlvh2
Z+sexCvOZyVOHk40b/YnN4IHj3jV3pU7n06YfJv3M2tpsAiZMIdKGvkSP/IHE+LI
lt3UvKX2Le0oSY4q3c3aEQ28t8LAtiuS/kd3VjblcVWvStTFJ+riUR3R2MNDiP4h
zvhal8lcB3ySjfLsheARyqUEySn7i4mDdxMzvUYv7QGTngTsZ4wVF+WEf+U5Z6wS
VyQzHq6jxsloadIARGTT/tlnbWbcY6BP+7fwRkeuAs5/psVztrnl5s5ZS5atU0l3
S77nuSMPpBkXkeWwkBPEBuTVuuK4Db8JbBgA3jW7Qw+JDKQU3cXcbr4NFK0VOs67
NQDDY0AeRc8WVNqT8izBHcIud/TWZLztOmPPwmUhCxY54HAVzl6yU8RUdkaXqKF1
yWmxtwyO1HSPG2yyg4xUMfXbrnb0oNMspkK92adAi39cVMNHIGY87S4E48VyK85f
UQvYJNcDaRvRqP6hQWQaItjemMz+RZ3M9OMysF5KE1b7bQbM5kWt/pEb/J3TZH//
JQClbGtcziT7N0VoqcjF1fBxi00+e9ZSZ7KiG6gFi1JlnqVt4PS6ejIappb2dYnO
rX/iiRY84vRYdnzHCE964SqwyTsPnzww0+hJeTxiiNQb6+RFCcEo3K28P9UK0WC/
wu63dtoB2Ct+X12vgHs2I+U2elUaf3TfQEbUuSIraxZw3nG3KIYFTf/9wtp7WBL6
vKTmjFkATeo8MMWp8Ok8IpPwujBAZMeQzFQfYezJ8pWw3nP4Rq7xARanfqoO6nbB
cvsdjjGqtmRlLJ/cAo5rKUFdQJxRg3vtYt6jhJz/AVSL5KZUQLIA6Sbq54+LFwqW
tUody2WTr5k4CISjHN1H9UfWXAVCh1VouRejlSW9MK4TWkOScjZzsfzmlAmX/nc2
8yRvP08p4gorKip9scHIYwKHxNzGN4q1p/zeocy8mlqi44JbqCvt7zi1sGRNJ/+3
6EgYedEUJY7+web0BiJ0P2bilVixpMYFh6ZzrDVHrJHBL3F6zMHINharqCODt5T7
+GFd1g9p+1eixajUDvlqHHfVJtq+IDSnvazavzmFPJQB5tQcqaoJVvh2uNoPlVb7
FIlMYiVW4+CU2MX8c6qE+IqbSvvxzAKJLe3wrAO6u8rW8lVZcJP3soHHhCwW8Z6Q
zKNk7oaffix+dXOBmnhuWgV3pdPf3pMYPfiKwZC8Xj5JsOWA16qPumuokwOQaoLY
iNPxU6QZ5K8MbgS1w40YDvRvlyJHyvsQfVr9oF4bEsodXIVLTKMSRduNvEwC1Mjo
eNWpXUqrs2p3NVpx4pqjOlL1Sk9uuOHAj4hK3S3+HSg6tksb284P8PcHWsITGOhp
uSKL7xmBU6P4bP6QFRSmGJONBY7C/K6o5+Hdntdszzz6LrDvMWE9mMIxYydkw+Sq
jD78TUQ+xemdmpKefwPrd9fnG+m21aIRif9lBut4r+6gSIYr4i47/u033Z+NVmkf
zKaDhQbmejuHk1Z23C08D8rYHw8+4sVqGWGnhwRY1fn1tPJ3XmAEOPf2dQiLBePd
SfTw8cHXEn8LI+bTcCwT8lG/RgVOyAUt5xs1K5rYad18WMJRlW0fp1bMlsw+ZeQ2
ATgj4eIJP2D4LzHU8M//1z3/xw7ZJdhgW7X1pXuN1Os04zqUtTABIV72VkShwZM5
EUa9CZKLktK8QMZfZHlNCBj7V8Um9mY7HxnaGkzJJaPZitlVNAHHLiyzmNhubPc3
YPteqtR7a8Jmx76A8i2crWxWWjWWcsS1rZeJh96Fdmq9vwQspPV8B3S++7drQ/mV
AGaVcaaXVGOCB2O8ije9qyQnMA34/uDY7jM7yr3lfOpL9Waqp0zHo39hJpYz7JUD
WB5RfpRYvFDga2WPO1UAFeh7PMUuNgOiz5uluH3mZBMi5bnJXua5WurVMJ9dUJow
6Lk6Yhw+GqEmJ00Yq4wcYPii/VxfLhA3pohVWKk0XFJGfs7dy1KZ5bJeUY3dr94L
EfPfKz6fiZq8aKxdgE3Hs1sYuDdXFtjmaZly4W6IqTA+r2OoqkLt/bjb/EnWVT6S
f09KyL183aoeUevZgGYALTYr4hfSeOP6wObqoDtdGNXmXQAcIL0VAUAtBsARNy7C
kaN2PLZdLYM0FIp732ExhLA4yzg3xSx/eDTbLr45fHca+kcszAcxGuCyFQ20za2E
TzHN4B++tmiRSqn1VnNl6QpPhpgp4CrIzdvvJtVCjAaVmYEcwY/ElzE9BkDpAEe3
S/1crBAYe6sVMiAohuk2Quloc8Pm8qeWwhfIakS0Litz4LoGSeOwVdtvhJTaR5iT
PsxMsToDvdaUPIGS+1M7iO26w00Ad9udgS5n69k22x/aEwNlcbc9+u7s1H+l/nsb
1heAmmJngy8YWfjtCjdTzT/qf8huS+R62DtEghue8OOg+8IlrcfmipXnk75dxzwv
GvSiht75VmXfn7YkJvyRUiMzZdymozBCVd3lLl8N2vlmqsp3tfGvvlbXIC5xYfyA
VRgyamiql5Tj1f3YkZ6XFIjOD+dtz5V6jF54SbSBGs+PL0Nb/Jbi/DoWfRykNKm9
J6oq70dT/UaCN2Plt8scVbu/c0eXe07x4Y2hkStTP5Ntgn/kFQfSNs3T2YF7F6sS
F4sDVI9vl2yvtdzpADTIQa3HAuqhbbuxzHEUEXhJ/OOKd5xqViM/9BRQLtW2MQoV
GJt30XmFnlRNNfwA1xxT3geVCwFhxdrBC4eQ9pFyRRvYCX4ycGjQfFjRTCUxwtAa
OuLtfGqZoY/WUA4IQU2p44qi4qqkZhQjpzfhboHkjb2rbrkmAJuoUWG0A8VowiXk
ovYSmQfqgzxMu1T5uvu/k0h0OBqspw8aMntsytFay4+r51e1dFhKbAs0imVFmvZS
HFVf+0R+6AILSBdRejBTMVUy4MBuAwcqcmyWiHiaQ/UPHZUv1x7nt6bxHi4kuj6/
utR0x9rUIl7SKFlOHxPIeq/tDJDRVw51Ht+5hcW0kHTndYItce5DvzMC1EVgPhFy
sc7tsc0fTGDW6TpCRpLl9XHUA2PCuY3rDJ6UIEljed2/HHfnfcIn4QvwZq8FS9qe
uYYgIaY7a3GFlsa0rWjlBStui2Ly1zuNxkTcL5CzfeABotKKSUOwB9xq7MKKCZuz
zQRhYzip5QpABhzBUjZR6KLN4BLET4L2b0mMsdds8CQrNYc37oj3Eli7ofmRDxsE
mE+AuUHyhFCWUsGrDaHM4k++VgC0LxIzrj0FCcDWKNVZ2PX7r+PmDt9SGWRdIRmR
qCpM0oflVSCJWdCY16C9mp8N4+lxLpV/MWM8z9M9fHqiv2lvyxFtqpQrhT5Tn6EL
nEV+rLcKk8SQNFvtJ4x2Nc/hSmcCbfmc0GUmsq4MGgsTbKpC60q0KCYphdUEDGWS
lE5yZschsRhBJJ6U18jgEiL3f7caogf6pF1lOQtHsd7E5oA7YThVKw7W8Atw5jOJ
FvSnyTyvVZ/4GUwfLjg/yzX0r8ftxluJFjiME50fhEPZx4/17B9kbwE+LK/3Vw9z
YVwY/hNAAyeQRoj7U04hhGu8dLKxY52fO6ZsvgHL0mSDmFteBH09OgacLpHICqH+
ONovmgZxzXcyJnHnQyGrXxX/Oon1G7pf5OE1AHHRkVotG0BN48L9UearfwlwUhJ0
XtshW0senXwwvnLUthzsFWTIRWbP+qbR+9dfytiVQeksHQTJC4ZRY0x0xMxqWaUY
sqfKok61DxuUw/MW4iyfI68JardTJ90dWf9Crdnm6gzBJcydBJYldeIqIbHSRfX+
QLuvuVFgY98FmBFX+UVgB2vvBVlDPvDkA0Vx7Shx4C7/ghHG+lQCYHoSGteoW9KD
A+By84Yc9lbzjXBPOxhvREFzftaj4ZCuw0EM458C6WrIh2QwM1DtoezaG1vxvzZQ
8F60fH/ffhOO1YoBSCd+ue/N42xJtY5Xth/TxWNp/kalx+KG+WYxuby+fr5klE1K
j1o04WrJSYS0qjpjXmf/7l5BdgKVMZNnpa1/5VAZrZEYXejEMrp6jB0I+T7xSmsL
rDfkKGsneS9ahMQzR4OZ+06XMLKPdb52934IiyzfJetOEUF1nE760pAK0Mm3jBi+
sL7XA9TNufA9WTGCp96l3I/+5VEECc1g/csaz9RXSoTdFUIWOld9DuhLiKW+JP7Z
EA04WyQ+EajyUqPx4rvLJ7bbqhgA5nBX4srnTyn2vqXj2E3R2CaRPnu4URY4NuDx
aU/WTXPddkf7H3c1IfzULx02XdtETVIpmka+f80q0zMwk6FXBeV67D3UYGwJdsP/
04jonC66nVBTAlHDzNqCSkKf5TVz6rlANNF2s9PdXDluvMxrmFAE3AGtLPKthoaC
OdPimbElE1zjfNej7Y2XeoWt7SSXANYzNIkc9ZoUe68Z6GOdsSa39hL+Z63rT6TO
OcV/IhJSsHqhvp/OlZ0oSrXlEYaIrwrLvt4gpLUx/YeYxPQJTo+G2KYMA7Vg2WBp
7ANkyK6sHziY5GHUOeKQwMLpziXF6d6NK4dwpTbv9yk7iWL0gO8Cl3FF4KUVIH/H
ajZXg4JAMU7YvhHsywu5h1xDgOu9kzmQy1hjHkdpxtQK6zncuaB23t3iqbmlW0hY
CWow5eeOs6He6t8H8tkZlpkgVNAvcC7uN5T10lm+SRzxDYbAqXTc9LjzGMO0j1l0
FuTkCtXFPq9ewYtJofA1GLgdJt1QkTjjxvmz3IXCxbYEaA1GxDkmAJa6oJjjeBdm
ibbJW9ediKyfj2JccfF+pzfRLHt1T63e0/1KudtsZftTayvCXtrQI5DlQKU6tWBu
gY8l62Q0B9Tcav+KbMUfcwHV7ZaKwbj0qxQUKcwNP/bDiACff5MAcXMNI87cX4FF
pqS9jOedRI358VDCkTfzGqtxCH3UFc6elP1gHu+NnW2RNmBdC4AmZyTbZ/BVaCnE
CVv2BovjZJNSIx0iy61H3UdwrLhXSZbt2DrD5Q7vV1wkXY5t9cJ5P3/lw1VErdd8
8Rt+kHxom1sXVmSvEZNjRXi0m3+spVIH1axzWiMBGyEqvGzCFLpAOSdBC7QeY4bW
sQ+nCsuZ3iTeyp8GZPADdw6GklOAhmx6UTdLdhB5FDnCMO0u49SenlMN7owzgZbV
tzAA4LDPz2jJf6z8BHCgP4UOCfMu4j64X+A2fGiIv0Zt1J29yoZ8xAIJEUEu1KNe
LYISK+naUNDSANE00HaFQ/Haxa1+/5ABybMLaxWaU0RxRIoRCVLfgkmqz8G3I5e+
z6B3QJR8m8VjRLX9XrLE3RfeqRkoWRiJiiRaER9tEKoPXKqMyQkSebeXDxB0HYcd
hDqMTJmZyx6yHvv/1AH52gOLVPCkB4V+8um2PGPQX7anDDZzTkf8JrIZ6rLgvhcW
GtNnvdo48vM6RKOuBvwNnu+eYQRhXD+qJKu3SBL/t4hhu9SfoTJpODTGge3cVa4r
sJ2WyucVbhY/tqFOGYGA89vlMkU8j2JgR9pzq2RbWAuZ9eu1X2ciHoj5YI51ha18
zG/NkQNPJeKM1HQUpX5p6ctIRbWDCsPL4aI9VNcbkxsj1et9Qe8ZCVm/As9chGA9
WT4ApM6DPCKvOOQBbzIuD44Dv25nqSZ9cHOcD9KFR52va+fcWSZ06lObY2bQm1qF
Zu6O06bre0pWmtVL22y4afJ9SEF9r7/UUqtm4pvu8jfUqclE5vfLBj6oKN9pmUIe
nr+8CjCyfXgosMpgCJi86hpIwKD/dS7mj+lVVMeDwV3exwGgvsZ0V+cGdjxVuwN9
LZRLjtXio1qS4/LjbF+kXUNbJ9Q2dJy1QLvVrHSRJSjx+ZEZCMlBrK3tjYAxH2/9
TNBSca3w2YwS5+SHkJMAHhg9TOyyMk04V67twA/FpbLcckhWjkWVEOVrxx04ILbW
011rVWTsEFEtI6IkvXZ7E/sDB9tmlW+6HzvFIHkh/ePrRPng7ySnOZ4DMvjqkjok
TaTyiICNbcatOZA9O8MMXhbaABz0T1oo0a6K5o1Qq/m4w95QdI2eKRH+jFNSliNm
K4ZqdLhNu9PjwMcbN67r1wreonKb7rlPQaHRK1RNLkw3R5niLxYf+zpiXeoDgdhr
SuiQHhr/PVnZcyn6Eat/oOEB1RzxtLV5xMoKrQdZ8ODHWh/JqQvI+mpeRIvauAPD
9NJGn2TELtVzIxKUoO8SfPjuBV/SIFDl48yEh5DnEoPb/TxpT7I98BejEJMjCeNN
AdKJEt9aAGkzAiC3TystOauYUjgH7g49ccslzz7lQjMoZl8LveEoaq653zY2GLu2
ehtNRFEhteJqe7gxf2j93jxKGRPRx4mPCprcIbRL3ESUhtyrXwfleLHUmUcad1e1
a2VWiHwL+w5hgaohX4dFVMO8Q/h4BSvsrHR5cLqHgy2jiEtQeVtEgqp5FIYQZYo6
JlgXof2o342JyPKNuM0b97p+/P378KHEjXEBXGIid1YLXMeiu7sKPiCImmBQen3j
NNvlbnCXSKJuLUr7jdbvuCqWwRtB6SPg9gaj8IOkCwmvrKJdueXwgxzFi6B5g0ku
3TUQVZsPL0LPbNeOLp6wSRbfZpHhHCmSkDukds570bn6mQgGkP+Hlsn++6uTLvDD
UCMBbCauvLcZ6x1jngJQJfIxXqrHIYhOg3zvQNZx4zU3ga1AV6tipGNct8EI4frr
lgQA4MH2cFMDkBhJHgi8EhKX4O2ukLriQvZZLGmRJAvX+Btz5dcI8XaKyVFlzyWs
BxRftR+dzEwUX1zsn94D55sY1xuNWAjhR57n/I1UK9+YvfYxQXLHjM6bEoHDDN/M
E00Ka97rj9Dw2VqUjfmD9JlVut3LiV+UQY1Vy8vrk53p2tedZa0CsI9/CXXOQ6Co
ehvURoW1uLfveE0wKCvKTpYkcINI0cHyxJhKgx3+sGT1nAb72F8LneJ6mPjPaINu
e2eh3Wt4ZhspeEYwdToUWz7CdFYLe1nFnzHY5LO0/meu/44ZYEmzvCPK6//63TXC
GHiyIi1lPlJ7PvADCF7HtSen6esDLeusuG+eQkA+BAwpJ8fZ+BQ6mpyhY88kb+aS
NbjuC3kEXw4WICxFEl88+47OCWawDo4r/xC5pNr7r0C/NPqRWPDzb0AEqt2qhaFY
S1BvK0+7aavqgYfKxpno00jaT6gfyF5t6xSQIatt06SSpE742MAAv9FBzWct730Q
KWBKwgT3OSTBevjcTt7W6axBXhalxJyziDZ5n7JtnrAlStTFMlISZJuZ1JodejOs
fCl2xMzxCFXjDSygLC/a1p5dV6vBwUtdk5ztcbBrECPpBYv3PX0J9fQjHs+hOWlR
7OCJh+xMOhekFvNrPyuI0c7aebViJer6eljLmmer2uewf5I5qSRBWmKqfMTVu6EB
L1zECPgwXhJfBzIjJCE+SCRaTLUG77rTeFG4j/cLeXndCMseb/uzUDLNP6kXlNuG
0zuuBZdZ5201obWI3iyILJdVlNKkCFg8XOooQbTWKud6EmOfOqsar7oV1emuOVlM
mClbDNzYWe3TMa9hCUutGtGzZ5xMe26mv7wDxeJ4Odw/mJrkKKFwUAm+hRw/PGBR
CbdarFA5DjTS/uWbGUbPQrOlnkvzZPwyChj3WRJH0033Us27dsY/n4U9s6MHPYQo
mIZkTykZzYJXNZtYycybOL5VSQzPavPa3vzsL8633Mjt1ymmE4HsfFvgiQyMBKRX
GgBq9Yt1Ia0P9CzP7053VFl30yqtHKCXotFgR4Z49foW7JzDHtXDEHKWT7elIEyO
DHffdlIIi9oUF2XaXj2nPkYIOj+JXIj+ix0n3w3SN9Dp3mVaVstOvcGkC7Pay7nZ
kPNBCCeEbXtg3eVF98tZ5/xSDHHAZfd5PmUz7JSxRdMIbHU5MGrEnDhkEG5xJyvx
6g/YqXh7ZamYinThBQwQXVAunANcZlWXgsc3OU920LBF9SISCRuNqwq03eT1LLe9
3yU38uLW4DCnrf55DspUux0Zgcp7aslqYqc/DHIDaIna6WzFtQRyO2qJlPXpAFEu
a41mpSq1OuS0SfP8vB+h/l7TiwDmoTbbZ5pHd5dOPNMoilFgXiL806lPYCg0u9Xh
qxmhR4I1Xde686aDQdbYwpBUYUBPyIBbuUeSWKDeOjOcM8b0l3O7frQ0/thn7rj5
YpaOINjjXSjABuNsrExyHq3spDf6eYvgtU3a2LFhG728lOMrcQtDq9rwlDQ1r4qd
EbnLXIgzmVm5S9T2EDBpzhQpGLw1a6cQXpCY1/uZV7H0670PNrEFin5ER+MLjZNj
fWPQS0+12krAyY//xWKcnJjFBsjjwunjmuR91YgCgELbLWs/QIjcjJutHX18TLAN
BTwy5xySrFN+yZxw4nhXygn37eCYv3Hb0AHJ6Rx/xMCcDQbyrbubNCUYtaWaKjot
TiD4APcQQB4TtTy4SvXt8kJhj9KAlesCGplE0YtoAWla9mjcTztGtevWYV+gqpj0
Rwuy+7o9q6WXF/c6kLpAbL0KAe7IVdNwZDO/ziCl2KtUgxGk+2iz7lZuttlDDNOo
KluKTCWtEW2jrk4lXhWk9piu3UHlrABsQd+qvVKUpELDfJIePWtrS3PN1C3RLmXR
vpJQLRaOGf8zIJLb7crcRw/aD9ykJr23BuCPtmAfRShKw+Ywh7hNb44YnszzEPQq
90zE2l998w09cbJVJtLxUoCbYU98KqNi7GlscKP8k2c7f5RST6/edcYhAiIk1Z1Q
ufoy02oF9I1siQCG/LRDORfzxsV2kon+U9uuby3Y3dP3USE1EHtGS5pirk5K6bih
rlfCYPy0xNyudNpp89CjDOQW6ffBxWT+bEiGakPMvbb+81wD7sGYnqo72lMXW2Sd
C9zKkV/g72Y4R+DuXy2EbCSIWVQSNAOsGDRCrXF+qys/iT6aue2HeNpmC0oU4C0X
YUQN8LHzxkh8h9MKD1b/a3v0G8upM1RXbw88yU7bLApxoT93IaK99viJiyrPThTr
Z+0FMw8xoROHF5t6IPjTMdBXVfZs+egU9jOwd3LVlJ79z71MUjeBMopdhJQ7GSNc
o7zYZkalWYJg9JiXnOT6ZyZoYfiKL9Sk/XxXIElN0gVfooVcKAV0rWWbCHy0oVqb
7Fvj05OxJu13V0O77pF8UNDvLvqGFQkRvIA6IAHFqQYxrBWErDSsS9UyTmRyn1Q1
RR3wA9X3k28pHfgL9m2kSYISBp1lcTEHuNJUWmKO5h1Zi5DKXvp8H48PHH0OX5u0
qWHO2M+/sKVyt1JEam55Le6d9nkNRWBAfQ34gZhDm4LjEvns4ilmFuBFDwM59/z5
mQ+7QeTepWjz2IjieSPRLw+n3W9IOILwY9gtTBbN+DKLGQsKsmaNA85mvlVmVbri
7wMdgR78rlGEc/L7WFcnA4vryza9J+eflcI7m8/7dljOwhx0mRiiGI3u83lgJqiG
MUYU+vh1m3cb91mmc+GwmDTQOK2l2PibgUgEn/A9o/nadW/KtbZFvTE63g+MxBbd
W28QAm4fqt+XbcA7/uq2LWsrFLD5f/TCDSvH3NYIacYhiQM63MLPMNIfOM+E/wbj
rg7qZRYamfyKPm859DIIGjectfGJzpvWABXkAsfKbtkIaocGPh1jv/cRjtCuo8Yz
Ky+hbFZ714/eTgsaDBEkKAZdWD7sfHJ5/WAQmnsXmrhZbZwe+SjtixyWkHMIK8Fv
/L5QY3DuFH5L2T1IZj0uyhLbIjfOoCnGkHR/vne00HyE/X90YnmsevbBb+ltVAFZ
88Ln8F6iL2Dakqk4a8mb9qOcHfgXwU1mAbidPx3wqh0J9G7R3mqitZGPJd33h8R8
VudbRLBCq1c2FFew2dF+F247SHdu6d+Dgin4UflpCnGXFSSyP2G+qoNHd8wIsDq9
QhIkFzdCbNGX00Cw/GbrMsAV6h/wM4CI4daj+bYQhzV+fo6inmUUHivAHAhubk8q
ZUhArnIHMqu9X6DExHEmv9W/PVQF2mORrmnur8bm8Ryx0wUFpVhQmS78K0VTqH5P
bj+GYY5VCl4CKgB6fNeiCDvzV0kQiEzEcap7DWv2G65pxATAz7sSVfWEMWZzCYgs
7S9gpYf+0pITEUrQA4BO7Xzkp6OJCjjsaEJz9wUF7IF1xzZoi1sNowEsX5GwmfEO
ZCWV2KdVq9Mu7ql+xzCRj5Y6m9yQfP0oszmdzvRNVcrL20Sp+MUuMQ95E1NnCffZ
pXdRb5K0afrZAFsRAsBlGxdvb6oW3+Tj7//x9pdABccJGWx6Kj2cLgaUVaS8dd9Y
RuRqeCdURTyoT5nEGmh02z0jkxKtusAIKNNY+fUBQCkBNawMH6QFlK3OYA14qu+8
p4YUKHUjLdZQ3A6WomCacKlnlSe/vEaG2i3pNrufUHUJd6nyAsGwjjH1Q+0/GrkQ
LMCPZdXFXNFqTbxuT2PH6kD29+2AXSEPTG09BRvfB1cLGFzXKwGVfiPXmQeDmUWL
G5+g7vuGfxqqdH22Ij5kZbyfkDAaxyneUyr1oHJKAkGLIjH2TokqtQFN7qIGU6Hr
oJEna6xh229SoRCei9qGu4NAwg1khWI8VnECgnrwrhjr49hJa4VjC5G97msYQpGH
ZGNfGyEp781SvdmjauD19Fx6LXDTErbBcrnvx77NzLuTjJpEx+CaWNgQbv3tFaso
HO5oYUFJaUSDxGFZ6dxklGWvlqDoKPk/Co4bzcEFVy8BrwZ2SqhqzCRj+lV1yhOC
f82IQoO7wi9fIXY97bqy5Sn7szPiDENRjxBZpfhWxB0kZ25PQz4w7hdGhGW9v2fl
aID856sMcGBepuMyh8ZjDBTIkzM5EVMOXd+2NJyMevhAH3JRXcVQ48q2xTSTJ8HU
38UIIlHCeYe/BOQ2NYL9SVSLfLDe4OgLrFAwW+cLQT5XXaew5Z0QLMuvrn/WDmAU
NrWP412VLndZJonFPL2Y35+iN8OG9+bxxID1cBwcBDjR189yIt/uNkMbyTwQNs3m
HPME93Q3V5gb0I1DzUlj1z1elLdcoF6J5EP7SEtG5yh9FKRlYshipssTUFLsjmU6
Fq6iNIMm9we2RChmt7QqQ6n+8jECF3KMrUxSvpJvuRgjr1zlzNQhx2eWXKdzZWnx
Z4KUfN6Y4CBFDA0nXLbaSc8m1q668ahm9tYFItKvheqDcEvkO3OX/5Vii+UB1wCl
oz1PZvPngRKYHPAYdfMoHl7lUBe9koSL6nL/giklQ2hF4AdtH1mkDz4YYE6tLXwz
JHQo47ybVzlMnVD47kcq55mybY6L8oxcNJF/prZXkpIJFH4QeYhh01RE5Eriq9Sj
ensr7ll9Fb9vC9V0G1xxk3+W/U9lb6OfnAnwZjGwu2wLuNPBvwHRqjNhX9NJrAjt
kFRk6znQD/kA6mLekuRSHjDGE+7m7otIJ+H3vaWQykm6a6MdU0r4FFZQdUZKBv9l
P84gZ1dklbTn8Z7yxoXtMo8g4bogYt1PWJZnBr2N/EsOKq8eIL+J/l27UeME3Nu4
5huVf3Yo/0i8OfEnU4FXOkN0KFM2vW8tUSRkACixIPghF2nCVHG+BUQS3a6JLioA
0ID4W1iKEI3nBh7WWkEgGmX5cMgD7+BBlaAKCR3frDOnU6tAKbzL9A9nOItcLQ8H
/QOuXU7Ksmm98p1TuiCAmmZQvNcd0HBOhfr3+U/h9YWJ1YbwzD6j3u0WIAG3DvK7
NcOwwocYSUm4v6a128jduNv8zRUddRCnTEIFP6J3ItniOdKq1V/Ux3ZzzcLmAlM5
MDNBct7dGm4FJhsP+7sbK5t4rjy0PAhd1EA7qX7EEF3IDD/DXSy2fjA6/LZZ+kcJ
uOjJLr876f7O5+fKFttnRJ1AoCI2ssvJlz/Osi9bCngDFoOGzpzCU+Sfhv6q57On
1hSX7MWnIyaMOnNkv591EtUlgY0i87gQS2coT4DetJoPzDBiLdBCSSE4e+ioIHqI
dbEjGsd4X1rRgxd7ygmb735W4NvuEDKhGNBbaP4CVu6oqqtt/DIJDuWMmVw3up2+
CPHE+51iEZ5a+l2HZ4aybY9kH2E3jmjnD6oATSjtGegaKsSfUGaFBGhbVBkvl1mY
uoTy10xeDZL5//P/lgHLoRiOUpCWUAxrcfoFAKwUxWqAnRnkGePlOs9nX5pTAQIy
++j4/hihsy5Yskk5ZDynbY7Gi5peqWhbnx3B4s0Zo7yYLH+bvHi2X4M3ydAEPupd
SgsQuVcTCmdBTnGV33X255g6vNabVFgNvEln/aUp43djhf8i0nVHFtcYYD+2hOxl
v4Kp2OrfwzNqEp3htQzGSI8v7S9u+lxW+OsojQ24Pv4Wqu4+m24igtqOweHUGh9h
HP7w2oiw8PzNrn4cUQOhKAFSw7bzwoZIrXb6PAtJ1w/LR4as148VxLASsnayqL4S
QJ3f+056Kk8ozfDas/xnjfpZXTPe/QEolpeXIdoGZMDPKdX5qPjwx/c/SRX93aBL
O+iZLI7GM/gs789Wb/S2fa6bQq1W8IwYjHx0j+5jFiaRSbJT+DSJgt+jpsWxXmV9
v0hDOpYoZwIOAYxrL5JN0/+B5UwJZQ5huhMX3rOUU1voO/giWlOhP0Eb/9LOhUs6
523KvrML86xoPL5L8Lh/nn8iK+uJYHi+/QRT+NP9unoKUfzYq2WrmFuMQC2cPzC1
YZcKKQ4G9f/5vxWlLd+MGNPnjRbahKDsr7ZjG2nHZioqplOfZBbAjL7t5xNgfczg
SPZFBTTDi23TpZHLtlwLjwygGENGJdS+CAWvCRpvXVT8q1sB3syva9gnHwc+xYQU
wKF7s4uWyZY5X2Xm2oHyLIPvHyB+/ECAixsrWOwXlQ1IreMuiPPU+gA71D78pAc3
5lcmEJ9L5U4kXpI/jzWKRsk54GoWtA+CaD2nRC8eKPUiqqLH3aNcJCJ2XF1Bxa9p
cpzcTlwCi7KCOuuhF9pzcd5xFFIVtJy3FBMKwqR9kkq6YENnvRXK45r+Lp2bdpzw
O9UJLP2A4vMBMj/BY6SANgRQHc8tdvxrqpILLHu1utRF6rVxoyIYTNWYxyUitZ/q
PZIZRhQGpYN9rvKIX+7OQ+ccCMp2qyw7U5CaTfxzQQn4K4UbRgaOXLypUxJ/UO71
/ug3bakZQKzBPEAae9h5iElb7fP8bSyxUiB0AgrCsWtzShWabHk8hY0LTRSAVOHx
lNgFm6uJH5V3awsUF3A+AunG4l/goCo1A+LrBdAeoc7k3I69iPFnAd32HVlkBqPa
/+FaLgvirSudRrTpymN9ZyQUMxoz0hGHgwTjTKrOe6onHgt7TTIEF0gRKoc33574
+ehVduToiyMQtwpetbhaIQyQ70MZYH687RH2psR2jQNRXseg6yJng29oDNs9e8Od
i2jaS+qZSVXOFAZ1GZDSvqtSL23lTVBgwlsRpKpdam0YzCBuzJsBD7FQVfPWfyxx
M3rPUTpfOioh4b8BkiTLk9LP8qhAK0ZjcwS7JZQOqyKluBFKUu3oR1T2vjf5loBf
f3owYWAuOQKc99uDJPyalnbJ+1UvSRPch74uw42YxEmCcm1hDhxcu3dHAnlP3HJw
hsnAN6edqEGoQ2GwgV8bu26N7fLC7j1roD37//1/hq5B7M6ZSg+9E7hpHSS0wMtJ
CrDqdxnXZN0eE2ZXYhkx0Tl+trGGtc/49QayteDzlWNtD6/e/mLQEnuqng+VLYCJ
CbbHtN1IUVMVDSQa3MFGnTHG5I6x3OiU+ZI0gBWZYMoVjvSgxXZyTwDS5UoVdumS
sxLLyxASkMdNNqUYYB/Jadtz/3P74o+4yH+XE442L70hSDrY4nCHy1Ouyjz+0+II
V4aUe4xIDx+/6BCML3h7JuXa94TmsnuUzviMumGR1FqU+W6NpkpAn2MR1+k/a+sw
tzQD7lKVWZaHOqSDDme3MCj5vrXO0K3+29qo2dOO6Q7CRFxnL4fNnpqZTxYG31B6
FahWwGCN8Tzmr5rD3I34aCgZyfPKhz5K0RRJEznik86vqWK6wIxcQZToqlqPjDSy
3oyk6INxeZVg+MTskx7Fe6nGkYad86LtINilAGWO/KwfpumzWOcaWUfrppErIMy0
dgAXAojTb5ipf0Sdhq2GLWcQV0o+e8PEkJr8sMk3GqQR2Zv43lQ1IziZ4elUBqkZ
DoRT227XZnR/DDbBD8cRYilzXDBic/nHWWJX1ke3iZzVyoLFd/NEJ5CPUJuL8dNy
Fd2TKeX/BxeX+pXDcGv01kLBG3VqFPENn+GjBo/RrPGvY5c8aEzmiWwDTKGcILs+
CXm5CtXPqtPo03RYFJmfPJkDqHDQW2VWZUju41GeCUUR+aa7Iu2oKCrykhBaSBTu
vmJiOytljS5OLHKpHFp60j0DCA7qdV/w99zKFnsWkyuLi5uo23ySWWDTQV+xPLcV
EdGMRvUlvAJZehO9MHqycay3MapoZcUXdHw7EdfXUy6fhjuoDkYNoK7UDqe8HR9d
VUBFGPWSrdLr4NFdetUE+4VKhjYLkmfXn5weUylRqhdD4RSIE+TLEz0XwJ/w+WNr
yG+eRPzxLRF+V8PaB7mAcTLqNSzA3XG5ahonr+uF/icwSrSugkswX7U8y8CkXhCP
CU2EDrEi+IGQPUKURdjltcIsVckes8wvPGYtCHlvGslzdNz3qGPS52ruuAkIXS2A
luOYtT6XuTE6m1uyCzauEvYmFpyFZieujjFReiuJcqg6/5/DHwVqRSK/O0CqqtE5
EpPs7hUstMPa2zncJldZS9ixoMAQ/LElaCsZAshhMtJKCoLrW9utkoqWEp4H5GoJ
F9dKlkaIjsBLmScHnDzHRGHB316FyXmqV8lWc9iX5SA5lKe+h7CvhU3Dkw3Q18Zk
dvvmIGU1HysIi7rh7Z7WyGFOPIYUrm3cJiiAZQGolZfOcemB8HsdBZz5aZ9fZ3BE
gDTWgYv1fHB2GhWGJ9LJWVKMARhxhbg4LMLc7F1Pr/y/cEcFsu+kJNHmIw1+8P4J
2mo+WY9Fp7f2P57OA4fIYOWYOWevnjsgffV3/kuveh79BNMOuKzWlQnpvN+HdDQx
tEp8JuULGDU32SN3u0hJgletcMxZujwbbJ+9psYfgPLvdKzcb/Qy2WEO5TSAhzn8
0dWIxMBsdcIm4ogNC5C8mXR7K8V/u8x+F9/doGuy/bO9jpnJygrwlHVZIKPiBa9a
2iEA7ZJRBAEbm1SWW495D8p9H+1xYK+YF7x0SlvXEFXHIjNsGk2fsseKnNcsPPCa
aXQO3+u2NKj00ej7tZMdNIp49iMFbiExQVUDOSkSqR6Is5NfI1oQVWxbB+xLMCG1
xea037i31EckJq+SclhBjNNHYH3cBtgOPEPE9rtc8UDSEgkh/OY/HwEywfz1NG9g
PWsEr9Xmbf6sWcpDf30Ach2EI4oj7XXtoOfwaRRsRdy0L6AMgi/J+VkGF8rJ3UfH
+gNit8yx+Abk8SvQtWNoBw7GAqhXwzZTYVFR/JOI0+xt+3i5ay148HqvBz8L/Kz1
zJH5HJFAhZBQ+e6eenSEWUtkHuw7886hmtPi1lgjV9S4abla/rbcLfaIU40869Sh
9x/wOKz+LS7T+IPBuAmj9ErX+ImlKcbM52SKLoY+/7XPNcKVMLV8UfYWvztNDwGW
etKCxaodWoGDeOAHnmcQqLgGFl+14K0IALVq2AF/QprbRe9ZvuUyLz/jUOsSkonQ
NuEW1ZTZtsO+PhoiUeR4QyCiRTdUZQeGKxtQbwJlZiJzUO1qXKnRGE6+yJGBLr7K
QLPB7fdgXLXDj15ORbF6UDz2b5H1fOmzdZDniE8ulikRY3nuUYEUrCeEdZByv6W6
hEPwgIeXlDQyY3GQsyi3DHgNtxXxRA37rExIZ2o3ugEnYjL8Brosbg/Y3SlAqz4h
blntoxjqyZKrxgMs37PpdGplpVce19lNvupBa+10gbzfqa6N5a/A9YWIt4VWop2l
ibfWEY6x3wvyR8K3yGfhdgq7ffLLm3bmUSlAT5JKJQBXEKZLUqfesS4TE/D4Xu02
vqlLyao+87ma4mabli4p2WaJ8nlz8g7xfDs2XfXqJLaDblC56oXvG/lM5tXs7+xk
Kd2PIDCbQDY8LWQEuWz9+HIBuq/RcJf5ERnsISAICUuy2Tod6GdVgn815qGR8ZLx
IEz4axEnEhPfu7cjrnHkGh1ZhmRACVU+Ewmfa1QNef5WnKjgSCMDteVfMiEdqrzq
oHe7/Xy2E46JZYD90SDeQ4770+rdbhxQX+iu1nRvV8kR8Y7gTdcRLSPaWMXklI3T
48urGjab0YqDeSSLxcfdH5SPFunyrmEqqrymF/+3ff+8vdK752e69rJfcgLqEzG7
XAyd85LfWyujeBOyy21hp3ZFlLDL7TVQtb6sWGeYq8WUatRn5mua3y3QbRPCwpIP
FdHktELbmAg0rofZetSFWpDD9djVSsNuVEWhyPL0ZlTfYLW8WxOAKsKN9Tv6PpaT
g8qvSftHd7KEoqI11iHi9fTGefHfSuA2fB0NbTFOqbeOFMMnuZpvtE3jvD2wz3cb
4ZqGO1izkiRXfB+yQ/1FUz7wcDSsqiqBDzxZTX+laUJVJwhi2UTJkHqBAwkfYBF0
aAp5LPchQmionD0YqoDJXQ7qbhquK0kjS1nLLZ+Tu0IF3C6tqA0JRt751V8FdqjL
26xjC+akxJ9CvyomjBROaBWnOMF1ICra4coGk7oOSYI/1tYlA8NopdXd5vHJpTmg
b0VpncTK2QzjdW2G9dis3thRpgxEqfUAT6MhMAfUNnbXlk09ozE06OWOaaJya/0R
0alZJOxOdMwCS2ZRib9BpE+OGYD7WJdbQdxYifZJIqcpNymDcu/acmIJSvKE9suO
jSMdBSYbFuemK2yl2XH2mZ6YqKdIuZaw4u4LtuYCvTf6CMypX861//IRkZEN/bHz
htS3yvzCmNgjub/wBF8EHpN72YVzo4qzILIkEU7sA1+2MykKfDrVnjslQSLfM+0w
Rf39Bq9fU5lsuwv9+mxyYMSvYgqCDxDIa4JCvSFtvbDNHVmDhr8/nEaRARUhMbH0
N35B18Ftwx2/HiNY9oREGyTCtccLV/1KTVau5QbKiojjY3Ot8mIh5Wengdg+dOMt
kRtQGc/SVknCjKRaix2xca/QfL/x6DyoxwyQHthSouwi1canMfeohK8wsqzQgKMb
x+fS01eLLvCj76lp4hgx4BCZ12a6AvPAyadvS5JGjx1wWYqZgL691C8oxs6alPEI
ZNZ11GCVRKy3S9hQ6KHPsiMAf3nfEx5R72wPftUjwHWRhOrqt91AkteeMucwlWCc
nsj6pqXbXcIEvYXPzc/CtYhqfwwe8b+4N5ImEFjRigRzBiLxtmO/reTlsxwmY+cp
QmeIEWBmJu18lonqM7EKFv/BF+nFNJK9h4HHomoBiASBUm1wijOKFfrpD+c8SQm4
uknRP8faSuM5eEBrW/fJqsvdj0fMBc3p564sGSBmKFuT6EQ6mREQABk7FfMqm8hC
6sAM8GmvRcQ0UpW/AmkeqnbD35ZaL3jaikMI3uqdFERCw43buy+9vfYk+FnN7ToK
UCleueKMxoK2kHZTFd7lDZTgTkf/TRIqF/Y/Ic1NmswUc0te0RbjyA0qe0mP0Ciq
F+YgM8XKrhksGxcun4v5V3u9vtKQhTtoO8ECjemPpyNFv15R7LkKlKGqhZPQvSL0
E6qOs/AXi6OUDomFsrtupdNPbbvY978+qlQlraaKV0+iAk2j4azJK5tpAaWNBGap
lVFeuCcXl3FthfDY2KzuCrPmfgWCi6ufmKvPMqwDnJgagZdRQn3T2E878uUvT4+U
b59E+A0wc7WKG9bkbu/gwe8tc9h2m2nNz5a6bnOCy+UjN30xxiS/RfRBQW7VpK5n
V8XWUYj3o/JsuEy5OvVg48NVAWjS3GiI13jMHG/Bi1dBwplp0Vss4ue7E/aJt64U
XxmJmOgP8j0LUZjwM+Pe2rVCDkXe4GCD/e3YKxpBPngZ5cfNISQZ2NB5zrwlZo66
tVhWGxfAOm05h8KmAB7nQNJ9FHYk7nAPvfSQer0Vai0zFcxGAZqXSSwMORuCvJZU
ItHQn8GTnwte9FDgUKtQMacRrWIB6NTW8KbyxvH+mJU2rDBb/YLUr7Dr6D+05SGo
yqSmN7Wj4b4RLx73ZvVLmzXGG4LaDanlwGei3PgkVeh8ZyuookelfSni/TN+osk9
uYGALpQlckDZb2GvMZTXqHDbL7eA6uGsLPoQqcOwWh4HnMCTAIJBW9vpNpoomHqU
ZCtmCIhFuUFC7IpiqPA6eD9Xp8M98u5HQldYHwPd1PwdZ6jLfee3sMXyPEihlKS+
RfkoIqQFKeln7DnSGY297AvvHHCtmLAy2LvDPbTequ6UKGBONY1aioq8+1RTc1sp
c5WtPq/i5msRH+W6vYYfb9WjSAbYcNatIy3cVwBkxEi5CiOBhxcdtyK6vdLsMTJ1
+U4YXRPwi0ZSKCT63Vc3j9G564bW/MLEDeixxJmYBKj6vOZ/1ILbPN5h266c8GNJ
1G9eeXO0jjPz34lTDF/je5qiAqgkYKDhUNW7b5kA46RGzLBnzX9lh154cSBaJ5lD
YdMJz6X6dul/cloeNS2omPOqoWxXhal0+KrqJrhBjfpHC5swTqCDU7EwpU2WRvXq
t30rPlAsqn5duAVSRGKOtgBTjG0uwwIZP0KDKAHW7WUtFomZlPoSFKe3UJZ9fkGg
7C4/XiI7eFNS3KkWlSx66LTgk508OLpTa4vpEcpgYrWxeULA2Zc6LG3IKmhKlazq
j6dBW/SD3IHBuAcBwIkQB/mb5yC70O1lVMTEfx+i80h/92zVQWBy26wy5MI8uJQR
XbBmgD2DU3P3FdQxC992n2HiePpQvuEnNeKQHJV7O6xAKa0NHyzo+0Xoa5oZYzOQ
37Q2jeYQm8BmRu6sNrKv5RrgEueDzQMgw4WtXdjIDIc+d9rcKD9ZPeBXPwAzKQDv
8VbPFbnrbVX+JT4+fIVf4pQM2uHn+6zHNcyox5+Ki53mI5AhO7ClN+PLQCMlsJ0p
7mlGVO6d+2fx9ZYeyxJqU/JTmhbKRYsNC9Vk5I5Q2l6qWkk7YinSv7hrjT6o4QmW
T3Mod5lNBH1LhRYC7vftLLGlIj9lm2OxUR6b1JHeBRyYSmmN2KgfrcvwvajiMTV/
4/FPNpkLpKaslRYgO8Cr2Uebj7OC1hcgqByZWPbvRE1TDLTfQRPBmq/6IbrfAEoj
+SNElbAFhxf2MWslfQ9cDuzT5nytX4nuyZCB704YD3cxGA2w2m20cOkb//f37j45
Uhy86whNvVK5N/3Qgl2wG0Wj12mtcAPO+AXp6CIWGB+mHLNPyEG6xLWR0nldTxEc
CdHN6hF7kgeRFlBX9Chz4/OgzftKzd/6wq8cE8GQxrHqnStxaIOb6zRobma1aS4p
vAEHDHfPUwe011aYm5mvXgaiMsY6roBqtlfLi/XmN/TSGsq5EuqTqXg5MNXt3N38
mIyZJy3BDLli72Rjb7Vn8o2CsDsp1gaVdZHBtaRxapwZ4RtLDJrHLrZoMXsvKcq5
COUarlZaudKKaoRFB1M7v+MCIXITKE1W6GNxTsdK0BydT4HB7+qbFKs0no6jirIf
S20QSUrw09Qq0YtfHy4RyqRiLqpmHZIuI8YRLUBo9nwDiqVpyIGeDo4CZaz4JVp0
JU84p61xdE+fVJFtczp0PyNDsBw3Uejfh5zMQWwvvPWJsLImNAX4vTLUqI9sr11S
oP7Ba0vjO5UmoMQCKw7ySWBnJfyAnFx3aJYNPqwBf7hen8OFeqA/lcQHW/5hrFtu
WlthXKn3pymjWuxzsvX3GZ+XV1/79UKe0Ln0fOG0nvDL4WmNYa90r+j9/+FAbc34
jwOQVGQXonilE6I5aa2P/SgrumySZRvY3mZBJoJz02PEGa+MqaySC7zv92sVBDjf
J4A2t5gshoBFEThxcFt1FlXRWnzqsY0E7X0zzOWprHprNeFW9aOM+WKZmZQGZ5bC
NW3z2l8he37a5PjGiYraCNJj43N1cnpqh1bJCQEHdAAkVDnQLSlIPFFkWHfJFjkd
e6e9m1P0tvaS265Bg0h8uMEs89gxCL5CuUsf37jkFoKMtjYuk3p6i32E3OqoL3ar
2OQfRXbnU4QaUUp+9lXGFu1KlAaa1o25qdbmkWTg/mgryNHudQWkIWTYKwydeW4Q
DVxmkZ4zV2o9M2nc107owgaH1DS8Tt1jC4wzou9qVwu+2swGycIFFQJ9DSmXLtNV
LDlegcKxUdmEq4i2hL0OJzFmEwDCevJCjMVOaUqYEKElfe3FHbi9HVbgUhsOk92l
BpgVO1ubgLyp3+ySWmQtOnd7KM/QI/HHt9cBllqH7ALQnYrbfsPPhQoCWpybSqK3
fvqNVVED3LoXzvfAT1asUZPj486TcH/n5yDwjAskKccF1aTeWvRnIWmqyM6PNWQR
lQ3Z0ACpCF2EP1zJswcCVVh+4QcXF7dY7tWnYDypxV5zmgeZdBQ3u0sXkzgiPhF7
2y0m34Yylmuwh4MRMZZdG5n3U5GMmQM7i936jFmD5arB7X7Gy/7l9A5Fm7Eqa44D
hFZ6WF4+xAGxZxX8VAwjbFnI295F/jiiglhxVxDLjLckQyVGDWl8Pv0w0bOuYesx
xefZrjhTQxF7GU4FOmHyA8H/JsVBYNpGnNJM7ZT2xSnr/3b4clrnq+KHSEGaaPSN
KFoAMnGzsHRGUkBb2zM4xxXEmXKbnAt8OdAYrFbYbQ5qrW09Ue1zbcKWgBk5yT1O
vuEwgKsw1VI2JAfdNYaAT4QFx/XIWbU71oEFGmpEi3KBq7kKh6cO4B1C7LLwZq3S
Znlr257YWnk0WBpkVD9trSdK3GMSVKjyrpJbqf0o7iV7E6pRlc1W8BV9mku8/NQD
GDDRIQoNCDQtNY15T8IJAvI44SOzrUhkO5bdtAKlMEd8lWM/g6wv809qVD8/4JeD
zACfIxesLaU42bpfkFSucmNPite9Yh7v4SmC1RnbNnfugHp4nMWSiCV/sPyV+W39
qjLkP3gtsxXeXUw7oSObrceNoCa92oLNanV4wK6tkEYYJ623qm28fj43Sq4UTEdF
JKYYGze/2b8E6CzxNntKaOV0sB8QCAdZ9Aypb7caeVQ5Z7zmH7f9HRCoZ4kWs0Ca
qURUgkPO2aOa+pSMwRlxKctrTPwjQ9JR2jy5kroDqNGeH719poqBamg1n/kUidEV
RxBtESORABxgt797IMuz4Q8127NZLNvs39dQoAWEziBJQhVaS/vZcay6tHRB8qQT
GC9pKAq/JsArxMDkar48QGJ5tRrZJQ5PMCuU/AVhY3s=
`pragma protect end_protected
