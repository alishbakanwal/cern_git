// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 13:57:50 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZGsXsCHxV8uhad9WvbHMd8gXjXF5zZD68c+7s/wbJHn7mLI2nGhVk46UO7A8qkhK
DpHL4gVylzd+itnCv0gcAFJvaLc0WDfqh/PDs8jp/7jgXghO3utfhfysoE/q0pHI
sxwP2KCp61xKncwZkezktI6wzQlwYUmVfQuG0bHk8vA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2352)
Xo6iMD2LiymjVCh/WsvsPnCbsg9AJN/eaNM8lnzPBK6Sknb9+gFwXydUcY1jGCzt
3czKet8lTVPcn8NA5FKsqsZJlZjvoxUCrO6m4Gi4UNDKpgZ2/3nfea7n9gfT4xdA
iGOFKbKewxWLlfmjuA8PKDPjoVz0nRxgmlPDj2c0hMKK4QPOD4rbAQzwFXNlhABQ
2VPoxIeC6OklZDpZm8WVC6hGEcozg5xWvkS7vTcgU8mmtTtS7Rl+aM6rt2pz9tGf
sd0ThcnV87kBJuXMOJSVxMLiJo2G7ti42B+8x2MYme8LTiCw0InN1nLXCmuSiVHK
ih2vOy8dNUnz4aBZBoH15jm4c3QwKUKiMG/hnCAd4vb1M1g6adp3Ddh1vwzGNkrZ
AzsiVbeYk5YzP/2ITR6dmq8UmM5VvUIFaC+OP5LlS2cA/4y7tCvd4AoeQyLIBQkU
KYz/EUJ88FzCa5oPx6nWh08k/N4laVKlARkETxmyQzKdkQ2LwwS70EIHu/sabpGS
i+S6BX+xYg3YkQ2Bn0rNF4Ws7fX3puCI3oWWtKGeV+Im+GT7s5mMZEioVceWVhrJ
/uDAw0AYDTsnlsgh/v3pAseOKH6uF7C54aoisemejpya+KZi66q5rDg34bqPuMiY
83FbdyII/0BWSbd1qkm2nGzHnB7iOqpS/AsuPxWEoxBDxT3szEkVf2abqO/t8CWW
/H9ouk2aU1WN4YbY38YMJvTcvcDcogf8DHzuvwBvIIVPnEvkcd9jE3TuRKD2eoUR
hRSn0MmKsbv/vE4xKKEPvh38CrZvNwU1dj4zIUcg1Ar4WzW3RxaolrNjO76TZsjP
4bjLzyrOlXrMehjrCcoM2Q2RG6PFPCAfbIHIRJCinhTdv6qsYX1eVwyeN4qoiqEn
TdMUTQ8R33nvO1ILSHpQJoQ1WvN7TeMLLFD6YaiartpVg7TfQyUfik3VIUcQjTwC
I4WlrolOAHe14DgJjKV6UyCBxSH3WREevNF9rcFRJW2POgkk96csm7pgkzvJ4q7N
VqJPZRaokZKneiCCaI/h/6TxNeNZS63KiLRfCVDOjr+uotb3EKINdTrDRGA+m1X+
fxJt7PAYMJaZgvAl2CNiczqyL8zn2JZqdUjJd1DvYCKuRkRo27bsC6L15ilzwTzq
oEFOFqU+6a1LzXLbXLUNVaxqMaRbGNCbfodLxz+SIso4hAeSkd2CUwTD+xg0lp1+
AgoKWIgRT/g/aTrmZZvzOD8utJHgXvq8Etbs0R8onYQ12CE2AsOw5WOxvJX733rO
hklUUsIqmsJHNSOI8hSqmYiCCxfeRI34p2kCjh961U1qh2AatwJKNGu0OqbI1X6w
puQ9Qlg65BpKsvXodZo7n9uRbG3zlU0xdAcBxi7Fxyk4F7o0EPQ1Wkadlxb+Bde+
8SOiB5KHBM3L2/glS4qzPTlaNi2DDvmC23ddfPqIsZZ9NXPr+U2W1TAvZMUu1XxG
VLzAzhBuECbLyReGmvakEZEiY2xHNzL2jJ+pABb9DMemtjgGK/PdaLXDbHOVs/hr
IaRKBDNuWssm0Hg/NCe0mSgUb6BCigx1vJ9NZWZETJPYtLGAZegJ59S53Pyv60yM
sjgwSDTQx6FbqaSrgP3vEi83YbiPK63d9GMy7qmVEHIdNyGFwk56NvR7j0MqIrn+
gEFJRSNVBbxtmHMFJGJS5WLpWBrHqYCMdP9BQo8Ren4vTW1W1la1xLVShVr1FDw/
Fro3rLtkW0HnJIJfrv7GFgLuLldQInwsMKIpnln8sLxWeNZxVge/M12ccDssSfvh
Q9Dh67n2MUnJo/37c2Zu6Nst1SJyHe/7fuKTbtQXIulDA9z+kJYGSv8Mi6FRMC7Y
S3Arjh0H5kHH30HO4CEK3pe86KSYtcQ9zFoXlNu+d+fJa1UhGcYBohpJxKHGghko
tEpRVDXyNF/ffJKZ5AeITOxrxxTWOs8hXAJBWKJm+y51tewwt6eyhA7W/iO+JXJ/
8nGbrbQ+q8l3fo3hsjhMfZu/CDdHWIVXY2Pxw8/PZt+Vt2zkvKIYrZqXng3W7LLB
DkHxZn0Ti2kEU15EKa5zrmNyO0RWWp5MHAPJGcSFQs9abRzRlMxoVn5C4VgfFV7d
D03geI+jOos4oEMtPMAIrvxsV/5eYxPxqeenzTHLsNBk2sSZBHZbJXK6i+JHMlxC
EW+39JUVuRNADEAtyxVS0ADSZRQvluDj6okF4EOLKpegnggVC+uUyTwdEOg7BQCM
oMERFrvGxie85Enrc9QSJb0NwBMPmZrrQDHXt0LO3efqpwSbrfwLte7cPedIrM8F
Dd97hxYR3F0TWwu8jJmZ3hIVbqhwVP7Sgya5Yjb1FDM5eDDRL21PZEGE5Kuk0VSz
GKvKKmTfh0f5RdUrfIqo3phHnRdy9hVhszy2rI15un4pdXm5F5NuR5JSMX5O/7hJ
HE1pCZCnYVO4yyyPL4kRIDDQQmyPQp9LeFyRn/jAcCL0ZeQZ+oaJJ5qdnniKUAQk
mCjfwHaX+x4ymfa1DNLRicqrmm/YKuQQVNVer63/0o0Mz/xSA69MNq96G7vuym/i
nk5aDBhcKtcSrr2S5R85qM/WDgyCEAyOzxUWDp9rRGzBNcQGRPvemb/hSHLDJTx+
4PjdgG47ORXyGIsGsSkh9jRIIu2WTZIO77s4OyJ6y/xAInuUXC9EtSOyd1x60SGi
CC9QsWib/Gp7B52lXbLobKuO14Ypj35ENQZNJh4uXFBy+gy88SUc0+3e0Qj3vo5N
4oFEY72KZtG16zcJo77OCqCbIkUYMEmat3rDIYoBuIWUC1bakCDtSmJOcV9JYOvb
JC9HvB4S/IXt66popm4bp+ztJGjR4xyKgfGaCyCOdIw56b/pgF1Y1FD9rDluEfkf
tzmSaX1E0kuYc2MRBoVkSl+cgCp39yVhQiO3rnWdsaG3JarDaw4bPifgpOqAkfQy
IH1aZZMWTmTS/zmQtPvyjy48CB+3VjfuwWkj7Dni7awQRVwl54giPw84+crr67Jj
Py69IZu2aLa9QchEnWkE8wr9jbxSnVdrR3d3yr/oziTr+Zv6cRLq9DKe+HhCcMwX
ZbH+KCJaPQRxKrMGWRI9yvLkJkL9an6DdUvNOk/W6VvDD9viBZmYM+OnEtCMC3LN
`pragma protect end_protected
