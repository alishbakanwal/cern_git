// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:31 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qPY5fciwy9I6eEE0obaFalR/Fu0apQQfF8xirJx281mZIaIijxPaDPRmlImZdOPO
cAoOSz/rU+6q892VoCc+Jj6CMsl3EarCdqxtKwODCY0FFwajy7gM73XsKYm2ZGp9
g7aVQMcWXoBWyOKJEiIcZOIjZV6G+NkR4jqHUhhJk6o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5184)
3Ts4GlODsh9xBsGChJiE5Cw3ZR7UaP7F2OurOIHByBIXH7fpd9xT7EDmo68s93wH
zxxuLfFUJFeHMJQgw5Sv7xTkoqulzhEYakzqo+2gGXTtt0upxB7uTTC0TClKoTs6
jbMU+0IeE70Ggeu4jmWVQwbsm5aNk5vy+LFvHaQGwozvSHJkaF5p2bewcIzA4Sip
dLi3BWS8a5HOVrOgFNDGFUe84EvHI2L8UNrkONM5GGQYD6yiMOf5a4PuQOXZwS3U
FusfW7CwDhOgVXb3pxY9TNbdRy0A1GyWR3WD3Rwnc0V/5zG1uelDG7PtD6i7cM4b
C/7pwPDZTsTULqSIYzgStSeCrHSE8sieJlXnZeL5GbW0Z7T0Bpgl1mFk5vSaOBam
b0iB12bXPZrcPnq4LJD9gF1CKxlVrcLqlnIuxBYF1yOJaMCWNzanGwoEIVCc09LY
MuzyCkKCDtbi9VT9aCYi6Gx9GBPmieP/FbRy1BIyacleq/oQLrZ7r4Oyzfg5F89h
3JK7bDIZFmgt6bYXKJK9JYV186UkN2IliA6FKY28BMqwl+YXCmXbXQW31OOK81MD
NWBfXvd3CpmP16sSEoHp+jw58BXAwDOgsY4AxUTPBW/gktmOqQGv2o4yKf8jbuJg
tTcxWK3hY5qrTCLNM1VbWdqeBF/bUhTtV8YCumrrMnow29XAzsNxhE45HSx3t3zY
/mMMm+egAoCn3ZP8hf5oY08ihJgjdBtBI+/b2vbzVQTFnV650rH26HKNFi2T89D7
Djy2ovcM5A1bAhdv2m1jC/bvS8+iPFEpdVBydWuaa79pw5dBab8TMAWFiQ30XTap
Ml4/iK825CzCrveMGsmdOvRz6oaj1wVtSeAedPET8l1V3zBF5RmVU3RDEnAdQMIW
Nt4KRN5SsspzRSFkH9SERF7Lnv1Kpl8WUPQjj7HKhy9ogTytxe0bY66NHefE3186
rTzdyC+ZU1dECbmhCkAegBY+ld+YLLsBNL9xZkIE0dvVG1iEvwDrmhHssYgJtCRc
w5A7IYKzlcQrcS1o6jaYuu8XnJ2t9O/r2kx8YcrX2cLrmXGUy1+cckzSmj7Yv0Su
xU58LUMO8U8qN/WcpdFuXrJxQj+RIpjf8yquQ7Zq/6QSs2Xc0Fv+PzZBBRa4trz3
UVOgDSPaopiR7Qzh0Y0q6+W2u11OiukYuNv1w0/V+VPyAQBhpjHtpOjDnTuMOUpL
WmDmROcAElUYwuaYohqavdHCxBkI1zAUjMGD00HfIdDBJUdrwuUn3H3Er6ovi0gH
ZLzEeoxeOw6UHJVEdVSh2CHMQoZOuheStieXOvRsAjIy2U4j1YokQqKC/pyXaxrN
tIyjzKCVPrUIzzBZwznYBgjDeJtbwduk0EXeykcKz5ySD8a+bfPANT9fqcT2IP99
FIwX9Njb5RS9ZNbFv6ZrDSNRgQolBkR51Q0hh/gGSfTvvJFm/H5mLeb1+1O0etZh
NF2Ins2Kves8sr+74Y8mo4BUvzsGOKzCActLfJu6U7mQO4Na0QcJShScvdIcWvEN
TPBh4UKra9S/2PCHpAXhRslVaPNBe4d/K6HSCzI9O3LEp3/owJojjLxEn+zke6ui
MqKcueyIwVLrPga4KG7rG5MBbJOqLahVC4tEtcHPiFUgpZ26yvIo4T0xMjL8RVwZ
xI1Yz2pYCDVPaZyYJAFn3564ael0/6yxfxl5tJKqYc4nwfdZXA4kvLA1YD+L0g4c
gUvTTur1R/Fz7J+fXgVhzimolo6ZR3d9xyvdy8qV1J/OLaZY8Fwdr1GJflcaWtfi
sPXj3lM/HDJvKWJdUxIT+MuKGIHRWanfd2d1eG+ZGR+LRNMlWFhXNv3XIH7e4ELg
uUC3bK2V1EXlBu+BtkrDL/eXRnJPQ0zukx1pGn2grVMT+QOq85miIjqGeukkw8xB
X582o+Myho97LbzgDGbCIDm5P3oFMRHIu24R4003MMqZdVRVCNh7/VRPdjug0T5N
+I9pvhi7f1vPxar1iq3PKzOgDttxePQbhZ1rsmw12Qkz2t+B7TzL5zRr1vhV+kBk
F14rb5ZgDb7Qq0PXUhawX11LP0G6muj7mlQ0MD3req8bOpJ4jeAJx/vIa5LwuTUQ
NGYan2iLtZFGvPbDUZXFyjbwwAXVcD95his76+Tsi1MBanOniJxCyxlO2kgSyJM8
kFynd7NWitpaoA+BPyisKTxb8x/4/s88RrDWEW5EqXajNQsBnz492Q06E4vA1znX
/n2ngt+kYCTSKoEGP2i+b6a85lUN+4WHaflNw9VWYUKMkaZUVUYTLrRyoS50zCBN
u0h59t/dO+bz8n7pVK94rxXblBul2khx4Ks5z3x3z6omzSsnWUYVLn2vScu4l7J0
6DtJdMGV+a2EQ9L21peihxxhbMmTke/eYH9aDN9pQKFhbGV0qTFG2IAL3Y+RDzut
0a5SQ2fqCbURIHED3I9yE9ZCQfJ4GBIGf2bHTor1Q2OSpwFtjCu/ZIJviLfGQoTp
n3Ez+XQMzVOyr2gxowiPR3A7De206Am/JQCq917/o+TX6opJ0M8QAgkc0tYJXCPB
aWqjH3P5b/48wQQARYk74BUOPs7ra2CBDbp7scIJM9rlt7lIqZWv9wBsoYSyh79w
cB3lLS0sjhNU3oO7839bhGScWqrlsElA+OP2n3Spx4t9fTJHqX2sDpgMZ5/wTyXE
QsthQ5uSygitjBqH4q0B9ysbspQ8WuMCJyonb7eAtDiVmxhJpvyE+BC70WgIPIO+
8PkIUTWURKcTxxeL9M8RkDuzi5/dIDpCgLg11OtYVd9EgAX7W866ZAeNNpt36CQX
Ps+LdTZM0sK45kGBlrN7CarWCu9p5g4RgfCOU693TTWSWGFWuPlZT3kFkzLhp6fm
Y7Sqn9f3+7iJElshpMuAK5DM3UvX3oWYKcvPWwPbki/jHoh/+flssNWrh1L8cQnI
nmgPrl9UCkFKdW1AVI3586zf3PxtyAHUbkoU92i9Kzmm5Gc/t4PhAp2AxfBqD18G
dFso6e/0aNdissZB5NyjbwZiVh9FAaX7k5u19mZU09f9iEwIuJGzfsYdiUT/ehXZ
k33l/nK2DImEq4xxFxg4Nq0NKfCxxMZlo96wx/XYm2e8SeB+IQ+7FffQtYNaLdzL
ZEs9sbK4y39tYyVpmkFGxgiYrDBrOYaJ6o4J3uKT9HLQlE6xdFgvStiGi9mVhbiS
BikM2CmXd8pST1eaV/FnRRPxqHIX2AE2+sa7Qy2nhzD7U0TcmkVprhI00MzbA8b5
cLwuxEMf57Xtvz8qx4iChf21IVWjuswCFi3BHDm70Q9CaUEpM+7HlSEXWgl1s7QE
9dJ6BCKk4/eUSdDjr/oSECoEUoMOZiygOiwb7qGkT2oF4uw1ifOqiYuSKpm2HkTo
wekj6Vhcp4NhEuOlFEGiE++avD1eLFOjdNWHkcGuYyecVOLi7wi1Jgp8fwIz9Xgl
ZnTD5azpA7XNsLcAnS89MKTpl3uGJW3/qMreI/0SFg+qDelyIXCD+5f9t2/e6nT8
+2TUpIeJl2Xl44K4It7uCcuHrnHYkP3PqcQj/UB/6xqMEzDKkDdp7AIe0krULKFL
FueKhZei4bZDpQ/CWWMRJQYHEvUNgT4HwwXLES1tQ8mQvWHXouI2oS3ha+qt9KUd
vpTpBo05HD9W+5ywrwDbHw6Sh1W52Gwyu/LIrpwUCLGx/Dt/1vQ2VwzVedXMVPUn
k+q2TpuJmUC2bVIANnVF6k9BnNdmeV5OB1rUp2rLPI4aiv6rPyISkaFNRFh7OI4A
oIqTtg+c73oV6uwi/GtobwSIvIj7PKtxB0kZG/HcgdKFqlR48Oj9VM3b5iaer2A+
ToqfyFWAewLoJ3Cj3ML52gvMnCO2CrE8n39od+S90wzEf8NejebM3ap80e1wdVie
uSyykJEJIi2PpUNx6VaksvKxumhBWVh41Iy8iXO+vlgPNanRzKTGQ6hIC6Bn6uBB
Jf1JlhIb8kASZgcENLTvaR2tgCeTSAptInTy2Kztd4SYnOretQPYts03YehdAG+O
B3mjpkm0Of5ZUZa+uJfhpm8pLGC2PW7EJCxoTnYSCzKfoNyi6i1YS45aJcrVqTec
CoJARQvtT9RTAIDi43eRxMxmLwwhkatq2Ccn8QguXQp8K+RPzKKSuQayL+xpkXbg
4xLpuguYGkWT9uU8nBrFHwhlEs2idBI2BF+vwzJ6jkZYltsI6rjy2X1EgZYJx7Sq
slstOo6xAlRvl0T/2L4ATD+xrEYTOp/oI9oXZVDDu3DaZj9bh8TxwUFkCitb3kCR
ke8u0eiVATdtuPaj5bv+MYZgkr2clTnMWclOQdlTMwLnOCoGCrf8Z0dvHxSJ4RMA
WNNT22ty45jZ55jDw1lgCc665n41ISdJNvK7koNinHfYQi0LbdzZv09usLsXOyQF
ZzuPS+ljMPDjYzkmfhFMPuyTQj9RoLATuLh6m4o2t8cSbSqdKTbK1LOFGCTTaDhc
L04yhO50ftkhmzPrZsA1Swq9w9mSQYbG+LoHqtzEDod75AglSu+8HaN8jitxQJwl
rkS4Fsf0+HAFi5WjiS05hYrndDS1t/Jb1EVy3d7DqYnQFppqdGuvl6+uqefIRusx
z6Xm6KCbMGamm8mi08uuBH3NuVouNqmgx1VTunTmxk2/m4Ag6xrR9iv7tCpThh+6
T2rO4DgOesrXHr1fMNsXXgEo06h752vrZm+P/YvtykmK7rw6c/UMM8jb9lqUunmj
+urRKZo8gOaFqKIotxKs9sSt98CDwCIiM9cXskK5NzrCQIRd8BxIjf7forJ2XhuC
bI1W9WmTLp9fTe8VAzbx44U7m8m5l/WZgo1H3zxURrKNV0CsYGBI847GP5pjoHtx
NgII2PSOjujpsjeUSUJlL/I73V6D/sABcEVdjmETsWP2IQRywFOOVYSSEeMM80fd
flUUG9txyiipk2LxJdDJLeM/fQOQ1gRJ9D7g2ovVQkEqMz/5i2MOtUk00vyZDWo+
KMNY9VtjAHjZJv3XFmpcYGrCxQbz4uGYOQ7UX10fJ8WfmN9T9d5r/lf8086LuR3v
XE2gRZoQLbB+iGPLza7nCeLptPAV9q2sC4tYXKiZb2OThi6aY//eNCEtguaTqKq7
rcWmW/t80i/X6V9PDC4jLmBIy1iyKu9nCiDZWyIPE2FmfXaC371U9JjEMWsMsO/y
rRLjigRFcwtgaiuZMp4IlUUpUzLNJAcQL7AF0ptgeJ7kYY0A0BUYGaSg8vKi95/L
XJvhoFU6U4ceRTXkRInCdf3XI7fKyBCT2y6vg5AdJo+0qc/1Hj+nWyl5ZBx5IhXK
A8gcnXRXrZaBcEJhqu+YZf5M3UY7A8S/Aipfu11WtuWjTMdHriDnDnWKWlD8m+DE
DPzXekk7LcBIBUr0R18MHd3crZ121NXFGYdoiXf7lJzVN6qV4srvtfZmgWBEfZgV
8w4PMA83OmUKWAt8+6qfDaSpMgZUu4fUP4ynSvV7+vPPRZFQRO9LjJISA1Rwdzol
ItBHx8Ms3xmDdkmOQelnpkuhRmpm5c7sRcnJtRtyBu+9us9RZ6RANVR5FhM7pLw2
LPAUG7bdZ5RHls3bjOGZkspqtVmc7NKe4JgogSbdOsz6GpxOBU6tn5fwCqcSuu2x
cRXa1P5JchCMWtJOjElVkFsuXhXWFfkmGPUEwV6d5PU0Y7foHkS6sToPZr2jvR2X
BLiCLH4sDX2uwN5rWL0evZY+TygwFw0LuUe8r8z0DEfm0dg0YBx4HAQ7Esszp/Er
cSviBUr8WAdhHISKE6sJcf2YYStVGe4hNtOJ1+5aLNz7Eaz3frXVK429DIt+aUEq
36bdo1gZDKfuNN+V6LKsggRKm4D3Cm3rvjkuMwwki5UUoJQWGWa5100S9FqQkdzw
v9reFM1Z8mYRobEn/C5pydzIyzdCnDHMJC9cRocdkQREYPchPPr0e6ZrPkbbPQlk
VKwT1JglZSMSCj1CBRnlH16g0YIEMEGPK8AkMBdBAkPstxS1+Xk2rkFXAv/wjYgi
63TAQ3cwJYk5mdJDVZKUiF5wp1y/UaJ/x3ybaAiEbvKKLecqscqvzn9wUBqF1Wco
G3eQIq3BWgpeqG+YjZJkG9JQJuS6gozDlA4k4tYMfhQqPjnt3u4x+y/QAme/OaPw
RCqKUHcsJTJrciWbCu4H201D/N33cAqx7SZKYyRVhwGODpAMZi6bbldSfE0offmt
EdIhnfw1fnPY188TE2rRC9yDaAfjkCkUn/SSllM5L3ce1hxOZdk2fsVzsNZCH7qU
+S9NRhVfikWJeQ0lsv6sY5cybx3oxmIfadm90ziBVhetxKJ+zZ5dcxykW2M5+2L2
Jc8djaadIx+h+0sYjxo7NKtE8Omu9HT5fqDe0NKS5YSNUw4MPkZcLcfpRzP1ykJy
ic9YBRwKRXr7M1AhO8Tjnof42iXe4ZIoSofcVvpZCIPUVloZWM1kXKRsAYbfRdeU
j540JPeF4O4J2PvLPmeGLiNCLMWhGogPi7siST59kES+ch+AhcoJ3Wf4UjiHzQVE
TIqSr65JONOvGgiLesoFwGiM/rqTvkGMskLLTbNbbaxJyHEVa8XerLfdeXRoHBKD
40tZ8CtwZgWTigoZEk5HyvJYJ3nMAE85xhIfv98nVIteN/y9JXPrLKhMNHYRe7tg
cp/XdWzv3HPqOIMRD75dDa1wBmauDFMhLAV7aDuZlEAwQ9CM/GN/Sy3WtCbYRQCo
urr14AMveE0YUkI0/TLT/OFOa8UpgOYsduhMB7lMjjH/Thmq0ybMa7eVOjVx5l2A
qVT42fHuXI/RxE/e+zzZzq+8T1AR+k30kdptDq/y4upT857pqDKIIAhnNrK0K083
+Acdqfa8X2uiZEiXN8Glv0wX1mtUDXk1TYV26ysI3l+LgmsApFYg9kxV9Cntrfdw
`pragma protect end_protected
