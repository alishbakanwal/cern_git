// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:32 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MqjUquuGIRkiu6QVtpKL8jWGlVfwMnztZZ9QuehiS6VfpG+n66BKqC8vzlZGsOkk
ciDKPwpQw8+NgENxzzGsgMAeDQoqZlBiNpSh3K4eA/fsdrpk3tInnDpXY4TWoMpw
1SBoMDZZrDB1TtTn1waoYxfJK1aypmWiV2Y31uRCzW0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 32176)
iJjYkSxmBRnA2ydyigXrRImJD+ASTcf20NtpDD8yBMo2n14IlbduR0uCit/zRpiD
+f0fdb62TaOBJXF7d1fEwTB8JNuKHXzlNhwcRgIMMVrPbrI7swLBlWZjpM76YUJ2
kqtdubnzHXmCDaqc4GIqlosDGeHxVQyOPzHM5i6R3ZytzlHGd1PKmC8iP8SZSK7F
aHIgmblnSSGuqDzCWdAVecfDnnIU6XlmczsqpJUo38EByefn4esZMlKkrck69VpW
In7pDSgJN4z40LTsNZIai/0kNl2HQclF+UjpSX1u7GmJia3upxnwIOONbgSA00OV
gZJNPLx6laXQXxc9JZuhWzLe/yxeLCznKneUZqt8lyaXAyxyXUosImtedywoRg+c
2/XgZWI60QefO44ZCQA9al+m31N/yf0cMbu60Gl5sDdPphzm9Zs9ER96hWe54Bdm
Igib3HXgI4nmVYTPS8yO5bHrqPWQkVzFEeuXBqtA5LyCrXjmEjHropm0gSEurb6u
gK6mSWjQyBHXcw/29ty1CnNrecaYJTMLsRxu5fmaqbxuN2aGhTVnCTuDlD7DJ3Ap
HtMKrdoriknEjMxY4s1RmknaWV6Gvul51zXgRTrvJopdrKBH0tRLFgWJfjiILGTK
lNe8hNy3ehH1Xtj1u3MnKKj8MP1FOsxaeQOtvG/LMqflsjLx3/fTxG+BHPNrUdeu
lTm7VJEfmgNw+0EHTFAiQ2vi5waVG+TfEdEArMpC1kfo2kFJvmattLS9tyADk+cQ
WZ5pG/ooF7mQ5Z+8cQDjoRgUADZBqrAB75clEU9lbirXu/UnKHzeKCD4Ju3eNFrb
OqDCyVahQh9jeu0+iJpJk0fpPOemsVtCfbuRjQFMQYN2eSIRl4eaVZirLo45VurT
mXMGdmG6WubmmSzHX2ZH2Er4hLyLQnCakZQQ1BYzK0Ak0d3gWLScSRfR71JXj8Qr
8XMnOS/IVmotcL1vjltSnyzyF/D7FFsiaLypEwe1qdfz0TgSHqXcU+NAfkIycJOv
06O8Il38XzYHW5rqRPAudt9JFhxmry8orbe3LUKobn7yhJJH6qNadMMDlAs/QNA9
ZZDUyHUAXdHUJyFRuBmfqGwiyFV9uzQAIsVrJwBFR3PkOCLQT4MkCtCYnQTAxlRI
nb/5OG7jJNEofOqOsSur0Z7D7mfTjYx8BC6PDSQpHkvfpo3SCaeLvdVSSJq3Fo6P
IHpM1K8EyxJ38LqwCB4+gLqloPzXM2TBcgXoUdagOWcBNpFsvUxhEcoAOToUuZO+
9W9SlpEgT+QNS8+ZQhr+709xQBm5hI8eQCKjO6+/waf9uSiuinjQPUP72N+4xexB
Q5COmtwW+4OACz9JgTh2xnR52lwyAkyK89TrQDt0a1gQEVq89+fHO1eb5sS6KRJ4
gTw9S9ASM5RtQpCTdoPcYrDfDSa8wV5FynMSogPqppf6epbCYp0zGVjsWpxKFCR0
c/II/SbLGyZd8dFFVt5CkSVbWwsdECpbsasaE60KeoIZCbeoVlf6vRYkeNkIDAKr
rb/fhrVFR3f95uZ0/ncHGHNoNG/TT7sEhCOW321yG46XzGE1PiTmB2MWmSe+Q4Dw
ZHuDHVr2WtiZB5ohJgVQ9fNdT3180MEuDCiEnncsPKLokACotNtvvwTbqB323kj9
TWX2GUwsQAJkPD9Os1yUZwHZmgMy6R/0R6kA7BdcHeNzpE+t4flXHEue9qa3lJke
ICMK+QaHU+806469Ufg5rTvPA702mOUkvvuHK2eln+Nvv1LsLCpMT89h0rsC47G+
Mta9elXZKxRKgfhnUhN/uRzpH8SgvuFIyhJOCmgwtPdoaicnlS2MIc+QLENf4Ibu
a1c4AGCREGpWdb3OlJrMsPCpYkCNTW/JEDzw3tr8l1ti4pn9+nXz+pKeKU08jyGn
FqtQ7+2Q6wRHDKXcJDD+SrLOtVGo3CzdovSr1j5blMI0h1oFLDfullxxvfwKabkd
Ys80vsXMX00iMMhqL4yqhHxuEY518H3qZgauz43ExdAZm+1Ns6X1hCyGXTlIXM3x
/M3bRDDOY5K2lpOPtwd2b7Nf+DuJ0a0K6WonjtHB9WeYLyBYL2qK05TTbG++wbR7
UUdAcmqBlX0gWnddEpTPjTsQeK/+nfw8VYkjiCMcKa2UKoylH1khkjbRroE2kRK/
O3fMSm7pjAuNs+WZbIyOwa90g9NecQ2ootedkOecBbphPmuocvsuI7iDmnLHLCGA
MoP+84JdVRz1pr5QJE4am1WaU8E5iRzlWV9liYkLFzjXHQXZmbwaQ/3T1tE9v4Mq
p88/nlUowiN3gJYzc0mYuE+mI11qs1AS6IdmJ3Fhf5YDbXAyj+ifIYq08mCVd2Rw
ONQr68dv+0sSkmIH1eeGvbk8hkjD/eudwvqn3Acs9J/spqH3q+VYw+drL6voyLSn
1rO6B3D3qUHUghGPclFcTIo//ZfkVmPtQZ4gMF9KsyaMEZDMOsD4mOfwF74WxUuG
Xyp7Nzx0h/qVkr2OgqsYjZBBXAx5ZpfVwU6KZ6lL03EipNzzEkzJoPlWTkloIJ7n
9mf8Yl07lpVxuYeRZUuYii1Nv6xU6NINJSjBZT6KpQY6nZ8hS/57WVFDa5uOsdh8
/nECndrsMkzFMF8+kLtfmRVJ1Y+WOz3CyEk0AUNY3vjuUOA/IMmIHxSj69OAEpPp
7C/29vdIbcUI1EnPK55ZauNcLwMHiFinU0VCFR7uQ4MNzT7onORKTI+vqTtU9qN9
uubrGwEX+aGFV8jxFlJdJe4YAJ5GYiH9bFDyRc+gr9sluytqsMH0MLTa/DvIQibf
UlEW/fYsxO/dDzRqpNF8hT/6qtAZ7YSaJgB0cSrld7TpM6Z/qxKibq7pkohDLvMF
lyGiTllD8CK3yrltB7dsp9b2ALDGDTEa0oYrT+R8VkIQe5T9ZP5Iw8K3a9YAdqXE
Ea3CfjixAayfnQoaXYdhwPn4Npsp51dpR6dPCy6YjHcFT7Bg5oRLSdFPuRYb6TIA
o9NLgYfRBGkYOtarS3Z936px889uKD7vjTJUFEsaq6HYKKj83+9YiEiGd9DA56ag
3GcHtvPYvS9tPMlceGiZUODIkBl1HYeV9f1elCXkdRqYMmr0+77VFg4IzgTzY4LU
HD4TNV0MRklL2ih7++SyGh3jEN74GNsOBtdJ47hzdQYm1heEG87pF1/lPpHyxUuW
NX/G6Lpzavb3IeeZdQzwMY/bA52Rqvj0XwkmVbxaw7umfFW6paSXcgPLkWoF3MAA
X2HrEuJjgwQnKavk/ko493AKgLhNRY37A13Qg6gJuDG6dBApm8hXBYrMfnA+2BAs
a9ysMrpJtHYmr/4zwMROZsWpo9KNHFCz0eLCEkQg42or0rdWIq4GGr30qoSz1tOG
uXCVfjhmHWVEl1DhryI4qSy1p1MN68vAnVXLXUkQfddm6QObRSdOAN/o2OmkhmIk
2qayAfyeczH57ocXDOH46rxHTSIF9nKR3DA89YHjVqI0jvt16udvRsxPChg0Zcgr
2wgpe8XVGcfAuGXAUg1C/rjAYDc0Tti7jSJQDALiWa4N7lxKdfasxWhJ07999t0I
sdz6HJkwSUcwGGuWpEhN3cIcJML5gtZRn1zYwmXKEmubY6bGRhJiRpgYYjoZIhV4
N28CbbEnkMzOe5DMO5k/KvccUCnQcEzPMlBKjHglQuoJscUlz8RCseOnEEwsaF9v
B43lIbW9HejWuHIaBwkrnNfAwaFYZBu9dDnBrpo275xTUhPxcAcOrirGQkeG18wU
PkX0pVUbJZI0UVDf/hnPsguEJ/Oc1sKtGkFnCFqU4MpXZvButn5HM5WFGgU9AK/P
IlRjYFuDnjnOKBl6ivsgxFfq5FcJ4uU0/8kb0Bl7DkyE3Wgl1dfV+gkjuaZE/zYs
ZNQmEDNtZfZcabN3jZbEaii53/dvAiDUJl+zuW4C6LJS35sGI0bRmh6DdJ60gbW0
cNtKYSuOXDPOGhMqxl3xQbhlMuFekIHXQT74Uh8GBVo1j0xuV4OS5i11MtJQMTxQ
gxKql3pzxmNxdCn09CLDxR2SVzlM9ROZi1x0uUFeQOmj+3vdU4Dg2XIqTUYq44o2
xIwuROuvNbQtYct8Z7GPPNHGayRb+IgA5jKo53sQ57//ty1xtMyMvBg2en1jf+Uf
pVRL45U4Py5VaVifOf1LeF/AZzttGlhU6MSe1p83AqVJoILrgZaOQybSNUqbA1Mc
ZyV++heY7lQYC/eOkZEP8xtt7zqsFHCqkPYD3ho8GCn3wai77gnKGunS6+P8XfxC
+TcuJMTD7XaUCQ3al5ZAjdEpV850zPZTAQbo9XvalQi24Jb8252XLDtTLmL6Fwzs
BS0BAzDrbSi29lTWG1y+y5oT0m3+6KVefoDkXTpk10gAP+FokdIPyLptRgTyh0HM
eBweI2d+W5dO9qlMiwteNKCacZbEYbwOJBjOtG7OumRIRFezCUO96fVKb72ZuD9A
jt16JyrE2B2TYcXw9JkjIQfztgrIdtw38Es3Vghj5Po9PPckNDNG3nhOkwzTbMfa
IAIaIfyFS05gNggTXyNVvM4jMTj2Sxb+RTyvNPFmoDmlDFb3mJXbBzuql5bes/t0
chE1d6Z8klK8jIwNAOK5wna6U/BBuP3CqEiP2lmoNejBqH6vgugaZSYYUcUggCW/
9WtyOQTwsxDZS0m3xA2jJ912RBnKXjuF3EuMu3bQiJqw3viGHyGe16FCL6pulDf/
cPNDNwPHWG5ZZ5vTxCLcTMyBYLbhfAZvO/JxoC3kPVKeG3HGXQVV7tKNs6obX1Fb
xIZurcn4kI0W2go9TKl7+ZYw5cQdgUPnQlLNgYY/suTi3KTpr1Y89iaIlqO2kmI0
TujBkywx1QZN/0M/ihlySdG74Qc9xu3OGy5VmL7SbT4Mt3T56AZ/11ZBCBSdYrJy
ftz3H6G1VtIa7VSz+DCD3eG3MmnF8+Kkbny/I+bY6Fl+0af9Ba04V+uiCF1AM4vU
ZhhZFWnRIzojzscQLzhU7l9UvyIlh2PfgLW7qZj79p7VE2LH+nMYAXBqoySuXk3B
nhEPSq+A3+8eMwV30LqVNMLsb4HfHEKfiR2/+DOi6zYK+prkmbDmSFZVaeiusHpr
3GKbLBoo69vtm4rb1CegyySokejQEUFTniJnRo8ed/sLEwP4QYUUv/FaYSb4RJAl
u3zL1HbaEkA9lsOTKOd/p6fkHyHBfTKlJNbdMTY1pI3Zf6Xii0hvhPZpJhvdhBKS
XfyTnuuyedmf55TVBsmF499IJysTgXtgDfDFLo0kHEQ6rtg4cmjaN0XRqzAgUaff
fl6Qo4cUCDBBtuCCWQHQ6osddjzdNG5jFR5iIaB+rE0p+Cj2IVVxPWhj0iGOhpJl
Qx/YrQ/dRN/WMSG+qAEY6IZqjMT7af6VD+3RYWK+cPVwVs3b82DHpEMek9aZ4aaP
JIFko/aSYbuwIxu6e4uRcFHZ+odKHTgYQiTnlOLWqJsZlqhQWbEBu4LEwgo8Iokw
GlsBDczDXzAG68eIM5BXrncf9pp2bmtXz7aEebaOm+/3Pg8x8xE4O5v1QdzQAr5w
NPMfriw97hlmpB7wdy49ykiLQ8KLw/BByvKeZjLhXQGuiCL1qIO2PHYTrcrqHl2U
50SIkJqv/nSmrBJyrVO9JkrHpy7Z+u7gIuxO/Yiob3qQdrLDdT6OVf1A7XIXYUeD
IALooe9ZylAGD+Fya7V6aNEFUDirlqB/1GsrGhwJLlipMcPOGcaogKc+VoZvjzq7
EO8+/z+NnnQfI1CWIZPiboqC9H8azZcjKTrYySainujZ+PqKJyM9JfcaJAmjgMsF
69ySx8yj78LgkXqZpGVJ5w+R0bP455Nkor2ak5UMD7PSkJMpcK9q5iYwpoNZvcNw
rY34pwBK1SpMP7AUZLD3JnjZxhY9TsrQvpo54ocKvj0OijCTVVC9Gmyse7HYewV4
/dkRWcV8mp094rGR1WpZBn5vfOaxWf0tzf14Rtl10sd7jpTnH1hPt0II03XUL7+W
3jFDy2pjWUE2tIskHc1HvRQDS0yOz6c7Vn34w3h1CZTP4IaSqrH52T3Hs48+s1yt
klGLitm80+QY2/QzGMM68fgf8vuinJ625pJt7VTfK+zAZRxfD/kOglDGxFjgboRl
ZlJQq4mbxIwuoWX+yt2CR+tNzkRXZP6V0JkfjRH3BK770ZaOb55mxs58rKdgb+hb
Noz6h+zor13+v0S5oYFOZkelamvhY+fgDjJ2regKhKPIFIjetv3ohvIHu1wtyfBr
oYq3QuYVL1k8wH5pO/IMPDL7C43dXMQm4rtZXxTazKMr63+qM93wix2TCuUZjgrp
7Rbiatk83IFWO/vNn80MGMpPsuyDfxhdmVHFkgEeU9a/4UaCJ54qzInh0oEOVKFB
Sqfccq1uPYTlgz+dXyeNoluSBKAtUpTuxdvkubgwxE/N6jCi6rVHda/Xcn6Ewx4y
fbis5qs2ix8ozfEG75p+WegVLGJkFv0s7VcwYWwMJoJ36pWoeZOBH0Ukgol3SjxK
QJBCJbC7c/N87QjjdkMiFudCl9dmHw1kDBAqMLVcdE27yQGPWphHy3GAK2p0Fw9e
ZVPY4OBeqkgRL+B0T817BXoQe8Trbk2LeF+H60cVBAhvEBR7/dXX13MOAiQ7BGg7
mVZMnVluuhtZJMP/g52v0y8Cszdz1oRJflAYpechfracHoNDySyEi0fWti1fj5/T
pYycFfMjPB6dKWOWq/OWp8VbZrDQm4LuPCWwf2HXPN2FMBJJqtKLSkargY0wdTk1
fjB6pm0JFPhw4Rkc0tF050xsuAXSx2qlMVICH6swIhnA1NdPVmwpmuVBCzMLqwMT
fecQzLT8LA48Dy+RQCEOi2J9mpnfxQyOiwfW9I3IpMoLFdSuS6qFhTCHwsYqEGV3
7jLewCv3IS8ht98VY+ndLcWX4EWjFpbz1erCOYvc+RY96VjxXyaiOeu0G2/SDXi8
5rfan+bHHHCY92fKgjDO+ebWFUPJfiKo1GlR8ErypzZNjF8X1jb7NhKyn3qxkAoU
WyYNMQ801NR5KumQcinvWStRT1P57d8xbWsBc8ZFSXM5j0QK6pkOXET0Nys8p6m2
VwxW1GUpzpR5oW3b+x8wHhqUfpvqCobEpGL+D/DB5t9zWvc/wBwIxK4O5wllAxgj
soDbeZLehtAwqV3nXfpPU/1DXQJ+f9+9wJQlTAwe4eP2fNA3zRQtIsd+OVWIsVDk
ne4rAoIyK+tQe8ubGoC2bVRpsvETK2fpEs2NNog189ZCYd4IyF1fipBpAiN+9ZqC
Zy2w+HRWq71hNWN1yj3b7AHMwYcO9icAZ1Tsv0DvgJ1Rxom0ocX1NhN8o2T+QJWP
a2vD08y2nvZfZHnt7rZ0eXDkB31XeqeVs0br20MJXdzUfKZc0s+2BobU8fVx0pxu
mlcBZULPGhJtDlLVRnyDK96OZaZlX8bMCLnNKLSrRX73Z2VPjErrB0qbuevi3q1n
KPhKHhSLojNx9VXj/WQTsYEPlX6g/gWtG8npvm3wmW6/XQpSqU3xBm9MKnQIMbpk
vV5u9wt5tDqoNzODFepLCY4o1zfZdUEDgyvrgG3pgEyRPRCEHElLt3F7ho0ICLT9
bGkf4nTx5LOW3ngI+Qw5gg6PEFYw7dtHe+CmdBuOWA/X5k5/KxBhcE+ofi1g6ixE
EzTnhDcJ1XCx3MOeN8mUj6I7F3Gh1EebqTOIHkPCbEMGFoO2447Tod5KYPkXg32C
7epmaeLCb3fpKGzui6gHJa9XCBx4e3MBa6B6uHqz3tOQlj4dxhk3euFVHqmgVuqk
O0OXhJJgzrAdlHNvqe/kISXw8Wdxx8BIW3Rlt7ba/w0EnGwPoqkBJazyAYbr/ua4
DItsoR7LJcYStQ/CeGHPVF5qqE77zjJvTFiz5CdKLNP1tBVgze6miuVRvOi1cD4C
2EgCoUYy5SgNoF4SA6JyqGHMH2EctJZExSa8UaBPIc7u2TaC/SBVlGbW6tFP+wm8
nSJTgDHz3hKsFvUZOuTAx6LVBAaHMmXe5i1XzwXavy5X7je7qpOxj5yO0XGutslx
M7VuAfHaxyqa8uQ2P8JvhmhjstBLR95eOFe76IrwmI5KoQrx81So+BUM3RToWv9I
u2m9hduT1GMACMo4rndtDvAN70BcQEcdfFNvNYZ9UExa3a+iBnZl5V16R//E/Xka
nbjrJIMGE+7zS1iLhHZart4JQ/2+nzc2D3pJy9HYs561PK5mHM4ObwQRA6RhhFuZ
rkDH+v8d7poiPuyIOjocbC2YoRwMTKIyeum2pbvZ3UuG/kD50eMKUvcuIhkV0l2m
IVSgLSMe81e8LTkHoBjaLAEUTNvfj8M+tiwjVIWAtA9EJm3mwX+X86HY3RFd9wMf
u+xE+U2B+gmkFUMZuRB7HKcxyEwiHHtcgYTGPqcB3z//yNPwSYHEjiVj5RR+taQ6
+8Dw3WdWh6FolUwD26jBVt8vM35sxo3yJ9czKqBCDQ27sR30y3E52cnMTotKIrMD
qZfjjF23+/asUSVuNj9uP21MSn7libYXvXsenbOAchuMxeUtml8rLkz7IoAj86Qd
FM5ymGPIHvKNdbfFe8oJwAITiSDccFzoBR77l5cuEiZH+gL1inPThUuClggVDLf6
w1wL8OVax/6xA4lwLfndMQgxnJ6W9yufVAsyr88YxzrbExUo56hBGL3r7KSR+3Js
HX3hmFcT+OBHNjS+q5fb/I16IWaZj8NIv8hjuUCcxoZB+IHVTRXWdOzXzOTTmG9+
fPOM312ppbSYln0HJkdoJy/eM5uqYYuftscfI92ud33uguv/Dleflj3vHcRgb23s
ltnD6ATydrsX2u/zBHW3KMwJyd81XODi8KcsUWIKuo2VbVzZbYS6cvizRB/QqoWF
yO17VoL6OhNdzj2YoiUlKAHSu21yjZfmwiB8UdghBsko85iJHNSSw0FVUZnZJRv/
EF71GmlVOHdhrg7RmLmo5pXkXSJWgbgBVZ2xEV22dgglkdPuK8j70S8qGiRAoIxU
y6PeTFiX9wnO5o7NH2iqT4zZyKQKVgq2T/mDENWgHpjj1KeCz+H5jIjAG8mzJAHl
F0aoCpookWEEkSKC0FWWknUQYFlV34sn0IcZuTAeY5VYIhRyoLqnDZ0Wn69qU7Fd
D3KwcCvH4ti46ULRvrPJaL198OLbA4T/9/XSCcJnbxVB05bHe41HASX6zMlth767
1pRergX5P7JW9Kx1NTBbcgmiMMScaSa6htcE4mo6Yie6k9dDY5il4y6qvAuIpN8p
00LGuNDFQtOKZ5111tZSLKw169oT6pecW+ZAgBzzDrcS4togCLra5n/uvjFU2gZp
XBV+aWlXFEJ0COJtO8xDbAQZXj4nkhg5RbR0Uz9OxG8w5QzNO6UIcSwWDG3HxfYY
MFtCvZpU6EXoB3PawIxY0Wx7agOjFQRUcd5H8EV9uAT853uWsdsbn0ndLsjcoh3R
ZjfvFytcIrfqieVe1LGI2PT6FDAwcRmMmNBXgE3stOZycHU/gd8Szd4VHS6RUMhf
t0brFb/bEOzzcMgilobwLC2CaaEToow8JmZM7DXTCKDf90UEtV1dDiYVhFVH4ZtU
C5jaNQjRt5Pg6/dqkOwRij9tXvws+KXcfm+TleWMrfi8fPxVqcLVM9hF985CY/Lt
hHkNHiVrFPYlTpCJvemka2JhmiA7/Z4mLr7WPRb9762uWT0Mv3SO2bqVCD3HEzFg
Fl34ohhGiggwiV9wKlQp1gMMkSGjyDU5RIAOTm7RD4Zp0wqcfbB3BCHjtG1EoALO
bmuYrEZg0q+zGGio7cCQhAZpbIVJaSa5BydT54H3baZObJdtQiLg+/x2xdF8rFEm
vfKaoLluzjEvvGQdc8v2YVyAJWOZb/Bm4pW1diHdbjBu8qNmb4lMSjBQ+EPUhLjZ
+oTp5tV5i8eVJUFBtf+zhwXoTEyHl9nuSJNqr/F3rhbUT3N/PW4j1Z3BA3ZEdbPp
Yz6TExTeeKIQgXMQgSEH8/fXsglQnOga37eZMf+rV1BVx1dkUfS9bWeIGJaqgaeh
96mILl8+AiN70M2WLbik24t9la2SKhMXWmTCA4lspts/F5+FDfTwTA7GJJjCiNoZ
LM4ySnu6z8DFQWvrnKdWKjqn6KqrYa+UQkx0K2phq6hgRlh+jkyjMbPcjvaHOx6e
hKkRYXG8sYAbwQE7tZ0lB+ojkJfATmiEgtG7JIsymPFEMqjQcSN51M22O+8mciI/
GVi+X77OSiPZAfRPGvHE3AQ6JfudphJlgA+5y4rJyuzAKrkhmfiRFJIt6GCk1go4
Lqzqv8VtCu6KUfBnTouRrwgKO0fahSL0mixfbqHLers+OQOX7Zg94uFXvh6M+OZE
RSSvQfzwAxlzpulbevSeb4moskxWALqKoPIPKnX8wbUgYKGQGEe4ytISj/bbi5SF
Vk7UvQSaruc479MPX56/BGaS9lfbCP7rYhgCSCQY4R/TPKF6hkKrdeRgwwMPGPWm
wSghp1kFI04W5ZzKY6iaIH41MHosjKzOUVKWxyp3fgoMYrsO2bFUao8Pp+rR+Ra3
E9ancqukHR490DcG+E4pwgsYiNjvr3DmUca6kgpbtlezUzLn1sBu4yUwKs78Er69
sHRbGhD/GxiNE4yYR9R7bx5/JTY5Otl4F3875BRpA/i7m0wk1hRLb2xwJE8V4l5r
93DlT7bpjmpnssAUu8issasW0gfeR2o55pI6BIVGMehgvKvVFAcUMt1ztbdMEl2f
r/k4vPqT8lDPz9Uduqo2nkoDxlHuo2VCCbImezx7QUBOqgk9c9VBGfa384iLFDg3
FyCaP7HCS8a511DMj+50yjmAauu3uayj2S+C/2dySF5gyehds31thVeb/k8NAstk
IMLzDoCAE+wKkJ0ekj14PGqJy9BGlURKPzRU6gC6XrKyUrSo0Fv6F5LAuuuse4ML
W/KAeocp7EseoF2Ii4ri/HmA1I1X0h8v7IFErhVKSp0Y/K6BCEkaZZJUl1oCwpwU
m8m1jL/lB8/DO0lPFk2MQVCs2/jG5YIx6Hk1MgvI3iRVAyEO+7ddPtjvmOEHIy0x
nv065VWnSc2n30Z8NejJUzGQC6bitZew3kYsW9gAYKZTmKZ5LDK6LSco5a4Uh2aL
U81cM0kr3cHslRAz7QrK26RUI1P5CRQdaIODSiBGmb4909gVTwgtTjvD4PaedAIw
cmF+fedZAxrth4wiLW63MknSMytC0/K8VFqIiGzTR9HiiUiWfUwN2o5rdMJTGoU8
fCX0HsvgUBK037EANMkzNhfiGpXX66dL1zGewzY6S2U3o2/32wutzE1N3PA29N5O
uf4a+nI2tzfHcqbcNcipgLfU+OPTx4HGY6YANyaJxVDB26w6PhmnTKKL4GiIBcxv
no0V/+G07CcT6Zf7kSnZjIx+2KRFreMnAT0Th3EX26nfIniqQU9X6XCQxNRaCAd0
6Ujo3PWPx4KLV+ptz8cjGIfKIFzf+bc85HPNSCuXamZaAuiATz6BD4LLPyA3XUMA
NDxp9j16RQLSfISUFt2jITbh9AKp0OSoPiV4smMjrw5V4ToGAUo9R2MuqmvMR3/X
wuX08Q2l6DpBuo7py6miuoL3FTmXqpTSmXZ833xHlP1id9YunkUtH3uCXU79kSeh
SNezbBqQbxq7azR/R66kyVXbEGAUyWWg8Di98+bX9AXI/Z5b6kuaqh6rtZpUCx1J
ZfU41ilwRDnDKqFkrISEPpNQGA1EnkbugibIbk6ZjRsnAV6N4sa+WVQxPdDhSaTY
0FFjyrxflfhg/Ziprwg/DnNgsG0IYk5eaWYDa8o0QOGSMwj/783xT5Q0lQ+pbTl+
509pjkBMcwvx4rme8gwhO5rLIS2OZG9zS+Q7cmXEGPgan6gY9PKWmM7N69jGTIZg
S7SRhNt6IBLldP7La0YmcqpyIzuxxL4Omsfmd+cDaAFAmW+6lCotaY6pK3nyBFRk
B7yXt15xCbYjczOXm+SwQcBkuACht8TvkCda4omaxkYioQTuHfXOmCsrZShlw3Pv
uXSX+jqjzKklgAZEB7vaBGLfmZ+fOiQ1rqrb3zAz6Uz6kUPKn6W2OXle4dqw1/vV
SECFBhEwVuKUaW05YebsSLd7rGbED5RyRD6pwYQRAlKJkTiSJztiVeOAL1+hRHxy
O6qulHcL4SUQVWtwYdelC2A8xa3qsdUH1KUX50BU2CJ8rztyYYZyQI1DRURHGENu
lThXI8Q0YABnWYUi09O1YPsHKFYTjf0vgSCgPskXIdcPxtYkc5yWf/nkLokj5hie
ba9MvkW5Cre1ULkKUHopyaZIBEelQzImoz/1Jmj5oiJBtcvGPBDfCzfv3cffVRi6
62DQVCh5tCOdVYg2p/rjlhO6ls3/AAz05DWDNjE+jASOxPB4qiqLFAZI+ueU2gb2
rRUJutJ9OYrzB0lvadNtEZIhIKCCzlF14/jOk0Odje/MZBk4p/Crna9a71uQYqiv
sLKtm7taovTz846Y8ujmLH9lcHoTtPg1oJSGSItwhv2ucsVNNS2SkuxlFr5MWE/A
VE+FCdKxWBr9FuObASGGbAMBbIS/ELeEXe0pSeJkUwE2oquIZ6ebhQznqIMZZ9+r
3KskjOk7/REaQEWvakYYtJWtVKMuRNdwdu7yB8mgXM+eZ+OY0LgXeCGEDslDPPj3
84I7QMH3XI8IlRvBEim57gMDhAJUr31SBdqSrQOOEQCD1qlXsiO8KWaALpgovhNX
Kdsx7sHJaaIy86dMaWKSjxYiDAJNXpncfn5bTHLEN9tk6tgBhu7OmlozMVGrKnZp
ySsN0p/Uxi0RgfrYpNX8GK8w0AfSNs8BE8SEaZJev2Njp4yDUIiia0fWO5LOkCBC
bVMTdahSuc61U7zHGIa5+3GMiNuUUlfvZdRamSpewdij9dBcidODVg3CNbQim/dh
8bJwXJnpRpA7KsvNK5FW3eV9iLsbi5zLp33MZOIx2gA6qMON0laBPpFeKqV1YIwS
RoqlG5Q3mJs3qeLBntboJJVQUgMu2TQA5jIOs2WxibkH1cn86B3Dn36rUKP0IBRD
B7kQ0gG1zjlXJ5dPsuGMtl3JTlx5fj8wA8Tx8jNig4TlSA+m6OF+RzRHH4Lr8FV7
oLsG7VExB4NfrDx+F8ikJarGBja+haP30tImN4e3thhkDiMGSLxZfkthHi39eBxB
4xBaWAbmZJ52Kfo6Z9UQICuuYKEIfavrcGROWibf4Uny8gWSW3qjWF3fWf+YIZXP
PLzR/3w/lfToJe+LIpcO8+m3nibT2PHNEYbeFHPnZRgVdFfcL24fAbEPw5/qZHXF
ExUfkt0eiNCmnJsFAln5YzuEQXVOE7zjj+HpqyORKxVxImILZTWor3NmA8wV1/IL
wtQ2Rnt1s13ISpB8AhGdMs8iYBKhLeOebkvkzdf/ccq/0TVDDLCZIdyOWcm35feJ
VG+NCcAR0Z+bnPjEwLGuTjfw79Cj6t9F49/KF+WrtWKfr70k2CxMvegJVeg1WZJo
I9vj+hySsTL+xOkuG64qLe54QC9w9OrhdM2D4ixrqOKHffTQ904aIySQogmy44SF
5HN3Jwmk3ZGd4KaJ20Su4nThvM4PrfhhI7FTP/pR+aE+GU1T6khBVSSBoRMxRapg
YZypSj2tQphji7UkkDUDq0TkD3hu8RNYkOs5iyR6PwdQFPeKOobnJT/uR/1sqnGW
uoFQkGObvrB+8snjA1bfZS2/o7oyLl++o33NSLygPcJisTOdDP/R8fWUw+wy7/g3
JyVUAtOu+VMaYRZAbu7zwFeP1/p/4xMgPGpf5f1vCvc6tfwmxADiWWaFSZun13+f
vQZ+/+lM8InZqvxchPF+gfCACY3lzn2BzTMO/G0WI6EzDo1Y9HqQ2oiULfvB4bLJ
TsA2bn9FfWdvpq6TeCMJf/IjWJeREcjSBaqQnZ7eCDwwdQRrhJlsnpAEEGzxkuBv
6b59GWJnvAO3XgJZpHbriu4MMRkR7Vil2Cmjgjy/0OdMbGCs1V+4dqEKGt82uWnu
zSCvCYhHxeP46l0VeGSlhINmJA0g+lS5FqKNK2b5URwSC7O7ymaY/8/qGCk9BVw5
YhOHayNaMdIfTqXEcUxt3GijS0vg20rFVUtsRRTUr30uwmwrFfD083VUKMgcQJmL
8tclVocffIdWCVDovEmPsNSdcB6ZM+tHkiUHp4dAQ/IPlukBd1m81jQggTYLqDCS
Qxtc7xuMMuRxGMiNwIE9VMw+QU1ffApOAIDZp/hP8by2uFY3rxSEMABgLXpXkeos
Z1atPJdCzesZ+mlHC68F6OJjd/4PF7inRwb0HcqNRHehV/Kte8KiwigI4Hf9qI8l
r0sHD0PfboBj/Exz2TqJlOEVtWh8ANChQU0mlRwkWz+T4jtAxU81f7qMOHcm08f2
4+9VLp3Vxmxn/tqWzAL5h8cD65BoacoVsmkL5zzSgRPSAnyngEzyervYqhjRf/Uk
N1yY+oPEmTDetfOwD+tZ81fEnrJ4LZVCMKHvFGm3GBbMIrffZEpsxkNA7anW1kLI
xam9FfGr65lwPFfyAlsEJw4a45ofszL8WuJyYGdeVtQNTKkLkZ+tNkJp75PYf1eO
Hck2Gcmai0Bay05f5rbyPya3lBOrPl80vyKAH/ap2JbHwag7y+9/pfbcNWF/qODO
eWUpQM1DCUs2Wadgljm/uLTqHroHO8WQX25ZZVKJXEZEvk6jYfP1KSFRNaW24qSX
OqWBzCfMFOgiaispsAfMWhSHg4UZA16M1b4fkQbZaYN1zlhskDNzCDqaFfsGLXaf
QfPtqYxO24C45mRSTabFu7qk5AYcBZD8hiul3DQWP76+ebQXucVtEZ8uZqTJ4i4g
Pb8+svsm/5jIhoDL41xH/KTeuKPu4wY+d5bHiHemLgmnamtN80+4a9B7vfCjVfnN
b44vvkYzVUZ3e6pjZvPvGrgufN2oNg3Ro7PZOoXQn3kDz3n6rh2y5IJHSoC2ruoc
ARfaX0fXboO6N/s6H5zqvaV4Q6KUJxdIqIIWMhyLhv3Bx3bgkWAPvbBuZNYvSvKs
lKLkkiOJ7Yj/+MNjpbIJzTseAlnAK+/s4t2ZpSqQ3JU+HmGkJ+/hUFe+6t4U18/r
Ogzb9jdoZGBO5vmMdCbBJCN9eNQoCyVkEM/PZbD2Tf3KYQP1JlVlHLXBO5mo6GM9
mEtlN4LXdrLb2u4NgtH+fpCpgR7XRVS7p4kiUuxaAdfOtmHbXcTy3xLlzG4YIiqd
6OumlsYUeWEkkxOaw/Siz2Td9C3OdGjdA+lrwpo9rys5oinXhnntS3P2ULtjDzkN
OiEKpZwGoBTcLOd/UWMXCTLIWojKwdlRaWu0tfjLsl7AjclVGpG83r6nn4KFZdIs
jbSBDl6YobGFQ927iUVekmu6ArYJqnCNzTW30EKHvG/GES5R10yfl6l2QWYS6vXL
tPisXWbxlj3PbxMfktYDR7kwijgYEwIm5VhelZpz+D3Y4neoSU5aPcAv8GSuqYZj
/HHKC89LWunIuvC2a1jidkpJsDd6B1+ZiVOqPDg3qp90lL5A2h13br411LyAiyfn
bm+jTSrvTbE8Dc6hOnuiAnN/YeOEGCaOqJFHPYONQEuJGeEm2alSh6UodRevj805
Xr9xPPqzpg3IejXEfrt5cebOFO17fKE2m1nj/Sd276sV/E/qmVlHy0d8CctZQL9f
w0TJNm9fXzDRqB0GC9yMtwbAejibAEXursvJDQ75lVPzZO4G6srOYonPj/c7kjtr
TL1jCB8eoeJF0vLB48YsgVtLGMr/BhFv1GY60sFwYuLW+gawtD+kUYxQRnayBAVn
PJAyAvdBgLIDRrqLi/kXpbCAxdCKJkNG0jSJIRX+Ck/5FYA5l/jIiuF5RVicfdYv
mjKAU9fEvj54QU7u/MMq5iXEKwq/cfIWyCN5+dM6PIsWYHoBZeNrcslAQCiRXG0p
VTWWvzXakHsoYiLV1gioJh2GicHvCRfukHm8HzWLKfigkCQ78EUu7+7dGxGxmcCf
2j8YPkRys9r4bf4v0VJBWxIGVKtDzvgU3FNDlt2UGjzgHinAq4oMdRSmWqesKd9R
nywrLz6ZlYmPKAbVsDTvSdirpc4iMAc5RR3VxH87f7QZp7ZAfSMFA5MQlY5WB3+j
4Io0Cp9o9M6KDhjdo4yezjp+wqMHImD1uV7ZSqCYdg1FUroB4N8EMM0NbG3oywBb
07nWBAehd7+EgCkO+Y/YqyOI++h4zs5EH7dldrM2LHnAbcV+05Ze+hR9XWvdYQ49
CSUh0l3YJMembhGZdULMc8krczANgbTAVMAGn4Hm4dOx3i/cfoHX42Gr47rpVLUr
KFDUfcuZMljtDhxURkCnZuG8awwtGaT/GlNW7JezEPhxvKQKtqOKIBOVZoa2JI32
NUWInSsX5GjwnkrhIbjFov8tQJhN56nfck120cbPeCjVJBcWyOz9B8qn7hcW9dgM
lwH+YqrT1rvryHuafGSQ0j5zQB9JL8vLZrpL76nDnmFz+Oo6XDhLw3vKF9B6oVVN
AvbpwolgYv8NuPuq+JnyfylXEgH5OR0fLbzL/SD9EcxKAkc/Ha6jebLmP85JKL/2
SGyQdN9A49gECBanFIrR5dsayBx0wa2ufLD3vImQx5Jel9KGt26nrGoQMrR73Fe3
vgJwNmtXaMaHTNvlPGRqaxHTjkq0P0Sr6st72IAIGl0kHGHi0/nsIaTO6FEy2sZA
bI1UNJkLLDN+3NAPPnQahJCv9hEqpc9JJx3sG9rS4q3kX06o7EeLTkXEhpl6N9Ry
aLa/mRCRGo8wqHJ2XhGcu/LkRmY4Ijm5CkNxqAQAdQl0gdspjuwsBsWtshY/8Elz
f8f0T4yLP9zSZGnUlmTxgmGpAqfR7RpVf5M56zxKhey88akth05xFJ/7Rp2p9PEJ
09KV9THGuiTM8CPiQJSuiplmkoulY4k5FKUV3JFImPst06azdSYmoYjOlJ8XP5td
p2oCaBGNAzGeXum8qS8SBurx06EvfAWe3Cz07M0QPSVvJpftdTLGebraREh/RH8I
W56t1tegnNyMYFcCOyIvLSPKoM6x4mTzAvnAnAsgGErLTdsBdnSLYygNqrQ2m6fb
jCCXgdvgDGy9h1tza1kL8N1aU012HwYWWJCqK5Kxv8LGZS1gNeLgxyt6j1aiyDXc
SeVRbfNyMdYNJn1l59SdvgnWRr6+0NnD67ALrgZy+l3+ke2TX72xA6xvJYI2rJGk
umKexkhgByI6+Q8CQPXIbl/05hgYxxIS4zqfMnppHvqsPnHKz2IXcFXA8052nku4
0ZM0+wdM5FJ2wYxCGsjHN2000oFsAIS+DSMC51yoNTMCiDdX+1HnQmR/1GNuLziP
5eDKllFULyEvWzSi2deng9pLnsUQJ7IsfrISkWyCtZudDm7N27Ghx5UaUPveyxUO
MtLWhJ/ceMGTc/jolsndpBRpsL2QtXPH/yK/6beKJNvK/Lnt5/mhYgzrnth/S8/1
iN0TlNI7LTyr4YnGn0T+HbPuSthqOu8j5pi6DushpcH6xxQLLWc7M2JKn5dH0oD8
K0y7amNCe450zUP//akWp3jSYLpPhiII4yxpviHOoQ26trE6L/wp138hmei+crXg
anpZKNPh9YeqZPw2U0L3qHoZiB9mQ2snR48oXN1QIZ48M4cSC6e2e/CFTE4DUIUv
uC0IafxX04zH6+d2VflFUYz6CMtDbkUPlI+9w1E8hLatB8JijFzex03vzt+B1Fjw
WUa7C54fWHi9nmR+K2r5JlfxJQd3qhNzro5rhcQE2onJl7fNY1nowptBn9vEISLG
zzKg9SydlZAYu2YtkXDlOuFCVQaytipMhGdDpQSQfnM4+975gZ2A/BT50Y5wRLzz
gvI1Rv5G7Z0Pk2MIe5v2sIBhZjAVXoTl6SMytrMljSo2TyPM3Kzu7QdfmTgY28bJ
DKuw6eGRa9OtDsZQqtxgW7RwyTr3UA+5ITMtbjOAEuX3ahGEXFFTVzQx4AdU73Ew
FRXOiWqoETiDk4DaJr5+HZ8xl9PatRIBXkJfFNyh0HS9rHJ4jNmy0ECm8aKDNinS
nTU1J/di0XS46ZvpYBX/JOUlJMnGTgBsnGb58j+Tl0dXBW/mN7LOuH6cN86MdFFP
7+M7S+NAi4u+uXvuyuIe5eelYfziqVdgZbAX8emVRVv1x3ueyT0VVi9YvMwY37Sa
vw9KDKLwGHVrnlq3zkkBx5zSkx5xfXfOWnq6jJ/cCPz5wB95i0Y9UoloiM8AruIo
0oM+65yr6J9StvMwCAr2iPoS92rW4k0v8rCqx9reiByU8eHI5+GAYXy2iKAOViwc
8xFdkXL1mRDsyDmcRtO+ntGGargK1Mq+mpz1FpmQfGO3WxXhVA2LMMt6mlnRA6I4
KTalY3fDMTrKQD/P7KOHQ7cvokhhbeYc3+bztqHFd30bQE8A5oT15ZYiErIstaMn
q/9TywixtsBObwrW1JrietJc0hNGh0ImsVnb6K28KPEhXLPMhnlIsoL44m5mZqnK
FVfR/BxW4JcrWgmzg2yfAu4lKmAtZTO0TD7sYfYGnBkO+RsnOl0UsIUfsfIPdwDp
2dxKNeOTn6x/8B8WEKSO9BbFx8TSuivewWilTe88CHsnZwUbP4J3a4NtDF/Ob4hE
zUkhtsXbLw+ON5s3mcqE/1jsFUjcpnfz5d8N6fASuSbEg2k0ZhUELKQ8gRJB6uZe
dA3fCj3C+yZW48oIXhVnk2t/ukU2X6b5XXpyuz5JOzATeE9+KEKipB2SjYJ8CkgD
Z1Es7pfJsbWwnzcE7shr26WqfLP0KwXEywwtXB5MQcOF2ewoHFVKQ/LV1GiPi3Y7
CEI37hwwxiWcQBlbV3X3FZ7YSBCmeWQ/wYcjZf03SLBjh0Vyz6rPNz8AnveeT0/x
/62ldt4dqvIZLw5fKkMrti2Ak1yu/Oyi38mQcf+WScPguaKLPuIvCqzBA1tki2eE
yjOWFs9U+URSMB7dcLa43gyXhJQMBmiDll6ufsADj1BIeJmmQikpyOeZbL9M+z4V
G6zh+SKnnY0FSUw1guf4VprxlD6kmYEKh2u0GUFyo2UQBruNpThNSmxv3vvP6PfI
F+k5ZruBmx2Aur0B0oUGTuHRMbtC+lCuH/NM2mT+KLuYsBR1StFSnnrXcZC9dZUY
2R6jjpnbgEKKnU8C6moqx7XIK1A9TiRBOzsH0vu6nSzQGRT4sy5cIoOETNGsQQFl
1cD2rCphhVQDaijChgnvR/5Ah7WDTuUhC9y2UWfzMInk4GCA/7N15mTp2MYirPx8
va4dpTi2nauwLYsGhLfZBPAxrrYI27vqYfLyweck0yjaTNDp43Dz4jPis5HAc6Xl
gwDnsGXnUW5WOEG1FvwBcl/gKUyl8CwBeDwG95zQnY1BUzH4y6ga93+4nQTf2vKv
zy4aykpqs/CUo0Ov8cJRR+lTNpqyij2a3k1tCqigvaRemp+F1P/RYMcUYG2mBOYd
CVKK6MGLfnsAQW4+0tcFp2SD4wlND/rlNCIfyd+slgZ47zidOXnVBdROoma/ZoS1
dAbHLk/EHyrCvlnPgX8q0oe7Q8FClYbRj1TJ+xL/xHX1TQLoG4GYNFWYSpLH6/ye
ai764LAlOKPJv7RN4U9RFECYTyP3u0FCK+UaHvmKHfz4NbByxBdd5VJvX37EQfKI
8S8qjaUOt+xrhUtksQr8zoJ4ewOmMpyFHuzub5/a6tx61MwDtS/Nz3skLc1aJjNn
kVNmDAuvdDiH+HTRLDvHmtixYzOr+eOuM/MxQLAhoSAB6KeWvTOso9RsFAuwHyrK
sy/br5Yrb+uoEuvzSnpNsUkixwdHFarCDVZq63mQ5+4sCEg+2X46bGDpZ0C8abGw
6rT2pGpSl1o1LgWFN/v/e4Pz3W95y1+hI1O4e5hvh0GltIEZ6qI8ROX8xvUpMFLl
T5/agV5nDUBuf3RoDYknGisKoiD+EGZD9Fh2sw7LZYVv6rx7N0TrA2IA6s4U22zF
LlScrh9rrDCT2DZSgbqfd9i/dE2zdojzADPLoQ14Z1BbIBS0pEboJNi9JDASVVBE
yzKflTCaTk8RE1cmrcbngHv43sleObuCmmFD9h/sjEWXqoQfJsevV70uWY8cnXM6
c3FXbxDvkXIIN2F17DK/cTmh+ZgyT5a4EmkntD5HC2YJaXAWhn4UP1oXX/J7pREr
XgQ70WmFyrDSonSj3A9TEMSrjNzl0J0L1GnGkwyvx08mwdQ6eNvqWVyctwUOaciB
PZz28AbtN/0QsGcpiXoORT/7amIKzbINwyQLYMLPrAwef0Kfxtim8IgP+QvWNjhq
NEWCF3rZxHiRg9xVWWPK5Fpy+2VrOiafrlMHAgriOqIzB9wyV8ghys2ALRbS7K0s
rCu7iHWYaC3iEyvUzZjogdGlm8KylC4JNPfgRrPdV90NqZib6mRDm/Z8eX5KXua0
QvwwqHTDRLPWVI7ATcs1b44VNp7fVBBkH7nb9skdS3SWqfmr8JQGUos57eOFFrJa
2eN/aOke+iFMwQ3+0Jl+lbYo6lGI4diVvTCVuzq/Fn+DRjCCxzSUOKHRGuLIsFop
cCxFOTxF0E4OImvYAeSavElUBBTG5uDz+QrqiNvUVyuY96sgAdgT0rQDLCwwhfU5
UL/8JufrAdtrsk4gJb+AEjs3dLrsHnDeo1URVUmke1UAWht30d257Qr+N2AGHahJ
j7rxEfU92waLka3J1SwtoqHq5s4UH2UxbANINL2vCFtngHrSOK6PRTkI5Wj79eM1
saiIh54F0KfHdqpKyaPClMX6yULe2zTDj6YE4Kp2Uk1CIUDXk687HHMLWFluKM7o
iqiNTOSXNTJ9EdO/oyYnNXdCPzgz7Pd1hlJyW9ZV0DN8ResBJPWlOkLTNwYz5iGK
S/x/I5y06KKUNMS3nhXoWZJxJ+BaT9maLOl0f4HfGtEuYyQsVfZI2w6FSMcnZG1O
R9podAfyGwFjD3IddDZd0fhJEz/gCpTd9GqRcPEKWpZaA7TddlZAqoDoaMf9jjcl
lzVPm8eu2YSeycXPF8wviiLJQOnB4wQ5Pk/8CuoRGPPO+sRMIQjWj+X2Rh6BBPgh
D5rYzRByAx0gxAvJ06SFuh7U2ZpNUX3zt53PBM01pafTZtgrTZxd7A/zpiCK3Lo9
sFvaY5sPGNqRw25NcoBsuGy/ZQTJ8JG4cz8MMx/3M8YK50DL4aqLXxoUb6JzPnn4
2CNp1iddimEYteUR+5pkx/Ry4zEelJRLg5uEa6W/lvVLzsS0mN/f1bWXgeqqjuXk
aFedVkD77/LipKD2U6A+bWv4++MrhvkidDkJM3s7tAZQa5zMFDhCELalYDYedqLm
jvQxumjlmfNwKOYGtrtReOcJE7yn5y7GWGowGvaOiKirnwu7G1VGnLriAc24Vrql
3PSbyLz1CAry5445gTBkxTpQkhHvuisZPZRrfhOOXRUFp+MaTKytWZhewfgmWdHA
+gJAONDPQUpyldDAAGcOVcGiSCKC7sRDHbL8o3JJLLGoPPWd75jJNNHyuiyZIttu
nvi7+LCazygY3cOQlp1TOQKxKoBO58KDinzAat9AUvOEBFNjCYnULMKtn/vOXQXY
17o1sxiGNC5WtLjzxK1dJ27iJllcnCuHHT7I9/hKbC12bjzwtXvZLpGzvLzeTNpO
29eTTmN/UqUc3lWKKhneG/Cj4hxbkQa/LBlcEw7XTEj7Jjl8bL5Gi11egEA+z4Ot
Mgs5xR/g7dOn/Epz0r8dhP0L8+ADyVNRi0l61piShOU/jyw8gxA0KpChLmcdGr+X
w0ba4kESA3DP/RIoXBL/Rnx0fYd7pBznruVxzzG8z6IiZQIZZdOvCXxi4oR2uL2x
LW6ofOZAtjDqwTZVaqi2g4sXkgvhCNLubF6eQ8GBa/A4vMnh1y1qc423l3XHyzEF
/EFVYq6/FI2ZEMVANicIExPxzOMUhF2lNVLvqp3QVcm79DCSSRXu39RMr+vVjKEb
dl04TrNqU6tCDYv+nhXK/boDxRMsX+nGV8AoJG8C7wbCZadKT4nNcUuMnuZgBVvO
2onf3nRMo5De0zoNj9YUdLZ6BBQfWflWGexOxnLIyKssl/yE0r/y30Xf9QUDt8Vl
IGK4SS9WlPVw6taG5mlG6/9fEaSEKtzGwNg3xwbOJozULiJC2wpt7KsYsPw370+f
wMF+shiT7MW/rmO1GP1SwahBPuDf09GHkq3vGnN7hQ1nr5Hpa/YD+9RfT/wrT8ng
XcohbEKfgnxfkxOih26J3uvhFnrqdzILpfh/VigkfR9sNU8lprB08ZLTWrBKptBA
EQaJLiYF5qyq1NbdTTS8/UOoZWCZ9Fg0R7EPMdJjxBlxKtYCA4t2dVC/4mCxaL4w
GoSKAbvFzsy4m2uqQkUfaOx65a8+fDN6TsfNoNYrAXCG16I53eIqZot8sb69dGnz
qchVW9364C0rNQnzLNMRwinmIKoR6bgsBwTbLRzeP4up9yd0WEQaDP+cOMzw2ETI
enwEoW6N+caz8lCQGye/ChWMcKkB7Ff37dbP6ybKUxNhhmNlCrE/gvUuCUf9bmyr
DwsTVA1yyqmW3ZFVzU0cBiDh7wBUmA82xaKkQc6tpYCjTrz4DN3IVV2V29ldQl4N
tdEqIBMh2fK2dFDZKVg1hj6a8EKLC2MHZGhlxEbG3ks9jXN51sHfFymbmhxfW9Zx
hPe9CnSJNs4iuEHxYQEk1snVAigUarru0S0NBsCs8UXJT71CrRyo+k8KgFmKsMbX
3lMCaa2dBIZVsh5f5UA14Y4vWieG2EFgCL4q7IZcJqduedJLERu9fHQPcv1+yD6j
8qmxcZ4t8JUBz/BbpKOqjND+mNWy7lYAOjFjLegQmXHTIJx41l/hGc25zxUBetW4
gQCRvl4xDXBbKtlG+j5M0yl7l9/lWX1ujkwY+6ShKEIZYZTn3EEilk56CVENvlbM
DTOY2m2GTsA6b/5bHX/dL+quF0H03Lgjmbluu3UO+lWyCdK0+IoTABJ/vkjxvzFY
Q6d1OE9wzR4ZzjCZc3Z3+AkBoj6PpZEdbYEMF5zDw5w1C2mCXSts2OqDEQnQKqqe
ZLHqaGBRXH4Q7iK6TlSIP3QD+40QFjDdA4n5+qGwSXhi0obWYkEv8nOeXR1trfiv
0W6mEA8BHt1fST1jsLtYDCcafkd2YMIhglLypgtkOXR9uuabOsx25dQMhEsidKrS
VnCOd2taKGwDKSHufFuiQXafYU2n6kxHoFMqWulzcJvjj9UEkNyk/FzE60YB5F0k
LrN16XlnhIrETD3ZBFhYMqLB/spQbdpamN2Kcrmt+r1PmO+ZNokPcTMNTTkmWAzw
n3A5T8otItjEzZG/LggtvT771hLpB0vvzORp9ojqdImKzRG4pH30znlNyhapKr7w
VWO4O2UZ64Fx4e/5ojXLW5Fz2yTaD0ibEk/UmJKSPifqqZw8qPsktjp9dqOVk9hw
Kjw4cSYgMgnDrayK+E7TCSYfgxJYJyMSKOH4wFHPE6phQnORd5d/RUtR3em/0x32
12b1T7RzmJ2+romqJ0+KB4cxyObaYr7SUWGWEeYjnGDVoGm+CQ11FUuyZGvv5HBZ
ofxtrgo1MnNMxcI9bSuJ0LChQuT1Da5Z/clZ17F2kwWzMVNVXDHbswgqeZfEw+HB
QPbTRsVjJOsAk+99UxTNddA+xrV1WZKgHDNCgRlI90yRtR1lyDyclnO+q64RV6FR
0YX1NVtY2tfOgn7w1zUC4/jcZN+3pblXDb0hk8YTeE8VeisxdHgZLhwG7I8Un4VS
eYV5He30iZww194J/aSCvqHiuJBLI7GOcqaRVGZvL9INWu7hVfLbKfHPag3Mrb/x
DbP7PQJQpkisqlGayAqe9AELibj1AKyRAlzwPD2B9PJg81RXuFIvl+xsQAFfFIam
qB4bQ3zgMBpmpDh6nfPxlQgA12t+RfHyeeSO91W9JY8vkk+ovp+Ws+Ol6US0pPj5
ZcW9u6TNqyCutCUgqpVP4Tfvxd9lLSmYdONA+a6KrmqRSsY/9QRoZ/ik9Xjf+289
BVWoB9Ub0rIIzQnMVZQNdUyu0x9eyEvl2mPqQWXRVUiihuCkz0UGsgQ+ptJK24Zf
smIZ/+G5ya7EXGt59xj2mdn+jfTqZWWHv74RCXl7fLL0kAPCPTXDV88Jq6l+xLLZ
SVqWr7yXeUgSR5DgoJU/1l+8BU5+fG5jPxnCaGlw3+khUQnhnHteDuVPnnHMuxT9
hnBLTnlKjgGNoRdHOm1CKvCvd0RUpSt79/A8J5WXMhV4yplEfzmbUBye82RQbb3W
BNon7gI1bXkg2xjq22z6cAGQGRxgayBk7HnpJhleJdgTcqYgS/wTtv1WbewuMUz6
/L5O1L/rkB1joEHebCo92SUq6SUaIpD8Qe7PDgLxId99RhmCrUa3l9D4FQz6w/oT
qscHwXFgr9ZMeksct7h6znJFkWzHxTDOVEOjjrXBvXClFb8f3oS7zXPcz7oVgjJT
jn94C2XiHYTqQg7kjdWD5FfPkeWyFOGOJJVsNCXK43mq/t3FTsDCkAd3CLfYL2nn
JE3pTS0utvlyrDOGB6v/JrIsZs0PKR2qetHbmweep1kpmCS8vmgoNsqd4CUL7TmS
a7Ay6DKpA7C0zrptLkAHrFQBlpFYQQ/kn2kfgIFGUD+9To7VU9o0sEnoctrFqBiX
zoV7w5SCVpXYPD5OCTs2ovdCf+cEQZ15oOdKElIAcvUxsqOmukwGZHOQ5XEspCuW
cdFfIfaRK/9KNT8hOo/LzZjOlNGbUFF9fU9O7res+52pnT48ORTdQPn73GL74+J7
NQYUY6urg49xd5OK8BgSw6tjmqdNE7WTsEymzoQmrmOjtS/2HEU5REhO2Zv+5Gk1
i+OypwK8bQyVwAKL4nHY8MhdhqRQYNlh2YluctlEmgPb1NGEWLsUNSD9j/HcqRmD
2SkBuQqcYyXaYCAlR1oGtdtvBxe/7GBSgASnXVqOUi3Jzb0hvCoFp8UYMR7bFWGP
z/dkK9hARWmNdj2uKfuAZfrhR1feXXdE3hjFqSoj4hrrEzihXZ1G/eN3Kg7Q7EhJ
sp8m1Qkpl5wpmSoN6rr6bu2JxJFl2Vh0t4bOolz0drkfxV/dyxQz330TzIw7/9aE
BiuY7TdQRNvftpNQb6Ei6RMs4cuTqL7ZO8Xs4kj4IxI7tFGk0x+7+ri5tBmWcFPh
lSm3+SyuwltWD1xzyOaiWfQ+0hrH850C3+uy7wSWdLk2YiCHAYMdT3VRNEjOvB2C
t1maLJVZQWPvDsx5A2xDQldR4NTfPxEFUlF5elA6DEzVtaKLEQgLgQh7UH3qz+p7
lRVkYCTuWEWYrTShItnFoeQ/+taBKyQ+b86EFXBte8nCzHk3cD9GBDj7v0EzaAp7
DtIies/EujrPHMtptB+rBIe7ZsMl6kW+ShW1BUHLREOliHVlRBm7lcRUixHpw7s2
jGZ/8VWOspHiQLQqfe7glrRYIAv2S5eTZHQIdZE4nD+TOH1+ERFuvw/XZi84dCmz
TqEOc/BCwwbiKuAyo9tQK2dARAWgNZBwsiE81FkNP94T+NczMbjCx35wB4zCRssr
evjHQ6P47OH7Izfn5crgzLJ+/Zd6shNqzY6NjeBSJDz1EmAQe6zVasCvaBECSMbR
8qMEgU7Tz7CquseUvDZpHib1vFX99GAWtQLonDIgDl62KMB9IK77/1o9JksErdwI
XVVKaomDPjfJVo8026J2fElq28dBf7Q+2rru1bc6ebSC6JN2HKJASMrLOBDAcBTi
iVgHd9/jfhrydrPceG54juUPsxZ8CJZJ7o8pfpx6BV43952kLLbkzTQNKUhyakpL
C6LUTsWlbdzRz81nFIZd1RySMU17T9Jd9XJES47Kr02s12bn2IVuVKLMrAUkaD73
sUMk9gXaR9bdCWRzfl9p3VjTKsujuiM9etUpADybNHJxvCoQPUuVcXNiTWrJ3izq
RsSU4fL2GtpShP11WDaRvP188DHQZ1Cl+7fpTf3/FUvrY9cvmVaOv81GYSCGcQGb
OjPRi9eACfMiwUO5YUmgR1/gX+YJsuiZvO9rPu6xPy7ApiY5SUED3jrtW3767NMD
w1iAFWFk6+PTq89njaf92UZJDFjSLy+oMsUXUTSgMbCJH1wwPMwWmXAHpjtCYrVc
d9woBaoBB8iU1kLuhSTIAIg/wYpGSuA5uONXm6Ur02KbtoJhhS5AbMmzf4H1Cu8t
yqt+8O9CBUgWW9USTMbE+UP0yVZwG1sEG3olETALbzCJYhMDnDbaKn8deA2i/2Eq
9yCL5u01/e///4snJnbg05a7A8NaIBNBXX5VllVixCKF3n7uNAP2ci35JAgJYTed
+EhWuZWRCZU6gCDSiuN+MkrcoYGDu8ZlxzYP4m8Ay+g4mmrN7OBuvvx2hMhgqL9o
hos/Ya+1MYXlzqF+9qPTcQ8kV8jUdMzvZ0zqtGM0T6WvSoNosPPm7UF0injJ/NuC
wmhFTMuozDzB7nQfOcqbPvf3DO5CfANrPklcCZ82fShNL5YHTrPV4JhkEA+5u+4L
itpdUhrsf2TMtXSz3Sq+kv8/Wd/78dBCwOSVxH4v7o/XCl1egJYtvZIUGt2tdors
bk63OEXwumR6uQ6t3w/raE62FYSb53CDtxbTvvUg1ZXjxIVOLCfaU7cVE8tT8tN2
cy9XnTXGlZ1Ny0z41s19QlI7iyWHrVXPmVBVMwgC6pSZER8LaQAuw7rHVj5GAEzA
6M1aZoDrDaNqztvEARhyPRMKRJSpz2LtVv11J63L8ZFqI5EVe+UjV82ieANRK8sn
EYIjM3e0rtmrEeE+f4m/gG4tzZ8Mp/fWGV79ezJjJMec5BqocCN8Duaa0XcQ3Cvj
qrcZ0fmoKzxyWIXMnRjk+nsjv/9lXv9j71TNn4N9bxmuoMbfApCgo4tpPDGRwbap
3HNG4P+xgMu023Ja4wIZFSaMOl4X3eAcIdC0fsBJZiTLczszXh9kfSQ/e3VdCsxg
Nkj8NjRNFQM3I3QXUuJAXu313A1Nt/Yj3uni+/v33SyZFszv7J52FKin4rhDR1h3
x0SMHadtSfPXwChSKR/TPwDVt6JUkOjJnlYVS7AWUgc0S1ifhe5ZTK+cviRaKDfw
iYAfl40Xic/vYU1MJBl5shQjSkbLZNU00nnwveaEKwtJ/R5G8TEh2SI7i4PCVnrC
vWeNHzypywcjH/zD2PLyvsBJY1eS6uLpjNA4CIL/IZwTsUCMTCRYUWRj4arAUoDo
bpt5+9t8nFyO+HBflUQy7pIGJcp2uXTBrHx77/U4IXOhrCH/lI8dIeWueqgQckY3
O4yM5YHAi0NGAXrlzYKAcdWsHlSRsB2JR5anMDi2oZs8+4cte+8S+DkCK2lMr3IL
SFQDUGtJHiYoMH59o35MzP1GLVyUXyg76dl15BFUmeVGbCJEgMB9WO65Wgzdeg0c
B3i+MLnMC2S9gzWRFbAytCdZsMLfwlxKfSI2uDDPBMxU2xTmISiqdzhNpg5Rw9UT
X22WjgGsbmhYhNC9mzQrR2CcccbZEcLvfGnhHjul9sRSz2i77xF/iiDrCq0F4qfA
oRE/lZmpSFwx9wYBZesVrKdTbiLNlW/mw7ChQZpYXAepi9lQXomXrROGkS+1dq7i
DthzbLOqRhTG88X8x2v3SxGDLr1JUWQAqnYNU/byx7iX975b7FBDqwJCv/YC+WkH
BCZApuVJZRSaytakboirPF+hcRFJo0eEfgTTi+7926hOkRRJKnfiIMhq4jF3bsZn
WRl1r2yUBeQQF+oqP9ajZIkct6Pw15H+HeYgCLi6nsfycXr9dZU2VNJR7FhMNWlU
C+Wg/5IGAlQhSgSlg0j0zhUmW9pggFv8daciUIV8+uPImMCjOuzssnybLKmxpvHz
slqpaWP6+FbRQPXMCw4BNOGCMUnylnlFQuaO0Unf9KgPkKqy7LdaB5CG4ehr+mtw
5szT/FK8fCNHU6rb1OJHdXSw99UNkuUvcZ89cHNz1ApPOXYAqvqZN1JRUUBOUB3x
C3bfb0AZoytzV1Ea9qbEA7kuqmFnsLymlMvlK9gGvOTqg4RyH4j5FBdC3R70NdTp
HrV2HK3PA0AZf9TrGfItUpHiayRTICrW2SLKSRI97/6SEMhDnjO1flNBeURJgh46
YOgUiDYs9pZkDsaUL7Ji7TdqjpXNgG9SqinjuBCFNDvR87/DJVe9rwhXWRp5u8HR
mTJMLxahYz+3wwh/WS/a7FT3ihC1WV0o02tpGKWoRhlP1081vOq2Ysj+NKIZPQLT
yxnbg6zjYlR+c0beu0yCO//GXeiCAOiS10yCd+wu1lVywZihICClzXaZZpQU/R+i
ZIOzaDZEB97IbWsGPV3nfkWkqUdbqpU8gJBXMyITAX8fvQiITQ16NdjQ/5R5D7d0
rF2k8pSfXc3EG7JOVqStIum2S1TJUaP2jJ6Cgl6zQnAsdloAyCVozGBlbL5tkNdF
2dvHTs/U0BYG/2UIjbd8vjaqsAoWb7Tqb5soDsn/h6ii4lNim3h5Bo9VU8ozyXhb
YdmVLLS+XdfG7uIubKOuv4WiJgA0lPbGN2WMxwsmov1WBagkY5B2ZP+aqH+c5ZEl
7DoESgNgdF6CCKRtpYDKjKQCTke8NNDdEMe+glTt8tBh+y7q+Lvqzz4XY820AULg
lRTtP6St0nIvUOq6DphM3FOQL6e2lL556jU27tWidxqEZ/ge4yfrzI5IQMJQjm0J
YB9hMhUoFTD1YNBAD/nHEBZl+YCR3f9xpS/YRQUEuuQQcCYiTlbFuiy29bX1jpV8
IsfAwueRmHrcZn5DQt5ITKK9eyvIiI3GTr3HINPgqxPYTIlFT0BUR27m7IMKf+gT
RtJLCEINt/Ubkje4/TORiF0xXJjWnXg5QVmfACTFLo/2lzaK7ap9pz7s3NhIrlHb
zZKkm/ucX9sYI+tTyFbQKRkXsLTpERnjqDZ3s3ziVTPxnahDWPMz4GKvo3mwsyUx
uLwzwSMb3tHi0qXJrqkjtKF5uGJqOHxEMfkouLiEwiTU2cTCzlPdgIEKApGKzBJ+
B7aC5ZCDWXQiT0fvKAPGZAx69/IpHo3tW2IUGgB3ZrCpUSGHyfSerPeUlnnuyJvO
nAihjBvgUTh/1ijyiF6hRZz43HvG+/sNeV3m2/B5G2y1zEzw5LYufN5vXaJq0Gvf
0hSpdE84NpyAZCQq534Gwa1NCfkevWyZsOKCSNuX58AIT5/ylKiPNy2JTFChyBCF
DtIqOuFL7JZA1iowGG3I2Bxm3t5uJZOIyvdEd29qNVkHoVaOeRE08WbT32dgTXxR
C+tO62YsQtbyeWsvikjKyQ/RWGva5pbgJZ5D0G8hQRst50tP66xwLhB77eEpW07z
7srMQz8/sB/i1XtQo/iIVqgDHooEL247ep/qEwp/Ev9qzWlzm0JiVelHp98TAtm4
lQYUcSNLIdOlMwvMS4PHA7PkKMJSbd2cQ62YeCl4dTeAccaU/wrxMkqXgR2bxAlg
fe0VcRZ1yKjY83qQpas4dS3BReOGKbxnyDK7tUhlFX5ejY+ogZMdRsy6Qklda0/E
xFgupSsLC3rzpm73R3zDuiiR0igZzJgZcJO5OP0el8DtVkOoMcngHudRE8McofhE
LNh8W7afqIJb8vZzY0YN/KD5KqHuUoypCZI1RpP4s7q5lB1dF6h9rCC0K9n8R3eN
C8yIR0mFJ8UfJxNy8uPKEqMBFM1lcKmQphW6SVKcYVW8FFWmq5LdEB/cQIzfHIm4
PoQQwMgMSaHABYuT5ngK/GzPVYooi9vpZVBgZ0jWrLBS+DYpkXeHoQVM0LB5Mhyr
E+NxDknOtblHYBtS7I73PEMPS9/4pzImOYwd4QUIGcp9WldePISipmeJBhexDBH6
85tdCKqK8+IThHb4bJIC9aka9EMxYxNTYcQtCGWSdKHOdARQ62MTg1jYGexZC7pK
czD+EroWP0+NYZNQrwpqR9mM7sjyotPuit7RTewpPFPoLqSXh7RhMLzaJMa2lJkR
LEPdsstzQg3vPFO7dCvelFFIP5Oz5G8LfP0/UBnajpiXUzdTst0JJqJtIxeTD38C
kY2T4/5fjzvUPiL3b+oqYy30SPkXqVI8GW6JIbGTfq5WDFXf7Gv0wuhjzSB1KWob
IK2rvdJDunSUQxPtH6q+3pHj9WIL7J8pYENznfYo91wA06P5+figdHYxSFlHvASX
+LPZh1qj2ma61+kuv/zJGDO4tvSsN7yV4S6VPKmEvH71xjaUsnxfL6mcgE5iu40x
4ixpo0TVXknasygdjfHMZHgrZjZcoZ5w6aO5octkf3t2a9pfdhER2kxFhRuc7QLN
2g+wY2/lS/q7yaSWssMPIicoLrIQyMcqzwbe7l344ePz9tBexYra0oubdfQVYw27
url18P943ct+spJyIEXGPETBOGlNYcdcC3SBBf4W8P7C7urJkfWN2Yc4vqN7Z+js
UzaWsdCjzdxgwklk7rH3WYUM6rG5ZjmToe4FortdjKBbt2ws/ON8nEokR09G1lxj
8og4ZsHqXezv5PvcGRC+LIlq06420ckOq+wQz+E+MpiS39bfPRUW6QejIOTv4pke
LQ8EcHnhOAYHnkGx9hHq3Hj9a/rItEJKYHOMPUrIRzgram+wA37YgpfmbUEAwW4I
iVa4QiXHilJxtGCpA6VqVokq8UWsnBkq9gwRWGmo1DNgDq+7Zb/M/uwocD+MuM3N
O8iwGPr7Nd1WQ+DqSGttcD0U2XiUxY0XTgmXKgO0KZ2mFpcZhiy/aZw3ReY84vVV
xsis/rvPN+W5GUFxUoKclNXvkM6VgsRGxSwfDAjrKD4qr/VsdX8ZIN8Guvw3y43Z
3F+sSDO9pPIbRJdbE+l4C4HPEGjNugroYrpXHKRajpoH0fDFsZI72xHbTnoRz0+I
kNfk1dwhdzcxVcyajEBiDbhNBq48IfS9dL32bRYxsViOukTcAcHkp3g0ba57P691
DNwkfhiSzfxqoFvhujZzuwEbAYTze5UebmXHbkGjW1BUTS/MZMuhHRf6vogKLsRA
0FulJZx0iHxOOFuqNnb3Fq0G1C0cRUzFXRTnN8ymO5ugrurQnVGZbHbTUi9kywf2
mArN8+8gbQviTcaObJlZnT4sx6QOlbR8qSvsdFB1VP/OHNtCRuci6037xR0GtajM
mO0gfulzsh8MZZmzUpjiLDhhX2RXylZm9kNwodnWGmCM7s5Y2BDWcYRsDJwdFo8t
mMR2+Dp/6uGzqpwWttpJUVqUMjNExzvRqkVQo0nQUIO5oO/2py9CtwLRophvp1px
d2yI4BllJb5EJq0Yak0EaE9LYhzLLeybL3u1k0HWs25uz8mYIrsFfzpwVQflvG8P
2JxuaJ5e4C+u61lb8OkpAm3sJv7N1Dv4+LQhVzWLDGyLZnCx4Ff1zLy0AqW9Guyl
vW072gjjYrY/Yn0KAFqmkZmssRW+JvwEk1NLMOBantRdCI7xF1/30s6DF529n8Lr
E3NDpHgZbCKO1Dr5tkDsw0i7oczG009owTnlLu0/JeDKrhxncL5JBo7sA0ysy6c1
cObvMsLF9wwWEWPY50CMi298X0LjGVkvSGhMcSctH0D8vUIVVwyKmGMaGsLk9uyB
juQVid01Ys89rKiC6Y8iI5nk1M1ANgMqmcfGq8rnmBzNvHhYGzeznEjUTG7vvkjG
YKkmNOstS0usmYfeAJl2eeg8MDiVhIt/9ZToNcMH2aQvRuVrkUIZb8lHfAEarW2m
DMCUWM9/Z+PUCSNI6J1+DSL2E7p6gN1VbhT5P8Ytggm7I/GZnQJGPNB1ZYFgRKPW
SCnVixWUexKF4oWTxlA+o/JcVINWGupFFWsB4VCE2JmFD8xZgqI3P4lQbPjgRFrZ
/NnAAYkT3amYuN9mwBONqf/iAj1kgtfUzSc4nSN90eDpfJXFqw33XH+jqX/GcdF6
PsiYKr/LhOfMnMWEHZGuSTDNDbFb2c6gnyeKQe+gc5Rz0saNV2IjlouZ0f48sJv5
NcKCqEcsagJP7VKQnxUyNTBcLZ8eZN1E7LqMe/3FSx6fkL0p9xHASlIdGprblwxa
8gJdwcbE9NCgOeEjTQijJfOqAcqQWwWZKn+IEIhPZrRJuHeib4QVqip6IaDfyWY/
Adbepm45hVXt+/LDVbb64avx3L4mwhz1b1K/jzZRUs1898oB1fwxSYuDoAmvtl0j
rxZkzm+4ncZEN+3p7bYwrRsEkFbAoqYECvHgoTAJuncX9NifO9+9u9D0SCr0tIO7
A3u0/4/UNFWXe59YOPES31HtsOv3REFBioiZkNVQNWDbsGYBPCXFEHmYUdAAeIY9
V8nkj5IlYNnT/ryKI4Agz+B0nIhwBLf76bHBFteEPnrYNZ/8MK2vsje/qJxlZ9Uj
SIm6a67OGG9siXz3R7y3UVF8qwALOycFmAL7o8l5OEq2hu5A/psVleENlARMWDc6
EN5VHDSAJRdLKBQHCOxOy+JSXrNj7k8G0mUy/Gzi0xY1ekMUvn+RizH5up1i514i
bX6lj1OGvemL0fPut/zXvTr/i+znlVi01GF8qSOiStOvquXIxvjPjH7pt49bdWWB
LmX73M5O2QxWsq9xSnuzmP18CPWUJkAO3RlYxTvG355IY/pzl9YgaZA1DCLu6Agg
pgGOMouQuABf+PtWxbPOQIXWH7Lq6FgGNAPHpaKVAIgfZeCqhssTJfFlnrMqz/p6
XPxQfCT+y2jkpF+McP92db18Ct38EodZN2FsfQVqRW7IRkC1AF26KhrGaad3zzJu
AhjKOmF/zqda3Txh4ZUTmMDrIGdtC+8ghI8wHSKhm7NjsF5Lrm4K2yrXEL9W932i
FfwufIuLHH5mIAEu7MD0BfERXoetB6QME8mY7GbDq0Kt+xQImABGwAlXJj3N3kl1
2XJOxFjojas4TZg3MqOMF+YzFc4DAX1bFOHJE77Z4aNB3dnfKEeo1CDHRlVntiMt
mGKiV8ZRMakiFGSul9K0kXD+DXOYQbOMmg3qey87iYxr2yjtWDHHxthL2+slRvqg
8rEwGSqBMo2nBXK7+X4/wUjhhhsrdzKFsuUsGB8N55gu2NVInwvJg2jP7GAjb2ou
ovuZQxwbfs85uV7nBAnTTGG6WS1r2lm98cMrpTo6MISNe5IDMcNnOp5jFGauC2us
UjqWO0GbAKYzW2/X8iKgfC6RCollNj5UBVfJG6bcp57Jdp4Ce4eykIugi1JaD1jm
EX8T5oV+grc1yRgVnORPFfmWHddqMzDy8kmCibB3kCFzRGlKiIqErmGWeA/lr7Nq
3K54qxV9R9IScP9FXBmM+AArPiNnNGT+IQwMkf6U+hyNE0HXv55Xoi0AjJtgYZVc
67g39bV8R8EowB9S4PBH6UYGlGGA8GYHp70MFFm3bg2gXkAKkK4t/Q6DDga/NDnK
uCGqV/Q5AStaR45HKcY0qUNzdm7ucXtEu86Ybs0hJPcV+z/LcZscylyAqrQ9WDEr
E9H/4hvTefaYpM4gYS5dNtU1+8kdxlobmnoQUW+D+gl0+dbtt2HWSMNC0plj8hMz
pdQA1iKZjZuC+pyGfvJjkdtF/2KXhk1hucQA3QzUXmViOpoQDG7+UrDxTv0A4SJk
eAEXcoC2Iy66CQuH0KfeUlcWM+Q7Tz8earvGnn6p8EtNX2vtWkmbSMwXlHirmMc2
jwk9wO2PDlIcXGmAeP5cpPp+XaVOxfM6+R7umWqy3jRv54dG1dMYvIU7juPPaxr5
e1BBSaLTu4dKMgm6Yf6jOLG4KUO30UDPoNpWpSfWtp2miw5uR9zyxC+MKGGgizM0
UxpVQnQaNlTFVNNH+YZsxb6Kb6Meu3ay8WwXjWl84EJX7HCstU+SlzdTkgy8uikC
uLO+qho/WCBL9+AYzqOcmwrYFnecuvEoxHHzdw8AbpHBWIGmy7VDlQQLyQgNjXvd
wBW3B/3ZpsKcNX4unsFfTExYg2gSVSl51SQZukaXVC5bI8D7pPBkFp2fB74xLhoZ
aL3/yYxsxCmQvNFfi+WEPyDM/ora18+CBktGperj4rNXi/r4EV4EUkUKZSLTvaS1
vxVvEYhob5GvCfBAy8pYWucqmR+umc9erhJIpleSj8YEtzwBwHb9s/Q5MesbG7YA
yFr29LjDVhVKKqlzzIlQK3qSXohar6mFLnQ+b10q9r1Ndy9gkllFbLHmpQmlsjHE
ZGdP+cmVSrd7Atq2r1raTdxnqo8M6XDMKUx+k4SZYvV+Lg2sWj7nmPZuWuIhmRJB
orD32N2zMS6qRzIZ52jPGl7FOSEMwPtb7EjwBmORD/gpY+/7f4vtB/qKeEASd4in
hvey+/nli/EpeLBoHJ+9Kb1EOfxmHU/5+AltTFz0KSAUTBOEAa1equ78quvc3dlA
EhQEGRsYtw/e1HK8fefYuSRoH6QtKRl/ebffKxFGadQykX4Q87JZ9bZ8e/Oh1gym
7NYR/uhSvhrf+7Axk/qrZ/1VdYmXXyk4xRUmZIealAlZqugjhOSITBJaBN3A9AKB
DK6zCX6/lmuKdFsPKMEWoiKVk1wTYqinb+9KpiCegd45yJqSJ9hc+ekAIRQWR/hz
x9nS10x5pPQJaBX8p1ZaDyR5QaKmGHedsuV2/YrfNdABikow8vSCHAi0oitAcy7O
TTZ1qfr58jYpm0mfvae5K27jfWJ2TTzUI9TxjUgbvkCmJJAabiCYclSS0a4S/vRm
OWfq/s/rq9tHMq7TmjNuMA6e5i2tEb8soJZhF/VjNwCydGDWjdU0wq/WmKSB2/oL
CCBxSbp8Vdvy1AOpLeMaBFcXL1cZt51a+7S/rJkwSCbxSQktVIUKNBPhKssGm4cF
qUguK7ShT7jihmrQbgfDrN4K3/Nwm6k2PCY24wa13uZ6o0gBGtF8LXykE9/HU/tV
HfVHSqE85NH0y7QVph88RkFDMQQTxWVQxmgh9j0vTDngVxLxTQ7zpDE21rJygDPx
LmbCyYGGAG7aUnLYlDK4Z9NSIPG/fTnwIfwZOfagBQJ6R1qsmQFY8gCpdpYWtIal
c5fcQ31vZV5pbj3mb2QThRUGVhDMGAS46WC/HTATByV/io6THqm3+yo5qYiDZYcD
K3RYtrnDnaVASPDbEhTYA3Wc1n6C9lOuOvi4XUBhM776rQsjlxil0+vHAIO4Lj0M
037pqDAJjWsKTWDq82tYiIBwljw/HKqHq0eP/VD+s2szwJSqU1jKYMaMs5EJODUK
n3QiZDi1GX1NdVPeTZFKwouHtqDoTuJqtDKK6UUjQqmAKq+hce9yiF+GFPI01/HY
ETVcMUiwEWArKy0CSSgPlP+NyKEaeMhUYZYWhjq8/1Iw8AxQHgYYPY+j3Y9LWmus
4kkHjfRq/izOT2wL59eS4MwWwlBp+D3QwNeh/eBSyl8ABiBklLUKsLQJhReySHvN
Yu+ZrahkkwbnDyXmepchRm/be9VuXj8ojNc+5t0qcL+1dE2b1hm2EeiZBH+D7NTs
hceiCZaM/PDRz8V3xNFvRsLzwiEGm0uAqQ16rh5vspZKKYvE91L6KFKXwkaBP6xp
eaXYEjn9Bev/PRag1tXh8zwnGxelQv04mkLcE9n8QdpsigWhh1+mpIKNG43lc+Ep
Kqgn1khHcNgKPqCLZ1ZSQknNwK7FIQhWhVmePBxSYBHOumLHajBRHiyqn3AIndo/
066FOUhh6b5Y7yKjFtOeZC/+RShZHgQ34NN1RDaLv8PwTO07G/p282kXpcDcNvh2
uFanC7BEtiq95z9oi8g2DDuFkd/WiNGgI2YmOwhE5qUJUD/qfy0ytZJfVmwBA/ij
nd5b7L1+whDmkf9p9OSVoEc8Gm04RuXZ4PPqji85B14OJ/erY2VTVFLWa/g6tiCv
kKhgpI1BK4LQXEo8iVfTdUztRecZD08y7TAFA1YYTZUd6PUKGD0Or+b/+s8L11qN
aPHLK9pYe2F75mIUHr3ewJ4amKelSW/Mwdo0xT4/ulfXWME5jRM+QCWuFigwgwnf
u3LraC1H4V/WtYmS6/mW7srcQrnKSxWdm2Q3U+JL6pZbzn+SkaNoJmbBxDLB94N3
nUkM5/5Ui0vWAaH8F4A6WN9iBBObCIri++dt240iIzHsxWAY1X1UR/TMHWNRpdfC
t50v6U6BncaVWl/QYHt2iEXALW/Gnq1NQVzbpWOMW02S2hH47eD4RVC4DXuSlwdh
iQAd9ZvwPM1RMaMEnPhevhaLaCQ1NkaM2R/2dgI7cF+8+oXNhku4fxEfB1PD5hNe
+JhQeE2ht8dZse6CIJz8h6QHz7Gpzkfi8J8MWgHq1zUTZZmc4B6zqMAJrhTpmE+3
s6v6EidKox5vZhK2HadHLXdndzvPNXW2jRz8JfLKLVv2VKCJrPX6fGdxFt8Mm2hI
a1SxuCruOwm7ndGz6zYl9HQPhLS6xkVbadJyJoaGHqylEaZRnY0IiOvpLmiwlwIz
hvjGH2nRWtR9lXdEkFf0mCT5St2L7wsn7kUZUo0WJeXUBEDRwdj+EiFLYpmAAFEW
YgTs53dZu8MS6QNBVQ4SxCR39X+GGCjE6RwwdPxz/leTmE1+rXmQJq0cPQz7JC5C
AZQKOfnRPOrJmrudgtL/MwFFPySikhX3ASEGAkwESdN+SpdSEB/ZaT4diHl3DpqK
SBeiYZtclo3m8/0dGDqr7rP1v2+dr/yoBLxCN92vIGaEqMbvnKgG0RsvxER0lENl
fjV/kRpwZ5Kk7HykT06okGZxwDcAe9ayxx89iCenW7iiQ/YB9rmBqSTm+3+xjOHY
i4eBFIylRd/thlDcR3UKFX7yosTfi0twmc1tYSU/o2qCMsZcZZQ8vezvdNfB6/mS
45bTj6BT0BrHBH3ziy5L5yO2zkiKR30Zp6DVjMQ5CujcWFnnq3eSTg+m3wzND06s
kmaSu+L8jJ6/F5U1iumJuaeWAnZxjujS9oIGtfugNu08ggWkz8alQpdl5U/FpGjg
PwLBdGTZyarj0zcKOU98F7klZuOEkW/F/0RGaAkX36YAu0FN7acfHuLRRrO20pIg
Z625RlxJYnfrPV6yQRCG0eaYS6aLETo61PJ6mC+JueWBIIvhKctbl9BolWRO3XhB
xshBchHd7tLx9SWgNkVNritESOJJCT3pDAq0FfjNcdIxciMtsy82wXg+McprcXSy
aVjnt/kPO2imkGTAqSP0aGM3U2y/jOhKaTgeUvjHJgD+eIb+vOUpQJvd4PpMwr41
Bmj+ShC2kHNx0G9b6Wdzadn1SG/+W8HWTjlp3ITh0SRjHUq5UbNkOw+VfmEuAz8d
QuZNyf24NyOhsbHkasFEg7BxhIgGSwdfdCADqull/6OtA1VAtXBsWxcJQZtS2xZD
JQ3IjdC9Y49Q1kuo0nDHQPWy2ZEUp8jqdF6XYP4BrztpRJ2eXRTP1lxIm/8yP0Jr
YMmefYyxqztnsptR/5U74Rv2AywLzJhPdFPw9eTtq9A0hQbRqBNrNarIK5t7U+8Y
48rzWxm/XUyyAM2WnEf/ePnlzNKMz3dIGzkRpglj3+1bZDE/5tLOARZ1F8Rdv3ft
MoLnRmfn7fRXR4HyhM/4hDx3tUfN8ZKqH3Wfl1WrmmwUFcy6JuWLRi1yGKwMc8ll
nTIZ21pG5jGsa13pFm2OfHusfC7RNtOUTV07zP6FIoUymLNSDdJCoI8kzOtlsauM
o/UG7cj2m+QLrExwJLbT5ViGLy+MQ8PAAZrpu8iJzVSNZO7aNP8qJfh1ikPLCAqG
flkL3z6PFlMKhN6+K8O01WB5ykTu7jSLb34uhDORSBcZ46KtuLZe6cu4EZjEW6Y2
3QHaX4LKi/kWkcBDQUqbOtRsOIBVCKfm/fy4RKEiV8qEf7tn03PpU3cWk1eAmeKH
eTv3o0yBLNzIt/HF2Rw1znWPamFYWyz2eMIh1vqW1jZaB4U1Vp4L34N/yQpfd7h5
qjKCIf6k4Qbmhh94PRgBaihZN21ViBzeWAznjAUU4h8OQ52Hf2g12fax2LVj6ghm
+peu9QYgoxP86tcDJ0w4mzu+IpLhZ7FHyHkecMR7wnYxjFFKQ7Rxf7Wa4mt5MfiP
Rl/0nGRshH7sqJ2/O2GPuaBSL1riYlb1da3jedoCpJ5ScZdx+9QI/ZXmrY8yFFpT
ntL/t0zYzd5npQrSIToiD82+0yFLYYgNhHHMEWFevgiQGs2MniG41eL+fhYvxm0v
/axaKfHsleUHKu5IQhEB0g/Hq0sBtTPAfq8JaDTQXJb0YfWyZMdflvHt8/jVhgX1
QepVnYAD9wgTb2bq2IuQkcMPXagQ+LiH7Dk0JvBmcElu6WYYWH1/3iaBVhJcWyN/
tvR6e3aWEkNkvhiWg/zVmLrZ1oao/YbSgirj6sKMMFgM1pxGre5nQBmhv9BFydLM
+Xl8TlLj93G+smdUcj4tq+Yb42j+a2UaaIOHDiRzdFlUBUAZPk08wjrUpyFYu582
W7gaCJHTjvHbUDRMszkyo/CInvZ/W6whV8ZB3fLKSykuRnYCDvVVRRkTpT2tqN3z
3p/lGDIhoMZ4XK4rGKPS4oYp2IbWQ7oBhg8xpyMyd+3EDMbb8jqCDD3oeOHBxRb2
CMDk2ZtW1OwkqOo87wc4IvG6NrfNdcLuMUIJs1/qZ7imgBBKnZEoVINOxjQYAjIg
1V+ucOkrvLpyGeJ2xe7c+VBAIPLN46otLk6wGpYguu4IB/gArDjiZKKGR3q47Yem
tESWlvpLCpPjTHuIPnmq4+ydIZr7qlnB3LLnG5sFoTuv+OSvA80z9966ePMxWepy
/p2/TWhyJBd/hZWtv3PkZuNu7lR368VV1hoJTPj3irdd7hrztWt4d2ztCO2sZWP9
pgrRf0KdkpzCRQWxtCGEguGHowjZwTlXV4axUqAiVLNawQmRr/OsbdEI8d1Ubnm4
V76QVF9unV5G1y/91t8k2eZHHGInQ2mizz7JzRNLpmQFVi8JmB+8vbmIii1cwvxw
+1KOKGzi1539fWi3JIN1X9/x3HI+oaNVjhmWLZtTvZU7poPulDl47HHXOTGjQ3Od
e/UFPO95X8ItjqXheXUfavR/dOxCNxQaOZtuhLmqxIcNOShkA7gvYYkw3zZK5iNv
vtsBOkZSDHBFBGVZ6esnkQnMRbel8pI9v831S8MEAk0Vx1waHwZ+3qnEoq45/ES6
Ln8b1DYcrW+hU50XUfrwBs/3bn63VtGEIqq7H8GtnyNBfMjbZcmTHxFAqNgVggNr
f0XVcJGe1KuDLYt77vzUI18S3kRdeR0pG3kX44oxHw26RTrg+My2X3CF1ma5Ix37
2JiUBbgSeXLlRtF+B5s5XmcUcozpnFBX/i5EG+4lAKJJBeATDir/5Lp2qQ+QoRjh
x8Sw/+3fbt5cGq5seyCYCvN/wPBl0UIGraSZ4xTh+FBTqO0Pw/aiXvPR7EPJx6N1
yyKjpk/KG+FcwN8CEhwLN+56DZm2U6jEawlJEOOkQqnMTmEBkO+zOiq35Bx36iAC
fzl5Z3R3z46nH872zVLaJJrQxmn7+hvNd2dmqgbHP6UsXZpxRA5gjG3inGeqWk/k
6H1BYt//Tk1LczSMPQ2dLZFlGhWZoKuUpg3D7oita99UlYLgqfUzh2skFjon0Bz6
g1nytR1PEaphR5mtop7YNuT7BgM6E2wvjHJtgPBVIj3cf+Iy3nWSUpxn5OFPo9Or
UNH4K63YKpLbX79kYyWF7mut+yMaMy2phvgW1frdC5b/UVKOIU+PSMWdnF11ddeK
omNxPgLJhgTexT0bfr1XSATSklwV3WdHj4xC+ExJm5LJwBXdL2wcXRepdSg4/vmD
gEdpl/J4LkTwbilmmlvcBnPUVfsqbi7VG4Tn0OAq9vmcsbUfMMQcUilbbVe57X/S
OyQqnck5I1c0z1NFq5WyjAuvLql4kI4IKT+lxoCnzHt6w7v0pRr9d+CWcKHpIqN1
YsI6WnG5D9H3H013TO5y7nz9UNK6xKhxxbC4EaDXRIOQpH5qbls2o9CiYbv2MCM+
cgSCbZnf2wP/ifl/t18aF7tlCYBoJCU9U8SYwNp+QFSDq2TOe9JFG8K/7w3xYukt
mpat7P/SItwtMxPCh6PXplJJy7vLiJzkuCVa0TKIYgis5rkAKvZUIhsn0rqswJ7C
5M5qyWfC2HxgE5rQVhGte6Yq2wrk2l477SjZpU/nyOJt/NwN0kZHenQR3+KtUcaI
nCmDygPjpY/gJ9CXpz+WoEtAfuKEZQEwEkDnOnEVhD++wVC+fhQaejn+g/838lr/
4bklGxZz3p2FbR417ZYm7rOJASDlSJeEYwJsSafEFN9ZBPx/MrZRMRQXhUREvBn8
LIidq5qYlqdtARiv1o4bN21ew4AMxJxd46gKJ0DC57DwhEL1xrlQPs7XN42zj96T
YhDgB7vkJzQ9ABx35hyLmFDAMGyyfGg+n455pMeuYFTcbxsS062XLyS+XP2xu0WO
gWrYHvqWnXz4gI33P98jBUN1tpZ/Bws0OpNRfOAwMfWgjYrUB88tzqX4M5Aiw9ze
22bopQMmzB8kLOTNbtJDcqrtDHEUgnK1D6qrcyf8fsDHv/m4lii6AyirHU+pXiuI
WyHUmx+60tNuXmt34iHwPrw65TE7wtImLMoei1f7ArXxpzBnO1QR5hlPrb00Bk+G
kurp3iz5tPfkE08b3BuuwQOfvDQSxn2U9W8a03xR5MNrqXhutm5h72WCT24zoQm3
VwuV/jZM6Y0JbKgxqjg7YBMNAhVuEekCYpnCaJBxKMT5krD68Qwtwwc3zNiYzFLn
9DEpLChcMRRiOygZWZeCTcGiWLxygRxaqBA+CI90GK9Kg8yCv7FBX/YQ3Wg4UHqV
j2zL3WsKLHitkGldnM6inwSUznE7jjjX1zvAeOKgCZ4s7rw8VeZmvpHVwJgfc3JV
RN5echGrv/lvI7UeXYyrQqcby23t9atGPJ4mKqxJuCqlo2KUQpqbtv46oE4d6RzI
/ko1trTCR7vkqi52O6v6LVd6FNKcVYyeM7hNxurvOfCqsOEw4w7YhZw+kMMCnL4m
3xpwjR4diEmsaAgLanRM+4wqySBsMXRYwuMkM+J35gszPAojtktxWeJlbUtg/GKs
vW/DJ1D86ZO5kyLVipWBQlSNYgv26FkOKoREcg3plnGGH+GZYF9I9nAkW1b+iODd
EDGK7nEmZOiCdknjYYlcPSyKHcY15hrB5HpPGu+YoRQYnHmYT//DkVgc+r2qv8m/
NPEixSP7NY4QB26RVXdV+3BQdWJcg8nBo+BH5qu/3awt4KEXykcFmyHQyHL/8EgB
oEcdD1YqfsfLap3lqaYO6wbnVDtzaR62igrolMGX3+3Ljl51k5CMlYWUoSHA/UtI
3LJt9BeObsFDV8YTAUglBVRha+t8hyIIIkiG0yfJ8EdtzrpHp62v+FVTK8l2gDFa
M84JwUS9ImY1FnEYTyzwXjsCvE7HsAo972oCCbaAFlVUNykDkCe87WTJggnvak6Y
r/CYXfiZ18bqMHUz5eauVDVPfn8lfPaNKdvYBXt7WAuAIrdu5OHRSpjZdWHa+0VZ
G+wedWaaOYRP6oAhlmwaAXdpavKpNvB6Iz0Q1Zq0LCorYV5S0EXXUtyfwVMNIw31
4DGeN1krR2NYyHCBBf1tGepD+CPTM344VOz8nLsE2RDLiX0SXH4ztZKCWThhe7yf
1YNNm0X4GUPSOUoSWkLnIrp3MLr5SqKfMpA8J4k1wxCSZPTMgcp8orafnJlzpvW4
e4ey3CvXpMQwCNoIzoLQNN97r3AZyYgJgHV8+EFDEAuPw1xrZUlFQZPf1xnzeDje
gECQDZuCjqrOesKetwB6HAFn4ETjKMMaa3T7dP6M/K/nGio8PY5I4VVtmkhj5yG4
jn02iLNTqQ3gk7I1tVa9NlDANgmyZzElWRfKl0QPS5JjiW7BalVOt6sLNLSQTfT5
Ne/ywGCFxIRKU2dx1tqsTLWeRSM9qv4B/voQXl/IIDFYyaiguxaOImm1w6QjIrUn
GImNetsrNLFGNtGMe7tL6DxAy6SPDLYSXjoXml+o+nxHR/iOQmJQH0Wv7AAPGF3z
RIozE2Ft3rUsBuEOTNgWNJ7s4mz/d/dIf2M1cHMbp9rv9p+ZQ9xnoapCs3rpZlBH
rJdLFuUCiRSu4mhnF1Qc1t3gux02Tbr8vZ9FAUPNw3tlyuAULdA90Mo4iHNlc9cs
UTn9IPlHla4RhWH2+hqgq/KdaX1o8M56rWKYq1p049yWYBg3EJUUbc/EUM3e+p+n
k/KngXT1l10tADtShcNQKjifpFwKG3vE3kPcjZBPrg1aLHByh0oQiibowH6enyOm
YL/i4xY5MJlKgQ5kXPiwyi3HV2LNl//mWOzs1Urh6+rDCH6H7K+hqZNcr/6H4qFK
vx3WEf9FHdTLaTd/7bjBMLdy5J8l4hm7PdO9zcZlEWDBwlaWcGahs+/7vzQp/Ogq
qYIwieBKkoPrIb+F4paAgnXasZydpB6edjIQGmBOVn5ywb5nGLp6VOJIIYNoydYi
/pmxXHpB/xzY1sHDgRiwsH8A1o789pZqj0nejdig4v+LmTn3dVvNMXNNtiOa8Brd
AF1OkV85ZRFTaeYb/GZBNx1YXGdLwg+UWpHDOXwqSKvGBKKdmJ3sYUsH5dzig9LU
LlhTzCeO6yZLCw8Lk6zSOikC1G9vzAe1mNxkmewRvor2HNfkxKPj8tXVAkGaCyGv
Xjm97/Rn7vq3xBHdIAOpMeGP5CFAWYHQa6ndeljvTps9yWqWFZbJGZtgfSWMyr6h
7M3jHSjzE+8TF/IOBouPPd8EHFTdBsuqObsUdk3ryQ+HfJ3L490yPdIznmFsdlxk
vUdr4I12ydS9lLBWk2dP/EwHUl7RB98kXTa9QwptWhZQjT8YZJhohxm6XyxOKQqz
q3lc8Ejj+NUtEL3sujKVowXn5rCTsYf3bmJSYnl4ZT8mJTGuEFAZf/s9TJH3LCuR
F/NCKciwIBdW32BpqGYANzqSzZzRKsVltTTbSaIdlc4neyKonDudM28e5wUEqwX5
2X4vdoEkJvltMQssSAxCfw==
`pragma protect end_protected
