alt_cv_lpm_shiftreg_inst : alt_cv_lpm_shiftreg PORT MAP (
		clock	 => clock_sig,
		shiftin	 => shiftin_sig,
		shiftout	 => shiftout_sig
	);
