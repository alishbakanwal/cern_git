// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:34 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
D+JVliQ9tIWfeLCO0hkKmzFwBs+PDviXhy/sxSMKbvR/jFi2YLKkZPM4M2LFAx/H
Ygsj/Ajn1j4wR5R+6fyO+IjiA3rkwDDS1qEhHkxUZGIK5BIxPFzxOOSBsP1GWeq8
18sUq5eGUoLsUSPpkipdvXdREGnj6ja3yONVw/YTFmA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 32032)
JFcNkxTx6a2ryc9SZjPH4JaSYwnmIzgI0tTkODEigABm+2FJzdvymH5IsRXRAJ/f
jURHaCSRC1baZJUOaaTtRQySSts3ln9QXxd0NqydJ0Mhwkp7JS0Twf9dstJB5AcE
VSRObwEsGRTnFfKtVliGITwBl9rkXoYI6+PaH9eANK8Ti29kInT1cl6lo8VPn2b3
yHYKSPGvnfKERMYszcHBb+YGDrIMnWuwLUVB+9lMSWQ9Tfjdi1tsazQAYyiJHbgs
rJVYpti+zLz4hDHYKZPxf8EbQJ0I8J1WYWVdXXG6Usm8y/RGEoR9z/VCqOT9EsUc
GJaLZkGgcHnF9ybO3uMCA8rpN/EqTI4qYkJLMPGtf88ll87h/v3hDyeh2HxPKQnb
O/BmFYYjQwCebkucf7SdXzxp28jvlTeCBBlGVhFaD5lcxodax/2abrCpGFR1RclK
SoHomxdQFn6S4JAG81VnGfwxY0f3ODUbHqzSn5T+UtWQxiZOlPjylk+zageCslF5
mcniZiIQ0MtWZbsvTFyQ+mtOSk05u51OArfwnZVgRDH12icOZDRKlIJEOLAZhi+j
8qSSp0GbyCD/x9iJrqktjNjwsEhrBlGhZ5HMATUc6pohczRpFchkjK2V3OCJ1iB9
aJTV6NA313PQofEQd1QSc8OYSUoR2TV88xzLOga4bXiOqpRjyn1sPvK3xp4nMMu3
IS8N9ig2bD0/9kUGxoyCFZhjCnwI5SX2axg+m86cl9SqeZv6jdW5xK6k45Y2/NGY
bej/QpDhJyQvytrlFnFIYneS1XlekTX4BY5At49XapPw6+cvZ+MPXLXqAmqJjMQW
FFtJJx7INSqAdo2/8enM6tM0CcCzNxnr/WAlLcL6atQKUGNX7PtPl+iRt66foxWm
W8Au7M2uGac+2kviVjvh+jgzIR8wlgYRkhc722lrCGWKl92yXSC6UIJMAwtjOWph
I30uyT1T2ISrU5aI4ePfzU3Ba4ZJIQEQLD72Ej3qbPHMHEkzFIUtIsoSOq3JJ5wx
Jym4LgZ2s0YqxrSj0lVVtNkyiY32PgDLBDcFQg7LwrNKJwwMJ7JPatGmuUCQWuwI
aXXrIbmXy7TVgK8jsISN7kapL+N4qFYDLkLeZA+wOxlF9sSMq3YA4iIgY28FFg0Y
mJPBF52Kq8/Mxj6Dkwwze//ek4D9/8rB7nYHj/7zEV2JIan9K9vnYe4a7byKkhm2
C7OlkKSUUQcfdTuSSw6BRnjYcvd4ceUi9rS6to53rzCFA0XFmuJm2x+MeQYN+Qkv
AjewfGRZFcTkiAHQK5Hl4gHme2P4lQ4rMmjS9P8o0gU/zyNVMO5w4a9iCN+n3JAa
f55h+1hEzZqpX3wAHODIeb5mDY5X2mJuDu3xt/7z3zcNwEX4ljmHVtkBUJw8Jtnd
/xu55Sy3sXm30dBLFQanVqGbqQxIDCMtCIhipOGEJJQyv67kacbdLZdsWYdwFI/t
m64Ke2pj9uiY/LSc5XooIlSD7ytrm4AEk0miti5gWloIpekr9YeL40Uurx2LF2Xt
udCSgte0Wz2cTRTn+7Tn+qnkwTKcH5weAYJKxsEK7fS80EG0xl5GR8rdWeG+odCq
tw9iAEju0mg+KEyco9r8WxHkeEYANiA1rjKhrXxv9Xg+MjXVjxj2XiJCyelnrKYr
57MXMud+w+42Z09eFxgPLP9LjAZ/IGIHpXxuJoGBTsXfE+LQhoSy+ji5tPzCFki3
GYT4r6HW2C0GuzXBqWXqzXmbQkOos3NKfhFDjMq1QJPGxpGx71hWiXRGUVDOojNq
ifO565eEB73qRehzkTG+hczsrtQMI625pNQJj13K+r0bjcfOVgHTnm09cZy+N/Fr
6MHo8ChmgbLicGt4tZtbpX/z8k8U93SfBW/Z9T7+eUcb/ZN5Sn6venYritHcwF1e
8gHrYoIK1vSKIpLTGPq7BNOekbKbQbwyfqlo+gsPw+5jGgdjczN+UpoQNAVHNyyk
DrR4qLerkGvXi4VWS8pAIGYD8DUmFgEA2ZJGEt2XAFcbyhLdJtXwijQkXr9DHPhe
zG4eHq92vXfh4/Tgvy6FzrbrxXsXr5usczV6WrAkR9embOksQmBt5EUrq599rjgJ
3BfhJHHIP79lbiuypIwkoA2VSBPcR6yB4gKythBgtRvpUWLe3GmHnJ/dCmGfZ6fx
zCJ289exIWnyNGAqD/OFasp+xAI2iEnISjgcmC5SWQtcmKxJqOhWGLjOAxdcmJih
Y2xQMnzhpr2t50cL8+ELWClNiKsQZg/O7Pz5UQ8/p5XCf8K8kaUuBxf0zTc8hLPt
sNZ/Zye9mj/+rTgWy3elNH6XxqEFOvgE8yRX1iwKlxGTX3L4sGkQLUu4d4B98njG
tacw+yMCdMUNgEiOCSifIsm3a1Vo8dxBKXcjW1x10CUgUq5DJegSU9ximXqrRuHL
xHnRBCj2ApqB56LWYqepu+J1tIWWV5KhPp+BMKrKweTq8A40LNH58utShNpXR5M2
0O3sx6D8GIowmwkV6qzNGD+oYTcOTktxmM0vhmGyrBSIlUrA/+zeSFR0KrnAO0BT
rjW3oUHRXMcVjtMJM65vdDedY5dLc1i4Y0nnPKjzCaapc6iV5CyYqT055MGHcE/3
313GIti/V1YT0p6mDULPAU11K4uReJZsEkLtV7SIfFRtTSSoqvMbQvVjVcQWtdNM
x9HUU1zwqcQWwZNHu8ohJ2Zgu6FVt19Xm7B6ZdSrpxsRXgpnduJwCgRIGXFr1qGl
8YDykY6seHL9cfb3VcQjPhLS5oGzN55Lfs5PKWN2sD3z5pJcsLD8xf9GUZev0/p2
phqzEBi0VGl6cbwnrohOIMEMTAG2FVnXMdAJYatG+o1lYCmWOkhoSyR6xbMhtWAI
Jl2o9dB9+WLL6oRg0zkYmmi+iy2FbtcMo2ukTopOhqevXymct4JlQPiGLOCIikDJ
Bqt0qfLzrpxu2NIj8tNmZjbI1HTVGn+vjeiZQ7t+5m3zZKIoCD3R1CLDbqlQr/IV
XnuZEbC8WiiOa7NcCruOq44U3UkMI/Y3/o0x3erQ5cxtnZj5qYyLjflaEQwZrozb
+XJgecWVTetRHvI0hCuVTPBY8eAgM9Vq7fhNxwN5c2u4EGnBxm9gF8Z3bpoDpYeE
N6hTR7ttCHXDKpH/pXwuCQ+a6LkRzKdAgL3l8Mh3GKcra6d15IK7A14vGLXJoOqf
I06d+m3vaQR47lRX0edzqbmI7XQnHyKrXhBdP2kZLhCNjGcM8QvkcXETTl9n58qo
mLy3YDCD7AIx/SP1x+QMb99hvzwB2Bl3vW3tekgNNV/2m1GK4bqtkhL/CvFLZCmr
L4M5Gp24PaOIwn/YrvGAODlxuRhzm5d1E+9JCiAsxwmxCkawdsP2CKlFP0Z7w7Mp
+M9nOCaTm1+2ylLFcXVfrCNzML5R0x4N8pVcZ5Tc7IBcBSkUbEMKLCnDF3AI1bls
pNcvUP0mseeW7qtH/7rz8d1RlzRBUTYmR3pbXDH3X5BmmydIa/jS39uQlWYGhr3H
8tyMDJ8qlekbmkrk/rwPJeJ7lhPSvpz1BhzbXaHBWI+Z3StJ83NofVytr3gecjg9
2FtxVSetZSFh1DG/hBVWyGjAOA+XFDTX7O3JsJz2BqHiS4CsVDxkUzC4pPR5thZf
Oxne+eYHsfjz2L3QuFGyN3U/G0mwJjMGj6wIP8Y2NualG/G7q+GQEnWMb5wgkJQz
vxy83dwgcU8ePWF0UWVKBSh1of9iWzsldmvxkYchKkTKO3SS7lRypsVN6uza8nYy
AAtiiyW9PF55h8gTJxOJapqqmTsxVfgpe+DENx4ko4jNYXoh9mCStVuUuqPccFQD
qM9HQtHF2cMzdgsIzjvMY4mI+LpfVLjJsFWi7bKO7hNz88W6jrK+9CHWH2sNbY53
5h5waN/pzr5zLW/6jzE08xZYZ1mM3pP7qriVnVivALckIuleSjybO0g2JU6vPZPx
3/dt+PATGmKkzS1FpaTF6/9Hng+17oD1CQhsmZkZfBAfmVSyX8RJPwQCOqXXzlMd
1Sco/7NyD/RVpOfX/MgLorwDpwAhsndyitDW2SPQczNx2zR3Q5wT/AMR9tqIiD2L
zH39en/LNcLChZQagqFh2N1Nv8/7dwj9TXLgU/c/0g3ywFLt+l+LWaWVjIGkzbdr
EFFB5jw5HzInziWbUMEOwmArfelRlPH5k3J4xn5++ZodU+2AmCHxkG3W/9oTnCyO
zSxo7jewnSk6Hf+VtJYLXkG9h1hJ2eUZu84SGvumdE8R7da7OAVNpIKQ0GIJUEMO
fLxsxdhqfYbrrC6BeWz4gaYdyGur/q4c7I0BOrU1YzrDMUAjaJ48QQmDz3WiS/is
WAPkp3jS01i6QNfhHEln9wnv4Z4LH+WeNOl0HlOGaSinSBgaCkoEI5wk202mg7p/
DyEEkA7bfYPPaiK8SNLBG7I4mJbtV51YH4AORQu50qEGe9cxjtQBOnwD1NOE+afa
HDJFgkZpMh/DlM9Mu9Pc7oQnm/RY6rWrdfk7udJq6MqcJuhFHWasb8SPuineut0g
/Y+7QzFAZgCnGqUF+COYstgw+wrjQDJP4PiRjUzspR900JKZTVs++1KPcF3kgcJo
5ITDMabMtiwLj2HVP/rSgLyDv1Q3BSf9RGAPDwBL2jiMk+11+l5JlirrhZPwLje8
rxiKhrp6SngRwPwPU0qNvdpy0w/Q32pTU6wdJXiARD8JkCCpSvUcorGvVnhNkC89
Pic47torRVYmWYa5zGMsSZ25jpEbcO3Uk3MzIdrLfV/WrinTtPuGL7O+YGxCaV/5
OPKTwJnJ1o7fTMSZVTDcsZlYQk8Ap6QM66MWUR+MEI24kuyzeosLUVqFoRF+le7l
RGP8u32+GzDW2MrpEDMO3OmIbCOcAp7hoOgV5FFD5VsBWhdj+sO/XqplxK+aWkX4
2eG4Mkm3yq+yuesnPkR/G18kMNrzdZ5d4I0d5Mr/H7ArO6ISYM+ilJDGPTijRSC3
StRxYZyXRkw1PxjFAVFx/lT4hVv/GCNZYd67QL5MlQy5x5obapYcDf8ejRyM2hMi
5yDvIBUXpXPx5dZ7k3qqjtR1snhTaLLdN0BvyvRUVreDwnIzgrKtZXStqesHcn/C
szwjpWNog5IRwYTRIUkMWoLHMNuxRLE+Gk4sNOu836JIg03UBfNOWJpsns9Av/+/
yNuS3LkrMLVGPJ1gQHanXTQNhrP1pVp6jFrNrUaVELgQoXLsN5OvjGrWg2dcFbT3
GT1JUyUxhhMBMLGbGGFmu0uKN5K6JXGq8dRvfkdtJ0sb62xk0B7AjFIlsFiXC6FJ
UDIIy+HDxdz9IUCGgCvSTilxaXA9w5qqfxui3tCH0rjGJzp2hiGGvVs3+zWi6u3p
osY5/zHhcD3k1wq9Af9vJIBa8tuwHj5Kgm5GWxybbnEA5SOguLMDPyFe6GPFLYQC
Yavu/R4Az24dxYMuIHA7WT3cgc7bVHmOt8r6w31ffzK4z5iNeAP1CwyLziiCEv1l
eX6Jqc7hkCkmwu/8f1GCjKFwgKnUd8oNjkjX4Td4kHaI6RMnEWmjbDFPTsgA2lg7
EZVh4UMbpPIF8B3weqtLj+hN5iWP13Rbp/Q5yQCTt/LjMTpS4ho9ofhjSj6J5o32
wvQ5VWa+d6F6BholMcE4Na1Z4ggj/4CHpDPrMF4yCQwE3A87+UZUhinKngdcG2hW
fc2aTW7B9cCG5xFOVPXc6dWIpH2LVqi17z/ZD333ibszZwiXpqAIWagM2ZWm4FfL
fw59cWK0A07gkoGDF9Yp1ZqYr9rpV/4pa8Rdx29CJu5ZczGAI+LbXjNXbjcrGf+S
Sd/V/EUAjV2OxulioRRuQEAR1/vXVlkTjPFLAZcYyIWSVGiazaBHYnVpmNIPNxyA
3EUUz/YsgcIEfB2z1tCHJU0Kwb/6ao0U+Hy4s8R0dDLHxZW1n6R4Zv2AqgxVe5/m
44eDRZ7wawco/w6GunS0i0R6hXeUKkIao5zPWS73ETLRht/rZn8xfbU4pJ6jZ3/u
WDrRA1Os/R77KH8mhR5zYjyUYsMQj6yMXqNYkzuXwkaXmVVkiDzR9Fw/Ks48QfLq
kO2Wq3rBf9x5/benW9MPUP4URcAS6+yR8PBp3xf9FC3ugA86R+ZGCie5pd0oJP8u
sL/Ajk0StLu9qnv6vJ1EUTfnygWpz785GxCvUMdiM73pJglyfHVscfO5NU5w68Fo
ix4Q1FqNK6oUwQ8m/g0mGUAMIpsK/iAFhSt9usC/0A0kBwDKr/NuceNzSZL2zCkp
tRA1TpAibkVJjSEb4h3QSZx+aTuRe3fJT9Mb3jtqCkubnRkkKlMlTvn+9t/eAtir
qUw5qLWOQ34Qt6GPxpiRe638vTyqBhSSOZ0Jt3a0wZDZq7ce/Ca7blaat9To/+XH
yJNdA3uHvtAdiKRbBXfyhMey8i8BQfqmZLZdhlhnh1z40Sj1klvwplberMN7+Cvn
aFfodzkPYEM/DGZveVA/OJSl1Hr2NzHQ2AZVEGkuZIW4MhzZui5SncPPTG7l6kY0
OL9zBJtpo3JOf4usvztMi82O8Z+QkDYQtyqxQClY6CAgT6tbdIGiOH5S78csfLMV
n/4xJIzXRKNmwGOXRiAQwodGZaSbivYDSt6w3daGe1kRC41EVm+azcVj2PpyDg+b
Zq4NGwLuOUzNc5b9sCyoBaUJoEL9ldkjaasBFYdlbvDM9sZALDASFp521NxW/Y6R
iqU5JGcq6sGmi8S2B4NJNrFu4iYGIfhnlt2aBW2InUbv+eZwMqljAFRLVgDm8vKI
zY8ab8xfKQz+nSa0WVwTaSPAspM9rkQZuMKncYvH2e8HETFCpuqKlMjCrphD0VS+
CGBzyEd/0r+mEoZCmSTScfKm9Kc7DFan76VkKex154VWrXP/AEkzfR9f7G+zK2Cp
sXKq2Mb5w7Y6mYXT9cCY3i+AE52Feh/u2bmhcnk8uOc3HxyICPKChcEy9aWweCNk
UqA8sa/GcWVi6b35JEIXNALQ5IrKqKPl2BMesPbdzxFZxHLYlagemWeuyPaW7jpN
S04fAbkYWicSk7UYTWoM/IWk7lBNQtSMnLIzgaOoor8n4gD2mZTWPdadz+zZ1+ET
X7n+Dj/+EmOlmZ8vxrBYLU4D/dwpAdSBbtt9JNzMbl9b5TjxSqt8PYjxR8afA4X9
DvfrvQaH6cyaJov4Eoh4/2nKaghpN81+ukMJZ1uEAID1Jv9hEcOvm1upZIiiVvp2
BLneAUSwhbtJyuzMopnYVdDobhdrwvca+R3iSXb/gyDglOMnCDkoADPLwDVWhEKt
+Hg6OFHkSTtLP9pvDtLDGiOSgitvNdCFQ5IOGYC74jAbETvzyFM/QDBEqdOeHMjK
54RwBm3bSZzH6MuYTiXSaW4pK+5XsY/R8FXB+gECGuCBGI6zOydJHXmuSOwXENov
atFSfBMTdeeSG8f1EGgr2xlE+0esRcgiwEXPnae9QSB/NzjkK1kFvJ7PjBusRW1O
EpXGDbiwIpA9NgwI+cATJwMicZ3BEHEriDuoMDYNZaQu0j0s3ytjgKJqW0hxsazw
Hq/iGlpHmyEiuBJIxQ0sTskFRdbN1xrIFMiwucq7Rs9F8D6V0dqJwY6P7ErZLZBV
4+QITrKUo+1KM1G3T96c05EhHeTjaU/kOjKUs/k5DabkkYU+NyAiU8kbO3fAMS61
19hQVXsT1vGz3TlZ+7KmELYfKR2Wr+683O97I//reYkXIUjLNMG5vjvK+GEIWoTe
Bsw1ier/dplpoLMCMKdznvyLle2dSTaFnUMFBOw/kdEuNP2FywO98SWQOqYY9CO2
9ummiLb9c91XOqqie8XTT/up52pebKqiPe4q1gPwBQel+lbmRkBb3Q3D3hGNDu/k
TziAV8bpL4rrJQKLl74YVtQ0bMVAh/cXKwjiaSsDC1poZm5XThl8/nPBrYMqFn9t
dczNhDUIvoJIrgLTZu6xZZLdmY1G28vbWZJnWUF95d1XqbQP9LT3dkbnqlblG+xH
0ZI4avMpLurSiqhy3FNh60XpcGIqqFji7Nf5uMnOqPUNvP98K6+3/M0omceUg3Wk
MibJgKf8WyzUaZnOJS/MF1wOIwXr8T9A1IrPE0cvgXJj5DvKh49vq9AFIxsJIfR4
84cQjlVnQ5VhQgHqLkvJo61ljisSM+OSmtIVr/hd4Qz2zxKpXzyREsNrRRdlZeNr
ZeLFCfMJwtHecjZyp6QzuoKuXWAnyff4Kqj/tFdJ9/rtzPlL2nehwI6wHfo9ZIPh
5JeV41B0cV9IiGA80fGzrQwOCDSuD/lbGbH4NXhMWb2lFVjtoyyzzuSHymEF19NU
V3HJtkjPpexaXQ4dgHW0RLM49wWoi7WwJKainuu/PO7Y7g7fPtU+S5zS0Gmr3uTp
Uo8+jSaY6vFVXmUZgKe2zKheWc7WNeHCTHluepeFZIoRSMi4jKzk8ElZz7fQZ697
RMHva3lYoajC/g4XXgHfK0uA4DhLDRjTgxsMKGHbL4BMoaubXqHAiKj3aBhFXgrL
h2ODXRxRsGxaFnDOAvYkf7uPrWmOQ3uoqsqmzGn2NasoxxfdsKVgsCxICNc881Xl
9m+sx+3cWiPi4b+bMINCvsjB5Uvzi9jhdTH12kNInZSzJ0V/TSp3ggrsictIZ71W
yzRGeedvyjRN/PWWhI7+XOM3KzLa8davIV+BeeRuPXAHHhhKOFN9B43+RwFu0Anl
Rt2WyLuNz4fSCjQ9X1lA4AtZHgaUNddX6KRUReUSqgoJIDIxXEoP6nviOWbAux9w
ywwqYvCvwaDbD+UBQgw0vWHHbHObJH7nj/9uISnI1vqalSdLcoXwopVp4ay1Xu+x
t32D9OFkWPeAp50qt25g2+zz37bo5XmwJ9plI0aXmi9oXpuf5T2OMDAQ+WuOnwgU
QCRlZKinTaVeUMcBiUI39MX/tX3qFbSjr1dY0eHT40xLrHk/730SYJ/HVfCR0ptT
JKut6cnaodT/+Y/yWK7T/Ps5JS3rrqdq74n2w8+FdqKunZSk2OGcZLtJv7JPbl4a
dM8ALWC2vaGC2tK8bk480DeytRE6vt5QuRXVUQXBwQmXqnL/K7bCEJTmF6iB4jNc
DqIna+PTJYfPBp2dHhOitTZdJ/xZc6aKTd+Q1Evnv/x5uQde7W/ntNgrkm2sQGnM
LTJzJPqbmdKKU56CVG3HOChFDwwOcAPzyjWXmjrHn7KaLcjF4GqvCv+UNTsCS5YY
KOyFcpDa09N3vPGrlBwSLzAtkMkz1GUbAMMOlyzvzJNu3xl1oUaW0bl+zhD5OSae
y1WGtnlOz/SNO+WPzIpwCBJMIh00CTZ4u1twkaxztCpvYKq5JtNUsn6S0Ly07Tcg
kyeNGNesMZJTNOjWBXD8+wEop09P12d/o1WLYLZBvhuMWIcwURCuuvMI1+GYI1Ou
BTwsvWspj6OALH4LdlkiT/Mol2OpW3zhd7exMbEwWGVSAeqR638dJBroC88EsXR+
cCk92jWdYAxBrSRn8G/xS4z7YW6Lg19fCpEDcUse8O+0SGymJF2zs0xCmNikNQCR
a8VY6USxmQ+vVXX2OOFYpdP2idl7lZzupjARoxV/Xj7K210cDvYUK19KzodFVDbi
/zMDzs8MMHXdg8vSshNAI+QbODlJO1suCZf8Rr74SKIGMt3MntDr05WCb6G/FLC2
u5j2TQprPjtkp9OwhmK4rGIQlWt6MiSW8x2HGGNt2vqoARQyYrKq4yAtsgtlJhA8
szHGE9UBSyMApgLQpJDigljIVmlkfQMJYGE1fw1Bi/2ZSD1nWvKPNYK93piHMkVV
S2+QCJO1FCA90FzslzvKRqG1skqnFWEb3ADhE+RutyeGBPyBDvobsUfaP8HwHL0/
LfpZGlf9IKMhA0+g4734tEOSTsLuAEQ1Jf667VxbQEjipKxIRMBb6L/RhVRXh7Cq
/lyF16ExgArNOPEQ0fNy7Absa+7ifNyDr0DF4lRr4gcUyPMu9hzLp6QwH/0j9Vu3
uzQNBjHIKExk8y3aPya3q2i9TXOOcXMdTND9D3JJq9vHAusfgxc5xWe8JVtDxZGP
IXwdAACZq71rZXSQvJMs3utLwouaDJ/kxYzxzJx0YgnuzQYzm4s8exBSNb3N34Jw
WYqV68xOMeHdEyGvANBUOGibAg8rscrjiaoEHNzw2LA1QQJlAopB8tcl7oQ6xFkC
l//00WMrqKBqwhtJEL+hkZH+d7r6VG7UhAYIjALWXKe4cEmsQFskfsnJQl8/9fnp
qG8q7qR3FUep8qnl4Bjxcgr0MtW/xJQa6DSqeXAXNYg0YAfxQRwbdWxNpf5M+qq2
ECiWSsSfDH3/t0JTvZgx+T3rhhvMPbc2DwZRt2/bS5rKk0o9xxTAfy1tAiE1Ux6Z
/8dUAgeKLFVBc2YCWMcpzr86Qo5B1qp2lziVSX9CknLaJK8jXTnc642e3qgIJ1RW
x30DkMb/srNpX6PEAer+jjMl2J3rhMG6X223jvJnQRr15/SpYHRJphUcgY6ZW/r7
aSAXlENNvv3iKz+LnxDRIzmme8YFWASBGmUoARywkkooqSsbiDOVW1qHnMCfsMqf
NPlVeAS7zZR3d9PfOW0Rr7Vjg1tIVf5wEsPWE5RjHhBAQXcQnsaVvK9IBbt+WwuZ
ZFutyQXKkTpx82UI2CRCNiNSIGFja2YT41Oc4n9Ves93jtqgOJ75N6WdZ4lIFSUT
RfxyeFu3cGblBmk0YVBid3r1eLaCy8MFf0xIBERe9cdOJQWYX62iCHXUqUpTufsU
qafw9XxoF+nw3OK8eQxCEnTNUsdleRm3M7+BQQdtlh9ED8Zd4g93Sut1pp/4dKmB
ZAgF2BK9WZsiK/MvS3L+vsgCMbwOrP9gizBooNi75SfssbUxTipzCegRd0m8U1Iq
q5qarBkByLnoFXw/edyWpwL0YakPMo5F0ZnCigcWxeKrmeGj4YGbHE4qcAJ7IZNN
qX4k3CKQsA21I0Uelg7buC1SdJdfbNbv2i9q1inPvz49y+1R/TF66g1fBPiyUCsB
bwoF+/op6tzJm8FOotRQ76E9MdeEMJL8rIYnDLtH/2yWUl9/r///wma13JcLjPFB
m/pvdpnhEWJjQIMzgJ0f3K/G3AoCMitr429aFLiJpNO2yft7+Z7FtyDVvVy3AwR9
Epi1aApub0cIfjxaz2VeEJ74t+haNPT/32MpM+2hiIME3tq0bo29Fuo+eyJmgtRB
lKN9cztU9kR2HBfwBVq4o05d3aU26VdNfvPiZvWA6mYydIgscVlEacD+zGaSvFZN
K9CsQQV1ZSg3MnSCPnelLOkEn3Q0LJgauvqptozaCBvT271UyW9+V0L/xhIEEw7+
R0VDyU9vYrWzh3RaB+ayLduqBDhmPhzqyG6Rf/iYqUrfaba/SuPFQSv5pJ+ViJS3
hwM98AGTxXUdlrJFAAbkBd2J5hBJmct06VCqUSFF35yk5HlTIic06u8jl7vj8RLq
+9dXqOgLUZ2sTpxMJ4Y3cYaSc38zKDovdxIQ/2KOhmOLHzIQQ9SJ5/km53sySWxC
gRGHFhtYOkDPgegYac8hZuIX24kyEKaJz4VUD/8yyQbKeMWeby42lpM3TTXDn9vB
hDfIaeRo0M3n9APqc08Byr6gifjb8NBrJ4x/XA6REkSnAdwioJAj/hLOrggzjXjN
06zkzykNVFKLWYpWA4+axBgV8wdv5DgNw5uDhGeHfI6auKOCPIzB6xQDJRSDyOhj
bY5TnAx202+kNV89ZzyEI8QkOoq15QgYwQ+18m4l43lBmmOsCPcW5I2gvokJI8P2
0/1Y6nJAPkvsCO9X8npaFkIBhTUxQTcIdf8+ylUefta+mMywNxLMzDLt8ZaS3Ipj
F2d9wjejsR1+BIlWcr+PUAl/KwafvN2+RzkV45BN4y88Pa5nJNqGYQvURW+AyOfK
OeIw91JWaT+9SDkjGv3el5+HbWPbFEFWPt8VeLmLAX/sBS8LKGAPmMyNcVJmEx8H
tem3OIVkkgFsN60HTD9YNDwkQ4jOassJWl/rTFhsPfiM47uiOHTveJziKahGcpRb
yVBQZ7nTib30Xu5GGRUWgI6Gb56z6+0oPGdhP89c29vbaf8nVrtnduZWh4jPF8cL
kza4RetMjJoRL6vV9kFk6oxXgv+I4DmRLTykmiiUBcN2vUwWR9z52WkDKpaqaGsn
HY9x5cwkNHvAr9DealvgU7Rbmycd0BoUykf6Hza0N28LSjFNqgWg9LlCM4KAlhwQ
yikkP1IsCQQxs+PNSssZwGvpu2JwMpl+iFmY2tscDwinWqvZkAZY9bcXY+MRlIsb
Paw92Eu1mH8rwXNSdhKhSxN+lnsoto+Mrii+WjrAQrJjOuHgx+nlWjsVDoHT5roX
AfkwtWEiKrogwoya5uK5iiJm5pA7NNnCy4WqhKPm4aMPfFcgHUQRiXuuHup0pJRI
ctBRJXcvkYKuY9dFuy7eIoqDs0F2oWEm3lrIn2vV7gNMC1Mz4YRrdpeXxnerJStC
0j0jNLnga1SnSOkUlmMmNE/eN9TEyjkA/gEwHDERg67iulDy1Rnd1mDbxivcs5iy
WJy0yQYrylPY3LWliqgJj8Vc7eV2UmVuWiaATNVgq7zLz7LkqMHO46f5DjThG3zX
ipiYJUEgLQLSTV04wVjL2BjUROVdRivaFsyLeRZovHgOyTvXiRnOgIr1tb8tsn+F
/jDxVjwJRVeBxlw19648rFpwaAXve0Fv7HGTSrqxzyE1jVSfz39tpnEWhREZ/LwB
gDCGVokm2iiDY2esg/bUwXcauRyBPXjIXMDtjzgQ7AAtNDBPB2ZvVmt+Qc2BJxpF
jT8Mg89KOOI1isyeIjMlSvbizpBoAdwMtrIbLp6NM/bHYYD1o3OTfatSMA/dOoQV
79DcDsZ5uE6/qQl4tt94dAcjgN91vjPMdlhabM70NcLPaVkVfj4VcXeafGgi+CqO
25Vs8Yoy6HtPAYuMxpDmfrfrr+GaYnlW8aSHFDJWrO/msdkO+4bDWJA/03gzNw0P
M3koJz73UmkM9HbbxeWGg4rPrZwgScbX/VkUpEkhwBbpEqroCH1DJrCmKsWSl/bL
7+nycYWawn+wcjtxddpDL9KmInOfIQl6uq01mdZaAa4qMlIunY+oFOmW4X3+W3YQ
l2MZgk+DxBtJ8idOoG16rxz1a73ll1zA0PISqNBJcPrMd0i2o3jcd8HKhQBylK0f
4PXLxCXVXphgFE0iqsNwd3OLFwJunLIjPw6GxZEEbaq+uAt8dHgIUkqbDYmhttOf
JkvX5vwU1PmE4MzU9pn5Ea9OgbVQOJbVto2BgAAbxgAYSiMfMmRUcVEOyEBtompk
AcYu9wS9CWGkphom5m5ENOxwE6/ceMZcXOx6BMhxcgu4drFcqMckBzrLdjawgFzZ
sWZfjzGuJ6ckYxu+oQTOc5lgU9RtUZ5BNzop3yDB0TFoXscwq1e8HRcz7i17Edjb
GOnOwhnHuGDUtdetGWqLwGuAnutSDDepWb3gm79hJoNRnU1MacUlNf811qezKhLf
TuB02noKSTVydASsaPSODmS6ICs1yGEI4HpLIIccnu6YL6LRSIyVVhVkCfjoWpKO
W9chDMCcqbov8557vMx0uUdnTZ8NYYtPJAG2ZIg+NJ82Yv2REzPSM6Zcz27KblJg
4dKPzIQeHQqUA2VQM9iFvfnmL6DSKP5msNX/pUu5cc4eRI6IyBA0bGDoDsp0rLhg
BDnJAyCOniEMUeCS8fFxgI4+XV9XHm7wtrhP2Ml+fMy+kq4T+NV9WFV8v7OHq9pa
g8rnVEsVtVkSq3el9KC0wwZpDDtsdyrFb9nwmRK9qbjwbNGLhdIWkwy6V7pcDe6Y
ITQgwV8DKLRvM8qx0L+H2Zm6vkdKBzi/O7jWPO8HXX7ahl0zam6EzeQgY24TxKi/
CAgEiKGqA+YEuNLkba+/u0jhOuK5tq0gwoINjDu9ckwtsnX8hJJsU7y0bMYVLugL
iwNSh+reT0g/rIO/1oDSHMw6FTX0ixuSIWncmJrzoCXOhN/EFFGD5MDxNSml21JF
kdb9FiVQmRB0U5SFfjKoMAwDy0oxj7nmQogc6xt4A3yVakCjHR/QwpcvkEfoFsRX
NNerjPAbXF8ksvpQB31afP7gjaisONSWN6+znvTdMs7rrbpIXWNUYOpl/QaU8B55
zPjdxGs2edUMI1kaMmpzN33iDij2a4B1//KG6sryhKTsN546r4CVyXgyV3NyzgsT
KX5nOGIkBoGqARw/PWabhuVRsOBRP+wdJDe+kQzFNsPEkjQViUF4rH5mpnt3n4w4
PsdkXxUruHtcF6Nq7AELGhmiRHgWSA6OZt5H37LRrweM3wPIBhzZ0iTDfhbwlbMt
Ccsfr+kO44NH3tzlPptqodlvVRAJQ6epno0fR+6+f8+sRybUCirT6OwZCgJpghHp
a5PGgW9vgLKY2W55YOimuLB0oSU786agY5hdp+oPda4AIbj9LI7O9Oc7rIvgpLJV
rjByjJJyp8qz0OUjhERmaX3sps260xuUAofpOCQYESLbu0XmXpGqyTmRjyPsEGUO
x08Z3vR6oluwH1PtRObQ0yqQaMnxWt2UkY1INQM9v+ThCt7x5XTgLXY+BLYiHKNX
YKeQquH6PqePwYTHB1ym502gs3ybiQ1kz3jsLGcL8oVN7gZ2PEuEsRHuKsrdAIAf
JmBUzq2Z7PlfxkOohsXCJAf6oDtCNz089ENJhzGXoKZLevNDkoXODhRUGPvqC+d9
j8UNnSNVmet8gkhty15aUTHN3OSgxDCvQFCkaOKxsvNqdXRSf7n+K6tu4jfDTi8W
C+c3VKEnqsDYY8wCe08IdKCXknPYffg6SldVf5TbojgtcI1d//3+b7ELUL4plfk1
4nx7UHe53qYiq5SWfJg/U4H7Qm0y2ewM4ds0MOEDTu545iaFjOGYVnaIS4khgf4L
epXtG/P8a4ZNP+1Mtcw8GNsxxHzQdafSV/LlrVEpsaQ+tZf0Lqib0+LOjKKaoZGG
oaj5nzWJV+uF46GnG1Zj+R7oD9L4679ETIHabX8KVzS1jSB8Gr7Ihb3/vuLdsXlL
y6bR7J3rkTNfkgrPzBI8PeTmnX9fQ7pAYIXWZgg6vlk0yYIh/DkiBvuaxjkmDsGu
u2yAEsyfqycPDCwoZA150kz4+dE2hRcPfQYJkppdyAtF8+oOpZLiK4nvg1nOv4vt
OmdGW28pgmXDZihRnTo2L1+QIyRB106xe4Im7NpRmqxpwM12VfN/9p/wAvS0Ywj0
4ly+4W4I+KYMVjO/m244iYS1Y7IDztptUFKv9RwDdFAaHOOMHyWW8E6zigVeVBWa
UhUkSF9P/3+73WvRGj80gEwnOGbfVfq4MPTEjBSpNCqk1QMKYoCZBwAYNStg1VPZ
sKCbUONPTLWvyMHe6uXXNeBanE2iykLX6vgi3IQp7hDBtjvoLQ4qideOHRMidYuG
AxrbeD9w7Y5N9rDI/e9HJ6XbrfHuT+NBJOiPhxEsvgHJw8V0zy6URSqMsUUFh8HT
9TBkAMHijlt2bLktOCKE290nwXAFUGQ17umZ1S26oIUp6IreWjQr1Z0mzuA6zqgd
Pb44EwNUrLcPK7LlJBsG4jlR/M+9fprHav/NldBYwCM/DU+blBi3bwi/RTOrr8qI
QY3D/6xocApX+NisI4/aoBxJLeStmMLE0PV7nyDNHv+dSn2fnzEN/zj8EcGaZzsz
XMK8HDt/90pN2KEbKdmT6LIzdXPwViL/8JY7W4ovpX3e6pMAKODiGOr7/CUByrUs
CABAkEarFnmCU4nasqPDydprLgNGskkU6c1qB7gw+C7mrUmKEymbxVuOiXYvU8kl
75KkZDWXIuTR4K032uCmigW+qa3F+5jpX71KiNo/UNT+LOR9oEGwdIRnXbyaFeTJ
/HX/JL0Xi+qXVUqkCrW7x3wdqX1B0yuKYN8m2/ZSsA2IK/aWSyQUgl3TO2cgBhoD
23ncRbd0W7JPWRyGs1Cl0Y6vg8ikhq2f77QydhP6K3+EtGPD5oAhN8gI1QD+mgxA
CHkbITlOVj8F2LscyiKV+vvWzj8P5R1zk1J5vispzj5oYTe3nB/LYKAom8V1vpoQ
Ng/9xde6ZVze+5K2vLIuWEcTuUyh0SNMP00s2IK+w/oMFYiUJ2jcs5igVxF8Bqo1
EfS/nrvkmNCgH9kHPlxp9oFhSDZinQEiFGcmr44LQ6veCcGkm08l0s/ZIwZ4cwvi
WW9oBoQ1wu4N50ntIe2uPVPv9EjGhcKtgdweP7SH89dX1UGaNevr9UsM6dGNuDc3
kdXbzxfDjFkA2OB88S6aoozMK/B/+XGmX4AfmSbFgkRWUC5gf9mqQk0j1CME03oi
h5oGYdWZ6SAU7W89VNzuuhClrnR4MGYF1WUlZvCoFXZVPaA/B64WhkqszxWhOkQv
2naqqOO/26DKXwfi+sQMgQ9achb2/fuu8mmzRvyQOMb3EwP/ECcsmVP64HZ93adm
HzsjmPiFqHjOwWkaK2/E7ItyO5sUTu+vwQEGonT1M48MCLLvBQfMD013zbWpi+gQ
KMvu887YebQTINLWUxxEeQRMSCrqDD+C3NoPl/gOKahsCdNrVIKEYY0qlQ+VobWF
HHAx8ExbEnFqD4dGGmahQSYZdrGW1wGtZnVDRfMju9x3OJyWJ/2lKzyNj7rB37uT
qZ2b0PIM9cIUUu7nGSEDyhSigBGcFNfZhAl14gRYi/C+vz63cbMSmahAjyP+m6Wh
bJPyVMypzjbtpN5uNlFaEHBP0yIgk4vZOBOSXD3X8brvhM2+5Dvz02MpPC9I4d6L
638MCNLvGC37sZkiCg26770bmjqSZOsUeU6JzdrePLpCeMXIxXuGqmF9wHpVkH2c
wb1stHucFq0jH7lcy86hXH/icb8I4JXfGWLP9k0PSdNRRfLDiTLG+WTnelInN1xx
mB8LiMocCKc9AhpnRKpp16Dv4K2tG51oe5ei+oy+Kf9U48dDY+9SQZltifa2lJDa
8tZ7Bt6xFxaQJQBOIlGJApc+jXMiz0h5nczyiBGuBOpPtKrDIR3ipJEH2/1zlwyi
ws9IgSja0HW0kmx4lCa6EAzteYwQ+GdQjouHjh5Ia3oHA/kVntlJF6fyrIpLuQ7f
eYLmrjdaVfYeYlY0+Ly9TCJFt0e3nbBT5RIJ8v9Vd7wu4868QP58demxaillX2H4
GqTLZXm0NjAIPiFiNQQU5HYKGmprP7vvtUchRkcxGWlaHsvhPvgkw7X7IFbVRCPx
06Jvm/X9Pez2Br4CY8j3XpI1aONs0oXWOvOosmXCJPCu3WxuriW1Mvw6V7cAqmgK
jNOdElJ3SW9blEm8AFbbDqinEF0PCcm25JWqfc94i7sE3Bj1e2XuzpZCIBn3XLP5
ZfTwRG3K5DfvEGW6PTbrxHBrPMC0HUofxz/RiPQ3BlwRpmyvTirzrNZs0VTvdqR8
awKJr7Iys/8808vHwMkyFbgsPxC3cE0M0u0qCFazRy0Aqw+dRY6+wbQhC/5f8QWN
Br4SWlOsOg6BYRM+f884sar1m/ZLVyutBSP4636KUKqLhAqAGrC/mC57FoGNwARc
jM7QtnxEYQB84trHDmOZu347QfvKPu+Q5fZ6XmvEWCXFZEg2KekFB9djYsIQgq10
qUPJ9eyKHoae/2dQnjkYkpJx36OMitVsgFLQHN2UntgitmR9RzOJTC7Nm/i1tZPD
XLehEwREOgdUf36AfA7/Grl2tbRe1IlBXzTh7YnQFNqoXimTI9l2a4p44pCz3CzU
rX2QDRNOfhIgW3lfbQVBGeHKyRqbbjnsjNT26cPiszzAMnj1F7zkRCcT0dv2gAXf
xwqR6s+PqV/ntJ94Nb+DBKQH2vCeI33dCVXsLccrV2m7TYaq2Zk/iMgr8XpE1PqE
+XN/C79WUFj0V2i1D2M+Xinqm4tU/P1TDGsv0xDEQmd6XWomZAMMzCBw3bjPyphj
W2Crb3fa6JKAfmn4AH5sdEA5SxJ7+o9iL3wllZhP0YmpBfn53E5tSIWie9KqHfep
91ryh+10aN6bzRx4/PYrEe/cASW9e2pgDc21+TYEXw0+zRK6cb6AhlAsDeEPrDsp
srwLbxOzrYDvi2WQqxhVASj1r9s36Jl8feQDzgMoj5oOVY1hEeND7WN2H9ETMC6e
Yzqc9WQmznNuc/97M5v9qYQIInzGg5Rk7ZjRB3SlJmfVVeqQ2oPE+a5AkHt8pVlt
0J3IPIPjE/cIPycukTXWbfBlAIXPm43NdvuglTM8n3Fg8zGmr+VCxuguv/q4FZDZ
L8vv0fFLVcoYJo/y+LnOLN1p9DsURqygcSe6mV3JqtgrXwBWNv4jHIJ8DcE2mbhQ
mgUexfouQKgyE9Bexiz+47da3sG4Dn8zrEEv0MeQPz5uoxK85rbbWgOfvM1pn9jX
DMTMoYowFJxdE8ibmRKxJFKsvFxj+TA33lZ+1QXl3DqrnIK9rIrGE896U88/HLVZ
5F7L/tYy9OXW2htrym/pcwRgg0YxavN3QvxvSA96U1xmZK1BXjlmjEN87hLysRWH
vGFAq4HY13xLk8V5V/vK8prtFGMJE6IRv275zbBLygygnMy+ofQGBNfyk+6JCUuI
sOwFgTVGNfXRLXIeIU1CKIQvjkEsT0rOK81g50QinC8NHgFmCkbC0riElAvjf7rx
vRNRFeFF4HhKK8v96HqkuRT8cWGoBsMy783SMG1rah596WVAyExSr41j8G8aIVni
GXQfd0VMCBq/A/f4KjdFwBGPqAdCAX47z9tHy/OO41h5hnhoEs/+8x+Zv7/iz4Va
wie3/hNR99BUpCBMxeyuQsLbC0ASE/5x4eoAT5xJxV/gPTOhCUTGfvaIupjPNUUT
/z/H2JM09VtL8gEkVHf6sERBtMYfUYVoazpSw6HXqJGyjDAfdxMF+sU+OPk4HEc6
2cGQhHde97hSbBWQR6HYMQcpI6qEEl/kBXqd2aUmChP55EL75BBkixh9Y74/Yjv8
QUBC44DiFWGPACyjKaNhwwtZ92n9yrL9rnTOkcoIEOPq3qzEoMbrZUEKpT5iMg84
2+gsCrcGdubl3o6gFaBeUSNy3kedefjAJtZkxc8zjpq8ulHxaU/ZPNW72f3Db2Jk
pcxdDAfRanhj6rWA16hl/wl4ZGyGRNQ+GBhM80joI7L1D+sg66RbB4skliO7qCDw
ez/sxmQ4k9Xwp0l2RI0WQdhCx9ljTnA+/A68pMWCGlbXHpAK8G5UgEyOWFwpLpRu
DE6+tGRph7ocMKERBLYDWINSa7TWQ3nBrCHpCMJ449CbIwfrCk5bnQR3OQELPVCa
WEfij9tZkGggJWvbVcQbrpGdcrNqdlmFqPeAEZ1afkTZ8pfVdndoQOWevidFB2wE
E95kydVbhC/wmoxKDSxy8jc0IExU9l5FqOAhfLvqxMPkqTkBK9yTygz/IcqkF3U/
DegCOcZ6A6qG3Fos54wUbHtyz3yiS84c07HyRYeN4eunlNH9RQzobLeZ0684W5J/
OZNW5ghXYXeRczHOF7kP4IBbkP4YVblReu99R2u2RehnhlUHpcXRb8tUdpIxLzii
5hAw+Hx+JYaA/P+GMzwKkvRylCFwdOwfvo0YBR6WwvU2GcmHnGiUakLnAMJcgQTR
VreTXt1kP8lZZuXDI1mQ6mUk0KYvOxJPdmnDvplhUmuMkXBxZOznPuMQWF2iVTqz
Pb2Yy9yE/126srvOuKLba46YCb3OU2l5R88CJBopWPAQXV3MfIJLsSMCWwEi7RXR
H6A5MVvikbFM7f8+QoV1UoZIfRd8mvg9mpEuFZlaN9NnAGsyaZoVZCPlyLGGec2p
6r7FTEX53GQ4CKsJKIZ+YhtJd5AFzLl6i7URWfV2Uy0eMtUpexRyE0/3oHo6yTqa
pSqFcPDQ+Io9Ah1zzky2FQ37HWitLgyAkJryJksPxu6bPoJowdT6wMnjWUeQvUZk
03cVwggkhS4S6Zdm0VYIwAMt4NvLY6m1JEBB9JWcPH9VVoIT58IckQzVmS2uiA7l
jezOd2YvZ6gKO9NwpBNd1o0zGjzkTE+CFA0zuyG43RBFdXVSpL3TeWoUTUSTHzyg
msiMIJ1M/3QZa5z1HJZqGYnuOfI1tivpuKlF6qAfZnNBWKGyGrsyNY661Ynvx6XY
+fTX+zf9oYwzrMUmMdhYEfTEnAlAsLOmxh06X+dU8r3nh3Gzpxml5ILvXDMI1jhv
IHIyNtWzN9UgD8k5yJkPdtQk1Dm4jVr1voL0joHVABXd3Z93PkVQh2gn9rV1tyl4
QO1ZClcJVuxB31yJ4bCGLJ5CbsmcODWD2gO1+05dD+aEZMbRowRmKwQoHhltW990
TwDTGv3gz5nU3iND4NFY8awUtoudz0tQ5TZIEM+ZpknDDsHslALrurWFemJWq8Et
OpTBd89sJ3JwSmol+wugrvFXUF+sBxkn0fThAEgPBwqevZ1Fq5gyrdOe8aXDUHEg
wTQ/m21L2tDJTj+dIMqdy51sPOcN7LFCcWS9UG0k/NDfI+tLZDN0JQ3UV2q0XQn1
N2gsURL/kWLSS2LjwTGZ4Bd9h1SNPm4zIucM2/lECfo5geg9SGfg2CuGEy6Jcn1R
XWQ1HabIlde99uifD/AIi5oUO7AVgrrgXS0cVsI5WEey+peYjA+E88iwOJkClvoA
o0tid5jrcFcSovINQYED23YeZDm+froZc0w6Lpzd+9wDgc3mu8UCD9g+m48b37/V
eraR2S8wOSUOKJw42DbU0/7o8Bb9LHIipB1G7+ToTkPIj1FWM2r1OdTkzx2bMdUG
VOoItvkfKabTYnswimi/hqqMH5MMb/wzIXskEUdTu8UW9/8XL0VGFDDtrPy/7zz1
fOgE0TdCowKmzNQv4FsKXI7TV4AhdtkZZWSYvTVh7wsE2fuYGuUxx3LYa2vLcIND
55BaXT+XpGXRSfIKj4ky9pNJTA7iXbQrD8FKvb6H/jykSsHZvLgxnYJZ+IxVSBXM
fGyfcyJ/CZjeCnor+V2lNhvAMxm2etaSYyQVx84YfMDK1+5pFY2sP38m/zOBgCD+
+vtoHZlDtO6YzicjdSZlYm3M6cdDyjRnV/2zVd/OtI3hSupVhtC7guRmAhHxTboO
W+y+1xtbhlKLSbfRP16yc8ffemjw4oGUqTrnQWg46yKJMbyQ0scMv1QS2gomniNY
DAJ2dZi3helZwDOA5M7RGV63yS4j6bO4k1AVNI0kAFmQGE+cPDgDUiKso7zySZXs
fMF1M+2b5/aiyNgtVJIPM/qIZ574T9GERg4pLi4XxE63SR6UXzdundo7NxYBXafr
XdKe4bPUxsvw0CHUjEAiBIoJ/eR+rcj/JookrFho6jQuz/023T3rVfDhd2nHMGzg
4ZdeOlFQl3gASBaNoSrhdYZLLgu8clr/zEn2i1FLjwTBjlzSKgnG3NMHRfYjn+9Y
fOW/dX9ChM33pchyGcPEn3e7oRn83QbPQQ20ZyHj6lsSwh+4AHhtavV0omN7KnqE
CLHN8WMm3DK6OUdhZv0B+LVmCx+JokmmR1xKMfyxzMIYUlIAqvcR8qmfVsAqe4YP
KOfJk7Ehf3JIIIzzMtkDqLmENm54HF58TFBNDTd4HqEpLHd9VUpRfMrCT4hJhlkj
ucmVa+EutXNcOjkS5pGGfS7aQEnCeyFslqgcsSKVkba7vHikYhUrp3aBVkn1ca6/
raifO/oCVB4SZPKMD+pNpPcVS9Oqj6hI5FSM6cWvnfRHa7Lhc8C4t15bEjrRk3nn
i01HJUymrc1I9XD/jBdgghJJkacnBdBTRJCXXS4xuKIY3vc8nHnRgETEuTs4o0OT
vXdo07TqQYFZFZOOmc2JMy+IZfqUecgmt1I2uIlOsuKrWZC+IvmbJZiDCOAOVJWS
H8U5kOOoRIAoFnE0gbRl3NAIijd9VKk3cxksQ31qITN/Dyvqgw9ztd+MHTC1Hy5G
Y6V2JIGdigVrphPPC7nehIAVjSQnI9z41JM2j2CuBMIf1lhTgX84c+k7iNDZrQn5
yyNCUcBp67QPw4dhMxqaDUM0/I8XkzEuET2t0i4ZQcVH6epZJVToav11rI0+KM61
IFnFiU2PP8RIR8EH6HS/NDgavl58qRRQ44lqCRp5QB/DPiydCgjuEsBCaH6gi5kB
7Hj/798TVLe/7PKgBwYAaX7HyrpplG9WeVgcfWKHPj3HH8N3iZIWvN2g0ol67bf2
p4ofzHJjDB1vhVi24xkiYChaJPMgYWMh6+jlnIQcP0QRuHZPCxUqP/Lbr9BFDuPB
3HDIsbva/mbYXtBXKK/VAULyRWQq9wLQkOtRrhoG4bqUw3d5I6t+rQfbgBfrWhLU
hS7n7GSkUXoe44RTj08IFnvnmIiMtku2xpFaNX5fjLoSSE6YJO7PKz8gTJxADx21
gC1IwbwodsntwRqnOpqBLpwFStIUDNZue69byrcGws6csWYR4V8uhTuV3k2QAltv
R3XP7gSuOiEHUMngmIWrEP3RLZJelbq2Qd1TrTj351aT62RGj3Cd/RgVQ27UPM2E
mz0ahQvZoTL7Ii/qspIWjwfO1jx0wd/5ysWL+7DYuBdswF6vFoPoytL52hS0bntx
M8Jm1F2ZI7BnlDSkK8h+gZsg1xja7GDe6u4iOyBE7oZei694aGoXvAPaAR+Jyrqn
GC8LjxDDiWb+mHZQUmfVzgKU8aBJJprPhR+5IOYyEsf8gw8doqMRNZ8ZAcq40DKN
ZoaO0zyUUdUiZ9b/OuKKvsBM825ZYV0NpVUReSV3KZdVt30hwZcybQupDIFtXLQb
oUCQTngBMJefyXIw5tkAxx4zav66ZKsVgzCsZqV72Yd/XbA4WBJWbwDqgdLK8t5h
gcYdu7bHR3Uln322K0vLmGYbPlC4zxA8gxmXLI+6OvqBgg0LgdxsK+kmbj0/sT73
fE+IubqJBfj9VncNIn7Q2Zt5YvU7Oz7soVmlL//QQn9XCGTZu2dcx6CtGVY9ZP11
gpg45LwI6jRsfhuJexNj+fWat43DjImvCEFsrwobbZesseJ66wa7HDorIUYTa6pB
zDR3edIpki8oqXo1h3UJahRudhMqrLiE0G0JI5EnMZDt6NO8jknh1qun1L7EAgwe
ROsUs8B0pJVkswieqNGZ2pOXvxX2/uomNi5YY9WryizQu2dv9uaLzU+NxKrk5lMG
aVVD6FVKuUiZ91hp321YqK6mvDOTLfBffcidumcnyDFnZjRzM460MlPMtZhkPv+t
uZ0+/D6ac2QhnwmetUBYRAMXVRQuWxoGiRC1dS3EWtfM091m4GuSY+kF3CsNeBsL
YLrVuStH3OaJ2MsM0z/WsvD70VTBpkVjQlt7MckvG69ncUpGEZzj8thC8xiuZH8l
xumWf1vmdNNDfY6wVuzjy+PKVokqNiW3bjsv0f3ER/9m0GuX4dIq/HE5z2WakBhB
16V7HuykGfo/IzanNnTcpCgqvnijwnqKgATjk9Sn5lkRGNYCzpEGtN24q3RGgTeP
wbjW3rNJOF1unMD2AnaZ6JHP+CliKIN9VH+GebijNDbOsNMOJGIAzst5FgcAe+3l
WkwdkofwCLgIKPE06CnqZNoXt4B5N1vF+ErKFm/D0jAtyLazDlM0pTcFJUaG9ASh
ZzbBQtW/grs97ZVOjcilf91ZTCwH2hhgVAichXEWu+874SK+Ryw+jNSG+NuFXvjz
juZU8N2/AkxM9nwN5p8FpZZqDu1H8iHKQwjKs/kTds69X8UrClx62eqddZqxCPyT
fiX12xEtcCcpC0CDCOiu5oGXyK0QguPvWWR+tR1PNzxz7WcngXvfqH1ahA7LDVL3
ipurvQuyvk/XEisVnpZQlr+YFXvZcSWPwagv6M5uMljf8TSRjlgMGFYmWfnlSF7t
M+0LvCKtqDIR56IDw9QClVVR3udYzYv5ts4Bw0pp/+RCnUgpDqP6IDJl1SDgWzK+
4p6IBv0Q8yT4li8tqOoJgnSlujIyAW+HxVIqYoxnhdFIL2NgXdc1SznPVyJJKxKE
IVXovKso7USmFsKBCbAP4HSh2CzhOUFTFYPO1ZuDZpLtwXVjEPOPiw+Zy6nJZ7vY
ymaoDSNOHebsdnPalqp3kB1/K3HseDMeOFEO5R7ttCmvVBpbRflHAqWSFXPc1GT6
/cQdQJmRbitdWxPzaXUhhUzOjeVWdlFqQZoXubjP8DImTGxSYuuDjXNIUYB7C76h
0ALeDBuNYRINwVuZzwjsHoLbdb9Qqgp8pbr72pMKCowCH0irzVFmE2clfvODevXu
6dgI851eUre01gREfqzkk+Izl+IKYg39Wl/OEqtrsUWCm35lS2ANH9dyBYc5Vpg0
aD34UiBhfhjFr/ZnNBW36zTrkmtY0WhXCoyYhO3XbSDUqyUIHUWo6CszR22Frwih
3SgO4uMi+5FZcftrjULbcKTmAIeNsDNqFAVFmhf4zc65E1CY8Vv3UONyLAJsFyqG
lgXU97Qh/6ADu3qRZ4imwbEMVBglKVDB45baCjjwtq8T7AykTQUu6n4sfBY0stam
G/qmWYOSbwJ7PdAgOGxPfMui/+BMWitJBFQamD2W9KysNXv2Ve30F3CpZrLjz91B
E2VUG6xKB/qlFqlVLUjug8KMmu+tpy11uU21u14xBSBQYndZFOE59cPy2k66WfJ4
1X6MjlUOG0T3wb4gNTtWtPNNb1uwIIfb1PDJbufHflfh+m/aPhlJhivczIexBvqR
jmAERyeaj+yjRmF+3OPxy/izyhN/9q8pOmk4/GoHZcgN/GZ9nuGCVc93uN24Yyhx
MGAc/OcY5bWzHKx4ys2ZTQJyICQfGEdK6RhJL/Wd3nMk7+uDbRm+eUxBTC2W3v4j
RDnEdqyRjhPBbtXFiJ15mg4nxsqgR1hH51S/ZXfgfR4PYosCQofkikTIk1Wm6y0O
eRsqx1880zHBUgi992rjQJFqSPlsbqRUA6EplA/06m9ezIiUffTDlt+eEhUdpXTM
f4j8vjYglvKvGDKN79qLSOchjhrcSAyFR3A0jELB47wSb0WNXioYlTH5ai2XTHrH
n43NlPZVdFg3dMEFllkJqqsJf5okFshEBlug7l3HIMO04P8j1OEYzhEEVOfzWbOE
D9pMPoq1szzsBOHhtqpH7u1dtC9GEiZy56Jzescl0AJy/JrpPsksKy7qU4wXZs0y
Xd7OI7hAimrCQ1wAKDT7Ux20WTGuJtXF8UGesUTMv5IXhlohbgVUDuRS9D6wls66
pkbzdcQf8k1tTWL3B67jXGGhXC+yzZyhppqpLvj6pvPABmGPQFR9V+Vczs+ZtNe9
/oy5a6eMkxgIHiUheZtCOf79ffZAdHir59jBbxJdxRYs9kvgIUlTnHZ96PPU2J+p
Co5sZsMH+/A7DEM1amYVFQmgfPpdrq6OWMfXj2xZxvnbafONv8pWF35bh8c9moVi
3OrM6fxW6Te0gureBn7QvE+B3eGos15hPoyl3IwMLt86pGAMNFfyQY8zIduaKg0z
2l1/V99LdzNMUuZ9JTJESuHZKUlHDhZaspK+yP4HBR3FGwTSbfYiR7wbTqWKZTFG
4I/rgB62bYjGJwn2C30RC+S/XCYDc6OgY+EiTuzChAytJmjPDf30dowE4WPJbZDp
o7slHB2xaR5bu63ez4Sg9Dv/onnsClrWrZ/1EaxxzJPAAFNjkwLncJvaI3WBG3k5
mCnGdwCX1T3+wVIrRhJtaeqFwacphg6jxaP3kfLFgVU6fiHkNntpJOylKME3PYon
9AaFKAzrvkU8ZYxXPEYIaDh5xDXp+G1pYx8+6p0qgduMzWPET608yDZBMfkl16hb
VZ13BwG5N2DrF896Wk0gXpTdyQH+aiNYbG1xzIVnt5Ug+E8wCnV609UMxvB+zhts
qHXUqmEB60hJ7eSlcxzz4OX0hQ+uwxC5rONGTDroIdwUyC72uLIL7v5J/h6QJokF
9a4pI+1KiKGI83BBTeVBG5+hJ8m6J9oQWYvEytF+VYsD+BFPWKwfTSHTcg3jTfla
LzWBSeiyUPl7k2Vz3XLYN6caWjYmt3PEoWkA3Gj985Q2x3mAeWxmGF2hvdigtpKS
axay37SNhwtuI2LgyHLg/ewVqqE3+vLFuwPJ9Um8pqgA/6svL1KiZCrnsll2yDY4
02sKFnZg4cBz9ItYmT3MuCEgWW4jxtZ4uMVS5oc8yky5vqJWyDFNvwhJVzPGNX9P
UHxtdbBuM9u6o/urPYjuD0P9sWl7YR/AZ7ypfSyvnvst5+KeRqTH3wH8aBFrqTPp
GjpdeH4h1Aw9hEot7t27lcGxAAOyhTnpkNtW/Ua/c7ShOD93f0Pa13OenbdFHlEV
OBN843GNSE9KIu7jqJNjgjOF4ucMt5bI3gOSC2cchavcobDcuuzffcja4FTIllmV
jgWUwbVxUNaGxGJuzJB3Yh+irch2UX6pXJ3SMD+UU+Wq3V6n8RuRWwqaWieGDqWT
awgGCf30SNTJtAbcUTUAY/oWBINcb4PXnhZpxcWn+3LM8zahtkqX0f2NBFKG8qJv
soPfrhACDOBC1NqWddUmKCAIf0PPfDd5E7YlZAy4oKLpY+LwxhPzt0S4u4bDJlak
6HsHlSng2xSqZSRkAg9B8NwMEJXksdp/Lawsi1NsbOrKA+T19DRioUS/6929x5Jt
xmo6PzE2VUH/H93/GiQIk1zncDAAmmsbZjBUu1dni3/B93nxtTlVvu92YTZ41wFT
CcP0x5IKaagfnfJP81bd+EEJ+cjca/C36qGd2eNGrfsGsyfBnynYnKEHz981fR46
nuN5NjaDruPLltpJcp5QZ7BJmCVRCWbdBJnQpPJz9l87Ks528cZDC83XmV1Ri8rL
K13rIpMd4eFyNzgmx6fxzSGO/SO0pMMehAQVD/AbzMi+EkRhpTeORzFCKFCeScIk
cMtlmLkj7joK+u+xXRlbBlnUqM//+OVeFIz4oghguWkHVa7PLIeDJE/aWO25d3c3
IOpS2M3RCKRGdXTGZv0XPL2Xs4hIK5LbZ7jp1aq/l/utsnRYZI6EMJYRmDV2IF0o
DfCeT9eVG6tsfHhhxIguB13BavrVkanErrIPcm2Ua8N5DTdf52P23PDDoGItH2kT
TljK2Yh2b2BtCzSigPzB5HGFq9fNIqEnlIZ2Webp/CbUtEAu4epA8E+uh5ufK3JC
6OKCXSJvGRyi0xTUezYJXffbYyWXKHcEHfxn6u5cJNhEmwphusATQpYtqAi2sCz0
UnLsj8Q3y3x3RV/xCc9S0hsJrRL66ojFsp14Z6NbI1wiTndLBXdbuuGCjLETYVsg
9SRaDQtt5WUNLqPso26OQzzFvXYWJWMZGJPelbFidVfWod8qv4EcYNSRc3Moa92R
s3pog67pZqTl4N2dn8nRN4BC+s72PA6tuJk67//z+YQRwERgiI2esKDQOiUbXmfS
m5DksNCpvy4GxAEo7a9zWL9GDAfMdznDZQYlkNdzndoiD2GDMIZh0R3oRliUWLdy
fxR0ebVTumj2xTRvVblBumdryTMW4kXiHOnUZjWqfi0q+z1mtgwiwQs8plAIuT42
P5cmOIj5cH3nqenf9V/uba3ZAZQpgmTsVjHCKam30HtQb5qGNS80LB2nAusAjmsr
MRpo4RwRewp8BFeibBem6A4FxBmAukpfJ3zlzbDQkMMDgGDuO1UqtrEvqkndn6mp
bh6k0F3MfhL7fXbTMdC+qL9QkPIFGDx8651KXdVrMNcr9cdFsiUB8+VCuXyU++nQ
LPY+hat9hNsykywSjB6zvocEJFiPIqIIhvaQ8Ih6aaSmb8FQw5CiQYigEptzQuMo
VqnlUCc4F2sI1hXY/JroQidCLFHr7QnhU6I78josorgZBNJubZTh/JNQTpNOnL7p
K8Z3x51OSg33pezZJjgb6BLUJ/qQv0yDp2qY3ofFQCPvWfBbpwRe5LypqetdX/rT
aEgO5cAOSGHRzAk8C8bQ95qPvjiXF2Fy5sKfiltjU2mepFgMVJXnRny0OOgdHUPH
0I+7U0N4OXEeVQ3FVmWLsesRwa1WFjfbeGyBMS0KbC6kOl3A83/enPNuWvd/mDY+
IXgLmwKur9jJoPAoGuUzpr00SxrKPxIIjVHnjPJ8R7i+KT0nbM/JchR4wk33Jmuz
l9tm/PF9Kw4/JYv3pjg4V6D8GmEkTaetMnMDqigx6ot6lcz60c3RE1/ONMzf6lkv
co8vMHBRDsfix58S/TRai0FJcVFw/cp+Q3qTOMhHQj5HLZRne7iRqnQApwt/dJfX
RaDTptxZgUspve0Co2zPphuxxzJjSbWU9EmR17i8u/syCX07+NAC8eDqWBWJpyrp
/E4jq5+Mcp4INhxgsx/tZAlYP1JLqEHdsKOdZqoG7Et08wrq4ZQYHYMiAuVmoJkO
ELYso0nkg8/LJ8CcTxFQNASoJfpqNjGnGqAUvjbHqEXlukVpFq5FTuDaFqvUM7Fb
RM6xwGH87zrAj8GQq9nI4/as+9tHx/jTULfTKKPEwfMwBSlXZ7VYg77Vh3XvgU3R
mkixI012UP9Q+IHfs8J+wpf2KQJ8pSF6ZoSe3UxxbP53Vun9t6rbRWqh9FHxMgZe
eKSnwPnG+XoCLi+B7J5VA7NtdQkNtDk5RewvfeIfcUtkbOu0AoQmtl8ysmzT/e5z
QseY6cviV4YAxFM2ncpJS9zD0zWYCYU6tTQMzo5igVnDlNczWOEaZfIqyN6M4sCf
t1kB/5pugDouSok6Q6xjy5nasCnGhYgGP6WnQvb6kbzC54XjE9O2jP0KTkmPZh6x
SqSTtkJ0PBJvetcKjYQXvzzWCeR30cg1/sxH1EsbkjcO5CXeIBPfMwMIvYlX1nEl
q8a/ATQRl4RHkvesJnGbzPT8BjjDuJm7+Ndunnm3huOeo23ta2K7imwpOX/pMA3u
x7Donbg2IS51M7Yodt5kxgaB9jfM/fFTxXDWVq6ZE+aEM8FWFvC8trREJ5amz6I3
/LRr/AZprnLkOQwrtZinHlHwNbt7szuzzHl9UaDoKtrlk9AqmbPpFXT9zaowncLl
nhjSA7fHuwoc0oJqwmvcbCN4D4gePXCaox2DQ0gnaPOkxIWJ7L+7qHmbewrjXlXM
zLuTz1LpqFZUPPc4qUS+g8BWBO/EQcXtOwnBEm+M91dFTOwfgpJGSDNtLfEDZgmV
tNEhOVsRqxBTpI9Hz6lAWuFmn8lFamF2yoEmYIRKz2isJclB50QFgX/fEOo8F4oe
KFy5ZRgopxcHxRKvt3tEKcekoykQ0bziCDxofxgaAcsRIkYwtIgGTCoXzNHGhrWa
lDH1OljYwekCEsxE+z0KBoK2Oq+z+wgatuQyaZMEaGlxLheG3CkXctNX7b66lOTw
N6K1txoWzvQX28ww+w/+pcS/+dH3mslgGKYATaZ8a6D71v3nYMdLUke6RtXNPhS3
qaJdNwXQOAVqFMSkFMI3C2IZ2rUQkS0y2a3TX6B16McO4H7XEqOEXIkkK3b1NP2J
VFoBi6AvYiV4dxLl540oHV6i8uQqySJGKwgbt3ZBJPykaQYwRTungDV3jugAkEq8
ilSB2kZLoUxSPFluV8pgYAkQk8sRjZO9zgwCDpjN5pbfT2/YqwlcPEUWUXbC8LpT
2xwmZ3j3Jrxy0679a/zEGvNavU0rd2FarS2k749Wa3OrWNgAybbIoumhS4nH+0DN
lkt1PkCX007bcZwhtEj9FtvevK1sjPJ012Oy8TmyruDBqhPbylhX/IUjbOcWHf3J
OfMIf5s/gsDcWOL9tvMqO4AM8DmsIfhb6fPlYU9YWMKMA5qC1bLPw3N2B0m/nbma
LafSm7lJlECWTPRMSduwIepvyM9GQiD46hx9vSXXCuq6jvUVbtD/k3XGJiT2Vu8+
TOXO3cNAuEtoLfiiaQeytYmObeIQtfsjBNUSXr2ZmhiO+77hoH7N4DS8uiF2e8fO
OWVDhFiokHi8wSBrEYi5u0HZgWPr+0UVfSCxdEti34BMz2wapGof1jdDWD0rAHCf
mk4nwDP0Ldi+1hE4seJgDsxGPzTTSyLO25ApnJWKxI5lRHv579cQMqTqEeIPGKoI
MCvrFb1vZ9ZgAidpCXG9RB89b4HDucbq2clqlnS9ro2hz7zgmkBGujP/06/yN7FA
utqLoaXzwMCfnh/saAmU+Bt4j1VAwTCglX+xdBk3ULqbFjxElKRlTYHydaKXwxkh
w2/4fAI732WKeJWyF9ivfqFxkmKk6jArC9qmoH09ixQEURnL3uRL+Hbync8fvnMw
coPavmERwnAGbUAKOudmXsQRQVGAO/y9w0/MGMxO/f3mzSgmFOil1R46P8Wbsdwu
LC0Qy1gZCeLwVyHTQx4zHJ/MCmikHz3cY3ZkkdC9T4HBJZQFXcFiGtxGwNu3L5YY
ksQy+Gjwi/jF5Co4JxbfP83/0uWAU0suf3iUdYG1ByZAoejPf0Ki0uo5qJn15MGH
NgT8i33YYsqkCpPtY6uhtcM1A9WlTpqsFnJrlKy5Pg3jjc9W3J94Nkry7EltBbkm
Kk1+l799ubhv8k7mQk78v9v2C3FbV9trTJ3mef0k4qVoanMGlHs6H/6U6jkZFtbz
gCDgI2IKyLzHHI2hEotP3+yzifKpMyH7xFGc300cjm0YojNn4BQMPLhtGIrRKKBo
lyXDvRxDfi5P36eiTFnhwJWPq5jsmHkQs95tj8ocZFfBtQnFv4OTsiOyEGuECTRA
8a2Q0hG1R0mk+giVJJsOb01/o6GOP0ey9KwYsVcaSPqKZeL5L3ICsBgiWHTz3eUL
0RDw46g9uh6uutpe2QNRUIvDfsAhxAKPr5H5EQN/AIMy5eBnqmJe57Mgp+LDpDjk
8vPKfCg3vNBF2bxCY41jsaKIkhvWorjTBzDgQUxbdlA5dNddFXfp6BWOSEzvprZj
pUyZskb4dWGQFh47Tc4Sw6rmQsdjUDz9+aghTFWt3GdY5UhUMu00/MPxAXkgGsok
WR6bDLqACViQC1LT2oUBoLSx1JV0w6GjFu1qgIIhxtfn85wpamK9KD7sTG1txYFe
bfgJcZHSMkUBhu30URnR3aJ1xdnV2aNhtEpHU8J+3fENgDpF+1HWybiVk/D4YoKl
4Fb5t+FULLHFWTtzBhWNDwJyNk17QDVGnfvIJVwF/sne1fgDKKgKnSWkl6QSVB7s
IA+rO/xyym5PX2dQsBEqALKrPF07tmzWW3yMxQwf+sTXXh1alDdI9szuYjVqMaY0
aoO22b4dNAjPTsyp21YIYgxe5dCORZePdl5/kHOqD2VS3ny88wzAAxwa8M1X3ioz
V9k5u2AXhyPPcZXqnFQgAifgE1iuVe2u833YC9CZLRgfPgZJWpdYb08Vc9ghfRo+
eHosH2m4jASlTYbziAyATeOy7LJJ/AA2/JghSN8FMHqMAcunO3i7SSaOGjqrlFfz
zhVBSvmOJIFZVU+Y6THYawK//fI/YJPLYj4US2qZtkD/JPqgkSpwJDINu4hcm1vp
8HZaK2Mwq/emJrgj9yqk/XZACwt9VDHvfderD/shfS9I+AjxPZN1/vZjUTLurE7+
+B+AyYa8s+fCZHi7sESkxhzaj1bMlFTAMq5H2t9zWZyjVosmAfzSnMSaDG9Vhlq0
hffpzDpv//FJBMqUl57bh2vgpvc7ZGl0CC49rZ+qePMPln9wFshuOfmxgwPzDiiH
Om7gs1NeaPV1K8FtkIriwEJFY90ygpzRgPGJ3doTttYB1wh43wEhhtQC2ScWzOpT
8f8O4/vlwM+lJCmBr2Z8QBXiAqy54a1rPfQqOaJzll1/MzOvcUZDrJ5SO7HenY7c
alQ1GWkrK1shjV4bRkDhH8xgWGZkLTS9c6h6bRdekG1jk26ta4Qsb1a7DIoYGbO0
A3aa2alMxy1ChZ7VKtCq2FemONpSJ3y4kCup7XDgnDbDLtZ6aUJIaEMQZYYi6auQ
yYzysoHLwSqly3Y/7lNLkueN3JAsEfnmTYw0L2KkIN75EXj72bFWSNqm5I52w5C/
L2tIRgXF4/QPtxBwZQHiWAdnQZFkkBaOpS+T25OEJNTF9gooQwcafRl3wsRI4ADy
k6YSEOM3PVTjz+7AEhtMSfmeJWuJFlUcFEJnkx0FaLJElxXv06exp0V9IDF/Lq6g
nYhp/vWJnpCDuIEd2cjzKaupPY3smMmoROJZyE8pGoa3wFV2x4y5+vOZMc7iFFPL
G6kWwJmrAmUtjt5u7ha15XkFKVszkAaez8XY3regNz80DVnORjnZDfU+Y/+EWXTP
DaHQ7ZXjT44KlvXW2sO0P5r3jSwjJH1EpPRAOLvMzKSBFnhE5iiXQG+Qn+3genyX
+69KLXqJIT7HJJ4igKZ3q+y2p5x5XusrLt01S8wHwUM21+QP+WhDboz4WFA79RyA
qAzgGSTpVXGAJ+P2VBi11Sx4V6BGGIt3kbV8V+7FvkuV8uuThX5f52ta5toU6sQg
KG9OvevyMN+Q+ti635BZj2n6NXBf2VaktglGY2juChXO96qZ1AyW6oMV1v8XCLHc
IdRk09hXwztDKsZsE8vIuhsdrk9rtXFvRBb0AGuAcl6LgrRadWoQS+Bc03ldmR6K
Ez/buXpAVLPcuX2wDEewmzkSgivR1S69v059luKMiDvKEIZwgxylLFDxZl+7rVhT
ABi0Kl3sjcHtIKoV6ujXKmmhLLJynOJR0kx6q1Z1t+GB3tDIyWL39DIgdbwUUAN9
HilE4v2GoFx0X8Qf/6kRaejP4kmorwAUAMTnEN3kqIdtqxHV1z2eEoDaHuEviSyQ
27A8dH3rp8nXSDaQq4mxfZY3uGtPM8wiFEz5jKHkpBRhSZei0RmdmGe0c68rBct6
ogIU3hauZD6Z4Eoue+JhvRAjO5CL8gOkx4hde4nexqY753E2NUaQOaiX1T0gs/gQ
MD0K3PB5jW9ZwtnOQguwucmpRNCsTaZk4mXODWBDbBxZX/QJt9Bpg89vop069Gyz
LZDxMqHhJ5rmM7vEGHk27rlfheYe1NtPraShmyS6oTuU0snkh7HeE1awIvvMFX2/
eNsfbiCMk+bE/0Z2KD4pYQ3M+7+kn5HztXKinG9K/18F0CU+u2Ye+QUSq70dkG0c
QkbMrSoJoxL3adNosGR5VU/K77IQwG5cPyI8AkhYolc4//0qMaZM5nCsd10aGkL3
fd6ZokyA/iEtYzhcFR8/BLyWiZA8KpraPzq+zJCq8f/gvCCKbmNbx+V9T9BWx1Fa
HmbTA1ByirFb/K18h1aLm1xm9Kb/eE9YPRSW8ZDLb+ueihErtCEh7SVvflIYkajz
JBVoAREIN+5EH5yu+OmIBLBK/DpFh8y2TC+1g9WpfiNWyCy/Mjk2+YSEq7Ic7MQu
ifXsNHK9toA2WLS3k57q53XVmZQ05Brz8dhAYUt9dL4e92ofOJ5nHE7nxvihReEQ
jJP9cJB6S8To+0d8PLedXVFxolzbFuaizayleJTGl7/mXS+KkOA8j32CrrEtT4P4
xbQ/lzW27RCya7x+vKEvoJWKoGWinfIQY2wovwH9gMzdVyNVr4siy7B1+usEAUTE
T9Pp49GLR5wq5lVMXlrwVOO8MszKz9ybRVknBcaFF4/qhaPxH7OgS2XAgo0xjBpP
O9PbWeIyHXBa4yO6FC5Mesg9crBf/l0sMemzIde5Cx6GB32qgyIojLuVAj8yg2Kr
Jf7/NsQQDMYDvem4H+h/+T7+rNueY4Ja+PDysrdMqV5aRJV1vPUK5qtwrnM8HqEX
B4zr+Kwjx23VKvTv3wvvK6P03VixZwg8FlNwEvKYaZdWN8+1YAe1SRcAZBOnEH4n
205XuUDRvUJAys+J1w1Ci+WXOwUOyn4Ieer7kjBEIZ11QIocMazu/OTPGB4ubIyc
a3AUyzfYvax0cA3FOJ/lCis/5oCCxQOX7ythshlzIAhzGvD6qeqB/BxJOkIdZI6o
4jPL7hOg+FOtQ3qNmbRbyOjELsYhyxHrwSFBiK7sBKaQ+4XqPSproeLQwXBxz1on
tiF805gZCGWgSGQl3SkzamZMouPMNIUmeDE1axBR5wl3qoy8PQBLLmBjQJTqwq5q
H0XM+oITz/zNO9ZiqWzgBVNGsCfgjiqt/VoOvxuWtoIu83Tr2bX4gMKDKk0CUqDz
0XICqPmoaDMw9434/D04W3BQgdLsN1VsQsNOtbjXDB9jfZsN4xvVYLun5AVNxihb
o0uNbmwnFUZeUIi7oOmT6RB3ChghoN5H7SLu6VNIgivu5uFxTrTj5Va3vEdUQDRa
ikH4uuPlwpGaHyYEdg0ErZSgvn/IbEqrGp/+m3eB+fxTv0sSTn8uNuKVk1QSHvyo
jD+dthKyLwp6IsjWtTc7408x4QooqIVinNH4vfEjRTZ1eK/AooRipTy8OZDHsarM
1P9axAnQ+u5dUQY6AMtLlnB3McpQD76LALdbUXiXeKYydCdZenmxT3MGfuuDrabC
dtRkH7/sPRCCjlPxTaeoRE/Zp7gC36k2j19IZYcw5yKFO1MjsyrmZypnV7M47Ni4
MkKRJl/yG0aCftTtpnxBDxZBcuFJfGjT6VVVPoEeoXil+KMDqw97JUNmU+5syqjk
StHPwJ9kBPl0ja3NtNKpi9MLfX3kHvzmr1FQQF/ZTiaIaH3Sis7AJaXlCsBKhha3
lU3TSOPmuJ8KaiGOBvwBnxnpqMUXgf+v0zPG8I068XQKY/uAghv8ORooKVHTqAOt
T9gHUqjCbys4eBSId1/GjwZDlFD9wvRyR0Df6uF7jd6HGEZpsiaOGTyTaBs2mfPh
KzTPtbom4AMMaa0DJ0pRavfshtHHlhFl97rEZ6T4Zja8FJfD7I1G/et7ev2kPtC2
ow+/O2idfhEv2qdXEdJpKSWcT+3iPwpJfXfAMVtULybNT2W7Ls72mJib4wnNhKST
nx9ve7jVyFeJrcy39YPhMJLcI83utn286A5fVw8RIbk5/q6RFWiFf/5EW2gLPhjF
2+qm01nUGb8jfTBZKU3bAyjwyqgkuMeCTxq2PvaVn3iY74sg0WJWMEi1V86TS+uh
nNohGH54rdtnNa1tO99/LLtf0VyCHcOziOR2gg4wa88an62G+j55qBYFbcwrJ+xP
pDQPpmW6ZsaybhgvgocN6062K9wrFLoUPvaRruz50lHCtZh1H7sZzFkNmvoDCtrV
DXIHVs4/qW1cVT4s7hH23NfjOvGYJ6EAtTS/v3lQl4pxU47A4q2HBPdtUWHsKeAa
1lLLW1MD2LYmy//87YrBBVQ6j3Ohvu9sTyEXAIrETjzp0mctrWXSSUd75HS2JSkD
Zq2xE/9s8nGn/OxXKjZfSrLl6N5qfSMuaFcvDYCfdrkKL4+6ByGAy5pwtZaAYkqj
en42/rU4YgS+bYvC5GlrMQ57IPC7BmwO5Tim7XM29Ubs+mSfQs+bgP8ll2CzCRix
qfP3FFt6g+NQlA5SFQavTIZdms1aLDIcvdTYihPzCjOmsalxpVxTl8Wyl5Rxmb/3
+6KZi7qiSozeXqEO1nxHTbsGfX8XO9BDe34bqcgBFWNSy4kICrsiAKKC7t/rIbW9
7wjd7B2DlJGDJMAH7n4VZwSm/N7E8mrE144QIvBOB+XpS98P7UhFGIpIsFwZmPKD
YNmzQFKx/mU/P97c9/4fxKLH+a5FTeDa1BUIhg3t06ZxnA2zw9/uwIpGqxCH96j8
rw/3bauwq0o0+Qz2QN37S1alBE5NzGhMxrCFZ0d3+2acy7Vy728mfkjtg6qMd11r
5LV/ZGwsE0mj0ofbpIITYs6FtFSxX3EixeQlwzMMpFsddeKUEKYNe5z/ZkcMRjWD
yNYd5TF+U/4DvHaL7Fif4omMd6d1qXDgobAMohRRvymJxKmmWrvI+396DhniMD5p
USexDNhlUzhI4Lktqd2QSvZw9Alhfjbrh091cKsxnlIVtB/wgbunxsy4UQv+Fg1x
Ofj7aTF/eZBdUimRC/FZF+kcO/CyMODffOrb6pkqsrjN8kLcUc7l+K7TD1K+DzN7
oBoAcZgW5Y/NpkYyoceDsTx9mf0Ot5SofKDWFUIGnRA72uWg1K2x5/HCUbSdK7jR
moUgo58Hl9n6UMepBCmJGYJh4UEVD/ArJ22EKBB7wxmUldwvI8IEHyOMj8rmyDC/
JN2MQiPLLykiUDk5XfKAYzbxKJp6tTA0OMFjzT5kr3Kq5tACGu/EVitAWPKwrpLP
uPBukzmRoVdc6CO/eRDIMqsMRl2C3qImwpDzOgV9QyBnZfPWxsW5vlOkOx7mG3N/
AZ8kHiHdwb2rMEfUQnvJ8Y6NTFMaloEu6/bogx7SEfSrQyFJFxppog7kp1N7d8fi
g+Lul0rOF6mdkVMp9DNpgMTYqwXuRNOJKzCeDOiVmfUqPpvXD1vVkv+SQVBJ0V3l
R80BgVMBpIQrCdbku6LMYO5pcs63a+mBwhLb2gF+vD0qyhbI0eAwxQGhOe7JQ3b/
g3kf0GjfJoTlAoV7pKBOhUFED+zAFMaMOVvWa/YBtyjR2zr+/uY0A+r+uogvx0Wz
9XV0Eaptevl/CWimB3rnS3/jWwMhXg5tXkF2/oXBJTeUhoyie7fFiTX9ir3l7Qyh
66uPXk+Fiqt4A2Tzw9HmFvCi7R/IOHZ0AnPNw0WrcQzoBVBKnjETETR+wo/q3Dny
zqPL6dqagw2TheX7IH4IR5TSU/EkyMf4VSmI+bhOba4ADqfu6M5zI+d4snaxlxji
iFQD1zGQQXMtZcrr/IUXavAVLjPmMtXClHWjYX2CDazUBcN7RoCyTOUfdGgIEgkO
w5+G1UlJuSTk5JNKo+yX8DH1IbirEV1KBWLqn+fsfCKHbQ0k2N7RkqoguYAGMA1H
ZwnoUd75D0VI3VLVEaqX0OU+PwqUbXM2tRrkcYpXl1akS58hVJ1/MFSqdhcC1moc
8qQ+NpDbxA+q8QewBIQ9gw0P7jRVF44v5o3y/XyjQ9YeIY1WmLuomtafhOic+6sI
Tfi7cOQVxSUGqMZsm/qTNdV4rYGa6d6WP22mgLOovYSU//fpuSSC492rH8So31Ig
n8Q/n019jTflhU3p7rKvrgWyjllGZZZRhUrRCPQbg5qJnX0780ZrN9cBhpL6wfPZ
NdjglFz4Vr0AEZzmypbhTwSaF/AebNyFZuOz0DN09FD6Eh7b8Vset1V4rEIkPa50
6F1fIJEJsD+BxVYpHNlvXHepwZCfAUt1u3rOPJoCSzOGqk37XJekvl3i+Y6OSVjY
/GlrPpA6EROmJtXIcLzf9KOWEZhrEfKVVlof54NB1QZ+cSvwRvS2hGweaK/4t927
WnLtws5d1Yfk10s4VHiaMOxbhJlFimlIpWR0h3rs2AudyG8DBLMccy62lnQG0O4y
3EJ4gxbS5Tua9EZxTHUw3AMRA7Cfj/GdjqqBC8tkZUhNmdOo1rrICwzp6mNcGPGD
WqC6WZYPM0M/v/sUFmKnKJLCryQV5J9SRrWHzGJT7tgzbeCBh5hHwsuzzP0kEw6u
hjw12ieeXxtgduDIHEhOH09+qlX5NLg1FcGjVGPu2rKUsJElkgZM/SfU9phxGv2z
1Bj4c35qPY7MGGGMg9PZC0xmdNe9BCgqiFF1MuX4CeHv3U/Q/EaFC7snA910OKeq
LsazI3yWJMuH68E1vEi7hl4ghZZ0g5VfcQM2MSFeo+KiUenls8QAy1A2+POBJ/xQ
VgC09zvSu2E5Esn6Dn/zDK+tbjC3hcZCRFtLjMyDof1foKKIiE4xXTXFJeMFul1j
TgrMbx9Nte/MrMo3fmPGJUvlT0e29ZY3Y3gHBst2K6vQHx0Dlhy1vIjqP42OKOZy
XFg7YqfpLaVF13KPtW8CY7WTZx6zUdHh6ExL2V86DoVl1Fc7JPZRwotp2RR7CagA
s2Aq6UsjmDZgdP3gADmqXuOS3yYjSwDwZ0Lop5aYY4mDVuY3OyyhycrcalT5Z/W9
So3+GLXLh11smz+D0EsQFpEkdUai0yy3MMxTSS00R4J9Db4s438x3aJsscp56t2L
yI5paPQuPEAsKjc8c3fqycHMe0kX1nos0RDohwC+u0tO20uby5Xdl5a2XeX9BrLx
U9MaEvCXOBi1vhJzXKuW9tO2eF7+vPPtRaz/iQah2/wvtclAsR0Kv0l7lO/QeXcl
Q7wMlSP9h3ldRcX6SruSrKbwBj69QZQv9Y0MPJPJHYtULBTLz7DDx1zCJuF5z0c5
cLKydpUUrax8Hwu5SrI5P4t1bCp+DAtjkrBTaF0USJcx1+tgVXdnfsPUkwLxFsel
Rwcqb940UzmPQZ25EGk1X21r0NgW8Y+wHaLwiZuU8c7LZuKxMo1QsjlcCENHDwql
7GH8Zjq0juUxMbQV2Of3uTK2LVc4sKoqKSnrePzM4JtgUJaU4PEgEZk52iU/zlxT
QCk32BpSF7TC/6xnfzb6fkIWjE4hlX5Z1tEAFuyeeA1Syo/U5zJzSd+8noryXggk
Had4cDKqYCILpqkk58d00qRYE3HtvHRBJYdqtspNqcOlVwmQBCC8h35PJHGAKC/z
874NopLEFpwmJ8bY96zjDg1bl9U49HoSi8QaopPrZ96QPQC4oPpUdlPNwdcKqL52
SkytJC4EPUSlTkK59XDgwuvd/2qdJgTFi6ex1I1quJGDGBu+9KfUd7DXP4T18fQ2
cukoDkTqeTjaLgWtFgova8dvW7m/ey/Sx/J2Hu/uj1or8FGB9yJDcVTkNF5D/JhZ
o2IsxeBAkuvNpYFEAbqzdRhVReDkdxdbdQy+jntT9qTU7TlKXjisL/Al7Z6QwcJu
oyJ9THevd43xsgPBjyEuY/462EhkGcOAmIDCCDjO9SixjoqpmjIPJ54TmpJCksaK
5dlZG3msJh6AZG83gunrrOTr6txSZ2WU/cyZU7WzseUQZ9L21x/wxF5dxktMnzWk
ABXlz6NXFHEjJHfAOcDk+qPkm3Vh58FZB2IYZhwpu0xT31E5dpZrH+nnowxVwz0r
X2ZD6Tn9U9lrILLG9VwZhdbDV/UphZgjq4G/HIEEWJm1VFJVGI4EfeIjJiIrLk5K
J1e/o5kViBLpWtd2sOShEH5oOWyDbk0fwELu8lGfLdHSfpI9WyyrtQ886aEtTMA6
ieWUqu7MrCgqbFjJudumEVx3a0/uT/xszbbKj9kB/RS6q5M5LsWrKslIDL2ENfWO
Qb/oejtoopEg4izjasVHITRASPa5z2pcAIGeWYvnngUYwhs5TmmmU2MD4GOKkJAy
Q9Di1QHOg62Itjd6cXoTXRWSnDKVvJXKYyYcYsX3hHXMSDp/VbyGTMUMHMfsb7IO
UwLr5OvCnUFLkeaTe6uOcv2UY/IY5nsgIm3CeBBKo/6FwRSHWxSwSbgmp6dIPucZ
+wkOUOW/7WJ8Nbe7J60KrTH8/XUOB8eW30TV12uFfI/6oLRkF023oADpWw2KQEFk
xtSIq+JDJn0DtC6URN/RIm3ZoZPsdsVohbI0iA1xg+P3a7+OKzPR9gctsdnjep8p
mmY68TYHMXvmVGy7XyBCGQI9A+kNlPu69Xzx0a+Vk4IsoF2iFrYx7T7++WuYOeaO
uVJuQqd4Ivy1nu/jopzdjyOwWc+3yEAnrPMvqRozUwhsAWNmf0fk9sZWPXhAkHFp
V1iLC0OJ/xaCTiMCQdeVggJTRZRnOsEH2rZqH7PdMPS/u4mMgrVSUmP4Hoji6zLB
kIzxec1qNj2kO0GbW0EcHGGe0BeukQSpcsFDed8qZj79ilcQ+l7jZLBAZvh9qX/k
zXW3c8dLwOHPtkdQLVTNkITKWamA36RNf2Wj/ZQIp0XmruA7BZJM47DRGT6lx9rb
lI4TRGhz7LwlG5XWsr0+qf2fG/PvHliI3EexepN5ddzuUgQoxbV9FdsHWQpXm/W0
IG9Uho1bI9rBFqFJWbcsIy79inWjgY5s4HhND9CU0KGjhLp/ZK+tyXl71MNrLdo3
Ka7WkR4UzXox5hJATV/4LjofIberx/AXt7c7PMgjOtzGQ6II2tBtaYtFGDlRnexi
8lgCw7/R+cdwCQonRrzMKhWV19NcMKeCWSCEPPjQc7CtYtqVD+mXMmwai7Z+aW0I
UwcZqrymIgCURV4lFmWDca8smj7yVCA3peNC6+U8m8u8ZtzDDZa4AQX6CAWJsyBD
Mx7QTJYiV+LBvvQop2Y9y2NCE83MY38mV7VROGHB0qy2w2VdUz9FsxmGU8Gc36JX
LYFyxQXRZlgMHh88f09DEHZ2T1SlXsCE9dmw6hVWIhlUvlVscds8td48pB6V6f4J
MJnDpB6rtIww1Cvv/qYi2mdHjif3CBMMr01NPCPyeGMjuc1/YInh5Oe1zD2x+tgp
UDOjtyBHCUeZ/26EFKT8JOp4T2jqFuaw+XwsaN5AaKUmKoj3Egel0rChujuULLuU
9qtzP3MvnK9/d066tFO4ttyMTh5F0yqOG3CDYDzUTu5CjIaXHPahWHY0Gfv0uKZD
XM0xb+tqSuRpV7SC1UDiG2loISmsdloSV1uMys0a2qPSD04JfeMXEdF+hjw+iQ8R
sASfBGgB8wAZtqbNm40vW5CvZCQUrbWOLK/5igsFb5Gbb5xiG1AZZmGTYpRPciIV
FMZxzBQimZY4KX8wWCfM6/l1DdRqFS2c0wN+uX32xVvYwy0FRzhIaApGTBOWZhFM
wAMgPcAaixMcuDLtAE3s1T62X966bXXjrvJYG+vm7/zFpfQ1gjG8LkD7xzEh2qyt
ZIA+oBSeyvS/mMw+CaSeRA8snOCrUXnN8J82YgNAu2Tc165IH8e8ED/XWsaGKszk
keMi0eHlQ4I/+Oj7+Y8dnjAULe5W0sHPVJbXo/1yXTgrMuQlXVAzp43VDyBEMo8q
rbhWIR1fRFWSO9QjL4z3zbsnGynSsk3yK9Z0yOSGqERjnxrY2jOr5DVsunaR4QwK
dkTuLaWvQJum4z4oq3ZtbuNnXPKx5VtBUdFG6LGywevD2kYo45kn5OaWWNuATnrd
Xn26hatqzHFh75bTRzOhakiJQ/jAXGlkrEvPwISFwl1/OuCX7tWABFLmHnn0aKL/
wnpx0t0q3aMbZQujNdWBoqKxSeAP1N2AdQ8NxFQiFpY791t6Gdo7OR49LNem/Aau
SLGvUITAz9+Oc3uux0iaTiHiEQzqxyj876rKAmIeM7tCBUw+vQBBlzNkzApwU/Sl
8TloPs1IGDDMEm3459bs6beY3C6/N31CgPIHr9kUvxAWO4kwpiU8xl6U8flVAJ7R
U0MIjSznp4V6J76dLRz5NGLBh2RH+OTuaiDAzGyG11c2kbSb+vyV1GcOKQBFQ/Gv
aWzo7+hcUhyCQrd2cH0I+4O8BGGH0+ZUznqutSZrrwwUX65Brx7zShWl8cai8/8P
XchHmVVuUbEgFP+HpQ385E9xonS0Akk0T5Yj+ZKrdz23Pf/jVw6pENlCEHDCLIw8
RINyKaA2Nm1JiwJUGZj/VRpOlTMZDdxoORNTWfIsfWfFa06hAYyFylWVVbXHgAQG
uvhkg4wMqW2ksTkvY8qUGQ1L90OjsdbI+0aW8Uw8jLszIpA2FHp3VMz7uMTeDrZt
2JosYXksd0gkMOT+6lx4g4RKtYc379FkCjhxaJCqBMUSdXalkikQAxbTW/9CeADb
K17gvSMW6Rj1pdGrD7xbYf8JWXC/zb2GLKeCjxRnxJ+x6kR1kGlGInOOwuheUr5h
GSYfW09XQMUrdFezDtMDnDbDlgzWQKIgc0dEkJV1BdU73sI7UYMP5DPVhjlDavIW
bw6AbQ/8NZtyqfuL2hu66REc0hNvLV3+Lp7LSgltDv1ZqUmEMQuYywmDmaTPwXgf
YxSRR+TEvqMtBslz5Mm19ab8mpel/DK1CfzzVF4BWWgHjPlryl5gXdoz2+FtF7wM
7LPOWUrbzioS6ZASJhipYdoymOaKklIM6K/HztM7mH79EAETK3cB6y95wKcDOODU
ClE+uTRQNhazYQf7RAsEVAXv7vHTXI+Q8xNS9DJOqCiHceNnvD+x1ysQphd8gho/
ScUXsqaJMtwhSoEE7sbAXd2AjDcZD0UXQ183VXmQdAptyosimNtdaNmKzji6HoGq
z/2fCDNQ2ST5Ut5REeO9KTyCZKcpFmaY/gCiJau1S3nGyn1IjioSjT7BcwFneICl
VYinnUTnYEKGShFmUgECUHaPKibaJI+NKTvREtuLxK/N2+DIqr5K+7DA7ENvUWJo
qEq67mQ4JcbbFlSCnZLlDiTDh08xw0sIYPFLDkMtYY6LEXqq7ssE3GmA0av04NTy
JRlMylABcRgd9PyErKcCrHukEX/70xrkwHljpGTi4mz4ppED3r4+1AP6cFvOQpcH
AFU8rE2rUrQiXsuKHuelfaRPXvgM0yrhQLICZ1ksCWazjRwZEymOCcxh//LX3Csq
2DjrvKO1echPKMBF5kdthyEvvAovfEbbIAa6GZ8MoiJB9NVmpOtn+R7PgRvtgVGm
7ZjxNu3Na93TjtJkyr7ZESJ7KehLpAu2mJmd5l+1WDHLbrdZOfRPtyByCIXBxwpI
12k9USpv0RUBG2FyhNnqwhHSOrMXmys2o5k0OGNa+NYb1840B6z+6rbKSHPlr5CO
rgzWyHzMmm2NcgcePLndcopgkP9TYkJjdURS2Ne4VECZun2CvKWs2AneeCCIn5CC
cYTrBHkBdyU3ZPfYlsnfk/gGY6tuUpvWytggmB1TkY0pT5zsgL1IzEpb7HCXvfgl
l0cDRjsV0maIKpb4RnTLMA9NsV/4VfR0c7hG1IMFZsSRMFPbHYg1hb9R2oj2Z5Wb
2b/ZrY1EQmaGzgjQ41PWj6LZ91+YzzBiQRkWHQQFhIhe7q4A//nGYTccgu0RNUhG
e7aVr6KaULt3pLDKa6evmkEuRifkn+488GKPcV+DNRCqJpGWl2/ATLnKOlhrfZAJ
ifWeN20kV2glCT6inC/nWg==
`pragma protect end_protected
