// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
p96KCfjA/2a5Ds4+PuORLlsKBVPApnhhmyhRACUGzk9DFvfoXl4iDY/V+VebsTvN
QebYmk3CFOTEctvcspzVcdLbOCN9ANKhfEZC4fUSWskmNCzkTkNrIl6/m0dcGKIu
yiZ+kN2B5A4w5cJL4W+4zR3B6CYf6/jKbECW/09mXd0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7568)
+RlYzBLfyxgb4zwSmjKjNsqvEimpUVY4Yk+DrHY/csjtM5EFxMEKeICrIPUyt6va
cldCC2Rl+f4U7l8C4Ex6BDsSnGrUn7vIUAeMGZtBKajmSBuwUuA1fDD6z/0hQhvO
hgI/Bp8IAlfiVmil+MPIia6m5TJXSvZL4fe0hKz8Nj4dqVGoTL7+5TfZ0Aclo2eo
rq+vEeOiwjIz+YaYAyLHXzRgJpXOpEoq2/Iye838uM/c5NFBt/gbPBiOcTUn/l54
TFtJtkk0ztR1seeAXRKP/12ibKmaYhpeI0KOOZ9uYKc68bVQmYuBx14tuWpI5Z6b
N7DhLi4M8r4zbi4bI4e5Y3mwcLkXjKyAn52fIil74D4XXt1DdIaCFlPj9a/rfIdb
jUx27rHKtSJ8jbGJntdP73XSccIAtdJIUHhGflyfwxOhqxT80zsJXTTnEOCzo9la
LQqIETJUHlDI8E3VWmMzvh+/fhb4pANiFiOzSPWbiZAXun0xSOTsMnruV4DDG7kg
ySn+GlnC/OhycRQyXaj/soJPsyM/8MX8sn692QBXnQRa9u1EtGWIjIDt+lPCWCjw
OOMvx4hCCqaM9ByJ6a5IY4mQy73KWY76ffdPRD42/gUcOq7RJlqSCFfs/Q4f899C
yL9zFzSTfFdJ1lyNZCy4wa96fWaoez4LrsxgTeJzbAt+41budXyqxJeKu4JlI69k
D3wX+SexE+NPeTp58gDp5v+0udJUMcnKsHjICJAwAAteZH4eM7PZtwogLDb/AYcQ
pUqrvBU85wQl+5uhx37qgjOiSNS2Nn2BqOBHQbw3S1oLHIyYcpXAb36wOMhj9u7A
aNAp9jnoM7lOvD5R+PeD5x9DZr7n9k1GEZmn2ANm8QSKOpwpOc2jp0dhk6oJFB6/
U6yh8urh0IHySFUPwygGz1yG/GqsKyg7Vx82btr1335maByOTuY7bouhrWA9+igT
uyUicopLKhsPFZdaWKETew6fDKkZSh45Gu/qrOBi0ZAbitqGXP6/JGLGf8iVk0yS
5Rq7etMYMB2rU36QqaFamlpNT7suDaLON4TTM0kxQD3+4johCEigISVurCEQcLOE
XxN6ETF0Ib+rkjVvQIG3ggq9YA7Z++2iOHO92eTPrUwotVm8XfDX4Qk0SJjfkHFR
YJW3BW+sNk1777VjEfmmFcbIW8NTq0NEswHfutEkVKhUQvGCmrJroHSpa2dhlb1S
RplLNdHwjIMZw0Tf9+c7Fstgb9C3eI7VsmSjrC9nJvuuVVo5//md5GD9/IB71HVL
dcoxsIAwYqIj9Mm+wEQupRkEhND3NSVfJBxvDWXxN+LF8UeGrXwY74IY8NRI2+np
R1WMAs4kzmy00DJHtAPatf0XiqBpVYHSye0pEi5d6ix613iCR01JwweTt/DHJ/RQ
LMo6QSTRI3NsQ7dBhZbOVXaa7M8awIrs6I3ZSs7d5aP0ZDQ9mPvoWsiYgTN5JVbD
/IjR9D5x7Gc7FE819m2q5+RY4yZXS6bMkG320uIeLiWgG80uQZTydpc6LRPZqert
URB4qPUhBzHznZ7CEXL7tUEqPmvPsJMcKllfI01PzVZ7yS+ZR2lSM5BkZjbktbOc
N0q/1KBKXPxxuUZ6nmbR6ZYH+ShVgQZQEuc/68lO3jYw3t2DhPHWSutGrGJpOOxd
UezP7rRv6VCNSsc/aLiefoswhK5VOXWJpZt3SOUiStzSIjUKSfbrovZesxxOhNkW
X4MjEyu+LLPivJV9q6LlgOTvPA5AFe691DvEoYViJIH1GlECh32BD+3YZ/Mv7p5d
IxeuIH7F2ueobbZNoKGpKpMVujB+k6+5V8YiYgPPXupJYdc9foZv2bqVg/ofQRxY
yuwjoLomiJiXnRRGo5F6i6OVtwjIUvHh4AKhdnUL6ImMTTBkNDAsGC5AF8XQTeJP
exnAHBkYEkbXE5+rcv+mBWi/9lJnBBQ6EtA4xunBIAycGHspsT586mSGEMwVTU0U
WO5b9V67/T9NN9zasRXbl3vlm+tNceA57lydVlukBGffT+jaXdPH11ylRb7Y1HZx
eS4Nu8ctXmgF/MX5ugAz4lMhWwRfXlesPIbNeX1eq4LOKeX6qCfvy3istU+QHQZg
DN1AQhNRo9kDyFoT/Gt2pAVIQojG8KGRL7wcPWhZuweF6ZtRmyD6A3pDbTiL/v2h
8xDz/LVpTOdZ1WqKcvSWhW4WgrF+5x55LpTshTQIIZfTmwHZ2QhEcR+jC8/nqjBu
Hdnk7Slu7Ytc+zLszg/wefrDy3rbzk53Oojwd2jI5mTYm0Di/cgTkvufRACR9IzO
v9NqiHvtE5+7PhAtWxRuNoaP9D6+P9sfbN2ju3Cpl/qiiaOH6VQuvJfQrLrPstzE
cit/zSA7CDuh6Y193x0uLSoNsYyD+epqAYJA30AXs1E8oXZnOMhd9/2d4rjE3WbF
dYsDgBpWA6g8rvKxtXsb+0YsDY4fcqQG6HuLqFfcPGGJAbjiWuk7PC6fX0WPAnNu
QIB/dE2UqJUKWunyVr2gjwgNzJ+TzlFr8fcX0tCLL7R5/tUl5ojOPLHY9A84KJja
gfZDss76fkGHSHjWKKuf9/u5qY5+ZhCTSP3g4c59Esb6vL9gmTM0DJub6sabSjrK
hfJyr09bHpGAXCzLkO+0csJsNeoFl2XRDIyp83+LOOlrnj1c6EBzFYdbVrFaEURG
sBL4yXgiKI2NRBccl1EuURheUXzov9LNvA2dDs9IhHsKlmDvj4nWZ7mOzFIxn8Ck
KdXQWA9CkJ6++xqeHYneVjpycZ7pOdM9MHdndBKTyU9kXuXtGcdKvptCKPbCCZzZ
vn/67ADswNS9KeFI19C5Bv5aroMFzUs6PcdRzFO6AT4u/u+YWCtfICQWLn+4ua1f
yJaytg+/1++3Ls61bRDxDnMxloLGzEvwHEL/6LbJGCdgu+bNhAHNMG26cH2Q1uq7
DsGaJQ9n0TTsUU6Us7XvhGqw7ZKl8tLbGUj+IEKOzt5T4Pqn/bpt7kr4SCs4wQyK
0xiXnbkqJ7TkZ4ZAUJksKNy9gnNc7j2iyuodE2+IGJ0cNaaTf+joW1jPzJlfn3dP
BPVBqmDKMh/9G5ZgkdtVvAUota9v8PU5rR3RizbOgZcdsxXr5iLsuDzegknCoCcG
0WcCKvVU8Xk1V97FGDtEs1LFhwYA+wvbE4ww2v2UU+jEH2V0q03VuukphT5TbQFg
H65vSwfe5Ek3ADP2ABvW6exKgImX4ueMAs+JB3ujuixaD+nINh3fRkLSxs7UWLuQ
z8N6VacYwrPOLnTggfAry7SsnWPKC4jGQ7IMHgNyXPTMxQlnJcoOgG+Z2G2bzNaY
ESUkp2iKHRBRyzGQzd7ZNnb1j4lucnVpUO37lYpKbVbZyXB7MX0k6PTEl5SFG9vC
23RnijtG+1phgnv41zEYZYXoH2/h0SSGlGra6Jb5cxNFs5I48en/CaCC7BjkmtOd
cWplWNUOwcV8UzEabS7uArE2c/hk8WGEtFkEBrh8hOLCbAyG5cFPKB8BCdkgw9yM
+x8nmNKmW9jrbZUsLXWP7h0uxA2cL8FN5l2Rbvhd0XFVCi1SJI4gpbhqkC32V4I+
/SbR0zvvyJheRw+dqAcqRbEUnP8ou1GnxcjAAsYu4/tsQArmFLBc3eYj8YrAH1su
MVhu9iCdcnSftsHrALjCUtJ+pK++fzqP52KnncjiwgtGO2eAx0BJmsPNpTD7W7wJ
oW1Verzf+b3Xun/fKZ8qQ1ZpqmqaudM7WDg4doZ5fnNa0WtBEU+ML1CIzWd0B447
5WfrhQaDgk5dIpEako4DcyPTw/oTDkfGtNUUtiTelT2E93iR2H7NxRkcMjJvx5Uf
HviU5kH4odJmnllraneCaRRm0FWfKotoytPLMxPmQTRp10JWMIWe1mBwLJNZB3n9
CWPwiuOlSn85X5cECcWaf/2oSXAWAGTnAc7cqwcxKi6y2321pKYYhC9bz+23gJ7b
wgMJHjzD153eaPjt+jpBgIBvjJ3NyW2gQYEX7It0rNzFOeCNDVqN/qjwNZHUUvTu
HFe/cSI8yAFGFGMPHG8ikDElOecxMq7ifHZ2nfiIkm0ZSaDsyHP0g+6w8cxC8xKu
iBiZmaVz9Uj7TLcQFvjrqVsCBQSyLXmMTCRCZ529DGE7pOwey3QBFtyKvWFk2jJ3
ROKUzAIPXycKzRc32QgX5HUPwfG2ifB9BGWNE+ggxmeoFJdHQ5OQFEgJiC46b5UM
my0H64TALeQ41oImx5IAhlWc+G9CQzP5dUI3g1I6prFus7ArWVG+9psLADf3ODrA
VqTfYyt0IamRACFb1U34khBEZJoc+R4gVuh3rw7raUhc0BRrljpi/n7N14ktRvVq
pa+cMO48/K4lPdny2dzFlZcpmAEsbIxUNQm2XFCmOUWKuIAmVmEqoqMVdZCU+KcJ
tYEjhN/cii/nU/ZWR1xhxGTa5lnn9EXABjRnl10hHLhRJrRP/4z2v3hfZ3r82iV7
/nV8Wxn9YTRNEwVTuKQ3rQzapkVB/hoG1V2zNepXQstodwS8sRQmQUID+yNrgmzT
CiiDYNf92zxGRS3bF4NgQ6xv9tIdiWS9SKuH+6pJeIH6Siso55xk02K6XCuSk+k1
bqZOjXzGj59/vL1UlC3mBF+ywru9+UHzjcpB0gUth75ryOmFolZvQ44n/ibwHzmz
RpARgZ0/iDOG9GTnaXI9/Ld94r/GUpy4Mq4iJjoDbwmRelFn5XkdComusP2p/Knk
4vBBh0FHIGggnAJoD4CtyvEktxt15sjkVjN+bwNvbaarGs0ycrUKlEI1kwjTU5fC
HlSgE3vCmQLGMcL+Wq0CrefFs8Jh9qfU7tl+d8sVd1X3eVR89bstKH+Hr9Fsu9vR
OSk7MOP6B2CQXZwJzM0rt7sBF4OhS+Mf3lENwSgiiMa5MhSDhj/FSdNFwZxTPKzI
oUTReHN6pYmpnRE15WfIVpRIYB3UDv/9P1risBl7qL/wSyChJYNeD2vNfJ/jX5Q5
ZzuvH3aBxCMNK8M3e2/G/NFyiybEHFqcyI+5funuy/MMlAoLiaVM2Jb7G+PYZ+PY
RcC5lisL3XV6peHNtm9EU7Jj4MqpaSCGvNGPQrs9MxPgfduu7227K533Y/aBX+qq
raKGSfzJ1ZZ1tAfrJDpi9z3KrAMyPquqS9ws98ct2LyzJkKf5pFDfjC+WJAPIaqB
C2dSG0EHBMy+yUxj9Fi+xioQU0H2sgyeXf+BeTIArf4vwWb6IY5XQA/tFd7aoEir
2UoSmwKRqzaafuPn02WZ8SoEqZ8SWpkT+T0IL3pdqMlOohSBGQEHqDdZVR4PoZvT
7wzFVBdlPpLJeuH/aUy1I7KreDuGM0CnIqb0GO7LSG8VXkki5UsHEHgpnx6XvMZh
iq2hxJaXfrBbbYcksn1j4kYyuKftnREF9EeWkr+FKb6BYHlWrzRlJ59MBWF4HdD1
0cnx/N3IYTrPz4M/Q2YDQPrpjyBEyQ7cz6U52Bxd6MmBkZhTtK1WpN96sH+vgNLy
wLA5mTJrykwPqC7eRiCpIi6dX+k33aDHmgBpqOx0nqqZLxxxVJCmt2AKefB7cxHJ
IBqiolAP88uM2O/FaLPcs1tgFypCqaJwCCNXK1vog/1PBWbwEBa6VpGSLXC8wdvS
JM9nYra7EPBrNvxXvEN1Rcps12v02NjcB27JTuDGn4S1TIErhScdfvoaHYrSonJW
ihgonjBHbs3CXB7VrLlGX6bn9rHygJ7OgqOND3KjmhFs2v/BG/A8xnMiqp3lwlpl
f7UxIuoTydsatyXPnNfssqGPeBnzirly8vDnvHhkJezQVfJvvpuSLU4ecqWwp5DY
jMBXO17cCG9FIedoJoU4yKWQXlZXPGq3OzsIyhvHRJAZETdidBo2ev2wzhlNn6np
GC0FgL8euUul/+9ktM6q8aAIlgMeU97hWDou90wC8Qn/XjuEwcXZ4qsG7eQNkcEy
h/dwgvTXG8Jh5X/rdfqy/OL9FqQPjOKzCoeRlSu5OicYYj2QAaZZ7ECi8+1CNpNI
T8/UB2XXmRpxg9n2dZKs5kcYOO3IC6r7hc6RsYKUAieJ3umSZgSVnz5nkF1kPz9F
aqKQNWrkgVEPKqJCzDOzjB0b77W48ugceBbvIWJWZjl5591GIgnD+T2rF1NlgYBb
1TPdKJZnjSCWdI1/XhA0UpaZeEyTrmPU/nAbVvWA+bEt9FIod7Mq7XWIUrmqzEwJ
gjyduS157g+eJ9iJfbWit1pG+ikJvDcsF5tMda5EteY0BkMioXxhP5bWudW5xrEP
xjKilZBrq27lwVVIp7mnM3vs8QCtjL+qEe6sblFCQaGj6mhPoG/zlw65ktjWz+vk
SGetlsDE/t3TiLzQdRWs/Cm1Bpmz/QHaYQ9u0P5xDKeG7rteVV1RJEPbvw9DEiJf
OcPZHg4UwN3c+TtHAW3TAXBlCbNVM/PlLjQ7AyOQWFI4dzmlCFlEpDjK5OE33h2G
1C5R68tM3yEARTX0BBojhRrO5cFiomIBqG1ofdoNVtHvEoSkbMD6N5f6Y6XWUc/6
K0aq7Q9kjYvHuf1hZlt/Kv/q3fAQxaUYNRCMhTu2itDlcWdGfxCR5YCBSe95kZhc
3NPPS3N09Lho65FuPPga1L5DGVA26jKE/vITkJHYrJy4VUR1i2qJUR6ssNBXPQIH
6vOd9Wbl6efcrglfYqQjsPP1XTNRTQcpL0huOjxqA8F+3cGBA7W14m7XR62JHim2
akfup3GGvpI3+FG/Xh3zNHmpqjgaSRDVYCUe1v8vXnjZij07GBOwPzN+83SkI/4S
kNbVjRrhoqQIXtsm90qUIbR+e8fXxt2+lt+BjpNi/IfF0oojJkzeJT/DrYEh5M10
YGhhAiGYfIYsKw/pk5Ns+g3Mem9ZUK8E22WNaPoZKRTqIEpx2jLz/464JcmwJOyd
SEm5Ps7fKf22aFWir83pffmewksg1rjuhkVipuPPpzWN3R/t25gRauCECcMRFO8R
/ocy196u+OlnsFr359gbJliT9QYVMe4qECO9LFcwI21GVWDRmmZGCn330E8wbpQ8
IQ6yjj+Y4FHSpB4d2fujbnB13Bb5TogsBSUeLAwXkNBSxEJ0vJhD4Ndh7qhKiZAf
bI8UVgGYlnJANmCu9Q5vuj+rPXNrGjJrGIVLU+1ibjDxHabAIi2yoRUwCqdrqm31
OZPlgdISYIaEw/uf4chTEvTlnG9+gy7Kf5nm+GeeKRwJGzqYXVKFlwWT38whZPoW
vOa9uoTfKhfLJJamgiREL2TkwZCNjVNCtpL41Ddoq+kSaeEcvOEBbPdVzALdBNeC
SGiD6IzE7JkyJ6Fl+YmKUYtHPQmrKLwiPUHkLk1ysVwNeeWAyWlZJSiT9eEjQaye
ZMInLLcPhAevKKHgZTb6G/FZzdBvBMxTrthp5p6Rv/tyzCZujU8DguzZp09s0JuP
nEBDNnJPElT8fjvGhnKxuKcaR5FhzhXazAuQXZfeP6zSwb8B5vFM2MrOsyXjp2eN
n5yurvTpSfNc3YXhcwGluCgL1ryQSKh4zMoUGRcVrZpNoK6Ujl5RaQsMNJ/umzvw
Nnv+nUvTne2Lrw/glz4YPQsNDPJ1PSpEIWjYezmQJW2oNqHimhoPFFXgfltG0wsR
P4HCpqiz+Ppyj4oSdWFiMynfl1ArNmTEHom1U1xCAcNnYKeKZQj1IgDDvvHaWOj6
zwKyOnxUSTNXj1agANsBRYQys17+SSGF6JfGN+6GzzqJZgqDvHeJawef8qkj/hDP
OlCkH0C9sDsDbAEZUyMurGdFMCj89wu3b9f8fHdPUcxJ84/QWiTEdJHQ4r/0igcX
LogL8FJeQEHPKYwcYSaPecR4YsGz2+F10ObKNkCjYqm4alUlhojzw+0ez8scb4Pm
ESsIgiLSmMNypKVN8VxiagVd7CknFFfH3vCqY3CURi1sfZipEwjnDdTubXuB1Wlc
XbtMUC+9rTFPdoom7Gg4lwqVxSARQABQHWQpnfuAZLa1Xe2ymE407yNBvxEISPbx
iza2lRECGVBPsqXDj+okzDgLXqyGdWgC278G7+u68o+JCC/FxE61+5iQOpJsGEm3
v9VeqlOYN0T/GjVZ7b/hVbS5BAv4ffFLJNtEgXfhPN9Ndap8Yh+6/U5Odd3fgf49
hn3ueRW/Saszrke2zPg01yqctBgLwf2d+KFnNf1pOofaRIptFZzLTwp/xrIA+nIe
sJusEAaomlunEr1TTtQl1pof6otTFmZpLDMCwSnXsqTUbrSfb8B7KvSX9sQTqeDg
mF6w4RajVmi4Aw6uxImjsW+lz2TlRqFCS5MOTaYlLPOuh1SzDDImYNaWf5La559k
Bx2Z1zBSp/GcWikN6gHBSIAecVo5pah4QgqmGl7E4Hfsv1mfzUUoueZOKOAfPFwo
hnxvL/Uhd8uLniim6fSnAKFFrgSr+TD6Bf0aJn1iHXz0OsqG+vwuD0sF6BDFMsRz
IE9ZafVUa51KiWBsuA2U0/faBXHeNitoI0sWtjMuyNyMf/Mprz1i/v0wLMSmqDcN
/XVcxT6d8FtUtC2BMQpcv06yAvnvRf9VnkiTRfuKsOiAGgFZL8Gr8EEKMjpvTSg6
MqWhi2F8h/quRmEtSWyyzHabxXPnru1/wWCd20jpF88rXydGkd6AKfB/0RwYqWDD
i8emcioi4fvQso0tYKWBwt3vrTBFQq5cXviRFV9cEduZ87/VU6sHmTQ7GH9o2rM2
h9zN7iyxQyZtDo79fEaHY9VHWBixdwT9jLVq5zgHtn9/2FlqbUVNR/MYX/XooN7n
EhKlikQMzNGoEgwWxL1ngisdEOEVFxiIM3IXLEQGL/2fhFCg2KmJGWlAOy9jA2A4
rhxdbh7t7WVm6QJIE1C6gLn4eOxPAAW2hcsD8VUjpQce2mPcy+k+9I5LcBmN9v/u
1k4jmTzAlGcZrrTi68YdvAuNxLuw/ZSJFDpaczSvynGJHL85gffZ++9sPJ1GoftO
YEBzR1HToX/DabMIkYpUY0xC1nJn5XlWqEDWhRFwpytWX/27pBMTOiApilt9MZ5i
HdYy0MVGo/9CaEXn5RqS4PJ6zTlAiT8mGMbdrc7W6Rk36a73tUpGQHvUSL061QaM
x16qkjZFuLKwqiBTsMjKhGA0WijBgHQXvsgYkcbAHXiprIMv23cd+W+KfzkcoJXt
CVwg3oTCcgQHHC3jerELV6Oa2tXPTUOM4+IDfZSgPAEj6biALbJjOdFjifzJr3EW
qaVc5hSR9cFP/H7mkOwXaZxYNX+n3FGNJ+UleMhcCYe/aJMuYOt5xnaIWiURzWVi
ornxbEHnCoe5IIIHVA2Nw3ZdHhVgaKwdfUwd3YqYDFONOXqdVaWnS6kNTUUV2Hkv
Ac7Tv9LOvfDhW52cKYZOhe38XmoHne5E2WiQCdpFa32CixefG2Yfc3LV8v0xIzY/
TQM8dVwkAtInFwJFUE8RLKTa6UroGczm0iKvmBtAgHfQy/BopYssSN43wpPIyO39
CjdkD7tcb35CMSj41yHMeEFkjgo0ftxpbtZBhZxyY4+ObLp8o4s0Xcss2HM9bmAp
MmJRTf5OgFjJB0gPZBKIlK4J28y8OUVF4mmd/vUsunIGSIy4mBeG6eBWT3IKmYz4
iOCgNI5nkxlEB/43f6p6d8or+GEpPzEttHKHKPhzaKMxdm+9i9w8A4eP5+Z4p08W
+KMjx5ksszyMxzHxQubHM235nk4CI+jeHbHPm+5uQrnp/fhqBoGDDUz9IkEUPPGo
+vQ+r1rUtR437T74TkFnbPagsKrlFM4NnrNIoMa1kEJt1fiHM9UKGcJLJ0zm5kJ8
JrA6A0Qdk98EoIqnV7PbeS2zkdlGCp9ywFA3clYVLFy86hr1za95kG7vuvau51aW
byULQ4A5ysmKfvPIvx97Qk+noXaQyyT3Iu5y/P+KzvT+YkaYb/ErxoBWK6lkyeN6
qiED4a29k/7RpJwQXPFwoHzzBOAppzfPjPl5Om39AJpHFm0P44gqjNESXzk6kjSp
rav+ZoA+gjUtx2HMXYD2hFe7hfVpbkqV/LjxDV6QDPapQal7c8vLzbJphpH2kNii
Gzsu1p3X+GLl11Yo1Xec8Lcv9wNBm24opCKhEt8aTzQ=
`pragma protect end_protected
