// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:31 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PG866/tbFXo37+KxJNpC3gba3sujzoxbJmpLMPOjty+xDD7rt3a71W8/9dDCbOt2
MOyvYSsIynMnjBcllobXy2hXeIhUGSRw9fEFprb2yQdfcC2Mn0+JqyIJs8D8OWkZ
MLlaw4vnT025a3feQXEhIk3D2j4L4BkYCWtP0xA89aU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 762352)
8mkeIpV9sAGVi9Rpj9dIN0En3tXgVtKU78zkP084hGXmbbGpTO5M3PLnCVN935BJ
6OlM6CC7++qUNR6JrMCnLia8DnorKjQkgKBXK2qurDYu6vR4V3Fe/jU/Z3vyzU49
/cFIRSrOuHAwpdwwUo9Wb+AGO/6ZECtZ6TWM+bdzNS5bpU3pXBhsh5E8qkr3XRHb
c2M5wLcTu3XmRGpb+GJSyxO8o5IlgKBJUz66TqWoXy7IILYmf2PIHKIZZWlXDIsZ
5X6EGuxo62UGeXYUMBILS26HPY+0SeHOt9fwuCiBtYWuYqeIgxZl7kyxm0x4/wJs
TMKkNHogUgLrHQAdQW9JtUNixDYTHOlO1dtUiS+ZP5O0nm0VYiPUa69mcmWe7INt
RBzl/kE43RJdypSf9h8aAoQ9SvBLVPmSDKnpokFOCTx0rWNfKta1QRdYzqCORIq+
ATvKgBFpLpZNPuJf7X8U9Zbyec+TEWCvG/vmj0FKRBnYwTvFXwd+sBldZVFgTxUU
XzRA4TdqfIHo41hz4yO5UsdfNSUGWrlqMMXb/xXGykRDCiHqzWoC1mpv0/I1k/VH
DYi2HahgDI4rRXO7AUMSfFEqtdkd0bKKqEQV/7NquVrs5XOVrH2XTTctU7XxPEk9
TIYSKzZWmrulgE6twoqmcGSIy8nDykWX5eLxAZOaf0lkxl/Woybf5dNfjc/Q+sNU
agGPo26ioOMduQqhkusfh1XURNydGZrXC05Oyh7559yxgYRi4dmI6Z0znY7NpqtQ
lzrLHIARmc3xcsb8dewjX5yoOr0V8yrm4kgMdb/i8LABUAQDn9OLfzJpDBeUBnhZ
HpVJUxEUFIFD6qHhK6SHHLClwXozARMcKYtrZZ0aqjSy0TylDjrcnxueFjN9JFaL
wmUJTsAttxtFdq6yzUcbhM74tqhTsgAGayaz+NeCMN/YLkQ9siKuvPgdJZwJQoq/
MTeGAYCnGeKXUngfJH3G32aozrLHqPzJ1grhy73dDX8Ry9jfspa4aJNcrFXt3r2p
UdzndJTCTZFP33DDXojO6ryOVrW/feeJP1mJdxv7A482y2mlCsDq9lQGM9i1u8Vq
LzQ+RLScFvykehKqKBiDqElsqgabSVARhSBsow4TYw2JcxDLyb5HwtdZKm3nLlLx
rY6tJUW1VQxzAgerI30bCua4LfjfRbq0zmjBs7tV//LWDlUsqw4pammosqGHgFQn
VKpXdCKIqQqmPVlNnhB31ZCvtw8y0n9RZST0xS/cqbZecnAI0PNlqe91pBBSAAZu
DEBxKWFA8W42fWwWs6Svi2v5fgtevKqWt3Db4weSe4ItQCWSITO02A3jwLkZd6Ma
L6pnyGc1H6sbuiT9TZcLB4TRKyCw/mpDFb8MF35VfaMIIC/17e67eNNNrJ/hSgny
UXGJH8B3t9x8q49THPMclGPtZIw6RXTWWCRwZY53wM2FlTqEERp5GdySp62Mb/d/
x25xp/ORo//poSfeQVEgmu3uVErt/+VGi4E5EsL3A5hAMoG+uGfC2aGR5xwspj9L
UGy1X51oag6H3zY+VyWKQdcGlTqbFr1KxmhGRVaKvRDco98N8Wa9CY8/2qOL7HLL
6lwz0PTgpc5Ml7NTOqCidUEbr/3bIHMyeDx997DDygQZil+OAE3oANJnPaNlfeEJ
nrLo3w/3AoaZ0wBA+Qf7KKzTXQSuZFS+dvTo2t3EJLhDkrWNr+PCDFc4argCPHVL
gDicPwVoFrqs+I93qGn0pTOtRSvpO4LYnFnk7/Jh9h/vjcQeB743wPnqzzBEpxno
W+KjrrWJsXaN9GbmpU/dg/KL9UMFDahE2Vwxo7gxuFO07Q0tSQFsFXWXcrZ89e9h
xDjjlpoHNU9Hgqf/kySjXbOcqNGBpNNYSev9H1RDSA76AbL+9w1Mt5U3bbBwuqqn
F7gZJP0nXZpP0Q+53j91P0BDxZIw1FEQ0ZlOqAhp9wKMHxNICTNnc+nN1CiLPIB/
EbjvCnOD/plpcUXIzpBMBMgSGC1oPljWaaJqwep8HGA+n0xaGLdxZQxRUV0JiXwb
SPmag1vre6QHlHnzm1jDhfQyU4GygEdR4rDhg8dd90ND6WKfLoCVpVJ7H/RGPLeZ
SvLeUcTSHswKJVIVYLnlDT6Zt36l0qh31MbnOs0iJpMXMy/ViNRx9s+3w3gVKVoz
zMzKLP+CHGJBmYaQ2EvToSrIrBSaPZyik2MTaiPpdIhFhsERljn5WcAsx2PN4SmJ
YAdB0eClrD9Zn2BUMlK/DFkCDVsO6TgQPiO1rrXt0Ny4QJaOm7Ye/LMgWCrYYxm1
SkjzV5VBpP+Vc6R9Dp4P5N/Kwl9jyd5gBkBo6rVZ74xIxIFHbZIUQooC2yhb8xoL
SBDaN3qcuJtV05xgXwa93pumWBAGYqKhf0zOf251vcobPgSDApvi3cxtPeQDQGZK
Z+g0kMRl3SeRY33EQLY58BUlQ3IAB384/8IYv6Xs6vxu1P2I8RFsKPs/zGxvPR7h
l3/32cj41csLMYap7f/HM0kdBi5vqswk23mOWH0mdxVGgPW3cKMWIfj9xlfPhBTJ
7Z64GbTVzXV4I+LeNnLwTewH3V+O2ztcxo2IQ39U1x27dfsk8Ol/Nw921n+TCuuk
8gKQfTO3Gawbo+utCPLLh0qG2VrhL7BzKEyn01iNZ+3+yOzpilCf8C64+AHfEdl2
1jCq2U+wD5vAZWvBp3zgYgYKYbO4kGzVPH4OLUk0PwmbLMO8lUdGmfI1CHuoaurG
j4RxeC7ru0ielD5dOJSNJgV5N+1pigmGacYwihpc+ln2/l9Qgj9UJ+OIcPDiMszu
W/H1QFamsSzg0k8/JGurpRVFdWaJden6vjHuSKEEh3stlkVkTB/nXUZ8MzYIQpL9
BhM9zO8CDitbm28ZtRw78oOmwJMc7nnHqrjTTvnwJSQ3MVfLji7vZ62n1byJj/vU
8D+4uRr0zfBqK/u7GQIrKBy70VGNFbmZJmItUXrczrvOVAQevHse/mw3twZFV/r0
XH8FKG1dHXdEs6NZs2xxNQSLhQLyQhqzB1nMaBH087jPwGjsYtUlxbxC8fb7GOP4
afA/+g4MK1w5Xo8f2fMSJRa1oRHE12VA4iBvhpnPlvHKWKAINjeIxTa8s6FKPIIx
ampdjQGS7tdF/2hHEuS5uA6g3wjHiom3flNRy9Z8llqj1I/3XoZkzA0GBnMR3mNZ
F/ClONd2alitGrVA0FuId6PymYo0+KBXs3YqYAB79mq07eFl8qgh2Hm7Q+H9cf5N
OJ6dMV/vCAnWHgiWRpDdZ2pwv92lZGwGkIuXFZBljFO587FWC4PYBHFOat6h/obH
TZfU10vRW6lbSV6CeuBbe4MgRn1ycxT+cadKr5Z0EjuNw4nDFg/kdeVK+hyBGEbe
DmJc+Ypw+GFJ01TMbLpwIQLVssiWkDuk2UbgqBhqEHu9v50ShXnC8TzjsrOmW9uR
w9v7Fe3DvevAEqOUzYtL0wAIx7jR97Lu32cl2vr//PtNPQCywfsPSLU/e7PDVnrO
HcJ8D5SKU1lDlmhFbHBBkdlWjL/8o3O7cup5Jrd+KHNOGZ+pYBVJZU+t2HSAvgSx
Wgq6v4Expi72K+DiYdKtBGxmRhFNRL2x2j7WAX89pDrlxVuI3ZJPlxgpF1K4vEk9
3gFAgZd3RKFRrS1SS5FuBGLvOYez5GoNbtysVhPAAhI5itdFDAoDupc0NoCAahnG
MLcmCWIV9Ci3lbgCTzwcA/BzC8qpgYuxFjegmOdsb1vxHm0q2diECs6x12LCXFCv
gIJSAS+tjn6+3/pcUjJeWv4P7uCgF9MZ6miD3K8x9+IEdH+ivQ9n9tB7IAaViiP3
kPKTgww+Vf0t7RWlCgcktWTU/OwwFvMqbUkAdT7vQXCvYtgvONCdSXOy0sMERJzm
pGtnQ0KL39IJ6U/lzW5cKmDa38M+PUfIQvJJghTU24vjKvy9kzomnpAFsOkBHM7D
6B+nUNjyG2B/RWDRwey18HYhx4i5fiC6jcCKcZEKf4isaeneRzWWrNQmw5UjQmCO
UEo/6o6lOVYrz0oQNX1P51ZHQQMvofqppfLZN0+2+voeAIFuQ8jQVhBLHj1HW4v5
gBhhczda1xWRy9M1ToCcsXSsZlOFJ+GgnaWatRkxFLAukWLGuU3E32psxoc7Ms/8
MLThBnjMl/5fagUmz/6llmezF2D5gS+bhmVr7xgXjgItenf5+45iIROvsi2XV+lV
5Amdxt5vIfO/xs7dEdOLGsVPwHDKUWv4igqA5jAj4ROD5gee5/90PXWh5YnNed0w
GCzwvci78H8g+p/jgASCjCcjavdjEn1Q4lbXJrnncWRO8p5QcTsznMtLjdNdGIpC
VEyJlA0bGtodz32At/bzV3Y2Y+PXCuISvLFnCirsg5bmEooCB3Ou/Ont1BEVmMuW
OAR1fpWLnix1FubMLmtmWTZzSEFYJGl72T0NuIZOBlzHwkFWXuJbpLZ9ldkVTEhw
qpvXHP0oOchV+esnjA1LHVvLEJuUFt+emg4Dy+nFrPmunYCTk74ffoVDtlzBD1ad
AORmWjOABuWXdrbA84ajOpejKYZprBWH2U3m2+ngepVGTtha0c2zjWKb9LTrNVec
qbdGwXNlX1jpWY8b02bJqnjdSIfXl12CxZZGw24XAve9f9Bw1LhwW6b1AwedGlXK
edy8z0wYC33vroeEsk91zgBGHMdHU51/NJeGNWI8eQB76LygLgxTlwo/JxxrcIGg
d9eQ60uok35eBi5ZxQeVhmTISJaUcjNCOlKYn33aPgjU4E2LxD2j5ZAsGDR4g1R4
JgdBU54ey+OkKrlBlAFMT6isqSk/SoiuA8Y06erfP4M7gvVQ3jZANMzkFwV/yC3Z
CWUN1/AVwAvye+ouTQTkGOtCZr6sFuong7XAuo3KQLb0iROrSkp90VUSm4t4VzF4
E1guvxlUHQYJVJl2Njc0x0Bi5O4sYFQHyYuU3POxLLY8ok/JokqwACtbXvAjpjhG
PhyQhrz5GroOPxYAQIIaeI6JHgafE80X0SCjwN1h+XpT+FClLkkbuEvt38a/6AXf
e/2QXgj0pouomz9GsYV+oY3LW3tfj/J46SHeXHZN9R/JgyhoqbyrHaW3Zhdfs5mE
drSWmx1bt71tat0lU8q9UoMfv3b3t5txljK+FPm/k5MfiitGUj4rsgm32LxyhOFR
qIjb0z5i3+CmhL9JWRxG/UgebhLzXLsBxVRMs7RGjHVeT8b/uHUc2E6DFj1D8os0
kgASOXDeVb0svd/piBNKwt8BzMHWmOSRVLryvtxqJ6nbVhAKGlaXBJH95VhkmX5J
udui9TLWBBj37Jeqwis2iN08RbGSAnXehoIWhIZ330fuA+NlSHwRBLkDA+kubfdu
8krU6+3BhUYR4GXMHTwDusTW9vLysE6K4W8hJ0yW0rEa8EoxwxUrhbdmVVif8KcC
w9Mb/9mZ88a4nxtUhF9E0cI+9LtfHu6LMv7Yl26ONYaVtKZv3N28cl1o/4jcju3I
v/0IhnhQ45sJH3thTVwFGlNdD46e47TYIdLvAA7/5xUDKzLMJmgIOqKgd2rGg/MN
iCzlFaHC+nm6CxWzDhw990zRKZeFzzGLwj2Qi4SRnSzQ3Ys2s7MVjMnNA5s1nLfq
cjTWM7lUHwqRaarCXrDofz3dL0HPLQtmiNnO5QpxjA/jpO+fJV7Q4lGc07HHm9yw
vxzYrNmrLEDBeTCAfuvXhLz92iwLsHbhrBnsgbHJOqBwi7Sli8k4f60E0LlVOoL1
tu05w2cSsrOBmRHXQascBgJELcZxtttBxy8Cfd44gLHNWebesrdp6+8cGF4/zCEh
GikophO2SssIfL6kJ2yEjrfBlOPwj9rR9pWnZTJyQundcazLL44oGcyDNj+Wmk/W
fjJc3kvhvJ9rQrLK2AoYaLXgLiirzr93Thjo9bjtoPq55NIKjY5yxOu5Pnw1QUBT
sUXfaCuat0rar2WlWM+ln2by8kqH+af8Xbc4pUO9mq/ceFHMs4dcnQzNLZzJgLic
N05+ivJb9z25CpVx3dH/cbPESbTNhWJEo8BzA7iUOTCZWxARCnvsSsb6t/aGU6tF
uQkyX08Zd+M3FAUcw32nDQinEpYSCGleC7h46xJH7UralOeMUBOsyI2TJV7RpwFM
nogwIpYeVVo5GcudzDVH6C0ePEmsrererkMFu9zSpDcq9NSLZAR4U6LNrSQK6N63
P56mTl7Yu8F4MlayUmxcWUrcgVIAoGyzvlAvfprmGaaZfAZgl/Tx5xnBbwk8kH5q
vg40nGkFxm9EW6K6isfe20GMnjM3Kq2Zq6A0wuAnMBtveXG5SgRkrSEWF979Bfiv
+3xMzZAdeQSm3I/SHKIGhMt9jEW38wcrNpYzQpzN1/YRhSUK0W0fEt0M4XEtT5bX
MWZ7BS+Di8tn2qbP1wI1BBomRFqKXG1e2lYUn6OazR3EDkyopkL8fE3fmnUx1sQf
PbXvg2ikhPH+C80q4kRYU7Mw50pt7zZlbmQjAA/H9lsrilFlYepXaTl1aWbo51Rl
YHG9RI4wnbv/eEB1xl/N7LwRqIGikFWgbIXjHEjoDFkBZXcrF3M+tOlasNtu+M8/
Cn1qDV+azZ0i68EW1kkOb/t0jjVY3uEBjVZ06S+fD5p68PfoTR3aJ585xjgYz3mN
zkYTxffmBQwM3C7/ZKO7bQAtDW/YsMkLze12TLFsRLzZWVNOJnqMWhE62wXtJiFY
QYHgAsgRD4EWbRITCsFb+WeemTU0DhnTJCkXTXPaVOHfGZwiP72yuhpLS9HoIHgx
fyXC6d6COT0xPeTgTqIsvlkUjc84447zAY2Wunu/Gp30PNYEMyZ6UlVJW4zNUO80
aPFsrT1DYn+cq5Jt0/TB2CsGvvC4ZjaMSj1imOM5KZwArd19T0J9eHxK/7iuWhm4
4IcQaiN7jQwhoj4bU28BpaRc9Z+PTquQ2zAy1c8Oj5XlErLJLQYQnKDBi8RpbRUu
kIiIM+lSPFvhNZ3SF7F48G6AVhLENbuTD9wBZ9YbMr9ArE9nO/TfNXrJtrQr2tyO
ygno5Q8bbu3MhES1t6Sjh5v4Cod4LAOEOSzUTbUIbqGNnCaNKVIVosQvQQdrnYbY
hBqLpHhy4cFKJmAsIKHlco1dU7S9i6T//wq+T7TtlE9cVQ99lkiF1yQhFSiD6nzI
b1WFUBlRQN4BB0m7cNHf5NlfSPMh1fXGgmo6tuhno8cXUAKnISaf42yWEJhnOYvS
xIv77mX0offTLrSRofEgAu5ycZd/WURYK+yet/QuzhLXwd/oJgzAH9FxH1h+z/xV
LdRbVy381EydGi7i4gO+AuF8yP3SCho1blEz22sMViNivflOV63cYyaNDyc8QOZY
SDb5Yk09NgSVs8Gz2vorTaf/RbSY/z8CAGf5CNnVHeHBTRcjlcNOhjbQ4uzsLGms
tJH2jVUCOS7bryytIz4zW2bWKeBZLJ/A5ZLtiOmr2AtsF6/wtoAawTfvfsICEoBO
ztCb1ABNIXYCyNeV3aOD0h3XmK2XDgxN0KD6VNsfmINUIZDPYava7jUIOoxsccqT
oVZUJ6bNbPkL9RU8jbhgS/Qj6HarI4J7VE9BoJW8ebwe//67Rnv8hNLdznas4aUw
c5KpwoKhKtCt9ZB7p01H6VRxGtJVmjsmVLs7qz6yUnviAMMs5QHhXQD9QlgjsaJX
eazL5cjc67IviKTAn32l7/Vdipt5CUzEdMjlGfaNI2MDNMakNl9ND3qQNne4U2DD
+n/wo+/u80/gaMbSRzlUeWYrFXTgrMJUVLsoXyEtl9PS0w/4OFeQteMlzzl3Dfpr
vQfXN9r8WLrKanlNzO1MxfAnttvPGwxqu0zTz45hMlb/VgD7iv0onaLys56hyTFC
NW7dQmAztEVRVm6DqQLOeHXSX4a7PHNoHauQHXz3yc06DXAYc0KnjiDEBAyefgpt
o2QwRY0RM+WYYsRcIkZxk55Hg7V9MQAfeWS840+gghJ4GGmaniW0yX6EIJIQ1gUt
il7DT1jp5MFFMrVbtwBKc3vosNQCyuQx41Q0K3GdwI6WRjUv9kVxF0Wihfq1k3RZ
bBQ4FP1/pwoh50Ven1RT6pQLbfDUeqjFRYvTWteorbzdd3qVS8n2hnEK7U5lB9KD
4qwQjjIlJXNfE0eIaCQ8SQw0Mk6uL/LYf406P/pEPNh2qSlZy0EUeIoVnPUzFNw1
NIf8HPuC0P1CgoUt2GHyJhnEjWzkb9z1VHSrTBJbjJVyvxQyygc/4z2+DiX/AH3D
6wQZJMRPtL07VMYaSiud27aWcbZTIvHMcldVnUUaxd5zPtwSvzxUV+/FAVUdW19J
SxE99MaBivn0/HmbmJqgl2iJ+Qgw1LIAaCOdXY3wNBgIHA5yIl7gWurJOugPBdDv
akxV/R80t1hKuZRWmC4+voyoAzidE1PkvcUQDYAKy/y5kXPpP+yKvtzvhQ+a1o61
pnG2Jgi6CF8myYUXYyV7cTglp8bfyTE6rmylQufjQ1Nlfvzlvn+3bwTtcRan8yrG
mo/4Y6l67aUOPHMEyACEaVizJrYH+KP4gn78VrPZI7zEKehznhCyTRfeuCO1IdTl
Fv7eZhtckhUnDZxSHF2VHgrcO51O2TqSB7wXtK3Yk2iXNwgQC9PowvJ8EIaUXoQU
cnf9i1USjHc8MPqmUrxBwV6zNdIRdJAt202/kfPfcuONwRfQXWUNLJn9EIMVg6zX
cmz2wI4SkhXA/dnSQ2iVq1XfgLuKI9sSPCk13lO9pADDKh2LpAugiqpUUOgpTRTE
v7Gims+yojupVAYJBPRYAq3ff4qXGy78NAFZtTzXwgugJmkNkeWdu3dxOGN+SKGp
3u1jOLTbS8rGb5ipD9CYI1cjwoFYr0xyoqVAIfbPn8s2qilt5+UKWVyr6TNFE0/B
gJq5oPVKoCe9LAz8k2TUH7fK/BzUMTLDh7U37hFgN6RF9IM/f4guFKxvFVCph/Jj
M6eor02uSZ06I14dwX6G4zV6seK7lIS0bVyPUMZsUXnDXRGXcBiKymQe7IXXhx/A
IZImnKfmZDs6JcmophHX0Ab/sBeFCd+4e5YUKZYeahbMDjG6DpHr0HxgVjIYBjyk
rORntAz0yxxnHTp9zSZ7wfKBSWYMyAfwOwUnfRpJmOQAdVD/0jks04mJOwIx2Fzk
l6CoBjQKxrqQ63sPFL9lh4y3KAqDFsTxaFcpwemjWiVhQFHol+vb6XdU5MaRGpOh
kY0Z9GcLZLZFLS952Lb6QBO53ZHBkKhfggWzfBCHL7/KEe2NMtQHADyKBeO4qYyI
d4zWVQ+Q6eIKw6mEiFsHz9btxbKlZEWpF4NO7JgKJd6cfuz711AZiv/fNUG2cuew
5ZaIDSa9X/5dKrJq9IdM1YiLbeeHHSkVCCjErA4IGpqHzpRLLG5eV94Vt5HCn1M1
ZQh8tRgVTcm5ZV2oshx8eXkfJcymn3oWUR1yEjWT3L1ZNWG57bgHWJjDDT4OEjk8
L4qR4ArCG4XV0WY+TlVXTdTwIi/2Q4itNwCNPPGhGUa3kOGIY8z1jXvSb+yeeoXl
K0GqvAjAybO7o9kn/aziF3Q/bX8txvUrqrJiIKwqDnAeQk2y/3zgSKdh5pEPZGrK
JO0ciuPYglKR8c75xtIW/isgCjNqAyomJNiC9iI0BfknUKjixQIFJJ7QC0cyPuok
WbfIf4At6WNDVku1ljmy9+wMDDwFRmxf99stBm8dl3XpDjUMCqpsqujK7ORoEl5b
0bpgVMj62Yvk0ZcT9ifTtBYP00jWbP6NRzHcp5YdPGaxl5utBr9rPK/1F2hVND3n
OLjzXovNe0/JKhntbXx/5wZwjg0GsSpyyLxynSaUUlM3tBq9NPtgmFszLZNdUSek
Dv7WnEHvz1J5frkDFEUKLj+8wRpVSiPvvbjH5f5ca2BOYnnk7aw7+ECGuY8S6lZM
84xrvA9TKbfoRjSzDsIFQEiM5YB1YWm8x0YJ2Ll3bAsVWWviXzN2/wJJhVpqPv7r
xIKxH3eqei06kqHr7wfBeD5aA89lMawP+VZkrK1e7CqI46chPecpKFykrlMNXedv
QHh1HEqw2y5oLyqMZwqDCDgFqsRsK2Jdt9Yn0xpP7Xt9OK7tLF2pRasPutYviUgq
bX0m8sHYgy/vobYRl01DDqoZunL94dDyYKUgLcEElHP5cEm81iMkgYtp06fYCDUV
9aOnPZ99O4fROpYjTmP8smWSuPMxG4oAkI2Hq0pT/Pm0jSYFv/bXQvBCE0MdnRSY
PyFqhIyhmREqiLN0l9wBAqARVqA3bjTS6xZdbEh6F4G1SooHPsBLTXr1fxTwN8Db
uXBzwfT7oyP7uOI6O05YGU5vda4x1RmoBNjOXGqMbiJVBkumiJZhPbIwL4f6aFAm
ziROVY+SohyCnta22mRGiMD73bqaFvn3+Ee2K+c+t3ysZu60/PNqud9qIrGu3KDI
db1+iDUnCG2RUboLmrqEfgu4xf4oBzdUUFOSGTRts6qoQwhq3cEwbkGOptMd0JUE
04toelDdEnWiRNfNuGQGj1nwCCSP6I1DJAneACVmty7JU4Voh097VS/bZ1Pjj4E7
WJ2YQuMhc48GbcHrgLUARDNXDeGpLv6EBFLoBrP9P+J+G9nBr3LeuwoMxzkfuyOq
m3ArpmGWOt1GPLzc+f5TW8RwfwVe1wUQeqkh0a4G+2ts+kDfm0Z6moHZGRo2PvBD
MDWtE6jELPRteTmvUGMvV8Bcpuonto85n6elI0Ia5UdMbaZ4hdA9Lc5DX2prQXNi
Vu5kcbQ3dz4whbDSerPTMenocXfAx4/KvYMoQLJwG4moSQGitNZ3/moFbK9fYx3+
3YCEnrLk2C+UAYYT1DjMGBf9S1eKUQcH67qalvdxX2QrneOiMbqfU4t7z4fiiDWT
HbbmHW2kmpBeoiFtXHMjujzL1KJ/ftyALyy+qArWPtrUukYfMkar1gHFSgSASqoY
IZr8yDidqWiT4fUYCxQzLenmwhd0db7VljkHPM2JM6G2W6jqgCYzSl00noPgnoOI
T38GNKz6EVKtwC8iJXMSF62hQmQykW+vSCTbdA9PrV2UlKB7fk0NuTFN0B2CHaEY
4Dt6pekMJIDNACAy5A5dQOmPmvlZA79elGZzBkzFlVYSYOYG0PexZd0hZDFLx9I5
rl9PNdosS/UOGShZGtjxvxKxhYl4FH5nBcfqh0DO45y9E4XARfEbRS4NG9dZNy58
Qj1Lt4ICc37V73qZi3R7rHpriyVV7VX7Pqd5W3+t8JE6rDmdyfRMfNz/FYiyMD86
hG8EdiJS3i7/U5dV0cPMczV5fkFBQfguW//ARWd/WcEsGextgTqqviNA3Elct8bI
menuixszUk7EJxEsvnJEr6o0ZmiKG4QFC+Lv4e1tQHeRN/mO/mu/+yIk5fHe8v5Y
HkCYbzHqc1fChzVFTrrVUeQhyWbSvoCzrFimJleC0k3j3aQLHxmWyhbA50++4PxW
/g8hTuisoGwBJaGcimQjXeXZ7Qtc+9NnXlKOxy0r4U7q4KUgg09G1zPFjdtryTQy
oRzeV9AO8nhItHO6zO4n3Zv7EjEvog86Yf71m3gTe1bJsE1a+z4xcUqaUSsudx9B
OMHlk52GLkEB14wHZ1HJz7DQFLlysgqSh86hKPFdtFmVemIJYIxxWsoQXk7+tV6v
Py5tus0qWwZsNYqzk3mD8it7kkZvloCo5n1pZek2GbbxfNTDFo3WCzLbwL/yOzvz
Ls9bb7ZqNGCPa/qxu2R/QlEsDa1+41VtuqQOpD99xFNB1Fi6JaksdVsDyo/nX7ph
sE9W5AwKwW6pHDsM62ZQ8Y4JS4P6P7XQsm20pMrZxcoWbhkExWsUxNTGmvSENIlo
TxGIL8KdYB1jxQlOLTdV0IUFalzq/poMwcMhkFRSNgyaJPLmDpD038xt9F/5u36L
6nLT1EuKkVHlEi6y3FeXbnRW7LpgjZYf5EsRXwEKa9wX3+wtg7HoZBuqNLnpn6GO
9yvKYmJvXlUfQA9V707on1DCmpgFgJAmVmAc5zElhcISR/Lvq1WBt84qwRlT05d6
8h0ak1t2AM2TVWek9j1FlUkPaiq7/9YzEmVqp19ipS41hSX/Y+TUlbkWfIkN2Kgw
u2sEV8ICsdqYslIpjITUH/huS/dDOjbvKqW4QZ4xUxs2VAJs9Jyr8WnsT0mpU70p
DTIxLPwy423kJYguhCWmcI7DeZMcwjOfOHprGd8GEhAp774K9qSpC6XbDCFJmpCm
7htdhSpVIimO4eRPDa91ExXbURIebrgkT5eCBg477wiBPbpxazFRE09IxTuc/oCA
GRc4AgXES83TcAmto9nkV4WM7LxpLjhDjOMddpS5mx02qxKfzKD3kKRp28fL8I5m
gO3YM4mfivkMY6vStCZioB2dikW2bUjGvMDuJ1c9w8QhBG6anmS0apo5VQ4waF17
9rtwn6H+V772zYnEc+wUcEY0rXgjJvH3Y9BLSodtOcMy+p8B4KkoGbkwXun693QB
JkTRJQHwZsdj8MVxH/rmPpK2OfAC5IbRAW3rGHJq+BDj+o3IWBdTxv8keMZPqJBg
P8xig/4ymM9pU5OKYapVl96xtyDDpKkhQ5NClr84FW2dzIb+y10U0B9zgdy79Klh
kMjBYVzGfpxcOY2hTYBUA2iEjxbGV8tBKK8QSYtbGkis34WM7pR/e6ZgfegTZS2G
HfU77EYYmTR5MFDS0XQtyws18OnEv6ovV/tTjrucie316qgtYHBW4D086rn/L0/p
bwTakrTtjX65KZemNZyf8ffrq3f7DJMw0fV6IkmdwQ9AkFp4JYCrJre4uelvsBEz
SZ8qfFXTF5g6CS24T1d3bkJYyZTu3Oayxvmnzxdjn9KGLRJmZd089TzHKNtluGr2
ArVFHHKCyWSDzxaZtP7PVip+bDX7dulBvcJMXTK3hgYeSBgn/eFfXXzSF2B5cTnw
vs/pVdjEo8bF5FGNtmZkr7byvV6V3Xms8ClkK4ghSJusNjwJGfg0Ym60ew63HXjj
Cd4j41g0uJmilD/isJroDN63MiLroVSFg+TXemJDftekzTthizX4e3060yUtNns4
ewpOKRrimkbDPsKFdHLrKjCyGQ2soa1SnY3CTJbcVBGfyp7TNYFJDaiutU41LnDF
19fccTiMUyw1sxwVnLcj1Zt2jybq/R3B+aXutzDzc4WGt/PVB3uDgjq2n3A7a2zy
7oiXwliBU3uHEYW8Qn4omZnCm5j3kBUk1HdynpLkCtiU9NcGcD5SvbMi1YctRikc
1sp//gGk/BjURWxQ0ffspZbcsHt1OBG7iI6icUF82R72B5XPGwqqUw/yF9SvJlUn
iOmvnuB6Xu7IrQAgLgcLmfeGIwD55fIeM0gNu+aLzMsgeezkGjLgEtF4Yu15VE2z
/vmkgmkuNELa9TD849hzK14weJSL+VINZ5w4qivYhPtKOMXgPTHBp/jQCZqAfibD
dQ4mWk2P4KBo5CgCidJcFpYIhK/d1T9Ewkj7sV4GTWvDaAfGQDTJUz18llNCEJpE
pgufZnbCrfmvfkqHhsDO/+pqvjJIgkt0VXL3i9wSjsWtRiRVxZ5rYSruSsTYFxFM
QTT0o6cN1F5vaOmUyrLgezbYdb39iZIlnyVgFNM+2BUSTGGJCgiwoiTvnMPy57G4
MfTHxeBYNMmKC9Pr/G4o0WwZgZm7+D/Q2OBqFGI0UzE+dhTlsXJcYl6oy2FZg3ut
oJNY06KW0JaB7YOpgbt9zAXQRWs0U/jrowoT+Zua92eUCulGTbSohUGnwUygXfO8
Z56Irq8XfPeLFUERnHxoUOgfUFcgM3w2omDjZ8i8pGXHswv6KGepEli7fz97+LqM
IycubVJqw4f1GuTHbagaasw9yrJ5MmatEmm2jMpAdKr1g49u2PsRthI34JJ/y81m
a23pZ7D6J/wV9g3VHYgk+lnELSSCJhYHykKTBlzGbncwehB5Q7ag9IS898Tbu6mk
T3tWjJk7eTn9pKUdJonlDSNc3weXiIEP/ooCxIGIkyuAHkpxI3vVX+c+80DgRR2C
W9c8T2byjYBOeUHBG/KKyO+BHfCyRsO8nbutDdFtXwOTVkg702OL5UsHxTrQgkUV
MhuErlTO+c5FsQKagEyqtQTYFDkmiCLHtYSBcxgdEN7k/cPpUJEyN68pXuvE9RUL
wZGYNS/AUt9E6+IjmaqSBcn7+qbgdEeD33kd/Nuvt1d1DOowSx7dCn918ih71kfW
HwKpX0Tlq7TH7CZozNZviVC9uM3/2vOLbPb/6ZGYTQPlIeNiUvxLUm89tmX4XJH/
i08VD0qctf+W8SJNHCBNoYsE/tbo/b/5AVf48mHIqS2ItPxE1U8Bf7ahmXw7ixUz
maglHSKJMJlIq6YOex6HDbCCRCMKw0X9qSAhpVorchnxLYQrijUn272mbZZbO4MT
C8fFSTlXqqvDe1rScajZ0q4UoLc+BJWF0NUi8V086+i8H1Ons2CxA5yrK20wrW2b
ifyfOUL8jarNQYaLZxcyo0bUUuJgm9gcL/bU+9xdwAAzf3Soqxx0/EPuDb0MkxgD
GBaZKgJv2r1mDV13+XgzB5FKpF/NkeRi1OC0zoscdkCCARXEu2XoGdUOcrqIq1g2
QWLs2X31fHj2tBxxRSjqVVx90hYYwFSkAWRoL0pbHYuTphtdKZzLKCXkqkAcaMJM
i9YuYCI7j+fSM9F2K1wU5zgErVg+v/CmDq8BV6i/iZVUWIy5pZAIUiEBC2brUnXB
NzBzHy0kfm5nUSsw187Dy5Iron1ZxM+UDr8T03vsYzEXFN2p2kBHA3EstOgm3yPM
CcfzZLGUNoew6PNAK4t5jBKmhtJLUp/aijysAopbD3geli7SZkXRgchliqT5hsQ8
+5AW8Se9/LSWvmxLU4S9N/lTjrKP7rYPhXQbg9YUYl5LHbKq40vpOiMopZTJoJfs
5o8iSYEK1aXDXJUBxL510h4fXkqRCj440rJSsxeJ5Zgszu1Uwj1387M5iU0msOAH
fYy5iqmwd/slxhD96NXgWpEezPU5TXM/fbaBbud9kaX3nPd/nQK0UcvlT27Aydc7
C3CQmhJMFTQONZIRIJKlGBnb0hnXWnORZQHclVsgeSKRir0YuNzVthGILxUiVX22
HVa/+oc4wlNj/coSNgGBkeb251g6gcnKAlVCFdNaD4Gtd8qX4ka8yfmvVx1KEOty
Yle59110oiuhMhn1xdLsDeyMfpUr/7vVknRNIgf6D4ZGV2NrkRsGyLt3pne61coN
tmpqT4pWEWHGy6CdF1oZSnBZSLF6IH9Mr+mhVXzp/XGY40erNlF6mC3Vz4rvrjBR
mJcs0l5k6cUN6dvDM6Nl68qLA4MjgsyAk6CyL8tJpHu/xqiVi3oQlduz1jm/QFeh
UUoOmQenG0q1xnOCBMg3TVii0zmGicMSW8u7eVbIIK7tovQF4webTqKqfN+wuJC3
KgpB4gfFepq4RgPRrACSIZQCYoHigSlzHbQNnt/C+Tpwa4PfCG2SqWdnPzFcPQx9
RXn1SM13uVtkGJK8XSK1AYvlH17Gw/q2sRv0j4n/mqc9hIaLJkHRC7nbX9pEiAmp
GHeG95Ba+1P17V4nlWe6lc3xNmwbtwklBg7q4+abMwGhXqtpJayixiXVlcyhrhsk
ehMij2oRRG2jT0+TUXKIns5In0k5LNWpf0CGbNw6ABbwW0spavbbveIjdwMkWf8c
AbXGucSmfsW2I/OkbFYx0gliIZPsWzpJAHMXtzgJ9WTThlnc5aqmpfHR83aJWuLk
zkcbo63/4FT8EHl4B/vN93yT48zEhF0BEydHZ2JXjO5bHuEfEBrSMHfGDOhqsypL
I82hG7xNQoLXebkpdFCX6G9rnQhaq1yMnY2ZbtRpVYUVNmda4sRPNndsXnZiAs/k
GDabcTrTzqZhIkw6bhy9F+sL9gMZYrToHKTu/FtICZlLmIwT0g6YDaI0BljKo63t
qjMpMR0rOAOMjWcW1YYDvmWvPF5qhfc/kV6WHKj+uUrdflInmc9FX1CXKogJQpej
6C9ajEsLH+/GwkADX7m0msgc1PLqZgyo9LUcmY5qOVthuYlwjCOFDcSAZ8vZgcRO
nCP3hDmMorXPAhH0STMp31QVPGzJV+SrWMtWSBCGT8cDMjcMMuTs7joWZw1hZdst
dV/wA9R4HWE5c9N1QpJ7n3VfKip7SiiCYIGVwSi583R5KrftKkSGx0CAnNA/Gpoj
NZfQIK2Y4fcPWUN++z97IqhzvRi3n2ioYWYumlT4XObvfNuleC4Wl+7gGp3wkuCZ
l+pyCq1Ce5HLtI143z5dVlvfKJk6zT+pcFvuMYl+QnWHZI0dCvBZVDvYaSIGBrxH
r2ZshbLhi2dFhT/uJKibrWVVKW2wLmmh3elkqC6DvxNdsVDfxHPw9d0a/vP02nUZ
/LKAsUqURpCkkV0Hz8hfy/3V6bJ7EuMZvDPDAIIsNUroZMn6c4t28s7iSFlbDqop
MgqXB+ky/OXBMsUKFI4RQJ9dE9A47BEZ+EG1QmYfF/HBu9D7Xxza31mL7JqCP0oT
N7aQmqEcd5q2TYS2Q8ItATXHgqZbEZYC3qBnqAQNdC0JcSNGeTbnEGKzWcNgKJz9
J/Rk0Gp+M2iX4+nJhfqsW5xk52nhuy/kv0oZcno9Ev1jcgajipp46hNExJsWSzY8
VnzhKWFz7mT6S3EZfmlxpJUYDhMQgmkjBzZRquaouBT2v2wpXKmWslrdyjuXwubP
ka6YxJItS5wmNV12SOYmM4Fx/njowQjGIowhaaSCO5T54zPUXFNQCQTV9nFxxHOv
lgxcF5o3CVJ5PiOnDaisME0CGkPylEPjYpFtYvIS0kHT9An73Vs5JBnTvcV3ZVRH
ymTmT1fJu0Hll7clEKgpqz4hJcaeL59s8HwWbkNej1EsXPYpvy1hJppN5tw8WCsl
nXzt4rvICfeN+a8zfRCDaezD4iIQntvskpVgM4+S0I6ujCRX/9vjPPl9d14B8BdI
Jn6JqV6NGaJxt+HyyO0kz9Fnd1NxMP9zRu6zGVPhSBFpvbDbv23dkrEWq8cyYS9H
MGFdmiGgWk/hzPSxAsKI+3a4xT0qWu4dYQDKjt4WpaA3Tv03NDO0UNWBKeOO9ByJ
f0oF8Mpgv8410hjKG/q8G5NTSuWD8r45yrS0VkdK+G2Zxh5sciqnFKqy3TIbSv0J
jlZQcY6crys/A4KH9EvO7TkE6HHlUSp0T+UYLuYGlCqN03xyPAO/bTda79eqh5+3
n8bq65HaFQLZiU/IPfi99P/gG6jo02IbUMF1usHPMbeuDJ1WjL/35WHn0m/2dwcK
u6Kb2BDq1zbdCAtVscIltLAoVRX31RNzIFkrIY4ti8mMlmNo263kyLOPJMCRsFRr
gZFreAYQD6thFRBW6NMVGt4CJRNj+O4fnH9Wf3XPb4u8NQtkfLW6A3tsttHnPw++
Nyl0Tf5HS12UJlwL2q1YW5Dkc/4fIPK0F00SyI38J5Vax9Sd3q6aSckY2lrLT4Ng
TzPTTnZf1y/foKNHLgy6V0G9UBc4lsjXFM6vJAdqFJ5vDrdk4wEZRjjFnxp343s2
C0KuKsAXAMw0Z87MV1+4uto351pKgaSF7ESyzwWEZll8VszIZ9vvOHI0LxuJD/Fe
g33+NyelWhN8hXaQCh93UhD2jZRhZ4nfSJbAi7pl31vWwXIlNtbQV1+0k5kps+sY
GkyP9HgKSMlrJQJWNGMC/U1bzl073IJ1otNaeqzIBfndDoMm+O7n0j5zVPqn94VF
YmjRwOB2yVvSKg0u4iIc9LJiCltFe08se++3o8JVpPO4C2k2+yGAuRPdjxBMK7uW
SvDqoaQmIILkabuNSKNh365ms05STDBkfBKQaTwGBekROtvR6+tEPp3/DWXEONLC
hEpmLxKJMzSJ4/va9iEQzbZx+lIxEV2l2QRzkwWZlrF/IBxpULbsuloy+S8g2jPO
FWk75OSO0mJSilO89SA6kVwQHzKjLTAqSsB1gyt/Tnsh68BB4KvRZyAiAlhkrFY0
bfN7ytTKy7rp9IKLeS10ryBgxLg0EdTHMI8b6rIv+EzB7YgnBzo2EzEzWE2weokW
rkCjz/1t51QkCoqFKxW8WWz7JBZF3dJGg0WiMDKxq7SyKa9S1IpeQFRb/LpUAEIz
e6tRPE8Dk+hmXoKZ6FH+GzOMu3Nc2YxrVt5mte4Mm/eEjNll5ytg0bgsbiHMqtU5
kzSoR6ZEk4Pmt3aMjQ6jltUFIHkEo+EZnf1A390TlPn1PcS/KzDfKRBX18h+k6jH
orsbR3Wmz4DiIq11gc1JbIp8T1s4PI72riQ/TInFZWLrsP5CgHtTfdE3xIQ93Uuq
XHDX/pDE+OuWU62MU72UxSUTue/k2x68fGOjKBxhnIY8bU5Hhr+BYtSeJr8VkqZ4
uiWl44QJToBQNc8+qrVQnrxjQ+tbWI58fV1skKPEPtvzThlTFk9SiQRpleMJhndN
p/WLwCrAIeu7YoJF6h/CibSOH4Jvvwwp29rtaDAziNmeI6OqNN+jxuZTt2Llmphd
uwVD5Vmc6CJZqrp2uDjrpIiQaJgv/F8H4WCANsCxbo1qTb51Pq/v5QICukwCrGA6
hTwovuZxAntB1PAsEgKKlJUSd6b38ymsG0ORxJ8U+Q8Z29/ffC3cHk9+lJprbpN/
S/DdgwadKy49tHLErLJKPcoNVq5iaL0BQnEHPAWXUsTrPLov8lYbZDZis6M4JtX/
sfDa4AwbsfRVFEJ3f73tNQR6CH7q2AzNaSJ1WLsDFvAXDB6PbhezVID86WmUVKZq
UZz8Gn7myvEDC44XnCgwQi6TMaIwWHQ3mf+tZQG3qK7gs/cC6OkrjHMMCzV5mkRR
P1fUt8VuJ/psLY1P1GGsPj7fuBb5dE138Is6+3kgXSxZzw61/O7lc0OIy3LOXscz
hvF8+QtxxqNtQnBOGIWaECbGpXBUhuRd95WUZxokW8PSFElipQwoh7zlbaFtDqcU
8DqYXvmYuVplyNCKVIQoWbvokvXXaszMbTyzWxRij1h0uoA+jIcaiPilh8xo2bs8
pHz1z7gDvjCxZ8vArUsuZrCSa9ZkSILEzqPY9Aa2r2uKi0kKgNngV2CE/S/JmBiF
R5DTxRHRyZrUmtBOLhUJN5Q81vgCM5B0ux64p3ArpQ9OB0FDSPgcsEgZ/vvOOkZY
d5wxQaY1xFLqVE3Eo6+OHgdFpIn3sT8yIe0pSN8rKX/Q3rlxhK2i6kHS7hT1J1ji
dIUAyMl35hfs7wLXEJ9KMXWVh9xMNPcDPwMOv1/t/dsgiw69iNJ2oI5u300EGYlF
eYkU5iUEyTIe0dlxVFq7pmFGQEJh7EPm/NTIRTocKI5Aq1H7dzqsJONkh6rYJhs0
AmPqFoCwYldgR+dqxylAtOmTiqIQgmpDLPDfFI61dZpOTBmVctAfCgMlhiTcdb63
akkktoKeDYN0ROVk4fUIQRtXLs9+WL0YY70gMH7dq2KAEB/vfkfGOjwNsZXBg1Oj
u35eaPN6nlxK8ugkTj0+O1tJdZ0955+5H03HfqG4MbeV5ecZldjD15vDKcLDFd1q
49LlsV6a3en4dr8ajnauEsL7hG9Xz5Fgu15ky5y4z8KLinXeqyzmQ9MldjUXLpXx
O/+4y3hgJDX9xrnMKfJ5c/zYlo1Ugqd1QHTrxXVwu/4Ut+hJTky13P+TH4D2izOo
QkeYIVJhSJCzLNLGN/gWFxZBhpPrd6/lkwPc0vwsioud1mWNFExUE988sT0nCtIj
PvXoY9pcKqU6WcER/7P/41BwX3DHDUoxPiMDs4XqpkavPoWvjV0OR3/1niXFArwp
+YH5y94rQqm8bdE/ewGFj6ab7COwro+JM7f9DVSvkvbs4iaVZsGJjsBks0boJEk7
M5aG+eWCUe4OfHz2DMaW6lmN6zfs3q6bW0lQ2Uv9Vo24UThgQ0PMnhvFOwyzcS97
TEXQDzXIsMoyYceAeui2oE8VUJUvm4h46TWtoaVxKkZ8YMouvaP7irjmWIAbth43
ah6BizIrlCbXvznRxYvQ6G+DjeSzwlq99og/F9VVGu/NkDgDOLGwjMLBwa9XoMwO
Ph16MSbsjJj6kzbZgh/KKMXkLKjWbFtkM4OsPupOdOkHb7pj2kO2DFRY2q7SYWjP
B5bANz452rfwQdk4Cc6dz98Srln91FoVLJlWK/+5QNF0vgDmQpBS9vSFe02vOsMd
9xeR8iDze/1JBDlzFCrP9OhxTsMl2HvbRFz9n7FbLwOXESwG1JxETP2FSoN9y1g0
/5XHQ48zRzKjIqRYGoQyGWZwV9chr59G82M0zIF64Y/ynhlwU+zk6ZbzQGVP0/MC
tJrZ4bhIlaaNlOIg72b3t5hMtX8Ig59LzZenNzd3sQhSizfbe6sYVBNGe6FggJTM
Ta4RWee3RoFHFBbodBa8nX4HUvZ+md4v2iiVA3lnHSbqrNcfXTWyMyd3rwZbUVB1
Oj3ZP8/Bwd0F7RtOFhI67St+YFhxKqFod5G1EINI8HRw3t4FmBGBj4JgcDDQ1H7t
gJRHt3CWaZZ7Z8WZteBYuO4ufnzp6oZPWvwQ4C8QGJzLcuC74kK32DjhME9NMrP8
XR5pGg63SAhJ/PSG8SHS+1wD3UhjZw8Lbmf4W3j5SFvPKCU5dizQ6gViwWWC8qce
cWiVUEChRCnL2m9+QVg53CY47qOhGpqNo45McI8b0TDSDG+kdbY3MpFzEO7/2ryU
DpjMni+XQtNnOUcH5ugIbHB5ZElSfi/AnZon+CBQJeLejncrTUWe2NP4jpFM7LIR
FVIFCJL3zmpnYwmSEHeozEht7Q2LlJWz3nbsvh5n2RWZD8i2RC1bRZiyIgGf4iHG
5Rta+b7/cxV8m+n7dMz/p+5lL3cjBmE1/Ze5LTR0EFTlwIGbYnODIZYO4iLvK3Cs
9+6NxTsMwx79CApGGcXa/BAEWFWi4G4mBTOYoblmAOnu4EXLH76NliHGfpIHN8cL
sMNd48cfLnrZOXG/n/DNMYBbfu2XSVxlFRIE0JHti5eY2t2QWZ/nUQVpJlH4ozUz
b56Y5QWtXlBuVgwB99gKBTPHyqoKPiufrhh6O3ebO9dSPBlHYrAj9sU+ARjDhZEk
T1jDBcaDMaPMvSx7VI0vZqZkNIzvR/s1rh5bUvSu58b5hchqWhe/AYVNGa+chY/a
5Ci/lfuW4mr115/w8I5A3aBY7yhKYPuOa+nXrl+1ZLp/uIX0CB5fEFDSv8h2010H
yLv5vEe44MvDhceq/YjBPpIWgf7s6W46fsxa1FghYygy4a/mdIQrSA2HvvFpfAnC
FI+FXskya7ekRFiyMud5JRYC7WagFshlcMdTNVMNb8w+6yR9hGXcNQEsM9Ctg+4C
hDEhqdMaFNuWvR9WqYYMrr524QJr1e4dDw2dQq8iiRUdFN0Br1qDULjWSjyzKlfC
a8u7tQHxT5OnqcFtoR5qX2vImPGxopnAFEC0A9fpZoQUQTtQmqlTdA3pMCRt1tCX
aYyk6B1u4M25pyDW3wewkpGx9vWOZuKpzS97Nrw3j21n8H2Vyby88fZ+4czHDpfd
9aKwy8TBIL41F5e13SI0WAALhezCNC4kUHNpclOtgtrxx07AsYMONohww/43M/no
2ETM0jVMo9c0VJ66ajWDauRbQI7Eq0t6L0Lntv7cHg9KEG451GQyk5Ic9RAi4+ly
Tyl7TM2iYA8fhHoem0lnaymlYe+97kB9nxG6fSGHkVetc0AyrwPznXLbzPCJUUmj
iV0WUwEZirML6CvR6ZgA4rpPbEmIppzWE2KZhQy9IH+6pM7MzLI9xWdqED0u8pCy
Eo+KfzXFb3I1gzm0t3iD5o8fnfDUF6j0EJ6ody1r2LSs3dkDuiztLIDlmCcrOL/Z
xmYvKV/ciAaVBduhLxRYHi9KXg7pbBSuWBcThIKvzC/w+JxI2LFih9tOSLKdJeSF
JGHOA+6PSRbnw7vU8q1w8rzdnvQg56xX/Y7oT6rgoXqOxOR3j8l2X8oaXNv/9Se0
O0UypP5IcO7xlirqO/7OKd/hi0OSRbS5QeHMEFvNpJDcTVQ96LLleaU72sTtduI6
1weiyBD6tVfLyiU2WsdVwsGTuM/tKSTqTdtLNjqP8iaj/x2kPohCHulvVMuka8bO
mSlWZeDjg4OeJ3bkoMaHm+Jw/H90mAQuQQRcLD0A+/AgHhry0wDZDkdQTQnqHTgC
DOuLCnZmrQBnJtC3NygHFiHVuswXjxkSQl9Ziv/0AnEowijyd8mVEwQHyZ39GsCi
fcwVXcVB3nJJE7eNlmD8mxwcgKjrB6WqeIV8/wXXRg4/xDdvTPNcUybhnD/zEZtV
EoxDh6CT2nMMFMGEPPiyOJYLYDPVDdSVaLkYIJF+Osn2r8Tw+OX4yJFtxTUxO59r
9/4KeaHjzsNeGn432tMNoiK+RuOJWAinHlDCG4F44nKiFQbPOfzcEnHPJX3E+ea9
kEblL917nR5eN8XVrLABawmNfdFVbsr4oDbTWPqtNquO8oBqvbtJjDy5buH7NNMk
HihEbKfP+XRqXks+loFPVldKTeCseO2pxGIfWwnigLXkRschaCbq0oxzd9453m/I
9/ERdGQMn5ItZfyt7O5g6o0Swo+48abbNA4lq5il1IBulsV6veIUWnpzj+FPMNTr
EJizF3s+/UNq6+/52kwCL3i7LxBaUiGaArzW3YUp69CZW2dQwQTIAddOvc95uoSn
RqVSa+1JJNUksbTVr5Jk+6fDgVhXHOWMntobGoCSi5nZBhVop6f+SaLdvniCJyJi
fXWAE0L/JnPjeWPF+ZWEzSP2WGhihhXh6fplhHMfz7xeVJsgaAQNwwxN7ElX/A42
oUFnEQW04RQaITsjgGv2H0z+1qD7oCoQJhaKZ5mfP88QQvrca3VMUd698b6H8bPd
3/tJhNPhGjPYjGr7QkB9RR+dZH1UfAmMs2koscibmxC9ZBynAG9hRjtqLsYYG2Q+
F6md5Pp77eAIB5MvTkNcG6CLsYQuEW6sCwXnhunF02ZzbtobhGXWNtclsPlC3OgI
VOoiQpSPFo6H0cvVgvnnE3x/R54dn1HFN3IT3Ev+PGgHXoVe6eHRSpjaPesQTqzI
KzQQf4GNGBxzB3Ek6bmrLOsOpRwKACXPobKJsWf07lprouwTRGpZUpNJ/+kNMid7
zxcIOYIV8QhF2poNvLKkHsJKqZvnTNdjFpPorlgt4agjSTFq9KQA9RuwU8O2yUdq
Q7TC86zoCXy/h+SHoGIu2ILnR8UHVZGzopHNBc6Ew96wstUb2LhaIhIHC3/76Soo
Ymqi8dZSBeROFS03SGRDekbAL9V1y10fLfc0rWgCFQXlsaKfsRn6DFYIa4mqCaG8
AGsDNRr+AVob+lFITuHDpZ7pbtxA1gvcT3X9v9MXQj9SIRJ4GzhVqxgSbEo0Gy9A
P3OhpciYXnzkYKsAJ99nxSAsJSc58uG7/ulVGqMo1wDQ5I8z+PMM2Nojomxsk/aN
y/XdCKrQ9uRFcSLteS78iGtF4dBJ/BWmp3klOmlKdwnyGIT/o+dUoTVgRnoHf9w8
RgyRXK9X1ZXINvVczhqGqAL4kslHmal63nw2IfvR8CL/V1bKfK3u36kHRmDpJ6Ki
6joWm6ts2i9uWhxq/qR7LWO8W/wNF0p20Uris4LGglNYmXlgi/6M+8i0P1rBaBql
dsOUF0FbKw6HGa+Qj3ZKnPyIMYsSBmrm8cTCXwYyld9wA9xorXeJFS01u5Dmt6S2
jHryAcuNWUuaIFB5hwVprayrozMnC6PuKWyFHMxQ6/Pd6kflmuxvCyNX3KJYv7vq
DzgLtdhTgr3qOFjLyD8iL5XPihaI7N+0mfSZSX4UnjAzBmEd5oItUZorVPrMTIbD
xFAOqrD/wC3uWrmK0cqN1H0ExcBHO33xHxikczcAIMTfiV6QrZd+7k8UXjavNgfS
sk6GAeEWzjDWkNYh5C4KD/arL7c6Shoe1rY5ixTDkLdQ/iSjSJqV0MAPi/K8ZYmO
56cnQbK8wmOpbZPDKR+FqEjqb0bzWkkHAn26EOI1QT6Uvm8VagrxfFfOG068ysGN
LcevYfBRK/ZEKtAI7B5w+dLAda4yTH+9dQW8VvNgrhsgzqsxmeQ6sJLUAk2vQEYQ
7l6HJgP70Kv3EKlMtoI39yyz2Myp4rhUKCXXvGsufvKhTf8pzie1JveO2xycjRW6
SiiWNArT8gLPPrGBoX+exhKJkNYcEZseeG20pVTlJI8zd5YBWxsdk9N1DjSdCofr
u6M5kdoqFTGmbp8c9zu2vLmuzQIy5ysQxeyMueUG9HpjK1cs1hhIptpTuihOrzhP
C5I3M/wl0zdWHxC8KRnksoLhLlYriXp1s8c9IcYxIZL2nvH7WRe46MmzyCt/XGZQ
+xRvhyUYsmJzMf2st3pwUGAKZUQF5diVcl1SDdpmYC1cxsuwv+CeSCaXX4gupdZc
mu7+ljD56EoQhbPlxSGhBCr1ePxwNmsdWdukE2qs3iXT8xPinZAcbA1WHKAg+qJF
VjtzxtSYDRTqT3BBypPmmFynJSxD6EG2hVzOmDmy5yXG+ThkKilYZRH+xyM27y7A
m4Gz85/PGBRRX/PipV/w2RP9Xhy7UetnC/nWjzkdiOPHFbhkE+T+OWaqjSZl1SoN
ghdgzClRMz/3AIP6n85F2AHwZLN55WxLePC/mTbS406249hLXzayfr6robtHpQs9
f9qx6CjG2ApCesnr6OInASUu4xHxCfQAFYiGyRyISCj3tixL8zwTXM/b6x98ChXL
i41qiRXHCV6VjyasLb72lYGeI/5p/qD8XI5/4JlNXDwVOIU9fo+XryqWUkqOdz+f
tr928p++BpOpLcGOdQlj/724BHMaEq49ZAlZGuO6q1SfsIsiYiGdqnbKCd/z9MHq
RgUPMgtPJuSNJpR9qIgJ7KOK7YUKR1d0iuZVAWjecWd/WcWq1T8qglrzKjOaDndX
whDQwjxJCQ9L63p1pCBJZmMb0mo9LB/F28xJQacVu1x6btIOD6EhR15oASBUzmTW
sxwylKjQl02YBN7Ss2BE9pQtNeTWlUfy89QNV55sQAFWJBy8tererFqNxVWDeAoT
W92VZaGZAdCroK3PK/UmjySZbADVIC2YQh8fyG1+pbSVyWQOS7jwdrsuvkBS7gWR
QUaZUKMTMs8P5tkYyrJtksOQOzaNXoRXMrKvoyGxvpLIVmp7W+IRsj/7hkz/PHSk
jFL8KjqOjEFOUfwdg1eZb8MCG+1TYtcwYjcYLbEHPNlxVPjS36sdBCp5MEOYjMK7
gvUoEZ8lBLNd2cBgt2C2c0O2b/K4Nzf5rHKRPH+CgDPCqhPlN0gCdvyLKRUIwyLF
MgosBW4SJA/YM80M4L5HMM9fBEqGCR4AlIJeNqvRIjAJgMFh5ru4Fu/V5ERuOV0w
Xof1ERk88ZJB6LBfbbSTFo/xwLIoe3YO8MIxdYlA/Sq1S7t5mQ2VPTHK5MeyeTmK
ImxgbtbRl/tvup63yqPVWKEY5K0DnSmqdlHXqqEQiPkwAtM3bHJd+XSlepStUobW
eWqMlzJWa1B6/+q4NRCFHWEBi60LWE90e9jfKnBOCvBBefrNWHkh4KNklge0xj4o
Rr9V+o21Nvw+3IinufpnWkI+GyhjaJg2zfb4h7Pi2Ns+k+eQqrju6sf6AjdPED81
iW/VIEitE9n1qCkmg/giDar3FN/329wW5V6bF0jj/X2oKJeCJKV0615h5CQ0nDUh
Q4//Z+wSCuPCwifgVQEs+CVK22Qm4J2W+m9/k/xf9i/cXVl8q5NTunjK6X1Qu/W7
qL8/wQUO9uh1BMBuGzeeQlib179YgoRNkpk58HcNgZdZ4PYgXUkb4d954nX1n036
KVXFvH7kZ2tlibHKoJIeA/cwxDh1zBCdLa7c03gqZygqovSUVl9e52KayldwsFel
F6F028ONXtlLbzzwOBO+F2CmljudM/Lv8Qon9OuuDmn/PCU7wbF7a9MzjAis2Syp
gMUCf86br4trZKNucviepX315uE6rFHaKhUXMFofY78cW5oDahPsbWAswMKxBUnX
qUTQgsCUEpo4Xq+AHZGR/4eFH4kYKd7L7b/mML8mF5aLzsiV4kb5QDq7un38v/pN
2znJyO9FtaR79XzStmsJ3XPFc8XijpyBzSbd0OEh+2iRR/Qsr+0okYBf5q95JCWX
aqlUw8j5CdxWbA0hWZqB61PKR8xnFRJi4lQzWfm5hZL0Rdc/cibGC0quuAWmS7qF
5AEJ+PwcPCJXjTjPBphzU5eIuLTLES7ZfwLxwpMhH+HJG4AGfCjXdGZdxn5HvGHK
zkFQAhsq68rX5QN/zGiieqPeLwLMa3VE9Mom81tmPwu4WlzvQMMWa8p9/2htKRpI
9BQrOwwy8W2NMt/y8Cp/ZIE30WGN3ZtLSHkrxt+VMUpoN4/wnh4qwxNb/Hdzy0BG
9fM8MI7WWZfF9UGqTNAh71irIssuRZe3dNlmK3biqRms0DzkQAaFJP6Bcg3OOkTs
D2oS9HSibqc65DAHUaTtrwm7tlUJHo8BLJC5BwHLV+HnHfjAEHBbmNRQ7ru1vE1M
YFgC2CoVOkicLCHphr26TUDshGicC4Zkdcb2/up2Lnh+3NhuPRqSJPf4CL6q3ck2
UWVDDKt8PXIgugRAQDocQzTw28NdzIMzytACy84sjAmI1Pk6AJqjv2CCqJhxvFro
EsS5yejOKhLkbcpH8ndGBpXp/+sMBp9B2aV/7393YgjwBLh5RhTpQs9R0aYl7Bfd
Jn5v+2KaArVrNMYUad6X56xWWNrDvzTkGANwUI22bpBkcEK69MR0TTNbEeqesOhy
tH+R4mUcqMPHJ5LU+zEfv/1a99BRwIteZD/aokTN6d2oUOzO3dUKSo6JJH2qC0Qy
gRCRJPN6AxwV6Ba/W+QLy3H4ejBdxNdUj5CQMvUO96ugOBXfOKGFLuyhTnHcox5o
HEJ5ntgZWhCZWL/5gOB1T7CObziKDsJA3I+64Rsv8u+chxeiWC0Chi5opqm+iuRV
NHGdjf5AMDsnpMGh68YNXX/imj2zm4CEd8hW0qDjC5USSZaL02W5oJ4tOnc0oeDZ
84efkUs+PbRbYaxx4XYES43V6y6Jrm00RiebcnIUlecR2mZrZ7Nr0o1nlZlTRHeZ
Alx2nYWp/JCu/o7OvM4dYgp8tPFI/yI8nkInbZpjPGPFO5RxtlWvcs9mKeMfJ5gH
MKNORQqtBkyBGdYCpEzJ+CjKEMD3z/FFPSzVtKd3Unm7qZ78dqXCTFLwpsX5reMB
PbDBk0AQ0mw822rfM8mY4X4Nd0coYP2L3fLTrq98rea59vZajUiYF9/RTbaC+TSy
mMXNjTcZRTw6V13DQ0bm7G3ScCVvJcRe6ub2l9ttCblCBcm1hC7iPNlMTe2IncX/
75A1k3rF/WVSaB9hIhsVpz0VuU8MNi3QD2yNDINrfxrT92O5kyC4e1OapTS8tUMs
/tIcKQ2C9cZ0GEdyjyKHy7IBL9lL68Xz1e0TgH5sPRKyhgx0IKPRgpBc7G3dDAe8
pfZpYM87lbwCb/FXY+fXzJ719nSq7m5fpHVXtvWAf3q/HWewl4B+QmjuP7KBbCsc
LQWN9oz3JK96SB2frsYE0SMkYV9qUfVNWFCCCvf6RpmDSSXOP0aVOLReOkM3fSC2
ONAlme2FsDrLah9FfHkLjxqEJNtD+FV806SfHArGr+RQlS9lWZycMhKQMoCDBnky
5YkXR7iYxLRAcnvy42pgPc6f79YkhUuD4J4iMWeq8QNxLTZXKE08V8m5WtbUNQ/I
T9LQM7zE5DQgKr5hH4eYqXNthCNlH7cDRPUmeLUCExasD6DmtnS+YwnfjfwGA64X
hnLsFwJYvq9eqGNtRZvul92Z1kXjFbF+sZE/EF+729WrZMAcC2/RE+5qpMIhawzC
qk2mW4YlLQuwDS4tw5wZUD6jjvG8Gee5Hm+6cjp2Pkw2DPWb6K18ph2YH+iAVnOR
4ITkFKJ4xSPAr4YrR4sspI04jMNKTi88eMC0KG4JIKzjHRjsPdmtwTD5bjoyUrPZ
1qdOZw/WXl09ipOmIPuXG7IrsUBrho/tYlSqhSAiGNrDHmylOqfcu8N6B4H+3Tzi
rtTzdonc04rY+EWCHK1q6TcdJv0M1MtsCm6VzmFg3Icx61tMqFTNMcMnkQ+NMscm
2Hzc4Mk8/dknVZAWDp4kQRKQBYaabR5vuSQ2pLjMd7s+//Zd4PjOFDBQM2FKn5bR
u91ujJfH9dkOZl2TbsSoUuF1GV37Sg5ToK457PnD/VERHwYYISyF4Ey5D/Y29ZdU
rHnFd5BSVdgS7Ty8TFwl8tiIZKjS21yeyZNscCX+7Y2FS/wd81yEHBN6/AvPQkC3
a+McXPmQne11LeVJKfFu9kcWiT/CsBDqrvCANaNwUQ+vkYtZQorsitb7LdsDjJo2
jlK0kRkH9KWs56Ejwo4AmFyDadkfy+R5sBoFr4JgavQQszYb1mp5FgtJKSjubQGN
DwyMy+inyH6gqJYSKZ1TyucqaXK4R/7Zt5riTkz+O07xLXmGxoiOc2SY+h4vgdkq
JyvIjjMkpdhb6qljnA4t6vtNSjzgll3ztZqHD7uoRj5bxEGeJIYT292CmkJOIhAp
8Dh9BzeA3REZk1gv54nkQ7S/QMy6E2YcObA+scDQe7jT6gDWEiSWZy2RenmzH3gP
vTSF4dOx9XCVUSe9W8cICQPgvQ6ZE75V7SCvkTp+6HJkr4qmXjp+yIsugJnhNpVC
0vnbRMgmkckcp5PqpGbSvDia5T/Yh5kpNcg9bXE7VuaxUBz+/7qJiPgFEhy69u01
jqXaBx97v2Dyk4ZV9YkT3WlY9OpGOAo0izWvl4GntD7ryFnNdf+j0nXBRzxL2g8a
NT9RtOu3skLPbFNN+CT75V/qvhIXZe23+2LHppIplRHY6UQUDltoDY3nYBu3XkB1
oVM1OJ1FyBS/zvqm9UPzNdVuFXBH5lJMf1r8QF0kLh215glbFJI5/hxpefOQQx41
Ec0eiQGYc8c+Iv2bAhHw59KJqCzqfBUJPiZOT0bYo7/sPQPWHiLH/NqtenltGEuy
6eB2N90gvPzsoECWP1JFSavKPK5Z7y3HWFwUoZwbkDtCMLbk+U5M9nKGqZbEp9Q9
ufi96T0HJ6HqxBsPK0Gng0Q20QFPnlOn/SFIpOFIUgr/rVtdoClWTX0iU9vjKX/N
pfBYgWkA+oKRnUWjl4QX9xv3bHxxgP4P3kv01znfmQPqYFQZpOrYFk5dCK857YE6
tVJ0Xk/WJ8mlKVBFDT02TEsg4jCE1wPOcKN/xnOLhenRYxcwwe29Edk4g0fjcdHF
E2B4HQ78hCo2zSVBtcwVOjMl6AXrvzKDjNCJ5dGke4K+9FqBZ2YUvp6F8Nwi8VCJ
VS5Kfm1/WrhzOM88MP9pWH3TiAMK1jT/nyLtLvXIWAtp8pHMQCYPEEyFs2fwJiRH
6Wv8zvhs4NgbbeRPBJtyiU3SzjZJ924pjGB11U3yC6MYclKfe7BTu4dYdRPudqrn
kz3W4nvYL7Ecdf9ulYKRUt+MA2h75I6IWWvXqNtaAp1/zQwo1s4tv6XhvTXZ+z8m
gsqRT6eHyOgY48VdjTY0xlw+spXvjPFVHdvBIGG23HAzpHWi8YGoNiwkBrWY9t2h
BgfA99SxiSKhPOG4Uh3G3wduyXr0IMnuYE/7aTVizAiLyx/rx9s6xLT+F1V51zC9
RdzM3gFmSyh70OsuwX9m8xmrLh5GSGyzzPnycobUd8F/uBSnwhlKQ9GFv+jzPdhj
0L4BJ8h/NJxAiRHoSvnVZliQNnaEsRjyd9QnamgemAU7p8yohCToLa3Jc5F7lJpJ
szjYH9yecDqcBE3TUhn9OaLXuQi8a5jHZAT1FbabvjjFQh9nmyO56vvbinQg7FkV
J3NNBUW4gPUCLGP/oyrAyBTfMQ0E2hMbYgXADJH6vNn1sT3daS0gbc8HzhYJRLNZ
XHC2BjzmWI70odeU8utpa5tRRy0PbaqRHn5aUTIC3vMpGPQlWQkhWIdfXU94yF2/
4LZoqXdEOvTrASmhd55gJ8kFdxRhboJaHAl+A3caSeYDHb6/xoJgdn8N4hBGwioN
FpN5BDwv96VDEPrAZ9ditRf0ziihqcUH0eA+yA1e7ahtjYA5oH0U7Sy2yq4N86IG
o7B0tou61+A8weYVnlxIeniv8V94rHvgNHzrq9deRB8bz5m6px3Kp97AZzYTPmZc
I59qKGshRWoL2jPmPtARF2DxfkqNvbpX+63SGN4p/XK5FpQB8KuoV7yme9gTgLGF
XMs/S6Zx7nNrK+JCr3vxgRc3cAl4wCTDRTwkyeX/nxR2zlql7i5z20fPcSTQbnkt
gWlgaB4J7ux4aT4d9QBuRElhS8zxIXefwoHDOoezF/Gdik6wdYI4wjs5WUuw2R5i
vHWdht274Ad9BAQjYx/9W3QuZXilPYzb1u60PEXvRhJ7Wdv7cB04EUeRnot/9D8E
QG969Lcz1qmqOQywUEHMfkGXcA4UyvP5LCMY3mkzmiVe0IBtejjauss7nMJOwDYs
1n209sxWkjDc0DKCSa+01SYHqvR6cYR86ZSYWPOkGpgFZ86CJh6xrVyNE1DtmJgI
nLdIcy6d37hpLktX9vZPHjAwJESGJAPMuNxQ8aB/4UosQomIcaTJAuDWVxZ/98lX
C1unJaW8O+gmGhKLEMNJQZ1tB+XUaDhPsV/P0N+qnl11KI/qxWc+ItHVzYIkxozJ
VClvG2WXIWUeBrBLCmGz15K//aBF5NKDDNZk9FOzlQIY/WPOKEMI0joYItkz8jt4
96TVOUFbnwXLizmSldeo0K0dCFXkrwMvUw3aB5c2KsCJjlo4HkOOLH5Zke3zZyC4
T8xNmG3XWeD+egRuG7b//hcOedu8mK92S4s7rLsxUD0AfsCfd/9kQqeOdTASAXYZ
mBuOUWrXkOes07lONUC9mTnlm1iD24KnlvkplCr1MYZb6rfOhFrUnbQdyE70Jpht
3jvQBmgUwlyT9j52zr21cdAwihjo3KbXLDH/v7jXDmlGSIqphtfq9F72Vzc0fy++
x5zvxLbm+lmxITjwCkSGzb1qopfGUmr4vzRePpfOC0cmMNnGgmMHQ0zCfv/Q1e+7
6W1PXU4b4cay+oEyx1j2guVBb9cbXtE8nYRFIhUK7wC9DR1jvz/8+cLN1OG1E2re
TX7YqsGu4BJkiq6E061sOtFAfwtkjxFaw9QW1Ikc1ZQUVFdrsTiKu9pOHR4WtOXz
rFvwGh3vjUC9FRx2iyPOmGwJc2zkZfFvBmNR6/OiQQelHJxoCHQu6xAVh36cvk/C
irXjZ7/+JRTI7uhVQF0Ke2wb7VnC3IPidkdbo4Ug39cqA7pZvN/c9tKa96hpY2u9
DCv8x4NrSOV5rrALG46aRVOt650mpcSy6qay8yCMeGEgxAzm38DIRdhkqxKiurX5
WIAqg/7g5FDu/fhFJAoKqUtDX80utPQpbssnJEWvk+s2HxCwFAVUKRCHOdg94Zq0
HzMtEDx9LC0DZuo4m3MKh6ppUOGUU0K187MpQRzeSOO5YDKVDbB/sKJcevFvxAMu
m8ElTkisv5hr2ieoRRZ+ZGyvXKNHiry04hpor3QFe/EamPmo52x9RNgB5AFMej2C
Se7dq/ZSulWbQvlaJm7e0yDTBqIwmswtBLBsMmClj4GH53qtsBsJMroY7HzIfMer
LKDIkJ2NvJr/b2EXPMVdZs1Wn4c84hB4SIr6Ro6I7gFDwvCp26o3pYJLyJm9NlKI
05uP7RKG8L+7wjMs5wz2C4Tuw8Ovap0rNbVnz1IDR9/awE86wW/tnk7Dr8CrvUdu
jxIrdIbUfn03k8yOIc+pFmkwVNfY1zuWX0p3DawLgkuKg56IAWeK6icwauAvNLFg
Kg/gytpytdFQmz575hs6LBX6po3olWA3VsGzk98HUp+FtHPXkX448wCME/s+a/2D
xbvWJpX2rNrSR47Ww8ioSKJ8uZccweV3VpiamqsVseRursKXfrIMK4e3Uf4BDkiM
DghQ0bJM9/soAUXjfi2SnFxaBPqK/RrNHcCoaSiofXWU4xitfCTG2ti7L29DPQWn
h8onY1P1Qo+CWvpNqqKPluSCTbIxH68pF4WTdlulYfaY0ck1BsvlOKXfNRrwqJCy
C/94Q1z/G0ihlgpJcYj8g9D12CzOzIoiUG1WYbp/gfSSHZq+DqJdA3FlVQrUbm+O
53sx84IZqbocW/ZjrlQei748rXpPdr6W7q7MGUi5D/Qa2o2j1wGy550H09XsO4ow
fxIYMQTiLHnqvx77r7PvNSRkOPq7PXkHA2MPfqI8/6syruBY/AFXqgI3RdHJD6ta
ROFxWcq3T3OYXh2aRMQkL4qTDVz4KXgC3svjQ0zFvjlODwCoUBfX9ALUacrRA5A+
vGpmjVxBn3XS31AXhBItUBXrX47Bg238lRjsxtcoIySPQilSGl9lQmsVxEFAvk7F
Z9ZnZhv6S4OoBx3GngyHT4tNkN/UvjSWkvNjwTeYs5/5aEbfn9DAy5y/6/ViASMS
sMZGWYBD5ZWscHoGWKI8fSM7slYImjeDkn1cjwVOUTN7uhIce5FLtr540uayax57
+SVt1ru44Cu+9TSaq2hHQcZZ4w7BnApNgZPFnxUajg37DzfFR1PVPI3hIw1nJ+a1
DseFWnAjQ/EWl/vooO5LUAOv6xa/geXtDd2R9VP7isN5teetM+lJuE7Wry8ouOon
VnEE4QZPkF7X11pga4qHW9zDDmNo+l7Mnb/nZLpT+9dNwV2X6wNQhTlwmGRQ4ovT
tff0SqVjmHIRfjefarhv2FhJmlA1JYEt7msXEnltI7xtAjabNvE9xP7ThnowBIyq
Fi3YunoUrIt3PJJS/wAvXKGYCgu/XkIiorHnRsZiVHsq9gtz9HAeXxJE5ci5C7M1
IT7oSzwQ98aVVbtv7GALrWiMOo+cvDxFUZLwwvTe7qKYPCIAtuP2najyHxHVyitr
t1zZSb3/ZaOmFTpq/ZeU9oKbk3qr/SwaUJohD49zVUcn0LRgPgGESur7n52Tjifr
LRkdjZUdXy16257evDb/TyoWGG0htL7YsRLzil3D7lbNbzurLRlYs/e0Q2PLEBkT
MnlRaFHg3mxfTVDDh0Gmqr4D2N9gDaSnb7L4dADPFCsth4or8GYhRLdVtpRr5ScN
Lz3IN4dHZ3AR0KrYinnpzoYN3YtkKWau6TPtlXtiZiDMdQs5NAKAGKjIVxyNWheG
fUH8tWx/sJGyL4+qrLPwsk3aYkPIiIOOYUOgUiL3Tij3s+fAzBGTBH842NKYfASd
ha1cnRgT1jAvmukWtH20ExDHK/Q3jZ45buVNeEX/MwmQjIJfZfPiN+0xm3lernD3
PwLCYJG90XdcmbvxS9BxO/K6Iys+3HAxLK6fESJKmXq27S5gnFZbI6+jPvObOnce
bVgCl08B0bdRwWWj6RM+JZKKasVPfFRQcfRQNjhCG5ZFMQbcjyd2Y+Japw7Xpiby
9G+o8kHzYmFQ8WQKsN+X1koUOYcXg9bloo9pmsYd05YRtlwgTGba51S2S6qx1z3y
lpLkZdQEnoOoPN2R9/DZbwyh7mtHVA+H+2kxHqj6bAPhzdIvbXm5+5dD1hvmgnlX
+cTpBI0bZbtXKDOwlCX+91WkhRa1PulMKrBgjCfhonOJ9nXqR1+Q6FrPn89e4kNf
NCmPXFM5Vch1nhcY+nfeaoqC+PIxGUdy8BHLx3jP/Ck1f9oWpiQfOqsjrYmS0MjP
7ydZUgo2kxmIKUlghH3q6mtkVjkkNWOZ1st9NqNZR18cw9FtlKIPNwFsfDHeLrcJ
dT/qQymbqJ8XHjySuBb73WBotyfVtdsPTYUMB6usbJPQ2A7Fn+uT5s3BGQf85uVa
/sMrKBrQswRy+MXy2uEPu5PtLM61/JEQOwEvNJ6LP5dm6WdAgHFp7Gyv8v9Uw2KT
N7q2PTU+x/r8/Ye0vjG2WpEEW/TmNyeY6K6Urp9c5eNMMcXnQMd6+hHzIkGtWMBY
cFQlyF5oHzVvZeyehimiwOL26BfYZZvftGOUC5rbtRw3QnLV0efXpZUeaok8ptyF
Alh9+WA9UJ4o5vy9cjlL3+MJVWOcINOyRftNoTzFvJnggiIk4HKpzPFhIkpRiayv
OSE2mVtDlZetKQ8+g2zWoftE8Z+Z93C9TWIqiZL3utOiXPjGt+2phQGrwgKA/6z/
oGv1urcGE3pTdO6poC2X/TOlKyiIt76hq4QJcE+XuOdXsjCraUYvdmjgDIby5r/W
GOCkKYl59mCVRZ3hvS83OGwjvOFVOjQU4+1K1d0XAhjQWwg+lFUtgpRXakabOwWv
EsVAKkW20VdR3UdEX0oGag5/ZimLBsOY6Cs+ccRLneYQQHoc+b7THuIaJgtuXo1B
7nplSMCKEwa4YuckIFu54vJE3o1omzRskOE0YeQKnk0v+6naxn8lxEReoxCTO6cg
IeBNks/ecvpj7vj5A77JZnV5YV2vwQvylJ7qap5w9dl5h5PhDQKg3CT5KMMO5hoi
EDX4cC+0zskYeZp8vMjVNAWRXVOwy6z78udxn6wEJ5izLYJgKweD3EFtYc3XDQ+U
FombFDKK464EpeSYgb+11xhYAd0bZBlq6sabz9JUiRJ+B9ITBBU3TL5eEsgG+9I9
RRXLrwo4P6dCzDqkRLhxLmpOqUoJSINtoNo50ed9VFMYvmoeq1uJto0QJmSj0DUH
QXCgzh8f7fOIgWdYZIpCOv9Hks0NM9T+N0ipYn2yIErcKE8txzkyPdpJJs3O8i1r
Zbsc64z2Sp6oULv8bjIOUMpAKFb0kHBMG02j9qF0JZxylDVKtAmgQB1lYd9KBClY
Encxi8fqrKmKmrsZOPgV1DFw5OC6bu1kfEgu38qxh1CEczq9+L5OTctvw2kIg4OR
l/A9Pvwvx+l+hAd8MeunYtMZwC32ikZbMXMsiNaUKsEzxhc9kSe1bXSGZE2Xhnuk
zOrFYtg3eTWrDlyoXwANKJ10ktqEhpsuKtn/RTbPQcDDr4mcl0pGu2uAGfepWu65
1G/X7YmIBsolAJIVIfGrSmitMEMS2+MtUkv+ErvpbmpVU1DDNXTGynrYlstPa89K
tQDHoWfcBgunNU7G8ygMV+EHyvXghfOD4bS7GEM5YG88c+VXDh/P93ddIkwJm/zE
5DGqurpoQXYNkT5oETiJzqE6uGONq/g8q13dDootleXJfKCHAffe9pT/aBdQayry
NFcA7fAtAZW+R496Vr8s7h4npwrygQBlFtTCniiGA5aY06M6/QY3XYkNWzelvbB7
ju0/LQcJcM2SDdT/zqVnQQHauWggFOaV6+kwxIgtH+zFfGIq6seBnFtsL5l9Xo3X
G5ox0dyuUl/9uARIFy4uheVqkgCxrIkbtt247UyE7RjOiKPxcPOuTl+uC9p/6rHj
wTha2fBhbPOytIC3ZVAjJwusw66mK6vkskXcd1Qq7dNUSXl6ewP7oxyuNvGKX8Hl
XCF00i5x823egGEnrip0pS6V4vj8wdWFPkHaesK++2D5TpurrF9cm5DFhUV0zxnZ
4UUGe1Qx+9d+rUJSI/QhwQE5NzEH71sPYH8bp3OA3XTFMMNpI4ueHvA1MvrLFGDi
aBy4F/enln/olTsWEV6KzrBjmLBQxNTn9D+ncMV7QHZzw/kngbrSbYCABGYusLS/
Eg6fwy9wgiWUdg8Uo2o9svQgSsDxEfYSk3aNZx18NAzO0X/9EkZ8wo5OulOTgmR1
WMKEibCyWoVVWhc4EcS/xVT8dUeWgFONjaiH0ZZOWFG16srWYnOnd2TEjDQZ/mMA
QU7TbeV8kd+fUy+H+nADCAyvY5HvcD2rfvWzwwzaiHBe/LMXSlcIZ1BkmMOgPjmm
MtwIeYUJLlm7yFvI6TJwk9w1XsrKWJZmXjJQ8SBln+7ygx9CmbtCvy9jqxnspA/I
v+uHy+Adu04GAw+dKFCR9JBcy0aB+7SzTvpxHgMrsYSdW65LTXmtuIbPcPzOAg4w
lKyd1CG6dF4ONvtgJj5FVUJmJD19/hLwNXosR8nzN8985ExtgQU7X7hh3og2XXnA
yKryhMUuneE5RX988ZEZdb5tNl+wa1T/Vbw3BGE9Ttjkkrur710/HueBd33P4NqU
9rHFRnky0ay+qKX/mjzOJ0lwhHJB1pssnmy+fnHSdvDeMnlohdykyWJ5rp4pu/LG
TmgzFfHkpPQCyOBs7hK2nh1QtgTTPgnahQNasq8cx1Q17bze/yS0I66lA7FO8t83
P9qb2VP10LV7WWZzcneWR2Aj1Ary27b0w1EZZR9lXwDUa/ncY6Viodeu/hRGOQtH
BDHNeu0GWCGKvsC8gIgFIZJ29/e0fuJG4rlBQbE5XTmi3MBkdXPJ2saS4esuhUeW
3JmUwKT3gJqSOyMXZEXAhGdFWhYRI0HJxVzxj5FF0WKzX2etI00OzlKeJcCry51N
E1pPhY4VYVBn97Jft04Ljg2gTB1vkT4d5yYjgpcBMRLktaUpm9kczYph8fYDzz7l
uduxbqwzwt6NDFgu3hTkPjab2kOX7n2GytGSb6B9pvLM1axgP8ehaPZNAvT5gLDm
zWf0UMCxZ87x1o4NXl1Iqo0tZm9vvaD/ZDzcvTYYoxp+tllgdoa4XmcXd4oMbYqu
hrvo+VOfbMhxvBPmzQecx503zAonlMRcYsnYoljLrSyTWal7mmFnQSHVhlGR/+wl
2yjrFmOrd6B4nm//kEbjU6WBR30Awf5yi7aHEe+wWjeXw1cM9FC1fvZQQ7DJB8h+
2YM3ZbrtY0dj652MkfcaGHchI4PY4UZ74ldCr7uOmsjPsu1ggOCoY1jCkyukPvAX
VhqYYuE/Ozy2rIthUZox6mK609XhPt4AB5j2sG5GJRyFOLGuPaExVxhePxnKUm/j
eaBn96csovr9WfmPiGq2MgdI8wB4EmsamDvFO7QElD9ooSkUtPeqDras0vt+nSCJ
d7bP9UAnpvCz1Ddr6Mub1kmex2ieQh8NJV7p7sMBNWxTco28BdpRWThQRCIazc05
UHAMbHYgkGmraj5n7tob0m9okjGDuja6mujf1Kw8dzbnGyEGLOEGuIPPtX9AlcI1
UxH3Lh56ma3OHh5Wviyg4YAoMJuNBbol+LZ0biPYNy3Mxm1KAvxO/Fj1zuo4BxMr
fiuQrqP1er4uAW/Wj+SOkEocfLQHpZD/h03ojgBaAXMPrUFLpo0XjCtEH85yigVR
ooMzGGc120nPw5PqsU6XfURmDMzpRI4nCyP6VitfRyFMDF/QJuCF0mhf369G1Hh3
31/5EX/VsOfol4bL4xyYWiG/QtlntfSl9dFZi7YO5CsS4pHOGRAmU1UHYaggWwAp
D7is03xRnPFu3P9e+yOPK/cMBXR+26emla13fGCHY8/8GUaClLgAHoq6iuyXo7R4
wt7BLMzloz66/1inn8qsxzLQ9Mt0Otx0aD4wrqsK0udw+R8lMVe3w/55UmPlyq9l
CBSsfEIL7PWJbjuTE5xaGxJlny+WAEWf5Af3iZnQo/w8Yd9VGqmt30XgZCyhVlkH
j/bZ+vK+Uu9sWltNW4fwqKLROZwl2BTzlXrToFIw67ggLA6fuYcLw2Uss3IJ0w1R
SFn6ufjiAndXR8OQcs/HSdRJEcJox/wqIEZ37LAWQkJ5Mb5D0KWYdofXAgHLLhxc
apE9CFFsdPazua171mKpyCX/VCRuqPMMy0eEej3WXCwlW16xtxMOCcXRXSnkDw2g
57fctn90Ne6cjYAMu9ZbEOTbk/pm6+TTREmAoml50XiAm0dYw3I3s1hIJNvvn6Pq
7WBut336nBhyJZ4W2rz8TrHfeMIY3K2IJy/HVex/YMDjYKojHfEsALdRvyammyLA
K6uGRNbnFhRC2J3us9n17UoXpCQB31Y5L27KhYM70B7qLjYvGN1oUoj+djEtoHmn
eN5vrjH/4Tzm71k++2DNbXrHiHDh3JYzITBHQZKBHEjvQHTdi1L/ghTJV5bKe66e
scCbhyABdLH4ombAp/d/wFg6Rce9fCJ2V6YYzYyFtVO+YMETYz8qtTcP2BFazy6h
A+2Imes5wHmRXtnITXqi0caW2XHnFviKZrBcG/hgLo/rLBygPQUSykQkkvcXk5jY
SHySFOw3zsWeuN8GLrhs+jMFOqoy8wnkZbP6mwF4b1RbuRLE4r+Oukgo8KQJ2AMb
vQyofC5cf7tl9DwTiMzSRMI9x391kKcK9k5wYe8QEg7eObzcKVAxyjrflPnobhi+
ZUOjFwnWyPRy6lZjKWuG+p8tnJTNgulbsUvLY9DrLeL4vtJFKJlctKQjAYDgTuN8
lFk2QXMSGPDwMpxTBZPrTKANg/u0sPa3sWh1j+dIeiBS9eOMXrdCU/tZa0kH2lvT
uBcBGUjOME9jzPFDYHsBoIoXDNFCLC+2iPwQ8WAQLsv+BWt8SrhFaFcehFjry3eq
qLyXxRyAC+SRv1Ml3I5ji7ukT0ySsRcFVE7DtnJVAq0s1mzSD6i1wIODM6d8XKfk
rgbV9QSgeuXbud4QcJVvRSJUmvTr+8ZnWAzCpzEQerkfFOLbGSbtOxxaln/X1OTX
AtmkW/kW908y7SpmNeNxbmYVZdIKGNNIR4zOrpEPEnRBC2JGR0mPma8baWS6g0SG
8CJm03uPsZDJNZhMUTWDv3N6FRbbgSOZEUpxT6nXHgMlogCRNKd4m7yYvUpB8S63
U8kPrmrjCx6GqNysdfxceHay3kAs4nuPEaWiI3xtYuJ8dHTtQasXTfS0/loULvYz
UlUCP5GXMfrYYkvHJEmddaEQhaAKRR6bbWwCsam4RhlCqMIdL/PnGZjiK0bqJGKL
giovqGY9nZOOOcB99Fc6FTvazOVLhOPEFIkIMhAm9Y3qo5JvZCePRc0V1Szew9vx
R5ONCnhoTT+8j/NIfEqjcGpHVgPTPew86445fLlMDo7J/dt20LClM7KtF+pbVUeJ
djbeQy6wqG4Xlyo/61qCubV70EjBq37yG2tgyrY1ltUG6a8m6aBQoT32d5BZSsHD
+CUGd08niC2WLfaHZGhvRIbjIeC/25F+Y7d6MkATjLhudP1hMOnPDxh4PDeNhsJt
p/J8u6aWjHGzNtWyVC4N7GTWK9BLV3m+rCBlCzvLJimY1M94/jYry8mqucq3c02q
DBlMHV/CcE/dnQIbR0AqZ5tDZJgN9jMgyI68qdrZ+WBpIztZ50ElORlxlGmEJvO9
ij96SN0mb2HxdmlnTTKx7usDTNc4aWgNkE69tCebiJGgN9H9sf9EZeM/GdBSu/pp
OUNW98ZrAWrFLMHIe27dZZxGr5lJjifjKT80kjWJvRz5JBDPxoGkqUJQJXToQKop
Twpk51t32pybBqbbve/J68ZEg5QqACvdsSdXiIHrXrlTDCtHC0LyYRHjzV5SuclV
4vZEXw4R/PrBDt36aPVKCKF5Ko9yct2ui49qJiuXbFjvvWdvIZBRdscrlSkj3TTr
JQm+bbaIkSm5LQYXwlf73lAlLd6x7fdeWeEzsCVNH++ePiqqNen+f5GDDThVw+Eb
t9341V3KbNpCyZZbZjIxpWXpg5vjVQZ9zdq84QE5VOxyv78xhg5dwoleaCZXZgqv
7Rgzi+q+zPWvi4QjTy6K/ELfB1d4ogp4gix2uGyuIFFv0+Kpm1c5iwdyji6yhryQ
2+ntpuWCS8JMi+9woOX92sSjm0Lr1bFIpvyNnwBXtk8p+trgLggzB6HHohDUDpUr
QwHmS8Wqs64lH8RYX5/MRGoq1vbLBxKvK24Xl6HuEQBll+h3U6xhUV209Yl9c9Ss
Z8IAzhXd+kaZQopvCKiCgLr+ckwpKZADvXhF5yl1s7/DR9jPKV0HkugFJBBLkmX6
cjDvzuZ76QoLQVNWp9VYVmowDvS3zFubq3KrvQgt/W+3UFhJu3x+oIXG7GMjA+t8
TJnQnYDxIOI579n/ze/bLqPIUVvrYiqgqTJBppJgLHxMq4XqbTKH2kykdgTPBqJM
bY39v8a7KxuQtJR6QsUiAZZ0hu4A2IB1S715Q21fof3Tg/WuVSpZT7BT7r0Y2sT5
lmFPgFHOIa9CuEqxpQ4BIx7D+7dz5DdU2p/v6Jv2PPycqO/sl6LM/E9eaHfJl/qp
dhts0UKPe8I4VO09h59SYjCWqzmfgCZLNPHNHAp/8pyrAb1UF1SUpBkDhcItgXqA
7eNa/ESDtpuXzKMbsJJxSVLttoFZh5ADs88oeJrFDpWEr15+IpoWq259hEO/0Pqj
0UK/cNatl9BL7iIusTGXj5unsPDTQELAxkDY6RaKSV1BhCi4DWc+w2+Hf+xGm3wI
qgXNmU/vG45A+4SraMp+n+02YsHeQ6QaGfFVAapbTHd8trgNX1sBbVP6gQNKLGxS
vXJQ6xyl+FCWkmeA0B1B9Ev+rCa5edfpXcZOXaUDJDRFmiaqlBSD1VDfdldRK4wd
MhpTI+S6Wytz5HwNPzI9QgWgg2m+1nUrAEipEOaWyktYfFPX23v2jpwwvL3I0aOa
C3mYruUq5Voh9KxXt0copOAll5xjAd0b1pksES3du1PVCKwGZ1DzttJUj9OTHOvY
lLbuzg5BMgdehIIyhQFTRI3I/SgmAHzhpCmVPQE1vcYfPZAnu8jJFmKXzgIDdF4e
LPytLs2Jtu48T6EgTAOq2LTyXLPt2NSJWIscT236W4W0TUX/CE3dNmt/fRolU22H
7BaN+KBqt5MeFhYz5OcQJGvd0Lysxq33c78fK0yI66E4ghVC5rL9L3DKkoWYa2Ho
6THMdsm51AChI/svvHHniaHOjuwu9W7ogIpAFci1oTuqUbj2BiOQHLf1iohz/hlP
SsVKQsDMsfFL6AbBBkWoZX01zVad6NA+ojLQQ32YoWjlTb6yIHmkd6zBf2hupeyK
/IEXblo9KgCoVqfh1CrVmoyVwE1JFZWXymY9D4PbHesg7hvsFXAcqDf+iUXGMddi
QtQvGaiyYYNVxRhd9qgJS6xpo7ScuoUGLEjWGSMbF36uZWj3acutkQG7KVIV+/kB
EEYZV7VS2/LOwtMYnNWISxfkB/gmZ9XVEQP4WacaFvgIrb+X8g1CQmCEcayZxELj
zdNugOZg9qleTkVyEKxW1U/RHmGY9z91ae/gZpTMybBXCWPVbft4uhlOuzlyFNia
FE/M7n6BIEG3R3vwXFM5wWW6BqWkCcQXoyIXU66e0iem63c38f93cQX5JDkyHadh
lmYYUajJXGCj4ufPCGZ86KN9b1qc20imXG0IUcXR7Poo1yk0nlM/9/ucrghGh8z/
nQnjVUAwEDIxHr/1zFKgGQVWWSIrpMMQ5UeL7TOmrFgmsMLvETEGpnpYIUCkTbgM
3LyBQbqXzIaRAm5tT+5fsEAE1fV1MagR7gGclso3CXGvPewFz/yD4OcRxTpZNkiT
haO79ztGXcWgDQ8dYFrvJ/cI1v5TB5kbXgwTooNeLxcGJcXjHgfAYcDuLgyU4YX6
qwL8cKLkwDJZediuRoS3LWc9T6Uir36ftQvcey3/bR1gx2bx4XdROHeJwN7G3rOl
ep+K2xCEJOdggmM/N3ttRIW3eU6hYETAWsS8bKStoY6a4UQoRp9YYFXVJLmsHHPH
+tLmTakewlBJGaYCGRRMK9ch3deHSdoX6GEd+D6gaqFBvxsBmhV7hvR4YIpW2mXC
GUTAXsLG4XAws9ARsoHzVp18xALKbUcRYgY9/O1gBqbhpVv+CAEUq7O0TmWzNthO
FhwB8m51G3BJ69gha7SwKy1oaRG/YhDnGJr2TvXWy0sXcG9QYhL68bL/XoZE7OLa
PeKN+J4WOzx8fbcbTTLYspbYAsu4iqEALb1e+PqmzYKjPPwU3bW6OqIxC5cFKwCQ
UBXWPSPiRFoIbLytjfQNqdIy7NYL9p4S3uG8L+/R/KNXEvUxLD+DxgCw17EscZcj
njBlNoxwBPvflVeNEbpI0XfrQ2WUv3aZYZFlLeTAzyEW+fqnZ0edpyzer3amE81u
uJwaqOTfQI+TUc+6UmIRIXGiXzIgKqEg5JI/H+pjBvEu/cEmmBD9Q2zNyXmdA5QT
WXMAbWWkPR/kUphXuuLrIZ8uamCfWjWL7IuDpIqwJKXd/ctqsb2ITFbU+WHfB9bd
Mwz1Wdle5G6Lt22yDLG3PAtjAoMKv0lpWC+oqt9ynbara13rmNT6G0fLZAm5UPHF
8Dp9KJP/aApoNA2KsKNrM6Kcef5zEeTOj+TEuvwR3bMt+UFFbHjVmZXP1SSsPDoZ
9TmWdvSQfrmKcFUyb+rdeaQZR8jjrg5m7aEOZ0ujt9bdeVuCR06YphzEsP7CQJ1i
le9KLnnNXKpUnUmt9pgRoTdYEu+gscL6c+q87aik0uQPXVVT5jaFt7Qza1OmT3Ni
OtgTReNVIIhYM9/i7X7/sPQC/ELT+XpQGSh6wEYIvvlrP3Badw+hAzJYaOBS3n56
jjWxx3PDA9tMbxm7iI98Nneq6qrHF28x95fHzCpVD4Yi/17jitGFQfIrWYchGzMH
DB4fuD1Fg45c7VxYSFC4xVBT0CjjfMkqgXSBfBtg9ypRNJFvcROTBI2qSBE0TPSP
q9niYCbpuFeZKIpFK8mhM9i8DcAEj3BKCmJ7oxFpDJJvp5qoJOb7phF3K4BZLKlH
PiVl3KBvDuMcs4GqsGN0rmGJF1YvzCsWetoas90X6RCJ+uCWpaTASyCL7In18C4Q
oZo6ghr/9YJ7ReE5wF0hcXm3aFAgTf1AWKtUlax2QKwKzrc/dVXEq9jgOguZYJNI
gJyHWT7Sls/CROXmGRn9ka6rReKXeG1IJFDDRdaWDKDG3dbbhHxbk9QrlC8+i1uq
TKFGgUXNRUFhxHIOYYg45dHEIFRwYOkY+tEc3XP42RiOD8w4QKgknorDtvDEgyht
v9P97Mvwa+cAstFs9336vUrd7E1ZMqnXIvE9CqvrEzaxs+6MErAmr2wUYDf1imbo
DSweghoNQi5HexjqnU0zSrgaXW7OXPz6exEfiXq8UNKt5UU6+WoIVnau7iN3lXx0
ECjVigC/JUN+F/UCWeUyg2etGrhpYyU0Ok5xmovuOQJVKbLmHd3imTC2HjdVhcFQ
ibC96KciRySjr0c6gdllmzjVDYQsJcD7q9RvUALFcctXlbOXlhomvfV+KdhIAdfh
RdM6jT5Kbba6/x/6y7RLEyIvqh47ZtxlMYx/RQgllIAQwJzmXfhx21tHWcMF4qhu
QFoy8kH87hZ1WpSG6uZXs4BeuiM/AEGYYa2celWEp1qqdAfdILmhUEgRmV+txe+b
CBBDPynp9azj08pCM9Z37qE7a/HSqujyAxD5uq9+xwRp/3nXWu3VdIuRkfBvfudA
9VkzDgLEedE/QgLMuxuk2nNdya06zeALyniBrJRda/xazvKcm9+wDihqe8/PkiUR
kVn5DTcMlvaxlAKweJ55MSdotDzLoWr0UCpZk/Hz0OrDbDof818S8FDMneBqipE5
meOJ0v7zBefGromeNsHGXWaM8Fmjt+LG6pwcfC3e7oZHOt7UPzNPhax4h34oS2jj
y80xLgiVwvTCojLnCSMj/3DPiLo5jnZsoZTJKdGYoe3S8nowyXn3KKiKg3HRz4IS
bjqFTyY7/g5souDuqk6f7Je4sSpGewjVilUMc5ZJUlpE1YmdUI/1MvQVu9F9TEqy
gBCivCMVCrIdfA5u3qk+U/+n1u39Q5WEWFArWztquVp3cccNOMk0DUEfAIg3LFnp
oojLMLdH98rkCeNTq+sXxoo/zsQyHKlh5Y1VxIFyIXSJM8ROfvI40cG4OMUJBnXm
IsgdFEyiBabVvz+l5+KKKj86VqoQxsi3sh5ZFG0hNXo73SnznK9Uav9lm2kGMAOl
LkhPzCFM3VfAEOyKWTvZJcq3YSBZ/friaebpP1Jw2lNPKOKZYWXmMluXvu3/bNOK
DAnCi+djF0nmhDYh6yQbjVIJw8pLF5MKsfsWHfkUTWSmR4y8Ahr2ImglaKSKgaqv
AQLAyNcZqIc1uDwG9AnQF+OJ3/6WvcZLnS3Mq1yEZTtmpfJ6rjHOxBrSMpDnohAm
EObCikB5SJsWqu6poGRiu1i3y1KseCqItWmyPOtQi5ie/g/ZHh+NiCDSfMX4SSv1
6+5p/+Smd+Zwr+fdstKVwhAiDpTqP+KfnhmHp824WBixgR+UDbfERLDJ0Gipej7Y
4Lzj9S3TOTE/5XfWHKHe4nMHcKLPA4T85Av27Bbxg3j9SNa1mLgnVzU2pdiJpBWu
ZwbPKSndZO90Q41W4tFa5YqswNPKWyl6dIxf2+rVz4r/BeEtztHGaIFQMCu5sKEf
MZl29VQtyacjodm+lETM1NrmAmVGYPDsjLPwpTgvdMkmqatVjnU9MZZvUpDX4/4q
pMjTO3KlJR7F4cLD98TvWN3k2G0jox9PjC/Gf78goGx65/qCmQhswNxc/PI53Q53
EFNeHfwTl2njQ6/CD6deGKiIi7LuzcqjgKFhhIdt0bYQQm3LHX48jemEq2HbNAF5
vanje3PmukZKO1qSzIGdAlBB2NIK6uqLLglMQcSU3frz2wZ+6R9PKhqWb2Nm+IVc
HswZ0+2qhQgGY5DHBBWgs7ASsf0qLgeJ/7IjyQ5Sm4YUpCNRLHsRz5FaXwjNqh0J
z8tZkTGm6frxiQBuw7FRsQzCaEqWRLWSrebpQn87XppvA6VWG4op3VI1hRTgU176
Jt2K993GQ9pePcb3/dmX5T4QJ65Z4A9fxW79IHSvfguDmJwNVXCPlnIRGcSTMunR
rL450uivmcowOk0iZbazZwiBGQMgx4a1gRDIlwlI/m1iTrG2OE4aYd5QwoWjH9gC
c+/IQHdWiNRwDsWsvPvJ0gOag+uCXdQ/r/J/Vi+STACXXz9bCXP0vNwIiLiLwU1b
q0vvhXTIR2H4tTyx0OKnuIqVWNzoyi+TRZ1ovCaV0r1ma00HG75guenXjvaejUHL
nd+0ioOJvPPe1KFqdSFTBc5kKdXjGvoZpxEMsAvW5KfIPdb+wfopsFXycsEW2rx4
5blWlUzGU/90aSOsJezYlradyAW522KtEpZOzIaDpCsu/D61/RIGxcC81nX8DUs8
sIHrOP0DQ20u8A9xZ6PPz0VPIFWyGdNCVisW4E3Sm/XVPCMNzQmgTCRLjxGamehI
NtVGjQUw5RJhfUxyNxkoHQVq07kkZUmMkuDCRFLIN27vB8gZDRSgMnVUlSJa3Cfk
smHUNmpNJ0FdKlYwZynOdrs3UrO67ntRq7GtZk+fRxFW0K18mTXCAJjy84vhXIO0
qroOGbSmuRiXiMiReZeXBJua8n370WlnSmjH4ewfath8KPcgFF13hVYKl9JV3Anz
hZWJIFqLn5QMN1Y4587z+bUHvh0AYvywBeqEJAerui1YcPaikZ0P5z7Jyzr9UeQp
3nokN7hSZaaNDYysPcWGYlkom3lk0eAQEFvkPNZXf6FQIoodZhtXZTRxFlIl2JZB
V/oMSaifW68ZLPnkXj0IuT71padxkSHB60iK0m5IbVQ+wZrr9zFZOej7VEgS1bb/
NDhfuc+WG5MWzsS2n7yTnmLCxQ8eqsIZ4W48PVmofPil7k98A3C9IVVv1q95QUNZ
V2RGQ2t7pgQXUb3R1quZV8g/5rcgK9dY4Yul3MXzLul6IF79NXokge7plCEoqHly
QXz9Rj5cNLLa/2Eerk85uUBUkzDVG/WIapfeIjfdgjKaMwB0L2acGeLZnnGrPEKv
rSpIqLl1cjeVFK0+LfWY0o84kYNUoJNb79tU3PXoUnSyLsN/oAwzAZx+2E6oLrwU
bbroYKTwnak1b9Xg8goBnSRo1Jgx1sybpoVwS77MkPAu99FWZFKgLwPO0LrarOVq
hKyU9I65bLR6yh2+ybFVC0tbZ965UKthB7SeNx+8aL+z3OYLsgJ2Si1vzC0C1SKE
+/KraT8VyJHIkmD2qyeT60Hx62eS4Tu/XWLAluJ4oPZ+uAB/JDRAbDoUztjLQ2cV
pi7b3UVvQYirnnsJTPdWrFRxjlwK50vYaNpDOs/aA5uebLUKGdeKJ1utPhHYxgGh
J2Te0cse34BAVTD46MyihM1qwgR+PzoP3A0q3W9mnoU6TGkG6GO3zX9lKKkA2SO5
NmvxVRjCbnA1qgd5n5OHrL61TDgx8MZRnWH1XwGIy78eIN8BoMjVI+/gUCt255yF
wEdJJCOzhZMnMIWZoP1OrhR4tiiQ+9NAC181il4xlDo4rFkgm2hLISe6o8RhPc0R
0+tIrGjwos6mlf79ng4COcZnkfLjqZYZYn2mPQkD6DAunvjaR8Nj0BF7+VHwHYll
YdJB69o2Ian37iHOykhhBdNIETz001+cLBpFlm4k4RTr7wzf5EKMGsmkBkNxn5iP
ULZZZLLjVljDVQLToHn6MNkPq55RCqyr9vy38IbnMIUWUyun5k4YQVvXJ0MPkQ+w
87PenjohWH+4XjpUGAZFaJg16SsWm7dkPI9F9JJCklnn9c6EnK4olMdiFbeHz3WT
LzJkHklThIJEBE8DgJ8rnbuuo/f/mkzu6ZQCjJRfLAlWsHxxFrPgvwzA0fNxnfc9
P7cgctYm6YU9Tejk4LEXWdRrDiBY6q0rjn6zyAJZXDzHIxJBso2aACwOzjef/yaA
2oFEpM6eVmUZsqSXKcmbSguxxz76LyyRjM+tf4yN4kNRNdvO65qthXSj+K9Hucog
4p5J9hq6X46MuhcuaHfqjHSuWTe7yEw/M79fewBBdoU89spogbC9caifrcecDetf
dtSLCDW+SYbIZ9VyZkoJf2RCyj9f85UzvJ7kavXIemX9nJHl41b3yHHjXFf5egQF
+8oDEi9z2kteAhgCAGKOP4hOUHonf8igSEWzljo0V/71vS0x1BAm2S8GKleRI3aY
PXYt9lrJu12kvStqvNVQseigRpJfsIE0TNdKOBa2dtVEQRpHNFYrUjOkZ2V5mOOq
QxePTVrHeBB4K9SBxWah0xiuFAaRFxTK6z/BTJIhemAdWxMsP9G/SkeNJPixIFdi
SM1EtcdrYTvZSMtKKMpczfEsO3Kg3+idGw959AGWt04P/7KXWewJrCXh4h6VT3RY
fNoLmYJJL6WxhjzTk5B5dzndv1A8aENNmu1doMkaBFHhQ92sQbgF4KjYxJOQsHtg
wU6Otq5IoWrrDUTy1EnuHgVQPgQZk/WWFtHPaoRAiFV/MuAkx1tascrOaO9uIUgc
/cqyf5ILVY2v2/p+UW4qQNJohcZM0Vsqcvar/1UMeKmJYxw4OQOIrwyQwz41oVp9
aGtGoKiqEhwusMXLfdM+9Dj/PjfLEip9bTJLjDOFh3G5o6mv4YlPXTOJb/H6EK9R
+/oY4VGwxUWyP+lNrkPJ+AMCt+WD/Nd/2HLTOrIlWMWh0ylkrpx5anlKRVi0rZvG
t8DSZtF509Gm3+SjonWeNvpjCkGc/sfgE8URQvmUTwxS04QRL+fPXciO8Htsgb5J
46kS4yPsy0F5Ks+SJH4mLQfSw5GecCZpaAKOtLi8MArO6UHb7TzD2bJYSpxNyfaa
76DdtoMnyFKgeoT0CIIV82fYadIbHi16ae2kBaNhk9JC3a+xDzbYZH/RegMZ5AQz
AEDFW1y7cUSaSg59IJ7qKcnkEw6zhga6xZvAe1NPjN6c/AjiBNhltXCTdla+xiSA
hBqUOIqTQvNFJ6Cx9zc9sahQwLwbcDFP/lRq5nUAhJfhyts1fkE9V8wHSvq0c4/6
N8/8+acBbv1etEj0DZnItbhGeCbbpDtMMsE7uFLqDnmvwg2OAzRTDdlkM3wmIP3s
Tnf8PgaO8ossj0rnWapqkfnYWihldwAi4HZ6dk0ybhqblnWJEalw7161kh+L5pYE
p2Ij7lCXn2v7EasV0Wi6jlfOJaVgsOzvNXRjTx3nd1We2vqSF2vXImUCv+H97qnh
Rly04M6pb5wBX72GtQZJ7x9fJbjrEN1WjTS9EuxXvlPEhnUtduYzpWOAFiEII+9l
bQDZZXRN8hIP5iDo6WnSDDdjV6cgzRX/lJg83RklG8WvYfXFy58Jj/Hp3HD9zJ9T
khF7YWrNcQ/5zZ+njSlP9tTxVSpEGKLp2WFn2RV1C7WkzmmFB8AULN6WW1DsTN2C
sHUiMEr5K4RUb/OxoECRFqZigxmNONcU7fi6ri9+Hazc9Cn6p6MB+MtsHoohcp6W
pI2nyGO0DM2NFk9B5ZFIXceJGxrlGJexo6IBSXBXhKAx32xJ+C+k3tbLeBvnSjhB
aRIl1aSh2+LuKKdUWnQGKuEd5Vz8ph9nBZIygVte5V+nhjNrb7k3xW+qMlBg+kcl
L0tadV3z6X20lGFXQMRbMpenIjztje+Ul0EQMhrqyLp18rwcSZOwK1/zUzeQStqh
yfoZV40uWbLA9uDL/VFyyY+Qcs+F9KDX6eFlacJjurlPET+El5cpA5c1x+YWRtQ7
TDIyATCqswn2WTcfoEZDeI5pJImxxn3SZg1R+dmNM8QFLpByPRqo2J25dzb/c3EK
QrL1yVWvhnDYPbbMmY5dqOH9KrvLauCQcL3YMzhuHjSkyPf2VY0RFEzH43YzG45e
P5KaExf2JXE62gQmoW6LUJJrgbWnCqPYfPyYbw3pjKIqesOV9EhftWXOzm/srnB6
pw3ykDeQiPFrfKQJxGQVdBB0pSoaHc73Zz8XDLN3zvCNsl3YecABJijpTbxR71AD
o/QO05eOCtD1o/MY3Wb152pyFuhspKR3p1jnE7+6fmyRE5+PMTd5s9ndpt9XkTH1
dzuxXQPiLgUaRK+tOgbmGZpqHkSeg65wN5WqJp76PxYTcQBrDTqMnLx+F10kRwaZ
2iSxL4rNuCfnuPDiiFcC6ogoCA+L3NOk3R7JGw3KFUk34Uhs8iSiSn0+ROiJ4SWY
5u0/Y2Cv2W5wOfl0FnJrSbauWAQgA6EEGwmbrv1P5xdTRbMCDBkF479/J/pD8S5w
CP3+hKyBQ0xtz8o2A0P4DCMRRfMUKA7RTX5Rok/wI4P8BdEbQG5Oe1Aonbx0GgNI
FeFeINc8qtQxlcTfVKEHgdAne9DJa9NZOTu4pgcz4fwDAn6Cgtz1sLS3q+uE9oRY
FDTIprwciMFo1ITm+NGZvpm0RlrMnuvA4+RXYsckSL+/jFUcYCwmbUuGYtJT+w7H
1+uqVngN4YchROAtbvLLp4NbXVNNUdd/CUrVWVX21W36zKW1sZS2lrDUhQCW6g4i
nXea3k8h2pklQFORgbGvkZIgY4OzMIFDNjkC2bvYDIRkAS4hNon9IP1cqsJLo551
1PzxY9nhYtAJSd9lnbFngd2myQE9LoiVU2k6VFhnGqZ5gKrMVzgg7u/k+zPup0Zd
BSt9eBNRlvGE9kET04Z+xvxZb5R/+mB7JBD3+Ezu4aQRU4xW+gSS3q6KxBrGiWL3
kRL4h5si9GoA2zBfYmnbvP6nNeNpEOHaFgJKWlK/RkUaAx0o7JSnj5uc5p65YJZt
y2u61dq9K1g/9FBgw5F3NHmyVGYD1sE9FrVYQt5IHcj2hAMGIoLKJSnrIDVnt6wt
tY3q5Pkqf2vHebSpp84fEakhvSwFZDEl4nxkaAz11g/f7IG+ZM3fwXbNitUP05Gh
ALnjOfo/rQQizpvfichupgvKzBJ4aHzgpeFtgHi9SiM8/kT8ezOcRmaomw1/H8Rv
/6E00Ppb1CzrGFMktENA0LnrKXOCaA4z/d72FXoaYzg0TTR4L7RP/iNNfx1mozMK
Ny7Bk7AvqKROWHLKnu+VoU2hvQopTPs8Sf3+XAlwc7j1633c1btht8vRFi7Jh0+o
FjfOlISZovDbUNHbFcpyA+oxdE7AB5rV2VnD0yZauN+gp5GZat5ZnabsYuP/Hl5s
JLN0As8h98IEHEjMOQSQv/lPTeIvK0upUxbfGvs+3TQNHLUKBKZDQEXbAQ+lszos
y9/nZ5h8y7QSpWl6BJbdoBNxsi8/BIlzYW+A0PacSq16tPR9Rzm10Am1Q2An9fFM
9jpJ7rIi+KrXKw4thYKso6c4Vge37maLAE4BlleFvM7qzCmlYmxdOoi0z8IigRdF
FMXJMD58EmqiO0YSkput5gjADCCpLL4/BIAmlw0D1mZ1GiVdAvV57mYd2qU/IcCv
73EtzygEWfR77K+ZQmhZdO9hGnDh7Hm6VHdYXmB7cXJAvZ+SlrqHWEwHiPjF1LCV
AIVyeWkeZ5pwUzhxw1DgdfDCWm3/7HUeR9jxwAIf7tXXcmx4GB5NQDXzjAYuGMvy
SnB31VWL+TA9bzrG5Gc16KFuIybljmtrrDDaWvOoTaeQ9zNQ3In19CqhLyhiVhZP
9TpQftQrwzOP74QrKmKd7h6VrjvB+7jxLTW727cKDNwFd2Ed2BUbgrGNylg43BKy
ZsSFtC60ULd8G+tz3X2gVRnBroAG+b4rakWLzKM0cI/5n4ZT162ohHXsq90maT2R
qRO7Mubl8Bo54ynLnARHXNauCQhw1OjcGoSl7baQtWW6Mr+iwwNk/SKIprYvGkQt
EZW3L+2rlv5P9kMD7ivfIyczT3LpNw/PdkKBsZepgnaTwi5dvDer5bNuco5L1BcT
2tfLGjTVWTYS2q5WaTYiQzIDXU/zJ95F0GINkW3tigbwkB+MAcuVIEO7Jtewg5OG
/S0b75qSPvmW92LMyid7w2yk1EY6I81UaeYUhWzPpbbatJofduGSAVxj6fwAkDN4
O2ZT8P98iemZQcB6BmfY4DbP/qLijANShy96wWl++k65I2+e9s1BGdRBA/8VnYVb
5uuy7tB+sr5/NPERVcCD60g1HoiaXlQgs8V/C5vkijY3v6ojzQvkt+d78K2imJ9X
duL4U1mxvvX39KhRFphbUiebP0jJD5S3HON+5mVy4ekWen1oQOYYVA5llMXCPEAS
FX5nyPgU8yXY+X1YUz7uqzLjMGKuNGYqq0Q5LqaCCkZH8Nba5AQ9/YibVvtoveoo
iSh4X9y//CWtKPzJLQ3gSmOu+wzUfF0ZNV5irAcxlnJO4Z29fdxlu85aBlzMciJZ
CwJtaPPOGIlvJTO48IU5tqL7zCCh7w2iyVENwz8eJJOdT8l+UKD+A4FXM5Mdrqzz
lulFyDr20FIN2fDnc5FCJMZprPNyuAuSDw8SrKOr0r5AGxDevH+PS8Hwz1WllnDo
glYfWhYp5ENONc5NzvmdP/BasTQNftMDuHRGrTqAbAUQBsSO8fd+bhSjJlb2abZk
IQOr410lxWLCTIVN06e8KBkeKV5bUyYGgqEdBQhhIeAjWR6B3Gf4UE+jg4aKIwZa
GZ7WaleeuoVIRUqo/qzBGKzLEWZ81fTOowd/N6ICI23pXykmD75zrFeXFrMaPDko
CApjqRM0Pfe08mJiYAdqupHWkJ8lYStc7VVS/okIwHRTm/Bqm+zqDOdtpww122aE
FwD++th298CwWuswCxzcwHk89wO6TL4pPDkSO5nxUWdf+9TebgrAfyzU77tnDuwp
/I+kpSyc12u1Km/9rEHvSIVpYQVphIdAbYVJ/mjgc0E6rbwo0kuknU9M1s9EJqZ5
PEU6BzwBbV6MyAHWbFWH9R3Z10ynALpyirlObXwrLrG+HabENRX1TNCFyk4KdRJp
HmtArCDA3fM9IdcvT53TDz3LCfqBvd8eBK6/cvtvXQj3jQEMm4uugdfT6vW7F7V5
NFJfnkYr52juUey4cigwY3YHCY6m/z+2mFhRUBKzoMr2pti7omp1Y5MP4t7pXvoU
G73ZAR3/1v6lwtpaFd5WKwXnzM/yuYgt5/o2g+F1LQ6spmzlXPNlowdXhskZo3vr
d13VB1ZnfyjNzf11LHmWoIGBlcRj5RKEhdWLqVdaw4VgqEgzSinc3n3qujduM8GY
QcheLC1RuNAMNZy1T1m1uGcv1q4l0I/z45AKDa7VNvlvCMC7tso3zkyBSDNwXybJ
9ScUSxV5+ROzaVo5rNHwQfQ9n1NDyDRe1BWORjdo+BVr93CxOruT90pMpFbnOV+R
Du2caxxn1yb/B+QTWQPlHNzucaIaQhoVbfJmGl+aqYKjfZLWL1HreFN4ZEQEJ4ht
vt/QPY/4Y6kF0yAotszyJtwCCnTrNvNip8inynJfvPFzRTBygTaG9KEH3ci75xKe
SBr22kFA4Z+Ih5fyvEkFgbvHkml84YjuRdRT4hvaBk5jSFH6Zn2NNeaQ6IRkbT/z
N7VE4csz+KkUiCU5OSjwhGNBfQ0Ti+SuYJgTydYp1hxQ3tJfDqmfBWY+lnHJhSzV
UdBPRwnlVfL5JOawb43G0NQnlmdmAgOHUlQagIHkPXaboidDffPkHvJBxRZYtqb+
YqJ+NuKmleSyOv4Fpf+u09ojewQzULMZxcoAKjfm/DCfBigb8hieg5WMiqJEIIXa
sd7qMXkTqIjfi0F/rmobJWEwysgWxZl/N01ameaOhuIBAKACUKT4EIfiIufkmxuP
Our94/pF0chgBED8HYvOEvXbFyyWYcDAoCTh3Az6kdWEdqYaX4Mw1QXKdharOzaq
arvEvQZbY9gYgiC5ZcJ9dgN/Jj+azac6MLFzxL/QRFIOsb1IjFxGdKBDy9wjtVrW
AVrCSJZ4kKXu8blvQWnogEQyEFiExnnOaQzjRnMgyzCZYnYI03kZMDfneDff6Qj1
oj4Orqp1aCthw0JE9YzwGk+IB+1FZ6g699cxOf/DlQNkJlvsZZh2PryGuEWfXDKv
R81pQWH9q2Diea3xxWZ1bMR92QN36+VCOMduOh80yYVUJZoUwAmtBTEsyHEFubNa
OeVR5RIT8Qq/tOacuJa212k7CyaNsFoDamp38N7wxPOkHqk2gtYUR/JVI2X6q0CA
RNZjX9YiIZj92EsnG345qqr4t9DTtwbrDw0/Vp8LfhQhiZkMLxt8Np2sQpd0Rw1D
KTAKo+6jlOEmZipWQCLpi9WwtbvlZPXEh3IPqbmvdYXaTwEO2NVQTqPMTFi09w9S
6kiBhxSsbpdnjvEByfkXNVCvb3cf58dW09b7hrbu0oTQNyTa+LCOtpuuSsnXEVQY
FyFprYcbPnEZhEdY0sEryk8a4yMpuJV6dXWcGvSCH7f4Pgk7ok2Av0u+Id35hD1v
7UMwcJFvYGQLKrhBVMDSeb7fEQw+wXAMghYDMKMT1hXDvAOuwfexsXxiFLvBO/4s
jD2G7k6Ohzjy1qWZbufoqUFSLA34zD9KEHx0/60BA6xhwqJx0BzaIDBNC8Uw0Wbn
xeQaCgg8RG0KeQ8AhEN/+VhrIiIszM8If5e8wrlujTcP7s8nGxVbklafzN4K6UZA
1gSSWo0q5vRZw05azjGwuZowlXExIw5IVsUNJkCuTXDYDH0ONcnRuJVyUT75l/5Y
ciV6MCJCHVqJVMe3OfARODUafeGsUSgBV0RHQdiv1qkBPzctVtTPUrQoT+S5QceB
Qfd59kQexQO/NVepOI3ru5Myh/HshwgRAyJze48hJyYJO1MtbK9p8f6C8DhKGG+p
GdBZXEqgfBZj7AyW2cnxWj/POKH9M1XbG9aa4LW6k0fHBWJQvTVt4oTS7Gywn5xr
BC/8b+MelevFjeVH/YyPqiRT4lILy5XbVUfVzSF+Gv1HvqT83CiF4NCFrnNbjmic
iIXb2wEAkWYFn3b0QlXbqngolGqiFqTNAz2jx19HMa1ql8KwWWhGrdcCApid+WKa
tRo5hpME6zs06BUGeGjG70RAPDGklHY8L3uU8CuEnN7MP5/ZBFOFUMBV1viK8tYZ
/c+677i6WAGnhymNRdZep2U3Np4o9SvmjCoVEYze776r+Lw1W15A4rB6vzdt630b
9adWqf6fIrce2bKZfGL/MOVC/rFRIWQPH0MnqZxEzkikoXeNIexLd0OkTQffdBnf
GcXEVtqz1o3oQP0HSnVUb5hmZwFVhQ9WxYYzGgNgKOrnJ8Ik1JlWMDIWVd3Rg4LB
QU1Ges5vEl4spm9RLV4eYtya4Tjrsg4DNgwlbKIoEaRbxdTo2pFjpclp8Z1tyytd
dr/+JX2vNC6O2hc8toHu5Hodg/sO4KmL85aS3nTGpxv8Tw5S96S53Kd7xmTDP6/e
ytL2NAZwB+YIu1gvKfMSFxZaP/YHc6ntkaMci6BrONA3xgVq+1Levu/kOoM8qqU1
nFSRTLObmhOaCF73vuWz3zBec868UtNqZG+lUFmqGF8fQ2Qr5e4fu3UvPjYAxzcg
yYZTqfv0kjEKGEuCxiawnGWGwTLou7pdgmpA6Tp4KWWplmJmtAqDKDUbF/bfuiPQ
Uy4UNO7QrT0Ar4Kevuqd8NSEuw3gIW+WoUwelaurWT8rjRDLJT5sU9oqBV6c/K36
/naxet5C44ZmVO3yFDgmRYGE7lA+1DCYywlJpsBPx8P9Pe+PXToZLkkH7eREbTQ3
9U7tRsPCGV4qSCFcN62XqWKpEzTP3Yh5Y2ldSYzPg38/1tb0Z19T6z16oEu+pW1/
8ymEQi572P/8VMtEmRqS1jtrVcf0mYPJJZ9W1SMQuZCcQsdcGWo+CS3L4GN9RGSI
K6I/QgUs0hpNioHXSkJo4X7+Am1FXDc2NDhhRp03CP0wScEFi2i5iyxxdmOg7J/u
VCCIInsfGa5bIjUb22cbbTGLlYEe8xliXaJg3fwjye6BpFBuqpD0iQDWw3eG9uMD
VMR1b8beG8PeVd9Qta/Z+h03ckfEpiwDNDhqR62I9e5eABqmqr3yrfJ8MYojio0f
uHS5Vpo0OW+K1NJkuvwoWspmGPNW7Hg5sv1u9H0ycw/WCP21S3iCFPZR3PA3CdYg
Y87gmw2fuJ9eepX+JXGOmeJMtzsv1X94r0BFcUhp6UkhRzJOyU73d2xJyV5T62Uk
+Qu7p78CiFBqJMFgRel56GciVYe+wdJCpe1CnQg+UP0aBy47vpNN8LX3aCG2c6gc
7wpCWlyUVQs8rMDSHkmczoVkApxIS5adZawr/7vEpFCzBR37wZ7YYVwn0HNmYZlR
2puJZBwT6cxGG6+KqvvJWM6pRpGnEu7XmQ4/bZPgKCDbvnf8eYOlqF20kQM6oX9j
IVuAWh15UMmqBbuj2YBcVJiMOr0Gq/KheG9OJEyyg6XkHenNf3yh5+H2A+L+tUN+
N+nGlmVzqwxHAryftrcQ4iyNxhIx3YKZRydoUac98vADNdDCKLvtn60pWf4lsl+O
q9O0j9eBCboRckoEipJU0UMJPwJuRXUHJC4/JEntPu4cU0vxC367lxvKkQ3VRnGj
e41H4MVVNMHvYSQk/1xx/36m+sqH9bM4ZZK/9wUvFumW9qJba6TyG0yc+B19Ni6N
Oxf8MUIWaOlwO/PTrC7kkGRgGr4Pm8MhGAFUvoIdnLMvp4Tk7o03q+EWdRQ+S+Qt
InDeoy28+gSArFAu/sC4d8czDAEaa7Fu3I3/Ay2WfjSO9iBEfuO3a5ty3ND0WuMl
WfDFphljM4A+Qv0dmGsV+Tzz+1XMX6NifSv1ii69zZ5IYCwfrs7Uyjeh2P6MZfNS
/mUvbC9z82qGRcdnF2Bmsgph07LACCJVyTwXWWu5PrhQFHviYrDhHGDMiNZnEvUv
ljw1rtKtawmMoqW0OiCi9MgLWIJEJrhgZtBzoz0gsHAbxMvqK2LYw2QFbNcrGs9l
NsEc0qcvrcsR6uLdOGODFO3bT4SxRwfWlIZvHr5ildHWF6a0Yk15oaJepxUIv6CV
nLNiYsDvv6aDia9HLqkDQGRmV5hbvQtHtvXokGW+WsQyLuQ9P8a9cYrynYu4mUMT
L60xWOyY52R6nPTVywzDHBZzBZ782bie79D46qq8EPSXEwwql45BP5BiGVDo2hZ3
Tlupqb48xKSXQR5/PrBfZD+02sUuaR0ETLME4wFp2QOgGZZ6+KW3GpUnh/hsvwUg
iUrmRTH4CW//ueR8n4qAmWKsvNZi9j0dbmUPk8oa4rqc2nQmSL8odpsDyoneb6w5
OahUS5pe28D0yMqf0QprjKRyreMfSIOVkltUx+f1kNB115ACH1dV5PJ2ZeLzh5yQ
8XHiZRSluqEeoldiM+wb4ecGRcwha8HLGbpaPm282wtCpKw9GW9fUEbJs+UsRRAg
ArUi78Y92MvdLAElXFNkPxGovtBnJcVDWDhRwSHN1BrcM3awQNrkdEJbIDOS19jk
s6nSQTnkIHJqHkrFOHId5aAb42tDCzom1YPApZMsehNTSFIAJ7yKqoUaWIrWymv0
EWJ0g4Riinkn06Fjweu+8mhKZZDD3P1iq2A0jtYqjIDRuf81pj+YoBrltr6H0Dvz
y1Pe+FcXWEpinXnUWNAtveOgAeQbrILf1uRbNM1qm5C9uIxNusyoQ8npQvyCazMv
TNvRgyKbdTlZkZA/wkXZoAdn2smoELyGyzWJhHftby/UuAyxMn7QoB7w7H+WC8Rk
rGyY2rKxyqR+YhiLIrLVTe4SlSgtlBY4d+4puGN1ALuXobQmHGAsp9ryb3vR+2M5
koxTFp7K7ccbyHcvRntEZm9PxdyzR+9XyepegmnngsPGACvcrCWz4IAB2J5CaPHJ
H86UVbAhbN7+/owb1fKiksR4iLbewdUVWjefmAlQ9+Ju8iO6w6s85e9I5HZQFDLB
bwVwv692kKf/vdPM5tK9vRicUewaq0vzO4bU3FGBmJyqAYPi5a60EqH1mn3Vderu
f8lufj2VVJ9nU4OYC8keFtTslQkoFQfJ67GC5znX3z1GQnImtdxHoUHnP384RnLX
0v5r0azBtBU3T7rZzmPRkzCoUpnnZoSYgUPUVST4GS8WfYZjdFtlaj3noFfx7tzE
DIFqd5MPx9EU8uRNxcdOghs/QJlEXmnCKlgF/6jdzNj5RgUxGx+mhuW0uhP4T+jC
KDVp5ndxY3dGGa3jKOyOdMVziS7BJgbQvIa+ccAG0DanpEiF0wW0gnZ02x/yYkkg
ZVxwm5CTi/ejPuzbRzg9UUTdZoEnv7/CzNuEpIwGyS/nhwkgKXyFQXUPyiKCJ4d/
C2vb+0T6PunrOraQs+N+2Jcge4vUZ7dMM1JTRkAvXpISvIgoxzkVGIraP6Cdkjyt
PwJaRvT39iHzRjId5f4VvNvJqcAW75fxNdG+wOfhyOPc4QG/gD0884Tdyu6QlT3E
y1XGQNpiTC9I6U8P17A/TXOPTgANY/WEGlvpECD2S8KstHZksZsehgsJZ+R6U+xQ
x51t8cPrhe8O2fWEgMVnkTuK/RaIuHhKQZoFyp3QekvD9Pilz9tqEPZccpbEi/b+
goQOZ+qI+mFnA6cIrkGHhC8OvJ36F+E1Htggb//m3uP1UXL4lRmCHrVWBlzUQCoW
fKcKJ7vJGB0P17IAvnjxXXbdwR+nl5Tzl3dDoAOCLY85ksn+RjO7zcg3LfFkJycm
bNZT/o6c78w1QevuRUt+NNlW+eFw2awz5CmIqe6512jF5F8vw5Wo//mltJLUXW6y
BcbABt8ObwFo+YdVhQMYALm6o8HZUV/Pk8jw7YyUqo2ZLEk89tKIV45NtVgm3JNU
6UTATeBtPkzyBW6CX5+2hZ/eMcAFo5qrLMiCJmmAYj4HWoTk6VZqta/YAH3rZr2r
U8KlpktF+rvNNKmv1YS2nFV5709vTwpbmfaIN6sqFYruoeRVFDopJifz/cKbHEqD
OWNPauVElKuGCUxQFJhxx3+6a9V0lShQ9PhthRe9BDDp1rdof40U+BdbXCZPx/yr
3N4IbyQRtonrBE6fEza355CiQGN7I13zAlunpF75BY8U7z8lTwuijzsy7EG/PMIy
sYPRRBfIae0Y3hTasMZWo00sm/fUNIKM8/3nq2Uxk1Dnt1w2UtPQ5Wi7fxVki58C
bOzBZlq9SPSI8m81dAA75DkO1U8BEEf87cP6QQ6JyOSrmM1VgDqccv37fNQi5KuH
zqF7KfeijY85Dnnlyy20GmL3rnRYWntPc+WYMEyBz1AKcELMqnMcoCtbbLyZnUWV
VT6dhWdOoPm0c98OCNLdxtzgOKrm2cU/vEX4OVLk2VdS+wgPxi08nqFL/h4CssB0
4yWtend4EpQ7dZHW/nVO1Pl8u6eKL3+0nwWJwt+mIPZykbVlUp+j6uM3wxHXh0Ww
NUWoiI+mFyDE6ot+KS2TlOfwug5qSrAHRKukgx2uw8Ys2C/2BTltlnMTLH7xRe7z
0yLVhQXldmbw+B9RRy+Z6Zyhdv4a7/VsQrv0OJFCk/6R+SA3cZeP41XFRYR27Hf1
qjOYdH0ruIZp1jvXXczZFizRRzs0adwiRGOZdprwx/yMBaMK7DvzrPCo9wo+XQBB
IbCYpeI8xg3mN2lCBw6FJrsDPaYepdfBA4j90s7LVMv8rPCirus81Nvsb5K4K39M
i+GV9Kyfium6oOAWv3V0FbtyntkCWORtJ6bGjfJBWFmYHJvf7+2RTAIPvnjUFoLJ
x+NAe5s/J7VB41rKLWra7KGm/0GvB0UGHkQ0GenvLv3DqN4ogVyyZOb5BHnQFAuJ
Qs3aUl/ZcBRv/Mm1GGiz0Dl/ULWB2krkx3tE8CGY0ZxX2lI2BT7GTl4uC6RUb8El
njNWYdN0J2O3SBtcLyTllxLDC+HAcbSoHwS2JyYu20sJNT6UDo4c0YKrKGyyImm8
yHB95kw27gNl7NMAQLdYp+vhX/hhB4PHmAkZV6CEwrIpykGggnlb8u3KNY7LKvpJ
N1ITTX88DCEaMOdQE0374zd6lKwB63VnsTDZjkrbHt6iB6vl0Tyz7CY3mD1DRoFh
FZSuXC7H9xoHcgyMzaVr/Y+oOB1Jyt7vVLtkksJ2BFtJSobC/7Ljy5I/kf3cDRVT
07TYVYl4yQQwDsO8tni5ms7hYw/mkV7LSWt6H3pvgFdMUIhKBJi6BPKOagLrTndI
hBIJXoTXntROl4Tbr4UTMETYSWpw8L9YUD7eyL6lohy5iivGi4Q/sucmU797CrAs
ThAwRbaPDsSUeTItID6vZMGHimDtxEdxRw7PsViA71q7cdKzcrJWqxWJHXCUxwgD
9JIAd7Axg9QPekK0saHvnBDqb6hSLSgNWbVXDAgt26DA6vpMSHqF0ZLGcAx87S1L
eE9TJ7Vm/P7b+mnjNJe4ezxWxUKeVindprqe6uAtgfzfg+kih0/PlG02dqxoMuMu
Nk5EHafSpS4Bgq/Ekmo308H5yc0InWB1XDDPGW8ctP1pecibaJi6bXR70+WN5Be9
h/9edM5scIxQakkGEGBCZjFmqr47xsg8YqxYYRD9mZ0bWmPq1LhBsethMcC9/Jch
PUWF+LSi8/vpPoOa9n7D5qMCtLXr6xQkHNxmJVsfjK7c3mvshod1m/wQyiHkfV0o
EPjup2nKBWzZ5n2fGJMkqMdvTfFs6O8RIkP5DuU/EW2+/44iLnAovtWvlNpik6Zt
NfxNGYP42zw+Yauc892qnZkvCGaQ7H35IBGzOED361a7haIpbm1TBj/sgedl1OtJ
M1Wu9eZB510QUyuEEe/zTrGqet7n3zrsAOtvQIKaw0CCkBnXuvSbkii08C4lYte6
6PetQa1puZ6NZjsYuABUpvPl2g0i+Zau5lpmQcX2tfCk2mDbxvjQ6RzeoeZ/iM/l
+7vCHFO6rRSA6auZUaEEEAzehmks5/YwqQc5PbDQ+ysUYbVnzg2JwRW3kWZF7PfG
Uh8rTVdqNyk/Ya/rv13ZJ7cQa8woN4PTVfUNsz2fxSMj3bWRT7UfvonAHGW46J7h
rXaKnOdWzPXaOiIFcrRySDVnfqpWQWIe9ZSe8MzwDCasEPW6nUpqQprXsO6vUqoI
gOg8OBm+HnXCegmCZveaPVU5XZNVjS0e34LHO2mq7pAZ9d06DHAQ+Wwp8JAVamGF
Zmg+xQG+n8NgaC6qoJUjaKmH4L6lc0dWA+i8kpFOasQNs+U621zP+bU3LBFC2Kkh
GdcoMm58jsIncd3wLAu4DgKHdMf5Aq9QJ71n4yXx2AWYhKhSs7K19D7f4xzLGYwu
DDU953WZUb4sNrmiSj10OLP+RhGLyOOvBuEplf4ho0hZZInieh0V7hKVOg8JOXW6
e9LD26X9RwURAHBtiClAtCVKyNjoLFYSElYzyvj/KTFreX9cqy/d1MTKfSlB15Jd
s8xIR0av0FEzgzo6fXFJCnNtKEoF+mt0noxtVFAJ84Fe+wH4qPRArV0k5dXxR6vr
cmMadbNtl25iVa2bUrdtbXrCLXxTlBOOtIpBjD0wGYiQFFAK+Nd9j53h8UeO0ZC0
NyNjGuJ0pSf1vnfMSLnQFdtSGk2/rpwdH2bNHfNL0MChWmXBRkd6227kbFT/xlL7
+6sH1alU2FEOAmt9HucRPTO3P1W4Jjsx7PgLwtwiFCszMXtGYrqoouiknHNi7poy
LTQSGD2zaT6XvsQNwb5O5BuO7zeJ9GGKS/L6n2ZyvF9J2Ua5COwXoZXXllVCOgK+
vCAYr+JkoReyjrGuqU2NVNn+DaL+LV/ntepJ6CdMCJhKKrpwlDWRUEon5ZyNogc0
Gxe+6O5PnL14/O5nD3SPjcblbDOB3BQEhX0d9ZHlS6cZinGY+kmK+GVaphUUTWYj
z+YY7xHe7KpiRGGlFEVg9tTllX8tvwWqwECZQ/1SUNMJkIHU7uF3jKEE3SmOFHf2
6YTscqE1a3oXURIrEJlNfhlJAkWXEH4/dUYU4X6WhoQreWh/zZ784NP+VONS0htM
Jz5+hNVPAVGkWmVonnPYiYWSmn6zd20l5TVnC05UtEhOa5ZXQisfRjzp6TvwltNw
uv2TFYgfKRURwUGOF3PW9EBHv/GbKn5S4TuAc079XXSWHyOIy5ywi5gSmw/XkJhU
9VDujVxc5yqRonef5f8KyFYKjB9vYediCNAAbIoV5XzrLwxLzLGKuw89e3QGIL6Y
HpVg3kzkdUN+b5LgpLJ0Yw7xOBZtA7eWMytYMSX7jaXWP4A+9Qp8hHaisHHMNYQG
2w8qQxzrSwR2v4oC7/gAZuxi+ebyAbdl9XFX49zti4kTLkBJdzfy+rjg41cEApb2
uOYB3ousoyJy83dRBjGnqybVcAbo+0YDTJMv0hT+LrfXmIMMJChDzDJ69Thf7krz
IiQktqOfnZQ5boqFj+xMUHMiYvKJp4FWmIQjvIwfLvD+qcftrGiNl/17ZYrDaWUC
i+pl/XnJfh20Vb7Qn6bFRoChvar0JDYlN32PkLN6gjme1cajIOFG+MQrKfw/+3Wy
VY/JC/BsVFUOO4ouOyEjpC/rk7jAxPQrY4f8582SU1mp5Ivkf1ywD1lAVq/+lRdC
RbIupvHPOSNi30n02FlyO8GTiU7sWgQxot4gOpEHNZYI5dKROeUVYbfUUjai0QSI
k/TfteD/NPL0QjXA9fbNZunLKyRiodigfZCYSR1nFJmUwMYwG6km5wAxxH8HWsp2
hDn/Mz40rWpEDfkVGNtbxzV049fvG9unRaydSXXn1Ac4O9TbJlVBA/FaHIZxD8u+
cy+RPLJKs5KCG7pTQsvOzvPBvYx5gdRkGD7KlU6HzX3J4OSwhxoMPPvCKGwEihFY
RNQUCejPmdmuz2S8Ev7Co1Cry6ID6NQHNH4pn+Vu1YJF6ktoxAeEJ36fUa3R+bkg
nfuIGE5PekTzXMuKbWxb5Ek7RlMcIIRzyvuvTPI0ArCOalc25fTMs9ebsC3mrakA
pQU2poH8y7EHxMsIk15w/vAvxpAzmBi0vmW3kpTFdzZnLldo2e+C5UqOY7vkOeGa
6pzeQpAWPabjeJTmDAS6gRUDiNYnH4vrm0e3Tz/PcRqVtZ8dpEqOJo1jMTl+KJF5
DwrhA65PzFqg9uusmLrx+rCNtSy6Hk8wmDO1njFpUQbaJSUzrZsvCH7vDNMJJ+jY
Bli51f/nZDboeco8rjtlL+RV3pnl7sKhNR85KpKuNkudf4/Mt8MpIAv38iB/4nlc
chcbVxKRjopgMLPY37wfPYAmxy2HDwoVeQ+tMyUxvFPo8N7UiJXxUQiEE9QkB9mB
CmNrheo9lJpxBpNK1b6I/9Rdzk4bgtmxWjNR8NWtEM0R6XkSJu8EDJJUIgo9q88N
DN7ONjNFcQnGpqTBz1svpBx0kdh8vzBoHrcmwC4KUO42m3GX69xABgesP4+L/boT
bnLv/OMxJIp19qteh4DGbGpEI01nf0hNew/yTvUuToCEv0bSf7bW6Zo4MAGeh0us
qyTI98v4BlLW+qKAve933bDPfp3UIvyiKxwDHe8PvgHf6MbC9rCvWHzZUpGSpawV
x8tWdbtV8dfXMJY0XOg2vRYSInl2lwsvmSWKAgLN2rHN/25mQfDFBKq1QEYL6e1h
0K87gC0jkWF5xCsQKQEOqGcaAi0q2o3+ahiuA27QBsE2zxFf9O+3Q2XqcmNaNyun
iIL/003qp9IycNV4rcxh6EYDT4ZjfpuvrM5zJ+GvNp3dDIkAEYo22D4IfBZDcdUM
WOyN9wsKUNaWksD2P/M+MwMj9zQOP82aGiS4Q6b/PZTE9u4pDzCUtILWBzdcaPpk
vZgvxDJzhKwSl/bSzpMpV7droXMXYE2bVRSKt3RHPJGgbTAz+xxkF7/ELzbB9FWd
UXGNHAl9Uaa5/jMv++W43s8DPktPK9UBDr1ntfwm1TrHTFiNTv6sNwm8v8hiAZuj
so2KbodLmOABcYxkxTVCwIxZh0mqWs1+4rT05scxgairoeZcpmVOrJODneATfPbs
VPgUXjctG7Nz+xZuywAyPmkFrwVCXRwPZakgGuMuzYIbuURdMHtdLrLttwlEHU81
gjp5MoD6VIY7oJHCBlt/OEuqiG7PiZMyLwE2DSUkRW0y4Rpx67QIWyBYUhNNRfGJ
/qj8nN0dadgQZZ1u37W1pV9SKxgH5zdIpw7OCatReG0F3fSPTAQUqvX7Yn+kvobw
6up4MmQXhW3SnkoZ837aZm2i26MgTyREBC5hEe8y7LI9kQQiGlhAgrtRtesUmVTQ
B43IdeAliJSrgaSsKXmHXz0r709jj+FjdzRJ9NKZFQ7AKY20Sd2J7TEVE/3kVK8p
kRvs8+LYb81kBmAmPFc+sB4urlJWRsc+zw3VugU1MEPWRMEVsgON6VgmwbPLFPnf
qRBSlRQ9B5HOJzxxLad214Vlzq5yZF2ExfVQmTAnYdxRmHBUSv8NylSyGZ0smSav
5oc55VfT34LvdbqXp+Xl+swCEpRSBpos9sb7E6675TE6hnujRazlHaPj0bOiTomL
ubEGmlo2ZNR0EopKk0bvos8mQi8q1LsMe6kdN0ouZmiIBF0lm6vLmk5giGVuXCzW
p/6RGteEVE+isb6FTm0hAVPW2EpzBvot/LNISHoRptY9cD6J28XRbKeOoVNBAWR/
8JaIBQX/EbsMP+AP9c1aUFmDKYKpWB93deGm/AGK5BEoWUy77tvjKQbEdIjtnKSM
ccPAaY4sn4nhMJq7P40lcJx3cDRcEtdz96LppmUKFJfqrnU8DMsnpyNAwz4cAJai
jT/WvguqeeLdff/rYjl9RO0Zn2sp70m0pfZneYt/ftqlLjJ/lfpruebVQiev9kFZ
v57cbmJUBuO4diJr2VbxZxxkzu4cw9IBenaiPpoDnppkAS7mv65127k8CH51kSa1
SwA3uNwZuFXZjL4oafFpIt2hVUs4A9G4omMS6nnkrQvelkgwFYslqb9Wz+I0ZvfH
1Fd5Iy4BgYXpH8GrVTtrYJIZs/e3GQQM2FJlP5W+WC3JQQ8Sl9O0trJXMfekf2kI
8diChq6layLWVcFivAxxHKTpWEB4wePHDaQljovU7dPz5rR9XeCqL5ZRVAIYjwMp
D3GkebB+LaGNJBXTI6W8Q43Jeoc4kondPEtvFAW0PSoc9Rs3uoOzKRPepVrY6tYM
OI1J0DVLsrPKVQLgGySqKNrZW1ek8wHw3Ief+N7pYc1p0upCfazWkzZfKCmkKQgZ
YiZWusnhikaywNiCaVc2R5C7svecAy5VBHXzNWyPnt5W4Cq8dyWx1C31EqpQMLxj
1WuG1Rqs/RUSi9rVIhEnvQqxV45P+1f5vVTciVqVRzlxKuxyhMixS9SUZseMlf60
LJEQ0HGqTHZ74SU6tPHtiIt4kamSIrK8WgPdkZX5TxJYDfHKANXWAwawZ3FQpAp1
lCgDye0va3I6f5oMB1B/yMgmcsY5kdzfvA6h96ECC/BswgUQyDtddY0bhHecf97U
KrXVNTzxOrd2bImqkbKDJnSRdBmKTQLkY/P8F8fUoiZZEjTjHES2f8k2JJifOKYp
R9scdjgc/evrOOHC0RXomiVXEbiSLCDFtjn3Vvu5nVArILz5jBG0ThHaVuyU0Qwl
43SLmAfb55rEPL+swhQsOK96uMr3CvN2oEjQRd8yEdeu30uQXxwEh4gH29gij1vT
xPnrUt65Qz66qIZTYwQ0Ya/h1fTmw5oWnLuBBWhovepwjF8bIdSso5riCmw7Rkv1
DApwdJ518nlXlyApCejZK7iASqaT32+BHW+H3Ccvbt3I6evVHuo3fAU17v0KRBSc
oOrTaUa8ysnU89PRJJGdQoHmUyadqEqh6nj58QjQ8GQhVYSpyuAoT4qBbffdwFOV
ts5WBoXVRZc3OodyEhiCtC8MahtO/3deWULHG9Uak0OWhDXII8Ou9pvuC/gWE/bH
wHE3KgMI8uqYeiBWBrZ+fuBpeh/BYdwItumJ7Kgwkq1ri8xbhMcl3y2XxtNAuIGk
n+UD/7qWmv1w3IMULik+wYytu1i1+tptkbX2Ta4BR5v0cm2h5hYWGQ6DMj3uD3ck
1D44dm6o3F17siPY5ExPthWjfBw4BA5GXmcpycveeTLQ314YTvy3Pl7Aq1i8ZuTG
35EEcmxC2xQGYzBc52sMRNKTDT5Xj/dVeFxyHSq1vJ6AKe+oYYfv8e6vRT/+CGrH
McXizOPdzuVYPbkPSIyF7RKY7L+iihDnZu6StmGHSqAl7Cpl4GVijQ+933XN4o5p
55y2KBGLb9SrjtQ7XKCsnbNuFPqCNOs5sE2XPTgroKWnPafwirZMhiC4HHQtxpuy
i7IL3fTWjVepAbwLdaKN1sJLeYJgIWZR5FWHQvqzJwhpSaAzwJhXOCoiYoa9R0AG
vmriBbP86VcP2Wd66bfRfoeQoUzYMEKq9Z4y9kVodK8gMlgG9ZyHsWcAS8yc/grh
PnXo1at6/VzfKqlG8g0sAqe1gLVMgeW++IDZ877ZlV5ee7W8yUw2HtTkZXROJx0v
SONXlC8DWx/rEiXkEkPOimjTBoBRuy+qXPk2iIthop2Zaeuy1daibmNifrvR45Cp
/ueU3eoppwkZrS7cffgxgyfbp21ivXoEdoq5ZAwzbmSA/WLQ+B51OM5AY2RBN1vK
5fmn/Zma3hGPpsi/rx5CbbAu+IPABnIe4nOOCkTG+mN9CQ5W209E2NB0wzxj6r4y
yFZeEc9uCEBQ6Fk/ZpPOZKKZ6Cz86/QjMRHV/X+6PaBlFkLjjnQ0tQC/YcSDZeSf
ZCf7D53EgOGvEuXcnB4c5I8koFc8ru8IAOLksvHrF1HBA9hINDEO2XsZqLjBl7nB
KSSG3PqgwatbMBW7/VXnGcMkxOVShhbJN7WrGAH/qggupuD0hwJq5qW02Q8rMR+6
n4xfTN3iAJd+7G7Taw9m4a33e6SCRa+Ob5CFXRzr3X6rCjB+wg0xui3HTQSReRuM
V14T1HAvA6F22etpGzyf6d1Mwu4CYDrDrntsP6HDe9K9JPD14ZUP5X1Ba1M4qbCh
sUrt3Z8T6/KxsX8q921Sq4r7z3/AMgssoFh5BSX/m5STzjox1xs8K6D45EBbSAqe
HLJlawa87Mbg27aBw/vnx6kf0jzp30nHjSrHng0WcbEerz4CidbfJdnvfrimJOq2
1dEhOzCOlH/g6ccFZBKUIql/01IfolRpy3yOYx+TzQBgzTZo0USAo1imcPLlEH5z
mur66PD00paLAcDe2KJOowUV76zjCOzTIJALmX/9iodyMa0AIoX7GrSNmFQoSz1P
VcClyTpSMOhBf1EyZr8KXxohn9G44/D7b2zWQ4XFzrDrjL7Kv8RgwzeYwe1kBKbz
WyOjipLgcwkqPQdeulZ49coChY/3AegWdNUn/m04SuyvIz3UhJAEYPun1hILle/b
NEh2oq9ubxwM/Z8lENZR+/aFMG8nxLiAp0qFUQ9Xj76VN6qsSTUkk6ePg7TzKEwt
652CV/Dp4RxO1d04ZkwEaB/BdmWEgrR/6YSZ27YITVzA7G7gmHzWczLWBjNR28qB
XpfirkGirdlhq14JLxEOuTd1vBEWUlXvynV2rjjTunGybO58kfvEl0cXXnj/xnjp
mOYpd3NEEz+O9W3oahY0aupsYm2YMhxmN1NTMguwtcwgCPFLiJ0RjWOP26RRgOys
6aQcVgpFSqocsEAIu2oYkobnHUd/7FKip7tSpr0m24xbxMekJAPGyWTUQJJGb+YI
nOjCGLLoyqMNH8RZGWZZnxsN+tppNYzwADNYUxwsUAcQLv1GBIYr/ztNfZXjSe53
eH9lfuxzWpKkmAlNsI2REv2jqEOTVYAxZuow7pDjfbI0Y15sYWwZCbV1ld9JFHxK
2tpvu91ZNpedaHwdoaUZ55Yd4iUiVriKfvOYv/fR3pMSnbtSO3zwYaD0+KP4Ikfm
gxooOWJLaFXaudFr+yS3picnxz4MqLtuJlAUPRhZyskN1jXZfKVRR6ZNECE8U5nh
KmgY32DrBe3Ftf2tD3XLz6Pog7k1jntz6etfIbDM5xQ2RwTxQ56Oq+YT3FO69Waf
lISmZYLhJP6kFd1fvDDbRwV6Y2CR5SgQR53aQxah3Kd/i1HTgcX1CrL0ljWo4+Id
bgGC3Jg32bJDLAB4mbbr4AmqXIQcl62tjGYHU9p6ubltkXwlPHP3AbwCn3lJHCM5
t4juuMaLFxXQRdnXifoELh8u3dHYCxgFGk/oSkqgipziww6+CLlgf1/2g6DOjTKH
O962U3Yfk3AtJZzG5+3qQuDfTaswJqXu1BaJtPUu1Ya+LwVRRp/CNg84/87UmVdG
pbJXCs/hRxD52vzMo0SfDWTdb7Uk9w4jmHSGSrtRyGPMiulQmHGC15K3mx3PvePt
w9CuHc78029CEKaib0PeQLMOYd84vRHO7s4qNA2CRMFmMUgpVGG3UFmroXUxpKnu
5Ikhx+hb8yr6OH7bZ+ZzshUctOU598n+F2settmRfLOBXogSFpPCzrpMw7AdYWUI
SEEJX84+XJN0ZvXMCRGxeu2cm1iCShflvZmBAvAEUig1/38cRRPlFiLI2+ayxxZI
FNgK0ic8eL/giJSCkhv7LtfXTSe60vo77fGRb7Br5BxC0X+CHxc6mzQGp+iaoCsK
miYFVG6xkJXPBP8fOtIMh+x6Zp7ko14zwIHX0pi6ZYLUSwrafkcUkHTw5SySBQ62
focDI+rQgXTHYn44DcMw/zp34tYw7NzVZHTWBevBE0FL9HLu1WLD1rUwPgVqVKPw
j04j9i3jbxGYASrLAFhiluUcjvucOtsMWi7S5C7G7A97qAjfZ4eN8eVW5cgV6058
mpGgMUbVo+uT4gevDMYPYrbeJk9PCy/NDO3mo6/LGfvFeFSWUMlmZQQhoy6Psdx9
CRVAfjbaZwKeUH69BLxRhe9zQBmEvJsdzbF6Tsgx25Eg+tI77v3FdhyaIn5CXLYb
SGr41qFTkFLpS6Zk51zUBywRjZ780m6ARsxKs76UMNlow6mEj0x0d0WYHWTGgKbr
7X+kIseisl5N8bV4NcdUpPkY2hFPkV9QLXFWpN7a2T4ViMqC3PfgbQW3ai3aWh/7
xudXf/5W64hhgAfDEqa4Xm/+H7KntKo36TxG1ZX5W0Bi0ypDhkmmGO/AvKZZfMrS
eHxdKJ98UMSj72VMoed+yFGDdhuox8qGonwgintw2hokq7KSLZHXhWxhLjJUhB6h
WajBxkMknsYrrmwQLB9Pk60m/MmLMsyLYPfVY2JX83y8ELiWwb/sQg6oKaG+FZzJ
3o41zLox1thT4/3XsGSYiYQaeJeJTP87Dvx78Z9wmkvoup/3OZiD0YUoC2XHhS8s
PBcjcat5/s5BbXgbYAT/pHVEk9Ju3j69ZiYcmVGUoj25HzCgQ+BDIeh4QMFUX1Jt
fAT+9dp/twUqlmDe2DFH3uu6pdbUnCwQA6lLDjhbdDlmQlJUKYkwufcPTFZ1cRcg
Fgtym4EyN9ZWZDyiDjFcBmiYcNR/Bdm8ZSm/DQPoHBRwkRjvb7bBhEcHYnh02b5J
5LbKWogSLOQpg2dFgVeQDjl/1AAFnHwviSzSYbTCrUwh4t/I1BaQ9HQK2kKHQsqo
YAdguXQrKaXWv7uxq473e9j3EwPuRO8YfHAqbxSPJNMOduauy7137LIujrAJA33q
VQ2gx3nzkOGd7h6Cz+3XGDG+nWbdmPe3LmcgLiNwdzcMYfjfeGnGvw+778zwTTqg
7x92GNCPvqXUf8MxruD5jSmdRlcd08NGUCMGUdf2PN/jCZrvadOoMGVRdOlMRjoP
FUWdc5y4JJ1yIFeH59ADNPacJNSFncYTbUJPpDvKIb/SkwgOUxfQD1SwUI7dqW0w
7U/GzwrcuL4+iBduxqWqv7PFpRyVsOfoCUzU6sxPbEh5J5v1bMTI/eC1LC8iKv4Y
GXzG1nbdnyv8ZJOAlSNzFcbf+WENoaSgECX1iIeeuD/UKRA0B/CKfrbHMrY0owGw
/9hcNMGzvfsEO/WdQh9rQeRoevojHxXCYiCAOiDy7NDNKL0MzVCECHyIa+VCIFDP
tX+MZC4GOtDmbg3ObkliJapDUi/Wvhc2qDw/Fx+11uT6ux5NyhGEiuUUilOP71mp
EaohmqG3j2ynS8X8FJlGd4WmtpXFDaytnapJH3fmmiU2eqC3t6qGXrOMCDiAmQFU
TsTxPRl84634Wx1NKcyTQjjR0RbZUFDQHfOXhC130Abd5DZBy5z1qq52CnUGIHkS
VAhrXrPF+LnLYf1VDf8MWGAeu8tL/V77qmH+arRfOtOdlwZoKEfscLxYHLldyfpH
0tZnOstYU9rsANOEDs4NXFNJI4ut7WkGuwWYOqBTGBAX0ZpK21J081VHGZKTQJXR
7g95mK38aGm9KWKQcIL5FIzWmR+z0p1HLodMa6c0JYgpezeEv6YOdmVgRyUIuvmx
AXlYVuCtDv+pW/tylMDvUXxMSDCiNusxLNl5iN6E2PXnhemE+LbwzsFxlYmjnKJ0
E1dQk1K/xBZ9POgyQjitJ9oxplyxXQoVkD7kLP9mtN2f/9Ak108l66+aGkKR5jjO
GO5BxjUDg8GAR6KqxunFW2uygpBumhDgf7kdf9Nk8nGNslXSu/SkY7WNEFdDjGjH
QodLdGGC/HQTVz7yBpvz5hC+E3f3i8lDOrk3TIPxADebIZNisUoYmFMU8QiHEoMj
g/T5S8y+lYHsxojgQoQzF5/gKhF80kUcDglRRWXE95oVSAuvQeoc+axH0y563L1F
GxKynmr6ZRNl92Xvw7B/NRDPMlg+8sUr7+7cKgYKd0nbjoKaK5sqjiwN57Srr9/Z
pvPuu0koTxh/pnNq4+vkWT8tSKH/IChTFkuIOC2fZbqF3FLOi9neHcVKsSAFP6TI
0OkaeZzFiXmzfL2YXk+IOCfnlmRXVXBGpbTA1DCS29ZcDjyqyii+85mlFm8B4BPw
1kJbTM63hyExbAJZ/Xv/OTXC6wV0HtTpWyRs9bzBpUpmxCmSSALS1Uafc1h2CM3K
p+I/MACFiia4jfNkoJbkncRbV/BHn84yO9K2PSeTCExWaoSTmPea2U8RGCTudS/O
EsctwDgaeUgipJPGonPWwXAU3ttZq0NBAeYfE/L5fVcRy8eTbz4sW+xxcuADiLtO
pFqUWSbajPj1oQ7jfU3E1LkXef3V0krtC35GO3UyfdJ1KE7qeP0mesKeNEQj1O2j
2/cBYSJDoWNZftCC1DAGuTqAEeCuz0ri4awzrK2TiCB1G1SwpQ2iNFftXMGZA3AB
mXX3F/aJaGZiZeKRM6u3jQ3iI1r3oaCQPDkWkwbB5x74H98TgAht/XVk1qVBbH57
k+RczCRBVg7gmPeEak/W4nmwqbUhxM9ypIsk0DExw3s3gYlcLgy7+64dnlE6OeOb
tbSM3MI5uyxXGTnwJ9jhtOHbEU3ApaNJLHvMDevnSxtXo8SQvgbcbb/9quRcTSKE
wKr4o/sa/AAe4U8K6QS0Xh0NPJhjzwY2mAjkMGrWFZrFbR+4BIqG1h3dHqaftNjL
hkOfo28FQ3HbG+YYgL7N8ZLVUNgufdyDWiJdmLYAbDEmk5aoDDbVJqbTIEoFCWtI
piSV6ubS6d4XdNiAlb+olApoSNhzmXzm+CRtLIM2Vi9/r0CWf+hoIysKdXRyhF0t
QdcMdVvApkOaBS30cGEN35ZawZkG6hCUhAQFANSkqmQ2HCJPYxlp+DwxHODsd21/
UrNn6YZX4yBjUpj1g8oJyVJLiLdt15qcjnaZK1YeyeU3IKaKxz5LYSS0E1IfUELh
DMMmZ5vBx11nuYnKQT/ZLuHA1W5/iOqAHhor1mmJZN9tx+Dd5GU8yNTUrAwlEu8U
diAU+P5nUojuVhxjpjV2zuhIDnbDXqi4BjiqJqTVxaCn8YwVwOQWuD0beym7xtbd
Jcbm3clyRl24oYOXWpAza3oGeS96ZqnpaWOJXjDfze4DGuuLV4jsj2pKma9e/jax
gpaiyn44OYH9rYBFkx1YOiS0oPH5vggj3koz8/tbASKMlO2I4eSxOmLC8KYQqI5g
1h3GQYbwlz3aXWWWwsDIpEfTs6kwsOEkV0oD3YrcNrZSgbolKaqDD+oF2ZMUebnS
/1XXuiOyFWUjNyrrz/t9QUT8F41XjYVwAhY+LwS41zXaITs6kPQnzYAS0ma4k0vN
4XV0nhYuehdgCS4FNFu3t1X73SHs0LsJaEkUDSbxbzpAuyT8TsfHEuwMW3kFbTjr
B0e8dUGlM4PwLQv9W2y7QDcRxzM5c0avjlrYEibN3N0j+dmbKW3DWfuwlpwB5Jd0
nSg50ynfHAdIaO0WJubqPIpWREddz69p2Jt5bO46Lv4Z3Qo1AxOobU7ftRZQIyl/
wXuqWFV5djKRLUupoK/5jUx5fPIti7wHvViVX43ach0lVMd3FI0oTgKM0D2T81Ff
0WWS6WasS9pl+cVaxR7lu2n5Sp4+IaLOeotGjxh7qZ2AIegHdM/SUU8hM9OEZh/t
KgQunrExjAhIYSHhyMoQkwmdxk9MBjZXyUQAsy1H3ShVYyqqbEKphwQ65ratIahz
nQzV8uvh/5orgOcIYDJIlvzXHA2HokJaYJO+bz40Jk1kmVJOoYzSVAeu1CBhpEeK
hhqF9IPGFqp8cwg/AD1zEm12YIJ8PP5eS7xqYzaj/JfQva+A1y+6afOFWHAPSRvH
hiUdFIPI2CBXyEPNsGqOUbD+MZN8OWmmrRwqeQkMdC6N+oHnaHIbttDQwtokEeai
shWCBzLQLUfgnYHwKOSSELLqVOVkMlwfP7SDr2HT83BRgNeBxxwFMc6o3aNQ77Rb
/bxUFrduSJJjzF+bua63pjIOVbGZwcwcfW4aZFmpFG/tPmu3nu3KjAteSlM47iEB
6V9pH9b6UZGUv32DR7THKpJmImABdx2FsjWtFGpImcisobWFFp/r//QNDcO5FIvK
hVFcHQz8jlNgda/Je3DQLt23w3coWN9d9dvCugnTbPXvc6WyHYlRmOq2VzqjUD4e
Og0KOK2d7lX8OADVuT8CcFhC4v6xdGbQ+T4pTe5K09PMQCiBqJ2YQ2Cesdc+JImU
1BnUR/FpUKa8wUmFh22DhFXPMlDBkwUf15QpB7zho7LzKE0XKB77NZdA71Zj/cBg
MwG6EwTIfGDGfercYtCoQOvhOvydYkOucguoBDKVGA26qnk0/0TwYJExW5lpOtyM
M6I0IEv5PhR6gChpekfY8pc/ViDiOeM+xSNvFvebVZO62Mv5LWJ27+gNExr5GWg+
xwvYdGP8zH9BJmilnxOL6h4/Z/y28pdrdrMXB6azDCmaKw01IqhbKXrjPA1jHu7G
Lr1Fl/aW1pb5nFEtNIwuKA1JhB4yBC4lqRcMor2fO66PrC8nM7fuxNB69cbrAGrr
Db/3yCc3aUvUC1zruTUCOm41hJBOC+ZJvFzvf4CT5ov/Y8DXNvuZ51TNWWeLdVpC
TnIfNQCz7kjLvc9riFVZ5mC6IMGqQR5Vyso+XnxRw4UrjmTdJx6gNo67S0NBJvN/
TzC6Uzo76jlDywraGC0ykuTh6dbDKZNDe+v12lzVqVAEqm98Mlus/kkRAirNQjyG
Zwmkv+E7zIxo27AESZC/B5fGRXE92IJ0gQx/iogDuciojPUb7g1dvM3Ul0TTsF+P
coYXIBy1St0bGV+7RBJ3xQqq4ytyFkHTZkFsvaU3CLYUajIu0G2Wt27c1Ebqm2c8
i7GYoJysUOGU3WD6aVusrnC8OQEprLc0ObJIMRS9wQs+sQLaNtnvcsDOxeTWeF4x
zSpCoMVWdjjGIcB078dxksRnEVsZrsBmDzVedzX1be65+JgAQ9crymbH+isvWBS+
++IbexcfVMn8PISUTneId7XCA7GvdRicCc1OphPQtlUYQ29REcSrSVtCTjFhYEpS
N4CjsWjU0dcex2mzB1X+RxzqrrbNcB/mMPjA5ODzif/5d953wu6YGJfOqZGmtEWI
KmBcB8jtfcEeDH0HlersoYhMH1sPKpIosD78eV0BvoER7AGa7RURPSMXEx4htOI1
7C/Pwh47cQfdFvL/5kkadoKT53bl1v1pectNa4IGBgwd2FX5ADSy9IKu6sPlS/hc
cDxTBpnjkFzxwFxfGqIS9i0MJFjwQHLADxZM3nVsxNqjQyN8qCpPhlVLne/aYY2Z
QAIKCdAqlFkjIQkIRxn6HIdDy+/tj/nb1yKXXWi+msonU4Se5kOPaRpVolMSm3VA
6rQnvdAOhQVSYlT/vokrCP5f71mIGayXyGayG/kzsfe5t8HdFmIm5p5VEKIRrbro
AFUtNK+7E/uBMAWmsj5PwoByllbz707eAYd0pTV7Ah25amkwdMUqel62f+BKH6SE
InWw4rDxnbq7ES16Usgv9W4r5qFJ0MserhwrLmdNSspTFajavC7kby8JTr95tp/p
wh8t26ZD6vsOk/dIDwtT7t8P+SWepFUaB5B+3GUCxgiaIlxVT/PbvjDmAVtuxjCc
J+ZRa/u8hjDx5qcs3ZVPbhxY95ERNJtyQp3lmsX59T7ONA+8IaKOst2fl+MK7S6f
Cx/4uITSMw9Ung7cpM4q3gKwDCwpJidfEtugK7e3DTVkZjI9Lj+Fv7ae2q97mjm/
WOq30VKTrikeuxYaCaLnK0jz1k/8VxHAfPLMp18+C3LDmxbvmzOoHbxOKBrBFjz/
Xcik1+aAr4trKGe0IpUAuO7qJiNVo6mi18doPAf+srrRBuJaa74eg5iITiXpPXZn
jPeoP9P9fRdA7EGhZX/48Kjzo5U8wzm2BbozmbiguEi3OCnEUjCoNbSEQy/mGzgF
Ql+h86GAkj5mOkFl0yFKOe2kg6QGu7+xWcu996sIsao9iqRsCZ82umJho4278suG
fNJ/Ao5DhV93kC7N0LuyuBMBqkzM6D09ajpi2s8IC3JhL+TpunxADn+gzsGpskuf
hYOgkgqDl8MFmUmUphdQFNe9sLR/jg679B3UxsKRfCLzisZh7m2Y4rsZy9GLhMro
wMJbpFvRM8AFRkcLoJYvKD0E+M/ukTwe5I3yT0f0YpChGnvDTtWL6hCI48Pb6/c+
Mqu8Gjq5Q3XFZlr7wj6D7ngroYLQ+AOIzDDf8xyGLac8SDlBUm5mUGX4nAAHS1UT
Njzz2ucsV9QP5HVA29EHx7iY8uXpjJ0lUbhJEnj4W4xSOEin+vIgkEzyrek2afkd
LRopYkK5cKr9RYxTq9SIA4xcz2fFIlDsSyP0la9f2NjHPXMEdeQWp4mDWOjUqw34
3L0Up9wiTGh83woZPdG1IO9kRWFKgrf26zyGG0/NwMqEgNSUqfJsdoUn7ODSfvsb
lG3Jw89L5qBa6pCWpOzQNq1T3x2JdcbobiwtYTly+vT9wEw0tBpkDo0lFDUeF6G7
0LJivXrfh0P6b2PaeiXsuF9m1ilDgBsahsmoglgJTCnUDCBHxyQIjhoFc8ZDXSQG
/w2DLuLH6UcQKPRHu1AuXnNr6NsGg9IB1lZfCokhXVIZtYqJxrlgxckjMqh3ForN
9GFyQEj5nqGtkVToE4LpVRQInslriR6ADTiKu2mbpT8le3hI70jyvU8ivdpQUp3b
WxP25wtCmDrLhgGaeNcoggoUzg2ZeBvEksVdTCxD00QdTQLSlqBqm+owcGn+PYxx
X+0Hvq09Zs6Y96F+dtplTGtUXeRLdh47VJiLa3RiM0hAZDFi2tJsdTKx89W2o3nW
dqQRGhiDhtNZhZO1Z4L2+wQ292o5C1MItrHuCHJ8M4P0dvE3YDjJv0yn+xFd3GQP
a6Kp4TOGYUwLp2rIx/wZj9mJ2koAgxFZudzii8np0spaUtou5i6Cmpmr6j3HpBC0
65bLE9e5FOjZEoJsa/6s+AGAXsAX7QfrO4TD/dCOyrit74EZUPUWLu9Asi3lv/4r
J/bxUG8R92ch3mdAohVI4UqqjXjG0RA9t5xbMdCzQGdjvlYj4k2+db79tSCr06Fk
XMUt2PF1iFrcWAm4UOq61oyYJ2bHL77X/qfsguqpsUvwf9klQgkjDwfGpE4S9YOw
ibIWsTjuInNev5BqGEsOmiYIMs7fum4hSLFmhny9ZDrcSS5k1nh944dLWjRqZRs9
yxqN/m/QdcCMtbcnkod/g+yblGS//FUOZV/3BQcXlPMdXEDnw76O27qvOn39NtAG
rC9DKgHYpoQghKZY+mekpOzIqnTF4+a1yLtBVjnmXtq+9kYpyMw0ht4F4fUmm9mC
fVRFr0HBQqdCgsN4XEGAWeLDQOBOon5u9XG1hkXP2ivfDRA7W8e9rIImdy7wI0Kw
AxFbin0pmjOYJOQEtPGJgL1a9UfPTkf+vnP680/e0DOMFhGHS9y9QfaErAb2x0ul
CJTFPVOXgm1ueGUSds7ZK8SLi0ay0pHX7mzu/PZ9Dboasdgk+FR+K9pXF14gVazv
zqUs76ieo0I1aiprlA+9J6ozeFOj8sTNwny+PKzKOwtCiEcoiQtQKTDPnlXg0h/V
Dn69hsUrux7MK1urA7Tr/d1cldHkj2grrcUm1AzVxEKR8US15Wt6c/QIUkACsJUL
Bsp7BkODdbNA9c6ezmBMlqEFD4NUwg+V9ReNhggmPYROKfKRQn4T7OYL+nrXJqFe
beYPscSDszbsFGRjUHqNtWEMH7cm3FZZk4bp2k1qiq485M1dfjxOTr+LqDRl6ayw
3FrqeT+EHWj116yK+mGpgExs0Aot03cYKnthNVt9fu7M5XgIjp+zzxpJ2W2lF/sF
C7qD7yfoKYJtkgZ32nlUr5KjHEWy/ytFiLB/r8rrJlqkbGrXHkBty0IjRxVgwyEy
k/5OUPfXewLByz+LXNAKq6pQdV5LH9j4rwC9z22cRXOJ9C8hKf89BWG27ysrTX4C
4G/DAQvS0o1nwFhFbfBKexKYAOJDyWn3OuI86u7h9yo3v0OvEqhPBMvXmPor5/98
8K3s+YESWq44aSj+1YF59oUg7Lyi2qICrl8T8Nvrz+rQ+1DGphK+8vZNEaoFV2fq
SUtgvYeUfQHhBW4LjXBxwO767KrqCGBAihfslsR1bKkoT+OuuE3QSVuc4AZGIHnZ
rGUTeYTtN2jqCZz62t0lG25d+nk5laX1sFaJQl0SUb0FMnNHgCjZ61baQ9OGSJ+T
O6bQVzyyQ1m+F/7k6XFcDXywm5m6D1hpH0xY93whWChpfh2O5mmALsT2LB5tM5Sx
KkEp8APn7SNBXHo5/cMNoi8gk6yUTWFtPRhnDTGeHeyJ7uYEGsLSAymJf7j67rQ5
bicJlYHbt9YQBaz/kGGNBdO93O+HCtwiZHk8fGXM1UrE9HztQYVnga8Sk6wCTvyK
NYhD+/k3Hbp3jlvf7iuBC3oSXo6RCSeDz78TUTPuYwiCIMpEG4DI+VzbIndfl+ly
ZfjctWeJqHDGQ1lBoEqROgZWrLtDzVo6nenaetlEp23xH0cDVtIstrBx2+gRTFXd
/Hug3emUNWyv1PdakIIMw1czrcTZmhxes3lNg0II+xhJkMwx2epjZqPZmVqldeuh
LoHQ8LPA87skfrOibhq/LHi17BU8/xkJM+H35ZBKtwuQ8oJ5+GFtufNONQw8u2oM
agbfc8Rux/eZG5+w1syaP5bXNNOH8vh2ClHj1HGkox1nW3NhcEeWDWZXVONZ0ig5
badT84zsB4Rq80m2zrEVSMjLrM51VtJdQ878y3ywwa4P9E7xrzx3fcMppC5bWfrp
ARCV9FwDeZ8Qlz5RfK32DFhhyibbDklygGRuHFQKvKaF31MMVulSLFv3yyi8K9Z5
WDoRlQs0dXq31lbrWcgK07kt+5VDUV5oygHI4PN+rbxDnZ+flahrpGuhtBqgD7es
Tz59ooz55qtf2PITHkGwqEshUKMzvpFHnueLhIYUUnoT+0uZ5eA4h+AAiRYAexZl
ew8FNlREfprCu56DyF8f4aiToIbhVePfUnuzAzoSqtxPYyzbZFzMphw/Sk0Zf5BM
sF1wMcXiM/2mrvs4g0j3E90V0wjCO4uyV8/iitmsPnrOiUr+FCLm1i1JfKZmq629
JyNa+FweXt49xqElhhtPuo54gpmAN31z5H8OhWcKTVea2yhCcIzPeeVnaThTrFP7
Nj+gBVFwCBP94+8svhzxhH3q2sjBB3Y9eEQ16fXrvEIBAKqZI6PuDYEeywQ8XzfH
fI6jUP3yZhmLFORjlYJ3eJmphfuDOOGK7lsrfKvLZp8rrBVQYtRNPt7UTQR1OtCt
HU75/bclTAxF+IXs9yPaAnmVMvScEDL8DBuZwkvyT7S9oMC4iZxfyzQPd2bPFKTZ
00NuGWsXm5em8GhMipzYAIX+XZUHXfUgnn2SgYsD9ymsdn0uavOQaComOPr7PfYz
5OAGoMfr2geJ/e8ec4HCfdndrxe/ZPVOTp5hzfROCg450YaG5gfYFYokIdWuz/h2
9jPmyh76EzfwFJr6SAMSQ8fVq61IQwGcRgRE4OMa5+pQyU15putkrhFKYyt6gWN0
XC7M+wCvsfczGzVT5tozAEsaZWb/s64YZUinKNkWth+91d6ezFFWXD/P/M8y21lH
UQ6d0EGv5ZcgmL2100D/ickrzGRCaD2se5iLxs7rqUBhBRdzl8GzfGg/na41BxFD
gcB9XsYk+bj1763qWTFV1YZPUbZCr7wn+hHO1xoMAPq6zm0wEMTbI+IS4xnZvhRb
82Wo09Y3xQJW2qWFApOwDeKvzn+NgGaXObrLFk7sVnWM9PLTYtB0dmmQTzYFmUpj
Ns8V2a/4T/dj/+AXMAqD3Wqo7qGuzmmb4F8TGQXquDsRvaf9xrQFNBTZmYXoHzbt
b9l4XyOfKIXGBGcu76Q9eUXO9VpIGEvpxTd2oimEQbyFor3c1FMCxyr279W2hzMe
+t9aU171OIH2tKk/lL1CwxSGa4SwD0peh1La7BDeK1Q+qwEm5PRtGIPG+tIHKgAq
0jSY3VksPxFv60t4D3fZtB3dVIH8GctuXsqMM7Qr1QqLgYSguc24Iy3odwnvOX6y
o7BcsqSAel4X3pTtsHFKUHMCdjcbQTDNTqnowSl2m3ssAtLvdg0d+r7XSchwUDDG
S6pMJnc7RFXmlmkudQRfclt4bvUCV0iq+iJ9Eet2B+lYI6hIH9YsimhOjGjCDnm9
pfEFBIz8JwJc6unpcYjiXP/Xm1bm1Y3J1vhtG8mOilVaa/qo+Ixwnhj+B7eVp3ZX
XnXl+WIbzPRqQ6CKD0gB2gwmb5w6Jj3Nze8n+y01iQXUzKHei7qTjywA/CAziw5O
pleP0RHLt8lkmfvVk5R2XV7AHxaLsFOo1wpOteHMR4y9l+RzFhfdzZATJKKVoJHk
4DpjbR/J5XnaIoSxASdmb04cnBZE6Xij1d5rAnwqsaR5EyjG1sXHYT9nJggNcILb
kczPnB0GL8YSeiEjEulSqPX4lO5P/FszobqM38KtEEtPgXjiO/QvV4nVRpeBM23s
yg3L0/Qv9V/y8t6ScbMWRnSs0J+69cZOJgStlt/jap+bX5lJpHaL+TCcPRtaTX6D
KMOl6/hRkmVO4P+L65YzSbci1h+vWMOvVyCNDOpkkXMDAeC2hgw2ltNZ+qmJrGfP
Fu3+9Jug2+XCO1J4sezKYQLlbddYiJsLsGo3RyR/akOeKBiOit3R0oEFApCT989R
FSNUde2MteIoO2ZCewz7eFbnK7fKHkSvA/sIsSR8lKeHfjGAvH2bqcB5c2x0gg5U
+7V1gYFv4GKHXnR2Hp+OZ9at1eet2xe/3VpkbXsWU3IZs0+YJPBlAABNCrhp+MLV
+OZHDXRTMZFl5FdP8GLdgTd6m+WACyYE5oVbSAPWirlPpfcoaKFolx3+bRWiAC3L
BukEE70aStPRkNvuXBHwaqgDHwFbcZ4rBS27m8ki3X77DI+OF9D3HB1d/jBT2eU/
w6dtlmjyFMtqh01ibowQ2X53TtNfjg075xVrNaO7zPHgyGctJW6mKAVxHhMZxgmo
n3XuMd4KhepJXkQL54o9P81QGexGJk+IeDcJBQo1IHA9/Em1wMfL3NkV+2tF/3gC
DV2iHHv0L9FRQM67EGYTurwBSs3ND4s0EM5q7jc3V2fuxjK4SsuJhpDpUEhq8BD2
EveYeGfvMQETB1v/yetAM4E8SU9bsgwvUtbZoPiOYjBH98orws2vj+tpB8iIoz7s
wTbPkiQa73N71eaR94z/f4B7j1zQrBq93NZ8abvYPs2EWiz5t3ZEuWvm9q9CiMKk
/un19y8r2XroE552Vx6QH647aARs4OuyX2YTa0WRrOhJeCAiF1bd4hnkX/OiCTUU
0359UZKWSUPpMFHKK/aNvT5q7YdkVUArTQxYtAFrFdqQcwAmPQrtWmpQ+64USEfG
Jgns5nJrMfjM6nlQ7RDXjs327F8OJdekiRZ9SVUYKbzJDqBNU4pNnS4+oP84p0XM
7Kcyfa3REQjg9IOCUNUY8XEIzVfGOhmTWrYDGv5RqV1NSmX+SBkOmu4HupQnG/fC
mGE9cDHsQ/5zQbhZbV0fZBPlcg3Ly2mDI5V2mhLCrWoLWSiJl91abl5W3YJERv4P
zluQZFUBZl1p4W2G3NmKKhG71nPcbqT2TaTzqEky9jhqPJZiJc1QLUvyx66riHSv
d6Kv21BjRTK6m+61CMpGODt2KAcM7jlmIZgNx0Vu1TirGZEpXvIWOo1rx0UbjyCA
ZM6LgLm1KNzHVycCwG2M3pJ2had0qyZ8Srg7ITVDyjnoI1tOZZEcObDqsEQHCr36
YctnU1ddrFtsz5mjyTs7HvgF2JO9O62qXolCwktNEaHbeJ2y3eFwGu2xu4J4ouOG
5uynJZ9hK1IzDQKMVwIcLb3xWJ1saUNEZSIRw1xUy/SBEqCqthYxs17U/Fht14wO
cRrdV3NGodUvJS4U7k2ccICMJXnS7xE2n23lrLUsiUTDz3uqUtQNfS1S6cCoUuAX
jrDMtxWXZg9C12ia06mMGxHVTmeHuOl/Ay5q3D2N5qd3bN9DUyQlIewkdOVnpGJ3
6K5U+m5rD5UVVXkrrlQ9M68xK6hYMcaY0N33XylGB11qdrB85lpdqaONd0v5wWvb
Rr4lFG3M6QdfsRdvlVPKOR3FoqmamUZa5ZSHPPUAgIv1rcO5Ahu3ELFPghLtBy75
iGciID6azNosSZ7zwE1/1MtbVgjrP7WL56rPmDhDHC7vuT0y0XblxbyUcoaFs3W/
mcdtfTgImSoQL1titMn1AsgKyw739t0i889RPdyreskIflzmZOLUis2d6hNk+jXW
gDPt66ENMDByRvUvJPA6Plyg83tbwR3GqF+xBNonWIL6Oj9gXb+bLmca1nQ7hs32
GozQfgohOJoohL8JAXXMH2CJTvJI1LYgT/2LBmfq/VqIAqfjYgVgapsAbj4k1/to
YGenglA3xzvkMqEs08Fx39eZAC3GWCMRBOot/BNlAG5j1sn+2NjS5dhIaFyEyLpX
W9NJK+Bdu1sJMmb60y+CnNUI7fpohSOhWQarSwUj6qXhRXgj6qb6gdCTvzZnTsUa
UiGkV6bb1iGridfzHb/2Ri9sriSKsDgTb6Ag+EgyU1Cnpevh+bbW/tju3Vm1mwC5
OEfmTRX3zRW0emT7bfj7xHzfXJ/pOEi75JgzTphQZt0qx0MLdbQnPhisdCRVTfjT
DG92DDscXa2hiVuxcZI95aacnf624d6tp7Jq+GZT6o/EaSLktI3qVdkQ11jvvsrG
fELvJwesZpJfQ3h7M72oBblxuz03uGzghMezKVE9BAXxUPmS9yJgR4cPvFqob0eM
nJYlVedkigJPz9xV3XlG6fPzk/w+lGQb8SR0uG1b6CFl5bCKlyKbWL0lqr/nuZwQ
6lCVlOFoxmeBtEd835gZ3N2jUvCozkHZrBCcs4LPCww9Mtv7gYOq7y/Imm1qok6O
sdfi5SG/7WD5HCeyAFzOwkIGtsW4x0REGtlzeABKrQFBEg0QR2ac2qiWq/yRJ6j7
3YnasSg9eCzrjUyOoga3adNMHVis1X5U5BitEXeOKDhinBR3ubvgI27KawqRFsuB
yAVJLxWkGPoInwgydK+9IwmuIlOR/qrju4rpwfTXM5tc63x6vJ1TV0uHIdDEnjG8
Gmahy/sjcOkrgHMm2zvyD2Zu4XoED0z6ri53s1XVdRmdokZjH+WZ6HF6TuYEIiIY
1wvNHXgnqgpEyUGOd+XpZR02xiETijfO2PIg2OXxaZWhcZ0zdayTRC5l9LujiwKp
6UX9eB8oV9XtNJ/uWI3K/SPQscL5E5U5G7PTovkb/EqwP9ed+cNxCA8eX6xrJose
gFDoD+SHc4y03snXOxowIMjfQnrBetVsJEa1UCcRaX0u2BINUKpigYwfjsQQR/pH
87WI+5GC6qBhx5PCTdnH2ueCvb/B+lmWaXeap4Q0/T8F8Zcs6wuJqoB2yYYBA6Ze
uiyuZTQ38FqQPa474L4MHiMhAPOTSww7ylQJR8GmD9MPgO0tp44fbhTXK53usLAj
wBW84JEB8djmj/vMugSFf5BcelJ2VyYL2/4UYaZXYFBLkh/ZknFku3zZQee03SMC
JgmD59WOVDHQTgSOuRnR2VILQKhb+VNwGjuItjAm1hpUMG0qpmZYGb6pBnLAU0zc
0mkLiXEMRponH2BqCPWe6Q3J4a9X8BBwz+ciWBj0E/hM4YpjTKFqDfQKDgzdLG8l
CgDIhvijzEMP0icdhQIGaNVBU5EH5QCHByPLr3u63J1T7m/sspb511dgonFeMGjL
S/dwiy66lwuY46xyJ1UnJjZ/TpIVBmBRaf2/jxs6tF0EhJsUSqL+uqppN2cJsfrg
s8BuyHbDyGDIkVghtk86+lZ4VUlxnwIXHCfzjA+PVEpWPDWeLrpcyBcOR/rxd7zp
iT4+qUij3Cin6kDo/VVb83+BtIE5nU3BfAAUQpjJwyj4JbvwryTv3gkV+S7ZTno0
bjPBj+HPQkd8yZB/2WxhUKIuKsAvEJ3tFh/pVpF3CxfHbd5rxxIcetTJaYQKSXcO
jgLAkJEfQ0FaKX56136mFPikdPhI2J270kBKx+1Bn2DJw7w9ok2VibaAKI9xylQR
uVJ0yuphtKvci/Y8IVBsoiujDnEmM1Q6NLuuFuBYNdUicrhccCtVtphZOLQg3BXz
xAgxaPNcQLeggAC9Exhm0p+u//DY+P0SeKvEFo9n928A5IoXEAr93zaZFmUOXtL3
NxhrHUo0elhWQv1TfvtOcN3mg/x1v6d9JtbjPWg9MWVK9jU0A/ZkFFwijukjFByP
ulZCaXETiTO1rLZ2cm5EauFvttWvWTFwIWirTIMcyS+DerGGZCTeLeeZO0JoUkvN
puHUKQLckZ0Dg8uA7sbRaKdyvP1pxiw8Jbb/C+1yUniR2QrLX0atR0Py1rxnr+nY
OUXgQWWtmaHVbUzaKaYxNV4pkLDtKSK0HkxBdIf1qFlt7ivEWHJTa/9Y/g1OmvE5
8rqVCWIi10cyhtQWtHzN1dvC8rVZ16XpkDcqyprKmArUBDvEK1qs2v27cN3nb7pf
QLWAkH8I3x5MjT3QigAgJR48Ri56BoOpyH/W05p/y/79qMpmWgPPjL06lSu2Ihfb
C0Ot6bCY1ERjda49Rr9m6Ism+fgrBkd1V5kE00vUMnzAxJEYNV/WgrHHkKXlEncf
fVYJy5LDVGTcUzebx6HxRphDWtqIWgGY/ED+O8m1lKCfZCmqF3TzmimTA0cZR52E
6cA1lq/IAefnDCeDBC6rC141Ncxlr60tEs8I+/U1fMbVfuRRal3rRty4d8tbgF1o
TgVMadH9Ztyb05yMp9HV5Z0hK+pfuOszaKKdF7vmAFA30WajvNaoQ91LlfgMvNAY
9FwOfzZyVWkzdcpWAjMBDeVAFTwnKKmN4R1be1N8HbVvDyBj8IMhQstfU+sUik7i
6fd5iQbXLii1e5Ybme8VGDLjQWxKoKmOlBeT4s4UFtN9BOBme2Q+RuXjIiB+Uh68
FrLANQo0IARL3YYxBrWaQfgHwsHFWRsPeO6CMXKZeM5KmqdnkhEmlUpsYcnd3b8I
+BN1nu/kFwFbquZTLaOSMKkL8DFpB2y85oVMmmN5im0T88EYcxu8iXRlqivWZPp1
PNTOMB6QK8WpCt89AoHLbhhSJ4kmD5BaGroSnCt8crQXUMGteEEcPnZaDhx9v8s/
bq3UdbxbcE8KlaYF0yNiCd9nDT8/HmeZBKRzngyg/4vQBySDRJzRaUB+jUew0D/i
HZrHoD/k8nf6WgJSKULUKZCdALOeu5mfNNb+QmxasUAxNyf6stJYrjFkcVH9d8CS
1tqjhbqxCZlswYGegPXyp8vkt1AIFCL4EcewmWboaI0IEc9yR68FdaU7AcC1qo7u
oWerna00v7irqveFKoTDiA4i7BCkg9Tjz/PCedwWFqN3LCfaSPgxAUa7+xETDfMc
CUeTmLZiXKbUDlk/Za3/0vb3xx9q4Xkla2eZ698Mlkz6dW9DBmXgT3dwsYyMF89h
+iocFjcc01dlo9p0yPPrEe6ejYFgICsHw59Jkhc214VGYzTg2kxamB/yjALCzs4A
r/WsRpgnjlwPYW1JgD5FLsn3wNNdjx/GYKMoxliz++54b7srWupnOvrSquFpPl8b
dRr23ICvDVkOGpgZApscEJNtrBithx0P5sZQCpgdGUlRPuEKZ+V4GMJ9D6lONh4V
obZwmPD6kQusnD3Xnim3j4/Jo+B0dd6rBR1/uY3R0xW3bf4yfJPJqKmQ4qnpBgvi
k0AyGiSrDG6WsdS/JIguSi44xyN8gqBU3SS8uSFEBtBxh6grETNUlprb4ewSoOOR
8GOSX2GP9meXDrpoj4R2q8ao7XlVwgdNOjtpQ97sqEzXd/9ALA9UnWvi2s7GnR2R
5JozWr7zKBaKVitIh9Y1xVN/SxdpLCvmRkqhP1RcOIhpH/xpN5b2/ngr7V9jeelr
cLyMj13cp4Torq9auG8cFLH3+GVWBZR65H18jpp4f/z5mVBvX0H4KmjDOEpxIAs9
oj9gZF8pAhUWSlCGKtgboVV3knB8euw9Oj4wybNWEU/RBo9XM8CWptlD7TlGsZEI
WU5KD7qXUB/60sDGu2WIHVVnVPn7CRnYTgJxymxGgJ67qqz6C1MLlgUyV+Cc7O47
O6jhW9lOU3+d747odIf+M+0hN7MxyUs9DNjTtdmagYtm6V5awf9cNEVrOo5p3f5K
Jj6iE1ixcQKziK7fEQ6l0v2YbdHTxCyRiu/FJvpQ2aL/QyhIdLZBT96+/ZEvufi7
VC1SfYYMJ/rPLmT/pvZ6N/88/nd+3jPlVQIpw2o9Gl1J6SWYQtzIOWVpZFzTPqM6
ktM2PuDV6W6CTVJPmHfcUaCr5/lMSo6aDZ/uLObIDF5R3sbwKvYAN7OnsvihqtOk
BNrs+YI7v9reCBVYxp/qdATEnYjG8pStNmOsPnXHnbYN85F5XxliPMG2KsT2DWq9
Pzl/2SVm02RX0QQoWsSJ+U/tvxoTQZJu9iHZKOJdrjhGtoWKY/O229q1EoM/t7EK
64qQxUI+ytB846+RILscJ2jv/Rj/zVoxl7EcGePj62MXKoGyRoJ49x9J4KHbva3X
fZtBfzP2oavsJuq50duBlBpzoPzmw3PLq39DygMxo1Otg0U6K0Zs7+7MbaBk6js7
/6TC6Wuj/TUdLEkAzwY6j/N4nUG5ZRhvfAi1tKMmIVuaCmKrXgMOTdHS0PZfbguc
S2b29tAX2KLtM1Mp1pbT9BMVP9uzTS/W0sSPPTAVUr0zfJwKHkmWOmcnxcbo547R
KMq0Vz1yY6NHdPIXHyg2AhjvVHjLzxyoiqtTjMLSd68kPmN2rHwRe0iTNa/PtQRE
FCqhEK/IXDjxwV6ELyWNI2vpKACduf185b1aVwifbWLiZYGLXr5vWSxa3iCSoDHz
wJy5OVaf6Z5RuIQTd4POlalKE+/nPDJG38BJFfEgYrpHki/KXU5LIzGx05A+u4Uc
26D1SyCSSX8TYZcWSln1nEw68P1JrIcKfupALqfE7zAK6HmN6gqzGw6Lk/l0rM8F
WPgVUV3AywHY43jfReeznM+v3RpR1hi4/N7R9RwlLwlLc/BVjk4xwpjrVvI3bT18
5beXqYEGzZ2noUqvGyKfbMpg3CUGClqvFBt5Tnczpzu+xuT5bO6Mt7AA6j6NOmNc
R+y0cFPNTlM/XR1yjRu/6UVKEXUW3EH6hKfulBkcYcP3Q0yGa2sJjIKcGENAEx7L
FpGxo5fHZqx+Xr2KpptYg78aez6N83qtsTN8QFjbjTsRXwJX20pGqNCUBMsZPgjw
JsFj/nwyTe24ktSbuPbNXbc+I5FKm+FoCmq2jB8r81+uUJ7IyKN5RphNQFXSIjT4
krq/V5u3qrKID/B2k09lZHbueFRiPd/w7iV3Trvmf7go7In24yMqyNIUwsK+ZRh3
vgesdvIwamimXHqhYjuArN5rrSs2gsi4emH6c3H73UWkq15GvT+SzCZ79wM4jeJ5
G5Cy8PV9bY+Mfbtl+MXa48ZOHMe7vNcx5+vH0u5ltVxe/FAsdTb1j2rizmj5zFvZ
O2xDaxe4l/hw91hMxSkwJbreFGRzIqM+FG+pb10WlfOLkJZ1EQrNs2baIJOsSU5D
5U2urnMo+7bAJ/VC1JtO5JzE+6uOpYMVlMiExDHcTc8g62puRbXn1YjIVhKt74Bg
M/c/2K88xyUhzysOpyVIWmCiHyrqta1JfR+Yz9bYUB8Ta+gzBfNl+0FBDRZUfeew
e80suK9kTbN+zxNyipli/uolnpuI+ISH/Dhp2BIbk9sF5FKqIoWdCsbe06LRy8Ja
u999rkg4T1eEZsZoDQ/ZJcL9Z5JHs3hvGJDmoFXfXOd21GCAkzCqekl3sUbiWyjy
yfC21Nxr+jsCHqn+zR3eKwKILCrqS0Glx4cYwsuz4fJ0TIXUK+rP6DIaoSNuQhst
j2e2ApgpGY0FH+lezGWwXV+Kj0vYHJwl5NjkDZJK+gK+fmskq3XeLjpPheStB0Nh
tgJO6cDtpsT+djTLFxVPy01bKnl+8T5ycuMZSsp3CiRajpDExqQLWPWBl0KZtP6Q
I2c6gHIiAG93z/qdK+uozG62BcWXSLJizikJ/c2e++X1dig7tNIe/gIgG4S3nNdj
mm5oI3uOx2TCZEyM9763WiPsWOOZFA57GmJ2xseH0PPI+bJg4ge+WopMbPT7eeY8
eKKb82C6JfDUmYetxopQ/jqQo+EsQkj3TRWrADPVIpnRqkdz5714lY3fjneVTeLL
cDxIv9OO+lqrDyvyrwR7s3b7c07Sn+BAFytX7Hhm9wtM/tiLfQXwI8xKxoXd7ROE
Ji/Gl+EMfRY1AKwJWWydgDQ5x7skt31MKLwiUM4COxhHhys50Qn+aHTPOBIhGP2z
9uTLe1+OZTo1xt802X7hQTuyBXc19crwECcGAwEwabZjO5sL+rnjNkTNA0fJO4x9
vGJUzqEjrteSlGc0CZ1sRo49c9MDrAzEpcnjBHdMIT+Y4RBMD9wUUHAVsidLc4GR
OiRftxRMf2R5tStUp8dtEKB5APwY6+N1Pj4pBAMhCCSMdEaDBXNLuAbeT2VsFvY7
UJVToOmGNH27aaNFjKu4ELQ4AUuH0Lq3c6YIgbztHuqRnMy2rykDTQqlBQLfwogi
PNsjbSXaWh0uoLAieGmlPUp2LOXkyc7DI8LFjr7/fszvRvPX0Bkhb+6QLdFY4kss
k9UOfDb9nZLeaR+1FNAKegmkuOnwfx0wKG/UzdsZxnGEwIQNFu4LKJIPVu6h7I8g
uYt4l8SvcDT2HvEZgsnoHVCZ7QzPXHQS4aEH4I/mYjJP6VkMjyIFmfkCRsdUV0Kf
kcckSwOvggx6v2Puikkt1zFVWe/zfil3o3diVCwe9vIp9pumaC+Ue8SX+ahtSSfX
65yD800XTCQAKQSxV2nZ8BQoe0KKNnVg7bfzY2NuYhDXLguRSQZWftQ85BblqHBH
ZLjH41Gw0zKx0VIjvke1Jky0lRpbwOujWcxbpiCnbYLIy8U1xDVOe2kQabC2iou5
HyN6GAsQjf5A0RUqfzFZMyfzHxv2MKnfAH9gx3LWpZfT525skMi8D/EnA+J5QHmR
tZvur1IyB9H7VuIg8x4DxdGqn17wxJbaWkOiV8xGaxC+dQkJr4GZ2fSZ8gZtpcvT
l/xgDEkZMtxkCAL2NRRGGwhQf1SbvtEBg/pTU/m1quV643G3c2pKH/t09h6owedQ
u+FADzYx075WGvyROqq9sT4shgqMlgQaIXJumVu5EvZtRbplQ6E8093SFF4cD5km
1cAcdeALOBQ0q8aPDPoG8sR9SKUVei2zih53K5KN/5x6vfgDakRPZnrL5VHQZYVR
s4JoR/4obQyz9QVEA9bocPD15ZI+JGTfTqj6ZmMnIJEY4FEn30hjHgMYd5flI7af
SJu9cEtCv0LtMqlD2WNvTCtmtS0fY5DDqbC+dFVTGmN77KIIvnA2yruJgmbU7zDx
NykiXC+p+pvcHFMcn79ua/pnDgchQLLJhkOkMwh5R8A1rjjBWGcPgEmkULVDIrI0
aeoq+OxWJo7CA046E/lMYKvhLWdbcsb8BoxWhmgy0Bp1CwHa6bsB9AJQogQJeNF8
21zefMRysYTesHqGUHL4/MNkF5xNidOvvGCU8iIz5yLN0c6bckpoML3spXRueP2m
MJCXvLqJgVDWKeqqfjhkpQVp5h7xegwxLeL8iEVHjjRLr6qVEdVA5UYquTwSel7E
UMZ4UtWJzx/P/T1NXhHgK5dxVKdbXSVn+QmAnbeV3Ba9fnO6HIEeKvuiVncJMJ67
WDztrd/k/CYl6UeuGbvFlWHd3C9JPGN7IvpVnotilQTni1veTNqJly1Bg1v/2ihm
o2j3GaXE3MB7Nl82KUzmRHmmV/BKqpGThBaRZEiobPVP6sVnxJm+6UD8SGtw29uD
r2VbqcRfZ22kdAxrVNt0JbsLrGKylRwmpP3FesPmNDR7kA54rmnbcSqjLD98ms/A
WQ3mflDv3HQ6cAK0NilUyF2tWdPCoGR0xL9KO3EVTjrMIPsdapalM3tNR5WDBI0k
D8WM8MUxG3ZbJWggtelrb/myW1HLazy28xefNZ24rs2uuCc2GUCopGQ2JO/T28JY
4pQR9josuzjKEb8+d/aAYitkXTD9mQqXEBFwAq49nfujBgNO/GcgJzCH1ndL1EK5
mExlqHbZG3NzonQlJ/ATS2axyPvRTEbJ5iFD7rFphLolGi4C7X8oW6NthYgAeqo8
28d29fc9LiYodE6LSp73H8DBO0Y3fdXwBvvl9VJh15pE2W4Be2AcEWeBNkxX7zcn
RvjIaGBRmwWosq/6PnTiKHzVwAfwIBZ5TL6ERBkRo79919MqwqUHi8htgaiIMFqs
Euig5w3gWVKJ6xhAqVgBeG2Qn1bHLxWgIKpGCVtZqLlmogiyVIaLBtpcqAABawCp
k7i86nbHIR/F6KxMhlD/vOkm04YcQpiV8TPwW+7ZR4lZcNoo7usQKAw6U2+7CNRt
80pomqjmjyYOffVwd2/3dW30gpVvFhhLe4i6szp5ag2NdXe6fl908m9WGdRaa+x4
bRYr+a4Indt2MfkkeN0ii1HZ9VZcLPPPTg6/BEcCKvUp/4NTTm2TX1dNHVFiqfx1
86CRwsbh1DQbpkICrUI6cWwwaaXadrgxvgxOgY3MZsxV1xQvF62+hYA7OeTUCbJB
QKfY1YCh0G/KhBJcM1XlFgdXfOF2+4sJqBuTK1isadAh+5JhIIwBg3C974dFTh2R
EO37r3n4ia1+ft/fK0TWF6F5gojllQbixcYq6DyUhi5gzKwaeB7SRcWDql4cAW4u
tS7MmXinHDUlVbck7vJ3wWcYvGrhhZ/vhOUSeJTJ0pZVPQ9U+QqFwvqZYWzt8FWn
2h6f8SJO2bdtRuljX5eJUrEX7v2VBdU8rVvUFmZ7cb5EUSwEYxnvLWgScWN5JdYm
TUE4RP7KibKD1Cr/TnyI6zANnJTxvo750u2Z6H5biSzLJ/iRJ8PgaVADBsD1VW72
k1mT+mTk+fo6U0iUF3y770gatrEftcfkzDdQvaJacUseS5uOZdYgHHgfqX/qUkeQ
7uTWpToQELu1PVVKKPSjgKXjVE+HOm/7J9B+qL2WwDo+X/CFb0sfzgRp4DioF+hR
DKoSROwk7m5JztIsUYDgeifhh8B7vbhL5nIQ+Bwami8Mt7EBos6w6EnrqPclFOn7
4oqQMizzn+qMGKAcd9LioeC0sl3zeAUoRRWG/UEkDra9fNvL+NIHYQDL/VRF4Xlv
VMT1kN6E7O6OPLfqBsZg5bhy/jeYF5q2VmtLSVcRUcIi/aR7g8V8I74WzHtplnMq
4VuLvzviw8CpLNphsw0CJ6aLQFKdRlLVD9NZL9GEktEvUWqzF3Ghahc8b5xzDyrK
1TVZky8XXmK+ftWY/rd8zaL7/RfcGT0Ufr3Spn05W6zjn5GoFArYm75Rz8GMj0N1
M3iHu7fUbwy7JoO2vlr4gUcMFjEfbdVfiDtjmWF+RKUqXFxYcp17CtBFlXfiCLZc
fpBh5eqWs7lk4r1Q2LwI8/THsnI7WX7Sf6qHa9KHIdx2F9FJMtEwQ08v0W613yIL
esBs0JJeUbJmrE8kyiU6ZeNINMG3CfdxX5a0f5oocESUThOR//rbxo2Yf6lfcM88
479MUJECuisJh+OEypOXW7WFctmLdHnyN1jk4sq/1nLrHDGA44lvjW6TAWu3YRQm
Y3FWhJyxsT9fPgINQiReHhqE7LuiXy8TPE2TIhQYWco/yUNc0nXsyOdXfJUjvazU
+wcxtzduPmLDLw/xGuj1APhxPR7dBfDjvakioEQglo3keug35VujjAzWgfXmxvvc
+47tRuC14WYT5eFdfTbURxiZJjYdrj0pw9VpQ+zQg+xedxNjrbOaUDwm1i5g5rxy
sjbqGmbA07H0hGAQ6Op26Ae1zcRbqW23DAuFaQwC1o9FNIdw3AygGIoppTyap4Kl
+JZb9tOjEUT2clpOuLa2eKBGrTuFbwNF7j0EW2Sik2csy7uGuSKxCwivisUQB7Pd
MT5cOeUbviQ67CdfyvqtpKLZdyMoI63znKpruy/fz2F/ElN8YOLKLBDYT9dzxm1f
hMDjXYSgSDFaQwetfoTxJRo9I0TNrxYTPtnrugTkHkCbjG14t2eEsNQo8FetXSjV
CndUOr6fVvYV9BOaBCmagea92+9I0CXaeBNGzdnm43TpaP37cg7Bf64PDJRrSXFf
hEJ2Ix43v4PJ0siX5UxpwH+6dUQs/FaYEc9cjlA3FXTpl+2JvwKOH1Bb3Nq6Ds0N
UgelKItBmVHEolrxFeVsALTfyXk7wdqHtx/QQdmOaecR86fKe0Q0BSXwOPMc5NzK
5x1bjfZ2+TWaKHkfhD7Bb0FPQJjfAZfCTlcQckvfPYAgyoKB27pYYU8TPz0Zdnvm
4HjfzF8rRBQU4faTMC6AADBxPsQXF6WWQXttTb6CCaGOG7cgAbrxW64rQiRwXNgy
qUr7IA6WbxBiWTLTsgz9zjLPE/rTMOGT6UDL305aHlisMauHlzO7GYYZNh7xRlLM
YjEiX/kOnKwniUPJ7PQnxXSRELBvZHl1hpXdrRgy0j6jcH2KKk4IUziedG8uyvWS
og+GYxVH/Nd+DJxc/vDGjKgJWdFTBtdngKgYaixH+pTtACu1AboUxXM4/raOUJL1
jEkCrii/qv0DLKIhjyU/Pl0Ux1Am8Vvfhrzse9Jy40ftYh5ENXwC4huJ0ZpBbs5h
7ATuJTbileE9wJ6YS/cQ70Vu0Elkp7nwuufF5W8e5z/WOzx9mqTanM78/lv1v0Kh
xStlXanyJBkCvSQbYcHW6LU2GCme4bP0DGM80pZBnR0agGVy1ds5YZF+e+l+wom8
Be2kesJ4gbz6N5VA7hg+CtGqaiLRBthUU9SFLqLZZteLbp0B7N8q2tOkL1gs13wp
g7deJ3SJN0bqK351xJww9tL1MwYnxiWX12Z0h9YEKUgVDOUegDeVjOZ4jDUIcJ7w
g5bXfgfd4LTKaUKSI75oVLodbETygMYeyRHbLeF7z39RVb/qbqpKjADhukd+fL/M
RKIJX+IpjmvcQYxF3XQkHQf+CWcC++6smNRiuoSRVr45IDM0mOCHdk8nhmsx8Y5B
CD+LfLFxR2IgIBB1tuLOSA/sblCXDhZ75N2NaCribctSCUCvaI2PqHZnFD6YPK+o
0CzZ0nr6oOMpnEH/DltpqGvvwmSjK11Go4X+JkIo5jFAOnechRQMiFcPeelhbyfr
Y2+UBx+6OPZKFduV2XjqZfRTPO3Hf7D9cJacYE4kQH1g9sRIla/r4q9o188gupsl
Ff59KlRhd38iJLE3SMcAnIkgoKb+3gtermAqbUCNtlDvZUTmWSFtJ1DBhJtsZV6o
qcHBoaTs6KOPzVb7fKebD8wsRtPztWrhknEoBdo9wUAaIK1mwKSxZf2Om4MubUu3
USNsARMtPiyFJu4/6DXKjWTtCUq/d97PbKtvbV4AMLdaMC9ERMhUrYXloEVU18ZX
ev8x84eJvBbS3cRBrM+jk1osE2sLIMHz2gRqBovEyW2aiAG75+FdMxnTdSojOWf/
uGS6y5+UXDCcEZGSVRwMXnU1NZ9g1FBfq/uB11cKqstcef9/n8ufNNoRw/+xWIc7
S+9Nn/asSNjV90wObePlS7tIp2dRIpJBU/hV+2RGMOmJowv1W6YzAaSHMM5Fxio6
H1SUsh3BttmVxy2uIV5q/nT+PWGdpfGe2px68AvEgEMEKBOThfkj4ZzOP6F6WKa2
Lv+K5NzPAq15XYnejRZnU7bWnT7W2AQKqvUy0qS0GalQo9GSiO+IsKu67t6lekqp
BI+JE0XysB82QFQeWQicNRka8G1xCTMAKgqDQiztCL0egTx9i4spwnVou2g+BSik
rTRotBDkw4FLo3g69oIs28Oud9bINJ4BRlM38eIUlqeaK1HnPjfUEir0CbRcIkMm
yuu+hIYywUfPVZSnt0hk+dNENw4LymBmCjltP8apHNdDLSvOeO9Ic6Udq7Tglk7M
S7MVm58hMhc8r4SqX3JOKWNS7YG7/ouzHozUQrWcVl8ZRECqrfZzIvJ7gwmzqNe7
JfgJfaiEqA1QQaEt5YUn2yNwHwUv4/HBfma4BIqDzD0DiRw5HPfbTcMHOnBNFz76
O+yEOF9nvEqqBqIzWQ6b7OxZmGfgbMnclIqgrZLH8ToXPdrcsdxzo8kmLlUj24ag
VVAQbrkkgWfI5g6MvQVjeU6Vc9HlETqtnG2rYxNasiZRRf6cExIxqHyCLaHY52DJ
Hp/7rkpsHftn5z65OKGUzHgmgk3ItqFtWk4Am2OufyRk80Xb8/rPTx/lli1i7cXT
aZXmfM9F6du0g7BuSD0UAl4RZPWRaKb2/9F0gypfblu8YTAbIKd37J0eEJyEKqeS
jq8p6ga1Q+1GW+qbBAaJpHMsgcENkM6Auv8vHRKwd1tMWKnw9Z3ijfX45jqD/iWY
y3QgQVyTsmVI3pENd6ZtO2dusW3bYLkaBUtayvDP8t+BYpXyDH5s8TNlJzvsFrpC
H3vAF7J8tnrunJaMVnYY0qZvNJMcl+0jpZg2dsVRpKwF6vPppECCrJIhhcX49T2f
hP+1TFhZQvl5PQLyDscyT3fKwtdF+OLTtsucVHeq0FjG3mCN14Izi51SaNznaejy
aU4c2QImJtKd3uwf3IYn2akDFqP4PlO/ZdFuOuD13SjCRPUwpsQmPKeRuVeWkkJd
crtyVBcb3A3KaSAuZ3uiG6YRvy0PM0uQ2CyM5g5s7jbG75ckMA0BOcrPbgYuzYfS
7uetz3S1hX1PRZvcx1aDX8ErYZBYSX1rbMqbxSaqETLGvnGti2OD/dK7errSoFu8
FfolZ3a0InS1Ebqc2I9RiAKuTb1+MnkVUONjVImnTkc4EX3wqtY81qNR4U+gvJx7
GzXI2seKbCHc5EHTl/RdbTl4D3ScATEdjS3KVU5y5QM0vrgfXqduhkNQQUAkiBvu
w9VPbLFbHQRP3fozv0LUrolD73b7rbUMAGIuf0hjGTAyOUp83edaa05Q+l54J0S1
M69Q7Ex5y4cqqcHO2c4PnkILt5q1l/MQydBEiASbbrDWIVKsCPkpertHji381KTO
BJmktUrhNoowxZS2A75AKv10XRWmcBW8nEdwJe0zHRUObHVJuUKWNrpo0ahXInp8
Gnbm09BJE9X90aWiTUaOhICyw6Peqzf1GSdrX8AeTHrKfMaYzwYbAMMAfPN75Vsc
3ZdM6umzCW6nBJtrslQwMrnz8kweS06urubambJo09dZSpG31fodSG1Bcvmu27wg
oJAse7IxM745FC+6JrKwoL2etdMHVqLLEig41MIjox5AvunVdqW2hLu4nP1QPo6a
f706xybcokN6MSZsyfXnnHKLjaamhqwdlhDV+rheidbdlSslMBvXm5S4CIXYAnlr
RURyQlvVdTJHfwuqfOttwSxJjWJUOvw3lPaBeXzSqauG4kU5nt0/jFK1eRb5yaku
0YIiDD88fDLgRq7VP9vzzAJyAHLqWMYabXR9AyCU/TReyivsb13xe9tZDOXWj10r
tU8R5yPu2FOEV3RyE5bBBaPkHofFJifXfWxTq4V43Zc3w60MBpRLcCcfZBnfbYFX
dE6ziL2XEWg26tK7xBEExu4U1gbo79izTRJ4+DrXNrb1TH0FUtIUkmBCGZY0CYUz
b9G9hixoTeYQYytAgjGaRu6s3kFMaYSIiH7pIMYWf6q0zh0bZomi1UKV5SZh2Vkc
KktWQC4hApujVvScy51eCMMoSQURrJg/0Flk06eukbeX0ogELpvGA/LHtWMLbOZg
12x6BaGUjYUU8Nk9UXAi/oqc9NxjguMFDPgrC0n8rHZZOOKrP10wksYEFiXM5Cf/
DwXCLte4pDuwhDQtnxRG3oWwZTkpKrohPynNPE7e40id71vBFvK+IsxZUziboi+o
fptd6PzMUCIec9gG8x2MjYi9xqdulHk6sbX7u4Jvmw4XK4gGq9c/+rLyxekG4D35
55fgmsVgA8FIZsGSmjIKLYHvJmh80226KO1ESt8sM/c0pXaew7sYJR9kPUoq22Ah
NDVzC2L0DYrG/0aDr+6hLx5USMdxravYeBl2gtl+jwgUqKFqewSsDl38X8nPiG9O
6xdydspbyfBjo423f2xkgHkWpEolvFbJhw4fv3cBZgv8gKRUjfDITIrj6xDm3e5M
vKoqGLdNIU6Kwxnj4DZVc1t7fWpWALEbJ1ZHCQ9q3uvhhGjFVexdRlxrhpptC71G
PI1vnJp7kbcDRa/B/FiJKqN3o8ipBk+t8x/rxDc0BLpJ3IPJmlMHZ13Xqz+2MsHf
yrrKnvBVEgnQ5eB12tLupqzbDQOPVbnsXVvkv8Tc75ejhlttMtuV2PrkoNlDfjAa
zUTlucaYai+ArUoqAU/sB7UH7eVQd5Jyd7UD2JUoDMnjw/6H0EIqVCv2EHGRZwA+
2LI2JeNpYMKpt7ygxZYgDKFLmgL0Z8nRSiTJ5D/mRQRqSxXhLKVaJmNuvlDzqkoz
agdwXGmBGCsX8ZyQRJ2Fk0hR521tpl7MpWOIGrAprtZPfRcOyRTZgcqwg50YpK+e
C8GVHNlEQ0XLZOtv/90W6ArzX0O1VG6IL0Y/9Dnp6VwJHHYEd+nQXykWpoozukSH
diD+Kao082q0rS7aFL6488jmu6UdJ3RZ6MzDSpV1Vr7FFBQ9qLutrmzDsoSUeO7C
JntaILEVYX0STF2Gl92Ndbqg5biyslsze9nLpwzE1W8dOBCfz2uhfAnRbNVfeKsj
Nx7/4EcS5sLRsVwW0lEB7sY+6dbT1FiHmyfpfFrO7drMyJkC/bkCPlpveQ83lbk8
hprMaB6Vg04OFl7xNfpb4Ut840Un+gTuzg50QUypSW5hFsYF9MNqyDJyHCuuQdgv
5GaePb/Mgd90HlZK96VSdFYJxb4nXWatGWNNRX1QrcCWVwyBZeQroaHjDds9uryD
iwm0Gmqn6tRPi0odPtyuK6zu9aXREfQvyCFqJAOl8vDpGHFM6opzaUCCJqXVJrbX
wZ/nANXAuaoATfUPztqfI1fLWEUY0XNM4e3ST8BloWiOLIKPGEyyh+M8IKSvUl3g
siUzlWszAWswxrhoF0a+UhKlGtYGIrwlBs3TRDyd5TZfSS9Vf35hS1ZLNcxvrFWN
xvvKeeJWVms832nCnSvQ/+Ku/VmXNYMwKmnNf+d+6zXbx291V7zLjMMS4sAd8+TB
oKC2TiOlkFpGhntWp1QZdhZLeX6aBS3YlP9hUTsgcf4r8zudcoqN7Vl4Fi4l0PUH
owQ8RFEGWC8RjEBzjYfHQuq/zdMSHvXf4v1wHL6OzNdzI3eNQYy6uR693AKyVqbO
gCld2ccMz4Ew/PoJHFxsb4y8m4XPN+mJn0Lxelze1btZ/JqxY/EAJ0OqiE+Klo4I
QcsaUyeQrhZzRJPqsNSTqxv7cwKNMNuv9I53bVp4jUS/9iUB1CpbQdDi7ecvBvJ2
y17EQWbKbeUl8zgPE2E02dmD5EhxkFYzb7v76gkXFOVB+2UhqjOhe7OeeJCb8hYa
ZnTJf9fu5rQcLqLwVQ9fXt0+5IVwGeb60TTa6a47tCXLVdNu3WshLavgjM/WFi4h
UmaVmZIOy4k0U+otd/KVb4Nzggst5qHUpX/H2JylpWrlvB1B2pZrY6w/b9l6h4dN
4IXMgKxFm7K9nbL3WEWXI9IuYPBfmKMPdVFE0RvtvH6lBSsJqbwN60x4qAYEl4j3
ZFZJ1TPf7cuARBFCxj2T4yERrpJODkaitkuTkfrJTN1jazyKRcaFEtGPCUZn27w1
OD0I4MUGVh82PaQPcFSmt2VS9dxXgtBQD8YeNm1QCbVE5al6stOodN1mpl1DmtUx
YHfLhr/1+LPSYJsNbjnVUKDfOiukC/PaipcYyjiXnsEYkSade2D5WPKWYY4M4gZV
KCpWk8w1vyX0zSK0Asxro5BOm9UFppBQW4pJEkGqKXonbDMJvZ2Yd7KK19Bz6yDt
+76AD+IMx633XIE3+1Hoy3Dcq2O8xVKpeUteiTEPcOrfPJP55ACqXt4jbfp2c5zr
zl+vFBwzw8UwIMmoK3yMY/X0nakL6i69DIDTHfc5fcOD+beZHfRFrz+qz4Vyf/kS
qHJpVdmxPd8rq1ps3cPRgzPaO2xWA6EWX5uAZUpva1NjiZFMJ9o5XxHvvV62UPs6
TPPtmufwJFOoUX164cZMFziDRs+Dh1M/nnloaAU+tobVI36aTg6r1qZ6pSXqPWAY
oJXZu1WCtefpXFsXAIEBNTkv7dF4MuDNOy5mn188nmq3SmnV+sXaA71DlM4DzfNd
XJQK/04zY2s2Xe7giADpQmN7OuxmZVJ05OJ5WxNnEZGYCV9A0uNpOWlFU+EJbYti
W8pdTKRxcfjzqJIdTbb2yGQhb8t+cE4gMepsslAsvPH5Y5nTRjXlAkOB0rGuLKbg
fnQDAx6qcLeacMVqt7+hqQtC/OeIqssO2yNO3x+jTAhBEJG3E1lL3/FTsLRRaFoc
LaPqZfsUucSPGXlX43mtnQjUeArDCAHReOFXxiG8FoPQwgiW3a+aKXLdiaTA6lLf
rF/nEuyZxdG45Bkc//68HOL/C2ZRucL+qVFvxgkcirUOfA7UmndBeCzz9cBvpgqO
NgFnNefCOyC3eaOHV74EEwQsGV8nQRd2iK2roNFunwH/2X80W7H86skApWlMtB+4
xCdeJFjwlHU80n0g3t0EpV7z9g+B90bmwznRPpeb2CLDplNOky1eJ08DWSNnbZbM
wfOvZyN1fctNjWEr6EOXQDbsmSOu4OA2/lGKLhTLqDQosScozIIbOR2Wv4BJBLQl
ZAMNQOhz7GSk0I/RGLYY1bYTNviVM6hy1lp5glW0pF/aFI7CIhYe8ReZ8Degvwy1
aD76zNa5PIrA0DuhoZKIeBYQUETCQiGY1YxBvJxYeCJg2wzAvsPpzcjiyqEESKai
CUSqesdSWHQS3voghEcBRQKcmKfa68xvrQvGKNGQYofbv0Bg8NHW7J9chBGHrqpP
G903eQkORT5NIBxaxj/9ZEkdwUjrYR3n4uBZGC3p/uz1YQK2ORdzVgFhYlbbbUFG
Q1Daltnn0Cfh6WQOFAs6MPvgfY4fO+IEThCcwTy9qF8yU19Lyh5b8iQtHG0wUfNl
N0vI2MnsxKprYJYvxjq1gDVAGiNnwo6EndKDMsI/iK95X6yytShBKOCJbuCNyCZE
BVF78AJ4kPQVgTpVfbQspaObfNMy/LiJpGVUI9Rfw7Z+4YJRUORDB2QexwCqtl/E
yFEbZSYYtcun9FJANRh4iuQXN1ZPNwEFrAW1S3luE8dt7ltKg7EDfxNmHB4s7R9V
8nphh8iKXECFiTXvCd93FPwkwIvCEuFV9iqiQ5WNHTk3uS/ocMX3MvuuCgLQuwJ4
Vhbi8EwvZAA8TyRxLNWI/JSx2s91aT4y0x2bJ1w9X7ka/ATt2W32em+WCXg76uA+
PFWTB+f5ptZCTyBIKVciMiocfJ/H7UP4dwP6FlCQBdodJJrCkeQYXtGIe8uQWVky
Y4FextUZvjZu7VgTGNeVP2nNmTtink0WAC0LQl+Zfi991v/16Z8BuBE71r1cYRFu
LJ+9T28rdcpV3FqXw5zppnpTazFq8f/DYIOlf6hy95Ug9JJPPPo9I1Bi7fa5UZ9V
QLWyuhRzLfVtBMM9uErpWrvC61lLuyw53UaShnLM4FndNUCLxjehjPGXqSIuNFyP
r3DzIrGKWtaQQva0IihObWBA6ndFhWGCBrM+zjNQFF0b6XFZOiWJScu3mbku4ISv
lkTq/mifsQZl0IB1yc4Jg661tMpoyN56F0RGPgBxrvi6BQUefVlMIa3eB6tdZlBz
aiK4StNXR6DBPgnTLhbo6Fp4+vwyQpyASIH0FWQgYXKe3tKU7uFisFwq4GKXUwMJ
VB4ScbTbu9o2W0XB8UUVEOtLXmr9opdTjZWSKKRch+Rf2mQVpMfXUKiy2mdDTS8R
2Q6uvp/tJM8qQjoRhNhAtGpDeGvthJeMDN9erCSFgDxKHNUyK2SObIZgI+LDQN9N
bGqqjRARQdTFMd3r6Wd7xXuZok3L2E4ksRmj28Lg9cigfF3813LhDbqWaN/S8M2p
oh1+TPOVng+Mnz86pGL0vTguO8pMzV6xgO7bNopPnSO514F4keJtUOT4xkgtT83t
VbEvgFKYZgu/pb2zLagd29sK2LD28xTR+6eCPrio47UVrX9cLqDz0SBLKBnw1Ube
VN9AYE7UFzANjPWqLEbI2QfKxjp21aaAhwZHsuOY7dFlhefGdZ7HI+63ecL2jGfB
B8rosv05syNnyI/Ag8ZWSYwgFipEOf/txEw2mSe9MSuvd+WAqMqn9fzajMJx34YO
j3PbGivxpAseQ7JF0OpwPf45TIe0VyXoNeXuJ6SL5Wo9lgRCRO8EBKV8oScMYVBH
lKhSHAxGS9jKUOLx5DHZheWNWQ3Azwfa5o5hLmLABeHnpw2Sv1evCWapoCExeppx
c+VphRbRrMAWBFpuEIXjH41RG1c39HgD49XCoW4hsLt4In+2scSJxdn1oMN9XHGk
rWjUWTVpRNajZnnEhfYN328oRGjBtRWFufJXQgpttsxmse08bLZzDQO6FB/wSGsY
IxyYiUoKxoAiK59uWv5NWknriieeoilO9IvGIEQ0aROPwLr1MQ7vEJFPt6ijmynn
rkaNUFmOqLkhueCrabnUcWwe3FLiUgUf+JOe2EMOKg7KQLCox548wkncYIrqvo7a
NCzXV2FIVDabNSVl/hgHeJ0AHUjbrHv82oda7rXluOWmSex97VAOiLZGIrJRQett
HMSD4qBskZDTiNWlY5Ben2EpsSOWLyb2HMYrxNBFzkmuYpX2QfsIpuZbp9FWQDY8
3nadoV3JNFfIvnZGLNm+Tu50jmWnSNnTQYymScVk/k/0+FLVKSrIe5LCqepldyjp
ewcjeenACWD86z3pWAb2FdiI3QUeN2iGSPcT389R+z/n8puGT1U0nut8IAUQd5Zq
KlUTsG/sxSw+T7byr/55+d1g/fd5e+aHhH6hdUMa/vWK3aywfmHAd8s7qV/2qXc1
GOBRyTtrecfl/s8UwDB7GZgJCvS9p9OIH7lqNnLStHKRL6Dqte8gagIJbw3VNlvx
HnZxtlBDP3fdobG9x7lw69m8ekItoSK3lUspj9MkQK3UCmG3ZyGcfb8e2yWa2cr3
prU3OAF4EY0NEoQ+F/u7f/rNuo2M4FB8DAkmEmieRGxPfASq8J4kR3eE/aXIRFzC
Yi2CEup10aQAYeolcIlMU5Z8iG92RRTTtt4J0/SbYPZWOljduycSaa2IRlzIEZhZ
/58Aehk2DihRAzWLN6W+h1MOAzwwAtJh6HDyJCYpWKSSO864TYwqEpNyqELTuRID
wDMN7Q+8mz9hZUTM8znCbzRpwZQOMuIXSRk7OnanRCIcQbHnFoYoF/TOtVyM9o7z
hVDaA03+YzrypB7LqyXeannN7MTrMlznMXrG3Ap4/zabPDApTwYCk55FakwoYdmF
0CdRnd2S6nxL00rTf28axwiI3017/JHb5/cB0ekHHcAw4jzWlD9ilbpVuLizGIBf
k5MZP7LwpieQo6iEYftua9VsYv+8Ixbm/2b96mhpLtsg8j+tBKqn9wJ4nKh5WKPo
G6FKfnRLpTr4NHQpHpvi9hiICc91dMC45MJPox2lbYMx91ZtFdRdAlQEFzlJBRXp
GHSODrKvzMv1LSKaDGkhX/Yu/GbuxvOe8px0MrrmhwYi3gh2P6udVsT2Y2GbqFJZ
tCNWKp8XWuyof3xQjB5AbFUtLvJ2WnQIVWtpalwB+oBMF+5lgas9VOEn2/ZXDzxu
JfB9uKRCVhh8fh356bfxZbpGZDbJinkCRADrqqelzFYg4/87wi5IbWDzpBzbpJLw
/iDuTPjARY6K0l+PeDc7qFD77BdomziIr6ad+YKxf7R2v9d4WxACc8/sjxeWFbup
Y22IDgneJTFCpHnmtuP80h8AFSqdF2kKhYFAPu3wpyJqtt2/niriuWgoAZ1U8ZUA
7Cd7rhyaetdf5kcA+7XvYxaeVx9lup2NH40nCo0XkEt+NAobJVf8/QhtYOK2bJVO
Lgja9aiSh9tZGY5nvCXgsL8CQK/+DI71AgySonEhpx7WrQBwGRQ7e8mwOhY017bi
uaBGZo773aDVPFML88i2sKJYlBsvxW4hAbBGK+q1o1se/BmE0UqhTosV1v8HTsGq
c62eip34arm0loP0kHO02kgXAxMs97lbI89oQzYc8/kQsxxUvyIhbFlX4aVTQtde
qMrWJoRVJOnRXTY14yoEfXBCcYKN2LIdvRH8q+jDB/ye2MUfXyZ+M/bu86cjMOXk
hN0VJ+39+C+xt67Qtr7PNL48Yx4JiOuBMxIqM1Eg655DDImVSPVXr1ZelhwcnBh9
fZlpHA3OSUPj1psDgAb6TYW9LiBRm8/a9gmZCvgQw9nJnJnzoffeoa8CCF8LRL4p
hyEyI6BwotQi6Abs2w4RZRY4MPOSL/RCP7IL1+xf3wvbK6rYqLRMFzm69Be9AluI
uSIuNr2aPGCz8domHWVi4AKzTOpG9VD5n8Xhb5p1nvXGBUHZond4NEPNP7PakZSD
J8+k681LdvGanAxNwhhmmHz9De0C3bZqUzGYP1Mj1FLQQzlDx5QRUITP+JbcCOXS
zBisCZNWyJoSdOW4IfHGjMnVtw2039qMHKyfmI96JfwC/EBwE15Q227TIlNXzGHv
1Ya5iGKKnJgbyfckS03lg9+mmbmdTF2AWQbiTBY8p7C6GnWF30+cYxKZ27gReuZW
xdFiQ3WyrrAsDU1icidg3gootgJMqezk42KGo+oFkJghmkSu0GyhlvbB56q5uxZ3
uhr2ubBmQsIPJ/c+fRs/ufB0EBh0byYa7xyV/ebr7JJSRtBysOmtYZvZazfEq6GN
/3C3ubpnOklfTbHoztRB2/2UaH9cuQMBgoYBiZQFCCqmgyqH5TVida9MWEJZayaq
QCD93+19h6hwrwKrarlrK4qyKMCPSrD0AA6mnevDp4lyfOnR++XHbXzHioGHXieN
wsPrxzaWMFVIlKlpnM7ewTbTXUAM2/uzIdVQSOXmXqroesUyyN1C8fVX28NK+N3g
tXqoK52tlGKIEFvcjmlnT52FScr48uyaJGJXQ5VhCFUe1uUYPsScSDbH70OhgKj7
sykMlB+LYDm5dZVPy4LBqC5tVR7QFyXLW4TBW/BF5p27Ug1RSkmK4FDXuGxuA33V
V2pPqJWM4b9hiQTN4DU/95/TODZL3kAfHujTyftJw3QgZBFc+aBEdxlbQ4VlyemO
Y7BBuxfxZk/ibgodKOiONglrgysSiVFAO/pDkP+vc6OQs9IysOXf9v0skQmtPE8h
4gRuEgg/Ge51x8Izo2IEB0c5tkxetEpGjTU2iz9vQBSdWhefhY7lS8zh6G2c4Ira
HTx4hB5+y9mz6cNRDWHc1nEBgeyys9eq9b1DzJLXvwR8a+uXNuSdWR7aqaCLk/OD
trQkscEGAGonNNk29leJIKUmgFVxvJIfjkcECIzoDpZHWBR3flwEjzpWdAi3dM13
w03xW7zFPgxIlkpW4H4y0iqks1W/DUilBwpxY7CsQQlwZLJ85pvpf9hcUKzdRk+8
nKrU+gfro4lLFUfzgKQOfXO10A/sibCsvT/vR7kw7Pk8yTUygfo15sZ+oVCIrnjR
GLo598NZKDLSoY+hvA1QojCespNQMzRrtiI/JqFyy+rph3uJpaop/1p3f688+zwW
CYBdWDLAxX3tD/n+dzTZwceyRxzc1bj8iscCW3qCSpG8DDXOLbp2M/AHwjxDQO6C
DDbdED/JJy7M8mCUXsFYLTHXW1pWl0QHCZmOZJsB9kPb2D4juhQRQXDM+ClItIi2
MMzB1FS2taUM6cWJbFLWpzxeg6+0j95lk6ZTHTlbNQ4LVbXoWakmTBGFccjeQeZ8
PUTNZ7Df+fdMIbE8BSNeSa3S/Z2vt5mMt2KaYI+4EycA+4ZObwP9Tne8PBPGCz6D
VL7Yz5vxumiWedGV9sEICpg9ss/o6eNWG3MCabD8hgFkOMUGKVzkaudeLCMOPQWm
CE5qfABJQOcmOzo2XX94ptg5IXmgDQQtDfA3yfJIce4b+FwWzgfuIHKt4jhsVb07
ekrHHvOxg7GpgsgXuLeF/AUhrYU6ONw1Df+2lMKOEMp/elzlna1eUiDvBpgG7xHO
ZbYwU3/UxuaUyRtWl0NiR0xb10FUztUIKgs2z8E4HpI+K1AoWoioWPKeHpNjC50V
VV5O3oQ+7p6PjpMML244xfVd1dc50SYytzpC+29rq9q3rx6puYl8qSXj9fsfqBJE
ZkROWXmz1oLLWv+GQQv7RASUwZg/UfRRUqb144JtuvE4ukIatpl4V7PhZ6Kcr4iK
Cz1OJXsvXRkE03teHqa8fRy1tFOK7iTy5QmEPCbgvztAtSVDD658GT64BIRlX6uj
O8Ck/MeIy6551bzrHc806ZrAecS+5S4Bu2RFjgOOuiVNR/HZbwHlW7jH7VsGo/X1
tX36Sx922oYZqY+UZi2CeYNI1ChbEYmcLwjYT9bxGrsnp8G5QeOwdNdW4H98yzk5
vbgY57HzhkQSTrtv+5hULKDUDnuPkoIbQ77UeBZEC+3YEGzwv4F+XOQvrq/9rhJ3
9Z08gBamlyRL5J2tZ+TTwLuuZ/Qhg6uoyLAZRwu34fHspyOKQtN50L9e3orbJ53U
sPj0akCMnbC0PgDrrNEI3Sw2NWYiiU6w8QQa8MQON3X8q7vIBlLqAqD57QBxga8h
K7BY6TY6xUriAIpEdZKdOrO6Me+YQw4/Rs07nZPqwxRlXI7LM9LMoMZ7C+GTxE5i
OykxMJAUzurFjiai77e4zccxvCtWoUQZmpQ8vBT5ivkul6as6rxsANLJOb2FhoB/
kZNxMYgwqX9QKeykHBeAHY1ZZj5ZdigBEKHUIru3mAFUbhqmK5wC5Yh6G7kKzKVF
dI39UKo3qEEnoyI1CHattdxr/AsOU5zj/4rVxFJ4P48qqYzFHD0ANU2sm/YTQ1Zz
40rqXSEdR/3JmaK1j28kia0wNo/NU3gqz860J7UNLMLJAEWNn+nNAfJ4dfg/vYkM
I2d4i3L9QxJxDl7ykJTm8z/Grh5FXpdS8h4J9V/ZJjzmXnLaLSN8q+IW9jljYykd
3LdJVCW2E86RpZPFYwWrLnh3w9JdV28nXRU0IPvo+3PYtsIH3d0ZL6NY9zq0oNP1
JGYvTlkUW3GVZMLdNoP7VveuIH7HAnI/2Mlba2D5Gky4stJCW5Hw7zrTdM+oumXC
3FuF1ubHfsNS2yaLgSk8kz8kBEHFBQMoq/UDZb3Xy7X+2cwP9QtBN92qh9HcP89Y
eOvZBKK9SmRcAuMUaZs9MZOWflYyZ5OVD1nbJwk8wTEgOgZTqpdRg6bytY+OpDQh
rZs2zEwtsdnPW+Zu7hdOKOpVoLP+XtBXr9WQIzVuGIPQjAeL+xkNJ47ZzRML7u4P
juOTUKpaDCMFkb4HW/d74bP6spOwfZ+7EwVZlx/WDVi164IvQ9tTUvGdPCicNzI1
QVzJAO4XwDcr4o3hvXNx0yaLYu9ba/tuRjSkO7jjg7JL/tKzN8kRGNPASPTbtG5V
knB8whV/l2/hZ/UWb+Z7sBcAFGfBxO1FZHlkLWPhP82UEFYtXKhtox5P21tCjbSM
u6nnVh781Mpd+SE5ukK7VrZFBaIixYen5kKU6ebxZW5jTlGGRMdlPz1+ZA8CNfF9
Ex7U1O8PR8UakM3zR2/QzyzGDXNtzuHfoxgKbN9xYUFQ7CQ7lAbOEEl14yl2uXUE
AufSHzjGpBNsnTZq1jI0V0z1eZlat076Sg0o4pQKqutaDNoDbVYSUEE0wQR39ti0
I0HRhfdAMWCrFG2F7fxSwot7CE3QNE4/j6hJiRzILBTfvZnR+N/8L8bZwCy4eqlc
w1L4DXGyQBQbRY0+B1A58Fgex+8jHOAVXqkJY8ZKcPhpZnn3mVE0wMd9Lu0koXMx
LqS5zDS+N3oOQwvku0rmU081QNaW66vfjUkoObs35s0Xcz1uj2/M6ibAqOX/k0WU
kUALKAKkEzOfR2DIQSM36jY+uAYALAHwEbu9F17S3FpCQM3476R/Q2+LO9FfTJtw
+OLiTLFAHEVVsC5gFA8ciK08VRnPjTMJ/Nf2rl/DkmoBVOyKIfmaqNh7JDVYv/P+
ZWAzHKdtsUdiQeSY41wsdIWraS/JiGFOvvNJT0wqDX/6VdVpykqi/NX/ivWdgtZA
/OgqegRRcq3AvFgVbfitX1V/xTjeDKQKyQpbDLT34Y6ZBcRm7Xe1TVNMiauPcUYE
+zpRz6dMngTle/HAuIRUZVvXUNCMbFX7WdhxPCL8rCc7lG9bzFwk3Z3qzv5PeqMR
qnqXiVWPpH2PYJoWJYDmRJYp7l3R/kG3uX6JyNIdiOk+bRrP2xX2y0O7b/vUGszU
lLSqTaaamN2T1K8Lu7ktR5nL8D2R28NfrRr52j06148Wm8mcrcEjFSqS96OUEede
DET0psa5rQFDq1R6nxojzLOVsUIlg/5oWf5qj9oTnR0lSLZinYGqpngTvt44Nnq0
DyQNOx8cZWnoYmkIOjr92R601K2yoVDSG5pCtPV/47+BVw4HnqUy1RxRiRmew1o/
o5YLL3ESI3cQ+JtO1hXz4cpp/GBFBwLTFhf1NwbYfq8N94JIv+U3S5SPmvOfFeSu
PDhQpbS1PAwzsLg+yxPTmUHA2wz7hVEUeRKjxEPtVsFXSK/9dLwc4MqfHDh2UbgW
SXLFeCaXqjNxFmoVEPNnFtLzv+IM5CdLatQKs82bFHCd1D0wr9rT3+SJyOGXnYjV
G3TOdIW3DetDxlJk51yAm2aLPeEnqy/JRXCbPtwmWmc+vQB9/oEWV8R6D8QAKFgB
yJ033esQMiDWRghoQY1w0Unp82ipuJPWpjbkSh8bpP4k+6C/E6iMYSiPDsN+Cc0+
XNx0S/p6bXZNWHBeBPgCdOOfE23VWB+YlXgOGLHZvCJMItajcdOEkFwbeE8V/bJ4
jG+JkxGAaZpBI9kAaNVpAe3TGvvfv2UsKjPFYIwgvn9C0lFpnXh9rnG1v+H3gKqT
dMNk392VTThydGCUFuZWdECaL08E4L5JlpZs7d3U6hbJfaDAlNNthuLO2tuv3gRC
FmSMPKudNbN1AL3UxwVNPeDqeG1TBCU9sljCNqmn0U4O/fooCwxicoAnMRVMCsIB
dYSNQnL7ZlWbl4yyUF/amwqQFHX067I7MADasQrPNukOco3iONMpe5DGeNWIN5zw
jXknjuRoK2G+jzJ+XZzjDiyR3CaRE9v9OfpL+yUwAQkd2H/geBbXyp9oT9TWj3sO
4koUaIRDi9jgZACYGoAqysnLfuIv36sXB9x44DPyRXJveJE66O8HrNhLXmZeeBUz
KiXqquZ3bYlM7ujs0fXVCBJpV2h0+YwWnc8X0MYkU2j3mtJRDL+UUE7bTdxtD8D/
l8wE5V2mOMZjTQKIZCK7gbany/kklwkwtZ04NVdeWBxHL7J39n7YNp38gdQmbMEk
Hxe2Sfs00uHPbJtAH4fojgCIk+LlQnxmQ58CDWGYzPOioMF6YwSLSGWQnK/HxT9Q
YsbT3uV2bl7xqGDZY3xZqnFIiorkLUunzKYmDRu8+nM8XEg8FXtakb53cyBojGg6
Dr9oLY9j8LWj022cLbK2fwvHlIz2wd62NEHbwizQpnoQRool6qWQWYBDqDXeArY4
NkXO+XIa9hcwT+nJQgQkjPcyLe4bvkXV0A+o1xAFCdUvbE2bEdhsibTtwhQkZDB7
HOdQPwgWOb+uX3VPN0HvemF/0j+c6unsNd05TAOi7gT0Xk/5NGgv2KR8vEaxxDy6
wtnxTGIb9ZdjQJ0HgHNo7lSx0Y0C/8NnbJrp3/sgvFpD4mHv9aR9fXSXyrjtqlWB
8uKczl9FLBL8hhq4jiYdBiwrRV2xO9F+mTHl5we4p1hbTVBiuHz6YQykGrQx3RM/
cSOmnsaUuTMoycVLGVO19fXuN8UBOu9bQSGzs0ozT0eg9Dtu1WoFA3B8VSFgpxxJ
DveT3j+Q+jDGvgsurWIVn9D/idG5Sd+iQffhvjqGhL6y1n9v582DACVJ7BRes5wC
Bk9Ttw1ATJ1K4bOwFsxz4jW8uM1hMWf6TMIWmKt1WAIuR2xv3+VUAd02Z86/txiO
JfZd8ncgfvtWacd0vDRCyRR5QVpNPrXeiXPc6WPL0jYIKqY+FKjesATRYrM/13aW
Ju4MfGKeYuPQZKoUPUr2F1tte8RdQtj6vtgLCAdZI8KeeZBeYUDhEsWwfmQurklh
JC48z8KAzXRnqdKEGa7062GROHUBy35Uu2ghWHPTbb2rZjKdoj9r+aivQ+DHKGCX
ti1W9exNKJek1W8+0MvAOHhIONGDbC7egGl+LY91Bpi/4tVSkNFtB73ki9asRZf/
5bezE7Kn7uuFIia4AyUVpJpAi+6cQWyM1noGh9NPRHzTjcvVKp54C6g1OkX5dHz1
Wtr5e7uQgTI60KkBZ55pefvZk8TCJTr0pEm3PZSEXTLOoPRJAcwmfpbZzxKP66/F
TD7p1mUWyYUdANEpE0JyKgwWqoEBF1fGoRoIfkm7D5RoY6fS3NbVms1wwlnr7nrd
TMvFGTxV32v8iDqfwDnRKEAmPhdGfINigKvJcxAUHNClSNI+GSfgEcIhq7bQrcB1
ZXxE0yDlz2yrAL4O5q5wP2vaQYYQEfDjdQfD3UVPnjsaWk5dN7lYna/dYPxVAStU
KvkhMIM3hn2eHoGC7qvPTC7WlqhUEJHd5rzE2cgVniFCS8FV0ZbPVOaWCSCKHcIK
vakRxA3FeaCnvkl1+qPLB6463VA8VY9HIj/j6xrVVe+9IzWaMeA7Q8691ze8uDyD
2skWkmJ6v1co++Z3zlGZhU4AvJirwF3O6Rfrnu5aYbMoGuiCgDdbKDDYFASUAX44
nJmdqpj7xq2XbRAOW5mT8EmleMwPNsEr7cAD0wtkyyDTjpqgLN27L4spZPhyuuNJ
7m2TrHPs48MzAFweDIFVtJ0uopXel+5fo8MqDsaF8rHRgQ1mlacSK80wORvXr1iY
jPTanlvqoRU0Qa2SD/KN+8YNdWTHmq/u8aQ3SoRNT4BVKXPW+EEPENst2+AtYgI/
kpbrhfrQ5StW1hRrrYKJJoSX5FaAoOxc3AaMF7uL0vS5rpQnlHUXKEuFPZ3b7YcA
BIm1qtOa7qC6Ogmy6U3IcJA5XrR++kekEsu2AwB5i5g+jOcz+gJ0fJpFyb06pZ9D
EWLbMqpnpJW1VL2ilQZydIaNlvR+SKrjPxlpkgvsYQz+Dpz4XrfyaSBuLEcNNYWq
wRbXUpuUXE8zWbF3fEv0v7yYMgZjZWrSxPAj2Nyv+0npjHScXjMMUp4XsSaZGyw0
osYAX7Y8SWjlYjJ+auqfZcLDqzCFZR2vUpjGsyxpVFx/4sUM2WzKCN1lQSZSerb2
DkYwq7GF99KgdcSn0NiPEJbRodLH+9gaJj6lnRjF8IHqGctAo3pYpAHFeVnRtrJe
OGEXlUBNMMa8oFOsIiGNVTsqOh1WK3rAwNmn2tlsGCzYehnUQAgp53KU34MaeOad
D3yYqo3vk5QPVXW7F39EztkWVwc6iiXotvpy4ICF2GXN5zMEZ0CotbdNZWbpd/Pf
jzefw35tn0eujgm1jYCYH+NuVTWVuAfU5nfNPIqsZexzKP3MXgOo5rKiGxWhFePt
rcG3StPBoHnZhh1gHXZco1/91DwbxSihf6+iSKvSfdJXYfs8Kaz47YlQih5FCVDW
IZYMEFNMqyuPJupw5EnxTbq8K1zMX1idKTnUzwPCIA98C8l4fS/8IiR23I6Z85b3
gMX0S3PCdGFVOaC3dPkQp70OOWA8tMqa+Gp25QuStx4xAdXAMN2ePMYaY5tqpbVm
aJ5ie6V5lDIIy9V3j0xpoWkH7/hg3csHGjWGWqWPxu+7KjxuqGpJjUMJCrLDCkJx
r5qoNHAce4yqyRvdQRzJ73zEbViG3L26fTVjRXCZmqSujfdX0nTe1FZ94Bi5rU+P
XMqfQ62sC+ycI3xYTKIHuBQjwjNKQC/PMK7gQ2ai9Kt/AVOzHc5czuROobNUeuIx
lavQuPImtYDGUIPyxBl1MdX+1l573FgX54LQ/xzQrDreopV24amp7DM7cpIlOtXg
FdxulOkpbGJ01kvFMIzxQ/3AqxOulxVVmHpKg1/kRZPB6wAIpKQGw6Wgaw3nbZby
hnwLAiigj3I4xP6aa7TC8Ul8ypXqYc8eBWp4GvNMXqIWCRFO8HcJBdZ2okrYfgj7
AGG8utlLmPRCzb4i6+cZck2478Y1uzaww+rEEF+3mBbE9gGv7AbcpPee1saecUQe
6w1cyMnlG4tV+ITF9+DgGQzctNyl12hhS/KlDn53XJnRGCPymFkgXRKFYP0eSeh/
NYRoiUQZ7d/SjfGUYp8xgYlRGdJFnW1wDNfD/mB3wnFcL6darAnSsEFFPpFE//ra
zELAeWPTgIXmW7JFRNP9V9r+0sEdNWbv/jbeNJljgQD7ihI8On0Va/hT5KHQWL4D
nv8LUkqIq/0hOE8Ui1lio+Y/dBCs/TzR4mi7ICM9YyGunMI6MnBQMZAVs242laUW
9xg550sYU0TjLk7m6FQLMZdD0TxPMm1c7UC00S3mnLScheNGCtNWcMO2lhO7Fmv/
qQOEyPcjyET1K9yRJa4q44p8BCbN4YPZvwKE3jiK3phnzAs7BL4tYcLp40uJUPG9
nmC2SbBBu/Ct7y0tCzOx/8Y6bCGIyFSBOvpDLVDvOoEsyNWK9tFE9kuNMicsncMl
PlbtGYodat0OUoRzXIu/FtfIp/jX48AeHfmhapZQWFoBTvQ/1dhjJYqK7ySoOquB
Oi+ASW0riAg5nxH1kl31EClvDuSpung+APKxaSV3EMvDo6rqb6uFqJINZGzW5AkY
2OS3HTZ2HN0uJ1iAw3DfQQ01m4aBP7+kwZfDJG6RjXsddZq4XVAkhmb5Osjsc3xI
e/A75gsudmxEkxvrSeENBo134wM96qAVC6GzEP7HT4pWBAKjX907c8STEilWvlbH
algh5EynsGint18YaCHY33SiOEHl3/rdnzgbDtkSbM7Egjr7fyp1u8Df6jx9LTer
OM9xmo/5J+H9f/BXryZQIc2myogtJ/41TGJoMLFUOpu1lsfPHfrZNjaRD+WQdekr
gMY01XhL2qaDQ5+S/DynFw7VokA7OeH2Fv1rBH3VkKmX9bzyJs48vjDGz3iCJTsV
xqG2Ax5o2RP7dkAzEyozreN3kecZ89EI+sWUQN5s2PvfBKbqYVVtSvEdQM4iwvxA
taLMoJNoItQwHyemVR0ytLWUVY6krmZZ0PjV5uhnnehq5SD+9R7AooScwIR0sual
1nyLVxu+g3p8XaSkw7VQ39S24tzcFsfL6UZZwXVaVVto+txxRbrHvaNBqi5oH2Zx
WhfvMryY6OT7Ja5QSaGUMbV0SWnseDdQDTH3j/t+M5xPicVcrDwqyb7JUXxWLhnA
41PhNSl+5jHubX+dF2uMZi/Xu0Q86X6SfNB34uDxBd1CUCA4WUcOY+veF75N8oHC
vc84O3Ti1YWL3ZpOP7cHkVVfAyPcAoFerd9KmolR64rnxhq+xYcxI3dw3rPJICPs
VOidJPfRsbW63cQwLTibAP8oNu4I88+2lhz2WsNJXwX3TuwPoY7LrCdnlB7dOOyE
4BnNpwntqCPYIb1DWZDXrrG/WcE0D1BVtyOVgKj4jKCUJ1SqeK2gut/CjRHnUcYl
wSgA3otnBiyxctZMHOgiam7r54nWTmI2VOlsmT/P8sxwZXpL9rmzdq8ktMqKC6tJ
c+oS0khl9Y4UxnW4lFeIPaGXNYSVrYiPnixQRKKaq1T7gulPlgHwC/Me1/A7bkj1
TYFIm7BXQowp7vQLuPz8Bgv7S02hDmz8F+9ipqdS50x1ZQMgScFUJiXWXCTqQJ1+
xcxTq4tTE/6/56AkiOlAYR9cLbd5cimkmhE6MtVdivj7EmnxKjS0Q9L7P/MDX9KP
caNxXCus/YPfzkR3iPlvESjHooS4YjAIyu6oruvFDaEp3o4JgHN0XsrysiLP7riu
pEom0mPYw4VDnxStDa1d2oBaN3iiuAJPhkrc/FN/igyvquIbwk+uwpxemhEXon2z
g8/6VeROArtrpM6qZPaIP2LL6Rp9W8DpeJA/D7SqQVWqJWAAkFuddGdV6IImotxx
PpAZgwJNgKMLLaP0TWKnM7flBEKjlOmRFNItqUelpFTU+nf+U6IoUpifx4ifC0OZ
s5QlbGc8wTpSbHd+Bqpgxww8RroRzKFXEIc8yp5T/jjBx7qxJglXxRFIOe63cbVx
bbS10Z/9ffjSqkoPT3AOOTTVepGTuAx5JOnd2xEbLqeuecHjdL9lMXZjaW54RCTM
wk9vS+i1eSaYRYP+6NipjwmBgnqHhPgk+UbNV1JjBmvsHuvcdWZ3oi9D1DHgB4rE
4ZWj5DxFOSjPbh1Fr4P/3RhqUFnyvRkry4AuU9/WaWmXSJpBbV5L1d/Qm5CrMmZ0
q7pZFoxYyKX+2PxsrBl8MAjlkes3F1MDzhgC58ZU9aKnnj3drhbTCVIV55ye7rD8
6kV81uu6lwD/pZO4YyjVW0CRU3whdLSkxEBahl4vIttw3vZ/g4LLiTIUjTIZ7hqp
zokj49LlOOGswjGjFqlgwrZrXinbGBt0ftqkV/385X/bfdJN/1kDWuYlj9jH4GOC
+42yhzFFCDSkVUWWBT7qrquUGRKBfo4XaVtX4m8EPaLrfxl8J/iVq3cBLtqgr3C1
j18gekdAlpCYD4rEaPAhJsEUrJFLrX3KTlbezDuBI13CliLTdhqhuFIVkvYpGoUg
ub8MpiWcnHdwIjKvo2K6ToGgyxl61Js/NhiiQMB+zGU6dVc5kfFsBtNmWtyxYmYb
rluOZNzDBIhYcRGkANCk7CgimTXLiSEWoXjoNl0nwzTa3Nka1esQEbr93Is4Ql53
GJ0n0LfEYuZndBaWlQbo5juTc8d66iv46zUje658mKfry2xtKpip2c6aXjQblZ9q
RDjgRkZSP4GU7VH2hSPKjoDmzzB0cMgrmVFkBjXlnpOEvF/f0WDw1eGa8ZcO3BgI
717DaM9qccOeJiWj9odWzgDSeWtn22WFdXKCnn8Xso28YLR4tnsacF1KNYHL72HW
jatPIFz4qpeZ/L4kvWHKpIOrO+69p7MrBrq/zPPx4+wL5vCRHfgS94eyCBEoYBHa
WeSu77wSaZc/zwNLSjI7vBwdzCGbmCHf5l6QmFEN96hUBEA1RtTeIPP5/B6YDHC1
NpD+CcBtQznQy2mUdcFPS22NzgtEBKeRH8HQEPtGvDOGCv/CSKbk0cRaQ8zB0kKZ
1jOPkXXh3afV/PBDB4X8Dy3i8lYmmuFRQUd11Z/JSD9R3DPe4VXux0u/qaiqxtWj
zegAhgcJdJQvL5UCUPrHjXVglfqjc8Zz5ue9uKI7h38B2FFjRaN9bMrCixs8Q6XB
kF80MA5sgWQwE+g2mbu/bfJmr7fiAQ+GldjFh1FZoYEXr0SUQ1SR36W5eFrktbfL
0GAdN4MaQBrF9C4ZWN1OO6dD/QY6MHjR9XW4gNKfb2U3PtTFfOcYDi5XjcjKz8qs
6S9d00FvV2gBkKJntk5vxOhco1u85FjMydLByrqd7ZarflgwX1t/I0ufr6prGeEa
Ed0etSRZ6gPBHIzlbeQVUEoSd9EseLeeGR5H4yPdyLUNee0nI/+YPKHtfF0724+k
m7lHi/D1d9akeOWLa2tuk+03cPdJhwYpCW4/w8gjEL6tV5G0Ky5tO+eJSY8/UKQc
HMinS/xuhQd6OBwRP5osPB4HWCWldHN7CUlMJtgnt/BXdPYxf5c/nqLHc6H3G7TZ
rAhDJISMjAFO1nmwgOabNrnqe8q1qzOyto8oFDXi8JyT4ClI/h+RjJw0yfUNZZWW
vAyAd9yMsTmp5rlPw2P6dMrcVJf3UXJDUG7MccZNtcaz+70RASFghvqAODBqxQ2I
xXwb/ssBkcd1rmhcvwy5hn3rYfjqMVWxsEQoyKALywEja/OtAWJyyJRjhrloCfcu
8alVjujdleGcF/IrXUtSszDMb1TZ7AmyixpHfYmRTmA5kDNoamuia5fgGpm0jLgd
qfSJ/Y9ghIJbxePk+xAnV297tOZzGFQDoZQjoNSvsazIvau/J6IwQWLRJx2gEqPv
ze2QxDP7BgZ8vM98mlnebe5bNKaose/cy7Kc1L3qRjJw87HPKwTUNTJRAt0vj8xk
1dQXpiN1P1DcxyrlO8DDoen9XrVeY2KxZIz8Ggxg0b1gjzpXaFr2jhR3FqX7YZWe
3IeYg9WhjD6eBOwEQ7sYKvfsaLXvsxdnUT9FAXRvoGMLI8uumSzsnVSQEtuxvdaz
Eyn3NqFdOuc9ff6qAbk0nHim79oS2BpGWy3+kYOODKuXvGqy3uPjrKGUvIhT+cPs
9ob8wZGKXLw+QzsFw+HW7AQIGet2BorYo1ytde3LS/8qwOpsKNQOOKM02yqVk+WK
ApSYR8ENbbNylqqCjKBUxTELMRviFAQn/5AHXrqVXLT1+aW5o4gbG5OglPl+QTdE
gTJFoBnL6HVxDtQ78TYR0CWwoQhfFZlWKweq1zp3TI0xJ1DSjnVCDZeP+P2aOSbt
84deiR/egMbzjEbkaUBLrwE5YXSmTCKfLqSw6hU42hRU+FUImpmf4GVx0dkwwa1S
/rV6x3SrA3U/HNUlQTtnPZA3whXE+t6YDRE6JGW5sBCLxyXlUGBkW1F3bSeyL9HZ
jMoaoeyTQQ84EAvCVXZX8SYpxAG4aOSDQAcWXpWIsDiAJSJXRHIAUjxGFnejeB4f
sUHSIuhudUKnsk4AdsTVqn0Jlv7jz0V7Gma3rYxGBRX8/TH/3CbBMSGHlNrkknjf
Ihxseu1Ay7AxOroo4WueblVq2jzDPZhb9JuvM9w2HIGwLOLojwHozWXBnfVPunZr
5O/S33WGK+WhyqhWCd1sI/qGt6Ij1hrb8g7C23/uf1r8zl8XVs3HO1RHXzrd2fFg
+/xpyuuCCVrzWMaZpz/oVpg0r1wUvxLGZnrrHsvrI/MYG+rq/xGtnC7OdppdPGeZ
oEOjit/Inbkg579KgVBXxZer7Qm13wKIMNugorcOjbiSM/iY0f8E6swtJTforJRW
G7JF5VrNjoI3joL0JlXq3rMIat44v82nidcA/drLejgktK8zxNPNXn7/gaXUbxOL
MpwHH205i2nAPkjBAKgylOe9XCt1JEODYWWZhei2P8rsVTEmd/lk5mPM9+suXJq4
jL+cIwvLdeFkhbSqjX6xZ7y6CqUWKgxIMd9kb3PjRRi6retIvU6RL+5fmQE1Ecej
xtdNOIgkQJ9Xmbnerp/ekIUbuf5EVawxM5ITmqn86ytqgD40Xkl4mvcGAiWsLP7Z
ieSEgGafG7019YCF3xjS999gogYTKu+sIF/6K1HyiG9TbCn3dStE6Z9bFCFbqABN
8XrZF4ClffWehafsHmorvucoy9ZNe09Df1N6K64VfS3PH6t/865mPnv+wX981QVw
R1EtJuDzGIaw5sKSP65EttJIJg47O7Z7DbuCrPe1YG5I+hunZAUt8Y4+rQjv9O4J
zxrdL2ME39mgtDV66DrHftGDAIxK9zDSggEtJ4Aup9sOgxdbpnrppDc/2G0BV+1U
FlmkSvEfX+9OPJoXR9Q14I/ahxRc9RVVBLrXiBSb3wlBcVDTUEUMt4oyesUgLEyA
MJny7UiIPaL8qWiNNOUSOr3WGFHTkkXhiuAJtJi6P88fLkN76Tw5hX5YFNGwC6SV
VRTvwQrRozYIeZGzyGTGtScRjqa5ay3GiwmZosgxfnGsH3i/sLopACCRJm6r8ubu
vmJe4qS/Ri19dGn2JN0cnTBZxh8DhdKE1XURFosGb28Pj+Wm4NCuGT3E0GBViqBV
ryGPb5hbjgSAPVBYmJGAZ+cj7hq4Wpgj91h7lazMftdPBBaER42s8G7ucYnKNJqg
SFfdP+Lc6Qa5lJ1DH1I09P7iAuPQpNr8zd1Qx+LZS8lhtUIR3Qhtmf8jSsSZBc5P
qSXECd7p25VWdlq/dSt6Rm7Vbz5pnCgbbRkpx0ltW/UqkmylZgZnCiVIy/dzF1uh
9xdQdBUZ//Ldoi1kNVk7VcJqTS7y6Cw5gcRCuiZkjOhg4Ym3bId17q+EFVCW54J8
xTMwlUnYwe5kajTqpBUCKzxZSX+8u3bYxU5iH6NGSxWD1MTuunKpVX+FBQS1o86E
Th1l0J00ud6f6k9D4P6xneJsULiBNC52ysvpNC+/xxZ5pSRibAlXOxQGZvAoAOtV
rHP0RuepmFHL3KXNP5UAFfuwb4ULFrKabvktzJFx9ybF2pXpOZGwtOzoFQd9VHQN
N23Q1ePiOSp2usSRPeakY9AGy7ATrAG1DDRm8DCO6muQzuRQcK6A+fSGvc17LuFA
/2nrOauPajkrJGK26N8+MFVEZA53I4hJLH2nxb3f+i5gSghlQjOXq/ag6vQZashs
sOBUjplsjnQYU52jwGU3XmWAR46aCr1hh6cBDqJuIJV1v9ZGtu3unFN4Y8M4z5gm
qwknDhcq0HwBwoGj0OcNrlFjzDXjRnLROdfC8Hdr3gHrKV3+0Q4duFrZuQEZ75Ni
Oj22Hmxhn+z/LA8fdgyUyaA1VJvamUikGGz93As2E7/vMQgroRfCJSFXO2xUoaij
b9s5+G0oHWANe7D2IfvajgUD5d2JeHk976M0I5X4OIw5SW/AoSWpGT3Gc53dAXX8
bxA5iymac6t4QKZhWcEKfl8fBBYUHAcChXn6kH9rBz3NacdwG2wtC+vgJU4BxdWC
r1fBFWPVUEqs0dTG2GEZPr9Wh2d/f91+kDtqGmgHlb4v6JK8j1YtMmb+5LTSil5v
zGwt+wQ11Y34/+OTmVMHYM/4XQ6lFVsgVL7HM/9v4fDh7zuLQ0fveNYdukZtHCVg
84OWz7WO1dJvldOl1rO4ItCR1DAkjxxqd6C1NvvJb01EHPlGf2ncFxBnH6AdS/JZ
rKugTHZdUdGLAwsNfdrXTrBiyGdMisDsL5b4Ha1+jYviXq3I4cq4JpedLD93XKlX
a1izLiP5v9pAiPApb6hP2dkjK5Xurb2rCLPalutxgGhN4cah4xtSb0y9IG53AfdN
/hh49TAI3RcgMsaw/k4oH34Fq7H+tHAoRbKI1wWVLSoKPZQDSfJM2YS08BxtlES0
sIfoWsu1/N2lo0Qfb6jydN5kfmxPa3VtNKeldGd+6JFSMzmkc67J+CXn9TEznevr
46hSTGdPr3ifgjoJdYWSRBl3FHxedeTdg3P7YmykHNZ5GTclQ1fSLlHTv3cBezZF
L3SkLr10H0Nl1vpuP0pdm7ZS34a0Trb3GmgevIccTtMbEyGCtoRIYaoDJn8sY/PS
MBoYjOT5+TAv6h9+jeaQsN2tvam0BdESLm+7MDLPztepCmqpvsR+QNWzWxl0ratB
4RzRTXJto0JMGHWnqgGahB/KFRpNDVRuGWZaMY9vCCYZNH6ItbncNT1ite8Tz0yB
x05aVve3r6cYfxqqFm24FzlK3iHUTV3DY5I7hqMzH2tIpBkTvnPhIKzLuXYYKkqN
i1pxp4jPKYvaFCr3yYKY2PccJtkRTwR5ozNw0tK9oxD16u90uoAmyexXuTC4vry/
3mqANe9DDbZHtifCsUCw/Ugxj1tPPzN+0Jy4GAnUn9YSOi1aDBKFIo1Vhj/EoC76
/LHi+Wc+xhWjJbBJLFT/XxPKlBDsQ8G/pSc1rDvj9iJc1PAk2atcdyIyTTMYYauh
BvauSPxolrbwD0teviOAyHwUV3Z8ciA2QiWGmc64sPcrFyDixYw5TW41TswYzjtw
4hEddTGGhwOzlXYo6TQ10z2wyrzRCJRjGDBo6SZtnD1xA7l36vPmaDMuqDue0kJY
tI54rGIlQAxeZAXW2hn+Yjrdd8t5L8E3cU89cRpeihHIBkv3jDOrHd9OJZXit0gr
zI09m3afcbAAoBLqdT8MnU2V6pMDm0/rggCoCmA0+JcaIdXY/8kDMoOuesFBEnNl
tPt9F4whv13/ZTo4zEAP4m81JGrmLEUV10mwQfVmeaU/c1YiYDzb78CzU2Z/7m/y
UHW+ehgKgoQ46FcOw0lx/qzr+KJ49pT8jebgiQ8ATHnZ6s6U3iGgRRjNQ3RWNF1L
azXWYrAqujMTsupuVry1reheZrA3+Xu1ZCK7uTowlcnwZoDqk+Gxe1Byb8eosdUy
pr7QXP4WFXMexUVs7DZ1P91EoHcjtcZzDJoGJM25i7lfY3ftyYsay4zZgApqCTuu
F2EDLrf9UG1fKeX4WT7NP4Ru3sLDUlGnbfAFs4iTYRbL89OiMX/Gv7qNFTY2bDvB
U56rQOqxOPPSzzKFlEutpzK+pZtAx/+sLKfGsfsxsuFWb9/lm+oRnZIkMwJowyQ0
iUJBkbnX81ZA8brAwIvIQRdm1ovH1xQ7RTxlRabdNb17FR9JcYLNzU3B5cqHooow
sR02UGMFe5WjDGoMs9a4YbPRT+a04Gyn5l+MrMiJ3P8REEyZfDNS2hMj5Tn/onvz
18xFEaY4KhI63sUevO/hP50HU9jbBYyPZ4KI+zAc+wq3M71GfAN/M4Y1k72MfP8Q
mSPb4p7V8E9MMY0HMJSnHnEldAH57yFhT7T+uQ3CQ0gMzrob0trlXa2K6x2B4EHx
otGuJDxL6Hk+KFLVQ5ACyWiCCC2kCbdDx79TPyQpug4sr0fK++EDBIhst31HvFbH
dg0jTz1y8VgiC5kY+thsNM6QQ55ORs2tYVCN/aL+tFPm5ZSIfT64b+G3H3H81x1u
DUCl0p1kANJKIt80224WRJQk1yLyGvB8ZnTnRwF2xeLmBQ1MCv7IOZwBVMVyt991
SMVYXlsFIk+9C445LpiYdbcSjWi7sT96B2008m3lj2L+iWPR35cH1KWW97YQIHYm
2h7mU3fFWdQveCXB/fMJHYU9+sI6CrDWP6LKyDXguJHYZEFC277CzQGdy/umFrT5
Wqv5tCt+l50toY1fp6fSJuuubHwtIht4CzRcZZLm7Wask6+RqzSu9tlhZk/YM26c
0r012AaK3ES5UpLt97IhygPOqnSdoZqPGuiBqOL+fg7EcJHV7hN9xvPB7w1dL/BX
vR8Se7W8iYPT5jaESO1sK8Mvfs6oapWl0svrGsAhXdenGQmviogW0RtFn2AVeUJD
BJ/pTCZqEWvJxUnd9FqN9yvfLEvLGTzGCv6W5Yy53SFHqVPvMoY2LDb+rFJTDJAl
X4bCIpl9yON28i4QacMZjH1oqxu/tbvVGvYKKyKOcCScbKIE1Bq6vmX6HDtLO3e2
AHndw6h6itFplGlJrF017IgBk7GUvlDMRYGSlo7BTU68jSvAJF2jPJig9ZCedGoe
BP80qczwIbLHpKBjhyNW60twS3hGO5bdZYaum1WlE9n3erbb+lUxzPy8xcOvQKTc
9lZNqvV6+HhfnZPkwObjpgBdr/ngCX0FXl3oGMb/TxopQKUzpJ6ZyOPJV0N5fGib
7gkOX2AlXnv3LTsWbDf0QgjjSE1Y8iaheSlUTN5mi+jtQIl8vPklWMTclM27l7KE
opm3p6hk6eL4OZ4TxUC5rp49TTDYbRVc3IFhqzKBtogO/jPsrFSSAU26vSFplpKk
3694ZdwOwmoLFZI6N+CAVBF1Ksc56ICpGWEm8SokQUSB8UkSQk9bHYGDKWheEv3A
4MUUVwt8OcImt0p6jaXkgzbcLMqTPbZURXqliQ7qu4pMaW6eWfFalddwLtyrwuG9
fEODtB2/nQKnQFGHnEOBkM4LmH/kIsPQeziYRTBYiloO6Rg3GOoJ4vKcLJLmrhnn
gRcBOPP5M8TcPuXMW8aRyhJkZYriFf05vfnxJ9oZqzQ3EB/yUYyRKPfI94hkOdO0
unkKl8LuabUCYM9+hyGNgOtEGN4sfvbNpy4HNJ2+Uu8MHtMbOEqPZKmzYR7gZDrt
arYSxb2Oc1LiVFlOv1unSm3M8vUCrBF0sXc+PlzD6lfrSo9pjTi/yPwTJzuujO6L
DmBlr2w2OhIETMjAnHuvhXIwl0qgcvuKYn+RqtT8Sc5FpsCIYto8vCmgkoomJyIQ
GFYBL5Xl0vTI8Eka/LfjdxG85/gBbiJYaQHmJp03RjfVVbyYX01GWb9QmK6HsXyR
LLiDJ8g590vDSUDeqmdn+0J/Tw+IQJ30F/P796qdzxX9pbQPV/vy1n5cQ7MERk6M
fCXOUv3O2/WQ2syGQAwgD+i/jvaasktrgzifQHtr9nigPVRcAtT5EOeZ70b5SGPX
SqZKOsfvyWrmvaV/PU/YgGdDmhdWbbaJxlJlZLWdPShevp+j9Ht6dvTMP9htfcgR
RX9RWG00YwBwFmIBAj4v0j36KvTUL7OXMb7BIY17dZjSd7LX2tlZmpC7unP1w1HP
+raDSN0E/9UzCCHibRtGKiLwC+4ecop7d2wn85OubVHRJyqDw5I7zxZwvTv1MmlM
3uGZJ5s3UG1o6CBWbM+YkjOiPDiFaOA01uyMiWego/dswio2SW1pLmUqQX6tu2LT
FTep8w60lenyQ8mkOD+Ur3zaGF5aGKA1Az8J/BmFcXLQ0D2o42iToMKcG0yP6mT/
XjKG2meUf5jBOhw8fGi0wizxvZ4j9iD+4uqAxmxjByTKrcEX43KY/jF6/NSDx9ra
fQCVkslvqU26z28RiQSd5TmErtnJWuMv7GtjNGs9DFFwxUtDVPyUrZO2IWPSr47E
rnF/zh0HQLdl/VBHYclUOQPImEpy+KTz2Zd1T9ehqeoYRDSglkPtBYW5v+tTpydM
UhaYYke1AM/i64vyL7cBmwFWnE1IGlSab6vUiM19IOc86gEPFjwp2TwW9TRfakAh
dwWKlrx195oxmIuZSX4u0r6vHhlkKMKzgdA2YY5ck0MT48VR5SPuylxKI3fywWBj
3rWjhaLX0OK/LOHkvSk89soKL9BamjRCvJ+fa3VeCS71B1TL3LJTuWF+c7EbeEuh
oaix1VzNFoJ336V3KE79zXmjodta5p/FP9/fWbCepglw43rpjEYmHDMpSdoxK1Ef
fdO9pppPrgdyr+o8vGkg13NxU0nydfDryRiRZXVJI0IIoW9ad9Qzv3gXphnpOmxp
jooAMRaABXTTJpAS6HXiNANHRc4vExUcnoj2/wCo5W947mjtS8RSQT2VF5ESQ3wJ
77KgbqZJ5M42oTYSQyM3rBILQRiaZCfOJFjg8He24PlkU1xQ0oVit3MusWgUU3yI
lOh5b80Ka4xMMmgHznOC0c9jNdLN4sJ5ezrYVSyCOk4A1W+ysOnSFcz9pRe0O1oV
2ejNrJslHMqM8UBewlgoZ4nO9vKS566yuZwg19c7hX4nnUlh30163LXg1b1SpD24
2tFGcAACMmZL/PhMXVlmXB//MyF1euV1RahTWAL6lUmmnrdOdiXzkvPqVfrGsdCf
VPY8Y8ihiZQtY87l6D7QSmqcVqzSL5YnooFxAbd0jbSduDsMhCBO4wckN5gLRCJi
h5mA/EzM/NiYsc4zoujwIWhIptfPBRz9v56z37hk9c78syjrvxcj5PcWLRmXmUMD
wbdn7KnME9gG+wQ8ipdZrzLLQpwoRGBj5evBNmYhvbg446EFz6ZjkvtN0ep/TGm2
4BzficAck0pt+zgCZCVFeRdgAEBhLrXi4bbRewCh3bxP8z5xrUQTU+PC5JPkz1p4
IFU5drFSyTRd2FzjvQF4mKRQXrUbAbllnI+9fDOQGJ6o86FaRs6+Kvn3CvmzmkPb
iRZ/jAbVARo8jcqetH21ISU8YxTVzTcTwhZiKHR3KUpEfdqeERUCAo8jWPmTRnhK
RXeNnVp5xJ6aOnCPuJLpbCdm8f8qNgWXyvPJP9GZwUZO2eMRSE/e2YLQkXS8FDze
th7qQf2OviBRurCKG/S7mcwwoF/famOgeSFy7f7WLxgvMJPq1LcVuH2Vr6JVJGyY
oWnwltQn9wWO5HKXAoJ8JxH4V1HG2lSAO0Z+nFWNe4Pby2XDPW26ZRvGMc6/uVFB
x1QOseVTqbsgBCvFcNQji05u2VbOe7l9tzd6zLZPEER676lmPLb8AqDkSG3uQdIK
NRPS+ofbFfkCTrFnR6W4CmPquJcaefDuLOdMp8SMb54jRKZ6tWjNz5jNLVUuWaOG
fOmkWnuDxwuRFokhPixcl3JggDJOUvJhrapmKIPFOc+vyE38LpnBN4aTqhO8YAHc
MdWEDomNSTDtXWsq0PAKHaM/AHjS9xrMkUjxhI+2Ywcht1dsCwTHqNQbM5b0PY4G
86HLDw5vlO5d7rw/cXwVNVrjVFj7BcRsn9K5YWcOqYSVcXZmdntdRiLBQZjcw1Ad
696BdWIf6jI1J/ARxSEC0ETo2x/09WFE9f24VIKW5Y8eqDoGeGuitIvtaUz9Ashz
jgN9BGENxxow3OJ6j2SLzLanbdQM+LqjDGkoBlUiFoeEZHpHG084a4CvjUHqdeSv
9lO2bPp69+95BW/hRjhdt9Lqpg04d9g/PpnhGPYyNgdwj4GwoO28cRRRek4ZmpaX
3vhkardpigJ2rCXRUm79NuijBqp2dIMEWdb4vjIiGqN4L0CVXhTgCgl0m6A2+19z
qZ0C6QKh+H16oF7MreErYKChQkmmxY8ca98s1dCI4fUq3k01kywNlUsWCSnVnLJX
D3roe5tccgh3HhtW+f/Cx+cYUzCmrYdPY3cFQ8B2CLxeDOgMYYLsJSbYqswNtqtB
ez+oH+jJuqyfXhF9ju2DWm9cQ1/MUC1wxfLPh/+UXJcn/mBReZBykHXw1CjRkF5g
W17oZoTJwJUHWWNnrDMca+hnId81mFU6Aet3QWSfpgwakFEHYh6Zligu4kV77OEK
apYQXp4g1GEhrlk6YQabRheEiArIfILSW93WAygQSPedHxCFiLkeVqOKlH37Z3Wy
/yrL8UDqiV3fN1L5A8NoCgI0SOdpLfPa8rFqK8oyIel/GNjDsVQbWUGAw4qfp5uC
t0tkFxAkP4EqxLGyEJ/sHH3AFsivul4j9lFkcCLZdrrg8sAAhYG+6m7G/oBvOniB
y+hGkVtusnh9aGb7GqgObwrALm9s6pVaMgVs9qDBhX7ro/JBcJ8ZJNORNEk+gIMd
lyCnga2o1JF9cAm04p2PaefloFXL/SLhFHAqdHDuyxjArxBLy0XZVBhTt3WXHtjh
l8RTrlpch/qaFAjBpSStojE5uop5Umg/r7oRvn2i0NQ4ogaUwmsN3Nc5ulCM0v9G
AByAaxajqvct3vdQG3OnLeiekRSc/PDKQ5U8wGuplhwS1TiExtMFTBOg5HwPgGp2
8kZhOELKJFuk5yzq5LFRQUYI8uwSZ7vEv80L+vSHCq8FyCZEvZALtzk5yk8NTQ7z
VF5S/Azg5PQ+Sk7AMimXX1An0DYrfFLDNDXocPVPdVLDFf1TlvKQrhayD7vriLcO
Thg1/b/u4dZeY9j4uffznicTOo472ZdED8cxTXfofKeAv3mzsXtTnvy4IpyVvkOY
C4VI7lfEmD7A3pEyOstELpBrgTJMpLi3I93jS7XFW1TySA2w6F8UXaarnezz6p2M
Dl9aPbosKMk9XWdKUVO3R+p2lkKq7RGAtd6LE9LMXK+uKYxXApTXIdrXD5b5nKqN
sCcxtjDpKF/4qSttW9WoU8Vu9Tr+YHXE0vKRsoW4SthGRPF7pft9CP80eFJuAR1n
aRcejQwOt4aUoJVPWGyty2B8GM4LTLCzGXTQwDZn/TGrd0bEMY65PDbY/XeJNWj2
VHMx3M66pAc/IJvFAj0XBjKU8JtrhCAcGGfFReqDmd2mM1YxMShAdZU0v4LRQzoY
qGbCX9Gy4E5GWCQMV9ATVIqD0Zq7ocqs7etr87AkVd0jTnCRbU2s6fMEZHQmX8T0
asP2z50URpQv54wAfolkFt9C05y540j1697R+G4xP+qYcVjSyW1nJ245PW95mVMU
6LxDkCuZd18uFWVUq3sd3iag4lCCiWhxYw0a1Axj5hFKsUG4yj9wLeengxhTD6+L
qSPCianewyuc3XKgs2cpZiDthYzdb3Lw3UlBs3Nuj1srCmvyXUvCRskjKc7o3zT7
4rbtU7qSJcsyXOd3f/AWU9+J8l7h6lE8i/PnL1EZMba2pEgsFIItw2+LEGqsjPhs
lZguH640ukS0rrzsfh/4mZCBmIJk3dJgR5mOUEc9waN1cTzhxPzBamXnNGwkTzrW
YKOoWxQKAyRUFmOcA4Vs5Qb5kBlg7G85O4CKixQWJg8gYxl6HsyGjdMTCdW1glB+
9bb674VS/tIJfU7KGMTkV2wwoAB/9zLxaOr+cSwyfrUtRTMHE7PK9MUVUKH5Czzr
iaAW/4MU6FEr8iI/8FRNCim/PdgbtgjttDXSLCDEkkeMm+2wkd6E6DOkXgxnE44u
k/8/xsghj7AOsRme/GT5arZFpB93z6rQrulo/sCo90hyBFD+ugG1BBVDMcOk6OeF
8NvrGNp/J92RLiyuBmL/lWoJ5Q2upN9/IIZudI1mrJOZkAUbkA9QcqHCDKjoQWR0
Jq3d169MQfiqcFI5NjIGATg9IG/uI6PSODMwu39J/pz7log2KlhYmDbQ4icexVut
8y4gwZq26rLwoYnFTVHXhLgeMcp9LrGHH3X2K6G3o5+2c10Uj6XPrzwxwpZwQI/t
qnAGcvfjdUxfF4ILi4vgMTI3JCy6KeXXTXwkt5JthhPOAEoFO9AidRnj4okVzoaq
XBIzhObCSbEXhAnGXPB5gVj8Clvq/GUC7SGuATTqRq+vuKZWKR8DVerZLCHdQyoK
LLHxNr546YZ9NK1Hep+dGxhH2pShNm7mgNuhX3MDFCJoXHhaWs/2YmYeeCNvAObH
CFjQkSkOAN3fIpCpC7AuTCi4uy737B7Id00csIWP4Aw1X6+N7e9Qt23UAKZ5vKHs
0dENgJMpDwHmJyokc/TXhC3YPSryIHo0snDIo87YrM55ZtZoWJ0J78BArBMGxFy4
xaIax0DgE0aMBwu74bTo77W9aC+duwrx5k/7BBlHFpQNwkhwXREHuUJD9BP2OLlk
Ir+6B77YrydZoziONheDu4lmSkNiw0LT1/9vcUh4PKK/rwDAlrvsdiqsGf4l7lpz
xmCigFcdZ5POSS5Ykjg9iTVBKutohAMbvChDzD1HBpsYFudWSYoa46SEEbGunOPe
cyhHP1MHU8nX2XOHiC43SqjMm0ujW/JjtZWJHnrAnYTFCJsSwyaOTAPiEWuooSJg
rdLyIAMGY299z/8zGQgE66pByMMsTM/h1P8zo2jpoyjXfBuCzNLjxLkMR9C81zIc
660Wc1AMqsYS+k96OOCJv2mKLzFhD3MjjRRN2eVITtV0A0rjGsT7UVMbF0OfZw5A
5wofQM8mZbEMszs1aCUaHpOqONDqnjUmULb8UuCa+cqhj338eEd3eQmzDMOQPS2G
JLK6HaUmL4NKWFFcyjMkiifhyoMOZbDZhkDPEbe2ZMz+j5plrusoV8WyOuGcbLtr
xhiZ69WyS4q9Ql0JGqZtq8rPUOM8NEtdAnZ9ya89yDhRAM25o/jUnMzZYa/t6wah
HkcgA6kcvKHQudpEOr0hUsiWyPsQMX8v/1ingKD1fJzz8VMIzYdzeT8nLLoOMUUT
Rb0PRCyhO3DDZ53mlVcCfRb7gCmhGc+CjqDK3QfWxre+/WA448gQ3uFYPwWTcyHX
XAqb6q0V/EhPUJvNxamDQzhQG6Fq93GybMkJaT6jz1/G+8iDJa76pTMXD9BeUVYN
N1BIKQMsFHWYxEnqqZyEJE2Qdu/aBqsBQawZQXPDASZ20Ro1peitSxQSis/qGu3P
LNJN/YqDsl39inAQkug8PibI/bQYnInFI+jjyappRPPjamiiUisGrSDF7PPcjQaw
CdZFdbDhVlDjeCs5Biz3Tr8IGiuFyIzj13pF4N65YR2ITWnvvQmfyUf4aeYIHnVk
LCNSxRS3OFoFH7ffhDmiK+AxsWjKVmVrSgfozN0OHPbI2qarTAd0wAhhQTvjgAhe
mtVYN09i04rprr3sT2rvilOZ8g/qntiPf3NbFL8vqF4iBCqubD2W7Y62iuj9C1l5
qokCa0tZOm7FV2qAH+tmbY+uxEftR4c3LWfanHkIigS/deMqLeTe1xFzUzTWZh65
YFLw4lLL0QCby8F6Qx6hvPHefiYiuhA2hh/GBfyWK2uH+TmDmb/wVore6wJdl13d
oqqkedz+50CmLxcVQUyYzVnSvACADAzN7lOKWI8QRqZfHsE48bz2yuGfunC0fpqM
U4KdOgN/CRKW+1DmiKEpaLMTR0YfGp6wdMZHyX5i1lPO11RdFV80gaZTGn+WsX4p
PJ6UezSBw4Pi6X+z+TajfyKvy8t9ebUSX4inFCjuYFR4mSGlapIdY77SkCz9Rswo
0VlHiEoFDbCzNYZ9STq5lUJEHxAKdDHLiRTzR2EMNDiaE8+Q24JXfExL65Y5y4Nx
+w0X/m+hSZmzYN/kZiYVWeVhhjAIuaRmr9GyWSCJaeeQQFKk5skjZhoyCgk/JJZv
HxERHXxJLICkKtfmvGdkOIZAAG+mU+LH0UmF9WdTCE3fKKLYIPk3Y3zGCQtI0pJa
lSki6I6kvntbREaUZoTi6JkB8PHK4piNY17X3rHYTxsVlzaWQqWpQYkpf6vhbVY+
XYP3KpiitB3i+942Zp5v8Uw0frWVGQY+WnY5Ia6DlO61MCyS79dqDNHowmWG/st0
InZN7oxvaeSVj3Ad0vrYyQ0/LrVGp6Da+GOHxK86mVFWpbc04+ZfM790Suc2nKKb
I3mk8FUuOhASBKm0DSNukLARBVCJSQsiwtQE3X7XJjyBS0JFwD2UMahhv8Tq9u5Y
SleGYp08AH1eQJW4homjYTz5Bm7pzg7nlNXm1QdElh58pWZG8anw1EsRM9t2Pvgf
vi+zI4H2UVd5gy7eMsfi9PuKD7hEUUUY15TUbHf3fMsViJvAKE0cLvVMChLLTIAM
/ysZ5KuLGRqW3AykF7xfxmWwngeuEIW8f+oqQFcPxtOgWmacI+GOZnV8GHr0kg+h
ghTz4yyYooa+aKZQlRwZRAB9fuAz/Ndnt84kTjIO7aYcqOWPJHOCQAhkYXleO96Z
q7n3UiVeMvWcOKq0z0ogqobXbptQ67gZkNq7/TV4hQPx0Dnaf78iglw3KIesQcvB
r1n5NEqDJtRYzibvwL5PXd0z/Y+Z+sl/u0sKZJZgjbsgXWmaekBpk91s+GvDABP6
FUeIR/cOLYQbcHpu8c3MZTUfmUhfh2hBsNqyfZjjNacGcC1GTlOFvk/vhgbgZDij
1n+bkkgPYKFAbb9ekFVUXwp4YRBOAA87OLTFCUPp1GyCaA2w7a1nFVL/Ca9zp55I
QsvMLExEjHIY45xDcXL4oqbW3StKjiaP3AiZleq8V8gElkiQwEvAUrvN7CqmV2/Y
SGbtRjOAvJtUYaVteFbJLgQEjmst6dCLBOkWgab3HV9VRwIBMqb0ImiJ7xMByR7c
bldwdvp8sdrx5qYrV6kVRayXeARkGRfpyGhQEcwzNDqeKoIt2NQaSaWo8CxtgeyB
Cql+0df4iyZgF5Gs4dyb/jsFZ/R7ZF65QhCzanyXSaymnqFEV6fTCn2k4+dWuHMG
BxH1ylkmqYMRvPQuGuckEZbqEn14GolPyC1g2+1ADiFIuX75nE+1eXZJaHhv8Arh
NHB3lz3kInCOGKpVc8vzKgG8JcPi6LbApkVYVJCVsAywuOb7HtXjV9dd1q0Curo5
wxSF8+3ebtyrvbghzD4xxr20+OYOFoUfwUA2ZAPOrs2QXiwuApBA0xwkTCbQnXnG
Dv+ixMFyHq9LcUE1A5r8DmaZE59i2ODYAnlZI+mMVEgCxhGMGq9eZ3/lx2/ptmGr
6u2/Z02MPOy6ahHA4Gl0iEYH067OBYtPCVQ+Nw86ITJ6WnLENls5rQFiKW9IkKEU
V+SQ1WghWkix8Ls/yFsupmRhFX1Jgm0ZA1HT9vJMnFXo8nr9eVFxabyq4kPiL8+x
RZ4wbIOhO+xf5tLOq+XyHsgLMjXNZd68W5KttkMu4Ez66NUR/09yF6uIG9zBk5mK
mS4ztp937UUyMkVjFJRoCw8acurXQd/AizkBA4E6sAVAjetJhcMWTumF2hPX0hvg
9l4yTfnEV3kRKvT1WZN+g7ZG4Z0h3LPlqCx4895kgYSGTGo5eYLYSNbGrGV2kzVU
FaMtxGGqBe+JSeDhkWxdObcl7qJABRsh3RxSpRMrr/XVu6d144AdHQxp/G90i/31
cJM+ixoW2wtWjtMit7sAR1AJ5MeAjno5gqcMXrWEZV7o6roiwMAbedUfiU4S3R51
2PlvPkOWI6sldJPZj1nVQF7GX2asiqAF/ZOye0bFh/6GG8C8eh+eTQ/EhOZb3XKL
HewYCpz1JBd2S+CwdGYDCBfIl7QVBS+hKHXRw66Y49HwBBHYWe7tcxWr3Fug41R4
xlmiXk9xTJDAYVwRb5Bwzmdrt6rNDil9dcncIPY9VVnpUvfBVdz6N6tY+4Keq00t
gKllVOzEYtIb+ryjoP8rQaWiR3ebMHEWurCzKiZP3C7rbXD+jb4auWwA6dvcgElN
oEPiwMK8KQZufHRKc2Ab1G2pETQFZC/DdVin5ITStnV3VPQEFP0p/pOKB5zWEhku
lcnsViOA+WrEJ7yKQd0JQvhVZTvz3sqAsqI5IVPZ8LVbFDKxUOc1oQ0rKWWvgdgm
ewHT+6CZHUJz+hyB8pdqaaOPx7i5IVlLRy61l4XOrpEMz7B5BnfX4gFVyJpjmO+Z
Lc2yCUQGJCW1MMg4WEJw2joxtHv2r1Yyu7WNcWgKbl+L1TOWaXCrE2VyX9jluTYq
90Is4DjhsFeiM7g3oVQK00UVGpAiHcnT3e6MNuXHaJsO3pbg6UoKs9IbfxG4mX/9
EhopUMYmuPZYcIyqkuvYVeGpR0o8O7Oo/AojG6uXqWrureHdsn/jdidgGHX+vEdU
3zavvrFtFr9/4Sl9DYsHb0hXw413SHUmwn2d1ma9uRO4BrYxSqZaFnSYHUH7OKLv
xjHovLydu6kfF/q02Om26+/CJz1AJJfO8B6HAdeFi5KjF5ywDjgYw8ZIcYE0Zw6Y
r0ribnIn/9GA/Ke7fKzu/yaz+l8bFqNLHOGqRnQ65BsNtftI1CvzJRtFqjK3ZEth
cXGTt/wcsJuckjHVck7QSlY27kMhCKBYtExgMhdBT5KUemDoZeeuoH5SNqEhXf7b
lRESEVCCeb/2cSwE3ktYamR5lfHg40dER+3Cd19WEWB2Loo46CPld/Y8JTbuP815
2zBv2SEUhVAenKIaIbXoG8s65EA+JaYStatIYdcqoJ4dVKfucko3iFgDw6mwx9uX
X+MLUiDER4nWijRjIGLZekSfvQAM6pO332/Enmwl61VqNtFN15NXZwBnBojaRcA3
xycpdFUPBXRj+uzjKCKPrdMeWQgEgw7K7elbPopPkvb0GONP+ah0mp/BSw5adg53
gvqv9z73gnc0l2rfk9XZ31hJ1F5Mye3ynSsDbFtlutHQBGUrbfjfPQXplvtGac2x
MpGa41N+ntusF1x41J0nlLVPQ3copZLotYDua/sIGNxlfB85YIsFaWwJseMkxKwZ
slCq1/04miIHjtiPbiSf6Su+E1Rgs/oQBNUXJWjZw+xvCdH1HEnNXE8DGm2Nkjyt
4J0XGaQm8icI3u679BZCeHL+JTz2tnYDnTw8Q+PJDAJRgqQwNFJFUNZNQC+RlLAo
GCL3XptOGiJ+0NziGN5cP7jLgAyP5lxnZGvCXgHjJ89dFO1CBAgWpv4d2urVl6FN
srCueds58O4WtuD98bL1xQi24WJp8MmnB9eLXIiqSW5Zzb3Kbe69cOGhDZ0vQP05
FmJ0A+23GAb94hGnqzIT7W4kVVKiXSTXzgxjx9zNtQ+aa4Mti7RWGAkJ3nnyWPyG
csldFhADTEtdtJXteWZicp8G/cwPA5vNqCHiFsIxQkcR5IF3FJQ5KZ/fiyg360dL
Azn7gVlSZCSEQNlERdWGu+ZbB0oQ7sXoYrxg4w2tMDUqPu5MqHwSDz1rZxyQYdXR
DaVMUERCz8zbCDL2qMp2rp4JDfZhyMND84ODQxlQ4PQaY2t1np48vbpOSHuPSlR0
AufKVMu+7NaJaeXFpinWJuVlOpgLW4h02PwLs8t+srrTQJu/vT4FNO7mAOY8mOnx
7sgz913m/ZCru/W/F/F09SuYMYnPvP1D+aLuuOhhHUg3chdjxaZ5rxhX9T6HzJE1
0AycFgJJCbFb+SGrXEFuKU2mtWtAVAc4tGjr0sFAZFqNl8wgBXWGKAEQPfzcVZlL
WdiDHqcaX9y8BHwH0siJEBEitPDfy5UuqvJBRBTeRYa5ezngAbvGPnORmTkjSZ0/
RHys5fbvCuSk6Edi0HO1FnkRA6Uz2b2SjgULSrC7ny+funh5IUMnP7BE/tM7ho56
2sK+42JGeFe1jzDyQcm/77UxEV6r/sPqb53bXD+rIfcn1KK3B+UX5qbjgc/U/tgP
Cj5kI9NZ4COMzeKc+3HJKSNkFNI3ne4PY/AU0qHwr825GJRXyWxKTRkxNPesLGxB
9SPl6FkSrcbxP8+jpYxwcD0tpyBGMTUBc2eJNsNYCwRyCrJ72L7+KVQ2NE9NIQLW
cY5dI+jFxetyfM/nDcR72ZwwVRwhv9rbXZuv5mw46HxLOAxRHLTH7Qq8lT09JVyo
cnyuDOwJb6rY4cPkEqoDvHlP2Ew8DPG5LQ13b4UpFxVL37sG2QkV4O1Bo/+eIC+x
h4ZCvEwdjy140PR5nilZqUrRvT+hTQKSirB5M2UQ1wsxz5IWw7Y7a12uIVV6Sjcl
f9Iqg8T05q/vjk5bvecq+oqhYc8XHceD3oY7PIO/Ined3VLC9r0iIzLBWEMQOrVn
0Q8WQbyD/RgYLA71MkPkEcTJg2PohTcEpWSGmhSRwLX4LZISdu7SfOgcEGKzVnuP
6JnfQNrLiHVKQC5rKyYLNz/WLbi+p8U7J5rk8K477cRTwuIYMtM72RSfdRicvubJ
mY/CZypv+1cThvyrViJHn27dJSwTRf5Wb/npOy3j5m1oUzkKGwMjFdrMrr2aTwpE
3h+d2U1WR7G1vJwTQ9lKiJVF8XChuwDNfGeOZZm8a20g5n2UuoJ0k8P85i9ctLFH
AdN8WjXGOSctqBL5ObgW1IHJenJCPLKXeDvkVdVIrqM+DKZm6d50+LjgNo5ISbuE
fDQocwyySKtf5ltZe2qa2En6fQdqliTJKF74/NYN9i4c8OaDzUEMb3knw5mlvvju
NGbF4/EjdjMavBw3zovEaF891hLeqN0t8/usfh7kR/nIwuPic84ElIpvttr9sRfL
iPF0uPZuJn9Hmk9JT7ZuDnTR2TcP73v7FXzqsZlDZayWVkWV4kEzTfYOAJ09Sg4V
kau29bWfuFvSysl5MqlRlKO5hCCXKrFjU4MGbg3/DfuML13zwrq4yu0rj6Sn7maQ
rQDYjAWG87/BkNEhj4cxHS8BnPY1/XN/JE6tTbLuxi+OGBUSQTZQlHHybJYM/o9z
FFEOA6USdQrXHf1OcAfzZuTYCwvZFN1SVTDOW3B9G7Dmi+ekvq0SFdiwWJc1CiVw
eu4NJD69V2eUii44msk40apQBlGLYBmZ2X78Ho7H2ZYwtaiftEGy/qmNeCy/QVfk
ouH0Py/9LXCi7CqC9d7ztd1EM5/01yGJH749AtK2BMt7bzPJziyaM9AZyshL3QcB
XqgE7pYMk6VIR08R2KlNx2A7olsuiL+ldETB7ULEslkc7Ul/hYmCLDJ7WhgH/9xQ
CmMCamUEXu1lMsoCv8pFz1/7m6NlbfcBel9npONhpuiFU6pRGBo7mvCC7P0qg/tP
wjlGNyHBO8kmEe7je8SNNepfAn39TC6/O2qD7qrn1as8ZrlEdVoCNjrR3/kUyMsS
ZhrMDx67Rk9m2D1drFV6JSqGzMoI/CfMEblekt6RSYBv2Gx1ScDiMH7JdOx03wHp
IpoynXkssb2bfiARprrPpxMNnouZeBE9DXu69Pk0m+ngxl1mfNW10uamW8VaHkGG
7lb2ZIpKEH/NTQ9gLcavdSAb3ZCBl23RyFtJhOADj53PQS7k4MPt2S/DJjey0biT
QDZhnB9niEsIQe/w2PV20yMIsL7GCjHBh85A1KDmJwyQPq6LlgK5hk8/N2cBLMR6
lywkW9XdA2/UmonImoaVFk8s8Jcm7UkadeSLcRngfKQ29UK7Dj2jesrhqFwShCQo
6JMLmaxy9hJ9xahYN/FVOkkqtvcM36oZdxBqYPENUqqSr2ES4vYznbK8g2uPxazK
R44G8Ncf3+YWLH3m3Gqtho220HzE6EuO9bY+0PVUDVB92+IpetEKOCm+4wEEycvU
3p2UNJVYb4SRazU3O74pHDqSoPTqppwO672znJc4cChMC2MrDI42QzsyUykBY8/k
qY7kUURG7XRLZ4gai7+Ig5NjigI3P71i33Q+i6LczmE83/IbGrfgDGITbG0BKAtA
/cWpD29Ghw4mdNucxCVN00MULkomlrvOAVAzT7qOm2/gfOpo3LYdCMI+DnuKRXZh
FmPOcnok3cw2CIYSxgZG2LYvPhdkcoX3lWJULO3XnBINYiOBMHfL/vM43y7wypZZ
9cTG0s2DMjrEroPtX/g6Yft11GfLzIM93RcP6H4UNeElKUI/C9NArs4poJfwHhnV
E3dsSmRlxPcwpiSBX1V+lNpMpZ6K/toEHcMYnE5/loeLOrnROXxc+Uo228lJvmps
nbR05174n3vaj9T7pe+YgpWFfXGQRrUDlMA3ndyBcIDpf1Q+HK4zwsYJC0mUBCLQ
8chSLzbMutmtjbmTmXgDMh+eQHlof+ZXYPW2pazfwMHOnti2LqTIJ/MwnKmRzCr1
5ZyZP6F3H8zYUtgeom9Nw4VWLWMVTbY5BD33mzo7qLUg4E7/DmVg2kFPtcYSFoqo
vieU0+bG3bVVcYb9sdPZqOmdNwQFw2ParR2sQT2y22Ri05UXEhnSbXuwr50Mlko7
oCHONm2oxQzHwrcj86RpPFa06GVcdBOc5rCrQsOAIdGmdW5Xhla0hQ9A2rAvno6l
betUwzle6kM6iihNL90cLHEMqvONFTem8aFygK+ahXRSXds1mXRCFGEWUw6tHcw0
80FgINaiPSk6o0P2vvkSfFMgH4G7VNjr0t3eQYQ3b2EOCJhcmKpqGIjoI/Wve9yG
G2W13Ch/h1YuR7sbkS+rEMGwGShIG0msC0nLFiQuCvHxrFK/RtBfB8OoEz4J8jGF
2V5CrB42qAKU0cE6/D9VWJi1aZI5lkrdWRoR2uNYPJmVZjjCiG+n6Ug+iaVvpjsb
qKQhnsXMRTNnWU9DzNJ2shyU6hW6dZO5ep5Ee9nYDnAzXXIho/x4ZteVXk+nZsLI
uvlVEMXSY0dILyMypGmk5lqYL5VfkXqYEY1QAzZ5o7z63s8kBFHhS6DUEoc9jasZ
J0OxQhHz6kT8gxtl48XaYnQVaof4ctnUUTJ0d/BNhyUYdb1GLbexDysZcFrzI3rY
RLaiXgJzw8k//QrW8fzkK/b52jswEo1IQYLhFiwPUtjBMJpMKGM3VqhMOG+myYEu
kl68DmkbPfbIIH24FY66bd0b7Ovc2V07aPmD509mG1PgUpp+lzedLRZktXrxmD1N
2n6fz8ncRRVRDdFqz+4oVfCKrd9tnN3NXKc1Qwi9Bgl9a6S3+wU1JPnndpWeW0BA
RI9tWCwe/PvBPJkpbtlpmM3TOeFRv1Wee7YsP7aCK3xP9xiSfZAzdMfuTnAmsHc5
iTXQ0GrQJiP8PtOKRnlzb5+KObBS2y8pvsCGcvFKP2tVw8QS3of17yuXjFycM4Yd
Zk1ZWcYMb9Bgjyk6UYkL1CCX0FePgPqVXclS7p1rvzyv+LkrvFEXJ1HjGO1SNGdx
/x2pZkwWZm31/Yqh5ce5RpJ1+MZc7v0hNKJ+VfAN2Jxru/B1ND78C8H4yTvn5l0l
yCFjXOEWvEF6yQK8beMUbIy3DyFf5yjbTmCdtUWlSiN0DYqGycTn7jFfjNSkos8c
zcygFGtNjenfOhaojibLfjL8niootOYfE1f+UhvRaeBIxz1WO0LVDnyDhagVb0fv
P3zwk/X+7czMfS0OlaFPtLTTeXK2t02WX4sF2N7Pt8Kfgsts9LgvPuA0LJ6kSL6F
b9KLVMybhc/UZG75f2eaTUBkEnnDkrBI+DyEDtgRuSg69p9jAqBlFeRgziFpa2vS
LGje8HNv2ig/S5X1MGEeYTsJHmJXmnYBWa41A4Vx52fEmMJn6JjBTyqcKlHq5Pgq
zOEMifxEJ+Yedyq2xIo+CKpsazt+nv669q1PjBdo1O0u2F4kCE/RpJjF08z69jQ4
acmPgEZe8/REIj+imZ2yUmvKFxNflOlaZVvOStJxu3wdiKNY/VmGpsTTJKsF5Sxk
8//jA/nc7SFQdhHQFerJVcKEWsTW/AqgmlMsTiKPJC3pClSBLS3KN5j8v/Gca6T4
T5ulPijWORg7wGKhcwJwZO6eNG0PTYCs9I9DO1y0ircrG8E10nqK5paOXDSHj1G6
7KKwi46MWuUrnYQocRYwP022NjOpp2KqMpWNACoR8VP17RYZBkPxqD7/nRNz4wbH
+sd3fGWN/td3jeH82BRGt3ZNV6/O69EZKKudJexIs5aMsgJ9nAVQQv8Pl24Xh4GU
JwM3KhF1vu8+nsp/K8NFlZSSfxnUOHR2k1xUmAZwsjBCdhY4QEYfpoWL33SnVpax
X+P5I3qhW3zuhglPLED/64gt1qAE0F53qmVy++B5+DiTgHkt65XYlwYzRRGWC/g2
YV86d5/zCpCSaJRhzVw6/BaH33jpnIfoDtFI058gpl0qoDgKFG1PYhJ4YF3nfrAe
agw1MCd8dFh8q0JdE7wVuYML6vncJr6ty0sH51/4VrqlRqROstP8fauPKHO4S2HF
es53zo/xjBHNjTBPd81uyva6mejySuBsEngB+6uBzgIbAMDMwYuEREl8VIJ5KFPB
PAbywtFteUE1e+joMLoln/ue8POKyNawVrSC0PMWND0QSucULmbEgWmsECdn35AM
Gmt/hqIQ1QxegDX0yaus3jRRLg7rDz49nE7UZ+OcMstCI+Crrgwaas2KkXtUVStD
rFqJdkU402kyLduYNYTZj59PwvpK7FvoZ2SWrgkV748IRf6wmuPuA597ZscsRWHY
7oHjKE67ahOyP1WwJZD+SOqKnEB482OaY6qUndhr5NE299HMJlzuR2UWnL8yrl1/
11xtWzrq2T+gKzx/Gubr6QcCeUvG8OZ8SZQd7rMb+ecSCnYFwzvX9qD+c25Iy13A
bc5i/a/UUn8+/HP9n7Spoq+WRbY6cNLKElo47Dp5IRg41Gj6Q8SK4wwjZffc+Suw
bubOfe+sZz4zYdjBKWkL+Am1D1/hxzSoLwcQ6fv8QKDDpmhK4Ro/jWsP/0SEtAuN
BLnSB+IJoRMC1BKRo/TGgNR0dyfZahLjMOdsVS28rq5LVzOYGB1Up91gOOU6mc1D
wFyIuO7TU+HT8Y1T0j7JE7sunYP0N/jVtW8B/VaVaMs8CDOcOqrYTSXTWFT1EPV0
Vz5Rtm026ko7fCW90T8ARvpOwBrxU41wKq5xgzyrBJ723kTCReFhAwUtm6yd6G93
OdX/tiVKA5Bhj5q8ORJTyDM8GUHyFwwVXVxMGLjni1a1KfxwZkm9GakCiRdnQ3CF
ddB5hVClaLFGDeEqsGfHv0wk3ohDdpgoH91+fSu4ML6w+Vri9Ywd8GfCi62oqbMu
+vsRBUs69BJp9dY5XwUTN88DiNI0Wk2QZikvqDfHVl2TW3F+EGWuoIE8RzS2ivcs
0SVFbjwQZwzy3/ABPOIC35gl6aIqSSJyQdaQFQ4zFEXNx2ka7GE9grI/vgb/1/6Z
C7lnOdPta/i30HcubW5wfNMWXOP8xVzMpg0xNfrUSKH5nNUINLLefUnldjFgz3nm
0DGOUEIeT5gY9TRvVXuJ5/YybB4ImpdMaXg9YMbx37DyoP5N5md5VmwBrTVrMtTQ
mh6dEVO0KqyaGdevLwh+6HlCDa90BLKi6GOlMZw48clvayYbKpNyW7gXfWiNZD/5
uOnhg1VYZb/HirXWyuFRgiJ7S8O2J/p/tCvZ/fSJKQxE6tpkNZlaVFAx5Xy7yjCv
NalNX+a7qfbKHgo1uIPT/12vOcsooserVZ2yOrmQ2OWy3jp6km2KOSsQOwgTEPV+
QuDs7rzLgwhlemmvKxTAztM7d0LGyhJjXQQNmF5dzzATSlYGxmDqvi0wKuv59Xmx
630dGHB4Sms6gG8/62xadbWSpusf9YZF4wsmgXFTnA4QRRicXLPZnJf7ghxmdg7S
2w6NsktiVRIICL/9f/9emOLI/p1fC0ndH3kiaqON4ZhfDuCuelmE/tviSqAybzCX
Jt4tzZSQBAGAq34Pfntv/2p1oTMt7SbfK2hiCvaq4MHjJEr1Z8UbMc980A8JnS3y
tpEBRCZv/iSFtODkvP6YUKI2kur/1K64WzA0cYMgHW5ppKKuMgAK6NyKtUbu2fvf
5VFzAtpytj4q5BUtFIgchM3rmrDEZlFhxQJYaJbo96wvLSSPlaaTGiZwfm5Us5Uc
DRZ3C9HYYU8oMZ4TWAf7zfPo3BQb9dUAKLQZ4TYKTgyBnT4UpXaWuPiEmTXZMeJJ
/32Ttndqg2yYOo9r9YKFfoY77mCKvtJWw/TzSqnpwt55NADMmb/DsMTpfqDUjUtK
CKmncMhgzgZ08dV387dCZt0Q7vfPHhw4ERCQ4icMKDQb1K6DASY9i/lMfFiqvx5O
3WKORBhyso+P1mWmge5IHwGqNl5X6GT5ZiaCfHWAjgyYaoUGyKBGqgeGhJioJdis
OrrF7r1mdHe4J6HZGitwt5IeAsdfO8ck7S8r79plhsZgninp91ee0sEIYcrbQkHd
e+AJw1ypjgbnBF4cz3oejy5m+L7VmUUbnIeLZDJEC8Lxfy+u2WAZiOvlpsYqemHY
YSdEC4HizM5pBgysjJRLIPwt7cTyhKX1smQOVz75SUQIaGBWhV9l+yCl872SQ/JU
+mXN8Y3UoXN+JFhcXC2nL3qPsWhMggy/sEujiTv9zihrvrsRE85GoDvCJtNofSG3
MYpWwfaCp3Fp8IkVEOh2ST2NXCKJkrAANK/5BFCeq7xHea1mjNSZNC1nJR6oZEUz
t8J7dcSl2Sc+ZiSxS8FcwI5aWD0Cn0pZU47ajaRyvrSu6d0icDTWFKcweQ9XSxJw
K/E3OwptorMpO0r2RJJKZl4i/RKssv7otlprChw50xveFYOg1SPOH/om0a9b2uef
l39VDP14Iag3mOakQSw/fLealIoiYOIrY3WrM6x6PxFRN5+4D30oacsWFCHX1ayc
Wa2zBaBDxHBkrIH6gWA1mnfPkNJBom/f6nL7Jaw/5okyjoANLZTPdwfgqruCONEC
ObG1/fEdQdlIeCvHf+Jt7WnXcQIqe6w/QXnhfJ5SNrWliI74xMtwi7acTh42zNWS
1qMIbXxjA1l4LIMDVfraPSgbBj6Yu0tPR3kC5Dg662JAuMpgLtieousmj91rrDWF
T4C9PVCw3ulNvAnFlLpgQU9WjXzQUgJKzDKWfuXwqX0n99CxvtbSxeqvcs16xHgD
0ENAYQcl8M5Z0d3QYGSa5rETFfblt9L9/gAYeOTMqAgHbGSJWj+oq/5LZhqVmNRB
0Qc0nndge/xtu2eGPhqVSKDuqZsBu2X+YnYLN2sOPtwlds2cHR65aSdxjw3DDTWv
Tmger/vLAJfBTQ+YykeLK3vmskDp9Q/zDLp6xgPGqSkkAdwE9LF8IsgLKqA1NjrW
b+tx6LJbXk6fODpjgZA8Iecyd3BS4nfjRc198vNOZZfxpEPDZf5Obs/WBHBTytzL
51ln45Os/bFKNuCMBvddMc5C2T1bTv9H/B354yOEf56v7HEdcam0QULszZxF6qEA
PxzCl7fFd2hvB/oN1D9pcY6cMjod9Npa9Gas6kcnhaItiF5t/gMnHNhtX/Lzxbj/
jzyCqTTvSpB6/3XL8y6OWdIeuODDzdYefRB0ALj8usx3jkP5PvLSLHeGWBCzT2m+
tth0fg7v6sv6M0LapmqAZuSqt9ISkC12Yui1ALakoAqVnGhGyJyelqOks4J7cO1g
qFtShOgNZc3ek8BV13i06T6ATdjgmI2u4vUsQCVxvK31SsvgK8Rume7co128xs3Y
UPbDkc7qvQYlHKCP93SUgIWpMb8fVaVoaC+XRUySK3yjC/zxKpKueEp7pLq3rL11
Fw1CnFEsdoDpfEP8vs5fofXgER7Y/thCm5t+yFPGNqO87JUUIeCOyQV5453iEteh
Z9m09vfHKEd5M3OoP5MFHj9JhEWxwjjb2XxV8obVr8RsWOYbcHHbu/aL5pPjbNJQ
rL+7rXgpgSzD5HnMcPAHaOJPBQzreynU2Sz2aKLv2fmBzc5KZLAj2qK1ks3abZqX
sapqwMFmIyR2mPn/g2PYhgECIP648RC2qb2illpfvRP/aH/QrYfV0zv53c4aq8fE
mM8bwDb+UYBQNV26/WWxEPx9TfshkIY07fViJtugZAsnSvul5ix+gcBIQ51lSq55
ltfdbjaebyae5nCWzHxqGPD19UNUoxQz/s2QtCj/ttbc8zyDiRcTaLBLmVlgigHk
JeoGw6UGL8Q81FnDWZdmHLteTXXcPDBxTMr+GfwPy/sDRBxTIrUNbWdbwbHIaJoo
ztMheV3rMdT3emRD9TlL/1jCyM5V3smu4prdjwTPfP04nf1uFKneSMbI+Fd7hKSY
5vab1jlVS60BVWUuJ4nXXWRWlhr4CFlyTLO4d/SDCsr70r4JWKuyqah6Q/XhCi8K
Epr2mYS+1A3HIfg0d9pTYruHkP+63U3l/S8RgexoJDadBzI+cRTFHV8PcjUG63Jq
EcI4bvASvMZIlRlJ9py27rP2qdzJKkjrIxARCC7D8MnzLmQaYg+Rh5pxFe2JhP/4
5eg1T8Cf7Eb/ZGCv6VBTQ1yxp/1O/kCIzFbeQhYP61AAL9L4y+mN02QDkr38CMED
2BiUUHY2QpuGlBWM/zVzh+t2W23TEy9qFUP1rXVMRQ5eAqhb2EDW97ewjo0RASC6
N8KEuNYW1LXckLrqnqAFKx87bo/fGWycYVIo4C+/R4NrvLgsRGMEhpO+9I45XJPf
WnStx2hIaReeOXcl0tr51T2+DujUvCSDMMTA/4gNIm7hT1Lh88nPqHnYXOMg9tYD
JdefiN1CULNxlH5BdtPtqsc978/+2FJ3XUeS4p05QL/HnbEoZHyAkgzigbt2IY0E
tyx/n5DVtqHbvRpcl4vQo8LUEX5zn7YCVL4uPgQG9vEkbznphmQE4kkexNbrkKlJ
qgQW6H2OXJtI1ZjMwOjajKqt0nVuAANs5RqHVaYo3CLQO2o5kjZluyE0uiZbZ8t9
H6tH5ce/T093F4cJFFiSCkofpaZyf4FslkKVc5PfwAum6FiHcIqHOArTc6KaUsKs
ex5zncsMYHoudHMtOqnZ5BpGjGQEqQSoZMhDaYOxiZmnRxJe0HyKUg34eEusqzYY
tMETMVk/mpTb3dqQBYMTTcCtaI22KSPFDzU8WBpHlxKS1ZReGUmMnBdoduDroPuY
jxcW878f6SaSzvAppqLIk/ZSv7Qn5BDfWaAd8wp+1edHmpZXyVKra8Nc/iN1Uj8e
vY0GuH3otIhoWnSMCPUfYaftF+uN6Z8gctlgMrRBEp+fYL8O5a9l5svCkTeRNKGj
OwlYg2e6QSibCrE4cWxFF+ItqTseLCSSGDReM7TQUPlmGDp3UWVJhfs8ti5WRxa3
L8C4TjjuCD92zgEJmATxXynmPrZj2bBTKtLTqCbXoJ/6zWXYzXru7gy+A5uUtL/b
xZBISFpkWvhYWmVHCirEn0Me4E9U37qQ+s7GbAHFL3qacetDOgIyCrpEqYksaxwY
0bcXrukxnkqExYfyx7RQXPj22QlMVjA8K7xHpqESUFfdiIfT2QyCiqTjFthf7c2N
6quYJorV+Ti4U5RU1og4oEXZKQkorBDvtjiUdPQ3MrOS4JJWjyTarygWAlseO3c/
syePluODa5ALMRS7pSzoNc5v3+dUCfskm2gHDFWZAevXf/9EbojdrvBaS8fLd2X5
pjCFkybkHgSYfSlnf2eIfQkqwhnp08QW5goAsj4LF5hrJoxdZcLgg+0AyQ3oFrUj
xEePnIC0IqfIONVrHjs0lwCRam8XA/QUuOEUR8XObQ7wAQnyOWA94UJ8eEAyXdNM
81KPOrgtKDksfdK7a1u5nrqYfMazGKL15AhWszqjzgZvfPIJPTY+NIKuzKofE0sY
FWdOtCGAY1l8c4A8HvzZSdLWoelLG2NuLjWtQn09RanHWQcyoQiDv8k9GEyy5BAt
APOhBUvolvruDw1h/bE7oCVI00OF69bpZ8/EQcC68F9qZpcFnkymxaKormCfNAZn
xmvHXg05lWEzF4ifLKakuVIwh+SuObE3xVWqGIMS4a7xUIDAoAKufB6FotOi0At1
8/0jKM/1WuEuAAJPJC7kfhxtZA38m0tdHNfPUMlTQbGSn3asD6Auj+sOCjw09Fxh
oSu6p2ji0i57Its6V6G1L28LkyhzmPZysRlcXJDunDFIoWW/REm6yDw7D9xNxEN0
PTvvYFFKoAqfguKUaexVcyndJX9E0fAKdydsiRtugueagARxkjorSoiUvNa6m3wi
8zFhhh2S65NQbJoBA5+W99R/eTu5kXSXW9GaMUofMb/tFz3O1MYrA5hrLAuRz0Ws
eBZACgE8g2aLzpe2f8wCvoUp1JuQneLk5RxAIkACqF0wTm3NneRuXqiT602UnXpw
t4Ohc/W4M90D4hBvNf631YY0TImxogQJ6ZIEqypQeCZNKs1Z3t5Q2/NSMNaKFiMU
N31Vg6PhwFLrBd+QkZnXDd09HGQowH5Ua/3YJh3IILNqBT4RfPOKESF9dyQGUODm
y0V9+Ja/hb8pBxEgc+A8bHLqpSD9FwLSzA8GDrZRIqf6xhHC9cXztU+LEnrNRwwP
xqMPQ3hsbOdOcsVZyF3cifKEfgzD6U5F12y0+CiKjpjuBmhps43/tk1qzbSPSvoJ
P2d6TPDjkyk/hVMZth9JSmVVSiZ09r8U/+qVNbGD8D3FYkfqULaHs0R6XKRknTdt
g5MzI/AINB3dhh/Dfar9YJq4N8iMZWUSCPbO6zKe6Et+KHTjwEgeeV91G5a9QKR3
/Whi6xVaPhc37uCE+agaXo/yViOIfVYq33+Nc4ZwBIZKpyqQ4WUlySVLIx1NAQNk
kCbvt+9nDt5ouqgQHJxRa5diMZM2R+e0gQ/ThEusad+JXwpYVfT3ZlVzaM3SsJ5v
rhdgDNw+JunZUffWLR8GLTn2+1wSthidh7Ll3NwXWuHDCZFv7bQQ7I42lLqT+M3v
iN7MgORyHv2R+w1q3CUg5iu6Ek9LHvdSc15g1Yb4iU2701brA9x5gYZKqFErHgqg
mDZgW9ZmjNNNuYfbTu2XBGndwHq7+8LdjrSjgOnTfkBJcgOyg4Sl6pIOofRZCI5u
oVvFVVARoig3JG2NDyJi4E3ifApfceMhLSFrU1ZNss2jexbtY1/HNGGOo2HY9zK3
OEqc2m27aUlRzdZd/j9Wv7GZWtFJPjBm7E5oHSwJoHSojXbMkkkwdimCY78rUQsh
VnEKoQYOfaMRUA+zMoC6pMerGhzZNmF7G7lxjysrdUY7OxkqsKYNVGuNSE4WFj9G
/2RUYnaQ96P4k1qTiQzxb3+0eAdEdzBzir12Whne/QyzZa3IknzVST14uqYrlJKH
9sVFAwiFbFAjMOCwd+v1UWMnPIU6jTy4Kwtu4nvwdQfMj8qzh24/5gfVLiIEWEb2
PACQs2GcTqdvoK9LPxRMySQ00s7xtl0i62U+qgFQqhzlSfVDxOkcoq2clzooit2O
UGjDSndKI0us6rS5Re3hUyvaCCZu0ZlXWOM4SFQMyufrH/hmvUbRmTZGxlYXEvin
JH+l75KrpVGz227Q4ODWj+jpEZIjoL0b4AuzxjXxv9+xGID45UXaUMI7QItXdTuL
t25/KtJU1afc7F9dIfVAQvvaUxfNECXXhQO5+XJ/Xxlwz2x1bz9UXH0MjkD+jWZW
YwjeCXWUf+ipkXJ4tiQS4ShqL7ksJ+g/ZtFZpH7XrE70j0Fz+VBk+xkLfZ9yokRV
srRjO6R3aKAwCUjtkTRzg5qbEtrEWATw7G3bh8Qd488EfqKJY+KB9g2cG078U1gr
fEm1/1B9+zzo6To+NF4f9UwcLEiiywPYY066WIzCFI8k/6ajnB0kByezuBc3kPGM
8KKCmQu0XrtHr/+ochdTgHT9QFJ+ta/erdXQrUs/X1psn5EvHNU3Jx8bItgHDJbp
/5DVM3Z0t+N6I+IPOXNQ89R6z/IG5K6x5WM21q+0p4rwDEKe+Pdoosyt0zB7JJ7e
Uvjmy1v/NnG3lbEduo4aQcv27sJ0NQ8+Hu1b/CxlzLB4ABdBuJZhjV5TvDZ5EaBI
BrFTslHK8UOh/K1ALSWplEkn7UlvaiFE6nclwyvbXaG1dPvjSyE3ea23YlYjDsfQ
HV1pEnu5Py/5cJJbFI6VdrwAXjc6YE7p1OA/euE8p8EZ+Fz7G443cgmk6tQ2uBpF
AAAU54s4dhuNlDrW/rhzB6Xm9ib6CrJayvbwPYipImQe2iaSkAGHyfPH/vC7O723
DiHjzI0fLwYttbfRCdvzrvcGd6e3+5urnM7TK4s7kIJS+Bec9ffKSpSpb563Q0G0
GIStr6YhEL3Q2enOF51MnjMmoqzN8suCii/GMYDGjB3rvFkSXRobqFf+V2b/anGD
AxEGirLGWOgVGw83PVmCrL0qRMcuPABVNxRKC+EdimzZ+EXC41ZKv2yGt1wgYi5L
mLPSxzkInhsmPNWOS5dvmdyAVtfrQiDdGniRgAeWeQSmMXEa1v9d8R6LkNfMm2qn
/gPdW1K+fNx37CPDbk4G7lKD7FXi2U0ufTjWAlgwLpjhvAz7kv9xDr5Ivs1Ey6fZ
1wDQAKGibhfCwUyEiE/R3r9DjKi/7tMNEBWfz41vfLkKTsyvZbeaKYdDkOzW82nK
L5MdYMkhus0FTRoofM3meWJjfFjC0srEAntOXLonBEWQNccHZAd98HQaO++zqDoC
tc7wdUaDEXcanRdTF71otlQi3RopsYNFRb4fyS3F1V5MMEm6AcCwnHGXjsQ7wc4d
/9vyTim1ANtCzoMey2gDJWEEmKFfM93wM6H0L8DXQlV8CbvL7a07KJpPXeTsTFP1
pHGKjfwLUlAc9B6jA0sD8/u5RBMns7E9BpPF+v1dAsy3qNiJFVrTrAT3C5cXe/OA
Hh3f2pab5TjrErCOggAa2wZpzwB803kgtY4xf2E7OJTx4CZV8kesubpHRwUptpZS
ak8COnX5O+40O0ZSZplyu6UcqsviIezsSH+Fjo5lEdTydNOhyQ3H+vxNI9/aOzvf
nt2zxZYRmevcmdMix5sAgqtRBEGMnZXaCUMi+YDJHRj5EoNzhCHCYoiShvPNYFh6
TwBIL+Y7YBqte3Dr0BeTSfCKLmgs5ZQVpq+azYEfWgySqSpIsesC98aNmbS+G7Ia
0zjZwTe6bx0FPFO7w5qIFa64SYq0tkku8Ux0TWW8AK8lG7+nk6HOWwVWDLSmkKdw
P8NhVou2+eZBjdrM4zbvzpnkVChGmjfOLx2Wzv9BbQSvSt9FkVJeyLmY471XZ4aR
y7HCmioOK2FpS9QlIdNIPnRdYPYGOckyC2FnDuo0NauW3Uah0wzKYeEf47Iz6GMT
JPglKw/WL9sCEbzqt7aqpzQDcDy2W2hCvwbDR77Tl7VdVfk/P1lbftXsUNrRdwd4
myMZuN0a43/Dy7rg1JtVoV77wmfjTw5KFblJPCaFlx2jD02jrmqqiNmCTun+s7EM
8R+gOkXgy5A2iH7CDzT2+ooIEYBCERss0mvGVFWIsHlkkbHRCcf/Cdi45JuTsEDM
ARDTGb1OJ8wzFTnopb0GKwnX0tu5sxIjxDb1e6lwkTySIuWIT3IXbRHZTaIjxM0P
qig4Ddoa2FxDSmPdC9zGgv/cc027z3whhDwXVDIGt3+3rCjSOJFm54UqUOmqp3CI
0gLglcSAGyXm2Vbv8AysUGpJnnQRUmPPBYPvg8BNFBIDc+BHzy0BfUXqXOpM5dzW
CQa+wAfSBpmbX/djSFV4mh+zo/xxBAtetMbY4UvKSAYkvauAFwMLqAUc0AY4g2jl
yqlgMGa3b1sCVU5rSQjc/xSFRMgSq/1G+aqt2T87MXBTnsMGlw9jutD+TaLbU7ti
Syxf0bR8ZvcD+Uf3jkrJJvjkgp+guGm8V7bHbFrXovzeklaR4VOjcL8O0ANzc97i
ZQR0UVJZCliLQmuWZxjCx0s2NBrbPmciA06dDZ0wgYqXhECCi/d1YSN8/88Y8l7b
AYQuUIfAEWb4K0VnrIG4gDq9D7JS/8qUak4sBu6tleV6UREkt9rrxq3mmIqX/RIk
ys/M8wf8dUJ5wHBwxorC3PgDnsuNHEfYBEVdp2l85Nno+ZsbKNfDQF1l4HgIv20/
jg7j9L3BrbjwmdHEJPMeWgo5wlGAslpLGtLObKiuRO7kEwxkCe3dhZblDWUVrGJx
R2pL7rFblv572FZF/38rZSnY4wAXrV1DSTKyYCUhsiyjLIuHNxu68tKcebR1snOE
rWkLtoiGa+sHr32DBrxF+JhiH0z75IIAtNZqpw19O8vGssHADlQZULNw6po/9b0A
oCDhjL70xb4+bozVa4NTTpod2BojVhaonXwJEFZJ7xyf9kOCMF7IfjaixaLfOq+i
kQ7n8uI5O1zTmnwxtrP19wI19ZRB5sTs7yl51WQRoUoH3nHWAWmRdVQ+89Y3zT+b
EO+4HBuA5oxj35tQNXKYI30MkPQdeT+Lk0fbO+oXDbLE8lvtIaWCkR2hJESgMfFz
o3D1BP4CWEeOevd16R3Sb9XZd+Zj0nq/C6MBJtKPv8hYfkSnjKg0wNw/cwEJW1VB
9Xb5r0c/7qJVGFjC2mAg3uii7/xJiqhn/ZSgE2KClqhDkKZoUzPZb/vM7vcDfrGo
GKNHXICK2C7GaHVmAXubtJFZbDi3VC4S+7V3zC6HwhgXwm1i+FQcn+3UBo4zIKbR
5f/NEDOg1BVLZPrsZGQ4iU01c/rcGNNq+9xFFOr6g6lopPkadwH3i/pgV8JH6ZSc
nTlp7ZUs/iBzLA+bp0/muxw0mQJ7p7f/LE8ZdvmNagBSYITbVJScpUqWo/Uca8mX
zt096lgIrLVx5j6jT7ys6iyTDGV8aD+farFEWf3iHzRsC05PFipKSSir9EOGMB8k
E239rIrm62lWmUzQ7sn1j8xv5XG5V+YvYISt2P4iTALroqViObgwq/xb9ddXxUav
OmmA++e8uR0GR6AIRASHGqB3zRYi41iwZfvGWENgG0OoMSvPfjf0oCDbihg7GFSr
AjlnkItYOrMx9tY34QrCKJ/IoAvFmWatl00jDXmjLwas/F/Q3RA6ROLSgLDYCkcp
/2HLGAmK4bKSxTQIryuC9lHCfU3lkc+TCU8d71wnEfcNWktOfm1ItjkmNkk1HgpA
ozSlcwUm1p7DTcxmRs8521Dry2AZXV8qjhftW3pczCr5wkwJVfH+LRs7YTYhrfWp
CYRrMfapvqQVtiAmsaE/MSTee+FX+yhOn54yAnjSCURXMTEwU2OYsjKMzTtOgbGd
eDh6MqD6evIaCCplCEFoUGjW9kjF8qmBug3aixyzJEjU8RIc3FYNA0uxl8ygBLDK
bI5R/oofiD4oOjZDOht3tRhQ6QRv8fbYDmDQz0W0nyXNUVrg5HDB+f3jLXYhpHRF
ub+SrphqPOdZrg3jgTvadfZbAGF/NWIGRmd3bFtGXtv0m4IOmcyNKlHVPLkFLlVE
uzYX4BxITQxLb6waChvHJXcJ4mNX8e4p9LmxDuhB5sV4eKakb4w2IKSjABk6Mhc2
RZoXWneL30gz6ow+PTBKCfS97AfbJclnMhan6HnqN7ahvsAP0drMl6nSY02+A/PD
OpY0tqEqxTjsrVZrlYkY1bTIzn+H87Wf5aGsmKGXQ7y8g9DbVrb6gBbSXn1Yn0xD
extYHMceq6iBcgN8WJ7mv6HC/uB5WYT2LqIkaetjirJt5y1YtdpObGfmVf7axtaX
/4MSixPwjgD072wHopw+blymVTKMY8dS7YGnN5IrcP+FsN4aPTR4BrKnVeubqaXQ
jUENZORyapfZU9nwJAN5iEacO82tBne1/ArmPkDUs6zq39uFtvaB5oE19/Ic461D
RJT72+feYdWqmHPehLdKgSv/eXFAU+3v5vZT8b7NVMbIixkuUrkMDX+ewooKN6Gq
NpdevaEGOhmMFFXYKZB/ZGNUZfL/JcBNCPtYjFcHQufWd/CplqbPMlBAhW59g2/H
IgwzYszOjcQkjDKhPV6uv92Pf0NJfFzh+DINVabxoHSniNxPfD1wfXLDEquw4qs0
bThKZUKF4/6NTV/bnc9JUwjCGPDaacFBFAgjm2xM9y9WqyCxwSr+nAcbijyF/N5g
TJxEjrJjl0tNB/atAojFe2E/h1DbL6bC7QXCM8bTPikHCl73MXH50S8uIL0otiV9
Mm0DweHprQoK+qw1qg2BSvlUvaq//LHha5Jcqwtad0RdAMi9+E7FlColF3Wc5CyY
VPp1CvH4lMfG+6ixgENflY/zK1uT6AIKEJxzc47UDG7kVQGaC4Tc+AwX9zX0iKgH
Hemo62We3lpFTKhdu7zWSvYEF9jYifhkKYQGTKMKNNmRqR9SLflZPnyI+QaNXe6Q
TVMegBGmUPSAkXI/h1IhNiHQNo0AT5iw78d5ELFGaznMkfc7iVRdYdEggo8ALdFu
1Riat3Eszf9FII+hOFDNCtMJkV1HBjvw8rrEo5sdYXDHOT0Rhc83cnZUACO2gfM7
SYXXSWRB4pIjwS66w/OCTYeFxhX04isqnEX+CWa2ArKZpVj9escDGPPRo9kv916z
kP0aSkfVgqr+kQrOnnhnLwKMUCMimw1OpG+QsqHeBtzotRPodhw408Lrbi7g7Lhh
ewxs1M0BddlNWHtzOvi8XIXadz1gHybiRiKLa2uLV9dmSjezM0WTgHlhKTnJFAMG
ULEhHwSDA2Np2izUfIg5F2gEzT9R7gjCfDyp9rD0JRaSEILz3bHwBnyOvAu6Waxf
dM/EomTvvJ/9NgP8yN5n4t4F7pk+j13kg7AegHp947TnT8y+6Tic/F8arykWf0JS
WwBgGBL5lf9pAB1UrrZq7mpHmDYafgsaQ93MS9ov96XJ79whuFi56MCJQxTnq+sI
L73ENQLwYah2taxw3qlo4uliWoCvY6bUNN/YVAvpjvy3/7v1GDg3Ih45n9krLVWg
rVj3j4JIv6EFl16hU4HUPWWxu8+3YnQlytJ7VajzuagnJo/CuikLXKGkkG6GHJfX
rSShE/tJguvWBQBCdEPRTSKaLu0vsHf+yptXVq2pzXhbCJofJ4eFaYFP8ET0intD
+E61OA/aCkJ7d38T7npW/FjVeUlj+R1XBb5JG6BreOmvFTKpkb6vdjNF6AVu/AKm
DRl/ZK15KPXt5hv7Tk0CQHciM0H89aeO3aXdOK9635ck1RtjKk3qiV4/xdGL8VzX
2Bz91eEqxbCVHWnGyOJLcuedIEwbiEcmTLZ5tMyqiz3Sn97EGuzuf28s2pv4wSYi
Dm8VBG2PkXP1zXV7r3EM1k+gT2QIugZBMHYhOGeLwXKhU8abjx1/oPj2ihgJUc6P
aaG5/6LodkZPYFocBSsyklUY4MV0K8/kZTkzK0h0FEezThphiF6jeVW2mDXuQtQ8
bbHuchOhcDZ77utVLLNw3dx4E2nsUwUIoti1M84C6yFvBcqbVirI2NyWGSv0JzDv
Mm2SMZxGO8C4jLIqpk0TcUAVtVnlPVgZjc/XGd2DefTKyCuVB/rhhjiW7LC14/lx
/gflAZ83cKu+Xb064q9BPmX+FyDQk6jKrN29z2vC6Da4GJtV6e9w642pO1Fo3N6e
CHPyxx7USMOijkMnNqjryTXoYstSMrkVSLkHM/tSiJKuFYKfOaEZmQvwxrREBX6j
Sg6yhF3SDtbTOJqp7QxBV3+oOabUCmH8oFomAdA7E7iSMlKrPsr5GhSWjjt4kgz0
R+ZwvvYRXC3fl97ahhIpcW63G/FJ9KtUCHB4pl+YqqdqRgWzKAC2JzO3AVgQQvg3
a91YYv+Q9gsMqlg8TX1vnHdjSEKjpc5HGho2bBp0Y1YU/XtpfOg03z/q4WwvXnGE
Kt1hwA76RR+1gmAhx78aQ1CORSyn07rFuudbJIcdF57JMyr/Xg2aLbh4UodM+o1+
THs2Ao2IDPa7jT4mIIfZKmEC/0ynhFL21iQFbWFwIIT3PZ2CDPyqnpkRbZzD/Hhd
9iGLZrVBNuAWmvW1tZbUP1zSN9bc0VR6AkstsjdNw39n57btItYwKVq7bTLl/DH+
l6/W5x/xXMp5Poe9ubtQ/K3M8dAIewfetpFLjjrV5lDBL49QgjxrxROo5+96L4W2
6b5nEGGtKFbzL4ValdgI9Lvw/zKW5iu0bu10kOinHZFUh7v90VzzGq/EamfSdeoI
4ezeRvyQ1ECEYdJWJUhWRzWxIUylsTtkoOaofs9immKp5NZ3qOwp1RV/p5W5enzv
I7MqeR4/8gxLHn+hDvhzCWr1w0wSxF1UH0fWQb0lZXVOuJw57tKvi2uzdgA4TzP2
TWuzc7gbPZW3xQzOL7TBEWv/3iIVW3pmgDtbvR3wkRnQiHIuye1YpkOn9Rb3Ws8G
lP78zLAPHb1gqdzXqJGhSAPt8u4AuvsfauCB9fKSgxWT7Nw6Uz9sy7JtCpM4o8aR
JfX5Na27GDvPFFeeH7DF7X5E3I5EYydu2Hg/BDx0fFxZQghYuQpCFBcLqkse+WE8
paqPDNDQEqX6owiDgF/UDE7rAHMjVtgU8G/WVv790Se0MEZpA03EYO79Rg3HgqOK
WJ0j8pX5OMpBPp151irbZ9wbtyU6zdSk0Zk6PQEUKlB5FwPBu/A5BMAhx0g0IVW9
zt7SYkBaKZOXmiO998JootrY3NPA12/96br+++/Mye307Nt9Xl92+5uuyE7SiYYv
vfqc2GM1SnwLP403470ncpwXiQtOQsd7u5JeofzGiwwkHafoOGLt8Mg8JCXRVlCQ
OORrJ5OxaR3Y9lqfJgDYmWMdyDuVHeJ2ZVlp6Yif7q5EyTG5uhIcXdzjTb5W1Jiz
CIIF3LL2Fgbf0MGUrMFC5Z6/f/Qm7fOdgYURNGKnMD3/IL4xWynANeYJxmsBHv0J
a+T8AnFjXfR5Jh4SfBiY6C9DJOtMYf6+pybMFY2s0rwvq3w9H/1/B/L9SVOQ/4/+
8DQLB9LWmsWDxVZYt0Q+tLVsDV0AnWbwt39Q14d0GSiyGSSiV1n0NaYLtF0y/oUC
NLVpTn8o7cxrWHN9PO7/IbiLQ2ZKPUaTcQJo6xfoOInXjrAC701Uqi2rYF6ADskF
9+/S/fs17c0j5wDjZ64qH9RnuD4HZRNk0pHxbacB70UtDUjy8gNFF9pXO0dKrgR6
z7vgBAEMkCQE4L71S0oKmFmWV/DE/z+e0ZTWxU1xl3H/oW/3M4zTNVGCb9AiCbzj
sj1vzmkbamyOscEXF4G3TbGABfRLYg7cWTrjw91jKaz5NeTEIkyO2ZVPWxl4LjRN
S9rgN1waZrtzwec79qerLnblI0jRoxb7vGZRYvtM+aQIGG8kQmQG/VhL2dRdGBcP
nMXOXNBmllHiwsIXdPK2PGLzEf9FtS+EN/ZNFWNcSPs8fEH0F4J2qXMPuEhjFhI9
LlAbdoyiuOR/7Mw3wzKw1gLKfCXj1AgMnc5/0obzQa5F0/6Fwjm55XAaVy/9fTBS
E6d3B35yzJyFtqzYKij2kefroy/+JgAwmdJprtQTKOTOn1a3zVez95LYd//xWFAv
gdGekvnAc+Se5nFBfF1XUiNz7FzzKLIccBb5H875eRRCztKeXdLn3IHC97a7SSLV
NX6pIWL55+3jTBcfMFywyIO/EwHIKATw6zx7nEvskNuT749uIO9vpEwKtFCfhaZr
NWKLzfXiNuivq1ABAxzJUJJtAPeIDRv0dDzRVejoJ80V+l6nLQ4uDJA94oB/DC8P
ApCIpzcEcWSj28yrfoy7eCSNYNHiiU9B1XDmBV3QnUvBjYZ9qpDFn3FRfQzxGrKh
H/KLVkKGdi//DGDRzVFpbw4J1YSMjJsDTI4ZKy430W1fwD8ANviJqK4nRStl3tYn
wMWQaetsu7HcxA6WmLm9DBQyVf/GSPN3Ufx/QWpoTfaLFuVf+sIV8+P+HwPh/jVV
auFJ44gyfn9RybqU4K4IfGjLjVeO6wmwFYhoMZP5raa2ItPJyQC/wJaHlmnJTOkL
z5tksKZnoeOFY4lmk9fm0URebbGCzgCjHKi5xW4uyuU1NgnF2xV7UEEwBPj9YiIl
ciFyYxZSgk77oKvEkcMKWNCCCco7OsnDdIRW3qepaPb3lYI0H4Ords/Pd79yeU9z
vdOvY0HxMsg3NFsJNmtwLysvftwcKYC8PjNv6l4hD5/9fTKpqKsISamxv5nTqVkc
pKxaVTv4NAqabsN7xq/SdhsCQdepeI2RuVZ/2EFwNU6H8wE9qZWt/a95gXkcqb/O
zmkI5188tliidmtN6GcBJ9TG93XLho9eCQu4tDlxIutRs6Y0NOt2kruLFTZOSPBj
jmIs9mb6/4IOhgJ6Yitipi57HPoiXWOLTw2B7ug3ozAjbbf4maFTe/MPYRj361+K
U8TWM5g7O2cS3SkwRk9zEhToCjsbgCczoFQVEthFQClu0JIpIUkW/vR2f2QEgVQO
e261A1P+rbjJ1yhQBdnbKj2RP3KD8yRbw1Ez0+THvT0vvt9wVz3NkqLxBJDra0A9
SdeRS8c5aBEJDwejRj0Rgk3EiBFwetYIvuf/KlWaZ/4S8NR/q00X+KLfs27OLbpJ
M3dob30IW9fYyI/OOby3kUU1+ZV+QiAdarOumzquWHfJKe/Hn/wFmOebUWk9uJXE
lkD0VSOg+IjBnwzMWn4vvrwFycOeDNiiV0GRoFrp3HDKQ+R2O51fOhCFkn5Uvl/P
ZQvIrePbII1uBBaAeXD3Q7G1K5uhiYV+QmjHo5cbxbT/+U8MJ++gHtgVWwKOQ52S
XIBhnyX9v5ZCot0TnbiJ4XB1IgjO435aSxUOdfa3EBuE3pin71Fos1scNYLJO/Sr
uOFIiNxkd/GM90u4Jzdp7Q8l3J6XRWZ1dZV40uq2my0Iwl9vFyGz3QlIPawAQOzI
A2WtlAWhA773B6fUG+JAxcB8D3gXkbYoK8JndAQ/hdugsHDWgLS59eL/jy9/tfL8
rRjARf23pdAMqCTgLRiH8G6EVHY6bKQD1Mpo319EpCoyuxuUZb25z0e/JI41bmbj
Fajy+SxmSbc65NC00ALbZfdkFI9VfMwiRsfI3KE1HV9z2cx4oVn6u6F6VqSojpM4
fXTA2ZeRNIkLNJ0x+I7x4NPqWMDAYAlZYkaSKCxvIo5wBued7XcbF01expmR+AlV
6C0WzicKxVcGxc3qSfQM5F0zXaqJZ1yQ4Pli1N/518W4vo9/AvB3ChO5U9dspTGx
yIOC+uS0pvdl/xzGCMN/KFyp5t0eTRp7Iqk2d6WF/ldAbJ9Bqy0jXEuhPxAu+0H5
Ln4323r3Duiu+UvBt3/mJVhAKgYOpCCiE4aH+CRDovG1O3FVLQVAyCOlyAhapzwH
SWJHul4Maxplk44Y2KFRsfA7IX3uz6ZtrEDUW2gbiQSDJSDsutwdnE5/S8z99Sz5
7uP1UfXIQfwMyjziAMxjGiiwlItsV/aCMvnUIPnVhv0jwwiUf0RkardV6ktwhxYJ
M3WYF/pVOdHJ/9Syc5Do/5uDqt1sUFPTzLD3C1Qcl6d3TPn3sve+EiC0kX7M3a52
YN7Gvm0zRc/u2ZiobgzEKVfm1LhVxAnUyU/NMU+HNySwN4yOq8FTRVeIQSDtuEAj
Zc/IhcBFTkWJLSWlAHIDOI2vMu15CSHeorku9wGZNd9JADgosb8RB4XpdWUKo1LG
+/k8z1DGCBjR4Qdj/eBLDgLmLzdIhLdTddGYQ/1KVMgZ+W7GTYX39MmTEOUYRLCQ
BOKMHsahvC0P7tly4FU+1LHMI+XyxqKDi4ffiLo9PFNlJhuT2uiptZSpMFyDioHB
OnZoHl462zXt9fpJEtgZvPKznDAj6cQM5PQ9ziezMS7WawShYchTKFwZ2UQWXqxB
lfvcowjMs9UKly5nha18YW36/EYA97EfeE8Q3WybJhasudL0tC4j5cVtv2zeNF8I
gjFqhY0DXysGzO6bF1uRA875ZFNN57ztVpB6XWexVBh6Twi/Z7oB6GXaRXW2Iz1k
PHuob7lTUJAlPd/QIpPde2+UxAI5G4iPhbkoXOyvqrYeHBjHeozvgTDu0mgnAUA7
BkOECmC13NwEZbmzbdCPDqeUJHBWWqQD+sTogUYjfCfYqYhlfwgKlo60uW30+1UP
UZckl3LJc4wUrYXybmjRaYBlOWazyRGbvdzO0cEnJoANO3pqZKVpVwUfIHrMNbh/
OoHedQrVxRFAYdp4J3U0+q84mn7JfpRJ9tQCaE1D0lBnWF6YGc0bkIJsfZl3LDjN
qMfCswl1mXiMTzfEKGMZ8jNtjPW3uI8ST4cN8Wfqld1dQSliDaNOYEemqu5HdLne
dHY1UaY/T3KIxMRwNsPtpYhntggSdO+e76s9hfeABGB54HoRPOMuw3dpIZBSQakd
Rf6M+oWDwiuIWzXIZpUuF3yrS3blhVKYlySL3RRn9DqonJh6Whvte93avvJQZmUf
gSa0Nu1lHKQIfzfjK7hVDtSOCjlclXH+7hfcwrr6AZwhqCYlRCMFISdKnLXDv8yE
o7uvPqma55AaKODWJTRsZtfw7nLWbmnoNtu6xhKyMQEEsePq8cKQ/ixNoZwc6N6M
dvJYadSMSks9AkJ0cQ8YfqV51SD1YLkhNj2Nn3/KLyQPmpKyiGMPYuqeFaOaPStU
Mn0Hf4M88/pXhIbHip0BiMpRckjj5QRpILYDCLkRovaq9J3/tBtG9NVNalEw9dMx
1aZekRr4PGVRagkRGHkuPzr0oGus773LzsIm1UpTMdm89oTXkCB9Dq5go4Aqk5xf
Muw6O009/G6r+OXomFpGEiOXyDZchYkCC62CFiObX3HvUbbQrQdkSQGb1lc6dx4M
ZrIJDMuxjnxfJo77Qjm6aPlWPxoNqATC46JY/ArtEmHp7UIRENBMIp/uZoj4wIGm
UJsJ0yIl8wsfc75nHNzeijaeoX4oIqQ55PWaNMPJ3dwQ7iS1d1T5aRMF42a4tfJ+
Nysgj7o4urZP5Vy2ohxEb9/VJGPcl8xNsCQM3l99wdx4DIj9WgF7+hYN2A9U9lLl
lFlLOxFUyt3n0UfUl9h54VUWLC2DAhcEW7tXdo6dCltPbT7DNm/3DL2IafyINF1G
iYgwecU0g/qZbqpMrvhTnM1Vn3WnykA6NrK7kjuD8803Zz8gTJfzGDzEmESBHr/s
quADwriNy/qd0RMHLZYSEIRFQJXGkbNb0sekV9aVqtWt/1brQRlugCfizOKO85bT
hf8IXjZMc5VLF000aEY28fkZn3M/+3cZXSye3osCOzjr1C/5lYcXRVPwHdJl42oX
Gm66LGnMy0IcK6SIG5+QAKTfplvZsVnG8RRoCOte16Lisx/6kg0aGRevUtN5UHVx
vemtJpeeIdnxXvidzF8uA8kG1IXj9ZnwdHHUxtvgHIr1nATlagWIWvb3fB5SlttO
OfOZJuBXBDSErQFtzmFjH3MGMKO4sAf4beUqGjTHn0fGFShwrfUpOyuLRJJA6kex
RlolPmncK319ajfteFAa1PksYHKiTVlxu5pWboYd0IqyRNFsvtrCNnFED+qMhzyC
w2vCknre0b2xI2rGFq4/iO+akVAq+UAaoQt4AISQ2VlWFQllpbqDS5KfVRouz6h6
bm7KS3NA4dpslsDtiuFi0QJFQDMT5qTmYADTi/YxPivtYTaNFx4ByVIIqowRNAjO
Ju+mpe6IF4OPVY0lIAtEOVKDOVRjF3puI8V2BeTuDRsWhhmOvLMzsn6AW43MX0of
VFeniQRkDHT9MjpJJNXarnrpHfqKj5KZ2tvLZSRY+MCD5tY3wVNKZx2EZVK632hx
16nu/f/XfYNkJvOA8HftRo0XVp0suUhkW7jp3pD6Cb0znxfdSJQPj0zp0jpFrvwS
eS9ordVW0Urok/iuh1cH94CcgFLNJEt+DEvcqVH0o9Gw7XRIZbnn/WxPOSN/C8Oo
RuKv6PnURolJ2+a3daqZcFSr/CErcxFPzRNljv2tJt1eag7fviVu1UvWHTBpt1Qk
QseRRAsQQrK6hlHQeGDkNihuZy88vxNGCaiFEPL1G8sLsobtRHm5YqxwlucYEwaV
fIG8xqcFoTJdRWM3QRLLQeb8RrVzxi0194twiTGTe2W9rAGeO3Nf3/E1Ssi4jvcm
3KKb9R2FbmaK4279mqF08CVULr+DKEhbLNcUQm5nrSndNvgdy8mCVrKUmsaaPTha
O5yFjRdbJrraO+6m+eVg3CUju5S9Ic1D6m5qaO8mkqsI+mZzoY26nETCBvWH+Paa
K08xO9i2X1+pDfK087pEx88DGiy5XSc1Au8txX9T1GEAXESBNIHySVHjUxIN6W71
nSSLkRuuDXPuhPyo9Pob6Qxh2Z9BwmcGIU0fa2GEJfQenSfI+OGrQTThYZLqrTBw
9HlDE/mRwk8rFasrpGYB1F6yfHRWCflBK/S0EOeYe0pQKpMmb+W8jHlpi+51kXwZ
IGYS0yDXniItXKPKKQXNtSxunEjZwfDi0nmla/y6fIoB1dLNl/k7154OWdokgC1Y
LUu5OJ9Ky+7lR5VEZ6qv0HKHXHBIKjXDMnOSyoVNunlg23b2JdI1Q9775TP9wGMV
gQIgDlIxFjKxJYuovyUNoLZhYfKP1xsv0SegumEuh8Uob9e4bzPkhJteARs2NMIt
J5BIyaVgX+iOMQluHFHRDS2sBHnai9xxNlKslR+uC7Uty0tbMsAn5k1N5fAt5s8A
YKWd1MrugU0TZwO2Nb2rqifxrMnDUKX6Wu6RzoWqIChiKqmZ37nWmPeAT2elP/p+
azzl6JZIsbsPNAmfMFMrhFg8VP7e4K4NlFsOKG6ixr0lmbV+0W/8cV18QS9NJJot
LasmgI4HtWbzIsXth4o84y+B3RadGOClLIt/3mTDG65NidqOiHIyRoR50hI4RJj3
kkVVW3saAc3KoWbwXv0u2zTd5bZkM3/QyeZlyiPt6PQ41RDZF6uPoAwkkOuEIZc3
K8mTJkZozQpsTvsFlcAa1uWMIebzMVENAf9KoJY3EWQVCregnPLvlQpsVu6GgtXT
tZHZpKfedFrEyX7CX4b0wnQwcRlIH/lxzKSFsKTjMuMaPLz8M0r4sHcutMAqyCfJ
ELaBObKFoztayAzMwDL/3LadUAhyn+SF98Gdc0D7g2pv1SMlGbGcVkXc9wIv4Um0
DJw7KRw+IZSr+2WFbikuQY5KjRvzEz+0D0xka7HgSV24lRMuFPQVDnn+vGcZMOjZ
xtsCRnVTEKuYtSiwJyo8GQ69/MYIwxPcN7LWBghVPi63acZ/UonzuWv+fycq3GtH
VgHDmCi8L/usv3WMSv/P4EsT6/bSfroZFw+bUCaZAOtfvWiuHZGDOpWxaHihxx2A
r8OjWfI/o0+DDSKzH5WomLNJIGjBijn3Lg1zzWDDIIZcQQniz9CPB9A/uLZmNFng
bf+2DsW+hiSUZh9TwbJo9dtCfGagrqh3pTraSwh88M2QLg5J7Krsk8BexbgOU/q2
+k+uNlwfQ+PWeBgKhhliQqi8sIFZjA+fVgiCKBS4iOvhX6GA8c1ja4UY/BaW7BZ3
DHXK6p1aQB72lRvbGDjfld6PfbExTB64vqm1dODsX5ePpJuC5m79U1E5qW+EXqHq
lJNGBAZTQZQfg4yez7DrzB5yieVGSGQ/ZPu6MtZb5SBp5F3w7jCzk34TmU2+keP9
G/18Ey6+Sp4U5rxi5gJbyflQ5plwPL88BoRH0QObFoouVLcYpAYZ/XgHah4Pc0hf
ERXBme94X/N3N5SqfRReTiQlg0eRZhHY7BJqDf7pvpX9DVvIm0YK+xhnw1c7sBye
3QrznGIsSkyC/c7Ej2pVksiWNpWZ4NCvM6zUQKyM0MIG0oAQhn5I6RDoFOpUKQqH
Ufeg1+ciAyAZ2TCPUp3BOXXCH3e7nTIllok0bT2MpprPCqGEiHv6mBuUjnzdd4sl
+P3epLyNSW21DVbIMyagb3Gr/QiPBCWWPbjO+Zo98ejI5beAQGYrNja4+byI/02C
/DleetpcJm/ua+1cTr5Zu963PgJGcMgscWS4D3BDu55TbnZ03PHB+d9up263dhyl
V2DnEnkw5Rw6nBek+b5tfwNEqm0eiwmCV6L5x+8uEFkh+dlw3CmuB7J5+gjlqmmr
qz4ADdqfpd2IxxsXBNDKEsvj+9iZXYIy4s3uPSHSujdfDZCwjNiEh+ql7UYX5N2b
EeT+L1uP+xewjeaoyIXHdW4WEuqqSlbyIBoQzPdkftXG98FLIvA4/ZBpGQjX8lao
xiKEIjRSyTzUUauic3HVECNZu8uTnNRqRXPEqGqm9Wi0HKVnWBZdvSimIF7ONwu1
b399NcXs4YjteY5x3ofPGI/noK9uh7XvxP9/mN4Kp6pDbB9vrBx2XjI4iUS1dUNS
WEj3S2Vfh0+3naUL2oArcoN7MDsmNVnazr87k8lkFhWBpRf+v9/8y0O83Rk4DipU
VkTzheMQ/UDw6PdL0wjz7LqyWGVn3r3acpHiz7NR6VInyLJY7Te5nTBejm8Iix92
lLR63dc0oZVsmrBb4RTn5sqG82YZe0E+uOiFQQiGEVPybMH/k+GDy+hWYrDoj4GD
Gwj1A3BgRrNP0kMN2EXbpggeKFfigrvwUfW87wXdNL2RKXLb8mIXT3pkvNqj+s36
7fHSexYB7YKaUc0QuMU6OZVplyAhNOF2KTPvBYAuNbBRflC1Ut6ioxAmfzlmRhYX
g70P9eL//mIzj58pdxK7fUKME/rd0VUFFLoQ8LcAQ+TjAacRNbXRk3pP2EhjwBZY
OhByZSnqycIZeqlHj975A+C5DrA2ACoNHhAIWqms2n2WGAdFN/YdWWvjZsB6eais
7sdLXekw3M5SONWoH/Wm/sYJwOQJD9c/mCC78i49ksbKtEOe6guqR7ytW54+VoRG
QFQ5BsITpJlVAXP9a9zcA67j3rty34nRrYCG2owbwL1OA6pVPVSmsZ2rCNtJDFfO
87LTfm+nv7nNaQkQ/0+l28EruMRdYAAx6lAmaVm1P7xjUFpfDRY+2e6h4xZM2+HP
EunjNe84cm0b6YzUjSCaHA3aEMCOCGcFpXxK1jBK77x7E+47AZKvNiuNSFlTmTiS
SOSdXzueIQ40z15xzsXnDSJj1tGdcxFKmxZIaYjysFIYsiOaH971qeb6QncOOtf5
cA327hVvKsTqcauMbUhOiXoBTfG6axAQkLDkDfcT587RrymErXHNDETFO3EtHdDU
Lr7zdhsRwuG+416dTW5qclZ4WE+GYm45PdgpGs7p6Yy1dCdHXVU5Q4AQ+eGPGOyi
8VTKyqvtFr9HQofJUHphmQ0isZuoXTCiu7lb1lWKDjoLpgT8x6CisIjiCZ99SboE
1fwWZjvQDXUDvq/UWRL1ZQOOyC8n/dMIMkhZ1W1LL9MRDt5CfQtVuZXPGPkA7Jh5
NmcKdJTuhQMDcqxjoS2XS3WEwjPGLWtFvpW4QztGNZUjSsdJk5ukHHJ6DvlQCEKq
3bL0MG0rG+lKdUJxVIj5ZJD/zqtF/t9XTfKFvrGK0mTKT1eCIrXEWWfH7M+ycdy9
OuC8mbp8e+U9yrLRdYclT8pbnhSTLI99pBrJp4rSHzMbnXT+9SsvsNi9UP/ZTXal
R334pMGXCb2WQ8quqQkMyfirrEbkBq1J1EgmrAPV8C3Hea22Jk13T900H2NK4zH7
PnwgKEJAxtEaoRRqquO3JYQ5WJu8KnBotA9jbahaxo8/HbnJrGKPip8tijfY1NYN
F6KT2ZGUZ8lz2K8imw1k99ZRaWmXgXs4/goahOC+LHTs1Gg/R4dXr3DGDzZj61+V
wh4eeZpNuQovWyxvcEm6c60egpBw+iMcCXmlhys1u9Hyk3RFqfNwGVA0rKhVwUVw
fYTU3rzypaITSTdREICcHesucsTyXQVcrkKnFt93c1dbL3lVXzX7As859O9U+LEl
LkjCWhEH+Fr0KqPe4EMONEpRBDIBiZcC98wETLlHpsf9vEEhyCJZ7zqwPSvM0Q+O
r5F/jwYpbANlTudzX5jPurQaGsoYnIeXc9lAyqVdPG5ZaXQKflSf0Tf3Kn74eNd5
eWb4ou1kGSBzHQ2nlTUWRpVUr6E5QNxdMZ99AXw0tacsWgAsT3jLrhLfrVV9CBf/
47aNT5FWZgoHPtKRPNF29Jc9FRXLItw8yFmei6mfnwn60VWRZALL9nkHvhMVxiFD
KEjPJMhW4UqvoVhgIhBLr1A7hVRTt/ozKYUzWGkzFnmwtxrjXMxMaaUDDdJBh0Iu
59Ns4dpDxmgrYQfkS03dNViZDN25xEDQ1KuoudWy8PG9GMBP6sYKnlp8MOSZwJac
Xa8Y3dDVXG/na98OLeLsG6Op9UIyu0Bg3wkMI5FmIk/YLY0W2ph+Wfy+0ot3Kxh3
Fb1rrGZ77AexLt7U2BcMVPzrCgNUZ1SeVoBSgQFgt+F/tIl53xSsfQZ12CwflKgF
nIuG5+iMgE9YqNZZsf0hzA2GqKe7pQNcscJmReTSQmTW9vQVvHZlUVWl+zIDbAlQ
J+++Frx7BX+WaNSct7U1JEifw8pr4inkah38WAepuVGooFehbAPVS4TTBzdiTbu6
BrfSSnpwH8dRWZLTbdg79ExT+Qy3I4Nwfvf7fXSt1JlqqMiutPqn6cp32/bUH6tI
k90ISeXiJwc3ceFmIFh+cQGzcNKyBnrb9qGvcqSSWrm50YkN6qZNsJo+o4LUU65a
M9LuiuU1+OefEIuUf5jDopwazYhTQl1K/uwmXnnisF2ITcFGROAMYASyBCoe/3QW
8vLPKrH/YbODa/mz1caS17eAu9D9q2D7Kjc6X3NIeLpObvXy0kHdvOJCzGh0YZyZ
5pm/XgsGbC44qhXy/clW/zqV7tsHyV3/twwwtF+NFmEVPGPqDtuZc8ShEouX10CL
Da95yJ91AIGmUX70RbV6ZHraNAbBJqtkkw1cHNCm2vAO9ovh+UBDyXBqSzoNMXHB
+sgNc4chREm50E2LmE8ul6ZGQiSyQlrgDUkinEefeB+gvtfquyz5RR/qXDyNi4qJ
rHgqxDLiTNhwjaR9kPZayLynttrP5ZXgsgvAg3bm59tGu5KXAX/uUyGzKIQV31FP
NugoY8G3hGtdL9kCV83zui7/VbiQSVCBBY5YyYvSP4ragODSBzjPG8xbq3ngUnKl
4RFHzuBgZiGT1unaQHGo/KozRFY+oOm1TxdMGUMDa58zXJx/qwuBNJWy2uq3KR7F
wX5WG014ZhXzzwW944QB1yNizqq5q/ZYNrfoz6UUmVx0/JypYVUSiGRYiibr0U5Q
bw73G/DsSoOu3fNseW12hvWpJ9pFMa56OVDu51yaphmLMMH95dvoybCohM3xEHwe
flETEChYbRap8+j+u0ncNWP+iGQ83JLdeY7Lt4zQcZEbyMC/4xvqAAN80vVmmVwq
kQCj0LkLtddvZbV9hS5TTzRuA09fcFDqfuotg6I1dUWS0mXJQLRRN3thuZegCAyP
fBu90eFJ8HGt6XvFjQXFICoPRAK06Y7kmrlZmzWneMMKuGaAcK2y21vSwEUkMZaa
CerxVwsTUBxJKXNOUc1PduyN6h2PbyM9X/WTm9iW7vWtRHveDdLKo/eLrH3zw3s9
/sNsgjgiU2YtFWlOFMLzGmasFl03TUYV1p8hcMNg+JBCrmAuxUN02I1nc9zsv10v
hb2fpWfP3/efGDzPSnSTXBpMmvnn12TEBHfscS96MgcxEkVurM8d9GtkmqUZwp1M
vIjO3DFvWld47M0ZH3N4fycI/VRUOV8GK1FrjTdKMfzYPMsvc4fMkS32Ayw3iHkH
mJyfuReO+Zsfy4Hy5seB7dktSxrTS7ebJ3VBteiQkPpThyvH9879W9DtVMaQEtjC
X/jyM/S8tka9veF/Q3rHYIYUq90mFSAXs9d08jVZCqlXVr3FIokfpSiHOLoZaOmC
4YPt6/t+1Gw/1u/09t3gUnK8AySBdRtfM8Sc30Z4YLxgQvhwLCvwxd7e74xA1oiV
8LqpxXKIioB3yywtMBPPI8S4zytagVloBcgcM0fStGeN+5Sr4/9EW0IoDz2Yn0cB
jWjOVOL2lZwKB4LEMm/ISCXIvbqzOPtK1vGp64jvadJ+iE8kyuDj2VKn72goXOQQ
0M2QNa+ZDTdGh5qEZ8QEedCfr4cohbBZMwasnlv4aduiskD6wu6qCc4PxL8MtJHC
2M3t6+NS9maRRhtRkusDjEtbTFep9wPLhiBHKgq7r/Fs3i1Llc2iziu4ad+3fU+D
udtk2K2QU3UTv5QcGETTC6pAGNd3FMCt8Okq0drST/fcZc34efU93L0wcN91Go1J
S2vt63nIIF/QbHVbuZUKM1JJGj/mV+cZyY7D/AiAusmdSsFnhm9kx1VWV9RPQFOO
7h9Y5oEBcKkXEi/deQv/jVVR5+uC5D4rTckhg2ICeEaAiKQd4TEfHdTVuC7LXSV1
xlk5CY6Ek5p6mbdZlUwl4xtQX74kwnuUGOhqObcexHh4l5RtJQ4ttPXwM5O+0K2A
XOTQoFu1N73Uec/I0FOoBvHpof/7brjkTac9ALS/3+ZymYcn2Qw8ZyFZCzGoOpFy
cYZ5KOOyPVtH/1sgjCDD+ImRtoUeyvZocl6iSd4GdpJLBOpw3BrJzqICYdkyLPAr
9lTmUY95Bp9PyvvnPwe540urHTuia5HWsq3vCZ+z/zlIxOhaLOhGGK8jzBfCca4h
F49CoNJk09qbAdGVshz2PAC+NdK4PLwsgWC1zdI4rh6jczzwXpAFrGP7N4g1b2cQ
5PCkgBYvQ+AWvZLZt7sGVB0Z8cMt9zuy2kSjfelhDx4Fe4zgKgx8PX+EP6HtjcCT
LNO78ru/+oXbm3d8rstXzqjvfH8wdZNkEDAu5W5o4oB/CWqkPSf/i3RHL5HyNRk2
Pasl7S/IJwRAz3MZeGtYm1k/bKWqK8CgFqOLlegl5HsgLjP7UHyguE2W4Pwrba02
y1DBq5jS71aizvrwG0aSaOxXWh8rJ85BIBn6HRLMm8bCKcjma3Yqrkk75w4UJub0
C1O04+jQfPS6wZlYBK7yqectE+njlQIIqjlFt/jzxmBTcQwC8xBR0pWSi1WEzsZk
j2IUTaPGnYvavCg0f2Ypff/Ni55vHDeaKRdeN8eoK9zdFosMb11ErCb+AjFFSMOY
hqvMhP83vNfSNOWOfVS9Rnq1FwP3JVM/a/7yZP4DVl/jSmPSAU2sxlaDz50XqkZJ
lWCaJO0GcTcmlBFgsnGIosUELb3H7vkFVtaJp00s1s8LXkh04ZNkcQHMvL9hIfyo
Rgufsy3sMWoJi4Oo2zb2D9XmI9RC7PgBXfoRz6vCBmO8TAfit98GrqdFjlv0n+hB
8DkSXAa+F6olTqfvEQS/amTWrdDEvDjicdqbOCgQIiM1XoIacTA4pQlIixSeLhjc
GHZzAHs3rcBdB7Ttn9skXrfu8dSZv63tAjnsUSgGLffxuB1YL7+IMN6EnesukTFd
PiA5mkjrvh4zJO0Yddc6nk4P0J2qNdCqbMIfDw4qg3d63wOPOfW7liv6Y5w0yVJu
NKhO6S6WTSt/7uD9G+J7jYTuQ0R9aS/2kQlEblpzWd8xV7VT+a0C+fyzBSqZM5Eh
LkVeqcJXJKkYQq4gAarpLYgVDH7Jj2Pu2i/zOlhGAjgUWxMRWdnju/AFyvqeoJQy
WnIMqbw4uTZnyAZy4ouB7wmhlVLkxpAh7MzXL+dPgBBUIf7SX5dVVmvmJQP2oCtM
EKEfNQjemVMJbbrKOBOxzbgWP8WNT2sl0McPiYpywHHXzSDAqtmOrqq3FS1qw1Zq
ei0iGhz+uliIYA9ppzcJG+kmADNM2A6TfbKo1eFm4BxQt7imPt65CHKsW1UeLNga
TKKt3WSg7KRM7gSsWQRfDZdCRwDnvGV/X0lVdgqjUW5IqP+B+j5HqNmT0XtZWxOG
q3gjW35PBI/kAiOh+fspPymTsLf/HdXaQRX2demJVcda+GHO8YTVfkm9Vv7ssxSC
ENRKSy2qxyvMgcWUlUZcqaD05eQ6+1XOm1fnMJGb61OVf5xXORbFq+uDdLhbTr5V
/XJFSbal7dNcx9wnBqOdh1A9XFjfC/yZ+aBF/5sWO7xxrHPzOmgesOBlNYyauKy2
s77QAn/WsozWoORtLLjYqBbkE5Ut2FLOHVSjxzwcYcmRTFIbQc8vVqUUA1BThqRy
74R8IY2ovyhQoSHl5nfaajSyYfskFrjRe8zQj8TgLiq694ehw73uc5G6HJqmOQIB
DaMMTQU72zl8s6dP1ZdRKFcUeUKBkBbsWumKSVNDz+kf1U+SGO1NzHf09Ef6xcXn
gko0jy512We4qnADz+Ctop8GRl+4aY5zMj3Xk4fsTf/p3kr0UyYj2Ju8ck72Zs+X
+92gf6jNzI6URxIUqoG0hr/a+tH4rz4l0M+A8x6ZwnPjlLW227uPl3DXa8fuL7KF
jr9TWdrAwcBdo8Z/AQmMiPsaMw83vqKIgREDt4AqGXRC5Rn9scQykTQe2HZd99L+
toGNHRcd7eHvSvRxrbtO56CP5+ns3yS9hJonAxoplzUcRB+N4QMzZEectxg/UzeH
315Dmyb/KqftWfqI8R9ZXRxZ3/I58xDjE7HyW+0oh36uTckVKIv+naVPI3d9Sy+e
ERApXTx9YlCIcdc4q0ekKPRvEY7yhmOeWIL4z5dTdyhbaVDqCIk2DutquPyTifDA
2nwkR21rglb4zTGBoKecrtfsSj0h7gGaQBeznOm2MEptKPVnvszp2D+df1aXF7Yh
a1quy5mVuu13zGo7+tP7oHbsABTqHmTl0YoSbtkQfAWlvPBiWnUxEoZ0zAHHpT36
q3e4xQD1rPvo3ZxucbUe2YTVC/JGkra0iqK/Dd/dU61rqGFxHHqQ4IHRWsxyqtxF
Cw1+FN/Im+6QZxuVvfPOnIMOTr+/+tCBAC0NZUcQSq46og9zD9073r0xDhPATx5/
CyjrbTq6YPPRaNzTQZJk/7LY5j7Tk0fXNtO5+V38mD8sEx0AT1pWMZdxrwacqSoI
lqccfq9MmVdXMV+CWRgcXr7TEODJjxbheJTLDbbnKxys9Vm17lt48g6kgcaBFZ/C
vbUDxRqv+EL/m8IskUA4KSPXqgO5qc25d0aZqUXg5TkkIS68fbRG6FrTkD0q6mPT
kBCYMmFjldkYEpHSTpBIRFCthnJFaYOanUNfN1DVS83QTo93d5RGS+6XtqOwmmTb
h+GPtrfXdd4jp3jAav2JVUp8uLyN+Htd6KDY9rbpDikVBej4QCDIflzTu4LUOa9d
f9zLlSaxri9OR6Xq1+us6aUtGy4MzTl5Pkt+akibHpYMAqgSpNup2pFWLt3YAai+
Z+S5RD4mo9i+LPLEc3gKQF1JwKmoxdWGIM/EJhM+7YiN/4j5ZYZAazhBPQ+ctfKQ
iTtGMbj7MgkjF4uOweqwuRXNr4Rq83Ov0Rx6ZD7ZuMr7BfDkBSXcHlIq6WwSbG5v
yGoCeNPXVevOXJADGDezOozkSs4+UMwtAj0NSJP/jN32B1zW14Afmxisk+n7nU15
99FipNYXjD693xw321de7VmNb3E3oG0D/zzbD3mOgpmO+5MT5X7ISmV9RpSf8rBa
yWpoPX9MGreIUO9B2sr7rpjK5z26LFTAkSGJ0Jk63Nyoq46CakWLnOe+K53o8qpA
Pfl6Psqz9H0UGClPOvOvbd9a84tNIH4lnLL+J9GVqq3esYTnvWsU1/tAfJFqVhEU
kfQWSsBAEU68Cm2dT5RvK5g6SoA7Fpdz3GztCuoCExE+Fr1ha80iR0E7q6wbTdv3
BlcVxA5mvhq/zpf0t46maf5RVBcsIG1AwJEHDyAOKy5GeUb0B31y0JDpFABEqyS8
jzDUFmtPkBrq99IhfQaLtpX+447km55UxFnn0KxzbYWH3UjIIg/onfX3KiD/O/Cs
xs6+d61t0NLR18gyDYX/cR5v5e/gCnF4KK512sUbtu+BMy9naDPBYRfT9heAIu0A
HeOm37hIok+FLwNs1DmtbMD1nzeROgTjUpTDRmVLoLaJkB1eLQ5BWykdQpilTfBl
ZSe9xUmjCXJ3JrAj3ZZNHqmYYp6gO7xZa3hPMolWl9VvH0VfCHdtwQwnkEbwWGBt
qUtjdYrj3jqhJ0QyZN4xJMvaGkjYpyoAl4i8lLGTMneqVT/12tD1+SXpp6PP6A/x
TnALLlQFgmyuTKLvHY8zpvVnYFRxewjVv9IGKJcNSc4ri7ecb7L9McQQPo6clT0P
lSlEZHos8tzMGOGFhecmCEHv4YY7SZRlZKFupqOzHKSbUq6FVTdpKGwQxsBDs7Na
sOnZ1lUNSpa/BXDFuSFNQHaKbrkpy5xYzRwe/5z4U3Oi07ekx5sn421L3ndMdfBd
Rtd8PXCsedeBmaSYMSlhMZ1+Ak+fudhxhAe46Ffg/D0xuOwC25N5hnuxY05/R6ci
VhFRQXndHmxajHrPAk/uG/e6mfqyElkDuR2UtjN1N6Dbza5llUD8a26MEv1TSp0h
LLBD65tFovlpRSdtnyJGxnGbEV4879wFRLQmroWyj36qNo1kK/MxvR88SUjc0dmW
9cGnl9uec5mjogOCDGgV+DYt1djag4XPcWs6lW59Ro91lP572JxFHU/RZ1W+L6+p
hlrn6TvRBHSc8a7xmZBUjJ/bb5uIhJUivBXyQV8vZEWhCOFM8R74RbjZ3VsjX4GA
wPZmCaOseQGDEDDFT1m2NCBd6Vtl0GS2MNHNvsrBDZEOAs7twCVWoBLtdH05U3Ep
MZBMOJxpKyhsFer8Q9cXNC8Nq2pgQnRZlPMbyuFx12xIdSHK1xVSGQAmWXtAk6Ho
YQOqODgbGXwTh6ULbvQU89pmSSyha6o3jC4pn/f6FtK0Qna1faxcsZ4Re/CCt5LO
nnXLVgw8FsoDvAzFBxlCcjj0ZnNxyiAcnU4lHPEP3giXPZUM/rEZJtAm2HUP5Ge/
yMaaTHaCJosTr9+v5NdKakoswHlGm631fNMxrAkGTJapUSSyt0dU8jeBuoc9z9lg
IIJevTjVuFZCTTljYsPGqKnkXHbS0z0/Wx2ug1xmZaQvVI6eP+4N9c/uzpHIJNOD
fu4NwgzhnEMW/OTNiFOZB4KVsUFv1bPy8IOE2bpypyyeZ64BF+UHcIQyo89m/4ua
T7+L3kqDzv8olk63dpwM723mwQCbl/O8myNqt1PAkErQPu2IKnfxt1Iu1JK2Hci6
WLmeHXyq526Sr9mcCSjvCAr61F93ksGKaV2DD0nPaKNgyiUfVC22ufxRuyIkkMcG
YKhhf9iYh4mAw92/alAxo7sXhxO5MDOvAPUxH7JC+pdIsywAW0v+aNNCi8VAP3JY
RSc/9CIfQcbaXpCALXKYISn8V6F9XLvm9473dSqRlYkGtXUVdR5CceZML6ntm/md
1vi8Sm3LjzArFo7U3SISb4ZVk9jef0VGrAb2w8noR9k0FhNnBw3OmPKBkIClyrzC
Z73iVWB9af0aUc5BiCrU6Yw5L1vQU2ZKE8IhoUFCZIWrlTUFMFWa++cYhgKGvx/4
BZ6MBVgPFXp7Ajel2sEtAlRoPiUDcbVVhPXmTp7rlsnaVRRhfKQSXg694jFOSK65
G5wawuDe5EMOc09sOTgIbrKtnTw1PbeQvuhjxiLmE/hkS+4VOU4e9C/uWPz/a7V3
b4RHc/LtUBsccNqkFozh5flH4xzFteF/wZ6Qw6ja7gMV+kpZz+1mv+hoEnqM4cd7
9TCyk14vpQ4NYGoVkRa8IuWI5vBpiheuOp3x6XUu3xVj1+CQuulBV1WB0IFc+Qn6
+h8cQ93+2PSiDrPYne4+/fkabcZgoej6oZG204qo1SbDaMzzIauoqn8eNS5d0buA
chqtmZJspZ6+Dxwo0tqyl5A9BR4dz6VWjxepIOjTOgWjOjQHMtS9Eu7eLKq9ZwAQ
8Qx6RL9fQ+w4CHpinOCvtDPac3h3RxDnwTZRwv5q84dV2UCaatAw+p40rg1z00RK
Nob94OIx0HoHKwXQQ9wuQFyLUYFGYl1FcuXTs83zQWEWYPUWgsb+nUYVukV75UNN
Go3hwwosrj+BxVf/ll20BnoQ13Bt/dEteowfXkcTTXSChUea2yoDsuYxVSnZIOdI
ThbI7jUA4iZW7ApeZ0kcmSSe8Qps2wT3SC7IVEAHlkSgYol9w9PnOQMHRbUsuaPp
S4C++5mglkYN/HLEuKAD2FKx4pwnJbbIewAgod9XUtCyM24EtxzJ9KDAdF9fATm1
sdU10LegKlXtM0KgQamSeysUv2cravlSFqLxUicm7282afkiFu9d6xGT4DMTCmDG
OxbKp4ptNmQ0bWdN9App9uRtinO+fAgOOEWf+5zXJluF8HznQrBVxCSnIcmWjkPz
3/bu7R4/XSXxBC8G9FqKbzDoZmd6uZc/Ch4MHNbi8X6dv0hHYtUNY9COSF24IcJg
LAsQqoEPYAoZH6RFZHR0zpCAModw6mSC2Ds9mXuTa4BaN1FRrmYumgA/cKpsSVgc
6R6CMnfaOSAlEP/4VQdfbQadvB1KwtSUzeJvecV5PXND+Fu7szfOzsGXqhSewfhZ
uAi3qje3k9i73WGSJYisQ81O5k9x9tKGgmE5zeos88LhkeeMfoMsT6OVC7nYyjaf
IGFBro5sYbio+5ic3epm0sjOrKN8cxw4THxrK9WjWcTUsBLk8SAESjx4YVwHt1bn
7ZUh11E+LSR9wDvwlXsEM8pHgV3bTyXR6Vh4qMDaJvF3cO2ZSHz46QuE2ip9V8aE
klD9qYzfVk0jB0ajduR6Oo+64rD2j4tgsmG5vdGDxZ7B723hSOoJuevAKbX3GcxK
tJIOarPfi9VBYEvK9H9RNAHdQGURSbwjMNw7d9KodmDrncyA/ZSBKrrA8zCsf3S4
GcGsVf1WoxJJbJX2Nbto8Ru/mYakNjXHFtSWk+HEF8wDp1aWT0He5Nfybr0UiP4l
sAEb3Oo4mVUkpHUa1S25gJ6x0+SBHAsFapduvL7gua13/hvDx74UXKbgIBBzt8s3
R+MEFabdBBkui97UcmqhnJO81qcsF9fHZ+jV61DLb9KCG1aVDX2QDuvtALLBOsrw
RQD60MUI4TkwCfAdaO5p/f4iRFZN2ZoKqxKaV8gJSSCbRZyi2/IFxmAKk2syGDm8
WJkB7i6lZ/VbawDTUDsE+s0exi2OGvdLqrpOTJV/wHbhHP4uea+T9Bic4DYPW7p2
Ph8yKs2tgI7nHaLyZiQabKI3Az8P7mKBuOh3yG8y4TyucVpOHx4f89ABNdhA2ifJ
6jG4PBfMkKH9HBGZM7GpIhogmZ0xkph9Dr9W5PUTVzrrNO5l0tR5DklsMT8WANB9
DvOMMbhRnOYGc0PTTNbnNF+AyPfzNjROXnKnSODf0nej6b+kEyDfTmgTU7iCVxdd
y+lQl/B1fpDgIpfmPkVsSbGdYLalMddKSdRx7vux3U9IfLfdjDbnUi5vAXxYdUdD
uZaWb5+fwOcVUwXN7mB4A5JowLZArT5LLa9v15/xDPZZnxMkgjFYIpRVBPXJ9Q7e
MFx/QfDI9mo99t231Y0R3OZyU+DYhCbxOME5lWqd/4Ne+Ia7gb/3iope2waQjjZE
t2/fUkUEq8qdbvq9Z5w+gDb7Yox5BrQbja/zfsxk9ZXdYCfcuDeqLjztRNC/BcZj
GbiB2/RPulftq9OCdVFkvo+xzErDRn7Z3GnuVgoHT6nst7ov/WQ1nnIvikz9A0Hz
ZbP9J78XzzJ853SAt6JvzjFWaBDIt6YcorrrqdixTM1U4LgUu6WGDO8/1ER4Z0kV
ECQrRElJqP41G7MGz3+ByjEAs+gbTuWX4ezJiRtG2lmbZvvLaghKV/rlRDErz96k
OuvAaC3UWbXlp0zUg8v98SbHn0MdIJSRpqm3s+CuRRygCp9xqx0uy4BydXbcC5Rx
mO3YhLfTxKl/nfSQQh2vqxHelCQPF360dBSd2k8nQmForyeZ/AEV+MSjcjipdfuG
OGfr1RuBOxVDp4t41uJx3ftynvRYq0enEbatZXA4QStslcLgvXu8dEg0R8yP9a/r
1ZnZfzUfZA6F7TvQcGaTeYzxidoK7/txHY7Eslt6+TfAbs7egRFRnieqknIzPAFG
9cPqFlvzE9JsHznO904J1vj+pnPWjpOjUdM9cIDGQB02tcAB58IgjROrY162sT9o
23vC6qztIGDXNnwonNVS6dGI49YYFmpWTtRlJ6NDe+eZwNnVgeem0432MPtrZWqa
0lNRJe4FhqgRv40Bgy3pBjrh494lYUcd5mSvaSoe5ceEkZTIQrjs/F6BrB5kOP1q
e67r4TuBH++SbH0rFQWbXUPNTxbZ6LDnvB5hYZIoHeKv1WzpptdgapAIGRiIxv5R
f5gWpvK2HVA6Zj7a+4HahvhifwLZDbwYGq6JXq8410ML1pPjH/cTKCvoJfSpXtGC
LiopkoOCdo0xwJHprJf9X9QJ2OFkzzCc+fhVR0leYIc42HpDyg2XIu9Bp1PVVxi7
PWLsbsDe4DSt9cEnnjF+s8t9mJvclN9eK4ZfVEItePG2bt0WRZHtJH0Hoh8OqKqF
0HWg3DVJ/0Mjv/el3jZMraIk56I6iP9mJhbOUAZFnQwTt/5sLwf5CEUXRfQWtNPu
SZ1XQZ/7NnCWyIaEPY34bX/5d5CSvYfjvPzzqrVmN8zrUVsuF6zrRxf74JFDsevv
QTRuBbMzesZprRAVGNUZIKzqz/wPJZfKYkx2Z0c+HMm+IF+EzGT/FwDM8guGfDrb
9f2GFP7FByQY0vIJaiP9AOSA7Lpjr83G/MMOTWJ0MBkaFS7uekZV1QwLAyyyqlPa
PNj+OlFDI1haxENQse7sLOzd4r2ym6TXG1uhi17qHQvzIAIInKqI0ARWi/n7bqdX
UyRiNJCXgATHg65PPce6nMvBpfIrjsYdyRBeMv9q88fK/s7FhWYSuQYRHKkHD+kM
l3loCrVm2L4q5Y518ikc8M1t6QNijuWFYuWFTw2ijl44UIQVD/YDCpYJLPki1OlG
sW12oyNC/AgJQQfM+7F1fR44UShKczu/ALvd0NEgePzm+f91BnleB4uI18rylXbn
4up/fQWMBMxi9RDH4BpeK3bPSZUvhKWA2t+txXsadgD6lOjjiF++qVwGQBKLKMp9
ueKu98WAc9FGM/lHqUzPykUdwPsY6kYdpvZZXzs5e412ZNvrRXEn49urJf1NDQSk
qR4MIX7Vkbm+7O71te6WP1cRviaERJDNoLP1lJQtPcbzJ00akbp1yPeuEqaU25T2
oKIQ3w+xmTmQSWuVHiPsQSFyKLaTf80PXpyqacMcfpqQQ+XQLOu6nYB9p9UdOGG+
V7gPfS6Mo5CPIThtmNuA07/ST0tOTpuz7GEISkUhYTQxi2uZjU0LjQLMUWaOmBZx
cTvxkLPoHfgDOeZNhHf1smkaAhV1gIAcwwRmwqh8vl07XMC7wCJKhRX+wHeLGM2n
rc0tgrRK4SIHZTFG2D+JUm1IkHM1PJVYFR3zSnszCJBKgmj9KDIsfgvXrxaQsRAZ
XwqfC2Dp3W2UkXROOhRy9m271/INsOX4wSPLXbzmbn6LhYiwXeONcJmIXXrFE2oI
8LHl/4NIcP7UAqUDUuL4miYVTTPc7R86V4AvBHSJGlsdswvr60ite3tg4blOWUN5
wEypi7f4aq0uu2oFf/46oCVqSAjMw2qhJeRZ00JpCEUE0/PjsH5gDh/1fBFGgIbV
EfYrnjpbp9+IgTOoONUaqChH1oYHle+///sJG/1XLfcZS8lKWl1uPvQNYcQdfIId
jBULkFu4YguPAu7UVwx8lS+0WSbyRXx5vdP2w7Sw6iEyNvEX6VPo091mGSpub7fT
aAo9L2v4SVlOdpoHG+M4HFRHFaoOHDHhhGLLKrY8ivmiBVsingVjJRIjkmXbNut2
b9ivYUczmMzOcJq2ODsmVbdrzHXBEX+ZKGCV/EvXYqCElo58lOpiRfTp59a9tfvf
bU/2mHaWfu2ylNA/qfiAQIgV3eYa7tQcfrGZJgvGgUCN/vqEGLPS4C19PW4i5uGe
rGvOwRuDZ9dZk2epvkI8j6frlsyh3ZZ1S1pU3qOPHrHRfpuVV5RUBF5jjHwcCTzT
4NK6M4dTiIazmTT2QUcILdQUy/QrJsvmmW7DoEI3it1IzcZCIdieGTNj49iXePn3
6pbamiLCSP7jSgJ/ESkMqmH4UTrX3rhE2et/Qe+X/uU6MfzqeIAuqFmo3Er+7jDF
0vXdSI2hK2kLK9v+yuwu8QJM2Lezwaaw3MNTDyOpLWVRRk4gfAAVXWwfrdkD+bK5
ZZOafDM9CRhEWbwOQN1jIvrt+3VDmAtbR3VTDrgMIAE18SVJYfvQcdwzv9wru+Iy
JNt1KRCtOWnnxeVtZXxsUdnkw3f/r8l4K6kL7CZGwIvgAE5OBd+P4Q7By5jxcPqY
ioqAMHvbsMMcRlYQkZZeLwbLnErM5xj1dc2UYf/XQQcTDDhJZD1iDkR/F0VgoC7t
SrSR/83gDz0Zy7lQuxpISECmdKyXpYMAU9cL0nq2YWjHpGimVrFMImQ4pqrvDG0B
IFGhIFE7INt6Y0E0iWTJt10Z4I4YLcNP2wFyoX7NnyyttryRyXLgcfyC5gNaY8B0
CIOKRObDurXdGIq5kg06BwQH9BfwFBlfKLqr1gukpWxxiG+zLh69GFuO5BSw+IUz
8YQlRINPv0dKzeshKfa0+NaecB59GkNaEKVumtBUXzomD90VrT/picgtUR1MzVzc
qt5Neh5gg/4nzrFd9q/Ov/Y5I0dxN6VJ5ToJxR3fxzkrjH4cCxDTS5I8I7t9S541
HbzzrCLvXOHns9pTCPR0b7FJxbXgwzGgpssktlSAUWRjca2sHQXzHA7ZujumRi/G
K5L2Ax6SAjRoptg8n95T0EB8aOhaoCNu0qR3nCN3JucG+pvePIOvX8aCIHI4lwR0
Fi4e8oVQWOqfJFEjk8eKLORUYX2EabkmX8N6S4yb1Baqs0Bhj5HwFbJlttkFUjw5
NPcAuNpT0c8QWTppHwHA9mF3CAVpr4Z499ikG4Komizew8k0vl+8miy1L8SqzsFO
RLLw8XEngfZzkTKcXuZPyaxupUgzCVFVvNkioH2t9rRJI5lL9iEy7doD+aj/2DYY
VVa007d4qVds9nHvb//TVDVD7EudRJgnhk/TsiKqpbo6mHvBKR7qP7XjahJ3Shfd
fppPEh/SqKJV4SnBh4eCk9q+py4DNEmwPejxiBLcfG8fdzxRhoRIBwxR3TZQHZGv
pX7SOP3nEr4R4RUw45Kzitcw+BVUiQpREmkbPiiJs4Gn4En3zr3SIgyd9B8+EoCo
jTKik5uk6W79dZMqnIHd18hQY8D56AYFEXhlp4l3CaRYlsWN82Wv/iFDsbGBTr6Z
8DnGGUWXRbXAyHLG9BC7POHHQnnOrZBng5ABRvyq+A0urvU66NXH692mYeNmf3eC
gDFxlBHTS5t6RPTgmsbarF3mJPDdg3AazbQBkIbpj9tuZAQgVB4p/Qd1YUzVrWi/
B4Ffe5i5o77uu4i7YExc9O+EaUyxImVON7XEpVOGkczXVACzvvQqqcJkYQMW6FQ6
Z7ameK0xYVHOu9+M2IewIFvrFmM8kIoyiWsZ4lbg8dYR8MLxPyc4m1CodZvL+iMh
+sXh6M2tydsEgQD779Rvg7BI8uthg82k0p6zyULjIe7Y9tetX+ZIYZLd5VzWkTdX
QL9wXwXUY5UuxRJEp0SZp+EjLdx/ABSS1zQ+kETp8RZHfIF0giAHzEYuhotpS63u
EPR57VmA5BBBcZHVTOnIL2WaRR+cVtn2N6+awXUAdQW4MtUarj0iC5rSn0VcPh0j
NnKgLp9uIfjT3HmDxdmlnBfHun9Z4ERN2tM8lzInWy4R+/XW400WcGkFEYNDRgSD
JvXQVMhYFJbR16XsbaLwROOyTeFCyhP0tyX8C5ediNia7NyCjaSPdyR8enrDizjl
XvqRew9+FIxVBaBCvJoAJO/5V7CNAxh9g/OeTsqAQrxBvV+lH6RcbabcdAhxKUif
Q3lpZq4sWA4oqaLL5K3fLgwQ1+DUKR+nBZDo++SNCGVKHkgzu5epMw0n/pNp8QIp
6RrgLSrjz9XG/jIr7+sNRkXf3tOIFOA3ZqvHAXGSAc5m3geQl4q0OkwDwphVzktH
ZLCHF+bp0rTfhILFFKwsGjgZrTLYXtfAfY8AgY42rRxygURNElVkBYInjzeRBe5K
5HrW3Y38ScqqDINQrjByOK/fc7IPxBZLLP1fx1UlzhNBdMM1jGngjt5vX+nkOsH9
Q6JMpNt/iQ4MYQoFNlsdjSFtx7OJeBuqpFq/Ll/u2t/djFCt50UvnGHthgIkFTsB
rMe8B/EiwqbSuN9CcYQDu7NTN6NlcLAb8f34/5XT0br1k8bi38e3hW9F14ZxLcLb
XxNdOMsMkYHeRXE9qTDpAvlQaJFI1RDWCE41rTr34a1edzbVwZ4/dpsYbBOmCkst
Bx1FKWorPAeDtreDXr4UmOzvBTSFLC0LdRtK4ovaSoRCCVpb/904x+0yRuGs9hM2
joXntOAT9awNT4UPG67VAK3WIUazS+uOxembsjtQE2thVwiuQ+vU7r/ujtIKEedL
iNQHwPz8rxlASvEYKH+IZHia7fFNPwxQpEuPAkK8BXOysRRJOC6Nh9zqE6mOwk1M
J6JSbEOMJCHlT5r/6hVNtIvszuGFGOPf1AqLBu4PWzQMhNUlpgVNJ/Y9Xr+aC6f3
CcKCEXEVKfGsGA60OzEnJ5M6l2/e38m3GuDzFK/iDDJhKUzD9uQt0FgqsEC9NZI7
kN/havaehoH6w7cucrVFZaOhEB7wYF3OGYBLEvHgfq34gTzAJ2gv+3Bg+bwgCzUz
gtiex46IeKHmuNBJRSFjISOdFTPouXziM8o3OjwcHNnx6m3VBL7Ozj6vEx1b9BVs
QmdqRQT7MA2HBpN8gkn2IhjnaPehWxaoDPCSoGJkwBaGpfmBWEkEKUfUEASUvpY7
6bD6LF3F0uu0Zx/zC0ETePnjrKH1ztBVix8Yv9xBBFws7TYiSbtSCM2zuT8bUfBd
xfAYtLNNhk3eqeiR3nH7q9rlZ3e54Bw01UWm2vBkwaDBDBlJxtFPC8uLNDVFm665
T0CN+5dcvZx/7pYd0Oqhdh2L5Jna6gn0k/yzvsMcDNt0SgBtgc8dABfnQwtD1JNl
JSItxIBD4MSS3lPDG8bfmv3DMeU0zz10XYam7EIWG45A6cu9FdI6pSmHfWXRgT4H
OMTl2R8OS0frAKsSvjsnHfyclBSkNzetgcJuSapUWaw1nzTknIksXsIznNI70X7K
P9L6EqqdWtcssCFdEGn/kkUyAcToxwEGnUptg4D3PQ+fGmzuvL1dJKF5foCfslBg
FdATVR3qFgxZQTo8L6SbY8IJI8IFydTgnDHEgQidXxGi0f7gRfIz3yOXfScjmNzT
ucVilaMmgWMXizBQvuvxyB0t+UK9tmt6vSIYW6IegbvzpYU1AvUkk6iI/y/CAanS
dkhYgRpZcNjNIv6S2wdFNxwjNq4U6FJITdl7we9rrApy3XWhrYefbic9DvOpvg/R
Xo8+X0CYbD5A3UyGPmNa9iuqXk56o66VxHPfCQq3p7YAehC+yobNuapkAKoM+XAV
ERihH1vgBsMXJrgFvwpWHsaDMJilIPb465VZbvW9FKpW0vWMgjN4dHRrelx+gSzw
uVjmTjBA91Uqt8eMoYKoeEfGCjTPr6YshPMmnbW8Oh1ycWHLycNTHmpKwsxnNtzC
qksxrcETNePCEOQY++qv/DuXK3GMPqr4pBUg2/qkvJ97np4DDS6YU3vNwI113Lqu
UUOjhh1ROBo4cUM8jK6pAPbi7ShtTMunCyGIjSWa0d1rpwtpZwj8LouYzLW8IAgG
ozCQSeen8pvjbi9pTWJuoGNJ2a93Gpb0InoOu6eK7LnprgH2Z8n7/DqQR9ATA366
/azlD2BGfVV0Oo3264L6kPz3kxiLZR31PRSh45ZY6+WNTcrCg8CDerII3SEFkGvm
muFAqnh8SCu7qKJ6dgbS+/RkAa5EG8lmSPULKVTwdivj4DSv6V2UtR33JjU8gh9Z
dHLrrVXvQhUMev0kI19M+r5e11Xn86ULiSc/6uc6E95wxaExitNxvry2giEYBlhD
lkVvvKM0jUA9LEgpCEZgW1TNL4M8viQmVVdII7RhgU9FtVkx7FbWnoQl/+yeb0dH
merCvlNdoAkThUqHWukZYT9Q+s0VHjsaxn1uVQUGVb8a9atUK9jBE0B+IpXOEVgP
DrEN+tTmZEmTYYAStFcemETNLd7czxVIEQ4l+AZcH8GG0qtkhL+11gkcFbMnu8KO
Ca0PMIPHuYw/e1JCEK8F0lJugScchcVsRmygdBR3+jCdzDfPdGhbP09t9hMHoBmG
bVajy5SKBO5Z/Rim0v1oHQBFe+ue4Zwuyb7p4SDiY39moH9lHHj7IxQh8vqBga1y
yEahpAUF9mB44Bur2Wi8al2mGsATZz3zZX59wGDWquCD1a11+Wugm3GjmmG0P+ZD
4vqdWzhdKzDUj2VYeFYRR25aXSjVEhjQVYAepB5BUMZIWjoYmAJZnrGBY4uKqzYz
dHnXt+OpAQQHIfbU8ZJwNjrzv7d8Pq23xtx6TYyzS7KOjq950Tuo5f2/6JvGXHCm
VPBg8Cr99P/jK8LVYqJJW6UnT6CNfe6KwYa6JHVKpfV7SAhmL52kSvDm/hlWirMx
lDDh+nfB9wJLuIEG1k0DP6MEwGvtlhgRY0S4mN3QqUNy6Ew1M0ap5yQcSLwQGfvy
u5ezUjbUXUeYCMlkJs8GxgFQKRmcae63P6wwxIKGaHp8Q65qXwcaO2vnPMm11zrw
I7W7jccNUHbgadOrZyYTQJIWvGkDqIQ4lBj2qoQnJKhoYD3KYas8mTT8yzN93kKN
qjrU/RG5a72oye4MIxyxfV4BOKIFSyfP/7W1OWz5qp5fACKl1d6ngA0eRur86p55
TsxNrllh0TNeTlJmaFw7SUXCMuvrx2yTYsGbPVR1qY4tSWJApnMsDtFRvEMQhjDn
Lwj48/yNW4TeOCIkJIhqE9QMjao7xrwQy1mAU5lep9uZtVIor3D+RH/nChPscF31
/h6hbgi4Rm5gt8XWtkF5kb3s0ScFGH83tX7Z/TcQEAMw0gaW8redYgW4A//ckLOT
Dn3r8UAKz1p1/8RdJKFaSMz2Hw/issLBP0CV2MTlpzbb9xHDT7Pn8S3TVwfJ8DuX
52YvPGzyAwyK4e5Hnf8bw0ryVHtvwQt/ppDcUDXdjEw3bj+8k4DBnJYa74CV654/
xxRLiehbabyB3BxDnwVA/05pObUjVhIXzsrf6UNLigygX6siQ02ZuXP0Pnclg1so
5bD3AxeHpwimyf/K1lbjzl6vCi/fkUTSfsp92xR1y0HVuvlX0ubAAp3/F6PqVZgU
Z148wOawYZUZ06wfWR0RUigNB12LeuBekWHKlUX8Rr8JemwBU3TJWTVVIOTQFvDb
Z96R76yrylgE/naRSz6nR1mFoU0SF7dHVXji78GH6LYtnPgN34DMF+46REeyQahv
VTzJxzqctkRQxwoj3xm1/rBYRZEhsC9m8nY333/JcpBvITeqRhmy1jh3pU8aDkwo
E5K8q4J16kvQKAua7GjF5d0SRVeGkJnz6jc+baw9vrdbD5U+JbkXQcdCgRh4iMCG
5uxTtxDWBA5eDFDfQiV0L5zVL+ua+9nrmuDJVlgQ7Kdy5loS8lWXZkV3Vt+gl/SO
O+RqpFEyuUZ6sMLgRSw9cEeiqN5jbWqYrcb/QmQtHt5+wR7h4ERa+fIrWi/1PsXw
KPQWoWuJLcZzjLwThERdX44vl/Ho6FH+/tP/dxotaYW9Jh9Sqc5MKOWFHn8i7Yc7
RxmW3Wkjc5GKLLefHWMFY24FFLR0Rajplhz+8yoLDq2pddZDvlYIXLB2y1jDZqhX
041r4nE4+8a6nzZEr/08cNYpPoJO3B89RXX8moxwn63R2raZM0emoPi89iW4Vufj
M9bh6wdcd4GaVMjS6lPJHGAtoMNG2sowk9bQwb5RAeUEIUF0wJdQ/TcWkNmSkQ4b
xybHFuwi8DQY11EQDbQIzs3RcyAdulr4wGE3YTZueRfw+8zYKg+Et4zBY8S2XDxi
5dJUIEe+k5k7vYAhCTAOxs38oTrzr8YFw+MJMEUSvNvUamWteghzaN5hrU+FUoI6
5W0XUWuuiTnR+lALbKe8ye0sr3k6zFab6Td436ANYseOs/bnuBJAglxRCG1P94IM
SGRxWf6wNy7wJsQo+Ty+0X8VMb+WupiMq8Rd2fo2zoMx9j9JUlRX4/LKxRdiSd25
wRmnf/cH3JWr1ODVe3/TnxhBpHQjRStojWdbBv4yCWDujoR32eH05eS9y2MEAIRx
36Nk0uMIJyykDvF+eUr11DCMo0OQApau60ghSIiMVSi1Z8xRBNQ3wgcz9y9OdwL1
j1xw5rJMV4qx9gwg8aEgdyQZkAoYvpQThLHbMQDMv+XpjjD19ee8z4GraNFxx869
xFHMWvido0+IsOLB9Iid32uXeVnJts3zAFjOWkXPza/Pe9n+RDiS1RbjRocf03Sx
Nr5AZBDPQa5nMJY3Ekh4G5P/PMW+km1J+cvnlKnVHbkiWEgiTaWr5ZWwoMc93WUQ
bDCuFqx70vGmFriQWjbZI7PvekBoPmkLa+j7DUFbSjx7jKOwbTXH3EY4iWjRtStG
Capm/vTc/m+aoQB1JjTLbyvJHzGVW4Wq0VX4ybET4wYc47C0CEyMD6kAYd47jn5F
qUZqOKKPQYv2B/7Q7nEyS1Ms+rOHoMm64KiGNWlbMz4WLY+aXIFXNoePtQYp97qR
oBmvZSZXpWW46xRh7NX4f0ah3gcWoghNpoMTzbPr5y2BQvsx900ucjYrw8wTyWtU
zPCgkKQAI6dpHvPhWpLYmdzXKjbO54xSpwECFOj1ChUYZOGBachhByZQmkzRiOh8
wP3NRg+oIlF7aP+yM/FRbNTLjpbj6IXw13OtE/jMuEftMQqnUi9xGR63KArqozsx
OZ20iJzV5vfCbVVp8o5aKiA1pfpH57aChYPIUEDsUNtw+bvaRt0LQyke79jsh8qz
1QRZ7LXY/SXd47ZJLGE+741o7CF/Bcn57Hyok3+hq/OrRx+BMZNquVThmQHN0KM8
9yTnHRLTRQwtKk9uXKHyxNOLIz82kA0Rr6dNnYXoFwHrQFFKtcYYfM9AD6nbxEFP
WYZOLJSTdPjylGVGlxdB1NVnAPchG9K2jMiJ8IJ4+B9fdzq6Eu8S8ohM1IkjOV30
wVkJfRFUg2kW+jUNKaDcyJ8cSm4PYb9rq9XutnD/yl4d8ESuBRr9UrZwCNv1/AvA
bsSdFTmedKUlsBnO3XINMXrU0rvELu7Tw5lXE2JPBW3Hyl5tVJp9VZlSorRJFAvs
soMg0N7CMY9H9QFo3DsiCB9bnIGWP5RxOpPs64MCPIZWdJEK3isCW3I1FiGKFOaQ
WSqqfjI48U0JOToM+RdWdFqy1H4E49l6634E8Nhn1blQaECW/oAbLM7AscLgPjVT
DuweSkjr9ffk1dPmJ7uCSeVJWwPLZtdRzlVG3Uku1gRqrnR/Py/muszOglbepFmR
GsTJNC5XicdGdhNl4c8dtnw/KlrD8j/1Z0hIknEj2HghoZnRM4BKsx+OHfoQv72G
EZruuPjIpFnvX8vFu4UeKri9XdC6k4tN/ov7N+vb1phkGYAssk06SqLL6aBYgpzd
R5YCKf4p4pdoY3Un/P2IcWcxABCKK6nok1rZMriBCBmqQYpYpU0lRdqvgNRaS5ob
XfFRUp8PVinWLhX5MUy/sMjdWvsZLfm6eLgD2x8enGAYvnZ29fh7u+9Sutxtr+C2
pspXIOBTU8HepJJFxflPPPzCQEja5E4DlWYrLnIkHMbBmHGOcRj6Hh/mHpINHGVU
7eMuePeUiukAbFr/Qeayw7cOceFYRSpCN7eAxz6QoOScI3f4P9/Pm3+rRYfFxAQh
nWPT9oNM4JwHy+vB7JeVUu5jUKAnJ60hnlKUL20UWvPRmdutKt45IxDbHCU7GPHe
trGBLr2p/T4IBiFvqifJ4epcQ8yeShwHCP1OpPZdPwHjVaUp+WowLtGNgKqYMfKS
LHzCS70hxIXkI4QAnTiBPI0bCTgMCAE+W01sRGbhNqhUlVts4LckdsghijLUOBkM
wRASvZc6F4Q4giCIQReFjlLLz5Y/u8h/MeIBCeVflKGeoVnbN2U2wPiFKPaJ4zpR
QuKbOMIsE5Xe7a528Pl3uuMAyf83rkZOVjWopg3r6uApPSi4AHoIzH6mXUZEjrWY
EiJoiTw98Ji+VNX6USYKCKaeDlUvfBSebst1Ao/Pb3ohrpL/hbx/5MERQ+ulijI6
cH0yMvHcErVHz4a7vMJxn/FrKvzQ9bLmJvyFt0IoppKx0awdMSj+gC6hMMWE+tJX
WNJfu5HSACpA2oCAFwxo+hbb1x93qXFar90RHvxNCZeH6TE9JmZJAa4wOz94+hcP
KYMLHOVBr9DjsyyeOpa6559rVjdM07OR1PcNzX2w2WHHkYXyUq5zy44VN0Am9cKc
NhuFxCwEUJEs58AtdExTy0d2R6owNduXx5TEl063uElgxU9e/LP/8+LsxpiaQtWA
Lgx3YLiY9Ii5rIo4J3yCgBTKKWoZfnsFCOEgE6DDiaYOBytd2hWUCx/VnkSK/4JH
PUBQMR78v4WifZp1eBm0luAlxxKB0hOQVBRA084OszbrT6HZwz19BA76d20MKazo
g9Q0wTJxJNf3vIA7TOSMWVmPtIDx1zGt7iSfQU+QL00Z1wu+20mUD9LhSdKwg9lQ
ZX4GfDqLvbShks4bhr2ZJ5QEDZlmEwPLToptMDcZE8PtLZIe1Z7Z7hlDzm+47oML
XRkhMS59j96p1T26PAoQhwH/ezJfrK1EStAn4+W1pHvm8aRmV64WuvA8PIRGN2Oe
uNa/ctySoiVemQnyZcN9pBcxewZZaPQkLm6mxTVSZmTXhjZJetsrxjafEr3GS4WH
9SvUaBAeJqEtIZRKyZ1JjiBOdheFQhfL7DgD7vDAQN5FviS0mdNagHMCQIGWVlGl
YQdIRYq50ZWtZCTztPHqjusWhi1ZjxblFpV4YfGbN5AfHIroe86/Noq0QnxasaAP
RG3fIUHt9TCES/uocNw2kzpTgPJqa/IU4lml7BYh+CpvKEmef/ouhC9DnoH3mZTr
tVB/5FF6BY3tlZJRIJ9VUkvHvJ7peendWrsXL7Ao3xUvqA/ViOZa/H9q7kVz95HN
qjkl+SO6PxNvkZlba1OlcQMJD95QF4lDmP/BLkvIdqW+UJlTdxUIVafkj+S2V25p
xoyjQIm04y0YtXZTck6BI5EfyzyDDUw8rL3doZhboNDKjF2l4F9PbH37ByCOtaXn
8r/MDdCLst1MIvit+XAdZtFg+HVvkWlR87UgM4xmXP5lCKvDMIZxZMjCp446ThtC
Pz3VBUKJPTBmiirPKTz2ZNix4fuSGuYFp4mQyFKzZoUmxqo8Xmoq2KXXJaSUjFle
G856X0/DXtzcgKfukDJ0AXrCceGHTunLfHHSFTlu7WojoMO6QbSWj+PQ7nL1rJnK
aJR4YZJq9uxc3vJZtcifr2Vyerf0LMK+wLVMr5SGV9lQEUH7Cfp47/z4HieYG/Rk
6HWp1eLTjzu8pmmKSFZKaTDLZAYiW5tDDzAsnXe4iUz2V/k46PiBpuY1ejpz0MBe
bCF8j+5Zxvo612c02WUFE3Kb6WaSA9wJ7eS7TXj3EE7qG1+wHGDgirZurdza2X5z
R/rFiRESsNItqMogRYANEDLQ1rd6nlWj68NT9usDMJcBOviEevZ3ABByqPP/UrXF
UsJswhwsG7Yv/9a71T4AzJO60H7usBLrD6I3Wa9UfKyashc5jMpvMdrmhC3MtxPX
al9BINZjjBMAGAmbPKD0XyiIxnmeZb1zp86xsYrM/ls6SXKqnAzUmgwcOKKae43/
KUMtIFVxPsxuRtlUAhxbKUzIlfM0C/2BnvL7/VqcywLIf0PiAjR6QEIHJV2PQuAq
FUIZLxE29FRdbmmwlKhNkWxuSeSLtQwfeq9GslGI6a2PNVeCaSttyAVgkeVuCfIa
l6Jjr69Sm0hb+zOoEJh3YBSaETvzEYI/yr9B5Nz7o24dWhTeETsu0nqFphwtgGNE
w8/shZUMPY3PoGT8+O4fmEYPqC/JvZKoiKWCx16BrunyRtReUOSUTcRtX8eyKP3+
KMAjPTBPZNc0g5eLSPsKifb0NmTigrzOCSvX6QnsloDuh024a21Hes/AW5XONyes
zBpOchhMMzr+V56zYwW2o6pkyoaKlDsWG8pMiqAdqLIZ+uJNxYzn9M0eCGpzZe14
BVd8joAw7WDBH9kgSl/4W38SI6Vs8iwc20I/rw7OiZqnfF4lDdgdmPtnYg7rJY7V
ZmIIgDu+RCXff7IejyRU/P0PrtZ9dNIJ2ldMpvGY8BiDKj/T2+lycI8UHgwSDwv3
Gjq08Wtuc85waBFnQ1zsNSjHGTHYyv/BuICR1wBSUb4jL3Oe2W6AXzS4L7dXA1az
dcGPQURMM0mqO5OVjMJyS38MTa6A4E4t/wVZAZXSF6CUWaOV/WBdRj2qsIU4Uujd
MRXg7EDrAZuowzGjKCbwFoEa7d5cZHIaZd3fRCEEscn3DXgclwJB2/vr0tDb4PVM
D4twXNj6K0/J28POgiCUL+FnHwHPaaA9jWQGQE09y9RH3Z3euWciO+Jk/qKrzP4w
gaXn+LU53VCNatWl8haTfANsk/LPk95Z39ni7w3oxJqT36EXmnB9WCtlnMH7ps8b
n8GnIdm6P+1Fzt8rFJ+y6dE0pHUWaPh7mBLkgxCmVECL7xd2fQiloy9LbyegpLQJ
2mcaJOVxuu7weu7f8Zw2F2wKfAYRL5DaihsEohT1+mO3BNVOK+Eb2e4R5N9vGr9/
EU5KBgdc/lDIIjSeoMC6E7S+VJSwhAml1fwTJEdcMkmGn5GasCxNMjocjBD+3uJE
gj7wPwCVmtKwVtc0wDT2U5QxjEZwBW0Hk8GibM9OxiOJOuIw5TSDo5bYfgoHXK1P
nQh/qjYgol5aRRDCXunEcSnIPbru0GWIXDSa4jiPANaSqRIhp9ROo5YvwG8oIAwX
b+m13JZFaZVdxR9vr2HA9XsyUGoNl0rh3iUk3jwyh58yBjcJ5rTgVDpYaxouSIrd
/G5fohwvX0p0NzoNrdwrGn1LNFABbVmcRPrE0EeJPLK7QVVTLQE9FJLpCRcbUzQn
mT/tZbj8SOAd4I1GBY+yxHE5GIsUAamdZYFdKrBl+hgKwwY4mbSBwKKfnvUezmcd
DJJLyMdG1b35PGErVN+/otyL883qpRWXhfU1mpHl4ZFUQ96PeFirw+nqlQkMmaU0
DvXHAbpnMs5fxFv11iydNGDy8cpyQX84rjMqhPmah956+otrmaDQpRTxnJ+FQZke
2UGhgmEqXC0rGPZ4ySFXKgcczayOLUR0Z5f4ClFQwRNd/yAMgSl9stMYPEDDCVPY
HdtYa1k/zXjqxfZokdZCpk8G48QPGXhL6oPTyaHDINCZ+TWXqNpnqfVfFPNF/zM5
vfDxmNQDJnjgn8CJsK3S0Kmtpw9vHOe3EvzvzhW27D/3NiD/kBfLxwBS25O5hj4e
Vp/Txceb2iDd2ojF0yiRgzooE+G7HJiUthZGAZ5Kd4EzCALgrAGntoUgzT+PWKmv
w/EypKbCs3cU8G6ZpPcSDjR/39Wh2pc+bTFGPKkN6nfY2tupX+OWRYbdj9FXS6iM
NBh0pP2U/h9MIXdKh5qAGjKqoehGDL/stOohb79M167sQxRUu9Y76Ny0nCTVHqqo
wTx+9p7X237FznvCk7BRvdsTnfr/oSpxAYZya41TXHS+PkzNwixwTuSR7WayvHar
AceAW9Ck8IrEArPc+FALbslvL0GKbYPArL3+R4RE0uHZmfHlJIuAfJnuMs+/0eHr
LoqpLLT6ta94VCs87N1MdKeYTAxZzjdlvDCrmy9A8+pgfpVGraHXL0VNUhAb9IAI
cpxSHiZxTiojKDFApMSbyIUCTSPeF4rgqmu2dTJYsBSAfAS6BaOAi0u2IFXHPkAZ
p5SvtlHJ/3kGlcl6qVIhZjtz4yAQrZjP16gQO7HlnMYVjh5frAj7uC9pOLfI+BAu
/JW438jiAsfnUIO+xp1OTHhgh567g1QyQCnRafoaSt+KLirdm/25v9DV/85T4+4H
X2kmT++C0pJwOtyvmHmc/Wt0Mwx4VJX71TJeAqXkh8FIlkwmxS6AM8sd6ORBu8Jp
NLiEikovHUWUB2c0BaiP5hwMeMOcQ2/cgJPRvtBNgwtwEI/CNlJRIvDqDU4bwNny
II8xvOV24pAh6J+eLPr8P553q9HoK1jR6MeSZfG+4mcYwrDNff3fJ2pn6r9+DW97
Qt34GLM60HxBGA7iqMaUO+qVUimH+G3lQDjSjlbYCiqkfXZU/m3MdF7VqZl1Xysw
bx2whfwNvlOr22PkEA+zyTogsm+oRdqVbK9VoFKKsCy6jQCqu8kL1N/y1op0ET0y
Nf5AAkowG5N4T3axj3fMo63bFk2n89ln+h47FNy95WP+TMK7kbHoNYyYzJkMnHwr
R86pdJXYCkgwE3eQRSNJWRK8DPTroIB3KelHZ+d9R+GVRZtVRbEx8Bv6hSD+tuPZ
R8En6ptE+z5soXvwprELu0MKsY3P0j84p5iwdjzk4qSI/mXc5vsBebf3TkdCnMdy
afks4/mH0SIoteQhg5kev/zmTHMkJ1QoX/Y+msHwc9fMNj3/NUa+IP/Q4J8ltuZ9
9MJTbWoQ7TUTTy8wJO8J02Lw3RISrcI4cGdvjNx5NWpUmE2YWw1ddDUl6cQDgisP
G7z4ryA1vjCk3WjMT5eGKZl/8MqubJd1XqLsmATuYmC9sGnij66wbl2QxkWVwHJ7
MwOovbriTxoF8VgetC8QPSM/M4tG+fG5DUYGoJDrHkWxzyTAoc0OCaNiE+AHCd+e
41RhMO3nnWLqm+b/Km4z17NcoC41wbIizdkljzTiziHX7pedZ/vw9VlnBQaHVmL9
9AaxNPpydb+Gg5OL+lcHdHzzeTmD6lSJdn7/bgI5G6fmtE6eGBTNYELVg5KW5ujJ
v5a+tZ4Jk0mEnHkcrupJM+sIoy+JQbsiwpjk8YPj9E6tf3173lfo42l212TaIgJn
0k/22+7a1tFjpj1z8btkn0SxVMhEUlW74jBZzcD1WSNpPb8csaSlT2hPc4LwPJUQ
bzPfW4cuBJwUnd6gBgsYGDx0KBebkvO/tLxjWkenaVaQLRuSTvZhBVV62C1rrzqG
SvGcZXyoFaxQp75aHEBhPwPT2PGwCvme1qFD0Nfd1C9hAQrRcpGscHnrZ19OvKZe
gu2H1eHc8LNAfIhwFBpm0fqCYN+5W4pA08+QBEpwZusnYg1gg1nYbjq4TdS6qi8F
i54NzwWPDTUaJrwzXfJ0CHJRizN1qTExys0xn5uDHSLw4nJxPyPUUCHGAyLuUhdF
GWSkKVIKuEOah4kY46Rg9yfqx6FYl80nH8B4oJ8rGntxI5V0/fNXwHOQa2oj9meK
MOymgYCFnNrW6FNnFpI3DoAbdyMvK/bPy3LL3/+W7V1Bv8po8HIDkXDkY2HGYViK
TV5BHC6dFkv+gtLY7HoaYKn0f+DnUyamY0byMlN1z8a1OdYKq+qaFhyLulTJpuz2
s7sa0HnxThI4KvohMxEmCPbC3Ge+l+FH73IJrdCbL4PRXc2YMaBFXlUThQZ0rPys
79oyaa87Ge0zVqbnNotLhoPfZELL4nTu1+hM53z2hrS/0HIFishyDKomRCRPyvB4
Yaoqzx1CC9n5av2XGeDrslmS3axGME3PsSXF3AE7T9bZ6L4dswjs9B2jEKbXCgNP
FS/0GIK8W9t0p7nDirhXp5clISYyxvhvZ+AJVxayp2p43g8wrQSLfNEdloAqtSVp
TMXuL6e5qHoMXwTEwByLDVk+Xexi/32pHxg91tDSldmQf525afBcWxjLDUHR6Lh/
9YCR+rq0hbrqev+1N31ppRlVDPcmnW4VObTo1/D4ErfFRDDbQXO3/cvheMT+zbsK
6IHckPSB/sCZlFmt8nip5zxzFDRgJ0j4kqd3qhiq7mhG4B1TsHQJhGkoriu0IKrz
bpnKD8Uu4FRHOSvugEwjSjAHmc1O57DMJejv6035NKTqLVcqnWeorEtwARAY3JTv
7Jh8bZIfX2yc5UP9XjqOz9+9dcTfUdKt6SUeUdb2zgazGlXfd+koX1+Sfui5gvv+
6ppuyX6VqdTi1yMFJCWfXvnkNkSTnRDtQ6F7SWY0qxu/o9/qdd/2srwC1gUb8jl2
WDZbQlP+sgjLGIZvXw46KmoKCd/5gLdO+ZsbavTUetO42Lv/Yf2nfQOaL2r5DorD
MnNp1HW3KtPHBVxjvuGr7zBaUi6Cbrr5eoqKtX9aIpSuFbqvOxbBejY0iR73lhc4
zQMNEjbXV7URcqCiKE/bEmp6ts6wosm39Y0MkJUaCEbTVvyPXCVZW2wnkNnR8k+c
IY2Kj6Jqfqv8sJNmcmGhgIpLk9YGlcsVv8yNXa3DDI50DfFZGVo2rYLRffjonfa7
X4CKyE7e3pl+85DWqxxEthwV1JGqrdZ9Yf/ZgGIq6kneC5hOyEZ6/hyCSLxHL+Pj
ax0ivFaTAl+IZOa8zhBh2mOPdE22HZ3Jag0IMJHpoZ01j8SGWVSrfiGDJIB4ig3l
8npdMrwljxnQGHRPHYD1Zg8w3Qcswqx9KuiEnxkY7c0wnLbd0XuPDoFvkJGSkWIh
8RGOEc9jMwmZYMitnEeL/TezUgJ/nrHKqXaihrAF0yEDZUsJSYzHEpdE2IEaICQa
eZgbLFZfeXu65D5Bwp++xzHKqgdP5CnUz6V6eW91hjNNMi47cgoOVQWTw6bGNlRa
N0WLKoL9EOtH8fqXE8BaOHpbAvFV1HPbqm57er8ajfpI0LCh8SYBGswulRJP1P9L
hBiWyIycL8OjzlHTlOFLRiB8jSJxSUlfeWc0UFO0RzuWWHFPp0Drh62dAl7+myEo
Fcka0VcLSI+4/jD99YFjYBlgVWKU46k0AKprekxEih0MEM/vXp1J5l/FPRRA7qVQ
nwhKVnRsbTWRa2UvXqrIZhYIuP2QjCH0h3iYn+OR+ZjxpJgOg3Xocd0J4XTF4RQQ
KhDVpb9u7Zluz7oFMs+yhiZhNR3y3SDDkyVd7k4yjOHCmEtNTncTDB5QPCAYFKLx
jsOr04KCbbz/HhoU6x0JmX6vYx3+UpT+6ehq/8kDpMQKkYhyoQ2ylENf2sY8QMcd
vIREQx8ES4n5lpoYU/LE52dn3+31VA3Z6oMfN2xMvvFK/DOKfzRFLzhz+4M3d4b3
Y9zW9zc6rwcpXLfrAzd6/8KdyXFTWrMaOR16veGxMXjrAE/wc6Zra52RcDlaPd8W
PzR1l2SLYuo0ogxwBHfFsRsrknF4zJl/vEYwT0J1YVWDhL17z19fXQluPqRqE5GP
ZWEyTuSXa4/0bFP/nTNV4Lso3x458hKVtLrmroxQaK166taXHCYcNsNrwOkVDR3Q
LaVlry6KYJDAD4e0A4mygrxTtyyqUunC68+B4lIga2eHdS0nkh49qDEs/AYVx6ey
h3K94rU0/TzCMoHylM5uCRFOr7MYFG1Vpwkkg86TlMTHnHgx4frf9cOoNPggNqPf
yCQIoQROQV+ZQhJa3co6GtB0xjLzGaqiu+vZfxZR1wNWWFQxIsQyyvlGl9LjU33M
cPSzqqVlrAYmWMdPaouyvLoBpZkCzqyTXFbFwBbAWFl0YDYCY7E3mr/F15F+yqvu
PiQragou8CujfcKxRmKcBlfYqA07r75B6NQcR9Jt13m8x1mulKJmE00ViNdR9+ay
bVsoAP344E84F6c98RhWXrI3WQoh3Nk//dO+b774BKo80fG1jLbM0WlVV6FY6hxY
hBD3H8i4VISN5/C16tB4MAccoz/3mIMb8agDCtjEKn6WNWsMp5rqeNxnMEkaAHrD
fDSLC6xv+4chVihWgIcBoyFCLNY2EsfpJ1oYc+xJrY6hKJ19sl0TaenxJ7pErybA
WGkqLPjnijfeg+RhYiZx/HMGUMFsTkYkhl2IYn3i1ioPM5iQB3bkgYlOFCBa4nb4
PCZbq7fZaC7mUG23fRC6L0zM888OIX8mFJtIyCVR9p9l935/0HZCigV/r32lNtjR
RsxqmNtRzdJlFsnw0knuGfIOtcg7r8jmPqjmpB1TylwrtZcM67q/xBuaXy/nLS9t
IjGXGCYcpm81+eqNJvSMzD/sQ+njPQH/C/aQ5uWvFrMquu6aC2ROdXyudQG4jo8o
Qh7S2A1A4cVgcJXPr7MnmL1h86vQE+rOXJN9Z9sdI7t3MTKzgnDu1FjV50BboZ6B
VeLWa0AMm7PwOm/UROlh3HaUwUbaetKCib5CveNUeP9KL1yR0Opkh5mh+028CaUZ
LWeu1ATaChbcpIML20/H3XcjtZNuzWXXDN32K9xGmVCc1XTOGmF+lj7wnnARh3k4
NHdZSGsTeyep3/CkVUEN6eTyTkLRy15T+OJyPgMIUdQU+m4K6NDSHVCSvmHfxGm+
9GD9Jpr5PMmrqTQF5qM7C2jJ/14XPz15TYP4kvtnyi+kf0wqg6YPuMAcK02DE1h3
5oiigfMgAnzCelwvgdMvcUYUlx55Mg9HPopNJ73AmQRycoBvkNj4Y/vIh5bmhv87
lL2qjdP/P7pXJ1vuLQ6X1jj8HK94cL2SM7ZOQCyEOtyVPts9dToZWr+F5h14NwdH
obZRtRq7+usxiFswd8ve41K6uwfxfgN4Rpsz9WKLSVtLxMSq3/RbKwOOgaillKrM
QQrt7ILYOTCOYASuyMPBmwc+VGEas/eNbTpZfyDZdA94T1pMlX3qC/Wrj4JeWfeN
Dpi9Srm8JkIdY903oc4A3fyXyMGm4g1sDChtGxLfu1XJX5dKuEP6sr2BYgv6XWSn
6lF3txL/muhBxuPawBUQ765JHb8h7WJh1U0AVHVOuuvSFhS8BCVW7xHZ5LziQQ3L
KjJsojRpwCK4eqnxBK+K6Ad7BnI6AbkNd7xIyFp5ks37J1KuHrtSb+qPvQmVcWee
ksf/6uIzgqvomq6M1FiZ4luRmN3yZrO3a7W8pNNZ1twqEzHHOaGcNU65WbDH+AHM
GGgluY5uSYwJbHMNV2oa9Xo3oVj62G+TJzNmS/R/R3pS6EHypv3v0+37wdFS30kg
PIaFZnjxTX2t9VbW9xTwbJdy5zjB2erTZuTkGORnX5w95sOn98I8rFuYDYcZq4aS
KEieGuf6nS19722516KQxArgZ0Ad3boumC5q0tDWY6UR4Ys6PVgMiaTvpZLI83Hk
yCX2VVeobDIgryq37xh7/mch63+XtK9o7EhR5r9WdnPL3v8ps4q3Bs8ccPiB0GrB
9bGvbIBXWeD5mE9JGt8SG+ZxlOYnQT+/s7hrWFxjXp2TNxgN6V9meKGmJlSs0zzd
A0Ttz/j/rP6rl1au4+7Vqjps6Dgs2vM/pqIhyyNDbJey080HRCRBXHUvaGIhP6U3
IyRBxx8ueYLeD5J90Ij+2kB89C+Rbc2tUdMrd67tDpgD2cMgT3uarOJAQop8ezVZ
1fimnrLP61/8BhMBj4fu+Djo44zDIt1Pf4pVHqY/b9ympYPLQVRkJRdexwBH4zuC
fIgeTZzjqMVIeHVpcfIx4yYtrE2c3AL6dnpRU+WVMTq9mpBYQU0sEui60EuuPgS7
HZGNTvVH4m0k/tBakiCxKMNTvaHh+OspNXPzrBlv4k2Owm6PqGcA91Ko+UcF/wBH
M1xy/BZsJhIwdJNBcRGCgJbF38XPol+y5I4F+t8XLB8lOfFaJtEyxIl+l1XZW4VE
1VyT6R8hQXtye5ZqEHxjm24Eb1W1JlbuNAMGIAufG7rK4UrPHmJxF98011SiQBH3
6r4v05ZJJn4BDGk76ru+zReE/o5fMGX3Z/XdoOJdvfiyDwBT/Wws6titUaetEArm
B521Mqa5u5pX/JWjecHnefB1zHZiX2hpEShf8sFOkM7TZg/sLD3jiHAwdMkBaZ8L
W37XBuAysj3kPv97n+JWDVJUTAggHznf+tI+9O+90wR2/5XQQxqRSufP3P+5SCAE
kQtP42sKHZjt52JI8ipcEuSy5SF/yV5Ru9ciKp1cKd83PW/rJFkcFSgi0RckHr1i
UEkVV3MXe863a7RKAOQ7xM5go5uEbBt38yXIU7khsP2bAW6yiX5lReKVVo40Yi9F
bN9CGMIa1KdsNzzqy5dXrZqYtPm3rS6oXrCsRLG7njHlsFREYKa0CFuM0wXw90Pl
jaoBxYiMHBGvI9f3e4kt+Vbe4oaynUUdOE28sCBSBCZqlKarRt9dn7Bz+P3xcL9U
uCGQDlo85bUzpf47+Scbv3sbqbstdrtDCmwvMydmUNEI/G8Wy2qCF4p0iAt6xbIU
+DbP5mwAEp/K3KUJc36J6UGzDS37Da31vFGw6Gs0sTnS0jT6xLKOKxY4iovRdvyv
l2y/3+FPOq0GxzouCbDQ2g6cXfKFVNxSvvEvJqBrtMGLejMMcczDzVR5eHWZV6+F
1VACWw1tJeXKVuPztQmmHf+J+me8NE3pPXLeomRJ6MMveK1jWetO1jds2eH60kg9
2jl5Kln/5V1zcnINuuM/zC73hVjIswatnhxZIbqJZOkjWDt4R0vr86qWSBaYLQVT
/DkxD8DN9rA3tNLFWwB5k+LLk4A1ciWYcqUW3AyhlULHatMiaAwruoCWjPZlCm1N
K9SD2BTtM/poleOeY9BfZPmA8jyla6LIH2gbP3KCH/N7SBOOKg1eSk+ZDuXPPkJJ
cm9mwzsMbN21CP5JClQBVho6qu0qYGPE3Z2Wq/IscrSUmHBcfQb9017CgAWFWQNR
9bEAsaMvbAEdX/xx2GPx4+B24w6h+rtpMNFSPBjJN8PjoV86epecOjekZFab24U7
rZG9Thb2asybMfxGc+5JK9BgJ+KR3/HrH331xfY4w/nUCT51UqWTW/QpQrbgbN3S
+5LTAMjQYNohYKJ7D/7n8pNGd25FqliDW5andtRo+1KPp3zRAgOYh+CRvALiDiHU
utcBTJ90OzuRCAbXrDNP5Pm/kJ9rxAc3eCNyroYw87NIc4zPKNykWdQxmgf3xq9f
Cay71heff4UAAEBOsWno0ZR1+z7QmtlBISPRPCU5TUWQN38NjnD7votySdpK38oq
HkZAJJernmEtLZoPo1JTgHZBOnsh7qO3FphHH/42+PxfqUJC+3PzF/izbDtG6CJb
2AVOJVAPH+KN9wuIseoAmGy127RBZcbl9zPVCbODoZegTvlWzmLpUZqlt6pOXHx1
aVkuwU2s4LVOVqKErRZamCs0GPzoCmwQwyBsYOUTPOVd1bKSpMlvEFZBeP2vp8gN
84DNgEWnyCbq5eh8Q7Vxti6pX66dVXgrpP7jCyWIRJ67d2U9IgbhwijooS4ZHRxb
VWp5mBqdXfgcCcKpTnIQC3ULoJKYEvrzmZoCM+oZzZHcpoc/0p9SGKsXGVtZlpEv
R0l5kFZMJXMokaW7f+1KR5i3yOm2wukrtM7gFnlXIoi58fHLmiH2qj+n6FaGeqgW
gPJ7HjoW+WpN/YE/zsytKtrF1aSpDYJctEbVq/+oRMLQQgMKF2OeCRqX8HDE8xDI
0qkP+MByUBzvKoY2yw4Dq2ZZ3RL2ELxOF+phGuYg17e7Jh1d0DcO2NvdNIxCTyJJ
ZJ/cbQC0rqfMLWTFbPS+DYytSbUIwVKVLT8k1aWNMfE0G7KY6RK0huWAsPcHpZpn
7GK8ntEcz+FfVqw23Zgb8nw6wAN629ms9S93iUP95qtMDpuTGlMaZIn9nKRCf57r
i0oxqzy5mKajXkOLZA8r6qDXsEveR2HSZ/NC4RtmkxFHM+USPQ/n+l9vINclfCfr
T3ZSFXRZmQ3dpYbKT66VYga77i5t1g2aVE+ko0FeYFQ30jK65UugZJWJ2r+0K8WT
jLApucUQ4ktWOm7f+4WqBGYEuCUYCRs/vyCASZORrLBbNTaftF3OTZXyTXyNZi2e
7FzGE/WiYFDWR8BwWNXoJsEI+GGx+5R/5L4nnM+V/fC0+M5C+tRqFz7WnxaDKAX4
yaS86runnTB1BxgzJw81vLF6CbscRFPx/Q/yLNo7otkBbQ408dqDI2MPFQ1h7YiF
ddEWbjlmRLB47QFyI+dL8XmJSdKVbSBmo9+svqHQI8cgtPQT0bPy5P85ed/3sZ6C
KZ9Ps7xAaEv4UuspTzsH4uQ9kgX1UCeISMSqjqPRsgUUVEX1Ut9oQnIrVxvtRbNz
A6cxXZXMwF3jYE8fD9UeK/SVupTdko/7scr4XTS+uCJVJinRNCbp+G59KIiol55y
G7hqfl/LKp2DSU4QjTDnEn8Ix4Z52CpOInwlRMg/Cb9K4INgYMGrgI5OJKo16kH5
RKeqYCtKmeKVJjXrTkCjiZ/Q4gwFOL6BP7Vp0nn+3yylYLPDUqUNaz0XICDyUeLF
skvHcoKlVeDI2SB8Er4ALcP56pF9Dw/sBYB80cM3v70D5Ttjm36hXS6zLe4/NuVc
oQP2/Capqkgn4R+9Xq9gPjSg2n65U3jKPNBPLUqrBPi2wKueDDIdzXVGihnDWIT+
3xSKW60QfGj2dqEBzm8lNSsSONFZfKj7bZ9W3YYtEQgqP5qRtzvfOkC77OJlGo0P
zpTGFi0akUM7aDHF78DWBja0r+QnPZnBnhdkQzdWVEDVE0lTZUsBiqT1tQyzADbC
ADCIAziESZmf77urrJtIO68LVViH5vhiMY1ob8LuZ7fwzU27bmV5/kssxnBwbGRz
SuU9df+C3hQVttgxILLcGb8LvH9BrtyVvCjhPveBKmzdhJ+MUgA6zWwFtWPHxDBJ
gfC0ry5K3a33USU4XSffYJJK2C/s8TCjN4oICrtTWTupfOU4aoYpK46bdeyvtK0q
PJs95K3W7d9w2cuhTPofncsiUZBZtBcGVBSfE549YZ5ARIHWEnSh7JxuBUcEP80e
PMt1CjTPMAeJbsGIJK4YkEXQszoZy1H9WNcRwMGS/eRufNJFMSG5ew/T91HHTdwd
gougRlWT8nvK7yvtnGFH/klRiJjsNdWNpZtl1uha7vLt8CTxXgzGikzNoatTXcwu
ETHDla+kZO5QTXqt7crixWNALVD5QIXgMte/rfry2Ht1ZZSum2KT9dO5BZWTSK8/
wnLx2buxY1ASIBllzP+9UIMbh+gryNZQLi1cLPDS5soRo2/2ogGHYmCDhytHrbj6
WLLNJ54KA3h2Pk9xhlpVR+9E6VB3F7fjHP26P9d5qLWVMRa4Q/lWaniiWp6r1suo
yIUuDxszeMqEZTSMDJ9+TQUIwXxEweE4eK7hnQ3xRY2HGFxi64y5I08iDmf/ENfG
mJEcnqLvi2zc377FdrVi55wN0M+OJugYKe//wbqKf+BhTId98YIaS3lXxv/D89rA
xj2u9n/Jk+oUASfKStZx2EUqQiLEGxblT+NBdZrCmLQMUnUfiCGU9ZcJFbrxiEhX
qJ3X2KUAyRWXakidfG2ZyZl7q+osfFkORg/u2vsWGVcZK7HsxjTumc8gUTkEP9MS
wR5vcF8MXpbYyF64G4Fpx5vXZgkVa92gf3+t95tZZiIpvN9sw5Pkei2ATdcWwT6e
w+sWCI/5iWgrA/GfVin1kWoTVP/iOJ4d3vKHhhcBBg2Yj+vDG6bSDcw1G4dHK43/
hUXALATwaiUWnBVLXgD6lKA2tb4BnuAgyDW/MmahsJOC2bHHbW5v32lpMYwwiOI+
zyeZw9Qv7OB8gc8rDiqb0/NyxKQZE8bjOHQAPFl9f8Z43q6SzhXwvPFbSL8i0xdc
+S4Mm5FOPbUfBfz66tc4lDQH+hAfLMaqT2xgiQCCdezMow10z5i31/IBcEJ4cvb+
HXPrUuc0mH7rUacw3vF+NVE4qgHz17fRcdMs1ydZvJ4/KY4Y/1ir139VpSl8FJlu
xbHt3YMQIGL7FH4/oIWnAwjqMh2GLzL9GE8ylqtYLk+9vex2MRcoEGMfJljCWqq+
9Ya1g2wbIzK4WrkgWPnt+aGS+VqyJ9f/ZdDjWXPAbHHyIIxAuBRpFMc3LoaGaaUm
n6lxKu+HDX/vrjM39eLy42lKmwkdX2vXBIAFEldfIIZY3Tof/XuCENPSNJOqTc04
RB68+LoXuqyqlQl6kT46YRcdh8/34vI5AdCQucJRt8bGLFNlhpTW9FsqRgbC9eVt
e7FKEBrKrjfYBCr/ytT03f1GRX8L2FPdDfKnFR0n+OiNY3JNusqLowIkMi9lq+mg
TO/x+h0lJ5r+Vtc9YIzzMag2K/U/Z16M5p9H6VM/W/vXfWYIg0fszFmY2QWIc4Ff
2P6/2WVG1ovh18b8rIgN8jkLtl8VNqz8z6V6FuLdznhl0O5zvkiZobxOYEkVBr0q
QGZYWnGGWegM5w4dPptbkBtbYwiBnPBhOs3oa+Q6qaLuCcDurviqMy0XQx0tFyk+
d0EqIh1H10Uy5LjPO51XSXqYKSMCGOr6+wx24l8uKaWxivPshLPvv6YVrv1eGxuF
+32wcDtPjEPx1IL8+Pbh/Gm0brHLcIXHWEXuZ8dN6BZ4qTC81L8FOMLTnG5gLD1C
O3hZbppJVyP7I/hsXDpJnL4yUDCYMbVj1Q9JwiQxL8+yJkPCXSI6eoQu98Zz6u4v
Aomy+rtIK/yUdOWVq3Fz63XzeQZrzGGEJ37oO/nZmMWZ1jEtqKowfHX43kP91rci
lBF5TBFg0c2JDJ1JNJw2QjYkhvyIs+uQrQ95MFmfu4EpI8HgFLcnxidh1mzeaC5B
b1RXI13X6Au70xsETBsAhBKAzjS40Tp6B1NAKLquQXQ/130HH9npnKneQcZSGrIY
uyOqDKYF+3jXf+RFLedOkW/7aVSb5H4H6Wy5GDY9CuVZMcuWMq054WwNC/8oWuuf
PORQazxQTeHBvauyIVUW+a/4C+vor5QJ/ZkcRx0qQFhMSlPx10E5krDSya87j9IX
gyRtf+LgpIYAe7Opuki+ZV3hc7RSlUFAxr2Ctsk9moO+WE5qGFkTa3MxHSx+ubZ/
cwoFVVIiUzAOc8WlWOfrOfWhL+pqWQIJxpLYb7zxDmXLQbAAwILXAoeGyh2FG/3N
J8Zg2rnJcA3ZQ6jD4wz+ycdooCk7aDRD5ENG4Mg/o2tl12YZnl6ASFUzmaZLqPwe
OgsY5prmLNS4Rp1FGQtUeQUYnSRHck/BocMpN3h8ghXPwX29R8DrordWkUydf/Zm
HxbVJQ7qYp4iIK05c6SwAln6Gjlcq9jRCgD2Tc5o7VusQOULWTmsi6uik0kzQcIk
9/8owj40hnOGbWCTq7UN2gKazDGhN9OBQslrR/L37FTkQlyweFs0NFGjwlxg3Q05
k1uvi+F093QToPfN2HnwVmvBwRJf7isi9FghVLeq3pjegGRM8wWMNThQy1HGbOxQ
hPztWED2kR0EtnO2icItpiBqzN8nY+ITHv8eNyqZOGIbM0vJ5Fol0Ae6tm0IBbh3
mFw9yzGWRXkUbaNSLyICsPRnhuYJ+Uv/enTyd4lAm0D5EiRRpFDY4jRLJu5vX9XV
JIkxNzqhg7giqtSQAjfMaD2dt6dzHNIzusDHwhXrUGXl4MHgKTM6ZxDugODl4ytq
UmrXOAnfynwJcStdoem5env+o9+Xbfp4w/Nc+QsMh2fnVD81G09RSHcY7Xh8PBhp
N+oVsFgG6F+2CxTHdsnfAsA0pFPeOD6c8g7/vZ6CYk3ofpA4jkjweDJVK9aRW8G7
bDrJkN1LH2uvlqHw8Po/AYCagptJOZ091lJDAV+y7dq5hiaiWy7Qfdu2DXCFrQml
lqBnA9EfxkLEkF3ghWN9JM2TOPbiigrsx8piizcK+4Le/xQm3iep5q0b25xefOnd
aJEL1FXUHfPGA9LNd8OJ8GLJe114tF6Jv8DtNe1jI3nZFyhdibMD6lV/IC2Oao7h
s72kPguJ2QHO1zg+3Y90XIUQeuMiu/zl1X/WBzJmzYUGdC3T3WC0VKGxvpDCr6BC
HTCfffbEZP9YAJLmC7R74akxWKXQ3yUQ3dRgnyXdjvVRk3dNLCyGcIe6XXhQ1Aqp
pJXyz5VqhzzaphyPoVsX1sseOlE72cMzk5IE+kzN4LqC/te8/0DJMisICCtNGKAn
9r81Dw2EfBShqSmmU+NvHXyTuSXBnoLWaL6TIk2KsUO7ikMINGQI/K8O9AfSREvi
wStZNnnQT8Bs/eNx9TxP2xfqmPMKdlrK8tJNPRaUNmuT2P/vHuyeNMlJTQZTrFJI
EdmPD0p/2hqw+eGRv9FNsOu7eSefh51LSzLGoi5xDH57Pxa+t56w46JltUxpfXGn
tQpMdbBakBAvv3O1GGvtCOTfAH2fO515PfCnpjNu6SHftiGC0MIZ9+ZeenGOEvcK
XHC2Yyb28c1YNfrik1ztzk2fHl4weKLpImfcUPUbUgqUxLnmVECfsqOSrkrpjodN
pS+oLFniMRtKO+cVbq7/IYKoqkZk1YmbeiEWqWYWo9gASsbY0ymVsJDWxA62Ny2d
UHip+MVHLGDRMiZOdopW9ug6q+WHJxZ6IRHSJQn0tDiB/s1qd7R/Cy8fgCQ3aAP7
kkDPcnGidDx4t1Qy1I3hAPMS6qlNkHBHzahbkFdzCG5qnsshcvWDhP9gNeP2yEiM
MItiMY1/bQpSMVq/51VXPZpljbe5yhvZ51oDe5GVLY3BqdXE1Xggbj/Dz3MhCdhO
qIeh2QPMJAj7sl6l5CQhQoZlygIB/8auyMXvwuX6hpZ5OTGqDoT4pacIp0BzkgW5
9v5fGLkxgsZC/DBm9FVCuz/J2EFaqn9KAynB6zNzNQymS0ZGzPWmwFBKddD3o6Hk
iPtO58dUnNPvjnSI2wGctGOthcogDShVvPR3t6vqx06f34zFyimLW7RoyVreriGt
CkEyKgKA/0Y7wH8zVA1YfUWtLS6LILLrMHYP9QrH4K9wLUtDdoa/45TCUDDukuhI
uj/ZGbLs1xY+5ciYx6K/ftiDtiOkcQ+tlHalGb89sIu645rJSOCcaGUTsERj6TI6
ygIQ98/9tZ8Qjwr1dxaQoySLKWIaFEblTF6tH822n/8Mmn+qt7l62GMXH0V3V8Vc
xifMh2vnh03E/nboU7BMQiHyo41aNU+YORZF2wHE2/r6V36d0sRkA9hptJ5Dzq1R
lAaTofYLIs5JTs+i/eIhZRRmCU0BUVDzUn3a7Z2nR2s1glOi1G0FlIJrGr271WX1
vN25kRUl/9d8AdZxazGiK97tPFbxfGSlNYXdjAMAGrh4udoLpqCxeF6HWWOlPRgS
WJrrtRqWeMGBGeADvaFw65sFxCQC0k5uW9cZUJvK3zEalfD8dM1bi/RDD9/wu97F
5271HTSrqwT7l2xSpoC7AOLJCyCc3gPxDRrAv+jpt688kyqaIh/3DBLNYodElAuv
VAptttUZCSyLSD4yiAuDz1RfJJZBCj4cZupME7GG8dw54NVME8RCiuFmMRsePlk9
uQSs0tW6aHatv2abqlaldfaFZfE+VS2E1rcGp8KuSSpI5xsC5ZJe6qf0wFZP6ocE
joWcwRn+wt2riAmpR+TRlLKkivmENHqD5NcBx7uytt6YztO5fj2qOLnmyiVo5P1T
N81d16xkguRZOalrP/5SdjWUb6W8Up4NzIiyUF93OfJV+l9AbUisL6aFZPh1DmSg
9HlzEHU9AQsjntpTqYLb4TJxnhXq99Sy7FXGbsrco7sdonP3M6lNNit5nvE/eh/J
tsyBBqvhNSl2B7cg/WGsOmdTdQn8ZzXpt3+GoLaNOajJl1brnxjUTwYz4ZCmXLiU
70+N2bqhL2WcqNyUCbQUhFd0t4MM9fHW//bm7Nk5JAe4Oraa5hzqDG3R8wO0O9Va
6x8csF+m+4vlSES9PtF4ifqJbVIuLZZjSSlyj039IsDwQJD6mIst4oG9ciJfg4JD
J23EcWsbTaVOKOFL3f/tdwL27Yyq64Bn73cwLDtZkfUvJMyUFcqNKb6pu4DE3mcA
8OO5Z8eOF0fi4t32NRuxdq1zpZZV5gcLEk4IB+RuXVNuz85KZ9zriP4lXQsywinc
GKhOaTJIPvnD5MzWUKuzqTsZfXdIhRjULfUr6D78TfpD0lhBbKy2C+iE223hM/G4
2TRz/ZoRiq8kydeTcqwUb33wnRea/3aW11GYV3yQgt1OrxLLE78wCGIJ5RIIqVSj
ehDvczyjFCSoEcgkUoXYO0fzQBveNNYDws1KXOU3Oq8VtC9zUVy/+quMi/Krwn3i
xSzrDjrOca1lopmEFX33/gJafJO8U5H4ByzMpNi6Z7kVofpPuVJu8+9XEGV+x2Tx
3KkmAZ8geoj9lLIFBQVzG7f1x42Y3liU2UdFbCO5nD0QkYlb3z5/C6mgsgWa3wmw
etOgMghWuxQ9u0dhUoNYtwO+xIWejDiD5QczmbHPjz0BzN1rjROk7q+y6L4L7xol
MUb9jBdAZpyU+sCRA6MlxgbzKRBh4ibEqfh4Tpm2xvIWhljQ3iLAU1zlmK0Et4eh
FOuH8VUkRP/czHl/lb7FxNSKyDE1DiTEoJzMZmV0VKaq/rcNwZibnc35jqBds7ud
5nLnKYPjUmOds8Z6S7sdK7Ia+2hCnq4WZ9YDOtHiKt1rMKa1t5P0gfxxqEKkFwBl
kvUhMmhghC7zkacFHDZxFoFZ33krTaVCKoJPOXEqyyLslyVwy5FBxK0a+b6fFHVB
WN7PAiao0XKynO9OgcZ/Iy6HGS5okr0hpSRLBoL/2ga74vNukA6UnECeRDnuSFdS
Hb8Ezc+Vyz0folAX1tDaa2BJkl1W+QsYqRTmBSeLyoUKzZni+eMeICBKYuhYLX71
xckJc6Z6oGWdyGvAKYTk0Y10C5odX3FEgeMPCuoMD+O3zAZEraKkJQ8YIolMeM5q
9uMHGcJb+gjIhxCijRSbUya/NgBaOV9yA/r5qSvr74xwlKy3bFJAs11R6mLtkceY
roJX4T1iHgx7AgaUfv7DUGrQyTGHOmZjgl4JAoUA8PJuq3NqIiIWmz7b++7xYuGq
E/ncldKM1+Ntf0DdQiQwmmOvaeFD7WT3bNyhx4CHVlhEbV63eCbSX9IDjGV43cSY
4eJSdZ4UqY0SP2DmROz0Ci/QnKyu0Y+LSfWe+NZ+hdySt6xab1RpjpV3j4LKaakn
yuqZAlD+kjjO3IUAV6/o2C/z9G5K02dGY2vMSveby1EjJHQpIaskfnqDn/fQK5s8
SpQINgXDkP0em1AEgjRAdnqnhEpVq+QaBNw5+ia9BRTvLShP1AVdhy2v5sN8lRti
Dn5C/w0wtv2RA3IqNrGR3YARFTeXQufBklwSqidvP38aIlKJ2adGZcrzfcnl9tHK
f103fYIOLws5GtOZREreAjg15Nf5hLZTYrXHGWRmjQdym/dkEY3bso7McG1iBHfo
ctOXXeh7AjacC/hX4Wkj+RwqdL8P2+xmVe6vWM1uj8jiLVcmuQt8Gg2mCE2csFsU
O7S+bqOdAW8Zy0VFnWMYi4IJyeQgTArYTBoQ6bSCQqzQ5hdhsaT4BNFp8IwVSQ6w
C69FikxPMdb8kqKoZ5Lw3YszkNtriHjM2nN9tf9KlKsnDgJmyOHJu2OMhVvmegwU
sts8m8IgC+UPmoMlpulDLLI4UyNswFmQZmsHZWnzyCejpkNP/2PY4+nnjweylOml
pAyOVdLx4qN0xUdJfpU9n1fNbfR3ebHX2xNcr3JKASj2ArIzrWj0XR7VGp15ai9I
meDmCX8eIz/PeDS+oB/krTdPz5zHhT1fWdnSJZ+BfMv68IMTp0a9Ic6OxUc4fXUv
zECUdrw2DXssiFa47VLEM7sH2JzP4+3NOVzxICVczzfaBIfP5Dlh6iV5uGWfOcV0
tGeWE2kMGC9wfBuYZ+k8wtmgJHLAuU664FOUWmubWQcJyZ0wtuyF3urYSFuce96i
nvVodhno1qE6d92Tys+l4cxuxYbVwwZf46sPM+ijvXkx/FNlSOnCAvG3Js7yndfd
2p1/3d7aEedKSYQULPSlXrSt8jweB8QjqBKJxJFh/ue0L1gFNLEGa/Zcw5ui0tgK
gQ+9u0MbS/ylcPXfwqTcUkOAlKKOu/ybnJMSRWdiGb7FmWEahMCTIdJxjFXmWKhV
KKpAt3lsNX1SFn8nqmS1h6+81cpEZn69G4gxzfTubZQONX30tCdfqIIeOoUY92IV
1gCTTqWTuDUjZ2YL+k6ZIVF+JTXS5JxolD+JASeGk+imxRInnqrQjKpP52lMkixO
UQkB0+OCLrGg/AAZcDYzdGFYgs1vzKDG913HrUNBujNiPOQflXOZsIaN5V6GYOR5
abvEv9NTg1RyvYnXPqZTgJBJtPdvWfWyMPi0XkW2ekWCtnMPoElnKtjnRhteykZl
8wQV1XHlNSrmOiclpT0pAWc9uDbgL8jDwygaLcMBPmTGNR/C7taKFBInNbf5D361
j1UpbfhsOErsUMzgx9qpi4PBvbytV4GBkKP7DDUN21IZTX3lS96ocJ7Beu8FjaGF
MatGYmjU1wGAwnaX8Kmqg/OoS328aD9Z4M9jOaNHjLzoBhDOH97DYyfniwiJ0yWu
TJ9Vf3+YODgJkJt43qjeb4iPl0uEsDlkVpi3L5MC20W3GlAWo9muUUHGRN9OtNmY
FtQSs8JmW0jFmOAjySmh473nADcK1cP/PdqfNQTLYEPd5C2DW/clexmATbTexYaL
xoFeL0A1YJey9ihoUEsB/qVKBRXav6dclCFzzJW+rik4/3EOvNRTqrWb4p0ly5JH
+Tmt/R1+6rTjp2Ax09XI3TntBawn6k973fvHRh9hUrRDkNn4fr+4uiQnv130qceq
CenmnI7t9wKzBFmrXseLIFaEP43BwSigZlQaEoC1nqUrgGEKNuZawkTJ3jR8uuiV
s1vscpccOmuyTx/1VLw4xiOJ+Teh6ZdDXtzGTG7glwvTFVWvn093sSLGYB3x33m5
qzzGllFjr/IIAYsG5T8rbCe1W4uWJLoZu44eVx9gq8Ij2+KYIeLLz4KAGCY0CDbT
T4u3i2s7uCqMZrlpkLGENDHWckAX8AHvlahS4OUOKPWph5qN6Hv/Zu5ScNFNzWr1
/VdOYhLVgljAIgFcAbMx0dMiQ4+Z6CeUPi3wer0lRGJLybcyckJXPJSeWljsm1cL
+HXufwUYGGePGLwKq2U46r+zuamorZGBiMEGwC3dU6HQzm2uEEyQbTnYGy4+llEA
SKSSm3wkISQR+5BfrabTEYiJp8eijK5dWb6fa9eBjpnsdlw4J2A1m5tzgkXlrBRp
ug8mLcNzbAocHH7yKoHT1hZjFOQjzg/djFBFa8nyDDHVelQX07FkuPVefRPlSb+w
WzCjHzSK2FHURqg+T0w2QrVZjRJuACaf/n9tCAtoGqPPvHU0Rur6RyNcQMCUZLmU
N47oMtd1BtZfzPrBvJg7EUd0luxY4ElDorb2UkgAjDarLHQOiUDOu6DS3Cncj9ox
mhVpzQyb0SelefMvfnOrouAQw1DqPydIINTtyHp/OZGzt+ESA8BqPXWqEX/Mt6ef
mjy+nanFmqgbNDR8026cy81rlEtdgqUmcODtBlccVRWSIc8QmdmPtLjB3Tz0gMdD
jqdwrqP1V6y83DvV/13in64a2krpGiuME6Mo3ScOFLyhlF11X1jV8cL8pSeZIXEY
wAFmJpuZNDXh59pmDY6KVj8p3OyO+plmsaP4MpkH4cN6/tz5EUEBSdpBLdKUAhQx
mQa4wHrvM18odPOe7NCIDYLV7x3FiMnUrBIPi1uFnCj/IewD6qCvyuvl3YNNcT0b
aG80dFYCDprgFdZqHKpHPy9v72btdCP3RF5CqUxJhsXjcLhv+YrjOrT1WYgczh+C
LSa4DvugKz9dxFAbf+EuBevWnQmtfp0OdFmngdqqJtaGqRViD1GnroWfGdfHdbs1
To91zDSkXxdJfdCSzwbDEq7+7XPiCxsb491fbuqK/YpGiqPkrrM7Z+fefHpzQd8E
dsNXO4mhS1DQxID69/HvTO/zGLVCfMGiRfQchnBD4q+an3pbibveJ8VO7HyboGyU
6xa61QKV42F5uL7DWAu8W+suLyKicd2J7N7mV8QqdgtB6wQnHbZGWxqacL7vtcSz
r0g/miDl2vCtQ/xs5m1RE34pFpV9wxWuTnBJO99slFWtvVaUBAIzJ6Tkz0kBYIU2
kOlFMFD0m45o2SC7cgJ9tkMwSTWCFQ6J8eSO66uz2sZYAAFVkeu4sM/n18v1oYs6
krgXw/KTLt+v6DwNVp8J5E4XbBhk/DnC6dIqcvneb+aQgdj9MXhugefG+1wiPo+2
c5Ooi2nlQoqUZFRQhv3LmAj9hW5EJiLXCFYtK19rCIXTQrfcbLNojo3QaDBvvsZL
BSQEeeFcb5Zwxx6RgRewVrV0TmCyHm8BdTfUXB/gu+3ViaJCYnqX8A8o+7m5HTLL
s7x1gEO/5zlH2uq3xx9klmjnk0PNY1ZEXA3fZut6YRw6B0UhfIyE1LCCM7HCTPYG
9qYrPnNOdG4qD11tLMERR6OCAd1G8G9tWcAdu/YhkCsUTxab0h2bao7azCBWaGWo
oAegwOgwX/9egk3KHovo5y09Y4PMBo8rh/omqnPO8MyoNaL19qjVbVS28/BUiHqH
M7GLxEg2efX/pRYudehBv8c4azHz+TTrE8iNiZHwC2S2s+dySIoPfOLD1pr3Wq3L
OXKd0+94sWTPGNTJ20Bq9j3turoI2C3jskLfgq9f0Wf/ulfRlayvP9LULjhVDjoy
UJ9/o1ia4BeLtMB+WCPvxWNBRv1/gRoYb1rDAudYw63iKP3Ih9O9R7+5Vr4K6m56
qkf4g3NwEse9gWzIqsivl35iLBlpM6Oks1iusmEQezl9rcoTSiQvNrSHBSWOGOXU
BIwFYhsLYfgi+z4zBZwzsrcnNB0SMoctRy7gN+yu4XYkx5my0+e9Hg4BadCTCpi7
LuLqi/kVk2kttdf93ukb39iFWHXuLC1kOzao5RAgrQ4rR891IYqP/9aqp5exxLR5
c2ypdCU5ac34TkCUi/MoSsaelZK6vNtbU93C8CeQPSFTXWzelHWdWq09nFc2oQTF
2Avk0uwXOqam5ZeQDjhXvheNawMMkEaZv5ZRADHgjIZcaWj+4PqF16oh9zmTIGMc
OBk/t3LgO5i4+Z5DkA+htHr1iQGvLqfRSrb5j2fKDqBXs8uNwZxA7lKfEtVcZv9Q
o9ZryDuDLyD5nb6tjJ7pghqDV9t8iLJBYw+Ev2kfcdeQd7YLVgT8Ig2dLODiK8Cb
Ly+4eoQ1eMj4Xf0rTnWDbaIWCbiI5bO2vQybEz7XOKDYMGscZauVuMnYYqJFkyyU
5ZA1K1rySsgIQuWNCJNUM8JsFl0h0wcc81WnVU3DwFQQeWAomod/XzjweNhoUMsR
11cRFJTUHU+TuW2sYsyRIWRffb66cBTQdP4qRK53f5pjM+4CuLyx7KMDWD5xgvVK
GW6wiZqN6UONAYo5YHVab2kw7H3DGcoBy9bVDqxNUJ9/gHu45wj1OR5s1N7eTqir
V2HHRRgz4DWDXctLOKTPsshike86B6ONfOmEaPBwQi0Ty4vXEYLk0NQsVLdHGTxV
te4ZQVvPtppaLMsK6a+ixbyLsnmkvAxcoiTEexho8i4eBvOQ6frJU2VLCTPu2cQ/
AEvpDbJ/V0OmYReNkomt3U3DhUsnSMKEx/5QyfjHoqt0mO5Ibo71cG9caQr3+a/L
eRQwV9C9dJs4j6SN/YbR2ljM1RL51x2L7W8W95/4zDwANxxLeN6sOZMp7W98gOAG
LaQq6EtxK6+Eq3HBCMB5hyeh/325a/XiLwAphcDmKGuEQsxSd9mqkUpoEBbDKiMh
FGSdGyqJhD3AsW1PYy56HIIKPGbd4mH7duv5sMEtKmm/kxPl11YMS5Nc3aQjfv2z
YqO/llbvAGOAcg4EquGLgzib8X5UA9GSvQisZcWVyf2/R0rBzCxnYdunCizWuMfa
QomxFDJW5K4airLJYvYfrKiJgMZV7iQO92WoCVGZkALG2NbM1lpsZp1LXIDk9rKi
MMEQYFRjkoY9qvMfTWXZVIW9caiK/4L+7bpdotgO/vVMGxxjlR4U1xQmOUCTmqaf
2hrPz5KSOT7lvvzB3b8Kjmnv9wv8u8ujARP+spZ1TfT+Pbqya+PEb4ZNrmmJILga
T4AOUgyRhItrRSvGg3KxSeXCRGspZb1VKQNqXAUgfCJHcOdNyVjAHLPbecjmE/xe
YidArQiNVWyb41BdBOmLNjP07xu6JlTWTUjoRlkMlT3qWzNHQ8ql0e3aZTU5NLF7
DQw7EWc7rFdEKhhWxU35mdCKWg4/RSny6Q0mgTuf8Gh7LVlwZzu5GmB/ZCshJv43
s7TV/P0ycLWTfDMhOyRgB/w55yAtYuRECIEYXSdNjdzMj8kpQalclpQx/VZkCpCj
vdiWerugO7x+AD4FkK0TsTcV5NI2MHHzJS37uY3Nq0uefesWJYQAQ+fdDfImGEMx
+UKkL3/QPe+NKZwNI4tvPnFCKjPTVC25hpCCYz2PJ8rtTkH6mlvjz5foowdwLw/S
p0ZjfNf7SQi1w5SW2HIEkeuurDK+sYqrBdc0MrlJevfYxu4t4n0EievT7q3u6ILA
7deSJwM1QmLTDH+OtBaDCaIetXQDlYitGMTHKyBI7ekZfa8jxRiSukwCbkmT0mMh
saj0+yRHVKPuTg/Ciw9ghgSDuCfimEEB9QKWtJ5d5J3VBi1y/EMifqnvfZblv4xk
Yd949jyNJbko+wbIKC9TONYdlMhT2uuzd3PQep78qWXHu8H/NINVS6fY9me4aISx
a4SSWqO5pDW984ai2xHnBNmqbcOX2e00s4M2LaAdBD8ubJdRLAUAG4fQTIRa70AT
fr9gpG/kWrYgUr8BDdz178YULSxFoR0diwe/ayfYEg/9gBJcrEZFOUFoVSCdD223
GqT2f+NHRtgM/k1TESi4Ch+xYLsCrRtjP5DgJ4Q2sfbUsHH82Vv2j0ouWz6/Uxy3
151a3xeKyG4w4OTyZFncJJ5qGFv09bUYx0QlICp91L2sWUNtlZyd8pqL9s22TGZW
PDjK7Q7jIiRAC4nnShBUDkYRcRU21y6RxZMu9CMJjcWkwYjdGmhCyLgmh2AsALOy
/glT35qx5PNGKQ/iUMdbrk/f/DZzAKE3laSi3F17wr8YWZ55WpjPqRVWlwFM9PuE
9Urugtdue9a+KIeiucMBG2IY3Z1IdRWVfXeLDCWVA9P3WXTjNas3NsCZ8QKNnfvf
tAM3c0DoUkqtq0sXB3m/SUlRaoq/PlNc9ZfWnhwEh0QvMyRM1gF1GjljxmJ1hUch
kRazMqsLA8c/9W5v7HFKMsi7jZwtXq22pQZKgQIIFWvy08nAEnCU62gl9WEmtiDl
r+NvQryohS8RHNyXPcADBn9EG1Nkc5QzzoInJS+7QM1aoQuXkMrj9D4d7paj4QIC
BUdcfREbe/eetihsN69bvaelYZ+QhXvLcVh/kzsC7lggsU6PbaYN3/vHZ01MFAc5
bIroY+B8zWoI1SYlK9wcp7C2uEzCTkWamTMBSQ1aofxS3HXak4BVdQ2IoCyyEH2Z
AwcakmBYRBMtBI3kppqg/r4aZzyN+A5PyneRIXD4aGljCi9nUczcGqtsFnPdcSta
GeqbCZZu96epICXoUmT1K5F6Sa53gBK1T1LLbKmK41i5eSWIJM782Z8hUmd6WOsQ
8uz6T9IXjPx9ub7chHO3kSlDA+eNc7sZOJVG7WYwI8mybUfbZ+wdTaHfR+lOcd6k
tZqgbkb30F+tMGL7AG7TMwwRKpK2Ac0oA43L6cVgXZehqz3G8s0vZL8Fe5Wqovkl
Fa3sWxiHvkrveL+vHLOhFR3AGQBJUnBTjT16LfWgSjv4qqQD89mVvRTy8R7OXKTc
GCPA03oFIcaV42BtJY4bdbEYe0yzzUUkOmB3NQlSD+XXlSgi5L6TvAPs1gnFLN2H
3eMecvGohVBWI8ex0VZUGaoKPWcs543W/TMvrv+osJP8qBGWVMqRFnvDjAAY2ULe
WV9ktmVl4KJMnPJRUrb15G5s3MezFyV3Gc5wfnBB7FYguxL4oW2B80wcf99P40wC
FZvyTohKqpVquhrO1qjPBCFUm8enp4gfJyeIUWlTK2BDKE5i/eLCigAt5RK6zOQd
l339pxYCogvFAin7YaOPZsh47fLDhHMugddbKV2YLOkT8RHDfiG9bHBaB0wc8hHc
dieaYU07+l/1OJ67LxOwEvtMcV8gAuQ8vJCB+jd6Er/mKVlCvlC7SwLc5BQ7dnaD
j/pyzO5v2QYI9SDLFd2x3i1mQg4PR9043s2aMdb+k6NFPEqjVlxPXIvr3pimAeHA
CAdv6kYbLKhTrEL3AnZXzt6aZxOH5sxG548CAkhWH12/bcOyNX6d7cBsbKNwi+Kw
6ssCK2K0kacqSN+xzshFxJWdvsI64yToqWFrn7cxIggrNPXtVlhortmF09+p5FTq
YnBa9gTJoqMIgsARtI6uTw2i6Te+Y/EpWEunV6ShBKpYO8RS6JnbqEcNa8gGekyB
FFG8dE3EQJ6cVM1iv/97KaHpCwg7BGdldMC+bAY7agpbnEAdcSG8gNFVghxzbYCa
ee//uEr5mqq56H8CKnATgbrHVlTI3HeDEmBXWSLYI1PFSE+LclfcFbSJ2S4iXBpd
VvWk8g/wupy6h7DBU++IVeLUXrIza3emHT0Rfwp1GkSsOY0FnuFqR9B2DQPZnugO
3RZE/S7pw5dTpvehzU2WOGWSX1VbcjHz6eCiT7fA+vuNduWvvUu6hxt4ahiD8lP5
Y7oJTqyTSgN238hhhVxuWmlqOKkNZuzRMU3D4NXEIel75bR8bK2vPP6j5mba+rJg
P/n4qb0jyEIvl8Vof2NfsNwtBpI1/aQA0wXmCYhQkzl9zlnr3jCaIvszginp+CrE
6rc4Acv2YdvkmNiuqSg6ApmNwM8poWX4bvJnOeosl2Mz3t64JAqNBShNNufiNnhN
qHxTZ8MdpSApCz0K6tpKlfRtGz0ZK60REnB7VUksWXpnQTUZnp1bZLK2xRSXtsa9
xkZyezUMkTfQetceoBCRX798OKs5KpXavDkHPthkclQKEx9XiLVnozvRXuiEFyfj
BgZNdhtFlE/KWd5IAKbopKXD1qHVzq19uobK8Ee2fDgta0Pc96rEvC0HTiubOl6Z
50D9hoNr56vL1YOKqK2HP8t8S2bRlN8C3edCBMyY1x5AMC6x0i8jD2c3Rw9cePEl
YKIX54MP9o9QaHYkFFBfsiN4Uvqic6vKl12PHutYC2RWsQJSG4dOSxgGbXStQ10U
Y9344PBKOiVKkuKXcFGuZ9FFogEguHvsNEEUcHbJDYz+IvxfPwiTJ44uUFE22w5Z
oFnLDbf7GjxsAcPg+ipHYPfxzxj6MpFZB4ZJiawhHPDYYsl/BxPVL10MbuF07fkE
3YX9fxKb/erlLC6B0j56XVvSR4WYLTk3rH/+WLinyXwtfp+pm7xH93vd+Ez8/7vx
cvtwMLaGtzCRMoPJAcPd4TjuwWhVTFNc9ueNtcwGRjS8s+QPbTb+dlh5i14Pbg3U
+rAibLxJ5Xvn379L6dAtGX5n6sGGQp3lYa+0uWlfpRCN02JleUcdczhCL2muNhYh
H7EOe1slBoHOALp/gfNuHCgK//aM2vxxaRLqPfqicbGTV/7FtNNqrs8OuucoNR1Z
jBefQpvtuYCn7DkPuEYmSBDPJaqYaH0yUBDAnHbQcMcJm96y+WOOFLM7d6mRW8B5
/suZqRNIG7J/hfEdhuGvOEE6wCXDQ7Hg5xt2vbQoJLc6YRxHCAEF6nais1vIYphT
aa76C73LezKK8gagk93FGUGnKUKn8Jxz5uc/os63go+rudh7uvZzcXv5SreSEgNE
wNxQYkhhOEvGzs+GumGNTUjqkbAe9X9kKw4rnJtgg648jrCaXq/rY/VfSMOS7ngr
Ga1ZI+IdDQGrIWWjipwmzAdl6Fqf2LIZwtflIcUV2jiuY/VIi1ywxN7PTisinUDC
QUkvxBy1TwAo4Reoes3ld5q4MOht48sev2mBqr16Ku8vas7iVNV3LJMV9dVj35o2
cFfx7YboaShA5uFuuRJ2aOdC0qE9IFSZc+TooGNvZc3I/A+pngcexbJtbS3UwWT4
J/KgaapnAW6gJ86SwQfSj3ezMqxlCwMQFGmUgZbzPqSCGtLj20BJiinLojyKfC5F
/jQM00P5SNfb5Anmhuxklqmu2eeJRsR1obvVHMhGSpmEgp6bUEhTa0NHva7NmkbA
iJqp255e8ZSN/uiJfaMkXypB4PcHkXHHtBCYL7ct2LgS8NSUUTcsLZU8XLjp5KhM
baZvAn3gOSvIsGLvhFNtuy1Ok6EO219iE8sy1xck0ewJoVgpIAfFcZMVyfhMt3TE
gAsmVdBz8Nh2AzPTAkLM7o9QWFwDcVZCPr+q08OrVL+kYFHa+bGYG7cu30UYNUog
cVHJIwgl1/cgrNu2fyOq7yvTv3sOmWqJE/5x373K6FQqf7K1eYvrPchx8jqjmln+
Q1uenRY+KFxmP7W3JMShm2JbzF62OTRCe/ow6xvElPiW1C9HYZhC4opfkZg/L3Zm
gasHtKIdq1433bNSi/aCo3S8zJLSEpEjwdX/sbapWsNUOxd9uLBHBkqm7LYA4NL4
JnocE8MmLfcIcuQVCdl3mUN5Nye1+MPuoqiW2N6LI6jDZRxmmnKVNP+IBcARgxbr
WNHfb1c6/3VwUFO+aYAannDtVSj5HJ9v1gVXdr8jIQSn47EUD3/14XOCkIg46xPR
y3BrT4tBaG1suFu9NibvmOjHWwAeKNteghwcPXTqqqh9cofJcGZF58ZSOQdWCwEZ
Q+8mAfEt+b3QebUjKKbbhz36DMwnWVorQt3gWKj9BmTptHhNND8h5rB/hWuhj7nI
gh8OxbFKkV9KjMWb9EHhnEY93BUleFGwlg/l7s5YoZ4ifM/zk/Oei3OS6eH+p/sD
DkqMiCmdNACKbJzScVfZg+j5sVqd8v+DRDatDfJa6uCsul9mIJOROsZwhAqxUrTB
eqAG1WTeSRHrvQPbdf1OSMVDQLqNsvjjUiJwk1qKnn3Xy2+CSUCSl3Y/VATBl4DL
lOu6+VaNADLqDG0FlJa6hgVDtbUvq4p+Et47soFxNXTNnne+NzOsJPCU96O+5DJE
ML86PMO9sQezuwTUx4cCY2TZLtG1pzJNTz6n9yJuh4Zql9obAMFYAgQicRL3OZwQ
u7wKlycKmLM6RcRStvY/0lrxEfLZ5c2Oq595xX5AxMC7TajKwkXkJ8jkNsP1KQYR
x1sbWolbycaIpZ/dsQioMAm9TDbsTtI/QAwyb/k0q0sfLsqS884U9mbu5QOiZL0u
QnVPFwSrvatZygRsE1Yz6qr7WHrSr45eEIyeiJsUX4jZarWmFyTurGyPwVXXwIxP
Atvh4DFwLRNKpSxVwWCPgMP/lYpIisiwggu5qV4ocHjzMIe2rXhOetzkmISP2/Jp
6lBwlWSWHXCmS5A1WmS3noZuQnaAcq5hXmIuWWud9XQW0EahqMnqEVI2+1ED2Ptd
KzgYcwGTUJFJF+rkSkVNVEzTG0kyDLCUtZuF5rWR88QPUNeHGegJZGJw85kfPJZc
OzOtjoGmToVl1JK6dsZ99P+OprW7eTSUrBi47TCdstfwcuyod+ya5c5iGjFFvnSj
HbdoFWv4OQAbg0BF6NwZfnrEmq0TjQ8D90xPml027cTPXYGW4GGTJCZtnLAVhM+l
avw5N7Ge/oqctZQ3R9X5IIeyxkNi1RQWhgcOElSbGnCTe37kECcg37K7vLipNGkm
wZk3ELD6livz2EX5wroJJYL8NAd/h0cFKyiw/DA+q+aBXuTwQPWA2VKg5TMO3q+B
IqjK59UehMFUzU/TQCHrTsjYz4eLszNKA1J2QJecKerRN5mq1AYmu4DWCMz3seeH
vHUJJC7GFtUSp52v16KBY12FzGt5IZnmidDER2+ZKHeKLb++9jhKqS3YG91Y++YQ
ymXqxQtS2uzRxuj5oTx0KaSOScTv6zgP3TfIPuY019q+cEFi1ORYiEAg8vkinZcn
uvoASvDnzwYrg3Torfjx2NEuq/SRT1RBdTFI1jB3luxkvoyR+4irK8Rhvci3pXH7
fTyMDYRN7ZkKn/6NetTNEHa2Xgz58bX/J8fgRANf3sDNIbY58C23tARADDKx2uud
0hikZAjZzjrKjmGwy2TEYpC+S4CRGg+bs5o76iLOyzSnGlYt12qVlQlddYakvERt
VK4oTRBjnRzJ+yXMCc831aFzkWlagPHKRoHRaqmDlivoX/WSJ0UFSg1wwVplkgVB
0UPqblBeW2NAcCuShfQdjSHyEBsyqNEaW2LpQkid7B5gpPWZyvwRm1+/M423YfE1
LeMcQn0ux9p1yNgVDXKLfqBEkFiHQ2JgUyRBVM7ZXCAjuSMdcKjqXkvxZI48AnpW
JZsJFd94WdTXj6x8o3o0h10KhKz6La887FzCKgneSVCEb8J9RvI62oSLqA4f61tU
qx7Lc413AwohGUq7YHlzjtVeMY6mGWIKEYldLFj5HLL3P97tu2xe3ulqtnRjb7th
Tiu+2PDe4NndO8/NL+mAkBzrNhUDlfLpN7y+49NrXi9l69zuqfyMFt+lKyRHc8s3
0d+wwJKu8K3s24WuInSFA2c9EF3zknPj+VANqfTJMaOTMCkE3fFE12QF6W1kWo6t
SsMCp4DiAFCIQxAd1trtlJcEbjmjMDfPixGj90znUVbyJywt0tHeBFoLFXuc6BFA
HZnu9QNn1IcS5fANQ7BKg+Rfqxgu6N3Nt3RIf1j5e7FWcSPoOirt8LVd01h1edQP
3fJSBlc4YlHTqoWRqwMLGNX2W9dUB9z2/mapc7xkhALchqTTkxG2wmM5FVYtVVvE
9x3ceiTdJH5Kp2aXwU5TjcM+LOs9sWovOc4KR7SvOV8jTfvP21Q1J6/uPyjWwfsj
L+F0nGnK/CO1a1NlMzHmSsW4QD/zGrssxq2f2WlWWOlOduZQ5OT1JdUJnn+QE8Yp
r8Ea8Ypr0j4AmciZJ9BTBO/r0JDm/n0bEMJs7sq51z+JyPuBWzkJOWTiNjFcM5wc
5aQe0RPwDWKA+tTbl4I3owEGH5rWm6gsOOTs+4qnxyIKiKAkC5CLUrCwjf583Tpl
cLwkNXBklxZw2V3RuoCJimqpRxTbClenW4bECwCl/XUQfGhnJyNQlKjK2DUFIPp+
K6ouxKf14pH0oNcD17fzCutx2FgElwOEm9gbrqK5R/sw1zoRnOR+awxhM6sSnchG
HjPlnI5m7gzUSaSy/v95nQ6mGyH3W7lKz/1HCGYw87IGAPBctqaWMJb8BYjbx4fJ
Zj8pbBBkZaUtSNIJJuOTImDm7vdjtl1am7hBbb5YmiQazv0FzTwJJzrsh12wGlEi
mdr8hXXMkO/YqC4QNov0pfOBf883w7bZQzvBNbBqJO1kBtkeBCpPijkH9TLrWPwe
KjTT7w59KGKRcC4Pbh9u4qQfjsE+a+rsunYqrVzDUAByVkyDnHTDOyPKFWmzdlbt
Ip/kFdvmSYCLXfETJHMw7Li4ipuYrCTipVOz55rRedk6lvIwpwdA3pD4gnquaDd+
7pKO+W2/npOmFyhvyTyeC5UIHUcLwRFdsZA05PwXKiqH+UzdK4Py5LSblRCp4xVY
lSqukL35s+oyFmbHINtLN18fIUEs9L5zI6Zhyz+ihJm4Ev0jVfzmyoY/Lszru8BN
/4R76woDcHLrKUPvI2kOD5G/IbZk9tsrXGE5uFpT0B/bzkO+qtfVMi/VInBfMNFE
ZXwmykVuvVHkpm8uFuD4X1FnOLwRng9Uaw3DJPo/f/zeBy8g4VdkCMtQ8L3Tvp7+
idASPv5VINR5k0owQlXavPJdK0z92hTr49cDQTmagxZ6bOMpdpNjOIp9uAE262U1
NHWLxjwIHo97KHLg6giiOvtOZjLKG8BLXVaRP3YfVqgAH/VwRcCh8SWgtGFwWdb7
ha2ihDEZuusjDSMklfTx0h+CAcCQoJI3rWZhi6zRT1RzU3jLjpai1QtQRCGSRPsr
HLvo408r2OCVROvydCKeEpo1hXEACyxbUKAdvRaOaniEActbIfZsIzIF7Is6XXtK
uEmLZ9Al4ltAA0xAvbhgiaksxxHzfNQrdlIH25srbNvgE8f+yj+CqluXHAasex3a
KezUZinapeOUHs3aQ6aElthSn7+/MBpbqQ4BfFFpaeUFBlM8Li+gkYCUEJIl9ZVO
FenikxQuHbQ1w7Rni7Jvu6ehfEd5wAcDoUXvqIvwQsNLHPMqqwUcA2p38yvqrzq5
m4T1gyj58UoAA9WkqhIWovPm2rG5HOD7DJTckz++fjNsN3hDzNYmOHnWegEzeCAU
NEqqo4a+w1RAwYH1XnOOKVT4GnEOysezS1k9p3gWbha4Zryb9Gt/1fS3qFn1Tbe4
JrLBhmLDaAjALcs7D/vTK7903IDNfgXkg9Yum366P5xusT6majCilfBANWHW5WYg
guDsW1WKpWBlCuhWw/oOyzrCfS/Tx0gCSiqBI/emiIiE6HhlVdB6oOgRyiVIZWuE
0bl1bKxj6mcM++wq2aJxqxh7pQxRa2oXrPSP4ow5lkp+zS5U3wJlDo2S8xRwG/fR
zZGdWjBE+YsXUlVN0rwcBT2t87sTG/t0WYIpLfCtUP1mbCPVoSHajCmgUTBRbDH2
4vwBbqZmL+gQVXDi5zzKOMdHmKItdglqwF9c4FYlZxTuS4YGJxdRwenaqK8LBaWG
TDM4qztPctQnyvW5gEKh4kKScpb0/P0wkQpaJrwc8/N8l6oAnnmJE9PBXq5mHnGD
ZE9ozDG3hJP23shGGaD5MnVkwv2DhZF+3KDFZhHUJfUbMFVBzSvBeaBLgAEHKsdS
ILskuVF1gXTy7DkXenGrLC49EGR6wa6aTr/Z/nipyIwiphYVqxe0eV9m/w3OlgJ4
XbnA8qFeN20WNP8nA23QntRX4slUen72sS671yETemweth3K5znKHTBS0ZoIQnu7
gZQX3QcbUyl0fmt13CBkO7NVU+XWwkNl92x/iKZnJgbVGlaKdSanhSCVbB5zKjIM
vjpprHm8ulX+MQF9wyfYrC8pRZbu3kfu2pI8c2L+vxxe8JqgovBvILY9tSPnFnUE
57+SLgh8+myYvqb1Qq7bWw0jOnEh1KVc4JZFB9tzaRGiCXWtkqNQfK+JpNd+bJWT
zzGVgp69nz8j1UD/5H+0r+m9Qyk+z4CIhawMb2kuu/5OTMW+7YPT12lZ5WqadoSi
rHjgotNquOI+U1NRyLb06OyvhR7bzgWfhEgRJ5rh8YwFirZXzh/S8LaeXZwPgARu
DH3zvXHeL2oX2uKAc4MVxc1gLqgM9Jihj8IDRL1Oan/NvrRrcPSMmtYfpdW2Vk0K
7wQS9frcrZ+6ACNIiQqCVRgNohi51+OyJP7Q0KTt96ryjDg3vk9Nefu4LOPIJ3eN
52m0rkxDRhi3Oeq7zTYcibZs26zsxuj5xI9EQiddXgBJPNr2q4MMWAr9jlM+/Xt3
gqS17J+PbdzeGcpfrSi/q6tW3w2FqrdwI9VYJRi4cMgeHzqjXXTAX4KnYj8avNZP
EKnlAfpfYn9aXYQo2E36W/9QvszMzDItmFgrzhi/W3RSEBLZmASJDOUg/RlJNuIs
KL4OHD8OXgL5MbZ5HKj50rskCh+hAq5r0o21JBqyeLTpwcS2XaQGzOHOAGxG2Sqp
VOy57e9WPDXFFPcNPpqPco9RvYkbFRugq3mYrznY6Y91biqHuYyEGQKCemfaMBDz
vlLd87OTHnyf43bohTme2axogjxJabxyh0gwJi1nrrTVA42bDq+Et4TISvn3Tger
qm+2PRz2P6FIVu8bVMoTHXdjYYuUMa0B6LOcRbg9Bs05UnFmGqnLtdHnFYXFw65r
qqUiWeLNIlvNusnnnSgW68Aam7V0Pwb/qlkLHmcOJORJYReZm3wrmc4tBNgudTPF
/32eeZr2wOwdgbA+ydRi4NzMCMPFS0Is4QHTeqTrPA0no3loOoVANwH1DYbc4GXh
hJZq25yM2KxhA1x4MxjEcM1nCAtmbLzPBOtQGAdbLVXPJddI8satzyuWQ2X9H6fR
SPAO5l3djcd/5eCAv2IJbw/yWyapdk9D4kb3euLXjROupBQGLY9j/EElQuGCrJAn
JkQ9lPFtYE+yJrYhlVa2cUkSEvl2xuif9Pzx+zRtgg2PXCtG7w/5j7OAYnMzlK1E
4l38/eIgZDhybCMbiGlkqfgCJdzgknCMam+o90fN9fvgy4mDki3lRUpBUScZUAqS
4EtecEV7hkcKCnH9JjNQj6CEa6n4RA0KHxD1S+QFpj+mCktguBxoZume38Ghxndf
d720IBqiFJ3xrXJcvKmsI6GTlXS9rhb38f+g72mvcWRWr/aQae0iy5OKrbMeb6rS
YzFyiknyztI84CUr6dogxapOdAOr47Zj9Gkzi7i3dbjci2S4T2Op1TdX17Mc0r0c
AHLbG/ledudQ/v1WoPKtTUYZB2xT+QnT5nT3uYmG6ZvOfP44/cf0wiQPuHValdyv
gbtmsPQZ1kPq6GXP3KXQK/XxlL3uXG77CD9dYwUIFlU+GyaL8WLH6WP66Rs5lD6x
lC/mxu64lZR/L1+p62MynOrTpVumMy8IVpbpSRZuXPbZZXqCfMGtBKx2AJZkDhFs
mHGmaEI/ikgm6ksqyM8811aTs1uTqwyeyvrxw3fAfaynUr3pcDzO3djYhX3XijCr
kmBrigs9uRoySVA/T3x9cA9b1ConOIsGysLdOUSKT5sV6/PIbiujhH41GuP0Fty2
RdaARkaro84xqSY7fVo8idSZxiHbvHmhBpN+H6f15uzfuby5cikLcR/kCZJGfZUF
UvTKev1XkW3lahfiAO48QLOtmRKZ2T7bMB43jquukBIWB/XWC7viOBSHEjTDV/qv
0GivxAaI8wltS05exdJDF3oVm+2v4glxDmmXf8UqUVeMz7tDnJq0oYRFSI4hrCP+
98HHJuNskKC9bP5MuHwxrDvIxOPYeM1e/mZ33gs0nurDyf4Sy6PVx1LMEHSyh+Bg
2OlWA2R9oXdSA4w9uazNhkozHFEI0v/19lTdjfLHzSQtdkpqFkF6QBA42PhLHiNP
48VdQXmwRh4o/sYWJYtVXWdFGnIDDiyBXdC3lk4xTPd2nRi8nXHkJExWEJsuwK6u
RcCE2p4vqgk/A5H/p5LTcovmaiVsA9T8QIcd+qR6egbViASDuHgLdMOmIUiB2JY/
kRFLuON5ZFvNY8H4KIVJxhwEuqAGfc2zWv7Styzex42jyB+ioF7t16CGmEWaljnI
6XCtzyoqi8DtOBQHMV37QT59nOm2x5wxXLxYRhJwhlTSIDRAA+1eW+XPLPMdZY/s
I9wZHzG6xdDasombFvZi9Cu8yoSVHxyPOhlBGmNXQomhvodo3sZ4E3ZuDJd+VQkb
5mnK/ZgY+x/UQJ/TY+5dtvKUzoWL6/RmQgCFAy0wHtiH2Fgu6AXjZQG6Ptgj5RdX
jFmvYyUsilcjiUCCaduKi+LwAlKi4p/2wSyUYK+ukrwgKZDCwisr0EZM1lMqJ/t7
VKNy8Cc1F/Vbq7oUdnqsvF7p4msVJYGhcSABnAPBJvAYcsnaxtZ/nXfj3Yi+Y4nc
s6+Sqxr04sUfCGESqHNkaizWkSXyNeZCLlaj9WIWfyvgo+UmCx7Xz7ALqpN5P0ws
Ln2ap6ZiANFTfvsWfZGME5azMH9FM6JQnrXHZuURnQajT/p0+S/DL6svifvvV4gR
w9o0WPpu9Cmkk51spbq+ZzGfWdan3P+IouTEWIvhoVNmN1oe4a3wCWihbeG+M4L/
3GSwmvAPo4Gb6kc0egEwd2tKPonVyv43tW+eft2UQIK6rZyUngd3dsAfsQsoWuck
+bHohM0u+fwxcOo+Np1ukqozoIUahI+nYabXYVnYNQxRYhlcgRAYGHTHD2rJ96dd
dOhqJkruDmpEdQjO8zR1hYy5R2y1wcxPRzjHuzj4yTpBPXVbhvqk3XgcpRsePwLi
tQQwvj1EKRDTbyHvLxcBtJJWUnfy4kTGNikvL1kyVeLgrmEbPhLtRIfmgYwP9t9E
5cg3RkRtieGMIpCGiMT7naRY2DA8kZoD2zVJw7+kPSRY8y4PudzKhpnzKAEnuzfH
zDEFkUbLCHGOXp3xMv5853Ij8MLAt5vvhttNJ2AhJUFjlwPUBZ/FpQg8KKM+8FSO
dU6ZQV71yevv1pOmFk4bEbJHq83X5TVzSidB+42MmGgl2SrjjKhomc6OV4QNOVje
bHB17x63S37UXZlFSaaomo6shxxQ08cmLoSkR/Z29WIylTbfhbDXJ6l/6HGOENvj
e5cxRSJ+NzkSXxZDtlAqMn5jlPofr7KK2n4AeMajdVBNxgYXmgBybK+0faB0AyZT
8Nx0n1YfGurjmt3IaXFs+giUVk+sGET4nb1c7j15dfUfLhkb+8s3K9+eHuzmrPyA
/X0SquSlpzRWhGx2yTZhV92531bz8GKXerkn6q7YSXmDWh33i4HnzLynB4o4DnPD
0tTn4FN8piLVa1WuU3mVmEitliFkHHyt62rwKKoXqWCxi5CJVoCnLlcDawCXRTsg
MFTsdUAhqbvjeabe3MdAOBXU50XJ76AftB8QhQhghB+cr7T+NmsRuUfTAb4e/ht5
cvzRPaAVfcaNJfXkvxB8qFCMc1uLFOgXcJAycmM0zYUbZSC3xIiQYtEgk+qFq2ns
L4TXjS4CeHao4MNJcceRSKm6Ke/HLlajtBlSbAK2stY0TTKQtwIBe8qMzeFVLQgN
Yc9z2cSc4e90WDEwM4uiexBseBIrNRqHV+NVPf3ZDSSWr4z5q+Vos7+Pynyy7VK8
76T3pK9EBfsk/MIc41iGrLpTxe9Oc/FdhbWQjwyAmenr7jj5DkZsQGJKR5LnnQom
G+LoHVih4Rl6YJTT66/aqM2JzHebQ3cJIyN+7H/oy9B+eBCDqoEhreyN+6wksRo4
aCw0rJ6e6IkD3oiUgjTf+XHDxXMQ8u4xBmoF2cLVhjNHv8E6l0uHERj/aEzazm/s
ljn6X49xZcMS3322RJJoHskJPaqloXNbJbTIh0R53iRNwFuVmV2gY9E0SZxzHWGS
ywABPQ0PftjdTapkD/H1sSe7a+VcTR+EbKlSfJMxUZazgxEttFKoTscPjs/nFVNH
slzqbyjyYvBx1YX3YmecQq2npy4w3DkUvl8uKxaQi8SAS7jfJfjrX3uKWwmCCYca
PWDldbCF0XHdZSCxFI5KLKrpvM09tMHmzouYLiz74NADCQEeylFXI/iE/cc9GfVU
YTIuZC/MWS6z/CQGX1Kky+7NMSHsJtuu6E3VWql9YXuSp8KG/njguwELKiADC4QS
dkRFanfCFpPl9aaZo9JlTf9brTqFk/qT5Q4PlKKbd060Ub81CufuZ4YPS0dGqI/T
c5rpc4IbJWUO4iofryxRbSnpbuEXGHIrOPcnG0v7qJZYqTe77x/bK63n4hPFcdcA
EjtOG9DQJCQm2WeXtDUnNd1alRTaQnoi2ZlXIW31UsGTbfHIsMAZE2iaCsGziXJi
2IlvsQrstHk5uJEyXB+2xxkh57kvLTt5LhIMICyjSZieCjLHmIGzBZU+DPfXSymj
dIaIkj9S94B3OtxnEMQ1Y5GNiQU7sxvZOTCwVn8emEThU7VI/EePVeLC74WhaCQt
WsKOeSEhnrmojcicZDn1O+HF0NB/eAmjCCm2zJv/MQWozh+A2wT/zE3pdDHY2/08
YtgJ3xSae2LcOCMmlTaHOy4i3UP20wlzu0OntoMHcyUbjZLMr3xlIF0HVImxhRO9
ZEvga9LrRqVCzHk3jDXgFHgdoFpu6Xfnsn9B0F5guuNz132NViz+V4Iu7t/WGQHt
7Ean6B0Lvq0bVg/QdmL5RXclOoYspyWLm5XiimKnRv1TnJwf0qQAyud0d7bokZ56
GV2g0oDAuCzGgflylytgI60ltrBQ0cZ4xyF84pXYOHFCsZvvnXHTfrbDfVf5sgNu
rTr5LVonq6CtB5DcMhlCBpIG1aia0wS8PF1u63orBdMxD7S+NNVkdzwOBOMgbolw
Y+ARWtvjqpKYAPGg+dqKiqFLN57w4CVmudcHs0Eh1XQbUIJbD8/cCSMofvWeBWiQ
4eej0eYKkKeL/oL+nHqB9C6iJdCWmGr4T0Ho+E3bBsi3JqRFfZ7j/juGtZIf4pJC
ZL+wpHEE6e4o9/2pVlEui+FmOYmAl+a/n/vyKRhskzoE01WImv+1mlhBGSE/1Alx
M3TywKGerpNfXvqc56exErvGOc30NJ3+IbvhoxHZyfX2Eu9/YGR45VM0+2qlgzwn
t7TGdTDKgwKVJOKxTdQxRyK6cmQRY4APAdaMeUkfu60KdDWKHCcq90noq85/icrF
ZZYuiT9feOlNS0kTufG2ZL3hpg+8xkjPNNMZnPLOD8MnSDA9LWjzIoS+XODuILT9
8ZQn2wPob7hYE6kN6gpzd+Ld4l0IeRIVQUttqiYzGXzk5n4JZjLr2NuCO8gmUXsT
P+ZDjCbBAuTLrBnwPyhogHbs3MWHau5HGTuaskiWEua1MX+LmeaxAaGzaj6x1SIQ
aWa10Qy5CrCUxmHZZjyH6BL/I3hsHzfUDDPihiPoj1+5bapFKnmPn4cpqtufVHSC
73y94/pyjxVm/FXpUzb4eRPjPWELSUBhPESy8x9J81/lb8ERgvGvW5koyYQHcC3H
XXMSDSQMGQLW+rq/T0Uagf0AKzJHQPEkQpftvmZJEDuJS3+bZNs08g3OAFIxjQbi
3AzNtbV6MoaU8b4nUp/IBUyeBdO40YBKJxjDqSA8oQsN0eLemZMJKblyDqFt3uZB
Jyk4OfoyoV1kjDS+C8pYdRbshhydnwBFixY1PzdO85bAa946x6rP0l9RaY983U3j
wKkEEct66NeaQht60CsnDWZRFdyG9z4jBhsGVlJaYJN8Y/6sXqptZzwFTlxteDZA
gCpiKP268M6kUtUnIMm6RJcIpUaNuvcITm31421deuy3OkxOap+ugaJfIAFuNV00
xhDJYHrOdiztJhQC1HTz4WiXUgCqB8wOmJRX45IIhVZF2eNQG30d12UiF11UqMKk
RaPNaqYbONQ1W5q6ZaHZMlLfYnkLRpJZzlU+Tr9RSZJesIHxUzU31Dx9uhjBW4yu
U3P0H92k0trs4kBf9Pi2jkhIbtf0fNXfKQKq2ZV7Y3GgIEbIsvilCokeH6tZ+6Jv
dePvugbWjOE3HXMuRwCP7KY5kp2RD7N7WG+kcgiGTDARtz8TDzvHIo3cuNc76BoK
lWSzyCWrMyxYzGpRWUxeOwYplI99gmHUyy8R64s58h33oWADlMQp4vhfa+BzBjym
Fize2/foFVlcdyx8e9oLX1dr9MI6wO6D8yRueEDrhz5OAWk0s9A/eCSNAKipQ4ur
QLudmJrxDBrmAs0mfnNh9ZZXs9m9tKQmOQ89qmL2GQEKyyH5L5UX8+Cy2+3LwjEF
SpJ4QkDLXxY9wLgpKEhHAbDk0QHtqM/Y8FmkjBSsM/8G+5Kz+m0JP9f6h5sU/OLW
O2nj0HHCOrtcjr3xW0liHGAGq7AAb/V+BssQA6fHdmRfNGn5qY7Lim0cz5d4LQkD
QFjUIwsdkzZ9NH/iyM79KjQ7IN1Hzw6YDoxFJchkyCSP0pzGq2tQjyqVc0u113TB
++Ymf6BYgkSTNOk7ojaASTfJPnylV195T239JGwnLdfxbc4VVtHOHYE969LPtKlr
ITkqV9TbUf61DLzAQTJImOuU7bRTKSQjoAV6X89WG/GJyUjKgNfc89XsFEvz2nYy
CpTLE8Cm9hYSRgOT4gInJg38hJ/PCOGOKUjttdNW/plMPeVOMHdD9Ugb5D6yJE0Z
q2gR8puC8mZQ9NJw3XyUaZwK9Pu03VW5djxuXVs6IStcr8886C5+AOCryeL9hTNJ
nuvlAHEcwORq6S2rrcTPfXg6PeExW068XheYuyThYagNHHZ/RpvJLKV0Kz40uLCr
nZnD7P3gRuEOCDRde+1E9ZogBhkAx9iNYkoORV30+KdZB5pCPFWD4Q7XOzpQex54
s5YsoT+Ok39ROjID9dZv294TbppGUN+EM4TYWveSQOyiEmhYZHPPM0irZQ2G/ztI
Dhal98SUzRJBXpX9ZHBlUCpgFl/wAxmRTAs4RHUu60xFFQNzABBWBAGQt6S/RTQA
EvA4RJ7i6iUQfxV+XciIDCgzs6ZPdQq9YzeKx8GwHYfG9/QucfQD2yJ3pSghcTbA
EEyORdi7PUvsh/UDB8SJkulhG3YAIL8XOqKfKw+Dgty1UPmL1n9juYeK4NxcDn7p
UmsRvdcfuSa34VjFyDpExMiO7v0syg6mm2mJXki+PlwXs7d+aUOOWCIOaEzgeSMd
B/k7v03TYQzxE51/bQ2q5uIuut6EfJXXAWmBM3Z1Ckd7sCbpeC1oxiFXUWHc4sre
yi0y4+R2PGzpWzX/VjZbs3MqjeaygsS1pUM/AUGOSj3jMIAe63Hgpt6xrBaTmdQY
gKfUCy6+42N2PoiDwnnfwmWntl3Dqlfp8REKysR5UMJpYq5CIE9Y+mUoPMFowHfl
Slft/hPawRFo2fICoz4UwtKb3FgwoGHAcZkhVg5cNLg7o9l7pVer0VkcGMlEgTkc
3pQTCoRWKiaCdAS1aA0AaWuJBWG5zGsCRw5L/PE0S13T8qBXnNd5bhvQpKG6lcpS
wQzyng5W2yEjbYI7g7SNGN8LfW0YsZPDQbu6wieXsZIO/wzvVoEb68zHxG6qewuh
SVsrQ5/16QXLqEO9yA2pw4mnL5GfO7QGc5YR/ZUqHWUs2iTVPMOfO7x3CGoevpUb
3Kz2i8LBIei8QVLiCwxrGGKiJSUwrTp/ay4zLYchxiueKWpsN78Ylg1DReBwPwL5
A5IYwOj/rOzpcb0SWYARQQcvJYEM7TSwZsttkcryJY4QAFfPFiQefWMzhxKXqjhL
5oleO49YI2XH+NU7Huz1a5iP/swGBzSz3ghMSi8lTe2R1iF2n0Z6z99nsLDMx7bx
/d0dAP5/C1ZRMOlna7MGok83J6wcGTmc/Ng3vnrAW7LZF7C74X3rLJrGWM3C04ts
nIJowmjmMm80yTCcZ2zpjZXtY9vzWLSzXLlVASV6/XyFG8H82m4OwKpSKzT59x/b
Cao/bFzB/0stJu6DwsUPeWjREInQQizcuO0ilK4NMpHmvoZRMV6K/q1HlAzLNgRr
a2V7/hkuSbcsDf5jCW+9rnd9Pos1uuIfJB09kzQ5n4cFeqFtX2GFkQeHpy/bkOWU
rD0y1Cq/5XhhnO7I32tV3QRrTgSiQD960/G0LS1rZ3TBLS3B9VPUSPzmYze5V2nF
tdARhItpD6yBHN/bOC+F8HdY1w3zRNWVE7KcXOd/c0fiatp3eGhTYKr0bc07QyAT
DDEkK/YUitETksXSd8pq0+NQcW+JJOr5qf4dgLetWr1MEApTfThtEM8YG1rfS+oP
4ZWkCDSFtepDG+UBGzDZV6zbTP25wX4oHedPaBn2BHctQUGKa8q0unVeNqbhUFtL
uNb7zip8m2fo7GWWlVfk2XQtYUibosr2WwVqyz86ucmM0OMHYQ6sbCHxOZK8Ev6T
u4DKwmvBroW8aEWa0liLXcKyOPQ3qEYar45aJ5FftsTyBtftMAxIDMZWP6VrkqPY
+JEgyfUGRUCFK3B3JWwevcFFhb3EpeAHftdk90e/m+liMmrbESMTanKtlOLIFnGL
d4TtaPMdLO9qa2QzD/3sW+r4KCpbP1Y4tqc0FdXj9/ydIwB/TSqePVKp3+O/TjAJ
bF2DgT8qhZ2BCounrcCQR5PKBSssAC7Vp/3B/W2bMNysvjwXmyJ8Z/zACYYk46oF
DILalhAVSye7HRklvy6tp2Qf2yZsQIG2dQol/RHKhi0Z/EUy4fAlHVzNMJuACHZy
686W+RaNPoL2Dpk7YD1IeM6Gx7g2e3YssH/eHkDoJtcKXQg47t8Tz2Ds5/uOgG+0
dbcd7MXzxjxBwPvPpZjL0dTlDZiNZRYTmkoJf8VB32MWdVNG/VSjrQWQTyU6JmWD
GmPHoXMK46MbKiKIFt8Q0vfpIHFBrsmQPj7foVQPbu3EnUSyraNTg3goIybc6fIe
Cg3UZMziL9z/NsyE9K+r4oXCInUp6yu0fFU19/r6t2kR89H4UPKA/yNJ0cW8I/GX
BzNAA01teuYeWpNohl0xjF7qAEvjmlf3iCcmj3+LE7rNHRQlbFUE1oOBBC80+aKr
dprzTBgVLGFaG5ZeJfkkSdGMDw1BchZNhd2Ju78paHuKWiwRiue0CfVJIaYj0/ou
5OMENJ7/UfEMkuSj/4xf2t2yHw1h3wGbrb4TEyN5ubhBeAZo5GT8MXk1W2pNg0u+
JGpMcqeqs6g0vtpPxKHhhdX3OBZhtW3InFy8TmoXknjPCUcA61X2KPpbReyb0Vbo
IgzFMOk+Q0vTX9b0+j+Bp0+Kgc4scPnNOLfxhSRYfJxTqBRYZcN72EYQ0VwK81yp
JTjEUtluNiFIFuMJnuJbTOqURu/Qqt+3pq8IWWVfGufaSqup/k+Ea7TDoXLoJyA+
G98rdgowOHP634PwbukevK5ZzjAyKNHogfc1lIOHCkG9I7leprxZIMDT00ew+Nw5
O01HMcWOyneIYavd4qnH/RPc/Br++vZqjVQrdbN/Vh8dpiynzfmoxwlm+cQCCO8m
QJB3oOfda5MEHZnMCC/tuV3g1ZyU3QnUZim3h3aKPf9iA6xh5dIFzxvCUhuYMksP
SDoBd4u6jRjXHVEhKw6hiKfC5SpggQso1J+nRBCzSkVmzDwUyNgtbBbtRF5On1+N
2rudyVBFoNxrwQUUwT/tWdYZxiye+EjNsnw4Lg7xybICGtptXdbRbnsNwyeOPMs0
4FITCbJBh588chtUcelcMg5MrHDNrZvNk2noG5kvcofG3jOaViPd8tebxzt7jvZM
DGEdG9i4E60Gq1wt3H4ChMDtdtNijKIs/CgXTf620v0NsSmOL1iwnz3jn1abGOOT
H4AiOEO8ro7+1xYtnUITVTCS7o26hR0ighj/zWljSx4qNjU1y1NsnMhwwiLwrq6S
ZQhy70FaAy9sLgh3cTdjoBpCvuiYJoyA6THE3Pp2nV0mtPmE7ZQq22yLyhAxpUFk
JfnlBF5BnX3Xcp/xFTvCsXlU4rYP+s6uN+4uUuMf4I44NuduaFaCGtLBZvV9/Say
T3v6j9440oRRjwVMx13Uext9ADOd8Q+mjbIyMmDsH3eC/62BZMQ8VRUX6ZqV0kKo
ZpnwrWTXXGSvr8SyhT3Yacl2vaXiuXwe2k0UBrL9DFql/FM5DH6k8f/r9r/xK8Si
A1LWQAoZ3k9ezQ2xFWfU7zkpU6RsW6gJOihXQ37wQq01LS/yWUWjrJmJHdr30NJm
gGFTG4aReei7MV3XSoBhepZOZ19xquCyEAL5ywfQBJE2e7oJr9x17mPfATU0gzLM
0MQirvkxPrPqFHUWb1C8uxHi4tKLq84onmozTbMjUJj9AX6J2MdmNYT98pEfYV4X
hNl5aT66jOw5l5rTqXUhtm42hQI1NUN2NMTxj+uzqe8s93hQbqTO5oXuxDiP3I98
BWIRK0G19JhJFsYFTn/9TCk4uMDjGxAm4jfa01q7+ZXvqPlnMFh7aiM4rHEWDIis
QUe7TwPiNeNbVmY04+6kjyxdnIqTWQzYqn8q0mAJaArvZpbxg+NkOlp9UasuwHfA
mhSJyveBBltqOUEtJDihOjRlYLlKGR9Nh5xcR7JCFXAQfSmU3BOOfZb3gKpiB+w1
VmibHsNHtNrsIs5rveNIEiNaxHAPPGRLLpNtYSIMB1vrIQKDEM56G7i2dKqs77Bj
345LnF8U5104qmfwrhHMY2HIVQg2M/76rQ/iCpizg2BmNeU1auCXM/BRhBm8+o4x
kHtDq4fgf35UCz3hESE9sFN6zd/HqhERjvmAxVd9y7x1L1tatpq1r5+GVvuuP1SM
V/4SqYcx2vNTWBohaZzBST6ZQM6tIJCUygOh2D9wJ5LACzU9jw9hxHzy8T65XiV6
u8TPH4RAC4m9q4V2IhvDhmstTSAjcBEBbTrVO4A2eFwPexQcc1hrMxxqnfaqjPiW
5OfD5VsFVOvrrihOEyHmuiv9m3KEl/0avGczeFKj+hr/I8tH27vdieVDV7J3PJS6
M/gS6EOqbBe57tpe3L1sk/6OlARB32uk5tZ+dOIg2o3WPj7zr6J5+TjehB1+BTfC
D18ElFr3Cq6BHys4PKQr37triqBZDkSsa+2fOvlkjCMVekEFPI9c+fWEVz8jaZIc
jcFOaVrU/qwogcaXfR1CoQqu2itEjT6QZn0l9nP3JgTEoq7NY7+PhIe1QuWoZUnV
GX+0iTt+5pufqIetwAP/wk3AOT8l4UB3O07Fb0MM/oHLRTuN5Rnhh7t/gYhEfc+d
92dVBhvFg/RpeX9m7D2YZi/dtuHZalrO93rFhQHv4bS6pyRky0Q4MYaQ7tDpzPzE
iJcTrZRNIpbuZTdKiIR9hn+DRGBT7vzIgolBLgXrBgBS+Pp5bIRC777Nzm3vfzmo
1pm03jO/5gCLKNK8mAZzPIs8M4flEZxL6noINUp8IfnPRnVNE8LMuVQoPSnCkG8U
5Yl/gh6XAN6xOpFT6Xh3vSWduHI0TspC0wjF4zlQYpi9U+CaH5KZu5CKh0jb3eJP
k9K7RYJNBvolJodmoZJD8r7r7NtzT1xMEn7f8fdAJO6kdUo/SjA5PSzdFYkUsRN2
Tt1pI0v2raxgYi3vQMDxooiGJ1AdRYcGRa1GzXLroB7tLvNabgcVm+6xJ7vgPHKp
RUnLeAAUc7M4QsIqTm7+o9N5+b1MDnKFEaocZKCxo7KdvDnNM8fiJMRmGyaLo/kQ
Z1+TQPZrziBo2n+1AXzx7HRMExUNtQ2z1Dbp9Ur6EYLp9WKkGNHvXg80IwhgKFSZ
rFTY91pJhURyeHuDajv4p5HSt1Qv09sOaASybbV2fzN7liFx8wrlqiSqlujP3qNG
th01ATRvLBWrMIgOTal/3nrUNEi4ZeXaitSVREmJqvKYUHxNZlK1mk8fFU/utpgL
MWvs/iuNmafxH5P/tcwZ1pUUU5HhXqRaFhnLRlWuPy6kyR4tUZtuVJ7uJh5nxJ0b
PDGYFVYTbuRGTslPdEyNnlX1ZTsIrmVbTlc7LJQN/0JiOsSiO5rbtjerNHbQRirI
N7/jCZXYFQa23Prbsph039rE5JDwbIQTWkyRGo7XUKdh3PbDwUJ5f5CV6wM+YzCE
RmTU7N+rY9a7Wa6zMZ4S/Wd7tN1laCKuHhm/oscRFA7YAjoEtMQ7TgT/JNlWwGPz
1c9oG0uMgiTtU3kTXjF9VlLFbSte6XdlHm/2Mp4Ppb3ZHXOwtIv/RgGIFUoauxRa
X87II+/vRGA2N+oaoIo507mTqMqbfyFWv/52iW/yP/D2me3iaF8/vYA1vsANN5Hf
Y2K7pimURv1cSCQstNo4wU0ray5DjT445JS+g9Qf1BXdYw6dsa49kSK6gfRs8NT8
h/TLAuGH6N4MVrsLez4N0q4s6KHUOBD0MgUgxw/1niQnWyzBs3E3uQCh+OvPOkV8
hnzbhtqtXBZwCjrZ6bt15ytYNeP/dGzPkb37XoGxCK77YUzM4Yl8eC8PmIe1OmhB
2xG2fRChTD5kiGIrhkj4hbC3yJ3BUt75DNon68YQhnkH/a2loQhYYK3J957chMUm
7O66hsqmwDOmMQ4vwokb6+yAcXpJSGUpWXyF48UGeePPCpd8G/Yetno+J3gSg7UL
s1Nro6r1fOTOpNO2zGBW5VoRJ9vn+cfHp83PCgL20nk4FatbYtNoW7ObemTLeimS
SpWGfcBmou4pSzuqo6I0ckkmclU4+UpOyrBt3oh9xNcLstxcwPSos/tYP5eT5F1Z
1xLmb8Xpyx/a0THQflUtDvd/JCUY1Dcj8t6rGdRCrsk+0UytUUJUnbjGvYP+S7xR
rMNv89hv+7eLuNN2dVqyRa5XBD+qU5/6szXM3DKfHUiFNkMROVaWczUx1Pp5S/IJ
n+YJHKnkTQdEcr4A5O5LgxjZWQV+Dtot+ojQrEcVQD/5IJKJX9U0S1jB8f/oPqUv
FFzlgfxefQW2zzjrYyAo9wYilqdlmIlC73du5VBzqqbwPbwpiAcEQ38NXXuGeeE9
SIOagYTF2ZakN5+Kihz4iC8RHcWCgdz77wPE24kf0J0zxk8yVwIODBFFUSYpxW+b
3CxHJPip3UeGAScgYlXyOwZAokSjG3b+Rwk+hP16In6Gg4paV1AhgHh/+FzG8qkP
tCb7Zz+BsE83U+CUE6lb04QXKF16jwhKYp6maFcdpGxKQyfucQUY4kukM68SVz3j
DshKtXai6CRpN/FA80EnaHKXAA0AqctLWcM8vW4PH1qctawpcVWL+piaPkezuIB9
SBtFoJrE+FTEmgN1oxXuXRmTijAv+MeGqMy/S+ZyxUt6pQFxrQJTT2PSsgNLu3V9
Wl1gCADYA/gzbeCyjAyUKzfcXsul5yiPC0vo8aovO14RhhpNahqkh2Oqb5pyQZlr
Z3UXa47y6eYdAMLW6hQE75Z782+9e4rw6A+PfQCW5myTiNKnnNsV9AleLuF2Z9hC
cLnKAtECpFlwwO+b9v3aYs3/M7pc0Kp+P3oNF597I7yxjYp0+CYeAr4OIIe4i9A3
Le+oPC9VFr3W3Cb55mioM3H3bUS/otxYFLGGuSteFBVdCFIE57/+MWTFzHCFzGu4
dWgXV4I90icC2a9XOLmcdkGfLa1F3A4x6lGLdtrQLFNpDtzqStZo0S4oa6MeTt83
tQdBKM2z3v8Q4n38vXFTiacbDT9aOW7MIHEQX5gnRIIozbzBB1rCXAZka6QK8+Og
zmCp61zxpRMRo9oR/9bqgCV0EK4evgsChjE8ZKaaSjmtISGeO1tjfIQwMH5+iT2O
pw7uIEATqrU0V8PQrpBgQ3dS2iPQ/JKBqpYnO2+YzBnj3o9dOBhqgXc8XulofAlT
EXYFzj6rUN/uBpqoAEV/YaC/lSz9S49nhGFvSXoqF51tw9S1TdkG95yX6x6A6uKk
3Tt+Z2XtRDJ9DfYpmLs8ZDcOtUAPGchWBu6IAFSrYSG3eIgRl7AqsCkukYi2xA5W
l9st/clVh5YUBcWZ0kDzloVzdAgBoyYLiE/amp3srtYvwjRPmP4gI1JBJyLoQpPN
MPd1jvexHZKrlk6AosGytOwaOJfAVvWNic7BqwfQU188XEaA0VjXs0myXQV5VTEp
ws88L36YUkdYZjOSvEDcHtIuGKBa664EjQB8V9kSqaigxsQCAVX2TewhBLHjAq7t
N6mARhBYmCMPcZFDI8qassCgshnOM8P1op+T0h7EIDIyQRT4Z8Xh+cTnxQDVzHny
XEgdWHvqaNVWCFDftZWkBoRYkLDibwacIPkReq7NIFjf4mtDVykztTfZyEu03jwm
b8jeZEOrztB6ekHQb6GZkOJu6d+RG5dlHOmQLqXSA9Xa+hMC/ll0lUwupzNMH1ET
V3TLiQOm7Q5qX8xLg3SW0QmAv8Dio+zC0kwxGFpfqlIsIOlHUIIoni4Y9TctMH3+
s4GA9X2+Z+b3pG2w5EjA/MLexOAylSGKztsfWQ5DAHae469XQT/YT6glgRTor9Bm
DwHUWXPu+dYJQmiYVKAqZIMptFjO+tvFROFrl1+N4V6vm/fg253FemlRsN7f1LW3
i32lgBuAQ7hXMQcob5vq6NIPHGPLqXDc5T0rSCuV9FSPgZ19ZmqL2ka4gnDF5vTD
Edg0/jdGUTp/dznRbFCo9bBk/XUN+BzR4aUcs2TvP+PCRi7dz2iNlrdmq9C/P3+O
VKGd7VXsxtx1jOZT7fQvwaXOlVyLFQFYQwyBazZgrzrrG2+EfOUwuDS2xGiDIHU6
XHRfoWC0mH4pVMc7lJqiegSN1iu7z97udbiVV9jDhmu9LAWIt5fL2pSTSh9Kd911
A6dezsB8mkSZZd/fynstSNPz4C5UoSB1yHiXXEmjOEPGlOj9hDtMv1LPzliUG776
8wpjJlsvXldCnz/b8HCkay69pB1yEjsEcaeL31cNcuE0xyIIol5ftRH/VG3fcs5N
niFwxVEIuFrRIzu1JQc32R64xBkfLdrCX3CykSwaloNBR3IIxVPNAUYRNESYKU5a
2wVwmlBacCRA8NN/6QWGDcP7XMmyCEccizQKpeQ8ivucQRV54Z6j5sWlbM+i3i4S
Osa6aLmrHNQwkBkvCxcnffhLG3f9u0UNeIcTZyGL4iaoesdOzq5iTCazXvh9dStW
gjm6VKWrkOZSs0zU5t1saiMWce/r/82u4uyvC44YwEXrzp8dcOkq7Njftws0X5tB
JJBNcdwd/bHI0kRpwfhPCtkNoZyZhJTidxHA2Qr5hITeOG5eme3rbZnZBDlfxYHK
wUK2m2ufhL4sX1a7MDMQ73UJsm9zDRBcnidrzr8tWTKdZqf0AaN2U8Lq+k+QPpC4
LzVrAXY7fYigDGRq1kJVgd+mDmIs2pgbebBCSp4wMJ6vrkF7T/1rxPOsU+ZWMcs/
IVtDv8sEt6SReEgtOK3kVc75HmS296/wwNHBD7DLLl9CS6aRrPegKhNvht/5Qf2r
5Iu7u5bWUhWQYDmaIpv3k4r47Z4tRH6zb3oiLkqSCmSyrRRVVlL5db/fkud3nSY/
wKyE9mp52t2KJJgW9N6Va3o4Mb5UTweYP4VHAu0GrGt4N/RAOysaoTaDY6omLkef
zzzCx7bH6SOEJenRymBF7saOHBqmyjojQqZCm5Fw2AHZ8TDpYFp68futfEFC3w+b
NF15Pbq8ZIc4YyQ97op13zcvBK4tVOfAaNd8/GOy/kMZpQ4wspjL+XHtdGrfPe5K
D2vG6BRzduR3w5wY34gJrzU5Y2xLEYLF+IRkZMLaesgyKvTpLX1Y5QNVHjS56xpk
ibQigMDnmubQR44vbfYH1P3QDldynoQhUWDxSWq2mwAWpB9v6uFDFYfX/JEk3BV2
3kE6yshb/btbUvwe0/TJ3zcTWvzoRrElEenXa7fbkFchj+TrKvACMNPYXlyG7rR3
4dbB5GHhZi4rwf99GnU+uUYmi6tL/FGawbSjUK/zdXgVygwz1p1PPSMNWDepbMvH
4C5OJ+D/aMjfxfY5OkOlz5KvM9rR/eY4PdjS0vfPm/fK+AfPdZuWB1HxDAjYGSwq
6AxCHNv1HOKcanVzZ/eRTcHoWBgAFojIQgtMEJHkrmROt/kD0RXRQLd9QxmcdBNk
uILD4P1oC1ygQ4XtVblduYMqI3FhXtkRzrJskf1gHgAEPI+YNoYNBxFA3hhClswu
/lwEuB35Yh8TgiI/2n9UzP3kKDaLcLhxpzSVgE1Rp6HoaN0MA8kE+yQNHQ25h/SL
vzlMSybVcO/VHhAU7kTaAb9clXy3+DkjjeLoG9IKmcT/h/RF6GRcq5IlkwKBe9H0
NjplO4eD4aBLkopQSFp4/3GfPjaOcXEvYKpzPcZO0KYYNfIVL9WGn7LfuY16HKsg
UIr4WTRt0vuNXCH1ueszpRe2SXFg+YbvzCdhb10f9V/0+iq/uQiezGpcZmLqfYmk
RsDAXAn0HLJSE3uZ+DhzQDu2v0UH398MkyzM1aOViJGn/LKwU7M60UT6fXzse7Tp
xg4C6GYIMzMJCXfkSu4IY6LGS7s4c0TCY6W1S9naNyCGukEiFzvgkAr+so8kgD2b
CvoNX9lpO95+u49O1lhCQi+oLhPo+MjBUizWhsXt6YLFoQQBdt5r5hQY5W2/YsVu
v2H9dMqqrEGnWddNCcq0jnwUP92i4PfNiqIcLX76EYW6kBNTGAOryUw9OOa8AkKE
cKytOCK0IBEUC6V43QasSoB1LMSLhogi0lMrPSf1lK3M8Kmi/D/tvqrlmNGkZZHp
L0c2ETBFY14/JYIndlNOVSYUiulsHVcBhjuadlcDU2HuWVwCJoVH6B1GZkB3cb2x
50gB/ztiu9TVktYPvKgBNG45ZGXmWDcInTghtQRt7+MXhVlHcMGhpQfrPZIzXBGS
r5u3VzGHV7EgF/EoWJFUlcgyDWSqmlccCM6ypfk43R8Z94lxL1bxzrgMETBnbXq4
18SYPNTiQPVVLO4ntGMXnZLans067xy9kM9eVAyDPCerj784aipEQVe4EewxblRW
4uEkl2z1Wm4U0Lc+bcma9yQXp/IpWVxsvs+zXJfXSYrFUqY9KsddlWz+KC6B9CcG
uidP6iPVR3tfaiZnNyF/NnbHE1Dern+rGrDMVaDpvg7nCKd+NmXn+knUWsp4qrfG
OFz9SUostFIfJbf9JW8jAd4c5/0O2oaaAvp7ID9K8Iy6KdWpbWReG6R72zYbrIs0
/nZPH5vaJdBG5HEFq0bf4rGFjPtevmcNwqYJ5tXZ6SmKz4oSzyC7QlE+cA3a8A7+
mHHrvRiuzA7wZ94huwTjucjDeXfFZs2S1u6QvxjWTHKl/d3nu7RcGcRiz1aCm3J8
het+MMqM9ygDZkQQOqIH2RMlcpARIJ2oRUOIClDq9Ig/jGMewm7otCR4EArh1V3s
XaSjyGUM2snyypWJv8KF8KemxRLIg7IfXgk6Bz5uveQ/IjCNVg9AU0bDHi2D0dYO
yPXvVO3g+FoxXNaMZeqwKfxl0A+3z8d86HrN39gdjHZqH9GrviLtetck2iS53szQ
kI5mlsRw6clhDD8fTcv3k8IVthK5W3zI3aWdxY8/LTfYp1lbKrQRZMZ7CIKII1gH
LS92PLcN7m2ov8ipOiqwTlYm5hLvhpoLo87fJKoSt0k6L37lY4MV/XBENkotPLe7
Y6IeiKKMEs/zJrQTJjCEKEHlRfijOyjxeY7NgEXAIgCmqzIkxSqUg/L/48mUFB/9
qX4/KpaFrVYAttbbYJxt9Psc9W7mHHsEDXH68rzFdxPd56jc4BYi6/9Kch60josr
NQoGndSa/qv7/fPeNmrBDm3Fi9TSSMhrSSkfzdmSRFEERcNK2JaDOOrf7Kw8KiHR
UVzMYNzM8WPtjSuh7ZketBZVmcMDBd1eI6Rno5e9plnJwWfqefBjkFDZq6IIV/2o
uGXtGXbTMLQq/Dv3Pk4645nL05LHTNzZN81s5Se75ANsFvnj8/Nzln8ef1aBu997
Di+X7qJ0ODGxn9/2TYkxZ8CFtv1JHWU/joKBANnfyZ8shxVAU6GMiL5KAaswoM9O
dGSio5EavnnfbmV+U0mAHa5r69DTvCdsbRqNy5P1abwpeheGHtLB+GwgmtEQHB4d
J5O0zhyKSx9/nKrKepjKnGZ4akF6Aek67JQjo4znE33Z8kCGrUnDweVSuU3H/Qw+
ASOfbOoH+I56RpmazGG+cmXtBs+ChqGzt3SHW719CYOfDtNHOImelbnkPhM8I7fe
7tyG6tqscx7UJWrca3Nnk5go/NTR5gWQfMaGrTjkpLBwtgnkWnd+HbtHpAzak5TD
N8x/wVb29anYpZRfWY+g5n/F4zl9HFs2s9KZtTIH5FVCzbQnqwhId+xkUYCJv8v3
VhfSU59rbM0xVLYrYyEGyV4MSXXgllQ7OPgWCokTsEK7tvpnzyDFhNpD+5LINX0h
HwLxsoio+gM3KgqMGQ85H2P/Y5JVkeP3Eu+BniGqvdyXWYlT4xKBzGtjFBFGnEAg
i5AJkt8jx5KX2DTCUqn+6CjKNdoUPnASquHjYB2336582HiBTtqcqTSFIDkk8CLU
/M1FqI+dXAwQ5Y7gyxrTRsAFfu72z3UZzyjVSc31zacrblS7Nb7Ux/ETVYJcI7Rr
PJvNnmkH19ZjaOiWHUWIozpLHAyCj0qIAOxo+I/bjUsZmE3bX/4vwT6aautD2CG0
c/wFf3FXcmfvPUe7eOkzs6gPSKkzylguJIzHPL3nePVt/oheukmiTug981wsdtCO
/mX4B+gRT1nren9VExVKDku1x2USPXjExHeI8rEV1HTUOLjGb0w75iwGA2N1mpUx
2zFEjCl97sWdS4QayLsGqSnn9/61IHYGAQis8kmMxDCKhF/+n5K9r/M/9k3oK27O
doUQRUCd6aT9Dm/UJY5ttcepF4+5em9zuMJ+6qSaQJtvl3Bu6sZo7QuwkgombY5j
ai7a2wyQFdBiMI1KmgYpitoYGNaNaD3lHCUXq5VTTkRnGTeD9JPPUvrUseuX9pcc
zAzJUzXf9LRMRXosmiqvxJTVGlhz2Pp1jFXEi1r7Dnntta8C7U61NOFlu679LeiR
AV3mEscZkfNrsOhNMg1dL+PyfKwv4XUow5h9nmSaOpRPztk7HZ6QkJmG1kux8wZi
f8h2xzAucmUy2+90NdubpgOxFakgkyU5xGrFTSr2VgTuDr40HTXYSPYatugDzGaj
2UoQQA6k1zLSo1uG4Zm0T3CMVz4QU/ZPigJc2quSulnDLNryvT8C1dBEIvociSeB
3J8YGxLNdWmjmjrDxQ3seY39ZxbZssjvvHM/V0fAbhCPnwPgEqVPEzFDHh8+s0bj
BrjAPreba2tHPauljoaHEy3y3RmPNf/Zx1ZVWQzIN7ljyTZUHoX44PgqRWqWp4jB
MDhBOarj0wp42K6xxUOtmbZ44BSCousp/8qIJAVHCmWBHYh9Z8nqsGCLAx8eb/si
BQSY1J/gJf73L2RW7TNtqEWDzQ6AaeuzNY1Ja4pQCMexPTCeoM35SLfAQVT1YmHy
D2L+1UZxCGxGpoUMvuNFIJ0rix/Cg3Zl0vu0r3rsb6+RsdmvxN9ldVbfvRRa9mr9
XWSj/VjxjjG18ErPGaIzXmYTTSC1+EyrwXI/DIv0h/pEL5jhzNuW/FPSCsbbiQDl
ctJej+Urh4KFjIsSnbibCaj0aHD2FVCJ8XJ1ALvsw7OJpwGfU/9eDTS1t//Xt5is
0UqXlX/XG56FsdYBNDzxSFZVg0mUlNnwuQTlm5PGht3q//SQICX7eZxmAdHwiAVp
Ec3eY2IS8OZQuGrdQnyrJLt+c/txRWhwMKsGOxYt+cFFNuc8FTIyRZscR1+c41Gx
Ib3GkV0nT8NEGnDdaCK+JkTLg2nmnb7iSE8z6969MNScBvdTMwolhsZO/zomtjeq
35vNakwqunxeGjCXM97kUoxpiN5BhEYi/aDe32xM1kQypFw+NPQqHeX6d3PfPrI3
fsoRHGhIZ40eQomZU6daPRsSiODj6agbOtTNUxgDh8xN663T9IUVKXNz25Uw3+X/
6FN3C240IFOWgwxIAWyS9V2vo60XN8X6JnpWLbAG6bpArdBMUJ3daKuxBiFoQv8D
/lQ9U4MjBVForKwsJpydONoSvVbF2k6PdmLbjrMUNEX6l5X/NN5QHJ2sPqrhI2aF
9+lZQIozT7HPZ7zhcFt8fP95ud5GyGqA054xGrXQJY9tQyPAZRh0e3kfzzMMACA3
r88hamjcVhjN5usqkSFhE0VY+VABhKBEpo2cQo7R6Xdn+LN5ez8xEB6rnJFb6PLS
UmUdkAQ4AL/smAiAFjgQjWh2q0BZuXJkDbp815FrBhyMmH0FsFwCDnZ+cI/x4MO5
8DRyaGj/yvrPpz1IlsqAjqwWqejeM31QDXjEgTfLtvuHjDgxkZ/qWYzAyd36pDw/
j5w7wtyGXJBuXeNCvOSfUieWiO1dz9TAZf8okAKniIp3Y0XeVN5zmXhwEe1EYh07
KRC8SQ5TgokXW/PyFhEGQ2CLAF/yODC30t2QzS7PsqQb6R5CahxFG6g4MN9eUOrN
K9ENtpOfwMeLz5ZPjucL/QSkyp3fJzVzpISasoSfxyGLkRKZsISs7NklorFFSlXk
j88eXewq7FUIGFF6BM9VVQB0uk87+Iglx0RxLCV5H6M1Crs1/1PN8X4RP9wAtWch
IYLVy2wWjqcVYo1dYp8zKEuxsv2tzVTtcCNxYnsRN+8I/b97eeBaAaAQMuh8wH6i
9yti+p8PxrGtklREgM8r7KwadKOkgdcgBdqU9anpl8w86ezpaAHmaDXqPYfRMkeG
HwM1046YsA+7ZoZoFIf3x8Vrk8DRESL2Hcv672pkhuYNISWlFmBhwIvCgP8xmdUp
w2PQTCDaiqeeNq/sjrjD7sV5dQkx+d9+XGPzvnldZ9fhklrSH/PSqjCVV8aLbkhp
tcQjLFeadfvlrvA9YGtYf+HDK91x8b7ziEG2I/ftUo7ooHfVkiHGDqa8uCPajzT4
pHGb72ZCZQMXWC2z/ksx3bSzehOjMj4g5oZAabju1WzPGeb6tXCY6Cr77AcwaAEP
24mxzVLNu+G0HLqM400KR8NCm51aqMN6oo7Smi2a6pm0WFpHDSDQYToF1LWQ0XTX
Ur9untGVkf9O0M1MJ3cWUkUdOH4wCDwJxqzVSzTdct/gSRsJkokguRoOf+BCKSTt
O6uEGgkNPhX3NlRGoVRWZ2CtXEk/cfWPu89mYrMI7JrqJVa8c7q+cAy1AKcPVqBf
4osLdKjknSjkQzHYyS+dHnopR9xu1w46hJ3esN1H8oP62u9U+6rSMd3dRP+MKXbo
KQHhyN7rYy1fUTRGXMjkabY7RG5kANT7bSYVYaNU7zhoxpfeMzngNGoHhHJpX37G
jQBt2ma9sdoX4aNBFPhCoVkKbVlfMsb6NSQLjXTjfFGF1PG/4fk90DfPB38IvVm2
evGTrNDm24urtlYPJcC3AAIqkKBWC4Zr/pyOuqVhysYclMNA2iIUuXp37l1Yk4vH
WOoPnyK0vxDArhbmhe69Y/g0yWxx5PKM28a9y7R3uKslKnMU6UCy7CX4vezhpx5q
/tT/z0f4kvymr4oobRCAl/6+INfC2gaClrWahJXMZFWnbUAKumop3sOCJ++8jf2t
r5E0vDx4kaifoDbVbjMxpEINer9ErW5Fam+8iOQd2Yma1vstllYj9aI7vI4h6SLi
WPe6lYhPMXd5/dgpyqXGHkrRz937Esd+nZbVDVwcTlPlE7KJ+skAEL/2H9Q66B8h
PYI75WMhp6oj5/a6fOp/Kst5rvobgALVl4l8A/fGRuz+tdKmnoUvOF7TJfnROReg
QeJQduXI4wHpli6W8BFQo5oNS8inLhHP7PnOjAv9qulynCaEioFehQOHkcCjtqCS
r7httYPuwNYxo0qIVlVeEPdWtR5cJ07nH2kKGGluxWY8dDIRMHubPqPefMDy30Ev
3KbWxZ5VVPIf/Ar9C43NtqQwfg18W79KH8g4LMu1rKGppdPi0y+KbBN+nO80sbZZ
CqePTtgJESCNZgKSATp4ogeykThhQT2UPDUngtMLek4tm/BBitmgdm/eOVDmgHXp
VzRCbmmoD0d+U3Eru/inMkNlSTQYp8etrtQVaTC/+A+VdPUtQC0BQ4b7hMVPZAHn
ewURX1G3Y46N0SnTDocGfLaO4cbmhaZ3QS6+TerpmKbOV3CBVPaaf5FFUf+oWF6f
3MipJcTEAm94UZAsCCoUtjzGmdJx1Ic+o5Vkx+vZS7y5o+wz17GG8MkxKlroz0xh
irrgCxu7GS9G3D2saqPSofBy1FDFl+aSUoClK+WEZxfC1FHcfeBNzneldUf2knZ/
PKFf6MGli2/1Aw/wprEWm3wJBIUuKfgFXmAzc3/NVg/szWJC97szzVwypcqxWvj7
/26YSWgjR50RxtJRJ2PI2wOS4eMLvjY4e1aOLqMY9sTCcFCaeh2N2r9/+RQYuW1H
XOkTbDrL2PxTLyVnvAMr09J8Ur7S53FYUp/Uniz3dNcviFymQESOpKvQTtj5N91n
wKwN91Xhg201thxTQL/MqeBqTXuJoK5KFkV355kXkgneXZHm+7SjjFjjbKQB/IP+
5/fVR01jUIeCevHz1Plm9O5/Lq3kQG9QZH40dZBOwxKBmBrMvDLqPxISAdoQ2OYh
RTLajt9AvD1MylZ3hGqbZvRR75e0UzDI+jYh6D/SIwuOY/2fx6Pm6eoj81VpImRw
qfxpi/46sRV4RrtQaqwuNoMLJra1oWsSim6yABv9PWMHFtLXzfC32U2URu7Ge/KT
VKv13DWsgdfIWpZhXeexyRApSrIzseSOqArM5J3ux9myYfcUWYlrH60713ZD5hLx
zFRraMy17vMqBfna5mrU9D5VVu96aw2SySW8EZhsD6tR+rQzIguE6XTTQRLJ75iY
pnlww/ntrqAgfjh2iRCgXQkh0gWrfvCl6v4ySJoY/pgvXqTx1YdmkpbPsuaa5+ZR
htWbtjdjrh/F3uHVTHUqEDLYq1zAwdMrXxE9yM5W3k15iYPgMNeoK7ihNB08J48j
WVDe3NLZgm+s1UZn+ikWd+CR3qpKlx4VD6bh5Bj+FTTwmTA6ABLQXLKtycXMWMBx
eNvEj8csxFaVPceZrN5iNrVClRVIfrsVnrc9ZNb51xvHUOty1xtoOjzvzCBhqWyt
bfwzn5javkYSS6A7fSFTHSfI04agjNL1yM6uEvk/xUpm5mEKdSeKSE6iSHwZWqJw
2Mz4l2xL4lCadI8fHDvrQUezhUCXpZzWQeL3184DCraRBI12UHrIN79wy4pACktH
YcW4BSUtPKHugAdgMVGNXFFPHDj9g4laql8rbxSHpwEx1ZI+jebIvTX910MRUbAp
LDXWv638l5JsOdj4Xqr0APjV4Sz/l7L3UXqEwdNo3YyRI7Ve1djW/FHa8VttsJ8c
dqzPk96SWtOYf0nQ2P7cp339K0dPm6DS+1tR5bnP89nkgJgnf6ZTzazK3OkGi6mf
10rgeDyeGoUv8q7cdkrV7QbmxHbZ8yYEg0m/rGM0s6fQsmAwdGByArGzsuWFEvuK
+YBfGjc1u6PiRLTo5lr8yl+T6yBgQBmE1yhf/AljKl4WGb1i8k9B62SgJGps8Ns1
6Cy0/gSNjZ61bNDsZ6HnDWE5MGzQqohkIMLfSKGll92xQjqMRIqMDKz7q3Irt36B
oQtOJilHDoRBgSwE7UOdkmRerduCj91pRYxwXzNZMaYMappypskn+Pr9jyBgTtfk
iJSJx7gqAKki3y5Y6HTcVbSFWXzPguNIBo/v8QfgA3cC9Bn9uI3YDa/uRTB27ZCz
dsIckEnLQUYpwk1yyUEucb5P8HsjxR41GhLXNhRQ6+ZjNFTgezN7Z1BJiP1SbYy8
Y8YOpmqos8yrJNsHzG2SKdLRh02D2E6++xjU9tzhjUn0559kqKDKsj7LozbxvD+g
YVoXqH94qWdu1Cr7Zn+DYT+FtdEU7yRXLTacsV/WgAwEEcAQQ4vdrLyRmukIbdn5
v8dsyHC+Tkrs/AAjqQW5hxe+QbKlqWzfrur8Xoi9HE20FcV5mgry9JI2lmGAUsKE
T6lQagxuJSALOJ77GO6H6NNUA0vltVOchlZiGFRaIkbLpFY7n0LKkvbpG8NQOA2D
Ul5TnlexfqQ0UqpWk+NdUg8n9vu2PXsFRSazhdvOYx/TzM6NVqj8hA+xww/oMjlb
gdNc1Ape2QmSlurA2kQeAvEUm+KaSeTW1r2h6Yw69F9aeI1m36nBKNbGdiIPVGWb
DhcWnmb8yhSKbsF/NftWI2OJVqneZV1vsk00WLBE+R6BGv7I70rEwbkgGXcd9kKl
Ia8IAf5sF+R2Hm4Sq4fwXpT4qD6/LguwAL1D6V3wa34rYJwff/KOesidyEl6w/2C
qKch6XvUJ0ATTpMyJCPkJfJLVUliwiP/sUeoEy9FIRtCdI95xtsj6X6sNyz1CLWs
ZIMliQ5Uw08G3yTwXgOv1AFqWQKGVO6xd5GRH62aRr79f70069li6OlB0mIlLoPX
GY/ogkHOsaTuWaiyB5G9xTaEbZ3KqgsYLwB/4Z+h49YkzaOykPu1Iy7nx36yyd8o
Oxcg6VctYseeA2uzOJwW7FhhRJafRSiw6quqYMc5kIMpFYgEVPEMxqAbu9J85Pqe
EiJbB6J/1ftoazZXnCPWXwXeGlbjC6xlJpNTzWe4Rez/+2+N1TeY134Gd6JexhCO
uKpedE8kXyHq3bJFrxc9dR/PIIJEh7tNeNylfKoLfe/Vq0SpH0EnCGbEB+Ilsjsc
BBpZUsQMvsGY+Im0D2Ys2dyUUSwV0/4wDEbBL9F86RJRyHHXEXkw/3ujRTqbja/T
88I+XF6CEnqmlFCmCEHmKwxHyh9sig7vdtF6hD2qdbRzqxbjQNR4GTKBzPw4hm11
4QZTNVx6ofLbmVYUgPDTnEVl0VAa25jeYzbRt5QyakI3+OjNv1IwJwkzaKvcGIo2
7NzoCAwG3LJz2+7Ct4v6lCBHhXnoxQHQyeE1u2r/9ovZWSjwoBTO+mKFCx8rATZg
rhIG4LCVp2+P1VsI/C/vGMvPFdwBek8jcQdvngobNBIkeYXHg3uwIZkW2AHrNLdi
fJDFmXWWSaBdOVk0SEczVqS2w/538hGn4K7b6/eGBydsu4g9ImrGBBZdE0B4ZSLR
Bo/wD1Pi+7v4A9tSKPAypOHgf3aY/1uSPrvuaG/Z3wmL1zpB9zDnuoPSdXsWe3QY
97cCICejfHIwIX1XUIMpZFwLUcPIyXzQFoBjyElJnJ3bIdH2bbeq2WQYtfh8ZFgC
oYgNkmF5jTaXBzERyKoIorSsz3sG7wh4pk7DLEI7pYS7j/rV0DfdsnNsNPn7aHTx
0qT3HzE2DsVx/Kok/S3ww78GmcLnzu31VuU0zdoTQHr6RiGPaW7AQpHQV95qmjy0
G1Zpq8ca/s7MQxHhNvAK5ijRKJULMMkBNOVI58PJvK96R6Sw0n/WEvjiEP8pqgWB
GvFWOuWiG4H0pj2Ovv6tA4zuAlwiM64918tcstn6GccRYFUWwmBEfSVh1tzkSSUN
5X4BPdf9ajPPJAniRirJDhz4HcKx5FXf84u0qKMJevGj6QyZm4iaY2ovbP6QbSuX
hdPnTNv/MHzZiomcThLhPbkx+WlLr3V5YlZJadU5u8ilygMyrY1QzLZrNFhhtOir
9pTb9hcj4WkX2dkGEFGbE+kdMQ+7CCXPMoVK3q9zkuIiTJlhggagbwrcp8JLs9Pn
LdUCz9bIxJKmgnd+XUxwR5gIHzuAiEgubS2kYmDpa9DlsXgydFkpRExNRQyYUz9L
frT18tAqxMd8+6hDDoLd+Upl0r0ChoqceegWFdhfSSDv4YOebWCVKYCBkwuFA3cW
PUO6v7+AaCD0ncZCSpKK8Q69pm0b78OpfPxoq/5XY4sMickppqxIN1LtMehukioL
3819yucrWB7J5DnFG9aPaaGeaYJQKBebv/w2AdnHvMg4WxI7/1UauUeEcgYegRim
pweYP4S4INm3amEjhlKTURvcAFYxi058nksckM6eppsrdt5NruCehwuI6ePgCE7V
Yr4VusOGKQ3x3MDG341bne75borXo10NZ+vMe+aCKcw/mQAbrReChjNn2hrMauMf
5MivTEn7i/eIOV+1y9HZe0DiNPZ8YEF1BzMIHuCpBgwmiKAeD6vIhRUDqT8i9lx7
E37ekH7Id5jCt6KGrkuIPmLtHsFm9ceFBN8DKQA05vpTD0dWDLYYAol95rUAzgbl
JvpLJzHSDPY+YVlbQDen/G5U6SE+gxmPQkrC2AwAxBvKy/HJQlaG81O6o3LJQiFo
B/Tdnchm/0l1StsEfHyz+IdO/HUC6h7lszQD/GcF5xLzx//40pEqz1zneRbHC8qZ
HoSiPcyZo0KAE/f9qi+5Dc80jJx8mwJWcfJMa8i9hlzdkl87i2QVoZPn8z8pLomi
4ALfigdaAcU87etXq2nf+TygGkTw3JaaCKgaoAo8R384myLsfl+8KmRtYedtysGi
abiGAnnAeFnovPfmo4FIYtD+48MSQTfc3oNzH2egyQ44e+0CqUxIz2WfnaohDxf5
xsMLfv5aiyZ6/h1snd9KTJtTC5Q705tkxS7xYghsukLOlpPfL2RCFR+nPF7mkhB9
6+foGepnO905SP3E532xutrOSpzaBUoby8GZ8VvRCLkEJ0b1RBdFu99ESGiZMzrC
tJuwZsggHYuNS06FXWYc8TWslcXfjQs7NYHMIL/FbqiW2YB4CnU1sd0cmbQmodfV
TFVcMm0gW9YrLZGpig7mBh61FaOF0xLWr0XOMresj7xK6/iHpR5nM7CKIxgUTHXP
Wx0jIBnxguoqEQrMOfC2NaLtXe3TgT3zu/kUCnrtT6XRiqLZ/9Cy3IdwkRN2vWh1
n/90zAwhGD+1E9+8ES+zxMlbi5rBEkpAWGTkDeqb3wsPAE/s0KMcZlzDC9kmvRsc
Ts/AkHCl8W8fGMaEiBzEsjDl9BUQEWy/8Xj43+yJbr75DE/Xa+nV0zrg4ps8tqyZ
PxJ+DbDYTCsU44WZudN185ZRH6XfEX7yebB+d3lxGTG1nT1ZDcZy9N6EcLegs9Dx
ZQveDlOzCWSdS3g5lLFZjEa5f2Qve5c/kW4uhECKYZoBFkEX0uZAQaIwUp3+6g/e
qvD7q6FjaUit36NG8Fz0H2jSqGheANPMlQHRwQxMo/FXKx9vz3gdSwKZwAtsATM2
Nakb8Nk240C8XVukVCn08zcu63NPBm69mB9bLPDX3MsIu5bEVv5+9dileJDXQoX5
n08ZX78g7fGfjwH4f1k0ry/7MklhMxo/HJa0pIcQ2ZSfwRdTc/Sfa6/m5bcY0QUp
sJKgrrbUZ8ZwxbJoXv52SyHJmH3a6noP3WsNquOEaHYJoaWuDtUreuz7BEkSSb31
sbfk0VsmOvarDPEXFDQf1NvCjBBjFEiVQB2AxJniGX/XCfI9IBGcLBnRywTQcggp
wUauD2atjHvqEfy6ivd5HkMomuVZJrqZMJV8fMD/c9k56gfeYIUlQdeUN4kOq+Kq
MoUgA9LwHWU7piWi+jJR4r980R59CgE07zXYe5YR94VoVfu38fgBBtLiXwSM5hw6
ZkTU0/GKouOOHilhgKBwql1MXU2thqr5hsdVkjXhZS77kvekeYwhb2iN6Wgtx4EL
3H/amMYWDvILbW03bmtFYvo1PRXTQ2dkzTbTml4i6FCSSqJ1gffRBlrTSFRObRSO
AfBFp6mBOTf626tc5vyoqZ9goLX42hI/aykaJrrgnWI4rIibhPXqzu+J+Kcb0dYb
Njpe1q0l8eylQcZlkt9wMd8Q8a2+qaQf86nfbqMOdDuMjcgPt5WmusgLwzOAltZD
bM2+NQ9UYE2V43iNUbas6sShKYoF9+wilNFei8YcCaPUeGveiXD3l5F96YUQ+WMm
V0S8q++J+tm787Gv1fLXsbpUOBDo/jFrUyiqC5qJvdOMmDUSItpFVRjuiRUpfe49
n1uE875oTjuz7O5UQLHVa56HXvHWGff6ybosHbmyb8N4zmdVcZvECUhbSgqaPeXU
oMftzP0Su4mk8X0MuNDzno+oLGJQQgfEZkggRYlDMbrzDS8fxQr3+9mLYj5jD1bW
k++9LLbZrYE9wQ5LjrQHxAf/KUqABIc32GfVR5s7bf7NDQxhaNX950NrtHQe7Tsv
kOw7TdXG0hi3KrdR4VHIPMTcpqUn0cUbeDi+JInWoy6xXE76mk3FzU74JZTJmCKn
Tgxx9C25839yrDn6+wRoIvGjMYXakElhXsNSwSVBwOaJ3Na0CvMx4M4oZvtKfXzH
ePMAQUy387RBpfRI6NxNKezA9je2qXNTwt9NfJhSXijL+bpp+dl3K7urfDvgvFih
JKUUCi245Pk5iS+C998pia8aijZYr7PEFzYuEOwMykbOKH3v8PkfoPo5pHFjTXFN
xZdd95ZYFayWxJFpVgcVOigWESMWysMGu1IlE1EqOdQV+YsbpCQyxZ/TOmw0XpvK
d5qKgw9nXKr6ZZo9i0dMWZzTkAqu/Jvh0MZQjijs1/xCnzmr/rv00beHwSw9aWCK
pnMV4UPpXr/gS5+XWeIndm9jNxDapWCKg8sD9KaZGzL3w+zZavHSVAFRHAr/ywg4
4aJz++cC1mHPs54ElD2E4Cjp4gCWb33oNaFv4DJyCGsVi0H68svq80EgsX5eibQg
5bK+TJ9Q1lYmUPbPYkDI9OFs2T/y7oDyeMPwlJrFaCBbVQoXhTONKY3mN+9fpQ2E
BcmAsNAY3f+I+STNU4DtBrgpi0ydldQvYZj7sLyB5qOQCHLeKGE2gZh8hRkMxyUl
D3fXXIZGZ9c3djcZZQp8rpHDyAvcfihcq6sfzMlfSvKfZTIX8Jl8PizcCz0rivHT
6IyVGQG3frNgfJ6M1cr4EydN6SXWfMNyk0fIQ2aqlTqXKz4jQ0Nln6rbu53YOmyu
rTwywvFYDxqRf7j0z1ScHh3epVkrdckKbOpHhGQH1VOEeuIkEFu8iH6aRzymEmdW
W+n5TjYMKB+M4Lwp2UODYhJCs/K4cDr7psqDLSIrAjfGvXeFbeaTvCuAq65NczIo
TBMxtYaBEZtEDfmhW3N7NWI620mJycJ05fjH/kprt2VdqlTaAwWz6hY5cYSegKpX
SnlnoXz9Zr3xHn/SP7opc4HXJIagiFGrE9fOFTvd4mBNEvUjxH9cFKyQ5+KeuYHg
OD5nz3k5M99JQlRPWZP5SxDuBBqVNoEDzYnLt/VNIwuS+FVTc7j+JCF6kXr9znw6
i53o58fowE7mZMWlr+dzNxwxRcXpUy3xzX4ZVh8mkJBc23Y38jaod2U60D1YQl3N
2VIzxzdP0kxQc4ds69WzgKuYfWC8A+g6/MgCrbOOAV9XPZl5CKFm8RFgAgeNSpGs
8KGB/WUJ1u4DBXkl7n/cTaUyu0hLY0XDoYaPQ6b7b0nC9jI5lypQSp5Blg7uqsCb
N5pzPGzZVeEgTsICEYJKuemxQLSKAHa76zRpGbYr+bP0woU+qZD1NAd7CMnOrpA7
wMomuFFOIXZv2r56wqwDluAsy84lPqLGUF8Sqa/zG/Dhl3qZfH5+VyHHN+uErEr0
23CJwD1Ji9P/bYLFrTHjk5j28Y9VHMAubAm4sUeiAQ7bjSpS4EQel9RcKhRTCzPx
1cWbyfvx6dmyHLOlho5XDaAmfGMb1Wj1T/A4gvE6Au7lJNW7RKNkZA27zFo6B8Bp
UnrEXlbAnusMfZQ2+V85imsx+ZF/QO+oQrwbydMjn87mtE7DtxmnyymLiL5e1mNz
+mvsw4zZ8eoQaPCEMxvjHIT8P9NNJISdPs5VgH+HOApCC85I0qiSXzPJTl1VnDJL
el9B5QOXDklUTqxTkzL73G4DD5fZJjud1jwtW/6A5/HePfYOylUeRZ/9euPKrhJI
S5BkMSbKicR5DUrJH6WVUGu/fuc6PJVy/SE2a6LlzaQtw99IHu+KXcKarljzAsUV
l1i0QYejzZtH4iOP5Ig3ugiUq5r5ceLRZS8nGqeDetWhhWGmX1soJJK5B09x7yhu
hupUiiRxNl1nQfiR83+o3q96wsURCl2BMhpFYRbJjL7NBHyZxee55ymvc1KkpIAR
0RhNsehy38CeCkPNc8m3wvP2UuYVAC6lOjOx6EJnF08rVOqPPLz28c/WWboUqO7c
lYCbcLFlblMyp1DgeQQpdHfSmZC7SKb9DHN3TLkmXbW6ZqBQYu4XIAdNnZCryw58
3TpCXgzM/f+b8O553ZDzZdfxZghpiShs3RcfMNesCjYfvvY5CXzilVrkOy5fK+Xu
wjSFcRPyuWJgjsFommL/Eioj1cQ5nLaTy6v72Utfnscwgz8NP67UwnozrwnzP8O3
bHbFmvDW9Px03WeF2JDcuGugfCpagBx3Ei4kya1uNdJizf9dpDs8C1zGQs0nyoQR
n0yYRg468RwiYn2UJeFlT/ukzO6dwNj3iyzv3ctg2Yv69ubfPccFMZbIL2ZXp3EL
Us2dC0jkVzIJaLIDa3rbZ0zgZv02+zEoYCc6wcePGGHkaWa0wiD0u9kTFox7MLP2
xHciWCILjmo/wVea8wAtWZXJBCFLfAO7v55PDbmOSjMTzs7A2k6eU9KaGvEBU0o7
TajBlzx8MFPFztau0aO2pft222eQFaosB6VtnRTY07RaqZRfIRQ+isyGlqcQR0xo
2IFIuc4Bxwofct6qM22HBF7Azu5NQvsl1yjmuHAb03nLMCUlB29cG0tUMjGfm9ym
N0d6O4lgrCwwY5otpq4du/ux32rrkhMdypA9JAO2ZWTgibzMnZDJqdRZb6d5sa3h
qqXvqq09OIU34lFUwzH9BTCD8FJ+8Vb9iMrKzjgSceOcUjFWNYBh5fWvI7S3spZ0
sGrQBv3Vy+dcs0LP4Ijqg5rGUx15LzhIVI5DUu7Ho8sETutEnb2xq4OGuhKBmBQm
siycwlAHhZ/RGqQ2AauTVCEs4z4IId9fkoM8m5ka5C6FmnfenAb/UQc9Fg7Prhn3
YDP5UlrXWbiDIIBhtPRPdkeyQbtLG7ULMnO8WQUElryx/0DGiX5rX8EmASXxpWZW
DXCuUWNswdz7Kj+Na8/aHxO+TxpsT5HsUVE4KGVYduLZ042bJVovwt34sM10UWjq
WH1oyRyNNcD394RKNfqutJQaT2iunExPQxSwCR4RUyCf3drD/iHIIzEAaz6nNX5N
tdaOblTx8LcWYJmSCC0rH8mMtRWnUZ3NU7D51FdUI3Tn/dn3GogVfLLHBQNrLBND
Kqqu50JN0TvA3YGCbC2roRh8tCimqdSv3GYjDD15FDk6IwivWKqx80zSMPnL4Q8F
/f8/MgXq/5uvL+tAKxCFBjMJPvMImCj7QrCG2N3o/r6idBahyK+KDENtuqa9WFSE
rttPip51hCbEF0kfBwVupOa9KLAIbt66u/zHcv8dQ+tcnHrS3U9iF4L/SNOhGFPV
AECWAbRDNqi3/tHoVc1lBDA8n61BCKQirXguTO0/zn5yw1qsaVJl2kTuRHwQ+Iyy
q9lMPxkwzWwbw4zldA9ADZt4OtUjyrNn/ohhrKFUeRUwu1AM9ZCVA+JStSJLdwO9
bGkIU+ioZlX1X6syVSICH+ajUgmpzHk7NPGd/DG10Zc1+heRbrB+rqEwA2hhgQuF
iPZA77bkNRXX87gZZ3Fi2Ot8uRor/R/GLexwAvGMj1ii1vpnDyzSgz7i1pWEadul
lKxLKGfierVTnp//yswXqGOQfMCHAi7YCcpwxl2jf3zumnrKNjL0m4x1zPaVW5zb
Jb9SWWh5QVOYoX+KJAts7ciuvrgbbdGauCLcCjW87G5+CTBfXxp9umbuaDyQlIdZ
q82fmPgI8hFi7RhUXCPSSRzuMImLlJ5qREjP9PXd3q+kXsSIIV2vsi9B45dJfOQz
IUYsKUx1vqrrCVoJl8UxrhjmQLUwYAXGKMdaL629Geq5340SzdVJpYF+7S4gA3CD
rUcNIIdCdM7tFB55YxZ8nARxu0bbLFX+NszeqFJiW4n1CmOcoG/X0FH6qd+ajJbM
eFT2SEN4LnVT2oWfZE03duroUKQl+jiHrtNXdMf4eeXOtG7gttb1RxM16DtAiR7F
Dm1ta8h16kmfE9t1Uzqge0Cze+WX6OTO5ZRzo7oiWx0MBGSB2dR4pzOK2uSDO6Um
5SMudpGFKyNwKhiTY3tQ6YyVis7pWJW6A8cKk8fXwmE9jNpp86G+OuaEgVV/zupQ
vPOa7VTQWeHRN/wu6hPSdTz0ippzMNE2ZhtcLZpr7VYyDdSYUHi2XTp2I4L/E6BS
UTUmXaseQlq8cPkYvTEg77rYQocWO/arctXq23ppeSV03Eq2SL+N66A2jZS65QYC
hWurncvKbGWWJ6GnNl5z3kFDeI+4gW4quNE2Ps8R2jyNYoRXoVInHb+aC7MB1dsL
JcCAdF3Omtfo068cfBBU34yihPtDEKAMeP+UzaRFRX8BQ0OfqUuSB9xyfNoqPu72
vSaYHeAikViYG7MfC0INdsmJteQv8Fmm/rnmjwSDTQ6iAQVllG1wc9J45eymtW2i
1xVvFUh/+XcO00u2Z5HVH0ceUlrARnNNy7UdwZLOhiMBCecxHjnint7xZ/08vyWa
JDnmeLlcc7DO9xy7cWdyrGGCgIu6NRCJxA9Rbjm0lD7lRxzUF1Ef1sRbsqLHvokD
F2zHYTT1rhr/iI3afRKF6lZy0Q6Xqrut3DlT9i5+UZxmBmPq5Dyjtd0BuzxbQNOP
4L9V0msacWVT/dbNrXD8OM48qJLVrzT0vC2StBa9vAmPRy1UnG+4YpoOP+1zeTwd
e32ciPY/6f5Trog86Br1J9BWCvHFZvCvDXr/KK37YlI1WuKgS2O0RKdLgezOpSMs
ZSai5c2srUGhhvBtN/RWwec98GsyMBasr6xz5H987bXSI6gfPJa+cRADgQrteuef
88RhdDI2C5jZQixMbYfxPGNnIguYtiuzIdiqR5M8cnkvCHYwuLsGStvC+5Bq8hTF
M5apxx3OhVxEwVkTy5y1zzselJdtjSe/GlW19ZvTR39NDEEItSDTJYabpUSAGV0x
PkGxie3J89E5cMopawCoeNhIjprYgakAH1gEFY7uGGIcdULkPzau7lDIFDT2G+Qt
blsydUFFkkHP0g/hf2VaIIteNa2NFuWsxw2yVOsajZjNbKhvqVV/dzXYXBvMK1Za
hXSvvFW6wq+KzRKKTcd0B4o/MHXnJ+tW+jHrmWGSNc6KK3iTttrQuyDZ//Pcy7ua
8+7IumQEZsyPkTfYZLhukzrPhlJEWTMN6o+OpwSZvLFzglOY9teZpzGAxkY7zHXi
H9luok70/qCF/n0aRMQij61VuPPQiOzHVI4zf+RKzWaTFeqUi4IJvEVUu9zqrQso
yedAj8DT8GlNLmP22sgrxnznqCEBu3jHtRHOa4KQdJ7y0ptxGOogFOx9x73kmtyk
rKKVVEeKgBdv/o4pn903hrbFwQvGJim6W9kBSEeJT1PqjJl4Ac5siROXbqn0NcNi
qLMy6uG71E7HyTTLoRzwbNgLCBZeCxmm0QvhTvG6villfABnL0XwmKyZ7PnMfLLI
6FEjapTgg9aNFvxzOFL6CSdulZqWIV92KiNrwErCxbbDCYyrZItUwYz5pfMLp9zK
6BzU93bvZuGbMkeNZ3PmKekrrbXjArY+hDsWVp1YZtelHJeENvmK2DUrngtbM2G8
sE7HZ80QvMcjrh6Bw1tGjBmqnOAn8z/IjfdtyIC8tMQdQY00mzHpZi44GvgChw3o
5adnyFJdFwnz4cf7rTmKY5Tb8ocbfmdL4cR++6PVL8GFWnWChIq20o4JZpJvEDtQ
WAPzCCtvtdSFepbyrT7P4Ygxzup0UDa1kuOiQpoJJ9DqWwiT8dcwdNdkIYDliKiP
vZJygmPCdulQqa4CUnrXrMjo2yMXbVQO0B75BWmLyFIrZqKNYfB3Vvs+rbdqzPVo
DhIpWTFSkavVBhKQeyS0YRYIz1x9J3c/NgMLou8YV7V/Io0I3cyzLsW1xZSfnmFb
sSlD2g56p+0Ue7wI/ejz/wvyJxYPys+kRhc6t8Hh2AtFLf+86YB5HX9KQsE+WvqQ
NYhvV0lwbp14J3m6f0VKYKtH4/qmci+NuS50hpkVKhTAxLUPdsJTEk24X5TjziBF
DHasTOIqXXYgflYcWtvJqErt+O7xZVNWdgku0QsJw1yGU0T4rClY08iO4VH7sXaA
AhzfTBHuKZbTTAvxd5elwF/UFBu2+fw5idw+BB/MaSA9B/KcPKQd/PqnGNY8Bc0B
3qCz1KS9N59aBgkx+IyDSk7nDezg9YM2C/F92zzo9B+NCC9BGA6lSpFylUdjLQ1m
TzDNQCBb58QKix+OMtMlxU7tzDMjXElgNYv9eRx+FgtB4XctXGJF7J1oL0xC9Rvd
fNonF538ckDk9i4GTsAggeIVRTiDOOuDEXiYcdTBm3BWew9q7p5QuE344Ejvg436
3k+noVnbboc7SKBegfvOQSZ541qDzQiRMHjhEW+mTIvFFYSyCk9lTZ6T2tY66Sw4
Qm/piu5EbhRPIHJF0kNqMOmhs0Qa9++voiUAeIWH85m5cqR070PpFhlMuXK6TXQm
6a8G7hwg++NCr5U+A6iXyDpbaCo6oKF5o+f2rqm4SdKhZ1FWYF5+XkftHtlGj8nS
VRjRr5xaAEdJBJynhzSUFHEHEDZpZEnZ3U8Z02YIvdar49SagOp+ab4/BVrk7wU1
G1NrDQZG6CJt/6B+oQE7X24hVExpXnD/J+kTlOGfJuipp+VJuCHsNAfs+jkq8Ygz
Yn8CaL+2ru+eU/Ib8wxTMbxAadJ+yMvJ6Dy/Q9RPLTeSlL9aTSD7/HsADtk0QJHd
qIq2aOCAKoJcWXFVA5kig1axrzG0Y7ls7T/+F7YJhblh4REKVAeuubZrii8A2P0I
I2oZPgN+xYy2MkYydSM65HzcHJSs6OtOau0J/2HwD6iFQ8DAnet6xlptwnCt1jhl
S75uF3qyeSvp0GYsb7dnocZWonij6RvTh8S+jSXW7BemUcZ/C6Q1pwWpPYyqlMkK
w9SBSNHw4FQG9G1MgiYgUYFrrCOWr22R6jj6kbCrNB+f+SwsB99tiqvZ4KAJFItt
cRK21RbnS6bG7wuvTWorj97Jidrvs5xjLGJjMxmsPYcW/2wuU82fBtk4WAICpsuX
75PqHe9zas5Co5AXUO2yikWfadUNUQ6CdsswJ7VvNxFVjtZJuJfm4Zg9WZVaCM+v
Zu+kLmuEzGc/PKFQpnrnEYq9hsjZ1BM6fBdodlFCLckz+rD5T7ZX/OqrCOsI1LHp
mP1wUp70n3zYn7SYHRlACYBWT14Rn7fhiqH9t6wzbJb+Eh8hulpGQRwScM01+jeP
8n0ux4RNkEeo2V6L+8K/TUvoKzVKZ60mlYMqei9SVDGQKEtqhZIwaRjOQdk+LsrG
DqFrr2pmH7ibDlczMQ3hSnlUp9Vbk3MLkThmv8a5mAxM1Ztq1Yq6reL+GYzkDzj/
IEUSIYYIcPYqkBm8mcaPaP0j6SdnvfKCeeA47A7VR1S+ZwFznLcdLPmTfqrqDBsb
ojgwXgP4a4sZ3mmUOaGa7iFSESmrOi4xnNCGscTZvtnjZTz9KajzI2AsVmZE3QfE
x6ELogn2AxtI4AO1jDLADfGtGUnkWSXHE6PL3mp6N2sFtgNOsCjBpK3rb7ExerPk
aDEtWdKaqu3XtvYnVU3ivigRaXMBzEUAB/u5kOJQbp7Yvep6M9zfITQ3jeIiR3gq
6D20n8IZWhkN6G+qGVVYekAmlvRdPpYviEydVOD/EnUWRsmzfUayDMWXyO9FzN2B
IDVuRRkKuu768SPUJL/5wJkwNXPMHt7JOUijG/GYvjK0jmoYYHOg1UkFX+rqZM8q
OZvUVoQDbeD30AQhotlU4wDLH04mwRTRSRVBfNGLYTQuPLJxG/7X0lFoBu/dwuRi
v53Kreon2WR9L8rlHGoUVlygNuePygsQWyOTlGPDBEBgO2oKgL4Fe0zCMDfCmDMf
SAhq4o3CvRz4NRI7Oi4HsxIQyW+224NeuuG0zFfZ6G+oQSeqKHeVL+bpZGPf65zu
2kez1u+zRTAq4kb+977+oWHcU5Jtw7eWjM35A7eFzBrfCySwhD+6DleSPvu2wRWY
YcI2kyflXAd8qLrapPduEAJfxFwfVYh2bo6CqP38q0ELFDLPGsvZjs3SiPKo+tOg
wOlUNZ4yyqC0F1BFJTmqUYUE3eSIokv+vCz6YTOmDdvFyDFWvsH/327R8sCG1yK1
LwwY/aiQlQW34xrxEYLjp0809MH9uJ62qSIYE8hHJVDTqhA1n+D7AXfWe2JrgDGK
zm8g2tJTBVMLjxVv7iE2Al5JWfG5y/qi01pl83a+mJLOlXHduehj7TBf1pFYr0QC
QOM1nw6Lk7klfRUp9+hvqPmhAZvaOyngn2KpvVbQPH4//X5SB6nS+ZyugGr8gVX3
fXwIWEKwcmUfFlaD2X6KzYuDM2R0W+EHsqI7xk088O3K+gw/zws5wlOzLZHJX5mA
zyQkHRUanELb6BtZNGuYIAu7D9h1MmsJpNyomsXD8MFeNtOAm3ThkwNJwh+VQ6fa
JUTJgCvw1WVNHqZzJ9mPcSMgVf50tRoWSsAM2Wu/qXSu7DsjQ94Sryunr8sRX+3X
g4EBaHTblAvPlTsArnUXRnt98rLuvpPdTRUAtdL/qVNNqs+CLXwHtnBLvlKFM9Hw
gSi+zZbmXn4YCTihH/QD3Wqi7DxZTNbZx4u9rf8LV5daUT70fxwOU9ItDcbXRXtu
QHy5TAf4E2z+/Hl1lDmSzQUNBoNjyf5q15DbCVkGEDeIzT1wpIjhn8L8qVP2cYaR
TSOXYUPbVoeGIjLkLxhVeSYtkXsa0GcldUk1vJvKD7pSHp1TtmijyKLz5GUN3wX9
aA9jLxawY5Q3WdBZf0ZDCvU3TmPMw/uI5pdPsvXM0T6OyozHAnYT/XfInlNZdzWH
WFY1QTLbov7y6/QD+2sXUU5Hw7vRXzItGviIJG/R2dz8gPX5HcYFrIbjZGjVawqw
IhyAdkjbQFBpEvKDocvEU7a31RbChEgfaZprFgx6gvpsXhDxgSkf1yIkJoX3s4Pq
1hmp14T34Q4DzEKRvsVxlt5CT4xXRkNUEwPxUEMn+Wal37IjzdEVmteVnMttnMmW
dskH++tBoXvJPktR8+4UlDATSFLj/PUzsg57/ZNsEa6N6Kp1ik9Vfyi6DImQR026
kIeWb/aQTCFY8ddfIt0qJZsq2/esxPQCKnMi/6POEvRRFu6LnzCXRWlNkU47FBOn
0iTZUpnTqOhR8lhZ56q8TRBng7/45kIrboemtIwq6wMdHSKwiJ8ORw6hgVqWo6jp
blr46Ok5F2W+Gr7z8x1of8GBSqiE29tDExWWF+HS90lZyRQUWyidalux+OjGqr4O
hYcJ0Gy2N//V3L5mBf2PW5ScM6blcj3Rzi5Tk3TmtrnPCkrb/vvX0jkVzTHftqX1
9m96dZI3WUd5OsJgneFMpD3nwvC3Glm005NAfKEaDzYzwpy64MsDzHGcgPwAjVgj
GbXbGPtL+9YNIYwVkz7fkaZcwTw2DZvYtMNciDxrj6gRqd0XyydUkdDl0WzJt+Ol
V2++Xw3YCVd1l5gUlgXrZH4Wkp4s3hDV4xuK6Ynva43+cE096nSLN+qQ8bxD++eR
T0GOlLLvL6B+ZnaPC4k5Z4+NdLBJod+LzuMZeW4kLwMV6ahsz890zcuxAHTWcEzc
4hO35mKyN3pqFu+Cy78xZPs4o8ezQk93zquXYzs5sOet05OB0vwqKwV9J0YRI7Sb
Nzs9LTgcKrgx7r1/qHCTSOGVn75cZVPXB2gcXgi/ddMEsNDfgCYRuB2mVSa1xyq5
qux7XTkBMJPsbfae59+yMnLF2DYbWGiJ/nGE86TJ8Hh302epSSihFnDUwL0zLiwU
a5Gl/Ba0LAH0iaDMvojwYH90gveZhwJFF3ZpIvNiB5oL4ntYf3ol8R+TdOS5ZyU/
Yr5RLmjtn+i8/U8omXjzwr2RzScFbknqjPmViplebmn1tUwqPEU8X0e47XuJDDls
GS19Qu1N7ZdEBK2R4JgV8eaU55GGbWhkhqU195pkKRxTeVJidiaURxoHqo3D6uoc
3qkDzZRDevU5xgz4sA/QoytlsNSPxZot1JUs1kuKB4l1kTkcHRcS4oioyIWMC16P
MGxUo1iiuJrRXc/cY6ZjKVE5v2fId/I2U+6HmfrKHp5TnzAltibjYFUruxRURBr5
IBwKeuFYob+WbolMHlq7Z9/itqav/5JOa65bgWmm8er+4iOCxhsHWhoWOnNXMtKM
6ppyiLmNt1hmVJLVsHrdlIS/T5nbDqP0LsVuVJE0lNVCjryCyHa4pE6Zw+iBeHXw
tX1XhI3P2QfmLEEi4Qz+dDYQLXZTVZgtvuqrQkK2Ljjun18I1wdn6NzTP1iRKLPu
kAu27MvAegNRqM5Rh3NEZV/FeI6+sULNyaDysNCXBZFkVqWoIEGiTGBXz5gXLz/k
oS6Nb9jWS5LSf///Yegj/fOmfiLNaHnkG16LsPWi5TZqh29C6aznxx6r49tfgTFe
iCN+rCOYPhy128bb2FLrWUHKktG9eORudxlm7DarALFmDIlRGW1IHdnvuFtlWuF4
JPjPVpAO/elZqQCsUa/KzKylBHm4OzqbxGTLN2OXCgCcPmt9gmUWy/VK4QNHRRZ7
nUqIh75A9PttULQ2hgvaCRc1zvHa3w7xxOOkTp7z1DnURsqjhITPu9mdQrS+iHuS
dxa0puxouTu4CiYf1bTRcZd8imYLYPEZP9idmw5yuWd8wG9sVK8dZHTRp8HRXVG4
imMlw2d7sRpCa84uUeuxRIz2ZxratDzx5DEHLpJpxGjUptV8IULGtczLcx4TaRLw
tVyUTJFgTMGMkNO50QLRYY0gvsA0Y3KhppQPti1sIUf39+6DvPFuu6bWwGejsC3/
j5otcu6GUYzFcA6ra2/CiIivye9OxmM3qdPxRhG8pbGvP6O815Vr6ZuZjIJNYC45
yg9vtQCLJE3os5XAbXv5kVMqIbvvPoqDyT1+ONpWHOGY7gUdapgY7HqiZQK8Ws6v
hLyncRP/vaQjYMW/stNtbC3BMGz4gk6kcX5YRX1Fo5nE1pWMFZ5lc4mS3zGsWO+n
ma1bWwHTEvMgKPymd/T9PbNn5NY/Su2/ysnjr6NF0YWf2WtVZ/zVWEvApkn/ZqUw
TwBmS2EAFW3zJzYISZMICDJckck2r+XRxeo36ujCv8ws23wXiFqPhH7vs2u1LEy3
/iGSN12O5ouKL6TE5lzmTxX3ZosqT4iBqp2x0q3pLNCIi2iiZzdWsBxI1Z3UWYDz
hfOw012HOt6eSasvsVSYcCCda/vW+EP4MwLG7i61eW85mAwIh2BmbcRTYxarxHQg
P0TP9xsiKdKdboXhONwY10M6CXNaMAX+xFJrtivxPo78ZbnCwkcvsIyxE6hLkNE4
DAquZmQOQ5ysUzcZ2DJzKReTmhWj53ELuIVjqtSyWUOQ8Jdkgv9E6wHOYG2DIzft
zmJkkKzEexSiwdOsqgWLmt53TISxp6S1iHLXYdfnKyAEiyoEHdukpKmuCqqdJs0B
0C5ym1y9FO5LSgFI07Cnq8L9vXkv7CneYxnVEHhMMkopdGUja5pOWLtED+DuTkAw
17zCNWRx3ifv3J1+ZODu+PRaAQbqs1eHX8Edb4jiYeLmlMmrQ8rXr21QXph168vr
yYqo7eq7iXLhsZCTpkaXmEZgRmrNEQVP8U8C8wsAp2ceu9czp+wln+lzeDsKgPj3
2xk+Dpn/iAYlK+a+rHYHGog8GmYwCDlm2eSglXPHKyMjpyQIKndJn1ejRfUcEinL
ZQmM1LQ6o61KeZoTfD1IJi+TZiYOPqJshyCVq8fNlX0+C+4GDOPP1gjqtVmHiAfl
Xati4mlAeBh/2XVgd1sGgUVlBa2NWWpHiv3d67BZ8V7CewQj5gXmFfLJgbGcjcn7
yF+F51fWohOPMcKcqr540LZpKq9Le+IIBLpmFOlHLnZdzJit/67vYSWP5cfpANSg
rmwYmJZAFxG1m/7F/DRUksNAyy19NF3f0HeJgYZp1ppfHL0siVARNKwnAiyMcAST
/rhD7LQkLWLR9MhIeSqralTD2rmbRNzB++sSIskynwZ+e4OD1VcJFhg5EY2CAPMa
hkdRN8rH87ZVtI8LyfcVTHtIxW7IanL6suZM9AJunej82nBPNgsHJbV0CkOC5tV7
e6Yds19g6Ls6V5ZkZ0szRFqZa6jcJ8dmYKjcZ+cgT3XAXMPkB1Z8IPkyh8AyK5NV
QfDBvxWqTjcCvPYZhvm0R/Ra/39tGoEiv/Ht7LTFcPfd2GE7w8/wMfBAuxjhPXeS
gSw0FdEG8MDAkE0AYZ2OM2GRh0nlqtmPu0xIxpFJldcL9JrDBCo3tqWav37+Uu2m
oy2cjFuHkd6IH0frK9Y7+upe2zoDFzwUkTSg68UuyxT37MdnkoEcNFdJm7Mpsote
7Acug65tivV1JJRwBZjccdZNsxsJBhhATgeMHiCu/PMxnv4wplp5MXYcthMw/lpX
OCHHxBrDrjkAVQcRztUdQEJUA6JoeNVINSh9uSefLw3C0d1X1qOIqtChKbulQaSd
lPc+Q9gOkfVniP3gl20SaD3e8gcU5P3jV+myc2I77ewefTX9nVqzxY3ojZHvYv7l
dBQc5cosNDCZworBml5VFfND3TaPUiV7p1Rbw18MW90Je5mtJxP9ygOGQd00iPTA
HPKHxUROWg6kqPw3W9GiinW9W4algtm2hPPV1fk8ddJZjhIPWL04WeZ7XyHkc/oP
6Nj+fGCE7Ml5NKlGtLlgwRTjki5hzcNVKRRWmv+NX9i2KnhVj1Y8UZbVrus0f+ht
cxcuak785JtNnC/d6QJMwbVSto+OniTVmVnu1qYvNPbmGbHZnrjvxJKCZlVcm9mF
Hae4Z7faKzlGCwBMT3yLSAD71xoD5uk2dmE9QXBV5Xp1ajoNGObCGRWr9NTMVz+l
XRfXe1cucdjZMubZljAI9Ju6OhYwrF7OrdMZ9CORCX/m3mKF9CeFTuviY+L/Ce+W
07LsJhtXp/cGq6/meRPBd7Y3h6S2a1qVMUnoB2L/HxJjJVpGz5Y/1c9BXi5QnAmp
Wm3gYWrErP0ijLv6g5VRCD2LVqk8ixAAbBi7JViwyotlbNt+T1oYdIY9vMW5ASwv
LBbTLazlARHI5ZiKognSGCDhsk0bnJzZwUFzLb2CZhDTfLwT1bRmAotXR0DxqIrc
3p7U/36OgPQWRIOqpF4Pi4Z8DWXruSJ2u9VVO1EHLrtWDYRw4I4zeRELxMyg3jkz
RsMx15UXDVf/BfaFYeGac9IqVil0x/KO58SEhMWxkrnq82mvc9Cke8PDwY1pLZII
en7gqWPQL1BFZrfHhR9+8/XUtKHBJA49J7/LuRl0qUpHtpSNDR0lNYFE4H/NaFlA
/PrI++pkkC34Q/6mIt/nj0tvlxO65S/DGXZPdZiuaF6kvv9hy/OnPYLjbQc/+1Ec
GS4Jf6BeNTsIFaKQKRWDp+P6XZcFImUF6R7CEtevbI5VjKAMmrECmu/xnhthX3Xy
3YvzXELcO3FEIa/12z2rNSaHRUOcPUM+52OP3ZE5MDmtLIqLVvd0FtvW5Gy5eEqv
AtlKPzK0C9eoTPNq8WDLTJ7KJj4qBMcmSz/TPHwtxQJWRCD9W7+Gs/bO/z2l2c1q
tIRwKkVknXEzaEfG+8siel/MflVUTjFTXzVdUZs7+BhUK3T7nDpcN0QQoA0DiIKZ
HtubBQ4Eb0po103eXDRyOqqV7e/G1c275B98Bb3Jaj3cqqNyNpB4qgFrM9JWTy8B
LUc3iiNXlcWhwdY18GXHxmGqa5d64aSetLhf7oE7kW/NeJIjRHJ00qP7Tcu7R0+Y
xM1ocH0fgxxRYr/+W9OmLGnQ5amdGetk4FoG+Q94lqKR/h9HXTElsO60Imq0qADH
q5T7eqntRgJMTvBySaboJYxZgzu8QWl6DdV91QUP0kiIaPwxQv+k92/nS4eGm0OZ
7aPqRPkl2xA+3rWcgCcC+EzTDhxpo/y8tUxiNZp6Xz9ks3xdNQH73yhPPAkl5Yqn
Qt2gyMuQUh/YjRoeooei9wePfjoA5tmjBPU4Bzn2KQT8j8+a6ooYeR6EDjOO1adu
G6nkrwI3KkQ8nqd/9oAS4eW3YZWNiSXj7xMNXOMHY5tbTyV4+3JQXseQLUNVNhT9
OLS3rYGWC69p2tjKQ7FAnUuI9yikPV5B9N5zI74k+G25zXLmpXuEFUZAEtKuf+A5
I2DkPe1B+f5OAWTux4tueEJBLmBajypiOVY0KBKH90obMRoQAKMVCYEnnOyCaoOm
oE9vUxoC1slHo4MQK7F050JRjffUtL8/CNBpzIQ/qTUVNFi2+ZQiHnixFefPHEHv
5nRUhCwK9zbL+rQb8CUrXY8ctUs7K4OkPnrid0I+pE5UJJwmhdXeA1fP1TTnxgWr
NSvf+Bt3deWhVgIgwbfVEYc8LwyOALg47Ax42fRRcDgV65FqqluYRCublcMQ35tl
IhR3vuiQe97ZZPD9rk0fRtNt4rQl7DJ7Ln+kF3rkMSAc5tEvt6cL6u2DwkTtBUup
mqrRJuiih0XibCDc7LaUmlOrRboAcjKfuUHiRIR+L3AhYeoJepCC95naOhXrtwJ2
mUmHDdAPQiu6wBOa0sqEdNltbIwsy3XeBPPCuIldd0gail2OCJMkk5PaWE1aMJTP
ovaUYk+x8lOU/EeafvDCNywFjtV1CA2nb71IhQfiyTidQHs6MBpalA7MREMqmfNj
22A1QbLmuni2WZTdHoZdclpZthugpghN/1L9HQMvqxf0Ss0ewGWu7QTZ+fxhGZkV
ENJ1ecJ0CVq/CCogA/qE9B/FvOZAXUvkM+vOSV2MdvKgBrKwdY9NbGR0JCurreRO
0CEuiR+pcH+6eXDdSMOjupAfVKmS95X/zpqSAabXv7kO/oD17R5ohpmow+okcvhY
UCi3ehgkk+dotyvw8nPLuPTh0w2AgbWPilu4/Ze1136BI9JqsHSVb8eVaKO0k2K4
MnxYCxYfftbbQ4iGHgFAsX7+3hgC845qqTycVRzkezWe/E/20GP3Vbc2XYyjowC9
34eLqaJYu8tkXtwFx4KvKyZkx4/YcFepYklnaHah9d6dfdOaWY8OPPzCYZboU+GN
ZbrE060EWvWNxctrLpD1OvmnJEEN7gmtwjIhLdOIwss5Duwlfpox0YUS2XA6MGTO
e25zKV66i0MgSWnZiw2w0kuiTf2+ifl4bUqYr2u78sAr+eymJpCS5uvfZuKsJGuI
z4Q6G/URrfI6t+CKP4nsVbwMIYoYTCMXltif5692pfX6RWg31dcJhPTXfaPDoGsn
+Etvt/FcqpfDZ4jexi511vVkEU32CnYnIpGP2L3xCld6QQf0CV+gUrux6aaLijly
DiNKWPEYYxrjwHIY/vlnLSnkNbbi8FAAmz3Xi8k2z7NGgqc1IMDgGFaMXh38WoFC
7IqmeOy33Au78EgKIDSNllZL/bRX91ubCCEnUqP3AldGdfwrPz6lyq2YNqimvkhS
UToxG8AqnhZg4SNxG6/DIjuSqF9ild+vdJ5xnKCNpT9d2GQC7wg1VN1QtB5UV8+O
XzJT5hXrKVH8ftA/Q8vxSAcpmEPS2aI2aUwazglva/V1N/77Q4IhzygRVY7Hq/9+
nMG2e1PMRL6xWX0RfCEI5N2iRUR8+m4zrcnPylyA4lDxwr2Vj7t816rmUStQLl9B
4CyhwaotsyjR+KA2pvydA+j07TG413PYbI/Qgrz7XsPR7Y6qls/cjyXwKtq+nPuq
Glh95n+RWSOxIJP3B2rfObDLXopu7ZhHzix8/SLUg8ApD5uatJNuxtb8zQ0bpRwv
WdLNBZw6U0ld1nzZiC0ubir07BNQ5fEjo5rk4C624PJYPySUWiNEgdLo/bc6uFI7
NjyX0Vg9Dv7y25TryjxAG+ltKLfFpYFtGzuReRKiADeJ4jSolklKYhfYqx+FVMgj
2z7yERpf+qVyZxyjhCTZajQRETvU4mKD1uj1qW6l7neccAWKaPWDE4XVeT3w8GQ6
HFxSStlTu6FndaFuICLWfITzS2jpRrFNRD0CXzZEtxGhmswMYZnJ59HE5gGPoVnn
1OIcDGENyCBO81hQJQq0hhJ1loh8hiKigKEvWRb/Q8LQ/09VM5HmemGDMG6hRsuf
HDvw/KiIKepE964UImR/ki92RPtGXNiKbqa5G+yYBZCf7u27Ol0Vm/Uo6wjnfgFr
+4toj15/UAGpOYzGOpw4E+Z5CF+kLskLbJ48tTidVsLlPsbjMJ0qUOefCW0ib21a
X/AXhyBsTKAawMtrdyR3+ECShqWFJSpimJiolyxZWp4H+Eq7unFltLTRnjnNy8S7
VDCYld1YJEAV72V0pDRNBbrO/Beu/y6LSxAAC68A+h44pbQTCFVH5ZWnh/W52mdI
x6hz2gPS1kySNwBoVnTJeliOVPgtw/hVkxsL3HBZBwAG2NQksuSffgMs1f5JkOPb
WHLN1By1ppb5N+pUnTQ+9KPHEXLgRoPKcBrYfM2TxuR0jF9bCIv5xR9QJG4LOkAS
Sz57JRI1Ppdo602QaIY5q5Tm0b4JEoivNk9/MDSaVFQrc2Z+3G/8vymO8jyAhS2q
ojD2k596CzAv7Tzs4Cudnizhkc66BYeeHevySsMpIoBvydboG3Mr8SAWGfECapAn
e6xnzY8JUx9qUnE/V6srPhAWkxQwrgvMoLoynnGSi/fgxp/Q4YR/z8mAuY1PCt7x
KaeQ5mcVAn13lSg3r2hMrt5DGbBcnrSNsMhdfgQJLhm+ZPJmLE8ebfmepSv37kjt
dtROvGUu2pAD8uH4Un2JiYIwZVde9SEa74yMVhl0sCTt/XlrA3qKSyelkFadMqLO
pxWQ/NkMCMIMzPbg3GsOJLTpjZ2cQ87sxTP3ERblU7E8o6k2xLdnEB+Ikn+X5E/6
Knni7ia75LurNM+fbGbarQQydhAo1na8hfukwUCwm3KrVkvK1jozAD6Rp5SEqOL8
gbS+pIoWiAckY5QmcoIRQ6ihTwiicAVI4LsfzCxAmLEmL9XsboWyauL7/YpbWgJ/
VE1SW/4GRBd3KBUp++MTTswQZn9C3eKq+euJTgb8ZJPfsv3nNb7wqFEvO0t2IlBv
t6exDjMYd/VC9JYKYKBKDOy4ahMik08f6FUHjehRNGZ71G3GtwgdLM+CNznjTzyF
sZAGEC80goloVsSmwbKMdSKSVXAaDveb26HYCsivXLIbwa4RNMxlxUYsJLz1hYVM
K57Eow7KWVQtr0dQse5qoPG+eo1f1paeJg1zlbOiNFhWiwmBUQh15nM7ZB3DTWbL
doTzQf8QGZxLXzm7HVPmeY3fozIC/ZQotPFtG9e4orJ2fKW4cJ+/f6r6fk+OdWtB
+QsAVxjXA85AYO2QnCCVK//xHtfLOGKFODMI9uSNoWVRicLUbx9p7k10iFQsuBt6
K2Obgdl3aOKxfvlD/QP10fbf1MoMV+VnpFBqoSGBU7E6C6SZYAsCUxWisZxQckBr
P3zILyV+zE2FMhUkM2dBwSQSZUjmAOKNIy11nTr21csqlUU4N5//6bD2ZiWs/DMe
wuhQsZ5WbpHKrmO/VaeAgIbOEVV6iOYuqLg4OaX0Zbxm7lJUEm+gGjKyXt/Yg+xg
Xu08quBPlg42PMt9iShI/YsjyQVgeherEwE05cFZLWBNNe48GTOnqdxOaC2Pa+ML
HiXjNQHyImvC+k6hW6Kos4vtzPMtJRc44TaI9hjvrWVtWu06ESOZHPtbNlKpqRSh
Aq/npOLrU1xwpQ4j7bwZB7XYqtvvndFbCjpQb2YmTUkIho4In/alS8w8lJDPqS1a
255mb+xMgeFIp9fJjJuVBjmbEAK6Rgkn+RK6d61BsuGDoewZYFw99khzV8HJqWNd
OwnzycOw+QZd5qze3WV4UlYNxfepcXWrES8W1QMoNQHR80FnNMDKFeYD9d4ugi3X
c6qIVhST/wCsNnjq+Q3uvi36QfadephFjQVJ9SODPQKemrds6dU+zkO+8uLh/woL
2B5NAdItnfB4Yb0iTVSjDmtDYDSKmgHk2wUXO3zpDjGCDPQWP4F4Tw0JkfBjYglP
pOzJAiNvoiYyomSew6BLpU+Y7/McGIRT0oJVE4Y8Qejpl2TPBw4auhn7sQLlLLRx
UtdRRwHZTHh3/XQ0oDsFj+7YGOvXQfmGe7+40KFRX6YWDIvZ+b/g4ydLTx+rJ6xQ
4/o5z/QUwTWMFBw8iMfpzslsBwo3nxCxvA6Mrko6cZWw8XRA6Te12xdepsjtK3Fy
2fh7crQcul1kpRqb+Ht5ZtCHdbciiCqOEey79OlfPAtvOQNR+7PuFc+yQWAsHbuF
nCi9vyn5F9mVIZnqb4hD+WzpL/BLP7oPYAAH/sRMHSA0jeDOBtksLr7tklarTEpw
AnMtKJ1pXP9CgFUMNHT/YhzS64YlhRSntwBj3b1TnYyIsoJ4rKEI2KymVMkfG4km
1Sy0PW3uDxM3Ol+wEy4Iww17ovXN6OosjwBoSpLo8w/5QeFY8If+46v3hTcKVMlb
5JWnSKLr5EOwAzXL6gAmkK9QRig/70K9QtH241hhkwuk2j0SMsnQolH+ARwV5yAD
srsK8rMWpSDtX1WaQJo41eUatvlygV9owDKARdme7RjfH1yCx2iRyNgug/xrP4Q5
kFD7qlKvjmwMSBFJaSOMzKiSmg/uR9SXY3lXCbSgTzHxVy5cRAGQIr6WbMOE+VO8
uQYxT7PkVKI4TIgfqwFsTK7e4FZgvQrH1Qu2HtBOL61xb+8WFi1P9XbTRrFam0sS
M3KltcahExen8OAIKCHvJbbTx2+dbv/cyWbBfeQQxXhpStACkN0yabbpEENs4LV9
2keXO4AeydYZjEiDHQuCw/4Ck9jVGxaPK0K0YMR2tufHX+3SDTDM7ZHoUxjLt+kk
MJdcAcVuadCNmah266VD6LOXUM3PjsUZi6SmjTq9+Sn6qwRRjRcncTjUxYCEUYK4
bYvAE1dmC/jQoNH2Vgj8/lYdLdnSas/OfauDHM2vRNIFmoByLDjVK+teNldArUbG
GV80XHRaN5MsLgm6bU+wIpoFWduyzXBvFLw7vJYWJ6Ulwrc0A/Nzz6wvv5iLUIwF
P+8/f/sdOO6zev7qLGUVfqiRiIDDse9xMcJH8fneHhVvAZCak+JLTUD5i2+47Hd8
Ta/SToj51cakLjLYKZkOFS++QdTYBLONKEI85U6kLC4AYpyczdL1k9J1g3yliz6C
3XgETrAqimEJII9M6lqGNttu5dNjNS3lOsfq/U6zkdNDuXK2A22pcqTi8I9LTaNj
ZwNXoODWKux1gA6UtG5HS525ePkMpw7Q5PlXW5C6ratGiIA3m4U9bVprqoX7RjBK
Cz2xjCwssRy5lCyMxKwyVK4kwPK20z05UJQKhIrlBdN/tMzMZ1w9LrQs7dw93Kyw
OIRtB21uAKoNtgRrpbMAMspHATYQ5FQP8oQfroekNy/xAs6pkRPC9MI49QPtzzho
r8Co3pMCSKWsSyLsaMMQ2XEcCuk7AQubOG1VhGbg1yQqJmn4emISu/NyEjd2+/SW
Q7ODV3D0FhrC6wLhoWwrO/tbX5zsRORL+Shgd9IRMPPz73i7XUmoB3MStpBX7YnV
3qLAHfnIJX7U9e1orb2WwImh5bRVWeNNb+4SLTCtscmn4aB1X19eWpRh6TPoBWph
Zl1iGdjve17FLyw1iLUeHScMzCF0qmD5qHmopI8lvhDGuorZ6HQQ7A1qlDUJwsk2
ZiNHVUT3hpskn6dM4X+4cyEIB3HnzPAcCGIVFQteozbGPCusKfesuSjfDwUEAm2T
3LOki8l5SH0yeU8z+HSyFx1mWMBz/38KCvo2mpeTt8OWKMmTq9P15RJ6EzsW1M3/
P6TAseDUTNaU74pNy4mEdgwkHBcOyAtlVdEsuI9YpXXRU7+fVB9Xgivzr+U3GmzF
MFhxJ7z+13UDbKQi5GBNwjmgrwQUHpGAfrbV+Dwd6iajblOl4uWvlb/QITwyO7S8
ZeEnW8IbHt43rRveOm7s6LbVWDx7nJ7oP9kzKl/LQb3qpjxjMak6wfPM0Hqu4gWW
eWoITIetGaOBojVkbJjWGn6hxz2dvXemIcjVLDUKrKaqo75XP+P29Ldcqw40OYUN
JoKFHoZY/3WpGLDPR9ZIVy6Jz7YpgKU4NgUsjVZWN9wdPJrm7l38SoL5LcjUZ+yM
WunUsit/CkC62upNA+uKY2Wa46oK3MRiXPOqBVKyWB7e3/PnpWYQg2pLuEEQyekm
8yK6ouQpqI5ERNbRN99UWQZoNnUBqkHO6ljogcMXIZQR6mS1d56b37W98WDDyc0g
k8VRWj0topSbnRU4VkRnG0wM3sd6yD6b/g5+ouPk8mfXf9uWerO70AFAShNIqDee
gP0vOgRxZcmhEmE/jOUMXAyqxR+ydSmVpQsSnkkoZGDa60k7fShkd+LPMwga9dP9
IhUwCCwVmm9TzkNa4Nh++7JgHOMpkz3OJvpmwuMbQps5dhludwRNHaWF5sOp2vuL
s8IEZpDLi8AFtajK0I4Sei6uLe3BHRGc2pflAEGZDxnWfkpGcfGmsRHjPjdt4ium
+6hu0qbj2I6lmn8rLsN1yqtHA8TkzXFjQqiRjCUS9EmiYy7dkFiwL6HLOU+V9GHk
ZXX1X1zsdJNUAvI0aSp8md427k2ilqpL0f37zS9gmu3EjQodltpDESqx8QlhElTr
VxrPNixa3XExOrCLuuqHL2sYzIcKJKIK9Ua7JkKf+qP+1PwzXsanTpw2T7cO6ajC
/kx7K58ZNfJOj+ViPkpYDOpOFBGljk/SkbFcjAPbwxyKAQgNkveCA4cMCE2BaWuy
kvhdXXu9AkouNftdXofl7q4lkcoXYczkL0WO3b1yT/JdxDGhfKNYHZSsMcgntOU+
WNXTj0PtKkc1+6zIyJDEG3ZyTZmhGdL6U+ddUYzN5aoOnskEd55Gjy3j8JVBY9m4
0YWOE5CihxVbQ/4nUdJcUHjYEm663bzDhxKrmSDYulOWDlHwBHAFvf+i0YGZ68oR
stGx1R3peSF/o8bGe/Xp7WwK/P1CJh24a0DujV7ST6O5dM6tidJj62/0DPCn28Kr
a9DDo11F8VlNA/3f392wt3KxUxWeLjKslic7GIv2jsdvU5pqs20EMi0Z/TNIPe+v
M2hE/uDXEa2U0oelNVMVbLceeYdVWMvxE6EILmkr6VH5GH4ty50BeBBd2j9kVsC6
UwfuGIJv1MT1l1aegYdY60XpYbOVL17sbjdw6KOnykybeRwh14toH0kMUnrNvJnb
sA0MjR6Kl7fFF0p5ETz+BXq5tqgELYFuWSpx0PSS/6JZ0nHXMPTHrtxjXo492dLG
Q0AnM2hEnkuI8cQENT3NfRB/Ax86eutvGFPBUtX0Pf4RlxrOR2qQoUaZDXO12n08
1sVCTpzWmIMpbujfyi51oi2ReNFnynuRXpIb6m0zoou+D4At49fro3oJs8Jlqxwb
yfnBH5mCExaShXtdZ32RIkLmNl0ksrEjIgKgN294dwxmQPV2E2UQ+Ey5v/tvJPn4
0C7qbkds+FiOf6ZBoMsqM8bcP8SPjpf+XE/bp5JbGcaXR2YGaNXe+93nH87jmM0+
/PSdpfX+kZJH6Ue682IT8ObE3O4fxmLhYZY0GIod5j1ePCBd5gKUQil8MyYrjYt0
zDSDddBP0XeI16WvznixjL3xtsKvvNdhv37nJSrCNoO57Qsf8RHFDNu+AlmCJBzu
Q0CSglVuEndnPCg8QCmVxlos9X6phfC4GTpjtL/QYa494D5l/5RsLiUJnTpyR9JT
j0dANmx/qm/7twKWSNIWszEXILlUngLSoAh4GQaRC0v3i+KUXwfKY/CKnL0C8K6u
89agr+eKrvIaTg4j/s2gGe2Z7XSrFjHn4khYJhpqPnsRjqKwDCWMKw3KGGGbyC8r
bd06A4CwmbD3EUCjFJmbeyG0GqZBEXBMe143jzKkL9xobY0yhYTQLZTfXi45ikis
YTi206tj+Jy0F5nMCRap/1Hqpv2qYYSVsxye5CChhN0qLOtyFHE1wCVDetYwPJEe
rCr3Mh7c7E3dnQU+pUhJVBetd+e+tr43IYEPiYtHOo//98VvAjZYeBKhUkhl5O+p
MTkBZmRJ73b6OknpYMYAHHrVi/j2sMURXiYWe30/GfpyBmKHvGMEGQBdHf3tVF1k
xjfqC5w3qY4/H0P60wOt2+680znuXDc5CognqODbFQwX3N8dYudcmTS3urby/uCj
fUXSyQDxrVLg6qwLFrI1+iG34bo0fMI8kNmTrRgJFAuXHrduVWqbnV2BdzD0h8fY
LhUGSE3w5VLPKjH3zskT9T+w7S4axROAnkpZFyXZEt/XnAgBP+ylWGDV2Jdcct0k
Ra/vkurSCU8y/mSuJ4jaDdTtwfbFpwWVjFWaKyuAsJtxe3RyDPykie/VKHsGtKnr
l7Qlm4101dGbcSAEJglrBeu9qKmFj4HD4CXSL75wdmob+g9oleZG9feM17NvHV6Q
szruT5aScLwrw01094L/t/A+VdRNcR0K18Iy4P/4OiHif9hajWMgONGqZFVtdx/A
HrgVPdUoprCvu5VEvgTxekt/2dA5gX1r5cElX1wm5kfJCMnrelzbepCvoCVuG97K
eLRwzMxwQsf8nGqyMm16OdsZpuzAF0HNPqdSMMo95bYr8se0FmdP4l1/P8IxnxXo
CtjQzl9oKwoLiJo3BdpGEE+pXB+OOtXtNQSYl0WZpwyX5c/CPhuOrvFpvwIl7JDG
9V8X1tDzsU8h/K/5TL3C0gcVF4w/l8AcNoIGPdZtoP1cDjJg9HeW290iW69emjeM
WPCQm7uTldgngFcuaM4JyRj3d7OGuBuAPR/QQdmZG+Pz0quporZ/Xvhw3KiPN7rL
OtZqQ/2qoouGfHQYrjVIBPlBO3cK6Ta8KLExFknHlrsHgfTioKLjmV14QgPWBJh6
wec/VHGnakjRGrMjLHKk8bZh30mGkl4G7pZE5zaixBHXHU4PYsPWjYvytXEb23N8
vfAiKkhU/+/9rtG/W9ow4mdgMg/0AlZ7yCjSqs5ebnCRirZZCwqQje5d9+4/6Pl1
/0xj3YAcvgGAg43/wERRblbQtx1fto1hldJAVOGx3/k0iy1u/eaLhCcWapINfDMj
wJ1HRQvezFOLnCzPUXEAdCGSGI39DPifEclcpCHLoE72focbfi6+VR9V9faP2VwD
u2MzZuyb9bviZUQyRWcAM/gxn7NrYhvsKRi5NgtX+z5x3BqAAujSgLb6icQHwbUi
Pl7d0xt4rGc8RfWARlsYaVenS8Wha7JZIGStCDTL0pWH/fEW9Bmg4iQpK2ZvYMB4
EPHHBmxVr9vd0aY0wC63JrEA6dT2AF5b0B/7mqnJbZRnfC4bUpBU7GbSFwYfruR9
VXjkvbUk26JIxs3jhkKx3zAndJUIJ5qhOin06uK2nRYdfXZsiJ0PjO1BLaiVGFJX
yJqOIwwaigi4Mzmga8I+3eobNzQTAudmWSz5PYULxdZnPsMPojmM3zUmlaZPuL5z
YJ4BNUSymIQhrdp6Bpbg0q6d46MA7tMVUTRHe7nbkx6wqfnZzm7oSiS0k3MQ219f
eLxBdws5X2bIhITzjtE5RciTa6CPmnSAcnNYDwBPgRTKavLBTs6wYjsiIgiCC/9H
JTHZ1ycrDpzAZ8MMjcwZPsW5riIwGOEpZhnSTH70eXEq4VW/BL6VS2VCrpTwWvas
RIKqM6uBUzcTv8tonAs9Ox+PepC3FlnrzUwchbAvCYTNDxQAffDkgS/deyl0huhH
/ACI9gXLEp/BY51cLlS9tTWTv0kRRsTdZMxGP2sORnLkvK/6LgH7BRjrjNHGiJlz
oCkmbK8I7Qi0OrzOJbEXoWrGmhiqAwk+sFqbN6iFPNg5qoBpV5Lb7fEcKwIHhcbg
YuUCysT/EzJ5YbeRoz3ZAqM/wjCzylZu6xMAO9P4as2v5ShC/sEluoHS4F22CQLb
MwiKJk+IQJCrvRu9ijymCOPRVdSRJu/9H/AluthppGdGgmY9NNt6lNRJauuijW8R
slctz0MeTMKOp0Q0acK86Vkkyl38iXO9KK1P7zFSpJqHNzQ8uBUANcK6ScZbRkv8
IrpOXIEFD73xEx1f2Lz5/ZuzuhhoS3ZelapQspKk+TFC1F/lKsq2sPWERDZKmjb0
QI7NcgJd+DxTukG4hyVnw12ni64Wku8kA6RgBG/f6PdfkabrwJfpZ4VpMJmnU/g1
rZL0TcBcwIQUhpCM+RL84EDQYg7h64WT3djofuicOjFLA6laxNbUaZ+rIHcbiCo8
+wRFL7QvUXQITd52qpxeK95t1EoFNV/ABbekzjd8c/TTM1/9uoN5NQRSMTEQF5LX
MrV2eKv7MuEfpoWCSNfQ8QYdJt1Rwp/2nEltJCt32Hhnm7YTdClBtUh6Zn40NA2C
jdn3/fBmR3KLlIE2SM8rgCm1YoL4tuLvPH1Nb/mivNNCgiYssVDX7BFcijMBdYxn
F0Yk11hCKCsvfSpsHbDnmw0kOpHUmPlqG0G5PHHFhsByX9xbyue9kcFDK1mM2EM3
MMcHO5LrAeU0xeUB3FhiYaJZpmVa5ejM5Ec2sDvs5EYtLWPeCJd72RoRjzaz6pyA
IHPTigebhTvBgp4Lo+jiuojfQz0Xbx67rF/san0/9dihr81GtAYpitErDcHVQ7sU
cvFeNKgeJ2CPrJo16akOuT6D9Kt2MaSJy7GFOtZGmeHwySliaOQgDAvC/uO0OCyD
oChNM6aOF8W0O9TVe5H79ZpN3uvu9simAziRgU40PYmrHTr2Izq2/U/PWIf5YQMX
/j4rH2/WgF6PmFL3AZuDXowVplRATOdfAnOBFhAVDLP8dbR/F/DYlkqoo2hwAjdG
BRDNqgyPbPFc6AoK/vaLOWwjwsXzHp+IaqcD8PTz7BKF9YF3etSiSkpqUMZH2ulp
4HcVmtFB6qeEaNl2cR66iJFEtcZxScGDla3tNdxHmm2zxJtcN/XZiDZFxg/9ztCr
ob8MS0bAd3LXTSdFrf6DWjOFCZfq2GFIhnytSszQqq1rB4ottGr9btOZbZTgZZXO
TbypNtnjOgZcvxCZRrTgnzL4UwaWfgRLsx0/Ckw9/9K8fRsfhs8eXyLgyWnJRkOY
3ReBBKVPH70dmhci/Krt8YU35GVN23VBCrdHJs6sF0smiZs9mNocKL5P7nQsPbMx
BNkrtQjL8neEMyprOnkSCwKoRWn+d8GjwwUoADjE5mmHhiMKPTbWzz2tt8llEC6q
kLWJGyayp6y32+CpsizUpTDqlura98qMR39gJ1RJ/lgtxG1Py4CJr0mFQkqiWGou
iELqShFir5gJJ28fc1bEFasEAJpvt1zT9b7pyM06EFSwuo8bB0ucPYZVrEmgFv69
ov6et0d4U0WNiMmsjZbgK506ZNyMG3AX9NZW90xksGvMHqxUvwUIVGDrDevrCdJT
HyJFdJbdVt3hZtQuUWBCN2def2WQaQ42jTI15imdGNq0wPc0PQSu0vNtgpGPTF7b
bOpU5e3WdT+uHyOTHVrHs4QadJU/l7yVIC0DexLMXrjPfOjoYSMswX2ZLHmW9MTy
K5v7u4cQOrSF78Jyvmq/cShyIjRV04xtlNqYWV2N0kevhQtLMtsE7c9+EJ1kbn6L
qRmImAlqe/ybJIJfz5qI1KTtRjh4V7d9SrQC2FKUENyv0qsw/0XMYatFdUnYCX2k
JD5Zckgn+jEW4UQ1ZSU2v7fhIKgoNrsQ7monpvrd/KhTgE6mtY4mlymd/sSYYQl3
U7b3E2mjnDMLW1NCK9eriSeGoxqiFKh80IBs8GHRcaa56ozVJbZwjl2wJow5FaX5
UCNpPpk193XuwrbwA6n4CSvdSV3Cvx8A9bot1SU4v0inq9zfWNfdhH+08dhCd+d6
Don5uKKqOcBi1uI/6hbk/2FRseIHe87wgSOvvvxEMJ19Ln0rhMXMA7Pd4lOoW558
noArBH8s7DtC3n1NlJ2POlML7nBoNOBeliMff3kY87V1XeFUa/JCuLpzbJv3ODj8
sCxwuB2MOb8ZpfcClLv/804uW0yOCnIw8DxUwoVegaeNBQq+QAFoYot38ne2n4p2
c13JQHvbEsJFwhc16Fi3MbdlOZSPH1JTVOoJB6OJBLUCEYt8tptrTb3ZDINfaDpJ
59QeTJ/noqvs1WQROjQTebgrCRS7wAdgrx5pucHgQpxF0TU5MOetV3CnyTdba7wY
wtGLe4GYFJHURywxFkGUear+ZQ8MglKPid9uk2BnSisUmFQCy4c8vt7SDZ0wq1oc
j0Xr5JjmaQleTFCYGW2WKjIcgHofeiRmrEzSco3tgtp1tTdBCpKcLnRpbGmzLxqA
HFcuASSK0g9SFPHYqUIppCimbp4lg4nyHhERjpI8YlFFuXtFr6VUWHP6UL5kTcPf
KJQ3Wcq7gmSZeg4DpW2XZOrdWeHVGt1kR0FQaD4O+YPVtevjH+LkhjWCXSoNlzi+
4wmOu+MlhfbC+uXyZTdobr+3OXRNOt1ihBcGbeU7dZnIV5qfUEM50F5mY7rn+c6h
SIDUh340fiPiHspkHY08xBYD4h5MZzmnAgEdSVMg5AJ8b5NBpNUvrtSeQQ9WHc9d
pM8r9FYKijsN7Wrahm0ZDQRIJ/WSgqVBoSzybQvq4KbAUx/mF/v7XldA8hFpefKq
TyZItIRTo9SkL6aaV4BpSbTIMXK2shDuRGrtcuqB6DJsHoPAAeJR8XUEtyBblRNc
v73PUoZxWtzzgqd9D096wTVEHMLtaQYTAnkP7ZfBN+DDCuAdCENd8BZS/JwOK4yR
84rfqtPIvgm2t2RZi2fhjOGw1fYF0YemNGxPmi22YvwcBxAWYiWHNZajWpcWWiXn
aNCEgdNcfMlGMvyqPz4QLpyrc8cG1NHdaELnkekYBJ538ZHgA6QIAqkZ1mbnOd62
ngodA+PO0l/HlgMDQ6XIUdE0Ga3cAy9D+2a9HJnDIjl2KB16Vz2bK1MNBF9cLOc1
ntCYigognEbKzYj7PnOoADJivqZwmq7mHhJxJzg6ewgaBJRxMyqHMDYiwD4V63Xc
VbP9FBTd7BZGUIt5MtmH8FWsZktk3bkhRqhhjbczFbKXLF0fTXRZ0YeloY5DruQi
dxEpKVSZZjElHYDX0YHCSgtVr+wUXtKBUttvsgNER4yvSezDXT9p2wTF+tuYeGTa
4DbpL6QGqCGAztm8YWsXbPC+pFP/1NffUrYfpPpA9a5iN1Eh/0gLQMnpJmW8f7/q
+W20Tt+BsitzN6+m7QOKRdJ36KKEBXgEtkj2Pb735fx2SkeUCKcJ3MIhOR/yjXEF
H+Wn7b3nzvAyqXgQLhT5ys4myKj7jXjYChlQf+5XSXovb/Q0EKPFyHJR9oQdp1vD
VT5CIXILOBr14mjTUWLta+SxHkXqJJbDs2GfGbEWygGiYgfFC5dX6rLhDHSMfgSc
UGeuoABaKdKfbUfimWoL11kEXUDwxNNRatDgZfKQi41bwZbdN7xcnHVJ3cMSAKK3
kQaGtDvUQ4aFgnL7xuaU4WyUJ/98f4r9ffSU4ja21M2eDT+szGWoc2hpClKcQJ+e
wVJBaGzJHkdhyIe5DoNEEtjJ1AUp3czYKvdfqKiRLKN0Z/+tf674IzttnKk33mkT
grx2bH+pBAKfb4uFSWcDuIIjxquKlL5frxohp5ELuOXQMq50OF7qr0QmkNaSG1Dk
mcGjQ5tavkayzigQfhsuEYuZ88vmNdhKklfE8m9sh4taFXGZQM9EGc2doL/QaDuJ
xVliW2+OZYjT8v6ICj/Zkru4sKVUV2LiaJBLnN3KIk40guvLaUDSeAzrdRiVN4EG
I5rZJ1SpFWVC7IUS1Ler95pVJEfvmGcIdhlCxwpjQaWYopJOVzgDUgFrSUbSE7i/
HXrItHwDME/0QFw1BnWyrgAKIbpZFha2drxnPHacN9VhCPHUtjIimRAUJRZOPI0L
VJlsnh7r0M8o8BNXNoUWTPUme9Peqkb4mklCAZgpzJbc9liQH5Vb1DrqfZ9fSJuM
4ZAjXJzTf2onua2P2WawX1NgDfLelBr/zMcMZtLtao56lnt4AxVcuNyLovAFbvf2
mkucTi4ya2vvRtecgBLq6FHhlvn9aFHAEJX6VJ52fhYxVkJfPRG4ajP+RNGgMKrH
7FUOBCOXPg8ErM/3SdyhDaCZon1hHN9fBWd17Ak79AAX63O2XNo+E20Jw1h+XT5s
xu5zaECBQqPLFnap+ulIUTgGZ6kyuo20X0ecbrU/yzL04j3OCPnmC8DYFTjB57JW
C19DWhhpStYe5E7wDEjw8qezjjjnmLAOmjpUvFjKLwAgw4ndvmbJMUmibtjhKHOS
5Wy/InRRqeOPUbL6WHFzHnZlE/WPIhj60gmB6cMRgCp26vqueJLIXsswQfpmtXx8
IIRV2/zA/ZxQBuBaFnjGZDbTeO7fGS6Re19bWh8/QREV7KJsg0qza1gqgJYTnhtb
i8zQWu2e5xxYgS6tM8tjzwoZHO3lDQ5rjCFOdMLHLj6sb8IBe0v1yt1bycBhisy5
JXZEEFoJovJIFsO/7aNduHFD2CrG23H77TbQHWH0YH0nVvVQ13Ln1cqvsKmyK58i
2m4ImHKt75B+1N5moWpt1b+IZ0S17s3ioBNRHNnV15Ed1BHBpsarWTAos9rVFYK/
xINvn9gtZCZ2wgwPMRxNg0ZetXCzZylpORCEPEFm2sf/gHumhdFjurno6yHvbGwh
pIvnNSiY8rq5dw/1cDAarwDJvxh3Ers6t/3ppBYyV2wGfq85XN9JWg1SrQr/VQBd
Na0fkw+K6FJazHGy0pclstS4+cdVoocg2dRzBj5xlb/5PbmKSTUXMihsMEkE0RLI
7vvG4ASewoqqVz3MrHdybwMUTug4edS1o87mFU4sSX/Bn0aqBELZJ4CFcyguqn9+
gkysaFQKWm061NFhsBrOdfyTB9ZiKBDw9yHseIx0cVK9N9eveXbDoQyNRW+W8lNl
yJrX34ja4mUYzlixRp+ipgx7dTpo8WWu05T5TB623kjxx9WVbXjOqQasHkhnxFkH
isbQzd38IKM76TIYwF8ygI6OJMYiQvBh+5xNZStTwNsBTQTbUKkZsVsKHzTNyBj8
qygBB+wLCQlxz0ar7PSAbi1QZO0BCMY15mO8gqucb/fC26VM2Z0RoBHVjYUfJCNz
4bzNG6VqfusSId1kCvR3BGM2yNJEp+kZrA94r15zlnHsoXNL5ISENh1YmOJU/8lp
cJ4wVI0BKL7x3s1mwbYEjgXBqVcJ2tB8d8eGTAOxIUU8LeYowYVrLKE2N7CKFv/7
Qb9xZyJrdmyyzcyJLTkRf7jMKSGwVaH1HOqB1bLxGQ5TBWavaVWWMgmwFlK++C9Q
Iyk/z6mD10iU853+QVZ1NNkS2DWTOEVHB/PfqN2avZiLIoVdbIr8KkI2DjxO24U1
ImtGoOnsgO4dpee/2CKh3Xvi8WLyKqSyb6aB0idCkJR4xoNIUzGFLW9c3OYbucZ/
VEVSlY+VjlsQoffupG4fLgqGTbSONTQx4zfoiw8n7BpRvEvOv8YfV4r74OCBLC+O
cYNMZPpwK/Wu/BkJ3hXbbBe1QhN/qk8TIl+IvMZy0vp4fiqbB7N5ACb3WQibmL6o
U2p2GRP/3K7pYcqechPuW4YzVuL/O2TSsOAQ3DHF0wG43Qte/gvQeJZF8iVcbkEL
GyyUocAoX/W3rojx6W6b9v7Bj/whY79GEop9iUcODXpW1eGPM63t6BaIPApLxcDR
l28z/suvDaDU9T15TquobGt+wnROOZICtprOuU49uIuSuZgMTlX8Siol7g5d5b33
mGi3vPHxmguxtQW3QeQvKot37Iynl4cAwv8lkfJv5HxsMhqYTxCfSJDdblupJgbv
ApIGy6KjLWIBHrlptusBASkK/PPwV5Rrmirn9lTgASRFnmf+j8nlj/RH2U7xL17H
GkCVR1pHNvOnZdNfpxHhydyS9trqniNLilNBIMpqiP3pGoqtMSyq8UNHM8T5o9ro
rhD2Omnmxtg0LOwupyNDgCQsYm3A/TAg5wpl5rrBeQcXH6fiEX3ZID6HcdDmg0qN
r0W6fxMdlrkwJ/6qyoAJUgy4mJM4yrW3awlco1Uhbjh4W8MvCAZdngdg/FQhHI9g
jmZ3INnGRo/F4aqDVXyyLiFIVmJ1CyB0AFBj+aOP947TdLvHNZyqQJWLxXlXbBTV
mktdkzxBD+cXMv/7faw+BSb9dod/nCMoUUyO6+mOA4fwXF1LZNFSQUoB4JpCINPb
VCUmHE/yMlFSZdRmXDP903NYM61IeZxJlw2IUVoXBG+2HWEi7WjAs+sAY/wXAn8k
RfTklSn8KdO+11DJ6EWUSbb1iiX0Nng+ahwiXMg+laYVMjouqH5LNDstldDXHBza
1MFexaa1dtNI4cNU+v+EprCHYJ6OhrXCBB06Thaf/DpaJ1DaCJ6tujH5us/wRREg
rgTM3dYNIO/GhM3ONlTs50DlvOqgRBcs5Zv4rzBCwbNfVCP5IBUIceLumoW2rDcc
APkDtr3loEEptAam/EMX16Ia1Re3+HolHxJJdTeyGqP5ub5noQHXijUiEbgEdRWn
5t1w5heCe3wvHq7XDwit69671UYuDHOPdVYqhSnAf5VPtcVj9GkpI0Memj4A5kw4
opQ6iFUvQewPrNCKXrHkB6pLtlL8T/fTek+RJozNGir1Y6UxML/Rb/GLcEzkNxO6
Nr2x86a310yq88i+6FquHKFLZpVcRrKmgxwD8tV0JHvkSFD+uYQAq+ZVasiaw7/t
8TXQJg+OqFEJsuzM78I9CgEi/MXja9bk6834McZFt1mINiV2JIZZs0qkZdVIA973
B0M/7zPue9jIP6EOqVAlV6D6SCrO2ncKy5PKj4e1xMN46fSkilIEmm/9mtJcFcDc
IXPknwmraiIz/jpSTrPbAt0ZJygxadY8kJcB7d+vF3ZxqFQ7WP2J5X/qGjd/l0YW
wZ00h/LBDLR5OC8kkZy488E2teWK7lcMRONsfMuUB52miGsYdRjeLVJP3PPwbaWH
2SEjWWw9QVneO935OzdSi2dXiszSohR0mIZ+OHuqmtBfL/oBl0q2zaJ1o+MvQMJX
6BUIqp7BbGTly9FzaQmz8ZlJ9kmGTNjGXAlPaycDUhx2/ZPXbfzzdlEqn9i4ZrN9
1JJJRIj1AFCzuoqw1GiDNyh6JECi0gvf4GTULwgfwPppSWRwGIgIzPYg2rD9inND
M3TKOjcRm5AmINIeI5e+sb7Ke8nEidqAISOOMksShhEue99MDzHDMCbDmFlsb+dD
7Xp2uYTFjwHn7Sk0jqoHDAwGXU3EyQjvqzEgysm/N12+ku2wp7lUq9lXh8VnS7Dm
vtSVCwFzczcCZJ6sv3sTuivtY55Xjkp44UQsygrTFSNC5BnmIw99QwIZwLPb5Je6
tApd7GsTNeBlxgq6kjFmgm456M4r2JZzhEgNVvwiTsZrdpCPqrRVNv7e4mMBaZ2J
rC3UYdZ+zU52Sqk7PE13mFquWm7wyI42V18aRigJ7WnkqcRdAQC0tRexwbOJ4jom
+H88rD9qoJB4wA2wnlb7LmrEbC7konjRc6MxoedTmQDj8D1J96kaKQS/7MEBVcQG
g8QDUfhTNE+yQ0UKLSZKMnnXYFv2sv/PWS1BbUdLLssg1rubO6UJnTrn/rWbchzj
rXruGPPq9/v3ZUSbPKBkZjZ8Prkl7BZyoZFztxwKDykFi46oI4ZJ3EL48wGee9nw
cHIlajSgz/jMltADvgBUPJzrVcBzPaLqRMpeBAeCWFfVQsCc+my8ybd5S1HUMTml
8Bfg9DQkm6nni2KXBluE9HAm0d1HzxcdLfVnR/V9FAECl6GcBYpczkS5+AZlE7FJ
J57aUls9tG8sUaiT0pYdA/mRtfy/R3Bx5QqeCmTEVdlD82uTvQrTEj+XrPeK8a5N
zDWljjYKrXQ7bRaL6UHnJ6eqYfTbv8UQEW1j1sSkgsH7rnuE/nLDspz9pSEinGzu
maURTunHv7gN2QVFwyQxSjCuv7LU9NRH3pZC9WC+t6ey0MhIURYmCIwjCwT0ienM
30G0FhIBzUeyIru729vz/upUcIiyzqbtlqbX3ftDu59emY2Z68BWMcjkKGxxF1zY
949Ctud8N+j3iZov9bOwcvwnfP93YjQxNb4VwLFwKReRl5B9objUykUuiTE9ksVZ
uzHXwSYEqeYA8J1MpQtwZYGCBeakFZYPt5mLDIZuRRZv3+i13oudo0V0t2iEX/Zk
jIAzCebbnrTAv1gpqCD/H5KedPa1aRwITDXdwcPmY+KdhuwJM2yCrZSk8/nL4F7R
pUDu63iygaRRpDueNVAp6/bhKxMoVr688GFs43myN4QT04904vrVUWiU4gkQq2Vv
170eHuwtf1jzz23oZvmuJ1duO/JDTeyL2LlLpO2I1Fu2igdX2NOYRBhdh7zTupnE
JdMYGfJBvpCqxi9Tw93CoLakOt48lupqzrYz/pwhWF6tDSu4RSSVCDoMqxAElJoP
/Hu/bfqRWZklDJXyHg95h5VHW59/6y/TIq9aivtEfryNa+vnK7ujH5mXbU/soJ90
0+VnG36DB293b33OpNr7scj2eipq7c0ywshzAegKSUVeN/5fv4a4ohQxFYxKg2SC
3yh/zecQ5MjANd9Hu3c/FQNIU2KdDzByQY5NsLFL0Iz/1p7D8VmRzWEMlt1PLV4D
tAd+qidIuEJwiMwAk3sEO21YPLOGrL+aUbJZManp/nPnO8RjgTUToOQ99QC5LUmC
ebVlS8AdMESqRKbHbkXxjRNZJEi0rvTsYZoQyOZrmjouznbqAt9ZKVv64RO542Xm
rRoyJyKXOKHaueEu5nc45BmjQ6LtTGQEyvJm323ZEWnO41ziACJuMj30DpuXrgvV
iznA7fqSRulburwLav9yWV19BIbGeUoEHA+Pe9Wt4tJ6DF/DKvR4tEI5p4CzbI7I
nk8MWFS0cvyLtKlnH0HZpgOf+SokW7v6CQ7djA6tD+eqZi5Z0iqmL7xitGi+aCk7
XVQMe9MIds6GwhgwOKCpF+c9VOsK9Flut5VkhCP0I1/0Ey7GTN19AoK29a4FW3X/
ogARedhy8PiUnKGuT7mtJJbtULMwGtAekaw8ao/BmkhvFRV2oTv5cLI16sC1+0qa
f52r1ZOfnpWEOko8hNQEuaBsyKCrqazPGJsKDsq4dj+dnoF8RUVQ4KIdD/IrnbpI
9w179XkMYwWM2i4GexLyOECOQO//EADo1A/IlRKro3bOLOpVl2rmhv953LlICA+y
dXK4Nqh2jkPfdfUfIew2Lal7lT3Q7B5TgQD1g1aSr4uGqd0leXZFaeMzb1wYcbTj
CB4Ws0/dPoybRl3yXjt7W7+1ljlU8i2fZbrYYwSSrne35hyyDwhVj1orAMh0i/Fh
srqfNwFk1QnUUE9NZazELLIG2A3qczqnn+ZDTMlK8eSnGj/6FOEUEnX4bUyZdS5t
y8UWM9YH7YD8kuY5T9HWaEbcFpbEbgdJmwO6J5LkpdZ7SleqAdsrBVLqbAj4FYk6
GgIpBBtyIozRaplMAa8KIroBwmp+qXcHKOncJi8Rj5WnkrMshoPA6JFWrsRqcjx4
z4zErOUMEjiEnpEld/zu7QKCH5siJ7/8czWwtAl6164iDd2F3kuC1q2jygLCg6s5
uzoVW7iujOisNKIOlByIxyxvGxX87Ne4yrGGpyQX2kRiz3mwleRLuyU4b7jMSFIh
6ii9FbVIKBxcRW8Tvi5Q+tVxdudSGwoEuY+OuUUGfoncFe7dkMq70m9uanoG3ZEI
V6EQCcd1sR5QDLRJgPbmkFXG0Tx3xHlMuLscTE3H6TGIlxVBDUJqDn92NitjyjSC
Y1I1smBfyBBkMLtEhsycvgNCIIvE91rwYxgI6QgA1UL1S23IqD6Hh9e91mg2EPl7
yyfjNzvA2X4H8XHd7eiXMZZofuBNO4z0eboS7CyxwzoznXbfDj5Z4xAr9fdxny7j
Wj2ykh3RPJ/VDb9tUvF4525mPV2fY+9r/Mf4liTbZwuL0vYsS4/zjp3P8E0kLB1j
vt3cX/eb6BkuGJd16AzeqosjXgNmySfVZj9PV0hXoFS9hm8NQGg+icZOZTAmF5+o
LwUk91DzO8Bhfy5Pbu4+6d0AYGJqA1GyK+SH7ntzLufXyyph2vsibD0o+BvZruwn
HWwrIvM3Yju6B0SHSUAGn9iIb+fljv3CMwdM/f4x21Bj6jj1eUvYdBTaOUVYCXXx
VRZvf0yupLIcQpDscbb/tOaMcrpW8BQ/RgtohdskkONRjWkMCFv8q6sFFQEhQh48
vUKEoqxNR6RER8ukf48jXBObg7tTr4aFdlKEPdPL4R6bzsG21EQn1e6dvg6d0up1
vCPAvrkB+iq1FPdYKQIxw83N9n9sg79O6Hm/rkwEth47sL/UlOypvu9DloBTorvn
wrcSrZi2v7xkCkXxavSOSAhosUGljisS47+WvRbT0ToeBfYl7up2sI2nibb6mBVy
+5zC0qtfuiATpqArHO+Q6wV3i5K/V0UymbTL9MDr2wreRPYZ356zAChnavKUD4r7
ILivQFJaoRong8Rq58Dx2rhPOc4DbQ+YjM1CuRtREdA8oSspvLtd06XwPNitQ9CP
BpWbfXIq5o6CroiF0HWU7l/g+nmffanazEIU5d2xem5oMbiTZNLw4+ls68hUGoLN
ulS2syQc1xbBAGBbQTxso1KKoFZbTYahUae/0PeTeVWdDAZ87O49hZlAoefTBnkm
DaPVJ4RbiPl5YeDVY/bLf6Wek7LfN7A8AHXFdwxuJxQdtOt4Y2FGRRUrTEGRHF7P
WJd7sgiZUFqJwAsS5wQByUZ5tm8eBouLwHRxzyjneD0NbYCxVqdOPsA+Ty/70oIk
OaNJnW59RMM4vywtLhfAOCRSM2s8s2BMf6v3gM2X4eVlpCb8LjmgO0baLv4akf2t
WnwKBmSTQtL8mj/QhbM0GbIROq77+LYcdi7YvgNzRUzLHhZIxjeRaMgBysoBTkCD
Bxc/++5q2xax2crorwdQ6vX6ZXP7w5tvrnP0rIuW3MX+5yvacXhfT+i4/5gGMUNA
Dj9RpaXyOjl/0I9XrpxjnMPffSAURbZYSYB20hT7UuDElxVmXW+mDiCcfMI3EEDf
KIuNCND8Eq7AhcWSVVTqpot21CR/mIVnCiNEAgWVze0zTAWzQ6bmq4TGmI8W3Srl
am/iVapW3A3mEvkmROPWqxozl5sV++WMsAlXV37i216y9D2a2FgiMH7Xkn0r/PeL
ba0FcNwjUuZHXT8R/dHTq5Q84VXjRy3RCjwGBLNImvMoAwDxWorxw0vMcKi53oES
FXTYudvVt0VXuXo0/HsMvN51X8vlJSYrWLVkhnLKLDsDfrKxCq9gKsOPQEM0K11d
Tj8ehiEA67Lu8Zm0c/B7Dws/Yu8/U+hOU9YE5Z/bbrOLGt+wDGBk3otPKgtCGdpK
9k45Bk7O+aJnu9fdUaLJXRFMwioXwBpmSi0rRD6sfmEx/nbhiZ1DhfP+ooeV+ALI
mC6id+L8jQehM6H+NxMCjSOw3Ms5fEgtqVrc+/PRe4IVQ+NPsODigXsjTZ/lAnGW
jJ3fRC8Hyi0IJ930q7YbDNqygrT0yD3tWT4A6hHs0l/cec34iCMgPduzrJOMygzr
YdV+eW+kOpPhwH/ELoy2DSTuuE0rWVP4G0moRO7vAWwoSry7ugEgjcHPviSoFIx3
E9Wg6+F9eUBV5hoSf/m0IpUvyH+sb5qB2mtaavTjx31628kpr0Ngh9UNnT/XbYY/
rOkcMskEDjcu43k9Z+TlehfPX+Dy+r+5RqCjEiojSOJnZOer85E5hBn6fhctzAZy
N3HtakhGIF0i5yLcBNT/aw66uz5DfKuT5OUmWPQ45WvOpuI35RewS64+5mJqUVhU
2KCRJSepeDUkpW3gvcOgb+Y+YonXxv8q4pWmF52TobkpYOvOJ17hDHc1cmAVOb0N
M5SRbXIJj8DvdRnfJnTWRbcoZT9KwcfcfwG8Kl8OF67AoeOz/tGbZoLw865G38mF
2OJ0Cq1TH5oBWsp6njqKoKaxLIzz0k3sVQptsQKwgC4RaEr+2Uibors/hq381ijn
4XBGh5AGf4PYHi/hx7kfG47ycYHwF8USSRUIBkyQPAb3TtcuS/1ApS19I7DI9d6n
RpLoFQSQklixr21+AeLsoRW/y3OrjT6EVcujdeAIKD95THoLGL/JKHx1Md6HAERz
Q9Cfs4ycM3aWhQuRTRs4u3JCMf24hVvWHJrh2lAs1hIqfq5LQLmkCoEtUA/gmFzx
kwiE87JzpYcjA6MdGYuj33r7thRKaHDEFZJowNmdW+7XI7LWxsFjELr9vBQbIsvk
I8TofzHMjVJKtEcD7oXDvRQ+oEpKvl1glsKc2gMEhkvVIXRlVsH+nwcrbSqCeheu
cv0d4B85E+tByrpEdIK17x8KKRwiPl/orVkIiikCkjNvvJbagJDQrQicPn1Vvrn8
TeqoiLegpDksc3go8xxkzG8Me/aZN0MWeh4zGTZtQSYxYhhTBIp8yyGHS0DV+bTH
XyGALS7BWz6AGc8chaMaf3JWOXVVcsrzv+W3EiF4Lws8S+rjdBqXvMOfFpsH15Mi
pGkJLI4YzozLj1M5y9XYXf2IP8D5w/NdVD4FJ/FtALAyW3S+SpOE6JohXKjN3q02
EwlrP+6nXgT9czm3pDUbZWzRRtZ7oEpenj+ESV2+mpnp3jaiHezBWjQHQKOpyhED
fqRYRPSd2c54Br1UdSTaHgxEsLNCTRjIMc7aJD/8tYAeVM5WM/6mX2quBrjrBdcm
KoU74RCGge1T9eq7HMKGWBOOVi1Q3hty4YjQHWRrhvyxt5wMW8OXzss76/eYC+hU
X06dj3OJ3i7NtyyB0Ki/d7F62wMUXFKb4KdNvQ5Ss8XPFKUeNzbShbsAhfrbUg3b
4wOljcjmc8RLGcqv8t7Bjgnjq+7XJzdNGvHBBS2sRz/+lHjciGdI5CeAaL/0p8+8
5QbxzEeeMd1m/waU+kuGxFMKgj6R1QL/hDsGX8tigdaliBXkNRJGnrWG98J8K3Zu
rzhmFowIhRgiIXnmDOiQiRAd63OuW3mWTSj+uLvqGbNvbXjOI4JIIQ3KqJXW8bUw
sFJPDniYPE5ZLLTWAPGRAO6y+NYCOhT9pVcdnNliPF3vRR4K6mFIW1QkwBk0JyJU
z/qzlGcvoyQC9ehpyR51zjwfW8OgjRiy78e1Xrgbj1EQVhU/SQG96oS7ynvCQDYl
zOvDCsQQ+I/jfhaKWWYbg7JG/NYVIiujpbUKLIZmUjLtTvcP/mp1illgNctdvOR7
ZZYrfUbqhUe7VPIj2WrwSx3XHe4U6gjaEVjEUBbTX9fEa4DLWUcSWOgSaeVPYtX+
aGf8e4mRrx5UciI8FCGo3DnJ9aOZaE3o2d7l+63TuHRgqWbwvyMkurHAe/Sx1Gnf
ULiWQDwQsUmLY4sUm676Hg8iqfqLN70TftdmZVvmQuLS9T88fLFtoeohkmoS1EpH
SbfNpsZ6PeTr1KgvHQK2OFCi2P4rjgspBY0qSRrjetspSDwmwnYNn6FM60Cx/+cU
kxTuW1E4mPjD4Otrq6dl3PsWBOYLaYYKrRlIGuI1ntxtU0IZIxeixGXsNupEmTFr
084knmwvhkQP98zCfCNA6nHhLhFwBhhp/jL0vb5dJi9lvbR/oplITq+jzqz70MBS
k4kwznrCo17DcBVGp+Pqfturt4ndSAYGdhNefi5ilYO94cMq4aUBrtDNY+BbaUBx
CEG0XLRda9tY7LCapHFVYIEnM5NLRQ9jME7lj94GsacoxgNaxK2UQhYl81NRhWZ5
RtOGhFmjnuAA2IJloQ6dX7AIn46kTh8SaQqPz/HfEmCSJKNbdOkherhEgZK6YsVj
efrJ/T0pUUbPixLVNxXXBSVV1fU6LQJltqV4LFD6y7P7MmMvnNu3Wtmn/I6851OI
Y32d75LJ/ddUdXRkscR+BC1DDC1yZ0aaqqRxsX85HiptrlLwaNHt2xHTvRELs7tK
hk7GJVKbFoTPAKMu8+EXdRdS/Rk6dBBDugWUaiCaF26ZsFK4gHVTEqx1F1lqsO00
3MCQUIg6/3hNLBK9DJZYOt4jH8h05u6zpvg4SUkIxXCSTYfEorSC0LHHfBeyVTae
qvjqbCRTd2yMlyi6fgMSs5FHc3y//gAwbgubGNvpbNL9le+pxojJ2FB0SQ/hEpVs
W+R4K4+gzZrXkNzNjYJjLtqHvbHR0kFkGvqjiy+4gMZlCJUhlMLgCDzGvAhHgqd+
n4hPQrLT9oiz/yfRJzOYgmM4OyUqNjtNQ052nl89WnFsN2QqWMwU1xox03LrJDVH
dZbZlPC2feSH7nlHBSSpj+QO/OfMy7h7qFvi4FHK+faRr6HPVC5GSv0RKlDNk/D7
0FAZJxN2v/BvvL1kJuh3EyLpVuEAa6KX/gq3GrMdGHmV8gn1uM6Cc9fTAEfsUXta
6VikoGtbs+uNMB82QImkhawxEblmBo9TlmTtD3yJ3AMbykZJyQhaGcGs+fF6QdAi
xRB6IktUR7l4E4r/b4W5V2CMaM4IINuxRDSRaSMpY8JHu8MN514D1pKr2AhqbIR/
BvOVeNJa8KMojWTu8zi1rogAnLlH4SN03TwSxfFLZox6QDKpkNePnyiZYYmgJUVm
jO69VbQmWIKkkyWdJUQBSURZfa6+emxXw7PFSfQCDkg9uaBNU0ZvR/UEx6yG1dsn
UI/kYm5foGbxOZzbM2sRihlCDI6tL9HpKuziKLUyGBz0oAc8JVyB9/LHRdsR5kas
iTuZyXyp8wt5SBV8lUByB44r671G5NuBqYeMsrPAVgDFbjWBXzVwc3YnLtJd+lcg
kpAvqPtog/VApgUMTYFOU/QaA4Qi8udGNGYlAiOAzK0UHTWmWZz5C3p4I6YmgPu1
v+dbNeTO32sAJDE6RwotU8BRdVvMTCygKF38an+qfpDhSK3pyKDXw3wfndAhuFCd
rg5S84pK9TooT594Z5pPFE7o12cmtoGuLpy5cjlHQjDn1Fxdpd7MgIBYkcB4rDO1
JdPNbUt0UEAocE3oDYPIUVQWh4q51cpAxEiU3VQ+/PnZ2KAlkvBYWz4EUhEmXPYy
Q83o/U3bh9b+sYGasUlAYn+cC1cMJV+yafOQITQXPbzOlnWIdFHHK+jHaZmlTeXb
k4VlxYMl1uM9kuLDQ6Xx0eAVDmg5/032hkHukDNLeSWG0RTdAxHg5sMCcTdGiDzC
kY6LzQHTD4tFNmGGbls+V7rbA+ppWGXEDHAxWOi+yg77tV8cRAolx8liG6qfj/93
IxGWY0C4zWSFVGCTPmRXypJBX3tOk7LrIYo6Le4QrncLzOyeP53/udSYOYLkoJYP
1gX5DpBVWEu09zTtLDWuT2jSTX/T1gG2BIGSfXaCm1Fa2M/VLk4lT3STZk/GW716
8kjvwK0ParOmCCW2wurbUdxgKp0vXCda5+Y67AEoInUbpEVEXebZyq7ptKaC7HRe
7UakLl6I8wQ0+OwfmQadiDQurNBnnJ7Hn8URPlOq6WlwjEFuYuNL7s5ZpbjCtydG
Rh5VtNJZcBMGLgHJ4iv4CbRzemGwIY4IlIRmdz5NfIl2qh0NG8wOqqjwtSp/fsme
bFTbL9iemnsxSkFEes5g7qUPiN02jEHay6aAZz5IhuPO+jt7Ml+lVR7NNPI34HIX
MQFcwcydwxDg27NKYciJAWmUz3Ge3+p/a7CgX1io1VRLWy4kBs9kaNr8koBOaSIQ
rgPMqfS1AoyRDiPCFexUUAoOXC25WYuTMB432Q3ng/tP3O7Ka7Awf/pG5icTnEM/
Lr8EK6bOpxNFxDiYL8PQdG14LYe4T+Inu9aIFMMDQDg/KOfJ60FblPrAR1Ohz/PP
P2f2T9mzz8Dp3OsLIjtTMytCorqNM0OG2MlaelITrmBw443/UdGbgLkhCknmGjyY
5fMwFlnWXw6psALfaZhsDk4Ir3L+Rjt/62LzZhR3IIopRJMut5ZZHE4EsVcC1yY8
UmBm3T4vcRIRzGKgH8URKDjTKq0RVP7mvuoc8SUkGMGgMaYcXii7kjPPvcOp+cQy
gn7/5sxtHvkPATffDletwh67wXi2HFP6iBomlCrTCYBIA+zicUKombJhazl5kEZv
+D2hU+R9Z6S2+LKhIYJTuVXdURrVPccaab5oEuhw8f2uxrpRGJG70NBZGpp2LKDN
pmoe19mtQ7nyP7pfM46XxRWTWGu8nIdchY7Nymxr9MjG2spoaVgt5qJExacuKVpo
H4XKYoycbGTMh7ihtUS4Cv204UmBpKNtyWIOSs5jlIPqJFZp4aiJOhFGLE2MjvRL
say3FQbO1PVh56OiFajNdk6SYVqeNt6HfsxCYrAS5Q/5Em1L3fQwCoPCYDuhw5V2
Xk8o+K4nvkXY93nhZrTK9OeL4tiQZ1agKbWrCVFL+JTMTQDgCvlisUz8D2JInSP8
Yc2H0dUf6VWSWSCbwlNJDQ3c3opNj06vgmZOycxBBd/NpYiFTHS/KFtXsxOvxgrG
/nBoWL6mzRDCvrKOZVJVerfKWkUO5AcfislFPGuyhfx04HAriL6BVzFkF4WIgXva
ZlbctwXq9X/xB7VZ4pmeNCuA+fOa8vPo09xn2CasgE6lfw5Wlz+Fi0t7Zoss514K
umvlxwmbfMpFYRO5z+gUjLmG6dJX0zvbRfKOkw4Q6Yau1s1YM7zQFHQ3vComNJjd
fISGvTEoJEyge68ex9kHaAZlkxzXRh7kl8t+4vFyC6uSxehTFFWZD9Pjfwf0Cd6v
OkXyYmoyDQIRin/yIwhAPLwnGYM99rXcZQkxmDGqIHO90xC3/TS/+1I/iNJ5AQ5B
q/2CpIKuolLSXDRbOH8DT+Tx9P21usMikBnCXg5MYH8OKclAmlxK1kVUDq4cAnhm
pZqlvqvvrRTOSk7coZdRA49/BvC+zu5Z73wTnQBam0ThwyuAucRkEWZ5VDq4Vlx6
uQH7Gi/cubwbxmOKeSmRMeF6EhdrtPufz5hXYlCzxgSnv3oRcummg/81MWQgiU3z
NqUJFtTRfihlhOjFSrgsvon7G1J5UnNaDwHO3Vt7Z1sLkqYH6AUVggVPRKsBCLG8
VrebbScgx4x0wG/dg0tDXEbw881C4rFdEjSbGYY4WAwQ/7I3qHPTm1ESZZF35qbe
W4yv69fQR5foQEQA58fxjgbmN3VUygWXteWge4FB6yQKA1wSI4mW20Xp6sOGh7U6
KOiEDymtlKc3YrATmA/A61gQtB6p7+6ERRJzOwaVr+h8RyTqMCoaGa4OFOPCQFV5
JHuO6WPpaleGLWjEl7Ida3k8A2uKlg9QAz2KTA5CjWmKMeOO2YfJ7Ky7jXp1NF9A
+a7THh+S4tNtIWfW/poT7oraOc4t5+XFSSMRTfS8eojRrydL9IHStsum8OjubgJ/
op9y1hwQ3Cjn9QuQFRfzOiYvC4GxNU0bJgolqhRHn0oiYOASJF2hZVilVuRJQ6qQ
7DlRk/1ZT3lqPzIGh5jpBZpiAh9KJZHaee8PIedyLICJeCIEJOhlSKra/fOT5VHl
VOd6CmNBlq6s54R/c9qBxjb3TLCMKT8Z00NpQns8KDOLw0F6P2XRpqSl2RN9t85Q
kIk4mdD0xf+dM5exbcmGGtly7bkkysYONMZ1mJwbLuDSZ8kAhFtsjEPGM+6jnhbe
cKTGdbt2QzJVidVNo3hkJwGRjBeXEzb6HcUG3LPWjSRO/qmiMIPb7nAz2/eTtv4W
e6+nhnxaV9OFtAX6vI5OErfwG666MySnflLeyM3i84IwERa4BKmyhQkPY+kwMeoI
T2B5eZGG79QCjnI1MEqli/uiwkQOXqjMQ3vEuzrVWapG5v7LxWbm+rsVOSePcvr0
Y9ziGUFugiX65TmzInLrthLxqLVT25ATs56gbqaVmFwt0VSYfQgLhYZGa3Ka5PBJ
RVlNSCgzkQNNgX8xCcIO0vFWAzQJsImnrzhLbvlNyVoPpPlAOcDpFr+BVctTkfiN
62b1pG4PF5Me61C15gz/F+1PnbOJwdgYz1gzxtktJnsaxbawEF0oIdg/eDUUyXvW
hZvM7w8qQc6erg7MrHkGY3gRbFUlT00Cn58OG1lVH/Mr7DMn6LJF9ln4y2W2RNul
IdYr6nIl9EvFCGN2sZpvNVrz10BLgRB3l4cipWCjMz79atjFwdSzhPzZWr4vDQVC
haK0pbEpQKK86p8GQks7H5PGdIzsu3fWTwLExyslUM98PUgyUtbGiMf/r9/Usn+P
qromlYjVbVTPZ0/ELNmYrXUaa5i9skOvgsMP1k0rixcLv/3e6jD5WxF87J5Ngr4K
xu18av+4l2PkhO2qPAGS6cjLeJO8GGvhJtg37swdSabNiDuPrw4pITLdEj121Vpu
EuSCKfHQoo4qUv3jmucPWxuZYjb4RycvVsRM3II27ffzsf/sPsddp9/qpO5ojbKb
XHVMwYFFG4xtP4AlYgIRsWEvQx1pBSgkNAqY6zBwoEawzrLTr/7k+u7twIL2Y0MC
9+3qUHEWLCgMxTTPgHp7xSfeoHF7fDWSpDydzeycGKSYeW7F7N7IaS1H4o2AuzUS
IPl2Jde3jsQl8vyxPL88o6huktw26qk4Jdk1xk1DCFh72Mo9WeLshnKYrG48XYZe
YsGTCpCH/TNZiu2RdWQAPEWsOr90NSdBLBxMpuDVtygajH4vOhvwR7HQ/Yu44c2+
qfd7fwRQ1h8AcT+JT4p8ghL8zy6wfPo2jrFMtQEN2v4ogwrjn4D7RfL1SGknRJwO
y9NYY0iNO12TGgCFc7XZbg2ICEcjSAVYkzZNrPFl1N52vZvqI9om9deDU0nmiATz
1vMvxw8sQHz4xJFvSwXSW6q/UCnUkssUyUH8qnIKXmxvRwwHiouoaUP8dF6Hgc7y
T2kWAM/Cu6F0hXokb/shO/QjWx6uyA9+hvKiPuZV/G05vMOFNtIzb/qJpTZlefHa
9OZqUyZm9KUhYXn3riP7+0hFrBciZS3FevFvwOjnze6F1hhPUOBqliuKuDpYWMB7
izLI0rL3EWH21WlKNBCcMFDFmY/s9ZwXPCntdmwzpN08rXkRA9Bd25x5zJlcW3hB
5L5q8L9MK4wbUW1p3vdLNrhtKtdBoyY36cWt1tlphrpAnMPq3RElp3lJZRf72snJ
uJyigpR9kyPOa/ciyjrcTCPvuj9sUxHtEfuIWYVhOpS3JeZ/yENiqmzx3h6Aeb9q
pOnLiLZzaOYx1gmO2LqMaC6f3z124OQrTBidI1pqp/izfoAWMdCcbKsZze2eSybX
dYeNpH8srTMm89VVWuBeZmjv/schTG+UZ5VEuuPVPGOpm8ZcYZZI8sAiQUVbRng6
f1Wq4qmiEIJ5qEIFtVsTlLsY7oXzspKG4BfxUPZxNf6r1asktfsD9h07AlfisXbz
X+jvVYcQFv/4KgvzkrFdsuE03tmSaqAzqEPpPlvzxqvJPbKBBwRKhejNl3gdZqou
mrSr5G03XX4U8GcD+MuQGv3csmvIyuUUjjJEyxVHku0gweIcLPQ9yQxII4P+swpt
Mpq4CzUAeLRkSgL/1mtUyNWZiGz+sfpLo6l2co5KE8ltK8WWErz7TDlWCTjl/3O9
iUnY3WY0Wcwwv+87+ud9XLerUsO0hsu9Z9rMNPs6ZC7Y+yjGzMNkT6Q5ymn3sIDM
Cc+4H0MwGx/vRMPWdnmO+j+UirxZMgZxMYQ9vkjnDmLdlrc9uXmA/lJC/JeNwpUH
2njpc4PLDEJHdM14opi74xXI1Y52L1mpQk1qyyx7/RCrcqkHRt3N3DsirPVtAqUt
GtJbzRMn9ZX714ZKSmVR1KEyP0mbvTcbeBCm102eQvjqFuvr+3KN/5yzaScm0YO2
CpNigpPA19iJbb8c9ni3oq9HMfAaBkdOzFZTARsJFqJQ2bkgsq/+LZzg9eRippTy
blNHo9zufhYnLSM0+xLfdsCE0rf83wTLrYzN9zEzVLENR+o1qKgJRDHXCRizwMSw
lxEmf3B0pDFm0qtEvq//WWc7YfleDZ8CjQZO1CoqYw1so8KTl9/cD2UVuX8oqwPz
Gfho4FrH9OpLTqUFu50mphU+ErYzEuuAf5Nj5PF6Ykwxlu70K1ioGryQvNxVDwdp
GRd6DFj+eX1k2KYbRTaVZkX8P4VCBit9hzB2Rsq+Nzik6sX/hoxgYu+JLZJCnIHY
jA7u6kfkInK9I7UTh2Sjav1AeHQ1/FXhIfDp7YismHtCbD4Pf/V5j9ZniymjIYbb
gRw57kl1vD9toYPDNgpQvGm/NSRwJzMiTKX5Oe0Oq5pCpnqghzzP5J6rR4JChCLe
uaBYXQzX+qkmxEgTeS2hjEoRQFzyWz68tO2w27VOZrWP4L5OKTN61XPYuKdpfdWS
DycFt6MEDUCGmyY+Fz/NxWV1J3D2W1azqG+uFS7wUqsqsdU8AEQUwIPtzQ+A1HX6
43VWEh7SXV7TZHegOtotrb68FrQpIRXs5kUgQSi78UkKeIJVotYsuEsxrVoQH1q1
RQcDfGwJJfdB5SPxNnu7NDvcC4SUDMB04JDOomLkhvYSXfA9T+e5EuwmD1pwg2lI
h5l0J0lBKLC3PIzi9Sqdumq86hqKmi+2KKXZ82YIs8W1/z+uaAUKrJIQdmcArUbm
IgnEzvEHKPkIhF+gArZovMnZ+09/bF/IA1oMJB3OG8xIuXv33uRmcpBQJhHQp2Ok
55RX3W+YlCQc8LsV6j2M2oT3Smw/5/X5H1YGmmiXyqfOEoyBYaqZJqsBFjRAmaxk
jkTKJEChZgs7XbJIPEBo72fnr4Gzn5Lg+x1JTHSbgmrdDF9EYu1CeGg/pWjd5f0Q
mfAZ7Eu3AuDuiHA2dH6UfStFM7Ss3xuEhZpLWY5cr+T1WB92ZCFcZD+YIz/cnVmX
/1LwGXDViplvzvTL2rUAHJacdkB/itvQ6YUvI5P3dz80LxfzovkBD0wJNlg6Xa1q
eQKHqNLminxUkBxuz8wEX99OKzZi3M8yiy00YuHORZ6NnhHUDVRA/3lfsg7xus/G
3/sQVIUWw8+ovcGkNeUtTr+mFuNSL53n0j9FqjtEFkvU9V8sqSwKd+DnTrAVlXgA
hBkZN+1GvP/bEWE0EUY46z+9gzjP+aSnycWhlcIUaAAq24mtOS+Zd6Ob9bZWYu8l
JTCHi+jZDQWIG41xHcrFCMMAuXFk0RncvbIqA+ScvKtfd3Os3Muzrud6Mj9XObke
tG9oHXNDZiUSg3ztx5vA9mtHAKb2FxoAwo9TEx0GSH+Jy2Q3Rvigr5xk81weEwZe
sR/kJcvHgsjndLNRSdte+mUPY21hmCdLiZcrKifbsYSCyh+YQRkhubmc2rQvSMsP
61XE7QxLkohpZhHbwa/xkS/C7s+MoDM7/2J2232lefwqEEithQ97mZFu5xEPzYWS
Nc6psAgbL6eikuV+238Y3mDiz0xSnaH9qHl9oQygLo38GVTGZX0aobs+sDqKt5ys
mdtN0OF2wHOIIXgr39MTAWukAcrlt0TX+JDqoKlIjYzMw4DsU3NX1GDLfAvpETwR
UibWX79N2eLQWIk3D1fr71GLEp24zEkTyU4njaRk49ICcK/YRWzM2d3Rkz2R717r
kw0tmqPiNHfIoNWqk8uNjHGrdWzHvrHZ/NV1eggwD2ljTeScir+22tfiw13i13bJ
KQwzVKaBukGRZGVYqn1dZl0ccJFYdMDburzW3L+bRpiXBDg4fTY8SLeFBSDpJAfU
jPuKhCYDiZBdkpvCM5B2/0EEhECyWxCQT+B6Tfe5lHXPeHarXgoCr5/PsyVF7PBo
ki9BeAbgIRFa95wHBQYPscUwTrF251bskfbkiB/azn1DpLgwMakXsXnJwj0S3pvR
xBZmPizAut0fUMkw46Hee3klt3NIgY2i/61R3KlpxhyIsrpwJIwbl5KaWnOxQoRb
sQWtqxdlHbbN27CKYTUwTf+a3kNLBah5bPxQ44u+g+hhX5yM4fHDnv/8y1CCTjKf
0WTC8Nqh7ZcZX6uPTy2x765ZlOxQ9EDX+esQXVdbYksfU91ZKS3W+wvjgQKbPQSc
2iTZN7cXKukruiFH/NI8qBajQQD1UH4NW3GW7wu6Rc7IVBDmCs/HJgolxphaGNUm
4l9QXyo01Mtm0FNvaL7o6yFN+PaCGioBVriOSAWeAwEKeHWsDefPXaJiSasSYE58
q6Vv6eayTFKUn2It2N7MTdolgq35qDgGK962UoNUXBRwlcvW/Z0zJ+FWzKxwu7eD
L1c4BCVwz5tgiilmjPIfim93YSOzVncesSkrupwLWFKErPTFAb7tlS4WDdwfPGmE
fZHhycgArP8Di8D+QgY8ktHHclZn3rNM2wS2AjnJ+rX9dcvwSyUT6blnId9PuJIJ
98lV8Sk6eBWQi/wQQryjDJO67g+mXm/phA580bWlzDjCfWR5dfv5ujhHoxOVwt7V
WrMJJFBehDIyHREqEkTa+QIJYsGC2/LdSNIVs6iIv8PaAseD6ECO23B6AlntWmWI
PeWERqvL4QfI0stU605qiHUIemmH3xo+yNVoIRW5IJRlkGQtQAHDWJAiGe5Ty91q
paI8/n76biEtLZUMz7HAfkKkYSuf/dxsIbwq7LnyIjYtWmvGxLvIqpdIWVFKZlFt
+HE+V7N+911JuHoNhLmBviUdRZ23MsgU2tAzrdNhdBQV+W6kjnbdYmh4H5NCuvlf
oJ4dpT0g+/YYKstnNlC8xQw/lrkV2QdEjHcwONmWS9nB06lYOki22v8swx8BjprW
ICW5jy7zyOlLYN0oI0m5yu5WFZk0wZa2i3TKnatSZvenrDu9Esft6tKLNOfNoULB
2iZ2ffPms8p3mXPzsYlqihV8uO+K+CLp8/UiO5T4gHY+HfthRhe57l0+/lYWsUZB
l2f8DDZORJmIS4vOYP4vmRwZS6FieQ2M3exWA1BDM9MyjrHetgorWVVHDgTyRohR
qLmEifHuR3pkldUAZuT43qQa40D/8FLxySWmX94dG8CZkgE71Z6cxLsDhvRyn0V4
2EBJcbFHMB9zWKK7urc9utckAPgjhqKxla2iKUYGK7nl8V9bORcsELSMGWf8Pnnp
WSQyGMGh+EDU0R/WQ1eQKOtPHLdS5V+62U8YIehrThgLijOmgCJR6YNciR6A2Ccb
gfC8Wad9qg2xHlSvk7RjtT4SOey+V0KDgzvxD+f+25LI5z/ps8pSR0xphek6qC0j
eH6V6lVyUygCwjzt9tn5GEdmL4guRdjLOEGjcs6eUrlujbGf6QKzevtb0MsR8A3v
V9Gb1x5aMCMgYfAhh+O/uuejNfjdwtUs0tqCKNhoT494Kt9RbMCNd5hcS0DouFEE
AfDK649PgZGsIb/LTWyNLiT1f4G0k3wTfDUYVU0jmQZehse7lH3zxIqIGKMh5Wqe
JdpgM5ZTjt7mmw5lC23NjsCjuU6EujzebcNPnWVDZIJfEz2sBge/fCUDx1PbW07K
ke9EfPuhUPkOpXb/x2DHzKoAIPEQQohXnDub7U4vfAp2n/AFLy/7XJK+g5X/vveF
GOgnkX0qm3PedgqZmgCg3Qeb4ji/1vA6W0hWpxxTYsTiLTSvjJjjhkoKnsOLqNyb
y+G/NxBE03k6Hx2eT0tMHfywYtsawwKafqJGOKjdaNU4mLf7TG6FwPfLFBuTKbds
LQHQohQ/im6Zcs4AeuXIKv6hwxf9wG2RCNUna08ao9/K0CD3doe2OhAoVhSa6u5G
/AtSJM+gW3cHu3j+NTUnugDqvfmrXtaDMYrQIO8L0M2R8eyX4jZHp59flvzX65Eu
hyeefNSxB/ng1TbRALCLFK7J+DHQGhs3F+VRwquo4h48NPLcTtN7X5g/ZxEgsKMZ
ptwg3d6afgaEyi70Kd7KRosb0LNb9i21dGOHFJioJpSeTU614Hkqrv/gGuxkpYHj
JogvrJJhgR/3b2NKvHAdnqZKO3fFxPf3EaoVea3iBwrkf2wf0EeiW3WUkd1bkIh5
YnABlSUe89ZLXSsQTsNQAKnCaokSq76Du5Mn0OpAJDCAjxZxMVek9G5YkG5x7AIy
zjcNtsmS7pJJJIhQptJmsVJL62vjk+cYejoF3PgMVTCfH3OGrKe9itpP9bQNO9Jk
G2loG7MGiDHar7xiWuBFONhkguyI0fqD6fLHfLRZxisxMzUsR3Hojz+Z5C+yvOE5
4eXY/+CrlvA0+mxipNjQdlap9Ezbn0qjHC09zYwYjS2p7sA+/9tWrfCs1wcIWpWq
foUybM7fqcKgzvFBioIMoQkhEiFXBY3lpmFHvjCJdFBN+Du7g/EnbDmUw2vU4+72
HdnrMbGnzZVNgmTqeC0qgE4b4ULOsxotUUWAe7pKA5hQqaPi6DgcOxumQD0tcQQA
/Bwe8c2NAnrQf1+akdtvNQfQL8J8H7GM4mbCo6Y4uklCgeNAb/S/qyYMX6oObLPv
QbeuYjiDhlu0vzZKY52TvK7705ce6T7HgUt3GKESScnP2u+NcLujYS5ePyjw6Qky
4+SMXBXPkkLGWODkMvpyQxvzQfB1epC+ZsIqTnDwNurwtEfbpFZmdlZM9OxS0M1U
us1U379dGppl4ObVjNaKYHD+Y4KxiPgjia7NHmGsBHTq4UTp6jYCwaKGVjOZttAR
vd3X6Z5JYFokdYc8dRc1IQ+rGAvZMUNqzAkwMFMkEk9XFOzEKxEQjsytOSkDV06N
aWXTNogIAh+VVsp6CqgOyz1/bNOCpx/3NuezLnbUY1O4++bktpUyezBpN8YWcREM
/k0A67xAHMz9yL6y3pGxtDkg2oTkFDftkW+GvY3Cms4YupCvmj7zSn1f7E2l43k8
zcPUftRrFA74ybxfPeBby+HHyU3yTzVIr4tJbemT4VPQQSAGc5nksuJTPheVB/1w
Z0c/DTrNT4TgmpQd1cWkqzERIHtAkpx5WnzCJEnmVLt4Ivn06/SM3n5rlHUh06Lp
XwlIsXa7wdb913C4EB89ZwVibd1a0zEpKvdvliRsrrKSsxCN63ShovL5AzVGnpoJ
8HvHx8kmBCmaYs7f1ml9ps22upsudqB1YLgjuEpGJsSeOmVewWW3wqisr1eWRHxv
X/s5krLxGWz23NcaxxsKXhTaZyVZaiNCJUW28z/86SXdXqbXjYqlRid4xNLumbj1
ioS8hb/PQMLjmmZVO8syiXeGksP4Nsvd885nW+4Xc6rVUkRntu37muYaVeQ2qscw
GM/qbj4TklX8nZCrvE73ZTS/WYYBOhU0sj21aGQgLYfplhrP6j3PFz5otSUZw4BT
UD7fdx/XsIvYaJlzMrBMI37NufQms3YlFG2ZP5+6KGrgeq9Z7j5fT0BlUuuRM+bE
S0DMtuNsp+wZ2wCNODSNQJUrOwqcVS/PCXRwoWkJZ842qy6knydIOUb/mIF9bTa8
xkhTkXtNDIJ8FqOy4uUvNx+LX8GGCIEktFh85g8nVI4VyLKVGrIso3RkzAjZOuHR
xwBpPEfxYUrclBG2y38aDmAikJGiZq3XYkxCfe2rgIIZE7RkQo3F+MdQHhtZjWXO
PY+G7zqt+GGKpAoRe6St4JgotrKSKeD8o+McEKF8mHNnuXL91lDMAipx6kiUv7B2
XdY4sYVBDkjrau0qPfAi01gf48ywWj2jY/wg6LzHtx1CZmom9hQdU1m3uJ5KWMOm
utClytlZ+xiT/L+s99rZl5T3BFu/qY4cdhpShVmmmIJsTYJ6pKbpjCYpiUr9EIzB
uP7ZpjH5PGVwjVyUK6GPPFLNhU8zHJoKBzmQ0icu9R0F3NfYUbfCm99vj5q/DAjc
eqTXWe1cIFNluTmzYKoxH8fhd90w3VQTLHbAOE8U4nXKPgD5SyXGlcquBuH6Bjai
sINC3tg8g5Q+tWViE5aHd6C06+E0zRvHA/1kuZ0XaFcJg5KT6iYsm4u9kXgw2pII
tuUS40Kq/VkTg9QPJTb2DNcE0iC8NhpW0Dz6i62kfySNurDFqnEYl1vloPkDLVE+
Cy+/r7MxphY/Dc7FqMPLN8DOK6ZIWXgl3nD7Me5Hyc3xJlc7CE2W5F1fV6PfLjbH
K0Vbe038QasxRwO44xThdkhyATHtsJqiGjUH1HqAVdeZALLnh4+X/spe7kMgoLxd
/wWeiWdKro3Hfo8U85UkfkWpadPkVAJwCOKWyIkGQjeKKw6J3jQhE8OkXrJC5q5Q
gVj45YlnOPLCQsWX5Kruptq6BuDOav14osV60ed85yiEvy7BBdPShJQK5SfnzOSO
PDSHpzZBK74QlxdYy3s2KHhwtBjp0Hw+tvxiZ4gGasHLYNdGJzDiF0cSxoLVvM/e
q7ZDe6ET2oPlEtV+3tcVDXm7J1T2QuWOYNTMsQi/t7FuuLtzwlaykZy5UzFRsnxq
93jNC14zRyxuZBEioQgVWgnIn2G3FBW2oOjRhaU2NEwd38OWdGhl3KRrFUWwoCEY
Ogb3E14RvUTaMCRz9VlKnpYsEbBPbYQg2ODdbO0dpej/xm3dWBH58kOOQHCW+crY
s+9wL+PHkdratmTvrdVfYBHv/rYSeTa6iTaRp5zkGVUeNtysFc0W9O4hxQqUwD1B
2qnSbQO7zaS5Kc0fYUKRAicJS7FPHA3K9IM5xLf2Nor7Afvg5cXGJZ5JijvA/yWw
HEtlda4/ZR3yZxoMT0TTxIsI/+Lqn6yoom/9ksJp0NkHoenIr742wQro9cO4Luuj
vZpKk+3fjTnGvPnyF7sz0Fn+OBjX0wW+XC0bxRyKD0c/JWJltrQlm/xbcx90GX8h
JxyBQx1fTFt8WDJkk1YAv1q4QcDcHzm10vFE27dSgP7xt3vPR08pY3hJUk/a2HD5
SdBJYkeRQDUix1SqMcaMt8rQCgEhc87PCRGu6QvzciUqyZsfjg/SowveYG8bPGjc
5xnp18ZKIYLBIKNiLurepaGv+3Tub9JIuSqXLjn17aX5lnhlRp8t/Zm/uSfCDLrF
eoGP0kUkLNR6t4FR1YRkGpRqKD2AUeBi2K1y4KgMS0IJMky01SQF0zypIvjuJCE6
K/2sV10CrOvn22Zh2Ic71DK8yJIVSO87bOCbg4/xqqsWRIRzOPzsthj4fJL/K+Ku
szId2Fo3Kjnu8TjcA7KJfL2ykPaVKal5uNhP5AoVwRCTaaPXxIRpI6men6e/zFSL
r7g0sfSQXsuT2gY5UBlwK/YCikItW1iadHEsUC6AaoTsy47vdKcXSyoYV99xidj+
6ZgTRvygYVmjzDTjr8gMbsfatwShjplGXbkFEugITT+qja/sMso+38jXyClDsNsP
bkkuvGSi5DM4SmbYWsewunc+d46OI1tJPKOpQvThnaG4xZTTHXfhvzZyaLub7YnR
py28PqAEhrzkzelCe8dfED0mIGB1B94IzDUMfdpdVXnEavXyS3WKFY8eTJoCcBo8
ZQXC2fhav9XDTGeVClmUif1Mo5PWFA42jG8anwKl2rwRqi79M700hqv7GpAztOm5
ZHaBu9oF/H0RTbH7MP12iJEJSFh/y5QvKiQztGBQFv6QOm2OupwjgqK4D1kElwOV
YDTyfu3HAdD/5L1d0p5uqJOEcxzNa/HnFdPmKaR2o1KoRnLbmvfHMqIszw87y+UN
gEZDzlFt+8d8AKWbtQqALmqnVubZHS06jA0COFrJFo0o3UkHz89PDNcDgnLh3Kh2
ktK5imV0JFpyAKX1hlJ+5VQjJbjai3RSEkfKdY/33F4UHOqTOJeA4bojyds/TS4d
RqmCsbtmOD2r/c044Y27bfpVY7ZqkH/p7eMYVEOvJv53eMoV/TeKmUsKLmoCCN6P
6SOuCKztS46n7TNo0w0Ti5e0XLbu+pCJ2quobX7cM1naaPC8OphBLPB/BW0QOpx4
SQZP3WueM/xudX2oSBNYbr7kzVqnIIYUkp2xidmAlFQLznqdK6ISpYo970zKoJuA
mxrF2XOQjsnbu37snSXQVDgrv5gdvkelCBU9Xub5+tXsRC+0wsVh13pBTgmgfBih
80SFdoc1qJcqDaK/xfoxaZ6mIjQzv9QMx/2AANf+sRYHlw87I3L0IwIGfSQwRuBQ
oKZWUzJ+y/ck+p8X3J3CFKzljQgfvMTOOoC1fHfhRbYI2JGboLMyc6NSAghuFYFa
FlFvLpdZuPaOjSA6FYNoHKjyVU+ZI5QAsqFVeS9ZSN1u799OMzC02CCsIqD+nxbI
8zNRXUNX5fPbCO84OiWj+aLlMNT5K+4PIlKs2YNys+MP+T2lLBa6AQek+tcW03N1
uZFYUNrgEMIXUR2ziW/yTvGk++OCI5UQ1MDjwJjLDcEpPwPn0wrgXf9GhQqk8kZP
0ME+4O+ntJ/en3SYEECUFQt1yF6vZOhxVs5vO+WkoUoXlgh6uB8keh90we2aKer5
ccoh4BMIwFqnymp4iOki3681BO3xNQM7ZLAxhffy4RCS/Gnwheq7MJbylpFW6RpR
+mhnqusMKmxgmwqyi3rfprgYj0b+9wagnm6ERmXFA3pe7C/ZbkVvpL728ToAYPk5
6+lKD5mvoJFGF4XT4+HqBmhOO1vhgJ7i7igO3gSY48Xwa9K5aNkNO4WjFFRL+jAX
K30lEdusCCNZ0gCx6pb4usiAu/zNITe930D4Wjx8dfSS9XWHoRFd1cCyaT2V4Ryu
jWoln2JkMqHYJ7OmiBD6x6PBZjDC1M3KFGBf8F7WL+UVzpBMeay9lVKLsQgRKf29
jBTnD6CKfXHXKvfaPRDPluLSew6pYxQ566Yi2lwxZGz1uL42WE3UX/wtKWZl1xKG
vIWm0JHtLLV0QGuYJ3il+7vPwgBw2pbv+6W38ZPOA4Mm0TM2acjajcpFjQsK9dKL
2pkT256CgX+l1E4Xh5m6bTHl0iv5P5YxxJ0O+5TISnLC+FqL5ROvI39LpmoWxyot
e5a72vXGb+1OJA4wZXgTqq5tOwS4541uJsqTFRmN0ojlVyMGxXNoGQRt32RW540l
hrKbsUYs249GrisLEaXdqP2kpArfQscc7LfiFNvOg4LioNAz/CLegeWIF5p/ILN3
7ZTQkMHYhF/tpG0mXYFFj6QfqKlIw43dI2tDaZh9Dgl8Ir05+pt3Pj542dF36doM
asq+Q2dOzqigz2RCK+jvybNSJLRRDUxSPeyCyAo3g6ZO1m2QFJ4AoE+fx6/EZPbu
7lVgMNCwg0jDlZ4dxhJ4UHkkWXQ+96T/L7lJFeJUxPrdj7hEP6Q0bt7LxPZ1Td0e
yZe1s83OSsTzCUUynk405+TQeP6vTqJrvftRrgMjxYg/wMWv+oZ1gzdPAaAEBDtg
rrfTs2iLoymj9ckNR8gZjq2UT7NiSMgUA9aihBdZGmn8ryKKllpCF0FSHKGzj6Db
E6qxoLhtm8oJhj6BZtewo3Yq6rxEzRGi6OmEN3z7PfRmaiZnyOMvCOF4p/1wyMwJ
ek/ECDO9e5vroOG3tpaPvzQzZc6FdYKqVJgjujG8y7x/70Ga1LrAErqFvq3JdAfo
6Al7A3cmmm3+GESGYs6dhzPi84ceOpMeh4flNiygdIkqkIwRW+qxXSSFN8eoyNgR
w+jvimg6YnmiYxnVsSDOvomzvhGoT6B5orcMUwlCWaXCzIOStxjeJaW6spxf1rGH
mTNvK0x9BuVP9LdNU+JG18Big35K3zdZGDQ8P8SbYjFQBopsfYpvFMlgJV7qJHbx
SF2j4st9YEyy66pAE7BhzKGJ2RZQYMMwon2PkJexBeXQwB8x+my/vRD1u/DuVdh0
SDQioklbV7iTj/eJRnNimOO6dARGlK5XuDRcM32EgiBPGY5ueM3krWcPI/75226K
XzpzVHyrcQst1+yWM8UEOrC1P9RrNmkJjJnHaCMivdbsjqlCdtrV+5DaNKSDW4pb
59HWfcQlGyRpK1u9xWG5qFJT6vCPkQyKcReeNzSoCMAYIscvurGL9GcPv47x5uu7
BxxosnlY74UtW8bZhIHCkmnQnRt9J0gzJEeZR3h/3WIoyHm5Y/RPL9fd+7Ni3X/g
dtBg2AZorgBVUFp5xX362+6r7UAlTtcnIw4xMl8Fbu1ifTy14YDuy9FNHH0yFWrY
pxdXi0/LHZ7HDJKnP3NivxTnFkuPBPQxtha61iFhAFVwJCpn5Bzt5US218azol8e
VgPLzjsAsb2DOaDiWZgM6/88jhyGpXv9QbyJJ+GgpO7O2RTPOesVy1LXF/e6ZS4K
z/i+G3CmSji8Dhl3gt2kekkqU7FA5KbnVufviWk3byqCRBNNr9eLTrKfvkpxLCNn
Gd+d7O8N4mZ1saKMC0X5HQeYEF3OhBcryhQTm11G8xy6u3D5qUMdxdJqJ5eYSlBU
a6SXyVyzVH971J5n/QV17YXENfkE3lC/dWqnhlbogD9MlLoyoTkmkL7F9Xta3Oxy
OFqOPOzydrSJdf6zaIwluCrUtgfM1k1XJnUqYaP8l5uKSFmRNmBvcvspSm8FgQPX
w6yGLifWWJhXagvXJyOENUSlREi8TVkpFLjZE1v6jaoJuZi25OSr1U3kM5KPUsrK
0Odduj/880Vnssoa6T9wZM8kuwWXC1Dzf1nlEdGVO0yAIqLxSGICj426GQeMZLiT
JhtOw0SySq/UREQg2/DumZaDXEV9FubWpPWwFueOXbDmK6IzSB//dXmMf8+JGvZJ
eBVZcaIDZP9hWCqv/A34VEOHKCy82WdMFFGUxkBkp3F2aDPOdGVpEovks0jPquLm
aX9f9sc/2xIr1DZS+TmZsr6O0St/F7GW0fejhB0XbqqYktaVJv5uZXdYfKizSBrK
8UzkQ/euYoDlPzD6mqO0JSvl7sreXnQieGFGYiui5xgQTn1RRpK89YO0SwY81ox6
+TKdtcz0oT6/L6PnvyhxdOpQ7dahfDz5swIbEaVWqco27HpTF7Dhfvrtu/+gAB20
40LGGn0gsZFrJ4O1gUbxNpDmBNY94YLzWR/pACRRKsb+ukZMa7yzaSHzwhEUFocE
rOFvZDREzU6d4rcLG64MHoRizTE5gCPFwV5JNL+xfg3Kk5KIVco0oNnxjTNdLBNk
8RH5fO1sy7bMfJLnkIwtLktewcmGGzDAVqekE8rT5vLZOF0Is1NaNmuqmRN0nOhf
IqBBGBuJ/yaoClJCt/u6okMBn2Rds9mMImEpbVHOdU8wTN2JDGAksj+bOCcD0UGb
/L5tJtur+nbVutoWYfN89FFpPn1cFeuZhOsC8heVW2OKA7VfQRgn9qhOtjZ6IPtG
fVmzCY+fUiOvuR09sKfIVPdlbsiVNNMSmHXzk6pzB1clwiMGZkNAtTSfG7zRY3vN
VrQVajk+4kZIdcuDqG/U8g3/kZH6LwbFJs9O0qD6Al5gxVNK5A6v3P+jH6P/Un9c
GXwzP0LGt5y67xSFrlIjQ11HlGjlNhNtrEusOxWqVKa/8IWdBA+GTpz+aYNtmhvf
01mL5xzHNDWk1AjSlycQNBEcF94inU+8f3/Li1eNEu5wgUh4FKW/KyfTCincgmQG
4pEoDNdsb8uT4zXmFlxSGTR85Vdp2FSkbCSF5JbCuRQ/59PskbW6Xz5qXf4xr0fo
1f+KvFT6rwmrEBe6XoOxyf/ub4hM6q1nq+S5v+caWmLH5GZaJF8ovCxGhptiApw3
Rxh/fNeca9Wjh5wVrqdaYZlbTXZkz+jeaf6UB0Xdlyqx9645UA9s8WR9Pfzypm3n
mlyN8XFCn0ZBLI6N74HKk4+vH2/VwpMv8MpTTCO6CWwlBH+G7yWRWztrzM879nC4
uewPDqOM5TEhTOVmkYDuNwPkorFXWmmlXcfj8Kylr8Ap0SarGA3hrULxtB9MCokW
+F0/yexY+kesnR/uVWRM+ollH1dFPk+hMcnTvh/zcxdst0jha1R2adXuc63zcfhD
uLIb/Eh9Su6qX/svquVprDrsAppvXhrdMfbxouw2Aol6URxdO+4e0O6bah9PgnzJ
VjeHSaecQwznPjuyF4EAkxXSnv3rtbyC1U0vsIH5BgDng5qumXPDxUTYbZpOTSF7
f62Nky3oEXA9wRVb/yPiAMuPbamplP59KSz7Rmqn7VVWfj7YmwsCyKt5u0aMDzMU
d4bGufLQ4qvDkeNnTepuzp2DZvRTq8dGRWmaHw/TMQRFU0F3ven5RcsshD5TWxqe
FJy8hzt/DiDM47IdOaKLR4vPbtWXnrnKQs+LqpKT371H+Y4Xrmv5mWMDlNxSVipl
2d/TjWyNCDNBQUCX8Zs/gkoxPjSHfZEomVItxEin4+NNp6De5cacBaPz2EmZVu14
SjB9Up838I6UZ30l7LJzUxYqyAexsT6yheGI/xNjRJgYfhWOq91ZeBHnntKKIGG7
4GHF2qY5HLcyYNLzughZv6yHOamFy/rj8XZIfrfNsA09lHspoeHplHqFD2FDb3Mx
9G7IRw775V+eYdV340xbTait+G8+issKTeOektsq08UgL2bgm3o1/upGzz7fgLvb
IaBRNOFv2ckZsgSAYHktYPrItaEyNcfHl2uCzhnIa3+gbcSU33+I/qL28RL+dUwh
lWoIrlpg66S35wOFFGDMzlGhepH0F2ci1pV/0EKnA1bwUhieJ03PPRRevvio7ouE
Ds3rsg4JNqtkt8G2t6V1/NnQ6vrdU6w8wiv9dnToFiRglNRhUmWfNSbYM4pCMvWU
lkHxe+M2P3YKtkRyZ5QjixqcxZNKLwnG6wbCiK58fJoJAOcMfp6IEKgyQqofnXHh
A7zEirb1PQk7GTvBNV0gynyWZb+JW7ZVNkqIDkrKWwe6r95V+RiHXdAQ6a0raTjz
QTZLKBu10sWO2M5IYV+/FJOT2Ma7KZTTHM34io6mchPxDzjWCMWVWSW9vTvCWZQX
N/pHOm+5eywRD1yxE399cSKyYVFYzN0b9+l+22EuZuEWlxDlsFsA9EJ01Z59F9WE
zyvyJA3hzYnEq6U/Ny9QgAZORCvG7PkNF0wn+TvTChHzOcuMWQWaHoHl1kIgUCZl
txmDALrdGKdIUvTdIwWE+Wbf1IZ7qiprSy8J4+przzHHPoLvyf8pPsLo3wKYMrRd
44pRKAq7KgRy1qNxZUUyUGQNJ7SXEcPhUVppsf0Dg6GJC7JScgO7iF+WPRWCKG/W
Xg7bGT7shHDZeNzRWLLXPc41vb156C1fIlsI1Nnt93GGW/ysF56tahCOveMhMkSu
3pz00qVBG8JOaZM7V6heBZ1msVpK8wls5qNF6ROQPlrfrZZstDesh/Chl6zTpOu0
oa59whE06MSqj07EN0J20JhmYVSjIn18o1bmsWzNTqRo6vGGrarC0D2vv0xzERLn
5jZJig8Runr7lebM0T1NjAcYW+VUlct6bDJF5FyKMKLwP7DmWEgwz3ByG3TF59AS
W/GkFR8PaPzbs4hxYMFABY0FE/4novaIV0Ai3ZsKd+TUPvrdEBOLgIQGc6wKXAEB
UhCbTRIbsMbbOZI4GRllEgZ6xizQvuUP+ItfY89xDG9kP8OMqvkB8dRakwHpq19U
+XuOBdcWZAOhY1a0/ctauoI+bahaRX24HfpIAuPYr6WWxJfYZb5k6HxosiS5K4Xb
6H87O2enlj8TNK7JhF0O97GD2QXzh6clfxV7j902aI9E7K6Op5kkigaF0ty37FIV
civjWJnuRyYl4WwQZZCus5IFvheg2zcxKIHRpUl/nGpUHb7YTloZsgNlt1Go26ob
/lgfK6OqPcu+vMJbzrzc74YnKvjyLs2T0cvQ1sbsKyL1ZyUBnc35zLbrc8jINdSM
IFc0RfTd+k7PpYXjsU3xPChlHu4ySZkXwFKr9Oa5ZDAhsuvnEhogQ5BvG+txabQv
LSW24ekaTCYVAYVjlKYM0814CPyX0n8Vcwwq+yEjreuGldmIMgDjLIvyf4Kz5/ii
Zl+R2O8p8xA0tO2lCUy/29qnHqYuAlYgi3C0rIrx9PHn292VdE+ncZL4eZJ6Im/2
oIaTwQqLHsxNbm1daqRoRUcyqSn83dyacepst2+mZD3vTXLo514KvUvV59KjUDcA
Sb5e3kPKQFZy3ib5cKAQzBLO4mlJApXM3QUe6CZym1jz2RLbdX9hPJyNpnm+jPYx
4by4bxKFnMlxvyINxMxH/0h4So0KWI4oEHFz854dMe0I0h+FKDrwL2JAx7tTTtO7
vP3RSTJYSvx8JUHD4YBqf5rGr/g86hNSRG56Q7jP+FZNC8ecLR8RZy7lyAiC8YfX
/Ty7KdZ+nB80TKx4ymlSPo6WDUcA/i9lr47lbmuXjhoIWgHu94HGB7Rb79vAIaJ4
eAI1dVT495CoqMBMkLhOi75AUIuH5JXbvBWSt8hdHYJy6qUHRtsBjbv1cewNT7FA
uw9UYRrN+wuzPTaYVscWlWIQs0rwthhwkFiwpccRxTLrnFM5yKa9uZcWRUEL6UMu
OXvuAGwv9i7gxDgwc2jTjYQR/izC383j9cnTcfqb6ygBcB+Ff8akgkhV2f8U/LzA
2FdxRSfPvH8XImKCirLjrtjWkTLGROUwED8Wo92YxWzJX/F+IzFJGvheid7K0EfQ
N2DXXiCrLw6YfAI6xGmmfARuKD/2gY9KEY2UAl68kpSY+O/eUkxlz5VhzERJQI1O
Uuaj3jfxPXrlw0cSMTP3PF7zib3l4+rNp07X3nncZ2RLGhU6FKoEAVMfziYEBdSD
LRDNYb3pjkI7I1J0d5IhyFvjdFNbPKKBKNUfiRn3Ll9BIuiXR4Z4sWFBKgofFkNf
YW8MSdM8EAZN4FfrwIZ79Dc2ggpVq8bHD5X20u64l8OYwZqa3nY3OXtuAdfEKxJB
/Eabf2ylIalck6icVClQX+HOyhQbzg53uKaaata3L0qJ8G+pG5jykFrWgIs1UweZ
GQmghDoFcU+goC+6f4lRtLFDIoQVBgCOqizZ/CwFiyhCx4bNNiUdmtrGA8L8CLgL
5Jjsji1xkuI1rDY16y2qLDJkjMiSIqd/n+aYWwI0atXkuY8o82u2FZr60lUPPQ+0
lLRcBYKE0cENiQ6qqH7aKol2TPlLCt5Km+8VFZi6oV2ICnRGfr5B37njrb9M4FBt
sxQaOFyFXd1qk0T0ChOOB+fVW0FoKrRM9TObcGTwP9bJsMXtuIy6rWyVKONqEFDs
YdUpoIS9lSb61gyIG3eXTE7dHjLcmKp9t+k9hPthle+OqkVZfFXgKq20CJjeuXGp
NAg2CiwbNWtIMoy3L9j/c6ru91DA866H1Od3EiT8JY30hfYsSOo4/w3DOoeSowEi
NbYYsQomo7QDn1dur/LJ+LwP39raYO3e9CrnZYvAgemb2++yPzS9Zklc3a1JGhM3
p2peq/jc5C1IKzMUTJWZg0EvamHIXTqPmLgBqlqK4WhniXPTBdBWz+iYfJ9F/Hr5
pf/FTQYe+eTyaYvjKnaaaIh4ukc6g4zaqhKvGHyFRtd6cwrARrp7noDPckksVGLq
XgITeK8a8wNpaiVton/KyH/xl5wxQ2HK2QS1/8VCJP+sbAJvrjKwTuQw8khu2n7P
ZUfyeYcGL34oVfNUaLGjDNTuNNcRgPTcHeX5czNYIF2YNED1MrfsWwYEsndbf6n1
rmJ6roj9do0QP2fmkAkP9gbuID83EbOaa2BkDCqSDz59cQhJ4lU3k5E3qGPNkabC
Io9hcHzWhGvDKr5sJo+r5CdYcleI1yBTuD6/ikzHEMrdiJVV/r4tVRXN3Bqw5gC2
NY0Y5HrThzf+fZpJ/5z5SJzhRol8hCP7vbU9ikcSNoYFt2Nr6lEmV5TIosb2WYHn
IekcuoxkyFvHeWOd4CIrvf6DM+dL5fnUtIEZWfqvaJvlLhUDxJt6VFVN7VoGLg5r
BUO2ezeAYjrauQp7Zkgb2G1Sz4q/1ZyXcZfZwtXHZm+H+KivGpGUcbDk0g1odWoL
tjpHEzI/OVb8NEeq6gSpaTmhWzGctLG8WI3a2WFH+42KSlRswnXzRC02CgGWH6wZ
t/UYKa/y423fPMf8osL9dLm5F3cg89c1+CxhFsvNT5btQAjLNUexmf4gv+xZ5hAr
WxTkh8mIy3v5nLd35lyCtaAlVFrkbFLJ8Tb1g6bFgCLsJfx9wq5W4pZbqLNKR0Wz
VkADJ4mIMSwPLTKjHpvxe3oSyKpuL63xJgErS8XaTXiKDgKCd9Zcxvd1AsUvKrt1
RFQhIB84SQB63UrLTekOKSx9oJfLPIk/e7rL6deQLObFfMW3kJCRx7HKLvGzMcVB
HveAEg/BkSU4D4s+48I1X44IfcNJWveJZaApgrwgDIpqUdNxrtMxNMbkhpU4M2gE
cKaMJ0+YenpWZjuZQBl0wHSPnHvGAfCRVQxHGCL1ls+z6c2pN9h2P02sse2RpOJG
tpw524FERsulGT0ycq1TroNvsnkRT3yrtd2T46uE6uVTz3QoAeKtd4U8oAPlOTd3
DqqJitOlMMfU+HB8zPHCX6oWnXiLLlX/gszOj1RdOke7yYH2SmfAu+jK9iZ53zG0
mzTufKRhhLiJWba+PwA0MUzZI+S6AxDGCPEkCo8mmQWT/XOZyQTLAZ+woaZCfUQ9
jOKReNkPVtMBNDEWVhPoTwoHMVFGxC9C/t5f4NyA+7NZnoL1csgOKfK84e72VAMI
t4GYSWfpBx12Thndjj8zt+u4nVezu5uoR1G/lgXxXZn2cj86MdDZokoCo764RH16
H95SLZswEcmiT4HxkJtBiUMImjE2TmpsDJbcKlLkq8ahfzQxfTiJ/Fx6SQrbApJu
J01B7CiVxYvMCdcNtklPSFhQHkf0EmAO4lHW1zuE8A7DERafj15zvcztGBaP7n0y
XKezcT7uEiDSY4Lzy1LefpMNYj3FrJpFInUwLKlXHAFxo8vajpLfcGFekw4nYcgq
Wf/CswtDmAdf2qpv2G4GRPZjpbsoAs0S9DAc4isZu/plTIMSvyphs1OxO4eJfQIN
Or2acD536trWzTAxvzDCbv55pVCOGqd3hsW/OqssrpFwAickLNq2wr4qrK55CKmT
5JLrc+4sFY+ZzVvQmqh11BjoJ5ejEONtgrId9J1j5+BQ04n+nNNSlS/zzzfaqu+8
ZaSPrZr70szf64oYQUfQ6N67k8T7eGg/BFH3ZAyYeGcGo270Sh1rGHMPloFUABa5
oc34gbLvAV0EwbaslconLvgFe5wOB7+4SI/5pWhYjL66LwtDNkAOAGR3JOwPrDOk
bUJDXmca5UDrq6OI4pD+JATDH0eN7oMIO7uxFmugGQQj7r0mfTzIMsdHQ0v5bTUl
S8dVJixlV2eEhFaTsJQS7V1Rqn4eAI8cpbAfvGeFCHmYRbe0+thw9M54ticbw6aa
a2XHI47zcBVgN43VKdLbQg5XXwAVRk7wRdEyhom6x6i1B0lZvVD3Uu+wpgY2BDqQ
mbdPBzsVn/2/DRAi8t85guCDAh0kEixmH0CjLZJaeMboMr+XcjKmAY+wUkuMoprT
JsO+5ubWTd0sqRNm4bS4vC5W9ZRbHdRyuMuyc6LDdXbXIrAF/8zu4mhcDj/YOW9G
13YAKwWo7CkakOVWnNjwTRhv7d4VOk/gnzyNQ5AuHeEvlvJA80x06nC7+nsh1CUF
QpbgpOfeYzWmHcvNMqzZUjlqqQRzJS2nlQ90QjB8XNZRonjQNdoJ2w/YCLwTjlab
Fo+bI2J6WpoNDldUJBkEjOeClHn0bzfz4AYOHllFehyksEFb30hetaXX0trRuBkE
c3yyr+K60jz419SOCFy/B+n+rFZvii5VbKGibICyEhv66pOkqx1IVbKijQ3A+W/+
faCmiBew05wcYwDCejVSw1IPNPeI7ym8vJiGcCnh+bvaGsbI+lUsSqgkbNJDeIlA
OghCFe56VeCYMHfbcugS5GdvQ2axzsi4Z6O/XrFc700V9yI/NIDjLWC2xh0KNIEG
23qZgxl8eRI332Ua/9QGmh8HqBn/YL+Qxuu3nEl/41X3v2i1a1zjq7T5TO3pU7y9
sMx2r5DcZiyjQRURWiQmrkPGuBBnjkwf2UfXRKduBzGq86Vsa1+0hqAR47AUvCjW
P7CHZiTA2abYwYOy5oVDLmybRc+OlYIDR84+ZyssGYupvzvI7ZrDmUUDdoE7lJEw
lLFbje5uE7SEYlcJaiuB86/iAdGq+dPf0w36YS80pwzuHOF5DhS7+lW1tV5QYrd6
lLh4mQ9s4ExlRD7zR4HqQVYvF29ChY3f3I3deeqyeFuUiRiPAJsMQGLAR6FSzTEX
IGmy1nEdGVtbDvDpbWbRVH7ZqVFyFWbpZl59ES6D/E++ynF9VEoTKSNK/RyJea1s
JvKyf5GFbc8zpeYN5Cnmfdxs7AZRSdQHgxxBG3OmOKrikfHGpt33Bq/zgr/tiSC8
LajQguXSoVmK6BXLJTjTUlaOLmL0+uCaF9/l+eEWSu3ij8C4Etv6nLxs6coxsmRo
prYNQdXnox3J06LpSy9L3x6ePYK2wOpst9FcoTrRt0qLc386yP7MBnxoGkcI4apL
Ly2OhShLlMzWYLBLTmZa9rDfxG780/Afq26yLI3Q1xq0jtOhK591KbdU4scHTkKf
P0KTRAtbkItdtFjRZD6iKYluiLbEF5+RacfKXy0S1TyGiVNJFQKJORZtpozyVw41
JKkqZIbrHv+iTIhgDPdXiMUQaaPCFiew+XpsxXOizv73aBtCNtBH82lFLVpCHtJv
HxUEfOIFL1kG0z4QpoarRt9DMv0wnCcugi5KYVdPW9iH8eYkkEOMeEF+S+1KxIuM
PsJ7bNIR8sg8CoePZww80t/5opw0iCeuSmKG2KSRrlkqVuTJ3I0ksvo9RhUwomYO
ob0l+KmSgnazBc2VUagnpoU2CqR/x6oZP2NoSn8IhpfRtMNyOjDBe6FCpXsTIC5U
LVjQXwSHvuAz3e7ZXgvcewkJ8q9CUEEjn6ddiZxZX8iKD4kIecdFOpRi7ue7xB1O
t6Vcf1UEr/+i1tS+Z+ug1lIos0GIedKLNc2+G5FSp4Nsc3db2vqdC9spHDMzGLsr
r8/hq+JakIP2qBjPlP6d3EnoHoG02gsqmFHKXlkzqpleMp7C25qGLyWCMHQHJp+p
doLS5nQ6bB0d5o3VihKOAAP6K2Va73Q6yPAgpvEFdGYS0En+htA1StL+5A8E5Ock
VVIXM2htM3LChPzrGAEVylkmeoL5bMhTVsjDzqlX5QE9bKPxiYEwFHxyogPh/hBO
hgLbvuHCSXZ+7jn67BzrhwCCFMzGiE7nB0t8g6iBT8C87Ol7EmomejBEjy1/Ayeb
CN5Yy+jVrGiW0/dSDp3Y1VNFpOuC6OdlxSgnKkoupS/E/MF7qViRWGsS1+0CGPO2
Db66mi5daxBhsNxdOlqPba5S48HO66xvbTdIV1iFEEcvXQyL/jQzrqudcFNhlTR7
92MpNWaX7X9i2hnBXUn/RjeAOLTMkghSFJPJ8QAueXG6fFfXLIFrZkRG4Iy/ZsmT
zloBRr7V56Tix92MeFgTTZeDzmv9R3mdqgRfTIii0HM3H++ZG21IyjSLEF+hiegF
gbqQsviacE13LzmAqIpojVYyWwtLoYvWvc2f4fnsqMd9FMjXhCjH+QaYFGkCbiM5
8SyA/n+Gw1t3DgM3R9AsoHtC6xqnToospx0py1QnZNL7r6OaUdnVRFddsmGVyBtm
9N8obSKzHzucYRiL0vYOBZXi8EccVXErDimIrrKAFUXMzke3S+SSYarK5Y16c8Gh
EFP1TbEAOzJ6H3bKueWxPS2c7/6my4H7CupAY1+C/IEzdB4+6hsQnA2OCN3QBw/0
1d2ZYikXZJO0YGQ+adAwF0aqp4mWY+zJFckGWDFlmblhgGu3GBvVVGFR+1OxwgTP
sw+H/tTteNZYImTrywno4oVxeOSFYcPf+oPjJoGcGM62zsstNqcKMIdYj0+PLNA+
+LtuOqJwIVyfo84+t3atlG03FNwyrdKAKide20ak2nS+vDr67po353KqW2GplbUN
7ZuspcHN5y8sOK1oOVOvcA6+Un22STCYVoK1o77ycSaVbDy9O5UZNLFdMw72GaBM
JkNscUaJ26AWSKexiPFug/GBo5+2KqgSM8OYo1WYJG4Zrnt2iMo/iRC0RVWKFk89
VvaGL1iYYQ6ypPyqhlsSIKZ0UccqEJCi4zqqFxixQeSu9OeTsbFEtJMWsH3FEFrZ
BFs+sfufcVZ97gVvD/qWldrUaxun1VrW2pwYixYdIIVbeUH4/cbKJfEclbBQfR4P
rxEf3P6GhYrXLGMrBdUZd9+xIBV9UJFHCIGZ8dOYqWrspthOsl8h7lJiESc0Sorp
vy6L9BGFechRiUwPZKr79LgVP4RTHyLnYr3ShAXIAAmVQ+uMIFhxZDrOG1+nwF1+
mI3Cb7Db1elAIrAUaJCuvpwTWqdSok4ASISObQdn3rnu2QyBnCUqwRlgByoXk5bj
MZrV0E9s88tmyUbPoKq4bLtpXEBITX4TIbcURwOzYH04/txMzfTV7xDZtEr9vmMz
lFSCPkNUc4baKGhEL+wrvIC+kb8hhgc4wepUisu+fmFeu9LTUJ+w2KEYGhQf1KHD
Fh86/vDPxUjDS4EsGML8KSH7IEfnPMvW0ks3adTto4QWej/YjHcRp8Q818tupsvo
IYgnf+COv8e+taVgk0t1pHYpm/fwnIQvC4pRUEb67pw/IbLaaoxYAGOvkh6iTNV6
CffAdnGIz6AWoVEDDuTlOA8Yxs5k64B+9ZZG7oPRCGrpeEiBIENXXuYsYTVge47P
nxr5jVJHlYZNeHPB1D6CSzS8yPJtJnjqwO2f8TF2wa8v8Jmw9pqtKtgKQ4IIQxkO
PG8ejtHiYcNHztjoKRKRhNiGpI7pL7DIhOS9XUFqQQW0Om+hXBoAS2u/F3hCTcWo
4twqZAfuIZebVs8CTbU9GsHUCcnWiDkHaHG3axOu3GlEREz2mBT45yahXNqXSaJ7
uUmyvH5zqgF2lUXdmlcSNbDdK5Kw9aXpu/24L8xcg3bW0oAxuBkd8ENnhJu5JwyS
6kMF+PICrxZOGrX0dFs2EwsmKbGEItWlUhqfuz7M3Ljme1VQ7yqlxmHijbvybH1g
xKlOaAHNAdF4eHnAOsi9GwsKMCKuLG1+s58oYbcVGX7Vonrwgo+9PkzZ5oogCqLv
rM9SiPLsg2aBHb6FF6hH/Ujom1VyL/Ciz7gJCQmxPlT6gl/J2fEoRnrpiGWYVXVb
UP4pCQbR1YMTivQK9jb2w22Csdpm1b/UZTXqOxYFFmgYGzpUAG7fsJvSRLymYv7z
vtoiP58uETL+2SBsvmfT5LOYd6pbnDylmbqLNsYR4K30Cd33nXsuJ0c6CLR0jVCN
mAyjBdifQ6pqyUuX+FhSi13X44cP34sR79fD+Wq5/XsIYQKodwGgqG0UByNvXxn/
UaBEd14iB6fukLCVZkjAfkaWBT/QTsZ1SZr0tbk4mb9hwGhldfgjbyJpwHsWQtop
VT8fWkmK4EA5+kltpv+56fLu6MfyK+k1WHDBF02/UWjB2pE8do/t62YEOGGp7jsN
LXIaM7HZRBwc51AseA79KMiLy/kmuIDCSdM70tr50xse0BNNJHnDD4XeYNeNoLww
4GrsOzoZvh8a6ZvBbNYFb3ummbG+VVNr7D0zNVTK9IO/LaMgriHWZtf4Z/BVSkiF
TPNtATuWUQ9iRG5by2KYsgaw8jtaGZIkcQxnWa9mUqWjeuG/cLXNSkEsqRvA00Vy
9IbdfOYsYt9GbJu7nLRDao3gnh+Tq9RI84pDJm/r+yAyvwVndecJqeIno2cfk7Ah
8dcJec/F4T3Tlxm1l1JaLD25IUIKhLOP9xDeqPX+aKt4Fvxr//VW3y6XocRpBIA8
ArH4FwffDtNQbYmc/Y9Y3R/Y+8tfBNoT7FGg1iHAccmvrRuaxOuWVRdZ8sudqa7s
8QDD1it+y7ZxcEOx5f53+ZdJwX+IrJZn9ScGyvimvDjzGida3DLVBfTpuRWAFvTo
Z5hJOc0UgCgVqC8WLQvRQQj3vznP7AYEmvYG1+eb+8zHDC3W0zJMbU/NPqqtEM5o
XOzY4jkkrsJaUK0duRCnjQ22YGC34ov38+Q9qgOJkhB1IQr/PBFQDVnayKLLqfg2
zwBo66/woD2oL/Kr4FMmWTtmM0JLNbKeUei8Nx3PXgCwBOyzpvhWqL1kqkH/ZZwz
uToBWl9zkPcFTk0dmWze5IiB7Nbi8OR4k8R990MTzcxGf8QB/fQY6eAVp4DS7KAa
2AicUxdaca/AkWVl2w5WgNatjArhQwXkceTAGN8IIXRbSvqQt2N5wl7ayGMWrUSX
0FTN+0FJUAG4YO5cN6OSHDyQwq+PqsCVI11gcrbgHD8Olav/6tn5PVkTaRa/U4ZZ
Tb/wD2rwheU+ZT3rKoNRClKWeCJz+bZSlW0azU6JRflMqevCFLhx0S5WVLD+xX3N
7WltvIlxKivWexsjfaGouILC2+IUNyC36U5H3hCvmB9GOnVDyhyWkvbpBQ0WV0FM
sRaogG+p+NI9ULNYTOOcTsLKWhholmf8SuuZLZT5g+YCUaSAr9Zhz4vtknOpAx57
EsuP9jLFmwjZNb1xH7vACgMHJkOYzjtHn6XskvyvkDbqc0RAcLaF4DmOdbRGgyqR
vrAe4ww0Ooh6aCn6vV8hKrXnGWKt2+muO7r52A/2i5A2/31FILpnzxflfjmvYaHM
LOMJ6N0Uqk/1Iw8/rbqZfXiAgtqO/QfPGS0cEiaTlC8Iev45JhqUEmkVU0kIk1oI
4lGLEKjoUCcXsaqTs1sSQC36gmX00r+NBgs4djYr62Crl0aEkOA0jESd18MqF9ue
gJPe2L7SPkCBNrfY4BXOhJG6HaLlbivYXhjYAXQOQArviR+zpwDmP0YDR7L6zUAC
0VpvxIc3tWhB3PB6dvoCGCmFHzAqUzhL/pLmvJ4EMyiuzpX5QNX6ZPZXT+fVpok4
ssPm2W/bC5vrcc8p1pCwchBVp5ows2Yf513XhU4WSdEpI4Qdirg+2IQY8HFxKKtg
InhNsVNHuA2GxfeYtajNGH0qHQA+gdUjxrC1k1RjNs9KOiileOi/GagM72OIY4X5
9qtYiY6bkPbUXoBvtznb9SNKT9445js3ov31eYtKKkcgJosqfcORQWidKAg9QTNZ
fhDjMRI1IHmVqa1iyDiY97QiHgZM+dTGBuzSB+Sf0Bw3obVl0IZ2GVM0eXEH5ltW
7J7uFfv/e7RK4v6Lq27Qz1lj42gDPXSCPa9dFdJpfGzneyp5U86bIimve9tiFGnt
+Y6w46zodroVWlynHiT48QTPxbgZMR2Q7mXQnL+Fus4+Js2RPMcwwH2ap2CfN0oz
ERCD6lPbeP6xOVrUlzK8xAwQm7cBTps4ZoeeTSluvkgJJARxOcx4nBbTpFGBcrdu
2FP9BtoH2QgIw5KpGJ/sDLzhfCkcZ1fOT6iGcAMmmPaBiwbmqRJysd6NuV/dN3Sy
eE02I4NERlVMe5E4vuzggUJKikMSG9+TdQMlI63ay3wIMjyLdp8APM2Vv9x5wAP9
4C1TSXFMumNgWJigcxAhAzUuCnkXjuNoIySqx94vtqCIbSttUGAcghfuN6M5hIa7
HEGNeJNPsliH/uSpWBTYilf2y13GbdSQCf2rjkJnsFxR1bmuCaIIVVWFrpN8BzXz
/tPrumuAOXZEUJoUlGNl/LyBOCbCtS4waxuWAbR8eg1+N4yEgm8uk7aS3Ql3ewlq
htXgEvdsYDvK4QVpoiCU6A33kG7/vxGBXmW1rRwGFZDDLZ/Y5gRyC9+/prP0eQ7x
i7kINED9BM+UxyaEnOTlr/8kuZiLMfRNIDO6BuTTDUlPPViKcDKjiR8fp6+qNhW3
WmZWkDQXkk8+WgEwtl8P7cBR1ds1pt3vcsWDPHd8jQ9utC4MST3w2jouFQIevpvY
79p2RBd1Bjlb77o76TbkW3bU2ujgvDbGXPTvQCKKNajU7yiQoTqbOlZSteDZiLTh
PtUzAF90RPdjMLVWFY9GDJrPCFxVcq14Im/+7hkZAKDG5DGrFH4NUAxwrHirp/cb
i4W+DDsCKXKm1eb2lzXDoZr551ficYYeLdB43upAe88MNXWFAVv1DDVZIZkHP9wL
BVV480caw53XzU656OaDS93FpIuO8BDpNY6lvMBWzwfsicFLV8+/WmKqwLhksmZx
xeLsifKojT9+yqllIEATu3Ba/XO1veGOm9369cialWPfzegKKLa9R2aU9ZX5d0wI
WmmqP5LmU0lYWj7lWsvARaT2Kxolb2L0KBqk/Fvo52sb7Y0o1nIZRhyCp09aLrUs
fU4XaYHV7O7fnLlxmWxc2yRZXb0hnb+KcO4V+1P5VLLVkKs+eYDszGHcoWKXuD9D
bJuGzVir4B6sM2qRy5QexuRKXENTAmvIDsGKubEzHwuIaGeRafWoNoaB1WRaK++4
LQ08m4yj/mziekLmLr2JEvxl6AuDl9IyqZtcEpztSylw/Oqdmmc+is5k18+vZ/dW
f9SBnFwp6d8vt50tiFkxv/CfBIs5/3VuiULV7Aru9i/aaqyiqNAtmrUjVVtqeeos
i9bBiHJvsIkEbu190f0CLnONoi2CXNulfhUqgqd0FfZLQ4pzlMK6biu/LZXsutpD
4u0C6Ju2aM9IdzaXJaXdDunW1bSWoe+3SZ1SWvyRmwp8fvcQHcgsL/+4j9wR3H7r
t4zwezlrujPM9cfa677aOcTmVDl2AY9xFSbGfYQmudqBUAUKtz9ycYjih5wkdPSf
1PB35D2hywgM8RvE6yVAgBoKOknsQ5zP/tI1NKrwbf6ar1TNQw3HenSdFr1hW95H
nWcF/zY720fWKoVW/QiPokJbFfrIjZgfONzEOng7jW+waNPJ1Jgsb6DbnW3q5DZ7
7ZC+0zF+LTUAYb5wWw98mvJ3k03oB5l78ISFheC1b4JDPQclzeij45PhLFBnvN/9
GTEhtQladykQX5vJnTHSUQ5BwxDgh3/ogJSIWvvpo4veN0vGmediBJiFJWa/fodh
qQDJzHEqyxHiseiFe3u+dM0/GyTT/5JVI065wsfx6+rRpStytH9297gjByp5nSi+
gxkRpBuhTlSEuyoQaD9XV1KGhw7ohSxRTcRB9Ha2PpwfVES4nSEDIDlYJgT+Yxj7
YVAfFDCDXVou9RIkvsmPT1WioAEbSezaU7RvZtrR/5TVoscpa0vp1ME9HL40H92k
tvHSOD8R3QHk3VCm2V6RXgb6DVBcQvC6Wgt1MOwfEK7XXw12uWzDXuiW0T/O/VIG
E6HzsLpmZOJT0ODA4C5b5+UMpBhG/AywP2FJJfW17GbDi6JJbL/djpvG/PcU6nLf
G1/3icsQFz6jsCaId9pTirOgv1i3M6HyvlUIET5iMV72Vr8od/mvYQBkL99vlPtC
a7+1DZKx2CSpa2g5aonvemBGzM6lUSFVsFJZJSu2vXBV+eJUL3lXOISAG4aGlTzn
Ci1dlddNS4+iHmsf/RbURHLI3fj7ZHqrVxDl+LtWCqkYSWxxE3xiXrKQjalx8V2/
/MMeEWore3l5JZME2KZ4uwGdsFrI8M90LVsOnFPMWAxFHCm0TwCNl4JbcSVRQUb6
QHCF+4yXbgnA9Sh9BhJBPsSkAhShuI1R9cEwIDboD3Sqc0XN0RkhRUs2ZNofoTpb
z3rWVeYb/q/O6uataqQ5pobMwEplCtqLzZxPllTCVzv28fYjq8qN7R7vuu6o1XxI
fkmEuYQpzFOzgO+vfVb9VI1Fznx7/En2ZyZWWNsZC/IuWW86SZnII9EBwUqqU7yF
CIn8NELEOjoAIy8eIeun4MZL1fljObAqLlwbx7SowobMF02+LZrGPEjBqdUriDIO
7LLnqrO9yhS68K0SiAO9S/ljaaZuciERgd8DFRxU/5eLup7xdqNx7eHZJWzgKwdV
Kr+M8gjvYI0CH/VzhzB2K2hPkIJYgr+IJ83ePSi5DkpdPgX2pbUNc5Zh1JMxiOEX
h8F2zxSVFfEAhAYmVAK0t7xlziYsq2qmwhrWWbdB4ZZJmmhNFCQ5jNbsL+kBJFHw
ecvkSXNztrxc4omliWhYGU6DRrFuA9YstdQwwJeTuSA3xDb6AvLPbaZD1j4T24uq
jgmaOiwEwEhAIhsNFuz0b6IU55AtXWR5Ugj+BFfzLzZ2jlORztpXRkJ9BtLxmnbr
4Lt6Pw4WI+Ku5Xa1aq2l1pcs/AbVmZao9QnzBWdT1Vo6/W0gKrNzxX5FltMwX4W2
SsgW4G9P/O9R/rxNkGxXKYtSIsCH+qxwj3+65c7g11zoBBqQbLn2JIkxeCpAQ62B
xmdhgJNCc9ew7Ruzz/u7/2IOS6I3NWS0thiVhoIdQzBPf4D8FvV8DBVQcZoA4PEj
jlgWXaPW8Pxc/7lDTViux9vmn3PYOkUv+S91Nup2eBLGfDfzwVtylPNjSqUF54BE
INT9RrM/K6leki3CAzgtTvM99AJOrYsivceI14lhMdCIG5nCE4mXq/8lEIkmn0ps
enpWD2FpOzuJ9k4H/cgmk+qSnDkTtTTptQe2KSV05pfDTIx/7lqcwVXxqwUKrPfn
dma5GKYXzTmdsy5C5r/LoaBdI/a4weqSQowmJUhiPOj+1fdnX1SHjr3/NP3eiIx1
1hhrclyfo3RAl1S/+T+zztJ78VIYOD7+ooORy4w9oxUYqJxGMcnWxGzmEDJbauuk
ww17+/4E9mQCfw2lMc59QDJ39TCCkyh2OIll9nhPJz/yr6viG3WXeYaDZbxnkk7r
SDFLVOKzpNNuvIBhh7M+Rx1pqSiepI9sY4I5/e8Qzhoup0crCaKHVRcd8Y7b8mRK
4y3NzyPU083aQAGN/jlyi8j0ynGdph0QZ38V6ZIOkdCAag1DkjE0v0/bo7fOBBKt
p7OkZnCbArLjsCtlBuXjKqJe/UAwyVSwYXjT52+paWlP2c6BSYn2KCkLTyl1Jzyz
4I/WQSavctQb+EvOCT6wU/Q5vUu6npI9StBVaOBJkV7pNO5pW567Unbi9Ejipr8c
BcAEqBPjk33snoO6SFd2GvrklKIyYITRVS9V2Y6sVr/RrZV+axZp64RRbKfSAMeL
SXeHS8SZymzmK3vs4nFjEP/BG/EXGxssv/HXkWM6PabQX21boVBqKPdwxKtTBNU8
8JOu4sg+L3/Dj+wWkVhJB3GqW0qvV4xG4yHS01mrgdM1pasjbHvsmvxDutjQkc8m
k8QBOSY7roe4Q6K/f39pKmwn6GmMo9YNgDwpVtWEhmgLOB86LTioYlIfSWK5ZUz9
Wu0GBEzMcw4ZMkwiY51H9LRIwfJtIEt4MmduCl/tEFAOr3hJ9cJnRq6XOTQTHypq
Mthx8Fdjp8cy2Z1iR92zsFMXwpm4gQLVaFJ7jMRTxI2Tbhor5NDOP2EQjY5K1tVu
cDZ9w0FnzdJhPbjndXL8vBKHkuFD7b1iwieg/svsYbggd/pghnCkTvhDfspxGuNu
wQ2u7HFN4fCOUZ/gzswyNGM7K25Nd8A5+G6N8UcTUU42vI3ZtQMpqrOeM2JEY6Hg
vb6hC7Dt93dMUwoR4fA2QphgDlyI1GhQpiScxM4exwm9uVxTxCTsLK046zNBYWrL
Oiy1G3+U0y4sXq7YW2jkF/dT+orcpeevra5mzO2iAoCFN9uFI6Jrn+OPMOpsGvX9
vp+SSD8RA3Xiqo2los5yV1KoEMVU1zmZ+knrX8St/UUBU/ebVSEWaxu+KIOOjKp7
DvD12JqOEaxBm39t3uiDy/2Jmfory45wam52DfJOTGZtVXD+B15mp2ti/etvWdJp
OAPblQlChbAnYrLnqylqie8eGL8sFfcrm0Y28lOu8JwKB79AxZ8SEYSxDgdLD0gw
I3Wy79UUdwOW/0FI7cG4uN7+wnrTKM0nwm9Zuisj11fL5w+IxAQvFNhovBLrsL7T
mNP11RbQUkyVp1Iz2mcOEt6RKKx7Ax1WLMXUnaiPUM5U6XO8wZLbNlQoN2I+LxEm
WTYVh9nm52uYDlvKKeZIIkM7yafkk/ul/ESffRN4VfMb9neVU05RxoX2Riioy03Y
lp/4q8DYW0dpKm2EUnf5lOThZde0iPsFtcj39xoAmpQ4LvosrDZh9VOj9PwzPrHL
84+mUaCs3mYkWIOeyt0ty8pSxfvEcM00cnBcAAdiDFfMm9+LXOZRcY1f4lit2skL
QkrgZTYasBZA3Veu073Mpi2hcaP0DDFpcxXREFCO35DHWvzRhdulUFpDYFh9GRvD
R0XCIcWMQ69/yA4pdVJ64XPgbpU4hxcb3EvVxOUtXwaKa+dcW3fUb7hDqsbPpGRL
kRBqJAJJ/UVb7VRGpZEYOMmj5tPb1W4+eU7/9itd10G1RNyIbSWIpdI/SckLfueq
w8qvZwhhsKQeHeGBfsL3GQ1q2p1IJQNs+aqjUfGnXT6ORHTfaXN7DBtFoTBsEZG/
0w18FAN/JZOUwjHzz3x7u8MTnaOhKmdQs6Dq5lZtWImivuCNO/ok/Q9/wc3IUEmY
WtZ57OSN6ix+lZB4E3jPPeqpX6/lOo6/x8TGD9UVsGaSjSvWBgbzvfZJXJm982hC
rsl55NGFGWuqcbTkL0DkxLgZYRkAFwk3fqEIqTTs54iEjiqRN7PJ/44l8PbHLN2M
cvYRlUU6lujm489XDcuhSgFnQ16UQTd9tinzM72/OKu7iICUcUyj5A3r6uKynsN0
xIY62AlDhb92hc/odmo/A7FOnw7qb2/J1fzCm0VqUNsRz/kVlYZxxxRKu8Qk1djb
NRWRVh4MIlcrzre68xPPooyJZNrfrPUFc2p9JEVgcB90QiJjzIB0P7mFP62iG3wE
4r5pfnHjTaVTWl0eQ9+U6/RnFrloTCH8vljJoiHGLt8QfLGF/3jnuU2azinKJOmx
vCFC983ugqECSiPPyZOHob8b9C4HQQytxzJxyAJe7I4+LDwZtFkkL7S0GayHoOK7
e2gcMJeusaJKmhiOKcRKXom/Elv+bb2+webUCYhNx+cnjM40+OJFZ29PDirUeu+w
nwOL1umQSnp4yDxIz1MObw8w77R4KdiP2i79g9YE3c5bwMnkdxpppkLdaz8PH3EL
I9OBVfTxnElUS3cXnaIOAYu0DJ+op50wcSHP5ScHOvWV9e5fYfBo9b7FfiZWCGYH
vhcg9wDSZj1BsN4B13zokoW/Fc2nOLeKQiSwJJC1EC9yOyuIgs+rmEczMqvkLJ2v
W3u6DPNd8CQSYJM/7gtlBwNhGKNhBeHGkI96HKvJ6E3LqAPf7rSMWCBccANTryuX
fwpdhDzhSymDfU9wl2u9KOtOFA9DaQxsSPJZ3aC8hjRECWKXVrsaqmCOlJeYVGKP
INPgDKT+Fz5Lfr0rbtLfZgky28L7tkP4AJmipmoMvqKsKjsob4zUSxErl2bY2MT7
U7qLRgoQ0eMO4LYU3R8by9Vb0EGgY9gIN9j0p9YDsAg/wDTYRnKLiL2+aro05/XB
bh9TQvobME8QlXN4PgZ5v4iFXu8PlkymTBphTHUkf/KzZjrro6ftIULVJesIe0W7
B5S5iw+v8GzahkS+CTZmaDU8NemS94TYhL4RYxhKCd3qBrhOpagjfcRGpLvO9bpR
B9VgEqM30GpMDmSlccUt+ApoqSJx+FhJD5TJx9BRj+9kWGpyt5YuYjusPnOQYp1b
plaqBVuaIaomDe6jZb+app4MmuU7IJ8NzatmtJgUVSC4/9qnWlWdl+wlnZnGeN7Y
puYqsyzUBckukqLHtZOg9KGwQ3IY1T0QYL6SMZQaFKlZaJYiHC/JiIUybu0hKgRq
CZsHPcyExafMZeo5lmie+9bpuVLvGXOxHl2V7yfgjKbWIfK0JW/M5sK0SFDj0z9S
IbKvsI+9eGUnQTaEjw5BSk2Uw4u9yTuAAX00tYXG8uwmRoz+qVUuGT8f4LHAgJ+o
TVVR8xWuU1zik7L4vWAA9N6VIHK2yZ+EGcZGD3sIExQIgnfdqMl+51WZydMrsyNK
+Tpn7yHksgAgKxjy4k2NTPmAGYjQBxqBujepO5FKtRrqhvObxol7eJli7Tv7OC+l
9PjDL4bilueIyq6Vw3rHG9SWzgaLEikSFqVRkDEfjJoy+lcxbxGoae+ygaliMk4x
ryzNAcrQe0oWDw+GDIX/KweCrpW9Z0+LzyBo6rXWVdt9ESXUqcIp+u9Q1MoVCD8a
NMf+cJ9/AmixVX492BU9vYY1s4ZeLy+nfEG7ba+DXICVoIY5tUhfPOrFMZPaWxhk
XJGFb6HFm96cm1ycg8FLvNstoFG9INUr+2xdQKhrl+EWb5UWGkMaj90SW1watRkz
gsFlw+FTnCi+tB+tf3zWLe3hR0EhWPVgIvZvXnmtuTfKK0HUJXnWEwGbomL2GAX1
nXSTkh+FI6O2k4ZSig0RYon2GvEMYdCCh2NsTJW0zYaDdIx4Ycs4QxYFUEpVdYMw
S2OFSxi/EFqLhKVqtNMNI7AYmn5mwTKjevcrieJflYMNZDwjpillJHUrLofYC4kk
aPLnFzw7YJujd+pfmv3HCcDffMUY/VkM3bs0PAdmuM0yPQCZ9lxYyXVjOOQXx70v
OdXJOUIejEfQsgsZX+6Van8H/5ABEpKZaRMkZxJPcvRm0yVHxOe4fqFs/5/1ZfaT
Twi0DJgLpOxQk+N+yXgu1iO1bxMRvuh87rUKNls7K3ZUfEReeJHmyVeneghqLfMP
XaPfSWb51A4OsOL4QP9lruJOKyayPnGE76V0h/x8ZiL7pcUhCheJJMeLXpKnrDPK
79ALAN0aluUGIP1zNvCwevJkcpKBzToKQ/xUiUrQ1yVX5vJIHEfi2vg5lZs7Y2kc
9JW+ZR32bo33uhuWrZ7DN3vVGIIicPfvmUKbUytko42TdCTshQ5C5NaT/GOuiKtt
3CWZfCq1CU+NR+UjSWPV09Guz+ggpzWlqzz9sdxZNpoxY5XVPxDphkoY0lWvlVgn
qgijxmaBqPv4iuCLnf8yEIbyK7rYEPeiamRKwsJDNCWhf1vnHOT4Pm5F5kiRcW0j
g6Pb3Mh0yRziIgxJEtc7AMbCmPt/NVs7kS28M9IKKsYJ8RpkaLW4yhDW34m2Pa6Z
EpoDBPGvl6Prs3NgWiNsTF4gGwg0C74MErjXKgdygUvaFs6Vj1EkGe4tEp8MVHQZ
jd+uj/KTzrhe7ZCoUm5IqfeKhRnYkWDSWOTjJO3Qo8dUllyXkF656dqJuljjE5Pg
xA4nOEZBD57uvGjZihuDznxAt4OxQYerlMsfol6fq0LRWV6LEp9aYKXDxDqlxR1J
V2Zj9gnfkoTpjXFOas/zoexkydgUhSNYzGHADR3EnoTD2GO0s2Tpx6lSRCUR/joM
RUWpx9+kGb5q/lTCtgj0xsJky30YSyTm+mcVuYFinyqeUJd/BnwWZ5CzMz7bQ12w
Hel3dRO052pEzrIHYQrNshjMAm1ihAzxpTpRqRs3jYB207Kf7+QCJSzUSGVGsTiK
1VKIz0VSSf35s2/+yNCZQz7iNcHjeuQfNHbgsFRaLt/4N4YOX2+Vgn/1Acvt1dU5
VXQIW1s/cbn27T9572lPthgHv5Dwz3QWGVez9X2NlHE1kl9FrXnHhHhEFy0shLxd
7OaQGRNgOvdgEg90QiMWqy5yI45Zf3Dqxe88cq+qzpJ4fJTANGV1ClBK2BaZUVsK
FEOm/+KgnIuKM72Mt+oLuClbX53rl+nZFBIcRYIgJFD6/7CiKgYm0s+xOAZ82DJR
8pzpZv7O1uPqfr3v6e3kkuaPPYFfrZvkJHfwE5kb7MHNoeB//r6axzEM4PcV4Ze6
qgv56VC6+BDR8VyxXJ6/xUyDwpl/lzd/rUGrXMtZoCa0ZrUbV3DA0nbxMJ9Xjcdu
FvwLib73W7LwKXWoQ8N+PHbJtRf2jxKn2ScMxx7aghifoPEsO9TnpvIJgDmZcX6A
hFrIr/z1QCvmQIzyuCiXjIlCN58UsuZZHzOHe+sZKUcmI4J3gcu9cdu2P/0PrQaP
lXs1FNKgDeenc+lM7TJqGs6t7y5sDlkot843BYDyenBxbMahxkYS01PvmmdtUWWq
Dv5gnrFuBz9rLV6OHibgW1GBPCY2CywY8YoELGR8fFjOQ0qU6px4aP/kSLry6FGF
bEAR6SZ/l70J9X02xRGj26T0Bfr14Q0Ig1ebjJty+Jx+82KMbRFSsir1jkhxn7vx
BtjCjzVopetH6ISu8cmQj1YXQv/T0b9xLPJxPenCedGZ2vrDkmO+BjtpBsL8qMWM
IHrbIoKnDuJZ/7GkcHd35BXujOxLbX8DYvRVkDzzDFLtDvYTL1UtrAQ06T6WkUuo
hKMX7mBaFo6fuXAy5KkEgRbbuGv6PtdL1hqusxyN2v1Rv4xnc48rp9aBSIP53DHe
oykoUHKcx0LhaMZiG7sl1Qxzicyt68Gwo8oMWA+ybFjnkViDhmGF9xwZAZkCr5Af
4F6yjrH7OugYCZQTTW+qtngiG+4M1jPrUEl5RJZNT1tYaHCsk9VLsFWZHf+m/HhK
vpMruq/IwKGTlTqeF89yXFiEv37+esMcHEwAdncGL9grv95gMSpBIFpexZNTBnw0
O25KshJor21pmNT/us+5ys7vBurzVt5i8aoW5sw7V2Db2nLyCn72iwtPzZrGGmDQ
UYp5xuiaAc4iq9XAC7VsrQL8Ve8cavw7gH7Epy25J/hNZzz60BqthFqa8OgFggym
Su8GKlNaV4HErAatSBZkh/3Hg+oKmosXDgLmUJeAk7FiRgOe/+j7u+ngrMQVzNPC
NQp5mTuYcJleyhTfz42i4TYeo+8G9fkA4uIEUw+MxuaUh9EDEfq+lYBAXOPma4HZ
+9Z6+JipRuxDZ9BhDUA64484eeyklWTZAKiHJ1YmlAkJWZYbmboKUR8fu0wkxfyu
YcYdC07s7ete4qsVl+FQz+vbyggf4KcXQo3BqPXEsDtvqJfvkXd3OcPNVfVZEa3R
fe/CWwVHlLN+uKXWz/1IIp3cHIwM0cJ80RPBlPay5HxCFkqogotY+elFxZiVBJc5
Xsho65cYD+9H38nrdtjlsK2C+lu6zZcE8M6E0+Yuw/XmMwXJ9kyQsL/ycFNxyslY
HeNR7wCwEOEaH8OpluwpFRvnmslvv7+xAZ094vZdXGWNvLai027pMOZjAeuRTkPq
MzE6JqVIBiDjvXX06FezcKp1J6ydWHMKNSBrGshZBoT59siZRulpL9wQW25HhKi+
Wh3B/wffcQ54T7IvNIZw0N8ewHFS3TYWid3EPk4JAnYyNv1he0TPPwgdIY/CRLZV
g4spzGawyWq3R3ppc95SDKWdWljmN2Y9++tMwFXJ7XrEHk8APQIrh05UNXIXvUSG
rrxy/VylhhjMejWujvwPtKA8Z8aTUA6PxUFuHSIjDTgcmNdWHeRsmI+I9opTlK5r
r+lUHBQRhUlxJql1apc0WFFgvVVy7F3GZwP16faEFsPkQ9CQ+zSajrN319Zb0hPt
izRJYPNPYm6qOj8r0lwnhWSPPrXYI0vdxKpYNloYcGeIrQZJAehngCaKvlQOlIFK
rHYYh57gmu0qSemYdrbdF26TMZP0hnrOc6ULohe5uo+xlhKarqE8FDfchg0P0aG5
clnQ0groi7LiwUnlUPoW12bHyTsmmToyqQ1YXkdn1E4sP2/UwCVCwfn/Kz2/Zu+l
mwOyjWJDJsvGP8IUB4GxNWxABfnzWl+HsVk+yfCUp6TbC3cwf7o/nJ0GifQIPyZo
qyYOmGQKzqeMSYeDI2lrJOQ7Ly/V/kGQpje197dTT68BNHuP7DyrElf7TUzJBfng
18GyZIUTjKnPRY1m2LYwXTHUnaGdyylAJJA6uH+mMCP3L69o4enMZgOEdYXv7mMG
tpbnFLGmad/IWATdr62ktTeLiqUlqlhCVX8rzEIhDifwAIubhGorF/Z4b6y6SArp
poC9+s08EW+rpWHvIcq/3bid+WOzb5pzxmtrMvRG4wpsgOxn8i1jGzvjLfPZ9ThH
XnK5yUN8jKZcH7s5kxrzj6WbO5vT1s0k6el8OvgJsZTOHUaPzsluXYTrsiYCyAaJ
a5xMTF+dH6wa6IVRYYDTHZ9SVGaEr1DB36fnkZt0L+TPelraC1kqmKyb3/euhvpr
VdXttRK0fcl6q62OQqA1y9xfWmOKPjKW/v+wXDsEHD4lS0Ybcg6mcmlyacb/aINO
tLIRsJlGSSIlfT7Q3B0aI2RhhJshAs+sCC7dB2wISNbK3ErgK764SpQiHlxDiFOV
aMQVl6J1MOHFLaMf0Dpr0d1DEerwKhPR9wdajYpFF4rvPFYkt1M7j5Oe2fmEK1RJ
8pxhlFOBRecgpOFlXR/mPeStu9iSGUcYHgTYfYhPtVuFq7hmAsE3MWVHC11N9WRM
N8hZYPLg+3eXaRgpbLkt+y5jo/fyAl4TKWNVZhHUU3DnLA3ZAEXypnOeFr2Ph3kL
kF2oA8LgK8fpgQBjM20wZ/uKG3KORfoOVWvyVLWkykBgSscnUtPt3vjBvjFjTIiB
xISKvEtIYgroXAbKlGvHBi0UIx7kPCUCL+DztdqF9ZO8r0KCQrI/nc9GcXh+pl2I
Yr+SJoZ7R+8BohbaxA+ASqnyxZB01V6kLL2FUVxqvjDEE9mC+S00Fa3KfN6x3DnW
a+IJxAv5hbMFklBXQHC4SuuwTJbOQw/F3f8dr4BrqiFzq7l+J5QgB5H8UCwqpAZO
NKvSuZbCbYXec4A8fyjkrKKhlJSC8jMqKpR1h3pOfCIBuU9bLPgXsARXqg7WnSda
si3HYo2kRnzs0FNAVWVstk8HckYUCOgIzGd5+MKbfpDGkbL04yCgAsM95LmMFUsA
z+dkefgeFNZpE0Mw65lqe1ubo5X0k51fyWt52aof2hEpj3wGLaQshi+DHfaL+N2M
RkQ2N53auCwNpF5YNEf/q9MkWAFy5kh7mFnMug/eolcVBfVXSGY7Q61BDYbUA9gl
+f0+ObxbWeW4gc8e4e62MAGj+yHwI0auG98TjdUxJIsCc7G9Qztck//VP2cAvu1j
2DnqtOS0uMsJqptBZU1e8EWD8EjcxfmhXSPc1j/jxcp/i69G7X3RZ+BE5R/Ubdq8
1n6UkhzMHpdpUjMvKJYOqXaCtJPltvPunW/WkfW+i9WdwIT8sME8dB3Aj7tLQ35h
wwBVxxFwaXlX0AZnXbIKm+Rh8P0qpbmRAMNkQ7e4m/+yqub7u3nbF4Pn47aYHs9G
9L9IWEiQN7sagFvvEFPB6V4qgND9tcrEeaO1BEIQrk/LbtvVYRfCPyP3le10h02o
itZUGE/iGt1guIdnzsxjNIzReRe4k68RiJNLNR6oUOt6AGg3cdFvf5wICU+8X4yZ
4FKTGPB4+IBxsdxGRiM3VonkMzX8kuWubZXML2tGksj1+XDZIg3XBKJIeCCsyubE
0mF6Cb5+ClxCLfPCZb1Cg7vV2Hum5krX7VliDzqwjfVbvBLlv6brh9N2gvJfbDL2
u7i7mq+Fps5taGGTDmOTPAlRWnEvrcFqNXcUUqzi6h4Y6lbJ9TRp+jxlix6fqAcp
mClWMuzbM0P8BsN/VYaYIF0quYxL6UViA6EVgKIt0ANzgOO1vbGEyP2KNl4AiWje
zyLR3znFadn0YJaklOh8CQrE2Q/4AbkQiAIKOzUcjhsYO03zBeN7xZtu2Hpr6aZ+
CFdXkLdcBlQQfvCcnVc0hLDMz7AhR/C+gyigAPVMc346XQIvBbGi86Ec+9NMDwPf
ns4oMV/9T3gkb0mos3vMzb6/f6sgYMM/G8M5jZWGtQsYfsow+NMFLxLOqO85ciCI
fMZeatKmqbajOHqpYlsrPDahqtkyIv82kH0q7u6u7GN/PV5bAcKYt+dwEOiijD8N
x0iAzB8BybVGpt0iIVNmjakwwjZKANbX8JdZ0TZQKnhSgOxZjo1Sp39nECxs4daX
IjjtMB4hA0bR25zmr1o6il89dnE3dmcoU6QtIWuYVtDdIsjw3YYDmB575Ry2WLmN
8pZTs48dFamvC6gMIBZOzQDnPI1NiIQywjCoKkt1NbFLk11YA2pzT9KSw08RaSzw
/5TULrR4YCMI1lBE1ioAXpjqI7UsYmuX4gPEtvxQ8123iHDjkmeLyi+1r/y/TyN6
J45m6ZZN/uKYlpOYN8RM5Ulf5SMdkkIuV1+DvWYdd8cz3W6cbZbOHKKp+zx6MNm3
hnJXBeznhBctW+9L1XW/7R6yai9obRMRwWBwf7n+DWevzohWowR4w/KxI+NdXYXb
Ql7esyJo2S/5hWz3GststUkKDh8akdI0KuY+HgB/68/nFZCvXXCDpMAE8btx5Tb4
/TXCE95M93xmoG6q9gEeXIWuU2h0zU+lqtxS0XlbkIlsVd6Pfxmg7yZeWqNn39Pw
EiT/YKAF9t1RXYoFfS7pwukaaTTCYeylTYyxOMj7tB7qioz5rOsNqfJmJ6wVG5pF
qvgjJCOF3SvNaTEfDSdW+1pgsMmo8NkIjQvhy4EhzHhtI7DfD2hssXsivt6os8KH
nnllaKpMK2oAsSz/RGouCGHj+LH+3HnPsHPvzXPYdbEnvejToyHub1pUsOIteQ+e
t/uTyICClGrVS/QL26a3rLXRCojSyRa7Ox0VEQz+lSIDTDZhneT3+fk9u+vgjuNT
/kTaf/sNjiWiWFD6VsqR1G0cRoK6Hx4lcWqmf97ob2T30URufqFet3QsxLxCcHOs
QluC+CrF5OIp7Fbr8KxuNDLmt/uiCn8/zVxscN+JU02EOr1lX2HmbN8/c+cEt7tg
Hwwg0d0xv5h1H33LiIxuqSzAQgqj9RBYMXYzZ6Z1+1c1ETFXakC5dBJ95XyEGatn
L8qr+B8Eh3jKbnPwMy1YpdEzRITqgAqMPmGAm/vVyZI271zqgsvUsKgWrAeMP4rv
SVZjw7zOYOsEyaNRhKY+ctEv2GirV0v12vBqEerYcAZIoPOyiVQwBRSZSAZqxmhh
XW4AXJbXJTIyFUJY3Ml4/gpzu4WMelYwe4xRKFVs0/3C4IC05aGX65n46TGZooTh
EqbdwbUzFxNW91oxejGmAa5Dy9+PXpU6RQHFPdCD8JiwPDVsDIAJNE+7ZrqgLphe
+Fq6aDb+XLPMxu1Qdv54RVYQicnTI8erV8D7CyegJI335RWVrRqjTIoj73xmhPDH
gdJm7mfVzlS7WnH+vE0pVlz/51uNpR0ZOhskDkOCHWcFXuiCvuYgC6JK7dVLHWv6
iZgDfkK7kKZ+iw8iFYKRYxey+gkxarpKnpp8X11af8d/EvsuCVb1KoCY1LfWEn3C
g4Ez+6C9jRlyfcyv6YlG6IRa1YKCx3iAC/PWy3JbgcrHahysRgH7ZHEoGackKUxt
rREHaQdG1plGxcuRLHbk3pC9oc1YyEmruE5gFA8EOt/ZBtgi5sz146KJ8TYWEqng
SKFt41AavcnC3579y992NDiiDqDiqv4zcPyKEPLTEAZUpRkRWomuQh3nnGZ1y7MV
hpPzg1YfJSpBqMLXFpSFZuXFJqSdYKTZhfJ1kmvKufhObxNb/zdVTmOf8LMETnS9
UvVtrCVWXLQFmAkV4ULQLV8K+9iEmiLswIc/n0MKmjkP5D20UkwnGs43gNR8uaN0
+fIt/yQ328a5Gh1L43nKAr01d5r8TkmaeXnIAcxnG7HLpAKKWCb82zVJSd7bmblI
IaylPz4dOg9cOdZLdS7jauPSx0SKsnD8xAZ2lPlPTgWr52gzXYCTeOazmcPIfEap
XL4Gy8fCsB6BSvaK4vZ3Fxo/f/2Obf9V9eP2hRyqMUJceezLjvEeuHIDf5BI21U2
69x12Op1/vT10VJGstsJwe9goW/7BqXrW/KnEjeEvcXRVt15+8OXNRAW1AxBulUd
+EvFUBGaFfuEVAu+mHfPZhbc5V9+xRlaxAGuJy0QYfxsXxHydXsgsXT9rlSp5ZlW
UAtVmi2vqZiQVh0pJEAseeSx0WhgVdyq0q4+x2o0whJuEU1Vw+RMfsiq5FiYCicY
d8mbFCqSFtkzmG14f+Ey64yi9D8esfOGjFlZWFprpWinRive1qyK632Vt41fESxf
qOFvCxz8hMxoBvz4gqCngufxPealNUnsIu+hzfdyLtbE8pxzO1Odu6cUSUtoTI37
q4UBqB2jYE+5BfydQlqY0rGvur3cQdzB9MQhN3FR4k6MctQZKglRGUwRb5xrt1Qa
gRY9Zd1Ew46Wwbeer9NTBABV9S/byc5Pz5WJhyazedKQlD+hjdz6Y/M391MUCe3E
1/gdtU3eNW8TbtTG+bhCh5m7zakRjmbu4IPgQYY6gleIFfV7iAKJMNl8z1AFuJls
R1UOqGgg5YibKxZXMNFygbzEbOOq+l3Lm2+fAS8nJzZwMELRxKduttU3K9Nrwrhr
pgYhhJuGL8HJ6lcEL4vIUSEjLbP/CC1KlMfGnjQjZ6LNLFdmNqp/1PjCXpiXAffi
4pYZbKH2c+NGVGQ5MZLdj//7dRaxaFhoJlOP3Mj4SZZBmKwhhKTLWYU7Hp0j2rx5
L9CriYTKGxV+A4gBrIppC9gKoaHmApbmz/jJlbqQcElURG+x6ce+aVzzlKpIXl54
XkInvrkdW0kVjD1t+OxRsbyEhQVUEMQmM5fjR5Wucqt+GAf+F86+/9iYUpKXkPBW
InAeDigeWVRn5yxB3DhWr+IIVKIIFEcP8XITraozoqjJX64PmT06wCqFoVx/p1A/
ND+J1wYEKGmSR0ZEsqzyV5foMUrCqB1ZdbgZMLmQg5rMCX6m7VAVNJAXy6AmUxJg
tP4g1pZt9fmFTlXYZkeI/6cnu2ovhFmwdcZJE3BLoTnIcyTemtqm96if+aFd+zKI
OY7LXVfo/m3zpyHrcD/oUVF7Ervp2xYnMbVXck1SYOi5e0/66j4pM0nKEDKUCIyc
u9k+HfjEv8iVS+7bE4RrRSxp70codvNwc3kaM9oYrYjzE1yBsGCm7KdYh1f0e+C6
YUsZxQqHEp9tjdZke1qwwwamZzYJueeTwi6b4iL6mewE82QZWlrCwTETT1InVCPe
BYkqvyxAghlraAszT+/av+da/psTPwONGQUh06LFE6cOpJXRLTWZUqACx6Gio7Im
laOopOaVhOFskB98OcbuOTVodG5SSyq7jWhVJiLGzvPszgT6QH4NTB5A2JmrNl5f
1UtpCn0AzoF5GtX+rtldWLrU5IqlultTQ6okjlyyWfo87r0V/b2CY3pRZY934/xF
nZO7KZjNcbtAOZTRfzy6afNkwlwidkUCjJnsM+i0H9cwKIF86UON/ANvZum2R+sk
D9iwqzBCxPQpdc1rkPVndpB809OfevtfVEnKM2J2ubuEkpLTPNqdIo4JzWFNH6Hq
3Y62E9sDHjaUjRDjd4LqbxcZ8kkxKHdGQqplsUtZXH0QSUaYYNJkacrDFFj7vUn1
2Olgrjdv3TVRS2ojsVKbOkzBLr6J64Tumi/HmIdlrRskucnAcqoul3M7jsJ4S19i
9m//k62iv9BgE3hvHPf/fKwojHY7d2fnBgWe0vuC+OB8IhdEYpDz9xWelcJb3JPq
03m7fcxQAGPL6OI79eIPW0WLKBcSzJ6K+zk+/7Yw3cP0QAyJzS9XUPW8cX1JsMti
Ng0Pv6knrSfQV5B4NhTRDpu2SRWuiK8PC77Gi9m4zbgeL4aOSG0kLKb8Cce8GJCh
PFc+Uzhl1uZ83TIFMddQq/N7cDd++LkYPwtIZGhZc9SOZW9wjHoVX29OnmAuOHwv
SXPgdccwa7NED90F0D5Oeg9cmBRMDVvBCfAIVE/0pdCTDg4f5hthunRY0vTG68jh
Ca0wB2bi/XaSun/z0F29lqgWfoMJNFqc+d9NwDyt163Y0CRtGBbFTt2Lp5R/yZX/
+I3cz7EfVBqeUgXhX+hY48nveRA0wBXv62MCGApdahMRIZltd5rBBzZDDKxbbjK3
Upf4FxB8IYxqaNOO8KEdWUE5R9QWYTCFtEqYDdXZ929/rEQ2DVeNyxqZXChwgiqB
BGrOSyDoCS/tF8ruzIch9QufnhjSQYG6GOrt7DPSONC2b9vJPLVkMbzwFwFE9fJO
2gL9q9tu3FfubLb3sz2CbQRCnMHXzbUfkAHLsgyKSP/884x78r+Q9SMGLBMaoefe
4QhOfZoi9vGZDT5lgDimv2Icchps7IwpxFay5t9CcXZs77xHY0cpg20o9opiWKah
r8SPQu4y966iEHUCWhMRvHFbUv2kq4LMWYuJP5FjgjQxk5xAy9M+j/I6tWcdV4o0
esxNF8P0xbWpnZrYJfAEfrKqSKtBSTBWjSs3WwHcAyFQWJydeT/ruaw5LPF++rhX
yRJ9iIJBCPxI/VE9q26SN0Ijqvg3TW9t5lNS8+3DjrNaovSt6GgiTlUhrkSeGwu7
P1sh7CnvzESiIop/gTj6xz+3kwINul8MlghHM59o5nYXRgtJKW33lm4pgHFWRHzV
3Pg3EMR3a6bHGGN+I4e3bZUCCNCtOJaZJIy8i4x7PSoNhymwbaeDkV6IwRQITdxe
+4qCN+HPAam+0G0TxR+q4Zq5Z6VVMOUd0TBm3kP3wpRnf/sh87SvJLJIBR+aVYc0
3vh5Yi+0nbZOPEfvwRu29rMdpE210YJztoE7veBrzCYBlNL7n71wowNVUFwjtdoE
27EZYTy/pRRY428d2qvIWiAvCgaW8NKTkIFUyePIW9zoLajAO3vd8AkU3yQfDIPX
Fvb8eHbplPhcdtztQrjU1/kGn4xJpOul533SZcS8F1kyOYmqKLn26/PPSHG3waRl
iaT7HhQOWeh23sU5i1ToCPaQmQZTD6IDfkWU2IWDspZUAywRgASg3cEWSvW5Xg7J
dQ+TwrU2SUP7xAWl4d+GzKqinhsE10ITXkh1vY1VeZGfa+Su394yGJmSSLdMXkpd
jpkypiNYXJ1IsEEA1NJAdv9AQIHiRNpCrEI3Mk0S7kjWnQGJNXc5n188NYBg3VM4
WGK7U4Uqi83SSENbn0e6Z3vTkFHwWcxMyKSE0NDgVSa06WcDxrXR6Ai+QX/dJIw7
nenOSR5pfoIsXy7Xofg4qL9sqkMb/kxqWZZrqEhOvup+CIurmlFpmyb0RdScWQKO
4rQqjqNe9gJkkzeRBTkCQQmkGQ3xJalsmxppFeZ7FK/VH0f+P6GWX3Mca+jVQzKB
XI5EFnVr8nSKMlA+XFMW7mQ4IDksQG5br2wsYOtroMN4mLs+iE+3xgXePN2bQVz1
B3Rjf3coUyYKVbuDsAddkUwm39WMORc0dSU74LLBFnnLF3ENilJ1kvGfc/gtDTY/
Re4BtoaJQ5o25tFKDuC1XoMy7CwTzsVSuGlKj4z2EL6CNvD7ndbsQQfNhJQieQ/x
66oKxusF5nAAOYWHX80cIcysIwg5SN8iZt0wAkeKy5Ea8kJyOGKTJM31M0ConPpS
Jlw3es31FnYA03C5gSyU4d4eFVPUp1UDOTLM3RVE1eNigv0+a7sAsetyj4p/k9d4
M5MtIbNG5Kw0XLcGq5OwUfLvdg0xf+4+reR0qot53G20K+ylILtEYOQk9snSt4Yg
umEdWGXzHjOpk+dww35p8msTD7tH48FUWGg6KhTBDHHyCOd5rullrFfiN2ljFFJE
LXg26MTIWzb8m8cBsUEM1qW5DiJX/jR3x+jsbG2nmocb4GnS2m22sH/xIU3MsPJZ
i9PHRHBEQXQIt0QdK9NMAcpzEGxXp0u9yEZj+fau4kYuU/15EDZzvHKSYWis29jV
y0vlRV6pxaLpCPd5rZT+itx9wcAueiw7QUJLGclp9r24HXgtFcuuyZnGBHUaohn4
3BiE2JN0So9pS0V0OMyMmjupiTCLd6bWgpcJfEsq7W8ksyQTeb36JFRYXpZILovz
ZJzOyeUpG+oq6iE8uTxbNoIN2F6tJjx6mG82dH+wpDHakx81l75Sh/9PwgBk2FhP
35QegA2iB+loJomyc96IvwJ9s/g/F+5+Y2+xYkS1z2qbjG0UKffaZWZTDc3SZh5i
y3d5XadDA2Bu2AT391V6pf4htM/8UOBQAqf2Qo/YJcVTUrnnEHz+02qr5qKli1c2
7b6fX1O+Tu2T+4H+oSP9eL94ZcnxXvJa+U6ZZ92yKWwhXNu8rviiGhPhs+J/WkgB
G4kGK46gCTm25eFlPVpnoD0Ch3fVYsl5XWUdYfaC9HZzwpQBTBnrEjziNpqFpq32
FGtmjHlyZV/Kk9cmOyw94q6uZ3OHO+JaBgQlKNFMXcgsXnJUZIPvD2Yo9Iv2oN/z
/DUBWkGuLN9QE3sNb6t+qiNyyu1tJ2gbBTJHKb1eLHaGXiRXeGS7jn+YAJPXLKd/
jCYI4PFBIavIks0jVej18OSpCispnSv37U12aScCXKTx2HDTgqIpzNnNyPbAZ8mA
h0OZ1EfkxXw28jrOL2XzNzzwHt30kSx93VodHPMYQ8408eItjQMUHtBsI6ogp0Xr
akHYDJQs+EED7+Y0Ymjqi4t/hlF7+EnxcN8CnMPhmt2oPLqqZHBCARqshoM3x5C2
kugbdSQ1yLnN6Zdh15jDv3afYiRENxHavmIzda4kTP/weKfXrbkld/Hm83aquLUq
Gnmxwpw1ws97hBD5I5+h+W9r1WgnVPvUmYPXXD2zH46HmGd418ocQMaciVjTp1Qq
tDI3OJNbQ5pXRrx5pynamtw/WgqmzHe9QIV0LCvb3M13LsqpcKC7ejtEyK5ckyGZ
YJ/wM50vYa4GUY7ZRxeHscE125zZgtYvKNecIlCHvEsuBBhGvkIR0zC+o0fTkdMC
GjCi3iXv6oXmYHp/IIQZNns92KECHru4qN6JB4sUVotpI8tVONSUj8jGB0NPM/9X
PyF/vrGT5udKkCMx5D8FWQekqDPpoBhJok+7laLNLzhpZzrQxjngZfXJemuPS5jt
s+lbY6PdAXawIUaGstM0Ld3u0n6iE9K0Sg9Iwd5tdWrWXkXw+7BrtdSIldNJijBB
TIzGtz4Jw1hpBozeBzObmPT6uz6m0+LMjYi7xWzEJex+Kf4uJYVW+7B/bwZlGeKY
qLcA6LBfPeZSmNe62kMaDwAYjdkc8WEhPrs0r/bE6n8kFVObYA3mEst+5s+Gevj6
e6+UOv7jq0/s5TScCaV40Vl0Beek9uZgL7yaBNG4BhkP9dsdYq04/BiABaBuDOTb
YZ6w5kEL4HiLEYfeLp2+Xme9/+/jzQJAsIM4bJckMGuauT2bjZTLzIUEqh3Dc2Yb
pPQoc81Ersz9o7G7bUPfQgu3gmAHtUb22F7m/oP+sk4GbMreM1lCRHkcrjWHKbmy
GxYCv2AEV8+2STD++yIswHAC6u+DzudUPuQpSLwandzHyk0QjouJGLVCAP46l80N
l8MSKfrg5SMbItxIboiAbZ6/pa9xGKq/PxFvAV8bY8rRUmYthyXHTh4awOzw1fnk
NEZzoGM09DtX3JAFrNlWtetSfTLKon0SiyBkU+rnzdmGInua9E5nXnWz1xyuJTsd
JojuC139cONt6kyQLyEXRvVDembAL7qDPB7XLgluZSlm8jgpRNw0QSOy8VV6b7qV
DLKh9sALC7Rc0EV4/VOyY8xJu+z1B1NBvZHG4MQ8Z8Nxii3mL/LdUG5u7k5/OpxG
MxABJcpLhtAmK0K9oWZML6WInfBiBLU08ktPBDBTk4V3aTr+0Gj9Jp9zotWhua9D
xcSfbbUThfcxsH44QQ7CpKpTPQsYy7cQSV4kHIPjwG3FZkWwB62JhHteqQdXZudX
R5au4FarSTax07t0uJQGHeyqDUUaRj9fZNhbcHUZUY3wQoHza1MlSzvZAUNGj1qT
LLvw2s0NOd4oa698agiSw73Yam4SJWXPnKp72r8615FLH3Qy2R9G7D7psyu+tAGA
cvFiMPMRe3VOmDLNl3D9/i4OdrBSDWQacixlFR4pYBkuDioj3rSJznTFaDtFxTJw
ADGnAHsfDXMKwtgqL/GR6zSxUz+1Jsp5ibk4Vp+O+724Df4EvPRy4lFhv5eOADHI
D3rnXWuNXj2iQq9zmC52zOdIygmq3cOD+riCAurX3pIAZs+L3t8BQGPX+2pf+ZaE
L/RZEVWMVRSl7Qw5WTlpnX4F32XMN5DQkZelO+ZAAZ7SRSXcHfGnwF/Ydj5+tMFx
PAgAfPM7twHaaCL7Zz821ZUIk6X+hIBdg4Q5wDgNhir+O+lr7NjjwUDGvi1ibbgW
Hek3mTt6WBpnl7FPhGQQ0wp36Mxz8rKUIEH+uspNdb6e5X0zaeepXQ/s3jaFSG4c
buOk0WrBOTD71nkpqT5IqNWoXTj0C64Gztbs5NwPsJ11SWFqjVyv19NoZUJUXLxR
rMyxqE7s5hSxGYYPX8PmdQfGa7cmt9eTBdDisuaUzzR4WEx5LbTD+yBupOnvCc1E
nxDwlP5LZMcGnskmW5Z0VRtYu+dw2v8LYpI34OA77gZtH5qGSIArpaqrs0UZ9TDo
0j7Ab61VhdaCMrkTalvyG7QVAFQ5+AYet0jZBBM9uqe5c3FwUPKfLs4kmHAZtfHq
7SVoigl3ApJW5pgPpopg+D/K8prq/sPKUGVcvTq+5G78bGt9CY/0mN5EjO/kEF9O
/lha6Lrac03nq1C+YlL582cCOtZnElu1YM6Sn51iYG32dWMUcy/oo1mP41Hg7YVQ
+rcCHW2HMgyNwweolpjE9U5+UvR3FpfoORFwIZ51dbl1Gs8C92xh49hQG9+RSObO
a7SQKBZGjoVazaYpdoSRW55uJYc1dImNQmjsMcNO6aTF31SGvlEppM/Hif+QVKn/
7vdZXCCCOGilw+tjTid+6zxf10bRmD7EpeDDbLiNq5WCm7WQhcBVGCOOYTRuGLI7
4X+3YcUbcLv+GoEMSOSHbn1fN3qPiaTTs3t45/4kOzHi1WRv5Y96AvXZiTj8rVfF
iWIV5kIUIdzBLW22GK87F7ktqpC1PyAFfYPEGM6JUNjQpjSwYal0P4GCojgRHa57
deAn88Yw7GkAPwPqQbWAK85O3Ye3GY52tgud7RXsIZFiR8Xm+JL7jQDRNd71iqmO
e7DnwgC1EVbnWECX2GcWAAtqM8HwNaLuPzYyGGimCoQfg/odWZVtO/MnLYwq/43h
cTpJb7woGDkeBvr4mk5LFa8m2YtM+CGYY4yRuYpsfsZdk/fz8NoMnO8gwV7dsEIU
1owgNAV/yd+py0A60cVZjXXApsxnLCvbFVPq2WL22P60/iP7ANt0e2OzcmtV4Q75
FZmMFpPtOM9pHYhkC2/BrXWwOngDlfFCXUZTZLZQ+wLwgBli2gZ4mqNJc6ciCZuk
p/ZYlruHAxZsXa0TQ1t8VyEllw+B259YW4URhpAzVN8hT/nCLdYn4tresjWgOEa1
onF0O7YzIliLcHBRCOvecWliCBBn7kG8ZGOTDpGfUVDjCW9gE9pu+yVSUTlvgnP5
9NQkpdNi2TTKbFVLykDmdocGkZMk4f9LuHq/Cq7j9sSqbuUGerKt77bcYU5msc5l
vAt0CALtCigrymkiV1B7vAMVuBzaJ79Xg3pc9CMrp323ZQGkP7AQxxZkD/P/JhZw
mTQb/YnzOj/CzU2+ipJj4HM/s1bufpUX+JPqq90m5EyIdcxSaerrwldibhkv50cO
ZJexXaLotf4Xg877RlCCdPkko5FSsZgkAKlfxxyeDEUyVGaj10ED25fUjPs8qC/+
nWNb/UoX4lwW2cbPf+2rLGY5HljED6xvi4+NWkfl6YBw0x2nUTjocsYfrjz6RJLt
1eP0pjZGFzK35RZOmHQ/F3wX4F89RBEywfub/oTcO6IWQIiGGJMQdM3iJqvh2Ty8
l7oo8C5UvpfNSt4aRv78zpsbyzhBtjW+ECSwt1Ajofet4hdbnmo/3pIVlWl8I+bI
//UtohLJeOYB0191yeZHlQh5sWDfTKBDScHkR4RXT0M0VN+hClufQQKuZkoAS4bh
743VVhpje6y2IVmglXDyqZmzbFlj40TGJIOAZv7UDCsrizmgQmqMOJyAsH+hK9Ks
iRDqQH/2Lj4073I/tFyPLkSCJ/TbHfKSORgjrLrwxD+rr3Wx2w2rE/P+J9o/oTIl
4RKgD7tElW8gmiuXa7pf+OGxtDJeQ8kw3+cahRrK6+YOhAPVdVCEXn3CZGOu5coW
ecvdPN7hCPOp7M5ANX1bHV0Ag1Zx2FegEVhMtn/lA0CXHabQ2+7/+gnJO1dgsMTy
7WBBWB2AI4uYgUWy+5o/zPA5Qe8DlXLdvcZP3ry+2PjYD8/95aKp5EdmGDMfxQya
gAG+o5m6IYHuZ+7znTNmX3IEFesKQfzLI9MX2/wbpDjm8AobngiS6ckJn8w2Jel0
yvgzbTszY4MhOXIzInmbwtzmZ2fds5pJ+97YoqMUg1nefPH8PGUNiS5ZueDqZVis
ZWe4zOwvg2fQaZMF6MXCFOtoFoCfs6GnXzjT0dIVEveudhlS5FjlUu/DdFFfltKr
dap92GIlR7W6WzyTJ0+9aKx5P0wCOTlfSreEH4OvJ5Bhnoz1iiZkKcyfOrN4thZq
TSQaudkrCZsOtkYXsko+hz8q4Zu7JXd7bHP8Pd3SDyBDORSFl8hOeu4r4HgEW3Q+
wez2rL12epfTSlnwdoqLIrBparZgR7AQ+vLzwR0xjRjTFwvHrieG4P9OK+NN3dKp
msXN3av28ooeEuTsa7FXOcXrt6qxGsUvt9LhnkHBcD/CseQqZv1KEdOmEfCxazQe
q3vW37Yy+DIyxhIcIh4vGnL991kVJkV1lVAWQXiKq8lObFxWU9TOv912E0qEG2Vt
jKfh8ELime8uEonkLpHujshwN2JBsg7JyuTF3iXuHOBmSKAw5I9kvnR8ltHOzGQl
TDoL2uz9HSlbDT7yt7cXg9gBmPcXe61TWmtNxOPgPdvIzZC140UtZjx7MvJsV8v3
abWdY+TetZ36lIKglyFBNwGJ/EB4A8zQqRe4mnNQzsmKI2fwDQE70syH8LPG45QE
gWlDehD1nPO4SMjVXf5JGdq+VQLz3hvFyHCFUqxdM96dxCC/JvOHoO4Vo7akLiAM
oI4/IdTV85WZsiKOm6RKTJz8l1BNk6DKYK8c8veBHMIWPfVYPIAiF2vMfNzFF13u
T2OizW25EWnsvbLtXNTBrUJt5zNHxJc5qRTAWV536DDQFMHTC2pOZxqCT1uDNPek
mx9SySOSUTOFJz3rHYIk6oppGgH0BXfCHfWq1sTBjoWrqB9jNgXAixINPE4ow4wL
w3Cu2zwcIQI5kXcnSsL2X1dcrN3MCp5fr3xsRKXL++ZhApjD35uiUb5YS56X5MKH
+Yb4hs+DaPp8rCxYZBXagXe/iXln7c2os8dTUx/MQeVGu1GiwL8ErxLWFAvvkiGY
9fo/FLaX8NVT4jJEwmPME7wgZgqXlrmRnoE5snr0skM7DCXw2RxUbK3XQnBUTQR5
uCCC26wKfYet851N3uarMlR9l5NUfyFWrWKIdB/mergt7aV5Tlf277VgZtgcZ+O4
thOat2wfjbA1fNb1jj7Dpb4I2mwOxEfsycXYG9pfcTdLwQAUv9RFPquHpmPOxdvi
wTegnDVRfVcZ8DnQh7ehv6fZPovqgcaPCOw7i+UWQSbGhjFmyUku8NOHKedBe1n7
Ue60C3BOXZdptvfm/TthVl1+1OIeXma28kD7ce4hBbKAgUZtaWLwS8nVKr0P4VMz
sf3U8INEg7FZ+tkLzLRC3fcx9fSk0MXQB9C4OPRq4/tPeYs69f4Gs1RlG1BtK/gP
8UsmGKCXKem3iN3reh2eFNggrSU6snBXmq+jz49OTWGaWCnbrVAt2i9oIHLGo8Y6
dBUmcgVq1MfOAQ5iV33/fLkPsBD7rfJp/koyoMZIH5t5bmgXcZZ4+xl8mKaKAQCM
Zdt8rcTtATKYEEmEwO7LY8UTuUpzjYIeKn7K8zgheXUrEL0y54SM6GFN1D6u/U/U
sn/DS0c362iil1/72NVQ1taF2JOSbOrr1qm3USFPIGwjarDjIvCaOpuSbu4gaYsf
M5tXprz+p/0P8LDtviWrVoVDXIF2D38OMHrwuF3DgiXnyviZKkv6SyExhyKbkikI
GzOh+5qhzL/EMFXitpmSf4vqnJ8kLykxZOsUSECcf3y/V5nceZOnvQTFDzwdWxnc
FXvrx9SJl+DmvarKr4RDrzaGHFoB9XeoM26v1L4NXN8TQf5hHohSwiUKNdat5QHz
34gEJLz1S9YE1MbALZgqOoekDnwTnNXeta7CFy3Aq8m45HO1MVT8QiJtZ2/s0xtr
C6qmAnk/k7EZW44qgltlV47MXAi0iwv1KFuwshO0t4iFySgWL+QixS9EFkUww14k
i6yuKdp5xdamdH4VUf3l0/oEaWLH88M8EXY3cN29nyslTefEzN6fAY/pOoKKT6hE
LSPD/OulPlblYrlZyYjuI5qJRnAIxWbfsPSe0kTZmyRW5jiArb3NrsaUqDyrsuQk
mHJhcxjsqf/UO4ANtEsmnVerWcNqUzK492ANya2Ey+Y3i0jSrwty8oGFhtYzJ7Mo
5LUEwZXMi2iWCzKPrtL4TbSDd1o1XRhhe91CQfz+4yPaCc1cxunCxz9PpZ6R9U4z
nMtQWAkqKRmF74yGR3u2lPR0C0wdhsIIK3kK0gOQPl1fu85mX101CeAIEg3MxgRw
5KHPMv3WYhgFCfU2lkTbY9z4yvbtVnVLVzDMHacIpS2ZGOVNfDSPJPZZK0urKZpU
VoneU6fzAKUZXnv83P5lRayJrW528FGX8v4iIP3TpLrqvYwBauf3p8vchNokgMsQ
MnJMfaTVZalsAZrfW2dE5Frix4+VxONBynb70X/CgHYSs7y8D4r6fWrj4DM/EJzL
rTi8OfDjCtSRljO5IAOcr4caIDiLEiUqUY1eRMHXyeYxn4JxRep3XV14ViUKz0Mp
c5n6zO/y7igrK1ImXKm4p+V7aNj+IeOwX/0dllUvqlpPeAmHz17E2jH2II5K+Eku
onqXWF5YZ20uVzPBNwYw1rSF90383EnDGuWxRNtdpaqZQMuwUjQPWTHeWHmsKcJa
o+e0msbg65vEBLoiX+eusm7KAHpbgZYoSdVc0HSDP5htxtbtVFONEDnFxIfnCaKv
SAgVjT3Xx40KA9+Jf9uaw7Bm9VDcd2Oh1wdouY1vn6NV4ILtMMgT2G2AXa+bI7yD
R3ZsnDHNIiIu5Tnl+hKre7BUJdvho895Z+MNmKtyKn1EPvmb4i2bvlCC4ticVRf4
EaJ+p2D0gpcf+DVKftvBIOmx+Uwkm/Djht+8jafBr7V99y6VmfqVxIooVWcUTUKq
3zeX6kb8QBtfuWryyDYbob0qDV43cSRMu5MlBr0Owh+Qe+iB13ri2tZVv0iRf1p6
wVskkzJ3j7N4BpgFZR66O0ZkBQQO7zNuyHXZP/XsOm53QP8L0NWP2/wBcwt80vDT
sm+HKqnx5+pbrEOj08470lxZqKsoo5YG7HMLxCsDjCPbLYpMg3dnZXbwPHec7AuI
G1WfSzvhL2+dPO0L7L7GUQ7FT+Mz70evsrOvWWRqT/spjRu4abmdlLnjS6pLtfiB
eWpb85C2UuasMv1wEMvdcPzAxXLqTLcjwPWaghSSEtZ39edO5LFlE5oDxAX4/O+7
yrlvX7h2TpuGidjIufUxIqafwx2w4LIr25i8Q8nGYiV+/WLTUgmlj6otjbsy1/J4
ZA19uwKTi+UkpWm9oQdl61ql0dHWKSWguMI3pu3N2jrf3vxFGwmrlQOM/grfKGQC
pU0pfKBGlKRulyA3ulBlJ5sTCf/tM+i5IPl0aAWRo/XrON6XyP0D5Lyex3VTCs3U
PFE+FkXJoEu0uUoulAN3+L595on38mEJZoL7ZMytJJkRy3YKT6USx1k7HIoYLqb1
u5LRkdYwdQYMowo+vXiohHilT5yYAQPwsJq5hBPlvappNpKk59pEAgcOY9meWxMI
QIZ+NpWLd4eGSHK2LO2xvt5zeeet455eX995Hy99x6u0UOuI7WCtAefaRqnuHoxR
Xm4YmK/cWWOxlvoKN6p0SHSZ+am+DsE4Sc5IuE55g4odzv5uL4NPp8fh/jEkMpFd
kNt/hP5Zdp/P8BeH7kb3ubdkjglCr2EoY71HgMZtLfv46ByWbTtPB7/RNbWfgC5y
swTuSUWv4GHIJ7vrNnAHabJQ+y0CrqOUuaP3nygvher1M1Hx9Rh9T0LmB54o6f9P
Vt9AKLg7bkUOnS5w6hstzCe/NPOTJlTbN/hKaPlSxNimPksn06zxwD7n+WwpZo5e
CAuPTWP88k5L9E8p+LO5Gz/aRHMbZy5ENv2vcEZwD8y9T8p8vB8a9zM+Q1b2o43u
e03ROJg9lnuWB3fi/D1UVCdZ5biDxx7q0n2Y5PxM99mRlighMxiIKdK1kTcQjEQr
fMztSVoW1l8NhFejTawJmkpLynFmBxXftxeUMueWUecsYAoU0hL7xNUpFpAT8AeV
Jcfbn7afw9RqA2+3v3IJeWUZZoGgipRBJSkpMj3y7b9u2TvrPA4M0hlkLWF5J1mx
a+5y3FF+l6nMEFw0W7KrDhuOQ0JbOo8xY1HafPB8YPfEaTb5ynUmT3vqzUlsDIQX
jC3hIUAF0jrEAHO+RZQE4gF6grwhSjZjQJd9sXdgCp0D09FfnGc+wG3TYK0UdRtI
XUkGQAGkVaLYFhLZ/VJ9F4iEx1G68mDwQxRiP1v/yBad/6jKYxHekoWWtHfo51qh
gNWiGDefr+nJpEUBtFRRv9gNzghl8ylGZY/AHT+jeK5TDL0hCV9ICsUtQHnocHMt
ZN2HgE8jbZydC8dClZqP4X/KxfC5zYbRbP436EohXGrD/P1BtXDACeTPlHSCMp9y
rGvK8F4Ya586aADatXkayJgBNsO5R+CAWkS0yvRUTD5HFeE5eHEv5vnLP5H1JwVM
DArSIr+tyBKBIEaM7UX87lIPxSS34F9MynIvZbiLGF7q9qhhrHxzxHfM7Z832ewa
Pq6uk65pp2P9uqOcdPXo4VKvHuqpIUwjD2Df8PVssS9JyDm+2wlkl8rNHIisCSQM
TPmJ1KuzFjDtrZw99kHIySdDHleFX9hXJSla7Woa5S8gCm5ZFMAQt0l2ovI0ok6x
FyOiwy3OF+y3XO/5c3AKva1brUoYN8AzJCZNtySQUpU8aNdw5GCoBA3Ljc6Aq4hy
5ZuJ8aDDnnf/3ctetiJNjUV718M6+8SjOjLogTyuVvBZK9/70eqn08Wsfusi//fW
TDAAGSbNv1dXmL+iAs9H2wOmkfd3gFPtqE3+5wZWpBJ6fCmnNO8wF3GyJidbzh4d
9SEgCKi8rbK90BXXqFUFVWmjlAJ8/0IpfZn5KNvFc8i/f5ozKf9qA6RfJ5YCiHTZ
Lq50FGakswzEoO+rrXSpQW9GbRka42rMnkHNcYjg3Lo5aRhoIPX76FMwxb7moEaN
RFBz22tzENDANZmgzgWiC4HhTFYXTIhPen9JfEgpvUfTOU4li9WHZmD1hCkjlAZz
3tllXjV5CAPi3bD8td+GmGz8ab5hY2by5Pxz4oF6FhFVS0hiuYF0KRJVLVdDzX9O
VlSnV7BQ83cLsN0SRpaBaLgJRfok0CW4rNvh3ZwyDKxTWNCv+zlefTEILiSvuc4f
klDLop8hqvBhMAYBmcvn4cTc6sIjZxUK9W+BcWa9DCTU/qObb310IeGefoDPnQNj
Qr0jcHXKY61KaVS1x6ad6HenRHZC+o8EMxM5NFiXp2igPITGq7pfW9OzqHfRqAzz
QTjtTF8gtC+NnpLX227TKLk3BWhxP4cunqxMxKArWqC4WuHffA97X0W7AOhBONcq
jUxbKjn9TGKtICJz8nVyNsqdBE9WJF0xz7I8K03Wu+M5NPq/g+s5q9oQKl80vsiv
RDe8uWv2qE57XHDuHf5sZEEkfrewKMZwXC0fBy5f+xIawzVfoQH+ricHTLDxA5m0
UMbOmYkZybV20aWtOC0I1kJrDH7HDoydd/w3fhA8YkFW2+N4Q2UY4AMTd/iyebIS
B/4mYfNaJ/f9MYO/caJAcbx6HpWWNVV919ArRZoVIp/h22yfWHUbOIrBzmh9/b4x
w5tlrVBGHFZiEaZgR2Up1K3kra5SEePI67iuB4iJLK860e9yL5gqdgxpe3p3zxNj
M9G8lT/WyBsEgW6uBhABrLbTcfTGke56hSnuolhuS+MafQ3F7PFNcNM1yANY3Q5b
es4Ll2G3aKRk4oQZ7t/ahSVftcQGMDXFn68IU6kvD0taxtM3hvY4Pb87/p529KwG
qsynExqmGlic0KpaofD0/Os6BwVWIGGWsSRKRjXAGwvk743+kDn6KxNYGlUxv8FN
npg5ZDqaTUy985EZClzGuj/Cx2rkTKA/Bkcol57f605UcnTWiF1Dp3FLDdZvQKwm
9D38bsiAlSW16vgrqIszx+mLEYUZmlQvxhsaR+1qxRX1hYzHkvv8a1MPCcMhnp3/
pVUxkkmiC35+baN8ToBcyh0Zsd2QstYpzGN1IrOb04fuT0wSIWRlfqFtgDywJhNI
Qlgu+GloagbxZlY/W97b9OyVAThihBJ55AS+NyDfHaHwArtTaSmMXxngABruupzQ
0xyuiyaqL6Y6w5sR+Gk4tuWRysqiCMNTKpqCbsmqoko8ftNt+0f1XSlCMDxYX7Rn
vD3/hrvdT1EXyJ5Oh5RXr6oYuD2tp+s41TwwVI+ZwK+/okghQ6KQzsIjjX5Fa82+
vG6tK0ecfJLt8YZeckdAXjpwZ8+v7T4tkGc2c4OWHWFuJsQgygfllFENs7f0uXuB
mRpSnZJoqvTd66AWNW6BAP1d1DjjLsOxZgBYWUn6zlX3iizv8TTJqLlRPseovoxR
l0ACxXlkerS1npYDCTPVyA8OcYeQR8zNC4mZAmRWEgQuyyxpg57ihisHLkcD0Id1
zAorf8QjvATnR3JQK2uxbMbahNMckyRdYgWmesMUCZobVTWmLkLUNIdtla7Pb3im
OMJZgKz7Eob0jmkm8yQhG9/ZYpX7T+CIZTF9sNVNH4mb4tdI3QeqMG7yfzr+3Z0f
5nNxK2OR9a1l9DRMlOc4WEs5eLMqvULqS/XIgVWDCInbO/VmOkrcxPHyAPa5rT/j
SHBTG+Thr8ImEPgKS9EgkVv9QTKKQgnNjq6qL4Qe00S7/swaqpibQdC9VMx7HhEa
q6GwKKRRPuZ8htgkgBVy/Jcr+vD7wdz15Mv+f8lnsnXFz741c8Ymwany1f5xY/Js
psBnedszhpwxRgqJarizKkBwwjT0/p44QZ1t0KwI9iQvghT/jVK95uYJb5Q5mzZm
e9uFyyOFLngvO+7IZosWrE+jAd7nHe9a9Hfx+yJN/PmU5RCJ95Wm4Jt8NTG6lt6t
DuY2M50GK1VP5Sb4uAdXa9QkEt7P0UclwaZPN77LF7SV/4KEVFOeXsc2bMfyJsnq
7CO+U9t6lUDPr+AoxHyBtW6pB/3ZRVHvifzg4lgYTUGEFANhvQYztHIH6lGDcyz8
LtYiJPNeoYs/fYvr4IzvaQqvuH/4NkORPBZkvBr1Z/bEugzVNiJ1Kfrb24EeMIrz
K1dZSULpoZoDF2dLzu3g3ZqGCEL7KZP/GAwbXRpLTfpoHuiJOtHqE/Scj/bHA5j3
7WWG8F7NsssLDqwJJHcMGDKS/+iX7Or6HDAcsCmi3a0JGRBQdGSP5XnKEvBIKS4v
IUR1KeAXtDThppJqYCsx6rOxnJbIjCGgSm6aioiKFSo8NrN2extUkEH8dgJvtIQe
oFVccWApbIIqTwAjDEc82T1k4RFvlwPWt/YRwjV0LhLlHgKf9+6R/ewLan7aaVY/
yshq7/OdzHMF4vud9o3LJbc1MCsWHSrh8OoPb02Vw8vxhT4Lrobt2pezjaPAQrpG
3pom1b4QVVrEzKDbp4ryO87+Q8n6ZTB8jLn8EQwvpPSE2vzLLJI8AT2GWcZQfkYB
aFyY1iNwSi7SWGc+GCHtFofuLfdAUjgYOUlAOTKYzILi6Gx0qwj4HNgY+hCZ69rH
F2Q/wl74t6fs3I2GPbNHSJ/WPGmr4IuVkUk59tfyfBxQxTyWySdYtoMIdVrDt9ho
LNPlaHDHZBmVuYtC2OAWN5JQeqTI/tO7f3Rv7T1MYREkJFtv/HK8d8waL7rtRWw8
UY5wiIacgSIJCj7XqoBowIXS3okZkpx9Sfonm+6OQfSIyCuq6mLWinTSTQfSH/AH
fTcfZ+khdbAr+9RqYGO1q1Hj4i4K0Uy2PcHmV9l2JQGJj30xyyhH7WmN/ozUQ9LQ
Qpv+YoHkN28KpJtliWkbpB3WxeXmx4ciJmROwEXMQtiXzM2Q8OFdjQVGTvCy/MZt
BIu42GV7QZu9aCa8iS1AgQ0ZDgDk+DHUNdyUlhl5tufYOOT5arRAVf0if2p4NIQV
V4i4unt66/Z6nibsCBAIaLAcGfvTcrhSzzzFgP/bhG7i0NGtq5S+C4snBQjjjCrT
B1EItVt1FGSuzTmq5IKMnAXtlAjNAIm3W7GOm4tZgw9v+TkEpojRs95FneVLHLNR
0Ar2a+gBFhS4HFi+JkJUVaa9D1Nn9wIg8IqCz9uJawkoA6wwz4AQnhG2UGitCHt/
+dH0M5bh0GuQai54N41cwmI7yMYOz9e9UlRndDUkPZS0LcukynXeVnp3GY6+XvdH
OvNDljFFEK8P0LXJQIEiIZ8DLtg2p5U1HPPsSmsMH7pslXhlwYxb9X6ct5PTTwai
+RECQemUiDbqrokLcFMyOBZ60K3clxCRooIotFloGNnTzs2h6iKZ3nnMShBftA64
yNuw0blZLIyuBdETgmFpb4w1hnuXjsAveO1ByRpLYtMtvIogqommWrG+7Zp2Pyzl
EHSuI9trJN0QSgFPm55+8eFEhWGWQGPUYWRcfwWWVkW0vAan1RJ0VysyZVPtPUHZ
KFo/DoJ6LH3gf0RSgdWlt4mWRGDjyO7bm4GFVXjWSy9BYmOZ3LS6nBQQ76qDe94G
8whToEqnmZC7MCuLTm6QhWHY3tQK/YqK3yM7buGlughe//1N8HrAV5o2bzZ8jEe/
YQ+acA4/FM49hOzr0EdWMM+1EicaYfRMrtkkJjxc8SjIKWBZwZEUDn4oLSdmfS0K
5T6oozsbjuGuri4Ms18HQtzsCm86wekKyNVO1tXAujxls+Y3TK0RayxyyvSbgjlG
3vIW7BYO8plDUqnbjhCDGNvpsrdV8vaVDzo4lf7zHYZlnlZj1//B0db/dJWyuF+b
2Wiz7BC8kD0RyHiWQIQwlq7a47cEisjrGZTizlZFF6RqbL2gyk1xZ5/steI2IikZ
vNksXqo12nypH5Pw7/aNUUs3NKT1ih7xLjVLpWwSG0jHwKmp51+ASBfMcEbN63nB
zNgz6xsxQUwur+971sPYa6EKgiX03De9yrtGq12ojSMOUaQotcHaUSFosaP8BSjf
zA6Y4w7nzZ8QGMfetl8kxNF1OmLkO8hBvR5eWUox/caXOy9I6gQ6pp6roc9yNQUX
u09m+Rd8LfaF4ux9aSarrkKsXLFlkS3wLyEZi0k6Ibp5vPnFiPtgWs6UbhTa2+DJ
mTXYSUCgwEnRItGgrnSAQ5fXX2V5V32Gv3EgDj0klmokMr0J5RdVlO7KUxm+LYZ3
h6XLC7A/9qikFxK72W7pwVno0iM8GN4yNETkwmOjL/pbBB3sZHVUmeVgRCmBHbUp
eMl2VY4J4Rnm7Yfc3WG5FxcKhsvVAVaDfeWnZcpFWwGU33ne5Yxifm/z1XD0CBqU
cyDMulpvAVA2+yhsVJHStGzNrYNDGmtPQlMItz6uf+t+5pbYN6Xpf3UwBvVW93YH
30Cv/MK0FNdqcrfBQ0532HI8VH0Wv4y9dcvYr00jr+qhIhqhxSzpETPv5SxXF1cz
sl4SE3puzBVbRX+xtF+gFwLSqtgnOyJW+HpLFHWLmS94bPnKs+vY8sG4FgUzYgiw
wvuLIxFvwuX/MHBy6H5BD5LH48w+jVH4pM2lKvYcTAVGcR4ksvJmF8C0SQmFXGyC
cDgNZMDF5iTyQuY8rJCTdmhhqnEjzKjDECl6xXHAzzwhJjRXfot1uTXfVmzKDfk7
B57uQwRQreYJRgPOift6SQobml0J8F2WWmq93BNYEOnrXjuownZGtFBlDFCmU/gw
03BxweThDCah+aWcZvAVyOdVv8Y2gz1amAXbLIMEafGamssnKx2jG7cmAqX5BAX3
URlsn/H08KDAtRtEOC+LkeYoojvDMDqeu1dFQoEFkeguFc8P2TRN+RFejvaB9rTb
de3mhEUHIJ7UeCHT1hQzsNG14kzXCxOHtls2kxY89goMVftC8cp89o0zfIyoViSK
cPYOJSkFb70HhepJzHxcPCx1sbK4T8+fiWoGcg0m9n6AOfIp/Hf7ot5x4fF3TiFT
VLOSv3WcY4oqa87y8STkFEa9nt+zTj4xwzJ9W2ywL0xL3OdMRUPhDFIvwp6YHT9C
8ORNJi5F55NcsaAxXk0uwwl3MOgf73W+H7xBpV6fsTcaYZxl081Y7ph10w7NNn9o
ic/Lhx+/pbcbIF4WFrC7HFQgqxfS6oXvcdHCODk1fUNPjNcVBDfoVw8Wt4ltS8oa
GIqt9h7ngtR9RYmRMNHzXOHuZz+5HbG4Zmf+IhUEFI/ghTnxmucipwczZFfc2xDG
jFjm+72UCw+YyTqBT5xWFcRJAGJgZ9NLd3iVvx9bwPPubExF9TDALDjJ8BB65yCF
UTM52M01o1KhUfNj6ps/ehEDXsb8tnclAY926MXQrJAXpvomwGDuptaproljEVFD
xzH2UAFQP6IlGyJlAg4HvyX17CTXTU5+HFbgD5G5MmictLebkLFsJyIod38m5uxu
2DLXydshJcP0LhkRwx0afAHHAf84cxzmVqLkmFSc6WbksIiE5U1JGWq6kmEhzZqD
59FHqjPH7BGqJn7bhN/njZOv9LIK4LK2Ow/5SwhGi3R4Ff54er3cIhruBCivYjD1
OdGzD7Xy3vhp6PpN9AX5VDby7ZCjvbe28bTyx/ih59pdOSTv3hSOuZ33uquJUHxM
8RWRjjvhhj3KfdT8UNgEkqHXp1jgIxLuvHqzFeALuwwqp0qgx96cNxqetRn5rSw1
udf1NNhWJaAsMDrJtCm8Lua8RYKESN6zClgQmesNPemZKYVmfH1jLxdPlSEqY1KL
M8XkI8uo6qBFgUaVWVjFTYwhyMnFH3SowUZ86CAVdYlUpNPDfCKwPgyngGPLREoY
N+AUZUGAL4DLXF6RvrIPXINNMeVbM6B5PZR7mJ1lFLGZel5yUAaVMdHYxk1BNLSX
bLcviFs0fsVm9bSOu5Njh/2pbXKghSX/YFdjmLc96Gfw6Z863J4H+5+qpLzO+5Kb
BCZoTSg0DCWGg1Zuk/3qWtCO3W442XxRbRfSq7NoX5M/iZeOuC+N0ImMo1DDvrch
6mDJPUAUst8jA7KeTg+pkQQBrYqDlexP0Xt+CeiFpeFMaTM3TJErGxzWduz+qjhr
daRDMywEAEPjpmefw+EtMSMrIwQKsakZ1qHAhWjU17rC/FTPh/SSKaLOdTEZ0UCR
5PnWLaThYpHQQAJQqEDg95Hp1Js4V4vbSy3GOKqTwPeGSdb47TIF3FQazI3Jp9tq
9+zELp09yBfQSFdOoEUBlUO5OgtRxvmGr7CERyddEI+f0i5OovK4epp2U2SU0FXd
1ylVNDReNx+Rxx5ZEuqZ1o18dNbD4uqBhKhIPlz27JD4ZGP1uU6a3RtruUYsgPr9
nx43IbuGXghjoI+K5nQwCvDPyQ9Of3LICC9Mcbxpd6nn/84r1BZtr7FvQNlkwSJT
XAce4d9j+/C3oNSAa7k2+6bOQrsDsmhASU9CLyAEKCjtTYpGvaqCuXhuWiHmMYI0
k7112r5DLPmIoizHism/sJwJ6hAR82XPOyeDOHPBkIh+GRJyRnm4cRatAD7IBIXB
6d0z6Vc/QSGbIFIYpeqmpY7eE37VBm4leky4bZgQENeETY2wt+LM2+/ciS1MwrI2
QfMvcDBpcZtrMWdTXtZ3ynm5C4DQW1RiG3eZ+2/q03wAQcc70dlJADOh3sgZdm/y
ZOxCK2VicNLiIbJZuEZSqGaDvaC7172kjxcUseCFJyF5ljwO9Jeb6NRr0bnHeIKK
Bse2bohtNThF+7fZDVFf28WdTmJ5GprgdOHestYCHZY7pe+gNhJQmVrQIFlbdGFz
reRSZBA9xmcr57wNerWC/zDbcsFup7fwIikG46o3EEJpIquKTijMFhd6cI0ejL5l
QFhLqc2R1yUrKY1RwneQgMrohBJv/N0idQ6JtPE4f9Bq5YCyVKsPmN1H3/tX4cQ5
/QGjOhgC1SLfogWv2fg2fiK0pnlHBkwvgTVmb30DPVIEBTitv4Qs/OTQEVF+Rfjs
u9u0SGURvXfRVjaWJ7Xqm572buQJe97dJ7b5Yz8myfn++xVzw0HniHsrSW3C5u4E
BVw38sdt+SzPNNZvjRnunJPMJJRVTOPQ4snLb7zCMPdbs4UYtMFW78qpHwWN2uPs
lvU9rnZtGP9FYElzvDNhxYNxlE3LDEf0/g29PCB7qSko/ZMBKkiJroJpyMFaU6Zp
0UoGlm8T4rt8Xiq48X4dT5bglyrGyAGd5Vbzlx+PIYRR4bRJ2ViNYYao5AJDPD1M
xTsNegfYj+Imfa+v+AEsBJYOn5o49Zkn3JhLhYI7JMvOLCqzxhQniWoVS8bJt2m3
zj2iE+ybH+ckgRehct+3bSSr+XoPmICmdgiOmT4Bgk6ZbyhmEGwv8ut9uP9BP6GN
j2y54/kVplEyvKRWMrS3FiMnPjGUy1/t2h4+qQRhYsXbw0afjqOt/8Qthz0ItQt3
NJPSNFraiCrDDiTq0nl4nnU20Y90/S8gqnBtScwaj9AaxstvO1XESECSRjGEzOIe
X7NOAqa6LtMIfZsKqX0ld0G7Y/y2XU8TpRq4SUOGKyptYWbU/bPD10lHf7ZA7kvi
JI6J/XhaXsIq619Dw1j01Jx0Oxj7JirdrwK41QQbbWUmeAlqybm+CFtGH8Vjw5Ze
bqeqZdbdzc1/F2kubjjHJvp1UwCaPQiCB+cTEYiTDb4tHX5Ar51THdJuvboSVfzq
VSVEm9jzUFrT15elYl6WsQ5A96lgo5GxV7dXOhzGMrY0RvggIxTg9j9gd420F6a+
Mvum/ZTrRowo7MuIxdl9fYUn0Ks/77Yf7aVen6+5RhEuFsQ6Zh4vsPvyrLX6BlHu
a4oIPw9/7+zyXzk45uNLoJ1P18deZtzaC+CV50BX6ZUMleM4DLH1MK9sgwJFNJeG
BQJ8y6wKTbmpXIqVdHvzljhAxw6QS54mqDSxK+bFOaN9afhwjAS0PQQ0V21k3OGA
SumWPyjqIHm4FvwS4eaHRs7if0GZdWQakD2gRlvz2pYRLhyyP86BiMxSx5nfpMp8
7bYXC84CNDMhEufyWspz1j5ZKAxgBfSMXX0DczzLnHAsE6h/2jOBQhvxua6Xqrv6
7I4w4S+7E8VuDotCX0/UcLiS8Ng9nmJJ9dm2TSPPDE8z5h+FboRyum+pgSTVKdc0
aucBpZHAVwolKm3ck39sYdLVkBXr7MRBnWV6kSmVhMb3UdYuOMWfpdDGfFKeBwqB
lsICOhAGw2qhc4IBMm5dzjtZLPRmtxvuxJVM3G10hzRF1nCKWPHQpWczBfCaXFbo
nzmVRduhp167QnzV6XWQvQjwfunvEe/+WY/HspUEA5W9aSxFz/HIH0SkRlOhsg0b
7xoqMybN1D3NbQcLui8EHb7wdCreSrNHHzuJyW14etfrvWIhXPP6ZWElhxIchudO
CaYVeEmSqOUUlb0CM9TY+SExwOhJEq2pHd4k0GHNAwDcUUNU06MR0STWAwOPNc31
euFWN58dfTgHL1CiR2fdgBYYmcU4+zMUI+vs7hI7PHYn2oZbU+CYEFF1NzWEhh33
aZ/GySmnap27HvYry8RE/UCMLFIP5XIGupDHevRi2MOO7AZcBlpU4GAGWUtJKxhL
Wzatryfc/Q0klNiqAb7Gt1jU0tb8vz2lQwLk18BH38IYw+wMZTjz8INpq/brnslZ
puy7M15OypeSnVvkaegdLevuLUB6Iw7xm1eQgxYdyZcKL0Aw4jkiocbxcP7cchNv
1bmZjSMTle/sKe724RtZUgsfCn5fkPaQyH001iZmx4Mp1jR1VQOd4QHGHZO3EHX4
xXOevur7MYEW8C0auKzRAZPpB1nLGO1SN9H58ztU8kwNyRdufQ7LryKuRkiPqqfV
yyPqOo1kKI8arAXpNXrZzUh36UGOOKWUQLXB2cH98w/S+Js2NBDVVr1yndTA+IFK
N6BNJQ/R7IaNkzxFUg8BuKSm3OCc8Z9U3Ix/KY21D9fazpMZjJWaRKjk7EUrQelC
aCh8tVd/gpA9f2k9V4Fnx2E1HUyOPvGjzxkfa5Sx0zilRhnvm0l3KbJhfczx+daJ
C9UgwgDurn9B6iVdrWDCKbh8dcJmUGI+WlOxhntPSxA8+Fe2fQ3t9fLDVhJt/awU
isvpmZovZO0AAE2jQmL+84YZ8W0oyC2HTr1SFpb/QcGZ1L4qfw2baQpp78WGCNDf
ugkfNgvzQj5xp6iZRB7UjdpP3TaM9PgJQ62yoDjNwWZgQCCX+yj2+PB7dnFZp2Rh
OBJ1DsZ4i436aGmDyGemuFiYzkpxoCEdFfSaRVKjwbOQQZMdyHFAbo8NTdLDbpzn
R7thR/AGVS4DGjv2zWQLFNzq0GrwxMkL44Qdtvo+9LKzIBmckgwmT+eCMdDpSTl9
cSLvwSn/OGPwrcG1A8yDk8MVXYh15ltLn5Pd5xPpskH/Tk52/5fHzsO21/03gopi
PncyEjx7AO2B0ivdDO5fDyDynS9d0O2I8TMoN5iQUniOsj59GaaNbkiRAnDrACME
mB/Hi9wRrd4f80BMpk+R7xwww987bqqg7PbLFuiBYZxVzRapq1Z/e9JtPteUtA48
cjLV7oZFaA73GQOvLruQlR23cpEq87a9YcckM1ylA+PSvqG6W7G4XHk7oaTmLkFW
JFUFeY6On4kI3rcxeQ/D/4UHPr9VFQbB+mDGCpkMXXT3DwmQMfMujOAmmE3wFiOk
GmVh4iVLI2ISlRxm91B8TjMoK/0rC3TM+oras2m9YI0UjNl43AfUKLmBSGxfSqXM
NSZey0TPNlpVv/qAlbc9pSTrDTCrhWTy28/AwtiQStnONn8u45P7PxHJamrwZEiy
9tT7rCQ0koFpzRRCSqlLoY36Jxl7Pk2VKID74YiGf8gsOUspfdgJ5HJZZdXYPeRW
Ox6IuBJ48RrEotb+VVKWSnujc1r2K8eGZl7jFuaVKsR99JBtVPYqiImiSDVjOno7
N3PbUgMXdQtwXQGlQNeVhWqgS5LtqpEkf4oIbC0PWTU49hdhj376qR/TQcVZV/FZ
NC3OpxcdPoXOxb7hqb67exm0RWhYENAcJ/KyrOZvztu8SI9lOntMcVsnOx91fyNi
VifcSWzAFPOO0v3Z2qSzhRv3bkINl9vo2XLbWcF/ShllX48L7+P+aE7cP5adJTF4
O1op/YnzXBi6ioixzjqAO8OWXylHGp5nODGL8a9p9F0pLxvwNYeEVXhu3Cw8LXV9
aEPKnRN8FGwm7IpUY9To5cw/Dw9UfBcrXnqGrkfxDuez4LA6x6UXtHyjS+p20OVA
RT0nUZFRK+IuEkhpKvs9kZ8s2rjUMpyz7Rr9JvBw1DzIJY8mG9KCSczGiG7+WCCv
+Z+enyah5yghs/vcTJFrBFamuk7B2yR00331v8ZsXWPOxHR0LE01/NS4jbOOLeVB
gAz4V0SYdYWSEKKA7x0tVC7aBUMKij0828fQV/LDdtVT1ETnzGzW3TAIfQEAE7f3
D1wEB9v7y9b5ANjLVrrzhRu33dW9gdXihH2syJwMo0HhZv8/k6+rjPf1HLdpUf9J
p+qo1Vdloc9UDfSUeNJKgDoVgNmLfP2l3OqLdazj+qZCzCyH7zEJbxWpWCefuRyS
7Jy9WTEY8E7MqPw8LxpQzva4SL+KIzEs6N7dM+hSJdROlHXJtrXvHNHWJ7uwVRiy
s44U0iIJNw5Io0ZwhLpfgqB0MgwGwhpGp1owj+zElyLdYNvqPTylP7uX0iMlGSag
PtgDcbsIDSMZXJ2aRyNBSEuZepfFDBVxFyGSuINCd9uh+dW9El0bYnkXzX8oWSw6
2G8qR9ogV2o9tCsjOz+LrzbhrgLCNF+/LIK+2XCrK4ZBPw2So0wHocnNM8wyfEka
zDYaVt9FvBqiGFpP0l6VGeufYiP8Qd13lTwjmZVzA9vVSR91H0aHgvt2iuXum5Zk
m/puzkk5aAfCU386ugPwdNMYBfsTu40B1oQVMk+WpkaRLO4QCwr0MLvLwWu0+naU
ZttNjiSAF/RBRWqcfYyOnzH6QxnNnLgKxgdhTfWQpN+55r94MBGF7xEYsfbilyVf
hSdodXLOO2ko8ptPv9rRzCaNqPiLwSXNtYsK50umCzEyxDICMxnHLoaed1BwLgu4
j7OqCgwQORKKPvOy23yBoVbJfNsY8Pg9jEiwcAP4vo1Nd1nq0FbRydiB2A9QA9d3
2dKMG/GZ8YxsvrZpMdTn+eWjNJ0lja9GrSaz8KTuZ+2Kzi171XYHw5hEbdrh0xst
xM0+ce+9fc9u0gtBPfa2gBMI+e89oSPRugizSjtM96I/YTleOmVwp8jM/gcFanrJ
hLEBVC/Z+rM4A0K9ia+9vY3BEMRDroLU+q/fllJmkLtQ+ICIaKENbfRd6aUeTjkC
sHFzYnw3TcaYEmWAjLEmWcfFlcSqXAI/t7dhgYWw4Mt9PZJR6u/v4lmpdEEsGREH
UQ6NTQihGSwOlnRHl9vPzuSqOPrKlZuaJ7rznkgzi0Y/vs1wtXAntuE+Uk88OZp+
PuMglypjq0SWRHWeXD676DAWZekzUNdn/F08NSU1c5dfXvQJmltbFG4eRFy3YL/b
bYlMf2apJDT48urTe7QrfilzNvfTJJjPevnd1m2/ZUf3uxPfAdylyF+DcjEG8UdW
BBiNb7HxGbE4rIZt4zYeP0A26F0ZqFzwkmzvvXqDWPis7tfLi2KxsG1xbFdmayNW
sI3rlwFKutKpk1G3CUwuXCuN9vlC8sPRrYKXxXyVflZXlR7gT/LmP6QTV6skhVQs
JOtz3X1X5YDdNZBNnVnRzd5OvWs7bd3wN3cz16OCL6bvk/FjV3ngPlpwiiDnr1rG
gdroS9lOZGlRxKCIOXO8a8xfBOC/yDSOqWXgerGZQtfFN+BF9Tipdk6EbcHpI3Ww
Sz/janGyLX30U1+Hzw1niWoghFTtem8IXuNK4j949JG9DMugdtZ4OOIvLx+Njpg3
SDpWFADVTvsygEvwvH9/bD5/efcKyCkJX121QmuDeq8OihHL5FJYcsBGPJ6QwnYe
+Mebq6KYHKhfKqGZfv2o5SyYwP2npP44LnFVnbaOamK2cySHCOjNBiJhDP7xBLkf
/aHwmdGFS5mPTlC7YZssKq+Wji/yomxoN/Eqk73twic+MEq3twr1kTSbfxUyfFs0
7gGCPJFmhrl+KKopRWNLo1C5ihkd9d6KAJD54ds/LU6ebjQ+8+e/PaWH6fej5Yf7
tbX/Mf3XU39e+cyvaVrfC4ChbzC0bCNN1W799zAjsDJpfjTqZxzoYWh0ZPPPlU+O
a+pJzUygtx7bJ5TvoSD5OYyEMZp+A2Ep7rNRPexqAoAX3dvuFoKSM0aampzX4LRQ
4pfP6HN3P0Cz4ZBj1/Px05P9mZv0KyyI/LhcexsMhN5N7PYe6IEmwvSFf7B+WGDX
o5u/6Inn0ZjRwBxLYcmRm3nrs34cZPFwLsDHCac991advQGtL/n3vaw1vM6tDM8h
ST85Cz3HHrjetYkZElueOjX4PLq+MH9RyZH+3A02ANzzbd6TAmu5tDhlfL6XGIcQ
vB+FY03LPT/ZOOmaWUCWpA39tpgsesMVbshhbLVvOJYl3SRcsW6ynRoSd9KDYCMB
BM56ARxGl9xIRfDuKdN3MpMi9yhutgDcxXVJMzdM9uUA8Fhj4iW+0/0P34JvEAB4
siKJaRZ7MWLn2meWmPCcKTLustOD+YjiWkHio2UF2fM2IUQXOVITsAmyUFPrwwrh
zN5F/vftlyo1ux5vKAX1Dg/KsrYq3pCaVXzKJLLfQlp5MjxxL9jmNT6PGacUe6CJ
arprSJhwo5O+JHFuSwkbneQGTAI0U0sAKMFaqc6ckrLWe4YbSqr3SYy6eiDzrNxQ
wB0lPEMG8E8HorOHM4kd9BXwW+KL9z9FnG1DGjXNcIdVLMkEbyhJ7jPSSnggLCdN
ITBU+6NiccDTk8JFZQP+UVF1S5HRmwKdbZHx7/umENOXm/xlS6sWvV9HZdbAegyh
mATS3/cZTwdpdfsy3uQfytw8H1cxZBSK8zvvawBNdTJFRYMsobIrnbR1DtWDDbQf
xlqgaC9k73KnZLLs5p8zKLUcnzQFR494omkOojJ4MZmPgyjvNIX1wIAPOrNJLgI2
U8I0PKYQRQ7dI7sLpisoZI8K36XjnL6/FIf4cA6TtfLmCDAhXpdvfL3kxrt0dTQ4
N0/aT3LcDbPdLmt5GiHcM6Hu2UdK6hMl6WfElK1SHLsiMY67/Rrb8vl5JqlFUJTT
SNEMJjd966oCnX7UR6WoUk8JSE5gat3UyqpkB8UDJAfz+4KW66e6ZZTie0jF6dty
SypKMoCbX1hG2CziYnYfoap/4Iry6vexCnZHmZkjCXXOdKdmWV+b1qVsQDCR2gpk
jMaHTpWgSNKi2GbkBU0fF34U7bCLTupCO6JpqX2tZeFCqnS7Xb3W1hTMQZ9R6t4O
SS37tOzCu3gWtpX+JCyrkh40cLT5InN4myS2A1K9yDXQV8jgN1AlXuLgSCnT80/1
ps2u2FZLsBZrOTufiXLyNbkPvrs+hAtwX25OJDKn5CYnQu/XWScFn85KcervFNAE
u4kFv1Y5PlP9SeHqMldUYfv7J8RKtG+7a8Q/otLW/mrqmO6LCl/kgbTEz4/ilWiV
++3Yu/Gfx2yilYHCOyEuWKzBxripmCF74dnTct8pOgzCvK2RyWlKxPxW/JOg6zqz
K7O5oW6yPDZ+S/PlSPhWJy1fERo8XPkieBYkqxYBDhVK04kew4ON7uguGThyimbC
qziOonp67Cw+fuADres7Xtr0Wvf76MLWmW6poRnc3xUhlStp481f1COxYvlov5kT
F6naXSUcCs+lol4aR8iMsF0JO3vTJbGKY73ENPHcQ6ZfKJddJUo9zy7RwcQI23Zc
24q22ESgqDfelujGS47VMAjj1YYjJ0LsykHhLcQi916Q2ItX0SpspcCdKx9nAZR1
FVP1T7Y/tjOF6ARU6mfqStmxh5ltzNzxnmpEnxbRzraepgC1G/IwSF7lgPcTcMYT
56cLfLHlJ4QZXgb73gjNzQQSgUeevdZ3Hgw58QL7L9xgjT8GY3ZnReJ12n3OWzQI
tYjSUYEr80YmQGJZOyRyhdes6IihtrX3Aezyv68W1GC7hMqL0QQ2W2eDsc3RxLlr
qE/CskNq8ekDgFrI95cAHSC7Z4QNK+sL1FsW6IOv2oyQ/PlvgV8/45Ozt3tZjaUJ
BKhvXrJjG3IAnkDFnsxCK2bP2FLukVUE5ManYc6zE02OsWuXOFvxMrDkQOucssxP
HhpEgbYvHMhyVsHmq0yLyoCOQUVoM3ZLzrKNgb1azd08gzlQ1gD7Etnsn0UKpCrE
2064QXcmZI3udHNleIHtDgNzmlXIhDPv48ju7I/gGv6NCMZLAVsLBZC1NSwt6YTM
L4Aplqmw8MizgcKel3U6WcMrUtb/lDc/N7MahBOG+ipL83ZQkkS1Rvn3IlhB4pWG
oMludcOqoB0F3cDFzbPxBAuFgDXEHKmkQnDUDd5ZyknFJ8BBsriZh5/qZC+0zYSg
TbvkjudYS4oOEBgdE5m8E9+YmsFRuG9lZLNop5Yu5+Lm9BgPNyuFZqi7yoPmtSfO
5Ju0lK3eNbvLeaRyCRKdUndSheEIv+GMgBOn//iTuh7xevXW+g55RGN60E1qnIGF
OyhNyEECMu3aorl5OcMyKjQOat1zRPZA4qz8jmLpDfNnMv2w0aYEqBW3ofdgXSsn
VBEr3BlGolOCn+L6eyGyOJgwkqWnsSrXUeEJZfPDNhb40UOeN63dHrJ2JR4LJwls
Wn89dQNP92iBwgiBhaSdgm5Ms/Lhj/KAePh/aFmhAUXZ/k2d0hzVQn3c/h4uexCp
5j1sAwzHsJpnW0z81QwW+yK3cLsneReqiJJ1e8i6bFHHUKBizPwOz7AgaBKY3Lew
de38VzAk780Qr244ve2RUztMy9oFhG/hMBO5SondV90NKraHIvIK7KUkwuy4Qy8P
P/ga5X+QYgXh3eQJpT3ZrvwUN8mUTRIT972sN9LMTEO5omtUunM0m2+Fj8CBY1e7
yspORiARUkUUZ0VXxso+jXrOkjhQq4w51dJqTiy8jLnOXpdsDAwv4MfGPuPeBfFj
n9YAPFWujST32bUS/RIlYV3htnbDn8vv56PXEb4xEUNLul0+gnvKEf9SicRqohC2
8UWCR03FDb8z/fkP47owyTJZUKkdfCzgty84FE8Sed+Hq5meWmkq855206KLboiR
MleQSQxIcoO4YjopoHIkaBQaHyclfY34QcfSxyf21JsE77dq3GAhmtGVMjoTi54y
ACUbqXewZIV3dF23qjucw8y2cJ0OcWo0a5qjq7r/TVcNOcXez/rZl0FAohzBxexQ
Gqwdrtz2eq4XDuI0Yf9uLvT55wwxdoJDVpQsNXUrmGfP+BJDiajig9PNUO+ZRqfE
pkj96RWkhUT1UJ6tec01+wrbzzCYDPm6qB00VXF3qJm5R0VtZewp/AKE1Kr2znPg
Iu1Eo8i1FP5j+ok8Zefj0xfcc4fc89djfY8PtIkqtrd4SicAndiaPp0aGkO6sk4i
7uNnx+wc2KWweb4I3aOjLdZBJwcIZZdLuyBEm0fjuIhkN/VJR5PPPfBTWvls33YP
kWyqEKk/AMMXCeRC8nGTmAPLaOKysw2mPlo7Boo3y+UVW/oppTLXeCJ8802jLT3e
D3/0TklCohqdOjpGiYLbAWd5zQZmW/0+t7J4kXTFv3hdxO8LvxsCR2JBD9mDMP2b
dzRHU21txNGMwnqZV3FS9zRBaFdl7HZjgG6QXZI+Q2sWR9CLyjCeq1nf44/k0sHc
8wInVyAOuHO67fNkg0aV2+qP4Vq1ZCt4uYQzt/a58+WD9YeWPbMIzLhxq1g52L+1
z1Vt1VtD294YO1HjalLQ3qXgQkPeB2UskyAZKo3fAeUnGPvqEtW3T9RAiv94LWht
RiqqRmDWupQXTnxa4DSfEbPN/9sV7UholLY8g7Rj9+hTTk33m5XlOBsWJbo18Qsr
V69mmq1azBzJ3H91vwr7A8RiOng57/ONNyLctmYNIqWq1hwbYEwEhRyidG9qklIl
SOr0xCepj77A5/gvyTdWiEKWQh+FWXqg4tgVDhtfbeebM4n9Asol0ngKX6rBzSro
k4wSCZniJ+F1tCcxvgu8UrrBCTI8LDTR3AUZYyuyScMGxXqM8fjBvEAxBX12mOP4
4rOr3qdUGzK9MlyY4k+3R6AbAnMB9kTht7hr51fP9u7m3zMn4GH6zuKA6jzveI2G
obhTID0hCm6l9HGazCuoz1F4iColYSCbPKESGAzmlDG1s6Wu61VmryBCCYKRzayP
zKPL2sqCcMuYTQnuiYdzj2dA0sFq325dMRmUBoHnY9yD+xSJ2RKfaqlXghX1yhyH
eosKU2F1lljWcj363nw54q/Ql3aGO9SDfQvGafATGGzPh5Mns+TPO9q1XSfScoqp
YMWrdIIOEm+x8DifHaeEu2wFaM+i/2H3doTXr23Z/rxC8qFIxnhvFqmT6ftLdt7F
v1TuDhiR5lWVl2s5CxiS8Y/+aK+QChe07+QCiY0saXd9pTWuUpG2yw4Nuxa32QjL
RfuiodIKpyqsIxf2Wredkzzl4Q7eo8Q3WkXG07VUU9hL9a2FUQmxw+ZZgW9ntGPg
tuEbkL+BEhX+FpjENNx8tTDfAxYk9MoA9+esPzKR5ATagZLCRIDJvDo1rrfpz/s8
S7PVWIbrXVddPCOZrS51nOiTA9l304AygYBNcSuoL3x4A29tVDlyWNK6iSvrZ9UP
tCK0HhjNhZwu5VPCV7McdngipDE1dkM4eAaTAFTuoaatLK03P1jNeYSF7gNtCXZz
iNHxIuhMDgJ9Ln5OHAiL2ZiehyWL1/zpoDrQWLEXu+T7RpM/Czrde7HA7qTBDDl2
TTvohEm1FrOYgQgYxT7zdnb2MB6yXF4gZGdG/Fao1/sknbj6bju3aDT4VbEibVed
MnPDLy/rhc+WmcIA3K//XKi7ygesDhk81XvXEsFFP+/d8RdHvewbYOkUIM567bbD
+XG1bFqVkYGh/109KDUY62D7BFfRdXAa6Ayk9fPat/xl6Cek9sytee9VTHhNM1MN
T9d5w//0pt4iPGUbp//nAp0KH0DGjHe1BZhlSyGxxCoz80iu04FNdjVEdcOSBv87
byTxPWY1WCzHDvXP6WMf1lwKgh259s71Lu1zVT81uMvn3g9pJtk2YGqnAZmepl6/
TXsCvJTEjxXyqEQmDX8Df3fSsgKvld37Tg8Kx4K7JQiHboHU9FxT6kOaCQuesiDT
F0SvysPEM+da9TThLOXkAsoD/uCby4Dy0oQPn+JljnrelzVNPljzupC4j34YrrJJ
6PTs4817kE1gGebF+hTOnN36Pi64ckhzlpZeQCK+oGNe4H01j15fb+HirvserXSH
gFsf3qIsgZlc47Hx6b9crwOPmmMwRGFqllKQ165x+Z+i/AdYs0FmJf/am8qsAoBt
EtCIZmIis4CfcPyPbkUMsyE4pbvYmbG1I7stI2QbIArm+d8+0xHPMrr34JpEhaL6
wLDWLPTL7gUehNo+fbV+WsMsJL3wbDQsI7nqa49Uc79tweRJK5jsifG1+Ir3IVH6
nnoEpBER/3A3NkDgDspCnXktcWAixGI9TsakkuHQhOBXEQdhpZKkoPr08KfLH7Rg
HssdueNtZiOfSb2IXXcSKdo0UUSopuRmHIe+2dso6CUH77rCY5HqHxtT07Ttrlx2
XIm7RDnkriCOMNYUrQ8V2RnNlGvkez0GbLI42D8ijAUwK51i1IabLNDAPc8eeM1X
Tq5vK1USLhvvCoi5i7KxUnkgwYG1qWCPPo5bG1bixjx5+2o9LinkM/LwPm6ghN4D
epq+iVpORoLLrhwbe8GS9NyW7CsY7sQgP0T7PmPpMtMBdoxx6LUVjJrS/wog0TpQ
1LBse+sgcIliuHMjtKDA7TmmcOwIiOsXaBd99RVVGxQUqyxE//p5WXQGGiL2ctat
Ev2EK7no0MUUpO6tYqsoCrM4sNyaqAelv0kq0KwerDdCkr4HGzStDt8PmeAq2FoU
oe/Mm112MJJZnXgI/8DS0tq3E7X9X/0A9B1XLMYY7jz99x727BX9bb/OchIAM0UB
K+DSh5tIfv/cqe2fYrFrjiaH4FAC5YvZ+VDNTFcJwETwGK1/H28JaFttUjv/nVmA
ebycPfmV1hwSNtbgaoWKy+ARGRdYA61VRu6X8YGVVbabF1ZebYghmopHwCpwbGda
1MDfN1iPGmR5WmCBW14zGbdLSsPYxzPlVjuidM1kKQdPdO7r5kkkYT+MnhUNkd+j
tcz+zjXwGODlJdDIw5KIfTmKufhpHSiQpLU9/gf/nZ1WohDHnUFwVZA9iBllf1em
naNDgoo+Py9CSa8rdR12o7bkpNpJl/I4vfSkWqXicu/cg7ESkKOvHZ2K3NlDhkd7
/VDMiyQr9yFDiueSXBw2oDVfETiw3Ak/3mw0pU7B2VQiFgbe3xH4/sehAfhwrQDt
RlAZsyHqr2f1nS8uLvjsfXuldJFGcT47+T3Dj0LoDds3bEhWCEGAUS7AhsYNKrU9
xG7An/e5UHARnvfknYe+77/J6gRgwfSNhw5mOrQNYOQOE8lwJP6N7mGgjpMXeA/7
3Q/btRvrKr1NjXDC/cqoeGauF4azoY/phfRfJkNKOOgII62lQHBFkEC8LEjfMHVA
IEdaWJ3mQutgOaDnLXfIXoVCji1BOPh7Pj1vOpGAG0GLlZsWThg4hTWY6sbjlMQB
UZepNiRpy3RR668ZxFbISLyNsHq3qAmWSJwUOTqUzdUu5iyjRcYXKiGtV5miO0bD
mJ/nQqndJ9TyrI/lm1e0VyW5OUEfKHrsx6QWq4qlt6vHyllXAEN5jqvEaCrtPieo
+tF2yttscfXw0nRxuOMLECZ/qI+woFV5AW/7ipKM++VMbYqDdWewJuy1QUdYC7FO
cIwzi69wae/HspTgWPpo6AgHfWDIZ/LLTcgYueAhW+9MWQl5ze8jIyfybbs+H5p1
WWw9wuAkIykUKBRwV46bkx3BhJw1QZB3IzsL29JwAFRbcusiCG5hzwg49zpOEIoJ
RzMKO0j+YX00fBxqppLLyyGbf06i+b0ZjAQ1whkLGKp++fmy/BCZGpT36aJPLIR2
6tDiSJWpKhcR2U9DUV2155l4CJ0FxXDEAj3Ni1suswXo2XZDV5W8fXg56nxEVRT3
Qu2tuVmGtfgh5rTDwk7q0naRKyxT99nEOViESQX+dD3KWE9TVvHF/LIRi/lmh1Xl
kQXuPOGZm6xd6Xn8jTnWUAQRSkSOGUsYEzdR4Q0HQydOYV36jVGw09kN1LGaF2ce
1bKlsblWooBhaSM8ITfqDrwKhVAs0Yl1D937fFO/3J95iejFNXRhKu7THoDLJ1FQ
NZeh/ixKuSsmVoj839pOn3vnmSNWWZ/X4bJdd8HoOS84Y4HOGnAfeud3SjyBt3kO
AfZvpGJRKisMTR6YaBWf7tYH4CSXEQvRiGhWSAl9zU8eai2l7ML6hWXHQxM14h9V
cTH8TGVc2qk/FU8BaZsjdQPt6btMpB+ylCjnGv0rcax3doh4pMPql0NDpZf4PfU9
a8fHlCxUxQaydzkTIPUHRa/XjDpH8uP1Ul5KuHP6uU1lAn/XIcP3q9t5yHH0niZe
3xA68jrjqZOm6GCywgUl89Y/jmuku17TQPV3GMDXOUKn4CpURKjden/O1gXBOmp1
YY2/Z9Esw3yxMJV4gUatey+Icr16i08Zcpu1R8nEMotL3DGeDAO4Wgjgv36jCWEq
qBta0wbMJgijF2vargD0ePET/5qATR8UQNs3msg+kA3qLB/I7SsUwtofcQMr5vk1
Hz3wdkpFZeVXracoXpQjXhEjpJ6uz3/22GoFIBITn+9W7Q61a2Z6sM5Ybqubg5ZC
vPYCABxStMdb69ujrEOJnvUZ8OQrgqKTvYjm4PLaQzNcoyZMREMDbta2TvVUAUC8
z74MPoSuCnS7OofYNh99cwnjHyFiGV9VH7ph+wFkd4llsWEsm0cxW9d2ApPrrR+H
arkdEmUwIYcgzfIxUYO2ZDrEFaMoQNWZJf/gr0oTEZ0f26WxiCSPr5RHLPGTNBtq
H1Y5slp6SG1WrJeA+0iikHDMD1FeteeT0sV7ASKNGfhAKQUfudyURtcdvP0b87Gs
qghjcSqBFjrm619SeGans0FjRvaQbl383Y2KtABwoSBcc+Lqw3WI7g8YJEC9KEQP
WVRJim9P7xHgJcFwOkURdaEWLb55K5I9VDBO2WSYxPHiNDjjTUFZ49C3HNTl6e7V
kwTzct+IqiBfFN833i1Pgv68scftHMCD0kqlJ4jdpjFaYzyGeZHrtCd9uyeibkn6
zAAuPLtSVBvK+EC13CTfsrRylqdEuVbn0SdidvZ3OH9QgojG8QRhaBf5oxeK/ej/
BgYqHrkLZBh4I5ATgbJxMRraa6xiqVu34utQk61+tXb9UhzV1oJku1bxo9iC40fa
kNnRD1/2yQq+GE9v4OY5SSbt4uIp8wpDD6ReEZ/Zn5q7Dz8McG09Va2imKWfbg+H
7jomXyx2MzADh8pCOC6sL1iDFyS6vHdZFNUEO8IZ52tAtmcho+lYrMtp5aXnqEI2
Y/hKgS0QTJwp/LiducFzcv/95TL0ixmw1blPY/5n5NLU3hiMMTxq+oGoCuGbhJjx
lw7FEN2hhmIr0Uy1leAKrqCvJc1GkXC5zKfaVw7jyfT53r9WipAC9NAN3Sf0mANN
PQfZ/nXzBDRUgb74r2nv3ydwdbka/Kyi5vOkqX15HQ96VY8f3XA/7keFDLPORV4S
vD4/oyM/uzRwIyuvcs6D91oEF05SwIdDYM9lQb4X3GKKonNVMXAN8W8rQqhfywN9
oNxPYYs7E+Sp51LtRPY2/b22UD32GVlod4OggBWn894cwm737XRDqaM72yUKY5/m
6zi6c6ZkipJ/9XmKI0Ar9ml422+knahlYWhWkQi+aIJbbU3dLekvvWpvYCGtl69h
0+X+v2hx6DFGgK52Pll71jqfR8kB/wDCoT4YSqOVxpP75IG1DI1inaUu/4hatDly
+YKQ8b4x6WGcOJPbkUWiUsFVZnCz2t9S+SanrrHoJCr7BOAlAWDIxSx7hslvoYuc
+naICPWJYBI+WJf0D4AWNDrCISbsXc/Eym6JSw4xGxCVh1YWX42cFFGvL/piNtFz
J4Yfkx0YcS2VUEBxVVEGr+4dP/cquxO3cSbTGQcoy0RgKH/zXHmWGH4k+wbrLgNg
ug8i4NZ05hm3j0aOK33/aOLXa0eyg0V175jkJiy1i7vCoPkJLssrhGdI7zlovDA0
SZ6N5xI/36MeKSxu8tSnoIjzS7H+P2du1ure//haZXVa4NXMqhNJ4TjT3O19DsQb
OW5/AsKyD7dTFwAmxaGcXM8OfIsy+2Nz/y/PLmQJIpuy+AzvB5F6YCy5s+el29Dh
7scLG+OO1c3dRnX3rxFDG62ooONVb5QKQQEokbvCo9tICNiNmZCI1sJAmedcENB+
qalmr2XBD9dtjHzT+8QINuljJbns53Wu2PzFT4wCwY+3qxtDBcEQR/trqg83Js2b
3iM5WoV2FfsimvbQUCD0NyDMR/Ka0EJX9Nqg6TgblE6bQAOLA21nxL9hOMTYO/dM
mRQ08/SLspo+vO5ZdJo90eGL2sDeeOJGenEZ7sUCYNydmn6b7rNlTI7TPkkPma2g
RbNAZmB41snjf9DlNDska0rt9iiQYVlj8C0UUW+VAuv7Qm0XdZRar82QjOxQ0AYR
h3fyTKqQkZuDRZolKVma93LXGVB8rHg8pbJkS6mi+2cqhQZ7e/2TPoIrIdwiUHV/
YZxGFUVNHSHa7IDMvJXk5Tq1mP+s8ltjiMQ+r+XQ1hMxXgOo+15XbbDRXab3p3IS
XgXryEbhuptMjQANOpEMqkytcZQE9yBzhqtb5sEyY546RqQtfCXB88KrXUCi9n15
K384N83pataKESSt9VYuzxsy0upoHxLe+4IMXAPpn4Mluq+5pFlO3prFAKh4/D7r
85a+0HDNn1EzE5iRazqaa6abeeJ3WIIKdPZ1Es6BBYJ1C2l0XAk4SypQLSFKD2ID
HSyb4avJI6vXToPVMM4ytAFlZAgxPxjka6bF3QyMvqZ+JZaO5afb/oI2/+iFe15B
LjN88nmDbQjJ8XmbYMtrGDNl+84Kw/0G/uVsns8BnBZ6hIrZcJD1ReqExM0OQszi
dpUANecgzsgafW90ZeIbF6oUJUBiNOrQSj5gsmKin296SZMjMagu9NLs9rl03d2S
n8u5llEmzCBTTRnQxAry0wn32eGWNiKSvDpXB1pkj3ZUotfsO2AXLIky1GyPLoTM
a9znKkjZ3PYBHAEvo3gEi6r+Z92IerA9/kMaS4FwrpP4/UAL1vA2UQQSNpkOS+Cl
ZjfVPmb6GTgOIVkkFKtMa50C+VuFX4AzhsIW0fy6439vUtTldE/6+mQIM+JUj/rK
nEWQOOwrns0iH8UVZn5hxByg7XJZRrazF8Z4qWloD4qbQ6NBdmiIaOF+xAC1fiHZ
J75R9e4MAjlJ50EFuR0vPdOHJHmdZ3exofAIUoO0fCkL/QeRXPswz1BCtdwNLpW8
kU/S/nSBhuIvzYEqnR6AR8JSP55ztwQgnZa/3cmlW9PAw6mp9ZVowBXMPCm4tZZV
deMH/8ck7HfIXvBSbEr6em7CC1o8/BBFC8Y22k3Gzug3T7xlP6J38sW6QnnnZzQ+
YDyJLXmB16o0xYT5DSJY68Fx131BtBlcJ/J+8btz/jijkrDfmBsMbPMTWtCXfSHK
mFegIuSXQ8kXQ0OjOY+HCjKtqIrzQ1v6iQnO12+6Q/et9fTo4JDHd1leM+p8sN8B
Wo5pitlE4vCShHsXpbRgDznbEREnRNrTpdyLkndNOv7smdzUhnMc75IHDyDiOQlR
2Hn1HDBFAJDRj7wsUReS6nVkAgNtf2gWnrtlpvhzhBaxJFc/4rLawVm0ZiXG6WV5
UnwmHI0hdJ/jYt8cGWNadDoVBTH0XfyvxZRo9zIL717ArJiw5hPR24DFL3azSBAN
hPdkEdA40Wmox4EMb9cWlPGKlbVG+2gkvo9tT8JbZ6WQczIGs4xlaWWoq8yc1I0I
CCbajLiKiCuMb/y89uQfk9CQkoBe26zc4F4yFRKAJ/YXsEYdhKPgORxsXdBzURRX
n5oQDiNtpHiyi2Xep16KTPZASR04tr9rRonCzfFievwRHAMZ86TzpxTqCBJJ6NJ7
/SHZDjL7So/mLa/loqxBOfudvrJn96LXWBsBttiDJfscAeD4+/GdYpa5Y3duEOxq
TzWgwYTUKYOxtslu9UZFBYw5nm8cP2GoTnkdk4610vTprj3Z1CtyWH9ErQha29Gm
u3Aweb6o1SEBEvF4Lu4ihX7g2LqoDUk2gabwK7RIAbOOMtHlLr2qPFFcCrIffv/w
1nXcb2ydet+Sp7ERhV8YmMq5IOxcEX/C1DpyonVycyRjcr8YaE/7pZf1XzWNcL/a
A/kHAV4ZGCshY/1lW0TfC77QBKZ0SUeKI01bF4jabYwaTMTK0j5PkM6ewCeFwDf9
1ttSTb+ATHO0XQivmhzKbsHdLGyWiF22kd81mTJotXTJ92xHyl3eFS21YIDulcx2
ZTJUTfXoBhzImXDavScAlRv0gxaSe/otBSrnV+SVU64nffjcbepmWqRh2rMW9Cht
VFw0BRR/uJj/QY0WLMA0Eemk0SqIBvroWrnB9d83dB9wk5M/DtHk/lkTvGwgUL9w
fs0dpWGkUklHoJU5s76JHeEyPhydl2C37oJ4PpD8e5yDZNHELFfm7QpVGvuyatvf
f2Swb1yUu5pI4PRaca3F6u0hYMgK8/o452uj/9FrRY+TRqiJWNidZr6fHA+hZFOO
J3Rp1aAwrvoIgfyHMMcMcZbeGK7IQsxebkzY6tEhRvitdaMpbYO77NoelFXQ1yzp
TPwZjsQUx3+GFnjKxly7sAFEpefKqrwLx1qNUrkkajKM1h8lRSCjUA81KABJsK5i
VzoePodE0BQwbDKzFutB2HoJkYh9NrPR2DtXkgeTcupMGUQCL4FPj/hDDrqrJIAO
/MxAqra6D56lfgfzgKc+gwY/DeXO2K3hXqeL0WuG9x75bitlGjIxkLYPBwOCEBgk
rc+m7zdhrChb/FsewSGXUl/YlXaX0hcYIL/jGa6n6H1WmSXIhciaN5ObWOVU+2wH
M2We8/eq41jNvyzkPIkSJpWe/2K6XARXK49C2pNa2XVTQh9MMSy1GtdGmSz4faeS
QI16y6ErCQ68TABzH2Du81To6NcpjzsvAPUnniFKYTtNJg2ksaJwSd9Gqiyx2zxH
39mR9PC9NEq7n2wxV30PFydBsbQDNJwh9E0iTZ6YA3IGSOPDFoQDTv79Ryj/Ch7c
VmYHKoNgeFXzTrzaXE7ZBStIsikoaNqBoE1F3GgNouq80rsDaLthR4s0Z4ZbicJt
XKQRsyeCSInh6Kgl/SrLogmePulNO8B8L0+VK+jJIs/JtlN0BEhsfz63QjRm52Gr
vj+dfuGhgZ8iAZvWAZ23o1WdWbqnJyZjA86S+QRW9tQ6fN1uzaOudHCWahmgcCKI
BjGBf530wrAt2aD2e53Re6neoYpc7ohxzRn3QhJkHRQMUx8MStGLWDz+n1fBwhdb
ybYARG1IODstHFQI0kW6hQTnvE3XEnrctE3w2d6JJJPAzkH7S2K0ermdsr3hpdw1
ZC+lG00r8wIYFMt4TayhjIFdWVlP/ndIu7vy7KB/GrY2OEb+4IeM2OEZZcQJwNiV
F6AnYE8y+KyDSRH0aFupwix/OKrbsCetxVsKgnnp6i58q9t+VXe3mUQKR2VMkc5U
jkyayHhLSm0scYVLbM6tTxjZcX7nsdTIDZB8FW7k+Hlaiz9qIh76OvTCMMLivSd8
rdtsC0QaqfpvuQS2nYBdD+zarE/RA/cBSRaATtrmhCI7Wxp7dziG7gYRYN3Z/A4a
jvy+KMPyJv1F4DUs7O4ku7Br9Pxajw2HWsXzAwq2v8L6Ws+lMsHwRaIoLhTHNucr
ywOpdCItMis9wJz8yMZh1kuAkRT4TJyYUvfvyd8kh9jDEOvutRK5LItRNxE/Hvlm
s2+0oI0cQrRwfgkCWRFZE0q6TOBp0POY7SKuVHEfHpgqhQ81LuQsP75tPx2rerdl
yoKf2WTWDolihNTJRK5N/oV1GupTq0xHrIRPM7oNZm8KAyte+OZY7E/NCG4nwhp8
0wZjfi1NfJS1yoanL/UGATNHIijTt30StbYYAZXTLFSs8fj6dN30iQ6KAeQNI4Cn
JggqNWz7ZwS2TV0a8Dsr1mVmxIL8GofVN4c/EheWEwn/8gNp3d8FKSfteZ+MRtDc
ADvG7nWvhdv2x2my4wpaX/HkpwJp5Y2KRS38bhC5UjRp71uaIISw38djQHgi7UHJ
cnI37OH5DrZrs4OiCMLbUkFhHYtxaib4AXUyjgzDaudH3kKasYoHDPHdn0LdyASC
xujqgjHoWXp2K3tnXqt7zj6ZMbR7IAB3nBkS0VqThKRXb59ACTo96W7DWIXibLuc
ZPA1/xMyrC6nMMtd40ynmjQLxdwS6azBo9RWawJi4Vxv4cocl6xpTvmaKH+X44v/
Fm4Dn4Cg/tUm++o/Dn6dKDJTocwEugD3g7pVj+ni/T/n0wlJLq2V+ypqz3hlQJFm
VcWFEi8Ql0TNDb0UacHrMfvqTyKiedNVJWiDKQe5eWqk3F5jHVo1Is5rvDQzIX6e
Q5tKgHApfSJDRU01OZiymWetWt1mSK4cwsko2oJYDMw6HIG7/zT7D+tqbvxpHhXv
YFGQhnHVTjZugU/7YZQCpTz9k0ejZBTnvxOu1Eju7DvVSamNrPH02uzYXtWW6o50
dhJ9Z2ZE6DGi+Dm4rs6ZU1q/TINGsN52JvOqL6qh3tQsyTjx17orLqe3BxtAxHmi
6qQckkkE5QuWTUG6ylFMQd84F3s4CH77eAoCJa4WQhlFb5fu23jl/IEk1zH/K4V6
u47wfp2m88bRRy3m66Z4COUAkUUH/nIsgF6lRZh+3mHzwSvbQWnD3JBNFyg8CGhR
MzBvnH0b6lMQtoo4mJzc6xNOqEI0zreoAl1vqlhAdmr2seUWTCiRW5PP6ljv4uGp
sXGjE0yQZEevUgXmaI8GBN7NUww0CrW5MA7VE4YIKYFN2isFJ4D0TPl+g6n5nmEu
keSISBd0x8KNsiTUtCSS6Bfq5GuFlhNxLztDZpfjvxEXQpnl9kEzQeTL2oF+9Ps+
KxTdtBkCZ4Ho9dKyIGeYpgAG8xecrxtbhiKiLBDyXr+GukPrR86EfWv/70h6IIe2
Ql38ppjUJ0wIM25gQfN1egaZ6+gvJhMuNULa7PdrEUz7CSLkXijDn/mnQ9zQiWui
N40ESNoi3olqyguXmHoiizQFENzOHT2o8yh0VJkx8CGD5xi68fcj/J1zba8JVYhh
RZd3RAc9hIoh8GL5eV5PynmLdbItFF9Z2q5zARJq86LO0xZCmKEGJFJub0rv+Wdm
UkYd/8avUtdb8Of9RV8w51Rl7M044LRVqT+rYLt8wGz7pOmeTwHSC8YuotfecvZb
5+AXGXy3HyEBYFE1JrbZf0gMMsXKx/8Sbw/ooSlBgXMCbFUEveFwElmgyIAD/ObR
Bq3lqN2rVze+DWQ1ZP/NJI7K04sWbWfwlp5llWik94HerAy8hYg+NOzCDX+VuVCS
jS2ez5E01CFoqUrYfatBctkYoF6v+7fZBa6kim0guuiPVNzxXB9U9jb5GkuHr0r7
cI5Ol9/Xk/jPWgO8w6igbdk4ccWFA4DBui8Cg0p9If3RAlkKC8Jiq3tKZT6RMP4f
mUnPxQFly6GIcvWNPJwMsXllELi14ojVDvo5zXPHt2Qwx9l+bp+eoTAa3cswsJi1
nKjfly22lH/TStNTtSzJXYTwrWznYtWlTWwrpdpvULgzdyR1zFL/TeqLuLmyaMsD
Sejvnz7SXSuHg8cGmw+/ojWjsP3ZuMK1QZTXW23S9MUJ0RxzcjXGqS7maurFjGeH
KDqlNAsbfLwIylYzvmpFo8MHyWCWyZ5bdwwpa5zlY8c4G8cXffNy+JCe8qW36eWx
0o1v5VXMlRxLCYaZ5YvyIpJJfD27RWNOTMtv3Po/TrqEVCFxEkjY4GN43Cy22pPl
u5zvjX9NqcywZnrWu2Yfznvs3gNNh7hDAd5QWZzvjaiKVd2MIiAIxdrKmY1IVZ7V
TeMlkBVGsAFQ0Q3WcHc5Dgr+2ZW76wwKwF2UReWo/LDihf8eG16zOiSfn6JBcvdK
uUnMrT1KP+yVPna0KFa91V1S74CYDft24XGOxJb3sWVbeoDVuzZMMYyl+iY3vjFJ
0ko1V+MUaO0yK7dMViJNYsPA0JzA8yo1rsmIFACybDrEbvq+dRekEGtrA9Qq00JQ
73WSAlN9iEC0CsbphKC6+WM1gCy5mG4N8V6n8Iriqw7hlEpBkQwiXXhWELrhYDt/
4kNsjuAgPyRlSP3DPrdT7PGGfDrBMcWQxYcPaNh1OoeXB0o+pZzwd/ZwvDe1oICk
9VlhbFWqzBBINUrQa2hpj3x+cQQPiNI3tDTgX2LO+pXdqZ0EpSpL3SEEtVtKFI0h
F0WZUuezh6vSZor/m3qtDC5A+2Lmu+b/3PLkKkaotafdNlmErC8QFtbas2is0M/s
qCBKcttM4OjRgkYL3sznzAfalKpZbTkmHJdxRNOzdCEYwaLIt7ptv8m4JmIVMjLE
He+Ti2SfrwacrZm6X0iFb+7/zjPF91dwyhc4QHWs3i4L5csSPWRY+6vBC572lK8L
s74CHKhdGVb7HC2YPtu9K5mSRcoxVbRg9JU+QLFlPof9Vt+FlvNqfuezO9iLDLj5
uL1APq9cSr8UTSkxv3bbcXobiZyVEDzlS5le0JlnuQbWrjCfA0CuZiiT+drikWRp
7kd/6Xn+iIrvsx2IPcoybotB/elroIIAKCsMqGmR77vcJFy1OZhKurQmKTQU91+A
8TnGEYZAANmzqIO2QGXn8PN1zCjgSec9CkhPWf4qT39OpnZqrl9Wxqb7J1n9TCOc
bCNFhglLl7o5ETxObC3n3BOjME8sGYIzSAz8g43+C/jSLDHtT/gvuHv1BFJyDcBN
/iHj0249pUtCh9ag59Q1mICXMhkYugQ9pm+Jo/T1eDPhLDmg02A0f+qSI7hEx4kh
SiM6L2wEc/x06k+llEoqJmZFlVmToTKaY2TuEO+ecg61U23miNbNnxFog6S9bo55
x4deAF74hQkhGrIpqM9xEB/SzpXg+FiK24mK2H1NgYCjoShEM6PqwQO/mnNZVmcL
HpiO9tEPT7lHkE91My/b9EZzMucCCJU0HRZ+6L7xQmUqErYvtEjknMCSAijOeSrQ
EC92jwu/lBB8mIsGyHDEDp4yMF6Bhofw94pGxqCLn7eZSshcYBz2BYscsdt2lc0h
sjYuNScl5xQPEzwTWRdvPzb/vLnrw/jvEd+uRNkq5nydwS4yV/sxixHVVi/lXzq+
GDlVUI0dt7JPWIlG0TDW8e0/jG4crrKcT2DOepwmFka9VNl6fpEE5A+7ldd2J8CD
lxZefvqZeeKI/fNGw77L/Ru3CVMEwWChQw12YuvcYNhdoFX6UW0s9GXKVvc3tjRR
jqmoiuGBpCNdEOHXWK3yKVC2pICf4Ka+DL1gd3vcvoCtQX7+oH0ELPb32tubVjby
9I7GZ7munwrT9HHiRkiR33BAoJ18R86bNvZhj9ABIqieDWjjyWVr2qINbzJ1+Hwz
AEZBXEBZlGa9G8oovF7nYVQOS9fGy4OKmHSPdplLW1GWO0d17qglSPMN7I2xzDj8
KwZfxadEwjLZwUYXG983TsN/0PsnxwJ+7iO3R0bNns+0+FlGSXB1c1gEaAyQo7IG
fzuY+2hUymf975W+wOJ6Ovs4K1OOvC0SZ59IOhHjMCdxi/gDLAiJQ+nJxIU8gMm3
2DXG+qrBkCnIMpuaKfl+EkMN/TU0LvpX3+Swf+2lL58hU+lmfEN+8uC65APovisK
GXLLIMqarqI1nMgr/LIXhyaWoQz/QDlAIJFtjRJJ+d8DC/2zllZXKAA9nb4GXkC7
lPk37rf2e6GNPln+3Q3OuHTbiChyTdouSeFCBXPOvgtFw1sT0y4sMnd+jYwMFn/I
rcq3jVu4+mAF1Fl0ncLhEhDP8cAmYR9JpQQDOtKjxRFw9G/EW/V+Kk7NdrEcX/At
wW8NjbGydpJVxZStzle7I2gn0Y31PPsTvZhcdZe0YnY+6MSHSG44sk2MYcvO7nka
ZrSY2XQFEflCXPQsmCADD7XokZoT4eb/4iSt/h3n1HlOudeIWH3FLYDoRVa6Vr4I
VniPjhMYQoKah9V+gOP5WVCWcs/V9c04PLS+38Tqg1/7GtJX2/CLoptPn/bcOGU9
pdBCh8+633ojrzGWvA4yKvJGYo2QcUO2bGjQGg3l35rl4rLsZP4MryHrvccCjO4e
9xbhMHFmLqxGk9xIqmVeZIYHD8gWBHjWs5pdN3dKKgMQG1/VosVJGJF0i4FG5SlM
9UwiOR7mNLQmBFD8p9NjYxXLAhFfuwFLEtyot2snUhhYALjg1tXzlr08FRjvMsvx
QrD8+w6Nh8+6xgSuVjE1oEXjErBefLqjDCSvsYlU9uQbGNeYrMXDQnV08u3MqUOB
QMjUiqSFW/2uNreb7UAAX0uIAYtPA7jLoboDNN4yjSKOew1pyFIb34cxZdu+3ibO
wf0z8wdwTlj7yvlBWJEvB7CRzviiOynDzIMCv17WDSmK8s+Ftn+NOsog1g/tqs/x
zjJzvq7QG7GXQtWGzb9ITZLU4UDsayp2mzR7LHf9J2yclUcZ64e/6KC7vQCd88SA
0D1eWX5GA7DgVFyCMc0tzQaY8mZPxA2I5rA6DLccJNCZ4Dfzfv69eXeVSC0nusOB
O4zpr75WN0w2HjjTyx76+FkhWVVQF6g5OD3NozQSVxfK1xxF+bOYYwKZwmkznK69
dSnlxYvJmfZ23DbGg44cGnTCeJBS8Nd/dO4Rpx79KQIITTqUw8vCrmpOYTjp0Of3
RDm5IdoHJ8nKICU4Np8/x/OR3IEF5ispPTPOIUgxNlZ3O+0WofSVTRu0X3D/Bi6l
iWRamfFh25zLdhc5o8IfevrDPNN7q+0lpOK0H4ilu0ohwiakL8QyZgKB6Pt4kZN4
DlrZs4kIkPQdFlVkwivoEjAyfKMneZCk2Xv44fzgYojihguaLUscYi6nQn2/LZle
Q6aBKz7syAzN1jexKpx+W98747jQsGRwwrDIYopRJJl56gM5ukWzzdzRCyCQrU55
BS/mgimjCFdakBHz66jlpJFENFzMK7WE96Zaykl8bGck3FcUoyjQn2APToCWCdgy
06NRL7DwBQhPQlCvK7ZvIlnsuZG6TtopdpalD+jspVB/DYKZrboXTXbY1DkMuEZe
GThblPOwiaSWceaS0w80/9DGrGzPxclcn4aHwiIP0fKtRnlkmURQ0Qowmo5btUTU
kgfuzwseS3ueqXZGDLUGeWjagFD80fQR5tUrdEyTATykZM89kpYyqBOSKdhXvSOV
+gNuRwKFRu9mwyMsT2F4lQ67+Vzq9Paz+VDyAmiRRHTyIKVKn1LkZG3gWuwgxUXt
yHcf+Lov2vhNgEAzrkRn1LxF3UlUuLcG2MEo/8+W9tVTXS8t4WYbUxh4UWwtyiff
IU1yewbpvb2NxNX+zqCWkNIPdRV9VfGlai801tkEA08dL6zoxufs3voH/weQw5CC
9maDR/6PL6e6twBZdcvdG7gr3uvzmfCdJCTfnUSSxxxtKcRFpI3enByyLMKQdqzS
ODpVORiBe1g/gMnzREV3ivBhjoAGQL+pndbtHzySQwrvVYB+pGNKZO8ZCqm2aWGK
a4INlV8R8vKDhm9cKwSGf32xoWWkzwAq5OBFN5grKRFClpQL3CqIdLjGgnbe+Y7X
Ne5AtfnJdIzYT2Ho0ozj7mOM3mJwMOgwq+WsaIGF21WaEwgB0R1YF6cjptgBhwLR
BQEFCuFD9vpafwlyM1/oNGQRho6grpUdIThf3NBO7hlx0gItL6bcTBCjeKEbMY/Q
fmtPf3ZncTGA37Y43NRBU5iw73Y+OygQpq7WuYS2J1nyK3Prdc3oIkRAyzefkAqA
tQOuO4/pySZ7DCjGmw74jR07yfAB6DBZLohUVvMW+POTRvcBWziBWEXc4iU5LUYm
xhaTf4+mKusQ6EosGJUJOS99yD10JtSXVEEFOolcPleKru5FBYSplagCzSvfy8TL
+VyWr8xrUNwr2ouIk02vbIkS4zeeKANMyP/1bIcQ7mGd8sitdqRt8kl4m5aNOy8C
jvb1rXJOnUd8ZCZg7SEx9ab2SizBYGAKhr1/v/fvaG7Fdz4d9+ss/oZwio6zWWsF
f6o6K1OaD6ZLJd47FXGnGtc2+iuBwZvnzlMzuE4k4DrjvBlnnxYOwAw+K9KGX/uF
kbUD9zB3XDYYFFsC3Lwo2laXXERSTRv0LexAnETlxZcrG02iu5VmFEaO1vRBVVTg
TzksIIE6GwVb/vHb9IJYgncKGgbV5+kcRm3Oen7i6rasaL8MnXXUApmnaEXQk1tz
nJvibalP6bZWYF/tfM2dIo+vExRhVj2JIuNKlR8iqf5npHVRmxXeVTkzixLp5sQh
5OEZbYYtbstbVjP+DebAVeyMC50/xpoAdpOSKFaibnhaaeH3ZnIz6l6McgPJnx3u
0NkjiJ726cEF0VMcdaZI68dB6tcc0SIm+sOQtnKmoQI8zauO2Q4s+jxm3DVzv5nA
9BqnwkVF6q/Bf4B+EfwdGhoXsbCKx6u/uQsw86FuSxpjVCJD0UYWx+C8uuxp7fPp
YdCVjgVOPPgOKmuh2UeYzeg/+bv1CDid0fQy1RV/U+HY/mXqf+pUia0hIcfxj1xs
1o6BVN5qaNgYo/Db28m0DzZwmXetDdzwu+pwJn5DZ00RXhZrRXSY0T69cNa1Mra9
m5oRlpP0aonJm4r+Q2CGjBYO2WNNfS2c5EjX7QzEeLUnwjVND0rTPOOCMgFM+Jpu
L4NUh5SekloD8lJaTFIWfqp0zKATsFamv8veA2Dos/crKdJ4biCbvqu4W8xTjcZJ
qknJid+Yj7zSpyVZuES0zi0OwspMM1NpvDRLIg4tGSprTqWt4t0dmw6u7DcC8FfV
uTKrklWbSQBjpPrkvtmECZG9wtrKqv7+hMWoK7Z19a4HRtrNnFA359eq0InlsRA/
HW86nP4DgYKtCnWnGGEj0hCDHHztD0mcBmT2OouqVZokIkK1MLRYz9qmmKFRuzsr
g9aManEQmRlfXSy+O0yE9K9giSx/dCTten8jkuJURzbhSYYi4exUxvxBKaBLLCHv
xfXQKpkWCbG6GAwOlh1xw0qse2Wmw/d6k7ViJedPv9ZM8Aqq0SEjS5wyPC9EGV4I
7Xszqq7B1wrm/KnP3EvQ+prM4u71XO3K9MjP1Rn0AU5vahr9Uq+UU7jT/eJFaAk6
g0eK07pjnT7k1YWR+/sl7RGWAYVQsQ3FvqfEj1MMcLPcUVi0z2V4N9V/kFRVN4H7
nRSvrSA18Z9lnqjuVFn2WlRMFpVNnhl+ogzkMujDIxifZMzi7ecEvV7+sHLrjHwf
kdp/9extyaKuQOsiQHGhKzJZwcyM3BQRJHW/sKFc1TpA3lLpQSE5NbDSyBEtJv+F
XvS5JeBjwVgs1GawbP6Dro9jiMS9nhO4JP4yZ9C5HRig1pavmphgcaD+OH0jbFpf
uPDliPx1/bCRHU4fHXSD57Un1E9+9whlKYyPVbuOOYg2gGG9TvpcDxJ+8EW1opgO
wXnGapmSEI6Uyg1xcDqPizpUWdWTBolkLbrdCGAzcyElONG450oPdxo2/zdbYSvZ
FqmKJ01d7CtO7MVQBkPGyl93EF+TFCSVhbcM3CjUdaKV0I2y6X125YDPwwY8QRxy
rcOs0ZUXcD03Bbzyxl6SCWh8dcQUKXf6TDdpH1XPJ1IvXzDckV4UlFzH8iu7KeJM
Kngt949Oad/4H5XJGChBoNuDukIZcvm7PYX4b0HW1d6enmhwy5UFGxEw+zr7/qAH
So+P6Cnxwcnu6JQqU+rVhyaAagnPSJTurogNbuGj8AKcEnhAaiMPQYGSCsVgOPsM
KMMxWGrKepztHgLDao89XOey9lO/z5kaxJc0rhSflY3Rh77jXyppeT8LE9p3J8xh
PDGdCl0Kywv9UgHjmb/Vfvo1JGifd69miZjZrvVyxPQqJIN9UsYxgR+/APF1x21W
4UokMOWbtDwDXTMaQVHdusVYum1KGZm3xSVKSPgSNA1WWBguAXVlUiDjhPqsGID5
UhGPBF9DM6vOOQ47raDFxAG7u1Qir2ToZP2O2k/vWlTrz7edJ44+WAYzFi7lZWa4
2uhzE+c09qTbEasHvmeM8sh0AXsG59LBLejv1EU3WwkenHOiJNRCjYgjnGYT3qHo
0OwBJ2xBNcmxIS2HZ4L+TAqBqUlAhVjmWAo4H5aAZEDVBQU9vKdqf26UBGdiEWKJ
3eG7qm8ypS16ZYCNEgA6n7GAWNsMnx+d5xMAeiHYgRtfQONQdLjdXsOB/GsP4/pt
7/n9qTzUqVDe6xooj4T5H343WyRGDQzfENiHkBEJ9zHXADxbTRKP6sswUF+dFVMV
RwSOtcqPUnyJtSdm5kdrdkvREfmYbdx0AUAuU3rv5dmDuoX4idDs8puUe7WrRbQp
5q+9PjwyX7fkgcZY3nCqk9oR/j0OvY3PSEUq+2l7pqlwyuEs6kaoNRINy75dPjuP
dup/4ANqBkkpprJPc1McicW/gy92k2tH92XOCAAY9gnEcaRcLI1Lvr/vxKp/ek2R
9YMEPJUDUF/0P2IZ+FOoxUWxNuuzz/UcO1WtzUNYvUpXUj+2PIJfjROM9QsJ7Srr
cack/OQ7fbh2z3FlESY29F1uWTu2xbEi13OiTnXAOoBTC9mx4Vp+7Nnuql2I7Rlh
BwPzxjNxqs+8+7W1O8Bm9Q9IY4GNnYYm7kYl9V/wab+NjOnwu9ZrRlYUMrxHrPUs
t37mwjWbA4gZ4YcVsjCKhFToCJwVPtNe4AAgNpj/L3uwJUOpySb6+LskQYg9FTOc
5KQLHAO9c6y6TlTqMtUBQiMpoMvoheE2dvEHPd9eZZ56uUj1Gz8aYXLnbku/2QL6
XO3VBur7VWTTdoc/gsp7ogLzcMmCRW17Tum+YfwuEZSrwZqy7JcZBT1FveuTVZdb
bZC/Rmei4KQIBfr9kv9fd/BL5cB8MQinCfpU6/uOeFX8NtaFl30OEyiTYX+SFWzl
tVj87rKcFh+gGi1cV7X8lqHVezq7e3LA2CW6k3q9niISawZR8QGSxo6FoG4K/GpJ
rpxURldF53pfbYjjowmd/atRvRqA8rJZdXBNzIo/tku7qQiMLWDxzUyOQlNFw0b/
iqLbPqG4wxOHdyMXy4qoYdhUjl5zd7H8hAgaZCSioqmD9jKFkyVJZnqBESZKRfXb
P6Ek4dqVCHVtMHrQDwz9iOBX9ENuiTQiQ7teY7J4Mk+/r3clU63j6RLdjP20dgvp
jnGoFSiDhK8rFA8u1tS/+05LBrZrgcDkKfi2BKHKwqWZy7fWqLdBZrJJmWP0l+KU
kyse0qrVWz79lCR9cl8YOexS1FwY2eFu7pc5U0F4Ekb3elCxCzSbAnGZbnHJ4WXi
2QhtAjyKnWLITdSFo+X8QIqYZdZrpSlnPWz4pOg6u+7WPQ+KSgrKMsoOF/uH03pf
ij9bko/E0GDO7xjP6hOaUyC9eq3aCNiWFZHWUbKrcv7olcCij9PzB+MfbqoWBW6E
9sWuuu925xkBBcRzlCXJqVo8lzdHZRohVcsqEaEU4FIv3ey9/AKG0VpGRT5JGsiU
51NAOuX7olH8TKwH2EKCmo+dgOFRGmFt24w8sCZtbN1tfxYpEHjFRLoG1Lxur8tv
nzjb2p5dH4p0jQKKNK/7AhcB9RPvN/nC23WJQKoNllZI3pFNCzQQkNg26INlDAmS
zl3M2tly2yrfmtW+FAoCNZGR03LBNYiGZFOFLb7bOWHkckPhtd4XtVTNtp9NeNBW
qMLUr+xyaRglFwAX9ZhBlCVCXNVJdOcSfnKJuvgdVsQfxPFf4hXhNbHSVeTrQWmA
gTdLQEfp288gDiwGF2RGsZVrjWcTOvEd6gkJqOgpDFB7LhSDjBmbqmZqCm8Nphhy
fg2Sj7pgtX3qlws76ZXw1DDCLzNpktIT9UkAUt4iDhWS8EJ/9/D5ybC9qPKHBaI5
teRDKwpRf4OglKgWs5nuXi4pW6NLe38ueek1NrtaFWctY15J4PK9/vsa5z0L5n+B
sEpfbfkEvpf9aY9ioPdoWpwyFAeNBQp3Jgd2XWOL8GtNKe6k0LaLBWJLHVu7abWa
clfF+bV69Pv3D+XqZuacPL4rxSd5u255m0j9knP6VQjyleS6Me99lWpnVjwFHFhh
Tro9dSazN/jqDX5Jy/7bwfpuRlKrlXDDGKVZMKR3w5OzjrQeQ8E8a8y2CwtTTgx6
9so3ZdiTw1ZvgageBoIohXjhy3ce2Tqn8VA2L1yU14iP3ZcZhOiXtbGOF0EaZ6Wp
kQT49Ab2ZlmMJ02EkE9bOci0bMYZ0FfFetAyXTTca4FbF6xpffiVbndrn2sQP9WR
UrieXpVb0Jw7NoiyWF7H5FV5RBav/PWo6AX21mUYgDOvmcMAGw92xygvpoFQMM+W
rYzIXfqKFbYNB8vKpz0mk6wtVjGN7UBuRgwe0fQYY0h4Zmu1i4kP1HAKMHsEOWt/
QdcZ1FGCv/y+gA9h26Gt4LYefCGQ5oehfTgPS9fHQNasAoLIXxN9HHH02o1WYGWV
S96bZieVnLRKeX17TY+eBzsfCuwnDIIKGGwpit5K+CMCCo2DETdQ1WsmvBnO1b5L
1qTb3gXqdYte8+rGpfsZwpA2wB9vQU/fhkRwemDIWV8f+oJYmwKBXIfPFrCEXgPr
O/nIwxjY+amKPbtS++m7X9Cjzv+ZmBxV+XM6YwrcRu1VthRv2rGIEFieueHcA5/o
AV9a45EzwPLY+AQkMVDwnJ0stCS10W2spd871SDnpERod6GsJam/opKaDfvaW3xq
2OYUK5U2cTEShSsTwHkp5kNCrgaKNFmZem0Zriry41OM+/tHYiwdjTSpDblAPyTK
XsJDRd699DWFptST69t4KmiJeb+Adqk5ztgSsDGVh5ncsSYJ5dhl3hmw1WW/2P2b
odmf7Pr0dqZ2IcQBgtsWr+EyL36h5P6k+oBmDuV6pg8hzVMyYyVz54C1PmQZXxfL
NPu/hleRTnIIqcMk5DYG7rB/Fh++4eVPdMF8Zne6hP8iYtWRfQgQXbtTCPSpjVEC
GrhZ/YelZppsKLGfT77LsmDkwCZYOfuuyUQSTJ0Lkp0blyYtODtR1FneuJVVdx9O
9xza+4yAT7by3zcKcACivJc5xiPXupoQ5mjUs15WjU0fc2yz9EdbFqTxb3kp6Hgw
Q7B3gp5UgzzBxgqoSOBUgwa2tVnR0wex30LyXi8UmafcJo4pq7z9fcwoMJX8Cwsy
xMLUqgvdi25nvvIYY8aWybZU3IcQwOjq9N6T3mAFDlLWZjb0Gpb6oldZiW3KWsq3
MV14b0x5aN0PVu6UCYS8iatLyuFXSIoyF6DUhYp3GqSreF/kjDwB3X0m3+oMACXd
O+crHSIsD/tVqTmyHzBV3Im17sKMIVx5aDNm++XKEDf4iJ4lFRJ5dmpiiDSuXip+
PfURrPwTDsT+wSljGMGj8ZYEMcxuUlprlZlg+o/sT+wpt51zTlNkpX6d/o4CHNgT
XVsq16LQv2fs2z14M8G+W3/oB2WCnKNnUgP6tbCXizautqZgC68Hj+D6WO9DDDN2
OWPPB+Me0pC8YLv4MmAbU1Ho2egGQF4S148EtY0+tt+dOtiUif78xi2QKYFUhJVk
jctoC4HW6eMhznhd7zkg7+Ejqtr7BgBMEtTDayyxdk5mSuj7AnVYnZuwI/djHcfD
GAvzKdOlBJyydDUunf0YjDAmpxeNb6e3tM5njNEAaMqgw9e6G9BL9apsaJGyobax
9rI9+pD2wc26dfEex4YtpqbgxioaV7z50KiFnuRDuS8t8M79KuYsnKC45Jj5oXfv
Af++fmOF/VDFGI5ESSBT+ryDGGRL189UiR2b2ptLTewKvTwmcqMxAuZsG5PH8m3p
/TwZhpITp28OWc5JXGpzXboLk4g4vxHp5IxE/szfw8eOl4p4qbPNN0GCZMqoWjXa
V6rcYondQEPWOvX2tAM6fJxc7nSS2XH6n5aki2h3a7DYrDVdJZcQJ60e99Wp4lsf
JRu9RNv66UpGnL+xvI/Z0nml3cei04CVupr7HJyojfk6b6707Fyu1JlHkJtzivIL
AB5djKhvMSX7pF5CIvtCOZIwlzWBaxIpUTw/DGACTsatAJHKat/672nihWpdSqzh
ONcVhdR8CgOXyulvm1hBW+hu4o/u4sih5WHm9LyjLB595uwFWHxDMUzLryKLQ6aW
PJLdAMaUj+KIJefnm9KfgECu4SmGpGGh7DZId1a4i7DdKTWAtjjcfJeNZhK4xpUO
H+BRMgzoum7KVqRfWIfIvXfhlhAo8R2w9OOWKItWEnH9+4fWgm5cM/+DK0rqAy6U
oFgvYxL5GIBVsJr6v+eSBeOt8tdHtKmeEjutMGnlfHQEOA6+H/9d2wFPULzolUAT
BVXKWxWAMOYXhxOiLop3yFEmkTRf+7c4R1mt33okNzCiqCbKeXklOK3SyP5qOlIu
+Y2nSnC5lA2U7NpXUqcBhoXoOrua1nXX0wM9KrB4HWvPEGLetBsMzRL4CIo3rXdP
YTc0vQZhyQGw66PShVeG+c4qHPoSXI5qkD7YsU4VVFHE0qqsFj4b1i7ZImSbEq+P
HoqkHIOmXMSDjLHopiAtogcMcbKC4FnaE2OJWqCD+i3ft6o7Mx03eg3Oju2rV5TY
W9o9bWCC1bCIjOCfqpF4CFIVJQbUa4LbbJhfT60zoi/PWd4vEDnVlKU/SbVb/kGm
CbFYXKB7yGrJDqGjLtSHzdjcoxh+BAFSwwdYfmA11KqrM37BR5B9Y8YhlWYomBCj
m+L6Lm2jjlUM5kMii4zK0ejSmi5wRXOmR5o9avWM1cC8bwiQE/th2HAjc6h951qB
9pI/aXi0bmWs1a7e/8Yn2O/1UvmztgqtuxSJOAtKquAv2X7NcL5HXUIUvN+Uhwj0
+9H6muU5LX6inCDSQGxjhif72iPoSdMDTMrn5/9WfWsdgem2ZDJkKX7tcQdv+exn
GTprWHioXpFYaDlfpOZ9beLyXm3c7ZFugNLhI45dkzD4xzN1SDTDShi7lXZIkh47
Gdydl9dyaGAGQvPwqcXcFzlBMp8Bk6dWQ4hzDRGphxKftpmMwFKYZmkUm/DYH/tV
5sr4xjAqBjbXAKDHScKju9BN8NxkpxiEKHFNZanCpzewXnqxXtHVENzpUYehXz3Z
ALZyt+9qmgUzw9URyYKTOU2Jya53Ji7NiU/xWs0m6ccoyB07ia4oR35TOM6COEt7
33WCc3uZGruipsSqIbuYBxe/Ohl5kVbQ/xjN5Fj/eM/EZcczq8e0u1e7paSReZVD
mQ5YjEETcEQo1OtDtzxd8DhE8CRobIqrKut38Dqok1HEvUFsYrzKIKKeF3wqXLEo
9KIsRl8QiJjzDhdtkycR0aukMrfGy8uJHmitSJH8faykaTehWnvzLw3HXEBZiFrr
/yDuFasRlNl33ZNEOnbprde30iV8TJWLAIgNSEuWqzTQhmlqhetkE4rP/AwpXwRL
6dBodYiIwqE155KRQKbpbEnOH0jMKI9g/0wyTY6tfIFAYu/RtkixelT26+1JfUC0
s1tmmRhXtP5/Pi/WMEoMwKjjNfcVVj6VuRsPZSYc3eJIT6/ufl6sgkfNZ/QkvEu9
YcpO7ceO9vH1ZAtnxPTWkVZKacPjwu6ari0JsFRbgjMh+N05R+7x/kdUbjowra1Q
wyro4ptKBjlHe2ycUIMxrOu8e/v6dEQU2BtcspyFfl87pmyLC8BuHpYyorGnfOWm
BC5gjOQ5XdCEhoR2y4bbrkV4MhzDjURTVBijs+a2T8kt22uWfyvPpEtgM1VkaCrB
nH3FPsqE+X1zceHRT76ozYDMZygxQopKluSp7m5PeZ6HwSdMsq95Ko+hz9VWDxSp
FHqBE9/ddRDpsk3FjHjO56QgxoHEpDqOHC7nrYc+JKY+u4npgIv5FGfqPP5eDJtu
iPINd22f47U3OAOvOGMq/8l3N8ZKiLNnOWfNos5994pCTPYhaGw7sToGW13COVg7
R/wqJN0tyj6edXIcX7UjwzRA/JxK9AP6uk4H1xLeogvZ/lR5aecd38OrJOyrqDR6
RG31rf+ri0uV5bMDz6Q42AXs7ngyhZIERJ7S/OZXqN9W4n0b/0+uUPrAj3CPr/ih
l1gKW+jtHiiUQAMFHTR7OyDh2AyqmQMJhwaDT19T1rr6l/hqVbLKPaFdr/SEqRQy
yeyk7ZWynBXa1TP19Pq8Wh1yczrbNQVeXoIL9jcur8EUSmx23KZheLYbAM7Y5/1e
XpDDek+3Abbd9bbCUo7VuV9tG+GNElVTQ2H1Q4zWDbkHaW9jzGIk6D+31tsgJkDG
KZqrtxrx9ArKnjZJPLn1XIjvcLmmRStQ9sfpbnv9b+892jMkqJgOnca289WHzKLS
y89jQAsX2tUKTECwU9axeGDrlJ2sqdtYeEthK/mEdNDjOpK2ZIPlnMNCZyBogp9p
FVptQnCK4uGChBCJfqCpYZORBGSdEr7krfHwHlKKjU5CHRKGOcnMKqxmHqOEBI+T
4Hir4o6PksnGJywUmhAcFDhOwD4YSImo90yZnyBE9SeY6B41h+BWcLohYLOrpIkD
azOs3H4YUD2SrLwG0XTLgEG2jzk9cEPTU8LQ0NobL9hBtWNX0D49fAW5fNTvhmvR
DJAm3oy0DhJhXa/pisUFD6G228Og4FC8k2Opwl/JdYZyZtuPms+yb1b/sscnHq1V
KU6cGC2+HNePf2XcoJAjZUU5AHVNQVS88qpnqroN8txX5CEnblSuDfGrZvLti511
VBEK4x1yndFXMbPTS2Vl/Sf+q8cfVyI1NAEOgxTeUZF8kiw+ix2dr2Oda5rz32YJ
o4/Sp9gODhO2oj9k1k1d7ialAMObJYHUhGp10XUgen/JOn572JsNR51lHIVnRchf
3lTgZArSVQGVR/jt89lr5UElU06Sx9m37lVcWuRnZmW0G7wdrFEX5SPx4hyG3UAa
FJX6aDzfMJbjcNZTHQU3DhW172higTRSTIoQkhu5gWHv2cS/LanyuCnIN/RJpDHL
NlBfsRAcq8rwWhlxnIimOfr1A8gEk27KkGH/dRYMVyjMRPm1u3cNHvOgckqppiZN
XRvjgaBj+dftY474ad+Gi8WExKOLh+tMzDisV3ljvk8kB3huZZPtHCWdj9d81Rmc
NAGYRjArRBnle9bOvbdwUw2pSRlgD20InyLaiKtV5Jg3K5i67EHQ8lwfNLGiISNV
elqFox4l7Ik00O8hybxmwPnB3aVw8X6xoqwL8IfSI8QMK34Nhn9tBNtNIl4C5GlN
jm9rRd6X07dt/MDzL8zrjMylN1CSxJAfcgqJzyu/ueEYbu094lvQ3dYMk2yeZQSX
bg0itpR8lcBNyMhNUQX5pwMjuIcsMXZ12KHZPWVpHKUq20LvHz88UiUro4cy1pJM
y9DMU6TMAVKg1UYL3A8u1lf04sLdXcdAWANDN3Lr+EruX/8rj0tudqeRdWuMUAR3
FA5I46zYx7f6HgZXLWTc4PS1eRkafErr1eJV5wlApOEUQxmgD266C65lrOXtlmmz
Rd4fTjhFX8dxH2zZoFHwHUjX4YUumzTDiuj2lUrTc4NsOy7YLLhYoHCkBYxTyMTG
/jODpmOzV8IebpDvybuTy6KA5hvPFijTt8Xo56brD82h3GHZFivbVbC7py0jfk2B
UEKmktL6mJUjsqFlQqI9G+23WtQknvzx/bhW5HCWhAeTtngzirqxt2MVwQygITDl
57CsI64JVkyNA+77C4FaFTGce5jvF5hq2acvOs8WhbVLziuG2HsadgnPxbmdyn/Q
39lvznhz8q0wUk7szsPaSN24SuC5kHxZ1Pgp78Rcyq6HlmwT4hVgdA1eJOsdSs1p
XehqCpomH5Cpfd0eC3FetQIUf9+fMtRbY8KCevu3JHjNmJNy+k0/eTxG3onyBZwP
pAK309f/cH61hHyD5+pZ5WGvO+jtpDQ6LZnc634UwPF4uQ5RMkmGClsJoZlXQTXi
rJ2rtLAU/ZCwFsYyq99R0O1obU93HbhrkXtZ3uoDS0AAHmLY3jm38qpTOAOMNTdi
bMZz/8onDg7OFl1iSEg/MYACAVgWJqu1p7YJLeALxBmQiQrioe2UBl06AZpvd321
2JtBp8V0izKqxSvuwtv25l7nicKDvNEZcwetm3HkNjedSKLYLc6ya0KNot4o7LSD
eejyjz8DGZY/tZY7RPRTwqEp8ANmMF3x5KPKwtc37NnhFQymcnkoDVbKao7X+r9G
v53DteI+qi7MmhcmGBBEimBZ140+fEaSjkdSHMcw04CV7UjpyJJWlMTbYJUmHy+b
Ooe6FFezPWJyiDwvyRXJJLmpWRMPWcQcGw8h2+Jo4VK2vxG5QqpgJYtw92C9Tgtl
iEsQYPHcSdS3NsDup3e/kNvkUQ94G/XoWmXB2U6geeQG3J4SXKdvQi3VvsKw0DQn
hKs4RGiZf4dsulqqub0BhRUVrimgbesn9VfdWw/MX0W3MWDEC1bnLl7pmEsRSfwl
drBPNOvF25mjKI2OwufDPCNxtz+weH/m6dXy8cII04mhtVGhK5GpiP7R0fic/UIf
F0TCCOzLQuNwlLrTEaqQ3C4ghVKvwJaTW5byEeoNr1yMISQRi+OqiXJFGXCEP9YZ
eAdOkf1e0LBG+QmfW+r63+PlETZRHtZm75EkUpg6sPcZWNPcMmaUxFlLEuJnjAP6
HxUFEPQhLb93E9OZs5Img5X1CIYR+IHxJjYw3oWb1vzUKCAMpXPxq7bxPcoQQXt4
CxA+vPeVue57za8L4Zf1AqBCv3WGiQvzaRgmJ3+OOGvaW/Mo83bV/J0KCA+wMK6G
HAXz4baVDqREyTLMa4kmwSXxphlsUIrx34LrDk2COwWdZCqZaexQjDgKeOWE2XnA
Pqg2T2e9g/ivUX6eo7+Q9cbigEBnpZBhXDws4WlqS+Gp/GHcRCYtaoTUFZaPB6l1
nN1VVqDOSgYutgfBbN48a8TyYqVmjsOB6VibD3YbnKAbqvn50kwBZ0hjdMRy4JQ0
4cD+rZ//QLgSyz66LJSecJkmxit2BYtnfLF198wo7KD4co+q8FOWo6B+ldByY4Ms
P9hIrCsuMPzLLt/LvnP1cahYVf+jTJOzJXEICQXhOoWKgHkZlj8dFFwyI1sQfEtE
Ful6z9koB0Hc2fSftEEUjOjhVtmJn/3qAZdulyrhoCiHt43lGVm4VfTRAcY83YH9
DBSkczL1OyynjH6cbCLp4KT9mu4hl1VabznsaMW6St0Zk9atHgnijeX7F79EkuRH
QGZhUgqKbTJaROOj22mG0oIL/HUDC0gLu6Rz/aoehtMY7l2Ko9fET+FKQjS8DpBG
Z1laP54zobtVmJcHO+IOIQB/UEAI+PFTfIIoeS92xPhzv89EOBQY+SRIzrENlAjO
qPph8EOC0o4tdhrl1TZmm0mUfFUp4PhDBz1xQFXGvvzmvswPzR1H2cw/fLMWz0Lh
ZW3lAYRav3R5wjHp6Z/dQ3QeNUCOGj0tHCbS0P/QiIn4s4V7czYFnxJEnAoW3pHT
7LQTtG+DMsN4QuAY+xWoF/PQs42CqjaEKiDHwIq4M0Fu5dNtaC5VodLHQOfeHdda
Dtwl4uLOfR+zA0kOfvVfOcIY1RaPrTOzmwz4YvDprv4IXPubcrqw8+WE20HTUJBH
yXJB/HOV/0E8g7RYgKpuUX5J/7qxKAQt+Rukb3hg75E1MV0jzQDmpchtFRanbEo5
nCYyuvl2Zlj83tkn+RnQ6BKzBMwmU8THUjTW4sWmU7+U6JHmyYpSoj6+BvkIZkz3
FuoxAlDqQ9cUrBKVwCk/KIQhBhJw3O92yw32k5vkW93MS2Vxb5prJB7RpqDJsu3D
hGUTpGvowrgUEL2l3AATsJOcUfxu58mimo6PJiOL963feepO/TW9Uy+1w+RVPMMM
9mKSd3c7iYxYrKzbhmTpStBQL7VGCCIhh31N67O8NNJrcUCmtVIAHBVp0HT5DJRe
5y9a0QGxBGezg3azUgFbZ7c54/USYN3SYSuwIxX+7qtNpM/+s65mBvz00u3ffRdT
ckRBSzVj338riqcuo7+3dT9iufbGFBBcrh2C3zlLJAyg7o1OwpxLwthQGLVYdwNh
4FfPh926sdYodJCp6Eow2lJDOa3WeN+9Ldg69kj8L1unfTyEnIaxEhZvDE0ukd9Y
Gndq/0FiIrYR1hvydJay9/QNpFqOjUQjB4Rdbk52rrfNlS/gohfkDRfvRr/75wrh
ANpJLP6wUe9vZRA9cCX5iHatA5ot6ZZaDAZTOw7SUlmmxhS76zUxymf+6C6X6hzZ
D1wvt8HBD5gnjzjsYkbCvKypsfYfHsnAOpEGAEAP/gWwk3eV2g4IXNZSJQB3GR6Y
kfofERjg1Uip3dgv4BSVqOivj0PIcVmg7xp/TFb+oJSlI8B9e7SDzLQK+qKIKfYV
1/K8w0yqGFS1PwwKDstfqXN8joq1+cny/rqNUm58JvQnkjjLeeombUXdGXrMTzFb
cozYcMOo3A6+e1/aogqzMW9T6AWe90qAFSflhFmcC0atyBLrUq7EvKT6Fjj0cKoE
y1enBt/c2eu7+hkeKG5RJoi/7NP/2pjWaJRbRkM7FhIeqtJS8AaIibMdLcez8FkB
CHCwsZtBWwqqFT5ebnQh7go8jEk5zpDQPoaOaeRDkEqtbCcoy0eN26x/eTAdv9Lr
IJsd6Z62m96R8OxjQcT5iuweviDGV4vLg6ifHeBjaTcSv6F4SehhCvoWFQhU0zSi
gxIvPpacNlYyjdhf/PyPBPGTsTr9l2TdB7KHd++JVydyQzM9D24hyrey3jU/mzHv
NSivno4Y2rj8y0qklq4Kgr6JOf8UqNrm3Fw4BzalXs55PE3U2fK/zIiOh+v0ypaI
YSQ3R4DBKEDlFKVuFL9ZU25fiSJDtTuD8UMqzCnL2ShIXXJLsgxnbpxw0AWTLSHd
w9QX4qpUC9TvFo1tXVC73GtqbhWSSMNTy5EKclOJPVVhP8GLB85ygEmRwbS/yAmE
IB7diPLP5NNNu/mciXh3x1L4efHuwFoeAHYf1LurAUoskNmC9l4bx/5Otx8JLVmD
Qky0VXPm9ugNH8LBxGR4WPWdxBiORarYbrG5hRGNRewaapq9WtIm3ukgSGOTDJFY
ld7XPR6rBc/r07U3rAzcoD2+DAu5VspIuyVPBMDLlvIAA5mmpCcCOoyF1onbYhtf
cjsH4j73J71oKFqZu3nJjfkpmInZiteRCQOD4CCdelbbMCq1S77h+PxvnyLFSoDK
IVD6J8KIOo0pdeTrka903ebVPaMuenypFy+cdJZTihMn2iXvtiMS4nxixI1t8qoO
NYghxxjy3iekcO7tldWB2sPtOv2biczZtdiEi8KkDaetbsPDO9blWoEZWtBxDPLk
AuhiJMOCG6RDuzxBTwSsbXtqoi3+hPmKeaVEjIz87alQX5IrrbBQC61/BR48BxRc
RJElGqlnSc1V82pVXSisab2y8Qfta7E4wst6OIoDfGCCAKF9R0l8a6nDy94mvRcK
Yy6ed5TCguJxVuuDiJByuXHrtovLqqFS3NjqwUeCTO90+Gmm9cl3knZUg1RFP0Fy
IEKS1QtVQhLCq1nw7TCVOv2lJR7V5LaNDW7qDguk3sUeaWeklsMuTq9YzoeIV+v5
KtGC/Lt0MWWbyXguhbh36JgjQuzeYkJAlC7fMerSXZRxwmKUnocmvuAeCgo9pzPq
Zv0oh2hRfd/v9y+rxB88q3Nz5tHEi4wIv/dQKGTTMSOKKXLSIguCseSxVclr0Pe4
uutTrlkTIN8jsHyp04zgJQcXrrhA9ugCoO75IXnTgnCAETEXTxSS8gL27XugX5gN
2ZCcRPhJWphY/XVPHz6bbxHaZbZpnZr4ZHPXPcfCp3JyKvtitwYOxPSP88xr7pv3
etLpFc5NSvqnZuK1IjCnENAcofKnXfaXLLwb9HC0VLkS/9nbSeSEKLAb/Ijyrkoa
zucwya7bQLTZY21hqySgirIFwZyzYHsa0/kLM3TrL1rjFPhDo9BylEFb17+oY/w+
qlf1DnIJ6572l5jnWkpeCuGrZgrJLc2W7/bGbvepYH0K3cYVZ0NbD8XXMeMA1OGY
DemIt+PKDIPhHQ0lQIT2sfvXcCws2DcU/U4+UJZ+fE/7O+ckffWCl6qn8V+dCFb8
razeeikMxZWyct63Cg+Cl224F3SuSoxcfVnh8jZNvdLdcpz7BUzqriC0ZdKCaKo0
4DCR0oxdNhl7os1e2DmuQjTJ11dH9dUy1VfdkKPlkU4j/TiEq/mITiRhtspsM+OC
bN4DV8V4TbKDEIWw/UbFjoK5+Yl51wCm2AP86e0JheXlsKqxlLZ847/bHfssShAD
S6KRiQQkfL9ijvq4xdy0o1z9J4AZ6Lb58j+SvtuGCmDaz/P9EfNKJTukJXLAoFu9
TTXZMPAmU/pm/3cXVGwZZcPODzi68B6whenT1z9NBaFvzQaxuhKaBY8K8XyBxji0
i6VO7sc2WDWyhQpElAmCcQmz6FEAebkq+K46Pf9IDU8zmqgQVt3fiDviSB17shKl
Bgj2jw4b1exZHiorh1UrACU45ytbBb1KNgdgqKPAJtHAG55icidCRnQltgsAqH+4
+jERK0ISb3/9BxsrMI6+pBsezcMimEyS2QJM+yA9cVbtO21/tUdlebUsAo4WDR10
kkbFFo7HvtUpL9eB/19BlIceIANKdN9K1kLxxdWyY2ITsZr5b66d+SJXwO5lJvuJ
IIKB8SN+6WPXJIMSy/BXKQ+k08ZmyLEB4Dxfjnu9G8hQzoqJhUwoDexRYjOeu4y0
dMYU7NuwZmCArIiLczXNh/IlxhOhr37FX6KgYRy1KHdKkpKz31KCzdOgJYwALQhT
nVZmpPsLaHfZuYJW6V5e0lE0p2x7TPsh9lcWZHd4A8IRFxbzWwUKLo2eVwYak2aS
9Pul9p10oqP9QeRf5al+Jh9uUFjl0ytll897pMJpYHt2Zh9pJ9eZQ/xCiBfutWtj
BUwktmtaoIqSuk79oja+ltB1ld/Z1xelFyizkKtqSkb7QGN4kTyBVztgfRctU0Pi
p8arf9jB9Q0B/82e8fb8+zSW6lzIpzJp+yYysbNtXtILfTvX6P1eyq5fn2iBH+l5
d4qqhBJkt3oqA/YDJWmqi3s/K74YMun5s2lYvXOgHsPuv5mrkMKl7dRbnz0yUYdK
AatErG9cgqvIwx954n7WyyGVmw66N6A83rcjOlbfQLKx01EfL5n1/qK1yRugln4i
F3fqOKzm/C5Tbn7AAzyum4MUHTQH1+gQUcXmkCEWixRfa99veKyzhdxVNNMlon41
/HLH+o0FF99PvZDBbalBIn0UB57x0zyg0gov3oKgUJFc1m8uzKVdmEJxxf/4Sntp
eEX6EF0Ynim9Nqmi+igE2Qe65N+3ZMgJkriKhYKdjODESPxyshDiJrShQBdcErQ/
QwenevX0pAc5Dr2l4CgUlRW711HD697jeYJbR4ZrzKSZX2LGQPhUTTyFnaWM1+AP
tFYCORrajRNa4U3zdIx8gfaVGB2ozzkgHQePT1fxTM8WABEdMb+Lmik1S1Wq41gp
vN8xhrWyRSjtrjLDOQAyP0KJavP+5G9nokrKhowdkIo8K0sVrxuPLAo5KX5gEhOm
ArSo8liWjFW5P+GLJsQeGD7qrCFZqm02gsJDtCmQRHYWsf2hXeYrNHwspeAgP8DP
X/D1N8IGYbzgiBIogACnERxJZ2gQcPNr3gPSqb2uby6IcCCDKW5oebfK8f52Zaav
smUa2o1NWVjfW8ac5s7pIbQtDo1vXEYohL269pOaQMEb5CQYa9mpxVExxXiagn4L
WeURjMk0VTpuRKBepQIampJxWQ2q1vCqxZLGZUv6qkiptRzBbty58n/eUplh+KtP
yflqdmTDDHbLMb3ANPFnWrCzAnfnECDpuAZKlpeNe2NvhJXfy+Jj86FkExu0drFF
RB1jZnSQzzyMMnATUL2O4HRWmTWck7VxjOsSpYW8HQCiF5R0CNkvUDTrXy/bdugn
ITcp191pOJpUskZY/lo/fjcU2DzAUI8qqKGhWe3FEOdOCKPQWYPqKNOsbxleF0Dc
DIQ1VZ4pIABMJvQDPlACbHAjHfP9mXUgZiH4/HBdysOqmzPAopH2+PVSxMjlggGn
u9akb6ePzVBv75fKkuZeX9CpOjPzahLOCCTRruUSa2HWMq4wzK927TBNmC1fD1jH
7DgBvDD0oM18mEDUp9DZsOubLBI3OfJDUIGfehfaw5d/i/RYidBiQGxEcKxr1/NX
mA5YROXr7Li0OmuC7oDVOFw48lYsi2YoCIxv1D98GQQTu5JPTVQaOpmFY2R+pmcf
dvHdI7DaeA4lNmUuT/uxCddElQzcAtdc5X+oUtuGHvHu1/S0W0WOHij/pkMWsPPT
VCjEZwNVKRQJWCk5rzs5Icw1g+EGH9+7ammP+sFsN+hNX50q3TsYqcZGPScinf7L
g3toSABLc6OgDBWHFSK5eE62bMQrqhvNEiN+c5y+W1DmwUY98CsKY2ZosNx1EPyM
fyGRCFTnB6Gax9TXSwM+uUoxYs+p3UdUeq1bDtsc1Rb4pVt9xsZy0ByS8Hep5/Y0
+BmZlmUt1ai9D2B+Reas1eL1XlLbOlebvuINKssOYolGpbymibWqQR4HInQstJQh
AWiEPaOlt2Yt5SAGbQUI1qKpaFoxOMA9TqG2DMdGzYgwU8sn2NlghKqqC+o8OpAL
FOlTSzJcGHA4uqMo0eUiTpbZJ+tFqvvOxwFpPNk8pvgJ5pjPAundTLjuK294X4x0
Y8bE8pMn46EIA7+yqmtBsTR2Cwm15wXjNCshdLmGZqREpJbn40fQSRke68bWLmvX
aO4Lk+Znk5jxWD+Gt7BAQ06wFLvLR8ecZ7P4mPRPDxZw078rLNt+blw4eHm7aMD/
pXCvstS7R6HuLCde8m8YTaKfT7pHokMLEyPAdfyjyPsZcKMSL3kjaLAwj4jSyKVX
hlXJjrPvCiZzgAr2YIbGOqtlnRWXMgK46HrAC+XwPx+Bk4maKdYYZ6TQf50EQMv3
mP5juSKYLbbuG3jDlldL2jxLE730RAypRsKPxsH1rR2GNxW20O/XU72kASwwniKO
gccZS1XbMCHfIIff7gjqXUASudXMAYxAVZsO9GjAurBc/D8Vd780Jx0lvCzHqKGP
yyRcGjDW3kVuYwEOXKphjNzayeA6FTanVFmx3ojS3Mk8S8NyT5r53aG7vAjlD1Ah
QURXcu3VS45lFc+g6+iRi1DpD3vB6LMJPZ4Hy1DlIt0aJqijC2Zww4ikpc6YXJT/
rpw83thWVbNUqQxYPBXUVzIqgvqAoN0IosmGiZ/9E5qnehhhg4SLqhCZWKjyzwlE
2SwkC6wOtux9KYUMYHHOA6AklNIAOAlVFxygtXBmHtcyO9/VvNouO1w1l+Oap73H
p1jZLUCCjfe2uvzIdyaaS+qZcIi8lGomnn7xm2oYt2SheC4cahe3yV1p7qhZR//C
BExnLcXEF7JeDAtJ+spsUXwGnEZNwi8M46TGByeEEyIdPjrLNELTBgbpX9a0+a9E
IzvrMvgRo9CX4crGf7VKaXuO9cNEa3hCGDFgwotm55kh6d7w0B8R0aO7d9Qul5Ly
EoAkB5LEtEVICfU74cwV9fiKB4w16n+IqqMsVWMZ6PBxL+r2BaDtKoBxLKSerWis
6qEk3e3IEqLrsTtvwluX2FA8eZFYwOi8Tiwgymfu+9UrNiFIJQNMu6cdNGwnpR93
jg5Br6mXHqhX1gnqBzKeCXBuP3aCDbpZtGmaU4KwwddbxfxNO5ABALzKdiWs92H1
I3+cnBSE9FcacnXK8+r2VCVOGHwjKuNvmGvTFtbHyfTqXYG9XALmSSm4bqygCEPF
iE2O1kAgc3tn5H844nXxtE1NxCgSDT1TQ11qlMqZEUSDG6QOg0T+EixBMCFY6Kfi
WsZQpoTR5K+jwpAv9qs/p4LNmuHJd0yrGYRljJ4KVUv2HZnZu/8ZsXu4tZFMZt/P
h4Thg/OOAqoMv6Co78XRxe/d/FxRcTKkeqTGlSstW9CiPgJwXAojKEKACOK5d8s+
4tNIf0qnnd7ep8iMkAEqH3NvdQdacgGGrl1ru68WlQEOhD5QQF/3Ie3tgAo6P6Xh
eQhfc2/R29yGVCggi9lpnWHtaKMZBNodIBg8yAjvNndRY8uGj4ViPG0qTed+qfrj
kskfy0K1XZQckbYpMtlzVpDm3Veuj0W809Unzo89HIAi8xzdwJz4jIjqURiXAc9/
rxX/Nr7qUbf0p7oIEwgm0ySXokWHZckSKRpfgQdphNUVg9vghp01qwS1EgfmmGYZ
mrQZ98J5DilmA4fj3jV7qvzjQ52jCxD4hsR5WtIJWCdrUdXRk+nGTsb672eAslyo
qz4yryxZ3NxWiEmRrjzdm2cVckvR6wM6WzwEHVJijxEiaGQW1SNWljI8Za7cvc3K
1OQV1FtGiKYq5qBjboQmD9CwFU2vjEt8mv0FxLHQQi6EixEOQDAHMpxxYMgGA76R
9pcgLvqmrObBlM56I2nlW0ArkJNjFspnZQFsZbv8c4mvYXdLePP7t8xNmCRWV9b7
cHZ1iG6193A2IoOv6Wr+OO1RBXrd7NII6VG8vcMaIDJd801NqAYAxqEBO7ss8pvn
0uf4rm8fl411IfpJBoacg1rQ+hLZGP39uy5pY0wnp6xL4ZfgyfIPzT5fT6DYuXXk
pGWceau9xdxsSILxRvddXx8x1v497cwPwb6H5pezdfp66tsjyxKddKbHGjEECzFL
lIOxBNRJBkm7Hv4Jp5SQKMpSrIDQbwJSZyFEskd+Zro3+6KNMsz4NztrLgnD0Eg8
neoXspmH2tNnv1RGzaB9JrtmOZExlmIdRzuEXQSeCkEfVYAenKvur4Cds4L+6sh8
Hh6rDtaQa32wxlZHr3CmhXZ/niB6biXWlQeLhqHU84X04LAYHPbCdKNeNKeZ+mws
n+QsEc/A2txh4wzCnmq66SMMT4msLJ9yO4PCatbe3Y1Cb8VPi2ykikEArdh6VEx5
dh9rNOjo8AjasYumjjdQ0EuEm1WOEMa8NpWHGdw4J4wnDoJw3qvF+bFeoiB7fE3+
zlDWv3QnJEkpNgQOg9zqjOa+9K129m9bKp7E6dPP44qz4r/lvBcGWz5WCta4n+rH
Grq6JCYUv0rZat/sSwWZDOYZDjr/+/uc6mT+UBE6Hxn7ZRzzCb76S8JXgtaHTWqc
OOSO4+o+/vZ8o+BKMTPp0ngfaFRJYZgjcAhvTh8zYxRxD5HhZOVAgxmBawD40Ofo
6yDth4tKaeigPUalMInR8nupXejYwztEVm/ycg1IfohwRn5vhA9gLnZxvBCz7YNx
zVkZopLl7stX7DL3ohrnLQT/p3fWYfsc8fY+hlgb+2ESu1jNy7F8C4IRVT5V+awp
zKNV0u31YhiCFISRWi0t4glVuwaA3DdaqgNpQPhDwITN7MU990593n6QBaGjnTGW
dLs1W9y6vZL2dKbWcSO7mGy31KjEkc4tshlmK6FRMl9+3QvrduYoc4os0BroMMcJ
ZWX9MYARWm9oOZKfIeBFv3o9bEGVK762qQCNLYJSGUfiN91tyL+ehoepXu7sAAmP
MaVF+cD3xmpF7CGCCIJVowCv9TLuK9AsqI7yGzcIpAGG39WqFJbgZNcqI3BZFP2v
XzTF8QJICpEyQEfJrLsH7fIfYLC66Qw+6m1wRuqQIYz+4CghwQDTPlnJemAz+Pao
kjq7GFkQshpRtWW0MFhs3dxatkru5j057rnbxEGsAdEDFqjp3wKZStNtOznRDyUx
1YVbO8qLpS+SZ3cUnV4mgkD2whNIDWSiTwvKCJgbvmtHs46F3d2TyOavJf1ljrPl
IQiwW/kDGFpi4j60W2vnbsJq22lxMZ021A6YXJPYGHy2lMjWWqfT6txuLenLBpDJ
ztLXx8RAKTnQxTGNYVYvoGq5NtspkSoPu+ZXIcivHy5RKT1wjuzeI2jiBJKT3IsM
7bTdG0n4ybhEQH7Djnzej+V1JLrpHgo0NJ9Ga8FPEQ4tSIghXsPS/gVPf2e8nVF7
D5bZQ9wDgBy9RLaa/KL5bi00a80vUlFHJN00rvjBWYRtI77I8AAktmYjlvUQyfZL
vKgMpIMbdfO/v99kw9JgZHCtFu+U9Z8UVrB/18l0EDnP+AY9Y7nHRIgHMBDZXTX2
cVfUdLNKRXXL5PF7KRR3cG8ytNieNRN/hUIADFfXDB+jSnPHiE0tjEw1APRWI35G
axvMSJ0YK/9UEKqH/cu8Cjeofh11bkTw4Ppgkx0xdoE3FFaQVgOemdYtnArcu9t+
ylFnX1pBRFN5+tqOwjV6BzMbIcahPEvUWvefp0RNeSAUifKLhP+eR496DDDdM1fN
4IiCdV2d4w9EA+rjxcVHNWOaBu6vcBFCy3RLtEskM9S727EAt61D3n4OY6IiF4tz
S2yR0tPv0SRq+UmaAQE/EtwBETKZjPg9LoTVOre+IH1wmpjPZtz7XnNriyAExFGJ
dxuf4PdgQ9PhVx8frQqnPTnm4Tv9XuEejUBqxE0zSha3f/NL8hgSAjs2YMuBpSzq
Tlv/zvlawuyFf5PueRCvITAvR1wX2lknPrRsVIol21feJCNtY/i3VGeMKqZbYuF4
zRJkXCI6+NKxkW1L1I09YeSfsrKZtRRGl9zA7scUkcAAdpu4k47QMMklwYvcoW59
F8uSfInCO4f1GXHm8Rjy1+Ydg07PIAOd+qVMSYacMmAKgaeDgOkFvdCX3Mp77NWD
TFYyBlhWrWpSbVIqe4Gpw6+YlG2Qn3zP4crdtJQt8uJY1nhA76YdAffR7f/Av3jP
tpvhzJfVDYL+fBUU8rzucp9G57mv0NM6KuQItxhdXnuQpy6jsOBxY3EdMYkW65sx
cyL30wy3rDh8XkG2s+N/QrSlA1fBpWMPpE2u4ObMZmkpgpAbsDgVRTNHaaRkQyuN
ftKGFbBab6jSsc9FSFEsveJSYbDTihA3VXAy/FJrJSJ20iikZFVl8qfmPn36BXAg
peoerNMROG4ZYQgiQVzmUeYnyKJNMy/4KQiQxi+Ye15z+Vjjs7UMSJ4WqBTH+fu2
ZAqkVIY0qJC4flvnEsRp5sHkKudyrddCymFQ0FIa1fGFDWp9xWvuOYc9gsujybDt
XhHApzasqArpom0ZrQja0HQ9wlBTVgjtc930qmmqkj1UjocAiPfU+6veonuqLetd
CJU5aNCqErqz1Lf04e/zpvJWLLj0EIIyenlJbb1fYYfpf+kgHFl98FXNfj+LW9l3
Orn0fcGPQUKnCpgSHnFibut0flEIKMvvfF6aedhqvr3S49xzCaMsOlloW5VdR0WJ
i/h6koG3Qgs/e+k8SauwQS8c13POsPTQIkt49k0ffux9A4D2DA2RAAk+TQpftD5v
qV1cAN8yEtpQgKoVln67iEWfNGkzESAJlG52IHfJII3sdbyRZ0c57huridzEZ6po
shhLc/XgsrTqeGT12+nGsK8OalTHdrUEyLGE+FodNbfUVgRSJk8gY7wY+NyDZfzz
/8yiimKtuz+hEQos5V/v61bFAGM0uRbsdLIGMgrXG9qDPOBGXzaK2rKiO00FKGGx
hnXSmGVZGSUnrDm7/k1PvKTsjugKE00or1urk8dP4OJ+04fhMplZ2br58EtkA2o1
BdzAM6+SIPC8M3FJMuIP9HGLh1e7TWU7BmC+9jB6RJ5oSDn/1b16IBB9CQQhqVG8
XpwUWT5FEP5jvsnlNuM34kSk55WVe9U72cixfS5pGVZJ15SxJZ9b9WsPdmM1IJ2w
jciy7R5qh/hFbtT3bbbw3ijIJ2AwKAkIhhYCN8mmXDWhZvSaiu1D4jtKWGyQlDh6
cTgQkXuVADuw7s7lEKul4BnsdTvZzPc/wXbq2nYggBWzrao+vQ+gc05++kr7LIaM
n4ERb44pn9cr6e8nzj51M5Ra2aJ4JRErRTpDZJlmtDaVsmEoreU+ywndecLyA5L4
E1mdpNDxd/d2fGSgmV1DWXT17CMpAN/4zDIwlhSjp0xSQbgQEDQJWK4FWz1eyAAa
9iHzqmtU6bIKOlo4uRlavZnwcf2qh3w19ltH0PCalrNF0vUsraMVQGnP3ILnYPaX
r++cRSi0axNE+nI8/cAnd3xdorLa3ZGYDK/vFF8mLTdJbKLJfHgcs4wyhnYkOIGP
F7H0bFjt1oiuc4hlubnBcY9C5IJMQrBMatLpTT0x9hAUh/RmYzkDGEFP44w8jmwG
gCvUAZQLLlruLnRpkxQNypdXAEwLDUvkh3A/Iij7xPgwJirRXdHykSkjGAk2hjEB
BuwERGhdExkkRtux5+6ihiVxJkI35cQtN9cQVbhNn3AQL1zlKDnj6vfNAFspEmYC
zJVj9UGoo5GXj2MGUaUl/MZFjk6CwktJjmcFjYMy3JYnJAggBD1T19eYXLHgDzYx
B0J2A8N4yhoudBI738XfRPo5w1p3hEoSSjY3b/oYvflS4TX3pq1mKhOIJbIZ2vu2
NurjXW2PPmtYksi11K3zKOmLjBKaDnwjL/kkTnfoDN8avOREhxOGglg8Oby7aUEN
ACZREcx1jRmF8JwPUiTMPaWY00NTRlPbklXYXnVFSrQUbAPV4g11bFvE+lxHqAE0
21CqFvHv5JHPsh70IBw+0pjz2LgHEQl1S6ZDYipuTIetHlyrjjCq84G0868rsnMx
vMl8r/b9W7uORhuwJzNvmO6M3JmMOt7y1nTIfbnf3cVXqx5kLHGx93HS+KtqIjEw
cW7FiRBcZqJfebeR2NFuRcYfoOeDLv9GtrRjmGlq4f5floz9ywN6+jjP5nK1vxWl
K8brdT4bokfcb60Xdy5Ff1z8KAD1dJ0BSWbJlglIIbd/N/VaMbjz+I2N9BAcSebb
aTAPcnRkAWkmALRCu4SzVcfD1wVhWIRv9DXLBKpkds6pXHSOVP8AGQaDB0c0OwSz
krravZzjAWTs74zg0eJfJrKk6YVpZwpzYkju2uS/MpfXFsFfwrERP8JORQkjL3v+
qLu3/He82o+iiYJvXBU8/+Z3GakYfvRTJhBiE1mV2YCVn3ZnbZ1B/SvGxJB1kOwO
363q5U/RRwmkvXe9a4B0Km+k9RL9Nd5Qzp5hi+xtsIgbaCLle1IQw/c+WYxJY4au
nEBnNu+bc/tO3Fv8/p/QH+9zz6dQVk+T/GhFFhKtwghE6Q5STKR7OEFmuAE7M/3Y
O/yaRPnUdpuTCaluqHYsE0clRBJXXw15dGKD1Y03S04/FQw8MPHe1YKnP8OEY+BH
dHRPCzN6Jmlx2Ce9LODOK3SZrx3cDklGk+ifY+NFYKGIS5uFnwD2RvwcMhZQhy6D
+K/+MdOSpB8Ycx4Gi3QT1KYtLM9P1GFJnib2ZKcYgjLzWGlrS3oKgKBzLG8JnrJC
R/5d1NG4nXB5Pj7G8CcMnXzoRZML3UHkWBiMjkhbsgJgBX6ppRaat4QRoOFkLMDM
xNta/kGSGEbHwT+Ex6XO1959hSHhlhm0GyJEvgws8xz6H4f4ogqngVT9iyuoCE/H
rTdrosLjG91XAs0QI5zPCC3oSmXrMoRo9bkME3aKV1auPIe4cwdLbIDswSE9/2tk
3nlq1waJ4mLXu1Rf1dwlQ1RBuJBNaofgLFKoJ/1XU9lErjtXzKEnOtQy53u02HaT
3/IUo3ru4Vo6Z1GX6ZUUa+Ln1yYGrvFbsQUic00y/fbCH/KT+ZnYsv/hnL1q4/wj
w60ihA9KX3t3/VD/PnTbzBJRZD9HAgsJcx8q0vN+0oE5QhLY2xnm0gAy2iH21eyy
wBg7IOYlM0CUTmbKlgU9tMdAloYLT8F4Tx4VeKtPxHH7B6hSJUhmiVuPUqzczvFX
rnqCGmYsOoVnD9KkxIjntL5uf+UTl3lfXEVzolTp8hi/JQmGXlkUOIAHwNdes2Pb
OF91YxWPRnxO4gGsiJrRegxXaFkoxMIaWe3g6uJzqeInR1Qn/kZ8vsp8vCKNYFTD
j41PCaSR2bbEt9crfk1b3MaS2PD0Y+JAq6KyFdTxunsiinE+4UTOqgtudKTAuWuu
ellsGjolPpPRVv9H16wG1OfKxd2qNyYwEInJ20q3oqZ9kLtKKaz+CezVz45gH+Bs
LaHNmA8hdh8p96xa/YvY9zfGkJoxf7KlkyK3Oa3nzzh/oocZA2sDeXwZdpKx8FS9
J+mdLibFRWO+vyy77oVyqHiyq0IG0TfOdUsK5hkAWSlAlxO8QBZePMCtRErmuIwx
yjNjz3iDOhT4qXQvyBP2i6Y/4A/tp3eNqMBnuAiOxXjxJPCQ7AT9/g1Bat9OU8eH
7O+HloNK1Yczh8GhY5sW8kp9OLWSflxh7GlVEURrwLGmqXY4C5wWCBo5w2m6em0j
i4QBLLUTUdQVpevY+Ws3nvKXmkV8NZadCPEh4yYfPhL8vcpKppUXMPKxJO6aZDNn
TUEb/vqvOU/AREvz3A3NhVso3mag5rzaaW7EUMH9s7Mwpb2Ti6yL0R8+ZkOVW3+z
IZwziWZqERcEv4PAYAEsIDOAdGIhA0vcYEhM7OE2OKk8DNqO4xobzj8KEBmvQwjo
XAQ05+28ws6h1380O1f9ya/1teyoHsNETDBciAKkia4wJKpebn7So8Cvro+WMymJ
2usTK0o/UPgbPoLnINhXElKsm+5dfWYofuZcUsF6f/8VGmQuyLFRet7pB2uR1X40
O4FliFkhTlot5ZtguEBaxjQN6j5apO2hVTRX2b2EdoFebJo+0MumA06WUYVLqH2o
wIXTOKmnQ/mBUUW3IrEBSU4RMLSS92IUQlBxhWyhhqwE/DzYrXABrcmlvRRiCU3K
MzOtzlyBnyOxsrlPjNpxccpd5n177weV6BdFv7/NnQmGK+I2DhJ4uvAI5TkYE6tv
ae8coH+Fm3fonlyHcBJzFwP4uato65KfUxpxoTTIXO7OHN8/d9AgcIf6D6CZamVq
GnUPliM8wv3FX36O99y5aY7P+pL3WC0W44z+oV/wNNSVWFdnrovyLjEDrypLaCPg
A5tGmf1KtgmWRBXk+fdv0IPWr1XA70TdpE7knZQooSla9LEhkcbJPe12Far3v7TD
3IDuKQOfJDfpoAF2Ajs7eBMGqAoNKoRS1sQEn33fK0NIKQb+VcC0FR/urBu6gSxm
YW4OwxrUyH9VAaR5VtiwT/mscftzXwU6FlXoB9QSJ5uD3TDP+WVbx4ncW83Y7EXf
eYxINz/3VgI7aqmnRPLkK+3A5OvHm6Eci+/dPiG3kApbuP9uWDGq4XBk2WEVqHyX
kzH4R6mumIchbcs9xKcUxG+ppcwLvybjE1KS8sxFXx3Fow8/ISqT+hkqaiTiEqLm
E9AAjaZBYDel9jRQxEwKh/zMggMvSdsdlBL8tNLBQYxFzyqH4nN+0ak/lpPoCoXE
a1z3M94dqGp3Mo9YKnkj+w/wk8cY24iHaBOYmJwJ9iv4VRkI/E3bwhAF9BGUlD/5
fbKn3zDDTNthBfYdtA2Crtoy+5uzMhmsovpWSRMW7yeX0PEVTwjnIohzLdRRaYuv
nvLLpYLnlKxqNDbSZPR+AZGJQlvpM56gW7CcP2GHGWYo6ElRBSy+uHHKNGrjacbf
iYGmSLToZQUF9Q7KJKIM850CUAcLzgBgRHId6muAt9dp710dcdte8GbnfB3sXzzP
oHuM+ojaQdoGa7OwT8wa3RTSDNxc8ZZOi7Vquuq53AxDdiTBw03XZDdJv0swggVj
58mLO4x152ln0+Uws6Bn6+RxAXmiSivK86k4FB/jjYqnyEck0DD4IkboyamV5SFh
InZIQdiGitGI35B6/yjdNB225DfAfa79lpWVxjJaUv3XOB7icHLMHF/AAUs+bCqN
f2hlYB7NeLPairFcD8Go43bPzh1Ad3Ihf0f1PAfzrknS1H0sEL9ObxssalJWy9Zz
dX9I+ScMNu9GOmsgwrDXEff9itoxvT64kLqVRtcrfy4KCYCSnKy3pf0P+P3nE0tn
4i2NdmNqB8V86emN6Jk7hUSx7TkuPQL7v2X86Xat2e2KiHlDHQ2tpSAU6mLYKMCJ
6QpeloTisJV+HdRsdeYy14z1VowzbEYfMUcqMxvcxGpYTkjkIZUgh4Jyc21DG769
WVmfuMGFvpxZjSPWSRA+bCKBaEAOZBaqbiu4XESQj9IjB9s7AXpW6uTOQSnIBJfA
WWBNYcuf+olHTMGoPYoWLndKt0xTi3+RtgShqtngJNpH3TFmKPZyASSmYFogMhEk
ePaV29E/sayeX1EApCsfvHOhKkJIebH3N2ZdCdnChc9zG3EELQLNDJUChG5jnp9f
yke4oxQEa6u2xEc1qyVtnclzz29np67DX67s9z1e1w37/bP3biPn0NYshOK1Kz0k
yl6MUYd5oMDtsq1rUhFzN5sRuY9BcMm5/BUMxm1+G0Q85VYaat6M04jLSsEHKH8S
6agrUHqjdpv1hUNjwaHd6+gf8rmYv7zZyWT8Q0rSsayfJROXi/VUbpUnXFksm5ZE
xfTkooZaGe6gnh20bNyZzBb5nnU9Bi/MMnWZCmCHo9JZrgUvJ0RtauQmm51Y9a6h
ODnBE+F7n7tMdAoFPF3VxxxuHXjNVaFM7a1iVinpEzuz4Bl4pmmdh37zba94s/Wp
uZMJJr0U/ciMppMNGwNFfugL06kT/Lu0L/LtLF2F1cbR7cjD+YWlJvzKBUrhaG1Z
uHZtbV8gDpZGgxHp8avDtjpOuJbwgT1YtToiIAwbvdqCRj1uJWvS4+ePyk/FWpHi
sf1Cyge3UCUdhnDsLybwJfpfybguKNb9zOaeV/aItuh4goFfE/p7MO+D57MN/Wqv
iGc+7JvO6GdedacRMB6GLgDzeHjzuwHiPmEdrYQOa1LbYpoQ4gsaiYDB2QTRmaUd
wt3mKzxPVpNwVGBDcJUdTLbSbEycta6/l6WDbyzHsI4Fp0/dZzBxjRZJ+h473q4l
1K5iorH4IKNTEHndn7TaVI5Q/16T17+sA1+Z/h8oJ8jBpgrOz3iCA/0entLtzbdx
jdItuXEZkZvLxxJgoZ7cT/nOGpsvV46k26hOlkrK3UB5LG9o224Qh/TqR/ypmaWk
ObnQ8pxUQtXVvqb+p4wz7VZLu9Xv6wNAnvnOdiuB8HoK2A8sLCw37gjI1OY7lHHp
LF3w1RKs3Ah+s6AhIZg53GqsnGKA608kS17BR8ZyKJcby1KpBxQDtmz/eP1jdtNS
nkPPDBv+Mz5XyCEn7+629B3+qb2Dqz+U5lCkhNM+YaIdCgRAvj/O2KmJWpDSmPOp
lTlTk28LF5wsS8b/DE00IXEJHcT+uqUbuJAiV6N64FCkH4/NdnJKqZKaqGdD25bn
Hrbj0b38aE4yK6ioOXGZEqNSZDPwO0kCLi1DGR4G8iG++gjd6Jw4uF771e/0XTCH
IqZLFMZTjQELhlD8iLRnZFHrR+ibs3208qCyEZSscFqPpDc7BTzFGrDQQ6PrlzMV
t/age6LSu76onIuuE+aHtTZ70Ut8bV+f89ft0BfvsXVu2IrXkY7Tezj7ub82WGOi
46kpQkl8Xjeo8UjIOlrUXN+3CKGBV//mT4xzGFdqvPyFqGPot/bFwQff/CcUWY7x
593rv/+CxDLpL/8DM15HDZ0dTpDfd2baxNPloj3LjHDUfrHPzRXbLbUXw0YVvALm
obOUVSDNZMZxyIwiU1VCOj9dZ+MdIifWNTbPPs/hZaEWRDcDs13m2suGdldFuGow
5fw4DX0bBOrzYCy+/H2I8s9SAzEnQY3qsFRum+eIhSzjISQ3HT/I1KcGJFs3YdA1
uzhO0GmAnjBGUd88J25gNgSosEOrXp2yoD4hOI31GC2vbzMg8ulmZG6tinRmTa+o
4/xCTOmLMXAJpqBmooD9+xfvHdY6eN5YSpcAdmvkWZBr6yJkhqSXRfM51w8g8rif
K9eKkWtnltQA8iQZ7sjpEqsrsAs6THhjXwsJsFkpfe+z5LBwqoXx/HhfSX2OHZVO
hTCsuKO9Xg4srVldS1IUgGaTDQnpdhxbIQWJaCrFjymGJYOo6+hA6cS2Og7+rw5C
6MVoxGDwsJMfRTyVIX5sU36DtmeX09nZQuFgUFfVomJssE2kcUMV7a8WXu1fkDAs
qNYPt2QQLLcBcIbhZnR0pwV3WvWSRwaqe1qBxUVJywf/WBZqBu4kYDGe45F6Y3yp
H7594Dr2jhO99g62OumzOgvZf56/Fu6FNCh0KQERB43p6RHdo03S3l1evkWoYEMg
dR/5l3CIbzJkivooSKGrr0IjDPZg+rm694M3OK4P6sqdSFxsAfpIHraWhNtXPqcx
n7d4H9wULKMC+qxZ8cxvyLej8vd1Zkw0R3i220xGondyrTScwPk+w9FWbiNLGRjc
Q3QQNJXsMK38CYTjJl0AVVos82Reh2EAgj1wps8b2c8Yyqhr8dh3pIfFq1VJ0dPg
pNnxdQ9bygePdLCiUO+IlqJV1doiNu2Y+nwHU7QnAlHPt54xHdHoeqrHGaHYufQX
Kjyd/l+3CU0ysIuarYj9g0iGuCF/zDn01xKmyUmScLtHxHdZms2JsZBviFMV/CkD
EqFVesVIKxHwHCucOQkYKIRvQUNchaibM+Q0WpRkCzL3h4JhyzbgOrR6ySLu2F2z
BwlM/PMGaRCz/PKCMt/2wsrNI/6Vwx6udhOcs+19GAFzSwFOku9pPiHTGdHhWcCf
d11CzV/rQhggod3zUa8JbeTbrH2VGs4ydhEP9IW9NlMmu26chvUniaWKNHkeYvEH
bIp+EELu3EcG2o67fn8chsfjHAf9dFHCf8bI/eDO82qmVsjwrG5AmX07fbKWRsFP
sJRT7M/Y/Up0SYtiFQsDMF+fpnmxn1Hv/7G6pJDJ6yG0kErhXLR5RNN46EvcnFT2
huSnwLDp3LLx5US2Hp+sqHbr+jzP6flZAtJpkt4tOKO+wPFKBvWK4QvoglCc6b5C
fGvZxkO9tBUKk1B40FdAxWxzxAXx7HLcPXRNJWXdb6/NZ+ch4wJWS+A9BCto7w3O
YiX15t/2NDtbrYGqs6+yps+FgiQCby1mBOrMCZbMpfAuiFl2VRZ3uzWL/alyq2/9
dYirqTiR+uC9tyCB7t+NRKQLMea7Y8JxFVJy+tr6TG45/3lK373BVsymAGhfazMk
wQ765CLP0/V5yCxoZCg5Wg2if7JHvdMGWg5gmqAR5NCxs6dKpXOZ4DopAlMrBlPU
2Xaeg5J2M9vkXLTGMj4NQEgSBJ2POdvGgQ2ucYeJXIa9lO2J65okXg+PNMftST6y
52AauycgRuCiozEBzwQ4qpD27p0PMYOPgWM/SAGAY5lP765v9KN+J771SRBo8A37
Zhj5Qq/aznyK9jUFcEueIWT+4B4SPeSAIpEch5QcGWdnnY+5Nt6itGN8NTqG4pm1
iYHqhmLMeGJS+4QzmLTKK9qKu2hEt3XPDBRc9/jezNX6l2NWg2dbJ2G0kjjbSfqO
liFhi0C/q1lUe8Us1A3oNBaN+cLFkRpwHeHn/yASOYnnZr1nf2pNKyukXhmNLa8H
/EBrC+rmhzrjWm272tc6MbSQ/rzPjOf/Itp/K3VclYtDF/yXA8Dh0oX1GMbYMdpp
O2B78nI5mESrCTxs4jxiXq2bvfDUi82vg91ggC0kt2xi8HbasV9aHj6xGHxIkxK1
+3xsUiKdKgkEx3kRUtvaCHTv5h6jWjzZelRMfU2nd/myGaicMxa3OIvdX4M+HPAF
gPGKb0b+3z6m6sW/cq+K4ownG8a+v3tptPEHQWGrr1t0W9UMVjxS74DysmurI8p9
G9vWW3Wc8lFBpA03dHEQzwrdhP+UjOTnidFSqlT2zgpHR1ocHyHve67UGTTuKExB
arGReF5IwreFlNpYJ/f2EUSRTjdpn1h6gWHfcmJKUYd8oqPnAhc8bqoR9ffsjqIQ
2BaMnwOwQNDexa88QCaoCrBOzedqrmHNhCc7wixi9wfe3Z8itZBDsiPkwUtjocyo
XLh+k4+BSLiVoW3vQnKjP9xbLDzGJDW4pvDEcO6vXbcMwvs8xRU8VXGra4UtPBLo
4k4bSBZh19AkcO6W928msALoBD5JpJSBWTPCEPJTOG5gy6hxPQN4zqZ8WpEO1UQi
Ayfn2VAAhEX+Os9shvskQnII08E7sDuzPDMy7K3rwnU2cwtpK1/XAcDmL724z2rT
zSJm+HmE5O17vkyBE63fi4Aiq3hQYujIepbBQZVemxaGClIh8t/b1gfwibP7/O6d
eb4GMVGCB4SZMaiT83gOFTzqdvhkIQwXCu099ETlwjj25hSUIaoX+kJOwF0Z1vYe
c7Kk+lJiiEhucv0n0aR+vejRq767j9iP8mdJ2P0NdAO65IqHcDa36SQfX/s2SKns
tNslg/4zSHGV7qF/ekSPwJ1tVRWhdK8MAfZ4eNQLBzgB4aIqHnIE/rWPU1jLaVyx
g6r83QBBjzgcHJLKtewHt1U3KL7queHT50tLVq0M8mkvw+nQwEyfPnVQm7aACm5C
By3vc9XjxULNMrZX1NO5qH9xShTH3Kmx1kQpf8v9vmhwq2qt7rRgHxPSGR/Ln2Wd
jDkQYcXUqDvKagAhpi6YF/5Lx9ZVrBadRaNKw/kWfquTNvBxhWeccvZ4csKlP9aj
0PGj32koiXxkdUwGf7DRSxsQMA6rzqBOywqPYkarPZ7bwosUbiVM0TDn9xy+YwSt
37Fc9CmewzZdU6SKhYhuGRgqe268+TOpN18OU7wx4BwIGZIjJlt8qHxuOVEdbOyc
E/wWNA4U1I/XJOI9Jo+tTdc7QfciNk4hd2/Puy3AqQip84cufF0BBRwC5d+q+X3a
7lL2GTu5XBEpUR1FPdkLPSmULLo5zwGTCGzF7djyFbYGQ1BqZysY6D7TqlcKtWfs
V3W1SOCG83keBzDt0ST+86PyIAh62Ji+12E8Or4jD2hoj3SKhxrFW7P1wmmRpDYM
YVunheV8XAyJBL6A7aszVk4pHLQQXqLEmQwhR7HuRreq4R2y0NScXirakcfGW1bp
KkflnYu9FKKtECnf/2cgLamo5MSHhjIRl6WkMZjO+jTdLGbBNnPFezKeZ/6ItIm0
oV4llWJVudOp+fOVSllw0L/4DzXxaq+OYEwZzI2TYaHob/ZAWfFXbbVIJILJY41M
OXqEVo5QVmNBTCmzcLlhIdz72Cx3Cp+zw9UWwv3hItAIaSK/5I2DvJhGGWQmvXSm
49iMWQaCPrUr4jHaZPEA97nooMDPdpnh9765EzGQ2MU6ulxGlckDl8hEJYd2+9Zb
8CXomnr7OgmQ83izmcWncEvrXseM4d4N9IrpPTrCvScq6zBkRyHtF6tol848Iksr
pi3r1+DLkqt//5X7t2SDjEUWPTpGy5MM/CUqkODfStrEz/tEZ7U9v9KKiz6wUjTJ
Lao7p/T5PXu4yuj+HKNxRx+TbUVu3F8RcyIfhGF5Jp9Fj0IxJN5bdy4ppTxjpBbl
esWQhCZ+9vby3cXnJii8Ya06NvxTPbqBfavVk/5C+fBvmd0H3AOHXMq01mnTTDrN
BRagqTAN6oE0Ig86jlvTfutWQpaerce7dIK+v8QmQf0fcqhdnTKhRbiz6hjuBoRr
fuMWzovlbQfOlTC7/me5nSsOwwCD0gneXq6EhA5Czp6mCLy+0aFGIPyN97pLyOKI
mtYqzsWCco7gh5/ByMgSYy1qrE+xWD7j91FfsMPkKugbpMV7nwvnMtSbT4uJRlTL
NLHjryt2W/NGyMwgs/eUtDOgeiXS5yabSrT5UJXhC6vsn+7FLoY3WIdd/yTqRnbq
jz8xFDphKgwM9BOFT5e8vOBitxtaTtONC5eKusIuzWZEGSpVVwNVYT9Ilvzrl+XD
Y0oFT0qxbz5wF3iAskBRm7ZvreNmiyf9KiFxDIh3yhaNU32OCJNQRV0JVsg4yJkT
3y0xpV+RPGIt/1vZVms+lalqfdZb+67geYbmLfbqQKM1/RxMBb7cbwANsjKtP0Tk
IFLnRByqqjaR2cNgC2g/ViDdeKYv8GbQ/wzuOJXuc8OUG9bYz8t0Xi+HQTpBOu2t
PRocK4jfIkG2MCU13uIv30d/oikKL0AhVl3ZmK+jzKipZFOtlFmo66tf88tenf9Z
LpJytDO8EsGxkHNXrQlZ79Mx4tojlsndJVkJPg+G0kLqbiAlAIAm8xYrE5N+YHED
oMsQ3NxWeYy9HqMcE30JblkHKr10xlWe4O2KYGF/nDQJlhqX3HmbnlDhZug2Jo0a
fmDqyGSQOoszza/TbBcbdhgE+AsrC6hDgS1X8MURM0FZfYcZ5v3qr/96z3nZUj3t
7zfEzGqtMrvAp8ME+MAZ0WpAvNrJIl7mEUwyAz7FbVKsLEatHaRZbnVac8JkGI+K
iCx98GeNuvDUjC/IJrmm1Mqi/B5F08+fxIQZ7i7S36f3sKkIRcdtFT02w327g/Pd
iPWP2yVj1AMYcSffh1DBAktkDvod3GAFkOtw+ubz+9Twd/EXDDcThvGHwKjKtQwz
gPd79HtkSLjCcvPoWS45pHfHwUf4X3vi8Hma3UwMRfpKqyCVIZnPZAiTt3846R4y
brgyPbm0ClJxzZdtYgXIfEHyCBGvom+nSV4YS4NmodCv/aM6g581zFvYGNA+TsAN
HBs20vmzzy5PvteJnn0Px62wDRpx6QsKzyiYRMw0Vz45WuLzrJV1eDGXhkRSYym0
umD5D9Er8pFR3JAtJ6JF5rkWrnlJhqcrvW3MX7gpFHKococ3vHi8U2naQPDHbaod
Y90vXRn9iHUPnBIeYWSrnj/8QjX6/N4C9Pw+xP7d5ChKwTK4BqKMpBL2IP2X8miD
U4Jirmzia3/JllU5wMjoHL0mbTXN8gS5C5Fuue+ehE4mEIqMmJ+SkrVdIPBvCUzn
3S5RG8BdFzZtnLxBJrYeuAPLFz6iNQm7fPkUAvUjj2pWg8uzIjLABSyhbWv8i8f0
AGNK4RJ4JPcYNoM7C3MV/B5iluj0KN8o+7SxQ3Epb5a4HmZDV/f1xUehkMFio6CI
JJWzGSMep7R5Xk2dx2+YjiO/AmnueVquY6GabQPEWR+ii38F7iRrw/aW38JxQaIe
mC7KDS6hRbpTtFreIWOMYR5mv7PGdLZsHskifK39K+AG1p7boUBnTXX7H4/wFnx0
7uCKlLda1pivUCNfPHnCKPAaUWhU3PtMWTEVmybWVVD8SDeNZozcymW88zHeX611
Hs1d2OBQsrojrMBMZi50faVEh39w/rXo6eyJ5oMsv3Y4iRKJy7oGm2uyEmOYxNRi
3m6p068wFK5O6eFTqeqR1sX33nueNuwTM8Hlz5iuxgTEjBlUXsGC7ZCe42/8fFf3
ItHxeD6fS95tJ2IrrqUKYRfIZdWcAZ28YIrd7hiVkUbSEbNM5OKkHP5N6uTOIN7V
b6btOgF5D6L+UGgnZGTvfoGy2KT9DnZ+04YBzU1eg3it6DjxLWdCEcKnc/E6VN8v
zMwCauU1SAG1GYyjD1Wpc+X7ylU/JJaOZ6/l2wss2Uy4dmqR0coxImmiQWk5aP0i
8mzqCsGerG9yG+K+77JQVOSRHhNhgRZY8H9ikmCr9UWpltOoKc7VcSJ2UDHgD5/0
v1pZCHTl+lZpsmmueOp5Y7IGGGge2REzTIkzHuxypnlixOR4l0DLRwNhCQZwEyCl
KcyLZDtXhmbdAYap2t2b1ECodefkazbMEifEQdocnGlnj/aQLlISk0IuC1XH8SVE
YnmNRH5JvLAoL324YJEenx5IVwQ1hEJ9a105s4MX9GMdrJTsCzAtrY/bacsLsK4l
zdYmpswkc/CCLuY6z5FtroiG1AzkgYyobMmeJ/7XtZf55qY7pj0AMdx7qir1HILO
2K7caaqhc+qzBXN0iN/rj2Du9KeyQzCEALOwBOVPUAmQydEa0FF4jsMGJ4hhcXAU
e2wvP/v6JFefu2ApbhJHosjSHWlq17nKYFRtVm88ypMf2Y9GkuJvF7K/L7/4hrOx
yIsnyyakNOesXIC/hQt/4ir454RVBObToNnx1Vv5jef4MeJKPerORtIwAnR+uNw3
1zHBZ3wVrK6yMcbopAwoLkuHCyg4/9bTx5RAaJZIq5r8YwkuCMZN0RcZax7loG3p
PITj8PVxDnr2ybSPGbBsjJN3GkQ+e6nHBAAs8fKMyLbUmyVNuVE3gjcwhgoPxjfK
DEUoriPnVQRgZ3ANa2jLlSosIOle+04pZNcOoOefO17Iew6OVL2bYYj+F7cPWtAI
RUFFWEoMoVldRYtjKZ9uq5zdhcRj3xAno+tpJf8gtl9mr6EF2gdRB9QwTRtavzxw
PmQ4q5ALgEi3UMnG/hvcoA23M12Bc5M2M7NEMvZ9BffbJ7t5esloR7KD9cdK3xyq
h4sgqJ3Tjw8YcHpeY+jyXMK/Kf89XgrdkvMBtXwPmLTn2rRBnYWli4XQrZm1Qo7a
redPvHM65tLPrJxezMLm/UmWL+0mcnTEp55OhUP7AjSmID4flRgSSUvoknXyN6cb
5Z4HUNJU7pG7QeaLtm/eU2EBnxCO5sUEKY+DAjVp1XGs7Q9ROOLZI2QyuRllWifi
S94XIF3bcJb53gI83WEsV1urraJM0WjZ0s26yuIH9cben6Dq/qju8nKF+a2Fnl4W
p09l9l7G9BvP8lZCFi5o8KOsr/JeOeUMqu1CmotiGwBCwe0bcIpHCNwrYzyOPh3k
dblbnDO47K3lLVM9FPwMDw5L1Yk9MG2yXt1LdPAKZbKN6kLcCo2qn9y0RRnIOv0N
MORu/Zo+nw+feSZ2Fy/fJ2uOC/xsrY5Fkn9Z2PROm8thKYX3XKc8J16d//dMgW4z
KRWqEXvz+6BoTK3BFLjmj74Of/jVibbjNBgZ3DEH1jMFlUJ0lMfiKM/83P5kDmCD
E1XxlngnXB8N/l9o4USJHEDm7Y1ebe0WgCRCuvupEYvObkYD6IvkBXlWlwYtnpFl
ub0/hzlFwNublrOItZu7YNQ94t8abNBLLiDn5AhPp3EzV34dzBOBg/a41W1Bdi9e
3QsIaBFTFclqo++Ns1DvQE0x0Znb25Nd8hnS9XP43MzhqRJMoblT3Tl7MvfT74Z2
Sifungx8TUmtm6+wSMollxzEI08DyC6/SXL+I4VNPapx1akTDCk/jUqTF6tdxVs8
S5QzsHVNJ+J+1Wex8tQGFSXjyfLyBSXqhBn8sfXJ1gtJG2jTOqaD1PnpziZXh6pC
6b6o6s4xZDdCR/KuD5z4uFnNKeQ+n/wgF1Ta2NKT6rUggDXXYl+vqxX0YUVI/NI2
Z/lfGl5LZr/tk6C7LdbVBTWWWfnFbllZsYXcNVbe99louK9nhgPU3zn0VsnFJHCL
a93pFBNCiTI0fUqM490uC5vJCfLTcfnG1+MtkBoVuZ/db6W0y/RK6RGRi/BfRPIw
sv4YE6UnsPPrZaX6bdAYejCF18811KaxkkLU/XCv4RCt4Fhd2M185SYeXzIWJywt
JNAV5OZwZbojT8iK3hoelagkxKv8u3ee58Auh+jexGMyOvyaFI5PsFNTXVla1tev
YhtdNIOKRbFJMSyukrLdZLq18jrpXjES3TdZQhrXw1v2EV6FpncJqU+V+x3rFoiG
N5X1uwHBEFniTPevMHv1gGkW8vkdzF2ARdMmaN/CjQZgqDv6geam51Rn5NJLDp1j
z0FaGZ0aPoFw0TNIPI8GJXB1MRU9wQ6TfiBm47Nyx2afJQdI9fXRqDE7fHS4t5wQ
xwbN1WWyGz0wiLahiJ33cxBFrVxvfyHz6sEOvxyRVywE6viUaBrJoICUztqe8TRQ
a1rSvYTj8I4LpC+cDI+0OHkyQEnblJDP1cv6wVW80PtSu4OcXt2VxWJOqQzoK28D
Tv42WYvVooSX1A4XVrs63gVRGoo5/HpFNhdI1lxfdoWD/NWVcA345Td3KNlN8hfK
FcaimP8K+bIJYusEfSimDkjH1LxxPV2OeI4PshqkpFA9naM9RgCxk2VbTjA6uhyZ
yySMk9Ow5vyWJoh0F89UGMILcCFn6Gvht1Tn+Pyi1Oe/bE4Fe8dMp9bUH2+fqYSg
Rmel+kqQCzrFM5iUTGsFmXlmgjT1xUmj1lDa7R13rrsIL05QlkFKqfPhQnn+BaJn
STa2AwrIgg+txJHOXCNk3NRZQ90wwQLbPyphr0cBOkN5jGpYiaelV+pHOEhy5zUL
zdt4kxMLnIyRpZiqVpDIpNda4yi5ohtnUe0YUz6bH/UsVlHWhoMJtBjenRskPj3I
yMNWsamHzS3c6nTE17KKeGf7pMPgY3OkjkegElEF49cKQi1OGOTOBM4zdbua6zE/
9nsvnqYzB9SXc9GLs9NzN/MM9fY3EX+Kto4lUFUyNx0nrxrYdwNku34QBtVIEJ+c
b2MteKa29aagfJuHWSx36TjMfD7Hv23CM92acsQpcHApkfidr0T/eJHZdM7CNN0/
NheDS2kDGOqY2yJiRGygCy+M8PMqEZOolIYmJyDldYCUOS/cL2jHvBxKgG/uMNe7
RV9vFPGow1osrUYO2ZQcTjMIPu2lbv2dXTUZh25Xy4RFt4Q2ScnpZhGkYf2tQikI
MIPIaM9nE8T1qNN9xJH9Phaego3uDgGjgih/Ydhuwo7z3/wdAZqNW9H1ts+Wglnd
StC+2BNFddLMZgDInxKfLf45k690pkmv8wQGu2wp+flAauberw5J/BK0PgB14eeM
7XfBzcf1JmYnoqKSXRPQM8R/t+Prg+fj2mB6681S91caxjgi5Pr2vdBGLMJS2C+t
10aQFpmVcCECki7MI4eMydRXQJ2RQEa9pvWjfaZSOXwMWOcWLtEPYT+5L6Q+r28w
H0nYxk+E5bDuM4IQhcFBvZxoiiUb5kyDgV1Ok0AgxeYJwBY8SPQmZrajMCXfmyzY
1y8XQ9Q/VljbErIUFeUWgN/NKfGkguq8wccFY+QU09b56ULAA9yo4TF2Ryxpi38T
9Gk07gH2SA2ZnqDC9Bcty9MklV0IvQO6ZFBXmerNoU/qEgJMAzEXgVKwaU7I8cgH
8c+tWkDCH4rVLx9KhIQQo0xD/94g5KaWDHV9lNPuDBLqBPtvPbsa+Zeqx2tHTAL0
TyfmLZoFwmv48wrUSEI+zCq/VbW/3W5F52mZulJZyFgOGJrnwz4WNr1LlcHPQy2l
WRZG6QY2frQnC2JP8539GATtMTMcVICTQMblAG4eHKFKLz1BIK9kqkWDkHxb0p2u
xV/3TncXbc/GI6YC52H5ZCA4VsOxp0U/y+2xBKMvw2Vi9SJZkKmPXarj+IoqioVG
zENxQa1q2h53zRQNNsN0fazwx1jmzp9fSuAkC+CvJwGbQWBY8SAd+FAENLS+Hy1L
eb1mVw0W4BiYerfxK8GEKImkEGvh1LTr5pwBkVUH4fR5WlWp0y3ILlqzyxhsjoIG
IWTHR/pXx2Kkwb3A4H4bm44Jh5emwKqx0m//vXoPLcz3jFRoUeNWFBONRc7UsrO5
m82qSFk75N7QYcVtDwXODvV6IzJwzCvBITEQO/H9/RT2Cf5WxMim6PuAcFmHpk8f
XFM3w3aGM6nBx0Vf+fAFBGjqbiSqR1piVrHtguSUkVQUuAhTtigvHmVWIuej/fXk
LooUciFepXotKNvJoPGmubhv83+PVe4cmwm/S9Pipb9grEZsqTRVApM64W+NjIVU
6A/b+mh2cFKbQM5419PIutObx1AznlyRFlylfgHSn2VdzYg56XUO73lRiB/P+8v/
VSyjPPT8o2GKpRhsimCSJr3wSzP97SPAJl+dQ+r/tO0paqtFdOecijbWWnqcTDwo
Q3mAw8BhzHRSDJC7ZEaMn/gYF/PKz9vTjs+IKoZE1WgM2IWU/VLYrruVjRLX1WPU
QeKNlyDjED3kpxx8SDsCxiLpoucqCQPRKbUvOLcjuw1aeZxEn7tyvDhQhzQtgpIW
EQWpY33Po2k8KU1iviFWHqO0dRKo1phgckWkzbbquW5//kJTJW6YTU6WhFaHI0fp
Sizxw1gp9mUx/E8xNEjpl3U0qJlKyLzhcT+RXRpGleWkfYvuoOMYv28R/4qemWNH
MiAfeQNST5x/fOzXpfLvpIyS0s0LlVP4pIOITlCMbcA7tLD2zA8PdFeOLmF8KDLr
jalLStaTWmJWgxMqXXjC1JSLFg4Bq36BFl2X+FHGkoS552Lcm6963hF8asfMFieZ
wqR/lbbSysm8GzXxuABy/jeAB9uAMqx1/N1588rTExMI6dp3ZuREtK6JbHAHcFro
vVNVc5FUPfJR2g3yTAfrB5MkydprkG2Se2hAo8CvXvclBwhVjyWO8m8uHB56yosr
sLxQ87UzRXmloAN4z/vOPbDJhGrGenNrH91fWbVwIg6GtHAp2vaN15uc0R6T3Wft
2DZ78MPSJP+7HjBDerWD+3yscMEWSQcODI9KcMF2IeofroOfdnJu+wAE6igsZ3Bn
llgD80QA9YreYKSG+4SraJwSdolUXSl/fDNqpbvs/pzVbirU0pPju3WB/9grLYiS
KlwFP/CFOgyVCj7DLDH4m6Ae0ZU6B6sAaWpVCU2O6jciEDnptp4b9ASyI9znSMqH
PtVu5jzqRjF9yz8frG2hJWUVvq8jJNH8oF8w7ZlkG+PE2fNuFr7HvLss/Q/ZqMsu
3BM8W5mr8Uk+T3PkvJUTGs2uMlRrw1RGi/xR9VxlbejrRA/xJaXxne02WTGEZfVu
5u64blbcvgiB5EQa5Zo36VHWxE3fUjPQ58IquvpjPRGHn3DwEr9yM40woCRiDJs9
esF45Mv/tPNPg2/fgALw2qNKgZ38DNv/ATFXWfe9z4/eUWjy8QGjP/U9jfiky0gD
pjU4/WnNjpTmienv0RsliWFEdAb8Iz9JSqCERrnCNq1tUOYpqkPlPtwOxs1Tc69Z
gWXI+7/bqajJIASJKGyjT3evDeQmvtCLNvKhksn2T2oxlSwyiWy2f1855Ejh7fWb
vf3Pbh12kCH6NzMnebuZovYtuK5BCkLScRlfd2aawN9aBxDQ+upk/aHP1VfrctfA
8ptdQW3UPfA+TUfL2OPerDmRcI3v9auxBzpbIT+KLsZqyfHyWDAcgJoWFi/thE94
G+Dqh3r13kB+Fdn7NKU3rSRTh+PxfwR/r+fV0UN/mTx7FTUUze4gdVImXRCP25Qh
220kRZ3MFpswG/V8Ndi0woW1P9iD1EZTEFN6f+Kgz+W39TjO5msWt8Pbr7K4ikWp
/tvwGM/V7KJkqkFviv1M5tbl5QRTUhOfFXVAWknInRMLAbxRQ8dM1gME0+GcsXY7
USpPV+uhOsFKX/KY60IbmZEa/TLBbl2iPR4QD1ew+4/hkPKPek4pWU7JMFmXnNCM
geEHPamyKTEfPw162AYbvjOl8KRzJtpYmJdi9I2wsP2w9dfBVB+/73AtUiUHKXtT
F/7U2aqYof+5eV+TzXV7PpWh6utA5iycRab2lr8PAi7mYxn9FmBIYSZlgsIujVbz
y1pBE6WbMAX21bN1jBJcJ6F031Bf/raXJv7UqjfOx9J6BB9Ap5755ludQf6IhxYl
uflyReCnd1kOtflltuC48ToS0b421881HNIDywzbuRMZQQUCictgN8DDi5zZD/Dy
Mo59FpnqbODT/0gqGbFf/YybnuvX/W94WsrNiOI6pShUQIA/qtYbD/7v1I0m7KaZ
xMPhZKMtmb+1ayx+AZvA91uQ0INxg8QdiqJId0d1WR1ZWA7nI/S+R98pe+QHCOLQ
g0iz16M1k5wj70jVeJAcULl0ywNr68bWeDXqZ/wniZCdMZ1/GApoePKU4gKOrsVy
/VyKyqUvRl9Ke8BCLYpTuzsApVgcGdOUBuJyI80FbdsC9BJW0rhZyn3ZURBc/aD9
bop5Myz7A93RsQjc2/iFSig//jkQxLGrEKg4LWYIYl+lHopMpKxVZsRrTr8BUWu4
d2InFcDPjXH6MFlqa3dLbFf+2siWzC5ryUQtk2mIJAQT+LW++DBEy0NtICWdzleA
S00JJdnUE4/zu6NPMWxO8AUwvAE1NiDg9ESR/ojJMTXMpd8AOq61bCO54LXf3hgb
TNJWC6y2hB5pbqkssPeHUpoXdInHj93QLdyXZCbxZXuvvQgY6iiUtkMmQv+KvbrV
QfWle8mRxx+oOpGFTpVMEbMUh10hNMbtEeaNk+fZfq5RH783LX9V3cuk0hFFccJz
0miaCNNialwAzU5FV5UfgPWbKtv35bk1VwXDrwVdsjQ4RYDhZnzFhTHhloDEQSqQ
DyYlPfKbf88AYf/dKXIndz3Shew0s/yBhe5wVelvg7nByd5VhICimVWBpFCUHxxB
IkJSx/UeeRSUwlVFTKJEKnWolIbD1mtIOYh7mhuPsA9DR//GV6MF4vNcbhLv3ZW6
TukUXQbpZBpnbXKKQzDCjWhPcuzKSuXANGObb7IU/MktH+T2modV9B8yNXGNhiJ3
zu8PbKvRMS9Ee3lZiMdemZiwHhFpYFFnqWxCsDTsdXAjagLvzShxZnXF65kOmqQ8
ZJDwNrR2x/ylx04qW3CQgKFc7o4RcL1XVr68nlnxK0duZJ58EnZYPZ5oY1GC/PWY
xwztZiKQOc4S2CL2f8ps6V0zTXixQ0v6+Bv3Ys0GMBZC4X3sRUeslqgV+wuPw9fi
vKuWzWTQAroG9NFtDEWcoyH7E1dcfJ9Cn5W9P59p8WCP02iism8KQHL5wscL+ApI
LvJh/2SwFw4RuJIhTmBEGthAu8TrLtIfN0ZvC3N1+3Xp3nDZXbGauYVweer0uInx
NjQpVhBLDnlff7f/vyUYcFasuu9DpklcJrCho+m96sAoYHX293BBlcx9AjsOdpxc
0uoVVqa9clKQg+AbQIC3wVn2h68uWrI5djZ2beeW0kNS7Zsc17NXfpq9iO9Y4IXB
SIZykP2QvrZRBdRyg0Qgn8NZdZBHF+hzZpN5ZimuaR9qu5DT3ZVtWAuj8i0uqgWi
xOGzE9EjGtGeBalM4liLkVCuNBHAl3k0hghWHGHGRMHlZ7aCpAqcGITjscBVZT0b
u6bpSXdGUf+Chr+MzaglCQeAEIMqbNZd+3ltqFP4u4i+KNUBBm9OlftBR1W2qM5Y
YEv4PwOW3XdZZQ9mcVru/sNWpQfpmhY1y2pnZYwkMU3n0Q9IXLJj+k4URjJzkILZ
Dot2qit5E/s550q81cy9Y2YF8/YWoe6v4/7gqLI5tORXj8MQ7+GjE+yg9lIGY37r
oNeJ7quNbFSTv6nfR8mVLw4Ijg5RllLCdLyNRJBZU4NvDNmCEkXDhcy8IyNDG1of
Z1XP3iFOvaQEKnU4UUkuHVzXcnvWp6yFdHKJfhOPso/9kIdJeU/g0EC5rzV02IRO
rpqq0QB0fAi+dILRXNGQm8fATO9uJ0Kfzv7c0F+AfOS4s7srxHCkGuj7CAiU6VVA
mBj0EegFRaJw//eiaUPNu+abmdUHVxaAkndR/QSwtD353diEY1cFFehEuId6fdUI
divzevbiA9MKduYNINswEtInBbT/AxgRZuzz8dd7cgYBahXqHiOGCb5IKiPVDOve
ZXWmunQEOjJQP2HSRwV+SgvNbEbooYJtp6jPYiYUG6o8C7aauPvTj5TEe3chwX6M
voC6fmNsuUVAP4OhrZjIyOLhNgwYvi+Gcfy6T8R53gPSfNNTeKZRFzHw3ctfOtLh
4YCksrOT5qeoL6nKeudQvtZ331kmP2HLGhEKbj3lqkHQPwdx0eez5Z+1DdPqTLI1
C+tEOpqjH99+cxNUPTXzjFFXveh8WvJWsrEeckut+5kFmazqh/ROUznV02iwXCvN
O/OCoCkhoeEmpM9cioDW9D4UzbYqo8aXFPJ7Xa+mgjHPnqLOpr4fzoYoz9QZqZFT
jJ+/el+Zz+JE1izPHAmkEWby8++spUTYPHuR805gce2OqefEPPC50gZc11tko6Mm
WFqopjomGdGPNicHJq+n2yWEuYvMzWGdjJFKBMcVAMIA34vKLp/aeVdSbTy+U0NF
PTy5h0LkM9UiktjWxULTDdMwgMGluZqfGxHH2QgEX7uZEuhPNpr06UJEOly/cd3Q
VkIGOch/J/9q9pRCx/SaeQQdUgtI4IDwO3xzguV7pXLNUp+95w0kEKZa2IFc/pA4
K33mRHbPkYJ8/baA5WhlG2+BHrR7AC5OSRcLjVouDJ/8SEfn13tRwU6MJ4TzoWn7
gw01cuOBvo/o5Se8e7IJ6W4WSdigNzCzU+7PqnC/qCyjKOnguA2qj6cQTqrseylI
JsPCiMfQ9kd8TqfY6rFR4FoulZN98UUllgXa+FrR0yJha+KB/sLJFSeP/3AavQ+4
ScF+XgMg5vnSKcO25Dl8euXg8jKV4YDgd4Zh/WCfLDLVB102YnxxQbHI/SWUUGIg
OhbPxNo3qXSn/4vEnBoxr5hzEU3oKB4UdiAFwsSWuapjUl8XrPa9hyD5QDcoSzGh
EAOvFy5hV2/NPB81+IX1ADC/XE2sdqgBrkbRpeT8m/V4LC8vhjezEVTPkiPlt3z9
4ZEx/mKYRmrLmFY7MmtGOxSfdp4rHUbalDod+2p3V6seLBu4ewsfy/KwvN/j3Mbk
JaSTbeJQH9Z6vKmEyXbDvSBnnmhbZOpDo2U8lEGl7aWA/QuFKcEA+z72PJW3ftC+
XlLuMigGH1sP3/uf0K0vt9xk7fgV20YYeHdY8I66zTpgqVpM38qBpaWqn99FziIx
KEDKQe141CQTZCc8/l/otirbOz3CKpslQ19weDrii6S+WyoTneUwfaApfCRhGPot
ZCOgvvmBy0JefsKwTH6VzM9BznONL1qSr6IH42dh4pB8trdb4Yj3q49Fr9xo3BuN
AaaK+E4wH5UJIpIuPx3CIBs2bpf3dwNg0FRGP0nMc/9CMZtygFZfQqFJfM65u87/
gFBmawQanrYFxPYE6nc9umj0twFoAo1O1rYXuPuf/PBs8XVz/7P3Q2GCsJnv9ZwC
CHnvOE3C1fE5VqeBSPIS1MXAdUewvxHSXYY/USycH8Ei353aNGuDJjpkDk6R0kSq
3LpD/ZgZK6Lpkj/ZKMXf63/x9gKEfL4eXLa4a4UGJZHY0Csz1erHLeOnPJEA8yOp
fdZr/lNYPryQNekGy94ktswpJDXsX/DZSCQg+ABn0eIbCaI4iC/lej6mgZtdComH
d4gYqNBHhmIYWCx9tFkn7couAF/wsBcTULCpR9xRqGpWiqMZ+NQLXHcpMhh+fG9A
RiqgPfoOh8mtsoWQKgJ8lrOKNN/GbiBvYjjn4GrxkS286WZ9I2Q7RuLEh95C9qkN
Xkj+hv1hbdNZEUTF8fsTOXTd4wwuynBHCqBDAfbZtFA1egNxiQIxJ5TBIMtL3sHf
dsHL3T+v7vdBJO4OmcZwBziq+VI9lY61ViFZ/2Anp3Wwz4TuZahmohReakkX5EW+
je4KmCTlzJWgR0Yp8Djy5lkP8IaqMFspHkAQv2t+QSoMDpxkvEbIAhwq3BG0jkjh
expPKI1pNujMt0y2eLLJBsg0gB69NO/PkOMlCWSSXw2mRhCU0ssoWesG4OMub8Rc
hUdTbibn7DUR8KbXwArBi4s1/vBxUNZEQQDWfPop3/HXyjbWDXagngU0/xI8Y3tz
hThDBw7z9kim3HR0Cc1Lp0zYl9+PlGpAXEo9mbYw+HML057SYHZu2I308kzRzlQc
FM9+WffcXBX53+Si4U5H3nwtmsa48F+5SV2b4kwflF2TqgBpT95b9Qfyv9ymDV8H
teYquz/Eme5tKMR2Ou5wYUDuFzwdm0FNH72PIGWJoatf8ee7IoNXoPgt1muhvkh/
xEJcNlbWzc6MNiCRiuhuQzUpQjVZoQdeGtEbmC6neUe5XnK5wzNgcUyJLO3insLh
Nk8GONt+tZUGXJEVuQVFstuYrmeje96/Ne6igkn+e0kOZlLEgVQP0bllEw/svXcz
kXIp7c7m/WWuqbP5C4zoInjL1jPRUGhw17cOdbDonlIKJ65aNzb9OVudkCE2XLkI
kwJLxjPQHrJPq1p+RFZvkLaNAdaFmNhLQ7lxN5cpokAUVn8FsKDYuvu5mXZ27KCT
0wEblzyoV2fAcqK3BLZYidC0MysPutAXwMB26KDbwE+zzlfJjNCzZHKVRUM6CDE9
Nw9PQPR2XcVl1QvOfYVigXgWBKOYQG3498BV0443D51wXGyXq/E3K9mXoaT5xxWW
JjR53DLwmpeNNWa5emsCm0i4yF6WkjiRvp1vI7oTh5SepbEjnYolAW4i10iZHpLZ
6qZTsdhDLj3uI6otNbiFuxcfDyC+p8JwZQaf19Ldysn9Spb0TTmDDWPqWLlvq6iq
TTspjll+8cJNUW8SMAL89jluFcYRGp12KVV/UgzlSnYJeNTCDiezz7T5E8e61fO8
OeYTYQa33T2nCwP/LX/MnIOF82xOtlXlWcro8CBwcMi5iPuCpk+5hC8P4u4GrYhw
4SF9e0DQVC6fXknALlPpfvJ6Gn7nydM1ylixRjOV9M44aSfI/RV49k3j7As54w8v
4ZM4OHpgun3VBU76CD8jl63XZv2dMVz/hRTxG7q1QoEvxLiYfp+lETmyqHiyDzTu
p8lHpyAcLEa22cW8e51qioJI70yxTPsuq4yBOY8q5JzR0J89MFMibSTOyNXYwHC5
ey+8AdHaNkxog7E3QO5RJwLAb+puo3mCdS+X1yauOyBMtwO7HOHcIn1m7D/Mci/d
mVmzKekr700t+MdIKD/opqxCPshUaO0oIo7n6+YcXCRMRDGivQRLD82Tougmym5j
GtVwOYqHA2PyTbX5tsD1oQdvxF9Pr3iK8DLCDt6RMgD6tzxqAr3oHPfRoQJKW5AI
2cCkBUgOoBNVGdRNXMDzZ8AU8dbjH0B4ws068Tqz9ZKwVeSgNtsUcCl5UgvYCUhw
KZoMxL2V2UtBDMTYrwYHJvWuVkJOYUjlQ1GdKs5hygBCFzLyRTrgra/rHdhbyul4
S4Unkra3pYBTAVPdVPv9nAAmDBVC0gXw+BpV5vrarjdrD8fljr85E5CgTrEh/0B+
zD3mgerfsiLHrMhEM/bb2YaWX705KxIELsRSAG/MwJXfTBFjqCvwX4cbiGMZmtcu
t0KM6Xyb1gqkVuowYiUKEKsltfkmbFmfx6279DsXOo3elFAD8+0CSkUZvrDZ8IhW
UxEdrfuanHE+mfZI826XmKyzrAmLGDAtgClXU+QUtLeRGAcyPeZduAlgizkWJklO
2dMujNdB/eH5SMUsjk0OtYWFwUDcOT8belu3X+fuDZUWyHC1LMlbynMKXUJJkW4p
rqTobRS3LoOSXoQY+8wsD8eNwIQ6jNUj+qHV8WMQSzeAJsK1cN87En5Ufmh89RMe
SyoOGD+VmOiL+rPfl+LC4bTRvHsNN6BTKjFQi1jcLJ0RrkPMeXHaqGh7l4IJPudd
zlFK39QWUUKNSHq6ezktSYIv6FRaP6eM5UdC0vBUQqpIeQJG6uafC5EjZcQUMjqo
pVcKd/S/M5vSC3+vD6mQ+td/EblQ+yeY+ebgSOXh0tVExxddh/iz9OF+2dyelb4b
7VhHeASSjJsASsrTPQ5eszPZjDr7vTr14rREV7fa10gwhyqb3RdzIPUUhXHdkUni
3LXAgSFIvikx3JtDNgskxKRkUdjvUo8FnjDJQCxx8mwCQVL3zRC/hoA5Xrxiv4dc
+3gg20gSQEJk+dGGdwnmfZ5oDid0bL50Qwqpj2lHC1i3doAOGUEMB7iM1Pba1LBW
k+TNIcm+jn5JKlfnT2NlUqvEh5lKhmB4el70tVRM+5l8Oys9eFTTdTn6A8Me2oG0
CK1C6cGwy6fQjBSNWlc6yKiOldu762rjzBD5EH9X1SJK4d5WBP3ARkb6nj9U0Fb7
wLR2GX0wXomPMAlEav055+fn1+IxsQoLU03U/D+5/+2cZMj67bqPui7MSHVi07VR
FBaGkxkGbVUJjrtNoWPPXFLA0zFoL3Yl04AoWmVlzYxE3KzyNsOJHlEXAMkLDYFo
RcMw0eFiV3+NiZbrZSlVzr6lPXMUsv4MpBwobzZ1UBEi3+/AQ4IY5rRGn92B4SSP
zJVbaiLGob++ejAs0Uk4qhl74ty7THj11Phmw4f/rXuSWwgq+18HZWgyVuQf9tbF
iwHAUtRy2w9eK5sjhUNIp9FRF05pF2ocnttd4W+P1KFrIgwy/Gx0XwJO8cqRJnwb
lv64I/PxGtFWoOMnceLfxdg4ejcbR4RWTRVXbvHByMsehNWmyD954V4RDL2FbqN+
L/ghmmGXXR+/e18uqTb5ykVtpMCEKJ1Pw6yDXLGLhXAI7LrAAQzbPS6jxdC60RBu
NTkf8uXKlarSJvvfoCyZh1F3qK0M9sSQnmkpE2KXQ7AsAMvUOQWC8rmVOW8CB5BF
Xij5CqEznWA/DNAwTNtJh20NbZRVlOIQaCbtNPYS7mK3g1Twi/cJJVE2O0A+6uUL
gGvdUj5Zy3hYxrUflVAPLUmUQo+vJRwYdBjiMFrcbva3Sd/n889vEiFJTN+vjE7+
GPtvjnm73V5+6T42MQJKu3g0lwwrNuy+Sv8uOv104QuXya1bquNpxzmVwFMEG8Kx
cca9ChMVUTkRWHhBlMwb36GjmPpq/YLmLvAKJwguuL58SR0d5mXInmKy0slL8mq2
xLPyopYIrolp9OIRNBbSeqrDxR1b5dNNSOgEL8Iw1vQxIYoxAut8TLHOQrWRNr0O
qXqW5Eevy578cD7omRCw7qcU85E2vv4sdT9pD1SpvilzQgdQTAa8qyOmceAMjFOo
/vpOLdEeNaSY68PWBwyr35KpVbTea9oeK49vvaSqu8WWYWOvbykcoiyQ7N1C2TzG
8jQzOdLgJyePoDAHXRd3qdPlEbIZ2AcZ9ft1AED0rFGa1WVookBU+P9CnX3JYhX8
/RsJOyMCJSbD+7rsAc/LdJwFRBgndHyQ+N2vBrbJurmYlFDTamCEyubkWHXdA/K4
CQEC1+FZTMZ3IMGlV82UNCrpgWt4qARFzDNc1sSVZKD6uDaT1duWbR30Kqqy//Hp
CM0DmPxa3Przcm2qFp8TmHvvPeab1+2QVRStU44mDxxKJLwuT1+jsT9wqPLhdF+N
aLj30MjUgo+QxKbJPo4v5auvq/bkblHJQabKzQ5p///7RS6bqnY9H+BFt+lpU1OO
0SuYnXcAPVNwyiGCdfjpgXlsYxT1Ia+hHTsNJZ4Zav9r9Wsg+JipXIA48Cua2Qn9
HxHrjd448zbE/VBWC5qw3or9o/gaZs6hl3G2l45Wp93oVcX8ml18epCG7sjpWyZG
/2hklsuprqmA0q1H4ULxa16/wi270cD0C3Ngi0zFxXYYYbhOJ9gc4rbwxPsySlWg
xjpfZOPZdjybs2D6cLuJ8W5TZbAsjzsk1l0IdWguugMKMJm4LmOwylLS5blpc8CP
1KEm5tQd7zzQxsv6MFZS7+03GjdF+b7Ad2ee2JDSmW5CE0op+/A+BfYccbPijdAT
YRqEzt/FHKKB698UpBhUDmKnIaOGom3/OqZJbwGkPvlWP4hIVdM4hwmSWQhme/Df
OJymY1p3VMURUd2mIc+TQ2DD/DIqClbkMr/eDxyG/+J4f62izZfPRFWds7HKNz2j
uKtv8qwSLYD2akgM78agAwjytxHvcYv+fqula9zJQUdzox9qb5RiAlfTWb0VJnYv
f974q0EBbP19SXINOPIo7v1Xt+YSL8X94MoJAYoQHjfhA7uWc6PIN3sJJU0oZiUl
VtDbpRdAEHUeMovIOO0B+WUXTltrLb+FQZy2whIBRdsYP/nVkDnmwNlU3sFhU60H
EadQBc3R499ydIV7+aY/mAg6bRLxYYUB9VqX4YFNHXZFR5m+gF+n2zgbGUQjyOnd
YTp2+iGV4AkKi0XWi8+VzcjsGdZunXDBuEIzMVWcC4STg9Z89dWUagVq+ZFkX2ZR
OJkGTAqwty35Et6vURI1ltYizIv4ZVqcgj2Qc5F93/iL0T+lAaKFPxo1IeLpG/bF
cw+1LH2du2FY7LipOkj6k6HS0YztwjqfBrVRmNLexhw/h8B44fzE3lQFLF26x7CQ
O2sMbbjLgpqSNfMNyvqbbhSePsixKKsXubc1SJXP0WZo/AKck1K3z/3KcYonjm7d
XWXElZ4DseRQ8mR05s9pVegrRWGBm8muRaDyM1E+gtKtDa0m0E8WPz4Ovi8B88vR
D6xpNDZWss2Vsze2ISeOK9ECEwu9MLxyJ9J7aHpRXVrYnjXsGbSCIUVzzqmIP9NK
U7CHD5KwIclik+fqoPOnyLnAflfp3ZERAQGK3pLG9/pxVeMP0cYGyIDMG0ZMyYy3
gz8+Hi6XsTrH1+zYSj61cnz4IWxUWyxKuFkgarSgn++XA9p1p5WKyKqxQx2Lnc0l
Ab1zlp3G0Q/KRZucyVuEf7QWUpRpZFo38vbevNfNloVzszFX/9ig+PN77rVHHbOj
quF+miwXhVYMVe6aqWjI3mKyaU/uJgP0xTXCHCiq9fR+tAjOlWYcJCDZox6XptYt
3zwKRlRmvNcItRyXjKZG+45Fv8rKMAnnL3ONLDe2ZJrLldMahKQlDQA2Ly7wh5DL
OctzKb4Zq5tOobAXFpvG98Rtd0x09Pm/mt7j/fXTASVo1Is1TBx3+NhHVq8Whh5M
tXgNi+OWuOJKI+/BQMYrKLotUwWiullkGrbe/tLDZvXRC6ZNx8FPdRlsmRo54NqH
ME8qlQlAmpAK9Dqgl4nhe+wRQox3U2TJhpOgFhdJoFcfzyyo7h9HGbRliTUUTEg+
Y5ehMkXiiQw+3DGBSePwD06fYatfvtTGYqsTv7e8RByKE1IdtV9ljN2Ylz7grAQK
4LfNHaSG5TkYG9WhKq6TITay4nQNTRYlIwC5gYB8NEEoDuk0WlczDFjxlzIWboyY
j4bl9dEpSs94Nb2pFCCz4hjRAuNRa+zqwQdJ1Jw4/kjBpSzFEhDaIqVbDlUl1NnW
fqmvYMSSMi3+lGq+ajV6vlqUzwmTfNKdZDgCHymxwwB3twVLN3vdGVT13n+TIpVS
hv+7jkMbx3kD2QSLWknTt2TkKFnWPIWfHfPQiJmovxNp/1+S3m5Bdq5SuaWMV74j
vkNaxGb38Kn+AMIscV83kxOCvkf14Rtlc7o/w5hygWvu2buJ/xk8Iv5yW+GDb30G
j6Rjk8pa+DLFeT45PQNVRJmuWt2/V3ZrWbVakijxpYCmZqszV7hovFYgh8YFoQCt
fyJf7dvLA2mjC722arCz2bHq4xjRCAsJeVKdbYgXOysfVsKvpq5uu3cYcjooC2nd
IMDTb10No0qTpI28uwrmmedWncqlQ0N1gShHaQapVEO9YWKPPUmQlsB7xv/UQhvT
487EK4GdyZjTSRkh5VM9jxSmj7OpNBWJeMSN2A+llzxGUX/h3BQEFfVypaGuu1Og
vn+s6y1TIVSebuSLJLRJZi4PSkUNZlzdY73SFUqJJ7Y5tV74qgdnGsaW/8pY1etR
kH7CZmzU1APttDdmGkYdlzfLtgB8UlhZs9tfmAcsSz6CpbwM3/aiQU2GkGlSlYOD
cMCfE9SQvOk4FMnvmF8kGL4fpQRIFudXph+Kr0v7XM6ci72koIy7hFhAbM5fI1ul
vJR5803Y9Cc17/krLgU3tIxP4dcSYab136/+HsoKbT/7/WtGLiwCPuEChUPdZlVn
+opzZPYw47+Za6DfvdV72vSaj/YU4/c2jvGDaVqd6+M72/wlEBA/cmFZXC2j+3S3
LDx9tu3k9tsLoO67/tpJcsYTXV4BDYZoCNTaiJsq6l80fa4dXoLkwdzKiRO7T+h3
YTcnmQlK1GvZAtAsK84RjktemDIWsojo1XUfKFa0A1NfUnEvnphCg7twAC/IP7fQ
w759F6rtksfiAhZajgyTmMIDAaCVTux9KJYrmv2UzJQNjnCzDku+mT3EyalIQbQX
dD6sVyaRNyGao6gwCPCvfyAxhAsBOse9jQ3W0r/IcwJLEmyKXES0D/0YhB/jjxwV
x7E72urHVcTPcoJ9kmFR0WYEyt22c117GRqHuJx8gFHyar0iiCxNG4gsqXhCCISZ
2Vy2jDthGaiHBMyPFi1SccKoClIcn63283O9HKSv7pkJYQxRk8lJnmUbN7q5hEC4
TkjJM4IZu+mNm9mruQcWWXCkKaCq3jB6pfwEK/7gbHVVeNRhRKNl6Gw3FU4/Z1JA
d/HgG0GYj+7y1qeVbP+jOb9QdHJ5mGzkN2k7+s+zYNzhiTTDmpIRuMTKmu0GDKPv
iy9QAFnfumlPFPoIUuC4Ysl/KE2ZeOLFLv553nKihfyagwqFc08oFGI5M2ojOFc8
C7FWXDv+nuyVaScKKuUhC12JOWJ1yoCZOT0GhcVEAlT6wRijmPrDR+ECYhpox9j6
Fnl31i2y63Glq891UosP3BwBZER0OLC/11WetCmhmwxORgaMHJuKCdrEtRj8reLd
dyy6wSqE9Gupfb8VHY58mBDIkyoudIikMS/7v045scJq5hu9+FeMNGOvl6qkZxqP
Jk8RVoPkg24JbwonHpHEl5rRLEdK8PEQeGHlJ4g3G5gFrzqz/gcQtc4qcTOFmg2g
NYETrU53J/W4j7OlYjsbhF/GbNRN411MRD7KVOK1Wy6ER4W6n73vCBvcUweGmBbE
AQBEmeRMsL3vcF+NmVF4gu5czstOeR2/pw2E5Nwxgy+x3e129qPHCAZcm1PUf1x4
E64P9mRjEFQYzmSAub/1/D010y24FY7dIGZlzl0/MbNYBUyk7xEXz6W4IvZqsDnE
ulWDQCx7bGi4Y2j4igyU+MSoG1vpMgmMf8ksvpGsVWaEt7sKbF1/Plp6nGbXnMog
GPiGbpQfq7AUdnfXdE4R08qyasF0rAWPSJGRrl/GA64gYQZo1C94/qb1kN0HwB3p
0BZB6QJwDM2F3TVdiRBmU3rj3kngGKTeyAncITKYelzl1h07iyCWkp3CXuQQ0bA/
EJaRwckUFYPn4NgBcwRuYymyxLLpVNCw3A2X5lMuO82UXqx04JnryaJ70qFm3aBj
koC/4OYhyUfVqCAuurro3H/1foiHHWsxW0tB7AjBrN9VSyVScenJ3l4vmUf9kkov
/u6kIx4LjuTIAKOV93JhqUqm9/UuhN0VTnyfEq8NDkCBE7YTbk5i8ZC6YwtAet/I
L2fHjv5VFnfyr/3ljipNqXFKYZZ1KRRO7g+PtLlxzMGdmTEP5iqQ4VPyvQ8/Xi8l
O4NglRxp2TVla+7yTb2QBSSZL/Kk8m1xBJYMVR+2atqByLf6qU5yNFINOSPDX7tA
W2M5NpYBhozNV1R4/FifLSNM27uPZGK4d8W8EpyX+T+WbPI/E7KsGKtQIEYM18Ih
bIUD7WOdBB0raV1vZGnlg24hJHU1pNM58gV1s0pMXnrBrqUXuE9ckIkNdReIEegr
nFEdpH7mq1/GNkBapMzNuUhlpizk3AqIPW4nNzJ68XsQsqZA3bCrohtDK/FET77e
L/cmpYp7n6xjRUOU3gTtRhaHzGUtLKRd5YGH1KTXynJW7h6ChjLy+GKpsvcvq1jT
sTabKMCE7Y8qg6aH1e29hGTxV8VHx3WAJozYTO9U8+Xn6IsMmZ0OKB6FTRJJ7D4t
MEbkmpJjj+OZXnCvJ1B0Ow8bnpVYjDW/P0/XsbcNnqI+iJiQiYyoKZ98TwgWjMvl
c3C8xlZrkk9lpzLyx6hrEryrvcxa9BeK+DCu6m4XoBYwG39DQDTPM6y/BFORA4/d
aSdiQX0y21h+ajCWG5Kbdj1VOIcjb1kAjmIih/GB+LWzs8QBlBMRTONyOtqwgm/V
uDI7+LMR1AaGCvfgyOKrpgCKGqsNULLOZ4QI41dmGU4YU/BlKkHMqwAlfShKRwff
3KOLgpGCrA9ETXnGk1814e2ZUFynaZ/l5yL6Uvrw7HnwrXq1WVwVQEBf2vxjtzcz
9vo2TbroXSiOlDVgttTjfye2BOOyuSBthlCa98x/Jx+/hO9tat1ItF/kwWmsHnDU
ufWhYd1kqPHAloo5mlO0IsS9KOtls+o3DBk4SkhtenxddX357kh4q2UBGLBKzq0K
P5qfonSkJinfjIbBgOhNGz34X595745wSipBmcTHR7FZaB6xgaIiZnw2bzXViaHf
ITpTGSFGHRqCWpNV3Ty6KS7zVW71DK8DQx0HCw4ATnsfnTjBinqVwCdRGg5XkI6u
hUN72Zplleppdg9Zjx4/+1mVf2hSzIortX6e1VZbLgArsJPtARaBj/Jpzc+CkQcM
kwiSE44+GIomoGfGlyR6+cxk6S0+mXLW9+DprIs+mCQgXNErvjKUclZ/IFiGMtIY
Q3bruRcmQrRmgn0H6RCOrVq6bdZGR/cqnTbeK0wl9b88tB1scJHPFZKOLZD5nQGg
frv67escDtVgenLOzErBDR2mVOh/58PKoB2FYjrG575ErLGIXSyK4hoj88AiQS0y
q+T5Y6OOIATw35rN35NIAatGbIVynE8cD08EQqFCga24FgofoHVOQ3itniwNOrhZ
gBhM672dMWEM6ibel8+Htiu4GqyJvQd9icRr+gcUNyGIZjAMYiFs7CXfIJ+H6wus
/0T+yWBEWP3KqO0us2B6rBNhyVpKpC4Sz9B6tucJDiEFVFTiw+2/Jk20D9cgpYbf
V2v5C6F27Px+Kn86xaEMd1IjwN7SUa/anIR95s2CReSJHdDgdhQ/2ZPcXucFkqF8
jCss9zIxCg3pdp+rlkE+puWIp3B6sX0OzWB13cR8ln694iyVnTVHMADphHZqm5D4
sXB0Kq047+A8tdvkKRDhGNmNtmu24iD7gI1DEaVNoGUhXC9ktg4rlXjRu5PvrXlC
mPnmDSOHkWlwNbuwmrg1elimzcXyuQeOegoMK2pCbYyMsY2LFL6rRDaYJMsip0jb
I4Pbsh6d6uDJoluqDisHvO08sp0hehLOOQM4shZ0fUMWpxjV5rps7Mu7YwspdQEU
hsXmpcJrcqM6rVgQaTlbc6b/EXJK/BWx/2Z1U5Qv/OvvVdfWwjOmRQaRw8e1hjmQ
GKhSEXBpCpjE2xLiZu+XUWEmYnCA2wvakyACHj+F+0VrnsddziUW6LQ5WRx2UE3C
7wwNbAK2IoAccoan+P72AJaMrZnb/4IKtnOAURZg8cnEAIGMG33ao3tcpmclYLm9
EgekBul2zGvJQw1x55y5NmhUCPW63TiMCGXfmAdtgqIjZKC+qWZ0dz7Xb4Z4rVxi
MAhoCuo32CzrjrZAftXgBXiI9m8zLYGhObpq4iDpl94fbTfe9W9Z3CNYZ0kYSwUU
50gYgjtj4X6yAk1vt3Ei1eXDq/REi6YLgJrU+aOJZcdlxOs2hEE/FERsv3XgVPV2
3cTA5qvSj0qF/kP4KtHFqgHNqZ6D19/ju8WejF16F7mHdu8w3rKrZsYnIzPU+yiM
pROfqKuBvNKiWE27OOU0qYYCqld3u+6e/HipLf7I0zMjgGl3f2gW3lYkBIOgi/JN
/1BczHaEhW7i4o8ooJYQ6qnNEr1MRAOcRnVQMI8dSgf1V/JyIRw8C3OSKv/9HFR7
CSCA67iM4uiSbb/RolX0Q+dPkx3V02P/gtq4b1MJ8ULyZHpkcPPEs+/cHN1fa9cX
najdO8cq0Lowkbi/0opxDaf5FU0VX4D5etGBex9wLhcxarmq5FT3mHfznWv2tLiZ
KooolNUPmm0wPtzXl/NFjkQPNuKYSv6lRFiSX3T1/YPHWAxSswlZioG8OKYpiiA5
veJi7apUt3AlxOPmnpVzbxzCcVDcKJ/v6jwt96Q2QJ17IHtqOFaOo/N0n5bznfS0
vgMInpBNPhTqI3cC/8TfD89Tb+jzhi2CODpDOfKupT00y4iZMgXhA470URFXlqu5
U4kSsdj6VWlotlODmAlU83xz2o9i2KVzCt/pKNwFk3LueN7NjxDP77KO6LdQb1Hp
rp4mekZRrRd5UmMa47V8QxKhDN/TH4XG/5YEwEA5d8FxkLezHOqGDDPtRh5OOTc3
PFELl4wZdo5G0sCG6oPE7OZoyq4eXAzqXcuol9agCDa9jsXVOjHse7ZKnfk974hb
FK1MCR0QFGhu6XM2sGMKphv+AdOQJ6F4Vyg/gT5hKZDLuzIXPriGD3HHewhhA/BI
fZRB0wzMLB+Hv87Tud+R+DP3feGYFeyQ5TmdBrDfGqPUUiNzrSc6tlL6qAZ+OIpE
oDUaSzlAyevpd3x0Z2cuhRfpoy1pFZUaSwJt+bk7u14cj0RYwvvdofCAtpbtsZis
7yN3QsKzlpIPxt8QgAE3WkcvYMUQcgXwSIkBbUvGtAis/mMP/PdD5bYkibw7gOV1
C71KwUoDrTc/al7XgOuBz0yz4WwMk+kzaOu28iFkvs9jBp8bMQdhluidZVUtM81N
VEkeOgw6WLDayd4TSWYG8adDJoeefe/Dq68Tt+ChorU+jNC+lRWNcQ0Opqp/8aJL
x55WXk3nb83U14PcHWA4YjnW6BnUIpd3BlAxaxlMgiqfUMVgmdSbvuT/rpFujFZe
/6VGB3NM2IpAi/OTL/EFQROuOlvyuujP3plVrdsspCSWBcF9NJfx5T+f/21Dmi4a
hh9bj+vlKrMTU4r4YhQJdVpVwIlFEYKPkfUG7Ibn28p9iBaNwQzla9FSuh5Amjay
GnLEsXho7+slaPYr6Bx5beXASoR+x6Fxkwcuv64TWaol9G+xY1CqLIRqK9yPTGIw
Ygidp2I3yT9xnN6N98u8mA5LBWdAc9rZQnxV98SeZf0eg/LC8pyKYBo7ryRqtpkm
0BTXyjvoe5PThyrCc9ufLWO7VWv5GN6UBgjyWn+3/CE/SK2OsiVzp0Ej6t/YhbjU
huB4+U+buixp9vrMAEeOmAiYYdm+Hqy/I+WFwQRpHHGAcSRpkP3rUzIoPVI4Miu3
+WAwPQXf4eg3ysjI1NN4qU5pe5CxQL0lPaBWQSz2HefNof4PjKpy/st6uRnnj0WP
El0mYNDbQXrMUBiY2DEFV2AHhsGwXxNfAHG2b3tUeNawXZjK2gQkIn0pegZbCHIc
Ip125nmqG/0/AhtPzt2d12WdNH+A2oZajfqYdWVHKiCD9zG1j7QB1iWYpDBgtWzM
++PtytxgUL7VbpBxmNjwcYuuG5OqSodw3EXpHymMKoHjDSXaCSZod8Z3ZdieCeNL
wCRCeUn7AYS5Xb50FBdCM+5LENtErElMeN1ymvSJnFLYLsymRe+9LWapey+HFhUh
/L3zhu+NUONruOCfks5ooMGVnoKEbdNFhs8nGsuvOYAUPOPnqjiYpfUsvnYzz/or
sKLbBIT4v9CAZ8GKLwOiwZhBzNVkU0DD4w9dYIqr0X9U6S03l6X3RWAhNZX0K/TF
RCrpgeauGawGTcfG26cDRPgPTY8nUARzYP3rpk5NqTc9R+rUe8ZVTaS5JOhCf7l1
VTwH00JkGw+N0ndZb09yKN33lowsipRNmkCwQoYNJp0FHMCLlay4+PBAvStK35HZ
ue2xWblG8K457vyrAda+PAU6MgTOOClO3Ng5qYrVgePbDY2zIvDP5Q9L8qH/4cr2
o7hXxUJlCXKdFKvStaQ/AKMeQGV5nKz/6iWsEOQ55G5U4Bq7ZFFHDR5T/y1m8qVM
ivituN6MFMQkPd6bF2MBEV5Sc20DLyoZSjpk69Qsx4ACFjdcl5k03VhDGZ7B9wJC
MPfgNmoc5RAs0KE5aHedGgrMwmJiMJU45w1yYKrstRcyjQ/1zoZU/Ik1/tVnLa9r
WCCAYnoCGvu+hURbwGRbNYJDqr0X49dA8MetwJJ+on+jqGMfYZ3/CapD9gAgZnr9
CtLiFpmP7GDK/+N24QizDrVZwviw7ToKNE7V3RHdGNr5SK7GfU5trW1bgRWHZUkG
2Ly7Dc6rB4gOFd3HLjBCtTEKEL2B0tS06YlfgoDpViepDzEP5nGlPmSYHWaVnnP5
YoSMJGxMGElr2d5CJbK3aPe+vbuKgp+t3nvMT6cAbqiBSkSKZ/FjZM8YBxB8UjmS
+I/k8eddmssB0i6xHBeJYwP732AT7YK/MRaKJUQFeKQ3VrRUn+h3baIOKR4yyuCG
12rNBFoQoui+bN9arda9lF2B+Kb/3a945q5crJihBdOAjTJdNIWEWLYAaSq2FvTo
OnsK/uLsk1Nzr6tZgLWV6SaKLUNW8xOEjnLTA+c65Pp7VMjvPRjN47P4YpVAXaMr
hbfT80eNIYPfYBGojRbdxRNChLUo73i4aLl5QwboYseg++m/yHul6EjnABO7gPQ7
jrZo/x3/s2EQRvXlGxptS0zfb2G9EYNznExWS/OTUIgUxf/mchL3Gn2SRee8/oUF
aPBQODSMnIHVY4FIMUGIuC2iCI1cvqzjW4tQFcAJu1H+1xdG/Vio8z31AKMOgR8K
pCV7LOGIcmvgvVSLryNijznindzkkBvm4OhN/yh87GWMUGAU2RTpF8yRS9bjeRt0
3+GKGnWvnCnSV5HEEcz9QSHoHyU+o5s+r+1mUVaWIIQc8AvQ/ZuuO9nyjaaeS/UA
/hpkj3DoWjcZvG2aiciHWml62FoNeAQuqU4ALCyQzXGgLxSln5RclggVK6eHlYqU
6pT5RK/SUqgjx9HYt+6k8lSzMkJOm49TtvONFnIFQ6HJ1ep62SXu/QGaTel3KWc8
Msdq0EV1gwrWT6E/4a0lVjILuSCxbraxOrKZXlfr5lDhO5V6pSoIZwDE+k0QrMFY
QWMgU49FtlPttszSqyQsWs/M9J8zRcjBL74Rf2NAfECyD4lDsQD5Flf665fKh5R2
y6LAhyqyXyoep2dlmHKmrtt/gYf02txkKCkhsLsHQHnaFojlbjXqrdYHQi3f4JBU
oOy4n60EM+3mA6JMkz4TR0raFqh4/UGffiZgdLyqWdCBT0Vw9T60RjpqkBNFBdlq
L5qnJtXGnKgKD5yjKhB9ojqoxYHdhUqn3LQKWng/I8Nhr1mFOTTEklQZap9cFxYa
08O5HtLqVDJ0GAUY4VxUvCpoxKxxCtBCH3neNYi0alytAcCNT5aejR53GgZhP1Vy
n44hItHYYcAlh+Z5XCrZ4v/Nxeiz6npM8XV/Yo3Ru+/XXYGzmZ2OHmVMDipGb0A4
QwtGn0cyvFJd2JIkpt1e7TIxOKxFFUbxUgmK0SMFEUek72jEggQhEG4gFk2a41r5
Vpcmcm0l1zBQ6zLfhq4ZVME0yPFk1uULdUlwS1yBmTwYAhJ0JVJv9+CptDZVS5XV
a4n/5s9f+T1eJNhNtdZen5BeKRjkhgBwIx4v9FFm/3Vuf7JLin/S/VyuMmeldRKI
EnZ34cpZH4PcSJoFhTKc3JcP1AT4WDXwBBUrfZNGEZp0ELCcVKV1htw0kfQrQh0x
XPLfw6lcQUHA5d35dL/YNFBxUuHLH5VyXJ271Jgej/iSleeCZAHh1F+gV3MnMky4
93L+VdFaQIsjr6Y1PNdWsIiLEfn94x55DIP6+fN+zW7KK6iwg3tao8PJcujqhx0e
CbFonwA/yziBTW15b6t+WzsMAd7BJYCblukt+tqHdXsNzgFetQBrRE5b8MLmC61u
JGhImvrAljN+gHXnTwLrKmGYGWzmofIPj7BW813CBTbOz5XUQP+u+3XB1l5qluf5
14bMfrNzPNJpnfu1i8xh2Hv37zFtJs0PgcIIl9GDG8zuJvkSHNsrh0p9rttX83te
1xLg0ZUDZGcpG5SpyFUfG//8IbL+2ZsHPHuoJy26vKgRSXyb4ROr06s67zhRYd7K
oq1rcLappT5CtsGxlDaTre1t8Hk1Jyb52CBJrNoxBQT7Ti9QmKSN3pZlg+zps8hr
Oz+vyjs9znTjA5JcLdqS8lShEmgpvnYU0huOZmLN1Xm2b1Jm+fK+KmwJRrCmvxoz
48dSMhq4sZnS91LqmVWmUpw2SFT50Pbh8xytXm+Cvni4OduwPD8jwFiAjxljRYUZ
935tJ88czt8NK2GyH8v74YbjPIh4llJCMBo537jZ6KhgFZAkvRTQYwygQQJcuAkR
ynimOqKCx/mBcXfRW19rXssH4j+5oNm7hhwxwrxEIqBBMxlK90Fj1KH78BF52gGJ
jztzoLuLapv1Ydk6qwS26hc4jYKEvmtkj1E9wGPIpgdYkUMBxQJBYkIpx7WE4cZd
GbJeTv/ljb3WvzcOubZVHfHKr1f35ukxYT4RrrS2EPXd8Dwiw0Leyqhcl+EZBu+i
T+9aoMR4quTKvDGrbwkzQrmiqXFG8nFimSB3XKOlPAh5hWA2pLdcVl05UeIPxk46
n+hzCVnP8tJt/YbEvNbk+Z1YluGMJnTgqqE5cNqgWzxzMVLp/MRxNNJV7E6VzcEY
GuERFOSkPlucCPobAhj7iiLpeIBDooA7H9bLVwgDO80dc0egt3BllV1Uo1LhGHOD
gh8oBvlWW6CI7q3rbRpWloUJCiTrhbmH4Rpg1B0RNP8mh+ADVpSasKdIYnfXDOvp
EcPo4p7gLySrcVhw1zwL9PwCZkFQp/m3tu5J/bt3mFqfF9nigS8yVpGcGxFIB/z/
Cbb5+VwHAvYF6SEaDlc+ewa5t3NYRzpLiLn9KGlM5ycbcDGrf+aRTyuT27hoDpOV
eAIsZ6xyt1P50PpoTyK7WGipqi3+/D8mh+UVFK9+dNLPVwMuIFX1cTcHb1M9XbOZ
wsVxy4kznaW/pMOHqnwKUCXGcenlIsL+MULVcVtD9nqh55uulFPQ/RKhPoGZCCdY
v+tbkfAHcK1b2AOI0+/Ljr4qbuaFYJTPw5icHG2TFkbDR7p1YZwEvCPLZMMhUslj
GsMqB/Uqw3VRGyCdHGO0G13FAjQWgoDWqv7wJ36ICkryc8QAspCwkwADWFpILaeG
QbQ8T/Bb6lpn6/+svcKfF0UV0KKZciFxMdmyQ8DSDhrIIL41GkVK3Yle/OUGzt6S
7MQv05rYGDFyamtHHC2fY/xNgbv3WCr1xbrbwAfUifsa+jSFgYt6jv6UZINDWBDl
x04M4Q2KahKWMwCLbLc+DcF7gt5b8QS/nRCK6dd3GPtlUfx3yuvbIY6jyE8d9MJM
g6a2V+rgJt/TKxzclRqQ1Am+lpQ9zmxBRtVOZEBc4vcjRWVBoBkXlZ8SiaKJokvs
MIUTU/z+RCIfv/jhSmP71yvPZoeS0UoGmG+aZrZvM0E5ihh2u8BntdZwP3CzralY
wuw461W87RhE6fXT4qwAOIwcHL+3zQXAbdA47nROTfzgC4q9DDOocal8+41r3Wak
13A+UoSvT/IddFFZ8OJUb6nS5IsdUlkusWAbaMorYfm1057t7YEKZRL+Rpq8m1pO
qObdxpEmTXAz3E2Lujw7Od5L0egJtptOEkfbltDBsKLUMB8MREDJegELWxj7l4YH
jnDqK8cSYMeXOz5LYE9cm5h0djRrDma5W8AVIj0C6OzvPzK/9SWXIvDMv/8DofuF
olY3IFyXWK9n5cwaTJxrd8PjHfBS+MaXmWStMlXzd2uzt+00vVv23SvBDq7dWy4k
u83UwelH/MAaephjVKKmU6zjOVX3267UgMKY0OO28WXiE6KGpLMDjnYXPtGrcHMY
zMgjC1hwATZDwi+ECxPIWkEdTM5nZdcjcPF6aPVZG46kjq2UXYeSFEFQuEt+EnqQ
76VnNDEtOb5hnznc5smjZ05ipn21dpaGws8p8rAkzhkRH04wjw2kNJoGHVeYCBlK
xT8nGMMcZUU6FgyzkK0l/ef8Q3IML10tAB2SG4ZQtVBAO/Vu1jip3XXScVcu+XCd
ffzvBLqGvefDt8t0UGg7OxbnVGkkrD8GJiN9Jv52d6V5jCmc+bo+GpinGM1KbDmi
dDFB2Z3AnnbFTUwAvaC5zxkvkRNlLnOwffaSMRTO7vvBh7NOZNAyLSVXamlJ20qY
yYF2b1U7XJ6t+ahitnvCDWSbcknxLrLKyfH6kyeQFy7muP0Mj6iIZQiHON+JnVmb
zVboPokaVoC3Z9YHcr5rRFS9tiQOlHwgzObtTp20Ak9LXD9d1Yf+4Y/e0YfCbPhJ
UtHHuQAGFviyQr+EOTCoyNSuVUQqqS9PwFUff9MYK5bvId4OCaB4aH0WyOP1U7n3
kfVrDtUcTFDZqT8w40UDaUOsomBJ3hsDXGy5h1lm3dO+h4yoUtkEnYTwrfEx5gDe
IIXcr0ClSanqiWdaUHbN/6f3OQ/ar4vnif3aKXEByrBMdmiOJCwLOSWReTAGTFSd
1AuyoQzkgONGbb/Re3DV7NvLT+yHyJ2fiOwwGFyp2DnD+LYhRSIUAxDfM3fdXbag
b6A51TvPCC9Dtfhrnro+h2fmdfEW+Dst6fh3rYcWdow9CRSst7LL2tI1Qk/XMadp
WCDTRjkmjak0rMr7zmODPQ4oWoaXHWRi0uGN1n5ZqtCHT7NVJ6FzopJQzoXbqXag
7QQWftejVhhwTrDxn/W/Apuylpp/JDYhDbu2JKFsHebJWmxtYIINksZAqJ1EuQdA
i1Z4scyQ4mH77MTYSn1bPCKyhYSBw+MhyUYXJKItGS86R3J5ahd7RGENd6HtV0eY
IVZm7SRDgdyi/dO7uj8yNe07IwacSwzI40fcOweEz3ttgAWlmgy8yK43vpYEL2YD
NiyMGOVne3RH4E2qKCmwZ7ef4j/WxuR6jJMKFyic+aqQ9cexlcPh6Ijlybrso1Y0
QVVCk29EgB+RFvCNAP6aY82PbTxXgLjEGqG/dKBZRDKQlWHxmB2qW9caAZ9bfeFM
R+4EXktVOwcLrHjQ2iT3MGp0d/Lo4qKRRVTDsF+mbM56WCRtAmIXGocefriSln4b
yjCAihlSDbJYcP7zeoKl16PNeYrYfsm+Whg66ILWuoXpeWs1EJv+F01OGUax/aQp
du9FUjR8bxoZiKBmRPnyffWEVzySIcq52Vzp8+0bbNIOM++UFgSUF9s4MsjT91qR
OqlBYi1GYALnIrwZz1OEkrSSSQNfzCpde3/RZpd4iEX6BBTkGO3oMERTNHQ3Qfst
ZzoPfg5X7+T2M7yPimzA6m8OjpZWHgtjYK+ZlbJ0BYzbww2kI+42c1ZGynx8APGb
ERvmkuRvrc9m8nU7QLC6akrGtstmiKhQXLk85Q40zuV1pzfS1gFlmMhHAuvS+C3I
Pi3oz7cMg6UDtTWOrY/dFh54jXQWXkPhwLJgY8IwkWyta+jwW6oFUxdtG5RL40ym
NLo7qxuQt+TDkbMjTGpIngXPaxNglx1+ZCbym+s7lJss/YeuNXqr+HDf/ccCFAQB
Jx8xp35W+CzvdHQcjXZS8J3MHU36Gerr/pK9y0k9PGzF8RTG33NoTuGA6nRqZT63
tgdd7FzzPkGa7S8jkH2ffrfg0v58NPU8PrufApSvvwv/gHPPZH1IQ20uXdqEoAIl
XX5Y34BeWAcLiX7OMe8yBjKG6IY+lm/tZmXgi0Hcvk9nI7t5uwIbiN16n8BY9DmV
TX+obY+aD8apiSct3CxKegKt1AVYmF1RexdE+bDSLiozQqbRiEZMRRqUNEsWe3za
WCp9+2iKXKDZr0JjplGpKp94frsAf0GfZ1H8uf6UqPONSTXxnNQ2jluAin3yL2o9
atkFkB9DYCMHnEyrX6Va1seYb+CFBPn56Hhxz8t+//gaye1WcBykIFbHXubrEctx
mH85xAI3koSEMZBq3AaCQ+B3gnyWwePkNALmlsykOJbCaZ15619IB3IX55Ou/k7O
XQoQk1vWFmLRSCvWKuE3tqy2SAyQHh+NXDsdj6qW8nz1t17tUEDPmrP3ClnQjQa8
JzFV8IljltK38ffEABizKjIbfm5Flf3uKlSyvshloFjSV6Px+IMrVy+hsYMmpY5n
DLAMQNpkrt0eCIYbtkLKQsTqIsFef7qoxIPwC/bFdd0lcU6lRtbOf51Y25y3ZFtC
DlmYok6xU43UATAzk4o6jTnKe/AwwV3IuJulsi0SDmq5QTMh+3QDIxJyyYauzvkz
r8lMw5JHYIDtYIeR8T3Acy3gMZMW3vvmuWdl03msptZNLB6Iw3bNcAjkmZf2OeLW
UmzsvSM0/FdoyMxSIdvgWKL1TXjvP2MUChEPVXRVb+N+YIog6cq6aceL2YrsFuUf
JyEj7bgbhKwE2wLZKqGwRkyOgca8rspTe+Vz4Sg5FC0G95nMlm5qaP4tPjLGSND3
DGGlPhi/jfgWvaYpaK7fvbGf1fqRX9ldytwxyiw1ljZv7W9kWBHCmNljrRWJuSNX
XEb/zFl03GtS8KnlCa+WZSztQoAuf/VgbKXDcGHdJmFPaJv2YAaPM/BB4iJbJOwt
U8KcJwIMCH0rvlh75DCcAeGTQORMIh8HqlKbgeh51yvodzmcib17j9Dqaf1Dt/ZC
WnXDHnG1wItZkoniF7+JuDnVv2crReGWrKEmQFzDFiVDk7arIopPmeG7Wgt5mJUB
B7I9XXaaNnjCirZ7Q1O8mJUx0iY174vVJzXrQ7ultt2l0xg2G0I9llkNjDJIj2Yp
cHmrSik0bmCFO7mEJel8X9a3FnDLU34liY9KW57J/7vOcW5VXebA6eQh1iBRd0nX
pXGKOJL8teIgbZVDgJNDnPnR36pYt9f6PBeP2+gK4Qa7dktIw174PRDeDNbJqwJ9
mUkReNmjPtBYyIXCydJmhS3NQlLPTGZx50VbTfI3rqb9pJCUk758/n/Mn14rks1d
n1s/l2Ir9zEm94kCYyY69Ui+Mo48/ywLk3MdiM48jm+F+9N3IRwAKWM1S3w1BB8G
grrdr+9hjMZ77fniDCMz4U8gKOJNg4Zy74NxT/aG0o2nXA0YbNhh8xM4XlIu1+VK
Gr/WxzN8dMXDd89V27yoR3Vg4s8mSGcJSYhAnfQ0v4aaZockUajBAcOGtOmftkTS
9RgFoTlFpHRc/rRsE7CsoCN6fKFASIE3QQrdLGvY+friOY8PEVqNAK2mUTPpZ9dj
wvYA9YH5G1N85WCVfw+/Mrmxc+XP55VtSMZzmUwXsNxnklezKybxQFlr0TiXgzBF
O/7UnFizI7RKz/VLHyqJ2O/7Y8BVO1RvpRO9a2plFs5ib9dEXBabDpYDM9vxFKbw
ZIwEUAgbrKEZ97lNuLDLDtpxCDONVbFgVOx1lW0SRrLB6+z0MlMPjeVw5TBDjhio
5nhmTdNPIW0OFEG4uH/Vf+ob2v4XVmzTfaOxbpRu4V4NDNdw4XUR42I/ioghkESI
R5+eXiB6Ar/AjyQCFIWwfoxyZmQ239bcCsHXNS8dJM+R4/ny+9bVmWd0QZDPT39h
Eo8XLaTvx1se3k5/faqcl86IGAPfsXtC2tCIMK0NpxcyIi57n4CasnfWul/j+6nZ
LgbwQ/74GZXNr5eFEVM4wytWcfR7Y2HNbTKrWFpZYUJPLLC6MOS4EqXnJlGLR2Tc
CBc6DGppRWKEFkA7YAKJiS1AyhMpYnX1/IDRDQqo9zxGy/6H9NBJAkjiYKxaUjvB
ySswrehKziNC3So8zLR637av9RvNVbdyzxZd1L2eV9A0XW8taf8kfmSO+21cRNkn
8UrxtHCwnJIVo2OiXkPfZwUSVCnfG+0JSJKSN3voHF82uqiZx46OT/nwHixZMeW4
wMLtuCxPWUFp5F+q3/B+rasXxy0ymurQ1mdjjVU/S/QSZobzsUFzWR+9qil3MqZC
2pfJgwFOjKKGCBa0x4lu2PgVCwHQttqKqTMAQ7l91gFd6QTttXh4giVH896mD/Yb
03mKDtQ/NW2/7ibYd437hxEDVAQ2dJcc2HEeUq+rXygtj/erCvRMhXtDnzmG3E5c
q6JGmzhREkAtSJrbmeAXdEFiZY8lXrv8QwYwyHWt46B9Tcuo7PndsuWzE73yoSnp
9ldXm7n6kdHtrq0J168HXoHsZfwlFKPgO/frKlDXlO9MTFWrY/J2OdoegrxORZB7
BE3AH/K9XFRa8ZbBkG/7+TznpCeG9iXIVlPnEseX0VJ6LhvCF/od4vpxt0MmeVCx
/9R+Q3ENH4hI2kC+10kbI+p1453Cmu3uJss9Y6he7XsMkAYmc96Onht08V5QjcJk
9DMShb8A/56z0kKv9OPbvFOwYwehjuDE1OIbeHMn8P9RzPBpaeY0QuNcJ+JnRVWf
iMDOYS+J3gPEtWRD76I/xVQ5CKjO2Uzp7QYDzkEb3vcLsQS55bduHo38lofh7mly
T1SUPXDNjc8150acv7OGKFmqC7Sw87MUlNdGHUmcXrZUbQx8B3TftKDdGiibcZc4
tw7bHNxwR5xdD9S0GS1x8RQK/b7MOdMclNaLGJPzQlZT7dbxfmWGxkHue153aYeM
rVyHj4QoMyANPGS+g74fxOtFBjzmC/ElRF+uktaCVTXOe4wwCmKVC48fSyAmys6c
GjrM6etW18IJW0/J2qiJlhIX05pq4HkvlbNF8+gJvyQNMD1G1TBLk4SGkBT4XwLV
N/b1b69825zI6UEziZl9w3guC6mrH0dPfSdt5wpwa63ke6oH5kMzHZaxNn6NCMWw
XTYlPqddbs1ZWPJnyKLCfbZELD3Tr/kbkOEzpyYSz3n9MAQZxpa5Cc7MrgV8hnyj
FDdChY3zDP4jgF7rFO0kWfE7Z0g0Aef++QQopiWO+fFkTYd/zkDjHrsqMHK20Asm
tyzc5uUQ46YzalJ52gQuxsfzM2ofh9MMqmeXFxmjK/7aOfwbyq1jm9MO0IHjc0x2
g3jHboJH38IEPLssU96ypIjud9ptpCsLZ/n9xPqwreD+OI57CDo6Rbz6VffRYbKs
5rF3eK1cGvZtD850eaeKU6q801k5WgKSDtwATkPcCjrnXrdvm5fl6/5u8Y2IMEth
c05LnzopFivD/mx3N19ZO4lH1rJ4vWcfNFv/F2Fo5XswZ00JsLO/vy1Wy886kNgp
ByDmiecn7gDid2YtqboZko+Gz56zLnouiIxWkkVUc2ASZ8fcE98khWDXy4SPEr2S
S30l5weCM1HsayDlazEWNAHN4Fi9lC6q8wAY7L+Y7rUCpcr//iSGEM6OtmWUFEju
SVVD6t6ujcUlWtB6ye0coeX0zanFMDS1Vn+cQinXn5tUZMyNRJTLlb21b2FyHmI4
PjJaAM/uILma6G1m72MGXMBq2KchrSa0M1bMGOOJ0MVIHSeSHx4oDXdthCKhfSgT
3End+VvhHQWY1lAthClSff1F3hpA4egY94DlZu2a3JLpq+77eYvVxoTaPnLX+Uge
SbRklo/w4JGbuwT4hkONiRK1Zr5Samp6I80aEG9j1OHBZVkOGq6yP6cyQR8izIjQ
czrfMGG2ui0e+5RaNbXEFcSUZpbYfIxVyhX4TyS762l1EcN5+ExoacTTgNFAloVN
eODaX9OEAJt3xS+JJXPT4E3cApJ2N4g0/G3L7jUVCn6oy+KDdH8Q6dLTuGhVOw83
E3u8L99Av1i7c8HkmN90axBTqWSAoy9pI3uffoZOse60BQQsdWNwMvMpLMD8ilqn
Gk0uypgvo0mxNar556XrFAFMSmtIUDbqhOx3MPF9h7u9smp0RJlnGBANkhc+CV6t
spsoHT7zl9KGDQf3DDXiU+zlhcHPMPCy+n8QtqhDfGwXNeoDZIPnV7jcQDOIHzj+
uSV7PO9Ic1IEJeOm0IJVHlzMsB+LM2KJlqrhiIfL/RdleQHWcrcEmUE7MzbPNk4M
e5SGGxfN8Y5sXM3VCyLiW1+XMmLeBAOWeuuHXe9rBllUzNJqwaIourVtQlxxwvDj
QGDbgQHLnD3Ghz08y2LRcbFDr55GtH9gxFo2MTfdN+1z0++SmIOlKt2A8W9wMhS6
81U3W4v0rwDcCEe2isJsza8KsM4CSWFXf2vsAuUG9Bn451rLr9MTVRuuB6mLQ8KK
rRLnngab7FS4CNnRua4Nd3YcIcX12OiTRf9kOkCmNLSiTeOlV+Wq86jcKT2TGHeh
Pfvc6lm0GA+3MzucrJs2CfhIKigyCNr9mypJ+yS1WrGniHePlA30bPiUjrtgAXhA
ROPTFpR9ritcsithZnew6HSm0dCqF13B2Q71AXsQFCwgQxYVVsF5YqUVxp1+0bkn
4znJi9+zRXBk5GbksEDbAf8fHw5LNt67kzJIU88lZPUrQPWS/OqOMzWAJzG2geIW
6xOP7qml5hKqlC2n/ypPGdFraJlOY68qiW/jH+YkJHPp0mjgBFUdkdc0piLcGr6d
KSq2ORObLUmxCc8YzC+dCfRJe6bZsrlvrIvxhOekHfuaxKuDGN1JHZcomCK+1PlR
LdZSFsBFkW/37FvgUxrmqmRWQOzbqH5xn/phdIGeyyyR7BjnWQeVOhEDc7wcknHl
2L300/8ScwjRGww2Egm3PPdAYLSLndmfr8CH9uAaEgOozX4kjbEmSKUX4N+pHFp9
EKt9+xItI1ouSJS89umxs+wG0gi2Cmu69sy07sv6YgFjrKFfpeHKRWvmzDGhh0Hc
Q4/IGUp+B+5u5o2A3DVOkwQBFG3B1jhazLUznaUXIQnpPaE17oYtNnrfglHMl3Y/
qY2pSYC+JaG1a4Plts1ITRiv0XyO2CvWMALh0qnpIJ8bxtm2fIFFYF5PLTEyU7uw
iyhAZbRfn73QNMXcR9ueprBbY259StYV2JPT0g2esVFXgimZ+Hfbc+GML9BfWo0L
kgZPe5bZMhSF3AqGK4Tb683IBQK6WwDOytBriKc8eFwx/kQ7wQ94cNPaKwXP2jB3
gINaQpPC/6MkWPOHcKGI90ZeE0FJHl6Kvvk49C1pCr8twaGrP4MpP5+Jy0rkzkoY
8fLHk0yyBfYv+Dw7idURflO7/rxuLNDeuUY0lFpWjuR38arjZl92M9LWa6LurwzL
ET+ZddOUAZV3Urimtw4jpZa/KCYYjM5yys+mzZ2v6GehKSw4V/APCIInHqN30ARs
Wii6aJQjDIOuDgLQsgb6Yd/o738QlsPIs65DlIHn1Qq7vSASx4ml/kV4FLdhoX/1
nVT+Nhnx/Gd5d6S7g6R4uzj6/fFGGs3ktyF0LT46HdDTtoeuevmritOHnPy5PzLt
rPtOO+6cImW6yCcGk9wGnIuYK0vdopETZoVrDB4gn0KCY/jzPQUQrWbQDCULiFq5
j0tDUWJukeWYv8HB4PYwkX+pXpnkv0JxF2yyWyy+jdBQ0esc/Fy18k/6h669dRJz
+XrLNNeCSbukTM6efh9CTgJ536CHPe3dmznjFotzvVaDi7qRoBGZRKNVCZZ1xEy1
RmhCzuuwYgMzpBxPGyuEgAjZ+8bL8KPFZsr9ODnTjAOr5Tb94t1aKLufO+gW86HZ
dAo4C3jVoGhJRk05NCxyp2j2hL5Eskq8xZ70oMWRCD91kg/AV+kvi29ZAOl1pACV
6RnOXqNfq8ZOre0Kukx3LZvrxjYi+hUKNMr4RNiwMjt6YrejK7QmVKI7UCCmRp3q
rmB4h2jds7JEYJzUuYLsmEpMEJ3C06fBVLhO8SITHIyH3EwjLZ08xhmg+o3MHf1Y
UV9eN+ir2erh7kzxxJGGov2kwoyv54bejY+lYK+ya+wmPyxVxRztY5j9GTWN2EVt
CfaVvhkoIzTsPulOAtwdlCOnwhdWTNzQyM8zUNgPqRqSPV3+/5HPPliv60yVJMtM
gZysUMjDtyhjk+ZSGQuVNWPmWtsee/Z9/XbCyM/jiqExHYtJKE1P4V2fO9RIsRbE
yGwjGCFnXMpzynZlT+nBJFQN54IeCOYzIjnOOG4lFkFnIfytaG3wT//Qfkz3ngCG
mlXcwm4HCct5513eAsJrzHP6dXamPuavv5FeD+nuWT5co8nKpP7TGhWq68k/9G0b
a3KpKFTEiMcpbAej+QSasbwFN8mPa3gJ/TOthabSjKmwcQ029m2Rq0FY7V+cZ/TO
LSsiiUWafbhTr3KVdtzvpn4LI/UwooxgCBYNcAVbj2BKWOzMP0fVsq6t9BqYBalJ
x6smyjcgmeWnfgSNBiCW9wujbslRkfmCTitVwG/he1rspXdBQFzMVZ6o3pH0kEMr
6AMeWaK1XJE50RBaJ7gBiU3pjduZ0tsN5CBrjxHzKXqS1dCVC4O29Y1+1NK9TQES
Mx+DuACXI5+ntC76hf6RH0VQzdNUtFWTxcFwKsHsX0gcd7HhF1Nw5VvCdvdxRmmH
88fWeGZJAAKR36p/NixBvVcS/jBDn+0chDfRFF2dQFQGIPtpnjOyAZvblkRq/blc
7pXJJ/90V8Ax3sZ6PdkdSH5hFb7YImOQH1FyWJDo50wMO8cfvxMsDVguJYW3yPcJ
SSVQUSqSWFd5yRZlr+h8gtPknAQ37xSvYcbafufg2cV2MNR1UQ7MpGiZaLjUBErU
0pWXhF3QLRJ8gFHNIa7o1qwyI8N65J6nxdjMAyo476bxk+GTIqUAmS5PYdkEn8Zf
zdzZbNsKTf6gzx2q/uhss+MRinsUoKS9vLef8ukovHGZibQCksi9BWDiOg8XPPH1
77ORtNj4P7N/khxjYkxUH6jNThLbona69gnZ/fy1tcHP3DT4UAF4z9qYUP4GKsj3
OuRC5byTVYyPY6hsHchWrtfZBG4BgaMBwr5eCaAL0pvEOv2UUuoDvi/eF4Yf/Pld
80vGvuuHr3zELTAG9nkcgfpUKM7LjcnS1leR1ld4wl9sI8+REZMssMVQjlAoMbYT
2LsxzBLWyknYTKJPbL9FnMkTQrSSx3ovpameuz0gtDHHaIZGncpPKqcoo92KaZl7
FMWChoomf+UW3SGpEWF+tO+30JFiUCBNGwxhStjZZzblvnvTwaIxGGrzc3balhtd
4VK9zImV/wqO0+EJVZua9G7C5I2+WVmIXsk+BDh98q1xGxtSA5MjvIwKDjmFmaaS
yBd4weZzd8DY+KEO3yf+zLBWnHGXVumyGk7Yp3Sp+bYqn/c7S/JaI+F5IBKsg3YF
Fnyas8SlRXkatT+LtoVG+rpxwDI4zKm7DbZotc8WzBxBXMenOdXruHEnTSlCsJUG
2LwexTEbOzeIAGYhhCzrKDXv9xKIIpp+6Q694fZJVV1QiQVo36Jw5cLGSW9Z51hT
JXMATO/XxVQr290MQnNT5nx5bkrXTerxo77QJAYqyJ6mkQ8GVQSUQE0oDe/ovyaz
oBFmM62r9wyMzX676ljGbcEof+pXBAtIeRbyyX2tWWYNVStYdmWKVfEDTPf+tq0d
zsGH5jkPE3gGPOrdgn7vG3tlYlMF/h5mwI9F7ImGCw6WCqidP3pYeFBoL92Cg9PK
u2TkTG8tLyhaKVQ13ckt4nktGdpHGJ6lL07afAgZq0rvGrZVUNK0VxmqneucdoM+
WSlSEb4cHAYjovD0XfA7Fp2AcoVMeI50JMdaLW60dQXfXT4kDY9jIb3T/rjRclpN
M3I1vpoJPH0cyyHD4c+pL58GdeQVxrr/GqPClYPUUQof8O9rKU9WSqDCfwAGpTUN
eBgTNDG19cOUdqi/Ct97Wcp86aj1IDq8My255LigAOY0pBNaziOQbmMHHPh/qB3X
NtqBpNsVsAJ+6K1byOjOZ4RRLdzhnako9zTkXhojvOWDBCg4RgCkG1zpN2Odxe4z
l0CDh3u2VSwXo7gDu79ldYLZhoHdPRsJwoe63lbXYyOwY5pq/U2KkwUN4E8AKXh5
RmMg9B50XGHR8EEy9eqC92t5pSuK4DG5EyqrFZnNBe5oHorwcaTe6a1/ad7sH+Nc
R9cRthbppU/AEgmU6UXS6yPrd6tj5RlVNu/+wibXh82++maB8quzqNA549A5Feeu
1Q9sL8g1O/DjGtJ4RooPNsFIFiJ4vnU11aQpw24zosXN10eizH43/KQRrBpeBA1d
ALPUl7zrpz2WWQbNCXQcVlndiqekcbNTwgjekDv04P2Ob94s/J3LHoNRMBKMK094
FEOxZzBxzbajoCbs63aKGCPyK79xDBPhHCwOikS1v3dZqQTL6zMk/7zNvy9mTP1z
XTv/Y0bVLZacqW9jiU9b7HyVpJ2+XxhtadnSNxv1XcL4SbchR9BMcw8yjc8zPKuB
xi9etfR+RIyJZu60Gqd2AEArASMubj/lTkwppdiO2WiQ87mR2m3d9h3sSMm2GltZ
jOP7ErWlPsALO9DVd6z42Xtlr7LM6yJ+xHYx6Vl02SdTX46uthDCohWq3anMC05Z
3f0VXxQq/9S7Yzu2o3ru3fkmdAaAY5YQ9zrl8fbeEswSrihVZgzqp6MkTYh3oL3K
B1Gr1lE/4RxiaCgbeL1muFEfGGeVkU8LEEsMDWpBC6hCwmLGl91EbtikUfEGK9Ud
kRXOuS+tmbp+qBhsnzdyXaiWnCUO0q0gkB3y5Z5tMsdvNRNX4sPRFkTOT9oNQSAU
GLKAqEfk6T4Dlii9THaLgRQZTtrK8/R2/mphT65KOq5GLPRRmpdgiMLMJ0gKbC9G
5HqJ/3traxK9EYBsOEUAh+4IBTe54LBQiyHBK2gzFUX6zTRIYtn69PdCiRZPZ1MA
UR3VODcJAxZvv7KYkJjuC8hUELslO/D4XalBRG6WvF/JyYbE0UDReekdyl0W1PNl
bfaRldovz0ZXsjcefAaCVbD46CX6/fcJMO3IDRsdJg0zkCWgEOJEyEiOSNkvw0JN
V/13xALI7sbCwU+B1K5e/4nTHAaZ13YEEX5EBYFJ0QESaLJfRPadze28qBvvzrxc
cJB+t9QIzIHOwXroc1ND7yl3LG+arv6RWmSrhchYrlAucg3SdHT2jq6JHVv7BwYV
NkVAP7CF//q3ILwhZLLgdfWAo0lhGp2W8fCOjFFoYkS6T6kAwojFdFl/Ps9Rr8/L
2qIOEMGxYyuuE+G829hFPQ79FspRidGBtYyUOokgdaIVrF/7CGDVoGKbI3vbvPtu
2oHDZmmTNrBJ3PsB+q9f7gGx1JUAmeZxwFpqAi+QlrueGwgs58XjkXyN8b/3Ue2E
az9pFcdVG+/c/haEsPLz+vVtmNqtKStyQAoZmgz9U7QlZFQRMWgcu014Rw0GrNd+
8jimX9odT7Oz5Bi2xCHxrwxXjxNdAt+AA8z3l0pBN9ik99DIX5BtsHbWIEeJlAip
0TMBwqtbPWVsmEbpkgHWX0GXFBI0MtVhtCsGW6EMQyCBpbYh2qD96/Tqs5UM6hVy
1a++qmqHMKUPHOzlbV718xTsp06+sDJ6oozy777qamrMJIeyVrd7b2nOxhsvviPz
Y8DC4LCur7dqUXlTJNDgCEiM7q9YVUjIrE83Fzfvjernq1xaARk+OrOV8uErAe6u
M8Cv7DqNhYVi15yYKrF7Z1rfrB0O7js1DH0UdTcwV41LVH5RgOkGTpMTZv7R1JlN
DIQdFFTBPm07x1UCAhyB1qZVNQYiFm6KUkpw94dvgI2QfoQ49I/VuVhio9JGU0y5
WlO5q6XyLYDRobywx+a9dEtnPiFEHCft8CYxIPQQs2Y/3wDuLDlnU2MCei/DdV9P
XJc1Fd3sa6DiQQABRdfhQbBOgxYyqFXQkvYQnUfdQpAIpS9d6RIuVwhRIFmH7GLH
tKhwQFOhl66FCA5Xa6u2jjb89Pv+4Oh5UYKl6IlEw4KGogQCiZUXdkhHr9B2kkLC
Ju+W9AqbZu0w8MXAnJlGuFjnfBlz1mQpkHioy8BVKuRiV5MngA5plX+FsqUheFVI
FRDKs6qjvD4F6PfdX9bPPQSLaHWDcGCORQRa398oe6m8eCEvaoVfT7HU1Yq8lnGu
JtuodGqh9QB/aUBMw05LyZd4PWu5FxoxX8g04PGJ1T8SLhfSieg4lKkjI6NiiAbw
yOEn/H/d99sIYDDO8WWxfZ/O0Jk3lId3LzJwVfAbhfBAMouZzTFrS2t0eezg0SLI
wIIxRzx7VqqZbxXuWHsOiEL3j1wsNbgRvFFaqBwn+BTWdAnUb0tz8D7LgDUUqRRR
oyApX2FXXQoIaZtiW5BEbjpnY94NugWUIU5NEYqlPqMCnq4UdP/Qlrq3PGttaq90
lw/PPoWVKGkNB+7nPsO5ZZSqPiEhh4oDLxg0ErMsTgM5eS+nIIiWnvNPudj3KPrK
42ZXNMIq25cQ12LoCA+S2gD1njbKtbEu8FAYCTvge5+BR8W21WShsawuSCxb7AFK
4WlrdMwREr4zt+QYdX2CS4wzoArnnJAzoBQo7SpIG2JpvDZuVJKnZQ904mf3N6gW
5NU6tPBtXsBuDWC/4uCyvDpY1VfdFb064Lbj5CJagxlk04ebGdpMmuWyg3JeZVay
hBwQ6vUfKGuvcKcmdihsYopRVeOnShC1yqhZ9pl2l5x8Mc8rclj7AgjEH0CVgkM/
QArhCNzD6WG6ipKLEego8kFfpOUXZ8C/pWSP031de7M9fk00CD9NFNpHEnB+baCd
6WvDoMgn+hrfJnDW97WGqfTQ496i6q+BiCdY6Wfy1tVZeoShgrNqIUn+BV3yLBmV
Or8fYiUd8/RtAQGK3phVL+S+V7Oi2RHtvnMjBbdWLRivV0YrG7sghnQGQrcZCMyQ
2IxUXj8NElc5ZkSczsbj0zxld/pn/sYXXHWPDpk5N/CnqyslPRwP3ZnqYnTaAe3f
3wfs09fXZ342EL1dX1jBIbTyQDKBlhqzM0Ps3SIeXqQfAb8lvoXBtA17FpKW/F0T
nLTC777jM8+dIZucO9LM9vf3O2L7Wp+rxgwuS7NHKXt61Yw984PUuSiza2nIr6k7
qpkHKZj63bCarZd2ORdD4/+ZnCgAmNAU3tiIo60JmW8eQ2U6eJ8mjhgi/NNMi2o7
GcSfrguas+zFDrbLyV6tnt2sywuk+V7QGPdqeD8kagTDrXZx26JmwIVvlWLOmdrv
nxtfoVvOwlvfHBedDUeQoGiQFRb6gK75To95HWJ8yBISQVohxJOd754wV5Ry+nKe
jMWbS9SuS468B6XyI9XATK1hjyv04Jf1gN7dhdujIW0Nq6VYVU4o+4PXRVYFc+Tj
iWSARX5S+em7TkzOyPWGTZvjsA0gqxctKDSH+GQTOjD5WTv6+8gZl3Rw6kvp3PQ7
cujEJJLbYrpKt8VXcOX7MMl7iB6V480MLXtPCoK8XrAGuOi+g3bN4+qFTyvEMYt7
Gc5vGfqstYF5kxbvnK6/MIg1CITCGwcA7SK3+gOka0zaRx44bxkVOwt0aG5JcsUm
ms3r8DiLUctd/8Ibl5NsxJTcV1UnM1etL+uxCuxnHuBKzicDPSeghnHAzwHb2BQk
gUzjcGCWBtsohVDB4Yj8DYd0AzIkRRDj9nM8hb0K+IVY5Ksj87W0RSHkrV2EFcfm
uivgyqGVRLp60pWi1BG0iGUWYQDB/m+gj5h88trDb49wYHGbOfsdOsQ6evuI7SdD
oxkkIx1L8nO3jpEJPIe/thvq7lstFyfz3DTGmHy2Y1wnPUl7wRlU2ddhFWPhg4Gn
S1g+LKJ1KwxV58kC6vNlyqKaCjrHaVkccb5V4OMR1yofJV3sJTUeTGrVFBhREDr2
ciAe5rmdhe7PkkJ0uxtZ/CC3VP4/G1vyvyo50sSzn7MSYLq3EE+bJ1hgqdqTpYfD
C7bGmFbnkY+EyVVKBnTx4ulh+MF699WD6g1PEkBnxwGrcGgUTqHXELDD7knBlGk2
W9I8YI8JRn2l8WZrjbZQzURnuSevkntMcUF8tyRDMVXjPVi2As8RbJAql5HzSz4A
qmzLzNrY037CvmFvOHiuEL6cp4uSSKi2Tom/+Z42omHRfrtoGFQ0o4+TUd1GTZL9
e3ehzH/Qrv7k02UzbdJFwBj5sdbuMiQ+Vu1PahfGvHJ0MlPVbIbgjXCV2ggds36f
zRmn0wVz9voRnAf67IJhHOdEQEYwI4RUQmGcKYAWtjEL3qP1mgxjKta+DAwkzXyi
n1NTXZvcS8hcRpU7eXP86fdSVhL91q4P+EszPBCccUvNGX/VfTB3zS5cHefBW1QI
7t/bFtaAk4LzspxmiTBDfUroATxXEtQuiBWdRrrmDuyaoFr4mUm5WRgaCcZyKSFv
ktvNrDOLrELNo5lRaZL4b/hEBTkPx7OaPkwcP5D4T0hvtnbek9h2mFk4VAMsbvYx
ZJLdHE1TrWu6q5Z04WPP8Kx5RTB88zL4Nxwt6cR7qxqM6uXeSK9a1nsNdzL6SS7x
EXQrURT31VBDrN/XdE/gSA+wkrveJ4/FFSIolwQXZZuB+yycVd0yzKr/pVZ9s20R
8WBEC2P6AA3s49LZ/Csccv+e7oJVoRNeI9G2sau8Rr9fusf1ZOo4tlU35A1QVMqT
dN/aztu1rA7IVdV53IxntvoXQxINdB6+ZFpfUkIrwXLizVGcrlFsmMB+TGaKyfur
eghxAzG2H92TdOqnoZQMPzCqCbLL8Agwuuid2OrM0fWA/0eBX4tOr0iFGCKYEG2G
EjQ+xRZ7xhAokUIiXALymvvUJimJwKS00NIKgG25h/2mZd6baXO9TK9m1dLSCVsI
gLuWTPYtIu77PGNfuHBBdnrkY5HaJXft03sI7yNu5774IX3hL9nGtYw+M4zPQfct
hUVWE1NnfAMDgb0NO4/0BO8zahjIUMgcLsYvpa+SY4bmThz6S4GywvYhyV9sVFuM
YwSWwQf8X4/oaB1I8xtYpgUOkA5hNuj62lVmBJBHEZ9F1+mr8x3XZaIk3QoqIX7B
3XXEJS5qM9EtPeIVVI2UDWh0OfleC5ppFPVoiTFSCs7UsPysTNQH7j97robSOzc8
bYjhlfSnDNMCaoBSMRhu5dYqVO5lnGVn07fJiuMla/mMw/s5Hp3SsBWw00vS4Tc1
qOxfijxJltAkyTl63HeOt+mZhTuS3Ao0gTFKpuxTb1vtItx4kjiWOz2DUGNm9neB
rsgbg+vt1gh2IbN410mqvHnA96YKI/2RRLUERUF2JNyE6OVnsEoKoUyYkn6jIofB
yCwdLyTLSKn3UZVGR+iKWMjAd+UH/e12Ok9rfYLMxu2h9HLfuXGJmgm3kBDSdRHn
dL+KGHccwJH+WxvLqWuzAftK2OEi5dgf8tNL1bpEFgODtFHmrLVxxVikoHMRV46t
SxB+sUNAQzUoeXN3VQy6o+3LX7rqcIbS2vnMrWFTaqj4O/N1/inlO3p96Kmd8ho8
DR36HSG0bZH3rsKjtFU7TjhqyDH4t5bBOmKexm56eEhARaTF2cFbOO8KnzwaYM52
PEMyydx1T7UU8xgYZJ1F+zxgtPG4HNw2ONGscOIaz2dGvbuKumKzKx4SPw3zctGv
lB8g9b4ctpjWWl78kci9JAW2VaaOhsyGcYMCFa+Tf//AFu7VfWlauFdCPgFWE8FZ
zBylXplbfsvvYQ5eshFTA2eiESLA0ms7ADsncaciCNHjOtApLOfR5ahINIceaOWi
PW8CbTvIAtP7Epl3KtcaCdXCsSdoIjZx1UAtbYlnvQyHYVIIXl4v7oY8dIijUNQE
qyMRWxMEMzSvexzReSKl4qG1lzjtcQvOyuqKLfaOPKECS0QT4sdH48HJbIzahwZh
mVIKoeeoj7d9XM0TLZIk1Mw5f4sDuMou5A3ppvfUCeKiU9DYsEpJ/B0hIedft9hG
iqXI3fKXFZCi9+KhePuqKupCFG/GgbixaGIwf86uIN3JT5chC29ARtttVAQRB+wj
SHm2U6S2R7NmDAUL/THsYogf6yAQPDcfOkB/ysVm6XlQxIDxGteD7T8kLbcWm+i8
bIR+y4dggNDp6XP9pR87X52Gbp1CvPsGMpZpzH9ti3kAU3GGomvwavRh+qApFzTu
byxlNPZUXjcMd0SKsL8LNce37kj834DLUlswoKFjefADj5Y0okGwh6VJhHvFwvxT
wEabd9sNH2eneaKQm1ubV7H45AKSsH1FFOV6cOyTHq88WysEDVHAsBk+dM+6uck4
ZqijQHvw5FyDKCRecm4tqnC3EXJJlmUt0RzwX2epaO9+5TynihYDxXxlRCk6iZ00
3jj+YkYI+JJAvQB/nAml4K2u5ozUzDxQ/yWwsu53tmyqsOlF7WNbYVsOJ91OB0OO
1Ml4zOeDGiS2EEyooBIbX8IJkO72BiwHoU6OcKtGk46FlwsQv3Lzy/xYeNVZJHNh
pwTZWpRlpin80jLlihz3qB19R0VEtaDnmKOX+fMOHJxMsNw2TUN1TfXBSrL4CndZ
R2bDYDlbmBvilfOUrj5Rrmnx/oJvDeOgkUybSmniFhZv+ct8l8x60U65Tcdaudml
PryzbCNphtaRYYYp9fk7egOFkPVI8ozWMWVTtO5rNozTRhQyG4OzxpLipbwmB5QO
NDbgu3rdeoQlzkRJye2gy0K5WxIgLKW0vFUAqMEkJJzbUmE3AWcVYgAIalomtigB
UunkbNiuAUHE7VWE08FPxiTE6Letm5jQ06E4I7V1PgtfP0oWNuO+bcv7RVK+5Y6U
bGV6xhuB/T3j+ysk6XnGDC7EInaxze/bvdOTnM0IvzP+ssr247ZrnQ3Rlq7Cdj51
TSNQ6HuV6I4huDbocvjVPo3hJEouJknkP/hNniD9sj4Zwo10SLRkTn5uHRH8xXAH
vgZaF+UTvhTYgLnQOXGlgY4A622UZXN4XEp+AtbKZvMWrCKGJ/LHiAySl1UqXc6J
K2P9i2Voe9CkjssqoLRuVsVJkP00A84E6NlLHptTzNQcjU2u87LvHY+an8TPF6aY
XKLPe+4u9hSf5TKLD3iXUzDtztYerPM1Cle/cYFcJqMyW9YgAItL4Jh24GR2Y+tz
TA+ZsTFo2csJyijbi78KdQBKcqbHGT0P9V0LCVjfbwLGptX9C8fRgr14H0uFq9zx
CQr7q1Oznay4GZ4o81sY82fFRIGAmtDtFk8bjY/mfxVcfuiL3RiEENYpPTiVitph
2AuLMSTZxjp++e2Tbc8KWKU42sfZvF7bteautmxn6ittbp4IdnXVs3QP6YExCuOD
SCZjjUpQ7KBkwGOoCyszNDl9LMVstnLAZfs7rXP7cfWu232EW+rhb/BCix5y7lYm
/tboaVARn7MTgwvPiBLqErPujQHmGKSzF9LgxvHUFHDRR4S4C7YLSCnLqE6Vgem8
R0YyoRW18GPRkxO6Ea/1uLjoi+8kQ66KYMWXhLBad72jwG0/SwfLKStMGIXL29WP
LiFsuZWrXglooKtPJwgRKgkLOUWGECN7S5cwI0S19bZ0G4v5KRcv+vGlc3hZd3gG
WtuJvXM1VoR39Tfi+g0QImbZs17WXpUVTHnz60qeq8MwoDbiUo/qNUKhxWIDqTHn
H5MkSPtrGfsGEEbA7mhjB4hLEjj0nCKFQZDC/+KeClIbOSjdW1L8zI1SRRLdCeU/
r4OxwlJaggALTUe53EBXFluwPfLOj41hSM3L54LNmrsyuql0ZKw+1W6+dA4+iSfv
PHUwQ6z6U/Mh47oJjJLEBGaCChtCzrtMvsajLMwVKYmhKJ0VxDZ7U+xZUY8cYwU5
4ikEEmn14YfM8m1CnSSUfGc8aZyN5vXyvYPXOgmCEsFB37rV37fopH2IF5cBbfKy
GdCEBIYKYqR5vDIisC9SIMq41E4Cl9X9GneKr7nwk6qBfT14TiysagHys6dhAWTp
ockaz4ZlUhJu5ZpGhMXB6noTJuAXO2SHoENSxZMnv+E99y+C71uRwAewAYVOjZUq
sBXBl7SZ+z4Ga9KefUBbcoCXmEu2jcjcUHFwoBmweYi2DLpvOIX+vCocU2Dz2pZZ
k7QriEEdSk+vMo0T6GHov2NRoouMCqhuksojzdMtTrgHoBcgABk5IhzuObKnsuR2
qm1AaS/WitrkxVm1D7F0PJZy1ZkW0OsSSv/3hIsJvSkK68aLsPYlfeT65eML6kxv
N99J6RQRSTjXkMdwYJbBue6y7oliTJaHwSyLfSDA9hgkkJTXam6UfGAZKozGZb4P
7QhSNyuOCU2UJvatZp9CScSgFqBQZ2NJb0QtJ2l3xFIXPuk8oTKyqzEon7ix3UDP
Geigq7rOKOUbS40XVzh0gkQziryRYQtzMFHwlyv7XivXUKSWMjqhlAO50wCa8/2s
LjzG7blmpjbPR9mpE0R5QeCTrM5cu+XjYYqKYGfOJLt8vPqDKc4IAmK2Ieihds77
L+YS0k4dnjryrWe6gEMT55gFXjb2IsgAxEfQiqRLtz1VxVXilmewQ8+I9MX27YmY
Q5XP9nBX6VE5RoEa+TIGO4+iIuv5IGeYcaaJke2HCe/R8PYhgNnHo15fOKGw/0Zw
c6JCDK9HfsXalEHg/DjTrlqXHcUvYUdwqh0OZE4RsNHWpROL8rx94U/HBUv2Pmri
BwJQ3rVZjc3sx6P/4EzN/LQN8tS+bQv5HxLMDbeAgNbRVKufqIE7Uwc/2rdlt7NF
0ktohzm8qOXdTdgJM9dxcOfhCMo9xvquI2lrhlurF/MTqmhWWMcrnJcJmj0ALGf9
hyj+b/nCZbhoXW/tHIa9fm2+Y3lrqbFSy6SO8Z5Fo1tDQ+6hsTX/jkavhIVpRW7I
RKFfGeFw+LDBOSPe+SgauVTM4+GTEZJdfY6/+IhfcOqEaTyQfdGOqbbPtyTH3np8
iM91LvTtwA+9fpSQz8obBnQXxZIf/kq5oH0OlHUKfEWwYuxA76njpiS/dy6swwsF
KSCF2FnR/mp/YUx+/lSAYR5o200pi6mzD81pmliR+sC/KkB25vmpvU7t+FsZaNet
CPdNnlVVl5DYBzCx/ZwsOJZUwQwxRSEZ/U2uIe4xLK9zQqDxWpZkImTIqsb11MG/
EUhjP1miWfN1phljplMcefOoSQa6BB5K/HH0izEag9xqkolJu6dTBOzR2x/XZEZT
BXtB0S8eIljNS54spJG3/D6KKVmZI2gAOfy2R7O3u1FgBtDPIe1ApqU6jr6OysiK
KoKDCcyV8XCXehY7a/gqbIW4/xz74dZ4eRfRlXlDbEyMCsslh+Z6DQA7NJBslftn
2p3EtEV8SgK2/1JDYrF8cX9SUyQB6bJ2cCyW8h50S7iYmVFxH56poJTxC02e6ZD5
Vvhr6vawc+f8bgWaJJ0JP7xeZrMwiiOREq+S3I2tH+0s15pQRK/if9IBeDyXllA/
r8NKbE7HpH7iih6aLHZwqGnRxNh7rRTIcJN+VTh8wj54NWdLpgduq1GNCi3J2/+v
6fXGigukrkflDg5Sl+NT6BrlHKx9fShKUmwXf5ShFVa4qV+YFEolO/iWFpc+L9Ts
WSRFDckUAkmhOc4MC+sx6Bni4rdAopoXbBEmedbZe0gL/sKPAQEGbgmx1pu1tMmS
9vJkARN4GBZJxHYVCLV1kh8raxFfk7pjqK+I/fiCzhamlvVTaZE20ZA8YWMseQMr
4qNxZ/jzeLQ+WTSMLOlbqaldEtjf3EOyJ+w44gzqBcMhOmIJj3qa/clpzejPeUM6
WCsHfg93aKT3w/AMO37hhOA5EuXsEFpqzcVNOpmiymaYTzOx43ZN8glKydiCNAJe
kPOz+uZ9iKGMjfaCJG+cqpOOv8+M3jyPu7jJd48xPDFbhtHZ9q8HR7owoERtM4GK
Lewqlz23QRs4ttVAoZ6eCDh0MpmZHQbnn74lP5jBziIVwxph3efA2zBprVED54U7
k/tc+9xumGLfmd33WtvqmgELCwWRRY0J87kqDIhsyiqm9A0py1GNQJtfQPfzVL9v
+orposJ4CmSOzIeDtcrzDMo+81e1vJrunjIME6lb9p0reatQOirKwyHgHvTRD8w3
Q5dbXV1efHKq/amM+WQTICglIBsjWkKwuqvb0neO8ShOsPcgBqb0IDzKiBI3EAUl
C0br+35/XG76qzPYQHaqKLM4cFvIkGFmUzeM49tbJXZB1DOnF2JBkNAuOZHGoiTG
DK+nJWcmO3ReAELEWkAZNSmKbx4xl1Og1AYHbc93b8kEqkeFuzvNPX+ZCPSZj3rK
PcsIu9+aiPio80Bw/cgwpWz3hyW/SOsKl7NyCiMzRaWVpecCBrV+FNKpB2GhqCHG
oG+QleTGRDMPsJYuKTvV2pqR2o5S6TDB+YnleP2gNAD8uziMzxjXKYIHBe0N2huq
Ol/2wosc3C5VIjKh/mYk0gkVxZH+MgZ9SfL9jyUXYwi6bUjQ+PQhljIemLl63Glj
63dsnNai/Z7RHtS5Y8YO1YXjgKMxywJQZUAIDewnbO4BUwRWuwx6cIXSK6AXjTIv
Nar7Os2NE3ZC32kJwhn0uwjZ0JCGN0jGhEkKsJTv2t6ZWkqP6fu7f9I0HrLxv3/O
wXGt0+Xi9jtKcGTHQzgRMknoHytjn+ToJ4jO+GU5ezBjNgE3D4cgXw70eRDdIRW5
3Sm00L46YONWvWf+SGIjqcFnbBIzyXsGQymKtNKj5+98AUD20oyVduMcFLbqaWgF
3A7ILnWDpW/A2kop9Y9YgfCOajd/70UekD1rRO1rXeKpBMtCyhdGaG0fCq7BeGds
XJ80iGxJeREKrtAb4t5J+8W/kyLJeZjerv+A5zbkZw2+LfGdRGcYgNkF5CDyWFa/
y2w6Zpd3x6DKST9vDdgHFsNBELCNNvb39lVd47WlOLJoBSLizXU9DQCMkrjVRaAV
V183CvTAIfGyd8q4+WY0Ujot+4WnjXik7o1eb68BMLi5sg2WakzDcdm/8Rnhh1u1
AW3ogA8dKJZwBmX7PAiWv5jt9u7olrWM980uZ24YlhGn7yWyHaztOL194qFYV0Vx
waBGGVHfL9w7U3/fGdvoIoGMFpPJtjWHm2Foahcv0+j+TtAaA70m9PGFRaHjwQur
hx/Kr7406uQhIh2fuOIauBCg47g8DpxrxEbFzZLSM23eaMVvVXbDcE4T2Losh56l
XaHbta9u9l2mDz60Qhcm1SzWzfq0+9uCuJXiUkCS7NTsbUSr7Y4Fchl3ctKN2oE2
Pdtndj4xLxSRx5Q94Jnx0QfU9fTP9G6VNdMTa62u3tW1IYjqMRcOEUjZC4tMjHsn
+M3jzKu95kErwy6esvc+totCZM7m2l1Xl6ZWiwEcvDt3YHxO3Q7uo6kv92WybIWB
UsqkxiLVTkm7xOeT8NxZpJY8LRgkK6WoBvVya+k33IynOvNzEQAXPRoVUxalm1bZ
BHmStnS8QQxXuYIyFFLI50JRlhwvQkdKiIkjSa26EewuxteXXOe7RE8LRaJFBTPi
feO8So/gB6iJZTTHt7RPwovjSt/JE/hZTAkkKRpgZDaHK+lkaq3X6Jf6cHoVmoTZ
IKC57CYWSAOTFXiXecgKElUjbGbVia+zZf9Lx8Jyvqx1aiifnSHHkIKKQRq48MNW
7EUqZD+jOzmxQy/gWv77FKGIg6ul3BENamHSFT1Z5FBuKbPDIsA6bXSsv33QRmxH
ZESXlRU27MXFEOHWdg96F7Jy7NZvOLFxcISexWiJjBMhXxFpey04WCijb3tlJSl7
25GIOI3bf+/xsomoNjvk6kbjTqGc9sIebhv5emw85mwhht7a1RX+MWtcYZfiHHOq
HK34hAypPDlV4o/9TkorBzHywdRclG+1MFXbhnq79/dAaZlqtobyaPytF4dLG/Fe
KNDkhTx4NliSWmX1hEgvVchm1cYbaz6KgKD6YaLp6rstLlNzuxxKxySfUGgVb/zW
u7FISL5wz3pyBiY2YQtG0BhjmcHWbJOz+6+QX2HhMRuDsJDtTf7WSj56pdJGtKQ5
vUC3FESU69jwxWjqJeq4FXMzPoTf+rXXTCPpUzUJGzj1pAtxakXn7PBMeuCvLfVM
luNDQTIIPQvPWmN3n4TIp4HICfoi9HdcYBCVoCxN1YVda/szMai4Cv69RCAsVURZ
N9mwFN9SeM76xofwbmMtWJwDnOGhH+Yjgwbr5Wfr7jGHOuWUe/fps/bIx1AMH05c
dLBcq3Opi0dEd73qyvlisxZukMk5rCgliqX0cFgtvDaJ3mt8dP83ieq3XLI+bWHb
BVCOxQ5012SCIkMgU6bU7mHCAkD9HCcvDiq2jvYfT/eG6EZqyKyE78c4RTPgiQtH
+yR9BnPu8qwnAZ6re3So8bFs9eH48rh+xcEKQ9gf8eVQLMZqLotmePYyuq4kLB52
iQz5V/QzUzvnbBi/Yok9rA7BVUOsLCCctlakxQmcX4NF3r1IIF8sDQQyjIL6LUdQ
FbuJmQTSQyJA06qPVxDCaEkKsamazZG10zGNXb0KDn5dElyy3lzi9mNTzGcERFDP
zXagedSpS7blQAY3L5saekWpg7xpMnoTCNNWa/iEzYYKbAnFlemIrE4N4ZYckfbj
iwuYQboNJCCZL0DzCxGTDcG/jhi0srb8g5JOCXe7laC2E7w2WPtToQ+pASCstz0e
ClOo/BqZMm/fcGARn7Xy5VJ7IjaXHsgX78C2jP6jhenK3aN6tDwl+v6pPYpxRdaj
8TYv1CVYnUTDrH9bk00w90M8icWRhKSk+kgX50wORZMXC0EyPEcTGvYz88bRW3c5
gaNHFgrsmTiILt0FewS+QwGV+1PN22gd4MSzU1AJuc9XDnx2uniV9PD8u1mq9OCX
ZIJAROba3imN8vpsTNYFUVM87PSKA0vEYp6rhUC3S2LfnjOuyRf3iIJzuB1jxPql
h8hAf0bxavz+frbEM7GgHkPl7K3cFlSVgEbxRypElmMfO4crm2xbfPz4TgCwYEUb
E29iTNOe8p940WExtH48GPujKPR9C4YNy1h0P4X3IePSdC0sd3Wcb2CSclpe8cPR
D2fE18/PFJKSGn3ffRmwa0w9uQbhJzfgP8sqPq6e2Uzu8EqsWXvx4ChGOelssUZZ
bcmOVdpKHzvF0Vx14yhXkD9qmHWP2kZTD6XEongjhXtzQBu2QrP8Ujmq00c/WzhE
yrGVRCJoKV7azPaJKPPh9i+yt+mQ+AdlAxy+XPTkFlwcU3QgLnxbunpAn2hlc9Tw
fbxrNkflV/RuMt5Zj7qDY2iDulyB0jfCGJUrPcbwz0+uzmRI/fS5qYjaP0vpc/pz
oPMwF1PCZNfGSVcNkh6nDpQB9AWIH6IEjcPAvk99C9bO+XhvKAK2rGv7/0MDJbkX
vwt5iICAI0ksAglFZ+qlPB2EQv4Fs+C0usS1gUwT+rbD38lLlZN/CW4qMkZRm/6H
dHimqXgakxa08GOf2SmG3LkdoTrfgR0aRYy9jvA8yMQXe/+A8CsJmssKWUL29eQ8
iox9DRtpwn0ZejzBs37ZGvI2Iviw6Wijr+kwzeE5JOWrtlzLfmexGAaCL2IoDzAz
yezoDvORsbwGpqIPppAnDaKpvZlFt40R7qA720IecLYOVRBkwSHFYCc2WW3E2VaS
w6nnEcdpK3bYE3uN3RHctREo4eHxP7Kj4gkw5EPkCwsVuAZBalgJtvZS6x9dL17D
dIIWVqBl59sXrPotp5yGi3zSH7r+W03MzslhTek8nH4tcK+1/IGz6a3x3oDNFyp8
3vONMbJGWiAg51YfFaILXHjt/1JZFx4LnaRGNRo2ept1mgXcFVsplzIC2hGzvg/3
AbX3A7tHDYqN3VdzpgYVYIkiNV9pT+w9lSEOUdEleIZe43UVg4QrOta6/Wd/K5K4
mHKyNf42KruVQqAOyogUmoef40+ptAl9QGJDF7UmChP87FtXNAbwv6KPuiCjfSbp
xygYeyJcwUtCqZcx17bRql0CETaOfcxdi9AfElxI5LWIRFj6Rqzd33bfVnHFGsQM
ikw1U3TRQODMO+DFH0poEg7aaOX7rdgBYqEfD6ZmcPvviM6GWVMRRmtjKgtIs1hK
HvANCfS27RgePJYTTq5oFOKrKHChwgWaqUE5bFlw254I8ocDpBQlsDfTqZt9TCFq
c50df+Zqzq4dyD/yQde2+ZLJl+mSv6myn41q52QTJGbj+ryWg5QnN9r/CCycOmxS
2OEPXyNJMQ03KGsR08DtDjfJdjowNIL0iIS3hA287HkLQAsSWWXI56xx8VRYHCS3
brsojXIIDEFOUmin4EDIgNLS8qn7U/WphTcMBk2saWiyZPA+/LbbQSG2d/UAWKXa
NknWYHWCqRALdf8XYWRlwbEo1GN4eSdwDGznRsqpwuj3tXT20II8WCbKYNHyYPCg
vyR4RkQ3Pi5Oxg9nX9y5pvj/9zHSP7IBhueEOxNUSyPFP607r8D2w1VuEET019+G
p3SppweUQr3UYr3gWFNax62Bq1tv+RsdtKsZkEz0QQmHmScB3Zey2Xnt+gJzIf55
hJHRK2K5atgk8YCQcrRJ8UlWQ357sEX7r0cH+f8Le5jTA7bMtZRPejIp6OaJYYXN
fz81XiukFTNBzwhqDK28Ul0C5SYMRBdKXfgFjaI6dsn+T+f4hSSubP9ZmEh6/6lj
iPW67A6FQXW/8sRLglbFJg250sK2HkNeDJaGI/cF04F52qFJ79BiEd5ja8IppDeL
n3a79A9uOrnAwkS0/a/MsSLdwDVcgDwBlLdHmPhuc09Pq86HsNtTyJoK08jYk+AQ
vLDCMHFwlqikRq8ixSoNzHvhJNIUQcudknpdu62velYDh4GPDohdMuYjVyXOHLqo
/0HqusnCDYeEIfkhOfwo9F0TMoWapKpUiP6jARaPTEmoBKOnDuAeVltdtAK+ECZC
1QTBfHFCx+ngD/ixx4qnue8Tlh7a+aCFfJSbaxcaoj97ZO997f/fyTd32nWn6CZf
eT+vrO9szCKfqBUFSOT1MuTwoVBzBzP7WkQ2V5raQIO+f01GVDDW05gUjFmHfice
jQz0BrK/R7Jsrs1IUW2ZYV/EkUqmlaH2nrk6F7ZKNrX3mc8SkWDogUPypMErdTY9
hzmL3HyAcPnMTRj+/1RVtMw77rBVt3i478OQVFycfSFIFBR03oADA+Nu8uqaUBtR
IvKXFPFPK4EBnkXnpkVV4T5A0q6+CVkq9viNOIEZOubSlu9Z4PaFzxR/gASD7I94
o0xl54csQ7CVBVwcwISw3TJRgfMytVg5qRsMGzXoY191VHnZD5FwDkpFoq2ohWmm
N4aJxqz8BjxSVDbkkCYd5mB3ToTsmDxiQv1JyPkcoRDDdh5zsSa64SYBVOlI9W3i
H9UqouWG4NZW+aL8rk7gLwzdl+RAkAoY6ZRe3v+x5JkkHO2olfoJ3FQW3Y7OmTcP
79hSE/lbLadiqACrc+ffJiYwa3/FgaTLl5j7CEtSzd85g83a5mA8PL2jekrQNHgy
anRKacXncIiatdXoJzMseYDi7c9sAZ60lCe++q5v3ejrmsFwbpChVHKH1tgPjh1K
UBKEHy0dgGK4Jk7A23QiUdGNHgoLV6ECM0cIneL5kqetdtU8W9eXNzip1NWonccH
kprQHd+D6tMF28PskV6fY79xoP17xn2zMOooqg9yDalO01MxJOc8Iqbt9aWwSPDD
ao2JTyoMCEeGsGuEt3mCfdBQMEUuopp7S+oa8oKMX+4ffalsvlrjJLmU0FEcgj5a
XhuKOLQY2NH6v45sJjEFv7HF3vejn+tMZZSx6FIRzb/Ov4SE9k1wicWtBeK+NYzb
BwVtm20z2RyxbwBu5rJP8D6XiIiTjsQx6gMWfpjjrAZuaxwMKjTfs6NmLso9fJ6E
61D9I4GrSVvh5hWAnoNBtcPspoyQ/Ym3FDJbXm2w1xliZkZLFBWpClXzyQNEyryu
UU7hUrd6XpoBFH3BqyJI/Un8jt7RaXZmN1bhpVTZuiUgMf8ZbwPrJ3oVM2DsLBWE
/fLBBNkkzA27HJ1M5EVnn55E753DlZlnlW1EPBks/zN+csa1gxqfVSSb5LGnNlyK
00ZSRVB5xW6zaBWLShI7SALtaGBnNajlL0K6lGq06HJoBf+Zkn6TpVPJ7Fk5+l6s
qkOXcE2gOBFGc2uPTN0KyDk6CPlqUIjphZAFiEx2X2kDXl39kuNTyZtVcE1DRV6p
4Ncp5RsZXFO/0ubx4vOWS/sUYEtEAdibEzt7444OpKEwwJzuFECA+sw3msFmH5TL
VImkFycVepzJp2UB1lGegMrLzHJnzP/tTd9z9+6Wl5+4Z4C11/H5+7hG510A8XzW
8vB1oISSPILTUpoXrevuzFB69bf+GRcXuRUT6gpAWGtT2s9aboNiafAFIdvW3ELO
D+M7cLslS62qVHUSCEiDTZXg71QKNQ1qFMu4PZO17sZCKYDOLO+2Dk22KdwTqpVG
bDmclbUhHHybbnNqueh9yiwH6GGzJoNTdfjpl3Zuz0aPrLN/fItTzkpBVPnSsTN2
lPdNxufc09OK3syO1l3pv37oskIwoP43HFTLErYzhd2mywYqqWfN2mUcjfYU8zo2
UEzw+vbUytESsMN4863WiSv2aN9viVyLcDrTXimXqnGRJn6pUSqKbkRLEDGd21UE
/CZ9v6Vt3bEgkWuJfgspOJrc2sdsCWPFRLaPNgH0S88PoKvtLIHtPDO+wIBLKUyc
vyGqCGyNkydQEft2i8BD/5eoW5R7l5q79Be03l4rOMIdatbBkFtgN+/FsjxFC2Tw
Y3NS7g/9LZLSt5VHAAJ3NhvFiY3eg1hdBLLOMOSflnt7syJWCWY51mTDlaFiEUT4
OCa9BqswcvAHfUNSeXyyuw4NWsu4ev74m+OB9yxGt4SOCXg/ErTNJ+IhUa/PCnN+
rq/sNhGPvFBUQm5doEmiSYwNE/7tcxqEdI6f8GnMSHI79ldNr3Uw8GN1ptb7VjEB
AGfU5gm6FxxXvcyjEnJxbA9Rrjs1RtgFKTLvF3oJUTBWUyfa7CSEJlQyZZJuEp0M
VED/+hvQHWK1i8+ti7S5L59E5npwnJkHJkQvwOEESFMwb490Tcd8E4uVLcST0RJG
Ugx1TN3OecW8rHLPRKs02MMtgNtC9b865rgI2YIsA0oSpUeSepR5BgoyHoF2SWih
rXPEsutPIhApwIEXwMmZAJMoD48ZFOSEleb/zug0qB0lyuIg5nM59dlsJyiBvLJf
E9r/0V4c8aApl1WJ30gCTDWK+XaTCmf1tCz3GcJAAjzAXsnhKVJM2QoM6lh+qsIt
t+hdrmQruVHbd6g1gV0e6SLS34i4hno6Pc3V3bchCrvvkKJfmtuKD54cJvSEdmKE
aY97bGeYA/JbcXSP2PJYqh1crpcPNCRK5PP+r1BmMvIUczpOSXCWIoZeMk7srhps
F5n4wfLAdh8yB1DSTOlew23yIXxHAcBI58rJl4aAAss2S6H22KYeDGpIrUA5Zp/D
i5Aeff7YshE7qFW/P+l7kUwkwxngI6PHBWrOBKTKT0mb1nY8/p8CPjV2ynROdJp4
vdNRQPy5TqfHsPu5pJThGU2T/rVAUlobjdY2Q+/fS24DNPs2gxkqlYjdgJ2Hlj3y
YizZ0w4PRg7bqRFQkx+a9HTZRR6FPxhZSo8hAhOCxext+W67ofeG5Q0v2bDrmDjn
gsYseT8qqRTnfJfPOn2DuhSIf30K39AeDCZNZmzvctPkHBbNG1fDwrVIbypRx+Sv
RIRW+O5A/4svwejhmg8fvfocdpNahGBvN+ilzCWWIw0Y6BSbe3bTgQlag/EJROdM
8IfURgVMq50Kvi22NCe56vVU6f2WIdOwJdpUZDBLvPwuMoX8ZoIt6QtmPTFtaQF8
M+Z28gh9hYLnxGZnGa0gOXqqIDNp9RrpCzFIvLtD+KL7RkzlF5utZiqod74Sj/wB
Eko+lP3cFYjMngCaLGR/4YHM5Ytq1lDfdy/d31MLJ9nRND1836etapPGobteJK5Z
fRPqQFxdqScRI8CbTIBzS/G7FzoSQbAtB6kmq36dIa/0IJFYFekHhoaokrUOJPHK
m16uMFG/eGiYNZ/kY3seD9Cf4CZNdsAws09VVGTEXHhK0QAu+PwPXD+Z6rBu0AuS
vjq8QFmMTOyk2KTaJyUAKjoAC9LQgkuDoxQ0R7Mf+hENC/I0V46UUyRYseIiFesu
HBlxPzCW5MZDRncC6wICKTxxAl+hf5hqStWWZxb3VFX4ML0eKkT9Cf2XrxNdc5AT
1ZCZLdosbAwqvGm5AcjuQggKRAUSCCUS+cx6gLKOnlHBl1C7iOK2huSn3FlIXddn
aBP/YNDb7VfN+5uyAu9LGMk7TPW+ZqyvIhyEXEag9M7uFoOLnNZTI3i7u9fy3DDJ
clUsSu6uEHxh/+qMCMMuT0kYK4ZdodiRPY1S3jLXCrjbS3n0ZoVVP9kfx5Sl+F+X
Zr5bdP3yA2itrC0pz7bvJq0CsMZySYYoQShp+3fGKBrLV115tZU0sj5Iyl6uwSCx
ONN+WnigHBdTc+zrj0w+sWrEtJwaYemnJiiFBtoLL/UOsdhF2YZvyXflMnwbiPIl
tq2Tymz3td5Ht7RNfGv/g626M0B7F7Mf/g8GZlkPaorB/FtJJmmQt3bsXaln+tqv
b0uFSHIKnGgYfuHA3CfxFHC8uWOs1uGvy0iXIXmA6VAGtljsKpDkeaboCl4M+VTR
7LtYwDAp9rdl6Q/pj1IEjWSWsa4iE+QNdOsQ7mqdEQUmr6o1phHhpu47by7NPwkU
/aK0FrmtXONvCWT1yAFfgL+xkfusSWtQXNd5mIIEUu6vSUgrbZ6ao0TMBJoN9NTx
YQGgcClwkcOYzsj1bQoGjyObGDsl3G8HZe9zlwuFTsNIp9ny25JRsA+wKm7x3X7e
uT1j6OhoUjgyh4AZpVtvN0K6dqrxbGHkPpdJDm1gBIJeWbbtPTXR1T/fcTHcCtvR
jbTJO4JC+B/tWPj03/j4hFT2zqSESfO9z4+sOYcFKEUAd+3TZjfUFg4h9oUCfnOR
8fGGtrM8Y9YCnq22bUSNbmNDwhggkNBFrXrULugRzCAY81JJLWipCPWPRIA/6Ij4
KAx8nnH0FzebIkcc4BMFtYoyRGdhvS7YpSOZsDx9d7BYvfFwqKx2HBbtiqdDn9iF
GJS/uW4ZwXMbEXL3/a7z4cAoXMOh55Mm9I2Ml5UAZYNO02Y80NuRo+LQMKYIS0Xl
FhXROSJMNkc5ELVxz6J516qBsIJiLQMSrLhNXQlznpSucPBuJ5l17coTNpupwoug
7bFYBuJVqfYtJ2WZe95B/AnkD7nC/K6BsZtd4IAziuBEX3zrKaH1pgm16YudlOa0
uvpT90NRffh8Bmms4pnWJg1dylKhw1IJ+UvbyvBWi2FDfWHOKYY1/iqec9kpFQQO
8tmsfCfDOWyxxmmaKKveJwQT8ypOJUyc/iqxTen99LkiStngM32crGaDFXtlgG7i
2M+RjKw471Fs2U9ahQPeZW/4bEJb7cfVYG+uYaBXXg4BdviFhAwUoTl4HKPPjLNo
wLCa00kxydKOHSQy/gwV8KXvI6PWboC91BjJfbpYzKVTp8Ewq6mQQBzCDdz/e7tU
3WISyYezdFz+pitRP65gHyozNfVn46awUb6RBLJA/lEoClRrmjYeeZb9Gk7lZJgx
zhOHev3IDKisNFftSx3k4M8wdTq2QMq6OiAJ6YLFGddxlji2+7knX1+mvn1qbRgH
2rSoXWUZqJeuSbgEh1UHmCNUiUxq9nf1E4S7V199/QGWSluzE6AM/T8xba25NhWT
ty8I7f4ICK2jh6r4F84SOxVSeQylfbD5JcenpLpzN00b773a6T8/+ogwtCG3QN/0
t/wbQ4E1L65vRsc0LCGSPeInKiaYdmif5tuIVlXbXIM2TaTcIZu1vwYu2hUL8yQI
jv8Y2gHKr3QMQ8y+TyxtoskMYb850Tnl7+C3nZGWvh9bMhhtxMW33cmiagW05Olc
uPBGVxmEd758wke2PF8jhHxUeMQDdTaY5d9QpqKhE1dSeLy0HK33XvVighlbv+l8
dh6T8xyoLZsLTXGZdUVTrFJqMbp19y9qjBx20c38r4EOjnbxNG9Wu+nr+L+yuk2K
23DLsKK5Vn75qrD5U0YQbWFaW8q5aXE1vE11coVL6GmdI7CjJIUV2T3hMnCukZLE
Z68lGN1wfNMz6Ru04bk63SiLMs1O+Kq7yaw/xDTIktgQQHgxHce/vI8DOBVByRZL
KVNqCKCNXxF0sQ3izxO2HcBU9qRCtAfNDUYEz6ZI7rwCbO2MqbWqKVPDCL8/z5Yd
JitVJgd2QS1uPTkYBvol3cgQ+w+iGQgPMUKHdJA3eI40cNmmjKiHRFbKCQPLQ2Vw
t9UbrJhHcuHlrgdYByIaDxGbwgOMHxK1M26atLhES54yf7C8vKm8z1rcU5ose5eD
RNr15GajXbngHeN0jZ5Zity9nibMNaA7wglMsHCabrhpBoKS0CIBD1NNklD7FQtu
C81kow0IwSqRIKVkdy2DGvoQHEaRewEudpvKhWwE1N+1Cca3FtLOSRRPQ9TYekwX
YmMFNqrlVt5fa5Lc4q+2UxFCifFWTp9hVOlS/9DWZLfQ6qbyzTrD/ATz3zta1YKO
zVPQLumK9xd8loil4TELA2h3eRI+pmTPiWK3fAkCHPNWCQa2iWbWRcxFkjPNNoJD
iR1ilE1l9NOjalwcEr9SWwvo5dUPf99G3GVnsFFoZ1uI78oJHhGjam+r4MBMmRy0
y3YSMGOnPFNKzHY2J/vAysi6kahRhQDsgZEBFULBhv3a60S74jAUpIVxQTbaPhwG
P/3NihMs6gGaZPZ2dDUCq9kXnra5RFjx9n98fJpRYgBPHKgGfsUd6a5uZ0YfRRXK
ximQ4qk+Y6Lv3H0u/C67+APynddSm/qVT1TzxZOo1xSvYQVjcU6iio+AxJPdhowc
ixnTCxSz0eDOY7of0YsY9q0ZhWR97fa47KcuNaFS1CnH7P37VtpUqSbeQg/qw15/
XbgYXqo2LyLrwGakwj25sA57cnD558Ar1ixkgZKTnBnn9tygW//lfqT+QyFBYHLC
k6qTcBzQZLCXppANeuceFhatKPEdSQP12ozjaZySmP2q2oF36Q/dtQvzaIR3dXYN
Tjjprj/UeL7A5KzDMixn0JyM4lsFTz4uNyD8njIOss5w23yrMA1hflhXoKUUaKkV
X+RUwZ16+6JLqrod3Q5Jv7VvFIPlQF6YfoiCPRLOu12WAf6WTQxr4fVW/9zeTMyr
0FsCZ4bDWsagpehz7+gQ9W9bdbCEzHbv9ELVe7RLFa0i5W16IyyWK0uDTL8vQfNB
sze3+z3FfcEPw/b1/iFrMdlYQ6Ao7rxNzZHo9Jvuc6gVaPse6wpL0KTHaQFiv+VH
j768Wp4jqXqbeJ6WP9WcweW42YkoXUP94OWVcK1JH1sWtAA0pyRmRiP2/5bvOe0Z
5z2KeYB+oFZ9DK4oI8Jfk/FSi1cFfRs9Rsp49yVuE0l1Wv3R1xBXEgLg8KCdPhIs
iHqmeNWKxO0Ivgb1eRZebuj7OwDch3ilBajOpfqPcPGhHiFFFBrXJAI/feINlrmq
YxHBhkvMa06XahzOLVHv0ZRmTGGlA9+bujsgygh0W9X/rgM43WC71Qvdk40Fklac
iEXv6NMKdeDJ2aHOWOnKG9bmoHQUZrppAInrrlIKI/BgW3Uawb+b300Kut4xk3pQ
DCu8QiqtKM9iAxFKRPHd8m0hbQ1vj0dsRbYMH/7XZhOrA93I6f6GZ2qAQObW0Akt
wW2Vv4+G3IjMFghqV4UyHP2m6cxP9pKcwPBNlQNzjMYF/qFL6gdWEKFG5qUa7sWm
RWy/y8IU+Y7Z7pKT6WwbmRvj05uxjosHC35xxvmncRwxnHGpLt0oKUQWKa/GKD1m
YJvfeS2NkUZDTigDjAeO+rupO7BITQ2CJcxSTt8nXpGmjL9V8wN1mkdFlcDyofiS
iEEEppg2ansVgCvV1mnneWysHy6tUKKq4aBoQDNwUC0XZ/s+PvLjSFzI33GgJoG8
EIHLLx286tFvZQovhaQg7eITMSxSviOa+zLCdCUgwacJaMyafnm2mGUFebysZt6U
aurwePqP2zpROB0JkbDAMsauY86WUkp7i9MLKM6SDX5GPP5gm10TGkbOwsQIvogL
TY0DGLtmXHLC5sqK3NQ7kjxVlLAm19GMFOuguY/rGBKHy0JsKnSfxWHcCXfto4C9
ScKkY7PjscCi/lbydb8QJHH2KMDMbwn+mNKX6VR4RelmpphWbMxOhvVts0zhOt9f
nf1T3PsIryaZiAdAXkFDiANAP6efatGYragvCpeGWG00g8UKEgAZgjRsNgy/giBV
r+sdUhdT9m3YsJ0yIRfwWL0F4i79dE9e2dUhauG1IC7TxztZ1Q8kC5jtHE2yjIc/
/DCNoWPLt6JQbELa2F76RheR86kBeRQ0sbGQrvA0W9s/DjTWpX3ixXvDttJnpRh0
0LySg1LJgwTXf4dIKxAeQpCqn+u/oL/1otqkYt3S3exqAcjDot/YBmRAiKDONzGD
TftPqqdOnP5dTxP1wOHw2z4DcDP5S97ITvdUnNdbJVIsEFCap/XRlG/XyLWsjizk
ORFwF7y/xXZ8mDskHYjvJ8WUmGvQWlShybFSg/raXeWZLc9HnwrHZZ5M3wRau+An
JgE6PmzTgoG6Y7H/IQ3FKHoDt4r9h1Q3v6+tP280ijAQonz7a8h4EYmHLHqL+8YF
uSZhLLkxAGBn/pDNgRWHHbjS8QxDYYzmxHJE9WyUWcfIN6kVWfg+mdxgM0IMdKRR
JuOk6klAoYV9ShoVCQQ5EnWkGzjbG9X7N49XFvKCcuxX4N7CkwLqg9ki5+O6bFOm
WhBI+5KT1OrWER+SMskurYCcgzhCClozPm/z84Fhy84om3pOvNqEgWcAVUJCyskg
GYs649sDaJDz2SCGJcA7CAbyeEwgW6Qq9baE/8BkTT+tUB24YRPKqZh6Vv0mVGgD
3cXIePiKa/eXj2QqNhhTh0BaXbGt6igD2ZyZ1aNwm03OHOBp9X4VYkY8hm/OEuL6
03sHW1TNgvRpwY4SWGzZvbwtM2kyjpXebHl+IRMMbBgwOx0fHlSI2E2qCsuV+23i
J2LtQEpXhPwkfvofX63ozwxqJGiAJooCNQCkfg7rvAFbelHaJuOqxpE23S5KLvm3
zMb0tGKPzGKCc4uk3GClVpShkSmkmXqlcdqNLg7iAcXhZXbwfOWn3GZn2GzAqdez
PaIgZKIBQcZmTxGcA2hDSj7icTmnb0JGm2X0sFhIDfT0nW9Ui9oW+P8b+X0xXvwu
CYCxfNSF2kNCNUmR+oSJ6qegaOohZiMbnvEHFkQL4WlivTlbpCsIg8v4GgvURIeq
RAprk9n6PTM4xTwZHBHeyhwH9ovJHSk+ZeOT1n1omqSGcLrFYb8kPUXxj6nENI2q
DnwOtqnA5gjvJzzzQwplGH2aRMdgJKpTmLu0xA7V+9u5yuh1IKV+pnrDuLtW+JE6
SrhFMOlPKtcAVfzWaJRpGZ6sjWSJSE/uJJZy5CtXdCRup5OAuQzI5c72YZeDEqJa
7HQ5FIBayHcRqPuBq2mv/lP8M1Vj+swAUIPKkckC7RiPG24WiN1+cIbHSwU5b+Fx
qb2e1xKb2jgW6J0HTm2TLayLlCZZzDIrozWaFCrJaYCULTglWm7sEc7w3dq4djmD
lNAbHqpJxL1s6qZV14MXU/QJeSIZjblEyut6iMPUqG9eUrb8atySSoGfgz9+RCUh
h4lp95Loy2oC1JgeALcC2r0NRBO4ZB4hIgoGcWqwfQzktRCc2qE6mILoRft7CNng
sn3x0aPjFulBkMyMWXMCIKcdDrZdptOlwCKodrCDWbEEFTL1KVds1R2PriMNYsnk
3QsP1kinRt9n/o9FzSPOtBKQrquAJtXXMQTIeFL6mwpn1ui0XJZLtCFGC5VFMKJl
wVUuHKmiuuT8fc3yqMNsK822a0maGL5hlQSD8oyMQFhP+13loilXrY3/eadQqIf9
tCH7cUAdW6KwgpPjXWJypnRpGCzWgM0yEErW45Hfae1vSqnfU1IZ5rLInLuUEnVf
GRjLWtgcw1DxZhRGT7GTOOt5a2R0ecqMdbHFjfiPfusVAsde1ldWvD43pFwZEdN9
VXXQSkmFk0naRKh19Sok3PLayhLJ78xtk/GSCvcJXyP0oqeMOWyr0XPravIjSzw+
q6fzgvffkpuUFfRCVXdp9/Hlo2hfunJYy13l6seT9FrxdYjoGmaVDDSiEJDWqEvj
uKvcEDZTU+rv3q9mSGmylo9pezjxgrJa4KVuUpYgS3FuwxTGKkXKHY9js2JUN7CC
969EdEeBnArZ/2TlGW5+kJGk6j5oSZMid7sm1SCPFi3wRaJ676sDudpfWBsEhJIX
/0vTqenE9dIaUKVB4NSYtx/idRhHcBVFIDxyet7xGNzRspTQ2eq/hkjE6KVidrGD
2zcwiA7MkB0P4WDL/yGcVFZzLcJoHZFlSBS6xzbcu+xBidjdXAhdbeMXPK5lXn4D
7EG3w/gQ94kHLvmfcNgmtEuQMtPnqNb8COHVwU4JT3cvW196P+TSz7i3xnQNMpWZ
nAH3qyx1KVfrZaxqojU+n20eo8BPzlbs2icyi2JNpkDW2nZ8QnvmFHWpMRFOI2vJ
+BI5XsizU8s49E5rOW0o8UahUlwrpx26sSQJYQI5CGeG7IddS04sJnWbmaVFfBSF
bp3TcrwdYfE3D9rBYzUGw37n0u6IHbStUc4vHq6naWnO+OU0hiLa2loPthw6t+2Q
UnKmt0JDJ59QUWl+mJs5eWrJCMP+Bv4xdIss2JbHyEe4abaTWrXM2bZqNaAx2XJo
5NDRGVab95RFI6Vhx3vhlH2M8LdqB+RHKebKBDPK89j0UwNf4ErygoDzZmay9q2B
Ai1gjEn7eFSpSw7pUwYmubyOLKrnnAn9dA4a2L4Dm1ElH44VcORmyrROW/CjkWGl
cRG6lo+4fCwHZgKMvg3Vvoo2qxUz8/71au6VNmfRHMY+gmPlan8lM2bNHw0dwW4v
4IzSgfR2b4LtzbJW0/w83Z9L30M5aWHyVQKAgQGF5Qn91cpNz/NivxxhPkVAr9d7
dv4XAp8zRQIYw42sbOhosvTEb6bpBoNGu/JWMgoiueI8Y44FSIyUZFutocVPQSJC
JBCf2XBLs6kX1zBbfoWDsJOvuvVKwuE++ZopRJTEBPzDdhCgSEhL+8vSWgdtGvbK
ojOVeHWsdGJj0lLGdjmPE7su0Fv/pxTUesFPPPyVQI+xDF3gV5AqPs3jv1K4RWxB
0GhvVec0aLHcoPCHj1n+E624QnxqWn0KPgsCy/vs/HD1fooKDrqcYuTaKDKyn0mv
LwJX7ZYuYOryvD9DpUP6R75YIlsNlag6cX4bTx/z2XCMAYxxmsyWBVANjnQZGbvR
ryKLny/w/Q/lmll479UqADIEFMEUEAUI8a4maLS17jXmu/ORazJ1eyMSk1A5W8ph
c7a1LByjnb9qO7E2KdjMBKh8GZyaV17UxnE1og1AOCbkgtjlG8ERey+RkDBg5CqX
CFOsvWeIiGMEPjAFQWBFEdln9nuDeGrDcr15tVD18gIaWXSdOyycWYaY7RyaDaWV
O6WMmkY4b2YyS7gkHkokZH8vXo2N8GHx7V/69cEoobr7jD5SojPVISho6SINOAzm
4jJQM6ObH5HxrVl5j8WxNjI2QDuXbINkpLMTNR3NsRAHOeIrXuXAlyXEYn3TgPy0
D/jKhcoQYLwW1vk72UTK8wJbsH6UtnrdvDVXtU9/f6jAik7mKgQCyYKTTAZtY3AZ
iM4uQFaBkJvMOQVmSDXWtesEWO/eLuZHTTTk1ynwxJGRe0bd3/FjK1M3LsR99oB0
3AFF3hex+i3rK4f138meE/x8cHjReBSdErTF0CsCJZO3r5Kng4DvY/0kQE7pbNg1
xCrs7DK3pPt3yvXX6idVlB05N4KvdLmfnmFf79qinm5UQ83qs08bizXyrYxQSNDU
2arJWN5kFHRYJRIdEmkr+Gf8pVH8NSkCLelW/sKvP863/rbPgVVImTql9kxQPF8D
yRg/ny8HFbO/fCYeNK2Zq87bHOs3d1LvdDXbK/9vzrFUeMpZSwfUr+TE3nThCCWT
2VZO7WkBRciBlw4F/RlnEdjre5iMt02611gCygoMm++3hQy3LTZKQ7DBt6PnkDbx
uWYSYk/8AL1QbRXA2xp5XM3bw51nB/2zPz+GCTro2+hHOqdeAva7b7VLt2kdc7ft
Uf9XQj3kb9JnGLG68Leey8+nnNzhP9ZR6OtmVpRUZnHpFgBs7j+Rnu32i64Qww6v
2n8HN3tiKTVDBCoL4wPrtX9K6kp7TBho/++NOalMEIYmN667+nTi09QJAILPtHP/
CdapvUPOcuYE9q1KO/b1viQxpFDFYZLZ9eipe5tCa4W2zKRV6qw3pA5CLejJAvKw
XCGZ4yObFv1nBsebaL4Z/6j/iHuRZ6e7mnX5C4MiG1yjAHaw5X+NoDhz6YeFkFKr
lBPMGcnFja8xIWFYyV+UoqfPzaJbITqg59ukJ/wnwW8fyvqSMnrktb+uJSD863bX
REHIWvzWpYNhkcqKwJpM5W8svxgNWeRc9/uG3GGv9S/dFjo7KITX7VGMczKkI1ws
CkHvbJFS4qrzsTBYkLa9rii/2xhU7GYfoWbYYg69wkJtInKv96RK6Z2l2NoAOHt2
NKOehvuLlHob8OOd0/w8GGwkXQvJHovusSLFEryZdCzyqm9nFk0mNsYEj+dSPg3t
d8mf/VN2d2B93goZ+quXIdFf3MdvmOOljReJofrvE5VWab+2k+I+Hg283uA5HQyx
vUWU5IOhvKxy3cG1q6f6FU5r4tLuPuBxo4HFt72UUlBsPX039pnYB7sSGe4TAAk4
1mPIF7FtiwMMhTMifc7Fp3YZs26B/2W5kCKobuA8P99ZASENNMZoNeu3wMtooFrB
eNasNlG1QD13YVTx+QOaEjHWqpjb2E3RHFsQu1UCxFzR9v6BjxXnhr2taKR8tArb
HxX47YHtfUC2iyQM591TEiRnnM0dfJcOwCdqcSNG14hzQFLxNvfmMx5CDgXst1NG
9SN3NXGNbWmXs89jSN20ngpJ8YtFomrKg+BkkSTFvR1i8E1v37uLK3dfz0OuGjkk
R2vVu/R15lDBds9JyN4iH/q76DmcUmvl7vCKg1z+ABc9eEyE255qpHGJNtV29ylR
tSLEfwI+hDEDz1IE7J2v0popH2JDIqeJqkT+GugymDrvoLz4VG6b8RKIpak0PoPE
5YmcUb0YMSGf2NOFlNjN+MqkRHTgwyHQ5x4SYrH9GGiVeuN1c0++GaP2bSo7NzHY
mBjHzkT6YeTpDMOGLhFCKINobPLxfrbcv6xm/F/kmEW1WAFmvRa+OV5csafGH6SI
ztIeXFK75HGKNbwTE22Kd4CBoby4o1SB3qZp2kDBrekx670LiBY3mxOJBBD8eitg
gU+gaKH7t908wZa8IkcECPtDhzx/CnDFzGzjUiJ0c7RX2Ob1fDIkbupWjFfUHXE5
haq63QftBAuof3P82KcaRTwX46CWtcvWk6CBuVgBHMLIVpBzGSLU7e+5sH3QrlI0
9769nJ/ZcXn6BGw65DmvoTC5wlrrI1SEqwqVUnJXzGGgdl1/oI/vLtzYpt0uCcQN
YK5Y/rmXepTWFVlgd1sx3PTkxq5a9OBLSn/Y4nDP88fukGyFm34ckZ5iursKFq7C
940mrZM0a4wtb05Lv+UeEV2aW1Ve4MyASVPJw8+yt0Z4zBZWGjlrbI8Mh+UP487r
xHXhityD+b5iKbZ2Z47mlWYR6Kaw6cA2CZwAhCVKWsg1K8rO83klotfngcT4oRiq
nx4rddkLcEVPFfyrfqxlqqYPn/IJX8YCFyxVxa3JFeynPx1pxY5zOCBnlelZxlqD
5pXg6MHUH2qaXcJ5dXSL1T+3BfTBzAJfY2NxPxyfxMWaHvGgql7fiNJLpJyAXHim
cZ+6rrkNbNe5Adc2RBup2uYKu4KwceYkxIBuwRaQgnCLCoV9PUX2lSuoLy+wjQ2G
sheGB90JQ9f1BFWY8XdjT9kWifP+82Cse0jj/6deU6ekv3vlrGv83Osv+751H7s0
H2gOUopH5GRKJDdznQr7LzLzLr4Bb100DoQIjwwuV1ZwSjNcYf6hyHVAumU9OScN
NNz6Z57M5TwZzdGjyXCqc5W0Mmn29QfkMzlLHnH7iXu6SxkrKg4u1U/grC+6ft+6
Wnn5ozvlvRG1Am7ZAnypHfk4NIJRFUOfhhrMnI1j0vPPvADFGK+1NLKtEiOeJLSr
JPEayQ7p0MOub0Kd6tMqRErZ4BgiO2Y8nHqVpDxLRxt69ygt2DAZlNJCatgx8aBW
mS8fW9A1S127ZCX1dB34wremQTs0q4tlsduIOdfdPAntySFnVkTJGs4v7/qLSwll
dVg7Qy/pbeR9bJt7IZ19aY25bVMcyCC0ghTk6OvAXHSDxBqKx0sQlzLw+thfisd7
b3lXohGptqJzdGBNw+AqE2TP1nbSPJCnuluyv320APBKoBx7KIYa0U1+L/79mTTC
4D440dhk9JKXkzT3Pn7l+UFJBNeS5mW4oxihIPWO6gNKVqfaF0eGtNSYSK44t225
ACHdtAw4V8Hn3wwcP10pcKSSa0RL6ff76Wi/GHIXZmgxx3bXXXkvD9Sn+C+ItQR/
ukDke+fxFhseLa515ojKLxGA3VdmWIM9HWS5ue+K+EPbAp0FuDFsTDZtm8KE4d/1
kvFT0RT58RYVR1PbA7NYBQrPCMpTfjBcbJ7q3ztXtvo34QoEpXknNCF5a4yeB46k
4FaEEtmAAo9De2mT+7llcydB5Pw7AmWtC8ww60mWJAIKL9/3kA7Qyh04BTis2ALV
quNBGQ4+eYeXcKiTei2hPWLhGP8kb+ta7j0wQK/Pus042+5HW6lst6leXRCrvs0e
CJ7vhA90ue4oZmk6kHlYNslB5e/61D1EUnyMMQGix1YurFR6iUMkdLQtJqsNozre
XXC7DNmfHfQNofw0cNvAVRMdaXy3NyfvLQe7isHVH3SLEywk7ZRxYvGOIoWhqU9S
D2ByixMsljJMSmC14gUclwbjJ/4xFnrwtzDlst1xZUtwWz/lIio6PBgs6AtEIcit
bWnzqcyhdX68An2NX/E7/mLbaPBGCKKuEUT5LZsCKX+duAknE0OpJpa4X7rK4XI9
8k/dzRmyCEO3/qPglUB8eMCi7ekfKMbuSWaUTNITTisFmX02jcWxbJFxnxS4oY4l
h2pn0DXK5c9lFE/tJ7QCRVYSPw+HkwhNgZ7GW0xNVuNQdRTE5KKWAVMC38eXoNwh
QvGnaH0vn3Gk9QhVBmhXwHRjn/YPMZ/c6VJV4gRbm4k83QkuB/5f1FQVo1DgKPqT
iQ/BBdJhF9k/9x8Wwp9EjhkhOqhyGkYpSR1DsQCOksqUosMjUe0C9mfeRB/Mn7y0
F+ajW4rC+qIjOBqEWKoN+AC/Dkw9GJyeaYZgv0sM5P6G9R1LgZJ5YT3wqq6NxKwv
mOwDTgeyL/EDrfaw0Q+kajmJZlg9CRVJz1TkanHvT9iwma/YdgeIAX8BJiL2t2/0
cQfDeLZu2CJhzG05hf+fd+nkl7dDMbmlJpVStuLt/5+uFgpUywjGoB4+BfDLgiRk
nHefwgsuDGiZjwVfrTbrn9ZzZwZkRaUgdzJT8N49PM7R0Uvp9rjgIUmQ7zn1akC3
igPLNAn+cmCPJjswJKP9pWajKn1mOxoP27IiELKwLgZCocmYgAAGs9NFshj0BkXD
3NSqgJryWO8P/GJBR+Jv8UAnX4F5yrdpLibS3K5jGD64YK4UiEc6RAmI6sKe7ieI
XEbJaDIKkzPTM81Ayu3UQ6EKA1YEyjT+eTHM7tEFVh1D0k45eIJnKsC4Krmhk7V2
P4/iwwI7diA1t/TawjkzLUXM+2DKFih4gtYSrptGApzW1nyjy88OLY4/jmwcYo7t
qCuCEUnsgewAAxGIbYMUMO0ZxptzLrH9NCy9rwG5G5K726ZJQhcNlUVnS/+hi7nC
Pr2z1V+YDSGu7dNEkhEivppMG24vKgdlx93EvJO8SUmUisEQAlDRUJe7FvYUmDLS
8SwnmejUg6pLnabubVW3lXZb91gzq5kYcbOI4QUolEzE8dbmlTdBBf+l9iIn+72M
IRcQ/VVEE9Dd5DA/6O+9QX1m8ZtD7yfb9aE4pis/ficygjO7nxZfgtpe3x9bmKoW
W72PP6Yx7rJL0EyHbAbORw0cJMX/zDtAITRmF2qh3rvVIIamLKSxnxDCvnQ3B1Vz
sIsvLCKGvkBVMfWdFLa8X4zwUTZAOkH3FcsxAn+GsfdmiXFZWmb4//cP/HmlGhUB
LtZREQcaSAjKCzmeePa6Wpyn5FAbGXr2KwimqTfT6WNiaTEFkM12cfm9b/OfAeb8
9VnuHJoSIUDxhKwMzUtFD/XEVpU2ItmYaDhbLa5mqYwxJSE+y2GOcycfIkD1Rrfb
IOwaNB1NPdgjzFmTrWn3HSGQ0C60ai2Inv5KKm+TiHbUj4e+lJ2MqoQlWKSYIets
SS8ZZP3tayV0UFXCee0GdZ7R0D3OhdmcFiY9/qfcagiW0VrrzHe1jH9Oqu//Q5fL
UV6wWGdtPgu7nZBgEUUS+V2a+VmYPpp2khH1XjhsEy7GG9uafITwCZK8jLuAB3/T
SXYhPnCGYuAiTVNg5VVdU8d2nheMvPMleOSDOJO+Vrtgsu2G9QZTwVqeNQLwqXg2
iuWmXfPt8oWOdXwHjDqsF/8W/BVmSSp7Zwy18y7w38isoA4ZZEu+/zXWFl8Aw0al
4sXAvGe7fvIZrwG8WWFjVOikyKS3k/SRyspuzVDXcv35tMEWF8qbS/eniVQW9MsM
zMbf3E8epqXGydBLlloaXs/btiVb8vlzh0oCoF7US3xx5e3rRt8dA1a5trCnj3oI
AS+G9VkpEs0dF0lv6RrcHlytH7/7krrkTsnRzrBqyGl0Nz/7l+/qOwJIay69N/Qs
7MqGH2DNkBaV7LZN3haYTONY8X/w3gShVl9n3v68L72OSlkQsQqBswqcoWkyt7+1
N7RQ2dkfFbuDJT2RpcQsSQSd/Omp6q6diJYW3onHtf1JfCAQBPWHbjucY63RRxCl
a7V9Q+u9CqP+IeC6QxqUudVsne57V1yUcXyrINl3CPCrtGBtRpJ7lxiwH3jft7ev
6/9W5WO8BEM6kyQpMC0FbEPCpk3wF4R4CGyiGZ1w9Ws58vreXyqfFKyoaxQyMPXT
JNn5wp9/O+qGIZqsVDQcLYdEyohM5H/oavXKfx73Q1Vts/Q9zbnJbCDaxySQApzy
yES/PHID8QWXoWrD/B2wM9duoiaARTPT6MSa/wYuIcgda86eb2mpmlbfA4Tw4Fvs
avNrIQhdi5lHOzn9kyge/O3oiqBXxgAyGjFpdTtpV7nLbJnQvuscOVtcHOcPd2jr
QBswfXkwbStvNo7cDK6cANDj9qvYmxCO4dDssVez1TzGlH90QdfZsWXWjspZwavn
1g+nevLyAm3M4L0Vpmr1M07NLiQKE1SBUeyHG0U2RwjjVg6+j8E6LNxB2R4sx+W/
GIxFTU9xyndzxw3ajYeKWwPcy7C2vxIAIBAwUNSU4DhfkdnzPhVRt5PA1LhqNtkV
pfR95EEaSiG+WhVSmKRsEWvGQUlvls3ZMTUGebW4wDiAYPxEeZF0hQ8eUtv6/2GK
tS5QEqcYPMH8QmG2jjuXQJXaqbDjSwc+fkY58vMwlW1ov6pFS7oDz5yKIz6GFg6M
pKJukI0a8FQtngrKHN8N081I5PbgmRBjrtPfNoXwML7dS0zlCyHSB42OeZ8VKUOw
PWi5kDjQMVk2nhEBNs62pJnBa0/sdYYacvwqXTiHkxaDa1xdE8GnW+tGoYf+uXdU
AX8GuS2m+reJ+6di9wdTvO9/+x8nUAD2YJ30+G5ZtQWKuonPrKkKKjjAXpsuZnPi
pN4YTj64+Ir7DbI59KhViiEEGWNj0aH2lPAmMh9YUQ73Ok50fofSUTNTnxxtZwsF
30UIYru0lx1z0Gagk9gqrgPOxA/vaSv+BbqmRMy2lz/4jwvaTZFlBcOJM6XvKE9u
ZVsKDXOWRNxtY5N9NzMjCOZmJZ/40ttmE8pODn4zstGR8163uM4iF0Q8mi6B4Glk
3FpLvf57+IDQ5zlFqiBUm6EQLXfuLdFzVLKbSekm7xNcEXj+/W0LMLV3So8mCrDU
lXmM09XHSFbBi+OBnzxoe2gLYNPdhLhDNESNYcyw+mFRCJs8TSNI3J+ItGVLWlgh
MkyjMhrw2M2uJw8vSFRv4Bk5XfuRky3hh05PM02jwwRkOlh8pvl+ToBcbK19ztfn
DLGs1nwnt8kXq4ctfHPXS7mpa39bOy4KzskfFmXt9WmFjE92UHN3eJREw92UkM17
DbsZwoauU11VMr8yFD/TyIVZmZhqHnysJxdJagtlUe9jg+VafPixeLpHuOcbNAn1
uOvoW8ixTTFsm7AMWVkFS1n6Hjlj4wpT9Oj1bMTK+7xdgGz0YL3WIn0AXOZwxe21
vXPfGpyNczl8G9MxkQYpzqZHbvugAsJ+I6yOh4Mxuj40lV38dTUrXjGK6iDDBqkO
jWvnrKzvmv0LSNEeh9UgPQ9z1YzgT85YOUY59m6cPyf8ENKFxrmEcmiumInYHZvr
4F8sUEo5S/Tw0VqRTtfXZ2S/EOPc+9vz6QHRiCwhbdVaDPmk4v5e8V1Uk6Ropm6r
ay0fwoeWDNk/LaLzo4vwIJfjgCR9fqcCz9xtnGwmlejSOPFaDJehhMbkK3B1G321
puKaJd2xU3N3Z/HnMfvZdYOPhoJfURADcjO0aQGZEoVmEW6TlyUueQQRpkUy+VA7
qSRf8g7i/CIE7D0bOPU9Fyy4eSH8JL1diSE0mYhO/4E17Nc00Xx+AjWTIPa8lMWS
Go4NzVm+RNyxvIL0dVWLU/lNcO6Bk/Pke233pgBQKw/d1S6BV1PAJNnnVFvkkfcE
+mKAauAbgL/ARyo1NG6fDGmvpQaoLqa+ZXXsSBNz7+LON3nOkAW9dgWtms7VCjUA
tIwi/8hu5q0lobLKNT1hFGQ7wFwt952LdEAtuJ/wip7fH+Iv/p/v9/O6vxRfkQr9
sIYRkiUwDfVFeZUPgTNsqH87bmyIjSXInQlSrxYhSRgpCy5nOEylHdJjhimh94Fc
qHtlq2o/0yE8mMw/tjpi3k3kwlCfuicldOwu5J1kbkpE9KVjdmuhtu0qTDj32b6F
zmaCj486if7NRpjRL2jDSW859cjo18kpIhApKzBlIw999RRilMCn7pDXPfkq0k0X
K91ObtVE9bOX3WAVsPIlhlE86ufM2QaCikNmZse0hRLgl8uvThDQv+xP0hehECsf
IRnEqD7Ab2SR7/p8sq/n+hbqL0S+mJjWJLCMx1CBoHcYbMgV/1pAs9fn7m75tmNc
kPHXzLID2eDqGkE1gNlkmXdTxTpEp7Cfq1imlGl7/FZRMmdhAqT4I+czRQJ6+1sc
doJ4DPHFVHQbq9OCpp4KWphvCf4+G1tzQp0Ism5awBD/bvuikFsR/+DYk2NjObJQ
VQVrV0rf8GRfJrvEmmNvXg/6ld4xftZmLDO8Sjzh4VQeAvZGehnkCwH9jJ6MSGq0
faGyM6OCu45GihZCflOfVNv7JrNMeUWRRxy/wgsH9g3hf2KICWNEe9aVEWt71cPa
3LPJk/3zuGF24GnmxDBZpqKDHbfoA4W8PFxZ6eLIS+988bwawuq09EA1Rl+JLJU2
bCnfb00gRVH4TZia42Qw9TfzZfq3aP3az9ZD1Zq88jtzw5AhyWgDNGMGEn4drnob
QICNkTN26uqR5cpMJm2d05AYodSxMoYeQbV50iuxzHRED3TIms6mBV7C0xXNSUvq
dOS4kKsergGVedjwEa+Oyfbl2fBBkS+HJ6SOTh07jD57YoVa3GD/npZkxwD1J6kp
xBU6tLPzxLSOpGxIiqMLLXv9+nYFaneXRuhRdi7N9jZ1JsSviYz7y/wUa0N+r642
4KjgZs0kduy2ZJWSGwytF+zC4hCQ4n184CffrEJuk7t8fT60JSg1FpiMl7KN6Ril
FXTqGCqxECOg9xPAxy6XDlsib9f9u1t0BeFlX6TrW4CxoWtq29CWyKYDRzvkC5zn
6LRdS+dY2fohSVNkWaErNDQcySlEtiZ2rNqegGaGgq6Qg24YMfN84jgpJAy9SfEP
W3kflW5DOSXWqbuRJaHfAUwBOqZp3jPH8cd1KNJrcZXhGF8XRLOzL2OjM09W5ZFI
mpSAO+xlCQISJCkPkF2938mQoNxlYPLm5WzrCUPpA1VnpJlb4rpwuNp/4eU9qYMI
GixVg5U2PX3mtYxalYR2Bv9vlRmEAUlxXsNiD5oMcTm98lYJ2Yzy7/M1Wr0qNrwe
lmMaNfjt5xxl2bxlGQ+820cq+OOyWgi80G+rarlk+YbNckvUuzY956zdXNS6trY+
0JIbs5xqWwoElBI1KN7BTwx9A0yTldeSVWN0rpjqBXvgjLe/PzOp9DKOSNXZ/Zzy
AjsodHTJlpAd7IgtVvtUO/7JzLkW6RbxtwufHGwhgXmKjcqVLmJqTfmVV5RO7LJI
GaPMByP3GgbItko8TNxiAjzRvXDR/N+Y/Ro9p5IEDGhj4T1TTIaYXmtkqKbq2qMe
YtFG5Om9OqewG+o6/D3EL5On+rNFUVdmU7W23PbFSLpYdnkR16QiUiFkZyXAplbc
7ggvKWLPIZ+bdVwCiNiqd4wwrHzLl5X6+sRnyFQ3vZ4REmY6cgg7HgHgDW8rSAac
Uy4RNJxRi3nitDOETsKgKZFH+fjsUXu9iY3lFaUAXhA0OU1N32TziW4j9+MJf8Aj
FdoWAELSlry/sUXjhDfhdlBU2n8kBemnygml6+56fYkV5OGPyK1Dr/IWJtWB2JVH
Zx7+DH7/ulwO7nehMqk6ZCXLuQNN4DZKEHDensrms9R0VqRBE0W+WuccjNVaAbfI
dj30ULPV88ShdoK6+s2vvLKL/PLVDvMBmEwseoE2hTFyn1NgUyGA9L6JRtBUf8ky
88DxPiPinW0Um88t6QgEjRipQP4MHmN+pT48IrOEQcdFxEWrXF2mKzVOgMEGKSPM
qHqljDEV+8dbJnoN/Mysb45v0YoSBOYytnPF+uVacEH1wL4/fqoNGOCnl2U66LH8
2oIa8ixlhWAV2BpdNlZCCeg9DVLU21A7pu4M4DQAsI03TLWeVrzNGbhd2pTEiS8L
wqXhRZhsC3hOGPOy9DYtbGcnPlRoSSjh2qjJNc0DLVBD/YH/IdxOJv26YkgJqFO1
bPl8VhQR2ew1xquowAFedNhR0PaSPFq05o1SbXtt1LHla/NnoVK9trSIPAxkJJea
BdKvWnDJiaZCvFw/Jok3wjM8ELmlaa5xbp2Hhi1QSLs+JmI3u3T6zTtiJg2ApXGu
rM6+0H6CGn1f9Fg7/6z68ma+emWqPIITqvNg8IjeAHaNpNWmZ5y6Ndtv1a6aQYBS
rkMVNAsKRYG7CCCDckAT0LjItzDdxvwl99o6Sy3aLdlQpv1Xdl5ehaU3Dner+QyM
I6BaDqFE0LJwnAGXbnm2K3vfe1fmODt0Me949HYkf9IrfF8k5lM543rkt0U2pEOR
r5QjCBWrkhP2ug2vikH1cAfm2ziwiDUwEg1j5QpD6p5WmaPPhzxPXIOGlqIAd6lT
i8Q+viTDiDLeH602jT0NBB6AUIzeiaJjoIpXWttB5uQ291C6hrE3aS8PPGHyqrTH
XGTsaUncLsQ4X49gwRfj+ocRGdGY9pEX2Aio54nRiUPQ13UMBpowa61e4+vD/Vbl
5wp/NPpEZj96iKYCFRJ2UQ2YOcQU56CfXVTQyUT5fZE5lI5HPP6Ma8GrKvCCrRwO
O3vY4wHd5l+Ews9I+PExIfxYRsHBtRTNofwFPOw0LoLwXePFeJzB6bORqPORGWuI
q+64MPVV3Eu5wKHqw4qedBqU3CQjyGBQ8TD4b7HXxy58+qfYsS1COgD9n3AeBFp2
VYOSMv37Oxg5c+Ykjm0ammPacLfuzrTjjdmNuUaZuSslBSNZXMHx+L+S7/HqzP+s
akxolGp8KT8HFQT7dEcoCPyrgUhouxQdgP3wTGTazKUe/FtDAYNLh76re7xSXwBP
oV92NbyiGRwZ1pBv+slWjRuszaHCJGH8exSDjTZ9Dv3WSHV10/caBzfWGO5Hwduh
yydtEd0m9ks17k9LFIr3aYLzuIqA6WaNBuxVB2a0z9hdMrmkmISa1TknOfqIoOqB
3vGlWtqn4f/0nnRVUXdCmFveeupJ9TdrZV70aAd1FWPUx6wrci4nQhqq1ok8zlaC
7AaDfkRsM3U51jMLKvGrnJTqQ64x7XusJEG/R6KSH8Vum+Cbk7JVayEjBdLqo/OE
V0nKgOylFesQNpU4NzW/TCHycjqD4XaKVaSmQP6vGgWQW9ZqrU6Q3yIIWZTLyM5V
FHNI1NPUaV4i+8w+SO3y/zLW/lVUXsLM58ZtqHUMy/7DZQi/KBiLWaGHjyzJ96qb
BO+JixFUtdoAgMamquDUVK7sMJmsdEVPM3fzep4LvTXpv2JjynUjzT8jJqUjZDJ3
GRZYVAdFJDHBzmXkWTUlBMhBpEueTp2lxDlH/en8+tBSIwWpeYQqeeF47m/IG+kP
keSPGnRHi5QAq7sNfaY3j71txHtq/5IkGZXN2E1c+zsxeXtZitlziKim8Vz1HeZG
d7vvTqu3yLLaWlhlz0CidndniJRQOeMDmp8jz1xSEFBdL6MgItda1o0V8maHIxoQ
u996Cs9IZuCgizdCmbI4PD3Eyh6yMxEVaxa83PGmpseIEIyMmrUrX9JGaV4Kpm7N
+z0026pgpn6fZwCZNWFug2+wNWKsdcaJVjS5jD5JSQZPDTBzXcODIX3BzSROXg1N
63vOxBbNGlbm3m3st4pS8MkZv27CTMrHg8dKYG8Dt4zMlJ5Oxl9qbDfwHNVzYoTF
X1kYeLodQhVfVJ2tHuqbJxQk1l5gzVMExpb6CsJV7/yEJ4tfNhGTe/isiiWtDPCH
xHNnTkHvnuCDxpoS7YVIAku4XVx7WH28AAXMDjdIKRAcRtgtMJFUz7+6Krc9KkmA
Ydz22Iov6XjTFWfrhJtFrGRvbslC1h7fcDVCnCb/DDOXsH4SIkqDDex8GbBEKU10
bGli4EIRGzqzPiXe/i7nC0wI9dTwu+lwwI7/XbcLjwOe3C62W47FFr7cOPIFPP88
d97hsV291TCRQ9mpvLPVrJANQ3ISxNt+00F3U6nCijZf5NJpJGEbhnBzNfYo8Sua
ntAupI4hMrP9IoInfXR+5qmjO2o4aQEKEviFs/ZN+8z09zbCDZF3qepUGIXX/x47
oAsL5VDOIqfXjvZVP1lP4o1tR2zZRdgb3HWXduJS4KWdgGhdCDlqWTUvCduVgemc
vU5bKwACgmERGp3JHNV/Qprh1+msIZjZi20nEfjqjWG9gv/Q0k6bYkBeljPqO449
YiGMcLtEVCDaNpHi5mevTJxwxKa/3+cqC2rImrIbWipQZbglb0SKKhq0GNlHNwaj
FTpeFPp+cD/px0b3efXkC7i/WQDlFKEa/Bw9v9G136dmRaMeUz+ReF46o5x/mfOq
7w/gEMkh37s25Q6x5U0PWGFJ8RqcStMeASuEOo/PTVycZzABFgndlJstx4t5dYBP
8kMMmeYC2m6OkRB7ftNAfRM2/WJDO2EojLTwRrifgkFcyc+bkoh4blYR+XKuuLCU
2OjhzEELMh3jXrAMmRzG5nD2LnrLAgKmHo9HYWdYgjPEFhRt8xstyykih/t9oMsr
Cb4KltGBSP1afCcV8MeqlMe6tuak9p/JyMaKJ6Ki3AjTSzJuaoz+WPbYjvzEIrYq
/88fQx11SpbLGbeI+o8ZP2ZslIKB0xm0h2rwy1uukos9y3HG0Pg/OB5nPbXbbQm1
g3O44xSnfVOGyvF+RK/X1jfAimeHQYyh9A0deoeZhBYmsRBHY8P5FG9fe0OUWvA5
F24CIgMSplre+04MLDVVJrNJc2/3xasV6Xsv7RFjZ7LaAirBaIhHUgNY4ez7d+ha
15RkKfmPVX22Tn36yB5dmfe1iJNgED7r83g4bdsLPI8pp1SFNAwZ+MPDs9d4t51K
NLFfQzPC/aVhMyM+vCzpqiJfkoVXaQsA1MIdWa8n1DzyER3zZw7dEKR9ajbPm30/
OiT5LsVFqUl8y1iHT/ImYEkqVtulcyTs0pNlJDDPExt7j0YhQJviWOm/p3Fx5bko
610vOgI4AMIX6eHfztLyVs479hepia4CKZYMf6HZwKwu6Hf6jygLSWmTeI8jovgU
d1Go5Rytv7i9s47Hq+Q6Rn012b+wscXjlWLLmgoyk3DlUUxwYKc66taOqrICddvT
+oU8c2SQVMJVzH04NX+IsX05x5DRlpbrF7ZkgBkQpR/8efnohYnEdCbmUqGDcEAk
Y6VuG+oNiydF3IP8sA+IYveg/7xf5bthKSalOpFqvLKI+lSvTs14nbJg/hbZRKo8
VFVJnXeAVzyK2zPQzYaqvBKY7AaEYsOW697e3CQx18u6HiXPalKwoAbFJI8CvpJW
9lw2FpdeEmxApnwF0e4l6BcmOfAsNOwUz5f6jpBpWpjtNG8zhrnIUbsbRkXwH4c0
Y0EjOZofGESkNp0lb+Z6LA3KWPbrAxbOqjjsxe31ot+YfCwyBIqzu/kR/ZCWAMyJ
42c6bkGlfWLNUZA8b0T1Z4JksXj+SvbYTo4wFajy5wViLHAwVjF+sHKFEdhLpl3m
0JkHGIIwZd6DAwXKp61Vx1zSFLW7Xbkw5YngytpTa0bjUp8ei65/hWF/S5Ar1JO+
/4wxCdQA/sqoHOFNGESscypHNRf/VQdcywl1sF8sdjfjrVjszxY8rAO0vHN3+Dke
fTOSpc/kR7613fEJNy4ix9WdhX1HNDOSBQjM0mVT6pRQuCbDjVy6SkPl+pJ9putP
wNHl5H2jGb8m+og3cXEXewiCrDBCwFeO82cxGIzfKApq7AxRYjtzumV4qDEL+HdD
rdPnSmVOZ0oJiAH2bEkldQJtSntVcFAdRqct801lnkHZAPbC+UdKVQN0DoLXWXT4
+o9kWV8X8UIvs7VzJxrrhDaBhOY1xH1sOCosafh9ptgupt4+89yK3rRXS/kosv7T
0LXUB0d40dO5PBoMRafjFcQg5VHLvAjlY3Pi+9VvgVss0VxY7xlGm7tNTekyAIET
MrSf3kGhCxheIVbxtTA3l0/X6BAa228dVMr0OCz2w5+zvxoh5yyYd837dtDBiTPh
1ldtP54TPL1vDzvosre2YELDCELAaNk2eT015o7jAEq3ZuClwZkZ/2busRZtT/rE
UCEY4qZb4rQsCPIkVMoLKQqRjmpicrE1pxpHgRWbVFD3z9uHnwx68pMd7sVhDhxU
oHAjoAh2Pzb7AOrVNUCjUdbO0JBsQpvwoOvBe+cZNvm3CzicUeNjYZ8gxbHZ0LLC
E+i55i9X2GvOIWhc8GvD21BxbDKyJTYQC2pr6iGsy1Ir0pWmn/XuZ4ypqDIhnvPm
KNCA3C9S6EPsxemWhur51QUr7k4nhBnTQKIPaHu3AMhoW+bPJi07UTzUJM4aR/qI
GHHx5iAjPsMZDSTWpPHbIA3/ipIhYvPtgRI6AL2YO2/yptvA6aA9itTjaqIHGO0k
TZ1czmNUzzQQh7O5hGRqAvQaJvbNcSacbGi/DrcW1Bfd2OBBxeAS9mA4HbJfcObA
Vuzpi6zcC5jZ4IKgGjsM32270joCq+GAJ7bu4wWii/ylI7j/V9gNfd49yOGZ6bTc
AcOEbObgy/abx56ES5A9ODWbzCkIYBKLhPEvnctDjCEUUtcwCTc+JoH5kJ5r0AMI
usnlqX+8pln41x+v0Ip69IwKHW2dIGPje4ft+gAoyQmHy7A/Mjx+niyr+NOR784t
Z+c2mWCGRoUqkxPQNuQ6PHKuaj+2aebZuodv7N5yK+GhM67KfllIxNipFXd6iSrS
r7XHQqhts6w9mclpG7qb1/kWGvQHW3RtT5XzRkuKebDoiy5HepFI1+KTz6gRRgRk
M2j4FOiqt/s3DpNSdyKsULeurgvUHjfbyzdWmAFOrHHP/7mvbvzL2Vt8Y6NPdQ2Q
qlF564lFRUrvh0mYyDDpDsoWkcDbPqGklTa5xoHhTiwbqcjgRKyLccw14XztHaBw
4wZQOJrs37yiCkjt9FEPkamyxjMH4qDwOaEfAif3LY0UltGuyJ8ufaQLL4i6P1eH
dt5Fmr5y5PDb6tEh+Nr6U4o5rwLy/UR8ObW3aZwh/GaCVXXFC0mVzRnR+R/9URmY
AtNtH9hDhzlopV+l03oy7GDxiDNibdQR6S509JrZEE6q+wrHMNs6ZjykCLK3vRQa
5Cfhe+4Jg3wifTWBm3omWyp/QTNuaYP4O0l8dSp0m2u2n9TTmLt5GbAPcYd9wUu5
vMuwj7PLluwlM5hfW59+oTSOWsLdUljfqNkK4cIzjEGCXgQAban629ieJRbZIPbc
M26eIVYGusfzfVcdtQYklVKsBWHlDPYqVm6J/cD/Pf5KYPHR8V1dOeYEBStZbdMK
mFkj8D3sk2HXC5PHXSiT8OX4zApBA4sfrGcqNIP302g9lX/fhkbkCpoj/7jlGN38
EBBjzg0lO2OuYtU1yG9vAaojtqbloiH4SUheKEWyiKb3AU8yBar11tZU93tcKhYW
dKorkrvFOgaqHmRiPIFRbfNcLE0IXtWzkRFHK13T96/NLdwUIJHlt1s3FCz+GWwg
4cNDhYwCCzAe/Q1N30mkw39eNGPLKcRbmqmIZKHqPQ17lvf2b8TZ6qdKW77k+R23
BA4smlIXAi1Ob200is4//9HZrOAj2FNa5NKo5mTTWSC1ODCpPuIr1Wunas2JPUTJ
aX2vj9gmPr5OC/W/14ZM0WOqyDJalM3ldq7pgJVbSfiq6HOlh4wK36KUSA6tSdVM
PRI9w4HEmC2aKptNqPtdjMBoB+tVR3k+C9iIRWOgKtCVSxuj48azrky9OTxylNd4
jG+Jx71Hh3lRk4iPyCYFXxvV7KbAXCsNRAsJ9Pwuls1Pu4U2ba/8/AJHdom29hon
FUM+EPCNsa4yHD7HaxLKmFWgbMa2pDKmbUz9sqqCrMBR3A6mJ86UoeN8Z2upbpKD
QZclTl5aFBwiRHd2y6f8I5FyChzSYAEItpr74SIgwsLM6LBDOa/veALT0cuwlFij
Ea7JpI4C6dLihUNnRsedM1rPHQAQoYakY67W3Iw0knVlQBKObQ5I6zjvOfvOBTsc
Y2ZFv/55D4NgOBNJSgWxyZqJPzXwnBVBPzqvXG63Vax6zvMefWNV6G4FS9Ngp1p9
9Zcz4Np+rkstS3Xq0g9Y1q63STHEPIKKkh7isPeEC8O3Yscg4swxy7yYS/IOzBfu
YdMlyCMM6rnb4R8jjIC0q6IaQMSLbUsyFfy2zYi5w2URHf/zZrmLIjdNwkl45q7g
xWpCMqPTitYg37ukfkyIEUGQrrrVqo+j2uabBNsdvvSdjFMn69m1nyWQdhFgJyYL
7yz/rPSjb/wlsYgjNQ9etRSZCZJ2ZVWl9eLV9dBnhshIKJ1XPqx0i7PMpgmnlDp/
8kL6J8G9MRfKZ8EphEIgpG3EHKkNgmM48DFa9EtYey6wgOSAnH+yFgpZB+U0t6+p
wAj4yO8L2jNkjxSTJlGDoY6GETnaEXv3oB2UpJeNX0+HokiMaj6N8saHlICsKkyH
DpDiS2715Rd/Gqqx/qKiw0UkBiCC6EtrGGOtObxKmLOqn5cm9NXjKEmUqT79Na6r
VEr3PHUxu9ZyRsXUa0SESg2HRirYn2QAzZNHysPYqCrIXKM8kZfM1LfvcAKjN0C3
guFDm0Y0ShL4o5HjFfkU+OQFN243eTsZWxVx7oUxRJb58QzSWcUZESYJdRBTBvzo
n1d0Hdbqa32cmT9LL7Bbgdc9P/g010otYUNSfdovaTDI08nRoOeGLofFY+7SeGpG
qWiea2/XysiZghzmTZlvQ8rsqypwoPrH6lo696lDYLZJyF8XBPbxGgXhG5rx2xXS
3Kp7r4eHv6OBiXsOgcQSAEceZRH5fLZALdMhzPvCxeA65Srg+w0LdownjRZ8qbz8
hHIKhnGhB7kLn6GMzo65k7Co00YdnoWR7HvsQ2qIhB/VEBN5/495LlUE++mxZ3nr
LHn8q4Cm2uQ0WpI4VPYfAxYVEaVEpzTIjJ2o3qnecnSWAHamyA+uIqj5D6gv4MzG
8T3k+WHWcEwIeFhfNeznZIY11GQmxslbZgMF/kVpcF6XgkyShCzAET4obQVE1FNd
aQgd1UxZW7C8nGf4XOra1ydhiNm5zl1vrrSgmS3qc5ZKAkXIC9YrsBWOlU8mWmJf
83y7is9+LZqGtCy1ql6KBi1wG5VEALT6bWkF0b44Gf/2Ib7RAomIDWxFvirgQpK3
9RjQPcZNLYXu5MUVsCMCtfcSGMakiAxHk6MEAraCO5cv2Fe/g7WtATfwccME+bHq
Zv0Jqm8hOPRB8zk6XL41nNFOvEHX74861Ev+UkNw7HqtdTmiv8CQBLm9J7qrPIeA
YFTp5CvXKs6Z2EKRi3P90QdJJE1IrHQKxjsIytTMRQly8l4gmTRahXNUeBLCi0QG
DmMyX+RDZoUPlRM4x9I3hszu1voaHWviAnuhLC/0WVbvnC0ixTdwrb5fGv0mTQ4e
t36CvTzHC9kywuinjzctCw/o84NvCQC3tH1JZztNpar4fJdwQIPnDY6az+fZM/nt
WDWiT1OWpY45Kk3LIb40IjOi6BQT/JW3i9cvEVjnv8XqZrZHSORXNYLqJDuhQlGA
wX9hGi2iAb6O+rsNOmt05z8AFf1TUFgJiOLb9BvBoZ7UXQxIIxdPNcEaHMNtnsZ+
yypdgf7lbbB2flvj7zgAzNwGXNanSMFnYl5AKeGEZsohyYHtIinDYEGG8AnsWm0X
hw99ntx/yc1gNg91vK2J3ALbdVK3fTj//fE07GCeHuJGSlxDD1NvXlSRkl2wlPfO
46q5o4jXwtOHAiSSTSdxWHfO/1/CFtwnSrJVtOvcNpkQBpvitPz0p6BQk824ryDQ
M6DmhcGp1Pciz0f0IbtZMVlXXTz0AfGAmB66zaBxdhgdSy8dEx5aAp+50Gi25uEC
GIMk/YwAgkxpsHS3ihB+TXDXi1PoMyoMJB4271Byw873cQHD8QdYtmgFl/wdhybw
/FVO/IP0ISvobGvh7IOa+Tabh7ohj7DaG3YGhUTBH2YXLyOcfM1MvCjBmyMqotGv
6SPxF+MkcUZ0+aE+mtU+zbdSIdetM4OmUKwSJCr1GdYWXnPBIkU3joL0Tl2iiqfP
sh9OKEJ1SABjjz6MX2OSJmllnH9syOw4OO6kpHWsWBnODfEczepBh8h7AXl+/jDZ
sl4LF1eM0J0wWDnbj5L7s/Qh6aV0cqufUjOJfFkjCiwQIY3gTQnplA8qaModoA/W
zBgAuUuaRJm0GCA8Nk9Quri7K4QMIIutjJWFFHXt1Yp/7ASqikgPwoNX1VBCTfQM
yp2AIU9OyHPfGWfh9PeiCYTJe3cGXdDthqF3jPV3CDgVgbeK7VkEKhGFAl/j9hyZ
e9EuvJhqRzCAzKWi0JPErsdD/Deo36TLhXY9A531LwvPDqYqxiXKLvCNYqgoDpW3
wQwLIzTgL6KcYVPb2OI6cbdlO07muAEhEmKEeO17zm40KeAI3P3ECNJ0OkF3QTjb
7KmT4f5Y4rgsnHEldmdgnjVutJ0mhvrGIOrn6IFy6HHS2HzcWLn7llA78kn1dYKr
eL/vvQuqHdg2if2IAEJ0TiyK0aUoAsoADE4qgy1lW/XVR9m1UY6Y6a4Uhss0CcM7
mvPUBhwPwhQbsBhWaJGl1kJxrW90tJdSEum8jLLYJGBE42oig0GTQWoSPwKR1USX
5RTGIxHihlCh08GDLQC7dkPzEjyptHSJMhFRfsjMsjQQ/rzlLwRGraSXQLMXAxFB
TIhV9VU2i90GQ8/S4Uvnhu6OR9fToaMHR6KXZpBb3DRr7/gkQHaxPnsEjdDkR5Hd
w8oFKavNJp/8d2jx3B5A8x26uvwtc2M7hQ5LHjCKlpks42WHtklX5rIt/0yGoz9R
mRCSAoNHUperW9E0d2cL9j4R4iyCJg7mqdT1/CTD7NcZloQsF0l+ebFsRY2MP7yV
amxwKWF2SKXs3uc/BpEC+V3HKy7TmG0otgQZZA+BEwKdMh032sk9nxC/muTUEd6e
1xlGP/5DrdzSLEp/CoHbyrrUfNQ9YAb06jVkzzcE555j62g9wXRUI17RigrSnTmW
2ALMbE2rEDr8mWoXvgqyrci7n6+ZVtD1SekAkgkmqpMqoX6oKj+up3A4B09E75sf
tKq/9Ujj/B+Fpj5q3kfIiv3OTbpWUXm09EHJVz00U9oOUwj/nPZ3UR55EwOQ5xII
QUi0L9pXSWcklQTx+exeQdinNAb0mD17cLcW43dhOZtukDkt0bp14gHQh+JtmqBu
eaTASpf9L9w2U+xEBamZmnJdnlYsQqq1isx0fDcKP+SJiPq3vPWYAiTXe3COy43Y
awq62x/T/waNBCeJefpIHvSaB6wubOY/4rkZUT9Bmg/5G9N9rCXpOB3FZG1B7mgb
7IlHzaJlO9sx9rVD0/vApou/0lkR3O2T9ljszIL7ElI/Gam7p5yaZ5uEd1jz3JJv
GKc9aF/VctbxyL9kAlOpAy/Z6+dUKLqUJscW2MsrZ/WzQk37ZiWPSC1Nj2SVn3lm
eLNontTA40Vuyg7T2WptFUqF0YVYky7kODcTEx0gZOZpBlZRjofBeoT8NFOcHA0E
xdoHV9qUMGGes9yWO3SRl9B36vXChobRkZPIi6D3/yk0KKwHRX4gLN5nsiX1XyZ4
b3jApDHPUKSA3Q4mXgnkekgwlX3HNUN1xAYXDD8OxM9ygOLUf/jaezIT8uatycFx
nodv0k6u1cI9TflM849QWze8ZJgTlMc+xYhrbR6vyvS/W35Wwg/0EoOM7r8GGfpR
oADhmIS7BNMJQqSQYHyKPpKyPuIthsPPuH1imECuoKUPUcD651lezLM/OYQbvjHk
zasKkV5eizhp9AHPDWnXHt/Krw/W9He16ZJXix/AMImcg/4qvyRgB/FV4gPQstVv
cWMQS3OEGRWiHTH1fPgkDymqByqT+JICrWwZF7Y/1o4iLeAZ/NOyJOlW/LmelQhb
E5uH9xtkHtVnnzV6/b87BSrosdfadbCnsqv5gjH3TJ2g2VKukilX8wzKEZ9M3hlj
UNEfq+XmHkXyBUfRJe8bDfuux9JHJegAKHBZ4bdtfsqquJF8wsdOUqyhuxdrXE/i
6jpeUQmmqBVQTP1YwTzG8IGLvb3GuTrYQLbX2g3qKq83vS1gUF2ULjgCQP9788wn
hKomq0BSz4in0+oThnchTcdkjO1QafQsuwmkTAA4WcXuJjebQxUkCKP9c83uXzbO
QiJuXIdZKY28+l98OrIdowtpCZ9CzMxQRyjcP3RqdjogDXJWe+o4a0jP8WI2Ccfc
otf1w6irMJOeJBUd5vgqU55ACdnck9Q6ScvNSq80uOuvYGkbBKj18bBLEYbsk/DT
mD7XJqy0GunUTOK+/eAGLGQjZflRek0WXGHhdCkDJGum+coso5MHdnG5nPENYsUk
9k1Fv0KjWBDn+jIbdpguRxZ9BrlbbDAdVI1rIKe0CnZH5GMvLwt/shdLme0G3usd
UGZoZ0Uks+fVA4ccj4hf/MFzppFfmd444M8Ge2KL6jPvQZsxm3bL6SrKj/c4WS7Y
G9JqNkJprBTk6hOEW0hBWPTSInu+/R5FDwGAAn43svfD0A9PARURWMzdUeosQfPu
0KermEdiHW5dr14AnEEL+byY1jsrHb1OGVo5Nwioy7t5ZWwhog56H9PRJf58ngrF
b3U6AmHzGvWjipTak92QVt8zqRTAGJAbxGsitULkofAox4aotjCl3leQ0AMxwY+P
8XKH0ANJC5kaC9RgOs2lW+uChNmdezibYRZI6xoVJHGOsKArh40VWJA9X7R54t3b
WDqh6ASwiKUILO7Ug1OZW9RGRCxuS1a5SNsOinshswpXPQq/AVK7W/mo51cGNwO1
1WPoIvHXlHRdaopQDu2qoEIQnGWxqjs1YfZvYz+N2Va6UKTu/roK+yWgLee1Kh3T
bXuzquUDOHXJ4creROdh5XlGVLGXdxLXqSuFt7PKw8bdyZN9RMAromNhLAmrtgw4
oM9u5YWj/e6Z8HCxe+K1ZoJynft0XwFG4kOePi0SQIythZX+Mn/yDQ1r/six4tpf
cVnt5N+2SUaFsJxpGBCDe3+vYqg5LVr0+pgop5JwhhZzAaYXOvzABppyFm7KxSB5
NYIGgRctSw6vOH22HiRf3sSzNrOZBpqs8SS7FiNQBgEUpPQ8XDMr1/nfyabCnBdD
Bo26Ho+SV7GPWjf7NFcz22z0I+C/akZvzV6OPnFomLPEdjMzeLc2bjKsYH7MD+7/
bdgWAnaSL52RjJ0H3Wd/h8fFWM428kDNFRAGwkYc7McftIqIoaNuZU7IzL6z4zur
vbScQ4f2LMqPQD7RfuXwDu6U4XW1v7oYZR+DWRiv7EE5NsjiZi2HvlBcZQHKAX+x
y6LFNKxtiYp3nivuRMnzrdazypV/Qswsv6R6wsV9PCBgXIUReKff4iZ47RHIjMH0
GE82/oEKODL8Qv5qpnGOsEBSJrXuMlteKMyHzul9b9B6Jgm0MSjwVRp/PhX7PTa3
pj4y3TGzlmPP9jwN8snhsCkoZIxQ7SMm3vp+b39lFkG/aMPBS5g0m/KZRxLd6H7l
jIyF3YLN0zXigQhridBqkg0LNu46RaA6id9XdCauHkOP8S+uslEpCcKlll2Wan+q
Rwz/VsrgTTjI+/YaCuS9lmvQG2nvlW+YsCqpTCnoOsgAY2kDiV3UJ1aFiMzmDEPL
si/ObcMWmLiDbAeqxODE+5U1FFvni3jJzdz86xNNNmM33bVlH+eJsARPynRraD3s
psD/ueMFeYcVdXxdccnHenDSE76QzMCnYNiC/5kHQFx037zo/8zwRJxeVAPvOzqA
UD4KyZadkSytkgf8L/qfwxzEobWg4U8mvAuypbjrSTje9scA1XSsjD/lWc/ylG65
9HZ880ihViVEsOpyCTw+iXgMFl57Rx0WxDxIJnbYSM/9loMxmXxSK8hlZOfvBFYY
AFUzqRRXEu13HQmhCDM36QwLEUGi0QY6NORwCNKP1On+v6lg6RqLmtucIcS6ivrA
JZ4EOIujyFTDTF4GkfTrxCn4gCb2Gf26NfAxQK/h793qXI3w8HiKkgPSr/RUq6YR
Iw2yaP418OwqOwYwBUmaZWgQSuj0vgvV5WtOwXYx2npsPoiV3Dc3wPlIreP7XMHa
ESCZj7Kf7Cg5KxbHnLPQ100s0sAmQeOpENA3FVqaHu+PpQAdR005zBHGFPPdGPlP
VX8YeiwXx2yef/J15E8wYgFASaiCJi6ob5Kob14Mx5DWevPZKqicSXMMrt1/Z72o
phs0mGWA+Nnde5OIzXYgANxYz0u6w0AEROqrqWMinEQuBPlwI5cqVzIXtHZoxIyP
vRMZh3sawHw5NDnN+KBsmvfdE+TFIwcTtNEZP8UrWAh2ifbgDCHwLEyY4LA8S39M
3OVZI/kZwJ1gs9LdKRBDfBIFwdbgQmBP1n3usPYjqorfwMzMF3inOenkC9qTnn25
IC8Gy7hGbfYvBmPkKqgpNaaWMgT9Y+t3l9WENLHNBwFD4Gxp4j2gY48UX/ViQt+Z
4PN2p20/IQvBjYw9v5gG3m5qOeO1lO+7wCgYcdJTnieu07J0H1r2dhAdXSgnZyIM
CDzHXHsdAFy3cQoy5DpYoRzvwRm7hCHG3k9Cw3z3wvxrkSY6tTcALM/BdDNLS+z9
0j6+rGe8pLLSOMzSydO21m3+7ELa2QZJUV8z6NudH32ygDXAme7UqTigOmEKCgPI
8p4ewS/VdWYU9IUva4o87TTKZSg7EZULvttak1PXUig//MGutMmSBzSjNfc/8oC9
oIhyO/jO8y0H25xsxbRZaqDjOpSx91AaNn4MR+CrwQzQmLOJjNu2KrDw9Ej22v4d
/wJwmRpNQ3BTk6sBkp5ua1Oq93ArUyoIPNZTX7C+ofXAtFRe+YTRBV/zJSQAg0zC
RTyx+7wRg49ON5wfKSKfWZ/379mntqmabiEV3mvaS83uEb4qq8Wnw5sAtZWyiVeH
kTgr5/jfhs8N2HfeGLTMdcjNgrPB9imCJQKYziDBO5kpwmo/1JukBmU1jkbdBqoz
23SV2KfIO+oMf3airCZ0WI5BKcThahhPMgBfeiX/yrzCPYbZg/fy0DVkn4ofkwYs
5BoLFVBPJOU7eoYwH4QRCdB30wL7O1uixMH33ImXgC8Grk61JaA2M9/93TlEswIq
jByikk2iuCc5dy5ARUcIt8A+BU+aqZUYA0xHJ6hLViv7d1tl4Kn+WDeRCsN6BVQB
STf2a+eyaAUVHrhd1jwN5yLayxrTonEPKdgcITLxiSibysJsp6J4kENBItoZWzna
52KYtaWIX1/xMNJEyEOhJBBoHyBJtQXL3PUrauXEHInqpBJ9xLRSlGTO8IOSJIPJ
UyvwP9AufD8hj9piv7JltPTli/sDKeOe91Bme5VYnl325js4WO/EUZ4FLkWg1tRg
u1DqXsusrSGnn/lHUtHy1/39dz/dzBM8EUsKWIn5eB6KTQvYR2mb4aXcsiATGCb0
E+QHapLy8XNE0rafro3XRFSjZjwIkRsfkVdPNxEDJz2MuiePh6nV0IkJh9jwwDSA
Q1JOkq2wP5QHBGZ+lqlx16X17XZsVw42eBT2Mt9B50uYGScmCmHncT5lBWWopL94
TnTzRfEvAGMIvREZiuM0UR70WuSZRVdXR1/UNK2NKs4bgJDxfal9IqTTnM3undFH
DxkzsIaMyBVN0ixPjY6UuTaemMCO1rzwIoQndRd4VUoDSI9MdA9ADxmNW500lLW4
kYlzcl6f4u6AgZYgkTcjkiLSoXZtJhkTgWvNDc/f8AlG6pa5UXus+EoTNTb82VUe
zdSPbrQgYh7cg1CByHvuhgEPzDMmAq3SLx7O7mH1tyIrKl/D8S3fpMeUfM+seiHQ
NpKDIy3WDZ82ovRvCXy4ZjWXj3OsH+NIyVBJq5QR5qAo/577+LIHq87QGKPuSl/s
qs6ISKf8T0ea3AmcaFGDzCId8bXXIF+LzRRYYJkMjRfo4NJTX6bg7pIqnPuFF0AR
lPOqQweydcdWYLFZqSBUccFxoBLWoZckCV88PYz4IiUrWE4KzFLb1Tqv6glffoie
es3lgsHPBuJ6NfXYd8Gs6rMHRy+aPEh9fequZUFJzU6C4XOFCriDMZIp2KJJOlBe
aUbOPqOztUp82F5r7TroBsNhHAaye0adn8774oStB03aYFzx1ECvS7/eO1zA5UWQ
r+j4gUi4iIdUP93yxZhbttwseoYRE7U7sIoz6YBhtwVq9a0aB3ufAiGnZ+cXL/LM
JaDwHXxXqqIV9RPQHuZu7c6FJUrbXr2L1llP9cnjW+1Q9sdQZzBUnqgCO9mgnu3D
0No6oAIeKUOqxFEaZQLpnh3o9v/H0VNjy5thjXOIQ6lViFueRuWK2d1mdWLO4Phb
x2KPUqa1bWO4ta/z8QdNxyWZ6CcUGwnBBTHZV5T0Y/SkcIYaFWS4zPSt1JZnAz1o
jxNz5hW1HT3Vpdn3oid18V25LhJCIVFmFghYHsdMdXWz/8iZfRUcokli1lXbGAg8
gSg8DkfR2DIO6rHqMeu7Khkdi3T4kp2AOxWybLvkDfgoennMXFvhIbdtQkvN2Dw4
uSOIR2JCJSjVRuWbN5eTEWt0xD4ScOPLOMRYF3H2VVhYhSSZFx8PSPclWCByDoxX
akVMccnaT/FrkmoF0+1+B3b5dHeP+JydQxo+O+dFdkk3M1Ga66uCgNl+r8pz5wRr
SMTBA6g9UJG0d80Hm1f4ZJk9l63woTPTCCBJ7HWWa39Geu2wxdths+Yjffym86pz
g2o277750IBwX34k862Ekua+HCckfZAy16cGk9/D+Dkl2dd3dwFttnExYIIIQ9l3
CYcFVQAamlj0rUas96R3/IeAIPN8oV/Kli9k3j34IB3UeL1owdZoXyYq0XAkTdKc
B3JYDK/5loDaRoKnNdvIYyRWaikR7u+/IcNn12lcMD7wAtz8YAosn02v38DTty+o
o9NAYx0UTMLKtGbtu5M2KXQh/SFi7qiIPgkf0ss3FDNjJFND1vgpoSa+fjFAoq4T
l7JOGbiX1mEcY7lO2tpZX0+Rybr79EWvi4j/OU+UlcDdEY2GnDQy9eT2tIkZytUK
b/90SEM9zRZ3jjd8vIay/KcaAP+XPJNBNhIgOmly8l6qkQ8e8mr8oDf+hML+nVNh
Ic08Gq5+zxc7UIk111B4b8vhty8D7QYNrUALQjzcyTz5ZZzUBKLpG+IdwrmNudtE
TxrtCVM/9nVOFffKw8YYqVZrR96wf4NfkiKKzQZdZ1ZyKCtQe4iFsJQCkE9FyM1P
HwFuBUNG6cKBCK8r0F8uJKn4q2uo0vGlKnKZFTY2Kt+uGlGpPE4c6BoddXY0NiyN
Nfwv7ZVWJ5bfYd4/ykyc1Tlkk9hzkehdwXpE+WyY9G5QdJICUSNeQQVV77g+gCcF
4nJUob45krO6/piJMQrNsdOPns+IKiSnGKLqAp0ElY/vLTYqFwxJDM5kEu1gOnys
7WoIXD3DqdhhwhF+VPwp1HUq2dtUDLLTXGPET0n3SwR6v+SV7dTShKbalR3IA/08
PhSrkJ7WahfUARDBL1CK5Dhr9SMmQGED7s943Ce/XOQIHs9Gpf41znf3ylYR5Wjx
ai8ztStTfEaop7H7cWtkQx8XR1HKkEQIP3ys2mPrSU8FmPkd6jG/NxYSUo4HxSFF
fIZHAjptQRtbfsTROSI62G0RkE12G8Q1I7HLkoSNTgWcgYtviPt82ul0cv7JQiGz
78OS5ju9Hdxq+yhLwVGMh+ZHZCXY6mVlVU0lzaRlNLY7RdTMe/de+75L2Cvv3E2p
VEsPJVAkdYosHHdlg+mcpwRXLM+e7CmMkeFu45+SYaw9Opa7X0xgZw0mLFBGhU7h
WsSdIUXyDF+2LCgCOtmbUSfip8UYQ1uaVMbVgQdQJc+CSqZOcrojU0YPVBZaEmUw
qCEHkXVMoQ9Tr88NPVmMHYO2IRlzjTdFtw8kgJb2XAs7O+L6F/jN9Zbq10o7x+Ps
FmCT6cgmkOw142NW2PSQjM45V3h/DxKWlIVVROUWQpU3PCiDO3eiL/URaEyv9bU7
Sb0shfCXYvIJMuXJq7VhDag0xbrTE37Haeoir6QOF4LHl83eSmGuy23AL/WPJu0t
0ay2m885MXkLydv16NTjbgzaAUqyt6vLC5AleIpYmfvagwDe14TRfKPYH62g28Zx
JTCHILRf5Lzp0k/00KcSDUikG2ZOa76NGEJCQMHaDjbfKid6RQI6+n9HCygbWoGC
TnXhKod28gBhQ6QU2zb20B9UoxJalyQ2Y8HDDA/RGes0UrZ9k1qbfqPVTqtg7x+E
RiJ1Siz3AbLJB1Y9HoqBrtEuXAjfJIasN0xfCnNRVrNc8E6YCKe32OW9urw7Qo+E
kx79PqSC9zakK+OVQIWaISQ4gRcusemhbikiQyt9IiHgyeYPguyymVCcuFKTfg0x
aZUHZnEgq7OwAu1LU7fPF+psjDMcXavPacQ9/b5W2dAmPdKzJzC+pkcaGa88oJSn
CnMaU0GW8xYNKYcfFZyAOaiKv4y+7WmUmDPlAhflLgRIMBYVhdaZcOBtfbLq7fn4
OXePkB+YTzxHYKhxNm8BlRn2e9r7etiWdDUs+J0xAePFS+uZHiC9ReyW2IREXTwG
95DZLuz6ITbFtr1bJ0cNUGSZ8x6mMWfwF1TP2dDnWwK/yQ/l//iMK4KyiuT7rnfT
CJ4edIxeZvsEwBhZGMB6xn6aGk30A2xNAW2fEOXHd3LZ+NMW0pbyRsd4T3UNv5HP
XvoQALN+g/U1Whm8E0xW7wwGQBRdSSnSthvgHr5b/5d4FRcgff20YURD/8k6Xi+T
8c0n2kH8k+aRRYwnvRr6MbiL/jgDugF0O5RR2s2nIEpDh7hkkaVe0YlqrK7HTJEB
Nj5eUJaz0y/OW2tIWuzMAG5zzxD2fHDYhLjP7GM3cy9TJLsxizGlP2gE1e6tMgoP
5An1NCCiZcEHLczbpj1+UWw2YZCQWmdp/yxx98pkLh3vM/i7CoNO2qsIVTZaqjgc
1pInrUObUoM9xHerTCv1Q91fD1jhtPdSj/m59Voox1A8ToKG+z89G4x3iBv4q8jq
2EwUmVkNQPeLOUGMZABOXkHYOw85MGykAnUQzpQ1rRs5Sf02eSqBXflBnIGs2mOc
DaCXIB5eDsS1C0a2YGPNQD2ZP61STw53jXDWGGELJ9UK43vIlJGgUxW6873aJP1V
AihX/UmoqTEQ51zmNiGcX5pMuXGWCLqUaqDhmtV3sV7iFdZ3r3MP9KGVpvgoDFAF
3b9VJKAi0gYwzouOVI3Z3x4n5cmfqt4Ar3Ycecp7fJ5MAs69Xpx0WMpodIvsE/Z6
zkzkzfygSiswuUNcqPlecCRrtN0p/WM8SMjwGefOwijaZtucRaZ4OE7yEa6CeTxA
9L0e+vi4JW2CYzzeQA+LyetaiLNCXAYdHE/TJVcH5kI/Aq4Acwqoy+yzstBPLh6r
3y+mMW9dK71+fQlJ2/b9sxOXQNPmmQ7bbHhwQR+lxqUxGS4ekV35Yz6fjCzAqO7T
VCJ1dJ+UG7wn0ofjCXAOsN5Uzd/PM6DynNQT4jKHTck72tf3bI8LaZPX8SYM5UX/
QdD1ZJGJMc1O3sFqVeHbV9c3uF2c11BRoChyozQWyMQqDl/mQjS2NCWTUPDKxpCt
h3OoU7Mp9gEhUh3dxDFZ0W1jbtcjUQ5TE5l5tXdn4xOnE6+Zh64oYMt9R0vF2acZ
/EWSPcicsccPhzeMbdlmRtoYioQCewRURB1fl6bBv8+SfjVEp6yP5QMbzSN0JyG1
dCsPVeLRCNWN47Blp3O9mrEy1WSJwZwnkUwcg7c89eWGxpXER+CJm9fdLa1mrWaD
kE8jTbOAmTTzp7U5GKReRfPZVfkJdbNQd7/o8z3gjQSil3Lutgf9gKdJh6A+Tgzf
5HHHKFPkmDsVZYJY95nV5fjjf2UHiiLRnjqm/f+HQyQKTomeCmZQrmplMUR0BwvX
MjK+/DCYOrrHMmQ0t9qGbdRB/4k1MHA3EJzQKbHHP4Z2YzVJnyTSQnaDfQKkcT4S
0ibhMZwZrdxdKG2homUYAeHKtaIMl0Rm1JeOXs40N2h4Yq2A2qeY9vW/8eaTX5RG
E5YlUf2O9riD6GiazUSyJuSrkPdVHehboe+LzC0lCDudf/4pUsAzjEdoL1VDhJjr
StAtgFEVCTKwWpKeycSx1xATiIhiGQhh6lxybg6UCH2lm6GA/iZ5gnWymHcK+f1L
cQL/pvzpzORuEbi3faPAIOv/VQh7SlMQyiDguQ5yYItMnS+4JxgwaMA/+H8P7z5k
xpHLPdLTg/BUe9gGCLrOm3b1fUGgJ0DA7qa0LZ+euXE8w1x+FpBpMYfXbuewS2tK
7YVU4hTczR1b4jGtZo6CD3juJFk6AT9decinWS6ONqte3on/41MlmJUmOlnQYcEw
J9gESDhtSeuYjDsC9FrecRjnvyfWh5JMO8qQ7lXf4ejC5VVgWYSP68tp7PMW9f4m
iry9xnRmLMOw/tZP6T08scWIS5Cj7jPs4lLkiVNS+iMZHSMILw2p0umup7gUo9E/
Zk+qWIfsOfFVJMk9JzFfDdLrvgO6SIbM1JTdsWtK+psAfpVKs5S5NIiGYnwwhw0D
Og/Frha+4R5fkueCaUcQ6hHYPQC/UtXSqGppNebHXarRfUKATDQvq9AXSjjCZtt0
IbN3iNFeIPBv7B1wmxg5nTCcCPsrEKN4sGJqGH7a/WEbAMo5i0hDE3umNJAvCwz2
xkMGQ7PI6Cv0CBYwqap55wmG8sbh1KsWQq0R0jZgg9Db+OLGWvk3mOq7EdHhhxEi
Whe1qGNGVvHQf162KSmWzjRSa8iGKjqt8Y72X/An6V8a5yvoVTs4C2SkwDSa3SAZ
q7pNb4dUMTp4ZAx/q8++5iEhqX4PdxzCkwbXH6UBhxR7nE1XCgTkjT9K9CLhuHlN
dARKNz+asOs0/Yj0CO+onqys3aYh3Z7WJ7vQbJ4YsmVGDItvzsyl4PDqufEQotCn
lRN7S2Yr6rmUDoV2EVjJsFpDMSGR0YlD3AWo8cDod9ajLLxtpM3YyvZwQ5KpKLoV
FUwfT/Fy5XZHijNKVsd0PP8RTdvqS7pnTAGNfEwt1diuJ7B//KM1RtkSTlVrHtj3
l2Q/6RFp+KAnxvbbQgMPscIptFlywUWcirWmUbesW8g7jCeLqiLkxnXrQJ2bsTfL
ZJWUN0tBBPSau1j33mfTiVvSC4L6coamRzYi3cgLEaxABAjPxmn2XKYo80KNamfZ
O0VA9Iz4Olz7w81jt4WaYVvqe5/oO5iAcRsEYgM9RUI9eNMuHHe7WcYbIe5UXFaX
7iKA/rocjX/pNrkYH0v6OvLGgn+mfw2QB56VvlGzzNSqZHjqiuAW7kKRWVUgX+Z9
YOTnXw7yyFBIqEqhuyYPwK0hmNfyA+FLEa4fVaLYJtcPEmIxBFcjZ2KrXypbCidu
+1zRk1wobrAWqPdcbltzpt6UzYjmx8dc9ixHhwap1fKa9/dLBDwSQkPJEYulfT1T
ut9u+iGDHVUJTtjL3hd3GiB1Z7Q40JPIiurZ51+vXNaW9GF1siiuWLtUAXXRQVJB
HBzEPAZ05O3Aod4jJQBfPzmCWX+bHKV5AvH1W16yAZO5slGZA86LpMUR1c/rnqmg
7M2Fo0gscnKJNzVfMH9cVc8+fUYqCTlj3ljuFwOVkdvRmsc0tVhqykqfVRkuJzKz
S7FOtSlHtQogw7PZ069KfpZKzSdwvkaW0/+t+UbmcvcNb2O6O5QT+1KD3rM1NbXh
PONCJd3qFtbkbixK31qwFskDfF2dwssmYNBr5IjPmhPOCX34Wen7FvFeMTztn1sa
K+XlEVyrll5YNoTzYTKpirm2Mfpbud2SHb8GID0KfyGTOqf/JR4qBNjSRfrIoOv2
jIBL5e9fjBOPFI1LTZp2ms6p6+3VvExpCbrchh8gjLOHlpluvCNSjYnY2+BsTgEl
0/M3tThEe9rBbXGIFcpbWDSr2hCImaf1rmnvaCTJBTDb+jiPpj77yYVjZfDoFB1P
kCD0rMJZ4DheAJLywu5AvEF7P0/kgeWRKTCEjvUIT6sOiEk9lJkj5wzjpdfyp5pM
gn0A2aR0criUeffmWgRDIBzq8CRs4lzIjyMqNhGmi/3mQMfG5E9zWKQ92EtB54qv
4809au+/Wb/DaZpSMIo4L0L9TywqinOWpvrfGDuOqcXqga14/YuvBNgQt1qsY57C
xPIkJzrI1/59wTg8dVMcd5f8e+UB68QUNuYhSBQnVsLV1njnhCyprIuTF4NQpMeL
XTE2nSOidq4M4qVPpzJC+nRksdQ6syqJJRwmasmgeJxYgM/ArTWemq5eiDqippZj
/XV0/X36Vb/231kdb/Tld35+cOmFP2ymhpLtvAlCRcT/Y6+Kfck8hseMwL/mYF7A
B1Qx8EXW+wR6U5XCP6AY4rCNO5nevRZU9e5DlMstl/373wMzM/VUekb8CGOMFiKN
l5pK2qEdvEvhIz0q0RVByhNwy7cdKac1EqRAhkhzABTpfrKDjeGi9M7ymbKnseyI
OEdFwb+Ga7oNNDFjyswmxnD9ckIimLX57RXUX4MIwPw7EyonrB/JBRgRFI+R4h2a
0+OOLazbHhfX4eXFtm6eTID26nDUyycw3ZDi2Nif+4rzyBgSfyyy/cKXNHMBOc4i
AYdcNWWJYVCfmkJU2boJr9WCbK5Gf69VR3COHtXp2uOFwiF+251P0HUvZ3i0CXp3
h4l76citUDELkjVqrqFhu5q3dBDSSlZEcMThoz+2vsI4VL/Ell7sZTW7JzyCfFuz
ObjmpOdnOE2hqUJv5TWtua21XLCNQot6ivtDxo68UyzuI6D1o5oNCdbsrKA3b0Ck
0ibUIJ5BWdbVTKsdvsreRCXDYvS23axRhHU2VlhqoRYkpMlH2kqgjRb5IrCVUfD0
9IHLlVfh+Q5LhIpglnSwAWLLAzJaLrOmDl79hak3oNtyCT0SKB3+7+Q9v2tr4ie6
JPWWK5rCA++jXdzYfqMXLnCWd7ljdJscqMTbmTrU49BPkft9h5tpDYMSp91WR5h8
oqBYlKuYgBE3xBygPUXJh8Q+lTiWhpDtGCmD6pxt0ai5sWQa4bSu+9v7bZzmcQuI
PfyIPrJ3Kro4/ExyE+I8PxQAkvvhUrTq0rChiAPUHzCiY5omthq8YvX+J+HJjvYM
XKumk0myUE8Y2XDw/c0EscDTTNcO98BrH6rswx78fzewT1ucvGiP04oohJjoV7hh
f4oNJdO7MTOphH9yoFlqXPWI3yqbvd/mAd0iJ3o87uG8f25es9ql9HUqq1U5R7XB
ZGWvNN0zse90od8Lybzfhg20EiilLNHt1pYxcHo0Uz9XhPSMxy2Zmcv+ynPXEg79
3sGx1YzkXuiv7bec1WG1/mF4rRFngmwgrzJ70WClhP3sELCbCEVNvfCGsEohpgcj
I+e1zmDFUtw6dQixlk4v5rsZr5qupIBwDdxO3v+A76Xn5fJw5/r8+4EgCDy5QPhC
I9b2trMiDD/7RliZua/xPraHhOQ65WtBKBaLC+e6mDsWT8+QhYvXrGzvleaGY43E
GcjZE72SKPtkqeMq2+88oJCMEvRANe+ChjjB8WEWZ32gSp4f6nCWm6MJlKKxNUtP
xf8kAh9fNbJeUJqLLwbcc0GwnuSmT7Myi6/5hWtF5aHrGf1+DaNTFQRCgv9x9Pq6
IBeZXp/DaMmW0DsF5Q+uPyv/iqcm2pfWw5G8NMpbabtw8cfnCcc15VvnUIOvVPRs
x4fOQVDAGZKIP4zsBIw+j/DgreE8naOSJZEXrrVruzs6LhjmPDof99Xuhm3Apm/w
vR1xlqqQviV7PLIPop875bAicY06iJK2+Thiozv+NLCXtFmH5DvTLO0qrvlKYCae
Ceem+9X8CDws/SK1arqTmVd/pYoCtj/6sBhFWuO9C59mudPLk/7RtG+Zhsd2YRMn
S+50yaoBojMfIVjBv7XklxpGQHl0cqP8Lsv9qYyBiwa3dApjoSRC7AB7EG4QXa7u
ATXKRYNOR2UxWfQNmBVdhsMX3SDTdk9ERI4huCFORbBRrxGOovi8GuWB1H2pfj4T
vbSCgnemUVwNk5oqZyw6zSSZA6zEsNpeSFWJu5tqur6tAj3s9HFOQVP5Pk6mlj0x
USSLMxjoWWDuMDkp+Ad7JOxPuom9e5yPWivwrQsaqa9tDcVEO9ug0mQ2Zz2xVQmQ
kXU1RXAiPHqRN67w8XCoCGZ+khd1yjvXvVtghrxb+opXBXlGzEkjhr6o9gX5ciXX
uoZJO7IhxeHiBfVYkvhG8RyIYDJvYV7U9Kf1HLsBBZIX/3EfLswFch+cTvU+u/F2
vpiK1Ub+eLpYP6sZHSZ6TsdaiyL9wXsu60qCO8RXI1S+SWRh1nPtlyoG2At57Nk6
2F4RdrmigpTjOXEOKjxJpIBDxeKiKPsu4eGrNKmSmpwXU68gUMlLey8e/Ik6BYmB
FOTohA1SxNZakevi9i3eWaIDoujlDlYubiEHNpXxcObzMNirVMelom/jwRz+LnIk
z3zazS7/piIFFTF2xGDqITh6Glalr6hjiTjcgpffMwKX8hryVNUcYPhzAB0J5K5R
PHuykd5PLdp9VXdOSC1EBW3uXYLuvAtMhLdBUpnullwPsaKy9knc4T3dtzlKMRKd
RZJGnbE5hFIe204z+jiX1PSKJ47/EKYsHB/VLK6Xqw9uiQyCcfY+8OhecYOtUOtH
vMfhSbSwFcp/hQOARIy5xOgm0NzdJoL1jnnOeR66BEukDFXKRGXelpRBARv8HvXx
2k3RiGzsjQ+D+jf2CpnIGQ5tEG2P6NNALI8EuQSWFLKsCD+eSRU1KQKKGM9BwKwz
OzYKZBb8PkjwXS7ylT6Sfgi9TtsgFP8loY/giBKdcyqAGvf+vF4gVgfgoQwmqqBY
P7h6hzsQyCkFo2X/gB4nNU2pBwsY5bQCei6ittKMxaA/5uTsXpDQMOCVDEt5RaXk
nU1i2h/AkGf4lLR4OIbNziOxiN0aQdwrabRRHEvuY2wwsU8BJCYa0WBt4lQayyYo
GvicXiBYcY/6W6xBGhc9FEsqvZ99BtlI9W9ZluWheXqL7RBlzkySsnWJyD7OxPPn
ZFLVzHjHcvrNHTZ4yM7OVoVi4AXoPHU12UxPqbVLDTh73jHa5vgY2wSSY6t5UTr0
oJgSuMXuTz41E6tX5TZut4KBV+DemdM2qh/tR76r2MnksmzJrJ3Plw2IecjIdy1G
bbO+OrSEZjMqTNwo61eDadz9A5+WBaAzLQ+WuAeQ3HscqZ4LYzUyUyoLjNdvXig2
ocNQburaGH5vAe+0uZc/g4OmSTIySQVBExS/061jdErrGqcZS6cX09sUllJM2/nC
NPaNzEXIRFthw6k52k6QZPiil3lPtIN5yYWj/rky0ybLo7HS/6wN+hZO/bPFTGy2
h+PGu/5BiGPPovCvKI8KT2hBrhnsQP7uNAUri/k8Yvuc4lPf+ec9qveDnMGdX7HP
3lxemSLcvEHoLm3Peu3g1ClzfEIm1zRZzH7rCNcty4ABqkwjYu/thekriiDBMrsZ
/7ppPaDV6ZiMp94Tmp0YTPeZDJDUqZoj12hQ5gy30Sf1V5A0r5ENGrrRn/WPqqxU
S0DwZlcQ0Q3+TINEpQj2+9TmEkhmBHCCSHzufU+BMtB5Cea9+mzv7S8tKchL7R0i
IqC0ZgLKUwuf2ZiuD5/3/l+ji5okduz058IXOaqKHmDShMVsA/y5sW3TCo3m92+p
Xa3B4XuEozQkds7H6AscK480sxcydk8cUfONhubT/M05LZbweovQpQMkrAZa8gDX
lKg3RYdYMrVnvJcuy+JbASWnypNuYVzHfI4+ITXceXorTUc2KynnvQDeGRA4iVwo
rfb1bYi3sfVuKXV9nJofVLhiVLcwOoNqf+RyYAwtzpZSV3G9MRIf+eOy1rvItL9y
EzS8Ara5gSnxu4gYsv2+seCx/Gb+fqrHnaTXvCzoTtPwOMmo2RDFDogrwJ64yBLI
1DlG+s2uzXfsanjIZsquffV6ZIuaWKOqClz05aYevW44ltFSEbNvpQ98Vod1d/6K
KBOIbbdidyQTjLkiyZcvaQmxdR5PYPNf1P++nfTE0v4cP2bVNQdIoSNGy0WjPpoQ
7kC6EDfkHpRbIWwUxoQpX+1JoDfmGhvxQIrThpq0MwpXqEUU1PtUShKlZuDZjK7h
gHeltbgRcbBFbPzBgQot+mqf0wpnCG/Q2QPZmlQdIyDhCfTjOPziQ/BAOxa2alHg
uEFLlYBFfKXwv18wVcDAPlXaXJ0ISZf5tV1qWhVa+ncL6Tw0ZPuovGZKaQIikXwv
K/ZNxYnUNVHwy/lhMRShOpsPMpRh8OY74dwbdTE3B73r7Z7hZbOg5lZfrWxTKd2o
CrpkitpxIcRBiqXCyWmkJ9BlqYCxR/MmX3zf1YQQBQGkr8EIDfXIrldP6C4QrZit
pp8zZ1KcAQ9+2Mstxmokglbxt+sHXCbqH/cgFuZaCHRswUK4GjW2kMQhzCo5se2z
tZy5o+E34n8mPDyiEVQRDDtBsQBC001pxe0tMdBIKYxNN0lGDaUZrTfw2Zr+gXOG
aKMbbvK0GmUCm/STgTJH/Q4cbxVkPUNVWZoP150/7cCG9BqR38mX9CZi+3zWglOs
Lwk0byrvxdlP9TFIsr8/+ed9MXQWDH/0uVzXFu7On8e7qror3A3/lJXZbjQb9CPI
K2uRVYkCXbGAjYp8Je6yHxrkSA170d44NGCMJCsQzw5dGCXJjy67+a8NYG3VheMQ
G7j8o54+wk8xuwZdhZrGXiMQSyCX6fGnsDEEpogaopqGucBwBjTZWK5wPa5bTUfR
uuiGig0w1sGeBO+pgmdsBSRECPFYva7TFXxq42UVipPrS6gROq9JD5osbI9pfiNz
QAHsOOfd4o7c0sFiBNGHmsLq8ugNJ8YvlXE0IzCVkYGpiC9m3PN6avHzBkfniCzw
QGnhpxVLgo5V/v3tXVAkDSFNHhTgI6b7W9jY31hq7wiErJUJ+WSaIr0Kn6oP3fs/
s8hfPZ8VJ2t/hgDTjERboH6FTnYvBbnwJRALHvm5zQakVn3ie0dyxXNfACCGUjxS
Fhcpv1l7dnbX9qa06f9mrdMh2ejWIv4UsBU/GKHrZVrF4vu5hlLBlkitVMG+uP9x
2I2QQCgftAYBlu3d8dcHeQ3FjoSXrrNAHOygPpW+igl6nDy7rMilKQvd6i9J9V5J
BOZDFKVTwPlKMTgVkraVHIEUwhOY54/0YMn73NxP5ZTZ2BYwYh7EJy/6R1FGX3Cz
7j9rOQ+Fo8jWnTQqZFM2fxSX7gY5r0BgeWmXOxqb1lmmAd6oOP/K67JQQS1oSpyT
cTtxOg1u/VnqNFANSdt39Xj35/MJ/IjOyCoSUG2kUBjVYsCspk+1q81Bmh7enUqz
KxQVZHqLQgNDWyUe11Jc1chogj+9b+Ctg52NyMQJdk73jeyXQcsoLgcniLRcAFcI
s5frfR0h/0J6I4lGP45CzonLz4YABbUDCEN4b8qS9XjJWMc8ti4m6JRbiDqsdGJn
aPRsuX1/3/K5f+feyphF/kskzUXHe7YKpL1z2HEOOsMlyFpDqeVYo1VK5j27+Pt0
3UlXx6M6g2pUa4JfDaKIe3sS8zOtu1gDmYJAgzvkN8BGOztzDBxERyKMpSKz5eZ1
AGknm5JGS2uk8cIrQMT9CWxOJL5f67EsPViJ2FAJLwFAVYM9DOp0fj2xsFMnG8NY
W94b7tRNoz4TrwLQBB4OL8WRgpKn3ubC14NRxIM+4gw2epoPYcm8WqHyJpXtVmJE
BuvooQR+FzxkSwJayBLIysUrfDwOSiC+iCW23cSM54BH3t2XQJO/0xch5aLnP+07
PSVZQgJQcHyfyVX6qfI6pt6gWxtv2QxTTidCXTv9NuVpV7F6QeeabWLHk1qMI2VV
yn3vP4FU+IeEwlfeHvb1wJ6fnumf/89UyQpnoCQ8j8uDMvilzxiUxCNRU1AjtdYJ
t2uOO96umvnWfKXT4AzAlz/oNjsAyF8tTJc8ZAiUMFNSehp553GUtNWiAYFFY63Q
iayFTw7CXIDGzUXNSKSKq9d3DOE37+7lhjXodSxKO8qZo6PyD7ZLHSDq2SeRM4J1
60X42QBjBrDV9B7A1JRpKzava/bdlZNPy9+MYjrySEmQn7SY+g6PXyDjWZI0u9EB
4vqr6M+WkOAam88KC4e1SsRir+GUgfv4rqMx04vibHr0hJgXrRob8ieteSQRfVvx
0a62HEL2giguPtrCQdmH8WW9ujicyS8shVAWGIWUFnVfVOUs5OBGsniwUBSTPrxS
WqpsCchybN0Xijk3dryZfwJfl56ZBTz0mz4FcQ3Pia/cC8i1KuT2Rk8j9xgutV0H
8Vcc/EWUErjqkOwfvpDAWom4l7Yb9ijQwEtGNjSHTNF/7uQoaHJvL3ecuywK+PDj
TkLyFPYq6d+Zr0XkSwJ0I8Xx7LHGrKo4BI55OF/UxLyZ4pPPQvR2ef8yLeVlqvZY
gmtN2MqUvpGIcVcxUMdDm/uX5Awg3hoswdnKdn1i7dGn9hocsoW9Kcm69JpY3J6Q
CZJBvIJ49zG6aBa4/9VDlqm4fWlROcF2Zfs0VRzXMPyelKmE/N7dW53JuHWl71Sa
MpmM08dF1RzlHcu+zdH+1pFqk/Jp0h24MOVtr116u9cY7Wuj8LgOgoPHsK8TB4No
6GTToXnurxNmvG/QdULcllk7xS4IcSOW4xj0SkiYA+S6bhfFPYQHtLW7Uuapy86y
nvdZxFERyxRYOEqbu0u6mx+JM8c1R2dc0LK4WqqO38EJCZasEU7Fnj2ARELPbPFs
FeDxgOT1xF1RflCdZzfdVlxizuH979SmTvkFXTrvGF8ZkTQ2FTL8+KWFtqiPf80k
Zfhe8zLrTJhw2L75GGBAiIUWFROEtU8MEJB8Ri2X/PjVKsLnT4b4yW+AyfKGVaDq
yKPbpvahAwqJq/0ZK8SUJo39t/NordseJkxBSHft2V1mYaQZIoyRnxjSNa1nOdmj
jB2J+NSSALR+92JGx4/CgFWUoAbybwxx49r4rOQ13VQmkuwK2gPLIym1JBe+jp6X
ks0wzDGz5H8sL6rFp/t+3IDqMcJEfa/a6GZT65TLJf7orZ4s2Gy1Ansxxub3qYGv
x+vEXTaQjEUaDpZ0tdq/SpmjctP+2b9PkF/3Dm2U0JeFM+Kf6fh2mQh1BjPLrUfB
7qkj6UxtR4+esZw7ZmjBHrbFjYMRUZF2c/OIERWfIHHDRGv/0fZ00dTKqFiaQAV+
S19u+/meEB/wVutPjuTvM1/OURH8V3iHCOTTtD6VJuq3WbdpizjgSK4GhvufytO7
G+95qr/BFcKvLhNd66pfQckTsJRRvMalaGeilJD89VGH3XKpqFgQVEwWWPrp10xQ
+RwYijN+r8wKBNQJljb3W4uQ2muemX2YgE84xYOKxlVckZX23zJCTKckESmRx1Ft
XFQCAYKZI32FE8gq6tbA/IdOwqmse4a1nnLHlU+LSHsdQN9dapfPv1voyC80LFCN
AuNM4iZJbM+p3VAqPQNAiMS8eFM4eNqxixZVyxuTgxrfMNLWIdd/i1ov0llPTylx
93vahudIZ/oMmHV/zL1sM3OME6aYUYvM0c88ajRq6TPt08vHhdWRzq7xDCMt9uYF
4iWN52ffBy3IszSXyFqtZGCJAVf8PkcU+ZGtAbg3aerWh6ppUn6HksubmMcHLbC2
w3mtmTxtK8TbFTJvdvVu2tNp9ocKtlNU7vyOMR0B2Geta5LD+jdvInonOJ0NmII7
lkro4bi+pdPobQQGx2bnjjdR2dXMBcGVWBfxokJUd5vgpe8NOsUwcXfQDN9yh3LA
JNb1umFpTxKKr9gCvecSv5cYxQfHAWPElzYCKUForb1TFerdJtc3XGpyLJUxPpva
/m3stDmF16FZ2P0yD/bKCumVUx2vGsKoAO8pliEJdgguFg/5Cib9cMXO/xOwqriW
jOflEsZTxnHIBNrKPSHALiJHoMCVHpVr7VdHAyGCNWj9cXPjCHvIj2918FYXW8mb
n+9Ygli2HO3eUj8mihl16990jZ+VEapFlKnHeoinkhPFjRNv53vZeJdzEu3Ex7ut
/0M/SsD8THwLEM8w/dgZsIdgu5nQrlGqMSBEj9YDyn20f9HB+B+4jb3zMqDupoiC
85u05rEmPS+0bWxUdzhKTZ1hG5KEWX6xYfIhzd0QgM7U4BRBMRqU8yW5mOZTvvFU
YXHtgNjbs/vgdExZgovWuxjO08nDQX0ynZfbfj5zq6I4EDW1CHyBeRthB0bgaWCS
qRYg56xjhPDB8TbKzJYcWVFbG9KVVEHQP7KyQUnOFMd5yAIJo/8SXid6+CbBn6ei
PQVvYjzBDTSSZBmWMO6Eu44+pN7B91uaLuwC1G+g+d3cz92+h4p+kPHJaWirbvpI
Fp9N+M/66f6qTmr+cHKf1vTqfwDbBDiDQEpezm4ruYPadZqOTYrAwm9Sd29IxFta
pm4DAejkMshYHr5zLFRsT/uya3kVJPon53mHjRfvy09Rwv/zMIxLXV0P+7C8KaZR
2vBOvQw5rAJJpmhDSemPiDhtNzIzZiTQGFfA9BO1j8hPwmFs+V1mhNQbhuKEy0fO
Wr72bBOkV/oqGfNFghGmbMG9YABj+NcPczZN1YE5aZEeFvWK7AYZ4amNuU7/iOs2
PLO9F2mAp54JqRKImh1XM6/HknfQ03QieL4VetkHMFWs8pj2q40oZD7FxRW+Xfhs
O+O4p8sd0Rg+AonS0Qj7JFU1i4WwyofKo72LuFO6Foz8UzQnXmLIlFMubzG7Eb4I
/GnX+jQV6mrR160THM8g7nFKzcdFKwf7GWzdRZ+akSTnPDwP3L9M3IrgwB21xm2x
3oXwaJTMmaUL9olBS7o8JEmR/J8+F6AhhYaJJlN8KSPI6FUwweopC6q7zbPXxJHj
7TI5/wisgWYchEOKKAWHSQKM48/VNjumKM02TPXYP741Q8rcVPKr+mFXiH3E9sLJ
enLNlSVAsjFeWW6Vpnw5nwlZhsAS0le0YlX6CArKK5hTW+FItefa2crRhgJuD1bM
bsnY338+JhMjA2VxpGuFNAUHpqxOn5ZIIU/+U+oarLLxQidIMriQeHSgVgIyVagI
iWnB+u+fAt2UOsA9+SxX1j3ZnXeTb6o1EtH8lS/wd8Ef9TvkfMaWJ2S5JAHXqJqY
1/bg7QO+xt0DZCLfxP8vlEGloQLhs4FZiR85uC4m5hBReiwsgfnmQ6yyaGRvqB3g
bB58qhnUz5zL7C6KVUtoakJny8w/MyHLSO1CHWg7SBJosvvKmbF55y/E7QgWUAFZ
7pNKYn0x5cgO4uJPIU/quqyvFLqKewmn8xOFsWHpKzDxnJ8dBojdq6AlE66C10wy
tLUtDBBGPvvnGINLv4krtqKo7NKLRAq11eqTe3MsiQU8ko7kWJagB9WOc4/sgGUP
3f0BYZk1rZ+eqmWFtPX3ItRhKM9iD440+bC6k/NkoIBFbZ4GUUp02yNtxIgJz2cV
Y+twHyYyMsKcp2/wAEFJ26bGGOQw514CmNaFtYAIE6UABprIZmregOnQVQ8YR+Sf
CDPJKsFZ6odZqOvEOdaxGIA2WwQpDA1JMdV2t8oOhOpox9HEcKM3QHZc+lWSFc8O
hqUHK8tDs2u8E9MFaFKk08y2SaiXRBbH29eGMpIFkh9A2FS8xDcP4a3Is0MRvps3
hetJ5RVGX4l7d+GARGLlgQZFqqOSeOcbZQV3fuKiAoASNCgXxlHHnGXxRKvwByqC
LIlusPjkUQ2HrKd2UPfmfrADVW6FEXx8ArcbuvFkIjMEA3dDMJeZzmAiiV3tx7Yw
OJauVig+Sc3zXrHhyuw5pafYTG3UJrxjL9o+4pftQfjwxi5/3sxkASDHP7e9Qc4g
CHUw9/cTYNt62rV1Vaasl2kD6Ey97SY7WGNXl9eEjwgJy3DWG0RUVuGWPO0L5zVX
p8AB/GNi2fc9SJDbToWbe85ZQ8ufpTUhjrthcs/LyJtrpaZCw27ppBTKJS1kjhs2
20q1Gk+Y7jyntunWhj6a/VKs6KZmsCDjgogHhMRcqr+r33YuQ11uiMWT9cVjKFZJ
Ztc3ANDR7jJ5qxRQGRl5zKbWQQly0AhI7Z6WxP1revWO4CHLi5fyZ9FadGlfAB/l
h3hFUtJS0fCBGp+/I0bNS7jrFx8Xu4pwCcyE50+6A5YYBhEnmIBOWk8Par15oFio
8GTYXlKZ9+H/k/Rp6gvXrym96Z+t4OfFbNY1W9lGn8V0YVQjZpQxGSwuLZu/TO4K
AOViMNBVRB0qyP5a/Zo+ESPgluYKxDFQ9QBNgg8qPLGSMnspfjaWU1x0vEzzOfAq
b8OVxEo3ueFeTGXlYou3QoMeFCMhCVR6j8KTDNfy90uB0v0PRUzv961pkFzur8jz
f3zG4cn2V6mfExWnNFnNiPPBz+SvSMXoQeRV3nMD5SBcHLdw3KyEWCM769jAVmWg
pudrjJV9cWhP4uruL8Y8z6TGLTYYEH3wgXxG7DxoeoH8MZkjqu/Oz44RwBVugtwN
4CoBYZxU/aYKozooKJmhYw5sDcx8wgTa36vOMKmm56gXzAViwCIvft/VoNH3j/kQ
ulHXd6l6Cq1a1fkyPCArQt6GnRNoVoUQ+1WCFhbxVV0WO/l3vUvWAD1SWqGY3PUs
5tULwgqp3o+S5KeSqM2Ngk/jFNKAH9N9WnaKw4jEjSR4SgjymmlVmnO5MmR76buo
Eacq2xQFbp+H+PWt6ZDV9gFNKAmQKKHQcbYj+UjUBnT3cKqFFEfPyb0RfgEN/DF5
l4uBBOflhTjwVNJLhiP0ZZC/W6EmFkY2d3y7nK1rRHn3M3j0LD+ZeVsl5dCGZqXT
Ne4auRi6F80HLRRwZXiPDAoFDH+zr400ETbEEFyK8k3I1RWmfREgkJkyPQEbdZYC
q39EUMnoeU32fpBxt9IEO6e3Xf3HZ4gBiiWtfhIAuu2U864hpj/x/NeP8Xi0DRF1
2g1Ctybk5spfgOk8y47cOQlpEho0JIgBjGNROxtILcC1lmIc2efwRPP+CiBAYZU6
OyLjuXfIe5EuMFcR+nFmkxaOJ2Ypc5+p9LIhHZRQ+qX1hWMmVPKrnGcwfNs1NLOn
NyvC9CClv45l6MnlxcumvYA9DaYuu4fNFpCSW6dat/ve2DvqB4LYJrjBfMGtQt4I
qA0yXGfzWuhbAKhBZ29Vg6CIYxW7mW/HN0ZIPIHJOPNrzLyIsy+dBJy1tsnxr0dT
PErh4AHho30mGYch2vYs6RZBb8nUpB6VdfWpTeU41Jugo7HveVmoo4/LoDjoUnBV
mbRUgIhGf0wQDj4ziNjppcOKE0hzFj/BTf8VHhP7nyD2Id5pZAREfaZMIuDd6jP0
U5Y0a+1Z3kt1nptX5+7aZxTKX5xAoGGsl0vPmBjPIg2ZGCg9UBE5Es4dYd/7wjR0
RALAZw6EvKQdD7wtpb9IA00YBcScEQ2zjid6yAkuQAWSgz2kzZhEXOLTX3CdvkiM
PrDHUiBqPMqpsu5PcNftaNExe+XqRh4MwByGYD2S333439K/Ojixh40VfStysd4/
BqWB2+cFgdXDf3nq7z6MDSjv4X5GCtGrtVhwsZW/Wt9keqqMp2FtyCkgLMOsowXh
6AlHRf7EVgdqkWZYC/cmmtfM5xi5WKoiPfFjJJzlD06Cog6YkVXsGevG1UaQIeCn
uEd21Bk96ps6/QqMBm1lzscJ1Uk1SxFf6lrc+M9sP1coHJhN013jahLaKMTSVhAL
BROzXdi1RsQmh3ay7XRoM0WtpIpkEwzjIf2oXQFc3Pau8C/Dnzv3UVbUWZjkTctR
d/+1Fz+k7iP3P/iOKkAXvo/G7B+uVh1hELxj6KYaEuGfoHqK5HYMTEfzugzUcREg
jbB5bRtbGfJHoAUPcDWW/ZJQYH/U7BmK218zWwmfCRwIeOzGPqlA4cRRJjqupmRe
P6SvOGEAUyoP70gqzrumJXbf1HAeBeN3/Q+/4hVbCKcTjuBIOdj+99Az6H/p+7Bk
L5/INU9mUUcnikmn0pse34O+4oR33vODNf6Uw02Ongn0Ha48MWak6IMl510YIEl9
R9pCXT7aTCZLZlnyOUN/kpgUKpdf9gVmcv0ZG/dL3lqu228icy3LqroBVjemqwaO
6XUInq8ceesD8fz5Swh4KZNfX3GH6fcsejoan3oPF+KnLV4Yf5kUROrIPM26sDvR
DFi8XPnSqW+yEo3Rcz+4LUhpRM/jKWDexs5IWITPb6ZHXBn0kem2BzdXPJNjmk02
q3lcJ6NIN1xCa5Ku4qzUvjIFJUcQjrO2zFRXrHdY4BISAZoBpt+R4MPUXHjMxEzB
4D/z8dBl6jL+SS4p5LD8HrIxQRffbPQXqKI4Y4XMCUjQN9mq9iuELHYh/Lt8pvJw
RLW+J99L3xnWhlk9YwPSSV2R93xSPzTNoKCLXthIF2bAXGDwo1KBKFONtKSV7OTB
ak4DuMvBBYvwWeGlaqKdFXY6Re8rB0gauS/ddftM+Bpv3814VuwvHv/i8mcY/FWy
6Ka/CgOSND3W5XXRuIw2vO7TTY4a018vLoJWG56q2RhPprhz+QBmbQD1FgIcoYkl
icmA/DZz5e8dsyiq92EEUBRUhmkOy+teY/6PJ8QN/QGavvAHvXfp4VZ+27UpZ/G1
rMvy244FnLCIhKZNVn7+rwqiVdPRfLqMTQsIgQiA+MvpYnc3HXIOwCfRxyAl/RU/
LhWffPQE59hvSR3ymN+89221VcjGRmumsyO97Qjne5D7eMyTW6e5wRB+6+tqQYZf
1G3iO1IBEwcB4dJXLEIhDc7l6LUPz6XIPQk1/4TG6xxcWkEvf21dnmS+QdOBmVkP
COzO9jcguwfovKttDSiq6DHzK1wsibcVLAMRuMwRF28BfE5HrILIJso04Bm4wjBR
VOcwXluhQKVMyrr1OFxCA8Ux76EPV3/KX51MddrluE7APhvbUhtgNTAQUG43Qfrc
8MRBzTXmGBezTaoHYHjdMZFEu2giDVD8M4Yg8n0FbEVn7NiO/L0mry11Zgmj+Y/c
tgEpqUHggDlXXUnPcJeV1mV8o3S0dZXqzEuXyYwnLIjYMHy8JD41oi8OGzS23bAL
k1zphwQvjKTASX98dF5EdEMVl77t/ZnIXdJnNFPSZTxuv4AJ1ArnU5pM4M3Auz+n
eYNeTeQtD59AW/gbJnpwmz33hAG24zjbwiE/Oyh4cils4TD/ZgDoFGSTKRLZhO4j
/eFzKH6aOBeaczxSw3Kea5c2XK/vNvOzIjUkw+nuLWJhRLmfm5yj0ht5D0z2DkHz
zToFBDNBebMWmtAz1R+4ZOr5yPWInrUm3Dypz7s7dY60TpfMidISIv9h66wxlKaq
42y+/i7Wa4gdK0fXnY2viygmitAWUoVRzHnGJfgZ5tmobrTWFI5Z35j3MM7v6kHz
zfeRZwMgKijmv9EnqCnUi/wxLQIp+vBFKyqNdsNGTGjFBdG5pu7Wuvr1CpWKiDv9
26nZvUdYPXAeA3NqGL9G9GVps1P0tlzeEyaBqQJnT8vHybE6/ETiCKxDMFdZFj+L
5GYlGNByQqrDCDd56SPvduBjo9FSAVwNg2IAwXk0MycTs8K+KhOOg7ifGc7JXhy0
xvRHLUwiwWgztod3wxezC3ev8bSXrIJmaA+zY3sz7Kw5vp+aUFNIbX4uk3yhPD6i
YZONCwyJIHAPRY3ggASMeWTlBYGbVmVIzKeBbh2Vf3GcemAMHVWxlAZAb+5XMSnq
Yyvo6MvhzSzytPh0mOWZdvEU88rdNzHBn44PpvJ5rIyU7GyOQnPUn9yxzr1Nusgx
71cPsiFgthoVeYaYgtq34OezLGX9/xcjopIRrAYGGcn5BY2gqdkj/fFAAh6MvRX3
DrOismmoY/arYCumal6SYOU7bcT0+Bnw3+U+iMQgcbtZP4rnQTL47sK0glUIm4t1
eBA6mRlN9ZCrD1FSw6dcvVdNOKDjsbHDotHadcy9DZ4tv/6iWi3W2FoW5PjCa3af
tAEXCd2hKEHUZVXqj4yIDJZwFVs7vlrYun9M5JBkYpIrGMUIDD+DUo6PeVDlQsYD
zB9G5KUFYnhqayrGlsOHZvy8VkGoI4y2XMzpENIKeUC45mQFgSHqSTMsWm8kliNb
AEygGj7wjaKUK97RgZthGGH72NPSTXQnPUHvn64jqB4s9satrrc/s6wg/CKm0Fpk
76BzmIESN2OzxirgZmPMcfaS5oGfkeZOpPXq7dsHQgxkRwHRpcn3Kt4xUi8BeRoP
R0h2qOHhU4SjYg9THKCYtO1yOul9cYnEMWo5Z3nRdTf4tZDDOR54dIkRLONKrAB9
OQx4/dZ+cRkM/yoz6bFAsm1StnDYND3gUIoXp336GwWRNS2e7KEQWI7KsNtNvN0q
Pz61zc670g88i+HghSpaeVsjmnI8rbQxaE5wIkcB/yH3DBfVaaHUxTO+krY8RfA+
aQ3nQT5nuD3a+iDSr19bKxQCugy0dpXQGHqCaew078NVyQMPMsUffb2/8ezAbQmN
gkFNWELvXEupggDh74QRTpju3Rz8leAijg00raCW2oq54e/6X+I6swUluPLvh0tM
5cf8z8xvB/W/PqBpOXNPsQIxHN2YD/fRdmMGX7P83UKYq8St7N8H98BiO5UR4ghr
lOA1aBUWCEalz8n67C4UG26BpdTmqfZJbRGtPy1MbIjI0O7f642me9/XqILaTHBf
9NTTHIoz+zURfoGFnsskGT+FhnNqzy2AP7O2jxXnm/Frezw5aUlQ4oxRhFOXutnN
8TAaNmrrEascU1frPbYyGmLIo8rm7OzgWJ2BOPQchhS4nnHOWpfQmSc/ts53jawd
LbIrV9LmY2TUe2MO605ES8yRg3yaeV6Yw81Twvyh8tJ3/9FjfAhk4TnSitGT8XWN
9CAc1xWIQLBedqHJvIKHA8DXfXImxyY9QJO3CbnT2SvKIpitoKeX7q+ui1Ej0XJ6
i22dOgli1qv2YdQkpVT8GfAdrcE1DbgUk6tInZ8yjKVGi+4EjHwQPMqI6nhoV9Bt
CSfqgHVKV7XNRHSc2/YkeNlquud1QYwZo+1SqJCOnxZaEBUg117IwCNipP2Fd2UX
BmL6CaTGUjQ82esn1ieB5oVTdxgXPbbe/I87aAr1Voq/QXQ3XRiNe4bPdM1zq189
pxk1J/m4DDuEFc5m7+uABoXbcnFjyrxJ2TRv6uE9mEcMMT93XasRHn33Rp2Ly/QI
k6wOqnw9a6qNL+MllTcRJLaiZZJMZexmFB+rIXsztBjal+fPAtkoY8dgFTfaP3fo
YJagLjkcBlI428JySO0/ED9O484U6oTb50cGZ1ujFwziwwY8cC1NLFgyRbHF/hC7
ceCe8jgCIK2N05hPY1LtutqSc2PCwHgU5IvYzk3GVTrVt8h6f/sbogIDjG2Ik/FW
fgcAURLqaFCqKW/4nx4QwxdRVcrujmuzitU2cB86pmWKHJ0G8uguJ1k2xHLQeAmy
uHjerb4NWMke4CflKhyK0OyX45zHvQEb7jUjBurTLVSkQzlgJSCnHWenquqBRBUM
d/NSsvwzkttdFRqNOB/FfFwSoQ4CJ+EbTbUzIqgLNo8v/H/Ev/T2j/2f7XrDTgjJ
9w7fzhGkE1OnYi1ieYzbKjvmHiaSQi6exYgT4I+VhK5CzoQFpR7bV9E8wiQ8H+z+
9HwxtpAeWhdpVox09nl2YDsVm2v+/IJ7Q7Tw72S5HaB9hznVODqc0J78VhZDQF0E
scGHCoU2N7XkUxBwCO9UMLecc1O62ahGUJ3e3U2tr9VNJpnlkhSvy84CYleUI6Sc
+Yr1GU+4RSLNzxXLfec1zOtPICD4bArkM/vkj05eAKou2fjQVZwwrmjmGJy3KvdT
Y8F+Kk3GweCfhd6v1+me7n87wh9sVDU1J/1aIKAptxmsXAaLimy1hei7J9m3lX6l
084K9jOgHzsityJ8YRlzA8BIE2qHuE0jKXIq13GEBQbW6NsR8Y1uuNzVHN1zDTCl
q9u5DidEZv1aHUT+ndfFSy6bVDQtTkcnuEaMzV6BadACmlLEqRbxgc7dn4mInhuh
qMxs7/lQEZ7zZIwaM43QeyWXFUoRb8/39MALq5TIEWCZ/ajTmIxnSyFsWIUy6Yde
jhhbv5WDgn6YhGTzgu/AY2OkMs7XynWfs587hjKJWFThB7CntqRH5r3jn3mYyq30
VFe2N/DfwM7L4ivPueqK4sHqSA2lVnH9vOCQBB7d0dnRSgwuH1VOr5qUX16VkWyq
wmSuSU4ZQkHBNrjikBK+hR8ovoOHS3Pa4vgTC9d8YDAlUNqsFsqWVwVnkzArrwf1
uW+Z6zCC29hMWrrEMNrXd9yjysNkcfwwj3VvIcbMKn978r05Z3tdWIIGQDAVZ0Hk
DGs64Q0BMAr/rlDbBpSQuvvH8Y4JmbP9xvB+nBm7ItD8sQLLqtde6BbRm2NdARIy
Chy0FzxVBiBslfQ+xtQHk2YnqUzglBIlxHxfjgn5Z+ONaLqz930VtnLvLPdX/aRl
sX0VlgR++7rpBCOqfDklpGQIIhueNt0iZ2cokOBXj5aLYGvf+gAATYUYmh6NIDoQ
fnz88N1B72YdeyxQJKez+mxf4/MBCzi0KSkmQBYRpCatYzKvev8VZncWx1yo4PrU
LZPk0aYSXBNZKII4RF7UWJ1TmmTyRx5jPf4WsyI2083hiqKgUrMQO3MOyRJn5CGC
X83d+jCKlZHDBiZC2kCoCDceiczrpfho5MboNKhg3xz76AJAX3YKlrA1VYvBTV1T
sSlGrjRgnmxET8C1etxKp8vYMMMO5HOG22JJQTj4/1RmvCfGq5E3pJKjQ0R5GsRr
TpFw071gbb3NdJJqJAug5gqX7vmxSvafx87s349ksW+lGZAWqXR9B4+vIZ/XmQaU
fDJP+rbKFmP1qWiV1Ch4ENFZ8rGCx10HVUQgtoU+LetQqEIOPuuQOR4nFG9qNgT4
U7gMtVs3yGmE/Kf9zEn60JC6leFDyUlIIiHsAuT3x7BTmwA3brdPl9YUsQxv3BPY
sfWxR2QHWXG73n85hs3nUISuK1mNnTIbpLhqSDZIX7s282FaYnx5usulhs86tbu3
VBVXNbKN6aFPrle6pFVedyGI2hBU347m/y+aTfJMCYwePpwoV362sENUJGrUI+I+
aGYKOcAE2Ckk4IYfPN2zb5HWoXfdlrJgxgOr79/aM3hplq471T8ouTpwM+M2p4Qe
aj/N1f7y+oVBMx3iSwNC2aI/zbT9zguEP7J06xxTGNSv8+DdTm3Z1c8bPJ9YwaqT
Fa+WgEM1NedhdKEzWLtfrW/rND/2euBqmLWoNCC5kq/kscbk4aAllIJDYvaLQpwz
QU5unrQ81C6au9M/10Bii+h3MojkLul8oF0SpdG3tDaUAljaBKqGu6Ao5JRZlFuP
6Qm7FcJ5zmHcvEPy92ZU7tcNm9MhyPH6sPhL0n86XZDyQDzoMdOJAVMSdk7NySDT
IGlnF6YwiBxxxMB/0Q8AJn2qR/0lmxD7beM31RZBws3ufwaz3z7aXeO2RIVp23jY
r+5tcFY8CWlawG30j+M2s89eCgmhtmtA+oT6uLELaEJcJ8j35hc9u9CaXf8OYA3Q
j6I1OQ1jsq/gGqd9Cl4mzjKOHNjM7cvcXcpYjLAhJ2LKB8SY7Se95k642iy6lKg6
B5ectBwazuDRffiANX078zizT1hFbQtJcsFkFPkK09bHVo43lzS9wPx1YnN/c19n
tE9zaouMkKvQCk/GEnmBoRkNn9xuCRO4hBKcZVCRKiAWIlenAci9hhUhDAph0YTi
LiqP/oV1OTvlXdGRobN1zpFLXDbtRf/32h8Oh0EltnyNqYNmcsHZOvkSvYri04FN
GLEBDHrMhI8fHaziituBlu2TCH0//k0WSV3l/s9toXjreTHun8w36jvizp9Eg/QM
Ns9O5ZdQR0x6M7X15KUlNe1C2B8ZxFakqziarTkLQ1CIB4TxDfQQbTNhMXfWfruJ
66/chosK6WasT76sYAuRqnxXPSn1kx3+1+96mVkMczwMLG8ExeTGFULPXd4nLsPN
E8KGq/H5SsdJQRSZYrUdkVNYoYjUOlKhk9LwFG4jIjwTW7weXrifY86GusF5eZgB
vY0xpg5QRluP44u9XeiUG1IsQAVhLwBH48zLtW5ggbXpS09f6FK+EI9C9oDo0Pyh
2xXhTqDtqlL+LN6F58kYMz3m8IS08M94ZvdOTB1VAa/2TCHAaZkYR91dK3FWKYHK
v0A9QfNOis4sY9d8pI1wxiCZJaBQ9EYvYDRZEpEp/fSfAr9vjTSwER4L8upPdjST
71cZEz/WDFCZ4hiHblMEh22xQcC9J09wBfVQyfA0HteGesEXK/OE5a+N03aBE/Nk
m3LmxTIpFjt0sCORL4NlGKWRgIsgbJ/a0Fgw8WwIJEPQJ9hjAMX3OAIeBIG9zKhW
ysTUo2SZ07Re/ahcujBUrM99Nvg6jL5E5wff2MF6rm1SZukeRsWHtsW18Mlsk/2Y
oe/ayvK92IZAEezE6iJStlBN+mhVXng/lSkXTAWSfKc8f/eXs8zbICh7gNfNaKI2
MNB9WLmVvP1vCdzBSCz2W/i3bjyZTzEUU1Ypglb+NyXrMCbSXozh7HgImFyr5FPN
j4VkfTmL0pKhgse0QCdPobQ1iyCX20N0HfeCgjbR0DZHdYpF/zcsLdqP4hvOSMzg
btI2L5y4PJWJqPnDZC2eMIebULVFYurEpKxY/raQeVvys1P7EeO+JfRbmNkEU3oA
xdfcGaFUbZF050PeQRgLRM/QQeob9jOtJoloL1CkSUOUxVzTMVTzYvewn2TlMoy+
X3OCCsBqhMp4KIZJrGsUxUR1dIJxow7Jb6iXTbVznqKASRqhQk/hZReZsotgSW3H
su3rZPu6EHxDD1lQhaMBh09ukwv4eNwT4GxtjkZPQvRWLCrD8pSWKySZlRgOMzIA
3WUKB6Z2uy5kv1WIfzzrwP3LVtecFCI9IYVB2bDHqAFKLK2xmg3dneVwrzWkuefp
8ULzYCzg8UCBPvsVa5mzb1MCcKd7h0yScAw0rir1f6Z8Qlu+fU3B6v+/9hBMGjsw
k23HXzJejSFvyS3GbOFkcX14obX+8V8RKAErUZ4r3a3klmQVz1enbZ9jhatD6CtA
epARdhYDUoriF1NJlmqnXvVtSx/ajuE2028KITSSyGK0CYTOjTokGq06NPEc3U8R
IhKhoGaAwGlQArykm/UideEPqjwWi/Wntc/aGErDopYxetQmRKBpyuFXGtWpj4Vw
VoeVPI8J+YChJl2iAwf1cN1nmt6kqP3Ay09q/obFRL8m+NnAhLudHDuegwc32MyO
ARsxliXyd+QrWEk3wUUkoOBoEFeFPVTPO75E6YnJF9VdLfxE541mtc+IRPHHV/rB
e2f2DgOEtj0rEVn7Xga0IubzDQAQqtf1lMu5OSnVwkkxdfpVwL4uf5oKnVxoqfCI
Fa7rH9Dd1CT/c6XFbIwTkarjlOws0D5/m+bib2iresYrAuQX+MjRT+fCGKHqEK9e
kFlISrGKPRviSTJo7W7QjWAFvV4aZ/Ae2MakRlaZf90aO98t+PFjHZwIGFLxxxoy
5tAfP3sUATuwh/oRs6971rgoDH5qO2pPcTsk3w+b9+sHm/C9SDjn1ItV68dglb8L
gQhfDZ8pi1AddWUlRITGgNP7vYTNiSYdSLK8kyQZpEewjhTqOK8k8amBKX5+yy6I
0N8emyiCjUQM7tocnnyCOfpgsnGY6GNWiaPK3jWBAg8BJcee7AQSeIQQ4L8EIF/H
IvAw0IuGFiuefOxs0oJZI/N9vX4irHT4zk0P3kWnjwIumdJj2xQvrOVJpJxO9czU
8mjaxESpFrGuqANjgPNthIxR3HqxdsuOfXyPaZWj1fGojM47YYBPlm64pSMoBmwp
aLLGDFTgN2shzoLMI5KBgZMfqw4a3H4gr40EiCyRn8LiCr+y1KHbMLt9PKtkNHNE
6XkZLVLgSjLmKpKlAMcWQL74vkbIbEcnW7gWK/wdsP3B+OA3GK0O61556fc0ALlB
IfRgz394KqP4V4MVHtBNkzDHS0hrZbKqUOD5Cfc+22uXSyKeafXxngS+hVp+1n1J
k4tBNLojU4zmCW6fyOz32VWpvQWUz6wgHuak28muk95uTY+ffD+Sp1Ubgi8nVKmf
0Rt8hT3LWZkJvtPLpkUBW/2KJMKc3IQa91GMwMc2a7OUbGYzWAkD6X5CKOKJjnth
K/MXU74eCVq1kBfIApSp6MB6EDRqLoTUvC4lxDk+ZWPvt8xcF35+sE2/j1ianh3c
s4X25PrekTugck4e5Gf449QJsTu+n23caMA12CxTy7cpwy3cCnQMVs9mSWHlOFBT
Al++ze7e4FJe31fPSyEVXjhhkSVkQ//NELpuZuG/82OT6YqUrQHXLeA2xejP8kXU
xkrveLQVViRBNM9Q+PGk0eQ8aU85JTABTnwjfwFEkya+f92g5wTWW4Uforps72yS
St3VL6A4AELEZ2tgKn6HfBO8esB2qUcwNXbzvvXw2PYGZReNALqB0JRiNmD38fGd
SIzQKtgUU6RV/NBORoxh5OQnvJk8/FqOh2n/C4werH1okU0/7zU4KUGGsnjD6JxA
xdaYjp272jj+fzk6nHrovcH9t1QkwEe5uzLa+eIdPxbU5qAAV/dHJaCl/apsUvTO
I8O6mpmKqm3QCUQvlNoSEOjZVsexsukANPfhkDptw2zEmKURlhzxcKJmiJf9Zq2w
JSc95+QwC0/1+pVU/WqMcJJfmVaaJ6Ynul9umEO9h2UZqqnklBTUAwodEtafplmh
mYeRafU9k5U0L6LpMP7UlJ+AD884yE0jvGGcqZ1oizruaeBDoKIJOqrSrZ+XxcZZ
/oecLeG/TsHSLsMu8/IZlczTSIYcVqgeDJENHQKuk/lFeDTq9/teABAc6418ANVF
4p8afx2+9GU0i4RdqikKQtZDb9rOqmOnncibBPEr6CHlICNqwMANyluDIYDYjdXw
/mhmDmc6LtIm6mHm+zXllXlXTfdqdI5nB/uKnoNRp6BpRl9r//n3vzevJMAX8E99
pqmke08wXDIIDKjgGXTQVNydjEov3yJwJvrTIofFV62K7M7+2dMQe3x0y9oXkx40
caR9GNKmImznaW3X9kUs+ZtL+4lDA6Z/p08VCZ984RJec6unC20BkSpMKmnZqGsB
Lbl9MaqGMGHSoVtfm99kgDCE52GykmyafAK7pzanXpHLLF0ZbI12091xTp6YjJLw
lIos/tTafMuZ1a3vgu2ifDb0ORouIYptWV/pYheLBne1bSdJXq4gL2gjX8aUTO0/
PB15AOKHa4NrqBbeJvThBN7UlJs3+4bEoyvpPFXZf5wo43XJv3WM8Xq2i8MrMXYN
RZxCDtxqjyEFqCvYIH8z7aqFnuR3XdYX/9ldGfVq7L8bkO+gdwDed9A+9xvY7aNu
1MmISXl66/F2v+93gTcND7YaX8jhCG+bwhSNlkHdTawNA0V+C1g6uDB6Ot6Ap5M4
6SHC1oR+m+xC+5f/RBOpbwEp1tSsN7XJ3DyvMUVfqm23aeI/+WZQ1sGTe7vM+RPo
9Rtl1w1XaVg9i425XmGs2xPNtYB8gtSukgObNRrrjLVABZzc1p/GL+QHhEV3shnY
UnMakiZERFmak75z47otBGJRrtf7VIR38eYkzJJUHYsDd/1xarr9f4dpc/IBMdjt
OPS2UJ+rX8iEEEpF+98f7wNTPk3kY2VmSok5h3sctsFDHFKih7GhA509f3Bx9EBa
fyQnJ1mriv6rCWa6BiZ8b0MuwTmCxFSpQbggJVAedtQAkPXvi4GTcGIKl6sTT27o
iuZ3akcYQcN5vmuQYyFPWSyCY8e+/4btHgb1g4YGa5IG6BbAR82qU4BL+ge1YgZ8
VUrNH4uRPscXXSB0PlgJ9gRBBjJRuRfJj//lhoxcCVPawiU3CwQpAoMM2z9EN8Kp
DLl9zHpp5ZiPW9cmnIp0s28FrQqMwCShWYn0bjPrUp9gYzRXNHr/Kvsyrk7TcEpn
pE2UKUVBG1atSEA/SXPR0qydtNmh5svd2Zs1J/oTmHeR6lPyEo8d5qnARMmpIPwx
jy2ZYsPaYyG6RwvbOaBsHIQ7wMHYHQ3oYY7Q8Uv5auBEV9g31WRAFWk4+PN/LDP7
H1U7q8Ydc3s4r7IM0Xb129RVj3ZDy45gfh/lExO8oVKxRrRBzdtN8+wlTgj2SEgy
OomD4/vkLr7k6F6fyveFXXbfKJV2af+C1bjuNEldt+yU4XhhlX7mFa5Ve1Qd/x4w
WgUn7a70NMfC+DjJk1eT/0BPuDDt/MZ4fOb4DoRmlxCd8ynxOXnL2EQ4jVYgDvDJ
YQvKhVBTGSqAlxp8HF6i4Nl6GKi1gKnAdvBqPnz8BPvAYiZIiZeCOVfaN+TGN5PJ
kiC1kImHNt06B0/Gbkk4+IiDkcadlRwNjGrZw0CtV4ejlVeoNKYXv20qxmXO7yxZ
6T68GLc+C3EBcz+/3Tr6NBrEjrjmKxBS1FYykYlgrRgJ3+6xhMQMyGYGOTpfMAnG
xSrJU5O5FKJOTMsyXR5BG8isWqNcshXV1e58Wjwlw9YyU5Myv0f/OyJ2QkKos/G0
i2tzvxVwgr7WQ35p0bgBp//NvzjHi2NFixs2ZT+jEI4qrlnZIvQCkfYEM9j0t27s
HxXEmybKYUPVz7vGx0EmtGD33AXv29KYZzLC6z92XlxQcM22OKbtILg79yt/m0nf
YB0245rj1gUZlUJo1McMPNMNQolPmeBTUSDgTdo4g+0a1JZ92yczmXJZkRWSQErQ
EOzeJrrsnUeinu5MfvnGABfiFnE590PM4EVkI+PKX50M8wRvCmgAaYckFaGf7TKO
1MEb6sD6U2ZaUYY01qlB1dwV7ng2kyqn8GQt6jZVci44jjIkGSI1Zh2UCe7lJopH
GQQETSmMFkObI1v7ix5CzAZK2BAIR38UbPvdrMft2UgKprmiaOyhL/jOv+yPqrCX
fFAw1F/k31vVMdPfWPqQZXYuKdDDNeyyBQ47RWLMJlxZQbjcXR2vp+amQjdWl5Wy
ng2corx9Kl7RgOq0wgJuV58/61HnEAIeIuZ289xbcJu2Oi71YkVoQBwLZD4bYVce
lb0uvZTQxmrkV58qIFyjbcsmRz/hSwtDklKl1pRHBVTmWm2cArbOoi29+5/g1KsE
LWz7RIuTFg+mlNngPCwxdrPWQXbM37TU9SpqFAnHCqsedu4VFE2vvzRwB3Llsz/Q
4i5p6pEHwQNWCVr88PkOmzLBqcQ6je2LO1w3NDzgp6+u53Sg/LKnNlJ8j3ex2y52
/4b3MkcvXRryS708l/CZcesBJqUahrwWi8mQZKVEV4DIKLgSNwiHCBRKHg3wKfY3
JEGXMpqTIYrITDzwjJB+oVg3derN1d78KDUfdf8rTfUQZugGUHPgjaugMQCgYU34
QkCsphFrUWQg7AA+KVovwhChdp6EpVFneJ2I+rGWGGrGiQyqqYNGSA+1eJAaqX71
0ewbMOFMe0DLc2P3fpTf2U4cZxZnimGliIyRtIkQVaPRganNukhbatt6JxKYbPJ/
4LsWueuww70b3+wsq5VhS7aDKuz92yI4yfU+U535w2FbMicHHtykdIJjex0o/cG9
MTIJceWNJ7MtCy7cHoVj/kbrTz293VWZ29z59GfWXBA4BJ5nQxmc32X3NODNeYX7
vzppIteSYNMyNDSr3b0ZiwTGLFvecn+OsH+o/lohniov7ukOt8dxFdexBxF04QHI
svY3WQRNWfV6JoDFq0LTFJsUNuSPFJUwMgnX/2UaFI56ZHJBQpKs76auaCbgeiaM
U23Eb2bFHB+suPMnkDaZKxvNDszXUu8lRY1AUYwQeUzskIJAtYdibwkZcUkXrAEZ
ZBZBEGPo/qpTTyZvXaaQY19AzTeGbel9be/c+IMykspi+tXHawSFdvjvYzuUfFK7
NJfnWkTtFQTWUEVr1B5S605gnajlftjbu8yFx4rG+tfwhvPexJ7+zI5cL9o9+US/
/kwje2Yot7NxpcrTm14KZeScwXA3EF9louY2CK6wgEhrSWZ0po8U6aYyh964TGxq
JNVYrZxHYsC/nNno9jh7ppfWkgMFK2GW6v9sYooFE6uZyTitA85xrZ7kD1yTxOIt
EoUKiYmyFL0FJMGoMzR4aLte1Ct6/8g/JScJXzHq1SsmMO6FWFjh4r3p5/J54BfP
Gi4fOhmc5bUkoVdef8CoAOFC8EmT0ccmJRX0+eCyeNsYBSBYXsK8d7onfE6nOb/u
gkEeT9AgkiO/qTUNuhz1NdDeQYPdwsoD0fXxGgXUobxzpCKz22yImFBOaSjaddrw
p4Van/mWzTOv+kh7DGOg4z1ggZyXrTUu2HLFM3gDcoCjxV8jGAEEEiDu80LQ12Nt
66YZ4x7KveQT4iqKD7lZ6UaabXalws2JK+x7+GWurSHuwWKUGndDNVT84QHs4/YC
cZf/AOrxpGQgweInToYiBu162q7grvu6rvepmZjvCy9IPb7/Vg38NQKOK7h1F/GT
u1NmdtSqLQ0zfpr6qrFeQ6vgzJhpj9WTkC6pcmSBct4302H2hXQ8rxTZhTK0aaP2
N8zOye4FoWUopJNqUJ8Fwoyq11Rf52TCatU/vMFCER9EbZa1S1Voi2+d7I7BuVWe
OSVrpqe8LhERsGZ5TTmfsP9E5ueMIgKxJzUQs803Gm83i1E6Fm01bOOxlvYiDgxP
dua7paOBdD1+fEdKPOr/o4qVZuQvE+IvtxAFv/dW/zG7+Ss/iHBeYRllRju8fdPA
TK7m/pJJSKew7MIbdtSU8kfNXu/5tM3Tbdf6azYxWi1mcG1/mR8J7Ro2MtkHvmLi
2LB696l45LC1Lr9szw4YuCxWHmP4/OeXhUwTeikP66eRWAACgdOohwWZXmgpU57M
DAZEyTNeChbFbCFBkrwethPMRLE4yeMoTFIRYIqnQcQFBJIiqY9Uvp7XTroMwDBj
D8elihJiek9FXSbuiffPGt7YlPj8nAiqBPpbfpnKs6KAPJ+IdJDGQwfvSBuBQfxE
UbxNBPLLHWcVadHXYTvqV0LfW/ve2Q6B5YOHnN2bN/8Pwp2wvliKAaXwt1xqUBuY
nNXReOjQXycHM7jvOkUbgpvJn2r3r3qA1jGnBKmRTTQqR1VDq63cddW66vAIcTmc
Yu1Egve1wAi/stzSQCtxJ50wptQRvSfV9KZR5/7SkF8LOmaXNdIFIr+XVJz4CfM5
Aa2yIiPjmrxe1xLohfgjnno1X70xJPWerq3olS6+rTzkdyGtafhLR4Ybdd3I18in
N0Zg4FLnQdNRCq+aQMIHWDJeCu2smeUIwwL5VwPlzgOiNQQx/ZjbPMGiYzyctvZ1
ZKjuo8UoRuPjgkhNFVA0JcNjui6mKHQYUZwz1roEOJ4ec013etrJyJpLb5q6lLTL
Me4lFTWECwp/ma/Ywg8hE8+5u2eKpkn0wQX5F2fjCNUJ7HwdHxOrLO7FcnDjkaHF
NB9QjHLmKO6u8PuyV5SNl3UfRJh2iSmyKxsjkuX0vqGNGlv2fwpWRUzzp81HfoFi
DFufa1SziR61ePVKA3t9SxSNQdNoI8Ci5JrUj8QEPKsq416ZKVOi2qGtKmTUASYT
PUbTWie24QEO4dBxH9jfphXjg7Q/E9LPMCeCEDujnWdiUs+pQx1dnOAVAnlXH/s/
5GjiJHrAdi9kFpMFx0A07T8PlJ+8vXGOX+Fe+S+FeOmzME63+ulqjKHFS7fVEZyS
gHc0cv8WZuektkD49a31LUPNHlrOufUYWlfafv2j97d9NOL8RrdIADgNSRZT+DsX
0ZOSBnWa1jjBFEy1LkGlYzdXZDWDha9i2CBxjdq/GH87IoPwTup9RIbh7pf423SB
h4a2Y+kopyKcpiUj2VOaLdKlgVorY+HmdE4qNlF02a7VVuvB/Zv1BJfj1tayEbHV
3+AEhIywSCHiJqs7NVUuACZbEmJT66qSz1mMQkyf2TQeGHecLH0vN+8z7696txVb
DlFbgvsWruIefDMQRLGmNhRekKswFJlbkteVw0ab/PtkhOB4hFkDQHBwj0yb6Yes
Setzr/lz9DfPKR2L1akLDfzq9cYqoZJZxFhflcBaqxryeR3eIRGRw1WK/rCy8A8d
3lP76Ek5+ShSluy5BGk1KQhy0thZSmsVmIwOXObv/p+wCZLMJk2d4d3z7tyIveEk
KQU1O8JL8CDLlqUOBaLLZs2TKYE0skcyOOiYpsGSiLwuW7wBwLNE+dR7oQoCoUq6
+oEgvnfVTdcSnACv6oyxR/HkuqvVJFIRKNNvgKkxWOtUc0ZHLEwisPwlkp1RMd1t
CAYLDbnClSGoDyESwZvvKJA+dbbzfVEUpOAtNJZ1//X3Xt8TmenLr26+qrOXlzPJ
SnIHVXo+h9SdLqXn60ELXtwUuYXnEfzLORbluk25Fk1NfwdzF+ZwQWyZT6dwh1AX
TGOaQZ3FatF6zfMo58jvqQPDkckzx81AMDqDYfGO1gP02mhVy6iYjH9cSEHOlcW/
t8nMmeH+wPrOJy/YZXH7IPGXDu91vaw0dlAftxOOA5yyHlqjtcKjeZIrdSEu6xqW
MKzAb+YBSQqfBmP1jc2yywox/FawbMtC7TRd+8TlZs2e/YPzPQO/txm4Ayx1ppYV
8DkHbCblmBK1nADXlsn1hrvhrnGXgGwqtUsw08bmx3Uj+ibcrfYfVJTPemcYeyyL
btzujGnh/ioRAKTTNCYlaEEFNRHcx2C/O4gCwVDZ87dk+7hyPULeX/8HvSHLhN2f
R226+8WSa16YTBzpqH0WL6sYjv3QKNR6ucBnI40prvLHD8Rxt5SN7w23C2SOINfm
DleFin7RBnYOTGi/he7AUMq+hJO0t3d8HED0gOJadPec4/CPRWdtPCfHc483byCG
roQdbSchwQoeQRI7tKPWOObjbiJAJuhJLl8cN6z1MIRaQvLoa9D4HqaOL/4Dfast
gphcYwYFnGCuZDOxXUXd40b8HYjWE7CQ4KX1uQsqhJuK5SB+S95SqObD1kRvaLJY
/DNQTEIIGd3boq83uzd+3bUBTcBVm0vMhvF32RTo6T9OVMiQ+9Koya6qm9QLcmVE
cPKFSQtdR4nqLhFCLVczFPEe/XCfmBndLFoIoP8/o9jFdxkLgz0lQnfc7ZrMZjQ7
AF7XpfAn2uG4+AGYGojdQHkbEgZ0IwqI8rST4TKRDcfBtqi1qyCo4jz00wGzLuk/
XU7bQhxkKUznIDhAZwFSS0wcmRuj3SJUXGzITCgza8qGgOSXBEi12zXs57Rm2Lh/
6jJ5z+9nopMLP9lnlqraE6I0pSDzzdDXWVldwcpuk76BZPZSXBh/8ZBJTIrU0Wyf
48xXZbSioIdrjW0RTE8MXUsU1eLuicACQtjjKXRay5dLuuFUp9IQMnuzfpIk6HD/
GOpSdssNoziN8lEj7eRpE5G3aiXZxl/qstDCyE7U3kTwvfN4HGyj6M+Wol4AV/KV
EnxVDcf4gjUiudwdmFAaRbp97l/kJC5Y9CGznPT34c9RF4yXIb9cElgoiPFlrleW
6H2dAWbANPmMUI5kCv6ghgemceweqLa1z0/bk3xhfED+IscOcy4kBf5B8TvwSaim
xq6TDhM0XE68ga9iQFURKljTf73+xRtA81YhSxlusFQTDsXqkaPk1Prv2Ys19pFt
6XVWODuExpavobSMmCQgj19W0N2vbwODzrL+4Aw0UGEZP5W7uf8prrF1sbdMjsB2
x7enuqMK38+MW5yvcwY3VESd8B6oKCAQCl0IU3yuUutRQVjTwm0aFaZa4axkZpg0
QVuKwDuEaCz6LBlK/LI6YIA4rI9Mg/An2HNFG4/GRA9x7tywCQe+mKooTRPkHK+B
hIlnqxDQ9U90SgVq1fVCjdjUvKC9aReBzSRkVKjPeckUFLfhOUhldz3Xkq7bWVaI
KuGmCX/6AG2JwIxwNneDCfrVzolzaHxhJsm/pogTt7NpSvarzJQFqaThS4G37J71
2hW39BUzuQtaR+j8dPVXgLIqmwE2FumEjtQU+oVruewVRRw8p9bWouQOTfqU8zkB
WsvXcvFPDLNP+vh0nSKmIcDCPDDROMXOI1cHpq2hMme8473yLNSdWLttiu/kDTFg
Ge5JettL0pGXOjIuuy4sCrUEPHmpLi1l2l7d2huq4w4O7yXcyuGmxOD43GNBPG6S
Ro3xfRNZ/HxlG5bbyCrbfvpEWT/PXESXpzCY8LJDnVkGvwdnOk9XE2rtnbTcZrt0
FDmqWYssrd8HdBsxQups0uIFCs/zrFM45swTQBobA1X9dksqYpnjCUaugYOx+9W1
uDIDShT1OcTb0nGO+H609/mxzdBiE+XajSXIeRULiH2UMz1Dh7wlk5Kovzl6z97S
qBecjsCjcOZscGoPDDnZPc1d67kTS+0j4uH9qN1O0THKTdVJjZWdxeclGUiqXT7g
vD3IY6RgF5GKJ4Gt4F5hxV5lNetxqhiJ07VdbslHW55xITXU/z04as2FKbDaorc9
qxO6Y8P2fK75MLoRmkgK6bL0bzoEc1V/3Vf7Cc2eJvXYttIPC7nuL6qgSkZ0dJeC
po1qLBCTPj2Fs00ABC6Qm1ic9MceD3Kwe+cEv7z5rVSrIjWc/S3UbceaYnPxZp6x
VijBSmw8Fn0T/+sosjnu6zaXCVdqdZoQSM0dI2ciwpB4Ahho+wKVanfm5t+7TiYB
1wJESXy8+OHVv5pz7L1Z85NXQOz9ybck81rDR72SUE40xUPmgItZxXn5Y0dhevJd
x54Eb0pJNEzsr+YDiZ1fWRvgp1co9kUfvuTsWEFi+g1daAdx1w1zf3b/kRp2bEHn
6uBAK2YZDMW/PLKR9sZk+kXg3wtHsn2Kt1qERCBdMlodXfLW4Ik5crNs1Nwh+lhm
IcAjycaTe5CSVcfzFy/Gi5Ib1aEGGy95Bgq4pAMR6BcvnoAZ62yxMiIRIM5hNjHP
SVld9yyjv7Ec3qJy7sP8nBRKqlSW9iWDU2rfcFwpT43D6T25wJXX5Klxg4M6PQ+L
XgiggvgkGOmLlZv+l1LUrMSLh291FRTCZza/U0NBiQPL1/kpSFWLBIGeZSrEr7CZ
u8pRkBrBtodASHPj9owGgCYWn0f71zY4Hw+q0PcJJWpN+UNEzhABbuBsjh0e/maE
5qr4J9dpz19bQ04tcUDIzBi+YT+Hxp4qDPKN3VyGhbJCDkgeAfYIlkFiwRM2JGhW
S1apFj2xlZrVM8pMzdNjdsEebjYJGi3c7Xyybu1ZlCGYReT42c/qtWRAo3xv3Gom
ASsRfbATPc/rate7ruJ34OIT4TZpsfW6EOPhILz0/1dDNqTyKP/Zv4w6Ia6UAU6Z
/5QdzhMS0GnKwGxqmNvkUlTetaKiDx9RMVPG1nNw9k9HZO64awxKSOTKlLL/ugfI
0mAS6s5VPx3PhkEV6KWorimYZXmPEzOXbaQEiXvFr4acsgs8mEi1eMFwEwt8oNoi
qZHGLKXB3/FCldEWnK8MaopfJ80VWqrTLTRIjHANQhDGZ/cUShi+t5v3SVfpkmNs
IcS8CFOtCnx6ioqBkUqErhQdYUXedZK3+aD8qeu70K9uMS4y8xHSb7T6r9ytcjLr
3AujJr4LFM2njQXvOCq4VC19Wkz7AxLG6kaKpAaj6OY5kPOdRdTdbOF3eFjYnk28
y9PzPdV6cpJ7gylSoUncfso7bEY4pmRFKoaYiRzi9lCg2hYSx2lrmTK3lga5iSaI
lmN9BCh3bBGQJXKJLpC0spcEvRggeauJ0N0dG9NnAc33AQY2M+GOO6bSzxIwo3hx
BikNqEDh8xGjokR2+KaDIF1ucMY9KDUrfh38PiDUfv0St1dkN+i80LFzY9JqNVaJ
tifxedl25QnIVJNw/l9TY5xyJdBCGZGO68+G0QkbIocX3PfSbR+0BYtNCRwE3BjB
4/c2C8DkBxfp/5Ybvkxxz790KGE37hH+7FMIniZpELmodUbdFD7OsQLd9AC12JAZ
5qIruJqb2K10VCsfANwK5gowNOJq9eKLe3P90OaXyADVZCVf+3a01V5C+bEMDewJ
iibmXMyKuN/Sh0nP6OM8pddcUZcoVzcDA6Y+UhxQN7u11GoOorINjpeobu4IeSj+
ODIuSBfPnTWQ9H/l1IG7eWKya1Eyae6J/7Jbdyd0zYECfz6Cm8bzhKpmv/zKEwZ/
0R3FAtXHZJjNUe70fbAE53F2LXo5z5KA7R/eMK3hAZtw3wuhksLBIBwjJTD4vVqJ
TZ7onF2xgIfXtjJTM7moXxX8rbKe0QVqbX9/fOufHQ0+ycE4BZQBEH4vtGm755cH
Y4KSeSXdLopAcQCCT8u6qTKOG9UygAl+iR9+ZHo4PyGgq7hLC8wDMOZ6C3QTVFYe
Ee8H3hZo5D7SZyVVc/lbnhMXQoPSH8p1ARJmjzOHCAqqKNVkTNiWm41oJ81jTJUM
whL3tqqGaZ1JBHGSS1xN5r5LaWLNvossuJIouL30CR07Gh3sTWs7sDNceGFgVrbE
aNm0q5VCyDFga4kqxoOvvJMuAx7PvCqcRyiEppMJjEqyS8jh+hBKtR7JLeXVm0qE
W5U9awgaX5HwqIYbBMfQj+bKO5faDIVX5SB/xzZT4qR0QBxS9UoUiqdOiPtAL3cS
CJBmTDpy2EEv7naXOcxlYFqmN+9l+q1G0/73GBkp0UityrJgXzBSz22b3/aRjj0s
Edi2wDtG8DvAu53HzpVasnhqMR2DaT9jLfskjVlMXBVGZ/j+nQmmsH2XEoi4G1tP
3LGfo5UngieDBUJKmBa8eAsN1uV28DfJdv10Rc+GJS9ogodsHeCPQsUP6FIPaBBv
Nhbe/3d13VaD9/TNw9cL3+2byff2I2sPOehAF2MswDyrljhnf0uOU3wTr06mMdHs
vZuRj+LHflTa6LOrs/F1Lxz+ON/1mmfzMoaBvwknL+qQS919u8AeExprEamoSWay
b//tPn9lznXxBM7T09PLupqEfWL9o/05MJ8UiYhcTX9BJkBPz1GubjZHS0JZ8AB7
xBdUwkXlKujLBW1ioEpRT/WguRNx5vXDqX8AT2AiaexNVI2xXvOZbMtcmq1A4TuM
cxKLGl3PrxYEXrFgvCbKeoiyu0wpPlCGKd6ljEp8befRMUUekpod5uSL+j16hQsL
vrUo/QySiTRQPRCByqNzPs0fRwWu6jYQoc9oVK8UOUh5YOJBmDUJoFKs5eo9nf4y
ERrfPl93vovOVNeh1u9uUoNUvSIZfIhrzKS6MoMz3AluXZTzLWrtDB02bfVjOodx
Q9fUoVNfRyyKThG2oLK3quls/6qDltdaTHYNDuCn7YGAmIerhcYjmpUAnToftVvp
WdXefEqEMcy8XZ864WziPyGuYKApPdvlfXUr9FvQ7vfDbtGAgSSSkyqAPFB9Qg6G
jIKupOctGJXwGyNTmlJMs6C0vsuElHF9GvBUQQ5p27wLwxsTO52489XY/Jr2m+/I
eJ74G4PFmnXpRjuqy2mZbkQE9EYoUFJVKMwGBUSWWg63TkXwiUwCZioEs5brixno
y825Zt8vqAUrTUKgdEiGs7sVkiTligLo30xG+1K1/In0e8p8hRCI0hbmvkEmJfbY
e7eUDN+2FoeQFfrdr5IbPAVlLLB/ivF8XvSipS8DtrXP86mX1A1r+f/jmRm7/ASI
CkLw6apLuiTDfYqjfolR5XQNcU6XEByA9zwxTlqUabvYtkri7p2NDxPzdOkvK2Q0
0InCqbn8USr/uQhfq+HI145OLU5rHbrSdKFazfEprcVEKpu8SvGahGXDinpXm9hF
Hq56Eb5OjIN4Fu4NkpHwLmduGQrnLn9jmEbWBApgc5rcHo3yqkRzZfaI3HtIoQKh
Z87IeKPgQ4eraMh3gssc7Djzu+Kxo7BBawZ0vkfeNlXoANiUOkOmvLXFjsirpIPQ
8trMqFdR+PZmOAnfJbgqwbGU6kYdijS17k4zDDu36CaJmkwAWBYX91j6dFQwaGa0
XgIOYXO+ULWfZoS4TsbAXwOPVh51UMqUOHbHlIYuoYXj332jG2Iy/p6cJHW1MikH
GZQ/JhhJt3ekiMFHnRk5I2qehWtr0HJv2NOV0WIQ0V6CQ6urWHbRKs8NuBrhQJRm
NmnfxiFoemLEelf8t7gLeSM8f7Bhquf0GffnFV2zmcMwo5QwL8x10ut0TRwE50NM
cdFFDmPDOw+vuz7oHanieGGL1TfOZ6jrgxM067VCMTBU3Y3MtRz912CnKW/Pg45T
1EugI+vPuEbk+Z4XLnCoJDftwIvBi6tGbV98QLurBzqNXIHum1GahnbRA5Pxf2Pe
P7uBIkz3kgs0Gmenct+uflWgevDijCrs+QEh8ooti0PjaG/wVqQcjk4ecS1JXeB/
25fNWRB9zznIXDC9Q3Ex7/2kTsXybBwI06YEu2u3gyPeYtyM8dyCLlmT9Il4U59M
FvJ21n+zynF7cYP3k6P7GDuhgG5NBTA/y6h9ySyN7YTysKU/HBu5yG6gOeGIkasd
5wQ4TOZixdIl6DEYEvVVRWG8Y8nVazBSzmFIGBsZdYjBuc+o6F7e+OJSiMVJDLSw
cERkR21q/xPzVnuO/suZ/baLbfdt347YqbGs2QqY2aQCJkEyLmftzEO+Fzog2B5D
GYh0naoqTg+sA4j1LlQ5ITDEAGxjASudczxKWwOwcv7wtUcQ7Q/Ky9ume95RSKLu
hDkqTOPxo0syNwJ9tl5uF4SXZBH67Jv4gQbdb7NX6dPXPUTNhAayxUiIn92xrtwq
H3aw1QF9lxupoyc8qVgopmBzFR4vxWtze6CWRVmax8HxIRcYBTYDu4L8AAlcj9mM
bry2imkRaj9Lf1EYDPnSccfCl1WQeEjeLn73Lv4zi2Kcma6P0Dd1AEKwrf65UMF9
Ct+FJAZBrsV14HbEftvsl1mbLFaT1R1BvsI+WFZFRrKjUWDs+CvW382rkE3a+08c
Gnix3njcOjydH32oXWLxCe4jbwvz3G+Thdaya5FBkF5Ua6t22WVpcjCLleOx1n3D
I38dzYBe+x3r8Sq+G+4G0tMDV2omVdgYrcF0DZ2qrz0wedPtpkSZS3jmNOMNCWdr
m/u1MH5ADScrYBLuvazliGkkhsCYrhEWo3tFL/AWMluOAtOsoWHfBbiReMiciYAn
FdqEVJz3Ub+c+jwcp5QgPq6R7vHrvj9f23UFOMANxv9rUooWTSKcUOC7UTpWKM21
A9C86C8QwH0MJItHohd9BE7nS5vj0I7qalKeTBRC/CXtr5YKrp1JUiaN2zFVKXgA
QQVqZMun2uSHmPV4H88Duxo48iKHhV1ZMeGa6aUZMYQMvaoI2MkXIxcH/WSJeTfT
oaMoAc26oMG2D8SGVMJ4vzw6K2yQK3HNIM9cJyiEMMflMmDbdp2oXYb5oW5VwbXm
0jhYMUlSW06xYkAn5Gog7MBnhGaKRvydk8hG5dxTNmuv4tC0h2SXdGofMsqEFqyE
E3PfXWT0uQa1dd+EgKs03zw7xQcy3V9SDMghxTjpWW0zIggdw6gJcamk9U9DXT8f
EQzy76wf0lUATk+m3+3sX4LIuqXfgK6Li9d400zrEG1UqSnLpLLmm3z0kq22Kz2p
vtlwcGdYrOhoZvJV6jEz+Fb7Csjc2jA2aQaa1gokxC+WaUCQzIWoNnwtYmm9GHWI
dNjJ2AF2x19o3NgmC5gCIWNXfmWHoJjkrVsOC1UIIWEksQNgbIzyGPFxMGvAdwLC
AiUJizcpqbVpRghxVW0uRAGozf/Z+g7EYu5j8pFczqYN6hYn9aLqZuhFb5z69VnL
X9Ftqs1HPQdulN3i22xAlndf0eVOu/r1mYWWxyk73yAPwZm5pWiVditT4ZRG4om1
n7YTfnDeyPZZGxNMtJSwZSFkZF+bV14zOULhAatEBMERYfXJx551Hujvnw1r8E/O
9gTFEFk7uLPHesStr/r4c579OYmhq/I2bo9aTDv+uO3zHtoFHhG65+3sJQQrYQdu
uQLuZPmCUdmx7McMTDmWKBzMFrjFrExpz8liYotPwqXg9iPW0pNJ6Z6/dx7n/HP0
qs3BUS1O2ILJRC1srx4kkJ78OPVvljQezCMEDm8I5qAPmJ7iKmHcgdiGLxL6Hi6i
JywB4os810NPGyw2+qxvA5EivuIyrh2nep0tkXXsXGzFTdTHM//41aZKojdK20gs
ur0iF+1S8t6Ro7qBDVsa2rHkfAHnPnFjkA30M/MV0m+vzPzmTyiUmmUjbIUBTBSK
Q+OHQfzGcjIG6so0NQNzo9Wz7g2JQl6S3az1xSN9sThk0hXpa+lQtiLY7e1GDm87
H4NlztNhLIzUXH7GDkvqnhqhrEEF3nG2/+hT/l+hyUNDGtId25TU594MPjhU6mNM
q+cZ5/H6+BhroJNG1IzkXFipZmYz5QrafGieOsMetkHXOHXhDg1upekq5EKrqpDo
O7IXCXgelpkD1FqydyT7UESvR8VVZtInkjbpvVEpWU7hweyiXO6V2vCe2M6NWc9P
u+0+EiS+WSvCh9wJ7jaa+Z7NdutMTKH5czOQ41xzntceCdKwn/m0a8Srt6k4fDp1
ZQ21A25kdRHJQ7PFj2twvjwDaIML0h4ZYVrh9HrROSkmOnXXY3CrgSixiPpYWDEN
a0LW0ZxlRZNjyg/AtfebGyMw9221dupW2R6XKQbhSe2uUrNyNL69F0b/T3ijwDI3
tr2ehRep9ziIdjjUdMFivA4mJpIqmRtIzC1yxyR5Phut1xMtG8ddHDnq+nGjqSVa
OR+UNbAuRwKHgTd40uPoeRH1/UI246obgk74o/8iekguqFZQV1/iDYOf4kmjGKZ9
iEf9y4IwwyCn05AzfQJZc/dKK8KpduBAdAjtapd93nmF2d/Z66VQc8i/itVOezFC
aYje9DIljbNWcbiPDIbYngW41LbIPouvHIPpdc00zPVHwNCMgyenRoeKIzEOhnxU
OWl6IJsfnrfyA0Ri7KvL9zWx+z4YZupyia/dazyGB5aNaMahLK1nJRPKKBAk/Afh
ir3k+fFMVRYWcz3Oq4i9J0Jor7payoy5eZiVRHIIYda/2AZ+HzMQU4msPI/KOLiW
DzDgqr0Wdr3b6I2Sxs4kU07rNuz5JonZkE0NS9Qt4r7y8bxzwSuSXeh3boJfwfl6
WTy/+Y0H+VNTiLCBbn0MbW/xEjCsi2hGXHi2QhbnsfV0JneUzjkevZENRTh6OwbF
j/CRn3gBUxQoZD1maZMArDrHNNo0DIm1P0FPYOWnvUvxQnQcKn90cZEdcoHNr2Af
t9iClHTqfS5LJ0GA1DOSCfIW13CYAPrNnpCyzX9XOp/ZXec/H3CCthPLJDk2h0H7
IfKmIYjtH/h8O076kW0MVJ8qrCtOf6ISrCdTnWEO/A9dWt5oKiOmlR6qB9LjcYA3
KGgnqKphKVa9wXHvV/u4Fvwh4yr7GdMRLzFjs7AOVFfiKT3pRy2HGZjsSp5IaTgL
7XbRrQ8ZRpaFtYtPFtJM+IBEiuagEUu511prbRw4V/mcQR/OvE9g0+iPygsCO6IU
hMimtXl+aSvoUR7yD9sdQu8iinDhChpqGSVauQf+1jxGQ26yZ7PZH8v1rHq6bQ27
a7/se8QllAXqjGaWm6x80Pxmkcfi3owq7Igni7A1zErU2IcBnP/7yDXYkRAMJEI6
n0ALWVnmz4THWpzGDhtrhNVWzZglOwthS0yFlJ9oq5ft9RGx9qfd9YnXEmDXh37d
dtEOt2GWrRvDWt3iEj3pxMCdUAaqhOq+7OExnkG69XmJtJVOUcd1t1am+lhSCp6h
b9e2qxg7BrsrJdlzvzc3exG1Lv05P06uYgO8tp6IaA5wqBGqROgl51RTSX3I/VSQ
R1GeDvimaYY9k1ZlaSZLQT4ZYnyhSFfx2sxfyiFJ45aqz0VC4Tch5fTqK+887/8e
KfVf3jjb2Vxbd7ul4U9VDqIB8XSTX0//5BKGRd5bcRFQMYoPaun/vYTw7l7yC3X4
ROc/0uiSa9RGU/mVAcmIWLaCvzMwd5hrJnpeoMEkNMY0N5JliGZ9NkDVBR+IMNWz
JE4hiVj/hWdq6UCT6IOVhBtRkM3WmGoBR/yCaUW4mDyYMoCHSYRY3VcUCIUbYhL+
VL5cjYjYsMh8M+Clf5Uo+ZVNiJt4rwf/AV0asmKr6/fDwDMXKV6xiuHsXuVXC/a5
gqHSx4iGwQ36ezr+3tnYYXj0EBCn7UKiZXWFEy6uxGFdiA92nNItYTlSssw1sMlg
3c6O4vr++w2V4MFnEBOZQkh9oLLLFy6bxZaQukTExk1ZqEPDba1nnv4clEpHS2yn
MK03NUCVKUm3Yy2Wu81HYoIMoz7hjsKpPhUtq+T1dmsItMZW4QmKRXBtxXtu930c
P/spQYd0Pi2QqFwQwMaqfWWG5CuCY2HtqJhtjW/ShivLHXrwbZbk2uIraTy5Cuv6
aq02PBdcB9o4cAWAq8hJgwh9Vgf3LPmpqvSX3OB+J1/x9tMHTpybnWKAN8blSl6n
Iz81nrXCP6BbPl7k+CwYdvzMfvogwC5h2s+EvGRYIX3mwy4kcDB2NXXUpHDXm2VT
jxwxbdgakdL5iXtPlfmRic5jvoOHAnzAi6zrrxkGbQHrmuDTl31U0/QM5HgPAX8M
6O7+9yfXFArVXhLd/yAjBv2BX5OlQ0BOZR13TZnWWwWQv8kvGJ2v29+bH5upEJH0
6b8w6vexqjaG3jTg98l9e1AAncLGdG0MM2jVksza8Wc6OG21SF/BT72beBpo97Zq
itVBSZuTGs/asGEuoqB+UTyx1WYA+Wm50k5YSPP1xIcgnX4hX5yZxeQiFpkbS/E9
he3HSKsSRAWYT5yQaKYBBoOUKLOapF0F4GiUo/VNRTQpztxzUFa64Ta2qV4aQP8o
6ff7wp24ysk/gUZqbdFudMih8BrpvkzelB3iUqXuL6xcgaXBROXqZw8jTMLMfQ1P
1lIXJi8OZumUHE8P0P2WGYoWD/7jofsjH7HxHfxNCxeJslrnAlCz8MsDhoyycdNy
W9MFDsIXeO1OLKemXTvUOedPckm1fCtX4jzoyo5Qv4qcotMajXowQqX423/uKzLR
5smIlCalq/T1++dolH4TVFX1cwqwgoRB3PDZCDvCqiYd1W50pVcgI7X0TayxVzHS
p9A8KYH2ijSG488EZnfHN/pv9IyQXa/1PPCZU97PdA0rtVXGCsSxxOuNMRa640JP
Wre4iRPTf8RUSBpCHO0ttZE+UkH7WhNIgQAAx+12rE4iuZO73iY2t8obx5QqwJSM
6roOvfe9EntV7U5RVd3dSoQOLTtKpfUhvuhWte6csckNZdW9ef6GIL46oi16dui7
zcz9pEpy4C+t6lacE2gQMVBejfXUAIqu3x4PuKRBlAknP3mHcW+9c/jOI7CTgJpd
SkvPZjCtizC7xzx7jz3zWh8mKDCOOQSex9j+sbiJDrze76Iqs129zCdYlKErBZ3N
vnsqzBGLVgUg8U5w6gpVD1SV1mV2+Ch8jWKPbtu27riunsVE6hdz0aWWlDQNowa6
fZHbhRlaCzJ2rGk42z4PaIC3jYgw2Nt8z3YWZi65aV4IkwbqURf0GeovDrg+2nzb
W2ldaO2AxDrq+XN2GFLfl7z/ZcgxelUbIcCIoX+Q63G3iJTQKgPx/qNO5poAfjFx
uoRnrPFy47UHodNZIYi85a0TxMpROlQKD30utq5n6hKtJcqqfVNFHB+5r7C70jza
SRZ5XQRGU/cRszOFZitxFoGwvLrt5oYt2nlqFMsQkm1c5/SjARBmRwtm6okVW1lM
+RdtJxjApVF/db9ce2ZchsC4jhPN9TmNU7/yrtAB466f/VQAODaE6NaAg27Mh1Pj
kea4aCl00CF41A1a5MtRAdOkB074bIpQMN9oz6uAXyLoNlFlcheU50rTFc2DdlTQ
6+9gJES4xmVuodYr3QPneMK5xYwsRvLyKbTp6BWA643l85+rpuMlAQ3uPJpxOckm
tvYOWiZA4r+k9pcizZOTILDAhRTtXGf46fO1sCcBvHDI6bvjZCudWBrPa0/h8h6U
vjUfJRqR4h2T9iYBDpSqEsC+JbElQL/nfbYr8Ue8+Yk7nbMs/5DA/vzPiE3XLWfC
+IvivVx7Vy6+p9ZKC0M3gXG2kaaSws33p4cjuFGp+SHjQAqdyWEul87E/Q2tU5Vv
6hKmwAEj3wXKtPt7kCY27j4ynAtlUbs7tVUM/mXdNHiDgtXeHYWIjUBxKZKybtQa
Qz89+uuoT1drthPe6CsxHq3Cp6jlj3ZH9a8BYE1wHQ1/zbS+CMiabqkL9QWZ+nAv
9W7NqDdV2/BHtrdzkZzcfxrR2m3l6FoVBr7gAiQpVMy/j4mo+8Wk/OYqx+5acIcy
St1fOv7G1OW1ohmTx0wAd0rVvoKxDR88VPkCEhJtG20LLuffB1we9CsO099CX1Qe
/TY0lieHnAmTwK/dmynwGqnYTdv+cFe2L7ujzfJiwVX/iQskbdR5u+AlV4eOp3v9
UAvqg7OUH5ihPoRRk2z1njbrHqSOBc3lQ+52Mjt1H3MOpNtH99hCnJ3n2Lo2p1JZ
2eLoLcjzHzjBY9TUGd3AhSeks0JDjVGjNVNc6g1tsF8wzzlb806EEmb2SUy4sD9e
lMdZo3Hy3U2FseVnZu5UrduLyhYSbxRbnVuyLW4MePvCazoBEzQYYLtRvjgKu+V2
CZHA7eK1fRaXbQvqNqXIYKHRka4OJktWzb9g77TM9aTMez8TcOkkg5/giRNItBfE
zKmilzpeWVjphU/lOeIYUwVdetlGo69+3bshGV9ikDX+y7XE5q/SElmlydaoAiat
U9peUvwbcJQUUzv+DUKo8FYfs7Z2nq32w8EB2OjL4fqg3XyTw7Fef3uyNn36J+GJ
Js+WIcFjVuNpegt/ttcT58KA8HUeJx32aKroNnk5hNVmTYKRyyyXB/cpbWSRzfM6
DqvpJYOTteazWjqMh7ZRwoQwDaSy3mq6PA6wSKI/sv1SXVfBElF194e15VQbIlPx
KJEGyckISGq8pN3a1R1v8Tin7/aFb5lD62rV4oTFELAAWALx4gxsZIOHmfC2IQam
+WIJs7kBGqni2yzla5S4l383zqA18ZOM3KoQYTTFiC05Pxz9SiB/Nxtq3pIh21zM
hXqm5+WCFrQCOFw8rEza5b3RaMX/P4xz4yCTyVaCmLB23Q9sd1jtOM33my7UG+cG
vUn9Eq/XOyqaEvtqA47CwTvHbodk7A3nCVrkggO0pMDB0kO7Gf43qWbC+BKs/6Zm
Ev7zien1rrp3x/qVjD53YPebqrm7XWF5UIBFOXyZfWpu/Zt0lXIM3ODpckit32Jb
jZxaaoiHHJcAwh9ms+vejdJrTW5mNn5ZFUQS6cBDr8+LI28ToZLb9Ug7dmfysy3C
DvvJJ+IYTekxjAiyyKC2rI0VlXasuL/U/Kb03I01Ec8Nx7h2Taq3jKKqboUlWzOL
iHGlg71FtrLhZmm2i0wtHih6mt8X4XMuZSNnegVOfAXQ532EcPmo0WOmgozY0osb
B2+uZy+9wGP/JafU9+PVDQKbPJvbQUtGM39UaQtedCzD6BaOtLTnUhfrybdSBIRG
iMsVX5xOF+MdpdGXTtf0/b2S5IWv+f0M1NdBrRd9LUDBfNoO7DH5BulGd4z4qa5d
Jr9Xh2CCwq+giEl3K30QiVxCHXonvPyCJfD7NFeDuugZRTZSmzlAtEt4NZ3kbzaZ
Sn+4RskevSU93NNL03Fx2enAE2BV8srFtdzhVup9ihtI0TXnVfNEkNSouT4RNHzP
X2J5KCzZDysYuqBJQInwf16EinUJeid0+Is85jesjU3lIAD4c0r5ehQmOJVQW5Th
n6yPzoMz1q0pJRjZXzKqJWAST7DKd3ScGUNlwGCL4+uicdXyvWTeYZREP2rWf7ji
voOqC/u3DwYfvmkLikM6wE44IjXr59j/CSnyjxn4U1PqKE35ReEzi40MPPVALjah
MmxEWI0WdGndsbtREzGHsJnT2sf6LRPmEjCdB3Xas6BACU7/rfAphRZE9uYfNG3e
aPs7i0fGS5ke9aHrldzj2vxySbWe1w/kbadB/KwZdVF2ZB0mPWfpb4GPtrLBZuZA
yT3VGrxNfUYZNaXj5ILFw3xmakNfBhvvbNX6yE1SCSRdEmXZgkPDtHM3MZOSdsQN
jmtkIiGZE5aLQXt8AA8uSynpNS7+vxWOSfjBLL8rrFmmLmxtFvjLA2/5LrANpDsc
yhX80e6tPoyn7yBPlAK1PHSUWGylhh+qggzd/fVpK8OxXgq0pMv0tGrD9y+bYhQF
wSsS9hgQ94fGGmn+2LyPoGwm7dfuZF8EcAPCxrGyoWQv/DcVqaMD0PwZi5cYdU5g
oygkEoOTis1bDbzwRx8bATuwn2QJrUPm6wbxft57WvH5ZD9ylu31C7ESpI3Q9ENw
XNasaFankbet3qJ3hBJ9v4O7rs/Ybt5GAYsvNHx9ExYj3idRHCxvXAQZGEKT95TM
UNjex8cIlmRZl2YsfFWPzDDmShyxyCdlm/8SBtfDH8j2jRnS8yaQ2JWbazV2P8kD
BY96u71g9UAncoCPxvl6yxlrWv/sYHCtVmp7czKHs/37iHaHvQNouc4ztmcmPjOu
bN54kTotvuUJpDluaFk8GlzraQ2vFLSnQIPNbWNgWP75XdCcnYWNDSEJTsYXdwr7
tqheboskB3kv2FIQReE12AqfGx9II0F2vvy9SWlvQ5IbMCvkKsFfHxgPpGBMAq6t
ieZaSenkG+dqMhGMNdeCX2t4gv85FCYOd++vb3hNPx2f8k9UFfVVL6LosS2KDxGI
B41Q4lNMKOxV4ubkAhnjfb/0P1LI/FUng40taAuJOQDY5F4xQFaAhbo6P4ha0R3H
WF3c5/ciaf3qsxUnbCoZFv+YlwucVfEyS7pKnfWrXuZtkvdkD5NDNeurP8hefkrm
hNeVrr71An1xqgDNB63lpyPwZZmHM969oNSvIhRAtbDUfb4OeiD4hqFC1mFajEJ8
JbgAYvDP8irI59PwJ1qQ0yfjWImt3KRaBFziA3MsXa+ohhj/oY1gw8o7jlQdCGuF
1ujEWhzy7C0qfsIpJfC64G+8vb3ESINyl0JyTwndGkBMiEhDZ0brWCD7HU3V9r5t
V7j8csw2GPPyBJZLGypc4kHFT2mb0n9RfZQjDMbMcqWfVV0L6ChjgPEroOJ46yiM
4KWn6/Kmx2YlqDbakXfFdFBioqEknmjnFi1n1C9FFHRhPqs9sDizXB6M3U+NV7vY
xeTptOSWqGO9N65Q45qUWNhg10JZH0ZflgdCXbagSSuoIGWWx07Dq1j5X3+auzEd
KXkOrsnOxqSPMNdO+WLaBc2TwcZQpEuo825+5we241isYuEotF+gHGO0TZtv7sqK
uAmQSwLjmtK4umADmzndSfWyG04+ysx0qikbDAkbV452B63aOVLgfZmhz3IUAYl9
R1iL1OtvbO+b49FUvbiRvFSQhlsJNP70qdh4gJduJ/9MG18LBL1wrhIRt83C29JZ
G7pGv+CGq3DXfggGMHExAXKuhYL8Op1YEtySny5YfTP+7krOx9v3A16vtNEK0mB3
IKotZSWhA0i5H1tHnP9njZgyxW6bEDjZFv89qFJZo85//4mW9yoTUe9QlifYxbkg
oMvszfFxRy4Brf4cXVUqXvmjzJZTk3X5nRYsH2K+himnAdSY1NNLXPp2/kH7m7JC
XDQjalocWSbD627vrFSmePOadn4aOlL7dZsMQGJKGQpuDfxtuqHOIT4DfP6dOKqc
BZkkogQAkIu+pN6Vew3q7hZCS3D7XBMKD9m7dwhUcA6Wz4BacsZrtherb17vSoGU
YoFfr0WIVL8AaDNuCFxgo2cJ5RreoEs9rSMNru9IXeK8ulv10is6Y1ufBcZA18FR
uzjke1HV0I9eQmOeKG1I4uyx1HVdLgRD8qcMicN03YK/wVKjALZjBtSm03XuK6KZ
T3IumipW1lYkZ154sMHZeY4x+hTu4v+PqrKuW+ANFfaDhxVv4qizGXVUMdO0lC9n
Tbb27I37Ly+OT7dqgx7lKMMCr2JqbFsN3lVMXAqoykBlVmVfqJZ35NBBbRYHKAe3
K/Ste/OpgcO4447kH2wiDHjIebiZXQBHH8ym/sZ5sjGTFBiWpVSRaI59/jducZAd
iL0Ff/sP0M+dZL3HBkwvdry41/nvNdE3tUAB2DuR9nntDBy/S7mdwAjy9pu6QlRE
S50i0DPzndL7nYkDEUU1BuS8f1dBXD6ORRX64ZOpncVm/RhOzx68NmDrG8eEF5LX
GHPARA0OUSpWRGtLWOabXddvpU+NuNOuUJQ5REzrEq91Re53NC8QvlUOBbFvwpqR
PXuPoWICMtI8nfAlT41vUUL1AxXp4gb2nh/v073JNNNH9DNBT9Antm54zinCdjMz
VCdE/ErRxt2AInkw5lumgkL2Iv8/Xv7qF2DD+sVHkWWWml0ZjHimUP+R2aIB7XLq
EAvHdmWqR29ES6khyyKAn090I2aMwp2V7NOxy6hWA5ao/O8Wj578kZeyA01cnwvm
Owh7ejSRetomKyLBb0TScNIIvjr1smR/QoLSHO3uyOkfdAJR33vJhggwnCq14XOv
mR9CyrlJaYtTcBM6ZVW8l9NLux8AniX626BEmk8G6LDVwAt052CbcUCWSQliiUy3
GN+GL5iNrYl0HSgfWG6MB+RgmAhIqK01WVsRVogCxfS+1yArmIiI4jJs3p+IKydX
RD2MLreBue0XEubH5GgSwMH0baF7HU1GVGOe8qwwdirpy0x+uqDJRuKlHMABtuSB
N96SaS0EK/7WoiZHKEEdE/ca4UHli4mlV8Y0J0s+c4eclpxhk9riGGf40uFTwXaU
WvkWJQvHiJVSGAw8xJeNc3/eLxEC+QtslEFO+ppI26ZBZxR1D8OzdrzR9UR5sNGa
r7RZIV9Mb9h9zWxJURQFO6YdeuwYUrivz7tj3SujR1CKMiwBt+TNAmNzSA1xsZGa
U+BLvKL1oznzSFbcd0mogWxtxJuZCz4pQt9ictFwQImQJU9yxJJfj+vOCCU1ba5h
tyTS6BC+sQYJ7x8wE+KZxjFwXQ4gDKswTLlRff7r458WxOvbMKZ+rlQT3OZIsQl0
BtDsiHmhtcImmlHbIExMXmheRB4EzeJiktRlP4Gkkt9p/kgJk4j5wQIVgUZfqlZ8
91M8+T/vWHEdC/AzJO83zt3nqBmNN9pfSE9zuVhWIuDvvb8G8iJMhkpJ60FI61P2
XPyxXQ/rpH2Mzzxcdv01NxbZSz5xAW3x3uofbhoNmfZ7ErwMrG05opP5IyftgJtW
8GFerG9JFdsWYH6ViYmnWXoOWQXyd2V+m8bUvKMXYKC8jC6rB+qQQV8extaWHpkB
kzlYv8/Rz0PKPrWXQDOhx5uYFdH/R9Ntkca9jkrFbaeO6OQn22Vg08ln75GqkuKR
paA8Mj5OMfV0dzh/o6MurWCdw8g6J1NI4EJxlWJ+cP3dmh79/pEILTN/rDdbmEib
4Y8tUgCeeDWBUTz5diH07Z+JiqzHGI7LKM+y9U6XtGFFDyo4ENuvV5XnHECm/mCe
6y7Wfk809nmuSiTGsLFWSCXtBZQlkfzd5R/QvHfdYLo2eNbbH0EmzCff3ptBIZIL
hINgQZpn9v7qe755eSvJQC1nkYRyagQdHq9lDzpyvbB7rnrRS/0VZYVoji6vatNu
Uyu8DCmhEC36ELhE8xQsYbyzn6uLt9yt+I9XxUQ6eV/4788dfx7v74EPXF5RE5bR
/PEW2598Tjy1DxP6QCcxumCX1HJt69X8x52+HiQIVndaP6Ncm/J/1ZRMsbAw9eDr
dtipldbRIICJkCOPbZnxItRY9MuwHCte1P+20xiPgJTCzZ4YnpTKiKmfvf3HbY9q
j6+090ak9G2lAFwg91yCrsoGf1bdUzXbwJAHaXNj3aM1EE5jX2Ci+zlRzkQRuRok
+C0uTXmnT+FO+08gpDvx401oh2xmO1HG0kbuesMl4pmVsb9T0WdPXrQJuCgRyPbF
wRIUunIpCR2J9gOrCTPJkzWM8xFCSuWdUx289qdWFRGrwXZCVPDVS5qaqbrTPgeh
jatWEZEPvSWmiDjDB0UWlMUZVTuWSkI3oOtAWIOn2+XjGZ69f66fii7YSKTHMFKt
/mGPRfcuC+WpmN3sHrUiEq/w52ZvsF5W3Kzm2gKQfRbW9AbwBuvBPaY6zPDzifNr
GT0zjAYX89zl0rQEnG6Q56YieH4tmdPK+cF8WyTgdNN2EyzkGUW7rjWxoqIO8iZw
kcPIRLdI0mw3EmnfBN2X1mEVdHuPBL+Dz7begf7KsOqXa1PgeV2DZN49nreVs16l
Idjb+ASRu0CM6cBljSCmNRS8y9DmrFcb6qERcBHnk5RotADuy3THQodaBr0SIiS4
Nwn8K0IzfxPo5JyfJBkNDuKkwMRwo1NUMJX+RPHWA06FSv8Hp+eINqodmpE3wXAK
McsRdMad2RZwJfRpAaf+0EiNCQFVSxFluWIOMT4n9gj4kZxJLPHwASGYg7cyP4go
1IqFRqFhmTfZKGx2NuI2u7bszi2EFEdSLNxsq64B7u7w4Gn/ouEjO0WWkiifB662
MWCmAxP0MpR1DGzFVfL0zBRi+jtnm0LKp/+krSMG1DMGGGalF/zMpcCGyRqtu7Hc
MxsF05rOedN8sKVvp4fJKxXnC/joa74nqyT7fOFK+HxBj0hEEOPjy3TkYYD59BdR
2Wkit+sKKjwYIsyYMtx85caYhqiMrfSY50KEudlYtbyQpLo+7TEV2xJKDfIPcivX
P7CytNOZjbMLywpoAF0CmA9lqsR3HnSKUy8XTnDurvhZ44BYKqJypVmA57Rmc7H9
c5uCoXtoTotdWhNp2FR+USbN0jSq356hQoCU3PKRIda94afaqcmGCGBFHEi1aJwO
9Z5tUK4m9eEADw+P1XaZLBJcGUOfcwCuJKjTBIE35zu3B3/z12K+at5RNpbUDK43
1KdERsDPONaPip0OyUz7Gdwt9UqUJv/F2chHQHVO6GX54ixGDRzEfaqHqQInxQRX
KJfxSGsQ7bemLXMHwc2O38g4ik+G/y+mT471Z5GsX/sQCnjeac9HTcLP8IGDMNIJ
XJJMe3QZy9q8QsszuF7+iLS22a4DPQjCtCBx4TMFVBlVd1Vfxjo3RhKD30y0zp2u
vN0eeVNzMCLVPv7Po2SqZrfZaEK43UUoEoIabVMOUybre/lAmg6FJXFjE9vgC3O1
PmSGJoPqZcQtgnPZOtx+KWZhdRTPH1eX7qIg+srWslDFMDriB/QjckgXQM0lDCy2
bvX/VvmDNmwHDPm2s5OOQpNvTAyeXZstJkBKqeQMeyKtOdInPOQYX+Y0upuK7aRG
kXbj6TqudbqLHUlWTUjkC696rHZvsYq4IHnAQ7Uz80OZeU7gdVkzL5GLIkQksNuI
MD8aqHKKj5DUk55C7VcYlFXw8Hqtc7vy9fYLdayPp8J42uhrnM+TdigeCClGWecH
Gc8zBOYmO1358mnvcQ0AN7rvC4Dnq81b9eS7/92nz1zTaJ68Us6QBNK1TiOp2zG6
33qauYro2VKN46bP1iuhHnTThBAI4lMjdp28ZJ3IgljeXW2HRV+XzyqUpguYOhPU
6BXjRnUtA2tRq2Fqo75hA3dJ3Q1YcODmIvc5DHIFpiLUEZ1gRLKt3gh/osj2p43k
pVmJwnCpddz+aZ61ZJ30jpU26gZ42UvNUmziAcH/e8kyTi3W2KUrM7DfmJJGaDci
FSs0fDN2nH2+PTcd9zvmTJMemaj9yyX6MjMYspyu08SDIamFUANXK/7oAU2GAENG
YyhANhnVJodOqh2MH0R2BI0ouXccYB5XZzoXRNU3pNpil6nhWgDYGzUFLPD/F9TF
i31H9L3xvKvWdRjJx8hhm/edIKkuVSsOkYOuaehgfH68Geevuis99Zg6hbv+nvNi
ktrK20bxobbjynsdUwWtGJ/tzJI2Pd5NDJuch/+iKh76Azo7k+NzIn6g2ms8mcUH
v1eImyFtALT/Y+gT0+5G0N5juZaCMk0Ip2xf8V9UjpdjH9pXaEKnLQYHhX6PYbCY
ndFC1cCZ9jLc2s+A8iDkoY/eZC8cttPUBh6zAlxUo4UxVpcZtl+0+D/noriQYImJ
NiN8Y8Enx7Rz63JHvdEUfLb+Wu1anFhEqgh2JSAZUmHmnHH7v8wDL6ZYvFarPyPi
tropW0FbGB5ChhFD9yS3oRAorRo9L6s79nYgPk0KYlGGQ7ohshK9oZUZYLg0Bc4N
epoFGLMCS3wN1HCFOXFbS6D1XHJYYthOt/rDHNd7UZEYFU9c3yLk/gTpNPjoPK8d
zq5IQzQv74CDvvlYQ0QMTJY/pZtaIgokh7Ebr/5KDGJGzZ81EDt53/T+6rrUedDb
yicbrwEwr9X6q2PMlXnRuK45xg2oMe14Awgy8McQrHYaMpql+Bj9Fn9LZCygWZkG
YpEsUalQvZpuZiC11uOHX14/FMwvcS3A2+PBqMXpVt8XSr9705j/KfIriZyVDB45
P1ZzJG6xmqyTuSHToLL/ODRqKNimMhcdNGvgsagz6xwj+iCBzCDbPSFCtZoRJXEi
T2FDsKhBqmlZJLPLHlS3ymNmvaktAf1WTkhCRQaguvNDEijHn0pux3A0lOhWluel
5ftEGMtO0MJilA+TnZdWwUSiX9HQiEOy8H4pLhWJt8NoPt1G8TZuSwjA+UaqdduQ
NmYF1iw/3vSWp3MN6+2srbAsIFYraV+S+VFbeU5CfcijE76zb89ZqW+5RgBqQqb3
paxAXEhFOgekLH1bh+apOoJD2H2RqgtXPhfilnYrpGAMQYPpedzRmLMQGbg1vQxQ
7OcDWWbdhwmoDZo0e1r4c07xs/PQuMqJEIIsg3viB/WdNCcYhmP1vEyK2i9/U0Zb
aTQhidxCVPCdOrtO5RRJ7qWEHuGZ0gXfQo/9FWmRCJ2v0vgT1M5m5vtq8moDE5bZ
PmJYP9UNkh5UkWgznfoBydDg5UuwX+Qm3eKkdOe9D3fHfI2T4dhi/+aDsR5laubQ
AqC/hCbatiXC5zHHeJmSg32Y5wG/a3OI115M+FrYjZNy/eC9MjI4P5dskT/Dhitr
6B5SESvDcYsPeu8yZRjdw3St69FDHaluy1peIihPRaUbrc+MbARmi5ckZvHowJad
GiPmVF4DwOZwIEMfKFJvf6nZXtQIC/GOLyZAjtheyz7dOIcmfURBL2XcbdfB244b
VOaIymjYGucOZ4DdarsVAPzM4Ejxl9fo2oKbewJUdUiZ+aDCaW1/hJdiFe/1MbtI
3MqjFMySxZUbwwie0Fs90xXIL/PJITCSbNj3XtJVyAKKNBBEOF1SN2wvbK0Q/TU4
pZRbYASp4XJEze5WDjGfiDJdNduEKNMj1BDpRHG1A4Vehxkm3e1Np6PCPhcO6qeS
EQRLUDQRaf4KyawlxgYzo53TK3tj+vhMDd/8yD44SJK9aru9/5xJMMqP/QkLLqnv
friKAUiwIrSt7zkCx/Kx0z0cL/l2Ai1X6w+nfdaU1eUyL40rZwsTbHt5Rq6L5Jpp
Q/QKJe2h9qqh2Dq0/ayfzt112aoXqMFbgHj2AeleKKG8XlrlLwzuqE3H06tNOL4Z
j/gOqrSm7+HPYqTfAnB1kurv2ibQlNJC3hlnZOdP+C3ym27kTetxeRtAKMQFL/f1
T14lFQTmhrFcL6tErNLxpNqozoyITOxL1rob+wUzolr5hKTgs5tbdW7cy7/Qvlsy
Jzj8BUvc4dzRM9FfHAbsJSl0k3p4nuAILMB+3mBKAGI7ZXTocnfNLqLB0UGzFc3B
GAJggFsbBQEYOw5ptIXutEsUBu0ci6+O9vy+AtQ5ypRQOyIvT3p6F36WPeiu4BzZ
Rd4icFbV5I0kdAV8XHr2VyR7UDGU/VkmIAszek5da/CcN3x9mcX4ucnQl6vYlo+Y
3lmekkkZuxPbnsnuMy73ugLOv6C39077ixRmplJ23imWHhOF1kL52p8UoUHwr4kx
5tYaQ8h0d2XV7MQ+Y01COGuvuqDYaf+cQLfPlLy3SWnI4fB0BanEkz3BtOpinBUQ
VVWXrQ90YLuRT6GIC/WD31c7ieCYKoGb2Cj6/DfI1UL4Zz18v30y16t9Gs2ZTmaS
60HbsC9BbquApzmeILWRAzAhBXbvZCnpDDLQOa+uZBML0KbcEvz7WXPtH2X0XVn/
4xhBsEQfLZYMOdqvJNCSxWFECCasFK35mNLzKLQbCYh20qCejC6M+MgQ/YXi+vKX
hO6Je612yIlmnVlROzYLVcIbWi+ktDnV165S5H8O3umD7G9MvIgpTez7X9q7fO48
JNNUmS0lN37zRIKDQ/luOjaECxjPeECY0o1pQhrAp09Z8SPcXW4HdzTxUbuRhBPn
E7TcZ18j2QVkqsvdF9esGyZ2h5TWsVLl+a6+levPYlei68aVl+AOj0Rk8pu5GMj7
rjyHUqA11chMza36j6pm7vE/x6P/a51+cElHo1i2EEOLFBEEN1jdyyOuTHk/2rlm
QoBcYBI4OzeVXecDbr11WP/D51NQWS4DWVnDC8VC1nR970suyoWFLYVg/eOfQuJH
xVpe7DjlAeBHpOKf8dMCJkWqECmWmklh/u5CpufuPJCT0LwRUyhLD+k/QTAyM6yJ
yuZoYO4XgvKG1XQbA8THz+SZByyzWSahi1uPRbygmCf1Rz70mIgkyo28I8cSCLFP
9hJ12qrUaFB/bS3Q1ZTkNId9tFKbU0ZKgqxM9rLNeWLeZ29vLnX03PqzWrVbK0bl
Yucw5th9NWrVRM9JxPlE1g9FSSdpC7G1IKjiPpQNLJ73t+WM4/0eIy2/3BGVafhK
U1vC+DbTkeKABl3SvfeKlc+TU7ppcbVEH8jTwg+A9rQz5WVMjc2JBabT2eRETqky
pibOSQUIAIVsg0Zn1wCiODn0TEeDDa3ki9SsUjRpmw3VCUkKAHNPO0/ycccTgljA
L9Iudkfr2Kz2NZLLL/6UwTg8QkSnFUsbVykWRzU/U3IRJLve8pBtwR35gGEBggwK
93d4IivFhTKAB6k/meFPHjhVvALxogfZI0V8dWBTrVGQxwFuBUwDz0ktlmRwewDW
+k384N0HDjl+N/s4qCdqwnAauEV3oQ8l2NLW5DuvB9cvja8g1yC2vkIRrW+LqIwn
lycXY3BUe+7uI1dJFJZ5p0/ge4FrAUopFMhS2VIIzw3KXp0wyFv61fa9ax6JHORu
KZxlaU79evCWJeU5MwK2rSqTkr8yR9zV/6sZKNovusilFdLgZ7uu6e4+th8WzPXY
IwjqY43yetupZ7Odx1+1t8iXtDTg84hCF4l5ndjHxCiVQvd+MADEkLYG/yJLWYT6
80hoatguMA+Y7vdZbw/YtDGbRfCI/h6ChQ0aki2hRzCu9bNodeOc5NljIDcX0bMo
kNmHEMQoBziR4+K0jDlf3L44/2aRvbJC7/B88/0xKDomYM+1l075jIGizI2wAaMG
SFSYV47vS7/iM1GV1VA8RYGsIKTr00Fae7MObZY6MXZbA9KZPt/huK65fKSTi65b
ts9YREuf0AehtCazxKL13dKOOLguw2DhBsH0zqwrzON+hmNrlkbmkMsF7OF3upe7
vSj+DEK/kVSogtTHR/ZEieRF7jSamBnuFlMewFBslwiCjNymR04snOk/cVbpHxeh
HQk1XC0PCmEj3gJRyJSGQjEg5WkQ+jGCWyUesKFUB0jZECkwl3DmjTQHh672BNnY
5s7+tVbEpFuubSqsbQ9+EFySW/9Gir01555QOU79iU1ZWstg8Z6zRIcMsQXyQsHY
HxykjZQiaxYnsavpU4bKhsi6k1QBLjVxw4OFl2s3opnKtHZFOUYPSN74aL8E/P+g
LnLf0hF7kzwR1mX4DwOG6gRjuthL2q7MkaVKWNNO5hu6l96CQI2XayfIGeL7v2Jt
muNEX1a9QJ7rPRE/dhZr3hbW7ZkTSl0qx9eAe5PaGyOUDlfOmTilUJYH1EKxTK2T
tCtdE7eGcTRAxM+tQjvdgl0hXoxrJuYVS89YvDOB0YUG7l3tkPImHfsCNRJ3E7po
qFRk/8mKpx6wPQJlUHlp/eDbJAR37Z5FaF8YxI+9dQ+c7jI3CrNZmFP0TRUDldYZ
WWcsM8RzW6Ip9HpLioo5jdfEjvWD7Aa9GEHQ3GuH0cQKU9Tb0TeTX+V3569SVd/d
KEZtU2z5+UnFuUs1hlnOsxs1U3hmAdH0T8VfAQIAINk1ZfYC/YOlfLU8nTGYNzBn
wT3zHmOQr2/8lvM4dNeOSUsObF8RE9SRcABmUm2hOY+kwMT0fQhBj04bvIs7LCBy
LLermxh877loMfkBue4avRUuW9v9fWMDOMW9zX0PecVXK4yaHaZOJViMzq+HWzS/
NULxEb+8Pk3hqeU4CnIP7RbGbCUe1kcCTSFxZDZoXdyZH2kK2BTWK8YXFE8M96B0
kg3KH2p1ntEIdKt2UffXvdYsYIITBuN/KEbPcOAAz5o/clLo6HeqfWdiPOjEXdnI
REscNlBpINEAX0CcY4S2YYGaVem+pac6hVVupoeuenIxhXP5OCck6mIlOgcyCF1z
uo082WBJF+exWHH/0pLDFlYeRELW0baPRXKznZbaUQIVoWq0x18ojXZCwmdvuWV5
ukAgcK3EPqhD2adJw5SZ56XBf5l1H60+wg1Oj43InOZdlKYHwBmUosDoYedszmil
jLef/sfnYgoYh+nJb5iADSIFINaMHqNB4sW8Lfzuryv+MtY5taI2BhoFqofLJhpr
el2Bdo/wl6+KOf6xJk9gyDcwk3emrMs7Y/U1CYwn/7oR9TWZrjGfHxOw9NIk6klf
pOehlKUrHqeIH3IxtSpiQ/Sii+TnrnEQog8izXvFRjhokgpGI4SncI3GQzO4ESTW
TMA9YJyVVdyGou/xlH3LjErw8qlr6ld/m40MXfGyvPQR8LMyq79cnCCDjZFZihFp
bSOAu8LpC2duRQyl6wGbcyy/GhxP8BVbZPPPuMStbTxFKUQEpmhFmsvmpOcAnX5w
xL81l5ayctpxHt+vVL1q4ti6mH8cdW1hBFG0+CiGq0JdmwwRdAV6ecL+OPKG5luG
KRvz9+9tCsW5XCsorPTWh4eozs9PdODFF0ZhE+TzERW17KnQielRH3Av5lcfmtek
P7A3YDUnv4wCHJFaYSq1sXzj1fhUWj4itNm94E7YK/TCyjb60SL9jyuiBImlh2l1
NTeKdd6CAsOTAlZcziFlDPimlFTlFZqR1bJkqwuNL4nbp+Qu7NnyXvbvNqqbUBHV
Z25JdN2kewRjOuI5weAP4j0svWf4OoMl7eplbaZbCLgY4AxdxkXx7qEKRrM4i1TW
99nFUCktcH4r48lIwD4T2jwfu3belH2qdqnNJhywTg9+cA6J/gJLb/v0yl0hbuho
0bKOXz5Wcp9+Nlya0ZskbmO7cnH4ykw4+AeKUCy3/1GXNkLC3ui4mjSy3uYN2pCv
1YDEmh6dil/cMLLgiVxpwbCFwWawgT8rJaiurwOChqT6Twv8zKIxVC6DPfKQRrzP
NpN6WPcyxiccbGdXINtChA0cjbOpkNNDrKnAkQS1KTVvXiFtVqOZIYyQTeue3ByK
qa1GOUwyXpkdhCIUOMh6iDftv3BdJZDCwVU5xEJozZKZBFngZaAa9Yjey3K+M+zn
NYutp77EvHg1pIrZKECgyduF4tZiIMKTGds0lf+TM+E4BOc1dezSbEOsDM7DHMGE
UcHW7WP1WAGzVBgfuZ/9AJfrnJ8hDqUcC4kEr/zxA9xqhETsz6PC8sdwlj8GVqUD
gvFeuPlr0NUrTi4CWL8DovODW9guQJkBn5bFlagUSQjF07OBKu/R/5jbfiPyUdmn
59i42ngEaGKUgc9OMbl49rOr/2r9dp3cXjfzn0m5PWoStKVi1ATUmEh89yvCgz81
eGSd8+b+jPCMxe1uPCwbbx4kC0dOW8XIOMvt0XBQsrfJNreZxPS2R8qRPd0/qoEx
llii2xcgV6vc9FBRKHVS8I+Gu+jyPGasx4tsPhussQiVLt1HPcytuRZlgt9jLf0g
k1BEqvmRLejFfXp57+l/vyMjQ6mWAKmD+WTHLls47PYGebwPbT8+At/qW9a6YEpU
VWGGMcjCHYX0KaIZ1q2AkPvr1jayHfrosqwtiYLgb7qht2Sc0TVS8La2Yi1ZWwCG
JPKJfEwxIU8puz3zSkA6uw6EWX/q73MhHMZ54ZSAtpy59mgv2pABIWvsE3k2CU5+
CVup+7CDndcrzJK0NyiQUOWTqzcWWovkYUgpnTmEBMit+0NnSDaODpOd+oW6hY/I
tYpRURzUoQrCZoX8MY3SqTqY0viYpx/TYe3j+G2xrr+DEMor1FKs0hYzLyL3aGQS
m31SioX1FXHW+AYPDfjF1FU6WOWvCdMtYf1vGLutgW6xkNJunt0ca+qYb8ZQjp8G
Pq2P48bnf5z6sL0Ves7IToR/w2mU9NqB98YQnRi8QdCd3Xumkk7aiqoyK+2WFkRX
8PT78dE5Lg9bvzxYLqhe8cffKSUv7eZCD0T77s2cZS8bI3kKzwj0usMkDGmgts3s
iaUTlT/hEm/5buR2inPk1j8mdHPzAL8Q5h+yF0eejqcyGE+6mOx0aWzAvV9A4qzj
JGRohEi85hEEFV4WNVaIEF6G0/2UsEYZbqKNHYxOyEswq1EeOj00pNWGarghhHcr
Z4m31KS6UwHZ8Jl6kBEz4nFVm2D1sjikfDd2j27RYdXB8E3KfTiz0o79kvEYOdZF
euUMtujhAYcRJ5wYQoVrvC6osLMjAz3KIy+CUjR7Ux92msc4lx8qH8He9mwNoMTc
oClQhptlS/ktD3ImmRDPNRBjM9K4RH8SU0P4/zkGwzkE9/xAPREUiQw0MsGPEWZJ
8jhP3LUFJEV0jIJA1Za0w3Pm7m1jiFW45Iq2VLXOwlru4DnVGaQM9jkDmC1wmwLF
I7ttamjq1zTBuW3zEECC1zxa18shUkbmj77p2Ymfs9wS1euVttYJ8CCsWcnXDNDn
WBcnuvSG3YjvqtiAJsCq0ofHOYx4rhtkgAFm0Ypr+u2WJZ6mW5wnNUSqITHSx7nL
DLp9cbQFVfCZV0yeAc76f2OYHVtJlwaRYWjEs60wHAlGlTIeGbm05iQiRpYypMQw
EdC/QwRNUoAuwT0Hd4xpz1TPHj0W9mBzHqpJP3hGuhEZrjDnDoN7O5+WrCB0UpI/
t+xEPzvPBjF0YasCwb85S2tp+JCyc8xf9dLpVVRNukL7qOcjNyqoSVUrYUOoxtMu
utAcyqu5nGAePUwYJf7XSFN4rEgntX6xBICWHr8WaTXSjRJk+k9dt31UtHcHIbbY
Hq0eRGnCazZI3a3VzyvEs1jM6L8g90o+/kp/qgzi2qlGhEPtq9tXeBGWs7Usd1DV
jd8PeKVIYnVrO5rfsaO9WqNSsVNu09Pn6c53jZ1brOh5nyztuqj2LFsXJlURzE7l
ClsjYVF5a+hja15MxqP5zEA933cjSXpEFYYUswYVAw7x/7Rsetl/e3Zyylhrn2De
617jqAZ7LK6ELNXe3Ik1V2ZmwYw6csJ0KVMnEfPhRLm2mKXYUlDpfw0xHdXNLlT7
uWOJzjHDppRyj1M2pM9tMERtg8WCqy5Kib+NpynZVMLQzryS9p+9t4bznViVoXPv
rpM9vEXSitfURlBrNjY71lgxz7HsgzO9RYxp3W7v75SHZYX9vMn3OjwbwV3+Sped
7Gnbg21IJxnWrmsvTj5wqQK6U2SZm9J2mEj6kIvLoLq0wiky1zXLfpNFExjuRqWr
slADLCt619hfFC0h9YO+VxEZxZkBaTn3/aKx1RwwYB10zpEH3ZT4z1gLf3RMeRYz
2cM8v0vgS+o4UsWBP3spngTGICudnZrz9ATIXNTvafZLmR87EsQg4sfCQ+lwxYW1
hd5JFXqKgLdQcRab7oueWhUJbrNfR2NxJUb/KdC/u0JEuQ+TIKsLPQheyKI5VfFU
GsPlPEmGjTaZpjZRYME4n33yF8R4ljqr0l92PeM/FsR4UflgAxvoJkslQAndpAyL
lMniqFaLyz682zzXdfHli90aeu2eyxIs6FrNfbYN0IE1hsTXbgCWBfxTkuem+pjS
/rE1/xI1nrhNccOBPie3MZeBEObAJnsfsOtEwp3YYKIwg3sQg2zgvlerSCkhzO3Y
+428cpEksUCz3+FSSMEPNPl3HucaRvhcJn4ztteqFFuc3VKT0fJrYHH3bHHMN2+O
FQzq7ffEYbOL8yGCLe0ORwZ4mOaqhtjEQGnOaZp5gxTjJrA4XAimgYK3FYylnTzX
JKSHx2pe+EsRZU7BES3kdQi/1aLnhv3CSzVT5f2tj24bBeSfU4qDIosIJMA/73ea
54wywL2UZGoFPWXsp6Ih+sedyYFUtTHVy4yijT9Wvl0j/X9fGN2lZiJ+TQLCIhww
/SWyN5yflklEubiEndZw5RMVldhP+mVE7OeHUOcVJwGr6u7XT0rPmpVqoC+C3sfC
A5QXEAgTO6yPW4TTMmJqGISNxivvPazwU0XPZr1fFZxnFrTzV9EkEby/5V+/qsBb
i0A9FNMSqMbPd3biZD3kFq00+O4GR8KFajm/S0qeAUpf1Qdsh7gg9eedWqgiRhei
W3R4YbjWNv/+1CytfTfqV2Jn/oaxlikZw7nnxPPILVhFeYAp35JGH7ph4uoKOohI
hI3w0SUFGWqdIWRQVFP1g4jKBwUW3ZGmE+GtZKWu9+mY0bLzJ4lV3194oauBP7Oa
5f8ueejA29xWwV2nSH5e6b7SjWeCZRBsjsdNCCcuhHrVU5LDBwYJ0TFWRPykmDJT
ptZQUsDxDKA/QKKlYUu4oD+6f3TJIZfAdovF0/JD6X59fDRdYYKkBUCJ7skpxWFi
oP+6pavs20aoL/hTLAHXtitxWACyee+4xE9UPQjXrXTL9glsH9kV3yh/YvPQpqGP
7xUW7pMCzL4jYWV+TZI9PWfoslqj70CJpPeuNZsqxexuJCMwREvRJuAN7lhjluUg
gsC1+wktP8tEOFGf9H5qGhI63XQCQx2qxBg+w+eNE2/bYWlvnVgcSMcCvwu7tDjR
T0T1LVi9AV6oz6cTYLhPwbDiKHk4cW92QsZ3uL97OSDbkC9C+Dk2f4kXe9G3II9L
aDqmaZhyq8eBXuEdb2/+THMrA0+vwdeyI+hpGkJEqPHQioO/2ro7Kh+eNRLOvZXT
+qdMQYDE3Wg6+3HdJSw0xLMlC9RVLr8YMlkXfgPNe1LhHk+vFE/4UIeKlfvl58DP
A5Dk2r5otc79DUBbAaumWCrlvCR0KgK7NYrrMgv/iH/0Pl6KG1pxU+FnE/D/g/i9
CkJVsnTSbmu2vNPKYkpDo2alB/o1NKZlmUbQeWA4BoCLvyMujA5vb3C4zUmSMMK2
x5lRbpXJBRBFz92E00rfnqkOlO3NiNzVlZ79Xze56+eB+3b9BR9aXw8/fEdNpBbc
oUMlKNtU/QGFrwLUSjQMYfuOezB2K5fgv07SheKI8DTy6/gLvZz0kcQhspb42n3i
nunlP9pxuMG9EE7RUTCVg5HegY5hiYJO7hZ1q1/OjqMa/90hkX6BHHiUI/bOlxzM
rpGERkvWccHKRM+ALb7+KL2ULYmT5Wc0W1TRl0VTGxj7re1tBSDXnBIvmbLbzDLo
yZo0Jr8VbjmuBcmV52j9Ddz2fybdmZrLre4JoA09PWKfOMHmw0EKYil1PbN4yqax
txv7cf6gWrYG4EfOccZKEDjGbV6FnsCPBPezCMbVH+kBhoSzQwCTTjTIIXBuA8pE
G5a0nfY1YqGdwFIvu28whVYLwef42/9YZyluPVWa59IOSpt/LapU7ZuU3JavkLw3
3vEITEn6KFJvmsZ2O7T0PtTpJfV4C0rEc4835mDIQACJq5bv2tSE2RYBhxUNJF/c
n9LxAncbXtnsf3HAtis0RyMxxn/1myir+P6FVc+YB1N7JSr+Rcn2ovTQkiotjJIv
ZHixP8s/pFaBZ2YhVJXqMnkYkKZjwzy7ShJquYqZdmBm1TiwW1jhvAM/CD4ek9qp
halCkG9HY8nbK4mVTdc5qPs/jYnrI1e2026tgzq7Q4hBWiwazHE8gsAaER3gYQiB
SkO9+6ldSrJEud9JHFGVKUgFDgdqj5F2j35wWVg0/k1b+oAV4UaF9/U1Rrepplp1
fvGsKVx7sZJ39fj+p+HsNzdFPVq9TkLPQyXzWZDchPcf4oBVUTsAOtsY/8LYPyFE
XxUHVEWjdBKL1VrXUDWpmxZtzy+K6y6R6htNR7ukfBGAR6CRv9XzUrNj+e46e3Zt
9sO0dP2bOdDSBWIflvOMS27Tt9wBi/zhuRV9u3O51vTjacgA/re3PFhV9yutYZoM
LcoH76vSXzZrJuHeSslISJlIonYDoixAip1rbz4fGcTevCmNMbYy5hsobhSui+qb
Kid0kuLSvNS3qP9QBz90ldQ1ZLvvlzNZF6h212eDg0pUsmLROjpWrkZicxpJW/Ck
CSXRu9Onf7guUdgw6isF5AOm4998bnuI4bi5R6HAxNM9zekJG8G+TXAAM2to2VMg
s7VkkYiHBd42+AQ9rvkCuntNiQFqnnf3h5JEdlCE/7W5Md9/oYzWLZ20OsFKFgRu
2cHkkjdQcGtQoA8XuDRlqmzjOCNU1gLNvxAQjn3eK79VrqrM68nCQsYWmlhDQ+HI
SCZhWryu/8KrCvTyxdRm2j65K/fH2T7iVR2TWeTV+bDe/wuTTd8CI/nAJPdTAfSw
olQfJQ18r1z6VE0IPs79oNEg02pwD8ubMVhlcvoBzAK1nXa0/4kygklP2rfHjM+l
jMr1zI43BbGjTNAC8UYt/JkduJFoyvwAI9RgTOqp1YAjQY2v2KFslFMU/2TmW5Xk
VXUAEDglsgKfjLlxz6R8g/R9ZA0MLj6l7ffM0qDBBHtbVNCSkR466toGRZryTXX2
I7IBUwcDpBZPrK9vN2W5WYwGKcoOYlUPB+Wf6bxJ2OkmYzEBAdTMOXeP8O+00Dn1
qSobqIMa5491+IRAJt8FcPdN2H3kVUoDuW/14XmIPNAldtPRQZWZ8hYl7hSuNsk5
3g8uVeeTABmvOc28UR0b17FwDebGbEDLcg0683VEIgssAcDAKFqh88/pKU5TTlnW
OWO4hDyqcox1aqrNU+j8p+fsT7Vaa7lk60JHvbrCIW8P9oaMsogaKezxHArjK6hT
qbdsPSw/SNECVTZOk8sNTUfGNDh6zncPMl9eiEDg0n5hsAWUtHZuMcTJibP9oOOm
9N5IwSh6y8ijWMmrIDWyh5f/r2wfpmbxBG4szTqcmDPydYJID5KLnTBfRhOhBMyY
cSeKQ7e/RkZE8qIgjO7yHsj/2oEBbQqJ3adK/xJBIUgZYHHGvELht3fgJMm+5Itz
jfTOssmt9ULxHFAG/A/he61wOgMZhZ5SllOXTK9I/FugRh+q+zwqvmvsBDKjcaV7
6gowU8VVXcoGQF/0hllP2dzkGvzxSlWQlza94SHwsz3IMO9VsIe249ipjVzft498
N2KjPzzqR+P4rUGTs3mhmnE/Bb13omoPtEGOeLkzOsRPKYqLuDNHovZ3xF1joBU2
AoVi6VS9EXOSlOQ2sxJGOIJPoo46ZUUGrLsXk6b8pG9HAw1ApjrnbcSQoLllNyj1
0Nfjyj19JxmkE297KlMNyt6yyyqRZ0aU0qKxcMpcbitlJU1/cik9oMKlBU+X5vjp
LM5452h7nkBynNNP8sdaHdJ0xOdRC6HjGwAYHt/cu+JwT6W2PKnYqMb7EGB8Vq2f
cAsMKqlX2iz+6JktsDnAccmYEFJvxeX49uEsKlTGQt3GDftQhEtqAWCJIct/f3qh
M315w5w/zkAKIxOdXUzE2X1QEfdeLTmELYzNTaR64LaPrNNPeeWbyyPadByKshMW
vsqnz99Uokm9eYl+i7BIuyVzzFQSUCnolQAsiBtKDzmYiREtqX+l6lwIJseET1M1
Abpvvv2scy0j4JgUR5EvigTSOcRkd5kCYi1dP3+KQsb3C67TKb6EWl4EWvLOZ28P
FFdWfNltqmXYXEADHFZ5nXkbho1QTakBYWNvafNetmX990XlHNjBtAkKBQDgaLLE
kgHTXDNjOHFLqXyAXMhCg8w2IzRKEgJUvpWrIjY26e0gELkNLUjktWGPJbu5AxK3
rlkkpgfnpSb8ihZRjs4Xk45rAV8l7UnkQgmmro520Ra3k28Uk0bHWvrhCCxlMeTc
xUNJVRKQzhUFplXoUWtwoBF8Uu0YsMDATEqPTtH9IgMxXIaoe/40AjRe15buivlZ
+xHP95/vm2LYZo1m1HsWWHkKcHPR5cJsp56/3esc0kNR7opWXZ7QHANmF6RJqLzp
+8JYAC/sFD05rY+YtacBFTH11T3DACFOlAZkbF4G7E06pc28mVGRqcXIvpMeY5VB
tLIMOP1JWuPaN7AU0kMU8udx7WfWEnfK9kJ8x0VjBfegXyuCYppUNRszM7qfIQWJ
3iGz849yZhVsXrINTqKItGH6FihrQQrcyQWAiKnHGOG/43vjBCFu4ANGfCqoAnft
ExuX+AQHTfx+BjMYDKCXmFSMSgVTeAsOokTkmBmN+kD44Me2KpQgYDKynYq22t+m
rJiqpVEX04cxXXTOJQnSErfjgA+Ra9eZRMtEodWwmcFSIRAXlqClkZyF0/IPPkn3
DeYu/hyGgE+UVES2iKnl0u0lNWb7CbxtxC67CPZxqbw/FGXagLbk7OnTIpv37vSJ
+T0MNBOGoDBGju7XjqaDWFkOoSb533hAJkynzM2XhEVFGZhn5bdK/55Ud5VnljDZ
/0FURjBa0NztGo5uPL/TneyQT7z8MdVInrkmoE4/Vgzzu34vgSfrduPaNlYn1UBv
I01vnXeJN3cMT+ffQZZHbRp2c/zia7pvB8DVxnxumd4k3rBxuXJvWVcK4Wb2hxRV
cEqdRTK7pzMjNMB+0Ii2UmQF88Xh0UXrpXxW6pg04QcX2q3zcFLYBFbRTnXKYAqA
0Av3I+DvG4mIzJeWaDt8lseJHzQ1gRT8xqlTWpEMyJUNWUbo2ubd6ldtWdRj1KXF
XpqaODgfHwQt34TrsUPxRIBBTlP/pLgmqqci3rlO4OY/fE14euN3SC/QrffxQJyL
j1LxWO759pFrMDn8PcES2KToDMX8q4UE3cDqefepbVmPbygL6XaUKTp7nFoAq2Lk
B2gXHrpRuQP9L+D8eWG+KXIKZOindDwwVl/W3YcrMBrGNxk732wTBwy/s0HM/0pX
6oIJoku4TE82HBXt6wqPLKhFd4r8eyziTMb2tCUIkEBqpaecEH+tC1hqZGXr73tx
yXYqWw0b+FJIgJ4eoEpga9SMC4ir4tbfSZkeTA0aadaeo00wZhC7FK7TjJkIMJok
UVLtgyZCrZMp0WqZUo9QfJ0vxsW5w0oBRwfB4bDAhm03YeQGAMftiQo6Ky4DC8la
T4rFOoo9bajjZ1Prx0Txp/SaWNiGVE4DLj/W/7iDLUYOYMYreMB5IZ6aOmQpGG4w
HYy+05a6InOTBqPt2+6l9buBn6Iw1Gg2rfik+xb/xBgn6M4BizOqwaGXQH352r/D
on6dRtWs5qGE3Uvo2wM8odhk0/k1GUhUeK/hqyUGbVp4E75ZdhLE8W9qeFOatY1a
fzKrX5XZewOqtJXyN95oflt7m3/iXv+mNP2mCeDNRM91eYSwotPX0S54MO+xSJ+p
DMg3UwC9Kp1RAAmPZTKTg/XsFNyzC3mugoUMLZywJkjrbCb2luiAcNTisUK1aOd4
HoYr5KDeViBXSGE8+3G7NHcwAzJOYeWP7L2sjhFyHj7KN98matDCREelU0ai2UMT
i5MTA3qq1VLo//qnfyFSeYSLzVxknGf+lCLx74vxI9sCBKZ95+/pq8KxcvapqVBy
8/50tXoLOHZcS884TGrOIINDXBhdfvlKVxjhg/B026AUuJBF/qBvSC99g6axE61s
DD07J22ZApb5X2J5hjck+3zAmBD/mhHXuxOmaTwOH7kHPfvg76YrO9JbPd9gVVRb
EdBv7jausVYOyLOpnbIj6ypDSkAXpJAaw2jYrhYuNWoWWribDX0nGqvUOnlYNW9B
UsBMWXw2xRuEsrjrPrk7H5mpWR3oC135dzJoECTvpt4oVeoSSYV8udbcY6EIzkh8
DjDSHLopRBApaR3MnaaQ7SQrH0LsUjjhFXcI4jAOrbvORTW9QRmdn1x0TU4XH1fn
gbhsQIss/RPknvLNosISvCU1GMC4rlwPbnZl/ifYvTKLaVKqEZlJXDFoHsh+5rcl
qvZwx+em79dFNAZmCWLmNlbMb+/YZfkJGNiPLtg6z2WfzsUaxLqjR3SMUpe0J9vb
CYfHzPCbvu4ALTMx6wHGYIy6oIsSA6zB2o7+AIwlIqC2nFzAXx1Ndt+MwmI1V8Pl
h4UKZpwLJxYbmjk/l4F82Uqa6zI7B7c2YKt/W6+HEeKwNaRVFlgEtwRTZKkz1ySJ
0MN4i9ElT7ChtgKQSiRkH7wviDamnl0x3dena3AWez2NorLmkZFL44guM7JMrKLf
bZeVEtd3dyV4jaMgav8tBcmsV73ErjqrioXPJOwQ5ozkE4NWa+KVcz0rl1p5D3WG
onJ8X6ONKyQ2wKORpz0VORRZJixIEUarTWQvfIBtBkXl5VYo5VnaVBLudEjHylBF
F4YEpT3yhrcWwejjCUmygWsyNpMsoUtd3Lt3vDZ4PFC3XrJJVFmTZdUp6GFWaQVM
SrKGq+JobgKqxgDS51W/PVcV6gjLa1z8vpsDAPdOZ2B3jUcR+zsziqkQonacINNP
l5RxzHLNKyzNLhGfVzdC0lEGabY7FD637CEIvGFwnEpm8BDVLp+EXXNoMvfd8LZ+
emNXHs9A6qk1/aLz2vHkDAPo4LZknAey+fYv8DpOI5jDDn1b21yUoEyFUAY1mvtn
TCpQhwV0zFzzxOpoyKh2IAjxXkwFvhhI3VMor7SLi1gOpZjI46imS4v8bMs7moBp
8vGCSP0i/iw9USpytCIPV38JIBUZ22qIk1TBD3ScJB705T8AzwDKsnVcTGOFrSJC
GY4BuGqr7zRNXl68bPWNTr8X+MXe2L7a8n+O5I3VRu18z0hmX0Oma2IyRXHbwGxv
XA0yevuxqmV5d592Mwx2U+OCxxpYEitxXsfarE6aQ4vg0sqto6MtO3hQJIaUvJ1e
azFOkwpe3RtiSj7jo/Cd6qtgi7+NrDCSs1rgEmwzWqFoils7vLEWWJyuBgLGaC/3
uqwBbDBVnX5aG30KsMbWp3kdzEb3ckvP/VxvaUpbuKWFzkkDPyC9U6YUzofencX+
034wqGp9Y0JkslbBslKcMOQ3Yx9pyK6FnRP4NIrjUD6oZDvXuBvMgpcKSDQt9YkP
SFX5xGGBkMre2k37H9X6HeY+scWzKwIwwB6YuQrgmeTtbh7gBQB5utb+85g7Vzdo
NoR37N8zAw7IKap1TK4MdRkVgS76VFyP+IrQ09CO20YPoPGisE/0KX+EwQ6m0eyy
oN2/zngQmm1ApSAr5dP66AdEniOiwPmJ3KgCF5tealiV0HfJw+E7QY6+hbZ5wzuZ
nwF/EhNuWdGAjmAOu4tbfhChQwfKI0ap2xvmzvTv1gd6bQ5UbtWWmDo7hmkLzf/v
hfykZeUxPc557U0a+LIBd/lHAKcQ3yrXmZIdbvarbj40YveObw6exGY1IxvmOeKf
T/38UKXg6T/riGwmiucVjype0746TFTxvMGISfzH6WzNTDhVRMGTPpK0G6OYC8OL
/YJQL60H58Sn4qwLxqZQDX2DOLjeOfoo68AIbBZK2+SYLfNBb5lr3CG9k4sJdd24
X60ecEuVkKcdwV5mtTUJks6oggi/N98nCEPTUi8t2s3Y8SvczQVYCGw++iPkeJBS
7gcZDlFG7Q5dHXmU/9n6SelujlRfBHf2WTlqk/8fEYXAFsmZQIwbgg+F/mYn3IZO
8n2/lwJdkmJge080YfMOjOmxFc2lTB3NN/6O0zz+ZUSpe1O1VRsU6IVd0sorcfjr
y1H30UnJZ5iEV/GYXB7DuvgOAaKjWPJO9WfnegPhAOeYIRJAhZzRUJrTv173o+OE
+S8L5ffnvS9WoMfN2e6adUjiVpR0YL/RudlDnFhBjEtUQUCYdLrV8iVS5SWJJj7l
iJbLEXP/t1r2sv1uiT1JnLuWPFYeWU1ekztnLgJ71cz5jeWsVc8+PdMNpqOTNr04
MaYBuDxTmkH3FfAPvVvMasGZkpGqFu4OLb+z2A+URmf6YnLptAKVCUcS5ebPnhyX
dJGoqkzXcAOl7vCkcz/1bILK39ATfJ5OB4lF3YgejbJAZngpJV2sC4EwCD4emi4U
fgOX/tbvuEw/aPXDFTsyECMFA51WY6zodv61C5IEvhPcapuu+6ICz3H5ddK/04ec
/cS5rd0Mbs2JIQ8hDN5COeIwHoaN86w4wO+XFMdgIS4vQHh0+TNUrqNkiSXwTtw7
bKHsO7kyDOAws+gyj/+CK/H8zlgJFCFIVl8by6kNGJifZ8+g0RRvxZDPHgWA4JBL
jMZnDE/Nffw3hoZpsoHuiLLkIWtlw6D5/swDunP+1XQr3RcuTWQHpnBe4cMNVwUf
ylkdoSpxieY/SzyOBJW5oa6ToR8Cpa24pFQPrKmKBUyN3FFGUosBO1syy4zFpqdz
kNBfqdjwgbLAh6rM20IK8TG1avdkJO7czzcRj5wuoTtTQOAULFdwgEAh828Xp2m7
rQ3b9dlyltCS2guNUhtcXRPWyYICz0bZXo60fWDLfy3BpgfkOZMg56yCc65n5X6M
eZIWEeV1D7Arc3BqEtVWxRCnYFmfUSAhOJcjBhfhEhOdloeJ4gQMuZIxVus/uwCy
qraqa5U1ePHCPHjbGdwwfvpqzjSQovcoVNze3j5VgjuhwOz17UgZmxO3Tokown10
Dr72Yzc0ey0oiOVlwV0Oxlqfpr+5DKcWLMF+XDCkGo3nX9gGOfx+mFMxUF34s63e
qIQ5ELpvKHWLvSkOIn7fw6ad7F+2dzabrJN7QR0gkbBvnbV6jIcvaeNaiuAeXcs/
2C9tD9qrEsngMA7do5Jqls/XT3jCZ+g2MKYQVGn78XaZac64WtLENUC28mHcebQM
9+N49ZndRqhEtyEvDuZMDea6p2209ZJPeZwIXSJ2llskhZQxjnDmNBwxiYR6h8nD
/YBA0GOzK2nAIH5a0pwKWG6RAH8hBOvSUuy1vnUQEvAIAGPUYhPlHirXBsD6G+Y1
C5ZZEmgUdcBbwZxs6u/x9Nm95sGrwxNmkwHlyboZcBoQteDg9oP//dTcC221Ez93
XkJzS3ygimAp+nQqNou2T0PrZKva5YRhkGqPrmnO6PduN562JEmsGbHva+28Sz/k
5xLmEW/j5RE7HDoGUQhQS/QVABEieVDvFtBjCE88CyHfITyuSjehf+Bp6cQ7CdTg
YsHO1k0Wnv9Yt4YObmgKOApXJrMsxXlZE8r0L7NB0Jwt4/GtbkQYBxIoJRFv9U52
pQpAsT3fnISsnbqmjWisyF4F/23YBebHJ/z5jGYe7b94N7uacFkTl8KFDKv6+w2P
Gy7XtE4vcCEidpuUk+ozZwA2dSW69WSSjcgtcWmzjsbAohDQsXb3awajg6dU9r6e
2v6XXskjhvI5M3iFQ28yyBnoGf3NcwF7xCkM8fP0MD1Cwa3aECqUrFQFwTbGZnRs
X7KNVBXl3nYwpZcnl2/je/F846cfTXhahABhhVBhtEYpNPJIf/478590z6HYsmbL
RjrCRVaVCvYsskaz2vgNW730TGnAknp3q7KQfGtRvRDGLqGMgcT7trfxWIqtvoDN
XAu3R/cJdI5QISciQ86FyenJVcsgK+vWZIg8nlX+l5HubA+uHAS9BNnUMHBtABIR
bTFEqcYgbHWNcRb8MI/V3pOThDCCQYMkQeRFQMFdU7/dIG15f1243UyA4e7Z49sb
AadhEqRlTsrjHB8EXIDdR96Ht/nOrnn1oWh/YMJSsIv50kT+gxuh2PAPhRpyPbPo
s99QLROoT3EM1llBt911w64OonkINa/cjEIZgbTvPUcuAL/8O6bkruLFeSRkKvA/
5E0l7cjavILwmephJEvomcJZmOh2p0VWqiJ5jdqSNIx1tAJuKag4b495tGdreRAb
s2XTgVR4U9BTpmuzOqUNrEkigxnHkUjAB5jxHE0r6Ng68eiZLdkE3PR34gBugCHZ
e5HiMBWC7gXnIDHTox79yU+LcLUKIjTTOg6yG2zz/frCUsjGv9JWIqYq+sNLdJAE
6dwzqUj2sHkmUq/cYvQCALwuM1K8+q3QENPvr1PvL3ZuhEb6tKQ9umJcACX1DeiG
Y+szkEfPdVXOiynegQkRFuXtPn2sd7sQNdJ0yWsJ88MAsT4D/iU+YTGUp7F3c/mm
noRvvnT1syRpUAb3Nrumony+EQ9xLdbkuGKk04MTfdzOHbdasSiO1hQgi5dGmkO4
j52+I60MonRNAWyvMNfcTTqpv3zJGba9vKVnNkFyBBCw9thcvQZan6gHvmCpHGO0
Fu0lLYaI2Iy8zelJcpKSNEKyAQcQgIksUgsQM1SkIgoZOjqCJ3K4NDKPTT39HGSJ
vnnV8TW5yE1AsjPO8MCKP8E+fmzWCuUOgTJREFCMXmqQHurOkTM6M74dG/q/DSX3
yVySql9QxYGxrKkAPWXqsikLYtqH5tlMFA+Ff28ftspmnUlsFBD9gdhxGVekpIvU
vOnZNvNzgrNl26ew434NyjlwBMnZsMMulblC6W2VhRAWdQ+Djbre0//bhu4G7yKH
JRjjbr77QRCMID264Om7oMxMuhJyh6ksRmVo7O/W5cDzcFthHdk1p0Yzq7SURUyi
bwYUI1RiMjfE7FI/MDuR+cexebxbxl4JqZV0KGiGazvNyXfff8gzcb2xR74Txw9i
VvTCKujUtnDCnwKbGEN3uF+iMR21DRR92FYXmAmAx0GGx8Pip914oWnNDsviyv+Q
7axA+nUmzgTgXozuD65v0HBHtkQGfQQZiy5+8OHZhkRFL4zr96hewFLu0GdYal4t
1Xusr0D3Ae9UZ89KJK7lbyj9PmB23wnz55jI+uPNYWASpeYHmeK869z5oSCSsh/1
KIRTjjbtPNbAlniwWx1s2SOcxwTMEW6i+bztrebgzC0DyoGk4mlhAAmvh3F30QVO
tME57dXzu+CAIFoA99q0pwsjzxmhYidalNk9VDjhNbaL2mKNow3Hspjc9UypRVm8
OLUlP4LtWgfkuXCXZiRAyx7/SAv8zRlf2Rm59oJC70eQdr7SSLGmrmncX5z4z/Rd
9wT54fzbzQ4OpJ3j3DZLQMeW8P3+RWB7nl5qNMDYKZOrBCqSHxUmSFewSNZFT5qN
v/HWZatYV0KsaHpo8kvYfAmIooeSFBQ7zjQyB8JifvD7k0FPqbgnuQ6hSpqZIif4
Q1C/r4WqIzjJD/nLd8A0ApN+a7XYU0pFGmXXJhCUm4nPvtCzFbj0cVyz452+44x5
qhEQ+nn3AA7VeqFo2BwZRoErsx1ZDQUUkFlzQBNkNcL6/B0vflQC69UfpnmGKzv6
cmtujagjlBm9yq5iWR4Tgyz2p6bzCuHqtGUKzfqxWOZejTq02jbpOefj0XpvruaF
ipysuNB1ChLdsKTaRlT+qLmR6DqlUJTwJ6Xs7qZ3NmxkuwlM3xNvmwMj9t1VWwbc
kjmJlE4aZp6+UPr0ngie8gNmxvKF4x3gocE7LD1vTTjgsgJD8qozizM57wuxwIbB
s48vLpEtZxolB7p+/68n0Wf7Nsemc5xX2SyuIz0aAD1KAco5vzM22C+EuRE+Uvby
qbAsqlDN6uuzKmexOc9VN8lp1fGMtcSg8H2c14EB6Qmaicd40WQ29WC5rgpS5BRd
qD+IsOwM7KYTZ/IQvKYia2y6Voo+j+v4JXAEPnPUAD5HPq9cWlYAI15HkWSkEYDb
aoMzo0Lk7qvSMVov520Q2mEmijqkRq54j083+ttoMp83BXsJEkNQz0ga/OkF1cL5
BoXyFOtpdbHiiE3i2uGgPJ6Uon52xLie+jZrw2HXG7G14frI7/VltGiFwDAcW5+h
lGrYdAVglGO7fYORmHlOPW8CLiBe+/aUa7cKj0fHTA3A4SuO5VAm83kMAzQGt7Eo
NVGF9HcDkoUNB5wrw9DUlbpBmstxjebIMzSU8F/96X/Gjti6djtQGHRHnNi0/JKc
VziomDe2INoAzitWd2ALBaeMlPHkaqvar46jmDKKnYYVoYS8SoB5GdMlQ4GZ78L9
PrkxTk51b5RPkjdJrDEFy9xbprtcyvyM9DQ8sWv0PrTsHhLadN+q7z8AZJiYt7UW
q2pAqb/SumGks7SWLpvmTII5tmLEWge9Hoy26HJK9CHu+9MoUDQLkEpEsIeHQZPx
FVHsXky9M3e8GcUtasAHXuAqN2RtMBaocVkT7+ok9J0hU5KZ8MqlJdTv+3h12Z7o
DOG0j0id3WG22QQPh3HiHBQK0dI6UCDu5NcW85aJuJmnHznj1ZiiZAX0zskEPHMx
fP/4N7hF40rE1uBwAFZrWvfU0DxcDsCr1iFDgqYgPwD55Rk01VmnV3N3siM6IoBQ
tsrkpSLfYJt8SLLOeDB5+nLkVlfK73rx1p1/pmEBZtnmVYalfTW7A1a/dV6egQd1
XDzPNi7AG0nbodlhpFenRjbYdMjKTxzfu69+VAJABRvgne8I/oHW1eix9VkqnSlF
ojnp39RNq64kEViEtFTtbw+ETcxxuELUJbRW+O7OOFUdlNbuCaVo7sM+8Z2U25kU
uKHMtxFlgdwL7wnVlfu5IbLdJibL/OswdozcFmKmLgdo4vBjwc1mU5tXuMpJnQw+
jAcFannBUyfADAwLB0gzFtF8avOtZgjY2RYoEc2emt5EyhX0GvImvRXPBrbAc4Ss
lCrTwEvIWyifserOVySMyctX2G9S22ZddT+VqTbw3wzo9HgqBlK7guFUu4Fyx23D
28P+dGKc87SdfXNM8YXOfUmwb1SgWvSDIuNCuXcSJQ0jm7ziHZyYn+XtczStMtuv
HjuBF1BdObAiHqwze5yfroEVGwCFI/P4jOVadroCeHhl792uOXytxbBhAEEuvCXR
u+8XgtiTSUn1BGJBRvcxw85SaOnvWGO34xrAZv7Vggz8OsUhBS9SH8M3VTm2VUyS
wm3/nJqkYilBCs6HT5P4veNFn8u3iLPDZE5gjY9Hdgahq9Hf0iYuxUt6EScMwCYV
G2Aaj59SyYhf2owPmeCbJvR8rfLdbvjrl+5C1rLuMP6EtmQSrXXGa79CaFY5v/VW
bdLwA0TwRevmNOEro9QPxj0YvLzt1hKT/U2k9HAHiF5znU5gGy9369zp7UeVoBOC
sjPCDVUHffVDEBKk+AUQMp99zJ998KAVOClNpYIIj2FRLwqo/+rSjDAZhdqcACi6
Tqj7wC9OEuE4wAi30T+Lm7rvs1QIxTIgb2VvEq0CsRR3U8hKy0eqZaH9JSuitpzn
JkmiTZLwHzJ++/yhGTDydXrFIXLf4/yCdWzV9ylPx19ibJCPuv46ORRN5vQTo93f
q6bj+er6Ee3vxIsyy4CHM7QCr4HuJ/1M1MaIar/0UiSp3vg11XX2EBgCGY5aMo3m
lesqaGY6MyEW10D0agkiU1xLy44CmEb1GTjOBZnH9FByhWo3JkO9z4sx8osG5OZn
SM5iu5dyeH/hj3i3PXO38NIIve9VzGIZ2hwkqpEMHv25y1pXZZ1wORmVSjSN+Ajz
pMEyJi6lUsmIScPYkPOlX7IW7htovelyLxMZfpxWABSDI6vEbiB3ltCHoQffmwp2
Dc79SYy9y8b0yd0fDNPhHK07mN3UqlrnryjyVFXQWPtY5nMrleUzWpHtFJB6oQTY
U+RRQHVBJlGBDMOSqB7gBjeDqQJdcY/W1uPS3N9uw/Nm0HjiLX2ag/hmWeThv+/E
BYpxXo9F4Dxc/XjjMEyd8ZOe5NBB5529de98g7a5KmSs20hqS8c7r57g5eJs9a7Y
pCHIkdmNEgDXWsfuLdMUBCqK4djFHw4UjkCwmQh0jfhH4m2lTIRXTif85EGO8fv0
ccLnPW7Rq3EtwKN01nM+kbS0Oh4OmkkqIuhQXgTEcO48ZHa93Azw/iR4Cjkb/OUD
lFADe9wkQX0NxW+50EN4mX7b2FfNtzbq3o1sa4ozMtSDerqBilZPuYeHwpAlKZZq
wZayHoiiPiMkwQBa/BMG5bviEJOsNRhhgunrYy8E5zhVWgd19XFeBMEzhiZkT98T
ISt+cIIoSW12zJiTTMOgBH+Es+KKsaHkBY0FIDS+uRxNrXMmSZOB7DN1BIFAd4B1
caTVRW/YPnolH1jevd9BSEerC58t67K9d2zpXwIkCSHNPXIidFydwMgGXFK0W8+m
RlaIy/MLrkzbBKnriWxd5cJoM3SatERuCCmzraZHb+on8GmhutA8SNeMivJ0KZdg
NO9DWdJrvyIO7Db49V9+E1hkdoqGObf3Dt8fVjHAf3OHjLqUqXQ0J+SAXaIlS744
sQZnlIQn/g+BgLftDvOZDOXQKJtokjB2RCNAFhr0Nr+1pLYyzlUHtc/msxmaY7JF
NnVawZJHvvwKClPzrgVVu2wLyk+sqxwql2GFcL88OJvFbCbDS6wArdX5UPYD3iLy
/rrL0TE+VNGnqYnOO2XlpM9GH8NtEZEV3xM5BXI/4OU4gj8/0av9LXRmexiPjY2l
RPjk/g6vEKjmy94eVpmQdW8S0p5WD92HsC2GNf/iop5ueXMDagBfUYn8ZiJ+fObj
CsaRxqzPXR9U8z1VpIihsiEUCUgU+IvvRk48qt2R2nQXzjjI/bQSgtjQqdp2jiW5
u4ylqbNOah7WyMZMef1aiYc8AmFUixVBCOoKo6AvZWQcWwRRgrJb94vFDowP6iV1
PcIuSAXAuTB19nhoyBkAVQ3dc2WEvK3tJCvEeCciicS1pNPyI+I/nK2CozSZ1EP4
DqvgUNtx5Ope5DQ7HvOLbwbyNDS0QwDGwqUjo9dHpX91RpQTY3tTgbIHTz8Cksua
0IhXtaCFeVQZQNCvzQ+mkr1rjRNaUZDcRR1SJNlBfbfmLKRIxp3i0bWcNHf5TnKm
BGFEslyrPOJAso1KOkPv5F6hUCS7HdNdgbdgp/D+kl5ByRQLd220FVNqVNtDJbPn
rmVGPW8x1eHUusOD5+WJn0zwGyhseVIXpeE6Eqp+DzD4MPq2kgBtn0OHnjXnbEzk
D4Lg4iwyGOoY9lteYzBqCHiivqDNpRkSJLOjcOFP246goTIp/03vSvWVNgATKYr8
/gaJFvMTC9sVvUQbf9mqXyhXs7WaG95QzYneqfjjcWGjvVqZuy4HPb3BKXk3EvOx
yD86+fgADG3Ipn5KxVqm3GDd526BseSzGtyfeDbEYtbbSzev3Rbh2BwVHAtA9KRp
mWQ6Gk2PXg7NqgwqMwgDaIGf95/FCLajosXv+MIrjzOwvXFV1Q2E31AGIprAoZbN
8sYqxUQQboOHWYN0kNVMQGTni3h3iTozCT6GRzO17OxVmVCWhUXatnewhhvW1wvP
awRbj/4O7m85Vi5eTHmVbsDAe2zGDWim2R1AGi2xpC4sxtOZuK9E9QmBDpTzgVSl
pAYSOtyfJMJvL7Vp+4nf9gJTaQq8sbT0DPdBJyw1tQ9HShKc+PjoIyX9HH3PNWs0
lCefc73vFH9kIaolb4092ZeTTdhIdeFqjHYeTIbXBvEJglJ/6EJMyXouFCV6iibn
auaitn8nRSgciz2CBYhMniWtg406RFhLeQhzzYZfulHO5rg7GrsjyPUgm6WsWO4e
KUwtT+f/+Uq1AnImysyv4OE0vWWBGbnXeiauyayYad5IjT/Y4iGpXvbrPGpYsYm6
z8YhEbQC1W6ruK7AZ9VfKcis+Xj0PRlPJWsxZ4yKskFpOpVcbj2zEbmU1qrCm1IC
EArP3gNyIBh1T/OhK7K1zLHJbRMw9qjENweCEySAZHd8BFRybJha0odYBrFcgp3m
G8hOJjqekV4wnRqllbZ32KI/y80G0iQh+1xSVfLTldW99Q7gkJvZUt9+VfpM1Afo
qKNGlV4ZefpDisI7NXu4DJWhFztpB0FULMDRSN25mdJSfQCoISrFBB0pgTnmj3dT
d6SLjVQXW40cWH6O8L+mgx4S7vKJ3SRkR5/jZ3M+BEepL46s/RtYGsvS3WTrtIOZ
KPYR6qQ3e09l4Y97ulYYmHQxwI94mEws7oVRlo3Mbti8w/ed9i/YRnII7POMU3pm
5My8LT2RA+LMmP+uaMM1KOXH/wfv2xFQuOrYlbHJz7/9ac9wI24de220iSPHWEdW
fPjbLghFSLZMyD6AdeVdChpitnzFJ9Iv12YAs9+ce/WiB0np1wmASTJD1N1gBQL9
LKaBRlwWz+VhOd0iSFGUzStP5sDfloBlsAe6I41LSoa/W43b2RnKW91CtGGLvXnx
LjsHCQxTik2pPfSkOMP4eAQRlRAKsERP6kWN1K9uAhO7Wd0A/VP2MkiAHjKb4pN0
76hRQDuZcs1a40E2a8WtixB3/5yN8b2jobqoabT9Y+CplLhQ9ApjPeABw98iSugE
h936rn74LZw4d4trOlA/HzDYXQ9yMW6XhrcZ8evBwmoH8tDtMVrqxR0yEedctO7E
onh/J3fbkpMP4JcmKduxrK29OgOGyburiKLOwtszuZqHqbcrIa4/zXTRZxLq3dnI
4UL4b/J/If74LKhBtsfkL3Ca8kCV8Joy2RvBvieXCKNspwBcvZuGVnT/gbfFkl2L
hCdSPsUsu5wpXeG8GmzN8leAiYe6FernCIFv+6h78jA1roqWnDk1bel2Bzz4V/Pj
aA9MIygaQPoEHOtbnR3uRZVPW1C4ccSo7Q5lJTzBeaM4U25p+snzJaCesby1F6JS
F1D2KhwSrwqiRPCL8ToEmo7U565BZtGgvfM21OXgWHbqlQVc63sDgC+eM/TJTG9z
OAJRbj5lPeJL7lHdmsce5LUnJcbfRw3p/fD/K/Ll5PfYxNqEmtYMWG6Ij7v5u8DH
mXgomxrPegZ2C/sZkI/y/vaO+Yr/zzfwMr4lk2JhxMs8fAKCHo5koq+fTacvRZhu
QXcgTDfYwXvX1MD8ikiLgyLzJxhb4Q6EsrqRwXnq3hjkGLcuufkSY/bIsSproOUy
x2N6/njUSrqFBZKWVtx2/WWbvKbAyZH3xqVonjTTLXApCsiZoF/NNkGF9f4zg4p3
NB/y0P0KhIajXAHIljfTVxYzz0aRQfZri1HUeRX1XCzskXNCTbjql9LT2GNBHTr/
X8UY4XMJ8fJtM5o7x0ORh/b/EIQf9O/Ut5c0Nw5d3+43FGB7O/nL3C8TUgj7J1ni
+33FG/eCO4jG+3UBlQSzEFS+qAGohQdu73lTkt2JiZXwQdlgElNRFKYAdIOnPZ1d
k39oPw+MzKEphDMoyvSGlcR3UQxe/0Dbl9aaoj8IlLcNEdrfSgfUB3lsyW2GpkUF
x31OjwFEHoQbHeLzeeW/o2f/eHOPxaB8wQvTS/y8VosULx3n1RjKIU0zX9LzMzq1
AUIUqmptTIoyc655MFhHMGPSbR9K1YY67Cn/WiNTwPhRVDlp5eNTQESgogyU03tS
v78ExRXmURHb0CtcuuIOoFrieoSsrd2MN4lDyMa2djiCdriB3ntO2AYWI6hUEnB+
Rz30asW5cWXpeVOGq6PWBb0BPqhMsjWVwuAKjg0/L9LnJECELLNycQnmcjNjfTjU
b7omcnfQepo6TKuPaTG7yZyEfQeAZ+WT+f7iIxKBtJisLhd7/QG2Sog32eUmnppG
CS0cKImZt3B6S61g1/xqiSMwjGBxsdkrCS7Qq+xaOHV7UZlYmyvVGnPSe0MXfEHA
TLUtEwyu0dojg7EFJTkXYS76cr0dvvf6SD+jtzPvKtu7iJgkThswo7cyaZ8hrN4y
9NB7a+7E6P9SQGrIupVUleDGGY3kiSmFtofhtxsUMus6Ja2+vL/VXzmkiDUlH9HK
fvoJpjWqFH8VO9FhijhPjcTXz6ImsdWExGh3dJ59GlohgY8fvGaY45hiJnhyniwM
yFPMtE+g4T9ZRew/+mma2b9CoVfOCMc2vvs/excEYQIGd55ugmK8gGGt7T4y1t7i
BDCKiaZI+glbkODfVYLSxeAkpefmLr1gTKxzBoYAgafCDBs8c/StzfblJBYDUL6P
7nJAuM1KLZE9no93TRz+M0AfsKjUtKX3Y3gZ6tBehn6zSoctLvqQ6EurK0uDaT0R
kDYZ/iR++cEWWhRoc9lJlOroZVnuFLdOhIkcpKFB8I/XdxbbxSLbT/mwtoIqf/k4
AeVgzYLYqkFXYe3hyIyif6xrtX7DE7gUxsbvGWSJo+g3s8Almm/OGBYZnxW7NXCU
YZ45kM0QeRR3PEnNvYWvxYLKudgtkc1uB8+NMspT2T1JlloW1ECcnGLG8vvOptgI
eY6luMZiszVPhzkz0oCEfDYWxAPSjjv6ZL8G2I4JdwLX+FL7u0/Px5kdH9oOKvGs
1G3afUyyVsH6Xejc9TtUH028A99iBrTXFwHP9cUdmY53iAVnsMYOuUk72+mwOKfU
bRi7TCg2vG40iVrslUQkNpWB8vG8PF6bmoPEIs4h/+VNF7xV3eWrtm77lS8ZVWKZ
WXw/t9OCHBZMIzcLuDW6aFX4ySoRdoW+0CqWZrc5At6LRAlXgXvQ5svL+r+A1o2O
LIo5S15JIkYVGxr7nmBShqfc3dDh8cQtmQ/iuf9jnk6FnA+vWjrP/8stEP1+RhUz
ycQGW2QFcufZyOPpQkGpRa9Uwq9a2oaiaRA8dPAJ0PaNlfoIKwBLaFLzl55pKZLh
8/bgZogXRsh2vL6Od2pD6u7E8El43p99VhEK3VUO7iOjei/+brQo0TM0cw3V1q67
RmfCpC1uPM0G2yk/YrfCThUfL7CZ0s4DraFSllo4pec9bqW23v4ochwSG0ACUqDm
dbGfZJrlgqwm/Qrnmm6hWh5X0G548RDg/oHtwI5abnMEE+gjYjxhYc3sobiF4NyA
xw/M2krSCNkA4E6PxxUxEPnRq79GoRs5TON99NuTjGH1n5uwWhrRDoVyR6cb8Wuo
3USGxp3/gILUqKH3+UXOW/kJVd1rrOiVnCinhfwGE2aiPUp7VJMW6BNGBXUhs29u
vylMPHkQT1svcXAOz6+vJwjfedd9vm/mzOIz3w3/RxFlRflGlaWfXaP5Q8yKhmyV
mbnUCWj2RS3X9t4yRNG/b0RA2ldReaLicSDkxw+XkmkVOvTCTiB6MKjJuOHCze2G
2aGsI0o40a+qtaHfwPuEjOxeXWZAHw7maCMGi3sE1j/WtVTtldVyUn2OSp8HMgfQ
SiPuPCK7i8/RO5D/ImpL01JMwb1hRkqeusRulYM+vgu3neKsgdoZgjABGuyqH3Tt
AWguz8hr++BQjsnIe25mlGizTEWOhk2YokO1iPD6QCze2xG//A9Pz7FA+3TVAXgu
LrZJ1jS2iSpUlLF4pPhl3+rrw0QHio9f5q9tPVamE7X2AsX2q/iyVq14p/MrOhmN
BuHib8OtPLSkwYAAZnElO8P5oGiF4qa4qzBPUFx/JrG4bBqdIGJrhC1czifUh7Z2
R0x9zLpfwJWKI0dKUfbaHiV5RpsKzG/+J7PluYVVCR4FxqNmLiXYfd2DE6cKJ3vO
RfHFzurNuLlglXFXH4L+zWVHacVbcXt9wjXnpGNBVcPUHigKJEie0UZj6sibkQbM
wqj2kTvvZXazvicjD6swoL/wsZdLmOycFxA0hWtgHPqZ47qLNE418sb3BxeNxmX4
CfMbeGypzN+v73ZjrgR4r/4uS9Pl5oQyjsnTashujeOrNasWuZ+GX/M0q7njmXpB
luCsKjD5KlIHqQvoLVhhwM1v+tudOpEUZEHI5uA8IuLg1QGLh2xbd6EFnqzK9hI2
biPI76dXsPaI3nP31SpaO48mr8GtrcSwNih+BrPIf6rBq0gEIJOwBrWPXeNHikzR
dekZ4BQP4Y4b1YrwJM4XNYarA/jTuX/+3+UtpWz4oj9TtV/mBF41EvX0j1kw2c55
fsbJSTfyInPyhPgsMfCBIOC9dOCQgEGPFBpjHlTu2ymuSYLKlPiVOAJT+bXgsT/b
8LhgnSikt1beqJyV+OK4rwLp8fKLpNTEbDrkN7PH+5u6PJ5X7pcNWthmRkVApok9
yvv9T+HXlZwoqL9cgQeCCpbk2mcpfcrt4MVLpghjb8D4dgXQs50EBlXWp77r/ePN
RptIYnQnH6jfDd92wqmFe5OydaChvB2FPafuh2dFiBYSHx8W7ZjsqDfDcMsMEHOs
O0rYgXSTSZ09y8ctDA0XU27dGMPFQwjrWUD7vHD9DajpwLu/PaAE6Hok1dQrqOIm
mPKU83odEKreYBjeRSORAchRkUPfd5J2RK1/icIr75gM6DgNPV9iwi74wXzGSOlo
IXcDSlL6DsQgx0YgROomjTG3gMK+Wqj3+s8jOlj9RakfvrB40uZqo+HHJcqN5cTN
iU6r7QanAtteWC8Z2odTfG9HRyZC0htTiTRDdhjLw2m3PENRm3xIp3AAW4/ghDoC
vcnhUMwm6AElDbhorcszBXE7uhxwo0ZxJFXeVDCHL40UqOqxTMEC+CK5KX++Ix/y
+Ix5hd6AY0XD1z9WxGV3ZaUc4FSfGnr/J1c88TdRD5I2bZGOPrxgyFT9vTmrNhU7
PNJRt2oSts84qiDGVTNBznJxOtaj1fUj12U6Lo5ytbJi0vyzI5al8i8I+m0+xOQh
emjTScdEnM1/vJEkJ3YgnXOyiWgd3sFzd1ZHBFO7FBiOCqKKo2+L9pk11O4g6Pax
AEKIgOv7UrMWJCEVTGEQGAOcehYiw1QSd1im3K2CqYEv9MZk41s7NN2xPMr7C573
fCSdcoCg6vlNt0gJjHZ59q5KAhpx7lBs9EmkR2CTcIr11c0Rds3yITeb8NW8Mbtf
pgubTD8Rr6Oa522fRL/EjPohVizUAaiiLGbvUbfQ8nn8KE1Q33RzXfuqFBLWydBc
dltxlLbRV+UttLFK0y77JuoqFW4GVLU3YDbNRJ3hJHhUdnQpJGcFuc06AQ+fdyO/
88EttWF2NEXteLY6mwFVi5I/msDNxOR5QkajlO5mnc0cfz7wSfn//f8h8RrYS0lG
bW/YCLaBhjd7JbV6PRajmZGZKmg0Zj76RkoVeoLuNFoaQWin0RGMyJ4EnSYkM8Th
stvHZFStDJuN2sNF+ipPVwTnyn6VmRxjaXIFPZIZUg5Z+k55iIHcwEKyu1sztke/
A/TQZOCtF374oUFqxUu1bh4Lcy+0HFNoxdVXWA0109Q3o8psvMhWt8ecMqY8EA6c
7PNgNVCSRDgjawstHiqmWrCwGwzwmZ7CUBtpeYvDx8nw9F5zptHi7qKbeLz6mQqT
cO97jvCpy91HX3D1/kfsxUIR4hVRMxIyAwGBS1CJg9vK6Lotg6EHhQD/QAvdGFiG
lrCntqhViGHnhJnzrUD8g7sHLo4vgz4kfvKecocf3aIudDj0Bl9FCu/DO5SCZmqg
Hw4yeA8CiRs+WYhQe8iKEbjzLPmT44EBZJSNgRdaukvQIQUx+Jr5LuJtn4Rkl8Am
a3QpdD04HOJlD5aI2/VtbPdymHQqOBfbPNEwaUp0FQR+dtlTgNGXbzv2tfD237Sx
UPkEesW70viIPSoNr6MGvUIwX9GE/Zx5NowbifezvFklsiIKEaWlrUewBUkmQ96j
SoX6Zb79UGA6dncvqyL/JK7VR0SSjzv2gDzhahHuFPl81bsKJX34uoblTmEwAsIj
66Oyx+zxAUxCfzi71iMsY4lUcyNnna0+gD+XBLUTcNgbrz42W+np0j/4Lt+vH0+1
cEkpAuCwQaCeSlEXaW0+7rosJMjI73djYvdSnLCckQXoqUEPoDOV9iD5EvLjB1LF
CJezrR60OtHL/jj0klp6fCnXDc2KdeBsoIq3nI/UecABcDedYY+vq3J1Jmld1AfH
Val4gUkls17K2fbxFOMFtybxG09jJc9d8vGnM3gadLdVFQfIlG9JGHsTEhjjCYbQ
A6dl8v8wrqUCA2hx8YP4gOxm162lXoVWfwaGydPHPTPc0wdPgdmAMsw1u+T05s31
hrxbEcSJg+QHU3X/1qRDv4IA1DYLrvaYU7mY1abqQFaPJwY6VSVSWJjVO22z/EXE
kiIfL4XAAralfidf3dVGR5aTE3YRZCvePh5Cs7VnTgJlFqvR2GWN2ApXxWIlxaus
qEP9QyJ+JPzMfak4j489LIwERa+YLdrXoYMsxfh4IHpoYaBcjrtGtFIQVfw2yoZw
RxH5xZawYwZ+TDugv6qZwsNg9a+Mhj6rdmpTBZ+82Am1P4EW9lTGTbKLSfRCSDOA
Msh/qEti8DOkR1g3ADtjIgEciFsqcIxBi4U8LazllVPQTumXwcxijiwDRNUiWlue
05bv5o6dcKoFkeg+4cYWyhwzYep1kpqVpiUI40gzg6eauPFk6zLvs1e0zRcNHtA6
ANwXge3mZa0jHsPmZR3+ywflz+g8t/BDK5J2E+/caazvaHEBQSFS/N3MCASLoFYD
HoweRkBHDgIDKcy5yp3aWOj1pCukZH0u1JO6UlBA7Yb8a+8irv6UV0t1E/BzI3ks
/KL+LlQx6VsiBkbAqeVZZS8rsdyKEc8Zs2IusAySEOTiYyt9rzOGw2GiMKqm+4wJ
AdLuxFxqiKHRSUYcKmILzi5cGHN5dyVrTuP1k1z0boJbcewOdeAhvDSqlC48aB/E
V0lkMBa/BSgX4Fy9YjYWeNEu5VfSjO0vkt3lFwibPLR+RFkseJe7MpvJGGhrSlO+
Msu52FdNLJCtK+M4U3A5biXQR4wlEilOOTykMpviPuVe/fG1xURgIaJHnfnvz3hi
aNFBQi6ICJT5LXLNuZbG688tjPxg6V9OXdDnS9JSv6pB/oSV/VpKu6M4gChCcFy2
Xxry4eAweB69Ur//ukteC5E8H1COfOyM9DNBymPx2NWJCBLfelpMtyQfdkoXN7N5
pDje+HnH+hm7m5mHYzjmcZnq788yHrJQo3MhxT5TKHh0Ifcg+4ZS3IthKfAlhaiJ
aLT/j7cUtn6rDofedE/qGAfSr3SODXN0vMkize/oqSuPJyIokwxO2wvpHeD5CfF9
zlPEh8QM10rhaeQvHaPQ2Jl1p/nfrq8eQsj7lwWqIZoZFTyG2iWOvbEM8hwrVpOQ
T6/ivvRV9NSb5b0gZ4jrGywaUXbQFfhH6mCe8uf0820bjJqjNkdEB9jaXPqkIq7S
12hI24ZmiYK2sYP8il/VDa2fyy6/VsjO5uU1wi/22c/NYJushlLm+8tHRKEho+L2
Ij7rY7cgWPfKqWFegKzOcqWHN+vRKdfvW/9vtgJ3p7neKiPChYnjJSPMQIeZzjJ3
LlpzKHFlISmSpHbQPqD7l95KAfj4YNYh4kx5vvgvQ6B9JX2v4HbfomxcGRtka5/E
sxOeEV2O/HDKFQExZVfRPWGglWJA7kDC+LnHwM47+tCKDVrN9BMBJkayFR0Jg5Zl
7L9JmtyT4fhcRs2nuvlhr91qbVNhIm09GWb4Xd5GaMxyJifmYbd6S4BDaZ0snmaR
o1rSA6lg1evrpB+gmN9NRPC1kknAWlJUkH8XpXYjw7UZPz7nivk9YgUhXhPWYUXi
hNR1L+LQSg5EUr3jHqQ3WlwwfbEb0VSg+6tN84351W6n4UTJmEZ2oCH09hY+k86B
f73YBtJn82Zw3ptB9vHdcQS8bNZfQ7XHpXuPu23jBDYmmpfA3VMU7JGmRa75BlxG
E5FJEuBxIjjtP0nc4Y7q7x0pggs3zI5og0c7eMmNzpI0KNkwL+bnWLw3a4DiZplT
RnqdF+MWU+GS5lbw67KgeQolkQoVpHAt0iawA9FVTrh5Lj0lwsDFXiSTu+xqCm1q
jqIqIqpTxi3hhkZuWDgmV+6q6r1S0fUBMj+GIo2ihso3Wxgz3ET8qADvsIbiOap5
mFEc7C+IHVxhbRGlHGzFi8EdrfFmXziOm4zXAG3Be+AYFfm1RkEogGwkoKVzWjy9
BAnbjafSn+uabemsjbKdxOX5axxxznlkOUQNuzg+89yezxHgb5KPmxMtDEgEdBVI
21QrBrjxzRcZ/hHkR9b2APl534SqdxoSz3KsPzCrRMpQpcihJU8b5dpLvia+ujBm
hKfxbARsa71nt4nvAvjWTze+oTNcmvu3M20rOCA3GErqn3QK443iO3vIRVbWjBT1
ETwyjJaJMswmU2Zk8RZ2D/kI0gRmCc370kd5Ri5OfzvWEqyDuFypeDv/u1wzn+Xs
uFmxDC7DFWmQ+3e4fu/7vMU+lH0K8304LCXtz2wHKGqaE7yfkOk6lyVOJphy6uNC
Rj5O8yzsUDr2R1CF1ZpSyyJcqix+Gi/OZ3CSxmYdNJ6uhkcIRQ4eb6bHbciC8VGT
3tDv/oVDWzHQ0R43U/HWDoHFHb5CDklQCxlims3LMHJOSv7RRotBaERsQDq73mNC
bbE9iLZ1gibRgHg8ToA0nsNdCxSZh4m1pyoe+N1flP3XQAjwFQh3UAY6IGKCV2fJ
inSlDDhMY5gZddjwd3gSFvIIqUpjuO0kG3IJ/I97BuXdpCI5P4fghSrGYq8jgl5A
aIstoV0VKyogKfm3nul83g8UgbGhpBaED3kc+W6ExoYARFF7lPyy2Vb8HGj4GJq0
Tsesqgi6JF2l13JeTvspNYwDN4/EvSvY59Nfpr7bo0Ye77Bq2aDeCLR00tPnDdie
0YVwMfPGhS7QRFla0gye6JZDF2/QcDQTta5OMkU1fsbOfB32dxxqgDnSjF4/084G
/TTOdw4t1oqYlfDMWVrFer7hqVEkTMiU4Sjg+WnCrxHjH27t5nz3i7hCs2PpvWk9
iXErq8AEYbfOW5bMm8rHCjp85wxmwAnBRH8UVVYw/LZKypO4PN5pWBUufOSsa6JI
4JVoZ9hk0Bnr7EbCoHmEEs0PbiTf8+1EaxRzBVWINOsruQj22ZSEd8JIKiIuH+k6
2fs5efLM4vybWzSX62oxWNNA4DhoUquyf8xPup/7Xrxvc/XmB211J/aUOljb7w+f
LVApLlAJoPLnuKuBFbNxpA87lDmsgQuzi7i5IfEcnIhT4YmdUywQ/0qncOf2OQJ0
MvzbmQ7g7Fo4Faepb/J1H/oJ1KcrCBnfxGMtuRv5BW/xW6TOYANCpe4MRtlemryp
r5oJNmsQkQ33TRXRa0DwzyEY2kErMZnCzAmijoZGUuXh6k7bibXO8jT/oN5uF0NZ
jHE4NfChi8Yi+2VeKKbx0NqnEURwgZwsjnmBl1fDp6p5czRH7Bb0jfQv3L4hkuFz
qsSYdTIEJd8Tb5RSqxIyh/zyyEEH745OTINcLtgV8xH3Wdt3lt01LFyTnTvi95j8
Fe111Kg1f9g4kPO/5+BXIlSuU6bVGMEz2IYjaRXoZNVIY5itsFQIhrqmgXbuI3My
tPYX27q9ocPtftKheRn+iPt2cKTdxkN2J8stj8VrUknKpbR84oT1ozZJpsWjyJIh
B+gebW/JUjKX/GQrun8UQEDxLfNjEk/9IgC1hu5aUTs6El8fRkfIos5r1QQsFHKs
MT7tkH3fbCqAsvxkHFpXKhhpRGBI4QI04MMnZjXhlszZESl1u2bk+P6dnklhZE9i
KSLUc0ZiDNENEytUVHTLzQoIDSPfRKDT1MZw4b2+e8hiqzcxMITkG8/pitljVptm
r0WyrjI6r7LpXFuGuM55d/DiEos0uGLVEuuky2GtL8fBizFJqXal4T6bfdgh7J2r
4xS5xkoAztBDZlgbNM6DakW72OetU2Oyh3dApsUjAWV30hntJqmuSLyEr1uTvU29
MOc83YPAPtmFX7MjSHywOKeUnYajfaBLUL7L0rY8y8ImJFmL1+SPksGROLR8wqCC
fv8QdWmqGUBY2n3+pklzNLxVnVXL7sZrx9LxSwBzw/g/rbVb7nkhcy+Y/ljkhyOu
x5EVmxYbyDRv5wEz8QKhtgDqF9MXLf8H+8O0ZR/HHAMG+wi7Tlpz9Y/8h8WR737w
+M3wm+sWhibkphQWKdXfrOX1qjgZmKyNDLJcg3F8FbJY2euZjX1gLh2qf5uKoIwh
2qU0FoenjCoxlneQlb36yxVO+hx0pCtx/mvtuA95ckVSHfCxwHiET1XhttRKCTrS
Omdos8z0ESZsw2hHobj6ZcWGdoQUbkjqbeJVphj9lzVFLFFAZdtqH3o/rSRhG3RT
D4RizuyArcSmnbuCpscu+0KOW9Dk+HFF7j4Z7prW9yjEU/YcN2FNUTKE3Uib/zBc
6MyYEA/wpcFoy7eH9shyf3VSqtYpbBDMlT27lrxTPDtJIScABS/vsmOgPKa0XBqY
CZ/lbMPQNdllAiTQe3FymgEbMcdbiA8YZ+2qzjpTzBJOSI/V/q1aXkxrebtq+kAJ
O6rpwLAeXiV6OixPAIcwpBPAY8Nz7t6/HEA+zKhDnCxCxxVAYGRSoCgzqW+gUYxU
f4317Mqhfh6+ibakEIuiTiItAPJ+h9FJbY/RqaTTI4qKoxxVRqmNJeqVTMYHWY4z
Aoj+HdQlTQqLyqptYReKOpHybECxGHyQ5ngJMPjutXN9bJYYswikhqa2n15lBkWI
U0QM/2iMfdCnHM3zcZccve7bPR6J4t+3D3Afbhpgnxjf7RqM3ycru8KBF5ntF1xM
KMG9Vp7MCePhLLiojTxBl+LzjsVsq9X9oDsYl5qgbxzNkOGdHmWHbXlkqlpuzJU5
AxMkWro3fH+t5PHOVWE/sygFz3KOx2r8lArHnc8ZuX8OIU5RSr50/PYzbHVdInRG
5PB6CXrbam/vvz8rNjsz/N78N0dkI5krpwqJgYJF8ayPg89K3HELEl+rQwPebJQL
ICOJzTYefNwgbppOaEv38bHiH8xyAxXOW8nP9IaJcTfRIR6L79Q1GiwjN2kRLqFo
3FM3c3beFbKrm8MJiEGakoEV3pJDI0g++DH6G6ZjBIHBkfj7//6/6PWyUxDAi9AP
xym0sGNpKTfyXggTT7adMrbxeT02DcN7kUrGdlxCpqHSz0KVsA5LStk3klLNpiOy
XyPhxCBwbXcY1Az1J4uXu3d1MSfLiCQcoc9rQgNjzxLb1nKDDqunkzX18PUfLKpS
sFKSwPywcayI0+fq3f0W1ED5il4TvR20O9Or8AqIxYUaeDy5l82brkS8cDcNm5l7
XSCO/fMV58BytlWLhskbT4iLyz5LQuJ7mrZZhs5stYUYtIUzago2GlspBFEBBWQn
bD4ysEp4DPivsDTdeCbhBNR0E9XRGZgXFOXfEeRlHIVlNa7TH2W8S8CY16dEvkyK
ayynZwqyrMOoIg+mWLFfY9/0E5iCZf76awKI70bAISi2GsKhU//EP51egeQ0y4cA
pngKz6ABjJn+n8m6leLvHw9AmFQ/kfRxGqytuX+mJeg2ka7he3AGublJRDK7QvAI
b0LC0HCxTuT+QrktR6CGkTVScnGqqYZB+MGgADkTaVhV1DdvzTd2mSNTzy4jZ+Gy
dpo8Mat0b6f7/a8s+Ly/qX0zNm7VyzL9+JLvOJtijYbBLgIN/UmwHiQp5vNJXTb2
Fk2HJk7tW5uljR6elX+V8Qf3rh8ragQ5NzrmDGd0RdHrqth7Lu8ccOmVlmosMA5A
leidqUvChND4oLkoBKTmEbsXCmyrb26BMb78Tf/EaGVa8W2dXQsZJcWzbwy3rttL
gJtmqpTuEudeIOJ9xkkneK3DZApvDWp4n0r7zkW2Hfea9Xo4KNsJijRUPj/P1zo2
4/FpF8kDAYlf7vfHCsNgm00/6k7AkwsOlc0eckS/R+sCCY6rq6H633dYc4wX+fV6
5QmPa1ZnbVIq1qUdwAC1pgC6JEB2neaIySXm4PAjgdUesMD/mv71HHwi9EnJ3R6A
6P1SG2SS3mbA21VC84QahMVlmcVIexZEXSGXgO5Zzw2h4o3sJUFdUbRSO7R/fr7f
V3AzHYMtgceMSKSIjXIoIONLCidFTDQ64yAz+3fQjRVXN85ZL6JVbFhRS4vOg6hU
KNdOc2Fu3/w/xgW1JbMlcUly2KcAz9hPBbK7LnNDm/MO6npJQP83r4iOW4F2AwKn
ZvpYnMa3KlZB7H0mPlCyTmKZWcexQ/j7DZxu823b0DoYCqKgNnN1SWsvEKXBx7tZ
bNL9FROfHg3JFuFs/poJE3O2bPsyOjbRqLxoxLzfgoBl+HVhnD9rys0D9fV2zXS+
cq4JAQpQ560WmjW4nMtNUHoxmZICu7cS+9IXGn2irocdIgrAOY5HG4uoUcS2uhwf
Oac4M131mNzKU/b8Rf0y1Zo/O5UJAoLFLFxtERmDnrslidF4fGk89gwCPtDjpcr3
u8lv/YczrMG1SHEapRDr4PTEgkdUqIM5a+va3CUTf+9meqfewYs+bt84/FzemLiT
SrunDASDspeZBYIixXDqSDIg0ozLbs9nxLK/Kp1bDZr4NovrefNXbduSyUaJ5ZuN
StFNTXR+bQZ1rv0gQvD/w5pGadOx98ShE8D1LTWlVKnnsUbsOoMIp9u22PZTDA7b
BXzRTOaGVjHluettBcDbIMn9I7Z3gqt3ymbUf2XYToDpsSmDgoqM1NC9owL1ht1R
h3YQzrc8YT0kZjvacNNfhG4ND87Y3FAnhW1yrPn1wnameRMW3hyj2bF5V/oBQzQ0
aXY6Uphd6BC5rKkWwVkNmTpxp0z7ldLpblyM20dldLI+Jt8VC7Yt4nHJVqdR8UPv
vQ/xi3z3Umw0ul82QDnb2ikxv9aExKXQUyhGsuC/ru+FjNZJInC3fg4rz19yF9Wq
qmTUhD7vm83gH7FtdwnEHS4+s6y19lorHVxKStN+4OKUpEbTRJ4RJrNeCkF08DZE
5nGdCSUEjpzVXJk0FsPG4ySAAWIuA6kI865weHV0MslP1p9Z+1yDKYpe5mVA303A
FwAcWi+3+QHJpqbG+4O0PlGzxEIDxcMdEJlC4KGQ/TuBtCbjCLI4lOGQ332GbYRm
5SWu3WPKWDgCjfS1UwFFSfDnmXuCmo32DYD3K1Jfc0UXYZwrqFRHx5Jq4lCKG8iF
mgq6jUF66NFZ7uUgKd7bbDKeeKSZWp4rVAv17gI/x+crOQN5mLd7RVT5E2E6MvOY
cBqJXc3CuaBnEYG8D+U6M3fAC91qNS6nkzL0qPCayjz3pAZZMDOpRW9a6V0Vvjtq
hDWCPxdOJJdvwCY6/sxUrnQJqE8OAfl4utUg2dORV6IjKEuCzmOdonCjMNXyBdZ8
5LWKhkXIvRCPX5UFmTUiYimHAx7uz8BHBk2NENPiAU+1f3n52aqZ1tVSpLAPC26S
wq+cj41gElODxXZGCOvJhF1jvW9S/2qPH/WAew4pOUwtxik9CMBbMeXjSsEuk4Bs
Do1tkyKFB/EpY/U9SBCaev9XWyz0j02hQMKhPSnoi1eRnPZCGbUjhGrSBjHIoWjY
AKB8HCl11oY+ORLnBrDMMWwYBjoMHdcfURe1854udhxxQcrONANa8wTHYT99wkBv
BjI+ysIdp8iIE/SvmeOMnkzttHCRy053oN0d9z/7ppW+6Ia5qnT3wXAwZYBTDp2X
ibLHPkNVD+QEl9vd9mXlmsWJUf2CjDci2q84Zuj+qpBPnAkikqfS0M+tO7sgAyX1
OthnO8Of2Vx1YvtXAbBWXYLpvf9UoINkSCQvAOvceO1beJ45boBdvo4QK4Mil8Pm
GFhUYc9fcBXpqbS0t4Co7m0ZEwCgHzb59ugSid1qfksVsCZrQ3J1eRFiTeG9+6DW
M+PUZTMNCJuxeJgKWZlXXt9UP3uhmmaJxEgFK7EUU2TOBe5OUqdp90dA/dyUJC3n
7TkF5v35keq4JsOzWAT3sJU701au/4II+4oIhnbVZ1wQ1cYOTLpIhKR9j1mvG6Aj
O8zxPyvFKoB5EAprUhpHP6VIUvxDq4yxUeinUw0VS9xRbd7WUS2iYst1V1yO5F4A
MqgFCsKVVP4M9UtvNBLtlGVliITOR9HxxY4rkrf3+vv8kq+QDZTp+iYAeM4e2pI6
tCwGReZ8YuVAQVS8nvqvoE7hGz6iqUGkCIoS+y01qkvkgDfsznWAZ9P8vII/drk1
L/xp53f40qKv3g1GDy/haX5HzuXrCY3jEJxHxpfZUv08/D7IgtdEi86oQNj+Jqb8
uP+ZI23ompjvIwOksOSH9kOtRu7tQz1F9kEsrvVVpZmZlk3+/MY2UCqsoS1eofVC
TYRTIcug8Y8ZQJkPJXsEsYPCo5ARh1lj+faCpVEpS0/5dxXhzL3s9d9DGoSBXVlw
AwAPIgdd5ZW32jS9BVIU1FN0MeZZHb3z69mo7JtEcre+2OK6Q81jM/u6jrKti8Ym
4xvYZwyaHckAEj9x3ZR+AnXZYf1x/gSId9HHgD8tOLwkV/3bgRlMvKj5jDwBIP7I
9amOi5QUNSyifBU1NtLNs88yBEULc3y6AbpIGhVkxOnU8ux+ULn+ABP7buBJpqjL
pMNJESSr9B4aWom0fH/VCTz3V4PjGlRwm9VD3KIP5dXKU9KYZgwxzitKusy1PGDD
L7kdodiLc5rNbdrnxRRyhMPb0Iyjyaj2tPrYcdYZJfIJ5gYQPyxsa68TiNTJI7AT
UV0HxZOV4lOH+NqBBJvE217QsXQ0nIGbP0xdTOBpy7/Kx0qus2YAXXOExY784s7/
Tfy0KRrHt6xx4XQxp1FNvAU4EnddSod7hClBIq1Zt4aBEI2hpkieq7kuZLgb8MCV
6+LczDvQJr1A6sLuTFjAkASbRHxZ8ov/I/ErAuqJ6zezfJHv/7mxvlHgwdBEBaZ8
PRS5mWreOXZvqeUM2s4kI5RhSQy3yuziHRR2jNo4AUYWm+qkL+jtXqhq+Ipb8d6+
JEfm6PA2zkqTUXeqvjAZ316HmXKbcZ+CMmLakMFQEIAZbSuaxVLk2WdA2YiuuoF3
i7zLrHKP8jvhz6Y5KGewNl+djSYHnD9XMtSZGd3bqI5CYAlbKpGjXdgONCUFG/CA
ESRoLnaBJuOpKG4WAIfsqyaePa/+M2BOACl3xPO1Gd82wZL8vmo1q2YvcKH05FkZ
AdqGs/9X6XYuEBGtBmxH9n4qxBGtmUEOumAYm8XEWMGn6J2BXsxfCIwich3+Ihm2
GyPeDlHVZgfXTl+G27y2EQJKHsuwgiev+YXM4/Bq78CHJO6mWuIOd1C33SwoNZiZ
frqhmT3EZavQs0mFpYpphI+mF6cAlIre73PptH2E0959OIpYLiHQopqY2i7TI3+a
oEU+Ok9rFxj9J8Hi069x3ZkQD2+ciwiPCkmY63xv4W90hyFAxRYLxobqQpNcZTBf
V1EM7sJf261OrVDxLRWKRV/4/trZGBz2QTVwlFhz5y4dn14YPHjOKNTommjznX4f
7jvu1+/AtdZAHY9tlLxCGy+eG+9GdL/uPrVJ1uPIglasdY7U5NUDgC4pQKYATsKf
JBfKmrLqdGY1ODD4eToLOl1nO5VVeT/6h9NjGJLu3nCLVUTNeNkewGGSk3RpW/li
TR51RHGWljMEExFEBvSdMgcnL5CnGKbbZmZYoFLtbDTn2JLHfGPJ/+/k26uP28If
2FWX1W7zp6il8QE/+KXOn7OR2bkUCyodHr/nWeU2JHousg6/2M442qqr88YLm2VT
cMoGxIZKtrRyaOHn1BCV4+c90pd7lX4zF4fXXkXCq/WgA0M9xcju4VysfleppIE5
ZexBxLKj3GNpEs3n5+FW1z1n4pPPCgmrIL6bw63XJyyp+vgzk6AqEXy+BgedQZzN
OaFD+OVwJgMrv+BVgudLhrmS7wETN1Il/6uEH0qr7VV0rNL9BX9CBk6oPCvXRujW
J3pnvhUIWgIfsshjg7dOwLFbaglYXoVpVF7ZBJvbmX9WOXCzsOl8B+6qf2TbWcLu
E4tBEaM24p3ae6SkRmQ1dcu/jmu6fk9zNpIR41b+Hmr/OyWSn8i5gCGMsxju8QGd
rEW6LHUOITsDcFpHqyDP/7k1Zk3RZZx7hg1Bcn+gYbLPmS6QR0KD2Wv4QFfUKi74
xJt7Zth+v5ONWvO8yB6jSWlZs8MU4aXAfYYtu47BZaBGwRCpOajNUUW4YTIHyFyh
2rgm1XzJmMqjbMQbyXmE0on0NclmdOCPOmHHUm4X+fZm22bNtPuVMsi+ps84iyCf
Kx8FJKGNXSlpIiUkJhfvqso9Fli2bUVobpm2K/rNeT4dVHIGGaT/OkxN8EdDKQmU
91sK9wG1KRn0q1FptDnTCdi728QU9sK33eXxFMfTKQjSNQC05+Ru8HlNuPimPPJ8
5FcBdDmSw1aiMDAfe/0sKKHFkm4ZsMnfaaTz6h/gypBD1ZIbNgh8gOQ8W2Mbv6fN
PEuScQt25XAV6wN0WZOfcK6R3Pf1sBjoFXJ3vEJiyXbhNSZiSWNdyFN76H3IWmWY
515ZE+U9H73TqFIL+F6rDRrVkezgUClc5VbWUgBflnvgzUI8s4ntFVYm2VTEaPoS
hsC4cxG5gDct0VGgOEQFJeGGW1iFIbaxs+ku1o52OtF216COJgZMnY42r0Zx13Yx
IHsfUJJ8cqOJqZ9QSrQcgNNy8VYTf8L/nYvCU56Asx7XNf04aWLPAGqr+vlzIIOV
uglh0QhPdXKCApJYkhuY28zNK1lkR6Yhio96iLE1JyNjGNDOFYdDTxU0CclREKuR
BMyvnqaLQbXjWBqyBOdnxK/zuisuGh4sNkkPFxViUyKR5/qCLn7Gf2oPJPpHW6R4
KSx5h07cfiGzwVQH8hUKxZKXFWYK85CfZGApgyM987ZJVh1cwCgqPp4GpzKqvkII
1TI0hvVxQ3tKUadxFpxAEp86OpPGu4FqblBeG07PKEmsNXBJZVWN2yugLMKfhWSZ
QP3LexwU4LoL6pnitEs4nTFoD1iN4VAHwLeu6KyZNhNen6Wlq9wD4f5IU/rUz8Y2
w4AfkDGKwzSAZqXa4euLdM7njR2KX85pPuCQJipwfQQi+uzNbZIGdLP49nL3mutv
ruvb1GACG4x2l4kuZv1FGGBCkcfeOj6o0llDgog3lJbl548aTHMCjEkL7396qLte
JiyfzqV6QoaVW4pl3mzndWj6vvnd8+j1baIhsbDY/xNCRtq5DQdNSk1JgEoxyCWl
bNPGbpUodjomldP1m0TNjFTigznaKEJWxR9RdCd/gpKaf1V6L/+rqo3Fs8vyFmF0
eanwUt8Lzjp7fRKNY1pSh1nSpcJLfHytdCqe++83SEgXth4w89aBcUKhl92+/tZm
Ierw1dTWjOpTYMce37sR7ARGMIeWye4awZZXs4vjYRltnLaB+r6f6GsnaSiXqBBT
EHoja9MqMGnKNQwAJvwYZhjWK4b5zEC0f73ADP4n93+mjQ4s75O6Jz1m9u9f7r8e
/IXJ8ey4drgDAENP2FsUV1m/atzkcLK1jyEk8KwSY11MddRV0K2vHRsNJTOKLI91
m5PXiEY1vgIrlXPj5TLnbbE/7gRlRCLq1eExxMpwO9Fp0DjDrcM4dvM5mKR6lYfp
xEFiXUIOOOE96UHUmRZkyKSCw7yNpYBtGGQX8nPqAhuyc/Sf0CPEqxGNa4kdroxq
rp2I0npOaJZBe/fARTY9NHmj2tUBT1EYx98qRT7QFm1mmK9jtHYE892oUBekkw3/
lO+meWVrHnNA7x5QFi9OVzM32XBtZPeNdPm+Qklkj3OQ0kOHOTlgVEAghphzaCqt
5RHAsnzNFI31SWKUcL1+gObSvKAX3+YGMhhCsoyqDCPq4q/a6jA7gmfmWVl98BN9
h9arh1URH/hnXOcwC6g51jA0JtYmCJmwNO18aSluYWMVOiuttyWzdW1u1nhhJITJ
su1kq7N9JPyvUpG2DsOA9OeCi4yznQ/ysX1xcJaM/iwBmdALKzMvx+UYSEvq9LaR
a2Is8G+cDDMhiHuEgQRhcts6coM1cKAtlZyQlzOzJoICIVILxck53nk7m4tPHK3z
c0uXCZEjK+pKPai5+pg+7Zs7SmRh9ShtX/4rCWZwL2WWevg36IB8f/msgM/cPSm0
WJN+j4P3lLk0For5n6GKlm6FVYL5Dkhr5bsd91jb41cYK4Y+IaUUCfDSLdxQoyUf
h7/1TR3VK/033bXWu/Bw3OFqAntoMLzRmAfigHFoIJkfB7AL0r+grQy4y5y3qfVt
pSReAVBu6VmI4bG/UeLfZ4J76LHP4w8kWBnmGyvGyk414vi3P/XA6fr6BgKbEV/h
7+RV6ceQNtdl1/3mEGvnB7yRUz32UKjKXf8ShdsbUDT9JjgjrhZjxngHUwbd+HkS
ryETD24VFPfiNJwby39ddRUOr5dvcXW1xJDWO4NY3YhR+nFbqY6qKnvHu4fK9db+
evOQbctQIWUQg+IdqZoY4U1lLKAfLQgfkA5KwTGWDSFgVfQew5iT3zfyNgAGNspm
+1aEVDrSghipCi9bIqJGJgJwIwDzix1uEcldzX32/FLGq5odiZnU6h6+32R4z3PJ
0fBDpGHEbOFzVMclhcumvRVxc1f0hP7ViBkzAxPii2YS4eOFOknsy+GQTcbZq4I9
qaIOdx69LBjd4+sp9ATtxJQJa2Uhph/VK95ZJaQrCYuwOVZwO1j94NZ3Kpvev7wm
W1hZCNakK3Iz8RjotSl2R8MCzqmaymPCaM9XRnDEjzkXPYX9ud1iGN6HmrWWk3Aw
m5MpRRUepxZ9mvOlRTfVe1AdgPWHK0EJrAx5HDT+9pgB4PFN7idvg/Jpdw1dgTkZ
zqzAt8mp+GH48NIy59NFg7OxyNdhmQQ+kQt8sGx4uVoq1If2kFkUnmhO5spyC8b+
TAel+Q0Yi1/RxS5nzcjvLvE8BgY+o/5rEMZ8fGyvE42NGnPAZwGSH1Roup9wzfy3
cCMP5aFB5N8rKFlE4vcjBScUk3htSXUpXtXH2HSmYHHGWrQspXYKDksfjVGzYXGI
RFmIOtbn22xzQwKejS5QmPc1zUHorYTYQbtRoXmTKNORDGoWFBwIXX2Q0ISXm9S/
HkOZKePoVaJmQDdHXhjLiR339AxpgFg460d61GY+OY4TC7imaS/HxjpXmatLw3xj
U0DzEgABVNPl0m/kAWzVjDuUxZL+RFlW4TwjjTaD8VgWbUQSiylDXxxaubKSlI1D
LB6QJKM36KMVEzbUyNXYvzNikun9Q2ABzP6h4b7RP5JmQBlQjcUow0GYnzkHGf9S
nOiqEVn+JYNIf+TrHgqOQhCHz4sMx4GbRa6UPzFfBJajK0i9WQrdiujvKUQqNhIF
Tk7FNsmD1pASJH0OTpIe5fEBVsv6VV+dT4RKJSE5ke6IU0E9saxrrMiJ+LGdjQk6
BdbDDxtjfncnA0ZX5yjeu8EeaaJEoecM57RJddPu3Lkav0sobLI4gM2tWh+9vp4d
7+InKzX4ni7ksuB+Ma/XDw88O6fohDgsacjx8lfPIMgT5reNisVEStWIW32xqGCS
MazCEItA+ZVih9XB5zoHK0TgjRCh3I6tBviD2/Z9cX0zpJEb973RWV74f+dvxEMO
+4/ws0oDKZ80Fv7x0SefTrxMSpshTdDaGcrzYo/rRUdC8PdglWufVZfSSg1SAXKq
jBlP0i+9GuwEpQD02bOhqNLmc6dV1GTzKmqiMBVLuuw5Jphq1nrk6egbF+ax/l5u
RytKi4PmGehByJajWfnEGzydO1wNCHw8NHyTClmSIrxWM6EhC7p86yvyHm704c1y
9HPGbaePNAIe57hXQ5oYtPmikm5d20v1p55T9KYrAH8+fzW2Y4+3YvbE5Qz2WXca
ZrwZQ5TwaGflbwRiGB7yMJnSD4cdxLa8mB9+74sP1WjcS5DmxBgo95bLk5/lh9Hh
InhORWV3FDAW7OPKgemXpbCTrnQIBs/+9QyBVW8k7g8VIQPlFOZR31S8sHLqcWSA
lC8U8ncd+6rpJeQWXXp88E4GCiiTZziGruo/UMDgTq6KwQGz5LF/YmJUHJgHC2wM
w5ocNhyHkbRTsMAL62WJUaJsi/F0J50WkVHb2070Q5hc5hQmp1M7TOzvVohWt/eQ
NjYd/JQUI3eQgwVXtOiNN35BbJ9MCqUzQEC3op3Z6yRzPuRS78Xa9anybPrctZXE
5jeS/gw4OFoeWCeQKiJVK69kbIFmSno0X4+ZJHoky6J8bhdkuxviwvdWKYV9C7RO
dgdl2oV4kpUr9vl9KSLRwZlRvc54rKxE2d6JyzZ+6IjUFE6XbU+cDF0J3mt9q98u
xVRBMtXIWW0huYRT9qhyXydU0Yuftv6p0yG4l+ybzZ2QZdC3rNTXdckHv6Enupbo
wsIo6Tf/fycgC/pb9o+Ck3EQavGqKcvEt/7ITe5IFMq9ordn/FrRdVV3UvXx25qY
96xuS36Uiy3LRhSWbYgmmJg4GlG5cdxJRqXWswG37neOX8+Rp6+u3kg8vU/faU7G
z9EVQOJR1VYpgCLukbtdWsTHiyUTYdxI2Pmmzy0XQCIW06UM5Az/bKGdI7/KGynA
6hXLq7XzuEPOyjhrzAJXTBSNhHm9GdptUg9JOmiXZwH8YDjlxv+wFKdY10n6PkFZ
nFsHUOdBNGqJi+1XoMOIzoiOSbSXz3mrgOrVfqy4cTEoFE/5eJB6MqyMS4XNhZiv
B7FubErqKIE5bRrtC+HB21k4J+F6wPk8/Y6VHLNT7PYnYy9HAKM5m4C1gPDlj2eA
MSWvPyfYTk+tUUtpuhJS6YbFTzvZvWt8vdfM08+ZzTFDz76QggVgpRA3b2J03u+u
QWBfpoy7363vgfgHc3F6nzHBW7thIuZ11/AM7Xf4pv8x+NfSBoRvevpHu1fpN7rx
VO+RmmzoH83zZPVTov/28Ft3L98LF3cdq1rZdH8m718g+PluLLiGuIsQV6TMR6MF
9V5EU0eWyKu2JJOI7zMLug+yEvAIqlxFUKxlbRaNsLylcfHDx8l5ZN2q1IWiQKII
zw7USUS7beeETphZyy34eHM2G/SG3l9xmVuM6+bckwZT4399o3jcs6h9AkwTtZwB
Hf97QnPDo2Cswl+zJwpeo+9AP8Jf30ZnKMNFaY3uuQh0587evdB/EfiB1ns+Gr1J
3BrTHSSMQgNfstOcuhT/C1UQTWpuDu4tW/9uiPlLGsAzkkHnO34aQYKi0zYgd+R4
bWNusnlGuoLvkK66HFx1yeabkrXrbkQga2TcUgba/LLkWOYNO4EmPNGEPPBzcZLW
hcL21f69LCgYIBEn5QODFCL7J4SI1mElkOZnhKmv4LN4BiI1ZzUPYRCWOgsFWJ3R
IEtNTr9OOm/BaihPHG9chvFB/ND714vsTc2ZhcZi9ekpb2s/+pP/PyVb3RL0ZHa1
DK+j1P0cF6AUY9Mxhul/TLCUdqJPG/D0mMSIM5jJudO6fZVuU/iLhIJzyRxBscOm
S6Dl0Y7zulIzZbYjVwJd8313IDYPdHX6KCnIk51P9fyT5+6mVp+2sWeHF7jxpBDW
ICmYQm1nw0DX6oqlCPGXJK34OCgbwje+p2jSHalZ7QP/uY2uCg43a4PacbKRab1+
eBWI9wSVS9CGeAxyljyid44453T9J2wquaTHzxmT7EdmYcZdf8fa92XDA+D/i+GW
AaErtXSNOM7qSGw3u0OPELGWuRuMDg0s07AUMkbrZ9fQwGvG+qsVu4WDGanJN1tm
A2CVSxlsHskAhbPLB/KZhzccpvyuUgrEPXVFEqpPTNtwCBRAPDnDIRS2IMNXC3D6
9mW44AX34bnML7Btn9wb2agfnEMb7vOdb1qMJEoBMLOwkDSRq5pLS/rctQ3SqsDY
rPcHm95m3yQCd97zfJckHjoXkdb2qrGu/t5EfD/SCn5BVX8odzb+2Zmnro4Nvs2U
GFesm7H9le9RtyrDBDf/w0ajvWjA+r6dliTChDJxNgo41yZrLlIIm9Dc2uO+BOlK
/CkkiGiaY/EFnkOmJequlj9y9NbqDdgQ3xv4BH6J+dNxacIbp1JOX2ABJWZLCwbU
WhsY33unCJXs0vIHPJnBz1zAyqa+zZ62zbikftuHk43z/X9kDbGK0fCeQKutySjk
Iu+brkkFGD7HOaPTOmsc/jci59Y30Ex8SnbOSOCBmoZkiGLpl6xG67hLBYlbmGFy
AmNrWTXqmm/YfKqXUXi/JkTRgexP9J3JHST5l1YGoctBuJ3iP1WyECmJexLzUrHi
/1a7d5Y6P9LifajvVHZNX/7Y7V5svBxMe6jWgXJyaxzD7BwM4TWq5ZVwjdG2DZDI
GYGmk0I2Us+yihAFm+lUzdqKTiKpnNL24Di11Uvda0xUCTVi/bz23XN/NPbDaHzF
ZDhLYGTsudX7+/Qmf18AA2VGO8abRv91Zcb2m5XDhQAGFqFqJT9KvTBYImCQBbxq
WtAEYmG8t03i7OPJWNpcBKErl4VE/mNfLobHok/58fJLq1wGwy+asucHcN4xQIQM
P2DJxRwfooceWhlMPEvi5XXINik9r63uZaPkOVgK6IpQHbFWrSdP2UFHRiHV+rJc
fFRYtB1mlwnvxmmbibBR7P5PI9PplvGBH6YzNboqAPp2pnNIMDmifhmZA/0CtP8w
chFh5hVKNJYV2Eqm2QLcBng25yF0LDsck+PHKXsPSJZk525LpA4QeBwoK4upvOnx
cb03lAvPRxhGMGertxqZwT/A4r9XD6V4dXJ3SaLfJs14SXRz357wftvkwIgAjVGE
FxnryK+LQuXbptnfQc+X+eAl4k85lIlicfAITlqJpIzGMRvv9m3XG4w8vl9IgPRm
iSWr6HSDRyuRY1kJxgf0xCh7YEtTMwTRlbPF280R/lblUwhVgXUS73kVdmM7HKK0
g7AtVDHfluxcuflD50H1vYGlEW2Ln7Z02Jt4HBa3vUIJGsNKZlUfVtc2lb+CxDwA
mJBvWFOfC4pQPktb2XtNXihf+FF+y6QleFdBMKJzImXcfUjgS58eLx96cR1iPsK9
npik4WOfx7T5XcxqEIKG9L0zIrGmhMAbNr84FGjdDYbSGN1sg34+J6lDobY7k0H7
dGN0A4rrXDH87SIQlHbm4fp8Pqofj51hT/9Vl2gUxLKSR116ivi7lmk0hrZQTLy1
ig+mj0NExmH2vQjmvSwogi/Lwi7bs35VgxPYh8XLdXcZxEqvWNqYzEs/w+isQGdQ
CjFIuVUT8+rQgA1t5w17UFJQFJ8AFUhdLCspKwvc4WvR2xEjO9cQBByS1IulD4ny
6F7NwoGntX7phLV0E8G0ZGG7ooaMTq9QQD/EhYa9eedjTDlCa204bnQXMfNu89bu
ge3goZmVIMKRkzDo22mLChZZLiFcizJp7/V+ZK8+ctdZy0nIl6VP+F4ueSKMBW0k
kn+UqKgxvO5l+QNwZk1xlV2E6mMav22zBpK5S7u6gV2qwCIWPFrEocyrD0XfEc5O
7iwbuJxPkohuasrQB3r5YoA8fweEJZyxkMEqgixw9AFheZyktj/o68zavLGmdLbr
73mMuki3f0ZfGZvEJBP+P5kXAxacGJFB6zQMBWLt4r0u51StIi2xzw8SmNoTyVBz
qWGS6KRbFBCAfDMU0e6iABbVkANNr1MvPHmQf2S6ImPeYS0cobbD+QDY5zA/X1bs
iYLLnbnKPIBgqLJhPWgS7NFgVL6BWUveRQ+mB+XVR9wM+ymlqdTadVtwpKqZkkMm
JzE0+7V7s7mlmwwk0tCYUfzlQ5sil3mTTvoRbPZMqeWR9jaEl9UhYbbh8DO2OxVn
QCEFwaMS3y5Ot7752NJ6saxz65HXoCRWYvybd14UFjgyVCljfNnVCZo8/fghZucn
JX+yqudAS5DoaCN3Nl0TzSRQuiJW95rzYIUpZhgEFfgtoYCZYNlHcauCKsNTp0ql
+ex558vtMU1lQjlUAOeA/9oqzGEOT/LMMms8hT+aMYX9IMGkGXqdpljrD9Y7uROq
1hUsgPwpZotjQ11kx4+FEkojUpyEDcihWKmLYi3oOL2SGjSXBpW90gnvYnjLn8Xw
kxBp1BR94Bua9tT+2Hs6gcmne8r5Qy0czIbqKGjvCKsqnDFTgO+8K6L/2bFNzLUD
UMJpj7pe1sM/HWwVwCtN+br/6/AAwT1oGFufQQT/IlWUwZrFnF/RlEtNp51hpIpS
Sk4DjlUXCxjHma+0203pxFUxiRNRyEA5R8hBRCzOVc0uaGSaiqXCgfvmP2nXSxRO
OK4nx1m+0HQii2wiqcq5r4uz0m7ruxyY66N5ejCYYfZc/hD8sm9lbIbzhcufeYH8
z402eHSUAxxGvmFJYCyWwl/J0ribJB8sCW0enA/WFqJzpWP9pirufZToqPEEEo19
w6PV0ZQaUJVQxxHb/X6Te9RHOiz4cjL+2U756knhWVvsa3+afc5z/zpc5gU42Sse
PSvCXlFdNC+DWvH1PWr74Fxtk+yKDQvSDa6YHMryG49R0tadym58F7Y+AR16Nv0w
0njb+jnlet3j4oe0fynFVQR32klFKglrSxrzWeVAwYNLaYbh8qIBPQ2I2tF6RSNZ
tumNd/zAfPdJbdy1i8fBbBBhFB71IAymvWmg7NleJvPr3Gwre4XnfSmsdhZTTrLr
k+RfR3wO34mabxaEhD66NXVEx0wM8hxu/8tyJvTPjjmF0XM23KHZ8yvXrrFFNMT2
ACkIrMJx5rmDaObsNskcZyOz4Xh6N2YfJO95VpDmaNcC1tTIefMRvKE7HpqYEv9D
Ra7rxD5A4jUwmC/SKvnGQd+xXxUOon+jUnTGJGxDrHM8I7Ofev6iw75vk6Gq/IdK
TPZ02GN5hQpeUZ02rdDkBrtm0Y5n15c/kBin+/HTbWKcArtEgbcZzeEJ6tnjm7UD
b7HSOSlS0DMKhLontzeTOIikFIfGKbrC9PFCDcr+oiG0Yx3YCxZD50cBFNHYTW47
PoBYptsjGy6vI5Qwt9TEMOtLsTl/Hxcu05gfx3NgT1RVYqvX1YqbSgoW5COcsdx6
5vY35KOMPfGBuJHo2xdsSmCrDPRrfZ03snukbT1SNjaWR9p4rZOHOIhYwYgTONH2
TWprGjkSyngSmmMIuO8RY4X38wuSdVU/5SUpLh6QVJrHfmYEk/l2LCQ3VLUBpaKI
J/VMV50Kf/zB1ru7djGYk/JUsyTLGxQiNokeN+NNcJ60CAK2i7C1DNDtV5qDuwww
MVf7aRkKwzzj+P5HtUQ+ZF051rK/cjlrL7dsmZMMDgj2ezq17zr7I3sOll2k8kc8
Hz8Dj2iJ8Pd06XGw6KkWNqfuQ9jSjOIv+eemAba2DASxxEY19/91QDoWQg4ASZao
vaogftWM55XJj09DO9+XGkO/jL2H66E8kp8uL4RcjYkLsE1GAsH6OUp8x7l/nLqD
vDJn8+xNXKRtPxKWW+2eIrLa/475c2aGQxoH0r3vgN7fWFo9yezYbNl1T1NAb1WD
jh5kZOk9xDuU35PLm7m5KiP2mjCVocu4bW9/SLDQwc+LU9aqJTtHMWh7AWS4MSwk
BD0AwStYVPf2EHWVNdFzrvb0wr4Vp9OpT7InY9Zz1hH4OdeeNziho5xCNlgHhDhW
z7jptWRxnDpn0bKUfrpaTIVQqYz/C8qqfTZ/rj4wo3AarfkD+6bqOd9Czm52ZB06
ulR4LsuBjmqervyN7Ag5GRqiWWBhtBzykHePmRMmd2Lp44dzVP0NoKGMZKXl7DTu
ivt2mzCWC/BAM81eek3VApem6ZqnuzmwZNoL6YPZuRcrF584vys+Q8n4k2g0OoS8
5mK5M0gCRJY9P+0txe3C7sPMXEi4o85pEyHFyx+vfGeJeCm9hJVHCNayP/4KWBiJ
t94EHlqteZK1gHTvveFNN/EY5RY8n0k0Sue02Y5Xb2gahJCEGvYFfH7IsYAMw4HS
EhO1JpeUr+6lugVDJoI6IpUvVVuwYKhwhdpC9zMwzLSj4jP4xKDT6b0EEymh4HKj
MK1A5QUxHSslw6HkqIKJwF9rwtOoM1PfP/XJU5iAjL1QWEBE5CLkYUTr2wylUSV4
aZB0M/mDFAEthkZMaiu3J2YoX18Ybqxfp5JAgzNVIPY9ymkmRyE7TDD3CCiyHbzc
u25gSB6CO4DbF9i50nK6WYzV7lTaW2jsqTuMk5IjVYatKe5OzGS/DFPlJi4k61W9
N9PCeeCCqWsSeu/SVtFkWt1B6SFCWTH8HMgTktVH9SDeZ581RN3tJXbqwyQkHI8/
BthB/5OKkob3DSszrU063LnP/wptwdLHichKAe6VMhZ1p2NxqPSgTeKeVrRsxqCw
56J05i7/ZQS2WvxQIOH2dnDKF4Mz4HsQZFTQD9znbgSm4YPy0XRy13rV6WUmJo1Z
Rol4F+hp/2BKXTGhvPLQe0NbYauF26G+ZJdj7CetkgMz+oGoIAW1guG+U5NztNtw
5AWcQrof/d1UHIMQt9btAUwUXkjYWT+HHJHRL5fr+ygVxsHdlbT/rjqB3T/SzaMh
vWY+BpXPyAuYZb1ro1h5EB5IeHW4jfoiMYT9OFpCZwvzkggAdi0CAE+6NzpgzZM+
kpM8HtS+kn9i+lXdOcN9FOTujeoJoXzHdb/lqvuAuGKaV5vF3Nvt58A/jxDZeg5Y
x3/lzpa8gClPMaJ6HPNER0ONMB8e9Go/h72t1MBvCfgUcXEi6NnzCmK7/dZaBEa1
mwvf5BsATK2F8bMKTI7Kn9Jv7eZPmHn37EXfTKmPcSgb7E6x0IaMWL2K2E4Tltof
zPdVqAqZL39pguEJTRzr7BXYnYqOANgpMjugP76aTYW4mbhC5cx8Np+Yyzv0Dx/y
/OYcylGGrDmE3l/LiT3xrjsY2sE2gDo6rUCPxob5Ut07Tw1rL8J5lOyyIlfkQUwp
ObJmpXGL292XkUXtIW1uBcOqe2fiwFeFDZdV4guFlAtSfmMofGpbYWPucWMVNM+N
r0yUgdGYMc42vN1K8+xlXcmAK5gVy8AuxBk+XWnArIbVGP/Vy8wnKObQzscOghQA
2tXhOtkHpDpTtHZGqDFVqOreSO+OotxEChTraKNSF9StUPXNyKqNKF1JZQBDlNIp
dxHBv1fqsTunCGcLU77M9h7o0ffJkK4dmsmlQf/VLcMlCIx2URaklzvNeqvW+fDc
7nPmwNZt+Rhgg+Z7eQmMhEaKuZatMHuE8yoz3oyMLUNo+2H4bLeQ0rd1YvoSK8Hq
4+9QP2i6p1oKtnaiqXz/TMrbHpZYktkusDji58letfAqmh4KiA/psxb9W/becNzl
DOYheppZwE6VWb7pWWI005xaDPEGnZtT+zAG9SbDANf6n93ZEi5wLN8Bsg/G17RB
qk/O/Lo6vGeegFg/FgNd3y0mkQjG3mSNKrAe0tWj23gNUTpVQlYImX3rpwRXqfj1
0TGscRrZRTHBA8lltCZcxQT49OQfT4F1rE7fRRAb/QJNjwMS272cfNS7/4tQqTqc
X638Ns+YPaMX2lsf0soqYOFGlI/Oi8kJEct7KvBdU5c5N+xGC/AGdq1wLys5tR2g
cVVjsX5SDSXgEqK8JH6ihcBAc/5qPagyGNju18+7Flxp24OryyIx6sGMpSPBFR3W
xz923GuS3TesOje/BVT2wjrVPUfr8rpFZ7w5y7+ht+14KKR1rtqEYza40mlK+h0M
BWyYKmK6PShrT8FWOa0r7Sv4nT+JCP1DnvsG6wYWOta5gYI9yyFmv4E7yIvGIj4w
g3cAbSE9ueDPV3ds2MYmAfUhJ2JdB7Qxjd3Ll3zwJ/eN9Yg065mlfYb1xqf9/sOF
NslaaaRWMDXRKv8xYi2FZqsOdpvThEGkxBOLwe7V2jL+mrvZXezNT+K2eHiKb6+o
KBv4L8M0aoVSxEXi4Y1AX09RM4SyXcVK9oRziK67m0Bgiwoj4M6A/Ru4qMnAsDvf
NNNUhlr9vlpF0XGF62hc0pXQ8/WBZcd3DeRWtwnrXzWi8sOwYYXdF3feIdOj8QRY
SgOCKjumoZGyDDb8jQWUGoQEArJDzM1t6C9Z8SmYK3Prhz60lKErNInFPVQ4hkkR
ISVZJTUP6Izkgh6K6OutNnUtRkVIkk65/o3JCQopVIpALsIi3C89PqmJNDH4i/p/
uzjUcWUuCm/vMEpqWTY1XSh19Oc54i9BuxR8gQejJq7BBJpTE3cn3KoTY9cxBKsV
CRLT1/XdGCZ216A3nb04Cw1G0EEHhyGSR6R4coVL5ByeXJhr8vFLKdLyCSMHhig0
k5iEVZ4f/wMpTsJ0r5TBK0tqfIge2E64PHEbCM2hhGLb5/TknnYa1EupDBbMxjwO
GQVTuJGCRoKiR1+XgtM0V4Ch6x62VPD4BnQekqIbTKMuAyWGR1lUs2H61cEnYtRk
a8QG4g639FeePHilWk9ehU1jsRVbvry+Kcj73xOqPfKVT3F+wUX/GQjg9h+fkr6i
fCajCkOIsZ37Yep0WMAnDxfhrxmJaqjDjueYgdrxnL5KpEDFrNnm6XsEzu1uhDpA
LhzQMB9XT7tes8GEHTJTnZMMb3tN18lBPdF2VjkFBAOdZFFhKHJPMBjEQhjDbnKW
2sBWMtkTbK0APK+oPyM3i6u8WWkhMvzxyLeQVfsfmP86abNyKyDu92Ey53meOhW5
XZXgjfOMXAL9gVXSS3+QgEtI/Gkw+g2gEv3+Nj5W944FX7/w37lNUgl0VQtHU8B/
rEvFwfVrr2DZYqes+kodyLCOSIvC4jMwtDnGAGqF4OvvmHHVisTYpszJF4VoBStD
tGzHNpd4MmcJDD0TpwCOpFF7KNGFHUNCPXwctieA4M1fZbNGbIOcPclv7kIMzajn
6cQ6rRwGspfzui5XKzjrCmV9eBntv6MmQaObPIkQ4r6wmQ/Kuqz4TzW7OAI5/Ubk
RlhRIO1CefigiggsQbO6brHlr38bdclaCOCDvh3Od72/TckoksE1Sm7aUnBgWVo6
Ly45TNIg9D/+QTXHzer3PZvDf8wmMlTjnKLQ+XpilEt/HV4Z7GmJiknOIKPwnE4v
czMQDuQt+fQ+P6DR0oKkOjbIJMvh242ynLjxH+vml5UwHPK4WkEZwjfPklIN/rwh
0EuQYLRfAYccHyNqvPj4B1wKo4aec4dM/+qarGlWwZjxlgY9qqNG/Tvlr60QT1h6
VxYLGDbqjAMiTy4KANiY7CmnNalEw2wreJ0AE92Ulf3xsP8ThzClD703zzxJPDAa
YvGQVON7g70rDyt1vBHGThTRK4O4QABNOO2PT/hTHGAS/oVLGNLdBM9ywN5+oemS
gimNCuZ3+SfLQj30nTYpsEj8BriuayICt5gXQFH2qYBAFbe4x3K3vNHEoDGLoCyO
m3/f+ZxPMyivCm7Brzx6O9hyc6gkLGU9gv4CizGGN6DMkVGFRZ7ukKf+8MYsHnzz
zE0sJVWjDzScRjsZz1ncUMwDOvUvAMrK6IyIAbgA03YWsInmCdpyDEXb4Gtyhfru
S7Siy4WBb+DrVKI0Hl6IJvsTRISBm4aInQ5yUQFCCO5h1kqBt6zHY2WC+bR925Zk
BgWQsxQ6PrEWumMWirDV/QMi6uWa3Bn0WWnQKi+ZauaiSuVkEyykeBBj4v7l2cyN
NokjgKZ7ghuLyQ76OOE0ghiHxCgxEQxfz1Dz2QcphyuYwrReqS49ghzAblYbiQCM
B9YnqsGx3cZ5bhx5pY/xrQhmRixCucA80Ht7iD4AI+UevUWgE0o1Pxx+yY0/jZAE
dmRPh4Uu1g92nxGWLqspsvwc9jNIW1hfAcicn5wELPH9OGANPgicdClzmlWS2Z1l
SX9M8UrMn/I6jioLn5xCHTQtC+45tfEj891JsgpjYlsTa5upmZE2XF9UzH8H2CdV
zo+dYNs4jxOc9/wa+sohwFWfnRMYR+WUgcpX8hZ3OuNQANWVCFA1SmqES1tcsGfQ
9DTPP3Wz2A8dwpLIur5mx39RoLeqYBAvZb0bSt6e25PpRRnPBWALg7JhYENDHKBe
CLNDxlEqoGAh7fPVH4mVV+DoBsaqFC9tHl+sybcgwtBga7NKB6GTb3xlEbnPFCdf
hz8w6b76B9EGTVe8Q2N7k0868WtXMCRVY/Avtx7Ll4cPzp3UE1iCU4rw+JWECZ4z
LcahvuJWrNdkAi+sKvhgin3cHRrSlcLz93Q5zcWJWF7yieDdSY8SY93BamSdubrm
IjkWMZwAM1+FNNW/jUEHIdgN9Oq+tb1A6immqjQ+/ifHp3B6sosqK4jgbB+YDFVf
l9XR9wFcDcHggqen25KgNuVI7VcYVfzW/i4L+J/Rw2JDSYQF1KKx+zwr6ucWkW36
7Qhs6CIi2e3mrqEhu3q99gfedvooYoi4YV+6DHxXg4Xw+sMJQ2fTCkJpyzzjd6NW
o507uTlk7NKlJbcIvssWMxGuvNV6WNimQZ26zDi3gwu1A4eMoDR6bhYub/xBjuHG
Xu0+4ilfOtZMh3/XMitXUY94GrOuKV0aUFO3WYBviXhPTeGfauZA0NfJnmp4eMHW
1lubJWzAhZnFs5vKqqQALe5kdjrNkdvxzXqsz4GlUwRhEu+YQzJpW3AogmEK0KnP
EYkLiBeIR9rBUmIEEqQkDG2+EPCrshlNFfJgI0opF7guHLlCskBtKJvOlex7hh78
hDXs9D44cksLz4piXIqC3J4YYdO4TcPQgloAhchjqYJCF/Z02M6vBYr5L6mQpHdd
G0v/dqavifMr6ZlLgQoV3c3hYPjtvNv47tckHjgLvNP81S5Opf6+E9ytYj6BbASY
yKlFgLSagr0qemjN2P8bFZyurD0QlMxVjQ+GNh2Zlv+fekfnCaYgBMp7EZPBYK7y
HSZfsdtyrMHn5wEE9T+U5LC987SrxZpPIp6XiTa/M3TQVtCsZEI80j3rqtQS6qp/
9WjNKGxz4THb25TR8P0/82RYrTejBKTdiX6SzUIiLn2a+9DvJgbTLNd6AgWvpNlM
XgQQPeUSg+NQl6n92sjBryblKmSYWVoxFhISTVt7ZF4bcKYvLH0BiLhcoyzAwxqA
1khLRDFQyh6JpEvfCW6+i69YQN2xfRLQlgCHKCbx1juQUMxXmQKh8eFoFqfkTV9g
FJCJ4XM8PWyavOlsQk7ljmATCRIRhmGFbdm7PwnFnWcaEm/wyZ0Mq8FUXeKtjmSA
c0lMFO9GR9Om5Shg39UBx4Ni2vsJyksAZFpwyUhrgEVAz5o5HfWwp4fITMXf7CxJ
KUqQSDjjlAZbbacDTGMGlCb7T9Jt21usSxv5qkNwxtBocsYfH84eeLhlv7EoX6nm
hat55UBms8QVxL6q36NN62hOxufQP1YZnrJDZ968ZKYK4+5eougODKaKA8hIcpMA
h9NAc4UHtrUqfJtn2V86sbXfIcC4rB7To38GKsLMaDnfTkUfh7PT0Fvm3hSsW7yp
XLqtmwW6O0lBYesh1JV3YsA2k44njCAyF13OjHQgBehqEWueNjfVlnJa+NNQYcnM
YH3Bm23nqAtO8IExL4KCmuJf3O3FSir3shbT9yIwBxIe1lBH4aJR8VyLEm9glqal
+X+/m70qgYlNM7Lc7rb5k7Hk/ZirkhFjMMaepuNO7VgVg00ZQQGmCMRnYYJl+5W3
2dNfLrQD2SlfMsVM8xVuF0zPCOpK4+clLOP/7T1uNABSrqSh6cAtZK2bHS2B51gw
CoHZ7VqYT8GvrPq4THYxgrT3HdR7qQrL5y4TPjrx1qsObzuRJOeQAsTb207s8bHE
it76Zz3D2K99q9RFFBTdAnkLYcrTz9D06xytPjjLP1YM0hSEvmMKuZTofy7MNTAx
EzdQBtJJeGxZzkHFopNP+QxQEI8Bxz660gzsHpW/pjd6rKuIySZLyTaWxS5ev1kq
m0bC660tOba7hxJwVhoCbBSQpOaooOp5nu8OjRSf9UHYNEl+f4fRB4zPpYZoMiWq
Zxj+qUC8tG/SXyOuNuxqQ3hZTrfNmX/JfwCSraHErSyDupXaan+iKXvgRxU9V+sV
yzO3PKKRJh/I4IRSWOzP+0Q4iOltNQIRx3w/qp3drj4bYmfMKPORiOKLI/UmI2fq
9saSjm81h1u/Q0pMb0gMjp9E47fBprN8ELL4Kg6J7u1W1FCLsGwO+9P+UD2yVk4w
1+bYJqpNY8ZbaSP0p6APkL7l7xCzODBb8rXyBFpBil2FzwWXBY5eAjkdX08Up8J5
iikpTpMeLbJAXxleHHdVJQxMUo49/+lvxUXVo0dOd+Z9JeB4l72WQEvvSmXj9pnm
MOHvGTUX304hL2UkSfo6K3j1fB8YYAkgP8Ew8FKWBGEgb4rYJOA77KFiwTbrnDFw
dVbc4BvgMPHaYuNbaBaa9wnT2zk/OutljhPLtN4spToncA940mjbnbcVmYQJFODn
rO9aehVSEsy4nrr0RSZFkGxVMC+Gqs0ejbCvrobla5oNaa82PyOr3mBhXAiFJRzX
052NXepGK2lDTIrFgIEPcnlCQ4PjJkNozmVSFT4MStxs6+gymF8AVeT+xhTj/kv/
IomxP5yOxE+A93J36Qi5eqTFiEUCsYuCktvJys65gd3E/5aPsTbG6hWuZKgYzzbW
8Z5+98ckMsyuIxJU6fQr0EemM3hAPcu0CSxzPSE+AD14yQlQat1eexYGi2D5zVXQ
SQ0C0TBcRN6EHuzv4cCIv8cIO52bW7ytOYTMCmZyASvWv7dvmJm2YvuyKdECdYK4
iTzBn7UZITw6F36vWcotlarVhYPQx6ZeJ8Ciw5e6EhJKSo/4kU+zgDh4xgsMnGfA
Z5budr9ULQZnXc+kVyMFNxwNg5RSyoO/OSOfeC+c3CB/nDItCQPYkbJjX/q9bNsi
+DuOz0uPHLKiZZLMfy8yKeXDUOS+GkoMFMD1TrveJ07qf7ZgPKrkPggJKCyq21jb
fDCV0prfZVsl2ihnjKftg355h+F/oAsTY+BUOQvoE3PRZH6zq8ebevkRBSdK8hac
mdz9i1oSi8cC6dBzbrtq8lWoIE97NNLINfiG5tLWTt8mTYn2KejnE1oy5CMKcFFI
XC421VEhlpetfL0NAOoMFwYiTTZZTZr1KstTrFcPKmLypN4GE2ahXvd1NWPPTVJA
TjWkfL3BrWnujOx6W4is30GGKbs7P1oZz7k67SD+ZTnGbVy5XzP9GQ00f2Y4rsV2
oUDEu8zxbXHW4XJdaDaZ6uUZqejk0igKErnUWRqBmrRKwBrV1I+Uw7wUGrWsGNSJ
OF3WIkxLvoa8UTx3BYLLBNy2wEv2H2YeWsYdaJYZuxhxheF9rlXpG8mYPQFjOsxz
7PHoMHMYGkvdBIS7Xhhiy6kc4eH0yVIy/n5QKVnQO+H/wUcX+JZ4Jdfp2yQ0rbHT
I2zPZk0z5H51ls4htRgHxpoPzd5eI1qgVEfFrthBpI3z8BY3vVAVOZjItKIkA/JX
AcRsXp8amc1kD5NM5fywuqlqv4y55qWTUWa8f3GDBlaCHhdyZ+kwHJP2tSyHCJZ3
vKu8agEsUR3PTdYCSojIzyUqz2wH54uZ87QLWQSkjvXDXncU9T4Q9Z/TMcg5Fkjc
lQAxXHy8WlXNvEXubsBB1cubLQcgig6sb0HRMNtsKcdunZhYHsrAKYqN6dF9Qmx2
Ep/M7qmZNfThjj4HqTl6UiYQyH3zMqsTcDeueCw+jCKV0viWXRTqjYuKPV6JisDi
IKs9w3jMI5f2ygxnzwcvu0Ml1TZGdpBoswQ9TnCdETpbfvMmGVa6PsscARH/sEKW
adYPExe+Umuac4dg6VjHes1zGRd2EPRKVvmPXydPhYYC8wI8e06WvGAmNWezpKKh
uLz+p0kDCWisWuQJdYKTF6s+VGxVeBSUggPfePHqLa4hklW17j4VQPj/Og1ZS08U
UX52kmMQw+1F9K40ENohoPV15hgIEOg4+RH80lZoDyviB0hCxKSuWb8Nr9CID2dt
xdfI7M/nNUMzADcmDAV2atq30lXyN02VxC2N1N6vcsS0e454JH37Gd/YuR/qa1+g
sx25mvrYIYp0dX3PgCbjSs0CkAwRoDT2P8ZKfRn9xnWJ89CmM4AP29NMzbQvpzyU
93gFXRvvyHJ/HtNs9x6LvA1qDvXmYVt2V1w9nSlrAL6zf8QB9xzPBsLp1/dYBLF/
6gHbzcxuHaaV7rKMg7MOz4utMec37jdwd4l5YFh6w/f2XAUg/d/O91T9okKkEMUK
r4L3wB17h9aJWCzCQn002uGyYSKn4tzWYbm94apyPtYt9hHs+K12QFaSYYSZbsxo
PuDasA+sOinIS1AbJCarbLcQe7ytLw0k61A+F64PLY448uO9cwczFhib9yuc+EzJ
k7M3GE3TjJ/vwVdAh6XOiqR/r/gdnX95Q+0ERrs1JLVjB7LDeyTO2mCPQzUCQNj/
TT4OF0jGvNUbkcoOPcpS5JVmD9HXFBDoxdy8SAg0yUoXbGgS0YN6E7aJE5sYgGoB
+GojV1o8NuO92w2nW98EUrM0R3wHifM4pFEJRA176F1qf7askREGEtStfc2DmeAA
+paoXhrU7BRcS9iu7pD9p8Gi/ZzPza4ZhMDeHSJ8ZEqJwv+f1VdQG/NHNvE6MXhy
tpxYo1LVYcBN1zoFOveVrvMnBJhjcGjdowwLRZCVxRrWOggkRFP2KtzAxnaIHK/I
sHANqo53yz5ZxByU1mSQV1A7odO6U+rtec8G3upeb06iQVrEZH6cE98H3p8OpBav
WNNOAN4JZ+NGoNACp/3MGK8onVB8n04lVrwM44U2UKvlMhQosOS1his05up5CJ+u
ZRHDMcXtwGfLF+6OjBQMTMuRDlOpiA4t3ggzpFaj+J+2+NfouHEhhgvNpxpKjIng
pi3pOEvv7Tlu08KCM3UAQ5IDjXZa+9zgAjdZRkWj6T0fbtLjHhskcCp6LBHmyDsv
/Fw+TDmx+yXtxFEGHENqWjBeq1j61xD2BJQdGn3dXxn+ioaNa37DXOtrA3/n6wrg
b5dvgXzraXqyAztDLKizp9ArcFcU6qvA8bU3zokFyL82BA0YwV/AvW38oKe9tdof
UighSCvwQELmTJBFu1cZ0STnOb3R0JSRV2ANd8KRcF008KODuZRqtxQkzIacIdI2
liRNfrE36JClBFs/sDzH5G7QOK5LThhwjNPB3Rs9CWzoeTQI1rgk8AZ1pZadTQYj
30iXQZZEl7xSZrGzRcjMV4kZ9D59v5nmTyzFdvTGf0n0myr4CPy0Y0ukrfYhLigE
eyipmLDuY25sMqkv93GIHCTTO3NWFkaPRRvrNGbiZFwPYhrzJh1E6CUbmIBQSath
qAjvu2WaPZPPAntkwl72ZZnQLx5PmYuaSMcaFFS5T0oPd4UJDDAfgSU/zEXHlnGz
Yz16+W6lP6vZ+xSKKo+ywww2JiqLMAgul3KKGTMQZf89b4wGOTImUt7DJ3lalJIl
GPwTxOkzlQc0QPwj8cBOcqPSt9bcFg+VrrUU1FTAqseLj19VJa5Swqty2y5d2KlM
Gta0TM8UXsj/xoNZaRlEN+q8qvInF5yG7kKrGziLaTCBqWiohSuTTQP1CIIuicG9
rzXTEPJjf0hiRdNvm7G/eZK3xPJgfVsoF5DZOfreXLqB6tFnKdgZBm6hBG42TU/e
tKqmirc6ngJMO9VutShd/7M1qiqNihsnRnZL2IVTi3armnd0p/4lB5NCuzXl3+X1
iu5CNKdhOQqtd2Czvfo2aO2JKZaYAez+oKzbuaEQbFgUNIbrjOE0qJop3eJul4HJ
CB2NT+tIruDUkoOjT8svcDzYW3WQpfRX7kPWY2r2Zj1oq0I1dWLd+/W0G7PZ+hTQ
sd5TiTEpGvE9O2poAawrmh6fZa2/ZtBZ+RG8+kMwMEH4ce6j6Ba5mPYHpV24JPXy
ufj79+mE030q4tEsXswKt9zknacYtDN8Sj+Ust5SKDyxB9IAap28G6e5dYOaVLbA
MbhcIc1u+YFZZVRA11fvQ+VPU4X+/OnIS9axoLs9+gtzFwxm2o51EvcvHsn7TUFM
OPe30gc5UL8lw1bTUqLJDsOqM9c0hVotqVgEmpJFvtBCVvxHa3lo0iaXGjhvRfk1
PvLIhRokwQO5AlAW+p7ADskBhSiRMBzusHIhrnBYFPg47nmyHvZuZd4D/Ci7i4gP
q7mh9le+1+k9FbKz3wZ8rD8vWiLG1/PcGcJvCIcuLrY6M0EEe4yPS+5sySKplhcL
Nkf4joBdYyt6bd/ELZ4AhLG8lNmjel1RrHLZ7gmjEpDtBkkRAM/4Wtjc8YgY2yOa
5xdnJtISQXKTVDUWd7tnndyjYbukDJwhEGzrqOqgXwafktIARmg4G8V7PHiHYfoE
ZNAf8QWeTZLMLMRMynGCKsDI96GP9KqigfkWR98HuAnRlBpQnIdyVPilFk8ohGxS
cqo1lxnxZfJ+4U+2Zo52mNdEtFhTLJMpUGj+Xaibxt9iPW63fMUUohDlA1vpdLj9
lxMvLmMtF23I9LsT1Gu4TtLfmogQ0H7iPOPMRjgw1w2eOhLHkXVal1moFdT440H5
w39m71BY9ohwkcZF6cmm8vL9bXygguSufLe7QE45qoPmy1gT3uwSPcBdY7BaFKsk
aSfGMuaQVrAiIxpCJ7UL8eiGkedV1iCUmLjONBnS7t07twdq6+IAm9vhknO1GjjH
iFcWsG5PAYeLt5dL/+dN9P5366QHY7NAuXCsRSmx2Mo70mz4Huxj9Car76SVuV8X
oT7ALuCy91kdvpDLRy0BVJ6qjQ4MCoDirWnQVGpO4iEG/4Tp+wt4LXMLma6Ti1iR
4fAwYVf5iPfSsHM1bc0gwJqKVCbqXheoJXvXFmKrR0e/8k/uSGQW+BdxS/7hIJul
vbfJfAkanhwtPBkFJRwC3K99Gr37YvctVtIRqzVRzk/OsHMbd5suoBrhHmDrhH6K
zk5KEZmWK5RKXbSj6ZEuKWUvPqq06W6kZgw9Wyg4SBek8F2Hrm4+ORBGL5PerxOq
PQdSLphamJzShn/niTYafhiTFWn14kR8fo1qcamHBnT3ZRpp4btlw2I4l0eZfwFi
+a/2cpskWyZJEzeOtSbSOfNCFQyqBmVwvTsRF84FHzJRKWAIF9jdwo+KmsVlqMG0
vzx0Pwz6tm0IyGz2GYeFwVNxK+7YhiFB2lyfz/ekyghK9fyxbPm7gZkIV3ZsFwws
2FwnItBGHu1tESZ5Z3yYFdbICesD4l5KOwLZ+5XbWd39mDOpKq+vMmt2YdmynCYw
5y74cyZuTG/cKKow/VEV8KkynXDJkFYS+baeYLXD/7I7zmmt18xcW+tqqj8b5f4+
/e0TqOmjSPbiURbxNuKsOwnVXhVFeadKZlXv9Px2YSmRilyJNCJZPXHt3qTzGfq9
lH4XlVcGCaIoTv9h/WSFQx/MfsLlgAc8HulGMPXZyG63VvR3IYfAplT0mqihJrtW
zimEIO/0sckPmjw0Sq0S+TofqAa6vUSKO+4WGF0LesuMhHHLCKz495Gyt6PylaoP
uVkE+gqmGOwwDnlZXE2eK8AKqkVbo7JrtLRSitEUIgfundzn+RzRdm5GzQ6Vw3cq
sSSl/d1bIgidT5Ht4OskR7EtWiDfJu9WK+tnGIVb1aKEfKV3S9zwDZLzmHoorWCT
OLUiHuuCX2RXuUYN0ea0BFkCQvf7Z5AAHfOGehlhDENMyUZLdXKmwYvfflU+WKJT
2xPcXA8ekVhjk/vToI41ODkx4kjkRxMmd91oI294hgCe1VdcowNVbrLviSiLqJrK
T069ALlTNWS9pyYKB6T0TL2IpUf2142CW1M7SyvN/pBNloB4FCHZlZqcxGbZ5E+W
dtucPcBghdn5fTvrfTBAIFCL1zyfKagkhubf2743KZhuN/aVBIO8qQQvDXOoW7c9
0uzu40c/LqW0NI7DFotx4gaMF43aH0z2ZHCGHFOyR0ewyAziDfssn1QUa1NWFpET
WUX+XfSvDGtjOli4RWacr8gZTskaoBN6WpK1D+2w6I5LcEzwc8LEhyiB8G3HYwk/
Ee+IQTbUlQABi1HNg8Zb1TxAgkFDWvEr2Si+Xl2+Tbo2R7RHCioTLwh2D11/Wz/0
rh7qj4AU5/o3QY4eEdD9pZQZtiX+/fY3OqygPdkZMAkTycaLhBuBHAzFNDTsGFHU
4wHdB6uZhH/41NooLy6k4U4XKeAYJp1/Aexe1uOh4svjNBQtCE+LGsNpXlGgSixH
N+IfF8EOBsZrnOBj/CeIJvk98or2z/+npVZ0Cbb/hL3MLgNNAUykIdJ8/alE78KE
x91tKP2FcfcCYPVOpEf2JkYqVg/u75RcAqm4M1bm71ieVrUCF4Zw57Hb+F6fSnA0
dhYJ2xV/7VulUpNDfieSYeNtObECitBkA3n+4MLDQ+okKfOHlPVs676+IbXsuKyJ
JrzT1aTRjiu6vkC0PT4rc/dJ8dDxRv8aMft/DV0UOs0cyJs7Nqo5QyEiuwXnerbd
6zrucUWNW17dO0NoZvciQjRIiRQkOBJZH02gfQVQVmhtzzqHcIPPoeEHNSWIkHJI
Qqs/Pk9sAV3+m+GBQCabmnedduIuNtb4cQeMockMyRM6fkPncAnzW1l1K7o0H7cP
PTWv4cptPSV2sKYRgBIh089RIgFu9PDo1B9vHsscz1DSnHXvNkL7YQ7AgGhwb1/q
Yirj1GYf/d1q6p0VbG5p9BIaPyq/DXWcyoFMzFgy5imbLUfHMzMI0xkKqM9ijuKK
1ptHglvOGvivxN0Py5zHp6HO3sJrD6mcbrPcGWKA1XAxUxGpC6fUAUxyyjuhNwhC
226oUhYNQ79c2VakO/3kq2Y88ztwNZOxiNLq7lglKKVWCIdYxZ3Ce9J9Er7WpC7v
jwSF3OM+8MytfaXSkOEpLhQ5+DZj2yJb/TlqVnjymFfaZINLSp8zzEOoXYMq3nlC
UutppwqDtCO3CcfEgx1Z3yM34abAqH965qsYUNyCzrFUvykvXj9Iq0zbbGjFJqvq
BytusFOyRvvrJGF7Sk3reJR/uv3ar3PHQiX/iyBYCwYZKF7H33S1UJ6bwM5e4OtL
d0yBoUx516vqcmWfHByku2VeTyQU3ejBP4cI6l3j9+r4Oo0QctaTlNEYQNzT2M0q
Ev4DganEGl0ZF64gxKJ20UxKpC2b7zY11fBJK5X149+Qf8BXuWF0tDEmI7hm778Y
hBYKKWLI5In6uc0XbfdyMtDmDyqYpqTx1CItFS4Sc38iDqeRG5kiSkJGH0M7OnFk
bwtJ0Xb6yPjLE5vJl0iMaLrRjKKKjWdDxoxDMyUSAUsza8kuTgpYTZheb4DJsRDk
Gfw+3OHZcVgNMDHdoHBH76/FdvfcseEDxfZD2rzjewrxcbg4MUuE+sXnzONX6XSU
q2D1j9MvO/6pb4at+/3x3SmIIXbvpQ7uaixrfvV6uRqswgQs/53dV+jAMUsK4jQO
Oy/0BL9OPzOrjH2l5Damb5CrPIBJTg4htCZ21VDrfI2sKLq1aourAPDKaxv3BR6C
+7XpfIcMrS/xJrmzlFs1LCkEp5jx2r9WIuPRV0J+0avl7PtBC0bwCmN2f0LLl0vE
MvRLfpskX5bTbHdhmD6ZoXmjaAc8h/xqldVNXthwBwL7bGmZkekOF6/TnQHAw0by
LcX8JTSAb2mVKAoDvvsmrB199mSGiSqnc6OjT1oQFu3WuaOw3qpoKo/Q21ZHnLF9
5+e0zYDus/9Tj9usNEhUJBbWpplSDsdttRwSX1kEVWt2z9hUi7+i9nEosLXefmwz
nqbXfVGjf+DpZWUj3pseN+yDexjeuFLH99c5klAxQzbwcTIbeL1xWie5OwAU2Gs5
2YpwxQ/hDeoB4zSNv0gTLFcMCFn7g1q3vARZRcWSNWXmYfYeXFrhGNt52MKvfgp4
tB6J2XgNwaltFsx7nt1pJWBYVuswv3aUinF4T81o/WdYAQJ8jYV9RuwZ91x959za
AuHCIkA9XEsRlCJRO+ts/KM8dx/QsmaQqlNbUrWHYx6uCuad2K//uxtgp70OL/qX
4go3Gr/pp3eDvJxE+gLew9bAr2I07sSVZUFJ0/YcGxGdQGS+RRbuqG21nlohLrTj
J2leMjdv4ycxtKlDG1GVPoyNGSLH8BDBuvagqJXs5BzrpCMNF9zdIf/EOG/ySGC7
WObl1qpSzUHfoE84mzOOQE8Wq2DVk7BStRx6HH6CwG/LcdCfLATyh9Xe9I/eruJI
AFEQd+a3urLyEtxi4gY6uCcdXjuFfdq9aDkLsQlrPtFv/a03Tei8xO2+Vu8MfgTO
BWrtXsrZyZgCbCFqhPoLElKeH85TtmnO1VWILccC1fzHfi5fA8HgbptZGvxdywNm
gMoiJ6/jpFspY+3MLRhDrXVbmsUpKLjXdjph70JkH6sr70FteazYLQaWw6e5VBQs
2uxvVHdnA8+dVxaoPLgs4XKt8x8IJCroPPM4gvV7hiBpcTk58fC0mSbACEuGFUzs
7jAF/+f5cE+nfnV/VebgoLcRJugqqaLd4tHHnZ+Oisu98hb5t4CJUdA2YEhbjmA9
/9FE6iDwr5INc59cEyrOOTU2GGM01+PtFydSB4qD5Z+hpBQjMEq4K/NZn+p1+Hlt
SYnjWh/P18EfN0ylfasgAzBitPxHQ/X3SLi+vmRDug5zvUfs3C1qhBKY/rXkzgcy
J4LVhRCg6gNCKknpidNlvafQu9Hzyw4wjCMIult8JpnP+98QDoVq90TXYSiGO89N
wLCNoo5sTLX37zYIrDrPXbMopGinXBDY36jpPTF7eg+cu1hi8q6R8/bRgelU8cuQ
oGiRwZ5bgIVFaOtJxjcfBrC4TuBUPaAzRycsHy4cHsPEwnD8MZY0rNU5+VSXm6mD
Tq2COVuMv6ndjGkDPtt+kCMKs8PUuLc0ZD4ZYIRYDIyNO8f7PbLUWV/bZ/AkaAcp
Y2hV9km/AuWSI6TlRD22yWL95bO3aSnvKWG/z90nBI+2KIcDrawRkOqW32In+352
7/rJVFht+mZK6MRVb2KSd/ZD10jYZB4yPK04LlCMZ94JeGSydSUk9A9tnz1Vi91m
5E7LU6WfCphb+UZYGGIZFpYyntSSrPKTWKvk6fUG+onwy+bHOASDSQdGSh/+qWXo
+J7Re1cClxEUDA4vdv8xTHHU+xu3V6rQRVWOoXVeyQKYq855267DVayNoAik2d/d
VXKmBn+fQxxroFBr5t543eGI+7V5xT/Cut5LYSzMTeH9dMgA/e6uLbkV5DPt12qt
ArmItWFb4qCQWQp4rUFVPWhX18CUY9rwEBglZ1/CVsQMTtifMKNjTUgWBw5rJn7g
8ND+GTcaKnwrStoQg5DgSQRHQg6443ueaavSyNQWXIUNrzMbYMZQSXx+9fjXzxE4
LnibZYEkMFOXmkXGzVRLPqmjG8FMbHPYkjaoOiU1mSoFMzcohu7MjCib8zpNgSoH
v8grMoHx0Tca0XBisrX/JzUNTUD/7FEWk3onNGnhLgu7ssis8hQjkL+taobih/wh
wyjsB/9WKJh2jTyP3+zH0wdYm9zNHJyQLShjmK9s2/kWA661ZWKx12Js0sfBpNyh
AobOluI940uHOplMTNhNGFjxleKax45L7qL3uYnD1LuJC+giGOHFS9NpI87K4754
pxnp+jCnuoSnTBgyB6h7IW5xi9Vn7dyuIns8NXFLhY+Z5asuQ5qpfCCuls9kdOCZ
TYBl2nJg7yjIGGg8bmSQeMruOisaYg4RmH2D4e0TYBVGZCIfEGaT/JreyG28gndC
Vjemm+4bXKumLFu7bCsTnnuVBMPIeslUY49YpIMIpAXe+mV52ETd5kTrlAyg6NNQ
Z0Y26p+4HaVrtukt3AkSgeKs/TVWZEuI6LUN5CrgPO/tscbCebqBJVHKMHkVnB9S
Eg5F3RBc+UlUZPqt518EMb6fpWOFZx5wfIP1Yux8yRmtTPj9asG/PJ9/tFR53wjH
NYLG20zqsTYwlZMGxqIGCNdxdP/1/2hAQhe79kkmXhu6edr3aRdizUAGkzX2Sy43
4PtXf8Qp4VO/oKAUxFtZWa2HtTg8ZTaBNaSqDGxzZLP4Ea3WfDyAmkJ9ljAL2i60
ZrjBlChJ2UjIPXC2MxaAu+mCyF4c7+Q8UMKS//5tj5uo6M2fUumigNwz4U3W5kE1
Pilfv2mCQZudatPBRWnxx6v7skjjOODCIvh0bKJtU2GwlXferzAXNwj/+QYniTZ1
xhFxD4p9A3qQ9IkgaJKdVm404JIZmxGSKT9ViSLg+7lcWEfd0fra1ismne4cRZYx
asuBKEki/UClZQlCxj/8qz5ffClJQwT6H/oaDLb7lFNylHE19VCSv7dAtiVx0Wib
lHdto/toVyGhNuAtyzifMDEryUUlMLz1GjJB3Jyu2WIStCo6ZtEcqHwee/7MQTSR
PZc80LrsFI1wT9X0IXgNeS3PonOtfgPgAayNeqe/s4ga5yo2cmfxIcoemNnhZjnY
2adl/ZlfR6eOAar5CABuNYIEJnOorqxecnNQkV0Ils+UKOqTDoRfZonKYXT2igbu
y5A5czw5N+osIcS2tXMcYopv4NLE3PVnHmE7YUM+ZN1Nnl85ULbd5UKr3OYuHH/w
uq7zjA0TlgGq0U2DOlK12YgKCtLzdp6dx++UgPv+s1LpR6GvGjBbQb3gZaeSAXle
TOuz8wt7HWze0u1h5kafv2x/3BOGO7tkZnBnXhSIEH9Zi/PIUHtPGX/yJujg/wvD
EtAogcXs801jcUMPdLnIlcsZWRsNiS0PMY8w1JPTEIZ0NTXi0w6+x7DT3QfXtIiO
yWJk+i24SEtlA4ZisPOuW5bHuIghePVlGyJedXVMrmx7WTJxAzvHch6qMpRx3x6a
fdgqhyL2V5YQ1zoAGabMU3gFEUOST/ZbFjt3QnrbEYQJ+2sldtQlmPfQ7mqZnUua
ESa2qQYly0VCNlHG9IQNeHS6OJoQBX3BqAzWD+sBXmgRu4wEZNOo1CpxzuxRECBX
wBzAwu6fWGiiU7Plsdlc/IMRZhrm85L4X2pYL1S+iSD7ZODhBX966M1jUl9gd8yV
6LQNSEsEzQRujtWK33IZcHRh6IU+VaOYjhpOFljyTBDkygKfYNPo20bm+yDkp6g0
vrTmdv+9HpfHFouPAXGV51/JfWTozDMFRELV3zOLtLSMpmu+0p5jgQV7V48mWF6E
3xjDne0qtAzvfFoFPB892lJtd4QSlxBszgfPOq7G4Rozdn0sGmCqX7NYBGC+htMB
oIJ7mw2VfpQCEE2iWL8U2ZTdRCe4JOqq/syQ08QZeyatKcwNsjUmSISzWBhrMZJ+
9pAZzPadrWLlbc0/ao2H/5AqUR4fhEOQud7vEe2O8aN8neaSzWf/BBnLEZarT+0M
2yd8vcJ+euEcZNBdpepFwlahlGHN+pSQIcSo1H17r2eHSsyK4myChhNZCcmiqlSF
yI6cY1XgpmZxYrLEihdZp9eWyiDnstOgaQyDdaI2SIcNpHYYBxXhdhljdyatM54t
TMUUZkdycm0XiD0xbEwXXHzjNuBWsVCgqQzu2qRT3XaXgab3mmBOh7220/F/A9AA
WLMvQ8HvAXQRDadtwRkcUK6yVMp6D8sfQz71HUXmsOO/LO8E+x6BK/TFEtACPbHr
kO2V58BTht3aLLsV7S+qAKHx02/K7+A/HbkFCZg++zv2vsQJGFfK0OIe/boJCz3F
665zxg0XC7BvfPzeHT9FkoTmlThVM0yg++ZaIBzK6pJ3wREjsviTwOO7F1sJCJbt
D3d/rDD97MheOl8MOLPQjrvcCe/7BnUsHgfxyMMGGRT3xp04mRrrpLlt9e6vkkzE
GSlzwEUTFjpnold6HoiMO7fB1EpQTALna1545izOZTWe+fpydgV6AoM3O7++qZdD
51sjHLr7PCPxPMFosyt6myuTOc7A8hJMt+RTPUepmirvVuW0JkKOftpu8/ZgmnfQ
jrMdsuKIZkvd0ViLTfnd4yIoAoX9ApmhVZml6Q3ijpwuXCAcAwrArnxp7tg5n17R
mLM2zXLQ/3+VJyDqJHeTajgf6X7uLH36+f2Ydqh7/vGR3e/PTnFZYANlrJIm5Zf2
I5buEMmBv99G7ryLTRIB3gXft/nxd3ALvyO2hm6j7nnix67JN7XsBlaSv9aUrz61
cg5frqxOXVsg6ipRkJ3jZv53AaqZxGAM4wBYOnTR+K2znBUQ4EFARXXlE63IB+Bx
Fab18t/pNzZLKcsixbwOn/v0JkhBvcIUZkBBZTBFnxr/SajOnaDzFu6lFGcDWymN
qQ9nxQEv9wfzjgMoZaz4BVmBKbRH2MGaz1hhuAKYvvawnCl2NC8qeETmfZVBm0sW
6Hl8eK/c1IUDspksq1uNycPe5eqZrdQKvaL3rQIomMxrpQw/c4gx2dRkxPHmmRpN
vm1cpNMbU1B7tJlWCn7qcGHq5GaqTvOmzO4B9C0KUE0EDFNHUcavOl3aTSpGVwvo
Umg9CCPNOPWfi5RAUsc2EkjFFlKbWWauH2ILCJ5EFRXd5QXEIcEGUnZkcQnzvdvT
grDOU+sYE2mOBduDEoZ8n0kTvJR6pzFFDC43hMmLK7Fk0gyzw8fNoHBbC89LAGoF
OD3uYP6X0KypYhBP7hO8CAtN8NdjfSp0M4JT/h/UN78RnMZufS2wb/EG8qHDn9uB
OhOnGgiAYMt9ZEd5lW+rGsrT2Q0tGwK0rlloFGaMMb8X6hPQHA9WzKy/e6ZOTz4p
9w4Lw5tXj5F/9omfuXGlC2jHlw5vQgjaeIJCXrblIiZXBPhHpSSzz+LX+f685TDZ
VMuIjK74IcwTr1nTBKyhVjWQndMdBk2jDRo/LzckajAzbyOTH3bWJOeGDcrRs8K0
sQA7oiqF/0qE95hld0jLRvhMMSioFL+7LBW+GrGUaeUMMTnyJvfLhM6mpXHeemm9
t8T1G7fFn0q2Ci6YVHKdj0lvqRSXwqz8m51j/jc9YZ1U+YaIhEQCmtRugrpVwHsO
pbBMoZmpU3Pa7QDI9zLLKXQWIJdfN/oDa5RQ4qlj77bcJfvcddwJTNFrAX2jAULq
U0leR5NFmIfDMHUDEx1iapf8POFDkRKTS1hg76k27VSwkwUNi4fbjffSjUWXz7Jn
gRd9C9r3FkxCserQ4qaecO0i19lC/wOWQSocTPGR3MnKUjKgimL3VKL9Qxq4jSfd
n35/rhT9gGjp4WGnWSoPrGjfPsm7pLDu/ZlDnZDeoWhmJDXxYSI57a0Otg8CjuXz
rtJVTvxv8np83I9d3SaKW45ehWzPoH9fjxOMueYMM1kPD9N8d6t2PdbkLGe3pTNP
tz3Ip0TUkV/ByNTQp8UFc1oK+VyncC+zAZjlISzv5w2km3Nez5l1PmPXRbXpfHoR
ynxZ1Ij5/Pnf3ZbyCxlSA7IJscoYKXD5i5z8ycXJ52wrPrnvGxchVnGWhpqus3VR
gLQ5b/vNry/6mTHSbcbdbmDe5O+OqjqepfaOAdLax0++r3nEhRMvMUx8GAetcRtZ
J8OfWA/fipIwb/EHO9+HeLIzasELLHkYqXx0H87fT8LYI4gDyOzP8tnhPphU2jWM
dlFj//mZkoPr9CEt+wcQ/12EcC5sfy9+TpoI/yVFyYeRBPeSbLmJjQAHx5Tc42NM
blbVP0p74aZhE96gePcmYm/+O2O1Ivd3BA7COGzDE702qyMCYX/Kie9srMZRlmkT
Gbj1xx3EZjD/v/liC8PZVewSwst0/ZyfwmO+dunsFbGKIcHpIMa31elUbEcAay87
3Ef6zTJl/z4UImkfm/WHOUGaJvpMW10bTUeM+QCBRlA98HkkvV0urLXazG+4vTG8
5giauAtvcmwX5opZjnEYHFLzVlNd53a5VDHadRFGGO7W7sbkkuCNbv1b5SBjxN6b
8WB8Uta3onk/XM6ht6Ij6EGFMNYkN+h9EQaLgzZhU0PHD8k7m7+I5JXE/dWhqdNA
R2xmTvAzzg+NrYySw/NPcrKvboAzVT/FSVbqWxreS7AEp/z5xzTvoyiAJEoW9vBY
TkS2POG1vqTfR+qF5gnoikJHLmvE7+RhBMkP+zoS8juX78cT7RTebRekXrhr7EyU
jiFBdqFZrOM5vdINrYbj2EkVUznTZpVPX/0R5Qbbmaux7SwKKq8DCf9u/JR63hNu
C0Kmc9ozD+PcLpx9/z2wxKCS2XbEAyevOF/ESg+dmEyWz223oLLE/uCMicDI9QW6
jZl5H73OMlfumCLbFBRBJ0G3HcuLyg2L/EvStBU190dTEaV3WPSwkbuYDJeXOSdq
mgOdNRcn1NDBnfksTlZCbbue57ZNrmVdzl6AmzHA95HJXKGYmB5KL0Spppx6WAHp
8PjyI+9pGbJZQ5JfEAxMqdYUhImp6n5/nrPw52gvElmoId7oIPBzj5mVqRmpQMCh
vyVraAJr5xGJ2/vuzEhOJ4LKaapN+vtCPbyh3UBePgZspCG3rUbP59iHY3nJzH2Z
I88W+NGLO5UsWSD6ZOKsgWVc1UZAf9xG3xzcLjp504IFaXYhzsyXpsn0DGO69HoV
OSZFzkIONS9Mx6xanptisI1QoJAbe5z6SecUPlIuM8/1jBLY+kfs3b3S9bbPp9F0
2QerGSm9k/ukbo9s+ECEL8VZFBbMyUrXnbZ1AAtEjfbbzodPEbJWu4ELWj4pedXm
DKMVZJYmzyHgkz9AhRVT1H1pic2WxHIr8KHJYZz9jT9W+F0c1C2vMASzc4LDafiE
8T6aMoksZkpK2OUHQ9InpRfUZozSxLTN+0dKqwddPl3oMtaCNGULqrY7AU+m9lbQ
aPBYpK6QaRr56bdYUCwHGchjdr83zHkqYqrZ2MnqHxHwd4d8GbHfLiq4TKo7GXBI
kRfJ8ozcNxvQv/AXlvrL/6GVD7aPPh4OUc8abehXbNFv3rRcWCY+F7w9oDIKnTgD
RrggJuM3ag06Rspt+06mvpHr/e5EvqLyboCzb3B+mktaAaWh1QRtT+9rrUlc7N9i
WWP2yYjCPxgZjl13SyGynSA84EQvboGhOFgh7bCFUK/qkAqTvHCb6Y/XNl3gAFVw
g/NgbfHFbI61cTk8xCoC8gccmBjapnhQvdZTQ3gbuQ4OOBJrUFha7jo1KHOEdEd4
BlbPHubJ7pD9+YK5MLb1a8OpHtfFyE7+wq4F+K5MATqcktvpT6NWI9afbapvM6it
338k/I2UPJHEKs6y+B/lAgraGQRN661anbL5H10CljVamYxpglc3mRM+we20KPC2
YBiEa86d9YMKkEyw2THYVsdnHN1niYVlIJ2SZzGsE0cqQ6NEWFM/v+iwSua+qCYU
5lo1AValTqpkRnVcQhggWq8XcN1TeV84/s6f6O3rNPyc4KPhrrhufotOLKCrrI7d
XvwrpL3xTdeqxzehlRpD69GGAud1+lYhf8N2K6QycQXzCLxP4NG/R22oSleRpvIT
kH+91vwUrqh0D+Wlq3GAIfw1l++7ruTvzahbdSYwp7gL3WpLD1PVRg7eq6s9WC6G
L8WMiD2nXm/C+LvX6Wd17w66azQlR+z4UCfvUEQsYMO2gkEXRx2xXTY9fk9CYacP
g41QskTePSjwf/ZEbkt4yQFlPqairY6XTkyguLbEkIc1DAoEDFgehKEn+JCQNvSy
tSqZkdfs4ALNOrfYA0j/JPPItFjlQJaZwuKvG3WQuIuXbu7pXrWYDlUB5PMORHJr
EMq1lUYN2wFDoeheBGNU/RhusI9uT+OhfWBrS8Se+RS8rewE/qcw38iyBl2brFg1
8AMsHpRO3pR+QUcYwEleSdRheFtwvLqFYrVRDFOFUH5mlIFPHpZUfJoG6iBbcwT4
NTTPpYZnhkcQvHewE43dDEJJvOQNNsKxWWb9AatsNuLRY3f4n72VSZJTqlfNNxYt
6pmmxlQAD95pdi7utqKNZDu2ZhUbSE1SXxNyVgtWNJgo6agpq7GTdEY0pQBfSU+d
cxNsrXklbgmV88PebhR2CHvwyE1zWd423PRkPt4ioYJjEDQ9hqzvi3I2L2eJKT9x
ko/bwT3GRvq5cQLWWGEBFVJ40CK2FylC0RDpLWFI1svYtSulz/YUzSI0bqgrSfA7
oDNm9dwe8pbLhWjXZnO2dQngaHaHQNsQcGtrIGQ7SVd619AFIHPmb5JvElX0Uz2U
MEEkiRTcNPyjbJru00Gcr/yCzxukkiVmsz1yYs5VSISZ8ZEoVrvREW6aQ0ZJheG5
vbxW3tX8p9dlQl4NiMne7IzVh+x2B/I6gMX9aHzHgWEthOD6ufHa1/PUb9tcihfg
xEFMwxOkbqZlzyMhXguVL8BMp24LneI0AnOqRGm149jpkgQAHaxYtpfs/wXBU15w
54BGCwoNmgLZHTzrq6UYY6IDCHWJ69mvL3anolVnRM7eL7ySaSjPx6caD7lZTyKY
GYuveL+ioYUoJUXp6CtajZm1GczYKhfz/yYKrqLfiY8PyajBs3PK9t/qFjeb24ir
R1paIfM25ibiqlM+zlYKn6vTwikt6ePhWGR8BgcWVUBZq37/KkeUfDNAe085QLLg
lp/WrNOIkIJjUWy6HiuexfqLygUmWTyzn64YnN8cYVMo8AHhQjfuEBO7/Xdk72Xl
j/9gptSvMASWDEWNCiQhhQN1nQ/kudYMDwtMKK/ubTq8jp63pi3xnV/AEbtYxMpi
FKc+ABCTYwutfiOX26r+sZJCsvwQ/KXn45pfJHEnWo6WBMiVzAjzBBq4wl0EmR4v
2wJvonnQ0k9VxShjkVOwx/rAMxTPvMqOPgwrIJ+7tlO4tK+t+20KwtcxihPJAqPA
DhWLqweCNQg8kPxJSuMO9bnIqsv0VQB3N5QsGqWvv0g1IU73VHuWPAfuHZWoiWyp
zVH5fZWXbh6eXyY2vVCEfckuRRCziH6lintj6dk+ufe5b96I4Mo7GifsdtndlTmm
hry/v6Mg8hCOvE8mkY+YgsKqjvVBL6IXGsQFwNqfb1NOdw7bMkS+NFgf3tZm5kWL
bU1ew9ORlHTSYLZ8tW3N42N3Y41YdceLrdbVJgzIJdJzbb45GyKGdsjneDwDmi6N
pieaiU5vY26+SY+RPG2LQMFewr6OgtQzM70tlb4HGW169hraTr3YAkdZxkWba1qO
lTiQXxegi41Khprlxv/vfBOVTNVBbwtzp3xUC/9eSQB6BhgzAPGZp4hZG9L6CxPx
WMif+d76kTK5O4eCO+HF7Vjq6f0GKpxKJVKTWnHk+dA7KOsdeU9ResktIe5SvZ7k
2FPyaCsqqwd6toi4PvYfhqoBtfdeYhlkv7IX6IFJYF2CXpTnXBcCsU0GJatpO8pT
6hd6j1fgcw5VwH4WAkWPkuX20gOlbo6sCREViQQ+9QfMukw0BeglIZ+Wx1//TzRG
rgmavqu6HQlJinr7OQn7zwIeFAQisngF9Ni5sX9gq4j3ZQDUsvUDFEM/n+vTjtBU
462T2fae4uNGCsJJQV1QWri4JdUg1dFBOz9s+xxvBaPGayAKzYj9agrkCHdTRtik
cT6jezFnsi1yHEv5zAYpnQadHogNGJR5EOAOdzncrZWSUoinFjqDL6iVz+9HSI+M
cRJ+yVIaDf9I/yj6G0IRm1kFB3/nPBmK9uwE84P1PH9bliBtedynQ53d0k1eLPYD
UUe8xCRCR/Pi3z5ppPW9NMQnRs2w5a/FP7itrlO5+0NtVB9j1OtuTkUshE9zLUa1
X0QzHVqya/zhAqnr+mrD1KLgIuOC17OCti7I4MrVmzttSTE3qTD9FIpUJsXmx6l+
2nA2k9oRq/Nt2mNY66rHscDiHaxdmZtwnJuvdsyjZvGL2btR/ire1sr6n0f90RWQ
RM6zcN6pHWbz9HnD2eGnTBWjQ+xhIrOGCjnlv/JhGp8P5p9izgsWkjHNYqTu6i9d
vsX6E+xohd6WyLxfd1ICeSy7pNmIoZAnf0imOA5zFUxQ7qWRSxkM8ipbFubdi0iW
uN9Ab/mB0QU5RRyletLZaonlm8slDsImTgUbh3Db9Nq74Z7Y8WdiR/WuzEuYU6nn
7W8g9RJWjIEuhakphVQ/XjuGiR5sv53HOkxhmejt72liGDwjDUxNw05GNtgQzUUB
vRyT8VhOb7fw5KlRxjMLuH3gH6ZJ632sZ7TVXXwZxSFdxgA0gSSRf6fO+w25Y6M+
BSBi+kx7OqVzkWG3/9OYptgPWTnItT7QiOSUK8f6BjF3bgdIicxxjQ/H2RM5w7bM
TrEdoDPRRmJ6heSuNyPlXEwTU6v5C3k4JvGzIN0AIaqubhaGk32O+irpZbIXvY6o
8v6yfl+HFgenxvsiaKm4Kc03jpaCxLXSHkkqNSs7Kc8zjILEkFdgBh/a+L7cOxwh
CuxQiIRbgAJabcZP//DddNZb7PAjjhyr2QYKd7T0SGs9pRqRKFhzKPrkNPTqDHbb
IqyzKGp74jg8yMiqwc2O7CTAXQ0fixe4Wb3V+nFYL+El9RmKqPdI9oyOIjYNckso
f1j7Y7kzaMo9f3c1GMSzRsd0d7gQolMDNBiUYfmq0HiUTYlHZj7Z1uood2TkrG6L
vvpuxh3QubGYitMunxye1dZxlcR39NqT8qBoKETVyUTxSZ6heTBz9BeUw8YWno/Q
Ys2Y1ZEf6k80r4qlLltEW/8f/lq892F5rqJdvhZLPjbIIxktSQFEyM0B8p96k0sA
kp4HzrEvX2r32/hvsZibgsbX+xCNiohnwNK6+rHAaGhsmWVxI0J77IsNKvH8J3Go
1Q/SSK4tQd82W/bMlgVLDIPsE47DZfc7Z5JnTRB1/GnKBaDlIEVzWuqTTxS8RhY/
gZUyhJb2gUAeJSyugTF4U4QLhJBBAWOwhHpx0VYIGbtbvY3qpr+oGWSmlOArbdPM
F1qSCUXudE6bsxo+TOH/MfOFEprx7++mJnOyBB0VJMDVs00+4iqqkKUfkljyQ7nt
yaJgqhepCl8pWXVle2yTT7RhpCLbTuZpYDEgCY5bWKg6aMxHFcSN5d0tzbF856EG
JDdMOGJ9ctBvnd+wyMQZvipubZCZ+IoZv+QUho0d59mPlsQfGFUriozRSp56aLOY
DEvldhaRHcZjOO/6x90JjZUSmiJygOuwKknb5VkrjOVwNV5O1QQkwU8QRPmf18wy
wzs9/vfBZ9B4Wn9niPlRE5Yr8Y/Y+QNlCtA0dONSb7Ac2f/Um3J+PJ4XkJP5MpOS
dngHKKVXYq9koI6O3q1GV5H8ScLiM+R3Ml1pXRv2FTDyC554XJkljCCNCGzEpYIg
HK1VEk5IP3g9baCnScubYJf+9JmzLXWmjmbzjF0BCu2sV/QULmLAUuCKYMlAoRLu
zg8YLly+0cfPpobW+klhBtmXJWpZvXsL8SCb/Y0F2FGLRILQ9SX1TW2DioMV+PFU
5hbraTorg4fVbKdMeQhO8KUyF88oLOA4VMOUv3LD3kr7ADv9nv/gMNYkpM0iwP+u
cErJ5HEkfYQ9dY14YXSYDbeDO5xKpCuI6rtEi15cnmQNN4Gx+hRXuCfQXV7zsBsz
wNIc/+kdiTIsswK/0c8UgI4GPuNIn84oyG8srLOqC3EKMqHbM4FIBOea9hDWEZ1+
I5EZsG1Dg3FmRwMzYknC6Bz5VwwGiq2a7aPOwcqojtnn6YSElCT4zuxX0DPFq1wn
XOYyq4KsnEJl5PHN6L/akVUis7slpFXoSB0JSIgQhDNuBvgwWtGRmmI/ndhydSzL
4eEUwPXIQ4IkDR9LchNksfodWEEnLm3Guj7IumvPVCDBuHygA8fEPHVDxmC1nmSe
6Zi9m/T1FflkAsnA3yro2qYkQxu77N99qeKOzl9+oeD4EEmzZ67R4k36NOLFHRgu
mjqVOneQ1naPnc8+hl7oT6Ythv8tf6pa+JVMSmZyXb8T01Se5sIeo0oiCGZULmEj
rOTLkFjO89qe0ksb2Lxge0SKNuyPklTEsC2s4FireTYeQ/g3n1In/xZ/COgtdOPA
P2xpBrTRdq5uNiWbAZXXeoW8vGIbGlevWJwk3q2chvVSXgI3bJRUDVdm0h/hhqmz
rtsalf5YjYW10AntS7kTBjF9+PNbywdnyqPkpsakCJteKQ0kVbkV/2qeYL5GUE+T
uA62Pd0NciT9AuIXEmxO5Y6Sxlh+kIBiURSJ7NSTAm32yN32LGZk3btkWD3Vwe8A
JSb5Oed3e7DTqE9SwJI3cQM2GAInDgPP3NXYC86wHNmqzMXb4Z9JFpl2kKAu63Xx
HjDVOtOi+R//uBVGDh5CyDnV2tnw7FtVfs8EDxxxsNogMSYwju1HYVMTndd3aaKb
xSb0g6dN3qM0srCSTycp9C7Na5yyi3FJjR8CTjNHh4+zeCw4jRdANieI2byZB4mB
lxSrUef7k4JJpCitqWnRtP7pr+IK5pHe277svjr8oJEwqjUQQAOH2eoqljqfg/z3
koaPk8F0U2/V9sB6mXw++BnMnHIr9gsOgScqG5QW1zQM/1hIcYy7MlP6ZV/8/tgE
pFvG7rbRmCbYbyJ1HkTHOZ8FMHGp1YdYOgcnFOMudcVwqQMbine8GVe6/1n96emx
e3Lzo2oZvfMrkjvefRyJjrTrgjXfETuqQtpzb02aS3vJzktLxJ2W4hIKtKiJy3Ob
rUhzAtEx2bdlk1d+VCa1xgNnnYuDzGGMrlq4wxY82WZos0o/ZT6Bzw0t51R0yVda
mo4aMHG+OALuq6em4JW0Crqs6kzQX74K3GoZhjsxrhpJEc+6VAM7YOUOD4X/a0bB
MSioQ6wPjQyclaGmOCr0dBt2gHXDIoA2GDtZXWZg5ApdwM1dR0EJnUDOKbQTd3bB
OYFoBbsWy12lbZ4P9EXi5BNISh3gyJE0lquzVR5s9lzKiL3FGVFDRhljzMOZGOis
vMRW5sXUJE5ANgxGCQ4xKB5XNZkfkNgeAOF04UIQN6pd1LnnKOcqXfLhbCnQ6drf
p4hQyH9lGBMiclclWAhMUGfRY2cbqW+WwzL4MYBM+IGzxOLiE/1FD69JrwNfHkR3
TqdqacyiqQhGC6P3i716knodw+godmr7fZ0yQ/UxIbQK7XMYeQabIWzY7tWnn39K
4lbPvZmMCd81Axb5l6lZupPRa8V+lIEt9f910QfSfEafzLEazs0nEWVG5JrospNa
5eRO+m4jPi7SVvuxbh9Z//0lngxOcg7tZeXaS876+3ZpBrOkIb0iHHG3J7D6Vy6y
z7Ikf+e4G1j3k6u482nKH6hLGRv81ZgoftXv3Jrrzwd63AYm//arf7YH/PuV/vrt
23SKiRI9KoiTSURjV6gyG10L2VbcHdtGLF3UmCzPllKobliVoDHNXUkqLQu5754T
4BBylrSxLsZqXLXHzcsNuNA1CvART/nrP1IfnnGtvOVsIoRR/eZXjwHZlSw5za8y
NvzXO0eas9Spy0cNGOtLqNqY1IMFiHU02GCi2ZEha7y2Hwa2szN7vaXNaM+8TNpR
P/C6A45VMqeoUQkFdNdkLmAP42HXN+8ZsGJWrGBqRVMNGzuGe07jFGOaMEzN1d5P
jMTRnQXPkzt4qcE+OiqQ/eW2pKtGRqI+Hd7rMoqNWjSoTU0Fsriep0ct/9aNYLew
DALKqW7qkiZ9bfFejGDX4ExdMbasr1/DYaypuyYE4XuXI67ghfo9sXsMGlwreNGS
DVYOdoRUBTGdJfRV5nczVQeapmIW1l5i6KS/2y/LOCkpvuQH6Wj167W6AsFugIPF
XF7AyaE+1irFwfmCu8aVDrYsE66G2BMstG7wkf+4A0fDXajIHBWd9geuw/cCypAB
mytnRBJfM63cTwP9pOh5pK6DQYu5qm1+7QhjP/VGc8GHIj8j1H6t5KYlzO2p9hwQ
15cWqO+xSJaak3EgRW8TASouRsbEUKtSCKvSYdeUCkEkd5S8Nk25WsExs0lD7xvo
fK2awvyr8kOFqvVtO+pyyFn89B6rjQ5aulhUBtkdQXNAub+kfqPRTeIuuHbd+DgN
WUB2KwI0dR7EABR0lW+ZXtFwuV1yNyXN6ueQlvRUyIGBAFwnrrzlCpVXKPjoNTGs
s84tFglg6bP7FaQQiB8McERIF3Q63/0ndKmFQkmt3f8PcOxQWjZ3uhixXtTg4rWM
PhV2sMZZauUDtKqMGdO64aD6DzC9CeJbxbiWY/yOZwXNiNDGMmtThBvkvvyl5Mv6
S3ZWpx7c5KEXdRDLQW3SbDwi8f3Pmvyhm6nTSbtFIae8M6O0bFFereMGZpmI6EaA
dEh0fkVeQCLGXeYHJ5AZg8sue9GTlf0M6du7iQDIJTR7CdkiRSEOvdUtch/hOBMS
5Lnyy2l/4D7MjrHKgdApuDZY+hypHguD5UWF81drE0BjEnsNTZtrXBdBEx6gIPIS
ihAXCxfV932J8K0kaxC2y5FbanHw75i19M+EHku/nTXO6wPhloFhinsEkizysHdj
1Ieys7p9cMQPUiNm6DB/H0hnTxbnfvmfcfDGr52RuzRo0o7RhZxDHQCWmNxxOdux
oa6pf99qe19X50CzVkjdVb57tkuPJPBpKR9P+kjrpBg6riWPg9NxXUuld4Ke/mDO
1Xrc0Ut7rjMDDR6jvBSLicE5ANiYcbh2OH6HrtfhHc16MmXCfP6Lc8eTP38DkziN
oZjqeqoYZYnWWHsHvXi3pFRgAULEHzCuxukbbIyF8sqex+I91SGS4kbAdh1LDc4o
LCfZebbhMt3zA5/k8bKRSX8k821vru1Qzti0BJuOS5EoBI4n24LodzfGh34u2U/d
Bp16mU1KLrvyahTR84zmTaYZ8MyXtTRok4XzquaPiPp/OHFkdgZ0D2+uz4URPlti
72Kls6i2b6l+Va+6IziEZp0gMYixR8rPV56pJvuSKjZE38W2Ffiakir3Hj1WYbLq
ByjMqjRU804mQVI4MAfXzZus/7Jt27KEvHFJ3YgS7cf94oqE137tDCwAfd3u3wCu
Qu2ypm9P/to2rGPuBa4GgEMRd3HrmtLu4Y+FPnPVRg2rG8nrN3jVRD+17uC0eNqN
+FUNvtjEo2NBrnXZMjREad74VJqHATE7nARim84ub1tKpT7oi8yuzc5+KHl9Be6e
AchvppMi+NDRgatN8QT3UX+8f3EfF/bF1cGJlN/qrHt8qU2UTDTJw1lBe2Qvg2DY
Bf6UCIbpIKDXl3i8hfkVE5B5fwJmt0bwo3K1w0ma3rYK/B19ZGoG6ny8UfrRRtSL
tSQY8BL+nCIOlAkudo7X7a3OgTl04yJmD6rmhIBcY/V0EhRLgaxYmqG8z1niglAx
w+xYHYS9xQ7I+ncuS3y4mlZBmdObZqSMPDB0kq3hqldwNo1OAbFYLwtVGJ8QmfzE
BQTdDRpR6K9ElVJL8GPJmaQaRhvSGOYf+b1abErwI/t24vr1m7N5tp4NDBWYQerJ
kXZppmHvSpWE7mIVr0SRgFOBXUPjQy5Q9RJlkn7+cM9Y22QrXXF5fAQY9+FrAaqO
7HvPidyvFGvR9NnSieMbHA+gPo6r1Mn6c16IubUmBw4pLrjcoSTlWcLhnPfzU/F2
MFsGQ2X6PKQ+iOVdWgHA+UWlrJPrCv5xgVVaHxxYxncKICcEYAaHuMecH75A9u8l
pGm+9ZiXvnnieGnhGh6mrIhk6m+4yANYi1PzIYMFWOGRYEZmn7qAuUlNSbWZ2UC/
CBPpDrstJQOTgZ8mF1wkzQiW+73/BZQE47YrJ0qUoVc+YOhGNdghbCqPJSoRk0dM
BtJwJbutSPL9/0o6vJJiT4zUmDrCnpRtpzjsLnpSutMH5GyAFGHYCgDavrYvd8ub
4uQSplLljkFkn50NyZ/HbMvigIWZH3Lx2sUko4pJ4xpEumJnoYJ53cgjtR/PqXgB
A22jBcxzz4Qe66qXBZOjRYLlHoLFMu1y3wZeIfieOyRJwJGdMT/GjUEr/UnxbtHl
ErLAgjqVQjVm6bRygLJvAp3I5Y11A1LueUdZvGKklVX/AYQB8ToaZLP3rgubUDYh
9JZpyuVIBBoGXrHRhBmqrTqPOvKzJaGTocMZMNQKoEbqy1GsgZzRcqJQDepqK6Wu
ioy3OBHZv1YckR6aGOm3nAYGD7WVxIZ12ItN0kbpsXP6qQIO7/gER4yckOUlorRw
YD0i84vUH+d8YUMAtOGA6Ar5UafcUQG0B9u2FEZyYVHUBDBnKYnRGiNrLgCo9z29
nfiCY+8EKXtfCNZMtxblzHoCd278vyoqXEDQRNI7ULCPhrRePR06tP3LtcKtVrVC
PGmI2aZBMZ1VutDASBWHMdVwMuzE2f/YTM9lgjyrG+BBg8JbK+3L6wztZ9W3RLLX
bIurRUzMoiKpRl7ZtJSs67qbAMTxZGtiInbleH7XTCh9LpV66sY76lFk7tb9xsgs
Z4DuNS2ZCXxSjCndh+KdSRp+wYZGuxjsXb0Bl3QYw5cKAetv9rRAvxcL5h9e/rz6
rmCoeecj1PPXOPzGI4A/r9kLo0Z4QKQ/XXx1UUr3L2rJrfeoaOi2H5WgywwIob/D
ZHGmCEwm/uRiqohB5XJGZdmw8cL/OnpW6wK/JFpvleyAvBezxgI5f4CfywjpEh6j
BZyhoeNPvPWql4zkyo8bNRMvhwkdx+7fhyHiu6yyDsqH/frkJKqUyvYed+MY7zY/
gDpp+uoyVF1wOmFvTd7XgMtBxJOd01tpW48zYnkEjqzExS/ChbJ5Yl5mt1NZsnHd
q5sI2VMvENWFa19o90400i/oT+Hdwd+5J1x4nwkZ2sQINcbMsCXmThUvv8xGeqDK
gau4jvgsYwiFrp2d3Oo5a0sU6mB8Axhm4JUr8z/J7nt9CUZNqBHnlXgnm+stjxNL
tWCcd0oHiOjN4elgd75DHABAVKepSWtEDyTAkPgINLjPLHP6QnGVqB6srHurVy4K
VKRJ85ecTqYGtCugooImjqluxc3LXZ09KDJSRy4cNj/DcJCrf2xf79n6FVK/lf8g
k83Bp1h5VrJi28qIFkPq4TbcnPOL0frZ9Qc9E+RtoTUSob+n0w1VEv5/rlP5gnWE
Z6gmjkNS6GgkopJPZjIAbA2Dl0PhP12wwUajpdDv5aAaCHTJdHzBZN/yGy5dfuK2
YPJ3LqPuNfniITdnNdMmGrWx0CQJ7idA1tr/nJ1rRtgw4h8X0OZCpN//371XkQfJ
/lFDQRU+thfV9GSqQWLdDc90BmYMMGXa7B6s/w4Uhhhnq9RMwHRJi9LZCw1uKrLm
yCuKKTSOBOIyHjydJVIarioers0ZIXDxIbJx2eEmXA2y3aDoQ05VBN8Yay6S1sCV
68gCRssUKYDJQ3oEltSHsDatA3IndTAwdqXmv2/pAtZLyNaarVGWcMLwCL0td6EH
KL2hFu5MssXCRhtU4PuTjuYfRhC8+khIk9FukQIfpUmwDZ9QLmlA0kZ0ynxjWheA
Lk8GU/GJl+s5o+pGPXQEy2mW7Zyvvww5TJNYGJLYqpMwxbI6Kyaq6KP0+FSWTxk7
zftS5EAnqCmQO/B3zJPHIGG3rdbRGGeDRs+J/Nk0WTWToipyvErtgx+MdhGBuWO+
r8Khpvqvnc/oAaJQo2Wa2JRwoqo3zdV4+IUWNQVXCgJdD7u+Ji91imHZeT0JXhdj
avzoVYqRSmy+KPGdqBaq5XB+eljohcp7dJIFa6uXDFAJfelApBwqbBdNCh/MiNnU
iJeWnugDsQg+XPam7YDJxUAfFuJgyx1z8HeyHdjIv82edfUXWErzFwtgm29BW5No
t1g1w/eX0oMSAaGd3kvjAQ8UJDbm3xb4iLd4mJVVK7D/RMC3tzCL29R/npHDVerc
KtT6jt7pKBd0edvakN3d46S2D9MUkbCEyTOL0etq2hXAuVqe5lCrwXflvG6KjMft
sX2P4EVjV+L04KvMfxChp22YedXou+SDzorctv2Zq8ouAEMO3lt0x0WbR1ediDhY
7YPtxAG1AXw+YxhGRwQwQfU7BcLbp+VHuuGFCE8zFBSKqh6Cb2k70vgZ2lSh99Sk
dRwe++YnpDyFDsZbVd12Mv7fTZz/JBlVHjcJLF9rXYPeuaR8e78hHTsmGdMqVbdh
0jNgqyeVpifcCrLTWike1kCFxc+GBdGvAd2lEciIyc6nhiHN6+KRSo1b80qRRlJK
/SGamVaooOuW6fpVfjnlckINajx1W8g9n8KjYioOvHAngh9sfUI2J82TPIMB06Hm
x9nvy/xoaNaLNcQJ09XGKxQM3PhsqrAJwgEl91XCYlg4Gdrnz5ZM87gq0aJ7Tsqw
Rc3IXlcVa8pytYntPOdyWxeHfr/JCfpH9AnzRPG5dffv0vJFt8p4FBL2RTNjg3DS
N5Z5vuOYvzaENiuPqVSBYQUEhGeOMnJ4fo8OsTvlOi/f8EwzQvcoo73Ow/gvjTEb
SYUWWXC1E6IfYvorA0WRRn6rK+MFiyh9gqZInQ73thSpXl6t9C8l4U/EeXLIH3iX
xAcrWFnMhqHDwpZkF/l9UT4e/3VXeDqrh1qyMUMmFqv3g7w1tzvjWlESkuOiy8c2
seva6BCechqAsx3UBNTFk6PrBD7VE8F6nJMUs9FfXbB0qeOOh4Mp7b+Ak13ZzW3R
PAM1d0tE+Dl/FyiyR0yZShVeIG72Tow1E2LcOn20oAjQq8JIyjzXD0mwzsE5hdm5
xwDtg5tIQKP9RZZVxPhtzYMs6RXt2voolygU8fSOry/Q9L4t9WFAsjxnTKKdwqjx
13BltQ1ZlEJKfFM76SooF/B8GeIFjCBYaiOi8G3K5QMV7w4GcPMgY3k8Ubn9fqx7
Bm0m8wkr45R3XtfLZU2LF/4lflDcpIgMP0GjEQXpcNFN48K3c+mQc0CDXnwr1y7S
b0ZTPgCdX12jRZzgUuNNkZyKCFATunKifwKiEKujOgSfIKu81TufURs2mZZL7aI8
BD67/f8Gla89npS97OtiljaAb4YuBct6VkF495rXiYHiGbO0XcGCfVn861idEUa9
mvq2fJeaUbKLL5JwexW+oYKmwGtW3C5sXxq8wT21LKCd1Qu3NkPbZAU2mgDrY1XV
2CnEkT9doI4RJAVmLyT8+gJWvqD1a6A8iWYRnQ7aj3ORmd6A+776PMIje1kpkv0O
ujjhq3ZzN+UhzK1fqrHI852U++HgAFPbLnkNWbY4QKPNUH59RSqeorYFnmTwu2kk
qSz2U1oi7OyzBqfYNMxNZ3pAVsnL8V64ZMxgmOSdhQhW+CzjXIskg9VMSaVm2qME
8+X7uXBnG71jiFqUYhmCOZwE/zl0PIlLAJg9nU7/o4iFCr1Td+zDXYLEFdp70iJW
wvFDo8GQ93E9PpmgOQtIQPlIgriv94IKdG4unKRvMYALtn/U+YJGVoaOHDQ453i2
YvBnrFQo/P03Vh+wisBIvn/W1Oxjo91fKm0vDpDr9h+mH0lLbJQ1P6N8/gqlALon
KbDe12kBR9IiYU8wWhPsF67yymbW+nd52YxYW+kE09oL+DBxYPn0FGlLHflHN6RQ
upacSyC/uQU/k1P/nyrG7QzqY3D7tBJo1hcFtubAkPjZzFo6InjMkSYDtzwZFdOF
R4et9etUMWwAz8pPfALpZ24tJlZkUkC7WG1IzI87PmmLKGpP/RzdPwH15sZQdGgZ
A7ZTQeOat8SP5q+Sw+GdweEbk2uFKDS4XWOS4VOKqgfAH6r28ViGfQgIvZppeB7n
GXlDrmu7zksEfmoiBth4+n+e4CBDkmXQ7GrfRlaY6CH0Tu7P4Vj+yL1OJXrglD9e
2TV6Hmiyz5WHED1eIhEIT4ZV8+yut1w3RTn8FqoWyxi+Ir10cXDyxkL7YGavdasm
g17Jo823SLe/8sFGZ8NGT+O4s2wyxhAHN09JB1R2CXmusl5zatFkTgp6qDLWFq3O
zar5TPaISoymN1qhiMBhtULY99qssU4LcV85f7vjbYDBCHsKNZ+XgFJizKQNXWhp
J8BmKjqGUk4b9p3EDh2KJPm8ilY5IpaZWRzt9D8QvGgniCnZIoh9Mxmpg5T3LToQ
XlV4WW+1/YWG3OoLQeSRYdbBDX/Jy9EIssSEFnNCi0hGFn2DKmlwVq42TJqlfoWX
MqnHkCbRDHA5fuda5eAitQmttyjCGpyR9VeRat7slLhGkJO/9mRAzCxSGwzvMEXS
oOrviLg53KwFtzk4o4ibpzYhI+hAnRZRxWesrOJxYiU4w+ZGoxUYgzzB8Q/fmVhw
I0f2bKBtgH5ZwyP1O+yvalv+dOj+PfuXdcEufGsjkXX5JuETN7eZnXTAUwTNJb8+
CQ14gt7V9Y5U6gxSElngUnjOk8oSQAfVS+WB+vUsR9qyeSBbeh9zpzAdIIJZz2+4
XxP8omcLv6GKsNH18/DrHHRprYdpH3Mn4koFY18s7tK9R+/gVsnWIAV7ublhBC6R
L5HZ29xUGAIBxXGPb1y3Cqs4kOui1KYVc46DPsPmwFlwxnsSjeJ2YRLUNICwpTrh
nm4ntHqE8alWVqZ1snVLAPzXizopX4lxP3HYhQbsIkE1GMImQawO45mt+5je6D/p
QDHkrCvfmGP1cICrhLwdK1EkbCuNi1txWl4LA7zY/4443GrAXgAPWsYPk39uP1Cz
0VfGiD94eBS/FfPOuyDdromp5oXw6AI851O8WHEMcFyRoGnkRycvM+DckQoehwjO
mHAtAAE+0ZZepx62aEZaPonlx8XQg1UtxGzakA7mB+4RPnfCClv0AWsdtPdd8I8E
hli0bZI19rHYw1sjufcGQOVX8FlLCdJH/O7Tbf5YSBoSVUPhKTPs7OUrd/clrT+A
o2hWWn8Bg5VNTptHUpqmPB18JcLbdlxNWEV+kwNaPWiTqZsjOL/xDvPiQF3LDWK1
rrzt8TDxBOpj1C+JKsvgPzo20RB4l51EwtwxUrzRvGvPTeiWiUnr68rEftPzcT7H
f/rOIpRzNj6O72gYzZOH3Xv38DZtNLUvtXEk4K72RzBi+nVXJAly7KJxdSuTq3Op
ImZnohWIPRxMRZXuyiMHRxoTQ01kWpmYeU1auNuoiyi65cK0Y4hs/ii7evsd1U3y
PEuIxq8VKBwfbFuHrfge2+nvC2lZP0AHJOpvL6kxCU3CEQTjQcJZar/DmdYqU2X3
BDmP8xbQkeszSFegDkObdjc5nzZ/CCG3RHu2fCy+8iq/+73vEzwBWMaBoOiI1zsW
X0t70jgvc3UBNK3TlMAZD25u3bIzTArYdrhIcTsQpimiik09J3Y/dLvICcj1XjKk
YFmvzk7z1U4zXZd4D6z76wQ3zV9Amd6aPFps0GHkXMWTAorikpZoYh+BumrL3zhr
zrN6kAclAQO+SzvK85wm8Hi+U7XPdfHvEtPzGG93nnZxipc7+XcRDHzz9F+mXlsG
PiShn1272Yc2Qy1CA9ORV2CASNY6Z/JXgbaGUDMacbu7UyZ8B/yd5LvEpOY4iNIS
TYipwrOZRcG9Ciz0Gd9mAymw7zM73N8iz9/lyxGX3guM1YMgOXgIJ0YwSUA1Hau1
phwNL1TDUvRT3UVKJSdBjfVZJWL4X/owM9MPJ3Y9QCQ9a8c/cbeCBmD0Dyaw2fYU
NU78eIqDWeVYWyY8O1b/Vg5GUNHpM/G02oK3UOCSR8PqwkdANbWNpJz14SgQfMpY
8PRaN9fYqEAxHizsVZBqEHVTevVr7ChsSvgnu57eXXw0RKQqTMh4q7sEVZMtOZD0
TjBOBGVlTRuTTjMNwU2f8wvczyZisUIVvTMFKijr3V3qYYWs+TztQhX57p3+ivMu
DCo9Jw52Fx8x2x/B5BQsp0EFTnEie6RiT8Dp2WAi7ZeOxSslwfBAXVswzITg2I3h
6VyO2XXnUvJ51SlgvGS0dw43kFThhGSFM8uY5Htuugjdyrg/CtMqPTLNfUrCiZnn
/uXuDDwDeDnZob9M7RJ5UBt2gLCWqY46WxgYHYyfSvUq86dM4rhDjdTJutuQO1zl
GBtuuk8oSmwOTUaYrmvzelZs71HK8bM9UemOlk5vpx7jI5Zx6oO2vu8i/w+EuphY
B5f/H11OoZLkX4DD8Nlh2Duu5E5DhJXnKoO1EgPILrY+egDODYNorXvYFb2g90eI
SbTQ1hANXQ88+/XxvEkF1C7mU0yfN3QNqT1PSm6ZoOvepxPLs2zR6aWgFP9qHFXm
QnDc8K4lJD9AJoxFv5T/Kldujoyyhkf+Viu1ntRP8tYkWQAAbIkHZILTPoaNHiMO
7pgb9X9ko8H5dXFupG/8FDQoH+XbSnPsQo3glzzUtAHJ0fm19vp7vlli9kcoyxVT
sb7YrxROYPJUqWRe2umy7aJK7xEP03mMcST17drWHxlwlS3nK93mqu8Q5jhArRgI
lGuF1Sveu+JiDG1C6gxiBzfPwrp8ESaEQqW80b2PDZshV4na83PyYn/7rGGW5JjA
YFRAhYlo9iJ25K6rOFRyouyUVsjOn5+Czq61ty7pzQxUr4RA6CqTEc9srt09l6Kx
S/aabK3Qt7I5a5KPyQ1r8WiAT6kFmRTWtTKoOjJqpGeTE4kSnQYGCbANXG55Woor
Z2bNJ/2WQP3x1CupXHs+bqbbdC/oLLiYYbSRotA2ZsjGhd/0xGDexrGYBCBqqNbO
Rry1Fh5UzYeufBqY2McOBCSOaTbVVSkJ00n7ijFhapX6WpM5tFzViu/UzM7DrSW6
ExDFYVZDaiQ1GTssMnYEcvCIOKBEUFV8E/PIVVpPqx59UVchgpy48jRv6/l/kS+D
oNxN2+N66AOG8mW+qNUgKgMTs5RRGlBtP6HfCMmTpQyIS2Yc5WTrkJDClyFuGT1j
VgK1CnN5R5iZmsuYvjUYBTnm6/2CvrobBkiljCtgDlnqiMkayUqgjHgbUh4DHELG
uncHt3oCxh9GvPJmVz+FbSgN1+e1oHc7hwG1jbYL9BAmUn9BOBD1Kc1jJCds672L
6s3zyo/zWZ+WghXygdlUZCTi7Z1Q63IA57j3mPizaTKirVCmhrW391RR/hygWLsE
w24fzoO2ojrc5U6LOQdzQkQk6eHUMGKzxfTBPEvnbUdX+7HEJtZ9nYvEkz2LtC/I
iT/Ewt9w4+aE3cBBLPKBHN7/jCL6jnIhuFmGyCIdEElVdsWkKjEEybsBUf261LMk
jgQBwwxWx90mOT3ygIsm2UC3J+StCmpqgeOjA+z65XYLsrMVpdbvl/EZ0yTqqRc5
EiD858LRi7xgcQBEJmmlNWrS2SpKhytMYK03kYGBpGgAy8D4qb73IO0w0U3UsaYH
3SiqXjZg/sV0VHR34zcFkK5JJLtBKo7vPYizen0sNjJN/gYucWMgBnU2o8LJlwcP
LPv8m9aUotQFXcOaoLBNZQOjBNTxbuoDKA4FDSp0zAxHAA1Nk3Ff/Z9Mf8CK71kH
QpADgl/ViV/osgYK7cmKQ3J6sRw0EXv7Qmv3rCUm1ep0ZdQ9kCPY0SOIcVT2Ybok
cI5k6o4whOrLyZzLSjTrgq9Ijw3iVlC7PeneA0Ng8V9h8pwc5iBEPzJ72ptP3z8N
MDaWy4p3DMBD0kjmgFYoIyWwWi5yB7Z9SNhIrdxLIjF2HEiQz9+63G/NCTn07o+l
OU54UvDj8kjA83cGWkFqH9WFBVsA+bdsY+JmMyNJDsfRAGvNi0Dq9hC3Gu/AK/Cy
qRqScUiA/UVQW8nQ1dHY/DcPK5hkDEZhiQT3gnE2kV+eDXMSySj1rXpKzYlBAbTp
4UXGZT6CbtkK878T7WJqaXLYSVOWleCmjvjXcbsxPwlX4h4470KoVPjPdACOrxCI
mRDNwozLzOI1JHHL8fvyJrghuvD1DWwUrPZiiSR8/SJLshuHRlawQs3iHpDvV52G
si7ji5FtDHnq9c6fnhAs3AWchLnMKu1x026k4DuR97LlavWuaQx6Z67TG8Ykvnt7
QurXDkzbqBO1eTVXH85ooDSkSTn7dRd3hBYGC7lJiPOYIYKVD25qUKji/hKs+31r
THevBgfy24uL+NRe5LkGtYYykCAgnivGNzG1k92+ix4aInXbexsO/b8D6vZ3ImLf
EQDaC7wEtFJsgNUYyat1dxOJjrelQw45dKzco0ueFce5XeRMTo11GLxKsSb57YYm
N2rfLIGbhXsYdeokjfB2wnkIpOtfFn9XfsRNzM2ZGbQwQtBxMQQ6P9PN/3p4PKoo
N2KjFqa6I0clguubZ1e0Q9kzplD4elbN+BI4lBaR7FJ1dpoUlPGP8RmJZSbg4QYa
tfxQgXWLkYTKya1UOPRufA8Iv/3MOX3pGAJu19cc0kxJFP/qMhGpO5OkPRyncaCE
Jou5DttC5MoMVQZE3hDZ+8L3cRPgx9ejg8/yqvbPLU+HHuugfDhxkvUws2aOLleC
HgnyEzcxbvyAYz5EiqyijkxwQheA9e2RCeSeGuZ6hPwtsHrKxtFF2ImcsUul0bta
d3mNXj1Y7dBCCCE2BZTMDdOl2H05pleCtmXXGmwQDnmyCAZTk3VWnLPIL9Lz9Nk5
ResjkKer60za2NkJvjewkH4kBJ9JBD/9tiV5r2xLtaoZ1FfdNWRN2Gyk9kxpK+Ay
tAsheyJ/RuIjrR13dDxVYgv4QaPdabKWk4JiKYEBlnl3Q2Dy/SMjkPWSI5+fNIs6
lA+UtSiGP0YMx9EoAXq4ntd7uV0R2ohw6KTsuK6AJyMBOGv8zFPLUhAXNkMolMvs
I38dv7zmKUPui0H81aenI4uAnJVvu77Ik4qHYckHUiQ0E9QFsSW3oYLTH1CCIHhb
sivhe5s2t2YhgGnZbcFDlLV11MDuqj5Z3oFyxRZz4k7xCAdAbEzKM188JTSNc8O6
IPM0vWjfvxNCwuZMBjqIPkb/9BJjtrb0c7CN9mwTbKkwah34raok0YHqfR+vRs8G
aXVIWQb2fZcmhenHEv9ADRwi8Qjl3TZAYji/ZoGU8+i+kvkZGK06eYmpkAh8YVPL
xfo/FSTTLc2oyncooNnfefRVH59BwdTx7RM4XoHJVs5+mVqR7OFhEKjIJO3mW2qm
zPOVnLWfk+uB9z7NegHJNUCyTOGN1Brskx+g3YLlaEE2TqnFSPSDlf2OSvUDTJag
i2VfH07qVT16HhKdZytNAgrgWhjZsbzwJBucIa1xYIff+umVPA2rf7YxwHd/DSOy
XdYi2tX/zfQDlKKiri+NCVAA/5uWKOrJ5J1tGpTJCVHqiTJ7hOedUxaEUSFhgw8k
T8zDAnhM/+k23P0i+PAneOJoj1gitRFCoSkZAl4aSV21SHTCyKThWqbl3B6f3t3j
jsAx0xKM8GWJelKNeowzHfwQnZSmRxLr22Nc+SC3URZwrJOtxNgCdnCpBss6STgp
YrAju/QILYFkG2W7kq3YbUIKSeJPM/QjofNXOjUQ9DmpvT/V7dfDSA63DTTGHjlM
qkS9tu6MZ8MqoiWg/0yzvVeF1SM+vAKx8IeW9rWICDYg+h5eHiyD+KGlSOr7gaVK
YnoYEEiKr7bnpLh7YTpZV5jHeA4eNOmO75+DJntjfTctmSTAe7LG0ipX5J6i8DK3
tMalLPyW+fCCUgn6w94eLGycgxANt2kO+wEqHiXTPsZh1BZEgdKcLtxDJyGyNbxA
apcMpFZnJ/cYMIVdGoMTXUjKo4fBXHwS1Gz/J+h0CwcP/dFyzjpxOX/yJPDbJKed
ijANr9lt7A+xR0CrQIot2aDnjHRdPl2sjtZ2L7+/KuM+pzvLuAtsm9UjrFVw6Uv0
XGd3oDEeqAhwB0RT6m9N1PpUC/kmSyYUW1ySptJos8XNSYw75Em+xgazDC1pXHhl
9CqGjX7LNVFNFcD2Juqmk+h9UJwXL3vmpDvRRctDVD+mhDRSKsst6EgLDRqVXN+2
Mviyg0qIMOiFqitNNSuM7BBWbqi5rAnT6MYKQy41XdzdbZhFmgc2wypJMNF7iDNy
DikSiYk/EFLuf5nBr29qhZYPkVyTzcrVmYpyhFk6/dq4VxnR++6f12imC0z4JptC
AZGVuDfV1Glcrh9cT2o99bw6o8qv3P0f8en8KOMuOaJEyvJRaotS7LCqRuprDxjS
pbBFkRTym/hfMbe1BqOk/H201h/bn7gn9qMPhhu6evY7h9qyfYNSqocZjT8Ixhvf
khTQiEJY15k2PcRCcWrMf00DAhVPP/r0o5DxmudZ+C75zwpTqDamRIaJlbW36Wja
jbZz0yVBI8Qmro+zxS1oZPcXmFcXLKp3Q3qWFgzW7KmtL7Wg1Q/JhVJ5EeFjt0WR
sC9hj9Y0Q7pmu/tOdGlxyTKS/UmTLvP3u5Qwg2sBqZSsufFFrGq+vuXIxYJJP511
+X2kmguEoS9OFIIibc00zpt8l7fQcnkcNdps+NHqYu/Jd6Bf3uxKRFjYUGk0Mas+
rM531xAw+VpH+FXsaPnkmbt5ha7533TQPN96mMpNDR2+1BVMxEByZ9TgBgd1mte4
WQHcgaMTxTAgCMVa564XL1IyBP6uusndC5OKOyX2gNfz8FX+obfwx0sD7ahCs4CQ
+fOXceKcNazzXStEHD7iT9jXrLXg8+xiN+FTqo/cLu6D45cUH3ggLHZ92xs+i8E3
DDXCqQhV8JYnIHZepCKUwLFqTxAzKLHIAUveVzYfeHFVdZqAz0wnPPMgwXRqFEFv
aF7kOm1pKDpov/n6JBekdQi0+JLUZYxH4Slppz+eO5/FBM3CdcmMoL6ZL2ZRXFTh
yaoMI15BSSH10H6XKTVdNR5HB6+MDaEEngTfViNDeYRU++X+VYTW9+82M4okCGPl
ganiaz+3lQU+XHqm9BN/hs4vuq5ErOuYhhaGrRJ6BFstpgTb84SPcH82oR2lLxGi
15lz068ypxMDvxYoUjJUtmDsXvyeHZFb9qB8U38146xl7Ru2bl7kA22Hk5ckzSER
hxUN74S1/nXjiEImX5Z9aVP0LesPiET0IbqyF6DioiEYfmi9q/gmOwDqLarF+FFp
hWSuADdO5CLtOFsliTdGbEpw8ZAzV7kvmlP/CvKIhcleB00D9kIG8bzqu7KpcYfR
rmxl5HG8lMhyGZENA/JSutH6xPijH+XHw/yGsTdIyeHCAA1R+kYBFKPLsrOR/YM3
3dVD231ip4J2nCuY1dDTIiC957firK3WyA0ufY57xOPrqACZH8SYd4qUKKfSYacF
su8QHu8Kuwpba4+nESYypUNFHaxyF4q569O5/eAPzzFTLkBhLWaQhvUHcy+X0v+o
a1Br6R7kfWbk4Yzti9TPf7W8Gt35EstRRyofbJ+UAmrmcOHQNosDtTHoiz+TZDKr
x3ZZZ4WtR4jGPzTEckOlwOtjLmyhw6BiouxREr/BWdMcEi1jLfGJ1xTUsjjVahFS
GZmLq6rmU/eyFKmIHCx8tE0xy1mWI/nwugydc3r5d8Zrvw+e1M59PlFM6sFfUEmm
sTlmn4yumElAkot/n0p47OyR2yPX8DeMxgwDy/pwYUIcE2AuTPU/9XcnMvSApuJK
oU9MtXVNj1/88cyxMcqfVyPMOXAv3LLTzDB9SyM8HadQb6xsnfDGNNbIRJ1mXASc
mtp8oQ5uwCTajdPIWV+NLdR8DbV3q+4h+5DsMNF3o7PLsxA0dHc+uB0CNbsalm1F
Q9eAQ/vFRG/hUc3VROMsOvLPZ0INrxTwRbubK0QlXFSikjFRuYaf6Zsjb/GS9rAe
7uDqeDEmmpvvCYaDepeSTu7N/11xxku7mobYO1ZCZI72ifJdcQyKE1Nn3chYXd7E
o2FA7hnXGHikY7ubiXiTj7e+jhr4xY8wxODTni1UFru8gnZgTlKeClJpbQxBpOga
Mlv2u0HpYvoWxszx3E0f9vjo+bTgaxAu+SO1MEprQWF0kZDvEXKT10Jfw6hm4ILi
JGgUvJkSnKO3iNkOwoelNUyhmPmG/nDsDoF++RmjOZxjb2suGUm07XtXh/UI9pAE
0/DSBoEjRMrpiqUAUfEnPdDQNrm0mciWccc+hq+tZKtMp6tWseSTprzI3KkbfjKq
QDqC5gvB2pE3FcV1RJhLVEjWpn+fMNi+p6qrDkiui0UQHaFDPRYGG2QCyVyxczW1
kXzJWEJ+YBfMNJKiGtkyDPxtOAlK5CeJhbNlU/Sg7JU97xU/VLwsNXeFbS5j3EoI
wU+jnv8AKej5ubjEtNgnHYDup8+jEy1qeWZAge9ahyulNKAz2Qlr3KBy31VLniex
uVNhG/MsNa0VHjxUn5th0NHaX+PxPhCyGnsUrxNDkyviiHlzm9p17zCXWczGh7sB
K5Qmh0YvaJ4Y+hglVVPxTNzGm/Ann51TwYadJPW/37e5vrZmYdGj1hUXUtXrDwZ+
Khr5z6OJqNRis2n4CL6JFHrxE2SThoY5zm7kBlC6uejFuTTNie2s5Cyz2Ys5gw84
NVodfLgudYVf1UVo2aQklMsu2it5OookSRRId4F0BwiTbN6anyGNVpy0s7Llyh9m
Mh8EeJxeN0otOHljx3B9dbObaZQPimZgXPGN9dHGZ+Enbu226rsDAyRStLhZM2nB
TOoX8PAoHFXh/5xs76e63y0a+l0WmkN0KwZcvk02wXBusnXdiKDzPeRG7uugRDw0
ZV3Fv9vTm3tSp2S+EYYvTf67vXmJQfR2Qqfaq1biHmiEUvzFmlFF2BBUIxV7z7gc
kqKzy6q1dneu1DPfh2sdpO+G+M8xVHHzyzkteFTfqDQbsdiGiOvMqiXqh8VM6xp0
HcEToetTIqSqMrNhtVasf9cTVSltwgOFsqw04tOT3+9M8tAYKiz947SdQKs7W7wf
jkgF8W0JBzguKawLjoGnUOKXEyfhyzu7wim2yTG3S1m7t1nFKBg8G9PdPIDrhPxW
YdJsP3Z5wtxS4ygUrAjenmD4qkwVd3S6kbofhOL7aVwJ6muOsRRAMzXOfHWk3Nff
UjMozxu5jHYmMox8ejN1vB2rT9MUeX5dYS2BGOAsfOTGjyO98TF4+mGZzPpQMl3c
cK+mHf+k6maO7WPeQqL/mA4h22sp00mgZdMvrZ6S7kKVzV6b1VPBazZXaRb+ToeP
w+kOXkio+djQuonrCdmZX7x6+8u7Fe3ZzwsjhDfwahIsCUmCIgcPRXbdwRPTkmJH
fLW1rXp8bioJhh2PcsmNwlgqoxYlXILPD4r7+KUBX7J4luLevnA6tDz7uUwk0AHd
0hG9E3LsXAfZim558iuNGZuLD6Q9+s5wfyhWiILHXL/oB8nximaqzGv8LxK+QSGX
97R8ZCYHrsAwnxq0fX5Ltryp1WsUWWq6yS83kXKHQ750QePlDqYKWivKGHEf1k85
FcrdvX9U6IvIWE3TtT0GmIzV6kQ05sY2Wfsjyy/mzS52IhSeIRTvXGS4zunlOIDI
uVhLt6JHZ86F0U/j+PTriXSXkCVDIyAlTK9R2Xfc1WEhmKvvKopqWl5XxFxfmRjT
KP2bFg41bJNx19Y/0fHscUbp07itg4ZRZFfuqeZyF0EINHq2tlmQpRJ+D4XJQZQK
hFDKpGZwkqNVPuUNjIcBhKCcq1mX0rHvq72JMNeeEwobp7yEf1q09SogC5sPQHmq
RwbXBHmrQwOa7z1pO51mjGzbPnPcStJ/NswzlnWMX9kWOPkhwMgrD6QOFWwHSPKV
QnZJccCekTexxsiNd5qH06HKajSB3/XcEJZCMDdFpXSs3aObjH2/UOvY715zlSXr
qVXQdQt74TzI+pnwQY6IY1+S89tlC8bWiqgvUkN1YFUWv+vV/JPfC4jj6l0Ii4Z2
dCGdRa3hvnwHFaB40Uj6Mo9L5ou0MuV0c538kSu5usGgCpqFnjHOBTZKdI3R6Mpo
dYqViDhkFMOj8GAlmdo3U55Dyg4GWh2fVt0qXdP3yjidsKYxa3pIERNrF+mmP5XY
QKtK1e2l6kozQb5HHvSCjVqgf53ZCHCuLBX7GZdS4cWe5FQHe+JAKy4Cio08hjJI
B44oBirAnHfZClsyzzdoxz9vwvhM0i8PJhN5MOhMAB3hPAvSijB5lVQ+e4rwKkCe
L18q3BldWfE6FMTbAVHDEtQtxzKC6OhjuJTz8sc5u2b6V17k4kfzzJmpIOIBDWpT
60EV8pLxYiG2QV3FmaDiHOY0vFMR5DPWK7VRspLfHNU4d2Sb+vNvjUMTdkgab8qU
V4VPrPaCg4S3ePMovZp3RV0jKAREt/DklCyrxeSsxgmBwlPl1UUgITVvSUQ9b98A
IXuRygeSE6libAdLCEv5TNGgVS0ZFP8Jhh72Cy+RSFUAjgtgmBpnt4vTttJVhvWg
Mo39Kfx0qmJ3M4LP9rS5zUIzhx3vZk/woPKO9QQGXKuUndmU6OwjpE+6DI614BSe
dctveuOjY1SQrjxnr3hUWroYVq3k4Eo943WBBBvNpyG+LrGbDKr31bVaq6Ui2oh9
6xQDhi3MVDR64eVdPcd79dXRDbpI2mhmDFUmm4J/St/4EzDTN3sVOTkUUolRmVKV
t0rgISpbBZ7MATKKhOJSmvcSMZD8lU0eW5tMi0ifH93MVZCItUjYORNzjRqJFMjf
OjzN/ySzt44kP1rLPTLAtTOHqG0xSM3a9tQ1yf2LIPaKL/e9VyECCWnf9+OS+1tE
KCgpwiSb7WadQJWRAGg9RKqLKwUU8lOyt5iFeKarM/ZZqaI3DTAtezhR3WhTkpSf
njddybR2Pn3BrhJNFWLCd3DUbrwCk3TgnU9dDvejHqg3yDR7hYB9baT8va61ZikO
c8DzyewqU3T+6cfmWZPNCzT0FHFScwYriCwqWPx0iVj4e1IXhun7H4Xb+j1TXp/8
j+BnF5kBLlErnXHq9ohJ9XlLZkdv80H/tfuhz/+ZrLHbbROPKoRFkc/+LSolDCrA
dMFC2f2gphBkECcKH9mpLBrnq9BGWtCTShcDNBjBmyHn/4b4vfAv3D5BXWbJfT72
KgFjbSswtgvsB+h0PJP6nhK4iMIJCVgCNaNByezL7Qoy54n4sK7ZXAIHn27T1fW5
8JjSi2IV206RYbZKahAja+7u67goJCdvGE53u7CwEEraxorh43WiM1TQUS0Z9y6v
X46bwzpkspM2JBdZKODyTKV4ZZVI8YN1byDx2jSpGfYuHqWH71gI5AqAloRjVbrP
ABx8xqbAUdg56VPuJHkflNDh4xuzZmKBtmR5quunHDSV2Sj4JSm+1KlRKPJKMCbK
xwNr7rMXhHHP/M3Y3tt7WglCWwG2c4yTY04KTyW8sXl1VFN5nKdT+xg1vsrWMkeq
GkhGS8bBLGbOYWvGduUBRCjGx6EMaprsbpIZK3T2kvZOfTAdY12wZ5QPjUs8Aay6
/TPX7L9YGC+PJ1X/EqOFEUc01W5R+fvYorcgXYZdu4WNipbnCYvHUV7hLMPW5W3Q
dzMOAOKeN0jSUzGdkiPkEWTqrDtM7TBH1oa5Rt5Nn3WwbrzboU9II48zLyyGpBuz
5nUwdNALGYsaKmpzw8QSHi7iBt8gdnpVjZgAAtzyWHqOAx5KZII4teaiqa8j5p8T
MeR/CODP5vRf2sTOYJ32vc6lrMId+vuRZCrYemLh8oTEcKPRC4dgHd0q1PENpQGp
P5++PMMooUaWTVEm8bcg+waJ2W/J9FauMcOvAvgqtnjUCVxlPIWmhuJXBiXKQO1S
lGS+vmTI7mse6tez48RkWaD3R6MC26tdaJ74hU7RApBQNtvS86lIHufOETRYMfUK
Zu2OUtoiNRZ6tMS2JfJ+8T0OtHyeDC6m2G6vW6x2+6yidZZERVmdu4Bqjay0xCMj
crmv7yAJh32b79JtTS1VzwbOVC7Oi8sutJ0hSMnRoD1+Ec2yssGUlsoH68rNK94e
8hAqVtI47zUr2Jlr5KtYS1FYd5j/co3jU+RO1md/IVdMXIh75e5Vijpxml13+f9a
XMpTXAJYCngqyvc+bF1aq7UAUWi3vlT3Rsobh5okMAWWF/TuBd/kHx94xW2LH2FF
yobD4of3HjTVZxCNLASY1g/Yx11N7QonLY2CeKr9InMwDGjAYP6cQb7KiEgNPACc
nW/60r7i2G3FT0YdC9/wk2qWY1jpcGrpigqgdUsAtjfqbU5szIO/o+kWqlKJU/10
AshJXH0UZoES0oVOEsGqvniuITuOBNkrpP46ATwnaU+1enhcPfG2893QLFIAZN2j
HFAjH0kl0prkAtYRQNjtZ68CikTW2r+lE/lS8k7aYgaLBLToq8zFWn/Ub360W+O9
Gw3KW1Gye5jDSGm0ex0fTZ6Dt+bwB2vdEiQH5t4pmESzp6ux1V0BIzpr6DCcVcu3
gpwLAJ9hN2Erla3awwvATRHcU9QHjNmQ6o4SAJGCpH3nwXvi9uuBCquOtkqzCpdM
v9ySIB+u8kv/q1SX7/J338ojbmoH92PZuN0lRI8lkKe+5cPlxhW6GBJpx4DIQUDz
42qZsK3MF2t0JkckyZU5+Vtr4zLulyaa+YX1jLfFt8F3k8+UGnnmH//ByODuZhPU
A7xHORsvGJI3beSKOIoYScYFYfwb9dpsNExNwWA+kTusy5BeVAoKDcxk4tI+r/Au
R0uuMDkHBPA6TIK5mWYN7kQionSwVHracM3nzZu0KMndCaCxj7CjFu3P9+7McYuo
C1AAWRG2LDusceudqv2T0qyF7OKWZCMm46Kjx8nIcfy+ClvcfEdxu35Et+Jx1oil
FrsYmSzSmhZCFXL6P3/AytEBx7DZ3isBzXTT6NrXVw6M9cBB/ES0O2pLdeFvsW1Y
JL1cQDSb+iGfaBxzGQi8i+CKyKe4Sqjy+46l5eZNVDPiQvPMpNbO7kS20R0isE0q
UEnQ66d3dst8r4ssh9kNgcI9urGdxleSHiNCkgxP6MusA7m26ERilgZAZHd7pN1N
+muDd96oGsOfkp7koX2rOBCup631J+0236tgs8x8uDzR+zlU3F6FuQzYLnKlckNc
dAh1MEklm/pPKVOlV0MFXyt/Ylw/LzCPkDtyXvTy+EHWN4mpU9sHonRtxMo5Lq8Y
hCAGYnOgK43erOAsxkTQcuHpY6YbEcu2V+tGKEU8JJChQjVBjD/rGYnxtHwEYSc5
QxGs1eHdagW01wLURB5DBsFsv7PasOjovxdilkfaLgM2G6d6gWi5S0eR7+tyFfN0
X7SUSVTGbPlTHvOAQc52DdvY24BdyZ1rTNhqi57jOHSH8HiwcyE7ZhgqQjF5ZZEA
XL6IFkXjMYu9PeHpsgLHHbqj8CPdxhX3Y+OixEFD2ag4ks04ks9FedfPT7CtKpIy
54gQg2wsJDVUJqx2+SCI014U40tXIVeyzNEve4QLDDIA72jDkufce15YJD+BbCHX
yNawYWrkqbhBpS9IrVHBOIB8PlpbRBHiurpzB9b+iea0zSIqLXK8emIweCVteDxl
eusORFndDKtgCP8flu5XW/eKOg4ZC3TQ17eQQTjAU6PVktps5rcX+1MQjgIH6Dmd
P/NjDn7m55D26WRT8sWRtM9TuCaO3O/hN7QwxD2TB076n0VTmhKbSapCoRZRBWo+
f3cV/rOWx1uEk5vuVh7121sl26zrFg5xGjDh7uOJpWHoxQ1+RYzPyHFGaIstm0ZG
21mGIqFaGitQY2REWcxQ1WQ5GlAuRZ9Jtu/9ydiHdpL8ooVSW+/2yUVEmG6bER+W
3kTZPcy7nGMSVUY1Lh8lR6G1ml25xCYq2Ykd/PvzQeblXKYxPBNf4hv1R06kXvnG
ZMwYchqJPY3XIEdyvs/k3QDBlsLe+Y9/Brxh01XjJo5L5DmnwcHuQF1S1WHbLf52
24Ku2uHran+usss8tcFx+kRa3+WnB8FjcYqgvA0Yh0M3SmdbODUS7cSQggoBzu/N
bm/BxrFAPoVb7cWGKbWF6vc/HeyIw33I+aIXfmVW9tLPvuQwW+6PM/kXvYY7wTVG
XayplKGsFApwg5KxE3Rl2XL9FFh3O+rd410hGojKRZuPq5N+1vEFU4osrzXf6jvx
RJ8A0zTDhXvnkvPf0QSFXBSEniPZVEjiIY7vRmyEAJOC6TPoU9CBxTlqJYr59v0A
Ypyouenechmj5bY2ZzK76wDfqIc8CC8c5Muns7J7p7+f8UqDtYfhTLz8BPa6ifCA
m97oeOUf+wSnwzQZMdMaZcss9E1LT0iOINXM5b8t0TSXOsTvim2DiRCN3Xbk+9ha
7WFKm6Wsf4SDPUWAtfOZezt6kFEgcLa+NfPQHHJKGW1Y273pUDFLHoXHEv5yQQ24
wi5LcoxFSq49saNRdLpOA+1jsVXy1gD2VQjXMoXbBUwSeqYkPjBBWPDfcys6P4BF
vgC6L+3532M1K1nKEQ5l+eFwHXdTYNdLnIIdUjWqejVc2+f2Ty5FMrwpQYk4Qx4C
QKL1T+g5+keWWR6JuqoL7qExRg7hOfTFd3XyD4jjusXfagcSt/NoznA/deulrinC
KSwIrtsnPWGbHuo2aVXNcGLniVspzBhLkhim4IH19SMvpxAA0BnKPn1tsMZ5SlwP
QZPRAcZLDlDwPXSokQGSTcw7H4zu8bo+XITCSdz8JRZm+0Q3IDJVaegTayILXWai
sdsF6c2qv1GXMzDhvJmm4g3aG7Z98vyBKeHMuukc2RikO4OOHR1R3/0A6MXPQ1B9
R2Zx8lQYrXanVswXe6DH+dCjejeQpC+aEqNba7RszSVymXet5QY4ryTF8Xeialgl
U8JRA0OxscwFd9RGrq79X3a+/MIPa9AQxqJ89pcV9OWV0id56EyNklEzb1y358ZO
cUXjLiLMZrc/muLRLjnDcil6c0whR3IB24a7zwYZgEUrw+nTgyDLJs6R1zNZRIgO
fqEmSgcY2nd7C+TZX4/kOFK2vX/cQMWxY23/pLvkmyTjDDtINjnasA2O1enA4IdB
ulC1yL+ZeXbMD/81UXJJsTOrHeuDWWIQOaJJAD9oCOBM0KK/CcpHWme1ZfRe6A1f
huxQ3yIBnHRpncWtuVBEcPXf9BOdoEoedlN2Rh6Xb8BMA0BO5qK1BeL4Kx8fnLOF
pfAakRQT2w2Qnz9+I+/g3R6K74hBKyGVehreyt4Lw8S2iKJZNiOzVskFYMZb7kJy
hrM50K6M3n7FSrVZkXB8KsZ25VjvivhJWiLMfr0Pnkrro1+l34QsKItXuiX+4CTh
/pifVn1cQbXcvNzPSXLcBbcmu45Z7e5sfQkWn19be3QLaoHDObJZ4J6M/2ds0gth
KZHeXto70OuMbwN0AusVtkWfgh05zVSOX1PjbSssWoSgzy7e1x9PCpHgpl09d9DL
/4HX/lGgO4NPNp2YhyyjSKk1s95tVK/01HcM8PZcA0Ffc8dD93dka07dzAk7kP1J
pNK+y9kkyx9MHRg7QS4LBBlQNI8/xqOk99I8HHSwfkzh2/Z/snZPTpv6GqI2nDvd
Je2hmfclRJKmtKrEjRwy5bTJq4ulJmPGi5RIUsaKB5jy+h/F9/IHub9ZezeSGK/H
dLUYSlT95dJVFkbJJsmLuOkNaeicZuu5YQiweJ3KGibe7bDSKIJN5jHP5EJD0lpf
pbPI1oncqazGZwThpdOvd4NUZDOcw7tndJcQy5cFSOm1hD4Q1sPiIR1Z0WTTQoTt
n1HIFMxIEBm5BINK8GThjPB72QE5yAj/kY+TEk2UaD5LiaMOIQ/IT29ejDFtwuaE
VST9yiX0mM7MryGxppspL+2ObVHNx0ZQdQXVEGKVZN/RTTNNosaiVHDQT8UlfGG9
ewNWf1Wnr9EvTaDIHy4QPNLFIsKUpiS05OdZPHTPwszZj19OsJfmNLEMnJzrhPns
E8pundS7xwOy2ZzvEQd1KpIdNn+RlaFfX4HKkEtkbXuWmAiGT/HfihlaqwED8CVx
J6fuXqaHKK/3URAdvwRRGMHWwkjGH5E8lLRUKigoorQ+Lnteq2dNz/9RcgCcKo4w
URO4kqSw3LhPEpiAzksDWc3prVzNtE1PpL2eLdU1I5HvwXjD60SxpHXxA8OdWJs6
DhmbyMUtoI6HHpvZ+Wo1oGJo4ElB1sgjayykK6EFNwrtR3uF/COb+DATgonzrtJE
wEROuPRH+AUsnpfsHmvTkNNDohC4E0UqLCtie99NjMe7UXJFHlprpJcAqkAcQz/P
gwkSexKycsglYK1uX3SZnYwUh2jKR5lTk9vcKacQeqoP9eLs7k3sm0mxasmcZMg/
XPcPpqmcohfL/Gqtafc+2k12hk9dQotFRFcBV8ENJsrn8Rckiaf9RT2M//oNagbq
EzFVTG1VzY7kPj24m6UovRb0m9wbfOLOLFRyDk27K13vVyUGjSA1W93eHqwcInfj
MdhgLYYK+0RWxQVbPn+CueqDcNUiiDgrNrS2BqeM+RzLe+8crBUtSHNzpUZ/xEhh
J4tL3lDXDsNcv7rg0bgu8c/NkfcBKFQ9Bz4VDHPb0d0fnwmWfT5C4te45VW6vM5a
X82sL2HoNCnr0ML0KV4nNtqA3eM73KkAoS+lExs9ySsntDSdMRC4S1fd8KCYJRFc
0tghWKLJftwFujLPJS+qilN2tjEdnwtSTgHx53cDkyfq6LutN05zaIVjG+Itschh
MhsbI7qbycYG4vVCyS8AfzwjylLDvlg+AUBuTyVRwFoIWgUEQSli334jcfIJQ33H
8qSK/REbpLRiFEvjk2GZs4HC9f6BIN3Xsq7KsmzMt8T5AD4f8q3OPBi/dnAfmECY
VIwMNejOXAvejlbMVUaDJFYU55hxS7aJrEBHuUgXQAWjtaQqsaO0yQveGpqlkC1d
wJSc7u0F/qfG6ea9HA9lHRgDuZ4MCyppsyc0PQ16tgn9l0aoRq4+nm43aiXPTZhQ
z3F/hQoCZRQfVUTQtlEIyeAJCcD4hJkmrIn1BYXS67iQqrZ8IBjCS6rCuLJ/odG6
ORrMjz0PJtZZ9iKJS9xYpeSoFb1m/lLQr8RPp3VbcdQx8erdj7U0C2ygtwsqCEFt
8rVssFhP9zoOYKpJ4dFE41aybOLRCCue/idoNzBZWrvWl834r52ivAr+WF9HLagI
TUFRELPRcWQDERksdPnDGqJyABLZi5tYwnie+PgOWIlli3vvz3GPdgyLJFuh+gEd
w/cF8SDrBBX+5aBMET7U+YKLmkM6sr7Ha5D+tQMsUpILEsp620M4Y1ncf/rgZVNo
ftZxR7FPQ7LRlUxwf+i20DRVC2xvZhugd8XQ6dpdkvC5MdIdK+PO4iWMWH07s07u
6fl+scdvvTlhTS03lqEv3Bp0YXZE221tTvGIsm3AmuEkmE3BsQe/ypYb2CiX9hH7
mCjCtNavJ3ZoDoYHAESgeBUw0dJMie2KYdLGMoL+NiwxxzbiYpo7NdYesWIx7Ltn
WXU5KN1GsaL7cBuSnm1seZ91EIlh/xlFWk+IPOSMoDWvPC1AZqtKaUV7G1YogRjL
rrJheO81q3ZopcRIYEmhKwXmfuabweL5iSfgi9SVvvJTFC+vZr3WjgXaSeJECRZ2
N1tPLQRscvGFums+xiGWfny2o30CgZ3LpI4eQZSBVc9MV+XIOBjjSyGfUGbrnXT4
osXy0y+u6YLv4o7Ypwv3D5+kWRRKo01unYnvKSKagNlw59zKzUM+gZ32sPjPPmoa
yUhdbxp9MKLU3FKR4NOIBGTvvC1fCYm/we6Xy4MoobnXpadzCMcZAN2EDaSX5pmg
nsDK1rIRJuAqk/P1c4MA3Z8okAFqgdhsrohm+OD7UgfXrwr4RF+nL/C8sXnDOtRs
giVeGteXhCj1/uI6WVs9/7Bs7wIEh2YsfKmt3O8L5bwSvqB9N4kKQIfs0jEJxOGb
Z0LlvJ+SqxehdHnMhAv8fl3WfHJSVhZPT4s71omVb/ayj+BKazfhm71x6o34MLLH
ejHIrbAkkSObjcVKEGwejPsfAOSrSI4XXLaLSz0kPw26x9hCK079aYcOKdlcxcVH
Qjd9EdXFpUwC2xdoEdCScCF5p/NI2HFPGko5j29QPZYpyILGh2xHmi+QUCoYfaYT
cfgv3YPFMgpGlclpLl3ByAbCCPb0OqSHYGQyV/WwiB2Lbncj9iW/etoMJGFu9Tlz
9tGAE8zhYZlPRS3gCBlirYoDESPJJUolIAVa7kRdqlJY2zpO9TSiDnguCtGLbDxT
t2sBOi3SZqMmHTuTd54HOP2WMcKPSucuPPpRJzbf3wDR0kz6M3esXUvZNodY9Re0
9Z2SMv+gDr/+b51BWWY8X4AFdbAmFjHpSfmg1S1pTBXhkh+oP9mWkqceA7npJaea
yuzmII6oSL3JJsoGtVaDk2oelmqaehViLSzSAd7h0nhSajeIdRtP1ojo0Iclt4F4
A5JHJVLL13pH8jZGhmj05obecdfiknF6Rb6amfYN3tvogSO47k/0byCwVwA/KWk4
JHiyOHPaRNzULuHoDfgre2BWUP3V4LjmBCOwrFJ5fOU3CXyJqVZ9ggMY04B75qjL
GzspjTKjIS3CoIbg0xzv1J4DOMKNRDJOXtjmLC6vTFxwMosH1itJO2ZhenRVGh1u
fCqkdV2sB/hWPMr+v+T0nm2TVuyhfbhlJ+9KOi21ZVECQrvIi2+/y0Gu9GM/bNJA
foFcfiIfpFjRjV0vU3qolvQeUsFtHk+jNOs9TREh8BZWMv83LPHEuvaaTHyvGOxZ
CISEzSjLDrMdPUreNkrf9X+hU7aikihm2W7MaskIg2NNRcx+fItaisWecYnpHnXv
SbeadFCVdWOL+nGQSYR+nnlkp/Mi0qK70K9L7G7cS4+l16dEixMer/ngNVZv8GER
ToIyWWJbmPKNasaiE/ahaU8XHv4RaraJQ4ll9gt5xSAOzm0b8sBtoQKGObt9QAga
wFc2wJN8YhWT0aKmLeueBYfyrvwQCQqyzcgVE+mKSmlytbwJ7ZeiGmF1fa8LoKwy
G9fhafHudAo67tTvk0iB7knWHa8X3ehpxxBcd7Rhb4K7eZFrcJPaeZQh/ZWUmcN7
e8G+rw1AIdrVVsXXNu/jTS1StrwpleMXZABQzyVsBdNl0WgwHGvQZ8eigGdjWvwz
RokphqfdPoq3uMRhOBy40kKP4Lk748/pn8v7FkNeKRuYyuwWR4mCValCFDALTwJe
0+E5l32ZWYJ0uT6DRf4iSnVIokRrhhJGbyWKeeQwpSmWo6mEI9zQ7xa4NVeeHXed
yCTgBGL1UoFEZkk4PChz8hg1oXWoTNpOTAV7AhcwE9PyThhPyyHq4OBidLjmqQOI
Hz30rlVXcXlhSM/fx2NC1P3MqE2goAxaELdIVa8NgbFU8ZoOD8JPE7NRwiK/T9Rr
+3ptaCA6L9Xced2nI4Xr5K+qY6mWj9q8TaRbqUCjUpuZLOE1G4NaF5y/KLEV6tai
qumTg1sob9NP0pCYc/RmxHSUNP5cwLCAsN/EKvd9MSorBZogy6LJE15MMeted7bb
hGkuhym9FIC7OZO51MHjR/TP651+YRZYVOfpeenZtVAG87LAL28M+6tPvjJomKpZ
U7ZKjicX4s7Ip9+l1PrFBxaX8TkJWYNGxu/r3bRyoq7T6ZdeK73dt1FSJmKEduxw
FUYfeOKsNxCfs/3ZQHLWLd3yZaSkXorrXypMOK9jG75teXgKoYsOrunHfvXqFYvN
aAtCj42fC1WHRhhRbwV4ZUBX9x505VkF9dfh4X3dn3ID83TQUQk10pQiEw9tu3e1
/SzEz7GS4DcUqodQCp/UzHbecKD582Pf7jlMUJ7Em3pXQwIoNpcAAR8B1gLX3kvU
EMexWMfe4u3JWXoJFz0ueyDV9s/YwB+sRzHeyWApsTmq0bpVxxrsF60pYuxK0qHP
I0iQlUkA5ceol9X//ycgrd7PmxSEni7Bszo2Y5BNr4KL3RM6TO4cZixkvhZDaxU7
HKlojLo7vYrSCHLqHdBn9KpguTve2hj+36cQo9AoL+OC11MMwEt11yYOgblo/bnI
xpoP/gwnUrs5ByXjH44XIPqZlc+yyEsI+yBKIGFqzauIsj5VcCmj4Hr+v6CPJ/A5
jQeDQZDMfq4ejkGXmlLgQaDLYLGcR80eKLhZZ8WO7OLAfWdOJICZpgQsDF9EhgFf
zOfPj3/SUoKdLA/K83UOUzQ1TvAI7Wm1rW1mNf0ovHm+o7FxqH1RCdjeGsjC8kqH
UZDsR+JnzzvMa/25idh/LptT4ArtQQS4qxFM1eckkoZv9xA/qc4Y8YecGw1l2jGy
o9RZTBKLgbV2go2/2X8Empa++JYr7TplHI+Tt1hUZbKDIIlr3TJKux2HQ6F2Mk2N
kr/C3M/nJfkMYStvRrT80jEnkyhx6Ut2hBmhVx3fQxG6oK3LzNI7KKfA1qo8UdH5
jMo5+A2R9g2Tp0GWaebKzarmjEfSvRzZXC7QK+BwIRmpePmKo+DhjBJI6GfPbKp2
qFacAG1Zh1H6I2woiRjbSmzpcBIxgc5rVmdK7/EHbkCwlWblMffYVvJXmV99OXdo
K4A9YrIvxn6q/nkF2M+suwtX5pd6t0tDzCBnYTrapHkTZAT2i1ZI8wMNOwrtKS8v
i43yUBoiB9jYmjMFeGL2MytB5/mECe2f1UFeSAiJXqDwol8ioAseFIR9i7p/tzdp
jCZ4CfR3WrjNSlI2K0qFYgxZotC3untzXln1mOZq7KxuqNwwjTO46CsOBb+pAQeE
VDuxZpPRInnTe6xS+Y/STmqm8i7SGPEro343G+02OtlRI/SctKwhN8V6kUabEEqq
/oW8JpPTh1FwUF9jXmJfE3JyMV6ALlw1qjfi2aLcAfaoyFDwS357ir3M8EcYcsF3
kNq6+/DEepWF11NvpX0u92BRnmD5DuleSh7YoP3OzINUlUheYIcjYNeaTjwTgSFT
UVI4h1R9c3R7q/AY2bphRbkjU00fVt/o7yZ/XdWSyue8wzETtmV5qAAaae31nytw
cN+e2hKV2vSbHTqp3Lm8uStVCb1LNtRBWXkMzsWr9CvIXvVFyyEwA/ZLLEbU6WIw
Lbw3m+WwFqeSGJmXsZ/WqjB3ZM4O3pP1G1Ev9MyLq9mjk7sQX1W3alPYU23wW1wq
YbTWCImOHLRMRGQ6NbiaMmDelKxTN2czqVO5ISex5WM5dHIVTtvqqPHy/FC6NrSc
kDSOz7m0z3ypoiKOCroIh86D6P1KAQvvKFoBlwu8ohuPI0sQB9GPelPGgo+tk6ZJ
7QoeKtuLPsd/EX5SVGbkId8aIlUKDHNimMLHpy8oOAkBgFxr4OZ5UwyhNDL+r4y/
zxjO9mzWARf6qgWBC87h9ZxtqfFWoh4jtBWdrviwqUev1wNayZRR97gSIu0nAuSX
Fj0UPiNy6LxcY1SJ0KdKH2KXLOHSyOPl5BXY5ITOcvlE0juQC5vRKBc0YyRdf1uC
FK4wmmuiLVZsKhyZcU2ib9PuaoNNzv80QFT8F1oskzjNtgpzwCvQmMcQeuQRvPhC
iWJV+SG21rTNHxbP7yEN9yRcRMc1ghg3D9sqmdrz8aAnjwPp57iHC91v66MLsl8W
q8FAyXbcErHMv/TujFYZbBlPdQwFRluiTbzc7dDGmBBJlD0BHMZmHdQoNhNMIlSZ
8yM/5txJD9s9cZ0mnLp3mrEZSArPgz3mmZTHKpvTnSXX2v8T9Go+prKiGiObLbUJ
91lctcbOSBhiv/SEnvCmgIaeiZe3x1U5sKUQKE5hR5+dyvJPU0KG5KZhGCYRvlzx
phsQWyoy2YG1+zWFadw1RxFrA/ltLmZ+Oy8ppoL1qiY+sL241cPSnv4nROfeuvQV
Fgn2XH7YIWDeDR8KmJbaDaKldNiTny/GmOKo8dIpCv0jzh6KjbCqf5o+RHJSQRt3
zRE8Kmrpd+khldpiKs9miPCBoulVx6YL7RtX7j6TZ8DwiZxOAwLcEnPfAkRgsqEk
AJRIQjsffWBtcjP1FT008SLazj2MDUam8cBpDOlHlb5yAhNLGxcasiSvc5/AkY4o
LxBA84EnrRrEUKPj1j4odHTWM75LHueMgCC606MxJ2LI2r187OTaC+EEP8A1ruCm
q/4fQFGzA7rGBR3TRAL1qcxJLLibitZRbbPkof1rJzEJJAIVbSx1xc9oEIt6nWA0
daHFw8N7wGo11f9NQQYB9KtWmTs96PwQmZoK/V9BEEArKTgR08avnbehD/jAz4UC
mEKt9nwV1D2IWficSYFIVMapCLZCDYPcRWm7I9S6+9C0ldEJYbdgfjp2rTfZPwA3
wAzjkoItUDfGRHXTqfbCexZyE/roN/p9k91lSY1fhvAPmX8i1RttV10iUgHeRyK2
DZz91ie2rcUqs25OZ/ANY7Vbiv24/6EvGxpM4Sy/99JO4DVRDqgxmxh4/Kjbg0z1
k9iANJRUXjlfI5q6fIg77ajBRiYKH85vnl6bfS2y+XzA4FRRaBuWFBoDn/W+39rC
pL5Hr20WvDIj7ukEvKiCClo3RdH9EJOe3Dtcr9bm+6mr/r6UcKNdAbsGk0Zv37+0
QJIjXpRTNFp8/8YBvQ8sY842/e4cLJCVplhbP+CM1lWpzRRSyirUwjYI8mFkpK9n
E9QNNfvF6xmnUBWR6w4KuiLyGY7kJFuYTIKgbqVrzoHFRUEXXWvzGc0E7dX0U6dG
TqWQR7tHm0cTRo+7jErtLWDukii3H2k45ZAFioJNtIDgXALoWG0ldrDpE0Eu1bh/
x6n6t75dquSsgYTGCB93zPcvztHwcZckSbaUysVHeftjtOC55Lrz/vLTj+VSKKRn
cMTENgRaCmYc0WmTth5IGL/X9ZOUuhYLVTd40vWWl0aABOgU84vadhBj3jLfB4ZM
TPYnIVOZatCb5nCdXsVMLmMfTPCKpd4FPXNQOsPWp0azLZkI800T70t+eJyMn7an
w+F/BAzHeauYOYll4s+kkQeepIgJuZZjBxpTQsXel7aCapKQFdlgV9qwFNQmPTUN
bzDONbYxKfp9Sw0lUR7j38IA1pOFNqX72nKFZ+QVi7Y0EXGCg4pL75en8QbDZGQB
gDWymnEg1EoR3lp2oNImeHqQg73jXQWn5IHDGCjLmyJ7IrT55FEKvzxS3xPY+xrk
Mh2DHDiTsk0TODFiKuo0L5f9BKur04oP4rJ1Fw0GIOYmqNrs2SF+NhaM/Rx6PHWC
XiOEF2rTMYRvk8sQAnzP3qGChjkXr2BFsf4OoiMR0Vit+T0Mx8bcTR9F8+k9IUCH
ejYzYsTjnaIX2g8uBERYuAUZYVeYvRxUQSMXohX1oGJAq1BfouRN4Rb8iZcvs7d5
XsdqGxDD74HXHuA7qF9seVh7ccJY7nCRe5CPDKCKWvEwydtYsLIutrqzTFN2jCVf
JDcQObwDXX1IMB2u6CKLLZAnidyPUx0R63WwA5ETYiH/7NzDQMtWnzjdBQMsX+UW
6WtARrtd9YQLnEIS2RZqJ5Nu8j7HI0k1cuxnOoHJBKKWxvQzg3cqT0LktAeYWdIO
R5x1vxq8SZdTy1UOUnMlxVARZ/mmTd+Y5M20WCRkRYfRf64tPj6+MIA5YCbXR1yD
LsGgiGIDa9li5v7+0Rc7WZsoBM15RY0DNkeCmF8YgxQo1tgmcQetX6spbpeqXiU8
wjGqFWhYLiz6pXzTe+PB8sK1OhrBetfu3LT0QRFhayPhe5SRi5/8zMlLR6MDmJ2N
qH2MAktoQbEtdVraACypy/O5Ya3sL+ighZ2oakpB2i6OvKwBzUYOK2GbvT+pYxNc
lkxkb18zr1TaRQ+pkDQD04blG+s3K+7Hsm5eAQgqSwFe98baAYx+TWctal45LpOU
eHeObeDugW1gClzc4xCLMRC4rJylRLiKU4HR34lNIpM3iwPJ7T0aiockcjvPj1tS
UYj4vwwjsMFEWld6LiQGVVFY0yJsbBtm7fzAZA2A2DB82LMUm7lINnxzZR2D+Ehv
bzBi43fTMwDs63Wq7MKzDB/G11JGDhJfGd/FkS71UUcdQXbsyI2gD9AqFl+Vx2KQ
Dk8BxDR6D23/0yDk+/kMbiurNeS2aRA+mIJDbrpZkdmWCSp2WgnLr4xSmV4gj9td
5zL8ZntANxyFHenJ3TMDa8GjgznIqfeHvIP1A5osC7YNCUirnCUec+dFTcuqi0gN
kUzPS1nnSHBx3V/OeD2bLyFD6xYkT7x4Ew9jCNfhH/DSGDzMXv2qeFpumsLUxapO
MMR4BjsIEotcHYunSNFBJ7OxThQ5VZ+J1Bwiy++iwewAs67kEODybqeWlgH2wFOW
RtWNVWTQ77bzxuBsiPU/Y5uFgSm7jDv1SoW+hG/Eb5ItfXST8eANAp8H54gNzC/T
5+Zzna57OfYKHLibBOCBUChT1Bpk5LOJq8LbR1c2Uh/fVVlUk3yoweIQDDmd8Oqk
0QE7QpgoCWUFMYIiqIP/qOw5RfUVNf5UqfwJItBwJ/t7K/iMsf3P7F30y3hAKc9p
L7vy7tYGPJ+GkDU28vsu86kiEvjY9aw0GFkPHe4jyzhy9iTtr7O3VeaO1IblRHji
3R3D/WsOEQ3mwzKZj3suXQhKNK+0BPJ7U7EKRy9C5pmuLDhJGBH0c1ygWsBWwQmU
Sly/bzszjRlhS2jYx116Bk/HTNgFT4pt370cNes47yTwPiCk30W7Z9BmExb3bq7i
itEiAcrECVbxB9OEz+cZb5oGDajiJsEYlgQl3Lkvxd5xeYRIB858E4lx9UsSnGBm
/f0Uolg5LZ259q7tExrV4TALwreqpPfRdA1pxeumQwmJL1CPqeiRYzq1FZn2rL40
xj3jfMZDznUz8K66nJJc0Ak520TvsaMBm2yn8yaOqjZxjrNbQbsCnBAlmIKKjKhl
QXLTRv6DANeMAGzgVJX1QsgFX1cIhKeSLAAdiXUG5cc9KE2CmxEa8hn5w4BgGgK4
L29mZvXvnw6VHlO99nVjxy1FzrMidNX8RtVJVgIv6ZRjSyy77KIcA953LDPwspdK
N+RsrYd88YcPOUByDWT09ucv1FqatCRC1dSzcHewjT/IA8ZaH+vVYGxxxcbiMXme
gQ40KxULeiGYI6VZWjaRJYE7BlO1yhVERPNN3FIN+6GXOX7dY3vDML4jVitzxOZU
d8k/dZsHxta+li2aPEjpj+v/qWyp8jgPfDA42b+KQwOgWD3xDiBKmDEpZaCKOqsX
N89XuxI+QPzvGrw1Y1GfZmd5+ikm6CNCRxcLBmfXwMNjE155MJ0YP1v+X9pbcb9B
L7epKCbqLWQHXUN5sPtr6/b78PGxwXfkMl3Zy5LbTt+8atmqN5dExfl+EBA+rmlv
gLgVL4+Xu2ri+jmjeqWN21I1yn+25X3pCW5KIov9rVXqnX/ifplXinhL/P49S/30
Fs8hmmDam9qK2seR3jFnUWtYa5VH2zwHAwiBfWVRbwA6wmYENqYahrz1dYhlTCed
C+2QsIXr1P01U0E6NmeJ79qUyXVc9/P5MQZvdqNUIEsvCcUCxB57kotC3Rw1m39u
EWHQ2XZlR8norqiaj8xWmZLpO6YL2nstfrcevGp7yXp66dD60QkQNHAd9ZCb7oSe
zFvzhl/dAx25ep3oeoqenkGyC6Pwe5o5lO8efEIOrNXWFKaCpQ7xm/CBLur96TYl
6i+aBg9HOP44XXvDEzoUo1K1HUW52m49XwY/CTJsBhPOWRqLQKcgIaYhGJKRc+Mm
VGtQVGh0V7ORXSUDtbtS3eGItBCZgECOaZ3hCy5pR6iohKBQQianQ12WWAv9Bbwh
HdSA6IqJbnBeOl9VNEydp4khBhPuH7K9xMtLj85zFGr/8pMFzrz/Avf2qmRS4nQJ
zfrkkOUetwlUM8OwTCWLufdBQR9+YTg/EU39ZiH9TR2Ez2MZYlqYVhSUPhqOo/3y
mqaMjFPPwrs3iKv8BY069/xMmuvMspapD6zlJIYxcEPojb2ZZ+4VfOsKEmJW/Nu5
zl3YQSdGNUj0MdEjITeP1bE8/lKLoUljzW/b/ymDInPo+PHVTwIzqmiTwAgjTS6o
1pMCxJICVbBvTnRJc5EKBi8ath1+wHHPUQC/gQdATXNhjEBr3qiuuvG7c4M5TLoB
UnglWov3VsMs1pNwEv+H+Ne8djFQ65c0Zt5yETeM0v7p2VBzW52tUgQqNI3VPQPd
FMZhKqSxYZGkQex/eT9h/AFxCSa7DmzF2mROc6YC4cIGDuJKeJyIFNTNucgfElyg
Fk6bsCtvBF4a3488wlwAUQ/jpxK+RBMRN5MLn1Vj2gkwaoliKFiq4mxTtBsmvv6L
Ap85PTC67ff1+p7dx6WmCrkKBJtBjGgV1gXS+BJi63JANCjyahH74EzrOJSKB/aj
NYw67DFUmxHGBXpd2EZSXpo2Cnjt2L6go4sAS1Qil5/N0oMa3sDq77M5oa/QIwxD
ytGgJSEZNu2wqx1zN5qt8MTVr5YJKbT59WWSLw7DStOqbzYGUSMpRaKFZtSXi3sO
VQTsIIrKxfFr15ucSE+AxHPUzepMC0XLBJv4CyWqWxguLdAX06SSf7E/yPxYn9Wt
0NmIZtfgLgAnZZJkO+UtlLwFkphfqs91Mqx1uZnV8iXW7aVe+9RGSLs/H4d1u6Yb
nzEtsoFlDdcXFsXugutsWUQ5wgOdAOPVeTAVGxjBDVftgkFjjMvo6wU59IQg/Y3O
oxlo1rvYilowe9BOVquin98rm3EufPpWLdAOBJrd6v5rM0aBNiBG0j+AgGUuVwx+
csZV2wtAWpQTCMCjhr3La7KLzjSWCBlwYKKAVa5R5hF/jzQBPW3a5euM+Uq5SCu0
6JQuezuKcqO19D6mnP0dvCSwaZBoGHNTX1c0UYV+gQzWriSOQqvZew7tUOcCD5nQ
whreC3R/wpMNUArZzjHgT2lTTn9buRruEuqwD8P5xrtdONiZeVucd/7e/jerE1Eh
/QwYZRhbbyLsbpfNGudd/poRdFijfN9XrMQjMKbcK+3AP44mWgTQWVyx4w8g6iWg
Xb0wBrcLJsNmxkJw40rCXxjVsxx7Gu4SN34ZJ4ay/CzIWkVHqDTlUqs7yiCyPVgY
sWqxUPN4zaIt0H5dxgJbTMZMkImFI5LGqp6iCCoC7ZqIJl2vWZBKhfcE0rZsbXuk
X6lRNsIpSi/F78wWEkHTo/lLsR7srtku37uqRmT5GLjI+76bhzfITCTEXDnJapQD
YVXdyXQvsPB10AHQHlPUUgzGNb2PyecAgyCChLpexEPl7r+dmPaGOf7z8Ov4m0Dz
ZE5/2LGbqj0U3rTm2v7HOUDXH8HaQcEV/UAyCTenjYqLQara3JfbfD71kZ0dGOYo
keDa+VP9JBfcYU5eCP4uedHItH7ugPV9R5irkP+XO9RcTHXO0Oi0U87tWxK6WAfN
2XjpfE0TUWa3jZ+5TUCVP8LQEvbqiJnj6tuUCe16VGeqAJcWKvpbmgJAHPFdBkp0
8i+FfMIU5EEcRTP+/hryBQ51IV3D1Ey6zC+j1cpU3oU3jlA4zftJwX19thPJmt7z
5Cs2Dc6iE7DQ+ccBQcoLczIO6BBQAQ/5TL3BnTWYMFmr5/MZQogGQLLLOS4KFgP+
3jbPIPAqXlBpEcaiBb3Fh7K3Jo4ooQDhKI5NIOmwZYeXbFCnq6dtGKL179D42yrU
3+mGiZ5/yaZlixJDhQ7lRMlIc5WtluoVsQ/FNfFktjF7IS3kVeqKo/EwSj1zoBIF
jrzQb3JpukqcXmx2ZtknsOsKqjuVh9pN7SZCF/6IGFbiLu9r0tlKQRZq/FKymo9O
cb8puIwqcLaekTmPs7rclcdB+7e7Il/IAHwMBgNCupYgck5n34yBHhFTW9sodDAb
13HLpwjxGvnNjpnFRmpzhSk1kTWKwo3aHQlHhCMA68tOOooDsglejBsqNGHFbU3r
ZEGnbyrqEc50eba14jBZCBTrx5LASS1Myy9p/VTd2CjmHCwJDvH3f/ck/mA01zT2
oZL8car1NpJruW0Pf369IoWlX9Qz3XVmfN5yKXIjMflv3yfT+fw3xtfIqRCs6YP2
CRn4k+M1Hd6mf496KgxLWCyJ8b2ISVXzyrAMM0Zep25Y/THtwe0zYsVC44V1rWMt
DMN/BTmFUvIeK+cde5t0wuzyQ+DT/9JnFmNAHGJfrvv+dWa0tXcZbSyhN/0K0YHv
tBpeyF8EGja5GpX52Ntz26d+w82vm8o0h6euNqsdyBWGH5mMWjBixgn0VuieEvsH
r1SV5U6FvUJaQNsFDOJgxiNkJ5bfqyiQXZrj2723vb+Lyc3eL5/YtGJp4XXrNhmr
HcSFx8lqlNoadLw6KWGkXPRdEHhUjsrRr6UAQ5u7WCKKsePemomvXpwp+r2oWwgX
zgX7LQ2GLuPzD2TyH9svwjaGc0N80RgfgGx+ZOI8iwRrUqienA8LK2OPODne4O5p
gAijx1krcMnP9SvvVSFflb2xKYsdL4BiIi1mvQzmgvVjPlzP2asS3AYAJrfsb6XC
AwLU7RiZlxPCGZ7bvT5cM/hUTh7R07TpF986TJGozDyF0PV0n96wsWqR9yXl/xz/
cXtZlhXQkHPJwpF5SHg9FuOpZDbX/NiMve8hRILxCySkSZYXVIh7HiC9ByU8SeCS
ciOeJ2cU3ChggH6e+TwcExcvCjnG9lu8UWZIV5DMQd6ur7bZusv25U3121eqo2n2
ZuOoDPWRkiqLW2yDwxBYsuQqhWh5pYkd3v6qdMQcI8eawH1ExfPKxKku/KfKlFFQ
y6HQyvUCFuuSPHq6MNyh+VZJknjqQdQGb4puDQLsOQ9FpytwjuixrmkwJ6ENebFy
/7no3ZgbkSu/3nU0rlNErSc25vJsiymOjvyPvPH854a8G/jRIPF2pXvaYxU1ZAzv
QevS0naGF8X16M4dL4zj8WR3CMDDIE1YzFfJkvhMXbhhK9w1dCfAmwJJM8CRi+Jg
yQghUcqowF7JWDy0EvsChjF6+StONc1PWfMMTgCoYr2eDD46nc4WihUDbzQwtZ8n
EN1O1i0DDPfTVU58ALdlJ5/TY+XcUQmXvnJSV3s1eeaBy/OCOKDogJUIZPzlAOHS
ka4ZatUc4tVKMrqsLPP14BXi5ccstuf6YapOQ0zzDcw7DPfqemV4skkOdPkznhYS
mjr8S5q2kUodUPEHJlMyy/WR7CbdVKHO9cO7pbKvd1ZbXH0Ox/VQFWznh0YnfIT6
CCpp0offqWfJHy0VE7IGbhW8bwOAaUKE7VBnh3Vcrs0+YTt8x5KTWrPeIt+XWS3d
AqV79SwlP9OJi8DOhoXrigTJdsE6oA+hN53eorhLIi+PAkqlacpguRQTyZrGdkLA
jcNB1xoCc1op7FUy6sRh9F0Jtq7Jf4VG38t7hZTNFwNIcTEPbytS5VGUfS68eio4
5plfIRzkqrhoj8msX5WhEjDGN+NkXjkxw+/5lg9sCU74UZeshPjpwczGAIRVEL5C
Di0TqBaelz5GQFrEX9swnsqeh6n4HbpWcszQgFpWUJ69fjB1uRiAN6RQBjrYLy3r
D2rOtjX3pVADCGw/zirHtcUbsm+cmwFvqD63GKTatjythviSQpQ2WYSsWRabllJs
3hz49Yz3+vK9UOrm6TKyMeV3H+udxGayDFl4DQTd4/6G/BmAuu5YipsLM7xlD/nr
eWVoYvtg1GjxN0BFaOfCTmIVttwohlGd34zvll10fcLSo5GeVSMEVA1VdTlD7ntH
VnvcHgbEMDMeT6Vc3NU4qKUBwJGeFaZtQUsNP8XXe51vjCwQwjSApb0igX8KN8PM
yHERtcoSh48dxoxlD0RKOfmdY7j3RsU0yAHXtEA+KEZl0qVMOI/lJ5qibZkWjF9X
tPJyOgYiPsSayCKcWlMKsyumTaJjjyx0YwqLlIguynp5KiBYiXnyODw9MLaRAgf9
8mGnS2ETdO1hE55zRVExJqRfZliVk7KK3BuiNryt4ZrrZs7Qxdn8GHWxDoZn6b2k
VAYA2IbyKPLuIHNmJBW3JHUFIlk+Aavsdgvz6MsRiD6UlQBkphSmpmYi9vVzfqyo
59oKve5Hb6nb3bua+zQgtBnpy800Ee3zKPtgrbywGudLffdxfu/xpkZTTIjxWwz2
mktbfe/w04PeMGiVp78LpySzLOMQk55t+xccHDyrw9NYe4snOnlr9W3Qxv/HGla2
40vuJBvdkgCY1bnYMq9+4ukZOsVed829GHthgmSQI0jGy/1KcjvTYEpMvKMy0oYa
12yONvLARCe9V/2E8B5GhRUk+PMwJV7ZPKLTuKT9dMtah1QP7mRYBxEws1BpNHUK
SkSRyMFAIcTY+/PEt78zHl4IXFdAxsK+S23CILY7k2nu3n+47el2twRYEKQltKzR
lC6s4jAlmsOi17LVmlKUCiaHbRhQz6HTpomUNH8T4S9NqLch+8zMSBD6ug1Uq+kN
M544TW2vazJGTm6vIP5hjc+GjvThDanN+Y39Z/h1ayenynkAm2EdIUED+DSHsvaJ
K5lm1eXsOk5p7U2MAUuwnNGykjwo2ezLMxzQQosA7T6hzkpBJo9iHyICHXg1DmQL
Hz6bK7WUedP/UKcPJjiBW49L+v6PCJ5YihLyyfykm4iigmA+U821ttAur0yqFU/L
BKs3h+9efZFpla+cpWBnZR7B93fmKeR83ZNEO0KX+sI8LNf6L2xwzycGQmQGtyGB
iRWReukHILWEc9lSMiGNOUzMGgrkAY74Xumhis78AvXsDtMJdszJ3OAkTRVFzyrT
qm3zl3FvO4pEefNHKDsXlEw4NmyEXrunYOASmtthW3q3/FXZre37RfK8C/pdiZbY
izLKiyr6NzZ8RCDtdqylxKJigJET9VIQ5UALuTbYA+zpjPFpUAZSDkkeHHESeYiq
S5Hf1ABaegTdcnB3kpvU/ijHd7n4/qDFUhHtw9ZczBPEbHXBqAvzzqGWZ6RvEqy0
9yQkutKHMJewV1Vq+Zcw9Gtp36HWnRJh9DXJ90OWmPmz8IDe/3iMjuQaCKJUBa5y
6OH4pRbG65wS4tpXZlkmrx9XCnNNuR4iuviZ6QPyKSItGF2fq2uUGwvdunvzwYeC
VqHUqleFmwq5PtLqBi0zbGPmUlMJEgJSFH8srFbM+TdnDSN+GmC4SV1M+eOPS7uz
9kBmcPcFYAh10idXDqPyY/rI/nGRaqFnagZoU2nj2oP9KdqpJMep3ucBnmWQJrm6
ocWyvaVAn9G+aEYxh4nE+8gI/z2zx1Af1yAxb4fqSaa+lxVpyG0ycGuxZEbLITZr
6ZY5gNzkXEGj2ym0m9sZdej9id4+KCgw7oYtaYXNoktG0qp5hH56wy/4SAscWtGF
rAM9O/+71oID0/zFvjJOplxgFBqvpDUdNbj30Ug5KdGBJ13SqqCXx2vgsH/YjFnY
w54p1v6CLP9xdXbWKc8G5cqiYI1/A9iFEjNoogDSmU6I4qgSG+AWTUypo6Wt14UH
Il/FSukaMoOwWGVDyBJc1wmPoUT10sBu6ZJmL2OvTzBBYo8o3EbY29zWcDXBXC/V
02QpobF5d+Y8bpyy6BCD3GuqUdOSe2Z7hUvmwCSmjvEnjNa5qilSyJgjs9fB7Ien
wMCmqALLXNFouFvDtnUoAG2l+XusW6c+M7/T508s1sOLvGeesu3al+OGdGIeBakU
eynqz7MxxWSyNOTnqUwWof26JGHiXSxYh3E8uh+x807WXm6i/AWQHFCYUbJhAH8q
9lBcHRLnQutIllCRSp3Bi+/PukkMIoRmrLaSazVuzxX2K/SLt9FtKurpX7Dfpueq
9ZwRzSMHt3CBPZ763x55tzB0/IZQOmz+WuH7Bzmx1J3k358+tkz/e0jFPJPWmXBM
xM1RPkM7jbpVTxwyGY6skOgu8HOWp5WUEp18q1QJd40cUFL4rxwYdXOowI4tBbCe
22RcZel4Ed1tZwkVYn19wgqWUOgRWk/aYdpKzf6lscC+xXojar11kz86xHQIhqWY
W+cABRQOkQGHN+Tgtfxutdzx5p42OMIxjRTpcdZnBfrAtc+WJcmYb3BJ1LPiEbNy
+gDqsCE408oYcTWDbI5y4JJEp7GahPXmWOx14BWNN3Lv4l91dNJM75kcptCz6TWo
wI1KWnxvaaKMxPDmvngNy3dizvJUb9lbysigXB3jlBXXfZKyoVhrNC9cvMzYNXiU
zW8N5Y/X94w646oCrOIM3kjyyW/UP9booxrvnpxMvTTe5xmsYDIC9OZ55peuguNu
KK2Pk/mbfMcigtXpLrrwsJxKsSCRF7uEXAQB/9kPcN3aElKtEloc0mJsxHd79bfa
uNcl8E6X6YPh5RLruw99SCYmeMZJH5OHLZlx3L+UX0/nOeQIZ/gUOjbIw4ZqnQxW
IzXgJa0n1HSsASMPnsASEMsbKTKu8D9tvot+MN3UHFX8ePfgkGl56gKouzoBpgjs
Hd2Hhf2Sl0dPrF3a0kp7iNqw8lT2fZftmfZ1oC5vcDfeA1QbIf2U0DaYv2RS2CGG
8pjxNHyFcRiMCw1uDdOHTdzCGmb88kK7osh5bHLtul9gbVZyi5+52oPoxTgZQR11
R1tA6SaSLbPDJzkNfFIAPWCXpIRyAujs42S8P0KUxhWR3nYGM3O2XhUv6D9c69nh
ZhReLWert0E3IFBTlLexuQLXdphCvcx4+7pGqpbWtYm0tuBEMYQzwq/3tadC3xFa
j5t8jG19Y5X7EY6zp7Qwx35QSibxTDJ86xQaSK7brxwYzzZS90D1Ahx++Qy56i0d
u337WmPeA62IGmW1IGNzSDZG40oaqX5qafrEUcrmYn9xnn97x5lmyXTlcuaAXEos
gxNLLlfDWa2Tf3/9J0vLrUKYgRVV7GORKwutk9gkbn2pb7DNaaQ8hiLUIqnE9QBK
DAmVJd+mistgJYCYIuEl8oSA+L5OZIU9o9zu7U6xWL/VssI5k6x1BfVI/63uGtL0
GAsCewcAZ8esRtAAr2b2alhC3jNtlifOLdSM7kZANi2VGOMNokdsRNCwCPI+0Nuw
JGDcDb6LFTMw2ZMK5lE4RK0NiSMVwwAHFHrAQCj+moEXDDdgAfPBR5n1S1JQht7C
D+73fNIUVqx/SsF7N7sFBGFdEzjAG4StEnX6Ox1sz9M2pjQpFFUbxg0Su0eZ3g+U
wn07bJdb7bFOIvaklDTN0y52ZY/lqfJtZ8Ui4vPnfCCrpKEoUjZzJi9712r8pWnb
eFgKkFtDJlPpOR2n/K+UC62k+z6BvpBIv2BC8gZczNJre6mqy+72fWdlr4hnwSWD
qzyNEx/yT+kBMv9YiD0kWdyU/RzJepRagLgZh+b3+W0ZGdN72WXrSRbZrwKCdkJ3
mI+n8vtdN5H2yfbmvnciDZBzVDfpFjar6v9JGwnqduBHa1gEFXJvUWryz2t6gBgG
WXsoJEfUEM2eif9405B6vmbg7FHTceOfZUbxdH3L+DLJu8mtzOqMgS02Ug2G8GMu
g8JzH6ggHabr4rY3hKTa22D0GZJvcBfrTN7YT4pJnwVaD/nXxWfFNsfbFG+gD/hj
OmFhuts0STAlFA/lIjR0Rn2vh8qt1fIbQKuVPu4xfAvfzT2/8Lp6rJa03eW1G65k
ATBLas6VYfaEVO9SYQoRNTZ9ZO+Z0elyE/TzcpaJnqbw4W/uMNdNZEw/8davOiCj
Av/nsfZOkPyvWy7OI2jErmABkq64biY2Ntuxg8VjmZ9MlPbjyUj3Tb9bRGYI1rF/
zlwibBG+MU7+2btan99FxArdUvhyVBU9/eZpHhvEOIxu7YWKCzsEVpRU56TeT/ul
g943ZkKf+L/R4Z9QoYa0izOJt+ozmDMIDRUD2T/Q9wS/of/UO/ppxvj1zNpwDX7H
WSr/VZO8XapnJn7fs0NWZaVdePkW7cEbtQ/krbzkNlqs5fdv8ukcM54TLaybtZDy
au//XlwDLFa/5NGBCwVoQH3c4Wmr0GdZ95i2CACanA460Ex7dxh8D21moXTD4i5N
/4nuAC/0F8QlrB/kGs5Awnn1LT7qD4uHp1HiNtsw3WleUeiL2JHbvqK+29Ipxs8b
Lyexymvf2fnc6QY8aWtTmkdOpT+fPTDyOG7hpb0ukjG1474GZZu+t50AEwKmDZXL
EF4tKrIk4q8ek55Ip//4TTnveW1subdS8pDjsv0iObCBYWtiFvFxX0KzV9zpfc7L
lODelFkhR8xXHYJEGEpQOcNiK7NuIgCtd6Vi82PCR/U2mF8FFdv3AJaAEkUwnQgQ
l0qfXrzPdyveiJtaAX89kQcaAMffr44NQ4pPX8o9A66mkCl90WK3nq1nTOKGWDsC
KSd6WmccV8pdeWarJ2jLNzvV3oZsx5zIpmvOg0UWhoBaq7Q7Xr8FLYaXNSDCaL42
NTesAPLGAUlszukt8VbtQRY9DDx4SiFK21+hoqCbvZVgbAF7+gj55W1MxvYVb550
424W+Yqk5JZaN1RE4vRpAkKvx29ZEQcBtxzY/j6MWmbWAWqqMPLbB11lj/Fv2cRr
uw/lOAt5KXyGk176zzfyWDQ+GVBIrKw0Sa74tVLw22vHxNDoFCABjKQR978Z2AxR
HV/lNhWfwmXJRXoFvOx6uTob2jNO3AxRGjIVxDgw6WwjJdUBLgrovzs1MI1qMUXZ
4VAkMFHPV1tlmd/gB1NxmK+iu+n5/SKN7zuhHRcavvlkSAjyT4sPrO1Y/4PVeOkd
7BK3O15KpmTvm0BvDndkUTWH9rTU5qivDYOvlJb8Ia7oDt+fA2OuU6heruIebaPc
JTYtyERhNFfHf3cLwY9pCxusUdyS0Lvp9VZhX+WymP84Ah75457h2wBP9SbX2fEG
XiXRCuzxmNbz/C3XSSja7I2/DoaEB7SjK7v6QCbH5SzBZ7zIvQNkeLDZREflLAWI
Hflcp3sY0tdViJ+oGLFs4YW46wWRFdSI1k6Z4PVE2He4GWLD/zE5P1Y+29U6L+FH
4gg62oWwMexaVtme7mUCNf3yO4TV8xfJhdFWcE/IjrkHsTix1DTIJqf4DqBj6hMz
63opdipSbqYLfo01eLj5U4gPlj7FOV5WfUOojzn56I5ROOTPAsZaWPb2a/GoDaYa
+hEjCGbcYK3nUMjzb5OXDozWKLHhZA+PF4bADzRLUdpDrL5Ejc62IE8S7DibJBaz
kFJ4oKMywFxl7yMJpn6Rph+v0x0Ge/EuDn6wWihO3eLAWajg5kLian7Rsna3bDte
Gw3zTuMM1IJVl1A36z2XunObYeAymmRfFYh7K3H61hyMZoYN6MA8cV+uL+TeTQCZ
UQXc6lV2Xn/RFno9p9yNkRx0Yn8Sge33NCUX8uxly7K/D9lKqkP7HPBr3QCGxwbW
DnEGECNTR1N0PEfnRJhWD74l94FLjPBL8ADMib78S7NTIFD7WpP0f83ywP3tJb9W
+d+QNlEsZjsPgnz2uBWNjg6SBzr/wKE25q8trzNpZitl4GGZZ2u3XfYqGT42gKGU
jEiqKC30KmZ0RwRhrUUt65AMniIo6NTus6gRii9mCQ379hE0cLcHL6Ve18Vd0MlP
WumeuCcmUb1brmlFj4aZ21Ed6bzOVugk5bQR/Wy1lepRMW3N55y3/ATLkT7oPdoJ
amw0EAAaqqYCsFwDVNcqJsQ2lOlLjDWkJ+K+rwjwKYJ1e2jugXZ5w7LuCQ/eVm5N
kRvms+wwALQJxt0yOTrgTiU9tAnZmzp1Ej+Hit2bIDSEZQrGB0fKU6vstb9m10lg
pMlZ41NlIpsVHn/P6yPw2MDiU1Zth+C4iDxGCJt6StTbUK9UcOGMzr3F66d5dtTH
1FEV+OQN6AmNRfgX/KwzwSgg8B2fp4WjIbMaPUlHR5jtMnjWhC9hlbEEHpWPhdks
lrK+Xekz7DXwx6mC4Dk4OCF+D1vEbxroF+I4x4QbFFbBYngpXLgxcKp9+4rZMzQc
6EpXLubFxqz5XGMdmoMZXE9YGmW//k7hGhW5EJtOLiIoFdGh1gj+KvTYWSzZcR9q
B3tJSMtu33dusPKpHA0tum9K26ka/ynshRsrofVIsUEQcLfDJIR6L2CH5i3YetRp
pSFkF6WaTG7IXPH+W4AKn2fe2Jlw+1LMXm9E9agLn7NNkGUK+azW5qpyfSH0+gDv
eh7d+DIPUpgjUxh5861Owyvgo9sesu9HvGayG41cRJ2D5iBTx3S8yc8dGGBCGewq
BeiB6xe1dAAEr4R+jKSL8OEvu7r4LqA3Tg+egKgW5urnEyfnaznrhIKiHfRvauxD
vMPwjuYTb842y4u+ru6xkro980HOjoHjNOiN4KdrkiTVu/uB6AFL7DcE2kxLe0Og
MLLjUifI2zJcwgeYWAuGzzCiedOqJKQXMW4TuWYH5z3QpmygyVzu7LbPm1PPjOf0
D0L5YVg4PpdLNNRlwX2uGGdJAI5kAo5KDaJ0NzYj5nYfSa65sXajCYwFPDcl9KjU
qixh3padl2SmGIwg5Px99THEiqehjJTZjiF4R+4ZjBonud71SQfsVdWHsvjpMJIP
v5S3/XTTjs9VOICjtn05zca5uxjWu/PXODChBkBCks57u7joY77jQbwTNWra2baM
ky5AUVM9hyO0bU6WRLFmUAOSLCo7haj4+3QupHMogEeDEWDRnW9Mh/Qcgdc9fpsK
ixp5VceI/blZKTSSIdnn/MiX6waUPI4MTjt3paztHc2HlCKboisD5GBWzKR1YSFZ
SHkWnCkSGJlnGugVeDeUP0UsAGHsLHQKncShEYglKbl5Ogl+LsHJ7wmLz5q6Dw9N
IdanNnEqrHZjaJhItA4IVyHiOoCFd1wfurBa5jaPrQmZUedwtIe9I3oZYTMNpqTN
xrDhy7mV0olBt/EC70kVORPP1BYCNw8YFJVaeQeQ+WzlvOjL5K4m9O/UpVIPerJ6
t/dtDomgZnbhdvLYDeuWwqP2ksQc46UKLEQttBdBIR5c0WRgOu7cYBEKpXhs8Gn4
wB6STjrKMIzTLgUi24oFVGeZTxJuvg6shUZ/qTJG06nN2HCuOp38kSYUdgefqc2W
QF0/DWv5jxrOwHsTDN+FX0iip9NJlgT+hdKzPeObFLtrXSFJUKz/XXlyA7uLaPhm
mKwUOfLtX5HEt0gfE2ZIPL3B/uYZzTAyXa85epLK73bt66wn7sCA1R7LNbuOYJT/
RdO/utUakG5sW1G0HrLWLh3sCZmJRDAFB6vNG27JLrwZ7BNT8Qkhb/3S2BX7OIR1
HF5NLcShAQTJf/wRKPDE/ODvn8yVH3bFmTIPqmIMAfignokTi8ElGDTZPEDFx9Jq
a4t0RscVLVXtnpfz2HtT0T7Ust1xW5ly0IASqPjGPWMXmYA0D9f1i5x+elFdZpjT
sTIlnp1yDP9PV2xJaVxuVCFpOHB6rnCc1lsQlyYfqW+9ziOGuhM9lB5T5BTLigkI
bg2zBps0fMd9wxWfUEONKrDogKoh56eG6J4LhYtH84wPiKQ9OdS0lr0v2gbSC7jp
on1iN69zDpbjUqLpvpjvZwwjZs0H7yMoGZvitMcysRPsh86Was71/WmmItRCs3w1
W9qSI507OxY21kDNRgKl7FDaCZ30aEcF2ZEv9mJvP2Ow7AWgwKH06Vwuqi34wP07
Dwws7+1e1E5r85H63H6O+oRSMgGoDmj4O/nkaOdO+uJs0I0IVmKpEzq7nOZuW36r
5y1tU+X81Ih7CZgbO+HNkzNq4aW2pvs2pig0mwfJz5KoVcIQEvoeXacwjNPT8V9A
iNP5SBOEEVLRSfpet+VKyMnHlEYMx4NUbjl+rkmqDlQnUeb1YpmtZNVLZVG/eAKp
uo+eOcT3RGW4cmq2R5yC7CQWB5I6oP45G1QyglgKUDRn5YBUy0T79bLUlkqQuh0o
gGhyxX6xO6F58rjt68fn86fxgfknNsWzGgYAp355PfCGhts/+v3/uqQm3uFAobPf
wLqwpe9X6WMxtPOrBv1e1jO0cxOG9lNW1WoIx6IuqtjE+AbwRweoJ/VpBqOXfvpm
RUiMyJyJAUHU3zV1jn5H/uNRgwO77jRHZBXxCn0e9pqZxhg1Vl5i0KchEtxxw8Vk
KVhnuVNjXXncSxdGvlQP+pDKQ8d32WEZPEpVskQlPkglt2lMQ7BA0Yvj5uBAZ1A/
VEjRkNNFwLfHlwaDFcl58nT7ybZv/ODg6C9SInC96Mb74LdInK9NsS3hPYbDLTAQ
0ZGn13Xk6ksAKrOmNl0wxsZpk5fnkQ+a9LuvTBhZT8+xBOH8fSk2dXXic5M2vaUE
WIr5xXV/RBpGcc8I6YF1qwQ/wCWN2IMVsb2lPeN67qNAlLClIOJ8f5HAD/GXtmFq
do0pagGGNvekPPfKx5iG/y6QsgSYNaYYZXJjecO5977iDce7dpxyF1wd6k7iPA6Z
nDGaZDTB1z8JIXDMevHejXI47XTzDqgBoVxTc4cea7pqy8Qx6ILXh73ROB5elAaP
1l6JS86+Guf1ouZMIX9Xky82vN4Q9G2FKGDfRoE8s6Sst60kXu84K9P5LO7yfPqY
v9tLGcJS/K0rCNh1yq7t1IpHgh3/e+MM64Zc7/lbkiF+pAnnx82h75kv9vWYVg3+
TjwiyJj1usqWcwZi1aUdjvZWABeGChybJ7A1Xun/G2XijKtc8heabcSfGBMMVTTS
jChOyPWZJhYodaM1DJD9tgOFXYKSO1OK17toBL7wpC9ddI+Jl/f8VyQaFhzPspir
kSnhRmLN7nPrd2R3+izNg8e3PNDrkmvupHCCdSNqdCpgC3EjT+j+OkguArJuqD59
qGRyx6Pm3sscWJGSQBI1UOnmps+KtW6GM8d7CNHmNP26xZ/kPMIqEHKVqPD+1ARq
0sn6EFzZ1oO/1e/iklIrPmkCHxjtTD60BKSzIVYcIWsLxtXLAlrjhm9i9auriA7M
rzH6eZO4/SoaJKwBa/6b+kCTLxRvZxcJnAGLQFtp5V9jCUbeq3j3uoBWMVhfmrLd
6BOKbj/nM1jhHG1lTKDm/qfaC3MOd8+e6s+OJxjSRvcDjWDAxNxHZhiOjrE643UW
Rhizag0vYWwqSDkMxvmt6SDxfAgmGHXyct0nUH1SSazFP5jTPb0AortuXiZOzL1i
2wHtGK9VBzhJI5DO9fJbrGeEmaKwq8CyJrUQaYBU1ARhjVEtMapq/WdkV1VcLHJK
LB7enQJNepccZ0y/ulI6oNwn5sucyAOKnu4rlRIQHTJmML2aDBwM2QEb41QIb1Cy
AqwQzDQagaRpa+46N5RAqod0T/poOAnczUys3uKPtOaK3Eew3XJzXA0QevgQBLMD
+FcKRwClrzIWCRxZkPyCSSmR2iq3KP1zBaV7rL5P7Ty8EGLRWAsB7wcxG55GY8u1
/SEv3aPb5gezVA/sUErgyAl1Hx3GFkg/gbSk7qSBRXyaqqriGibPsUXev4UenChw
XIAk0SLi6+/ZezN5Ei0dgYGTwI+AwReKlm/lBFKsS9htUVxu3zmH7Gg7lsTaW3Nx
9R2FwNg3HUZZlKPQVNn10oXUN6EjjOzAFckWXKzXpK6UKVT//dX+nPGYttbLOLcL
/cWoutEQt0dz7JpMJCbkACdiT8RCboFdTE2sUCehrVKN6ZD45dB2I4Jn85g3Sw0F
6Zh8app4SO5U7MzTvVBu08sUmo2iqKFAv/vDQLfhhn/1DyDdCr9iOsZ4Yam5Baju
KG+YeuWNCkx8vvEbLtqK6Ow5ehrCyCpQkyVDziZPfP8Zc7neJwONVKEHT3g8+zcY
WphazYPmrdjZQ9e/8/XTpUKRdXfq/vVUWyP8tVy23O5wK30AdWlpkRi4eq/HNrWS
nS3iKR7jUliVL9uBuUD/53dzeNqMzi1SYxpwS3IftnU6dgBT0td5Y0peG3KTilYY
OzHW49hMcZHxzzp+oE2l2zw17VbaRNp3gXNWHkXh9ZJiI4Fwnn0y8HFUY69RqH4h
FCnqHzLuWIsw000+pGieAidKMP3vGwZKhIBIsoraClMTKXzuq/imb3GFBHeQqV9I
fZsxlo1Pm0E4RBbEZx7Nlhvs6uUerVBXZbM322PY8hTDRDs+olGkUe/dEbHXVw62
4vdEMMXl4dE5Kbzg3CncE2CK+YrOoRcEeIpJP6i/XQHidCHOO3lSKYtk7/NITiy/
peyhHaLf8IkaLfdE75li8G9SFpF/vZRGFXXCluJq4enxH+lJKouZJBa4gqbfivkP
8bJ4AvrbGesnM+JHIw/f95uvaHtSD1oM8I3wdzXN34BcxcCnP0Mm2k1QcgH5XRgs
C6iplp+YHgAAJcXoio2TjClN47kdMX2dGdx58OtGmcz6bUNwaCnSPX4hRruKy6FG
eFPNLVu8SsGCERp1PPmT9VdQ10VNQjVW7Dw0TSvhB8mw6aRCrCfSTk5V3Abg7XZs
24OZJpB38qL16PA/OJe9eh7k7l7qLVLJUyx6xP/KXdWagjrWm1gDAFhGFuo/f9st
fRvohu775VCoYwgR0YJz4KpEtIgUu2MC3HcCcHR1jY7i5CMhuqykDb/YVJ9vFeV0
Oj4F30QRbbaNfHJRxxI8Kmw6qkX6xPKe3VDFSoiKyjqeG0PLFqvw40QCyQ0nKX/Y
CxMaEc/L3BkZGwU9mfkqly8QLcK4EmDBc5ospA1d2iUT7vDpaECaDsQNyYuuqvdt
ZbGxJe+MIwLxZPxjOoB2V+WRetPMNct7QbQjWRQYM5dwwRy6dGS3R60tbMmaZx9e
nRezXjjn4Xxjagl8/3yJFmylFNB5w5DRkBzpOajy5yRX63fVWWNSA5noW/QtiLJ7
nKegInXelyDCuRtApuhj+VsjNogLIw0pPyWIpsOFPLHSgsWvFbigxTIrgHEkjoHU
6UDgZc5U6xJd4jbKQvWd+HiLs5gc9hn1cJ6naNtvTCFsccbXPP52HD1pFrG6Y/W1
INC+n22q/xiPc9zwKzvCh2vVZsGzq6odWHAvwZFeMXeVyt1cLLAXyxikg/jFe7of
OEszgWAuFZr7dWDvUswsLTCJedBvQzRVO1HG/p+vevRVxW9PwC+8St53pi8QUIwn
+/6TCoSEP/Pvi/c0G+P3wn7/YS7LHjFoqDFiuetsEavJMfse0QPU5RKR8MltIOa2
PQOFMGaPllA+8CM4JvMERXeVQJsd9G1TYx5BllMhwJO6gtRLf2lZ8rdNRKrnEKjU
XU/Uk1LlBf9OV4gUMf+WHmXpITXuF8i87liH6RoKikK+aH4iMj/+PSnmfcJDnmB7
WeEM2/fKqf4fftznYd9pQJqS9SDJajgTnrjF/KPR+2sNPU4gxAQuZlGAodh1CgMU
q+bBQx0JF2Rl2NgoFn0yeGopQEKc7fF8+HYa189lL2CRL18fh43W6DuzUp4uf3x3
8xi9EKTW9LkgpSRJ6o1QZpdZHLIXnHEiRyGE0RlUqxPYBMraUerFq6MQbhXcksoy
a83+yXX0cLXyPyo7W73cVWQNNy/vlT7oK67NShlIQfnL9PNd5rpT0TakbQGj6mms
RqsjIn45JpgN5sno4/nuY8QVS9lixfahvtjTUUlaJbaIlwmmRoOdJKaq4+u0sQjb
zJJFaW3+uzDyPiUHlKmmWiV2M07oiwVxmHjFTcpz0BTMUuRcH+bZxx94KWe4fu9D
fR3ymhJzlVLt9iufCC11Jt1bASzCrs/tEOLpY7CSgsNyd7/2L7JAApzuA09z5D19
fg1juzXkfw25VW8+TNI4cfALI08tzO/LPQ3FbdFiDTHY2fSKCxHqJgHBxRAzxOoG
MacytswAtQIta/ec62GOZ9O0eugt71tkLonAE0wkP8Bcn4Qd9U9YFKAbiWYtjFhR
hk5T/p3Vnh0RahysShYQLMnj3gqAsh9Octu5kdM9ctMsK8wLCPWqn8PP96ET9CLT
vOd0D830wb9dStdLNTh+yJZ/0Pe4SjTqe+WrD1hwTzQ+o/AszO0yS/ElA5AwXj7y
2HYlChnTepJCEsfnvZM8AerEPjEgVOvmZoMbyHm6mZVf5PjggkHxEtLpZsKzM1qF
SFqL9RNc1kp16E4L1CHry56RhA0PRUEPqqV6Yffy7X/Bs9Pvo82KN0h+3XRhnPaW
m432a8rhWVCDgVP1i0/AuCgDI+HGAto1DgtvUkeFyrgUErIf3+1S6Yd0c+sep5Jt
P8BXbhrpWWI/WEG+gQRAKWiWRZIOE7yyF3LlkV31CwDsY/o2zQuMueAPYG7utQhv
glEHzWcEfu0UXrsINyFT2Url2vGVsM9QcYkxkAi9pNT+8qUWo1QMV/4MFOEpokU5
Gz8zGYlJLbqBbcfNoy7Md2ZqvuZuyROGMCN5AI+Xrbwsw8ZkjoDG1UHzODj6nsmQ
ivf0Ot/btG3WxZDTM1UGRAQmLIk64mtMUdz5/8KNsRvSQOSIBsp2YTQs7/RfxjBO
y7v9dnIWsYCDudXSjU5GE8a66M0Z2SswNE4yvPAVowSTJXQ5w9oU4bYnD7HADJKc
40bBOCnAEQjm0v4YAWDps7cTuysakoOoiHhreSuuRiUJFgpD5j/qJH07lfXVBwEM
Z4O2Ab2r2Wbto8UYdCmwPos50a7/exdI9DWH15P0jsOZJTyDbUfAoKijH++oefGu
ctUv77jqT1NQfK3SuDAL2qw2DfX7Bu7bDu3JVr0cEAUGnPWTk2cVaEuNqPERpwLq
uhBWXUGIp5P6DgQLX7wFIrAW5Kps7HdcYWnrChvd7/KXl2jHfWmDjuUgWw0RtSn4
JjIfjH9KlrHRm26ie4ZueRZa2dtC6KoSGpBHrZiBZ3jaGaKOF2KxW5/UQxr9WdPW
YQiIRkbyvEm6tNENUFOsZ8B8I27KEL0DLX2wINdyXb7v//9k5LFkUcV6Ay5pWtS3
pvF+34pgGE88sEBgNK+rJ0+1rDWoqOzdCKvOG+LuOwlBneub1pDNX8CROAv8+UoH
MHX/iySYwUyuTpJlWTJg/BycLa7qchBf1nEPqt/OiKA3iGj3c2T9St+/15YyvTtt
pqIUm+QPRsGluPys3v8r6PFB9fhFKscF4ajlhJWIgbGyNYZUWqbyJ10GYp51yxWD
/T8UzPdJZzm9K95RRpF9QF+Cax+oiykz8Q8Zmu7A1OIX5ZEFPZrsBYp06eOGwqqV
UiEYsrGUwAjPB4q7caYpZqGl3FJiM5liQ+7jKw8t/Y8O3h/gmJJyakNkQh6l/umA
Dk2cIJAv9D67USluWiJ0G5H2DxDrijkL6rgLPk+ud+T3wB++NOR+J9kF/pzRAlLI
AGniICfgEOVsU2FaODybNejeWRddolY5jSNIJ5FOL+42pivKBXPyQOBCo9Boxl+n
gn69RtX3/3Psv+zz342KPFcXgmytbBXxmLAtQyjsp/stk6MgpAv6/qez4Jo644x7
uBOtN01YzAOskP2eKBCqZy/wEUy2glH8LR1L0RJJf1Iarwmwe3uZHOzoendqFxUW
TNAYdl/siklOP1fIkGTlMsZ3Ee+xRpEkQvYrUii3LXLOTQ9Tj+3iPARn6uwZC9VZ
WcxqGPe7Eba4vRhZz590cDK4cmkT8GKJRlQuocayYBxdn0QUNwM5WmVUotBn6qBL
BbS0iT34wPlvtSqeLHC/2wmmMgmq/GzzlGX+BIYxDAw8DWVLxoU0o8GR212OxLXL
78HnLSiK36omwf5+0F1BVUQPqGYMFBZuZsF4GI3OmeBEqvhrK5myJJxAyVZ3lCH9
VzSnkUyTz4QWG9sL08c8vVpm8cZNi1rlnfxWj/cpw33kMNSMxaLSeipZZukjDZWM
UQrYdhDRyiYAcyO6mxhY0vzD2o5gpweeT727kFmnIZptb6cUVPQ6Khh+IUQUX7HK
OwhQwZWB4klbszBqVYuI9OOnvgmQPpZ+GU22+xMpxIXQP5hJfgc0pMY3Ktfgych3
MRU0hoBduN1wYZg/6EQvQ+Eihm0z0RsreFsItNVH3dH1XKObuF2Y5ekoAJbpXMfo
fL53Bzl1b214CXKBDBE/Yp64/2q8TgMSMePJ6U7OEdozNPsZ1lPuMShEV2hOPfXq
EMyEk9atUIuW5JZAyAcs0dDfJxQ3/iaXj1+FiGG72DDXoW8kI9pRGJUJHRpsTHIv
jhlola7Oafu+mRTyzU6fruFVK9q9jweTCH6EYBVs8+15z33IZLyw556OLh/halaB
5dIOQFf+Vo7m6aANMphRy5F+7kz+3jCBRI5ffhQXr7KMdG0cx2CAivSetZLP96P3
C7vXEL1Q+Q2/3nLtYKUv9cVbAlfu7ZOvi8AQ+oJsPGYVx9qyZNuNChFnjCQUsJu5
RnwY5mGxoqHuv+lZP8uTlQ9m5114xAlOr6r19DoXtClX1GpcHjdomJ6DC8EnSpKC
/P/ZJl0vYAhUw8EIjJ7Wc+qinS7AsP7KcAGNrF48ZtfRW5jwQAWfxd/zaKoXZOEI
3nA7+oGMmDKG2eelGuoWSV1Yy/kG67i7j8YN7HEk5bEt/O4CSs7kNVlzcl1dsU+0
OmZhIj2e7pWGP4XL10tVvEOFTZTJlqpCUXD8yNsJKgAQGY8aFkJiZFCgxhS6mXBi
3kQiHBwbN1ZWmDyCflYXY6rIP8hU+zAIsFK+W7l/4NuQpoJxo5DqmP+GfDUF+zhJ
QAcOtolJhrN8ADLf8+extDZZ+OQZy0Mjsb3ccFx0ISp15O0QzUDf49M0tpav/GTu
mFGzfzRmgMafSi0RuaxaQwhNVqkYB7pwsZdq1owzzVb0VqMuAQkm5zftqWMl79F0
ZXI1WNAiaWVR9Aa/bv2x0HF+VJuumvTFmP8Pr2RVAyBwi9FHynL0+XVVMEV7WFad
7M9EFGFk97fUCKRFz4CUEh2ntHKCs3sDCdQaIJqCi6h0t+FCh4sT0SvFKrktUzIX
xW+3VmJHfEamMSMUi1EeqARkSGly0PKYnE5itLEvWBXSQxxB6/phIP5xCY1/9cP0
nC6pH3XqUrrUs+30NChGZDZRm/W4sP/A3uNuJ2oH8vbjXzQVQn3/5benOXvzFvMR
2YUlF2UWvca84eCoa7Vad7Mg2KC/hoFgLCsS11ZgnONPzsyoiZb6Jl8wqUB6N1/l
DS0clo0IVFJwjU1spmOpkH98qJ6YzQiSda/jvpiZ1VVC0TObkTihN/TTvsUw5j0W
oovIOo9n/i9bseiwJHiqJ5z91iNn/t2hLHDsO3ywBvL5An++nstxHb6oPnwUH4Yp
lhiXZBRfi8u4wYkwTgs6LCNuc2IaKQb9/HcYW29s0A9eI9tH/gXNN4WlU91h9eye
j7hgpplA9NiWceIcqqMRkU5DxenMEQYb1MzKRAsz3LxzNZBGV1v8acUeCBJb2AV0
oKUmSk5EkYAQ3zfXDyLb053KmWOH++90Z3Q5HHL+6Qnk5UXgM4bhASOs3rlJnx9t
qYwfLeZXY/zBI5cvurUig6lpEZSVd55sGYywKeoWFAQSeDkeCO/U3OC9fvouy0t7
OqGriyzuPWH6FC6nWJtRLED+XXhwkqgOfc4trYfMCSYxxKtBVNHQirSNmbwSHxg6
QeRtDdxikhw5/IqsjXsn2vj0sDgFAUSihNI0yEigHYWQbGQkZgNZgg53OIegzJAa
peGUAhiD2F+9+TsetXYsmNqYG98OaR+Un3FUWcIHMmWBNwRhuDvPN7ntwEYY1mI2
Ccko7S+KT4kpbrKc6TAkKO5E4c8O/2nBA9SbN1zn0nwI0YCtuwnLtMA1Ba2uwK11
9eMFBSB4ma2evaspSn+KUcAargxG0ctjUGB82SynHAuYg7/SvRhKvzrxG7JqfKfM
Kk8XrNptyNzStPuepEQBP7szDje4l70TInnX6p9XDRTZ0xxK4oVinMsPwPZqL/0R
dCKP5iygelbv4bVJ4YFwVOi7Z+pM1w5BlGVCJRHaUe4BJkqHtxQmESNomq5MHcSU
Y0clWEkAxWNNaQCjils4eREi2GgLK+dxRkhkcdLIfbKejdlWimTPU/2e5u8wM79x
zClahNeIe6pN365qUXhe6n6hnTaJweEPQe1qYXFf7s3j6+IuB2VFud4pslJT68d5
T3mwV/NC8fZJDWrfcaRqNIcdCP6ZFj0SA0jYfIC+YUWy7yzKEPA4N22BsYKqceRS
JXcWkxkHlvFK1R4ALmUHPbRoUBP26FIj+ynRvdZKETvGBAhSZRGLJbJedhL9jJsu
0VVpPUR6hi8ptZL6CZLyoLQAztftVTpj98VB2k2ujLbbzrXvpqH6lkl/cKcgsdDN
c1j5b+cqy7j2sXR7yhGgeaVzwYG9bzGENKIh+Vev/DL0TIH5CVsqc1x2Vv4d2LRb
TxeHwJyQg9sARp9TAwcftOfBPF4Zhg7BxzFIEhA0BHIzSpGkcEUUdWmjdC4ifQHy
EYuolksqLE0CYnm52az++uUJkjjW1rSKOVNzDRaqTyK7lXX83hQUS9TUWEtFcoD1
vp2Yl2NSmqoooj7xbHPzcOyvZN9RP4ntWV/ROEY4AHJ1uNptQrmrINvEWSUtBAX9
kMHRmU4MfflshW5i/QkmOGFgr5wYJKUIkj4acmdgBnANtM/cEPbX4EPP0jYkphIg
cJ8TIlGNjO0gwF9mjDVLrQivl7pgYc3RLEsNVK8B0DvqrbuGqBWr+0CAEyXB66fZ
eweX41nVwMhsIVsQhRwfuQ3qoceGnKZ4w0PDUhxU6z+vRYLyALGSNAI38BdGm/PN
LRD/P/LuJdEtNjO/RLBRQ9tB09tyXZIZyn8Z/LVL6Km2PTX/whyJAOcIoaKzJOxG
6m8ssHnHn5sTP4AHIHdYn/yYksWvNta879Ja6cMc7sBNNUBrbhgk2BCYzxO21NWw
349tW3Tt424vv/UvAr6Qy5hqyeBdjyhe08hdIbo1a7+/jGn0ZRsgat1KkU/5QecP
wNo3QkhtwcYDu/M+F5E7i/GoT9btYKS5njOq69ErRs/lNV3pZB9+4XSiLgrb2FS7
mkuEdImc90g0zeKV/yEkGoqLDC0nZiSSBBEzCc+3Umwngigv4aA4dUwv2rPDMM0k
3sZe4YHvbH+emDtUZpPUO0Q/bB0eGnQG/tCPHZhSkmqlmDGO1Qi669y88GK62lWS
BxKNq1jMkg+m/pNnPBgHYAdebGH0YBcBwV9nY4+GUFp8WnbDO2QLRR8lodlCai2R
pSKk00wip3XbVz81WLe1RuA9hodTIKXAttiGadCD0dqNi6cXdRu+nuDlAXnKQWjN
ElVlWUV7iTjJNz+c4mdFicptoL+coq8rH0+bN2SCKtSqvJfagE0sbOi+I/KTj25k
tJ0nSKGTXP37KIURruhlQjpZAtbW1PIbW4ZBoh+XAU9Sec/YJjtsxrhNDrSeGKQL
G/TGAfzdoBOHKdHUa8y4hmetWIY1o8AcOZMuB6keZCyK09PEBBXcKLH9mNoUFYXy
JCIVCSloSyki0anp0EczeXulVBC6KXBbTWra1PePZNzzTJJlTsOZjxnU1lwHlMFQ
QhDkw9vrb/9cZp4plblxuB8sQBCBJGjMb8CjkCcisoKkLDYAv5j98VYxCJrFzkEI
wr4GQd5us4zuIfOtTstRfjDZEpoXhXrLtM5gO36ZhexOjHmgQpxK1A+A3WefeTsa
l+wqG+J5PB2vzQAquv+4fHln+f6km2ihPdJOQPlW3U2nURWsgSN2TBHsbFgJpjR7
ib8AHgKlO+opxm6SZKx7LreuTy1PBL9P6QmLOFwEdVJiSrMUHtScxFBw+4CEFo28
JcsEz9ekwmYMesuYGuWm4E/c1C+mKYVuQlJaXcbJ/HxfCM+Al9Aj9FZLYHaHGgr+
0knE7VtnIcjDxbS1gpByhdsS1SNpgOfMJ7YOmdzMHQkLT057646fvwJ/qr8Ns9Ix
p26WkT2b1tFWjfHSyD32Tjg3XuzeA/xr2b7aAD1ulKihi84UkD5c8Oy3LxkJeqdK
mMljij9/D7KAdN8d9qIbiZeV3LWZ8DxR2ixZd6F2Z/9jD373wyfRbJDBy+fGtEfa
SCvc6ovljoud38NMsZqzvq+jm7C2hgeQc1qjd3LiGhE6r66Hrhl3tx7QnHVe3z1j
iS35CZG38P/XLxnr+cdrg3gNf9/I4O04ZoWMf8jFoiNtWJaUakDRxKt74j+uNpdD
F63rh4agukGcEZwmuWBYcowswSSPFJatnx+ONfQd5uVv2hbl2mHZZlNux+6bkX/6
CYNfZu/sE4V523cytGHt2gWEbBnVl21oeGMFO3EQ0gD/LPKMcCGNUigh2GLx6Q32
zI3QuyCd66LmZTMKVvxBf3BVDdQIqVMaPMKzR+6sOrEsgCCzmJeRnIluBM+oerP5
gM8AOUuKOxvB+Gicbm38X1QoeQXLjOxuZdN/JYTU1ESutzmTM2ZpnyU+sw+gjicG
DD5P3nOEqFgn0TD38mABgjpTmXI2l6f791vWySwSJkXWsc9r31AgkqGMkQ8H76bz
po9ZQfV0Tzd5pKLhnmZ2VJXEc2kkBojbEOdm8af77fYiLjvcRJwGdb7qwYHhHV3u
0RLb3Eis0FsoMtF3VPrNwggeHevNQz4MkS6p24lxU63IZc4aCmZzgI+9sl2WcuMP
ID6UaJ97DjShyMsiJti+SaDHpjzaCrT2pPYGKRgl2377DiNbUP61Uau8uSQr27M4
qBXqRCEc+4YAF1baXLaQA7ScJgmFSofoMiRnOmd73+8u4jtYsWxvARrM7RHZVaf1
KG78TXtovAuQJveqOi2ElCwOBo5zIkVQF7sVfhcqHZXzx4SmiyctSBJDM84IFsNo
9y0wkmDxHF8VbjHxqYNOvVS5me6dbw2/pZwUeric88y2NgFwwUfFjZGafUutfU0S
D6us4WjokBUlii5MRK5ZC3oZJyqICv7rDK46N5FZ5atUcrL+KTVpzO+nE1iS1HcR
izrpWyJKVhIXvxO+HY8cxTezUXGVjPoBl4yxDc3z7obXCDmGuciKqwGoOoE4P4au
2wia0w8+5Z3Dt0dquN07xa1N53ZFIdc10UDEB/x+jAYLnpPzbBl5wOLd2Whc9++l
vPsvzlr+Qv+fBij6gXmGCpjt+qeTx2KAOW+0AyWgrhDkspaQVfDHKbVQZVYjn7ja
vVI9CpnfE5mRk+2AUN4lG6O6NBApkAI1t58p+2kIepMoG26GiuUjDwpyoxtxk9k7
lKuxRr0cqUyi7IsJwoeQTbFuVJCiH0K+Nln3k2Yw8mtgsKwW73KzYi65d8Eqrohg
ky/ziNDpMi4rA5seMKFX9Zc0R9Pt0pNwUqfaXaB9U3AKW25DMR4ljrFFz/zDfOHA
OAFXyBt36JWku4g5qcnQZEBfJE6a2oNcYkcbsIczpmATK0U+j+j1JFFtE3eX3qUf
9DVNvCCCJ/W75TFTBVyWb1VpZoUdQ+BKZY3JC+rhpi5MbQpCmlGLpmxFOBrF0vx1
XA2LVY191TQGbDUHPS5i9QVUZ+k9nj8zLUMcdg6Yk89gz2trU62as2teSvJF4sdp
Jo9ITUyfSGj0gWN6RjfenGGPCJU8xLPC4fDB3VXWYoYHVZuq/TYtzzHCJ6ZEf1pk
FKWyJVcAWG4durap39pnun2PJhW9MyvE2OdgRTSt2zu6acx+NH/INJvPV023lIVf
zdzSwX8Oth1TbA6DQYlJPhCUvu6TBt8HFbUqEk3IzpJUIb8TM39rTHsQtLnba3bC
dwy/UHrzmyahW/r6kKBwoKhQHFxHDGZWXqPIP7UTnhH37vSqzOYEH/qGXZgxCq9E
sSPgSpbcqtUkyY5r5sdD0ODG3OkQiVUR1oJ24+nCIIPp/3vWm8UMEnEG51G3OcXL
2zacs4tY4Jmr4IPLnMYqn6PAsSE2hqSJSnWraBtQI4G2gqbskAtoRLHYv3JIjn26
ouXgVmb/pLgdPMo4a+esUU/TH7Ucj/phd+PcapRetWsd0mF5ckXEG9HFhg0K7+sN
jWCKrSgv/31JF2Q4G7iZISEGDe/9kY/aw2pl5kKADiTpKs3EE0GNvOMPwgxORodd
pHloFQ4b/EzCk6eBR4PVzlWvaBSbguy638u5WKGvpC0fa2trKPZANgYhsxZtueOp
+9GAp5SsQICJrMrj23p62eWsQ06nwlNHYm5Pw1nhtWXxrB2se6eE6joyACN9/5mK
O9bg12lcSvRigm/o8gMbOLmu3zepnY9/2RoOieQV1lOZwoQ6674wOGU0qnNqPs0b
HM3YivpHEZkc5hz4AK9bahymipaCl7DfQIYs3EMzuHxpGbAz0uphJvAEm4nlUbT5
Tr6D88G2QwSUCBZFQGjV9HAnL+v519t3W25HBxv0W6YsJJSI11q01eDBNH6S3zXo
whIoi9rNyClv3hMPY6j7VN7NalsajgPD2l4Na6ATBC+UcoBSSscf4CJ7v1T32pTB
f7uLfht4XXotk/Afj5W169arBuDMA95tSHQW6gS360mThN8JXxeS4OQNjx2txQVi
3Mr5P0Rli3lSLn2i3Vmhl5/7Gxm5HuoqC3a3rr/z9JcS0ywiGDlNf5FbRaFdfV7m
Kh3jxnb/EgcJXIJplrAVylXkWnWquewYmCF7z8mmHRVbr5/D2gor+22AThrk3L4X
y2BzVPHjw8YNiUGTQ+CO0dFeuTgbIs2bKv57Ey/n4hM+4VdaEQjL526F+/kgUSWH
DdBzwq7js4S4m52bNQVO7pjtRsDFXuALR1XhoOll2MzOXqbReyQ8Ke3AQ2rZqIAn
MBuHpDAi/jn1OCUFTx//jmXX5Rg5UCvoLk1CMPIOIfW3dyigt9FscnE4kkvOXmve
obRa1rxjd6+ZCx4YOqo818XOuXFbm3VwI4JMpD6Yge1Z9K4E+CLjz+wcUWOPSg52
yJQeAknRQ9dYXLFrwvy//JOZ31DgPU2YD20IKGpmYhVUvAXQ2E793+EUYS+ClDeN
Rr8FO/8blXMIleDLZwcerzrGoOuRNBvZ7utD/T8YhFx0xEapsS80r9lHj/tCSYWI
dZsQJGB/Btum6Geermscs9wlaXEquw45dbU/na2I3p9sfnk5CTmkCxxYYmpPvI7F
k0j85rDvmNYu6NHkLGiJjMcLhiUCOecmhq7aXQbmCcqTSF2UO6IdF6QdayvGoAwf
+qNHI0jmi+hH8WS8soydPHIpjOhWccgxGVQV0ZMKFDrgWim14P8QNH3PXtQIQ9JD
JiQO/Sx070WUsk27ufxpmarLS8zxhpvB/dkNNc8GaC9Cqb30AFSKcsKMbXhmDLjp
7zp3Gvb6UpF5VnTozgDvbjlZUf/IHHJLfW5OIHRKX4e/BPAck8iFm14XSCJHs0Bw
+25N8reHet0kIA5NkD4vrSUtnwVm2DenLZIwawxGsFU/0CQWUoWgfVsIf0dtWbTw
uJHzHM0u3I4f3hhxoj0YplGVPHYkx9wkuePZMWIRsbZfSb7kHnpZdgF5dRIvtKXw
vQFpeslXtZyKj75JMXQQFv0wjeA/5GjaNGKmW9WsR3VAPu6iqAZcjvrHhZzQoHap
0P6B74t3BsNo8XDS2b3MXq/LDzGa2F0IbEridfXInOlvXG+idyn04lQhR7SP67/d
mG0SPHLyKvvTC/AoOCRnyDM49b30qzWiHebWz6dMb7hrPg3M5nMK4EwPAxeYObH5
JxhPdfnFfgAbFI6KrGWrhABE8If+7xnGsrNRPeo8leaKJo+vvuEQVrCT8Rq0/5UG
1CWuXk5Zoh96uv3FD5G6pMWaGDKwuaBIkM55fEURljkrt9x+L6uXe2QI3MxOXFAv
UBwnzerMJaxvJFULohFJiSMFVgWOOQqhJZxCZityI6kNfybX8q5ubTZJdr+a0u7t
30FhKQJ3zie771VQnFkhBr1IaXAszhtQ154Wdr/HUJFk6Sh6GRb8+YSBRpEGYh/Z
EzF4NiRiPs2R0pL8+yWYMW3EvNhZ126vCscHiM5MZ5lnygZqmmdmDuBq7j4CR4MQ
yBbQwnJSOirMf4Mgid1rBxZau3Szaq3mwAjStiC0bojp4MDu278GQUbNUYANwf91
sEouwIRJfVGASJwMTfeSCKdc8dl0suLU0Lzxsms/CberLRMo6Tqz0BKyYTdF7Kv0
qmc+OvMYGyhW+y+8e8PmCH303mVlezeU1wVEWTYDH8TkRLUyEWwaxZCnkkHYjnc/
I2V5MgDY6/L78MsawlzDEexpTOAc2ia8fBBtQs2kyFeE298pVvxRuF8qoGYgWlLK
WmH90v67QqeWIVEOiXqr96nKp6wtWkYRXINw/dgDoEr5j5NmHAqu1ACsnoKxRs2v
ctUnPznK+GozxN5w0rhG1bTBibn37LFprQ2NVckzy26iD9n2U3FJG2YjJR/av0eJ
cRANqY4w+yIEJ2/iBgfNK/sGqKUX13sFfRA8sBO6qf6wFmAGjPztU5qJTDWjKkKE
1OvW2+h93oIwjQlMY7eV5acuUOr6hGz1jjmZIlx+OdYxIAm1/NFNYBMPsO8GGULc
wIyK7N6HnOjZlKc/o3h5uaXL4aMPd/AzlqvlI3uiYqr5afYTu+AH2xRxk4PAy+34
3JZmFJVwOa1MFg8MWRTHbXaUj4UDZFHR0q+HE1oKCKzYOrONU+j64bJPOzC5RhS1
rAJb8fOoZivfbypwLu9V9vTtwn5/OCupmqpF2+5AsnXETuiwyPFe4h3BYevf43cX
cTw2Cayd4znq3CTr6mjIuNQeGRtdRwVovSJ4mMHYV4PTIT58VJifyKEY4vaGSKBy
ZifsrdlIg3Lf8Jr1gXdbXtglr4vA3SI8QV4tkX8Kmw3zq2KOZ6tMUGe4u2i3QqoP
7qckkK3hgbSlk+MrAdonqFE3waOcI1NZLexkToXvldzCAEHE0HDn+PnCuCvZZYB/
zijZip6On0MgPpLAd2HDXePfWxCrdrCtACdWuYeAa9fLYNKoXUWMnDMW8rd1Qid3
XEYNMLEBUhc03+6FBsavzSPgWPZ+ECZhUFoJ+ah2ftz4xWwJ+la8TOcnyexUAMCV
dPSk+B7Z8ppkWEZjGqrdfjlb5UpnBQLztEJrysY/e0yM/ViG4LjqzWEC1RlfjR76
Nh9EE85hQN09WHxmLRzg/LrHc0JUZC/rK/WmyoROcq+hYjD30gFdvAjDEnxn+bzQ
gE+/uC0c+ZOZkbcsL/kXc8FXJg7B76ifaeimVbkQfGJs2RN4pmYO0dUO5M84QDJv
1mPsZY2KNhb9GbAfYtGKjXNR3eYSwtR+k3Ksv8j+COhyVAzxPlWW2ED+U9HmxE43
pjwLplLLA9FsA1tiCT8P9IIsEbA1fEkbIoOujky/1hFQ8vl+yeJJNMTzH5Xw8RwG
IGZnX+q7uYHhtq+kHDLLqW2qkE6D74Y+qF+Q7fHXSkxh9KK0G3Jkvw7Ij3hR5pZW
aH2nL0iB+6XfFbwDdgVvjc51zKBeRlIXm0OQ6Hkyy//iyIkRwSrw/h4miNWf8YQs
dBR6BOekI+T6r9tAeKAq41piBR/dhqQkmkrO4mobs2A8FGWgiWUuziQlHbDaCqab
8NWKsmtL4DnVlOkH07sdEBwKjLmkhnjCR6K+ceZZAfiafKS8UWAvsDi49tlZGvUz
1uUrAzvWaSQ1UzcLUJBpc069f1QfAvS63JSGaRS9BEuhFtQAU4jhyNWRChMK+zUA
qK57+ayiiycEHye1ETCetdE7su3xrUcSlECqLbv6dCP1EKy0kcBDUvZR/RtktnIm
rVyIER66Xm83DQ8DSGj9dJesWrVSkfZhd0w0Vd/4YG3cz141G+80Ir2+hYGbcbgq
to39RyVxgBHM9FtITkdYFkXtaydcRehcSGtWzd4fn3NO+716vxBa8SpD2isQD/mM
1FOGy7mYf8Pnv2xk1fAyiFifoOt7t3vrRY1nYYxYhRk15p5yciX3jBECD+JBdAvN
on7As3a9QbGEAFxfMI0n1ZHwaS6opRFvDFcHcryQO9yXH7od9jmPwdHaOjEO1Dpk
6DQjA8KJ9cDSnjYox/vuVedMTPhIbMxi8kIDkKqlZUBhNy2D9c3e2cf3nRf8Smph
9TZVzu0njOitkzENAv/e56Z0XYYwRO37vkZOIy6731qHka82tRIp3UnRHZsFnR0O
NS9psET0AcjO4ngjELcibD7lftiykhzfkudMYwd0xIZ/EPtIB8VU5QgNSLLwOxDE
hE5yzDAUtYjaWj+3nxJedklcgiQC2DgEbBcPMW8/aT0HCQuaoF3X2mEOQiFF7ocm
xrNm9xvjoqM9+2pdDviUnrPFp3SV90FrNgxww09xbC+vf3ufCtqTOAlPxZlR9Vcg
8d9vkWBV9Kh6qPwXKFypQFqC+Abo9MZBiHjzrxPTIYphFN21pAE5OjjKGiKwWThL
NKUK3z7+yc5v/HLEhhbcV/CuPI++iZtARhfHZ2UKVsS1rUlOEc2jRh5xKjZJ77uk
/k4Fgx1hAhIgWxqK5juTS7cLTRJIkbpzo8HM6utB2hyJKbLcFqRRNd43S73v0PSK
ETVcic7PJrsTqGna+wbe7Ji+pAAIwIAac2s3e/Em+nHM85WQFOu7EMIUilCCU32H
h0D1HoUDeQ+9ban+1+QCp4AN9RZ08HDuFbb92fKQY6kCguilIrlLCaQNEuXHeA99
VAUZEyqe+8T/uYTaf7pTVTWUcVbeJOd+CYbAQmwRhUnibZv2OpcD+aPj4rS0CYE/
BgpRBL30ErYxs9O6d8XrEwm05uYLud0mO1a9q5jxb4uPR7nl1MAqvoKSZFa06h1X
fg1aV2jwaC2GMt0Dg6w4x39yCP7t/lHQziernCRG8zdvI6JRW/kbdbmLyFMrDkW9
E3ZmTpU5gnW33/B1ckzQ+hr+lJjYzA0Gf3B5FOz9yKO6pfqhYuqwPhCiSnLTbs9Y
tIegHuhj3zK/IjH3IlpakzyGl3b61U7GCaFg68UVaPjUwHPPRu3k1CFG8+Y+RFSK
tEIHOSTi+weooeAAHvo68isanLnGuS6/R08RNuRBKXHXaPSe8L3BFnBOc1ObGaCb
A4V8mep2eTSrFwJBqy6pdA49/epGPUfkK8FuNw+Qbwh9d7TE7iahFY0qfjCw952s
Txd84eaNOutORDNC6VjwIzoYS/UUZGvOwMTk4BnzUiTTMvVrh8lRvvoQcEgiwIMs
galzRaZbhlHXV9xz5iqZNQNMeKYe9Klc7Ccu4Lc3enuR+SqfQelHjBINgTDXuwsJ
XWmR8kXIR1NgLkhs/Khqzm9T7CwUIeDhad8FpISErAKvectpQTrACZpQqoM6gSwy
U2w/h4pBBcHICvf+ODuXZiEipmB3yyGWQGz7OeMusHCqAglnh/XVN5WaprYNGHXd
2I79n4Mc7Y69/XpWJEMITkrMFEk8J58dnCyxTbrs0zSFEjKZrp5AUzUfRVb22Za9
fMocHXkGx4gGkpjonnZ880uoGhX0Hqo1Gqcb4K9eGL33OrD65gIjCv6DJ+hNuMXe
ShC/kuMk9kEP6SMzmcJiU/k/DVXR6d2PHLqG2y++tHimA+WvOf8D0xryqdVKatVd
RgeW8QMQgTWgiOEp3VHPvAm0/Ox3ZyKpTo3Td92GnWylQZn2n+atWf2W4Wbn2yzs
mlZSL9hoJDZ+1YdihjE+GUhNK0Bh/HPCwzh/YMOSoy+0s9RNSpIugeFDV+3LKDTa
LW7FaAga0FFwD3kViSmTKbF1Z6IJaQj/zB8yq3zTk6U8OmUBQzEzq60K+1EdnXi5
QGSaOnr09OO+FGSY+rCzHPH1Ft1lu4ZBCZoxxu3+t1JwIbuJCnQZWi+nANq8NQ61
5SsC6NXJNWIY6cOyUYl+Siwft+CvLGHbOVYko6qC3pvzxWqys5b/+ll8/rCVGB/y
GWpVd4iXbQitRaAlnD/JIVMAE6Ct2nQUNOLYlI4dTzzAkbxgUNx8VtrbkFS0KkCG
JoSOiCOZkBgC4LtHmbP+FEj0H0CLnDLqwHt0JfYlKaZLdXW85tDZsnC2+i50Hzsj
AcFsDNC6YBE+f3mJZcybOH+TCprxB0IP55smiCKZlFr9jHalx5U0sjVQkUG5WcCa
xHxf/UGoPOkU7y4rISMvnzNbBVmsXCYPvWZ0in692URMRz9JUHFvriOGlNHAoN5F
6ncOJ1SiIvsjhvcjit8ButfGmSTEtWCO5gY2UiY8B7ozoNE/3SQoRBohwfIlw6Sc
8dI2Z5m9JIORjpbREHSPAtQo/KlEv8+0ftBFSr8xlhwsHvpJgE5j5Q/DrGDgltKz
VXany0rMHB4oJNzBEM/OeERlTQIgAKoacN7+75Q/MLjs8eCgQzPp9yXbw/ry1VBR
b6EEbdjj+dpb413xGLaCD9oxtWEjG3ot4jFATBpwRytiY1H9pBtdsVvAQ2zkcrFk
MPWGQ5L/RP9cQb41lmsEN+zJrebEP7lq/sIlCbnB3GEVvyjy2OiSxhXcZlndJNCV
EQiwcZeK4K6tdXH/2l0wJIsF5wUlUz6Dd+UFLSIkr1547JGrijmhMqpW3CO2x3FX
LiG8Sej9U8aRZcG0CcFx9ufbIeIfW7Fe+oTENoZ0FVGyyNCh+t/3IlxCv8iTzaw5
JSHan0dh95jpvyGhZrtBTNZvW87acyodO3W4j+WlzUAektbq8o5ZZMof2GASwlps
HfSf/uQducQwJ8KQKDC7OaGRwtW74CGzCEnuym3gmN4sXMSyDyV3qoZ/0s95tnsg
Yiv/r0cwZhml2+d8sE6r8O1raKuc2DTLCyGzol8O8GbcQSag3eH8UndWat7okEDy
Txu0gXCOy5Wpp4u0FAMEVOjMfnwjB5xbfM06kZT7gX6NHOIhDH3fXWTtMEoLX+J3
S4zmIuD91ttaeay9Oi+03yH1OVKWcZmzcT9EdZ3A4TE7ikv06TDll9B65A4hMLz5
qvr3qk8TQfN0VWks2aOq4czc60dJJfdG37s0yE5aW0bKqe5k+6QcNn56k7nSdwMK
nCw/SOUNZjyuIRBs6a7qQQMxpceffYAELd2/g9RDeD4fXv5JxiHwnt6wFqi3HoUR
U7mv3153OkToTafnqnP4bIATZM/9TssUdZ6zSPJpjbdTq0EQuXxXOVF1BvhVhonX
oYyBLWC4nEJkww5vJQ9gUI2R/fpRvGgpBN/Ty3Wps+spS7GQ7zsYqSgYaMNKJWVA
sO3QCA2q71kv3a1efexONtlap8RGfMw50Y8QeUjxLYhRplowu8UcjK1fYIdwn3WC
1lGWl4I1CN/MYroMrbJcOX+7Xh3gqL7zw0eC1X2dkmTQRO00hjqqZAM/NiFnrLbW
oisDGYzPn5NunWkELwEX0Ucg1mMrxlmMhpTI76hfDvaSXaddO/Cbqa26Xf15XQpn
ChYvlWrHFn3NTaG8sLGaDFT26qZ6ZA3Xp/j4tSRL0eFAVtuUM1mp7A0o8FQhlfsO
lswREh5B5wwSZn6ucdOCCraXU2lIRTtzOAHRiA7knj+v5HOsyrMuV6j4+GR13Zl0
EXF7Z980AmEGAqyTmveQJrd4lN7GWHMhsPDoDpuNsTcQdZ6FN9OcEgl16tf6GI7t
Xfb3SSsSJL7PeCY/LPbNtUtwO8BUWWMOWy72CdYSb7VqAz259p36Ddy3/wqGorKW
4NX54OyclWr3Mfua90DoBMQ+4oQUG2Etona+DYkC2IVcSk5FGqiPZx27HkS9+zbw
8CRiFcVpgq8De2vKPsjg6phlJ4l9PezwEJO54SN7+c2Ixny+PI8VlPNY6G2rGy6I
p8ySqsBX+RbcQWi9h7XWaqZdnVurtPvdVMLJBQU825TKO9c79Uj6N41ca+uMW2o5
IqgWpo1xhDnYus5thazlmK7dOCWzAxvKw9N+0clG0Rk7/PutnuvmEQh5pF1kQrCR
Q/e8F9VdM2sKONsJVJ4Cm0bBuiLJQoK+xQG5PI/R/gzpwPwOaXVXvT9syXSj5qVK
lMLiAWqGk5bd3sbbKjkiuvJFjMyxTgj0ZW6AFQ1HXPEr/C7a53rQ7Mw1FS/E/i2z
iV4KazMJjSMWBvM5VvBEhQ7slvGWywzOPHKnygA2P8dB7at4AtO/+FNq9TrAXD6C
9w0mQcoNlrHkc4SjW3g4Tfj0Z6WIVHKcLz+NqqrkASLu69RT/VsmPxvUAMu3N60f
RBxp3LrZMOeTmpYn+qqdLSrbyQX3tUKil/oMoEccu27SMabJgoRcYMWi4LPjInvI
pvap1qo73bfYpqCaKP8ZgUDG4lsYXoR5rhwLWQ5mIcGTnlvZaIbPVnUSuGvPH3fo
mKAJAtWJ/v0d4SCq18OMAllcGQKzYTc3WFz2zEvfV1xap1/5R4ZuKv51fJ0Vv3F8
RyHN+vUoKzbOaxMQzXbL4dEq01C3bRnB8v1RgnFLEtBcq2dQMckbiSXzNeYUg17g
Mbq/6tU7NaH/gfq/RMWPTcf9EeyCyQn20aWBB+daGJaodJNuZWRg8K1vMYGreGGe
b0kB9bROiY+HXKe0B/Qgp+hdaCfBAVHafOk8dQBQplaSj73ffQr9alOPFGPN6v8s
wMTXvq55y3OW5YJmZBHowZZt/Byn7jf2OOxXf101rD2Dt8IXBHAeTLbOv1naKE0F
zkGPfL6uw1c26SOUGlDu47SQ1O9tKd6n2jPhOvsRKWpD4t+VP8VBcHZ+4qLvsNCr
u74DYpK4ZQoxtBsbNI4mwBXz3AKIE+kX6W4LIhXi/L3WaaykdvGf2TXv/aUa+vPI
8g2NxYoi7er3jpe93RKjqhc7rkInhNdHL2A03o3XWXKZYi2F0RAs2bkNa4XxrI4P
7xk5zyvLp4iCnoQdXzfsiX+PKpLbMh0x49lZNZlfIc3+P0RCZjOsObY08FYlHLa2
SuY3fqSucTGxwlRc9BrJ7c8Mgqs432jfWyOwpSrCyaIA9iEv2u+y8EnwxMUKmM3O
TXJZr7I/b6f0ri3O3RNy6NszmTR9xUr8kw1oUSff1PEyypBKtBqYcXnJk+H0X/yk
bC5JfVULSkBa7aACcibw2zsIu9YbShj2uvL662AkbfGk4+Ay24cTWcoClovduZkt
GIWUcsma8FQS8xzEYsjwrd23pK3V/FV/XFSVp8y3aUGgs/PXE6YEqdAGKt2TvaT+
J+FGTtu8VMMF4eQpXSLZjJ+FyY7hLG+dvrgbtu9EGZrAGV4fjToJaJAcRRfnCrxX
Xb0W8JIpxr0e5wQtHyVnyvcgQOCBhcEKrMFKqxJQd2eJIw6MPUDTlPcO5L5yODAa
Q4mqhoGBDS70iRAHlooMzdgxIN3BlcFqMxGIPW7kUeIIOgzgErSeVGc6iNsuciD8
uBLf0aZeGgAG3bJLYJ54lzjkLzu8wUbdT+S+F5SIG0+JEi+m8iptLciLthvtV3wt
KXMSJOy065Ah434TFhI1+cGd0GqZj0r19n1el3wQ/kctPF/4HJLe2FlOnm+wOG16
MW8oP09c2bIhzFV6ft2Rrc80Mwk5PNtgATqTVGQzATsELnXeinYZ6hiCwoYztcOz
jaMf7x3iq8xLDxS/ZgBiXdZT9JwQRALpOa2V+D5eLHxmC+YTGAB0hVtvzYuYXIt4
82tPAXeu7xvg++fqHelm+I/GbJPF2w4Pi6WNqVOE/iYQjrJhMSytth0zfdvw9qU2
frk/q+Fr0RnNA0d3udZFOPyT7/bXOVa0NwOx29LE6CNN01dyFpew42RrepwImQhK
l8OrbN+tI6IMv59z8kK/XlehYImZj4CXczHd67FUkBIxsxq+t+Spx5QyXrpdVWTB
1ZsDK+FfwFvUY31C8f4PN7HLI9lVAihP/IzFO5qem7jSY2XMec7AYGAqsETzOeJG
etUixtXhBe9J5nylzGUhQEO+a/mxaaCB5Z8+tznpx4b83H7Uwo6FpWwZAxmIbnsJ
gjeeUpqRKudFycGPVmqiWTyFI3DB5HE5V/uJC7DxhEHpWnztnAJoAyAlKGjCJUs1
bgQo1Bg9qgUr4r2fAr4r8D8Hgr/QY8TVUFMmGArcEekBbpmvM0y4ZpQvo57GxZ0W
EQm569kb/DlBS7Z1hT/GoT76MoclItw4sthyw1DpZT7tezQfCek4kkDJckjz3Q9N
knbifd/WbYrfSW/aJF4FmIeu/VyzW6XVSQdOgAvuRFci+tNcse1spx5LDIwj7+Ir
JDT5myXNHS55t7sUd0GrlEXjNAGDFil2TCsX8nnFp6yEc3YH0ddUTY7foMsrW1Fn
eNorjcvjuffVjXZWRFRHWyPQ5zabTtfQMbPU2tDH+aobPBzH+J6hSrx2WohOdZGL
zaPLRxD1o/IgqL1khsNXp9pjxn81m2DxjC+PS9wXUcu7pF6YWHk1XViC/JOHmeJH
Y0QEMss7FNQ1ANwrRNHVoorFUa6oG02u8tO47ePH8FjnlXerSa/RnnQjLwxNv+kJ
42qhUKCY0MexTCZsXkQ4JdOr2abjPx+g0pzyjsiOYCOONf84sRMxKjgwxDahbcJw
XzT9BojMjJnqX1fR/GS0L4n0YQuq6jCescUoZVSgXIN53WK2Y8FMZmMuoz9DusRz
9Wfcsn8XDxfZLiVx2RvOvmKtSLxEjDMXFqQphkJUJfJfTib3RKKLKB3ecOXHC0Vc
CgnRFPQ2AB9LGBhXtXkD7hrszAqG/R/IOtM12QyooulnEYmpr/H7MkvIqMKZ8tpH
wvlM0WiMvJQYkeTfISZcZxBD0ZwC6EM/GMhvW18mSwlzyHVJp1+dv1qel5hBXAvO
YssVB7IdAVBVnhAIZO+w8fBctdkebOiMvPjcJbzOhRhCdoTI+67tCUqaOeQQr3YR
q5dQLwWqbTkCl0hmNUzL9CmX2hd6kTUnrDKaGxV/5IHJoTbtuSQPgP0oBZ9y2JPJ
5pL6kqT3X1vxiWKxGfnqJxF5CAW/bvs89DBS3UIIMJZcz4fWyvu3zchgSOD4Ltyl
V7AkCH7PCMN1H6cZFA29gpDZ7a0BpNB6SgHkjAxQjD3OJI8qUVgaXDLZ6JS7hQGC
9+fLy3cN16bAtjAAmCZlhyA91Spw1X4+Yi4BgMQniSUB65kYpU5xE6rxZHMFG43w
w6fd/2Hr7Rg5G4nSOfr1ICJIFfKBygOANa4vsc2Z3r9r3Xlk2eOnzImahd2vTaYp
rzlwPp+BaK/6TB0GykJz/AyF7n6Jk6eyfIG2txZo1LKmnEdZFRkg07Crog5PkK5e
ghleSCNU+3AwbCWXdvhjsq/vozhX8OYVFtpOx4+Eh/y+gROhephV9JrBB/u5iEpg
It4yrIwgt6qrq80go2yJ8Eeny9yLyGm7uCjBdf0byJD6LzMXLt6BVvsuWpaEIZXz
P6cgh5ngWOV/Lbe4GDWiXHNoW5MR7oid9JWiNBsNkmNeHXZn9nq3hCgPYLIDzRI0
ZprTTMQm7k9sywV8kes971KttuhSXEHFQ/l+B+zuQISsfDt25Bm9+gj89Vo4T+JF
S2SDF+fiWbfPBVJIl2wxyezpVjJ0yDzV4DQlBWth0QNgQ0zHEDwYoy9BOX+LU41r
eGIs0Do5++YguykKaQaACfntSvdVmliZ5y/zmOVGgxK96aurF1ttaBQI/XMFBjjB
UBecvWzhEriKxFI2dpdUJMQWc8YHwht+54dPV3vZ9WD0pV64F0yZ0IaMddjadRI3
qQ2mD14uQ+f5e2uqSahp6E7aR19AXI6JzwyQlzQFOgUuFH14iHOGHN7gUU2GRV96
rlyb5dGWc7oDz5jr3pxtZjb7EciC5HMFn2eH1qzlzmolOPUEfMkQehUbRcGXLYq/
mvtj+xMOxhQTtSrzH2N6YPIwvNKBUuKD3FnkvUYhmTTP9jhq73XRPs0hOA9AAEqO
aiUx5Wjiix2cLO9vU65hpQE+2g7+m0Me5JppAjl7yvmK0ibJOBcPriEEnZU+UXBi
2q83r+QNIptR2RfgVZBizaI6fBYLydny61/WLk5EPHNjk5kI/fy8niKX4+nxBGkI
ePLVupRnRGr58SjX8kzrnJzd6BOeeHD0ShuFX3wXsc3nq45KPb4lqk5AgAdpjn30
UQ3BZw6MGcEwYkVEdoGCyKTUOsla8FgkWjQWvU9ocdE7nCxyTlFdKNbzuego6n/Z
UQ89IrLyIFAEOMED67aOFAkq9t6Wfw3JtHS26R5HliSap65EEcEiy+ma+9DDbCP6
ABqJDOClLgopiFjzy6pOxZ5kE+z6fAQJlV9MsUITumsbaI7y/h/tL0Sd3lwYHbOW
DM7fZXu83Ch8DnCTF67wpU9ZWa44L4DPK5zLx3UAHjHbcWGcbDXsmPZr/QJYfSk9
OKV/QcxaTX953AWzR/v+iKEb/UmX7l6c3EV8AxdUselqgkzvBmG8SwLF8XdKSuEi
eJ/kEj/4XX3sh833CBdHBlJEQGHgwrGLz0pMYXIPn2bTCbRF0WheDaqYGuR0bSje
/Q+eoQ5Nhyaj+HXpawV1Xv+Ge4nLfnwqm7mi+P3cLxa41DUp70KuBzqJdyxUZUsH
/E2ral4yTvaY6A4XwkwcTNS8ViIr7Vdd71241lhdWfmoZANLAoiSptqpcqHXs7tF
ZzH7HoRXAfDIautRagsEJGsC+yKO8Q/0H/lvrqe36eC8x0YKqBhukZl6hfLcdjn6
Mw5ecbF3iF9VnUd3cM8iE1B8ud1MF2Hq4PS9vFasrzJEFXvs/gMAotezQw79mVI+
GTQu/ATk3kO+9Q/l/JibD6692EydQsOdqUUlblaZxhgwK10zIEvZV95GwMTrzPUE
SqlrJPpfCFizxQM6RIpBig8+BySK4qjakgBJw1oCCJz5bll3WtDeJgGZ6CdBLTzB
IArOp2XQXsvo+4cvLQ/q8Ua9Mxi0jfsC3WmqwOLM/eQIKaFs5P1WorulalY2liFK
dQy6Cfd4nqQHLsnW/VZ//pIYWmTuHUnJ0zbeEAprcW5nPslgKgZ5gj7K4fxlSOhO
LLDujG+EKeLqXbTHfx0uu0/hYzyt90bhYJ5DufTJub+b/w5O0k9UwwMMQf9PIC9G
aw1gNbquOkwl9ZxR3WNlXOIDl5hArXzO8SbfOU7k33uIa590Uyy/uEjjj94YYZZh
us67RWUtIFU/9a/kcmNIBdIvv+VPgSI14Ezq/EVrF49zTTyr39I5kcM0HZn8642k
0WsHOOH4ldye5cekkUGxqkv7Ar8lpCIjfo3vcG2BXeus9qZiQ8Se9e4CJo0G3vwV
CUozv50f21ivqdLz/I+Yrb0gul/ebKkxXx1nOkdJn+MYiWAPr2EZQlqWFn5RX2Di
beqkct2hWTY7tTZbUqQz0/f2uDWxwUzOIdNOzEYCGP3ExycsvzruxojAXCMQ/HTW
ckqy5nSJV6P2+EI2Gw0aOeFG9zHTug59v9A98DpX79WlBGuQcbAka6Xa/4tjCV3v
wGx+hC5oCYfuFpHd9tGsgikHU/i8gSX9L00otM1N8ok9j1eGVGEHQfDE7j1bAhm/
kGUy9T9JtXj83yJHBn5Qodei2E0wH88EbSb43R/5N4w2btbGqqQwqhXntPXny7oN
tsDNRaTQPy1biE4vsm2Vat7qeq1iVaSS1lbc59K4RGxPDwxclgJRIXu65KyVQGT+
YQntcyNy5oNG3fcZufXXA8XH5stgwThzuAgcYdpr46M4SOO92OZR9CYJRkHE49Fv
qhi/TfB6kfJL1W3hEcczr2+HAGstV3sUb246i4rUieYk4YYR1iU7m/l0x5nINlBd
nUUxsFx9hG6RClu79p10Ew+ysoLwoNmIqF0+S1eObaQ4qHjBKE3sJGJ1G2Y661fl
ZxPRnf+ia6BPA38p1keVgO8swyII0BJtA6cka+7f/U57FlcjuIVaBRDof9jShLyN
dwxoBKx86oHjmUrhEn0fIiFQ+UDjzQ1ZGwBto0mTfQNfFyliO7k5K4gy48yzIz0/
xhHmTWiqS7zLkXIm2WObFXLJIUb0AxZxqQAaEbosbvg8iQNkzqQwOJ3y1Lqn4Hu5
aWskPz3SX3HaSsfUefyRav7+gBxCIc/JO95deDT+UpCgKgVbMMfknYJFJeY0gwF2
uIX6VGBDEcYNw9+Y+vjH95mbE1WY9wnqm8GBd8byk5EaqnEzh4SxOoBp2x0xyF9k
+MS4qWluqPC6rOcv7qgwkRKltGOegfoNIPlGUubFKkyexi7ex5UkU95d9+bcZgKm
+iNf9XtxDwGXXU3PJYx605noVVT7ZCyGWvF968M5EFF8AueEhMVXD3EaCQ5GXpKu
v/jgvRDqXZKazRM78U5TWiKfj0ebd5/nMk/Cdv0s/uY4Zsqb1BpL2IIWzzjTdRpE
0xLPQbCpmh7qpFaWprD7CoIk6WcOdaf477q8AAdI0Bp7okr3Z01NSnG4I9m7CSgl
PW8B+xWpGSof6+MeO0TUtE+eMfENGDtMX0S4jyWVKRXTB1avxiYaKEtEANQddgSu
gv9p8fAXjcxjV5+VBRZaCfB1Wt/L9DIKr42p/2xcvuRefscwBNu+dXCHAmiVPwCg
jZ8BV5b+JOzRVRqNaSuyNQNDgGVYzbspY82C8nOKjSWOVwPxIGLuVytwIWVOMOvh
LQi0zyJMiCGmRjtyzrqNgcJt0YTzgzoC5G00gZPbsNE5u30NHb7YOgc5DdFXSn38
K0tquyNNbcK60RYV0HDHdaTOvQ0Mntu5d9rUFdUcx2Icp8wlzU+fDyWDkqOVS+sk
fPLdZ5Pu0++BfKN03ulH3qSVyFYoWh4gSp50T87RYJWf7nUHdfLfXaLQx8MkTxD/
Kqvf37iQs7oAHF3ykLg5qTOwyDLJ4G3l0rSLwtY6fKYdac3C0d24EPfWSRUAcknH
24NAP4M2yCKZ5ZHAQYHD8E5uG6q249Y36tX4l4gszVgDEXtILC4J30gyGV3ONBqi
YNXTm2559KITMij77P0JWa7QlN0WvDWA/rify50WVPlC5IeuR+iNOFRVWbrLUslq
WfX/W4SBLhUUDbd02PGRieTtVrtTEV0inJrdlaH2h6idj4veAHhd1R7ADkWYi0pR
zNGVcFFezSnr647qIjG9MMwAQEHIwJ7MLQyzPA/I6cE2CvLUm0hKm+wwT8o6mQbe
qvYQHPSnowerlF2YLJden7loittOXd0fHs/U8D7ZrE9K+dr0LAIyhL76DfXEtlDZ
RtDJW/JXsOuuWQz/QAy4geIR7LFquEmJqnT7Yka/mzbMCrtSx9Kkaljo7t7u+kt/
8U2D3VlCy1ehMz1eU/kCRfiHkTBlcc5/MLhQSbJLqeGJj5+TtGB43K3kKaqbeQwT
JcL2cbZbWXKRVWDAEQ5TFMorKyFb3vfYAjHYOrTuMzCzdfzDuj4nrlNWsJCFKt7S
HDSkA1yKIlqpTW3pGYGHgNT2QfqJyRW1p1Qd6Jm+3NGnsxebxu2GZGFZsDqQFonQ
CpBO9R2GqVxfAczw982uBKmkWb3dfxH6RQ7FKzjnZRN2809Z5XqYx4VXMx9u+lV9
XAgfzYn67sdolqJjQjEjGOQfjEuOYXvLOpx3JGZgCLauhLDe1uiqokOCvVUfdNWy
Y+8mmbqG6mqKrvaT2joR3JXMjsoocugCpFYbN+FJwC+UvTz5DublpCUVH8TL9Y6B
KmunOgy0i34ynz4KMY2cVcUbAR5Y0+BGChLNXgQygiJsyL4OcyGgDUgRrnlRSgf3
Pc+VPTUV8jLqFtQAk+etIsOL9lqd7uIlaOLWud0TukHZBimv/jTOn4m7lUIvd8Xm
azjQqiRoaLDUfmqicbXEufK4TeZEaxmNL1RBbE4axX7+s+dec1+TI+9hDjk78EWO
dXQe3q4Iq2g+XwRd97ewmS3rLqAio25ILPiT3ppckYvX8Jdnf6GgjPo58FOTBUS5
gMvR5JXT5z8aAnuxCEq7k8MtazzyOJIUsLsQXUU8krpFsJioKaXfgTpwbOBmNLqc
STgK0ZPuFcyW/f0IFckausdcpmA4xVrwUUQPPcIQPGvezltyvOGtb79UJxSUV/p9
HcVn7kSoPSdLml6oQjM7qSZkLpx6SMsoKunnynI4TboSE1nrTsY+X1BC2SBS2aa8
7BIDYM+iIgXavbkHGlBqp4IgiLAMug5LcS+n1M312MuPve+Su67DnDm/vD0QrRSM
dcFTzjh1T9Wj2O5UTgrN9RtPKqxdWRMEcaJp0efakIq4tXjoVwB8qSrkRdhX08WO
2MR0ZVyy1eaQZANZWtRhBSnYHiIzpcV4883mn9qxrkbEXrVzyEDJpNeR0pMCR1PQ
sI6UdmjCdeuIhX9ahUdWiIrXtHjS6OAHh8xkyCEpVLh2Fe59XC8JwfqkjlLHlA8t
vAXvG85dRn3pCq8u4+DC8GrWD59/r0bN/YZPxbNpXzVL4RTWOAewJKOylxye7DwR
epJKBzlfmv9SfQ1sZ4aI9rOCNkXw3ub52zoqjWQpENU/BtEL4LPXQvM5vlkqsw7d
8uWMIelXCpJUUKvvXh/pLgKxRj9xPO/Dv1hCG+u6hBT5xSMuN3ZXNKipEeMc+2ej
0NH9+DTUwtU9Atp5npCVFTjhqYFQatlQGgbt1VSMdf9Dekq4nyVAmvjC5/1jWhbs
plhElJT+X0i8jNz1J11Xan6kvV+MTR+8K+FTkiZdg7X1H/tCBLPwfmsABFXCc2c2
QbakneILP4LdbB1Wop/F2ibt/5egEOmFGagQHOOrT7xCS8GuKCEYgHWJnz6nxXTh
9zkslGkaBH8FZiq0+oS6eocYQeMMI6O8i5wOxKI6Vjz5qcjNnWUVCY07gQ6jg01+
AEnaRF+ezOAIsNA38JJCsYnRjJnSDj3vCeK+cTPlnkqFJgk5dRc6oyrv2CXZGlnG
vJx45B6uIv8A//pVWhDi0quJWPztm952g5KM9mqnQTzdFic+PVAEoXgBcu3THPsu
UEHaAp9duaUrGlhT2gkw8ocTHcmxfK62zG+mIJgB2oTUG18plmMyJUZJ55sG4jAM
4j0HS0Hju83F+pc0R3/zA2smU0smrrpxhb7IchMj54YpUWKDzKv7LLPe60ZBnR1L
Q88tk3gVmrqCe+yozhjK2qWXHgg6++Hv4fQ98KXxlsjWIWEYdyf9kxZketR02icZ
vRTvL3yn+krQMbV63DMlwvmyLh7F+HpxXrENJS6g/JFEfF8jLq5ktdBAmRh78WGR
UwKb347rK1RG+rYkef5Avb7LbYn/N13LwDLkoXF02tJKpUetgDuOXWEZWnkoVN0I
3Nsv3hJg2LdnP7CHMXtI9gXyCtMeU1v5d6u1nMT8ZGj1yExDLXiQY3STbm6x+ISi
IW2HHXuE5cUpJEAXtOItNuz5mkToGnfks6pJ/82zyCEIBkiva/bsdw9z2sgXw72x
N1Xk6A3IOmpca136CSyXmsOjDI/rn9warFR3OMrUQdgYF3RzXYKs0O2K1+kB1RN9
FtzOTUPxr7FPpu1am8Li+F38/b09KAtisaS0cOUxBgQMd++/VTn/4j2pJ2/GSM0c
jdF1b53eIxT2vIzbz5Sk1oGHVKIlhLhJ4iSlBfAYQ1DJtHFuqMNcfe/JGnmBYzFy
/xQEk9jaXsJEI5bilQy9jr1E4BCP+fHuFwrO/DQ53jhP8Jwbh4w9fmHha4y2DYKk
g/e1KzntOYdCAI0DkQZoxeaDaDrOy9YyO5S2N9IsLbNaYzMcF9IrCWKckfO9YVOj
YwazLLdJ/Em904zZ0w0fD7SP8Cg6pXa1YhJBhMM17wHIi3cvA8lIaFkV+N8CEgA/
YD5EZvnigk/FpKChd1k0HjFlRKAbNZW37pTFuNkjVsUcdY3hjTBi+IAX7zY//8d5
ycv1++CBiujrH04wcWhLgUckGm28hkWgxGmd49FCzajeJ+fNyDKYVTV+ZufY81TT
7I4VzbsfCgI6jhWDgwADV+rY0aaqPremu4a9BrPxP4WidEDzS3ipKPWKmpe9pIaU
2HUUIeVTgsCMIvp1h4tc1C4PWvENFIi3i0QlmWl0LKQkgX7Jc3s+F0OuhuHSx9eb
dCNtMw8zuTjAwYcmJqSUtF5tAl88shib6ypmXaGnh1JcF+hisy/EFES1/AKyw+Fj
F35m4gLBhtB+0WPHAV7iHSYIahFfXL9VLj5JBjMTJOrKjbOpPFXD4SbTHKfQ42QQ
arSefLvpkOfbhLrfgGwXPk+fOiHG0HNGIKz5UVEIiQucWlO6D4JL6xmRFiqot39V
XRHZO/1zx9b3GsVs392J5Q8PRehSfgBvmKObX4oKldtN0zTmE6BAyKvt4jqdF5IQ
F+kqv2tauFoX2jjj2GYjeteH8ig4AaKtaVy/fejYtQOsWuNGkKE0aomh+zmDxWj8
X1QP564lAK6y0WqDeFkNXb6eKTCsHXYQcuE1+ekGseo9Bd8xJQgtRsPnDYyKHfG1
SvvbSRHqyDHAv8FkuDWcNEuDJioJZey6TS4HpbHA3xH/fWsLaq6oaAtduPSOKgra
BwJgDQlPJ/OrXue+TXPRxOeTy0fcGUFB/JEvIqHMXlah48oeKRXabNko0sJwSPEj
ofDSTrp9SMFXjrpoL3LY5/ZVT/zY6QsteY6BBtJnbanz1IN3yzL+UpJ+Dw4k/h1k
a1WPb/FQeAwjnWUh+fSyOI9LNfRk1yl0/XiMG9PCzC7xemocKJFJjXjA6h0HJU6e
bMVUvLmzm+L8dpGUgKwP7bpXRagEhfOdxRxVKhzeKkWvwwamVWBR8tSnaJveilXL
jTmaF15OietauccpRV+UWoBa5veT56j6jhvfFIg4PFyThSEAPLSa0741JSUrBOKT
uoClR+9UzbFtSc/lO4nw0pFk4ALNKDq4XDYFtcr/D+5i0oqmrNnoLW44sDDLX4Wn
TQ9rMFfE4VrI3bmrNuotbiD/gG5NODNqE1tIrHbmgA8P3Ofn3WvMmnwCkg+5FZTE
AgtTLQvJBhDNOIBryQdlMBkGICaqRQ5eSY4+2VxJAj7oBaB68+Z5tOCJZ3OkiQRB
gPRnS6ueI6JXJUE4kIrRp3E+8L8ksNurLrPUuMvPXFOrMbGDWfNW2CV3xvdCNKsc
m+323pd41RSIJhBlOB3bAn24DKXQIMu+GcvzLC8TyCYPwasakhXb9jDzbwnS0146
dfXd8aX/ICLM21l5r1GWOWwrpa4SGrMsybJuTzEty4eEIViTzR/5ieGtao9dhtp4
j3YOPBONdtAJsHDHnnI9Ei1VK57Kivj4Z62JYZKsOvhhFkL4MdQ92kMeRIrJ32bB
ZiObQJsoxhHLzXjAhmSfa3NukNG2L+DhtWeUGNaO/q4mnzyBSVgA+0OxaVDpyv8D
Y6YbwDcihou2QrSfS0J4x18/atiQ8uD2QmzLm7ijcf3QfCcpnB4N6DC/t49Zq1c/
w+EInRzGuXJv0hGOas/k1PbPkWDqfWMXbDA0dl0FcW26b0neGMwBKGWvXyS+Ui2o
yIkOt9zu5ssQTKb0dHgfyxjLb/095YqnwPeC8tHqDna2hx8QdNeIrL1tkxKiPjrr
gUmPGT2C/BRVlT6mALI7JbyQmi2JKQHsB5A7LAwr0NlwiIqmcHjvMXZVMqDx41Xl
B1SzU4d424wVttUP1keN+vYw1uXCwODO6uQNPxGfFGryQly4Jxw91fv5s65MQ/wy
9itWFTaezmgpUonC2NmWv49NQ1weXgPhvOoOg14iaPUvsEjm7H4hpB269kUeYouq
1ebolIdZzbaSbwDEYmlUHHT0ntuVZIVYG0XCAo4fLXs/xXXv1vFJ7fofHUviPfST
BWuQ9eSNVKTQ6uOGm6N/0iX/ECNwnH+zezYa7EZq5mHEKLTWF8BuncV+lZ1pZ+9v
U3J6/2+HlSmhFyGbw1ZJVHZ2/oPJpkC++Q/rSoPY3vCbbwI/XWCGyw1wHZ4M7c4P
SXGJC2Or9xOwaZXODJzZ9HB6ifbf7hu/6GcgqK6EFg2E+FFU3ktEEjdClYdaD+1b
J/ojQQkXgTHxi70N7isz/TdCwgkfXgfEAByiIQdFNr5yuAaIC2MCT8ZmgXhhCnqx
kBYyrY+TScLCRp+MVwCuTmJ8y4q3YmJfvaUvIhEd+/nfJ/ouoaM9/OFbM+7EvzcV
/0hrA5xGRMlrB3G11JmIF2ta6UK1JmOQNEdlEKkvG4RwIMIgJCCCFZjrO0aWpld9
u3AftIkw93C2MX9K2qZkGmEwrRoOMc8pbcBDdcp+m32WddvUev2Km5owo5hlROBO
U7qSPM+yfAf2ZRowZ5SxNJOSTxlBQjtgYtxdvHQDwot1CIy80Q6VKcmVFIR6g+Y1
l3KSBpnxDAKGHnLTTiqQE1h7UuAig1AVQvCVQ2ucqpGtQI9pdhv6ALOKY+EZMP4P
s+i6+EzDnb3a7QjI9qUzlkWPIqPXMwHyhx5LGyXNMW2A4t3kXDO7KqUYK42MdzTB
BhJWMjXkrkQE6brVjem2vNdrCERCVzKnSnQr6txpgFHsyZXlJ/rvTP0U/lpZhB1R
5NbwrGr6qMl/gj+wvwm0UgfvOvRZ+EkVCI6Tkn+dNbDzra8TFu+fWUgmidQ1sPBT
pys+D2klFvTav9pcBxK3ylclETVYcyLCJYIFJWz5r+JFMO96m5jyXLcVCOJCLbbp
+2262jLIDJn1Zd+rZ8BJsF5wwbgj5Gfpk3qKYU89+zzS2hyz/lsP0u5eOBvK2MSp
JXDNd4HXJ1iUzrp4lXYq0TG9Eha4EhQDaGlrtMZyXWnYEV0dgJyAtlOHvuyh+136
ksW2OSBJPh9fVit5mamFa3ixpGN61SP2uXYXdE0dr9nX8XtjpH48Sh5/6q3q3+2K
zFHlCYM+1HSDgbW/YIQFShYluCzrz/T1yoxmMtVsmhE+vlzJ6BBm3+iOdP01FDHS
s9KDUeC+hrZDbf3UkS3ZdEWy1OR3PFnXFrScZezMHZTlF4BjKpql+fLHa4zoFtce
g3uFTMCatpogGR0aX+AFBpoS1YrReImQvtSs+fD03IxRqZDn/m9mybYCrZkeYtSl
4QC86uDQDuUnrmJJoSqZ3hg5jFnBEAXia4xmNwifJahF1dTYtEOunVoIE1pCDiBn
dPYDx+RNBU2ubTuFe7Nt5kEuoP+QHSJGgCu7NtJKR+sTumhFMnsi5kTlGoTqgake
h+UW7NFG3bqM6JFVRAfGDJoGh9jy33bTzWbI5k/3qCfpbW3Oe4uSzIJH8IfWk/Py
lVH9kPk+zY2YAi+OkpYDelaJTnlZvKyl3fMSQG/picNRj+dVLBCkl005dVy6TGqM
YtiFXhLeaDARGpv6hp3F+LCqECWZLfQSZs4tLzMrxanhp+1votFj2oM7LEian0Nb
6CQwK8k9JNSvJ2SQn3LP9uCvUuS7XbQjzzhJbVC/7r3HaO+hm/nGP6hDk/rZfbDC
oCO+8w5RhU+CsApZU1Da0VUdyQaqMzZqG84r9E45c7mj8l+ejo4O79SnC5I/oKnh
WRUidj7WbfX9SNQFrte83R36gE+JNiHA/E4AxUvwb+1DMoqcL5aMpFCTqpdqBrbH
fVSHLQaBt/Dqh9WcSZzX9zyuPIYKgDvBvrRAL/IabgAZPwxlgNQds9+WO5lERgnS
Q6tsmVYjraR1YzvIaT1UF/ScqrN4TgnXjdufrr/FlOlAi/vkcOv2/c++acUlADDz
1KhEL5A4hw0uFQRRzucDehcG6Esm3Yc0GOc6Pou3/hLTmseqPkZ7QYk79I6uwMMS
rmWRX3AAscG0s9P9p7Qw2iac70BOvRsqSy62DZM08+0X4C+iovmAiNYxuWLXPTf3
CG74eAePgd1h9uXwpUw/DYemZJzSuleBSZxEv2mZW0W7tTsp11ArNvTorA/itJ+G
KVmrAD9aKZ7DWZ496sAuo+z6+XHXAA7j54oEzQk309N8rBRBmJOJ2rj0jlz3fm8r
zY4z0wySPpMdNDmBk10s9r+uWPo32FD36Jmd2nkuRBQ5LgMcIWrrSM/rk8QP2bKa
w8w4Qldd5KJJn1U99j0GAmDW+kETTrsKJpMoPC6tXjC43k/tJsWle1TjISuD0y7y
/H7s+wMRnM3ZG71f01OLORmgyi41bSBe9JegyUZCmHd9f8H7FuNHZfWMzIWqJDFa
sf0LTjjOsjenePFoKan7VA7LE5UlaD0j0/Fbx/rc0kYN/KAVf/+ErCkNxEBh9ZbC
CHa2dX864nZJ1XyJhMuYDAUB1J/f46m/1jJGsYVm+yUnu9bJPFfpcqxMlnZsIt4W
ZGhHMwcuFj+EjKS7z8yY9SK6NGVAVZhnAw0WvEdU3I0+FYNd44O7JIQ5Kg92O5Qp
4A1LyTP2/0ECWpv5EhqDX5sDMt0Tep+ixAR7DfjccZDostm5YZiw/jT6tS0V3dWU
nKAAcif919PFtTkwKcDdBoXSs42lSHLahOLfDtor6U7ZY8CWUTzQvz8aMuiA9hsY
PpiFN29ZQjbt4bFx7nlbU7n50kfqYXGUM+I4zXQPo9HhzdAdG1D5qOJWP8BYO207
QoO04eb03ODjCFtOqiCiazcaZNiMlZE4U0y/1h+Ww+sJFQL2xX6eQWPOcC8VSx9b
J4u02mlPCKKj1TSo37WsDtzYWo/5dRQgeHgvulmIDXDTGJoPpEu7niEwBWa52wtp
JQfDBv6WMe/qeS3gX3t4SJZdFEzixdnM3rfBbiuXWr41PsMlg4lox0lRlFx5GQIc
OIfawwK/i0ZHnQKEnjMfIjmC9PkRK/s9401/FzXlMKJMhUHUJroDn1xIvwQ1Fs5V
shlGs6IusOgv1iZtVLarq2fCNaDWBXE17PDxU4jvDPjh2TBBOcaJxwBAeX9rfQ5a
BntrGbz9SO93yGuRxYsc5rosBIy3DoNUbdZyP4hL78TtU2I24pe+AJ8OUZE/Z7nN
/mFhM0ghU8qqm4IRQaeIouAGC5FhWjXYYaFa5xkH7/5/isC2cf/tTaY+7Pvwar3w
h8Adqk+RoM50b7ZRODPmy88P0bfRFx+B7NTxONvBzxVr4iNfE5n7pfU0sEySIY5g
naNuPUWdsJv0BeSkAvHLY1o0sYwfhgqEg09W1CHDiTwA/lDJDU27zATcQI/178D0
RMXF/nt5ootIfQzFEUohzwSIVReShZ4UVtapx6bKuNC+0Arwu0UcChVDAVI1bF+b
TJTA3fpKGeBtDJrapvTtSO2UGZNzwFbPlkKsuCLmMbeM2B55lN2sFPd6rn4qQDPR
kYvp5Pe42eRUybYeFXpcd4jqlm3a9Tj+5c0cVgQthrdhaQtgcMz47Vhu1T5gfsjQ
YshtPDFI+SxqX5mlkeWzJOcOXSl9tiN/RETb9pPFj8emP3TFaYPr6gfna5HkAdWP
t4+vwr4ByjdL7NZA5LBY/zfEIz3AwxBHV3//3tO09wPuyCibTdrzf46qMVP8bT7n
oZcTFRPXF6nUkhTiP5QDvuIqeeMs6eB0krgxcEBfViDqJx8KIqq4SVb/X93c6WpH
9ly6DCuPJiuQ2pA5FB8I+PYo/yco1g2cCLcMVKUV1pxZ62/1FOFWwbj9kKyxH+SO
zo7dpTFPkLYp0/iombW9rPb0hyr2lS8iA82ugHCzXtcH1VleAyu1JMLCwe9q8Q8G
3y86G35fhBPhHvxbaxf8L96I5L02H8cTPA5YjsYv/9zKeP15wLfMVwp9FCUG3pLr
srUj5qCBXNaKJ8Jg2/7YWveGVB3rHaQNTyDEfM2RtEU0mqvPGbqYgTzJ79Hazstu
YQKufRRUZGVBjPuPFHStlZEWe6WZKSJ0z2+QTDTe7BcgZpCmqtD2G1FkTMJqBrXh
j0Fw3Yso0hzUkyc/fTq1XHL3P3U3JAlRyxlQA1DwZH/EzMiKsUKyjtql1EhCPuEh
DZPvW7cvv+nKSniPZQPlUXI47r0gaLHqwYZpVu6zx08OY62iMMoSDGaQb6a/HIUA
gwSw2xfXhMy4ewKLLNUXvNlS0okVXOfWx2UgLL+MnQrqiwU7Fd34UrG1C5s6wTRz
ugyI6tVx7Y/GsNhB9kEdXgdIIujdSjxW13JfFdOiLAtRKxcrjiZ+J7XxpKOIWkG+
Ol+V2qqw3XwaqfqZooy0MqCYfZQQYbvRlmEoB9dmzplaqphv1APbjfE4/My/VIpY
2FI3xeK7EuCMmU/dSS49LPQsZg2thOAGjcdFGEZq2xaFVJlDg18+VRada3+oot8d
utZu3M6EVNgdPyMtkRmCVDcrBZIvLJd4g0DeiIqc4VTaHQU3D25GsRdZVhEg2a+c
OhK2Mq9/3zZpnHg20TKX3uGSw/IWGsm3i9b4z3Bt6VNVHCTAvn0akNPVcfITM/7w
+NIYOgk9FxNWKxMryUOxck3cj8gyo+PCMxmfUbHpsbMx4uLMLEjQI1Z12taFQq9h
VeFMdg46iSP415eTbeIfADxKFZI+F6fvR30lv/vSpaQvT6nzUKc525qSVeesRmg3
2iCcMCgmb4xrqkLqWrQ6RzABjFQe//qTAI+zafbMXwcolHWBqWiB6d6gGJ27mijS
XDVXcUaJ6hnVdu3+TvutpXCHySg/HYJl1HSO8a41h89X4o67s3pL8b64svHXZ0sn
Lk+ddVpDtOGN8SKHYSI01cSVkW0NjejCOkhnrC3Kp3BTkRtZ2JyEUUNXnKt++pf0
T/zVgaHVAC4lKovAuS5WDhIc3mX1dpgzomUKfj60BCADI6oqsrPjIbUP0Wm/KnVG
PJnRNfXSjZUDkFJfdcOe3+MmzuCwdVf5V51OBdx4ti0SO1oi9p9aCJy4od60AZ3o
jKZcdXlnGJUh228AYQB/rSRMWInA31Sw9u2zISSD4tCmjkWlvnG72EOdJk8RhciZ
S2w8Ppcrqv/8inLdSM2TiawMCcTGm4WT95GOCEnHDDZ183SbtYdgpufbUSHKhg8g
/5M+t1zllTxmb5E6rwoOKGiRx0kDDB2y1zIyVK53s1cH6C/t17UpCMUKSaj5Ppk/
VNL+dpIgiP0q+CXP0R6lqmD87WABOEeQ7Gf6qg8T7psvocddlkjB8SL6y+18R6gz
MCLfmQRT0malV4gk6KMeMaC6q0pAM+HQIS/BQglQ4/Mdz0JDB6Rg4YZ7V+oCxKrN
O0D1Y/5vk4+9jRZXOpiFKEd1eHunD8ItqxT8yMXXbHua3nQd0jfYIAs0iDFZz/hb
InB91D2isfTYyReFvOYZjGIhpxxHNU8q3C/AlUc4BJePjfmIPx0rIf0TghcnaHt4
T/ezdgEjEpx2vvN8V8tx6SPW0SqLmU9FqJv4bqrxbU+GjH3Kjn7joVUaV+X5ina+
A6xPDRlCvPZ4NuNEvn9ldrqqclj5flrpzgBLKotKvDDnl9IyKl9fmSpCc+24Av2A
SC7M/hnPeXgFmmm10S3aJq7SzoQKWkYvMtDc4wj0oT7zmMWC2i1Hdhkq9iA+TIIY
y8zcuMiT7hLvHkMGzQE3LEpWDZcTDva9iBUmwZ8/nakW4Y2pF6YeNs4L6HUjQ5vS
z1T31YzEc40Mbx37jIwaeNlAuQus6l/V2iilhc38YpE7YCOP6/EgGWE8bEI49lLF
zdO9XHCbvLtSUqbSMPjzPjQ8Du4zDTDLMBQk35hseja1q8dBc08hdp7vVLOmoD8c
6faD1vzLlg7hgAc1t6c0PifmW2AD0mAR0GrS2iZwVSkuQNXuqIGj3SWH42MVVlKl
PEIMboozA27FiYKEnQrllpDx30WS0ko2MkUzr8186/hd2GeujpZWhFG4aMy4BQAN
2tL/z55qL/O3aEe0NR/PjYmoVutfAqFOwDqY6C8Xj8XLL4v2LlBFB8xqgxdKdVxK
GcvYRHjp3gGuxyA0jCBlrwKmX22bgxecD+w2hvtF/aUXc/ypwYdTGTxVOX3OrNOV
fxmaLOndG3bneBrHeop7XzX6OpU1UQgHDJBx+Dtymm6qkbJY370QAkikBZzsBU6g
xMa4c3CQDx3e34tTvD8h1eS/ECL+XfxFVbzwKt6SN+5roFStZfqt1QTE3IMPFsj3
R30BQgB+07hyZ2CDE714vSCLbBtozCv7ZTR/lxQzf7vfcSJV1VmGFjYkEFutMh13
nt4mQ3wCq42iEHII03p0n/ww9uIPkI8fynoPv8/uW6qc1aontmH2+6zztKLLyQ1l
b4DRuuTWiTNc9PzQidqWPsuOKdDqDIJRPsG+z5eNSAJ3gysX1TnrxPFas73Vamss
vloEFhjyyowjJ0ZyOGsRNRMO0/IgaHQXIiYg0+6tgak6mg7RuI4RAYe2IO/ab/YX
cw5QcTgTd/8m1ykVl15pSaSmRjrl2C9tIjRiMDUAQIObIQVCVPLkgelb+0N6u8sH
6Hy6/8W/7B0l7NV28kZvuewmJPHQrGUMMS6nkdoVwTspM5+bzbGyk+AcCgSyQ+T9
NKaDLxFv20GGvaA/jGwM62qQgdzr6Jz8zMqez5RAgXOpWQrcSwzYWYeme20u6nya
2ma60NYZUn0bS9/peYCCHRfZkYWw+OIzAJGsaakV7/DKR9FlvCWl/8loqq4K700g
hWP9eQAdK0Ly5bKOdChMpmq1guqfi/jfLaySwn0SF9CV273ItWrDQ17HWGXkVIx0
fPl1/B4NwsIugk9wCYbqHxUTU4zEESm5kkGycVOMYwRAGS1E1/2+WgWQucVgnw/R
/CjRlrzaPMsxchOEf4kYmB23z8kwkA0V8+E/aqWG5Xynnn3AxkHA0tN2Gcty7A8+
Kq3/O2i1diZesqGcTvGJN7mv0Umv599cNJK+5+8KnKA7GXGb+Lwf8oXvEkpiUMOp
56jo6Uk1W+fK7tdQVjqlrlANtxm/MOIY76Fq2awOQkYIM50VkTdMFfH28wjCrK/d
HCmO6RoPQNs6/+p9jFQMDZl90rAA+d0YUfLQUu+YHnlAT69E6ByUoCcR++QCN4Xa
WfzhvhiLTU98O7vjWKgKNa+pGMB22z3mmxgqxC5K/U+bAPE+HoCnBgLtH+3G2Bh1
tdPRPxcbftKDteYTDoXI8qoP9SPwLgVbfCKq4amljVIsCMRxlzXjcH0+hXnnrpd5
FNZAW+qba2+nMWSvW5zMDwAkbbNq7aq1YQfXPVqbuPXaSEe0T/h9OzLNtsOcdyef
MAB3oF9Nw4QRab9yAVrDfoTh/pjrPGSAltD3puUrEQag76fe2ZH3ltv/gFKWyEPr
57LA4SVVpMNe6UuirJYBcyqQowsFMQHK/pZRTOb/kKI6cNCN1OsaGH3O0ZZTDcx0
yAIrXAm3hV1f4UV/gSsyg/Ubf1buOf/cS7b6SZDnma+p50j2g3fLDT+SBDWwlwic
X2xMoyGk0hz2m60lC3i9/JppG3BbF47Okg8pOxh6d+rswZwZXbQr/bXM5rEKkoBu
lhJvwLU9TsRa5pRbehTlQ7nHVBR+WjrEKpw2puRGAYaBQs+Zz/N2CRKwv1wiRauL
eevp+jYo9r5y228Ntot7W/77U/iXWj77HGTJlckQP5I5FPaWPcc45O2e1Qrhti8G
fq+3HJORMRFiz6ad0w0trz6qqJIdxWRgPccgJ8AYMyQOc5ojn31iZRPRgkbfxKm3
JpQfMijcFEv+Zhafgmc+si2aZBFRm5N6oXdNazxXp9njoZJkY0m4E5ObLfJX0rGc
05D8HoDSkLMWkiQpRnvDW28FTA7Q/UgF08RCjOXbivOzbAfdkCrnEBvW8MK/Mrlq
X7tVHoBHtWuBdtrFRFboat4qK3nboKu9WYcx0bqWKDlvA6A/taRzS75xCI/4SCT+
FuTS24pRVXVYakZKWz1hUuQCMuIr5d3/J219+/d+EuJS+aBv0xwZcVvN38P3z4wf
2GWBFkR3J++k3fMh4K6Ethgekf15eOGyponv5L6WjnQdQx/Vz07SgJZecfzP8j3g
mpLEzbu5d6w/dcX7UrqHoThiIzoNG+scYTY3GQ2v4nPLdzTO3quW4wkmdB6pKvQ0
OW4PFcbEBCHJ6cK0Iihf/E+lnWSd+Esa5ps7CvuUYJOCztIg4n2jMhf3lMOOR1P6
qPB2awU5ZyktQe6UkVrRFW2hjR/miCck/b+PUHNR5HJMOfhtyyX2C07JpCLFZPqZ
02UFggwHBayFtyUgzugJyAaGQSiXzSfSYWaDtAP/0CUcNkXiEy6mmcg4SeFDWJrL
XrOfx7Fc+Z6Cnsk6UkEndSYrMoFeyjwnkvfcM3Fm+vaGSlwOn+qDi+RVPvlLxOc2
AjjqRpyUNZ3lw4SkJZsASpVx7m9bF/QJnO+V5zvjGUUc+WghArgewE2jGPAMD/03
4Mfk2OANt8/SOA7OjOCRrF8WwOmeJ1cK/QFb6GCwOWDdL9z5a5p2MNdGCTNCXgvo
jy5y4nZuZvWUC0Kx5GHyuBMBj8w0yvv+k01dv/yApChNWJHS38BcW01hWTyC7YbT
+bDAjxWb5+ZuvjqHUHdDF9VT01cJdlxXcRrU/EUJOLrH+EtTOaQPEiL30ohS8IIg
6hVzwTlBvjtlEiGsZnpQTBs3TcmPAcPOz3yxQhG4eYRxs3HAANZxvymavfs4qKgA
YRRcgBtpxkcTXOhfI/R6FE5V05UBjw3XBbVLZ6fUOuSV0Llnkx+ghqm4XMC/oX2T
DXf3A/eoVU5kNvn9RY8zS9FryqS5HPIqwlc2iuRKxmXzCjM4ukzHpqHcKWPkpory
dVrbI4tsrpI3edZpEaIkKtu1Hq0fhIBHJd40EL+g/d5WBJO/zgsNDosZCE7FGzlD
e4k/6Y85iTQJBrEWhn/V8pkkN4I2AbFDlMVkcG2TW8DniCICAPkYJqcib8xf0yOF
kOhGbUPbIOyxYq8WGNPdg3gXDsx9YwlQitg1rjv/uTpXdDhUwA1iwuVI/FVNBqme
ZNjcv6QhqKz+4SkTWnJBUGyW7V+YIOzzkAuFlfq60miCZZbcwV23hwKCi8CBTpVN
NzGZbXp3kdqaeDW+VGWHI/YzFH7BwkPmLZe5ti+UrZ8IzNXkaPy5axqQ2ExrNN/p
anibnmhQZNd7EYaI4zXbchH0R61nm0ljg1jLjIqmiaK8NQHUc3crLkGobW6Vom+a
gn8TMQB3oeaqlLrsxPrc29VUN1gHK+esYa6oc+JcOhMY3NgyjZoi6CcGLwmiqVFr
ssGRyPW5MTYtPbNJGdGyBqxa5Bbh94KRKVzwkjcYA4psyHb0d/jr6ZchLQO5VkdV
VfeMPXcAugorT9KxuJ54pSerrmJkCYsuwYGuQQ+zoU5NGb5Gu58LNpgo2jnPj+U0
AeW+YGWgW101/yseNLOPIxjRfcIIcfzKR4UBrmQQe9wI9qRXErwXz4rjnMefAG86
jPg4fjx2fqrTrMGm1uqDJPcgrk8vmLB9e6dm5KgkfSNBGy875uygf8VO4/pXb0In
qefndSw7QkKN2soxBFZ1eEUg9QZk3x6M9K/63eTlQOPBcHLZ3Q3Vgy6Hql7GZWK/
Rhzx5R3i+RvWIkkpLC16CUtJH97Wdw8p393O8kU504ddiFkIbDQRavmY4c90xK3k
u7owcFVgM2a+Xn1ur9O+7ipS7jPvRyjQ5knCzXm/Jp19WNQVsOFOZZZSTcU+PcPt
rUntXfIkMvHsK+30r/d8xv9Xl/MLbEoIUI9hksKQ9YrPxClgdmSwe9AQxXHXYor7
SUkCTnLuQQSYxGf3V9dw074OdHV7Jgl17D4ECl3hKky2dU2EPqcoNSN2FtfIqVGh
lWSKx61v/KSO1OTo0hr/642rQTvm4CB2lB7ArbruW2raDXDJDMUaIYut2tE8aUp9
DBjhtA3jNdxFMxC3oK1K/Z93U8zF+HWiwafy3fijoHbYqx0uTbRcw0DtGqlVQTxP
kJCqAFpgtPnmhAtXDC5p/kr1GrDd9Rqylurz4ahql5t6+AxKNeLZwbx8pTWG0YTy
IqHb6uwTfjpAmax2iBNszWr0wzHok0DB+w1pNmNHy3tvEU6HwQv9j6RNvebH3hqn
O43ohhwHTH48ulgqYm3L5hTY4bhyUYZlGgBq6hgz3prs9WJuqL9QCTSaeJZAWqc2
368Sxj+gqs1AIlTjdwobHIiTz4bNiTzYPSNV8VSpv2pm77UViUZgRRN1uYuGpndM
BfQGAzFOEK9dBWcLUu+s7+l0RfqBMxnLEo0XUXMJLnVQRcBmm45rPZclY/lrvlcP
D1M3JgywerRauaXXg+rRhiCeHhO10IT35pNk/iVIWvpD59vQTI/8MfneWAiclanN
4esj4WTJskpsSldMKUJV7wKLalbJTPvDbIJvx0DyhD0stV0QOZiy+EeRXg1Fvl0q
+skHNq8DQgVG3DmMNqQYLD1AmCXILSVMggYBbFmb0IeVIUGItIlJezwZMvWhwcn2
PjWP7LYtcvG28ZpdnzAmwkO+XCVfA3x9C4U2eg8i4kpTDh0cB2QibKkE0F/qmF2s
n6QRynCXUeOWEi7ZS3AnWKbE3f3z1IUV0ThjfYMoosw0zxqF5I9mRjMYsHXh8P0o
PxFxnAtcbvP/gJLCTpNY+aJFylopALS5INeuv4t/Pf7+wiVDEqZW+cm7sBaGdnJs
fhbYhF5PrwWbLKRzQa9IevmNKrfi2ixg+ctR3/u7K+w2VGqUPmRxKWrFKpQCnAKc
EoIyHjzHnrw1I3B818ITU6gGwyrtKk+ZbM6za0pLiqwkJ0pgnNtKbPn32fF6fl0g
KGpwYB3fPZzzIu5Oe6FU5VuYxgB0aSRfld8nFvF/MEHnjKlOqiqoGFCfMN6HAs//
4IOeQ16RsNGXuBlxa+4Ikke5bwUGLn8fniqVFA94p4OfWExe6iBF1a/yyjfie1bh
rN90TY4V5kGLs8Z2tW7gA3Cqb1Uxr8ZovvqbsMG6dQBWjGse584WYPjJobcpXJVi
Jgm+J3ZYmz7WY4/gFnEB4lBnMEVEbExAEcWveuXspmFUVTDvRuDtkr2wH5K/yi6t
b6hf2dPyvNffxDlhM6ChLhTX1+wQwi+qNSpDfHZGENpfDSBg0WZ8oegBU3PbqwEH
Npby77FrjgLANwoPuFEolqdGz5E9C0ZelSOFPFoYYBRAakNNqP28UmMXFbusVS1Q
/ajpFEaFcRS5U/ZdyyRh9L0ykiUtQD8d9KZVt9hHTw0GTJ9u7U7bD9BOOVqjjETG
7DJYFAGazb4GHKtOMURUJVgnmWQtqvcOJZ+mBlMAsj4Qy0zW3MP+hBOq2Jgv2d4Y
GIdvcmilSNHTraQizTg4HnKl6PhBDz2GMaOxcTwzJDls5BPmDituonq3eLsXyuNj
8f4YaIJpnLZqbUprItpLizW/zb5SPeSVbaMWPDGQtcY0/Fb2OIBZglhgS+mYiJLk
C7o9NYKOZ4H8f9A313PARfxpWGyHqOAO/jef/tLSTvd9rJZe19uDxhYSqXZgMOlK
3yJxqCnonKeu8ohKrs6evRVBc2dNIPmrIW/TOqZ7nS2NrM0llxKPHGbEu6/or+ZT
x6wOJHHHQWBK67ZHOAkrrpzfXit8Wp9/YvaDAXEvbRauN/d8GAWuPaakoNQZh+6T
VlTzusDXeVL/sZjE/hD707tcvjf81ANjex1RyKgMDZewnDyYFfgDQf2xc97dSaYK
Pz/Bubsc+f6KzqqcabM1ooYnXKKqUm9Fc6BypSo/1tUxj15YAzYLHILyk7SHPKNb
7LftxH4jlMGR1/hemjV47xwvnn+gH7nFr0RmGa0/W12S8gWkCrGAQ7zF2kNK/nc6
0SG1P592ptADeHpTZnZFlS6QsU2lrJk4ZPpOVk0J/t0K+BDUPUqk0rTYM0YLTuBq
2e0nRTKdOIxaT9agDmpobvLr/2SFCUpMki1VFJ4OMlfnZ6ZAlvnQzcsmabiQDQeX
HvAo+aHg783YoKsnVFfkTFmUxnJk30jHowsANVag1UBdM9IadJd9XrVe4FvficQ8
nuA3Aj6nqsAQfvszhuFYH4rOUfPkwSRBL/9Y68fzPqx0LIpMNDO8Eui+gVU+/wzb
SVNPPWLXTtmB/gCXyF6JOUOVREn5nhbntdCySrf863rwTAgsUkS5SvpzHRa4Xt25
xJwVe7nPrXPndF8DK80oCiGAVH31BHBw5hHg9opuuWqo0d1FfTECTPgnpuBR0z3M
rrg/Ng7km6Vj6FuLSc9rk/AIW74TFqChv/FFOlvg8fY6vxU/Iq6bOwkg+XKHtH4U
d2l3WwPrNgMeWn+mNXYIxdvD2Vtc9sdn+9ovYIMA+jfpf4brphhVXOSCKJ+FoZi2
IQyoDK9hyBqr1eK2R8ka1++w15OId8GBVwufZYX2fSdTzqLCUFqhqBN4ToNLpJyI
dzDoI/PpZFSh8QqJwqjjdkxlxz3L/X+ZAacC3n6CEFISvGktLoC9cFy4wo8yHtW0
Y0ZvsQD+eXtwucKbsev9CsPYvsCyGp9QsUg6QzNPe2aLObsy4ceZ/cl/OCQz2KXE
bWWzHkSTcUZ99AuIcuFR8N1hgNCt0iCiN2cYBjcJKBSWbIqwuUoQzyZURMwgftP8
UeGRyczNeRKUCdDgyaFiKxkRBPu+xyD2lNdX49SiAQ02W9p0LPV/lQGSzabETcwt
bbsnEWcA3oxOsLYOgmuOyIEipyOE3Vv+8akzTzocAuC6rULumOrX4TlLXsweIa9j
RbF8iELesuHl0EXz5oDXxcBQGwPMurjsnXk9AJPiWtAb2uMn/28pEk1MC+PHcL04
qlyPNUM1iD4cRt6rY38fWXglKqjlXaahU5KkojHV/VXm5m3HAB/xp+MCtwS1qKi3
8YWT3dxeU8Ce0lW4ZSIqcFMdDlnkJj1n1GI71sKU+nv2qhmYyKw7YNy4/Y67PeCc
ZaxMlYB//8Ip2QW1vsqFpwWWnCDJsT/HmiqbOXDzNQKTxRpihXR5nEosYs6ZfQmz
48hP7LlyTBItSTiDLCTRU7UOU8OlXoCknVqTL2Aq7ZLVJ70bWWLfJ7LkpKOLR9cn
vLWGlo8lwfDH0aUfEBSv67e4mDw2ZbdXO8LeptvYe6L5IJwAS7LHBUvM/GIgfao4
8FAKsvMziaKhshLrGatzQIZk/BULcnKvUcrQzXXF8Ie4/rOFAXSk79nWJs33w1BW
YlmrTBDIzmKK/Wj1N9/uymlQgHOcXxj3c7zkqJLdWAgLX8fxCCxYLQA8JblyENzw
DwZQ7Abhug9ch2AFkVn0kZmgyqKAqRu7OhKyxQqaJDE4hRd0A5w4VHnV9cTjOxd4
nVrU9ASNl9hiio7SzpbWsGWFUke97uMeeuiWvVuKQDvZwX/mtHDUSMiQCWu6BK4p
WnGxZZRkJ3J18vuRqK0tDzFWMBq74Fl32OhFt5dRBkfHFbuo+KFLuWwmOf3RFFZa
+RF/z/SUCn7hloRgEAYolO9QHZGD7zUrD+hBkDq5BK0UIEqf3tru8n0JyzD3pc9x
mrfwth0VIQq6y0P+/vTi74F3SwRHpTlTQendAXGXdliQHHzUGo9rchwvIB0CLvTM
BphVUv987PnTvaLVd7qYjRq4sd7Q8cPYOEQ7G5b61WRWU8B6wcz0ZV449PxpLTLb
qP4EdGR7Avdz0/kUDxKl+uggcyh0YPXecm4zd8oFAbm1CeHPm9FwTa8KwQWTWL4t
GwViQj3QcbyoouTcG9JLnGQvlMQQ0Zr8j/krX0W1KlUbbBmBWynbOHViBiTJwlqz
bJLN/77bx7DyUXBOqAoC93xeq9kNpZ/Lu+1xk9ubRVBm5E0WEswAxQugaUx53yDU
V+yEQLEJ1V4CeT1mT9k/mjN3zxnA2WU5WLj5hEteq2NWLMZZG+1DflgnZBIv7Tif
gYBos+F6K5+6cKqKny5GLLu9YVQz5t8oiEBE52sgiB2VMMlfPMsOwBJ70mDOe2Qs
mGKQpZ989HIxRcP6VgUbqaNON5W1SwpDcm1iyQ32y0Lyyvtv5r26RhW7fjPIZlJv
lc4blgjniN0bMn2JkUiQ09lGLPYbvWYxL5ZjmLyGdaWnEplhXaAW1oP8pOtZzMB/
vv4OWoU9upHYODGqbRCM95ViYY9xplR8/DcqLTtLlLw5tG1XIx5bs120ZKKyxCEy
ExRgUd+GHhVT0Dzth9Nwf2SRMRMpMsPbWmtBcY2km9gAUEf6j8KhEpPT/HF3tKUM
BFspY8F3kYkvSc6WffpJYXrnIgI998f2Asd+mc1PY23Khqjakn+s73MvVgvqisOb
MwUhVFINkAxMYqL1KmXLkEWdexDKGaWL3O8skklO/14Q0yJ7QAjCedSDPJPRfB5h
McolsrEsDLLEyFav284KswHEKEEPDb+APoPxPH6bN6h4P0D8yRS4RfkmIgoMVc28
bjrHSkVWZyXs+d8oLAmkQeonWfIyh3V6gilC54oAdtqJb83BmmcAC+6fATAl9uY0
K/DoJukqS3IDX9iCIFn1+FIF1dxMiMwiUuPrBF8zuBbybKu+ucydKHn4FKe1KNGE
mk8Gvd4Eq/D1ffxx+mJRXc+LYUGkxDo17fm8IlBfKtGzn2ZyE3zBFf58e7L/be8+
B/Y5BGhtnaFHFadkVrQ6c572FY7d5H3R5c9Sr3Akq44Zceaw0BRYOWMWhEKGHN7j
rn786hv2Wlt0Oy/kgA0PBmm6aJBRCFhmcCbEjjpSDnTNC3wgSKbQDnf4iN+nUc2h
AlNvdjGU+lAwMp/uZKHIGtKS9vRT48bzsubdvTn04MkpSCDnmjQK4PPg/XO4pmQA
Jfd3RfXlHDq1KEVMWtVB4ObfAJOWvbOnMMjf59pegu1gRJpd/qPdjL0+Z250dsQW
U/resl1exOC3tLVpEfuOkBVVA9sFNgeMLYqRkFXF7uTF8WT67KC7qSf7WNFxQIu5
VpdqTFuvYwqQw1/KqvbXdnuwbQt37dADcGffXhjg2uI+W2n2pbjlUwFGiWjZmNIw
gzfEjTCvcarzGIz5v7O+eqjPYZwP9jwPsC3x89q4oXQ2zECkHRyblz4a6taYc7XP
JfINAoCl19tHxxikuXiZKSOOk4LEKuMeJfcSOMo+Yu13IQgkj24vMxkslaE5xXRu
dNkNvKDNPPTfxUkvAjVCLTq78mujhAm6BIIwsqTgajNbOU1mK66WggZ0l+JdJwnh
aW+TUwzUtr5Y/nfQmf4SjstmMWVJf78d+mPo4WPZvMA7ShV/nmg1HbGjCxZZQEhx
2AKSMCOopKo2sZVkPj6jqzUTc9nO75PX0Ssr3yx9p9HKWtrRn+eCwgtvPVHnIw34
0HRHEJoQ+9OuRPkSL9Ru6jIa5bIbfs9/8u2Nn+zaLLtZK6uouTnsH3kqXVoFb/dN
10sGkLwbnTptH0GqvsDSq3cJTS+ySOEbgxdCEsJD6anCN+EYO6127RzN+JeJ0+6P
kP5DwFFAVqsvSsUsDvFpkVhHSQEnO9tu2EufvwWrl/lWJjk2R0ClkRR1r7/wBXxy
oEToOvvdbENtBm2cihAoMPQWyoUm00/85nR+dtlJngFrNQC4uzZcmpNWry5/zTjQ
/+7wIJi7iBDGDvi79kAUcg0NF1R6vwACWuSdyXKzWemzE11WkCa1GiD+BZ9nZxQF
UnX1+CGPTDsSglVnJVfM1K1vWp048axExKbpJ0n/omt6aUt25zc8T+s7BMWc4hup
6i8T4lf5wl+vBiVRteQIQVoJBF3NX1Eu+1NE08AjYJJHf0gule9YV5US1VAY3SnV
gL0JQ9jpJwuYH2D+Gr5Z7OMEjokQvR24dBLErFr6X85KXh72JIrWEkJiC63Aca4Q
tHCrxogXsrotJwoq3U05m9qHg2Y0eeHUztAubaM/1INenglNe+2FiB2BGqw41yAk
8XGdAA/7d8djTmFXt/ailc85loYCaorC6Xa+4GYGTXCvDNldD7jAzsinz407h+js
SKlGFHE2SQ6OwAOpDvPLyeWvuwqFhXWFhXVPBfgET1cky2IsTkO5UTEeM9A1AzRS
Ztsu6wEBzMq9/klHF5tbHp+G3vfsZ4drO+vTPeu+dg/ebCVKczjf8MJbm3yzZXQ2
C83ENUcNOdWizFBbE9EBey9IsSwJNjjvoasbRWmTCeBdGX9ClfdHWKOXslEJtOUh
n/8f5js8lBYzAufyHJ2C04dSVcinurPjbe+byjBKcd09tvr+TKC951UrVKPdR9pc
ud3MQD+/ItQv1OdBhu9Lf0fRD2/Nq+nGyJ/qOIlrYSUtMfTGrLeNokU3H4AbjlZq
ZO2tGbROmLy6bumNEDZySlHnZovpnV8gxwqszhG8u5W9BTU2WRasFBk8OD1WEXiY
e1Vkig34ajlZJ/fy5tGH+0rcW2Jcy4wCVZ9pJIKOkbFtJrTf8I6RKelL0lKzUBY+
CrWJB2KvhNPJ+06FtO8HyaCovs8yw+IxHOzGQNsdVgQmvBViHjc5vqmzdq1ifUzL
yDawCnS86zYMpJq06v66lwuVdgz7Sb9hv1wD4ebtnCjkYp4FECSK1uaC6mCWme5O
4oiV7EwdkD7gNe030aEwExBWRCZjYUItyk8cetRAocqFNAgRd+qe1b8E+8cnDjh/
38g9Pl7QTLNyb4Jz1VVPzcC1CtGXEHwSG13zDHOFm9QZcaZqEZuoPi/sWG4XxT2H
9M/Kb4M+llU3Sv81W1LCC8pniFUuH3W41/xcPWlnplTByr1u8kasbP8nEOsVVczI
Nmh+3Cs+4Zi5DN+hV3N7JVeBdwn8LyyxkbLnRnUD5a5eHncMZPD/b9jdzGv1YOML
LLBADUF4I7xz1fyByP9RKHMUckpwzGB8Hx6fYdf3h7FLk7nO+xCrLM7twQrkiRG1
xMtbVBMTqHAYCd85gcljOk1oZr3gvKElOxmLq1mVoYPmeO39OaZhfQsLAePlPPlE
0K7H5EFLVO09fm4Wk7P1+JaOxFxIxyYKJzvNZ1+b0ACgwWOf5i5OBL0suH+pGqvf
Jsab0ChzCpD4+a1n0qAdPm3QHx974clWNi9teE2snko/keA8KW1SIlyyCw6rET9y
BYLR269CM8ci9/GA2SHvng7/GfznEl491g+mzwVd/i6d3ZXv/yhT/du3k8wH6dS/
vy36RN1Tu08079cuAd9TUQjrtWmtDrWQSBAAFRX6UCHQmS0i9c/S5Fzteiwzm0En
TaeDu9Hf29BAeaWv4USCDT4aIDw3FUGWGeu1UJO8cvR31NOU/4nVtPZ4QhZyxMdl
Vior3Gmi5WEouL8nFX79qnK5MUWJZf48svvXWOc7y4kh6oXHraSAg5+++K4ajL8z
pcAku6RHsfXcd7PAWC/HyWRKeuyOcb4hiRw6SvrRyjdAEKKirszr7Csujd4THQXI
aP7WbRbH+X6j0GtRZsrmoZPEz4cL7MaWodewkvTDv0QW4dBfHaRJyZEvckIg1ffP
sHhPKZJ1b6QtKiAArwAgIB8xo4PhlGYKNuBrEK3XjGqPz2q2idlVg1UreGey/KiM
9MG8jTv7oIR0h8hWTtoq9Qj0rhO8hmA3u3doOUgQ3w5nvJNFuSbmBf8wBTaE5MJG
aGm6kX+3A3mxgMZz3X5iuNf+xdrXKjZtubH3G/m1z2pwoenua5siRFy5cB68ooHd
P+WN4QaiHWpaZgptMq9flVeJEmabcr2rNK75gcEoU22QPMY9c6nLbwTy/SDgwJ06
xgbkFD/wAgvJoqbru7j3PcqxagNOkMXGSeh41z5IT6C0UikAsoeBdCinEMwE4mdU
KgMG9/wjeeG400JQP6RHug5M/deVE6gHgdCHHTPS1PMHW5dUfkaOrfxll4oVY1Yp
xloz8GXc52LfzAL3qNHyE0G9F7E1HsbQwCMYjzvufXsERSRIE9MsMnEOIqtvJFse
S0N6rXVQQ/bR8T746sPgDjSjEaKSZno+RA6OrKcmoqXG0qkG3cZUYNwEEhHPzDvj
FgiOQE1VFY4WS+9q/ArWRz3Sm98cyoh5nhSZkIaLJ4GYBbzDqgJIjQ737a8FDMKC
xQvDp5C13CM4B3bNMs4tN8EDGf1NghTIGX/DxU14cq74UAbQW9FViapktxCUMLXF
aJMmHn3ioyWpVIDV+tMhGCaUihIJV5SfGFQK0b7dvWozgnAVDxpXAXS7Cmz2k/BM
Ui8jsh5l0/bxoRyyYELPkjHVLCQtZrVim7bdX2UHc+JLletWgiYHpmXSrAf7Zmg+
3we2/4ReDQhZXIAzlZbP+qE/f1JdFLEsqXN6aC1bTO3gfMf0Tti9lRvc7ir3kQte
x4jT7iRZWhfRKaDxdGdHquiBgv3FYa1YcmRnEo7/GwKaajYthx7j8Wd/02uqNAfp
T9OC12gkk9p53FQYRNw74iIOyuoYJejnuX9K7jCouJI0wmfaTeZo5y1A2xZEKNAk
vR6ZCmg7hUI8vMe20O7CqUe8mS8X71+cOhmWrCYjCIaBUiidqx8tUWG82jrkYWSx
LyS5zublgLxr1TKN1gbZwA3pC/jZNMKDzzy2IupRBEIK1ovWSwitxhOpSHLdGAV1
TkEGD4QFasirbn0CgE3FFzLcW1W4AIJPMY+EGwK99WuOeEw0fRo9dtPmwOGxEdvi
w468/Ssit7/IO5ey29ueNB3cPznXLwbLRFk1oVOvUTIpqJgbiFguVn1vxVIGxFkT
Tz1WVjgmEqg/U7FQmv9B1RKXvB3HhwCpykCgAwSMsUSSGfQQK3XgBT5at5OKs8kE
56ZrI8D34+qTc0qmBLeEH4Z/5mEdyuqNrQCAH+0RpkNwSuS+b0Njz5JfSLpbiPen
7HiMsDMlLAN9vFvb0GCHZXQMdijFcou0rFFWeMDeE/tn92mvsHx7+bP0WcFc2mN8
tiLwQtTS8m748BGm4dneIkGeg6e6yI6R+jEvZTKMkJ8rXPgyGBGMDDYfXotX0M14
pVvv1dGPxJ+UsiS2nhuYdVfxPR0CicalyjWLbDI/s27GRDMaMxzw59SbuwXNEfmy
WtAQiC7hMQpX5ZU5NBnevkPQamu9jOQ/DmEZOszLc0rfr1kY0JzMlhUCdTOtWfqN
7g40vSYXhsABFSZQgnp5350esbmlo7rd81BZZRTWZqM62uW5AY3wSgq9tX2UGztf
oYy5tnrl8CUtC/pgMg3xZOyDIRcYP214iWXGCVpD4AaEK1+WFmpLlgvBC/iKxImD
faFSwYj+4OfshlQiqP/zmpIO/WhsHT1V9jC1d9WRpVAKa6y7ZrGeuCcl53jcOO4O
t7pD2DqL47sdt7eeX6BKu+LwbFmNHSCAQP1RMSGTXnBXjGwJff/YXEI/84aMk9x7
C8IAZWa7cEHbMa3A28Fc9L4Z/LlltwL2clcFwHbIbdU3Tj07ihcy0gOZJzE4mBv5
Eb7iu3+CQ0YdXlhRPiaXQQJjdjsqG83B/urU027Hm5xuwI79rksNs8AOTOPTHEa+
wCtlqf2+vqs8HL+SNgaVzH2tQaBSh9UM0i+i+CudAczyb4qlT9Ozjkpq3zWXqE0D
pzMPEcZzijGIwjmDM3K/bh+JJ8FmiOYMVCUSlMTMyxB1EX0hjVaK0/zWdHP4A9gl
Bp1tgI+gaXg7yAa2zIR30fHwDW4+hj1rj2DMMJ8cza5e71HAnQ6SBMK/D1w6cLbb
vE039kwoSDKJAbDciy0OVKyuRmg0MKfcOYyEifssJjWs/UbueyObNTpYFjK3j2TK
RKG0UNbASxsBvCYhauUu9Z4MMlojDkfc6tT6n10ZQcGDl2UTVTddDan3Jlfgktuc
pBeulRI4p2bgulYP6ydazUVXBvYiRePY6WhifzQ88mmacrPCkENqLgdUnAY0GBF7
yO1/i22+6z+W/M5f5l8LVJJjc38QoCMHoOohFmyryjHz350K1hz6M08+XD4GuuB2
YqQYcSreFr9fDr2iZBID2AiqxTE2HIoG2M326ntvYmNfcEVxBQQC36r34ljZKb+F
+vmfwIvcPEv3uElBDZ4yB9e6HTb9ymt0erjo4DQhaiQV3JgTK1aKGuKV0U1YllU+
F38g/pE/WBRuFTYa+itFrrN25UgucGranL0RkIdG/BuRV4IKS/cA8m5vfipOrKhG
WHOpBKbsy9mDeOCMzspMzhJ+pnF1Xmx4lK7REzEC38KD2trQyVLhdROE4ZkZbH7w
r/S1c/RbHdC4F915zFs/bT0qi99sikqzKwB0s7N8Tz21/GgQ1ncwWqvA8npkEVPU
l1Rat+wuXflrg2yY63gOn19l77peBY1hTFN0iEM1qIbjM3d2bw59cfPesJ4X3C09
bQHGF1aQa1sQyJksv0M2U3ObpYNHnn2O7gDeCxD64IbOfwR4fh0tV1Dtn0sDuP/2
tP1Tv9MHMIRnagTbacJweMQioevFYnTvh5D1xMgkNwOWjRDgo0bIG7uYVH1LhZIS
y3yOz5PGkpNq34ysA1x1WRzFklqM8f2oqpOavvkKlUbLrzTN4BctY5/IcbYhfT+T
pieT56RP4e3MgX4pOESdzVNmDd5XjcY8Y6DWRY5uPxtZACIi4Jojv8EQ9lq19IE5
0HrMgm2xV/QADkR+RjqS3p4U/QO/hjjXyhJb/njOm9hUMqCF+rQlGSdfZ/TQEkQh
VAEQYFeUeIg6U8sN+RvmuTIY2mZ8CvEmOcLMIlbPNgdYJdNuuRC+8VnLgDy9WYo2
tEkQTPyQmYruq5OmHsl3DpmBqg+EhAKZleuGe3fza1RvF055daT6fzsRj4nBwj6o
gFO9WBo9O7gJSSXA230uOcNBc32Mp1pkTLddoqEgOUkI/XMhxrIhwkIVnR0hueDt
eaOG6EEFQjubqzMHO2X77P7fHZO7Y/ExdJDQW6MGMMIe4cFu2Sj8gH57uXVpCAbY
6JZeCcbMNWpL4J4Bw8qTu870onM6LM2EEsZEAEUHVqOPbUcPEDdJdxcDLZyNiZ6A
j1zOTdyAb5kZ0ciBwSikjEVtSkR84M0WDGRV8u/4yYzTk6TR2+GrbmeWMZKXFUow
+ftfRGY0IostIkpxjndS3T4ps4h8Dm1BHLrWX9TEuAiNfNcE37e0dnlnGAOupi3u
ro4eh3BVR53qnok7r+FxaZAk42ABDxchB4UI/NWkCHB4k+wrIU/IQTCpZD3hXPvx
W7iQcoBkWr2NXbh4t7JQdoUoxQEkV9lWa8+yA/WtH+2VtGTB4VVY+mU1L2f0xEqP
n2vjhv4hVQfoS6aDlZrzqZgjFRaNXBKG2lHYGd+yPtOw2zLi1tBE/ZFYz27hRKgz
0ObWwwUfyfZjc6cmmU/tM3lVXXyC7nDfdPeUwTwUxsiKPq50gPBKT0X4hUpWxdJ7
jBF+inc4d3U7Xx3KL27zsp58boBM01W7Y+COdvvODrpOOA9LtU06l1qKMmydUDMd
19HBHQ9tNexZHhpvMFzEVmaTOSeUlpUDn8aEBVgudrnhbyMxFMbVvCO7Jhd+J2FV
2SOEaBEy6h4HBFix/ucUALpwzNBRtnNp6ouVXk9DfIfRki/WKp+dISgXOGGe54ZV
I3DCTHLRqFWFPip0CrLAHdrbalEQSGpmhYG4XIumZvR4OLjBc4M49zrX9Gz/to0D
eCxAGLw6eGjeorrKiaqc41eBlKKg0vKEsa+WQf3vvtrowuq4fIMLa/djGHZde6vG
t+4u6udaWjXSmcjSQYMHzbUkuiwkw4tGSAxU9BpjvuOQoyx3oLtoTBbVZOfOq6Iu
3qy2Auq8IHvnq4HOwWsEyprVD9eTxwxNjZnN4WqGB2clYG7VQGpG8j9yoX1U5lTy
bgWiB3GIz8SvJoxMPm68SGuXGnRqiwaLv9m/+hidFZgmTd1RgVqcq50oEV2LNYBw
m9l/Vp6dSPb0vSMHObAoy/TmktF6ezVSIfQnY9uhvdBCvP5fD/F8UZgr3uILJAVp
hOyTvd8uuixStYb2/W0k9zOjDr6tWxUieFiJ4fWFpLxWcVwIyQJjWsIpp8S0ONuw
wNqW2ei2nuQBhbyc+F+94bEDma9rqdlX1osNlXVEUTCK273+98+8HcMeZYeQjf4d
3vU79cE/opjabkJWivaLL7MVu+plluCI4emvfpsDvRyKJZhEKShgL1fwiGvZGQTd
JRPSkgGnRBS+kZkrFurBhXlK9zWblb40K8I0cBf8B8VzbnVdsOMFAfSJrR/MD0NJ
xAh5fZCrd4FvfpLpxF3cNsyKgbLimPkPbeNM40i7QJdixAW7P5N+o0F9scOyzuMk
Iv4+v3M9A6OccU2CCngIf6yCo03yYUvIC51kkHo/7jgwwPAvv9yN7uqwJzAJ4FgJ
QCqOuwYL8OIAm8zReWaejBLi/88f72ghGKj/YEj1BsirZxDsfezTkDSL7wrFaPE6
QvBV80IvgI4XfvvxdPJadJzGz0Nrc9dqodcSe7T8oQvAHHogQTFAm2DAnqEaQf73
g9xA5AjEYoy6L1PFH6W6ASUuCDLzDCZpjdV5yadoOFKa8gn5Xgofs/Vrb7XT67NB
KMTO+KiSxU7OJnlmPrHX3xdr5KUQjt9slBrWAlEMKUPwhTgV2CzwEKakCZGyPdNk
unVU4p8pL8ZXrBVeTkcLzz6aHLPFGjyjvTFvpazhFTbtJ/Uz6Qzv78YYn/lZyYzu
M2nxgU0Y5wL40j1hIa6qHKhDnSxod10ICEbB8ITq0EGL2LR7GDatHixJmYHha949
8HjdkTQ2s6uWzBZIIZrRcdIwUAv7Pb8XrTk3U/nn+nC57Jn3FG0coJBVnAjgyJF8
sSmQ2LJ9D5TrmQjFdFWcbsyMJYri0bBvXmmHR7IK79/CCLNJBfCgKhGRXY1Tyb8p
0Sw1E2kxMgGjWRlx/iJ+YMzNl501jIcf/qZIgAOxyhUueiMOrY/ou/0BTKrYq4QI
he7d2ppT3SEMCWcCBSLVrCdPb/HdoHceiXOsvM4ZaB7jRAStwzjeCh5RAsl1FwHo
QNg1Vxte31EyKzEgNTBNQzDkGdSBTIOrhWgTKYYDyfRFePcNzNVfIjCOTIiLEVvi
LQ+2W3QBA4qoyFAVvnHL1jyC8xGP8yVMBLWTpqkql8Gy0ZmYkhUcf1m5l3XXXPr1
4UTUZ5Vzvu3MpsLN3jaVkBMQIhmBI3MKRdW1jv5hAtnyN99ZUI5E/scIrASixJCB
YHYOf+GzOmJJM3xm3+DdQiGzfuxUDsZb8K4GPMMOUrgePg2Echzq5pLWmCkEGdQF
inNCAjB22AeR3/HZXEcxe0oB5Xc5OfTLwOju/hEJ7MMqPbL1/sC+25tzJJhjNYjV
PnrOT+IA7uBFJEtyHsm4BaAt3dxwSbWhYXOAT2N1ZaAJAsi+iYJyXANaEC9NSPfK
R14MXVmtmQ+DAo6t031octSDb4+j0gUJIcFSmkfE/EP4e82RuVBWNZEeU7PP+2Ex
64GbduyvjT1eRnjKGAYe9+TmLIUVvvazzd34gStW+OtY8jdhf75wBNzfj/LcneUy
Wwm2Z969gv9/vBwSeYnmlAXexK1q2LY1DCK73zBaV81chu5Z91zFasYL2n+3BrVm
BhBY7tMa8Vmj6wvz0lt/4scSP/Cw4GclEYe8o1H/9iYlfmRZMRwfaZi9okCGLid7
uQrHn6KdX/A17fX00n4CaOnl4yeT58gCfSUcei28A5/Kp4gZKlyVL6jS2GGYfpl9
QAN5l5cvF7HhXsoGryj22bELJZ5iT0gL4HEBvqNoTYHpu+OSMcTkyNMP3jh/PiZJ
bw7Z43vsEeBlv5niU1K/K/iw2miHVmrTFkE1Z9mV9RpN8zeriDE2nT4uJts2TZFF
6h8QluoBk9TWZNsyecvHOwFsAy9BB6X9Zl02egjfZqDicSev3xKLWGX7TzI1cl00
s85b+AAaT1+0xnDLARhLdFdpkz2yoBh7yC/7I9flfFI9ygVKUoI0MSrip1zfVJBz
ki8J2MCqGjFUA6QhRuvKTovESyPC6rcfZatZJ/cxU4mFiynjX9x+uUlhQXrEIoip
z2eeQHp2pzco6I/XP1kSaGV/9CpHdEwyPwfpuVLuL6/zMkhGtx2W3O+FTdR8eitG
hiZK45Lb1i2QJBYouqkepsr9DGKJo76b3YkcUiQ+qPlUGmk7wsvds70pleT2KexU
J2JGnP+xm1RIC8IWqiy/dAXHkQohmC/leqtXDDa3pmY9ztW6scwAs0xC11YWxEpu
SW+CvHRJ5YlssgW79GfzF5L++k+KLqmKwwqZtEPyhZgFW3r7uCCs/f1H3JOcv9AO
EII9zkuPK7s57l/cgkyxTPG6RzyIcc9pSnXrSsU2HQlViaqyGk3xIsNLb6zLAIzC
S9H0WOHPj35nSzWzcncs4uJjlVhtbhvYSuDj1r4e71g4t8w5ZrcghDEUJEKOfWqP
Id7HMOaj6RMY6Mg23kecrsPL+urN02m+FDzp3GXvVhIjrAe/FmyH4FXbaRgTE8eK
Z8S9s7AZFdQiMJfpDqRCN8XLxCidnUvew25VPZN67XntIRlqIamQr1AxBXFOoUEi
AHH0vX4yT99s6fq9zHhahJGStghYjg8rzpQ5XSFCx8ex5Q0r5WvYXAll7aCyMZUV
BYsKnI92FW5yi+/KgOk03OwraMmsViMiUz08REVgOolKkjK12cSl8ANF/6oCRH6B
9UMo3RPTGbijQx1+GTwWmQMnZCOCKnpTIDBkCJAvkSab7f75abCbb5LIqDaYAmPL
pb0lpD2tVKNUQnSNsIuZiyuQfu1NP6ftpit1m7MlcLtA502DqPHFEvDv+2hWF6Un
23sr7FnkdAgx5QX8H5XwTfJ1nZ7phBDPHc7m0Gx2An3kfF2J3YdHKp0CDa83qtRH
PZOtD6osjmqr8Y07m51J8wQ7/HM8CaoOk6neCRyEpQupVptJTi7/oNKfqW69MJM7
MhkqVlHSQh4+EkQmmQUgB6aooKqdvBv6lCWvBxQeDgf2FhzzmOcGg/X2g0Ohvb1s
rpXjS5oNPQQClWQ9VjCW6GwdL4jzTPudnt9Sq0j3kNP+8jdQK0EpPAzSjyhMMRit
Mkv6ES6feDTw+KdvHa4crgl/43jz0yFld68Z2pqL94Jx3dTnefHTb4sEPUEhcXBX
IPM6ejKrG4vBQxI9rQF4OUAKveomjPun73InB7oyUva8lXbnqxo8jLPb9FU9gBPD
k83vnaaH4cMI5Tt6wt+Z4kVkBBGWeqd3QDs0a7cYYhECS6PDYstmFg9S5koCQYML
Q25mfLGQJCSCInXiM4D96ikXuI1mRUPg5/DLKPjuAbxZHQJQ9A1DufWASOgVOao5
pR3/vLPK61tXKupqNPQOK8+X/VuGrjHH7AjfAPoPi0CAj+EF59xi59PzhrQMyHkd
6bTylop/MdQ0gz9Eft8m7/uwmAAk2XRQlvZWAq4r7U/0hRPsQw9KVcWZ3WNlwf5V
JzM/N22ZVOOZ7IeHFymv6aCPV28AYVhLqFCT7cFLCaAV9X02uB1g+7HQsT9/HWDw
xQRQnwBpRG3I9drUjk89/IIZ0hAQM85CnRUAGLBhfwHbZbtQgPdk/T0hrCo1eI8y
rUkD8Akgnw31FHsoz1syAUsM98N76v40TGnTJqNf9YKOBhUXky+ffk2IFo4R/jnc
+MS7uN89vddgMTEPat9CQ8AcXr/f4k9bTZwgUU3K5ZHQFO+/c+5ausN0B8AvwREL
8wdj+wNzqtyM3xro5DFBSu5knHs2nYf5TqCa3gNrZns9vwJjdVCR7iHjV4F11hcd
GjCTYptl0Gj3B2gX6+pbPfYdz4DclaT8BPMbSSy4/NN1G7Ee9fWg2oeccpjfJpJA
DfeDkPhCI5Z0JJkBqt9HxkcSIdCZMtExZmZ40LuCbkHYqokkeWB3j3eTJ2fo13q3
Q/MH5LIUqbba0xaj/+sCXU0PGHc697PV0mJKsdA4IV2CPuv1Up05kxl+DZQP/Nho
u1tCB50BLBHhCP4YHx0mb0W35732nKKL6mSuZDOBECx0WWMyw3YN99Va42R6CqW4
sArx5oFJCu836CaioOImO1WqEP8JXsEj0dtkTtRW/jhZamRRrstr3sZ9XA50ZF5Z
dlp5I8udL8UGNvkcyBNiLc1Ci/FlcOfnUNN7rd3tlN78EpxvU12vyEMdO9xSlLx6
mjtndzo5RzIBVzY+TBekcZJEaRJDgz7+FTZTD9/XW7DZjYAk3KzWVvEAHqAjvCwt
mhEC1pLKZrfrdkg1IrhSu1oCYsMt6Ji4axAXDPBuvlEQv4PPn1HcagBzEGwg2VB6
846K/O7rOEXfwjfpuMiSCzRpYj6DsoT2jHm/6GccRIO0QBtvbnYHRDfqmVnziRcX
UEz+AVkNNSGbVdlF6DVzS+5Pv0UABWhgrJDJ30LTo86zlFPGHfGe0tIkiYQ82QSX
gl41mvOr0TiGbo0Rg0UyWGhnpZw4XNTGgKRnWoTFaVlffzdjHTcOAU25XtjQB9cT
8vfvDWTzxzyCYH0ilC4tNqTgwjIKOEXNAuYcNTN96j83wuX37PXn1wo4MdKSbbNS
bQVum/NgwX8zHZ0v5Wua3U9/lJGAyYtjAIEHtssSokmAgnYEMrBsHJ75F1cStrtg
Mv0ZVEQ+7pY1Be0aKMf8DmxJFYkn0bILyF1Q54X15LauWbvErmYIZdZJAGnylbIw
H4d7w2pY+elbW1URHpvLZJ/Ag1XdDHQTZfVWpFl199FWLOLCYoobK4THkIQfBvF1
ZLs538mGzXJr/Q5fPVA3SJiR72BhK7vno3P3V0dZCOuWFSACIGyorzmXjecQmoMT
jsUcrWcEPgMrBp8KAwaXCtZoXVS4r+p2LU3nS+T+dj9zCqeY0hSdVE0OIQsFMbAs
MfJ2m2AkSs+8DeLCSmOLWXoji4d0oLhsN1jAJsIfqY6qu/iVDmiIKV6lgFZNcyxZ
vZQKgThR5Q5WzLKJXZBg831Crt+uq6UyUdaH3w1aHD8Y5koyQyipdu7L7KmARyfO
KvUw8V+bWT3DQg+F6lSx/qIDw1dl0RwLhL0B7Z7qERTR3ryFUa4yyAaPj+woYtQi
yYGTxignoXrVDCjoNmJIaJ1rzxp9UJ5/Yqh/NVyCw9jUthsgtdIhSHyxFfy2kcxK
Oltm9e9RhxPejoJ5odULad9xi9KdjeJd8bQDJyLLBk5sViaZcsStcL+apmN8s4yO
U4msvIWzYAe0RTExMnMazpSWJz3EAPtDMApJKTyZh7tUdVCnUSFcePMd9h/Bnqiu
Vwuha7BLxam9PYoEKDAyCqZ67lVdUxKHIXOf3tbJSeLKZcbpbe4qyArC5Y50bWQT
hqE2PdGE/XoC+rmPg5pRSZ7qBjiBB+yvlZXLtn7xV+CjF2kLmm1FQMREe/jqMAi1
I4Mxhh817XCxA/eMPB/AJKrjJsf3Tx0Ifl5Yy662DmHzrabx38hMiigv6nPDTyOu
9W5oBDyr8GjhSeN1PZ6y8aihBC3aHzFhV64Ti7HJj/JXRBDLXg3Vrgc0gDYL+GKt
O1uuEQ8sXpK7I+7usTuKu0EJIt/NaoA9+Zc1wYnSDL6qj80O+EUL786nja0YljqU
BgqU39Wx3jxT+IV3/coMy1uUjWTEkYdSo623HCkSe0ubnP6Qti4UfelxOFhwTn5k
yYamHfD5VIgkKowCKDtRu2c8bxOqRXiVqqKil+Nz0cXOTnM6xsUg515p0mdtov0/
eFMLm+l80Z6/51PAu8SObWcNoHYKRRL4rvWRlNgNdmePc8f7oQplPdhRto1LiGkV
y7bm6zQ+Mh0vNlRvmZ8PnSBUXuiLO2/4sf/tvTzDxF8ELdGshSwWJlmpUip9HkLx
OWnvd/yf6GKsKT9K0WgCpu3aBfMwJ4qR7mtyJLWIw6MoRJ9wKDke8bnEnpEuPFkq
pF0H2nVW4S2WwMzyN+VW4cmUg3H4E7647+CxHEI5sY/LNROTCCcYx35Dhu46j15Q
FBleI2CDoVc0FlRb+2x2XCBr6V4qjEYPuk5FLsYQjZU456FMI1IwZ2hUGSX0PVUR
68US62pYt6heWHRfvtyks/DyCfOrJOqCzKkg8VXGCJv77MHb7opSoqg4SfEmL6IK
mandumxv+bDKbYlthu9IBVqTZqWN283sfUsGO4tieD4ww2tYSBghiMWazrT9DClC
4s46vNRMuUnaO6kptoGSVBsZ3znOhVrHwEjjh/AWJXs/FdhjXC3gfyukcDZY5rAK
06tpPN2igAmbFX4sC2+SeA7epJ/fW2xAjQ81LZci5AWW/5cZGVpY+KAmtQ3v3o56
99PvJ9hcBamTbb1kdz66f5cnE35SOCcmlFmHwVU5KTMk6QkwGqaZ5xUvwes2gBZO
cG9X5uOadiItxE6knPFaJVcc5DgjxVDt6/xc9URfTh9wNrwl3La9V6rjQY4a0Jtr
F7ZegnJgB90XUckcTescQeyCseyxeE9rEfjwTrK6DaCzlmvdw9iOUs4a6hZB/LSX
alUL53W5zOBDdveJByYpDDtasxQw7cfw3ePPDO+swRIenOoCuybN2jAJhGTvy2cr
NPu3njw5rSCJjaBm0WEa7DM55ZDi7/1+IDJbwLcJFLpEYdmOwVOMvtwWpoukSrNj
Cq5XXQhKDYuIUgyN6OWU9ixgHMPe8fK+8K0x/SpEUWGme7itss00zOWEmewg11eL
8dF6VnGpoz8S/iucdQ6mp4I59T9rVO4HIqk0aZlQMZu1UfH7aKxuvzSogJd2+Wsa
6QQqnGGFlNZbKF86D3y+NNvGBDsf8C3oi6oakkgbGkgRcgBGwTJlE3qEEsJmRaEW
xTp/UZpXFQ3IRrR1hy99V1BlEt+84NKxEUTobD1xe6ORxOLgCtEm/h7m4ROjgjYG
wqCVWb8uOGJfjH1pRWjVRBEtp66vyghaq9jOCfEPNssYOU7dq575BZ5u4b8N2BAl
+ZbsB7q9KEIMqNvaI5MdFNtf7x1PfLlyZnMsWYnP2p0Lynlfp6uQTPFnBu6Bnruf
io9Oc8CAB4zr/xGBLAiuFk1QYFvIFUopLr/gETqAXlgoZd2EZgjj98CvXVOKtR7L
zk9wX7OdeUcKA7oygKLefRWqOcjszmJR5nO4ESO529EJiSRsWu4Wh0eZ2Ra3NJkd
oR/JmhtGQ5qDzGPW7UadMhaKEy91OK/p7OExtaagv9LDnqqvZCsZ5ZrHOFW8ML2Y
ecJzQRcH59EklplDrhk41OY6OuZuBWwssZ+UCBSrHXQfbhWntsLOAlXKm6PEOaLe
kf1o6x1Dbjrq/56B7BHEy2tntgbfnIPwj4kB8TmaSclrNHs1R/Tyk/rmgrRbmBHn
19RKFXpbQ0UXNmNXojpeCWXzb2uNHxnKDdhCKgG6iouy+/0pFIZsmFimZTZKpCrJ
oWNsmjAcoEux4+WTYXjQZ0aK9XwSGcAWKwlivI2YfsPwsaH8LTvb2RG5Psvhfcxf
4knZiRq8ZifhFH5mzXRFaiCvmHTF8NNCAQ9eh6K9m0Qvm7HOB5umtfxZT2D9Bg14
+vNV6AbjHv+/7qKB+ASNoYWwo25gqJWbmaYQ32pecez3lT/g/g5svfgShQC9BR90
Y0vSzy3sY0nRjIuzvj8UeCRF2VCyL/2PTUxhUufzTS/wx1xiNyFsPkLLCD71Wm4u
ad6yMG6wbNpoUQe1TL8U+wYd265+whWcNzk/yTLwuMMshcTIeVCTTBe70PSUD2zV
X+Y3wnzbdLRdpHJ5U+Xe/eiK4utCj4it3Bg3YGA9BH4N79qvB3/0gOX8WwIhBely
x4ccWl8+1U+Br5m7lLHW3bIokX6WbeXC4aRzY0yejQPZlteaazY1nvf7YDIk91f5
FfoNtnmD7lhNRHyS0isqAEx6CFQGOhBgRhFNVAZL5msL+1lxV00fbTvayMwCheub
7ibZqfe6ABJqZUhvtKXZr/31/broK/cW6yCs7b6ukQdv/ejnDtmTc1kJE/gClFlA
jcDpB4ucMsHoGzTSaSF+TlLcJb0TgkAZ6LAgzYvJQDoPJGSqqeePLK4+C9DwNfVN
+E2wShF+dzmXE/4+92SKfKKPTr9YLD5AIYij5JoKI6dUSy8nRRjLEf+GR/3MKcvw
/zSIyxZXK7V23ihFVqpAzHHqYQaDJJtPiG+pujna/HDB/TcmTbVoK6mtJ5HL604T
nyeQ3Eb1OiZv+egGkwZM689FTOC8kJgLbVAUuy/fcUjxej4qc1F5+wpWqF69z1os
ht7ZtEELbyOqWYKa0nd7N3tG2mB1cLaduChHFG3FPVQLs4EoNrLD53ZKXLbkAXRj
M1lch7g/JbJzdef12Vu9N0cdpua+8ahxJAkVzvo3AOYour27vdbdrdnHKKsopCr5
BISg9jx76wNCZi1cXZPguYYouUsxwNwwuB4j2MvGMCVdkD+p9HD5CoqUM6FlDTob
9o74dT4rUm0N/Z2pLBoIkYJLWK/au4zBDXQzdr8qoeIse+yJbiXEy9qeXoPwJUaw
IzwGmcdFr/HrsxyD/aUBn7RihRDdzGKfsmfwaYj/DC4kDJJp02aRYCfUZwb0+oa+
aDFfkqck3Y5e4W+kjANYh8K595O2i5dhQ0Y5bojEwar+6ZYgqH+P32r4tOwn76We
Q3KoJPpmeZDSLKXLHDGKBx4EKZHEUUxoz0J3KXwMCz0ElLk+KDc+Cf27/+jJOhSO
EVWfSyQVsvOgycLW1uFulhyhrCkup/2RTXHZIUl0Zb3q+2IqDPWI41+QBJWQC3TZ
DQbDn+CAGNMVwDIIlyCBCSrayH8kD36rFyr6MkPWW+20qKWuc8byr1fifBf0Vrtn
wHCgplA6ET1DY8dFgHP/sWjBU+bSUJOgU9FiZTHKAeSDL3gdBN/MItG/1HFXGR/f
dQIN47Lz3KRylwla5weJ87fHfMHeJ+ebpr1NfKq9ndtyeWa+sBgg5zMiQdr+Emlb
T96CsACNuuQ1mT6Gkwszy5axQhHWUAIbcVhjrSIzIGfJnqQ8uYbvMMsW6FoHsv7o
aMr6hqtKOdRTBu107vZuttiksLgL9xKlcSBG8DN1b4oFUWaHtcQP2S6kGSX86Iw9
IRppsZ0VtQHYrP+dmHL7bDUSNADk7IfZ9El9XPOObtqR28ozVIfbCvngytevxBu4
FTSnCDlXxiCUmUSqHdP3SKQ49UEXaMjHfPV7IjqWG6U+LHnsa5GvL2+ZrbBrdWE6
bKTYH5EAHsMvS5lc/v7wRarvhZeGYTBRO8nFSWsVZg19/RIEwMZJvTwtjNF8FSXx
dh/8KPS19ClP5x7xpJ7694vKVHcrdUyTf0cKFnxCEhP4LA1dVGWCWsg6f+qpdehm
O5GzOsM4Z3dK0W6c9qEd7LSD9820euS6IlcHkVDwTF5f4haX6HVExbpWQjvUihvw
F7AZQJGsgiRS343AqaURy9PGUF+DDH5FJ66GCPt+T9NEzBYIvwBjv4LV5yFDVUHk
u1P0W7w8ar0tAIrWIC80Rxl73Mmd+91x6hdGSTYcQFMweo39gcaK3LLu09yjejIl
AQo/jLQ1EEVJEkWpVIJTxdVJBvTOSdaSzyE58biM4GUb7SDRcuu93RX7CRXE6RGI
CK2wfvR/qY5wdjB+3QaJhYFjKr16pGPDttZBnEYNB/2+Id+XMqgI1K7Mehczwkvx
p3gPB5DaUGaK0DrzQoTJLv42AHs6aBQWyrn1jSQrZrhfN5NW7CJpXazvDnsl1cmv
oSAdXakMGfSb4B57ou5HnygV3hxpIvhR4658e4kBlBCHe5OX17MvezLXV0qRzZeF
IJTMu0cwSnTIh5vEOgHV716/Ek1B+8Zqzlmw/Ux67Go2spSvhdbPLOV1X9hxxfZK
1rQXBDudOxTvsS8coduP7ffYqLG4xLFEHp+UJEeaX5CKGUdHzLRUPFrZMMJOja33
EO1rZFi1MKmX8m3Dv1EgZH0yIZWR1yCtYXw5S9gNpvIOO+i+tTwBwQMnTVbdpJ5S
3x/KM8W/BdTbC8Ut1TNu8oVZpaqc8/1UtUVFKHtGb2O2KczeneY3vsTRs8wc8nO4
5JUfYypAc3R/lXNT214Y++6QIk1ZQa4gEuniDbJgcnTSFuTFo7xqVS4D5TKN4C35
19iWrdK9jOfJ/k3WTYj7gGKdMGfCL2bNktEzKwTlI30TP3gZUPniBy/ulbbLlIbO
+UKoAc6EIw4CcjmRwx0tdS8/JJL7LveZEThtYd2HqZU+3AXxNU/8PHaHJDkUj5YF
5+O35zRZA8b7Vlaba4gVua7CIxBTRX8bCbvRRC713n6K7eUyOeaMmcdQdxEzXuPw
UlR2LZ9sOEERXvRVnwnuQ+C2mrpLHMGfTQqWqclEKIwS8nxpnNYUerdqj96vVWva
e9z0vs3h/ItjVycHSsnz9vSgDGtBQ0TQagT8AorgRztE5a27d80Et87PR8v6+OGI
wrwHpGqm7jrCtRFmm1/RjiTzXISYCCpARGBOpRjbC1WdXzN5BGLOIl0ELABwhAaY
0NIDctBnloh9iOXLENKxYQy9Xh/5Pjb0Dke/+XYFL9Op9cPQtR4Vez8ZzB4GTH9W
jmyZbBYkRChwxRG8jpT0f08wPQReRYH1z4O1+96EDhCI9drR03E5X/4iFMc1jjrv
qTVwMHqoSSxxYe8OPGlSd9t8pqjkDspO7akt6T/5uZcI655+rJ9pCCXQ8cJW0l/r
sPjmdSKVc4J79rdzUotjn2qq/2mYQ9XTeUaHHDHI/v6LkeD/4TVqAIm6w10ebTLD
VjvYRFMx2QzpxmC09dfNIBV5z/LPcO7VcgnRzef7FlGN2yo6ObXADkVmiZtsyw2+
ldnWeG34A/I+Ebr1qbGZaCv0bt7fxY6+tAsiltl+gfARtct6YkWQ6X0OGZQWW9QY
pQEGKO6rXcN/moeQwpuoqnv1A3hdGxttLxZwwAFlMpibAJF1vs/CBa7To57kUemj
L4MhXyme+ahatiX8GXLcdqUZUrwSr6LwgvVqjcToXr0bhxlvaOOQsQYiu0S2GXzX
vSBwel6Qw3ta8WuCLkmnOFc0c2vdsfDwcSvUUnau9hD10R2ayC8TWNPc0Pa9KWMH
81lIugMRYtWahN7AZkTz3v3novxn/c+zxsdEJ2d3dvW0644TQfbJHR42I+wrYzON
ro75HYxhY3VMbyzdh6k6RA9P9PcZBTg1CvWnS2AuSe92zC+Bc8XOjOqdzcysFm9U
aOAa8HvO7ulDH7P3JkRbZgLwObZWR9m87/jrMj92kuZLGbVuxO7ZW31O0bz+8Aa3
dVPUU4ipNtv7GCRhDuRQznXvA60I5zOC+Lxat8vEgQ1vsCKT92FyIaghNpFyxItW
/ei+U4tBzZqqwEC6EjfnzLMW1Z4tvvDAJtO5FpTddO86UiFnzUXk9a9+4RZ/CxHY
Pygaga8mK7LFIROpZKslm8UyCKE7lM71FdBxkwiLoRitInl3lm2HLEpghEHbkShq
BdurcNJWiK+g2V+Wz7ceIwH4Z+aipdFlgoxLaKeGlTH/cJD2rCzVWc6j/ByBrykp
bs5fiZb5//VtIadD/kOXwbaai0GK1Wwl2Jjljbp38iS9o5u3JHMCb5FC5NX4bppG
VIEBFXXLYx7/9DugQGxmIiBhCm5na+75sQ/6rvkwlCY+CErp8sHMFw94s5v1n1SR
cy2ICGNXuojNUx+hu5xpG0i9PKL+rfQBaib1mjYDfwLgUOL9Xg1ayHZbgvUZvANu
pX3gop5ObFbcxeyeBLnP5CjoINNMjGB3fu3yZKs7d1mb0nrpN4Nopg4G0iakfQUu
lWU9yl42L0egqGPKJDL1/WXkl88MfCVLlxMMkameoMrTYrpFyf4MRN3ECjjxiAa9
uZ3aq9CdokcL7+1/W3kRq8UL4uzMdolEQEF1F9hzbSggmUQ0eyu3B7z0inSDn2fI
Su/8YNAQQ2g/pPMVxEWXSJAtbmOAclNKNXKAlXXPhmctulkx5KRG/uVK2qUy0XhD
8Iakw9SYY3l+UfPbKOEV36vhTyjcHz/DD4PlpMMy2A46xXEWgmF4MF3aYbKWQcfl
Gvi/NocmHiP9l3COgkoS/6NZ3oEDmz1K1eOOPyJ85JNF+I8KhQXPs7QjaJl3UaW3
V0VdcI5xEaq1ewvCQYCNFoOAgG5yRewe7weMXrUVjig/nc6GGdIrGJN6OfeULEFz
nQXSvjAQtLIJQart28tAgZLf0f29DclJUM8OVt/iST7PPtTG0psPB9vB3lTIN9dl
Q0lri4s7vK+hHplSJ7vf+VQ2t84hsQprYw7MtBf1x/Qpdi+BcCnk6DB38hSLwdqp
mHiVtC+DBQHkx/3RccvakLfgUOzwaNZc9opk+tIoq6eMhyHFAd6hZYQ0WhynnJmB
OsDf1MYzryedUmQIhvfbZ2Mg4hIieDewb1JuEifR3gzp5qAUTj7S29oCd6/50ypk
WfL8uI5u2MebvlDOD2E625PL/TiK5MN7EMjOCEzv7X5OjspbK9pvIlnBuBB1LAUh
7sqmxuUkMoiFshxKTE0zaui8wPz+IL7S1TPVEdaiC/MZR6Mqm+vUqbXury14+8GS
Tc42WxBBiL6bhX8qw5drxwgPjWES5ASZksIPRlKFRtrGCvAO6/+LlyTOMF890d8f
+8A53CNROY1MEUNsxiX8WqJNEZCZku1tnKKh/X2EnnsA66SbEjTXeGfXQd5ufKuW
wkjlMXrLWtduCsvAe+wWuLr7faio8X1Jo8Dz6aURHJh/aCzSkR0NV0+MODHQZoX3
re4eC8ckhQmia06PKlitd+2w+8JsIKx2cifR1LsPZc+6AaQyJY9ZZ9S5DRz1SKxu
bQS2r/axxx5a/p6Pg4gRpZ2SHWHbymxxty9/73k8V4OSxHmPDWRQFjZrENfwZke/
qikW7GRAUMd4B4mxVxddNmDMphhf0bFOjrrD5k3d22c8QKw1nhXn+HJFdv4P9jtB
fxVuLotmIi9uy95FT8mJMGHlzDaw+PgFFXklt83qXc/CV5+CRx2CChgluXFrOidA
0e5vHpm+uV+a+Wits2rZUi+EOyZeYXLwhg8njwwZr7aVUp2+TIZzRVx8xp8t1w/O
zwbCQ/kXY4CnNRmL6qu2HP7dqDhHR8xv9skW6RlmJTiZLDNRddGGxbGZwnS9HwyQ
6VViDOspTdvwN6SxDFw4/fyoQXXn0vBEBRnohIz5slmSWfezwh6RJnOXmhf136Hc
faIRMn+01MZzxDGNCxRhT87V/ZFrLaK0iDZSLDH69JEdhcka7Vt7ka53K4mXMOp+
Lr8rQjeH/QhYwc8s30wZlzVglretBRHO5wHyN5+y5xkdNLroNGT60ikYC4Z+fXMA
7CnHw2mBNgU56++28yGUH8YARx414qf9jgXHjdflgM/IrrPl7wlDYgOmVcaRce3W
w4OGrsVbxIL0Yr6A8cI+wNAlqWHOtWgbKA6TrV3vPg6ZoFqvv6joNqohS44MwuQ5
uhgxkF5jmHsF8odxPu5JDsdF77JCQIJifOXcsoXNxM72Z+8rIA1ieF7TOQrZSiuZ
jSmzZR11myDR6aQSSOzVZoxNyRzkPP0Nv93Yi6Czq8zxx5GK2/npIISzBLagmv0e
91Xv9MlbqYG0K5g4E+SwsdaZwzFkQ+BZ0YjTRpt661K/LgX4FWKm6wqt9KpJegfQ
x/Ih7b3CdCCmsXYwnoNa1KvZ2W7kfJCvIIRU2xKWRLGza7DoaEqrF+KRF1U3pwZv
inCxLGl/Ibl/YuY7ID3bILsPKtdrlVR2ANRfN16Rbzm48MpNlc6JERnlaCA8fRSI
ce60XuyxQcW0alCq7CLocxJGPF1KO2TZZBYiOMw9IL9iqmyl6h6dWDZC62vqiYgE
xUUiPifZSc/28MUN61vPgtYiupwc8nI7T67hdDNSeoBbtuKlahZOh7jhLLC9MD6P
kN7vqM3VubqTwP581kvxMezaKUfo4RA5IsmfTMfqFht9hsDX6eSJb3H4Cgwui4VA
zXhKUeAIdKOMu49rHet9McVG/0MprczfsCYYnx9tdJDa+ZpN20/o2H6uIT9VG624
A+hS9wB0ZDmGL9Cb8pE4Eph+aTm4MCO1dmrCJcF9dpxZM198ZOqFGKz3hcElrcua
AFNNMOo5r0512jJWAJHVXMVx+G6m2ORtawhzcDYGDUy6g5JqGmTzHO6gjm2StF25
9ubpef+jId7z6XDIX1597V105jnDfDBFH1xHD5RqJABC/fpXBHzFVQ0ip+01DsOH
k8aMZ6DhoHf+UV+2qAo6GP10ABMVSMlRcJIZALorSIjiRD5oCLcgesuwYGXyEzK5
HyndOgs+tFh7gYvEsI95LcHY4Uranv+NovJhod2CEi5ziWhivz2Qki0Y7O4AlvVB
GSVNQ+AY1knCdkH3ZcJ1MqsPPeONtG4FYH97bCeloJNDUiX+BHC8r+/sZvuQmuyx
+QGZLP+EhUHWM9pb8MsjA+bzIMKpINgZate3XX1y18ZJ7gXJBjTS53v2Z4KUaZbK
IvB8rhmLJgiVHYDGy27iYsEU0ZPBoq/0T2vaOQTv8VmBbXlYr31urY1m+7y6wmHg
RH9fJNh7MfUz3rkySwjsxp0piAcgk7l9FbvNwR4jaxh7LO1QuNGp+nFxkOUcnkEe
H3NaESspMtr77D6mCQe8Cxqe8VBJju0dxm93BsLKk5awZmtjoOUFowtkX8FuhOwS
8TqE3Szht2jg92v1CsoIilby1axQB8roxC+w5iV/RMCfDFGnfNNUlPw4jK8lGed3
TIlLP+Lq5nzdh+VZ4mx2lIVCmD6moegNQbEQWsHLX4/aVIPPNQOI5HYu91znf5Cb
NLy3zOAV1CM857Lr7BsUW+rh7qEci6jMl+po5tx3ceYlFRvOitHqf1VUVYr0fIEB
05cCrwnHNesE20kTegqRM9j/c8S7h7CeY/9eqEfScan0MJ3NlQ9jbKCiBNrDgDgx
myhpiaH4OzuvNBEU30XqNTV301NhRCqpTHCnCyeO8epj8COQhKpTM7tMsPcKfnqA
AFbpRuobSzYBPQsAf9SpZSl3dx4clKXG0XNHntlE+IqefWtXSBvx2ZD3N65wVXFY
cpA1H1hFAwWBb9KFtKHOFFvZ2yKwuAbl0yY4oxFuDswqIr+lDwFROeUtCxwr0wxE
xpSdX3SbYIQVWIzNYWa/9tUSlPQ3ZHKqmOAtaB7ruJdQDM3Z8RwbI1ATJnHHRFyH
KGnusxZfbBFEneW10zikLtf4j+FiPWCkuQmenAY+/nXyxAZSCchnuSC8KaG+caIx
IWT9Cj9OmP4kaVjjU9dWfMvwqmoSvAiahb0JeS+dP7SZIeISXEvQGeStxy9bqztC
yuBmwiwXod76VU3TeL7GV+jO/msdLWH+z1J290NALTQUuYaqgk9ZMbxexokwQbKi
BAtbSC+9sekTye1aV0ipycCJIHmtGwkaewUFkaAZKwNq+TnjKaGlvEoNWKrakXd1
doy4AlAJGJCNREiXDcuRoHRn/N1Lel/7OB9lEx5aiQIwejGRzZNPqCOerDNfpm3q
xJVlGCCR5WudzVmiRlCUiSRf/h5+dm/EzsOqVVb43tccKR+cJ8UWWmtPJxx7OR9a
LcNmKRLtT5khrJsCpiVxGHqJM/YgSzrFKtMSAYMel9Bb2NctcvJzRb/n3m9cH3qw
Zyv/EqchoXH6Go28+gEPJWjNJdbBtdUrYdRYjoQhO9SN9EMbAImkbo7H7atLdB5O
9He+duKILZaT+jpZE1PNFgHqQXGLLjbuv8GgJdJaUHRmcwSSR2fKLjEM0/LV4Cjl
LazluKac2eLM8dfao+QZhKgEl8kb0PY6mB+2c+LN9TtzbNg93LB8xRBO+/QHeX9p
KRPlBFtGSirdwMoc8GSU+2CvDcgObo9dTkRAGNeosnxz9LuhBgF7d1/JZwE9+fl6
pbz4NHa7mIfEGFlYULT5iE8Fgfs27dyO2A4S9HjNryuwJbhC6X21dD+cMQ0WGtOC
UloQDfL/4dVte2sm8Bb7osFDx5/4XSjj6mu1ylJ6hknrfcPEJAgvBtVyyqjv6C88
42uBICJ2z6GoKCiOUDjcAcWCq/UZTU542lsGyfwD6p855VASDEnp+y/FLG/0Dzcu
2K3lNR8RbT00YQkbN/ZP55r5oZ1Pys9juafC2lafVx+4MomqGN/YfZ3HSmdY+NhE
Pg3FMYF/5JqwYnEWI9DZ1T60n97kBoRRrHpEvuajgZnyD8E3W8DYvCfVyjjVMHc8
z3ji84Psz9F/65tL60cwb1sDiS2sBV3ppjrOIsLuP7disUTBTeUGv1S0AtoIbF/5
pghLYWohCCp6fy8SwJltFQ2ie5xpEkIBQd5owird6oWQHrWgCeN81b6DS2Li+x3+
fwA5ty8PJktWsyfz/gSmQylJ6X0kVVgfF6EAUctcgCcY9QmiK8B0vmidr2RgaK91
/sJB0eNCLiMd9jvCi2KBmrZ4+hRtjenwzmSeeEW/ujOkNmYFkFHd8tJXyS7iyrA6
nFBgZTFRoVwHBlj9lZcpxl1XCybv0MkABrB30HvOl7zwAZ7Va+uuoBofBO6430dC
mpXjWdMqxKgY6LQ32Caf9zHUXlSmrS5BK/HPJl/hX9rceV33Vf9mK4Ra9fQ3sxOQ
VKPbxYzT44iVT08R2xtNgmsPLBUlJI26jwV0ZRivi4GlTa5YB1sRIxlJKgoniwTM
wB4J9bOievGliobXQdp6cnyb2+sN/Dxmj9fDn5fATEzsmPzqNi7Ty0+gkm4BWZQ7
hQpVBM/0I4bTmexa92/iDsr6AnAufjea6EpmJoIz6KidZWqGH6byaSnJfTqaL58i
7veszlDNW/0jd0pVkShtXAr31FGNcWqJFa+xKdq0otaHE4HqVxSkZbRMkT9noq6x
WZ91N7yKcVWOU3E0sTN25GJ04wvXDqKLJYke8N9m+bB3ngoZuPMO3RhT2n91n+Ep
b8GMZpooa9a/0i1zUlWOc1bqaVvcnrUaZoP/P/gpVR0TVunA+eLfRVYApjhs9LzP
Gb3Y37nDT/rZgXZ3LoMqZ/xZe5GfddNGUpxCGqxyRa2/bSSrTXa6ggXm9clTf9BD
q0ayLjOpvmjXmaSr47nBJDy7G/jEN+SrgU+YN7Af2jQJ1Zv0b9wi+4eZJCTEVWaf
KJ8Vs1puqk7v+QfJyhUhNB/r6fnWdVlohrYj/saF0RcU97r5k7kStdBA2jH9ARzB
ec2svfHW5vbd+uJRaKUeixqab8tkW0fAyo4g8EM7YmQ0VXo7JhJN/UJpRp3a0GNW
vHTneLx7GeS1rnKdk54jcT9C67W7BO6/Gj9j996BCRw6pf7m+BGZn9mnwU50Ebze
4/m4+5KaS367oESgxFNoKYrp0ggT7Arebwcs2MoWDk86UUmwjJz3bAv/vandcLT9
6R5kgIiFL9f34OC7IotH/kezzMOjjJdI2dtpAzK0YjCBDaoSnvaPRQplqMSYzN0T
tgVyktAfLGV4K5HSXKyxSZD8zvXcjq+KFBmbp1SyxkkBfM1AehoLaZTQ7R8rm0Zl
m4PTBmzAPiDCc1LgOENIV0uDSy7NoqX32XnTaogjn7FUtbw9QJxxw8rD+Yu9/4k+
bac0ptvYJrqj1f3Ivj60+RwJWL7/okOmbpunycQKkodkv0KHEtMiaGzQqqNpYqgI
Deis45HxRKDA4M0wXTkO9UgkW+xyqdDfahmAAb2V+lUQI3rR/nNFGfKcO/8KgYIr
6+rdxOuWMYjzaumOs3PffcsUtCuUvp5OpZzqn09OXYneSFuv9GbkGgRBTNj2CQCR
nMt3mB+F+atqcpcOt8JaaJV1WwpxQJ9pv10R0RML51GhfrXiuYtIvT4lCMtV0YBO
PsUXM+Ux4bOzpeRl6A9SOo/XoUFXv1l/g4vr1915dR4iVQ1ZxyP9GC30z4p0XArj
EbyT3hxlEJVjwl+6XvOu75LEmxOn+PXmBgZuUTROwCqYUmlDJ5P1oShktUrPzrfG
sCkjVANIUVgmkIflnU/ynBF7wVGwGkjWEXMKFKanPfOrbQrB5cUsmgNf1K9Fg9h1
m3b1tWfTRQ5ri5pmsYo90RFci7i+h6lOJw1QqUApQ0yoAZ9HsHWF6NAugw1g/qxw
rimBLTmiBEBbZC5hzN5wt+mmjmhXADHXWLT0kwp/v4I/9wJbEEv8azzMkByJdmcg
RFsHC9XHKA16iDVNsx74rDrueJo3WBdXmlQrf/MizbFDt8IRKFCZE4Bp2vtsjUC5
qIquzUSfMUZm8a8K61HrfFR0tHVLAYB7gMAh9Iqj5kcxidL8Dd329UQnQD42XFqE
KzxiuxxHYAm0gssD6UucdVex3G29ml6XAOKgFm7ljNnVP4TVczmuk6XTzUPcaG3z
uWljgHpx9dbWtP//BMkFTwt1EFJtNtZRilBY1lFxlikJ+M31n+nzR8E8FLDIQrZX
C+hnKDmY1JL8Nw9ouUoHQKtYPHcyOC7LKDNQsQ2xWmjv3TDJjGzHowyMV+Wb4Eq1
BVHyAlM9txUHuP3LVfxXUmP6OLX012ztgi0OudnurEGOcSckJx1Vd6iXGwADQeu9
V7qHU4a3OEVQg9aMW0LRrwxGFdAvaNSIijYR268hukOHTCIcHhkM1DCX9qSk2Uty
l9tX2Hiikxu1ycIiIbc91WlfQWOnIwljXl35xHcLmGqFKVjQJjvXQQv6RgvDM7MJ
9CxuvpxZ68qbYqkoKJv4SYvK35kr+mC3Yx/rINAFpRcdpVhf+urmLSRZlizzAA3R
xJaghCN5ycmQ/xuoKf5KmZ/CJ6jZk2ENsKdSqQPCstvoLcAxwjI0lzeS0miSr5SG
hYCE/xUq9zEico6MF+KlscNbV4Cquj57K1FbVu8+/slVNoItCZQdZO+b8w+ccAZf
TqTSds//c9nhbKQEWkvNGkfspAodqk1dkLaHjHtIGZvsSWNISIl4piT6KK6utZbN
JvTecBYtXT2GeEi/SSf52mQ1trOw+ycVsQCazyKptnJvJW+1Cz/mgn1kiWd6T37v
yjlTP/UyIfckWMnNQg/POa8hvKgGhYJos0//8jGjaEG6iCn04gsRmqDtc3Smcbta
iaUZ/SLLrn36Ie1qJK9luLr81Oy31vnhJYRyCpzz1CqaNE3Uo6nJBoVOYZQVYvPp
OducUs7XfK3pFnADJI4u61gioxa89qTw7F36BFdstQgs8Lu6HBHVUehlKTNrMlPX
GAFA5LQiEqJDB1nejHFFqdR3S34AhmvHpHXr6zc9uNqFkLUz6+E+fzcZ14Sw044Y
IIGO+KVVcEMpgbAbymhAPx2A2N6XiwXJ3Tnh+ZzJafju31xhUweYwQ732Tp48FAu
pu7UTMSQr1dlRYIfoX2nyXeMXHLp3Dtbu36hdf39paY4n4HTSuwtPU129pUivtPj
Q4nU8qCn7XjeJ9js3qCFI+MVWHCGUSf2jFY6M0fOlUPWt3xYdPWpf3Zj7SOcyfNY
XBfhk+X+xcjjxaQH6dJIqfbOjzFvQ9/Qz5cNbjv4EjQTAwc2hvleWDMh94LS81eP
cnsH/oXcu2l4TrdeUlpktBB8aM+vNd32lYQ847dFKURKyv3za11yjLTT7Hk+ERQb
A6PTMWnObfy0ShBfiyeqWE1J/sVZE9K04E1MBXrOT5QmyWTNmcCehRD3ygQoX3T7
xb5KR2rUMqtCwyc9z3USFdcyAOqud+c/irS3SrVPWX/9kIgga+y9oiA0DgIDqCp3
hAUDEMwh1qZEn3sOtFHTbnv5wFa5ZA9bjbmxcyprwYTsHCBX/565BFv9x/twAPpT
vUJjfueDUvkZheQzLn3i+Le0fsHR74jtGZcveGa8hfEPsf3mk8z/JhFYYNg9hCXj
kUgitcRrN5ewvhMmZMbhQ46wuzYTZXzRT4Gz9is4pyaE91OUuBhP5SDcoLoJXtWs
8X2gmMV8YTLI/M9r7Sw8CGkTP0GtL5nXFXtz/nYK7DqNWcV9V37fN/yNng9jmU4o
yFJlS9HMUB8vO00ErwNvpfhoZt7N8GWsu4HTnmaP12W9aRMncT+dhqC0PfupsDVj
28bjGL7cUu5nfbXM4uiD6ghZRVuMchS8r08gNwRmJtBDbWEcRM8uFcRzNg7j6tKc
iso63D0MBP962XBrJe7mNLXZN29rfw8m6bGXqNVHHjGCGcUrk0c/AURjdo7KLzQv
A3tv6RudfA8pWi2bjqMVIoUw+IJOE074lhycennr1UBV9KDOyEgVVAJXSkNPQ7Ic
Fb1ZK0sXEhJoWuQUmBpWOxcGAkb0LeitBUPTFvXrgPuNeP3JFDgYVr1+niruHMuo
0SQvWFWuwNB6YZn9KXQfeto5EohOwB1PKWUQoVSEIP7T3grc/WCwfffuXbhYuKxr
Xn9xw47gHGlZGofIvDen9QgaZBTrtAMJ5iWbxvlEmMGaE12W4522qJpYSyrlLq85
mzw7kkOVs56SJwfg2F3h5l8pzuOea3AjIQ+aGjyabQSWHFutlcH5IUJy5xn6ftdG
+dvznncal6xdIBUPlMuiB0L+MmS0TtcKIikVmJDXYkyLztmqHXivXW3iYokgzRYZ
1j0LTBDeigS1gqMT7fQxPkqnkzGBCnnO41bxS0L2Z8BCCxDWsBmWKY9WaILVimEp
etVvTTXq/0VjNPOqP/y1lZ8oLvPm+NcPXTFzrpwmsi0Xh2r7uiPglsY818Fda4Z9
ImtdrZX8ZA0SkLR/SMTkbVP1bDtUAB3Mv5ScVfpmr7Jhw/0MN11NIMac5tGa35Jd
M0/wviXNyNe+r0E8AIHIq0HH31K+sqOEIPJf1ag/HWAGjwTIF7802ITJoJdnpirk
tP854jXg8LQ9ONzZbuqnJ/PCvUd89gTumxZJJaSrWaVGFzvSOGhMEzaGsmm9WgW7
Iiw1R9fN2AjdxC8axtF3M9EEexBvHbUk/WjONCKVe7ANjOpajSMzkw0U0Ak9609q
bMrEhNmcewuZTl4Q+/Ew3Wf+31JYZoaFiXAgyKUlu6WMfmAfRMSYTz17qGQT9/gM
Ekk3/RYfGWqErGeLqZYUszziN1fMReaMuFyQIGssD01GlDxd5hhw1AC/lomDckXB
Gs1gHltRtjoumt1gqB2UDnUkoa8CppVVdY+J48f+wQXTsAWe3mEc+QRvkjSzwgNL
2IBBYkt/+cZ240pFlTc9Ftp9k3sgxsSWtt568YaVBVBCMMWygf1ihklp2kZV4qOe
S/w5TheKMM4gfp420KE0Vnm8wvKZSKFvnd/h7MkRyaksMwUn/zJpZjZZjxBS6jYa
UGw3ozqN5oFO+WlZuIhqMomJy3Z4EPmomPTyecj3IOpDhhrG+H7NNFB6Fo5NojK9
FlzkAVhEYZWzg+WQNeNYtvruMyLsZmPYn6ykxmz5VWwqZ5kE6plSDRiCsyVJEuyi
X6QERAP3Key9YEYp6jMxC1KcWkCN5gTPqMslT5jTkOPuTgB4J8YKjfD8fM/u6XNm
Nz443ysWKaIi1Jb178Hc5nJmnTEURmvl8Fvwl5+EgT3aG0ackrpPuHmz6tewohNa
A1FY/MYLJWM9+5SHrr3tjYNmIQh1lt6ERv/nSLpDH6OuoWY+zafIUlIzJZVdvFZ8
xxRBrjPieuRYew35QvqbvVZVYTEVula6rnoxmevl3lRRbnjxdcsp1Z4i5qxDXoyq
muqbzOqhJpz0YbK8GxrzhgGBqXaWlVQqkAc0I3vZmeBxbwX1n9itJWwg0bpjk9mO
81DlxGn3dZqx1KpS+pxdWYy5pnKvKqTQKaafyX1N0IOM2mUwzkxV8ZEqiXttQ4wc
xHqN7ii/3p8gHtarkhLnylxouBsEtK7JRmrl2C/d3g5mLG0thAc2er8foxpyGut7
mJCjQfjWwbZlYpP5NFCAGSgFrIVDEUMpaqm+3KRcPz2bzXiDkcLHeon8b+aqEyC+
BeE+opsFSdU8jot/ehQR4x+fnHYdgSDw81vG4wZF/n4xGhRYzRpvRMas9dwJWdvh
s3oVQsUxF0cYS05Pp88upFAnPlo/jb/Y/39nIwCVe9XgZ6G6D79WgKTtHE3ziCA5
p9pkiVwBM0M+0NX+t6UuA4ndciEVj08mQueA1W7ET2fRO6LJjYDuJYbHPnUWANhW
CzQJSciEn3Cw5dP9BCWMyrawYhKv27yV30OtiHnieBvkeaWXEfBeEJfTa173CuMo
OZa9/nDmgZaZL4KevGM5LLar+N5AoxoICeHvnTboNiQsd3u3SHPXVwb+t0jjXyhK
jtij4lnlA8vmzTuwG2YqQPOKzcYpD9GgTv2MnH4o317iJ6OUvlJ+EEYSXzprv5n7
vR3hxf4fk5qItGbye5uJrq9h528WtQ/xeHFFFQbkC8TtBTNTVT6KQ+t/jxfVXtRv
pt6dIpsAmldsx0vDwYQ+aA12xPn5MgQCxmCKO9kKCguoJCOKFt5/T6+Hg59n3K6r
i7Riuc2W1VP+non3aR+kWhldlMD/+ocAtvIqUC4gnnpnqLYHpzGhAspJHnPpIH8C
FwDlFe9AJrZGI92VHdEHcsTlGhI4bZBD13BSpJt+FCoRqspahr4qvKu816ztwqr+
LwXoRwEdRtBogymdO1iOBAkszaM+DvWbqieLSSzQBW/lRgpnNwykmstTazVueMXm
vJZkJx8+2apINIB5vqmuIe9K/A6K/memCmny9lsmZKtUPIYCdXiSbDP/BV2bF/9q
Inw+BaMR46rcKnpVFMZrCaIRHb9H4RL5TAf6jvuXf2VAbFu0ygLbsbqQUGcF9wcu
hrHDTdTOJdkXwJP8YnSyHQHP/Qumu93ujjQ3OaF5PVYMDzgheRDIldDdam/QN1lL
XeeqwgyMmGaJF+QVKP7qR6M37n5ykXbSzg9B+jPKLK3AmiPhIA3Nd/zRgglgw6bV
ZVJWOj+SW5xJ0oSUeQNa1SVhsXi6AgHxE0n1uyWDe/sPt3YUXiJVJkRKFk4JTlNR
nfK/TpuVDH1pY9XqDDgpqngQ9gTdUFdrIElA1oBeLWKqdcdAzjsBOL7S9UegeMC2
aL96Y0dBSOW+KwWEMkQATY1YszQCsaDHL+TZ+VkUI6/bvBWa3d7qv1rFKntFtScz
r4255B8s/IH2ItU9cU5U48NUHripOK2Tc/uQNMKb6M0joTyDXjWJ4qBk0pTdbGOf
H4WkpgQJ0aE/ckNki+b+a5fXQgo+DeDn9D7eAxF8ORlD22BlMxt3NU1L3nvoFjhT
C/nSACz8ucaHS1HOwRuIh0ABb988f+jNLhkeJJcW3dUm7X1XGo99UlBQVh8kftGh
9hIt7GUou8cDgZ6JB3mYstYhMQmXcXxa9IC5UMrZR3oCOvhCFnp71cnW4uPWQuJw
83Yk1WvnCYmr+ADwis7B6Ud6EFmqPM6PaojgBg+Nh8GgMc1q5HtYYyEbO5Ognfgm
iqhJ+zP91EEJJ5HSLY7roQBtCGmedgTarKCOY67aqzR6QbRaSZSP2vhVXDBbmHWG
XPp2xsk0aenWFXfOTDKDC7/arVTC7RuSeezsTxnexxEJMSksfVMffW1+kNftJTeW
jJOL+ClLcUKr1uZiiQEIZ8Q/Ghi3EcBVbrp6mL+Z9CAK1kHN4ivFhDydNn/WkmO0
vWiq7fuq+PzVEfMAMDuUEKrMxY26Er/qs99r5w/LfFAVPcRcF/t81dXBe/7YqUQl
vejTyEtW938nXAyfEDt0CfpJWw1fd0WunzX4OX9kjPy2vSRNdXEe8R03Xzh+sAK4
UmqhNL8sbn2GNbxVepEsJ4pBkcuaax/qWB5M6jzoMyxK/zVQ86rOmFuPSE8eqcV8
RwsoDXXAv+F8di5WsaXKYndR/OX1y3as6y+Plagz1k0qj0x28kl4rGGnXe0nHmfF
sAk/k+gjPOg7MoEyrGH5m4FMScP+ZZab3JXGOldTAO6GSduE32zrgnuVqih5lTQn
nKhIPK02uOALEim4GY5RTd08ziXAsgPpHGALFxcjF7SWBt7nkjNOxJplsLFaNnOG
HrTUtrb/+Xrq8+VVXJqx34E9fITHJ39pbYt4l5U7Neg+6ekGaEzZwqR6c7EmBW/K
OZxNy9bbQupmI28iJHW5ZO8RV0bdUGUbYgDspAW8lx1MSVoH4UhlkbmzGktmEuK4
x7453LuCUDe4Dw9oChcJuAbbmfUfOqCgJu4RdmDfhMPqjTtEsp8muHkWjlmKyMNV
hs5vVxDCwB0Tt5yKwinVCJniCYWWq25tlzoMa/S3SFtHqhMTBQSArNFgxRzIS+Gf
dHxE9i/R2CJCwTkrxyZfBc4G4Hyl0hr7j9x8YeVxRIXw5MBzFi0PiSqczGlPTkoY
OJgZWqMVgEgCVivAW0XneGSCnqInGDd9s/YxXVLjwbRO2iT/mHngwMJl309QF6KM
ZABX3k0m3DOJxoEYlxhnX0KVKkX+T5enL/dHDMPIwsJ1gCDo4aKZ2ByExo5IpG9k
iCa04Xa3QFfQlHqsvKw2PHV7jAKCdkS2Yj4d46uqj83P62crOenjUe+pbRddf4C/
jVNNtn0SG6HVfIyTFWhnWxeXQTFpgWNn+3U5m8Mh3yQvzH6ie+ydgZBkUn2Ir3ue
aVGf37HDmyElJfcTvRaKz5Z6j8ht/Njk9rOtPdAb1EGkvzeOnq9w9AQvYF8jhRm4
etCS/ujTRdHIvVoKOTDE7ovhqSiQBMSFdt68UDgHJMmxD+PcHMv4/uA0pbaW0CnW
ppp622pABg+zQKklN64JZ3wHSIPwCZ+hSwC/QLwectW7sldb8SP5TpTT3fvWr6Yy
vhjJErJnRy7yzsGjNLRRgZpiBJAVeVQP81DcBQVN6T1E+L12oWu0Pm6t9rURRvUr
gCu8lB8BIzhMMaJNs2WoAQZLsl2J0zez7CWWs64uAMcSH6BxHR6cMN8g0YykSjda
FeZwbqqgaZC94y4xpkqvRjqjtNABYhMxfyYvzH69Y6vEBnEl2TCST7gRviQvpDSk
VUfrwWMCkcBPaHUXoEDhCw+WIjxhZN3pj7Yf01Y7AVsH6/s5cy7NT4PO2GyJubTk
8eE6fv3u1oqBQ4z6pgkaP9G31jNmil3aMevZq9KAYLTbK/9bbq8KmLlpXm8qXFwT
rLfB5apS/H6+SGhUuHP2OSFGXg/sdx3ftYyUueC8DgGNj5heu79h/Zb9xQJg3r+9
qwWLnC6YOSW/aykJRgg/XnVzNN0lIS/6I1B5tf6I+3bAm+ZCyVQlmEckjrEVmxQE
LL5FHpkej8d7/KYoBtHlMpPO3P55GN6IImI7EobEwZQ5Cr51RlHW6Rj59HaQlz48
tgVJoFLkAr+vEtlTI4+azh/t2YbWflQeovAc+U5Zny1r1IXek2WzdZWP/g5z71Dd
mRCoIw7iv6luw6rOCo9AwQ24cLkx64XPrrV+6R4kUneaoKX/LIHUg6XKglJGf+ki
B6nlw68JSPYvwu/E89EOi9RmQqoOdJiXYhxOLyxn7Wbh8NwH2HVtWZ7Ne3naA5NW
e5j6q3Glo7swx24d9WfeUGBg8hsIZs5x+XsMCejmUqs6wEaggnIWLNJkWYhvJ7FM
MRyGz/CGjbuB7wNRazMV5+HMT+447gbdTU41AdOXQzDnwdw+3RwAqoWasyJ5rgLr
/1Qloaptzx+FtIpar3V5ncJlLuGL34K39WOYN3Z6XjWC6cljLapPFrjRXdf/veU7
nyXS65aJkxP3OMroFbApuqkR37YuBJYOs3gZnWs8YNwOGmHEI/kBnY9JdWszyMnk
x7nNCDTOh/KqUZjrpRm2WKijziq2LrTrW0/CnfvoT0kyi+zzsssqUnVmAxAbJpeW
fazMRzStKOSf9BXTY22cty+2hSWrppM/wslkd2liNGQQUo+IIS/1W6TV06WW7S4E
+5g7GIk2Eh29H6jDkyu3qjDpAyhwP3xJ4yftvJ+gyPBr1thpc6Vl+R90pVahirZn
Rzyv4ruEV/wCND9/RaSIGTnw88WhrFiNxZFNEAx2xjKI7XnW/eZfihPUAlq/vyHZ
N1ZRDNXozhDFbK87rXdkmIvjG4UCylGOTZwvk5UuANi04TVpgKCZtdNmYMDP4Oec
MH6aAtFymAyGlsBX2v5tCZ/w+04O6jwKR8VgBymNA4RpofImLiWBb0C/EmTpeH1R
MbdtWeLGT+bEJsNxSo7Ih/zTm7mf7ZdfYED7rEHJqj3fyfTqYfKhsFAsf6v8OVvO
bUFf9X9MtZbh/TU3X++43Bvlj0KHD11Tb+/iB+tOm1kpKVSunRzWDqU8p4ujacHV
/n7EIiuVyYzvfP07tMq4HqB89kWcvwUWpOINxzvLxrLFEV+GdAtS9WFly44SNf6u
1K1b+SLt2SicLNr+zLsgs9e6QIsojfCnNNwBTfK9I61Y0QTFce4MTqnvWk/hZROm
jfPByB+/H8DzX72IkRe/OBQmWm0tAYTH+7GpvMCHYx1K8oKEKkFV/CXOxUsdZLu+
MVQZyQDufu0yMDXa2BGo2uWn8rWKuDQkiJZ9plbIFkbvX+TBj/mhnReOvMqRbTzw
SSP+ZYhZObpO/5f01UTMU9PZY21fS+vypfCHUr5jEsoWAz3RiXt2GIaeBoekOk7b
KowRazg2tld6cURaPZPqbXKbeJ370e3uSwMnRk1SKzn8EgcnFIv5ZKPuNBTpVgZX
ItdmrXphZzflWmW4a/MaFJZOErWyfvu4yie30iwU8lXcSJXfAdL/i98JptdHQxi3
Hgi5rJSUJB5gcjnL/M/BQUQHGd/YwOTx01bg3SPkOMyXWKkNJZTCxrE+NcAQLJ/5
O6/paRSEZFkZX124E5abI0G+GfTc0rNl1D1+ZcevYcQm5Y3GPOAADnpLk/wB7F5J
j9KwXuN+9GeQ0xL774CJsEI9qV1r156wDcw7d7tpLtE/QCF3hpolTyO8nsEoc3jp
xcGTMTN5FU6ln5X10IITk1tMBjyWQr1rxOi+nj9mLzLvEyYtVp9skAMsh18p+Xkt
lQFWtUEDWdzA3u9gUEKlYzOQicPCeNLYn4ky4J+695GHQT2xdrlPwDhkEXRAIsJS
y1OIJmlsjp1I+qbxSoWRVcOqAnsohWBmQJkmT65HT8lcDvEuaywRExJTE1TqIUT/
y/HvGXVKil3ySa7xDWQiWdrLXH4F/glig8hJy17/q5p7XdZwQ9oKMjnpGqnkk71m
QmdPkbHJ+pYFsgVWTeKaocA/nuNx3gvtcHPHuTIgG8B5xZEdcJINQfR8yMVdodw1
qc9m2tOrnYNWS72r3DfaJzV4ulWFlroONoY7/T0+I2uMNSp6CvSwrWYrBc4Mx0om
SazuWBO/Ab4B48haZHxNjbIwGym761/U4VsgZIKWX5pFRJg6xncI1WRZV494wOSA
F49fFLZ6J9xdg7YpYeK+qVCi2FSzBAiF2UywgOcx054FNctKuCrhO6mIEPLBfkU1
03Qbof1TT9X8PMAhCGyhVUIDc4HlnP5eTgpOb9MzSAX1z+BEw0aJYrV1H5qhU6Au
nnMX447BNErwxPSXNNVZ0I3CXMa1anYKfBoqLoYW/C+UEkpyqfmIMIFPG+PuUtNc
eo/2uwhSy8V+v0Bgs0s14ePbXOQ2zIG0V/huTy43co13TWEkp4o9aJFg+aSZHP7+
PJFaxukOB5zCM9DvaZdXXnfbm4AzN5U6WMZ9wngt4vEsAPjzkp+C7FbFBOntV2DM
UGRuTHpU4YYjLHO4yLIKjoPFz19tqDDs5QQsxDB9wLImg1yNmV4SU0/Jdy9bZk8Z
hhaF6bfYe77eVWQ/acqnkYU6xsf0UOaYkc/nyHhLP1sB/aTaAruXuNToIACnwzMw
V08VvvgkaJpXFBVmVtwkX1iJsZhPvyhoHlcTQyEv7NYRgdZXI4t8NqCHrdBlIC7f
RoRchL0VU5aGwPPl/0XsxeWGhhihS3/vmeDm9Magf15KwQ4OjaQdiAJnMDW1+45v
n8pkG8npqBZ2fwdzWaAkSW7iDLn5jDv332KYZoPpB6spac58/qJw1ZgVVnJMV0m1
ta0xOdtP8dgXUwZGGAMGrcCYUFYGjJfBNcqyZVZlWwa9Shd5jGKXkcEoyE77gj00
82HJA/KNNuk1R3RbnjvbXgtgijn7d/4C1A8A8v0E2xyzZCVw+3OfksuGDxX5yfEj
7JjrjLRwhLrY+GN4OP4+/QztE+KFq+OHX60l+97jK+r8n5k8WlOa1Cmk67JOmmSp
oh30oCInkvM0Ke5UWuCdYGggxYpjzLTDRiMCO7L/U3I6PFFjKwexVB36FdrFdbcc
rVyHy5MdmSsmAKSaDg106aYtK5Py8iKhvIZHelndbz8QARItAreMNb28Cp1tVf4K
fABdndM7U/n1FbScRgOlBa4W2w3jSIaVK/UM3byYl4IZNi4S4w+tHYrCKk8D7A8w
XrEKXK1Ma8xYxjc7vXKB9gC3XgB5sNS5fSt/aWKUNvbe6FKWRKQVYC+PK8fDdYXo
E0HDbVrKJ2GfqDD97ZLFFDNPUbagvZm1nWyIBKuZFaT6VqyhcXpelFt8JTftOC9o
DbWdmdQMvZo2aY3PYKeU38WmNFO9lS/fZqWhJF5GlCDtOknzXw66kNS3u1gPRqpM
lJ64xqbWon6WekOTvwV0kSfHHIPUOg5WUdMebMOjXD3pzioHouWqVPOsZhDC91x2
/GQB1XMzFZgfoovi4CxnPpAsCt2/LCORl7OsacWQnsDQ1gXzC1k47OII8+KXsaX+
vUZcuc9ZouM9gkl6g9Yb+K/C20H0SMxl0nlwgFWCR4VR+ZeKYCsgUFCAoC/2WrEY
Ldai8AAlNDW2D2mAep3isCpU6ka8jEDBQm5NuaEX4qpQryOD32mlFRzvtjP8fiWH
Minx7Yj4PfuPIjwD+1lYt4+eCYH+NvN7bj+rByibDHViJD6o4BT6qknzmIEEbNfH
c6ZUcnY+csuDnCJ7NcKrHXl//+/htlQncJCgtgSLNDkjVXp/gok/YtBY+EoiUPAA
jsnU1HH4Mopsqz2hqYCeo5RqyVIyW5ydF1w+FglNXKTPYel77EPOuImb57wclDvz
Gc/+I9qRHorA90hbx42ugH6gHf064gEFGMebUzUbXazgaJPGBn/NRgeGVPBbzCqu
APvT2U8IZCwvYSe9fz3ESRLCxdnbPOhLZn7FDjhBEDZ+svAZyH1/deJuBXz1USw8
pTn7E/8pGNt3wuz1XFED0AR0WVqHVAZzFSilsg0DCNqM98EntJKMJ/bQ+Ot5kTWP
u38JNN1ziVezNSAFIQ7lRmMi2f1EImiC1e70ps4+ImvDM7W1GP52VciWqxaqrlfT
cOmQIGrAlFU14GYkW+piuFZf9z7ozdsplLVbJ+IiEv/ocQZoumyyeZE0ryJ1x7z4
caoo/vlOzZbVToCilxEfFfdYA/x0VGBJ+pqMScg3WOuRwm2DgSwUxB76RZiAlws7
n7sC4r+UZxzPIPEa8Y4DQKND/uecrqww9JWWmUianY4/yt6q5AKfbvhr2UOJ0ro4
BzYnOI4Az2Ej7jnyaOumXvqomJlbGy/PML083M5JGxD71Lt0DzOy0dpLrCZ0DAvI
BhKcRNEVWYZyqH4PMLcvMuKZ/Nu+tzCGfuUOGBOBQvacWd0l468HppEyi63RNuie
oEo7UWT8rJhXvUCIAy6hGZtS4wjzcuC15F7i1PpmHFjYTr0sR7iW5PGCXjm2NaVo
3rsXGBE6RCekneCsRSHnWbkMt5H9Xx4+LfcGg2hl1mpZvNO40wxAhtqc1RQLR05E
xmNvg2ELhwgEYAsc2BhUnIWpGBu+9Mu8pbaz5S+TTA4cwgt+cVA/KnAZvAbepupG
dVe1VS6ys9jT60Cb7ig3z9MLZ2VRfBmOzB6vxJHbVM5NPvBWzUuLJdtJvjQh+5Hz
FMczTvNOebnv3EolO1w/RYKN3EcAy2JWAXWP7URNp4S8+OWMLezo9MUP3Clse0MW
MkEbj9u3mdvVzRbR1eoJgAIZcdOued20Vr8UmyVimXXcfsUbi/ly3zA3fPQgLKxa
+cmiAezLDj0bBuiwDK387Z13ZXJqqbfJeWU/MVxT4cMNkmvKXFPPvl12YNLSTWCc
5DGcAAp1WOxLjjyAhd4FYCxQ4pvL7WH4tC1zaNuJd/cDa91/jLNZ4uirx3i9kEXS
N7dKhRppmxr30px3X8TtAW5piJSr4saK0ZE3l+cfju9a74eupgEZvsz/DXPqPd/Z
3/QtqK5Z7scYTPl1NDtI6q6MixmTS43gQuni/kM0lL+jSGggsYT9jEe/2Y/9J6o+
0ZSnwM4nneGNfzwcesnaSQQ3HYIq+5TmOdheC2i6bq61N6HkttspFxGTOmcoRy0n
hoo1EprCDrAhrKD1VBT7x/hrN/MJOHgZugwYadtPIK7O3airJIMJ4jG6b/0kpqOo
miw3FbjbnKGVPHvDqXCJeselOHHELIjXEDpesoTkPRJKg6h+zbrMBs5QLkyN0xym
d9nIolDkz6YO0H6FYkTQBABTJBYr4ir6E9R0MHy0JZFgcH5i8YzIhOTn0eW4D87l
voqBF+gFocegx+XHFdaPAukC46VvNQmRPWZEbpj1jGiOdD/FesWmaoWKONqNa3EH
7pbBTnOHsXgMYklV6+RR269m5wlArWJ+1/Qr/9Pz9MN/mK3xhizhAsJjbXO1KqMt
cx4AeR5Oa1n42JQhUJboLCzZnXnb+lb7axhiFZ09HGRUBRDKDFECuGPElvoE4QLD
1Ctf9RBe70w8rul4zPEuVh9qM/CAs9FMaS8j/dAtExn/gBVTSgIpqXM9fg2YTLtz
A+9hzbnGfqgkylCOXuGCjowiHUcDdrm4+59QLtKIDL4SZlT/JQUpe4oG/NuSqlrz
wJSItfMOq7HBdLuOzwgZG6Jv6FJF1j839poE/KzdVgE2GTRoAYuUMh3QElfGUxDj
INJc0fov9lGpd1gtnAyONuGr0KZgMsxlaupQDKZUtHYu5ho4eHpfK7HYojAu4wlI
fO6BWg/eZE8imofQprPcqh3kPJjwCuwSzAlC0z15jBUoYM5GENUhhNyDKuuLAT4B
FG1soPC1zY7ZME2HBk4W/EQJrs+Y+RITxGOvsKqOaVUikA6eCUhQ/j76vPXXyOK0
5HbXdwCfpbewiSFUI21Bk+PwDLvjqwsdNhDkIG1AgCIHgeYZCr0FqOU61ul91BGM
3fkc4NcVfoeAxifphjA0XbyacF+psAS9Lm9bBqVTDzdvBFqnl68ekGfASnpxcBDE
n2gg0mO7/SspwQYPK/jFxJeYg/1Ns9wl2icWPXHB+TImF0FPeTVu/4KRAL09G1GX
vveTAd9+OPUapFsxa8HPzhrm4zGN3LeUc8pgG2t4s6cs1uI9eRaKpVWkymE7K9S2
aQV0Ca8yQ/orXipQGW2rO0t54LqjXBANNHgpqo7z5PCRKYt3vl2SpBeVtp334QIZ
3MeSXXuSVYo0tXTDCW2kGGhZHmCD04/DZbUHVdN0YPAsjdKG0PoCyjOumqBLWHUs
QZbX6PNgfTNEJXHBQ5T387S37KHj1ovraWLaE10kdvjrZA8167K/wst6bjY6pyfp
Je6P7Y31w5OHyCWmPJMAZ28pfYVotMLLecXwOPqI4SJy5zbcuz69Tom4w/sKvfoH
X2XgnjCYU+b348zwGTXG4C8FMv2LH1LOrcobzDw1a9wIDJtzp4qinZ3iKjbWPNSk
ZcMgDM1Ux72vWeP9wKgU2vkALhAk39OaGLicXPmkIitzEG99Vu6q+lIl8QogmpmC
YU9VPuWmHPEb4HrzO1BGwZoqvViCzfMBnrSg1TTVuEdPPcp/4lPvCn0ud1Hi1qRs
JVS2pI4efFTIZCCQO4We2RlE+rxcKvA9MVnUITJgwmHXMQzJDR8LTueZ9rZ3kWbM
HHVHDawAIF/kcl5EoRDjsFmlzLj1pW1k/0rK1QqaunQvadwR4HyM1I0bht4+NeXu
FWX8TDyQgebF5q70fFV0Y76LgN7xOp8b7KXFdN/YrgN8fXosI/6GRu5V8nnTU0no
vrDaKbyI8dw5cT6RXS2IujNM2683pINQ6MBfzJP2T9IiTAzoPeYoiscnL0EAQa4P
NHcJ6dylrzHXpdr4X8JbDkBFcB7l2tDw5VAjiDCfC6Zzco1va4dDjb+tLkiE3spx
6EeWg9mv02ttoaFq58JfXRmcEFMsXkFFYpk9NWZoGjCkRq2UyXQTrbdZF41p1/XV
IHdTwYG6G/wCUeYlXOqdkYtJmP5FbXvJyR2K+naGBChofRy+Jp8p8W0kJnjfMgF1
ESB5qQ/jbY/G2DSpTg72bGyzNjiPAZl2tm9xAi9/5WFYwZBEppO7Jymc3iTAPHeS
ArdfzZicE/v1z32zeFY3eu3w8+rdyjNvCrnILm7a4/OkONCQC+xuLk1OT+0Obh/c
ltRctG4RUIXOQZ+NkVnC4YDqekju551WMYEJ+I4XVwx1b9VylY4zIkaVtgUD+BOa
U+cPwvJzZKpcbmQsfTHUWM7YFtDhyvwyf927sASa8AXKHkl3o0On1Wh3wSZ01qHq
iH07/5MzlfHbdys6YomtDpTIQ5PBluRWG15I8SHp63vgpMgMm4v85DVxs3k53J1N
JFfYPZJHSc34jWWbw4H0tK5B4/hIzxmaHIw2309+MRQOIs28E/x9sQXvoywBqUiV
eOPiAfO+0ADkib540SqN/HlVHxD5+OIvSrdxOKEZ5PqueeeHp1XIuqzrjXjxLjlA
jNB8CzbG24/nVoCtXnbeY2x0r0k/YaJ6o3rN6ctoHxe+9ZRrHZ80me9S+D/CDT/s
FpDf2qGxEwZkD9bSgLybZaZCzsuMjPpBiXFQjmF03AJVOUkc3bp6N3Z9xmCu6X58
mHEUvUmUjrh7LaaOU0jqz9OXPRDNR7ElqQlN8g8R2zH2PP7C3YqZgt7B+juqSjWF
S+JpF1LVXMz6AjHoHcguqfAAVeY/nl7VAD79faRPc5P2Yi3tOWHr8CCogt5d2AQt
lbuvZL3ShFUSPUe4iF9UmwBgORflakqlaRiOYERckwE15M5BChHzOcNzNZaTP8Ym
NSpmWTRrzBzDU0+VF3BrUtAziouWQwXmJ3UO3Ph1cKPiwTwQPid9rKKT4WiHvO72
BTZyB45FDvy2pks0ExtQWsGLMAFPh2D4q5GDUX4pigXvY/z1S/1EqiW8+4OwGGxd
JY0rDFBmZPZ/vm7cCEFoyfom48H7U9HLRdYtOnIyiKr2O2WHyaof+R4BRAMWpeMF
jTGGBRePJDOkxKTfSscwYgH0kBfYkTZU7e237PGQClDTkM2qGfJZDLxGd5B7mo9d
fSyvvkHnJLIcZeoFkenTpcUYeRfhHLz+Wk9RcBWyFJqg1E+8L6+GZd+nTCnG3EBz
bKzfTNSoBT0qJE2f3djoSfanNja+IxtHLKM3rgaJ9NyK0XnjQysI4DXnJeh/8Uzy
pxCw2wqXm6lJmPD05rVxGS7uRCMSXQD73eV/LODrzNJPX3nk3KDXfkaUunCPzpq5
8z1amNStdm7YP2DtD996P2xS2i3eDURaNyerI6p7J/63klMa0eVqo+tMCW6yD2uq
kDr9DWZrs5btyCoKlkGZUdKMXp+KxyNWksm2MGRzs0Dz/RTtHhYKD+6t9dpv/vMg
PyjTKlX/9XSZ26YYzygFrwkm+QiGl4NSy+OzdCE31nALv//gOjLzut4yNPu/hN6R
P7BAPRxCQEjuTImiBKdMX8Qpl55VhkKXorrqEpW3IMa4If2VuW00YLNW0iLaBDAJ
VoYaSW6PApM8D6K2h3yDmjRuVU6VtrWHxGzUOKuBpzXJZFI6cHV5ppDyV7I7ZiX3
jA7MussmbfyQ0tTCugjiKd8dKMGPGEGdO5Xfiz5zmyqMjQkXLm9HokwBmmMIOCoU
5dFR/xfszXz3cN0h1kO+g1cwWl7egpYRcLRhBRySsnBI88Pzumd1BYqFglOx02Si
/ijqG67Y2OFg0aU72B2WHu7ImK6+Drlg02J3u0tLyfdK1uMELgql7UHjnJmDZ4eo
VH9sw8sPiBlYsTz6+qYfiteIBNa+4icBjm13WW6GEeEzWdfajGokgIKVH9GP6zhj
5p66G9cewnNfZwg9oMX7D0OzcuJYhXXKpwDOo8reSKyGHmhJrq9alPk/Y+iu8+vX
rj7XDRaN8CBDqYCNsoA09nGfq0OgxmzWktC+eaHwLaA3GGQrEUD80zHEYTLljiVO
m042yt8aPylWCoZ+FgeasMvrVqI/EMQ5REGfuw8Q7xzDxlMfiG97pcQ6lssU3Lie
tUejYSkevEWNY5K3JwwxsuAK95F/fCQHpPESx2G1/x0hBo7jaMXCZn2irHj3l5Zm
Pm3qpPsICbdDf1iAqRtGn2ts4j/cGChXsdycvj2urni1HOEZ+lutGWwSkKevfe7l
c8rKOdbd8RBIlNb/U5S7xgHg7OBOXaSCkZ7M+nxn921g11IZRG82zpAaEwGy3TF2
DPvTY22Tbe/c+S5hsHq0XdBVKuu68bBMw01BtOV0+dyfkFOBEY5nfs4J2LUQrIgy
RToha3JlCzzZgF92Wh+pbgQjE1yacdXBk2l4xg6W0xq6HNSdzqFKf24d3C+aVLjo
Tl9XTwlvt6vSRlf1QA2Pj+tpcqE8vLadC5N09IJcqeGSCPsTOyXzoXg3KsA9X73d
TwrKjDcyloGE0Kh7+VSVqJ3KWMU8eBdi+B2EYZPuDthDIyry5q5IsaGNDlH9MXL6
ybo2QE7Y5zP3XkYnaRExDhD+iFfBd70+M9JVURbAUvWWnUbkdYEmeAM64kC12laG
EweCktJTXGXfKwfuJDX3/A0NRV6TE83DQ85CvtmRqUAz+9jtMhOBf1QodqkI4I/s
yYNrVAmpIqhe08sKk91pJI8yFsqaknSmzznoEXto9yX4j9QiQ2TzhBQbgPr11h3f
AFnMftOhqZXIHlbLupWXoHUaNJ9TjzWFB8FIAFNoqpqeFj4cFor5Vep+9oCu1MYo
8mwlAMUHuCempAloLFBzm52BwU8H81TUxb2PyV6YV6n4K09pwmu7caZHF1+fnK3O
Dp1Xm47mFvlI0Bg0GBQr/iNLnhadIq51e3575sE5mmjsEHoojhM7lwYCZeC5oEdY
khCI9Jl/KcZTP8X7bY3cm7WJdfTW8Q34F1UDlIU8SL10ZMEtqlfMDx7JRSi+SCGL
qN6CAQMx704rf65JCZsE3pS416E38StItwhWhgnRIxvExOL4QwjgEPhxtPl8jrlz
pwwdKCz27USKHv12leYxMbTVxN7m+VoliJT/ZIGvGYYbI8l8suOdK9uds1h1s6Kj
ROJ0WqOjRrQWS8kFpzumruosNj53oXhgX1bJMSiyqVZNGepptvyLcs/8QiGuhco8
2O7qG+cyEFXzplrMEaXClOdB/ZGRBzyh6KScLbOGWd7NS40Rlgodz5h9+sCXlN1e
drAPImawGpdCyesnCNwuiQcyaR20HLUkMxgnAu4gA8S+JOmc4jJ6NSoja40oSyPC
ux7HdQEOxIAk9io27mf9NZaX1lXHTkOw2D7okYqfMDEbuJfl+BZYUImO5MlSCVmH
NjncFDreHyu5myqCDmfBcQtfjCuPL1trxIps5ok5uyPhKnRqQk+B76oVK3ZoCPAL
W30KrIZ2xcJL+mnsa58PnGRM1xH4W1VHRyFteD872DDCE0pMSGh4nfXmo7Akp76t
P8V/R2L857pPUPgcPZRiMhXPjb9j5fkgmk4XSajWrJu2jT73uapVQa7+Mez0GmtI
Fmx/ztWyYMYgB9UmfwYApOvQGB5zpS0++RfOZXtivkqQHgLwKfQKruTAY5rOanHl
3xWo0Hbnqo0hnLzmhCEx+UP92hzj2a301TG+bDwGSVWUzgD4AUim7NkcXGglKunp
1PicDENS7yTdwbgKXJQl2kDbjLXQ0y9ZICOPZbGZTJa6YdwtK9a/V4uNbycHlH+G
66LQ8Mk6opDPa1erIctQwTNCID3YIlXVmHNgqvWlCAW3iSB/c0IMlvODmcpzyss8
KOGFKZh5+FixOSooZsRFG0EOon0qXdhk/CGpw0oupE82AxKLhDPQQ+cAdINEPEkb
LuSQdmymCdrD8gApE6+JfAhBudTo1Uff/KqR7D1VZ5Z7zaVywnxjObggkKbCxFiG
YQc3O7rgtuUPNxpDdsl6eVDIf36Ih8IQ5trpxp+FlSYGIrwPDbJLOv/N63dFYcpC
OLN53v3pLEpQ5oHNgPOaFsgpZQ62RkN/dp2CSdDoOmoSaTpbgN2gH/Ozkg2/2QPQ
mgpQvgQHXtC20DbtOqoACuV3efKkxviFESpTQlNlFCAmm06eaSDCfhBdQaBApV/t
vkN2Ed02jxMv/bCYO1TFI+MgAGylTvR0RKxefY4Y2neeY4feoqOrrQDPtS3ZkIXf
Rq7DcWcbpnZKH/1/xwn5qyaahVpGUUVYuF3YeRHeOL6L6ggLdzWhkMm0muNsJAyk
aSnsXVQvR85YeJVXwN0PxVdL7FmFb0lsthyiNfXl5xhGU7CKUhknt2KmACQZE4BJ
roKkGHVJyuRAMZjytQgpFo8hegLqnwq197iWFD/aa7roYlhry0X4zlqOtyNZPsWV
WeOydr/3lTqzgatUDceGWweqfZgyPyN4ag2KSeXAu3zfADV/X4pdYM+dnXSAfC4N
NjkJToRvx4cyJPKbzPyv62lZL+ry5xudyOLezL3wrI/YaWB6D4vC+CD170jqWL2i
eJUZsy1W82mNuqeemwla9aIRQWu7syvMllCr4SeAOWrNpj6zozPEF0QrSGKQlzLC
qrNOT+4eDtYBRGgDfLuZLioBRckbZaFgAICXyIS5TJIhw9OfBIO53halCzhqH/Ii
rfhX7Pa9kdEs+JFjlX6cLqbHmPtKzRlVwAGZYptuZDYAjzjhCnh8zBav1d4nFise
YasvKsgW56oOIVrkrWi1Uq2T0HnPcAX0G+Jw/5hBiKrB2zXA+W8RpAb+DQLHVUxA
E2E9yE/1bXeSjoWgfvUs2NBiWWnPwgnnBfBtbpPAsXNHA82sFjgq1tcd0ce2W1nL
N+jBeGerXdAn4ysLRv0k6wzn93BTL4YlaelbhKnZZLpOGrqq3uWfYnEs3h7ZzAEz
SLYqJake+HGgPfl41mXMlBSFgNXGHOXyD1jf3FzdNpNLXALdWReJaPRS1TWKOz1I
ZkWpzQvhckhI3qkm68gYv999d4TxD7xD5QxQoWEOroM3Cu60gpwBWg88ZKy0OON4
sw3IQ90NtXLQXkqL/4R0+gFQzs+Csz/cI9gSS5aZKNtuoU3CVR9kiFHua1DhwafB
tbbDWRtOXUjuzvz+k6aFTE2C2Wdg/a5+fAyYf6Cninrr3H1bCy659sCrCMzyHCiy
2p3ddEVdRRQjnJ3qgeFbgCptPU7xzPYugi4c9RKXY1pf535Julji1c/AUQ0AdWQk
myuHozjL4hyGkeBD6w7LepBqNrfyOt4ApGLzfLmlAWCzM3f4hiMr0f4ShwEVBHBs
aySEVuNuH2CPCmS72dWqwcH2gi++5sbyJS7YXN9A0Wu1y02PwRGRfoDaQTHopOtP
6bV78/WSQ70CC+BXbDz0202HiOjrIk6DNf2J2ANjSPt4WGW5KpeZO+L5yq6rGSue
+OYB6PnhFyD0Im2wF7gF+pGWmphkG50lLeF6XJpEr9Vjf0vad/hmwJj9pGxWQbkl
HYTsK/+4QRb203HeoCkJl+05YZK4ZkrBYEWwoYjC23bELUQb6NHdl7clbsQGu8PD
+o/u79maEnPSEPBlQvuUipeNtRkuVUw+WbMzbpb0GPqGI8bvQUg7kyXUNXGfPIMP
V3vtaxdigvEan6isP/IVDRgwD2oXtoST03E7HIQ9C2rxOykCtnzplbr0tGwl+CnI
RP5KRnndOSNVg6nStd3k+y7tuG0wpiLzkd5IrapKK1muxrAhf7+Bc+wfhLfCC0pr
VwoBFmam4tVNC5dIH+hx2VSN7Ghu8SdHQ8H4UnFh4YwFvP2EGlIAV8njeUM7R6ov
l3ct0A+dhXyuFPmWMgsFolPWIcuWcHsCRCFO6DfZxkSl/Q5DtuzdpeGwl4mkE+jy
uIPKmJx9ZrK2WuYVKdjXBYLHx86mRCSEt+u/M7QWPgtFC0o3Jk7R3nZWkC9I7SYt
3jS+mZmEycJONU5UrlVnGhn/bf4swmRvubpRp/gzHru0kKji7WnUTFRn0T2dxJB7
Mn1iQyzNLpfJixoNKb1oeHX1vj8D/lZXr/V+HWVYk8kS4mv6G6B7Z25NTDjcvAId
He+z1tFEX+jFTZAXc+J9sBtfwaeRk3L86PO+zXq29dfraXZIjzOUZiD1u+MhkHAD
4GYmCAv+XgzUKscdxZ9Zasi1XN5NHIplgrNMYvUHHwVuEkaAFtM/oYUEvDnOhfG8
3qjDrblMecLkChhxDdQMfQADItzq012PKhSCNvr2UcKJkaik1DMi/OTRfj4kNXW7
EvuSq9P1CtXAB+I6b26RoMHZUoKoKLFfEihDvFeTojBVO/mqPxc4oTfyRR50Qjit
CbEqbuzeL9v3xtZYtYGxqAg5xGadMlJmbyWisvAzn4xpVmowCdtbgasKlUH8HIKc
unKsUJwMkwk2y8/vFcf2N8I8GXS48JMdLXTrhXXyI/c9IG5EDjVSgKIl7xmz+51P
IIU+FEc3Deg7j4dTHYxIhCidUcsfRw9AB2VIH6NaKQIKSNAlsGv92OZ4eyxz+EZ6
2P2ga4HKGcamCkQ+eTvEYQFtLNN74rkLUu3s5KVYtn7J7U91K+hfwDmhOrxanVIA
E6KAgZy4UQw17Zb3RMMWtlT58RNlqxI7QuYVVrHtIB9bqP5/2vXRqjZu6l9b258d
zJSaR9UalkV0Br8TuAj8nsl08y5K/wJQowNn7Sow2qcdYYu0e0PAzYqfjKDxDc77
sdryWz6NpGleWCX0dxoTvEcYPFVdMJXIgLZvRTnA1rWrujXNtsKwORF7qsvD0jMY
Vw2CS2QNKACYUPl2BlZgGgEh8yb8kqkQtN9N9RBYYoVW0qQh1CofvUjP53jqtPaw
Ra1n8Tlpd+1JbI4+j0eboxtO3N7Nf8YS9l2L01MVYb7vwUt2OaVpKZZQUwjZk3V/
zbUnucb6jERgYl+kuipWSi2l6rXe6r5h6C4qpHyKEP2gFllNBicDa/1+Dvep/M+o
qpDBXPNVZsSvR+ngU6tBjQ7nzRBdomANCf6Wj8E26bbS7iMwjnlDHl2FZmqiGBCT
/6yCCMf1AGixB1O2lb3QcFxqaoH75V0NfyyoXVtlJyrPrEshg8WGqWGjLmf+iW/g
KrSEvzy03oSY2QI6BQMBTuMIvYIT+vEHApGYhwBVvzQ6jjRsqvOcPF57nfPDXTa6
0yS5EuaEsMduyvjXiulahYYijoiymz92icsKaENmS28OltLFRec1h5YY86Qzo4z7
QRpr1+ZSrpAvxpmQaShyLH0ipb1FRLhr+Ep85hD5VbpyCDI2fyCkuN5XXx2llXvO
c4vdFFKP+AzlQt9iLMMEfAgEgXdRd/G4fas0cpySVGL6RIPWh1NSmlx1j5OAV179
ISYOpvGV+RDHa8oU6QZKrFMDOE3UCiej9L0cw9qASzJyfEflI0iYaV0zHE2+vK9/
VTCn/AjHJ5us3C9Q0vmi1k1JI1txLSkOxBUB85vWqa4wbT29Y35MD/xa2yvSN57i
XJWiYM+okj5ehDOtlE2cz0BdblVdIwk9P6TNsPnrz/leX03MBpooF3vEwBVlru9G
rY1oYhf/wy4WTXVNUbJlWqcKJBLZDIB7NSdvdalB+O2kiVR2Js3NQBLtbNzGI58i
DkyocvkCUM9BpkSPXKGocxOIo0ZvWWeOgQh/ilSartwtVrUG6rVNaE3MVGB30Ksp
yWTdtM5XiFI7y9iDraM+zlw754xEvGCuCx5xdMJ+1cIsIB5o/OlWzd/90QYg2oHX
S8mmr/oO0CvSruOxgNmiO4KxueTyEzJXULLEgDkPYmId6eUocbch7Prgq/m1/z7F
xFMH49OpeCY12sCs3ByrRth/AyZIj0MZUhTkXzMm2cUq22PSs6U904rFDefEUwhc
eCQEYX5tNySqbfweCbnEo7ufWNSWwrwQREyF3meDxvBzD/N5lJbdUAbz32sG0C6v
HP+jgYocl+Ad3u5nqm4WiM3ujcZYc1kAePKHw6GTRidXaPG4a3dRkgXzj+rC3w8u
CsET+7K1/EBDeQZgXu5LRxsZlfbFq75KzxDLhukB3KTTG7fpOYuf2Jx6en8fK1uD
s2VcxW++Sjf/0X28iESTycBgka5hqOvGWKhFiVXpZM/tog6VgtAFYsNuNVC5VD35
zHRi4DBnZoTkasS50gYlTYrV3HQ+H0ZiAySOgh4uxw8zz3jPY9cd3ckivHt0KhdP
bDYKcPKEM5PIZj5TrcyqD30onoUpBs+sSiueT7gE2rg/nVXPi5Zg35XLvxB7SJiF
LtJRYxzRzoKngefug+oFcIlLhw6R91SGdvf7cSgVpQc2Joy3FGUOm1x+F81EKwlD
PUSfv/xS697uayN8+Gxx7axn1Iqwt/j3urUg4ldmqxR4BljSG2ImTezeWe1+kcqo
CsZvMx6FBd9bo3bNicGtZv7u+bcCJrcb2y2Sj7cfciSPfKwvsqHlrA9/Nk2buwCW
SCrc+XkFMouwiVGITfXF7MbC4ENU1rgDMNYK3KUm/uuNWjMnCYdxIPLqH1oJRnYK
AR567iUiRuGay2ZM1PcmB9VIkzJfYGxv1xr6m6b/WOuTNDAAxQpFjYj2R7Bl8Bnp
AHS2EQ6y3k1S87pRtJcJ5sf+kBOErSGubst/AeMzF15n+ejntFyNsL5ZMeuIAs5v
+c3IHqeHUrDC7Dpm+IsUybCKSU+jeiOKE166lzy/G//bs2HOEQIaZGvb53rrMATR
Szfnizpp7suCxZgdNCtGGnhGsT7rn590ptmc9Cd8MrEcT0db6Txf+dFtQkyKoIF1
Jg3wRxgtiorTqSOnmmR/Eg4WBQBId4fGjNzdVXVP/Yi9RlvcAO26e2GJA/6+DXJb
p57HZ1FSxgUhHYNVDuUXR1NeyR/yGEOGV2ReFFQNYU59dhPG2S12IuK4jD6PBx0T
+08l31C9T3poy7LghU5fBPSHYvve0kHytqdmh7uA+gw2Cw73PjA8yq0sX8QoyQHO
dcJ6UVtDRfTao0Kkp3j3j004VwhsLB+u00XR5hv9JGqEe2BTDsSBUgud233KfHFl
M6LcSDRSQ8w0Mo5Qsfi4DrkFkBBxIHaCurQ79J5FRYdnNDqDIqZvYzgERIkUY20s
H2P2mORDTXWOjV8w8sYL/LsWz8aNG/9DcHqsrFGONUVVPweHIyunFcxuJfURyFOB
tUU49dmGBN/eR4+59eY8EjQHfkJrVzLZVskZqoGWEkU2q9u4+a+TUNYzj99Ercb9
DOhOSElgOgBxjM5cKJQcDsgy9B6tO4z7qQ2GQd5GczUU8q7/dZ2J0WbAdZpO4lQg
Pb6HMdwIaVivFLSpODgQrXzMCjSF5nj+7fw7XJiNp92PNJXEoWaabJJ3U3VRw1tx
9NcnBnkIAnQ4dqt9hOfaPgOjuJZat4vTVdyc54kn4OrDMaNGAp1wtvG02YlQ6Z5g
SdGrjCHwNIrtVoUsO+cQZW8fgejwp9VAnqDexdtS3wqDGrlfB31F7/OA0LltxUyt
WpH+enfLswXG5FduATwvk14ebUzAX9OxX+A07LogP+rGaJgmjKVnqQUZhROpG1ad
QLG+yYm/2LGPnqsN6P55lUxi9qY4VzuFT4U3S9ize0ffL3COX0s3Y5NsI/yjmDV5
DqV3v9QajMeFQHkTwk77JZmhFjmumBfnhQU4q3bu+3J1t9JE4TRDzYHrNrPFij0S
rU6610L9bUixf4FZZ4KVdNKNMeKpYzaP6XzwbXTk9+hckA9O+5QgZhdOx9Ib4OdI
kRvh3Dz0llmUFp0M6nB0m4dYVfWOdooea1RbqgONAkkN+blFSfq3jOiVNcZ2QdsI
R2hSFk6GPaH2fYSUsKrh3cWygR2ULvTB4/xaQn5UxPbXUoLYLmePDmVxYxIryN6S
DnH40xq56l0dB2D4w8ak/D6Lk5YTSSNAX9Pnhc9C5jecpkVYEJqLIrICEhx0b2WK
AksjpL3pJp554+4Sp0KB8QXdEMyXDZkxps7Sh5dvrQklDaZ8DLRV7Y6XDdBTXax0
+22ipwJ8CQgmnVa89Lb46k+0fdbJvYUIPWWy5RH0w9xHLCuWdktrqinfhOl+PAjx
ij8EXOWbtE+Stvv20cJVF1a+cXEkwe/Eq7X8jKO8ZamopF7jB+6AXSyk+/zy37s2
b+oV6HLYOPJ1z4SzwB1h+wtZJ4qUqtSPvBayuJ/+XPvnquJhmQynj23rsAMHq1DQ
gwMHuJRFVdxJJnvS45aI1rRAejRF4efxs7L4F13D6OQkQ6oqpJkHWOq27l670Srn
W36goVmJAS9Mr8WvV9ZIxNpDu8duqlRck22O2Gdw+QvY3hgq3J0TS6ig3q41nGIF
zqUhSxfJWxxn7lhES31ZnAEO2PlDKFHEuJF6TKhlSBEh6jLnUNkwmQLdVgsm9tuL
f74wna9U8xUiWYlTlc85nlN522ydQd/Pj5H+21B4AHwrMfCRGBhLCFwfQOPwQtIq
m+fO3ftbM9NCLjYDOyXb2FfeGkHNzZ7VtYCtsu6xmMmh04IPJjLv8FQ5q+yazByW
O1zsSGxE4U6IHgJpYgZsydrqomYVDYZRdWuHWRfu/3WjTpcc4P7KLusxTeb6PyNw
ps5PSIGTyELu9VR0YuDt9+rhGNrrmi5d3nidvhfT9QSsa2aWfQtfOWWgwKc2X7YE
KDzJUirYpoavwa7yKNLomVeVVF+aYX2swY2xygmLqEBTaDc7/jBhb7BdJCscY86M
B5+DC4WLb6Jk0cbR7rH8ZAM74UZ2pXaTCKB+yuKSopusqReO3UEy8EhBfN4XsdOd
4K6qP9koC11Dhh37n/i4uVZNxDsRvemq/sskbBHaePrjFgJg+yPp4yBBFqOUW2Ao
IUZDvN5Y3mNYQ3lYe54BcK0AGy8ZPyMKTzxfQP1x3UtGX2b9RPHmpVQaZt0aCEPZ
/8g+U+F3ArxJPdMLw973nhS9WRHOQdQgwG2PnIy/RAbhde6NnUHDmlF+k7jTNmt0
vHYquTOnVvsNI/y7gnLwdvuWz+P1748l4jUrfPxMjfUvoHR+R0xW4Bp8V86/9qSW
Fp1RVaUN1PyceF9z0BxpJRMvQ8rFhQ7yFzXrTQxIg7OeHFsEQvnvgj4ZDRsWZSw/
sZOReUS4YdXhhJFfUBK3OPqjTXvXIfvo6odm5nFyzwR4q/QdEP6zRGe8iMwOKPlR
moYaCCVQGImt/h85TOkrEM8FuxEvk2FnLnaV4UGnE7BuJpIRgJWSyFrABtCWWLMY
deg3G03UE/+35ybhpHJ5x0Rckt6k+I+bIcIdYqPqMG+AEFhhIs+u7hRmhMdrLnD2
LM1F3ip27EnJPrCQwDStyyBKTTN/D5UtBB7akAi2WJZKNp58PR99ivVIop7tLU1J
TdElsUxdH3shG4AtzEtRzDh5RbO3324rZNCiP450krOGhgktLltKo2m9Qh6n4rN6
82WCVIi1lAkdDjpbXEp+LWzG0GChuEQqpfPzktL+PspLXdJpTeyjLKGCAPOGoLx2
1p7hGxAUnlDqyROlDvWhlysQbwUtXgFyUWkQEnKsVbN4Y+MUrw1KYJ4SaFk4kReK
myaZXQv9krqcHjGGsBvFk5sClyUzKwpXgOCitK6+9FiFDDqsa5A9BsALm7rFN5M3
VGwNl9GjdGT/oIEJj7YVIC8fl6H2A5yBrGLx07rOlVjZS+DQddEx2VXKtuJRnfMq
wa00MaPh82U5gCjjEMcajMpv1P6Ln9/tuRa17AGawFRh7rk4jeduSdBDZkGtt3Aj
llmvrlHaHf85XH/HIZ0LNV4Dt5njDOOf1q4L1LZOXkq+vx7jUg2c6YAwOQy3eKnU
T6KbC5Meo0LPwKZyz+LIfvI0bTG4KTue7jsDSzsF2CoxizilJFjEqFM6sg5UHZz6
43FIPU32z205EjOLzQ+Ei7g3VU0wyq+THiWgADMCXmz32SL5qBNvPUxzhMSsd6JF
rpx5zBJFvH4e8rYuhmKx3E8wLdD6e9ck2N3Ots/aVVunx+cZ9THUJZFv4b/vBkGR
te8ECl6iseNiS6SkzOVIAm0sauMNjur/MigiOxZ7gbcvDtj39umUYUGqTqJNDNGj
Ez03R6VX6R8WxkEGH/zwiC1msCUQGRFXU1tUu6KM1cViScLt4rhFmhev7call/1z
w4PXh+2ZnbwslB82X32DaCe1XMYTEpf/jrqRUn8Xu5mKYmcU/0lE6RY48WzSgx6H
2DTT7WGpw2Uno1xoDy9QzdQ3EFY1OgplMExdIy1aMZRgq8HdcUb1cPyrnyrpqwjd
9zXQXtJ0PSo0/cnUSORiuFXNGbivOS9aIYYRh3HADRyXrmf0aI/Cz06KSWF/IEKe
s8clUy3Y5H7mL6gng09Lrp4TckOVyyiy0WNMkD+zkcnogNiobMEdFIa4MlGDFCFi
npipSVynz4D8nnYZlWJJxfwRBsoPqdEWVv9EbaTriSbFmsEeT/1VKEwj3f63XByO
BmO0CTNVWSJ2SnojSfu6A/tbO5LmLg5DlFUJk+Crh9FuPLqBmwuOF1IP+s/MZdVB
nNKI1FGiNfi4nMVUhNh2/NQ8mag1lWpZ6ki7XODMLp++osUrx8vmoleijpuqBvEQ
5Dw4clvJurz8o4mDf2FWjHQYqJKN5PYUfvuE0k+ko++q9omvXfeYKAdTJ1YPQWuP
s74ydzgNsLNTu5S3rfoN/YSZn8fJhQPy8+O9vIIkVmvD3u04WVXzlIPuf5ULIRQI
n+EzKVvGb4gzsLM2yGfF/p87V9xzPzTp557aOmFjMGI2tBt8RGtoNvn1Q3fPyOZR
2a9Z6yFplzPll9GsjiMDhV38v56K2AP5BQyf9svyHIGtz6YkFg5P73kXpPZiGTFz
OOZIjnDRW21ko6nsjGqqlS1EZHJP0zauMi76HdkfBLxS29mnmAfYXRKR+VLz23hs
oWaES5UxupzS/vNnsBhi0qKamVndSV78rAdPAUM9wc9xG6lppuLOm6wuaoXpD/rf
Sl73o+8nMQIxAH/uSNzklY9PUKX2YfgE6qmpUCZeqPY/+x/k3G/SjApejZRTpsOH
ZyhHt7BWIyMXya44jlVhQOFNwa3l4BGSPtacUea1dHuDDj0sVqAZQGw7T6laqwO7
miBDaF4tPYu1luUt5/AF5ANjewM4rCxztAXfbKgCkWBPA5yBtGzaigzAKyQvimnT
iFMFu9ZwqpHVmuOiqOw63e51VIknS9YMv2l8BA5WyW4qylALjPtNm8C7nY7BXdpP
VthTyswQdfFd+Ae3nkYilIIMsOdPgxu/cVu0yRl4knLCvtr9Cq6yvZMb1hX9soJK
D4D3CinECMEIUJyqV5m2cEkS6pu6kbw1pc7f48UcYoHCNdxb5owDG7cNyzOKYgWJ
gqa/rMurbFnNCR3sdtnmpkH3th72ucUMB39PXxfmfHKKMgjiAfQ5sbrkFpZHsMnr
CqUGggIiXn96iRdg7BaqqADj5CVOn/tdniK3+eNIys1v70Gi/qct5ZzAlgzErVbL
YfcEvYQxoRRB7dWuwmVCdkg/KySv4GX45t1Lz6VlGgSmp3s1sIBbH1lB06R9n7aB
BNzQ9NBJ30jmOooFH7XU02PbWbuW/HXdAqfQ2JKgfHDziPbK74g5WPTeJn7yeq1R
7mYtAh8xSPDLGdYsYzCqbhzw3Tz7lfZkeZIOyIjMQgoHAvEqmfVNGt7p47KDT4/V
4eKMxL1XaQJpZlr2pe9kS/O8EXNAYgYk9ghgh/8d/gBpCViwzcv+ty6Sv/xePbcj
lRcu644DLX277B2eNy7neEtXxRlBBerUiXs/ddXwjHm/6nWhWfaYbwhxSc5Y3Vrw
Ak1UiPLsnRmblvKVYmmRMMzJt9/JVDV+4OGEB5bF8KPmJU25uWVbkeK09kcoM7Q8
6H/yGnWpWMlVrd3OABbufFtZQXM1odonmB07XiBu/xv5prUU00n2dPcLZ79LNbuu
LsCop7s6fX4emEHp2QH7vdDrBkNe9Qjj1+YTHmEfJP49lldFBdvSDObI92cF/gXN
Hd4S7wN0yEHCsPGRHnUsRPqqunL5CcQ/EupaA/yxSRXuBGlYJw1FGtExqNPFHURI
6z0SBzd+VoeJvAMmQpjDerPElsMyvP0J8L65E2Vrt/Xng9X3lcGS26qNcmHZjyFw
R8X6o2P7ec1zDpJ87Gaj/4ImOuqC8zv2omjRJd/QbuorsNHU16Hgf4HUA2cHpRIK
vm+E5KsH4DbIT95IiK4PjTENTfo+IVqDCJV63EN5YQvfiVXq18gTkAYeC1HN2r16
BOcF11ZVMaNL9R1NM9QwRiVHo/bQKEeD8n0xgNAMRsCM9r3R1tr1gbaUXN34Isj/
fY2FnkMXXCVQ5ExsLfE9+dJins8Lpfb4R1cydpc5aTKJ6HCAIMzbYwzKFGlhV9qR
sFIFvsznJ0RVg3G4WJqOfLTbADmmGD09sUx+dgbvx/V15ZOWbh1h6wQj21YBvorI
nRLqRuTv+wE9VSFI1kBI3PNQ81TUA+GpsiUnyCMUYLY93kX10NsHP7gLZ4Tvebdi
tYakZVl4ysTLCqdtSdcXrDqPWSOIkb3AOP2Pr/lzE/qGhAqErKQvRNkgzw2uLwxp
Q/anH6X963CKAd0v+B2ZziC/2X9iY410hYpmPsqhwWt4gXGMUAH2du6snyj6w0Kb
gi7BrfMr9fQeF/TYwuGqsW8h48clesK94Pn+HSW31feRL9HsaUmRGMk2Jv89tRPz
nUgltlZz7BT68Hpi0qOc5MCU5Jngbqnz+yiqtQQg18TFrRuTy5jyH0yVgKTca+zu
nRhyliyG9EYX8CWFRjzDS5+DINwZ+sqBfIZr1Ae7RmfvzRJovFdvy1ALF2b9R7q6
8kPYCwZNsyHJQ9nhKhFfIiZEVoNqgKc1tADjLbFuKfpwMJL9h5s6gxgMqAiHzaCr
ID/IvAVk3KXJtrZtwf4UD1tYmxs1iCasj4ZtHOKvgThjEzgUkPQVN85pdiqi1wpN
//gy7IKu4KArbqmyopLPX2gLgy3ig41df+jChb8JTDTnY0B39Jgh+BS0FanTRUur
2pA9h4WnMa612JNm4ZY3XMbeFVaF3OXTTwKHGPkNzeBrDuzS3yBYr2/Xy16d9F4r
vOyWItB24uP6r9tM58Zsal3BJFuxld/hnsSwnMwaAqKH1vXcXPFEFs49WbjGUp00
Q+eAMx4wGITq5o8ygWWRc8GLwn8nEXzSAJfSBnKxaGlsrwfomZTfGGAW/U2NCQSC
x4Sh3p2YCTqJvEfGhmUvYU5Hda7X8PnA0glPnJ49gCvtgD004q2mor2tJ3ne02ut
dlbYyBfoxi0DdtMwvN8DtkvrqYLbOBsWQajyTFhS2Hrj4oRrVybcUklZtEeHrnNd
3RQPRCJCvufTkBxWqR5f2Hnvxu5Wzv4CUpzkAVzarwbFsEvviP1Dhq0+OG8xJE7d
7mqnzf4P/rKfRzMpm4Ai6jzwxnAs1yHL5ZlvhEOIMQijMlck4D38CCyoKp5pIQYi
pA+zkwyQsoZ9NDXrccobKA3uWKKSZlsfiXU+71vFJeODwghUKIpm1MJmlxWiPtEZ
4hYCKy+dq3u8+MjPK6sNrBsNN8kTQ6hEF3x5xdJ777zEUDMgx2rNUEZ+nwMq7E+4
sF6h3SXyqV4OrnDmYM4DwTyI8rRjCl9EB+L5wlmBLdb6fgfuRYGlP3KDdguXBx56
DDhuFjeqDgLXMT5djHJYisaysA7IMJzfA9RW/0kxdnGzRaGVRv0hKtyCBkTN3fD5
LmTlJjDt7hCLW8vUrDR3NBQi9ZhrxtEpqU020Qb0B75VhOWiwjq8UTy4dtyxmI/y
eUuzDj040zrhLmEZDwu4Dr5jCoT9IxJQGdDoxOsMMIg9oLUCsqnYrg7CD7X4gWhs
klk2FzsQ8Htb+YFQ9JlEQxgivI+GUfDEnKT6zrGxM2t+5nSE4ALpfMFUtR/5NnOR
VinphSWSQ8z7S6B+hciyCxIBFMoYOi08wx9+KUmVL86H0zprK5+sDc47kCSS+Jmj
UvWt+r2PdzfpBsh6UIge3PO6AvAa2vag5X562xOK80sNJXH/L6t0Us41g8V8MbKc
vK61PcL6qduuxSA7PjzZ2bPAPUEgTEMMpcoewLkvI+xRcdfqeu56KsskFHKoERvN
4XWPYbRdjsHLvuP/gnmYXhowxy0fDvouHLKc9GcgE5J8G6nJ6yzc2jLtLEYM5Wwk
k5ugCaMbRBrYdPDqLn4n4YVubf/lcAtxJhTnRR4xSVpDg3XuDFh6gNsY4wTzUi3i
ytsRledCEYbhLrCqYn24EPdBHAUp8tRYQGw8t9VnzpQw+MYrnHDtYKj8V0VY/xux
ZXfI2pawCcAjMC8UOC0+0+BfeXYiRyBYFhcpSlFs4jOyJ9c2nIl7MF/dGLr4Yaxp
qTqWgkx+oSUMzOX546itVjpf3NY58qqGVfcmTt2GV70YwJmdQby51uR6fA9wawIj
gJ7bWi3oX6VQa9pdkM3y6H4Ov/cutJT1/Xpjil8ASWJ2dvXVo7OWWObl1zNHCecD
kSdHtnFdiZbVSLvZTFzA3y4wqhosmXKLIjktQwd9zTlodeMJU3QAXnTYm63SYQi4
9EqR58cOC1Y/bdpkat338aMPymfkRwH8odL2+WX0Cq/jdiOQRFmvrynspOybp+hD
If5eauSc/3wVulJ7hv9uCP0S5vjjrL/N2egYvLdxkTdlEbcjL98gJcnlhhifP9tP
jb6g5hMf0o/oM8EptccHYRBYH6HG4HjoTaSJpEwA+R9Oz6oXUI2CBV/2TyrykL3m
pGi7PSzB6K0eXhwkDWaKq9IP0R2Sozs9nITJy9vFOCeD1xsX5QOj5tqscrDYNhRC
v8Pw2YZvZ2SLOuavMgG6C2uj0qByg6ZuOCWtcwKr6/ZfT6XUfj/CE+x0EWYDqVM3
/WAyqrMTMqK/zT+1brexC5C9aP2/DL5tEOFAiwKfGSZdY/XOKTE2t3KVUAPtlaxT
iZnpP3fmx6cChFmsrtYyPCRPLaOakQmgooG6oPY2t/0nciq51ZvKBucX8kbDPBG0
v0uc/qk3HuE9PwrH+RrxJuTUAp6G80ueg8lsZCgKZ0LSWj6r8a9i138iR8sTI8hx
662fismLDjqDathn+242O78+Y/ZmcZD8b5fU5GIub1shslQmM0rP+SdC3Rxr1B5h
b3YHyqlmZe9bM2z1j3ax3Y0pqBknn0g3yvb8L/sd0S9OJmB/Lh35C2TPlHl/gF5+
pCzzaYAu5qnXrlRFjBzrSyESD34rsnDS5I+ckuxf/bdTLwkemj8DmIpT2Fqx0lnN
ZPaMSK0xBDE4TQgxZH9YguPQ/6EvQJ+RFyWaGyjvOGnX9Oq7k1f9YQ1aS5eT54LE
3dHHqO1EnXdvxX4pHH3GIRKVqHfg9QwrPPwoJ52rMrlh4+Cwkqh2OFZfaAm7Go+6
spPh4DFuWKVzJVtidGNp/zSUPiUCCLq1+jiP4pzxyfMjTX5UVyJS7jiCrKBRosdB
0Et/ZqccIxxdL017RWw2nvsYJY6MW3jqjj0p4sN3uEpUhhDNHxvmCPEEtSqYUCSq
vuGBDW5KhyvcfJcnUCzIr1ZZu5besHgUUypBlH6dODQO9z0kpo3Op3T0doe/fNyc
EZdnIi79s0OLx1gwaj7Z/NKWsebhnsNFgE4GLcOd7kFnOHGxfmyn1WqTxKoIFiiZ
+tpTOU2hYE1KZIZpDQmV1h0iKT0/LQAgPfy8Ar0boVVQSUIDoPsV5nL+SnGeVlwt
cgooTQAMBVWCd3tCkViCeLeAJr9wEhBtx6tlsZLOAfZKHgZxf54ZRMmT1qduD3SN
/ElB0kKdbbvC1aNGrMZWOuK+Pk1kUOok6kV3Vd/1h65IbS/xaPo2wiWTpIWUHPBT
KFi9YRGV8VU33XzX1oFW2qLFOVqAWBgSQhCm9EjxFF2ZlQQVQuBHqPjM2qd/+zss
R10ysMwwB+RBNNHavUcsRYwiBwBr1FWNGqG8hjpWqyLY4K3bEabKSxaLPsl6nzae
ZeHWGjzkHQDi35a/kTI5k/g7vVAKem/Qiy9s6ZJoyZd2TthUMhwfmcaV5pZaEUQq
r4bCSmqcUwJavrF8eBco90A1mKaSLz5/QsQNt8M5gxOwRAQp4q8frktzES4+SemS
rDn/PvBmrniHAp8CVFBxqwQOgI/lWmxC23Pawupbdqpy6/Z8M/KxvROII5BZddHL
SwsStB9aUoE8bSlFyQFTDUrqv09uz2AmuYwKnf07vGB7jM49zMKx67w3rGIXJ7Z7
tdYhu8fUnK0d2VRd88wplSB6crABxWvYj94r0PmMcxOkwvXHaRYYjwU17vCBVhxf
ON0aq70NT/105bYjkzCEyyv8yJfAyYStTLox5E3MHcuZumBiidwcCG+PZg70Lm3+
G+5VkBDV8zAViXXjA9lU7BHGsXWoQkeeZTKtmnoaZu4ngVz3yLYKWuWqns8f8Uei
bYoR3YlRJKXgP6SwBMapr9rNLNMpCavYvQByuAIBNR5s+xs4Fk4WZByeEUYbQ0Yn
A+LK4X/7zIxXD2zak73MS7vsUn18ihOhlwEkanRfs+sGrtxEyXQFumOF/2XmF7/0
wrTGmC2Z2Clokl5e7l+JlxyrkqGotwFVvuNVd+jHv+1xMlBhvDs5p9407rAB02Rj
mYUK9cQET2L5gM0i5Ls1XBE7QfSrvU53ta2X+6kol1MnCDcbIDMjibxkKg5rDhNu
U1urAddfFT0Qb8MXFuTngeecT2zAWzV3AywsoqWQzMa3maLZbLdK2n+zEUHOXxUD
3K3uN91ooepKPsNnw/PVBKaQWrb7mkFseK4xC9cXPxZNk7PuMDVEDGuiHV8VKpNQ
kuUcgEEUOxyfuPOPhvTxphfdGHae4cxd4fF+CgAT896pwws82Y8bdaHT1oZqzNWB
5QNE+0/7ZVbzM7Pja+vvyaNhX+r4a4xUX/qItgsZmxnu18JGO5L13kKNJh6709yk
thV0CEN1yBu3NsrC0ev9NdPOHxO5IpegG+L6QijAxpnRyRVkCcTf6lououaPNMiV
DBjy3IISDsOXyQhPVlJp95Cw2piT84n9VO35kd3SKNftIaOfzus6r+3yE9AdOWMJ
SXN3eNwFwc7D/dqHSwyO6zGKd74JcBw4HrUTUGRP57gE+jXD60K0veY5bzMRmJSH
4/5xP//mPCZOaEffziFgEo2NMS7jHMeAHqpALVy3WoHjyujdvNFpWL25ao7zEEFJ
pjBbStZPnfHoYv8eugFneTyq/H+9EV+BPj0ph7NglcAn7vYA3tpJaHKBBCRGGFjf
kwF5PRi7/7IOS/ISnmiO3HBChWYV3nlQi+xDY6V1DXAqoc5XxSnvUZXOVHQ0yyF3
cqChycxTut2+RrAZ+TH+ELHhBvE7NhoLzvQcjOlMkSHeLd44DdLLxSWRxyGDtcif
9m2MCn112785K2b20FCjFxMoSbZTgf14IPlHpfv/TI49nMZcnQLHzjy+cj0d44Eu
uGJF3A+2hxuD+3ZMmB+GvDDBsNNuXzCtMEwiXVQDk77m0pXEqJfVxdg116bKxqPD
OMIS5moVjLUxrB4PuueG12NGrtWeA1VtG+zYY0qvHEZJqrsJQLiSUyLI50NV3alM
OUurjNzolFSQwPv07o54tvPbqcpSJeeY8rCRCI7G8CIbPF2kcfCVokaOsBAdr/1d
zGjDPWCJdu5i1vD1vrDXtFqirgll7jsSz3l/nQIwC8oEDMEzy/1/TM2ZekI+88PQ
mvJ6D0adQ2KRSQx4YXMjnCK7Y39bffvOSP/sFA70oQ4+fOVbT3TVk0jIjwaFiBkf
qZjlej+o6/Y2uzJOg2iB7GLpK5UAHahYERRhowPbev006HlCtrmVeNMrfNHIsccA
oJJopluHkpO71uZiTU4rBiwD4ZgkHpht6cjX5IrJPcv6c7SoyhGechlmdp9BOAIj
Uukg6XaXV+JxW/oHiB0+LGxgYCTDk7qUDIKlUhDccerFjuGaVWm1pBkssl66q68N
zxxRLJTnZMCc3/qKVMv6wtswS3a3lj4yrjtazU4604+Mv5ZouxOZ2CURvWWf5VQW
8X6EiOpkN0kwXrDUjf3V7ezfFzelzMHGfGoKYRmNHJGlLtxiZ7ZzmQ4hn1j2CEef
9UvCT6A8+duxegpOiSbnUmOrBIKPsTld7IB3XTsLQQX/zC2UtrPG1wowUUTvw7ui
oTtfdDDKABju742UUO4h2R76OviCJj6VzF5ysuJhqGZ6qc5LIqbo7WOeApRxPVvp
D3wmU0cElbWImmHXsyx9KsObVKTVTiCe7kzpwJWesq2P5BOaJjs1Xv/RTM2plb8V
clMbaMtsqkkn3VnCX4iAWwMV/Nnq69e9UB2JsvDGykozg3ygWsai/IzPxgD/DEX/
lVsDmn7j8e2eTemq4gKTF4RtwfmDK5ldI4Z1TAyMe3/4BGeR3IBpzGYsVUTrEnb0
9XIT+s4h4rbaoL8p/83lHUxII8JdnVU/u0fBS+sq8daI/5WyKIfFz6VZvQeY6UpX
aDKtbV5B2CUIVOPR/R01RsHATPBTvyN2g2dUvjwLsZEL115K2A3B4vDQMVjf6zl7
ycaOrt6FSyLecAG6ZWNKWwMc8jtuIeA2dnpLQkvgTMVfwCof3vzzo4I19/7qt7Rn
emw8ABJG2DDByomUBnDyzJvHU3pZM5Bv69Ib/BIIee1K71POA0jPkdcfLnTqFiTx
Qsb6hPW/32Km/T7jjgYnKjDMVaqY56aIqSlfiGhYbHBcvc8uvcLEe8sDsNB0XEot
5nf0jZA4qmN8j7S6OBeN3S/5UJ8EqvS92HVp2KExDvaWo7l28m+TRJ4JxbMobFuD
nUTrFKZFwiyrW7P/JMIZ95u5fDRIP3V2VNCKG5ej+9bu0JjCV6H9no4wWOsBWYUB
XpObDNXy5SerDEdTidgvu89ImwNOk9EzJ7Snlhhr1qjthbDH778MkeJ/Xb0Wl6fy
OZG0FuYCWgq8zSxO7jOzg/N2cbj/3qR51GS8kIOmctufqnOcnsn9/NWtelDGXgFK
lkc7XSt1q6/LInAJ4FF+ElvINnNAiyl0Pd8zA4hmUgoZpyLJuldejVyLTCVlex7I
b5mIIKgMTVuWmx5mWJkOG7IOOpJsciDEGOZLSjgtz1dQn95ue1P4Z0PvlB2xvfdu
zFf5Kfc8GKvyKjRXJdJBRc4ryTAjtEk9OZ9eDvC4erqj/8IRUdvoSYNLjdXXUoHz
rGCYSpLbPUaqTWkVF2ne9rAYJBJlrGH5TDdZU1YoYvCswXHshwtuHWt3zJ4+jPr3
M1Tiz2F7ef1xzYQ+1mfk9pH1guroN94sTp/2xfemYU88qEgsSuxt6Brxrh8w4JxJ
vIgpJfRr2edZlAhBJ52ESwwUBjoAcLdbE6WFf+kB5+P01C8iaqvKNig0T583oNNZ
Rq7N89m9SC/IArZ9a0IrcNwZEJkL9AkcnPXyzQbNiRviqFpd87QVozoebzoLWMNN
TYBu29b4e4xa8qb0oLlt67Z7tX1ceo7k4lTVV0mBgyEpF2QWSKZA4yKvFP01t29q
be/NFylmF9BIwYhn1tjrdgDilfeHBw3bangbEEBEUGtcXJXhJDNBI7C6F569NGW6
Q+e2RvVAF1LHWOVNrmOLU9/VupekiYUCRkmjzICv7YiwsBvaMi+itE6HMmBahpO7
w6zQxZZdjCQqiwOyL9Or1KM+8EZcQxsFIimgkh5/pWl16zjL4GSmJiiBOY0Xe6A3
TaVtKRbum/NUP+y/bEbJ9Nb5xyDc95ChEp8y2xfbuneS+ltYxIeZDLlOrMrAOKGR
nS+xBpMlB5hOcsG6dq3QI5b6I+ycCvSzC+BhVXaqUUoEbAhB/yWvl9b85611jp8Z
dQMePafhCdvZSMGtiavDIQIfy8LJUp6GtHC8Wn/r+zAAZO+mJ6UkL5R1nc3SBu/2
P5gkTCOKkxy8Z7fOTujGIFTyLl9QWjlYrKEIi4PZzRBq7Jwe05M+vysYY1ofEWTv
Ng7tPwYlz3ex4BMAD8O702Nm+QRVrUMSRRj/xe4IykShtYeUPOT9T4h8phoDj21w
jarpneTDRXdGBCOhbN5YD51PvDiFN4pt84QWuQAY+Tb07YlY6t8tGpCGbiukPa/e
eBd6igwcN1ZpTHYbyky/Wv4nI3M5YDucLXLiIIKlRMhkeKuOc8fn68JBQpzw/fB4
9dEltSYpl+euIDE+lxKbKNfHqLXqyHhhpAbILazWBP3+wfrXsbz6IHS9xcMvxEhc
tfxJ+nBKEq1+WbY3NuPP/+b9QOpC7hAVtKLWfLrZw7STCkltOG/X2WrQN9shIxqW
yrDoUcrbHq20qjZGbWKz/ZTE6w6QRD+wsDQIKoX3fVspXBEGw/iVxS4TX3yiMQjd
e/k6K/mbwnWB2GeHWr6k2k6onpFwmEayXrg68qKamX8hgqtw3diaBtvTVtluKunp
gesx+8l/2Co9VQd13dqhCc73cvhZqNdvAQWMHE8A31EKpl0H7ZTrmjyCflekftdg
omLMeY6Go40PLKSE7GYWLpfPkOIBhB8vmMx6+9fW55Vc5kt78qO6naM+ZpCQVLI5
rDQmUaRJaOR7dlEidoAC5bCD4R6O2B4ku2lfhl2EetBN9B2b/SvZQ7hChHRu7z3w
aYo64J//ZvB7Sgt0HfrFaaiasKbDZqtdqix8US4+LJnEpSTk8MNd+Yuh4Nh/JR+6
i+WmYyFV0cGd1vacucF+Xb5mcdKsuKOnMoyJBFAqcKXnoS1vv3udJVrtliA2YGZt
hkGIMlqQqy7DtQPyCwZLzmInNfmq8h83mV8wzyl7/EEx/jpvSWIdi6DyW9eb5zc6
bniRTYodwXYoclsFgVaYs+99cTGP1ENtUWr8U9E5ZrZuDKJ5WKjpD4sPAzu0zPlN
gQe2JXD2hRGyjCMoGv4JOLj2zXdDn6d7s1vKLqDDUvF4OXhnNyiw2EYieErPdS7v
QvniGjDJwaVK3iDDijSdRwbiDpgTH9hNlG+O6LKDTeHhQzImqcTTtlShlMDMXUjn
Qqfo175IBw9togMvOctYXrOdtXny0DIXTEdN0I7+AYYwxh5y4g7LAiRcS9Dj+7CP
ZdFgsHSv4CplO0M4W0QnCsET9nOrFJxg9vmiCBFKqtcQA30nl0gClpE9lkoIzG8h
X7QQTU0jG7DAftEWRK8RM9bnzDyvWL/ehb38sp/3+67tTUsZSr5JEd7ajlR5S0ZY
Mb1bw9/KBSmyYJD/agfAKaFEzEVjtR11HJldM8O1xvsLGnQqnVB6QtG39JpJ6+PN
Xu8F2gD58FFcCemXLNI8NfyFFRf/8VoO/ZCe680J5zVAbP9d2wJ5btFrbH6h7iZO
PnaMFTfuZ6UTjIkcRWk2+jeeLBda22sd9TA4TqsYbcNpsWdlRb58KGs/YxIoYmco
P3jG4kSacdcvBSc+BHXxpTyiuxwco9/MR+s/rvaf45icOJjUUNoxaufJ43RYgn5v
LS8mTOoId3kck16RVEnjxuruaVy8UoDhNh66Z6XscQleJgtNlQNgG3oKlq3MiAxk
GPnbSktpygr0bmh3dWk1zP+JuTy1/yeaafL8yRRzox+42LPLyi9+6xJ856G/nDDm
0qGRE6qIPjzSZJJusNMHdsXB8Ls4GqDtstzQNaSkOaf4/MmVx0RK599jQhZbrWcu
ApdUkKXNm6X6Uxlu4PDrOBl3AY/a7h4WN71lhtUhdipXk+Wxa6BKvyHO1mrRkObZ
ef/XqvmZpJB23UlQub/6tKQzfw9gJJvQmsnlqrWDt7rWJHS4qpoQ/5+N2rHGLKXz
InEJl3fv0IIoj/CVHLJKfNcq2uXZMrDmnBinmKgM9wIRWYGL1X6Q1SOR4J8jHxPB
aitKs9dbmSx+I2cyXyxt3rm1gProXoBpqKlOBECrbk6s1KX0XD//Lgn5qMiNMbYB
nACP3oKcMZpUvNYrUhP01Bn/WJRGFL8zYMlH0q5oRUOUIORu5Dz4xHeQJdAsnaM0
ODRX447JnwiBZ+DbN89jU2/l9DBb+QRUC5VDylqOCHkePvLxdxTGkLUHvbAamRe/
1mx1ndsbvXfDb1ZjFhUdkbBM6lLUZ46+19dsC2gtj+5gUg/tUzHo2pZNX/Lg7g8B
gN23sauVcr79ujPOlY/RtTpUgtuZydMs/Pu1m0ys3omX+gpzpeCd4Rp2BIU+hqWV
NfPgh3ZMpJf3Yq3PYO1AjSIMToplIdlVq0mDJT3MGHUvj30j33Xlh52U32tc3fWL
fgOes+eNDhgKqoKea/W7XeL6U5k4EOtzYr/0DxK0MVYXzX65Vqs9FnFbjXqM+6Ex
CcdOAa/VNKyULP/A2IN/xJJYkSQZh4CEUP/bzTNTXoZNmxEm8s/a3Nd6LMF87WNi
2dqjzlVvjzVisFF6WL9q7GfYHskWvJ+oLbWoRkrj5ndg2266up44j8ldURxsv0r/
ldvLpZC+KmzogUPBh1HtF1/lF0QjhNlU5nH7AZ6cs9BFZCNiycxOVBi5FLsmFWf3
mYVnErgEvz6r6oIjVnqNkbbNc6JpP6q2PU74xJqdCZHZ2GXv42GtGSMY2nFxy+4U
GchA2gcWNUEmwb35Fgp4gO2CRMs251xWDKC4yDtVbHEcPJ0YCpmleHKVwo60Qfjh
JK5Cj5GRG7sR3LGyYdI977TJHsog2MSIXSVdKvtqY/4D0XvOeukK9tAY4nUAep1b
XiQH5+Ofh40FFLmut4+AivNwkLCkJpsYcv+mZLpGH/dqtrTOYsqy97p8e00VoQjP
L1JHIWRX6u5L6GnSzHB+5CpKzZpO3N2BcIDsyw3HbHUJHrIKlMBXgeyOkVbVJGgI
CLT5CPG0vJppws9GtgokE4NJkmgZk8SL6ZsFq0qvVq4Hxvjof95sUNKVb7/CCIjB
LEYOI8jLpXX7IDzZUenB48qWaBqJ4PqEFwKiGbmvphTo4Iyyq8CKEwePY1BbZCv7
WGMWDlWLq60D6YiLLu/QK6RrM/nRX/7ADTagbTYkclnHqT3xl1McS+K8q6OUcrFa
wVwrRR7+Y54KRiqR8hdxQy5w/IGFxNDCSZJp/LJFrG+pAmhVm8fgrvRlJOSc+2GN
8CgXtWmQxay0PPdda9S+5zHXu56S+YSVdY0nV7TUXLpm4uhJnd2sAC2fsSJurTPa
/cbaCW4xqzEbxEw8A7qZcFoFvRhEMv9Y+Wj7xGcOD9KH87r6ItSYnJY1WAOyb0pC
R0EpQtqvCh5cVKToC0OuvgXboD9eaPaEDC1MnMT6VpWEAUDxeYsmfCQgiR/aWzih
Vgp+9gtGUQRKBm8u1r1kB7GohZWBJ6QmB7hDco7mQDm3a2TCSfMQ+ioeXgntddPN
6rCGQaNmpO8tzGGg/6DarDPbZFVemWRm9516eZNlK5qYHE/3L7/WNMa9OwGFnLxI
K6gk4MiPijn8OXwXgtYHNBragekOZfEpxRAg+qa6YDfTi/is2CNhvCNuMDfyheoU
VLobC88anGCTB5yQ9gJFrZ4z47uo1Ayhr5QDRcvQFpdzSi3b7W+/ywMEL7s6xPsl
WekgdcTicbamLG7vZSGhPvzLDbfKaJiaPRnzpX2+kbdSKDqEsJjePTcJ7gjFX+Ki
pw6hePvNfDcsy8avqAsbqSCdRpWJUZod9VbVEVLSoXOpjfW+MFwt6jeZGxTyvewb
kCPJRtdNbwrhRMvsBUem9PgI9tlBx1h0KlVc+seASoqgZJ+TMhCKWn23bxue+/6I
sFBK+tFlx8iDMiOclB2do36BBZEXdTMeKdRtc5aCRe6PwT3r99n+ToNW+iAfmz1P
yncfS5guGbSrx9KAjN4nWlXmNx4a/0obnRN2+6/uaPxPnjCtz740zF2IjQWBHTR2
Pk2EtzAr6gpn0pOpCiavvTuLtD5GKji3EX4MttDy66+eyonP0VGaHLys/0RoGVae
RogRe3dsdIgu78/nkQingmsmogybYITfZP7HXwlRlgUdVvdhVqjuZz6jV2a2RCj+
xA+J5O8ZHpYAZSkvx4+1qMOt/AZ9u3obAofoqa+es80+GSo77o7wObsgD9lNBK7i
zV5o/unU+zXx/0OyUATkqwAvM/YiOH7PmzAI7hBZhbJDie3vW+QWflhTY8Pqaj72
81+ZqVpuVwIvlurFNuwFBNWf7031abGlhSqIqF1Jl9dryVa7kJyB+1ClxBQzRrQO
4vM7Sw5DRhT+KuTkzX7PAA+Lpt7D/aOPZhrdBxihphzGC2ti2byQ/UbUrTMhXrAH
LmFJU8ZG6hGoX16ki9+yI7pnXJLncfJDRFlQmNxatoV43kJ9Y2GsOo03LAghME5z
B5a4Rv6xHII5VDshY9OPCCuzi+2KzEpfWjky5DU5Yy8W3xKSGueriMvd2YiyXNdk
0RL6fnkMVCZK3lYKko9+n58murr0ge8a8xgztAcN7hQYej3MK9hvD2P7/Upjh4sE
TK/ShkSZ1KJAX++eq0lWD+tnBIha+6CTX+cOR+mwV7U/Bp6SAG2hkqT9xFEfAePK
/rVCcndKNyMd7B3EeWnyL7dycHUDYHuqgGPyHN4u7x1PIi9g93QEGBJ03k+NIG5j
zh0EzOL6xTLVonoRC6qOjctAm89tBfRin7d2I7oNBkuyJ1k1zzMr1dIfGVWN2EVN
2k4TSXjMeaO7XPLRkbSIzyC8I6HZmRC2zvSEvgqhthxyfi8IloFXEp6L1siTssfA
fQmXQkrXizHet7OwNp7SP5XFPacuUgEKOPWhDYxhV/KdIa/NvQam9qih4/rSxNsv
iVwG8kLN+YXsq+6yKJHbD5ThT6spehJFAPxfuJmWDtwBLI87CGABbCNkWe7q+qsd
yBAaDbfIJt2HQcL+4hOgtUBjn1YsZPx/sXk59VM1Ln0o87NtrTBgYIVVNErQiAOH
ZWPqwseE3cb8SauyKhRtoRXvm2UIxd6Td4wOzpo5USuNChJEDu8SJA2s7cI7m4Yb
MblR0iIH6QxSaRByC3GvJHfBoFackKfPpRmghF+4czDcDJW20u1+CN+0pXfLu2m1
K4WeeKWmV/pzirOtBJWxsytDrWkANzf3mZ93x6pz//rS5Zqe3kUhLq9uL3qNtQYD
bLVdanT9hRzs8HcPD0Wi/q5FmRjzZGI82C5Esg3qMjOtoT1N7L3qs4ymMy6t7br0
7FweiXNAMvJUbVLFV4InK6/cRTgvAb8f5Sh8jp/Hsc2i4GY7nZ/G1DstIAc3PcQl
7TEqlz2BZjM+XWeOf9RSwfEQjn7h6/f8d8KSpa5gM8froNZRmqbklY5gaOTrGjl5
jUfeuOhsbBCTeRS3nYz21D7KxHOBzpFB6Hb/M0FXl7OwgNLAW/K35YPJYjV8No0J
r+g/AuwhrUwF0kKejyAUaquu8ax8vW7wt5ODvOwsDHF4+TWskhF/kBasVBaqGxVZ
3puZC6YUO7vi4KWrCbKm0vv33An0ln6gNcnhM05MrESK5YZ7MTrHRomXhBddhLoX
sowfBBPk3PBsow1t8rCraY2Pe6WiRATjIYNZs1/i+mSm+/TvJgPQQg7bF/Sdwuxm
Rjt5mveImT/fKQWJOuIvkA4v2mBlGQwS+hTQzn/Bwy3zH6+MytC3nszt2zeAfTcQ
DH0QuC34+yPPxaHrFMcptylseEtHRoJT2VKXFupBMaLXwYE4sI5XUgmz5JVpIrKR
bws+KJOhH4weRRKmK5bNTN2Mz80plpxkjmAt/bx2EvBm9tR1zrv4rOeSClqtKf1o
DVSvz0yDlyA21IvmfpFf8IQzkXxZu21j/Sv0r9ZhcdCwNFZSe2Z87trhDmDjkZ9R
X2cPRrRkJBGSHrlRrHeTBT91ocNbslulramm5Yv4xyKJZyzsoBHSNYGV0nwK65LK
eLMeImAe4nDJdvGSAc7bkmjWc6qIBIy1lNpj1sQSloqXVCsgbZ7q7QukRqyZGjmk
CPY5j1fgO1HkgBLwiqsK1kBLNoPRLulSZju+vck2mS+pygWgwyfWg4I2sFIJKwNp
ISwztPbPqJFn0xSsqk4pC6R9/oi6KmEv2Lymtk9h54nzzFVsIN9KllN860+qDkvF
6UlEipljlxGfUy8NElkXNBp9CNLP4v6QS2t2fV4CD97XDvv2vjPcEJyKh8V8zMw/
Xz5tW65SbN0nyWHUhkT3gXFFZ4r95cmd0cW8vbCzK5tG6qIKeNZBxWqAwuUH4MdM
5p0FA4UjwPNzqywOy4Dv2g/8nWheOp7X0AiYNW7e95/U87YPjBygLEfBPJR7Gy0Z
1uJ5nPvPsKtQc7V4YHNGRKThLVp0+pSBuc7CSOaIZbCr31+ZGaKUUnCUTFHpUhAw
MU+jKZmURdEaBifLEoR0D9MEMAbI2iTQCoq3EbI9PyFykRSd2FoNrAX7kbsV9ZVv
HSXCNYwiZ1EX1nwdxbOSlZrqzxGNusQH6FmgsGbMZAc/GoFwLv4HmUp8TClChAV6
ecaB72FckpZNJt9oUEr/FIzUXSeYNI90y/89Lylh5+0ndx69MAIkpN3s/v3nHFJ+
eHaZk7nRnJsQ29c3uaulYogdvxhSbcwiHHr17ZxxBC3x/6EYAynQqlWtcBfARBCz
54RH7Rv1bYaweJe/s1dz1v6Le3DtFMZWr3GK6wU5cNLaqwpp4NQuT2ZQvA6ThGSt
cFWTqBN5Qln0iWhI6+4UdnVHZhy9OF68RL5IG7h5Z8oNn0sKhifYRjz7buduhDEH
icuSPGZLSjmHAl1Q6QsUMXS21ZOdpb1PSPZ/wP0rKsWjhEoSGoVxN9D2Y9tUUW+0
YHR54eDJfBQptlpxMHCldqqRjoHRoak/Rlq2on0Yn44yoTz2qNN54XGFdvTKYtBS
/ryQ5KSrDuakfF+PS5E7x3c1KMLolZA2e/S2d8PAMqTWAethyy0R42cev2hSHtvx
acZlCuxOOxFsEWJEJtPYh8Wmo+AvFpSmHH3hkkm7bqM9l9hsTyGY1MuKGvi19ETk
jFROwxBv7oi5wCxDQHEeYwFnqYb6WnGStab3ZI4pmtEFAVlL8YxVuGdI3dDlSVLQ
CLlLpF+nsK9wnVX92AiqahsXSbADfSD/74ZHWsam3reslZm0PWdgT2Rn3MW4i48N
P9DsFo3KWKIEShAlNhHTnP7iDMFs6t0FbItIJbZlje7cXGtTBQw8jK3llr9XKvQ+
zDYIKsfOadh+U1a3hcfGUWKWrLAcQgRErZbEjV8BMqXu71H6pLrcNxuT3OqUnoCm
woIxKVCiMoA4APhX1YFgU3jIJXiR6R3Gh0cWY4DibFpOGAZsD30yXOKKaweDykW9
/HWMMJOUx6y9h7EN0visJ5tjgqmiLc7CTmx3zvTXTnCd9zjNSZ6P4LDxvtSm2lDm
mks8JgEOPQUmjAtUcU0QJ3vAliXLqCo7U0OnqxJMjd087iw8i8qnW4+NLYwV11nS
dWxAtTBKFQsNczRUGi/OHykViNeAnHMV1cG6iIYCphU2FaH8M+MzXd40XrLsIIps
kEAk9otXB1HJHM8807x6JMfildyGq3g2HNlYR6I1xwyKE6AftxABVKaQehXUXa7w
rd2MnfeLoPlFSwBkdTJlmNGCLO0QSWPMhkYGFQSVLljgJLEEb9a6pR9TtwZ9VRLN
+2wZnSKrSJIoQfwPkh3hiRY6BPqhC0lzCxvJW4iuf1ptkBN7GUNhrBbxiqIXFfgW
CLxsIl/NY3nVAb3uSxvSGS9CjacVSIG/CXgyzRc2jOzFtLv8rug7GfXPM4i3knBa
I4xj9CrqQKSE/moCG06Z13kqivCAwqWV5EPhPHe4CfEKh+HYpjaAmMaTiDXAd5UV
ymJhr5kDRzGkyW/y0AkXO66nR91NQKfnTje+NFoXVmsh21zFOqgcI6J6+9kh1+S0
nbAiUX/fuxHrulg0u0NHx6Qj6efqvkpIdZoxbTVwu1Wnk6nYh4jYy1u6GnshmtDZ
lV05FLOj5H/hyU7XcDQBerMPAJyqNoe48pmH9v2PPnnxN5r9uf7OTJ3BLRl7xdBa
5u7NFTJ88jY1/xH9QBJcvDsLnzQCiJmZQxz0qYucFwcflql6SvgDlVWd7kf3/R0K
ft3l4HcIkVZkhD9eE3IZriwZUY0c2VY3C0blD6vlFpG/jFWLirFpnfzs6JEcMFmJ
DjSQ/8pDSwP3FFVTvzBXLIyPGJGJVYgENMq/2mLLqLbMs5jbDZMyPR2uDUdtCYxR
5ZDhXhTx1pbRQS/Eux6S6HLkpiTAzTZnIipvOhUZ+iAuioMMiTaSn4WKkX6OB2ma
hC45vc1wDLQyk9cb2Xlf84+GIJanJQDS5bzadXuK84AziMXKeBrNDBsoTLTgSLsQ
g+Q9mKh0giPhnP90O4l0eApRMYTabfH9s9/x0x/DUDwUl2Ot0Mh3l2YyJ2yhmah9
MpDON2DBHLWoF26yMp7snAKHxiz8mwwJ0c/C2bLqtvyWpPC/sEmorUrdxIYvLWBz
hYgBeRxWSC8Ogwz9rxhURhqZrcNmlCXtTlfCToTvEqhSaxdL1iyzLQnopnivjoHz
sirGzpc+gw5Awst9H/OX0DQTfFoCpNpinVQRr9nodQECQoMOmPSHUx0gGIV3ddRH
M3MvbN2B09RROKhq/5RtAtVXMDhE4oakVIlZ+VhbiqHFUgiHhUDgAAkfSrSb86iu
9P0EDOkv53tzCnLuTMbDcqi3celIqMp7Zg1zIuMgp4VITixO8QjbxE9pqQoqr/BZ
nKxr7CXAp3/QpH1J70ejv5qoHw+86NSgSW0gO1XmmlklbPqv1bEiw3rbjUNQ3YsR
jOOhDTnDm4g5OJVDSsW4u53MXR5hOKmM0XxBUTB2XicG0H+b6pZnDvBILfxNI/o2
87TXKpKOiUTAHIehhJhwvTHL9BYxjexyKO9CVaDOX3uc+DbVDYPlDfoRG/3ZVipV
wqtRauXbasUtQlyWQbCa6hBi43T+cLZbAZ5SHJJKcz6TDPTWmTKVE7jJK+dZqtdJ
sfGlJ2B5Qil/WMJ5u6K2vlhXaamvOZAmH/SLN7Qu3hridyMNrV4QK3/FBK++nc6z
h4Y1D5JgsDzXNLYS0rnAqVB/bTVmvpk/KD3jbOrdmtKY7+0pWbsjEF0EPdzVYoEZ
HvPcigIo45Xn6hmLNEzGJWtNEN58jeOnapblbTW3Qc4pTjahQ0iVyVlESvp5dAlD
YQFmCPeSK3KDK6mgxCHiZ0kGIMbufkLPKYhk5kUo7hcx0S39voK2coFeM0oN5IMg
GdaBWCOeNJkbHxQ5jjqC0Ft47KjBgTIl3sdFTxCCb4LE9VGv0crhdM0+GLB+SWql
+ME4KqpQg6i8OpZiH+wvmpIWpDF56wM6bABLkb+EK8tppfyJPrXxVX/sP/3WPXpH
nwOF7LN7jmAvrFSuMxofaw2kVeIuJo6r+8jiUb8D3VQSGt5sdblPLPPoE9y5URF9
WE6vaXDAYZH8anrlREHqFjRUoE6UQ2VpSaWvln3hM+Tzz0PT1EZvNMPjB/iKLzn0
aWebMBuYfsyEbORvyRiaV3sBud9WwpsxUbpRhoyu2Ge69RmnFx2pV+ZDouKbT69f
6YH4SLeWVxTTurF21KhKoOKdO6uI51Y4osmBqtV41QkWxYm4CIJOIUAvKZNSpwC8
PS12AK2fH4icCCXY2q4EVQsdjKo/aRRvsZ7HNkgoTAw6HptGt0uiVBqWbNs45egl
oKD8+Z8Fij7LVqYUnF7Z9eYqIaJ7s60czsT1xrfjfreqhbuuN+azb9Ja4dJR4egO
RxXg+ne0gOa9iwjNhxM0TMh/gsMdErdkqHJ/enwZtu4HOwrCq/EOUXn9eUjZVVMw
8HZIkjvvHe0lYg+yphjBX73gt1Wm1Lps8x15v5F8OjXPAA7UKcHU6/TLCYdbIHa2
HP0YVVLBn3vIYM7GE106B4OhriqU9RUG9wDsnRoSIlf50cxf/yEg3niKX8s0AJFt
4swabuVnS0Fjmv1vcbW4trKp2yA/iSW6JUS9Ji5C82CDipuzxqRCm6gs+HqXtzx3
S+pNIKKxLZQXQIv97fQr4IWQkBYUT8x//rbOwS8t6Om/INjxhphbYEM9SxgQ60RR
7hsO7MAhCcaE6E6uWDdmJRxsQEuDhd4HpVPc6Xne4ZSw3/aNHioO9h7F+GPilfAc
1BSktzOdZ2lwkyEZrlQ9bLjbNxelllpYGUQLOsCL8IsPWrTn6DZPib5MQpHy/N1H
w6PE2lkzx1/cswcm7ZldnKlQEbF9WvzmoY7Hsz2t+zTokdU8n0zVo4xgZcZSx5td
L4jgH+agdNvMPA047GAwH9Vecid/kiUkMvCJgaAOAlP3Y7FEes0aqOjnk03TXYBs
qlBk+yQoYAV0gBMyCK54pKciaV9FpovFPiH9gd8tjqXbJ8OShEOfHgM5yeKYVeRU
ShHwGXa51WlttK/bc7fs+FdQucMRDeRCwt6D7YA0nUWB+WnQIyQ1rrkYn7kLfegD
A9s1iwGNI6EkIXZvbH/aYOnvye30HMXFYbWtTn9PUaB9O/mB1QsM7ZmFosbt2uVy
TyPpiIvrjCgcva1MvPhIIZzB7VHQEe07Dw79dNVe/scp8E6clgcq2w4oxn7mXEVP
QTSunTC5oGCuD+EdPgaPBNYXeD0StSyNXaUTnv5N8+81sBJmUP275CcG0qCk/AdM
SGVJBUUfuCg0LMLAA11gn8+5dLnySEc+tRHrtsGZiVpuq5jaRMDpS2rAyv2vuxNO
SnmVWInDW2F64fnARTsYV5arKJ80ERqttjnWwOdM+ycBmkUOevA38Eyy3mQG0Vs6
zZOhPQOi97nFdXwTsE9Iy0RZIrzGLwkEHh25Dr6dbw31SH/3BMnN2y72JWa2yxcP
5P1TUfCbUtDvWez56RgwEIqVPIi+CQKGkhmOfftorGnXJWSU5yO+XvN2dlpOoVEt
6Dfcu3fvb2oakjJUJPuVzGKxaLeuhRyJnbJhAZStVYwROyijfKEhn1W4W/m+KlsF
gxpJwtmtcjVPG4KokbSX9DiX9s0uL+inPz7UNVzIkwrcR5DS/tAO8oXIwuQ6pD7x
cuSYzf8lQp0eipXiNSK/9K42ga0YZRRUQLO04korLTvcJUxVRrbz4cHzAm+g6yX2
cYffKt6uKk7oVBSjbEk1ya7o1HfF5hVTYnPOxH7X6kpRFf/M05Y0MRBz6Ha69g0D
9HdYN7fLcKZlCqZMXOpV2Y396RHNORHmLDDEqm0nDwKna+P+G9v3Xbm4HdmhPBqz
QvrD+ekAKo7wkTuwUEAxWNj4FLdLnJzYFkq+J5fh1JvdTwreiLc6ZL0OGTOthX1B
CJtK3stqhiWJHPdcDoOIHfyzbyTm1HjyAN0e0soix0c6UWOATw0QeVS3/hE8x9Lw
guSY8gkHWXR15GyBca57Idih15P+smaR75UtwybMmRRX43PcyKe9WGo5w4dHTVoY
mD3J+cDFDm8VMLmaOND98O7N83RK8ad3Ua9AST4AA4vEAleREDvpWxos2QiuXWAb
meWGYRvT/ECv+Emc7lufb850tpwvpJws7DQISPerQIB2egou+RjLNGspxvQCgeQQ
gP6d+mRPJO9Q6XOtt2o2c9PoFTK+kWW3lvvISV9nDaDiljjVPifXF7V7jqrlcPzA
XTV+y3bV+u9L355JSYqCSV4jDIr8mqDI5haHFHSsY2Iud3W27Naw0uygvYrusiSa
QTHeba056zmB+U+TXHw5vWXKRYU4FBYVyXq3GuhBW9rTlQkNXwAvPx2RNrVE524a
9/GqRqy1fGL73BwbWp5CjSz+nto6r/CF1fmbNiGAzXnt9ZW3WYsFtG/pHd/gRpd1
ZO7wqXTI5+gMR7vVUyEmP0Pv46moqxHYt083gZFJ09SLttBv3i+OK/nropw/qyGz
6l6m4YDU4b1S5BGQ9fbzbPGjBJfkp+X7Ah6tvdZb0WA/HTH4vd3ViQAf9MDtZ5Gp
jWmCqT8hLAqVeaMSn2D0N6onHBJhL13cmnPchMrcevgLXDNsIh491MrOKP/Yneb7
hsga9Mg3CRmo8FyRt/JXEBk2OiOnUCcBKKI+FZ+TkjA+8jxeE8MP/7mEa4pZpStP
yq0xXUdB3YRSy9JMAOwOcCrjWISr6oYwE+B1LE+Z0XFFOstGVa7tiicC3hi6LU5Y
6qivWGsr3PXz3wqgnVVb89Ce+HDq3NCK1l1EVnBiOUjrSJoYLhSggCyuec9XRgix
5+zOUBRElRKiL46lagJqY9yHAfFdlGzAjYRo5ydqKyfaANc2yrWF+Z7PHtXeMbPU
TsQwhJFkxtL8FeEmVAbo3bGzRqvq/OBX2B+5Cg0rMgUoUQ0s79B0MJ+13+C9BN3N
ox9IMmy/tJau1oTJixYx1qH05+4/a1hj2ha5IecileTxf1dB7xSo4wJFC6YW4phh
TlpIJm9d7wcUjvZt/qs4NM0RUNMICTPsDKqtij65JfaR4b1ym1VRvLteiOiZUTS8
UCiFgJkz0FPW1sgd/waZ3aF6xnxrDlHvWbHzq3ZQCIaRoxQT/eadHOTftqXSR1nu
ztAthvIl2wNUN8GESrfZNIc1vhQer8jHn3gX6I0nN3gUc/YQTlh6LNsNH7ABu1XC
SLbJwv+rh40BsDSCbbZTXjRqzQTeBvFcmEcsQ/1upzg4TDkZbKdexNm7ctcvJvs9
Zphr37mG6b73Ox3nypDJZkU3Il/640wJaQOm3yoax6gs/w0/02EKrGTNq3K7WzXR
jFpwjUNh7CsT+4A9ODea3uvjkmBIbViUPLjgVUeMtpIPMB9lLUM/zC67tgF+i1cN
zUiE1Hd+UX5sNIAMmLXIUP9e30EbgUJR9MncFHr39uRYcJmznA+/s3yHuOCj6vlj
2gbCaUK8vbrtjydyumss+EWrFmTzRMxvqgJSjb4vTxW1/T24cWQ8YU9frt4ORarm
iLduzf5odG3utvLQAvD/xwIc6WQgqmkmpqHeJqRT7B4XuvaQo8Y2dw+fh6N9WZaR
9l2+aT6N9X93JymQWpgQW0kfpFzz29dvXGqXFzhsMs4P7crXp86EJ7xbK+4mTvMP
gwu+GB6Gkyx21q/P7Y5F2iCGoyE8wfgu64X0m83lmobVYPu8qoVedK30zoUvfUFj
K4NCd7o7NN7JKw1WfAAuWbkputfgZnVfxBx+ZVvmomMO/sMLgGfnjz7AXvHRCW5m
ipnOA70visvgPmlR+2Fpt9CUWaLUJKuNakTVehnxpFagwc5tD6L9Ao8wdYw6Nbhn
CAOUWvUAFXb0VzDGCRUGLOjHkYtekZuVPi3CwdtY4+B9Gtav2YpsUYiJN7/iwEZb
ZGBY8CyjPciYDAAR9TlKqmWxNeeuR3DTUC/Zno1pGhrIqPCiQ5t7Zre/EeZWlApF
2q1Lo85S6LnVqwXJ/phttoX5WvHkl2e1Tk4aJgE8o8Ea3c2VeyNVeUBg1LfVhr6X
/xUZiClp+rF5g49mf118GzvAcltuzZVnsi595rIOKkTjpmHB5uD4DHZi9wKxqR/M
OR5VgTh+NiDQzlj+Kvv/dWzbb9nN1WeNHPCpqO8BFjRA1K/ZZZBgf9xT7Caub8BP
1Fa9YZlA3+69IbYwiwMrWE3CiSan0yGkydz4DiCgB48ev/Z9S5EcB4TocuuENr2f
57RGDZeH4kmcSxGAislty/dWuXhkaA+g5ICrPuFttb4coteWjb+3uMVNAqI/ETR0
EBzPOHDQUSQ/EECev9RK8fX6YlXiXJwgR7gfhcNpG6QXUdajZd2VbxgkAdDECIu5
DeNFKd8v8rzH7H1J6Ypftj8IdMgxP9836gK6nknEWCRDZjY7l4Qr8tHR/VtFdeQk
k+BLFk47yVzcOkQVVMqx80tsx2HXlffZy7Pf9ezbm1BpAWl5W1zw9MhFgBwqLoTv
GIXO+tE94LuEx65F1bXGT9P5B/qK3FZsezyTAkPOkEYW6EUWDIW5LsgoLfVz2gNb
d/hBEJXc3+oFZMw0/8UlomfkSiry+wKhKhMONIkaPo6Y7Wy1s0/kESIkE1s2uXrL
YgkBLP3yWaBwEKlrd3/Y3+1QHXIdK8hT2NaxqiIjrjkM0+bRjG0/fIqUzFMTaTD4
XjtPy9ZuijJqv4AY0JlRQOncizgEgvyAC7uLSWIRFR8qj3TmQIU9nrMcUWvTc5fl
CYu4cwWRnglzGq6PakSw8YtBFaqMSPMmBV50Sig18aDednUBgyXBaKTyPpTjEcYL
noPI2MH9fvCAaOC1ftfdIm2HXVggQxhPOlFCMkGnlMBjsjNSRnDk+WH6BYkkG0on
aQD+wqNibVwc26jEhs4p39NvpFyZa/jJfNw36/rVGW7jxAvfmAvoxSfgmTRwMWoI
QC84gkEpqwWmLjjNKhUvNVAkETaJJO90oxtNtpgpYqXpjG/aL8o73fozvORtCFlI
oMBSHnZJpbRRTXICnz2maaSATBchVepDLQJ/W7L8gixTuPu1bKzfaApzU2fOumND
XM1SepiDhttYe1rA5Nj2SyjoXQCA+7aMpYCPFAycH0mDBrip2//pvfchXTjMHsR/
Dy0m0+tLv4bliYkcCIAPFrPRQ/NfIOIU4iIMbNIBc96uq7BJKBjuIjNvgOTFlyoT
7Swdx8we9UyxJmH9KhaMepCqJdWmN9Rofa7uh3HWLk7fL979iuRroLTqVDO8qzi3
OiWkeh+ONr5oljppwjGm2TcVP5qBFu1Ru5cbphVv/GOTnL1vs9JhoQVNbn5WhAbW
SJ6tVJXB/OsAQ3VCn/rllyq6uwehAu/H9Z+Fwn9DxR+4yPvrKh5GjLnCT8xckElC
MMNZsxXqDRhg/Z1448dPLRvOPjKPVddaTQnou+R5t7BePz1L44vkf0f9kczh/hS4
Yh9F18ubnWgZ393SgoXC0aeYxbSmca6qF8pfgdHT/P9NFjUido++jsqWEbEujl7g
7DUIxsrKb0ufm6ZdKKIhI0Sxn/WUzw23+gWxTgDRH/VZdQIchRhG0yYMliI/MkmN
cjCtEahl7lHsajAxzWf/qfPTbZppmCF8kC+wwYYwbcIs9z8lAE6xnKhxv73geUkf
mZC3aDLS83zaHE31Aaezn0Ov9IidNk1t1VFBmibjLQOQFQ3f5SYIlTEJZjhBKHyU
wApoeF2Ri9uOVSlZtlqKQB7r51Al5hUAfKWL0DmXk9XPtvbCjxDOPa4yvpsZit0u
kR2junYZncSnFIHKmYcdgW0oD/jDOPjGYv6zXzkyNkLUYO+8crr7DUy6zPfZbLK1
LTzsePdyVjhCVZ6Cq28dI55gIVWuATl+IRND708NOOOwkYCETzs7IvwCGEZ+L7h2
mlzhZILPmEPD4G2wRWmUgec2iM8aGNHvbdMpHOqgMSrGyev/Fp1BKdELK7db2PU2
44YyzgpKZL4gCUbjgUZdDsOwOSx7NBF7w4o+aygs78nlW1n1Lbl+gaGWJ63Ilq2N
Ia6TLqmZyAm3UcB6nv//5cRH2S64Ltx/wmPelRmtfJvauhfmh2KPzNcoDgRQlVNc
d47LMvwS1ywWbn8z2MzH8tvYiaL3WNv8eG5RmLwU5vPPrEylYmXGvcgbnOe8UiJO
ANCwe6v9i5Fv1gXEWi/8PldAb+fvOLQqh4SpNwcp/eW1ahg2E33/wPbsPbwS0fM1
q0FzX74HANgAN+2GYWxvg3AzRViGuQngHtv2oeTc6KkWCGQICo/8VGNDrspjmYOX
Cp82fl+Gg4syf/ReQp8UXlpMZOe4q2VieeYtj74GYAyO68YTv9aVhPC5FezKvpRK
kUETjCDNF0iN83vGWe9wsTHXmITsKeJQyL/ZEDYNFHXRM2c5RlNGX+vP0NT5ApyG
ve5kBFuB8NzxzGgnDECk4kntR4zIyUbKn9ceyT1owS3OsUKC9aK58qZ/X+x8am0v
JiwG5oKFHjws9T9eQq9M5f57f5yj926wXMz5MARkMhT9GC54gPWcgnteQDtjs24O
xGylnsgdvszuGsUoPMPURMKVL0hFSOaADXBPnJPe4nLUtTSXaEtJHcGuGu6Wmxlr
QcvgdEr1D7I3k4h0dpFXL7en2JRne2RXhWWGHbEU3sHrj2Ec/Bv15ZG9/6JACQD7
LiH67ggOSDCjfWMHwRKJI0Qw++EZwmozc/dLlt2EFpfqYf0BzM7nepE3VrssQNCK
scpqf+cpTnwCOgqiKNZFi71yi7o10TB0RvHGZE83NjMHYKuMIg1T165/Yz7V+bv6
/5ZWVvaD/Sanc8Zgjj+F+Is5Hdg5kOlpYtfoGwvTWUI1UgtF69aY/St1ObF0CmUP
WUSEYQtf5uSH5v2oYtR0Lcwu03AhiL2aAv6QVxnQA3tXwmIrWeLIZrdwmhh+30+y
Ak9uJLdk4vCU5bHKrpjKinG/sneymb3K97pNRE6DcsQp7V6VFdjtPaRuX7ktqWVU
Cun+MeaqdfnpyUl8odwsA0Fi0ktVzziXD79vJH1sVgjPoLfSzvjJuczFDnx94r31
CIyDBFE7z2nQD16WHnx3JBgXNmd+0O9eVy0skiCj0VhSN9F9utgxCEhl7ai4zp0v
cuYs+LFRn9NnXGtw5v71pjLog4wrZtFwdRKLfpsz/UM9mpsEoSxdG7Jg983UxFUl
M+pTOtpDPM35RE16z2tjh2D6beV2tBo+q3NR48Ylp5qWGXHJASx1sM0Pa+XjG3BB
yAqovWx8I+0UzlyAq3on2YPdkNle2uhIC3frsYJ1Rmfdk/24znyawuKvDCD5ee3g
IF91hvK87DJqq9L1cjJd+kBwGa1l2XyYbPN/W+VQLqPUggi7KRrwznRERptR0V0e
m1MXuhDcA/MAAA2Ir3R28XzZYC58+5lPkhJPs6QXVf4gGi9fSmJ8TQ/COS4v13EH
kYnVmkohL079DILTmTCEiqYQVuWfoNa/3Um/vUstiRD0bUwU5UUWqcQhdzOZhDWl
lpKyPTB2Lzxr4Q7KA38s65xF60nDvNEmLFIzRMLH4aW8mNrzcVojQ2BEqj8nTFSu
t1WAthYc/Sdt8UWvqEp8g23TGtPBMOwG9UsUNDLSeOyPyK2S4aRobQ5tMuN35ZCm
22CX3rA1GqM0vmHWF0y0ud2vmEGbkIZHrKCPs2N+gSlDf+PS3lYVS746Iah6Xq4Z
X4PJamA9pwDxfrcB/sV9/8paYgKhZJ9R/bgsFs/g1D5rGl0rfBFoqOj2xxMuKMjI
rm7vnVqCqcZYiddkVAW7S/mGdFgUHBq+5EqLRdc9R351f88/NLXNwPgWIyzkYP92
yP5/n6P9d55r0y3e2XlKcgAwoSSGuU8EJ1V1VoCfuDHHkEr/dyGx5J6+kE0DURTw
SRKwA4ep78uBReqknYH2odUubRb/p6asTqWvvMubCwjN0bZrN1jjsJQW2Fqc2cDy
uDXDOS72wHmZRjREA26+CHkGD5SfkMkod3ZcaOLCV22RtTAJsWO7yJrBH89jHnE2
nYwXGBLLEyoFAqQbHVcEBiH1ls+QNmT2dg+RZCsRsd4gU0CFvcBo/q9w6/31PVnY
7JhoCV3I5BppBhYQ3G5GmrJAWxMzMLxVha5sv8Kny0w/0ytx8/ThGKhg2QfKUau+
X61COZohbrtfiZUim3nEkIEAD/285TqF8CdEHU7SEW1IaoZmjOS7Wwf12TXyx+8n
cFM8yeaDwCpCV5nO9iUzw8ihAXM33ytmyOCRknWj8Xzo9qyb2auMcDpqboAfqtJP
DoRRwAawryFRJmGxWwrvGaWQTNOTaMgW2otWDbEOuZWl900wpxDc0Nj0eaATAAQc
5OQaMDAELXB5+CXrZqivWuMhmCD8D3b9GYhjfnoQrFE45Y8TaxV2Ae9SH0CTPUJ9
7obfF/5LvN5bSo7RZ90ftMNElzNsaxs/eIUIqjzA+q4bYbL/w2E4BpaTpHZrj3sH
plXoyPlW8uqUwN3H/SBOK/pyqQ5AE+XZsh5E83NK87oYagS0eh5bTgZ3X/C/Io8g
bicUgl0IJvWiPdxHk0l2BF+pjmwyDf5hxIUPsUl8xlL3xrxfV1MaP/QNIMG1pj4h
BkhXjWh+QNncpYUhCjJYgRPFXilU3y1c9ME7GYX91xiMVsE1ZC7rnPm5MNO9jLE8
k+2Ooh2VdqfipaspZyuobnWbGS3jsZsU9NyleWDiW0L3G/tchgkQhve782z/c1/1
t/nvH97PeT3BQUUQ3ijQCicqXa6FiVncbRjGWKiyyHVYosb6DEpm7HuHDw+IsvOp
V833Kbadl2tSmS7gPAJigD09/wkT6oLMKMKPCkx1qi/5nvfArL4Z3Mou1IxvWkr2
3ZkhNUyW0p2kJirJSHdoPnx/Hgi/jSSGAAuNL+201sP1kRELUxOV6IVrAE+r045F
GgkbWtolBpvfMqaWE8XTGQXszaQqSEq/WDZ9rvraRzT1oWxfnjwr4xA+wV3PMcXG
clzzwAHwjxBnGDJ9WKTJSqdiXraOvlLBVz0EFsNwPSueMlPqV1tfsNgS9BQAmH0q
UPAtvOzoIhxyTacJxPNQpW4ZyZD91lSDnu435wsB52S4c7pahwYVhTQz+RKfQhGt
rf+q1SJ0TCSEEuaMc5yk11w6nThXokedHREStB3JDdcyLiMAmbJX6emBnOFZf5yk
EHxczqBNB8ONAtZO7deLqpeRymyIB9rMcJ3FAzetoEanCkyCJ2A+T6KlWbHk3+MU
WP+W5N8uFYFQFRJDE1NSetJoN8HeQ2yaI8lKp3bzECL1ddrY34jUwSAQcKuLRXWI
GVTRXLGjZH74+MeB6NQIsVwAW/Ca3SqoqhN2nQGJ0Xo68DtOu0W05A8TPQx1To/A
4W3wJ7DJfq1Bk1jjfDNvwcpclAVenHNCxFtHmM1Ekd2jYf/ffdxbmMM/sP3kTTbx
vuQSc2vPrOMUHL+WcxA0dP6AGZByQikqW55PNjhznvOOTEayaZ5Ol2hlphpeejQ0
9YjIHvs4Qf9ai/yfZbOzBGuqC2r8LLphQonftZLQMZ0FZsmKtn+qYQA0kNhT9ZRp
pxLyHdJYyNx9IgFQvPPVHSDfMnFdAcRWNmDiDv3XNMb+AQaivqTjPL9tPLnY1KJv
2rUQzgXXoCsOLnHd6cOIKZW80rypafqYbSTBs9WBOTyQmQOl+1oV/6y4sBN2DAGd
TUd5mcRSKwvwlxZrzxwfaK6G2BkdobmmCGY8SCpEVjKY+zl8xjg6cFmrD42ekfvb
d7B79+zFqwLUlpY3WfVQ1UiBKHycCvuMJh31C3BNctYu15JBTo7G/99hY67csnI8
xcWeJh8vdG2fOkA3HAxBwnHPBs0uHn0jkJqtXP3G4YIZC2HjFt55WHKSCbmNyY8x
gCngOSHaH4eZ2AoLLukQQrf4j499MvscDoSdFA1Cpy247860q8vxwKvsscgVL88Z
rq1UjIa6nIeqarQ+WADcO7y3dUlObFTYNsTHt4KAIElpWDY1JQBV/hRAxy2Utnbj
8f3oRf4W71+iejEBanVtB3o4X3u7LDBM9sHZ26VnUYLHQSiZMmVfhtGWd1cvpD4n
3bAWr7yaBkQ+Nl7EtfpesehwrfRYGqjapBWDFWKxFNsPWtAZ2QT2MZNmOiQ3c4CH
+6lLcHD3ujk9eA6xdeVCa3C/giUJ6oB3ABCkH3/BQ16Ocw+PwDkai7lBok/sqdx6
82eluMxZGEr5Sq1ZE3+kC4hf+YI64kEAxjh3CQcaHfXxj5H96HlB+zS+dgBt/Dd6
Xg6xpfxPvh6+mBiWsaLH0jcWzXRxGqgbga+j2ghG/JgcI8whDclzRqVZwNOxweo0
GF8Oz3J5vhrfhdnKL3c4otuqgnRUVqB6g2dKSQ7YvYjIG+u8jPyf6WvOAnMIJmrQ
Vdb56C2FIeppcad5ciybYYq9TlHyTGLVGjNEkl2HiXT2gF3qwaYtF0IE3Xb4UoO3
gUF63ga4EzcBdUSk91RcOR++sYLEjGBpKPH/O2urLzytWRkzyfpf+j4rxpDI3lDw
1fmBClbb1+9lfyjv7W3pD/S1m1ZdBWd9mES6LR0Il9YKYqTC+Kxvk6lBSQZU8zuE
EE1JB8ZOmev3lEilkteLoKxDUHNztMOM8bHPuYTc4ZpnNvXCHWQyQwgLL6PmToQ2
jYParhTKKFKhFST6h4C/bl4k0xTkZrPr7pe1U+HEI24cAMfoPic4hwLROlKd2HCp
VXCdZMZHdj4oy3LT+pX1tVVPuTA/W3GRAEUB5QHTN2rhfFw1RXhvvIhokuVzVo3p
MR7YbIfRuZe5jEb4Xr1k2Rk+Q/N7+oa6jn06n/MNTvBS5q7mrbgDsRJKVa0p+/CC
Qn5cFLqU5aiqjksmx+i/jjPekHPPC0jb0Or1eKBp3HQxZVIU5spX+7YRQoKZhJY0
zNkWhxpS3MTCwmSoeENRvqDX1raR925GiMqHuaoXs67WSXC15L7y/iaGq905rJjx
Fnlf0NQswBDVn26FsxCaPGcElljy5VnhzE8Ub5awkqGORiHQOX7hHTZ+ct18QI/6
HmHp2K0EYmUVZXOYnCaCuTYEdmf9uSxE3k6OtHnYe6DGHYA2ZF1onF/uVjohs4IP
RRdTJ7+L6U+AKp6/2SzWYV55knXcpcOZfFjlPUuART/m3IwHYM8HCpeLQDQlgObS
3zmqX67QKrbKpg9xxPaEyUeY/Pz/Xt5IdscE9aBdUPXmSQ7ocMfI5Vfc6nafhWSd
NCGLgDaMelQKD2Q9toFK0R7Ku4ojVMU/9aYeST4cayM94DDAx1i+wOy/Cv7wEv2L
PiMNBQ9hLaqxKb/3QQ0vzLo7jXMvZA2Bd3vcJVh+2Nv8WKTIpS37UiQjCfFb80Pq
wa44wuSo1AXGEy9EOqI9MMRNGyGphvUI4CeueHqmAM//p0fqvACo9YMNNkcuMtfw
jTkyTssLToq/EzgZtI5ypFn4csUiunWc6qPbLaIpc/R+LmXjea5V+0bMIIts7/me
gTbG74Jjb/6Fg9s7GnMiLXfn4dkAz2+DMBIRyifqqWZQhgmsXncAVLZaqILg1Fn7
98BTBYpS2QPZaEJF6cF3xxlU+LcnC8VCons0nq1Etw8iceLFTOSicxWtltiXQvuu
9r29DHVM6E2xSb8cNC08XDes8Y7604nTWV4/rc2IkKpBIIlCXNoCYYAypZzaR36y
PZ6gDXbZ6Ovos7EYhXI7qgRpUDDnuGpztStM9JWq6EqXn/Rq0fC/lOaI9cGUWJNr
tHmMcavQ+dp76/x5Wpek+FCnswqIvxQR7Oyu2a5kzDdiwScmkoAeKFLIox2iDe+7
hmj+mKZtqTpYVFV9n1hNDd8uQ6SZj3uPr0IbTTfZKEiAD3Wj38Lqdg+XW17pT3o0
InB8s41bUhF+F+UMO8mNLghEee7QVjwvz2zTR7N4YFUKX31s7HMlDeTn0JdCcDNC
3X9/xrPs3KxcTSgczoECRFyt9ZJoXMbhW3HLNFqvgHTYioFgEh7ivkkI215gilBx
rxAob2h3AmZGg4mZ2M9j3cM9d16RkawWxRmLNcHJr9cvdVguzy3cjyuyxLJsw743
y6MbtJtqqWRqXCygCUL+HJWikmBEWz61305hcxbH8lKVl4ME8+8Go4xtRWVppvS0
U+nXqos+j06yiQshcyykmkQn7kx5rYs06BI6yTO6AjCruSS+kp4kMbLREddwyvNu
DLbtgLVocSAoeQTnquLW/W5lsko+eqNQZNh2hAd393hhxevXALLTFHfbIjyjG64C
8kw/+pmXKA2m2SFGHsRleKhhn0oGv/IHMqgssN8rWnqq8J5S8e4vA95yiBgVcY+f
DOiktJ6QAP4qWP4Bgw+hnAP51vlExpq6dPCBOUgr8gEldBGGbZTwa478PYLwMNKK
DBo1XYdGxkPRhe+F3zs3oobTcO69OP0JvYr1AHrU9hQ6MHdkw6wZZw6U0w2S54kL
WysGj6A5MgIdd184fkk9Ia+/cMnTX1j+BdjA8O5uSOnN7N9o9xer89F7wcPkB/IW
wlQKcpcoVTbIFi+2aWuG6PvwjnmgQtsfktMDqpkS/S0F2FU7jIBAr/BgP3ehykvC
WvaNqi/9t+prgZw8n56JN4XnddLNTd7Jvtjr3UWRqjbR0o7TjNiht5oZb6Q1rNHx
JzOMSA4UDsk3Xx/BA/EOgOkzIEFPTu79AiFv5CHGRiCft94ffUEx9FGj4a23Iyr0
9ZzLH1xu09Vl7EeprE5rZlHQakhh1QBFjHu3DV/WYUDGQ3VbcxO041jWke0rJaKj
lYI/xFg7ohn7PjR9s2lTBgkPUk0dAREZqLhT0BJxazKr0REKHmP5Ddibn5IjVyM7
w3PTjCzeY5HuRrSCIxyF2rnc4FhnR0Uk6iK7SBhd21T5/2SJruSMWqhzWY4dwuSE
JrDs9+CDAnncMlo3Dhp7uclGmTIRw27oFhUNgr/M71GejaFkiU1zx8SMcsbqRhr5
C4LYHA8oTGANqYgMCKNlLwvURwg7U6oGCXzif4K2RMfqdRsZDZVku//fGU74KtUi
62qjEPZDy5iZ+YkaIQMVA5PhRYqGninNB7COs1DccWXG/0j0dPAbQ4NuMWzJat6+
7EtenOZcainFHftHtUgNmq+NhUtMbsSw0DAHTPdlUvQ0RhruCne707KfZ2CXJFVS
EE2uUa3I/PWM9EgUH5I0de1I+m36sOe9ylO+fL1h5lpsc69bSXURSNUDIox+ed02
N3qdUFfN1unHVrkxMp4zmgLQNik7wQu+EFlFe1m4Rmrqp/aMpvjdNwPPPXoC2ElB
eTS0U/9SLhKdQu1+evrMyXZxoB2vVLJ8ihFasmz1Puvmt/rPB1nYVXDQG+BX2Evz
tWf8268secsktnukIjXk+cVz9Z8nKoS8I8xFNKRPFldzNo48aLZd4e5gGth65RUJ
x7DXbA5yvafFtlJA6WDuhfpBmSu6hmVc+BpZsyRkvaLgjwDx+GH8m2LKfn7Kpols
kh3hvt20fDG/u1yK4QtosGa3f6EvdCZkcr5VnQf/tlnFPAGkclfRnD8SxVSFfLvF
j3mRwCHuw3pAtSUDy580EaxoEoOkWryNMcq5qYdVb4e/OQ/7fqXcfo06+zBdXvAh
229M7o+b64oGbj3oKsxAlUAM1to01RHolO5DTUciUSuJd/bcyOHBSqAR6zAwj84B
XWNI0c/5mGA2iPQ6C2yEK/KaU3dzR90CjzZPU6aN5CaQ9BGjdOeWALff88+Dvj2Z
BNdtJOQ7KaC3Qp5aki9Jd3WtAfcQt5TaFvyd5S9NHcQO4SvuGplGpyYxvw76CMep
i4P7EEveGSbshxivRnkBYNYF04WtZutJGsv56JOrM4TjXp0pijpyOxz2YXDUWRa2
03me7ooVy/jQF8om1eUX7G23H4C0gmcGpNDrXDZNjVvmcG5baLxH8NIzRGetnohX
Y72iJGglP6qNIDuGAUWy196qlFa91WVg+BRi53Qh2S0NEcv5mc82rlW9X93CMi/S
CXpmP3VbiumhtknqJnUfX1gWUPoBwotF0vs1BiWGCCQFIQjGaYWqsKnsEgmk4FIw
pKGO6r3OQp80kG4z3W2SgEmcDUGebchDSYbj2UhPvFXEPxNzSBKtbhsiathwMPgg
UgUrl42HCnW7gON1Fafuy4cJGxGer3Tab6jYUn0LMNEUo7U8DpfQofgEwvBqxAAu
4kXv7Bipf02EbHu4DCBQl7QaeRIz0Tj8h8aD0Rus51WF6gbhvRyaEa/DaMywg32U
9MA+0qmQCoa8DMEEUZPkJX4GtcGD4YEds4IBt1p9I2cK7PRNXojxeDBZX7XSWG99
nsOsM4WSpQzbuPPM+FG7SjpQAZdvzaIb7fId9FWzretIUbNY+KCteZxphbX8Jmc5
TUHzBpvUP6mRGbJlAl/ZhHqXf/M0Oj0QEQeJ2wBuJJNkaoBcU1/gMihS7YFI3czb
uEt20cNyZHku6+y9jHENYrJhNp2SCpUGV3KXbx6r0JLoRkFxJGwbowDRZgIpMmT6
O7Ym+a1BGR9tJkDnXAz9NPCDkRgUyexX9CulAwSQYxmV+tDTkWjNBAmPwjpNWnGF
01+UCEDyM7IrdHfQeGfRTQnaf+vgXIfVSRTx8hGWSDBM8080Rku52WJy6MCy4Iwv
OHCMKF7DRcapyJCvXE9SOtzjktBN3Ko+BCd2N/Z3lfi1F+VTlT+ol6L44UaIHm56
eQFXN5lWLVu+uMDtJ1yFHR82hRo0Vw/ePLR2iEvpomcfU/nmVbgXfTYBYb/MUoDP
t8G1e1T/qfa89G6gxnICWzNHEiHDJNRO4nyZJ7/QZu2a7ShEWxVq4GBcCAT/Oqlv
b7c5+GUpKcatCbKd7q9BsD7wzmEErwpNyDQBafr8TQWOzaLqmnCOfoJ0lu3zGyEP
BHqKwajIdHIDpCiWquSiv/JpCrh/xZvOZqs9mo1w/PCyTcP5INOukkMZqlPj7k5p
etLfocyELO3LtnwgLf9BU9rhJIVHYJzC2Eez0utBVSvWWVY6c9QXRmdacLBIcm9O
dQnLs2T4JakTwQY8vOzdrIvlqU8MXhmNZE2+hL0QE7NqJ55Edk7J5Il8pmje/Zaw
SXA9PlkJcnWhoBwJO+bRfqHnuIUcKIpfvJuBezzG1fprlqPe2Sm5b8Ze4n0dUbyE
4O+uqhTwIcHNIJ/xm4DNfdQlx7clrGhSXZHObgrzYDp4Zf3yfH+rjDv3Twva4C20
IQEPOpKMFIDbZX/m14SHbxpoGuAIS25yMO1vyceYqZFnOn1wGqUb6TxoOuEnF8Zg
83Mfm+Mue+utk9+vmyuklBRYK5ccprc70F+2/qyeHNPoT5rlkcBN9My0hnFwLKxU
hhc4DCyEoSpk4VFCP/9AcwY1vUkG1jx0VRUzCx2iw6/gNpVfCT0BPvBvjNUFFmRw
vShovpWH4g+KTntNGKSUdX91gRTpNLatXgub59GGER/MGYwVkIohB0KKe2PQf8F8
3B0mT0GQEq2CudBO2ALN3PZb2rH7UFvVB1i739qaYv+vQ7smM2+Lp3h9lGMnpy0y
8OyT2i1JA8NrqDlf19ea1xw6LkyU1mTXbDvjxpvROHc/vtYkMYxKyp+CoyJ1ywCI
UtnJlqa2gJgfh60c7Ohq76ekbxYoLuHsbfe1JuGG2ziZMC6LxW06EyicIll4TL9k
naWnvxeNceVJhH+DGNgmFJmD/n27NpgEsw+/jn2DmFCUvctnK26KwPP0nGWuaZpJ
CpBBgl2GMWDOH4s2Rsun+do5S5/DU68fRTJN9dHEXe1q3jY8HmMYQTx6IGiLX0Py
04VinU76j34jg1ij6XFrybii36IaqsGq5x6/b5kRMDqhkEAXTLtP2ftCFZ26MVMb
aKmmFu438Zd0sNF098/Lp7uHRffxsFVtNdMZly2Gs10amLmu1HI8Uta31mpslKI8
egeq+yS0cYJ9BdE7k5vEiRCjNM53en3sIwWPqeYYVcTuI2mRaRLJm/nhhw7jpFat
PDu6DhiS40wpn2LkVsV6N/tzTt7/bO40p8oh5I7DBrNQiLrAqkkiUF70u2B21YLq
68jmkudFg9XAcxFyzIaP7zmqrCoXqE4BD3kPfU3SLuJ3oxkJg9JuncSB0HoqAShC
QzZQ1dQDkfhWoU+4t1U3eVfhQlwBxgrAqbIuQheZxyksqgL7tAYbVrjYLK/i4nOq
VMSOgGYHXhY1r0zIzSs49NGvnI0zFk2uW+9qrbd9ZyWfK1zDduV1RnY2gHwRzhnz
NxL7uOsKRCUaKYu/9Pn+ZFE7c1uYGLXz/Lrm80cwnN9ERJtQTXykOeBCHqytp6ft
mBts5x4q4pshRf9KfK+0LSCHN8a1l9XWZsrW7CE7ZaedCIOjCqUM4JM9pDPg0eX6
k2VpP9i9Au6mdySHDREzedyCgsNFlYcgY0Mwz25M0PODlhA73jpImftuNdXB8cs/
wVt/Iw/NnboM7xobZVAsVA8ucFoyRoxliUHm5PMKylWPqgS2qgs35yEE6YWeKnbu
ZHRJNiDAw7WEo2h49I/rcRGDiimliP26ND04E+NrJf94pPeZfxLypS+zgQfUoCbR
g1X/PlsPrqcVilutDS7rb/Ez+qnHyOflSCFzLyw9s14qZzKoEhQtBRQ7bSMV9Lvo
UVNpwZqK450s+E3J1bgNrz8+hzBrDckCum+Q3FHixXYsKF6nuWqQjAGO+WvEcUuE
m4/9yXSA2+K3xSd7Vo0rjIjIPPbxGAdLeFIST6QxcoEzjePNaEaAgmp6EVnLopRS
8M/1daI+DcPqO2S33+GLzQindY3aeK2/lI5aQOU3ncHmHZryHxou74zS/vkIGOGT
SwO8IygX5h2wNkKxzbjxfFALLSMIGBx823TgopjksbrLRgIS/Vqc1EKRijKjFhMC
pzn74RQw4X/Ut2yKwOAL6ySXh1/IBjXCY6GlojufrNDDnamEpwmRySPWGVpJw0Xu
CxJGmTNqipVW7DDD3mui64lapYDy0bDq3ibzK1Z83/xZFPt+zGIOWH2RfZLQINUX
w0QZw2iNJLU3YLwMv+oCsfSfdu8mOGjIdG3n8/YApdRAY3nMxgEkHO46OQT7Rx71
oDklQ3M1v6OE9XMnOQavS4iXk1fBDeFx6rVL35lIIyGX0R/iEoI64c126MjcApIx
rOMh+DfIj3KC0oRdE+saTHsd2THlnnPhFMIMNCWRcAjbjvVHMsvJEllyJmZeeH3O
pJt6gscvJL0x/Izs9KHqS9qXZcakp9WiYoS57nLxyF3tLCEJTubYtcz9hX9ediRy
FENfUZVIaww0BnsDhEIx9KGSCKElLRs6mfsOOu5U3xYn0Rkan7hg92Rr4sOVV5tw
HamBXuMtzxkJ9ccwqjC1jGMsQRR3H+bp6eDPkHRuYKYTwmp+21vQcN4FaLk7PuIH
1UA1lcLzrm6si6u5sRi/HkViZopXAt6kwW5au0zwU9Dnaz1Wyqd8OgcQ7HBsgjhb
S9TwPlH43DTsoCZsrAsTOIC4YXtQ559MWfTfAyGh/fRutZKqaBHNPZaJxFXRK5P/
mzmxPSPL0T9roxNiu98xo0tis4hovPJS6+QMIxoeZF4AU6a8rkqBmDbs3vtuGEpd
xf68zjee98nq/nA9ZES7lSmjAyQDF+2IgV3zScJwa4Rm+bkhu+N5iqIro7NDwSrT
E7AOtiT9dy47HOwTV89ikXMhafmkQfL2VrrX+xa7lyUV2oPHep0pFvHlZWyGDw1o
1NoLzfKQyOKdci1OtB5wOOxYKQcsJlOg6+hAnfp24hjSR3HHarFoyybcXAjBhNJF
zWmGnGhfD3WKG0DwVcNSjt5QSIs/c6GP1ivsQ+yX5D24efw0CUHIzhkyknhlv2KA
/kcHnWUAJJRDiUObPlD61R+ivLuACL2AGPXJ5dH7Up6WRjiwlDp72Yu8VVeIqYrR
fDtxF96wPU3cE52abQILe8FjtEaP7iqZB2e374cnIGNc2VVfl8ZkoEpK+xnd2uzk
7i25ZesrSdboHtKNDbgoX5ehfLWYohdMvfyOLyhUNwLZ10LcGuK7uosRrpBy1+US
jOVL9xvXkBqTPxY85TtmA3uHr+t6uRk0Kii8L44545HONIn46I6uhP+Q2kMOkH3z
BnIxRK9ZdUkdXuwVB1lxueAlCFuUSABew+6P0dJCNzb5AOmX2tBvdy09u9F8bAy3
tO5DcvEBxguqprheWOxwCAvDjjHstyf5fS0EJ+2j+NpyWRvX6e68f6zaWI+CiD7U
kZBcBJTQMn0R81pyP4o0LlW1uer+sxh1c1mzuQSHZQAnxOC0Nj9JYKMyap0SHS48
jHY10RPdXn3NiaEj6Bg4+JGGqNmhM7RiXN5/25+n1TQHulSANp8GBjPGZeVNsTJ+
+MvUz66bnDTS3YIV97Gxiltcb2AKPtfvqPmnnWd2QlZPC4/to8Hb07WzT50jmQ3E
TXtBTXL1GD/BXwz0wvhYjwF11uwxdjB/I/4UwLG2aMTBsUVDc5bG5u9kS0jjgm1P
3bOnqk97BWjjpoJl5KyCC/lFTd+spPqbMdZ8zNex7v2SdyRttYy4SXMy3Lnxtn2F
SW8PrO46K/lN9ODOiCfrCGMY5xrbakH6YIPFhgHVos9LvTYaDfZjc3aJ9e53sCJw
1E6A7xhhJ94Rer1QkkABEwXm305L/7zPTRD5wVf9fcidndVUOawJGr2ZYyEtAdwN
tp5ap+UK1td/7CGOlP/WRAgWI3LXpt8oe5NIG91KochdmLrPqPLldLiooV2V1A/a
5kRvqiwwUGpQbcgVahg2PfZ1eqOJEs+wCu3csOwKLLlFb4nwTeQ19t53ixAoCB/a
mutBj0bvB9tMp2Y8NKIPTGPafL3X1H2z1fO5oYQyR8CeU6vgCW96ZJCXXmrYLXqE
gWY0Evmdi9/xjAxsn3+I5QD3ExtvgClnSV2SOaADn+nd6zyAtZSGpi/pQgHx5TSj
TPbx7PC4T0cx9rG6eTC6yJrQox0ls2C6DBjuKIzTMroJPXLyozJWI/kmjGvmzCEQ
IzxJiOQIGohBRKZO6QvLHCjuk0EV85290ijR6c5bJjKinw5YIV31iM4sphRovnaP
o0c6aNLM6sl0auN7phexmhSAdhEu7OnKPNQ6gKTFOkmEuQhHKB9wbGZUW5PMTrzG
gNyQxdHhyZhdSAzcxd06lBILqPSa8qGeH/Md7iecsSjZJNI+iRqNtEDvCKYTJh2m
oN9moWomdaCaal/Sy0DjzkmRRIHgAbngwm41ZCDKhedvkLs/5lj+rj4Xh5nweDXR
mr43vPcpvRtfcomhbt9O3tee9TKxb3hIzYkP0J5ivIhGK1RLVwTuIlrCNTXr4UnY
6g6LD7FsscT2HlKAHDYtDlhgMQjyJTY3QyABnLni2dRASb4bjPYjw35ccxK3uDjh
d4vED65VotWe68eVVO8D2y58/5Ap7MiCN1lExu5KL3H8jEjy6vGNet+xnIAfk4Ig
RkPQxH+lm9vbznVX80i3p9oyrd2KABWWteqPa9i/mXrCdLd40xBpGffC7UI3QkKz
Ew0rHZBNkRkRjSY7eu00ngURO2qO4N2lGBrnV2oT9o4ztJNn5rUFJfLNmqguIfyQ
YdVBaFuLnbZ7padYYzQqu1J7B+ANMQ+A60vCAxMs+/GbWOgdlkvxsezmBiHHZ6Up
HRbNzYecUzTaAr1U754sd9fJhA+MgMwJWk+zT+SqfsXVgf64gFFbXBV6I+dAPKXP
QhOX4ljL7HWoem2bUXFpaL5toxWSFyIvXrHmLVgPqAu+4xXKZtb5NST/idDiv0OF
7jNHrM01YkzypKCOOkLNTDRElOuvE2WbTnmZKcwKc57Cy83y7bFHI1QjTqguTXHB
Y+xwnv/cLTbOA1gNPvWGrYDHfQELFBYlZ8/sLhU5PnFBUXelqc9MI33BymHo+HkM
BhRmvl29UOgZ9czaEPq802xFO8UWe3V9MEMqN0D3Q0ksuvcAB9tT39tgefpsSLRf
MrS76ke7zMrQcc6BzvP/sX4+Dz8xQcikRVY6CUowSusVSAS7t7/cFRmaqnKU6UVt
UzWiEALOdV3pdyvh6wyJXAjK0aGKKbjUT+D1uLYDy2bWXwVDALbxNs8A0wpzCCwV
cDXmEVkOoSGKOS8Bj63bp8PHjFZ6AN0I8HJu7qy7nX3m2FXgVlg1zRzS9MtDhmRh
HZB2X4emEzYgY70fM2ykNjO/qNBU5wc8aaTkMTt2dSpu5Jp0KQ1R01rtVc8Ew97I
BBHCKRTiucFjdoBIS1hl+1n0FyartywBYwXWiKi2FHNyhAPgJrI7Ro3zLbI/WZH1
d59fzQ3gUW7/yxfWWobjcDf1RKVDLAv0r49if0leUVXin+4dF+m0rCMzL22MwWM8
n40KmMRWR4khVTSrW0qmVq7ckogR81sCBEHAQ/b7uhKQCp0t200Xmr0LIw5/Y78R
q634g0evMhX+uQUrE1tT30Qnn0cnQu3OpHdvv5tk0SDzL2MR+201cfImS4Y0jtHl
MJ7xtb1CXF4FZQgxM9DYKngRM045Ydm8whZ/HXv6q/TpyHxc6q1ARvxi/6RiHS8O
cDohEBPF3XD0NNXtlJ6FXtJ1zMmjwUbgVsqZ42vrWHE5xAG3guLFkxoCtFPygn2v
I0mzTA6QafqkeV1lKoBv8c9f0B7nlGv449rNMq07LCUx+abU/B9KcfEixeDXFF1c
Xt9jF8kh/l4jRieAvCVyoUg40OERhEEsp+IdsriydEnV31GkRVd9V+w7kkLjxsVj
Cq+i+2QK7jhkgyv02i50NYeM0B+SnWbKZSlvH2VtBF4GuYPPze1AD6NBvFc4Xcnx
Tz/OsjmEcXTttYLShyib73uI0eqZRkWxoE75chdBCLr35saGFIjT87OAM6G/US4N
oJXg3LZ1noP481ZvGseT4OKBet/CfWacOe1kFUuJgjOC0i4tmG+dHNKTOpzA88cq
N8VkCqq663arFDpeVz3sCHU2u0Dw0VdQeZAwgJ1OYijwwZ9qc4Gj4rEzTtBCFatj
5L84h5cm7ajuLh9Hq4oLr/uZxEYylvPdS/HA2yFnGzZgS0VpAyR/q3Zj8FoGQyoM
moEEXXXuqkTuFLu8Hoa/vRnfXNqsTy8dp1X2LNumZUGx0D78wakZWHVxuJljRVJh
zxBxC8QHK0N0Eudu6HPvUzEazsuQPYC+cW25QTgXU930pkcZzZxDvTqt5QQTZlzW
VUe5WiPb2PvoAgTaqRwbclZtapv5xtgTYc5a9JBYrPBJNRN55VuBasUFtFCQviQr
qAEZyj90hS++dhhuMevBtAEoS/EffALOIQ2k4mHjo2mC8m0N5HUaSBEtKRuhDTSZ
3gdcD6ERK1mt9lbUoNFmoGs59dfbDNd3OIuHBviPr76D83N1tnsDcLXlaLeRSvXK
wj7B+XTmu06MTjk8/hsy62zMGt63U8+68faiRgtkeyPJARM3i82ORkAaRiNefs+J
ZXTiSZ+CGThHJPcJ2d2Dmk557UcxrdgtOH/JtNpSdP35hpcizo49DcyKqJERW4mQ
J6ya6CpZdCHTLTCYr4ZBVR7sUAeS6BGccE+EtOzOwMNFXRWxtS+xisTtcMddBRPO
GelIU8EuFy4dlDMdYeaOzyDvtny6tIvDxTJNxhxUWaiJ5mZo3B7+XaWy3qM3Fp2L
0YBes9LktSfIxorBSWpuG4P7wWGw5py5lz1THMlCo9GaCUJhkaFL40T5RdUNgNLP
u4L9IW09dO8uVCO1Eul9BZqycTq9VdH3VOKa4rTyklWfwUx48nX1qO/XgVCaBj1H
E2prSY29Tz592VDaKYTPDtgw4bwdeOAePTgVIf5nbo8PCOGePPYXkhJ4I7EwR7oF
iQ9rQBwc3M+8Sj+eiFRIv3vCAfu4pSmdxrFvwRnnOzKr0VL5+yOwF8KH+05dAJmY
1gUtvbWAhPKDlsKoBiupG4STFhMUkRxKHgf6Tv/65wgegAJMQzF5xDPqxAdxC1qb
LJTYML9f+k47p7+6hPa2ByXT9i++ET7fniuZFAbup3NfVL//oWgujYhcsbeHpQYR
OB/Kfaj4lB+pVFtbVCo6Ag7ux1bCjB7lKGVU/g7fG7ZVNglYsTfatVjDwq2L/7sP
vInCJMSYdDLqjj6zaI+iVME5uWA8z/2HIGHAWsTo788i4QNNe6rmH7M06vM+1/yx
0Xz8QqRIw7qNkK/+pxOGawo3vm4bchQ0zjKAyAgnTCBF6/ciSsSXakPFuIqtPWV4
SN4MNvwzsvyj/5jptc/J7OQrvSMjtaFZ0/zUjEUB1v3xur2emfd6Y4mnPWVnb8N6
WAp3G+JzjFkrJXMMpt6VmCSU9xKpgLVBROSPMVwFXhk1Qrh1TZ2Ovb/uk8odFiT2
ePba1e+hu634wHsX/GGR7WzlWmrc92NjrcUfj0xOR3yDHdGdWY7KEwMyFhqpJDp0
NNINLD3gren5JqcinWZF++oA53+YRKyKIzwz3UD8mhX9xIsE9tcNTB8dSDo4YDj+
ZArGOtqc6M7HhB+I07aHUhKNWt+3SB9xkKqoC23uU22SK+TdhlWaH62J5BNVSemr
2LLh99a1VOiaXi/xvxgpuABofuBzRVGeRK9Wb4qwVGnK+gejOYN9BfVFNks0Z7KW
VdOa5Nv9oZaDrOeA/POT6h7VI8cd6JJEFhJWq4G6SFMO3SDkB3UqG7D5lhmJYJow
+XYZEhbmIrVZMwgHkXGmoedF4guUf+JJYSGU4oENc6AP8WJ75/f6B/EjL24UleCu
YaPESbqNbFd98YFTauZVJtZPe92HMVF7JDWCmEnxEQl+JpLv8bsHb8FF1f/eu8vJ
EsqLJUwVnq+Mz4qA7gs19AFYoGVItRFh6kAFrEEq8/QPUCRrRpceTvn9ZNoPMTfg
2nSLic0rEJrpuwsNwlBOMmq2+tHbCACadhDo02IZmO4QIrWbvOakb2IIFwL3S2SV
iV7+XTm+peujc6C+Q0xKRkT2c+lPj399Pgf3Psr8bI6h/1OHauPJCK0hEOgituqM
cfeyMbUi3HaxNiJySDwZYEIesCyFogA/Uqk9B+I+MQTqR/GDWTwkkpNezWWNf7h3
q2yuI9NnQfG5gGdp4Z9/F+KvA/1RDS1ZtEvKC/ESS/V5zWP9fZhVFqRk/U6VRou5
2Alwg7R7Ecpa9AMYYrpmmUxWs/LRsK37g/jcU5QyT+ZTwLUXtC4CR5F3u4WZQTnk
yVMel5wvwG8xX/C3G+XMbEkSufnSDxM5MhT254Gs49mwK/kuVoWYkWsD5f6EG4wN
vVQyp8/aZLwttHcEVDpbTI4acJbKOSWUyZetPXemKHjG+MSrnyrYQenbshCZrw5F
6tzR83C9e3GaZe4gqQwyqNbXi0dtyQw4jHN+kKmJOrKEEjhWpZ+6fHeE7FkDl+H5
LlCHQE2lbfXX4wXdQC//BQAuwbYCD4KqOG4mPcsEN3lmGYvFytzEdVW6sl6bIk+L
DzQ+ubD6naIIySFuAhIGjvaoCHW3qiYw3S9sbxl3ZBw74YrTsE0iq99ntzSNvAZd
fYI54a67df/pHE98XdqYQaIFgHxWvSZ8QPrcDJSzbk6qOpw0RNCB2bBa/Ve4JI3i
+6NCO2m5xy3p/H4cFdWEuCCvKCcr11KyzuWV1oPCSyrF5PCG/sywTez5CGSibrN8
Ik+/nvkr5dNtyoRD+HHCo3Kl+5HZovddW+q7DBoU8ayau3S15t7eN6wmIyI18i8B
93kK8NBcw77hsp0NtsGpug6xuo25c55sxQYhr8wi31Z/hh1uiH27pOUgeOfuiPpR
kl6igTEgTbkQzQ/PYlyB30JRCcZqAPVp8+atKJso1Zz9jsZPS6wwTrY9soKd+Jy4
O+qHU1w5jWjCcKv78Cdr7/tmRZcbn+LIVxiKxfBB0YuAJ/T1faWqBrywtdOv2v29
N6e7908FulzSSu2wSnMnLSzgymtQlKFXlws28Ec9H132tbsvd74q2NW4nWun48Hb
AxIfbtinzcyh3DBJMd+3y89J+T7amDcDkUOjZzxOd4zZr50GnvHwiMSeasyeXfKX
bZlI4wQE0+jq+icwdGjFxFJZ3Ysew7pSD737BdEP0YO0JwFwD6wMKFuAv55Kz6Af
SYxU5jLehbaSwZ58CO8OLEJ6js7u/Ezm5LdwUUI0rak01YHHfXEJMkODGqcVTELk
brucVvEcqYEEcw5ckA8w696sm1tg1tMtS+za/XAYGgRA2ogpHv7g2E5lB8I1BEk0
jHMcyt5JDYbPb9diIFHTVJY7jOSPcqseGYfCpxINztCcpv7628gMfzaOtnqzgeN9
Rw7NlqtY2xAQy4et8swUEYvxdrsivNQlfQZglX7C4CDnsiiP88INi5ksF+lsYWyq
69OtOtqkRQ5JIEbN/Kk9fEqrNphXWm+fkEVeJpU6fbRbF/WXQyEGAi5kiccOdU1K
46m+YGshTqsSZCpE1bNanH5qOyAhrVDdqP4azfHFR3ChdoeuynYfOQjVCvHE2bDV
YXmqnXJVmXcMq4/pJBNLKXsd5sydatjZz9Yt0bBJLcjZJaYZueT32bdYVWKxSddh
oGprgfRxADiN7DiLbtCJiWWSQBivI/EPrDZkO6Wlad0HoYl2TX+sTP9m9a9eoFjY
xoZl665ansibfGyNCX3xucMXo1aEI7mbKX8NuwcgRf3DTHYTYz0xr2JM3vDr5uev
QPqlnfPBd4YcHFC5lo16Nv5/oLT6xpDeT+myEXYH72lY/PB7nQGSTLhPXbxhzomS
mVSB2K6pEil+2v80cjNNnwD0K1b3Pq0PEZsIY3G77J2mPstFtpkhAuRC9qIxU3xn
u/Q8kCTOCqNiwDHnmScYXmp9nm5/tAxmNForiDeBFDCSwMJqn07lOLVFzCLUbFUE
3ypMTOMQgbn5p6ELTsXdqyjnzCKXCiJoKGF4gGZw+L2XKfMUupRNy57LyTgRM5EH
P4ub7ujgRTA70te8iRj3jRDm//jFC7PgSKl+AIW+P8ZF2oRQK0+xeLsDuR7MO0Lt
oE2JIamehIQ0VyD0seuxf4TGDIm06+0TjIyENz7jQcS9DRf48ztQJHW2Rzl7+2+R
eZyRf5X2I58iK4SFBgYOqmELErulS0S7vz0XMT4OWAExCh+uk4IfYphXokQPMJvn
aucIg8V3JxiM8nR4mlzH5yftJw6cr7TiN/01J6SXTd3r9l/M6d2Mr24cCZk6VMH4
JBcUp6CIpgTq/8KtSM8M58TUzJRdZunIbJTrHQ9ckdngOGMlsJlB6WHG1qR+ayJ9
caoZXHH6hSvJGdB443G7OwWI4qFfL1xf9TyZjk+yWkRJqptGyMj86o2wCLwW5nt5
ON02DmcDQtln4+Bmfeqz7++eVNkzEFMRRPXAHTuXz7iNTnVy8j13NPWxfM/CADMt
yIWOCJ+3ERZsMV+A/WL/wZsNTG8XtM2bcJy/XbgHqqeC7QPrOQwo67bvHKarXRMx
Pokd3Yd/826bC/7B3CCIUqSWbWCqbt3n+03Z9UbbkNh98ALr79VsLEu/c+pyvDSd
LgmEGAPTWbtnTvINfsU+gw+LiMFokK6XquR6ge0fpoETcZ33fo1B9x+dEr0t/dYJ
lV+MPuKHcoEM9+PowmkkoeKYmG8Nzxy1WYtZoPjQWZF0xDn9fmUFX8vZDZxf2f3Q
Cri5XRO7UbZlyxtv4QoyUCtb4uAvu+EM1yxJpzmKifh8V0zY8GfAede2MY8qGKK3
bVcY6jDBzO1gn2LpMV8xb4wRiNWJ7RphowoB2Y6gLIXedVX6jOg6NnKEZLFpa6em
YZCQn8Pvzpq5owZSwDV2gTzYAXhjDY95+j7wBbUMFWLFh0XcTI/Xs87MfaBUWkmk
qlrWz9ladLbqhc7LgFwTEm8RaV8Fakd6u7bTcXPHB3BcE8QGa2P4BZdziUokStCd
E81XAzw92YDUTzIkqG8Dt/EUrWsfDWXgEiPQbCxTpJFDON32eeL8/E1XgTn3V6cq
BT5ZKEDAIoDt4hHdWELkXyQClUNy16C+LTRcfldefyjvdrMWTEkxiHsCQrpvT9XH
9oJhjIy4+x6YNz8Hrmk+AtX/+dpczFPTTMOeQDkVUhoFJ7Ha+++fJvvlzr152Bdv
jV7Lo6/XzbLZmWrvefK+2JWkOuV5V1aeULEUvD88txufTaWrwClb718K/ju216D2
tCU6JJ5ejIVrIuLf9Yz1c39IXl4PJZfIdEoGjN5bLtSVcizLHF2kiZRLbp+Arq95
+ciaMnwwVufEFhEJAD/yO41dIIu/vmjZDKNNxDWYZ36giBShynmIeMlzFO6jCE5q
BoaBujmeKaS9kWVmyu+MOJAaoTuFcwtUSFND9Nr3AJOxYTI1ecfZwI7CgWjE4475
ORic4D0xsZrM8OMr2J10I57K8p8zHLk2FX2SVdXCjg48WviFTyRt9JS7vGLp8/eg
q3JvSRs+ZskdX2D2dAp9q9ugbQG4onMFxNJxsZ/z1q+3nIQZAq/UkIoOGyUcLkhR
ptDSMgju9/EKYvR/b9cVTZ5Q45UhvyUxMufryIGzRxLOadvhPRGLolIlrDvIAVZG
6lLgfUgriaGz0qJ5wL9oxlRyOnb9D9pqfMbb15Gew2h0pzbiftX0b5ZtAH4bGVOi
tHXe10ArcfVh5gudRBDiuLdWQwzpLPjPyPzxnM3uJVarcPkHeX34KxgelTvC6y28
53Ybo+Ywbg4QwiNIRNqfQxdnl0TB7v7gSvJriQxJ7PcIH7weF8Vll3kzL5+S+924
5GZfBWJHU5P2umWTkqStBVLc+ZtBIezqJA+RrFXjRfK0n+1MWEcnf1+vv9TCJhu0
4wADDf49VbWYT73V2X3pXttqo3wmC5Bxs6NuP6W4yz942d4VnKL8C3Jd+Rt7h4A8
TtA28og7Yq/LyN+opUBxzV/+Yd8CtHm+6X90bkGz5TZhTeUJGSY+yxYujGqVKQKJ
DsYVOmEhRURcHif/i3zhT0JrqqRUx/ulio07G3vsMS/vK2rdhzZgySiROrriTiD3
MGeqAP7Id2w1+FH+XC8//zcQdkf61mDxRRRyIxf3KtyvBk3WOuGRgcsTxMkdX/5Y
pT3roW6Hntc3z1r7P2r39ZBpiCqInj8SONeLu8p57A8mLjU5TZDkMeMXkNTMyp/B
A065L7tkgRhtTA8/YZsiszATPLIJ2rM4atq5XhU61I5WC52hl0zrtA0WoH6uq1Ou
wOXQEKdNoFEJzmqxb/SdVYONoC/boR0gzznvcJ1j+8felEsh3jGfSwrgfstbA4YK
gNL3FyMb95dd6sjC3oLYjV98kfCC9fNN8z5UjJEo1RNX3vjhFcKZMu9R7Sn4vSqn
ZJnvikYGQYDtAqUebZuIWCnoCkBhcQsoU2gMbyotwvrqlqP9E4PgtXBu5FgwVIW1
WHjRUKTP+9EYA2CWhHEjModvNa0sfk8AQfgEuT93mpZ+gS40Hi3tOTGQ2Z6O2AvU
3/f4LzenRAgI38hTrrWP73JXsQ4hX04TL41SpbB0T3yvPL6+O9n74iPhvmjI6Jy6
WtUQhCOj/Pkq3Kjk1iNm7ksQt8qrgSV871NU0SiyEijWF1lZE9bR4WPs+K2FkuAx
A8LTuTlxjSgmc7X7a6t0sB7gMi+Lq29y9dqRFhJ/rD4iiRrPOJ7RTxaSxCXfM21E
6oysN0trL77d7jIoINw3sZeYkX04Q0x4nARwWjbjOq15f0qH84aAs3jtpn+NUOJh
m+RpsTjM9RWWyA7H+UgR4UI/HjFq6w9xYPFqj0CQ+I63CiVlD5YxAOZz0CGoIV5w
CjgR8NKgT/xhKMkj79Sij6dJN6WUvh1np6cnUfV5JSfs7/6DoIL9oEv725W879SS
+0dXGyYQyotWXl54kN7HwkDRuIljJNatlY7mXUeGAsX8EXMcF35TzeYl/qaagG3e
RH4NcwMiJsDyb7FrctQXvuYX6uwprO8dC6HauDZ4qRhn5uxSviHeS+SIHWBs3mSN
QyR24oQIsgIRD+myvScaeZXBuBXOrXQdM2XA9DZ8H/PMn4JOWyM7DOKSjPyWP6pM
QbQyZwzardSdw6NEJb6PGT3oASib6yqznfPCrYIOsDnG/m1fyWAhyYwAcxzLfXVH
HfkpaugO8hEM7iP1KCHEoZy4HZ7H+xYXQMt7taCJFi3+CSsgW1KKMTGRjN9iD46f
FT4887SzSgd8/lBfL1ZxYpP8pKhmdZIe9ZTZJRftmIDQYCtF9JAFuFUqTWPIZJvW
kmAX/TzmMSH4OAS1VnMtwVbt1Z1XtFLqFY41LUir81S9hFvGyRSISamqVl4LtLb7
OZeAVzpnOWJupti3S7EvIC53/tj/KDEN0LWILS8QDDVDLxIYGo96APEb+yENsJ84
w2cNpBlkhBbcAZwFSdWOe141kwgZpsbI1dVOCD44eL3B+ddleUqgCVYgMjD32Wpr
CmbsgOd45eoRd6wa2YS3D8s28rQNKnXqVgRJ9svkICRAzom1zBLNQtUnVHpHsjj5
xfStIyNcKQhAkKmC16gULo5W++nY7xIlgm959RZRXORqoWiq99AvknEa70IL4apq
q5uO18xx3rhvg/xeMS1Ug9OGASFyQTER2m3fRxBYnqUjVQXsVTVMeZsStB0ybY8X
2RsqkldDrhqxoTFPo3CkkMS+Rs2GdWvwsbsIQNegeLEsgs5FpHzPWYrF8SJn9X58
+S5TQ75GH5KRuaRtWNII1yJ65pfH/14k8FCu2z0H8vvVV+p20p7BDnCbBH9YwYT1
nX6MMuxUGiKr1f255P1QBL6ndAsgYkbb7ef9KViIGLH1wn0kNAnhDMZuDyvzerRD
s/rbypibiiKlonYUMlvEEPqhhscb2kRZS+bUu/SrhpP93IdpHCCLYS1iafME+IbY
qvbNSxWI1gpavZzjqRIp7cdKfcFXWN6MyoLXleYUQYYa+YMS226QDWf3Jbjr4BU5
a5vH0cXEqZjsdFHfqcgG4fheufNJPzLZr+zml5O8Dp0AYBXdNnpHDci8JoKj40rM
/1304l/2uwX2a7nJSWJYftZgQ1ZxIHQsBwnfO+FXog5zJe+vOq6Lrw8NNMMN+43T
OiWalwfbNpijn/Ph4vxRKpGNoa4R6kZypjkO/It9WGuyAd4lxlC12aYiarSzLXVg
e33qIQ1W4dsmikq5UsPPopAOc/UOq8zaAizYJTMzvMtNTY4HmNpf7COUckznWthZ
E6U9oFiaFWPe/0E1UAJMb6cUSPQVPor1TWUu2pS+ZwTBANHcMRTpOE2HhZvAeeQY
WFIuWSCGOoOFDK6mCCjgiS8Ubl0bL/io6khGApNxAy2pAASmejCsG5u1Rbkcvy1u
RKE25vRd/tIaFOtAEf5K+imZMrCuPMlUty0avjqeEq1AtjceiuHtpbp5JFIIErO2
w34Oj5hEcva6gWvPfnZkPgWQb735k8eRZYFeXXyrIQCzAD+KbvqgHqJ7XL/iy3Bh
ezP5KOrVb8o64V9jU7Jl1rvraAy7f0RPNHx47d9y+Wm1J5hQmPx5zTXJ+q962H7m
py8xTlgk/EXW64IyYCwyEP3wWfh8Izmc0zavv6IaUiHcFLYDrGODZhaOgyAu9tuQ
DivYP+xHeJoP3p9aPxxt2ahXV0ZJD/H9hcw1fhqF5yPAz+cKDyRcHZhWPWgGoxbk
I3gpUX+abnw74cYBR4e994pz+NadpN0EatS6yHMoTVl2p4U+9JgqCMa4U0lr6aLt
tJZE+KH3Ed3azF1raxurY+Hg3GcTJCyIVICvsc2CKZXd3wczvjyU/SBYxRrORkVk
qIG8RQ4u9K6GX0MhmtvAI7Jl8N+kHv99/qdsRhKUhZP6JcPvzHnvOFrR53PUVtZf
1nCsJzOYf1+1VZaJsIiWUUNSljPLcAcIK3CurO2DhmoinMrhSxEHYX9uFHHHpzEP
Q6Oh+N0UEpkB0Xv6gpObaqXHl7oa6WlX629CFU9jvhIwPMh44U4GwEtgBdyVYF04
NL/NB+w2TDEeM+QswaG9zAbFMesCLvd/1SW9T1ZmtjMjx/IhGAKm14KujO3o9mkd
SaH7hmrpQsXgK7qxAH9+Tjr422k42fBZ4U4xjGISEPn+08UMsRaebAjiEO6zlgoz
89HbY0KljGDh3CRFlP3Okz0Zgxfe85draDYz+uBU2HXKVS7CbpmcLQxz0Z1cYdtt
76l3NuViRU7dHnJLefMehCvnP0JVaXTbk5o8ppDKgMboOUo806Kw9bMmReqD1TTq
55a+3UqziBLrHt/zueiE+zYZP+Nupr9XPnSFwsMO+tPMiHtFYdF2uR+u7SIY/QEw
3SqSOw0Rnh2p+kgMa/4GLbMvpIwuBcvap578w5QIdMwLtQYNg1Y0tto6JSYkh8Wt
uKy+6qjCdFWCsSTLkwx/d8k5b+WjSZhCf4YgQsyFLjQYPzdGnGLvJ8pAhELUaLNH
2s457pneUJJ4j1UBU4jlPCNb1hZQIIR3bIRtkFEb9vXf0ElsecO5OcSpM/SAg40W
rJl7FQQpjKfKMt5onhi1lra3Z082THp1kb5r9MiaVW+sVbwY07tefuFrea+3Es2C
bFKmKSnAzgKUoXXBezb+f+5CxjNJVvPcKuv4HOl5/x6IPA8/CWEbyMwzVoLg2G98
dwHul6qiGCO8M1YuR0k1VbMayyWJwPROVgkhbPbd0R1uapjLUpLRed7nv9VMhXwx
FAoVjiDFJbDpJ/Id6wlJSb8LAioOfNY7j8EnZ8bJmyFXuxh3X8O6+zikn9FfFtol
dUsYz/hdPiImD6NfDBRfFUpA4JAMuqSL+vMqXXekYSyY2B9jSk8b9r+PQoubyJSo
DXL4zkJd6aJXnAzvWT+aVkeliH+d3Y70S628TFbCASE6HjVY3vryayAM76WQaVGz
vaGWyP7DDJkVTGoV6ZoGhCSJQyKdvRTDYS/T38ID3KuEyZiG8T74udpezjF9ze/b
ONWnGu7O/zqwv8k6JxgmR9TtLpUyxlrYVwYB8ZyPxW741gOVcC+6owOHMVplCbBE
tLjcIr2AKXOMAo1+Jv+Q0j4egAXZ/nodboTgI1D73Tb4+/+LZgoHuN1tPsTERuCr
gsCLu63ygMf/oMBq72fRVFtmVm54AyaI5K9nne3h85TSgC6jzaqp5ASmudxZFD1D
pbIJp+Tr8K18szcpHkKfbMnRreSgBrF0Hce0AGFni547zjf6AUbrcuWGkmchTGLu
KC2gjcW0FzeW2/zCW+A5ArtZqnrnRl7K7OvLhRlg0wcb2Yxt9DRuoPeNcTwOqCEx
0cmsbIH4xNoIYtGdzfqMLCQqtsSh83uP3UOxczeyBLpoYOiNl0PFCA4PNQML/MFf
uxdIftaRt9OUFbVTlYj74QXlzgKL7R6t5NPl8TmL5BfLmPh/FlusG82Jn+EZ63I7
TS8rCvWnLqRv3ENmAWKhbBeaPBLynifjRNPMlJAK+WVvD1weZRORz48GvTIyB+F4
sw2XJInDb75XjDdQ4KvVlnY1nIjmKW2KO4ZvSuXYzX7f1Mgy6kKBbZCGK61lThlA
FzCADaGd374rTnJAfjf9Lc4dDjCbSlkhjIPOyeQQ9FFJlYuHjJtc8PCRP8a0ZHXy
zYkKFrVczwMHp+TmlyYQau9AO3gzkjEuyerHkSYz0YkifdGmr9shgOxbXdgi5FhE
6PZmiPDCm4ImQhb0kzckZkZnYo0+6uo0pmjKC9rEUnLiejPypwK57krsJ2ecgevJ
TWbZZfMvtb4QZH4w9HgqrlEByUnAxbWXF3Y86h5jjsKjD7dlLcrIz4bmr44Nn1H2
caUMMH5yRjDHnhwIQXIgF2wcHvKhKr/WnNslda6A/7JZIy8cBvzwa4Ur1cwSjp0M
4WK0+iBxzX9mfkPtPXqimvIY02zHni3FhJKoIr/EU9G/5eVKOpW9WobHuH3XJnUj
35ZrxCTfrhf5eunKnFZHY7SczvlR13Xkxs2nyS0PGB1E4xG6MvdgC9TOKBoItewC
sFn5ZxTWAfmkvBzMr1kgDhIG+M5QsPvSSa2Oc126ptTCfeUEtJyTdceYPnhc6ral
YDyAu77OKQURWLHphUDkFulU6z52tPu1iwJW5ZHm+SSEMJIheWo6aFIExBi1mQ3O
CNqVBlOdr9o3tOBCv19JCgDBKIMCUC0sil4tF5dlY9VCp7deuFTyvJnWAgOhZlRj
BbWDRWVvw2UwfIIYWBboHyDGJ9pXnv4emLW2WxGthRGdymEj8P6v3SBnlrXXhK04
xncknRMja1IVBFsTnvC7ycFMYWmHZvjveKfHGBXBR20A5uxev7bP75xZ0Nr73Aai
7eBt+9uoiSZD3VGhsl8NeO3h0lC1S0azEua/udRYVYOfWrAbcHvb3sEEyvHpP1WG
T9ZftyKHseMmZmBbRuvdYEhXmIqvDjWdek9BpEcp3hagw3M3gQW3oaFCMDVoRfOj
XhskyrTP5LEPbHXuCx9nyHwAo5oxRRZnIjkvgnJO+bpzbIqHeRfURybf8tY0gt1o
f2Cy0PiFa9dERnCHd1c8DBsvv6irCLXq8Jo7LfOb72tS63zhPsotBmrWdM6JV9qg
ch6hUOBZelQtsx15XwC0t79Jt3yiUssVXH+In3JBgYvfT2rt3MyETMP2ym9xPgg4
w6E4GZ2wmkXBCNNTvAsi9jeCQkar14Ba+JQkOt6K8fTnCG6yg8cUmNF5rPwGbE68
A+ej26ibZlGm/UfrUeoUh9z32JxWyq7zE4Dus77eysuDrlec4IzNZYlUE/jEbA9B
yDg00NOR2DDez6Aymho/8hxrY6Am/WlW8SbxZg3nG08dTLzHdrBUPtKQ9fwYlo+w
wce7eehDS152ZiT7P4HtcOm08wIYR0UXmXAuELBvnPFsxVt+pJrOQ1V0j+fX9X9V
r/XbsK+USEWsfL6u6uskopeqFwdY+n/UvpzUBV/B9xai53utBhB25/BX8q3J6jdC
rlXah+cNFXDjeblfTrzzfyoDB1FxiubwD1XBtJSlUlYQRwj0azNeWjLUU/WE+UIS
TbuuttzPXgpdYt2SOTiOCLGpI8KfpaFfIyvDG2iw0BTzmuTZyUAnlx4JoQf6M30r
6umRcGjkEazlgC6i+cJwXBs+epwz/qEc13iKJ+SHMpn0ZSSHscLcPUJJpUpg2B7S
V5k4bNQsm78+H6f7C31TUN/qc5SKkvIjI+zio2/jf9SUKUCUwsLlKrhwVy416aZx
FmundfRgm/xtY2FSbGKNwZySncPcpXVXM7HSJPKD4jECeNrGtNV4sUYrwizjlVDb
72sJ22Wyofc72RYvokUDR/JYUX3T0PWMYd6sJY4PnmpGjqiI9PieHJANjSPB82UZ
G81N2JdIB6uj0LuoqTrWETKf1wZSxbRBSoUOSBSdgqJh+bh71ktgvpp0Fu43b4pa
aK7cK+//BjWiMWm5EbkjW7fkc44PBYDI7hPSDQLwWshxmW6YZI0m/IyEZxAGZJgi
EvS31fS48sMbJBOqNY6uXNgml0UW9zaYvUkwqHJDvpTyjN2l3ib89bJKHwIaSgOi
ioS724wn+Lpi2FzvvaaHe+ceuhIz+DNc9dle688yGMWkhiZAcSy8DhJc2P+y278M
NLeG5sTV5DwDHtAoSo3JH7ZcChFByrXMRIvOecbMwb/hZst4cdNgl9eZwPVABu9P
rQVbspgd4nURADom4hE7HQhrYhAQ1REVPdjjwjBlt3T/ydjC6joTmfs4XX99vsqY
I4T0vpCD+KC5OoydgTMXR8hoBVPoSADhEFHztacTPL6hlfrJm2s6kUHvuuFoGJhF
xAL1cpAd8k7clq98vxRf4e2FzGkb13ISh/qmjTsP4sPervmx4myJozBZw9JU49DL
mhdhgHyrDiiCUVLtyhS9HKmYQHystH+vfQuyb4jNGlzfcHl7CR2jkGn4eJfU0tbV
lzNfXYU5uLuHxshO3JI24XQr7TyFkMoiSrXDCbHnKTMKJr1aj4a36ELls9al+Wu0
9uv1xYd91R9Sq3N+XW1Rvzogz/8SoBE3Yg6wwCcRCxRLKjdBZZNkYqx3ZsnWpe3I
vxMBBPWD5fLgKs+tUy2W97NJl87Xsp1v+wKkzqlQc0qVCO4c4oXTQrN/2q+ot9Ce
xqE69SbEsnWge81GEN/YepXtKMl5YNc+W/y7kMUNgT47IWRA4biFJGKN785iAkSb
ErcRyrIxkQxtPkljm0yihTGu8BTdndwZBYc57PydXj/zDgXb9hHibyY1agkh8XFp
c1S2niXEbGrX7yNCZWMSNXmGIVdjLkA7ELMTQsktnyGrZpwnoeF34tkvo0aiwnEN
GrB96PB4h0C5OHdskiwVbu/zXr0flKi0FybuVEar6+EJQdNPdATAJ7KIE0C9f579
y+wco31MNx0NkuBuBop9dlGtZ/7qhUr0cq6Uu8E27btcTltin2OCrnoHCdgd5VmD
MpzdEnMK9PKZZRRSDwjaEQnql+wvko9IH+81YISECDEmWTrV/VCXknGligAP6n1n
pwGQonCm0z+C5Lb9H7A6rodYIS+7UzJTGAR8owwEvPYBGVHNU0hwbw2N3d1bVjJ2
/gk5buOpWErZcUo1UBI+VZ4Rrw/7KvJ2dYo+c4kxnnp4JyheBPTEWdypZEkwRo9o
4t+51BQ39ZkhDNjN/CeyHaPA+VNHK85QfST8VYAWdEN0MP04Pxk00Ii5pyWFRAtK
P/U3BGZJaol4lTN0ngKpivEZXlcwtN4/1Ro0/r+BgbQD+TlqDXXqHh7ZJUKkt/EV
AJXv8tZuxVJ2/fMEAcXkE7dODzX3VHEmmHS+Ea3rRxLLsRrlB+017/YO4KW6Hpm8
6el717f+YGBHmvexYhRuI1xeX6dOJ2i8i1v9g/NLKuv8diGHANZB/eR67kJrkyXt
hLbosLikgzTq0J5oDKMI0S74mD5HdULqxJlN2Su0TGV35bugRVYPDl8Vs3YvVm5A
Izs5ylOnjU/TSbJqeuO4L9UhVHf3wY+HMjRPPOv3YFQJkoK9AVsRCSYX/BTSWOUU
+w4X2Mz2WWKju4iAKMcdaUlxMHN0YsU+Ev0+oxJaFHkcUbRlREXaxf5u9DFe7ahr
TVZSNKMBpDI37vnRFYKdr0a2nQreKajmGWca1GAx2smHTeoHWQTq31eIfhTahl1w
4KS/VCmJR70jf9Sqt+//U+MgepZQzU2yhqmjBmBY2iq/b7BoigH1guRCRaiTlVa7
jBdEF7v/5LkHJd0b+8KHo9o0hfNk69AbiBFFy3s3LGQtD9uGz91FKQBpWMsBAT/x
UxYeSghAjyGA1O6UY1XacOHbsiix7qoKG/ja/EQ+eO0gPaAwkspME5tjBLViLBBQ
D9V84uhMUWiH+zzuVx9k/KL1pDuNJv2ndiTL9L+kn+XJB1imxC+9U4YBk6XuTQdf
/F2fQBHp4Bru4qsDKyZj6jQyXoxrg/0gWct3OR1pbhO9tDMeq9JqOx3uQ9HH+uWB
QTL4ksA5TGDNZn/KrFHh4CwOEtXQE4kSaWW5IfoCPXosfv6ZKkw8x86GcDS/v6kw
yQfvU4LYnKnHbaZqpkTmAZTGQkqkXs7Fmd2mh+w+bZQkWtnwEsO3H+F05RK+fRkw
DE0prRL2uT1/fF7o5zLAd1nnf87RWw1194S7pLBh+TrFMpj+RdC+vZvK3NLs8ik1
Pj3IFxuOy2zrR+LwD5dMPnwdBlqc6deJuDpBK/5+8GLSL/qvC/kCUuY2sHJr86W/
cfL8S0k3E9Opnsrq+UQxdPsDaLtQiz9Ou/3sSWMC4IjNMobLq/m+AOKCpEbwso+N
MGNDRKO/2rKxv6IDm6X/3bzRWhxArcm6QseTkEoWdZipo0o8K3BR/5LwN0zpWjP9
PX9mP5rcT+q+co1VpQ4o2Ywtp3CQYRRw7lPFtFQwQ0Fcwrdzsj7ZU3Sl7ZE8LOih
n2UCTwlxcwG+fJXKDRkCjJUHY3IoNPSzG+t1XczRvXN/Cz7zCUL8wCQ6xU6E8CbU
RodLj88IbZowKtbqiZpfRp83gPR/8G36bz+a8eanyRifPD7khjrOBRH+iO5TSssL
GJvQJDclOliSBgT2Lz4vLwmFhJ+W89NmfqGfWBOtHC+I8am69dVsTu2uPG/BzUFc
LT7Xpa9w+a8E6dY5cMIAVXRYvK8w7E7aeHETkFbIo+I7Vfr9I+f5U94HhYa956XX
qpnktIpf0PBgE9cH+bjZNL6hoEwrNB3++vop9C42Bwl2QdANNezuoki3bIE2waL4
YWuk+dwR2aaZEJpsYz9hZJx6SqYmvYhkhYXLHpVpvL4z4HJQqWykSCEhEVjUyV8i
e4eqnmyH22gt7dlMwISfqxwBSlfhwVtxEL1q1ugxycjVpBv2gvKPG0ItwDO5kEYW
mF5Avd6LVMT1RMy+jn6EjjmumvcJGDrr9jSBdsuRNu899plYlBdxfpW4azzcw9uQ
w13eQ8eQ0917JcI+1j1vrQgqrthDLkIg9SvKK36HN7Z/YcOxH0evYXq9Nt+duv2d
sjeby+fwrrZmwy6eTV4dVovyA5o2gG9YghvDk/nDrkki6At4WAWaRe1a3+JuTUhq
y2rg2NMIGcnrDPqxYZJtxKUnc0HTI3P0yXgdTLhIe++/ye6+VC5UvAygTWRGvi6k
IzoOhmUED18auNDBqCo/0D/hQlEf+8KxBl29F/wrzfSXtosxFQBA/qARtSU6BMqe
jg+vLyeymHMFopP4StXf+SmRWwGDzW9Nw7jwL0zXyHDWy8c+q2CBjlVoklPf4X3B
B2oErIyabEfG/GUiObVbRzt1+oRKdtpn/NPEwD8WViGfzBVn7UCD9lAranKM8vFz
FtPk47jwfmPHIBwaJ/diCfHPXEKrN49etNzqeXKSB8Id4ybkwGMJqJ1tBjVBotzO
Mm31pXN7dzF7JqAUMHRkcmBKpI38X3VLF9sbFUbG0cgJEskyVjKar5zqBWUbiZin
QcF3zzXCVKsmSPXDwr2HR7pA1vkf6xMLpFWyWyGskdka3YCP7DSr4C1sLyBLEv04
H5ROuAF6ZtKHWooq/nPdRo5IrTofiT9ZRDoDwGfl6SgeoZoRldr4PiLgz/3JKzuo
/7ghh1DvKU23UFjx+rlmN7QqS07g5ifu2khCLROPqqIRkOjCQRg14qQQgYixGA15
ZBnETlzIHeetfKoox/E6gr29rKLmjRnG4jcz8nxSPS0V8mSnISu/ZYIoLA6kD8rC
JQj2YAsNfPOaOTYxyZRS85OPsyVXwbNVcmCQedDa2RqH9UZiIVLmE3h4W+VyUAvw
6zOX04deQtPOPG69vdueS+DsGoKZ+XNzYJFYMLWqE4l4dgFukY6E2FVOfM+Bl2Le
IOt2HzDrBd4hfyqZzlEVLBsVRjh7+jPZY3Upwl5H1myZHILc5bno3+xsWsxO04Zu
/7PpplttnQtyHXQn6tw+Uy2eQdOpic6CV2A5wT0g0UKumCAe5uyznJoqWZ2JgSj/
02QRqrcewVTqiJuQtbOxkbcYSbfqzfcd8drcInxCCm4XHdP2SXq7tW0kX2xjjybT
qCD5iljj/6EEaHDDjcSmu9jzWJcc6gKGIdtCcN4WKAf+H9Va64YGcvpUKsNPmiZO
Yaaq5mR7EsViYtxKNJpZHmEwArvnSMmAoIoudcLZ/kyXhUHYmqJBtlwvST+XcPZK
zab3BrDS8GC3W0R4AJQmjQuqL1GSUQJpT5ojkZehn2Z+Pfv4fsH0PqdCJiN1Kskk
toetWFnnmJwGXX6Dh28dAH02tZvW7cwq1tkeVCuZLgR6OHIuHIMmWWxHmOOrNMcR
7cCaVZmJ0fiaoHmtJDk50TTWPjEumL1xvxhGMWl+Ur5z18D8R/8SR5Ux/F/yIctP
06ify+xNHmtlQX/Vsc0mvEEad9xkSQG4AvGBERh1KZIcs5uxMrlRj+JZrA4NNiPM
bao3h4NFQs9Js1P2S8WG5H96efsycVpdsGJgIMpItLsrrwMSsu2YeM/Nav9ywhq2
Wxl2xnDHBHOSmn/mDCnEB35m6cIzIzszNPl+EGX+oJfxp7fmrHnLWiiKqZCNljJT
nqQDBKmhsdD631q+BeZ6Ql8PIU6EYVpNOoQaSmEq2fRj/SYpoeXgDBYRo3dHB8fT
gaaqNdAXPtqefArM4T/z546IVPragRsquCcYH5cxxGyPlUOKd8xrATKmBP75SgE+
dQbWevba87cnbRgtyllowU9YSK+vGgtCu6Fhl+BB5gMl1G5+iZauiEJ5MLaFPKqp
747cvzDo3yBDP/JusdCqisGuev5PuCAaJXYyTBdvO4HM0Q9MJKqDk7V1H8hTWh2T
akwWY8DoDSd0/Flkr11KIwDY7RZnNlWoLxfSzHnRV/SgeUb5qZTELPVWj0f3vN5C
TpPiTI4XDVxCsawDm5DIWEMLaoqFxULoqGwAHi/p5qgAiUNw3jCy2jaUtv3vezJW
6pArhL6AiOSJAeLV9zxsh7581uvmvPbhlIzs8DBvNpDc+RI9HBJTnVY+fdlj+dHS
smWeuaz7oh2otubVoSK7BzYVu1TRyl7ceLVT6gAOt4GPlywoUMDmvuo50AVQQuVl
hZICyq6uyC0RPIB5mmb7gZy61ETRGG975kd8V0Ad7kuZPzKypmxFWSF7kFVGw9Yg
fUXUuN7nIX23Oc4u7XnmpWlEbioqP/e7RCA14oGncPxLDEHeGiJjBwT7ZEZaxDqK
idgGCJAiamgQvKcV6VPGmtfv/rs6WmawEj519fUt9Fjr4TW37kfkh2S31pIyRONq
YSDmzRvmz06SNuu0Ol7a2c/TRUye4QMymokY9wWE4WPtXeqGP6vh3FQc5EfSn2/x
pHJSzKEpKaJ78hU7k7rnumsqpYO6I9vhTK9SRJlozMXBWiWSB1C7V7SzT9b/xBGj
vC1BiUP135pSs37lVC+VHzSEU3oLsMrCNriZsGz6bLwnkAF7iTB5vft/yJzf0mNx
ttB2LluoxH9PiKUt2B/p/JXwJOZiyOStOPMnQbX4DZkzwhE6Um/Fe9nxEBIvSfqR
nQ3nYiMhDfK3piu+xOQmWkHoOXShYKFXlsXAT50pkZAzbc7vaImLQ/edf6lpMGnz
LQM5lyh1/I/PD3Qo/iqfFyWgcy9EWbcdabcz6TumvEEEzkZu55tPBGp1ZtRFJHhg
Jkd8uo+URZWDIXpK+BGaTI+OCLUBfVxKX1MxhLFbP8l1SPfj6Nd3xnwwMO5aSr+t
UEGQa2IclUVm1SBrZbsOO1o+k2NZ0XPELTffkrbYMfPeeRgzaqfyiY6XV++RDwt2
C/y7XgsQwdFsrSvX1Y8kOM3PDTt51zVvEQC9uAdwsg0zNYEJrcpZEzEOXaL5dAFO
iBCMMF4Mbi3X597HGPhGzRNDnmUVKYDmJzADsNJdZuOY5089J8X2/VnTCemomuC5
LGE22oqcnhIWdzArLqk4cDUoU43VAROptNqHnhvX1fThGuRwt9FupS7oZGPpiZEd
pv2/tBZ+EBUyylYJvTRfyVAIMMo4m44sZEKBS7hTpMwtXB4ofDHruVkEymreOOAi
3ilO7VHDulTfoN13SD6nOoTu363tTBpnfZfqRK2a1FHKWb2NSHsLaZ+rC1+svKNp
Ek5Jreg/NCYxfVvSlD0rjy3jDeqMJPnTJsfZjen9KkD9xCrfj09FG7lT1ZuGNYIg
z9bRAKrtiTJNFzM8RhezfIew5h9UZgi/y33V3Y82dtIez0G6Llb5Nj9q38rheXn+
Ojgql//nKLMlqfInFmNv7MSPMNA6DB48NQRQIWu6/GZxyX6aHVCp3Sv2rR+Y8s03
uqgG6J5DvoyOOYKeUhyTG95QvSjU7Z41JHMdxv++KX1VPu8YD2RwRkAOWoDi+XkB
NPskzcOVjIOCg6mi4J2svQGNXyQvGXLO1MypZn27A41wpfeD93sypcYUuSGrsvTi
ge07ImgT3tuWp8jTbKCRmIyxPqEfoFOihr9NEp+YQusM2dj3j7ghGKEfO6fnjGDa
wJEW8Nz6FniJGRpMols/G3sTvkuXKkasCNvBmy+ci59CzWqHAxP9XgP89fPsPQUc
CSzPlDcU+tlm0e9qOUpqnvgH+fNrSOeCJMSD15qzNWfs0siC4hayPym5PfoUecq0
bHNXZRizdmLWp1G1+7whuVK6/pPxd4JhZEuJfW05q46T6HrxQYuPo5fygnMiArFk
O2QSWpe0fC6Wbv4Def2L3UnG9aJWsqcWG+z0rl+Vhre17h7OD69LbvclxSiadzer
J4PHcudfPjLGFTa2CSf3/IdF7qpSiQtLnqv5Ubr+JGJtEIT+Epoen/Nx6oqLvNiI
PgI7HFnpTGw2hE/xhBfs3acPGPo1kNoj54stkOA+psiFouhjSyAWQ2FhaKGqtZQe
c/1v3nvJVXO6fx/ZTOrrAJG9v6G/EBGYHHoFbfyZ9posvlx2wGe7NFa2Cz8mJpY8
GMTt+8PCn9FWMs13REMwe/XgLTMD3O4nnxjC3zTpCiayHpZvI/ZWccSnKlqQ+E0N
BcjipcJ4Qi2h5K+CgCej4mZdN3vafjc3mgrbgBolDtzTn/3gZPQHUe0ynmkql1a1
wNIs27yonm5gYB/b20W1vn57elK/JveN+s2I4p/2uGGy+yFxsvYoCY6DsGtOv5VK
iKl+6EFZ67sWqq0tegO7F85Fo5u6v2Q8GWNx6JAiE1ovoVgadhPM9TCSusGps+cr
suAr8WEo3e00R7ZMUR5wj2CXnccDHzPvJAvp+tPzlkr+W6x/sDYk5x2mqE3SLLU/
Q68l21pnV7WzuVvfFlsVqCYmDfBNkzjlymfLzx26nTYQ1trNxJ3VYJYMZFPr9YTh
5smV54clZUYLOZiCFeOPLGW6zJyZXmjAm7dGyPrRxo7B8iOYNXehxGZ0CP1XVl9b
VQjgixbdl2+yDK0dVTrBPDmRhyc6r+kgPybEMCliQ7bkWjfu4ox8N0rKqwqKt6RR
F0Guf8baVjfyJy3Vxqr8vyINCuuTo7ZGRk8jFR80xZTrs9X0NHd2T9n5/8yuvorS
ycw8O0VWy+IP4E+B4Ty4W4DU2B4nm/Tnitl8Vbx3k7URlKjgJtDNPhRWmEdmaHWW
79jWReIk0wjR7ZVuiyDW2/z8jLdCek+D8386U8HJZo/jvTqEaIxIHhZa8GCupKDS
5PLh5YOdqH9NwNWmNWTqPCRPbQBjA/scSn/PBVn2aogfsc5/OSnyz3HR1j+7LDLI
U5Wg0r6PqtzivE8J+zaH2iJ+aE2z4Ohe/YicKLpbAt1gt3QhxJQvaTRvZE6TJpdp
FaRwccn1K/FEdcjX3X+h5WEE7759NzwmQsem4SHstwFyiwWI+uLKnDEFZo5skwtN
kYsIxEXhyLlvFsghfBW3b2GttEDW2wQEE4rmJBjQWzwd1vMa3SOsOVHHveAIDTNh
yjAzOzKd554jAMxrAo/VjHFR3kmNyhKSywGQZK0SfEcQrQpnXIxfwyyxYVMWvIim
p/iEIblQrFOmsu7e1mWWylJubjylweHBOZODiyxCND4bl6zVbp9J7oF6NSXNlfl5
FsZI1z8Um8w7Gp8t71hMGAvIOZl+s1hlpCXszOfSlEcXKUagEfcxX9OeD6oR4hQ4
P2Aq4UWbefBL9IaWU1cxAe6tEJX3smPKmueey5rOjGFDxq++mFn/YWxZKCJhLEcq
XVrXSyAzIjpkJXagNEajiD6QN8eTR3qTXHqtnE6N3HTbzQ9ZB8v5o1Ogwp1HgMhV
OYTRfFzkAGFluGlmSzTGabdAwRTsMEjhpN60KSiRUJkpN5nphXp09wzPJYHJRh0A
hpFdAOLvte1N6PMtxs4RVyqnP8te4mItgnCTgc5ZSyl3Lg4e05/Nhq5K25Uo7yL2
bEK9xTjffSXghWN53sVd87rjAv1mfBLm3YQeHZAjOCdx9tpNjBs/O6WL0uYbSkC+
MzSvSsD0qlUkUNMhUGkW7YrYwS90T5diJaeh5DQ5hsVHWEuACPqUwHFtsDN3IQBv
mG4mv/qN6pG3KzJmTJ2Fu8hfWNiE9weFpLKud/qAN2dq7/0k7jgoBbBUZGH7FAY1
EIbEzY6FlAAN/fAiWTfOmGkJAWfbD2sJUj2GzKZ+r4Z6ZZkSVHnLEpuk5f0IekLE
dg2o/673/ORsuMVhXiUizzCF0kDeqCBke68sWlf81uPfYvMCXSc19RDAcSx7j6CQ
zSF+hq+ihZ3gow3Sq3Oc8wfZ3lkRomovek+mzYSlQ7k2fZiVqYsORHA3/SzzQ/Ge
rlsfNJHmQPI+HtBXKhDoC8zn7I5BH6hFm5Qn2UlefsSgRe4ETQgwgUa3Av9Zxehq
O1dkUUT2ZcYdTJfoyjI2y8y4XhEl4cgVH8hh/1vFlasGOBXi6E9g5GpldMjDaGBo
iq+LLUygmD++5BZDsKKBb0HvH9sjNU42bIykaJAd5TGbi8qfFqAqJLJIwPzGzZL6
j8aHUHqWuYPLqC8CoXX3vzq3aW7BMLmfjpzdGub+ay4r6R1FpoonpBzUUZqnqzid
mIX1X/ICPYcGG12P6Q6ep8dMgGapCDDBzhyReF5wd8Ul0I6kfPfgortmwzWDXfUo
rbo8hn5jrq564QAhQjv40pJiAuWSfVQ++hd2dPjBDiuXFSWD2GFq3jhmGGEJpZos
i8UFPLsTh13otI3xGiRORpyiGs2x66nAcykJRMROC77SHPeKYidSHF1s8R1eiMfT
uTmvozp6iqq4yPvSWGK2J9iz+i+DJU8TVRfOKcxhx2/YkZmwMlMWRdG/QrKQDp0j
pojqSJ+BEqLUAw0LWqxF7JmqV7jEGaiJAwlAQUSTGgt9g6/blSS85zANxiN0qroX
B2Ue4zHffW1qNPvPfyZhL3RIYvHysSJWGgJdL4uFxDDpx9eSjPd3ye+Tqj6P4fko
D8EgQGfzzkQ6sCB5A1K2QFBUt5TeOzFSCsoD/1pGkvbbJzJF9qUzggKbv3kanL7w
KtRIqMgr1hO3lJQfa/kf0Q0Lq4VBGMoMQrQ5fDKWfjlGjCuFHPWk/otPcSHaAHRq
0vCQFMUgnDS57sElvP7l2pw2QGLGhXa38QvURVW2MbKQH2fJw3qlRK675klYXWc/
7qXFAVyiACq/qJBLBsQP4Z4xEjUVfokk4WOFdHVJlM/ANneW3/+pbOHXI5KmVYeC
v5TLPmi+o/MhTYVLI/8NaOgQw85xy3tFU6STA3pTUfsCGTD/E9F2m0zLm/98HE8f
mDcBWY97oe6M4Crhgs0vXb3rwdNvT73CbAQZqzN+zMYvA/37ZwsAZa5569nkZKbM
dngOVWgV5Pex2A7rVtOIMDC/do7KJSlu7iVEpSkvfxDDgGI9x2KhWt75Gly7uFOh
fuAsFobeIx3wW4t4HKbT/V0v0G2LRNfuXu4TFxEc0budLI9tsMmH+oZ2Kv2Dfkrl
JoI6yBOQmNvAeRIDJdYKLkCsR7XYPw0LiosAnuzcoiXe3+t1J1+XiG4qa9nqucYZ
o8E38kTBRWqoquCpFNWX06WlERwMtC8VHavrf5uAHNdTwVC2W6a/qmgKmL/+aQCG
U7VTyTOkW8qQFI1/5hhn1kaJBQ44PGYJE/il82GF4Y1LfWJRF81Rh8WIOB4a55NU
LZVcfg5qeULd6h+mZQ8G8429HdGVS/f1aBLI26bkRvXiyeIhmVl1fFmYXGBXzY4b
C1QJV/hFIhlRUfIbOyXutP7z2/4mV5S9nsK7+UM397L0J7irnsuWQKAmZ9CQGxl+
/uTMI+3Zd2FOY0NJLpLoCaT9VD+LpfgTwfL9oLMqLzbiQx2ByXeh7aAXawgFMKuu
glUDqmxpW49rUTFLA4inozlIMOwVVAhiiOewqDPtuWrKtrLwTxT7b4KaiEKDSjmJ
Rh2czqMvQiEYcIl0i6rwwkB/nBPFiHuQjE+b4eKdycd3EoYXwG+KzdcDge0ECvZI
+0me1p6kMOYFsbwc8dV5oanAynVZ/aM2HUdM3CJZfi9sEky/cLv0UmS9G2eg558C
pNbsGAAfwVchbrhglA63ifZBIoDCzUoWaLqJMzR0pM+FsklucA3YU4ySVXAlCqC5
R7+XzFOCtY3BH3y2wxpkDA0NHpz3GwPWg/D5ed3dvL0Ah9a4mAgS9fvgnBe4sihZ
D1jSkMobJm/TMKF4ccPeRvDW9NA3u6eL2TeiL98N/jV5gr7SNQ2JVPWHluMYsYYi
YqoV/yp4rnkURFJOGcE66V7BCOhxIGBJeoV5+KAcAkANbJ8oPq2rnOdsPQOsR3ag
nhD/praSKUX4XIECW9HIlervDYK9SxT5IY8zSPU7ZZn8HHUWazTGVj1M/KEZnwI8
5YGL5sHJ7gzRcuC8jiygU/DqIxm6LnDPOw+HT5cCeBYAbS1Dr9G0dRu0MU9+iyiY
iMTJIZ+RRubudTjWHOSfSQbfeyUihlmo1cWjpAae0zClShZFiW2ktFm4swUnGGW0
7qMHLVbCe7nGibG5fD480bkjmBNA2cecDngfjwai5hOe63gWmqRg3bJiDiqVK9QD
AkTya1lXFovwWnMJ8i7gLogzkiAMvCvgPQx3p7IFJGsncEIGSg54i3cqxmcdJimR
ImDjy3TpcdGqZTA5aHSA2PFboD9+UGt13fup3lwjcJOfSroQsODDNsdkM38FM1O1
LuPqNoets2sKCC/TMaU/AXtZ0skh6e9eJHJRkJd+IGo4mtLzxkHIttWVUcfFkGPk
sKVT0BCQyVkQqrJq8W46tRJ4hAg/m/sNxrkdOViBmlPmVp0xCU7M182CR8zJLsXk
UuXZXK2+foQPJSeSxHi7x0rrwCh6bb3FNCScfWgthQu1G4kFmkaLkIX8xIxGsmrO
m3ayT9YxUgui7vpNWGbs7I+jW51g70akQr4A7X6m1NUP36dyTioIioAzLxhS3tCN
A+2jYXs4sFcvpWYc1jriTfv1YGMQr0LekYW3LYVOuL8hu0OnUGah25GUL3rhKLqM
eOBcQsKFg9SdYr91FRWyvaTPxJRmGgxMwLJXlW0QiZY0CBk2zYMrsRHD3U0nIh8E
CxHOPE2bEg0TkwpwmoCFqvM303KZs26SGnJSPD4Ij3Z1Sn8quhQXfrpPzg+1gDxT
npYYElFmMRih9B6hOT+wh8Qxld+nIyJLe4SKfEIml8o4FLdGWwMprmsgQ79r9x03
9gvuFHUsbNO/3UiBuyoNwkIEsTgrpESm83KpQz/i1TP5I5kR296wNIaYhuYOoeQK
zVZt75Wk23W00+XVBaB38W62ho52Hi8wdJh4sVQRc9IgbG19H2Nnu0LNWVOx6FLL
4ccXvZyLlcUoS/hS9C/175271MQabShv/2jLtMMtEhwUU7ZxZtEoxleuSGYr4u+e
hJlNJ6Pvy7pZzsWDPLPQCg7ZJd4kRVKxBjEuGSxg2to4t2FU4nDrzYoqvx54iCWJ
+V2jNgNTqdU1Fg5Ia6GNlFodq7sZxCvZbLJzM+pUY4CLC3x4Tojt3cYgkdbXkFM1
7cpc2hVbp9qUr9RGQU+edISZmYPJfxrjDf7sfHdRCwDe9gBuy+dobfyEIRVpVJjN
PiTyPz2qWom1Bn7E5NZGzO9izWJlHW7Hz+3Wb9FfdSNchpdMhBIa6Ryaq2/0bAaB
AfBtv4WGxvsxaOF8jG0JUoY06eujk7pS5gsqTjQZ2rmvCDXZ2rcXtWHzJxXAaEFS
d0u4/FU0TX5VMVMbReWkGPortIGfGjL1CMZmTxQBpJ1B7dYMJBZyWf6zR8Sgx1BR
iv92kRdrXdQi4XfTf6Xzx1ORuFQJ87M0fnw4y40omilJQItw75delNlbq+YGGyFJ
E4XvUGwBwVXxzFVga93Fmb/hfG7SlPmJVxIuoWQ0kJmS1YYh/sp4v7ZxI86074tB
n/6tF9hXCuDTp8HJ9AuX8DX4IcK/CjFZA43+fPiSWIDeQXAyRyBID77LZilDavFl
V0NjBVJLP7c9V6UYLWyVhhiLkvjV9aXjDBDmJR0wP+QQzuhUPmhEoBv6nXBWHK/e
uJPY+tXL9FgqIxcCpaYxVJIqPKPszglaxWXwKtJ2jiI35mlB+XTp7o32p59B2G66
gZd4eSGydifRYga0TjkgllqixCiYHAWtWXw48kpq5hFag3CB96Mx+UZ2LaYdsF0Y
IrJWaBId4noDjy733JCWT5Og4vMwqVj9qN7nC25OBFZdwCOQBtwhLQUTwHWTcOqf
bby7/Q76tOHGWzNCjhov9upd3SschE8VdcqNmr3qD514E5aOu7vxQQYzwy3ZXE77
u58BGNldZKH7kUufIkvDQjsm64E3pwEUg7yUAWJn9jKYKceNJdSOI2B4qkUIZX42
XQ6sjH0DWjXEUxGlejFMrFuuQv+JyydSsUicjeo7ik0gDltpEYxWcFMkIL6onQNy
Oxr/cqQW//j7t0BGdz39CuSasSHw4PbSWnSFJBl1ozo5JuACpYIYbBJQJ+Yfnl+S
xneO5s9X+dKKmcfnAHeObGsobMyIkWejyyS5YtO7eidiA3/IdFr9jkFQnlplFNwn
fgR9FuAeabqLOaegJ2takbw2BIKXm/xZNE6G1dOvmte525Nr44VXWNpm0RuSaq1H
7ukmX9SGotPryqd1LOy9Mbl5ktIvcN0LtZSB7drYmXolPkmIu5ziHP/BoHBJFH7f
SG22Vg2q2mcx8ZnOfVbVri3tfW8N/y+q68urplw5YdKFI3HMzTX/dMaBpEaa3yPF
h5qBhmvTNk4biRBz3WKWD9gGzcntoHkho1BVpKXXJ7IeGE50EL9PIi/DapCYSm8l
+wMGJG/Z/vTVXsLhJ+WyaBXFKqo7k/vQGXAJOaIRiA2x6cMsfT6t27iEP4ZUrRJA
fVCunH45nZNxwSBsDwJBlhtEyTz7cc5xDXh2ps97+z4uKuxOCdJY9+u0XLkPDnJX
S23ZW8cGQ9Ws2XUmeXLpyP53AiPvjNtlMvQUKIeV1eLOQvaGoly3Emu5IItqFGD6
bO0vq5WIHwTVeq/h2lYfqneDXZdn2B7b4pS81tSjrUKFku3UgL5ULpLPjZo7zzCV
r16Es3Zap1U97BVPiB/6BOI9KMZQ9g/einGFsFalxFg2mP+zcAnPL8LggZTIX2Ic
wo9NdhAV4+KqzYRPSyWUemZuw80LCvuuoa9Ebw5Gc8uSJZ4c5/G2Kt+X/aPpxKNz
XXm0JQZoZm5Os0GWgiLC+9Mnmogm2I8eMX+biJpI113HW4cJdikcx9QgE1oIF6RH
XyszriPXXXe1f8Ee1IV6J/gJp7AR12aH816CmHN4fva7zpLtVYDJHaFzsQMc71tl
UTrAzMtet4BlOGy98QErGo0iHbfoz/rE9Fg/VHsOPYaqDl7K0cdlEhPtR/GcPOh8
YQBpu66b8JV6NnPQCZNs4Y/+W/UUSvoDyhygolX3VI3aIYN5/3dXI81dxYi1Np23
41g/f2jVI6U9l6TRHfz5qBqfEFLAEN5EwmZOiATPXJ3ryLR2gLVcjbUAAl2jvMER
KiVxCK9HKkxfWZ9U0gp7Rpzlyo/qw0jdm1F34JKBcQjOpbIqbccyWjcThnFg8NP1
JforAAnrDZ80yWY5J4EOzbezkKg1hzyY5ovwRQW+qd0dC4p0j/CPuc8eC/AbJCFO
+dXoLgAl6N29OhViaofli7BfaN3dGB57ELUpEuisIWDdwBnXF6Nbvdp+4hCVjiGJ
6TogbvW8UuP46LhtwE8HOZOrSXZm0NILGpMuXwSXV4rcbUERavR9IRu6LUALvYCy
Rk4PoasO3yDuc1PsaVKq3NvGN9xF1+5KMlXGicXWhiKsthV4gUVzwJPAKNcPre4V
NWsqD/5/F83uxVjE9P076kc1aiXYDCXF4hUSCCIc7uNi3KraIwdCQ9SGTNEompQ5
TXyCvevsRCBR9d3fH74PFqGVzJKItP3gqQj2jfVOG0C/iF8CPYZ3kTiM1vsXW62k
wbcJYexnlph46meCCB5VSJmBnRv0C6A9T9hZ/snmoduSwNrr+6QCWtHIED0SHHDc
fRFC+7kZuS+FfbIas2zRex4oTV+RtgSYWbX5X3DcgFLc2xwTFU0k9gEC0kNYBWxB
5Icwrh86Jwn+38WqgRsgOQdRL6W6t1ugcUkCsUi/RSJbBbUiFCK0FMZa8+OryOII
lZTUJ2Q4ljtNYD79TyqbzMLgjYyD7UONnp325t2ylf6tpfxugwL4/HdePb5r7lR9
egvEsZ/799ShLYLVbUW2Tkg0bJkeqOmk/QdWr0MTbeEz6iMPTzKI6S5EB21pUcwt
jB3x4CxU/wo4cXVMPjaq4uddIfk+ztw/rstxsRxxUV8nXBOgyya6JLFHCFpBeKZG
W2CQOCm43v+hPKMsw23WX2Lh/NQM89YLItojjr5t6eWdwQCBl7J1+dlsM6gNhilc
DBWTFbrPqVh+SopbqsSKH0txJb64FbDz+kScfQfkOJiswcS1lKYNPb5VuVB1h0+P
zhjCINvZWNl+CjkZA22+yPhIWaFwL4Z0Bd9CXso74fvgiYQwAhhTdON0u0lYPUA5
yPoe0lQvBpVNuxJWcV7s+3F9Z1WvvruhDvZ+ap+hH5eKHxMD3DN/Hkcn6VQlNt3K
x1gku6BUxi8RVT6CXf34lzuCuhFgUdOwUtvKjDlS9/yDHmTVKVds3whrOsruubQw
SA6AV9sHKR6rloFsanXYk4oJlPdvp8jXkVXQlQb5wGzGyzf59JJpchc5yObDGSVO
W3ldU0QxCzh8nMR3eT+U9NObm/wwCdgtRX+JJxEvifrDLVr2sbuLomlUkxqcm6pe
NBAAKQF89NjHlJ1W9izPZdt2Z4bT//w3IXyzkog9Z2YPzQiEUe/lT2YDR7RvsZPP
+UCEJPs2rWyBm9VkNKw+25AOebvJTaeN2Uz0eI3fKGVLKt/4E2IOJWS+qFmRQKli
vXE/IiDKg8WhpBmwezFbT8x/OSq2DOh+IZ3SgqbZcCDRiYCQe/jJwtbznTQvWLf0
n1Fw0LsK9PBuazRMLIRxS7xhRt6tvaHUMfqjQOwZtflw/wiCPlOzUBI3EJamVWY5
fhOk5hanR/Z5vlTtboTHsnPZ9pNZAHEQVv7MSZFaOhXRlFRmY/NwDsk5LMBuvR2E
k6A4PVq+XlSEObHt8mMLNd4upHzG+tHd3CMIQM2/n79F5dmNOMjS6hzrWk8VtKiN
pLdQaxCz1pk22VF6zl85Nx75SVTkmXr1vh4bv2kq1ZSB3G+Wp3z/+eNb8xd4cgxt
glhXD7Ezww4psM3re8WBmhB3iMnEXfh4OLtFoa3wVVo0AV+CxQ/OvnQeZmdaGiPI
Jl2Y6nIZDi37/bab+UfTUVKMG0XgZE5DdhYalmhBV1SNcxVjtaVUXXyKrXz6UkPN
EPwZOiEP6oK7oy1qItngSnw0Edxm4iz7kZ/VHR/IljA0dYjBPbUmQlABM9zK4Er7
1+AGGjoND1/+ntO3YTtLVUHScr9Z/5ZsSkqkJCHx63ZneQlcqbR7CMEW8mWOS/D9
0FU2NavsVptaSYamT6Y6Q5xNh5n8OLfKF8jrTkELfWf9w0b1x77y9vXltobquWeF
Vn2iAFs8s31ROGoeMVrVYjyZQWLLNY8ZKge0x9GPiQ0o2gkmUcusF44d6XS1AWmW
VVF3/9RuWvTOPU4+ssTq91OrlJW2zzj6B9OFmxReTkoMnmIep4EGc/M7NywYYW1y
mphjjrGkXeap31fmw1bW/HLdRmzNq7i7J9LsgbVbpuTpa6Kb3pac3NguxzM3Umd4
Zn50kXS0B5iiS52K1i7SxjEmoxC+Oaf97NTLd0SBlYSpNM2lvzilEx7gpqXN/hp5
PunlvDEpSnJZzVKCWoeGbBBjDZQ+DzTsIyxccsSQARclRSeVWtH+JzF00tZ7bbGf
Y+c3DDtm6fb3sgnaV2gr4clB3PG8wbyd2mbI21wS2pv7pFUYhuoh86x66au1Yfvl
/nMadFTeF8OkkbumaTnv9/06WA8DlBD3HrGAeyDOrZOi6IHgVjayMbENcdXqdgFm
0O8TiENyd0i1DDfPzVXu5SMqdmjSDFHQiLLIu9YXcgQNVNu1oGCccvRo4QemqEcP
MBk9a3c6ZQJTQcEBZewgKNjDVrIk9uZY3nW1NKmrw4XuoyALshi71SOn30AydzGo
Pnga7KDq3jUZYXwBzqRX94QsNDhLTcIcwZ8rS6KLBLlG+A/M/F4PnndD7kntvSIJ
fX97Rv0tD4STVUn9U2kq8R4X46kldTvWNLdktB3CGrnlCglVLYjVfM0DWCCr3kwc
7q7wOCOc0B5COif3aXeO21idH/A1tQTH/Qe05Wy9lqMXkySkYsF0W1TuooazttPJ
OfiTemFGmdHCbJfl6snjEyynNK8R0asJEBD9gZddPZ5F5B7zK3m5Qf8DohAfbbVN
bK0B/0cN2dZuWgB0MJHSvCVV999cHA3Dc2gpjSXayA2jQHZ/2IaQOKK0OhtHMx22
pvCJ785R4RPmxBnDo6OARrjKIeCdfdr7Q46Krf6dUcn9Aimds6n0Mj69bzD45/E8
QIdwBh6AIZDXdnzotUEToA9+l6G2xQJkJRIOITdTLFYJWJGiewIglBr23+UWG/qe
GzauDITgs4xGiEwCEXGgUI/q2Ipai0pRQ0rHH+5/OiYN6O0qmjGeDJaejQA7LisI
u1Nsgx3RwUEnTtvlZ83UbkoMIJwq5Qya7VOQKV7dKPuHQmHrEirjbZkAfHgeL4RZ
Ek+ozX4apSI422xjvhxqR/SvwWI7fjHQ83pz3d/MFcF536qg7x/Kgo+hflOP2oU0
q1WfI7oH2Fmrx0uGkS4Ayfq9gGXvQHmS5Trx08uK8h/84JCnSVvfEA+nFJuW4/6s
kTkyU+YFdlBMwugvFjLhDbOv1xraK12E+TTzLMHhr70/4HlRv6TkWc9oI+jmjy6D
l6J7TqsRxv2nJcccIStjE81Ok5+MvJm4o/iwEj0jNbudVqMte19xbXL6cnH73U+N
MPOz+4qKF9VtFwYF8gDmpecLRYFdYqN6JsKzlWoA3Awj4nq9pAl5XSfJHSTcVfXa
qkHL44tKIM25GdzDJiLamq8oVArTCNV5KohnyEFtIdmwaW56GNMKF5YFe4XoBgyE
WLe791FOUjH5/P9d0NRTVTMjo553uDRdK4qffrP23NHd8V0cv6pmW1Po5A+ABFm1
3aNangYGyWL88v3aqLFB83PY3vS4TRGKBrPsUS3hAozLtij3ujpCfrr5e61a2dJH
nCLw2TkQPbjzFkBdE9WSf97/ycXaw0XcMNwotWOyHyZLP3l5Q16gO1BDDhybg4rP
uOq2lpcKM/78M/Ux5IyAKB1cokNFo0+gYNqt+B5LDK+2hy2uZcoL6vvdTyWYNvzC
LLlUDTl3W1h0FHBP405bWpVgDjdcbGiqF8x+Wnanoc5bluE34L2aDgBVgYxb/tGw
wPAmWdFk5Wf3fS5MDcl99OyPLQl7MJHZe3XtD23mLaKggwio6HzyIBJxx6pqQvjH
jRdGBKYxsANGzfG1QlRoSRHxpRc/ytQoNAdCmMiTFYWT5OQHEW71oviKVEhGPWvY
8SVaxa3qvvJgjG4m0MDBzwKLS0XNzQL+0G0FwfY1rXy48rWbz2TAyHa0bQKOv9Nw
8e3bt986b4seNrnn1jPc9Cp6oxU8pqDBGsiYJ6eQmY9CjtQHf/6G2ItlSOkhQ+VC
KEVWwRUkSgcEypZLmBkgaEwtTzF8/8y4VKR4ulcrhx0c1qUqTs4zRdliF6rebnRY
eqeRI1yKS0kZNkA+yle/5HVeFAkMi+INMYbSBH8m5TGbWcR3xeycGzs8pPTXx+2d
AE974SqFJaK+mGzIw9mHrDZV+Dr7r1GFolTqn3EWj8fV32hi3xRZdUTC5AhIKwBj
zVU2t03e0uHk+y0107o0RzLVp9wzt+v65YWAz4WcuEXN5EvRRWrxQ6jt/ucju2KJ
fUXCBO4sCmOwylvgqD4q5L9ZXXR7avEheF+z2CaYrcE+b+q0bqux3P3T3K+bcW4P
1skRZEe8ob4aGMhYunJfSHwH2WyNT6/uul//3uQj6NFwuMo4Nxoa1vcALw3i+saK
Gr49ShUnkOc9zwxrHTytbPtCsjXpjcyiCGtlErhr5pBFIUVLgAGYRQso+Rv5qPlt
fAcMZC3fsDBh5kp8L1cD606SMgCSxQoZKNULyTLpi92XD0vCWqLxTA5OWnYtpbgi
juNbL6PGudvnqNkE5PX4WtZqTqadEbs14Tj9+7D18qoLeZJCahN3OemtGFmJHXT3
D2SfWtLsDr4NO0W2fOVNEaAv6XUKYIFQZWw1WQbW4KGX/xJvFui8md6t+svIpQWs
G9sIdNW2l6iW7FVSSrLaFEvGyJjH7wCfCQdYQrhM/qQxLP5IjcOSmGE6yjPT0EUo
d8dtVqFin+8FpyGiyKfKJ4TrYKFsfq/M52cBJrfWetFIGAijtU/Jcq5u64mTzlHT
GvRLwhLc1y6zpcbLIaDOLxJ2Xfz1OyhlFFM7wPc4gxzeQ6svx0KrmeaLruKFGRl2
2VQBcp7C0+LHDI4e6qSNgXACXn6hs+UN1fDd6zeXDTeDwHEBiKYnnzwH1+/ewxGU
E4q2jgW0tZDfzYpfPhvrSMxqSHrHm8IUbh2fhUZ7mk2AMbxysgt8kh8xldrGV2qE
sO2kOuN9vH1TvhPQJFOYBjpR92Y45JWryEVqANuFxVEnK635WskPDM/WR6zJptdm
ysYIy57mKTBZ1QsKUBhxlHifgPXKQZZafeZ6MOp34KreijvBUIn7dyu3akWd3ryj
DfKleXHMvDEplNeFJPUrAQJNX/2rc+uwQ7wT+G7dcyAQdVTu17p8eOb7dUEY/cJ/
NBHzjYRoKUaL5+UzmABqqlbpDNXZ40fSeXz/3D0UwIzSsoCBjaX6ReV4L1Gf4ELB
MYX+ChivfdwLhsO8zMDKvMtSiLh+B55gMyOly5NJpwAMwp7runPD3oe3DYeZpLKj
wWScWyMnBmh800LqR7DHcFw7sLxg7pi0Gdsu6Hf9cZYiHs5nhRdW2ZBUFw99i3mx
0ovldPq8Py+hWb3i5wFFoEYb+vRiD410mLSngrNttI5OSCLsGdAdEKZ0MBLNd9ge
FOaS97ACmh0G3OklFmtaFpdu6z9808yQ5qyMMbRjd5V567U28mJTyBdpwZBOjjai
aMURngkFXQqw+7m+02t08rgDeYEvw58gzWOB28JgPgceHWaySwx4hgrH0fyFdpRb
mgN3w6PKvT47879u/mZkC/cRkoTCeFE+kS+8twPT0MyAUFVhaidBxH5Bv9Y9xImn
ige2co6/sRUFNvM7xSo3UXx8keMD+RMu2ySVEAtUQxwwEUyfPJ7cB1ZSIi5FVejh
FNRp9uURubs4/mSh7ecUazaili/tv3TgE4P9R26oZFWa+ZVezIxWnhyv9UXoZZUx
NAm7uKdsAlpLlH+6y92Q0Pc4Yew1N3Gy58Wu3ASDXqk9PbHkmQHA1nJYhNdyn+W1
ZaaOepn+8xFOuA0fGNANLt3fPK4mYpf4ooXIZIUcb/dZHW4s/KA2IgvtLcLrIjT4
ryQQFMH8zvq5Fb6AfcJSG5BnY9sKi8pLJRajCjkMB1LKsALXNT/4Je07tBnT2KDP
Vw4FbCzBS/oxYYXQW5l+sHzRoupjGEf6kITDvhFbY893dY3nihVrXjaxBR8vKK38
zfWrFCclP9m2GV5A23xzw8DoWZOlXbncNhV4unn+DAE4/Eeqs4QpwJ2vPqKAgjKq
HlN+3umjWGMAuXG/Wx8aD4/Ik2b5ON1U7zYgcn/CLEyozqkcyPomzYcPXlGGW417
2bfMa0OvI40+BSb1XvvbI8dlQ84KKy2QloXMG0SwJac9NtQU3kEF2uFGxcgkxhkE
my6GLs6fqq5GZJQdpNkNc3OniffrzT4HgOlk11e3sDMNVbXVAbT29Ku1t3vdAWrY
YbBrc/SGxTsuYn3DxBfEPpzQ1/0a3Jd3p3Wd+eHhtQyMzvyXoQRqsDF5UZPXQA3g
8Wg9dKbLYt4djcF0s62Fl2okDHA/w6XE7QjozjVig8hd50edPVlCOQ+fObT19aPj
cL09nTcLVo008UCnrW10hz/vxJocNVizUhPgy8wRos5cdxqH38seig54pA9O1eia
UGxnKAiNl7gyATjINOw9xJ4ANZpe/t/AF03hgLW/G/1HrtKDthkPH+oGVoKG9wBx
Gd96KuqL2Qaq3Fraz5P2ks6QaWcK/orXg0NFLnxvtJCVZCjwd0vXOsRcJwCfDNsE
S3jm6AIb8M4Re+REjU630RQxjSDmbg/ZujDK043mk/1aZWM2gq/iyCNXnZ7WLre8
toPgcnU/JgUjh1Gf183M7mH3hKoZUAUnHR3veyx23yDnn8EzIkASF7mWlXxgy+Pu
glirGmU/Kr+WuqPbOq5BDLyjQpxrK3pQ+Mdwo+cFfA9dnqUEtDr+LbMAYQFyPW8L
MlI2xBSwz5OkcortTVq9U19+pjJ8SS082RLl5qS834yKKE9PA/7iQy3u2OEj7zMl
Da0DcWB45Grsiza7Akep6k5Oda0Z5GOQ4Y0BUWc0Bo+6Jy8R+rqHr9INFtw6VyPb
Yim2WZm3/c/Xc57v+lBp1UATNeWyk+bmQ63PeT5GpBEq2qZkwwJJcRcdMyJOt8au
ZvNOw5ICTH0CELnVfzJDLOOfu6g1sZVZjErEAT3FiIfnSkovRBOGBpC08J8WxSQF
BwB/KXNQWpcdEYqrF3t7c0lPWhTrLbJclZSWpGlXQ7Q81OOISymXUPAC113tMEXe
L8xjo/xmFqYWu8K0Bd10Zdt2erFqWLAEguEN6Gfhj0drBjgtcC07lWicxrTlczml
2RJIAjIOFqBGhXx6P782Wdj7oNcEab1KVaR/+iGak4zJk85zKP8A0uc3/q0VVchy
iwMLMc7l66mefLlkEL/abXwUEKx2ZTTkAHKO8O+wv+EuDfuGMc+iXiQT9nbtJymt
8V2hvnE+9A6Wo+jViqnpBaWvaSAz2IIaDsGA9rGQEK8WfMxZKEZlBwY/blrnlQRV
X/N2m1uvCRehqB8FJA7gYc87/qHTIhCbhBaNO0By7zWasULhu4i1VO1FMro0fnUr
ZHzJz74mT+UwcW2bYBNe6qh3ORwNjO4cZ5nZyQpNvPMIrZk8vivg5C507X2mfRtd
m/2YHF2pcKct/dNwwgn7o+RswtxsJe4iGUCfnaM6KST6aagNc7Lh8V3B47WNfP9+
gjLFuAr920u262Js1/42lOC0LdAH4tmIsS61SKpzWzAqUwmnh+2Giqm/S67In+qN
ZkdEwusH6zVn/7vjJ2i80EcjhpqTQyhFsrWlXwVYYA0qccazv8G/3Yf02dWBgKpH
fRIHh/pSxzlkhgH1ZtWJ5hTVfpyYyAKzxL71gBwY0ehMMUNBOcnI7sJcnKqZShEQ
JonOgKYGIQEtC/w/4k7VIeEliPrQVoMul7Y0IU6nE3jaok/eR0nGk5r4bwdpom7n
SifIz+CTyItvb7PFyTuagH194iWZ2yfS2EB00tHb6BPpLB88jYzDDuM7L+nLMbYN
5SewryVuycmkGw6hXWg6IyIFI0XYNS5WIXVQDN9nOKMYQ81GR3B6MpOhXGs9Wxey
ZuXrNQAxQFHmvKCB0/ELGZT1tOtjFRNEM9xgtPLJ3CB3FgBfy8Al3q7XT3Kib8Td
d7DWZTDb0LdfDLia/KtgPN0pBuSFuVt4KawgKITDzyU06fAypJM7Vt+Fs06vbrsj
9CkN0NbsGeXTOk78DEIMEhMhWUI8fcgno7h32eWsBICWuUQFvmWUdt9Ycx83hqMX
5Ue52MmaAI3j05g9gL1+obvTOrL/aFQSNeIBRdA5QDAZ8LP5TZA8zyS3IEVCe3o/
IDpn6rT3m7z8SfAO8CFbIMr6iZpoTt6/usiimBf11TzAyQiR/ee75ENXrU45R1x/
OnyB+FTS0eKimLnqhwEYlS07vZU4XZLTSrRZPlV9hxrJ7Ibo2aycqlBvuyHQzcP5
Wt2YBwm88ocIKpgwsLgMXOvHidSlIGd4xnealuWjja3IJnUcc/1S1psk9sgXYviL
kV1GmPnTEMfgiXztA0FSq9g9bMH8Lw6oYjyWPOeBoBVZcRwcF542i0/hmL5IQXcX
XzwX8HEIF9hWXiSdDycCDyY568QjBCfara/s7PviSgQtDkHtxX0nxiF23HllcQeZ
2d++IhunSWUVxapn4uUlH+6NAJJJNU+y37KlDd+5V0W5TtPZwNFLEADAFwYxOfQD
rk6Uqsy4E4LB80dnku/NDkTOqw2JWcoUlgrf0QWI9uLA8beGChCji1+PEfI6I+e5
3VyzW+DxxspP4BfHi9fgMIDlRQDsjysDzAAU6Wwt0I6YVqjBYfEx1rknQcaxUthH
bOOM+SuOwH9Uou87BbxkolVoIUM7ytzDucSn5dFIbfO53v5qnmggy3Z17JcnXfGn
XrYASiK/B+RTI7P5FJF1MFBSwpawrOoL3iB3DihV7joC5hQAbXKqNQlGSpnNSbpA
DGzyCAaFGwFdJhFb77j9Yat8YKupdTGnYlTjBK/Qjq2Cbe2wXZjkZ3emMyTNbk4J
5CP0OBrFFS1DjXoJMQpNDBX5E8lBhS6YMrXHuneKfDKgIN+z7xgVR4cdtXuvu8Ug
FPH5YyS6qpqP9YvCcHJG8QxrA0e8Nf30t88jH1QK+iSOX/P5E3Em63/61bUDP1C/
EMI3R64ug4IJ3EPI+hNLDzEvCXqUUJRi1I7eby+K/WlwGPR2FntMtId1GG9tE3tw
+vHWFrjzs4yIqVf0RxdqyWeNK215bzpi8ixiVxZJNczDY9ktbz/aXxP0hIyjfSoP
vyq9aE6Y0VW5h3UGlixixi5YkGn1QmML0A0bG/BXtgAU0C7d56+4xUS3+WqlFBoI
eUx8OBXmWRgmdOGXNABRmt/g84WezM1KSMOFL1sVR6gSVxt2J2umW+eCDUvvMUIk
SYNsKhsoag5tv17Vn6Dz9A3fk+DHopknDD9iUE54UHiYaskpgxbYcSmIFKQtOgn4
rMdfNf2RocupALUHPpH/2/nakFW4453UDd2Un/R9Rk/j7OqCYvHpC9tyozDuMEmp
xJHTY2mJG+BIgsIXW8gRuObtlCcdNXi6n1YnBivD7u+2evOQRHwq29CkJ4Ot7ext
e69mVKaUqXMsCgoqdDlWHBFrcqa/Ph6ng/xsgNfXFfhhnQk2l8+k2e+DkMLeiiHp
HpLd74cGgzTXSOdu9J27O11mUOdT17GF+NxnPS9is47kDganjVIpF4MRwNrwkm3J
BiLOSc5UUZ3JTFSF90H10WDIUwYu+AmlJgcF+dXQt/SuENioUuPGzR2/ZSP2xcjy
6NC7jG484hkHQcJ2miRcYouSoG1QMyUlOrTodsKuAzgAB2lRmDXI8OlvYJnGev67
8WDWpAVr/iD4vX2phiJFCLWfPggHNZieEPqO7jgDrPdSjjJI9FPvkAU89iWTv6Id
qbQIfORtJB3m4+Xx0+DfK/ypM7l3I5ynUflkMt+nbmENGB2BGQFi7gRS9MbWaDWV
K8G+njhPWtK/nN6RY91ACDgbsJcKp9L06+6+GyzQJaXfqVvH+PREBPgxxjVTU32u
wt8C4OlxQzpjEuNxawOB7NjcJGXAzGOtKK9s2NJT7qDy5VH73FjgMrcSslLoL/0c
h0HG9aAsYrHyCuEgiIZpXIZAcip6Co3DBN+LWVpsayGBET9MxxQ38lhRkanmRPEc
GwGze12hZy05EWqA3RFYGnNvrk/dyQaxWlTIR2Y0ExzLJVKdIRau8vTW2RUSxWPn
FErwkOndGLpt6E965nS0+c1ZX7pw8Zjz7uJz+k90PCKzHI0hAY9p+043p4L9rrwr
i828jIGEzhDwcIMca1jOsP2FU3rRfkqYhAsm8LeQys78jRAEbbnwN73/GGbuOy4q
TzjVQ3hV6DGTq4HlSmuna0lRQiry7Qnm7AZhVDjlHcXi9/y5HGwa3Hm9T1YuF5Gz
WCUfFDxr4sizpZ27mei+O75SJS6K7uGfIlysSwR/7Oyhu5N0DmuY9FgZXM2F9xEJ
9+w7UxhFb0cs6zx7zFQLVyqDEwCtlfFA91S6C/WBUUKdX9UZe+2zGfbu5M8u+L3U
ycCFJtZc15TdNI5AamSK40rGvB/G1om5gSF9NP/QdBimbglk9rEOs+JOzVRG9ASo
G0GdgagnTUNyw/XQ11++gsQ4H3D0IzHUvrB24EOlwoaLNqAkjTgv6FmU1DJnKXLc
VnxcBbTts40KCMx31gtV0yHwjrENbZ1TgfNoiRMOP+UARdUzOEyTJ+Rdo9G3odjG
lIiNd9Iwexc7Wx3OF8eywA6T5FuN34yp3W1AcNzN07O7IkMhdvrtdcnm2utnvNWK
99EwIKjfzYP9NNpWrX1D31m+jzF6AjS5VdXwMrJIr95x57v6d/yG2juGPJwIb/oJ
Aw6jEwtngohXd3RmELSWiEzLRqGim1FzuanRrwbbVTOPGHN6tOJ2iEBmfOu3YheB
ZZB+ca4UgpwQ0CfKegTzbOtFv//O9gkqPY5KcvAoSdzqko6jlwzxIHalS/2WD93u
lWtF1OFn7PoE9WXYmx2tcjZiK3hp5zEy2mYu7sVGNq4VNW2yD8/1Gqv44D3uYmY9
SRec4HGUF528v3vCcDsIY20eV+7txLfVkZgJExIcpPq+gYLd+fAHz+qEheY21NUL
EGOMQIQaTEvx670TX+6a/s4bpuaASgDi6ReFAPJanCtsOAR4c6owgktEQ6nAympz
DUoKWAFkbD7jkDfv51majNbGhaRw+CPNSIA8oVz8mG5K1KzNVPDyCRYSAkmvTSqP
UsL/PKYlTVHLYiiUkO+4e6xpAJZSfdi+nFMp+nPco0uZgIxAQHV/hDrwI8+7gclE
tGCnrHqdyuGLnEpd2iqNKFFhxIQgUuQGBfmtRAaxABifp3j9N0PIdFMDRKRkIchc
SEAUbgBrs4zXFfcOfQ/TgZ/tQv4FX8pg0WwHhHx0QDFopsUb1SoFW2eVP41Tjgzb
etkfQUVFKGJsYNvlctNWL9JaTCkHYnTnczzORcM1JbDhtC8h3dG2pFqJymp9qcHZ
GK+KyQQurKaizeZGlvUSQU5d/hqFAmuDHa5mkvuWaKeDDR5TuB4Iqf7g1JVcVjLz
4Pat/0bbU3UKpuXtScKHXjNXVhN4ILWLCVgNdni5JnVOxtAIjSPCGVcUB8XSneVQ
zGn1wLo75vQ5/oRhECpVHvEVf5fAKNfHBf50o9DfrzF0ccGFIccuTinzt/Agev2O
NCa0UQMx/MOOtXLmMdKPUOk6wr7mj/Wp4a6D8ol4vXBZ4U2dvRjewxXgHb/23k9E
sKni0hzhOrvLcLbyK4BE+J/T+w2OUst7FKMFMYFOIXZ2IVDuAv8VDXz8t9KQDhEW
iQq0Zxh0nEJrSRV+pxn4ZE7cz5FjjJar0Ll92gr0033xaK8lrN7tDO5h60WRgKXv
I4tCCIi3r0EsEk35RLJ6RcDWsnXjRMh66fLwXzb3Oa74yiVYN3iMrWJD3irdM7Lp
34FWijZZDYiU9aSy8Fx2W1uGzz7DLspBzGb3cWDm6l/b0qoBba1PXHtkuRUvRzWv
sUeNj+ch2GWETnb8Vk7aIyxpCCvVMMS6qMtWt9c2LlgbonKN/XKMcGHhtlAIHHJm
fU+XeE2vbqCXsJdEirjEv3gS9WZ391eRzhMmNwOU8NFGIWbPaSmH5FPtT+2Wxkk9
kmCjJv4n5ifUSRakkMKCHXZ1QqyNoJmQQ7LD3NANk3aEfX/3wmW8s4/M72u61Q8P
RMpclLoCqSvWKrXmJffsy9fNvWtnG6+hBxjo94Vj2bpor1oWrR76J/lTlFunW7RL
3WLhQ5+teMI1HmAawj6+zO4lr+lbX1XUGV0SHyC1+Q/tKz7dDjQnXnRqsU4KeHHK
pqnBbmyV0HEdY4xjgg1BDZOsnreXN1aVCFoC/rogf/QFGlEOYGnMxwnStWjvVetq
aCs1fCLItAaY4qL6v/wHUXW4kopmjhBSvc1vD61OUXUsz9zLzaLFLP0gTIV3iu/U
WVk4l3S13Tw9qT+WZ9Rncnwau6XmGPi8eyIsc6oREoA0R+wNsf5Ha2+7PjyW6GIr
jH1fXa/UDlHQDvIb4/Yqg5czT5qKXWWAX4Wx7y+TFaZFzXoGx5RnWbdL9kPVPOMu
rVTT67BxcizjG/+4TCTDi2/Tgmv848EjZf9hSqj05wQKqbptQ8uqlpKzNp1W5XN0
Rxoe3lrKv9eCQyGRwvyqOA4qO8zNe2t3uOPP375yhkg4K6P2YjBgYDUuntLKIiwo
i6RydiUs+qNuvYDbgP63w9LizjSsOcpVo9sQnmPgBfqt/+LOFioLDzh8fr+JAMlg
R6b4vCZSZDl6xsVPT+/3cO0JYXKtYiztxajrakdaKui8MzU9nRCyx9GPUzWcc3i9
MMFiQ06y0+TkOGxbrZpNOMLp/FhEHqJB9HGqWhcN4vXxHLUVDZqZRTg8lEzcItju
mHLuwXDeZjtAJgn/c50W1vKSmr4pAhRmGZ/bUf6rrAzf79u+1hUUdgqjoB5eh+5W
ORDJ0ekKkHl8rSd/Kux2kcEclJM+flk5BcHN34TuBfVqhYgWHzYuZ04QQ6EPQCQv
WdjFeNB9rMuXhr5mTVDeAGrcJbev36ySs9e4tgITzsIYf/GTwFTu9LyZ7qIdBxQs
B+pBQTreXwjZZOXeiL28sxTrl4v0UKTy75Ia3mglxFY4XFX+P37Rzyr3YM4MRAZt
gsYQg0Au/BWx2GEUuiV4RTzYDVTLT5t7JyaaSxwrD+e1q4WgRjFcpm4sf1pGgzk9
EZV0XhKgmpXma0RCZZmYYD11ZCcFv1nsfHlmfQ/MHd7aZFkL2h5cfWp6749CCx5M
Y86xXHnNlaAD9xFi1cxR5RT9fNJ3EzjTlT/1k6WfNJP6FqqhnuClUmnq+2cDV889
s8eH6B8qbMt3zNrkJJ4I5S+wgsxhveqYaxMnjwC2ErPGNLm7M56OwcaIYZBIr2kC
QC0XnJ3OyLjlYNxSrg8/u3yT73K1imhbuwANydv066oxbmtLYg3IjGzpyG4/ouIL
Km7L4sEC3yRF8mq1SFwZ0U01vhGp6v2bM2ci0sd7YPlXUDyaw9bgx90kygypxWOl
2KrQc1sanGaYaVBxjlX+GxnFxqXUXBzVpx15JjaWJR/TZ6gwjykHof6GjmhDu9wH
qG4JsI49kubOlM43+Ct9rfMziT5ucUW3g7OFOGMnYO8dw1B+j3EZQnmY6iCUKqUf
qUJSBVZJ8wdyhj1h1PJ5UGp9MCk3bJFuFR1ckLbMhjF1Fn8ILgux0aLTNZf7EyQg
69Zz90he9NUvnOnxBgIn694hFVvd8DhdcrFsCti1iWtTo6/2DbI83k3evQfnvt/t
oEsb67vqeOo+mG6xVwlW2YB0sE3Fp7UU+8MFva4nhpqmt2OmaWzjBTNZhaKmfQ63
SQxtazWxGY41ud4MlWihh5bwq58wGQbP863j6SJCoQXqGMXcjEY6LWO6Fa8SRi53
guu2fbXgZI8NvSA2ZL/fVMqy4j/CijZRXFlqyrFlCFgXB2/Wt9RfbhBu2uIKvUMo
iQw7gKtMko5qvBNTMI6cHYzNnLpjznNVwSuw3BgQvlCPfggsaom8zmQfaZnkSS7X
FhJVbespVqDWJC36NfxVGA8tISvo98rLmjnXD1/M9Ehypg393ddf4VGOxr7VLxxa
jBWr+MZW01M/DchkVoF4WkIaCdrB7g7cju5WPkqZLW815PX1RTqqzYkii4EI7a9A
6MPfLpj8h35OOJzY/NcTG42w3ysofvjRB1n+BfK9aGBqGrtmdrSE9gN1mttwogPU
KEnJVkklqlYi7S+hKmCCGkeULl+04Tp89bpv9WVXnohukiN76Ha3zeaHLQfpdjyk
s7Vva2J5D9BQwE1bQoHS3F07P1blQm6y3pEnJANvw0CIPEjgf+J/PH4VOKf39QmA
mQeLRIu0snr7ZFEZRETC/vlvJSkYU9VeJ3rqg2YDmyTcDyOTo2wt7Km6hYC+EkZT
h139XmDC8zWKfz6E/PdIfiZVHlE9K2oEratBssP1o4wZak/5i0WEq+qbMJE7VTNV
pjxqz2e5LMj9SySQBMvYd8Ltt/SW+fs7mC1PxumgozhRFn/VG2wGlYEsWHQCeBkP
xzFyPALSOpxQ7WFfmt591/qy2Ed7ia9HIqbz525AmjcqHVP/ZTMNp9SrBKeEgf5M
NqTRIVvih5UaXe+UrWEpFfcklOpmk+qnbplMk99pLJu52FEWcAkVpCg7Zh0IVr7+
PLzuoVFxEzZT2Ze9Msf5KAJUNzDQNGvrqP5t0u6VSusShTsSxdDZLEq7fENshfmF
NhLHJXCdJoeZ9mhM7w1XUOOeyt2utAu6ikvE0WOIeTZUNsXbov6oe0zUs8yDP6uc
aXgMqWo+2iQQJj+cy7ztFQAjAVmQgYhyyIiS0iGNXycFbvEWGPDMlcyjDsjyGdl7
XXNEa60avX7eqJ5CYfdaFKm78qsgJgunETreKl0cWLffVQ4C8UAQt2yksLOHc4B9
loRXyJB1pCxSQTEASezW81OwQZJVPE0wWP6Y5Iq+g6LFnhzrd1odB/N+46Z/zeVf
WDmq1HbKWr5gXHomGO/NgCCoX+xN/X90Fu9ZjdlQ++xrGO4izBn8ymqUgSGmMrV5
21HhcZYvRmAGIeZ4yqGHQOInnPUlBoJXQ5scXFZH33jvXQcR6o6QXqiAJR6UZTxK
vhQa1ThJgcqcO+tbRO/SpjUFNMwXvzWysvKwL+z+hAR0AQCWwG0wzm8qbz0nLbIB
vPdMkkhZpTmn/FJeRMTfW3TUp7EpIL0ge+N0TP9XllSc1c+/nEReznN5av0rrZNm
DQaf3Si3RB0g5LarJYmgJc/ZqTsg+Sr7RwPAZPCmNahTku1/xxn6Y0bc0SA5y3vT
cA+XZxFZUR2JgltNDZsVwtz19srC72kra8OKLqDFPsGsOQfOND32uK09iI4NYm3G
SUoBkD+H1pLkO+VmbczS5/EaSO2ng2uxZmZEJZ9TNKTfBd/0OiSsly+ocuSDr72C
fVCwOadDOlzuxKH9TOonBMSZG6MezRCCJw1SE2fsh5RFhAYCNakLlZNo6rAAc4OX
biaOUwB6RNSIfJNP3KawUwWj2lxpqUMb4ZhcNBvHqVXVyPg5CIRHM2ffdV9C6e6H
tFbyTlE7d6LYqfWM7qjNmd0pZPGXsBccwYTlveev3GTuvlukcsq2dVS3ubVSFRzk
ur88wPAg+9rKtLgU5C2m7wjcC+ycZmFe5I75jZp8BjsCMhVqkySmVBLbud+X/b31
QaWHDOSM54lGUpH6cQLFjzxAotY8N4NvoYGZrZrVgv09EYSp76aY/UXSHS0YB00Q
Ce62XAauMhJx2o/DVKGPGbU8XhVnuD+dXQzQfN/gk3NO1b2sZ0bja1EgyCm3a9jc
iGneOZXQ14b6uWZ807lQneOyvDeAQAUVykbcfsGHSG+M8UHkJs2sfQnKvigXhzIi
E3fT+FiM4/TLBX+9NzzO3/u7bAZh235TsvEweRwue700V+mLWlqJfB8Z0AAMOrao
DVDitAb7PD9JaHH90LzE5b0yr10ZBxYk4Eb6WCoeHly5U6q43odPD9dZboJg0UMR
/UGSqJeA3/MRbjXmC2ctQo54J58P3E5qMJmpEyrOP6+M6QneuB6Nd1EuSaUco3Uv
saDaFAF/RzyxcQD4J8jMqQfEO1WC2YHrDO/qz+PNng4wtpTOxooxPw0m34i9S5HH
ZdCRTN+ualIJb71nEq9Z30tzrIiWAWsp+IGPIT/qR1Q2D0q9Y8+hKbCir1CIpD86
Jy9Ll+WYg1GXSSLoQglRoH6dsGPyNhPjVaJWMa8GWYV/tQC/b8AjMRlZYmOZXogP
uvpGu41NcyPQasKw+8a4YNhYjQDU3ySSn3o4MHdU0yEj42+3PQKy747dyCKMHKXV
g7voYFYjy9xRJxptgx5X3d04pw06tKLS5vcwZVKUmo5pywTWuPdYKpP+/mh1vlWz
P1NKDozQSTADQT6sIjFgYDhJ9ag/2Dw1mY+84N6L0ExbK3ALy122hxROVqVvC4Qs
hnnLfWStdWrI+R5tB1plxiFJobZ7PZtpmaBLIwDPsITbCosvRbIcO4mmJsFWNI6d
CcV7gD6TLE34Ugz9l2m3eDsJGJy3PbT/k3pY1a5SnUOvlyihCUfHMnbfUzz6Mvmj
opStvmRKkmMW36PLtMQQWJ0i53AfdrkSOR8rqAzQ5wwhNY2AaJJRb2WPit9KIsSt
DT5f7WuvbD9FF+B+VQkMgDHZyy1puzjckEPudUIePXrRYSUf7kSi9ihq5yKuQgbV
vYbgmO10w/GMzfGd750lbhxxykBzAsPNTcULZD8wMCaSEaZRPpr69617awVzn3Ti
jqFynSN1FRagkNC0bBvEDNj+GUH45tezqbpSzslbevEdCQB7WRjzm97ubgGFt+2s
OCWC5yYB6z6AYRSlKgo08CYlsMw4QSJT4D0NpkG6ucU8KgGoY7fDGwBag5KqnG2x
HKS7fLrJLNCb7BOWd9bT+CpYldFFxn0BQTbJtZjokO5KP+3atFFiaulyPoZA1DHo
T2NECCzVnt+KhWKo2FDnDmrP2rWR2/3ivUgRlqHtBDEmzPWZES1vgJA4EEOliOPj
Waoc/MY4n64YdtudMgLMBzHfHow+VhhaNcD1Ld8SU0rjZUoVs1pb9fiQndxeRc/C
j9AqqNz0KLc6n9AIr2z0WW6ISAPjiM6VafAJ8YtcpB5m8VdePiY7Oqvvf4i5OqVU
cgV80PnB7uzXe39vH4f6Lp5Huew/yGit3LFaLdOiKEzk3kNI8CC6Ezondi919WRB
rSErvh08EtPJjlsdk6YiNsiwtVwsvYnaSO2cBY/VOZAz/UwuQPzDy0n6Z3x61tEQ
NKoAE451wo8vz3LyrOPoCYJ5fNZ1xSXtKBWC7k9tOXzq2W0eZ68BgjSuTsZaONci
e38a4lb0gwqJUK3XHrAqc7TlXhFi2YpOcKrknIAst1YjCeiOz+kktmesEGPsYLAA
Go7+ueuJUt3In8ovdd0b1SQUbdlwN/d+0LrfR6V0IaqByzrkDVAYHfxNyPx4gZqm
K2shaBWBcZaJtvjK+8qKgY5pdK+X1fMs2TeLwDKctz/do5c5Lv7MW0eSdor/Wa/Z
K6fgmbfxvJevNyvO9W8R2YK3zN9lYl/xnaX/yxsfxI1kPcK3kqsiGzTlU0mnpW32
vaKiIBomeD/vkNvA5a03FY5ajW4XRXxTmAlaxY34HpGYeoEa4ZaJh6/uJo9rV7Dk
Rm+H+AcKqm6xSuQid6tkgPcWhVag8YHijhhM71/fZ+1UPd3+uk/XbS1i8BQfQRyZ
/gsM2UFe8Eiyv0oT/3gahnD/4DlAXFG7XXgvcQx+K8QDAbwLRgkGMUXHVG0edHxU
cttC+cTL59X3qy9uTS84r+pfsljF+JVWLj1W3/1QHMqTeEGzP7mwrmYtPDk5n4o7
9Vp27X/3ZGMl4DfIUu0hYlA0k3AP6UlBcSqUnniWAIZQbmWqw2iZBwOUyv3ZMqFO
70DU+0J9/I9M0gwNRFJ+9yJZr76/oTt0jri8YNP1mlFEwSpC3UVWFSUe3J/eY9dO
t6NoiEMufEDWwSHsnZ50/ID0XM1nRdgfC089OkIMV4w0iNyEm9xKuvI5p7b949D8
ea9wqxo+C5ucT0qMZL/FGmt/ZLgQeTLB2p47xnX37dLZrDf99xya7HGzHWBLkZKH
6M10PjXJu43SQBZV0ekAMDt70//L0Uf+O4K731y2vWeDaahRX7Zc44U02DOGE6gB
qNO5Fc9RS1DaduB7SYQjA2eCnTp0soT29fqi4urMkMdupOP3w8+P651VxN0qKZlt
Pa5azbaPpjPk6uNewsEnrNgWTczFUce6bKE3DjYAAnTPuGORusFkF0rwRcI3441M
MfRjrBZQu/l9uy4avjHesKJ5GhqpA7zgkFK6vg8ALDm+w6R+dQlS0gVG3EK3QAoN
EkM5v1JArjKwOElGNdjorwfXOdRf0AgrJCm2ynslnsNrZmL3CR9sULfUo6kNqzB6
wmQndQajB+GQeq5+ue6k9I2/UYr+Ym3K6McoavhcykWTZgehnpAQs5nI80HMkj9N
1Y/b5emOZELeGPTGkELe/AqrU4VhxxQppSqfHQFJEENJ8dYcpmk91iP+nMp9TUWV
WbFbDixdcKUmmDNsjqw3zYituxvm/tYmRozz9CA0dpqfc8SDTXkr1OpDJOA2AY/G
sioNFx5X8r5OJipHCBle8f/M0I0SHdl8cHlk3L6DGBKFGlR1QSq+cAKe2LQMctQ7
w55V373Fjccr9RFKUXF/Q9SEtct/Q1FiGjKjT4gFFc3nn34IMSQAASJGrpown5wx
3ux81D0RAXFfKp/22CjBm+HVz1qN6pL4TOdc/GeioiPNm7EOBA+YMslgZcjLIPCZ
jHnZDAj2C4Pz9jIoK7wuoX7z6p+q/rKSIzzMTrDsszm5qkwZnJPeCXh+6tL8BEMg
HEBdvBdoG8kKyuYuYHIjGUCYnT+Fe7XXatkHByBM53LSS/51lVZjuEb/c03hWEEl
0JrXyvmbbFVjuWGoD+sNrIRAw00i0WxDjlq+aVuJkBD/2kextdpL4dEhQqZGC7E4
4KT5ussjYtm9A+idm/ZfbiknFMCQEayeYTaBZ3sDEMMp1ll0csC24k+R+Ea+DPHb
J3X80BpcULvBw45u8KlqtQBBPe2AhbA89WkdsKssU8WzIKQNElzsfaV0Ufixtu41
Kmi8pwSApXs56aNDMo+FoaB2l0glmXRAqtr99ivwIqg4NEKcjOF9QitU7XIte0G7
uigmvTkKZjCvyan5AhmfLpObmySZxvhtV2jUtXGi7EaMyffetFDj02SC3TI+W1M6
Q/wevtFtqz+HELR3BDuK5G2vJ2JfsJAWXAbo73VLZF/I46WHsSm07dT5Dgw+qCpr
mjKt7Su/Bo+tB8UPqLuxA1B6nkafFY6lnnM7ty09Ydxg/FOUHRxlZCVHwv6WbnA8
OMa4RiS60YcLSEUzt1WP/48rkFIM2LOt5CPXGjOpng6viuIhQz+tfJIShLHKR8BT
Z9gT8z6e2DTml8/DWdc1eDtfQpEAQRrxEzeCVlbWnwulb7d5stMHGYMjnCeNF3ud
9LgCDHj3378rpxVXRV9JC3FnpX0ItqkQwHgocdF9kaqi/sO6h3cVQYnRkK8VnO33
p0LQJL1FhJSTSfezX+Xqv4W8/JHn826X4c1q2IMV8QXEChrdAUygBet+IOBIwOYY
/QNLh+ktGevpieNRcCzy5iZct5+C1tZBVz10uFQowvkOg8SpksBtXDg39GAcX+eC
HNBCQ0u+C1G4FqDVY1RjmxZta9ugGsnUHf6cBC0r/uukPw0OWplkLuHHfIEJypi/
C8yBacAMt1kpKud7wMV8+StzONtMypDOrnGUpgxOF2lsR7yurQsYk+FpNEDhlVo+
QM410R6MJ9brBRjj4gbh1LmTdZ8tJi9F+w+RSuKZzEqzUJ1ACHxGvnDmHbk0mkDf
+Fctt67B4VLrLdqSCIZrW0C3zjhxZ2zlHgxsn1W5yidJjJkmZBZmiTEu5CyU50mL
4xU2oF8bWiGeRjM3JJNVCtAakQAbf/ysRtaoeITP36gtY6hkJm8otayzAMY5c/QP
Gc7ZZT6XfqipJe3+/AxqitsakdrlU3qOLR0bDS5trkh+jjBjqSDkNrYIRiP2/jA3
f999kfAp/MZIVF5fBgTmEro+PLc7KOM97GnfXXnCtfdnIKtSdJ/5qCpcrPp/T6MV
MlmE0OuFFUFxUm3Tg6PnzYHIMST8plBXBKOXUSt9BqCMve6Wfa/kDUMBbekoQhjT
Z/8E9WiQ1L5cIeF5WllYuC6E03Tn7XDWX5Phw3CCP6QyIJ52C7edRO2cTb42sTix
HoDBTVWYrnpsyXh8UA0IquUoQ8PYkZn4nVE/mr82hkuzJ4Rsx7bWo7sWhooaQRTv
O7fqZtS1/NCAp1ge83HPT0qhSJ6MyNgfdvy8lwmYzU2WIAeAYPocgfjBlPFMr3y6
iV/NG2glfXxoVn5iXpYVKPLZ/OqUb2QT3fyy3TZy4PRMKAvc9F68GEQGD3kZoOPs
QS2z6ERh9XCtZctwewo4O02F+V1qRGW4Bj0EpyTzs1wOYcECcvoZKjmmWU9hqWGL
bRV77E/b0p01oz79qG19qC5nIGin8fYEHxfPSfLp8/bcETByH65aCMtnnmlQv/po
b9cRndRRnyLNhthwAwuLxpE+rnQLF1RWPRIArdvw52Sk4tvAYtJNmynNA6APxETx
PTN8ESdLia0Kaf7ytU0hsx0tS0NkUGDa7YQkdQZmkleNBnau75rEEClFFyai1NKN
Xm/CFcqmuOy4bSsIXF/aCQCcKK27V9HhApUxrMC4ioyjQ3gJh9K8oOtHeso9iKMQ
BiWpW1U4uiPNYtZVcC54jelFo07+0/nW8njB1Iiz/1USSbDt2S1ms3I3R0VuM9EO
2m8DfZjzv/TNZ+J8jIKVv/RbKM2kCEgeoQCYp+SQGwWkScPXMKWUO/eOREnaqDoc
WNZoHF5ZmuVkruUGsPdDDw4lU0YyAnwueZ/72LlS1TR5TtiHqSNjOgv3Ohawp038
h1C/KKeDN6t5MVvAR0eQN+WwP5aHjcOX+/EQrNwmRGRv1uCzuFOt/VXUZo+b4v5U
N52ROBVe0H1nbYNOSzDXo1KwILiiPqgQqlQbK9B7VOgH02kAK+DSvWPoX79FRqk0
LqrwIozxVnSL0WNcA7N/aasqA6xNFYQ0VrVgmTosd2YNCTd0AhM6BSsNN50eAnmN
s1N5RZQL/bNlPkYMiQlEBfiH5LiMXVHcY7jhaiCG+aI9hNLF8S1mcDF5iAJfGmd+
KDZC0rUdtZfVJ/q2UA7hpWgk6fg4f0lYC/Pe3I5/jjgL68h10rg1Eg3tsG2owuu0
i6Ecm3+xDs/HHxfBgFZezHUxPGvZsfdxmDcLu4Fx6PzViwEp5jIIvrWraeZRCtCM
XObtjmt8rRtHKvs0Grp3vjZnKxv4B04nx0mveFC01d/bxYxRlkjEdoYC1HI2mAxd
1UJqCeLn8N0e8O1cSge4JuH8RCkHQcsbIIpzzCMbw0X57IAAyVuwflZinNM1h/2Z
djkmdSMRGx9dbt0U803O5XE45imCB/HbjjLMocrvOOzXEfNF+1/Y/oWTlXTpyOxU
itvcIhYdA/NjnA/eeQ5C2SWRvl0AODFIi1UF5GRG3VwBJ4m/TAyAxTZ4piPc3nDh
/IumEs4g09XhK6IzkJCvAI/Uzir5M6tbxbj3sRCD6seYC03D5n4j/6KkM5ogIlRC
/i9OizFXCOLKIUsi69QAVhCETwZlzCiycpZNPzcVpaA7sJEoIVzhUP3PZ2eyy/le
N+iQP2aZn/s1JCDJqSQkABZGGBDzRvXU9aQdC2eAYEWzfS341Vo7QwzLKCFPNcOz
dHuadI3E+Wh1owNMF67kelHugEmkN9iTace2BqQZ9HeWxsrp655xhe225RiXAkMm
OFLprsCL/tcFr4DpX36tCb/p+ADBl0tsZqJJZ2sI8OLZQRGGLJOmF0SXGMt3hgxY
j0DUXEqLI1Er2okBsZ8APi6bM/BzW+bk9qoXI2jSLno07Z6WQJhhWeNGHPVxLhOy
YGB69teVpQmlBbTG1/4eSKnJTLQMm9wyra0y8K4b3e9Wbpn7laQ2KtYTkKyuXAnM
coHHwfroqFzripumQ7x5cXpvw2wHhHQ2QuA6fwHMxJDDRdk1YYqdQ2fmQJwhUjXx
FguYVIijBty/CjRbsMMuDJ2+oQSeAVgL5ZNL9fwhcF00iMnAP8xfDE183qejbonb
ZOtevyquS4yZG0z4ztYPNM7jYtPbKpqDN9F+QIYyNwi2dZrskCzXU8w/vfTplLgJ
/DY2Hz0TyVA3csaoXF4HBcCgtdz5SNbjI+mJYSgIRpicZ+tAXFSBf4Pv22J63+O2
OABTbV4Aj/jwgER3jmK5w7mA4K3MQBd9Wr2YxnmKVuYmnEGV4cMCUqdgCDIWrnij
Kq2W8PZ/jxGBTL3nF5Qw0OC2JcFHrhdRdO6DJ6/QG5KGEl6Uxc4aklrB8xcejrY6
NMnhMW8AaR1SCGYF8r38yiq9mZmVyTOUk2/YZGkW6dtAUm6mnRQzU4V13h2Epn9J
diHus0xqWDWNM7Zw5GM1e/5SXqeglVDhpiFWNx3gdKgjuH8F8TwbwneAXZenU4g5
AK29EDZ8295TO6JhGgBtDb5j38ITMQ+7CHth31AM34BBatRhcbHbLMi1vmVYjbJY
8IQTnuCTwy2tNwbpAwQfqBz78cfLhn8gU5hhDI8oGEwhTTugvWJPVWZKIw5/x812
dApN7puSnKMUJDj5KMmJRR1WHlwdH3xm2liRQ9xd+ZFiRCv7RumQe4lSr21hBOwV
QoC4LXT6/sI9hPW2SUTGrKM0ziFRWfl8AukVjP9wQrcXtLtgKem1PLQJdv1WVEHK
fuPYjwpVHrhivLIRG6pAN6UcZGPK4CByraYqPZXgzY88Dc17iOV+dSWSw1h7aYvV
wBsJa8opo2KFFwB8ji5RPmiGkIg8nMiEt3uz2OcXt/EnlpJsdAOVPL3FwtUvBXqm
jLTE2UE+hiU0gKWD13+C3wVGSV35oBW3b5zuXUXApOYpSmI7cXWC/Ed0gJa3nh4/
Bk97t3gqYOoPd8sGwgpDPWd+k2M7Q4TiU5S8kGC8ndfAxKIfoMSd2a5C2JbnrUkj
IS2TxGEFaOYR26heKjf6AT7eUB/+UAFdnrl+5Vbhexj9A7K+OB03VhV0pJJ6sWEg
/k/UDQK7FRDaDzt0e1wfI4Cc8oZJKbSO+2SNfm8N/wY4/EurTGiAI0GbXuhYjCF+
/bXwC6eozGBfB5hH6fn6fytl/gZY6sWT3TwmOWI4JBuuNrXLT7FPx45+AArWMHa7
AZf3Wugqk7OrHD4pwZalshZyYMh90tUIxjXeFmcFMK9iyuTOStCw/UDg4qkHiyzx
DLCvSlV3Rvhhq7akw4t690I2675Fwkj3QsBmKtmr4oXkzmQ6L6qsMj2kUCCtkDuy
ddbYz1QFJBPhusY41r3Atu1mHqPcR9CiDqa1t1Dl/weCdJ4j7y5EfMen0lGpFcu/
76iaX6Z7IclXZhBBfuRrsTJbon/cPfunK43XISDvTlSgG3aZhiKvDnZnTq8RyjbZ
Q0a0o/ybdRE/ehgRZZmssHuywwbF8jFc/0fc93UrblC8U8EMiswZ2i+NaxMHD4oK
7Cv7tNJNc1VVfxcFLCZ0qGQv8VSSZrc52l54PmTCALwxzUZH4dvVkLENFODJYk3S
oOXsU4Z3IZn8YRpL6S9PRmIbB+mq4oxLxMng/Lc7wZWnUOFGMhmf93HD7X3Kqhqc
RqFZ3ug79XHLlhwgk3NxWJFjDnq+eD1w+gbRGcs1fq/kO86Stuomeg6dngyPHARw
Lr+af1PgH/D7chvhIdpHSHfZJjqoQ8KWE5e9WFf1afwaY1sCwpsMkehu4Qf0jaZV
yRwwaYUjJRZrUKJS7ywolq6AmmtfRE33WBX9j+bgqqk6/mSWyFE1Nc8sEMB3qIDC
wf7Ivq0eowZYl97AUc9c+QvEr2BzFeBZEIm8MlgA5O/eV0Ftoffpb4nUxPL5jzSJ
XZn/ZqAR8A35At8wn9IuuQyWSribFEgUISSvizl5UMTsG4NmjU4wfgX+q4dbEcMe
w5BnXdE+cE2JsSpGPqIJhZ+O0uF3P6e+Mg/sk4/blSwP5/ddEXImw37P/f4eZw0U
1HTdPe+Abp4eMLxsKV61koNg0dv50p2cRDtjeK2WUQlHYNckL1BA9LDDDWLPa1rm
Fv4sDhMBgZwsBHozzzKAMmebhSCg62Hah7xiSUAaW42wGXhgAN2MUrjBzL2SqcAZ
FhDoVbTvgaen1jOzn2Xhzw0vBmCzNWVhM0lqedSMsVUZIBv4EBPZisJoVZoRxIik
9O8yO79EsGMKE38T2YSg0CT3CYw/PUgDawKpgQq/3ofR9cp+06zWWZLKwAY50/WJ
ktLsR8GphyRx0eiic5pINlDwUfOuc9XG/l9VyAdztEq6Crk3we6RZ8fwx0oWEyR6
RK4Gfs9M/JoM/tpEpq4CDYW8JyZSuU/DLCeFv5K6/wf9sCpKOytGUbE2pS51HVZ0
s2gsCKyEcOLQb40Rqu3ycwTQK5iSk+3w+37C26PAX0D96MN3YHpKJTxjEARZBgJf
RR8hELOHqIbMUnNcH4ARvM0LRPDr/JcTvVUpZxxeGrdo8ZkwhuEwMWxs4tEbItyv
oQASxMgg0813kzbOw6fZhynDKqV0GcKprDe15gjY3Qx6k5UyzsxVnLf54VNgtIdN
khgrbEhgxWIMg/MgEWn0ME2dg0k3IYtwwlJgbpvN1LcJZhS+3b9xCQJd22uKZgAV
apBc60P5NsTWE4Kx5BWQOmHNXbAMsHDiwyzcm/yVzXhVzr0JQT8TtYi94Gje7i0W
COxJCH2w/SvBRBRXjkuPZ1rTtE/3r1BFYIWIp0hajFgrIwCIgbDA+xgg5Mm/whBt
88VTHZ7CWZv3c4XA9VcVuZg53tK6m6l71pHGaxyoKhPa0Iw3iX2O8lMM8O35svEL
jbLmuvu9wyZtKtJz2W+LSIhWBUXnPCrX9Uel/oKbMzvW1/Y542x0LKiqoke05EbF
TFKwM1JB8nTdVDenpFG6DCdTAuCCnHkHmH4yfZ1F+KJqSZ927RPCPYtcE+BaQeJA
ggZe8FGos4XwSWrqTi6Kl2fVr3dW3pQ3HQTl6NWYLvFuHETNUR25Zy7Lezb/ZSnl
Y/ncjOyB3HAHVAKfs1Y8QKC1Kbjyx8NT0fWgGzLEBjPdG6c2le+2ACZS7g96hFDP
gXQIcjPV2+CHv66E8I/dI/7m0rDOI1Z5jy6qHjsZE8q0AdULAO/aywSZpdMzBI11
J3UUi8DvnDarQqZm4Fo4NWloNJbSZxEj3cOfps5doJ2BEnv87jFDTTNI9zn+L3tq
2mB73iniySSpDhEbL1bwCBzkk6kCnP3CgSdEkkGvmnWBVDewhbMNloLmDvlJ+T46
74FEMgpOI3fyLqGY5uMeV6avZCoy0Qa86sbI4HnW3xfAu8weP4e/o+BPTSW1B/vv
IQyRnxTsaKDavBlwpd6o+jgUtyxaF3UqJDqdpfnDjGIbwh32taoWA3hc6dKmAlUY
BRYV8hcyWcUK8vjILE8ADGmmNx7vGSeNFAuaFhiOq3NocyLq7eiNk2U5hXUBZlL5
t753Mpz3AHDQbw1Flw+Ik2N6BPPjSwTV6kZAVIo/kQ5JRhqT5hvRLhlLoPJoH6Mt
CjyealoUjcS1Hpq+3EEoxWcmdBLYi9u4+HFf4sFtJzefG04GXHghMKuueX12uU8G
phuTsPVu3yJl/e2bo/3phj/xU9GakP5+44u2bm26Vh3bS5U38DHk3LpMzwHDlPw7
qmv1ohfMRq7xvkyUD7ixrv0xY+gRcx3VSXk1pegl9UsOci0zEON4uIW1M6ZbTuwm
DMapGltiI8zOK/emY9MpmkFzgSz4sbgtD4OwJBTzcHi+nNJq9m8PCN3kI/dSqOpy
H3fjnzTRwsQ0uPw+TYIguaY4llqys5WPVvBqe0BQkzd0HW/Fhfs2aEiwgpPVTEhi
0HeLO6wLXL7lFmryVQa48M2/jPoi0R/IxNlIZxuelwRAcSAhngtZ6upTGEyDN4Mt
A9CgTqqy8MO7wYSXj9AxbBlFCa9OCJ3iThYbTfx/PFbwCkXB6JAeQBvg5SxtMBPO
K79FGwbo+1q7Q6N7j6qPz3smvm4ZIusC9MpVsJGa4j1Du9YHcoYWzkc3yf9E7U2d
7ozTPVrX5ES/nc3g+efGWdeHLntRXusPpv1m6Q2a9pFJHD4iebYgxY45dwgD5J4b
vsnvK4rolmiWMdN3dEQTyBtXwA76NBu1gb066vgDNTc08qhzsWYmQPcY7/RedNXn
zUQJlss6ju0LbpjZZtGrL0BPFhpKsQDNsQyTfjFRdRu9NltC3NGBU+I99DO7zuEW
44q25pliRT3fogFgvIRJwdutgXdojFrGxOVjKLCKTTY7fc5qZMVsPtyfgSd5CY0Y
pl7B2M7SqgleHIXBbl+DR7XaJQbISqjY310CRGI4Kd4z0ouJmiK+rd7Q3d7hFHZd
GXzfFudw1suFOsCXg0DQPAD/jj3A3obmyYjo8cAn7vDVrnRAlWyKrPi1isIKQNyH
EmjHKvRUtDIcErdVsYtAE3MKKX2fDi3KvKWmyiWw0jMjn0HRI7IHAX0WKCytIhWf
uLIT+H996qQqJ7HxeqCoOneZ1PGUmhF+rA1yw/Yg4bd49xYCoClUmnRk+9yZErRs
QZ7+eH+nTjmX6b+RJ5PU2jn6XMr4Dcfes+XbXzsNgk+GrdfVo7RZ1aqRvvbvmT0R
L133rJU/es26NDklsvnLazWs2gb6vqswocneWiOF/nW2UikC7zir7PEdo8S2tBeL
wNUpkDJEXIJ4V7gb4k4gH9YlbPMiOLyOPPgEeXARRaylqFLsSpa8uWxDolATRBCG
1hSusFsSQUCDwe6QJdDOKMy5OLNzNbECRpBcQ4wVq4fKs96xNtzH6sfU1y+q7yTc
P28NXMg1wOYO3kqFh/uPXi4B99gwqJd+LCnsHuag8Q0vp1GHvzXLeJ4xJQnoXPYF
I2OIsEsnkBdQFN9Z5V3V398YaqhVEbxyMWk0+am7v5T1m7OkMoirqQ3PnIiDLORd
yM5ERzu7saQHZDcV5GeOMV9B4vsORw7uNfmNjbNNXUHp3GADBQlly93bfsBmHhg+
fKVV5IMZvOfm6fF+ByAdH5AWZq77AtaqUhEBNBtXLufOx7Gruq5rxrGB72m1kCou
nu8DtJUqEqfOMP1oR/jJyriMttLkcUOsRJ/ICIPLytIAmN7nLSHEf06+TmPdmZWQ
yDv/RHRQk7ITpKzTBqENFNeywVrdd1OBgByLMVFvYlqCPsghHJDNoNFEZAbOQISa
q+XtYfu0vXjQctNeRd2Hn53rAf3OyRbEQdLvVV3uXhxu76DpyHnuGipdqPMAh1I2
9YsWvpsiXdp384WSvO58Z+1Xx/z3JaDCdx1CL/l22VJG5jAX0frABvdKzizUBeqn
3w6dn0/tlXC6uFEUd8/gMIc8cQnbyMPTBB1puqMxXjF6GripKzzyDNC2WvJS3ec+
uu7SgHA80ofWj5p/t1Fjs8n+LOEionxkncLSPRX+3PTyC/79phScCRxdkatlcmZG
flZ1vqr1M/T6PzFK4sxpNJ7DgNbl1FYnjTQjZiEFQYXr1iNi/kUVi354GonsJeko
J6YfaHpvQOWdPbdf4jf1X5WPIJNue3rQw7UpN48aHsBMFWB90go+RVyCI2rIF9bq
bMeD/xN6QpNKkY1YcVcp4QihEaUoHDdbDJ512YPBaaUsAAk5AYUrOFcTlv3vMQEb
DCuCXYpxKgIavbXpl1GTa9diA1r+mzyVFKZobe8SVTauxFq/DUVFk86xq34ffOSN
81QOAA7GBSdh5T+P99NtIZpqOs4uAZdXvYXaMuhHVeSZD291xrxyfHOp48yfQE9A
Z2Ky66qE/dzxakQXFw6j6KbQHvreQNGcAkeVCQPJXqtMmyd+eL1iyr2+fgOEFbuP
UpUKCGUl4Aalpbudx2GTAQ/rcizLyQBS9wlh2beTdyjmlh7NS5cSo9bVnDHPKE6N
1IeHCQCEfG4fKbgoPP6OO3zpjLaDMQWUiTh/xrOGuDgiQrGHhNujf05R7sT0t7f5
EXLtXUZLwW1P7/84dPsOGTQ2ftAHu2JZuj7MuQSw7H6WMlUoSGcrd8psu5NzayxQ
Dx/NHAFI8EK/6PQlS5pUg1DkhxbAlGMS+UCTRe7XopxQVzEhN/xD/PVasC8ni8+4
scsmaMZORjSRQynz5zkj6s3MzuEwkJUdok7QZILlr4DYFzBjbjkmTQ5UKnQB2OaH
yysoqPPwjeOsg3hve6RmIqCI/9xMexBBSvB4Ev0Tui78X716pv4zYqifUAULwn8t
Ap1rN8+8McLpKeIsmkisREuN35vCssIeivkve5xg5t0q1tGuCGuVLsp0NFEBzyPD
pmXX4l7dg8ZpMp7JYkFQDudnI1WnEmQfOH82VlR6rLBQORGrBCyCzwAx0k3MH/+3
xUMl7q0H0pJCNY//1X1OM9VYJPHr1zo1SmtbGsWsake7IBzh/XTuCuDsHOLYyreY
gvEU6JzV4j7i/FW27R1x69Wp0w9eQmx1Oetur5kwJK8s2nWGKmZ1ziZEpYPSRePI
rod5gxyfxP5coNy3ZWfn6pK4b3MDSCilHrHCQ0mCFKIdf6z7f4nO47ykqbiRXxnl
BZdHlhrYbRVoBNBwAG/8+ETH9gfC2EM33J19sd1ikXhl9rz5fWFKsB6R1aGso7/G
M07WxfWE/ttemXoIMyq1tj8SJ7g0y737M9pCjNpIGEA8aQF58LVAQ/3zHjHLb+p2
w2PwLaO21oGMGgfX+9VN3GmROchATieM5LdNJyA44dY20NpOZ90KbaISTOc0//kf
VuBFtIRys3m//ay+Y2HtpfhNlVW2hEbZMJ77OYO+atMKkjjmumf8TIEsBq3NgOne
BSP5BSfsou2uy6ErdOhae8QLjfpVxk4r7wT+5Z10A4iISA4+UgIuz+razbiRjar5
r8iUCfVpiDYSw2LfLYjXb5VHtt+b7HhyznylJdDD0WhEOW3s2ZqfjDOakt4kUqKh
ZKGX56RhRYttU3NZyOYdP9egRJvk5XUEjflgcr9IpdKT2ORp8NsNdziyNHJ27jTW
9WzRYjB5dlFRLHLIiKpic4P5T5deELfw/XhTjyEv+NuWo4nkStF2xriTsxNVdzAU
5dy/XFz2lA+Ts7ngRZJtfdKGc7xhzS+tLn3Is5FI3MYAEgLePGQKf54kED1hqCUX
zc8e9S4QaKfjUQwMNIcjDHZxehALWUXrsEWwj654llKwtAN44CtQSB/VZOAfN7z7
N2pLH4F6q7Yos+qcMc5mIzdV3I8nxTmGXBuWZ8COTV5QsnU00G1nlpxL//e7Wszy
DNGM1qOzp5ld+XSdv/akFNjxRMlYHzledjU9nj/CMv1uHLX24aU2sNHHu1pXDgXq
qxQKUcFcCZusvesNEITaM5SNtg9dk2aBA/NOn4c36ys2bjviYC6+06vIe33pdlQ8
oEKx0CYW8dwmDrGWbNOL7gcNTzQgkgLln+gBVMgvMFCjLVI1OiPyR066FBjTKeaK
n8f1Yof4JM8U5XfpGjNBBPjdkyjRRMrWWHjJwJF7qoHevM2HFdrt+xvr5+ZyoZqi
h1vjgin9ZIxHUJgU83SGtALdZqo0kIgnoRxEVoIHM8k4/IaRAI9CNyQbjQl/xEgf
Z00vP66fO0/JmfvPoHpUYGmyjZnBniV7ToSk7JrrpY7QyW2HF519ZzPgrTXk6fe0
ryCgcLlDxEeFfp0pN7pZYf0RHO+a6qcOSLhra9sdCgIsl7LKE92WJGMBOXDl66Lx
tWPPPWLRaah/1HiEJBsUyjI9OpqiHE8ru6ZSxICSPzbapKozi0weN0KuEHjM7mdk
Pni68xPrXdcUv5iEx8XPYYDFM17BnX5L7Ovyo2eZXV2+pCw2jYoQs3EKQ8k9tV/U
4zLbpGfeKkQKmzvRJzPAT80dOskcZItbzMgCw8fD+wIs+tZO3VnFEsHht+L+Xv7m
VwpcCoU2hRIOdX35kQAd4Tjg0WrbtQkb1ur/LOHcip2Tle59kwEVWS1/zqEttHhD
qwAk9HS+Jpms8pAhIKqdS7Np3xQs9a1Z3rzNgXcutsaXRePyfu7tQMRBEu7i+BPX
uGMTYOjQux6h4fjeuwJavHkzobBXd0jBwuECj7zuoJTmrPebm/z8AtA4htPcXDtC
K0C55OpnfBQ+InmPWmGEa5Wj9I+szA10+Pwg1oNWBCfQDPv40m2p09BdhArCfKNE
Bj3DNcy8ScJmtbii6fCVSftzhk9YTK2MB7KyfG+Kg+cYjed02OdDYXGPYl+GfYHR
EbpGCYJzob36XqHcXjv139ekm0pm37vZZUDv4yuIbDnnjPIBz8aN2wQ74vYJCRiU
OtJWXl6twFXRBWx9Ji0JX3s44BnCtDBJgv7ogkimbLhSkZ/K5BBHuoxW9FrpScx/
HMLwksql7D7eXwwVpPJDca1KrhzL/Y7lOx/1QcBdu4KGGHmULDWjpDRNcjBGA3u5
DnJqLHPpjymb2e9UwroTWu9l0WasRjHXSJ8ez+lh8m1T80fVPdsfPc/zK91+suOG
DyeT+NfnOMeIpz2X1WsXj3mp+8TGzhfWbpV2kowTxV+erhEl91VC5jNDI8ZsBWvm
WF/ID/LyemED5PbHgIpN9Kr/O6fBsTx0Pt/12JKAXstQMm2teDrg4Gr+ZuYMo+0H
dulXCzc2viHDUeH9W3XQmOFv/jcImOUOhyKfmsSfokJPSqLlR1kL2pI+7G/wiq7U
Z89DWOYH7BZlouJr3BZXqcnJj75VzDIMAVLN+d/Lg6kgrrxIufYtrdop/Z6/cVhN
QCTaoD7LPNs6WfeXL4VWIAY43Tv2WFNYf7g4x8aRRpfF87MavaszTFdnPvRBb38R
9wtxt7gieJx71qH7Fvg5wKU3MFmkZOT1BFpmwWbaK+lMjpqHqyEVZUvfB2DhVEci
S4KJih/Zee6cgZm9g/64kuYu603om4GMbstHyo6xmcztKa+4ByI3IZg79Ak9cXMR
0aHvR+1yvU0j9jeJJbc+iAECvyAnXX0RMQU0DwvkfRqaZFDDSO8bYqzMhjhdOYda
Bsit1Q8YcGD+Aboy/Jjxms2vI/KTjlFX2wFd0DpN0V2fD6oCpzEskhdua2KHzJbJ
4jJCnztqOSssuy+uZsnmjCewJyWwMJZky39UKA7C/NeZeQZJcpJqKEUfZgcZJZxA
wbTwC1+V8lWDXSbXkizokptCWTDoPULHHh3KIcMxmplGK/0xEnlQ5/E7Pjhzyx7G
bSnF/9GWUueCvnXC0bB7h8eKHm+vCB7H86WgY0GolnrX4Jr32zx235zgiIzz4QQv
UI54Nhnu9wuKjdmkkQkr5gwWksYZNaoGA8OQ+h2kVxUEOzOtW145oZbg//W0M4ck
LC9w7X6QVURjhRgtrIEQdBYVjzwInbM2FcMe6/lo23hxnr1gj4JGYT3uVu2x+E1H
z6sqaWkpIDpLuEqBrUBeO9oKYFy0Q9tcAMnEvyCaTdeoc5IFbmzcQrTQdBdcyAxH
rn+kofYXT7xxf3v7lL+JyxMjC/iaYGAcWUO4SFzUthB7vnTlg3rf5P1JJ80rpf4l
mCdEqgO+4ugY8lCtoNSyOfoBkpRKNNMGtD1fjejxPze/q+NeheHFSdaeiXkuwM7y
lYDpZlwLcn6JzGDRee3KRA9QMZg7pcEkUH3N9iDvEMsXTw8WD2nIZhTI1P89/fwz
R5urjREgwGNobfgapicVmm0vExgkX6t3du+ByT5jhbECvPRAZx3gMyFomejdcdgC
RQHem7xOMjR1QO4VaJ8Hn81m0/vnDsTzAxmy4MO7Yj5in0oAVVXWeXXsoA1Mlp1R
+fCThi7V3o6HC/3aB47xWyBUkSC8qVeX5t00/5oq8Slm1vq8N5cu5f6C3jbnBPxx
1AN5YjCvWNtUIawU3ULboYKcQn/klUKsX7+lerveS8vB42dEmWZkCyHWwaPpghnW
6C0xZpNQ11LDUkY4Odhqr3pRYmjRdrdqDL+J0zfweWXbzpj2WJYbAk1ZcsI0dKOu
PsV+rk26qj6sg0+VH0yLXgBpmynIwD/hoA2YTHAHYa4MRn1sxjWWqcET7izluAEz
Zozvm05fl7yhPMm9a2WC8EZ7u1owciEMBGnU/iB2PiOBIZHdEASPXQIkTMU2PB8t
QQV/Ngy1o4QeuLt8omvcPCbQo5szUvuZ8BWksSaL5lkY/LNp92MlcOu5brSDlH3K
osrhZH2WNT/EubKqVf9ZNjHNk+WoAHWY3D9mMEkMwnrMgnA9ccF+KcCtPIc51RwS
NIY4AjLO/AxIyBJtWpO5uu88gobHJbmBHR6LkC0LlIfT8AgknMR5LAMYTLoKjHYR
c/FnMaYxvy/5qukOLNJtS8x2Se3ZHENbWR1LHp3pXgF1lSDbVIuARRSXb6N9O8q6
CzlKxs2HxjmAFLc37bjtJkIY81Zp4rt45i1ewQ5pfFhiRcPflpJ98Yhqq+28hEtP
U6ebjncWdStfzT7k++3FuMEYFYpVB3eqsKTRV8WW2uQEvb/hMlBrPxO941aHXZp9
PEgMnlDxafqpi+13GJnYi7Km/JN5PSzgUHadPGchbvOTnj2eJBIeakD10q+I1VfB
DisMZAGBmyY63dfVBfB9bcNdYrFnVA1MXmpf08EF3YNBb6gvqcM9EpULVOUrxgry
QhQdCxdVHFtCvMIHrkI1Awjx18EirnKic7jHcZW1JYv/BhuwP/sJwFNtW3+eGpLL
VYxnREti39MM2Tucj2OZ092ppokMst07nUJtI9fRHDxQEfX0yMOGs20rXaARwbMm
3780e2smr8ICVb/TNLoXQ4otuouG53WzqbH3Hn0XGg8TJzF8FkMQYiLRXCvl+ZXU
duMNpLIwz5GFCcxGNSGCHDZ3eOLf4zPcom2IA+Qr8/s8yYBt+T3GI26h8CP664tM
Ds7/BpQJ6u56MlyU/zDrQYFgT5VESQ0D2+RApCXI4mDf49QMLfgMI4g2KqvwNVAf
AwV1iR3XvsdmKBhlVuHRKMaCJnOE4spmVZ+xXmyLPjkUciZKD1AWUM6dZXtFXA/A
bev+BSzMUM3bxj4xaRtyHzi8BWCKQvuHwUVqUESsFmlt3UXRiw6MulykHJfIK/mw
xP5JteV/3OxssY/4AXV5dMOp+FbbVN1U6tWZV3iIigaW5u6kOjZjwhOClXJxamUa
RQj6bxN94Jhl+xt9EnNYUoKH1vc4BvzRsVsisU0mr1Oth7TyS2rDnGGCVT7Mkvr6
DqCbtOVLtqbEQejAvxuib3lEwhV1p46zRPWOqMgLzeDuLI26x/cq7kJYlvPVul+E
5e3E4YfpOAW/EBRAaOdJTqUZkz7Jg0793Xg7D78fjBu1cYNh5pbK4Ma7GgA+oYH0
V4YLGF8FqxQIyxnhywu6xC/NQ92CdIJ6APyGYdEYR0uxVpKsggfo9Ladk4E+ET1N
czPuFQuL7YDfFPIcMDKk8kG+26KLkngtoz0bN/kIe0J2XeVMT7feh1m3sgkUK5GA
NpaoQHfAcWat300OrkwDHnrRACFUGG/5febCugYgvV+CK5GlLV1VXYTYfOyZQXWH
3zgYbodlYyH551rwG0Y5sNgakRD6aAcj/aRQnXex/CFB5nd7hZ28ZNslVhG2T5GK
F8hd/xrxI1MTrxHr41SosIwEHJTSbEfvA7i2jtjtNOgJzN5wmXCz1tvONYFTJsBg
LdIYKDTiPCPTd8oNrRRkMVO94wWVO5IoRmwfYrZA37axXYNLXHkdCfoPsMA4xWpe
IkwUVAqFdFexram1W9Jmty5zNpvYScY5f0+arNhDEoFx1Y0RjPKupOZr2gL0STL1
U97jGDSv1YIO6F+ebsEbMOB+f6Oqv9IDKQQ5BN/melqEtkOrU8/SzHLnl8LIczYY
QSdRHfhistOQEasvoQYobne+3jy/wLgJ7BJRgbYFx2s4NPV6BvV3zboOysXMLzqd
MaRn1G8VFNqb6xV+U+Q/JvgVI1Ul95CLD++KdCPutOBkzyIRNT/Di5kj5r/dU0OD
noANI/GHfn9zosDRapFE+kq+sOvXM/Ej8pKQGa6P0JCHhD3vazv0mqZqoJttBIYo
oEXGRHV/fTjm0LZ4abnq24/RH8KuzSQ6tgwhFIFQJ3j2sNEwYPjfN/bHh4lNkHlk
cmmg0kcI1LyLirnJF7XKgb0KvcQoa6j7CKBk+f97a2u5XL3smK0vIqvYsJbZd5mY
FpOAc2Oidx0OTTiHwo95zK/jS8u+DMzrWGtxlfEKS44adp65f7B5tEMUH9n+lY0H
v26NfH/jrjv6QaaewzB8wqQlNmepcx4OQ1lYeyFeBAfHa+qytQXQL2trnuAbFJKF
0L9Oo6iOrpwZ5ogDOthFM2W2NAc1o5oNbwX3b+yK5y2eXJw6khFtzvROz6r/qZ4v
IhUkeF+FU9KOUrQkOJEaOXKGhoWHokokOAaFZ2bgWJWWAt2gL0YgPL1lwLo/pkiv
dIpU1oCIQVMTivAlXhkDdSfW1hAweBZEc/oLPsQZF1Sb1avABKdZsNbstXenjfsV
Hr8Nb/pGAXMMg0YzTXiBarNgiAohRJNc0wq3/40dMeoUnSew2X0FLv8G8YpS3yh/
I/mpr/XonTj/WO/cMPKZ5JrqlPo7/23OWnhmhVoYQxzaecSrj5As8C7ZHjf3OymB
WNRFkRiuxFQHlQqF9b4zNre3/E8KSREJM9V4wetDyxT36R9P+miPnK2MfT64WJvK
M1GaK6QYDWq7ND0LhGMPzrGVmfwZduRZ9yqradbNmCvVybVKKvxPFpaAHaMw2e0s
I8mo9N1MPEHyyNP4KtC5ybL4FNjEpxI5DKLfmW6oWEwchk9WdrCynZtDEygywpD8
+E4m70xdWwXhSkxu7PXighlKqP+/Fther4oCUCZOP6S/y2zQRZ7sMU+H8fc79nak
Iq3NspI1grWxtOoSWgbZT8VkVKWcVElcpIusUiZ8I5ZMJDvCuZR1CpkLWs6lKs4f
QRIxkvnCboz2CxGdEKEt988XKD3t3pfxidSnIBLtqZTotFSQD6dZmFz1uV0R54S2
FdfmHqYarWzoyq5QOlWaMq41+mG9EC4Osy1rX82TjN3DvkRENW6dHRWHbgHsLy/W
RH57H8wDuUgjsMKtQj/AO0F+XVF1SO3+Fw0YIISytj6EoZeSAGufpObfgy/DPywD
lVJ9ag5VNXRMl6a/fSok1Zc3F6YkAof7JHJORK0zaNj+GFbE8CqdwjUCc8C8rlbT
rP2YnygFUb5k/XpV9DGY9zrldMXh+GYSyKDNXCICdicz3MdRkYo2Ox6US+FSdYex
Elo1DJErLZ6S940dMzdRJQPYc5KWhWk2H0RY8+qld7RcJe5VIG7DhZ4M6d6E8utV
deUr5HuYHtoH+l9dMPuFWsEgkodXe68ZqHm431vhsXfGQMEPKGZcNpAF3j6/5ZsC
a+QHRoxqKwjZyd4Xr4n9hm3sZu6B12YdRZnJFIJ9CSV3+R5d1+WZbQB1AcQQqYmh
ZK3HeiDfmOPzxuoq4GUn+1TukBDstkvyVS5YS14coGSpgo0rszd1VORPdN8Qhz2x
cXRa+PcXWvP+eM75/rmMPH7PffFu9/7f9O1Hn+jHUsvEDneZn2sINkbE8ZYMmXMf
8f2q9PCrHc9iyU3I0k5/BToSdZnJ4siilAujJpNcMBBDn6Mkj/pc6cA2sXIs0KtD
rgVqOu/570wJ3CzNCjOA/Ve5A3dYs7n253MeMhCbINWsv5LYBdBtOBggOUTrCXlP
L46CYChMlUmiMdC0qgQE+d9CssGJqz8CD/0UiGFJfQcEDr+1d4V2Gk/f1Qxt4eoY
V7WT1przvAsgO2pTZpin8K69EjYkXMLqZU22zbz1bFhy716R5sYea6mNvH84Ajk6
dvacUUV5LOcKJCQYlsBVNrzy7o+o5E/1iaq4x+EbQ3jdhXxUEHhInqh3SKPd/940
BcC1aI7UkhPqaSiNUrpERmjZkd/7CCw9aFB5UrDxvIVM0reNyyvodZQuy9NaIuxu
NCAHoW4+jo/tjvdlYMNKEW+QBJpt69mNRiBiURzYxaVYaPOjhs7IY40WyIcEbsja
inVYNGnEco3rzuzL4e4VDrasbGz4KAop2RAZ4fzknQGCB1qCTZn8Qqi0+Xvo4NeX
k1Xn0QBeCS/RP1yOdohX+QDnHexQ/snVlArF6IFTJzqmhv+G3tdI1pz6O8Uk/a/F
nrAdn1nBbFPq6Wrv8lm+9VP6HiWxrkVryxMVBoFoGCAiixvDoSumgE+ZeryZy0rs
nI+jFmZ6t5VWH5lXHIv7tu6gmWN4qaEXpbAQ28AidriEmIbWoQwrSU6jsM7AFTnv
WHifYTAkbQqSh8mmRycb7IeT5+Mg1BkOCq5AsJ8uwVq5Az68AoMU+zl88jVO58mR
SNlBWzVscT6MqrtEtCFmJTiXdLnEAM0iO7lkqKKO4SRq4fQOKhxkQDcmw7i+HzK4
tYBPLd2CLn4J58t+VXmMhnFXleippFeRS/2PbGcaQYv1K5Lr/5bNGDD4Dzlshhlp
GeZS0l0bfgBbEjSlQM6laGYbKtYQ36wh6BV0LdtWqs4YXOnWmVgqkgJjXU2U6yFC
TYUJm+OgBUNi3g+Gyxrz61jhBiwIanEqAiPUTNmMgTdpP+nsKTvM+nAU35N13Vy7
gcj5zhzFpXvx0WvGdKgRC8z4ZXRPTrdzfc+ZSoyk3tB7aVXAbpHPccwMrUIOweD0
iP/WW/fC0x4ZL8l4E+5EO4XfUMDngyrfkSDAdbx00DF1je1gblFF6JcvcuhoWMFw
qNaPEe/uic2Am3Y8tF7FQdyHp6yHfjEvq8MB7gliq2ZjlRQFWCbHJ3aH10Pkj/C3
7Q8OrK2PV9eJVrRTYXG3Sz4CQuahr54WS6P3nr4N6RMEbZo5EKq76HfHSO+vUgD+
Owlk9PTfTUhlNveSoJBgo8Owr+V4rb8ssfPGsYkTasALN4seBJweKVoOKUuNrwIA
/kwt80wNIx+WFpNtyTqntABcu6Qg/fsV6h76BpXkbgHhcW6dkH/c3/DGZHnPYqem
HfHqRfoWBkjBQ9ITrPJQH91eSdn+Tt8PtgYHPUuj/4Xg/dy86Uxbe8Mpu4I0pMeC
0UNqwSCRPVMoGj7hKqqe6LvqoG/sHJEYoUYaTd8pZfgALw9iS0EltOfnT/jBXdny
zk627lC2dpHSr5wkDnJjR/jgUjMyq/oytCRKHoP3WGVL55Bke6NVxbcb8CGL4Jhs
GBq9b5DyRZIDlQKAsXd1tPDSTle7O+Tvj+x5lw3fGVydvYgcgjAxvIRerDtNIj+O
wxGMmB9BjWjVA67znUu/olx9/UzFWN/o7BNUdhzC6YfKpOET8vHk4/E0nRdAcKYd
UXLdGfAKFGI69a2j0Ug9Ei1SO88S+Pr2ToBLHGTDNyZlzStzKPc2rvciJWOOxjpA
l7td1IPGZSocjOF3H6eXNNfElA4hojuCRa8Rq1ulusFeiIPWa8TRozQtdifn4KoO
4KkdgEDjHf2VsizBVw+aX4iaeb0EVSgwubA5F7TjvqbTGSLgyjGYfgpJM2Yig7yH
OBr0oi459IJlVri1CwNEwk9d9TCknN8MG5p5HwRpspgWJxBmC3cD6dGrmcmN2nO+
h4DaUIdAw8z24O+eHW7r5QegVLgFnaswDd+hZbQDoW10kIYhvf0cbE5OWbKKw7MM
GdHczBIiXI3tDarFSZ4XrWBCDbrMXjqDxnfNEkRsZApbDBYCPjW9PjddSy/rvhe4
4TvobWSpcSFxCdO+HuiS+PG15Piir7NFDejp8yxbBdi00wLxRimpLqresAo2ydSp
xb776sAmKy0KTYHTC05R6Gih4e7zn8mMB5L/PK93MX1NG0JwsXmhECfvTN5Pz9lp
sx8evEJai+hOuW+VvVT8nlpxEUdkrto9deSf4ZF5D4LYlipivxl6sNZcuU5X8h9t
ZsbzSD5D0kDBs6+MHetCzi8FKsWVUk51t2fBB039rJGw7I+n+QV3ijMjn0zxHyVq
wY0yVF/UiFbP4RjuYZ5NsTXc5Zwuro2PtDWDfegbNX323ED3F1o1+gx4w1IbZQds
hQyvSN6JpPIn0YYivCGx6yeTmjOQKN6ZVhWCFXVBS88D6ZgyZ4Ar89YkCnAvuOkR
BVBgq1Ym3jTRDUlgM8CY63lWXcYunjpaxkZ4W/di10ELesBc8D3eCuQO+wPF2BUo
0x/u3xIqXKdQnZXzYasyEaKCdQllJsH7RfD0Ty2EfKkkvLaBaVxTHTh45Oc2SDVI
jm3Qtzwq+nB6Hodu5JrbGK+ySpjgNe8jfwXv2tD5ua3YnMisFnDNDhQHt4owjZAo
XvkSJIjSA5DMxGzYwP9/M9lENXdRGWJ7JjnCNPp2nO2cYc3BLuCjotZjsjMRsQXv
L2zX8G6ldnW8w/vZVpy1E2mjisz29rTkMsy5GUbf4Rwyj/tzEQbuSKAhlUbcfFq0
8YW52xR1Mdho9jImnqwak5MUZbg/nwX+HRH9vDKRouQHfHqJbx4Ug9OnNqLSefr4
GIjjcEFNEVJwiF2JtSkIsx4RPQbeE0n9LbtqpQs7xdTsWsjxFLAbIaZkalrmTRPW
be9+W9x5ew3L6SfUsmjQHZaRv2HOXltevHoxTqhAbZVuvWPndx014rYy/CbVNynZ
r9E92SUs09p13/qbAGjnxg0oVSxudX4TREuuBBaFIEp7frM6L1I4kyRhEMi3/64a
IlVyqWcQ9/+dxhgZZqU2TfoVTj7qg5a2UzfArxCXpUv+G6eoRjosz4JViv2dWEDl
pkFaH0WeTCGIJ4JLiJ5fPpnR2PWyd6l1Lp3MnX3XpEc8iLEjggo+r/91xWgutyNb
aWVFJJARakgzP/h0QG2ypm+hBpDggaKt9kYF9brkvoLPB3x3uL3MYHfjiMjw1BWZ
LR7seuMuota+7pJgu6utpGhCAHg3rF+W9zSFo/nK4gcrEquKKPIqyg+MV6ZANFdz
JXtS13CTKWGpJliuTnR8HTxQQs7GHliAQ1H2FUwIVKIRRSDRjK4OLcu+K8UgGGed
pnarqgp/ksmrcvf7YiOcWMJ06T4EUd8m3tMBHXRIAUkyI25Fx+0uY0wcZewekWC8
iMqMwWZvkehQiJa2fA/3Xbq12hQh6Ok7p0UxeK6ejtgovVPVVPw4W63ORXxN8w2f
YSFWRIwRNfOdkrIntbGctcwHxQGYBsncaVXirlKA5yPDDJS5R6rUxozk6NXBB7j9
SUm2OPUvGYzrvZUPNLxl/WicpZL5ogrXdF8mu3gwg2hG27OOXGVpFlvn8R8HLQiG
9mpzjgIyu7sxGwrGhHAsHM8W892UOmJYi8DcLZQ8zVIByM3aBne6SaSDGFp5QVsb
8wIllyBH2ZG6UrdOaFZ//0dPQZHT4bGBRdyfVWOXW1R1MCskTWNIbYWsFNMN7lA+
gmHQbYUkQEA2N3bnEbIAMdk3vn00o16EofdXD4EIcBoU/GL/emLq3QB7BB4WvUXt
EdsOlSQWWj8RlJW7dJ4tOX74YKn5UURzDiH3YKL5D6/b9pQE7IggKcbC1aQR7XdL
+SmbQZ6PJsjyellNsLLvkvMpbmA22EgL7pX+RnDet+SYZGdafIrVCrv2N3ZEd+v2
BYN/VXwrZzVarAYoDTlHoqMnHWJGIwlA9gqInOfzi9GITGevYgBXQ2zvRU6dXTKX
EXYfLEE+cwAHNc5BbPj/ViGv/VwE5u6Nga/KfpveKA+YR9p3QQFkRFjFAPSmZ+s0
hsW7eCgyxy5CPsKAPNOFvBT+YKAPD1rS4zuSADgA0SLvh3fEFKiqwnmVQwF6r9Ca
7J9yHi1ZSs01L2sp2Mvbhmh24EvSBcy7vAMMz2lnOC5L5mI0bpBMMaTGnAvv+9bd
KlI6zzQC26rSDzNHf00Lw52w67eUbTKmnmd9t7sZyE+aXT+QF/oEbByLeV9e4p9e
KgW/mS9P3og+x+dG9YGQ+lnZ9ZGXNBIPBGcmHbt/4RHdFdt98f1OKFBgzqsg5UFL
klLTZEGZg91P6LR/TIF9ngGwAfFQX2hxOLaqDzRhGGQZmnI9MX43YBOXFlS+04gS
WOvvkHJTzGg4uWTgFFL3PRJyOC1L/mkxDGGwDu1Rprr7pQEaYharBG9+TAGZwMv2
JjD0FVxHNEFuCh9fJW3aIaaGWqWOHJ0OgoIlsL1Kg/B1RbXRb8oujwTb09D9XIgV
c8QyNck4li8BtQpHrLrgBl71GskIMstdI2OO05+jHjiv9QFlYxHE8XqDa/dMybqA
873GccFkUYjVkBGnZF6+63cIR3rLWDcLvuBc1c3WrGWbyYm01CpmYRYVXWm1M7rC
YONtUql1f069wli0dyZ2ijQC67QM4hrOhxEzFE+PFWAGhSMn89wWUJGr2NIJeJ0R
fJNXEw2ZnnaamQOhAtM2r3KhBDznvAbIeS2HJsV6Xj15ivBUKuWqiC7WGpYYkRck
28oQg4D1Yr+7uXrGEYB9r6aDLFxy7j/jCX+Crmw8bzEQNRCBYt2mOIEiZzcWEdLo
yYOYUiO6x5uAyPCkbSFhEaQkfTWM+aFdsJ0K0y7pLg+UDEqX5erXPvz4HsLm4aMX
MEV8sKrD2eS6dR7hxPcb32F8knFVNs6yRNsfDQS2zuJCsDKq7HqfrtzEY1nZwd5M
uM7lVGqnxo8uELRE/uGKNXgubtjEc4ISWiGMGjme02wT88qZCFXwTdoYvRMabY9l
UMZeJckxh0IXMs7IEniTtNitLsRG6rFB8CTmpRUFYGC9DTUabJPJRfxZnPW/srQe
Aox5Sgdhy0X451Q+VVe2MkOIpfZipED131dRqED6VDgsYYNquGm27SiMm8ckTC8t
1HjURu6P6IRlI8BYi9rNze4+99i6xm5vv5OBQ/m0xqFOffEum8vSlMbp7XWbkAX9
zDtybDWaZhc2lHZ09lGXe+X0mOSfhALVi6xMCmr/LG8N+23VSfP1wXIFbU3UpCpi
PUmgmgwQg9wAKw7Y2+6ezU5lDUow+FfJhPfYRMGaumkZoFV6SvbywHUIDX/tkq3i
b5Y8s+xIiLc7pkaaEhwgoZ1oa9QRHWkgA/kBosjgAFTP61/yf98ST+qoeJTv1ouH
dwVj5rkV+PdLRV2lJJ6+5+Ky4x/yCioFRC9+9EzGX7Pncxel9Uytxym1PNUBQW1M
9+eMlpsjhq5DfoTrPLwHokkSoMhLQRol1DH8yk0BjYZ9W9b0bw5sSiJwBG1zN0Z2
BHJUHH3NMYbzaZShP5DLWchro8gJbrHQJDlKJBO37uyGwKaYSh+L4ibfW1hWxxxR
33n+21cI2dcyXYJEljyMJrTTB8E6DZV0dkRjZ2q0GoGBspziE+TgXzpzkkWpRy6h
ooYRZiA6CQk7OouX+j6nauhjlCTLnHN4g7O2XmZ38EelLRjL1ffeF2yyhSEfhhOV
l8FkwSSZZiAgCb3Bd0vLPRjaZkYAtOinsoUrYYowc50VElyBEydgRtwAgaKx0Mu9
ueOEnUt2ti5XMRX4kgLRTHmYx62VzIBWCvGUFME/MKAeQAEtXZCkGyAz0rf21auC
xEs5zbWmk5H3mTSuuCDvK+mJZBvaAmHaMW61yI+MWwI7+mSOB2qcFgaqx6NRX9Wy
EtD+iq71dYHh/TZISDTh6BMxu5QIh+R1ssP2iT9HazV6wxGfm6uuLOC+djk5mTsr
iu0o1JXXGQ/lUYP91Kw35W6CfCN4DXxweqRv+WfKW3BnOUtVM9iIsMMEzZ/9hLoa
o5FNP/m16ZQ1dzllNMDslUWo9r93oTrYMRSLs1LyiX/kfyIsB3GDfzuqUouyNvaQ
J3105rm1fDUyEnjZHUN4/54RaXFQpjbYP1EFMNbsJz0/5B0bDyDHmO+zkK+QX4iK
sUSZq/Azfg8xm1nJI45Bb+C2ycBsGmaiMZOWCK0rN2nsdmjC7VqNeX332rJ4kJCP
uY1lWNNO+1HzzIEMYrGD9bpI47ECphk+drJRnPJ8Q2RrTZHN+hIUZ0lXJtMyBtjH
hUTp1+6xi4IQZTKfu7AwLqw7ULGzpVqvNXhAQVhNzebnK+t27ik/xb5+ZTwv4mq5
YySFbugdaK9MbV39k/DUd3rHlIHBSHJJ7r2JUqz3yAbSfcMFmTpKUhhaMUdyrNff
HiJUmLkFsfmI/pmOQz9w2msnZvjAm2HRizVeHvijSSaDrJ9vfcjPTPMXZvX+imTg
FZfSwKkih6WQS5toqxmKlh4TrfbzHD5Ter4sxOX5FjhFNZLa5PiozDjSZM9WFi0d
1Di8tJI/6kCp57AzRlrGPwK0fFd8Lvbqwep6rIzHYOYp/xWqr9L7essmX3CUgjvc
dBeF7FO52zM6J1exRFwP8sAYsi4mLIHDBJ3ZYv6i8e3WQF5YndRaOlXYUNWf+wXk
/9waBqE+gKaFbdfVf/2/OfO43xPEj65FAXCcFGJBGUIpbYZ6EA2Y7+q+6HgTItmT
aYE+bhJmC6lYFGAhRWRj496vQK2dNU3Z0NM6IWsAoZrQDRdKCUhbiwfi/iSgF5tX
ITLynC3HBi6RfaZx++VIBM4vJ8d2g8ZqqMl3+d0treWLxHo8f/c8C0BveseeUr/e
IlWrYfLeYuKyOKCKTdot18kFwr7iY2SFoAprLqL76+LLMBx9thgx75cCtv/pRdPU
Ez2SBtA3kanLvRh58Mmj40CDovym4/yQ42O5CynxZ+1s4BU9FDHn3x8Uoxq/UyRe
RUMCxNPZZ3bFPuTmQTaxp/yUXg3DSIeXOBzH2MMJOOr1AYasH1lUk6L8PDABtgrr
dwz6QW+5+bWohbkMUqMMx9ZHs49jkjN6VLjjO8GDqaiDymSuariKaxGBCjlIVMwo
nTofKJZCc2utgKr76HzvbrbiPtqZ4WoRmsmYSw2tVwpUqd+V3TqI/iJisxT9bwcJ
UNsUb9RcUOlsw8AQM9sEflLBGf8mTaI0RDHxaLznMfN29Bf4K3BIzmrx8rl0J6/H
lYefKjMOEfGkPUEK7xLzTJAIznD0Ibtytq/XTlyF8+nqFmYN+99RnvS4lKtrR0Sk
Y9rZbtJjFvINMm52e8tljOJRjrApnfeRXGCZoFdzAIGvuIm7Z66S72s6O+15oqv6
s+IyDMzKeRTX31I/d1zHGTb4Z5U9QC504fEewiG+VRZFWj4b4IVpDgzW+fa/Yn5M
emONqcdL4GfQ+NOe90vBO8URnnAIYXYo9Zq/OtmGDuv7+h5QUltu8y3Xs6JmVALh
GIEVMtWUilbLaFEH1XND7A43P/ZSMcxPZRc3FfYCkOB2To5NFPrQXI2QoHjUE2Cm
6ClKZFnL2/epcZfo/WV56qoFxwZ7g+krVLx6iwzr4t1h42y6e4D2jeLGoKwcuY8g
Z2//hic4acg4kmPesTNFdIqQgZKL9UzZy96FeEjh46c7TYFRnBWMXLh5+jqBcmRj
X56EO/Djh/TSlEwj911OyhN9HhwRxBz2/ea/JpDUX5B8cWsA5/nVQQ4H8zUYuFsY
O2qh6H8HPWJ/xUid/DemNNsBoTIillJfId06zcibDG+OOi3EYmSZBgJ+0gBIBcqI
wqxNTWjsv9oG3+pb4nvaIxcnMVZty3gXmY4bySN83hNWgqYmjNtiXFEWbZEgIfAc
CMj0yr9oUFJNFPhlNqfbNm9Na2N40PaNySU8FzzfwjkvEBeKzrs2owdY413X+RNO
cuhkLeYaqDZQY8OX0dWisj0+fvyMx6S4BeMXyiOJ5VFcRJU9BysS5P2ErLXHr+Hs
fb/Am3cF0dS3IkPvuJfG5nNpvK48MCwf0VLU+6OYrB3tc7FWLGeNkIVpZ6DIk0YA
KlUoQXQgyKzu/5jSAaGGwEza2P+a9t5nW52xTkItyahFjEJj8k02Y7Z9K9vfxeCw
H8o7N27mCU9577cnZSf5F5jAv8ht88NLyYtttT/FAgQnxkooEURVTRDHB8F6jveu
ejpx9SZ3kjmMKjPvgNGctOF393nqY94HpMz5p6Z16o2WemKsBwX4k7kMZ1zqCCXS
Hwge34VvhY+tHST04xDLDFbW135XIuQzNXK7cEYT3WsKNyfE23DyROxEKds0CNwY
SqbLKPA1L9uZeJ79lTy5kZBCVVeUwEmKsRPVFrciG/vpcM6/jVVTxx2bsC9mErqJ
ANQurwkNOcJmbgEceUu8RV76a4vsuURPuX6iYlDCiy2cFyQuEAGXVL10ZuombPKt
9/eTWxyDwT7o47lJah04Ct8/jZHlTIsfFISGBMq3vd4U/YISR5otlGbWVvzq7YEY
Wil5+BnqU2cLUCgkbYq2sebOkGvO+n22aXV/XfJiFbgLD1WoDMFpANAK9sx4Eftu
m4o7mI0DROb/leFupHfNK8mEqT7JRglN1JL1s7lQx36xK5mdKvwO3Oi4I+s1OdZA
s93RBU+CdpRfN9aDxB+txVT1JRAgldACVjumSUGBVNFusRUopjhoTUeMp8nKhodh
5OoovCK9RX6dzcAx3zGDVVoj+9ib/sHqgPPAmc97H8tsIR5cMRSRN24M+yy1t7pa
HLwIBGo3IXptk2+xKl5I4PYKgpCFNiHmcBn36g8rLjJddQkSpZUL+NdoD+OkOvh1
i2Hw/KKv2lExqI6DgMoZh3F3nnUNVWakHlHjcytCOT2+QkiHS4vRLYc5bQ6lWKCW
y6qWzoWqfxhSOUQggn9OIAiPHeeTT9ePflYXAigD3k8kKi0hosKblY58O5UM/J9B
zh9UkSXVk1KBk06AiHsTmUOrmYox9xJfo2ynSI+plaJ7qt09cKTvo/6RU2ylW0HK
EC2hrBxwOhIJFYhaMhUs4wycBoIykGOzUnBcLEatKOHz51Gqk2BrVNWhE7MvAep0
1NhxcDy+GOP8jHbQyICqQpeRDer5hlxDIcEY02gSriME8oIjfHf6qiFFACzdX/JL
G7+t9wmc6pL2T4H2grdMHlp1U//Fn/97lneeec1cUqvlnWuyXHFnNQM56bK+BzPY
KgHn/KmKmep+zwA1mkyr71xXkYvndEyQluNSk27/iv3wr7u4tmeYwhUWq96ymnYJ
oxwJHo9ggSUQ3UjD1RtaHhu7TJsYUsQWipEivZSUa9x1E5QgVxYKqy7Ijon4gEnd
sonOPK3r6BH9OOPNdTa2ENx9yvcCvard0t94LyGRi/wE+DWDFFDgZ3yuUmkMCIzv
Bml2P1hWAEA1MyQ8F8XrYE0CFxktY00LX4RtbY3/ATKMEgCSwyjSPp3Glo6fCrGj
LTAQefwu8fvnjp3AycSRKCkw6462FoYtRKGzT0i6R/daoGjoex8zVYV63SpOpA4C
FX6outTpvUUiNw4TNEcmTo9ALKsAk30Q+hhZ4KCzBtrnIklQKzN7m5qzYYwDKs7/
IUAQTKxBNawWA5PUn7ykSb9eNRbbR+vcgmtjcDQFrNartCqoJCkk8VjdhaWnxLWo
jLi9sWlSUq5cFkP5JJinv0gelAd33TIhvPydmUoY9XtrFiUzu/TkywNFvkD+SOaP
mmyi14UWYkIEGjcx0bokKrFCb69zp5h/Miexo7i5WmAb6B7qxoiWg9B0/JYD9/3k
znQJxCkxoqj61vy/I6hnSJ9AChWuEigMTCNx9efNvH9UeMmD0QS6ANkCRjbu7JQp
X8ifWE5j0ZT1ycsWOhKK6uJ/xxSA2Uq3CLkTyVV74H0VVMdFAs6/ACLto/ymbQTP
C3JrJZxcXRlDDXFQ+eLywEH5VlAoJG1KFTMnc0Eed1GBAtFkyL3hGFEMQKLQpQr4
xGDj7ORhLwn7/kgMBmPgbXH+BP0q9vjDOS5QbVDfGzlVQvzq172gnSNz3GUivQSM
4azlXKmV+V+/2FfnDC339gXchYt0GZr+mL16wj5sxRgAk8Y+kSOe8dZcqwTTQyJ4
ArqtWxyNzDta9nQe+4SCVCtoGpi+qrcR9JHLTzhxAkVxkMnnkusRKJLKHWGY+gNB
QLbfRRwCQIzOp0TwliUqPSAu2nyvb3L1UzmUa+Af6p1phRobX+F00m0oCyv+UXSB
doiJ7IusVo5kBihduFkyeyvm6MrMVhqqEKLTwCFGO1LEghKhRAZyDLm2Cek5XdBQ
jRtirrLLTz+DOHwyp9u6G8d68gbS3DxViR1n2MFiiRTvOq8hbgBt/YKEJB7TIfrQ
OIvAYdyc7GXmfUMFC4930PNPyEXiAw5ITGny1lYvJRHp2SvoGmqck5K+h1h+y/Ix
8lqiQB/25Y3j3XYIoh1/tvPh6oSg79isFhudFmqYFRiSRhpcV37el9HdPSjbgoPM
0fjgbQZasMD2aW8l3f1ylgeARqCESkVJmdxMRtACxt+Ty/w3oIQVaFE/YcgW+RXP
0p1aFbPvAU7QGPVh9h5DEHaxVAC4P1YOi1Hg9Uwq3vp7iZcEDhinidvAIddWsjRa
5iiw20F/0na/zE9kQOIqgXXoGG8AVq09UktOm7eY1CKzy1009s6qH3P836MEqW6t
4/lpSirO11LuvX76Ytq1oV7F+BaINJLMtclilMm6mB5Qeab3vLgWZ+JI0DriOFKN
1ScY/XPN2YssUzDnhIX+/HHUiGKknLw2JnNQB4atUJyWOcwGhCgX31TWnfesOY1e
15M5RoegGdC0mHSskdnuzIRf0r+B3mHBFL5C3jbxHIdGXOmaLiqq9VuCDJwMyg7+
9bGUwbWvylFL+awLqVfnvsXDkoUhG/Wr0UqVacBpqCtNTibAA2Aj1mA+fSG1HQqm
K7kClIVB9C/TLv6AOUInbJ7HqUpD9v464STBvbivHXVYDZ7JtLPGZWTe8rMmQkP6
Lksjmkh6QV4w5vsJDv4S5piBLJq2SyBMYIo7dNe0zerVwdq2suOoQCdO35jGLLlk
BNPVN3PqX/ydjWm2VEsS7R+ItjnKIWbGU8oTW7H2J8l8XiQJNVZ0Iyy5l6Gf65of
H9jdCPNw3E1H1LUwPzco9l5bVDuxvIPteMLhi2nWuH32S2pJFFL6pNR/uFcGSz6F
OyOFRLFS4YThszvvGo/H3XfgzobKHd4ghUgk2iPGcqKorVVUdq7PpOpY7+Yp9hQM
sB5KlZiAowFKMEcgubQ5WJFTwm674le2cyVl1oAeRIiQg0G66HYxBZ/L2VuK4+rN
0D2+BUKuPt1aZMj9xM4iU1vfsW3SnXt1iTx7wWwx2ZtRYnZXAGMSrMSl6BYGy8cJ
FGhaT8k6m2HJWeWXpdVFK166K63plfNINlI4lODIjqJxIodsymcwpouI3mZJpt9t
ORl9axvjLRz43ILCHd8Zp+9UKOcFA5xaSatbaXBl2cvMVmE706b70i4bCeqnqZ+s
5QpmjC7wEdF9Y+ukuv95G8FzN9ezdvTtwNpJYQMmz94kUnuPoVzElCkl5HtDlY7D
7ULqDr6pvDbF6A3CvG06bqgW7fbtKZ4f2dFrrVVHVsYK2LlcTx1MiDfsOlnll0qa
i4u2bbYi8fxnXmQuLOb0myTbt0lASMVwpIUT58ct2gXB39AXH0f5rZsKsnN4KbAA
grrzWMv95VAb6yErx1fPKYld8R9hcnat2BinUimFN+zKuTWNUqEVVtty8RbYpwpr
nM3Z0j5jO/09VFDh9h6oRDg4ga65CbOcIZ3uh0HnZuEQSb8sBrho/jkB9uRUoBk5
dLMXAmlz5xZ+oTFkqDAwxgE3lM1D0KNMIljEgyOTw38vF1IlwBbF5yu57H67n57T
hOYGgKuIREsrpIOHskWDSXmcoV/eRol9PmN4/YxVifYJRnXhtowjHfTuIqJm2218
99DMC3Ol6LFVV/m4K8CMftYDZX4nwPk2FNwnp7omfkqYIsCrKlHQ9blS6v9tdpFN
PooHfYUTc0800n8cB/QBlDbiYU0IQ/TFEJBmyktA0DeQ1yTJnW4xfHPF54w2VotZ
AlQXdtmlEgYNaLDrG0Cgsi0U/qdmGfBknouVtohl2maB96ejSC4tZMc/st4m/lE1
298akXgR9lFEdlb6MFaG9Mt6N2ZJoZEfPgboU/xee8IsxWZVguwNJAuSjfOMJnJ+
guKukTeqSnr/o+izBPhhVHsszOeEQsMsIxu0/19VgcGJGNHA3qE9xHTFKAtmiTAC
9Ti0PGxgLKnpizfEhv8QFF1+kjSK00YsMue2lRYrpJoxXNG37CGmI4mo6VNg2lr2
FBaOwMhI6+wXJU85fH0srTa+wPm1UCgWzU2oR6q9dfGVbNeZoNFta11Z3P1kJCDA
AKu/4BSCK7zLAYDZTGEhDTKev57U5OnCZzR1ceulIgtI92Ba2uDNOaO1UE3LUtEo
Ir3IWb+ktdKOa9vmv1HPlKxaTqgng58mdrvbRqzWUzQItZQgSKmG4sGk4QJJsQFm
2V8kD37RJBldWlxwXaDh/Sa5LUXek7lLqJi13dQXJl0VfFJZxOV8dqtGk62jL6wH
WaZMmr7TR19apwmlYaEy2TaUBm/cSE5d+AIAnSuS0AA4xmZjinLAOmRfgGu7uD4V
q8sSUjTndnY7t1zLLU+2COiOwjG/gDvS4c2hAa9IFT9JeAzWt87YF0zaceWcvlMt
DxTZ2UTJCNiKSJe+3SEGzD/EjdoC7bHbEaBgprz1HCrQIuXYzW+Qk6zog9HFmKnm
1xbTJPfmmQu09MVP57VTo+/90GUC+69AfBous527PqOREkOwy4JI/nVSCWTNur6u
fcl8ZhXfDguhzxeiWDj81TBqEc637HtjmTeBHSEgMGikXO2bHcdYwYyGX0hYBSib
/+r0zNFCxv3yH515qulE6gnX5sWJRMiGO4tAkvkPiQtnrwT5tZSWv8i1Yu/viP/i
e38Ycu4hPAd04WhulOkEZ+tx4eiWWdvNcXsqc4hp+UL+5kKrm3UIZPaFd0KmwmsW
+rWYF5vBnGWZylnE/ztgITSyeBxuN4G3hOrjmr6Wz7OMEj42AxTtxVCInGcZ0I9X
usZV2SS8RIgArbCZh4EKKH+extHHmjaquQZeC6EzHHvGC0SpQa12OjU+EMajfrwY
bbixNn3o1ltGBPPhBeYkY0WTgBRSFuRVHD7CSA93PbvXvqxIG2VRKy8Zpbl5fNvF
IZqs3BYCMOnkGO57DvE0oTqBq/WfIMuuX4q769x8TaDwYVIsXBZBJ/uRY1kPyhCZ
/pLp4SoO59g+WGvADSSYxDv6PcQj9U8l2oAwP0meDfw+nf4SU0XONfw9+jJrOtbC
tpnGcrA+QeyDB2yyXNf/O+enGjEzMdM6cv7g69SZXdKsvMq/PI/kff7BhjhcvX3U
l/3G+o8c3ORgg4SfVa/gujoVWREcB+aSEauaMpFpid3FqB/8LwONotu2x9gU8BS5
gJm6kwYFywrUL6aMTmAENkx/9HskGLiKLnIajTuFQ7QR0ds7h+qC5NgW6zKMMn0B
3wOq1uV8OyuqjWyI060xPgI2uvuL2jaZZlL+WqZ6/KVsp37fLCNl/aZO1OSPxKZm
kC5+8GllwJuB0svjo8Fj/G90hPkgI1LhqjHCIQk1/cM9qdUVkcHy9tnB+gph9E7F
NFycp+aTfV4v+0eIsq6S/9uP2XWVqQSnBFwMXB2c4hz3svlMKyymX9zv873a2l+j
BrVCu9lM05BWgROTBSQ+52Lbmbex3E79TBWkqGhGwkzLwFca0REiod2XF9uQMEgj
TKP2y1ceiUbpHHyYv295sgQN6P1DfYFF53UOnQW/z7U6KejTFlpLjSqRv7EyXkNT
Wm+DzSIlehqwPKPLdBfGDNSbvF8c339nyUpPh3L18gsiYPiFZAzD1eJWZWIh5xWO
MIrysP7FFIdUm6cShiHpZ56AITkXg1UmsYiMXAKTw4gdHokyh9PyCdjKewIk/m03
/Ah6cuFTpcrjCOqXzQIW7UcRkTHID7gWieNt1MU1SoP2xKf4ob4oIValW0yqcu8q
6E7aP1EMf5t+WX/z6uN656Dnd1zA6xStSyf2qp7a9R6G3mPULNdftkyGF6YPHfvz
yiQlWcFRgTaE4RmAPV83NyyHJZvu6jjoi0GcRKAM1J9uSclazGKE+MiT3rr+ob2E
NpakiWA0c4uzsTgPu08TiAUs6aV/QKVXM9MtnUZRhOWsxqbNIyPSd/L0anbpKblt
TFelB1uonWP505+QP8dqLwVFkNSupSRc0rJlaAYuJDbUpbhEQwSnsP/7tG84jUhy
EVLpEJxwMHwoyRaLkRu4BBgm5y7MZGf4PzhV/U0qMwgz8JXhgcLeNig47eBAMvWS
DeNUw/C8LNopyWT/g8CLwFqszJxXLF6sRAng9HPw5A13oXSNAQ7iYHSeBUile/MB
NHX3uVEg/aeoCGVfUt2a0FLT9IEJ79SA62SGiiOA0OKP19YLa9LLYLqQDavsT9tZ
5znoLKsDi4EMsBUd/kLNxFNorSdfHaELf2hbzHmRU23K3SPEX51kbaEmWXIC57e9
G8BJ1wUKWPlD3mICmtKj4QN3gBL3npJF3qgFf5O4lZMP6U37Rhvg7lJ00mYS8RdD
hv4UW121sTSWgt3wcwttI1tvRdymmPthur+x2MeotGuLE8GW9IqooLcKg8GCqucc
rRV3MBRehAtp3SBUqD9o/0TCjbF4HaiNQZpVlMC8O+Roa/EyRrXsCztDv90YnK1i
hr0l/aYhOPcRHVl2Dc9VySX3fx/kKar1kZSTjGoU6o6CNvPpnPrb5dkMnEw50pEO
EaNEs+CjCpLrd25rYCB1B+6joE/ZDyftQLx4EfEuGNDWSLvmVXCZqOBZLxllTsGn
S3qQOC7G4SVVPtH2El+XutD9edkLJnSbrOzj2MD2PkCzweGf3yMZ3kFoIWpAg5Yi
5sgrG0gMKFiK7m960IrGMTVM0t6ztUCLiOZrlWTfy8JqXNgXdgEO0f/I0YMWv0f/
9z/H/tBdBcM5r0Q9cxTDtKF1AU4o75eAf0XXNpjoUBeSfZYkDZdJkdAX54pnZCVM
8PVDOW/rDY9ktZGdZv9uTsY35XFmWj1T86Br6zriSmOJ0KgaUKd7xAjwvYax0Mp7
ClqqD5Kp3uzcJvd0dMHSdgkkyNhsDmitLOV9lXyzHC6AvR9GoeoFmSu6O2J+isx1
dzyvldHeTp+mYr4oNFnPA0uvATCSAt3Tx1NFmtvvLMKheodMvVCH2tTB3ICifA3g
XM+UXgIa9rqF7OUDxKVVjqF9VTucT4RhR0t2nbd1JYJjVnyq/9l86rQukSjFd3SY
o/eU/auIuA5QzQWvpNnpMSBv/kDgme/82iHEwh6SsFS93k4YWjsw3D6sQnA18oUx
HXJD3pOli77RhjN8kMJB3ew/ognVlw52OlyoU3ieOwzXCWKhX/TUK9pug30tckqh
evesqPgwiNpXyegB6GbzEedp5Phi7wZ2uE7jmky9wuTblX2Q9S7nAwSy/uJ9OO5t
0hntV0e8VE7OpuUUxHXZOJy6vp+DO/udd5zKuQEJK6+yhj1S5tP/IOTJeISv4wq2
l1UIuIx4w+/42/57Br+uOJBjY+Q2zfujezh1PvX66N+j654X5CBKoWOsTvp/Upjx
b5j25VGPr/OYnW/ubnrL4eEQH8HGNuFHWsZwNltVXJJKXSaHC8na1w31oXEKl93T
ToqTd98+ndNyHSyzQHg3JVDCJIie/tVklib/BheCIWs1ID0WwhlKDri7FGiIn7ZH
CWWWAKGhLv5S+QcN2O2yHTWKbw6LT4zudU380HwfLTUXKTJp9g2nvqFugAXVG5zI
NpEPba28qkYSlj3M4FwYw6ICGuHPzyZmqjXVu3zMlev91fR4aWAo1kN8mpRNc3oA
tYvjf5lLi2TAwZd0yLarur/q5jQK0k2kC4kqgmguyq4hMl5tpQOhD79IO+bcc42j
ie9jMejUU8IU60UiQ2jlUg/Pjk4G4BzmePu+1Xg/zosMtfJNVe2sIzMrffQ69vml
myt2vsAwUPoqCjhJd0KxDi7F9+uyt3hvgathN3+uDm731CEJ1GqxSFWTFNaeWON+
8GBRR/9ihMUkP75Sv+MaiP9J4ZdmI2H812b06uvDVHCJ+VEpyZBNkqiz0oM3bFBO
Wb5eoD8EDiM6JlTBu/tVuvL2vE04kVk28Abcry5TRpuC6SsY5+Xy21Xqmy1JFf/9
DgWQz9mv5JAonh39sskYIZYJrzQGRHqVNG0ZCeg/J+U9DTSHRVAUeKo6U2wztkma
Vq5TyiI+rfToYkR/DAeR5tKKkrc4t/veUS6BtDIoFiAlBszGgC4aVKUDq0EH+4sl
kjkU2f+6RKXFpFney/yakAwyLxaIVcWeAmfIkW3IyxdxjnweqbVzZPT71gTQQsLs
D4EMe9vt0yvfXWZle8eFE5bp6ptRO3joPjnzD2Ahz48lDBP6G/oHgRRlVMRSgUpK
4HT93Lj7/1acOcjno7TYhbkEeKeRRg6SNu1K7iyLKg7lH6fAMAJyjBrzTifBSFQH
7QzOmCVZb4D1DIKjWB5MpmuO1gn3sBL4nRAwCPcHIxcqFj+K+/ZryG+4J0q/LuDU
bm1S/W0JqG//I22OXt2See+U7Gtuut+JsoWgIzeU44Ycrg4RelRMTI0pKe92fHLM
4TgUAqPztm6Jmo2pqrpsNfho1WDU++mjp9Ko+lHBT6ezL7lPnOT6Ai+EW89Akdhj
4VSDMubNUz8954JgOIhpFJ3Eukj9hHHABKNX8XgeWRhIqLlMXdxibshU2yKD5XtD
rSjDbquhMm5Pp8QJW+YfZ7TQbtAJW6bbz+Wd0J9AWvH2M3KYM9LKnIdzsXXjaOV7
/0VNR5oylHRb93I5H3La8AGJ20b5BXXic+wC23QRhxSdFhKzvMvkBNcw9f4NEl9M
8KROF5TZRgtQPEWGPAvY2yyJiESTt6FO+GPL6oU6BYbUFErvwPbWyAXy6wSNF60R
c3AZBM7WqFSojVWbBvRalQoobECoiPlSnga25Kv3VkKGQDE+OnTC5gAZf+bF8wMU
WgvK4pPI+Vs/iUZmXx10ohzgdZFNftja7hKBVD1o0QJveGr0Xix6bk2JlmcHV+sj
bTDACBk+nCJLLnj6tJZJWnIoPU4OuTsUs3JUGi+IzPilb9XraVZu1OzVVOcERvZ5
/JkHDsZD+wQadFYajaE3VHPFPjLSksXbjF9eo2dcRo4TwDUGH3rGwDrQ5i5Uu1ii
8BwsFeer31jBr5sMWL8663WUqkXZI4xjuCDMr0nFk5k2Y4nBrPUfUzqd1+p3Imo6
nJCb49B+aDXq+bceGgdaAPjpKOOQS7f7m/Fh6AnFAGlUjNYBhTDuL70NHRr7zPPt
7r7kIwagp5DgwLxY4ang7T1xSkf/PZhfLmXk9Dcqi5Aq/+cjnvW7ZiSn4P8PWzrX
iI2+C3Uz8eAi00HuaQg/LrCg1Js+Y/uCuUPB7KP6cqUTPU2HusnF1OiQVsk8VvWF
dNMSMtMn1Yfnrhw3oSMkQDJW9g9e/qvoyxGxazK6szHYmyHiMl8Njwj2qQjbI2jN
QA6t+Vipk/NnQFWQDY9Qr8ljPpuzRunAMtGoSXO0hHhdTikh+UL/Lu+hHGODgBSB
EojyjeqeecOQZQ0MLpkJ4sS55nMEKKPMjIN0eUYJcZZD28Td+YM0uVdswfGRd06v
MVQhpaxgO0k56E71VEADHK+udI6pXlpdWOXnxW4gbgj5W+/4CfrLLabsspdPUGnZ
hxaWbWoOhdF6OnNgk4TM4TAWryHNvBQX6/3homBlkb+At+o0rjnrFGLRMB+1YGEB
m3nDIRf0DY0+S2+QlYH+GwmUkr7u0opX3Cckb2/K02CXn6Piyf5t6pCjfkPy9AtE
3sMpJJB8If1Ed65HlHRPsyHKKNczuBikrYiQHitQISBsRWiQaNCwpsSdUCrNaKNS
D/JBeHzibaUxE2Fir3X/ebf1qpM4HVodVKuJrXsTZf/616tgpF09QR9XZMc52b1/
+j20STN4+550ggOHcAu+BWquHaDH8wOk4FFaPc2JPT64ITb3Q0vP/TH8+NgR7wnp
pgxqp2z5QwUQMxypJ07pu/tvtbyivXh5CiQlqnwADY8lp1WuKS644GX+JMzHmHpU
NGvVCdlGNlVPBHA1gGbJGGy8wh0gqS9cYFpmz0Gx4rqOG1GkxTbhc81pkyqVg6yZ
rvU2wGjkyTpKDBy5IIEcUgoHOFyCiV5MUibd5BGxP0Nj6H0GhV9jSIVM84b30bfi
RGDUdcQvT9nA5nAmkeZST7sZ8Dn206F7tTpogDOf2v43x0XYKt6Qhddn6S5h/BZB
EL+3R0mX8BLvbmx+T0fxn0bpbeR5WfDg8z0rFTBJXilNiJBbS/3cU6RGqQR+qbhE
bryAAApCUtPFyVwdCDwv306HSyDmulvaSyW36BwUsYyKxiqnmGWtuPtIlSTNsE0R
vMOCBMQx+j4CBClMUvNF+mbnTidfJQe5j+8x938EIJxacCo23+9oHV3/w4wXULHt
uSuSZ6tdxTu6fCSoC4O2/YFocCkfo9iBYCfhRIU2fBveDS/u+T+QcFN1ue3NTme+
TJ8D0f6nhO/tR7r4rDEsyrnBD7lxjmxSTNSrj8jl2avVMt+Q+op3yIOg3SB2TrwC
TJsYuzoXZqkSVZdiUJI4Di6hgyQo8TraVLSLSy+MHFRwOvGWeeVbQi3nimCsVvkA
2lJteSb0vMJ7+Vcz83eH89VOFQqg6hchR8bpM/1BJhnel1tmXTaLkDiDZwyJ/S9P
P3RT8nqqqA9Q5g5p/LUMlzmV/2qXnoN+3pF1aaU+oWuyvEWOpc4z+4i8k5QgmWUb
pqSjyrmG9PS8wvysutpEBfIumjMsmwuta9ji0tqfuseZ4GJXZKGHXmTJdiL3JPVx
sLI9EmX9Bw4pjZZtt+PxJwweoqD8pnrxJ/PTlDQnB2/MERky51nJiG7mtHqJOScc
xfVcxmfZAcxot5Gf34VZ8WiVhggAK4MQfiruZ3PXRHUaUr4C+ph+BYq5qLEO3TXQ
rwZjfPz94NVSopQLoziGBpEwlLUH4Znm2Y7a0LLj9VaOgH+0RC2AxvtuNa6YQkRY
TEC/DJczenfymAMdrOPWOOmtnccfbDlrDBHxUxeT447J6zIv/fe1R1o4IFkW+lLW
JEpE2vJEp/PbA66pIXwoJCJX4jk59oZZ0NlpzwPQGtLUWxpw5pGUCQZotRPtQSiR
52eS3FVTgyrtbf9n3xT5cnC3PYtzwPce9/ZLNeV9ZewxbvWthDbQ7BdAjDahb+Mj
v6zi6tMTgjp7p1Od2zi5NLJPuQH9+4IBaprnBOY7ET6Fmx1sx6VzUvAir6FqpeQV
mrbMKyqoFJGoSNlipmbc5R+4AkT+Q70iAsCUrTZQ0Vv2BCxs8rMsDTVAYHG1aTnJ
98QjNDQR5yuaKwlW8Fk8rvERd0YgqACOVzIOFRv59OIGdn1aOYq5lsXyUXoHacR9
QzPHejeg6xLcQlbL6A625QQSvL4iu8xA09p6Fy0zI8yQTy15yw9CUXT8fYQeKSkE
HdrambebxmLXdcbRT8xvtpzS/ay8czdASc95fhUpE35an0nMrt9gopLKPK+Q9DjY
ned5kR6LcpZz0gq5+k+o79VBO6d+43OkTHnQYiKynkfbPAmcChnPI8dNT+9ZMO8e
repDw0dXnpn05KuwVKfSgbbDCaoLiA4bezu9BO6uUHkMXElzinlSOlUQX3Lwlyl0
sLvAdedH3Kg8xRJYSu5tWWBLl01AKZkJDocRV6VQYUduL91MpsyPPcF1FhNm7d7T
BO5Tsptucw/iuYdyA8ZLlD0pRVgEwooRx48qoJjXG/PjUF19qJKACjV98scRogWG
hl0+A9pOgdodSXcp+EcJKEct1YUEDfR8i/W6thngQ9B/M7etf4ipPxGPOsNNSH2c
JSdBu0IgIKYr55XqFjV7XQGAIGzFunR3gduJT99mbw4PqhS6AJc+ArCcO8/53ci6
OPKAiMkt8SizAafz0XF4OCHKa+VN8qm1VN3gdGwkxuuz9dny6g80ntrGt/vAiQZJ
h6O/0DlFaGc0NKCOK/LYwlv4PbLYV4b7UrQhgZF8hwwOhr4F+TDsLq4kgyJxhBRe
gDh2yMWEKG7eSLVQhuIPVl2ew9EUsTbsL9Wq8M4ABHFBtik+9l3I0xfEUEGLX9op
uT9VzK6gjgxXcusTxb3mLVJz9WwYEZ4b9o8NHNRL7xo+KBahCiRzzbiabO4WmKjO
JekWIZiW7D+MwlxNYj7J8mzKYrozCWfZolznNaixhgO8P5SNjWNUoFz78klHcd58
PjaFMZs6ZwspDibgEn71DNZB2CCMx37Kai6A9dji9j0RcZ6Pe3cn2rvhtPgIszI4
vxZmlmAGcIgCir6JkI87F/tKBbvdtA1BfZ6m9/9lUotjtImS4/8VtsyvbaP95i+/
SGFX3xaBDg5KRwNiaL575Fj+zivFYCmq0eO7Q2PFz7Cz03pSPUbj2mMhCFy0Rh4q
eiL3HUr47S2JkwwdrFZYIYS4q2OUl5cAC+C0UjsrXoODDa7icHtjceWYoUzv/G5s
34JjW1Ut7moY/0P53L1/V9UMh7TueRsBevoQ2TyWEmqT4fiYO5631XWEGKi5S41j
zT6If+G9AIutt1+5IrznqZZyyjrQN69nl6wJau6wnUv71eDXsZsVbn5YV5MY6cv7
5lGW0FyYNBt485FRIUzCargNw8gQyJXPKsktMb0L39ToqlFf0chMvXjRSISoAp9H
OHBuOzTxMJ6fGnYlJg97tGHn8VS6OCw8kflwlW3PQcfss5PsyLjr9X+PQY/4UYxT
F3bcwQszHZuJ1H/hT7ddHo8oPegg4VhOYlbjz6IUKkKEaeTWbsdgE+kBQDePjJd7
akmIYUIL/L1ow+ksDz4TZsf93+HSGwdqNWLLre0qdkhvS886g0Wt4F5KAPMQlayG
MuGOCzEGRXWRuu8NfBuTWu0BQtte5JYmclbH9Imh8PRC4/X3l+AsL6JqxamDy0bE
uMW1zSDrO0yTI5jeayqUPM/g4YjGMkfBYYepSeNmZBJkUCYYE7hioHbZqCS2iT4b
cG8OBGiYadBzHzrZ5VuUf4hsHqaSo1qma18i38bSahBHNr/i93pwyWgZeZ+0szro
TxFrfrLJOy3oVt6SMgI6a4dTNWErItySDglKzXtpzWCARyWYY8GQJFVA3YqDd0Af
U8HncdtmgUiy/CBfrT5+wr6/xayzDnShsF6ks8HVvycyBKV2QcMjjHLMiRcuCgLE
z2kLVIFUH+0dJow3q3P0Ogoky03+lWBD4GepmclLaelCGfpGmGjwa4O05pooeE+x
WYDhJ6/S9tHFoCYfNvXUJ7fKP08bBgSWWKpu5uCPeraVdUFy9q5Vqy7poR+aFT3F
XVsiuvzpT6gl4BJjN153EK3Qf5k7lMHFIfTLMBiFKN/jpr217LNayp49nrFealk4
zLAYULOD+yvyD8NBu9kOFR31fi9ZQ50M/oJTbBQwNH2TvlOeTaH/0WW6jwxpNjop
FZcP3Uj3F7CEhorFUaharDDkIPbAuXhxleCNTSTfkB1/x3gmYDiRndey7GDiTFFw
c9LY3a2gtmGcN/amqrN07GV5wslI3bBgkbe1BiLG9G7feQ735HflyCKS5gBpqWbr
yItbnuaV1pMAzAtnC4IvNC2+xhgSQwHf5G2d0BuzZyv7sWYlUyiDLI9mW5iC4rVG
gfVIRWAmN/kdJjeIoBHCTEhT5HsUg/HVTr0cECAUU52NRNyaBozvjYkwgXmhf7Q8
e1ZksH9X6qOqwiuqwoJpGEQ2YL9Jk4hdBBTnqBU/COi233nMiOj11tzBgD5nJpxa
OPUmjTlG/O7KyLOtsWCl+NQ8TS7mIBfkmTFM/Rb8sVwFr+xGK6EmlT2CJPOrz6K0
mEIoBAjo01pV//SvYTqEbECCCfRmTg1S0pmgg+oAN3eGekgzcVPDWDmUygAOJ1lb
/oal67SGV8m8SMLws7bXBQI7EWRiFwZCCCbLwRcvNl9Q2MHCglv7drA1tem6pxn0
zAljjK5oUDMVoNaTnIEFkdViFq91tD/EIFiJswETlDFQe+ITSeBw4ljLoSxdWpeN
KbPu5X62KPpcNiP+4rWIh6b9IUzG+mlZ1oJe/P6GXtDgZ5rH6Ur+mXwb38JgoQpm
orK1cpichazDVwQI6ycIh4UxcdreUL9HHN8jQEYX1DS6Qo8IaVFo0qv/QW5u2SDw
uSwrr+Gkjsbd3+29UhAwOEt9l1CiMXoLTsFVVkE2DOGIU47E3Rkmj8xbjW2/TKFd
CeytMCTsQ3WFmjpUv+0+4IPxwqG4Un+90mF6WMmH/YXp/3kAmbXNGh6alya4ctrl
hPF32PuOLp9oK99Jd8ZY5LZIQYk9CkA7PssNsr0mgCzX0/xEAnnDSNvKh1kEJYcW
dP+E/Pd5MEr+HKEvri9yCN+p9r5TNFDVYIqsc5IarM6Q7W/DaKjGIRJ5LTwauOyt
uWkl32Ln3ixCsdILZ6xJzqU68tjWEgvO3yITXzX7u3kyXOG8BgiLflcib02oyuTN
rH7mwPCCLeXTqlqBVk0c2TQowqAFSda4Lkih/GNp5PQrEVrRo/7ViGMNjMtTbD4H
IUUjITSPHi1JNROpKFY2AiFCnYwYYyNeSINze96JE8tgIN3VBRan5uaBpQ29/ayz
LVCMnqHa5OXQWsaD0o6OHANhHPJTAGvuhI775JHOmnyKJileP16d9DxEbqsucF8f
BrdEe44lZmmQobqMdsj1+bKuF6ad/izMk8TGi3B5azf8FzDG06ERGe0au2PUziRW
4Jpuj7L4HuTzxb5OpwR0eAPlqq1SKnV1d8CqNuiybIAr1Ids66/pewBX8b2FbE9/
i1Nxiv8S2gIF0VzJFqanxuvythQ/3AScbHb5ewp7jFQOTOsdttoTG5nAb9svbvfW
hY15AydoPubsJvp3t4FZWipt/TjoTja8NNFOHp9SohPHQF1M+new40weNv789r2a
fNShcBJz2FOgkVZqg5QTo30pSCEXK/SzpITQS3uO28GufMqQVYuCzinsAJ4QGCHa
LJk+voKwpLRVW1Te5AMZhWYykOYZ3m6S6poRfJT/Y4CpD4VROR3eE2ukXc3J0rVL
aac2modDaC7cTuleGKyVk4l1tY9FF7CvZk2qboeBwqedA7uKuuu5CC9FIR5X9fLW
pLku9DJRle/hYASJwY6mb9f6NPZL2sSjVewZgjS6gtMDztG5T8NwMXMWhwHgwYD4
GmH/zQu3ajdzGQDWS74Dj7Ri1zSe4IhsqX/IzbGyebGq0Hld2dJmiwiLfjZ7w5LI
PrLs95DKUB2kIfeU82DS9fs3/P9gOBYchrGJWOcJ7tjTcPP4ZbZ7r2rSPJJr9Ltj
0OcGTzd4diJkaUHfOmMPMfoDNAgQYsVbUct335eduGu+hW1e0Shy8ijrFbgn0te9
T4a6s0A+d1TzsWQdn3Uiy7SYqbuiddu3qlYklHHa0OJH+RoTRWysg3jjeB33MIeU
wW4utSx67nfOtA+zVrDBICKMQCQNdoT0jevkISjwJh6t/ZQsR5MTUzemYAiaGCGL
YPvGhP4z1u1W5Ezz3WV8F+e1lDMJqnwSgRFcJkkhhU4x2RbeOopVeTGZrGQoxeHq
i1nYg/eWVHbhzKcjgQeZUQ4GYxTPWcAFmhGOimjs3nyOQ1iCr20NPStQHcu5Npky
OPL83tOMtpeieaFBTybn+81RmwIocewxwbdV1dJ1xIasVW5sLu4B1ngaocR8lPXE
q7DT523zPeXrWpg8nA2/KK+36fCnIKCPgMmmxWABlHAK2r72CSLspZ0WTwgZHv0s
TqRNdhsp9e44CP2mnkZnQmlcL5pw/9hxU5Z/HjZdbaDHdlwaJ9XJRQNFYnI4X9kM
oJuC+CQ9hO9pj4Xbefox1VxbpgDcEpguga1rFcQNkCG8Ltp4mUpESz3IbrSoqXL9
U1kuMoX8MtZ7Cf27B/L76jXjWL/BS1vObs9/A/aIzGLjmfp/aU14DazAEQPaMw9K
7SR8HPqvFmgHsLttT+NaJcu4aSXJ0IcC7m/iVS/XmAkL7Ck8wPMx6fFnYthjEjLh
n6bHcLlSUWHxoM8Mg0csGsr4FyzEWZQ5UlcyGj4/JlM6sjrhHOB+U0KjKkWQJKIk
kg9cRdUO1z2v3+2S5skFl+2cyPaPSLK64aVDrN/n8/J0R0w6pDw6c6st+xB1lO3z
R1lGpicb7FWEZpY7p5lK3B8cAW7NOD8ZDJZBNnL6Clr2PqRTwaH89mftAjLz3+7c
sKEEg8P3mZbGNRtioesg/bEvBLUTBY9gEM4RLJptagqyUoXC4iv/sTtvjARyyLAN
DPRdsk5L+FcfoqPhynvEj65/vfuNVzkZqpFu1JCOahHKTuiY1RGbj6zAUPa5RBo2
KESOGx7i2uq/8cQpR5cLb5hTlqheuIZSf1aYjhm50v+9OzFm1oaD1fbAsbHuPYzf
g140eMxZP6DAxvmAmxNNuWjbEoJMQk8ytcJxvHBTCNM184scVWpdy9FqfAOY0DuQ
ygPl+/7j80obKT9kDur+qD2v/uJrqprzGLaYcEKiBNQ1Z4jEqsF/uCbG/icdmUN9
ODRHhIwXT5Bric4EXq4V7/GMOH0wrZBW1esQdOy4Vn+AfVOMeinDeheRHgbndmPW
6mGkczr3X013uqB1+EHWxgLUvUltYSvVmOhI4Kjm1PJ8SCfyAjZ+ASIiwOKucCt7
JFrZmBmQV6akDqB9sJmm6bjei/njpXY4uu6EqTzgvmtUNEMsyy612qaK8/oaTToq
3Egbne/oec38xLToilkfhdUl4Jr6bhM/hnmjWFMaQLxSLw35n0USC+IEnQ6Qxqrn
3Ob2k3Rt9cJAGCKchHEbKTQffSTCQjmYWchQZEQTyMFBRRVOBqcVYk+LWX1Z4aUk
jw6EwUBJ42EhJmd5ZaFTiWAJyP0ZS+63WljTD5m2IsPQ3N/p1wFcY/96EZEKxWzH
cankFLOzQP8ynw/QAOE4Upi3+aXeUJqDpV5dj56tqawlYOPaTXCPrTeCnPne7m0X
3ftMvtf5sEZIJ3b6wB87J5SdOEuu5Hnpzx+VVPuphNXeAq3VZsOxm0Ws4EQnU6/0
KjnvFJyr0cRTnwYF0p4fe/saeiDaneZAGjKlikVPuTgLXBQFlj69FfGrjlHJZMJa
hv3ECJDu2X+qos1uqYkFLgRnyyt6SM5gJiwAB5OUyokiLRfME+hi8ONqwflep/tV
2C5oBWbTXF6wToATjr0Ku7ZraCVz1H/f3n8mkh9cCKK0/0u8AjYJTvKzmynEWNHt
D4GDKuoyfPvKsyOLyAnPSFGu9PiVUVA1hPmab3KDDmQ3k2Ou+V3eHfciIiZDuB/C
v8GUor8JIecBMyOcW9f8c9LBqWDEIVOPehEtVroBVSj7tiEwfXmUXjks8d2Y6wuD
915phrZ030SX2YIN0rJrZ2sHxbaX6RUJ1Xx18O/+3i6mEkxOWPVF6FahyLAGN4Zq
VDffK9+yrh5itFlgqdvnW6WR2aH6S6ZBQbSP44Ks4IT5YcU9vzMPHQmByP7X8XFh
YgkkHJeGLYMSS6m7MQh953yJoV/kqgNj1Dk3Aqhw3Xhihk4lBIFvKArWvalsLv/L
vg6GseCJKtvHNL9LPgMmRix6/pDhmhUkqBu9iwaV69tIsv8XL5Bwv/KHS0kZSTx5
xyPmd8PIBWPvs+uG9k1dgxU0cVYdRt6ZaOjuWF/jEtrr9yrXeAX4HAmVvDcy6pNj
2RVdXO1tZIsSB3jdwe9phFkNwapbNisINe8/NJjfagtgJ95w2AlVTBlg4H4Mxyjj
lKacd/9PV5+CAd0jkG+v7jbPtleq6oI6ZkTYq60zkWo4wfCvAAviwnqEp0GiE1mO
5yMmer6JaK6ksLM2OjXX5VZR/hiU8Hg2WTGFTDUJOIHpPe1UQ4YTm9Td0SjBFIgR
JLV36OTbGKK+SCCxbxLXql8ryeKcUxV/eMgRmdIAncU8XxYX0aeBeBTFwJupfzJx
tbuI3jh5ABbENmwgciR5Wotb8xwoSEY/2+rkiuoRMQ4LTi/vRmmCAiSxMchkQ2pf
0nc3IY8zH9doTlPToIWJ9bd40Zv2rS9Zg/KcncVRIK2w82WdnoMTHEYSnfCWXOOl
ux5mNbWo+/7x7ZyH8dJV8SDIAfnTg9pzW5zkhIOUV1UtJ1hc9dN2GCzcBijOpY50
zbii1UoHKMQ9uM+u7lGAHDHc4Bz/gvZkVRKyj+RbMmxEDMK9O+M5jhS/td3hmDg4
6vehKEm9r3s5Ap2+bGCnK7wn4AnDYP5tK8Gp9HfdjQGq5t05VeVwhBEpCStkSKN7
dNKUnr5MwFJt8ImgIEd6jeB+VLwIMUj/SxGOtN1biPlEhsqutUjbpHoOtdiaRIKJ
x6gHhZk5FE6ZPZhdUFg8ZEjKw/yTLXrmo98Vr4H3Y7vXKtOQXUoJbsBsSubFIBaQ
kfROYQOKsC55MtQL2dtHlqxOEQ9Cms5WsMoPQz7Yhq/Cor4eaNx5PJBLyZ+8YYzC
XPuAIojw4Kl5fWnk8Tl3i22evTCABfCveTdLXdKA1bFCnJqOf1eqM4RB+Gq2XiH/
A1L8nPjhyvqPRepL4kSbhZiOuiAvGuNZrDnGZfWJjjzDorgfeP2bqH+boG1WLW0n
TKODLRuOBFPsJBFzy5Eny7YZfcHoFrRPO0T7QCpOnIlFT+GqDg9tIPqFgv+2JbpN
yH63IWG8AauTuQtJ1SUdocdSrnTH/3WTkByYGVT/uN5tuOAZ+eeJjeXSoUSi3nEP
yJrHlUk4PUK5RRMXXKAJT1UtmlfTAzhEbJPm7StGeWOmqdKEnoW7FzmFRr5k38hl
B5qToTKR1QxW0tBSPAVu16Af81HH0lpAMo+9PMqfZIKPNzeHdYvzUZ2U1kiU/oHj
wSxqD9ywrOhpFuvtZA4LUw9a1ZMDzc1LeTT7XtV1dhQbdjGWZnvxwQQAyXTrpdXN
OnUzKkiQbnPRvuWv99faHVpZfPhRDo/upDGvwkgzhL64DPLHEsgolN69/b4ATImf
4PXTJg0OdFBYyRwxP72SQBgLvWwzw3rkVgMtdBL786MillMOJV7WuTbdV8vWfbBW
+MVqJlrSFlGygzWZkZsd7ZlvNxlGS3OhXJOBAb98aLvec3IphFUViQRvntbU2LH1
t6u62BTKVK+Gt9Ux3sI2cgj2ynyCginAqnRF+KLhP1SeuFENxA1tP8DQOmLwJmY8
POj3PWWciZcam05GKx6UR6poGIKM3fVSNRq43OGulQs9U4539BBxjmR2WXEehTnr
M+QzYsxvykYnz98/zVpbPFHneIa+w07L0wvwYuOTRQg679hN3PozaEfdTftRNQIC
JkQrs2EcUW39PUelEiQcYqvC0+EDMObJmx4JH/z5nvhlTtPYsdLnzUFW/JCiGmfP
xRkp6MJcHuq8NN5P3QWUZ1xAk/Hki88LzsbUkgPahcUVhrKNvo5zA+oZjoX9MdCj
sUru8KGmu4oDAIJU9Aj4iZ0mhvg2BFYP69OcOif56SN7ffvXKN28V2vqfs7opk92
iuOzCBv/LGFHaNNdF3/jtzlmZU7dxgaGGGuU8jdm4Z/c74cK9GmGJhzOpRtYF1Lw
RS/jztecjr4IPSEMYBK4rU2+JLThKZLQHwSsmqCdx7XnqQUViu+j+OGO4hCl3gdL
kdtnsMhZCE7X2msqlo6cTCVtnoEAyWJC1PGnKA7Cqj5NGCJCYFB0S5g36Kal0a22
FlsDjhEkC4UOEDtrN9FLOMF1mZZ9q1tCuoj2DvnFN7N59HWBJEfmF/p/t6WGLCz2
GO7MyNzOdFT8A9JFj8QWUvTMzF82voAbAtN1gaedUWqW21TfPAxtA4bASryPfn2q
PnZ26TFHuUcr39OluM72e7WJcFhWKOZQX7pMqskfMgUFmPdu1ZdIUa6GSNDasHPZ
K8L0T6JLBr9+VxPaBfFaLH7MIQRuX1FWCuI1/TZ1pwubKldut7necBmNJymsl/T3
GCHYVRY2ZfMrSprq+PYMaQmyzEMyUsi48IulvM+MfE0eataujUWUadvJOFTUmy7a
Xch506SLlUmmf3qlFs/NnZsM7weYZjWflJSDjFBWsPmnRhnyxZDX5ItaEPvyqGps
YEp2OmtvsSTX2zy6lXj2W+RjO3W0rTUxsIt17KV9MdZ0hfiRGHl/HsjP1GjFD+7y
K2XE11HuQcyIl4dnim2+73m8ZelZtRZLy2aH7TRbsK61hiui64BMd82lnk4qUw6R
ovSe5cIj7UtvlGQPfazt89bsp60SJOsbvJkwEfLDhckYkOwA8YD2E4O1t3KDBSd2
LfgS6FK0H4643sQ/NgKQSjV52jUUDEFKVCv9bssnzjRNMigBpn3ZTYFpeAihm71E
1m34qIUxC9sFnnc5ox2Wbr/BQZwaGAbOdLczOupUEeP7MXBiZWAIZBhn2lqHx2ey
QhmUmP5cGlFFII/SiYyA2/Q/fhoddovMzpxNVhbF0hKe072F+cpURkl9Be5QF5J5
JP65yNqgTCdFHK62Crudi3b2xvg/lbzPiKJO6MPzPs/cz3VNzm43CcRcJS5tv7xg
SWTYOeb1lKxOrY/tHagdYBO6kAoV9d+BSBZLvFBt+blK27EUV3vpFJHNrSS5BF2T
ldmjuHIitPg0MjNJA9LlwiEjRnBAUdai3ike7ZOHwpWopp/7T4O1+w1bQWjf25pr
hDgux7GsmUtgl3SXm5aaLh2+Q5Tpv9fIKlF/zM95VEYh75DM9jyB29tTuxv2QRmt
UNYjLl1apNMeX3dbm8VzC0z5ROhy7YjC0i5GIBEa8XtHxFiGF3qNsteqMG1oHUlx
9xK9fdaJ/eb01uDCWDlsXVqp5bnNOcVRzozXyrf+MHx5pKUvJ1bUQu/x7w3fmlJN
LmI1RndF7vi9tBfZB5XTHoe5HeuCjnTDKHpwup44rWJmUbiEHqppVQ/nF1MR9QTe
8u88xkQnFGpvkKycGuQgRYbyadtNcqnq+Mdx4pq4wWgsrKlL+eCdL1o8zexp3eCP
Db4tbiaHVxoFruNPaoOHPPc6N3eLtE2qZEhCk6lAkW204G+iTEN16XUsuwppD0Z6
tOKW0TkY0puZ/9ZHppcxVL8hzNJBYwb+D5++7g7pyIZxWB6XfrqAiD0F8AKLCQuw
MV0NjBpoLJk83EWUDsGMFkJ/YM0SfzKQ+AQjtYbgRvvWT2IPt2CS7U7NwX3N/6Xl
QOpHOReDrHo1pOHRzFnbvO/gJqT8KIWcXS0vdRD/1weCkFJ0aBfmj3jhNF/ZLwG9
5+v8jbhcK1AJ874totoeGSOefEkJUqp/xpvNZvXXcDMZYGxo3ENIBbezDfmlfG6Q
dDt/lV8L8rVKVQxKxT+5Y0FbpQ145xjDJROwx/NjQAWUFWKzIoP+0cyubNTeWV6D
b4IZQKSUaKXkEAqMSwx9EVGIaG7iZyktgbrI62sYDCmj2P7ObJFKt64WyubUgkPZ
GY4Zuzm3ZcYXYo2dEZ/ej/oyqhgkq5+qHjoj9t+2rIU35mcjglIvzRsSY1usAgv1
3+J7xzg7xygyDcbFoic3A+Uo3RwqTci9zWUysn264W3r3k4ngNSEjV2Bodrq6HW7
BBQudcJI/tZMWcLnQLLnYFwv2jelvcSv0BsB4MMTm+WFJYd9u7iiu418CEMpfn75
JHMzA4YsLinSHGzaLucHeatVkId9LTwtSBmOxPmscMPfO9DdlLquATTPOGiYNGGl
5Qmo+P9K3iCVuIUiYb4qsIRpbVAILe2Q9yo1lwIRgGzs0m5j6AeOCpTHImnB9uCM
iFI7twaj9Pwxd7sL0VG49xlK2rNKpDV9nk4tG/FHYlFjbnFbAgliVM8lUIyDuQv+
QRYjZSMt/2et1N1/PG8cnmjGCNKh8T6vObKEycgv1KKZ4NPu8nhix+Lg/TPudwol
O/0PgbxC/Iix9oH8/SY9o8jQx5d3RU4DimCF0LBcFsx8IdvL/Q4tKnLDYZMpl0P2
dkliUPZZkTZs0rr9drZLdmUWPQ/4h7oI/jnVU2pqsB5nxMtgiduZI3wpbF2ZiNBl
7ycJP25D8Qytm9UxiT/YNuWZxeGYnnBZCu/zzHAmSURsGt7pedNZ9yFjqho/5MIk
XwChRzGEbm7yq29imWEZ0UF4XywK6cklPgjSBXieQbVTlLXGzhpDAOQWKq7/Q27O
QlCURyucSR47NOPFAVuDwWI8dDg0gt7CByOTrid24fC+5fBn2ME2qVM4GWh5Kmb+
38GPy0Q07ZgcSmwvPKbKmDI1xy6iNzGbbR+ipuA//CDMNNDzGNjePJtfYeb1wLLD
UmRdsvDfBXVDFJuyGi6MSAA6MihMQNr8wccaw1V4RECr+5YX9HEMsEBLk6AXPNM7
0cGNj6DPWukDnYRZNHBJnMI8OCsp8qt6ZYP7nKlqEmaYGNBjYqavZ0X1YbHU4zoD
d22fR68nnoFUmcEBwfQRHSbHNsra+ud4eezyuGHJ82H/RA8XHy/4mfY6dBamcq7w
+UC+pKfKGe8m4XMXyyqr1z9HLh5287AvcdD0NotqHJolgf1/ojhT4XvMJELqCbLc
v+raTtbC+laI634gklOxm8OZLY009PlCK1s3e9aNeTqkcM8eN6aKxPpOsTXoS7B9
+vzQshunAHwcZz3+4tfoVXELxyanNHLs6AmXJHQRxzIwLsTObwNT56sfXuS/gdhH
Wlp2gqFFCBCdBCe71XKIu0JX/v0lsvTJe8yNeJD4ez+SsPD/Nzy3jlBCFXYmhJmq
xUXc6EEz4PtNPkEv3TZZ23LcYd0R5xeJLANkLi3EqqFOG49Xw4ZEHWjjQPPGKF9w
9Ji95/z0oTAhBvYPL4kJumWXe0O/7Uu/V0Of2OeYV6u7Z+Z6xZu8gcdyoKukhMeE
xqsy0rwZA8SNRgIeKaNphnkgy69juH4oRXfU3chEcUb7a1mwoONStpX8G7di2VWJ
mi2jxq1ocoYn6PW/BQB/KVp4WHhs6NdHyila4jkonfxbzOllpFw8x0OP9ZwTnJgS
o3jyKZ03Gd8u1aNLbygWqRz/i+pQjOZCl8a6o56NZIkm15S3FlUl81Tcld2xLV5o
LtjJDivtehJW3lihwEYNzapOSidhwODdNS7k3ZaJ3LyIScI5e1ulFZzCuMTi+AYh
5mgCxsfS1RXznVraWIO4975TL7ZJZdnCuHQovuSc6dRVLLHW3j/D0tPEWfZeZii4
OFo/vGFhEFCd2fb+z51tCtBZiHL3AG+7riF0UxnoBEAxHhqP84DCUCmoG62Jumh5
WLD+L11sW0WYHKY4oy7e8Q+xILyk6sB9DEyNTF8X38A1+RwdcfWruC65W+aunfMA
EUQEnG5tq8idDOdyCfFCGPMSmONloBJ8CLZIIps7ShC1MM1HaP0Cy9JABgYRHLA9
oI/1HlKBrp8Ko9V+ZVxMoGYtu7+g54rcomds4EnweOldath8NRiDFL3gfbZQnGEy
ILVo+ZoIWOcZHXnqzrhxA+VLYV+yS9M9Rx2O2W19ZJYZ2t8QN6XNwwJwvEJY6law
KBikswSX0MGFSHXEVLkvbu9AynsiIeUmHdaTjEP0RQdD3tynk6WpiRc9AgNfqxH3
/S/ox6FYIBCnXJY7D2oqxOnL3mp21yecbIKuxvPMp+wWPdFUeLAaZJv/iVDgyuCm
DwQMM0AgsCCFfFO9utFohNjxwaSNhymm8X7d5Yva60zussxeNfo6pRqmpnhmhY+c
zx6s6PYd4GeAdL4CFywFb2/v3E3i66hmUY8T3uEzIy2lokeoeWQJZ0SSnY9CjShA
GQFo9hC1YmJ/wN+/iyU10SSmyoUGGo9UDa3P12Fx+ROvVzkOWNDJ1PWKx0pcEe25
/wtoq+thaUelZojz3nLJEiui7dhyS/g5sKlvd9Y+FUCXVx8uS8vVntiDOz+q1l8Z
IZGwNPUhM7REe2+cESVi+/zjxmeGLaPrvSIUh/vaWcWWRHUQKW4Amg+/bB/O7J21
/Byv3BL9pIW9YvucZeVBinar0GDuzlX2zMik1AbQTmi2VLhOaQG8VjUMDhy1yPME
fKG0V3ErY7K1QczK1b39+Nk/MesUlH9nS9KUWilR8epXIb60J5VMHepNU7OAlxEA
RJK3mdzX4/IKRTT8xuOJ1lleUuDC14RubvQ7yvdHUpPy7gvmEwUNRjl62fThlS7B
GgqDpLWaBoNWg0YmkJJ7Gqr/X92JkgGbghcvYJZAchFYvB8kupoon4+wpOEEL0L6
tjCu4jM3wZ2KXEek/E5xM2Gk7NVb4+H5h4FwAvBwSydR8d+dSj29zWdxwT0uTId8
GBfyNXbtgTWsEn5TukSifF6pyo4MhOkFr45IVcqKyehf1xhZtI5HKLH5bl55c7Z9
oye/Ky3BYJcCw0BDWLxGeEklzrFqXBapA+988aLaP/a8KbfDudy8qQ1aHqqHKWkN
6e9HGwEx+sST3HI5aWvgcUGTnrvxb/aLGSX8cBX0DGOYTGw7g4AzADj8O1/KCpAJ
nY0mchKMe5OK/MYE3oUm6HF+Fj34LarDjJTQX/FkoQkMmN1TmYiQBvlhVESFvSQa
9fzh+aIe0GfJ1sLfOf8oDVhq6Btu0buR6SjgsaTlLQrdIRXgI2wJmCCRMUj9ZQLc
AzNX9xLjFnHSC5HJBnjyB1cPK32tcOGdjIq7OFgPr/SOMMIxg85NaTkr59SniHPA
vA1pK8dE8hgQnqKKGWXVCUXx+KIupTP5N64yfeFv9LGZsHZTHTFx8RZ7S4JYSSpA
XLDhja0IvJJUN8vWu7mM6hFv0kH7GEGaGEgCmVeGBGAiRrvU4vJr9X/hCSFtsSoV
yL49V4l3tchLIAsXgddd62oJoQC/Tu8Gsa80gmeY1J4OPgxRt90fQBqoBung+2XV
BMNxxvDw5BrqiWBmfEJT6WiaVmkrczSuzLyTMRk1AINrJmWnPEMcw07Ywp2W8RPs
WcR4v+8aaUfFgq2NBbiJaLDTIPdNlq/E26zCidlmFs1qPVTPEZhYVmoVZLn6Ru4l
FGsNfiojiDxjSTTWy+OVzn8WJOegxQDPcbKObwfRBhcSNRRSpwohiCkp97CbTxYZ
/xfGrW1Z6yImFNS1GTv5n5wAV376X7mO4a0K2ZupSYnSwaA1kI6Wh8eyGqJaHOfy
Hml8j3TC3AiRAd0QzRC9fPbm7igjZnXiWQH7QaTxr5k8YVLV7oe1mIRUoA2ClbiO
N1lYmWlW5vVeknKJ9hXXl3ZtWS5zheVfVhVn50XyJ1uRJLv5H8EFjFZ5RBobeisN
y+aA1ZZQQ6OlGnnvNKCCDgbaPZZtAjhf6GlD5wow6FF3UlO1E/QsNxiT6wumq2TW
4yMxYQmCRH1NXUU9EsnjrnFb+cCv191lUOdVPaSH9xTUwAf3WNGqoeubDrfIhvaI
4U5iOIljJ2ng9WiQBaGQKDC95AIDmR52/rV1efCS8xkU46klmsBYmm8iSZQyolVv
JmicSF8eyfFNLEIc7tWmaeVpIlBWxR5OEqrhpjIiOBQGygEmU2ASCadvNQO6/W7L
WVFDmHWV6PKVmKvbCNRWfpL9FV88Hge+QmuIpuxPo//dyPGvr/we1QkT4OzS/KT0
6mdbfe2RLZqQtMQ+rFZBmGM0df7SdPJp4/O9I4rrTOIdhAqnLal/GauTiL6YctJN
CFNM9nNQtIonvVIkacfDR7Mq6SM/NGwYD/L8yYBNQJmpoc4YObrCkHaR2OfplIAl
bUnBmGgeJDp0223k0luaLTmCwzl84unOIbZpmyKKAzUYcssd0oevLM2JhNKAwOyy
1jOKpWQdMWy1nx59HL+HWtfF5HP6D1Zlbn06icoABFAg61bi1cA1cHV6Tk7w2VKh
iceIjY316DDeGX+6wjE6pdQwNO5MVM4rxbnLOAktj3q/t5gn6OHAC8AwaeaAfgj9
Hx/klr3fb+hcFsQsnh4MxxGoY7BSc9/vcvQ2gfsQ+iaLy0EFNTgg+Nr/jnWvT/9p
z6s5DcXeWKvjGtjRelMtYzRTts1p/nY7LnogQJsgXg6/cK8lDLAx5ecDe64D3cgq
Cv9O5IkiWHnyzoUfRsD3+B6tYSbfnNnOCmFqRUraDAQ47TjfYYvT5kRiCQEEKuc6
r4r6qCFm+ML2VSWTCqLaTcSnMIFMRiU1bSEziVat4+OnlTqAojPGvQwf3+z+t56k
ASNi7wxxSvSMjPtjRkYIEy1U6bLRVKBUVAUEgseuDedWwB5fUPWArEb/SBImMRhp
1rGGLL9AjjCAV4cz3dkBXahp/0Z/KWuhPR9BZ+15XOikDJ4jsgwwo86ulAi78+oy
ZNX130ZDVRiwxhByMyfISoS8Glut8HI0iDLjQrZ5cXdb24/P2YqVRQ0dDYBb3pvv
2s5zrDOvXuzkZbXd0yTWc75PCbkPBmPSVkM1dmmO2wx1Y8inZvBHhCftLKPr/uDs
atLsA9jcFLz+1DmppIfFuaSfu0NIgks5lXTOSa+UqX1oz1o4jOs8Ak6s6TVg+RS+
CojzyMmjtkvbvsfAFFpTNXhznUD3xdFQsq82FdNFQ8bqlBEBqMUbMOiPvT4OIQbo
fcHM0TG2a9rIgjGCwfDQ7cH/xYlXS0hgoqAp2r6Ls5SC67KT6hh3Vh8HpXEUxYo/
xsdGon4njSA4g0jWdDpPgObJa9wNMArjSc1Ba9fCpl+aTHJTjdA1KUf9T+ZSe2dB
Lq77/NFd1DrOYBwjUh82mGG9O9GvhnrW9zOwv2X5D8XLVyPMRkipFKqYe4Pg7UdV
iETyP+PIjaOvXCPlfwbmMtUZ7OWm5Bet1RUyGsEK9Tanrj4kVctr6LHuIFduM+sw
P61LKTAC+2lOX7odYi58GyWYsdAA+vKxDdbeUp9oiF65NsRANz51ha5tgJ3GCuSt
8jbnzhd4lQG0fBjdeHAe6/NP37fBddBvbhwsVLJnd/WmerQWUtKwsNCT3atLpTW3
SdSEFMuoDZxnMVZq+tAWojUp5Jzdc0lyJLOCooRtKJyshtAQwj9WjDCRLhqjqQeZ
ywcuKk5yLfBxoeAhMY47XLo3WRfoTGs3qPkK0TDTKyuCTDOEGxGAKUnGXxuFiqCX
e/tksBoIcgh/H4GHnwWJRrQ/gDW0w0iA2WHh78giLj5eOgoF02i3cppXMAwtMYGp
+Odm2xGXs/PfQsI8rFb0/f40OPEuT9e1PW5RsKBlSzuyArNAR2QVIWe2Lo0ESs1O
hpyxBVA057Qg4ZXmxZRiNIaBT++EG+yk1lfxS2z2hpBqxMd8/pEbhCZAn2VA8xQs
BHNdt/pcaue11VFvUBYYqst8Ta+Km3NWJePHDz/6eu6rq/tSAn7QKQr3dZKruxm8
LxrComMV/TprEpDrjdiBiehfGOUE6wzZC0VoyfDQcgqXwmuTFd85P1bWSrfL+aiR
bqUTxetPweOBaY0xawQGyjC8qMPQ5JfzYnxY3kHFAp7a3Brvl2ymVRqOTHUixyTS
V6lJBlxR3ZXApwpNbX+BrIKmVvbmG6Dom6xvm2fvI3NWXvhwzHz30dpOp4/OMsbh
s5ikkXE0gTzRjB090EQ7oTHhAk51nGZjUd9R2Mj8U6WInsuAHQ9qVOFaES4sceZP
tLspykCh9He4isk8OW7SghviXbuI2c+G6uLTecLebrK0aeir4bTSQMhesy40WcJx
g7wfKrZaZ6k/30ZB9AvEAHxzgj1x6n5jsQXyb3ECxUtK+eBUybva/A1+LwirPGMB
I7zPGA+Z7mFzmZwOlbPEdK76HFd2VSdZU00v540/1PS556ictXOSvdJdsG8aghHV
YtoZG5L72iXZvGM7ISRe9X0BSN661MK2GitPUijjK540/1TA0a6TahvghYmt4opi
OQsCnlNNNS91WpEIUNc7X03pOG5T9utdUyKcSifsSlkH0HflFguaH47Z1Igni+Cv
IrVMP9XHsSIra0Mu8L1Cu7AfTx6YTq8ZzUULw2WkZ+9Cmaxl5MBm27P7Etc4VF5a
2/2DRAcO1AuIhYDbHBXY36FLFtb04DOkAPzCoHiK6V/p0V9c6r7FLzLpawe4np2i
CprtaOYXc98qT0fjQQgrV0V3i9wCNZD6fPYPJ9brqBBWmGdoqzs8BWz5K7mpHWNu
StXF0aZBqrkzkW5EH3m9t19nqrsST1vwyoZg++DXdO9rpRqGW2iv+xgdjY2WFkRR
t/WfX1ka61vue0KwE26As37dGRWrJV/7WHczt39Rlh1KaK9ii3VB0J+7CDfcucoS
gCpMZdIn4NaO05d1Qs0bXeC9LKzkrGzvgs7XOU2iboIJh8zm+bvFWDtX6LSn3rdX
HXSk5x2tzvMUqRd+WqMWWZsCPZkueML5cJzq1ttUDLZ5ESNUJ0ZX+7umVKtxEAq3
wX4oq0utX8wuHmwRlz1jTI021SGei5xdJc8E9v08+jZc3lB6ZAFQpvu3FmJF1frK
w1X6lk+GxeiRuEzHKgnMnw42dgR1n8kpo8BmmKvx8t6fBDG0fSrO3L1RzEeWNwWT
zNeyn4oL2yTRazGMfqy1WDoDBa6YLej8ESEHbR51E6DIPXGasNWNELNl+VBcKCkm
0dhlt1qn3evMq5cmYkUX3Nmak9qg79cXjWY5ULJv3lHEn0XYpV2DSQsETPnbtK/4
rQAy8ApcfdkvE8v2s1kr1r3AFzEwEpxN/HE8oDtsQnoW06vB/CAgXvYuzZvDh4r7
53S/JcBVChC7dYI8N+uNfCnkyLOT+qAmoVM3AbEiBbwGb+m50d2F5icCMOphqMlt
BXU3Ot2vJsf1It3G0XbHVSLRyQgadtP2aJ42YEsFKg6hqsM1W2Ju57ZbYSUpfJ6N
G+G+X2kW18qFqm/zUkRP3mKYL1XUAVkdL/omlCEv4zIIxXxRhJJcQmk6LeZNq5EE
elNnmtkn1x+HjfB3QVXYTA7cITyddokRi/SYXi4VyuSJ4HTE32VBGOF5Mlbgvs4g
IX4tFeuJ4s4pKEiwtZtazvlQREuM6kFaZbghfXMzg1dmtGn96zs3Csnd4HwVwh7u
Y95pf7ma+Uyn1uD4t5FGwld3MkYK+MuDm7aCn6XodL604LOBcvtlrrI9jF8p3AC1
sCTSV9KkEUgTZFc3qaA1H+IibICLKvAPmZfIpAtTqOviJp8W/W9xMXokrlmG5Jc6
wOJpI0jV19Id70SxDWu99LoMKnoEOlrxZLhPEalcJxH4MRSIT3WZTk3d7CF3cXrQ
2cAIh15mCynrxHeaMXokDDATVDtr91C9sjv0QAmgybAMsb3cq2U/dnA/PbD2BvcI
JdYquU6JlDwMU6hRe4VYYAIZUMV07sNEGRNTuDUiFKoMSYoson3LN6n1O6eeJswb
zS7yREFV7rxjJ8ZTNY8NmEQdyYf2L4NIHFj7zj5Zk5sWcOvavlRh7UEbcZo/nUh/
bsLGiKcv9I09uFns9mngGlKTK484O2Wp3aF7KcSoW2mCOPBu/nMZacpoefFFsXWn
r075DLf6EfAMU2IDNIsismcvibmmanMy7vgpbginGoYtZCnEXFrBTnAy2W7NV4tZ
YxuQMX6BOcMrkHbmy641RYI6VM9waqOy1zGIESQrKNDEJoSUzxkDBGsL7zEJ5r8u
o+ht5oRxncGLN6ZMA4m4A/PJ5XqRb8MvFa8MjJQjaE11XURZeziANI0isNhAvf+4
HyLhLOgjvqm9/TeXWoFWUzyf8Bk90gW8M8wE8ZM+FLt9cScZcI+Lp+nfVDFH1gHw
hYDW8XIHh3DsqTeVCwsmPNei5CysRzEDx63DD3MrBnt03RS+UMNQ9oBGkFjJqmmb
Vecab4y8tlcqf82b7ue905n6Zdysgh/nS87xtAxxzPtcsbi9rgsa2F/iLshXB0/H
mTRySNAQ+wQIeOlzfeZgZRKKkVixeCttxPk8l0IVbyQ/OApi3ayh/M+erdbUyzqG
srfLkmG0ot5UabuG+TZKggYmIYi64YKZJ51t6fJnIchh0nuNW5qP4O3q2abioaZv
f232Lc2x4aCRkQKxyT2+W4n+s/gljnvUSayKq28uzC+TviBYm1SsATBlWxpFlcL2
8C+1VRRLOY7HMJGVvg5SdysYRpfrrQZpTulj/A3gb1pWKtraJLgKMUKH2CUQkap8
Ai191QquWDyEIwbWgWu5tGKFyXb1+8Tsq9qOWM3WWLsbZ/yQKxbx01dBzd5yCcZa
kwxxFVFpyPLd7jDjqgTTq6olb/9OpGO2593xwVE3j3El3lUlU5uEU4sUhuRyivVz
EkEtX5gP2R0BF5sIIINIBG4x5Bo7Yf2RK63ZJjrXE0LXFa7hkwsntKEO8BF9Y0Ga
JdJqtgY/JtBJLRXVUfVPD4Mv76g7BKS4cEDvYlrDuy6Z/l5cB+wXS7QsDXRd58pv
KARzcbFzIOIwuEJZ3zUscYAANxCvAySzJX9tH3pCcJ3ZIdR8yKiuTKOKRZJkE3DQ
U0ZDKmb8IG1qVJyMwOU3RMuwYW5MkWU+sS8W9rcY9XSMyUGnyJNeSZeRcsfPSWmK
9HK9vjnPHMz1fvrRFMjjES3mxGVrMZN0+ekW1v5O2B91szXv6ZgMXFqfuJy5yqmj
IH8+Wl3HlA/cYGZ5xbGUqoS2ODI13m6Le6QaP2ZBuP2+qbnekc/UoPVIFPvzmxxB
Svm0j8BGXyCXE0QV+Y1EtPnFiwXareaXDBWKBiEdnYeg4owiKjspn7YGNxDTRG2l
097t7B8Vk148LYo4eT4BUhQ+jerm2DbUWRsrU0ymIZWcuKKod3AdLP3MTUkerigR
s/DBUm4Lr1pcu7qHCl3/2Xu0FN0HpVZkw9lGz7oS/QBHv5t8zPqoQo3ozUfwIah2
OJyB9r2VTWGCjwp2I2NwoW/ni+OcNpeC7dWhAg2+maaEM9mo7fNND94YvnmM1F7e
3Exe8/Igy4J3aWqGsn+jSwn9YI5oSgOjHfrA2+m/yba+qVgKMBSbegHqp7qtAv4w
TsKWRF301kpeUMQy1CJttE8lWVyixlsAWVwc0tTfZu8vw5nu3TylcxqMlc4ksEIJ
FQgeA0xJq0QLsbUfP+SHmIYDxtoSt4V28xyfc80wIRTloDW3LPiaUJ3EcHNG+KwO
EMYQZAZad8hnPTtYVn3sZoYn0J+irHBtZ0Dmvh7yMOvzl76vNoookS7sfk/mwLju
DCXg9eVuRf/SDJ3uXE5sPgtzQaDbD6Mo2/lBe0vqlbfYJ6j43f9QXiVzcC0Esya3
IBpHsjTZX5WOD/ciyNE4zGdqJOkkNb/MsyQQPReIrftdK9x+I1M+rz7rFZJsP4aS
w3dbCXViZmNMQsbyDaYVFC0iC/oXLlb4ozr+qKOAvrSieiahG5tvu/QxrOcDEWHg
+lcDPF4ogA2ljjApGM6rk2xOeHczXnAQqCsigrphMEof/U4kKozW71kb7j/uqWof
s/WQ0FYPuq15rk6MM6AJ76h1thINjtFXGtQeSHYgzP4LV7huwewBGCqTu97tGyXx
9a1M86V8VbFNYljPS5MmpynPiqgThwsCSP0Mg99rKage6ecZky/ib8Ft6hFYtwPH
yAfeLmjA5bNyxpA2mJJtsAsD1+riy2WBShWcxHC0DWnh88lv9TjjQqv4RmyqgenS
6n492OwuWxw5cUsgM5wgbgo4HvhAPS8XbsGDAYjb/0V43pkJaLlbzhQCleG/29sy
Z3wrY2GwZngy2HU19oaQYVUZTGOZqTs5AHkF5WMxUSbk5rewbf1SM5GhmJL7GzEB
pdPWd5M06mR7CT6MGcQ6ZDeYNkw0LaRQ/hYSxw7VERUfdZGq+IFj8Jw4Zx0+wfRI
/PLFUXQ7XorhsRzb+Eq8sZ5UwKnZ49XztYO8zTo2/YXfRO+jW4Gt2rbTpaxTMEUM
fbpe2yEBlsIf52LUzpSTLzIcXxUAUAcP2KIReYCDeQcJzVGtk+Bq1kTFF0PDB67O
L9qy+ncdHrJPbzl+Qu2x09XFVWW+J4+SxxqPMMc/f856STKHkbEuHRDDy2vKKAPC
w2GDrx8xmsw2HxQcu40sGLLr26tE41K/7KWIYflGXjtcLbsBdM+mWD5kb+Q+s6W9
YcYQgShsig6H/PDPG41QVt8T087/20ELK8AFCnKPLKYR7UiQwZcZ4HdPObC23N4k
2tObikU4bJKME5LkT/1FpFqDCufbZPSc9s/DG13pT4gI8AKxkaNIb4c8ps1qsOX6
pUsFimzLtD0VL+tB4f2xLyPyN/Ifi3Z52NVgbVNTn6St+/osGRxWK2l37Ov1rloN
p5PhEm9qrXdPFAi3qVtNBRrtBC6siqQEgD6v1ZZIhfeSxwXeYeH9JKZAAQL62Cpv
H3a7fruVAe9q2jDiEaJo59lRga1Fwequbd3hZPZRQai8xpFrAQzaYuYyy455d3uq
PQUag3NW3oiv6CUTV0ZEwLTBdy7QofZtDDMCMH+GwQ75Ihd6mvNPxhaujJu4wMAh
/Any6AL0dbywbhtbdbVI5mseV6kBgcb4vtRrSAUd4BT3+n5fK2e9KH1m38ltGkzh
AFcAvO5FcBuONcKhIqv1ypt9+fHbtJVZ2+ayt878+6XAxJZuV5H1ng8D4MDbvnHl
rm1RqYHsGCYTUf/9i97T7IHZ4wKobidvUqW+VesuvFEEX+0pxK7Hkh0hHM2pcX0t
WtdxrQjhda8dZFq1h1VTbxrCCx+myjXKUkjHWz0gHEQsAQrGojRFjLqyazWNj4OY
adKYsMX7fAlXEXJP9/kp+oDHwBzlDu53I/Y2i1sJJwPRODASBxx/DV1BDmz02wD9
/zGa3kX5DY1qthWILwGFJHra/hWkN5x1B3wCRW7atRhcfsblSZRLQ7lmaZ3HEmwo
voA5Nvf+BVM4yX+5/K24/rHMdrm8eO4XaLeLlPmO7ROOIiC79d5Bg5uaDtwLa8Rn
FR2i5qr98IKaD0BlTfyTVz/srhfXoM6EWQlgJBeZiH03jAtF+GuEWpWvCvC/TCI5
nX63D+S9kT53SxtQrsrP1Hj5yn6qnFsmj3xWyWk8k03vZFTss1So2p1T/7JkDcpI
9rjgKOJVo971x3NyQRPq6lwpWas+SqXA6DkawgRp3HmupIevArxGhsSl1DgMnPhD
NXvS+81yFYqqZ3z6ckV/NDSWyJTfth2PEj/dRNTD6s3hySewrGHhwZ3KpoKBGTRw
5bwtnZJ5Ipmf7zTbuOot4nobmk9p6U4l79PPzNJtejjABrFTxLjM94TnW5MwECUZ
smBPSNcZM1R5+q57vq6hwYPQdJXJvTric2R5BvH4F2HDwIp/y+nkPLnq8rfmTbsi
ac7Q89d//hqppZ6iQ5J/nEtA0eV1rFGgpZFCpwr+piynZBS2n7VumGXJ6MJNJLS2
kbY1KyUBe9+4rXcqLen7Iu/G81kDRXH8xnGq3OhCGqEyeyrRxJT4T7DCn13W1T/I
o6owdD3v38UNop08V4F3nFhc/An+B1qjV9tWIeVlzbvuY0WwVgfHiKr9/JaOp4U6
bFbidFxr3Z4IpSTNKgIP9PI9+Iy58lyThzFAwmNt3dI0yOkXew7Wx5sEHxTacEAt
a1/5Dhhfqs7DH3Sg2p80ohiuFCeXAQ34ooeKq2EoGJsRJcQ6f+LBIB3fBUE/NHu0
olB+HECGH/8Gbl5IGDqqYfbu1yiqsU1dbDiaf4s5vFBAZtJ71i/XtxkTuLiTCYDV
zmjjIOBmfxb1YByjz52paiHCAhaFgDhZNlzPupcv6L+BuU6Inx94I/3ezveBMxL5
haVvcfqVm4R8jOED2bfoXZxPhgpjK5f/vZ5fmdLAZR+K0eOrBxMnhmmiBBD6PgOH
xFLMHD1rUrsf+QmfaRJ4HNKwdaFe/F0mJFHOXdDfFbhZQf960UDQV1ZhzEZbCCYg
15ii78YWqVfu3DS6pkkd2Md+/pL+QXSSDcueVqCOf0RexrGu1NGAXRE1utQs5GXR
CfkpTvrZc/MiE/hzOrS1iIov6OIPJ0h+3EZ7UVw5T3qLxfs8aPrN0C07U4v0Ir9U
Z66zHHgwjEt3omEKnsiceFFP7GfivyITOmIZcSiQHDSr2zJLK+mKHBOyWGmB4Maw
IJQN9igghHRZ4Cyzn630Ve6EqlfIF61k238YbI0QOnSnHBsGJFi6Gn+w/gih2RRX
ISHBM91/f6iC2Y3xjrh3LUpbb6+ZtONcZrdIFy4GpZIpld8eD7CAYy+Xs3TOk+FW
FCVOGZcde28qa6jGeK0K9+rn/Ukvss09aJVO7Cl0NTXea4rvJascmVFOiDszND9f
4Cfqsrts4fbJb5YWfaYSbAbvzYzXrGBqXBP3OAWxwd7H15ESgq29na5ewHCv0ioY
1J4VjfIBORz1rTmj43NH+vR62+gtpsZg37OB9VWz1JZ8YMEW5opKDeVfZi3Fk4v/
+2DaFJmL0w18ta9cQpPXjV387jPikLRm2f6c9bd0WMEsT6q1usSaKLrwrjkpfzy3
s+RIAWHixb4NTZY3wTJnAlSPEeznZ6hn53Do9pg84BVzoZDWmyHdXd08QLfeKi3g
spB5TBRxP0cEJ/A9H5qHB87wO1WnSZk9GtKh5RVPaStPP/SDf1lt+j5vvN5G1hh6
9wNSLWI7pC1Q1+j2lJw+uvQzmOEvfGHammGOjt60zDDeUiQke4K0ODXgY1aH8082
x6TK7mkFzCZD2sqPNS+3eWvGA8ZIFQV+EukYcEBGqaWpePlOsGu4SbwE89SQQTrF
JyUJhZreZuscGXRIyXuhVHBX0X08aczIYkWh+OGSMO2kmE3FOnt5UAhUtaxyl7WF
uaOvFcVn7YKW67gsy4xwRKPDeLQDwoVcF1nZHz5rWNl0+CDgaOw0Uht9/Qkb06eX
rZR4yuBH3mlTpiGgNnMUAETJ2F868IQCqH72kceZowETIXmyK3TEMJiYeJxH0rVW
oV5g/6056xs2iun8MKK/+nU6/rXKQ6Mq3ruDF9dg2igSD5qkWnxk2hYByBSDch/W
yCPBKFIMPtrWWZYDUNRu7PPHuOjfDBk+XWxwPB+GICVb9/2tEzDyPZtJPlj1HwJi
HBye/E4iSH0YEwXhtpJKd0icTm4agno9Cp7qDJPZD5BrsNzVwTiEVtTYwO8EspJN
CwBxeUt70qAJgE2VqORcIou6SwjnZoDllhaeoV+jDyzgz6BHgYktiUy58xkLt8lq
jktT5igboBIbLIiVE3+6BBYIxX/P928izcqr++TOmwUwW/2Kr48s3/ojc+4x7aJe
kM2K8EgDuxZO+kGZ/sfCCHtRZikPJ5L46911Q/l212WyZJVi3xJLS91YssTponNX
w07PXhBTNA4FiIDSUCvbxcfMpEE+lYjidkoYLFlo56mGy2J9aAvG7p/24N1FjUd6
Gh+CfIE1XQDOOzI6BdKD+d9LTnn22ed/sKxaqCCYuSa3UTGmEdCJpYOqTV3ywrKb
jopXvDqDRadkYqTbKDUjP08oemBhNQWzLdV02oqD1E73Q6SQ9R4VDByPkWLs5SBM
OQkCusE8y3J4LmI2dKelAnfUNE2EXqPywcik/cBC7TuYTJWfoZJRJWSLoxSZZ+TN
sfltRDpPFj8q0tbOamKaEFt29ORIYQFnQGueIvhG9tcfuubfLVhrZqF2bXhGx8/R
yavg3OxEv8bXhs+WJBJpmEoEe/yAYRHN042pNvtOOVRgCH+utx/G3yidsixllQ9A
THre9+yf10BzgK7flcmNTaf8R1rQ894KqIuzdc7umE22TLDjpv0aVwwoI7BL1r66
oawm7ZBZESFEPE1/gYy20tO4mCp867wDaiSNuJANwGORGv+s41TB/HhFRreeAyTq
0Zuf5Y+r0CJt4+0eDKRFSEClI2AukEmXEOC3pBPNgJ8/dxRnyKKBLfdaptaMB10v
LKnSbkgYQuwTWh7eEP2hOvnYs4UzFvLKrfmy/XnSloWaqRY3Ee1QXeILmx/rRX2s
e5d1VqLvdHDsBYkOOFSrlUYoCh/6xt3mkiz58HG4Kb/+Om05jmiA9IgN04rBykhA
pUL17cm5EC7SU4bIR3anfZqA5t85hjbzvNePEdbP/KYlVDIU8CMi6oMweqZSmd1I
O3NUvUqCEKkWQcOZR2XRhg/V0pdmLhQdJ1V9RIEL45sHray6MHN9nTdUZ18uT6Rn
Mu8rm+9HZntSO9vARw7ge3JqKsgZyQB9uVkqi3DLcn3ADDdmJvbHGtC/OZdQl1Xq
UF+r49oiopJoll1eQEmva5/w+ntQhNmsvs0oVQfoOYGKqncwW9XJnF0FDfSMIEhq
CxTN+Qm1UKsxPau6UlemuNHsy0Jxtrklp/FqJajciYqlSIKIBhcKpvaB8MtvwwOR
LTu5d/M0Bwju56DUcS+4joSuTETSbhu6iMMxYO1rN028SqNplKBI33AmC6Rio1W/
3vZMVj8QqZHkPXmc1o67AxG6h24Gaec6lV10GE6RLjR3C18HxCxTFrmbfNUuvYGM
JsAEO1Er6hjkDyumYh/n3yXn2sTkZTP6qXmzSzydz1lNSsY0g5XlMzS54PE4X0EH
dsnIYr3DIp0o1HZyNlNRyvOwPMnBrzM5TxQCe7+aqx+uSuhiYaSnOkoot6T2D6lV
ORBHu2XWhg0zSbrDgKA9YY/T3HfcsDAqyqbq9lyDz+APlnnhxW0l0D9kB+HhEtkx
Hi/WbfHZMZaLC/aqoFvtvFB59aRqrZQ7sghu+cFMMY3yI9ZYsM3cpIi4Jde0cTYY
rf8KhxLu+RFysqN9NtGz3x1JeGUF86OUo/cD0uHl/UQ3tHw3cqKma7F0k9S+PSan
uu0jJiBBHkC9mJ9DKjUXsHZaeXHam2BigW1S+vkJpvZ22zUP634L9Q9hVEe35d9P
PEzAgC8adflOfu/T6WDMyHwbCvr4eTQ2ihD993k4OjOXeglUqebY6hh56j5m9s+p
KWg6q0Jvyy6sOVRFvWPAGggitMq6BMkMrhXbTTD/TLUokb8boFtmgyPu7YgceNS4
KlYMW8kqAkgfzfqZjAgzDu6Qn66nBHoFsKgdJX/jTs+kajp9AJH5HRxe+t1g5f8H
fRrIYC1u9moD+slnty+RsqR2CDu7ySvQVV6quVUSip+AVCRehH5+uU+Tw/kAhIw6
95YXJ5rJY7fXX1M3dgMWGLnxaOnPq9JDY59a374p45nBmkXdJ4IQtg57NcMICSQx
6s7+cbpoXYC/Ni78qV8rAvBoyOVZB0Aq4rJ46m1t1QQWzuk8otDGcLHsk5xxODVM
cGgq5XVhjKkKw89EEOZ9cv+GUBH7ITYOEXHwuqXfTm8OdymXN1huz/FI0E6fN1/n
gbQFsv2kTz73EMYdYt2G+RyHZ1RH55bCwpqiBD7INY8qnGtzrMRfazsHq70CqRLr
NtoocuJrj4Hxd2XAoVRwdZeeC63EEUmjdh1n6Ji00ytr7YRysAQ8rBlxZVgTtanK
/A5iHmv9BIOoLnK6mIsxFK3rMfBA/8QBYeOQu7jPtfb0oVMaE2O1KTj77+B9AitV
+QGvknxh4AR9vP/Mjt0DFgUkMN8GCdZlr8hj2tJGnWlirWQrdJVVBcL2CU07trT6
oHH5+ow42ODcwVT/EtU6mmqc7Q56CSJ7johfTFf9C8SFUyyXiYA+zrLqvjs19d3Y
rqwX58qBVwfLKx4zUE+yaGGqVXppTCPFvuKDFFtigpxzHwp6jO8+N8uSXp74q0FS
+hLCMaCx76fcQxCPrD7Z2w/dnBy8NjzV6sS36pNYSOMONa1WSc8TASkHscwUVb+R
K84Zf8zVEYaExW7A3YogG6buROI1Mh80v3Dif0892bmc36do31/fOZnC/s+60znn
Er1TQi7htE1KOECBOWdIlqDp1IMlG97edq5Nr1RqTUhw0QgeXdkLaLGWwsG2hbOF
VymQKYQxYtjD+GNCWpG4qzUpUyfdOQB85tX+IZBKSdjVMvAo/4pssRNWwbbMkyEM
3cZIKhSfcudtgMZcXujXrqI2iF0ak/QL23pCzWq0c37EA5zXM6Bp9qAkLFMEsQJV
4E1iZbYhHuiUCbhERxCvOfzs7/2xuTDM0L2DtszQVAX4cfVEbs54Gj0wmW9WpU+R
P7bGQtVJ4WNtYO8Xc/U85QZ0uRueZPLagSH/S2LkqlVPGI2DYCwyKiO1b39RhC1/
tzJdMZvFzmANo2EOy83ZTl8Xxv6fBt8CbfzwoaUCo7iDuhE1EsefcvC3YBPzM3pP
i/XRFglkNiAMHi5na/RB9DJE6mRKXp31xStcyqjR57FKpOegRpIcU+NmbJpCpdLN
0xMEW3GfdgA5H5F2RrI3bMVc6iMiGL3bZznhHJFbBWkMi/98aUHXAzlpV7BgGkZl
LHYxvui3u/+hX21+XTz6B2iU55UM0lbE+22lBjxMtiAE4ncZ2Rxoubu5hblWQpof
+FzJeeL77383UWyPTSLse1ImBXAt85DsPzl9xBHXbgRYViwc50mRELRUr4UYzdBN
yb6wkiejurZEN51oDqXgmpl3FW5oS3b7tOTlXzsC8whO/lrM+naE6enn8qPOZA8Q
QdR/gakx3R2cyl82r8UjuCubjOlSPRJ5D0sY401Wob7mJl1ZCGx49EwQjpaiXeFx
dINJ5SZ7gsHF4luHvRWEZ2nFg8gPvkbs4Kk8n0xIDAxmF6gnqSLaNgGjSmD3jv41
6wiFKQ4klduwlP+Kdjf9ABeOIQLBpPNaRjF6LRsoUwwBixqzUDLcI1SwipgQWtW/
+btgY+0UXLRzuzJycU1Q2Z+SpQxYr6tH9dpVs4XCJo7PTMgo5AeN8qM9vqlfO/BK
rsiFBSNbuNITjZOLF9HBJUu0mgz0olR++GU56Bg6VZdRQSBqnUoGpzh3YtPTku/5
6kHSKtaSfAC9fW0bO+k6suatubmn35w4O8iGmpWSKrnQMc1t/NzqzuC6OBWUBMTV
lHAM61WAn/+tpBQQMyDZGZDZ38oJTdCTeDGyfchDbTgu3mAtQt1wmlKInoB6yPm6
GJ3gg9zr5N/7fcnnDfIt+cEkapkTl6Pobi8Cr0bo9WIVC7f73Zzn6H/t1hmjWxu2
A/ykP+iNi6Wi9OPmeQxLqrCG+quGRqRE9pt0Vvu7e7l1Aag6DCClCnnTXxKZxRRe
xUPEhnIdy1xN8UYZ3BPBATB8AoR8xgWcwL+ujr7yoZ+t/BorHsHe9PVPzlAIXnjP
EzkXr03bMyQRyxAHlvYSgoX6oBF71qY679/C2/m8CvEAlDxk7rBae1HZLS3xhLAh
hpyWY/j4hAH8/flDfXSS9eAT89JDcqKdcLHNy4YFlEQsCTpcFcl1j0NUDZCMrOfX
7uGVFzG5LykLw073IMl5WMq1lbybpAUBI/EAYQ+Zj+4ktsaQEceCpm/7Qirr3uKX
0Y0nxpjfQDg+1p3O+S7DA1G7r2UKcqNis7dwI+rQHXLXhoRK3krcCeUH8HujCGS/
S5ugfaLN2mow4+HObRIfb1K2IPataZC/3LIegaRkKnYUAjl6DYHv9rk8jQoXDdHt
AMR7eBENRFGnNnu8MjLNrMXGcCl8iHMmZXklMH9XbjyczQTA8aJMHdQj+iioQIgB
Wrc2Yq6Rq3NAnkGA0azWfB0v9s9zS2DytW5IYybeTyOyV9yKjsxNI78Rp9PgO0y9
YUSwC2c35LJFAFL/o5qy0Rj4dIlWMvZMUNrvpw0RgFhWvVimHKmvB3ZsuNCTX7zz
I0mUeivch/IOIq7G2ALiwN1+ZVtUAYDZjtqRke856nUAr1SXPB5sUPBw6xsHIHjZ
efZJC3eXxw6tMIV3d1N14uBVAGDV65deUeONfjk04x0RoifJSvdAJkOMV5CpNt6l
OAeVTknx4rl5AUXEpHqxJPF+8ykeUnWt3sey0ThcT55ORqISASgMQvRLHrrBa50b
hMVhvWsuioHEiIoYajkwU6QVQK1x2Tm9ZQmITDFaWP/TjKZaG3Uoe7VVUPwc/05h
YKz3oZ0Xx0O0HkrJf0HEZFKY3iCP6i+anSM7vhUrW35XfuELJGJLVzW7ldj7HZv3
HL9uDCZpCznNZ+S3BvDK09fnvXHk3uuC0o8K+p8aL/sWVQHuHapMPjcRnB5FQuky
eA7BLkbTOY7BPie6+Rz1iZUAlN6LGSogxAY1AwqSGRNF+kBfZEgc6GHq4IXoBynQ
o5kU5paxoOwNlZ5FZnzvIadlUxc9/n940M5dKw829hOfem6bQ2HhwfeIZfymyM1e
ZeEXQPVkh1bo2D2t2T+AFHh3+FFO+c82pdTeZmO7ykMPWlajdlt7Gmjemcc3YmHx
7mlWsc5Ra4ZXHmbnEnIBGEhSRVo+eSbpsVOvYSgL1BI9HlHjPthLIHk3YW0cpTzY
yhF04jS8euolHfv4Kz6gBAk+5T9HJVOwnfbnt+Xzq+f1ZuOZg1lXNd6XoQtyZMnl
KYeAlJ3Zty4hGefMiJA+r2/WVm3hm23MYiLeYCdUsOVgsKbFLfgyC9+CcEslIPpV
MgkWy60wcyMZ9HOXL6EQnxea4RIXY1SPQF+zv7z9+JFGHWO/3r6ZWK+2PXWSN2G7
5raAepKUgW0Epbr+bgRcAGRhuewzXgyGOetoPvS/3fNjx4QnK3BYKw32WUkVjbnK
mAybUJSECWRmx+NE2/NqXRghlsOFKwI49kBVK0onRdXYU2DfWAxFr6x58MQQHx0N
q5K7u06x8OBHS4+D2vu/Sjmk3RgvGChNYU4iCHdkbSA5ZSFZMeAYVCfOlpVB3G9P
9Lo2k2AU9Xsoe82iPTN04/y66O74SX6otRcyyUN4fAU/WHEHeiCpKgE15TQlEIE+
a7/oczIZLfbCDiyVpQ6zDx8MpxiPVQa2E0BLno1elyl/YEIY22/m83fHBplmiINV
MEtBHSbBUZzUZGRewFxLHa9ifLNFSSKd1lOaynzw1qUefKNGQ97kEyRGuT7qjH+/
fhyhklObDwbXhjmr6LQeo1eLuP63YnCLyT0fasUTII4bqO94hqeYqlsI/kDZSxCh
Mb+ykyD4208rAK6lOC51HsRe2rEtK+fVmOLqhjxH3DInoRCocrv8X0xvvRW8nscO
NvuCxqu/2CbU37ytQsxu2krw6ZjSQSRQwX7cccYGsGpXDssiaOhAxiBVRPnqhcqm
9+hB5I6dmidVojCK3sr5beJwcJ6Hh2phXkfEatw/JXZOn+Vv6DwGjRmlPj+hPUhj
A5zXCAoFDf2mLNGvQDbs0hjSPXuLszwFU+BAS7dCnzBJh4yDH4G9JnL2KcxJyVeH
WIBRcPeGIb/QXzN3JrAijnar58ep1XQ68phnespwTMeZv/5Kt+3fqC9yt3fu51X0
4vQtpzVeVvZV4+Ie/KgISlwHNWqpek7Kqo1euhNDgZYULIu80bM37/N5iORIIjfi
zV4a8vzXWI2VFz3WP0FX4QY8PYsYCr5zDgESCGK1qP6XtRpXYxtqr703KBG3OIHO
6oDr/GwZ+vXtuA9PSbGPhUeYHXGV0PR7w+sEO3w/9wFRllkaz/9X6R1/vQNtHBDu
5i89ATdMBhLcnpg2sF4G0v8zY77bijRQsmkzE57/feEBoWI1mF/yepRs1wItrnZs
gnWWC7dtDXw4TqD5ShpnXU7CbDFVA15xUNrWs8GHUA135EYB/76rKw6z4p1OqG1+
wbx1Qr2wlSxrB+0QHY4XJDiF2fOsjCRRaqa0CnCHjm5e+iUel4C7Ld2pnKeWof87
whs7cKBoDReydPudr7Q4Ti0VwB/jhyDWYaqJMcGtCLsBVADXS6cVguB6LXDnKP2o
seQmToF7jzmtN+ag+aQis5+pXVL9YOG/QgTWlpbqo97/Nat8g5mzc5mXh9IB4WJq
8hwHsUqZ3MIeChO1udZUN1KelP1z/H3HZzz7Xln1VmOzc1yPCCe7e2x1pK9pikn/
q4LZVBuvCU9BnxlYXmKLd67ehB7Ipuey7tmBvSwEiH0mkeop3ikqGmKpNgnfOZYL
PQWmQY9U5YDjrsU1CfDi/ujuc18jyPh+cR5eXfiZETL6Uv5YGE2ynD7bJ80UErgX
z6PAl2oC6WkLhMkGu/WwODzKcwAeX049Rf2qgOrYNjqdzAZWKb0t+1Hb/XsNjf1k
xrn5cO0sgwscy+3Rq794xlMnxLitmZWVSfEZW63sogx2ijf44hR5xb8OLR2lA1kQ
Cvu/aoGFHjvR5QiRR0D17NY9Zg2VowcMt/YIWlMODoE3k0QSvs3bhsELpSYJ9tFL
Vgcly/qfKEuIXPTqd2R9IiTCxXkHkKxOQ5TqSl7Q3Vfl3pmbqgOH+APf0fpbfATh
ObuBlujregTW3SLc3rFTvSR8YLa+06mqYhNzgSQE7nxFIMqIPVO84peWMWI9d+Rr
g5MGALt5qoKJ/1i3fwzCU+3cNXql9rfoEd6AbQvtkWI3MLvGIdiWor4HYAQdfOXn
/Vbp1lP6+UCDHlHO/gf8TQEOES12uVGixclFfQigAe5rEgCT/WRxeB5ryLjBQFlP
uqbdPPBpq6k3+m1TRP25LMXye3/ucFbMzU3QPSvY8VrdCMb9PqDj0VXYUYPIj/d+
wPZZHFbNxnnEJVE4hHLf4zSOVXleeJfX3u5rUBURxch3NK2G4Hp0HO24eoYhbKg5
reYpw6s1BtIzs0gpLCGLRCl2T9+bl6C1budWPZlOyt6zn8egy62eYipQ+vfGKtjI
ur+M76yS5pYTD9V9Z2AQTgn3Q1Z6d0JMhwZNY2KuXPiDsL5pAQSI5jlPxvOzuEys
ePofQNIfBAKOig5qAhUAoo4t646KAJbygAcAH3qrrJH8pgDqEAJAIHF6Di90sszO
y5gF/P324oDtmZnBNAV0MA2Gb0nazuqEU5pE1ukFPpP/cWZZkiA74I37MTQAU0nW
Vn1CAOSAmtpynusyCkwqqFSr0k+3/CZVUe8GifJln3jal/DlauiAoFkm70P4597K
jsRx3paB9xJeE7Zbj1IQdmAa/hptsWhAR6sfFT/5xoc/1aikx5G86Zv5sykUgQTr
VBp3ZdnpRjAPl6RtFamDldLpoYmFQF58QfRw7gNd4b+5+jkJ7nbpSQlkdnc+K6hN
c4t6PYQNL2tXqbWbsS9unmt7qoV8qBFdOak3bm8VZZSdJGBAPu/RdrxV6eowF1Ao
CWl1Hgpbmm6kF4LO2gv9f6T6Y78E1E+Z5D6OYdN/YpWt6m52TN6MrOFrYwgwugha
s42KU+cWGjt220dgc+lKu3BkUowh1uwU19b0R3/y+KmtFykMjln2XoHF/GaNWPFg
cgEFW3CqbspzjFb7Y9NUmttma5RnuKP1msllugm9JLkxJjAHG3Ux8+YjLjbl+dl9
8HfzscYwchAehgW06u7mPNyq2NXv/wK7iKBJ+a0BWmz7vjGig2ahxbP99jCU6f6l
an8Mn+jBvLGJtCyx6h6IqPyKL/Vf8AtdB4S9jUJa+8CLoFNGOXXsdBEtjdVp4JiA
+lH/FQdT5Gc967meIMoRREDDOBJIHgTwY04PlrDsYCPW/F09dWHiAFlmOkovJiOw
JpIy9KZ/fH/+34VpLMyTmB6wsPPa5oTSDtqCuHcMs69YVsh5NUFlYiBRI9KUuPzO
7Ol+wFLc5L9eLr3WXk55IQw6dygMUu0ZzCcAwNC0ttocL6iuk3jvhZ0oSNI1Oycv
IAmbjD9mSqV9YK7rXnZn8YV3P5HjlU4SPD4i6yk8QU33NY6l7Ld0HGOJaiDOLWE9
TmtPekVmyMyTMeR3iiD4n1lOm7YT9JgLF5RjjekivxJhVEiXhZkB+Bj35Mn/0cjy
ECXpdBhMMbTJRVv1NnykZ80ZLMbPrkiST2kpHbHxmcVADL6IzNsTiOUQQUigLLaz
GkGqYeGwkuXbSAyQSamjcM+cOhrCEqrzAUNO7L3uUZdhJvXrNX+4vwh4fQBcF7BK
yJJtPfB5zS1fd6vwnGSSr/dXe/maeofiuo5mzi1Ez9Tw2uMUcrI7V7XR/nRgY3zQ
jJwYBJuRP7pHubOwIXMeNC8JNMPDRNfNg5emyDhQ69Sht6MCCh3kfYSntScUviGJ
QF1LTbfw2DndSbj87eJ7XQ/+fLRspGTtViTh+Ir7W9zDGZIKATl+09UA80rGm3l8
2ArCFfF2ZpoFnXblYkvEgkkyRnBE6L/2INJlSIsy4NvI99V0T3aSivP5+PjPmAYh
yvWwcUsIusUo6DrdilHW1C1OvmHsPirXA9u72CmtLvVS1eFrWN61qOAMTuorNv8B
s9I5kIF2gAENupP4YMZi2geAGaYK/6tPc9tlZcG0Qj+oQuVGSfsBWuiLXzu2ZpNl
oYLpjHBnDYgcEhtvzZ0h7Q9eOFfm49ak6Jz9dGER0sQIhcnkZS8gqki+cEmK0hmP
5xmUJCVceuPgQV+2i6xZFcm4iOfwrhoiloao0Xqh8NqmPZ9Ysmzi+Buibh3Daz6A
G6LS2fzuyDgkXp91ifv8jLYab6rBimxeLQOsM8/xlKBdm2RcmQNbtgiTyv0Q26fZ
jhu/jDR+h4slK3LFYKO5SGGPxNwRugPbRA+lpGShyQQoFTz6MSQfZb37tO04nOEU
hR3yp5wNeOad4ARhLY86jJEjdaSZh5f3fmzIlPthseKVJE1nnQY4RoSkdjGDXmfH
N7TtfUhgB0m13qOZoxE8DMDhBiasJ30zlb7M376PSov+z5Meo5MxiXff0uv8dYAQ
KuJ/Or/UcNP9YZlw6hdfofFLVrKDESQOcAnNjs6vgq9MeoKv+ywFvoVNOOwXc9en
uzVraYi5KgsN53AO0pM05wEWRnpBwMzk/7BVzg9WrzkeO2WSTKqh9tEDDzAHfTJP
RXzruKR2/UB8pnQyjHABfG4NghRpPWjUnzfmG6ogeVxwdFrJUs+oQwDmZ1jZG4Fv
hqc6mbOjYIwY2w0rDY3cF5Az062qCt9d3vevmkqZ+4PVDfunqC9qeCRMiEcmGMrE
d/Oh7/QjYupjZXT4fIBLEMvnj3NsqpYOfA+tXxv3TPlaPWrZGaK9F6/tI3U3RDug
bjq7kuDPBoZBh8W1lkeEs0+t41ZU9T04w9btS3VKVWbqfeQ8NNSq6DlT02HoqWjS
vLikBmU78owB0/npXyGAt823CjZhdjAdK1tKYyHqwW4C7ioEomvSP/0/eg+i+4c9
eVtFEAzzVZcd1j3r59TgVVBKFKJfX9diHqw6dhTpLOx4IBbBnXkG7ePG53kE4bo/
gSVAf7Hl+mJtzPp8b3MaZG+0T33C2DuNpg1lvWl1QTkdSTGeQ1fUWpeoisCq/TSB
rlAvStiBNWHzlMv03vfCo/GFAmB7tFzJFmX70CVtCvjjuii4LgM04cP61Yfoz28e
Hj+6Wp1E3+wwDhDDp4r/SDshhGqlv1PsuoioTHXwy8ABR7g3APgBG981zIQ9NiyN
khDXZAiiFsiF0xomIk2qzeG8Ppo5+a2CGIYbBc3TKovym2oIh8ymKwPAyM60oT95
Y7q56TdQgyAduxMFXqY4QRJAWmOJf8sb4F40CyeNBU6oUrCCI4hGTPmqlrgL3YpK
R7dZeOvHrNaYtw87DieRO5ydl0RSX0XDS601qO7TOVBNCbpMVQ9Zc47F3vs8GkJj
CeG0sJ1fdp3To6fMEZcpOK8nzwxpdwbtSQGR5oRFQrwxBjpGPHgNhbFpYFla/VsY
LYMxMoEy+oJW/rGWWMnp/hHwgmBIh4HkFDGHFqTrECj7O0xPru/q9dr2s+ISnBZw
oKs8noClGOKLk3OyZwy0Esym4oF81xUuU5lOdrdJjHoj2FIQgxhl2GICptEX/EaH
C0WbgEKbonx/UUVxo2Tpu4ABUoMC0t4G+j7Pzak/2eywhITzFp2MNYeuSuEhWjtD
ftsPuDxb4090XaKJtpPRZff0kWtlPbai3u/uFX/MZe8nCZxhrpLdgogiPAqq1rNu
zzCd3Xh9azuo/a4mzPsQA9SNfk8N1HcculQ1x/3+/B7BxqIlkOFwwDOZnSN4pL1w
fz12qxi83ol5Ye09eVk1gcFRQZC2bmfgoghF8ewAGDCe9VLoHA3L5GiVtjOJih2u
qcd4JDpvR4s/FZbzxfnt+mtgrV5ez24hACbZpSVN7nFiEpKigj8hargZgYzKUq8F
fCUPUUk9x9CkNwc8IM1Cu9AjEwQJ6mQJAxnMOnW1uMeAlX5VAgNnoEGfomguENuq
yxnM4k0VZmq93XwGSoEu37yG9hESzyCwMYsU8bGHQZOCvdDruPWE6cnaAZRiPQy4
hFhfPw9u9FMWgrqNPCMRgqhro60gvX1qv6+8XvEoH2I5GcoGOfBjRA+9k3S1zo4F
p2XND0zqmatoegqU27C5Kihj/Qxuj/Ul+Mr0Be1W8ERfF3FpjxmjAup0AuxOzJ7V
69+KGAbwyBQK5TP759ZX/Gp1U75lwe4ZjZidHic/taVLIYnHHEkfWqHWd9iljoMx
6BG66jB3WclSkJ8cS3M6uPrkx7TbqFTv2vcHQMrBFwzvooe1HpN7QNGGIslRQt6C
oO9Esok+jEn6ea/rFGk0xxD73GUS5aqG/Em/HzxGcgm2zOeWaSbpKxvSXZwq95XV
3i3xrf5WKFlF9a0exnVbToO+hzc+Z8GACuSlhK8YTdjf5QeOEuJX+CxrkEZFAmCC
5J4+lsmr8HDvSOBxb4FbRirW+Dsvm6OJ9CsRc7EMxxpuWDYTZzb0DE9CswLqrPya
3nxeH5Ojfd+SmbwyYUCmFxmoe74uoVSoJPWyT798Nc/xJbLo+9UDrB7aaT5l+1fJ
1KEyNGNaWvjeXcCgfCeX+18WJjQwEY6yHKeI/zz7kB1bznar8w2+QKhj/7c+6v8f
5c0G4U8uhExVCBzDySi+DRXKV7Bmzl27DZkYM0+ulkW/e9KZ9412OaCrI9kgKVBO
VEQxswG8i2qUIeb2iJqt6lARu1O65Oz/gsZZHUtJ6G9VZ4i4U3fz9JHftqOlb2jr
hKBPRn9kFr5+MU22PNxSmJ4Cx0dl/lS3xvgdBl7Lvto/djtzsmPhnK3IISPybRC8
bA3A1TICCE/mepvkb6489jxDfK+R1FM/6xpjVnmBhNyx6GykmAvfO9GDAYz/iPnk
1j8YyWyE2yEn+oSFl2exzPsajW9SjUu/7H1Uglz1hC4DO8kM7svdqEXbTfoF+7WH
qZiHDBvI42iTpcpZ4NcWyp8/6y1YRw458CXMFAKlhV3WmrDPUdafwHkaPiwSFdkm
NC4JyS/hUjcmZ20bBMGKwbf1bjWWzCWvMptrRGQhi7SkOAhizcXhaZkVy/mOgbCp
9MZKpENtiZBp9MbkSX6n5x1FLY4yTgq+0hKNRfG7JewhT4+E2OQRmMreY22+ttnQ
1WCYCn0etqleHKBf2DwnzNlfr2Dr2JvEVLCDLlk8v2T3fj0+PPkd3gl3flnXKAr5
MeE08ImSz6GXIqKfOtIBrzIFt5WPEv4y5kNw+/1bXodAJfP/ipuhmEYX+Mtjr6z6
sIx8O/DuGs6ro+fQbOF/pyabFcgvPonIG3yxYW0ceUvI4xh7pku6rlPjyGWbr4/H
oG5UJGAGi21LgZq7m0mAaELKHWAXEl5E/LvtNAKBOXWYVlfWfPkvapGiroSATYvE
aNJ6g5gjbKeKGJTzL9r4PiUj60tQyrABhZoIbV4OiRE7w4fEQMkQfBq9yTatnYpz
UMx8MSYRU3+KsBhFQTSpIRlgTsKUpgsJblFHTW5YvOHEkWr4O2kh571RNgNisgSk
TZhuenyZYCOfDANHqSbbY16GOmUOQ/KaDzt+9Du73XjTfICfBJRbjZBi8NwSrb6D
TYtvu9WO4Pwh0JZwGmEIwU1naOlGpXIdiRKX6Gd96Dwy5QUUAc/zStsuAlh/6PDB
a0WruIaiD6kTfiKXFqUPm2Pn0RpO3snt3QEvGrCbRftkPbLGp8MlPA2tDh3d/pSo
HEY+I9aQGRBSRhqxZjhLfeWu7dVofnvPJcw1O22TltIdKd84N4EnUZensEDCivE/
5yqvz5VfNdKtreBPaZtqwPska/37jM6rAij7GHPhhs3kI4lcL1zIHy8OT5Qvo48T
HGwaPMQCW0Crrl9FLlwt9NwDfdc3+l14IgArXzqcYzm9qT/CfWp3tBWHByPxqnz8
GMPUXL49LRavDiCbGZwSUcmgW4N/ej4SBePnOjQHq7FhjD1nJHM6ihAVIoOj1mMy
faDqG79T7nuQgn8lk9j2DMUQPNoQUZ9zV2AeEtZ0rFXvyI3Zsm7GiFg3gVOmOsDJ
y/I0WcJv0KjsLuedxQHeWls+uvVQisQyAA8hKk+9wS8nbDEcsuG5CHlaIe1QiSvY
3rTIhmGpI7b9dQ0Trb3SSU1lEXF8S8sUpi5i6+qtwISWxtZoWhgPJNfMoog2EFIi
a7jdLr5PEmAhRTZnoKLsl7AZi+tg0/bu20PFFkYpDWFgg8q4omOly/BctwfA6eIO
0qz8hX+qz0ubJCKH0dS5NhsynGUYgz2jmWVa9D2OFQl/mn40gl86MJiPnx45nov+
GIozd1zPoJluto4iFudLglfYkTuVWMkA8myDPPiJCBDNe6pQyHlKlone3J75HS9C
g87qhFOML+mDlOY781kTcEFlCIOto0znshNKm2ahZGdTpd8C3w0XqN+ONB+FbuWA
Wp788UPAHJjdFmpo8slwoFQ0lR0mtF7MmisPer9JnKjAStgTRG1KPPPzPBJ5W03k
RpidT44MpxF9ayC1aXWgRn5ofWtinGiXbz+66+Cp1WxY6cDPg3vZeKRWPZHkQ7Yi
MEnxc8+3XpJhC1xkPk8ir+1PQBgNrROf/p0zGrl+Hbatkf51dK5DUdczv2K/F/DA
Sw1xMsCWpFXwVQ4L/PIXkPVRu5FvipTueqe7RYdH5ivtE3HegY+b+vOsLAVLrbay
6cDoVixko+1IJXZDG321Sc6nCOxfq7Xg3zhLbNGBmpuopFIBXiHVsbWA0iVram42
8gqe19FvyKg0fCGSlrwdzJlOwrvpnGXBiSbGwgHoh964UoFACygYZvV61Jc2w0Hw
M44LjPeqbyOw8wcczsCFan3jVlOhy1AqwIF1415afyKUVf2wHhsp5I/0AS20Y3Ey
1X0Tu2klxqzv6wt43SyYMJ35NgMnnnkjkyJjUUgYLN3fV7yi3pcgQcV/J6U3HvWR
9ZId0Zzkehlf0uhl+A1KR2KVy1yFHNhkhP7/Bj4Qm6z1BM+eXMfDbrv7KAFSymra
qHaJXnJQo0azne3NDzo1RVtdh0Ih0DRjKwThGZjhOjxyEbb5NZVD3+US7jk3pFif
IPVGWF+KXmBQjD6YCbm4FbSslZR9MQryDFqq8HZYi/h/dUroGaQv1XOCWRoMQDi3
Hut+H0G8yyNCn5/X8A/cXiHvMfRTv1EqhYfO7o4L0b2WChz6c6idbvz9qe/lF3VR
2OgDNlnsMltqZecQUs9DR6Sh3w2cC4Wy0X+Fd0OdlTtXTvW7BLdCK2Bp4YXtvuJ6
JE/yj/nDzWzffOU8oVEECt+WPMmyRojOCINvxstH699ycOdFLYo+pVHlUGG1zHjf
S75QUIjnUc/S2fWSshL5cUGjCPYecR/bGgKz9LXsAHcfjwExv6efFUnwldj6Sk4M
II0T+m82fJq5oaVHVj4igouEUvfE4BjbBUWoghWPqA3p3FsNHMs1np7fH7waUrRE
IXPTJUhqKX825a0sBdgwVJkdDN81n3ytVHBEImOhO3rXbLIzXpa7CRd1fLXiJntX
UsfkxrcBngExAiE2tzD9EKl8HUq59EEOa9f82hju3puBuP1pVZ7rnOdsYR2jUZBH
qDz1GpixBwxsssQZi/vHGdmkSGYAs6AMgUaW34MFuxdegLPCJ9nm38OJSQd8cVhZ
nIaInL64wPkcXFF+5dY/DaMbqdzD3cww5/EK0Dp1dR+D53zig9rP9lcPGEZlLeMt
ADev++kjzqY4MS+PLDsh00ru5NJ0qMopff2F46462mCufWT7iuHXu1qJgkvjtg8x
eHmlbpyemF2HRZr3QyfzDtMvNBhDiDlDIew2Z0/gnrEWf9pounXbncgpw/jinWRE
O9Ak8TExDhpGILZwlue06Fj24efLzf8p6YQr0GFNyvYQZbhW1ojR1k6+zWkaLsJG
QVAxnXrUFR6M+lmwCBk6cmq5NMq3a0daIZt7H+13n8skcEL6/Nq+uSaUra9QUmWz
FhEGLICmvKlFgyAW40GldHU7GrCUL+TancsNFOM/ITO7TNTOt6Mk0UktWykcTy2T
4+ViRTktVag8LRoWAb20Yq52m194jf8Q3z6lFsUgsMfAo+n/AXLvL/taDeVbILSr
2LiR9WFyDI5YfptPpvn0kFC+iKA/F+NoEabQ2ZZsbQej+Fv/Fdxqfk83uAV3rQR8
hsl4Zc4FD+6wzmKZ6YhZdceK6UDcI376rrP/O9Q4JZvEo796Wj10OjsSeXkkkNIc
gsEG2wymN66fAQx1tKVk0G5/FIMblmnKBZf0HuA9MRADLvcBzX5tp/UJClGBfr6w
w6SSSZL8MzA58urxHXATKo9kMMbzIndZnXTwx/0s0tM16ibS8m9U1Ra8iCKSoksJ
eD7SSGs9BxDhAj1w+lPCseHQGyIDaz+pP49iAB5A9/KIUgBzUWcnRXdZNsA0ocJl
PUrVk4qwEQBKlT3MCY8JuDUr6v2DEXuUApR19IvOxjOD77Tu3y5HEn6CYt4V75Bq
KuM1qfQ7axonXFpH3yCHyPZnKJb5Um3KyWJSPnlcmB8aFAn+7pbegIgE5XtQJaCJ
AZ4gIClHXXrI5yQI/mZVm0PuZ5SnMbMeWGO8uLzL/zuXBKB6u7U09OScCM/tBQL2
TRwTH2Wz4S8vJvKend9zEEkZl+7B43vpeRcD0ZAUyO/FbnH6R7U237d1djO6/jiL
srFM/gIo2pk1HVXV4VkCjF6aTpj4esV/dzAgUKAq6ztXXMIF4+kEeHTjn9je8GzZ
asoiNJr/L1poqMlRSSMvRYhQJIbtSyC6UgEKirIIvYZMg3d8ovWKUp23Hjuj615i
Y2Vl4RjMXyVbBaIS0cNCAuYZ26daZ5uVHA5hOk8l0ug2a0mujwkwJsLVA4swZEwY
BHccqZFSczT6WZ2RxiKaqMG426cAPW1xo9LO015DnKsjIlBu1wJCxkmqNMlW4vNN
mv8KJXoj2WAH3LUb3czvikM/ndGn8RJzMuB5Z8bjMJ4gqOiM3rcTJIYZsO7xL96u
ZXlCtqcaafOZ2kW76k6un2oG//oksa/b/Vqefcipjp2geMtSl24EjbMHY+b3LOOa
GTUfsTMoGvUe+uDKaNTY1JgbCC+g2xHDilwTjhjWiRPHp/QXx4lSoeUHbZYC1vdK
mBNpbjs8BRRBvK57xFsflwPcJcJD1tbmh41hh4YxfPDi4ZeIV6ypro24FYYoHRA9
RmrGeSVi63+syZ/KIlfiZa/56XxQICZHJr0mx3pfS1H8gXoiNAOr9wn1kMKGsH/k
tvUjbG5yuSHnKpjOcbmowjefD7+/SWks/7qQ05Crj9G0L8SJn/+QQkkV7tUFwmto
opCWUh7hmpYUogxE024TDaUMzVeg8LQcD7exWEKg3/DVdxoOkEJUirebZCxAfosU
YkumBN0gxEbjO1F/1rbgHZ3V8LsQ/eJZKHzsMrVuWlSKZQZkjDk2mzHqQ/3jMdOV
R4TQlwYR8mrJOhnpGtfySaDDoMzWRX/GTfL0GIYCI6B1l4t9FLIjOktpBmN9QGgL
ZSHc3swlvGdh39QW/yKe7blgQvqDuM/3ALvYpOFH29TZlVppPpEkiN6of6xFemRg
/1UQRC/vZ20HT8ac5GF0czjhtVQDVITSYQlX5a2eDLe784WIW03xDwL5PkXFUjNa
tfPG315WrthALv+q+Q5xtIZ+y1hfxTOOHjAySuBTtKeaYQjzZPQqyUiBLWNmb5hk
NPauPQxBkJ4XTWy3K0WtOk0AVSfm01D4CoPaYrvzlzMXFsmQottGQxwflrm55wqX
JglXRcWxnDJ3QHc/+oATtEHLFjfL0AE5pT0e0x+YD6MfktbhdVyEPNJPnHCIKTbS
7+CMWF9DrwpMEG5zgli+aqbSLfnoG27W7BRy4aAwD4y4c0jCu76rhNcTbxBRr7Aa
PxzugDQ+6xh22EJ4ImrAdBNGp0NPMmV4ngplpSRtiPPB4/42pGM/v2GELhJ8JG27
nSYItD708aHrACnXm8VvYO8/hwsQUV3ihmhSeRZ6/FEedxo3uEto+XU2LQkmzH/F
ypXnhKz8d+odzG+lXPSm/TEPYpZReW1mfL5FrVhoUO35M+JP1JuO78LgSx7uiyZS
+FcszXZN/zVn5t1o81l8n87A9VsRUPqdKXTeiYV3PIwEF7c9JVETdLqV9g9fOirP
v+w3alnIQJPEZUUmvqsVEyJesuhlria+tPlfyz5f0W9zdIQW3Z2xiMbnzsOLesko
sk8xrhHd1Q8IZ1SyQSSiIAWrc0b4/iaC3efHUFO1baw6eTgbP6TRjfqAUcRZ/AC0
A+rYehjY1wzMpNTQChyIWBrLD1qZ/A+58btiWDn66LMb/S/CWiaRXkkt9OrYushf
FwfyeD47HkLjD/Ynp7bcMzzrs5hhi3qllYZrV6LU1kwv5/wLsCLPepRvXywy5GnZ
ATjKgQbt87kAIaMTPFj86y6pEzVJ6ipKWepE225CjqUEM2uzop3BqVtih2XYq0A8
5cV++C3XmLqA46I4Q/M53Ffw5DnPQRv8E9rA57n9vXxsGTIzsQyeBrIMLKz+7Ymx
pdQDHxVRfZNyFYmyLiJInN/r9a/Wubp3sP0mmeFqOmR49KDoA7/iquG4z4FnmEMa
slx8NmoZcZHWRRU4ktAHiMdiHNT88n1pjwhQ3pQnaFUJKo23V5i3dKx6cFMgj8TO
WQAbHOvmKRT3W0tuQyHAwIaA1EB82Ze5e+TXl612KG+W3hc4U4jtF5ztqGcSjS4g
IIEM95mRMouLBaEQ8vsFaZdxQe7zwDx/fGkZqRkCHq6e6FLRQmgDgfIeC3lNZ5Cr
dFR8Ikn46o6p3pA8xSauVK0emVuejaTjR79WVg0cuAgghY5rWwRT9kobOmlvpY1q
bKg91YFX/dSAWSblfj4gRCLO0MnMTkHvETg/6m+dyxB7zPljalfyaaXGaxMep2j0
pIBINKerGYCNeLi+ztKW0DByuK5YqzwykCKERDMz6bhUF9r5the004Ppbcj+mjGi
wZD1lRccru5bCn6A2E8mhziRTXhvcniGKI5++CdRMWPhgVtSLSdVnIghsT12uJN2
HlzQaLqNakWMtymdMyquTFNJBJBHg0uV+NEetM+Raz+y1u5A6r9e94UKyskasm8p
3tSPkwSMNnWqf8lTKHWl96w0CJsrv3mjbQQR/ERG7FMqgKyabeDD/2aqchQ8sRzE
VIXK8IQb98FGyoYMn8U32XrFMFlkcTRUsJQN4YEuvqhUOjRQsNRHhuHe57pUh/xW
465iM9G3EB5kFpha1sf6qxIZyrehoQJFRnNkXBLlT6wOlM7nEjntIEOjsoqdcnUW
rwLh8Y3rM3WBw2AFhNcXOAJR2rsb9V6YKQxRsOO9/LkiJ/FlEn7W/2YDn1G4TZP3
7P8+Pe/ORFGafDgGOhRECjJDtZi2Mp2gv8I9ZyzYIbg5TreZ5EqgIcv7AeQkgK6I
27oDEQ2LGun/6Af6QS/Jku8fx+QX4+lVh7MHiQMReszgs1Z+AenPmKjq7zySyMHq
cg7aOQiE/wcn8Se4SqCW9kHvKTBymcnbBntBWF/aLBsMacd+H10dWwIGyh1iMPHv
0KY9r1ltj5zx1v4T9J0frulHSZ8cokXupVaDfVDaXRdkoogqxuihxeZESuYCly3u
/NHo38gewH/VsOxCg4ZrBoW3dz6Q4Mo5NaxHGRNOLnPbP+/5vj8AJfrshsVYMIgl
ZYC6kzVmV1KeyKJBC0KYa98/h2cPJE8UON0YhkxfVdamo92m6yDYysDVRe+E1IPX
tY4Wch0p6tTLLHxXL8EMoplMepHvROf2wKljekSjDxewbo72roTcA4Omgwji8CVk
jbJ+L2A32/yNI18QvN2/LJITteG1p7Jpy2NudfqDbo+t+4ZllrjII/DMpYx3lMKX
WUDvi8QClzIMAnwVQetl/P5+7LGXcXDZNSf745NvTbswnRmqvXZLxE7sA899DlrD
BTTqMUCjuBumEATwFSLINBWEVDDumIc8xdwrJYgjXggaz0sEMo0d6gtA+L2p0Vkp
aBZmo4VktuNqoerHpdSKRvVXhoJJPnH8sZ65ZsGbQ9A/Eg+oFPVzqgzkDpt8hKiv
BzhFkr9rxDO1zp+n9654dTBLd7tvNaTBDqFMz5jte4PT14sQqq64azv01TQ71s+N
+GGeqYjaoNSTk/11e0s5UOH8MCPHL8GU0xVhVWCkcDAVWPY0NIr87MBcNw5NsTAM
V9J2UizAm+BUZ8YxxxURDbPHJdqUU7P3ndRHWJL/c6yCVvC9UmVoZlGUw70CeNMD
GRJM84N2LT9GFsielZtzzlQxTVEXbYxOezyTAu0wfT0pa7bDgNmCqhjAYDl761ey
KEMMVIs6ERxS62OshPiWTj42o+CWBT3+M4G2KrpJ9QZ91t3VvToGR3lEU75X7rc5
kOz2QRKZ+40gLbsSyrYhyj1J9OgenA+EDKzFVbaB/AUoMafgfDhm9H+so9Y60L73
auJQZPKciv61selR3MVxA1tYtbUbVrMbm84kE67diBIz8nDbkAxOg4qRjMki24Js
GvdacpjVHBJCe+SKnE9z4xQNJA7yEQdrAy1oHjncEFy+ja1QzzUhK4epSMXpfWT5
di7ZGLA5xiUFgjbdI7C+Mr7BaK9TESR1B/Q74JcTqbGZIAftau/dzH6ZCC+FNT+3
jfvij2voAa7Vs6Ru7muh//o0Ns7osqQNzYgJBMEE0dTYH2OKUZvV2Kq4f+rVTnU7
XR4oWhyWumdlBIIGQmOx0oQ1IN0DO5e3nrrRKVAdejGoUwxLnIFpJMuHSRYiwhvW
Gntyk5qP/A8jNRAezkf1A9mI4w+tUiIQ7dBfRzEHhuRcRFzVBu0NFwpoNPqlhIjn
NoxNu9DTeoL9xTiQlqu73UUMOFNx1OEgRwEyvB1889WiFa9oFEN0E0Oe197iFQql
dSMDp5R3AJeQBZRYx/6300Uci5Z/rtiZVHE436VACy9gvuJFcY9fOTt9HyM9c8Uw
LABUrmMMMVci4d6RFV8+MBds7uDwkqtkvzAvuy6fX8+Wl/caVsbu2FABtNbJE9B+
9pkH9wSamaLVmfGNKeaQXTKCjIXWpSYue11Uz+MC8m3IpyoQAXRO9HHBiv8ztZdZ
joBavixnQuRNQtABhz1Vi0/erUOkG3uCylzSyiA5eOvlRHqhC9sVUKXzPn9di4HS
872rQ/3SsKguOOyIls4j8Q04j0ohexrHHb5e+ziZN7gbAFXsV1C06Vvb8Lhkt9o3
VhpCbJMsybqmo9rp77Ilh1XweU/TzPynqYPEXlsewZoljqu0EcOW3vYcPlnVeduu
9P6AlPHBB6dwc4WRF6tXNd1IM7xdNhUuUKdKdE0ZXAh+//NFAAsIX13PrhO94KMB
KqO9gnvRcgnoQHKfKMIcJDIvYGkURGvyW3OAjdvSqcpPbg3pS56vrvY8CThn+M0E
qHflu/JbrfjYQnQ8OezxSMIstQ/5GdQlO6B2bh1Kyy1/tg2XA9lPYcmjsHhNkgg9
N1EXn/6HsJLPiU/FBfeAgWTxJAP0gIEBj1nsO2eutvkYjTmCw7b3Dg13TXC9mpFL
SeICk3eaNm0aFmnaZAGKBIBzS36SXuJrcJ/slRqHohSSmBTAb3M5X5ej3SCep1UM
DOYorJyUUwJLLOqHwPr/YKmqsvf7cPKmp0t115YYJl2OuweHLokW22XqkDiAmQkm
k2gnA1nxGf+CEDbiVICFd/0oWLzBbPFro8BbRY0KDPEgmBg88Ej+BoNYh2AS4i2N
k2RMsIjCjNxd7FOs9TwuL1RKAEh5z+8fnuMqbTsMY/7C1ekCLFmNTLRZBtLi0ySD
FBWgsj1eEMOMujkm5dQ0O819froBUHPdtSjkd0z8wcFuWwOAVrxgJ2j4WI0jCqWX
ZiWK8CKsq3Z5n66e0YR3MI71avJSGpgEuQI85EHkwMEUA88itpBUtP276YJE7E94
Y9EQQd4G6TszeFHpVG5ATCd2qB3hyko9l8N3fPflv6SqLcUszY+RvL9kKbwvxaxs
N2V1wCVQ7cX3kgTBpwAKzwmAqYAY1B574ss47XMpks8YYObVAk4Dv5qATEfbtwZY
4rS6KPKTIlsPxRq9hQcGAd1rxayPvMFMVQY8ek4GWmg9kOhXB/UsPEnAOXuT3Sf2
3PV7VHLSKZaOxt4qv9eMFYmIrlb6x1Fnl+bT+2L41YLlt5ojyXFXv5hMR0PJe+nS
A/TIkOKvlv7wW457suJ3pAMfBVRJKodiW8hT6ysS3RExMsaTyAR1B/CXDDwhTEbb
AMT616vwY8Z5aut5uw4eLIZ4NovyVhg7BAOEEoJ1Cx5vkUk+XlFaSndyEbMMh1FY
SeJRoB8VTX6z818Mx1snPZlguiwvSNW01GMzitAmLLDEKowj6lJlcmzgoh2TYz24
iJ6O3ux2czRN4WpoeAzE3lxyPyHffSaIMGohwMszW7KX+gCBJB/2oE7ut+hMEq0A
c8QSAURlJK2sx4bs8K5WRdLBZ0zTrNR/3i0rDzt0SPU/CnFrDg0ApSwj/pry/E9z
hqiLF/HQAhl3uVc1NsW/gF0GzyfqhKRvtA/IUe72vTm84bKzbjARcWmqU+N7AXv3
NI3h/qQXuFXB1ggh49r+yQbiJZrIu/BWxabddAHAsxocrka8frbTnvR4s/YaXtgP
WDvGThm0qYaPtGbERyGsEbjOnR6vV0uucIS4WU5A59JczWidxXw6FKYiqg1QsmKk
7uNkzthsopVxNYz3JQ1cdaoThKAQIen7D2WKd2XFG410vEzfieHIzqp8yHNlaudc
2T9nIy1Y+aizva9iiKohg1ZOR+4FrNt+2NYn0W8kRth2O+rohV15s7niejAI1c0L
hLG5mfk9Bwqvk8sJVL/byJRrLld54GVtQNgqS/cvP5aST4SaftCKeP2oYFSMAS54
aHgXBByPlxUtM4i9JLkyDrpw+oajfUcyzA3ym0NTZdc245XkN7grj2mv+75guLZv
uEEZwJ4lkO9XcLvNpnHl9ApL/lY0Cd4iHP//7VOhaybaPNs4KV3/3aRNWzPufqRT
v1ZUryQskF/IZbPJfdBdGaN1hKZAK6Jzq3mLPEMmpjRvVMiCkae7R6bkCYMTLObL
7E9E5788WHvYEiH3i3kDXZnUI+284i1k2eeEYLbZzr4F7Rhn1trjB6b7K07jVBS5
bQpzIskTyCuVzwdph4FFnAwrP6tmyeJrIrrHqmhc6IiApZpbnXoCtFHdxvaNMMh2
20t9s9bXeqwbV8X7OYvylUyIt3/s2ps6EQwIdDrqPlcNWam2D/BkLLtaeq3g/Q+Q
/VsdJyKog3OQs2U+0osu9iQ79qtg52UfxWiJ0slBOMDj1aLj4ox2ljCLLuVkazQA
PuxG71MFBjBCMjKLxmioJRn79+1eGxPRJ953t0MMsq9RpFM9HcYBIidF2bKhe4m3
AdzTrH1UFzh4eLJDwLgfXtJoBhZkqOiIszpaQRQCkKepYxnpBrfTbN6yZC1IAUOE
QsBl6xAKSxExULcAmSIZzXolsgjAMbTfLdp2xaFRwvM1laiVrgXBLrdTYuEg88Hc
OaSp4lEqK3CtOJ4XuYhUzXsPAdnpoNyv6LeXUXo8qSZvdncI0cttDTFMDEeqDRkx
EWn2AdjaonOvvokcSh7Q51F2CNwjoWd+PB06WA1wj8PiqHcaxufnD6qLrYqdAzcp
zOm2lBy0/c1nRggasdOBIq6BNWotXgJa650PstVBhiugA63fkEHaZgGZiyDXrytq
k/5xq3ZrjFMrK/MtLngmYVQ2eSbzVN1qT/PDy7psfTkMAOtH6sCFFEoNbpGNZ9Yy
ukbmIRclERzdmg+5JBoRVTaWNhys6Ttzxd1Og4N6AZ5c2TGqR2La7xFVXnrdCIMk
8u4b/tw9eRDOcduP0fwlC7LNK6OpCKgEOrMy3uL0TViARbBjA4Dd/aPoU8dMjU3x
CooJqK6xJ5FAbdEGhlSaFPEooJZDAGk9jT2EszTtG0CrQO7lRxql04lOvPBhOYo6
o/grSAAY8uMFJQiCWc/3SyqnS+F/Z6XvGPh2yRE5YrchICRK59HYTXvmIIlvPofn
QqhzI4YDbg31rKNkovHrxvkKltczmVb3ChLWFrnB5C7AV05/N1KGJ3zB/bkjYaae
ZjnRYEk1/wH5gs+keAyKB4Hdzrd7TRIKQLi73ScnTWxtZljrvbPb983Oz8l9a45x
J9RlHPZ/g2LNDzhFUrE9OGjOVsryWPglaDDy1sTZwuBSr8i/zqq9/IESenSEobsa
e/9oFJ9OHDuCPdhUiIgso1QKOLYGGXrjkGHbkOKQzNp4l4/O7Py8XoC5pOAzhGOH
L6bDtBp5ckwDk0RgNKvmYNxNs4pNw3anSbybPrdmclhqrHW3jvBUFXhmBxx0WjMn
Bg2KLxfVpR8u1tXeW3v04OCifxtHfSX+5rsrdkQZSLxgHVWQ07T5P7JqiIRZBKnT
dBjBIMAJanz3QUZbOizVbnQM5gqZdyA2w+ZtMZMzZYAA3vtBv3W4Aq2VlaRNwhEj
75XabjCzNJdIg531U30lVmufRrs1TG6uPnkJSeZO1MYQAGdJB1iqWHXRR1t02mPj
OLyy3BDfKWN43yTvt82IFSfBqUIZF7apx1IZMF82xystTf9LK+fRW56Hs3qedOop
xCDqSiGyaWpfamsHF9yUzG1SZSBxxvQEesruhVdfBxEcYHeOapHqg3AxOTQyH4+m
benDJFyzaxP5kiurwbvVCcBKJKN8SjxzAboCDYEPOqWlpB5tWB4MDE04R5xg0USt
MX8aYkJqKgVG22mIsC66+FCmzK3/9ypNfq+Ubs2JcSCxMlirsrtMDNpZTBomHgTQ
pE+5fVA/tadIWLdUt8liQlZRayFuJw2sDNjDvPLJPWs1780P3WEdy+piqszdFk1q
Rf7WRG7Yp41i8SnOqIqJLLrXGP9G3wZY9TFbkkM5pjG8YpTCaRqO65u2V8MWYnzL
noC/GXebKoxdXJ+sJiC0Hm9QmvmMYB/mpPMyx011/mT18l5oDlL5mZ1EU7zkP/x3
F+t4u3IPQP17J+oUu/R4Dz2AjvhTxbXCFJSIVN3WcRezHk1yEMD7obH63/x/r36h
UZhTGcmrB5kcAcfgrT1qP/RaQFHXBjTuOZpGUDuHpkC1NTGCmS5NoNCxz4Ii7fJc
3xzlKd4yoqnSL324cct6BAgd+DE/1+VzLGfq8B7s3OXrgE7eTykBgLSMw2CGrejS
YdlSCeE6Q3ocgNxn7cquNRF+eDI4O59Cue1WeOPCIqO7thr4vsx1pHgvE5Q3pjVP
6RJSJm/KmX8q0w9dqzu3VyuICP4EIisIbDBrLZNU6uNOrGkFnNBpbo4duFZBtnT3
6GfIxxZTDzKc9KOEOnr/3MGiOVm1OSa8reQcghSqnEG1Eo635hW47afG5njuz5yz
jxQVLrgJTxr+VXKwjeQ4Dr7YPcNEs9Q88d92Aj/jFpdbVofMIKOboNeFPGdsme/3
STkSC7LqanyhHAUTaF2faHIhn7nKnRfOjLeVMu/p+/CBlH+8tx4huXpb2NrS7Llr
Uj1Gx7rJw7lsns2JoAYiR5up1K1fSQbfnBZukEJemHNbc4aQPTC1aruPTD270Yz3
VvQTPuCrUpOEe9keZGK80gB4bzB7qEGYVetyDdtHwBJSgmpVUGQ6MbYcE/eyjSTB
BgAt8fv+T7jJEg0fSLCZXszRSGk3S14h1Dddqsp06P4Gfoai+7H/7Vjiceg8/T6N
Uhd53T3j2W0mzGZAA3siThrqZW/KaQT5O/rP9DTVrD3PQ2M8shfdhKEJXEyuxtO9
N0+A+dNvNSKNeB3jSyMv/sOLfVpFUvQkN7Xd4N4sor3AlK/CWFNLDICuPXl7NTXH
atRdfEPMWQ0iVJLW/ZaydulUUf4dCtiqx39+/38qc3AQayrgxRx8T8rKQAjrkJjQ
Ck21siEbZMTGe3cQQGyDDXUiJKSmzTzEDR1KUmeJjVCTi5GfyxltUAeQiTCm6JlY
S/irRZmMOZwWvcNj0iiMCEvM4ktXTOjmjG3tBrw3PJRQHQ0d6hgQRRJIWKr2GGjO
7/sUCAd5angGgPbPsCBcBbG8I7DEZl6SMKt78wwZ4x8fWLMIkHQ8VvbM+ly4h9uz
OUD3+qmgg1+lsGglMwxXtEV3zvsQaVOrayN4h/tSSG76FYLQ7YQWtZMLXa8YqJdN
1um4lj1Zn/quNIL2shJtdPSPafOIiOdg+uiZ4Nmblsa6+3WuEmBP53X+Q2VW0UKE
NKSVnHnJ6Qy7BDfIngxiqSb9nnk2WCt5xByWZf1UvjpNkHIAL2fZKPUUZTvmduXa
DFvnScCGVD5dglNmPkYa6E4gE6zx2yoOifpFzGVjiJ4NgGZZT32fKRQVpXYmUM78
OH7YmY92j5hMfENZ8Hy0Q8PXEo3P0rZ591zooH97x9DjgH2dfveYEQ+wWVx0VxRA
lqEWPkYEHbE4+dTnc/pR/WmPl1LmP5ct3cWdcVduP/miGSLwwBVh4Wb1tp9gaIRO
mIMBF43G+qmLAnlY+02KT/SSrQnQAxrDdKLg4/rT0MgBYpEGVBYtKizQcVI7bdCT
ltOvkxJmLjfEMROlxRS7IyZ8ph6Yie5xiUXZogrrWACxsMPNmi/bmYvXonowMwYr
cryZ0TTY2zFM6nNM9sWhlzSu9VNSV03YAMLbQulLh5dclkO2IBtxe7+yT+G3oXSB
THmah/A1q84FCwRwv7hmIaMLw/UvvqVXQ/uo75IlzNLmpchMT6rEe6+cidxKqQVP
olOABAIGnDG7G1uPn503UsRypwTqjsn46b8XeipeqjE4DpefvolBhYIoe/nqCSMS
paLlKV/hJo8MTbWW2dDyg44b6ob42SrcrfH1E4z2kvOHiZyrPCJsXvxKqHhjhzHH
lzz9fpiEFLoMvo4AF65cHj6O9Z1lA13pUzXkVVQu0HcwZZ0SXHT58FD+U/WhIBKf
/q5hsY6WMHQxpqqQX49t/gbvZD1soozdDlZzh10CJzLkmJ/n5XfKupR46KqCkWaG
HuPSGWpybccyhJTxFoTIXVDemqAsR6euVJaf1+naK45tUjYNDqVLJoaDhF1kk/Xd
ldgP08pPwX/xArCbAqmUDr+L/97yYSGUHneeWbd5R6Nfhk7tJh2BziqnVIuEFVv6
w6KN29zQgYnXzlgBOXLXqjXmyoUbBWar2DkPWu6oJgf+JQGRtChlx/fF4mgVe7SW
FZePJcM0WxDAkimxt8swZ0aXWOnZ0uOGdDQAscXUr2BPqgNF9HhpW+9bvzaqZyEM
V1IPQJyS4XAkV+w1iLljbjR6eRGJ9EVQlz235O12k08j+Cs+WJPe+mBat8tQkaWb
6vNE9Ja4DfssyxMVYuAO2rtpf/On/8okyJ7A7iqP7gUd6HDox3ZpdzJ8ZXP1CFlx
x6CO2v0nHjO1UidJkEujg35ucIDzvJDVSFtkYbH52o4KvP3v/BG+qDDSwibtV49R
9S5YbOCVz6ib0IPgg2ElWwatjWdJyz7GbxY188oJ3rna/k+c5s0hlVm4zHznjg1O
Bg6Q4BrLd81r4gHoasInJYnCelSWfk2pPYK+InnvMhZTkuCU/ra5VBNX5LOpbBph
amsK5iiw73WR6iZUsiNP275nU7Eurpo/DOGaca3V/V1/iqxts+I5vmeV05dPsbr0
EwnrpfUVkFhqphcda4nS16SA8wwuI+iZEZZ1CjAaXKfh1kEwsNLBUbFDgRhG/OAV
C9AzHBg5CE8U0bzPY+xE/uRlPEAWd4gU3TfZyI1MPcto0xAdtXvTvK976ovUzYOZ
43kFw05HD/N14tOyAXGCBFML3M0abDiof3oPQfjfneForl3Ah0425UOjRccSdVpo
AW+4lPsvQUFE/IlMxYvi+GDW62h3Wxn8zyYdLMaQSvEEO6k1OkNzDDLD652opLTg
Y42itdEC02sXR4TG87z2G7Qfx2zkz4flRbfojcufOKiaCbc1t2RHFmP7hzKXsdsB
EoBMttSO5q2Cyub+vjC4Lhmop34WD+jZO/py/zk54kE22lpdMz3RkrwbgXYWMk2E
fn2yPVCnaRG0ieaX5+JbXexvNXNXHxBreeyDaF1CKLXhMi5B6/ktVHEu9gPy9+x3
CM4Jy9TbUOBE0NNcahe1TnfRZ2Uv8Z6a7g6raxowrZFibS/Tlov8Id5+/dRb1otb
CEMkbRzi3cX040wK8i8W+RmzmoknSsOwQmYdDOpw/PaqoFfSgvtfhN7Zihio+JZD
fToYt2NgX/XAVPtrHeO881JT3MxrUU/IJIm2s/HbJWQS630D6qru2Zyz8ixmbJxK
HLZRNvM4H5hdP+UXM3cKcdOLj+/26vi704KTYx/EQA/MojzJoyuXdtzR9n240akg
ABvtOV0E4dNtYptGEZ3A67fnt0fYTdSrhHlDbucNmeqOHoIll0aqEQXNdezuzIDz
wlgWdkfGveQpKarRkj8x/5EQuWPbMHtcb4Wvm8BC8c13GtB/jiwQrkCVwzYsYw54
f5ZZPWDkpzKbgQOfBeiabnWwag7rpvSTZEd+Rbxc8Qr7re/ZyPG/PgLJfniR/j5n
FitmMP+Nhz8rSmu/Li0bqhqxhPJdVHe5UDrGbv3n5mBey8+jzdb4grvivZReUNmZ
L4OkzUo3YdkncQj/EW8P+tnDwrdvqluiYnXo6M3d63OKKKbNCRWbIQQ+aS7x1P0H
eP3PW+rQ3n5VFU54AATIlW9OTuy+F4rrgJj0W+TL5KkuL7qhMu6ZPt+xKjh+Egnr
taLzgJerBBtiAoAXqoaxnyEweUvPgzvZRheECE2q59vMN01Pmk/FOy/E4oqNLT1l
mIRv4fqHV4qFzpN0lGybIpL5+Gcrx4UlIvBjakkcz316qZADjaizrUqnclsYSH3u
ZNJWQHvuu4BdZIcGFvQ2Wcq/zyjgtM0hNqFiwHYSfLHO+dPsEdFVbpXPCAle4kLX
1zKj7QmSDgcFE7cDutjrj/GD//50rNLqm0h6gJkSawBAVmuQ/emLWD++FsxmILNc
KyyKS7AL+0BqBptvTCKcakLfAnlRBNjL8ifHxc+XhLUL3XCEYnYzs44PymbBqtsJ
tfH1c7fxrfjN1+rQTVbnNA8AnOZXdMlQ7B86l4JlJMznd4BEUFtpP+ArhwYrX79H
4ev/pLA6620vjC/tZtvKFOJlwXYKDZfldtW2YDllcAZDCnKJncbVAQk+GDvlb4Au
5S0mbj/LjxkDSPzRHVk3JD7biaHzO7Z+dvErf5WN83FzRtSF3CDI2IR3k2MSqVhB
2601kunB9NBGPerCfMZdAL4Qhd64Q1l7DerNjP6PoA3CPViLZYXbaeQgmJCf0DPV
RdtYMOi8p/rPDLy3lKUWGkVTkoIMXbXISXJ8zeg1PZsNLwvCWcSww9KO+FAVKTGQ
XYg8Rg8LRzMCpwgA274xhRXNV0rvfzq91XbcG8+5QQ9uB6wlxjYVo9js3ctL8+V6
i4ijY8xfC6XGi76tfVMy1ffCdQVsbzccgyorxpz+kx1orO2IXydVawNvYr87aIhn
gskgzs65vRerdfuj24tKzZEbp7EafNEk25mY6UoMUKZwB9Tk1ToWCoCoB6z4lvHA
1AyQ4BV5mP7Rw1TyuuGypf0dVbfFuRDvFQUUYvZ8NgDR8KXON4h0yTGWrThNa24o
5mWZfdTAsR+L1uqhKVvVqZiz9DGrEzLgtLiW6U+alW29PDBLfve6+ChvCWjx2aCt
sUHqqoIjPmi5kVdxXjU94pEwe4+F5Sq8FuM0GGh+b9fOiHpi+LyFJc8I3meSH2d5
2xE9l1BQ9ZpnnHySN61z5ZBb0qoaSh8XShKbQcmMNfdToOcvbAn+IToJ9OthuS2d
AHr74T37cdaS9kkEGCdIub0Q6xGvnniP2cYYx1gBQ2+LVJasuCCd7KMHFI55cptA
g2h5TSnaZ4euS2aR+fcKYP1yPFW/Qs4tOttjqfh0uCwpSFiJvs33pISsCt4zDqcw
gcd5Dve6gtYjIw2DsWgcL56AbRnB1RFqUxGGPDjicEtAs3Rt/hbPaaaKHHlaf60o
g5ltH7inKsmwTavBdaUllbuYkuuYKnKAPZemn81qS667XFXB8twbUDPjyBJJLqfw
aE9N7IZgUrUOpTXe363o4IY+8EjG+Fu4bNKT4DWcIrGeH1HiHTW6RqOtDroDdH72
ahAtMiYTsklxHvL24wVB84Tm61vjqqTWF6FrLLUxeDuCHaxKP2Fs9mbBllQE4bwf
MbU0ruXjHTAkS3jWsPIv9eERCjBm2f0VoEkQyRwzW8P9Zsp9kQ4fJKpbpIvPAFRr
KADCDrJvGzKCLLtGOK1MfC/nPbMnMXNKpAZniN8SChA7i8Gw8WlRuArnwhil7D45
zyvGYMaW2ThWJ6dtY5CGa3NFTjm852MZ2O4E4uR+n8q1pNnjKWwMDcT+pCn8qy6i
STcO6Is10LN/Gf0s7mnuXCGfd25H4v3mj9m68axOsgh0/zliGDvwQR9GuSJT3QI9
ocnp4fhU2gQGgv4BdHXav7EGZt3KuRPA+dz0TGA/DyPH2yiPVYRCwtuxd/BQX5iM
Rt3vel/3A6pSEXUO5A1hv4+uYPPCqlxiAPl67Ls8IoyAoh0vW3zyHNXUcyBorY23
ih8m5OIq+AMIDAGugNUBv+Jlo4QQIZTWxoOHFjFYtDKtKL4jvwsMT1PK/1MszEkB
kEAwyfUQKkQOP0r4TJA+s1EaZseG7BiuItffQxqI0eR5amxl8bzgohxmGYIkMOqy
K3SsTkCjs4n439gJpBZgXeWkEyKjnEWx+p8Q7jN+3hJPOEsgfQyRla8G9HSqPhaL
C9ih0Ric1FPG+bCercz4CNBsjPIKKk1pKdhHzpAZXDoaFYkdfQNIs9GRXHX7Z/ED
j78wKzCLV+0eBHH9gd+tkx7bS7bzXGfVtJ6G86THJf6du7VUJ8eQotIUXMCbLEks
8qwE38+fZc7W7kCtyXoOJi2SVSX2FvI+Bkda4JBgcVtsNb1NIfrisIQQZoyFB1Al
NMyCt4uRrpcm+wjH/tsAh8OOrmWrgc/mohs54brwb/p8Pt3M3FATLqSyoZh5OSij
iAtCMu+hLNr5JcUVN5HI+6nutgb0FFLTqcFkAS6g9NsrWKzPLeZ0SHjUdlMzGExJ
z5qPSHGya7OoXHkuCJQJXhBEpEdrHjFUPybaqsiSBv4cZDSJieFDPeqWgVGw/fiC
PVWdlVQRQf5B9VpK5os7xeEAPeY0iQxdJj6qOsXDUoH2vYAZCWhVijYaPDwCGXf9
cCXKkGP1uf9uJWSTOUx1YLWyaXhqkTMLUC6+t5KPgOmtPYpMrq/+b+qOOgkE/+pZ
872jZmgnoXhGbR3BFntcwwy6BzIBOsjarRUoevDBlQxJ0azduLngLprQO1IEk04H
oyY3efvb78i2pNGiFCXDTv/qBPQTQk2n2XWktTDp3a5sar5XyZSmgZL9SRm9GyWb
3Q2r5L1LLkqTAb/ra90CAZxkwWl1G0KGRVg/lCjV/Y4LsPHtx6eh0gFMBTtZg/aW
q2rubY2cm+Ao1S0e/9ZoBpQavWe4F/gGNJ3vuuyDVALTPQGcsax26DdF3FL02250
0ReW1SoJlyLqIliZO/+kzVAawE1M035rJ7RMnZ49mSgmuY43W/bHJvGghdJZSaL6
8QkAi0nOGudOT8MO1TGqM3hXRNflUZ2ik3q0iWYusYRFuKmxqC7AV12Ntphf7X7m
eRHSDX7l/6gKgSJwWh4aXXNZVqavxW4hwBryyNWlEeVuAzc0zVmUT6PVA3j9rryw
gLcX/E0m1BkkS6DRl3WDlVMo3Z3pYHe/w7K0YwBabMZjtumsh9/7oJS6+yc0iBC/
T5dcuMG2EPqY0UIoshJ59Srw3EEy6EVa7/oBlofgyvobjlkArO6tH13ATj41dZ/v
R2+aheQs+fWtbIozGrzV1Gz87ptZI+H256/2tFzrlQtuQY6LALNKd5110XswBSZr
1GnX3U4hTssDpMkXP2NbSHAILt1U0+ZjTVo8WYrjE6n8p8u04XEuWJgy0Ka0zLNv
frzvw9aLJUObEVE5jL6EjGUhOpVOQFfPPgVG2zeSve4eOZdb/rZ5H0vYwYmY1Mlr
aVhYx0OyjOh2jE9MaFmPiqluKbahgMWS8GzggqJc5Ap9dydNTmJtEuutepvNNUGH
ws9RoOrlOv/JleELEuNI5wNnnORrrKGimiTBCMqDRjFtYh1iXXYc3dmicWAsTT9d
BfYdK78/oW/CtYD5AXITPuDT/9HNHFmvh9yxC7l7ZqWiAJifdFhE6J59Xg8uvOPe
tV5AOotmtSJh0OLu/rNBySAdAhmSbmKH5LAh6O3dIVdHFM2JES/7Lla5sZhHr0Ws
DiAryPGupJ4To2tijwQWpvnINcpTZVtrWXWy1PJvvOKxlCGOPcolnRYcPHW2yQoX
9zd6jJIvfjuTaGi6YqeABGKZgCNnfQu2MiaqXOyF4RE45VY9/BjmUZA3HMzmbtn1
CUsOwfcrqmlgtDW55z+Qfn57Q1bfzFoD9rZOWxU97rhDg+yDXy/mPikCs+8C8pIv
GabRlZEp0WTZaX8f0Xdx3f2MDgcDP2pzOFj7nP1KUdzjC85z4EpRKwmG6/dM1KVS
w/TkdUfwbwF727HRR5vyH0utCFWsl171z2lpeoPTHv9mq7SQdJSVAfNWznawrIpj
EaZ0CSQXqFnvezdc/VIoaUkKgWlM71rFqmitHMQXe7/zYfBrNJm6FI51gWxwsdgu
2jKR1oMYbpCllb/R1Ne4Jxpy5ClS8p68D04msD3wuLPGqmeB+RrTouGGm0O912WC
3ErVoKkRtpMRQBnPVpcr+3lAE8es6W2L0xdSYwR1nE4i2rZQJF7d0VGsN0jC/S8P
Mwu2/FjeYyxCAytUQuN+0AGENm/b9eGWacv0nMQzhcDzYu7xHC5d7EobGS4DqvIk
tkTNApjpN92ZZOsNjjzE+ZLRWMiZCg5U0nij/R3DPO8NFfWDY8IUebl0Fw6peC27
h7Z5jrrxek2BfpXjkQ9Eil95KSp4wHrZy6sx11V+Ysxh4r3HJnzMxHJnI6qyPuNG
CgpY6W5L2kU27/j7sgWdu94ItiPX2oQQ4u10LUgD7j48VyDxG1MidLqb4Pst13GZ
5ucvn33KMeN68sfhkWwBK3XrVs9UV5lTN9JeSoZ91IOfkObcMs6lpEy6+B146BLh
yjWAClW8Skl2TM/BkmPeerghZHiPKoKJwOWZb2shRkfk1DCLSBaUrqju2ha71xKE
Lney7IvPapiIBbgPLU7Xvw7Uq69jS8+wrplg/J4A9rpJSNE8YrlYqtqgFRdT+HY+
Ucygv9rsSSsVfKB7fRqgyVfsIf+Y+vNvfgBFEynRIJhp8gnYj/QgNjPy/0RZ2mR3
BkMebP4dj6YGJ3FtY85qlZhpguLS+KVm45pEXm0pYY7eexh2q0vvA9+pG8S7PU4z
ryRYpLM+BGpzwfzSHUPqS/oK+OvftusJYRnp90j7xAul1pmnO3GPG9blYxlGF4cV
Y+YY+me4TouEZsktpQB9f3iHHA2kzneyRYv0rnPbqp0o6Y1+4Xz4ClPS89H5anDF
APtk3NdzaalqXcNjPsEAvpq1PoDV7sRyBKdB3wSfXx1hj3VkiowA41zJlSrm/Zo4
y90DsGSYjAXnKDtSwPOQi0i5IBvsy8cV94mbN5vrKsSvNebJRCSfYbxv/sKTFxZr
fQnkMigX1Pkau0YNOYSxlHEeDUuOiWNCMAeVglMKdOIXeBso6IxID7W7nRM3/Kej
4fFKjT3gc/KQzg4Z3DgJ72WF07R3xxSU7RWgEPc9wlR84zTFst2zunzMp1WlDahx
ZURgjaNXpQbH1VSV2tYsIo41AJGzsLrUY6usmq/vUNICiAJ2MSu4gO0MYUUvUOH0
YL22fO4syhyATJSlGBRDbZ9Cnc+PAZuVRz52nNwjQRDAnbE/xvSf7X3q3vNmT8t2
nUw0DiyRnuODzuirOJ4eplwZuDbz1SNVokTwL9loElb0yeFH4FL/HpHsLM9Vb/Dn
sEmV7VYMbcmsRERksfKnfV6wcA+dmE4HQHXaHJfClRlgH31UWh7N0cL0lD2FGtUF
6+gV4KVzAqUNbkvGmi6mkVqq7K5pY5v/9oagS90nYcTzb5xk3YBwqsR5O8xVyN8X
NsgGtK0yCo9Qu96d5TxoMyOr35+vLhVdL9nBHxod+eVPGKZNrtH+998HE2yESl4H
3KF2QNDrvoSDT9LiofBQxL6PBNWraB+Sa8X8Sr+oTQ9VquCR0VlQvTLnkoYov0QO
GeP+t6VPtrSkxFgA5ynWaKeKhviVJfpMAInzzRJNltQzIukA5Ej/436h1+xQQoE5
s4kCgKjM3YUjhp1wJ2FPrWbeY6cNDGd+wi/4DDiB59bbuZW7CDZIsNiFInW5/yQa
jc7sR2kTeLryczX53rQsrkRoWItnPOeWEGx8hmv6E2UYLk6y0eNmh8xmznmfgcE6
6Obq+0uBrPUP9yNSHTUmesGbPGarpaRo60qnHB3XZKGMHNYgaNYt4w3pexPHogJ0
WcdLJGoFry2C0vsIHgmdt0i1NVSlSVbOda5iE6OeoyrAcCi5xS7DML3S5VusGwds
EVsx6zOz4aMGm4VJis15IDxDJx8jD2q3trA5PV5qwLNfSVOwpInR6byxPLhdwKqo
iw9gtMd50R5pdRzQurweBWdZyZ5peIa69k+YU6qwL06EaQPVQJ65Lv9dGM7FhlN8
EsRxgM474bbhi9aKuME8ioRPSLYhKFEWeKtDu16ghKz5/1rCsg+MjGS1TpfBDVo4
ZRf4j77taCY1KwIZwtdhFTbuqgM86IxsODw1qP2kPD9NYXcYigFtBfugrell+zjO
2wUpyFgjnrO5HGPt6NA9lRwc5qrimGR7f1UcHClwh2kR2g7MmsUoyDm7Tp4UWKMY
PnSFyTVqmDJgLHdJjx/U7fqenv2ZfCY6t7lpwPUcMeAuwG5sVMj5TTL6+SBVQ+8a
GyAsK4GwQmPGykn8ENCAXA5zTPxiNjXCuFDgprSUpvtMT+rHSUS9HNBZKcf8dhsM
Xh2CYHAwt2XguyW8GO2FANNHA7OcItY40xqRfog8+fOL6dxHE4oYYaLZS7EiBSmR
44KS4HoJqNW7Uu5zTtJ05XYXB28l6fjY30cy4QhdLyoDeMtmFFRzGhD8OSNnInlY
1SIQGWag3KspWDJ0TWHn/HICFz5jzQTnTULQ637UwRrmMoBjalLD0BgXB/b0arfj
B2d+NX3TNRVplSVpVvLK2Hjy6qgjhzboz/vpHtwKWDpiSHv/zLLtiXqurRfybUSc
2G8ePzOsraEbGGl1B8R6b57LCtdA2ilZTnDPMk/MRgArOHUMX0DyiJ4X3voVoO3i
kLw7FZggDGfpMVay2coqf2rW/BEsdJ8VVFBJ0vX1MB0SAGupiGcPr5QOJeWHiXcz
tuVpNuKk5A6uE5NY7XGdz2zMGumb0wHQW2iib8fEwm7Co//ZP9b+QijhmCbiekNh
oZrJgQo4+vjkX1lYWyTVrnSI068ZzYugDHfdA572je9tqpd2PzzO2O5qsHofcriH
sAnpvpYkQMHEpmCS4bOD8oDbLz8i/Mb39c5NyIpM2jR+5mg3D/OoYdYJOhvqZzgA
3i2h+ROaK8wt9WtC467ySnmVyN8DTA0zgXhtdxq2GqCX9KFu768WHYgfR0P1lZne
k/AGGBpDfxD77v/uvulFXwwomPhQoJWHy328SjQkSpZrWfPL5/SnUtOuwrYokGPK
dFCiGXHbe0D7UhJkUTjAt4M46WwIYiplG2FymJ8T53spjjQMHy3lKwkWq4tl4se4
UIQ9MQXYX1jg4avJZ91h2RNONfEPk1NgrGZ+zvO1ZWbrz2tDtB9f1mDFYPpgXgLQ
H495skmCSkPFipYDJbShBxBzd8Oo1c8irtBLVwV4SAHLAV8eJDCIiSXdjGRn6itc
ogSs5ccXsBEYsFWjZlama7g/FFX/wHKV75hExBmxZzpG9ah2eUoz7Aex172mig1R
gPQrmc7B4DFx9N/hVxEZOVEIZnAQ5FbPLQIi69pELfZXnMnsN2rg+t2TXGogwPNr
9tayiC8l87TlkLlPOCfIZ0amr0xHvPAk7pJqI0hwcI0mywsfxAs6WzUuF/+O6/tu
pDtMGaq/IrDwYXfX+On0H5qLw0fnSbh7Z0uUBrGXWQ/Hc7nYWImjHVkdrhlZpsPc
PZIhIH4ycCDZHqxOGTX8V/dDesgCpAP8MKsv3MZ3AawdG+Gw7wNmE6wZaDOyCMGz
O9bAaAe/is36bQXqoSpH5rlEsY61LN84z1fBpSNSCHCUiEd7YrZnaKaZnw2jyNTG
rqHjnURLKN6G2nZQU7D0t1oCSNhUeVvuAn3MpbrM9nMLphtKosEQuchcgtaxjU77
wOkGM51rJRMy1O1xw35eDzfpSGYiIgks+ckiWg8S983ufu9ZkCeAEiPnCQ6yf0C2
BuOpAucJ+7v5tMJOInPQ3JjpFCoNNp5EDD10tSPRXyph1CEdFHZTsNSWox4CPq8a
2v8xWnD1yh2t0Xm5f9gYF0UFGhvnXq6vET1X5aY7PSKwH5l5C8i1uKirWb6QNe7L
NOYLTaXbR2C6UbK3apnm934Px+/lnR2n21wq8vtrPDhdAPwHmlctCopvXPxfnHC3
/kk+Q9FgP1qG7dtO4RjKyPgzpvDVc3aUpNkTGGiWRlvSDHyW0OgGD0aaGDnNvjvB
1oCB8nkVX6VXhYmc+1JRepPSxoMLXQQMLkr4cDSZ2/A4H/aYwslflYb1EBupPNq/
Mu9aeWbkCyZoMoWAW1ahfQm4w8f1PZmByKGLjJb+BRLyKrbwXg5MnAw8bbeYLFcJ
nfpgGP3wpZ3WztQT6zxxA3E7sK/RMMZJvy0ZLQnyNMB0hKfk4F3LZHQSesHT5obG
MnWiaGAi462qrvyVfLxDex+kwZBWX4vRhORpvn+o8Jgj9nvOI8QL57nO9sgfRDDx
EpASCp1IvYosGwiGHxC+XkRRXXFOcfuFH0w3fM31k5Qqcg/KAtUFkyxhApK+3rNI
bSS208lZE2oiD0gcdUL1YGbHzc4F7mzvxNscLWTJF5ieEkT4RWhiLdFZqIPwzbYs
gT26zLO/tYxGsP8DfcaoJcpad72f/+NSu1dcE5zOwH3wV0OFiVYbIcIF/yjsZKS2
Ptfntg5N93wBORzAg2CxwgVcTx0Pat5VsqKa6kkXPHDV8Gyng4959/fdLcYqFwfT
LJnnTB8ujl3Sfb7Qu20uLiJaSBxaBOYpuI1TNYxiAkcc0CW5nA6hMeRk7GkIligB
KniA3wfPnb/3OiLFPfbgOlZfzWJO4tx7O5bZUzVlpqvvfeAlLoiON5uwgyTp1rAm
R/0u+dywDG0E1h2BsE32NMzGMb7PVdDVsvB/HZMm+tYHMjl+ytsgDYlWth5BoI6t
r8jlPXon83SQcCwnSAgDnk0rIesWEAB5T3oztEX5E0li3g9SxSbt3KaEi7uoI35W
8eL6QitQEq3oYw8pI1V4B57AIR9fqyjoVAyh1oRuNXSfS6yvkFNiRyvBDT+d+EZL
dtXDBUYkeGV2d5DS3zKEDgoqHtloS52s5toCgl3iMurwocoqqlnAJ3+z6x2WMHts
NgkSj5H7Dno7bnOklwEkQ8rAQGMN2536dbXcMR8TbBOnXodDi5imcHQAlbSn6SUi
ZjDQwVDWIJhwmrRQ0nG0l+i6p1L9BGEo5FUZT+0eGQvVXOMwd9Icw6aAyI51MKwt
QZ4FLiGIyoILWczDO3c1l7diLonQqMcIac5gy2e0xF2Lmn3rahH5DqFZuWNa1S5h
hNXSIHsPx9TvIZKe2LIuR9ccxd7UDSsRjEleFYa3h0kFjkCDLPaSz4ZfurzyGcup
gZ5IBUE+nHGS7T1eqKv0/EJ+NN9CJYNeDNRL4R187+0kLD26bdJm+29m+9heLNnV
yN9Ac5bhzAOTO1LBwnMB23TSKNxTgecaMsR5bLwCnd3BvTjMkGjyhNPwwctXzJy7
vvMwTlVo92+5h9qWdgO0Ty8dUYmlgk3IkK0esh52aKBans00+71sDVkoYIcgElir
kWIM/6bLYCpfImglWhqH/tl9JINRO12jYAvrWjBqyYWPlo+rv23FVIpy0jPSuIiQ
3LjAtI2CTiay5QDIINj/5ax6mQReaXtJEEFSrMAKA1ANDghwUAGMEnaoo+H1TA7R
mXOD9EQXau7B/jE38ku1MyLlTGTHe1F4+MNAUyaIZV3CtlQxV2ROjjLKsYTX26p/
MfDdSzXEziVMO5hJfHYCalpftcH56xsvvk9DtdAPGuLUR3aOrXr3zubbdZh4NecI
GDfeMq1cWH8qNyETH2jxlTHS2K4Y8qiWfbVsUZL1ncTPzlzBiGjW2FoH+PdYfJtw
ROJzr/Yaztsrq+uvyA0P+edFT0kmD8dL1SWR56rDo9MIY7KmyXH17wap4XlWkcmi
qLUO7EGKuI8Md9OqENevAMJozdRdruRcFlOHpaGbMbO22joIP2rx1mYmgBaOPVym
VFtPQ2dwzEAPTuAvvyNcdmXZs6VjMunxEUmBkFg/fuZ8kN8NGV53+3P+P3kbrS6o
K3GWMDumQIjMOU4Q2hcswXUqtH3P5taPrfVn2Bry04TcG2ddtrM1zJZBoOzu8Bql
Ykv5eb6FkehOvAle9zHNqucSLtd5FD5qlbPIl3/UY7XOHm6/rwmo0DbPwSG2e+Tc
PL1gEwrGa/G+Zbx+GibHs5OXsq0bEDxBF7ugKMCw8+frADPvhUT37Rk4Qz4KDKrM
pYcFBE2Fn+NdB602Dy1o8u8rjb2c0i4MR8EmYLHPHFAKVkpE9kCC9UxTsLg1a7Oi
36hh/kE5/wZc1Tk3lAXc36AtEOdnK/GQalGFw6ZYoBxiuq7O7QtKCrB60mw10JrL
bJnpo0a/8TvUO1rD847lFHS/ul9IT0ZsIJtXd6ZNAofgUcgoZjzsi2NThCMzr097
GZ38CEu+dLp7cGPeym8kXqvzbki6YFM/e4Hhu3GU7pfMvosZBTUcOf5wvuBLmCkl
26c0S9R8OcYtZkTzTd8y6RKJIFqKQ8AQY64KDaqL6gnR1zcSQs6jUbnZSKxDYZ6f
Zq/YlR68V13/1EgFGxNX8W5Ih/WdEOpzl5KZmKH2MpxVFfUc9WKnk08DsXsWnCGO
r3XI2unhnZlt9WFhuUoopaNRxze/KTT+kP4QhPGClivYFiLYYOFJGI66yv4scZuB
nDBfpT55yig7HCBMsOCbu6/fmrgQlgEnLQN8MNzAyikdQx1xBf4Ozt0oHUbuKZ47
/RHSIeQe6i2TfOvIUmlXhOYuUPi0TrUwwAwHQdrNoW9H6KGsOAUzNbDRdHq2CSZN
msTSUadxLtw7eL4oNNgftdC6OnRlG+PYgFRRH+0NUqiSpYFYAF5PZSmi/plA5uB1
2rbWzwtDrlrHhgQqdgVNMmGnj0CiikFz3dspE4GwePuYZNKE7Qwz2Z4NxEtIazo/
ktJvoC6kWHViB5eiEp1NErVl0xWxL11Qc8D8nL0YuRTedb/jCoP6fHP6xXz2L8cS
qcML1GaIpJuyFCbYKURqMjOAmDjigSU/9U7HUYWZ9W/FNGEkw8ogxWmhzgsXfS5N
F1ieYYMbwfSDLNb+LsDyffc2mOYOFhYyzupKH3bJCjW4O93ZHaaXQlOzG9RJlPgH
/QAeRv6jdk7HpA0PtdDzy8IXlE+c1M1F6OTFd6nUoV+SaUns694TKzQzhmjDtlLl
f1vZvyL15qa/QoWVT21a2HhZ19cbMDznJm6sM6aZ6qpc1xiMkUJaWP/I+uDGMq48
vRkEz4deZUvstWcFFvraeDkkbDRVPiad+BlHACWV7eltaCs+/BzpB7fr7rculYl+
tfnVFX4xGv9ylHKSPX03jMCjkVAyI4V+8OBpak0GZhkWiIFhxrgUrCnczuw640vu
GdyLkuBITjdq1y8D+DALimh/7gku84T/fbueIfBsvI2x6OV+7LxXMEh1I5UYeRoX
e4xGsgqk7nwG8rRevFzfYVDdixMpjiMLz2goqXnitwETB7rJljUlvzqDWN7QgKxS
OUcVNilKGft33jeawo3x5WL+RQd+CfljCR4x2pqAckAXerNCP/LATQUEKynbm96P
aLZHqxvGueJmIO2ToDTGspR1s/e0bMEMmHWeJY0lg5jHtWbXnsygmv+x3a3K/YZl
dxPHOh9xBaGHfh+sWggu0zlADtA8f0t36vh0ivhZSszesflzAFtMEZHUQj0TaCbL
LLDNkShV1BVe4kiCuarHOA/zbo5JLqprEFd/75N926GVie+/OPmJEzZaBxOUmAv5
BmDbx80ulvEv5V7sdoVH2QYhx+6RCgCRxPjYDVBOsHyhGuX95zl0lNusJ0Y+koyl
cHkifYV3grK3TSVxfEmRy8Z6NTGtmaEWvqf6En5FAPojAzvlIKi+HRTLWw4vyN7Q
FCAT8UsNJpntWTQI7+18sqr24k2IAUsi/B9mTnDALQv8W1J3JA0Iaj82WvMbmmMw
g6IWtzdc9DeCfp31IrN+lVH8s/r87Y72PjbHryyobOxcOrtvw7cKXsFR/Q3obQja
El6WU4ZkfnHgodKuk+KK1/jdBW7JSqArWmbY6d0RqLs/zX7RFpwQNu/zp8zY9EUs
CRE0sC9/Oe63L8/Cq5HV52nhKh6RHjKH3jxCgp5O/ThQ8ew9HBMHHW+/+M/0Mzui
s87NCDQ5PlW09I4oc0Dq8N3VTZgKdyZipv7Aea1rpkwkbpDyNcgvxUskahvov7cd
xe8HM0ogW7vHuKcCpMhvMmAs87DGNFrYLw0y3WmNxVdgCp3EDMVEZR6KjAGB0xaG
AotPo0aNrNzUezHMBWwe9hLSE/Nk8B/UUb28iwVDwen09MkSmYElNm+1+zkLH80A
w9CE27F4Ek8xKr/HeeyuKHutkE33Iyjbx43rsvZTSL/2wckBAwY7bu8YR/R0Hn+V
Y47jjdPKqKDRJ9F9CFpVKwSDaZaJ42fq7Dj76l+94nnIzRo8/iuHsUk8A/5r8qQR
096YhoU+/q4+uvK49zwU0WY4lxs7ef1wF9d3vK6OqoNAFlwpiGPQxlMg1+JrBXTl
J4SRUiwilrYfWTid9TDieNHSjRwgMuLZ5AJYHIRZ2XkwxmCgH4Q6HzaeEO1zCAPt
vt/3Sz+rHwrYM59+eE2NYS4bzIT61csoV/iUEw/Y419Lp3VUxNHvJ6wxQkMWvbM4
AHmUBDbt/rV1oaUewhCcy+Xr9f5+NNwzB+vQlJ5pMT8Wpl58MX0zX7zxzhX2tyqm
VYAkOZmRlcr2hL9jJepdObk+zAUkT77EBBlQ/flpKiLisP2eM94KrB6Dz36nTfjQ
f8DdknK+DidKT0mTlYnHHTvSZH/qKLBvMP8N+m67oTdDJ+Xya99d1/Sfc8dJZ4Q6
z3nAQAMuEcz2SmmUxuHbgwIAyzN79/U3dwY3+CpZlNAbLleHyACDS0hDtJj0iWNm
QSCgBrLHgt1Y/xYlIEysMwI/QA2OCvDNu7Hic60SW2KjUPyVMzom0zJb9Hv7fdlK
BpOESs7GQBL4VHmkTGPbsJAOQ48qmtGNG/vaWwAVOkyhin/BR6+bv1OI/QG7RoGP
TV6GKTZ2vGPDmW9EdrE8szx6dXXprVWgiK+/xh2gupSvxytz2s/cZJDaqr5BtzXM
Ca6xD1XhOxYNql8HeIFS1hPtpRt9u8nSjfC7cyYu10Q1RGMNRa7iISHNCqlARod6
zsPc+Nzsui0YxakxjP3jdr/CXt87cw+JlaRwFp0jbp09MKqNONgalbvIm3Eaoyv+
VIGk51crDPHGiz0jLRn9ZO7qiaegs7EWKlqSvPYgyv+SVZrleHf/98c9Um1zG8NH
Oku5ObDmIZbxBgHoab3xNSvtN1p0bvElEdq/7GFZiJPW5iFtycQN1jfWM9JINc63
N50VZb3ScBrG8LKpEqHDTLm/QUUHIAdeZfeUYIZiIecaapuCmBGUMZ1I6hUG8sHO
Lj078hPJhyoFTo9jD5k62fNDXiZ1Qbk11yWM3C+/jImB+gcJYEcA7eA+X3hAM9xw
Tv1I+Iaqt3K/4U6XavCFJk9XGPREENdlqOXHRHhxb2gefC1tnHxQr5bM+UWdDbd+
K/Y4YksA4xzaeamC5whD0A4ROJnWraBWnGRBoKVjwt+v5BLCt/7gtkAvysuzNzps
cyAOrmFm0h09ng34emV8F8GyF1Vgfp92NxOVVhLZjLrzFYNWZoQGQ3yFgqKtY3Ru
inD22GJFtyupea4+EGm6sfXUMHldQRY6OAEAmWPFTaIACdtSLJgC8J+ZgprEePuV
s27rzl558XV/uC9Wz5WakX1ErFHmakKgOMqUUWckW4lkT9lwEF0S0MtFq+etmZYa
C11ze5YIp3VNUIt3YCWih1cB66HYkPX7XkOD0ZNbYjQxJZ1OewycCbI8b4KwsW2n
xiNgQs1i76DSdexPAph9vFjy99ztIPv7kNaqtCYVlWGlBu2rL/qRluJHIRxA0WL2
0Zj8AuYhgvpwg8ju563Jj7MMue7j6oIWBOM5GRSxLGXavrCK5bDH5Z58Ea3WLkyS
CIC4eyTtQs+Rl+7xrp46lrgKHpm6SthDMa+z2q/ITd1p0vnOmOM4xu9ONJ+5wQNO
kEtXCoPiyHyarnny/q4RQh0Rb65tQc6pAiqW3gflWjuWAuYIEM71LjY9czIhjAB5
i/hbJX6nhMKhTacRzyoPn5EI7VXeJtWMGO6cSBlRqS/9uMaTW9QAHjwWcqQWuIED
Wb0YreM9k1Qyqna1KWSPkIedizoRF4smP6FvMh1Ie+S4Xd2RYrOBFhetEFtCtbVu
pZPwAxazt4dkX9HnJsYzFHGWRtlPkEgj/S231Sz93hQhOF5jlCnRHqFIPwn81nxR
eskVRbHCR9KaqsmHs5Qqw0p+IKP6S50eNj/+vNJpdW4YV8UlWLavn2iyUClVlDiZ
S0gKRg4Oa6rpziy8Rdy5wJ6Iwg2klyg7nqCFmUUaDoYRo3xRs1+h/+8bZScR5+JE
5xsv/0RNzjYfbXH8N0kJdQ5hzvPw2SKHyGB+aLjH73vI+EKpnhj2/pg8ZCdMbKBk
lMeOXU7zLBUVoXAhKwKkFN1Uy5Fyc6QXeIMHewMUveA9n6WLfk2AMjqzhPnSwUJR
utenfusjii179EtXl26t9Q9ggaq2WdYc6VVl3FLSnRQFHlgG41dRMx5MUtPnpvxe
8Kr/QMreVCBYmAKoq3b8TUT4Px/mr+qCoLKuIDIawoqjvcRikcr4DtIVqE8H0gCx
IyoQn1skQDHxlHApYkDTfNwzqpOYC/w5knKUFuKItQeZlVd7IC6HsN0TYq2gWbCH
6pYeBtMklu9mDQBMB34jDXY2XFzGemdd29cW0nN5CemH2XBbYdLIMPtf+RIt3ue0
nx/qgBPxXR2niza9D58/PIGEeaqczJwe9wRIuz5WpQJXMswJ9XxFcaMxx4n6f0Kk
SFp0KDHVV52FgpUs3aBxrnve0L6a5QFceUm3UdTKiIzWjUH47R5Mld4jGOVSuZlo
qgm/DEel2HfrgvCM6HoA9k5bJcM6BOL8Hv4Zo3VFSYEsF2dGZ464K+3FrnT0hINv
noKZF8FDLClUboNp5ez12KYxum+oLB1PcszoAqWzZBIiCyUpdTiHs/luYlRolTn1
2mERjE6GLr/L+q/RQ4hO/WJe22EPtGTlEQn2OfY+4PsMBTvvA5re7H1qleFA1VZa
av+ItBf+tWchVO9ZKWSCjt3JvpcAImT7wu7ybSlxFMcK7edFiPreo/j7tejRrC6H
86WUo15ikTIVMS9QeC+ZH6NgxdfULThLfPRepuGDwpxqNVbUUxE+FT0nol073BP6
TF5+SZh0v9CjgvOynP9/K1LlY22Yn3XVFeFaN6xfzIjkBd3i7oF3wrOcDu0pY+Ar
ykfBRYZ4qprIW39ek9Bi53eHUIM04jIMh2M6/+KKwU1AZlKyOacFlbafxL+pWCaY
SuHBfduJVrjM5/zmo+FBFUHaickFKFOzb0edFtjD/1rhouLSCXlxSy+pm6EA7m1H
2Y21WbjlWcp9vqgsG8FzoAFaJF0x5AfvY5l9soIHe55OjgmgEFSsi7HVvzzQQjcX
hVY+MSFNx+PNnWPq66UuW8CPW/yJJkCfe32B1+JFaZn4hcjsff3zM46eb9GO1FRa
UMUdtzGII4G+0O9qNs4k9X7D+570bdh+inveJOFKh9L6BkBfxMA3gWD4KLAZcx7V
1MGeHumkO9zWRYsu2LmixSVxQRK1W5+hr0JwYXrjHCzrJcXE0YrXG7zSGNSJohZL
Hv+1DSJHiy7nkzqzx6Fa7qCsaQvVIK7HtXV82DF9TPdk2TxvDH5PiAWG6Yny76Oo
xLO3EcR7Kjo9rb1nDkUL64fWpz+kd9OPinWRpGqpeKn+SL1u0CJbmobHWfXb35Kk
emvM9GstZa6uBfYWCg4C4ZSpeKRI+8R98VPrIQ+NcW7dU2snZpQHKQDyWtP1I75D
nt6Tox0JrwamhAylmeEVOFnBwDUhh7dXlwkzymeQFlVa3rF8IRSQHYMXflCQhjQ4
KtwJPhfCEJY+PrzOHbNvuiyJTtGWFTlug0fd0ij/CRAnw9/rPxYWU2ZSLgExuQj1
exyux2dTl9VbxLEOo3/ZTDR5UiG/EpeEB2O0NkCAOyyMRCAWmgjGaioAIHBvcNLK
hHiNTL1I5kktiukSxZt+f7G166zwWLoMNddYDdBNjPmfx+G1+LXVIJULLidAYWtJ
mKUW671EfetGZ2+Z5nSHX7VuPl9GOh3mD6KeI5XNCyIsyJ85ZNGQTTHt3M4oPmKl
kR1+WfYm2f172Y8+8TJltZGETGBkdSdB+TgnHisJYkw/BPgPvIuRATXDTOtphgrF
LudaO3HsGp6e9smptGHnn9jInwHdg26yE5ro7oJprq7ebSV+yWGbYG/TJXCANj29
IJGBozQCfEwGUd4mqoYGGsVAwSXFTHhU6mgVdHv1MClrJ7/Yww20F9921h7NEQ8X
xv7LlvcuzHQa4aeL2zAU7whk3D7KA7/d7xo0bTi5fLIyAvUzXds7uBsbgyaUxHPm
O5W+TCXx+EdYk1KNsKatXLG01icTbSIomTb88DHvO2rFhQUC/P8dWy0lajiD6rNp
+CnruN8Bv5ycJixWO8ySlaOUOE5ciu/CHcRJR5JYEAhDWETjvmM+xoIdk7vp5tfP
QugAyyt5ggZ878A/Goa0AXRHQZmmT3BNqPiKp254efCYpm9obnCjw41LLc5wBC87
0fwmkKGV8+ZFWhZaII0PknrfL3bKseIzXxQzEAcZXymaxp0GMIMIgyziC5lYYcP1
/8CVP6E9jNgyMWrucvU7C4zWMT57Ligr1BVKRG3oilhpLi7FoL+//lIZ6W8BTdfT
Niktgdko2d5WRdijRXJ+iS1FJDv4xb+6ODuLXJuatxvt34yFY/3Y0u4p8BziSrnS
5H/nmSWBNESHGCzwXCUWwM/g/dGTAD6KlpwER/xBE7KKkIKVvV4BqF3u7Gx2bN3i
rcLZ2Fr4qWFb3F5IUL1wmEEJTPFMLs5xyJ+FCQFjYHvHRCD0YlF0VLBvODfK85Ln
/dO3lTB2T4HHtZy9tNJ4u6XLLyvkTtvHP5QSCTe75jHbmd2Z4EBKm+2qHlUS1DCY
7xmRsf2tSQmBixjngo6jpqmlU4HwY0XBqROPg58e4kvqSxfh1lTq3ky3VfLpw2+W
y+ROBy+21JsdXg2Y3Q7+eq24IggQWa0BHS5c2/KHfIqlqfQKbfETFu/0jQi4TUGL
88qoCT45S6/W91KwfiQ7o7PKoXgM03xoeYT4XZeXXUQPzt9O0io2Sw0JfKHKQT1Z
sVLGQZwlOGKsrS3dSwitxDR9ff3pLdlcaGpzlV94QUHwvFtunn4VLsar02+KTsUY
+3NJopxaK6gJwXsbOFFqfaVeT1VNBKk7l0ipdyaTh+sY2fZrshlPac9X5k45srvq
UlpZrSaijeYjvhgDyvh+yMTA7gmCdFvriIRIfTKin9uxozNEdtlwoCbmExGZovsg
8ujnPc6bQ/Bk4xd8U19y7oleWzbmrTX/2Zn7pwYsNkqFn03TCQ/MfcSP9qQbnzhr
s3mmpC/uBXnfcpZF0VaYv5xA1/aoAUPtAZ+KgGPKJAnfzftwtZLZgsl24+UjSySV
l5ZHwK4iTO93dI/jxEaoL0ieDECt543uIV+AhMw8T9ipl4/OliPYPAjZXWY1Kvb1
jE53N7MySSibXCQVxYiJucPzo0K1XzZD5W2f8sDkFx7TvOLEyWHThFzVCsp4UcKh
pu+oNMstJLT0goG0Ku4afvszMhw5EvnYyG24RKqBAz5+njJNOyQW5fKugqDO2TCy
TXOxClNtwTQtq301qxwQfRhziETAL4FcdH3QN0O0UpIGUWke9IPxnhltoWeqW0fZ
8Hlcj3jDf2vjB7hNOWglVZUxn6eQukbTdgwO31PhlfKHUZkndSoZbB2YtQGWT4y+
k+D7HswInL0n66pWYHPpDq1Pi51YECjE8kgXOLngTq7AAoBCatNN3XAl7Ir5ctDK
Tv2zH7FnHOPPPLO+DSuSU9T2+X2Ub/OOwu292Jlcoqdr5v87GGg9Un2c6m+x6xX8
yGALEmxK/yF8WObTsYHyQKLJHfEsFkkj6FDDl4ecUz/qpJSv51TzqDflVODSRm6D
zroWe5qDa31GH59LgDp0q5XQ+UL1WpFH9LH4oPqmHKMm181Qjyq4MZqN5nheu7E7
y3c4noat3ehyI4cVKjtMjIg/0A5oV0oBKGwEWyFQ/zcqbDD6hWnHtjf6hfFQiSkO
ejfICs1pby04mQgXrgfN/DZB9eUCTK6NS3wkJhUaJTaRgukLjURhq+szdEN3R30F
kuBG/VxN3ufgzop/tKn4jlKyNbfmG/8M2o7Lr7Xe8RbLH0/tYNHXXinuc5+yYNLx
sre77G/7E+fNUsEbUyBGwimreEgh3FAVqRlKDDPfMOkaKByr+5D0MaH7mz7xkm+u
ecY6OSOJAoVb4ZcAm29tiMXOP+Y6dnhakClOvTGCJXjJ28U2ZsVMNGm5+3EShbR2
e2hCJO/IshN+I8JOQUNGqytNQ0eHrlWVsQyDS/B1T0Km5Tduhp9FchC+3W/6vOiv
memNdQakyU2w790Go238dW4Rd5z/LSVPZaG/IOPkGJukOTQseqCdHf2IdUowTpOJ
c46j+jQUYoGyiNt/HD9YPdZSZPkkr9tphfc2mtz/RCbx+CctauZexQ2eJLRoI8oa
rhazTen1F+NC+d/xdsU6bmjr0lqNrHh7bcXrS5D0qkelHea+Y8Zv7Zw4lbByeKHQ
Sop+8rxrS0G6FcJ51nSL5RHV5SLAc8L2HflDMfghTRlu1/Wj5BpxBSRPVy3x6FQe
A0xv8HwzRMytKhFcw/dJ9m8HdvjMxXkpz9Tppw0+/q2wm5nGmoqijhBPqo3sp/Yu
0g+VpgnhxiX47JicGriIUHqflcQgJOJpPf26prQJapo0l12+lz8Z1IY8OnDAVzRa
c+MCSz7CoyLvZ5Q/Enoios6At4kCKmgvS6fggE4iqhZb/9IFGJl0NrXPq1jGxVR1
glm9LXrvoAneOozE03DnuAdK8ssMg9oJEwVWKG9XObwuzooA7dCWRwo0VZUPq6YI
0lA+zdVdNcBfvjJ/HO5nk8unuqmsgp/qX0MY/qqOIbSNeP7Ok7DMuKf6C0v7kBfv
Lvk7jolQNP0eFQKS0ymOP/Bch55VLhIFAdZfI39SQQfnoE5H7sWEwpIAXfbjyBY8
lnqyLD403xoLDURSRbaVZVmJxAyEbS9dmA379ZJ9VzR7hlORONRHJrUpJBiPH/s8
CsPdRjryS4iQmtzNs1wPV1mYk3FYu6Q2I89ltPsUDjc/zUYgk1hbWSRiTDqM1TL9
Hdjj/PztFgZkjoZsJdV7TmmzFUmn5EhsTsNfu7busJiGLkV13miEpQqXBunYc9sT
a7x/zdpncIJLNYYDqSsV2YD3VoiFfjhP1PrxZmI/GUMTiu6xG0kwpJ5Danvt3/pV
HqZ54RaKBS61M9EmfYwvDyd7h6g2axs+MtAAQjACh89PGc/rz9HBR0w6v5FHrzXs
Bc0F+Gb9hVpoAqczQUsEK8Kdfr5otuz4Xj6JWJ90EXcSzgiFOXStnZDwmq1L+VwI
OrHmw0bZovtbla2UChORtWfAh+imuBsTd7kr7kA+xWFmjcVjJ9UTJAMCA+I0aPJZ
sMhLat0RBRyGC1cvHyyjy8InJ8H4DWQ6805Bbf2Bt02cbHfgjRhlskB+rsl022+c
yUYRuKXswbL+4klONNzXppwW5jZzPhet5fLhztVOicnJymMgdiNNTblOVdxk+cbZ
fsCVws4I8iu/IqC6tt+Ofmv/MkTSnNBBjWzeNWikVaq7ZL+K3cerSEhzH74lIMBB
BMwRstz7q02omHYq4ZKiSyxDVr4z9RC2cb0Y04+SGySENsIoM9e/Mk3Bgi5duwuJ
2ZDPOmVzrvJeXzwRyQc05XEIfTvm2mxAoS5QlE7TONshvI0MKunVtxWVAf+xVTMH
X4snTUjW5QFwzbKxj7kQBwyQCKgRG+Y9SZpHct3zpwQwYbaVCRGXqjb0uL7DxIyd
DwjV13wRNckEWGze084FYanpjm90qhDLIFjos/AdbFFaoPyS9/RWWTSlWjrGXPwY
h/IByvGMCAo/OPVzLojBPfrvYgRbaVZaWyIb4YaDSMOHkPA+Ya6g+Y2Alw60ZRkG
Ua2o5jR8C/Nm6UR1yahJ9/lHpTQIoprLKcyoRRGblli+/ZWQDcW4t33/AlFeVoHi
SqL+8ryLsTeJ0hyfsGKClVqXwV3vMJwBBj/eIdsUD5T5p84Bzw86Prq4sS5nI1rf
/A6jeN1lJfzhm+p9H/WTzgGhzOFSWVrBucyPjBItyMSthT8awfpH6FWQq4E7ougC
HveO9IxoppSMdhCI3SUkGlUk4fGuLdwZPIgpm0OCJHsy7PkEN3bmSM7wLxIZDVdw
w9sqL4CxW97WeT0P2qCZAywOnv6aBgI+QNBUxJazfMPs7KBF56lcBRSvBONcILCS
/4mSskiG5MDhWYJGu7ATnZ0eejsz/2cEa06DDyp0fI68HNk0zJGiIEkovEA/TZgJ
rFPdMogTUdpnjnzwXv43f+J6eTrLg1D/CW5ZoXC1sUT0ZkoW8eSafWj0w7MKdfeJ
UchyHibud5Ymto5zMaTqgjwAk6Yh21Qdev4FhbWsHXrEN7cCfAckkSbpyBASbSaE
oo3hC7PoSJSu0gIKMUux4NfoAXP70iCuB1anSn+CN4qdfQq2FzKitkgliMhU5ZdA
kCrGlB51kmRCK+4k6l3iM1b+dYo4f/5woQDjpCD0WSF/+8G4bE1xupkN1kl9gi55
xu5EXyHPW/1436QVmuX7O0jJhVSk0GNZGS0ZJZOi6xSNUd8fAJfz8IJ/7+HNgaSv
jb19laaMjzHpY385eV4RuMubNfwXwvGgC7Calukz9lBfMlEXAEw8wcnAtUEGWth9
t0ClUVFx7XIi8mUEtrbePgv+qeYxcd2l6fWOd4LPepkNsFnms/rOO8TuufK2qD/+
9r4PNVR2LhYZBS9K1194Sa2Mn+idsbhPrjIGV4MOBtbuf07+pTqdSfQJycQjErKW
KhIt6I4ywiHk74COUZiI5ZotgxNkjLR8dokWbQaV6K97jZ7T13xEnm0vR0b0PIh7
ROtoh6iKZVZ8zqw97KimVNZamFuKWChij2KNXw3VimEdSEH4omkmrhztjLi7owCt
mOHM4QffcBDwzx1u8+vvBFLIVj3pIXRnUB0YDNIf0m5lKAhNHS+9gyyP0QcLi9o0
Mjy/vBNUHsyHtwx5DQsyEd8X0R1x6oSpA6WHYe5XhCBrbot9CTfgRbGsVyaJFP32
dF/3vq6UrHq0K4wE+IYVTPpU0H4zeD0eEGfJstMLEq7h9HMIv8xhswFiMhU4fjYr
sZzcWWVUKfqOKk+/TwTK1AGm7Nyn2WbbXZal3KUUfywbU+iyZr8aqvs2229qbRv7
ZnEjT6qzwKe+tFaHA5D+KhmPBUYnuGCarqdzO3dk/o3jKpknEd/F5szZwVl28xqd
ClozBMPGhgAfH0+iNVQtpgIerNhfVSbHLXGIId1TsvKaT4i1JRnk5Du57eZn9Q38
BtxoAi4qDLAuYLkxKkMPYua69ph+HCUGZ4so41BM8iCNZ3xow4okfhZ3vzAHErIj
vgw46YZntU3MAxTEveVilCyOjk2vHPith8jrT6+2m8HV9ou08sPUrSUOxE46SvwB
kHu+pbdeNauuvYCLi2peE8KXGyIIIih762IgjSxnQ5+OXoSzsAu92LqkVSCq8/ju
BLx+pMkTGQtL1H+2d47KtPMlJzreGlfwbrz1Ixw3Ou4aAuQUGEqUWb/iJndmOMb6
Dkpgu0W59xxPtHc07AeULQwPJenupWkElLOFca/HRj3VLF5gCsAw7lvhySNeMs3w
4E4M57solbmNgzRFfzzT06zNGgPAVqLW0/tb6NqezIi/bc0Nae9UIbNuuneLizdt
YFsHIbOtgt1dDXLHNY/ibORVx9gXzlYBBDJGjja+r60/iTw0o+PCwaBetQHcauXK
T6rcU4jKsVWlnniKsy7wZzl+reRwpl/tVWfTD/lcrfeUqW4G8y0dBsykx0W2B/BV
FxnYNrgWOaiupOGdNB7v3qJBT4SMXnTWupSNiH/XTfrDGvb7jEFSQYgzAgh2Q4+u
pa+/JbW/sDzWguGRul7nrQbRKx79iVN8IJ//g65sETcEZyuipm86bzFngvRqcbHD
zJN6cozKvcS53/txAJ5CZAo3SMxWzVEmiwgtvciouWX4ZGik4PkdHstBMr2ASxyl
o2jmKwlcAJxOm7Q5iTaO5U95ypACLhc3D8U145lIV2p35FgzJG8+w+zxIA6zgNpk
3rY0i7jnG+PcnAdfXUb4WEsbJ/gySpen4TyntyNuS0vfyxZhWz3QkLO95OhO4AIl
/+d+0uiwnzBfgUFxBiMuA9W0cpWVQBrFoKkZdapUVhNR6uyRN/707NZAHTP+keDl
OfcULyfa6Mvi+cNsmVUWPLGDa2orUNnwkr+/UTHy5EdRJPc0Q1Vp99VI+d/9s+D1
CWxHJoy4Jt1hmMAmxdDEHg8uV+K+y/c26NtxhDgK/iGKxHEwxIY9n35CU0g/ItI9
VnqhBouIH4LQ4NQ6GhGQmnD3QHxiVq0s9gXX850PFIGHVxs+vTiWKPzyH33MRv5C
Fl1cHd3TgGW1dmQSaEqt/zY/Oq1yXYq/bhM12ijWrzeK4nEki9ekHSAa3cpl+yMY
or9/fHF/0F/3J1bAoeu5PRAH9VxObdea5zOZZjCURQIl/842AqHHW3oc7M89WibI
zykcqr2KsUo/ArLfNGXoDJ8ImWSMGtHlez5Jzf6d6+Kix3U7Zuo3XgOsKEQNY5Tv
uBpIVyLf3qPFb8/gThVDFjtSmndzrqh1SIpV6fDMvwwyEhYOE83cMd9I3oL8Qh4S
dpD65ewublHNoJv+dnyIV4EcB4ItI1nrr7K5DScQOkkwpl3MqFJ4wFSIkmr1a4Gr
OeRbTmkA92N+cQUb6rfaxeqk3JX6fJGQiU6dI7S6Q4loH5JOX1lN3y7jYIflImsv
uclpF2cGDdMvBaWqHwSf9YDYyDVF3wgEKlTPsUsDN++1GmjmM2FNWnRz5aC832yd
w3oUcOxpqd8xLW0aADOIp8sSMHnlt/VtQN4LcVRpA0+Yh4Y+95ukdG1Q21M/Lhd9
k0kyXfl/JdXWQ7aeNMIEwPhMOZMnmOHK73dAm/xsDzUuItyMF1mK++b25etEcGsE
3fMRLWDAwD3jDDY/5xjFufi6v4BqnZMqEqejm9AedKacoDokFSs/bWEqYX+la8Ku
ZJpXnfh4NvPUiNNysCYBZqqOrbSgMK0fYZQK+1SRJi2fVt189f9Twq7v1WJMEILn
MTGvB1SvCE+kyviDpairNv+FE43nVDyOwCAS4c/dAWFiPm0uYTNz2mX0ADSiuVFa
5NytDT8Tro3J3yRmHepUJ+zA0dcX9ym52mI9VzJsBnkxx8yBmZ46R6wnVhPJK3ju
/dbf+MHvMs7QHAzx6D1vQAhRUYj8lYWklflxUjjuon+njw1T7u2Ffvc+FrF3pYZA
+WHfyzUcQMKL4J+JBttow1LFGRPpPYsoIn7mkWDkcIbQXc4GhRZqpWMBpt3ymQKn
3GJ4y9KOFvgPvi4A+tur8U4f8zKrr3Rqy6Kyrwf9niRpRudeZSUMCl/woidbETeq
GMgYBgKhm/iGAry1cpF+wDmzekj/I9ReOb/fLYEPKQa+ckdnS/iFoPxv8mBn4yEk
2th8LDXbyAzX+G7djs702u4UjAp2KKoCZUHWMt87vnme+EZLRkOEXbyEaZSex9L3
XZPsqPa5EoWLBBKprRhpochO1IBEAVqQVNbczF8OAuJXE9L8mYwhSN05+ZX06m+z
gkmWIp1lic+u7aF/xpD7qoZQJhD8YRGxWrN2Wp8spRjOWy6DcZYyrjE8xHb+snsd
aTW1ez+t3r8YDRCl6/G0MuROIhIRwC/wHBDy4QbyZ4iK/w3V20CkvH+sYLhcxM0L
Rvj8j2uWQJndZsUWXoDrn9QF8G5NKEg65YiCABGTf/oxOZQjI1PYu9DA0GvQBhDv
pE1ru5vOF89eK+gSJOh/KZKXnqlijEr/fGc+ZIaHL1z1zYP7RAq5+8VwK+2BWAhZ
Yr8xwNp5NRxRGWg7iD0/xDNpvhvgLQ7hZ/1qlCskfWFH3x7ErHIDYntByk4U82t5
l0+6hQ9Hq6eXZ+s3ze8N7mRhDUF6YCaTgj6lc5qEGNIRFDnRN0qvbVV/1ZKR6Xm/
pYAbxzabSRALFUz1mfiBOEWaxF6LMs5sfOvxoESg6vDwPCeZTNOj8Ahjnt7RFbH5
EQGanq+ZGGRaY+p9WbXqfvLO8FSugOSeW1UcIKVdXijBtWEsUa7KKd8aMkT/xLxp
sXUXQgb2TztxjW83FSTuhBVij3eooKfyfNB7ckTQBMel81QugsuP919HwZqKnhnU
bG87ri6/QF89lGXOvrxFd7cS76ZCFQh2o5dG9+UTb4EMBQHEVwL5J5rhYTTo8cMN
kHy+g8hepErx0PZECDsS1Td/0Qcikqwn2gQBKYzBIsGaGU684Z7L92Avty1fhUxu
w/2ljsoQAzKvGUUAYRFeRyLlbV9xxr9QZCL5VOt+w5kvkbmaeM7G7ax9HfSdq8co
IST6ywq2eoVysYn1soxfNcTA0SRP2dfIm1v06qKkwUb5EzqKw3xkGDqOgYzVIo1F
AOkTaD4kc0Jj0cXw5O6B21GSZgCMOKmY4pni6QmHpzrI13GNPO3zyOBB6tR0REY1
yIsuOq+CieCTxE7SFIEXkZ5RYGcZLSlv4YT5drFwdQYs5tVQ2B5Je1DeEJdJCWPA
5rlAA6jSzmYnNx7ou3Lknk1KwfU2fAOmM6i9e1N2dJFQZQDaxQKVoXY9cNVzb1Ff
NDjzVQf7pwBNl+KTbOiKSfeZJ+zak5BQvtFhUsGre1DaAb18Wv2DFcfHn79GgNQu
pZL4LoSGnAqG9b7gTB7m0OFS99s/iNogLvyEj4WBvpQeZBmDY3x2YnPv160q7V+e
6Ko5SM6kw12XqtINA/XrY2oIjBtg5NU/HkyDDMlvvVfWRWtCnjofQy6xlCmxM8be
/fksKhijVybSIlKkeWtoYMxaFTU04mL2q7He0WXAsqP/7is9LuOrsNP29a03lI5s
GiHUFNjIEnR5y+v6/5w68L7xTrRZINfE24hlkuFNqkJ3hx6aDrfpl0VWusmeIjiy
xTh4It6BtZEcj1FYqMl/lwIOqv99V8B36IA7WlFlpOZ+yFi5JeMa/Uu1JnlWA6PJ
k0cmkjuyu1MamKnnwoi5IbYGec/NMDQySlOmGXA2HcupvflXjZbobxwITB+2wkWR
5QRy7XiMM1DvADupNX6qLmsurUPKsgVMvYBgWv9/KBxWeJXkJMKeaANXIE9pP4rD
W/aehSiOrClrNwoYcz37xUR30Z+DTRLt6w1b2X4dhjiYU99kW4y6kcMMNg06QrLc
ky3Ce1VajCNYo2lyAhIjUk0fB3d/7hw6T3SuYiql9CkR6btXCuAh8juBQxOZQfVM
sP7fyNHg6Rpkol3QyxDTWwcW3nA0qO7fvvOa6OvKPpozCgRiCBTS0prLHBcd2KdR
trokB3oGjaNTcj5o6BwFf16y84leMTlGkcyoLPVpgylr1eNrI88vH2OUHz9aO3j0
onJYgVYizzljE6/6yTSI44Hb+VhcIHKeRFbSM49NoNQ4llVcU9rXGlsnoWRDjYZI
06KPQNIZX/ZzUGE6aD0XS4B8yOtnoNDXMMBzK5FjtuFbbec/9Fj1ZhtgQnoGoh7H
ShKu7mDQ3LN4fHfxjZ2E/HvyB3YSdTarAU4gBPu8stR/RUllF8c3/hv5ay5ycA1d
98zDF7L6/Vb8UpzI6wd5rzc+wEB7jlg5k9AcK2NtJZlfs/wWmIbYF7lQdiX599/o
5pRVxO841LRVHACBxkrwIrR1kjNd/25AIIesm2ObRp+VgwMPZr8QYWY8oaG+ZfBx
oD52qN6yD/aCnys9YPpsemaB6DHYU4Qv+5RJ8jYBCmWJ2DFN7fYAkJgZGlJbAqpA
//qHZyhdDdr0yzFRgayZXlZA+QVwUEjZDgurw8WM9QkZPttf8N+4Mo29815lPQY2
WeVueSjLIz21dR8DLvLQEK52usPHHKLpvFVmlI3u8d8dzcFkGMF9Qj1dQ4589ZE7
yc4q277qIPdJTVmrCCh0UHh/O5hGGZIZ9ZxgHk6YvoHyC3IxhHo6GZ2Paow00rHL
VscFxgcpsEwoTB1z5vz/5ZbJEPKZQNTWq1ABKFuEucHUaJtN9V+1us70SLsEyl14
ChuPh+ui+UKZNfOAOLbeq1W+SS8K0KohE/DJGG7vjdBztH3zZoAdVYHtVlvgidLl
84YIy/N1LWyGSU77SjSnNc1PW+aEEsaTnShzLnkTemY1x+5/XGKJ18UUWIzZMgQj
w/SS/57cm4fndT9TfHfSJqzcs5Ys1pmA+srCjMCsody3QOkSq5bgjMete75MVAZD
CkQ6AMndFqRPM3GmfWJzR5aTBnYZHpyOWzmafSNS9SEhvv4253XRUSExA3Xwygz2
vfP1NvOkMisuJN0OlBj67juIxXUFOGv0kdkijp0ui5pDX2yLthWgJgqcdcfsXWAa
f7N8Znfr8CPMGqdh4wr4si6IubV1AAeMl64+iX2beCsTnvSl5qY+Xz/NzDbi53yR
ztJJvizSl3TjAvWReeeXppg24BNIX5F/UtCn0+8ZjSxnQ/b2PYzsadnYJKCu82pq
U5VbdOlTSpXDo8ZRzhhC27N7mkZVjyTnracKoVHvaNjCPD/1B//C5ioTPT6E8bW0
ixxW5YSSa0Hge6QAzd/m5+EkF/3VoKyVw3ewY1zfvgTBWbeLq0ExM48i0+rIOdZz
98DLIrEGWE0rYyuD/7YVgF+S0gvxHT9dCXqwEFsu4y6Rn3ScgA3Ym8VV1Xy3QNjT
uplpu6zkArmlVGxj1SxIgl3ybH7zP8j4eVhMC80t9gARpz63rZUTN8JsANa0tW7C
rJZkXG5mQ+gFAWrvb62muebNXYjXvF0M5oN2+1ypaOPJzlz3zcPwDcflG+f7+QOb
IXhDQM0zh9IMm0ggrt+qVs9eI2Soakuq3BSOpkruMcC5w/fb3NHfvegzKPqdkCcW
+uAI5Y+9VHQqSEd932zxIBZUUF2jR+EXCzfwl+8BbcpESdd8GNJk2lL8uUJo5751
G3m672gJEvsfOenRCIIa1smMQJPjR6OF9Iu/X3sVV2f1f15aEoJp8JDxPqzR3rWi
iiCpLh4Kiaj5EU21eOs372K/5V4SWtl1VbJVPotaKhlMjTwxJtilEihhJTKndYCg
ZKJZ26s9+Sx2+Z9/JJ6Cso/q+oeSJAg55uIdPxwTpxZkkEi1piHg8KHWp1fT1FCo
byfwEPilmWHahqu2xm1Boz6gUHJs88jkngssMwIboyb2R9hK+6qzil2eeHrfdS0D
cPLpTcbRSlgld6VrkJJTVoHJcMbULmFdi9EMjKjxEDfS+ixFcFAiKfusFitqwXCJ
fzpL4CkIHScAXN5LkpddUaMVQY5hI4vkuuVu4BnCnyIfcSnEvv1uKXhLsSaJZaug
h1f6reR+5FsESYg7G+8yi1ZW+jIBvsjFcJjJvgyBoKrPETSn3JYUyPER9m4QP0V1
bw7yLoGc+PyTAeZLCPIn5Wy7BCmI6zdwhSqeUDCEZhvfy5louxXrFdvQHaEGNnHX
n4XhhgRVrp9aNmQiV9FgkhMxsEy/omYu1C/oaDJYdim/qirzqrNtVaC4q74Znzl2
T413gVnHZHAtdNXIfiMmsGucxtZFdk4+fT2vxOmj43D2j22b0H+RqdfNT4GHXPbJ
jb6Y3TiUmyIlPbnuihyzcY/4yIc1aVTdvnCA30m0cWVTjv+TtPeU37U/Lk7uPJoX
tWG5CstOmnMKE1YQ6weAqMHGFsAMhXkkVC6gICTs0CvkAh6dBzWnX/tpbE+iy/e8
p7XzooWriR74qOQotGeeVUk78NlU+a110e1mA9y1wv/g8g0FszmCDm28joD28Nk/
BWevx6iJ5HKD0AitCuEDPDtyT0QpK2Ay8d0nCrIzAIDWIsXK8+5g8sxe00AVEPAT
I/xOTJgZcKs62kAhE7XjzVM6HGia8RPl6QmkbwKZvwdzRqs1dGqrA4e5Qn76KVq1
epl9ACx+hVfupVXVCea3NoerdXV6hetfF46WMxdjHQxPrRrWO8g5SFh7nsvOr2RF
lbjy+1nDSZQFOPwMcJxiQ/UqzapWnnJpIHpgeFy+kalXxHikurw/oPAJ3JpceVna
J3+evm9nLnVrqC9RMGVzHWclzpzZztu0MerPI5Vz75CzWc9L0MfV0OTPiTq0fwZ+
IlUtnaDm2Q0cS5SzMuKtkLk8PyNGML6RR9ZaMfk3eIePy3iEUdw2aDS9jKNSA4Hk
27w6SmmB8blAl5CWjsbkqtvjvtaCTHtlytXqnvzt3omVo6DzBYF3X36yFftxNvMu
Vceh+IVNrCL7Th5ek32euumyAwc7sQWhN9xdYgafPDWoz2eKY2l44MBOJb2uBofn
EfsAuEJzsYVvHUbGJTRP3oH4hr4PS4V0SO8da8z0AVBXH7lMc11dFsxk6kM66org
U/KH6/3dbDn5g97kvSINxXKf76DJQUDfdHJSCgRtmSbMXcAuhryGGWyhXPX52HiL
JkEOiLCR/loRPkWOAzoUyeTk1ZCT824qUAN7lMY2rSp6G6CcFqGB/JUjwyAyxbkn
Svp103sVblqipNPxZQ/rM5k3olFhoih2ZsaYc6BFAPim/qAqf/HoEUMxMr61tt/y
tHNUgH2gY9+UJlOibCf14Es8BfcF0XW+A6+mc3LhMcEyops6agKNd1Kz9G02aGbH
Mbx3HKqE2/4M61mgxbR3bsFG32iFvEDpwK/H5zhU/ATjqXbW8az11szC1d10X7OM
07Y8fVy0LXdh7xM1rZkwBGWVT+czcT4ERbzY9RKnTptVkMEEnSDr7KuR1actS+G8
jQw3moDrvXNXYjTlZvYjpJDc9PHAnD7Yd5UpiFhznURbWkHInRrWxAbC2bteV47V
hD3wQmEpXLtuDhGiSJOW+Py1z025RtQP9KcxF+7zfo/nZ4amLqkgnsZ3t0qomRij
tSzdXmMj4Tx2V4to6GPA7JIodIm88ULJHrSvnuzWIKdBYixOfvNTd4UgzWFiySUp
VkM8hdYpmyP39mo0G9II5TOTrGayrP+zUcb43m+zuGkl4tsvF3iR9AxPI5BYnhTQ
dzz0/4N2hRsrUOI8vqpu8Y8470uF8UlJtllL1uc0G4wqM6gWanZ86JjBGiE4tv8x
033FZ6+p51rFF3J3un3yvp1XC/qTn/ySh1uspLaVVP0nijtvunLbTO9arfBJGmEx
JCbzq3a+iuKlxxrLpsXkZxUb1Pjz09OffKNiC4a7UV4c0Smab2G5r7rw1l0an49e
cnc6be4CWAPJKSq/XnTFMvmPtQzYQ3XfZX64ZY6kChJ9inhwNqQxtLIvHLbRfNpO
iWAoijUaqjuCr5+n7y4omqKiSJBnUTHWqhh5zSjsJ2PB2wjc2AsiJcK5UuQloB8A
v/lmEiadZfS5qLZKqPmpdDqnAt46o4dlasEGIDg4uJVha1U3rtRJclYOIt7AwNAj
9b4CbXYdzlR5TvuqSykM3HJiJ0uytzJJlkpn1lU7gmcCw/wSc5r+/trI/h2rqXOp
6rl7851cVfB3tOvYk+BWjntBlH0lF0bDoCMuU9pkYbKJRc6VwWSooIjfey0v6xmt
PoHFoFOr33C+mnnCVswDS2D+HyaIR9mGQjWByyze8Fku11DUcxTG6Oc792Z3SI4t
58xHsavqwU8E1JFFA5tkk0AN0vzXxHJdphScML2Np5GkiqnhD4YerBXtUQZ1n8es
TG4ckjNP6wsPDKlDDMgt776RZmQZbHR48rfRgLv9BYEgPwsA3/RDTg34goHYw0cE
JYY/Qr9jGFi4P8M6MdZWWkS36P9mbFpiypVLhg1zyzeQymQ9zujzmRe9ey0ajq8V
tNWZvkwW7MekdtPWvOMIhCGcFquxgw4bHumZ9weWI3mzOLOF4DTlTqlrpsnaAhSS
lXseClJEe4BpTnNhXlrb/4a1sjVzkyMjh9u1+f+38th1TR5yWm0L/by8+zzD3tOw
7JDEA4JB1bVKvVzlReYKZarU6tqPt7SKR6TC0abXwO6ixDVDFmHAIf/GmAYxBAQO
UwZ6Kujf82wUdaAVZL1K7COA5AWZC4wbmdtfzMkiZeXCQT3lTpLZFo7KhIUTKJI3
EjkaIggouzu2WvrSUC+9T2/u4dO+9HmyhxOxk9svH13SWjEepQv6bpWqvXLNZ+LS
RSPYU4JHJH8hLJ4qWwO0zfkPPIa2Teulkt1LfWXJ3tHKGV5n2meBGlFnE72FDmDW
WHERJucL/M9sdrYqtNOak5CVl5qQYFqP/wLKiDmySsrLvzTSkpU7fZ54SzUuNbwA
UdrCbJfNDvT6xEKD0czKnXwl642f0yDevtZyvBcbCUrz2mVHnI7XOt7MPrGCCFIn
cwC24H+QeY55gAyYOL/CxCMdbqSWO/26gxtVmcPwnmywUlGE5iY7WL9StS8ET7BH
8fF1b8sRbfr1PyjjXoF76k0mm+0Z2x9JD8dzaons5Rodl89bHHQUgme1u0Q+jPk8
Yuydj23T/5dva4Db9v/NPOQTcHaWy479N/lRQySKfWc/60kX9EPV9W/dOSJEn/Jo
7OoYS+LP0JkVIF260OEirNm0usAhcZ18RrlnUpyjpAiOakK5SAb6aw9UHbJl7Wai
VTM7cozbgSuneXD4l4pAdXPB7bqnqBLMWR8Mt0vsHz0SBN/C5gnUWRn0eOqLZ9S0
PGh2q1NgCPvV+NuOh2hrjaQyxEIefWwvf0vLnKsyKVc3bcgXJhhVpELVXKVaKb+n
WkaLEEZujYHoHRvJ8rBq3u93j9VuQEkeMBgfJbYy+7A6iEdij+G7lXdrifY4Cpbp
Z1mW/VXcfM0hY5MxPLwI4XCefSk8x6EO6HXvvB46pbW1lnIYePiTJW0FNC/PVo8x
V4yLLMSrTXJZiy8ThgZmrv6wsHfu6lLoJx21Fei1RgZwl1S+runJXLevDfJPp/j6
YwDZi2R56rWbefXX/45MMXhJwh7+bITPiq7V8j8z4Gal4LLEaRXlrUk7VOXIXhvo
AhWaCK+sdpTfCk20m3pI66wfGSzMPlhSBT8uTPv+AmtpH6mHRD7CTgxjrtlBoPq/
TxviCA2i4kcDGIvpU+Ucrvk6I2JBkNIXpzR10BsPOdk+y3S9BpCaQnAgo9oELgK2
vI99scFQRqCapFVlBJXF7g5BVYLl0WCO5KNdOFNX5AL05FhZJC3IEYf1XiDLZYti
0P9djrCULnJwoI4FpZus9y3uuQBhnrHqbsXfRvDCVqIpRXiHTMM7wbGKeURqeLxc
6Cd0ibcYru//RXpBh4Or0R95Qj557yNMQ5Ca6IK9ENyRpshE4gytNomJHR+fj6MU
qyhorCyyN8DcZeWEFAm7LQdVPyxoDphFQGcDk/AUaWl6t5onJCTAT5V1sK5++WFw
fapBU2vKJ6EofLJwaEUYM6QxVUgibCK0wGDGnnYF4lFCWgfT8Pw0Cm8OIfZMzRgj
+M8KfS6eX7Q/JAPF91u7Vy+2DrBt5oKjkgMbxUD5ev3Eo5GK6rwf8GhA6aQLBRwv
uKHDQfo3NoCLSiGbELOG/rJFyjrftqTSwG1tk1vfIrHVUnlcQgC1BtGNwPLdG7mX
hmtx+jLYKfTe+wbIwPGqvDNmcLZuVu45XnOHXa8MLAy0Ot1I9UkQfDn2YABAMmoS
z7ZkHn0y3t6IqSgO/0VqpbX0ire2o30FL0RjIy27S6YzW8r28p8jU9VMrk0SdE1Q
yLk7lOAFbQGOPimUepwbidXp2hTJQAXr9IGI492LDdukVsOC942Ole6ZueTC7WD8
kwdi2phxXj0eQF3u0DEMZVVdjo0pB8dZGDqzihBCW4e6oUx9UCqaudZBhdZ6lTXH
aKYcG2w/VsJAJSHLx2Jelgef7Xg3K80WLp7ErDkCSP0enozq1s3hE/BEj4squujd
kqyWQSfi52xdjK/pJ1XBAalcRf/Yx7dQHSF4Uov9dRQPdlnW4oRK8xYv9FVfeptb
o4H/+bdNPXwH1D5Yja4827mH+tPl4YbawuPIdYQKJuzeDUuyVDXBZTGZI3JD76pV
KB0ViKWLYQHA/d41G8lCmmuY0jvFFFgayY4CJUjCmdySjl5l9Ajbub3iLvCXZ+fP
hF0rcjz52Z3UpBdGoapW7ITm8D8voFMtU0lPfSUb3F1qeGU/q92pHWrBFJEfDwXA
87TzWbyDzNmOaAAwuvewvobzAKemdmCymTyrE48+SDjD+vZLihE3Q214dUr7TE6V
QHBlN1kU16xh8fZ+9AIe2Kke4d7wchJWfgExjxU5ScVu330ODVUpAhyG3WV/VjaF
ZKfluTjMEW4ppDmw31DPwXGAAiVQsGTFv4bPFvHP4HzdBLuuv3Y+Gm57feA2T+59
pK35yhmI5zOoO2usL2qce1/aGlrhJYy+JTN68MCRIwqhVQTnSJt1JdFa4uSuP7q2
EpvryVC2bErptbSHlu0FoMgZQVr18aW/bxLA1FB3oAd5Ud7Do0MqY2wstYcSryDR
cKkqjExsmpPvg46dqNvKhiLpwK0NlC+LTxBw3oGiO8lPCP/UI2cUvK8exQ4d5GQ9
K2Q45F0ETGGYeI6qVtOfbGHhAPVxJe1PAEoyEe3gTnSHDphB9BEch4ngPOJ8jyz+
RF1NkTk1fyIwRriM2TtaN2qXxKqpxlXKIh41Uv79AXMcRGK+M1fGdJ6ZDjMISTI/
1ofu1K5KGdLHrfGiRxRJyTMFsvHubD+a1Pc+ZtNGznFQOmXRMSkT9eRX8rLW0lXu
jsKwGOEgBa3BZdoSetmotylndLwWBquQRkL1xR0hKKqnus6l94WV9E+gHjEV/0zf
EsujdpfQpr7ilSOAOOIUkHpXS4JQ82Yl9awPeKpocls9tDX66znbcCy/K0pkqQ2b
qsfAtmShssPkwcP1cz9NZxBo2ETUWkYI3vX2lDFZZPSFZf25J2Ej613rZQxHQjdb
SImIjK1abh+k/ojJIjTQPxIcSoaAHgfR/+BWSJq+x2ml2vtYx+1jeVTFqFcPhWKT
XQbZjltI0zuRt8CyB6ZCiGeCbgs5YpqmpKliV3JkWPvoSLcbFzGjoFrQvdKjFudZ
B/refMQt5x9Oi/UzaoBOFj/O2tzHpCrc1O2ajYMN2T5gOLK/WTOZJUWLLnM0tbO0
vS2EQq4O7+RsWnH+XB+EEGIHDnWvf+CKnWgzwYoN7nfOCfp3n2YbNHsRO9VAW48r
dCTuaq/0x5B2tvSQlGkNZSawyY6D6HHeog1BLlU1NJx6sWNy30H5Beoe+LuexcNo
n0evTGYZrULKrFx61Uhz6wfc7J5fMpzl5Gu4swKZxCN1ADOV41L8NbBjokEd/7T1
pAUBGp+zl2PIL3UlvP/Eork4qpS5RpIfMUVCZFHhTK4U7/pqMM47hboHmKaDnlET
CMcwS0HvEFV6y/MPeNy59nwce7q/sw69VWYMvQD7YpwifcxieO7FbP2LX2nf2kZ3
66IeSDWrHOb8hPSvb5+hnU612rB5z69dtgXSCGkB8Um5f7m3v8eOj0P5II1eyqkD
413HYjaTbniT1mMCvwmG106GF/jMvG8CyeHyV20dj3REmI2Wi08FFrttw46IYCfr
OB2A0obk4VdZ/QIf14BJy1lg37egST99dStG71jttBf3viHwc7kjEg62AVsP1/vo
iRK0ZxKm3gKmkBDYP5tN1fsxaQF+4Tg/TgMfBZUxi0oUbJp0z/Gs3vC+nW8YZZ7T
rEcO09e0tp0s3HSzMxabFhbOpv+poMwA4nKgzwa4bnCkMbxBDEvdp5az2QyBSiWD
z/1Cl51emhntQqhXX5bILs0IapBWJwaNh+WuYYoYxCNTYGcmJtHl5ncGsHmN35Hq
XqmjqTBvYEW29UXcwtNeA74NQd1/vUnUSTnbfbVubGbczMGGfcrrPBV1ZW05DWfj
vZIuslqdUL7ftHB687CN8KhwEX3QcYHj0mkbRPxBsXua4TorVK1mZH6zpOH8Y30n
1zS3HBv3eMEdpUQMNrsuSEP0MruTvIijw+GwcBn1L/jnO4lVaVI/m1O6HY5AymjI
BFDTYbaWR2vvxPwvHr96f7JzBPn2FuVyZATq1DS1uJ0vDEAu2KH4Se9WzegqjUpG
3xn6tUBuPvbeZi6NO4JYSbULpWw3JxHKUbFdElPkP0yTEZQFmlFAL0/DStFslGyv
guvMefJWJkqwSJ+ZiRnxuz16frv2FDSSXprsU7GhjupqQ3XRHrJrXcLwIWWj0Sro
mPKFadAjFcMRq/y/6+CtAXv2CSctcuDFHfbCewUPHkb0R0SFVeFW4rLNV+3DGrE5
41/gR7t2Qpomem6JhMFRIoJjBvT80rQHXWbkn+n/iHKao2tPUZgXSJmfMr2nJcCi
meqGhAUeyXc9Dl/JzlzZCpF1cQQCtG+BaYudm/Dlh5Vq2SDUBInHecnf1nx6HJmh
xr/Vooz+Oxc0qcdD0ySOR0IjagFnzIF3VO9vRAczkBmupQ0lgyXVgMTV240y+NH+
AdBryVrrPoURaxPxJWX+46TO1v9vB4W4/TFm/akQTyLzVxecVwef7lHgPudE7Cvv
e4AtX3lZ2ZP4fLm/Lz96k3dq472Mo4dmWsMd1iNIBIQJmSb4PIBsJQhn2EeXzn8k
0xC+rpWBjE6+olvCkRIcJv9XLtSWKzk+9g2E6ZdW8x1k5tqU8YK/Wr8tfoTtMlAp
oCqyEoUD1D8YubbuSdDqZxmFTJaud4n/xyWI/ZScw7QeJ6fCHZwG744PXICPMm7Q
ZSNkL02BQScRWdxnUgBhWf7oQE0TnUW7GcTvQJzl4HODXxi/B5UTsgHkzR3LxVrO
2+dzxlb7VxT1IKwB6wfG3LyeIn9OWCK+Qq38hf6jTaFPZZx92VyWlOZ8H3OzvMpZ
zswRNk1rdaTgul5LIwozfne0XpNtlwLa7HGrS2U22HXOZPDvZoY+6Hk6oTne5yVd
ktcprDyHSV/Z6zdcbWZbiH9fYbiWeNuN8vrUMnKRYiqzlTQafXkPIfcWRXHSNYnx
d+4PC9ep8sgz1BEi06pAs7/ZXefBz8JWIBY2tHfxsTeqazUk2X1BRcK0E9nZKInw
qJ6vtxPf06k2O9Gv44GWdtf0jXYKoTWi/lOxIG9xtOTElD2nzpKUU1B8DQmSO+Hc
nchxeSgcaYuTla5aKRrjDo38DwP3xieWKkN59X/O4soOdTeYkOrJJbO5vQ0FhZhe
xj0GE/VrEwMYK3dnnowXXoAkMcp9bqWf1VmBEDv0mceeHJV/hksiQvyRTQ44uLts
VYpR7mmnsS97Fc7o6P2yjuvI/20LAXu2BZKHgIiaASeExGMv8aam4/FQsqvJmbEk
vHRGySf/RE0yUdvDEULiJWOdRl9MN0PKh2ggF0lfzHPnimg3Gxpb1zHrcqY8nlcU
t4xvLm6mQU7Tz4cDMc9GQqistO/E23gGpvexgHNzuTA+eWKQg7hwpjbA4bN1pCvb
v/V/swYWux0MDj8cDhgysNsO3IOkYLfPaJUc8CfjUqNqic1Q7F5Z6K5mKDq9nee5
/g4lZVQQ2NYqYH6ltt23Csfo/Zj8jdYrA5UNHeKIP0e2FXyaaic5mOoLIgxh6S4D
L5O1+Rju8BC72OiUcLR2QvL1Xef/fZ4xUW5uPFT+iYATcaZ5fJV5dvzDNqShusVT
bS45hOwYQTF6J5F2pKlNvzGgk8y5uvVLHmtaZMu/QZHtqIZIVZW5UZ9gyP394/db
WRMN8BciIU95V+zr50CQOT7Gb9d0zxWs2VDBwkn1ejNwZGgG5XwKNOwOK0zlAm4H
B2wDNMkZvi8/6e6JjrQneJz2zp8gEw9t3glgvECLyZ6NLYzCg4QeChmgRYE0wk1j
lqPeahH4FC8SIT5R/ZwkJKIUCjTiWNL4cy7Req2cn3Eng2bR7o0vFYrn2HghT1uR
KwsSJji+TyfRBzVd99ZdJC6833DojxsOW5Hwa4nL1g4KXEjlF6oBWyusFursoiBe
qvLckAtFlhqgmOsiz1LgiGuMjN2xWm+JEgo12q6Xe1yG5OUrqQkzm1VOhNyyLBR1
ma1LWlzglgJq6jwsSHOpwRIs7xjpDYCXGqx+BUu5gV6gQrL3jcXjTAHVO/C0DYnX
kyygWQ0EqSH07M+qhulso/dFyU2xfF7K4GbXw9FShpGVY7NzIBEUBs1qDHBTKU4o
0tJGIEm1T0oZ4fv0o/OXiHgqB3xMEFnn7B8l2+TYDsxjVbzPJTQL6D1v/mFHfWtV
YK8n9RonTvsC0rippJ+kTdgYeMybnoaTfI2nmGQZnMR01oPfbcjKHPtU1NkZhtoH
VrEofhTGIzghzpIX2JldpvbBFEHgwUIUFV/NioJFCqaVaoCBLCi6evA4IcFh/wde
zqvdc3twUHtKDxRlsra7Dv+Yso8JnMVy2vU43ok3gpohj9Nqu9APH17BcwgYWy3O
wcixOm98XJwsAwX6KcE7rBjDYss0QxflFu7avEkQ+/3spAv92UU4DtMywrmyKw17
EkIjhILv3y5BnA8+Eogo2TMdHAjK7SwUE3oOqaIwpvVdGq/Dp394bg6nrvDFbeeh
dkMTYTy9r2v3g4Kt1eF+54QnXkZjuP3dkrgOBaZxezG+489wpNs9moXox7H7IHvn
cm1EnCnstV+GBC0NYX+mUxPKRUtMqaeOutQxCcMTFe5h2GXgEeoadE1JAJOzYpwu
+6wjG3VPXB3O5GkOrNTfte1K4kxy/STn49HKwXGw2vJEEwVxXG1UYTpLBoxiE+Rc
MnU86piEWiWWoAy1qMughGfg+CBB7TXNd/S+C7ppieLLnVRxFAUMzsM1bpmvNaza
ap32TWRzWjmLNY8CHLRvYSJ4v0CcKyux2UhIFf7bAemu86WhAQ10vocSxFR2PnnS
Glr5JtX7oftiyuwUWp7LzbNHtppk8EK5dWcdVgUpKl0wKdWJuhxf1PFGYQQge7qS
B5yiUD3DwH3sq2KMVbmlI2FYDCytsOhziIFq4aObrkY27XefafASj2aKViyj6woI
bPRVg3cnC7lNbqZtR2+5xjvATiTS+G/EWfxL4u7bRG65wklfsLHDlPTck1JKM3ru
24d9lJsmJ2hXj8Be6PpqsIRJJ8mCRE0KMsKLr+w2N8AcYf1syGdKg3ZE1bmC+vYD
ZKoCd6kY63sd1fk3zRKyx1yu9NMPMTFznRumoohuzLTNsi2Q+iEQQk6LPJsXXuFt
oAYROdzZO5X3Y86gInf9imjNY+3c/UZzLkEUTtjVfQz3VlV3WsTQNHJKdQbS+bb9
QIxNEmTFvzIuUjyt0jhPTcXea2fStzzaRexl0ieUuVQbueAUpor8mmExn/A6712/
ZbqNHj3ziJZAIu6JqBXLs7YDkkQLsA6yO/sYLuZuDfHWYMdUszmZ7qZ74twwE/ry
7hS/ODxIa9qmNwRG8waNsW+R8/6vwQcPNaLdPOilaZA3GX2LN6adMpXmRhjUNxPb
vENeL0Kl/ZzQ8y9Y/0omzs79vSb0AnmOFOT/EGcXl260zjjmrdujRxQ4U0ZmPThJ
ooFQmKNyoSOyTS0YM1mRnc1rIC9Wy+aZY4blOFt15NzZklrKMuB7185iW/MrlqOE
EPotp6SBS4lHYAN3QwD65EUH1pp2AQ+fXJ5a8+3cMzYpiXNDJO6WR5aysflGXaOm
x/SjPJcKMN973sxp8ToykMUV1qX9umDZZwrsTIFxzchOkteyEAzRoilCVYNYqD9B
2Fji4C6uV5UOZXO/3scvu2Qmsce/5wqhOe5AHAVA1Hw6R2hXEvVOzpJkvMtAXaKl
t7RhuaNtIT0267w/EiZH5FEtvjRsx2CbPg5zc4pHInzScrrBkSTJhSTdbvI2zAHP
j9dK2dF6TfvDdGjFyAeGK5znDaUEl38RTADJdNdoFC513lZp5qByHBGZ3WJY0qFB
fK+8B3VWiLyU0nW69L6gf08/c44qbk2sd7Sw/dpOzGFMmNpvPmkV6oMEMZJDhrDT
m0zADL5i26JMsXFLLNbsMhIKi3WKlt/ZOxbYLu85Yi0GVucTNHUWB8+3pdeF9yyS
gREvebjlERqPZxMHW3GV4B6qdRpaqiOGj9I1H6DclZbBgE6ucfO8a7PojEbnrKz2
mI8nFcDismsuI5im73sCXTRk1qdD9NNDrrzcwj+AERbhyWbZRvgEX/Ay1uKpwMK7
WE7jgjbpGiMO6ZXepqm7FynvDWFS4hg9Aj9jgmhVOgXNZHaBf/MJ/cbIXKjqOhFe
dDzkr7JEmYUr1ENGz0uyNQG63NxOOrJSmpd14R0nF2LdNgonF0GKYF22ATpCJD/6
Lxho08ZsmrdPYNrrybsFywotiTKdYe2bt/pmIO7M9pkPEeKaACmoPoNz3RJ1CqKb
dNbxNFoyMx9H1l5NxESqAusxo0q/3B88ZkRfeP14M8jiWl35/DEC4Hg2YaQ0HIMV
4ZGqlbu73O1/3jDXrN0ZCtAionRVk92bPY/H1hg+l2C9GVAsL9t+qx7skIcxF2gF
3KcJwqJGm3CnEJN2Hirs0gL+9UI7UIfrBl1NGMyF0Yh/uacjq/zXd6SJpjZmafc2
k9UFEg2G8Xmn/6sHKLZ8GkRZMxxEfuOKBehMaKBQKn7UeHLtO/dyNuN2Vc8j5NTe
ZdpvVi5pSfyJ3AwBMK9a3X9zQkRXfEckLYIwLWY0RwJW6oM505Lb8gEadmSF3C7R
A8Qcci7D6JbSm4lxQ8P7oDtWIkValqSRFg44GCdJhDdGm9iDWCc3aZDDkYlyXbCS
gBF0dahDgCGXTr342Ocs70se6dYbAZloinLGHZLMnxgvgMJATAv/cgO23QenJEzY
b8+eXtPy8h7+Jbf/86A6pKCNdfOJ+CE6+cMluyj8ywbXbCAoioW3itX4ydrjF5De
zqervPKh9ZNfySQ1lUFeXR/DrdkAiNnhJacFCXVB62kO2iPUQCxSHj91u0WxhdQq
y0FhNx54W0Pp+xLRdgEO90HXjg1Jt6HlJ02/lZA8k57j0nNaopnAzwbBhnBAJ7vb
xkL6prUiub6sR7RXwdYHi+8vMK0uTTr+Z0m/WlRBgjJl3fuQANPfgMelhuwcl2j+
LMjlfo74hgW6YcAfpULTm4x61VlZF2P4bZO7YnOfnk4GM3hQ4mRPDZatsqEz6XAm
vuGabV+oaC48LqBP0lS5QEiMvQwrK2S0fS0iJj6H31ZOGPgKgbTWFt7q7Yxp9R73
GZNpuyxZri3ClJpaT9rtcEH0vDBqSaNpZ7b45Z8lxGOcPcPLznUVyiXbhDTe8sbk
Y7x3DJ5nxy0glyICFcZDmZ2M/daqoCpnRVKcVd1KYRmJUKdP3Tc10/JGmoj8SALS
0G7bqZ3vjqtl6vYpwoO8H9OX1YfW11hoRfCp6xSS0eC/VBndjqBCiYfQVafPxaSV
uOh+kBaXqKotHrH1j/TfFLyJ6WwRc8zhmY56AmW+EMtVHHBjrfLq3ADuIzieb7zC
Q/NwIjtfGyd/Gt3e09+ph6AhDEf3oWbru1syOQtu4YtZovLIfkfr1in01duhYjZp
b0YeTxFxEhkMTyLH1MlZEH/yY1tcC+XIYegXTC6eKt/Fz+sQAZn80O4hPmWfMvKq
SopONC4M+6Pha/zYQE9yGFzaJBI296xWlhOko/7m6QqGLtBoL1ade+UdEfSEcQgz
Lye4n9lcMMaTbIAdAa3/5xCOOzP86QXtx5TV47S3D71q+dnMjIutnR9iur7hLPUa
Kf3OWT/BHu06tJtoE7VA3HOugszntYJCQJYKdIM4hWLH2yQa0BWx7HKpGWHb40fP
rHfkL1Reh6UIq9ZcBuZWeohV1z1GC/I21j8ZmkzgN6bvyDAJHb8rXTPmlnkKuGTe
DAbkqE0gyQq93qFYTz77KaDvSUUW6vBC4hXl5zrE4G5qqWvjY1z8Vqd94VKXxwXG
pRX52O7zc1slGWfARfDfJPDA03nxRrlgnFr3fqC7LbpToHCLzODlRQD+4gs3qb/f
/DsMN4DEcFU+vFI/WFEtvQEHp+wX3FjqrGsrxBum1Ew+EOdJCYKvJTDenwaL+Mcb
+mPaRxzt1+wQ87TRK2qV9iXOe8C4vgxr8RVu13B/GvNrJETwai+DmYk+oTW5nAq/
GxaA9eE7tHzrVgu513u2ZCnaiGdh9a1XND0iG3CEFr2JHIKL/5zhkhzd0zoGDTXA
8Xo/vfsPM1yL30MoyjHvN7Rz/eukjR+956FEMZsFvmunwbyvCMeRCVt2t74BEKt5
rOfSrf1Q8FNEt1mS7FMnr8wvzPRyVWeJFrAujzm78GCXUGkQZ15xe62WoigmYV5t
tj8aKLEGD8jPCQEMqQ8CB1ljBvSwinuPbCIi9U/Bbr+dBGdTjV20pxhdixhnTg9v
Locx7QPmolhdFcVAcpXh+nVxpalkrflErY880g26j4xQl4auDVn1rWzCgyOqFqZ4
W4MFL0XEp63NteLCXpXTg4eES/osk87lScZbB9Qu97o6o3zGerM8NjZh8zP/EGG6
15wRbdW7cdgZCzYGsbtbCEyJkgsnZXC8fZioLtBpEsnc7T8DNUgwuGDHJHCbFRH7
L3cYQAt3qMBGRZ+Kk2HCflX/SxgDxjGlwr8vAldRvxx3GmHS0hw2v+4qwp6yf1dZ
by6HQpXD1PHprs7jD6i8DLA7fAVBf3xlA7riac/naKUeRNfblTbZ4dyvlPlH2+xB
4foynogiZ1WP039QR9jpYTRz2gOWQjVtNuejf2inLms+YNAH6XkAYKek63khPRbe
1yY5NkyZD4fhFy0665QyXPUYPr4pbYrDg7FSDjtTWMLPCdx/LLbOZtFKXPV2Vtt3
Hix//ogfoV1VlsmeFQTxbu70+1q3O4H5RuMkFoiFFrMPFGud+75da2RDzNPyUulI
4AfLYEYEzzQD3YHdkV3lIFpLYCetI09VVc26dP5MXyjEo9LhXdYyU7zGNjdrw+Rv
C4XQ/5y/VMCFPYRudQf8IxNhFNUCUYlLyqVvIHwH1MtSkGaoiHaoP63jSqHd/YZO
E/LYSDOdj5xFr10W2KbPt1efkRuRXmoPsvOgTSBBra6/lTyPvwVJUHNTpujxaOQh
TsNe7xkqkSr0PcouQk+3Q6lqD5S+puSnylTRMPy25zg6///Pfu0lMuXor4Zx2q6U
a6riII7Ju0T7JbyWowuf8wJj0WOyowNiFfNLBEko9RKMr11noLM6iQR5Ma7isOaw
vrKgvaEb49ELB89FUPSG68jIAwcc7gecuSzH0ELWY8odnd28cWzVHP2CIXmF42JB
64gMO1C//kQ+TxT8+wpFMwxQPiJO/panJExG2HSnc9rmI+Akjcuj4CqfgfOw7S3k
jMsCwQq9d3idFmKM9skw1++BEfectjNqfEJvJHUs4KtA6ucCBn/yOStFXKorrUpG
2zR8irQNM8EWg7W30mPWcju2evy5K6xlAPKA5n1YAS0jkvNyVWACPVZQ340q6wj1
eSXFT9d9FXDQ8u4Exb5Q23eGfl1ObmDafCexiPL0Kp6lpBpXwHP47PFajuUHeJJh
tPalDPV1lWEqwsxuUZjiZV50EtV0BBnw4zZA+qYJrw3plsRo1IosQv/k+C1ZcCRw
Y6Yv8d5jR6iOokdnKoiaTxsyy0D2jeHhIJdxPtRXro/zJeqXqtDzkyHz4+N05iCY
kCYa6p8dhKwIgSn+qxcruXhh9gH5jFZLu7sjzwRK7O5WnTEYpEn0XYM3XSSgZ5mB
0An42yxzaydHdDGvqWbjhchZY2Oi/A3N1Gd/rps9vtwjrABUcFWMBPp0oA9HtfXT
HPdW0yCPbQgcmXBis86PyoaH/ryMMsuhxAgV27tWA5h5K1Vq0A6ka10PLKKO2GTf
rWNczJq2EDW+TyNqcyqXBIBRHDE7gfs0ZgCfJyv5eVhiWQuJ4lEXJxz8XJnjBTe5
fMhexJJ9fb0uxP1P0DlsK1/55hlIh8NfXKbLWjI918EMsSmnLFQufbX2K1mZKHrx
jKkyIMQeQ0SqpBGa0VKC+yObEs6BMXJIg7q74B+jg+PXGs9pCikM6fGR7F5bQbhw
s6pbcbx5sNGTXbKtgZgoRiiPjbIvBTbypUfU8+p0gUEuXE9LucrQvpIs28ETRWJ1
IKiPpHoifJnPJEsJyEdHtzEJhR/jyxHPGBIV/U1Bb1MH5Yr4nD16zYljBOPg3JuO
o+fTjSyHYFxOsoUnlevutwMwhmu1iplWM32QHfZJV7LntVtRVrYip5R+0yVfvxwr
G+pyzGDbz9oPhawKf5T2weg3GWxj3IgRHXrE+ljbY+bzZdI0tN1P/0edlp2x60pp
BmUiGgaOL/PhojQkx8+EKRUZC5AcYI4iDnZjTa4adszIw/Rdug2TLpKYTwJNMdnp
CV+P0TSAWzDdbLFYwmtNPipyfx0iobuUm0eEGTtXg1M/V6VmGkmVgaOLwNKfatqi
FBMb7QywdM4TRQivVK5WHxbcgscNV/JnZGgoTZB0qRxFhigCvVR5TzwWAUCVHFGS
16VpSkhRJijahx6za8NiHuahfwSr1bU2GgLpqVZd3V+OZ4wminhDJmHdgiE1Eqyz
er3xj5ITQrSIT/Fpy7/b0l77TEOUi9NsObQ01oA1+9+rv8GK2BpPam2hqspjgIOF
QUbEONZztI524dfA5/4hv5kFl60Csudpix1Gs7EVyorh3V9FrqAitXbfr4zY0fVn
bEZB7QLg4IMhy/yj+CAY/g4W7jrzO1S0LY3y4Lp8myZv0CMsy3n0dj/j3LRfBhKX
ui2BEHKZEBidmWrplew07bt+PE8IZ3uJN25hTmuVa+5aziEfi6zuxnj5RcJ7WvKU
cLhhxsEQY6xoLc6FL9s/Y+3/JP80zLNy6Bt21Vuw01eJYckDkHIVLoIC5wkFo4Yx
D1CAXvvsbtQqpIfEgTXZtQguY1z0K4lPNfQN79swXjs207Wk8Q56wyvCYDkD92ya
i7DfIx/fXmQvR6WLVW1LUugibjZf10SrZktk7OnjXYsafJ+acbxyu9hPXw3+qgwM
ANNdPKoNqAm8BODKMJpIjKPLRbjSWeBHKOqRx6EdnbAwgS5hm/8P9HT9N7ykGKQF
r4MxOnk+H3FRJ1+4HL0v3pGIoGE+wUG/+eoXpueOjSxjfsgo3CoaVXmHrnOORBC0
om8RXw7jV45tCinQlgdn0Q7UBp+vT2/N824DaE2hSY1QzlmGTgldf46Ii6H6Hlt+
XJoTNRjgKqF14hVmKCw3ewzVOc4Hlgw72mxDfrKcrJaMY/kJsCVCrB5PF4nSUYGF
f2zfaicRmbAU+Ic3BdzM75Lnh6xoDxM4PkR+Nhh2N9qTVetMHga5CtZ2oYOGmhhZ
v2wU/kGsGFACdhuaaCoSeOfH4MSTJWpHleWuUnlbQ1cDpqvYsI4okZsp7BWXHw6O
6PqZzr4ysTRRIrLaVxanX94ADTZJEN0Bmf7hUHaROlPrm/56AnF6O7wVI7BY/1KK
82mjLSpxmgvjHYsSXpxxePMnytGWryaV9a6qe8SradnruccVNiIOc5Z4JlVepYpb
ppnciUa6J8vhmspAhhgh1X30AEXvTEKnkiMeIAA9Cw5fMW1r7EmzyWwxeMJDiABr
L3JX6qvmYmmoPYYh5OZ7lKsGj8rHfKB+/VZUztMS6zEcG0hpnCcV8qPWSiEHgP44
cT5H8KAbTkAss5gR4dJ5EHE3bFExBwc6JqlQ2DmW36PtYwqhJ8QRWIOEkLBE5X+K
XxyTLLYbMNgC8+w27XqVNSUVaJBQobNbmhfxJMRqZMR1kwebzS5xx0vI21+cS/9g
WmZwLe/8YfkWmlNFUrY3B+VOm3GYjX+Vphx+dmV9e457UN0hAGn9fZugksCUpyNh
ntxehurPUxZr8/2j8gwzWcSas0TbT3eLnBD+PF0018C83sKlg3DKObUqpbK66DXN
oZmkCft/xgAlUgPI/iKdxC4717UH3kuaiTIjeYPcLar9U112R/i6TUkwE7wKUygc
914yzpbLlKhsnFp8cxCn2jVam4PPto9FHNRo9Sf/Kkp08p8QrhrHEe65lxUTHfcf
xY+K/IWy2oC2o4qDKwGBnOoVITxOvqTgwJfGmjY1S20x7SCN8NchteTtXuhyRw2U
P/0VCYDma6n1xuIxzQ89PUwrW6FLtqWpmAfhdLVRJ1VuW323ave9g/d+mTQtreHO
MFfwxVd1B2QD9aTNve1dFQdlYTI7TovxM5g5xMXh9wC8NuWoNnGNrbAgfMY0DpBe
GNicJDe3SPXq0GAXzMrN1QkZ+rfXk85YHz/g01sFZ0tkaiZ8+GZHGBUNcB9MaxUC
aYeDSqfAFitkdY/rLUHt5sRlS2C4XSj2yYt+5mIyH9+Lfp7alBlDPOCIZmfaEikl
1mM/YMEQH2HdwkJ8KFH1jp2g445jf3V6/GBOABLXktF7ma15tXYPUNHOStQTg6FO
NKUbmequ6FDwqSz6Z75KVuNFBX7zrQjEu08/5D6sJI38ZPJ9pioAEgadbH9PaLWo
Zp9UCiLg46qPIA43h130D11ZcVaJTqmjsEZKLVZEMMtUYrFLMMe8VQT2Zs7aA1KB
/GIHcZNE3BU8hu5OfcPSau11uWy/CIR8gfeq76bvU0ZOwYuH4WQe9S5t7B81Zcm+
VyZSX2GwyZd8K7DLQZ9B1R5CiTi+exdMBZf6h/C5b3+oZMUnWc+e+og529zOLGW2
EEYe5ap50TViA/e05Vwuv8QwKJg4LoRRJ9XyK3dqvHN4uMC2Kg8/xtWOrlOKkCju
sqNQUz294KaVuTdUrp3/zCOLPr7KHYxCiGuFbjOITFUUjvijOJIITzujt9TOHaac
o4yFDCjPl4hT9DodgsK6+n6ywxjiOkCEYmfmVvOGYRP17XRwWcqQ1ISYGgyZ7gbK
QSW9IVX0x1xaiC3Jzdz2mnBc+ajssB8u2PUuMc6xcWkJsnIuPRPV1A/1MfVKQSdO
28AGDmuSns6sggr5QWcNj7bzwN82QneBxpFEYqyxyDEnnMxMHvqC+KE3dp2gyjuj
dao3cK4NKmcMW/FxRvCveQDi7LtUMZnJoY+q3hKnSzEpItkBn8euTfacaIJCVzAb
dl5yzdCTtlzoll4GXlR1e/8rv/xvG3h/xl9x4XcTq1b5k62SmI/y0tvTh2oXdZEX
R33BEgtNsnigRzLp/HiTqFu8cwRNByVYC+P2hWRK+7iJQWD32w3WqnpBqxduPF2l
2PUHOhzclhGJAlRmqhMz0YJDaFhpEKdVQBICgVcVzw1SSsSPMunxd2J5vy0i1V/y
VhtUfcA1BkjeUGafawWohCpnViCreHWExk+nD3sWJzYmPEAHXt0Y5fOEdaPivfzr
62Z0jICAd57jMwaRIRnQQX1ubYEjgVl2tVcNCLJDn6TIrQFRoqcqSOhg0gjhcGD0
6tNWGWy24Oerj8OuSr9rKJuMQxAXwemcvFyT9Gf+cozGBSBeUUVEXXGDF/NMFatv
3ZcYLC/nqhfvVVgCRVJO6IAb9rr+kSq0knxyY9Z77brAREVl60mconKYVsPl1Wpo
vy7OHueAZGyG0oR159is9nQ+3MQi8QI4encZmlWxhnd5bKUcsrgQB5Wel0SeFW2f
IMeWMexknW6wt6tIrBujI77peXNgbSjdOtTFLZRc1yqlK+ffhLhq5WoykO9MShHB
gEhhFYxsjLtakDDRyUhi3qj3xD04NvKtHU1RKGtkfu5DWXVfNCR5yu0YR/oRSMoq
kv5x81oVPzH79J4Nsr5PoJAWeeJvMUyWdfCTIUz7PqEV0dAHRJhnppK6cVYIhV3y
EG1FycLL5Pr2byaKnkcbKm+DIawPimGb5QjQEwgzXIP6435it54q7oMESQxIiqwm
4pt/3TXAWn4lBnE8WpegqTplUzovgD39mYqBvDaCwEWscfaCHsEqEF+j8UFYEBxC
ZMC5H03Bf/2l8ONY0FL/IPBUtMmjPv231nx2YJb/8WjTasWnMOxdMKv4XwB0hIuL
IXtlgTZWJeE8r+4t6JzmuNHXAleQFfBiORiImUlQdT/9f6QZp4YPCy1GhfNGYhnc
1xo86+ctDB3T1eF9W2fYBPC0ryMznudoUrKP1fZr53P17FCTVb1KSyVbjwfLeCNa
6fEmR3Fpl8rOaMnL70Q4ZKLtoqzOn8wbAeLoIU1yirrqPlo+uf4IXpQoIEmGSRui
XjVAZ6WyXWnOab3mHjmNfAemuUIcBZlMczIzyKbSp6rWW+h63TmdC5YkVSzVwbO/
2m8A/ZpoIunzHvgIvOXiGc7z6Eo+d5VUdvF8R13yWeIT88SDSuyOVUQqg5qsAHO9
VPzwahyHsfvhkhpoONWMJOeJb9T+FYEbIe+vSrV2gngKyXBRMNF9bs9KL7ql2iC0
WoM9QIZ6AWpvbpclDrBIQt6aGQZ2M9SU8XQnrp0naIsoru+8S8+8pHwDE6b7nQB2
o/jQQzZlSNguCDBtaYuUBzHcMRGRXoTq9hFBhOBcC//H4K4ImWGl0HZnRviwAqG1
Y/svJz6KJ6HSEv9yPJWaniF84avG/poWOEjUkNVHxDsXdxWisGVlfJFT92vx2g7E
u3y85+3FSYyzZl5OXKAt7ijLMkoc39apEO8u/T91n4ny7tETsyKPmImK9yMqE5fl
DQIR69c7ISjEZLXvGE5IKH9efIxwQifHL9qUI49X9jyGRGXk2YmePJqOC9ysXcIL
l6wRA6MQ/209+Sleh/L0ay0o9JEa9SGkoQ37L0EdYSc6BkGFlTf/zt4NXYWyOdO/
atZCzi7JRf5tFc9LFbkR6j6urYfY6CwvruPiWEZ8vkNDepZKRxSY6DY8wDUSrYIl
6HE3eBV3wF+mDeqmv8IJtuz/LqoGvwyY24HX3dGpmKqU80JdDlTfM/MovDJCwQcO
chyT9edn4IxL86/rFid9qgzwDQ8cI4RZKCthQFiecG/pZjyZHlPrkZvmk+8G9X0W
N35a2Tp8sgNkyMPDWAp6VXjYvRGU2uTpihcaBZo5sUZN+w6/8P3H2drd+9NPGy2A
jT/t/bB2jNxwv727g6nS0hSKip4Cv03t6XaFB/eSOcAQjmjxX2v/TPgafT2UrjVm
+49HGj+BsTL7G0aZAgMXUHrsXb4E7ic7PlFz8tPU9qQSvYFX0/B8T9FVKoRnhZpG
zFLACI0nj1sLj9GXNbJaHDCBTr42ppJOEYZ3WCkjKHaKUGYR/hyNrV0ICjGDjlj9
tXA5wD+B+zFVKMVurMjJNMnSShc6kxG5qZrV4WwlqtV+OjPpjc7uMgx+u0Vja7ei
srJ2m0nfd9ANU1oHjaDfGDPRqZfEayWEKptA6XwZ64APrkHdjrG6rzyRDdZyny0y
L60l0qWPIfi/Fad5RS2PLuR3yXifFVgqiFKyHzCkrZJJfeB6kgzgst0Fe0rono5Y
4WJOb2jKtMXoiUddydgKFL7mRLyS0jIhaeqpfrQl4ynx5H7zs2Kcy5kCiHypbbL6
lsP+DTzaLC48WH2O4cxZjgjz47boNeJ6LOC+arwhe59lHXV/+9ULCwYQ4FDeJ0Ea
BEoYid46T3UHqmOo+3t2DUC4J8aV5EXpO74Fct0+uDxQApvcm4UlrQyiUAqnwKTV
8PCqVN6GhhTrolGo6YOFWbGzw1qw2UxYTW9Fnrji6cS1i+OhoeYr2kCit2klCnrZ
anHQf6wc9vB/fhgcR51K+vnIVQGS+E+nX8RX8GRKpJ5xchmioHNNtrItmnlQ1JGU
s/t5XjMILrnnCUfQ6dYCJeE/L/ezZM++tkdoz6kvMcf+ik+6tCOIcgf1+WByEdCD
8fkI2obNbwj0ju7elgQ/OUMso05rspfYi1BZNzwqq0XeXW3w9F3QJQLAAKB5idFZ
s3aVP5X8OX9jx9v1f+4U77vYE64hbJn1oEqiRB9V8k/hXJ6p0XCICMrbrxwN94AV
yylf81rlf4J2PNzQwKwxYfYZZGGYQ0rd8/5BgLQFEOQ8fmb1KMy2kOsgHeStmErg
7nrKUaPFAYA2S9nOEeseUvGkQkpPb51tIGDnO86PxtyGoJ0ifd9Vdns6lh0dzoLc
Z+Y0E3yNdJyKERFSa+QMab1zNH9/HZr/8IVfbMA//43/v4EhkHKuYwRZrN2mEe5f
BLuhTdmfQvh/20byyRb8aivDsCYa4/1AKmi7IrHdQn2afHUaZu38VIgDrmv0Qgvz
RFAZstjWt/PbXg3flr8fbEWAFiHxMn1362vROlENL+uAxSS0qVblllRIS0KMbc2L
a8l0hsKIR49VHX11zzM5c7iJibXAndFg40KHkJr52W9xM05vk6oxiYxHbPeKF1yD
Hy1zoKGzRD1ZiQgV6BqPGTvkUiEsFCnLBJvcChIBUF3lk3kCGsjj1CqwIV2NPt8o
716oCLRPIQGT1GwoRdlo9xcC4p2pog/EQWNnGjdvwso5NnEf8h8fCw8Sv3gKu4xm
xBe0E5DrNlmuRD7YoMi4Of/CWqkPCVE2s+Jxc0wXVHKFG7mjj+6MvDXH1i9sjGu7
JYua9pvc/Kri+ZXRrfe3EjNbGUQ5OJX/0gWv6QnWgxjP3nQdx7DWyQ1UnJMP9hiQ
T3lbYJT1odP2D/6v9UltIQtrVu4Nmo7Ke0PIdDfZkTTevpehO32jsjz0rjzdUicF
dMWg6HQbijZzkdMjHWiZT92EHePdYwlLuBqHgOVDTzgGgdjcpdDEqzgKt9UBQsbu
prY7Sp2wKmp2qUaWeTGg4qXdl+MM+zdo4Fl0iwuKub04nlbDVA59JqHxEwq1c7fg
KWjMFtKbBmmuqWWI+6oE77JlviV0SlA35qcU6qrxXGlbyk6OSqHaIKL0cE2Pbsif
U4GgBq09kLDQ2U0PLw2phFYkRJmzmPQ0u/XUo7q2XlanIBKJrtPtOMYHK2FG7/rz
lmDlGfDhRwUtJWGJsmP2UuYemhwt1T4pytLoc/bbPXziBN3m3sF0YuEarps2UO4S
ftCjeGpQk93xSXD6maE0lGyVZluWg7+6m6QUwks3VZY93WkuJoRKlckrylyDEfso
svwcEbO7EEf8h2pV5M74ScYZFmSd5xHg7xO/MOj0cxt2apsEY4+9H/RsAGhpSmFV
foa1brdDVzByBQDfEXdUpcNXmHiffqoF0UPZ+rOPK1C9YxgopQAh8GoxLQKjkkz9
lDIcnWGX5Ut42+A5xLUxVigoKxvYG1HyA3v2pgRGNw5JHMgBxiLicw1u8WH7U1q8
r58dMZqcQpeJeZA5pWw4j29+0yAbn+f2RwmQqi3OsZFOBXf2vcB4Ei52TGvTGLdi
vw0W6W2P+tE7GMNgXzlM27+Ts0sAkEI7gPbofXc7bf4K4LD6VaWni1XPtKMFg2g5
Yan48fAsP/mjL2RJ0x0ajMS91Kp+q8dt0mcAEZKIiX8t98hW3x/qWHoZXHgRkzsn
V/Jj8qlmR85MA9zB+I3+nRhm64TWt4Gz2qaVPBzbsZSVME8gQESvhpX1k1bEqT9L
qXCNs+uVMXwNOnjcW6g7UbPxTH6WwR0y2Aw9h4zmbWn8t84ZjKnJj/vZFJb5IgUS
HrZUoqyatCg39gGy7f3NkdIkXIMvKnvT87exLw/uafkBnD4WPfpZZgn48mYahYvW
i0ieqOWRw8puRgqxPrw/5yp63F03cbQwL2CB01jnyBzR1V7iObVxX654LZZeloie
B4ZjU8QqW4Ftbms6/E7gDuENQ6JzPhKtGQGesgEl5NKct6/CpXC+HxeObVZbfSpO
8fdxIPhGd1DJ0y7gm8leD7h/lmjzDv7Azw5z5Votopcmwsjx2+PWDs5+q6vmxXR6
K8EDyWQoejizhbYZeFpDJVF8Qw6tv7nd/l4UY7YYQcvEegjn0U5h93oxkUge627H
FCNG6PnZ30PQ//W7TE7237Lr0Dt6ngRPDB4CBmNAIxlrsSRiXwrh13v9qo6zXjWP
vjRBsfnGvi/2o3hJQ8K+ElTaba76L3MMXK+0GoGYA03EsZTqKgnRaytBt2BbfCps
rTDW0goLkVNO+QgCCJuTqWoNFh1E2eTmReTiO00lm7K0v0CHGGJVCZ8H+nJJk6iB
vuxVGgiZ5FsGmOF9eSPtuifHj3DGn/fTDQH7KXkWwhdwUFaIIpbvS2Xn3A6Fnafj
VD+WoXWtEyBYr/Rlga9YRp/3J9VPW5KJ6OKL636ouWjmbU5o05K6qZocE/UzUalY
3escI3urUS0QZJ/EG3aFUK7OSeaYgRIOURmE5mhnJ0WDuQjuuxaUwZan8mtxfBqm
P0ufxdemJg9vsaVQH7fqX7hb+cVBTPwysa6hkClGlpQK+N7cyZcgu8BqXvaftntM
SX9koaLmJjEKa+lg0Wp+maSsZqQTeXTYvwEwcMrB2HQU2QdwOJzzdNR6+H+ZKlXN
0ra22nGotO80dKqWxPDLzr0QCNmf7Tmbbfv2+10+P0VMlU7hPefmxebZK2ENFuXB
I1PxZ2gjbVIgzMqXegYEA60iYgZdIpkQ1eAWsNeAcVZi5K2N82v07Fbi82V4QMNV
UAREt450zx/pHrQnG8IXsVVsneF9u3thw5iZI242ow07NTKUu8LBWcI9jamXW8V6
japoa2M3e1iMherr6UT3hgKZcJcNv47e5MdCIircMNBLWrbkaCtkNw3zY/oYbGF3
IWtR3o/StyUn2tFUd6uGKIfFM6b5c8QkGczHhdiA/BP08a88+ATKSOSsTDkYZovy
kDIKf3EZMuBULTwCS2tCZcxuVFSqexQ+lhcYmu7CrV7oY/X+h7rebFOTSv4+sUae
jDrwfaSuBZnKozB2CFY3oah3OGCTw95YVx/jolEvHV6AhNacrdkxLgBb5ttsyQV7
xujKKbiSh8X8QuPzJACjmC7t2G7sc9WjzAcLBYYoXmuYiYT+HsjOq/2v2bMjitl5
a9CpiPXsvR31MFxo3lGDQYY5oHvutB0hD1J5S3dxdMkwVAL64FkSgC7HCo8s9Dwu
W8Lx8jJcer/4wDeXIc2VGiy4375XJj9l0U11ZEOvz0/BQth8KU/8YJExaR0VFwZf
nHdoR5kAJJY2Fu/LkAU+waJoMPpyrbPlzxGO7LEb50yfEmWRqOy9Vw/UQ+b0SrGg
kHLyDQV65lS2c42A/7MdGq/lPCGBsIkhvhMI0iP5BYtE1wTe04Yd5xluFOxD5OTd
Gz/faFq6yFwoTccPLAnczcdPJlPajLdo8jHrknsIL2kz5ypMrpFbpTHUQ06xYPs4
uvkMuBvcDizjXlX+pweu+WDzJVs6nphLoHPd826fDNxOxXS/URdxZMc97O0dzgux
EWlBpCVxqA8zfhFb+E5dbJGght3wFERzmpLLSDSlHp3vAtXN6iuSwWSWCc9+Qp3T
odGbxfd3uz6MfHnSQGA+B/CyrBghVB1LWHqP60z1gpJndlSIjmKwoq4iJUuzDeD4
vcPSurfoFdvDrSTWtOHVVdVkPpvX4xFYgQ8oHQb1X3nBjbW+HKnDsAx0Ii8XwIUB
/FtSXl7sUnP38QM4b+TA8hxA77y7xwtIZTfy/Ep9ZjfHgtsB7JYJkKKbnwE4Pgl0
sGJQ/J1oezVwh623T8JcLFGJ5uCOSp3qvOX+5pYjKNSDbsF00U7LV3yP1w92krTl
Xdrf50GSP17MUHeckfvT/E8H2uACD4NqGS3nbhqFPK27ocCUtet19H0unfyvp1Kt
DEaWeBattwYcp4+4LG+CiyyX9OBvTHB6hxCRhNzpcI2nD3Ec2Plh1zKhlyETjcZ2
hylA+brdeLiPhcjJylmgPDY7zfUSXzFhF4YxF7gNq+On4y9+aVJySsMejuSDdBjj
JIQfXrOwRxOjlTK+oUnrqxoi1217xuByP610E6jb/Y16l/rciL8vAXHb6j17FrXM
jLpNH7MAcFrW3f/TCOUpzYXafzzkK8erJcmmb4vu3bGxAOkDZZRtrC4XrESgv9e5
OB0a16v9nSgyw98G/ItDNiUw2At0Iyu0s2ASx7se1icdq5x5obc25J5EnKvIv344
RBlU1h3vBG/QKDuqie1Aq5kCwEBYF/DN65rTAdYweaXePJjcaK9/i9drTdfUKwi9
Z9tL2jjo557fpRbLgoMTyUAvGcyNQgM/hrGkabsa+i8mPrdZrwPZRWBmDGH2mW0A
uibeUYhfjb9Sv7uRHZu8cPc+3vnOpdBsAY2Vjd3h6uAUkz/bmfeTkyEo7rJkrXIl
n8ioQSTTJCZmDK+dPvnvraggPNI2Qbs8tQYYNcVSVDhqxLyiaHk6JXm6avHOQj8/
PF1IKjSElwL1y6m2SjLXnRfpzx6+Y1mV38eQztt0UtrBUdjc1ximKIXn8yYww8Cd
v+Ypg0vDsmdYRPdlHpN8ds+fWQlMySp2l72hHnAPD0W0tZ6YpEY5OBblUEUSxTug
CzrJxhTdI9L5XHWeg1TgJNoDPVC+CiT3CVgCFzIWsAlPIdwuV2rjhBZoC4f6omz7
ywyKsyt/aHofegG/2uVoxJviha6liLH5/ffMSb1ohuNueeN3mBuq0stQpVrZO9Wd
Z+xWqHm/2DsOci4ckMYS2Pl4mySAMWM8xdcBm6TNU0IKF82FQJ3eR0Zz8x8x3ss3
38X/KDT8/7T9bBjke2+yMdVpnZ5s1jCeZOqPheNkhZCuM1iIERbviTztVFMHHxAZ
imdhSfRayu6VExqLZcQGdbIXgXDnfgSNUN24W1s1wJIsR6fwDrBU0lGkRnCG6Xzl
RB388qyWFxl61y2sUamDHddNWvzFzJAam/JA3zUVAQhagyNPFqO70X96BoJyvM8v
VZwsgr/b1SD3eCxiZwJLZqFartwO2wjyn2hVcE6eC6XU6YsQL6VpPgwNk763NJVc
NOUMNbOyEc7pejukPsYzHzogLYOOUwZEEAgQKx1anX98/MGB8ajbhAlC6KDJ5zby
ZVrTEaoZ8YgtZEac7DTAQcBNmvRBHx8bidgZX2sbWw26L12guYAlIl2tdwITb2xh
eSOe2O94YwzPzhj6hxBXngFI6enav+KL3emXZ6kSDxra9N79MT35SWEAz7WmocPX
45Sh+1xzb3p6iemlrshJQ10u2hcohb2oIQF0/P1GDS4D4IRk4wW1R7A3Np+NzFjV
o65/uLcihI6Xyw103WevpvF3/iLqnoNrES0j7kcbc4CuujWmEb00IvlAAHP7hyPJ
898FZMr5x4mKhVNHwlIXSpCk/oiEokq16a47Ud+dUrXOsAezosCvukTD+BxUIW4y
97msYdrfOxgraYCt103KxF0Hcw2HoiBoG0Mrs7BRAPwCYlO/zW/Mzr/TWazfLWKc
Qe+qz9G5XhE3pj7dTzLaLim02ieeOaJs0NpCAgy70ow+8QB3HjvNjST4iHL7dxey
LZaS0uO8XCBTj3Xu+58/vYW578ka8r1OxkWNFVnJQBFVbe0K6Yw5U6VsrVjqNOz7
CJbqkbCBY5zzApsfJSlUzgN1nI/mqnJGgLSI+E2xBucQO0qG1Ff+TG1wrnUApcro
pGo3ycWT5kTURAQd+3Bw5q8HMrPXOeCmpDjNwXZUi0ro5WCdTLgt0lJwXYXtKzZk
xUyym23hUa240rwaZWGc4Ha5fKmzKQzTPw6/fCXSV2+kz7lavoNnHdcGyGf3H0so
hu49Joxx+HF1KZ1G3GYHoIy0OPR1O7w/VZrUMK3nQU2OmcTk7vxRsrytUAvzm5N/
8Aawc9oXYoz7yvmNRKG4eoa64NdPN2N80gqpDxwRNn2hJBukAMACOzAluV3AOcQi
7EBord+/LAdn06s7N9amRe3YX1EJaSv8XMxgujEo8qGpk41C6vkRena5V48Xn9gA
ZtZmeOuh1sWO6lUtWYujEJEo3pqkMuxpPMb0kdTrPvOPt1KhjI8sjl2925iv6Dit
+4eXx+6EqVI6fvdWYUoxpzt/UBo5GRrjI7foh869fOExdVs90Sin/n0ZqpRArYDl
aVq52lsUURvd0qWyrSkZZs/N6H56Se91wF2zrfLj4f2ABkC7nSC6gxCEXzXuswTQ
EnTgSCejtWiP6YsZLIGYJ+xAPtfT/oKp1Cl0p3H3dlzF3IJyAGsgnvXy+ixHyVkh
HkySdgFLaE60UmYkFNJGVo2Ppxu+UQlPfixxrRdAbvrRi5JBBv/SG1Ol18LcqDLe
170Yt3NBDTr4yXAxUKysjEslnU3sn1ZsVNZJ7Mgf2RAWkE38GvCiYAN/ATaRqRSi
mxJSxahmhf+QSu8bNChMcpohrATC1aOZ/NZRGFEKsFBv2mHROyi372o3Gc22CgEf
56SJGz7Sp0nKIzXbxa9U1WXgnNvevLnxiP+6SK/YwQY1L1NFdTT0vmxYgUCWEJc9
C/4Mqp6KhY0d1Tw94spjQ4vRhDF/HS6b6Ce52OqQ+FoKFxbxZo/VlIKjOHo4MPsh
iqrQYR300AGP6fVlYChCOocgn5m2DbAJU64Et8/0lYXpVBPwRV/VhM8Yav7Pvt+G
a1SRKptRAR7tQfnGp4fPoRpCGyVnPsLB7g2o+qgQH88tYMZ2crO+XobL8/g6ZChQ
lbYFmo1dILLVLcYdXuos0uXAoOMDPrIyRhw1nZ6pQwvDl3Ssxh5O8Tm5XrEEasZA
9eKL813++vqpHxkavxaoYdXOtwW8YoeA+hnCteQSRX6xuoTFXLwPfBPehhMjDGW4
Jvl57gq79JgZPs/L+/qq+wgN2fAja1qp9lrdI4CrKl7YwBn2Jy9PHGed75fwb03w
pJCdSwfc5cBdUNhfNvfRhj8yNcPy3OQcuKw/saRRKjgvxW+fOj4SkLHKbmShubhP
i30/37/7PSPNhE4seuW8YvuqGsYnQEpohBSXSaS97Z/JLXk7rGgMB3ovYHZqRsng
yt+aIss3LcMC1WY5rOVAh0nmMQ5428PajjiegVG2uC1KI9jarXh3fL6AEte6i6KJ
UGoWEgRPpoKHgj6iAOwlP8rCuT2za/0zUs670KiELe71r3INtIKuW3CUL3Cam4pA
PG5sCPTA0woIPfT96FbdlaBTkFsMIH1ivcxLEWGmml9ikdgZSsS03inZ6OIhdtKs
Acj2iGrfY+AalbtS+nunfwOFMChZ0pltTh5dTzWrgRURnDE7gW2xK5utqdaer1YP
kX0pQ6Zm6p7RhVCw8mofuj8ZAM8Iry7dX//Zo3E2WrFR4jLr5sB40OYKKEJkmgkz
o/4mbxtFhUwznN9WIX7u+PKsUjLA/IOOXj6z/Tqw6AKyrYqIq3rpg7gyABke2ei1
hAOH4u8yroDsiIGpksBZvkhPM2aRowgvJA0FxVD9l3bqstG0DLU+h/FdgCOLkvDf
kIVX/Pm1V1dBDMhH+KP8chcHMF3yYpzc5fTffl+oo6HHrxgZ4+YSqXB65Kdox/Kv
67Jr93DY9fExbiBrh8xKO7LxE7EfDWyCdDMzzR9tNkOU7++qvv7z+XzDi9aJn/+k
u2NNltxYiUyIUvEP6IROP1a/9cCYcgJ+KNw+q1phXozXaR6kpdT4fNOOqX7CWQ7d
vRZSxNZGXxlaHjjRKsyu0Ilvnfu0kmvRx3PbxeB8VHIT/SVdTCTnhmAVToCWgORT
7AD2AKwtLsn/1rAEaQfsCTi/CdNL08u/lWb5FdAjR+DD5sSOi64DjVbCHmLmZ5fP
R3L+3cG7thErNyoVO3bumGMFyemMimodV+Cb6sP+gRyPhH3Lt/34gzvCjD5MGrwv
9WuO0H0ef6wi/nZnobpm2J92ueO4S0HPjyOQ3STxX1/AXMcfhpeiQLxCJ3n5nv/k
s2Ghr9yHqaG5w7b+QisYSYUVfKNFNfWac1Q2AV2r1AE5juv5xF/dGMDIXDtPrmgd
Txs8lFC1S2RW95MMZ5AMc6zojRJEtJGbZYYZ5krFtkzhDK7gvNvvAjbFGdidESFx
54C1ticmy13DBELAMleIIlmtstqdE4U0TzfznB0VvlrRkFviYdLOgfc3g+GgKtL7
QniagK3IBGJDOxbAHNHkEGKWZ2gvahHla1QITt1GY3NOtr8nSkWDEI3XAym4gJe9
bTUP1SWL/H+UQrQsX/w8839/BMAHvm2JsvUZW1PLn0C0Oo/Yk8ZTP1ZU1P2Qwonl
+JiGRvhxN4kVV69vNVi4oJG5HxsdaHQBvQxjgc+y+wb1vJCNB+vH+5XraM6pEDjH
2vGQe4+x4AaM0e5KpbAVhO0rBEV1JUHr+sB5FYW20UKmddFrKhFlLsAqO2D746LN
n5kDyyvSg3LJWXcWPdjz4l2JEvs9cb3M6PQ2dQU4bpVDROGmm441Sd+GmcMiimdp
v+NPTQK8u3kR8Ms8kFUaqQnrZplCRU4MCzJASTwRoo+R9+kWC4xwtpXOORr1Mitg
gXLXDTC4kWDTK/R2ECCvWwO6zY2P00iJal2C+U+gR6yRbc3/E0KiKoedpBWNF5RR
lftTd3eYdmQueES9lvauIcaoKJOqdxffrj3oMDuLNvJTJGLaWCPYWNLlbfdIMlTA
Af7lxwVYGM85MRHq/HBdHye3NhwPpLkdop6YxzTJ1bVGNsGV8B4O97iybTfCU0xJ
OCkO0ogl0wN31cOhQMwHzSfpdSCjhDn3KCvYhcu7KtR1s/Bz32fM/YYSw+IMEq3l
FVrfDBaBZYvLIxib5oW68wepyh92FhPYQzkZnG/itOd4o1c1zooSkHIlA54zrvth
nH3XW01WP+1PwTKtrldzH/kGVPVKkhxG8SUauHe12sJY2bocF4TQ9Kge6qcDXqd7
oXUbaIFzEfNA+gz5CZRbs6ia1YeQSsFssS9RMYlh2LGjl/hkWopU/hkwMvaiobEN
+u7mD3KThZTfYt3/tB0HeLsl5PWHasbDka5CbOrE5BikYUdYWb+oA/qDzQEW1hPO
NB/IMaEYGP6jcVGOTdmo3VxzF/ywHM3gE5lv3BoPB5b/dxzL1EIe1xY7TF3TJQ/r
f4ceEN9Y8mQZ561R0dffLaMiAhyYTfnCo8XcWGXItJwtfgpMgnxVX3At7mxqhB5a
/kFdz1ossvbkjB4ZZghhhBYkj51egYm/M4LEeGApmALR4uaaSUkVz5cht6chAaXV
hPN4GrrxNiPKEf1bF0sOoAcYwLyvbvAX1835+4QhmVwhpRpTMhzlykIaAB0emgL5
ADA4oFtrlF9GI8N+RnCa1Kg5enFsoRcM+AfMCHtG/edjzlZsw60dpiy6g7kp2URl
N7iEodhs4e8V8SfDfGPkZEhotPkreHeNR2CrewhB5v8heX1ETSB7j4BqjPpTnmgn
3OCubGzn+EUtTMDVwYpFyv+VaZPqt8DiBWRqSo7oBsv+yXfxF7oK4QCLWwC4gTuu
wa8vSLAVv817fwJlF3TKfQkskYJjaqm7TUeHroEF+C1lupsgNaVWqsKrrrKWyaaz
hA/Icg/xuXlhzUZwO+A3byl/pZLddK7OnEZJhocKdinC5iKMKMi9RkguidsREGJ8
KhB/eH1CZh+xBiyjIHGmpf7n2+O1U2fBBEXSEd+EwbesfXEavmMJLzTZxq9ILL8s
0UMh928xjM984pZpyF3/spvIt0C1JHiIAKifrQBwN/oEhINZfDDzvZuBR5WF1PDH
qdpM7pH0PpIQKALtNPRsdDL2WKI2+C7UNF4D46bLpB5M972pkKjvCi9AzCaOIpIN
m8wWU05LjOraORlwN+cBIuvrniknYRK6Io9mDTqyceJ+s7xInZXJzBZjohcjQjjY
eaKxwDyQmRMFHaaq5Ym/j2T2avDdl/q09m3SRSq38Rg3a7Z153wD8pMIkIp66bGC
2SMQ25EN3aLgvlppVY7qE5Je3UAz2OV+riAA1NqmUzgP8lJJTQfdvvHCzAX/Xmaq
sTpZKP31Z3X1dyabadfhiZbkZ4gHBu6pZX9PTCpc2+ERiwJHSXCMQPkWD2I06Gr2
FN9twKdi7BC+U87+qKGbMCHU2fyJivXmYYxdYmdjYbpv8EZSFIg652/9Kru7+USO
6OYgx3pcS3+avAX2vGZ7dPBz6T8QzKGveaPgHoeb6HYpLTaon5VRSaM2tQrMWmos
e11rYUgrxj5UMepHSA0srpcUdezjVTjIzmySo4G3jSNKPtcvZlAWoetth16wUlSZ
e6y82+LL5VtvyJQVhZzs683yP3ZCIlUcx/T4V+MJbPT/i7Nq5wIitXCiLkug23dR
UTUg/svARaACnH8hfExLiS0aen4t6+JoJefn/nIoToIOFZLifhqqPDuTE5fTGKoN
FlGCPeE0mny6bQmt6HgoAddQHKNxzLl/bMHOhX6Gv28Dtd/dDt4eD7Ux/ihkHsWs
PFJu/PtR9B27OD4wyjYJgYkTBu1QXOafwCkTDc254Je/eBh91ODwZsLaf8oPfVt+
xTsma+KHPvocgtwaXRajsawewGdy05CvGSEA2ULHjRrTHVbB6dG8WAVpEBKOlgnR
XkbG31+ZrzIR9BVjzOtaJv9rQ+HGI8gkAv9GXHCjYZXpd0hjM+PhUTQPvv/5ebho
tmhihrygUCDW5JpvnrefUHZ5M/BXc7oKhVhlA1HhENIb0ywnAf9NjTc2RbWLkQix
3f/vrro/MhBxtyzHvziwySuuqrHi/P8KsCGe9DvOIh8t8vlnZeDIZlGMO3uRGUCj
9fN2USlgRsZ7cre8WaJS5patCAnElA+T2bPLUCIIPTuJ9r8BxMfUmTDR6XyVxZTI
dscRQ5s4/z75rcEYnVx1PXiio5MEl1nAvd4sYAGv+BkhKA+K47X0SN6yKIs3w7/c
L5cG8gJ9HbITtMYgdm/GRX1kt8KzI8292R0+j2BGZh3Aq2egAkQjBrUoR4U98HMJ
DiLQCaotDoVzOoGA0HU7OzgpXScJ0U981NmumxrAokXTZPQKvuKo4xg+fZJdJYvn
cdRtE0d8HI1QcjpXVpVDZW11x+J4iKEFH66hcFNaXXTc5CjHXmb6VuibLRxlfXsJ
YMUlNA/kUZH8Zyf3E7HStoDCDzbqzYYUc/hSGI8Y1Ds51XLXA2LtERJ6m2E61crq
280R5q0qFGHMu4AOWjA4FysYrV3tyUHWnIfVHJmBJJbo9Hp5bY+5g0kXSyq/OvGq
3MRk8+yjjKF9tRR/wobTwjC1PYBcreJfm8NPJ+mXM8yfnPDntA5jLqw5jGYrW/oL
Vactbzd0jCIjcSKt1+l2DUPKM1cI9OB2/EsIaImBO8tHVHbpf0EzlfkX8x20tV9D
ss8AcXdh0YHJpGdHgOJL9nlR+AVI47xVUIwkQ09ZB+tf9aoPIU1BGnWodfL5OPed
gwvvSR58vs2Q0GTE1G2S8g4SBujifp4ELH1g4nLpRtDzjutYI8d8sIbeKIc4bGT4
y25UAOwHi5kUFYf8cov6t741JTdQQmDyoRjW6Emxh3O/QjXpuBax/mkSeZaa+g2D
KJms6DeeMYymihMSg9xpmf+wwy2o3Sgd1rnS+ebk6obo4i9u5j3z9z5A86FfM6gj
ObCOSWaop3L7QLcr1H7VZla9wUqpF8wdmwF//5dUtOBt19eNda+Pd5LFaaADs8t7
FfDmbkd68aCN3MAyHAlUltZ4ZqFlyeCsK7pIAmiJMzOZBq/GYKK/h9e/MkbQfmac
nIm/q+o+KuyAR4ERw+GYgAc1zJtQmsVQfitIfWf4s8unuR5KEqTcKE1ivYfoSTPz
r4Ya5/N7GKi5Q9M9f3tEaS4H+5QqeF0XBf0hnc5tKEDQhULW/rnOvp655NK3ynda
p4cp7npVJYOhg1NIlFznvLyugRtBn5psSjJBaVFrMUvsdtGSxWeS/0ujQvNLNl+t
LSXJo8/bNuz9gHRvRMdjHMKpl/2EZ6pEhQgaWCILwO7nQ4k2Df6GGKOpoVfR2qkc
ZqgoTsBQxoXNuzlI+n03wms3CUdLm4tq1tT0VrgnAJM+vEsA/fkGOd2BJi8X+Blb
x9yML0hRYyn7+AINHojQHHRhKptLMjRQ3XQeWbS4ab1R7sLoUUHBIVzGGj4kgi5x
nSqNy2T3E3d2IZ23K/WVv3jW5dvBdaIjyrX9WPywDIpruz9D7w68pisDQy0RgmOw
H/bt8LCqoeG/RxtTvZqBZjxXY87kWFDWyUUeAVb88diG6kjl+uRKKzgNlYbn90/7
aPlVLTuYqAXSNShT+D7+MX+DQ+i67Ff8qVECOXN+8xS6sZ01ZwleVI1f8y+wk96r
KttD/jDLdG19FimA43KUXzht1ISSftH++QO0z56ap62/EJiMTOUa+maO+d44YQa3
Aw8dIdsp2kCDHesNjDLvLQPY3byg9uk95aW0sdVpNly7vGEnnHYJgMdPfgeCKzAh
GOljMDJjArelZC8yMv+eZ44/qAUdSRmIVLkMR9u3HK6WUplSe+HbkHm47VRxe3Qb
q7nRBK27C5c9ATmeqKJskTRp+sLAfbkZH28wsTC8YropK9td0+pRfEXtDBRZnsYW
Za4KM1TSG/k2T06b8uQKBnKHpsKkPojPhWfmPu3Qy5JkjnwtFjmZPiB5/mtCrUfg
qupdatUajvVS862uXL6ixbzAeTSgvaHfqLB+fck0/9mo8sWnL2Sty3EfKgJNgvV8
DMFTKI+ULuRpgBvGndx6aUWmhw54Cps3mz1rdnIA2gniGn+QfVe22XuwM9DuB2N8
33VrTZ5rlkimz+X/QUkGAcxPs7bs+dxgfELT8WotCYpMfB7fz4hLcArveYrUUukT
m1OtQMm6QFUud37lFA5Z9D1jE7QRzcXqi/lzgYog7pNEt69P7DF7sFoSnb7syW+y
mAWA/BDsYG4r2Xi0jjKuawQ7GlqNLRJZjdaXkXwA1gr/N6FkyTGshgF4ffANoZQ/
qlFbCKWu3n7MBpPbWZ2jvPD92jCpJko30f89bUgKZaNLLOU5xn41oLgt8IRltOLI
YJH0PG1hSbmWiuFY6tXh68BttQDN2G8R9Gy4+UN3G6uNFDi/+qnf0fAgZ17nqGK0
gobYbQxUIz2he/IXH8HXrP6rPwt9lauw3TZSIksWj977ddulNQ6vhFJgEl9sgFki
N8/LG3V0BPkxzZYe367STVz6UFNIl24dzjFcL31U8AFn2xhS89HJs5CdnOpXolpL
LimdTQIsDSx9hbe79Hm+Xvg/MNQ/CVDUbsNCKp9Rrdd4otwCOz2CrVs8j5nM5czV
D/OCL8nAX7GAIl2dtJ9MPw1d15WR6dq2HIQE1k6au2JVhy254OLLVwYFLWZA7vz6
7930WdOzcs5vNFCRapsdG184sHU9AOfe9J3J708Jw5T8Ctct2VV7qUoN8nmBOg6T
tXGtlr4v+OmREBPuiq4R1M218kv05e+PUubZtk4B5JPRoGGmQFCCUF0uQSIASAE1
cr9m8VfL10LHQRnHmLRLinYtAdBeeIcfM3oF/d/bfBRwAy8smeWGmTCK6csdUXRU
zEE4gXfDG80YWwQ+zcVRBgurV+i8QGN9DCLaB+yLq+zdR4K9yd3Ag+8x1Vemb4hu
9zZ0TmwSHGzidK5A3ZAJcIweenDar2GzxKXpVyF8k3m3Q1j2x7J+LmX2UADB+0Lm
Ye3rqlrgudDD4Iq56UcV2EaPyS+gspznBNksml+q9cpLkefHNgqP0zYb9HpTmz5W
47J7uwy9c4+B+2pOOUJPvxNwMN0saGMb5naBUFxrtec0wWlCB8scrlws+dr6TiMG
marjSkaBKoiHJBAdgPAygP/20mbVUYuhx3+RJlslCaGgosO9CbLyE4i1IIPhLJHZ
FJrXjJXf567np/OPLmKo8jdT+QzgLMN8Ca7DR1pJjXI5PdB1NM3vHJeqUEK0Soi9
jj0qUa9IPKhGBOSzGFWC6/X/ZTGNUNl9Pak3Fwh/13RRnPMmSRwYhYseox5yLin5
QqXHsFD7v8WqH8p2vDRYVTSFrmg8o0WSqmkz4ibsunbq8xQ34sHfJs5xd19v+9ol
p9aPeYrXHubUQPAecChZYnUUMG60OmtDbTSipc6Vp4tAsNyrIRx0Tjf58kW0veCQ
OrgLSJSgkHDF4XuruAuatEeS5rlhuDIE9dakDvcwj/FyoJPiXgOyaXB5xNcykwL5
uTEdK41CMAnfjBZUrQlWIi7IBubsUWpDGz3ZljJrX9+h0WPjmfrHN2vaVpuRN2am
pNdrpnAwt/DXw9QY91FiI/y6HMVqO1ZR7QtAjk83ctdIzBFc6y7PrqqkHvwMFTNK
UezyrPQUI9zaFgAeJCdgMC2j1Wma7A7eWBsycn2YQ9I50pDCO7wQCWoZ9D/SC/gM
6Bl/9Drymf2cBUi8mTa/CKCBgKgqF2B4Yxtc688UuViEes3aWpPQjN7i/JUoPuwO
z67zk8040tOhd3FEnrbX8v3DPLsxPUZ2seMyc0bv68zQi23puV05upkrTEPfVa26
ECFdLsGcd98t74ol6cRB8hcIiiFnUzHV8tR5Ck9XnnHrAJSVr1HLicyV+u5Nn2TW
QcdSznIGRYftGA2iFtLX6dtb5ILJaQ8/GJ6eYMkPKUozUC/gWRp0IErLPhRk2hnR
fXxkIgsczO/4GAJF9kZo0aExf5pifiGqZ/m1T94txZd3N4U684FnSn+o4Sp0jnhi
Kg7RqF1WYLwuTplJFxh6uSXtUMkDImhmdd38/Im4GVL+6syY0mX2VnGuf47wF2xL
l00ts7yW64BR99T5/ksGlkcbcl9h4uKZWsy2AXVvVe2UMcuu3bQyuQJtfhMZxWax
ojJCckrD4Pq0C3PhyXUjwkTcaM1P3XdoHFjoFjyYaOVS13d/yWXvfTcYDm6NMRd8
SM+1MWP/qDUmIjcOz6aMTtOq+EFPAuYP5t3m5hFPolyhHf/k9lzeDIjb40V/rcYH
wrvECoNK9QnOj220Jnxkl3u29/6gR90+OKoy996IEL22XGBepfw83WObvSbr5vYC
1T9Nb9AffGwXWYTGGU/+bKJ3vTqGoXNs/NLZIJIFajSaiHicf5mp+23n3gTs5L//
pF6WfIkFgkY/P+dwVbiyd49fvdNSeI5L17gdnoyqpIvAJRppiEhts7L8D1dZTa/t
DHGh7z/gOSEVrqJviyk1QoBewJpKIwd/QjvhNBGc14d/9Wks1Oce2KZ5o//qyXdq
VhH1Pq/fHjGJJ3STb75y3Vw+kutQedBotvUM8B/GxWr4cJe0S+MK66u+83SUc1sG
1GODW0BQ/+GaI41PGj00BVWl9SLd3YQogdDOxiSg98NahMsA7FbrbrWzAB5QP5rv
cZFRQPuY3N3K4PUMFSJWARQyN+UYIZLzakXPyviicSHhaSs2wDHIQqyqDI3CxSe/
YSxmpQywoHP8BT3iPHhvtjcbz+nqVVQ+4/QmjpHsz289RZqh/Tt4dnFbWWbwx3UW
TJjA/VqEITv0BTjeBKid5xzI0RgRPt0fOaQ3HGnOi7qlDDf0EmxfNN4G4In3JgQi
UBNlqUkp20/YYnGe7nOhr0cRb8yG2OBOE+Sddr/sKlFiSb/VbUDm3o1YJ7+M0t98
awzI/cEpSXd7RB2pBOYD+UYqH0X+TSHHccxzhGc/pBJUDurmcZ7FrjKRgfvGDrkt
V3n8IhZk0/Tstm1beXxp1RBlhNGcSisYHsg+aYvCkRRqGb3UGkqaNd/Wyg+LLGZ8
ymwvTBmVa5cHTbCjMgXzlkS2Zqp3KRTyVFhQZBMF5dYT6K2m+lQdtq/Aqzr2r1J6
gEL2Fr9F3XmY1wGGlIq2Co6etI0sp+7yEbZnWbqkfo1AN7BLWMeMVRHEN0U772Lq
tD0X4Yo9B/1CscE1fyyj+Pi2wUu+L07Wv0s+VG1Yr8NgZ/IgbrW3V9EIBHP9lCY+
LM6O7IQobioqriqGtOI4CBFbd8MZtU7zvgojGIf6QHJxOP6QuTmWet3373aoeHqn
S1o4C3cuGEH6lnC2B9KVvbDx3zSU+Qh7wVZU4mwi/VwJbCEjow+N49q+gPiDzB9Z
AMOhVUNuyz41EWLBQ8CZEUKSlg9ejIpbREDca5wb2p7tUB0RROdysxNZsny40VYU
me/IyrMzRCA24i0YjLGbW1BlW22WHfOJ/Xj7rNEdQ+7fw9nTfjKXc/DGBTVvctBb
UO6rrDpjW9ArDaAENy8toDgWKMDYrePRwTuukvarGxSdU/JV8/3s/G7O9qgbgO4/
F72mkWN7uGCCxR3KCa5D3ZCH01D6Sxt0OiVrYfNlx6pClN8A0oZeY2VhIHBudrIY
G5tt8/S6o1iCXuHgNGgtdKohL9oJ/uib08CzIgb/atfCPn4JrBJ1bI6zCBHQFaRH
sXVsDmOEwCqatqR/WNoCfRNHE8khzHETTS9WQvFFSdJy2mdpFss9mNsRbsSxAvvO
fa4dX+aI0e9DAxt0PPfRdidAu2seFgiCImqsV8jkIowLKtmQ6Ayyu2pnAU2lYmGu
RTmTvHk39jHxCTXq7BwdfJj+6bXtdiF2iGXAsv20GTBzRH1aDlYWteg2SP0TUqwO
jTUP/NQm2eaUdZtf+eEYziUcgJFHudvqJfBk4TWzI/1RtwUgENMD+aLFUa8wbXD+
mJCOUpfB0jcPEMk9eE+5AzDQqJTEbZAqNRDU3NMq//JxFPTG2C4MuQ+Gsvwufc1d
DV7gxB+SPer4+r73Di5TF367WhgZuQmbih9CaTHuHuJE75jMUYii6cChT6U/isAA
4QNkXEWp0midNgEKRHBOU7SVJD2PVb98OG0ZqHedcBPxReCm8uCTSxZtW5uLrAFo
RHVI5/wYiEH2vSrh6uZ/g1BSSptvQZU8EA8k0+gr8uJzaUFJQJT6o48Xk2pdHRkG
tVHnFv+PxmxIS6B+hbZS4Df4VpCXQnULYGxll/q0T0TfOTMhVyBoRfDt8dDzO726
XzpQPWxayO27+14W5jbNjQtu6zFcoM7Za7isAZo9Khfr068yWNTpnZRaEzGtgpIU
IG5lwCCP1dflWZse4t/kMGKczj5wz918cTCgzvMN6d6MLntMfJbTGq/MS10Rf71t
ul/dsdUJnGJoAd2M6RWVsUIpYSlftQYZYkXypuqAHNXnPK8M68sleiYnafWYs4Vs
MMoA7V4FIiSXy0eXVyRdxYtA15USYs3AWRaMqwLssMBsNWr8EJLlpz2GgFiQJh1f
pbIwQ/1TTJFur1q6tF0dnpfbnVa7Hk2r+/bCza5wvwNISlpHhsEm7VGzixKsiavS
Nc6fv1KFtTPULjK0CMGug4Rwvu56+bgSSNOQb12XuHKA1QxcWffvH+hEPHM4d1IN
Y2DltF0jW9kD5rZIwPEEeoJOT0H504s8+xQaG7E8k/S2xaWc93joDV1DfWK5rmLV
1gZaI0x/kN/1RWz3+cb+O34zIeyvtSo6eOvRFT3ZZDsT+B4csgy/YKgTzSPLfMoL
E7VnD+Ft0rjyzArlknKsgUVmS56/EEO1TfuxomJXrHllUYuQHfV/jFU1b3gYzbB1
yLgqvsLmoxNuSqxXYhVHGpMwTgwjs/RtEXd3BsDHtlD68YurtGd87sT1ah7mTyWH
TvclvaFZxAz+t4I7dgMLHq72dUdvZv9ABDh0GrT/YG8YJ1w8WiphlyJ1D/Rv3CzV
zfylEqLkk3jRlObMqmn9OihVQ23IR0f02np12SPYHAy1dB/bQBnWP+IuZZpVD6NV
G6LiCn/TOiE2dquOlITi3wVJk4i/USWM3zqkoLhVme4wcoRbDYfUInPs+6+sGQ9p
+r9vO7zis6VJLls97mflJYMIFulATjlLwBu9QIAbATcfYHhW8/R9LR7vH0m7+Plm
glYp2+01hAWx3gFLdP4UHhwiOmIYLh77h6Nibh7XsVc3S1UJ/Ph8BbA9ao+YM7v4
PzWw+FHCSz8EbOW00u8Rp2DGYOVvqSfWs6SiRAdLdFr3IqESpfPjNuYviKAWN3xx
/AmhvesbLg5ldik8JN6LrIs8QLutEzia6gRtzSdkD340BBS04h5qkVT2oD8mncam
hCV1uzJ/ixXW9TW4pBT6wWYTWcb/qyM30n+Cjxqz9EML9oAJfECrXgmwsrF3e/7D
BVsYG8EYTuAtmcNYheoVsUY9i3BbKkifrP37Imyx43bWxb/ls+DOrskuItKKaJyu
6fenVyZDwg2T/C+guxxQ0OfTremfDw3EHv27k9wp5HW4m8OEgb9exlqRF95beuTZ
NCyCnGB8KjbQQW1mMRk+qixtocXuXrVmIsj0BAdp9z/31bm1SFDHVy+W9uRqrOr6
3uvbfiRu/ErRJgmo3zM1/GROimX8llDza9sfKK8jAJSWR8SUxSdemdDgTockRWJM
FWIl/q7a9pbDgCV3QaxaabEKIGuEQl0p/r6gIJAM8l+HGHeJBVbc3so3rm+v/3Vn
4mqLrxPbtjkMeinIlWjgfe04GCRznOEh+CM5DjSNDrN/9DAbDd24D8Hr8dBMv1mv
1M5AX2HbeYfRWzry1lT5LQQf2fPHHa+AhDcF5ef5tlkFNDw4/UoKOKDWY/f+QpfG
zPAn+wxLJSoiu8eyeEVu3+h8A7fvZ6h0kzkxyjg0QsA6hE/ZQD7ivEEeNV/v19ci
1vb3Y8RSc4lI5MY/dG8NkQLbBPjaHyRLlAEb8wOYaoIkMSJBtCf0sRaqsLAFB/nZ
WHRgHfB7rsie7q/0srbS9T3aZQFZxaBDt0xoIQs0wI8W2q2W6UTWhuGa/GCUQKKa
ru/bIGerr3Qis3LSR9ruaAD6SHX/2CezTF3XJhvwbGBzdh+/Kq6NXhrZAz9PKgQh
jZ92kq3aMdK/nqGRZ/2ThNOwiGGzOJQEuQ7OX8JeyOw4SzBi6p/4VM0ynjZ4hW5y
/XZ5H5x/8xM8oLSqxsPGbOMuHHmaPnqIz4o1dR1+bkLJSsXwcUZyTskoeSOwSYEQ
q5II3Mf95+tWPqTDIuesafBsvTQX3WIqTAm/+iksoKXOKGrgtqWcmIybf6UwcH1c
bITBt3NV71pQ/rFg2EXrvXeUiPgrNvRo0l+vjtJi3hrZ/7FpFX2CtQYOZaEwfcFu
2afgm3gYYDZtlusEL4yQWxbnoSnCEzr7hrkrtYJJq4IJk9OIFsH+2fl27ILkdkQQ
DczZuxCK4lNtvyMLkZ6PjrPLaOsX1HNsPTWxnUGJcSaEK6e7e6rSHmdaHSA66hF9
/BOsUjYFVWGEQ2gK/pdaQay/r/7X6ex08/XrvvlyD92THchH5L5zAzYqM5IvV/p/
6O40cFNaTlg3rksAjSqVMc0+0dCXn2rX9xaK+GL204tOL1syifYcxfXkz/TCEalM
qO/EGs1Gu9BTO0H5nKTbDeqntqhrxL6bQpFiE9IXgchsLxO9u+FVhuvfXaM0qlCY
O6cy7VWDMkpmWQGtYOr5OVvI21sCG9fyCKhJdkBOqq47qZb+OYSYVzZKm766bAai
eCOLhA61Pjh+8FD84nQnSl2Zey8J5TQ/KsK6i4YisskrQQAxgMOKDGDeO3N4h+5L
ZJSYnsYaWAj74YMNQt3gyqQERRAwd3twqjCCRALWmWvypE4/z03A5B2/Xe9gmT4a
YJMC7gFsnHKpRKYV+pUq+WKxbsVZkhAEY+wegO4ao++fJuNq7PuFCEx1pef+Sewe
unrl00Yqc5nHm/wDGKc70wlm+dB8fcY6YcZUwwLSv6MvYRphgwpQK9otE7RPT+nI
rgfJ6+FicTJp6d+5Va/jZXNhQPMyCt0zJHfYnVVDxfjgp7CZ1UBzmNK9BfXrErlv
VIR57cWDVgk45VGhHkEjr4H7Ig+SWANv8GKMaAsAmd4ujzo+0GbDBTAjdgCVjLsu
nYn+InFJLLot2IBWVkOGS54EKraNpqW2kyczrQLOfgEfwcJPxx/hP6vPacvV9d+o
+C/gcWSIAXDmJ2y3CVGegS7bWTnJ7yxJhzi3nEkgFEzAvtn5R8LnwnSYT/p5qh4v
EjfDl2HZdXAx2ZOapaf3w2QtpHN/qN557ZJAyGnkCTEJvju7qMXhnP6iAF978FEc
ef2QrRSvZUWKQkoK3JZaNM2ACIcNjR3k8BXWKi0FK1onS6C2E5gB6mrnTMc1qPKi
Eh8qNM8CD147tceE0PKlivdhbSk7bAWKdeP6fiK4iGlw7ob4XaXFnN43I0XdrJ1E
0XSufqYMlY+igE89dGCd+wZO0uoovh6tMbN/KHiRNNjR5M+KhM+qpK04DqmPKnDj
rlYdCJBosoNfZXwwzjPr8l38CcQ+FVeMouqXp5ED8tVbLC5Q7hpJ7g4Y3YvT7/1h
cTwVhaUVHtLKwKQ4tZvybOaMput82youw2F4hA/sTnF3aF7vFGCtT7Jo6SnQvkyM
m/2TxZhS2cwfabaCsBQo2jNrqcfPlbgXvL1bPy9Z47WkASA7GD6wFm6GsqsIepfO
wfh6f+LLWn0QNt3WmuFfuYUOAsOqPBLhbe/PmXrI0pe0kIMfz0d9cCrN5dhZUJHy
VJxAxwLBASsqMDa/jFDhMHmlEKgG5UXw5L4OAh8/JkTIeTKt7jtD9aIgMGu8GwGP
CoA4+PMly0doss6+YqX2D4eDDERRQvTScobrtZEs2Xo62DdqSrLbjXM5sYQEjCN4
i841LqWmCy08tP26Nj5fJdkNGykJoo5AiXZ5QpTZiUDJmEnVqD9xP+hAV/YoR/cO
fIRgj4XRPMWNGIOYXrts52F1+Vb5TqOE31E9xPB9xRKSm9b/HD6CVF6LsMMF2eUE
CIxY/BNNKJ06db9IQSMDbxa8SVPiQFLTh+/ZzPl+uPDUcT8KZ31ClcZm6TZTtCBB
+8Wy7t0WwZeOl0cFIBaQ4q4wPYlLEO7O2her091nmiG5mw8ebxLfxy9tmQApBQqM
XSzqDbsK63sgPHh35kkdYE8nJBfTNE4Hj5J2tKNV8Mg+pdXRMpz+H1NOlNRy1+le
pjnVcbfbutv8XPDPfe5CPswkth1tUJCPmfW5tlWEd5TJrJ4eHLfdDPcfN8gSYMwe
yQ2vq3MrGrzC0vq6wPlY4LrKPCODNl8TvwemChB/ajnwYhnyCz8x2Kmhe14TTKe5
jE00IN+iWhSFGP8DcgaMRpgJxaTOgUoReuA4qmpPtHNFImkiP4DBUYeYaX3ji8un
cyl+9NDZd2jCIlRxXAM8KJ7ic/Rg4GLGQ7dVdJKDsmxDLtZPdpJ0lOX8efZsAatN
ujmpC+W/X8dJzRmSo+dKx2TfE6/OB4nNEjkBuLh5CjmwZ2JNQzQbpjn7IDCifBpk
/jvr+wuOtLzsQHEMbS59r891sqYRsH+L6HGsXA7nOQmkByehTlHo6dUA2jza3j8N
UWnsIo2FdevYdS6J0axOfeTpak2psfidf+TMXZ+9vRdCq4IzA387fy5aTqkHQRI+
O6HHXlvTpbPgXCNHF7nDUJ1edZfubxx290kt2uBljKxM5C9FvrY0JVvRo+CLSxNC
nuePsGbz4pUzaZGDQc+kgrhYuUyBmZ+vb1ocpei7GpEe4I3+H1m2DtrJYYHOBvG8
pkzCAswtxnArO9VmJOK0bghY9o1y78wq9nsFVnlSwZpENzV58SZdrFkQ6UsbUO2U
F4IWu3BboOLcGl0s+xzQtqHXb3iapMm7TFSCqph2nytePeliagOAfCNYe8zKYRbg
oMfcQpin4fzNlI2G4waLxT9RSf9/YW/zGjL3mlpzRDhd5ZCtQpG5xgSLls9m6/Rx
XsY+aZPh8a8Txdjr9o8eCgvFUHD9hYfMLnXZheodQ5jL/HjWpLyDyCjGHeIB7Ewm
HQSfdeihc+YHlofhUF0aYODtj6SWp3VztE7qpsUdCPdewC3zSSzpk9UcYdVuraTi
CMvzPV4uXby5kcE82cYR1IssTYziJ9uKu5KyTzqg1Kc6Zhk1MWm0jRHwagU0+fyP
zRaRmgvIHUwk2J2LzlousXaEamNW3lPwsY2jhluwjsXh9FvpGbSk1TvlHL4R0pww
nFAYTxVMkbfqrDNtnudXWIK9qA/g/tt+V7VxQmI+a+jINIRtLV4n/hBmmJ++dSVd
iNuWdRexEk4BxDdol9ChjkygfDvFuXqOHiGhjnQamw1KuH9gOsrAAclAgK+Qqm/5
b/8F9H5Oe9NzB0BQSQ3F5/og5TFzqyu6ZBNV78KuNQJ8WAD0UB3Zz1/F41Tgzs2t
zY1rXxtjbA+fNQrC8Q7hNbzRsavuct8sa2bbjEGAaSmfsY+7h7gXilgpDdN6B55O
XClmiG0dlzTmXplCS5Nn/TfSazJqnMyfR/tArz6iO+GMuuaJ0qOai1PEDVraVizn
uq3jbnGjCjhB+aewFSTipT7hWP4QE+NYB1DlAsWgH6A4fHOH5KZ2ec9LdQfe1Irs
GGIsN6er7wQDIdoom9j5nKbC7ymfflezD88DyYnG1AfP9JklbX0UXnq9hatif8q3
KiqChqqHwd7rHIXaguONs+PrjYm2ePKhRzcGsV6PGtRd8rO5IcE0+yCqkNKDb0r0
uWZGqe4lkXqcWc2G/9aLa37wn092YCmIyhfW/WQ4/gOlNQvHhsOYFUz6t35DBSMF
urLtzfXfiuZq9i/7lkTBBNnHSvOGlPqMlnlA8ckzmFmnvujN7HT6O+BE1nzTXLID
he8Q1bpnyBpEhwSK6M1N6Qy9qImU/vQ5/5Zb7SCLQaG8uNVjLJKWWjdxJYBWfP6O
q4HF28l1H1lsBXtK1zzTEjORgn2J74wviQPDSqmFve5LeKqPr7FmKPEE9ajSC57z
6oe6+r5R/W/Y+TMneCAHQZeQ3d1dOiuN9+X23y4xOcZWpdnMxIedAjxe5SywL/ZL
3IoiYqmhLGSXFjC0STdyIRnqfCJcnNz7jG8HrNCZWdmf7w7YPL3GkdIeR1VZigM4
1KnTgT/s0e49Euw6ckvZOeEZrIjggWPFOCTYiFuLtpAIpXhCZyphBgCJ8H0eJrw8
gQisBK2nxuXTdvJtbsCcgqBAMUzfqsrWmVs8WuvNjs47O3PZRLv/YMTT7Yqo5X9g
mef0D92EyHpdJAwiYgnR870DWWuX7bg2BpfNwNI3lhW5h41WKLsxA4ljbJ3QPS1t
S4NwfA1wScPTwmSh99vR0AYaSy3VhA9sDZ2GZ3UT6i9n/+E4qdPfNaunuMjpcUN9
yaS+vU+/Jvqen2LzO9U06qC4cck0DL9vGQ9mGuWllW76RWc4+TUDF2VqeEnktuQD
V3WDszV6KejGTHoBA+5LFR5FUPMDRUqG+aU72ATD+OOrk+alX+PHv2L5Uw6543GA
0I4XPqZfBOQ3R6rjAVhB+iH6oNVWrTBhTBZ3cl5ikozwn4i6nz/SRnMdqYp5cZlD
lpx+rdqlOwEdMZbDIBgUCVtexBssNX6KlBB1KYgl4zM/fM7w4Odg1pWk5OR5k1DZ
+tHPE6X2BwnTYjlwc6EqS9QNyEf1wOTLKfdjNzi8nabo4iXNPKAhO2NG4zY0wyfS
ATscXP/9KM2OTYfyhdJpLtLv08D80Nc1cGNPsbvqeMcluBqKJgfnElf1FD1/xqZ2
qOcW8an/tZzBPIIL3SW7jyqJk4Jj3SL4oITWYzSuXaNCS610FUlhn1GBIbNjDxJg
y1tgnWx/7PiRQcIlprNnCWaiwGM1q3umknC5brK2SujVvPO0cz6lQussPYWC8TQW
F9EwKg4xUCTtVD2HWVXhvU7ZvBX7ByGubO6v355/zCFsHYD2jWMMfs5Mqkpiodc8
NnDgamD9/4PYL2MfCKu2Nr0v6okqXMOE9oJ6rQvCEKG1O1HiTUx4RWDcOgmBiGY5
LTJ6DIH0L0xA/fv/SGJzlVqv6FCQQ/f/vzFvohCfLCpgIVVUdon6v8EenlhR2s1v
LrfFF2Wdvf7KbzV/o7YPmOtpb/Jgc+V/5DvJI/UkbJH3fds9sMezr7bntwKj80iF
B9yYaPjBVsnBjhq/4fBArcsZmOvdjrAAheSFjg4r6L1XexWdBuLXzRLkLpcKMgAX
i3hmZiNHeyKjqFGZEBXaeq23vOfG4CFZ6iCz+pb92wYYcacT3vCOHkONbDJ8Ktq0
0ArcA00dV2QuSIWrZPF5EMS9oTh5/GLlJjKTZ55pYq9rJgnGrV0hPPNnJtBv+JKf
9orjTg5A8n6dFuGWz8wVqak/Zuqr4sH8q8cwyjZ7geFyezydU35Ts4hWddOPKHGb
9nd4DU78dEl1hWN1C/4xOx/dIntKMjAhsfWOGmr8fBNoMNKHNGfadDBWkuh3WKKC
E78lmxkPqPVt2UpidkLckC++LhNczov3StLoUf6tLs7JuIxerxfzHdlkIuEfhIV9
pIiUDFYLV25KTN8zj6JU2yH4QyWdWg+bNr09IlmQoEnQH+X4GJkzwv7ypvtzPWSW
VenPxq13smhDLmDlfGOSW86ZMZsHr2qa7gkYRq1U/cQ6scvwZ3UEl88Jm6CHmkbs
0J5YwEM9MaE5TFq8+MNU92oBJPdWN+iTjnaCJeLcl9/2PVpkfCwa5yUZewvtKTGw
m89D0sLL88IJ4Z8c3pY2U4CDg3kdYhEF6gJjhwAJEbkkOGvmNTEsVljPGnxEmmMw
zpoTaNHhTKRN7RePFN76iWhBXfzgNkA+WEcn4ckhs0gl9Z8bYxFIK+xiqiT5n3rn
CzE+QjmnOjiQBpkhoVrhoKtrkAv2MKu3vmMCQtrJiiANb5hxDyYFVmBC0e9l6YXL
hNcIAaS9rN64q9CuQ4PxrkeKA5iAUC7UL6qkgMpUNRXIGfsAwOF0cQlnWhTlEQO2
B3PqUpLY3Qi17Dh5JnDO9c4/hZXcmMcZ0JMR5BawI8FXz/4uXlwcndCvFT+YavVx
ybaWWlhlIBB7crHOQ3Og3weytdeqwtCzr14W2a7y3C8drHbwRMY4yYFCTtTIktss
lSnnoPKzMIBE9DPpk5QGtbUN24Tj/ZAnWTDuCLXtDjQQSnewXCb/i21rJbDSQ/Ps
iG1ND5tEWg56CbZuExrKtBAUt6sgUazGFZ7pUS0k9CpbswdpoRwTQ4d7SYi1rWsb
UR2VfXp5cE13vGJbZKv2gk36H5jzgmphAQOW41gQZSsSAQ9GA5xttFVURa43dgjY
qgtpeSYbCP/skiOd4h3AOqXvYgbzsvdbE/VbCWfxVhp0xAZKVl/4pGwQze8uEKCU
fRZuGKMn3yvHbPORGEiDMFYIHChOFfuRICIVybY2u9B43Hqm1O90H6IsBnelUaox
3Hr49WQuKrwppM9l8bcBZENr5GfJM/46fu4aSpyZ+8Q6OzDL/YWmwe/j1BKQoqIQ
6Gkwogp84FjJ8ruEyjX9r/5oAmxKrqzbSEsZb9BvUMLetB0PaA+ekqOBKsy8kD2o
KveMbT+bzQZGKoJshxv4GQc3UelZoNj07nYZ+lzsUK7DwiD/r+h2FbMQaqkbF7x+
AIDLDfLDDRTItf2OYHkpTrwawkhOL2LROMtxabvenEt32Ijavxy415nlxa7+NA75
B/7vpG1OPc21tWTV3OOvK9Z7pJLwglK/QrZBdkDFbrvF/2AHdlb4y+tClbx4NnSA
CAb1I432CnOeguna2gFFdfgvjdfo5vEPXEC3hORz9DHnvf8M8utwMtlykMb0Ru9w
fj39HW8zZ9SzL54ATtOJful/zkic45lfamXT/SxBVxK7m2Vf7bhBPZehHBib23f9
6GsBM+uISBh4GkYzl2wZBVcPA0/70dahoXAK1jR6DjzggdIR1c+YpTfi8GBopJ95
/k48Y8bL3yUzJiNvCZFrxYcv6b/KV8FDe79yfvWzJqpNtVaf2EW3W07+mZbzvqDr
1q9gHCKTTswrZa3PymNUFe84QGE7tRxSq2emaHui4fWBk89I5rcB9GoSFJnUdVlN
xEroBl6BI+WCZpGOxLDzprR6VRxrCML2Z6JbsI/HIcReE4gzPqV7nN49I9/4wQQ5
vTqmbFk/0C1qmkJSOU18pTScJaVyMe7ZiVfv5itxY8dlu0r5r+6KXrl2ccFMJaUh
jLukvgDwHJ3mazwLIQRKuj9PlTZAmxQO5r/dZlvkVb6PUv4VUoGoHrxwtDc0jemL
23QLttOY7epjgRTNeyVrrK8Qr9Ft1bZt+S9Q3Ys6KOG3c3tvJmUyOBDHux8OBHJ6
9icafilcVcFe65fDBQIe6HgWM4LqFuL5QNGRIuWGYyZnbQFL3Z2Znoi5E4XniMjm
NYsqy3MlCDMm7NhO1YZG3HZiIyQZsMpmRjmYsKzdfQ8Czokz4asWj6z/99GH4P7d
DLu+Zx/SaAQlGDuHUSF4WhyDvh8CCeiuiSIcqkVuHXsdGWJbwaR9MX2Tchka5JBR
Pn1/3kVvXQaqAaCCx91fcbu14U9EqGgEaY2cS5ykipAzfiRhX1Op9XfSgUCBgpNT
8nPMle4sjn76QsNV3qSzTUz+UeSkNtXXxpcrZyPBxcnWn73Ot/sFfz4F85AsWTy3
rVSPHF1Dm7Go/1E4zpBTVts8l3v0Dvlxbscpj8RarC88eaePXBOwkBF9Mql3hIb/
MPAIZwDfs68g38bNhQ5Lw294grfPs0XV3oJZiLAWCgcmUxZNVZb/KAT7kt4DtnY9
QWx7djFAPZdYmMX0tXFqNC++SYjIyp1kTTulQF5R2Q+Kslh53EFi2Lsf3wGK+x20
kJhatCoy0J7RzQE+0z5EY1UeBpQxNMzwVmSQnWXZ5o4fGCeKikqrzQrnMXstLTyX
u1HUCVy/YlRghJ8efHu2W5qX5+oaoVHCgwOYJPCyekfx+5fm9tO7O4zDNRVFoJEh
OgtlplKGf6pClTos+9GhJh7W4tCi5YbxL7vnMEFK+zkbiN6k33aKCXQir4b5CeTu
Jlsot8gqTHKJm/kx7wt04BakMuVjcfFvu8io1jEwYrYK1hPPgeL/VuYZ7HALbmEn
+QDbDtZTC8awxQahJ0My07cyLI/02mIQYlndqRHUihphl8+chNU2+7AiGEvtKjp8
pZHXMlscug8cZYMKbY6yYpasT3jInIC8BEWBHbNw4ojo6cYIWqiOIxMHkXVc18IV
UoqmeAYBcTmi+47IP1CjvKYl7MOhfmOFCKmiahijHoYuD77YWTk9XP6zTat2Vywu
Kv0zxLN8elMcm4TritcqW3TpmNje4IWmuF9yRHhkED12FGAa0U9PVboiXrkp1LHN
oaiSeRalLZoIdpjmSoptV0ucc7xCBg2cjars8XUugYJ5tWmjeAg0j5PnWnpRUf7W
kCGPguBQuKsQOgUGbRFCYbFb2DzchsSHoGm6euGVEH8snqlslVnqPKcR04nAe7Hg
dGLSjnTmYLo49OluWJbaljssFTEE8IM26jQaXSrqKZ0spxWt2XdS5RHoGYA82IXJ
HXiHT0uomSkKkTm7lbe7XkmwOMMP5cHun/yAZ2kaJjUxCQe7RE9zWZ1b63hvBiMu
kAc84aUDUFt9jWVdkULhT6Ldq5I3+Xa6BlRx5+4Ls3h4YhgU1Omchym/gIu6u80B
1NxVb+vDYqBaoUNVHSU03sNue6q2ILGKVBz7/7KIQId9O80W4IRtMP1iEAPWF51X
lFEwu2jLBiQ/AcjZcgvxYWl00QtLo2RBepxkoU8cbE+hT+IwSZoBEh29djl+k8yE
5BVogMFv4jLLsd0u3bbEX41crLm/KFKfYjEGIBUS5opnCdK857c0GVoioNzwBv5x
QEk9aFNtZl8M8R32D4mrj+pEK4HZYkpTb3jaKXlAAgKVef9mTBIRjKKN8poKq4cL
g3rzjNXoRaZOzdat25+sdCXQVt6Jqiy6/FKfdKrw3KaN5iT+3FcoT7yhXgtr1uVX
7tiAdlxykcvptTWuZKm9FAhrEctvkEQgkdHB5WWcUs467bP2i2oqTaNfr4OxjHQs
AmgrUkTwgYztNQ1OAPBBPm0qFYWul7Kp4ezJ3QYcJhfB1IULdt49hiy8wjN+LetD
NQ6wOMjpaIKHQqvk6UXFzts9i0gy57Mr0H88YHulFopvMeOeyp78E71PGx3ELaSs
WyXXg8kGB3WRvoYH8cPasaF6Yv9p3Jb7/I0COy5W5UHgJMLlfh74dlHPgYO8XDAo
BmwGVa9s6IseQB94swCAh8mgOZrp3N3oovNEu/QOpy12z8SbuqEmhxHWtcj/o2zF
kqdzaCjvnkaut+4/onzSTV3bC+udovkVxRXjkNbw4vAUQ6G39Ot9zFYs8zt7EWnT
tlRI++xY3KrjGxoWRMQ0cjYDWQ8E7jcrs5y/ygakeTmFue2wvxft+d70RCMG01n0
3CK13Xs4vTaxFNml10pS7vJPTIsLJNbRdLnVMFtS3lHoWZuUcKcQWIW1Fd7Zy+Q7
DaV6oU9sZZZxAfoD7osmOJ4oJsdZyH3Ala9IK8aGHrKXgf0PNsPA1RGvVHBsCh4C
CWOPaq6SqvefNZxuD6AqGlnroicsofYLXzBbUc5qsJrcG7dP0ghHhmCzC65GmoZ+
5x6C3XYD6nVPt+rxEElwSlMClMvyyvMMPLTSki+v/WNUyvuE5sy4lRAVEznUvQPx
JNRkphv5uMB+BzQNniBdE9ywHBR6GMQ4Agg/nDwz2hMDKtSxVf/s7+jXGJBA/L8Y
IbaQB20LReEaoWY2/4NBY06i9JpG2PYsI0WUnDS94YkU4bmFfpUEFYaFfdDm9fuD
3idxy2hx6tcR42uTheCA8Qlz7KCiubdHw863N1pOYRdWDuQPlCGjHN5WIaD7ePx8
8dFXFgNZHFznW4PolMOqt2BHxsMZBvjZNLpVs1D19pyjWNCctRLp3+GwQQhGHrJZ
i24WBHlUgoU++K9OSeAzWNraQ55G5eonUOEmq1zKVHBLEgH6KpkPCgUhkhzss/2k
83nx62jcPfSadExV0cFy18lroTT1jrbYWiZHYU4jIfpU8HMdDy+cbmWQdVtzmeKw
U9EhN41gPlDKSf/zUZILAGsdOPFN4xND24rxvMOS3i4O4wKPn4KUUMCakzBSXX7b
hmpWVv68RNrWItA0cV/+NioVZuqZcSG3p8zrfrW1CGQyK0mosjG7PzLOUN8t6qbB
XmneLT92wkkflZAkqqiK9qufZI15bNdykzMQhjH244L8mMkA5TuRzgu7RrBPJSPc
N03RlCI/sOLI7iHsAmibzizUdqLQSFWMduy9NNXlCq9Of39MiV0baUgkMOr7axXu
h33gCwTLbuAqBx0QaexWxazrd31r5yJUOFjSjhuamFPMq8UwCCGexUUXLsszBbeN
fmUzfDASTEZ57b4rSqDqvXv3V2oQjBd/cEGIm1Aa5RSpsoTRLrM97a6isl9aN1vQ
SL3Ni5EfIFC61loG+dDk/pdPGOAMUJrlFSHXWZdOg05OBm9g5Ol7IL+VmxizAyQM
yLxjqxEsNfLj9xyNxbqIK0/4BOHdcRWnk7fIj1mr7ZSFq+3kavsMbrt068AaARn6
2X9NCociCXunxoJid3/T7X2Vc3mfGmP7IwQLcMO+eV2sVkzq1Eo3f1xTUv9MqArX
N1J78DnmKDrzTIEa80oJLtaEDkCqZzupSSrrEVsLCa+OWxn4LNPfS40lnWcPOFTG
hRAk7zu/qwzblJ0KJagQnWb6l6kjkKobYXcbBbcNaR2G2Z4eXi4G2WIEPvEx9Ex2
pYt3D70AmFeua2DFXgP8X+GaqOB5SpedRKvz4+oT+v5judE/2sqBXnDgCx43Bv/L
3szdfSgPbUfrqq+Jv6j3eqsPZUSvF6zCbdQpvQglOaMvhp6YsYOAad9tPxZSxEJt
OnxK6f+4nfFwev2IBWZ0fnGpdyJVjGu/kTDTzy8eh1DJBE6dPEYtMKYd+de9h8Lk
Xcw68u9O/jzLIK0FdpfeN+NUWl2kjQxHGYGmDBDw9juEksZeFSwG9MDAAWI/YySB
aAj+LBnMZHlsWXX8JhZIIPUPYa6bOFflx7Ojmx75btq5BVZaMBA7NQPpCiwgqw57
qFG0eKT5nwPdRHp9d4lQLvLLaBI3OQtHKPjGJaVqp37TPeNF9plHyGbFv8uNJBaF
Yp6kvZJYhFI8S90053VhLaF7sYtBF2VAByE/EyiErHFIvVnCJacwY1YCpr/8gNYq
mIrW4T4hzjrVxm1QqS09Kzxkdy58cfm6HkLZaZ0kwuvenphOZbLRsBFWrYNuItRJ
90465LhzfRxGAKPLquvNz4afiOSlPWbpPZdhuk71hfNZUHAmJkcRwHMC4VK1obHL
W+mjQDUpXSpCU/BnZTlGwLratDDJeWz9VQYgB4icsaSpIxTw6+Z2jwORl04rikMr
uSzUMe0m6bavd5NoDOoHL2I+Nw4UI3DZKAx7Yvgnvzsqio/lmO3jfdlPBmdbM718
oAPKny7QNLzm5hxpdDtDlch+pWHko+GJjKW3p4ZMDjoaY+ViugZ4shxcJaRfO118
8TvPUMYdNugL9rRrekRJyvDvv+BqP5F/75dLdeZkktxPnmIDNNfZVVu4FWxmXAel
N5zkj8TSpIlxO9ghpnV2CZLCb87CCgYVyXiSevlG1cbrDQdDyJoSaEdlVLnsBwv4
KeoZwtQHQB9W/ABO8TnYKWK25EPhp5SR2t+J9lB0RhA31OoYOcfxVv+JTJJmLtgh
KWImk7SkA/KOmlvquNstZPAj70aCDkt9CqzaJnnWnTcQVEXHsTNPkmXqUZe2pV70
RzSrOjBTzRm4aA1G3wHbYVv14ZRCVoANeuToxQgcAGZTKb0yYikjAw7V0/qVzchX
v7PnBmYSsnTdPFx0tC4qvki0Vy8SH+TLxi2R7arlP4SlDT7T4/5u6LM9jZgYev3M
DGvsEp0/eJAgboAAAyzjhJCDj5WV9LMRIyaz8OTIBUniC+xazj2HhvBmUROtABsx
NHgxr1uKP0Q6L/tI2ZdOCc0OxaycHuQ9Lyp5EwEzeEYrZc8/CC0TRspJvxWA4cXI
bH6ArBeWZdxwoxNlSDlMZCh+umJH2gcjoITFsmW6oMXRtNghlKlKSiW2H4AUyvmb
Xo8liqy72q8Wva9RBa1mowHuY05WTq2PWYgNKH5Plhy0WlV1GQPjLK5bcvM9t5Xd
hFKisf4ABbMIxv/Uh1F/fP3uImEP6AlTilZ3V7OhExRLdPAlprR0W0ghjZBq6auo
T2WVlwYMFdPRSB/lbb3Ge3lTU2mbi6HTZ4agl8vdcJ8cZSXqqZnhZVitBaGl+orT
vGjuCfoVyL74gmwNv3LOAQ2fKJfNrzNh2DjYzFed7jSNNgTVCzz0AuVEKUs7Hm2j
44PEf3dLn+gWo1nGrBmAD9+H81WVHk3+1fsS8aXsCx6lKD/fRQYq0qjVXZH1F83N
rYgvOF+5v7KqKebbpXLESh0M+T8U1lF+G98SOI06piIdv+5+uAEQpO9V50uw+KaU
pXVcSwCLDS5mTd0QHxy6PQLXVfiPM1J9Wo/2rzQT7Zwcer481618nW17cEMuj6F9
cqSe4EWYxTby5qeOULDaRCSApyqylTBoUVwxScca0hYmeBzzJnpoimWCIeV1pHK7
ibRU2pNV07vHnKwL7W6tANVmLuAdxvqkCWf5EaigkSJRV0tDZH0j+UK9WDvuou6L
1h3dtVBJcTxpgiCpx1af0SlkuIO2hkuF0Je/zCNq0+BLp4wawaV6Inw9aukFxLkr
Kd5KhOpF0R0QXmI1XOtK1Vu6qQGeJTNL0wFhPmGOXlUbYbcoa1L0ycAGjeaQ/K1y
INcwoWohBruyKsrNyROJnLLMC8544hrA0JM0oFmXwUW2fs0AHNHOXL9h8RycGleM
ALqJaxe877/xUZoD2wh63EaOvYYJ5JSvLkFwveXa6d/kmcUsuMQGbqtqAXn7MVrn
j5StsdATsROkvsD2MrCzJLqDfKcSJT7JQgQqEVuuTX0BOFtobYkN8MRZzQ8YXRFU
SxanZzUX35pvPmhqvvVHPDBAuxIbONDyRXWeIxSxrV9370KySu3Dtfztddl8YB9J
VVM+KbfbaHzerl67lFOPBk21svZk8qFLIj8s408SLCadekjzblk0BuRsKBXx+ctH
Euy+cqJQ68NHelEMYaiMlJZFB4yg2Cua61QGqBjVvojBbRZx8agzs3LozDgPW0rT
SlmuvGaJET/LOmksytl5/I6/UIUX4BaoEbxf57aogxMWWeGdzhk+fyhS2OUM0GX4
o9Ya3ik7Vg85rorWNuG7Gzb4Zn2R2tRUgYbihNL8rY2Ej49dlxFAhkma3wpoVTHl
4yfWYy1NUhLOp4FRkmf7E1179/6TuPl3am7yHDIf6T8CZR/8q1NboM4j5ryNGq10
eWEE0gzehx2iuYitKIT3kF0BL0bVMy841xAH1f+5UbRfrFER6J0EVD5F3pMYoB19
+CqoMP2hBvJ3UQIqtGevImdaHkkbjLVP2+oxsMbNg2V5S+ipW+Ohqlc4pTiKftvH
Yav+F6BEjDV2SEBTQmYbMoMgE+8RjCbqh1xa/LfP1uPPeb3bRICA3/LEOsD6ZhB9
MmhQnWeLAWE6wSs/eYKu8+2QgE7iHurlnnuWCczmMAEsFWUyYdmnXstYu784HGPo
tgluylrEFM49IQEepIgaas68ci4zUFYt1++IN7dbJ1EGVNDF3YIIuUDp+1jDRfm2
GHCxG/ZWSEgyB0pbjlllsT9tcyBSSuXW5umNZCa1n2Qq4Q6mCH3E5hKgoF3qhF9h
ubURDczD7zclP0/9XJBS6PNI2DSNyR/omTa0aeGP3dW+g/klF09G5WfdsM54l9sW
0ZriNc2NlR7Klgs33jqfVM/BFAlIXu7raRdiwwndWem1d+W9+ObCtesPdsHey9yf
/KgBYvQGoDXlZVtWov2PeHWny4mqnHEsr7P1Zea1BcAYwflw16Bsod6M8N7zwdiw
i0jQKWVfgStCbCEl2qIEFSGvgameFA/jzIwj3w54t4/f2AkVj8fDTSjXkvc7v+ix
8/Qa14Iu1ls8N4+DD4rZ5O6f1dGDv4xiJNGs3vBy16W88WgCQrpDF13+KFCRfdJQ
Hxec+Ci24lTjIjWRwfhzMpgYs9fyO/nX38ITTuoXpMt4N7VuzxlgZejGcRboZBi8
LKbyU01omlrrxIULWYI5m28eJCWrfazRwt5+l8A6KPcbWU3SAKbWcVWiLpTTa5Nx
Cx+bVVqx4NSy+G98c5Rc9ZigIgKei7R7f73LFRv5d1yriA8QTb7jZo4+7GvFwVjW
DZeh4UCUzNq7cmvjOPk4tkXEx8DzWvTHJsTQHV/Ko8SwQgBfseSt/Zy9U3BoVvTE
10uNr8sNU0mwBXp7HmZHwsltRMd0KrcXTyM7ipmBqx4r107kHwGex/4ZN+QvlGrI
RhKcylLqp5dL81HV3hTlCZpD87MzeFPhoBf48qOwPmbmMzSJR2F3T/GzYnboKw7w
9s6tVw+nGByJjv3jt0yy2R6yhO6Mdhi4lVIjRqg0xto6mYywu7qX3gQhzovOh1Dp
sYjaJFM5l7/jO1blZUG12q2JNG4HY1/83JUInwt8uoYDQ52ylR1+NGd6142qn3ml
eRIDgLyKaB1MVy+UkC0W+QleUfNYCxqNidfWTxECLBEHy9xy5g1jCHUVnDTR0jut
O7ZQIzfE8IeEuukTO4BmYLogh8vVUzxyAJs8gQFBr2/lslSzvwpRd8P+fYp1Z4ks
VGVAXN7o68geSwEjo6Kf1qu94MDiTXhMkqy9yFvB2b3QKnRT03oskfpJo8D8KmzZ
76V+Rqjcdj0hLLX6rFn9K3H1DF/asJNs3fEBRXzrKp+S1LAnFLwBblikYT6CzR61
dNQO7hK21IJbqAjhhCqnTBmrrfUb0EG4qH/JwvRWTTqHmILEiOjzWcQ8oSvzILP0
4IS5+lFkWiP80ATJSp3j6F4Yr/FJner4pmMpEJJtkzYkINxyj4mjdP+IkAn+n84T
haLsULxsS9ttubC75wU2cXC92/4U58cbJEhUEfH/RAHbWoriARdcD0oooc92/uAG
ps+opR4lVrvXkeyQjbEIh1+qGnqHhEpk4+jLDrNQfqnUOrFh5axcLeYAaa5Sn//u
Uml/sFC+iv8gBH2kvN3QYwWgsuVxqoh20PMiyUmhlJuOafSKADnOkq9LBJ+lOIpd
5tlbQ6ujucZmFrDtxfG91Mqn8kwY3F0v2fDVdzNcKiiV/WG7kIV50UKalDAMMB3y
6FirEqey98tqTeDBRjDid1kqGJqWU7ounFrc5/zjtb7GXwXpucc/8OXWQxjunUBl
EdAfdZDnxo3XO4tk9Kp13YStd8ZeFtcBSpKaLuZkZh1m61bvitxKfGMtXVw6xifA
mIyIlCuUFgomTWDLtZqRvlgk84SNeujvwdOygQMtECNf+IsXJjsy8qOupmJ6OInW
wqYEfJTTiJqCxMUPSOrjznELY/z1EtMQc2KfdlAbYTnuB5azywXyTlNyTCmSGmbD
vSCvud2Qf+GV/eEpWpfXgFIswQcBwLOtLCmO7/mWOvwzGkaFMrOMF/VyYOH1HH7g
ohBsKT1xuBg2kxbpgn8fL1JOsT/O0G1JXm9RKmzVyIsBo5ft52anJl54xhycBYM2
beJAQU3JVT0lhyZZ9hTqrOFdNdGe846Jo31CiTb2drdMYcj6/e9UrcVbaO10Kjh/
aznNy3OL9daosqTrTudD3eVMa9jDVFC7XCalNlwqN+uWofS7XafOsKtvYLHL9vZz
58T+87TxcqtVv96ug95xPn+FvNcVHmWFfmIi/e9ptUe8DEU6xOz8q1vrw/ooBxN/
rGyE+Th05qgRbftVeAds+rDCODDNha5d2m7RCpEGXK178N3tn2IcZgC6XHJ5OXDi
3PCbVduzXVle0nXxNgL1t96U58oAp1QCyW4S94ailSeAQ8bW9AJ8USYazNx6TECa
fOIgkLU+1mctabQv0nw7rkS+fy40VM2M4649xIAHdaIHitaOYk0fO2G9Ee63cUeG
cQjxQYovugFPiAru+v+UMtMZMh34TkTIcDXW079ZEligrHFM7sE8RAEyQ4EXqHG9
tiX+zIbvcnejH389sUCFsSrc4d5skv/+/Wl9YGA1EqNvQrmxRkwCnQlxSKz2LjhA
skLVMfoILGAg1RIjKtNcAWnCqFQ5agxFbwYESsROVJkmA9k4n+yIbQqmyUkPL25V
19i18FgLoOLcXmvUtSYh6+ljSMO3JchaAEBsC6GQ/N05PWshr4D8TxkX4y1pJpYJ
s2fo8gKAIjLw7V56Lixrhp5ROOWf811RI/yWsIUnrVuo5Djd5FNlPh9UMOox7Jdh
L30JA3Qu36Z7zAJm7TYIau3rmalhaEgXmw+Va42UbSe4FB/O/CRb9X46a96tfCV5
59fcxt+m0qtHaem5CUAk0m6sHQPfYd3szS6bP0HdaMwuvCvdm3pnKBo0N/hCyIxG
z720aj0gHzjW2IBTigQG/2+zagofGUTjJpP9Ye5fqzRbem4bmEKnr8VJd2p8D0wd
3TBZxQ0925SbjvedLaF3Awtj27FpiCo0Xe14vDtkYHnA93oFhFx8+v+e9TfgvGW1
F5kqQ2MBn5HvmawuIexKvQk+Y5TyU4EmqBzfStmmwsDRSNcIOjtK0opiOY3qeinh
lpw66OPMqmmGh95DTJ/C1UeXrZnNO6zAIRsk2E1jANgb1ZGCKtQCtp2uqhImJ822
xp4FQ7qoP8Ay8qHi8f2YW/+N8l6DLx2s5MSjCgswCHcmMQHPXoB5PK6ySseZHSq/
wZgU+ShNKxB+4xtFSwPTwpvilZn/7jXJyZlLVwiA79PKLY/ogGhmVMuih1RNF4ik
F+7bCi61jFX+7GY6vL/SBLcuL3ewoW6ogQ2bKFKnMfdC3Kbkc3OymiP8vOVmb46x
+rEoNDqYqu9sB+mpoRsJ38u4kpH47b262PS8HfECEf04lMtmFYehZNSsPbLuCMiK
2RL2bdXbWNzIPVX8qzZ2TTfluB89YfceiMG8kzA5GKOLD0JeOr9d0wnE6/cOVqW1
bE5337np3Sh3ycjkYQOJnXX4U2nMTXjW8yVnHoZBG9D7f7XupKgAojSrI4WRTT3I
z6H3zMPYlFYUW4c336aYiCw6A+AO24O4GFyVquPLYd6flyIVbWui9j9RdT6UOCuO
uOvcTvjPq+LO4T373LD6FmbcuAhTm7KfTtT+p8DqCAfnJqC/bmLa2rj88GbCSRsw
t4yF2YbFS9woMSI97GZAgdq80PMdcXAVhztLNj9zRuPS8+AJzTsrFhnfFW7HWjy/
UgEwg3MPnnEV1eFZHh0sxIFnNMaL9Xrnq1HPK+wRRR2mpyRPHZ0q53f3RW/lzwmN
RzCFjY7hgjyCi7P4xWwYJts1Msx8dabrOrac54rlo+3U1i+p2j86Imb7B21dnMX7
QAEWUskyQFFfnY9O4fvFKlhx02uucDIKhhineuqTzqf3sxQiRDcoGZFk0h030D67
oaaYV6vcue/hC+J2QeCkBx+hy5mH5NNCNL/TLpAUyVI8dzS4o2ZZpMeHuOy9V+FF
CCRyK1n8j7l3FKujfMolGOVmSDFwolRxwGd0HKiVnpW14JNaDRcAfdphklNnhQF7
qj/g2EiHHHZQTPGFAS1hA+B+eNzw8WiRBnaxJOTbRTGvRk3CsQW5VRR4fhnFQBBz
uJtiowiBIjiyQVJN6IU0GV9tibg6J3FT5mTKQP+4eDXoCF5qOEI5lVLrmrxQD8BE
0HjNQfLZc4SUACUU6+M1W4+Ss7l3XbV9tHOusMxcj30JUo5M2R1ol5RNSirB1n4G
SCDs4aVUA/R/KHjsO4mEVE+zRenaQKqCi7PG/cFABpZu30angmBwaUuimMesLngK
zoSFFpEgKq1fVr4kdSc67vGxAdw3vEXaCDmpGOquvCrFzFRu1TpEslK1QeorYZgR
wYzqk2934uO7YuiyE0uOhr9K2UjgHTCK0KE3VG5YxN8ZzU70lgO0MXiqIv0nJfiy
nNUfOL7MEiCQL+tgheqsjzoz21ISuRB+IeRSFPQcO3qkCZUu9oh5ROxwLSmEup5n
EBE54uoObxtb6wu1NPoOf99wEgq2NHesNCrSRXitUY4L/Qo8ZCwYRSz5/DVTYmD9
c14q7hba7iKoJ2ywS8ggQlJPBe8N1/UKJ74yRIghWp5KNsKoFzstv00qOYOuwK4g
LvXBVDWGVj9vHQlyQA9XMjht/pV9Cob8nZTzeId53iViyaBFYQBFM/QlWgRM7Qz0
y7jtMc4pradD5RQ6Aql2RmGjjVdF2qztR+0xO8TdfGVjfKYpFxJo6Bf/U57foCsI
IXHx4e8G1lPl7adz3KUbkvvyS+BVuesN6s5tScZjjxU0pmMEWLnbE29tqhlG+be4
zTW8uW+knI7OD+v7hiFEjlJbAk/CbOyAPqUtPRvSr33lebqDln+TnOtvtUOdpTg9
ey9lKFiJ2lmBLpbZ71gtbD68MWHZbsqA6+NCdcJ3o3USFUk7TEhuG0ikbwh/kExq
Ya8yqQBv9YUFR/6aufQdUI0xCXydWUnxPUQKHLzzsvMWTJC01zqmbyH/XIifpvUu
K0dqkOuYf0daw3WmzcKgbDmRn3lkkKlwd1dr7RPO/kyZDgO54kWXSw0PNrjQyz7W
FE2w/kriX70y4luFY159kwSOzFVTBqqj5TdiAgBOTmdDCAjvDd0EnsaSp8gPGj3q
+d1QbzmPipnXBM7N9+Ak6rDaw+F9wy7a8ehmfcrj64B3lyiV8OICN9qvNEQDtHMR
RuhcfGMwb6q8TI3ViCql6k3zhy4b2Z7h9zZ5x+3MuPh4+VEBOeS5vcesJaPtgZDm
3qvnAbsbWmCMoc6kNDLtQub+lXZkjrzoiywV2adRlKq1DmT8RrCFXPPAU2uXMl/4
VwEsdRnoknyg3TbvSubpVdOVuGf9zXzefsjitK6OgZJjzBOlJ7M3JynDhIzICJgf
GEbitA40TPUlqnbg6zW7ukybd3IGxHi1TtuMPwujqqKX2xDg2scNnBPOdHpNynY6
ynX+3QyrRZK35VQH+6V4gUvJfH1MBair9KIRpt9rBlF093mWJxV8ohFSv//S1b4R
i18KTzfQMLuMsU85Cn5hgX+Nen2pK8QSX2x0OQPu1kNzn0x1TCjCE5DCg8YskpZH
6uai5VFXj0bJ9YEHm31c1Vv8Oy7e0+skfiXgYDH691ZBRyS3MUBmKGjJeSkzA4OV
sk3TbhB3L7MDiP60zYh3IzCGLT3t/rRngqNEFgBspf+OHRhgC3nfbQ+pHVNA4PRl
b12jwbXcVee3dXK/adxJ7eELt9VOOaiHkPzwGTLg/YP1pPcKQgwukeEaDhjQC8Pf
tH/PpdSBHYdMLPq80vsNLYUdTFxmZ/spaXWIL8urMC0GaXbff8PBfuU5eFXk6znM
AuIkFHkpxFo92CWfAx8PSuZtiHon02Op9OTGwVJL9cNkwa+hkx3l66b+lfxc2tdg
JkwUOp2RAjOs6kLzBVwzRP/0EVa2LtLhfESqp5/WrKKgvhhkRwxvtvjtClNtTouw
UfwX2fAZxfiBukS3K7t2BCBQb1hfaG02xh7Cw+jeGTsExdEL6ipt5jVXK49/nDnI
rYPxAAwY7fWY/5mfyW/GbTV2vu8YBTtad2E+1hbene0Wx6Fh6qZu8kYrBhpcJM4k
Pi4SHFo2w3+uxvP08fFvLpPGzisiMUW3FX9KnO3ZAtktku670LVvHVT7GfdemEfF
XGMBaWBWIdvzHCuah+ujmhDsCc6uxZv7TMxhR1XqmV0dBuA6Lgy24rrFfsURgDvQ
f7pZbC50do6gpgAxjhkMv0/6sOikl0o+BMkAyQmQ1EiUNoENDtqyG5Mufd9z4/ti
hEv30syR9HFE6b5DZ8b9FQ3+o+cqVs3YSl/7QHeUC0O71opsLLCJ6ChMDEwhzDnR
xIlcp9Xb+T1YPUmXxRNhSlA+Qa4QPqNnLAtWJsfWaPYCtvkJGHDSaixbZlUDkKKT
p6usbj7M3KiXq6FKZmah+TACH6NpWqpyYQKWV5EEzl5B0s3n41bc1FBJ3UQHNj6s
ZyeKxfEEgnFemK+3iYJMy9YPhqDvEUBLTTCZYCt4B9jDwSQHQ3P74KuE4IP3ej7V
eVeAQgaF0WgASunoawvrEJEHsAfQjAgNFxlGaMmSWpP4kKzMJXmycbHNl50V/yNM
iDM54sUMhC0YBO9nyGjAdUCDehxitumbAs0EFcen1VCtuEmnR8+QwFbCOJsi3Bsn
c0/IiLqOmW5XV8OZMGYZdQsrJncOXdlCZZ7Z95yZinYHBFdaOnG+S9lSt1QQSFfj
2MCthO2FYBzRfHf+mTKD0UHBCCofzzcre8hz/vpt9oJzbMFQl/pz2rnpaW0xEfbB
RxXIXoMrKKiggU/kZyL3NuQ/K/hzAPqWIeozxjO+QawuqKalu99H1Ur2KcHJjGYv
WDYzlwhidRLt8A3mbDg7rd8Diw6Qz+mNILh7zwLI5mNOE9coxW8wopXengpSfgJG
ci3HNWd2Ca8ci/ZBigqpg5Du6dX2F+35L7K+tFSB2JCLzI/IsZsqMCA50SqCrlSe
Aj8MgMUDvrrOSF7ESCMEHOLqXcjY3UJkiXy/YO07FwDi2sSynmijoQgJ9n3wNsJZ
RXwjKEwkvzhvI9W6cjqCOgzlsz/2YUWTm2jiOjFJSYjn9asan5mb5ben4wmMw4Wv
i7rjv4h+sp6AIfJDAFRViF6sFPwdy6GDcNnzBygeavKKSav1PMCDJIEvb4ZuU45A
DbtSH5IIiEsFuUsaxwsNqqT0Icd/WhIdrwsF+W4EkkdlMMI4Om5D5NveHNY5masj
L/djx51u+Sd7XNjJxmbpvgsby7DSo5SOioJA6hzpHyRO4LQkXKG1rOzjTjrwcG7g
UF6alM1w9G4TnidwhbHedvEs3kiDwavVSi4wvNQGmRMaQjB0ORJ1aoqv8Ae8xqcc
82EgCuptnsV9sDF4lyVJZEJVzncLnDLqjyylgofqU0TSRjiAvEMKd0Exp+MnQNoU
ve2GN++pDRVJM4KHkQ780udfYXu5JrJtCJMHt4VLOKX52ueQ4HlzvJUBfKbx9lzt
YnnpZY1WVax+w35/VYHdJGw1j/F3hCHBdKjavd3uPuZGRMdm32MBeU3eXP821cKp
G6SeH0Qebejqnzk0HTAkJ04Nv8OcTzMFYg/LKBk4O2gfgswbcUB8Tew3dE1aNVf2
xYTLCt72+gm5oVXxjN02LpwWW3a2NulZHmOZyvmEt5OeC052gFqRwPDL3PUsAjDz
rwF/njkUQiUsMBfH5kOB6eCmugRzs6dS/2qYw68Bp7LQ3EL7C4gO/etArJDYIKP0
2FXOVG0NyDXvXD890J/UNkGD9tC08e6yKJeXNAOymGRLgDKCKumTAAnteiRrCEMp
dn2RIpO3b4xRV65czcMHAQaA4+oxzZQ9DrGmGHjGV6RfHblPaJzUIfIDm1XXbrAb
Osve2UB2R7ImKS/as4J85PHQ4HwHiR0rKLP1KA9MQpddKxreK5LAPEr1aV5wKJ0E
qa/bvxJ2bHH3lM+9UbStFN0IKRKs8pYQvtuCFdRPn0rac9Sa2z9VmZz3J9tX2mr5
G2MfLUwrxYe3mgzmfuxVknRmTm3++l/o5X/kTyqTuFJIVP0NHQmBQzbUrnD/ld/v
5W+nfZq685CJ3c9ZTQAagvR10SUKK4+aU6obbNNJX0D4FBeB27STGhByzDwF8TIr
HQVwqt2jdRjYDwOgI7E7gTGKH6CgEOrIi54UKwsZR6kKIhMWR4a0CM39xzrAjb77
rIpzidDqlNhXkdhXJScpCEl52d9ftzJnifamAWH5QLz6xaxmKrWHfxQqlMQrXLLh
+HLd/ooqPVk7drKPwFhGdZLCKWohbLsXX6dpEH5gXcicSIKBoTDbWfyiyNE/3Io6
CVotDoKKB/e8U+TS5nzJ8WdecxErKwOVwF1zK/sNYKOCMvKGC73HAoHlH/b0Xkol
vu88fm4NdANavDlEe4Fcqj7jK4ZFTIHbA2EFDihWfvBVDQsECxx1ElVGfG49aHm1
FDKe63wxypSMl0KUEG0UleO6wBeymip4rwUgEbWj0F9JD6ZczeJA6M4jf7KR9e7U
tmivUuIbzuoQoU8uQXCwTe0lruz8wuDO5yXJb8+4RJ2HECfdrpx9dALxLAtIzlSt
L7Myo+kXsTbfyjOmnt67AqG+5N4h7HSPXICHMwfWCUByrd0RX8q9QTknIb5y7Bg2
GDP3IylFUmeESnLM5XhCJ2ReMt7RlggSpvJywvO26B/wRqYo0oP5Fm2CNceivU6b
X3LmBfPw0r3QXiVHh+j3oidB6nT9s93LvwV7USTKn/Dp6lHwmTtPPIW5ZEivKjdl
Fp86RJ9+iKvI8sONDm+hqxEluXsftzyt2AEjtvYFQHReXuEbByVSxua0Um8W9w15
SbkqdWqOFujrz2O5kNdhqTT1dPedK3h2u3TojGOJP0/QXlg7+9SnUex79i4Do59v
OUby67+FHV+j8JwW73Hq3mAkND2hiuQPJe8uCcykOT7UbaM8zc9Tf8uzVXRVl/yO
cDesRcGAp5rOQrzJdp8OC3gCZwVRuil3r7d5npZu5/0h0oSaV03Q/aVE6iq2D/aH
bK7rHQBRIdFe+vjsH2yD3YkqJzRMUBudaNuxyhSoc/hP2VFVUIFsKGHqFVFczTaQ
OyG1CgVQFVPc5FBvOxDfq8UzGEO6I9KR4iky+KIzKFY/iUJdand9tQgPb17KIxr8
PIn9mQzHYRlUe7jlKm2eTQOWQDCevA2031LqZHUnUTX6x4vXq+ZDPFhaqxRqFmkO
+ewcfsqvOuhbYqyj6ykESANY3cOQmjO8L/b2npT4GuOrpVcnQiNFVS3tWfZPLZlP
UXW+2ie9MieYeT3X3p//WSTYoD8cSFLGYUGfbWtyOsxR8WAJlw7l4fUByfFShT5y
onGS2tG2I8AvPICTlngZ6GWU7bmHkoNu9gsFqF15ObtFLKWFyXLlpdfY/h+/tJ3c
07ad4Os6BG5kdxjzI99NOw7Jw1fr09M5jV94AO4BDysCixtlhDin9rBrT9lvACNe
X7owO0TSfcFlSH0nTWVFVlgqlF8/ZQYa+A1I+wWOUF/53nqTpDbuT/SK7r2YxkFP
bLqE4ScNLbRa3W3DK7b9AoIsT2JTUB0HoiGCk4GSZLEsSOfuCLOYs1oVwa7RVv+V
cKefKRfmgSEKvUwudHIEVZxLDNDaSDNSb5L5dkBbyZ3as1ysbRM9Yt37YoX4GSor
SItmsAL2SNTtBnxdMpEWwyJRE892FuGF+lGJAQUwPJBaCYL6dHLZQJFUZHSDN5kT
HCBDQc7DJ2eQbjfhUHEgpDyaH2S80Abnorm0hIWviMUdtlbm1uRezIo5NoLB9sfH
piz1yj/h03qM43YGV+dpl08bx0GzP+n5FOAtiVViJHjTtxyxgCqeegjdaA2I4wXw
0kdv7f7s/dXIatcyFDsTDqqcTKIcUNlcJHPX1gytwxKX9RPjoj7RXTyASriVKcKq
ctPL8PHsvbwa5jpAJIkYNj2GVujGQotSvhJtmFPk/PMYbNItdovMu6r1dO1FJUI7
Hj6ooYZOGIE37SWZEhn0i+aToq/YliR1zfwdce8ZRfB+JHxtUjlE0dVKYFEIv5l6
D3s38OnHQqWc0zUiDKQaBH1uE7JOgvdwCiHdgSgkKM56O8oLdGJy1ZJ6IYK2hx8w
tFOZuTwyy1oGORVIztnI0A6E2+dXwCTRFvgVpq67Fr3Gwbpm7Tf6vtjPFDpsofN7
z6oNMwyaKZvfjq+kZh8XiTsvkqc7iFF1D8geSln8Vs9GUp1ST/Pql/x8pLNcLCtd
d0e3I2jg7og9uYrBC9gGaryWB622aB32HdBb6bX95w6SgOfzDAWaDiVUdf9SFLgx
PTNR3nFhfZDL5nlTwhwxTFR3JLkJeUx2WJKdAsLOktUDIgu9a7GBA3uUqoK7UFpM
7KBM02XgLqBtsVeZx6TUqsQGzM1unapcHkDcQdarZgGSGAuf94iPPxKgaMEVEOHX
zCW/3KoSX4/PPAM+sewpbSqY425SS0d2MVQQ7LLCggsIJoW7b+CBaBNZaQipHn9d
0ZTZVVFL7neQqkX+KAOhuGxE646pOW4hsq/t6yWkisW9Wddq8FxwpuuF4GFLoz76
iNJhKKCk+0igr8E0auZ2KOtWnQ3e9rOSkSimKauuexNXidBMnoZhDhc1H7lVwKHH
FzgYPhPNU1zFUyMM/hTmWy1RIvgTcPhF/h8Cgy6zZO4F8Y9QexUL8LS0dp7rABwn
AoO0E1dTKThzZwrPrZbHJMzX8uA5o7NKbPa028vuGuxzyrnodhE4aFk+blh3ZL4Z
cAFbaTt5P7ysqrgbaF1xjODJtb3CasXRVqHxs/bLAwg8IR/cwcIOfX0EAylKBjse
pvL5CoZA2+ZV+z/88ohm4rnu0RxCDasx0cZdEEBq3HYnDEBziuCz8/JgNlmpt9/m
0uWoQJ1LvAKaGU4ER2dIzvM8V/LwwVWgKf+l3XbyXKE16NtaCFY3bb59mTB85ODp
hG5M64lD8ZZhO667atOhAKLR4Ir9mKxRrNjRS2lCHQkieNZ4yZWQyMmFxfb06r4n
vGFm1ZD5EZL4apUJzVPx1lbA694Epq/ii28rU7HCaM4YEHmspjYT6BCtXQHko3Ek
B6+8BuRF55hJkGuNCtYXhHOJpCDHe3civMDPeDj04JEMLHf36NrOX08rdcIyVIT3
wWmJ+4Abp6W9aBmEsRWQ/3dLkji+cemUzpiG3pruV8Si7YxnTfewxhOXqvehZhkR
su5loDc2Vn4p4Pac0PFnB14O+JaXtjnWYxeM30l+orbsEa14Tp7Cm0VOjVAKiv2s
MkfHFbcCDa6+eC8YYgDHKk7OYDgcFp/VOr/xMqvE7+QontrTCm5DSQZLTWvd/8dn
2xGiuq121caJ5oAopXlaeE3SYruwJk9AkEUPmlub2+WbCn32uu3sNVm6UwZJO//H
TRbeUJAqC9vehMjF3/jtO1/pOohz0YHYpjCqtGyaes2+06Gy6Oi7Nq4I1wh5m65z
nFZ9B+0wiVLApHgTa/84KDsR+0pLzkymIZoUxyoo35P1c3/J4OmjocDhXmi0xYAn
rcgSwMo98BxIXQ78cW0U7/VAzypJtvX/MZHszlIu33QhMSbRwBM5l98ypvUn5Xcu
PR6NgBvffHmVJkGosYPBDQuk1R/dXSsAIBYmjrYFo0cYS3GfrXBrwm9cTCGoeYNN
0r9fbdlXjT+HNZf8NVMH6thVc56Ol9BVVySuuSE1lUoUT4VFsQE6iXW1iXHhJWvj
yGmrd8OyCrB1ZKs8x/HkGgudxp3YyhPuU6eloaZ/oH1AN7GPmfea41W6JTeiHxmT
T9ywJsshNSBE0ZS0VcXymaB15FW+SjS3e4KCosF8Li2U70SHXnD3+/TwQY4CaTBO
bCx7fBiZFgz89HUXRd36FfAwtdQIZDndjSMojRkztmFS9PSQmTvs7hR2F/7o7Ah4
fwkeFDQsaL5o4IfkZE4P8D7RilRS/zHLlZWeIojIeyNERm0AMNhkoXgcN5+ga4q7
NqH9aLQcGCUioUQKx9BWYyjoFtUdf7R2U1RpHrXzttGoApL0pq6T/gw04/Rsxb4d
GYL9nk2rwrmBJyLDs/oNggB8PL1S52HtsEEvFLbE170nzfAAnEUUqjzllojERdrS
ztx51uqfjbY/UmBdZrCbkUit6K+DGpQS/ABSfuA7fFs7b+7Ney3cAeVpfzCh9Op3
DihDkX/EZrSdEdIWXJMx+ua5Lq0vq+UDyGI/uYg5LhZdpVlqk7O+PCALhYSnyPk0
j0Jnfxdlr4YHSZpjm9++4gbK7B4InRzSxJ1Iw5nk/Cjs8duJ/Bd8UObf99/S02Ky
SHiRgqJwfHXf10of76ydez+bGWcvWTFemDvyksL8qUYSDWw0GQVrkLOfSe0kowtg
2zbIJFus/mPS1tWMNJnrnXSHsbkh96U1I/RIZrGUbLJro1FxrMLKAu8ihhqZGAAQ
awU3iM1mB7XXbldYrefBwTe9izWaTFYiK/xoKE7Wv5bIxc+furBuqQ7eEFDVeP9N
l21gzbHGS6SACStwhREGvvduAknnzpmAo3zT52Svkat7pqqo4qmAs8qLR8jTYVh1
3wrhj9098qmOmUDz5FPPxR7TFBJyMcKiRpvrKAtTD0vCexEcEK9Gu/kbOU/2tBMS
GxicHrTtElQ5bSE1dYiL6O8V+/rHyqbSti8KifTBIQ/Lwdu6ISbj5mZQt74tzXIh
eTD/yzrnZdf8E0255Hm2I+KdVlcJyDTS7QZe5dr4ogyFdhhMtiAUsse6gw+plkWz
63hvdm8DxWut4lfVDcdGh7PxDFzFWmtRGxbOTYo6N1I5Ilzlg4rcRfakex4Ti3xi
piGIrE0M3mSI1uwZzseqLVFzMo54RAJ73y3ewrOfy24pn1cv+pqLsDrzaL4hPoxp
qXWeg2WnXGJMO3pUW0r22JoRCslq0pLiUBZSzCZ5OG8ZZLCEa8FixKR48ndoJg1D
0SP5wtvPh+JYfKjD7bQEu6gv3AmBHBHFapXf/8YYkhjmd7F9HlhXeuX0Y67pOrQn
fEemPiC7sHcejr381Cdj+vf/A/tHzdML4FWBGxUYXdBo10UTU1iYzKGIL1ElxKsH
jruuffvBJ52OzFxQvDdlPDhDko/8UVdrtzacZyImAqsqGIUSLPVb2ZdGJSp9Q24N
1aMHIOSqldT8lLphKro3euY0HEAGgtfc9SEvNjEP5J5EzqjXbf83xRU5ReEen/xA
nuKLywinqMRX+ZFOo6BD73PIhsdpZs7ZbDcHKWflxYXlk3TU3Iajw/hOYi8PtDKb
4PqbHUdTGN0AqlVWXYQd82lfGf5H571x102HK4L5Vc6vulK5ynQrY4UMni+zCNeh
lhvtWUUt67c3RWlZA7AsaCp1LcSnMdri1/4tTna1YI1e5eNsx0KpJml0iiMDCn/D
AyKP0/tFiwREvjmFD31HFWrUM4P0kIvCln7e8CAs/O6VMUoP0aJptnBURLde05YC
ZMc7Oggv5GE4+ok9ESrWQPVFKtdoHnSKtoMlLln6TsKf+rjTqoiABnCvLWUjtR/o
i1Mrlbt15m/8h1vfRhI0CYd6djlIOl8GmUe/YWCDYE3FPTlZJsIrs8jE4v13qZnQ
99xVmzgmnhp0Nj10+aQxbMQqtc7D8o2byyeXtD+uVW1DHBSYDfB5OPOPGN8b+4jH
wbarxZowwGiHLJ3rSerl2KRDX1cX9ZnCRGRucsFf55fSp6g9owYyPwYL5AIqAke4
4r/A6qIhVwAUfEHNDdUTgsKdhe2eVeRa3sUAdJpho1vWHGruDUE0KsA2D2XBIJPP
B5jySgxbzfUWQ6HT1Ydp6OaGaB0vvLyEnjrWyK/6eQJpGENQeS0utOz4VWD4dvsc
bbBCLvuOKy/VqTU8RGxclph4rnkQfxBXtDV0ZmqXf9OqlNsSFimN2+yjeMPzzwnn
IkJC+89WEM3iAydjoX0Kq5bTKJcdzr6fUKqDHkOUoBqLR0ODBnPv74IiZF6fRSV5
xfunJ1T6/rRG8sMIRn6wkZUkX7odqlOkr0mViD+H8I0UCOXdcKkcfyHzo1bUzBEW
5I9Ttx9CWS68bwOHXIWdFEsO3Rfk2fBaQk1PojBKuqd38/BGrds/79R0635CKdZG
6ccUZjjcCqPtbxD7tJGBZA==
`pragma protect end_protected
