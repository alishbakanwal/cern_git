// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:24 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Owr0UTuHuK5vnxchQ6SXlio7/rfaHtI8mHUs4h1kCNtTeGPJIyt8ojoWZ9VuW/Z/
glA7O06rwqeKTWjeZFxTLAxSNMb4N8ttODfJ78c2K0f9G/lAwP8D8nVMcHLFL7y9
4UiDBFPh2b3lA1H6k9iAsSXR3KTz9cAgDjxiK5fUvwo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7232)
c6JDbkbm5gFkGe90BTaUV/CGI0urIDeqKtwp7IVu9w337siOBFqmK7uFue119WrR
ZsqLtrLM66xRH2ixrgoivCNBwT/4AFxQcANGBpjKzwz9agZjfGAfHizJ/b6CecPG
IV0vR0ulUYShtj1Oxjab+P02W3sbddGNfrU2HHlmVn/Wu0HoywiagzizfJw5HnJI
hxtTdAPl5Kdg/IbAe6zBUsFFUANoPc3+1MEv/00podvTbA4s5/Gw/Q3PTtF3DLQ1
D97ZXINjYD7PCygt+Amqevvh+DIVkSH6QknPUWwaOf30pkEaypRby/0Gilr3Wsbb
K8rJwp0wb6U/TZ2IZ3F/CVup5TbrrhAm9AMi/VMn+RZi5YPYGYGXeog50FhEXYwf
yYA3vx/sLR0iY2moVU/CZW+BzBx7WntTKmzmUyK/CCk2KwCPovSSOASbQZLxd4AP
JjAmjsLe/DFA19wmp69fbMKXlWyVpiW8dzIYZk8rUGjhYB2QFtHWxII0p8EES5JY
zQmIvUh+P6SNatg30d2Job6/b1PymUtugWL+P+zi+xBVXVlpp9+qqoS3b7URiTbu
FGb4gI5BeHZ8u/s0mtaLMMYo5QrniLkb/URYn+TxKjJPfIJlBJReoTFVYV1g+eC3
4Mx5eZEwdyz5yeFBB6QtbkGz+fmRZ7Zx7dN7TxkkEV8Ho7R9k+MRyDLsNLjp4BEJ
NxpWo4U1OLajXp4Io4JTGZS0yXIcsNq7jcmKTQuWVgruViibmiyezW0krzvJuefX
lYoNsrvlwjRKlZvQmouJW2ioGLQIt6kZhVrRc4s6/4tSJXS9HpjzSrRzYwHlgQ+e
7b4ABrd/lnXXw1iABaLNjKb0uDzY5W8CBhnOuqzZM+9XZIeczMEj+aWu6VDB2/Qh
G5EtTJZH/UX7MIHhcbkhvW8VNwB0YF2PtCRXLZaDWVt+RXPhvNKjWEbGHigmROPm
/tvz5WIIcZroEGpvtFUo3zfhnvwC2ROjXBSuk7ztMiBr6zkrcU4NfKsqd53rbgru
lNY0Vse7KW9mQtQuMmcgsWwnD9klBdar+jb7cghIaEEt/LSIUJKqFXC4nKo1svWL
YROTzFnE2JQq+i9rqmUKHdrNKMgU7N34uWuJDUyeLFqG/jKHdXAcG0GnP0D5bB+k
CvCp7B7ioapXbX4cJUBiYhj6PRNsiWmPTy68ZVQxuNDnvGz+vDO0owkg5E1wW/cI
595pjHJo1FKXoMC8Nz3rn72DUetuDql+OAN/hHehztwbzqiod1sBAgBBsE+tTS7K
gPGnCna//e/aaly6Di/W/2omyFxY1HOHQ1lo41DcF2otcItGBTi7GoGwK/1HCxu4
Bps0BcbeWZXOZfbyBVHlpCbnUOLuHGR0P6ydIlapJRY4J536A4I1ZJkmwqo5ZLWW
B3QYhJee+qHmJ4J2LQLLJbEUslUNACsOj72CbxDmzSe+WL5nR7lOL6bhbPklC6jL
DLPuvcM2aKPNn79gJ504LWISOqPwwHAzJ1VD6qqcC4Eccyl2Le3p64qvMJao1h1h
gagZYN0jAGKDp06BPC7TPzRZG4bdyos274i9P1UwVM5Wyl7g8BPifx1uOZ8PllSq
U/6d044Pjd9y93VcffPL5srqBVJxuwNS15YgoVteqY1sgfeee2Yj8upXfj398pvi
TOpy3XATT18C189xr5mGOIe5CmtDjwHM00BkY/o8msU/UhwWr1bVAxC+QkcBlplk
658lnkFcscQ78qZaggEutopMg88YH69xp01yo2OO3lQ673pYvV4aaRciZ7tZ7GAS
HzDzHUoKT3kJX3gk7RC062L7L9BkAiK8OlHUdqblIc6uml3zeMjzjskMirz2q22n
fknv8/n0N4UJRUxMn9t671i7xHRmxAnXNe0TaY0IgXMvxdl3MN/X3dsTqf15BgWt
KiTonhrRBjIKsVhtLaT3WFta0XC2B16hytc7bfSAnBfZf6vwFuywjosag4e9MDUC
JBfAIY0eF7SSzhSXAK87suu8nhchTlzfRP31QckOdTJZsRMMhwvGhRIrjhDeqeko
lvTCutCwWmC59i6TGSKcr+nUEpOeOSqr3gbIdmZPvwH5XKKHy/ISnPrJh7VfDDSj
qbG2y3BqYWMcoBGJ9F6yo/ICqHzZTTjMWsNo1E+8lAgrc/cDsCeebcq7IYaRcG7/
7/EVINBbxqgE3okpmgwiNKaWhnhCgekLVCoJ+LDCvYrdkvjSLvwtcj3H6QAGKgP2
Ic21eKfcd4kCwZj5MpPEFXNckW00CzT68k5E4Km552lIyjhZXw7lPJIJ4lBIdZS6
PDFyf8p54HNOEMUtB7ZQvsfeWyGDPqjeRyVaLoL/RxjMTY/GeFOryUkGXuwcE3wh
xW6SyIcfCdxQMyS01tTxVu+ACzMkqHWQITFBrhwU2fAzfMDRJoTCysBTNAn5ktAr
CdNmAqZ0K8NLN4OIUxE5OQZqG0kn+2UD61Tjvszae6kbNGXCsJcu+sOiPQC4OTQ8
V8CeYJlGwNynpWIPDWwDi3lTJPFr+HmaTbwYMayf6XOYP4iMZ0zWawfpBYRvfQW8
fzlDJeLKXt8w6gQjvkvUqifz52sQKcXyt4BfgZI40ukHBA6NFWVb4min9tZJBZa1
Ch9YAHDTTn138u8OGTGniy/X9yGBlzZnIfAmO5o0mokOhXMvGVH1UW0Dtv/FYdE4
WfVINj9ahKhBr0aANP9WvJ9AOERnIM8heoOWk0jKkURgaF/n5Jzm3cIYlOhi2+ab
87R4LLjOeVb1q50b/a+OIzIW9usvb31/hLjKaXR4jpcoX6CwZaT9NhMSyM/QqTUd
+M2eQsvP8JB+ktIUigR6PSiUGaUffXg39eDdGBbKRP5eLwNgdZLn4dd6HG+1JdIM
zXlgosppJ0j4ngUG10ul5emqHUbUNa2iWtlJgOUBpkqTrGo4L9nWbjETjuwMqZ1v
Yg2WaAXQeDs5B/xJ5MB+vkOeUSKNPv9sHwukt1MYkR+f1FhF+cRv8Zm/C71pbLB3
Qfl6c/r3waVd3LpNAg5Cm2KxzDVVafiVOYh0p5F0hpSkjRl87hXqG6mqtNj1xIQR
017iuKLB86Sy2+zh90CycEyGWogdRficUNvavHoikolaXD+HhUlKQS/71D/fFaAS
8J2wFnl3zGt63CCV3F6/Whn9bcQzRbhCHXgeHN5jo6FYeHtzg//EpgeRyI0kpff6
qNKguR3C4HO6OD8kGbOERuIL7laq60XQQ/hU1VO86OL1g28yvcrga+oX+j2SyQpQ
qsYJFjREXBlUvmxc3PDnbg0PLREKXHi49YMGIe28AS1RjbKT2xK+Tw3NtKwVYv4h
pqJFcSVPqpmo0eRNQw7C6i/joxIAKM7CFHvLdHGLpI5rNoZuRXEOeWX6f+LfUmi8
UOaUp9Xu8BRtJ1/1/qKlFIMxtURNB0rX7Zph8LzrGxjeqfKvtMtTE+ITWS3bPoU7
ZGOjb7iva3Q21g2I9kNUcDBtF9TQc9lo7UpyFlKKY5JjkIgZzQjjz75rBtOHqK8C
eROZp0u2Mfs06aXsKJXbuLSefk4I0w1rRu5PVMOm1dPrppmY6Cdpq+tbXc3vZ5Q1
u3B3pNYGmmhvsxdrQ4ylgarhiewObf9Ynn87ciYlxgGQyv51SqNOyPKS1dKu9DRE
3sabYXmhPaRcD7lJ8HUrotPVg3autux5hThE6RrJmwJLzTffTiEZ5z2/dXsg5zWy
c2urW2hrN7dlGHw2r3Zre5BuqvnO7WcDDF08AXua18RpAabCZrsMJXI9TP4xoaiN
WbjjSFn05aUvq2Kh7HBWnFMi4vB8DGC0ApxtzOgtc2eygccmg62Dob5bYL9W89oJ
i7s+9qJ5njG4MwEV76bI5JTYq73zd3D2RFiQyLx1eLHTOULV/I0h4QDfYFf0dLG7
mgzuF5c8N6YAgscIBDlxZbTgdRg+MgfyfXAZTzqf09evvU9J5OLhf/Muj3ZLlaaQ
GOx9zAGlYYwf03s+h1DI30hGIihpBKpsuPgBhC7X0/qX9c3op3Gw+YGrv0hISmTm
bqf7X7KLJrJ5R97spmkxTA80z7uv6Ew5qTioiPymIfHuYM4vObp2iCMYpqKBU0c7
omw1+oT8Mk4ZY4cNyN1037gwdOKQ64B+OsCcjaB/0K01kf+xoMzsgVJ0q9BHSczs
gFFOD7doklsYcy6F/SBNTe9zOL8h9VwgQ/crdlHnotfBPARvaHo4Ag/nsXfT7mnz
7FNe9bQ6QAxCZyA/P4zfGBJcGJNYdcs0nHpim0hmDSlC0FsiM8TPxOVRhdKXUj5O
rSttrrDzE8a2kpFsG8BppCs0TmDAyEEPHoIvqYup0LgnIeqMJRIPaJcNvXmE5lIf
rbBZL5W166KyT8B9Ly++UMst9sUUi3MJdLngyT4wMWW1GQy4fu0etKCE3VbpBVQl
ihvlE34nS0Q3gQZw3B3vUkQvwZEEMjIinSMRSdx6yDn4hQecoRo7Y5FBbCVjRhj4
aj7b3JtRa6Y5XXONu+sPQLz7jVeCFFQjolIDhbFms6xZqu+tZGVz5U+4NUWI+jS8
GG7Okh6b/MymooBBOwjkX3yncOM88R3Isbf7fBfoDjsmMcPPHmU/T8OaQgtYQZ54
HX+OxzaQWrrYyk3PllRI5HfFQoysPILKfPgZ+OViVoS24eSmkQbR1Onohj+WMoJn
p7rHyJbO7MvLRpAPfiV/ogi859/0EDz9uAehQ8UAL0ZCCeKdrJ1O+MXHx/pcXiGL
/e2QyaxhdKcMATkPGAdHyV4HNVMbAs0tq3Gd1VHgRPkYssYDxeZ7Kfk4v1JfIX+/
0yq0fmAa0uSSNHB34xGn4daZ2yXp9CIrRVymwTR1JUnT1uBV21pxz/3Z6YQYfDHI
tcIJFLKhkZVKQXzWII8P/UQ6TmNxhxJvzjB2ns4A3GW9GxlPckUGkgMGh0TpYUdl
KtEiwfM1LSi1+i/P05EKG3bFRHqa3qY2nSVKARrMmeseyN9GJq/HnsJz+VS7vc7C
FmhCKIuh/gwe1StDeKp8AGcBQXsCwr6Ad7MrERyZpZtZc4oxUMSbQEOH5N1BWClZ
AnDtXzoUZcAevvmDiRZVzcZEZELpSolrpNKxLGclI7DK4vXptzsMAL+eu8pG1SQV
jM7tUOJ4MQRv5m/qoR0DOaSJR8eM4z/VBUhEsMLA2H0WYd+YGpvF60Lz8l9bqc/K
KDatZQmBD9aA9I4aI04QeMxGV6v+9suDJEsjB8pXzITnFjtkuUn2CANYRbEkXvTs
STD3KjcCFRrXQm+5IkOywbLym7APHRJeVqOdPpqVdCwXVQaPyZX47ZRWmTVCWuN3
YbySQy0CHtLktCpo1HPnKDnsPhQnFNn30YQplaIjmFq0r2zhz1qGuoIskO//gEVm
U5Z9EVeYmX9Xc2i7KwdDxVqISYlx+Rklu3nxhFnnRnu8h92Lvf0EIeovrDSSqj2M
Lx1+3gCUsiAxJ4/6vMSJ2lIu8/GME443yzSq9LE87NkTY7fZCqHmlwyKXLiv2fxq
91BPlCiN9G0y/uTKHiVU1m9M7+rtqp4KPXZrLErjmnNaMDr5TojhI1RUvYKK4qxv
CI9p8R4+PwmzrjKN3mEkkmD+bJVQiGr67pgI11GR/vTAcOOF5aQjBFlUxqNnockX
0Q8sJtYq3gpriUujrfg0+uRniUZi2+NDDEtiSbeokUNI7iu6dpKB3cdODhPqxp7O
s7kt2X4vBisiO/NkWmuTVrwUllyPxm7aoGcFSL5dqmgNIeGuK2qU0deJLzacLkKd
JwgZ/S7caL0V/RrF2Oi5qn5sXkHBYd78cAs38pmB5LdXXuEPDeIFgcn/TOvFmdEc
4U5JDfWHl+FNd/wr3GsvNpjuF6wIGGfjcLUMWPw4RTmEeuB7gDwgxPnUJf3TCCff
RXoIYRRF3RRB9ge2l3d4xpQPSs1ECvLLouMD1lWKbuJZrhXA+YogQBRljUqI+fT8
m7rbYdSbOg0S8twl7jOYTHpB6wVhEkItQfkoE2PHpx//P1TxiM1/INfkytdW1hnj
wQt6SozEYN0RiOH5dhMUjGMn560/Ep06viu2DpiMbrs7MfPeafjP7L65TkGUqlcC
YvaDzQoBX0kKwOfEA66LYlZfwW0klPMrh4CccMbCgVwruJ97HTr0EwwqJW32FcFq
Hs5mBHuZA424dHlwgUQ8eyJZrewkb/Q2q5LJDhkus2BrWebWtiqUcLejLRSallmr
Vd4TV4uPI7DP/+QPL46SuxtQVrDrgY6Xw2j73fGLLhMdTP8tN3KqRyEdtQrDok7z
8Fu/xmiYjmvC8vpsggE5wT0bQ+I/JXxkrdyDLEzqrb+iOYAFV2ldaL2b86OOZvgY
G+CYeWQQyzo0RTeG5dDA7GLMO6WOa2Fi0RvaROn6pIHZXs1cgeTOBzIHVwBb6cuZ
9HWr0ItJoNBsyXFkCTQ7uHIgCbIKQVfFdlf8bJvHL6r8ldLPnTgheSKkNZTpmDlj
ab2a8ihABJMHpoYed84hu+/uYC+H7YEHrPTY0VkB9gRj38VymLNjPhV/6L2fyLfQ
d29sqFJwMtYNOo2uDHZRuqtIMbUjQGSXifWHOgdDXoneAr2FyIqZs8sqsZDbgCN9
i5RGTO3FTr5Pa5b3AoVKTAl4CXflvVVxoP+lrDb2WTlI48Qb/z9FqjMK487t/6Qs
AZx1FVaVPVyKBz/w6U0UMw/fFG+CSk39ukKv5BjDE4QO3GkC9rdZhVpg0QBHiHnM
9w1zA0PJv2bw8smdkHNq+wT104NCg03d8maiaCeBi1ky1m+ebgHdqb0fee5N/2EM
QpDQUYj78APfuBPiA3xwdH189G6YGvUhRlVnd45HwLR2hZcw7tjvsRdP5U6TzcPJ
OouP4RJW7jRVuIKV4iN+80MFr9KtyzuwFDbN/oF9ZI05j3aywfXrDP1QW+o8aWEo
EcipNEOSpY56/HGRlDjuUMrDRWBIBvASaZAW0Q1qfwiUhKdY6XKxm0HH7JwGgsQ/
47wXEOmX5sk87xR9rJiabKteu6zLsQNTEWqG4XXdiL58gzxiD6IWxXVn4hTxMEyt
7+Z7Za+zau+HsiyF4pMEnNsPOskdQfTeufct022CpFwsAe1R89MgM6OxiaedgJOp
HxT5rucGOoIjgGSg3GDgW065V3HbOb7hdDwkFHXzS7IMe6cf3feQpQqP08mqan8E
+TIsl6HsgNMgcTsb5ElSRMMTnzIimF2EQLkqhouDI2hTSJrFR7yToVxoXFDh6Sz+
UjYO+vrCowDIB4MOVKHhjfhFPeaXu3j4oncEfQADmAvTaKHqrnrxzbg1+TE6Zvz/
tTp2kVZrNq9BEG/l5nunwBHzd6sz6oj0LX7A1D3LZrpdKUdy/FLBAcBEVUI6CeJb
xTN38MLKQeU/iGK3WJKvTXAe45RI48ABI5VBU1TLmT7ZXT45rCDFnhYrEkpKp7pU
86B1nrjJTFEYCwF1BPwvFyHZwzHN9fIlbpr1I08N0/O4+JEN7gFYJRO28JO0swnD
nQ2VI7Uh65vb7UZabYgUYeZXNh9XvIei56mi09DBUdmsPPLNNL8cOx34YSKvKi/x
mu67whxCwj+hoCEHBw5r7kPaBXTzW3iKOdYv0DM346/aLr6/9Wg16g7Bmd+l1kvH
BQg2d6IyphvXVGAFihYesEB05BWADHxO1y5ADK+fF8AtyJ99Zru3GzbJMvActJ8z
DIqQpaqSSh8gkCN8+6bAtJskg8CZ1XmXee0ZFKXId2urGBQ4LDht/h6SWat38yRn
l6oCtRoB0RiBkTui953zB3nShZ6biVMjn49xGA4xINtBGdRkHYh0nZzh21ybPVkF
iUEFHtlcHSOmtZFUmwzEdVcZsX2d1TVJdWkjbC76w7i8QChA8DtWqhxH82GwFxg0
G3EsYSuLEwl8UBB0LvBJ4xaPHjmKsBH2AZws7Tm9Wy8M0OwQ5lr8TDJAy/xXGTDF
0rD9DMY630SjSRmJSV807XWZWlBEMB0XfmRnZ+0pDtT1/EAGEExsyIXN8WbE66yr
EWIHb/Z2eD6d6fk24Y+WCo0l5TPWQ/oSrsdBQAYwIbKyNuX8ARptx5QATMklUSSf
0ZlKapymIzYCo1VZt3WcQ1Ce0/BcuFgum4fX81IlU0AyVlpWdSMINz7FLy3j2kIk
zUpj604M44Bt59EbHv/XNodpnK2lSEJVu1Te0RTwVDx50IP/WeFNTZDIBLQ/Q3yr
Uin90sNIdDifS6ptSS4EUDKiFZUwC7cnNvRhy3fXRCH56Aj3SLJe+X8HsNgtdURQ
8aQI5KInqKGEBkvwMh+XZNZ8Q7HmEXJ4od0WWCaOeXdAlfjHKAJ+P6mmTtyW9XAI
0sk7M3EWrBwzJh0lJe27Uji3Z04noVzR5V9IKo9OYVqpx1REROArLc/grN9VCZyb
STOs1RIQOkBpp0leOniXW+vOX9WZoCF0W5YEOITrkds6z8QcbxGgm4v5ixhbaeOC
KGsXpDfnKO667V6c9mBV0Quq/X3vsf81pWlrgDtaQjvxaOGKUs9IFhJ6gOIeNDln
0zD1QDGf9ULnFermTJmfby03aATmyRYvR891nqtm9jgO90V+9m2eIV31SpqRaenh
K2RDGfYCxDPxaaR7plktbOPpi5mGmthU+nAYE8yCIv1ZbyJoROA38LCgpRB1c13X
OvDZOcLSxceq28MwwskRZbJE8FKLF5ZVwrIYu1c+jtGpxmQlJ5ElUSoDCHqU9JjK
WCUhUtLTZliuhhgf5SJZ3DvwROCgdaOoZzdq9Ym3sjFMCYew20+FWAoQzVZ3BW62
Rx7J/+GDXpZ74Bfr5XKxOsKqWTjPm2cvxkCBwXFC1ZzMlBAaaD0L2RpQ8LoVpkDT
0C/VF5kjtP03J3Q1Fmv0p/dR51du9vpJdoeaH8t2OFknf7nnFNmd0dje9tRotOn4
qTUZ3QB+jvNl+qYLR7IIRR7BZluQGsJHypsVwSnazjbr+YWuALvA47hCYuN/mGHu
Nxuw+ngcGwG1jGFt1LJchFwMMYn2m/j4wnUC1RgU7AOnXdsJNZi/G3UDvdB3BNKa
kauWzcLSRFiSPnQsZM/1KNu5XO/PPqnuQAZINB+ehvtPG0vC+zp9jVps2NPfxPt/
iOnM3iz1qZDwsjVkSVdFcfZJH6Yrx2smG6s9QYiZxcTiGrAZGj28tc3Jtu7H5qnh
UhNp7iCnVEMvq2z2VqCwcl89OXAcP7QufVH41kQmDaz7XVofrJRz0ALB+9BC4M2u
XD6iwZ5kGH7K3xbajF3YtDyNwW0AXjEyrT8Zc9Q5DZua+PhPYAkKxi838RabZtYJ
lap7CwXCH6X+7LBHgwalBIIIzK7flVtwfglNPAWPs9ljnyxxVpzUfa3ynYG7UwZf
S2qoJ0ujU9TLkdf9PHXPyReScMjTa1GvFS423cyjpNSzJ/QGWXZmAsGTxJleF1gf
YhQT7L7PU1H4zRtui2yx2SUEEQXOIyu/XoRPlTmJj+A8DVXn+Xf49JMO/qBDHWrx
o+jx2Z1l7VsgDp02mUtUqYNmCyr8erH4BjTYLbkZqm/A85KrpdxYcyLkx3v/g/to
wxMUeCSlJKqWP96DV1dEMbCUIVn2sbV+wqG8cXaRsWuHvYgl0ffRqZH4q63s6pl0
gVdjy+EswVyLn6WwpWfOKs/dG0lOGcW5om5QtQRt4Vk=
`pragma protect end_protected
