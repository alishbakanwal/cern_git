-- gx_std_x5.vhd

-- Generated using ACDS version 16.0 211

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity gx_std_x5 is
	port (
		pll_powerdown           : in  std_logic_vector(0 downto 0)   := (others => '0'); --           pll_powerdown.pll_powerdown
		tx_analogreset          : in  std_logic_vector(4 downto 0)   := (others => '0'); --          tx_analogreset.tx_analogreset
		tx_digitalreset         : in  std_logic_vector(4 downto 0)   := (others => '0'); --         tx_digitalreset.tx_digitalreset
		tx_serial_data          : out std_logic_vector(4 downto 0);                      --          tx_serial_data.tx_serial_data
		ext_pll_clk             : in  std_logic_vector(4 downto 0)   := (others => '0'); --             ext_pll_clk.ext_pll_clk
		rx_analogreset          : in  std_logic_vector(4 downto 0)   := (others => '0'); --          rx_analogreset.rx_analogreset
		rx_digitalreset         : in  std_logic_vector(4 downto 0)   := (others => '0'); --         rx_digitalreset.rx_digitalreset
		rx_cdr_refclk           : in  std_logic_vector(0 downto 0)   := (others => '0'); --           rx_cdr_refclk.rx_cdr_refclk
		rx_serial_data          : in  std_logic_vector(4 downto 0)   := (others => '0'); --          rx_serial_data.rx_serial_data
		rx_is_lockedtoref       : out std_logic_vector(4 downto 0);                      --       rx_is_lockedtoref.rx_is_lockedtoref
		rx_is_lockedtodata      : out std_logic_vector(4 downto 0);                      --      rx_is_lockedtodata.rx_is_lockedtodata
		rx_seriallpbken         : in  std_logic_vector(4 downto 0)   := (others => '0'); --         rx_seriallpbken.rx_seriallpbken
		tx_std_coreclkin        : in  std_logic_vector(4 downto 0)   := (others => '0'); --        tx_std_coreclkin.tx_std_coreclkin
		rx_std_coreclkin        : in  std_logic_vector(4 downto 0)   := (others => '0'); --        rx_std_coreclkin.rx_std_coreclkin
		tx_std_clkout           : out std_logic_vector(4 downto 0);                      --           tx_std_clkout.tx_std_clkout
		rx_std_clkout           : out std_logic_vector(4 downto 0);                      --           rx_std_clkout.rx_std_clkout
		tx_std_polinv           : in  std_logic_vector(4 downto 0)   := (others => '0'); --           tx_std_polinv.tx_std_polinv
		rx_std_polinv           : in  std_logic_vector(4 downto 0)   := (others => '0'); --           rx_std_polinv.rx_std_polinv
		tx_cal_busy             : out std_logic_vector(4 downto 0);                      --             tx_cal_busy.tx_cal_busy
		rx_cal_busy             : out std_logic_vector(4 downto 0);                      --             rx_cal_busy.rx_cal_busy
		reconfig_to_xcvr        : in  std_logic_vector(349 downto 0) := (others => '0'); --        reconfig_to_xcvr.reconfig_to_xcvr
		reconfig_from_xcvr      : out std_logic_vector(229 downto 0);                    --      reconfig_from_xcvr.reconfig_from_xcvr
		tx_parallel_data        : in  std_logic_vector(199 downto 0) := (others => '0'); --        tx_parallel_data.tx_parallel_data
		unused_tx_parallel_data : in  std_logic_vector(119 downto 0) := (others => '0'); -- unused_tx_parallel_data.unused_tx_parallel_data
		rx_parallel_data        : out std_logic_vector(199 downto 0);                    --        rx_parallel_data.rx_parallel_data
		unused_rx_parallel_data : out std_logic_vector(119 downto 0)                     -- unused_rx_parallel_data.unused_rx_parallel_data
	);
end entity gx_std_x5;

architecture rtl of gx_std_x5 is
	component altera_xcvr_native_sv is
		generic (
			tx_enable                       : integer := 1;
			rx_enable                       : integer := 1;
			enable_std                      : integer := 0;
			enable_teng                     : integer := 0;
			data_path_select                : string  := "pma_direct";
			channels                        : integer := 1;
			bonded_mode                     : string  := "non_bonded";
			data_rate                       : string  := "";
			pma_width                       : integer := 80;
			tx_pma_clk_div                  : integer := 1;
			tx_pma_txdetectrx_ctrl          : integer := 0;
			pll_reconfig_enable             : integer := 0;
			pll_external_enable             : integer := 0;
			pll_data_rate                   : string  := "0 Mbps";
			pll_type                        : string  := "CMU";
			pll_network_select              : string  := "x1";
			plls                            : integer := 1;
			pll_select                      : integer := 0;
			pll_refclk_cnt                  : integer := 1;
			pll_refclk_select               : string  := "0";
			pll_refclk_freq                 : string  := "125.0 MHz";
			pll_feedback_path               : string  := "internal";
			cdr_reconfig_enable             : integer := 0;
			cdr_refclk_cnt                  : integer := 1;
			cdr_refclk_select               : integer := 0;
			cdr_refclk_freq                 : string  := "";
			rx_ppm_detect_threshold         : string  := "1000";
			rx_clkslip_enable               : integer := 0;
			std_protocol_hint               : string  := "basic";
			std_pcs_pma_width               : integer := 10;
			std_low_latency_bypass_enable   : integer := 0;
			std_tx_pcfifo_mode              : string  := "low_latency";
			std_rx_pcfifo_mode              : string  := "low_latency";
			std_rx_byte_order_enable        : integer := 0;
			std_rx_byte_order_mode          : string  := "manual";
			std_rx_byte_order_width         : integer := 10;
			std_rx_byte_order_symbol_count  : integer := 1;
			std_rx_byte_order_pattern       : string  := "0";
			std_rx_byte_order_pad           : string  := "0";
			std_tx_byte_ser_enable          : integer := 0;
			std_rx_byte_deser_enable        : integer := 0;
			std_tx_8b10b_enable             : integer := 0;
			std_tx_8b10b_disp_ctrl_enable   : integer := 0;
			std_rx_8b10b_enable             : integer := 0;
			std_rx_rmfifo_enable            : integer := 0;
			std_rx_rmfifo_pattern_p         : string  := "00000";
			std_rx_rmfifo_pattern_n         : string  := "00000";
			std_tx_bitslip_enable           : integer := 0;
			std_rx_word_aligner_mode        : string  := "bit_slip";
			std_rx_word_aligner_pattern_len : integer := 7;
			std_rx_word_aligner_pattern     : string  := "0000000000";
			std_rx_word_aligner_rknumber    : integer := 3;
			std_rx_word_aligner_renumber    : integer := 3;
			std_rx_word_aligner_rgnumber    : integer := 3;
			std_rx_run_length_val           : integer := 31;
			std_tx_bitrev_enable            : integer := 0;
			std_rx_bitrev_enable            : integer := 0;
			std_tx_byterev_enable           : integer := 0;
			std_rx_byterev_enable           : integer := 0;
			std_tx_polinv_enable            : integer := 0;
			std_rx_polinv_enable            : integer := 0;
			teng_protocol_hint              : string  := "basic";
			teng_pcs_pma_width              : integer := 40;
			teng_pld_pcs_width              : integer := 40;
			teng_txfifo_mode                : string  := "phase_comp";
			teng_txfifo_full                : integer := 31;
			teng_txfifo_empty               : integer := 0;
			teng_txfifo_pfull               : integer := 23;
			teng_txfifo_pempty              : integer := 2;
			teng_rxfifo_mode                : string  := "phase_comp";
			teng_rxfifo_full                : integer := 31;
			teng_rxfifo_empty               : integer := 0;
			teng_rxfifo_pfull               : integer := 23;
			teng_rxfifo_pempty              : integer := 2;
			teng_rxfifo_align_del           : integer := 0;
			teng_rxfifo_control_del         : integer := 0;
			teng_tx_frmgen_enable           : integer := 0;
			teng_tx_frmgen_user_length      : integer := 2048;
			teng_tx_frmgen_burst_enable     : integer := 0;
			teng_rx_frmsync_enable          : integer := 0;
			teng_rx_frmsync_user_length     : integer := 2048;
			teng_frmgensync_diag_word       : string  := "6400000000000000";
			teng_frmgensync_scrm_word       : string  := "2800000000000000";
			teng_frmgensync_skip_word       : string  := "1e1e1e1e1e1e1e1e";
			teng_frmgensync_sync_word       : string  := "78f678f678f678f6";
			teng_tx_sh_err                  : integer := 0;
			teng_tx_crcgen_enable           : integer := 0;
			teng_rx_crcchk_enable           : integer := 0;
			teng_tx_64b66b_enable           : integer := 0;
			teng_rx_64b66b_enable           : integer := 0;
			teng_tx_scram_enable            : integer := 0;
			teng_tx_scram_user_seed         : string  := "000000000000000";
			teng_rx_descram_enable          : integer := 0;
			teng_tx_dispgen_enable          : integer := 0;
			teng_rx_dispchk_enable          : integer := 0;
			teng_rx_blksync_enable          : integer := 0;
			teng_tx_polinv_enable           : integer := 0;
			teng_tx_bitslip_enable          : integer := 0;
			teng_rx_polinv_enable           : integer := 0;
			teng_rx_bitslip_enable          : integer := 0
		);
		port (
			pll_powerdown             : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- pll_powerdown
			tx_analogreset            : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- tx_analogreset
			tx_digitalreset           : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- tx_digitalreset
			tx_serial_data            : out std_logic_vector(4 downto 0);                      -- tx_serial_data
			ext_pll_clk               : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- ext_pll_clk
			rx_analogreset            : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_analogreset
			rx_digitalreset           : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_digitalreset
			rx_cdr_refclk             : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- rx_cdr_refclk
			rx_serial_data            : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_serial_data
			rx_is_lockedtoref         : out std_logic_vector(4 downto 0);                      -- rx_is_lockedtoref
			rx_is_lockedtodata        : out std_logic_vector(4 downto 0);                      -- rx_is_lockedtodata
			rx_seriallpbken           : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_seriallpbken
			tx_std_coreclkin          : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- tx_std_coreclkin
			rx_std_coreclkin          : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_std_coreclkin
			tx_std_clkout             : out std_logic_vector(4 downto 0);                      -- tx_std_clkout
			rx_std_clkout             : out std_logic_vector(4 downto 0);                      -- rx_std_clkout
			tx_std_polinv             : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- tx_std_polinv
			rx_std_polinv             : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_std_polinv
			tx_cal_busy               : out std_logic_vector(4 downto 0);                      -- tx_cal_busy
			rx_cal_busy               : out std_logic_vector(4 downto 0);                      -- rx_cal_busy
			reconfig_to_xcvr          : in  std_logic_vector(349 downto 0) := (others => 'X'); -- reconfig_to_xcvr
			reconfig_from_xcvr        : out std_logic_vector(229 downto 0);                    -- reconfig_from_xcvr
			tx_parallel_data          : in  std_logic_vector(319 downto 0) := (others => 'X'); -- unused_tx_parallel_data
			rx_parallel_data          : out std_logic_vector(319 downto 0);                    -- unused_rx_parallel_data
			tx_pll_refclk             : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- tx_pll_refclk
			tx_pma_clkout             : out std_logic_vector(4 downto 0);                      -- tx_pma_clkout
			tx_pma_pclk               : out std_logic_vector(4 downto 0);                      -- tx_pma_pclk
			tx_pma_parallel_data      : in  std_logic_vector(399 downto 0) := (others => 'X'); -- tx_pma_parallel_data
			pll_locked                : out std_logic_vector(0 downto 0);                      -- pll_locked
			rx_pma_clkout             : out std_logic_vector(4 downto 0);                      -- rx_pma_clkout
			rx_pma_pclk               : out std_logic_vector(4 downto 0);                      -- rx_pma_pclk
			rx_pma_parallel_data      : out std_logic_vector(399 downto 0);                    -- rx_pma_parallel_data
			rx_clkslip                : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_clkslip
			rx_clklow                 : out std_logic_vector(4 downto 0);                      -- rx_clklow
			rx_fref                   : out std_logic_vector(4 downto 0);                      -- rx_fref
			rx_set_locktodata         : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_set_locktodata
			rx_set_locktoref          : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_set_locktoref
			rx_signaldetect           : out std_logic_vector(4 downto 0);                      -- rx_signaldetect
			rx_pma_qpipulldn          : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_pma_qpipulldn
			tx_pma_qpipullup          : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- tx_pma_qpipullup
			tx_pma_qpipulldn          : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- tx_pma_qpipulldn
			tx_pma_txdetectrx         : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- tx_pma_txdetectrx
			tx_pma_rxfound            : out std_logic_vector(4 downto 0);                      -- tx_pma_rxfound
			rx_std_prbs_done          : out std_logic_vector(4 downto 0);                      -- rx_std_prbs_done
			rx_std_prbs_err           : out std_logic_vector(4 downto 0);                      -- rx_std_prbs_err
			tx_std_pcfifo_full        : out std_logic_vector(4 downto 0);                      -- tx_std_pcfifo_full
			tx_std_pcfifo_empty       : out std_logic_vector(4 downto 0);                      -- tx_std_pcfifo_empty
			rx_std_pcfifo_full        : out std_logic_vector(4 downto 0);                      -- rx_std_pcfifo_full
			rx_std_pcfifo_empty       : out std_logic_vector(4 downto 0);                      -- rx_std_pcfifo_empty
			rx_std_byteorder_ena      : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_std_byteorder_ena
			rx_std_byteorder_flag     : out std_logic_vector(4 downto 0);                      -- rx_std_byteorder_flag
			rx_std_rmfifo_full        : out std_logic_vector(4 downto 0);                      -- rx_std_rmfifo_full
			rx_std_rmfifo_empty       : out std_logic_vector(4 downto 0);                      -- rx_std_rmfifo_empty
			rx_std_wa_patternalign    : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_std_wa_patternalign
			rx_std_wa_a1a2size        : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_std_wa_a1a2size
			tx_std_bitslipboundarysel : in  std_logic_vector(24 downto 0)  := (others => 'X'); -- tx_std_bitslipboundarysel
			rx_std_bitslipboundarysel : out std_logic_vector(24 downto 0);                     -- rx_std_bitslipboundarysel
			rx_std_bitslip            : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_std_bitslip
			rx_std_runlength_err      : out std_logic_vector(4 downto 0);                      -- rx_std_runlength_err
			rx_std_bitrev_ena         : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_std_bitrev_ena
			rx_std_byterev_ena        : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_std_byterev_ena
			tx_std_elecidle           : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- tx_std_elecidle
			rx_std_signaldetect       : out std_logic_vector(4 downto 0);                      -- rx_std_signaldetect
			tx_10g_coreclkin          : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- tx_10g_coreclkin
			rx_10g_coreclkin          : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_10g_coreclkin
			tx_10g_clkout             : out std_logic_vector(4 downto 0);                      -- tx_10g_clkout
			rx_10g_clkout             : out std_logic_vector(4 downto 0);                      -- rx_10g_clkout
			rx_10g_clk33out           : out std_logic_vector(4 downto 0);                      -- rx_10g_clk33out
			rx_10g_prbs_err_clr       : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_10g_prbs_err_clr
			rx_10g_prbs_done          : out std_logic_vector(4 downto 0);                      -- rx_10g_prbs_done
			rx_10g_prbs_err           : out std_logic_vector(4 downto 0);                      -- rx_10g_prbs_err
			tx_10g_control            : in  std_logic_vector(44 downto 0)  := (others => 'X'); -- tx_10g_control
			rx_10g_control            : out std_logic_vector(49 downto 0);                     -- rx_10g_control
			tx_10g_data_valid         : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- tx_10g_data_valid
			tx_10g_fifo_full          : out std_logic_vector(4 downto 0);                      -- tx_10g_fifo_full
			tx_10g_fifo_pfull         : out std_logic_vector(4 downto 0);                      -- tx_10g_fifo_pfull
			tx_10g_fifo_empty         : out std_logic_vector(4 downto 0);                      -- tx_10g_fifo_empty
			tx_10g_fifo_pempty        : out std_logic_vector(4 downto 0);                      -- tx_10g_fifo_pempty
			tx_10g_fifo_del           : out std_logic_vector(4 downto 0);                      -- tx_10g_fifo_del
			tx_10g_fifo_insert        : out std_logic_vector(4 downto 0);                      -- tx_10g_fifo_insert
			rx_10g_fifo_rd_en         : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_10g_fifo_rd_en
			rx_10g_data_valid         : out std_logic_vector(4 downto 0);                      -- rx_10g_data_valid
			rx_10g_fifo_full          : out std_logic_vector(4 downto 0);                      -- rx_10g_fifo_full
			rx_10g_fifo_pfull         : out std_logic_vector(4 downto 0);                      -- rx_10g_fifo_pfull
			rx_10g_fifo_empty         : out std_logic_vector(4 downto 0);                      -- rx_10g_fifo_empty
			rx_10g_fifo_pempty        : out std_logic_vector(4 downto 0);                      -- rx_10g_fifo_pempty
			rx_10g_fifo_del           : out std_logic_vector(4 downto 0);                      -- rx_10g_fifo_del
			rx_10g_fifo_insert        : out std_logic_vector(4 downto 0);                      -- rx_10g_fifo_insert
			rx_10g_fifo_align_val     : out std_logic_vector(4 downto 0);                      -- rx_10g_fifo_align_val
			rx_10g_fifo_align_clr     : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_10g_fifo_align_clr
			rx_10g_fifo_align_en      : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_10g_fifo_align_en
			tx_10g_frame              : out std_logic_vector(4 downto 0);                      -- tx_10g_frame
			tx_10g_frame_diag_status  : in  std_logic_vector(9 downto 0)   := (others => 'X'); -- tx_10g_frame_diag_status
			tx_10g_frame_burst_en     : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- tx_10g_frame_burst_en
			rx_10g_frame              : out std_logic_vector(4 downto 0);                      -- rx_10g_frame
			rx_10g_frame_lock         : out std_logic_vector(4 downto 0);                      -- rx_10g_frame_lock
			rx_10g_frame_mfrm_err     : out std_logic_vector(4 downto 0);                      -- rx_10g_frame_mfrm_err
			rx_10g_frame_sync_err     : out std_logic_vector(4 downto 0);                      -- rx_10g_frame_sync_err
			rx_10g_frame_skip_ins     : out std_logic_vector(4 downto 0);                      -- rx_10g_frame_skip_ins
			rx_10g_frame_pyld_ins     : out std_logic_vector(4 downto 0);                      -- rx_10g_frame_pyld_ins
			rx_10g_frame_skip_err     : out std_logic_vector(4 downto 0);                      -- rx_10g_frame_skip_err
			rx_10g_frame_diag_err     : out std_logic_vector(4 downto 0);                      -- rx_10g_frame_diag_err
			rx_10g_frame_diag_status  : out std_logic_vector(9 downto 0);                      -- rx_10g_frame_diag_status
			rx_10g_crc32_err          : out std_logic_vector(4 downto 0);                      -- rx_10g_crc32err
			rx_10g_descram_err        : out std_logic_vector(4 downto 0);                      -- rx_10g_descram_err
			rx_10g_blk_lock           : out std_logic_vector(4 downto 0);                      -- rx_10g_blk_lock
			rx_10g_blk_sh_err         : out std_logic_vector(4 downto 0);                      -- rx_10g_blk_sh_err
			tx_10g_bitslip            : in  std_logic_vector(34 downto 0)  := (others => 'X'); -- tx_10g_bitslip
			rx_10g_bitslip            : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_10g_bitslip
			rx_10g_highber            : out std_logic_vector(4 downto 0);                      -- rx_10g_highber
			rx_10g_highber_clr_cnt    : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- rx_10g_highber_clr_cnt
			rx_10g_clr_errblk_count   : in  std_logic_vector(4 downto 0)   := (others => 'X')  -- rx_10g_clr_errblk_count
		);
	end component altera_xcvr_native_sv;

	signal gx_std_x5_inst_rx_parallel_data : std_logic_vector(319 downto 0); -- port fragment

begin

	gx_std_x5_inst : component altera_xcvr_native_sv
		generic map (
			tx_enable                       => 1,
			rx_enable                       => 1,
			enable_std                      => 1,
			enable_teng                     => 0,
			data_path_select                => "standard",
			channels                        => 5,
			bonded_mode                     => "xN",
			data_rate                       => "4800 Mbps",
			pma_width                       => 20,
			tx_pma_clk_div                  => 1,
			tx_pma_txdetectrx_ctrl          => 0,
			pll_reconfig_enable             => 0,
			pll_external_enable             => 1,
			pll_data_rate                   => "4800 Mbps",
			pll_type                        => "CMU",
			pll_network_select              => "x1",
			plls                            => 1,
			pll_select                      => 0,
			pll_refclk_cnt                  => 1,
			pll_refclk_select               => "0",
			pll_refclk_freq                 => "125.0 MHz",
			pll_feedback_path               => "internal",
			cdr_reconfig_enable             => 0,
			cdr_refclk_cnt                  => 1,
			cdr_refclk_select               => 0,
			cdr_refclk_freq                 => "120.0 MHz",
			rx_ppm_detect_threshold         => "1000",
			rx_clkslip_enable               => 0,
			std_protocol_hint               => "basic",
			std_pcs_pma_width               => 20,
			std_low_latency_bypass_enable   => 0,
			std_tx_pcfifo_mode              => "low_latency",
			std_rx_pcfifo_mode              => "low_latency",
			std_rx_byte_order_enable        => 0,
			std_rx_byte_order_mode          => "manual",
			std_rx_byte_order_width         => 10,
			std_rx_byte_order_symbol_count  => 1,
			std_rx_byte_order_pattern       => "0",
			std_rx_byte_order_pad           => "0",
			std_tx_byte_ser_enable          => 1,
			std_rx_byte_deser_enable        => 1,
			std_tx_8b10b_enable             => 0,
			std_tx_8b10b_disp_ctrl_enable   => 0,
			std_rx_8b10b_enable             => 0,
			std_rx_rmfifo_enable            => 0,
			std_rx_rmfifo_pattern_p         => "00000",
			std_rx_rmfifo_pattern_n         => "00000",
			std_tx_bitslip_enable           => 0,
			std_rx_word_aligner_mode        => "bit_slip",
			std_rx_word_aligner_pattern_len => 7,
			std_rx_word_aligner_pattern     => "0000000000",
			std_rx_word_aligner_rknumber    => 3,
			std_rx_word_aligner_renumber    => 3,
			std_rx_word_aligner_rgnumber    => 3,
			std_rx_run_length_val           => 31,
			std_tx_bitrev_enable            => 0,
			std_rx_bitrev_enable            => 0,
			std_tx_byterev_enable           => 0,
			std_rx_byterev_enable           => 0,
			std_tx_polinv_enable            => 1,
			std_rx_polinv_enable            => 1,
			teng_protocol_hint              => "basic",
			teng_pcs_pma_width              => 40,
			teng_pld_pcs_width              => 40,
			teng_txfifo_mode                => "phase_comp",
			teng_txfifo_full                => 31,
			teng_txfifo_empty               => 0,
			teng_txfifo_pfull               => 23,
			teng_txfifo_pempty              => 2,
			teng_rxfifo_mode                => "phase_comp",
			teng_rxfifo_full                => 31,
			teng_rxfifo_empty               => 0,
			teng_rxfifo_pfull               => 23,
			teng_rxfifo_pempty              => 2,
			teng_rxfifo_align_del           => 0,
			teng_rxfifo_control_del         => 0,
			teng_tx_frmgen_enable           => 0,
			teng_tx_frmgen_user_length      => 2048,
			teng_tx_frmgen_burst_enable     => 0,
			teng_rx_frmsync_enable          => 0,
			teng_rx_frmsync_user_length     => 2048,
			teng_frmgensync_diag_word       => "6400000000000000",
			teng_frmgensync_scrm_word       => "2800000000000000",
			teng_frmgensync_skip_word       => "1e1e1e1e1e1e1e1e",
			teng_frmgensync_sync_word       => "78f678f678f678f6",
			teng_tx_sh_err                  => 0,
			teng_tx_crcgen_enable           => 0,
			teng_rx_crcchk_enable           => 0,
			teng_tx_64b66b_enable           => 0,
			teng_rx_64b66b_enable           => 0,
			teng_tx_scram_enable            => 0,
			teng_tx_scram_user_seed         => "000000000000000",
			teng_rx_descram_enable          => 0,
			teng_tx_dispgen_enable          => 0,
			teng_rx_dispchk_enable          => 0,
			teng_rx_blksync_enable          => 0,
			teng_tx_polinv_enable           => 0,
			teng_tx_bitslip_enable          => 0,
			teng_rx_polinv_enable           => 0,
			teng_rx_bitslip_enable          => 0
		)
		port map (
			pll_powerdown             => pll_powerdown,                                                                                                                                                                                                                                                                                                                                                                                                      --      pll_powerdown.pll_powerdown
			tx_analogreset            => tx_analogreset,                                                                                                                                                                                                                                                                                                                                                                                                     --     tx_analogreset.tx_analogreset
			tx_digitalreset           => tx_digitalreset,                                                                                                                                                                                                                                                                                                                                                                                                    --    tx_digitalreset.tx_digitalreset
			tx_serial_data            => tx_serial_data,                                                                                                                                                                                                                                                                                                                                                                                                     --     tx_serial_data.tx_serial_data
			ext_pll_clk               => ext_pll_clk,                                                                                                                                                                                                                                                                                                                                                                                                        --        ext_pll_clk.ext_pll_clk
			rx_analogreset            => rx_analogreset,                                                                                                                                                                                                                                                                                                                                                                                                     --     rx_analogreset.rx_analogreset
			rx_digitalreset           => rx_digitalreset,                                                                                                                                                                                                                                                                                                                                                                                                    --    rx_digitalreset.rx_digitalreset
			rx_cdr_refclk             => rx_cdr_refclk,                                                                                                                                                                                                                                                                                                                                                                                                      --      rx_cdr_refclk.rx_cdr_refclk
			rx_serial_data            => rx_serial_data,                                                                                                                                                                                                                                                                                                                                                                                                     --     rx_serial_data.rx_serial_data
			rx_is_lockedtoref         => rx_is_lockedtoref,                                                                                                                                                                                                                                                                                                                                                                                                  --  rx_is_lockedtoref.rx_is_lockedtoref
			rx_is_lockedtodata        => rx_is_lockedtodata,                                                                                                                                                                                                                                                                                                                                                                                                 -- rx_is_lockedtodata.rx_is_lockedtodata
			rx_seriallpbken           => rx_seriallpbken,                                                                                                                                                                                                                                                                                                                                                                                                    --    rx_seriallpbken.rx_seriallpbken
			tx_std_coreclkin          => tx_std_coreclkin,                                                                                                                                                                                                                                                                                                                                                                                                   --   tx_std_coreclkin.tx_std_coreclkin
			rx_std_coreclkin          => rx_std_coreclkin,                                                                                                                                                                                                                                                                                                                                                                                                   --   rx_std_coreclkin.rx_std_coreclkin
			tx_std_clkout             => tx_std_clkout,                                                                                                                                                                                                                                                                                                                                                                                                      --      tx_std_clkout.tx_std_clkout
			rx_std_clkout             => rx_std_clkout,                                                                                                                                                                                                                                                                                                                                                                                                      --      rx_std_clkout.rx_std_clkout
			tx_std_polinv             => tx_std_polinv,                                                                                                                                                                                                                                                                                                                                                                                                      --      tx_std_polinv.tx_std_polinv
			rx_std_polinv             => rx_std_polinv,                                                                                                                                                                                                                                                                                                                                                                                                      --      rx_std_polinv.rx_std_polinv
			tx_cal_busy               => tx_cal_busy,                                                                                                                                                                                                                                                                                                                                                                                                        --        tx_cal_busy.tx_cal_busy
			rx_cal_busy               => rx_cal_busy,                                                                                                                                                                                                                                                                                                                                                                                                        --        rx_cal_busy.rx_cal_busy
			reconfig_to_xcvr          => reconfig_to_xcvr,                                                                                                                                                                                                                                                                                                                                                                                                   --   reconfig_to_xcvr.reconfig_to_xcvr
			reconfig_from_xcvr        => reconfig_from_xcvr,                                                                                                                                                                                                                                                                                                                                                                                                 -- reconfig_from_xcvr.reconfig_from_xcvr
			tx_parallel_data(0)       => tx_parallel_data(0),                                                                                                                                                                                                                                                                                                                                                                                                --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(1)       => tx_parallel_data(1),                                                                                                                                                                                                                                                                                                                                                                                                --                   .tx_parallel_data
			tx_parallel_data(2)       => tx_parallel_data(2),                                                                                                                                                                                                                                                                                                                                                                                                --                   .tx_parallel_data
			tx_parallel_data(3)       => tx_parallel_data(3),                                                                                                                                                                                                                                                                                                                                                                                                --                   .tx_parallel_data
			tx_parallel_data(4)       => tx_parallel_data(4),                                                                                                                                                                                                                                                                                                                                                                                                --                   .tx_parallel_data
			tx_parallel_data(5)       => tx_parallel_data(5),                                                                                                                                                                                                                                                                                                                                                                                                --                   .tx_parallel_data
			tx_parallel_data(6)       => tx_parallel_data(6),                                                                                                                                                                                                                                                                                                                                                                                                --                   .tx_parallel_data
			tx_parallel_data(7)       => tx_parallel_data(7),                                                                                                                                                                                                                                                                                                                                                                                                --                   .tx_parallel_data
			tx_parallel_data(8)       => tx_parallel_data(8),                                                                                                                                                                                                                                                                                                                                                                                                --                   .tx_parallel_data
			tx_parallel_data(9)       => tx_parallel_data(9),                                                                                                                                                                                                                                                                                                                                                                                                --                   .tx_parallel_data
			tx_parallel_data(10)      => unused_tx_parallel_data(0),                                                                                                                                                                                                                                                                                                                                                                                         --                   .tx_parallel_data
			tx_parallel_data(11)      => tx_parallel_data(10),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(12)      => tx_parallel_data(11),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(13)      => tx_parallel_data(12),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(14)      => tx_parallel_data(13),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(15)      => tx_parallel_data(14),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(16)      => tx_parallel_data(15),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(17)      => tx_parallel_data(16),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(18)      => tx_parallel_data(17),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(19)      => tx_parallel_data(18),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(20)      => tx_parallel_data(19),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(21)      => unused_tx_parallel_data(1),                                                                                                                                                                                                                                                                                                                                                                                         --                   .tx_parallel_data
			tx_parallel_data(22)      => tx_parallel_data(20),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(23)      => tx_parallel_data(21),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(24)      => tx_parallel_data(22),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(25)      => tx_parallel_data(23),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(26)      => tx_parallel_data(24),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(27)      => tx_parallel_data(25),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(28)      => tx_parallel_data(26),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(29)      => tx_parallel_data(27),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(30)      => tx_parallel_data(28),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(31)      => tx_parallel_data(29),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(32)      => unused_tx_parallel_data(2),                                                                                                                                                                                                                                                                                                                                                                                         --                   .tx_parallel_data
			tx_parallel_data(33)      => tx_parallel_data(30),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(34)      => tx_parallel_data(31),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(35)      => tx_parallel_data(32),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(36)      => tx_parallel_data(33),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(37)      => tx_parallel_data(34),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(38)      => tx_parallel_data(35),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(39)      => tx_parallel_data(36),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(40)      => tx_parallel_data(37),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(41)      => tx_parallel_data(38),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(42)      => tx_parallel_data(39),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(43)      => unused_tx_parallel_data(3),                                                                                                                                                                                                                                                                                                                                                                                         --                   .tx_parallel_data
			tx_parallel_data(44)      => unused_tx_parallel_data(4),                                                                                                                                                                                                                                                                                                                                                                                         --                   .tx_parallel_data
			tx_parallel_data(45)      => unused_tx_parallel_data(5),                                                                                                                                                                                                                                                                                                                                                                                         --                   .tx_parallel_data
			tx_parallel_data(46)      => unused_tx_parallel_data(6),                                                                                                                                                                                                                                                                                                                                                                                         --                   .tx_parallel_data
			tx_parallel_data(47)      => unused_tx_parallel_data(7),                                                                                                                                                                                                                                                                                                                                                                                         --                   .tx_parallel_data
			tx_parallel_data(48)      => unused_tx_parallel_data(8),                                                                                                                                                                                                                                                                                                                                                                                         --                   .tx_parallel_data
			tx_parallel_data(49)      => unused_tx_parallel_data(9),                                                                                                                                                                                                                                                                                                                                                                                         --                   .tx_parallel_data
			tx_parallel_data(50)      => unused_tx_parallel_data(10),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(51)      => unused_tx_parallel_data(11),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(52)      => unused_tx_parallel_data(12),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(53)      => unused_tx_parallel_data(13),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(54)      => unused_tx_parallel_data(14),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(55)      => unused_tx_parallel_data(15),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(56)      => unused_tx_parallel_data(16),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(57)      => unused_tx_parallel_data(17),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(58)      => unused_tx_parallel_data(18),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(59)      => unused_tx_parallel_data(19),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(60)      => unused_tx_parallel_data(20),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(61)      => unused_tx_parallel_data(21),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(62)      => unused_tx_parallel_data(22),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(63)      => unused_tx_parallel_data(23),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(64)      => tx_parallel_data(40),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(65)      => tx_parallel_data(41),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(66)      => tx_parallel_data(42),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(67)      => tx_parallel_data(43),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(68)      => tx_parallel_data(44),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(69)      => tx_parallel_data(45),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(70)      => tx_parallel_data(46),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(71)      => tx_parallel_data(47),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(72)      => tx_parallel_data(48),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(73)      => tx_parallel_data(49),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(74)      => unused_tx_parallel_data(24),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(75)      => tx_parallel_data(50),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(76)      => tx_parallel_data(51),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(77)      => tx_parallel_data(52),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(78)      => tx_parallel_data(53),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(79)      => tx_parallel_data(54),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(80)      => tx_parallel_data(55),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(81)      => tx_parallel_data(56),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(82)      => tx_parallel_data(57),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(83)      => tx_parallel_data(58),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(84)      => tx_parallel_data(59),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(85)      => unused_tx_parallel_data(25),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(86)      => tx_parallel_data(60),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(87)      => tx_parallel_data(61),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(88)      => tx_parallel_data(62),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(89)      => tx_parallel_data(63),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(90)      => tx_parallel_data(64),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(91)      => tx_parallel_data(65),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(92)      => tx_parallel_data(66),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(93)      => tx_parallel_data(67),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(94)      => tx_parallel_data(68),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(95)      => tx_parallel_data(69),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(96)      => unused_tx_parallel_data(26),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(97)      => tx_parallel_data(70),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(98)      => tx_parallel_data(71),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(99)      => tx_parallel_data(72),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(100)     => tx_parallel_data(73),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(101)     => tx_parallel_data(74),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(102)     => tx_parallel_data(75),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(103)     => tx_parallel_data(76),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(104)     => tx_parallel_data(77),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(105)     => tx_parallel_data(78),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(106)     => tx_parallel_data(79),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(107)     => unused_tx_parallel_data(27),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(108)     => unused_tx_parallel_data(28),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(109)     => unused_tx_parallel_data(29),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(110)     => unused_tx_parallel_data(30),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(111)     => unused_tx_parallel_data(31),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(112)     => unused_tx_parallel_data(32),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(113)     => unused_tx_parallel_data(33),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(114)     => unused_tx_parallel_data(34),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(115)     => unused_tx_parallel_data(35),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(116)     => unused_tx_parallel_data(36),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(117)     => unused_tx_parallel_data(37),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(118)     => unused_tx_parallel_data(38),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(119)     => unused_tx_parallel_data(39),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(120)     => unused_tx_parallel_data(40),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(121)     => unused_tx_parallel_data(41),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(122)     => unused_tx_parallel_data(42),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(123)     => unused_tx_parallel_data(43),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(124)     => unused_tx_parallel_data(44),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(125)     => unused_tx_parallel_data(45),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(126)     => unused_tx_parallel_data(46),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(127)     => unused_tx_parallel_data(47),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(128)     => tx_parallel_data(80),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(129)     => tx_parallel_data(81),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(130)     => tx_parallel_data(82),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(131)     => tx_parallel_data(83),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(132)     => tx_parallel_data(84),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(133)     => tx_parallel_data(85),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(134)     => tx_parallel_data(86),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(135)     => tx_parallel_data(87),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(136)     => tx_parallel_data(88),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(137)     => tx_parallel_data(89),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(138)     => unused_tx_parallel_data(48),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(139)     => tx_parallel_data(90),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(140)     => tx_parallel_data(91),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(141)     => tx_parallel_data(92),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(142)     => tx_parallel_data(93),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(143)     => tx_parallel_data(94),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(144)     => tx_parallel_data(95),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(145)     => tx_parallel_data(96),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(146)     => tx_parallel_data(97),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(147)     => tx_parallel_data(98),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(148)     => tx_parallel_data(99),                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(149)     => unused_tx_parallel_data(49),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(150)     => tx_parallel_data(100),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(151)     => tx_parallel_data(101),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(152)     => tx_parallel_data(102),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(153)     => tx_parallel_data(103),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(154)     => tx_parallel_data(104),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(155)     => tx_parallel_data(105),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(156)     => tx_parallel_data(106),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(157)     => tx_parallel_data(107),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(158)     => tx_parallel_data(108),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(159)     => tx_parallel_data(109),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(160)     => unused_tx_parallel_data(50),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(161)     => tx_parallel_data(110),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(162)     => tx_parallel_data(111),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(163)     => tx_parallel_data(112),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(164)     => tx_parallel_data(113),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(165)     => tx_parallel_data(114),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(166)     => tx_parallel_data(115),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(167)     => tx_parallel_data(116),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(168)     => tx_parallel_data(117),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(169)     => tx_parallel_data(118),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(170)     => tx_parallel_data(119),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(171)     => unused_tx_parallel_data(51),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(172)     => unused_tx_parallel_data(52),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(173)     => unused_tx_parallel_data(53),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(174)     => unused_tx_parallel_data(54),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(175)     => unused_tx_parallel_data(55),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(176)     => unused_tx_parallel_data(56),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(177)     => unused_tx_parallel_data(57),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(178)     => unused_tx_parallel_data(58),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(179)     => unused_tx_parallel_data(59),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(180)     => unused_tx_parallel_data(60),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(181)     => unused_tx_parallel_data(61),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(182)     => unused_tx_parallel_data(62),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(183)     => unused_tx_parallel_data(63),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(184)     => unused_tx_parallel_data(64),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(185)     => unused_tx_parallel_data(65),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(186)     => unused_tx_parallel_data(66),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(187)     => unused_tx_parallel_data(67),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(188)     => unused_tx_parallel_data(68),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(189)     => unused_tx_parallel_data(69),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(190)     => unused_tx_parallel_data(70),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(191)     => unused_tx_parallel_data(71),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(192)     => tx_parallel_data(120),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(193)     => tx_parallel_data(121),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(194)     => tx_parallel_data(122),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(195)     => tx_parallel_data(123),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(196)     => tx_parallel_data(124),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(197)     => tx_parallel_data(125),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(198)     => tx_parallel_data(126),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(199)     => tx_parallel_data(127),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(200)     => tx_parallel_data(128),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(201)     => tx_parallel_data(129),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(202)     => unused_tx_parallel_data(72),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(203)     => tx_parallel_data(130),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(204)     => tx_parallel_data(131),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(205)     => tx_parallel_data(132),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(206)     => tx_parallel_data(133),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(207)     => tx_parallel_data(134),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(208)     => tx_parallel_data(135),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(209)     => tx_parallel_data(136),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(210)     => tx_parallel_data(137),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(211)     => tx_parallel_data(138),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(212)     => tx_parallel_data(139),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(213)     => unused_tx_parallel_data(73),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(214)     => tx_parallel_data(140),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(215)     => tx_parallel_data(141),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(216)     => tx_parallel_data(142),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(217)     => tx_parallel_data(143),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(218)     => tx_parallel_data(144),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(219)     => tx_parallel_data(145),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(220)     => tx_parallel_data(146),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(221)     => tx_parallel_data(147),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(222)     => tx_parallel_data(148),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(223)     => tx_parallel_data(149),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(224)     => unused_tx_parallel_data(74),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(225)     => tx_parallel_data(150),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(226)     => tx_parallel_data(151),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(227)     => tx_parallel_data(152),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(228)     => tx_parallel_data(153),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(229)     => tx_parallel_data(154),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(230)     => tx_parallel_data(155),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(231)     => tx_parallel_data(156),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(232)     => tx_parallel_data(157),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(233)     => tx_parallel_data(158),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(234)     => tx_parallel_data(159),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(235)     => unused_tx_parallel_data(75),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(236)     => unused_tx_parallel_data(76),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(237)     => unused_tx_parallel_data(77),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(238)     => unused_tx_parallel_data(78),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(239)     => unused_tx_parallel_data(79),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(240)     => unused_tx_parallel_data(80),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(241)     => unused_tx_parallel_data(81),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(242)     => unused_tx_parallel_data(82),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(243)     => unused_tx_parallel_data(83),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(244)     => unused_tx_parallel_data(84),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(245)     => unused_tx_parallel_data(85),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(246)     => unused_tx_parallel_data(86),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(247)     => unused_tx_parallel_data(87),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(248)     => unused_tx_parallel_data(88),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(249)     => unused_tx_parallel_data(89),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(250)     => unused_tx_parallel_data(90),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(251)     => unused_tx_parallel_data(91),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(252)     => unused_tx_parallel_data(92),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(253)     => unused_tx_parallel_data(93),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(254)     => unused_tx_parallel_data(94),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(255)     => unused_tx_parallel_data(95),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(256)     => tx_parallel_data(160),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(257)     => tx_parallel_data(161),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(258)     => tx_parallel_data(162),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(259)     => tx_parallel_data(163),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(260)     => tx_parallel_data(164),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(261)     => tx_parallel_data(165),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(262)     => tx_parallel_data(166),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(263)     => tx_parallel_data(167),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(264)     => tx_parallel_data(168),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(265)     => tx_parallel_data(169),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(266)     => unused_tx_parallel_data(96),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(267)     => tx_parallel_data(170),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(268)     => tx_parallel_data(171),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(269)     => tx_parallel_data(172),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(270)     => tx_parallel_data(173),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(271)     => tx_parallel_data(174),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(272)     => tx_parallel_data(175),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(273)     => tx_parallel_data(176),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(274)     => tx_parallel_data(177),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(275)     => tx_parallel_data(178),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(276)     => tx_parallel_data(179),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(277)     => unused_tx_parallel_data(97),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(278)     => tx_parallel_data(180),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(279)     => tx_parallel_data(181),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(280)     => tx_parallel_data(182),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(281)     => tx_parallel_data(183),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(282)     => tx_parallel_data(184),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(283)     => tx_parallel_data(185),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(284)     => tx_parallel_data(186),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(285)     => tx_parallel_data(187),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(286)     => tx_parallel_data(188),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(287)     => tx_parallel_data(189),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(288)     => unused_tx_parallel_data(98),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(289)     => tx_parallel_data(190),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(290)     => tx_parallel_data(191),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(291)     => tx_parallel_data(192),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(292)     => tx_parallel_data(193),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(293)     => tx_parallel_data(194),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(294)     => tx_parallel_data(195),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(295)     => tx_parallel_data(196),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(296)     => tx_parallel_data(197),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(297)     => tx_parallel_data(198),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(298)     => tx_parallel_data(199),                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(299)     => unused_tx_parallel_data(99),                                                                                                                                                                                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(300)     => unused_tx_parallel_data(100),                                                                                                                                                                                                                                                                                                                                                                                       --                   .tx_parallel_data
			tx_parallel_data(301)     => unused_tx_parallel_data(101),                                                                                                                                                                                                                                                                                                                                                                                       --                   .tx_parallel_data
			tx_parallel_data(302)     => unused_tx_parallel_data(102),                                                                                                                                                                                                                                                                                                                                                                                       --                   .tx_parallel_data
			tx_parallel_data(303)     => unused_tx_parallel_data(103),                                                                                                                                                                                                                                                                                                                                                                                       --                   .tx_parallel_data
			tx_parallel_data(304)     => unused_tx_parallel_data(104),                                                                                                                                                                                                                                                                                                                                                                                       --                   .tx_parallel_data
			tx_parallel_data(305)     => unused_tx_parallel_data(105),                                                                                                                                                                                                                                                                                                                                                                                       --                   .tx_parallel_data
			tx_parallel_data(306)     => unused_tx_parallel_data(106),                                                                                                                                                                                                                                                                                                                                                                                       --                   .tx_parallel_data
			tx_parallel_data(307)     => unused_tx_parallel_data(107),                                                                                                                                                                                                                                                                                                                                                                                       --                   .tx_parallel_data
			tx_parallel_data(308)     => unused_tx_parallel_data(108),                                                                                                                                                                                                                                                                                                                                                                                       --                   .tx_parallel_data
			tx_parallel_data(309)     => unused_tx_parallel_data(109),                                                                                                                                                                                                                                                                                                                                                                                       --                   .tx_parallel_data
			tx_parallel_data(310)     => unused_tx_parallel_data(110),                                                                                                                                                                                                                                                                                                                                                                                       --                   .tx_parallel_data
			tx_parallel_data(311)     => unused_tx_parallel_data(111),                                                                                                                                                                                                                                                                                                                                                                                       --                   .tx_parallel_data
			tx_parallel_data(312)     => unused_tx_parallel_data(112),                                                                                                                                                                                                                                                                                                                                                                                       --                   .tx_parallel_data
			tx_parallel_data(313)     => unused_tx_parallel_data(113),                                                                                                                                                                                                                                                                                                                                                                                       --                   .tx_parallel_data
			tx_parallel_data(314)     => unused_tx_parallel_data(114),                                                                                                                                                                                                                                                                                                                                                                                       --                   .tx_parallel_data
			tx_parallel_data(315)     => unused_tx_parallel_data(115),                                                                                                                                                                                                                                                                                                                                                                                       --                   .tx_parallel_data
			tx_parallel_data(316)     => unused_tx_parallel_data(116),                                                                                                                                                                                                                                                                                                                                                                                       --                   .tx_parallel_data
			tx_parallel_data(317)     => unused_tx_parallel_data(117),                                                                                                                                                                                                                                                                                                                                                                                       --                   .tx_parallel_data
			tx_parallel_data(318)     => unused_tx_parallel_data(118),                                                                                                                                                                                                                                                                                                                                                                                       --                   .tx_parallel_data
			tx_parallel_data(319)     => unused_tx_parallel_data(119),                                                                                                                                                                                                                                                                                                                                                                                       --                   .tx_parallel_data
			rx_parallel_data(0)       => gx_std_x5_inst_rx_parallel_data(0),                                                                                                                                                                                                                                                                                                                                                                                 --   rx_parallel_data.rx_parallel_data
			rx_parallel_data(1)       => gx_std_x5_inst_rx_parallel_data(1),                                                                                                                                                                                                                                                                                                                                                                                 --                   .rx_parallel_data
			rx_parallel_data(2)       => gx_std_x5_inst_rx_parallel_data(2),                                                                                                                                                                                                                                                                                                                                                                                 --                   .rx_parallel_data
			rx_parallel_data(3)       => gx_std_x5_inst_rx_parallel_data(3),                                                                                                                                                                                                                                                                                                                                                                                 --                   .rx_parallel_data
			rx_parallel_data(4)       => gx_std_x5_inst_rx_parallel_data(4),                                                                                                                                                                                                                                                                                                                                                                                 --                   .rx_parallel_data
			rx_parallel_data(5)       => gx_std_x5_inst_rx_parallel_data(5),                                                                                                                                                                                                                                                                                                                                                                                 --                   .rx_parallel_data
			rx_parallel_data(6)       => gx_std_x5_inst_rx_parallel_data(6),                                                                                                                                                                                                                                                                                                                                                                                 --                   .rx_parallel_data
			rx_parallel_data(7)       => gx_std_x5_inst_rx_parallel_data(7),                                                                                                                                                                                                                                                                                                                                                                                 --                   .rx_parallel_data
			rx_parallel_data(8)       => gx_std_x5_inst_rx_parallel_data(8),                                                                                                                                                                                                                                                                                                                                                                                 --                   .rx_parallel_data
			rx_parallel_data(9)       => gx_std_x5_inst_rx_parallel_data(9),                                                                                                                                                                                                                                                                                                                                                                                 --                   .rx_parallel_data
			rx_parallel_data(10)      => gx_std_x5_inst_rx_parallel_data(10),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(11)      => gx_std_x5_inst_rx_parallel_data(11),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(12)      => gx_std_x5_inst_rx_parallel_data(12),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(13)      => gx_std_x5_inst_rx_parallel_data(13),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(14)      => gx_std_x5_inst_rx_parallel_data(14),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(15)      => gx_std_x5_inst_rx_parallel_data(15),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(16)      => gx_std_x5_inst_rx_parallel_data(16),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(17)      => gx_std_x5_inst_rx_parallel_data(17),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(18)      => gx_std_x5_inst_rx_parallel_data(18),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(19)      => gx_std_x5_inst_rx_parallel_data(19),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(20)      => gx_std_x5_inst_rx_parallel_data(20),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(21)      => gx_std_x5_inst_rx_parallel_data(21),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(22)      => gx_std_x5_inst_rx_parallel_data(22),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(23)      => gx_std_x5_inst_rx_parallel_data(23),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(24)      => gx_std_x5_inst_rx_parallel_data(24),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(25)      => gx_std_x5_inst_rx_parallel_data(25),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(26)      => gx_std_x5_inst_rx_parallel_data(26),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(27)      => gx_std_x5_inst_rx_parallel_data(27),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(28)      => gx_std_x5_inst_rx_parallel_data(28),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(29)      => gx_std_x5_inst_rx_parallel_data(29),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(30)      => gx_std_x5_inst_rx_parallel_data(30),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(31)      => gx_std_x5_inst_rx_parallel_data(31),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(32)      => gx_std_x5_inst_rx_parallel_data(32),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(33)      => gx_std_x5_inst_rx_parallel_data(33),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(34)      => gx_std_x5_inst_rx_parallel_data(34),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(35)      => gx_std_x5_inst_rx_parallel_data(35),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(36)      => gx_std_x5_inst_rx_parallel_data(36),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(37)      => gx_std_x5_inst_rx_parallel_data(37),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(38)      => gx_std_x5_inst_rx_parallel_data(38),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(39)      => gx_std_x5_inst_rx_parallel_data(39),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(40)      => gx_std_x5_inst_rx_parallel_data(40),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(41)      => gx_std_x5_inst_rx_parallel_data(41),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(42)      => gx_std_x5_inst_rx_parallel_data(42),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(43)      => gx_std_x5_inst_rx_parallel_data(43),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(44)      => gx_std_x5_inst_rx_parallel_data(44),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(45)      => gx_std_x5_inst_rx_parallel_data(45),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(46)      => gx_std_x5_inst_rx_parallel_data(46),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(47)      => gx_std_x5_inst_rx_parallel_data(47),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(48)      => gx_std_x5_inst_rx_parallel_data(48),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(49)      => gx_std_x5_inst_rx_parallel_data(49),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(50)      => gx_std_x5_inst_rx_parallel_data(50),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(51)      => gx_std_x5_inst_rx_parallel_data(51),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(52)      => gx_std_x5_inst_rx_parallel_data(52),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(53)      => gx_std_x5_inst_rx_parallel_data(53),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(54)      => gx_std_x5_inst_rx_parallel_data(54),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(55)      => gx_std_x5_inst_rx_parallel_data(55),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(56)      => gx_std_x5_inst_rx_parallel_data(56),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(57)      => gx_std_x5_inst_rx_parallel_data(57),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(58)      => gx_std_x5_inst_rx_parallel_data(58),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(59)      => gx_std_x5_inst_rx_parallel_data(59),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(60)      => gx_std_x5_inst_rx_parallel_data(60),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(61)      => gx_std_x5_inst_rx_parallel_data(61),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(62)      => gx_std_x5_inst_rx_parallel_data(62),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(63)      => gx_std_x5_inst_rx_parallel_data(63),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(64)      => gx_std_x5_inst_rx_parallel_data(64),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(65)      => gx_std_x5_inst_rx_parallel_data(65),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(66)      => gx_std_x5_inst_rx_parallel_data(66),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(67)      => gx_std_x5_inst_rx_parallel_data(67),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(68)      => gx_std_x5_inst_rx_parallel_data(68),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(69)      => gx_std_x5_inst_rx_parallel_data(69),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(70)      => gx_std_x5_inst_rx_parallel_data(70),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(71)      => gx_std_x5_inst_rx_parallel_data(71),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(72)      => gx_std_x5_inst_rx_parallel_data(72),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(73)      => gx_std_x5_inst_rx_parallel_data(73),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(74)      => gx_std_x5_inst_rx_parallel_data(74),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(75)      => gx_std_x5_inst_rx_parallel_data(75),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(76)      => gx_std_x5_inst_rx_parallel_data(76),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(77)      => gx_std_x5_inst_rx_parallel_data(77),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(78)      => gx_std_x5_inst_rx_parallel_data(78),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(79)      => gx_std_x5_inst_rx_parallel_data(79),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(80)      => gx_std_x5_inst_rx_parallel_data(80),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(81)      => gx_std_x5_inst_rx_parallel_data(81),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(82)      => gx_std_x5_inst_rx_parallel_data(82),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(83)      => gx_std_x5_inst_rx_parallel_data(83),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(84)      => gx_std_x5_inst_rx_parallel_data(84),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(85)      => gx_std_x5_inst_rx_parallel_data(85),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(86)      => gx_std_x5_inst_rx_parallel_data(86),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(87)      => gx_std_x5_inst_rx_parallel_data(87),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(88)      => gx_std_x5_inst_rx_parallel_data(88),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(89)      => gx_std_x5_inst_rx_parallel_data(89),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(90)      => gx_std_x5_inst_rx_parallel_data(90),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(91)      => gx_std_x5_inst_rx_parallel_data(91),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(92)      => gx_std_x5_inst_rx_parallel_data(92),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(93)      => gx_std_x5_inst_rx_parallel_data(93),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(94)      => gx_std_x5_inst_rx_parallel_data(94),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(95)      => gx_std_x5_inst_rx_parallel_data(95),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(96)      => gx_std_x5_inst_rx_parallel_data(96),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(97)      => gx_std_x5_inst_rx_parallel_data(97),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(98)      => gx_std_x5_inst_rx_parallel_data(98),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(99)      => gx_std_x5_inst_rx_parallel_data(99),                                                                                                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(100)     => gx_std_x5_inst_rx_parallel_data(100),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(101)     => gx_std_x5_inst_rx_parallel_data(101),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(102)     => gx_std_x5_inst_rx_parallel_data(102),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(103)     => gx_std_x5_inst_rx_parallel_data(103),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(104)     => gx_std_x5_inst_rx_parallel_data(104),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(105)     => gx_std_x5_inst_rx_parallel_data(105),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(106)     => gx_std_x5_inst_rx_parallel_data(106),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(107)     => gx_std_x5_inst_rx_parallel_data(107),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(108)     => gx_std_x5_inst_rx_parallel_data(108),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(109)     => gx_std_x5_inst_rx_parallel_data(109),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(110)     => gx_std_x5_inst_rx_parallel_data(110),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(111)     => gx_std_x5_inst_rx_parallel_data(111),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(112)     => gx_std_x5_inst_rx_parallel_data(112),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(113)     => gx_std_x5_inst_rx_parallel_data(113),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(114)     => gx_std_x5_inst_rx_parallel_data(114),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(115)     => gx_std_x5_inst_rx_parallel_data(115),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(116)     => gx_std_x5_inst_rx_parallel_data(116),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(117)     => gx_std_x5_inst_rx_parallel_data(117),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(118)     => gx_std_x5_inst_rx_parallel_data(118),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(119)     => gx_std_x5_inst_rx_parallel_data(119),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(120)     => gx_std_x5_inst_rx_parallel_data(120),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(121)     => gx_std_x5_inst_rx_parallel_data(121),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(122)     => gx_std_x5_inst_rx_parallel_data(122),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(123)     => gx_std_x5_inst_rx_parallel_data(123),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(124)     => gx_std_x5_inst_rx_parallel_data(124),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(125)     => gx_std_x5_inst_rx_parallel_data(125),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(126)     => gx_std_x5_inst_rx_parallel_data(126),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(127)     => gx_std_x5_inst_rx_parallel_data(127),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(128)     => gx_std_x5_inst_rx_parallel_data(128),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(129)     => gx_std_x5_inst_rx_parallel_data(129),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(130)     => gx_std_x5_inst_rx_parallel_data(130),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(131)     => gx_std_x5_inst_rx_parallel_data(131),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(132)     => gx_std_x5_inst_rx_parallel_data(132),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(133)     => gx_std_x5_inst_rx_parallel_data(133),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(134)     => gx_std_x5_inst_rx_parallel_data(134),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(135)     => gx_std_x5_inst_rx_parallel_data(135),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(136)     => gx_std_x5_inst_rx_parallel_data(136),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(137)     => gx_std_x5_inst_rx_parallel_data(137),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(138)     => gx_std_x5_inst_rx_parallel_data(138),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(139)     => gx_std_x5_inst_rx_parallel_data(139),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(140)     => gx_std_x5_inst_rx_parallel_data(140),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(141)     => gx_std_x5_inst_rx_parallel_data(141),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(142)     => gx_std_x5_inst_rx_parallel_data(142),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(143)     => gx_std_x5_inst_rx_parallel_data(143),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(144)     => gx_std_x5_inst_rx_parallel_data(144),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(145)     => gx_std_x5_inst_rx_parallel_data(145),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(146)     => gx_std_x5_inst_rx_parallel_data(146),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(147)     => gx_std_x5_inst_rx_parallel_data(147),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(148)     => gx_std_x5_inst_rx_parallel_data(148),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(149)     => gx_std_x5_inst_rx_parallel_data(149),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(150)     => gx_std_x5_inst_rx_parallel_data(150),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(151)     => gx_std_x5_inst_rx_parallel_data(151),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(152)     => gx_std_x5_inst_rx_parallel_data(152),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(153)     => gx_std_x5_inst_rx_parallel_data(153),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(154)     => gx_std_x5_inst_rx_parallel_data(154),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(155)     => gx_std_x5_inst_rx_parallel_data(155),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(156)     => gx_std_x5_inst_rx_parallel_data(156),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(157)     => gx_std_x5_inst_rx_parallel_data(157),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(158)     => gx_std_x5_inst_rx_parallel_data(158),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(159)     => gx_std_x5_inst_rx_parallel_data(159),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(160)     => gx_std_x5_inst_rx_parallel_data(160),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(161)     => gx_std_x5_inst_rx_parallel_data(161),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(162)     => gx_std_x5_inst_rx_parallel_data(162),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(163)     => gx_std_x5_inst_rx_parallel_data(163),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(164)     => gx_std_x5_inst_rx_parallel_data(164),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(165)     => gx_std_x5_inst_rx_parallel_data(165),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(166)     => gx_std_x5_inst_rx_parallel_data(166),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(167)     => gx_std_x5_inst_rx_parallel_data(167),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(168)     => gx_std_x5_inst_rx_parallel_data(168),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(169)     => gx_std_x5_inst_rx_parallel_data(169),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(170)     => gx_std_x5_inst_rx_parallel_data(170),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(171)     => gx_std_x5_inst_rx_parallel_data(171),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(172)     => gx_std_x5_inst_rx_parallel_data(172),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(173)     => gx_std_x5_inst_rx_parallel_data(173),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(174)     => gx_std_x5_inst_rx_parallel_data(174),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(175)     => gx_std_x5_inst_rx_parallel_data(175),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(176)     => gx_std_x5_inst_rx_parallel_data(176),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(177)     => gx_std_x5_inst_rx_parallel_data(177),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(178)     => gx_std_x5_inst_rx_parallel_data(178),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(179)     => gx_std_x5_inst_rx_parallel_data(179),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(180)     => gx_std_x5_inst_rx_parallel_data(180),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(181)     => gx_std_x5_inst_rx_parallel_data(181),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(182)     => gx_std_x5_inst_rx_parallel_data(182),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(183)     => gx_std_x5_inst_rx_parallel_data(183),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(184)     => gx_std_x5_inst_rx_parallel_data(184),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(185)     => gx_std_x5_inst_rx_parallel_data(185),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(186)     => gx_std_x5_inst_rx_parallel_data(186),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(187)     => gx_std_x5_inst_rx_parallel_data(187),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(188)     => gx_std_x5_inst_rx_parallel_data(188),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(189)     => gx_std_x5_inst_rx_parallel_data(189),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(190)     => gx_std_x5_inst_rx_parallel_data(190),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(191)     => gx_std_x5_inst_rx_parallel_data(191),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(192)     => gx_std_x5_inst_rx_parallel_data(192),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(193)     => gx_std_x5_inst_rx_parallel_data(193),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(194)     => gx_std_x5_inst_rx_parallel_data(194),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(195)     => gx_std_x5_inst_rx_parallel_data(195),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(196)     => gx_std_x5_inst_rx_parallel_data(196),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(197)     => gx_std_x5_inst_rx_parallel_data(197),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(198)     => gx_std_x5_inst_rx_parallel_data(198),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(199)     => gx_std_x5_inst_rx_parallel_data(199),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(200)     => gx_std_x5_inst_rx_parallel_data(200),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(201)     => gx_std_x5_inst_rx_parallel_data(201),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(202)     => gx_std_x5_inst_rx_parallel_data(202),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(203)     => gx_std_x5_inst_rx_parallel_data(203),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(204)     => gx_std_x5_inst_rx_parallel_data(204),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(205)     => gx_std_x5_inst_rx_parallel_data(205),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(206)     => gx_std_x5_inst_rx_parallel_data(206),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(207)     => gx_std_x5_inst_rx_parallel_data(207),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(208)     => gx_std_x5_inst_rx_parallel_data(208),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(209)     => gx_std_x5_inst_rx_parallel_data(209),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(210)     => gx_std_x5_inst_rx_parallel_data(210),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(211)     => gx_std_x5_inst_rx_parallel_data(211),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(212)     => gx_std_x5_inst_rx_parallel_data(212),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(213)     => gx_std_x5_inst_rx_parallel_data(213),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(214)     => gx_std_x5_inst_rx_parallel_data(214),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(215)     => gx_std_x5_inst_rx_parallel_data(215),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(216)     => gx_std_x5_inst_rx_parallel_data(216),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(217)     => gx_std_x5_inst_rx_parallel_data(217),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(218)     => gx_std_x5_inst_rx_parallel_data(218),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(219)     => gx_std_x5_inst_rx_parallel_data(219),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(220)     => gx_std_x5_inst_rx_parallel_data(220),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(221)     => gx_std_x5_inst_rx_parallel_data(221),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(222)     => gx_std_x5_inst_rx_parallel_data(222),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(223)     => gx_std_x5_inst_rx_parallel_data(223),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(224)     => gx_std_x5_inst_rx_parallel_data(224),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(225)     => gx_std_x5_inst_rx_parallel_data(225),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(226)     => gx_std_x5_inst_rx_parallel_data(226),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(227)     => gx_std_x5_inst_rx_parallel_data(227),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(228)     => gx_std_x5_inst_rx_parallel_data(228),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(229)     => gx_std_x5_inst_rx_parallel_data(229),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(230)     => gx_std_x5_inst_rx_parallel_data(230),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(231)     => gx_std_x5_inst_rx_parallel_data(231),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(232)     => gx_std_x5_inst_rx_parallel_data(232),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(233)     => gx_std_x5_inst_rx_parallel_data(233),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(234)     => gx_std_x5_inst_rx_parallel_data(234),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(235)     => gx_std_x5_inst_rx_parallel_data(235),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(236)     => gx_std_x5_inst_rx_parallel_data(236),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(237)     => gx_std_x5_inst_rx_parallel_data(237),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(238)     => gx_std_x5_inst_rx_parallel_data(238),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(239)     => gx_std_x5_inst_rx_parallel_data(239),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(240)     => gx_std_x5_inst_rx_parallel_data(240),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(241)     => gx_std_x5_inst_rx_parallel_data(241),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(242)     => gx_std_x5_inst_rx_parallel_data(242),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(243)     => gx_std_x5_inst_rx_parallel_data(243),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(244)     => gx_std_x5_inst_rx_parallel_data(244),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(245)     => gx_std_x5_inst_rx_parallel_data(245),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(246)     => gx_std_x5_inst_rx_parallel_data(246),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(247)     => gx_std_x5_inst_rx_parallel_data(247),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(248)     => gx_std_x5_inst_rx_parallel_data(248),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(249)     => gx_std_x5_inst_rx_parallel_data(249),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(250)     => gx_std_x5_inst_rx_parallel_data(250),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(251)     => gx_std_x5_inst_rx_parallel_data(251),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(252)     => gx_std_x5_inst_rx_parallel_data(252),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(253)     => gx_std_x5_inst_rx_parallel_data(253),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(254)     => gx_std_x5_inst_rx_parallel_data(254),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(255)     => gx_std_x5_inst_rx_parallel_data(255),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(256)     => gx_std_x5_inst_rx_parallel_data(256),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(257)     => gx_std_x5_inst_rx_parallel_data(257),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(258)     => gx_std_x5_inst_rx_parallel_data(258),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(259)     => gx_std_x5_inst_rx_parallel_data(259),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(260)     => gx_std_x5_inst_rx_parallel_data(260),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(261)     => gx_std_x5_inst_rx_parallel_data(261),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(262)     => gx_std_x5_inst_rx_parallel_data(262),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(263)     => gx_std_x5_inst_rx_parallel_data(263),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(264)     => gx_std_x5_inst_rx_parallel_data(264),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(265)     => gx_std_x5_inst_rx_parallel_data(265),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(266)     => gx_std_x5_inst_rx_parallel_data(266),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(267)     => gx_std_x5_inst_rx_parallel_data(267),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(268)     => gx_std_x5_inst_rx_parallel_data(268),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(269)     => gx_std_x5_inst_rx_parallel_data(269),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(270)     => gx_std_x5_inst_rx_parallel_data(270),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(271)     => gx_std_x5_inst_rx_parallel_data(271),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(272)     => gx_std_x5_inst_rx_parallel_data(272),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(273)     => gx_std_x5_inst_rx_parallel_data(273),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(274)     => gx_std_x5_inst_rx_parallel_data(274),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(275)     => gx_std_x5_inst_rx_parallel_data(275),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(276)     => gx_std_x5_inst_rx_parallel_data(276),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(277)     => gx_std_x5_inst_rx_parallel_data(277),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(278)     => gx_std_x5_inst_rx_parallel_data(278),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(279)     => gx_std_x5_inst_rx_parallel_data(279),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(280)     => gx_std_x5_inst_rx_parallel_data(280),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(281)     => gx_std_x5_inst_rx_parallel_data(281),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(282)     => gx_std_x5_inst_rx_parallel_data(282),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(283)     => gx_std_x5_inst_rx_parallel_data(283),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(284)     => gx_std_x5_inst_rx_parallel_data(284),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(285)     => gx_std_x5_inst_rx_parallel_data(285),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(286)     => gx_std_x5_inst_rx_parallel_data(286),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(287)     => gx_std_x5_inst_rx_parallel_data(287),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(288)     => gx_std_x5_inst_rx_parallel_data(288),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(289)     => gx_std_x5_inst_rx_parallel_data(289),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(290)     => gx_std_x5_inst_rx_parallel_data(290),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(291)     => gx_std_x5_inst_rx_parallel_data(291),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(292)     => gx_std_x5_inst_rx_parallel_data(292),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(293)     => gx_std_x5_inst_rx_parallel_data(293),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(294)     => gx_std_x5_inst_rx_parallel_data(294),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(295)     => gx_std_x5_inst_rx_parallel_data(295),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(296)     => gx_std_x5_inst_rx_parallel_data(296),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(297)     => gx_std_x5_inst_rx_parallel_data(297),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(298)     => gx_std_x5_inst_rx_parallel_data(298),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(299)     => gx_std_x5_inst_rx_parallel_data(299),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(300)     => gx_std_x5_inst_rx_parallel_data(300),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(301)     => gx_std_x5_inst_rx_parallel_data(301),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(302)     => gx_std_x5_inst_rx_parallel_data(302),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(303)     => gx_std_x5_inst_rx_parallel_data(303),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(304)     => gx_std_x5_inst_rx_parallel_data(304),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(305)     => gx_std_x5_inst_rx_parallel_data(305),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(306)     => gx_std_x5_inst_rx_parallel_data(306),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(307)     => gx_std_x5_inst_rx_parallel_data(307),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(308)     => gx_std_x5_inst_rx_parallel_data(308),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(309)     => gx_std_x5_inst_rx_parallel_data(309),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(310)     => gx_std_x5_inst_rx_parallel_data(310),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(311)     => gx_std_x5_inst_rx_parallel_data(311),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(312)     => gx_std_x5_inst_rx_parallel_data(312),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(313)     => gx_std_x5_inst_rx_parallel_data(313),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(314)     => gx_std_x5_inst_rx_parallel_data(314),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(315)     => gx_std_x5_inst_rx_parallel_data(315),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(316)     => gx_std_x5_inst_rx_parallel_data(316),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(317)     => gx_std_x5_inst_rx_parallel_data(317),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(318)     => gx_std_x5_inst_rx_parallel_data(318),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(319)     => gx_std_x5_inst_rx_parallel_data(319),                                                                                                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			tx_pll_refclk             => "0",                                                                                                                                                                                                                                                                                                                                                                                                                --        (terminated)
			tx_pma_clkout             => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_pma_pclk               => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_pma_parallel_data      => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", --        (terminated)
			pll_locked                => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_pma_clkout             => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_pma_pclk               => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_pma_parallel_data      => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_clkslip                => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			rx_clklow                 => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_fref                   => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_set_locktodata         => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			rx_set_locktoref          => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			rx_signaldetect           => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_pma_qpipulldn          => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			tx_pma_qpipullup          => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			tx_pma_qpipulldn          => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			tx_pma_txdetectrx         => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			tx_pma_rxfound            => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_prbs_done          => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_prbs_err           => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_std_pcfifo_full        => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_std_pcfifo_empty       => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_pcfifo_full        => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_pcfifo_empty       => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_byteorder_ena      => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			rx_std_byteorder_flag     => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_rmfifo_full        => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_rmfifo_empty       => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_wa_patternalign    => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			rx_std_wa_a1a2size        => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			tx_std_bitslipboundarysel => "0000000000000000000000000",                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			rx_std_bitslipboundarysel => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_bitslip            => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			rx_std_runlength_err      => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_bitrev_ena         => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			rx_std_byterev_ena        => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			tx_std_elecidle           => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			rx_std_signaldetect       => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_10g_coreclkin          => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			rx_10g_coreclkin          => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			tx_10g_clkout             => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_clkout             => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_clk33out           => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_prbs_err_clr       => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			rx_10g_prbs_done          => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_prbs_err           => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_10g_control            => "000000000000000000000000000000000000000000000",                                                                                                                                                                                                                                                                                                                                                                    --        (terminated)
			rx_10g_control            => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_10g_data_valid         => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			tx_10g_fifo_full          => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_10g_fifo_pfull         => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_10g_fifo_empty         => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_10g_fifo_pempty        => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_10g_fifo_del           => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_10g_fifo_insert        => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_fifo_rd_en         => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			rx_10g_data_valid         => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_fifo_full          => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_fifo_pfull         => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_fifo_empty         => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_fifo_pempty        => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_fifo_del           => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_fifo_insert        => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_fifo_align_val     => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_fifo_align_clr     => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			rx_10g_fifo_align_en      => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			tx_10g_frame              => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_10g_frame_diag_status  => "0000000000",                                                                                                                                                                                                                                                                                                                                                                                                       --        (terminated)
			tx_10g_frame_burst_en     => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			rx_10g_frame              => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_frame_lock         => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_frame_mfrm_err     => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_frame_sync_err     => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_frame_skip_ins     => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_frame_pyld_ins     => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_frame_skip_err     => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_frame_diag_err     => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_frame_diag_status  => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_crc32_err          => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_descram_err        => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_blk_lock           => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_blk_sh_err         => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_10g_bitslip            => "00000000000000000000000000000000000",                                                                                                                                                                                                                                                                                                                                                                              --        (terminated)
			rx_10g_bitslip            => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			rx_10g_highber            => open,                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_highber_clr_cnt    => "00000",                                                                                                                                                                                                                                                                                                                                                                                                            --        (terminated)
			rx_10g_clr_errblk_count   => "00000"                                                                                                                                                                                                                                                                                                                                                                                                             --        (terminated)
		);

	rx_parallel_data <= gx_std_x5_inst_rx_parallel_data(313) & gx_std_x5_inst_rx_parallel_data(312) & gx_std_x5_inst_rx_parallel_data(311) & gx_std_x5_inst_rx_parallel_data(310) & gx_std_x5_inst_rx_parallel_data(309) & gx_std_x5_inst_rx_parallel_data(308) & gx_std_x5_inst_rx_parallel_data(307) & gx_std_x5_inst_rx_parallel_data(306) & gx_std_x5_inst_rx_parallel_data(305) & gx_std_x5_inst_rx_parallel_data(304) & gx_std_x5_inst_rx_parallel_data(297) & gx_std_x5_inst_rx_parallel_data(296) & gx_std_x5_inst_rx_parallel_data(295) & gx_std_x5_inst_rx_parallel_data(294) & gx_std_x5_inst_rx_parallel_data(293) & gx_std_x5_inst_rx_parallel_data(292) & gx_std_x5_inst_rx_parallel_data(291) & gx_std_x5_inst_rx_parallel_data(290) & gx_std_x5_inst_rx_parallel_data(289) & gx_std_x5_inst_rx_parallel_data(288) & gx_std_x5_inst_rx_parallel_data(281) & gx_std_x5_inst_rx_parallel_data(280) & gx_std_x5_inst_rx_parallel_data(279) & gx_std_x5_inst_rx_parallel_data(278) & gx_std_x5_inst_rx_parallel_data(277) & gx_std_x5_inst_rx_parallel_data(276) & gx_std_x5_inst_rx_parallel_data(275) & gx_std_x5_inst_rx_parallel_data(274) & gx_std_x5_inst_rx_parallel_data(273) & gx_std_x5_inst_rx_parallel_data(272) & gx_std_x5_inst_rx_parallel_data(265) & gx_std_x5_inst_rx_parallel_data(264) & gx_std_x5_inst_rx_parallel_data(263) & gx_std_x5_inst_rx_parallel_data(262) & gx_std_x5_inst_rx_parallel_data(261) & gx_std_x5_inst_rx_parallel_data(260) & gx_std_x5_inst_rx_parallel_data(259) & gx_std_x5_inst_rx_parallel_data(258) & gx_std_x5_inst_rx_parallel_data(257) & gx_std_x5_inst_rx_parallel_data(256) & gx_std_x5_inst_rx_parallel_data(249) & gx_std_x5_inst_rx_parallel_data(248) & gx_std_x5_inst_rx_parallel_data(247) & gx_std_x5_inst_rx_parallel_data(246) & gx_std_x5_inst_rx_parallel_data(245) & gx_std_x5_inst_rx_parallel_data(244) & gx_std_x5_inst_rx_parallel_data(243) & gx_std_x5_inst_rx_parallel_data(242) & gx_std_x5_inst_rx_parallel_data(241) & gx_std_x5_inst_rx_parallel_data(240) & gx_std_x5_inst_rx_parallel_data(233) & gx_std_x5_inst_rx_parallel_data(232) & gx_std_x5_inst_rx_parallel_data(231) & gx_std_x5_inst_rx_parallel_data(230) & gx_std_x5_inst_rx_parallel_data(229) & gx_std_x5_inst_rx_parallel_data(228) & gx_std_x5_inst_rx_parallel_data(227) & gx_std_x5_inst_rx_parallel_data(226) & gx_std_x5_inst_rx_parallel_data(225) & gx_std_x5_inst_rx_parallel_data(224) & gx_std_x5_inst_rx_parallel_data(217) & gx_std_x5_inst_rx_parallel_data(216) & gx_std_x5_inst_rx_parallel_data(215) & gx_std_x5_inst_rx_parallel_data(214) & gx_std_x5_inst_rx_parallel_data(213) & gx_std_x5_inst_rx_parallel_data(212) & gx_std_x5_inst_rx_parallel_data(211) & gx_std_x5_inst_rx_parallel_data(210) & gx_std_x5_inst_rx_parallel_data(209) & gx_std_x5_inst_rx_parallel_data(208) & gx_std_x5_inst_rx_parallel_data(201) & gx_std_x5_inst_rx_parallel_data(200) & gx_std_x5_inst_rx_parallel_data(199) & gx_std_x5_inst_rx_parallel_data(198) & gx_std_x5_inst_rx_parallel_data(197) & gx_std_x5_inst_rx_parallel_data(196) & gx_std_x5_inst_rx_parallel_data(195) & gx_std_x5_inst_rx_parallel_data(194) & gx_std_x5_inst_rx_parallel_data(193) & gx_std_x5_inst_rx_parallel_data(192) & gx_std_x5_inst_rx_parallel_data(185) & gx_std_x5_inst_rx_parallel_data(184) & gx_std_x5_inst_rx_parallel_data(183) & gx_std_x5_inst_rx_parallel_data(182) & gx_std_x5_inst_rx_parallel_data(181) & gx_std_x5_inst_rx_parallel_data(180) & gx_std_x5_inst_rx_parallel_data(179) & gx_std_x5_inst_rx_parallel_data(178) & gx_std_x5_inst_rx_parallel_data(177) & gx_std_x5_inst_rx_parallel_data(176) & gx_std_x5_inst_rx_parallel_data(169) & gx_std_x5_inst_rx_parallel_data(168) & gx_std_x5_inst_rx_parallel_data(167) & gx_std_x5_inst_rx_parallel_data(166) & gx_std_x5_inst_rx_parallel_data(165) & gx_std_x5_inst_rx_parallel_data(164) & gx_std_x5_inst_rx_parallel_data(163) & gx_std_x5_inst_rx_parallel_data(162) & gx_std_x5_inst_rx_parallel_data(161) & gx_std_x5_inst_rx_parallel_data(160) & gx_std_x5_inst_rx_parallel_data(153) & gx_std_x5_inst_rx_parallel_data(152) & gx_std_x5_inst_rx_parallel_data(151) & gx_std_x5_inst_rx_parallel_data(150) & gx_std_x5_inst_rx_parallel_data(149) & gx_std_x5_inst_rx_parallel_data(148) & gx_std_x5_inst_rx_parallel_data(147) & gx_std_x5_inst_rx_parallel_data(146) & gx_std_x5_inst_rx_parallel_data(145) & gx_std_x5_inst_rx_parallel_data(144) & gx_std_x5_inst_rx_parallel_data(137) & gx_std_x5_inst_rx_parallel_data(136) & gx_std_x5_inst_rx_parallel_data(135) & gx_std_x5_inst_rx_parallel_data(134) & gx_std_x5_inst_rx_parallel_data(133) & gx_std_x5_inst_rx_parallel_data(132) & gx_std_x5_inst_rx_parallel_data(131) & gx_std_x5_inst_rx_parallel_data(130) & gx_std_x5_inst_rx_parallel_data(129) & gx_std_x5_inst_rx_parallel_data(128) & gx_std_x5_inst_rx_parallel_data(121) & gx_std_x5_inst_rx_parallel_data(120) & gx_std_x5_inst_rx_parallel_data(119) & gx_std_x5_inst_rx_parallel_data(118) & gx_std_x5_inst_rx_parallel_data(117) & gx_std_x5_inst_rx_parallel_data(116) & gx_std_x5_inst_rx_parallel_data(115) & gx_std_x5_inst_rx_parallel_data(114) & gx_std_x5_inst_rx_parallel_data(113) & gx_std_x5_inst_rx_parallel_data(112) & gx_std_x5_inst_rx_parallel_data(105) & gx_std_x5_inst_rx_parallel_data(104) & gx_std_x5_inst_rx_parallel_data(103) & gx_std_x5_inst_rx_parallel_data(102) & gx_std_x5_inst_rx_parallel_data(101) & gx_std_x5_inst_rx_parallel_data(100) & gx_std_x5_inst_rx_parallel_data(99) & gx_std_x5_inst_rx_parallel_data(98) & gx_std_x5_inst_rx_parallel_data(97) & gx_std_x5_inst_rx_parallel_data(96) & gx_std_x5_inst_rx_parallel_data(89) & gx_std_x5_inst_rx_parallel_data(88) & gx_std_x5_inst_rx_parallel_data(87) & gx_std_x5_inst_rx_parallel_data(86) & gx_std_x5_inst_rx_parallel_data(85) & gx_std_x5_inst_rx_parallel_data(84) & gx_std_x5_inst_rx_parallel_data(83) & gx_std_x5_inst_rx_parallel_data(82) & gx_std_x5_inst_rx_parallel_data(81) & gx_std_x5_inst_rx_parallel_data(80) & gx_std_x5_inst_rx_parallel_data(73) & gx_std_x5_inst_rx_parallel_data(72) & gx_std_x5_inst_rx_parallel_data(71) & gx_std_x5_inst_rx_parallel_data(70) & gx_std_x5_inst_rx_parallel_data(69) & gx_std_x5_inst_rx_parallel_data(68) & gx_std_x5_inst_rx_parallel_data(67) & gx_std_x5_inst_rx_parallel_data(66) & gx_std_x5_inst_rx_parallel_data(65) & gx_std_x5_inst_rx_parallel_data(64) & gx_std_x5_inst_rx_parallel_data(57) & gx_std_x5_inst_rx_parallel_data(56) & gx_std_x5_inst_rx_parallel_data(55) & gx_std_x5_inst_rx_parallel_data(54) & gx_std_x5_inst_rx_parallel_data(53) & gx_std_x5_inst_rx_parallel_data(52) & gx_std_x5_inst_rx_parallel_data(51) & gx_std_x5_inst_rx_parallel_data(50) & gx_std_x5_inst_rx_parallel_data(49) & gx_std_x5_inst_rx_parallel_data(48) & gx_std_x5_inst_rx_parallel_data(41) & gx_std_x5_inst_rx_parallel_data(40) & gx_std_x5_inst_rx_parallel_data(39) & gx_std_x5_inst_rx_parallel_data(38) & gx_std_x5_inst_rx_parallel_data(37) & gx_std_x5_inst_rx_parallel_data(36) & gx_std_x5_inst_rx_parallel_data(35) & gx_std_x5_inst_rx_parallel_data(34) & gx_std_x5_inst_rx_parallel_data(33) & gx_std_x5_inst_rx_parallel_data(32) & gx_std_x5_inst_rx_parallel_data(25) & gx_std_x5_inst_rx_parallel_data(24) & gx_std_x5_inst_rx_parallel_data(23) & gx_std_x5_inst_rx_parallel_data(22) & gx_std_x5_inst_rx_parallel_data(21) & gx_std_x5_inst_rx_parallel_data(20) & gx_std_x5_inst_rx_parallel_data(19) & gx_std_x5_inst_rx_parallel_data(18) & gx_std_x5_inst_rx_parallel_data(17) & gx_std_x5_inst_rx_parallel_data(16) & gx_std_x5_inst_rx_parallel_data(9) & gx_std_x5_inst_rx_parallel_data(8) & gx_std_x5_inst_rx_parallel_data(7) & gx_std_x5_inst_rx_parallel_data(6) & gx_std_x5_inst_rx_parallel_data(5) & gx_std_x5_inst_rx_parallel_data(4) & gx_std_x5_inst_rx_parallel_data(3) & gx_std_x5_inst_rx_parallel_data(2) & gx_std_x5_inst_rx_parallel_data(1) & gx_std_x5_inst_rx_parallel_data(0);

	unused_rx_parallel_data <= gx_std_x5_inst_rx_parallel_data(319) & gx_std_x5_inst_rx_parallel_data(318) & gx_std_x5_inst_rx_parallel_data(317) & gx_std_x5_inst_rx_parallel_data(316) & gx_std_x5_inst_rx_parallel_data(315) & gx_std_x5_inst_rx_parallel_data(314) & gx_std_x5_inst_rx_parallel_data(303) & gx_std_x5_inst_rx_parallel_data(302) & gx_std_x5_inst_rx_parallel_data(301) & gx_std_x5_inst_rx_parallel_data(300) & gx_std_x5_inst_rx_parallel_data(299) & gx_std_x5_inst_rx_parallel_data(298) & gx_std_x5_inst_rx_parallel_data(287) & gx_std_x5_inst_rx_parallel_data(286) & gx_std_x5_inst_rx_parallel_data(285) & gx_std_x5_inst_rx_parallel_data(284) & gx_std_x5_inst_rx_parallel_data(283) & gx_std_x5_inst_rx_parallel_data(282) & gx_std_x5_inst_rx_parallel_data(271) & gx_std_x5_inst_rx_parallel_data(270) & gx_std_x5_inst_rx_parallel_data(269) & gx_std_x5_inst_rx_parallel_data(268) & gx_std_x5_inst_rx_parallel_data(267) & gx_std_x5_inst_rx_parallel_data(266) & gx_std_x5_inst_rx_parallel_data(255) & gx_std_x5_inst_rx_parallel_data(254) & gx_std_x5_inst_rx_parallel_data(253) & gx_std_x5_inst_rx_parallel_data(252) & gx_std_x5_inst_rx_parallel_data(251) & gx_std_x5_inst_rx_parallel_data(250) & gx_std_x5_inst_rx_parallel_data(239) & gx_std_x5_inst_rx_parallel_data(238) & gx_std_x5_inst_rx_parallel_data(237) & gx_std_x5_inst_rx_parallel_data(236) & gx_std_x5_inst_rx_parallel_data(235) & gx_std_x5_inst_rx_parallel_data(234) & gx_std_x5_inst_rx_parallel_data(223) & gx_std_x5_inst_rx_parallel_data(222) & gx_std_x5_inst_rx_parallel_data(221) & gx_std_x5_inst_rx_parallel_data(220) & gx_std_x5_inst_rx_parallel_data(219) & gx_std_x5_inst_rx_parallel_data(218) & gx_std_x5_inst_rx_parallel_data(207) & gx_std_x5_inst_rx_parallel_data(206) & gx_std_x5_inst_rx_parallel_data(205) & gx_std_x5_inst_rx_parallel_data(204) & gx_std_x5_inst_rx_parallel_data(203) & gx_std_x5_inst_rx_parallel_data(202) & gx_std_x5_inst_rx_parallel_data(191) & gx_std_x5_inst_rx_parallel_data(190) & gx_std_x5_inst_rx_parallel_data(189) & gx_std_x5_inst_rx_parallel_data(188) & gx_std_x5_inst_rx_parallel_data(187) & gx_std_x5_inst_rx_parallel_data(186) & gx_std_x5_inst_rx_parallel_data(175) & gx_std_x5_inst_rx_parallel_data(174) & gx_std_x5_inst_rx_parallel_data(173) & gx_std_x5_inst_rx_parallel_data(172) & gx_std_x5_inst_rx_parallel_data(171) & gx_std_x5_inst_rx_parallel_data(170) & gx_std_x5_inst_rx_parallel_data(159) & gx_std_x5_inst_rx_parallel_data(158) & gx_std_x5_inst_rx_parallel_data(157) & gx_std_x5_inst_rx_parallel_data(156) & gx_std_x5_inst_rx_parallel_data(155) & gx_std_x5_inst_rx_parallel_data(154) & gx_std_x5_inst_rx_parallel_data(143) & gx_std_x5_inst_rx_parallel_data(142) & gx_std_x5_inst_rx_parallel_data(141) & gx_std_x5_inst_rx_parallel_data(140) & gx_std_x5_inst_rx_parallel_data(139) & gx_std_x5_inst_rx_parallel_data(138) & gx_std_x5_inst_rx_parallel_data(127) & gx_std_x5_inst_rx_parallel_data(126) & gx_std_x5_inst_rx_parallel_data(125) & gx_std_x5_inst_rx_parallel_data(124) & gx_std_x5_inst_rx_parallel_data(123) & gx_std_x5_inst_rx_parallel_data(122) & gx_std_x5_inst_rx_parallel_data(111) & gx_std_x5_inst_rx_parallel_data(110) & gx_std_x5_inst_rx_parallel_data(109) & gx_std_x5_inst_rx_parallel_data(108) & gx_std_x5_inst_rx_parallel_data(107) & gx_std_x5_inst_rx_parallel_data(106) & gx_std_x5_inst_rx_parallel_data(95) & gx_std_x5_inst_rx_parallel_data(94) & gx_std_x5_inst_rx_parallel_data(93) & gx_std_x5_inst_rx_parallel_data(92) & gx_std_x5_inst_rx_parallel_data(91) & gx_std_x5_inst_rx_parallel_data(90) & gx_std_x5_inst_rx_parallel_data(79) & gx_std_x5_inst_rx_parallel_data(78) & gx_std_x5_inst_rx_parallel_data(77) & gx_std_x5_inst_rx_parallel_data(76) & gx_std_x5_inst_rx_parallel_data(75) & gx_std_x5_inst_rx_parallel_data(74) & gx_std_x5_inst_rx_parallel_data(63) & gx_std_x5_inst_rx_parallel_data(62) & gx_std_x5_inst_rx_parallel_data(61) & gx_std_x5_inst_rx_parallel_data(60) & gx_std_x5_inst_rx_parallel_data(59) & gx_std_x5_inst_rx_parallel_data(58) & gx_std_x5_inst_rx_parallel_data(47) & gx_std_x5_inst_rx_parallel_data(46) & gx_std_x5_inst_rx_parallel_data(45) & gx_std_x5_inst_rx_parallel_data(44) & gx_std_x5_inst_rx_parallel_data(43) & gx_std_x5_inst_rx_parallel_data(42) & gx_std_x5_inst_rx_parallel_data(31) & gx_std_x5_inst_rx_parallel_data(30) & gx_std_x5_inst_rx_parallel_data(29) & gx_std_x5_inst_rx_parallel_data(28) & gx_std_x5_inst_rx_parallel_data(27) & gx_std_x5_inst_rx_parallel_data(26) & gx_std_x5_inst_rx_parallel_data(15) & gx_std_x5_inst_rx_parallel_data(14) & gx_std_x5_inst_rx_parallel_data(13) & gx_std_x5_inst_rx_parallel_data(12) & gx_std_x5_inst_rx_parallel_data(11) & gx_std_x5_inst_rx_parallel_data(10);

end architecture rtl; -- of gx_std_x5
