// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:09 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
caE6kBqqsc3Zhe0vFtP/H3nJySTBDgkWMd/EgLa4aty6oeZQ2E805SMocalZileK
2E4GNhtKdnwS3Aa/L8p0/DuhqYyS5QfC3/L4Q2q9MBNNP6Yqfg6a59Gf9HXXGaD+
gqPlXbMP3QqPKJ40TTlPDlVogGn1C+mbUrSlv3kA8yY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 104704)
T0h/x8K4hYyPAsyEw6iGzQTGeXmVA11JXdkhi+c5uCkhs0UjBoah1SyQrX0lyR3k
MKj2afuwpVRMvCpsHLvAgTJyT8gpdee9sUCOlu44UYB68LPFJy6Nh6HBJkQ5qkBZ
c9xL5k61MByjvckeJeu8C340kJq8tAfenuK1ZnjWlpq4+mmTZZAeMMkYEXjIbb09
PU3hBEUHLlbs+nyCjfOoRYi+2Q9NCJy6ykMmr+vFzO88AZYBlnF5mDy2O6Bzz1x3
HAQxUG4DBlBO2yzaslZAJWlYjLiNKDAwOZT2mwthP7HnZIpGFJzm6mGgpDsLqfNn
vKHCqCrmpIFQy2s7DFAzM1997Fs17Sc/Q3WPUlN73bh4WkOsQ4KPwSWpHDnG3WNt
WnMFmQm4R8dUd/lc4WyCmHz0On5vpTv/PbiHrHu80cPP2NhoYrOZiPSzYJZwbE/a
Jl9Ellviyh81M7B5IWGBxZfu9nwIzgoCFPtz+6b21VQUgtXDEGNFanijnd6sMLOE
Eg9X7yibhlyemVJVYfYrPqjjIM/LUrfmXzS4+ldkYGfAlFU/nUHMq4WfBtIPzTr3
tPeRDalSBZtbzK4nx5vBohKZhii9cVsak2KPniDsEr6+RX+5tVkgrPN23Wrj5IHt
Q1gaRDH4ucd7FnyMVC3iXAai4GlR9cgKxwbpiq+GMWItR+nvYoyXY6WqJTpF51uM
+/ofZJwuAtFqVMrUbfYJDSTTKLPTbZbN/RULTXYfkcLvD9Vgp7manzyvn9hmi719
abZ6uSp7X7k1vSFB0MUxMIXNvCRmRCD3KUw9Az7CXSN7fbk60SsAAP/5UXpWfL9s
vU+DR2QM31uXX5EGrdytdFCUaRSRKzu5udjD27goRCq8tYvRA0Xv9ZxE9nwMbalr
7knfGkH/ejRzS3IcYMC2+KI/A7PAudzPclwzNGRatYy0pWwcwhyR1Jzxkr1g/hE8
EXis351T5Hjp2qSysXDdw9/HspxNYqWRkg3qn2vEgbMw41I6znjaVmPM06YjHVKm
EHDH+kyaGTxkZlFXMI5aHASWQjigePBWeNOArch2BKScABRL1knu6E/Jvd/eWEl8
xtGt5iJ6yznIhajsNqOpTwS0rxsaZ/eDkvanvbBxAhvyU6WdcQ4kJP31BPLTSQ+S
W45D8Yl2GM42MWiRyzaAnvLXsNN5/LnWuordehS7yJVntixtuoCPFEk/xlM7Nt9N
81w6uA0Kz8zTI+ZAC4TjjyNroofMeHm7e4jpm50gyGF+8+FZN8R1oyYWs3Ca1TrY
3wixIDZ6GzIqu6GFOyTBNOvD4LDUX88+A/jRsY6QlUXPiQaI4XRAyAHDP2bxJue7
9uljZKOijmsWMSiReo4IyN1mAd1/b2S0HGQRIZMShLv+CkcNy+1ESTuoqJQaAWF4
y+qtMiXQDBx5I7FSKghbte8v15Woto5McrhWZMyxFqUBB0KNbsolOZWYa4d60zEv
IE9OqBwpPOvVg2iD0J8Pnxqus17yVjfBitI1eUy8Fbkpssw/aDBtRLUXyLJJrD2m
HHF/TI7Jnk11f+TeBt1ZHAU9SQOjKvO0UGNdCeLmSlTuKBMnByPA2ymckF4F/LxG
sYSO6gzBOyIdkIcdIg1trp7aLIpjHRJ76dcXHZzmyaCXQ+xZBIdMwQnYpp4uOXO5
/pLzoNL7NWOQlJz3m5DNGE1Y/lFP19eGmnvlJZ9azZsfTHKAiSDOklSwTzQ1Tx8a
po3OMgcts9siCV4WdDxSdB0VRktENZvvz+UdKn856dxpZ33kMNfMYY7TS1msTb+3
edYiFDlTGgPjKCVt/Nton+OrXeVIUgPLfPVmwqfMLOAwTMt6/kTSRWO8CgOdRh+F
0qnQhVdCRttczPJpsRwe5ZDBFLtYTZ66OqujlfIRqI/CJITjFunqW4XUShR58YCU
/rGzMFwVRDWwdY2VUAcvizV0ik2yVB+pFwViI9WL32Cr0a/ssYEjcdF6SPWqdmd9
0ANrZV3AFJSy4+Kfp/bRZzkxB9rEj29zLo0BOzEGlI3esr7kqOo7iIcrsea1lDCL
V51A0c2ONDmn6DFakHEVqpwANv6hcEy9x4xglYdkVPEeaRU6UHcuh3R4F49RiIQP
SfE8LNTLP/AYo+oOkTzUMDh1fB5+f0eXyI4wubhSKr/rHfMAJQlDUCJK14Go0MUk
YT9rCBVMNrVt90Ndeo75v4hFUuxaP4tjrzKN8gFUXim/x4EVjGc7WBkselEv92Pd
f8zjtabEwN2fr1U9BNIWLdFMzaQDZ+O4CaLMy1NQXdyKCGz0KHDzsOh4qEVJCVUF
CLiv+ZSLhHOjlVzF8S/d01b6E03GFw3fShAt9IP3FLgHwAW5VDw71k0jQl6VRRRW
PX1/jwSdlQ1VHZ8XM+qqHkOjfypkCwMTWMh44yVA/YeIQX0Y1RRme+I4TvxQv0pf
IZ9F/g07lpQrphKWbaF3pn/YOSR05SjCg7SWonYYcIaQK2FMHXvyF0TZ6teR2897
tQXAzSqxXJ6CyI6Km5wAfu/aQnYbPQPpjmP2gmcmg2PU1nNO4pQCS5eW+VFjyD+X
pLmOzKpjiiOcvtBaXifErzqNAT2mWbvYz5CwSy7VIJs85fvgj+GFw6/j3kDGo9TD
AdTezZZT5uEDqLHxYDfkP9qFAXCrgjjaGWz2/ihsy7VofSkLQVoERrXQBvTacJSw
Bol5Z+OFYc+beGuVic9MQ+AdrRsTnShPR38vLr3DDF5ZsdXp4cBZptE4f80LpN5f
ckLpErnp4O1ymHj1wfok2F4b5qFDO0clq+SJ7GtvcSi9tV9KcK2HZ5HUYByNcFoo
BAM+S964VpbGi/gXe03+oV1pbLfO0kkXnWuVPIpzFvZj91/FEy/pt6hs88scb7Fn
3FTm6KU049iWIjbteuwwkDHiTMkKbIoKDAg+r6hwrAOJirVVQoUI7RNhAvmfnRis
mBcYu6yDky3y1+Uaf5WuJwiq74Ksz4rT3CnWkpMDg64QhSS3uqSIrg2z69FaAGV8
CiDk+Tpj3v4h07y4Y/Rw10bxVlOeJyHSdsl5K03Kk4Gc1ThtN2Zpbbon7OS+IQ77
R8h+Oq1jvdxjlTc6PiQNRwulsWQr4LIu8JZBxrgwv8jWMVwpLNl97kLmZUVDxH1R
mVAd4b+eyOTRBa/DW2Eg/nBIVyUW4seATk3G/aJq4U+D5BfShrxYvNJ17oWbDUlW
5A9MVc7Vz45oa+RdXd4WR6Kw4iFt9Xvzmmy9155IWm3F/SViduGjgFkqRpWuGVnG
BEVFGpSpuQRGt+tT97uuJYhixZoaleO73Y7boV9JFRUa+YHGkTyXToGgiLCYgvXD
lqKZ3phnZvPkSdTFki6GOTi/imcE4Bm7+SRmpEeH5oRwDy5k7gW6L2jdhxqEcLO6
lcnVCrh3CFvpnzcdGMTIMHWi46xDSA5qHxQARDvBy+3EDBwF7yVz8MgAFhWVcvVL
vbfPNxByVmPhHmqE4tDC20GTr75ZBvqX7TEwrMa5/UPH8hYZZE6dFBsPAb4gNjP1
n4ecrTEU1eVei9AjJixh52Sgriv3m4p61cM5Nk4Tlff52B/v0bI25eExrO3I1O16
UuKC8LQhQIGKfVdi/3VciALxUG2OBUG9pQc0B89Hgy8Bs9LtV62up9k5zQtJguYb
6Q+ue1vXo4TOGa6obdx4KgyYsQpvgvuqCt27EpjSdGxOI/8bhjDZyX6anYKIEN++
NOMwpQbxSp44cWXhFi7fbQgIsgX72SzssPj1Z/NaZt+naMvOkLyw4mH7pqtNDuH8
eXS9n12TAb/9Ymq3FSOfmB9XCUly+1+brdClIJ14EHR66If5v/N+5zA3rTj2eyde
fByxZs6U0y301oJA89aoX5fo2iaXy7oU/1yNkux64WneeuTyd/hdV1/9cK//7Fdl
JbbkCkk2XruRiLKhSjPXoyEq/elp3+dG7tmlenS8XcKSZQjDuQ2VzvAJ9rpqmqJb
NVgfC7jqHkpIprofvUBvHpJxZzZMxn/H3Vq5lvZcfZ+vPjUk/Vml9aWvaIYCoAux
pBwJtaRg2qpFksqwV82PpUt9qB7ZfXme3C5TN8Q/+nbT37fYd69XdbClIt8apGY1
QbpPHksbWzdAoxLYjN59lOrvEML7Ev7VfXx2kPXMukCGEWzFwodrvlGhWl/DstRG
MM+kIUSXPAJisKPo8DWL0st85fBs81/neGHiLq0d6rDjUwkyh+ebUkRuliCSWsaq
b+lGsa0Xs4HEoX0a2zlJ0TrbfOEytA/+H/WxMeGxj3KrBu0RcVp+j7acc9kTgbYk
sKXZyV9DP278mD3//Dn4gI3SnVhc62Uu3Fs5vhxsvmq+PaS6Y2pHrIoYMo792l9h
DXZP5E2IOSvctWjl3DJz4eUcIyOwcqeSGtxOMIGwr/wlRzglg9Q54Z8mR0s6QfB+
OGwPVfG6P/3jylGBCOVfXskGZjKylP8jt08tDfQWSn61kjFEX9K008fYnDkZ0q1e
IRhnmBF2YOyOWl+jfXV8ojcH7u4GMSLa8AsyrlDy2g/k8x2wVSIfUHpaaWQwQnAi
8Ad/8hze+TuS9vH4J5i0vZz/GH7iPC7AeQjjRkzW6Kb7TBRXDJCkOgq3XJUviGVt
vwsw/Q4XuEGYQSkYtuo0PPUYsROzmxwlXc4VKsHvZCVBXbLIkySCx4bcSbjMFSdh
Uriz9LCT4aWDg0VBsAWEGLudpN2jSTZl0ACs1Yyd+W2wgx6MVkEoL5d40VkrT0B9
bGza/utNVmgUfFbGO4kHO50uoKWsJy9/sN0iy6KUVEFEQvIO6wuhqU7SNtZIl3Bj
H1SVPUQ4Veyfn8hqF5SxzP84taeNsXHpCfS92rRtq13SfyjNmPhMN8NQkpPn0bzB
5BTpAsJhfB9dBhjDl3N+c5AkkxiIor0JNqroJHRFqH9XFfT9YCcf6yyEniiSwMy9
H9pxaOOIZPda1ttSBYJGgtYyRnamTNUpEuTf77ARLtMbruMMkIIsZI3t5ukaCOPF
3MCtoBTv1cJPs5Bx9uS1C/JEFHS6TWfpdWAy1sLxm7ScWivsBZTHXqBfWitREvem
+UDT6/72aTeKl19kmMw7JEUABHmem4xFIu8QYbKLHvZyLAa2v8DWqfGQmvzISxV8
5SlVNdVqRl/LwoOo3JTQqhs8LQla0SwkAGnmnEjpHcuHNSmkYUlif7IWZrPm6faO
YssW8ub/0h4yaS0yZvSaiT90uNez1mqNAZpoOyu/CSf93vkNyuzLbbva3vdX1cmT
1sMdj8kIVGVR0/5mbuw0nFEnm/ACOtSMTB0H1uqWwtcg33RK+Z2QnHwKeQaQ0yxY
YM8VR2i8qorntphYqloo7ihf13qIgLmwZdmwI8RhgWprX28lEpwhRruXnAuVJM1r
qop15ddo3zncabVLE2MMZJhD4KSxzSdvpE4J9LV+0uszIa88mwEKAXpdAPJotlmx
NWw9UOFY8kl7Qm7mcvo94TvEOtoSjGnEJiqyhN2IDLvbzIGlTpVGkGaxylHFwXXw
Y2QLrYWyzt/YJLNANbPWb+eM8mFbUeM0B90n5DvJVMDsLdun+XmkLFEHNdaCzaZB
sG72G0/2LiTORAb79FNIB56nZS4w4vFmLBvbquEge8JcoHxQIS/QV9N5zYhHG0lz
O1tlUSSKPFFqiu2c+5JYMMy1fRBoyMiML0RrgbyX8yh0bO4K4/jYcNKTUrggwgm2
NlIzSOIpZXwKTErd4hUI7jIXzPO3GYVSVukgAbrwa7cn4za4gmoQAM1hzADz6Z+W
gcOl8aNZnF9aGRQd33pRJLVAzhZHDLvV3fiGoOypV9HuwKbbwS1OLeEtK3DyCoyl
4I6wkMFjOKS+rrdfwBOy8imx5fd+yMrUsnmkhM0bBDLKiW2RcZYBfXBU/7PDXXg0
8MiYVIce5ngwQhOXWecW+4TO/ZMaq5aFfPvkkfp8JEmu+DjaE5V97jy9LDPcko81
CIICW+AOsMWJlSvlg23PlXtB5H1MDEA8CHWHH02Ao+RIsOtEVK8mYvx3Q0TSgRpt
12o2OrE/N7eNLgC98bw/MrF2wc9Im+HTW8VIPYImZAT3YQw/y7sLGo019iJiY0aW
WjRnYVf9a+uw6+dQ9817zhKVzz3gIHosNds+K4OjuVbEMzWHBfIkRWwu+FCq62HG
UYed8NeeZl8AMKKgb8MqOBwzl0hPs0i/8L30+HHCW0MqnQ16isZJwBSboJpeYsvM
UBztF+Lbmh9lZUQozHsXF5MJdW9cp9t4GtzChIbevsd5QfOevwXuTzSRdAD2my3e
jDBlnWB2CR9RnEm0UX9ABv+RNMIjNQwidXG7vtU6SeDFFQ7zPPyGQlOz35J8RQ8H
BsO+Y7rrKuWlK3xWq5nus0+yCxXDalLYxno6vyGee/Uc+efovfdDNwArvDl0wrGu
ehRp8YuNXQcd5EX8/KbgUHR88I17YZwwKCDRsbd51Jv5qkIZkwbDXeOaaRmbTS5J
ad2kunJQd1KxYpZDhjjZuZW3Hjk38KpFjTnaGX/40ce6C81KUPmIZS2Te+snVaf1
zSxWEbWiys4yG+rANt/rMqft3c5TYdCiVsFXT6hmxFHmaHtQpQ3DjHB2BwRnpe8Z
Fo0gOt8hWLxQL9uKladu69/173AYkMEpaLJ+EvaWobH8NhXRhlh/HT8oo/bi2q0j
UwYSej+1uNgOuBfebr3x97QcpaIEBZaj7g3+iq8bHhStx4ou8YLeXTN5oxCCz9If
eZWvDT/G6AvotN93ifA2ywqPy2JYlUxGshbDcM1IbhTvBAColTauUqoaerGgdEVb
WS9lhY6oxeSbFbpmjstQlA53mNQeyJJ5KtxNQKDpeVHQpBh+QeCJmFZB+JMR8XSk
QMKbKqKj5DN3ikhBZ9lJTzdCVG8wibFJ8oQhv0HXJpKgf90IHubht5JcByk5kBSb
qiCWtmVSOQEdQh8zjaF5bYk5+WfG6UKpjn2EjDakblncAPtkUenXaNOyXSw3EeuW
HIFWVG7zMOZnbXQJxUoowahNZs3mKPq/5X3Tk7DYyPTv6kM5ac2NSodZrCf5+iBG
ATBRahB3OmOVQ262x0jYmagPUcZHYJI9zbnhVTYCGsN9EWPXDvCdCRUKh0YpsU2n
au3IEodrchdw4N805ehCMjGqXHPrRNxDkRajCjnSHTdfRd/XiQCDiAheAc8EP33R
5pMxE1Zs73XN6yqC9arqqFrMmG2D2mFntPt7tyy0Y3R0SEvsgtMvx/6Xlgj5t0em
j51L1/3jz14XfoqtO6TtqmjKVefefKsg3qRC4vm8M2cmQXH02sUn2PUleiTSPNG4
ZgZ8GM2i8X9d7eC1kML7f5HWhWtS2YjSTAWkVThQmCc0RJSLXo+zdMUIGi8+GDsq
Ja3DOzfEER20mp+KmcLZl9wjie8m9gdS3QUAJdCcmwcHE7YhTeVft7MNkTErXAw2
/9z52aACRbK8NTlWhwErChMAgC3vNEJTEyr1sOliJhZtKprXlIqYoqP2tPd0izzi
SbOsGZqCB8JfgW+B1ODzgodfpQs3VUw4yZRiLX9x0ZL1Ene+crOF20zKx/kWNEZE
39h7u8e+96b14QJgYuPCycc+pxGXF3LYvW4pshVLzWo3rz9iBzxYe9Cu0KU+gWUT
EmxtFCyQKPPOGSZH9lbRzJCxo8wbzww317UZlu0zT3iX1sgP/KirIMHVuO5KP+ei
KHsvOS67BOHgkkljCLzUB1RfFouBRs/XO8SD2z6icRitlKRx/2/pTmv6QQjknBfU
DzX7HLO3JccdPiV+u4CrlSYo1/kPA5qJu+GCR9SiPa1iwnyDLucgfo8CNj30quWz
69iRg6dNnrbNcKCJ+bLpnJmnVbYqMGgA7Ck7qpADpPIZpI8vKBmSgUD4KmzdYdtD
Ylk0iM6/UMTBB6OBUWCvzl1isZ7G0rxeEWvCbnrv55Ta0pW2tzEA+/rLw+Zdv6z5
LpBnyP7AKJK/8BKkM6bTo9HUl0q1QJfkyKugDEREiybli3t9uFhP240CdpDY7ukc
3IZdwmUUnfR3CpvRMeF+9B2UJ6B8ab+8Nt3O1NctJl+cMB5xG81BFKz5EncIUolz
b4VfxBwlM0wqG82xAtfwuEgIwmR9Dd2jXVBKC4/4eQqWtX1YxehCvmh84/ABTJ3m
QMq6zi3YNsmBKtxwgPIHPH3LUwbj6i2PR7UcbwnjySBpAxBXlB2QdJro9jr5ORxv
hv07g6/1Ou16oj613aAzZFS+XmbTGnO3r4aQXspzE8NErEap+7zvFC4FtJM+pJA/
x0lpJqYnp0gS7Cmysr5W7dlPL2drn7RkMbIJUQl5KhdZmEheD/WxsYxe0wXv5iFJ
LoTHoppNGoughTbJXCD2idNVFZ9f9o+naBiwl/uHLkY2bVKUjrEH5YjxmywXrN3m
SnmN1hmCXsokkGH/xk8vTISZB2o/5xW9Q9Pm5PGZ8rLP3wwLJikkvPvWwnyPJnhu
rYDJySBKq89C5FSBG+IyLS+Lz22S1nkq2vVjMDv9eP3WqFVBFwqQZZUkLWZYIQF9
U/d33YyCnfZ5pejoPNerBpeehUX9KECV0rMAZy0yrNE3adDnzycgu0QPNZHWva7x
T2PUXDYefdBCo5zecwwPlt5FnaBm7UHQ0cgc9Ktkc1xNSvkLMMIvzQkqWhhuwKDD
iB71cXj7g9YkLXr898SnsgS76qXfmv/1QrUzX0eHNKlO6Aj692gNIoO6jm+4o4Qc
Z/5XoV4/ToPlf68qLcsm6cJSUGQLV+FFDlfdMZr3XhsknF7psFoMNc9rt1lqobiU
QIr84zHwICh6xenv+faoyyXaPCrhZYpGEsJ7kdb754YIgZMzBnEyvuHjva8y5dBw
nwYhGDatOH98nvz2rPa4LNQs8KyzzE8hTJhj8qrEyccvmJ5xCKNk6vRFFT/XGAxI
vguc+XfrfAVSRX1IkTboLK+0+iuLU7VqmXbio1CtQU2shxn9K94+IvLkHxe21M6n
iW5UziUN6IOCfdvCXC1UZiH4aoeBCF6PHSUdEDJuSDKl0Q+jDlMfEHzH79XVhviZ
5F88Ppblv5xEXSqPxkp0KkhTaPc4GTW0sF50t1FJpE9ZofzydMLYnBPr6EM8tFmA
D0Ze2o9YC7W3vwbMMYQccYsw8QZNw2JkbC4EYRfP5logmjqU9PiJ6kSseXSO/dnm
WQv+FZbLAZbNqNsj3osRK0ThtFge9WdAquR/EDovpdnNWAGNfG5pj/nxQmia8una
aykbnlLlGZG+QCJcZ9Nv1TAhzOPYl8FzqzKinuerDy34XFp4scl5eONUfWr2wRuJ
RImF/KkbmDJy8p74qJwAr1yc3cDvOERMgAzZZ50qWDTJGukb+9T44hSjVG6B5fUe
qfbGMc4ZEiP8B5ndUn8EwDqNJvykfh01xi9TH74ocyiniXIB+T+AX8QIAI4DXNRh
cv2JSkyoQrxD5GKgZFkDANwW0N4UkVVCW7H4mZAdhAsNLVotB+YrMLUBhKXPGZtM
mM/LLvAtIvtUsfN0wYVOGlAt3ZpZpAA1FFAYQn1rA6QlBksBQWo0c5GppfzCGp9o
e0PjCweye7ewNac8QVgCN5FjK3enZl6eBNVG/KawQ6Ob7+GS5ucuZjfTEOIAS+hq
CbMp+DTHBphwH+5DXRfURMCoAx2d3g9zCRSaxOCPIlrk2hyc7Z7S4gUGaV58qItw
IjRGgO6KF83p9rj15Zg85IMqDw3dknyJewnhj7+pK5OkP0xgBIi8wCHnA/bmmeU3
v8IQ6FOW/xyqq8+6a0jfl1ClBAix3gVM5uskK+u7gLlIfc/g4WLRtcEmuhMhR0Y4
Gpc1xkHkyE6AfD47u5Sg0Aa4Re+vagsjBwm+XBoQrctnyiCLdYsvUGEKLXOYZEqn
0aYKB/wyGN3ALlZcfawhWvBG4z8+MH4X8FCqRf9WdaM/5Zmv/1HcDt0fpatgrtrv
sdpAA4Uq1MFAYlLN/eQOb9DAoMANOYN/K3nPM4xK/h5+TcG/MzM3JdfVwSWUSdBA
e9w/g0NikTXiLE/SY+AMTrxasRcJQZNCLv/udKm4EO+O1nL++GLcaN05mt1lB1En
g6EdW1WHEbw0VfoRykdNNLfdG6lEoMH6IbWwwTZy8XsZ4uuGlLVJRNA3M7+pWECa
B+1a1NfEC+ePIzbHRYSggPZDdgD1F2liht4liMXFofaeqlGS+Vw7qIT2H8w/z6Te
TO4XvjhZe4asLjG6Q2oUTLBwZCdc5N2cHklfE+Ey7/OoMxWOPz2rJU7gNz4xwCOI
W1qkpQsSwcm3r8X/rrwKjK98sTrtrmXleb/xKkrzeIIoqSYKhcbuJbZylG8ClNik
vVEreKAL8lIgsvTo1IIwUfsuUQvMtFHOLFWsFvRV0Qkn2LpPTTZ34OrL8182dc18
iPHqYALoBNQg2/ye/TWmAYYn2/35owLr3yk8wVPxMslM02OA+b+NIsCSuQs6AL1C
a20dQs2IZ6qk1nKATdg0cB50B8Er+GHtLgcjT9I75vz1UCoz9WvSyGxKjvIbllHD
5gLHC2PfL0XpolB1xbLNl2J7Stdzl/gbZs51lGfTUCbtfQreqEXM7e5xert8NEDz
W2xCJw+7n7B6FzYKd/XR2ducDAkKzIkBZYH9C3afN6jtfjyCoJ/SSpRWvN4/217O
mrBf37gPQmhrqNO2fb1BAPnfd6NgxdCybyTCKznDQ23M+JZGupHUQcROK8LYs5Y1
W5MkR+A6AWG6y7gtYA+d5rKigyuiwq8vBYA1p7f25DqXVR28jWSvo3ziprj27j5c
tpi2dbSWT3rcpwDznps9nZZe/bT8BIXL+bcGt0yiYdSIKJ3QGvPKhFK3kuL3Ywl/
zYt9XzcXcFi9DWKjtqg9wJp+Rr6wU0mY/TzPYYqbp+6QaOwzsV9l/q220CUUGXw/
dZ3RaNw1roteTvScgMjBA5lTlI9J101O993xkrtMCGnfIjMlUpMtAAPLHHK0jrRz
fdS7oGmBkDGYnNo8amEzwi9CpPzb8nKzKCbsmqZ6F6SibwUp6xLfOPXaoNdKYJG6
x3I3CiK6Fm52znimpnU1q/5rzuulb2MyDR5VpbrAZbYVv6mB17RAJLPE+fYPH4rR
cbBUz+RM0f1K6ZyZX69/v1oI80CHoD7a4DvDIG7y2xu4YoYPsHovm4k7hDJUq4pu
nmjaQeemo0UyHhijvuBUKE8EgaY1n/CaZ6vB4ldsLY08IL2A77M3bA6kccIzOKRZ
xsIXuRN00S83ROHvk4cFJfzE59Ok5mrYf+H4KtcrUU/XWjTGme7Lsc/Nl+D1SW8Z
OR8aQyYBwtLe6lHoCPz8IEMfNtb1w9oRtes093pKEtBFyJuMuPwG13AmBnClvzho
F3dPiszPUgvB/GKTGa9NU0PCkTnwnkVaYFeWc5EQWUbBdtPKmc3gyiTsH+5unqzJ
w4GES0CWXYifGoDTlivaATDHIHzhvqaRYne/z29kS6XrwNHI+Ym6vZ4pRLSfW2Hj
G+0FeQIRReLvHq2IcL1dHUt1kowDfh4AZFY4+nHe8UIWdc+aryt+GWSgnbRpviih
t8Y2BqCt2Kut3nrXhI6fPpp3GKokBCD3HXXFIj/OzAtsBaoti31ackzyBUwX/GDW
5MAQVL4BqxwZodqkKuiTJ+pCkS4g2b6ZXsmMrHMKVZaXej3G+bDBFkrE9Y4GqVgd
0qP6rVNnAwcyYruYVHLllWZgAnS6SAvifDTQyi1+C8aafbLjWlMCrKTVSBpMqke9
Ut3YK27BWK8CqYGvWASZxvDCyiIaglAWV2SKukjWzIRHa6oI3E19oYRx/6GhtWGx
6sMppDturgucxJ2b3M5+DaD0xxY9rVH4IhH23LUzsaZDhtdfAQoLmvMQbPCcfCa+
mlNIleOpvbn/MCYnyT6CJ/QfT+7Tw/B85aGrRAg5ceQkIbqTwnrmzfbb/6gIUaOQ
cLMZo9uiScRPJN4IcxFY2KZxMOmTpY+1F5oAczC6c0F9DfPxEydm/de1Tb/vT7O2
4FZ4kPjs7o/AW+sMomWWwGt2lmlGOrGRRqaHnXBiDEuEEtCFTw/v5Ti2WKMVHZJi
DTfWSegAhb24NN86C/zbOd7TPLGAkPXSI8KopE8V13fcO4xSg+ni2c3jWLpmc63K
C6C/yek2WVKuBSc8oOVt8L79K3Ru0yVh1rMrR0GRVAJBI28BwGrY6bsUZwRfbV5Z
ne/q16xfFWGT2XmTOUGFPoAzCidRzFJcWM9+f7OzAVWiI4BgVfyB4KQdbS1NbEOX
5Ky3ZWKqTdUm+QH6qTk2Ky3jln1Vinrly5uKwDfpFxv0axlrjfjixSP5+k8nrafz
1MXsbfoXiT37ghvMl4Gvl6UQ37L1LmcWXxPGgXALjlumFGQFSup6177pciI92cev
7vU/ISfsVvm/MtYskIHwVja2+keWxPxwqFtQB/8NFHqRphFY9Gf0YJeL00Gq+nF1
9r3OjoBZLAyk7z5JtggqvcfDnOjEu/6z5eqRbA5dHfc2jQGS8P/xnFZRiBjnYIQO
q3Tr5H5IGVrhZZZCu++kg/0fK0O1laOWT9cH3IEUiXwbcBSy8/4e0gvqnsfPkDug
KZwScq+3y9LaTmjmUUm6dhk3fVq2GVxrK1FoUlz5VF65H3XNbnp0IJ0q5Dkucgnc
9qV/2MgVDiA6IJQiVGtyVW7xsrO4ixtScpqksQ1wr59RJv3RlF0OZaLMGjmSmbQZ
HM4G1J79TQthTJDlrbgivv6T+8lQUBrip32xRLD3ghojBEV0oh+leWfv1xXUHDE3
AhISMOpRFXL1lgiMZeo5koUnLeDy5PnD2zjFNMStew5F/uuwOrfuYOXnxiorFPVC
hc9USkMrg8/DmxkqhBzgg1kYadQqwhDBg/4JzIru43aLFGN2zlgmYTKEEf4aZ7pL
z1ZOVqjhwopX0kb7LwbNoL1y197qNuJtxZ+j06eJBnmADigN46Nnw2QkauSSxdHB
Ie9QB9kehONeK3HBDgJllMjBZKMA/hZmU2FfGDqigWc3iL6dp/PAhUAVVi1JYTk1
TYJN8WOrLNGaTVwUE1or8e8QVYQSjkxN0wBqqFy1c5RykT7pr3RHpUsbLv06/WOb
U1WEarJOxQ44qWpjMu0MTZFNYZBXk63am8b8EzU5+nT4kpPEvLgbezffHsTb3WZy
G8yUqN4A1AOiY1EVx0bfEIbIWaSZU5bb94ZTVei+NKJ1/pnESvVuOMWmCzOMdK81
Ix3tuAPPXbMnaPviHCDDCONWx1QQhiPUMbdqkt0Kffsfd9+Z/aM4TS89SfvsbTzd
SjKDPuMPVjL+yoK3/NjBwiHBWLekjtcbXfjt3qj/i19hcIVjY7j2FGjFI7OiELjO
q6NHhPNs0TChhWlJblspmGaFUn1veQqCkr1jUrgt3sVATyHQAoSPB+T3sx01ya1K
5sttUuMarxUgkZuKb41NocvW7mwR55eXQaw4zevwn+cx+EAdkHOZaJ36O9ncSyhv
xfhhezF5lwQRc3qFfX9xobYssV86o6vmOQI37Mffa/51yOSmFZ8za4N7Pi/Ndn5g
yeIywMlyRo3HpxEC9FB+pV78FJE7e4dLtOmpDiU5er8ItKAeQJSHzg+vN+GLf9ko
U6myPTut8onUYY3/x2KYPM6tJUqdmhcKDMQzy1nAvLwVZBoAiW0mE+zps5YOcZ8S
TohN1fStXCRPnpWYas1rBQwMQLVN5XdQTN7CMMXPMf9TevRKr/LSphs7OFAmcFSx
aKHdRxSjqxvXR4fyAQ5J91GyKzaNMieJ84VATJHmc8czAsmIcATI2ZnhdWl0w0+6
x2z5owAY+dugVTZij2P+OcTsd2yuKtXS9Zmd+3OpVuvpaq/ryHJR0dOSMqiAJ09G
T3ZBh5wD2uE0eamxXLp+9zit423woP7i06YkCB3xTiUOnKJAknabJdOrLKVaSTZz
MjuR4VjNOC9qe7N53e/g4KO0J9GWIJXvU+KvkgzohOmGqMakEQn4F9UDQtqZpyub
EzHwmKjfrwoPfJmxLpz4CNZ2XFXRgQKnYD0ZLcSRFptC4Z3h/De8FtOcn50a7qaQ
wARtXboug2rtiKklpPH3bHS39z6a6sTcS5ykKJvl8ibs0zjLF0vcdcvmfHiJ3zXI
eXC+xeeZjLtYlrd6gEsT6BX6x64E77ZzefZ6oc0XAdlf4ONXtX0oISTXFqe5Tdnn
HMBhc5FrB/+SrXmRQXGCLB9ViNsYf2JEFiDSRDXMcZpf+C7AfVJW8UM70LM0sP1h
c4qp2OfcPMBIJBErbHfW0vrwIvkix6XlcYoh2zZ2oHG/Xp6KIfiKbhsCk2CW7G4s
5OrtJ+XGNjPk797LguS2Kp942QA6b8c6XCkl/kMT6/JavqP4DeCSF7B/1XHskhrK
NfmLeiMLSwHCd/EBwB6wHgYKmKX4TE48QWCJvCWBQuAci3HD0c1dPsAC9I+OpiMV
Dxouu3RwYO21g8rsto+Bbfde2bJzi+xg+YFumpxGSfaGB4tEP1s51fZ7ASYoA1mE
2tFInzMqnKSt46+6g1qy2O0BODpyJWviD4R86oLmtMeoLJmkKqchfhN1ss+3e1bP
cmIsQqSZ5WC25Jp7BxEzD/1E0wQdo+ILOFZagBoySjmRTXXcViwnZUIT7opEoRm9
Dv0V5bxKPnFr4qVz0qa7TuApTG7PKusqG7HObFmfqXnATLpoeen24ZqgBHek9kOV
2E2a/mW6/nveP67teMRKDkjn2Aij/nRPxMJLN1LKnl9fynY7ba3N/c7GsHiatJ94
1Y3y7vwgET/SjbN0YuKzA0BD5afFwpGnZElK74r3Yck/NWlh/sKU6/VyTPCMeQL4
ubl6Cl9RwWUwi5YnJ6NAnKlI4YpC78E1boE08Be/mdPkD+q4RTaGVUDOQPDocYx1
pvhzJTLFFu/I/n/WEvVk5QtedGzWRuc8TxegHBaM1AO2fuPMtvgjkOwUIVqkwvk5
mZY90wMIOva3dAeUuqxqJlWgII4htEXHHlNTILX5NOejMyOI/ew+0dh+sdc71Oq/
kcTPR0QvEC3e8XL4yZh0yBo9saIdoIW/D73kU8CuvhIjij6fGQZmxnN97BKt1Sq6
31CYJwlXdALcKgtUoCMNcMfjjHYUxjYFULi9KlSYHGnIpYgNY3pnxlqG1Z2GHUqo
zKRwfXQg3oR4oRcDBFkmK1ZbwoK0d/rJdBfEHFOHpas0RnAZrgWrh4DpK/WKMR3p
dm8FVVBZV8L9eSTGcJJUezZUDFnpZXmk0AYgeSdMM4NOe9i28RBsAiVT4tzLp9s1
4XUPs7DLzPvjUo9KztJEn7XNgtzCh/8t3c1KnmEOzOQRMJ8wjlahHSc5quvEfghA
3wGtZ+U9uCbf6kaZ8jK/NgYphtgsJFMTBuv2YIFb0pKDsQPWcFB7TjSCxb4ScUEM
K8eOG8ProAlA/YWHgAaIy3GkOE96+vdhhcjRv0fELQSfq8G2qM87GDmu2s0WeF3B
bTKOcduWBqsDvc0MaNV2pa63YmVLqm3i687JBVeZXR1jL0eeXmPq68r3eVnFHVCN
VE0Vbhq3nhL8/2l1Ybod7Uhje1rsyGB/IsJ52TYDnAQYDLtVFSH2mdNjcwuiFhMx
KFBCvHroFou0sKzecodVPlqwP80pV9ELjW+a9L8rRNBPRCBrTtX8GRRK1JJUJQ+t
UxGaYMZwNYxLDdpeSvrOtIGYg5hQaODhESGVSXy2itPQmpU/OUAEWtyQNalrQSz0
2r4A/XzQxgKJHTMVXQoUp/9iVu+nVZPmiWJBi5AU0tFw6NhSeuBvo4Ic2N9Yvtu1
TPNzL4BjasZmM9dS41V0P8KUOAFw4wQH+ijzjZQRi6fabDeMlte5H0ht7kucP3UQ
pwh5L3O8ielMMs51HVuMotTzgphhdDUK6YiRSDuNrfKYIcW5tUwElt5Gj7T1QPtq
CmX6OHWAavNnCcgvsf0xsCHM87T3V+GaN1DYilefCSal5zgrOwoU56aiYdqgfY39
xjO1xQRt9K34ILCJR6pO4Vx/fLYGPO01LG0iniWES4124q9qGysHYvl+ulqq76tc
TAUyECmXkYc62Gsg1KwOyAGi4n6fq+9S/a2qt0/iFqlCqXwCnp6HkYuvfhuI8a8B
EU+vMncMTIbLvtqpXc/5TUYAE2R2++GfaHv0WOBweCxmnIf5vbZyM+sgulEv1qS0
j9LncIhSb6Jz/awpCPmkZh26AQqoPaU+Fd3pSiJsohCLmn5GCYNVLB3DQsL5gPKP
qLkaB54fgmag1Hc592eujgkDPq4DqIHJciynjIBwWw24RBAV8ZAdM4awjCJtPgDu
91Dj9VP0dYZUJ/lXdhpvQB/NH+D4x3D6RxrqSMjwhwKjn/TvolwY/avQ6Abhx660
DWWYYWiRgJDEvC5l1VVPpqJW+vKvFuvMJ3dQzxNMz3Hv3lVSvHS26DWn2w/PQq4a
G29THssREno1W9y0FLmq+FRnj6/g8SlRt8LlnvuPPM9pzXWNZi5+j2Gx448XZNMI
MWAw48V/QPspAV159s6AY0yytczLi6aCa6f9Vcjm1ZMHB1CkvUbDUeNbY0El2z+I
pE891QEMMZXffUNOn32Ak+8GSRs9lMc6HordgaHof+pwtsQYKaRAqEDg8Fm2Omem
+DHxxD6bWb6Z+Af0mbiQG7atCK87Z2YFEKvlUtgsB+XwT6RyS+zwIHYm0Mizx5yO
AtMLAj4hyr5a+y1OIZUhZV/wZNVCFJMTOwSQWOS5jpZbdw5prW4znhYSgaP2kEFs
+wkGzNciHH8apJV0fWSy9q2o2XjExBhyK+8lZoEVtrCDdHqq/gZOalPrF2aiZEyk
BfUNWjDJhnTRLqzuQdit3kIkoEbpM8dc6YoWwx9rxRDM+TR8+5SJHoswU7A+Xrt8
OReqvUTcAygVow98YAWLHVm1GldrfidvGmbXwHHjrX6kkgm0AqHb8iClJrVmrrHQ
W06tPPtV0RnTSxeOg8DxG9XHaF9+2QC54YIfvMBJ/oRtMDOuBqjprHCkmEYAUN0I
/TABD9wZ77U3gCH8eralcwmPULzmURgSzk8rYPJjY8bAnSxPdKB9yg2ITZRJ6KC5
/lvWJO4e2+dwhFZ88Fmk8Uwm277EJrr/aWiaD7GQTUELXD9PdTT5Tpqsxue0bhfw
epxHuIT2c8AijrNrx4QOM5w+S0nn/xUePhqwqnfY/s23kplFGABZ6mAP+MuLdohJ
CQSq1uwGh+34Z+QuWQAXoJ0ec5LjTobMbInqpsq6hJfo/659jxa8xALIFvpYERyc
FexZjhGwIc7O5q0hzeauyni8XPQhVsguc4DHI+hmg5GQQL2sTCRSGPkZLw9OlF4/
nO2NsTp023d6EJdU2shyGSsjjXmsBgG3/guOk5vM5/ArVzF/HUGoo66Cd1h0ui6L
A1OgzLg7WxjhHGxP/TFLl02foelmmfDcckhl97XNe7wA6J/NaQkjgc01VlULgW1c
pgW/S3c+PBDDuxpt99mbvCK6Ft3EMGETkcfmFksUfqjgWccxr3TQNnZc/gmTCYAI
TMRqVLBHUu8jrznOzUh+2xVRuj9zh+6VCyTJy1a5kyqaNupcCu/8OXHfEIGtPtkA
3bcRS48o0XA+JEplNQIDM+tbFhYccx1pm6ofytxvUGwsQi+5OOQ8V0LJA206CGFG
qTcPeB6d7NfzDgndbvuocYx/ZmWBq/LMdy3h/cbag/10eaUqsTNnnDxTW9jEHCcV
lwg0fEk1OxGaK5HZmdewB9vx/8LOSpSvWSvnCdDomE78uVuGG5Rs3IskMm+ft2fQ
taIm/ti+Mr3CpzgTBu9fKlgSISvXUoRRh5yYKgxI61r2WkDPyEBPCtgMkrAQY2kC
DzhQfVw6czPSicm4bYpSqXtrACxWVyjQmLgMfbg73vht+0Ol8Fxw1vvtXN+irUvx
sbpXj/nzJuKFMBxEx6i6vZ16SdCclyUUAGmVcOi3kkoTa6xhq2H8XeSwbENTHy9A
dcD4QvgjVB5KuYCB6jQ7C7p/4Oj1JjdOvHZyprvYD1nQE9Te8MwudFUYZhtSU6g/
IPF46Oh9hv11odQ90T6f3Aj9y35vmv/CBxshg1523kGd5k2/mGMk3qCxD7tugJg3
4M9S3Kr98vALM/VBGbZaqTnxEiL1hu7xJI8NTDEL/h9W9v8XIbUTvKKHE7H3gAFg
84OKelkOFHkd7xMOJ7ZF2WcWCV9WDsfe4/cO9p4tpBHwR+gsO6+3wuWCz0MBtAHs
88KyAbUOxoEE5V+ERlwLG2gwCJUJYdx75ofdUlRQ0kdc/hRo9LhA9/hv9gQNApkr
u52xg0EBRaO6dqS0PrOXFlgNOyaxXFMAtj9hz0HQJR0h0MIO+L2/D3I9/FepTKXW
QNyj/g3BD+FaAMXwUoTswG+M2c8a76Qoj0Y/bF1YPeHmPtK605zstJwrb/9WSIwk
jX0bjrLx+Z1i+i+k7GrMluCq7pcOK3GomnttuH3qH3LgWqGPt9S2l0+swC1fGkm6
Gf3H531JKqG4BLwLweOkFcCEFp+KFp3LvxhxInupoB+4O+N/JfxzxoSkdEyYci1d
Zr9xuH9Wi7GQHwXf+f9d8rt5xX89/aJt/gNHj8pZW97L9xLO84lL4JOcSQkYiiZC
n1AgQe75IiE9VIeCekT0evyXHK/HhY96EWDU3kP5LRptmQ3ufOa9zjSYabiFiQMP
XuaCt8H6uth3QuZAOVGR1aLog7sXjLC7VTPx1TRDKTYapTz8TvQV/WhXSWRPzQeC
qkeJU4BVvUDO3CEnjdI7gWmJvTqnRk+QM2Y2gFSeqNUYe7CpDO8qiDzaJK0ATjbC
8Ser+3b0MMwggPYR9bsNzanNphfXA8bu8rRXNzwKDXW7xn9E+bT+VdHcXLpup6M2
W+J1vultFyM8bpGL0jlVFdrIR7Fco3rQUkaCx3hQYDhEp+/Tpd4Rpk4ZI1AO1EN/
bs8SXIqrqMxBaEBfflo15f5z0hJpA6Zwx7vKavls3m81anT+70DogIx5FgHmEFa/
5Hu16xUkIqMHnARZWMBezaXcwjdRfA2gnzHw3oXZfBhWHqxo+4+ZeEJW0h+of8X2
kYCpQnW9JICjiUJ+agfAcWmT+9LgEeomAsHWimjLDGZYOgu5/GC2aPZpWKHsR8x8
ntypznHkvF033yUTaNtEN5kSj6b5A+cJ/PYQp3P+30jsdpOmeFOc1fh3Ie/R/Ocl
XTpqMxGvLhNJz0TK9bZcZ7TbZ51rvRdF2tj1yC4u57I/X8vCIyCnNxMX1rriL0XF
JhCq+Nrz4V/DiWjQoyeHu4+ql9T1hAze1k6QUZQSjcz+5XDJiuk20zXuhfQix9lt
n+YvVerAilz56iuN37t4+vgpHg+x6IKZMqHNvIeu1VwnMN92OBHN2fggpNHxjBbr
65GcATda4cHG4Ip4UlOYC8OnkiI3qsOOlxjUIfrQkKtbzCA2OpIijcmdeFRddQY4
ynQbpo7CmVAqEE660Dr1FD0lf6MRilbZ0XJhEurUJ6cx50r+8LslWs1/fneKs0Oz
IZGlHS1RCi5B6xRKc+zaXPtB+McnqCUUnDRkji8N3f/y3rpEwblcTwM48N4TtDB2
LkdplVYmavJhUZ0s+8qS0FkXjQoeMW+j82q+nhK5Nne36ZCYYZFZiX59SF63ATfA
HO0BnERRc+xbSjrt6rwJMKN++IN9HfQNK/fuTL5vdW4YvUInxHQr6jaLlGyZlTIs
FGurIIPPCNJd/0WFXlvtWjwE9fRkP0KiFYxN+MMJDgnrMb5wnDAJYl1CwedhJjng
Q3KZKnr1MhTwwkd0KgewOyusx3nC/2DcAd97058ImolZRtwwwGMMp7yA7+ocP11I
YqLNxrb82BOavGXVwkyKhmX7GOd0Bu7kNc/KSCXYA+hGmRt1LbxlaNF/8YlzbKxX
NwCNKwprqz+3MG2lZixIKLzqyXi/wn7D+sjln+P0UaqO9noUzDyb1kP8mtrttbFF
9sm7pdE2hCe9s1Xz+hbOePiricX1uGFao1btI1LPEF7Uu69OMe5JYoQVahIAc+BO
3o+mvxXfAcFvlK0yittuDYnueNAmzNbDoWLifl2IOPzJ9XlLOoXmmw7QKDnJBztl
rLtKBjtUR0hYA7jLap5QzF4GZweJqdw5P7vK3cLHihOt/RX1oWTiBlFmrSj4PupT
XUReDETHFTQeQuVT4ii/kqiaUHur4KDIphPfKQVLDmMvIYd+Cy/RiSKu3T1eTYj/
M9a853rNYfnIxGy8IOGd6sjDiEP5Lqa3EEEWJ0YdvDCY/NQpdd76fiHVtpMzw02m
TXOd2XHHxVslqiHt1opeoUKYNjBnoIWn8+16c0kb69kVNGY2OqMiXd8758Zr/pjy
usvNFJ9ZyehXZcRnuJl09ltHsXcEPJ2FCtg8YCZFbbKfYLNMDmhdcsNrtAJwKzWR
4Pe+VS2yakyRg0m20ufnrOxz367HQlyr/tRL6nSUEWvYyWs6uu1A/xudUvH1+M0d
75IefsWbcnVlif2EsV+anACHkX+Ao5TBCGraC68DEW3Q3EdPis6xa2tmsOR1ypT5
V8IwAa0thIYwbsa07v46UK0WE2T1tko8S7E1K5mYtjFfSMH6NoUQjZKEhFxKvEqD
4exSh9sM9Aihh0K8mTpDVvxQsqQUMDFwCFgPtnJIwI03Tn6PNK0ai24CGzg5Uxxc
3JP59WY3q39X/QtOI+dx6msMKU3CTjZR9hyfXXo/pw2cp5Fpczoz+7TjuuotdkCk
/XmKd+yTsQWytG3zq9snoIPejcXSU/y26CG9xyR4daUQyTiYSpbKKOSbNLQjmi1P
jlGkMX/9HIP75mj0fKtPSKA980PZJf9YCi2BeRkY6UCRrA5bG2X1o4VTHtDwSD1d
2J5maP9qhoAwJlPfNrn+WKOYakuo5Y/D1wxokQxU6mH/7If86UWhCeH+n2Ob7THP
kjsQk/KaHCk/F3uYLwn26/j0i2GMXgMwoi5V/0csgZPkkXlIZCXxCesbPVcz7Zmi
x9U8xzvoccuInpqFoSCowCmAiVI5myf9vmHGjW/QVyOKLjUyHMqbhB56BRznLsTm
LZ2WICqYj8TMGWenoL1NRDZPlWZgj2lUH3vcGtdbyO9jUsaImmhkOXiDi+MTDuSm
DnJh788i6F4eNjQ4k89gAafFn9AqzQ5cM0YJgwi6Xn5xFtiKl0AVDnrt1ocM9Taf
EJmh8QSYAfhz9nUSc8Pvy7AQQEJMle6qRs9EJdWN1xMqtduqGFs/+VHvpX7NIRB9
2p+hPmKLR9K0o4cskTJlcrPzCqArnIOpaVQ/Kk/NCT1X+h2Q0t31cbPYhZvJIAU/
6ALHyZaKZcYzmIQ/Gc0kl9sUHzhT0tiJhj0S3o8xVYCjHMaBvJFitQrEaEFKq92n
SohwkUo6UQC1bQRc4HS7ZaLxFw4VdBy4dVt9EZKaTW497jbmJ2HYIk9xnFca5WhQ
aTk+KXexZ2xsQo9sqWM0BwheNl9xLAVHmIUXD9izHvOkSkOWQv8aQ5RkjFjnm9/i
Q8ZEvanJKsCWhE5RgF7q1zM6PEjTLRUfVYcAuR17GrUYVYKqH7NfFOAgOctLoycv
tpSA460gDh3xEGjgjv1Sbu4SB0uDeZcfZJfSmHfbAKTS69NQseOTz88xdpgUj7NZ
7C+PH5eX9VQhYih4PdhiHOj60dBsx3FRzudsrWuRalbGUNwE6kngy80y7oX6eWvh
2r7T8rEghGk1DRPwIVgxFq6fK3dexj0QnZjb89uQtQGBKQkYuYFdHfWs8y81cC3f
4sO0tJzTTX8n740296GFTOfSUODVTEHYpYPtF3ZnkqU1BjbKAZK2g0I+l6Qqiuj2
IVzsUaH/K2c7U8h5RDV6qPNfGs1ONqdYrrjWo6nF3Pjb1NPEdpIgJwxuUUWgg5RH
uci7eNgPX3Mj3Hk9qU/uIgVKOYu//AnAChxRuFQG+ZLifAlkcaG50XzUQ/f35uTn
u37KejU8TpZSLFCYXVohP05fxUsGNHbuRFHpjcfZnfEZ5sQI7I2CqRSdA6DqzbVV
ldfDT3CNgOcl96wSK6PRX/ApAh1oIF/cAdNqsFggJYNONu6Dmylbeev0+ZE71Daa
wEjFUoZyZwh1kZhVar+cVE24hEBTYJ33/NgzC05U6PNBfEhn26z8ZZpkbwDLofsF
sZBELug+kTqNsJeuPFJoK8M6l3Gv/cZMi3XZAnEFhIK3KWkpGg4l/ObKnUr3qpr+
+bBsx9+90h1fCi3cCefIksZAWp9RIcbQ0OsZ7+7zp+29e/DB03ouuyANO5I7ucvk
rICPScWlUduTCBdjv5razw0PzQ60ByHFfPT5r0215QESgoj4z+yzWcMzQsoQshtp
/vlHSpxSIr9i+Lt2zWKFpQvLf6ccXKI/3qmtE2kXkGCsxsDGFN23NSuDi5MUpSWg
1UBCFyD624iNFI+bdMmI88yvuL4n69tryb7HrgvNIEh5iP0dxPCMFDsGB/RBA837
6cJYfwScyCTgjAP1VpkxKBOwiSSK6oMDEbDckuWCO7WNv4TJg50ncp2PStrheJIk
+tvawcZI+HMjMS9ElsuyCHcJdSU9Sicf/5JvKkSU0D3jKUh9paPpgCn4n9XQ5j9x
dEwhxIsF7bk85bmjYwp+MoIQhY3YSasvwXMbhrkT+9Mc87Pkp3zZLH9ES7yiWQjF
LSqKH4e1ABovAwTmXcw/z2O5qAQhomlaLPJ6YjymaSnPRvdDKY/U+jZ7IQ7WxzlW
x28/nGy9/w1jYdLXen+vByqnA6zYvckALfhD4OyDYLwjQnrEeILkJ6bXXV4aBBiJ
N5uVv2dmhW+hMO+l2fBUGswHV/GToutTTt8Uzpda79gqaCqCICUHWvTwUx1yyhzK
CHcJBjoSwyful3GqPyq9CQRuxa23VyGBcO9WP+V/LGc8BXWfS6/h9QhUlqs/yOr0
VfTRDB5bAi6cqZJA9DCyCSZohCLRqaOQvdg4SZwqa6yfgV4XphY5zdBxxqQPttmV
/2gTLhrswcY0C9xXTw+XoxdM1My36Sglnb7LI38tdwCYs/lTogZygSu02Efjq1bR
rclNNp/jsvTnSxG44p5qyQnAKbCtS2DDJQZewR0PeASHoWwVW3PtujVt/p7vJyqr
2b8rKU3jCkePcWjlyoSRglxzJ/YdbO34OA2lHtVuCoIaW9E7Nx1e4wkFiMJOAa/9
8fLlEYSfPFkvZ9bp7JMCJtiNOAhMDMcvbRjgAld+80fZ6dBg4v77om+S2EmkMXKp
YYli0QNGC5osYHOR1kBxnObyAzGWcBkHzKclesHYTxnncLXEUDV7GI/QFFlwkY6T
QYykltrIl0I3kiobWGZikqwdyRv/+68ai/gSkui5Csz0xBm4/2Mp0Z/HRheErN8+
VgyOkP1r/zyCLKWeJEquFEAsecT1E6gEBpRaFzYi4ifH3T8vWFAARvTWqRP3RtGi
kaKclw5xNFf2qZTFR8iKVum0b3KkwQRe6q0nJzxo/pm3Jnck/x61qTEuJ9AP+5HB
l240CZkzb6c8BhDc/XqITSOMkS6nHerAsP3Aw5n696+GkNMKsHMjoSU///b2gkhD
xo9Xkqev1WNSqL1oEMK3C/u7paxIfCRqR8uC9qq3LaN2tOibTvgsLG80tq7Mdtrc
9tEPx/HbUVLYLcZiHJYGVTYSZ49MQiutVulUFpQE6nJUiTeoLul6/cPW6rvPCVwG
XuO5reQCBMn29EmG2b+whAiXZzNKESyFA1Twr1h8pgGIdqUVqiur4Ioq0UcH/5oU
Es0fMvBFsv6uPp5QEH8GvyYg60FpAyo9EXWQrfTUtbVLiXZAWl1oIoQt7LgzRqQg
uSQQosMZORQZ3JJOcdjmy2r3f52TxdsP5kjQiGuCkJ1ewydi2EwkSsE6pibxIeso
q2hQHDi9ZDcIKuA5JOG0+Vf6du0HANIHKbHEUeZTXW7OGX/kaUYvqkl7sYx8DuJ/
T0k2bG0KPiiAKiSSfKQeQMe3IbhEBx0GQylPNlu1wo539VH3lAjRlDrQyfXM4Y6t
8CfkFqhq97bHvcKSzZQ6lMrAADmzA0oV+ZU/JANuimjj7NSIeyNccPDjTwMTp27G
16lLKMEKCaujTZGRqyZOlGfaLQPxZQjP/AF5rI9TppOKA/aQ7tM2GlwG4k96+kyA
M8RSwVrDI05IcY1K9H9gnaZYklg3aRsvI+hsomvHapSe8GWltmrLXkKVPzxLf3iU
Vm90pHckvFtWbUXfYRT85bulYVMSB21VSdM0D8UOmtGrG7rD9o9W/hYZ7wQAyBza
NKX6o9Tj1WTrlIZJ4AO1yXcoXWTl01vVzP9ukxWPk47BDTltzvBKDLQYT0uL3c9y
BOvPs1TGuvLR5fiEQUWfKtEF2lIQE9bNnGxAn2N7qcr9PSNBIQzh21ORjKhvdzOF
KTTATLp4yqQSaxs7p9wJNc9I7dATLwBP9MCw/Yj95hkL736EWXN9RSgQvEvpea2U
aEeOJAKQVPS5obmx5/gP113S09FAPrBXHa3N31efIoX3a3VsbP9V9SMUiunnfq4N
2YJfKlDoeQ+y/xND8SHiQ6ZusQUOLh5rn+kxLdsLGHKIIb47XhhPZzfMEwGbsKDK
S36fgnrxxbBYZYi0u6264+BXpnzr+QizXFaAUea3i1uMK3o6p2PSJ2Z7m518cBCI
t1JJ5DwI8wwySNYAjEuoAvVI0X9T2hfhY+q0I6d3SV2nGlIvyaS9JKZEzabWFmvp
zWP3QOiUbGhojR73Ga6BUSibSCu6I069lmYnu+6H2Cpm+HFmd7LIK/ogwvP0KXXz
tw2P+S9weqAjVk48lH5WTM/fDiqqRFltePuLWIHGmbjM4vy6/Q36pbYe3g9GgzdO
RQmMOCajJMkjWaqEjc2HOnNEOXsSq4uw1EWxvBxOL6T82YsONPgJ+0yxxMg4h2RE
OXnHPdMsCEpkwjbFPSzosopizrR7iwiMB9+YHmGwFus/qS9zVCMJf6JAfoU/ussV
VVtCY8tVW/lx34tXhNkEIPYyAwd2GI20yZbuw5EchyYDjqC9biuxHNtItU6hsRd9
sAOUHPDLQ0Ia6dm9XMTdeioiQUeSxMpZjCgq9Rre/JCaTqprkVz15EzwP94bD2Hi
Ga1r35bHZ1/bfZBjJvTSdQuqRpgrIKq87VGYnYy3S0m+6W8nohBIhpH8vhlM+Kl/
CFg11jBHenDxAXzDLJg56T2+uF+CplZ4drPabSiGLQ3CB06gkY/t8zqUxEA1963Y
C44BWa1RwxBzgfcBYOr5ZSNlNGgkMEjADj0v3Qmz4kwO6U0+hlyxhfd3AZeHZPHn
ltqM/gQjLkIbegSXF+V+7QCZLzVq/+mefQ2AtlifcWT546IoY57KDmdXzoxuOFAi
lwgnAG9k2OBjMKoZ0S6EhmFM8ybg5ANcg+6Ssl2/WczirdryE+8l1vjxze7y8Mpl
17KaQV2iw6ykEoHkdJxUVRp3YVozIVmHLzKeCzTZ1D+aBM5Q+yPLjrndtd1wxm2/
eledhqVbQHyDlTmFB0IGislrKFm8feV/VE+ll8dxBDrDz+hAxjzkI8OiSl0RUEd7
p05C8D1bke7KTlMSDpiBRLLeM0PEHFjPAF30HnKyFwKcSW4n8V16hOcRygS6yoED
Ugh1mttzITnwpbdGUofRCxelr4rLMgew2GYFGHMyd6ipPlx8HTZAWj4MvlymFt/K
/b3HRQ1iTESLWVSTdRh01vshfUSta+F+lfvUHHx4jo4bjCiJV008bOM/Oy6FoqwJ
ksy7lzQ9516ZgQg+nJnDTXe/u7bpsZazyd2N4zVuW8V9F+A06PDj+J6uj6d3I6sT
g/w2sdFuhkhIJkqf2GxWN5KV/cqZc+FSy+TFDPQupKmJteKsia3H3EUkE6ENl4cy
OiGF6q2ykCFssekAAf8/WYuZ8kOb5prqfsWRsbDXVBbaDxzsW7j6BAXOVxW7hhCR
sy+HNH51r72Cyh1cr92dnLEX8yWfAntQaC+AnHlkISRqJWOFWcS206iEZZRkpSbq
mYOLh4rpVHlemrlD3xXHEiMCVLKiDi0a22e20dhVqSqgbBpH3+ElYXo8RwI6Ci6q
lYJmhzSdmkKFV+ATaIHZExjQClExbwVbmuHdVqvW2pQDfG2RPfkDO37wskoT9q0F
14FNnr1y9gr3X1JpKzvcZbBMebXU1GYB9hXwhLgeUOkA0GPOqHpmvlESapsLJZms
doruTYbTgiTjCcRhWAr89Vy8dlpmaAyoh+qTJdfjxF2Hm69CQRVVAPyGZWVtWDkG
HSJwodgE4awULIVhk7lY53bm0agcwvOsK+eV0mMU7Z2M8mSbQ3dkp2bcI46guuQW
svlt7gqHfSD/eCd4LVNxfiEhL5njHinOjIrKcmlewL1zEh+hilVcBJyjjkMMaJZ1
rogcy1iQtpm/CrA0jKP7rBeI8DjDatphydcvkWWXY5RBeKQ23Qncs56+h30abdni
itL5gyqsakn6dPljlEV6N6iI4cUn4E8EkSnulK08WdL6G9zOH+OTObTfo0NgDOwz
yhYWJJZ4sHypPLfaoFcbRCOJuFWUlQ7qlu6+iht7dw4BXjGKJb3Xv/9NBN5O9kTv
fIGS4WACtxfLmxzbVgRfRuOhp9W7OyaSrU8WUatf+8i98Le3LSWPt3TiVTq9IrpG
KpjIXd+WrBsdDuC4KuaJw4aYsvVoRZPxzmizjrUx9PoGTAbv30dSZkx3916iMDg1
eQxpVxn156VXygCkh2ORA8n4/8Nh3ZD9o8K6nfNaXB25ZkA0XTO0EzmkYEgSji6z
diuAEdnHXC68ZjYLMLO0vLFsT1KBTnbS9hGqo1hXJIQ0vqAGTfIinnUqPaj7Dw3j
rL2YrvnHv30Wvm8iLgQs1mb7S9sOpUP/4QZlOYMQXn9/OgLpTTUD+75gfyPL4IV8
BPxAv9rst+jCHIoJ2jh8RiLnuQMzdvCYnffhPDYcAGNMuEJjkdcfzbduCFjcOhlb
fKy6gcH3pUBuk61WL6hlm9FWUWZ9zpu1Wry0JWfIFROe8//FaxhiJANqXgWR/cOx
7tLVNyE/0RTDo8Kn1elVDtiO+IK4Nu0pBFGIBQNhXBWozWkZB3u8ezO5KDOVaycY
sUCjRGPu0d5cw6kHf7JC56DPGulSg0aBYlPJYw+NltBCFSSaKgW6sr2Kejoy1QWZ
smytwk07g9vCEx8RgwRbG8GXf1vD893gQnsxMMFj1M3KCwj82IzucDF3MileVm+P
LYgt+GdXfb2nYoEiX4H7apocmowzR8epP57sIMXgzNZiTP8mYU9nGqX8onRHmPo5
UmqEWARnrJIKMd1XRMTJek+uSnn0AVqmKTfhivzy4OOLXRTbCdP5Wsu3VQH1suQN
obF3Kk17X5GrQvCb3EAs+u4w2AIrzt6IWXtRVUF4XZOBCSPrlFvVPca1hvzKNCKp
HCmHH9Y1QWGG8Rd0c/40iCxStE2nciF4Cm8ukmL0QqzYL20UsVBNZHHIU8ktOrnr
MxZS0QQSAfARhSA+ZI2y8e4dWS7jiYXI7tLUt2T/+nuNmsEgdlzyuq8LbB0n9dMg
lsOv42R0I4k1suzxXV89BryP3jcuQEKG8saMIsw3okAhNsNoI8K4OoSuubZgEsop
aWudH5tn3Yk9rX5DUFem8vtSk3Y09Cc2BZvalBWMOSoY1iyAz9zxkQmYh7yTzjQ2
O0rGrqcoUdMc5UzPibc//ZQ6/NnKbhQ6AARfbH2lUWdxpN82Z2OK6CwNAxrmH8gE
Wp+Z4CKFFgRfhBp7HE0e4r+jG0mtuqelF7Ghw0arjiNIPABmhgwrltWAIQ68xUoc
eTFM7v0bkO/9RfLs/u1ls09Q0eof6evvbDBmbKBYVoAnk3zlDOHD0XoabXPCvWV0
RriRMTY/GfZULcWF5C34cfit7vEwtejgDp1IVO/OH6E7ed4yKwyxtmzegqjsUTHj
suP29jI+gqsRn/RZGlEMY06W05yelbnglRT74S25cuZPBpBVKYmKh/pYAxH/nSFW
5tFtpDkawAuzsw1al+EtYiPQUlZOKN52FTZRObQ3Xe52rJJstSvsxZaxxUZNw2st
dB2H8AySMJQLy6bjR2SIJ6STB6TSsvzbWneUOiommhvVqJXLFLqo7d9j3HIVmn+G
T1K1oKxjq4Ek9F/nXROnw+HEdWyOewYPHi6NnCxn2XCJLmvEmGbvtzdObGpzk2EM
gabBobAvqP21D1J3gbSjWaHwXrRV2QUNuXSFnzAzT0/yS9zBKNwIjHCZPKGMf1vV
TIjLjTktYxxnlyE0oMqsjHNvBTZqduxdUlZhy3nBOOzY/TjgQbK2zUZiYerF4Vx6
xduKQ/hL1TdpaBhi+E05oQAskpx0awVUJtNMyva2w0sy3LUu+195oQttboPcLY+5
odNPI0lOmSyYfaPDSRIAeeMKV3GUBGr9nJOqddUMX+IF9Lz9tkYcD+V3VxiTmtqG
qaO30gPFy2d5M3oYna5hnAogpUy9JOWDO7uPv78z8Cpllsao57d5K4GOXBD6f15M
NYc26pSXtjcpZZ71HXd/k4eObLCGo3zKkFefFydIrP6miSzj1AuR1TW/ehIsFJz3
BiX01vvFAbc+5Axafzt6iVrLyucluUsvF6ULzADyqhDOs/RI16k++vPEJW6tDKDG
AB+V6nbW3BD1AG+ev+0ImfHAhPX8Fog/6V0PGqrrtig+EpzFF2uRmrrdYf9KCoVY
KoNwvY50JCLj11ceI9NTdnLAj/Ha73QGm+KUKjh5qSCffbmrZkXheaWVHS/06nxB
H+VLROAaBfqw3mB9T0918A2NAGXax3RniFe+bWLtrglDQXjU6PXZ7NAGYDDlaAzL
xZod8in3Q5QKVEILCPfp13uQm0lUFOQK/g/0JECuOuSMZnu+5ucK43diELlYA2Cd
Cu3iKO/nNCk0dSReuHd7VjoLFIBNqC2XVguiPIx4VjsiWP1wwP+cNCbDgbXGy2j3
fiQbAB3j2pRxWYQkOudHjdq2N9uinGMl4cuWjtmiKsI9Q5yPc3Q6Uuch1VajDBVF
B0+aYU9AzX4hWhndtuSvMVxDcssxcLsk+6yDlm9DKxYDTgOJ9O7bWov9WFLHHiws
FLXuVHm3B3taBcJcGtETwjclZfe3JHRZYe17lOTU04r8KKzZWiALNifqoka+InHK
R+jgBpXM+97K98+803CK5Lu0L8V43aBU4aLT7WSeifg5bbgu6yckq/De4OtYeOVr
0K2zvnBIwbeXx/ziCm2YhRpPvXN7Xi9RSjOlBMd/WYudLsSKy8oORgv06MuFhDk7
H4vLBEBHZiyb3HMf7wTQK6AEbfFgpaegjDnZZAofNSa09IuTx1auWakvj0FiB9ti
Xbo5WosDftsarck65T/wWPtczvNBjFInsczdE5dseb4QOXcpTHJW7duTP06/v7E0
JWtrLCXkbRI3Tf0gN3sIwweo1xdLVTAdCHrJVshUXdJVkfPh/VeHFJCft4Inh7Te
U1wkY/0IEDqZyCeESVolog7k9ZnwrDVFyA0CfJpC/Hz1n9lXhguilSGU+oGhGe/4
uYG7/OwjLzbMVTGM1QTB5ujR00Ce5hV8dYbK9OSzpICUEyMvQxBVBqBF8cIZwtZA
TH2UUi2GsAy4q412kcY5vKTuENHsVfy0jyZkeD2T8SQqRgKE1GZlT4et4rOi++SS
0zXFs178/UtlngJ236lvvoPtf+WAcTYdiG4T94p9rxW/EOyG6a2N0y2iNVRaHjAD
+MzjKBUkRIL0c4clkKt9aHBuPSUSjI3FZRmdRE79pJzp8Yy0w1FKQ1msjAEml3Wn
AHqJOV/HkfHfqR0wGErJAViCpSRBnd/xohMLvzBrI2AIWTWw9NDXjgJv9jRUdYds
GRRyn0tLr0t05NUeJkVPkK8iz1r1Pe9osUxnyoWbyR3QASDA50dyPPZCk5643i6y
E4XG+KpDI25BuIzzQgZFknbw9y/H4qRmQO3Uz3Jt4uAGk9aU9Rb70rHF0e9hZ0jY
Ujpbxm2VDRfOQW4D5kLlqhOlSqTLZ46ZK8NtjjtJH9Knkuo/MrUMAZWyZcZx3twT
CQc9l5rJYTvNlaiUOiKMPfBAMmKGmW3KhTLqH5/IpG0A9JetI84qsLlenbr55uD5
lE/JCRdltasp5v24SH8coIrFHko3IBAviVYzdx3flF/U/plsOK1mUgpPRYs5uAjk
3K7XHmxGToWkiIHjShrkLc4G2MvvNqt7zjN+NHOlAq2t6FWpflPfYjxa54GpD3g0
xUcPdwqhQjCoNUX+1YTEp1Ymcz05rvfrEK+Jx2btLgeeFcglTZPeyx+y/yaI6agb
TEvTyaElKozbFc8OmQ8m1W6gp/C5sMY4cYnOg8dVVxPhzKF8CsaFX94SuYUt9D9L
Ar7n4NmC3MxZ4QROYzAUUjMDfgKQDDJOD3GeCUHp69qzaDOwSZ5UVur3r7XdnOVk
AvVBHxHagEbW/vuR5Kt8fyVStJ+orw6LF8ar/TmupE+89RegiYvbD5hHnlqwCSN4
leYFR2lyvtZgp3C3z1C3DMrAaeYoTwjvq6A68bQKL6bUs2UjWXjoHX7sW3tdNEZm
8i+zhd8wNO9UAc8xPmtmLfeJQPF02BUBjH+WIAeL5B0sOf4mUscCyxxtDfYS9im/
4qWv8R4YOFt8QyZiD86OzO3UEEfwg9c8kJxyjPxHXE0oJgMFJvKnaaF1jN0t0n6q
q/egeV4VdjtyNjPwWSubcgzH13p/Zgr02b9RszFueGywuvheo4iN52ol61iH6ZFO
ghlObKdGR7TEiHxyR2icSWrg+qHqIgJAYB5FL17TQzMoKL9DQbp1QKLYa04S2b6v
uEW74W4nqS4pyztmq0XJ52khkhgiG/Wsig5tsGWNGxg7z0x3rVsR/EPy6yvoTz6v
Q9GdE4b8BpmtjrPZ7J9b5lXQyvDUJow1+jlbEg321r4ksqnWHXRzh+wOvXayxU66
pD9DK6k63i7uEksm+4eDnGSM4La1CuJGCnSCQ7P2KqVIdSdWzBlOssLLFXIEE248
ZWYAgl5tIVmnntNetBgd7o1mxaUihNjQDmBBqIjuMk5Lgdzge9V3884AlZPS5aFa
8pYQQlNwmJ9wIU6WKioqRmapToE7k1DPu015zgplTEFCBui9+KYIqBqj3M3rUysl
0Li6M8fS5NmH/vWrvA9ZKeKb/BYiGAHS9d9YAFELsymJkvlfGv5Ma1yEBWxa3vzz
ZpDwrhKBb2oaLcLJXpydlZ+o5K0fXO7LyKM6P7Gec+WjQv+HH0YErh69SKfbHuGD
bgp5/2+X55thq44hB8mwTV2aHUXaN6xf1NUzbV+XS4LqlmveYFfyhCmoBS1BFiPz
2E96cNMlP9jqVLxBu9nS5bfyagewrZH1f55HFbILLDzfncdVQHhNvQZ6Mc2vVm/g
C71TIWhpbi8+HvCR82aN0EJmNPlW0nKWfPlpNQy6eWpYLDdeCUi9zxo7IbUj6UF8
zAswH72iHkS1fuEYVByVdjRVm8kNm2GnziK5e1/QJ51IHGqU0uYZmsXNR0zxatmw
iYwchHKvlPGvY9rgUdrj3MWTZig5KVGv5+rxWVwoc9iOK36+2d8o4IWJ1brKeK5z
+/YdjGMLymtshyqnejinoWwxg2yKyaZMYwf3rJjKx8je6SIEOD7SmN7SwvjyO2fE
oXgBS3AA2IZF0ImzwY7sEvJZe0QLSSaG9x0Kah0y4wRASm18pzgowNgYOJ7TybRy
SCoxlKY0lv/W5paroKJDtwwifzk7JDHJFvhynU3UmBNfkv5OgIIgYAN4QuLaz7/1
yLOUaJiM/HDFYU30gS8AWz75gWJYCCw/kq5QAoqzHC/AO1U2ymW7d7SRKKcJT7Og
bOsXEeCy/8uK1DJ0H7vpYMF0sOd8q4FoaWxBHwQ/3wnczjLgJdzgsXXjquD+niUH
zBb0+8sC8N14tSSEAl+ZXw+MNies+MxZZDwuhh/iSV2vtPZuxVo9u248TO+FTzhE
wx8E5QkM814K1WoVz6oLjjS/ULiANl8ytnHAQ3d/oElPhyMO4v4DcMsH37Lu7yr7
eITLfpLD6BDyLrdvkpDNrmp9t9kuTx7VZaMvt7iIIdxK7cDPfDJSuNJfBy2w4cL3
buVTReEOZEFGbjHl+2xePt2JNncfPD9XzGTwJQFLgjWgat/WyeHO+FPTzf7Kwo9Q
/8/dC4qydpmBxzkZD8Jc1Rr92FAT3Az3NkSnO4lkX7lGporCmTqdFGhJp9rW0JLW
tDrtA/96EnleuN5Ip8aULFRv1bwlgo+Wu4j1UI6VxD/pOdjBL0fhet1EMyATYiM2
Oq/NpPQcUd1Isb8uBZe2z2LVY13MH+9jZTZBd5Xwyhr+4BHSGDbP/IyHPqc5xZiW
LwCYKX3M86wcoBctZqDrkjT8epp5bLU+QfG4z1Fg/H5ap8RlgQ8nj6MFVD0PmB/C
euVZREmxNPMEHxw6vZyT4X1iDTpDDgEmTbjq1UdrHbQWmBMOXgVgUWYi+NgnAFfc
nl9ltWMJqH9NcQrzAfq/BqmZ0XTJj+KkE8zR2EVzM/t31yEfbHsF7F1mokrA5LzH
BL+wjM0MptO6C7mEDfe9FFgqZHlwCNG+9PqxTjdsPQU/08OIVSKoVwuDrvx7Kw+n
V64CYvkCGojNBxsxXDj+CK8an3GEBa0wgiMjKGWY7y0ZHt24xc8dlIfkwBaNyI9B
7SPS918gUmGcS/dTzP73FhdfLX77YZVx4vy7flrNt92SM900eWiUQdU1QxMsJhKZ
7eolZXdV1PBk5Mgq6CrX78i8LyTj5BhuQPGgaEpsw1l9UG7gdUhBJIsyDYgONVDs
mP7427Xy9T/UpDpWqKufu29wcvPKKYUTose0pvlRMHpzP72HeJDm0chWalfpKVJP
cNjrHz7fs3nAQdBQnpBm9lCJOYUAmO5ljHlITmqd25+4g/mgrosuM6v/VjaxKaxq
sx911FAaKDGV9+7cuVwQ4gtVbVqI2IaR0Pjs8LFVPbaZ6dlIIGOse2MEI3ZJjTdV
hCFh8Kcs2cO9rsmVUa9z1kroCKJTr5GZA4KlUnAPMcLvppgkpLHM0A5HFJD6xrwY
92I0IA49CsqD7RkDWMLSlVd3bb2rn9ZgGH80CPL3bTTF1r58qCPXYFkFOu7PbhUn
r2Rp2lzsZ/9nMTRwl9y1+noxMnrDHIl1cEPKA865hhIApJMDftI4yl4ZWtfZ2KrT
pMclca20bynysNB+TCk2SIPvKRjiLWvWS+rnrJ1ScTG9plbiA6lWy3oMyHJAlF9w
VgTItO4XyEItv8FN1V80sSBeWv3N3mYgzwjFfbOVvk0k0vEypS0NCt65U27N5Nn3
X8f3j94b0SCA46NTk5nFx9BmQxLzCF9BXaVguFYSUkRYEcLCi5rGv6fSULGe6wMP
vayCW05Y7NMeZaP+KVt8utg9ruvsA4LzOSknwWa74HgMMIxgTB6KS7pf+sPV+K4i
Oxb2A8OghsAdd6hRsmVVKVUXaAio+5W60wLRBqjnhPJyGMXKWdDVhoBjqvZy4Wbg
frdPs0vJQsl1173ouO1O6eINc/q99AEb22FVp/U9dqJftvkj6C+JoZIYk5W5/3wD
AK9xyHWjBK8QNyoGQvd3Cn4Z202QuGYkP6fQ8iVo7jBMVe48mtlgscV0w/AUJSb8
4ZRxF/j3jUn1NWamnrOTyCTqewOVOTcIc9HIWX0vQcr6iXzVFmkHRj8U9db1fP6y
mesY6NjnoTMXt/yYYa1t1xfSzRmN+m+wyrn6YUpdiNangX/LXd18VJG/dJWC5FMp
m/BLyPVVLAy9vDnDYjoQbeGKKiI74+nGWIVb4dnrcmAzvB8Z+kquD1+quyO0MDwU
4RKBeG+ifqOPVUG+ssTA7q1WtxBZMhM9fPgcabuoZ+wY2xKQjX5MhU09YBM85Q42
e8OiR2hP5iC8F2EV6tflxlW5TwW+5i0Ljg1vKkYr91seMeTOIhb0LK/exfI98TE7
4OrUDu/9Z4fYmKVZ2znoHyROfmU5dlzhmB1eVl9xlsdurBqC6QTepd6mvBELI6Jq
jFetPxPHVR0/Rer61G9PRHXiRQPp1TOWGGPxnYYxmOqYt25GSxc1c4kqzguAd11V
T37bStB8lTaYk27xH4IrnNdrD40IbT5G9UtyQFvK/jGmBKpJm/qDBl56p7mJXHRC
fmK1QXwlYxinzZkAGbzj3joZ5uKk5nOahtVzhKkWV6HDnAlDQuwRGc3OmhfiRnbQ
5PArZqMic3cmldbb5NFhILlxWRkESSjIJAk/qCAnAbexo+BUXHp6M16jbjCJRRwP
dHnonzkMXa/vQWLPj/XIwpwsMay4C5yHM7u0Fj5hyOEkW7ORdV/AQRs/9KBo88D4
ZxOkk0oi7uQ1/JE/fsiA/XRy/ix/si7EZ5rmfuj7tlBYEoXlOvbl6AOqw853R9Sz
WTlN74q3RmOQVOCZZa7kt/w0DX+VyrOUJroOhSM5W9/NpmpvQOq5yvRo6MF5ZXzW
tvhhgh0qh2Rlf7/nc1kTxEuqyZDr51n98O/Ngw9eRHOMrrtvtVUlIsoScVAodhIg
jLswG7Iw2QWnad7n4kWWfM7tY1RfT8ileSa2tuBFaIsc15XwtNtNjUApijZtMUD+
gM2v1r3GVA1QhqOv1LcPLMw6p46ggpJZcQRCnMpEGES4pVqM/3KSLpndXwd3dHmt
jETpYTAqqGzN0GPC31PdGbd/WnGvBcIBZZ9iDhZ3d9mXYyGko+2EEKzQQIv4pt+E
DTloIHSarQyamtMyq6UkLdXMMMYRoDpTnqEF3VczC+v6U4UM2Y2r6UOzRHG2r4wO
PVSk4F+AHagXLdsNrD7oXX4xHotisEJDnuS6HZYFH6oh2/5A6skXwRuPz4/pOFx6
/4wcYjIFiLJ5J95dY3iqaBjMVW18JDyyb37uJ55rKQjtEq+F0LqiwXtviMWWh8fN
XHqNJ1vB4OBeuxCIfa6/IBl0bpSRs9sWAwJNzSm4QrqKCXYHmzv7dWPYrGHtlXER
3UPhhPCmM8qpy2TZXmuFRSwWGmLSjo4yT87lu5FboIZNf9Fw9iUc84SmD06AQcEF
lWpAsPXUvCAKYUZ3w1pPU9NfCVRNNpa6t/7cAmoV9S4FW7mFPGb81HaUGhY0IjNY
bIGyF8y/lVXr4UFv5orhGTBcihrOTXLoFFVdpMDvYcH/lEpVgRwJQt+g3vpqji2M
T7bbB3ZoYTk0giAPU3qvIWwHnyWRuWoRaB0S5nwGFNSKgMlD1+UaHmz4WisWBYG1
HM8tUiWVJ/CM6oJNdcD9uHxXB6qdxqkE0+spPfHXV0Vsy7aYVoz/NyHP4+iWYmZT
gO4ZEm0HacY73kYFOO+KwucBgD54UcnuLX3ysKNQxjtiqHUeAMLEdjdiLuONNwms
ws+hrYtWxHgn49Sd3weRyOmY1REEP516BO9YfSV6tsVXq1+yrkdPQpfBqrC77Wxj
CKKNcSIZY88EQH2CpxUag9xkgiVyNeZh1I0l6XxYsWt4K+qRUfx4QpOBcoNF2D2v
USOMqv9Dw3AFuQ3RWRcRjf6o+bJoVwSkfYj2J0sKFtMlVxphODJrY2nA8c64ixYI
A00QY/leGZag551tftVsIhTRflCSE3bbjJhgk+Fkg0aXxuiJIxbH4Z2TrejjVLOl
EITD5JZMVke6BnYlQVDTnZmR1dnoKvazVVM1Zt/mBQmlCI14JcrXrnjFB372lLlk
3rBdn4cWMt1RjS4IvlKztKdWqMVnkjZuPQx4ZWfQEv9uiw9uS+8oVJl8opv6cu2F
gtpLUbXIqRPbgXkZ2yvRlICGdBVq5Q/qBZapLyNF/4HkZ5IVotFVWUPom+VdHFCr
uD7+wUiXVnsHiC7ftiSdJPVPYDo/Pa5HN6HLHlCqjz+MIekucJTYVMY2Npq8syWh
h9VMswny4IilrsV5QdO7RpUDiq+lpmA9jirQIUkykzQLgyCLXhq7E9UAddHWeJfA
CYx26Q7rZVgUMLagvTHaQ49wQx7PnA3ispwa8mKdXhQUfNpVjBHMtRz6KRZaMJwu
D9shOPhrp+doM99R1Tg47aSDgoILjkMngH/X1eoRXeA6pcIvV28SAa3kz8SGDD8e
F5ZQTbTxe5rRW2S4GHSb0c/09IYnFLd2yPMMimBFfdRZ3CK/Ydnx/L+2HHEjLXde
fx9Sq7saE0Fdk+m1gUE+UcTXQNYrQCA7n+6blDzayyvHaD5cKsw7gz0o7H2M7FiC
bzt87kSdAM/eEXmFvpej//u7QXZfMHC/SVfwLEB7HRO81hVSWWLfZsNMSGJW8Xh1
ENPpB/zeccB0QbkeiZcv2/USz65wbP8Vh3/OFvzq1ZIxgsO35YR18NMIPFNhISJx
E83jFnlI+XY5yzOsug2MP8maUTxzaOTq1Uvo5aYDrM7FlKL5mhDj6lxyxlZdoFEU
Um5FoURNYtAO2jgzIeG/YHMDqKwhuqMTR6u4Rrh9pUg0BwE6+ds6YWpBWb+QIdT3
Ydv4gZJkCSXKwCPQYgykH5m3f8ranNNBAXtBFvojuQn9n5bgfmHVbQflaLQnsAJt
Wm0HefcEUlYK0zox8QE1RS3SnZaF6vXl8KiF3dO+n/y9bpuTavJcZhbarlb9WCzZ
mz06lFk1GsP50fG6g/d+D/Xj0amcaAvD7pHNE6pH5iwyWgPwzlue+yFfsWtqGdGu
hDwScURpxuPoZCywJE5Tdd4Y4ySfoGY831a1wIogK6529FLp0EvnlnWbg1f77QuF
CZPOwp+ywSY46s/tnnyEqBwA4TPKBhrUud0FwkXOMCaPLoiunqXO9Pr0PRxfaKQr
tuTQWIjrJ3YPmTY5fimcr+D0iW01xfICg1HtCh/dV0EZShVg5BpdSAH/Ha47RWp/
27cEjVdqY3UmXryjU6Ktts/aQlNGPEC10ARZHDJWchHugzTQtEMY4K1W7HlQYRDx
wswZF1fEphxP8LRAyfuO382zGZws0BwavtSh9q8KZGRQq2uKSXi7OwEQ+/nUydKl
kavwPvXLW/W9ceKi8NEQ5tW3830ZWv6P+vnqHpSHsnBbxKEwZenUSIVl/kGkD3BL
J9ZycHtcakW5Ssi4m5PFQmPaj94fzaTCar+zxqqt2yNx+a4RW8infj9tqSSx3Zg5
741CCko93CZ8NmuQcPel1jy94LOhL3KDj1W3H1NkiFWpo+vb2e2brcC4FwxAgnXw
BHvyPHrcE5h3Fr/LUozdg66V9Ffup84V2eRtC/jXfS/irP4V9o7lVF3ouwPYyCsQ
3FTqLETYMhjKR/4GhfczUvXRAUesZAiNrfO7RZQ0W6PRnRK/cYK7/9dLQybqmgfZ
Ozs65702fl8icjzVoQBZkZPo3ptYdMev0/Nj8rem0rLaW/tv1MeedV+T9MsSWH5k
7YUw5s5TBCIkwU2klDHIMyXaTZVXakoJw6+QWaRC/UMysgvGxHc7x7lRw1q4Wbl4
h9Nd1s9MrH071whd6oTeGrtinZY0TYkITvx0hWLIGTB4opUTbgNeZyV10Sd+ILHS
0vtXX6uAAPYa4wlkdQuwPbWo7VKv+wXFbrYWdOa3+y059r5RueV7cyA/lsOa6unQ
IfLfhyQiDAEmVBvj2zhKJT6uXxZ4krwbsKrpkjctHoNIJhEHHuFHb6L14TGGfqot
3gL+J9pbNxbYpCtsjFLR34UbfhJ5nTIop94Lr8qpvu3rZYTLW5bgMaqnIwI8NZgk
JxrIm/HnKICP/E8D62Bwm0mKIRv2HXEybe+u3nKYBmePykIq4YEromnH1fAMnmEs
WB3BS299PAwZI2ng6Tizi/HV7cEd8QAkqZylXdPefO1a236HXEMaRPZDvmOQlfoV
nUk4SRM+flIPqeV8G6vHQTFiutSm4GQzxUT1m1h4Lxc171f+ZeFV4Zw2R+pv7L2y
lxqxgJA5b7oiC5yu+ztsxm8360RTt8n3nOah28oGDcU+F7ljX0y9Sr9FSirrC2Ll
rG+y8ILPJ9YiewM1s9EnXK10LIxC5nzvZwgGeEmpQgQjagPQG0qS10XuPOBvChip
9g/WNxdek1CYhF3TYS8ajrnx3Oq1kOVaA2jIJWrnOkrShoaT97okxhF0cxCZiPZq
Qyh9hmecs46rNKBhptGhJVeh/ZcQCn9pb7TTv1whigf4F/4X1wwbuESDw6FWqNQ9
Y/bk5B33JsSarMifM9dm9Q/bmEjavuooZO8if/5A5G+luTNjG/qUknRrobDdIDFU
WA5FWGVcQldeDQDdqBwP4TjxfWROxZe95JolST7+9W+G+61w8cXir5Z8K/IJdphk
1ylQmgTr8vLwq+fhwTW90e8xw0lHY4dH8O7zneWtad8sHug3CU5vZA4URKs3LFgq
btZ/FNEk2SyhDvNXpIt1VJbH4/sjavssUWvB85rqvFMU35VCFJqdoiUOS6gbzIO5
6P5Nb+FUEvy7eX3xb3J1vHGxrLPvpDJkQflc4KQxj5UL6gSY01a9rEvcbGW4UVh6
DdNTAV4octVFAtx7TeEhT+KxQkmgMohuMoSJv4hdhwNCvXCULvPBHB43KyfrTavr
QCDSWC5I04Rd0bgucHcxTngooZlCAXaFUC5gZCQODPqzJLaFfF434igwCCwidqiF
0/opKTaD76HhJ/JDOxEg4UcJmkbOXibgAdSADtrl16LfCjPOElEF3cuskSv9xPYO
voi2XQULr0GIiWAER0U3CZTc4lki4AkoZJyM4UasZP4/SJKnUVbJnpwajr04HJtn
Z3qKNIBfN5jzggw0/kpBasVFZlVQw1hqHH4WQ5tzCcGjdipOlVLUmTRIXHLWL34D
Jt34wmD7s9j3m+ar0uEiX4DjWDVZzTQjXjJ6bAzWlk9XE61KAV45w6FWID7UTCIt
IoQSTpRvTQkqxvzISCAk76MojXLPum/qxJFU6bfYwpv9CJqTmdLiRbM53IO8IU3w
P+LcsQzLWggEMcFvAXkwP291SJq9Knn1/zOVHYCAJri5IFPMFDPQ5fbrj12W3XOX
N/SWxZU0LJKf77SJXoKxbv0m1tKDSzoV3Qw7HvROhKP8hJ2eqWY8bzr0kDmw4uAG
KpjVzMZ3xQL+PCBDJmBa3h8eJXRZZDEHIZHxuOFWLYuuLzvmqq4Hk9gmWsii7xuB
0ysZhOkkiub6bEHCW5E0XYNXacOTvPxNtGXINai45wFQ7oKzBQjDchg7bmfogFfw
bF/IGFqOoDkic17tjh1M6WcfIEM+ev156PJaJm6atyvVBdR8cPLTBkjbn9IeBYvP
sfLTc42zShhRuFg6EmxxSWgKJbinjnGvNb/7UKER53prNGKc7FQFmMi6evxnIH0X
vl3/vhPHLST+gv0QFX94xAY+75xPgSC9oSBkXo+AjGnUv/qwHt63hj7pDz3XNAVL
pbZQL9ZlYe1eEx5l6OopjRKcSh2rmFQdh35D19xpejTPOPm7KsNxI5iWF5C980Fb
DAd1mMZ0PwsIyYhUclqW0RDQj4eJofeXuxrulVIte5nIG+efVkQe0zP8kVCj2s11
YwZBbolYJhRznoKIrjEpZyYnfZctmpw4O/9i4g11ttTFta5z3T934KP0fRwcoxig
la3QarQniX5d8oN2m6gY9/Rfsh6dbQuMWx9p6X3q2lJgUR4q4mzK38yFdZ3WcvK7
PvohL4pfCNddWryWp9Mw8GIQsPSVyI4wbslMyIv3P/KzXasbFyXlY4JHvEjdKbJB
Y/Hm7IxRBb/fM9GpK+dUwRKM3wtNoobo1tCa8X+tKmoflNSLR3Qy+b+le1yTc11h
9Q3jLdX7os5anXue8W/cxHYtBDyQm+b9akuB9r60GIpqj6dujNlrNHC50rVCFzP0
bFpdCkduvwdVswIojFIIfP3X9MjCnbjJYnKKHFMl2TLVlRa2AEmCQO3DqYsN1IPf
unzly8OuYOs55IDE8QJDIKERY8RXgLj4xE2KoPBgz2bNBxEM45gWmi8uckPRV68l
eQI3leWmgD0RNnmNFwoPNTg/1xVY+OV1tv1JA6PGL/fniBGx4bH1/X4BVz5LiEDa
IIC1a0PqWPwS1TPdXWxh6SZXln9Lw4ssLwcyRMroW7EGJ/KZjAtPPkUO9XGjfmu7
Ysp0gjdz+vES51agHDxPRov9RDS1Cx4UNkpQ7phaZihzQ5McNeI/SH9zam04m/Sa
OzSRzhTL8XaS64fCUpy2a4pUDEZB42V/gGwYjjv74VbR9NH5rgrCpMsEU4QknfbX
o206FwiCovjN86mOZzPsj+nhkSd7pcUHpqJPtV/oPusOARsO9hJEDdbpjMILaQD2
bxfHK6jW3wYdnUack0qDZYxyzLQwWK2KpA1ndSqr6FyXYsB8EA+6j7eXRE22oMn6
VeWgyuYrA4vUJIglpL0xRiQRUxHS2evGiMAHqlklqLdn4N8PBJt9mSO+EXAB+8Z8
n9bL/C2bjl6EqUmtTwoBLCbJvoFNa7xUxeliI80BJjnfN3w0aHCs/i9Mt2TCZYUg
W8iZGyxshyKCUqJn1EQmtekDnuFMTUDCVBb3BkOF/2M0WYvKbOFPo20xdpEXrX98
BFV3DZh24qI2YfpJkTQLLRbW/aIAWoNQuF76lj127oHDBgWh3h/KNgZUQYIC2BXw
UcIdSZ81nilZjQDRhUhPBkTTLuZN7Uy+uJMiig2Pd7vrodcoQG84qFVnyvTnvNiZ
Ch9Vd6fjMctY6Sz3/RpmcECcL3fO41v2xPn4Q0kfH4FhXQvyTI44uv7a+NlkiF8m
r/1UznZW22gq76vvyWKYuykA+c+/AlxxalKXERno4dSP4VWBqpRF4vX+ooykw4bd
NHwQWa+TeLS5vs8xQv0ucTA9F2aNU4V+aWdiQqTJGy+/Wfo5PplF1SpU619K1Lmx
a2T5d5JWjLdlkD9+CbqSrRUipevAnJV8RM2U+1Uu9S18gxK60m+JRMOuh0d483pl
0YbhzcA7+mNXdpiG1T+o102NBJmaSc9v0qJ8a1qZshkBQieyxCHrVhnlNvuXAB8v
0vuQtQ6POfq8wb/MNN+F5lEPVib/FuJawq4HbkUs6Px/J4LWxhYJjfERgrmHRUWI
DEUSuNdfBv7KIuAk0nHlYgBE7ONV73/QEbqDOk1d5W5BcYIuEllR7/L5jo0e1FEW
qIfOX03EfXu8hY6mzKuT70xd15ZnHeLYlMMjk71Hm+u3kAv28XfboCZs/hvGx8qV
G3C+VND+vHBXbZ+ZcjmvnKv8LFYeNI7kE+WsoIWF3vfD0SOZXsi2QAOa5ZWVkqMn
JHfRQcid3B5jJ1xpBrHwhwJXOolbayfqaX603mudS5EnLqbtDMS22BFCKzi5IwRG
aOk98mR+eaM9mn5EVY27ZbU3zkL00DdPpf2IkQpqEcJCHJDcU8Mxpdj2KEbmZHDT
ybeCpEX9sJGYgix/kEE0nymusYjLpMSNYO/pRBj0oHAUiZ2RG/MbH2DoHq6DYGjg
erDPtL8jBeApI75BBG22dEjx62Ud9rt46yDGTGnRzFNru6EXuQjLCVmyaMmxcjox
GyG/KNKC+18AO0/FgyWgvEWpvlqY8szUwoIARI3bFWXIHUE5Uchn2owpVuQUEhKV
6DMgR4mhLUjncYFDFihGCaVzF+kLHzKFpPA78nq55/q+6HGMZ0xTm7aB4B6t3RJp
R4dsqLarDWUJ4sf0k99M/Ywck9GYVIF5pbwYXfgrGt7iEx7iEluozBghbmTzskB9
EazL5B6cSRd0jiDDHQXu2lTyr068W9ffwAZ8clj8kG38EUBuL+xhqkuHr9Yq6Ymg
WDYAjB8kCtK5u6cfibGDPs8fQ0+NVSDaTVEzuNq+zuNiWA4khYXEWpBq30wT3fPx
YXEPipzGpdZCs4xcTtQFxJzDimG6DHJXpJDSAft4c+Ky5gF/YDGCr9TnFdXTo9X8
psOHku8Z7x3GC1PjnMPFuMcnjFZcTMYQtXSyMlrWcnsUkrsaTgmDOdIFiA/GORFe
L+SeAmEQeosAGoVJwB+LbFYAPZxPj0m6yJj5vpv4FJ8D03PpNlCBlOF2uxDmoadp
AOiilcE3dPQrQQtCcrmZB3iFS16LGjrxmAny/Dr9eq6Y7juxUVt8UhdZ8NKAvVVq
jYaa3871vmJL8DZOlfCaspy7DY66Q2xeJ+3eRgMpO5r+RnuMmDcFssF4Ovm5DdOm
AEP3E07HpEqJiaks5N4JU82n/YbokJuTRcKLsAMiY/jAUfLr5MzcphYS2FTNJK0s
1mCqzrW7dxMzqKylpnXxRa/+L4VrfSATdKZakgCrnPrSqp4wfhcvUlLxHewhzoRg
TauFvaBMD1FAVFvVV6n8yZSJvRXgwy3UqQmAmWIdI/Z8Xmkq8GGRbRSu9LlL1my3
/hlhL7ibAFA9J96vKbWKAL1UGIP+OoAbYmc3aUtCvN/qpnwflKfRIACR9pPmZTap
Vx6OINL/fMwE8LHrdVHXHgupctPKxy9HLdsIAvaEZc2tNKeWDTZRDk+Ke5sk5UIE
j2yE0Uxp/VyUjqtVcO0taCKsoA4fs9dzOQwUT52xxBrwM2tkBsclhR5yoSCaaA83
Oy0Y+ui5y+/SKVra0y09O+bppVaMPVSUIDvUXq2cZ/fnRFtafORJLnxNzpUwYh2f
g+6l8pDhaocKUbNpdMJK76to6ATDxgluH7ecjXMSIg4wel9/1PEC0EJX2KGGtdCH
+viwizLAkkWMkhmcUPLNAUssnvREL6EPqr070zzKQvhv3IjsZRDzXkkFV2bsQwCg
3GWkZRmYT6E0p3XU07BptUlFv+kFoJqY5pxUKEJPE9o4o5BTlW0febs3bYnmpqFb
wwtodl0m/y2PvcdN0HbMK4JmDlRagm9quO4pDL9De5QpG/HZircKkp6K/dzD7aVG
h6J4ZCinAig77OR6W1KnTBVIZS0nyzSAO7h1dO2nj7DzMsEP8rg7VEM4tYCxeC+u
DH4eE/dFs4LFUZoSNMkHFUs2ah84jdUOOXV1CiwAlqTAZhdXbo+sVd8avs02iKFw
5ZAtw2TcdA2hLkeOunXzbYjtaoOjGhlx20aeUnfZUc0RGQKp7IQIjgCMQ2GzTB51
DvvE4GaC5/ZgiIhy82+iR9DhSIJyRufnu1SLtOHrT0Kvjni/i+ko8uphFE7e4z0Y
r5tPWNZ8SsxBw0aEuRU2uQw6fzq0x45dIjb/V+qCtqysuZJDHJlQmsPialky6J02
BxExyvYBkRqY9VPc4poJpyW5QAabfjyR6HGaGATtvTbgWpFaLcr+Z+NsIgC8wKld
oWnd4Lk90ELvLdfPAmLWwT0KVDee7ZtA/vkhyZ4hHgJJwVVOcf0W+OB5nSJ96OA8
KXfskCsKxcGfsHcdAovpTZS5H1O5QNvd1tbBnu7YzFH1menjzl6jMNufX1Fju4NS
7zpB7Pd/+cgzBOHkN9MTCbRBAbzxDfC0zeAHlB/Y/kIh543VQiMIV+ySeUFwQqr2
nkjc0jRMXIKB+Esdz1ro5RllS0weE+dwV/8Hvf+1qgBitRdurYC5VWYt0bG87KIK
A7iyU6IRrFFq5pVIoSsqQTtuK4uwT0NkBCi0NZmHKm71GVyWKfAD5LrY5ladDeSX
1bS5zifX1RBzpBAgbHyfhzK5Jn/c0xzK9qKSIL3CUcAD4aW2OrLfn7QmXRWbVYlM
HfHjNDsYcLt5MgaANpFvSuo5GL9Ou4gEYdyF/4a0FMUPi0sNCGSx4zQGtpUFMnzQ
9gSDbKcV17eTZT1yQqYX5k0SwN5PSB3rvsyS8P8bd04spu9aiIuQe4L2oHcIOHhm
A5s8h59HDY40nVsxhebmOm7McxuOZG8ut3KIMgjol+WuX7IKxjcgwC5pu4hH2pVL
fDN+ZcJqsMfaVZljtuv+Ufg9AME0t7ijEZPu7qGscdyKJA2cPsS5GxsnNN0Dzkl0
sDx6kklhZhl90TsRqID/QUFZi4+kuMtzecdNnzaLmEPmJ89oaTapHzBcElEUzoUJ
c7whTVF/7rk2iRpg2dSoHV15ir+wYxYQsOzyiPeNOo9z0Ab9XYAUpPDZxQ1zZiSu
i6ABv79Pdbl7geuUcWkNiCowuwNjhYUcWfs08iV3XAP+6dpO5uXRGwxNKbRPOLH/
xuxsrj6d7qzU6LVYLm83ZKfdrzfH1OQ/9joTtxpOsaCMo+qaFc8IGK0cdnc8YoAo
E2aCLJRJKhz0QjL1wnN/GtDKvYGemjlreZ3QoWWyfMbpm/UFuS95edEe2CPR4d8e
sxEhcJnxwQCbL0RvJ6e1VTBghi2YCvRr0Endz77TtjakYRKF3Lj5sXsXECRGEf8O
/8BlfM6QduxjVzvs5ZKMtZ7fkJr1YETvytpHQfHhp5a9R4mR73wYeuD58mfMeN2p
rwvkdc0sp5SXxPD2LrxDDBg8dJ1EGmDNxHy6+oRn5Xho59t3H2t3tknN9fRC3XrV
qUjfH4jDTFva9ePzO5n1ho39mzMgJzpuB142vj3O8YiSgOrj2brLFD01Z29g2y35
X6l07ztsA7WmbtLXRsu/2vASDv41Gder3LD2jN5hHY3if9Ayq6hVpVErfg46lJ28
v1/LrV+O1SL7xc1AZOG8vFQM7jUBrtbKBWhneo6XCOxdpWm15TaCJKtfaJ8ntnkJ
znc9iWbfDwiZ+nSwmHxNQAm55rPTfR940OJf1MBeRaQWShlSWd4fqlcsVnT5L+Uo
m3pyTH7x3ya20p2zXxYcv5db0eFehZPmtUI2LAgIJ4ptu3jP06Qs4jNJ5JfvvddE
fzLk4HFu5jGI4QjkaqylarAaavCyef9EcLw+UssaJimIHcpJRICCj5WX4WvRpG09
XvI0M63LZjHGnXDcBPOXdyJiUcmmZVmdv/5aOS1RQb5nFTBzCq1LEWUL00bm9maQ
+dyzc8wyVKNPhsoKIJbV2JtG8nBjGjN+T+9Rfs/tXU12kC+22s62OwOz96JQajQ5
drLqEtalPcPikZRUfvJIjtWE96pxDigFFrQWYvQTUEuXLS7uyJCihIUe2dOloQeE
QhSqN2RQz6FXp5MBxaGA2hR/7+LAz/xBzaZy2I2vc5eR7+dtUWTUrIoO8dx2z0U7
TL0rOUuAilh5Gk6h3HUb5NW3H5QA+/mIivU/dVQlH7rYEPTEW4ES2n8gdjQ/51Ao
64wmu4fX3sMZ6WNHUkRJKF+Y/4x7ErQhVMflLGiwvoWGpWku06ulHr9IKxU2+H2n
iBAh6RXUl4n4gOx9YCm5WMq0nYvQoi8JdIMWPnPz5IL9Ba5svEY+MKYyGTGkm3u5
tFMomUYdJRoqDWnEdS5u/YZPR5TIxGhZ19x6FUJdvxmQTSxY6qKQ5MAbbcoz2tBw
J9zzLu2dcze6B6iaKQcEfvgqWzX70AWQWAo/uOeWg/BPrNZUcUpt4/7ocmDBi8Tu
KQwgtKlE4J/+Y0c2x6qgFkH0q/5hVHWFAEDG5RDXZpuvpMshYhcjYDjUI5Gmpokd
n+l8L4o8e2yXSFoRrOIyrW+1DDkUEie1YW8Pt+DM/jxTEBfNYVOunxDw5dthVQAn
HHIoDwPSlgLCDa4TBLYGXJ4WUNq8jCTOPkCWCWlgXjxpBlCWX7sUZIBJkPPPfjv7
1FMkcdiVYsiBvBSOyB7nRNfqP+2usP599+p9QsNi0afr0M7nEaBAFrIrufspyOPF
ipRpf5IY6ZFkWiXjqw35YK1gB3hM0e88SSysvmq2Fotz6gH86r6GznB2SW9ND46A
/gSYiRINuAX6Mp9WkGTH+NzeG4C2xsZYI6Yl+uggVgfnD+FzM4awdkEcWCV3aWaK
maX9bkxE0y7WuNoKeYgGvmgopuWvJfnuBS3WCaiWA955LkmM3zF1lpABfGUOBxNO
d+djZ6ilCTN8TNFK/UoA4qziP6vkht++16xSduytBi4KurxfJP+BzHNI4O30h6+1
LFz5804SUjk9J6K6ThjRP2az40Qq1XVmohe2N+X2KtqIVJaUtFUcMWqrsoi97w1O
M4T6bgGGM665zPlNQfBBuBu90rZC2lk/f+zxnUITrGifxHihQjORfAeIeJ6nXANL
qGE75irDMCLjm2kkcmK2Ad8/rhYZBrqtKJ6AZvQgaD4Ihrj908yXoYCP2Agr6n6a
7IN4KvAuhliW/j3QwTe89NmDWGh0E8DpdHdQv3MYvs0rWsioTtpJ5jvrP0y0wIhd
dFWlpqQvRPQ91CMEQlRdjD1/c452BkOvgjWZcaIQrI2GxL5CT8rD178e237QAItu
KECn0lWCWZCeTLK+TqIYXApsGU91iUN2hmAxuWedDL6uor623XKDFPPAOMulIo9z
Ru1r8eUwua06o0ec/UQzib69hL6XXLuAxRRodOMOBsS+N74eJ8auBvdSxDc97zLi
Z3S8ia6ttKvp0nPL1xZb4JyZ9J+8lVRrwmTMvkWlMbzLMqWoLSttLjFtfch2zqAu
bkJAWvTfthCKOjEq3fgsYsVwOWo48FeUnQ57Ur6SL5a4eM2na9j96Ici62FfACCg
wk+v1KJ2znhZ2QzGta88lBNeQq4Gg2HfakNsFJ8M6i6VxyfXJo0EHVFA4EBQNLRO
miCdwFILb03P28ZDX94gkvAsq+daoDmwtDpNBWieX+kUNTTnblWHEacJVqcZ4oYa
vx4AFK5sfQXDSYr1TxpHZ2IT2lfrEzsvsxqLz/q5vd8bsv1E7Mf8TQ5w/IjnqLvH
edv3mjYUUnIK8v/8oCRp1gefzTMOYXPDPpY6WYEfs9t0F+hzniv43+CmLgxw8x65
3ifBnTeMRb1yBceJsbL317Dbk7g8mZ49P+tM0MtDCGwoB4d54DOwthdyVe6bAtfL
MXfrbvMM6E0WEioAGO/TphLdQX1QFzV0D85ArUmknn/QPns3jLs/TCTYsu2NdKlZ
vD8+SiCr0o/CGq4bD2hRwMpYzixHXylLIMlc6M9jj2IUvYSTrQz/b0dUm0ulolMh
FCAszSMJPXI9df4XD0AXgKGiSFNyEPbm2zKvLfoVtVs5emQKIE69pelxkt4h/PYe
qouyUS51iwsjqpSejNSbe4OUbw9uOzxsrmsH0azFE/7AJcmcSsBrXx+Q0yiljPTd
JUIMLk+NbDrLPZ9BFEi3GgCmZobtmG6nttxoiGk3xd3Cs7lUUZsT3yNGktqzWjJy
BqKKPqQkPh6ATHGIDlq6Ht31Rr+j8vU4chhXwtw/65ZlkEf0YCKK2RKJYPwm2QQQ
MMuO91kfDoaXj5uIX6a2HeOV0z17eXEFtPQmxT9KpLulmgsjg3P4QdD/4guj5l1w
Sr4WddmCkkuKFL40QKnlET4s49zzlPQ+q5K2L7+sBKukmRkSEhOwTtjBIS/6A9a8
DKOKgszKa9VMAOD5jKZAs7fLHNknLg5FrjbvigucvQmfTsvgLeneLd0ZcVCOD8EX
BLukrtiVgs/MtnLawt+NTCNKhWeSXa4j3S0RJjVagEO5RzVBjYADRhp8cW0cwijm
CxqrQHZOHx/ri9hwnxMEfm1HLhVamk0fw3cs9Fiv/Qk8mz2PUaWLWZyAITi1omMc
0xR803Xs7bOqm8jh5s7jEGQ5jInTV2700r7KKOsVXR5mCJbvzg0OESFvzQKD0R30
T76h0TwrdpkfpCOifmHxpU0AYhgTKyGc9C+C41zq4g6lOJIRMeBeejtcPB+aX8o6
bNBgaees8Y9SFUzfFWs9mw5rOq9po4hlbKrEXrUjlq6zC/NVrWyCqnf0R00T1aJH
chpWVaLk99/PrchapNxXdLaGBymjEo/n1vRDzZ+gMKHga0erj0QMGvrNCCqzpTlf
sPPTfLRa5uyxZEYxV9yB4mt4PDOG2Mzyf6fMrMmij/EaVoFzAQSrUZNytYS6nE+c
gaQhXX1JKZxzsVz3NfJL84KMcEpqDgJUn/C6DrDKBdp9LDPxdUWOvvL+SzI83O6g
9Iz+BkW62jB9bz9YzNP6GXQqSaJvgewi1+kx6NSQkZridN1RlppfJy00lCZjRK6c
1puAGJasZ4L2T+YS9Z8KgOBCQMSWNH3rhqQ3wA0UvMMTYy90Qwuvdr3amToYoxDP
ZKVjr4MN0gTalEYbzxDIWhX0JiZDchS9HMezGGUP9f1o0L8U+7Y6QBzx24o8M21G
7zwHm6R7fW9aHZUOco4T9MMWbRUQXwhr4XLh1MxkVNFfjWca74SVlVcmaSCtmrhr
PJdLB3RfmyVsi58c/AxP0Ji/3tMvADNnlZ5hBAwbQxKoFqfReutmafKt+PrfYspS
FuDCOH/Y1lEVO14a/1isrzTy3msJcTg3B+Lk8Ce+UHeRww5cAZMgk3M+CcJmLTcg
b209PKIKSQSoaO59nVYQLxHQqz8x5JcQYI/ltdF3vK5L7NuuX/UZecObM4V2DxoL
ihPxOIeP31qbYEErkSjehszW+/zYjyzK0NZTG9ZWLkCGL0Tq3Nu07ephq1rdwCGe
tn20ccDqqbpjotNeZ0pA2fw8aXtg4QErySAQ6qeGe2j+rmnxeyP+pCyhlSX41TM7
MtR5TUHs3FP251m/LMJU0e34lnXQPmqecNGx13ttb5CZn0gs+tZm5oIq8Dv6riDS
85Dt1jXrXQTJ5BkwJqJ5RmBQyW03g1nw2CTwVvUuCmNVKOhQc4EfnAFfNdvcsLz8
BMes7n/LW63EtsQqyeUfMopUXZzEczQ+GuuRA/5XJj3qanSVZQyQYsM0qUfxUpWJ
/TTo2kxgS5xZYgSXdI0GpOpe4x7K8r174UuGuU5Vve+RgMSDPwx0UbhACB1Nuadk
xrb9LcD2O3IRFS5rgAKRhKdGMje+f3cIOIR4M+sBgLbXK3XtayZYRLe+BAszUl/y
d1e6cEzZ0ebxWwGGfptOy8VfMkrr+cy3T610azHxo7k3fZNKgWL21J5QcGbmgguf
oY+53ectro3u22vHdaR8Zt8iYsj8coRZmBR0z1dlZ1tm2vEe7OBfuIXDtKGGOuKj
/n2quSeCRWVbg0jM1dh3F6oK3kc4W4LIJc1QRzJ1IwtVOwBW98AVdJeysNKfBnBR
81w2pLkr1aQ7zH5z3ELWrYNAZ8/xJA2A/lYC4XhhwpLUBTpTFBNdP44gWQisXHLY
HYhXG+9pDp4HeyKV+D90wUtVrtDcaUJSZVesrXnC/1vuzBimJQJE5c7Kg2GnzGwC
FwYeCh2tZ65fSvAjAziz1mzaSKCr46I3Ixq2CktEUmGUJ9/Cmgr+ZAhlTzlyr2ZC
gIjQAIdXonBMeoC50cddUU232qB+na4l48wmAX3BuDbNSOoK2s7rFVAe4Qy80zMT
E/Rr8HH9ivZm74gyAdl09Mgldm8HFDXntzAqHpv3F3zgYrkQ+wB4T9OygOo52cty
M1UKzvAXqBxqqiDc9ggVQQSLfdn4kAvGhuae2iu0SOUSBhtq5UuXSr+YPhgL6kUw
NZDlE8Nit1apfYUOjJqBBxiHAgCGNpwlxXwvZqlKP8zMP8wi835Y3ZudLYd9HQVB
HinJ9bzqnZbpfyyPYeXA5jo5wZgCTZuty5DmpItEJeUjcAYLqcWftUi7OYL3U7Od
3bAGFwKuo4827oxPwqaTgr2jd9NHp3OxhUJ/KwGyVeV+H3sOBbNxP6aA6g58LVif
yuAB9NgxAnwUZoOFSVXPurvrrg2eieBXsqF7dGeD+J8DglU0LslJcG2tniosHoXv
fFe8pigsci6AbNDrLa/0+ZckvbQM8iwr4JJTcSNBIvnQvHRewyfrfGf/ebAqjbEK
fwnUthUvjd9Dk+0kTQxgGzufhLsTD4BTZIXkw0124GaXqYbiitqmRy8cXPBxD02U
858V0ZigE5qpaB73MzJ6SNpV/UCUs4N/TJZHlsVJfI7HoytiaGeaSqEBeuhE5LKI
IUtWVA8Hb/tfUs+VpK78V7zg1psuVAEqEPSEeEkmZy3eKP+8QhlL2YqbMvGf/peV
ZA1UtOaYz5fMgKZ+FWSYRmPgJYVcNEzfzVl+hKrEWp+2L5BOC0jW6S5XDXteRgCA
IcZ0rcMHdxa+QvwsplXaAPhr5p6thpLVtmVmMh4t33Pr0Eid3uaXsfIE1TIMIXcK
XNL4xm5tTlC82PHdY8WqoeNSgXqnx494VL8nmpZmoWv0OV8kzMZTcnWFeha1MRbS
L1GwtCVpqjhMKJL1FenEjhimsIrYiFJj//0wgkB4BDjYbvd9ymGJoAPxUaJjDKTY
EY6mRNrzuH6h72B85Mez601z5RwKY+ufM/L3pBMQajbJDjQVyjo8NoxNa5OGRhOn
w+73h5zJV0pdrO+uwS6lWhWyvAI6kDrTSi1nFC2/+k8PxQ1VmosgAQDGrGUT2vyI
6pZFYTMeuL5J3uRi/4cHUmrycYzhz/aYkZwgPSFDGROokf0Jpl0PY+OXh/r1ayu0
mQMwiTzB4UyxYQIKzr6950z3YtxQ3qHpy+2iEvLGI2aoifLESoKMXbLBRSRAVoNf
l5dpXL6WpJdcf9zy6MfFOGJSoY3eEEcxxOOqZvPwxDB8rjgTzTkLvsEVuhtr3S7W
N8Qp2PPlrblrGGu9AZjyCkiI/MI4rMa9UJ4YtdqLHEVRFbCGSy8H8IGVlBFgYFJf
HHulI8hHGQgmZrHXENS3ZNlMM4gDtnrD0FEi+3aoN/y43g4U1vP1Q8+z/thDfSRE
T3Xx0aqRPwzS3P5R0shXERKOCaq9Q/HS+c8X0hU4Q1x1AOH8BkCbvYg251vXFztZ
JL7Ko39S6nfyo9V2y471LZddKCa4P7++2ofQM9SJ2ne6FuZS9WJ94K3MosLc8dYF
HaPedMgs4d8OmfNmkQ3RK1yG49qG0zqAYweqysUmsYmPxEZavpwX9HUZacKUkUXZ
ntX274YBaFIBg3ACsfiJV+TMYiyqvVCUEWDNjobRkxUmrPp5TmU/A7ujbObwhSIP
EHAIZMjxoNdvL/lZwPBFEKLAxcw/p40DikUb1fdUCWQ8HTgfPGGO2X2TVeTXweaj
aQ3vZEKWr0EjVFvykyiH3VwNDUXeS5U8RhDdAwKFat5jylS2EfTFnJXpYwd92smC
Q1NutZ+LmSK2Y2wjCdgb5wP7ScA7HbYU68uhvKRT2oyDxKEjIndnfrWSAuIpCJer
Sur2mnZm9v+B69rOPBSdM4T9Nv/NBTyUSCvKxWQ+BHak5sn5if0Wev0C8EC4fq1q
fGIkVpityasG36AI5beUL4kntHEGd8bVCE6/MEcWLz3UTe3MfZo79PZfLT4hpbmJ
U6q3vYcvM4+vJPEDn3wtLHchrDROp5zbXTpB2+ROMU5v++6x0MtRGBJRZxfSYChe
0UbztzHFcqk30YCjuVb8hoeCg116FPUjIEnjg6t1OnUpVL37T0uhfWAcwafhHUWs
x+xnkfRg8i3BS6tGA0q7Y5kwlYJvBH1YNcykaT5VsHZidj90SVlHvnMXirNl/v2j
jYL+hcWbp87LkaG/gtsjyH4q5ZvlHBBULIsE6AXe6Ne15uT2ADjcMQFlhYkB06Rd
QV/RAS9hMOmoOW3jMdxeZcX0taoiALYjH+++Elsq91M+PH+1i5EGFUgbXBoyZuiK
l8kaTQKPo04d6CQrj2v+jZmIQFQOFQLt1hf9t2dwKZh9f3SUBA75uerHzVD9Xu+m
+FdC1o5fIYOqpHseSkTGXmm48zdxtBPuFaAervjELTqxAe6vMktLxEVjs3if/bDm
upg+oDcw69r2H28kmGr5zZzGUFes5SXpB7Lo7rk796uHLMZybaBTzAES+/5j+FwM
BJjpDBSKzaWGy6bd+BpPHPBWnwBHHMjDGxyUmaNbopRU0llqxmxlXzUvMU0dZQux
YEgxj+sHPnA774UIMfj9YUwMqD9fIT8zzyCfu9N2DuAQOE49ZfWoLjN3S7yPmzGF
49dg1cWFvEbAuccaJuQXceJRDYa95IguKavxnL10Y0ogxV28zPFy4AkT0BpJvNs8
bQbBG0N65ZgOjHhg7FdU8wAwMSd1xpTHi5/1HpAYhKfp843Wlg1gJP8LG/qYy3hO
3uMW5iUSyS+OY+3iu750qFfIpWKfHfA1T/70KtsSUSpRuvK1295dSbGY/zEokGGE
f3cFsvBGeMANB/wzaLNVx5dZ/C3bTOs6x7f2fcL/obfirRIQUhVjlmBwqbOpDTkR
UFph1VP9Kd7zHyPLPBh81yQURXooguZmKvPxxoYFVd5kXlLgek1IY2LAcaplfadk
PjzjIsT3V5ZNjC9ToLZgy1JIFBDLWjyp363oedfl/PoeynUC5/l03aFN2pxUrBFb
r/ngMXKUOPjCS87kXcLI4wIRxm20Lm3HRsEmqulv6Ns5L3VWVoRVIpNE5mIfI5It
IZPfKVcZ3Zq47w3F3wsfCe0QyeA3wgiXknactHicIQRKihDpuO47Cz46x2cIougZ
2JQC6AB4cvD6XaD5Ba4SoWEAsQhErsEbEFwHrF37M1RdmhW/RkaZzE5JQ4S2PCmr
Jz00iUXufGtBKgG55U+WeDM2zqZKHyb8RxjUF2705ZXoy4TMSc8+GhW0oBo1pdHJ
MTXBtb9+zMyA4v5SVQq+fxOmiko3AgqfhD3Mywez+RMRHF/cBJQ5kAHIGBlywPxa
M7yW+tAvX+9GjppR8OyJg8b7zFWCT0TyoTi668rHZ20OQyUYxkV7qoa80A0MQZ7h
5applsHvapVi2gFMiYPOdWcY9FpGpuzjgocroQwnQ0zeXjf+/HsupvlcGZzF1e4H
qyG5HhhZ83VW4iFW3/amAu9nbGpGd/nRZzNL7bRnb/Rbn2fAB3VhLZoRRjG4dg1c
GI1e5SsOIwUCwKrToaLclfIxzrtkeiRxutrEYap6ya6sZ8iRkqAd1z3OfhOy2uUX
3FMheK/+l/si2QQAN+ZPYcBICFOZ+ywjwgJEQp8X27RI2Pa9Xe8o1Xu5t1QxXBhr
kRtxnJDDZMTeboCmnzUC6GZwzz/seC069voowua7+Qz8lXGDxkLxyGWkjg+5FyYK
J4CAL21yGmabZ8Jg2jNOqapN9qU4k8OeZPGubIAFT7+AwHBNfzjzaVFdrpGr9vTi
SoAdy8EWMQ7zKxjoSuzeBCVMN5D/jpw79HNzcjKvKL1mUk2LpDh/23VbnlVuroKL
pBS689IvsRBS12jguzeRQaS/loWIVo2ZSQbc50DhK4m7h6pFK4OMqceIAA0nhBb0
KqoT+yfbGZJypJh7loMbUqJh9YSOJmngBR0Jz7OZaIXhR5+hA1dqX65USeDHFnP0
kS42v5Enf6LHpOwT+wI/GVXJCXgo+dBDLHW4heVA0MsGBbse1DOCaglj+gu7NSIm
pHS2CTTyn73Lm1uyGSp0jgXCvwQ5yl/3/vBnbG+cxLJFr9Zx9ePSvhz1WzpGC7uW
ngSh801OBjYhlKG4CkpekuGXRYmxAOCthUGsoZ0G15x79Ryymp0N87rYK6bQv15Z
2d3X+RRAPQlw5FhfBuyjPfsdjk5TBJ79lfITggLdApdfKTHWFoNj7NT36R9XcLdH
kWTIMnSKoC1z9rsxJjsZPstRqhvc+eKf4B4aM3/pmAgeW3/PgiMaTAxKdJDc2kW0
iNAvs8ywJAYxtYsXu+3HqH3HKF9qb6jcSpxkEPq1az/UuEu/mgIbuuzgVzplekaM
8iCJOfsqCl2YaV9v2rF5husCZXCROJDpUD+v2yHkBcGrgnf2fc5RJf99F0JGcFF+
o0r9Mjqa0DxMdpaG9MXx2VwPlBQ6l/6pvx7e87FQFcL3Iawf0gqQPJGauRSRtKdp
HRB+N9B1ENamT0ISUBv1qfyzOl978V2OsKK60EFpwrFVBYA0UwCjSaLL4cUQl3it
VcGH2VYBK/tMQhLGGIXhnAlBWsJh+sArzC9HzMKZVAMiesYU1lbWEEA9xKpHHAae
48S4/TpfZ/mfTc4Uj/gUor/aQ5NGgOuG01zAZ8BslSOjdQUaRuWrcV/cudzYXA/q
rt3t+VsLC4r7Z19iwUq9G/MsG3FtkrCSVTBHMgueIenHP7eG9+kqgUK1WAdaB0/p
fvzFwrLeZwPZhvkOrxW4QON+EkRCKmc8DI8LTIpsUoAlaDouco4z6Ng4uDuHFMKz
BlGp1z5552e6+9j1oin5XYZAeWcElA74+TOXpRxV5d6V9dGZTl2ae5cUGmfd90+z
OrNE7D6SHLo6P5i1VIKEezSnm7w9hsUsnUUH4Qn/in1/2mozf4zZPkQhSihx0Ih0
vd8arVY5YvwKMgPeR719WlNMJPiBZsmew++QLuTa2dWSeIcACkpRxdxy+GFH6GKm
NiZGEeH4Rii5bzpa7fdyoWOKdDn7vNQ8scw1ypxgAeY7yETEqN+r2VIhjLtFK1S7
a8shyu0pqzztVvgXbmVRI0d/awwxZNkuHwI/CkfDugm1uinaSx9UkRcpTKStma9h
5pBBez2Vyc4Yj8leln+3HV9Ibl+Fil4S0NsTfkEc1MskAD+3X+n0G0pF1rzftGpM
ZMF4ToE8xdiOeo9xAKs5GGUtzSbEhCevij3N9cmZhaAFgZrYJ/K34WGwbxOamfg9
NRGLCGvNHEJWHfsIunrrvD3Lz4fdSpfK73XiamFfutw5WIgRnOp2tlvplPGbQ33S
Kv2OOAWBq0SN9iPlhQGqlwAOuVj32+m3TfIKokSBa5hHVt1x7ruHbw1BuNgJ/mcp
7VmYmbfEIazka3gM0DrsIETzxPpzYdcLXF84HHhPnnc3uqAlil4P18Q9hCqwZw80
8QIiY1Y0Rqt5tqK+5bmipiTt1PWFRSmjR/F23ISU8SxFyWG5+XVeNfkaSCWs+AUf
vor38HKJNz0o/evUg/FHArcx/Zs4x6+kvaNahD6WoW+AuoO/+Kf6A6fgUZUX5ZMd
K9cz4/Nj5mekh2TVd8PszJ14KZM+xyGR7AbLUTScr5feh6s2vnTzxWLsPpms9syA
mJ079AkNF5Wz06X68Mj+XVNG+WIP+dx3G0OWmukojxn9ow+LaNvbf+0lGXTD35CS
z0fp/omXyMgr+E1bqLlsN23JA3qAqIesYgl/TbtUJDt1/IsdkW/1iDxp50gV3FwC
fiqggscmsi7O7hj9/3u/SU+2XlSUImbkMUlSPzYHNOnW0q+UWkVGyvslBgWW4cpt
GoBEzT4/u3WqDZ7kToAQ6MWeu/gvtyH7CC7tztYMYHkolNB1SApPkcSqrG7PpXca
/ur0WFR/+AjT9CVrxyaHTxqQuy44BPlBrnLW4x/Sfww/LWN/cJUvCwKyI2DgHM/b
KXGScZYjEuaWkErHTxOH8hkVdRWqEjeCaLg6y7PRUMwGG3qe5Oq03+HcHnbSYkZS
Sg0Lcss36vuCghYFbdhKVvScNnd2VTH0ED+YotlAHEc3JRNKH1wxR7kBkhqdGZXN
4iaN7ZNOn8s7dI3oK6Bw+6pOV0OVFrucEqbReD4gSNGJK5BiX4UAxvxbnjHy+3Ir
kY6qtcaOrK8sq7OLcPyUHJOeX5HlH8PVL/S61DoiLuLLdFwZ6GYSxDerHZs7tZQE
if4lo5CymkjTJRdfwJVwWAROKe2oF6uYSlXAyVGLh3X7AZVUs0kBdAsG3wQnxMKj
en6IQ3daTlsrg0Bc7I2kabqWQjGcRrICbZsTjTIuQISGuwt3aTWi7mSCWhnufXBf
xchLLVytyzgGkUZDIVk6IACXjgp/AMAi5pEWiHl+fsejCvyiEyKFKsY7bF3GTaun
DScw7bR+3ydFA4sjhAbQsq5WtRqwU6gpM6VpXbJS50oIOZ7wXPN9QKyZ1qkOF5Zs
ytD0pnXKsGPCOz0uKouHkrCxPtp8wFz/kbX1gnx3wc4QHmi8vjjp6IjHOb4CycgF
RmUXA+7W6Av58vVQYQVI38X1YMjODl/ez/Xa9mSvksf0m9HskZa3S7b5iB8W5kv3
+mg8JxSuli9+pOs7yWUNHLKqBUmLVZ1HKj70kNBeMVKsLBc/CaXZEHie3Rsn679s
jaOD6UVrQ/QVYgkCD5krKemXIK0EVQ0Xwk9/5umCZGftDMwj5s4CerODhwyeKuQK
Gtw1PaZnwEnGVeaAA8e8Ucg54EV4ZvZammZfuzIcz8qbGuRanmi/jpnFf+yoUtg8
7wU+O/lCe8MeQXX4/s6CPPY6igwNAoe+YeO/c/Eb8255Kv5h5zdiZBsE+ZjidVRL
9xvdCJWSguQED1uVuDwdW4JvxUhHauLYWoE5MzSpc/PqCk1IWICGRVxy5xgijanP
Hf2hSPEnR+uMZV1TyWVonDwpGLlyC5J4ovxgeRZCUxy6O49j++Xn/5JQwgqlirfr
2AegmbYDVYlHu6mbrZDppyrLpq1fSGSdp53ezaXDk/ce2/mCpmu3orB4xm5OGgpg
vM1rwjKL9RQr8mvG+V1x8nAWnax0sek3SlkeSDvAhBAgYfM6jMmIELOcvLOt82VL
wVPvzyoLN3cwmFj5NmLwuaPoOYO9TAxKP9HsRM18fY8JwQRvbMoKJLSwgJvi+FIJ
qn4HK1OgHdY7jZd6nCkyk4y+DK3nVcuzlYc7E/9z/lme1arQ7VXZ1v+kru+wHlG7
FUJl6sCIYrhEx4+VS4467+G//agk4Uwai09MbUYFXVcbF56qo3jqyNogXNjFz59V
0axbfc1/LDkhFAcq6dHZv4HuvSJy4n8Uw6kj19Hf6tjVmcFhc0r5rzZ+sSRaI+jR
b7MI3gDv6J6ysFLJcbQqR8NyJrdm5nqYduOyc8zksWks8O7QLB9coQ/P3E8KWOBG
XuC4dgru23+K3v2KRD7kBaSIe6N/n3DW6yywHN4/iQ6uS/XmkXeiadpV/a1mG3ry
lUlGCE01F45Ip1JxlV8snUp2QLKY6LI47Sk8tfqO4moCo+AOCQY6inyl6NooH9NX
cKHwoqinDm5dXwPggu0lAzwVkp9IyQgsPYSUrrI12TB2jYX+MJw5qikLxKzh0w7n
/F2SKeHYA8wks0J+scJSu/iuV4tchIugufej1zjr/k8OXpQiDx6M224MUiq0GXRH
MjCMH8906DpGUDFDa3IR3RPmTJ6vZjVz8Yj4Yc5K9DTT/r1UBx8KBAgBMYgczlK7
wN+kNBPOuJh4yGK3PCrdWOUbPOqyKDJZ33+LWRWP508a3yFAeoVeTE35luwNH0wS
UJX/3hqWuO/wn1XKBH/lZEhF3/LzVYFEi5vYhtvz6iNepe46jZva/EHw23fugnD2
MuHS96zAfpglSbXWqBM/BnNLquiaxoY2OfHXLtS/7Y9YQTuDUrE4wj2k5hHtyzoC
JDdn0+wiw+8lxisdZhK7GqwiUcvYI9JZl2b7cpUsAlglJH9PA1hnUNSSNIQwtUVQ
J7E27RyIgT4lUTtD6UlLr43VijmIldvcXvdUfYH0d1KHH6EKSnBlHvDyoJp5wIFO
7Ej3EGVmGpeF+XuYgXW0j11R2vgiHUXxigVyxHBo8is1VVLed4bCXqQvBdjbB+wD
V5VuHWQkLfsx1pgYWPGy1KjoZN1Ff+kxwKPmchZ2ZgEy/Jvz8RT4dyrZtqHPqd8G
W0cyI5axhaiJMmipv/I7RqNxljHvsMxsgCe3HXrJ8pEXwplyxxY8eW3Wxc90EoDW
LRJO2QboQWEyx7KdTSvidKUtjucFkq+MKj+Q6qxgaPxf8YhEcDMELjJmVpA2Ql8V
f88gR/9rxoLxr0lKbHsbvOPdxfTlMap03KTgoSaT8Ek9C9iS13Q0nXjR6nKjlotU
lxUEAWdxNQleftmpHZwq9BLEl7uSFEtc/LTs2UWL7gDIlRSxnBFNRZ+1d9mQRcGN
hv3yrDco9Hcq+KVCU8t25lBgdbR3f0O3bL2qgywWay7qEjwnt4xMrvG2SPuZtgwL
s/+Jd4XkXwzADTHtUxD+NRxU73FBXCg0perBMdalxHhAQ1QCN6kZWgIkHM5hnQWz
qfpPtp7LhBAkUtR5QPweTSajOLFLwurc4XNwhEEf4yJmK/baMfWSwydh4B3iyzPW
akyBTnvYer43ZGzzwiWEp2rOin3aTii4r646/tr4ijY01FPC+WfOOSKFIG15wtA7
jiagzK+Yrn2WEE8At/p90sho9vs/YQi0rPgptxlLGyjh8C74FyRB0CmjQ8up+VJQ
gwLnBDpd9wpcu196v4JuL9smHrOgjVnutL6Ck5HAtgD6Uy8eub2u+9Bav6uDS5oj
rIHORSWTFmrXLFqf0EDjbsnYWuH6wE7xeHI6kCYcbshcVLy/IuTTtbTtgi6NakoS
M/fbTK1nfAovTLB++OVRYVpytQlcGoUegjgF0yU2lZfBKb6MCrk9PbJbFLE8GV72
OEGwW+TAdXnrTQ9tlIm+z0S2/eTg/X9SE0E71/eynnvsCvjMVpwkHv+inULW3mHF
UouqCkLLs0CpqaO6FlZA6ceA+Ngry7Ffd02nP9wxXy5GLiL2FxrUR1FQMtL/CyE2
0vuKm/ejfQKqrrHuYsJ0Q5kF3fuQ42bgd5qeVUfiMGl2823M2fmMkkZKphVVMqtG
UgJvNxbaiTW0SF27NbE3eS2zAz5YMCfpBziA7iUZjjALMzGKNUUmvcbDdwqi5sI5
Uldf4Q4d1lUDK365hpjBn9XHebBts2ckuEExPdxBUNuvAUq/2dZkxOWHwCNeZyyG
vXyrEVJhbcL2beNVwCAvz2HxwhgyBbV2G9/UHpOBio9zmaifuLl3sNBtzf1Qk6jZ
oItpkTdwX+jnZM1VnzetqWGlL0yM1HVSonNi7XB6KY/1pO47eKwawDxLukrTY/Vz
nkrNGMBMkSM7PWfg+dyprJAu9erLmc2GsjbGkD+/HYysD6vqqTvosK1elk8l/yqA
OwJREHg2B0hfSaoFGfF0x/wEnEe0bNEVWjsotidmV/vnltKJoScpET/dmLMH29Y7
eVfDbn4l4HLoNaEC2FULzM1dCU9qga+uVl6knc3wdchU6kAb6AcLr2jz2a6fXwJE
r3eVDW11PtUIWdLbNzmrCU+uxbuBwDcJ8gYVh45x4eZBg73vcTOKMaJQF0p40eab
3hsytm5Aq3LhKSdHFvF1MpvD/YIaj5SMKndKSalxM4lacnEFKGhXaVz31e5W374z
N1o26IcJ9rxR+vpBwNJR/sr5jFUjB5csgh4e1BzxFSXDcz9bhyWN6Wst/zvjm55h
ZzuFANhDvV9wc092V9XML50bvnLFrVmiZVtO4GlgEKn2UMHDY5jd2eij1WAYG4md
C7AwSgbv7DzMtTo4hf5+lz89Q2wF7VvYk8ZDLZt0wosklFgQhatkKud9kTh3NAgo
3vpM6CRXTRuCW3YkeZTohgfYYV0N0uQ2u9zlxTRHFnXTVyaM74frYdlGWy8j49hV
LkjHhMMFxI5hQrWQSSlFO/GYhk3AaVK6QZjdo+5EwkOJoyoUIV10BA/G60RhuqZ6
t91vnNp2bVd4olxS6fvMqS75yGHHHRqjDHBqKmIcYnvLXFZpTqUSLEfjpGfeaf77
XP6HsqkZoJgPMrr0oPcvigcJSzJTX65ZJFXcI0bffUH9apFFNAwGRItPuTmFUDsf
nVQ18uNQhR3532b5OTyLZLg5VkSUjE07dzxRmn0WYTrxldBvUXRdxHqgmuQHOiZG
SoaCZ9sflEl6yzHFK/MSpWjk3AGIaZ/+Bq09pxjpGfB94cxCt/bOE5tR7cn/PS0N
D/0Sja2db1C8l16s/k7C2m8IqIua6i+DW+YUhbkMzSxEBXuAtLfBHrzZjltJcSJ6
oX5IngpQAAyMs+Vk9Dw3JflXC4EL9KZkfh5fg7XvcPzpo66KI9M3/f0ND3gbeS1N
pWjLhi3ps6PBmtZDWqwFRq0tS1w2gTEtN5w6BYuCiRLvE4AJT4+sRh2IlimpMxyu
mhEuYmDiIUkwKuFN91eECpRJokQ+FFw1WcbFGu4fBT9d7i9hZTM61gfyyRp6VmZB
82eYUpY48M/4TfGSJx9XmuUXckz7l5Of2qzIi5lcmk8q34icbqtHHcMIV/N2nZCF
kj9cUt3vwKTSvqjuqUiGXytJ2XevYTC6OeKcGI7zN+2JPMFY1tFIFBD9QWjerBxL
izzLHTnMg/0wVjw653Lj6v41mgc9T+++rtlKlgf9EH9Xue+n942yFluR40EZr3OI
CG2MhmZrnrkPHTGCgaYogH5gnPjYuajNTj33203Kpsob4ENOwsgjJDKrMKXpnxq1
P5AHxUwo6kURRltqK44nAhAxxX5ji9cHdhf7F9a4eM5QxCH3E8NtWqDp0Mb2CzGJ
3IEjrDN4BHH5u7cPGPOZvZLTYcbSi+UzdMYDuCHaPloOZIuZv7mk94Vara1s4bcz
tsCnJMJzrAK9Sr9vLJOygLHdzRtQg2wT03xzy4JOdid6rYZYEO+MRqai1Q+qECci
cbuywZsbAuUa7CnWDbdyc4AUti7GpVlUa4hkeP+iwW7k31enH/ODC8iVOPH9t89b
BW5NxRES8thS71ZsSntXrHZ1o+YsfEJPafDbh50dOdNejb+f2+l4xogFrimdh3eb
ylgECnWpznBMzTFJ4ZB8DYFhtuK54F+HGVnsGuwv0RZuIWUW21vCk9cH4oRPeWYs
/zXOpQwP7viJ5vUPxqPIucroZ1hbxAt4XukLmOQ3ptskjZPD80rjiOCnFE2xNcun
jr49Iv8o5jao5uy7hKJUGjIYoPTvwkB51yEYR8NhGFaW6KtfvCNQmC4c0EXp5zhJ
wRRiGmFSFICbFZRmcAUgTswqZ9hqn9QSTCV0FD1c+0Ycfs7bZjrN9WLZZ9brlDuy
sEhQwi9hoTh5sZ4aPfdet/yrNVJIU6VuG4m7I2ORSjxFLy46c77xnQRJHON7iisW
mjN0M3dye83l7rxSZZ9KaZev4kQbGYu+/tdFGx/IiDQH5TgYQqVZNnZDeN+JpZu1
+cdNh7azcokARalPqr2sw1rhKeX3va1I4qOXl6c/zh5q7CAkPLXWKXPJ3UJO2Jw+
GiQr8dCGghehYVsfXrWoISVlD6nFguK10pNCxGKkZqDayQuD46w9IWr8yxFf8UsP
8hIaIxMU03SNG2K10/lMfYAaEG4Y4ECew5XLORxe7S5zmh6DVtHdUiTudiIWiGF5
qSq/1J/VXQ8Z+TO6JgUAe15Wqxdg4KSQPzyjOpwd2ZEQr8lka9r8thZBsQBTacTe
Vi2DnlpHkIKt31Hpn8493dvhDNAp+2PhzXmAcdysb2ZhwOn9+iPAOQxLVaC8NAxI
o/w6L3cyOBSbXtmoxbYfS+p2YTWOO8PW6oXnIDJYTXuMUwXGAcpF6vmVcowukLKg
/Z3bGaEYZzqerSfIcS+pBxOkr++HuujX9t3REm9nDsN50ywQq14DgEegTG5CNcf7
uxzoIW1I8xdmv/QBfAEUBaWFvBTJZUM2XQl4bfpd2/qDdJyLCJp492Cr8O3v2jSo
mzkC9cHl0hYo9a+lx+ctAD+wZSp87KW//yijJA7k+hrdn0EEMHX9d7thLQQiso35
mopu3jaP56VeJEcyYHP6BlILA4VUdKo/vTsxbgTJHJeYAnXxxURUfcBoyStYDOO5
J4yIrF90qrljgsw5w51G9uHeDsjd9m/zMa56FJX/ltz9sh4Q4Mn9ZjFz7hk0CLE7
tgPR0j7hVi59jvWDf1IVNNwxfIabaXHvS0iojIv83uZfW0VUBCsCx9rJ38JtOjvK
8+Zj0+/6/yNHweqPKOr9lAdZtF4RuxR4bRkmWx4ffxF/iKF8yZbGqbjvth8t2BQW
78Z2duWLziFYS7WN8q4PviZNdJQK9MpQpjDPN+Tn9l4taK5JoZdS7ve5uBvbP87p
e6Moo8dTDhwhl/csyt+U26csVPaX0DRrx7nVmCyYuS3zwGKPnuYWsC0KtcJpK1O2
7REA1AMAtwDyPdGUHtL9ieDntx9KULC52rUT9lI2jnOD6D3lK929sgN9Oc0IwXr8
ArvxUz8FeWOz6RnhZxfgv7GvIUYe63fdBdLX3Yy7eUdkLCiYrJXol5LSKBaRf6ve
dOEjQL8yklgba5olJrbgrvy9BrN0pgbRAtzu1IE5C6cmursMTtibQaWcL9jmpJFp
VI7Is6gm2cWcwtSlVUjVF0P4LUEPEW7TMZTeRyR9BAzZFZvf1s0MNN4VTgnOT77H
ZA55+JkQSErIoKVl0KnyALDLSDbhV8g9WpEgOsbgTczv7bvw+Psw4NiOzwlrLypC
pqDAa23pgCK2LP4yYznWYnIqS3MHONBKX7I4f5PHrj8qZ84dLJ6eP39UnFhAwGBl
Fz3wrNcZ6w5WReAigum0qa9cWtWMZj2GxNQaJTi+oy9WZhAwjRm4yTfMZFPhNt7H
bNuZqa3IYtn929wLnqW7k589VN9rUp09Iu1MZDI7a70UK1JNYRyCHdOkh3HHFxzn
m/ONvuUyJlIk8WRXT/4NvwJTeqfKbNJpLJF8PzNOdYE4Ig9YrD+r1RHv221qtosF
oM7RKffCk8a/qW9hz1Beg/yEhq96SbnXTFtvzugxGBduE3Ja7qIYanTSOopaC50A
oKuOjcmmf+iPqcE++jY/KoCX79zWmBVAFYZ961e26coHPdhcuDHTwc+WpSK6EdHo
BSo9vQp7PDk1s+BV7YjavSjsJcWDatIcvIy/tWfUEaV+qNn/hiuhWflC49N6fqRS
JDMZeCGYTD2yAC94ViW2zo5ZHo1aDxdwRcLOWsULavIjdrkH1voSRNS/wc9ZRoF0
DfF46liFX1C7XbaE3OSAPvKuyLbXblsq2NHFNQgyNczVoWD5JaCmXmTp8Ql2qu2x
j6dVgTl1vcvkL/YX9HWqCtfodxYloDaHuxHzOoIZWfXsh8sJUorWVjqZJn3tWfqm
TWQP7MH1rt79awLb5mTSWz1C11Aa+ZXucLv0RDVnZkOUb/+Zk0UfMpL92UAHWUuK
Tnjr5J/AH6HRunYb9qq3up3XAkpT6FTB/ang9qFPegMQBBIiVL5NxP/jTbVvjOhC
JoMFD6Rd9QSiEt2PoOc/vT1b50TIVi0+wxDfxzcx+iO/Huadk6itD3YWcdDHDAoH
H022I9ntZaWp7I+yJ/sOqrOEYsCi9WzGv5GHURbwEzdigv3UvjYfUK1UR+yy6Gz3
FWljjZzWlVlvMj5Q0bvrJHaLFEqhqZbdpMUq4/iTNJgxkKm0hSFxLXJDWPQI4/RA
J1iMy4pfxjOD7inbmUmA1O/FTBpB2uW+9YRbV64+qwOR6/1vGLrBjpld7C7t/pxs
so3Bfs+KcGCQWfZEFrZpTCjzbaGP0E3qnEh0u9Ds1GQwgDDENK1c0bhkMShQbjzY
WmsqiUbfTKdYO+SXulzfbEFH0dslqIAWwNELuy2xk4aeMpe2DiA1EgtYGyU1kni6
MEDFs1SYFUmPO1epfmXMNlqx+SmbOwfkpsp7hed36Sn8dENdNRYJbhr0QtnxIabH
3ujjUSIupDelpZrzJnjBUepRZ1+aXq7osY9N81BAWI92O76EtWxzGrAoD4cpnKjz
5HH7V2HGXPbeaMLjx29ca/tCwQY+CTxOtl7WZ813cuYz964LdLjiM3xxzH1cyvzh
prtey6VAAzjaoAXxhZvFkf1JDU3GIuOl8JQlR+tP+mqGF7r6rqFYkDcIa3oDvlGz
Wx4ghTEi6NNNsNjrMZcje+WNfJV5YAbv57S9JbzUguxCIr9uO/rhf3k677a/HcTx
7wjgTlW0dgeAHt7E2q0R8HO7lJa3FKjdKbKWLmMivVEFok6Cf1mVYcvDXUU9CUGJ
enUcvFP+zsRXS3QCp1yEHqmHvWHKSa4VjS769SOr/VOFNvLkt4RMWQesYWfQXArB
F3lSdITaKFFA2NQ0UuBlrEmpbbV3TDCmXXzmDIk1Kkej1PzkIZbaJZ7mwPsFwaZe
yj+HPbxWLimn5tlZhwOMXdXrbRsC3jynY61HGbIX3EMFweGgOID2tYqn4NpMY6mI
jvc3DHnjal2h1cq2lT3qIehz0MGMiTnUUz5cJdStxOOetdPyBcfUclmH9J7ogVYN
UTbuoGV32y9f29QbvRir9AheF9wbOo0IoKJSLHvmWsgimrmFytdHLLidtWGikHU6
98+4W7zdp5udET52D8xAl6QsF2pKCR8IS2y2x9nrb1myhp2ZuLuXJEImExNaMieq
PCKo+K+5YjGKFVPLglC5yLZ05BA8WFDQD1+sWUJmVUVBXZ2bRLZjUKkTC1inY+7r
nSxZwoTvzxd0t7xGh66wda9Lmv9PhAEgLyJQ3iGXw03BN41bVtGCjTke7aXzNrzE
5pkckAIZI/nKMgVNXLFqXYncUSaOTNgdBVmeMNUTo8RF2A8cu01+spTvPdekAnQv
sFuj5GfejbZCmTCwZ9raQ7faVKe49xKAhfz3gJoCLkGLUVTSCK0ngO8nZgOqS7m2
d8dRd+VvynMw6CfUijjmXEjg7zkiSdvh/7UobBHxkbgkXEfVV0iZTwaoMmX1AF69
P2aKYX+zjfvQ7Q0/5UXjgi+noXGQlZbTmJ6dzFshWOF0hfX5QCXqf7PptSaqtdns
VWDoYtR/XElkZ25QMDxG8vp7AVuIcbrjMWKvyp0EUjFNRVV7n+KE2FSKaljqTDmW
aKdN6+DaAxLugTw0sgri6+w4CfDHpIdaKw296nvbe/KZHQ0k7ip/VGgmpBMe3VWZ
+zd5h5vU3uEhTT+1GuyeBx2OERNzn8TEk4r0n5GokTJTuEZ5659rGjqWrIiNtnL1
F1ihV34rPYc39eHKYMgEnRRfjYyXxB6qrXZWiVawbCY+JeSpjulFiLeUo/Y2LlWu
TxOtfPSOFfAtTPlvLDKHRwnzwUF4ZEurSkRPLIzcHSEy7hVMqFYzuZG+MP4ootlC
F8oWLhO7Xc90RzuZxpf4X540wr5J9zgtJYM9SOsrXViUEAmcNiWHo2MTexj0UgaW
IK0heQxNEj2ig8A3sRYDHGQaaNt4kocI2XtpGQAlXfmhJAzcGL1celuVFxLEOZhy
xNxwZg/0R80PqrslK13di0UbFvTNZHPphVIpFdG9njmPD8HnMeAyz/mMBgyZdIEQ
eAg0m+Rux9SyCcI9N23e8lCDajXG8w7fiwoSGHuUqZgH85NdLPzkqG8mgf9pPhut
yfj647Wscai90lNcX9uXQpApk1yi5lF4jB53k/YOQz37hc3Ini1Jcf2SQEdZksCS
YQLnaI/1YBBvkcFKqyyNkDITL0950WWZGG6zkbF/jN6N8eSa8Nu1nqQGqgBQCvtE
mm3rQ3MRwVAYB8oPmfNGelib7NmklmzXUOWdfQp4yms6nrXO3mBP4rWjvpPkpOb/
d3xXK1C+lNwMKgUsnW1qIiIcxFhgtQOLc33sKwN3VhIPhJhdXNk4yBhIUCm/5SPD
SNqOU7vXvWcX0B5APSBgkfXCBKzrNgQaU5HvPjTCTYULf7bKZ9zD6VUhUjinzIBI
27qIDvKfI9jkmBsBtvneAl5Zozu2WNp5crDWhNu14rM6JI5JzAPHdreSzhJWDolZ
Ly/nKwl0h5a+M7nRLlLlv3fjoN5aniQi5iq/1NmdWej/XvgGPJbQNNyeBB55mlhR
Y/FHsjpYhHNC1vMi41J9E6+Dh54D5SpSW8ZjeAlbZIYjoq0XtSE5kGT5Z0YLldT7
14wARSDWpq/gla13Ui5m9TCeR2aLQXm+4uLAdiCSQUAdj7Pd0l2AgIAzTdY0LOis
a/I5IStA0d0BPP+2GGzj6Bv0YFkZ6cyUAsDVqHaA40c+4oaDgmbDNM66vFQJHquS
HW0bVRD2kSSE8GlVRUtEnO2im3bZh44CVyiKLfbn6sI/Tyz1UF5pQlvYONQyp+/C
WuZ70YJXPkxcVeJLQ9LFfQ94D4ED7kz8azWp61JKAP3n6QYTPnaWy0puJp6lzFlm
xtcFMAE4Q5EFkyPjJPmWcd6ZYgFZbMxHrIvbPVx+n6nMJ6qHziKgVCfxDIAP/BPc
QYRRoN0RuDwmFGWFJVucSSFxWfcAEilu1F8+2kOwvTl6D4gfncC9UBl0yXENNjd8
Ju70mmIHAh6enKXygHf1hxDOZgzMlthTtS9BbASRo5jTtVa1R9lcYigRkpTmK/U2
amNfxduJyuzwdFKO0OGw3GeWurg/DHFsPXR7kwJvR2b1CdZdAa8zzJ7RChLAuyRW
KPyhcRx179E8Z3f6PR+LB5iL4f0f2USZz4r5flQULZrfYJr5X1tKUnrdP1q1Wjsa
YTnWOQVzkWFPQ+dYviwi0lJ7VbFcspJFemn0z0Z+ky5mpH92t+mO/9I145lQMZgq
Kis5cqnSg0wEVk3PLo5OyiJVHfqeutWtxEYRyyn3sMp7L+odAQ6AtwNcMICfjXcT
cqTNDnO1WweG7imgNqFHGfacjNWnRHtq6YgeYG6IQ0Dln7UF/PyVnkZZuw6RymTf
0EBOVjB82mD3sPN+4dSKdkyJ1zqK1CCQ6IvoekikebtKG0UmhvrLY3s/kv2xRrtw
7UiUk/8DLd9VjSdHh9Ixnt4YhBifRUHEcWPd1YB6FYlXleWnBjUC9xwfIZO45GI/
B27ARpppRTesrpMKLZmjsiic612G0Zrwbv/9ms10zN/K/y8A1F2Lqu9DOqqx7hCW
/N2GqSSo2pXdF8VidMmIXWdXAy2kgxyf5/xSv9cM7FjwPCf1pImsfdPY+lsve09X
Gn4q++ucuwddzOgpMLnKT2W1qvfSkfS/W+EFu6d3/Lywk9nr7cJQYLD18w/+qMQT
HbqDigNpdHyix2JiLd72crTcPEmj/K7dw4jbDLJ7PW6Tq+FmOKGcq7lLskuwzWc+
VSMZM9+vTiyRDJAC/dT36uv2Qj43LN+rQ9oLA/66MJ5uw7RrxItXVg9qMjVMquKj
7dQ6ylr5NQM3Jc8XgqWcwI9ktHeJ0FYGxx00yvvvDykvTB8Phf2GohE9Nhj8063l
6z+V6a5ZSj3+Auabyg5ainFDG94qW+EKGMgwuTZOhxVB6SD7/TCX7rlTZzL89n92
FtZQeF3k5Hib85NAyKY69UY3ZJG19d2P6yg8wzsBjR7n4xRMd1YQAb9yj3XrJZ6r
tdrv0eqcbKEMH6zafNuu0vJCgt7Fzfel4bVMtFlIBTCzGBI5LE4LwsTSJYfDJ67J
NBwV2JAhr+sUaaQSKEnmprl5JEwC8cGGIHjf8PzwrMhB6HSldJzML2zt8kNZ64XG
E5k/GiH6qY2CESC4NBu97fFgulRSF+DuqPxUD+EvrzDFF1WgMVLOOCeZlp1cU7Nu
NWAnoTcvYWiYqy9pKyfbIqYx4uSI1E2IBMMg5+CPivI2IJzYI5ElXxfDvKN245TD
tMcl+VLoatPkqYN2I+gjkIMkfFRVeOSY/i7daMuPZztyoCojikGRJE8dASKlHBL8
PCXQqDM9bWFYvzh0p2Y+A+m+7fTf651RLmbgT9T8HSs6i8u067h5m2d2X1lZOFpx
i9oPmEHZl1/eU72KQ6gP6nsa46tba+O7armQ8O8MzgRa+ZMk99dbJc0r6jekKRrn
d5E/crJ2QHfEqXWK5Iu8QWSl+CfcwGsZXhc0A+bCKUborcq2tfv7pjQWaSG1bQ0o
svAgg/g6kvwUC3e7WFwiZL7A6dZlvDKVsVlyyCnWuDdvScybU0oshoq1WSV/ly+t
s9tBcpmAqOCF4giY8LWvpgDw6kv+JlgHphQwo3PK319V6GGK5Sou33sCZURQZRS0
GlZZtwc0mIhSV14PRq0dhiU7btgoKjTrIW2owwuczgJToktr1agLU2kKInWQdTkO
9r2KBQdBYfuDfPbqlXTYGbRUdqPgs2xi8JUfdiu65nW3IYZ9UfnCI368j8t1MPUB
9mQM4I7ZDhO5tr5a7Z+GstVQz8SyCQts9ymxoKaQOt9cEFDoI+XkJZDYrUNKT+NE
SX66ueo8iKlcrusR0/gFIOWNbDMTfQCkKsssDtb1Rjdee3fhd5XQvctbJ/ShdQb8
7yUX3euo+WIeg8RWYHo+VlLqIancNhbThfKLS/353IYGnu43ur19GM4QJB7cm1Bs
YRpyF3iqXNzAh3/QSZZOaEbOL1ce9NW9XgvDhcYMBVwVUa1M4ttBOzVMJnrKBEyE
0tNX8J/5BxDibV755FYRpLvSkt3AQYFFlIS+QoVEKijLCaavbdF8cYsNCCb3oKLj
fZTMZsvjb4EEUtSppziJm3oMb8Lop9geKzFHMJ+R55u7Xdv+SRYW0gJm2dQWmEes
59QBIvRgXbjAtXmOCvBDqkvalil2YOwKpcmRIO+IlgKIcdoywsx1irDA2300VXl2
5KweF/vTF4Pmqk0iwH6oIEi6RgJsjpTysknyNsR0Iyi7pa4svP7Zmmema/3PH5M8
yndon0vHTFLjuTfV/EgPDHK892RgZWycuYPwqcbv4FjhG5B3iDsu4JOV8amyb/Ha
ow2dF+U1bDnWbEHI/ThZwKx+h5dFgy2WC/Cc8X8buJiNuJn/yFfJVCGTuP6SFyFP
MLK4H0rgxBKRcSGJZIxxQZPcKDkSql8bWzcgQ5o1jjitoFP92V79s5MBBWnTYjiI
6bXzg/Zs7bUDXHYZ3aWbCGORWhLyAMU9Sm3sFJkhoVcdj5ooIZsfFOLXa+sldw76
yIgE/6qaCNl3t75YutFCJeMLsH1UCwiiTn/dcLejMnDzFAucRobpEmX69uF826ea
9OJXMOiMEhdQVr4D3Z4Y3eDP5FiQy7C2A7DnD3+C4EYCIpTC86++KYU9ZjdknW6S
v/nVJ3BRkeJHzLz5LIFcMX2dpMPYSOKcB8y9M1fPHTFG2Ha/p85KFa3PFF430oX2
Mq5nNyP4HYRfAUQFkOzQgXPWkgkXLz+TDrJ8MpoyMdz9KTYL0gsqvI8pLfaYOP7y
97SlHaZ7sesMwq20S2lNTQ9r6lxbryhE2RbW7GGz9wy11t15JoOyzrrVKk+NJ55f
yTJ/CD8FgI/kgqFThbfVSN3/uTT+gQFbDEjeXUZ54P0j/9Re2ZfLM6dzC+epYTPN
VWf4UoxWhlO5v9m519QjA98SOprEYkzfTURFUuPZ5dsclpmVqMKzBYSigTbJmvkP
XoT6gT7Q3/HSeQMAPl3IK7NsgbCkQ2zfMLwtCrBnZqh7EfNHdpnrE8YyCgICwwSp
EaUFlpUftruE5NFTZN3fvB1jNh5QYt0vaUm0uMua48MXJS1ZApLYXKxot9sdaV/m
kdqtdQikBVpCvzvi18phhduYzadyzdW4Ix4VOoDrr8Cjul2gvpCgk6q8FevmQlsc
IDWg8N5Iid/NiPDWeEriOHfjV3DZg2DeXmNW/sJRiUDV4ERZiX0XfUs4W0MtNQQ0
C4VvsEKt3mWDpPnveaquyIT8JXlJffbnz6h5DzsWv8Ic8Q63sL3Xx92V1zPn104v
9GyBBMjTKKttY494qgNT1hw/zjAtdX32oyfizZbCBtApA2BQNJMVqEf7AZHaSaUZ
0LmfILWvt3ImdleCL4Q3gVaG9cORMlxsd3w2koVFRpFNWqaaqsCNDiWBGnN9oNsm
giCwh83AmC/8507DzOUaArtas4ji7U+AS5skexCy5kW0VzTdfOhjeRISv9s0FfiJ
n1r7lTi9ChNz3WwYxnxOG/Pb8K2WOpZDU6uAUVqhZqspM03f+UGiMSKXg3DTQdMw
+xfjF46UusvFMO2k5z/tty/kX3ZoeUg9DCFv+wHOLDaNVDMUTSNpvNtmzrHFCyXd
0bE7LuwJ0VbA0G08SfIS8OkoNXLitryKctFS0w7baHHm73nke3u40JF/wuEjro1P
vuXGwVpdyL4ad7ksU1ypvZ7plo7IBoAf9j8mKn2OyrVEHHdmFLwTt7UxuxJ2HPTg
/569S4t7GOoCngRxYVL1a5jt/Rmb/Gpmv4i2JPTCLrgiELgoyK/gU1eInymY/fhY
bH5mpaerTC0oXx8yGFI4rtSNOtgO9fiJRM4Ja/jIQoiBFzSMbsNZ+Dxitl2xZHWk
BL0l2fy2ldmbD3v7e+pME3ca9+Te7mtWO7Tc56tVmFG9BxJEtCFBsxgNcaHj+BDR
y999rJ4IDU2WhvXjuizy3Hb22YPaMkvcCWYD7tEEzlc5lIHIjt5401mtZf7fzStp
R4GM2bkraSs9E79LQrS3qSgPiNXST3FXjTsyLn7c7Cs7umdmENEN2XYytyWKZY2d
NiCD7/tWmzBzjH0BvohdxNRJcyrbb31voAHN+suYNXDk6o7zyPv7oVg8VkTiTPeq
DGxbNO/X5XC5/qFR2v4g9GSws5ssHgdHt1s9SCqUrp4wK3WDC098n8sGLNGQ0ki2
hUkonc9icAJGQ36AJopQ7XnlvpedFQKzvL83mDbaS+Ih1ZTi8k/Gvwe9eooINh7Q
QnhgNy+0JJin4DmJ7I8Sh55rQnjs1IRiYaQEpd3T+eoYxIkqws7PaE0E96fmU5VZ
WKPBl28ni9QSkA9xTRJUicBlS7/vxA9LZahek8MneFN6IeI++l2/qdpAG7Jjg01t
PC+cKSlpyOrvRYn7QOzJmh5RnWNVEnx78938434PyUnBCpMkBrrI8eNpbbt1IDRo
Fk4NpqV3T2fRyQytVPHJ3O6Fa5MKdvSfYh0QXbY19BuK1uREhhgUYP9gVAiJMq6o
WIGW2D6DmEhfMP6OV8poxd9rav0/RcrnoMkl2r9+hQmGoJ0z9sWmpvrN/2F5OcSG
EaJCB5p98glrvEQLo0+5uzsUNMbxnfQPdYRwVJbQSYe7UyraZydjKz4ojNlEkmG3
30/zY1XlbvcBGkZKwnNlUU6BjaAphsaSbqexoHpVGwTojLnDldfF0b4L9CFBKFn0
0cqj5KfYfCKHzgOhRyoDCR/HU+dNNnd6d8pQVi2/0YV0IZdyotgNqLhPuCn7xzcW
qOME2bxl3uZ03DadfqqWfY0v3Xw7wmDXa1P7u7PN5peFEap2PtgCMwrQaiHmxe42
sRPQW0Y1g9T/QuWXk+tD6RKca1ORgoNwXcL7qPOgmubz/5LgqRlRUdzWA1rivWfo
5BfhNIjakatgZVayskjPNL+JutzF4FR1Rhi5cMNV4CuR8kbcWsx0mHQH67inL8/+
EGzYUg0rl5huFL7GuHY2HTDG4Bclcnwvok+cYGbXqCYycjtXzMsfdzBFAcUaxJDJ
xSqxsSpGgzjgJQ8QDx1d7k0mXvHDhe2NOUfOrZc540u+IJg/YG8Ammd52h/+rE2m
XO2GYaF+RJgwYoy1S5Sh1W3QcqtGqIvr/csaGG1uN7C/+1zT+dlhxMeI5/Z7MbDb
ry2QJGXAdXxtgitQNCnOEf9ckX/qdXpfyv4qADJoLCO/Ma15v/k022dL+m6ekz2S
HzIyoiAivfsvMYj/TwSK/7if+BzQ9WMmWCu+VDfen8WWPUGO6Q9DLuRJ8Y0RpNyp
ev6nQMubuY2bFOt7n8CoAwCuKQ9yQkVXN4pI/veA385S3fsfM9w2u5B5k1I7ng78
otILsAbtQb/hVUgvLonvhc8UIUv7NWQDb4JUudvys62FCSNP1JJY+tzEl4gqPcmt
g8xXFyhctnE1hnTq3gHp9OpJEX6BxOBb6XFNr+6SIXVCcyLJ4vog0gjEquClW2EK
TEZ+8sJ/33hBrEVo6ZxMlu6K3HA/5xvI6l3GkytT0G/oB9e86CX4FvwFZldKZOI2
+kTVVacIvUv0hs4egCPZtzSAwk5XDZQ8Uf2FcE28uQS0Zn8bKHMx+BUmhQ1jykgv
JXVyZTwMUb+r/PH45vM3hVf0uWAIoLyqBMPYX+2fWZy/jGw10FyX3pVin9OoXp2W
15g9sPOPBqD/MugGUBZqvF8dYw7Xfrn+yCMYVS/oZTnPmhxUX/0D0XvXso5cg27G
nupMFdaU66UFWHX1rtqQxujkwuxOZlNhH+mLuowu1px2gevPuiglCEfN2aM5i+xz
9n/crOV235FP47acHHxbk49b4jxj2jArt5pfSoo9YPAzLH8M2+OBfVbqDLlnwWBn
qBKnGwSc9fVgLD6UKLzqhAq/i5OxUqKA319XCA9+ui6vAuhz+7e5hA1FyHHBUGb9
ijs6xFEpINpl9vLMpUcp6snNXBiH3qVFvO1P2XWmCBCG3cENJgFedOTDdqRD1GsH
Ch7b4L5zywLqilF1gtgjXNjN5Tsa478cKbd1Skm9JjRy/lzKvD5thc4aohJ4psqz
E3hX3f+W3jRIURPDx/3/egUQ0r3V+DKgOQ/2scIGFqCraHFOATW9Or6XdgScACgV
joos/NpYe4F1cdkxewqifSZ3br7zmCLz+Lt0M/gzn1AIi1oi8jfsy/Xy1bBbuNXf
g4mRc20inZki7MJJ3VdS6x7G1gkNZCAZ9ZLQKZyPCO7ZN7tnzOJqKcuU61hguUzH
/+HrnAA+lIiRgI1ZVa6kAMjqijnGcetViWOd+GT32lUjd1mqY9xu0jXvDm/pwc03
kMCT8thPkMnVzuZOXlARVYObeNOVrNnQvoMc3E6fSSt3seMciAbJrSNSbdGA+3yC
3F21Jw5AzpjpSS93d/GgLO2rbYreE4/1EFa/3954I9mWlwQ3NSx5o5+SeTr7yfVz
04vp/yU8mXC2QsCklOtYrHlA0DXbgl4i6QFJF20hYBGrC16AlgQG7Za98CtCnrSe
JT9Upll4TJh/0owbEi+jPmxiO2Kp7QlhhHzKOjDmc7/PySUjpbYYN3hgYn7v8b6J
MdAjj7E8+jj7GXk4olUhchrbJaYtIzY4n8vhbIrgGECuINIbNeZ5vR4B81uXWpj/
LUtnyPBWwASpreJvLR/fyYhPBtT9vcHGPy+FZrEo2B36N8blYUn13jKxUTZ4Qk8b
RgNYhIQWxxLTxonAw3FQqha5j4DT5uVoN+D+ceItLZ+BYk7+bOc3Ux+SAQyp/x8M
4YzSfX0fO/TDL1LbRJ57dYj6PXV6vwEEbt4xXhNNgam+goeq1dbcdWY5t/349jd8
Ybng50PdZAH5bK4J8nr4cvsewk16Kh02bx2nC3N4UB8/MB2HkDhV4yJPWtwrG4ZY
xg2v9yGX+Lh3+86ULw8ESEfKR9lnbWCItYBPjki1O5TJild5UBKkI66UAS9Ot8XQ
xY+omHIigFSAXB9FYpBmkPaJQZdeUoiyBveg1eopK8CwOO/Ar3+MadHLb8a30ZuR
QkHNtXvAbMIM9JzYrECtofcAechUqVWe/6a551/eFkYyS29aLvKsvtMFbbOiPAQq
7T1yZgyd62TELKTsMAwE3ifV6Xj9j5RN8IvvWzvNOzMFuzz0kENwak/S+b8Z/Q4r
z/y0SU8q4wRXxb1lV5kFis/PJaD4RQkWVd4CChk0m6R4iVOIKdvlSqqv+OYpnIF/
h9H4dFjiBHQPc5IWzDcQeHe/FzhGtJBqykqhSPsd0eZsriKP7z89DKgfutd9DxET
FwAIoetHT+AXpxE7708WufvEZJfllTtVRtXvgx6cWDSEs/02zPGIRfRWTriHdnKs
uzhDkEI1P31wnJcGV7p1WNVl72y+MGRedDNQxrdUt1t/WJOV4ULtWBg+HD4v7maO
IQ/LbY8lz306OGcvezatH0kngQaPj/lqlbY/fyEm1DcCuDJXsXxmz8dPF7ariThm
Ew3QmT2SI35lY0yF/8NCCcSZCXlgZyPUGu7ZIFgUCM6BDOPvlBCHQe2CTnj9tf1q
DJM3Sglwu25cPy1kTcdgeMJu3rNG19biul+/JKcH4+W/oSEDZ+fpspWwj/ZILiDD
U2OwNHDVXYacdCRWTsZXYzCQOztOZ/DDqGYuaLIhSWp+d4jboINxJWn0NAEw2HO3
1d6sFC5NoRktUOKwBkJm8O3975B5ZVury1PU0KuBPAPG9HmAL64aErxnqmC6Ls2P
2UaQdW3arCW4oIW1nhOvJnQDSWTGwXBX5Cz0anR1GkMMwuqO/3bjwZ+8GSnZ9Us5
FJkJS1zd9iqowB+sXV9hxM+4C/P213OVEMeOq8Y2Dj3f32LZKeNIuHn/ZHIn6Dbq
6Dodi48qHHDtTNwN2XEsa+qrEs+OZYzUXHchmnFWE3VLIgEdlZIgxZ00+ADRExaQ
I1zm6MigBcb2kX56CeV2NgbQM1i3Aa5b5U1K8FMpdJhRD/YJIfaW2QIvCuRjQnj2
gFnGiIBOGRtFg8WvkYPtJi/0CkGEi0kP1WcZRokpvW8sOe7w4AzY0j01ACDp3ukT
NidiQx8S+Jcoo0/ySAqicknUGKTtywANPlybGYcYuAWqp4JYH4Nj3VAdBlv3OEPw
Hx1o9d2QWD4klbed/mo/tpZR2w9cLFmveRRGqZCcg4erqx0PfEOnO+yTecXokgyA
2b9p34dX3mbrUinw5oS52r3LlOM5uREwibr7FERCey1WXjHwZVhcxcNFd01zP/5M
8SxrT3ib41Ws2xaCTiQe4kxJrNF0n/s06ssTqpxzR2fMsRC44ISyr8xhpfaoNZPj
soTKJYyW+rvtx5mKsF4dWUbHSTeAZOL7SgF8E6Z4lp22ubEwY7gOwNGXEozZ2hJ2
2n3nTSFmFqLL7a3zNBCMXxmxUxStIyh/AFJ7msSi2ghEXvX80aIVUPhYoFpjWhkZ
ks4ts+35ys0vAxVSa5KZVEeLrpDEFg7v/cGqSylutp7I4ya3VGby1znZOtUyStE0
/wp970T7Nnd1tdicHeMmZvAg86nbyrgmA3kjQmDRosCedeOoNhaIWS5y3p2JobiU
qIxBNpUJvSGXzK7cD9x5vgMunXHdxljLWuIRkI3Kkv9dAErmJO0xi1BM/Bp/zyIR
OmAfSsBplBewoOD/YRVCNgrMxEKkkvx8j9dyapvsMZfur1qyEohbVxe9G+xXMnxc
40yFL0vFfxewOLl/OTYogXw8o2JuchXu1ZrmQDTnzfTlUUKnOg4Yz2oVevYEABHY
W++z+G4iDHYKN+yU5UaZOs95jd7xTYVsG90m0qbvRlgNiV+LWi3QjWoVc1hc278b
qOyPnOU1bn1Sx9P4a5c0n/42S5U2yUvRUm25Vjz5OGsuNZw0v98OOtCUMBhqPPk1
A0249aGErPqbU4D3cTOiRbC1GTQ7tH3B6/PiDzzDgJogdoGl+cHf6ASZMhbGpUYP
TsXzU5CpOJNt8iwILEqf2G15UttEm8tK/yIOJADBhhISJFBQcyxO335dhrT6zsor
kx8T92H3zEIcNnWhLXakSU78i0FeigbrBl/+zxpOqNE18iIOjqZfFLMQPR2Aqrg8
k0TsrIlBfNkK1IpgXwtMTayE/ynSOhY1cib/h6gNToeYJWMHUGur1NzyOsNaTN8M
CGXLr96KQhtWAUq/0KB2ssXSuTSBflftnl5+yuHy+qLT5crDujhDOO5+Nyfa5re+
OptfiddFQneAMz/MIe6JSkXbXVHdWjNP5A+qquakcuqLWBV7qnqTM9AOxEbX1V7b
oJaRhxfjaVzVRtKuxIRvWBj3nbYcT62koOjEBaIAiLMKo4MCvSFQaR1jLVZJqbo1
5V6Cvf9FAp5wTqbjCCYwjhJ3m8yO6Lut+V5ntfWjSPbz8UhFbBGwCNxDVExm0i4s
XMEVaFnoUZ7dN3NlIqsOAblaDKUutml3KC/3HCYEMGPSP2rKuSi9NwcfXlyiM1nw
S+3vBDegzsuuWumUfnWtXDSLUWbMOvD78IvRchbcHmX+t+DqTJrmeKNZCOgp4gED
5OYSGSUSB+42AHJPxXgZgypuQT5kY2Dm//AH6bDQAhYghzYupQ98d0asqYAyvw47
zTgmYHrYqBq4ZNVoOmo1/ykgi9M6ym58q7Fn9S08B62Ng6wvnRBg2tEqKtOTLgQN
i+RzCm9xrc5KC73GKcDW4YsamBf6p28Ap9qD+ZgYmyK5MuIgxgfBhi//6aIg5UyW
QylcH543l9t+0yIcs37lvOq+l8QjBz4potodRXSCM8SgsXl4IsDVvKHCWLJ18SW6
K+7MpVAj3lOd1kAkQu8RJf9G32oytUVgdLSTT3CBCh3TiXKUi6OxtyxSghd2VAfi
nisvyclXudYmVbTjIwgVwJ8PXSR2whuoI7uYi0LrjprTi2xuZQd1/XTwcIIQ6/Ro
H8evlzF72//L1VutIj+4+dTZoaa965EJEt+lTz8sc4/R/AoaiAEeJEZbotqOwYLs
R7owp3T4VS4dIYCuswkHjFk3VqIVOOHxV+rquiFYfQwLFzEpprupPABGB6OgWXLV
/+9nUe4x/9p6HzSEQ0GvnH1PLvtATK0iNATcFhtXswTeu4smLSvnPajMkM5vMAE+
MmfNJMquol9KJJ4RmiyAVLgeQxTathiszCnu/DbHGkFtQaesvI8nKbP7kMoFnnXO
xsH9rgpjiq++0g4f4k3BKMkMY/sCuKSS9oU0lJa4wnGHiaF7ZnLOpSux3GroS6pP
VNxHbnsLmr33yn+beDXscPsWM0jImnspTQp5hejAz9FIOLY1TrrVtD1CuWy7jes/
p1A5PRFARfzzn28b+wAz1Ojy09zY0Mi8XJD1aI2PMGmYlMVdnRoyAEMrcC+kgCuW
NJHqKeRMk+VGJPNum4yKxLm6w/b4K7ryED5g7NDDThaU20HPzOqKIw1cTwPXgXNG
4SbnlJUB5f3TtZ2jI0NZv8Y1zsReuva1E1JnB/jxLVy2+7lx9y0TGFGE3QptEuE4
MBdsViRnD0mYfg7lfrJDQM3dNJ9tI5XMR76lVOMusNltQv4rus7/l6ct2HEX0zGD
WDUAjHHSSM0CyA+pwdQGqTOk2lfTSQO8m8HTnbNNQQus8NBCPwx8yWNb21l/wIoI
sGEzUI+U7L6ws7LiHXofKXR9RLETOYFosA5iuVj8r2R4r4x7JU1RMt7zasIK8tCP
kMBe8N1BDbyBtSM3umKFQlw7xLw0NvX+QrVCuDW9pr1n1ZW0gRfIu/hNUD9ZthTe
Rh70HeRR7W1/tsumaN9ZPR8imBBI5E3noqDQ7+95IuUhs4+GWYwIIiCNDy4YGW7S
Ojm9gyoZJcxxcxf66SDSnH5aeGLSR5kdiHVaV4I14HjcAKNR33n128Jf6RXnJs2J
aFujudWNoGG+hE3SfoEWJeiK0+1hcSD/CTwnCG+QGZlwXrj7AYv0oGwn4US/+U39
rmpdDRrGlPzpgwftl+FqrKb0NO2LTYqL+3WXqwEtLILbv6Uhxp78QES7xtOw8Fcc
SXHaIqSMdS4IdBzqp0TkF+BxTD2qJTLwwFvByKkg1SyNNxtyufSE8XgK/DKhhBCU
bCV8jVddmuoVjvh1bbBXz1IcFJEH8MDjQuFP1+g+GfFBcBJ3ZPGRpYxoprLeb36y
xm0DZYduuIQsQZrrbPCqN1e63x33JpCIjGngWnmb5zwsrpZL1nQZzMj/NdtO6loC
v80o+45SXP3KyJ2WRHhFjSBWXgwnWVyJA8ltZutvYt0UTAPaarv6MS6wWCcI2pmH
kFhfOZeiqXsC/fScEbXzpnls6X52XXCCbbhns+h5jaGRDIC5jL2TVeCyJYTU7lXj
+S++SPgTGcJTBEUyNNHve6VT+IEBM1QDtPqZkKuwkyYhf1QPndbdHbZ/k5+HalNi
ie7/X78KEefr9CguxToaPEbwmxSsLsPAYTTO82YnZUnp//St5qNtVjILYHajnV82
Ira0X4apCreI9oWDyxG7lKvazixaCi4kxUkaEJK4OCHbS0c/FFCrXZSfGpf7n6IV
nqMeKDJ1YyCurwjGEGKkpJO4f3FPamhkJMQUtcdHulNpEry2PYpw4WcnxVIaiwlI
xRmFtLEwZ/vu1P99v6lxuQ2JPkTqvsQrRNWeeicRtDbBfBEfUwoJSedZsKuZCI/h
hbDs+ZwWIJPNqEI/mghGx0kt2cmnz/cBFJTPsorCPB16gDJv2sw5dW8Cw2RCzg8Q
7mPs42RRh7+j1jqvZ7iAYjzuztKW2BloRyJkLS95c4Uo8epB1d17ynm+g8fbiaKW
L5iBtNpJr6vB8GgyegFO7XU14FYn/u4OuIHlbAb6tXJLthG2ZSjBhvCMUJfpvHsK
PQVDZRK1ovpTLSLJkJ7hZrvd5SM64vQhH4uAGslmbNQhaH2lUz9ryw18azqeddkR
JBw209HejWaCJ+qI4DmpVrQcf0l9S3yNiU3ERs0Nyv+daiF46PSle2EZNB5RpgRZ
R3SVlAWb514b4qOJJMj1ZCiCz0S7WjtT31LDFYAH7JXotrmJau3lShUqxaBBWjGz
lYeqrjORhImlJbtkxW97mCP+XoTQqttN63/MWPzk9oJ9yESv8Ch0kNgYnbnYgICf
C7SuAVVw+N19IgPAXM0Vvg9nE1zUJAD7jpd5ay3SCtS5VI5Wrt4ml3lXqULUk6k6
7TM1qpqN4Cd8zOxE58HJD14HNl4yYM3rlRXGUnkkh+aDk+cV2k3I8VMCmKAHS3xw
fWJiyBQGd0sn/6SXyd0SowJWt1yxGYBsJcJuVHNraS4fTNCv+6iQGlUiAFrOgc/i
ko2tNdLixrCypsYZy2WjWVUZw/L14LpDEgNqYdUU91ZJKUlmGPkmuy5r8LlpHL0K
aPoGUQKYDptasSybHp7UAKHk0JO1YRfLuxjyMEJ3d2QR8OotzWqSSZB82wTXBtIr
hyIprxkBHbK3tY+pcqANYZJfCPJzbPC7Hk7A44CIf2wxphmAFWHbl5qAUi5Sh5N6
Zy716WmWPOj9c6mZQF6GOR1GsC5z79Pxr73oToGg2nvGXc4iUNvUx0drorcCczXp
iH3L48GYFAuR/k3Iqo8eKgKp17Kh6z2lVrqop8fXgd4E5vMQ/bQpsVJE2RqXUqLf
12X9B2LsPH5/dvRpU1y3CTJTeS4MRSF6Vgv+IGF+oJ44Y2AKI9BDR7mZvupefzLj
qWYvZsh1On95lq5KOOWkYt0wNwD2WmOF+WsGPR4CYExZfpxcPL36IwmBrXbQ5oC/
e7eq7z04cE6yjTJloMNWYP2gwBqlGI+6udSlcv/N6cdc7gDqav0U9n/Tr27udbh5
IkWDHa0j7nqr+4YshOmZjWMwCpZgCN7+97wFB1rmoMA1qnX5VOzDjgM5b+1vCAKA
X4ADZZW7riXRrXEwFShdUg5DPkQWJe3CY2Oh4JRvDpYEjJDfUzeLMSrd1l4BCa4B
lzAuQwfG7bzPSjEjgBYToXxt4JNz9aRzMtNLYy/lhatWqAeOltZg/zX0G3F6Pzxh
CBNxA3irWqdZe49Epu7jyN9cY3SWAlMUAjSLfDnQofJf56Y3Icu6PX27T3aLdLzp
0oJ1pBx5o8hth+UEKBPrnMwewxoPcI85DrCnOsi8R9NVT7k0ME6lQn8SkLNAiFyb
6ZF1IJUFZuPryzP2Lgzz+RRyOjQ7XUaqa1CeEbP8QaQSESHlnvSYsnZqy430jZdd
1uZscAteLA9P2wrPM1+uve30Xx2WqRMkPoYBvxyYDCV70ndbleNYl15eDKk3y/A2
RpI3A/OiQEij1E4FqehZZChIvWI1snahoNkAUDnSFz1aKULKTx6/ywoGwDiYweUv
9/qd//JJ25sx/lCcpFkm4aKPzyMhlR2trO7QxXw5utCmh07zOgmphf4+1JaCx9gy
HlG0waowAx3b/3ha7K5h0/JAlhpJPvB9dbbc/cb7fP0cdSH/FANiIyyh1XOw2Byx
hOpD7ZY1zg2ywbhOcqUVUlLjGJT5R0IuhCifyoAoUKqoyyLvj7koiF2O9UjAEocI
J5NOIqVCRlZ/7PcrFELxMu385tDWZEZKwNHn09xfjJcTLcAxoOp9SGyTOuUzTb4h
w3lJSNgbB8O6vDoGq61sthBYDHru5EdlI+q4IAoOCyYjEfwjoT8+65iNGoBuJPy7
WYMIJ3Ojd+LY8mfDnJmOtNwOm+itrV8FpDug765z32vl0GwJHdS3tQ5D1KWUgQcr
hQdjV5AyxLquztrh0ceRHwJNzlxgtPME+j+eUcxO1C8yTSv1d8hAe93csmWAEy7S
t7g7kYdfW7AIVw8JbvPDwMhY9o9cV18zL/zZhlGv2DHxR9vx6Q3mg3wufUTgv0fx
o8SBu34e7kL6bKuTA7z5PK7nL2bn/Ziz9ct99EXGX7awyVSntIgrxDS7pOK/aCDJ
cPpOcN3qNUzg32B2WoDwoir5Nc/adVpLfZcaRoLOLQrW5XguqnheH5AxNphLT24Q
gw91RlIex2MdYrRbCDs0lBT4LNjN9Pt4hYolGzR/7n4qWNu8YkW/9nhhtnX60dzg
RscrfTOboSVx2QdfcRBrtVaNVARymhgoYy2jdjR2WC7Nn1sdHJXaUypR7W6985rG
wwThQkwK6fHuH0JuD+cNVazPhyIxEYyzfwYZMvHAuls8DMN05kzmlI+J7xEcfgFy
K/UnWDjATDnl0bV/WokUB8NRS75IGt41YpFh3TeAmfpGJHqCplSdgYIXYbgeSAA8
lkkcHpEs8PqzlKuLSq37toXJ46q+A57UZ9DT0tZn1HyIjES2g2CEuWUukxMkkDMv
+NUsBYz/fhMy8jwXRom/W89w0MWN8VReDk4JK6ucxBOEZNA2WVSV4/bKSSJ0YpIu
KpV7WD0qN90OYTLT1uGQQ5Cbcgm03lcUHc9fvvpONfDALmkNTFA7swmzOaQWEXVk
Em0JbylVagv7LFiq6m7KHNKA5cQtGtT1DMEqg5QgGbLOGFfuermedRCgtMANYJLq
n8kzfl2Y6VRR5o7KqwXDQ7aWeoCqSlfap38adyFIqyfGGnBKh89JTP7TcptsmnDk
uoSQPu8NJeusp1BjWjd1SyhyQksvqGmbp1p4AIrmSOfarUQxanlxcgzX0XkjwiLW
sFuO1a2uWj316Mi9uSw7QtPnAzI8oHlJ1CMeDAMPD33a2IqfuUXI5DWV7vv4NYR9
RjqmzIdd2olj5I8yfYaHoPjTpsK/qQn3Xvc2tg8th3f52d2M070wxQmoSDoeXGU5
HIgqmU2YJbpUuM6yEvPP+nvMaTxN6Oo47vYI0VfMbEIN2XVeaxQgZF3jwerHC9pI
pTBElNC8ngtP35fRZapH3iMxtFkSuitpeUTDskrI2a2jxSCVfJtp+8r9L0MTBOgz
b+lKZ6ghnzTLmn8RP/wmzom7bDxwT4RA5Cg4QQ/a+qRgjkUxdTMipWMRxowRuqRa
UzngXcjZEwdl6fGVLfh8Vqi6uz25v4p8J9bEeEVkkDRJFK/nJX9BRgOwynoXnGGU
b0oJGzQZ3YBJ8XGhXrByOFst2FpXewW20+oltg37+vuyCkFrR22J3fV8iGcDsEka
Jw4WbVa4jzhI9DAsnvRxivvGfjrCwvOK5ZSpT2tP5zXtNfYHcyGxS2lCDMXb6y9A
1JG55CnxZo0ABD7SqLkj6wPSr1vh3IhqW60MfWRjIK1DEofjoWMDelM6adB3HRI9
Ra0XsjvXvNSZs6qjhqeMMe5/zw806F9oplsZNC4XOrkuM9Kp6Y/76XsrQdwO66z5
1DFF1FL1Bm6n+CxxlMXbd7sKyk9ubT6XLOGro4sRQyx1i5YsC1eHTL/wwlE766hP
stvIOqpVcXv8XkRHBoeM0ykj+jgXMcIP+1/vGUDHxGCyF3EdfrkDyKPCUWfbM/hs
uXMAajLDMhmROH5KJIjTNUv+Rz8uJ//rvEiRZ0WFknZk1K/0UjVWaG/b6N5Qapd4
Zvc5NrJyN/Vv34M9YFktBJ+zsRGzfgkZLcxRt4rJqzAJ0rDqN7avT9alvwvNyyKp
sIGmsGo3JbCO7zekuYYqRNZi0EKnw6luT5PWu1fRoQKlQ6/xXnoqC+dtTFHlYKvs
gJgAgsgtc7F1wPLVoGO4pYbOhkzZDeudAfYp+T9LK0Nk1lNFk/9RCHpR7juiECPS
Y35QjzYwdGVAb6w99L+9pZLwK1L6rrQFsS9Wd+7U6XfGCmnsyiEwKjdmEazpva8O
u14WCMYr8yUfV7f6fy/pNlV6FHWPxIL6Jb6jfhcxoLkXiA5Wcn+0joOjmZ9jT57U
UHve6htZ+DZjh8Y9eKr6T2y4p1eDKcrvOrpLQ0u1aOK14vrGQ8AxLrsycaA/6Og/
tTereYDOrhuyd4ed6hQEKZQyPxnzB8JIjnL46KqRbOIE7Cbm6MO+eTjp+5ZAMkJS
HTwXxyKjiH3lkuxuUeVvP+zjRDy6mqZveqdrWrtCRq9vOLIsRzLofrIy/b40G5yG
r60dh3sPHyaw1fNprZrKeIx4puoxWSXoMrCQj2JbY8aVQdS/k/UumTBkLdXgrtHf
USVkwPqQK9r3obS/hlCb6VahSbNJDiN3wW8DGxGdAbCHv7eJS5KpXn6k6tA6yLv3
XBqh1jtBRMAcXPjlY5YKPIs/X5X1949r2wiZRmicdV5mZaNbH7GUNT3daPMFLqr/
KdoWN02z5Z29W1+d0qxkjFmMD2786bW9GZ6Wj8CIEiYDxQSgCvY/vJaeemXwiYh9
NVy2DNNY1jGdWHMQPfMeo3SZrTZCv/0UirwpgRO3s269JF5ay7OVnfpXWwn1LScf
avE2vdQRABKDhrOGUTwflDuqyUDfs6EZ/mP/K4d/O66T/9CjWPWhImG+Pyb5Ylop
3NjC0Ra3rcnkGP64ndBNMSFnxAxmYpm3IaHLzWk6gukXniRtgac9dcYmzSZ0f+dW
NYggsCJrN982Nhdrf51TtZmf7assNNxl4BUV7QCSiPNAUGxw5QVum+lcIz4xIEUY
rd7MqzHa7bMcHyDdmgZnRnWAtgxUq739FiMwpEBB1Vt5l+VsOBNfEUVml6TfHubG
N1FxvgtaSNTvWpA55BcRxzfdmVOM7LKifr6fot9JRIRTm0cXl1jC2mRzsp0Q5uJa
iB/tj0NI3xDcjhm4UEu1siEhFd7o78mCMnHeyvD/mfn/eMv5YHp4ziLdt/FVWKvA
vigFaCAvE5wvwJT04pjYFQzmgcDI1aFqQHJ8QAzDr1882z/YWxwFxqsBpumAGt8s
4o4j5ElNAezb9iSlOV1QUi0Uuzq9W+SzN4Z9WtARp1yCYimhLgWOed5a2Gx92ecJ
ux/lTxOTo1ut8elUB6kXwtq+ov3LRedNmBUhy1gHDUR1f5iwigSgROt5jOelYRx/
yj/pjU0Gmy6h84xrAW3XpfQSm6ihq39OTswuilpy8LkuYclwgy936MBDYco05YLc
TKtuptU7cdWllyUfs4SzUF7f92MssNVofz4zFsdpS0B635Ef3NudNMTlsk2i/vrJ
KViIrO45SmbStNJuzWhoQEOrYLAoSZlVaRfQpAh5kBd9CNkb7BWxafG2sbUR2un9
+rml9tS+mzilMHMN5hx2dYCgaDvELwwUNMNJqC5znijWOsSDILPhAIbnZzD7fR4l
xk+y5Cn/jFeSmmHzD+dOLHphr4GDx5xnloC5dst1sBz8HhGffy45oxm72le/AMPP
BhqW/9E05l9/3bsZWTxJG6r7mfKF97uyjc58no3oHiVKUSzPpP5EH3b7bnfVdhCL
yjgF9gsOhX2amkRyiDR/pBkm117FL0Spi+A967eIpeNEc55JlHzKOYemm+jfBrtu
uaN8rHjEA+ihQMIWJMS5SzrQPodVFwIzicZiamh/AEdyJ4zuhZ78zPc6DvaFabZD
rfGA1feJTu8cyS/Ol57MbDl3NU+agc/0Gb5gs/xacMnHcMlBQVYwHu8NhQTBCzCU
3lJU4adikj+LkoZn1BxKkt7TFRmVqt4hhU9FzZirUjDdxiOaibpcyIVuQ1QPTGGF
juetFaCAzTzd2qk2Xdh8Gr3ICvbc4jtKBiUFE/GSUCjQwTCFOV+NbctwPpvmTzaI
fBijiRxJ0OF+I46PK/0Iz8MVrqM0qtccKUJYY9c9ITplz2mKLUB5njjmkhjmCb4V
LbSAWs7zYEpawotwLlPO3e+wZhWbED3r5s6ee8nWrQbtt/FX3xiMOdcztt91SWb6
kqXnE21c7JNXNyz1jjlGdFeliMknf8r0IXqZwiVlWNcGIXlIJ5q/ZnKi14Jl1iLi
HkmsBhE3UHOlrzQz9i3QjLF/AXPgy8QgSnqXkaLKZfJyykA3E6GFEEOOMXj+tISi
I2HsOmYIqeoBER85i3Dssxm4/m1iXN2QzCKf8Xgs7ocytOc04UIquc6Yh1tbu6fV
I5khK2Hy7q5Yo394Hh4peFsybxox+8YgbfowSlqDKuD8hWXvkHOiU2aEvmsmyHvf
NSXKjIjXjalL5LELmuu8lUEv6Z++5tzIQRi8YPa6NOPsvqgvOm4FKZJoLpbLG+vg
EOilv06BPnV8liFwYb/Sqh/oYwPCkXpSCD+Hm62UKkY85zHeBuCUiMSwyf4F1tlK
yOKj4B4gHFuJ7a95bsHB3aRWjzCPArzTmEkvfBHOU2BU43f9q6/4OsFoC6l7PhzW
Rp/XLOhwpJG29GwuMZam374YM4lr2BggPufApgmOxpTfVyzBQ9HPsG9pctNEE/RM
k7YL+WND+oqVqUHWdAxTzkqwj8yJ3TYLNWUscta3wPVQP6rnX80Jt4PfSpEy0Bs5
Fimxd3lhZtiTizbHPOAFDgpdvCxSfD7UzsCy5MgPcOFniEDtQY80h5RZO5k/Wyap
CfA/eUNpy9D7TH7v5nRJNntcob23GV7ae7ITyTCbI/SLqB/BIBSU8BDwO1Ib2H7t
JCuCsv20J0PQ5ZyoJk3rkfGGlgqDRGF+BStaJNJXDE6tePKO6ED9jBvWAVRZ0i/K
4YvcoquPdbF/rqitmt6g8LSNlQW0oURnIWS4893UEYz8lxkb90wAfVY21tgebEFY
UgXw5xdqXaVLEj1kXlD2z9wfbokIhe7He+3/5LcoebOg8P64ScnYz9N4yL0SEQGD
MqWnvLpZYpkAqOXBznxWpmfje5yvajR6XM5xfdVr5E+3QNiVvpdlfgsGjO9F5NEj
A9ipStS8gvKZ5UZ0D3JXozJCy14oa0VTM3s19p02DF7bdL2mazLKV9e46jhC3Ee2
19/23ZB66SGRGJ0DG/y6DY67DRX8NRDM0immOEBmP6jkxebbAINF7M3/WTnZrDaz
XJOmfXKc8o2GiH24NQuKlsDDHrj4qJ+Z3BYFM4Cp/ml9j5sefzZBUiy+qu42y479
UzFJ/l55MF04bolvdB0xfvSk0Cp6+2CZ+2Q42IvdLbHmCalf2T1a2QmGu6qkk6bV
4y/G9WCj5XsnLeVTvB/+Sgv3AQIVW7iTq0Mjqov5615NBd1W1VkMGyPVya8adyYr
SBuBUNDPDhuYk47hEA4I/u8KZeohgoCQfiOXireUgQ22/VCbfqhKrMfzkp84bVVT
cOmqPM5ejoDdc0YpIaeu055fy05m+EX3nPybMoWCz3UMAmAonOXcUTHGmmXsd6zs
gIFFFI8X7O6HPfx9OKATLk9VOleTklLxstpskPHtPCIFz6/m9LKgkh9Edp8MVOCG
RKTvH0gP1e4yXr48r7jGUGDTytkq8sUNjcX9OdUvc/mxFY7adxkTo+rYlQAMVN8E
Rkts7uZaJm3cj1TJdHxL00j4Xd+QcGyEm0GirNh8gYzWw8BKSidEtOQ6AUBo0a/D
ZWiIGpqj7Z+oj0eBRXVsvSTDc1M2Vl2y2n/aCmxKoNiv3CVulBXR+7wYb1ArNzrA
yVdPMGiAFTeU49AWlkY7AX1MfLJVzrdJJWaMzNZcYi4YGQkE8GsZb0TtLoM2TnSZ
uZ9GQrWbh9l7Qf+Uu9m8WBxvCeaWjeB2K0WgL9MchjVSeXhKHMfrdETN/7/javnD
raKkzPB3S5q7Nlkupx7kqHcC3WObg6I5/JgRmN41uJ6pCzM1aUYHA+nMbViMsOZd
pWpoY+puEcQLbR7CqnFbB2iLUCNgDAZIpfPEwtpNwrJn5b+lTllqXmG6y9Q7fx1U
nTiyoDLC9zItNYD9u9TIYEEsfTsDJ/uF+TZD71Qzd4PKasM6fPzduckSyWDA3WLQ
JrWXosgDAFFPWXwIkzZoRkW037NTOCewxmPvao/rDtTj0xSDys8rMbqQW3RMOzgY
wCQZQEVu3RND0089n7QWa+p68L3dWtZNJn/tVdDU0ZnpGaWF+We1SkF29u1oFYva
uqNORiRbS64cdswIXiALOYLaYQy4RqjS0jc+wUbn4eHpeVSfYKhLnQfa6QSO86MB
6QUctOQROC4Gv+V5YvkyoQDbyG28acf/JpYyE32MsyqMc+kO/8nnhlkjQf2QEKZp
WZMIP7lXcFxqslwfHCTZI2TXhFaPXbv90w3OIktZe7mclC9Qh/uP/jF6SgyhFdmB
Pmb3AE/uo4bpVpUnq5Xf+jm5WI2bSyC3FYV1UtEPnzOlrln2Ib3fo10QFQFg7aqi
M+kZi4bQtm5wIAQcwxiBKlBzxzuwp7B5Km5F8O6BE8nzBB54cJJZYzaDOru7K0id
+TWqxkXpxUtiR2s7loHuXVJJZfDqT6P/mQUTzvodqafJxOo4IfLSY1rm9jC0Iz91
PMgogmyKHs4lPXKKLcffSvBnzTQkezFPlIwQVyJKv+KANvgn/Jifls9r69EDjvBo
ihu1nHykO4lKYkjt1XYMCFu10YF+6K8SOEcsuHS/kzbOihSg01gHVyUg5dNv1M3Z
jkhIJ8b01nz8X0MFs809BE9mIGzz6koRO83eKgaCVqcdJrAzcKT5pIRsAbEODKov
LbSyQSlvD/pM9oMyJHVv7Pqdwv8yyodo8HiApPE+K8irIwVAWiL8Rgc8amytqPgX
Ja4NSkDI7oUNQ7Buo2kfJi8d/qk9FSECRHUFkDu7PQc2vphRfDvk7/cQ6Jvqa+op
zZhZSKDP39eROIuodQh2DgaaR90rjQf8HLKRExpM/X3YpgeW7REcxRsD16pojhcL
dz/qufc8FYRlPxvLkH7nberh8ctyCuQIzqWG9LD+JWKA1DdY991Xe16p/lszcviu
iNkLmREcpRR0XPtbMEzUhxlLKMje6DhrIaG1CjDKSyMrENa2Ee/lzPaPU+7Shr52
gVWcmqXTu6y287OfCdPJBW5gwx9y6vMT5K0n5vgFB1KdVtCVUUOwFhbduUZZCkx/
HgoIm+HQHeEertopCgtoGV3cGf71xcDCQaVsrb7cs2ENR/S9cxE6d0N7oGIc5ggm
vXrcIw8oqpFgEfzzI0XZv3NEEiRP0n8x0rGexbHYydVSBm7KsgWbuRw5JIb5zsdi
v3jWuBetweW5+K+nMQR3STUwIXj5L5R2xMcN2R/e5Nidn3UGXWk+sLeXt6ncOe04
JzeAeCPyDExMaibTNZQ++IrhWeUJL+qd6Yc2u/aQhlGyw6FW26t8YRrIhgLSU83M
+m+VPs5pXoxG8IKruvzgOWvNueMvtQuFlfCJYDCQSpXnZaDNNCbPrBtY4b64AEu1
YHnBmNFadVc+JAmreDKxyWehWv+nPZRCTo56w6HP7/CBVEJDsDSaAfEpXvV94J75
fotdKElGscFFeHFnKYe99LT9YwkMUY6zSTdCPHJhEC9NoCVR+zyOf2W+tq9uPd+O
XpdPZQgxO2WozCWD/i4jllf4Q29cKkfdq9KpFbVSFxZCvM45Wtx/+JR96ij2iQVN
LfnbH4me2Kp8o76iM7C3yCv9kEe6w/DG2NzndTW+apmf24NqwCFfhFIZnpvoEMvW
GRvCl0D+EUdvgw29P9HFuMS2Cw75ppxDAK+z7AHytmrKxYtecDk7LldXZMURtDR7
vnPkyFEoMiAkGNUckBwTbusuJpdmKMkvlnJ4u8HyglKGAZ8q6G0TjIuUS5Ij22XD
PO6+8kC2sBjvuZXTZGRO1f1C7qWI8Hp/8lpjPXPd4nwr9me8xMBPm9XPvGEpwHBu
aZse7rzm5Hq6d63jjuIh5cVEGtLwGOwwH+7/Lq8oPmk2nzkmprVt4Z2FO4TwZt+J
QRm+c/ITZmTmMtnSFumoQdBnijXMJUhtrWN+tR1/KglsJ6hqJj6p2krolAxGFRqh
3poZwKBnu7hhH8Yzh/NLK0ru9p3SeShfMrSCGMZ/xgBKK+avq9IiRtSaQ0JZJn/4
bIJSLkAYYJtLbwzwCnzwD5UGbf7abckiCcGubWY25APZKIGQJC+w2yaGBYxLGnXV
z5516fLap4y1V8W+lDTVUvy+59rC6s+Fyv/92hH/Mdh+wXYvHOb4JbcI7Anr21qC
WLD2RvWmADrWbsiPLP72ZjnQ2oUF4mUhwgukDS1GOmQhUQjl021BQfjFxjglPU6w
pQCSZdj7PjO5H/jMXOE7/AdI0kNa2ONZ+EEtfJ1+ghbCD6q59WQxX0UG3D0t9ExR
3Fs3TY6mINS4dO1zF/l3w1GmjBGYEYTeFokmKhEZMjySPpbgSIHEpYprwuJwUpMB
1qljrGI4K5AOha3NUje36vorAmAQGhztbz6Q6r5oZeWVyJmYEEkEChWoOzIRcLCh
Vy0J8sPxkyRV9/kjPjPTpMvdJwDZDxCjrI4KPYNtGvgWfEAA0sm+7IcdezbjE3Fs
OZ2D9tX0BkTSkWttHno4RJE0uYk7rbeJ1xGeBS28AAYejb7SCGe3CWman1ypQx3E
UnrmrHL0Bppy/X2GjK3UWR3rC+v2y45FipeJdbkLBoGaM0zbxDB8SmxkrvqFqEEb
EOP6Az1jM2e7EIODdoEyWy85F1Ykuf8bXGzUukDsIDKlNkzJQIjw4VjalY1wCo4S
cQqW5TeB1cJSeL2y/qA19V9LVgbw0ZSaXnuWnVhET2yMHzgUh0rHovY0wuazW8JP
hC9GH6CI59hbokNK9BucEV21Zm02lX/vM16YfeiUvjTRhwuEqLxckBvCuRlU2iRU
9cDTkOY2+4Ez+AwQUNdXs4B7GfVgEsMwQTWQSPlhj1BveEGoyobbHE1AbeOgPsYq
F1eEqi11Le4KzSIT1d8mGlp63VITMOM4R/rhRQ8/UnUed/CvMXvo1FpAtzMQLpzd
22X183dipOSZlrVaUxkQXqmJGCCF/zxcFFe9Pbhkzsq2wCuT0rA7nuMI9Opjn9Xt
xdXHZiESagMV/REGl85bIdrbLc0G4nh5+iUYyXqs+XNCX4z0QPgm2vwUZAOxRObt
orj6OFiSS+V9yPYK1zC0fND61S3SF9bz6fFm/R1o8p8QkEsgFYHwj9DKk8+NYobr
rcihpcPazuR7EO+KqBP7VaLhq/t+aEDREvWqAD5ozN/+9d/Csz0LNUZn5qYlqLLX
u7wtWM7UO2MSXzaqBlXRUEO+kklPQwDVxZYyqsHzYc++wkNXlYy80xsD9oAvAcr0
x7zM0vkgKvsa304UPQn4XNwlbZeDdSiweRVA/W5MzYFAQpNDF+P08EkVj0CUSLmE
vhL7/PCtgjqCPkM7o/vM9U4HWMFTyhLxW00AHh6eWp6jGRMH+d6lJxjF7OvdRwmM
wE+fOhBnmcrzo7DGLjPKkwZE+EiWd/bSrM+krVlnuFzsx1bw55gi0AaVo8DuXstc
ir2n9Umqpkf9DUqAX15BhNzInknqNPG6vf+zPlbRxug1zjDEChG0O6gflaBJvEUI
tKrmvaI1SMC2SDIIsMJt7bYUhRfoOj9ipqTpvTUVgn2cCD0JghjYQtQHL1VE/qV6
pFacr1S9HMztD022Nh6YjjF0enp04UY3pk8uaKkaZiw+M2tG3IN37PxxaFRrdmuR
utztV/IYVsJj7b4zwkwgMjyAmeDg4LcUng8BxdLC5GdBD2ly9UZeVU7ss57nhQju
hFP2YNrXoucFdyRXxnri4yzgswRi1ZAtS1soTxsFa10E8FHCJs+u72gl1Qz6sjWz
jL9AaxXeqXx6kHZupjFKcoEg7Cna9bPBqbjXPPXXYDqeJn9yC1UQm6gHjVPqsrzt
py5Mta2etV7BeDBS78aQzJ8SLXsaUp8Bb9Igc/sF646Nel3WvhZCoa5+oopv1Kxk
n44ldd8xDbsRue4k7CQF/icZJmVLVuryaaoApaQi66QlE5pzAPotxekU9qKmCMY6
1lqZw4KPKlKO4i7kochMUpqlz71iqy59ScaJWlZzNKD/3kUg/I1sU4yzn/b7Z/XY
uGVbfuHZTz5pyfViSAjI+tjafr2Aief8zmy3R5kC3oF5FJ+rq5E+NxluTSRrXaL3
3ziVQT+qULO8CQls0Y+acHq602xRxSpiEHMmG94M6yaMpdmendMRSDccGhb+T/vp
3SiIMHaGV98QIcvyVC7PcPwKwmQ4L6duZ0XAdrHdhm6xtoqURkp7kJSpYc6g4GYz
ji6+tgMqszYpmPb7Ie62Ebkrys2Jit844sIXUodUeTuoXv4WXMghTvwn6ZHEgNh2
osA6Reas2VmVvb0QJLQxNDTvvCbl9iq8gaineU1Fp0r2UxmjypoozEsY6ZTREPIw
q/CApaGrzssQ4yZHRzw4+agsdgl/eRrZX65ycJhgIi7rkMG0S9HcqcLhUm5iELeW
aLN5C1ZK4mR0+b4ebWOTXj0/9iDtKO+v6WfYTWfslPpm5doQwTht2Y3mmzFxwsdF
y12XhkZmmIrdcSZtRFaX7GdjhsMdFMFOlwXZD+lHjaVLxqN6ZW9NNYWnwaOYlOpw
EdpSxs/smznVuHoOtsY7EqIxYeB8RAotWUTkEp37FUjmt25lNeHb4zdg/IpwUni/
cEF1/lAPCj5vTz7i1+GkOQdhz+wliJkCjSe+rPnk7Q/AK+tbFsD1GYyU5hv0Mr71
NCLaoBZ5KUmmWwqnt9kICpHBQs2sUoGAQFTgnz9QsARpbDt9msfH5FBMyuAG1oc/
qmZgI9SAeGcfF6HHjbjH4NpENyQzKdnPhpPn+wcmvCzfJ5GJJWnBO8XU04cDj0Lo
hlOLzTcODYdTeRQgajHnULiPRBGoPSKWFNP7PmxjtPNtJHMLJod/mpFoVnRwiyzo
isI7vH5HFsPbxyQ8Vo2LQFVp8kk7S2hvHhoG+juMuxWb/BARaYfw83eMeId6qXZ3
Iebh0GTb4Rzw3J2j1Kczsp8nV3vJz1S/Nr/h7uKLhveoeyKCoib4T08bm21t/uTx
z8BUzyoIpREdM8ps1F20tuLW/q9LXh4o8SoIaaLY0kwuNxMVFIDwHitDoGzoZEnB
UpZ6kuwKNglTuDlpHLs9MX92fpUQSf+hCNyWC+TIAlDa5BuFebSxwH70mHlIqpLT
h1uNzo11xnx1tIV5G1rtb+bwLWjCw2wsdBH/IIRah197YjVqDnbPazt6J1njaj0k
FVRKlq/pQ5vsnKb0UGmxvSb99PbWsWw1JZHl7/ffgpu2ADGy5CXcnSa5CcZIDY43
R3xdpwKbHzHdodW10UjuZ33ITb0CeKBUSnGMMnWuIK99KGMjf4XzoQ751HGGcwPK
pOYJE2HbRuPkQTXiQprQskDp0A4mJQtG4MApVyNKo9UMfZ1MjqWJoopCTs+6tNpm
sE8QvcgqO4mT0mxHhzh6yr1/UxG+/sDXeZS8+1i5q41/T3xSxq4/op0xP5S80E0G
kF3q+Je6TInb/5pXNXVDfUhG29x9mBndpKvbDZoEYVnvmyzMwrYdONaYrThIiSx/
DPo4oLGaNwbqNhf7r+Qbu8MJeVJGsVu6IHFuMJxBrhPON8kIWWfWRqBhyF0huKEm
RZM6PF75cdl6TpCuLWRTZ+nDP8jI8+4kq7hROy8MgpNO0YguWMICV+hR71RHjPDk
+Q//3/hvbGz3JmIL6Npx4offXnvLcPsHnQze7iKF3xVXF7fMUsmCrO0h0e6sQTCP
PD3eAX82ntQwPwXZKjkL3FyhCmCUpTOQIavSjvMEBmXC6oAd771W/CKB81LhvixC
kSDApMQ+oZSI/orIsKoQ50+Gt9HbkFkJ+njsBF6AuUk+FlOpzkxP1YCk3w/RdOzA
MLCSltGrl1p6DthkPorZZy6lNQp060/UC1lBaSCB4IoBEGTu+7TT5HwDnhBvek94
j7hXW9pXJd2fzGr2EZYLjoJSmaUnyU2E48yPRvBXMLV0Z5UdRP0MLgVchSbFl8Pe
VuWLqq0sgoyUVjPsO+3DNXbXmlLKmwW1WVQxohYnvHpcn9Gn17CgglN0xQOVQucd
gJiqcvgmEQ79Pa9tCMQYe2eMPHbcGsIFPr1W3Z+WLq9StfpKj2h3BRFpx6Gc4SSg
0FW7xtLLN2LX4JwJHijodfHl1LbY1pxWZaNIk5bVfXZJEKok/l+Eq6lDQPyJeGga
Xx/ieuA4aoOYYP0sWJw3Q9lZcXzBxcuL37JQNylIabr+WYW9WNlERqEkKwtTJmes
TNhF70mmc/OpyWJ06dVj0sHBr+ZvrDU0Ka2zLYiAoE4/FpgtuSE154l2DyhJZgov
oW1JL9i6ex1AA70vLMotxtc6PngQS7d+5zuucehPRZJbhCUIbsAM6uDYnR1Iosne
KwmWy+UmfS/IY6OHkwnDjRoVXiBS8R6vUUnSgFnTGrggYsYbcGFFJms56cdY8rJJ
Z+uZAGWgVowlbMTV9Wfc6sGfEN5/JnBp5GgD36VNF5KlPa8CRnrlBxLat7a3dWZx
tXW+83YM05ACRIqxjWMXP3stHAJwcHVBPEhFUhwDBbauQ9Oyj1WroI1ry2r+2lN7
c3ncOKWJN8NMFTAjngmo1fiwknKWOcanhIS3AwGNeLcQw/nOABppGDyfvWZyGnKX
Hcj+xcCD568r+FpqE3Bgk8muqo+3d1k8wGNfsb43NTxGy8Wzwu/dim59rPJvkUUO
cEhPMk0TBVFbfYrxpbYAC/B1EajsnpWZp/wFsdzrE4ONebS3fqUXnsH8ta00NsF8
Avp623dSgh0MiMpYxdjvVuaMW0/TYJXAlVk55y/qhLwehR/pDA5VoZ7Tx32hYeMF
n71dx5PuhWyJQC90CffdtUYvL8ruN+/Hu5luOJ9jSFm5Jq7Q/TTyizPw+m/kvSMj
VPaW8xt6KbWgyRX9Z8qV2Hd3fwwU8jZhy9pQqvKR6caL5E12EQYL8Sh//ZdiZRdF
Z0ctIwWoKRMSNqAJDMRrr9tpALPJVY+fJuFpAkfiyfQUpCoBmsaesGmhzncUs2jm
fWEeCOSOeglvMJ7Cn2DdGvmyNSknumZwWIx0GlpeJUo1ChWhH0Wf9ZPOiBpqBEGJ
NrqQ5cxH4oPo/DQcGtpBV87NfoD15/9BDOWxz2csvLQ2jNeRMQqOY3fm+WkpHcYT
eOn/sLyJUqRjqaLOlRmZcdWKs6MKk2Vo4a7uSX2XFdA5WzAZoNieHUStHc+j9QzU
Q9zsHC0UN0uwBzVO6hvOaUK5eL0I/2pjqUQpTcnp/Pg8Z6DbPRvWs1VEeSMDzG5t
CxGed3SIfW6/BZ0jQYnN1foRJQ1Vo9Ce3zFCfPwq3YzljHXGljyYeal6rChgdigY
qO6pc+8ysKaORGL6UjxHtHDGeNCk9oZhq7iiA/79SOmJK8F8xi4fgnQfEynAprtt
WFY4+Ph9wXWuEWFpUKLY18uoCyVISZqbvyxLtTyOxX06CLh31lo2iRoP2T3iioiB
/D0isVj+ClIY5+9+KYwlUuovwceJYx319Z06V9ZINubguDr8Gx1yPH3FonaXvt5k
EjK5weooRuw1sVM1Ap2Dp8+nF+iqLPymxTSKdXq+Vp1vNx75QMXNbQ4iyio5LaJx
Wdi6o0kUCJLYiZIXquBMHxcJC+ooxDgcre+g0TVDRtmGORP6SUc/P9lfh1S1tnTv
3//cXTtXA83+h2smlSsLhAgrG89RRU6GyyfsMLH7cBfT7vlDe9oaApAwi1BAn43d
XqliPS7yahIIkan/adyV5CarCi5LsYqNZpaqw/4jyoZZKxv3xitzP6h93DTk7cv3
b3xKKP8Vg5LkH6VeIBmXpMsi/YCR0f7Q1I/TwhVmOJBBJCoBWHJN7z/SbCIft7ea
Lun4a/vDUGSrvIO5qEsjLXvMKQoo8cY21bXeRVkrFHyLfRIbWgsY3Z91AZUM4Jhb
EbaJc51FWAIlBZBOcpD4hCC6JMTOF1addwDljpdjITVzMnbBq/RTzLkFTquCON5o
oy5MW8c34w+PZjdo9eFzxukeibgtKcfzkOl81f8CcWtk3BhSaFxlUrqo1GlzFexH
fB4GE/DjstiO0V/llRoLXUq506h3wuTbFR42hX6chRt/tok81/zlWnWhXGFQmTRl
Whijoyb8keE7YEbbJK2HHrt32h7wOKsNqY9fkWYuXepzkqBz3vUKzAKukBJLfO0y
Fwe9x/ILrATEZmjjYXBeWvnxhglyfRijH27o8f6gDNr2+vxnqyYFYlFqvALQsQbN
eQMRgrD0HF/uPnjv6Kwy+AZf+AqU9DdJK6bSo8sOiyiJhQLsa/JxebgrzVwCEESP
Nr/oPCheKPyjkRhczXlzm9AV550KwvIGxP5VoDZQliPD4mg2OEvTm0C4HQ0lGtxm
H0EM/bR5RNeVX4UKgyipqzNuXrAajIPOp0GQeGLOakV90Los757ksY42oUUg76wi
l34Amqgb8vb+5MCCuFkbpuyQn0cmyb0FyfzxS7ThVePqxYaW6ZdT7jheXA5n32ir
N9F4HD9Q3McVezKo+7Da+5x/VhE9fALYMWzpSlcTulTu6yVquEHla4uvxwPDC9u8
g6tDJD8Xoal/2hLbWw+SSj3/FL44ZEVztbZgWLNCPqrLIyfUxR3/kSlM1g3l6Gna
/8RlTuqewkT5gTGI7j7Cr5Eo4wK1fdnnQ3ZIFK5qdugxfngNv/rgn12QbLnAFpMZ
YnHId5/YB2cHbauWx3x9rttuw+bkDlyx841daSqe4Q+GQmF2B1y1Fp/MgU1OHbd4
tmqpgvaMc9f+aTtceyt+cdVWREocCVrCPjBmEuyvwYKN6XaiRk/cXvzvNuKh57AZ
+3kyx+JMzqq8QLRjw1psATJfFLX9rgp0aZ4ndEYdj4UdXpJw2+3L9p9v5g3ePWI5
U/VTxdvCmGPvHDUCaJsDDtUfugqyYBdUxvBHnLsQlo7lUqcp0MABC8Gic0yc78k2
oYt67JHj1q5xTDqIdtQ0nf5OsS1vr5kjM0bsWuucLyy9PRMSo+8O294bQRY82TnB
ex/5LZ8SMFIj/DKQAJzaHGCQsaWLvfypTc7+9IxWC8IZMudPBj5ltIii0rayBgKg
wB/aYHLfroq+72F89TgyclK5xXi3WJxjkrcVlAj86DVa4FeUS7uUV8/bXmE/UGsj
GQOuNrlc8b6TKcbdzz4e4h28cjKWhlzLah/3Zs6lr7tAni39PVlfJdCXBHc9xCLd
XQv1+PFvHlEsAXIXsOe2wMSVfLcUucr0w64AFmjiB6CwQ973oI+oQIEBrLQOfjJC
dmwwBeOIJnYFezzF6noiYxHXJVjoeV/tHtapMJYEW3MBmPta4Dk+JH9b9PRSYn+e
/M/+9YgtxFTLcmuc/yeYe08a/JXJ9ifUXrFOSFrkI/mezt2ogNBig3PhrL0qOYU2
5r3/zTJWbGMK+jAcl9HkXEuhscG905Pr1VkLWxz8qrOMWnK9QuSMvDlrd+KmeRM5
ZG5sGAazSy6w+9KfZISMeouUnsoF3z1UxUokkXQs188uOeU7TUmSWO/+vaIwLR3M
+lhbunT6aYPSl0aGNE+YRWtafrh/WcgkkE8FuNfarhfwgBu5CMNQAnqgTA7SvnAX
qnFXPcy7r/LV7xFF/lMwzOdkKfzAj02BcWPEMx2xGwaDrOxVmsk6vppzerrb5x2M
bV6YC0iBgNhZlMlc9EYwYxEtO67ZBKxXw7Ylb/mghicCVrKjeJ3/OdS6CJG72/XB
LykKCp8OiRY0tQkDlPTtKFB4Z8iIVqFbIX6xKLiqSTkhAg4BebB+eAzeBtatfE/e
N7aY9+KakZYL2NgQWrHUwI4PCGyif56zr6X1G3GsEkpcHilJW+W9ARrC7DoC/BMn
yF39uqVFwp3sIDYJs3dP872E0fQpc7e2nsaQmE107pfbGj1IPcdJVnFg8KaR48+F
PemEVapZ3tlPOT9fhx39MI3kyr4tRI3xU8n4wlQfrpbqjFS1y+wZjc6QZOAAkO3C
Qm9ul/OaIR6twSRLxI9fCQIoJqjFCudczXeIMJhUm5DCFsbduIdZr9PEa+UcPvKZ
jfDu4BmdZBSzGMB6cMMY8ylwY+SgO4HLodRz03ckeAgCr5PGZVJSJnptKEWB8/Mh
vPlg8y/Xek+V0TmClPDP08hL8o0CtD/xeIwoL4546E3t+OvyVkS1J4+w/Ud118Do
M/Pw6f0fRxfYtPpaCGZSO8647beyVxkTNq1XOtZ8fazNc9e5qUCGiY/viT48VcjA
TjduKjtjJkdrwUiTlZtIZowvdnSfb3lwDFubyQ4IsX+o9fSvV5S6Oo6AHVyB0Mwu
MxAV9isj2AUa3ZY4Wn2rU2J4WAc9AJ3cJQeeSLw89VjKXSIISnguGAI6YkMqNeG7
MQQcTUbnOVxTK2DPFoE5qv8Z3LVg8fO4sW6q3FUV7Dr3czMVNOBwmpjmf8ZIeEsu
uUWpACKQnGU05vyFfeJOrU9wyaTGA6k+bPi/Vnfh5LGkG/7u4mS3WhG38JqJAlVa
M4pYav6/llgXoHv1/f48vdqX4vCZpHQ5RnOZ+0m9dWgKuv906mczGm1elQrk9NdS
PsfGfiWPbSzxiRQG2xfqunpCQf0GRX1g+mY6TPnkKhzYbyxeLCohu9LdGg+4ZZBr
ZKZALXCrlePrE5RL8q5ZqUNeV2XyTJ74J0jTTvpz7NeyhYHa69litjhyE0Th2LMY
bs6vmZbvy6N/7EYADbly17zAGsoRQK/CbvbwcHqLHtJgIMt5+9Z2lYMcLlSUizpQ
85XrkBnzL2sgatQcpRP9y/Cwbi2JdlXDYDG3bPYti1YODfPhp2KlTkB9JaQjCTPN
0TM23BfEjS5PQEdvdraq8tgPH827ssu/yazM/x+u6ZFZm/ujGPb7AM9nmuu8ALn8
fKP95Zt4wZvKJJJNitsESyQvXnlzAmX2ylO17F46XsUUySd+kjqAfpDuazCtUHcw
qqLinXmtQ1n0UCRMx5NDsk5vc7PGhlaQxUjVS93+UEp/VHA/PC168eEmTdc6CIIm
7IO456bCu1W+8JLajWaCw4mtTqvN5Ab8DBDN4FpCPQ9GpkWV6nNwwwHy3L3H1Iwe
U0CXOH8bGRaZCqA7iQyT2STUHvWAz6+jPYc2yFCSRnly2VlvSXmxt1IeQJjMlMSE
B9vdQXDLnJNPwITDi5uztb/bSLYSaML56ng/nHmlPi2Qzq8oSLLRWMM3PyNPn1vW
GyZjThWYBsCWjnKXrkYJDuZDDGyx/dSmOQXmO8Vo0Qfx10qhnCRCXUoKwvDKQXQW
6GtGAL09caljMR1CFjy7jmX+qfFx+U8/q+IuBA20pNqUfWkFZbh5xUvkaOpbvLAk
Wbx7qRGbqmrfUDen0f2HGxlpjDz6cI/CF8oUbm7nRjHEmJY6BK2/bZJvAP9fUtnu
fLFeMiozL01f5RpTib9ltSjB9iYP5nbhnHEV3z3aGDNC4UdKM1DNljJyb7mcWZl3
ZPOhCmzO95kjQ8UiWpbMysXxk/M4FqBP7tdQafARPJePVAwO1jb6vkXoD7UFm06a
10dKCcyn04BX/Wn1D81hngCkeyQWmusxXuhWmfpGzmL8SUFYHxCW9ghbNlFuKkAD
Br+wwznUEFA2buK/WDzMftV4GRwto4cBfeH/GVwtZFk9khWkPQHhXhfwwfM7zmdF
/CQzXJajecHCLUf7a3Gw1t+p3+/uch9Fv5TA7m0y2bHTtEhqw1Ed/z99TusW+Za0
fYG22oshWdTk4W5DwSjb3+uGuR2hYhC+uXpVVWbV6exPpCL45XUBh4v4epry0zD0
VbxkdzgY6uCDFidaBVSOjbJlo9DTLVcZmtCzY6+nVkdTnKwgB3DN6i089TKMuwMy
QGshIuUzkMV/Mi7sclwdpSUQ0Yxd1cVKIILAcB+aDmC3F4GxFuRUWc9vsKG77OIO
+GXjMC3jSMCdc/wu7b9T/d/UdD17tkX1ZOcgosEqs7uGu3jy+nKLUE0lwh9SviFj
R8CYAZyNwWCaOukF1IixBIsyEGnEwWHDcQf2IgpXjfpHkHM1JFnkJmyW1mKCG1Vq
i2rcHgBUlUc1L3owR1Mqp15XLCJIIUMByGPdkGn7yngz030UjZaKHQvH9qsGi6zk
rKPGR1dpEITj8LXJhpaGZM37DqJbq2PZbKQQaSxVP0Eq5PQDTiB0mqHjYocrzR9m
m/yfBKi11yWZPS0mp/WBwdObmDlMgSzeh7T2atclJtXl2g3wF8uZIKJ69MkAyUbM
bC4urC3LLHbdsPRhd95zSPJ/eCdZaoXr9e0IdaTvjUH4gWsX9wNPbzYp3AeeYbBK
YB8lkQgJ5ejPsYZwKOpx8jpD1KC53naCO4rVKt5dww/tgP7wdsfXSezInw/pYaqs
D7orlP0Y+LHepQ4Ickl17T5kGMWvgrDn2klmP2syEnSN1b+X/kfFzkP8cP1KjSTy
FdlBHsxcS8I3rjBof9hXDhbRSLYbvnyx8VESCApWp3c2ou0R6wvaZr/KhUnAmo6t
Uh6p+FtSg9iXkoQ7aj+/Ptkp7RD+urwg4V5WeeN0FmWamqBv9SgX+NLP4TWSklQQ
z0nuO/sb8JssbESo2QhKnYvSdsdlymQFGIZ4xTdR+DRLvq9A/AudYVzEGXafa7C/
7SdrHIGf6joJVKH88A6lSO6dXyzgAJEKBqIXV6FRGzIW5Sd7vEsKBLqj3o31rPuF
oK9VK+4MmUB2ZskpbibIpKx5IDBnmatFIFQrmLipHd8VDpdbHFfCpCrZlqCwDXv6
kQkd7fq6o9R8wQQqnxcFCGFzIfxueEBvUGVFHYuzyTQCvo42NU0UIoDLjZ7MtyxC
RSDaREhtWhqqdsMhq92QC2Sis3+QXwGOOvbJfVCYLtiNMyd0B0Ielhxr+8YbNFck
T2/YN1IJilsdNBcO4zsT1MImRUnCkNuMyOhqZQFr8toZ6SpMDwzrrnheFJ09PmZ7
H9bQia9CBG9gj7xDT1gHiI+g+lOSfwd2IbR4DMlw7VJlL5n12P6QpTs7rVIU781z
TB0BhkN08chQeSbzmAf2VTcq3fUn4V4hWKGmKio/kA5ztm/a/Y9wuw74Ht2EkTyp
zAhtOVODmhJEj5qyCJrhlSj3wfxSAgki+lNK2VaAhQvju7Hi/UrxKzeHl29c77nJ
R6R2urzNQiyQbekAPtH2fZMHmCxlhtBx2xVd5BDpYROqQYN8mTH7kQ0WN8TzqipF
oHTsHcnacRbuqdYWdOVUFi1tnsrJiFNTDhLDUB+EAEEf24fuB7Iz5rVfIHX2Frid
Ck9cwrjVIEcdd4nnjdHXPniq/vZqvWsgJ6GXSTTY8lcqya1SUocZFdh+3zEwrOL7
myN9d6o9oEO2au1WB9lUBe4YRZMUtYpMG1m3N9+nY55K2s1ckJWlH23A0C29cqpp
IdeskjlqiPngiVK9wy1+YJ/3QrIkJtJFkqEXiRGdJBbUQDQM6yzbcog5wIQt9o1D
621zYcXQF1FW+noFf5uARQd8Np1FbWNu5ZBrPs7XjMzZLqN11f57nb0IIH5zmeof
S0ZV3S8fpztR3Yk3/wNGrMdDwppVkumBrejem4yTfpqo1bw9ywSFwsrnHEgUNfoP
9ObEOgtAhwQg3ae7jddFFvcOrT2nckfb+rdQANNcAttr0Bu//rLM7xDLFHB4NnL3
sSKl5mCeqOw346TUE948IF0O03t+b5Lk1KSEZIMXfa26nRdvBOOWEIEskTTzBNUA
TRUR3WmyZlG+EPWb7YOJAJb8qxuq8KEP9CEr4QTeAEs4vh8sG8ARQK4m1WCexs/Z
nZ0t7Y6wh0udrRhteOtdW+Y1aJzHTboEDMRWSd4RDSTx43rAMbp39Ik9YqUHDi35
eB9KPVK2OFigEzxhRvAxgCjegLXbocQcPzMcx8E1d8It7d5PIHJV8T96ejSmdK+j
BvfKn9itenvm/ZmFBGnM8ZKJnCi5U7Dx0PEnO6LKZbj90M0QXZMt7TSZrpthmHZA
fOrbdPsOCmyCDD30kakriqcEG02JE2dOOckSO45F9KaJONkjVXpgTZ0OeG9bTYs6
J6qYIVIvztbCnuH7U5HigCWIbeSOkxaewFapawTsnX7H4FtNP9mjBVzhJrpKJLgN
5/WYbbTY80BWcsqdZVrwMXStu6KlIFl1xzQtUGQ6ADKnjheS4AAeRUIAtLcE1OPu
c/OwqjsCWMUIrvl3BYeMAOBha1vwUF0gEH5jJLVJJi5pid2FR4WYdY6QjzidRGdk
ID/K6b56SneNCZu6NWuFh1m0INnHYUSyL+1+Kq6fDyc8qrorXSILfMU7rFTb9c6P
I7NCGC0dYwo87twXtRaDs3xhG2874+TMeoy3VA8tB72QsR/TQupeVHdclcvCLN3W
Z8QAOLZrwS1d9ErO6X9GmYOs/WWGCYFN4sb1xXale+LUMg+szbiEuUsRjI42DTpy
aBXMbs+dLJZn0GjQq+5APfdd77FOMD/VgdgnJ6LGTxkMNsmQYAkSvkgb2Bj/IJ58
ppdjvD4h48rHxp9H/1nSpiswbUUDkXhRj1SrsVShME5Kz2naOE9vYh3HKiRhPu3H
hAXWZbqbg4VueAweDS2EDamOxYydhEYucUvdpzEP8bivUCqYMQumZcJ6G0sR/rfD
5kimqOPrv3T0kMrFTj7CT0PU8Hfz3v+fxJzGF/BC3AYVoHyOLgUjMgBAQs3CDUpf
mbiYBADZr/oPvjYiXy0Gg88GJldZ9zJm2jATRZ8uUO5auEYgvm7NfIDzVUfBoJEU
Ftn3rVs0YjPBaV/WmFhffmSW3D7/h1WezhV3im/jEfg0SY7a97jKgQqARM5yEhuI
Q3j857h/po71cDkrA5kpNKyFFJsl4VXZ8iZxOGubOIg3kZAhHj22bxi1kdrAypE/
YvI0nQmQ6o+lD5hhLUIezfbI2PEBGy0U8n9Hvd2CIzu+P9xPaujSSPvtrxwbHnoU
nWQzKfkUoZ2jSMgTTU//jCPqYXGfBunoyQeSyf+hG8HMhZjz3i+Jof+WzMvuqc1U
TdnUYlTOdciUr1M+d9P0Co0omKhHuvKnEa8HXJcL8mXJKP2MVtd6hPV89LbaG9lV
eaasTsCbiYPCPtOvfXaD8SqEG7QHl5064lETryZ0iknZ4bsyeRhd8MDKU/j+3uyV
INtZoRV/+Jdv688LwMeEByUKL5z7eNTWkQybutsz8wXQ7FNfH2dFYYntdiYj79zZ
oIG/kIOzL+J87lGLjTEsQFFXnsGOJoxr3dsMpHC5Iok8vOSd5XijL8NEDdocVgyr
kKCK/e77W6NyDFyEHCNT+mOnIebYhCsh+R0yU4VFCj/NCw6eeoqo17Tb/YTsMqk4
lIsYDKqmOtVAx9MrtQX4C3t39qyFNJXnTEwOyJH+RtZ00kheIbLLpLy/qFHa7Yzl
L1V53zPcS4NbzrIZ/0Se9vqAGg5EARfBkPvZcWO+3zWFs1OeoKY7bc/uAEyaQtmM
9wMWMNCHtSedCpNqrbP2GT1eMARsPRyB8GFeV8whkoUr6AsUf7fuVcMCKaxI9g6/
5b+eA994X784Rbiqu2oUb6add/iNmggehjr2M2Hv73DSojlY7yDtkC+pSfyOJR3p
THaKJ4HHhfxhPUDoCJaoGRmMdtJ6adTiQs2EAVpsROz0QGE5J0tTaTYZlGHtNqUA
zsyVQFIEtvb2iGSF1KOVzbZosT5EUt+NzeoEUTOr5onb/CPFSxc+wor0FJZYUSkY
lXgzOQiNJcWpu2w8jeOPYrEykWyg++MtGUlObNhkpwutBe9UpEUbgun/5diE9FyH
tSIh8G1xQGCaHaOEK1WhMEHAXpxB0/WznKo8IcbZgKb1euTlz1kyj9bld+b2/JET
hK2VgtuaPUifXvvidRE3Cy2C0VOhmvVTtVON5931dGRrHUm4VXaZJu88ERGQjNd2
15ck74PnFrOrmlUCfzPmqQ66u1z1YisOB7tAKIjO+FARji6QyHCL6WMlR+F3LfN/
pkhBpNsBa/rwQIwFbVQ0ED0BK7IKYmAfA/LFlHpOIOBSnqyX7CXGfFFyvzrPG6XZ
c4q1EgBklCKgPHTmUAyaRSFwB6qL1WkAU6i087ldEaVQnotM/EjfSVNwiZ/ZdXlr
uujEJP8xN0rn5DDWt4NhA9QYCqZ832X98MxTplsw73HBxt0fMs+cGyyR/T2PhEVF
rsYKyk7uVmDx83nTXzq5dL7ToR2bLVQHKzqDdaDKKhIokrizR/uev6FNo7ZaYitY
0LueX53EBZFkXTC0L5V/4e+8gwjb/sliEx0ISVGm9cNPnfYoXJQdTKKwQ0pint0t
uUktETIX/RDIWXMLkaPasa6DrcBbSsfpzgqoy2Xj5WqchfgmUebAYf3jjg1gStRS
5CAEc95AHkSs0zzljR1X/fDLNQ0HGMDGa+S89usuxvMFoktvIGcpb5nXSLctgclP
iuvMKbzRfP/LvWTeqD4eJfbMj5LCoZDgiWikXgHgZFKTcCZdeofjMTfUZucNrYxx
0YvG8bgGeotPcgmDnXOQwSCsFauZPjWlpgGvttf8D5+O+tn1uSK/HK7+M4VlBVn9
9jo6wR+IBd05n7VnKAI65eJs9TdS+OKMWvsUgkZwB+bj9Rrd/bRATisinjnUEQpL
D1D+MX4N+VjEsw6v6PcMt+AUfSuMj/KHbuIZ21dEmPYMznU0P3utG6LdjYxar5Tt
VB7go1dNxU8lbD+3cvcJ8qhXT47mQBTwZ9KXIGAvGEKg0qR5L2iTQTHKgiEf/E3W
7YizyIjXs4+04RSaai01fiO8HqQ5IYhTn/zGApC6vI1BM9AfpYoU7sB9MjURCuj5
QO/jQ/W06y0OcMlCFzvI6CP76KaQAlI5fjD6VMnaPvh06D2VjlS51lcIE0V1ryZi
hXfuZEKEQex4t/VlT663luNRo52buSGVsDRw3DCr+VynRkONaA1ov/14h2OzUVH9
dN+dJPqlMthngLC/PsyuFmoJF0IF76TU7iFuvuuhVko+nwOwe6Zhseu0m+Nqq3k2
1NJp6Uqrw0nzoFiXsB4RBjUMn/9x7YLjrhufQRgrRjtM8ALUMs/Vx8Q/zM7YHD1T
MW9px3BuCeArOCHCoLypiJIgSqukY8PE6UvIVF/nbgm3ObyMk4SpcJMZ+KPTLl9e
hl+WgHYTg8/PT1uD07PClcParQQE7RHMJ3h3M4DBmBjTDgRWmKP07FDdX9d4Au3B
7bGGsbHJKemPzfn6VkOqohNzMI8Gc8OnQKVhMGexIft/OLhJSgKaN9Z7wD3vI+Z+
m3c0ydFJ80m7SxcrGdRL9cTVVoVpf+5S9/jl+4SmDoT4bejg5nAi/2VSFQKCCnGo
n2SOgme3VTJ262xb+j96MpPq1YIGdC+AFfAo0F1g/X+SWl/y3qbL1vy6kQ7HOAf/
NZozRVV0l8rV8Ys7DQ8T3nUCIi0jTUZCn3eAauj0SfyWjD2aFHOelzpn8PPMaeTD
ymOxp4IyacXvG/zpvMMteKF0335wND0SyvEZijGCe85HzOzmT6+EHQLfHKfpu7O+
RA0UWbbQuq6YUuYIYIv+FXwDJJtbd3qGu8SgDHzOGkgbRp5Q6LAfrj59NuNNSb+0
/xKHlomRy8gdRAHOwoUsqmI9utXbOslBO7O8+FtIN2IaC+XYMe9pWNCOJ1+qzc9L
zSFeRct+kNsUJlTeSEqaWVIko835/8izdK9zZnKL1ixyjDihw6u8HTpWwIA79wTE
A5TRwh2hsIKoYGnLlgJV0x9PBi7udmnxUXpLmL3p/VI+4hcxYe1pnOHXSJUzDmQ3
noNP9QcAHICn/3IMv+pjG4zHZChnqpY/+uN69mna2ImjMs6o7FEIUNy6f4swgRUD
4nNpEquT8g/9NumtNrMVgn50e2O6l8y4KrZkSY3KKYPGZGwdPGg/HmSgmqEa7489
aPv+V7hcFiWfKEXoTmenurYPGnI9z+JHxd0wq2/dXCWQcHqbN26vMKY4FKfTVTyP
d6++jZWpB1IsVZoxtYJenTMKfEJG3/8qkCjHTAejAQH2bQg4axb18MDkaDem2Wh7
scI2U9g+CzKFFpH+S+etx6NN2OAxz1dHGHYwCjf3GJ/d2afXojL6WZfY8IShLSYX
HBj5ANrj7sM8apOA1WPu7+25JClv8sDSt50SXvxzuqQyqZjhaJn36/RyJ4adjzkg
6Z+zPi1zTUx3MSZIAAXgKkj+PQaAMGI1loON5aU3kx9xvXDLTXi8osLJi0mbSZrg
Pjt5lrh14lS3Km+tXlOIRZddVGogtIwujFu5V6hQWR56KqJC2LNsS8Cn43WUppqj
NtCI7EfMTajGGTliYrhArmpjv9huIRMdoMe6PGNzg9/K+c/v2DZr24tbGnrmDO5i
M3b1BFy+axlaar48ir0ay5adeqNfnHe80wgL+7QrDsDc2Xjtiyb2zO0NZYlgdizK
b0hxpOra3vH7X1x2qY/4FSs9RqVczegHHZ2FPmkj+1yZXP9GAAlz2ENkHnaiC2+9
GzH8HmDcZnzJRn3PHrWH3QRBk96I6Az1onmbOZAuJDv9z659SMifMoMJQc9yB13X
ziUEvD4UoW/qC/BDQMmw8oXiQRSy1Yjbxk0dVcxjujVa4T0QXjpVPW/TL422c6F+
fFpotLNCEOD/XAc5dd7gojvtS4JAk/01XjJ7ysmT3GkVP2+6nqMmhcSeFUZy3skj
TIpygt9+I0FPCKsVzS5UkR+4+Qi8DGC3gSq62Beu5Hy5YbBz/GpJeH5Q88EO+6UG
80AOjacuZGVU79Ym0FIvyfuiTFsfyrWrG8U8dIDms5Yo1ABoDsLSd8rQmA4ayEyj
lFHfeqoqY/Ibr7o41ykce/zqfzfqJ0EqvWXwpxjJ8zLTj+W2AEg8CvgjApEgst8+
BoIsLGVy6E395cCRsiiLgFZO8FamAYiO3ifAVdQch7gLX4syZhoZvfgF9VXarUw+
/ukg8GlP3hCmhweFjqoFgCIrvgr5JIEc/Pg2qqlj7zceLU/5Z7pGhFETGryKasz5
6fpgIYEPLFnwHJL+KrEnHUQnd3Lqj90d8OCr+MyUtBj7Q4WT5zE80M6+PgoAQsKu
sSmLXjUJP0JRIlkNqaFdl+lJlI6NugIMm/JJ4da1QxOW78PltKtInAxFw0SNv/BB
68HrnLpriKKK7m4w8j9y8HQI2MIGEnbFMUXqQSgqyrM1T8YM/4QU24kHstpxyrny
eghb3mu8tbribbP77xpf3la8gFY1xO2pwg+VYTQobncslq+8ADCpip8nHZe71zsh
PHQ9IpPz8TUoLaCYzeqkY8NLK0H1fcwGl1q5PGg3Exw6UOGxie99Eixek/t952xP
nXRI/o8eaXmPiBlz1EuQOvRXyw1ZecvnAlFX+cbVMc8Xy9i8VLLgeYNZ8+rXOM8+
OD+09MP3aU/ChmBDZDG+WsfFlZAGFVi3KfDpqOOsP2Kaxt2A/TR/OAXPRGuGmPmB
c9S7TrPUxXEFGtZgCD0/4WU9u7xbYWsqQK9daN7bIy4GDMAhmc3ULGEaiWnlW3ki
3bGlBnMOCJiZ9wGlmqmEq3jP/tKCXc21GURSJwiAn1GWv81kNwD06dUXtpgtYs3Z
BYMmUVYKSKFo3yP4H4gP89KCDeXris1EfDwDMHmlTavtj9P2fb20i5YfXtGpXGq3
88d7jrzheXAgPJEzopSWpKcv3h5m5uQk1MQk8MGkWQYZE7iTLCBPgVO8zzu+KRDh
hYAvOoOWvfOqbvqkZtG9UKESJhMjoZRdOQSw4kFeXbtfgDwqOpM4hqWvfSBlZ3JB
4YnUD+30xl/sGk19lDZL1QRORcRsuMa8ge6MCGAI2ZkCHthk9VE8w35gTn0rKCJJ
LVP5rpnUa8oGJkQu5Wk8Qbz/2aboYkgxbuMkTGYlB7TxNLHhyZZbJ6s5t5zaGSUq
LarOHM+yRgi+ut5QYr00nMH9rBJzko/H4unq97nuXgxUsXoMku/M7A1T64qV2mUU
sT/Jkp1syGujema85l/aUuPA78eJIuhzfRWSO/8gQUwNgJ1JN+Uj5Yp3K5HngxFd
7jydbOkH6gWaW60fto04+MOfBx3o1sZ/uzh/Ha9bOqv9ex4B9LmKZPuCn5/Dw+km
F+ZAnW/9x5ggLUShiucPAD03a8W/3XbMuS0HgiIGTsy6razgFhaQsJlr9ndXoO9q
151VyBtNN2QgA6lvTOQXm85dya2ZNnQFpnpjb4E8hSs4laLYLyG87It8YkusTaOb
GyagF00u45kQjCgClHBtgpZWfq5rYb6TKMMrATPi6VsKGkeQUPIT0kgTxQb75BXJ
yD9yITqy7Ms8PKMfTaD1PU4pPU85C+C7JVzni/1cyBYEswneeQUOTVQdR6zjMtZJ
9wqVuGYEXn9Qe4C7M0KzIVQ94B49t4NwxusmEMSQH5ZGvSUeVge6Ic1Z0/hdbmXZ
DpuGV2t0aB+30htDXCRW/462Iu1n2G7f9fUpIAPIbR/O8HJLPwmcMAo2K/2HLqJx
KpZRWEc+f4350wacH5Tt/+CmDPSb22os8AK5hq9asBk+s/i4haA7RDVdf7VT0CDo
mY4aUVEYiWhwt08gSezqT0MUsby/UOqlQOtbcU//dP3Vhp/mQqt/wG+lK8Gesrjw
HHnt8cMANhE32VZ7SnIuGaSSWzdu85z4HNbhISb6Gh1DgtkhD/vl7H7sr9CU0Yaa
V1a0anZ7f98ZsPWzuO19BTyz86oRM+USRfj8Kctu6d+zKDgb64CUQ04Q54vJDBxS
RYj6peuQRThR2/oqgsaAee6O898RVEyr6jvycIXAudRIn8eBORaYrFyCve0YkM4d
D0yoee6xgLDxW7wpZLyvaK+QyF6liobkOV4Qpxr3I3j99aii+obDeghgIy4kkvp4
7HkiLG/+nq1kCK7B1UVKmuKuIYgHH5xvxO4YMCcn2bZeO25p0LpsQo51z6DYjXkM
4CBmyeqsJSos8Ui4aE8nHUuvqizh5auaN3Gd0dvPSZMgvKA2hNXMsG8ri/wNKXEp
jGnQP+Jhaf3MTTJ3CT/W1fLgNs6TitVAYV+MNTp/0ow6MkpBa08zBOZUaIF5hpL0
2pqy1SYi/AD0Y07QNeggXl/VGeroDezSq2+8GiZaYVOrA6t6qxyu6NIFQeGvwQJX
69qGgodP3K1GP8ena+jcs7/8pQF5/r1kPfWaLDqp4KHKI/yPoWi7rh7jQqeSM2Zu
WXaNfDeUCAhX4sEtO14SBYT7E8KX+bvNRbwe4vEuyMOLmauwW0oXVtq8nDQJQqY8
u4MiJAEh0EsVU8BcNLgpjZgPu25VA1pI5hxByojSCRSu/Yj+KFD7qgIsXeDdCHhc
1KEj0R5IHI3qO4ZaBzy9kpKLjSaUeS1xLKuxnRdPQh1FnhwXJgSKY1UC7ZBNuFZk
k3u/0C/H444h2WSHN3HG4ITCN5VsE+5maEjisYEE37O2qkv9f87QK2znbqaYQTCN
M/+FpcFwsM5cjhY40yNFdaB/zYWVByRUiZmdp39rX4vVXDraMF4rkqED+wQAU83f
rQF8yfCZCBRfFBPVGRAXg5dhw20g18vSBcGH5n9cgUHw43zJqursmZ3a2JMUEsNp
K6PwbY0zirpedVdvDqMDd3UXu+EoREwqruiOswjIdjEiVw1D8moPWqc1fkZfQPGd
7cjFGbwh1JmsYetLvCX6Irl6COhx/MIL6JopGppSBNa/Xs/fhg5j6Hfd8L0vrHCn
8EIrBO00HtxchnpR/BFTFkkfkoqJxwZWdjJK0x8yNaVwGAAGAiJkq/tZvzP8i/55
EvRjm8TUqX5/m1nEis4YjuxtJL93YOwuXCgTr+ykl5cVFlp2vjVYp6OX6ToYQR4r
tS5+Pp9aEQuQ0HQuWVS83so6+Nn6QWJuSgpuHcIT7iNLPLd/7MGLUuN1tgvWy07O
tJjRbAA5eSyrfJYk2iPqLeAN4xHZn6qoVjxVeMfZcqqqYddkzMqpPv3BXFeCrrsF
bTXCR5U5Vlj1YNNWyELzhSEqAJyh2GGf2R97WKZPYbOFzHO9zTzOjlQxsxQZ+TYQ
mNaGwgDYiK888+wVxaGUiO1JWIKBxK3YQm/uKbpp/rB1y+1U8nTuqwq7d6WIFPPv
62sPWJ8OoHGAlYjwOlhpNO6NNYUgIhQ9Ry4G6nKk7fDiIk5tJwIemFi0Vw3PzQdx
B5e6SuwZ/JxUioVb5hsGhnNhPAVI+CD5pCFY+d0hFAW1OVKxnUvhyvhiuuf2/1f+
70gD1U/Hi3dO5bU+P1dIs1MqT3katFLTbFLNT7ZKKBnvZ5QSDgP61faEwZ1P2eNl
GrUEJLxd8j4QFpbpU488S6gdmks9U+bH3UUHaoq1d9hylHyZZbi+3teld9H7EqRV
kjhjZyU5lTxJYKDy1c1JbyR59ScgH5smCSYXbUMvRiExCdbt+tmXmxlMTeRh/c/W
u1WRtuYYix7eV6/zZ3U1Er/Ja2aM3QvEawa6Bd2SixPbepoqvQB9kcshKHabvZnT
s1S/eWhRMQE3cqh27eysyIwpolZz3WfnK7SnjMRF2BRdjuaMMQxS1xYvs3J7tKkw
d+SpIe/0mQYj3e0PjzbL0BMBVzoyYqjdjl1zxsUkbXPOxhjP+0CmMhtTZZP1JdHm
gJsD40EqA5Uunvik7jwsbIrand7CkMFJ9B8X4TdFgAz8zZ5nt1zhdq9h36Hw2WIi
WzTXu+sM9KI+R1vXHjeq2rShmXAnmn2RTuOsXbnar1Mid0duszm3TLrzPrGAa+mN
qytZPMnir7M5q3+IdDBdoEyk4jGyRAXPyunPJb2UhRxd+hu/QE3cb9PhEeEa8ERk
57aQmfRWHa045N1D6hMQVK1djecMlMN8Tf3qERFDjS0J8x8Ny8qpS1bI+7RKNU3w
UzDhAq2wewl/DdBWFwWtnJNrgVwYq9KN1lIxN/KVGCQ+zCI+WEUvLTCuzEv91IcG
sWr9Rh5i5GP3Fob3DO3+gt5CjWB1+oxBWK8pe6Qjn2K1at4WklKpdizEf/5eP+RQ
cBeLVMj60c+brqgEFFn8SP22pD0wIf+g8py1jsP7a/5+w6MMVzqM3ZkrHzuG4JnZ
S1WXHOv7Y8c1R2yM4tGck037OU9ZRLW1k/Zd8PmO7zuEqwx/LadQ86mjVwoM7fpG
76VcyX0EXxgZnxVLvDqHAypSqXlEeeRCnGYpDB5HjoHz+VrP26iUCyZfADnVpdad
eezzacKBJNrLuN+DWx32xE8CLDfZnbbOsuYDTrJLmmT5uqnVIjgoBsCiw/3CpHde
WnVo311VRKkohuhF8yKPAiILBrq1762w18eZ7LKTvQBUt/+Jbq6TxUTJuujsMwWb
hxg4jnhAF+/SRh2BLdaOG6frhaDR1SrXiHGPtnwhf9YcitvODH8CItqlm1cocR2k
z4KALbWty7qzMdT1EdFGCNNT4EuUk/FSutmbixzaQjg7+7rhGGPfRG172B1Iv5SE
dCMuzsjRkATpwKDC9pEqvel2p8Q+P8jYCAWLMEMVkP3qdlGEc66SWcGQarNj4bfh
4aFDKODOV5UKmwFK1/ZVzdN8kE0N/UbO9unh9WC/eRMA55LVrZt5F5+2tTwBQ6hu
ZeNQqGhigXXkxmZaoIQVEl/rNCllkNc+wOKHQMeCv4cDahvoOAQWa2kgzptfMila
mJgM8SAamiNFHZ53rdaSGM0dNVVcS/dJ7IOE/cHheHPkoytH1Jh4EKp0gQAGHZmn
v0uCwPxqW55d2MeSuF0EYTK9sswipzkU2DdhTYL8ywdmcNFJhJt/n3tHdPaCuVhR
1Xf/+qwloOI+9qzvsXZmzoVmUZqqQnlAw3TQDIwg473otbXSfBgtjrt3ZKf2akUX
rxlatJ0443n/b2ga6ACxPC+Po11SB97vJvItnPPmJU+XViDe4K1G3OZzNsZ4vRzb
w+VsAhGasdcXCwl1jhJPuQvgqzyWALtiHGtsigrBpftRi7ERH+DGWDYSnsihI4vF
Adwtr7wzTPuRT564aX0q8CyXEKr7KSQEAhMWHI+WdjL5zYdVGyEhL8noDxoFpkcq
EfTp1tAg4YZ+cDtkjyCpwTVjps9TObcsOJtMbWPWsHmoqnM5HYHOu9atWQ5PMeGT
cUgI7HhWRa/o72ZB80CIikbK1yY3Zi/D6CBccMU0+tjej0N1XVnaMCl6UwXv+Neu
n8kTiVuFrEtQmwZiOJYawICiSOQubcf/hW7orEk0EhyhfCq7xeWhU05V3N+hCe/Q
qvP8NfN19RsXbHf3rNoAxXyfCYlUkrXHOyGP2USJ4mGo1+mKa3nPdjP7Yg+SB+Di
O7R44do8seXd+UjI3hgaoJz8YYemZ9RoY4WS1s7z5V8Hr7sBchjeNEfHObpwPVl3
05mD2vBDgJRecrENdPvUiBrNknNYHc3AdGFWkDNtckUDDV23K/zv72EL9kQL+TBb
OGweixxWJOEcUJueeYqu30fxYeBUXVj9q0AS8ceOCM9GZVyLpXzuvRKdn6OVVHse
vIKbQlELdZgWxz7RBjkCfQZCIkS+oqfxZCfioFbQGlqIcKmvJfR/8185913bfGTq
sqZRVAU/E6SU8EcYB+qSgQ8OfDsx7e2c6jri+ZmmLthmMy0WkS3MSR2EbIOjjmZB
HK572PBH82SW3o/u00mFTHlfmQuZDuyhij1vi5QCfWTDrcp0xToNg6QiP5JWjt5x
w0W10vEfJky7+h0eY9z694P0oJfpBL5RadAfdnR0Xo7V0yMxhf6tO40kqOA7MseA
UxLQ84SUd0bCPMbhPBV3MisGGLJZjVlHHCCFYWWXhI55URi66r2MYDyRuojW0aFg
SXdS/MFS/SqAknHi5A7MkG2MOt+vLjKtfEA50M+P0jUdqtociAKDsLBpSDTkg7hQ
vOpmtcVjn6X2vzbLMQ7grz8NcxTVbo1BRwJAmrA/W/o6i+VE4M7T1fdd0WTE3fSo
dzYzx04BqvR5BP2hY1CzOdDN4HJYKwtwNkpzkrKk8iKMJKw/GqmqQ7fR4Ajie5gl
b6eDZQ3m+/FXedDDhTc80VCgZtoPeW6Gm451Mo7ftvSSp/R2B9ICCnY2VvLwk1Mg
AOqGFdQzbJ/sZC0+Iz/dlXjxJJhEfZsYjubbQNZ/tf79JtG3hUvvR8bvuNLO52hd
XUhpeZoMKiWO2Jwyx99UCsiwi+5aI8fjdc0HuMzQuTWBTxwEUFlCRSKcRdP6PrNc
OhJmow1vqUi4Q4TYUSrYG7Ttj243CpMbNrgQHsYXv2Zv3A+SFN/7EdA8G5OZgmdP
TgcIhHn9vk2/VgnRHqUZqKZVDqSnDHDAL7ll26a4JAbGbe+YmpT3bAuy3LJggduD
jSfwvvy+NrXgcxL16PbaPEDePACo1xgWZKGWik/GnmorqbQKczp3KZA/39fEccf2
oJ+XrpP9rymXJ7IIGN3KFlSKMGTTXYwnnC44BVxCOb58/i/DGVDPrVdsJnAajvkh
IP1vU4pgY956+XtXm1Qbfphy5/1bSMoNApKYv8ZFKfYk9LxOEhiElfkBv3tOb62j
dRcVoRV4S40HP4+SARARpDgxLK40hgKNBMjcOw0eIJybUCNPyWUJurISq6t+nFvl
KNQ9TE/UgL7Xj5O0SwUTPaKE9zFDc1TEk8y1YWyJQoaH9YgjzXVTSz/CVhmLp1uz
ubTV2S4dSkVULWDrHaNz4Xd8XakuGk/iEISNLeeBpY+uleCMpNqNqj59sIir5ukV
BBndSKgONvOBKzBkbh5DHo4VlkxNCBeCayiWpYoO2hUUhhqn90VhUQrpPVeol5JG
TtgZlDAAU4GLimw9vu4U27DSOUce7KvLs2KMyqWJaYaUvLoQWos09ZafNYiMsPRZ
FPAL2FRmem/UffLs1DSrQKcJCjnqf1yj+oJ1UqA/6d7sU4ftd1wm7lIzssaFxZXF
DrDNLowy3lDwisVa/iph8T7/JwCyAbIZlvxYysRdPGKv/6hINWpyduhafI7PUH8E
SvjXj5nhUYbC767IaT+XHMDOfIqnEC4nPtG+3N0RLKDkBz4YpeXJZfxBld0OTDGO
bEL8r3SJOWTS8CxZFCu5VIkBOwsNtIYgbBtxJhzCB91XCshjRYWF7YPFIwZlxEh/
CZiVfLlYwx6jOZyMIjvsJQ2fUiZa/0pyFPiWMpY02ZNLHcDj5MZn/4SuQE1I9y3j
71cMm3FmS1Q7NqK03slC9bczwZ/womCC5sfkPlXWdx5NFLedX+8YE24GkCyr4xOD
SYomCUhl92YEDeFFEzUNVZBuqQgyD06s9E7J91sR/j9xrv7vuDTpMjB3PNM/D/nx
72E0LWDon9CV4FdY3oQCDTl0JX1ZNpLIKHvCCl7tw54Bwl6HGqfaumFTU+hf9en0
sJX++aKIdAMDtoKrf+zID4PITj1PP7acMq1MkXqcEwWJ8I+fzW0o886Do/MBvnIZ
Jkr74TPVkUe5UZHupiGXbFcIXvkvcT2PSVYOtgw4aBJ/fVWlyz/pSDSwHW8hGK7B
Vz4BVC8wWxa6jaTQjSazid5mEQ7/joGB4ZA3tzVs+2W2q5JZr7Fk4fRTBjDrFpQZ
1n3DD6naezdSjw+r8zXp9qoqdSM3Y1EJYn1Brz2K9hpsSonj/gVv2hunpwKdTQQ2
TK1t+3HpY2jN/vkQcoVU6k4ODQpS212doSHUxOY0/FkU4GdUC4lVFVKCoeKjm7Pg
2Zd6435EcoqxOuiDsmmzgTdhmZtJ0iesn7TnP2qKkLZp+lfCwuiYLQ92y9pdO46h
DbIrHyFMNDcT6uWFbOQmGHl8IQSoJxcpmB+Ee8acdXpz9XDTNCApsK95SB90kHDG
igDSEEsLVQ6qfySCcJK+7NVSFdpI1gy7j+3C5k4YM571T51aqr9lJlui11Pa6rGl
lg1DOGne09AOHqgdyfl8K0rhbmpneA6yXznZzSgIAiJGgBQgmYc4YNoF/4Te5OZd
xUUKhHVKeYhqI/oxWE4Jv1+AvjvRUutWPJfKtVj6ZqcfVydKMyOL1Z34CpvLI/qn
MfP5Jj2I7p6BWo6OeEq9bKwNXZGH+kb71MUep3Ixih50BJmPhy7U8aj+fEXaLYiL
aNizd2bEbsm1K89MpVKpzEyN/dZjsgqfJAPZDhW7Dmhv4tkNDr8h29Fa0MGY22hK
Biu0oDrPihvvWdSfB6UhIM9sMWIhDi/SgtzeSjIbjuPFv6kAgdFWVioCdXv0vxH0
IzBniWdTbh6SZyYoL0lKWlfEI9Loj4vw/IqEqk69Z/9lXzVlpkorgfQfI8+YgjIA
3zzYQ+g/2u598Gc+6QBSL26Lw0ReYrcoib7Yky5Et+gLCrpjbcbr3h/+2iOnprcK
QtztTl3fmQfc8cmZy2LhCu4+t9BAISloceANZ38AQ5Uu/HlUt02dTl84qK1zlLP1
DuV1ImweFAsNCY5wIGHjSpqSLGla7l5mjJrSLCkHe2Z5kGxEZTJPv8R3RtTbrx7K
K4NTcXJKJcVixn6Q+Zg+IL+0ZClT/eJ2JCN1piAL0ZckbzUrXrnhxsFqMWQTtgA6
8k7VdkGkhmVNg9ACTOMDSkznRjws5bfDYSV5eAa05zl3R/SdfzQNg5DSU2lTp5W6
kEdNXhZUHq6o/q2btxSVZ/NO9U+dlQBta5561jEn+3H8SkiTpdkCWjID60coioRO
+S8I9b0bm79a44gHo6dhcjYx5tY5tsrgHapbhHGqP/mRpZ5ix7ygdi8HW1U/73Y0
8Zi9khUGnVFvLIbwD2YnPaNCQHsOq6cqc+LWaJxaJJ42wrhcFFANZ9TmTHRE2kyB
OnGRrjiSov4yPC/DPdb2vdnlx3H+3URVo4MH7H3ScGDzBjDsE1mIBhTO3bX5qj3D
StCz1JCuFh2kQLZsc2bNDmk4SXAO9/wJDnI+gUvait2FkxO7Sp2gdQIUMsDm30Wc
C65ffXI4wzYdLIjdcxrnv0Isf3YPqVby3Zzd+LUEfuuG0oNbJbNY4fBAy9fOsFYp
Du4OyvjtZuowAEZrK9cchgaMhlMCT+UM72ZV5o2Ep/nvIKta2AaMeppAPoZPLeBr
M/9QNCrqDzRFMgvHBfhlanbmsD29XXdLr7ElrkDg8rXo/bGZrMWvZ6xHW0GdBuJX
JnArrhd2TNi/nCq+BobaH23rmHCbGQHX8QzWXtIjgUQuYADlZyB+APN49J9pREif
Rr653ZHaQydCb1PcBy+x5vCv7hzWaR068GozTIZcekQKZCxGOlhds1uM1XO+Qgzz
Jt2Wy2L3p5F1uwkIFCLuIgbI9K48aGssV1/0Z/X0NlhPA7W0lCODrbb+fW2vR3VQ
EDaPe8jEGxLSc+Nomp35pPa/QHtI5qveVW1jeHqWOPjBKE/6ta7UnCybdh5C5ypo
fKo5DY+ewt2Lkt/zqIAw8W9r9UY7uJ21EUxiOJR5uhu4APD7nttg85XKt7jhUx7W
W5PJm0mnxZrqx50pJbojTpX7q4i3fEzYeT/bz/H9wlC4qWFtd4ygOoxQX0HpRJ1h
leLihflZFgR+9lVjsUaXSA/ZXR6Nf1pKOshlD/0Nn9sHoErhYKhL6c58Gr7jAy2M
CqBK0Q7z5oi7o9CUJGKG0l32AdWM5IPXauvNotKf5jFFuRjG1otox8zuFdy329zy
TMGFpu26ixvCH6mLuCKBGoUI+3p9sOb1sOe+p757+WxZP2M5ik6f6dGIJI9lmCot
k6eG4DAx1S/w2l9PJY227Ybjqy+tyM79dZry94YycvYzQK9pTSpLV8WLl3zw/GVI
Hz2kHCIU+/2lUM7COPWPfqACdd7tgidVCH31UmqaUmbCXotOuzBGpSkwGmXhU81l
TNz+SCv8PYsM7B0gY00TAxUL4jfuAiQjuSA1oMEYnyo3cDUbSYXCHx8VB/1M/BR6
05mttqpa2nb0fT5pkMX8U4QBS09VP6Tz0KLdpf3/ocnJKB1FqJHnWZa1F2tK6uTn
54JPSp7Jho+vhRUhYnen82THf+lJ5WL3KZpvyphM9NARXwQBblPtShhjGNPy9948
VgUk4fliTdfVViT4lGDin6mn/986e5XZFA9mXdCafoaM13QbvjEvQc3t2013Juti
zzxXt8KkYjg19LmV4gSB+X6Ay1vwFSNnrsHA/073mKlicPTSsLMVPcszbLwKyTy3
T+P/OfzF2itsT7Dh8MAsOsW0EfGYfDaRAgj59wsUabQ8lqpJCZxpbbcBxuq8r8t9
kPN17+rvG3LwvIL+jpEZR+Dwm8A0ZYcbgX/Ag4ZjR1Ats+9TogZHMEkRAyv34k+b
xRxp8n6vGwzIYkCCv999xVP0+slav404N92DbT++GpZ6xetdR2dzPJ9szp7I0IAQ
YsOvSPqoNQZHaCgVk9rvzf14+sdBzJVvnAZCwzDO2/gkWeWVxjaEuRss32WBmWLR
8WZpuTMoHyie2pHCs+wWecgnOgdNfR9oNhut3t2NFJL9RYqgHSNCkIkzmPYiz6yH
1WwKMC2yhzkgbCpl2QU0L7c//K3S7Z4nnsHX0K1U5lxPweB2HmskHAkNg1Ixf2ez
+SDMhd2g5xmVF68B/BVJ9rY7JM/+VEPxIgx+Q94R1UwUBTRTtDhVz1TaxUVqfe/h
vEYIWEZS8viNgoB/cVrFWYuBR1ZMHScxJAdhz+5ctNlP4zGsh9uqAN5N3UFI1of3
P6D6tX7ubTYYceR6MNUwjGgNDkhofMakUYdPy4mciPoxE4t7TdQRAueGwx6dV/h0
Zx46c3PJjvXp/3uJeu3XPHCf7X+4BFwsrr4EhT1b86K4589loHN7Uy+lGqLTlr15
gXHUvyF6PCEoC+6OltzLhvKmnz93OxyNJ1k0hRatJJAXH1zYWvEK6iSdnSMkuvJ9
rvcPYO9sRcryGBlmSxgJ2hEmrQl67lB5tJhTVQJtQsFMBAWq+WhhFgVBHh3wPWi0
33UpnKtB+e79HBq9rOVASXKDmWEkPc1+T7q5BAa5FhPUn+7irK06Dy8tmqzrWHjE
qw5Ae+trxkqj8eKo61UQU9MntU/hQzHM209cpbI1lL7NdaBqHKQ4d8VaXP2voWgx
rACA94zse+bMpc2/zt0fp+wy9zJSQhbB+2/gcWT/vnNpH8+t7rYQ+tzcH/j6Ea5d
5nIV3zZcR6rajF9j2LaEDkviAsNfRQ+Tt/RPif6tC6pHaiSiN8m/sbqDHXcp0PQJ
ExzKjkpJyAJd/1CsAOp+Ud27hEBPDQGaJ/SDrsH/5dzCW8aiYuPNsQoGCQw4l+by
9jvpc3M7jZazK8kYmymOmjzws8whCryRZdXwFupnvEwjjGEpg+Lxu66EvwjTDoET
Z4ssFq0Mxf+USv5ot/555PR+jt5gtlr4T7W7taZZekRhFoDR5uMSEpAp0uqYasPV
oW1OCI2SBH0Iq8D2a9W6LmLKcOrvE/A4iX7npYHxwJihTjdNr7SSh8iOsCVQSDi+
qGDEcqNETriJzmoXAiZLPAGe4DzFXezOU6V0qNas7A95+AgEHkoC4RUJtroIRqh3
dzQsRl5xmt6/WymCWRwsf/bZjOPJfmd6tXFpBGKd9CV0O9jcn+DYknxFoUHMqMn6
Vw664+c06QcimSXB13/JE8lbxq7+q3Na9uDYf+t7vQbtw3DzLxQR0iaRJWb8X8oL
NcAzXGIRkKXcYiJq/bT0S1x8ul7l9tMBlkiZqqPsql3/Dg8CDe7n9Dhr1WGjvjkw
fnfj+fv3/zAVxsTq48V6x/rLdzDs8BuSL8HR/EyDVN4Qregpl7miSzA9mAEawjwe
KZsu+yV/7AoOdbT4jBPQS/SZhUOADkSdsuAZld2KHeZkvZr2mKMATsObMkegleDz
njmiHIZQKGKkUoAS9et+JaJZPfHh4mhYgEaaFr9jzjC9CMCYwvDPW9v7+T+vp8eh
8Kg8nwNbEq5kRtqrKDvZY5qBDNi4nwcCDwwOIxJMF8Uqv3C8822xM6vG3Q3ZeVQm
6Djc61e1j7jZTAD5OBEG10Tz4d6xpZz4PhulIuMH3IzAruTCCbq0b7kTGcgn7K8Z
nHkT9Oa7ijxMqPP6jdIUb0uzA5UPV80Avl2U4hYbYKH9sHV0KsEBOXLquk4Zg15t
mbUk7KgZlBQrlSMY1noWPmDQPqtpF4CgkEj7wL9dxaqqPN/Fdyz1u+kGQfNccxKJ
nHU7Yg728t5pF5J6Muof7ybs1SBDVscpGrim6iSR/J6vryzlSc1k3hzgxki1/FUh
ysCGd16SrI6e5gPf7T088/wokqQIZe4YxKDzW4DVipS47270JQgmCgvoFWXLPyHz
qbdS85TNr0HariWWomTonQJWiptQ1PFGyjp4qilGtNwHX9YlvvgHdvfeF/iMHf7N
xF8d4/55qCzjdWPCd23UrIWgedKrU+I88355PKpxbG/PK3T7r26Bqsaro5yCATuf
YCpUMisUTnU16eDVa/6QSRlmEqzdBszWRYbSHE1HupqgUWqZ8EbCO2LbQR+bnE6B
pfR+6e7zJXnl2c0IBrdClLP91E7U3V16XN0xF8feUCIyC9EFmJG+GBvng1x7BbrE
ESQJWioAebRJXi40ipZDAA2Jcp9sN41ba44wzmrOs8ne1eM7Es81x91PXb14sFkM
vjFkI67+rJVUDSTPsv76nERh5jGX9WO91FqfSMIWCUAGamj7DPVBB0Uv+911gOCQ
hpVO5wbFadmmNT2HGutoCboBS2hwQEDQj3C2jFm1S09JGMYhWEH6+Hr8e8Yd22Bj
dJUrHimA2C9vfLG6jIYe0s6DUHShjxGIhlyY9Bt2Dffdnb2PSdMDSO0DkiHax8Bx
5315OEEfLZT4ItlcUWGC3fBmf+lvzu5qptkiVIEtiRdpOD0P83fUmWiMP+E0+g23
1UCgKgCjEYxSwi7cZXfepu6XMngZeGi5uvGkROF7hOKiQAGYvMyxdg/6vVdEHPIm
CWvhRHTipqmkK/xz0Zyc64ZCO5Idg+NHbbiWLUzMHJ2t0amnXr/9UPAfWl29Hcka
9H5qjvk52t4xQ5jwzJXzgyRVe8BNjUrz3o8uFWCeP8M5iLxZPK+WUJ7avu/T2FHn
8HWsI7JE+DjkKJUTZLMaYKwszdvO0FByy4LKzGJiJmwqJ6FzlHwiAmOAfMWepuGY
a9l8wSpG1qTgGj14hcfG8KTBsbKNQZo17Yh9t6dkdE+Ef39w1r6xtcrlPphZhXKU
Ych87RbE88rA2KLGsfqj85KWuQh1X+7Qp3DD1jjmt6mpEyKWXDauJKtONiE8LdTB
TIokQD3qezZLfkrDmbxnMibvxV5hmlt0hFLO/PR+CeyMdraBxN84bX7kYKW2Ma84
rgpzhVPNqpjRwEKYzIImtHHk2rDNjJdcIfycoK8VIKPlOMeuw1a9LGaPnOG3eN3a
Q5s2V9EPIQZgBFRWoD7EyD6Bn6KJPtdMSZfWatZUx7NRnJigsHZtTv4gOm9eyb/9
Vv0prhogMawxjzkbAJwqYP39QRwKijvWEyGANMZebPgrqGdq6p1yLMf0hQncXS7i
ADCxtoAtCIFjea4C0IzAi/bw3ROhzgoc2OxJnYAs3l8vJfWeD6b80gOOMNaqMOeB
3sVV47Lsaytf/JnQwVAjMaO0HVqFhCW2nisqGB+NrpHOuINrLBLTm9PJ/4aqBnne
4FwH1nEsPAN1QaruboNWl9JJDZ6wTho7Mq1thXSfs6O6iNJiYIUXsDRte1BisG3t
wSZtrTjmPbmj7p+ppbesqfX36oYErA2OchDiwJ4vTwCp/Mm3W6kDAdQ7bKrttX64
xSoB5OIyxkbf5NsPNsPR1C3PFTHusYdbgIpWoiaQPAeYKGORSMQu+HhhZXBRJZFY
DPi4ykuTzuMEt+unLH0MIU9OaH4bzTzIiJUy6RFFFIJ6iUViIa1AZrNELdpqoZJh
K0WVizpWQIb9g6BM98If/xGdtil45N6R0UFl05SgeJobS3k5rzrf68XE6sFdPsXv
lictYTjnV4DENFLArPhFhhJspEB0aEERfX25kGQ/G/q8hPPLNZ/LiMKxULi47s1p
go1nKZ/VqyK8rLjrxTn5PBwHJX3fDIHojUp6nWYP3wK1FhaTWNtJf52LGXVWpT8d
0qNGubXlmLNAQ0nh25OhmC4cBpHNskMQD15NQ2Q8oCqpx7VjdVxJ44RdpkwnCBai
52ppU14iWzHYtugqXCGvY/T3ZeoB3nhgp8mdWbAvpS3DX43Y8JOUqxxnDHYvLcpu
Jpf/mVNPAYQJYGVmzgdtPDn0OhzJXiia9yKe3rHXJ4i4YD3+0K6MEbtNXsKoNWLL
tCV5u7cpn8qxtUM8+J8hxigkRdbq+QTuxNylDF6J1430CkJPEr/++hohQKX3luIH
u5nUKgq24MmD3OATrMvcB4owf60/KXlFBbZV8paQ79jfubSVvneKKnLwBGY3+6zS
+OiUoak3Q9XOvuXXg2R2Hs0WpXQRxx1fESlw+8T4mOxgdoKtCg6TtpKFX6kgYuGb
UoQ6zfBs4lx2AKdLAV1ylZp1Z5cKGXQaWD/+HwLdVc7QwZQJWlh0OqA/6JnQVP0o
42ohgVDacFfCiVy3O7ONCPBvdmic8iY7Js2uRRjZUb8Ol9oSO06ijeUmSihGZu87
fwTIFZNKRffP7wQuceLv1mZGvJuid1q4N1B+bEI9YUVmE3R9sXRc36meumioUutb
FNpIH6YNncGhKVCGJ1LaO/K6jb6K/ygNkrd+S55GJ5qNJdY5LAY7p+IyI+qmN6+9
wy7Bg5BwHxuQ7CyUylDrWku8Z9GhYSL//4GSF3OvzTued6xZCU8LaeXoSGofqDQ4
065tE0i87xd4x4CLinvcRD6FzkcB+7wbDWJJYhCE2wxDotuMuHvYn7l92xUXFxrP
KatJtgcR2A9XOtR5lP74ZzDxd8KoTntUACJADDKjX2QJrv7VPE7DtMrcYyGaX4J5
I7u/MMP4sFWtDpnnivJH+KyjkwbfuKh7UWR8sGEtsyPlp7C4b2l3EgDJRn+ebB18
XqV5hUpdLHdUO3FB2RsWqWjL94yXj8FLNyvwnkflI2jNdCvD9v4RlMOICYuzryYa
qkdmglfrAoNshW5LgDgOX28PE/DjNP+/Bi55r7a+ro5SD2+LuegKCpRtYwouUvgT
CBimwQLyNRf2SCZkct3vkSUN9m2gVwxIX4n8RZFO+g7QjO9x3n3s7fzgHufwq6Zt
8ExjSpPCmhwLIvkig/zzKodsIya3awztupWB4uQFp5w9Tn87qjb6fGmDw+8YC/OB
rf7e4rT8aFROk9ko5NxJtAIVcNjvLrUmM2zRGrpHJP3r3oDWVbzxjcaVa6+zOBd7
iSVYki7DC5XGzLmzvvZ0eUCOqzl0bdOgqE1GfeASU/erirmbpIKh+yxdfkek9mLg
mSwwmL6HK6upQ4j2UCDHhKQiJsBAsEe84UWK7L5B8LbBAIQd1F6hcvL41zM5qiZq
x4E37wdqHhL0vPnD/udQ+nhowngpPrD6Wf7zXyBWwhgInkdq6J6mwjsQ/Yl1wn2o
xp8a1GtEtNri2eOG1MsxxrA5Zu7JFrrgPBGmwTMkuxgkwG8een6c+7sCp0oKHUCT
exHZcK+bwCtzq6SV34XYWnINeewibp4uoKs5GKKq7Xzio2PubHJtIn1xG9tih5uc
3xYMZeaYVhsfq9JYzDd8J1EGuksgWFY83nk3JPxIe2xvh9sZrRoiU1tRaYZw9Q4I
nDZH/zZD+ZXVWXEMm5j4199FqeFdKxUcg1UuPDVf4Led97ap71JVEBhPxJ4ydsJL
T3G4CY80DudSg2rr5PTqroAd29/f/H0+/CVA6uKGLVSOb7bYrU6oLwAf90KH6jFk
YkPYioUlWvx/ApRjQthrhbk2FgqZjL/lZque3rKcymzMd6rD4UqAUa7ot+YbwPGv
wxpGz38BwdhbK+vDf6Wn9/CQoJLbma/w6wxj//W9qVMqt8RlQ3Zbhuj10+hwLeBt
RtMDTBnvhBNXIKiKY5wg0CYc9mXAb1l7vZPvajCQM58AWG2A450vb1cl/zCXmyxm
QKnm5r4SUFnBFSSqYd9wL6Q7vTwyHRqgVEl9gEky3soqWzaL0bc1KFs9DeYS9jxO
SuPbRlsVZGqWJYlXYIcQBSIu1pUE1LXpxr6bMy+0n28xXAYk2ywpNWTfADkSngLz
2EKNeEx3zjEcvOCvO1U3QcPm7xlUpQ3p7FEwavwJF39MNQJOmgk5lNi1LUYgbHuB
hqnNjj4IT4kRNidhWQtQfOFvlsQPWGZDWgUi8HYrGIiD8uLd9rckCmaWyYri7n2b
ki0w323mwAHb/Li+Dy+CnYOx3w3HrTGTgCbBLwqF2Rij5tEHjgLV4dg142F35VQO
CqKRui6rwRKop/zuWNEwrKABCFsPLJ88LB+afsA52kiPBnvu1lI213H6jcCW2q+q
tZGdlZn4CzeTVYr6stbOFb8lWetYjrSeCZAMYiqGH+vLu94u7v9V9HPEXKkRaWQS
vnkvYwlglpRKE8Rr7peDd/FHzsjBaKfY2CXpTrdFaG4upnBgILcsJpyJpSau+bD4
ASbhfNMIs1x0r3j1015UyzHEx0pYB3wAt3TbyLc6EfpmE5UG7u5i40TwvMIrIS+c
eJc3lAs5GNvWCjzyY1zsKzzuEySaETyLMGVtc5KIc4mYiLhqdRm6btkXN5nMp1A/
KjSBF8xoLk5sbcL9lZvUu+UOQ2N1E49NKeUfcbb9svTglgwk1cgcPHnnTpwIhVzP
I9bn2Uf07EIQthbyGQ4x8TvadJTpT7qaZb5TFPE9Fz/cLC3UwNJgmGlNqCvVJWpU
qCtS23Klz1+zO/RemwZs2YF/1af9Kr5qQ3UhD9F7RmRcv9HwkMzdj6JYZ8/pe9WI
mcLg6RRPA8tFTxlwjxgSaUGzEOAougAXFHw6CgNzHe3jGgNUVSzZFe3qpjscTsfW
Rzs5qq8ucP8gTaNcmSk3NAJ+GNhqNpLGuS0FJY6Nu5q7xNlyWLJnkGr5qvPneff4
nAtB7HeTodzIiAK2xmkqxdfNQeREW5puUJQs7FObm4+29/Yq0CsIvIfE4x4MezXN
NtrvC45RVcn7z0Ftvzl55QgA+vB/KR3RvzBeithR51BRLZtT09nIWgLWD2GTuHZ9
aY9yTPtKOGEQD38JYqlRlSw49wUSeYwncmiyibFvL5LpKtFPAHabalP43YhHdEgt
ePUjybRL5rJKozaxVOZrxmZWt0jy3eG1Rl6iOAa1tBtMAZSzmgcbIchHtOyCYG1k
oSyxte0U2ex4IamMusQvKZEa22IclIU5DLjQH9X4Tvfdi2+oU4trIw62CDOiqe1k
XTcf/OOXGijr1j1nXOJJoEIe6XOdRZDM1h4On6m21Tcn2Qno0uUFVAqyonX9vbXb
jm5mPwbjwOp0Fby+8EK+dCLVjBPMlH4LPEu52CfDDyvR/yuYFtABqjXwn6Q3TXnd
vo8QSVGuEJhQuzh7PIFeZzIAx3Ud5p18+TLDZbGhi2184J9OPXzk/VDv2hBH5M+R
JBhd4NYnkxdDX9xZmksGRdPn5b/V9//juOy/IB5oXoLoRXBOY/P6KMybNlxIxlHg
h863CT98/HdJHCzm1lu3MLXRtN/0F1Zq/bKZr1DmLQMBnKy1hXxaRUna9ZmOL3WK
aUm18+Y91/L0mDGug3R/DjAjwCObcVj1ohyozRljotZ5R87diO+oEASS4nCKIphB
+2NHYVStxvZp0laHlwSWcswXLavGqdMpvyeIjXHe2kMSaBiSH5rbYSAR97Y/ZO/s
tYSv7c34OQbsR9G3DsuflgmDuKCKFto9uYacjaEWanyDZhlJNlxb0EWhja8fuJT7
JyZpqas6kFhe3EYwHwaRwKqbb6Keszw8XMxI+ydM6RJoV2VTOgCzZ6dVTdR0vPGq
aIQGZc8kSQxGalH14zqSbrW0ovmHEveQGy4UljnnlwxhbFyUYCe9ZlEZykMlWCx3
wT1arzO6q06yrIlBVM/9p4oTZHJW3CRv9J/6nk17OBF1UG1gpL7f9rWwcbf8xNxS
rTXjGtUimqJe/J/69sp6HSkFjM15JfcDiYa8tFqa5IkIQDd3BEJfMTnLv2Ax1XPA
FfSZdGtnOIfgS3bmS88XqNt8RrQ7a/kCTzYNeqpUFEy5lapNhwQQtxHBA79y/+vh
CK9Gdtzup4nwuy61T/9msp4g5qit52ZRwGI94UQ4m3mFrBYi93dQFiXgPZilLu5G
TJeQoI1E5X331uSQkiv1plhvbXkt9psQTMZpxzJCrQQFTmYXWFihI4TFompCvnft
Dx9L6NWhvMexyJ8OnY8g7xQie3X2k8oZG3wkRpFfNLgTLgsxDC3rYqJXGkkibg8P
Cu4ciRUJOF8BhjOQZE8A9kHuCrDFgITUKb7NvXmyzqhaUdBWXJHZfxKJ/0VRcSaZ
TeQ8pM2gq1RrcQLpGeFFqYPtjA5dWeMHwSj4LhUu5T+Ar/HaqfLL1MJT2pupsQmH
LPPsgH7tXmnC45DDxKePkVRuCe9tRSshH1uAyDGcfTaaHzUwK98BJnLcOdkO/1pd
eXTZdJr0xFmEHskmOIeItfo1wH6yZ/VDtxKFeUjO8zf0CZCMRpOSfcwPima9DyXC
6Tc1FHktTEUvrJpA/vuzAqP4aMrA2odYTovQH5xnrRFoWyPW7CHiqpd98aT8T+dx
ZkYRoMkj3aqzb85h2rEu1q5ExzzX2CUUzWpE7rM7ygedM9kh3XYTJxjh8sQO4Bhc
25teTj36b8888Cyu3zwzn9FItYQcQA58MUV5RC8u3rZfLavxv6GL5Px9/QboZoQP
m419fgvPQ4IQG8ECIqjOQ3EzUX/2ynEjdmOMRjAlaJPXzvxMKSrQVeZcO4IBN730
DQHR9pNGkEJDCddDZ40MaheaW63ntd9Ynvaw7RKxeoXsIBSwdMwSKqdXmeTITrS2
bSFNruqHgirdIkmlTHFvwDcVQHG3c6mcGL/I2L3XsleFKz7FBdiyVKR56x/7EPS/
I+g8K0of1KXPJMOcYFKo7mVibQDsMFAtyPFC8OnPd1l64eKIY8QLml/9NF/9RX8o
cmS4LcR7y2R4oOljatzfZ6PITdVC/E9FhFvIR7h3ZR4OaEWEvx69XkR9qMTzssdX
S7cEo8RYHXRgVFy2q2swZdqhC8Yu/LlNOvbNXRdbX9yQbnDHbG1JQtycm+N7+s7m
z8rjlzgbtNFhyqi0BNiiuAQukrXZdH8P5f79n9GSc29ALXNltbrWPRPQRGDfJFKa
/EfiAPDt3wEK8fga8zra1UTELsRgJpwF1b9nyizujhrM679rBsZWPXPyJTn1tDyW
nWHmZ4nDir7qCnh9p5r0eBZAQSHAfy3nhaXjsZ2TFV50nIjRSRqvSE7I0XSHgCLv
J8Y7HUg5hpQPTCISAj4PN95KxBh8V3c8lqn5FCwMfXPykXkkWMOSt4OUg+CWgTKZ
V+CxkrXraLww6hx4G6s8lV4C/UuYbhjqpzoiDhKbZGy8KXAdjLFBFD1OkM+5y2HD
5y7tGdSVx0Qw5uvbeFB58wFvV5pmzXJ1gfeHULGODCVxcrmgYKzgoHpdCUYMIIH4
wECkKnb47chJgMFgBCend4mQf3T1oD9SndS4/yc6YfYY3A2qvttBGgcr7zez6Ijz
ZbPb/QpSg8FWYUksVbikloAdrZsHvLwDc1b7qTCWg9kivIwBwIUiM/7azCaVZCKc
6ny3OGWZf9ZSLYbIQRkgAbrJ/5QBARa4ee3xf5PTapwWYH5eBy6OdCWoZpSArtpx
gCxtZlCw+EAoGMWs9MZqa420P7PT6GbZLzVfIPckvVNjgvB5MW77PKvrPHjLviqW
Evj7a44e+xHdM9PvcSFT6GzrTV/ENLZO39BIFRSeAWdU6Y1bq/a4zjTnpX5G5Q1o
kDp08/RDpanaFuOm+yd+yADEiW4VykR2YoEG20CT8my4ZDNuUQRCd5FrOTHXgVWw
YKlEmZ9wuPHyA4nCrHcbNAGRlDJM2vphIZ9xQLUQGpm9lbbON+PCOSr1q4OQzq4q
u/KE+MWKLOJgkzJ42UZSjzj4SoGGhcS3pSc5udOUmeDkoEVdnKImfV7OQQkTlFGG
o3l/cClbc/BiDNLO/qjWBvI+v59uMJ+/pJNZyEVFbRx07G84YykuA5ClvTBVdbAH
zOXvu6nDS3M3PBbpgkSrLuTQ9PBrNKeJQ/ICOUixzVPWQvhbKWQAbelI6x4nz28G
7LLA7tANsBl5070rKZm6Vbw8g91L6S8xw/tclbqBGsD5F1h7+uCw8p3wT7Hp0Cq8
eM5OWxH+6CSjVj+qbBnfobnzmVmaf1o9LIE4c+qQWn9WXJh0Kobj4PoKEuKkLJhb
/LIxFA9aOJeG/NtEhIeklTvkKIazRxmk7v/YHNxKwhYV86QkE/yQQXYiO36cr7++
Yc+tRznBfKpI/nXLWISuf3NRQf+jIejArd71JeOODR9E6MmlLVHQVjWEicHVPz3y
lNHL20dPOUEPslpXfi33oC47y9ZzBGQdbyvh6FkG2TxBC6M63VEOvaxK4Dui6nnr
fSg2TXimeLYf+8lFglvzwvDQX8PhDL2e33krHatcvAkgza/IB5QuA9BwJMb0pdxA
F2YJfNPsvrxfcSG1RtiUw61qeMsqOZTVN5NnUBJ93Ds7QEwMb8KQrXqQfeOCPKb6
SJbN7kHgevZym3lJiqpJhxq8FqOBCjs+PS/MXXkRS0dCy5zPynFTuU46uFvXgdPf
lZ4kCHuH/qV1xvjOuDmNDzMZ7oW4K2FImB9xbcC7NpUVHCV/ayd/xgLAgzEKstlW
kkhzCBEtkUXR496sPWfyDTWKh9lWyWnhQ+93LJC//qM5gm2+hYp9NJuaN6kzn1+N
l9vmbTEeDb6PZITccZKPnq3iUBOocaay7luFnD8A3txj33xD78qO7djbbqOOS3ca
V0vY1/+16Zy2FXZDMgNb6+/RhZEpYM3KzdHRXPfFjYVnqFup5XzwGTtO3zGiChce
ynvw0Rq2hPYWcQC81Cm3PYIjiL1AoefSIC+04v8QKJZBLD6me2McGp5g7Ii/FCNX
SZIqaceHbGuBvQHWx6RxCDbeR3sK3RKA58uI2cjuNN2CFmL81x4hiQlG5gvENtWX
Vgp/Wu+RR5S2d49t2fP7jYEf731vYdoTNSQJaal2o3x5rcgc2PWAi2YN8G4IUMRu
kMtHG8ZAvBeROfb1CqzjMuZwBxh+FH5vKaCz9QKskC0Z+oB/oWbPYjAz6//xYcPl
uKnIwM+DZQU/v6QKIHe+ezLr3mxDoqce3WQWSZBgbQMzwGe3iuQVOSj7fbSO5nGT
QqPO4UAbiT1lgGnGSGAyNr/AdesoDjq0RbA9HrYDfMAKrWgRyxyOjhUkPhQJXg7o
OlZdghxrOlUBIXdq97sFENj3eX1d7l62XsyVfr+qlDHUTYPJMC9XGZbyXI18k5X8
P6j/HSI7eUr3hwI6BlLOjyztE7efDgzsBVCkyAG5V3RzmYYHGkJ1BYC4d8nkofb4
7GijkTpNx0b37gEFxtuO5cA65fQj6sbYfFv92ywZwgtvqYezHii+zcSSUrhWCOVI
XZZdD8bVZVo8LDN2z/4zuVm8MbQRz9nolGR4nxq4FfutSDBBWa5YLBbJv5w6+7to
DWSJGihXKUB46zrANzqYza1xjbM2s3tHlqWuOJIJ8N4p9KMjrso1CMiB4SvHu7nj
jyrN2ekNPvudDfn1x8rk7ejc+yagWvmliqrRNcvCYaapFklLRVlUH/EnPDGzFFQ8
u7TuJAssUPXy1h52WswUQzoL4ZG7bs40plW4puDB8L6RUOkcTBevhbkUdP90Oe9F
BlGRYktnBQJYClB1mjS75rCOrVasX6maid2hwts5Zoz6VoDqPGkZixBwFgtFmcyT
DNz7/67IQ0y9oS8+D79pB+rVwZtPGBz0t20N+jqI+XiJL4HwIqRiNKWAh5YSu+WV
zeIgEqqrSeFOyiQlaj75c4tJ/s5rKA4yDKAABq2NJRdzhgr76cqIHIms9DgvwWIx
1RHnuWZ1z2HMaHbmSwOstKEUOrX5VN0woAu67v7oo3qZPtZqgjytoELxyAzzGQ3F
K0SbBq0az6u1ykBDox1QrZZn+y6rCCtFWkqhLEwRIt9O6sFGFLMx+JTvcCnE422+
Vn20ERZ+qv3wbMZWqT7hP7C5541Imo6eiKWrsQ3f6euOndvCbqdmg9nDcmaeQfHy
JqATgHoLrGFLVGqCCavNsOE07oAheSIALOFQeZl3sLNZzq4lYA1jxGKH11gDJWgD
wdZZhxGsErm/xoi6sqZ1Z3DBfTb2v1PjiKU1BzT1Hq/lqZDZjLEodFRanw4IdxOf
KXWTPk3WsL3nSo52fR+jRnKXkoKWbiTCA0+W5u8uHFNxkukjQ+ZAifkoN6yO1aEW
0tSpx1/I9ksCbHSDZT1MHH0TczDsoWgrkNRMzWK94UnAR2FMyYsDRWTCJr+EpNNG
2SogLedFt6b2E5EMNpg3WJAVShF2BbCDCdR7wOmelIyIkKC66z5UvlhVECO+9mp+
Y68uPIBFYenUGXiH3sba2o/xJHYikgoDiIpqZL2CSEf3vso2dXGYm1uRGavaGVkQ
WM/jLUyqAatAmlQrv8QKt6aFxR3B9TqNDfK7of0bUqUTgx/usEDyWe6cdnSFKno0
OO5xWofZDfJ7LsPwEi48djFrXCm670SMCAhjLkcCajKKDgu1j2CAxBoZRtH/EQ2h
nNpBeR7bfSNaD6cDBm/cpgXgcjWn+E6zkzNvNs/x4mXMTs+6o1wJi2XkRYXfB6AT
L138SLFBL+Y+y/mC4uU2yDNsCS+pVYFwClWzbnmts5dWngqlIA2Pew58AobBbByW
NYZEWbeWaL1/L3ygqeph1obPLcTtgcfnI2J60v9To+pop1Urn+xAveSt/ImUXrED
BcAZW+oPIDv2VmS696XDyBC2HwtXE3btYX8bUBVkLS6RB2qRDYDum2BEerHa7sTz
bWJOwc38A7UhA77sKYy7F2FcbZKca6b6Uc8xIHu8fEv5xQkyu2lRZL2HsnnON/V3
oSieFfhAThpC8jwrvXNOLt3cdEAC2mld8N3gkKX6kD96bx6G65rA9GRfU21bsVni
Piem+ZX3heWljhGAL3aGhLnEM3bIq+N1Wv7hXPGoCRaeiKzC4dGy7S+dT18WNtj4
BjeauWGkKt25xcD2YIdHtoGeYBHEzu/bK85lucrAEM4gK7hBkxARnIYXD5SmqQr8
hGGIdWJuQu/7zt7ro6aTSWrTPuop27eQJLZIsAct3IK+Hv+T5hqGVqidknxdmMIm
0/jpc6zIq9/uPH5cJL3px+NFVNHKFuqrkVlzdGCxkW6WYR4r5tWUxyf11JtmLl4N
l8abG2ohYEas2dfVt26fITkH7if6TuXubKLPcZVcmiymv5SbaZxlEizRfhv4dJMT
9QLWXHTcJpAVjnDFwaWo1luf7iC5wXtx1gWWHVcr6FChnrFqy+LtcNM0d2eBpBip
dkfzoEYK4hUa1DOwQVNsv6MYiT+5ybYc/K1IiSW3H30jP6Kt73aatJY9p7CN+bV/
5LfbgQQktL5myJFZtpDf0Ldg8UpG5QUxHtFTE9OYshlKYr8M5bhWmx0vQ2InQRUq
qUvIh4uOs8MM0itxXBi3ES9Jtv42RWhEl6za36X0zqgqHcQS+O80ZXrjUNeBJWRQ
sbxB/hYPsCkESkwiSn6iL6cGhtNChcdcCkXWGTb81zaXcLk4PG0DWPyCsNBGlMfO
2izfNOMWm/sQYP9dTBV0kngVCOz31b6JWIclD7+lklJ0l+I7DAnXWvkswnbT7xrw
XpsTh19GNW9fdK6+nbPmCqitgO3E438cLWqaiBMhWHLEdCahthKFK0IR5a13177d
4lajEu1rtLmG0CQgXb/RCY4rFQyU/sA+sGZABGhbirJo7h5R374dGgDVbxC1GxiZ
ZnOXuoyGPAj7grlQN82C8Vzg9XootVJhCx5c7CtpxJ02qG/I+IUkw2Dv/4yZpcPC
YEoI5jdpEKcLKM/jYpJf/4em6Df2onF6JLj4550TTFlJENFmgWvH1bQd7yPF+A8a
qu2Xm7c/sKZfqUkPA0NLbzpnJeDSvjmD8i+eRFkITgj3/wrAh9lYPF4J6PYQrTU8
EXrKHkSh5BjrQcKq2kYMMe4hDV+2O7r9BIFTzknZT/aUT2z8auhEC3PVCIIjgWlA
bTthYQcXiW4/5F4p7l94p/inGFBURW3s/qNFzujXd+Lu/Yq0zBEonnfN/yjVTu4/
eIwJgH1rAV4YI6wAZuVxTHqJtpHS935VpyYDLMTkPkv5jOoMJ8x9+Wq+kPDcE7cn
YRAvo2/aZ/0jKEx77qeKeWcIbSH7ZFs9RGADjbq+e9PpvTXAiLi02LQUwrXPoHl1
fu2lJtHKqjB1d0RVZ7xz9bdnuELi8SyqlIRMoJZIxfMus+b6zkAexBNw42xgUzTn
B7YVmkv+zhCz59lvAGw4rHBGUXO88u4sFm6DeYZ52Z5F2QvpzbYpWfXgvmxi3+14
x6kpLXveSGBsuG1bLQ2RlVzX5Y6vQSvtWFTalPDryvwYS/loqy2mlIw7PRuoGK8p
QFRc8Ag4pmpfOL+oXtyvuTFt6YoKlBjNvss2s1LI7FkuUUA0yZdNVT44sOl0EXg7
nx4/YQagVrt/gPxd2Kig61e659SCRifRAm+EAd1Q5Eq1jU7IKbrX0pjMokBPeAdQ
2K0mSsr+Rtc3anWFtZ3JzVbL8G5MgcixdH6yv3OX5WnNCkkm/mc72HVn9/+oCtRl
1/+Bm68PJgwWPbgNlVS9+qAADxKdhwuVLhKUbgF2kh8Bw+gdVthlnN3MgNWJYI19
NYIAMH0kUqAwLdDuzIkcwl/q8ZamCZT3dG8mJkUqPrQ2KPK6yCICprEstguaBEv5
VeWACu643OMLT1wG9tQKDYQY9RXRnwtWDFFvAlfq+WVis5+IvxFuN/VrgaN7qKBU
ML20fKdSDZGFgkmpxKlp3hboISORXtX002DmURYxQgnYKYK/kcYC0pAjNe8qoWP3
vrJvQ3V2AVbL8oiGYupSkihBEtyi1cGJfrHIiQRYcgeZwdqC4rjOw8m0UakB6rLt
Njk4PmJkZr0F8kCLXtIC0LnChRh07MtfbOEqgrE+u9PwJXXqC7zGWZfX+/bCujJ/
QpvOvYElVi8ieT6NYnUTnvtHvTXqDEYlAGQdv3CAokM316zUWQ0fWan68BcdaWXv
BPTOzVk+F9DFw+HW80/f/DWr6n2N1Oo/IT3Zi+RL0Fh+6hpMnbS1HU7Ci0AiT0kJ
k+AD5GlwxM6ZV0HHBfBQthgWGzHOufChZSpj+jjz6hx3JfUCB8s6ywwTxefdqqZw
MW+xoQecxBQHxfCTrBZNOIxMltEg28H78zUXqAKi1XYkPIdiQcjOyAp/lv8k5vTf
njyO7tseALzgRfMeWfOGeLRQUp9UIutxUpWfbpTm++Jhy/YMVHOt844sX0jnYPuw
2O9O7bG0mr8KLyLIM789LgpIuvaGe2q4au8ROfP4EiRuhN+bOO0M+xBZ6S+fA/mg
bnDLTXLt5G4TrXOWXcIpdsJwvJnE7RIFobsFAGIAl5Ggx+b3aUEBFXso62WeA5DA
yNLvUguU5s/AHzGh0iJXEx/2dsZbCVucEMpSe8tGJ//yycVOhkVI01928Qn1IDn8
7Tnz2bCq3eSlneUUlEXCbhyk8JA3QWou42lfYY9P7BXiRh05dzLNL3UWvdpxYNAi
ojaSAL2SFO4ObLAY+C+Keee4OU1xIYYOfjabh2dMFjlllGsz9+0JCx2whslg1hzR
/JvA7QfYW3UIjgeJwrBhaws7ytXLohPsODASeVAXRyu7L15eLIDnpZ/VaGvq6Cmd
peY1usR3D/L+rnD6B5bjBmryWURWnAAvAoGFYy3ZxckFw2OkB5l1WqTFc2Qf5orK
6Z8YhjuyJSETMpmYJQXjOyeHRp5HnYg+OSFYLDw6eg6YNU/ewux3Em1R74QsqEvc
udT7Z0DJoCgQDlWQCmyro2+Cnd43MNOUO0VgMDVnOkLQljuc1OOtogmLl0SmHzc4
jRRbgTbyB31FBhRaYseSamFd62/E5jD+ekVS4Iue/IpKiSwAegw+sVMtpF/kxHAU
Wen5wOR+t9dAMnQs+tHDvyBGlg7SKRCLKWM6NuwYgKp6NdlvZ//wTBGiHh/BvwOh
BsC3LW/dV9nfQsFbCDZudYWn+0R6Fl3kBtdjP7d7nFiMoAlWB3cGz4WnAUWZYYqg
2uqfNL2e25TV0j5hzjt0csnyBw93OvQFyE/KI0Q4//EmSQ8E7jd0T4Pv4qov3TSE
bn0uBxkgrPGbCkOfi/0/GdFzOLxwcfY+Df+IDTm04e7xXM564OsL4EtKCM6Lpfro
U2p/6uWTw62+y/WWPtZk5L5KKJXwxhKK/CAROyZuaKOU9MSiCNrS8SH2TYbKtlzf
HWapproFe7ngDw8lx/JsY/fyp9Iqh4UIr228VIY3mc6xfhUjVBnviNkTdWwbslbb
0Dx2qWkpJMi9TqXI8A5DKiFEYRvS9pt1Ipz25ZRVk6QmLXN/U9YjySe0CfJMnUqr
sxfuA8cCQRT1ECr01whf0O9D1m4helBfSMw+5BkU+wwsu1jBGh/Pt2sY4xHkE8O9
g6QDx+B/zWhlVyDRclRqoLJ2Cs8Ikt/4jpnmVzVm/ed13U0+n8aGFyT/NmeEX1Fg
OxlcU8RnKCOQiQ4hgK5ss9JfQzPCbZmm6ZHyqnKPjzbzZRCJCK+yfSJZcTzr0VoY
rJ/5xtsGjfL+PSVZO9UjQqjsSp+USyaYm8YZRmN5Ue7QodKowbJ6q3n1AOZk/FIA
3wa8hTTVZHH5BIhT8Bs8OWcrmE27wwAikYfN2DN67drblGZDP+NfDGtbW7yVD+jZ
xxRPoXCw4l17XkDvSfwYZRZhrMUHUI44mrciz305wtJLoDcNGcd0FAY0em0gF+K1
qeGS69H5mjM/DFK3YKPEdf7IGJtBbFfS+y2WB22v1a4c7a8ABbImoYdv9Kq9lIi9
abiS9RBlUXMWSvYMp3sLp6wO46qHAJRBc1H/coo9LSxqHnegwFATUgzGt4ntyddr
yAzbkYC9BtYjdbcDu0/7H+Aa2UukEY4ZfmOmgeZvWemwbldofTz5T1QRGiawJLdl
2DGgxcES+AIx2kl1V3lrC1zj12cjuab0lZy+8U8lPaasn/TKWfluqKEmZpfZrsE+
9yE1mtHlTDd9lnqs71FbRskv9PQYmaODzsKuc/7Ai589Ha6PoiTE1ueFsYgr6SZI
TLWVQQl5lEapeJ33Ko1TPBob4kcieC7QtUkYdWCcrW4C2Un6yb91ttiELF6LD2e3
YZ/A4z77pL26t3yDmJ2lJmTU9VpiF5PtRQVaG8BqwPzlD20uX2f/EtUHQsO6mMa4
iiN0Aq76M9gLgx+MNEXY1UVo6v4b3lpMyqZT9pJBX2kRBKHxIwyHAIbvxW7do1/h
Bg7GGfnwTIwXPCP+t5/XLPWdwkVMUuC4IBZiNpqn2JT01Ou31t2qhgZ7w3JtFsAi
I4k+Tf8MH82qkBizzUR4AaRXVEMhkyrGGSA1bNc+VLM/MTv3UTYcy6qYCusFY0K+
IA0quzx6GlalG0gheroN6lDSDxfRXkNw/GLeI6+EeX4Ts0qiYBl1DzJU+7MdNHmh
3ekiOHqJ3s0FaV3SAplBS5W2cGrAducQ7vP3qCb5w8XPYSQe17G0Jyha4PvMrZZR
lZnYc+tUzBOwQVHjVwniz8aEKmPjO2hgjS84Nogdz9r76Drfk+3liBShfTYFFY16
iF12RA9iFwK298jlxZe09sVljx7b5ktyzgfxuuFRMtbYrP9bFLJpiTwvjuqeZo3E
KQKfXYO3BwEjXW8YyBOpvYhpjEoUq24/xscnP3NP1T6ds8qpkHIY5LCt9wq1KVek
plP5EYGdxQziw2p5O4nchLnA0bO3OpIB5fFyK73BYBuSGLBc8Ow2BMFYl24tQWIg
LZT9CsTVkavxLdiwzTyqmVrZYYxTOi+U4IRYhG3IBuLQ8syAHFSyweM1TEptasvc
WPqy0k/shVhcceEMTwgbgZ+T5QmP6iJ8sZXzbUEqPTfBXG+E5Poepw2Z4M+daAUr
WFjF6oSYkehhXxx8xwnMniPBRGpS6JlBlKUOwi/1jbOy/tR2BMn9c3WeMRK5ZX/1
VdFG/RPLfxWuDSWYbofo+jQ/oXfjJspH27/mY8O2gMIjWu8EFJwTF93uTkZHPg25
N7/BXS8Xb8Vn8Z7NSTYF56KrpFWghEikl4B5NVykVxsI4ijreUHsQtGEn4L+bFwR
aIxRj5VaAXgjFJxD93glHHBXrIJrs75eauVhV2ODb9tRpyKTbS19LNdiletjhl58
bon4L9KNN4zwOYgb7lQIAc6xkQiPmN4zfmtl77ZuCOeRw1q4oqG3E1pstLT+L9s/
OxYM32HlQ6H0eR/LxRTMSlWnOvvyzM92FMhcPeCURIq1ls+YA3IC75Sq0rSqhse1
Vn4/exLEKAiDwRRKmClM9onfVf4F4PTg/MfDTxuD3hMfHRz07pmDXY/+9bcGuvDT
wZnKQpCQwzlfSRoAe68qkkO4o1AzdLrknW5ZlUD09RXHZ7RWpQ/fQT0Hi7sLcMuf
osks2aLtS9+1N0+7v1Bps5BxfSXaS7wglCN1rNEE/9tSMe8ITrsI8riSserMPRhV
4TDFpqsulU5QVmVVkGuX4vWdAO/fM71RS+fviQ169qjvXBAoIZcHwynHZPM199yS
puFsCm0CE099K6VLm6DevWUR6WjJ/h9J0Trg6iWnflfTE10YGG4ISRCkZHdbSk9V
XNL5SE/5ARlzgJp0bCplKhm2qRHRKQ+cKCBjxMCz0FSvwPUKQHVBmsSNq6aUijbJ
q/OV8v0FgsWcmaFnIvhdXBkw2Qf1N7gd5/rSAN16O/4fWgX3a2ZGF0pOI3AiDssY
nG3Z13zExTqzCwcHc0Kmnwarhav2lvKB/1dpnR2zZURXt4K6IpYMusbEcs2hJVWX
j7Fjom7Stkip+M1y/kvyzxoWO8hk2dSfCyGsITMS8PfrIuG9xBHX9P/a7Cc+fBy/
ejhj35thZAQqAhFC12dj2ARHUulbVHPhF0ja4Fu82xw64wMrDT7+V0uC7UNKPgjw
+19c0pGJrwUWGOBvdBU8Sgmmd0UzJuudaroLesNDFrkC7CRT/CJS+5atbqrcgglm
nqY7FN2dFUMLVsAkpgwmm6hX+ylW3OzBo7rNET7T0EshBHRBJDiaV5MbP+TlvK5N
oPgvT6Nayr4ZvIbVa2URn70m6TtM2nqOktn5t3z2GYFmbWu5mDhWAi7Es4WDjD4R
xaSpJiJTupqAe663W/3bYNTH7x2usQnlgvgve1PwTftpxb3SFGNI9jQUsRhr60l/
FUYGlqmtX/7x9ytcyueN54QXbVizmGGDu1tEFPlgX5HF2RkRhJ6SGG+lKuJR6Up4
f2uCF8vEdk02ELkbhcceDDZk80DmuU2noJDssLd1hsPwFvbzLjNDEBAPKiDDPAXZ
NLAmUNXMIgu1bGHt5KbE64p1+VrdZnqL+aYTMGrm77LvXZ0LVeNnXI+C2EkO0oRs
dCw7Guwwq9IuQiXgCYhfIm69SF0vXC5Ln5eTL1XCMBQzv6z6SSGlAUg3sdtCVvg2
L+umhGJPSuKufmGoMEy4337VL4Xpjdg8u5C2LGhDsRxGXH3fiEPs/o242HSqdpMB
4Zqvar3DJOFyKxe96O9BSlwZ4B7KLX4Igywt5zAysuBhfGg4PvVLXzNkXOUx8LoI
GAut91L0E6EHMjkJQ9AmSlCivf5m0i3yS4Btgt5vIC6lHI6Nf+h+/m5HwAfzzCrf
nqhKZWg8ukg62k1pRiTOEBC23qZojcFpNopLZ1o7MvOqcxbPQHduPHz2d0Vgq6G8
8uMy6X2u/12LX+fy9tCYkOWFvP26psXVZa+xfeQwZj3bg+I++Niql0Fz55wP4Y9c
MkE2d+JghuQ+4BR7xRq9stkZvfg7dWHVar5GaBHvOxtWJ789h7nascxCwymSb+3n
ibcHG94wU5Ag7U9JmKTz3zZLJicz9tmQe/YyJsauZBhE4lWBIs98zmA/k6GTiVnK
2aY25iUkwcZy/QqzGNDFa4oALOfpHNX8dqNzxtakB5eEjzGlDvyaj/sqSuPo7vx2
TMQV053QkgzR8nYTlY9rgUjELPPt422jgmxAox4a6m3bir3fJZHgeRBWJ3NpwtaC
1byooU2J5+N8/1MhGWWIP6emm91etnR4SdtaepRCR0xxAi1+IGrfziysqaQK1pxc
ug/0IU+QJxUT7tCKbhKXkqP2TVGTdwaoIXVIiR1PM8zQECZ8GUyMakqtQ6GA4MK7
Ho6n4y5O3N1xrgMhQLFECSB4V5sdPyl+6+HyF4e7V2JrzTXszNh4P6C+fHQIDnDm
SFxpR6uypdyFaeN4YMa1PfCUD8o3viCPIJSWLIV7pK1DY1isdFEuk4jNp4wSxtXs
fmgjOc4psy20w+M6wVwBnUIW/a0Qiewe9E560pR+bDmq4cfWop+72YXPAhPPPNtV
bEILMFcd9Sy/Q8w9F4ph9GADkfd6NBJDwSfFHP9FuBuheq5avDR/L4TcUT0Be50Y
ktPtFkyC+1Efx+evkUhPmM7Ji2JHattAFK9P4EYZ/lEou+T/UYZb5rxabotqmN4E
dDfA+Znr6okI27/jicyUl0As4v2yAZNDId/FbsOWSe/wRNjNz6f9j9DgkdPx/JGn
QlSfnpYjeVPFDMD/KFoSlEQ1jWsOisQwi1L9l/OmL5MY2LeoACD5iVzjorCc2tTF
R/vlpZ9KbPA5Zd0yMXBiGpsiGX3VnLtbMDS1C7UgfSQg2W9U//qBCdceXu2VjYI4
4rg1pMRLx3jSJxfnZpTlNtf8Df0GOm07hn7RKwQDaKPJy3pTdcWEDgHCljjqxrrV
iVL2ZxhEgdFZkNcFbGOVYwrunpN+Fa+dh7IF9mb2PYRnROjTZMCGP9/f0vbjA7/W
qn2hDPjZAzxE+GhSiYKC/nMK/S3yiwr0Cen7Enp95CQ+9NWpdsAGBw2cvNdLoZ8K
If79mRgW8ZLxDYb7DuqXBdWOPFhZbKRaKIUXYdkY0aMP5UEj6IbA/EytPO/7aC3W
f9sqjrzKY3JE6ah+lMK/KurtgybgFhI+GOf2uwJh/T8RnLEaYKQbms/AisR0GRgg
SYM845UT0qTzHO98qfrzzViSvzyEHQFpePqBym4TN4fkLfQVhcd9r/RVlNl1hBjb
Y9jCrdF2BgQC/wPOe5HOF/w3YHmb3V7NfsQl817P+wpkBHbk10hfzD0WfGhKTlM4
u6myrZc6OB/dj2e3NzhnNSWJDyuAsEKxqwn16bmhHbRFjavwxPNY5Dy8KyDXRXIy
0iNxU+xSqIUoIXjNf2NnEz8pvGXTYnNvhFqWuYRa3j3YyoG3cQTf6tQg+4q4TP7B
n7cen9zzx/pRUdyfBnT0bGs4Pye64btNy/z2H52T2hX2feOqRzd1cV2Dcos934f6
8FpjkdVT+DBZrbqGIkZeCRkUUiS4vcY9FKjjVWYG+JycNw/PG2LLbhdJf4oB8Ptk
6BBq9BtmiCjkbX9dXihXulefSs6B2Ac7InUau3iDsbDa+2aI6h8g8kvTRf3GXqRn
N/5/epb1L2m+Ck88KTU5AD3TwGlvBGqy13zARp+knqfHsdfzrwm6aREu1Ky2dx53
+5dPYNuFHjYV1VBimoDyVrKkCxelFBvf9PwAabGQpPnUppQRNje3Enr5T7N2dtly
0o/fKLFD9d9AGPOXUefsKpW24x2ldeSms++mEpN6AegP6nk0ZQNk7GFYBY2bLVeT
ejsHZPRVPWkjUWaFay3meNlOlsagWWnF+OyK45CAIWgbL0chvvTs7IYiWo8uaMYp
ixxqqoi+Rq5T+RoIS2SHhhARFn2VUWgKqauyZwvceAvk/R0LJcnuTkiC57yuEuVZ
IVZkkjsgFcjc8+ch2hHhG2GpwESxwZ29fLQVcptBwuzGn3D06Oi3oJ1QPpLVhm5q
ehoitDcQmtLCmpIwprOXgXfR95V3JiLpK1XUHK8kX36Oy1jFy8ycguQSZkxr5lKS
bHLyn7s42eYAmZOPRytlM4NGwAKswlxE+EgWECgTIuOp3O07Qrhby+vxd/x0NLJg
90Mli2K0wIJSr6cv2uxZQ/DdB7yIlYz/yy5poTdPD7Nz7sHuNZUhQhxTfaD/eL++
oWUYvNFFq/M02GgYDpqJIcINFKm9gVsD/mpp86E1PcDf5YSinaUlFFmsac7AJCzY
bzHgCI1/CPWi8odBAeyNV7/KPl00pnj1XsBo7i9fXxGtMGAXQmnvrMlRa/+Ty052
OtOcxXLyT3lRZPvMO2630QP1ltNV+jJ3kvaC3HVQZlL89b++RI4oxzdt3+1Kf0jK
p2OG1Ue8JNx2+jSpVtbQ7KToSMaIFuYmFPq+UzOB5cwBEamag2/0R5dSDkoHlClz
rcSrxNm3YvkoOmm0cBzg5qHaHOP4xbll/N95VTBKwuSvXmCAEejv0it5u2AKc3Ia
ZFxeixTTHvIBx5FWneIHuOn0lD/45UvZo2O5boKAKBt7BP8VGYvMqR+PVZSFKszu
W4bFea1UqKHEmZ3rMEqGC+2fdk9RaHmsLVP0eg+Ewoqieu3JcSKbq7kjXrj7hb22
7PSQK+CFToeYDVkLHJy41MzQJWy7ZGI7WBHB/trBxHG9urRAa5MdKT6/tmDQ6wqR
x4ebuu1ReQvunRkonEmQe0AMH4AIOroEW669TuGxBqCdKTe952DrPMgjkJW/0R7b
qg1IKcAR6WKzq1cUXtgCekLMSzA2lVPZzzYCadvPyLfmbE97tye2+UfgoR87bm6a
X0nPORf08cauI4VPI4aPUwnCF4zcLMWppoTQ9izHgn5W243b/XczlAhXn+YCUY/m
Y7MC6MKi2jRQtmXEBo1rMX9x6vxXru8qb++L7n0+qKWqQCr6ghwLXaQTKGHqlEQ/
FLL96mVq1EmQ7FO0fqsT4Wmw9sdy+8I3EobkfHPTaDbCCGLpWcBY1GyB9ohW+44o
IeDZPJe/hxGDdqrIUX1sDNIeVSeeLZGdfsu/w8z/jKFrgybml5ehtn+8vsJLwq3P
s7kRrLpiMD4LzoGsIUr2hPifEzf2Hi2DEn/QUjAc9StFbbXBG41sQzdTsvJneRUh
lub3e3g42LTyPWvxGNOWkA1iWPrI/LsKFw2P6QeyijbcrfoPh8/GAOLw2lXSUg7I
djlwPF1KFbwkFa+BqpQsWLsi5us++3HJ4/XQF+w9g5hDxgwl4O0qOBOri0L2Mgi3
QGCGOjhDnuW8lVCuXknOgiF5aZn+sN7SIXwhc29qQpDll4rJOFYXoX+2P1BqqCZ3
hF78vyprV2hhk0SNO78Pc6G8/sXdHybUrtRceo06zPyW01nPWax4iBN1QFlqp8MB
URnW4CG/7yNadoQYBtXnQ6F22tgvVzVLXiF2iRBMJkZOAB/vAWFCwzG2S7BAIsjC
Qa3cavenVeTX5tGuuA+gIrwXExf9GIsRBME8BEJLjX93nukL81ruQeY6sPbQokrg
7K2E2BSpB+6/Xs0Occv+ZcLKQVvEPKsFuDT0Wg9o/KwAt/CS6jDY4882m6AbTa3g
eYjirD7OKa7nh6EcoEdc0Uqtf/0vAIkp5GVAI90OruCFY+1m59g3Ik7PV8P0aeIA
B9YvvapYTOakJnvzciJFJzMsGIWAzxkaJiEXUSCmJIl6lr0406h6fgONcpNRb3OP
dCPi1mdmBiQWfllvKu81qPWT4HxNEGuKUCti05Y7uNgqiSipA1RHSWCL+L6ZBY8Q
SisyrzLKBDDaRuz8n21NsFW7FxNdclKLDUzl0vdNjqy3DbbYUGPzHR3fNcxKrGWl
ySPLxu1AL0Yxasi9B/8HYW7YUn+46gXwtphxJx8NYKiaWIKWVr4mXx6pOyR0VE2s
oz0YpD8SIsqBeH80hFLtGzr1SRckxlAG7AmJz+sBe1/WazODn7Kaf3HXYL+TilpA
vDc/bpV8HxmfaBZSdF4f9NNDYVMKxS4ihVDc9Jg9J2bwxnMpFO7hPYmdIYR8zLdr
YmXfshtIv0Jw6SaEtkfaR74i6sRVAm318t13uTQYe8lQxlz5dQODP0WiRn87EhUv
p1MmBaJkTiIbcVMYJdIqjvuNWGjcfBHgLm8IPwJOjGLoHKH5W+ZjC0+Hdsw9O/S2
Iwu+qXLq825hi6djMVcq5VX/Q9r9zgPEKai4Bh00rjlKPu2xXwo2zswnF92gDozB
ktxGwNem8RMfoJPYcOe0cidY/enm3loW7XyQNth4UcMXXrtFeq2+wmU1qDhPyzLD
8ymRnGed4YdR8/FfzAwpXvQMCLsuK9NbYEhhOvdyeGBmdzu2CMOdORt5M/M1uV58
j7SxbB7dW1RmfAVybZpE8Q+ho0w+mIQKV1o4OMWJTyvfPKfC9wGy3xgcn5AUkLpO
V22SgMSXD9U8QqpjfzmdTrV+vfhPTklqjLuwzXmmOjh4sBOsR0hQZUI4Kej2oT9y
pEGckTua+fXVq/MMH7iHXMS5FP3cgTb/Kf5oRP2xAfBK1+5BOktceZimI2z5EWsn
OWIoyYroYiSa7TgvpM1ACKDsuHtEXq98VX1MIVYRbv2GHM+IXgQS8V1gd4KUHZ4m
+qhjtMYsF5MDYpMdJXHHJS4hkYtC8Oites2w/tZDLdzsinVPP9apMeIJvV5BwRPy
MR1irR7alJ/l7ZVce8H3735atZRLZ9xlTqCMGSjDfV4V6QyqRL+P8y4g3KNaMTVF
w6rkSqIM9aBhLw+x7nfmXyyFzFYbZt3xp0HkwC+M9eFz/eSiabNzJ3y/DLcoNOiW
CJXbh6+Jo1mKpfnzT9mv+XEKudbqkRUwhD9oQRT52qqgXROQRSErBYiIbhKJVV1J
xnnIXPmFJvLM/jQM2tfUY/C6bSvhIztYqFBab02xtwmtbi7Z8OMWOH5fpJfiKBgb
gVZ7TWWsh/Su4c7J3xenttUJSlmmQOj81U+7Prm1rKEoHfs4HWQHce65id4ZkecX
cOKdrDEY3MrJSNSn4kbaBy95Cz4vbMIPRyo2hbSWIcggL8ELlLAUG7tSuXKxHGPO
nAkJF2Bd+bJqVKAj0SqVxPlYRKkQl7aSGr2XTVe96l2aM/EfOg6ztNUnXtjn0nVB
mNRVghOepaKZENwTD9ryy1aavVDd1utkXNkv9Tlzw2LtTvG2U6xT6F8pbGDUAPa9
a3e5OfAolRQMnab0kh8XOBwljNIMSzMZvZTbWbiyOq3oljmDQus+YePK2O98GRE+
v/VSVPa6/pY1eojDLJGO7Ob6k9NjfZX4OHxbWmS5C+mFR5cEjVW6SOa7c57NsQbX
OcJxKz2GSuxL+3Mkn/f9FiC0tNrn4Hj9SvDqvjyC77KXO6bb47kHLjuTTflu/P4p
IUABzftC61AUUfxFn7ndh6e/mSucwe5r1CmSQRJP5mEphBvmjsR5MsFyY7SM2Mka
K6uC9B5DaEyFRFjO1G12sufjaFMRtNhwSjrBrnwZfUYljHlI1wtf36uZ2J7p3/Z5
qLsnRzuirkXYslj+PbsEXpIF+2gtY4k2IMa7uZzFxPt0pdTAmoo2JUI0gj9rvflr
7C0KuDyLJgDYzw+xVoNyzLVuPEWUaZjjTMKJEYDT5oHZav4RwhOYs8i+dScZ7uQm
rZatB3sTJJxyMnFwRRgcc5oZNxUr29ZMyXeouFpCuEGfLWJ4mb2FpMrzdh9XdpIB
d29u0fkPBN6cG5vikzoKjg==
`pragma protect end_protected
