// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:26 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
EHrGl37MA6k98pvnZ8cFuNikASZm8kQCdXXZSXztO/aZj3cGRT0a+Ff0zBVG63Py
e0hayNy4FVigkP3+pQKFSZR0bywA5qxmfm4Gj7vGmCyZV57FGqP4cDEOZdMN1w9D
J9IqCRujSm9tVqsygMleLjKl9Ek7ysoIO1YmBuDxkZs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 762704)
Qj3vL1eRKQaiQioHFcS5bF+KSp49NRua3pXVZX57UDSaKwDWWdolt89Nw77PAWMK
Ij4O8hP1bIbdT0LRZAnzgYHNgXofNntZ/krgdz3DMPGcskEVjFzkB5DZvtIsjycj
F65Fn4RlHK+iK2PdeQwWk1XBQ6k1N+qo4ejy8aUexs68sa2mnzVqjQ2d3mHEmNlU
5Q8UWikUK2vseTLJ2wwDgSFROVWWrggXJlXfR7xbwrYsrBrUHTNHB2iUOeDLLWeL
IaaXPkat+KlD2aFzuSicDYxnrOiwm7rWb6uv8+NZZSx6Dn1K0uL6ngJGVf8HRAun
IXdhLwBO7jzFH3LUpidY4H1HGKZH518Md7C/C1Oyc+1A9QKR1UTM0ooARHXkZiUD
m5vH49PZJ1FtvQ6VkF3gFMWsOnjHAA9TrLxaJ7AiEXL4DbBY2V+s79n2gW1Seywb
q2VJbwoXJdGQb3wg5NPjvkeUcjueWgTncwIf9tXKZgPMcP+JBx9Yh1+2HcnBdB9D
38lHAEgZwWeMuB/Om1lXSJWCl39ErhBQQOjfw0CuICKMW18n8knC+QVk+/RJM9kF
XaXuRumSSQQ1LkXBOkj7O3LbbnFhfQCAUKQn81qGwR9O1lIn+Hi2M0Z2qhm2iEFi
R/SgxeZEJNC8FF7tsd3mhyk5fctKJIUVrSIjQT40krY6y1SSTIYLUKhT1AmQFh3s
1F90w0BJqpgewpQ9TQafoALrT8DVdhNzVI+N5JfFT2XR4Va6iSj+m9RnOzjgzpVL
K3ZJ7/hSnXyGQ/ZUdSc7WxgG1WDOWQoD+7Gal13ycZPkOc7FZt0nnAAb+Bw4r2I8
56FhO67QAENP3zdTgunjRYUffumW9STEVRYijRqMJQK9Q+uOgSDL9i+9orxOzLA+
Pd9DOXS/IunIGr9PVtNp12YtPP9Bof2xcxx/XkjFLXaI8u86Fcvd5N114EzG1WlR
izeC+0U2STsnPcb+FLusxsv8+iD9ODRVFrNs7jS/Vi6/SGyZeL/m4pMOHPa8UOkA
7cqNte+eVffBxcvQtWlDWxfbh5l8QuIQTXhr/GbVpNykOU+fU89VYY5DLK43zqpm
4DDbPowhhVMntZXqhMtWVzvOylH4oB0yqwTDbDehPHZUgaM6glNkP5TwO9ZIowIQ
75LrBPTfqfDjpQwII/Q+BXzEjKYa+axhFCF7E6lV9vkKnHXyxXEr/bETsm/E55Aq
f06dyxJNEKsrO//eot4Q06gaLR+Akg86kBYVOEaXwG86/eFxMPDhql6yEErTfabv
ymvVh5YjxEUXS/UA75JBnHRXljtqSpMhsmhR9c2jQJWdKaE8qf71gQ8djCY0u8R1
h2m2ny0ESWwENOPGaWoGn7sjiTbmMB+UBywwzEdyGWIMZQshovLUabyAeciJ+on6
2ZGYAWoem1CehfCYOkP4xoXkthwidy0zLst/Vb7k6/BPLwBp8YYf3050iblxsma8
ctlieS6Vr74ZH0QfYEvH5kSNxbuA7b+q+264dvrEhsB827RJVDVkkmTkFDScQfAU
HW+qhUq2TboBHEalsQ428abQBWlJWYV3htmUiTha16BnV/b7tzil9kUyWNCe/UrL
ZZ6irX4ndOIzpaAq3wSFBD48o7l/pLDhbJWTMJNsEL/Yia5pJUUONTAGPWpmLp7C
IqsTOBVRVgQx5ri4J6sfcITTGKiiuzOxCj4nWZ/74ARHghczxXEWQ6CFOaMvdjx4
U8CbqSnN93py6fnFCCQW37rz5ndCZMk1p5U2wV3E1CW0eWqZVA+LLuN8jZ3K1pSK
uknq2J0JWG8OgaGrrui3iS5peDohZMKlE55l143ReB5eM05batp1t2ZYCQIQFNxi
bd0q6hEdbBnzxbPjSbcBs262ST9PqfAoYg/3LjI5QJUJ3bu9vh1NuqkPgW+PEPum
8neyhAk3tPWNY25iwacVh7KUQPXoy/Vd9EznkZNOSyeoKe8B6IHjSEhyEHOmxlfG
NHmkrOJLE1GyIOC9BfVoOljtsByZCuYa+PyR1rGaYxgWwJ1GxZCrCeJn0SuHzCxS
28/IW0dlHvF2lb9rW8qZ7DXr4lPdWCt5IYDILrNTmTvrRNiPHFbKR1HK8suBdUrC
vyobmNipto7A6b3F7nUDn2BAhM3jkN8V6gGbyBV4+HnQH+8oaMIBfyvxxBI23Zc7
luVLlKzS0uABQe1y98u9PE2LiC4MtnrgxDgjzTQAn65g5asbCmFWs2dBhyFXoYZA
6bvwVq7opXwNwiVbK85ZLhJVXHAQFjLqu+K1/DrdeKQDjGHgADwR2W7ui32398yc
0lCHrmEX/0E/FzV9pr8228OQAA8PX/Ji//rxvXtRsdYKVYhYbMtIoqTYxi9AryuN
1oJ9tlVUQgtFqX/eHtsMX2h7D8asx5QifPHoE6slsXMvRziLXPGnx+V6aZX805h/
cqJ2MzKYLMjScxaBegsMJ5hMpt9rzVjqim5PgiXiEb4arlbq45Kw9V4AVrwlQWh8
7W9dMEVoTv+Wa0ELVvbEAqFlI5FPApO+gxXNtuEDmd/42uv17G1J90HNcVykWi6/
bw7sbnTdwnw9fvOLoBVEqIoZAP0EH35rWvGsRdjvEk7Sc7eVNy5MGXjCISNE/iNp
NvHGZ3oC7MWb8JSs3VW+4//d7MOvBfmuhmXMrD0MGBvSAauBcRQFbomUpra06UgK
hyF15mHpIS+bxyOgulO/2ida0C6O0/AMoBsdVePmkGXWvZYOWDT7vUVV/QN7yphT
E4wtxo7v/1R/3P/BkUDTdScbk3XPP7vvNvkOmFmd8wtkuA7atuAtyibLt6djfLrK
jPBsEWFj3FUiZWej6K/6x+gJk7SooGHPbtcbEEKPF5CqKmGO8R3rwFFgBHqBbwDd
kLtk7J0myKuoclA8VsWhOFw++7i2grIkMMayBJbF/7v26WlYY6rnVZkcLqy9TUXs
XxktEJhhlIDvjbFn0yvlYMJAntR4m2EJ2I/nmOV2juwIFjT+pGN+7VP7F6arTybU
5lCAJ4NQZNYzSFE7S8MnR+8NUNb2AoepSZTkiS+xlQ6yntpamP7GiNDYGXjy0nFO
fwUOxOySLnZZ1EICaUHLrZY36sj0K2DGpwpBbAmDqXds2Lan/YeJc7pUW0mr8BGD
GoRRAxuVDyZXW5/07Fpvb21D7anW0reLrifwtvA+kKVJCvqXNRQroCsvmylUthfT
Pmcbi86Qvl1XdQWH1AKWjfK88g92haclieck7CZqWRjJkIS/poqxohfcswJMN2xl
qrA9bWVNe3Qc4DOx9B36FFqNSqUXe5tZhOGltlf7jzZsjRVg3+QE59u5mQ1uVFT5
0z9ccQMyOqf4QZnGegSUUavEUHnY4xmlSjoou8ms4GZ7v2+tvTFRPZFkgjwgLaI0
fz2OyPbb0Z1dF7zvi4r5iLQIkX3qnfS57SUZ1BBr/gdZnwdqvAKCUs7mQ7ZkVFni
C0fXug+xyQDxJFqUUEuDiNZbWd+P/mcWDHLpt+xBgPILGi/nHSqXBgK43W9G8OjE
7Z17zwr86YMLz1+qS35FUKexZYZYqBNgSWZUQNYmRp9J6uHKA9Zw84NbqBuT5N+S
AxRjyYIDqTfzu32UZ6vd+lfH//2scnMrBjoHscs7D90zIrcA1vFscHsoAGGl9V1U
ffOHTRzrHGUSwWa/neTGe/ZsUzOsCnh79kP315WhwzwRrRhMLr1Oh+xH877mX5Gk
dNQfhT3sXL/fNHjz8CYGGMBOcf7azg5B8g6uo1GC2/RjniYYGkS5BpaekqZTBoB6
ZgGScU7I/Zwi65VnpZE/WXzk6GNU8lLOJXyjn4f4x4BAqaZ7lvVOqVJI+P8asgYw
NHXhIr9f3neeUtHOecxSYxmE9GEXfeuPAw7bAkI1t5mcmi2vXcGuOdNquanCu1vc
ZMuaumMowyRFddOE6jW3zx+U3PIL9l7+HWgoXUUGUu5o15ztyaDivcIJ5GMxtW4L
s/cw1CzM+FTHYXKiAvmLPcd/D9Ml/uZtKalTx/jBhPK6hmOju6RTxpnZElpkoGor
fROaO5rAD2K2p7s1ZtOOvkaAGPskgdFH65bQhskUdRKiScw6dWyQMe0JFcaVdsfm
2Lp79pEFvPsi8NqlgPKqdHPhkY7kaJ+6iK4SLv9tpNTo5bKQij9JuwCebstPlLT1
INsRkDPRy9yErymz/JLeu5VGMoJb/5yFMCoQwzMR1Hby16Ci2miikTEk6RMxO39J
pjXGOCt1HQ8/ekygTtujKt5R83ZDeGD53zyDbfu+Je8L1egi4R12UPmKhiodHlor
5WIroBJE3OpkGKfObVf3w2kUCz9Pbp7Srs3plt6GdxEH0dUOu/VDKhb8zjtYK+f3
n24L8I20kaGo43N0y5lVxmDBXKE0LAT9R4x6pttVfFEZGUvMzsbGXfD0vIAb8y5O
qhHWVsgITx5My2DOrPPu7L/jPTgbqyL3HRl6QYyW5yoBYghAXsTZhw8NoeeI+JHQ
aftKi0TXC+q4frr7rTzvt1Ze9kEIHNBSwig07ZmryIKL4ufY7H83VujKq7VJqC/J
GhMGYGjRcCPp6fgnqFnI3y3fzDdy7a64OJPNF1rmi8nGjGviMVXMBjkYdmtwQE/o
l/fJHAXk0mZ16hWIkBz/zaQgr2FJh3r84yiJzcwIbyZa0XyK+TdBi91fArL1GLaC
h/wmnKZmHcK9KS9CD7qwOgOUrzaMFcjXzZOX590KbPEQX2omQD11P6QZz2KLw44G
pzwSbWLKdYwOnqBxnmM5WD+vkeja8VAQdGPF4GWnupE5KpgUXGGOUsvmBP8WeGDU
q5EAthHDklSDLon3RnEC/Ql/mTOpBCdMTNOKs+89QDlLra30T3e2TbknyDXFRSIU
7t8gfdj/Spcmh3J8B6D8HmuQ8tXra61fKl2/REtsJzJgx3qWdbrMTG45tc7RIu/G
2j8wroBz+lhmcFRaIja6zygI4YZjQzjl9IqzEXX3Lhzwgo+oWnCz77usxdZbfLy5
RSL6FXb+bOAIhn2EJgL2VDlw1PGt/m6nlXKVFLkunMmlYOB9vWQS8Fyqv5a9lrXl
lxQThziKfnsQ3t/PDbFKfVsnoKIkQ1sgtlIifPx/oJA65OURulTFvS13SmbLnQqd
SMUVxYeu7RAHGTKO8DGPiNPZpuNNKWeFyhBYgz9U1XszyBy9OhdlptFukXRST8RO
hUqQzbtnqq4zvrm5DtFUyi3HOSsh+izm0ybAVdXRxSlpe2Xu2W0hA1tbqgJGGm0w
A+A4QUhw4CmsGgNzv5+f85IU0nMxbEz3iyMXN0W2euJH4xtIgXrrTXpEpK4vieNf
b467XeCKGjAwMixjNOR2/Q3rdObO1WcvMA4MYxCGne11EZnF8uvUOpy9EmravMng
pjTVgl8dP4YywOXcNaGM8TB/enhrroHqFzxbHqAtqiElqZdtrj/JyZNsTDUryttB
u+PIHlsbiF8B7LwFi9YoYYSspaSuZHeqChvYM7jv7gcleSomFiOoxe9Z5pgriCji
3k8JbLwWvtIRt5G/GGZo2Ra7oVM9gAoLVBdHmM6QhN354RwFo/8PtQIrkjkhyPuv
8Dvk+0HpiUHgj3fwY+UotwnfBvMkBnAChHUqKdOAsQLBbdYcqhfVE46t90tjkmSW
hcB3ZLOH6EPTB8XOUNa/WKEwJY1HJsaDVpUs5kg29NYKbFlZLcbhLDZ2DDOE5o6q
jNhzXA7DM/PnuDaX6dSClKdMuFzmevDQsK2YkohPOePJNiQuMQzKLI0xm0TxxWcE
k+2eC5K41OBhPDpFIdgNwHE6Zyr4TVI6XrZFJISaAO3O7/0ryc4J0ksd7gNu5zXm
ffBuSddm2UlEQY/Aq8NzVg4f9fmOEOg3Nf8eu6k+xNiZcRQVLacQlT/dvETjlADd
rT4yXz+QZn87DDG/uJTev1QfcEokRcAw+jhKuyVoieGibbe+JUuh1Nmi7w0vWGip
cZvWYEUDvOWI831GPLseEU7ZEI2aYs16Nea8x6JcaFpMbspofGQnaxoNCTn4vmbx
rPUKDWtYGZ19KDxu1jHfiZGK9xWX29lTVbWlVtO7JO7JxdDIS4RcJFI7o8PCSdXH
4gqPmz/6EBELnYKc1n5ptDCQ3xNZdbBAi2pOLArtfQ4a732iNKGAplkcNXBp5wG8
oloYm4/48uciAhaGyR7eJUYVhEwJuZHM16iuXH9lO/Ueii3XFE+TNyH+qtSXlOcK
T54XzoVXcdPiyT3m8vz2KwkLk2ADCq7S5nGqB7Hv71MbQhAY7XtZfLJ4963tKgaD
8g0BtWL0XeKJMM9VbO/6hTvnEqsDWoDy9hYlU+lL/OwsujLGxy0w+YrJGy4L3g6R
XhXrNMg8gtb9mU7y8fe4AyT+rKdWZGb3NehYvzCpgyqAusqJbBTsELmXdTkNmWkq
PeTag+qSOlypawalC6KPDctuC5o8AxdGsh0aZab4h817XUctdloFkTGTG97ihN8X
5+zu/6T/oNvCwyyk6xWRkqVhguj4IdjWdELMb+oKfK59VZdQ/klSHbc2HLqeSwVT
bjHGqdSujNUg1oAP4pUiKtD88PGe5ApN+WEtbDYiI4VVNxKrdlJmsVZdK5FrVWYg
g14IaOJVAFu0in+3pDXhdNSKZJ+qEcYXdmpI8HzHFC04vMVkYw/PmgS40rSrmNkO
FWVuUmb/koFCgXUlJDMyribWeZlcZ62LaorW+hOEA+vxFdVVWXqLbYbT1pg4qrUr
3Du18RAqHeUcFRyp0sDOq7GeITVDnwU3IZ5tggHQH0afiRCsoNyL2lRdq7DIHZwc
2rDNMftTNgDolCcVr9ebuAzYpHi0+Lhhtn6QICB31wiNaL3ULlmSBznYA5E1Xfl5
LZjPqyB88CtxYdp087I92kEfCG7+p6TvE22bmoVzABu8enaWT1IR0dU7c8mrrTfO
ZfkQA2/og4ON9kZMyE9gBHaRmW5fhO3Ht+nXd8u2/8UsonqPFwqyyZdL9KBY7Y17
aSzB0yik/j42DYlnD5QzDAypFF3dHdMBhlz9Hz0HfrMd6Ji4cHhZKh6xJpZbfCzM
uURQ78ZF/1/uI4yu6QBmqD/htszNl/7piCB/Hi3uqhRoza9RD7mY/sgi6Hmp6sC2
HZ31SWoG9/KbK2Q4bUaIoh+iZkwXD1aIF9g4/HQWFx6hbGHnBNhuadHv/XPlYKMp
xuNBG6KuD2IMPo39GhntxRm+6fUojVadsvObEnpNBlIB64EWdvVWg1Lh8dz4B+WR
OWcd0NdgawSDKC5Sf9lbzVPEH2M0EnOhNeq2I/bbrW3IhB7tMlR0BQexgdxVTDAN
cZpDFqBNNQOdz6nAvYmmgDFG7c5WB8y8xqelXay9uddnbUvs0TvW2IrsCbvM7ZXA
oS94UuMaSUL6y/R8U9dM0qK5UJCpYind1dPz3o/WEfWcqQWHhWXDAp0MUyATgSv2
kp3vDqCjbwxrH8IQgdip7c5JW15sgi4MYmBMUnCJcb7L+AGzYsAnaE4BkuPHEcdw
EeCGhVSQgN69t3Kvi7EWx50/W8XO7sjMR1uNbdErP76KXGyTDyjn13RD1fzUM1NV
EGYpcon2YjaBxIfQxmVz/Z5dcDhkXHFiYEujd3l32aaVp5tMTBn5jg0HQCfOlFvl
SO27UhAdVGftmcmbqcrL2U8CW0ADUbjMKIMwSzyR1mYlycSRXHZgTColXtrognGg
syEq8A6BAMoPnwmJfCW5pT2Mx4J+BGHOUtZuf355+zrQFr0uZCyztuN48eNsOt3h
JuVBRYday0yFMWMDgTBOH9WDO0xM6p2uCpRq3uxsUtojqeNrATXfXAlc9f7uWPSR
zqCgtHCGocGZ2Vns0HP+2kBgG8IAgXSt61O92ePPGoRCBwMaYJ7XGgFcCvCh1A25
xRHTeQUilMDjrlCaO5/w3nkXSLxzdruv8EA9YG4pR7wJ300o17sMfvjudLN+LOpJ
o+twjIMDTwoz/W79035TawW2vhhywy1tB7o+Kmj5C0SlwEHCLbjOrwUfj+E06Nzr
DYzJ2dQI2P8uRZstelpscJScWCeaBrBsKqhhpfDbQTZYEFozT/is0GY+Y9zCn0Dk
3d5mt/8qdtdvPqaBe1++iPpfB2iJTo4kxxpDxK68lrYT+DpMY0f6TF1R1dPqcD04
oDV3MzXmsn47xDAl/suAqYL/efG6e8NWe1agqI7B5YEKofHnonuHn/7//3QcZm/N
SJQ456xb2dpz5F2AsVT+PqIz2opRMcmhs2fSwnQJcFystDC8IhngzKlAyIzGxFpV
T7/6dAOSeILaXoMdbp5bM7H972Sv68sNEawnOWs3FI+dZ6A+dZvMmptbVcOjy216
kXdWj7W5S4iWEh/z5Su4y+p1sz5skYMOX1NUiJMMNlVSAsm3I6TCEEMmvaLWUODq
zHnPe+0kcKUqDY3seZulKeD3r21NsRCZnP91XVSxi3ZxJfn3wxKf1V9a+EGnkEnC
ciDZdsaVS3VgIgaQhvwgjI0WVFB7Yzy/stzEtTkxCbjzATsTm8JpgK7RDSXTKHjD
sCfe1nxd125AsTWa7+DzTnad4V60ckcmF+fBI7HGZJ7OvtMF1DHhuV50gulCwT54
Adoiu0aYGqgLhtUxQ8nj5v4zEPnYVvlLChajKoPNbYVOfLQ7+4kVpYVDDchnczQ6
M+H647JJNNJYD7DYqjEoCgnsNDkyB9anEDMrV3+AQzU5atQPsDFubUowWk4n4wdm
MhRr7K1pcAoU8OU2PSC25U3IMNu+Q5MBTw7BgWNIbBuIFjMsOQqag9pJdEjIkRkp
KKxReAwxQHbJJ2b8lqgOKJr5TwfY/mQj99B6itjhGbt+LMB4HPWe4u22YbtmOF/t
Aot1XmUz8tJYBaJA5mBNE6+ysngNXWH34IHVtYRZuNpjFRpcYmkwUvz+29g1bB7p
H6j5yoWHAUgbL39v80Scs9X/R9PicPH/WCd1cQrcJwbNZGFhuPf5F4vllxy/YdxC
OGXut6P857NU5N7hHSmzr98lsRoWHeCKqhnaUZQsshAdT32cRNzOs18rnjvtpyv0
eqeFrt7dbJluzXWRetbsgdPKAPZia810+rzfjzrAsBWwJqU1GT1JxlXt2p1EYQMM
2ILo/0kJ5M7fOif853hfxCVroF1ZNjJQaNQ/EWqalRejqakFBLpk5ObS2ADhpEi9
Do7jpaHatgj1FwoJKxfm+4+P+b20CvC2a4A3ozesxkB0RvOC83GitKYtn6jOc6gh
tK0M0CvdHYf24kr1fzozuLQCtQLxpyUP9nQ/o26Xedu2hGamTqLPAGZWkBCpAWmu
8Lg26bYJXjUbG1q+xA1+PAoklLCreGSo5E95yQx93FHvtfHcOVBP4rt/jcsNWU8E
wVs1mLQKJ9hIJjmLk9I2gSVaP+kN8tLIvDX42wsdZTdvyy6TFs4y/osqhvLivHDy
rYhX4lcXyGEcxujt83tGwysR2iqOC+1N8H2E+eP5CFJZ2fGCVf2QqonKdpcZ1mVv
NmyudYfqk6VRzOZNHVhTevl3fgE0AKuOJ/wMUUT/ljyf+jMXq0kyCQr8yHGBUwYm
8ctsN48Wt1mqhpZvUSdovmx0/sICPgXb13iz5bQAhp+C1UgGHAzS95ZZsyWk9jGv
jn9OpdON8LzwIgEsaQvAK/euRHOg4LVfbv9sNS0vbmEIh3cx5Myzm2IJdwJsajBo
o9XtMUL2izyAe6Hqn0ZP5CFjD0i08ceeFJkFpKd9dskKlmnee4p3SY8VeTrjeHBA
mZH7AYuiOap0hy9t+iWTUanUkScxq5zj0KJmU0Rr80DhbdWdhOmXgoz0P1FL0m0g
wMaJl/KeIOZaD/VG2CZo8MLhnQcQ+I2cgMGwIedL/h5dpKs8YWlB/99wFG7cr1A8
qr16/BVvCGhmuVATkU8qaUBhq7K7u2XHr45XRXw5EzumqNmtF51d/B5wa2Wvb5Ti
70u91YPts3P2xxRCwGxebetKfKzwUx/A5N+rRZ2fl+WeydLMmTXfgSE9hLA7nbo8
XJn8UaQkhkjzGapFHH/wPB9zvBw8jWbaZp0lsc/aJVUhzbu0x6j0cIJw9ynmAFzH
rkXj6AzES0Tom98SaRQgarhnVBZ2hlNWBhI15Rkq14Y62suJgNn7c6fKzwUTbYfe
NJmKmnZqapV6k3QXLksIHx1RtpMZLBRPsrCbdEyDlFbm0L5YS+ynGHEQmFMItp/A
gqNGXrzceRDL/g1lWcqVgHChZibvGr1kLvMsI/hKGyCQ1KzZEIdavSOOVhzXfccP
2Ks54QbPtf7DIme6kOmiz0/cmjmLE7hJ5rmRK7zE4X2Zw41ri/ojU7BDvaSr9Drx
cljHpTB9Ft8mte9nNWGwHAbOt+swj0d0UV46EEJdPuDAexrl/KSvueiqxBX0Q06g
iwiQnwK/X6MM9wCjHl3TkOWv0wSj0MejTvr8YtHtGUNXyWqDix5dwql7MnGSMeoi
m5G1ccw5fzXupl3kRRIDfoVoqngCwjE+Xh8MfJGmr1JpkmUDl8pakPTAv2km53pC
gnpldfj+pFgnT50YxDrpN7oRDEQsrLs1BPQ8FmZQT3JfOEkwWoxThUAYlUvcvUB/
7o1P2QbywXI3/hxCYlmQylucaHYMutImB5IbMmY2QIvvFEKEVZ2m+MgmcnOXX4c2
1v1ABNbDmnenb5tIxNLYTY2DrWgXr7SalnfnS2XCLEwbB8O4m9aZQ1mdpEgilhn8
mpKvDnJWAAulg6R5CNUi1eP/Qas2lBZcU0hBH09JyQenwm1de2SgE3HctVGiYFFr
ttbIieyMRaUhJSVO2ICvnd5EI33GCp30m5G6xlxfFsFXOcqe9jkGFGEgrjKXQ34h
jOODzS9PQfk2/UPV/6n6Vt7/nA72yP9kSUcug8D9d29WvcK7j+hHd8g2VRfckqLU
xCiv8aBLx4qwWdAuGrtHBmi4YzWVGW+nn+dKMYsPoab9+eZLq27RKeGyncLYgdFp
9HCQhURuzOoLdlEOE4FSclYsYky6tCXDYp5ndz2Vy0gTI9YthjYV5TP0mhq9lbvp
5p5uyJ2TqMB8H84RdXDYvYBAQ64TJCVnjftSAK6mUlxMN2eqaUNaZKjvQhnBc/m+
9TInCxGsU8a5hYQWM9JC6PBiB0Axog+kls1VcCWmi7TTpS8D64/zUX/fXHg+O+0o
55vu3G2ojXx8rfumyL79mAlbegZZ04uG0/fEjf9HUXrwctToArfxy9YNfSD7B+gz
azSvySonaoQamsMdxJLql1h/O+jThyVeU/vdd2TTQP8LW9aM9MtG632hS5tjE5HN
fpZckOhh941gC84lk3DFHT0/yA6pMpJ3bcFWgTvytfhU4l+DyDgFILV/gqfKjJ5V
5GwOL4lo65zojKG9uNrkAQkdpjjqhytmFbCQZNJc2eIf87mxlElGOT27DOPlwXaE
NpvOK1gtTLHNPhKZo+Ix6k7twvZ6ODi4g+nxKtfHjxS3BDA/lFBLqibLONJWmWai
4lQAYGxJaEycLUP5FqC2KeP+kplZ7/WnYWS91NmHNFCRxcrGuKy18EXyrL7Hh3Nv
6knrJWXiJqXOYuqTmpxdArnFflykeXf11ra69f07hW2lhEtmlBdhKAk8DR2hAwFL
zL67H3NABaUGUkgS8rrX2UE9kyAp0hSiKiSJ8nDwnyIvxCni1dRsjOm9z0Hl/Pu4
B0+FqVaVmVv7jYwE5MPWUaliI09sC9qiOnrJIBNf2tEZ+gnr9u5+82B8zsm80U8Z
ZXDcHwjO0QNElJr+qYkQDhGAOOSvSRSExo9Zpy1yZqOMpJDTBjcH6N+ms3Yh7OAH
1xuUucGJpz6wbpdN73oMuht6/UeI4XbvrWF9R9x079K0+G04VRfBd2MTZJrpG719
hctR3w8LqJPmt6xDdOmZBX/TqQHRG31cdEVNHgxVn11zz2epgJXKxaat77LL3wyS
ix4VWSDcz/nV0R2vsuvoXbF3IGb9dgNkEY3rMKC5tYmJ3Vkiy7b8PB73d7k898Qj
AgZfI/KPhi7ynLTP1Ewk4LIA7Xq0P+2Cql53WjyO9yOxppXiM8bxaynnV0Lj1+Cg
YgIN7SmALA+5gT/N391D7eJYEd1InzfHux3wUQ7M6SP6F8VlHAL97zWbVzVZxQLP
CzCBsgLBSZcgz0zpqGPhmTzVEqBRpzSxoot2cy3EFvKn1cQ/NeJooUdAXorx4Y79
kufUAJbNmZTe2Nitvf38JHCBzIG7NoRHHtYGWuQ8qiNZRB9DjWd3VQXCBt42201Y
/fjymjTRQaz8H1IZ1hiQ5Yn6z9EN4J2jgngUUEAbQr9aSVjoDHohr1ezSwVQ3vUK
dz3KTd/vz4v2O5N6QA3Ny5BExbbqOwrpLCEQwlujaDsGKwxd/WBZRWpgolZ4Q74o
3qAzR70arQPW6Wfj8MQuOVeClV2/F0Nsox9fdAFNkpHS17IBgyaoe9uY+J8qlOff
Smu9YHM55pS84/YnREdt1cL8HHV4rRgYXnQEGny274Y6QUoWgEAOIC36IUEzLDyb
xulUQqhjBRi7YY2xf2b6GZJdmnwG4GiKdAJjlVc24eXjz32VqTnMS9vbxhd4hF+o
MDoPMIDslKZKrFhuGo3Bp7R/cCS1XeL7uvBHx8SUOsnRCrcak/avd7Rm5Fmy1tdQ
X9BGK+UTizCmK1yQmPQdOpgomcff4vAJYr5W3wLUlfjmPLRWnQvazGQqqgyjcdBq
jGLEMlZ+4VglKrgMpSZ+IOzLSlz/IuDZSyUV6XNtmkiRMdn0wD0vFjb8WQiRNUCT
7pvENpR84vCoBZOaizIiBpEgB7cr6mEjF/Sgau1X+6vRSEDsRhaWuKFoUYMptnoK
4GhXUXOhlGf0RdSjcxTDa9ZS8K6B8IWE85teUNcsi7AiJ5MBGfwmijyuEzfiYKk5
K7BpK72etkuU1O2oRR0HdtvgVbHSSDO0Q4BYgEeLK/QYwK7+g1yjfoW//gUEYdVt
Ty/Z+NT5t6srnNGgDnZNS6cXWKa7eYxtEETtE0umvcUhZs0XizjVIk3Pioz74L3d
jK4UObV2kdFJHrYUQI6HkXl73AI0xYMyR04LiBRODbTOVs0JMVCKxXdi4GtOFMGI
XZvZlLLGfRkHC9HzFCKjAm9bUEr+3QiXtWkxVv5oLbLeQjcHstb0lSL9Dw67nGuR
Mn4apYCQk8bn5RL3oFuWZvgsed692My/L+ObfhGqTLXVS2fW4QRibBYM2qEDpR4h
6UYZbh8t7yuKWfVXMr4/e2nfdR03rkZOq3Fr5uiPiQ1eC4vThQVuMORo01q5EG8S
k9Ehys+r7OdhBfFuymgFoK6zV0bC9VQaWH1hjOHLxSRt8k9KXZdKQmEfUrxftHgW
wzLuGdV8awPqAphzdAMTmmmpCrqFOgM2O+KXHkXpt+enWJNnnL8x4s5Q7+oSK8XS
uhWlhNNuR3sP0mCwMFoMr90LNswhK151n6aN3YRd2aNzOPXhthlUDh1tWpSa+NW8
m9qr7ucpEyr7tndVGH+bZK9kSQujnwUPYdd705e7FvdPweKr7y8OSEUCnT1NgiwC
oQGmF/1ZiKRqCXkx9OWOHN2O4MEbnVYnRP/r0rCvM7FR5jpesxyN/+fkMV8ud6G+
RCzrO5VI9R8pAtKEIYwg2VnlxWyqiHhlRPV2/PrCsW290bF8EnzX48WekvZFChs9
qDGUJvVk2sOBQfdYJ1oHpDDgb8VBmy5NWbHsnlO3mbtpAXz8jW6uKut1PuAaUfjc
08aA1STSoxs9P6alfeL3ThqxgAn+HmZnO8uspkCchDmQF0hBZzTFDGdKkMFEQ4hS
UfmkrKgXwGaMxOHD1CEiRxtUvI6jnRs0K/oeQa3wGB38pd7DjJlckPJlpZduGGcA
Dvmop421bof4eUzO+32iAxYcWWFuG0IRG6cANC1XgJl0o3algrYxV8ArzedkBqbq
R1SmcQY55NHDWN/6p9hrjUEOTwDejN3hJW2sFxhdnUhl29kVGioByu8fCXD2tuqM
jFyVvs3O/xsxB6d1Fxe027jye32LrbeADfK/zEbBfgpri77Nlof31B62qpGMzhS1
wJjHO5RHZQHgZ6A3yUzpYDT4s/buiE5iwVSYxU3KwAgbeNbD9eWul2BOMN1f9xlN
DlvQiyKa8+5OWiocThFi9YTW9OWRPGqdLQ+x0+iEEIvs/vyNQc4wYdaki+Zy9kQh
F+bbTaDsx1EfJ0NXOgfWMVfz7tv6z2Ch1Cm0SQrM2AcO1R1mX2KXRWHZjE4MnKLN
qXyFHdHd0OH7FoBXr2EmTXBJsE7jcQ7fRA5kIqNnWBo8cFS542KAIvSYdWDaUOLH
oEY2QsK0DWzmQpv3xMhCxfqMPZMk3Vs095GxRZNtrSkj4gy1qScQAt8rlmbmqcsu
aKlysMDzIxnL4GUlQAAGo6I54zSQDPaHKVccu0+LSZfHBQ8v85nqOCEVc+ERaRm2
n99VQLbokaA8wqxr/t5appE5EGVAbFwLp9QwxYBUDYtm4F4mq9vUD7Z+1k5tisfb
I8mflZCP4ODt34SEeqHaz3jNcwjeY2EXmFpJ35v7+Rxkzfbx/4Naw/f3sGd4cS15
MUGrHYucnaMjGUWV2/RCX0jaZAP9BRXNk24PUozcqGvlC6xI/lyX0ksNekGYXQSB
IB4WNhb3vch0XKph3UfBObHGx9fu2JgjvtE49MUcFbBtluMx8TnlU0Y0o9Diltue
fC0Q3gCg7nMDGtQBs1U/mfrChP+QRVz/EnF6UnarNMMabzNJ3mwOE5eZUALs1MLc
2bpS2Id55kFxNqIlHU5xzoZ0NNMG+w9GQKpqIerbkn9YY+hQCf8BrdUvnHG5Yl5v
9angDoobKgSunDehWocKAwr4NhgVk5iwnbwVEWt5K+eBjoa+2MAuwmdLXpLXJIg2
03B9ZCeCIE0Atn/zbz4FHoH/tQBWmcE2ovR0ED3Sh5UIQ8C21UpIkbkcFPj2gfCO
NawvRSxpFntcsoXWxH83Acs3UELCxncjTma5njIkKTcujgCmLQJhVOYBrDjFfkjJ
aTHWPGj7uHdV1QgfRNb0kdW+0uEoWzeEyEZoI+od1A0JtcGM4jmqa6mxgCiADP9o
/IUQBi6JF9mmFfDu8sQt5oimJB27Zg55x4cjBSOZN50+PgnS/bC5AeHKjHMgk44W
IHLYGzn+xeSo2XMle1DgBHroXPPOEp/N0sOKcdI/VvSwdzx7curPJvIeIeWdiRaW
C5kEG0rwEuU4dO1+p/b2Cazt/f/6/kQ2VOGyHj8q7oeUMQ+jAiSWQ590HWL3WEUM
fga9yKEEn27duTTxlv/2JCOI5wIFJq8Zdkdb3sHaWgl3IoDqi0n2Oan3sSUCqgoo
j1Ypid8hmk/p1mGzXCGIeYEPdNVDj5LExOD0/YstITfpiNC8ZA+jxiYeNODMscxN
qKy7/Jv+7mI/OEE5RpIY05pU2iEKxTcUz+iH/FnuPtDyb3+dIbQtITxrv8cVfs5z
tLschAp4vNTx5iB2pz2YtOZqf009w9EBwdpR9De0pGocC6b78MoHik+oHaFgnSvn
yWFkWI6B8g7ZMqyrxQDgEse8xxTWIvtjy9YHtVU/xtnmCo+/chdNWgC+LtprZaIZ
vRxGaeUAORfXd3AjnSWc9t+0RocjyoY58x6rznDMEiLodRkxNNmwhwSqZOcwV2jZ
6WWdxvz24BeVuyDxO8coviN1eP57RlRKLZd/IQUWxDZcp/xGDx5mmCDrIoTlU4fA
SJtUSyqQvP/WJ3ADdiS2wr9s8h6iLdSl8//ttXcToirW/rDFY52fumMywDAFMjO/
yFjWxfGJh4h+KCWGYjUin7tQ92xXq+KMIhVBCcskn6LRGWXXS9X0Zv/ZpVpbeeWy
snA1XyHOMyee/qEJGvrDa7xDosHQegb94PhfRYgW74XOZCBvFPFTh3SO/reMeQVc
WKYNKcKYRYRlrlFv7N62D2vFUtcIt3av7skdlWAB91hn7yH0ta0s84kpCEfHApZm
C4li7+hQQTLTKAeEaZbH5BYc3XtLPO0QvWLzmWe9QKVr9CTax+HWHKZlaKaaVgQR
1DZz6nDld9b+g/R9ZaWqZteI/IOVci+vHYmhoE03q5C8KNEBUJvQwjC/bO53noUN
d1oO1frw9YXzsnuICH8vrezbhIRHCrng8i+/kBO90sw2jVHq2ou8imCH367l3yNG
QIcaNKcxEuaG6bXQcMBCQbKN5gZJTZZy7P1cU6r57rBd/bOv27ZnuZMkbs3V5iPz
I6p3m1p0XPYNiAevfXqtEpnj1QACGRKkMTyqRExZDzsVL3XE8MwEwrFhI8P/Ck7O
KJwA4bCpfb9mNR50pPZ1Yl2t1TMdtg2gaN63aS6B4DyiBf+CHMAmaC6FtotjYK9j
3bmuz8Bl8Js7G60DRgMzNEMXUMWVVxkxfpQBdiX9wLNZITSVLDc/UiReh0DBB+Xr
81l7fgGHVNmzQWTRfC9kUOwt5M2EIkeHyeZX3SiPn0hxLWxDKjYnMbInyzyO6G+a
x02vpF+iYiGZU0mo1jjIPD1uMpkUiJn0tyj5xZ0RRyNtIwWz9ELT3aGbIw6BcHSN
1V7k+lTrtGTi0kotshQdPeDq86I+XlsTe/6rv0IWAekHA08QmQmoMgmjkb0BgrGt
x5zXOgm6cnaErrCRGXKwAVElr7aoOemjEWdfumyrT/W7yl/VlGET8ltn4lYDjqVE
YBWX6SIHCCsjEB0A/qMwIeHPs5136ATBy+tPmtg6CdY/Cgi7o8EkdYdp99zLwXXH
56e4c/eeLa4kWIbL09W3fQw923+NFbRNeyh9we4+LCX4Zl+cfWQAzyZRfNLpGj0X
ii8k3S/e5VfyszLboqsOm3hh5jsxQttMYg+Zw5reiOPcyEsnaaW2f/JUGVRr9ot1
GUd/SrZim/bo6086Y7qkGe35mlnsSkvNsjSF+oKDwrqVlaTWKLdByvF9qkHHrRuc
ZmM+vaPSTzRuJ+ppqelYzV0t+AHgxD4NrvcEY2ThY4JXoqvVHlO9LCy4cT8VUCdt
jWbit6qGoK1zgITi/ivtJUG5HxOJLZgxngWjgwO8DZYN3wotq2+yU8PSG290B1p4
qJIG4x1vjvFk0UE4Irpt19UUWo27t0J7+s+NF/bynTZMUjch4+OoZ0Kuk3xVTDiz
JZI5FfYRYD8l/LX2BXsdb1PbBlaR1Tyi1Zu2/BRLzifMVs+itNf+xd0SEydfWULz
r84P1bJx5JXyuq1OxZgqDHoB9LgZ1txpKJLg5xDFqarT5m49D0CmP6wdv4ijQgmT
zqW54SJDVDCEl+xhysCekU3K8NhO94Zuxsm2WGoyvlTELKIdzDEDQ9ZnBLG2AZBT
K9p2fQExpWULGj3UTCQDOQ2d1rTSYA2emWc+KiFCAMGgpR/XUQFWkNL3d7gVdsZy
9gVmdcswdlARKNq0zP6ei9+0GqBy//+kbget2xTb7NyoN4nn8BLex3jQ29tLacA/
eTcJ1Gp+2Lg6LrPEP0/EifWUPGY4+j6qcqY5G8DAJvQ/uR99efVQfbRUyfePqDzp
ec78ztgScl4Gs/CHdOdrZ6ljt0lRg4tJSmRqJkLX8V7D9o3BSgzXmQeOmO3ckj1v
/8SoVhFaYjyrzNXLKsfOnnfJNslUdhI3yGaYpY7Umg7yFvmG4m1mWKFTAc+su5Px
8VK3HRHm55KGKXBXk0XuEG3m1fvrxNU8/8fjcurIeRWcwcvvyOJSPzbH3gMET7qA
Xs1QUfnSMbjco5QL2BOIYKyBM/w8hkwTxZl0X90xlXxS6f9k0w0b1fBu+WS5DDdc
WvtkX+CzB3WlBEwNDuJL4c29T4em2fPzFc1mKQJmUepY6+DJmnUmE1D1BIwerPb5
J1MlXDWBGNXHbkIAJI1JlERlRA/YK0zuuvSbo1QiVCRAawsCOyY+qbthUHVdwR1A
vEnbybSdxMsW8EWv9VchfOjCg6PPje9WejdYygTdRlsq7tVGZ7LqcIwOcTgB+Ygf
9XeKBxGYn6TP4mW4u2Q+LVPBJsvi3NcFmnBb4BK0FGA+QJxVZVa2lfLUYB804Eam
K8tqDFbu0FTv8OF4K0jn7erp0IXQ9x3kt9rj0Tf1oWv9KFZE3Nj23ARFnHX5d8XT
dE23xxKzqbxybUmvbp9zm/nVU8NtTvIbyNiHq4WNSe97wFKnyr1Hf5vYD1bE4tRv
Ck25zUn3TDOigsde+mzSMTvJyaOz114WsnqTeOMsyE491jlgFQAn0vYddZRALeNW
0OjRdEotrRJLMFzR5glR8ZR5Gzm41WSDivz5m6mHIvD7sWW5uic1UvmWTcUrZWV6
iv29W8By5CE9LPGP8icVTHRdsiID/Fzeupk4lIGvPVZmKCNK8PTrjbPTcRayQ1uv
lYX6T7Vh0UDm+Y6DHch6qyVn0xku705G56Bs1ojjmGww75dZcVNpOyk2H/l3GAIm
sDgB0GZhTVlLvHUbtrerAs1K0oyt8UGt2DwUI0YldQW16ASshpoFJvLA1Hc8hRpH
+1b01enzFhJZA/yqKUKc4XCjQmZGpCq+UzYA6VofunW/vKlhCudbB6CxgLgjXh7X
wZvfgmRMvF+dbPAIsrAGr9phe5+PFzM9xhykBlJsX/6o8RGlFpam73G1/VmvLnX6
GI72oVR3y9qeTM1+iT+fhQ1IzR/+SMNGROuLzUNR8tpLYg02qA7fYW4IkrNnIiuf
m89ogSdS0qOMCYQCWfQNHoeNZVj9a01qDiTZ4WmjQzozUYq3V5zcY+91sGa4F5HV
0OMfkab1t3vP5C/16s8v86T/51XEdqj39fbG96SuPu8CMpUdgSZ85b/wDA0fFr3R
s7pIHL/NwCBvSG76M80SBinQ/QyHbd7n2Tf0hGWCEV5Qn4O8w0dkcYMKhgQRQX41
NvULhdIX3UAPIZVYAkJmnYj9u72kxYd/hWoU96LC/D4yIDN9WUwe7PPV08fwtOT3
CEZLuGhiKCBa7VPbZGwzZgonNZyCsROHy0oDmEGOn6QtanYUpFkvSsqp+hJqsUNW
/C8llIfceO1D9mhLgnJZmxvziFV82U2r3yM2tXg/kN2v0hhlmcJ+SYARF7e1jj4c
V26sM0t7nn+pc3rS26xVIyVJFtFL5l3E1t1jnKBs49U6WTnh0GFoqRi5osxdQSS6
XG2bheIHT0U8YnchRmzSTsjYZUtU7dD3pytP9/EzYwswWfKrFehMWdoY2sJZuM7u
5uf2GO6B3Jb81oG9Xmd94Zfuuf/d6F4pZE1ZyBpUsyq4fcjlR4fBwJuTXqgwP65F
Dr2nzwxQvci+CoWnrmzm7xwbAJqf1fx8K6yfg07oTdmHyFvX0UD2gfoaDJ974QSN
yp/GWL4oUPYiSqgtDXYrK3Zl0goMXCd8BtIp5JI8BkKBPb7JpadNDLQk9cZc/SOD
QbohuZH2/gyW/8xDbb8vcwPCCvAaQCBxXcBP/4bK0MSfcwaRdDUOqzqWq2hhhvdx
BpcuyPXPcJi4fY/3qCklvXnOrR2xgc1c/GQMGu5XizNk8gvhsd1g1T+iaesHT0LG
aDj5iyGMGS7gnrRg8fDur55hFwe8j1+esxDocSlCJ6x/s/I4Dw28AbQ9Voq3n9Q4
9h8TdbbZ5Edx0Ivt0b3FZ5WirPf3Ss4YTZQFsG782tZ9jDqqom3QZECcfUzJSeZC
JYqt2K8DWHtMaxnooXz0rL+7ZuX27sECh8bDkm1tCg6pudequW18kv9HERc5d/cl
v1hvNlLmdJ8vkyS2cBNGOlEukgYd4LEzUfmKqEx+Uo3di/IKOVdQW1WrYleL8Adi
wl4LD+LOETr4houaczmSRc5pbkrh6kQqolLP9x7vZ/2z3p23AL04CTW3pXWHjKk8
DHfmKJMQ7IctHmZCo0w0W/HFjFVZfzSEBSZmISV4p0fLxF2Ds1MCSi64/OrsykjJ
0z5k0cp25n+ub7yHVNx0QQN3Uijl4DVHaheSfptcUEygzvBSefFrUGkJ50gMrGgS
8hYVSJ0hBv3OKnqYt+LM5OWuEAil+/CAPNsL2Mu4bwQSa6l9xjTZEGPH39W9tk4D
RYZl8M6ZV5Ae+DT14eMDl5e1kjy3a1SttYonqi79Hl4jIhWO/XKApY26CY4gsbuP
68qWv/jiBFRkqMH7NYjGh3wODHd8fAuUjZAa++hHxbZvRTyH2l/zz5BaWj5g+7dL
pRultoHC0hNnA4rU9tFkJIzlZrpAh3CSCtSKqAG5jIB8mOYPXmPGXgY6CMkIOCpa
6vg1R6Vb7odi310ON69f84YWxrtg2Gxg8DYuttz2anmCvQ7UHxvq/u1BfOnfOJ4H
WUxwboQMhCA/9l/Hojat/6MbwxTLoKuobjjUGJrp5gH3jl7fGeXM5SdqUo56P1Kj
I4/FK+0dSeSuU8O3lJYq1eXNSLMw1qfqMmDSUJpxiayMXuMhHoU0J76WEhH64A95
fW/erGTL2f9ANfdPs3rwWPmOEcuI3umDS79wafS4ZlV/9kuh4Zr2BXU7d4ve6iXx
NNCGOcOY0AHSxO0ndpdzFH/NAO0H5vygZlf01ymzR5r2tc9Z1dUPsZIjEOWsCtPk
73xG4I4hoQDt9rkgbhwex0V7zWJR534NViJG/2eygeQ3zYu/197pCHeKb3ZU4C2j
EO4S2bJmHY0OG/a5gamt+P0sxUoikqdgIIkvZ4HcK/wKp5mKfTDJd8av9e+byIlN
pI/QN5RMJVn/mkBLHB63IJ0slm/MDMsN0m5spzmrg0aqlXnyQ2xQnBCbkifdpTO2
yzVYvaLYPm+N4aAra0NlnB1jsXAXfUDK4q4qT2XYZ4U2dYsJnIiNdXWIFEcNeXQV
d9zmsjTOsmoLryKsgGOyO8pJtwZcufdbkggd3ITMuYIK2q55XRLQwjkapo18KOGa
V4883ZmWwkF6qLurTX76PZDLiRmwJNM2F6ZmNZT3V0xU3iiB+bb8dKhNRwzhRdVK
oaNIu/T21GQNzh25pteh3JrXGn7joNX8JIl3YyqIy32sUlH9I93U94jaUstn2ZP7
oJxTqAIj1W+euv4i2grY4KJ3SGaoP3eRhC/ohhfkjdzEpjerh4/Q3jxWhaQKEgRi
hqfI9t3Gtuy5MEbh0BpiCqfhpI5gVQmAjqpP/RMtqPoXp/sKDCFDaRP98lh7qS9R
NzEYY+e6l/+DdQSQzvQ5KwGfy9S8yWIpe4o3S74sKKgzFtPK1p//0LlW9JqOO0Mt
gtr40Y2B2hbtB+84a90TgwGuV/ktA0Pb1463Cq1hcsHKRRREYQIXz9P7t4C/mIgx
nmqqcU5cXOeKv0WaRZHutvJmAytqIqxU4qGN8U9Hmy2j8a4OaVLIpL107+FsXv7k
hcNsUgVFnT+DyNTG14brB6htz40xoW8hOw6nh7nMMQKt+mNDlbuMQSv6ftFOgL8d
ISAdOqWSXSbreJbsgMVHvn2PzHxlampN7jpDoh1XBxVlX/h7wp5RPlbn5h13vxSf
BIzG0ZqMq4fiXLxZEKCYQPa3L4x1ZEKHdQMGWe9FxYdaKOJwC5WDpdc4HWozLDK2
h0gLnAOCgYBZLJ4uadNKJPDTCg1oeXFedufSoTxQa6o/GRiSg39h8FkY7+fz3HV3
rnSsL3Xy7tAHiZpu6RbktrXWuSHhMK7QnxBE71RipCM3cLHC0eFrIFQ66yfgPkOS
yc1OQYgA0rVdrwwXzil/IpODfzW4MNKHWzoiyACkapQhbLG40xWvxHrDE1tVXrJr
pqFX23zxvYqgeporQWVfrAJdYU2fZTJjgmAQz73WzsTTGMQP9ykf1KaZ5pBndue8
wc0CilK4p/qpuY+gumqtVfpwpoNQdcV6ukP1TOB/pxY2ZI6Ga+iFJZvom+3GA8EO
CXIF/gCBWCbqsh0y/zq+PDcrdg1Jfc+wADPDZHGSWpJy36PVdjlgU7s/GXnCNMxU
lFDZaiLI37y/+8cIxPk4a6r6zF8Q6KiJi3ppnshQQufb2i9yCqHzUg/LBImQ3+4d
WYdjvG43gtJeZMOYcTc9uPkoKyOr4kgtZiCVSGWtLidb1kblWecU7+GR3eOeT4UW
Wo1XxfY3bESoCjhYM3nSi/W1c8IiScGIWvo6z+p2q8meNcBcTKnIpzr5yTCcGKCs
hXXtjOUKS3y+5fFOc1qDJAxEmzWQBDJYjby7+YBMXa+02b/reg+Cc3h/n88OgS19
beU5jOkWGcKgYtzg9JyvgdNG6EeyBl1coSK3cpXK0kA6vw55YLWTP3CPA0sGVnkG
KEC9kqlXK2z7+j+BKBzyeQg01/FiumVAx1QJGH6MhhiLESLJXfPw0mtg80q5OTX3
IWSpa8QQzgkYaAcuTuTnYQeNHfiJx8lVfU9ULh86UpOTJOBEryaAmHRmclpkRsxl
MMkGWiC1KlFNtRqcRhgdXRUPOkwCZiibWS5J4enS0M/UF4vKL31kry/M4v3JGsuN
Vd6zmnFxTZ9U+XwMi8kZa2tSPWytsDtA4bCpcTGlNm5DjheRUkp9FcM89+14i5Gx
yiNqUp8++4pBWeCLhNWM5nliP0SUNa3/QGEEKnIDb2d3yUlmjXOYUvFQUVQCJ5ko
kgPLteFznhxJAUeuOVMp7UKxdc6UAoz8wu44klOXeYbhipFnwG+vqKSig4DLa73C
SGj7F3oxHQ2TiNQ2vJaGQbZjVlwXbM0WN3YlFKIUQbVUKtCExPgFyKqg0Mcu2XMO
LN+jtH6mFIFRlYNiQLicHY7KNnhhk0yIfMiIGgWchEPJJYm/V7UzfR/AjsHQDZwg
4h/QwPzrRtPy4FwONeSxYOoeOXjd3ttiil2L3Ol36mWI21UDCye3/w5g1ue7XOZw
REHMNPGp3+AUvVFrqGZpok7EXoOgdF4VkkgcrU8a7uH2lU7dFpoh5K1UvCjx1rbC
KUhI0HgwHpd7HzigIlzaLBNaFH69dJtqEtViQWffpzJHpZWB56W756nT6s+kI0oR
Z8MnwNQybuUVnPxKpU609ShdMxlOI50fZVamaK7uOmNohk0nqURFXN5P18S+RU3U
GWi8UqESaLVbBSWa7r/BhN+kevxYyBkRMPhzxb4c8lF6H75SdAq/cTVZO/sYU9nU
FeA22S+0QB1+IsX1zp89RMPmfP7bsXP7hRcuvve1aPrEXI79LH+AptXddc3ycr/d
LctzfnyDYLpIskjwpgqeyLYRVXwGgZy9QTaN8pWNVs5rgoKdDRK4lEECkBtmhKAo
camJzKjZCAPjxDw+TUnTgXo2snoCSbmzQKEslUIZK5Ko6wQNAW3tb7BwutiKqj91
3hAYwQQoTUIyhIG13dey4Hf8stEtaqebzCgVuEFm9g5gWTGMPovKv7MZXtjZfHsv
8wuvvDWJqpgkseMv0ErXu32Z9B48UbnHriL9n07QIWuFbKobSxz3waw+dUz/+q4J
KSjP7r7kfK08EQEOKdPlJWi3SAxva6VaXypQRw0P88EKcQTDFS7qmPr5Qjhx6H41
NxHFLOIARUD9PeyQoCAr6GHINxzmNU2xSMo975we7JK4+zMMA6SmZq/7xThFj19x
ZiUj13wk9roqCURYB3lOScpYTKEnQsvecZX9ELQ1p5sajL09yaxmRAfpHCswj4et
W5JnctpFY2njFO6ND+33+SFI3LcQ8PALEMueuSn5LkC9I5hTIAThevWtlNUrq7nB
2DbRTE1Y6jtEoaB5aRG7h87iCBg+QQdXIpPv+edjzCEA+Eclv8TDPnAN2yik6c5L
5LJfbxEx5k2cJW+CMhWgBDBVt2hfYOPodleGR1mWbCC59l/ueAV9guKCFvzy/cj1
cPy2GHBsWezcE47TO5qQ2wYIyBTTRlzbtCA7Iz6GnjIfnlKrAeKA2YE6qI181QvW
MS5xAAvTTjD3aQwLFx4iDtZ99LHb+KuX3V/0Y1XqmTO/mCGlaFOFBDmzGheFm9m8
6UV79wCGRmZunR6UlEvSic7FD6sL2hjEdHU2k1Wo69Wlq+1LjIzEK3ziEHpziFDV
Ou3/oJ2VzthDiYEK5xiJjsJnBvbSTXbvUio0COPXeXlB2UypC2jOdm3KRNvNHZJ3
LqSM2mLGJwWgk/IY8/u5wGQ6UIGDNYBoTTXUax27Vfcut5Rq38u3z4gpq95bNX9x
2hKf4aOgZE9kxoKaakdgHjZAyfi3pSVNkTdJO3NNubPuHd255W59x4edMelRmAJS
TKDNydya8LKYXRJwy3ES6Ilmmkssx7XM9aJ0jqI2gUcEcKUDaEhfMQF7tKSSqUL0
c226VT+r6mAkdiXLRoibApGY2wBGLxS5tpOujlKOKc+3YvzoOxgeXTCmoxZ3B2IN
mLOnhBC8SMAzp1MjzTWHzpJ9lOnXrJrtX7IXzEqEwIVkfgK0XQCYyix5N6hueiMQ
64epd2o4nRGEmTe513XJk/8rd9I4s1xnjdlOiFHBhYg5Fee2PusOjNs0osVu+fXN
/I4j2VG0wDbOKVj5tLqI8Ybaq+0wR3+uQfKG1GZA91cnfDzFvAzzjPp/k4q9U/v9
QHNlpYxU9mr2OpUyNPK/7+ny73N0ixe+PPwBnzt9E1REqVbDG0y3S4fxYhIyRJv9
Nypm6qgKa/xlPmHUnJxVA/I/7GYRII1oNmB+g2jFSXMVSdKf5OrwFXKoJI4wxTJf
vr8YsvNccOVMtQ5iWuRrpE5dYsiqUntwHNxgGfXP2AdskA3ty5KPrAFmNA0cfLOj
B0/PIrE2PH/nm558Z8Qejy60tUsqMu5bCyuYH1KM6bvuKPfxGNa/cDn8FClWxgfX
Xspr+s0Op5dVMHJZEpaEdq+Tmw6Bgt6bAV4P/nTQkPMVVWTFTA4qOL8+cIuZnN/o
bjR8k4jghXL9P48aGPvqOtraofAbNP8Sht99p5E1S9vcTp3TBeWmFgGTZXLBkThz
PlTOKt06E4shQN7Is83ktN690DeQigxSL94ZEfoTFEEgqdDPvCmzDIK6ORKSpESP
YD7mWP7OUEHdhvgkdG5hLRpeDwLUzcoBuSoReMNKFMNpHfzyyNxFUew9HOMLPlUm
XkX0bkgGuE3Kl6SrebY3Kiq+AesoVm2Qlm+IyaJWECsO9mGY2/8yMd7HJrl3ozqF
9dP3Xw7vZh/51c2K6sQ4Wioq+Bnd6wCgEuRGEvhw34Xp2fBUtgFvrOPniLCvbmhE
CP2oi3uSloCWwG4yZVkfepahV+ikYbVeJUwYUx+oGbligPgYBSccLHzmpcgL/Hg0
Vv4vA4GX7z6qQGLRXA3pTGq36ZOcA3CLts5GrsUNlH73KOebcqsaDbbPwite3Wl1
9Zyl/xr2RwmjaJJva5YvrjX9cZQKdFcci0QmWeS8+EBYP0BwiGYvsrcz8V3yVqW0
B1Qjp7Ijcw4OmwFfDBFKyEoqzCjbgAQEmfbseWKaybsqdWq6//lh0jzpnSBhnm/2
kW5QvX2G8jFlZ3fmRx4q3JvH708cMO2bL08HJwmCQ7I3iiuiciXTTrBE9PkehgNc
5JhDTBpadKawCAFqviZrgKobdSQUDDDz5IQ8+s+2QHlmyAghMnxLi0HLM2TEYJ/9
1CT6mW/DNgSgyKHKWHVxXNPqMyReUdKYtJeHmHKgrBm5Co0KW2yzCJPu1YSjIxT8
D3LUdzlgPngEH5jDD303ZTbV73loXARMnvlUvoc2OYgDeXX1Df9YCefPWpEy4uTk
UXneiK8v6TwzEPzzC6SW3GOPFEkdz1BiPv7n+huA73DhfW1ShBXkSjBUa8VgnbRV
ntTDa2xezKufMlt3B/AjVf3jb5PfZSwR5SKqi5fLwWp+5STLvVS0sAoo9uB8jhVy
s/giPeVhTslP4+2zIlC2VgUYXxq26zr010uSPqJ8ri6YVEtxQGN3GR7c1nlIKdxK
+r0ZcaHmDVatfLSMJadR6B2fNi+kNMrxEhAw6U72+9LeqvPJXuj1dyPlfVlxb5RG
wvdyVP189cTibbhaoPW6TQl5FwoqFWC+NF4xhFiobxKLD6PwPpLU/k7HEpVFwekD
YPTognzHKz8slVv+27YL0LeuyyARu+LfLHscyfMFh2DlpLDkmgk+j2oji+83ocb3
saRVDgvFaZghiAz7/sdf8XmP9G7SvWQbFFhWZTeV2V8jDOFpXTMvHKTTuZpMrnRf
UrmmCC9Kn1AyYZteubkUy98uTkMSvmMoQP+JS+H9l3KsJ+Fk5z5VE4slls4IKLKa
o1tRb97h+laQbPbLBuwzl4sO0WPg92+dok66nxSWvoSMvIOkWK5GowzNQaMf+NjV
2sB7CDpQfwCT/5HspDguwY66ta/ad5A6HID0wlPVDGCVjUdqsA3dQZOqQYWE/FIb
021pVQrojmV0NT645jdThPQZ8FUt0ewVMw2TzDdurh613lt/I3lktUoU1kjYMRK4
dmHwPiXCtVYLhW+qcttOZN0+57J+s1hd4MrDNDrWV2smsgm9kWFpsgY2PAQ89SKC
SuWACUdjC/of1Q4GP9zgsEEkIHHsaN+zdL4ElpA9/Z6QMjhaEc06JVd+jRqsqPs6
+DGDMx4lNhMWrW1DWf7Zjnic7gY/oq7AhFfywsNtVjlLjTwvfgyTM22NcgwSmw8s
yzuA2kJXBrs7+OUWAvChQ0FzR9a9YTl0H7xE0n4jSYVrWV7DXldqdGCCQOyQAO5b
3GC4ctmBp11rMns0vCfYzXljV8oX2S2iaXw32Jt7fEgm8j2Ke8s8xxLzTvtA+mOQ
bU0blm/+bq1RKhHKvMiV9G4fxQZ+gKxLrtbKgHRSqzX2jQcV8jkjxyOmY302Pz2f
ZL7rTOZSJPTiLb94pV/o8Gxlw64mXv6Q+THaqxLfJIqIq1olZ18KjBvfsAKDEQpH
v6rssak63Pm3+nP+DcewF2wa33eI7LOv2J37y+XAxJ5RHotQ9zu8JQTAIYsSRtka
E/m3B1UY4MxNFlwjFz2wIUc8nQIujsV2bZioBjVBk/yRaJvLQs/xEzdKQ+mms4Wc
3MnMUI0t5v5kA+iaA4pj1i4irX5StLIzq0DlpECEJjLLuEmqbAgy4waCWMUayEDl
tiJwnkpIWCa6nu9QmcG0U4J7auikT/aJMsJQwzRZ9lp8WOkziKlT52S4BBthhrNf
l+cRcEXq+Z6FxZYBobtZkSpZ3Q61xDrpAAku7s4GMuURTB4Wmj8jjoqwpva0M3cG
FyV4PCGVL9OkLe/72uv5KaKgvlXZaCZzGqJ/C7JGqcvWuq8gZ/uYsIlgUtAfp7SG
9BZdOJJba4ZXMIlLkEBegqT8A0sovnMlhx1/PZwFt86Z80/YVd4oeif9P3tXLIeH
hAeaHW9TMcSs0K3VohXloJLB+MOJqLNqN223MUW14EpEgCjZOnv31KB5gUJBV7xe
5K4Lg0ovOF9La+bUQhFTOcX+2sFc5tmwdHBv/Yz/MyJ3w+HFjLGFahYs3+4Zb1T7
Py+HZ95Tah1UmdmSYkc1qiRWmA80p5lzmHp/jUFFFiG0XQSugTaDG8tmByGARwO7
O4LuTw8mDAzHPJGRV2uc5uUD4fZ6nYP5v24FtTDaEFljBJALJz3HaRB6XFm2O9O9
kndTDHHEuEogio6zMmPLNcmNKdQ9fvAcByUjOf4POZZzzixHVed2sfD12hQkKS67
cblEkqTz/GIxdbxblY6ysk8m+Widbt/sbgCHCc6FFIx/2dNZSstyXys75G716BUn
SKzo1szvCYH8CJbnhLVaab2/FTr1BdT/LQ7S0f7keA6Gp8NZgMGlqgruXcP1J/qt
ObHksS2rzwgG2Sx+GPyO/lfYI/rgG4Zfsu/ctq2ydHWVWDe4lBE3CV9l0XXbF1o2
RJOZoPWq1+CUrSwNxtjQmxnjLhjs15E2YRZ0XFNMm4UHBNJkKLJJgyrYiGYsPz+a
hdh5VL0XiOpfpe+UleHqnFRVNH3/Sm5F99ocPfXvSXJ4IlczZEjMyOJAwGkRrp2o
lnQdferXPYLp22T2T5e9DbQou9Ml55DKhzzfH8BspdIegFfzue/XssbU6k1xegup
sFTFXQtCc7exuUTj+qPUw4iRabgsOTwyOtxBxWBwe19t9qslzWEusvBeWe6cCDfb
j/Y/DgcNr/FQ/he0rhAOQiqTDDvBElujxQhK1WZVSqkDMTGYpGMi1C0L1Ya0+DT+
Xbv/Lt45EE9BMz83D9Svlq+dP35vNArAS3Q85u2ABAhU5XUCNTUgWgnSR7wvjPdp
uF7448Z8Hxva8X8/95TxjtFmnocIDhuS3QE5z8E0E2ZHWFPfxd+vD0etLXd2x1y9
W8q6gioN26RhL32S8CQzaUD+xeee/qqLKGeO1K9BO8uSIvNwxeM7oaVpQaS0vCmg
KMwkykoJKb+9FByhjUIzFdjqi8Y2vfnwhmNyIrnke5Ukb5E+HbsgSw6AtxiAH6FD
+IvCaFOhiT0BNeR1AW0UzO6hc2j2KIyv06zmsxXFpeefulWKh40XAkY8q6GcvUtt
wgWVJGot5IqmF4SdzwoKvhtbrNdkl5wa+6+NYlF7XhL2dVLLtzqv73y5oLUTwqdN
nVxUVWwmjU5t7mSZXgzASDvsC8wxAoqJ/pr8bPqTXcS/o94Ds0TiPCrUfO8kk3al
QGyeIEhCTC2mmUv4Nhf0EC/Q+3qzX3hofnP872EZHCwDZcgo1KKUKuMVoTRcPyg3
/qrBi1itKiixTqa5dlJB8ayTAOp/+hxn40EwN8tQhxEOa++bGlrdNnpXRaLq5bi1
G12w25aTa2/C1yQQSdfSQQUUfEia4lTyDCD+e29Tp0j/7BZrbIkck8nhxkDim7Cp
82t21D6B8suP7DNrZiQk33T6rnUFvzkFpKtIDfjKtf0bOOCYo+MFwvr41KGop6/w
95ogPzJPUGPwR853R5tXmsQ19GsRMhG7lpGJWVHd3PnfmGeA1h4W8oDlXicwHmFm
OIDQcvdavQheuQEvxm/NsI1rgSA+cjoVmkUS8ks6r0ijBAD5NvTiHeLrJwynNthH
riXo0LRSVk2pqWHcezLXdUcciGsoEtKyvaYYr7KXTMyK4vok2xFSTMqAMmwdj2Hc
NUDlAjRL1jg0e5QCyOZUt9YpIKL1zZ6ItnOAvFaXYF/XxPZ1eoakInZMgZPdOmUB
pidafs6SUZgLuLR/ZDLxBujJmBe7Yw0KIEanXfaSJOpoawpuXeWln5hpJB0yoNZL
u6MBpIEPIQQ5Ytjv+c6bUISrKAqOUTfOwVIeIsqpQSfYFAeqkj5W3v4PP+psX1g3
iCVouNYTwT5tv/gryG589kfmkz3PvZ9poAFLl0Je984sRnmYJTTIInApv5G5LMmV
oPLxPsoSzmALkeNqfoWUVpdw8qQdFjO8/2ueb28+mcKSl1jOOu8YpjtSaDkLgw3L
/AoRArNhDNw6R+HL6GWRq6RSQTrWHmtBy7JWodhPbTaWuWPMH5P7Hb7d4N4KQJdr
0TO34aQD9e+UT10sPizRxnkZLPAX50ZxLyiAwhZu8+Wnyy80nLxrZ/AHIY+7JVdA
Xx3NgzZnHU9sOdGV62jW+mXp+3yjd+Vi/ucgI9JBLdCkU+k0yPIw1uKvWqk8aKEL
VwKkB/D0TKIjLyAZI37B3ZM8u4d7FXHdXa78tQP1QOZRHqvOBnB/mlSQ/Huzuk0K
rdiVrNXgq3o4DbZwpUzmDW4w+/ppXs2rBQ2Il5pAtB993zgdfP1N1ooScbJQRniz
GmQHxLcL6BIWxEL1zQ4w5FlMBHWH53nWvApdJPmSPBhw2FycUko671KI+Ps7NQQL
nY8por1p0SFxtVZKUvV18N7oni5jV96IYY3aIw3LXLICYpQZ7EFKLy5YEGQM+6M/
3J3gd0U7vENmKjHtw08/jbDfTDpkofseMvsY19jTnRsTd+U0SyjfXkcKwb0LpKCz
BGw7e6IG6wzXufJgO7JuleTmyWpM/9dHrcyUPG+zPUtRNraO+FrjHMdSMQ6xPkH9
uJJS78vh9ZJBNBrhp013HR5X7cjNKe506afVkWwzYpr9IWjD6kME0lGjw+IBAqOI
ZTsJWj0zFWt+y7JLJvU75ugHRWdDpbeh8DAlCUojONIrJbYt4YEuqwgcKSH+R0Cz
yaCZYEnNmiDnswgwNL1YQ+Jb/CvH2Bzfz1fyU0w59tBbLs0ioWibk6oBoXBrb/vv
moAAqj9IuFzxkCxw0X6SnUULgjwOh4wneo3tdqPku3071RMWqjzZkxN8XPnMd/G7
ZFnybHmapcDiyrX+gecgUqwxoX9Q6mUMmFMYmQwdFZAJyRGMkfeMj2bkZ3B3YhQX
Cmb7K71MBF3b8xvA8OqCNYUVX5ugCwiKIc+jIzMXzwsPRzYUIymVVoL4ymkzYjfs
cy3v9a/kPt6GTwGW1wynIhneky3fTmtnYHebMXX6EuGt9R/8MVCQoY2PMIHDJXv1
Ezmtge814BV/q0vHalxwSuUHXbc7AxcsedUSY5FjUwd6rzDFJgOee5zhHxD5SjJe
MgHPrDhrSVNSgAxcHSVGITnhzF42n3dVvJTAU8bw3Jar8+qo5za2a61QGKoqgrEW
2iE13m/nP4zNDSoZ4YwkHyZluhigqAMJQqoP2a9rOpNGV6L6AeIYEljYlPDR6l3m
Jlez88KXcCmsgp0zKwQV4fnIhESuztEJaN8+utPVC7AQIw+0iD67VfLguTRbj1Lk
PDuS8BD/JY7PiVX88ZmD2c2YpiXRdLiBzFLNlEp/dmOnaUk0j3Ytk8S7FsMTfzAP
0BIL9gQ6oZ9Z3/UnusN5QO0MBZqW9j3BaL4vwE/jwiN85YjpBIofPNlQ6TUwt/C6
f8ERS/lZL3suE/UlINO16U+5qu9gnFRKiDggqvKWt3GlzOjFK3mXyYnciOAe+D7b
XkvRDbZ1uuF1++CCcq/D7bHB/azcp8NF9XYxU10jeg+5p6yCqTfMWpa8fA7zLVgK
rwYAHrcwPmYGjcj+2BGRrprJ7oe3F5+L3aL05hyx6HjNrRvXokmsSPk2auVRu/Lb
RRYNWdvoK7iCqKR21hjS9FwW8XEmNcOjORJNSRoh9sb1OPSPmRGv4EskwqOMLFh+
SRID23fyLE7v72qjs0/6cFuL1j+jT4/qs80iE5bCQw+dgZ01eARJmOXGCZDpGm7a
U9yRXxV9tnnSmN3chfUwCJWL8dRMzvlDW1HPJTjg3rFo9qSEc4e2tjBQ+i/kOx9s
QmeI5RTrKANF9idOHLDGiZcju61++4WdyEKyx1vp1OaZLw232v0vKwItiMF8uDwZ
ysfE0HWgMowHtyIkScG8kTRfc7BU2nd9iOGZv/y0QimMJSn3+JM6BA4PQxnwQdID
m7hxr3P/vD4nx6QmWVxHjQYMrlpXfh9jXMpyd6MmuJyNR8giIVJdUyNXRX7yc35G
xl22K69wVT7j63BkHKyP6SKZWGzAkzt9JeBw352W+xT1Jd0cdPQPgpW51hWQlWPc
8oPdNQCErsZXAwtkg1rb8FuqXKyso9Y/7Slu3R9M+GLJcGWWXaWrBHBOO4siLEfd
WrWmpGorlETZAzDiSnuv/yOSUhavvrhnSv+NAq8zct2TOw16vLnjza5HRAy/E7kn
kQdrwJGoi5sNg+TKIhlN5Cxi3XiXL/UMBdL/VysgqOviPmyPkp0JlMSKGGa2tEFC
jkXhD8RCizU3CDs6aabi4vE6UFxpdOg7UsMCDf7BQZZdB6ZCztt8qrj/2VMX1vJo
vfVFPi4YcBRAkyJapumtq8od0bDvFoHFjnnphsWwfwSDsYRUuSsoUb/tU/FehF9R
ndUHIyqpA6zAfo0mCjAdfGPnyepORXVBjq2uP+/QT3oce/+KrCggyj9IVDvWAAe6
2KCKlfbwQ6D1mDbYHCUZJv4uv2O3nO4ZUQnz4N6K3ZHjGgR7BLBewa1qSpmUm+rC
fR2CPpKxgmfiuiA04Nxjbdn6xl17bkBlxzi7EOs0c4wki61iRv+Yd0BrpyFr0yrZ
5PQ9SjbXT0VOexQAur8FjCeXvuA+3GqeEmEOr0KoU3/yxGIucosodFMIG5XWR4K8
n2NKb6x0DT8yka65x7ZvaJYEMNfUkWhOaa1KFmSRZrPrv+3EIce8ct5Zcbqes7YP
KO0iQvF68Z77j+Pq82rV7SZgxHQ6wQ56istUQ7hF4YBxXVLTJautr21cY1b9jH32
U8BsUvbtebShoFJso5R8YJwkMlDojADUJLLOSudt+c6ZyJi6g1HV7c0pzvhb6Ho7
PF3vTI8HVbz20kpQFOfWFgvBpvapgu0X1HjFKiwBhdLJLMSF2HgWuyChgG8CW2mt
WqbVD6VBP4BcD6d4ZqfWx4+2GHWQbcm2fYu4B0ZjJLX4nFBkowtr2HjEPLa3zYma
geHYpSsOBymRh5/goBaS5KN9NKGLX5FJtodBjFV4qOyfEclWthj9RzhvE4d5gLtE
NfXaFHRCMzg05PtTM5LSHTrjqYtavTQzYF4WWH9OVvr91/7TQ9VoXJNz/pdp2feW
0Eb3KNid587PmZF4YOuT1PrurTZkuofPO0xAuAypwHEIw0daqyy5wVfZNCrmN5f0
Mrc98aaGsrofL8Fr4JLqOi+UEhqxi0uXSnvXlRPBQRMoA2uio9CnzNKQU5vT5ol7
hSvj8JfuTsawaqylEndSjVQifytzMBG4KyE9l784n4/rLF/3nGiFEm2WGP5SAsVI
6ciRRr8GcF3IkqfBnLavZY9O6Ui4M4sGTTJnU9vUp+B7J66Pbi09nXKa1fOdazZK
u6aFx6eT/vyOaLrAQ/F83tJUM40wbrvC6FsQ0RQO1n8Or5BBvBSwdzMNcID3BGCe
LhjOVEjraTA4LiJHq2AWTK4Dryfu7u+OUh9mk7bfOmIT1cVZxpnj83CrUYQ0+2s9
hxDZxie8hG0d9drefCeFeYm9oJ8+ngfIb4lPc7YhxKSCwZBCy178EBSgctMFF3i+
TS2YgNELF6K1YbvnYFVb6PGqxXo46Mt3Q6KnzXjHcyfFYQCl1AWYorqpL/XECOX/
XNd+AezIANd+qN9RrBxvuRcD5x5ZqdvZXJ/inK8S1cu0I9UzUQlE5XzftW/E6M2N
IhXn8KxWlf++VgyixOEk81IER5Y2sMmag0NhZbCn2VCAYMBF+04BbEewNXwxzldE
0rfOoTonV7TxDtvX0gTc+lifEaC2kg9w8DXmNpq5hUkTh4DnWyVCddzUjU/CMf/B
g1s/DCLTZJmdG1GVT/RYsrRsdSb9z0IAsb25pWUFJqK0CEKJ6ZkQ+o+f3tBTzhP2
UPTtXmdgK06sjLmkL6XPIE9eXb59qPfhrYc86ARVxCi+b6bV9StG/99cZUyqSeZ7
VXKnDwSmEWiuDGqQC9p+tpchTqweTjcCzyaQf6LyugoQEvUx85JNaFz3fPniZKfu
YwTfBm/eumKSDFu72FTrGopuMkPcwB6Qg5P7iuMBo7PJZxeQLu7au4FKzk3DNuFX
M6/EcdFtwXGBrqeSOoyr74b1KBQTlmyby5Ck8Lbkfte2n5w+0yJW+QaMArRxwhqi
aYPQXI209Q1Uifr+nAbynDDT25UaB3SZzQEddZ9/01KOP8w1WNWegHejPJX0fd6F
z0hrmVUM/NnMVPpTJ2ra4N9uey94qo8ktMcl3w+6JuAtdWY340y5ZTCjWv1dL4gm
iKTNNTd5GhN/tefej+5W23vjBV77GVMhlLMupiw+y7ICop9TUXUV+eqvvYShmvuq
JTkwVu8nkybYt+x+nY5aUR0SUnWYCK2ovJ7UE/hA4wm18oZ6O3QfUswSXBA8paBg
TLlwGjMAau6ejWQNHOzWLUTILpsTlM4ya12O+iBwdC4J9dXANE1RK8ktQq1T13Yj
q/sAkI3LkxOOKRrpCKvN9Q7dG4q6sLlpeZsDCFta7QYOsgDlIz0GPnSCXnyxxlbW
kOT3tXQarQmwtSRiOB/8wJDvlAIZz/ib6/yWYxPLEjTmnmXyd4VhjszYs0lqB0q+
MJvWF5eswbO0Hl/nfbfKdE66E8XH0MZM1J+aReutVEPGVAfESqVgZxESaIrmfj/2
6z/X/y5utyMXliniXkQ8XBAo9mjcL6rsO/E1p5HN+He/J6/fA8aPh1cAD/fEgUT5
2mxBMux6oCMtD19auilf/cVNnZiPXhE252ksd8gC7UJGVskk2Bri12EuXZYqMf+g
EtsLQ23sjh1abMRtwf985hn9Qok+eyFxD0IU32NIEH5F54GIHH0Q5PRIhB3QmH7Y
/oyklk++pUmpm72RFfptZ0AtEPoccXRfHW7LYbs2Tu6voUyFgdIRWd2Z4dVwP/Un
I6qtBaA1+iewtQBUSf2aStzignvMZfM1HJw2btJKWAnPp4JvGA+EB9m8u5CbX4lt
T1VjznMT/ONtPBVw+jBFjA4TGGzcaclszoHrYkaWGV1UVWC/RYoDrxSWu2vtNvP1
Ws8PXMr/TDOVkjio9i38nmv/Q7qS5CWTVurV61iEVn8Xt7Do/5sYJtTEzEfP8fKE
aN34cASwZT4QgBiDfVQxJyeQEaoREHhBbre8NxNTg0h5B+UIqSQNlbkNFYW4QFmI
2qAgnmInqCxxGxvzlGrPV1jq0se9R7TK0dlXOdT7tCxb4O7erKj9e/4cp3nj2Htc
5blkzw7KfypCPjqHQFD+OWbbHG9iC6lx4NgbO3q547zdqy556Onp3HVm2hVa04dH
b4eZYIun961B9QrBXf/fsN9Gp5EFl5nvu6tmzfcEJTuB8cENzq8Pe+eYEHBoyYBB
67zmvTc6rWD4NfNGDev5y96S2wUQLCLn5pZTRJiq8DqAQJxwvPbEYm7M9gLFPHDr
Qz0izhZ8ZkhW0x2R07mQJIpZVcnSTsS2J2JICa+JN5gfRjDviE4S7ayeJJiSjDtP
yYX+oppgB9hDHY/ioXN2V4ALzuJ6UdnTyCUjPDq/970K8Xmd3Oo1ba7gX3jiMlta
+0pqQY5iDVUNkIg1szs+5UwMSiIixZGwRtCzbZnvXfqnhdTpwfRDu2z8vYxkYkdh
x+ODqN9eW3kSs3b/7xWKeQ0hXfHcXyCQjtz2+QQLKwy9XnjTYnHX2c6o/0TaIWRD
bY6TnaKAPpaeUcGHghIvXJp060r5tkvWOUZH9i+zmmK5fpkwzbWN+kmEjXpGtmu7
qP8vwdOcPCm234h2uDPQksmo2cpqCKDsU5ra/XTftcj++W0cgVA28OGbZak6BIpl
KEpBlNhPYPwO33N6CKM5lKnOK8hL4yRhPF3coR2FXvIHPUI31KXOnLuWrmXUPTbJ
n7ZpKY4FNL4OHrqaX0yoNlzHny9TZFdEpdtuCxqH7TJxmFQNXBe8eAKVy/bSywPz
f8f/TI+sl3m5u9qdZ6IdGdusJNpj3mTt7/2Sp+8Rld0ZySFOcvfKXXYT2ADvW2iy
2m2/iSIvWPOFL/JPYxo5Y2/MXuDAat2tuW+dxgOURL897zVqHWAs2HVZC9TunV3D
wsJ87vjuhVhPYhpNUVFpUTUsQ2jxoc+isFl3+TdfOwuPqB/eeYqmY4D49d04TP6t
PfNamLepddqMbVGWp1gKJievY3jSRPPrHfEHuo36uprX9xMD1coQGYUNfhNKZm+c
KGRRJoIDAZtUHxnuxqk3esEq9lZ+DdbzEja2GJctX61+TWciPZ5TvZHOzpDXeO4i
kx+uW2BhFZQNYV23wWPO/dVz1fVkyAT54Wq15I13JxTW3YafRXeLi2FGZxYOtRUR
JY9pRvph11Rs0zBhC6X0I+nyPrhmZzDYZUbUw5ChQUmrSFYdN7Cx34PvfkmAJDN7
wHxGJd+NSdgP4viiWWcB2OLxGkf2c8PPN5oUg8D2skZjFv4cVsoMwxp8obfQxthv
JLOzHeVp/L1BzYjq9PwYN0UFMfr+GnUClv4RWb5i86gJwce4JDW8PjbPkPNN8gLE
lak/2Ad2AO6/lXJi2+JMB4mjclwZ024r09vVYweZ/pk6CYhTxsPJvvzzwH/DtSp7
HyYLSZwXjHlhJYDCAy/daKEZUdPzjkvAOjZGEmHBACHpjH1BBlckf+WHwYOMiQt4
0CWM/TTL/2vUFr8Lxl2z1YlRtfE8/Nl5KU6VKJ0z6+RWiNFJc9/pECqhD6l+yUQX
1X4Oj34yfXi/lfIdqcQJ4tZQWwb+TOh1yJq2MghWaF0iH4bZ27A2sbQt+eXqhPt4
fMUyvotNS3Ib9oQAsr2zCeX3LBocf/wAr0IjpN5vXkjCIU/reGMetzWBJkKxSjWj
EdKvBHRuz2OAJZ+zHyG1m4fS5MxiFwU3qqjX45nAsXWZlJu6nJKGOcPNxhbIrQnb
MsLgNSkqtlocgURIyka/zIhAVaM5rGtOhFqnKHlTfxOtcKypmwDfVkx72adEOAjp
eKNCW707YgjK662b2s/4cNIHf8gt1cCT43T540p94lvQc6GmIKDNxU9+M4JlaW9t
BkoH526ue5QmWjqG9GsAFeT0UjjAt9vUcXtVeip3M8AUMXb2SRDwGl0H50/AnQyc
lPH4FplUlDUBnnSldo9zr4Awfm02deKMhIYYvjOCBmjx8IiNIpVpiIp3DF39M9pp
dISncA4MxGy/xWDU/u1WDAiAcmCsxjb3ZPwDAYACl29h8ef+hjbCI4+valc0TmkM
BM0jaf8ShzRggn5zXfVFcYQ3fo15HmEYKA4Vr/tGMCmAMoWR+wQPn4Ye69M21DsO
H+deypQfXau9C+H/Ikm+/+f+S8tP8+nZgYhYjSYphjactXxHXyZCxt/5UyhpBx7I
xy/doXb3NV2RDhY9pqr30it2rJDg1hz/a5SyPSJA63DQVfHvnDDHllONgJo1l+5M
j2CWrlzo5qu+Al0FGGfnnIfAlx5D0M01c6cKBRzdj/kSa4Oqj2lhyC2bt0SJKLCX
goWCTHoHev1MkNj4FnPeqCCLrMLNBVkbn9ANfJCdchAWSi7FCC/plFyVFScDYp6I
/Fudxy6DXVAj6I091Ne9piFcTQrwx4JfqyxB4U664q+qPZrKZTG8IB1dabjNTNaQ
BUcGK35LEHs2Po/J8EGnanZIUH+7bHTDRfUIOlkoE+T43z8ysMnUNuVGLl+2auBv
EF3rRnCiD/zReLv9PgEcDwF0Srdo71/p7wpX2TNtfKvuCgnpmL1Yt9sTjwgGM0rH
GowaVo6PAqq/wVHspgT61IADUUeT/fqhfP+a1HEpZSL1v77L6aGXdz1pSOF28P92
tICdRo8SZWQ0yUPIkIqfF8AbSBWrU2Zqx9J/moOAJTVlAjSohWk3DxIEyk+zzHOX
xLpQFnlLqZ4DKRoMQwB+yfMejrzWpN31sjjdtc1JbcXKwKW85tGf8mTcc/3CCvpQ
3sQ9O9Zi1pr0PhkMiNxgmwe4+NROZ0tSIRCcWe1054Sal0hcmgiGlHWURnNA3F61
nA65enrYgDYmlasC97QBQaB1qwxWgJNZWYmXQy7/WOwn0jc4cLrWdkNNVZNTcIHp
PCo4u0yf78lNO6dUAQ54HjFVyaF8CG3ne6w5useJyoMYSKNFZ40Ily0L5WOB4xXE
iWrkfVt5y7PJCmFZqVby4sPtuZdN08qk1IPbj+wXpg/5BJBda599mcTpLxKRb7tB
b5ev9AlHh595i04i87Q21eJFYxPsIzM3mp+Yp+XeE214AAGiWMJh4DZ7uAyd946o
4ou8W2pxFyCTrfPMLWueipmVvV8PMga4Tz68FUWOqHtFfLwZXmiAGTMyjlWbKjqZ
WZ6scc2i7CtkdAAoF4F76i9WJLNE7vGZstJSov6Aqe50pTfMSyJnLjdzHgD9IlG5
XIFXMwg4rcHeNyQERlQi+yEaKC9SgV8D9U6ZrXinxWmIf15nIhUYO+M02dJNh+Qw
O+uN9eG8hn6MG4LLqtYiFCTfZcmH+XRkAUlPo0Q7DAlwykXwybm8W6M/sq9jGy5u
cFPtHAyshBDuNxZ+IX4jRDW+ibD3hepLA8ocyIm6rQj6OO8vfjg4Q4VoTzrFmXR+
VCxWaLzNsK5TWxEeVRFFdDZqSN02YRFrv+2Ca5LfELVk6jjysw4i6VocusvSUxIC
SwitR0ceVTrQ80irq7VLU9JBWU7LCQX1+CLuG39C/MzAKLOhimYq0vXUMwSR9pjn
0BcLjFaQcm8xVDGiBwjhTGoKTg7kSeItBjCqvQ7xgC6TDqal6j0EizKK4Y3SDuXt
584Qo7quV9JcdTpvTHZrCjEsWK4dXO8jl8dHAbJUMmLEoNxijXxcN6gM3Y9Q8EZJ
HM+CzENUn9QxRbxS4v70tqx1owvT20yY9JDbrcAdE0PuCO9VVm7LKBlQRPan1Ggt
vQ63b1gWHCMJ+iZFRD5yQp5BtfyY+J/EH8oBGR3brWt6QgW50j7a8BKsah8C8jXj
tTDq0Xz4ZOkVR2zUp4517PuW42uNLH2MfCJZ1kWP00IRzhv821RFktroIN5PYq3h
mPtJZ4XlMs3MuHcNeZcsB0IgEW0KA9K60DJB8fJGcCjzE077OMNBX/y8G5yUkfSy
NkoCPzFK7+ONljMKrZOW9I+MOmempUuEiUJQXiT/IzNly7CkfsHsV1N/xFg2nYK8
eA9Naae5ohnpGfaHutaG0cQr7tQR8XLCA0+52k3850LCiMMtu99QaVaVKq9CYG27
kktPERlX97hu6NYLjyvSihPRuzzS3vFWrFIf/84IIcBlAfhbjT1GIqJ2v/7PSh/y
0zWMD4qIW6wC5pwBipm1M7qlFgU5iKb/yBumvgLklbs7/yCDXat7dGf5WE8FiqUD
GZ/xXNiPFLE94r0dtur/Yx4ukQ5GMpQ/UX6jPm4aOPwumTCR9RikGkSTT5Ftvm2k
BfnMHP8mSk9lBhiJ12CN81yxlvG7QuOx/RXoGRzpv2WHwFddB/XHkTUACyGnbVlN
nvNU3j6x0+DCFo18eBIbwEtgP1crKzONwYh3gDwj8JjCg3UOCRXO2b4S0T6PFPsd
kJYj4/1khS9ot3tgTD3jDeN10QzNynlWAowMFJ8lg3/nL62/tqlQ9oz289RKQBwb
jrEyJq1TIsTodyyyoeW7omUH8vpI+rbva0qzWaifexRer68puwaZtX+ywoCfwi2f
Ki1SHSnT/YwGmkksytMa6PlH5Gy7+rRzibpzP4YEFWPY5KFcWq0Fs28jAFnrJmuM
EzlEMr7S6EjVXcjSnwPjqFucEshCqLSMxzZ1lS3wmtp+7mrUnWf0nqkpi9WeY7xu
z8Si7IvlkI8mALTnzMZi3qxlPORsDPKWOMfHfZcEmCKiv2/okeTUqDJ3g2kwDqK8
WSh/PV4i5MNSNuUnc2ZK/bbFQHgQIQm+JsI5OiNLCvi1w6oQWb861h2fSmcON7TE
n4RER5dNh2o/ZH8utqCiMqae6Z7k8UFbRsoRLe5q831sH+j831Rtbg9fzvNp0Jsp
UOVGT+nG2rzoD/8PwjfzK6fMQIvkyLsVRJVka95/YOzBLcyCcHhiNzavD8szsR+n
7fJVdfu2UPVwlKHQCIXCRv4ENZRoDycvHeLf6lti9MbBVIw8o5wPlN79bqOysGNB
DCEYfc3BTQJ+CbDDJazICaHdDduRqYbS7Ax1bXofCbQtp9wQXBd2LkJuY7NZz5o0
BPZUo3A5PiinANG6Mb1kp4N+i0UPBSjolTTVSSTPDiSLuUrkdKd2q9AR6wp4Dy1x
dlZsCMxHNwJcGWxk52ukrVDc0DaXwv5hOdHzpwSH1yVrOuP4RwSAhEAOypPQCLEw
b0VTAmZmU3eh3GA4RMo4aVEMNdwUyJvyoSVOjnyxPfBvxndbEsXnSaSN5OKKERS8
wLy+FUdPqNf/HPtkUQAU/VjDFcJgvgISRv/iogSFhsJf45OkXU5MLk8T85p7mbPP
5SYRJMKBJXq7Ec9szGTGfnhduoEmnwjTZ6nnG+gp6TWNNJmdK/p6vnRRg3DhXj1l
aj78iV3Ek+QR/Dd9rRsIzJo4aBxKgvQYdlIVuPOX7539u8GYccGUcU2zNFtjCWLl
5TGjWAaVdRmDLia5Jy8rD077qK1YZRg+DPdkO/qk5KMWdAi/bcU7FdzYFPOA7y7v
Nfd0TjkB6vFokTk4YSvo0LvqGLnT6G/LA6h2VkBND8J6H+GQR8UYWrrD7B/AL5B5
PWj//GiW6tAIc3SUnkxkhKOrYy5muBw6phj3IKZY0sq+q/knxgHp8jTbU0ZGPBaI
GMb7ljXjaxzWJ2Gi+Zdlr3m4VzGc4mLcZBb4WBzgUh8dWbrpOyYZHvUy7qX0RTWq
LRkBF9aGY555/T3+FX6ZGLS0kF8HVc8eda5JX8CgR0VVol6glRfN1XS6RD9vZTEm
F1k9L5sm4kic6v5U0EmHgpnxH/f437Le7ohVjc/n+xfV9TjQBS4VIG+AcsQvu9GF
vSubkWeg/gGxP+icctBXBJkEcnZF2DeDaDQuvOl2A4wPrd/7A2JKV1HLQa0Bn/fG
ciXQBPHrijcZNVmt6Y+En+dnjVkNfOmu74tuqEXr8t9UowNUOgKHEkisuTbCEj7j
U9Oq7585tN8mGdwrdnh0m3WnGnq/DMYAiiaIQjeTAQlwgSdm0deiph+4cQWa2gL5
Ppoc3JetMc9gjGkKCoAdO5v15oPBi432qPcx1sI983AybqC9+puH9ruKLe78y1mF
RR53p6qMVlawOvc2CAAC/9fLSTrtVfPC0/yQu5C9pdj0ldyTbwsx9UUkmCAOdTeE
LY2GvUkbFmdu11tE6bbpASRaW7W04+ZFLTJWJ+G5lIfs+SEXIpw9YysgmlCbOEDE
Vr9W7/iui+/2Uyzq0woE7//F6sSTqAlyJU1YU1cKYI/Cgci2x2zi1BicQX1wya7A
gtznZKuY/VaUJetB+7sO6VrOcMpSh8FSy4Vh6j5+L/1NCyp6+JsFXOIWW9CUBy8d
0mZ+Xu/+3Ddndj9uR3jWo1dGRIudEL+lzZrtJAplGQSi31n1kgMF90Zk80ONC9gK
FBC9yMoyC/ZaQXcxlpW9mq2thMgMUGxSgcNPI+PhZzBVjImxv6px1emVoe0ePpOk
MuoW5HRKAUeWMd9idoZJkKpMGG+YkE9OB+czyKw08tsbEO3U3+8uVriK3W4NAReF
zaTa9XuNRE6u6gZl2UqETsDgqUa7dvsK9Nb63zd57X0TrRBPhZaz0/DQUuVCnZed
5IAHZC5oBJHcPK91vTP4euMf7ihvosE6fitUSpvZRkkKJq4eTsG76Pk89Mu90rmy
z4ZZ63gZoXlkYW6VJpD8DUf7OVPND79AGjzAFvlGA9ktc+gGRiSvZOC1GE92X5Nn
oThn5Bh7Pcb93Nx58jgU/ULYmPWuZlXZ8gcgzL+84sEkPZw4LwUC0fz8n1/+54Jt
o3/ZKFEmYpnfyugMPpFwqwMqSHEzmW5AI21NBB6lNr9bmkUJOmf7f8ROTqIYNsvp
G/jDiJMdjJkS2RaZQVU1hw1FJVuiVVy/sMHY2EOufFrONa4kDVXWNQvhChN9F3B3
swEkTpkvCpAXVGGldmnRyDP69LcCnSjXPLnrq7WkSy5Lc8TCAmKePfoFTrhHKz/K
cUpKwrC9gWSrStGjIED5clbjvPym0VUJxNuJFPoAakhpURWINw+PoUKP7Uv1giiM
1fphqfWVA92b3ePnEdrjTDLA13KHMJnBwYRNnxAIEw/A3HqQWycQUIMfKxjmqsjJ
DtoxtCp4u9R5KbE4hDIDqi4ghdyk7JkxpMvyp9skJ7Gqjx++OkxkJOxG7tWmBXb+
e7slYj8iNHPGhMmRAyAFq2XIIRpN25XUAnYn3fHoAqpXXhB5DDqbcbWG3/0hB6xd
Ea7kdltN41C+z2pJ0NImCPFNbHjsoajYpwJoMoOCF0u09LJrEre5+0vgxz1KtPCK
ov8z68B2pQXhsIKzIADZGpSACMPqkMNsuh6qm5tVn7HsdHnAHVV+IVSEcyPQKpsA
0PAX4Y+PotJYWE8MKqgEOWsUGu2bfqnFDsdwoUhDQHG7EnGJtQjQF2MwL9RyDCYl
iyWSXyhiduTWxYYfvXLoYIjh7BroWz3hTBvemQAOM7wVGKkFkLDdU0LJk9f0xsAl
Yei23ks8LyVz//MzdDoVb1K6EYu37k/kOAD3pejyAPgpfVSA0GSptS7E3o+UhcFo
RHNi7N1QqcmkFPHaNK/mgBW73nZfRDrlBko+wROZ/KuSCa/IUN2z1+mjkmjEBjwW
HD7CVANjxGkRUI8AjeHHKJFXwKGtx3rG4lBWA8LihcT0kL9bIWVRhRqs4HE2ZfVF
09H4JATR/AO5oecG9TM94u7NlPvIXWoELDAssIYoLZAnpUfWwGvvmgYeL1i66gT3
SR/yrdTkXZAec1vRLttDAuOesBS14CB+ejCYPfbfvFCtU334zECdaccG6he9X/jb
idM2u47SnvQIsBlzvsWUBwCCWD8vSO6UtSDQNaB8YGHgMLSgodeCzQbPDeSvgVVm
t687Kv+T5R21+ulwuUYhg1o1nlTo//TrhEycrmAh8CzCS9nwg8svd9KbUD1D2aoX
HY/50bu7jowP4OqUaHonNoIIRoYvxWJ9NnPoCO2iN44q4WbATxFpVx1lUnPpMz75
l21WOl5ZWvWCfQSuR3UmilEJUxUCobqUXKylPVmYSF2U1z3kbVhHJS15XT2Ge4Gl
Z6YRB9kOuQ2q0sFtiE6iERptP32fzlmsOHRS2gYnOp5T1h/9GZN78WZqMG5HQPj+
DXB2ULWy0nNGIRdbYzEZHTKNe016uQrFCX9LqpALtCJcY2n1xbRINmNUtpBDtOQb
4iPjp8u+9zuJoZDWWa7nd74YKktyhRdZaGk8pYBLv8o59lDpAYl2of5IkCzNBnXe
vVOZUMwYWzFNNFUohSlGNnWEcpRb7JmK28BFVJcPwICBZZkT3Gcd6q7A/MK83vOJ
S1WyB+VHsqJnM/VHsW8a2fTyQQwC9mAKWtE2iBrD2FH6H1KojYtFeJ/zEHvFi8/c
pKSesWPycKz/EV1ykTxh6xk3z7rxjAbyDsMa9JQ/Km0ijS6st0CD2VSkqKlCcE+H
j13V39O9046SUtBcTN1MAqZo+Zi88o46kgk4iUxAHvjdYm2Qa2V7F0kt/EY0CM/A
xC5MmALX2re/BEOJ5TdtCJ3C4EpnURTwSunQxALlwALl7qiEmKZ6fyJYX2dt5Su1
dw49hFJ8zHmVFWxGZpc8H3Jp2Rl8Xazw20H8TpZfBb2uvMe+UdmVy90qZmx8rEQo
tMksCKK5hjRUt57N7+2AQJo8sBmkyYXaPl5QAGWbKqyFUL2Drai5+GjvFuISscwH
2JiSTEi+9a1lLZ71n+iyHLStwJuv+ubHw/UVQUJo1o/z8pyrCLsBfyRaduQHmuo5
4n3/sDcVBhU9OyPJlzM3/5H3dsEcRwCgRrbyK36iluFyrSLAFDODlbWlqEetFAMs
aWXdm+h8stWxd9+Ffo0lpK8INEE0OjKkhaa8w94kRWqwFxyQAyj+CPZsNkLZNGeT
aAZzuCMCJhocVvFtZ7EXs21q+ru6a6g1FaPdPS5Qvph0WrH6C6y5ndfiXF+18lu7
EOZbNjy7KTjII3SfB3ExPLDy76JqDkclDZjDbwOtrbEEL12gXs0BAQNWJRqFu388
wiEP7drndFiM67ur6Tg8VcnSbEUaeBNlrBIjHSdfbtphIwC4e487RSbnAPyo3TfZ
gqYDd49bUMOCZRqzypDbGms6t82iZPj0HKkP3j8wQs2mizZkNqvgQBGKZ3lC48Sr
m37yZqh3FtInpiv3E6WdzeUx+FCt8587P7uex6fAd8ZlQfg5mnacg4sp4KG/44Dx
8LqigGOg31YibThgV9YUpWIWRlJc6TC3k3iNXHXtsWDo0VnRq0jG/SDL9aN3RVpx
/rX6OyhmE8X/cPkcj7LhAVomDY1YarsP4KXw3mdWNpn1T1vSDa18zJYuacoqMkPH
yWNeOJi9OjNwAdA3wl/SGa1yw2mumR3cP+UoE13EpolRk+eV9IiCPY7HHjmWytvD
IM7OCngyomYxFXfb3BWBDTlgeVShQSd0rtpe0u7zzWQo9rNBahk4zA3aHdGE0R0g
IzNxsGCXwnuR5tQ3GZxpa9nIGL5WyC9B49H88+3T7FQKzV+EZVFyADm+ZbtzgG3Q
lohD9lrmIiFHA0cPuboSybl39yedSsYIFeGf+qvZbel6ZamUrGkE0AKIgXtJ/in6
IpxcCpvR0YjJXnafaH9ctyN/yGeiadETEBT1O68xEVS9QutrD6jCb/qxLwHILRUZ
Rh7BzmiaPETPBK6IFyOVAOTgOuZceJjBilsk6rUvr1aYDul8EPixRehLCJlWOEfa
oKYTAd8IirU1xF272+OdGcScfZSAs2egks9nXHcxOjlU+AErn6fHucaO9M0F74K7
SyVog9jaDgjY8XM91aEIEog5N6YbI0Yx1jyxx0fhfDStO30DpMrnLroKMVw9/tGj
K7LjFQ9WQDV8BvocXG2pJEFaUxxTVuwhH34KMcjBO9cUA7p7fFYHW4q6ExfNjZQN
9S1nhXK4s2DJlgCyoBJudPlA5Cs3aSbx8Y19Cc/Z424QFjjxIVAtdk4HOXxQjNPd
/j6Fnzr/0zp5LwfWjQO4hMT6eBo2PH0qnWJO2bqCFUGRvN5/5VrWzhGyvrYekoGp
yLvwvpr8QVzciQv5pp+DvDY7+HUAMOIRnBIIX8ojmfQH+7RS1E4aMZZ7IH+lXgck
CENQ24Fm1WrnWJaSaw8faBk4D7wbKA9vEBQPoEqUNT4Xwm1U67/7JapNBB8s3JTL
bn1DXoKffBHwTh5iSjkEG5otWKY7wqTPuAl84yp3I3oGw/ty0ln/d9vEQ7X/GGkt
wHSWRMLdfLVpiQtVavBYEU2GIrJ7zrjEQJzkhLZHPgjYrJ80SxEZORO4bH4BA1wq
D/SWIbk2HjMS3Z+Cr6nqyyKjD0lERqPGdbXvlC2giIYKsdscYETefJjtuRm2XP+M
NjHLXsX1DsjY7SHQIHFoyaYvdsJlyu9qzki1FDu3MJPZSXrHY/U7ptmBy8AXiFC2
HEnSN7PRBQRxEEliXCxAr2mLWZGrxOaovlcTX6cewZlhA2AB0LyohGqdqS7bMrl5
9ypKuhnxIbOQPjRsbmUMOvFXEdrupdDbJ/FWcutGWI+qnRFmDisDmA3v8FVQhe2G
XyNfLIlk1lh1UEkfesiAxAZo7PwNl1d4Y8s7ORJTEN9092m+IK2BFwB/z8M/s8dP
2YQRN9fluSglnhtW4N+ySsyWyWFiSuk0po2khrSb8R1GpWgP8I6Fin8k6b/1HrVf
TOQrBr5OAi5r1dNMbppHoe+XDRYg3A0KcyKAo2tF9NpGq31LCbYavZWJ0exC6NHY
qzisJvCQ9NMj3megMIp1WdmGvbhqtLB0YWhqdHJqdDvHFOe7MyZmSJkkVS0qx7Dn
I7Ao0qVErfkPGOSu3yXJ0U9U0zKSVOc7ppywtHLmWIUHg52Wp7zFe7T6JpuffAjq
sywi33qw4Gv80qwAoegnsqz46eqKLLMfLC4SNSOawPt26yTeGLYUq4Wf+5h5oYav
kUOk2heRkvll3Pw+Cy5r0fuLjg909yU+66TzZOoQjd+f8Ziy115fJAdp0G0cb4lV
dBj8yHtV+4sOXOZsHW5IkNt5jShXwkXJ+tc80N9DbcopyOvKVvQbhC+lVGA0h4Pp
M/BcmYvTGgjTUKMqXetwjsr+77R4Qh2eT0dT6T4p7cCSWPPD2yRUJAC/whx8NNgT
0a1HTDDDkfovibyAHg4BayWGRtcuSa7vSURZKd35gMPhPx9sV5oAgwoAr0Uz+1BV
Kty6HOA800BmbJNTV6he0Zs2+OHwpzo7bOxzSeniP9L8vJpCwVgZVN97ZnXzHO+M
Xf+RtostxgXFSCpu1XxWhg2pOn0SvgJCb5KJJ4RKnKEQJUYZqCkZ6kmZ1WoTSiqp
XeXYmSgmQi2bIzI/495W9ynNlERSuf88uWI37mdhGkVW3stdGE8bYBN5x0+Ypc/I
hU1Ssh3h7k40yGN/VYSF32ENtdQiFJBjZPZK2x+0JyMhpK49GVbQ9dT61OBGA/nV
EedevkliQGOvPf27T6Dvl+pWxMUSfyE1Rp3cdFKCAArJdV41MPjKEvhLyUZnenQP
TnfpLQDR3XwUDco/aWA6XAeU20Qzi97i6chWKwND6K0y5MF19yj9Gbpx4pSU6mO6
9eMs4qxzRpLtHqu6xi0EGzkmF/85vadAulzrHiEmvNNXJs0+jHLDATF4J/gFkao9
IzJPyK+2UFRFn0Yv/uZ2b1PBRMK+gLVx69j6Asafh1wW4YULt6KBjwcR/9AImDy6
jEdt04xXS1JI21pSWE7V/6AjY4lB4nMi8gHrXQlzhMDbd57v60+lZGw+Q9qwdixh
Z8d4QmeiCRuE5++M8FHuhQQxgdO63FdwYR59jSLUZ4dWnLnzNxoOYB4MdIg6X+cX
KXprzxWjzoi1iH25+Rxf6IosPyGa/bMRdFX2Nn6XNdaS9/pl2epxNd7i/9P6DIVU
bO7/QHqD2ZQOVi1C3NG1lofhGW+ohHKXrGwYs/Jbb3uQh2fFiI7K+0hohnZt5JRD
HXHR6YJxUx0G/t650HLyOjU/sSnFkiOvUV4ULS0V1Q136b+WSQ7DNImhdTXNmv9N
lDJTOjvqWoGwSBi86sWjuYRogC+YrjmtCmuJkJdryoGezlvfClouhIWN4ZwUMoFr
nPwdfghC2izCe7Zvo8SvK09HT9Givxj1z3FGGyG1Prod2BBa28qqCiL6j8NY1h3R
gxR+BpSb67KteaEiTlYk229K5AJ25E/iHR4mwROIZ4+Fyin6JTc8T9vAIRX6HjUZ
dNptogPqoRC/pGRyoJKYkH40cRLObyINZrsF05y4H2zDKS0XpNHjNJUIxxO3kIx9
EgQMz18BRIcOu5q3SRMQ2B4/Kv4Be55POf35g/eHvsugVJMqyirpa4ThP0oydzrl
biLuHXpWuBu0BXRyQr9q6sLpebNIK4mUn5oi1l/ERWcFd5wmH6U1LIRdsq7J2fZI
ifAiYY2r3ojHEqROekW+Ksy008lk+HSD5rsCAfcwVwIBx8txw376qSjDaYNszkR4
pJBcDVnHEQo33uuT47Vz7CbMpjaxMTFekR06O3lzKobpBOx6yIMKNyuF+j8vxKK/
vKd6IicTIt28gL7kcJZII/HoqIKLPkY+jgoEHmWLC0PAf98AhlWwRZvm5RcSCZPz
fuyZS8kYmTzvd0di9DYppx2o7JjN7txnqvpE8M9PQbWKOkJP4n0cPU52g5pK7nA/
J5imdYm6g/qVF5DbKlmpUeenEgsY8G2gCJh4lJse4frdBAXmMD66OswzwbalG90r
4U+h0SARyb1E0TWjpo/WyeXy/Xl0T/dxbZs1JdvHd9F48VqQ+Fq46PETFQDy8Pvt
3mZvuyqLRg6sSdvA3ZCiApmUMgt0BWbUkPEQIAuQU4prnPeMrr7BFeuNf9+VDXM1
/UDY8bSYjeLLwKZsNEc/K4+ZvkZff0hpy7L3gIy/mFNKOnw86WSqthnQZ/QUxDx9
Evn71Cz7GrJ6ENrxIXOfywnJ+WMHl8ManLY3HqJoJ8by87aNz2LWDp3QYJGD6HqM
FHpLlyyfW6CkrVRvOt/DnqOTeQrmCeHUC1g6sGi/xVqHPVoQog8igugDi682G4bx
Vb4IhG+v0Pi48yvJDPntNry8cyStwKl4jW/wHZ1IYGpGutYHGlmoFZR7jHiiKxAY
2jXBXmKsjJoVHA67HbY46GfKhT/ieEwasw4CJrsG8yaDAmrM5jLgyKLdaCXxWZsU
Lk3u0xuYuby4f4tfofJvtzDddgU9N9Rou1M8EpZmI8CZrGaHL9UoYI9T9+pNlYd3
M0vnZaWZ2GUqhx9zblDFQiyztbQKJGRgKlkLlGzvIZ2oPo1D/7/1BeFZN/dXbL/K
7UoyaROW/x5Fac1FtBpNscYuv41yfLIm0+u+pTidV+E3Pm52bwHGqgvFijmsKHlj
7xn+V1zwKV8o1wH2ROQuBXz4l6IMGuitiHG9cpAbIVi52US84ojmXxoDehponjlw
YmOnKQlNOtrrPzT8q1jGiMq8pTR+LJSuvm19oZYNcbYvL50o+cxpLE5fN6huwgEV
aPAMPv/b8KpWh/xk4qi1CYs0Em1Tlr7ilyFlPfbTs9/Gx5ZQkjxuBkfIUMCIFDLA
Da333eS8y1Zz+xCPMElRqPvKW9FFatzDh3meIQ80TpqyuhLxR3vjIkZxjWmG8ww5
nFynyTjVPxiHXfAR+7DKRs4vPzF7lPckeuG5iycFtXMyqC6nbkrduTo3GCYBfWpd
oOjFhUiOdFM+vnzFQw2UJdFamBsun55Ilzb0auwMaF1t7bSpwZ3aYvxcEu1XiWEW
hjmyN+6mPs/lt9Ii39P88rAPK335zXBPPhzRxrrkkqynq789FMssELjDGoaHgCH5
B8q7m/JPiLA2iQisPAMlG9QAYGYky8+HJYqlYnCpL+RFlIDUnbOWIuqp+HD+vkLe
hIQ9wnEZ8TDEIxH0wGrfdwh9otdOA4+Ysj47QnOXaAdPqIaUyy2OoLJ2ME0ktaSE
CpASGsv2I1/fmTGLVS/yHcYJ+ibhfVXn7Aiqv28j64vN4E73VcGhXLv8fIfZTE9s
pLcx51Yim7MhpqNgvg2seKMCeN8WsLRTjtjI0Csa0XIJxzq3kB88+HxhY39q/gxm
JwPQjObcawKr+BUOXQ3wtFsyAiFPLexuY8ABZIvdMDLHl3F7WG3idrq2XEtqdyN7
IivgxLU7WHX4ipLTZQqniLaF2p03GrXi5pKzc+HIKpYywiB+sdyz/ZTBftSqF/Js
m2/pIT4jxdna/hx2NLvvdFFNQWquBKd4wZv3l6t4dcgv76zEdE/WMhDZxEFWqzZZ
8+Wm779R1oMkMyFFlo1OEvyE1Q3yXKCTH6JwZjLTm6HuGvOF0yVhrzWbsSJ9cpK6
SA5iDDgyTwqfF3Catw0gdcV7VertwIknGY9IdT4eoQkHBqxrRfDjgcMrPBjumQqe
ZQUH6MeMMdL4G63U1XE0eDR6RBPzAflK8C2ZL97y+0X8ZHrL3XQpLHcY5mCIbWlf
Zj4+Gef5B3yvWP3rW9WDiH6ozVUbLAGBw1f3gDFK1REVV6urc21miQZsB0uvWtqO
t8Sb6wR1MLmRlklWbvjIE1kxl5VVxNLHit7ZZS55xRKj/DK3S/H4RcMuOxBVk/91
CH78tO8S4vRT3OBVWf9p99dpgsqwRrKGZhCsRwKp71P+a7kxW4Elx6ZJm7Y440x9
PLOrp+juYaG2uxbSHNvX6zgwKB+RTXniD0/fvqb3f955zsk83MPFdBEH/g9yc4BF
mXtg0+n9PhAA9DYc6adcM0UoUouHv8RrJWd0TvTzQnOPYzOpaSLVYAZF46mDRfjN
gm2Mfuc4uRikLjTeMxcG6+JT9zIJvRBF3yuU2tE0BOsm+JjFijtBncs+NDmzu5O0
IDVir/W5eSm7DXdT305y5UM6DiqPhUwOn4JwFb2ZMb57vYa+p/3zcji3QmBvyjb4
P7ugiK+TiAcj8pqYCc34+M1e3SEJJYR5XZ5jV7fFdMPNZ1iKvPNsmi8XHCy91NW3
TlS+8Rb9781/qNl2h48o90FB9IAUXNdS4FwIf+6HUjQut8cpAaC5nWflJQgYdLnG
Ln+CGqiZcwAktJBrZ6GVWonZsSPwws8W64GuCzDvppgvyalEygwCVVT/hzXRxwWr
v3ajhHiOUz0LqhvL1WJE0OMDC+kJU7WJl3hVh66LArlniwpDHIYF7dcLnEuGySRo
9Ninh7HBiDr/kQvD/DkeUF45g8U480Zqu6+UHU1g4H3rlOQRfQu7DFpc8GzvpR6N
It7xO+RYcupaBbB6pJAFVJ5S1hyqjCcfHiqyRCnBUyK1GpfK2Ij7K2p0dpAeV5vV
iWIpg4nBjrVp3+y4TVt/E2U6MmXRt4QbtVU4kqccyC7/aCTYxwtXSxp0QG4EL5kr
aBumRJ2x6rpLWPUZJ9nNyHUKeiHbbZnMBBueOUyvTJcTv0vMxf+7okmdmKMekBcp
WM1PveN0fY3ManjV3ihHGiTVG5K6DcMAZt3+yRioIu35l3o4pKrWgihy1opBHiXL
AlVw0p+3TJdq143xj5pLeKGkH8aBpoQFLIYqhsiaIhX90AJLhctAYsRUAckEpJja
EvZnZFldcJ2e/N2bT1Tlq65+0bVH7KuY11ikqCjfyNYiIXaeoLY4zW9RGRm7OXkn
hJToLcPoF72hP+Oed88/SuLUEoQn2BWETeD8b4bvXGjJGq/BeLiOusDX0qFL7mD2
CaEwlwxPDC17/OBmXlpu/8a9Wlq1sWLZiumyep37vrzST6RIVGmKDxgSCYQOGTsj
SzOgUK7z55qUfMHuGikvnoQo816mZmchOTl+Rpm19nBeU4BzSBCkuSRljNHR8IEP
sxCqt/eKs1ok02QssLssu3I1ixsgp7xysmHXf0cEkLKOkePtyX3UlLXrMzpLysOo
KjBIoG4p+GK8MnFmtTIhBBaBNjOs3jj7U2TeDlkP3eV2h10ucEzQsp6y8iCwYV2a
GUgBMgtCa5TiHxAXkMgzbybdjGUGWbAPCDqx7sdTWGGYsu9vNVKXooS6Kkh179na
bbDsYTD9dsMqtKHOhfXxbERk8reIHXAzSCvlRfSTNP0xxB9hAxLfN2VGkNNwAyOm
WWlj2EWOwKzjc2VAuJFB722XbC4jOH1vXNHuhstbWQ+QdY1jNcxAUvUiPQFJ0lSo
9mJPzDoFX2KOnRvcebm0aUIBzggN32E5K8dAFIDpiSPufBXHmkRL7fdLmMe+ii+B
DsvpbporOHOgQNXfp4Q+3sVUoLs40D4t1+FYaEVdqlHy9lCW7/srhO2NB4HLG7QM
im/kaqv9HxRH96cFVET98FBrgfpPE7/X/51gdJ+bdoaNxv3zexsj3xf0rIwo+4Wc
5vCViNF4IU+UqrPal++PDSHiaTh2vQbfV6UcTsds7XM3ChlqlUJjmwdk0ZTxWkS5
xI6VXcb/n0druaT54At84Zn2pn3TpugytdnoyvX0iRVzlTtDfQrFpbxDgXhkPtWh
CJPyWZeimoMAEXQm569h/BUzs3FExpPXZ0azush5VrBS1xbQqnEOkrwfM7IRSAGo
5i/1ttxkawv2XDWXDPY0j+E4L++cVhIbb3md/643RBofo1lRKnMohygVw8h0/tm9
jWL+Rj88ed+oxq7FkhqJls0peGdz3yid0vgMORXarqqN6MtSmAR+BSO9rIzsxYdm
ohg6anm/qV9qbiAoCW9CE6HsYNO51jSjhTEHS2g1ycrcTapL619+Bl1LqMenkfYN
81E6hLOvkL21EOhQ8h9OJvNITOTV3A9ibkTiFrnZsE9N0wjeIK2etTCairS4ZOkp
eSWiAQueT6ABko1JNEqmSLXTbD4Xm7ajwkFRcwsX3fW4HuJUN+8jTj8KvC1Ub9WQ
UUXqNxLPi8x4bAiXgsz0D2lLhWkSlk5wBfROOuwAArsUcxZZbwVqX0WmKJCmPFXK
mvdzOlVNoFyW1H2ZNBD+BKKt5k3ttHewudB5Hui41sp3QRT7Py5K1+SLTWcr38yq
42o0Khohd41OmbdDkbsc6npBhteFP0r0rRPVL9UjiPNsquSTTVdgdJrDC574nzXv
xzdArTEQOzj6hxRwpz4Jljb/u18KUL2m3pYHEmuw4Y7/eMyVtd8ger+Lqg107uAk
CHgd3jbJ7nWTXMAFv2gCtrQ8bVPxiNjGcuzefgcHj0x0fWcf7EogXokszLIpAiSg
uBxymd4dPENbNOO90xENuAl0bWSgVeKbgjKFzK7iUoMpZkdM2kpDXXZtbtLMJk1j
An22ncxUUg9z0rrp0WlHnpTa5S2amJVfb2l+8AhV9Vp6h2b1exY8aeVDA8izJ/CZ
HJjqtWCdm+yfiN15taIPOYg9jbjEDfleKfp7YNgnMN3lqKXXfC6fr+fnhH28m+5T
y86UWspJJigfEgcpRWJ0cVniF7QrzYJmAIqmk+U624qgqzFqcb02DwUwBvfNjOlm
ZN892DI23VRQCgU2QQziw2DgHirLwLuBAgvTH8/iC8UBw5ZSupdplGsbtLCPceGY
M3Ig/zfGT2A1rC1R9O7iKLbJ8p0ToBTzYTZ5TrVnxngfyhX7HwOmF1p0sao5LXjE
/F73Vrg0dxEBME4rxSuBEsZaVD5vdXNZ5kEVbNp+i5RZKe6CTsRyj4hOsfMImUKh
cDrzdLxv0R3oI6NohTTe8eEmP69pcaGvyRrOgyttmawLlIqMQpHDsNxwMyj/ALKA
IlBABWGLm3oN2igB/JR6PzsECu4ddSdjS1DUCYYtiIzcQeN+Vp+autB5/32TJni1
yPNma9QkdXnAHrNqLMQ7bNQiaCOT+W24697aSvOOluv2IpwFHO5h35lgK3e9Ve56
1r65dBiwvc0RRTtYBXQXUWEQdhXER3lnRE/e5AOV/Clz5rKKV6UQyPxucqms9BMH
JPT5ZIbIvm0LpWX94YzY437857gh+25xUCiMkCnF+zvCE3ZnWEC5/TGx8b5M77qf
nJycExCj7bvOu+SCol/OoNT9W7gfmQ/li9XWNun7kJEd8EpNCZgvm2G0UTKm7aRk
xy/e1CDG54NXASXFnByTuyCjkpkA9B/Q7yyfkDEostqDKHVl8bW3ygj56o4Jq0MN
OmAPFLwqZTmzou2gEWqpgm7SsRaY00wkbLIzr/kJYcy7jZdxfftSMdnGLAhblGNT
WHyZv9G1V/UHm4h7qFVwuAq5VqLPsmCV8WPXnChADvueudB0C9s/XtUWF6meh8kp
qYEC2tq0JKei5oY/sr1I3aHYrn75haeYuz3bcCYo34sD6LDAvCnnUkvSv9ONFXAk
AfgZhQGkbA2VWUR7LIQNEFR/ZGBE2EB1wz5Lj12sdpTAq3AaWNg0U3vc/U6sdB2H
ULRkHoM49cqzdB5bDweEQ0JYnzFhtxXRLBXGcwxWzejj/UxNfSkJJNvkHsvCk3T1
GNZ20ICX4suILxLTsCk+YCh4OsPJPXupIHBUqGvxyZ3L8WSHmGtcQNGlUCX2qgUP
UMxFYRV8tDx16haf3z6aD+kUzu4q2PaUQz2GPxIoyFI/XYCnEzNB3KIrz+ArdGtD
4rZx8snjRUud6gkpIuMb4A9JuXX7BhPWTce4j6quS7gi/9eIMVe78fSHqz8ZBGUB
8MCbD3vsxkEfsrQoUlSlGPzU52MnVl2bV2CgW0CrLXO1rp+nFoORw3DOQRZqAl4+
Dy85v9ywsf1oBl592152IyTl1/9RwWF4Kn6dEWkjiHFGxi1ZxicHX6w2mWn/DysK
GhCCOroyTPvgpA2i1uSNQPW3oINMR1Rj/ae/XcDjRoWpKuJQy34UFXU6UTQSmhyy
pbepUWI7uimpz6Vaa6kLaBrS25ENPqA6xP9QpKRvhqS9WsXHOe7DMNKYlp9MXDP1
fMLo73cA3oBQO4YbM7djk+pz6Lrdvwhhq0eklr4N6LoZRLzQ6p6Ht9Q0rlE8XKZ2
eY+2ibCVv22h6qP6xhx1iHQj4c8NiAgldoG+UDZcuPLXEYQcmmceBcdnC5LOoDQ3
5jMc9l0JirV8TZMek4ZFgWsWD8r2TaQ6kIHYZ8/2TlorUnqqjIkK7kOv2pgUqL0t
wtgl5EDCb4nDyLUj13qD0GpcNQ0PpAG3GTZVmWcFDeQRiOr47b+VToKqdU4v65ai
9F60SY6kIVya6Yst8vuA6jJALZx8J7xIsC8EvXzuxof8GSUCRnrBZU2HnvYiuyvP
++4JEmN2+PcFrLb+mKpYSdUctOYk4H/QHOF2ysNjDZirgE9KuvmICBHcl9VST2Eh
INb+Kj/9nESmzDTfmS9XSIMIGmklBjqIG9tMrWDU1bY2wqlwiskXQ8Lv5KElbv13
KntP2vfOCd56PK3fkfOuQItKw5RkkrVeJbW8Sq4brIJlro0tp2VoFMJBZlu28E4k
SsGFGYpGCYP0YVC/CW8NIydDImk/lX8zgWMHwB/UtY3rApRU/p9c3uNkSnP+SFTH
0q3JLHnFlkZUh4/15dDp3shSiVz+xm9EdA6YlqyUASwCEMlqG9gStS3IkogvTSbU
0w4u0PNH5QHEgZaZp6JvDv/pPsOErncp6RgyAIT1RHt2GJVS42I3niEWcrNmX/3K
i+qhcUv/MBVXJlPgAtZKK7T9ASeRBvZVmK9EDdHTHvLvIrD02iRUF6JJPsZje52b
EJRLQsTVtO1FVF9513oRfNurGTSDQsrBf3krgpB86pV5G414BkRYDZLhBeGCCG+i
AM12ACZt3CMn96gD8I4Cr9+qQd991atFJH0rnBnKHiGieMHC5qtWVgeZpoT9n7ye
9N7JdF9OvG3Khjx4IUuLk0XIbzDoQU6nrvzuzqUvfVvfPRG5+PD21ID/lQyG9OhG
RdkzW9bBE8PUlyXPfsyBUU/rsNYDldLjneuh+cc9hoN/RbtgIBBaZTxf891J/RSM
UaM8P3XLJyA8zdRr+SFhXbJBTi5xmpSwl1KvbUk4rELC+f04yd5ZWOpPoRErJoOb
LUpPXv0p3ZIFz8+M7JSj78VfbDQoiDydm/q+SpHDgzn56eVe8HLbHrDJ7anrdX+x
6dscsGIsRkCiEmXrKFZzLvJtkEjC9oT7EwmRXuxSXWSaSsWpRuoDdgXDq9auSIWR
AvDyRPQDQ5FQZpwuhryWbVvUwYHM/vlPHWXbd8I7mtta2wIf3cUmOEUD9mqMrOnv
DRZTMbbQgVbrQUzErqGk0TtwhExHAtbojLc+7piiT2Ykz/GWRoTLAXGDYqGThpg9
M7sL5hU1jvo8gs/nq+X4zVkvcvB05uZHUPmfsN95Lrt/FxCCCRHB9dJBqabKrfj7
w140bG2cP1fsPmiquTcjjn9CRY+0FA5+qkNr2EIqz7tMLtd261F2K47etz8uspW5
7VdJyW04Q1ihwDZQunY3wyzTZkT5Fh+U4matthapXTZWGbyZsvLZkEXJ0AxgzLLj
Na3XSuQKsXMiFa/CMrvGJ29p+QP8h4/kLD7hvPDVr8UChbFlQFugRU9FysP0gC6U
dWbFHmHCKPOS+f94HAwfEQpXTCn2Hxh9ZyO0GrCfFcWuzf7XA8FvPG5hpf8ekkiG
u1VzE5eHzJ5fZzwHemg5BoYVnB7UNz67uOCCqHS3NqodrRZVRCroLHfOat9ZNuo0
CQyUpEv3yFZK6vDZLzdTuOneQRsJlH49RWegM6YEWZlzYQi8K2Hvs66d2rXxMa++
GrtQINbEZlkpDJwoi9tiwbLUCsmfNRydj9sIP9DM9mXrw2+3Ehe6HGf/J4tPTpaJ
ibIVOrvfcMZwHk6/Oyb0X0uAAwJDjr07h2l4E42m+MHNnHwzcPhYlb6AJI2r6o8w
IqO/mhL6XZ5vwQP0U9CG+XGLYazDJX3bshJYPBIzun1Tw8K/Z+H4aZ354gZBlLlh
HRfxAqeYMrimRkYioPncKjXqNyH/1Q/Cd5GBKLGcL4taFnL3xREddU3gwan2dIY1
vXMK4t9/lvsvLJinN2GFC0E+FJ55AloA6yAZyV+j3YdTPUcdphsTNqHHq/GgHmSD
69HwGROIEXevbQJfqWRh5zhOWJ291cZm4vBbV67X46wFyiqBYhAmZsTGdqPnBXjl
t5TID7SEiD9d5n3FkNhc/JYnqOSm15iGTogT4ZFaJTZOzAXhy0I8pUMVyhsjV41D
g9ZPkZsLKXOvQZYENkdMjxv4iVvnDQky27Cm3bL/2BdrzuVJhfGT5UJXofM2HRCh
oOC+uk8zl/spGgsORhKvZokLyvfHLFFSPJxhFn386jPjnlvgxI2gHCEfzgpdkpH6
vDLqab3iOH/hE7q7nPx4Zg/Pgq5tWOZqOTiDOjfCMffxGcs4C4+5a5jRxYPto2Ey
l/d/rGngbd2tpm3UU0EDm3l+MplV6XhRXiTXrIK15jihh0b9XRrsek1NNFFXDUqV
KL6svOHnkJ4dvwKnggGLeNovhjHkIvYTjdpenJ6lpHMkdueiryUcMkth1Sc0XE+w
R9wxUnC8cmyT8DCyRDkkpstT+epL2D+F+vdgIMlX7TYVtRK3Q4MlYmsTmOsS5rHM
IwCamVyMxdbvVqRw20hg8Bqlqx7QuXYCUC3Na/mL4dtLAKFfFpIdUCR4NKlEfnp2
hrcDdx04ZZoQA5ghHNDcG4RTEVP6Kf07MyssnqeYBRRG+MHzuNlj31GYYrXdGYUz
lCFejbGfGYVk3+zR5aDYvg9Aw0RVywUqsvhljqVv+3mxcQDQ6X3WNKn+wyUzT2h1
FLaLA5WuIsj1ud1tEQ8pmLSEkCe+XfFu5+9gg+roXT+O7ivGH0Gsz/Jg3YjZQNEV
nj97vdvylbggbndJBcHU1wg43LjcBABQjdKOi12dTLpLEuFv+SfCVk4zHYw7bs99
SvEWWH+ccRS5Phtj4DSyhe+1QSm/hquYBvYKh+eU5p0UqTrtZ5TGF62tY2EFRpFf
gzCX0ExlE8fsEj3Siil41ZohPZ5qrx4wQ+fsdC9nm9ocpz5vJT6KnG5CvSoj9pyg
m9r746qmaAuW8hyCmREwSLM8g04CCQgpD61lAC8rFQDWuyyL3rq0PFQU+8BRXs6W
uU4TCVCwdo/UAwAHlkClYh7MKxs2uA4nzKypcaCjrnQXsktsoekUHhaFjJpiZF8+
w/pzUepA7RbI2BYcD8VLR+8wum1u9OeZ9vda28H1vdck1i36AB3H/9eMsB4M+2hf
fQ1CA3eBg+0KLJniBMxeFdc76wIHfI+QVdT/rwH9e7M9MDz2/BxeP1jo/H7cfHzV
jQfzuhRMOO3q3Fv6/8gHvEIEtp8VEqM3louS110vEbLLuCn7WA/DmsiYHf075bXi
ILhkiRQdYa9jHvvZKjy+1TMgJ8NoSFzS2GO2z4O7UQkd2L/x2S8L2BrOEsJrjgiL
3gAgqpSI0jUGGGSNUZmvvbejsMwx5ueQFmKw9oUjUSiWmISXwrZUbAN0+63RP/i1
pJSMlWWt0pGOa7aScBZOKs6wZ1GxiYJTmoHsh+Su9Yz1Y835ObzY5U3l8xjT34jO
QstGIcB1RO3NlNTS6Dn8HhIkBjCG22z5R3fzoBn8ef6AxUqnN5gvy1N+rYuDZBGh
I0++aYn+rN48T0d6pbbn1zAmP1rsLCuuZ89MdkDMubzC3zId/8MQVwLYuI+2T3KD
krQhqV2yqBrUvNh9j/t8HMCPsGADPJcx7uKLv3bDxcW0KfCjSOmN/V5lowWX9ZfU
sdauZ6rcseMUXxwMPD9f9aqB3MoPIBrA538QqlNJaIpiYaw4bhZD93HTeRavEiS3
cbJ7DWoE16ujnkv3nOYDapxhQiBLv6v8oCLpPsHGB+LNNG+LnNNlsScOe1T65xjv
KeVPpHCNUOmKeJba3GLkYHuVsK0BytDQEQbm82Ncr5sSh7bB0mWQwHHkhui/GrRj
eKK61cWZEdkhVZ5Z7bp2DSoab8rAkW7wXnUuZoUDb5IfM5CPvKp1IcQwOOF5ScKr
EJAzsjUtkD2Wov+mTExs3FCE7Gs6W8brxXBcbwoHCA3BAEPM0vi8r/Pu2fnkpDo0
Ytep3z7CtG1m9GkZnlAORe8/Upz1KD0gMq4aJGKOi+yf/M05Y5VHfkkt1xMQB1f8
X0ICZffUP1ru0HjWmyWc0Hx/njRv/6JkjK59/X6RhpV33Up9FAKeJoOm7iZHlRZ8
z7Rh46/O5QiS/eva2ae5VEWGRA7vWQvD5VLiKF7vDrVKKySBb55154FxOY2TJGzs
/Cq4/OEzFzgFUzgYGqRqVRxab09h070gmEVBChSIxu7GrWsVgdwXeRB/GLYUeY4A
+97A9l9vNGgDWgKArmxHUeRTMpgI/2CLVCG18iul4ozi6cq6EjtnSgBwmgrSpR4O
T6o69S1pwLppAm9XzNlJHI/zbt/L7ezqLEeIGv1zcXs9CsiCESvn1BXE97Z/PWEB
i3xA5hZlRLSvM3TIUhv6knfd3ZGidB26VDSSCnyF6wUF6tNyFdtfh1Whkq1MUnnk
8fEcx8rn6+rP5sZGq8u3m8r9Glccs/qAtMVKl4jA4BlFHgBvlo9cqqD5uN0kAdqw
e9XhJ+gbUXLb20jtuKuSYY87JU0cPnIr6gfRNNZv/TsJ2UsIQAJ16vbvndeIBFdm
Dl5x6fJaNq0ogepisAw4i4QLM/l6cqWiOPFgDkzFQzpJSBfIYJH1D+HltJeUdy7n
XNv1JDdVypmBqUoJi+GmamTI3Ndtx/PxPZAkbpRTa9aUXeo0IY8Nr+fktN9UHBDB
h+ehH5XXSyGVr65NSJ35AIahzmiZq9duKB79G4xXdo687NDQp67ibanc+239GlZx
pudpIJP11v6T/VJy5y1E5YOxH1T1dazZRpjnpURKrevS5DFUtV5SIMwSENOuHeIB
TwRJGA3AIfmkLuHcYId4UjXvTnLQ6c1C+cwWIQzsP0z7kMIPJfPbVCDLCq28mig6
70ZikggRNKfXekwQka93cE0vE8fOLHK1tB8IRozsuCAop3kq17RVf6OV8Fo0CI+7
5ogtHiw1iJeqCH6R0IDjdhHFA0SlDXHPZBeLmCyscdZtxzIokiegvYulBNJBrGMI
xWjY0TxaG6qqbajFKFOp+DJuP/D+xbSKExnLAU12ItCZlHNiXD+tbyRN5hw25ilI
d2zZK1OfRMoQLkxsHaoYY7FQkKB+LMKT7AwTnmxKCc6KhiaH1HJ6AItTHUfKAY/T
+NOycv6bVilUD0R/yQwjnHQAxb4NA3y5jR/dUzePRDS5IiprsGIzZotcYlV9D5w4
faynJr6lK5Ri3ML2dUEeNMXk2/+YtaV8eBNICz/4LoEJ//MvXDqNNg+qA1ePeML8
78ReHco/PXVGrAQ55sb/fMk7PuXd53ET3r8uoC6cNL9wNaa3uSvM6MRt2O9PAQtd
aGp+vqPNRtDETBIKvqYLg0XgTODMDknm6Wj9hAm5DhAySvbex9vkpy+nHZGYsWTq
cwnGz/MUQZNXakgntPwLrNID2zXIO0zXBzXtnRJjVIvc3TUtFVXFRoFe+A4+X0LM
cjibQqdEFrKYAblJRC8xcKSQKJoTglNrjVV6weoAtjiWv39Z9s7zY2y74oCIUkvG
p8mWY3FmVofZTMuqrk5D+BU8FCnFV/fbfXqsj4WFjB37mcmXqobO9puv1pHSDyVz
rPn6ngsEXOygLGONLxtrVqifTVUFhozjsAU9xS/7z4KdcHXdAji64iIAnOqZUWFV
5V/TmPbiRjcDlU1iO3+7XrF+6q8y9hQsLD0qxzol9BTQhmtmxb4nJEVByIGa7niY
A2GF0uFkZVninnhC6idNDLtloSD67GGuzFkHC5zJLJD4l20heqESSVYkssWjebbd
t8Jj/ikc7pgMUvjfstgf05jx84bSxWnsPA58ZUzSSYkCfk2W76U0Bw95kCzOnQTY
Vo9BsQVvcxza5ySU3LG6H2hcqRHhIcRHpAE8u0C/dwgfI65mW6IEhDFdDPqxopCU
Vhy2MkmBwqf/Lb5o+7gERz0hVUd4vNLJ79NfWoBxWf184NdnDFr96mZ4V5L/VwsZ
kVJjzbkWbXckvdMsD4NxDpap1VifINl2TYgrxmWGPWQ2jx1lG4ExvTwuGIvT8Fyz
w5ZpZps0fkl5m/KFGYQvodhjkM8Av4GggO+KMuDlnPin8j47ITV9bx7ovjKjRovy
LGF/p4bkxmCHPcxoMc4J/syloD+gwKp257sJHGSSMWyEyBQZmCH/chUHcR6oUGHf
eGQYXYr5numGIEejX9+5fm3hvl1cUkEX0d0wxyNQMmw1O/Tgdssxn1yiMruAUA3t
aq4o4SF/RQ458uB43SiNZNyVxJ2LRbrXay3SPku6mgVrg7n2W+LFqu2CS41NyuWt
74Ot7DVmZHQnSkSZTc0A/wCxEsK4iipmHYbnQRatCcn8oOMb6PHg4ceNTlKdmssW
eyluiIRdu4ROIFrVvDz35lYzo8arX8N6+Jvum2mpGo6jmDM9F7ZT92bm5f9UosjE
2IfVS8FVMdGjqp4xyFiWhpazXbv/2KOaPvonZKiYeQgUl55LBae6ff/rsBRe2lKJ
mB2SsW0fV3yz8GwHQ7MNq9Z78pgPA9zZFq5BjEjCyMXJGHAhzq4BQWPuf+cSyI01
cErpO4fMeqhyBBf+IiycEXoow6GcZWd4Mf16xOwXTY4OO30iu43T1CwsOpq6vcro
L+ZnXNu7mCwzjRW7ZyHnDeR4ZxUCSjvXd0C6cCvFkJ8VXCRubp7ARoX3s5QYnybw
64qQZmpWeH0tMimddqjLQYN3kj3snczndG+9MZWxRyTZDx3BKNglFqLFsNq4XIPJ
tppTmS4pnboUvD0DuHsmVQOZR70shg/7f+r12eNmnz1jwAB86AKsDT6fXRLiwpkB
cSBGa7Pt7l9TQYn+V6KmMyswjsH3v7prBCuBStgwzvlNanF2uvPUp8Ss0D7uQo3i
uI4t1BsWG6JwOjNbobmiecCO6/aLYBmE4CHnq33U4pL6s4UruDupvbCalRySZ5LH
EqcKsxu+FjGCEzGFRj1jStb1fjaHXiqo0bWmJU75Y9I2HDjSepISEOK2AuydVW7D
seK0sELgdfaCpJlEOZ5NHeFv2oUu0jlUOZLXE7iGG0m4o62epkPiq2E8kos2XIDd
Td7FmpE3fskfRRCUvLdNt+AUzBGYtc3hcL2o8jKMTbJzUYabZO/geLeeyhWdCdDu
yMlmpTp+otUmNIt4Cr9VLekWmnKGLGKJf6ENN58p5cKRI+9PyYxmWkZanAdwysgm
NcDocajoGdVZGT0KwKRzao9a09JOPAU3vDi+SyN7PHTM2DKep/TADml9zYG9dmBh
npefWg0sqzXeC0mFZXXJdmqzkWPAsozhRSAEELxoQ5FkmU88nDcA+elVMda3tnta
tp7nXciFUE/pKb9Cvd5EEgr9U4Nrb/tUTYj3JDIDTKuqenDFPvRwwKkkpul107FN
h2rULaDXNmFrGne6EH0vbv+W1rMWHX01S1wFkiDVh2cY4DCw8tCstGLHvGH5rvZH
7f5wNLeTtAkQXKk9uzW+3SG6vV/Ei+7HQ2YjlZf8yFVDtidoQAv6hAi+WO2JRf+B
z5wmAIHqbk0O83ilOBkd6BfgdZwrjVSE01fPjdNeV6/c6fWKlAyfD1uHBRFEppea
i/Is07fsXPOWZruiyKNFHDkLULGeVECBpmnDP53T1EDNfrB05ZaPbolTV/Jc6nkz
ULORV4MmRhu3aKqgz4zMWvo+dkVBrlK0GmEnxSaRUqt7yASXr+ecAgxqBu9qwN66
CQVczsET2QLAIiowJcbnx9hkXjbnVk/YBjCL5TW717aXdIdMgqx8Sjs0M6umIePl
L3rVS9wd+fp39QYBlvaN1ZmJhFEqMPF+8zN3ibfFC8zy77XyZ7yg6PTyKCVstAPG
8RA9pZYNrHYJINEgn2Zx/DjZveR8kaQlxOdDU0wJPfKWGtI6aTWA2MYE5sGllrni
2d+VroFyhAOfGbYhoDpcDMVSnqymi6KlEuE0YzQo3bplbxYTnbaaCyiwSXW6UhwE
U5CO2sW8+4anbTZN41BqOl9/awMBphEZOFzSlEqEksemFJP5litH2nQdsbRYuGjm
BhwlK9cMPnOWcu1g0n/F1Jrw5lkLSfkn5JjuUWN0QBOzzVTQSAN6AlvGSF/QC0Yx
wzg4q7Sy4XMucnB+7nrXxQ5XkTZzWb5XAlx/lrKVHm8F3CJUN71HYgjF5jk6Db27
dcjkctLQZBSzJjEnGI4yaQ8CBBZinGUdKCBTSRYfm9SHNoufEr3twVS8fty6eRb+
fvrYqEMdNaC8cN6mcBYCtmPYJQ17g9vl7HEjc9U8xi2Lslca5GnoaBHGDBxQDSwZ
b2dAQk09qy7N0XFaxzMVbb8r27DZD+yivxgarFJj9HTmZKlFobVITbv+sSGZtP6X
Oo8psjs/hJEEIAIRZi8TcoBs1R5TyU0MlSzQvh5kKrgWVGoQ3ju6W3+fQPLAa72H
GGbZwm1QGC9Fc4uxPoiBJeE3mZ2yGCMkmws8Q/j5c90VZ1YzkquBSrc/HdYzDN9O
Zr7ZH9bJJz+IsX8pcbDaryEN6dWS7OBfXqLBQSiYNST+52uj1o34giaxLwL5DC4+
46p7z8/arO4Tf8yzCfCsHEi3pNtm/DAtwprP0xC0jDmi6+CUfeapTAtkJsIq8Y0J
ZzGGZkQ7KRE+xAmt/HtXuCTkjQuaJ9ghO6fYbKhMV1t4ub4fU/T1uObC+N2DuecD
a5sjP4sOjokDXlFXqo2OuCmc7zBL5PW1i+BCI2YpG/QNNmj2NuGOAu2xm1gaV/ny
MphcQq2OgLfeSirDfzj9lBkNJAsUDvyXOllWPj6dhroaRuB4PvnKsy2x/82xdlHR
zwjfYPywB7xHO8MLSeguSRNiM760sjm98SnB2r9yJmQjoGRXgd3j8RD32bw+EnHF
kBzigKOQ9s2isPdQV91wSLxgssQSSSs0i+p+GCcDeSIIh5Fib39Yjpa23yibVxrd
+bLTsnJ0sVG6aX2gzcte942WHbAg2bRjEvHsaNw5VU37ap/YIBmdEFIwhIgL3/t6
1ZrYawm50Yg/PTAXlTdZa+e/lg7UQzHhgCWs/1Psk47/S7jPTiVY4c0s6qBeedl7
QItbZoxjoULiY46alJi2MJc5Ql01kibe1EGf8DRC/bcDeHs28PsxZq7Z3SgzI147
82gkvtynhzUyuYkSHL0Y21XxULOf3klRdHm4u8fL2LT/p0hnA/0A8nkJUo/ZwV4a
e4jqLBxF9aGnai02RtAB7tEW6KiWUfmL1df1DdfiySOD1pgQ0xLB0ryUmiCU03fd
vUqLg6Z3Bk9yX5mB9cx8IZsu7IMlliRoLXgGvBOHfXqwNTtyrVeovmEyOBUSGm2T
wOUBdIzfYWy69ZZoAFV3pBTYInAIVYAmIaX26mbXPOZH8Lhwg6uFHtT03KLjriXj
9B5CC3bPeJ0cVyBsudbkThlLsUgPwFzfx+dpb8cFx4laX4Z/tv+aNVR0nRx56SEA
pJnjf7Iiw5Q/YqQUCKfRTHGm+ieBGM57V9hcyAy+HXnboKAA80jhvNiOY96M5jnB
rQjOb7OS4FetNPuHgiev34ZXE7K2gKXk/ayGHrrXDaaGJPOrbB0XLJRdTaHlADbA
T9itFzHC0kLeqjnhIuqpaYd/UvZfs7pssRIXrPloGlDjfsbU8tPu7h3NBF5lQayF
1eEc8bUY65AypqXTM68ScmweydWt0BnNMDmPJxubd2yAIr/ZJV8X6+jP/94GKQeJ
aS4PwYRyGfhOX34G3c54w58rWtxLP0n9JKWlC0HB2qihEoFHxMf2rLpxbXkRfjNt
j86BHZ6sRGImKlYodCvNzt4Y2UqvP/IhNSMsVJmq2B/KjpT+FJAikCB/ma6e8nTH
mOBCkYJvOMt9kZE++4xHJkSJ53GAmFkrEQIwJ70znitCDkYtotliOPQSFv0lrTHv
CEnFrCwVYwbsc60c0CC9NnxWgZsafbbWutc1Ndm7ZzZEX6KIjbjSSgw8kVi1q7/b
4c97b2xFVOrgzxlpNZbZ744JbCGoul/V5ProrLb9wdsRbzr3pm9xBGpI74zsfOC/
APponv3NP1j3vslf5Maq1PhvLV5q9qj7la67hV5k6uI6gTdv1pJx6iExX3J+Hm2c
kpjvmLfuPYSaf/+y+mzZmO2JpPmC9ZZiNGD7q4/w7qndW7Xg4lIQP/OWX7FT/+B3
qOtG9NoIx6AqjDNLI184uk9k+6sQUdCY5bzQexYjHbonHV6nsTeRwnyWHTm1Ch9V
WAhOGz1I0B5TQN01K80IdHIrnFDZzoEEMrtGqcubWB5hd63vIuxQMeR3wTLa38rS
euwhC8sXgVvBRl5FMypgvUo2ehbn+cFpYS1lhQ8ea9El1I7bZKjpUzIws5tPenbH
oEDNuzIBUKsuMEwzvx0RToxgtSb4tjNjqgo/L83RSUy8AJmguhPqKsu8dReOGsus
0zmgPJR5wVUpFKVWBXZhEchF3moac8nR+84exiiBU7odVQLmwUzRwFeX8kpuY1v0
KJi0evu+CpbPq4rLJpENv2vsZiBPtXopqZO708mdzYpTjohWEAP3RVJGpskRj4Gq
dvuoi93S/m3m/YawtIRTsHBPRAT8Z2DbAh0TjhrzRa4d9QfL093ppUGNIHrLg869
AckYjDr1JxbFGaL8tr9YXWzuUYjCkjome0rzebkSrrRyNUOGF+aYhIgbplDDUIW6
ygySFeawOuaEXh6YXNHBOJrdoT8KFFInZj2kbLK1ns6QMigbU5xa8X/PsXVTDlOA
Y37LqCGqthLBE6gY0K3DU2+C6LFwpWZx48p/B3tfgIgScrYf/EUX0zfGp+d1PKtC
mPQiGc0h8VOjB44EYKlPRyR+kDy9xCc50RDtT+gyTezXt/KnXNdDr9nQJ3LzIfNr
7EXX9FM1LFf/WyI2YvGgZAUQZa44FiNAJ7mS+VRi866KsckKK4Xt43XC2rRuleDr
4YT9MSkzm3T3YSKOQkdCYKmMs/ESOSLNUj0A0L3IqOmxgJeviB9fCdZVWVBfYmWk
4XT20vtG0Y+FF9Cag0S3rBMvthO8qKKeamUDvrrUyV04MaIFM4tlyFNKZBFYSxA4
nM0gtKzMBOQzT3zZmKz7nc2g3AY/woJ+3wyvegSd05vowU1czUW2yEghS9xFgfnO
cTk2KRPPaQLFVyePfs9SDgD+Fps+eT0IFO75IILvguWuyTBI0EV4njm1GpH6Eze1
q/dFf86K3aKu+FCO09ONbnCS/iZ9SizmsvLvl21sM5gQdIX0l2sbLHv7F2CD8AY8
YWd4lC0sqbONEOMmo7QzVREYuxU9JpioKGy19Lo0EvgHNxrTugVp5pH3oPWX/wfs
YEJRS+LRgCAg8h8qSuilv7WAwTkUEfDUOW8bwrJFmQzC+q/QhVdjZXLaqWK8St6s
DOFpc3wLwzhJicFyPcaYwaiIAE+FaOKeBMjKPpTEZBuOpEtRL+zkmc8kykoPd+kJ
A7668015teq23haMcajSlOi0+kg7XLSRjxGPKqenVEPstDgQHfdBm1ld/qawmZBo
qu5ACAJeVmQrrl2WyA7p4EZM1xsrOzt5UpVWe2hqooXo/fAF5hlixyzrQILirVnT
k0V/xXWeAqv6udNyhRVxSGzZo8FDtpsRUSmWRw8B39C/eT4qH8OEf47bIRNLHw6j
m4ZTi3zn2dmLNVbTuLbhB25xtOYWdk3YS2U8lcCIHcFITS6vn6BEOTFoIAYueOHA
9VwhaU/tOaHccR+I8XnvGy+bXC59434pdD/yuBhTENgFdnDRyvaCYkeZlv2liJJ+
aKC6P/NoaevnT8QU0pmv3hry7e+40Q1LDnXK2+9NQ6owk5PXqJCXuFSnnkf4aJLI
DOzhTzeJ/b6xUI4tcShjjGhblyvTC9hc97LVQ4QJ6z33qUgM50wlekoQ8AuVQfyZ
hq63G3kACyJSwZc8wdWSIhAvGSCdmCzImbV36Wxm9Xqv5+eMQznwKNX5yM33Bdm7
ieZrlPbvRcglVFoNrPoy7ebWkH/pzFBOt+xj7hUryOnFrmmBxYC/shOTjAtfbvE0
a2vb2QTM7GF7fk8Vfi52woXSRWEJkq/P75CM1FTt46/ZMulUP5rxewM4NIsnhoDg
YCFuVy+fNJ990CovGPPA+V9svcx7xM48Db87QdDwDeHY3WFLNLG4byBV8xIQW7o3
sPpvUAE+MYvcJzI4B8a6UUHDVOOqhM92SaVuXgehMxil2gMnfAN+W5HIPmXJH+4Z
BjPfHbudZ+oGW0qgGxqYPDbUaBeg/f73yrptt2utDMk4cYfPWGJ85KhcAkB9uKKE
y0oE63rMH89+m+txUy5gLETvODV9d7YSL1ab9af+u8UbvZU+AyTw6jL7MWM8qSAN
JqydrCdgZksm3h6FdYfL0+vT13RzODQqKyZKieoJow119lRsgjDOahQD1TEt9REb
MbU9nQbRt0CbDmZ6mDsmL6CHxSAdJu6QSqb1cby3EWp1bMLQ9noKmgqYr7LjYCw+
kzZkTIfg6TT4NgUL9rY14zUR8rfylL/de8Me+SnkGWSW0p3fSAyN7s31io0QXpDq
Q4SCzunpDC72xFr5SMgBUyUcIDJWCHNhGB/vGdyXeN0CIGV7ydNXjFA4eCxgyeeI
gGo/LsFC4QmCV9R/Yn32dD6MQI3uX+7hGLxIPYhgGueQVbt0DWfVaFNZqZ97a6Vq
Ho2PCt5MnZjqYPtYwVvfxSjG+wbKXQKiEynJitgXAlpljfX7fnc9ndhgDYhv69Yl
Pk9tmHtcb6GOzZlTXaXKC4mcUnJUahgCARZkt3HKnJS0NgrCuJpZORPvHRFIUa9R
9i9rQ05fSsD8XpKTS7ZZOU834YAJKReCzoPUbjqWjkWddkIQj11vJWZU8PnGJK5f
oGdxyivbqhlm870DoYkXB4akE7MITif25F3ZlE5CU3rQsOEghWu3t0qLkXJrUNJZ
A3JvVnsLLbfqmaFPoLRYMk6rgb1bYKSoSOo1Y1cqrLCTlryFPmzLPnNpUE+f9QxR
EHxEUnBCrYpOvvu2wNuSYLHtFaEdn+/mtWYBTXiojZKTvh6+mmhctmFS1ygFc4v5
JsIHfeMsn3JPJtjCKPLeQVe8FIV100mKmlqkxJ7bC9A9vUh7sA0wsJT+GVJFkHtd
o0G8jMOmZzntmlbF1Z+eGUNxaVLXb3t9czLHI4OrU1Gvr3ddAAHTQqbdBEFP46wm
7xGehuIqlW7sGtS7ydheSDlzi9RZAYAm9Ytv02h0XM2kLhKzYeCXF77SNRmT+QfP
e2ct2GvmG+YFk7wYbTigpI8S1FQHhnUVBogFEcRkiSW8O+GhTSEs/09NE9aKp3Mx
CJhyzB94pIfs1tUfBuK+cWdda+rCrmeBvyEae9vNK2VGyaSRtZqOP3Olth7lZ4Cs
ogWKtm2c/I7yLlP0Jq60elMsI+IPT7dqzdGxONW3nUHsEO9Mo9GCVAE+89aOUIGB
9yVIofU7CebMafa4YEsRmRL8++xtptlGRL368X3LtS4/T/D+xV077VA6Abr50MHL
wdClmhcHgQABiCVRN0NorGLmK0lhM7yLdhCYOIauQ2gDDk4grdSIgWT0jh43AREE
zrVusrQb6EnjECFGGCu/4c74iPACluO+JKNgZ+k2xIFfTSpuovXgKHk6K2tmJu9z
H5HoqtU0R+El547Nb03TUnSM6ezK8ueR/n/9hUuUJJO22eu3HuMydmKWXnfUlGaX
d/tUdD2iR9q507TkAwPGAgd0ewmIqtHe152BDWCb+v+xSdxJXSxkmMWKo/zCVONP
K/+4CgZJEYsRNFQxsTvhDzHjkpblZ2v5En4oi75H++bVpvuz0hCQ3yPXiNZJ8GqO
eFmzuo7KcZJlefQXlBC41KLv91JWHlRR/4dUG04Qtsvi7tLBXGZ5qLopWxNAo6oN
bI/tgS+m/GGYnLnt5VWDWua6mGGCYp+8WyRyAajA86CnRo7OJuw2b5hD+TV5CZfb
Fj+Tn1d7PoiiHR7isRUyB3yNWgOlLCF2bWoxcSRVmQSXbDMoFCYtuzDykrqw/M0K
+CL0DmL/+CK+8UDkt8wdh6xiVdPt6KaLo8QxV99wL813am1wTOoU13R/985UAKuC
2X8X3m6rXZEutNd93SA0Vp0cbCjYix+CUXU5fRYaZOePuMeJDbsqlEQKf1eLSM7N
L925dPVM+eakGJ92PTjwgMJWadeGq73RQ54+TKkRJxcUnfmn/nn34NC3FfzxB4xG
9uZ5qp5Hp61TWF1NxC7+1MIgvn0g+vOLMHbSFRl7BbURNLW7TT6hyqkDojkatklI
pZCPPfB1VaSDFfzZRYzlPyETIWGBaV/O2NbGwX3nnGMRRy25Vj4JNOVlsvwZlSuh
kqRhQRr4ZDjJDXQJnWaJ/FttrVpuAa7at+5wE47XIztrvBY1jjkbo3KOBjj91eIc
18qVkTmpYyft4vqKwrTfDKC86c4lSQkFPTQtffEyQDTOsk8gp/IpteNX7Za99u0v
k/SFSXAIXIsOO/fR7YLVYFg99aS4jgUdezYcWfYwB3aaTzUj3LuB4kuxiU5Hmy4X
Xo8gziRmTLfnQxZQr5xSZFcN5/JDxO+/r+2fGFb9QcRbTDhgZYA9sze0EnjeUdbx
8XXA8YLHK4Sfievi5Y5m3Ia0I8BTUp64nmIudbgtLiBkDhBCUE/hL9Sm83zcoI1U
YFWA3T3ppq/+1eY6Qa5I/QmwbLzB92RT4NGX+t8b5tLQtnd24jhMIdRLfK3z+cEP
AOmSr9MVWY1F9SgQvGqYzHFt1rRfC68fkRfI2OSbsPl41jjtT9aKqB+LfzWAzqs4
9DdOXWjZa3LYdIn8DY/mS9sah8/QYUkThIwlIF0uoZd/iUxv4si6qNSMwqNj94HW
XTmU29ALDsT3OpQyCcy18IdMmqz3NT5EktvK42f+z3ntRP2EmLVnwguLHuRaJtJw
RwCQIGu4IUjfqCuAs4jjfSCgz5raLuwiux7jTmkGutL72AZeJkvnbUXY9JFNBtaY
WE/pWTr/ysb3mo/NpHieHwzdcdoqwH45zktiCM1drp4hTfymaUE4OvJ//4aJ5TIg
RwTypXxB7vXbpnq6jXJZx6LHDpuyqjjLlgssHW+932RtWj9Lr1rMt/mjt/H7itwb
zVqgusm9wXkT6Pgg/r2DFGkImW3ikt0jztkNuKvJupvhsin19kN6QtrkkPkGipey
WZckyAMGthQSflO1VLa2uXfVfIBxxpUEisvdGs0QUoOYrD7RYBoXDlxmxErAsGrs
1Q2vAc6/PeTjOo1MAEyWEW0joJMwTfT6x4+vmXyNUgtsP5qUR9saVpAa2bVOwdbk
PQcoAhdhFxkE9/+t5AoHsMzhKcckWQ4grUz1jyRDRGa5lOW3bzUPO2N1AvjBnz9M
BHGqzlPtYgJbttKr/d9dsrSsQNkbi/G6+vZdT5HyLs/Wi1FA9VS2dPo8KtDJGIQe
CC8EbMKESjnNH+iX4TjA2gLRKXwNLjxdL1CEI/sfpcNF/gWUOiqg4BprE5WokuFS
9+AoDrP6rQ5KDrPk0nbhPm7EZYtE/FHujGT6VJnXSOv5IQBepBrWauwf1JorwOvX
RfhHpOkTVlee95prIuO2gewVtdzKepf4dBHvJ8mLpP7tQjKtjfc+eTXeaY6/cPPj
sUjPGWCzrgNNU7AxpROMfqV4zT+ZeK/qM60lz8x1RsUwjBeWjqU0KG0SvHw/ehkO
niQfrhtVWMbI6ycvegu1ostDDhyrxY4CLIcQZDAJaNN6l0927ho8wPntg8bWKsmD
crPY1MtydXN8tsObg8aWOfik165fg5F2uCgNhLkprg2Knug859XQdbgUelqU5jR+
07p8mmih+LxMVN6F009PkdpsvGCmc7mN4atnafq7KA/pLfv3e710QYsognAX/bbH
9mjh+6/pK/5ixuiZrbIPlovmOiEALILWhfIuAbynw/atAvBCPwXphr6RS1+zc5Ma
KI/vS0aAAVIp7/zSrinqBsOSOyohRX3l09XZvRms51095YhOsfo5mKHRzBskXf6p
4GBJDBx9rch5uzgiwtyFEu5NBGmND0Tm0cz1Oall7SZX2M1aJuz+8oKGunJDnFJ9
FZZTSibCd/KQBDrdejT+8pfQ7n06wgbmTF3zw8XsWx+zm4MXUUBUB0BnZv1kgUvR
ekFxlfyQmPeT6sXzkOiPErD8NSTpgGyAezIRTSfIbjxW6R6GlWJvSaICGyg47zlK
bmynAAHaHAjYgqygckICmKds/espBtMHp5rvsQHSGDhR6Z2RfBK5UJHIXAxe7IxR
NMlC/uf0989v0gkk3MfP8m1pDFXBh3jHS0+bGz5t0DTP3NYASwzDexKqfKV/H9/+
73E+/lu7AEIqE4cdMiiZ3480eFgmG1JRkGtIH4RKg6Iw80kXiT5W4a2L1XyLsep/
CUFYzKjkjqK4cpOy6hhi9Yhu9Wj3JRQdqYKhz/lWWAoswXWyORUsNS67dM9riIGL
xPcQ4+zzAWZL3PwtsvNxdCVB0RKAoLXli//MSSSUddt7eevI+dI6d8woszCYJA5M
9jXy7ufqoHQH28YiJ87k5gwfz17S732EQBP5U0unRkpNNt60iK77qRo+yWw7nwlL
XiRy972e4//WNRu3sUmUzFz2L1dQ1ydvn6AhOKSDoVphEzz++H0oojcC1v6mV9hc
bsX01JBI65E9PQ49mqxwJtfjID566eutqjAJsm+JdJwksD6Med9XTlhWw8QbC0LH
UmG6wu0ehUN7Xt7HROQ3ierfRP/B6fs4AehVniKNEcNHzpmJk4BW1a9m1NJOPma7
LWB8omJTJSiY5sEfJvqerwpgXWBAAOiqTRHCU/zMoMpkV/23UPzkxDppXIYYdb78
ZPYvfpl7UcB4qAALMR5cg6zM30YGVlr3xfjt6Lry9TbhPKZIUfhJbv1RYUzDO9Zy
IEzIfXsrvBNUCwx8cqqPw4PR4ntWj3wpYMbyQtMWnmCuTePvj//6l8+GV+T9D1fS
QoUzna1O7HlS5YRQnTVDTC3XE7fKysdAmDHmPGtgHQRTWLAvTkelXyNXX0mAC+8w
cXkmeM7ZoSeOSlxrbrjOKJZw9q5w9XOWjwJujKZQyR+cOOD7+MRY8DYP2qFg8l9K
KqlduGKSomG3ZScx+EzG73AKTh8qQejKA0jHBLmaDuwyEx3WfxW9sLVTe8SHDmgI
0EaIoOkHp+Yel/BFVkgXXelZZvk9L4+xhRmr7rSKxJ8QcgNFJq63dH+xTIVUu9p6
s4NQN3CywUpIvkbaKTBrgbmMethsgTj1gyuWR4SKK+zRCCpHiLPBwgYn+x3Ay2qr
SEvK1QlDY87eC3HHahb6UlLP/1r6sXam7fh9saeXB+IUszZUZ6cb/3rX4a5+pv8P
3daKJEheuJWk3t0klR31HfEW0DU3x5gF489KwFu7u4CGXR4V5RKRVbzLBBlpm/fe
ooWZ29H1mRIaN4ZXFBzLmKFQLIDHbiksvRbuYOlQxz6lF4VpwpC/JKJnHkLgH36B
xkMvBsiGzXZhuuSmFECLevCIa6Eb/zhTaIOuLzzv/2/bbuboPSRSZHbHskuEVuLn
MeBlTbz1RGHdIXcM5qaso7y7jGaA7UkDsS8GolRaMdUc5cNnLIf0L5FqV/TepZd5
2hJk0mKE+e49dXi+Hh8J2Xh5zadkrvrcenNw9y3Yw2W3ubRoshp020W/PyFSrA+U
E2Oet96yfmDG9eD1dfrFFBeNmqnHZLMal2T8VBFXKayIaN09VEGjQrR97vjiAkvq
4W/dyX5dEbnVHIyivP47ZjJEN629ipdkBg7u/x1uFElUP4VtSr8eO+gV1Auktesk
oCxYEUGJUOeMgmCwbOWjjvfYsuzOeyhO9WUKUnvhRihwZE/vz1t0hp4CQsZpCBjP
Ttr8+DlUr22au2GX0pn5MVQcfmwDAR3h3R/J9paRfej0Ya/jDfMfVzNTtutTonfc
cc2mSC5HvOXaenQNtS2jRTOzoo+kp3deKUWNrF6vS0Xy/+FlcgCfMxirMGWkb4eH
nzH0vFCCFVgQcdFl3KNHbqtHrNCETBZY+b46BiDKaPIzV3qyWdCtZXjPFZYLK/UJ
BxqxXzo1ruM0NcvgoJhtyO127QVG2Vo1pZrBomrWpXzgMVV8tVLnMMpY95kA5W/V
N33PHSr5blqo3bTZLG+xXgy4GP3sNMPGIe/jg+RhZF7dlWZKWmJfCTGejy8n4nn1
wGpn7uTDfjkS6EnG4FeFX3sLE26QZUA9EAorarKcdpR+/1ePkEt8bx3KFtBcirt3
u9ThmB/yMgMo6PwhfH0M8CLUybGYiDCZkuc9bNYg5LCS80+3kwV3HGzX/d/DeNTF
uGH6fVL4VOhZzaSrdquGDw5oq+R0yJtllQ5TQ0A17kozfq3TRFDHX+w0sVNGngbW
DrLKx9s8ZpJv6ToL6d8NpNMvjhWqC1F2kGLT99r6AKrux/+n0bfdx6mgEWgxF4fJ
R3rKV1/mpcHNxCQW9liQuq2do7hV+7he6IpN9vZqYb6ZbOvCqlhdORzwtAwJyspn
XWx7Sn6ULJQJv80+oDPYAtH6CoclkqC4DhrcX9GTDsD8WHuSym16xG1eNWWmlK2S
XjXKZlUZUlTV/XQmyFxvbf1KoLtJUxq6Mq6XpSjpDgs/A1LSdu8Q+2KF0Zgd7zr6
Z7RFK6r8dyDu8fvlOi428/2HAQ0JUNgl9V5T9kX1SdR6RPApoRlTk9TlBnG7Uq/j
xD5yGdgU4ESC+HW59WU7SRgRHXc/BtsYfuyH6C8jh+3U34iqZPlMN10EjGy4Nc+R
sE3wbmBmBXZ9cDz65DQiZT2Ek8vCGG2fIuzSFRDP5NcDjGgfjyat4Yn01kE12R3B
ze5SNi3i2Dln+GkCPsjnggSfd7UhCsI+MwBuMVxIP4/SqiAhEy+3FXgICK6Wn8A3
KAyvSguPvMM4MVfCLaK/nZof1abYo6plGcxzGlxRzbY3Mv9ka9nh8UkbY0XAoJ2S
0RbhAHBptuFjsoDNGp3llwLsvcyWXvp2+Tn2vpSmJoa/uyG85UMu+h10YfcgCYqh
EUsepF9eXQyTXi8TwiVUiYwM/iDpnqtq+o225yt4IZRngtig35sS6Kryc1FMLshg
nIJElpNwtgVNOblWK0u4YP6hLhww4MQj1DUe/f2k+6cxJuEi1OffGcoBKiaJmAO/
gtDrmxDebu1AcL0n9zicVt5p2wD629dTnJiHkXizbWOAtVMvhq+hJ7i5YY/fPTPp
SD2r7KbmKwkhRHiK4rGZgMzozJOhW387DJkX2VKW6eBE0Pg2rOSFea2yWTNTFWM7
7aN25HudUheFJLut3Axl0Md/dnX0HBsHP+77K0uoVIBw8OzLgdVJYEG1JCxI2ZXA
b39VGF+QQJB3RUWvCVqwynccSI+AxjMPCpP+C/v54hH8oc2s4XOtuynfX5hevfQu
H4nNLsR+w6t2qvxp7M6t7iDgjwtYcd153RCiXzWgdjgB8iBdxbX+cAiQV0b4mzgh
OsoREDV9e2E4zZolBf/kRFFw7hePF5EYIFTMQt77ZvrVGj1PHLWGUPVXEKUAEKmi
/z+BVjeAKIRN3Fan33KBSLMuRvkGGmT6k9rUGEvEZR+3D9p7z4H1Ce2IANXqYSgK
KNoZRwk4Te1dTn3bnHQQPlyXMzYTaLO0zTEU0JqhRF5QkVEUvhMWRQGKJSqmOZ8l
Px47Bc9vo8Qml1x1SLQBNQ17HOGVE9JYX0lIyfOWGjaSrcDzhAeQoTQBpk1BzIv6
mULLsqamGdpzcwE+nHSA5cCbBb32Fc9yp1Psz3mmMnqqSdNMuZUYh2TnhuHW6Ql7
cOf0ZQ+63iPlRkHM92xYsrdS1HCg1cO07vt9r7YEIxhDRK13HLC1Mycw9lJFjBfO
InkjXmmogVcYuWQvwuwLoyPMimo8CboTUvlaUCJ+GtFcbBNrD+ncicmCPNRfbtLc
XEe9WL3n7Ip3udoSLZLdX9bxq5ezFqlnb7v9DByOsgfwZOy5WcPiTDYRe+N5nlso
oxDep++XOMx8bTDcE6115i90BSz/S/K3OWpbMiJ27ew3K8b7bSkWaAXr6fkwGUae
rdNgD78YzFiDWrEC3wTtvwRgWnXr4CI1Ug+yVIDza1Bo71UBBHnn02EuDfWelG9G
uVAWpAis299bRyPML2Cs0M24n4SOuOs3D+e/rso0TwCWhl7a/vec7+js0rvoP1V3
K/KpT6mSl7QRtrl/BUSJn3bjyHZlN+2zIx/ChgEfbaFRE0Hv5pnTovQUR3JGKExD
7QHapiasQxDQUAMQtsiRzIkNIhI5XX9p+NUSguuNizcMvs/cE4jPQCLxeUAZIsgB
6yPQ3qeNd/smNOLDzuXy3CW6gQlaZz6y/Sui3vNeCxhwbzMDZ3LB0d4rvDOCw+RU
rKP8ATct7aPx+LP1d7IAY0B6qrEUQvtchM1OQIxgV9sqGX7u0q5p+6wkyNCUW+FG
0F14u+xiVQCnY4YuqYPOd8KntifaWwcbB9sbhHsi3x1bMQOCk9n1aneFvsdDpXcU
riQ1s/keIKMeNQlmoh/wzWfxeZOXvPiw3RVSVGq7RQPVDLViEaY9pm18XegLf8RD
MNx9dN3WiuwF7hOPyxpMXTTn7U6I3EDPmZO6bGORnne6Y1xuhU2S4TH6VmIFTxnC
A5Ti0Fer8wQx43amwvdFk4NYA4r9yrJ9wUizYlaBWO+c3Xk0tt4ucCqxCS8mg6b5
tmeWTRfjC4FvXnMIAo8J1AiWCnHPGTGwgLTZMCBv4047KCcANq7lSWtkihy3i3qB
aQFJrhEBQI0tDqsU+IEmi3KgM7Ks//QcYez5Ry5E6iS0ywnhtKkMGNQqXglN1rb1
qIygEI/oZxdHGe/xMXQU6FRCMoincx/7PAUcjLAOu8dTyDkXV6CDnRzwZTrU3Krj
ptUbi3k6rY64W7i2N/1zp4Sp4i8YNpZDe7+4jwMRxlc3fTAz75aDiWcbW/sKDQ4b
JXMq7dYHYNSlGLfJQgrX/6u6nCTwi/5vEMZ9jf528T1tl2AzZpNSi/pktgiUTvNT
yTUq3WjlbdmsJOTnt5LbJr9ViflfDiVynbQIPutbURCxutRMZCzH0va2tZgMTzMN
JkNVcjlf4tDa1ov5De1pjKJ+6kNHTh5f5tGurdbOyEKQM+tlvkdJwK8O4gVl/Ar3
g9NKQScjUdGzTox/3fUUOcQ4It0c/RjdHsPxkvGVRLmT34jReEOm5h806X61ER+s
fkFdmQVtGiPoIJI4mYx3RP83nIULQgn81bWCt01Pm189V2ldL8RjKKooVXZeD512
Ni/Vmd49lELYQSrCfnbBdPDyedoNuGyjWxMEpQ9QTOul1GmgadwO7cpHFM5oCunG
hsjygcMLUrCgUVtnA5l1HBjS8SAdUF1DF7qDwlzGv9+JNVAMmLvPzDVQ+xCBs3k8
qrUr+GrBmdkiZJ39wxurkNhUzBeehknfdSVajYvBmHr7dOJggSTou2XqYanxRv9O
/kyVBgOR+Px8H6oHeHZd7aaVTv8QFRY9eZwco+xnhqeB0/NpQdLheJ9gQ0ghCwAu
yWwytLVqMBaAzdxB5PpmVdg4OegnvrKTF+hiS7jaIV/M5jqAGl5Rh8IxKDH5MQFI
PyrfgHY+hRPEQcyX9xvD6tdS4UuvHXHC9ojshBNaO/IbjgxBilw++cJAfo0JmLCM
FOdAAmGX6dR3x6+toxLVW76w/mwWtga9vn5R2dQYJimy1JcnyaADuHgNCZslfyMc
NK7wG7hZzDnNXeCW8v1TcvFufk99xigbh3eYRADXE77M4MREv6Xqavdn24+Fk2WH
E8N9TQxWSAYPSI/1d3MEgnhCFhM8Db/pTc7lL8ACD8G572/CleOv1OEsk7rguSPB
CgxJjKkwI0hR/7dBRXmjpYBGdwsrWYs0ysOeQDYobGQ1awhpN29BQjYLPRsNclzD
/uY1CZVv039SvteQMzoxdNmvMKQTlBaB4Pg0zPTmPxkHVUqnvDu7/QVo5EMjSNHB
XqOMsmH4zr8XuLUiMR96wy82ygeHvTmPVsiKTdroZBWBe7SSHSUO1uz6hpGyOdEb
QU4nay7xFYmp5qzCzq+QiF+AtWvQs2bGHvSvjInPXlFWVFsNO4p1P9t4qZWpZbn+
Mwp0EZpbBJQ58iKN3rRjI8VlG+mS+mgb/hxkuMpTqUcUtReolttBUgxftIajmS3i
eLLAghznjcVMi8Y0IJU0qUalUs774YvhKqbr8t21pBYZAYkoAWWtF8Hjy0jKwrpr
nzkW4RwOab1P8Uwo14ak5syMgHOGTtwHvOv+fi3HqbAwCvvSCmc+AerZjTunA61V
dKYsxmf0qx9yNv/XESxheIDi2Ta+6eWtbLKI/62BBpKz01+Posm4MIZJbvJ3WS2Y
m6qaQrfJIzlVD3Law5GL/ofzlfonikQXDtYvkP1h4jpW30CZfiqt/IS4TgaAn+hs
JjDBc/zC5j84E3zXYCHK0aCFXkn3c1T5UwyY5I2/4I8IV8BUn5E4pwAdKuG5C/FS
i1MaHBNrxypz6dy3rHzjI40on8BISOxf3Nvu01jO5KvZTk0eBBm7UTL9c7UOOGh0
Gte5Uc/ZcuUhsiGVKfMhQ22htebyvxAxBhrW1Y2ZNgoj4lePKADaEQT5hCxcS5wo
hjjmOnyCBq33ohTde7FuoPVFbndnpwnaLmzFEXY2KSDpncGbwAMNItJJ3BDPMzbE
nl8vtY9yL85HvK4bUr/lJVM/0x9citl2p+DfTpq1++Fzg9/wgWaCx+D9vOA1meWj
6w4vVnkT6b4IsgPtAvFOilqI40lsvFA22c8qM03EcmCBcKx+e8sdpH4hg7FYK0nT
/+XhjyZXLHnkFVNsS5OWdtwsJHYUmzMsMg8MWSVpi43Y0aDhbIH00scxg5IwbiJU
MYn/gDd2NaKOk911IbParbEI3nYPjLTxoWj36Nd0mH7OgEsZTzOwwAQWh9xzKWvX
2caZ58zhWkP7c4yGqb+tui+oW1Ndl9glGiExyEhXkIpRycLfCVdkOjDcjhapeVLj
ksMj6mka1teeelesSwhgzgUldlxvBQ7fttpt01o0LrjrAyKx4rmLOuep2EO3yS4X
e9eFuFdBtAuvkl6I7kszqDf/OJvW6AsOdu25oHHyfzOIrF+lwM8gCbCWH/dkAl+D
4jVOI49q7yO2JAro45ZyF8fQDP5ux7WrQAC3bp4EExjeikb2ggBoeyJAkCR6WyEc
iOHSVml9FqwX8j/u59pIdtBDcWHlSeLLLh24AQub89VXNUFlYls4wX74RWXoGvZv
FrlPYVOJDrZAN0TTTpVRzL6RgFkEXK5emKhT1oUUzKESQdZJBVy48/ILcmIDtNLF
8Ki0Hx4JAeUinSRHqgQR12LMGToivlZtpNgieLjc8ZlT6ub1mYzAwHwcruSAE/sy
LRESZUMokZ+J1ypC8E9FPW1pkP7g2SMHaWpuliQVNLpsNRDQdpvll7/y8S2fBbdJ
IdZmGIXZ4gQLO5IMTc18CchFTxtEeyuIFET1N/sTvdW/aXqGM2SjnKr4QP3zHjrT
H7nHSaeMS3hgSlMl4ydgUbqbLex3+ki1KxH3WoLZhVibLkrLrW+o+IFu8B4QflVW
nvXyk9CECKynlwNh660AfB6CxjwK4YnfJ+eJRnxApRcRDv42W/w8RpZ7JHe4vPY2
8EFKrbkuCaz0bYLNxS5y7lD8x/NeRG1NKyxHBprZNMgieruQWaorEvg5f0giyzKF
y4mKyYzbZOpxsDY2VRXMuM7djVarHoLfsxaJ75GMBwZC6OLWXpeO/3FhSSAVxOLx
VCbqcEq9XslITg6eilmopStD25H1NErBT5lz5PRpThpvaw1d0PdnAsczUMfqOae2
b4Qbibr4X1kfN6obwdKknQ7IUUTuVxxyRIu0PRMaQZ6ot1MGlea7KLBb5yyleCkl
IW/Qw4VidAlYcMlA7zgYKN7/1KzfOvrVYCPqvf9/ZN3T8BPuF7FcmQG/wi9uH7iw
u3cN54ztt9ZtYn7v398BZbs4NoDnKNzRGJTVPWWSoPEI3zrOWxnlZ19zhA5nsgVW
V7CMA+9HlRIUy38Db5P2Rmp7r+tzIZ9AmFOeFWQCJA0CSJz89BEMUTY6HItEEl2E
hRYjSgZJjC3NeP46O1K87VeBlWb8GbQMmlTiHyvTXEL21Iz/Wad2O+bpNsYCx2sJ
1X1+/hDugDlN5deg54MeyAtfnALF+2QmsXJ8QzWZYxWKghWM+3QMguIrP/8Wb27r
RPiAYVB8UZuuXFmklfpVS4IQVilGDJM2lH+ip43LRP//5HOz3tfxJhx+R2zCzaCM
zN/hwaydbTSdXcO0rFpkrLqIlUIkumxAiiKolMitPCq7Uh2sNz53p9NQICAW10/W
PrvrW3TndLjzQqs5F+W98UTssaYKIYSEnUeI5QMI2upcZdGG9nC2mLXq/SyCev1W
bODK/RmDedLaip5aw6F9co7x9gzH6XOplqSAszH725C+4nXd5r8mbXCOHBXToyiI
KYKfCZfuF4PXMP7jeif0KhXtnPUZXHpX+c67VTD+mj5mX8Y4Mbf06UEETEiPZClc
7G6Dv5f/JfCs1mGA2f1n8CZBjb8GyqPzI3tDwibYjPEEccE0VfRwhynQHPwp2YUy
ohQoX6MgQDjK5Sh9NkO6hsTxyzXT6lYjCWYnYBbJkARLPDxWAx3EBXITMoam5Yjx
lDo+cJagMWCI+dlpzhSz4+HyFAqFjfEHpuj6XF6g5PkjZ3js9bpFJ51H3WBi0guY
WVME09S/T4JtpYY1qDxoRApTCDVZl6Ih3rJ95w9rMfJCTMptCLnDDjTvwtlmXrxC
lLNfmRD+tposj6nA7OBo8ZViosdzLvxpxDQQbySw91EMPcx8eTzfLO3bV+wq4cqU
nllXk79EnSgGtbrgNGWdC1L2w7QJl0get+NBo+2PoxPDFsr2cOmBHdQ2mCyLHBDo
8S9NIZcjftyV6nMYpqzKvQ5iWq1cppHC4K4c0BSY/IgBiS3GMxAiT9hsNfMU7jZ0
lUJt9ClGnrn2zh62X/tUYvWBx4SrtlxTrgtP3xdsWnTyw/MyhKPGlnP7Fs7ZKxkp
QHqhecZ3USyTEuhfdBhdEAHakQWQIfgLMhBYO2//65JsigqP5Y3O53RPdWmZfO/h
mXr02V/sg8pW/YylfnkTxKgQIgJM2sjgw1Z3jt9eBSqNri3mCwJ5U4vTQv6TfG0V
/Hm3FR2SAX9mChBSa1B6hRWbopMmGsI38KDKcsVi1UA9X0o6xZV9hOclFfPLcqb9
ioUKY33yzOyaIkv92lQpSLvuFjNDEbFzGtyBfIyhMfiO/NkOeIn4iAPEfwQfjs2w
zMoyQzvVItgImdQItZGIrIUR5t3EreAx1l1JTEmhetdFm5pg6KmO6yuQZJtEGjpH
ppq/NlXwnxBpa5u0QsIEQO6vJ6zrRt9pfEWg+p1JBmcM37J2QbbW8WYoiq1T+xWL
o29p1qIut9FTjR12nXNYhDwjrhb5D7TKkyZhUEh+wjhNPNEy4qH1Xkrb1e4qCu/P
sLuKHEgW2q3Qf8S16ClNaNk49076TL7LHA8/bg0xTxCWn932rHT//A2ZaN4YWqKK
QuOdUh9OBQBSEMG2L5UZYkDh1ZQ1pAZQyITwWoUydIyQ1ue/d8bHj6jem3RNeMC5
ACBlvU+k1hekQmupl0swDphkROICTMgpYakzRaft1zglgeEXMsLZE5xPq6/YcCCW
0pANCz6SGQ9t73UOHYC2rdzO9n1QDh3s+p//yq5Fo222upNp5I+KvVeqTtnS12Zg
BOcowZJu/8PnZrJn3DpdTkUmMl+XBYFzZ/b0TlrynITUY5TYPETD6qCpOR7micrb
zrl0yQZO+Gzo1kk0EjO+Cd5I5UsDykqCku4A49+Wce7gnCVfAiyY/HdHIognx0+6
sR42/qlHGHs2M7InAVLy42ZezdJDWqNN3sMnzyCUPZlSdU429w5zoqSrMdf915HH
SLaKsBe4Dy0FNirIb9gUcMcWQd9VkWgfcdVXlu7PUpihhgzEh/xKI9s8WUL90Yj2
GbESiwiRb/PFSEh7eOLERftd5m8cWAp3VnrhUMsmlW1tXtGOFGQ0ZocqnLn1pbLF
x48fETsnfcnynoDcNCWvhSpM1zin0zSlb9cxW+L/D9BbL1zvwMFaNkIOEA9LMB9s
0wnQTYA/gRueSfqG3acI+bm+jGjhHR7piWmYaK/5VNobKWKFdnxHSh/iZhghiO3e
+ELrzXaUlI1KBBwhjxAgXUH/P2E1TrbEOMFQNO7kgDw7rfUfJrW4bKVZWHE2g+2/
h7OsBSd7M2/sPfGWNB5CGBOMm2vxwIPq3I+1ho5UWfegqkaYwhURoHeJoHJq2kDm
q6Le+3re/SsqVdOkbaQPODIbircxfb0a5wpE6N05X+Q+C1VXPP6J7SpKzHzxp14h
t50rhQM8Slo+M7mPQHd6EaLrfoL4eVuGNnANCRou2geYT65uVNCLKPRmdDI5FRkc
06cwq+MrUi9s/QG6rjREb5NiUZoVaV+ZHrO7FrJW7hrLQYJzAhi6IQ42PgPUaGl9
MHLlA0rWt+01SWi+hH1xPas71G3m9/BTmajL0CjDRv3J4rdKN7hCuh5ZTTR4Oj8i
yZc2HTmgAm8msnjt2UHTEiMaEQqop5sCbisnT9+V/YNS5dqhghwoNeAN2+Qtw+AQ
CwaIoBQtViWPXAw3SvlRdCZtjXqEmHm67Wts/78EqPhkdhiqduW0Tky2t8e9lCjA
lmia0WGzojxaYdiUZfJN37/3PoeheGEU0xlJnM1k4nooTAIftvYuqPVjBBIZA36n
8lYDvwFFM5dboH1YLTn6yx5vt3rOA5XkUF7wQqZvZCN8BRA8eHkiF00Icl4DGz21
muMKAubYknpGdXUYoUT+LNGvh2wzqAW9EZcdikVY2XognPVYPdURPN7jxEncQG4c
ipj0FLNJx9G0bARulEltdEkJSNd5aDMyxQQ9+VJAhzXbObo3gpT9XZv1IIrNfvWr
CJzIvXjqwhXK2MRqLfBXBeALlCOHtgKPR+NawXb8Xfyopi3ZqcpsyUDj6WuSEfOl
ZGm196Vi1yLf+1BxKT+lHk4KXjdRphyGgV/DNxIskSkuRcXtYVkZZh1WWgmvJ8Vp
p42K4kyqjs6bFWAzh1YURJEu/bHYF1BKKLQhYL8bZXZKyCBqZS2KWA182x7vjIeo
kXiCK/4ynGzsUiPnyt6uQa4m+zFhaBLaTZNreGUE1nOW993vQyJXwdh7Ofld9Ghu
oYQR0vMlXAXJGekW9kf+i4+YPnv2MDkgjeNh1SPq2kquetIjxljOEAKAig+OdVAc
YSIiwMbxe6ejcaJBBNzQst5Ed4986r5gUhCSWRj0iay1iGBf/w/v2p4f62qM3nyf
iVNBFfWaY8Ftyj+vZUwXO+bMmNDd4oFvJJY4dsI+OZL/TmKGTtU9ELFyRFw6eftf
kMfG/SySUlpu2XWKc3N7nquyadPyiD5nbntlpeg1wNtFPi0jxb3dnEyKb7T9WsN4
blusC7P6JwDgaCOAxO7X+m/VZKpsFKSCG7I9xcs330UvI/dtf/jwyQEqFottHXLe
MxFTEZnFrLcBs7uLRHvfCA0R4C4N1hSYZI77a1ODpC404rzFuVCpECOKQ4KI13I3
KdzESPB3myc6q6UdtN1/T31K1SiYrVG20acIU9zZVYlBlkxNaI5cuZpSZsXxjI4D
SwYVwWIxDMgF2/ON7Txap0JDSvTTP/+g8OILPJQVC0d1qPqikSTEfCdXMvSgWtkM
hFlgK8vealSiRAvM6w/aeidmA0xv0PA/mqv9O8XMFHssQUiRh8DDu8n+6utE2ox4
W+IFJmCMy11XXNNQ5MrgT6Zujnp8x2NQDrtJtz/tEeS93Wn8JUaZQJSNVwGrvOII
3iiGwF2DzA6NmP+879Me7SDNDQoZVBiJw0idZH2yBsOsMo0E0BbJ9YIXvPpxp422
/ZujN0H7uwmX9Z4dFK/R2SVWgDeUV5Y+YIfZdlZxd+M3pSMyKbLLNg0CGtoR8nW9
bUq0ZGGAKmK80pb9PLIXIfMucjj9tP42aWfr9EJJ40UxoqdcaTSzzc8e2d76bqoa
bHjEMNZ4wZNzeBakDHXPr/pucFoLmpWYozgUrU3oGnIglgAPTte8e9pIPSmgtZIA
YH2w4lNsvMq8FwryMes3nxQ2OcnJyF4N9beI0Pao+/XEsblCaxJAPsCC6HigdJH0
4PDMlyeTlBz51khz99DjBfkRfllPJDuFrM14YknJJIAqcQNNgKenlt+9J0Q8EaIg
nPUDkTESEkx2BDQGg6z+Wtn4+elGkr7FjQTe3jGRSJRBvO/863SeciGHS5kCJiok
yCt80x+5mR1PkyF3JCyO2oJIg8yE44HiERLyMp0jJn1XvSQNKneF48Gb9AykJyrL
DMghA73HsjNa3ncOTpZO4aY8gIMwlquvW4vaR5Js1nigljNc1GRr+76mtDvtmnb3
2TdIAp9v/HOWd8toar0q5LDi7GJxSJfkt+uNdmO2oLPpTsDVh7BluDYdM/GieBKR
UgToS9ksx+7L533Roil3BQDc48rILeQvm9zwncYlA79YuEsqkDwwFXfZJ1ga35Dy
VXHZAbQZE6jXDidQ5D0337nD4MnsdEPMPgasl2HesuUL3dnhukLQrcpISGZgQXxR
o8uA+bEeJgstdUd5vfphvGK5P4k83DGAl/c5vLOBBTy5X2f77/bVcCRNMR06JMiM
Gq08UaUa5K1bNYGrV+2givZZzl9bUnaaIQWvhmFcJM7ZIyXyoOahyYIGSoGQM4X7
Yl8h1hYYVTAjjJaKKoXAzO2twiPRFM3SeGLUK2kmzhWFEAdIvq1nKvscdYqCu4WV
TG43ONHbrf2GUGlN3rYZqb2tXMUPYq5f1On5mgsqSF1rcQX2vYskBjYHaDm2rqAi
e9NTnaJzSdR2qfwdKTJHmoHtI0oBaJIRHcwn4Vb66R0kGmTicFS0w7SzdoxdTEoL
+JuQRGD/UaaaUsKlDhtV2ex4wZpaENcihXtkkf3pFoJtlMdh3mwtMQPzYVILq6ek
nnPLU6fP2Khkse+ISX60KL+8YGwBN0llyJjl35AHpYgXWJQNlIT7TY1sLhaWRpRQ
Z/eQ5K1/JkJDc1PNC+WF/Gn/7SuiZCUfeHOoVvqjX9xToqWAoVtnp5n5BdABQVPC
Kx/sb/Mt1rb6es7yQc7ahhabHexAEE/luvNiLLlpgZA6RTF5uOs5rFqXg3vJaARU
SH2zBG4jNMFMWx9P1sHtN5TFB1pooG6F54OsiIE+gE453t3g1MF4DAucItKgw7Un
KCI0URmILaQpItWrCMxHpfbIRSImwEjrTk+wWTSX0wUQpQdnb+rukq8z/1KpAFql
r57fg7iJ5YuCStLi1KpnC7QncM5O7LGI2yJtaqBFxCgGZ3Y1CNnc7deeSXwmPIRC
/CUo2sOOvRrFuQqldDm4tiE08Lr6UfepQKLIlHmSBQbPzT3AHECdaOjizdIDSxkI
CRc5KtolS1DL6mJqLDnbp67d4lScticaFs5YLS6iYnjG1X4KmBGBpN6O6s+D1gg1
Q1iB1q2peco5YmFoeQkIjl917q6A9CBeRU24VdHFhEOoXN3hdu2KIBhicSuI5quY
8o0IuHOvvdbOkgBnQwhIT6xqO+G5Mi2tNcMDLwgNns3N7Fw497ClZTLD6oKpmL7V
5pjih0IRWCT8S0TzOUqHm726z/jZyufd497QKFDsYDbuCodwQnx0fh1Q1bpCLxpd
EPSho+Bdu+ChQQYUsPqseyE4tZZO0Rec+p8t4oZNJX+A46ngZv8gBShdRM7tyKXi
tXXo8Tvu51Dy/F0lD/1TD6i0zjd0tCkG8d+QmdMT7U8VWXQ1j8T43YdxBBveWMQ1
+pNasJinNoXMESohKMtR/ZPnmhZCwipTXy5RMBD6aBChe1AYycg8OXGkTOp5plRA
EiP9YwtgiJNVEj8lTQ2YXKoSb0vwjA0767pIKPRc4G8tCn7GTgg0MEm3UxzbRqW6
gYuN5HFp5LSrPkiWHVx+2svTQc+KbPIttwOmjKcy/OblTd4otxtXLZ8kqK/PzwY0
i12j/dVx/+1iM9i7wXwDzoJ79Jf+I9dzWHZvRztqUYOagqiujSRI5brvViy6IpMW
dYBT/gxp6t2sAuS04ROzS3sSAkzdRxF87EW/S+6B80FHKZWtRrEdeP5dd/Ffxu2U
rS+WTEOnOndeR7+qnb4NS2vVcGUBayFFsxTpX2GBBIBgImegRoCCyRqcGbz8vDWU
bQIDP1l5KBcmCy67Y+i3cx+10hvo8EItuwSVMVuEWYzOipTHvA0OY78fA2+4n9ul
9HkikbsPAIEm6BEKEO2R53U+2ENSIgIAO4Ub3+pB8XEumBwsNwzXIa95o9KZKXOS
fCLaCRVeM8Cys+QXXpr2+FixyzT2zr1k2isMGDy/FjzFizYkBqgL8x5p+l5AQWZL
7eItdB1Vi5T0d0b5DszzI6gAyU3ky1EcpEh6zjaAayOrcZoAjp3KBxfwqggRE9dO
Su6r2kPPv02yernjwMCWOs29UfgTNH87aRs25ieTLFfDpOeRpb4jmL9o2pRo2m38
GbvzLoIadx+dgWI0tUXfbc2YqVaJYsRCbUAtl2CqSY+smrbS23/k3lFa6z7th4Y1
SasXfv4mm+NprDm79VKYbtWQpxSrMQsaDI4s59nCq/wN6TnBxVOHqNkxiPKPsGI0
hwmorMorBBU8BeINeX5wF4uEUU7aKBV++7HjSbarFKQ7Zmr439MMlzsJeiI2ZEmq
0l4H6DkcHRhRRUCnlTr7My776IIdtoSbKwQRZvUyt+UlbWMRRTXUghwAUqc91gch
I1rDM1pS6BnD1o7ZIESmsEx6UdWfjkXA8y8WAdWistNYjb2wWz+hcckjpHP5HYo6
MQ+uFWHfyikJK3r2VKY3UDgvG39zRBcx/76O0+XXbDCv3y5ZiZVjePwK5rnjnooo
ysJBmbSgHCqdAcRPYO45ndwmxAn8ybD2Lp8Ny5RlXD/BN2Zj32zPGGh+MYxQjSBq
f76LuNDHOf0joY+vWMmymoybJLOP3kPq7BB5zSW9mS754yrkYb8e7USq+8N4AkkG
rFvUZn3aNcrTgiLCs1pN3/MM0CqiPcCuSaWrWp4wVhEd6gOLZx4qE3sn6XMaN2Zc
amNOQg91U5IfwyoC4Z60A8A/mZCMHOm1+gJCuLvsB/BYWn1Y3Skm2VhMpQEzji+J
s6O2XqA/mkYKN35h6jaXfHuPTX5Bg5btS1MS/eBnNPLJNsjIzr1wSWwpVVSg+vRG
WVjeBAsNpXQmPIXZtkwSPak+TzJP6AOmTN75Vu+wBFSoIEJRZ2yWdR//a5A36W+c
OTaAy9UxASw45Osf1rNJnSf52znqn0E6cTHMVcn59RQItI6V96/JP+uA0AsQpMSQ
jrGyEpzlfJ5ACjjOsmymg8Y8/7ft2NxfvyBdOd5+v2Xs5kbMeBIjICNNzEAY8Kwt
YKsfWoyyaH0Ml4YaJDx5nLY2qYWa3HsbObDKwUEjjYrgx1NyxFUv2tljiNUw2V69
jF2EH6zWiBnzFG/95+pXr9PMehOInxZObMEUxa/OIPTXchAazIQOpFDMgCYWDW4p
HuvWpLYsdObE+BwyxTZzVqfm4EHLc1YHRNI7w0huSouo26mmkmZVQ+4Gg67sOA8Y
BmqmF4aaDFqNwk1sD1DFCGns3uqOsGd4E2CPJpR9MAkFCVe2x2p3CIAJ6xbKAC5D
hU5hSY51Q2s8sDL49d+4oe9Tspm156D3eKsjC9i2iljCLdbNWeUthxPGYo3COMQi
9LwN6TLGuA9LMIcnyfekhVUTtXy3oOshmcELf7dsWfymFYkZoe6Ol7ZKLPEDVWGL
c0l+jJHq6DAbErDhzEYAW06oGGqdZM5qMGipt/EDhYLYx85VPkuWW6fDZpxJgrE0
/VS8LzxwawCVVk1b3p+mRUuN40ot8/GPgFapQQChzBxrosfNg4x/Oe6XrXXWsynd
sQZKfoz9BWhh96Aw1o+BaL6SDyAqaFKKgxw53ptGNb+F499tBOqXmSLUOe/3apsO
zF3bjp3q3I1tO3gFSdFupnFYr7eym1hYrmSeqGzu/fZIqNlNJDnwky5f1NgyYckk
1v3BSRY3oYwNE4s6iTtKoDAb3R88LfZEuyUEjQXLymL6cCnkaZW44MoFCsnddsFG
rsJofpEOiQZ1wi9jLsRZJwzRkvN3l8+LuIRV/EJBwRAZvwFPmPda0PKpwrfcRWOx
jktfOh7PpfmKrEU+t0pnDx7X+CxA9k9V74kJ+SARoRbPHXWDGXADEjQ90OWI65Nh
16LRt0OQGrAEreO38BIikfjMm4jxrSeePJ1MF4CeCrVamlk5gUS44og13xgmnDBW
W/JxBDOdgQaARNwmT9Xz/mMtJ2v8Iv8SOBfm/F3HuJJgXraEosEyRUYeUxNQVvFg
36dM8rcZ+pr4shIGKO4DfhGB+TZAnzp3qZtbt0g7xcoNRRooBVCYFmQs1KwY/bjV
ttuO5mTbdKnJyW54ItvA4KXuhfgM2bK6kYrcA0PUtIsx+332vI1gMEk/mhCaVBBi
XxkByJEqM1F9pnM/70ctD0v44a9/ROHZXECaYVALbPmkB08/zlg7rfrLia8xJB8h
90/ktnZ7FRu2F64cBoyNDVCK3VKAGmjigvpx07aEe8vbYJaMTlOa4AApQQQ7v+tn
Uzq/KqdkgPJr2AVgl5sqprCBF5BZuZjwN2yyxVNEcfEXlXJ5n4Q5DLEOHW0bJDM4
z0fA7AdUovUb0qaHKQA2YHQhCJqVgQyWxUxvw6nEofk+vtBN+wEmsy7/28ysiOMJ
yywPENZLwU+Mp3kt1MhJniUHBCMglR9burkszHp55nrV4sfUF3bfvw766MxNqD/E
9PBU2Q9C9huy99JopDWxv2FXLsXOl4mQVtQ8xAq1nLMqRCduQ2Id2+HY4ZkKz3S8
3bdiMyrhKJqxmkGthR5O0sHfgorXLDm6ZvTu/Ax4mMZ0y/t5P1s9Hss3YGks/U6z
TJxj2dzT5FEtyNZZX+TZc2/M1nnkbKYWEaMaIIvkWyoZueI5SIqU14zPGjuWtoC2
cFFzW6h+2M74ksSBo4wAh5+0ugvfjdE6dhBY+Ddybx6uDzh9UB1iVkHaZKKcP8Xy
kSKKZSl0fxiAktLUIF7dXpfCOmdcImE/LmRFHRrRtrE7KteF0xGBO3NQYgLUDCfw
tHIwPGTqFvTfN9Qn9DU4GvXIS+kRQl95gX8fJ4G8dqr2oBwP6AXraKO51AXdIVy1
1UupemOoKE4t27QYAnslQ0NHhexmG0TpKQK7ujJX5u4k03Mum3JylF4Va5Es7jgD
qxoa7qU/i6pBY8JrmTTSjaBiKF0CjN3LSHrGMMX9rSFH0oXTgAK99Fxz6gDBhfex
wnYZokj29+A6mSTn2YyehG1G7OPqbDlrVtTZJ4U4X9sEC+bqT8QYAV0io3r+tU5U
timI3uNQfidVBvbOh0ZG1TBkSt/aUc9FlZ6m4DoRbd/6sFc1NQuTuiJ6X1jU0xWn
23Ul97MbZkfYm9MwBqhefu0u5xUyYmUWBJNDio0sp5t1BYEEq9F9H7r/rrxM0v/q
YxQIbnYpaZl8uRkIbncGama5kIq27MyGRvczMQqtlCMA6/31IoiHEUjiSIy3zFE7
rexC8TdXUbBR0jOXTl4oM3Y/CCm9YCKrOc697scWTGGYSixUzYhanx/qQCaJjwxe
+0vWNzf7Z7olvMrwEwdfkpBgOxmap3xtARAORX9wWhaSrbVjzgifzC28rLW7BjQl
vxQxWXkWBxEtzXIqd6JQ+Yv/6UHlSG7OHyA3rGronnTZBk1W9/FkjtQTdLwF8Z9Z
Nt5asSZtioY9vJYDdGRAtDAyPjR1GLLDIBFQyrzQpbwVb849myD6DPt2D2Usskff
YfrFa6OCsFY04dIhgogZaj4L9zSXELZRlYlEeZyAZNrmgyK5KFNoFjkqDn02VdNx
PFmFhkwdNMHbovikt0qbCAkQnP68EYnOXWuJH887nOyJC3Uzoz8xXbRqXcJXEwCJ
S3LEpC27WTfncp8gvpW85ycWb1x267XU3y2POcA1yHZtiqBUcuBoGV0Lm0TUuTkV
/3mSB7JxWF3plZthJ8mLEBHh5donoKQTifN84P7Cj5pUx+U93f0XwDhXySwsxdm1
5pdnRc5jB8KQ9SIDQ5Wlkg5Hus0qLnYHLvwA8X0+uOeLvTSgaNu/ViLHCHo/cAAb
QN2GdRaKmmGhbu7VC6sbN8RVNi7IfEzEzk95FDYcfSDKbFwxLLq8Otny8lcusK0y
hclo5hR+6HxN4ol9kz+WFFEuCoOyOgqU3wzv5NEnq+nmNoK5oT9/ldE/qqfAL8De
rJu4MNwdvxvzPqnKnsOcNggYUxNdGYzRJNdTJDVzsEG97+72SiPWm5Kc8cyOivcr
D9xAKHaWVE3AltilZALBXKBUqoYaTMNCMe3eOaJrOdRDu3TSvi+VnfCV712g/wM8
zBOEb7FV0p5EFmRt95j/cfSA2yaDjpw7CqZXMBFrXl7YdnaSiSR2XmK8J3GWr/Qx
O/Bnfooq5C6PRuxotHsfUv7MVq+Iec5Kkq/QkjAlQdbMs2G7HKXI5OaEdZIuQpND
O0qpoBjxjnymGRif0mZlxTFmdRtCD8XKwGrWd27dHgIa6+LlINPGQ0X8VJSPjfn8
4oALt5jGHxHu8tKTaEhJheMU6kvrTtk8x0kL2rj3O7js6Xav2UYAKi4576kum9yj
Z9QSrYEe9CgNvmkS+xVjt4ju02K1FFFZctJbh147KxNyfszmWgVutKvgbDGa7do9
dogGpKwwIk+pcLAoT/aUzByOilNzVl2t2CyjYUOlLgs3gFo2VM7Fm4+Le/HM/I+s
CH1sYkvxwVfWWlrlSZ3mg2tdOkD63R+sjXwz3KcCFqbg1vLca+9nGWsOyPpOdrdg
g/O7sq0/WxYV2OtU8/Cf3UlG2vP/ytz+mmHzWpP6UBk8ofQPUqOT+48kb/AApu8b
Wxs3KylALVTPnCBkGFRlCwLaGn+Fr4CkUgWd8A7po7ARGQGNcCqvl1/IchK2MDfR
a1TQPqescTGW640HjR1nqq94JAacE/Kvi19fm+ijFkbDi3EjdLLzafOU4XQrNe0m
gJtBjiLHWXio6r0QLFAkjELzxJMaXsfMDZR8w+Lyhd1XJMvu0lsOx+971dDVpn+a
2PUSMM6nFyDdz0TXR0Ic9y0sw1DpiAtiwx/BXKe+Q7IDHZGEthyl1lWorZQ2Mqk3
NaL4XupVp2FOjZzACWUrkjOeqnsSa1ids+1+OVCi837GYHn36er9IGEOZ0Hh5PV3
tLDLRPIua5eRuoKiwxkjtOqU7Sbw4tWXS7+LQemLoBJvAggNC5IKzniuiwLxKzF/
TD9dMvPVeQ6JNT7phNz2RGJLTrqCGWmkGevcr6h9ydKJfCMVik/FKHigyqNCCB58
2YmH1NagVFw4hA9/DFSw64oF30dsET0409ZNgiQzKR0z5UhQLXRtWSrq4zAFkUSM
XB0DhkxXqq5H97qj/Xl5KS2/ePqvwlikj9VtTMFMfjfMqGiyCDto3Ll2wCWLNJ6G
ly9Wwg/bh+wSCuY7WzvchOts76zhhDzW3giniql+OZLSqjIRRrxJ2N+7UfmOOouD
IG9K+vBDrNN/relyIwCwNNZbsKqVqejVvoiqpZ7quWKs/XifLvC/32SJm1/nsGte
CbjdUHaF3PzHIgWpQmr1CyOlkItB7zvBa/0MkFU//GtgdzqnWd0w06tP2OgWWeP6
0RdG6+mp8lzViJhf9TOFc1wol6MUjb44SMF2DzG9CFIypPmrFqR60JCOojd9mURY
3xQ8c0YLCU6KM8QlPdQekncXtT8YJ9LwhUfcaNQSeBQv16JmTPUygAdZfyykhbjj
wpNC3mDjFse4Ldw6kidSdFJi/JYXOdJ4iMvCeHHd1sHsHWEMj21BniqTuR8EfB9Z
NtLBvq4SACazdqRsHMWgtf9vCBK9fXqqaHQrhHNIL5LjuCDoJTn5zb9M0Un4oI58
/fLh6ZgWoLC007jmZkPWO/WMNz/MpYBkdRIAH1AKf4TgMmhAzzVXDjOi0JDLm+4l
CBd/yNT3cuZWdOb1evoIkGLJ7ScKAeCEBGG4pjYA1wsbuaLURKQ1k4z6kAVTCwDI
MJoq7qA83fK3f8j7wyHXjdAxgAn20izIwZJGyGuQkDybu26xviESFeaaw5RAJ5m4
of+X4OKS0XvL1gQoa03/hzjx/zU/hfxD5D52a2/GKiNAoXnPtaUcVT0vrc7++rpD
iT+rphVR6d+snqXGKH/HNQspe28CjlvFIkS8cKKrPFWQWoXmpgkuS6Fx8QbLVT26
8qjp3axCihtqjvXg5gdyf28eA1aMCwlRDlmqZL3tNLZ9YatARpNt0CcaFdY2c6Su
IGPDw2yD+Wy2xDnpSAUy5PFBZH0dAPurzLkX144VepvIsoyf3xsYshIJeb/HQ8iU
BgEMtIv2GfwVZzS37GNU5n60uiOe4GPtCh14PDC9ZcRxBNnqQ6qAYkFUgv9Ochzw
ZIfMmjD8Cwi+SnuY+thV3fKEOY6zdNXDmQIM4AQyYQMznnrsaLBbzDm4anKu8QMn
Udg8Nj8a5mzkI5IjkbDJUxVwKXD05zn2zBIICyXomUIe3H+5f3Yh092tGgrcIvau
JJuAHuFlwzQpPO0RPisvT2KGAJ+fbR1KjZOzRfZj8LM8h4awzvKariMHSVtlwJEe
zwqShqd3jjC/3jtunE9QQW2MvsJR1WITBjqTgvOCP75gjHgwtO/+VFagu1QD/Xfp
AAssQzXLm65LOFT18qMovHnzN+UnKdZUS3ap69yJiiweRcEsncs9aUEhSfDL3uHi
4m7E0Sa4Jp060ZO+LrkBce5xUSS/0eOc2hThv5kz0V19TSPTqMvinJsrdnZTSOc9
x+xoHn8RJ580Adyiylm3nbBlUd6aSVhYxCHiyUw/vWR0xD81Uo52ikq/+tL0WG/z
pGDtN2Tjf5z137Z/dbJifaXyL7pwmFcJaXrA8WTVCtceJONcmRk2kxvrm/scQIWF
F9/jLN2DziRzdAVfah/uHqUxouOE0BAEV+wit1JvJxIlXKqX+TkGdZEKu/2Zsbdg
vQjIxO8HClBk6KVA9Na5ZUk0CMEdWpq/ObAB8eiktvzgFvVeBbWT/mOM+k7rH4Kt
Xq18q/9NtQ3+05Ast2M+dg7K8pqd5+0VNFpGYK6gmG7HJ6OighAydd5Yb/ha3p3g
vTu2ij9jdv8yaPZAQpdyIZBRYeXLVq760HZMsWJQLZgH5Tu6EKQnb1IiBcP06HqH
vAqnl5r4Ch9FkohpDcX5fasONQGtvWrScgWYVUk89VCh5KtzFaLpBRC0WtbEDdqY
Ni26Mx/owsQkqspZfa2myyb09n1PgE8GmVA6Ur+dgCBwRZX8n4ebM6ZKJ4dQoqJY
JGJ7ruXKE6dCdESp+GY+rB0NF6umJxRryZvTiMteb/TRWxwrdIRPhzbUseHO6AAH
lRWxJfyKici30orvnnPFhO1WSEn+cyV64nagn6i1o7APcTM/h3VZDC57wUKMWh/6
lZi7nsewU9RbLfu1B5kw6SdgrTqac6fFDuve+Jb7p9Vzn30nxksTWxUbviGdtPPS
2ckchaJ4cbl3HuRufGbsQEj0R8/3vzcZKC/kEDFQSobIGqAOilUk1uCa6C6clvxz
2qRDu0ydnzD/5W9/YqJiPU/WNRbz3NnbDJeP9k8gc5KbwXKg7CGXgd1efV4rvBCw
KvZLU3GSBik0SI8oEColDNuk9D5Tt0jmIWG2FDxiVdph1SMSZ7txaIK9lsTLpAgL
73BVJpSVyS7UAI61rEfKU0AQeilmRYXWMnsKsZ7ziwWWUdDjzDq6BSGtvq1zPuq9
YUIgBUF2c8BprvSeR4dHLhFcJzskl+Q/PLbDdywy6/rtkQ22eEZsNenrK0XvnLFy
FjK/UET3NIRWQyFbum1ZsF+Mc6ypx0VqbETZYDTxYqgy+OKxOZCZq0z7PwOmGIsn
EkwMuX0X9VQLPA814/sOixwpDenyCdzPa/VNcXtwtmlPEmXf3mjEjXdyWZAYU0lu
K2IsaLArzzZHaHTLI+WKc3suxjSxasyc7bbCsAEQ5DuCtKQWb8f0+a6k8GFOeXnp
naPN9dpI3k0XTtiXU2Pwxm6pwsAmM79bEKRO2KZBeiBXKQgVaSgmRxFbgyJR4DTx
D/MCNxh13XB5Z1w0Qq5LVvWV/NlPv3oi8iWFgoISknY/br6ecfJe2ieakmuy1oiS
R3hLGlmptlLYVbDsiPbHYpUDwrajGbtYJ9S0+xN19KGZksLFiNFnYvu5juw8hfPi
770rLCMCDH2LFPN6upPTK0viRmMfFvpY97591WajvHb6pKAqQ8P9aXQ2fFjW8sIb
2EXfi5ReULJhYe7qSSmsSS/iSDDD7MzZuNvVfV8R/ij+eD9gGjdA5mbM86f8T61N
cFT9iyYXx/EaI/md7GBwQkftjonv8up4n3jvRo8TSbTRcr2yVrYsB4gpmy1Q4k40
ncHRZrXG7dKuWWuJBEnjJRvEOklowxzxtY21OG7EVZxHXSDNkFqfZz8tejzYrZq6
BBEdWy2Nknrro7/LVr0Neme59gjCq2PjTDwv770zBoUGgZy6D0J+Qhy/wfU/QXC7
+Xt6V9utoTLWKKCLfwlNhvwzpYeX1D9RLyrfc9m5iLY7B8wUIqsnkCww+eJOP/JI
yrgKCiQ6hQnjtmOk2Ol3mXmVQeIphCWedgiIOQi4u73RDFSLIL/yofB1zHEzGWBS
v2z1p3ZfSdTaEmu8JUB+3AuIp5Zq/e7Guky3VkrUXxJyvqmMB6cEAEHacbKmGpv8
cLoTvbqorCS7RFj2VoLr4bhhpo8xeeNe3r0XKGQabB35oXjFoo4IKPRKRKpbnyRE
DVHhjXwWeaOEEsLCY8gL0VDCPQfSuVBHNq4r9dQ6lgeA9RAxIAXDrezfPxkrXIz1
QUxGY4LURn4ueUku7aXt5rSJIioOiMNUMxHHGhRXnngd1vh/iPYEJdlqR4tqFz3g
9uAf2Ro+VTiF+6xgN04B9cx23LJw3tnH5cjtsdR2v/r1ynYdeuiBoNLxNLB5atPu
1bUWyMiLJq/hIo3PX1+ScWpO0KKsEpv2WjrXVVeS0Zmt+k4LDs+URAJzTrHqCtfV
4KSmq7H/mtc2T53Jzzd5P6Rm7theKBWGUcH55rBe9TRY9dmUfcGgHJTxB99MFgzH
XDqkywB6zxXDAn+zVICTGib6+1Gqb/ibwNf4qacvyEQavYfN9N1CQBlSxGDlzaeL
+H3eYdiMIsg07hk6BAfm7m4DccZmrp5bcnuQuTfotK+2E4AyMOLoCLf6fsI4yelI
EKdB+yq2sY5blFunmkN6ftlqsZcA9a6z/IUocdywOoS0feXfhS+wI35jsDykckUE
88I57SXf962G1Muh1L/ob3faOCM3PMUzOeuUmPkfpSy9i5sQU+YbTfTQu5NRB5UM
bopE1mLyiA/jw3rmBgkuqMoqSQMzUYMY27DcmozNOw3dsP4AsRtDZbNVfPqCeK0k
sqQXygtLQAD8+Ha37EYLCiv0pxEQvllDQ1MarJ4N/P99omid3kpOtbXRiYZ3RgTw
zJIELL/WDj4rg3VmeZogCEKQJXE8xnGdlthROGXOyZ8czdf7Zw5dArG86Nxii/xK
pcnyraQoCN0TAcheVT6ACy2V+nFKdbTRjdfy3a59AfBttCW6/HmGSA6UTNlbU7Yj
N0hjccGjPA/jR+V6LK9MAD37tPQqGc++aoP2Yb4Tf+09yvCNK62TBZwccdca3QTi
gOofm5ZSob7FOWPH2KuLjwRkqJooqZrAIoCLdUUwgvf4bFi/xgd/GZqTcjizn7ts
g3oUd6Ado6NvvlIPd3Nf/BCwLlWdfYOLcyAWVQyH8vn/yZFgJ8lz4nDbtWYyMj5+
E6UxLiS0n1MmFerW8CESnh/MP32LneWCgZUy5svPGEkYm+qv4DPSwZmpyEf1czbh
bs6yAs2x9LlMnAxo6f9aN0s4IQBR/ws84mCzOehSdgb3ZgHS7meNPO7Bbvk3PAAn
/uGcnd/IEYVpkLFRHFs7BPe9kPsxnXZRlE73HQi9o1nZux/Am4x5xeZwGJq6uqMK
FmMobJLtAoxmAR0dFTHWqM87G4OYRTXHRtfyAp10zzyKgwoQ3oztLHm3SU8+o6cU
0OIlPekS00ueSt6CXH34hii8/qZKbeM56zINHgswsUi1lA7FTxdhVbVgDahidkQR
8T+Vmrk9qli4IsUFKVVf/ZYQZO4Xpj5cbn/aJocaIcoBuHm3psRO1PGi1qmGH7Wq
5fvhlpEIRE49gMofVqyhCWqLo7cM9ndn4CCYeCyLRpm5kawGrEyfBVqRcVS3VXJd
IAnZ9eKQ/eiP621DW+by9YtATtj260WJgZk3ESkio/aiskt8nc7odPczUiTwRnmH
iDSsx5gPFJnRJwZGkSjc4Sj1qPbjbDA0o6SSlIF8KsRt9/SV4XSez9oaaR4bfoVM
iGd/zFUFZH5r1/PuqQtVHJNOpHqFEEeAv9atGob/IvqSH0aGCDJnKxcHKem8id8A
JXkOLYJaKB1mT3zbSdf2r+j8zf89lReJVs6Q41Me792pITr0q2plSd/DMcj4wPCW
l/9RnLcoN6f6vkbrdldDwc98cq36ph92DEUqnyL4Yw0ARPmvrmEGRvU4um+R3X/h
hsnrUvcJhr11Vp588mLOOXyNbroFaO86RMxar1bE/PkymQbeWxry2nFojaOBw8uj
72YecypaEj8cX15oJmDodpk9nMxT+lIDtI1SBadRf0KcGbxqSiErpLyiqz2AAM47
aX1sKUiGC8t8WO87FjI87SHNw0fn9f5kPseUJ3cnzVrNHMISj97huDzd2HH1sjSu
xBXWZL5bMmtdrF6BQ1fMNSVrCaza4y/e9gNR1HWDPpttHJbqKuY8n8B1NFHBpq5x
XXPQgSWSm81bM41ejPNqibSv9cI87nSB3AT+dPd5TMxg4U4DhyKgwpt028jMy6LC
FJ5T6K+wMMlzHPLniy63kbxMnXzbpRRjyNwATHCcjUiQVo2mHa8iiZaRU9XPGkx1
0pC5ZbW2CxrCisSMRYXshyBXeQZm3wx4VBkpDl99XsZrT8K+XnI9o2PgqfpJX69O
6aEAMCTRCKvfcDe40EJigPRNjQb99M7YoJHvGsg5mZvkgVQRErxKNfRI/ekMv12d
cC8c31ByEF+Y7bKvOQmQbC0/OH+pUJFIfseIjLM7L8I2AZclpQAPEjWDG/vMDyLK
XdlVnBx2UDECGws2uq8JIxLXulNHfcbs/rWquYGZY80fcNWnLm7rQ/qQu3JLND3M
mOoX6tiZd2LNDu8ffPigwmEERTbggZTNoMMmzlaGL5vQubQ+48F3iHaTc08S23oJ
i89dYNDmliCR0Q/vnsfrw8xsDJTqdJkaLz722mcazb1iXWFF2eY3BzivyYGvjtTO
LMUOQosev0+vd7GJ59wK6lyrbpqvPDsY4P/L1vcVCA4mo8lUKMs0Z+aXL+GAeuXt
lJtfFhw+u8/0Oq9cpEc7gaD0Vu1K53BQeufZ64Doh9Vs9jUbZObTPtVhAXV6gK0r
7hrlfILfXKN4j1Oy7plk7XmdpbaGYlYGbJLnDbe5z6kVZx57UeuYCVFrKRFtjJEl
tGGAyWDLsSK5t40LN8NVD9oGa13L/fCA/E5wEqQfgeMocSba5I2PQLLhnm1XXlAE
o/JEAPvW2LYF8sC+mq27Oug2n/WA4bjtOT5LMxKrc7fZoWTlWqjGvv4sUO06JQ9O
8gwk4zQmH3GTf4skjsDx4Gy0ylfNvvBXUERvHq/WOQve+MgDzJ+4GgjkOs4HZLK2
9oXEbkhNhYuK8VHEzCewa+ed261LD1eZPJxcfIROY1XLhk24Bbqkkgx0ameCnflg
z6iOsJILV1PQolLOq1/MwkXmTdvIG+uw5i7yhKJNg4MlfkvwmGrgpZFwJpVAMip4
l1Y9Q7ARZ8IbIzvnKNKxNkF4Kbrb1Ya85ynfYoqt6dOD1XqOd73BjT+akht6DsUe
IVGPb1MAbIoQYZ/mHAQb+9XcP2CKN6uMzZEhVSuUdsP8k3fbwZ6B8wSQh79dFKxE
AevSuqROmRBTBg2V7zzor4yhDIK158IePFoXY6HmlJGGbm2E7lCPwstDKQa37x5J
IN6Afx2TLOOaN+WjPU6wx+m+5Qmaxt5YGjoTMFJifI09HL6teQlqbPTHpc6OzGZ5
5PyyGab48xtdyKN1sB8GC0hWEeLKBPbTHGMziBAhKhB7LlpKlcaIDE71BPku9J/g
+O6Dr5e7/kPMnPGSTEvGnTv+pVmkd+OrwoZpWq7MyaKj5H5pYvEMUxySJ+F8o6k9
lC2l1eWe9tUlMHktfzgSy+OQhcc/fpsqft/XDPfEpXDP8sg/AngK8Gh5msYDrVay
ARbI3FG/1uTHNFJlb7J9ZKflEhuMp0aH3+sDvCfe8OfprhCFmaGJYktSBXoeZ9gp
5K23IK6z3c6iJDSQ7EpgJxPrrMm1OG0cUvzc1YVAJcf83/gt6JMIFc5tA/YRHpCr
MMFjcsxjxjG6bMcDD7CulOcQFrHwkzjBRrnhey25a67L0nHk3LIK4BTHvGLjLgW4
FsCSCDq7+cr8CviVYFcgVrpDPlrdLtUNch7j4YICw0XTK3/KFYIXVyaqX8BehQvR
iQfqCJBzMxu2LKdYqysoY7/IuYd0YUKT8za040Cx2phSQKhYRpp39xdQ9IyTLHjW
OSr7BD+Wavcz41JFjmpJ0nkQIoDGQhwgT5lpDKhgEbmPsUfy9wNmYAChcMxDnZEQ
9uKehVKfZ8mDTA53wz44Vgu7MrVvnYtdKcku2PRma6B/GNHiBm2z58yQ7gsy6OXe
V8kr1hYiz1f39Usp1noN/G229FxDeCzP9YvmwVHEWbAp4wiZiQ1BCkjlhrgr6aGP
e12G70Q2gcEGZ/JJyVTXzoGejf5L/fBsPM9XIAgPVyo8aKI46DcO+we8hJQ2ixwd
NsuBh9f1iT2tR6A5YSvcmiq+omTfmBGOnclX1x02uWj/R/zb3rkqhaqY7eXS2MxO
85Ms+KqM8EFkaLX8iECJsjVIQmTE4Y8xcY6D6j7NS8QYuq3j0x57JrANUgsNkxWw
lPFMSSPGlhPTBFMDN7S9oyAM5Yh9ag3Xriu8qQCJBX+jyNtysJ6OETHLcKOJUakA
PPA1mU38StGDg9Y/X3ye+SiumGdp8/6mkYR4wbdxheUBqhcxAUVQGFcnT9oFAhvy
lzxzE/ktcQk7w3CGMPsdUHxyZHtAN2Fdj4mDJp0QGDkPuIDJIyI5i0+kVnbZ7z4W
wyOP+8ow2wOdQWw1Oa590DSY3g4TmktjK4lPpMgzrOz/OIvEJHBkWXTtik9rwitn
r3lRrwNOr5hzTdcfut8OJLwOBVTS7EnQwbyXPDw/1MLlWKBsDmOLKfCDn/PdvasX
A4wEAR8a7bJIre9X6vch5IQTGtMHzXkMJCtUMn2Y6nSfJApjbvb0Dp05bvIB6lhp
/WfrS5+DdlIBIm3gT4xP7ngwvlV/uWwbjg3nmHqP+JuUZrdpJ8pNVj9dan+/aX4i
Cy6elDvrqgIHdb2BS8H8oBZU6ipBadTQXozW4sMbmogLT3dDC/s+HWN4pIrsY4QK
rR865oQuOmuLpVDq+MYfLEr2DI/7FFyCF0AmRCTjRJkL2IsJOVuFGp83FrYG21t3
oB9Xv+OWYC5uZLk+P7rlW/Jr/lLIiIKfQbE1OTUhJ7NJKKQT1ASNDDA6iEsRelX7
3syZnDQN5o8OQH18PzUb1KNdg+ALlR7js8EkGQDFrk7X37LcXbRQR4uyNwDOY1Tg
CjKLJ+K8vRjEaeSkpX8TOmDVNRGzSPDst0aC7hbJ6E6m9qKXOhtu0e25EZNgODRC
WqoNlYcr9srDCDFaAtiw1faZP3aAyWd1YwAWG+ITjvisLO7c1N73HMB62FCgtm94
BhtvlR2UepegLF3Ig8eQVuOTDhyeTx+N6MHZV2PzCTsUZHKdtqhgA6JL5L7TTCS8
37cUvfC+C+iMlXio50GNxowNCN4L5Fh0VqFCsAR6GENngobyoWj9urE9FS8PViib
utFHSs5uVn+wXCjTqO4hU3Xn8B05noaLHmzmkriJV782nnKIgpJOzY+0B1JrNXVz
BfH4qgEajZotS2rg8U3BHmXNSkLikh8lKkAio+KwDjf+JSlMn4r2zDaDrLU2U0BH
kXNW8wBnTzztsaNddLAQQZR9Ns6GEplVsbtAxk3eDsbCSlKEZ2zYkRmz+HQHAtZj
WwvCX1QYGkNziys7f5+Rvk2E/dlp1aRHTXrwUDiYnFDR4rlvkQObhGX4qb1NsZ/1
K88viLLz3RNPqKQ/lJw09RhTC+OWgLB6S6kfonkMcVUvpTAxfUgWWGAbhl4/hROB
uUoglcowp1RNbsglU4SwQZhAIqSVHre0TI+fr3SB018I1o82/6Lv5L7atW7D2BoB
EDfJ9mzQUt/Mzxe4VEW31NL+1VqlFVHgv3Pewh4Tm76d0vikRbWjInEhjAXW4HBv
vWEL9aGqFwFwTYW/dNmlIrWJqbr+NMlcDquOfLBuucez/3N5pj9h9AoOHY5785md
jNkCxDgFtXZ1OjvJYci93gt53oReGyIDKfqck2+TPFdQ0i4IDhTNPJ+vU4e4Y4gW
HYoyhzc/Nev17+ywLRDK9p3ZaGFfKrXF1/oLr3ZK/sMIhjhym1lh4jPF7lfdBHNX
8EGLkXOD47jKZH1ej/+/tc9GVz7yIRe47FUD1Qfc6dDxD9aFxlyBTcVuA0Ou+pa4
gN9TrFps4IbCRv78MA5PslTzq9xXXCdoWjm2b1N70eqOhHDg24IvgS/U8O2vjd/0
Pkd38N/o77mUn1MegUnP6/Pzi2k5/fP4l5RIwkYfOfHf2OY0mchcPphknUJ6O/6C
ke0j1A7F/XACzDCRGDDXMVAjUeVgqnDae5bsw+kdeTHg834L9gOX+HE2Fgc1xdLZ
v0L5awTZvMXnQrl5TwpPbKw89CuGRd9Knf8QGIWJu29nFqwhOJt+r6DILmW3CCC0
i08fJCusrMzJVlo3UMtVDtTQZfQ5hIsRrM1CoRTK58J8s434weq67LHinPLowUlF
eedHSVWKFGY0W4HoPqD5UNKWQ2A3IptI4iGYHhQBHHlTR838Q4AppXvvaIkqLJRD
YOXTEccQrwHLHyqZ7MnrqTaWkjGrHmEmiRPvJm403eAUgg4AuUDhFWm4UAldXiq1
Eb52e65rIUjBLeufJS5C/tWpVwIFQvi9rmj/7hskU5HJ9HSFBESgqtWjBmQQRMod
vXhSnCq6UxoNEmkf8+DGgbTWjxWKjE4M/p3tw16KUfcpGH6Jy3xeyakBdxaQ21an
51z1desdOyhbF0UwuY3e1LwT8s5tks5yIjB0yuNCs+oBlsGwLQ9dlknuJpDxjEXc
KFIwd4iUTAssSwiobz8Hwyu459vOmbZQ696FkTqgXY+XS1sfVZM3a6I9T6cP3CQQ
8+dzTepLhRPsPBMqTPsEOW3u+J87RwdtHOb5r0oKJRhco/rTh0leLdyDILIIbhhL
PlHeBeQJMBtO1VaaplpFlqUvPSrqltTHYCT+xplxY/yPc2dE8oLe2SP1M8adCS0S
Iwkv/ve4sQ+tyz6Sn5FW2goj0/zrSyOeFLqwQHV6S8webIqUK/uZsB+/BBGYnEkS
knf5qx7J80Ep+scp0JRMhwhBDNdXkv6TVHMM7nglw1Q0hxaDd91sIoMKLfpEDVBW
DhmMmgaOKWsuS7Y0wUf4PJ/Z/UAhtPJwCErSblygCE1yiKIk1NyEldvGI/UvgPNw
FGo53MKEOc05l0TJFQFTFm9YQE3FWdw15hVWHWCr7N7TgkvUt6Nvfr3MmkKJDPWA
kzl69MAiTxjj+jAhW+kIe/EbfXwxqGv/kqwYgeLpnqJ5KH5oCtrQYDEN5w4C/vO8
tTBUSJhYuDVN11PjjeSsHUcBA5EKcAW1nnRKh/v9+J4CoOstB3mtOzz+/qRdou+B
AZnMeo69aEPyIfP82CfqtorjOfQfJQNjQL1hTo6i8xSHshIl3NcrOyJ4vOcxSAMK
aBB0JHcvKuIQIlaAmtq4SVPKx3L5HpL4PgYJdSjdA5ZH3FO0uL1+NJA7OXDvy9xQ
tce4eVOaQ5I4tKx8Jz2xicK8pqDgYC+gkCKHKJWDcrm9suLgncaOhugqILvN1+bD
ZCWFLgjLw6OL+2uBOgPs7KSOrom5RenHeVnZB2gPMcOaY1ULEp0WfgygojwHCtIu
6hLwcMrsUOEvTpA7uorDraxZ80HPPNDD2b27SUzoL8xn7ZKRbauT3X+scFSmrKUu
6j9a/hyUbm4zE7Gc9d/cPj5Aa3CEaJ44lxKWU/WRMBqYn38rIWm1FA59c2BI6++t
jNM0ooZTqUw16sNyUGgo4wbuq4aDBbUGfpoRHCdPRp0u2dw9mLH9+xz5QEFSXwcU
qfGbTohSxLKtS3dEUMeatEi34ZuWG65zGispYif05yND+883NxnsIZDb3vOesScS
ZYV6J7fWr3RLDX5Td2j8IEkg3RQzDOsuVn1Lj7dIqQ4sn0Lpmf9xyVHpBYVebKJs
1l4yTKviBEKV5Co55y7xSOwuch1BPW+CizS8FHyQbBVKkFvdagCJUQWkqe4TOzio
3wB5XddYA19nWA9xFKRozhe2r0XN37gplUOwKsuE3jjIFk+mTOQ6UJ7mMHB6x90x
DC1y4p0oAOkz5moaNlGu8vpRrWc32P1e+1Etnj0RmLkNCD2jvo/P+MBqRpr+/RxG
bLHD2DfIlMr1TFoOXoh8VAkjOl5H9QP0ZqBQWWCb6Mfbt4y6Y9mitpN/g4xZVfno
juBjkfMFvgUZdvrg4jlMnqyHktR3TL6Fo0RTkcWpsk19dSQcPyn7n6DzeLDNf8cF
vAij5RHq4lH/0PGhYsQjbDyZlLUQSpaAs3K7y5odqw3yev/rPU1UmFDKkrJKfJRK
W8AjaYwsd9gEYjjnAHChQGJCZhBDUOSs/OxmC/OKZBvDH1TJIweQ/bBD94+cWwjO
J+7LO/0GSrQntevn52F41oBM3VpisQbWE/pC+UGLQGpGxINMewLMbhwX5HGQCxiN
AoG68BQp01UoYOz819PCTJsglMo7pj32FXplBBS356w3w0C/cgn0pirdLWfatdl+
buP1AS4dUZ0oqbPEayPkAJKd1xlDawUk0f8j4qBlyp0tXLCmY8dnWBy0nl8luI2B
u/Au/v8W99isP/d26oaCszB0bUPzrjnzjIPc5O7DrtlzcqBWgogsAo9+bAp2b+m8
7FOLMHZFGuP/8Kzoyx4w2nB9rQdvkyGGhkfXvwBMpTCCirgnSSGvYQap6I9XRgoH
ihics73eSyV8rv90O7yFwKHIiKl5sNEJEQvmg7wauK5CSfZ3jo6UcgL99ddlPJtq
hGvQRzktIfqgSfTEZJYSB4GgYEknJnF9lkhfp5RhOKtwyRAIeW4Tnnlmzch5nrRO
KDWoNkr3I9jTVNTzKvTg2zoTu36QYFzv6ZWy6HzcqDp0q0n8WdC0cckm0JEpasmZ
+X3/2nukqzbSd3viqN5ZFEBUE1NlM5MI0V9dDvfRzi8wwTe8zZQ8h7Iylqdt3G+E
STj65B6r1JXG5i3UnRSMWKbPy7/wESnEWKMfL5k71vb4S2C6/HFlNT/ESaVj+L4X
Qz5JPlSntdz7V1HzNcA05s/zxysWyVewLidfEG2jKtXicF8rSZ1T3fidrTpvLs5U
WWoLX5ix6+HrE0vVdKmHehHLYkJ1b3KE88KDRA4u7bC7TQw+z692VWuvkb3wFhUD
jMQjSisZe9KrRhk2DY9RfILk+JUckhg1hpMYtXN8h3j2ecHS1TmKpslpiSZsOd4a
GOXM5F2PzEWGQpYUMEc9TMW+Tci2lf5Y1cYKXUHiuGO/dOQc8qrn02D6yJx8SyT0
bOanR5mY9lho4PHFxCm7thIIJ+h+ctIy5SKnGhjuz9FI5nk5OYRHNhiD2yDLoMNo
wKMmGHN1bMX2bBttDxnx/GGyUDu7hjJrF5Web2Vk9h0C3gcLWghzkfShT9H/ydWV
Yqm8yvdo4YNYD6w0AJ9A94fytZFqhBWXWxtbhoi9X0YukiOxNdJaotpTOdu7OlWx
FfhSEIyAu9h2brrpM1hqRb5hK//5PMPa8rNMS/0SG0IiM+CYHeDQgndi18vDEKwq
edZUB0aIiW7+PpYg6iTMBIPsEqwQY2Lt+62wwXVxh7Xkwx31BaN6B4Z0dPjohASq
em2fJWxB1IPP+JhXnFGLwF4sjj1AVNimrYWOTA+aa39mFq6zuXuTs4wJsB3lttBb
/46P/1dTeLO0HCy6UbHgty+1ZrmM2InCTaJ5fsRAlwReJKRMM9V+9W0bffO4n+Ml
Fd5LqEojzfYViSNkjo2Z+Gl3n5aYlhXcRmNsm3KM+uKDZffyzC1D2fsnYxmcONCW
1uSXkfpN3K3LLSmQNmSmcMNoWoC5MJvSrSSB4nfijyj7OV6z+4zTp62S7GhUkH8i
/uOZ+haSf+qucutmMB03A2ggbNkIvlcTd4nmEYRX/BqyYAFGFFZ/ZonxtxWWRzwJ
QKXk/F99STmymhgOhfg8mgwPUfzPcOORp+0uj81b/c5lh8htfMM7A/8q9ksPvlL8
UfuMU5Cu4j99I13StfgIxRcC5aW+Fr9QrQJLDz/DaH3msS1+j5Gxgl1U1BnWPvEJ
FY6Xxd8M59+Ovv3+JxwtXVfWbkIykgVeU5EfUsuPj+Nw8n3flVA55u8kzumE1Hj5
BTKoD362YDMhRHvMLYyfb2eiNOvxsiiIm8v3/esgGOaLJbDYtd7FZdY2xpRi/ndY
Z0mgmkgqdotQMifhmAFt9GBrDZlPsXXXmzNMnV87W7q7CUgbXQHpVrHgr2W5I3JB
CFd/x82lKbjz3ju9FD+a4xfoYPa7603rggdYDzBpOQgfj6MRXGWti0WYS9QosQBo
GozWHelwg5S8N/WtBSwoxRPu4gV+JHHgMiVNtbUCeNEnyYpGhtKmSPHQf8iIvYF6
v6h7bd/RBRtdBWUCtvUQXcFnN6ddEbEnFUwarNDwyNlyT0v+wMVXftV1qAvXlSOW
wBqqG0FXec9y/BblLMdRJdC8A8PsGwdIwoPPWYj59EO6IEhMuAof8XVW2Cil2Eno
rM/qmdRq0TD9qzOMUxVXTPd4YeCyHrZ7srAJEQnTvv1K8VKMSzjRC9wZ4JP3xaSk
iA7VIjpIxGhi3TQwR/6GQ4eiyLxWeq/fL/6msFYmVQGmIIGslxXMzDL+6fLUIifI
KNbMzJNEXT44VtMiIn5qxSYXyRWFQ6lSAtL+NDsDXEBazmhFNBmhvqPPzCLuYQYb
/1OMoUlxviWuJek0KOEvUqciAJ+pjuUOtFY2i/Vq0nOmCcGX3vDV4BtGvhPtFdDU
wtLA21QneiyLlZkvcc7/kbrc7vRBlXdXcYSSobndGX1yWdqlhx5U4558d114boJ3
uz+KDhzD2UO+JNITl7b2xl6w+ZdAoPCJE/UxK0DKgSTJRik3jeR9108S7nkgSDai
OnHaZgWDhM2r78Jhiw+CYlJiQq8+SDncGOxf7Y7poH94LLpurpAN9Pe5DrTkfODl
E5X9O26EliW3y0bS26/htNkrCHlJl8FK+z8o9ysO9Ba7iPK0JSssJKb73AnfKZCN
T1sm1oGfhx53kkUdJ/+dr35TSyWeRuOgzJwl6VtUIJ9iXpGw4rd7dniNErnANxzk
fGFBV2z1ZtsR/BAJICXSCK0uV2hHj4U5Y8VoZJxV4Y+JqoSLveQCAam3+Tk69k4G
MY+T9gfJk+hFhbDojdSeduszVAa/mhoSmfGChaIQ6J3fXdSVpCuvtCxEe1uOwN7M
7+8D9rjoqOr7Cgcbzja3GxmyYQ2KHswMhPN1sTNlkOLW74CNY5kgTBzWbCHQha1t
us1t7Ex4QJJ7SbDUy4VoyW4hJQ2LEQaVqJB8ckN2iczxldUC5E9CmxbZVkhTvTqp
83mxcH8YQxYBwssyCZ0Ukwx/6Pp+XLcnGDjTfhZHmiej7VG9gWgfe8dhXHDalvHK
O1DOtTOtSVMagSTm+uoGXRvru8dUFl1FlH3rpqLDjoOFUmwXG0duT+bS/M88MjMS
5PXnnT9vHmarVERXypEQCbN5nxl4wm7/g5BfPqL2TbkxqZlXN65wY/jIvhDSjVDJ
NiypT9Ai7l/sw+p7e6MHZXd0QJhT3+cWTZfGpswsLmEjBhVs79HoEc/WSyfzCDia
UNlLLa8tSu2/ZjqAITlLfcD67E5HdfnVQidf0vtucA6FfDIpzvYSQBnmc968TwBY
66kE+AilwmPvjlqQOYYDWZhtq5sQMP5rAj30Z6T80ZDGuoTVJ4Jky+3RfB39EkJs
ujMD6GKB+7MIzH9SLDUEGNcza3N56pwByvJxAtqGYiLyYNRYcWqhWbXRsNmg2LZA
sU1yHqrkBtMOnMTep7oJyguMwJx1uWtsSpmv2FvOL72oaRnNyMtQhcI5sXIBIf3d
Rvdi1YeidbwJcdzAS9MAJFf9+vSlHcJ52FqDG88C5K38WA2a45d6QmonmnrWw38t
kDJx7LDL6s+5XbwiOfkaX1mLfkGyfNZdt/tYSkLK8JoHfieKopaYJD4g4y2l9Zft
9KLY5A5WUjzzMZXLQk/kBtBZpggjF3D8lX3DSDMjFwE+ZF5Yq+ORZQwLmqp9C2QN
mnhVpjRSwijfiG9xYHIh/iwOMk0tX3c+ObqZAnifPlouSBTvMPGm1HgEjoVCPGQn
OYWlj6n6tVy2f1CPur8dH4NVRxhX1BU7eOo5IW8eC0G15mf5BeQ9iT4uMmsoAp0L
ALH8ke3uqfesN88qzJ3FNDnqDhlxfV5BYw4pzdhR+Ky6efwCPIDGKdNiYYZ0Dx/Z
u/uNMgjr5Z9MJuP6vd0ctaGo3ZYA9jVhIdsE09ZMhMbNNnSugmFYNxufivmEOWBx
qn7SVS4Fme/dM25UF/IkAjY2asFaMQLYuFfVtXWGdwe1aMdsgRxlCls+lMW0N/fw
ntuH48Mvntbh26SEsWL3HqO7dgMXztdmC/lbOSSsN4KcC3HGAp1n1SilT3L13ngL
7PV+jnu9RteNkGORWwrr7N79aewvpMnzKR38UDVVfpGdS5xZHN4Fa5cpI+IvmcC0
i3mG1dPwx+Vgl0AAYQQxRFSl55QOUkqTkaCqTrjaSaCV1IhLUf9WFudiW6wu65AO
SSXLe2wapyh6kY7Ku2FR1+lhuokYMw9n3e+Epz2ZsMHvBKU34e7fB+gfhWk3IA15
vPdaKFI1sJjJwm4D1qH0au2I95DI7a+nk+eglPEoU3FlImSrHC1W3ZoJBUt7xDuZ
5CltwfnGb3qvaYk4mnSAYDAlzYTt9XV0yp61EDD+gpVvg+pzyp3Sl3IcIPFsWdVs
keF6h+PNLzqPJ0Vp/MKP3VvAN90Gy6WESFXX5MXg465NDWZbZyD/WdnjsoNRe4sy
50BIT28q+ZBfApex8CowjdOPLRrBLav9EbqiVtxq3uCUVhuxVATnwMvg0cIEVaZP
uz95wUxlmssYoGysZ0tAWXlJKohEWGOIRfAYbBdGbN5Uc2YKClkNA6ApNMJU/Ygk
mcj5FIrxzYuQ0hpl4ThMvh78gbuZdGcD2XmyS7zwr5fOCLwjZ0Kg/V03dfD85pdx
PKjswn9PR+kRyEH7elCQp6DT6l3nji8WBBlB6mqqLtVAoW1A3f1UUqcx54JS7vjs
QYetXKpcYUlgVahiax+sbVeTBCgshcBjOk7Mn7DjF/pFR00wCfFHc4K29PykKYSd
sNXRnoXmaDPF8tU5Jl0BtA1rZv3fVAEZeHXWmrW4iKXUAU4MDJ5zjTQyNvQb3PI/
tXfH8rHyKj5rzyuVf8VB4fNZmLQQqimCwLl+XdYWfKP2oi8Pg44q5TuVYaXR581/
MyQM5gjsf4ugf0coN17EHU2eg5jNWv9XJazOuM2Iiu6fcTmbVh/hZy/PuwUZOd0F
Ui5NLNtwi84WTSY88lSU1u/0Q+vPIon/qCJCCFSZcw15MNaEFS2jHoSmzikaS0vc
6pWf1sn+xVpe29kZdpFBoSBjgP6IrdrJoWxQwDg8PoBDwDGJYD5Q3KP4fTT5v1vU
Wpb2pAAcOEfmYg2EwrQ9Vp0+lfWOIjY80HQZVgViUU0MujYht/vmrULhA44d0CJB
fZ90xc4+hNG37adV6n8rINHZjXZ+9xOz4iqveB8nfTTRst9vBt0FHSheSUBJm5sS
26DoDJwpASEkGIZqgs+ApwqxrZCv8DFz4cju6RUAYgLJ3l5H9SCqeI8Y4oDuHxil
NhwVtnFqOP9Rg2V5aOauQyFkTK+eSyjGh823T9tFf9tosL/HmbZBEToRw2ki80L+
VKBNLVsA2V0JuvDKpha3qGy9zwyJmPtvE8Jk305qRBZVNHs4T/lgjPNzPlsIhkvR
h7g79BcNNx5p89+5pZnkqPUD0gzSmHu4bE5eBeWAOu3KYx6EMZzq5h2BtVqa6yY/
SAtsZVvD6ONK6O+wNshArkqgmOneQa57HWz+ZCcBzGAFvEL1AevkoZPNLRtGlY8f
jU0V9msgKsVDaWnmjzNmxeK7/xV+37KFBfkKcwQ2ao2jPr4lqhaFQVVVnZ81rQSe
d0x0kGcyjfeqc7TJSqCjNyx6n/n6iPy7KycfOIiGFbpwF00VpI5rqk4vfSdB0164
+mg1caC3xtS1uYkDZH42XXCZ9f67q15AiouRJJD+C8gz6z9feHc4tS9RUZFnk1kO
Wy9gipWSSYSMCgoSgzeUfDI+vwmkORVCdb7GZna2usxy8jnv7byNyNvG0ckLg8Gi
pVdEOYBwlPU/fBnhjVJ4LTIti3ab8Qtl7r7k/gh0D/aktKJ15JhQgkjx7GZsnJzD
Z9HDr86ccmkhXE821JICWcRUbRUIcw4wwd9SKM9mzuDdsjNQpY2zOoHuJ5NMrKA0
RGEYL5MPaX5Lkkxt1xYbUYw8+eE237UGgyC5rJ2LOpdbtmljz2yaJPZMYB4dcmIz
SbJXqY1/qx3OeWzUTWxTe5AyLOQGcQq4BTa2FIR0etn0AfGY0Jgve6I35E0baZPI
R0BdFmGW4vM2F4eEyBp4If+GGcEthbXUfOQ2X2r6ktt//jO/X3vyEUSEjKu3Y1dM
Iv66Z14rATn2RUpkz5qJ/f0cRjhmftvgKSaEjKEQAlbPeTIAj8pNRrIr7T1Duehm
u/tFZh03MohGsFlaxNryWkUnwXR0KK3euZw1Jz2QDdJlbnIORprIFQ6XRHuWOkTE
M4e4EYbD7HIu1rUyx+LosmPNEWklbSbQbZT/2ZqIb+aVxzg8zigLVyoKtxDlpNCq
jhuWBo/SYGwSj579pS3qnlnSeAqNFkjxh5sosSCEqhKwMCVsWXpkW82YwT6u+IHJ
FrN0Qv5lDOnj6vG1akzzaBR3TE/dwOHNFo3hZnqV35jCtU5GxTpSIKrnv3pT7YWS
o7QMKDGoHq+gbH3VcEY2AvWZWTObimntz9K5nxae3fQtkQmuEOhxOW6mMsL0lHFs
03DyPTw9RLVPc/HrN5vYvGItnbzWRudmNuglGEkQSdtUdN6CnZQzuI80fhnGNm8k
QFWx3FFejg3BGkU0tNUGZNFk0sW0/i4rte+jeqLwncLfHr/EUubY41H2qFIns84G
nnl/6xXiRc3oAbFtuTI4nFIi/wrnEZ+qffojnX67HX+P5qA+/DHGfx84EEst5oyy
Fe1Uq3ILEpbv+LifO8H65gCRvSA8YXu3lzLrakWSjZFx8ffrQJ/prK1CQkiaw02T
X1mTtw50hWAFx1QMJGgDMu0rEYSkfUU9t/+bxZVcV5egJ9C5B6J5+cMWrjxQJrGJ
oENHhGdQ+aURTqHVQwtgrs5EzBTfQnLdVw6asbe+riDWHtc8TnkK/hh41PPvQH6h
ZpYYtSTQVs9ve5tn3zDgQkxrz/5LprRtIrqkbQn4lRgzC+lGH1IsRY91n8xXxccC
/u9RL4cV4eEwoZ0CpZVYawQLoYmh8gNq8K9AG96oVo29rKHZozCGtXwSb4m02Yxz
29Mv/f0zopLjwwy317/MNMjCEAEeIrIKt3cejAq6EOWqsd6tHRn+IkofOVlCD5EA
1d/TIYgd1h7XO4HKAjaDoElHYcB4QyqihgeKZuTsVF9W0yTlKCAc8+HCdY8iklSw
IURm78T3d2IKpA9cI/0HH5gi9mnJn7ssR4bWilvit5F4X0tAmX9Lq1reVNBovFCM
aPlhJONfIT83nPvbLbzmxNvc+2DU3azp+tMTkBllISwbqpc7VJZL5XpDpxEsuYRm
qrLuz7b+7/EgbfiVotHPRqjAd3rJ9sPlquFCG6Y0fcDCPuPO/LnOmHji7i/lq/AQ
Pw62jG+EVAkhgyhWfBHg6rJ4IR/UwqwjI1g3rmoouRbrmTzREknXcBPkpSmZL2Cu
PBfmXvA61MpyJPVh8ftrfMVHFYVekBL3kEDHTuvpztdG77Z4Fi4+CzEWm5YmS1eC
OmUwBzf2xdK3lEZAZWh8b+1xyo5Su6bp0x9Bo93aE5CUMzLpKOfW5pzdM4YmOumH
cUxxRSVywqUnPkVlNlv3pc5fMKVxkUGRTqU89VarZrpZ93y+dZR5suP77+gN11XZ
55ECyiM5bw1P0jEFEc8ILEjt1XNxCXJKJJFwdo5eZi3yBfI3xEaF6IwqiUFEhhx/
/2+OuUTCh7KKMqJUgTmWDRQja40k9ANmLg3+eJeGIZ7LahF15E1iZEJFA3mdWFk/
HAATYDs9B2j66YW1h1RgM8MNRSQQ5oUHFlMKCHXWUwrtmIgLLzP0Y6xv7bsHqGRt
Lt40zdxsUaDRM1cdzQu2JPCpniK7gveJhX0aTRCsigpbRUJUN15TMFTCl5Hx55ol
Ir3cSMawDGB6eQi77OFMxQSubSifBt2UXZvV2Rh4SpfbxZgu4VloO5z81qdbDvfo
MOzuukyA9PVVvqUMASpbeaFixnMNEWuRCzEjjHMRqzOu7crJ9+7XEoTupEVPvt9R
wR4e6XMjvNCbDSNL5bXE9ATya99zCMMA+ntLCzcaQtMreUNTQMh5J9VnhU4btc7Y
eU1M2PujJRH2mzIaoR8GhIf72kn0loAOA74w8b9Tk8BrpdRpY5wx5Kcv+J3F3L50
RK7Q4bX2cNQsXTgbn/U8+cQ99+cUj78qcoawPC4edMOJWoZ/Ezb6sz6prUj2zzwz
Y7J7EkUZ+NfQuG4RU9OtzInam0jfJOJwQNg2sWA2BmPT454keE02ykZBbwsxtedd
2I8UrLIf0s4BcieC62ZMBz0LmUObev7z062VfvPPaPqrC0NHEA3RbZp+uOXJs7kA
9PQRsSD68EwbusTb++zUT2V0+8H7KwKUl2VzerxWTmZOW18vn/WNBYSzw7Lwg8OF
DV81b9wlkbBueqts+pEk+cBsiQeGmWYaA7BBjRSRxfvaMnm0sBg+I8ffpKFFi8M0
EujRyM2zKMuBi+GsefTfD1BQYiMNlhiISm4wDtP3gdHG3g5J3XpWp4kbLlQsd6LQ
ZOnjv8Q9z0ZLZNDQ1mCNKM55ea3tLc3YMHvUHmToevQJWU5KCDvYzYFyueSmix/Y
zWESn2pXkL8HGvs13rxRt2lNS1El5PDEutv8iyHMj3jm/QddNmaenxL6P+QFcszS
oan4Px1YSWdnudeYRFsH4K6bx0ioPFC/eQMbdx6LjDKOgPWfzlaWD2wl5hLmYOlo
Z93RvXPGYPEz0EnaGqJFCQ0cCe78i85R5IVpA/TFUjnzzhPinFtgzd0btmK5QGlA
xbcLL+CEBzk6r9mrAyCXeMrAEqEtWKq0FI6lJsHURv26TnHabHiZxPTVh/o62sLq
23H5ttHR1836qOaENhXOQfS0RlEJO2KGzXZbXV7kM/d1YQ+ZKH8v+cO7rSKi55/r
2xfuid5QkkpBjAQt9CmDo6F+BGJa11jvAAAuFBpTKtvMCix4LnwM+BAS+GvklDQY
klLuS+z0uqxwphs9Iqpv05npABuuUo2QLn9zKPbg9uM2UZqNpbqaIyOScmHTO3yy
fcoX99LNpeFIf4G9idiwCx40G9ANnlUlSyVivA9OKwAIOcgKoZPfhfA1ne0woGHy
EVpeZkG01cXg9oX+nOiGAG3dAvYKMm1vCpEDldGQehRIXwsy3VPVM0j2sWZkonpJ
dgnDWTrcvPgmhg2FJmY2RzUu/tsxeYioISZmGslHGfxQWJ1YhQbKwzoNdm7ugNVn
a9d6sdE3XK8pKYnTvQIqcjypoiZuLVBHqv+8oF+qkAUshTDZTvIe5s2b4n5ug+jq
y7AMxYA4Sb2sH6jy4juUp7mG0yfzjepDWH4fokrkaTn0SgmeXecJoxO+e5NM6E26
EcK6lEZdnBed3tRAOMzpj+d6dSg8YVoI5ASpQfOPh++X69pl+c3xulCsuRz4tPni
3w4jGopMnOhbTAJgNmak+rm6HnLjsCF7JQO7XwFz+Ety4HGu5HPTjFFoWopvJcMA
gLbwbgZ1craXjERoMJNXUMfdXFiVTxsPVw83fwnItPRX+z5bx85QGXoMOYUEF4cD
Xf1mpoVQATi3vlB1N4XYgzYnm/XKuhRWjRYW0PzI/8vEvsM0xXzqym9atNXw+0Io
TOTWy6QX0bfXAr9WpxQKEKgTeWmyP7KHkru9I66NWkzkR5l6xUxxg6p5yy+52TVQ
G3Pt3weEr3BaJImw1aFUxD6tF00FdktHwDUaGlLJr+mEVlUpxPvml1nGsiISnV1a
qR6QLbMiOOnWPYH1KrjtlmPKFUTy6+qjzjxg5++ZLcE3qyuWdSBadNvrMvGXHOE8
4USEtlj524y5LF8fXYXrKHRWRJBYFBMkIV3iQUNKHXgOu31hsbuWduwr3BsNMw9H
IipRcb5VsjGwHt1kQIgZ+k2lcjAyuZNjukSGeS9g3JtpZgtU2WwvF5ib9BdW/kKV
GtOQi/3Oh9nE7CwVRUL9qgtX57kfQWd85s+SvSfdbBPnkkzLldxqWeyHM+yeEV+t
7aL1bgCWFe1J12nszh+6mogbb1O0fRYZ7xPSFFpJlFo4PBhmXs3PodnPGcWe15kS
j/xrC2rnkWchJMYb5g663TUHwaAiMNCiJHFi0/M/7Lc7sprkRZFB7aNaJ0ewIIUF
NdNzm+Oz1Nllnews71Lu5C4LDZkMXWwJl5ZpATm1Z3sm8mE5Jhr1+ESc1dEjI39U
8WKB5yIYLYzLtMWHw/DrHQc8fYxe74Dy8dcWBmDhmTFNX8NGy1W+qjexWd8MNZbz
IoOiOL2i+Bb8jM4Dhf2JyNA5MzCm7Et/lrpUZCWVTAciNfBSX0oRsKDZNpbiBPic
TpVaukdaIlzkLjvtfJwPeMD/t53zmFtJDHxVd+GdnLjz9tMLuU1fc8211oVH2qNo
26AgqzKkt4VSQxso/rgm594/Utmrz211a0I9efhCD/QNy4zXb8/kLJBUszhHvOem
8PQkaZ5C6kfKoCIasFk68L4QgyJ+/64QfTRcLJE1IL9LGQAaLfxDVwmDW5kzySl5
USSWAj2KxIVaakak8kBp1ffDv1/cGM7pjGMPRiNyvL8CgBfL5jlRbecnoxaSCQ5d
M640GUM44MWZ2OHfffMPmoudNXtmRGb85JUDczwT3/t1iVoYtBrLVkeScjRlCn/3
DwSMEZFXR1tKKqiABJQwU9fdaIRnJDM+Bb9nuBpTGsjqeRKzTwc3qkDXKMP9o6US
UYCXNvQ/MRGuJIvUVjzSDaUNGsA4btwja9zouRE8B6JPYyA2F5VAq/PUzsQ0xEuu
fyCy/ebRkJjKuZlIK/TFeeYio0otMF5kjWv2uy2BIEB6P624a5x92C6OpBYLDacP
rZBN1PGKBHwueMX6WWJ8UCCkBw32DSr2jHk5mtDiZ/qm5Ibi27JGOj2OSAJlRqWX
eRJLLSvJog8lZPKvVL1UI4jhQDxekw66gRpgy4STm8mRv5CdEclvonEd3E8uCZ4H
8s0XUp8crdrQGC+3il3BqGGpR9iRQnQ464Q62uY/ntir3SJUP6oaWTTTYi+/Cm1s
nJqmkGYjjLdkSFc+e4sI7lSKdkEy7hgiSKLkNrmpqF7wapmAgCLXx2+Vuatgpqn7
tBoF1aJcIowNfn3N6Apf/QwnKSpmvaqw4fqNhfu7y1zVHyqKB4DIyYi4IpodkSPD
Hkt8/+jr7bwe18GOYPkKFHBINq89bS1WvrH81QkeU+5cKPF7lrrnCw7e2BIUzXDw
2Z/uUCaWS4V6bl5uhsmDQtkPeYB1OF2F86j99hrg1/NiwVCrc+PEsSnOV2IgvqCn
cAwKRBhJfkkvDKK1+jrDWcf5Y3MTflANtZmT/xjpMnJbgKQmIMUlS4vKXy7QforC
7V0Xkufk94Y447z9gP/MWulxF2VI9GIiTaSgzbX5WvOr9Lc1g+oraXHdYUjfM8vs
HtkMbXCrWowZ0kqKdxZeZhvGUlRsnZKtutCROmWHeKeIrYALz3SE3l/PRSVPrK1Z
XKSz3UzgFnN8WWKTpNtCDcV7nhSmrPRaBFSDdmmKcEA9wW6x0pdpt9rJvFRObz9H
tpL0QYh1lYb6b70UIshOv137Wd0aQw+IV4VTrYRlr3JO3lTFZ4T1YMQYgZbLk700
qkgBPndGWuHZaWJo249zED+fpSxp6wIL6+geW3yN1JoQo2IZJQJ0LoSCgb970YHS
Mu35WvziI6qMKEnKeSw5FX2IOA33Mb2Y0A64FsrSDojD7vh6MI3XJSdyFTaj5ixN
v0Dv471YfV2adss10HO7T3pbnGHnrF0EdPJ9FfjOPmS7RvirNPMerMKlRcjvG1j7
QC6BskfUTm4jPMoRqHRxQlNz3dPNk+iDpeP8lXOkZcWdb/cVeJvjr1b9pHucTqe8
kPm3tho7MHYoowaRSpgBic+7i8JV58iuFG0LD9lQp8fRTKP9sMNaXbjlHOh7wyqD
LuUR8WcMjbzUS1gE1LId3Ccrwg+udhMRTjITc43ngcErWjiV9EqUNqDxX06zy3jf
2MbpxXh5reEsIhaQGUPLWJd+NAf9mo0vsiCf0UnEfat0o0K8B3tGpRVwR46GvV1z
W8kvKKFSD8+lAIyRnrFmqFjdVgM3E3nT3VoyLTlsYjK5lXoNvTCVIOdzzdxtZ5Ov
K+0Lud0DYucNeQs1whuoQdI4wcbMG5+rdpqBjwoINgSi3Rmu5OC+I6OttBwkh3gr
TqesAkT+IHPYTJou0cRTP27fUHa5IsHOMRjTgcC4ch5tsM1xNqpQtIW0mQ/NcBkS
QN5YQs9vr2V+TW4PryNsz9lRNqCtI+3gQEOWmRkiFjw0uul0X5IijkyoFrsNjxbD
P80gSeiuzI0WAcW5MY7qc883Fc+wwfFVc07VP5SQJhucmCOO0ezND7lbbtrg39/K
o2nai68cIG3eolFTpTm/yqvDphMrTIua7YB9TlDj+a9NNYSv5aibwHUnK8bLn7Zp
SLsBbzW+HBjWMJDKfR19GuzS7lbmwtCmZYxbP9aSYnhVwI5x4LMwoUYLAgrya96w
7qbj4k0jq83dve9bAY2TkfJi5DQIkE102QePuzew7apnjpiKCbCvV7EADRf8YNUo
lb8Kb/f1wX4+wDAivoqlqY5xdXfqoVWVV2wkH51il+dPwgW3RaboqAm18uktoO8e
WPrcmgKGIEH2wPb5NjyJHCa5ewFbmmXb+0zDwChQ5nQ4sQw16TWUifMzvMNugfRT
aP3iM2P/yMAEaDrzJ44sggRhXtj137HNXZK8xVO/tcnOZbT2zwejy1HFprlsQE6a
WV5scU0I/Ed8sFMFSbOK/QBRLGYYSoLOSyVhdWMBWTDmhp/JittPmD1f+SI9Iv0s
CP/1AcZug02VHdL8+AdkjuCXHaUm2pVsfLkJzxLGZ2dUdIXrYRRADoQqpb9Wfgax
cH8tbgd6iTCZjqW88kKc5kwm8S7hnHl+gIf3itaKvc4MwE+bpbzUSJPc2lAsQApi
CmhwqbrEhoNJk/7fb4yYoF9pCue+Tc7RV8I3JVUTk8pG3l7BEW3UBG/pCVtghIui
srzp3qFUo1Ja7Mp7w7DlwewfwDHztzHVUESeSQsXzg12O2RH+0ZGOnNCPlz/amtr
39MdFXEvicFlpbkG0GZZhQVUKKSkq+D8kGDiZIbxLWcAXQyFTQK0dttwKmXS9Kke
KXcNK/PfQlI1OXxqhx8vF1XAe8mWcywn3+YIFU/zN3rBNtnJt2ylP6WHd2b43ld5
Q75hcbOvxN/NC7h7wggO2Q/9vjxNKImN8AgKF3m4F2FqVDCvK7Hp3drLS9mhdzmv
O5gKa0gYr+XJTnpB1MLviD71NosPddkkQN37Yj/V7iGkGo4FHfof4/Y7PTEZF7yy
Q1iZ0MbCxJVA79IpGTENf5VZAUuE/fRFoGKV78B1ZX6qYIVtWYAeZmcutjsix7Ui
RV10Tu1tG0yPU7LPXbcmvuSzdl7dd1e0CdQ4JM5dBfuIsXwYmMC55S3+r0MoFlqx
KbKlaQaG+eHgd/AU4UX/FiTHk/2pkyszayTmgdzr/uD1YeVcNTRh7aO6oF0y//XL
OugIE7YAo/cB40Lf8Hs2ejIBIEImZPBDeBorcrGFmc1VP8wxRoqJf9OFfBVu9C3k
3OCBy+HUyW0BYrJeL9y9LUpDRmHuTDBSxZ87umZ1VRuG95eDKj42Yjp/WqZMQVMo
/bRs+DysNS2A2/e1WXeo2cDUUYIpsCqxPubci7HstJu+Vt45GlXu4Ir3vTQzawgl
rOE1k1icanlQTqRHun1HBgKRC3cDj+n4SyUudFsLgMhcTbEwYy1b9JO4CWnLtVFt
WxVMkoj+ECNQr+FCnF/UFeQ9gQw3sdFM1QnGEMGWc2f+X8Be8yK0zT/iDbs/bKMD
aFXV5CgJM6yBEDPeMjrocI2cMnmDu1TQMk+oZJGsxxj+w4+iGDLao+OzxuqX16EV
2ZqSA3WfZSe4RnprUtw83WKLlPN82tX+cAcozMSYv7Fgbp707hV2fAfq82IKrU/N
aG8pUzzKb7LrzDN/Aq1tnhee9zja8rZjtG6qsXf/I5oEnRWdmHsacgpY07CD4Lt6
ZAaL8nQttdzGWmWsXAAQwkcULkjI7Vv7r2v1HSvsh6O+Fcf26JyjGSIDcOMN701f
2ff26binwzM9RRsSdVC6gwEgMF4YOnu+V/hGIzosxtvwkkVOavYkgImz4RUSOsmz
OmGZCBwFiaS5Qp8fzf1miX3JlDF+DsyIXJmzLWxeyJ0z6NKEnkA4LY4s5q34dSQD
oogPpHeFTP7TYbQnStdoEA2PDP9yGSynL4ve7cy3n7s/ALdOD4CRDRDM6PZIF2z4
tfXfFd60IeTMd1T/+7u+0IygWOEOz3Qg5sb2FZ/PR0Wh6TiWzH4gCSJwQ+4iJ7yc
LMmE99g1RIVOM5nrdEXdsaPmCW5dzultUA3gB6nc95fHrSYNyEimoydiEIMY8kiQ
JoNG3u+al5cxI7OHmOfFX2wEaiL9SzMcZu26kCic27Lc3xGgxXnydOBCOFn+Q/q/
c4ilsjhzi052ya28FzQfRkHbFpPobPIOjHVurZ+sHaa19xc1xOZWSvxDgiljj3H5
GDtxDk+mFxC1n+LToyeV8tcedaf1VZXB6Bu35P6Wr0Pi5P0s31e0PhtlFQhT1aXa
vRrOwXFkeUEyN2lK2KBHIhNRZUqSAmySy+NdPBm7+7Q06Qy9xV+R+XmYXTobnWG7
lTN35GgJS3/LEviEXUpEI8+pWASx2L0H/NLalc+on/zrPgr6e30pzSBGnko22oUy
9CT67D15Ey2Em/mBFvOttGisJ8IsGKChvBJBj8If7VJ+B20LOUugvhJC0GcvkcbG
mBbophBx25wfc7uOQQiIuNFCArPXWycd+9403O3gbhZEampFqBxHe1iU13/Dd+Wf
Lj6TizClfQEq0uNF2rFVAWW4gLOOJnlydLdl8Mz8p7MBbgpYZp8gK0xpSjUnkDY6
7aCUo4A0TSA/VE/pGUYaaO7XGHnqNd03P0+CsxPlr0iDFZji/0DHs+3cnfvQTC2x
3ynyutOilwbkBKWJo4DWtuTiW1uo+3Q1T++2El9I1n+OH/LfnHsC7kNGCXtHS05O
+/C4I3jHHQqqO+f0vjwYONOXoOk/4t+Fh5PY6oKVe6pILib1AcdbSN9z23iom8vf
j8xxp1m6a2wMCwxGerXqt39B+BxSdCEN7D6aL6y40D6AAKc5k7352F6sGGjDkyof
bbLAcqdkzhzfXJ2if1F8WV4n5qQLI0OuS+YJM/37YVla8DxeleHsIGZYxWM1XmjZ
ThkMfbquXtWKzL1zIJnrASQoliCQoJ9hrdiud5mTjc29ERd+CfvoLaXAkuI2C0T+
/xD0SIA/t52O5jcsDi2qaKVxeKpeaZO3dEXBbF8Vil1aYQgdeN6pFGykbvavJ7Ag
NEzpNone7SHDyssZcRxG0+LSyRia2VdOcH0+kMVBNfLVCgHPCAzCF9ZEafo62e0C
bPgfkNyEg6FJ6AJ70/LEg48VW0A117teMfUJLsXitzX7zU59li/rupimpl8lyzvQ
Zt7/rRYNRed4wzSYl/F77K2tRft/kypirXN5CBhk4mblJkIrsO1MUvaWVjd8sTsv
87hPNH1a0osSDs+O9s3x7Q/5hT6wXZcDLjyarKG+5utaagNuEX42/Nhcu6LhKqH5
E/DUbQRCbqEVHoociKM5fTKrE79EUsb6SRUvA1QtD4E8EWJUfs1cLtWREy5Qpx22
l9mkCkOZ7k5eVCYHmcOPdIvbYzA0J5iXX/p1/NsS6ElfoopvgHVh3Le9sh86WjD8
2HNx36lZrkHid+nXOojTQhtKGGr3RStm3dDFt/WeqZnou/rBCHgX73B/5qyLPLkp
Ludxtu+XOh4ZPSpnHCilldaM0DmTsPtfb874Yc5ZcddEsk5FKYEYEpWsgcp9H2Vi
/s2mvYg1hLZ0zAzmEMYEWh3x2asF4pzZ8LNgdJE2M52lvFl/BIn4Xm+1nw7YbqND
pwnW80iQQHhSDz6LEYQrMj3EzQJijsV9E9hjaC78bKp8cs4c8UQHIAOSCZZaIEc5
+y9J8KhjEugS9f8gP4vccnQ9/XWui6KCdpiLzwdGmzxKO9220T3pkbn+dUsgDQqO
vodLl9+V6UNVJnkXOXP75xot2x+ta/6BqhFhkvXzrEBakJoy5tdXNTjoNELqfKOU
1Qq5fRbhinym4DzBL0kz6wW8IxJO1h0ntQFfKs4TNAMvMvoooOs7KG2sHj5yK09K
vgpLX89CluQ4E8paRLcz/tUxeLPsp/wMbz1vvmUEYY4I/SlKwgXTVn8eY4eAGRlS
8tj4QczpMIApUy/68/NzmEydRgYUjWrIJc8W/ubcCcbTPUXf1JmNckzYDk8i4fAa
hhGaC0iaFj7/VOcuemPFXxs4aT14hGT4C1n6YBS6ccIxuV2FFQia82XGvOAryNDa
yi4wJp4F/mW+m/cgu6jPLwDUN1YY6gDBuPjGqqMCsh+Fl5zgCPADlYz+plEvz4Ll
v9fefPc/pd/RgRB5s5NGZkj7Yz1ExZsEDA8mbFIrxzyqTbABko50pjeop7JbeOpe
3XenTUxbKzNMEwQZ0hfWnYXC1TMQK9XqlS5UtGtL1UQPo+RmypggeR2ckKlXmmSR
2pb1y9Hs9fUeZLwHn/78F3BKZdDe9ByTDj43qKBVrflNcOkVG58LmYK4jSldz/NW
JbrnNRYlACrUA4TWkZTBdQkrPMZcvxl7nn+325t7hMGZ5B1RqyTeqafpo0HWsIvZ
mhb9S0LcXWcNmwj4RuQtHxTwHWKXAdpvp+lLuJekf9fW8uHsRf8ZLXTkVebm7tTA
B4/Jy5QoB2/k3e/djmX22nqzff1FWD7q8g7zrCPo8h72vT6oWF9XRReBIpu4DXVC
wv7PYvsdn7RRj9T0Yb8mGbJ35MUJUsgSTRvUIDg9iTTmbqA2xVak4E4mlhdPxCVz
JvEkcvXB2A00ChxdWm5CJQAvfuq9PylrikGaBQOe1KEICndmr9upQpg23NsHv6vd
1ashlfl2D/+G1xbwvA+0G+aPiaL0Lz78228/PXe8AOcF0o+qZ7G9zuIZRPWZq8aj
Q3ir2NyFLhUKeytcYUNzEelbgBMuzrkIHmnGslZipfaQUsUVSMTzEW0uT3I/7DL0
jcVTuYUDWsSzMmQ55EF9FGfZEvh2LIcieC9dcn8xxu83LXdVGdljj3xhDQXJDO5p
bWOWRGFnk3XMqFjTFg5MeQs0kJp//v2UKQAm7RfxS8xqwIzrfGV/qopCHiCKsTIN
U/HSC+QSu6cUuVI3AIbWQbqAbUKK349Y1eC1blb9sNw9Vu0I4anmuJEErBXPS/kl
Sa4MaI8yljTY2pAdfBvUYA5mUB7tc/sBj8fk0E8t9xeZSzxVO8QudwJ79//dFD/b
M+DFhn6ypBRNsDmG/Su9cTGvH70omewWaqIyard3ccq1wInjGWUioY/oUU6GFSJE
60tan+p1Rg4Ma7/H0zQpqByXQBoMBDncypdVT+BIDRh7f4JWpcVQPZTzf2VM5XDl
/dStF4VeDsvlQW0Y5d8MMt9/vn6PYMTGsBkFohmW2wqs49dRDE7zV6fEsXhes0g+
AaOs1DLH6r83lW72CVPQNmjEYNJJgNXoPnV3BWyXpDIDhvc0v7d0IwJviXhG3N7P
X5aLz1b6VYNNg6kLFP3yTbW8B41+qPL+O4tm6L1KypXZNgwJnPY1N9E5TBzUeRMg
OnaMzuvQOC09x7iW6j3fAT657LisuFkcpA0j15nuPPNlhPAxqwp+kK2Nf1PQj4P+
VjAwPXBgRN39hglrFGnDP9J9WlTn4q1GRRBinrpJzjb6Q6VGX16Sy+vixldRnxb6
iwrhONK+Oar+xGofBwLBYEntGA2tKQA1J29nfW7dt5pp8o4GMrxXtf/3da6asKn9
LQcyQoiDgpzd3cHxQkbkl+oDK46kvSjcnDfHWH7e3ba858+A2+qDjD7UizsEyXT1
Fi11STmVRaljZSLfInAoCHpH8C8FsShylRFrmjCUNLl76ebASbPM5mT4ZHLX8azy
TihhWwrf6qaNuaVJ6LBMdX2cu1ASo48PxUmKyjMOldiXL8y0XPzQYSL1AjPqadsl
dsm+bKp0axXbazmZojzentjxby80P3txc9kN7CBp9rIfUU2wQs4T1cY/aAb90RPp
fN/BWMDGBlBng50dzMmacmfmBlBBCwFYd5P3tk728dxjpJBUFri/b2zXvemU0JtS
/J95kGqpiF7KJiLM+NxSPK3tLo9jGq9CzhlGM7x+a7bO6tcwaSvekNh7Bd+X8fie
q9Iw6PkRB81pEZMOFdg2rCizxF9v1EyDHtexBOW/4CV9pmFoLoK3SCeJJgxLEl0g
32gNb3Cc8OMjt+Znzpp2aD6mnd/bu+tEwg/hsoRBo48deF/7hZmVaChY4JjibpM7
U9sKC0u+4miI4noQEVws+aHrr+Y/DGZ+GbHKyEwae5iKx/enWqg3va+PoIfHGU0k
uFTYydainN7OPXlOWZoX37s4QDy19CbL/7oJ45gtsObmEjo7BIT2/dHIjViz+5RN
2GsEzrlIVbReTKg04iWZwEO7S1Nuv4/3dW23jsp55KLosZymaZXKHAZDPbKqL6fz
Z18z8C8eRoFgOtlfQbeAvmlRsAaVJYCBXhlf2XLL5Doz503YzImwdnIUZKkK4k2u
n6TWwbK8PfEnBdLTC7fP1Z5VZa4Heq170z8iSBxmBZgvl7hTG4f8D6DgCaV+YewI
4AFvCd86n6H74eRS0bOonZpjjNAcUwuvqEejMosnDMUwVUxnxTvYvrrUhHT4xTNm
rgsrlybUvTBEz0uXYF8yMmBwEF4cBVHudbjAp/FYRQChEeQpHMO0labDM4UuN7/m
4RBv+47yjG+f6Gn5R1uOTlUKjBc4NcebW8hhfnZRkb+IJvBoAE4O8nJrU59270+l
aw29luOZH2AUvSbJiwFoQ9bry2BIjyKufVG8Grbgr1Rn2cEVtdLjvFj1J+gQgEtO
dOlnaVN3xrfLQAJp/b4Doe3sStbxthxRenoTjA8s/KF3A6zexGAbOgCvuD42pkav
TgFOg73MhHNHfQ2HE9eiuu1yBxKiDnOMohf/qcm+WUK2RIyMzxwWpLZJeUluCkfU
gMfylu/r7tjb4YJEgCqhprB+/lpeuzuhsuKQUYgkchHnkFqf3d5yuGfrS4v3BeXv
xsazjOsL7+/yc44OzeRG3CPVQgFQPj1TtzKyBBXIlT7CrtTKZ5H+LAeYxiY2xdX2
kqKpX9mjY9y0w4fIzwyw8SQYOVAwqqwfiD0y+jv2ASlNuCSdUtXuMxuTg0zHAQ/A
glIVeiSkmXOI0w0EwBv7G5IWXLbtvMoEXY42fw1maZcMFsnCtnnF0XOLCLr9TzPo
X02/2Sv9QO9vr0didrp5Xana8LtaKmYP8KWtk+eoyYCIRO6YXgTiQHnnn4HsL245
aYrsTX9g7nix8EP63ebKXAFikaZntctjwJimAeuO8vJTxvxJlEsHDXud5uH0BdBl
PVm15gciFZtoYvry7tNqjJo27URAMMnrHcNWuPLpnUr34El4OLL8LKo8XZMs0miY
QJaDh2vLEfCzicdEtvzI0gVmg8o/ii3LrluNQN5OjRsz/UG94yY/VE7aSZP/Xgwf
vABw08yxMovxAW0ef/vEN6hwpyOvnnW3047D6CxrhJhz78r7IAeNptfPgH733GmW
iXGfcX7FcaqEczXD9YZKygnT0Kc/BZ5WAEklfweLQHX2ug34kAfQqh6TEEskZcEK
RlzExpPjwURZ+JrvIYQHTLKSIKxJU8/fGfgcX3tc7X+89gtqVXsOsg974dZomjG7
SAe8d4BgXWrs7xhR+LSOjeZWz2+NZmahdNwSAxFaChCkKSwbUlmoYGrFOfMBRk3c
EvupaDjKf4PGwJ7zabbD42j20d6zzL9PLOdTip2++oUzx2nuGhXVp8/TXja8fcGr
lp5pDWwR4mu9wYSaqN9LUhagFDAf141ZWqAIKFAIZWYCk9bwt+1QjEN68N+339Re
XMj8BhT/ZcuE9QGt8UsckBTKq7VoVfUFkgUlGYGr2LpHN/TWynESms2Tkh93pAGr
9cmnZiTHcTCm+bgh16Lo27XRqs4KOM1cq4Y0h5Bq54mw2JrbkhTAMdvY2Gw+u7L3
miPLDKHlwD/URKq52DLgCj4VGxEjogYur/q4oSMuosh0eSwdWVVNOeitUbzYZegX
tuV+N6/yPhwhdJlOtwJeDyVAXCHTSL0itwKBXKpO5FNby5a86AVDYsho18r3PObX
KcwEcCmwsCMhwUkkFwqFEYOXzg3joCmhhijIx01XSuKzRKAjaT3pz+DRn2rtLDJH
YikfPWNp1vBDfwJsuwOw60uc95zljGkr3TNBz9VQ2BAgyFIMdN4AKaEX+UuQ0tpO
pJc83WlV3MffkHRyVH8dym6CCm6nVFjhGNMps95JKvf2fgeRqMc1bKnXGvsgefYx
DHfeE0LSRXY4N6EhqrEd+2m2PIvFzLJA1yXc4VbBSaaxx6Jaj+zFTjMTUGMARlUm
zn52zVM3O7XI+HGLU23gZstYL3QmwbfIhQ8dKchhiTj6PhgF9OG69xVlVL1xU62V
QjLK5jQ72S/YQuhCElLu7FGJqCh4rRC68s8eaVy/87t5gCLUrjtKjcvEm3pHG9YG
MJRhkcYU4os4WYhAsCcI/yh04kNV74hXhmPnZhDb+sEujSKOhfy4Z6YvyTnngILX
dxIwIM9mrvyieBXStDTonEtqa5y1A/DoXMc7XaljzJcTNT+oIz4QJgs4I2jFlK2R
623I+Afp1j1YHLhbVoUCb14T6CdH1t9nKtwzhHGkL6x+apLQS0d5DnpuGgoYKJd6
0HYsRPJmUCcnHQaOqgKpMIfwRxym22fXgLFRVY3F7QQ+cPARjsGoUBAv2eklLdQd
XrxTvLpQSm/VZ7SRUGl+4YYQ4ZgxUAUOeH+7+AHevOZRtjd91wQ7pGznvChF/Q8f
cQyHVy+o1e4KMtdrzz9Bz3dYOKJ+Ov6jkqqtJ8SnUqe4zZ4cR6dcDdnUF0g4DHKz
GqXmQ1C55iB0IWwCP9RWK2XvYtdT9oI34ntXtIal/O8j8ITgOGjr6QOOMU/xhE/B
sz/1EPRzQm5Y8KeRTgeRmtDIQDpvx6VqWFBMjnWmsFh8Nji43luInFx2TvCpiqg/
PWQZomW4HkjWfdvaLp4sxgWFMTZErb/GBqJK7RWjGZBxkLdeJgk0aIeZyOmfHm2t
i1c7hMLE4KtO25KFlHZJr6vyXFjQgHinP8vOCk2qeY/H/yrxFRffhgHPOyE0LtO7
cFRf9bWhXc17BDzOw+GPL/MnEcIs2VDnySzCNVKvo+idTuNlSMgeDWUGONvpbAdE
mUzjUv5YzN9JXmkw7/QkDK9M46h+IForDFbJ20GqEbkTgw/+n4O012Ct8SbrTw2Z
PI3Na6pSThnA3YG47TRDvR4zzQHdiQ6buZ7b/njNBWZLRqY32eib2APjvr69LO+Z
6Xu69MfXdAN3OE84CMlyRDA9tiQjL3b9m8ygK51ffCkBuAdkAfc14o3oYXoXBdYk
DPtIhAVl9MHogZTJN+qxcPDB8Vq/AjRjlRH5yrmzIyAp8ldcuTc9PZkkvLWwI90H
TJ/xvGUYYUOpqDXOnUXAdvNnsRSrkye170SB/45CdMHgTcwntuDW7Q6+8Busx+UO
GogyhvTuR2eD8G9/IlUfcx6tKQEwV+Qr/6sBLoojstZEQd2/ELfV354xMiyIjm6V
WoLDPUJA+qfp/NYb5mhOWnx+ea/hurVaC/U0ViGqiLOLXzEuwo2FD4abyAEM1hnJ
f23ip1p4eW9Ru0jNi++4zg7BPA5+b0JRyJTV+s934m65l8cKq9cdFUTeDd6LSuWK
4gA/W/sNnx6kTaV/cfdVuNbQ+yShUb1baX85MbkiUZXv14x5bi5BUQfp3v5nOozo
vpCp9rEZ6zQ8MkvfBeVyDnmA+wBDheDHDQ3ZhlwornzkkHRcoJ8L0nb20uwwuSxJ
L8eSMIJJBcY7ZAU9TbaRO0hyWU/FvTI2IVb7pQ/2HS5lhwBSXbCir/UHAVqf6zgm
llgRDkG8vKmOXgTQ/P5iJn7aFl9SaujA7iXX3sYcEPxCmUmdXWGoBQwEv2qCeyrv
gDJosYB9PArg7/aAaqXjo3LiG1NGRIvouu27E3Bs46lkiIUQkoXY2+dWZZFSDAT8
bQfq/GoetJZAOUbCNkJosDm9Yar25MxoZqTqsiOQC/MO/y0bqdTdy8QCLfnUflpN
3RWSbwKnd+Rz4MEifxqpKDZR5H9KqAoPPleOZ3Mexq0TM5p3SfT2JKn6GP+5B9Yo
3lE4GWwDlMBbe5GuL7zAnoEXQB4feG0DcmdT40QjyvjH0g9m5yXApcWL2k48DDsR
8cxKqGhfNY6SBuWzlU/tWFjNH2D4GO1Z2QkJoNjBdcnpiA0i2i54UqwtHq9HvsH1
ixWfcheg88IbLlC+BzedQHaw4bJu6/x/3LXHc1AaX/YD5RVeqVLLCfi7aV5eti8c
4XW5y+L9roQ5I3ewERxR9oy937dn/PZCabPG2/dJfi5+TmAy5U2zgE0dnyd/boht
N5UU73yOryEnDSDDt43/V9Z7/q6sv2jopQNlYh3XkI/VlcTEPHsFzl9MmBB7/WlP
bfEJLKvU77X0XaES1IviSnNUJnyQlgbPJH526IwA+3FuiPbReS9S/DLLbz4KPQOJ
CE05dHafglxlJ6ncjXISEzLE9NQSQq9Sfczl0e9bXefWIBzoilXEjp23amOC9A5t
dyn24wXmeFSXrjHTtueWqc2PR4RIVnCXeHrpIXBZaeoS3CItp/8iKY2WDOtCuwNe
+VhFvv9kFUGF9dDxGfTsEWUnoMEOxqs4HAv63loolZ72bOvBvgSoQSMhupVpNAI1
xiFbNQ+mDAd/AYP4pkYMQ1o5TLTdQ/CAQwWGGthMHrTEmSIse2u+R8z4xPME2Q7w
S4zUvvy33jvV51NQ3GegSBiaI6/l4kVNIzMDxsBp+UFcPMn/yuzP15f2oNxIsj1p
Gad59bDIF4W/qaUfDTPTzflAknjp/PwkKnuHpte/juDq9TiWfMSEumsBtdEfKwO5
vnRiVfK2lm9+o3HcAHiNjk6ui83fMtKyqDY3AZT+bo0kxHTRQVc+UyLFPjemWA22
+bohq4El1i2JpU7QIWqyPEVAAu0V0ABIJlrimrtE/X/NQx09SqJTxFrBRXoQhdx9
jcmFDSpMg3Z7OclyLNRuRZkH52b7pGJdONPTzrvfO1fggO6C7kk9pcMcX/p08U2A
lOSKhxjSqOhQF9fbI2IYTlAnLKU9Yuas8rsH96A2pfvSzAGC/Tm9iKnoILgygdF5
soimpw8fZQBLcw/mrVdUbkI38VTeUwWNtG35Dobcbze/v6fjDm2Po5xX/QcntS7Z
mdztGUnoUHdF/dcFRDyp1xwfpEkHEHYSNj5ve+EvW/82eGvMrosthgC2ZHI+MBCH
CatoYA6fvIRb1sJqEX6Zbtlex+eCo08TpTwrqJ7e46fgxP8AEjUJ6plnPmHOIjQt
xWEGl2JF6YD0wYW4SKMNX7NRxcdQldce2y/59IgpCqpW3m8Hv7LaalhAJzcGhD7M
PlYt3tCpL6CfKbUa7TQ0OOtGeKaQqZa7QwqOlEhYIlBUVovO6RLkV3BOs5ObyF9d
3tEIzAVpfvMcykiyYwnG2JrpJvIF66rg70Iuks0UKOglpO2MQg2znRyHpc/9UMrM
vjADOCD5l7ciFBwlGwuOXm9xf9W3GEOc5ssDtJ054wSx8Kd7hVU/yYwMHUA9H6mU
jvpsIXkiONzqKm9hGT5k0bkhOxovET9A4848p9KHuKmzVwh8PfYGbiuBgQUHIBS/
fgf7MEGsCrzLvgObpdQ8WiM+7gypXcl9+a29E9smjtCMQOBNuAOxsTpbTwz/YKG3
EWQhVVtuxnnAi8l0fONTJOolZaV9Xo4cuQpJnrf5r9OW/CJTz8lfvDhv3FK8V+Cw
gnrex0DfazfkgWcAppJdNhK71NTJ1kwzjgHeTKEUufZG1zEt9/npQW3S7ypPu8i+
UcseRcy/bHc9DmBjhbz1yXE7WReBBE+QfwWz0aDz/q1xYKLP2tQEoR9h5BJ2Qi39
SVou9wpfnS15co4Fy/jKeM1uQu6VowphPVcQStazJ90QJ5Pl7PoOmLzA45WvIEu1
o86trfyuRbTxWQJD2dJc+lp1cfxZ2AMwtXHlAbZlbh7FCo4/QyXvmGJXu1cutqzq
ntqMbSPtrnB8pgNxzaAdkz87Zx0Me8Sq1EolCfSP5+t9JX0W2b8p/36nVMHYOT9n
6PZ43zRA/P788j49eQAANCl5gvrHn7+VAqTEHZZW67v80XJArehN4YX6qIsAi12p
qXP9QZJvUacWzKom90liMzWrdGqav6GZQ7FcpFKgsWYk0n48SIiVdNTgWVBetM61
FzW0PYRx5BjgbilVZMlsPuaKDdQug/ENcPQQCap2xE4Y5LThOYwQVUfoQoKj9zDY
3iH2VDLJQq+SesWBhrIMKJXjM6iooqvxdO7NEt/dyTl3tRQ4+gGXrh3Avi3Es2cW
f5uPZeMveFY1A87jCVF4Q3rTL4HngVCktAG+tUM8I3tXXcNep3gGeTTxO0G16z2M
cCQWqY9ISzf8nI72TrXUawpKbrlViQhPewHHzp42v1bAHdMzehliBQ/c8dEghtFJ
LYHv8JKMeH6GgcEVnFqDdvLIS88MOX6oOoJXbSCXrB6P123qdOo3/00oWFuRL1Tr
pD9EQRPf69ZwMhj6bhHsLoeMkq6aK1ZNeJPm0sMvNfgh9TNz5kbBRyiFSj75TZQQ
L63Q56SqIrxntU0DRrqnBI1bg/VjG+PWZhwxU3B6M0r3iuWpGw4uAnAYyWYuJlhm
FR/dwUuvzUusxP+kONwJxK4QrjoZtNs2/BQy8hYE6RvGik7DjM79dTgijdjgyelH
GNs49DBmZ/V5Crja5ZYSUfcpkU+n26tCZPK64yEohCBIWJvaMypGjmfTs4yifllR
UuRwPQfexkFYEHWiEgIDf7wq2D2U9T8lYcZ7JZDHcsWL29d9SLv5QeOAt44YBuF6
10CHoiGdlWOqWoWhWonBn0h7ma7F11AY3STJwtPGXMpuWJR8ovoG++z0uWvo7/eb
dxY8fI9we/6rtDmiGKTIE3RDXDZg0JK4rQKua0ThMgUtb4ECB8K0FIhFP5A45k2C
u8gQdcqTray52RUpxEqB7lXSmHJ2ff1gU4QfcmHfTdS4tt66W592BvY9I1dJ457h
x5P2ihWpwvY6V8m4Z+diKPkPkUfiQwpv85VmtS1bzGlmC7F0lloLBmkxEQXUVdwW
kvr3IZHMJe5q2gxo2ikTLS0YHQf0Urx/nQdHywaTH/lR/Hx3sa4+WTvhhvbpWull
9/uMhQCEhPIi5bKy7Ey3PADc+WvFucQKiuwpXjm74v4m0E61o/dK9dUcQOEe8zGt
wCjapHhTpDaz/JSVtYp1ekevM2nqsq2A+iOCmFgK+kTw58EvAX7gxGXauG9vgEIy
D6Z1S9Dbdu6t6Pu0VkG2PvRSPeMUYTDWg4z1wOQt1oc+FshbX1pdjVi4Ku7vttEO
7Pm0JVNlff5yJyyjgT+Tf6oKnvRA3Ek64nSTa9wHaaaBWRRjfpfPPw4M2h63BTWY
qSELTygqx5jwswdDH8SalmgvBnB/x35QEv8lv1UTeEewNErM+MszzfJ0wlhSUo+D
HkCWu9kP2MCxn8q0vEfSel2AgeFt0PDSXiJKyIkc2sxVJrc+fV400ZuRaz1T9qcI
w4UMmLdkaBNgvH8KQ4H5qM4+4iTb987UR8WbYg79bnCQGF8TxsqXCUSXZr/fEv5O
7fWTTixobdR+gfIgSSMwnGc/ilCp0YkVxyLV5hjvB062bpDNVXLYbnG/4quLu8qG
h3LlFrLd/m9B50aCydeKOIydkS8Wsf6Kwpg0rs/SMlYolkKNqya94Tw4fcpf4Jt5
F0JYL4leCTOa8UregxoDdC8EakWJdRBMwosn0XVoFGPspe2CrFVCt+bpzjhD0JZL
mf9zB2TXCErYU1ywSjA/9b7p7AIz47pdtPQTzT5DDHrvSGySiwT8BzV10DJv2Hwb
EqVfaBJuHx6HSaN5hA6pW/Bnx77r+4mZSgvJvLasjMzpO7KLwSACXehyeJ/7zE+R
qjqpIcq3Okc3pvt5OLzkVjkKFnYNFH7h0h6hbhTS9wQMpi256yJFjJLO+tfDM+Ql
u+IL1z7ubxkAgGTy210dDMoDsGAHgqpCKTC3qFOQHKTd2oIBFb9nxP6X6q3X8FrM
vMX8ch3Sw1tW7y0G8yJYV+djrt61SPV3TpIFwERwIwZpjqp/oHE6rXCmDiYzCoZ0
hqLnGSGiPUkdR6taFkSAqSA7RAN7ubSH42ccDHOcgZVU6hHcWearcVdKLCMRknX8
XY2ldMEbBEG1mT93vCV8KgWrAFwPgIG5HtrjJoyc0aZKR0llre6EKgW4Vt8He0/5
snHpW7CwGYFAU0uTGeTl8rr8nz10aRbft84zTH8xsPPlHh9wuPrB+TMv+OqQrZms
NRPwe+KchqZD5QDUwQNfMmaXcp31YKBucSv85UO4F4ZyJq2LTjEEx/w5dj7M3br5
QFEzgJ83gidzrpduf+xbbEfJqpPlDxm3x0HDoOdMJqbh9LsdbFvlLC2+bRY/cs/g
2uiFOZ4uUui0K9dOygufUPNAatg1/P/F6Q+yvWY/0b5Hm9ox8cBC4ohGrXgESSDK
BeQP27TnW75F5hNIQIfIhvTKkpWQKrIQiF3naJfvTFyHVwba6O7q/Nl7Tcip81YW
Rbatr/4O44Fkhz33oKPJh3BbCIp7J8ieIE+KN499QnUXMrEX5++5dGTdhmvWuUMK
OVybnf+1U/+gJzfQPc7V7qqUfOBmwy20mn179d1g8tA8t9A1/IpdPAes9nJqbpDB
DDb8KSE0yLZNHYojvp8CzfMaPeNKEOS9SymVqqHX05vVfiRH3EkqJX5cxmiyP6yx
utTcuvapmTpnUQGr97bUMAzp7MmBnAakvyjV7FKxvVDtkOQdy5yvyTSVAujxUlEi
zdb71xiPxsNKebYNxkY6xt1erSUdIdXW6KwVKdyk1gAGR6ZvAb5D+pZlq0JBJVKx
xy5mLvUBhAovTNLgcSFHaiLi8KE8M9Ki/W3Cp1GZuv98Eg3B+7/4ZkzdtLYYk6AV
GAB6ZRbYS6bRkaZlYz06/+EMDVA8sgRiWh922z8wFXf7ky1FB1/KWvQ2624O/Mkv
YQjA+JMmV/T38LE8HFAbvJrZXPfuzf2s3+GI9Dw/9qdHW8RcLMUDsPHkHg7Ki+lm
SqE5Q8jzLmi0U2CihTGjIfU/TlqIknUidvu1U5otnjoBMqGUc1h7vf8LoZmaZ2G2
/vQttDD28JJRmkY4KGStn5rCdGhZxuDJs/rw29degH2exNervxoN6vFL5kC99Aan
jY09zd8pzv8dcoON729wMlC13dYuzrWGKeYtwoZYADCwJcWIK2/VFgtpQqIrxNUU
RaUlVM9MNBd2Slpiigh3pGGColbU8uA7gL36Ib0QJSRKZ6mEP3/t8PMy9o7KGwBl
zSLJNFjDB1yzNzeGQJsq5bU5KC6YambbXQwE0us22y5oSWzhTerZFQVNfoi3XgcB
bcRJPsHdk8idYc6lt1RDwUwfMvcNrT8ihrCPe7KszOvy1axrBsEyhfPfXLqaBZJL
e94/DlY9uBzij+caP47P9rOEUdRb2DokCrTsyObf64yLSVTQl8YrW6rQI7vCruG7
wvCiruwC1cYoiioL37OSEF7upXqzTpK/Hp3aOvO2dA0tFkUabQJ9QE0buhRThn/f
n7eOG8fiK3k53tXCZ63i/6REGMSJPP1hpyVV4nq6K4djipvnJTc1S6DYne0B0RXM
AhJ+V7OwFLLLvXgDZbMBrYKi4FG4U2oJoIUTynv6qUVW1XxzVEF8S5f3hw7zfIcH
9Lp/BS6ByAMCcm341dKyv8+E6z5T1A/RteR2g4sA4XWBDnrNx051AplIbwySXC+K
PyT+PXHYnSIl484+zffiEzkiP4Ipz0aKTTPGQVAgeCmxYWPiRy0lBnzn4FXAWthh
HX/u8hk2505wOXg/IxfxCkKmtU7GwS+6ziXT52DWQL+3w7BzIqND0C1tT1PWfLzP
+f+qwpVSsb06nTPDC2rHfCbJjwsuMctVA1OqV5EG+7TOk8LjoBC8vsyEvCtTGJ/X
F14c/mhuzRqmT/mT3WIHGlcJiHbkcSxj5B4e47I6hml6QXtI3b+Qd7dR2KmNChw1
bUY7+1SK5AVFBrFMBS9R15l824eYItrPxz6mx2Cj3D8z0oLLiM90RiB0waXL2qWZ
GrR4JNVW3m5lr0AXlrPp6BkR9+QKcQxiT6UAh+JLW4k54e8GbKRESHZ4ZQbv4WmI
Jt0wApjK4bTeB3QRdA6eGBkb+OrYyoCAaXWoM8EA8MvlqfkjRs5qyxBml4lIRsr8
qUeuwKFLLXlUrHWfbGFmzsmrYf/Pbb8oejqg3zYRo5B14gRBl57aeWJrVQ46RrY5
vfAnsygKs5oVA/vnt5z5MFo85D4mbgI8MU1ZDkwKz0zJEBAXdK1jFtZiu3txCO+S
dt6kcRDrbPLQVQFAkoI9MKJMNuqam9RWjmGprF8hZJnTL2LkWX45riG6X1oLj8XT
CovjUTJt16Q5WjbxwO4/Hy3IGzSlaTENNfcxZCMpQ7QKDlENQ6FbwF8JLGQCXChJ
fNWzGWTdiQ+TmTrLjAnNHPa0k0aH3M3wU+Kr9IRmvB73I+PqzWp3it5wy3VZsszG
5ZjP4+2NaPXBI7Unl3eoOkmrIoU8UmdqdAt6ViGjqDfcnbWG4JkH3ueiRTwtQSA5
YvrJULqnslTsgwgTVQlLLA46HtSmngKW/bFHyuJcWy3/Fmp+gC344MSNGqzH1CBl
FOU+LzLFSo+WZny3LWbDob2gedeHNENcbOGcfMsfdYRnuY8qa8kX+5uhY87kM6wr
grocmDsAX5yWCARG2wnVAxUs0e7JcSHwNe09j9zIZboWu3jamBlFZaQw98miSvM0
9AwnqMigBIPD/ioIydurXOJYEOtOq1qUusymyxs9esluNZtpeWu//VrlLayc1H71
yETm1PF4mYaCB1mQ5KG43/TffJAsm2rVFMpmnEpIH5yFkFGdlvt9QQfr/+CaSx36
p/UYUYyHIyInZQgPkEpO7SJORr1XK4VEXAOxbXqNP9CtxJIk9VG76UIeItx4uuSO
swDeSv6GClSEEbXIqriCoYVzQdwYG+9vm9NOIyHYDHj3B+8OM2G4annM+fsoMiSU
Bim2Fm1Y0wGzk6ERiehkCjOHSdWeLcET39k/rSji7OkZ5wtgwBZHRAgRA4i9H5/e
G0+mL2DNw14f2TEmWwX2IIfy7FCl/D8K//inuKdPaZaiPhQnep0S619C63602w2s
3jg3ACEfJqudsP1g33D1gO9oOgTb5av7pmp21gkVurV3ACD1TLD3HXoMOZ7KBCB7
73soA17rDfscQ2+gG7c0IhOEnnIEUhdwedQZCVyczj5S8P8pOeLz74tD6k19WgGS
pgrj97rxNeSbiHDurcnyP9R33+w71ZW/7jTirSe0KJRy897A0KTXV5MPsHuByS2m
cUnxrP8gLv8elwwTLTigvR6Lex1EOpARzAIgT5IINaZ0IssdQk3BfNGpu2oUisBU
l/wtaTI1YEd8h2ePyUirhryi0hq01sK/3GCwKWHgrfHrYPYOD0ztNp5RCgTzahxK
sWxo28c4wPvaz8eXW4SeT6X42H8WW/dxsWkRQfW+VL17jCywohehhf8XZaKbjAlk
IU3+Cm3zXDU2CdU7nTtSzKJiQDXu6cXePWRBMSkq6ksenMErHM8il+Rt3ClRecWv
4lFQsu7eX4KVRfC+y8fdv+1MutrbFgXUqoiClQzR68HIiEWMIhkASWyN4Rd/DcBF
/CINL8D2ZKa6NzkS6aP1f5Aqm7FVJmPmyTvCn8LOZ2T4n9xuuEsIbJLv7RpdzaWe
leMYAn9N+QL7Atkux8QXzDrdbj/F+tGZvU9yuR7lQfaO2OSCzVCvjZPwXAxLzPLC
4m7o86OXwJysCYpZkeyqkrY+DnYtC34BMDhvXY0tFwYqn2CNOgtpHzE/StCuKcB/
ZBqDZso2cx5f9Tv2DQ7yv2fglUU/kCs5Cd+p/qzWAPhsZ5N+7JEoRIAHLS9BPQ28
PGnzixterD+/d+RoYORePup7nbg+8miSJNwwTiQnXlDG0zEdDRdimotfiouL76V2
Wj78sp4x9C5VLjZZHIBu/kefrCdQ6tx0n114pVW/SJUFyA65g8GICCVRQJtpOxWy
T0KSLxHjMcT5fMjCYBBC0Wf7v+TzzNY9Mq7plPhWNmU+INvOkXSHlGO6R5LxKqoA
1vOSQ0V+LLTIIoQ1I8ePUosdtRwnlaIvH4lxQ0Rs4QRXz+idVR/YH2NhoS1iaYTX
l/DvnwJ44yGKunN+LZub1IWY45eZ8mNB41Gj/87gXMnMapanM5RBcrQe44TqzIFN
UOLccsjtje1OSDuYcPBTy64dFivnpWmLeL6a8B7KSjXR8cmvjM+m6hCNSgcg/K0Z
oNDD3jOn0D6eR9yebqgBv/Y27NY+RoIczNMKCuNFjRQKSe/gV9cQYWMhz3dAyGI7
5amxW/PJvLK+c62uZV/B6wHFmQJKTkVp+hehcfdoFKUKy5zlUTgLXbr29Lqrvn39
FtSxlK/AYBwwz7G23prYXnQkXLTvvZjS94yovJ3YzztdBDtCvm2b7KSsAj5/oBTR
7u3YYg7vYi+9K6y3D59WMzsJZraMRWcDGBPyo57ib/IpyomjJgnBM0UOe7Y9sRwY
c6oAMVd75dzDunVu5azTqMd++EwdKBXkQW+YsYoPorB2p3aiJ29QZCUpV3iskj1y
NuE02fqEa7WqDcCjPm1lgesfoEFINu0+obfRohQuDL2V3vZnH+NzAon2eWEB5zK8
ZtPPnH7+PnlYJn3wtComu0i2Tst0p86Oo7xGsQYIVtaYUvolqYK3PxiPpJu+ZAQp
nQqDHl0z13DecUiueNgPNK2nVoCt5T+B1DeZHA5RBsUYgJuS9gOZ7GxNBqyH0iX8
ggCCp0hC9UXl+obGgcqgSCB7oMVXc1OEz+nllJbS9RtrvhTA5zg1s2HRAsYb5MG3
o+KkjfyP6hqMD48xEquo4vDUb6G8GiH3DUy7XO01TzmEHIEf8uYPdWlQphwvGREj
/iNzCMyTiQd0J/VK2QnSN5no//ysMZtHkGI41xlVAv5YSFXtBlqMp/8+no1EzL4a
HQlzoSgKJNyq0O4bcAxg37zcriophoBsj2jjpfMLk4O1jl/6qj8OyKJYcziPpqcM
OS8N6720WWMIaIekCDkKWyqr4p4hQWgG7CtOH/oPfRsFsZoGz5RteB/A18n+jhSA
nYQq5CBG/Sdl7y8LeAPTQ9gl+m71a/GVHV8yWIbO+c8zwtdBaMARIf69w+LRvEio
y3h93uTetkVIEm8vsOPnZ8fben8cv4+o6WL7kCRn9J1eLRNK6fttlvgoxGmQLnww
nMsHYRT0LsYe1zAU2Uq3AJ00ZzHgbBNsfAI2efm8cAvUeGVbYwrB+CNpkK4M2Ztx
w+muJfJFL1YXrxnK2x8MqjQi6lT3AP0HLpGmEUXnz0CcD4G5Is/mwkvKfS+1WSC1
i+6Xac/Wg3YfWAM212gmxOk8daZ5LIf2LXR8tEq+SEJvvyZXVcYoPa2Kpx3LXuzO
AFWwt5scGjNdaaFt1g2W94lKWZIuxXmzo7+ZVsuxJ+a2tLCGJg/dVDYg0mt+olo9
RYD/VFlEdbnCqxP3eUPxJK4WZoeaU5+wwP9CXsbJoUDQgEaSc6uSiue8xs0mzGrn
bfVth+Q0qBuCFxICdh33Qpye/M2fJN0hRBEbeZ1I+X9OCh9ukl665ciAdaaKYig8
JzD+adNzocRH/TpBGv17LQq+ijYAzTjxry8MGUCLRkv/py1oqMZLHwaTQElQ+yB1
/FWhUoLsdXzNH9hqpj58o7Ol8bxQCJ6/yiCZrBgg6OyFm1rh9AtF93VkccuZXQjj
EhgcC+XU8/L0AIEqexJCAVCvhTAs/JXWDB4fNS2J56hdRzK7CBFH3t47MZXSIwju
wkKMwh6c3cQA3zX73Ri2zSLh8XgtsmwTdthI8yqmEnA5qkB/OJVOcmHqKWitZzv/
q+J17HOlMMArvY7r20hACvaaM1MMR6yMksyCSu2JFeDf7wxbvAEXkafSqDIXVkTh
J6kxPQSLxLtbasePnpFpZx2C8lYKPG4BEgP2Si28li7h6l82c3L6qlOVzs1B3D+Q
kKToW46PmpPLsGPVkovlvs7Ee3b1uophl2NaoRZxeOQE7fHe1RVl+eiOzx+a15OV
nsCsSY8Q0epx8Je2RKMn3WfM2pnjzWWUB5RoBdVI+qQqHs/LlldJeHvFJgRF9LrI
A1L1UrjPA523Ry81urqHWRIkGc7HMmxbumCA7xWnxKHFbqSMw+DmKyHZpMk8d0Ej
3AB4j4YQBZGih3ZS8Wlk7P23aDB9NHnAL+5Ww1mafI7zEOb67hwrOmYSMlHhEHhC
lxmDuiwWS39pv1bAj/8PdgEviLie619O3I6j3DvVZarpE01J1j7wJ873sqrUb4zk
Pz6fgYtFfVTnvUHJ+GEMgwJwP0jNnjZ5qRbisAflSKbSEeoAlM/DAMTcfRYJs0OB
LeoXnbfxiYn217XrfFi4P2OBJpKqwucV+Zcjuvc4yJ/TvcgUE7QvdX6JAZtagPF/
NcwiQV/g0Q1L5sVyGIFc0lTOQmWLYy2lXxHzy9XcCh5q+/w/mghhC1SWWxTn6t2c
faCOobUVJ9GU740hNjnKwNrjDqLY10JHj6BgBsYfAQcnVW/hE8/+VPWsgiSwY8Oe
mDIIDTgtLlW4hN+RmncKzvpCQ4/VSxWIbodGF2pXp/garCPaP7B7rtaK4bfm8H1s
DEloBne40yn8i45ro4p/qnJ/dFnDUhA+hkdc6yBZi1eZEP7KzaswpwWLYGV0zywZ
4/62QXCbOHmLd2Un0FSg3ZnUcgNHDnInPquybrUJ8iPGK/CgN/lJNYvASizKcIly
nHJOQxe2ytj/kxFxBZBb21mVC+jQo5kcEDIPHMGWghuCtwBRXP2m//dcpsvxNbFX
p8eB7Cd+aiRhTtGfluD/HlczNWLw7os4tl3RVQFI3wvBakVdT0CkYEXZTVwSiyvE
uEeK/Hc78TUmX6wMHzELTAyKlSObN3ey8FASXRCK6Ne9E+4+RdKyvoOlJQdlJm/i
Y54paDTtV9dOfWs5oDhjEjXMM7h7j94mJUcp1mV31PIOlgh2IJDUpFIEiroJ8mni
43SCLkitcldNNzXwc4gxBDiTCqey6zwDy3xsy0XeXaGHsFmMqgmKLHQX9/fxrY+3
SKcnN4R98LHTgaQ2rrZWoTC3CMrOvL2P/2mk/2csDdCi+oxXYCkguqDtnpa1yjeC
xjQQEEOkw4vUK0+ALTnXDueLspkYdvb6EgfxeVni8BywkG0Q6pyqE6tUbCeObUta
m2LKS3OlRxsPP3Rzagz3+2WysjPC8HRiI1zwKqURNMv0wDX324gznhKJumwP0T3i
N97Ur7zIJUqgg0Cvwp0WdoZKv5YaDP5SbgBTS+imwwuuTFwxp+5Smg7ztW7TQGQh
/o3qSiR159f0Z/WIy6gxvL2Js1a2nA2RiR+ionGfVAiMlu53qKBfZAUNvbFCD63I
WiOo1K3EP71l7oU7tVNOzQZsjcdLvZz+/oF9v/VvikdUZcnJ8yrpeFZPUKCS8J+C
lRTTBl5dgXOzLofgJNHhbipUeyuklTNVxqg3fydoQFcV66HieoOE1moQub4tbtfw
ErAO7jpSyw7Ebn6tMlBlG2QH4taEg88qD/peDA+AGFNRSi94o1kyPK+4w8r1BicO
vnZIrFCLSoF3WAEy24f4PUUwlIJWI9c9Td61B4rPDZ6YWRPs30hLSGrePARa6+vO
U6ouz6yMotlmRlouRzRV1OIasL8BMvxrZLFk1P5rzBWSmmr9fKVhdwnHQxZ0mG+6
ntdV6ZzDt/gKdn0E7Z0yo02ocXIqiRRkvyd0k0mQWWeNPh+Wi2rEdqn/nB6Pd9z9
5m/t2nwRy9oL1hwwnqblJls+EE7vitPJyr5swfjmHVKlLh8egSaTje1EeO5Siz8P
7jMsdYdkoo+VjRziJazVEuF05bfdPBIroiyHroJi3pKedII3+ufqtBmc2Uk0pQPW
BVvHrBFUI+a2DRGol87XPdeW+lYgf3fkDcIeivbnzqlyHQ7XwjuF2bW1MeM+sdpD
FRuNKvIE9YXH5hdIgBrjBMyxsCuQs5XdBoZef1fZ4bZSntfBExQwfkl7PH+U86DO
Hzcvo3iPV858C/a6kcLjKMegzRZCCy7XfMvlavkeZTDj722LsfMTUp681RdUznrg
yveg8+MEryowHxZIT9qOA3S68MDnNB17IJBaDvoma/cfDqoN7HBWVnoglBcPlup/
xr81m4+QJXtzpSMNXYl36QSSGrisiR494BJvsdN+TZ79yCSUMQ0TyPpejiCxGJW2
pxRe5hxmiUbmqkF4S0ZukDM0rF24CvE7EsU1jKq8QCt2B+L4PyhkDpynyYhlm/uc
HAmAFJKAUI6JEguhOUwZm0Ln+YkMvqLIujHLBuOANoLNjajVSs41zvmVuRMghNQz
PmXNXr6bXnYPweyWN8JdJW0UMSo08ByB+ZiT87otq9/TCGUmqFj08AdhDKzV02hS
1he4kx06MDKY16SLGJ2qWYJgl+kL9tP3C7gehCVgNU+NdABX49mCo9W+fh6DIBVi
/FKRSV0jv/lBbGNhobzQ04a7UEKa467xbIwWxsugeZJOi1096AwcUfVbczyPU9yJ
sTDVPMVIuFv/x5Moi5I0zetX1NS1HxR+nyCylADS/zucdBWaX04psVsoIvvTZHZ1
acWVzeRpH0yTUTBCPfXAcs5vLBZrmd/Dxs2/3W6iX66GxF6KQe2+oRQxFRD+TCKd
hiTFChE01bItZpW1dHuYZhzk90XvNj4VcHJ7wuLL65Xon6wBMDunqx/R22qUBmTp
LR90CwN0R8PBkmtw8McfYcMVdj1sSjUyuRevma7mDw7lATgp/fJX48ZtEpVfNeqf
GPUkLiKBOgUH059VMNZSq7UwQ1TQGOmdSvwuBWT+mN1cIjX4tD9w/Zj+8BPjbHxC
F0py5r1rqtB/cTvJVSxvrAwSyo0B6svNoECaI54pE8XWPVTXGAUdMb7LAUD90P1C
Fj+vsZFthEBBaw9YPdhYT2sJdDlGN82TVz5WrcNfyLDBOPRwMNSvXPTLjra4RE27
N6bVAYmDK/9c7SeDahDiD6f9J3O86G2Kiew9QOxdhes6Nalup0GZ56RGwEm4kgdy
6EX4YcF6oL+SLNGi6jlX1c0SOksZ4b3jlAC2hYSOpa48htTVsPYjJEdSFsMLJWAw
aNi+sXJ2QB65ZmKfQh9ySxCkoMna7BNHk+PHmgjKjgiLWRaSEVO+1W9uk/u1BPh3
70wCe60fdVpy+JP3bmPHai+bJjSl1KB804Bc3yYq9YZ2L57VydE3N6Dd+SsBp+xw
pVAzPXlMdFv/ZmHOQxo7xjSH9J+tTPAyg4O3C+97F9sPy7/7qvc1BQ69okFRHcgW
E6YH2R0TkUkAShSPW1jE1HL0QWwf/5S0d699IKRYY0X0FbX1LQ1e0863eKHfmN5j
0tq1esIhRBuDFdt4lsG5ufwdPqY7N/I2kL4jWvVPBzN+3p0YHFddHjDlZq/uYEO1
zAckFeZEFJCH4fAG3PaazkKBD7K5w/RQj5VlLAkOXirFWSvCNhdOcVlHeBz0Dp5f
aiRg4aQ7fbWjr/1T0bZS/qVbfb1PFtMeeIAC+2hSN/5rA7996xAV/N5YUC8yNt26
pk/XMgyBoRLezU6CKaLF5hs6AuuLRfbUgFF21cBXaMwMxPbfQyAEREJfZg8nVdI0
Qn8DyG7B5+GiDQkCXbXvMegE56RwrB11HEqxqh9JYRQDcf/+HaKK02dAWcaPNHzb
YbYeEFKcmBHUI2ofORWivQWAHTLrWtCGM+7y0H5hkqBglh2zPU9Ag2rgjCG2E3Qk
yXoBTJ7RlA5bWXVFO0XusK/Bfc4cv8xLdgU0R1n/YQeWsIYuhYNJq/6lRdWlSzX8
w/rntLPTP/lpU44F3ZOIVghwyyhGOrOoS8poWOL2KpLAC/23lWNXGpt90/lFII0I
m0WqgRWsn+VhLuaMC0qzMXd98p16wLJcEsJkkUKXrB0SkaT4hi2Aw4864XEaytY+
mepjCIS3G9xcRXkl4/H8/bTR9F711chvU+2qzEmoYj+HAbXN9y4uQ9Zcrxv8uz5G
50lxv5qekCpbF1Uwp22pSfbPECzIISmLoe2/7k9AQ+eJP5JU6OJViHSZzAP1bvAD
sx8KaOEZs2y2D8NyC1rEzoJxDK8NQuWGu6FV38aeWjV/TB975iilFLZPVYAG3xU/
uBT21JirJqkbEOnVIj0cr10bT0+aMGXe7WMbi8Vt2zphgZTz0/faZqnBUUU6p645
Bv4+7yrSDsoqT/q3Lzh2vdMd2GLo8u3HgtsrVa8bHEvCzPHQdauDa96mHUAbEACd
IUfVWZPVcNUE7rE61G3HyifXpB4VUl6gA9kfFL084Qk21TkHwiSWPQLenZtvEHBC
7Z9gq3OhyY6q0otNOdHUihNsOFhd1A/6EFnuL+76FsgI0gcUKh6VJ+zVdAqvBsDn
YNuG0sPKHauOD0HmegIgmF3CW10ubDgGxRuYFdiwT6Xoz3HSJBC8TICZ1yseOe3U
MrcF8pUFlVxJLw7fX1IFvRoms/j4w6VRjMkA1JnpYKgcVfFPS9bdCTcTim2bLTVz
aF3yuuDO/P96/BQQO2ZEaOjnh9dk0b8/Xjq+OE6JmSH2Q74+BUZk+qeWuaFx/X9U
cJv//A0i85tp3MaMJ2Ru4kJDMZMLIwEKVlVO59Z56c4DXhNidSBDBiiaL1L2OvZb
fKIu/NI51M4vB1bFZYe/Ycmzf4hP1jMuvRWf4/kheBA4g6LI17WeA1kxGPj3mNw7
dcaSo0ldn6ktqE573mUAibNHg493xkJoLm/FFedv4HaRbD5UyO0AjfRNcuJj3d54
RS7iuA/0Tn2C4LOCazz9IlUjndey+7LULek4euQnndjbS1OrxPOis/lEF9SreXMj
0+VWUl5ExkLU5N3SGG3C5V5Aia7LnkmKAti29z0xykwzK5jy3QeROjmkXSgCy4DC
akOkTJHA4KMMk3asF5iJH71YdRfiPMSu9l81igPXZJsQqwrXDPJIh5iVwJmM8TLV
WNTkvC1/ri6C5u+4I+kFpWxsvBUv+cAJs7YrGhtDsWjOQpGf0ttuTU/bH2rjrc86
jPmfeqVg0pRQCGXQSw/EIBqRqKLSh9DK9X9a1Ka4OooNgeJ2uIrvlC7qMmy5iM1F
Sv5X4qbrlwSz7TWBVLf81m2UEzzbrkOS/HiCndr9aljYiJcK3bOcFeRdjCddgKAL
xoC+ceZ0RW6ucn03zV3VM5aR7amOZaRsevlgvrKyIlyNXQsfnutCcclc/cQdxoxJ
3MMPCqO+q7ZyLmCiyHK6BnbrJyxV+es9L5Qzw6/J+5N5iRhWH9uXywRevesHbB3Q
HtUFevNkgCGHOq6quDbIEZX4l6HOLNa8F0GxNV/+7fzEtByn6wtw10ZyXhVYUbXO
7UHaM4oHzD1CLnSaN7Hbd63xAkeGg6dhiob/YFWfcSdTWvSLFLHToEOwCNfhifuX
2X8agLN4kq/QlG/xgpdP3OSiaeekowLI1OLM9nhNMZD/IknRFNlvY0wiOaUeukbn
66pj0dvZLoglrWbia4Qw54DNYcr/hDvGlJStSBYRBLj4KeEon1ZyE6OhhzkkVq4Y
36sjMdbqodiTcgCgr5V4PRGlqMY9kNEgXjpFaLKgbJApFD4xNg900GCX1eVNdD7M
sXsGMdhxpYhyxjyKsG2r7XjZtOHbH5+KOsE5S/Kc0izBggIT+hmcikW0mQzkg1f3
Q/4TPkRcUYbUcYTM7TyKBGVG+tvnXOtJz+9xqGJ8KizvoF8ecr/ZTGiu9+H1++/k
Dii7tzm7rah8cqSr4Qdcthc8EIyFzJqOUcNutJPD2P59R/wuhcvBiO8ev+MJwjui
Xa8kAbtoyCDDfzHLM8T2Rw8tpdHWoEl/kAJgmnkDSlNEhtOWnckK0xShyXHvflmO
5W9LLjjBqL+pAhKAgnkd6+hLj+7hTpQp+1w/UGOVkZxjocR9iypaJEdgx6AchHHO
GZUclZf0RGuGcWfWe2Op2gG1JEBSeaS71SuBAQG6o872hxWcJKqn1FB7K/6MUnc2
u7zh3b4/Qxanu+tcVlyDsuBw1fSZFq3ONVx0o3QR1izujROZFhCFo/phuoo97K/E
AAQ83jcN9GaWH2OysKDRktGfZ8wM6PXgcQcp0HQelKCCj6jkMmXOPfoA261usJtv
3O8j0NV11WApJX0z2ZkRO4FWeLjZ3TMpKFNTdB839pg/dcHpF1Knwd17+1uhVmI+
EpAllwT0hnorH6L+7J0ZxQICUcdeo+uaBKtKr5N/mEnCs/Hzk77NFiBvxBMrrBih
mGbgbRymqLl88vACkBeLqncN5xD/lEjrcPZ3rfvgA+MzwXOa+uWDT/e4OyP13GpV
ofgJWzLp14aY7dVKI9Lz/CPq0NxIyVXBLgXAuQo80PTj4U1HgjO7QZDGRnBjCH8L
C1U8fZoljuEk1IR9JHTGdHKTm6tJwqP2dPDTE2JdE4XU0qPkRqcZBWVb6Y2INnen
hoyqhp7QplgIHZkHo9yAphEKFeeudI5KmdWeaLh694O4HXro6ZVcEAHK+z/ccQ9I
Drp/Smnx2GDS1Yb0yiiPUqsPuigR4mrBex6GZBpaaZEYNEsfiyNTbKmpV0NBg+2M
3PtYOnShWhG1t5Wcd5TB9H/vRgyFQHmpjbfWd29rOliZ4d7mcjyW9jgxqgeWZwit
mggVx0WbCOeFYnFnLWc3kFmD4QmwLFdlTELYVKVKysAhyBVJVz0jFJeGgEk7Q8Zb
FcDgggy2b1qge2PQ7cfUjrmY6dTwTdYkWzCiWM6bE/HAxHXRzUgboOcAk75GYb5l
3lzzeCXA6xYsdKMBGKwTRMXYATMX4cKzYkkE+sXu3rJC2vJhix0BsCcXbK84v/en
VxG9DZBXlEM1UxZGVNvqhioSi3pMeo2UnnAkXKy9ChkUoiPjs5pr09mnvweCbuwU
upcrHh6KyGoBJVjVNnvY8ZWvx/yDbFPi/bm1fwAwKoyFHNkyock9SJFSC4PDrcB8
TOPhJsUdnSUwvs3ZSm6PBkmP37CyyFWegrm64ZtJRuouGs+eqqCVICvkfWgM1HfQ
Q3fa59Q780ovffqHwDQeVCJToX9/M3klNugyHdYrJSciijb6VY5cjV3Imbi6o62m
jABkVZXLPk+Bh+cl7ua/sbzQuvicTavlGbG4uubHZf4RuiZWZ7yTzt4Ls3uVUUbw
voppiJE8286MUqUFwnV0FzuknJmFDAv+vL4RB5K98V31X6ZKmG1y/c6uIVnZhQ+A
OAAGqV7sQXdm9WBGYjhrZdD8gDK/dnlOLgoNa/D9s3hh1jshFuoKPgEDR9HiPrlU
Rl/h0uag2Pk2myK0KsVwckAMBC3szcIOby2i35z2tiKeQrcdR/6ge4uHCzoux7zv
SyagHZafF3p8o0kEl854jSsBkSSQm8jC2R70+h1Jov7ILVDIiNtQzoOXaR/61Rx/
6BsAnL6n9QVQ/LL5llk+cGQ0uXrwk/EukrgOabhwuxKnSmfXjm5I1kfqCd8mM08E
/gr9QFdXV+bp9Hjd/VlQmlUPnPwDa5wJo269SPsBltAY5NOuWKJQZN4UpfSH2NM5
CfhwVbxb8gbyqMMtl936dsTJ/iOhO10JwfNf2BPwyH/VsItrilwOjPCiSTJax5T7
nN9mpwVWFcayQQ5XGfcdEsobkdA3ODe+FfstwZMgp4qP5LnqwQTkcThbSbKzcv5w
3D1bV1ytD2Ho4GGo9rGU4L3NLmbWwGlUTuYRRfXHJe+D0wX5D48N1NVv01WDkPFX
b9uBrGvh0NtEELZG6AzdQ1s8nbm6cpvIR9prGhv66zbjaXbsUASE+apgKPrbW3rj
SmJfnnnt2MyJQTwmt11yqhf+c4OSWVK0ABRXpA/wvALLHtUhg/kxK6y9BS2iUnXT
xee9Px6IG76mPGYywPI0uYFC5iwEmM9LyBpf2pjElxsbb4+NCv6o3WFPKvcSBWSL
Z8xhO+Ep2NU70Hj7qo30cqVNtR9SGcBedZFSFIgQV9f7zPC3ZkRzexQXtTCbqjhs
yB73y6+5jEmG2zasIDXfWfo2u8mkrET+seC4o38IiDJYOJuBxRdTViIhwhwuGG7j
VBF2MoVE7srAuykaMKfCQ9oRewEfdbV9DEYDikjFUamiZidPbLXXSZnSHfTNaB5u
JJO85Un470S2XIZ/GjIeBF1PwfjL1kKDNHdSIcOck8yWpPMd8KxrBKtT4QpiUEjF
NoZfphnqlMGnS0Fna81hANZDj1/RNi2SdiILH/93L14pOq9O0C4dLW9Y8QRSVklx
MFtKaSrR4UwMpyOCMxySr3AOajwagNDc46kJBXk22B0KWHbM4PMlTXlRxpkkIDRR
tT5AmWA/HfPA81UNumBIhrkgyrgnxVb/qFyB3NssA7aZ2OTMeOfDSVv1F8R6kiAp
ilmx/thwbp+JcsL7az2GyLijCcZAFfT5/AG0C/gDy8ea3hPjvOkkNTipPsCrVpQy
RiF3yR9TZnR1tduqkFSjuE4DqM0At60CQnK9rG+yNvUcateWFIUjUTWzh0qYiKwI
yZArTH3CnhMOKr+EI9YBTp3G2dTWfcdZmQ2Y0VndqUEgIr9VPk+26hNEATOChhvQ
aQ/JVF02meXZn6RhlRVoVUKNa05Z57QPM6AIM6AN8ijXCFnt0z1El8lDkPX9nOgc
sQJ0szZfhJKpthf7lDfp2y+yKujXHbfyrkjwwOsy0LHIyQ3/u4vdmBqpkGWZ0OVP
Px0Dv6wLavSPh83+XwR3GPeWAWvr3ZqKhcc3l3b0mOdlL9SIfc86U8RLiQE1B/IW
RNodLN7AsMvYP67ZirLjzHiCQ/FFDfP/ckmCuMgkuXtSRqSIhd/HAfxwFf4Pv/e5
PAARZTCVd4KSH0BLtg592kLph/ICMR+oPaVohRR3Fb4HYr2C8ZKrKUbBp97JUnqY
l1aGuizAsG6+INGUATH5LQ6mxIo8I6n1jWLQn2X3SJ+6NX4fSU6Bx/14GVqREy7B
vJy00Xcj3wMcRnzLdkrEysLBZyRebOGQQy5TQcM4Y5oYMhauksd8fiC3TG0xkio/
z4WDjxnv6Aer4mpIZ4menbQxRahDxsbf6Q4R21LEGEsICUnkMXFafiZcCEwVmTF/
tmyOWYOO40BC+cB6+QF5r5Qx1YkK8WeYlJtHpMhTuyuSqg7oNBjimOR8hAGPphCi
9aEbeF1r5pngkMhmXIyr/ycoPbpFexT4IuWSRnkrtv/e3onXOXDy6X/eTJrNdQuV
Qn6WF+DexKkrjhAVVkLcb9yHRLjh+M0v3YsYhnttzLOY0PvClthH2/5dgf99M99J
B20KtnVLVVmowhH9KO5Z2T79YiXNC+NSuSFt++5VMTau8UULimlGgWeaPeI3/lMZ
PlwfvDr9OfTkcr26H5ESCJ68jD5JNAZggb51NBy6XNyqRcurvj080xT8ODEVLpat
AIBTOWvap86JLkBnMW7yVDRZ3/yx63M/i3hlh9JNr7IoD5FIDvvSK+k5K3o3MpAG
lC8pCbEfH709tYY/L7L5sx3k3F4wW5dBwGLfx8YCWGANlgU87QGnGCtHB73cjbhX
yZKUY9p1qX66Yh53PW8PuH2vDZPcztcHIdBU2HWVstJzpY6xRW0rLaUf0N4FOYlQ
RGAVTUlAwjmC6k10N32MlMNiwRm9OI8CJBrwa/k0TuLvGM8fNNBH9+V/4rd2TXNs
yn2fb4VB3I+x9rYdIB8JDRVy+5Yr0SWkEqGHDHjR3Pk8cA9+GW3Ld0i+5nkc5JE5
P8eWd7uLf3EsDmlGaHddQIyFJeEkEnI0tOj7tK7XZCLYUXcJnoIM6MbxHEaRyStD
6WuejS1qwPkykePiY8H+JVs2jHNJnNc9NZAsnIJ6QmsEtdza5GptqSsZ9ydZuuU4
X+b0De92biRArnDudlVceQa6H/jvJZVY0IFRO0Fgmdza6SjSw4iVSf/zq7G7+MbW
EcD5oD1qiLzwO4YoEM8da7Gg6EkNAI/vzCMEghVCRUenebolpvZyfAEtiFzi0hQl
j6v8KLD93JLZ7Ww3gIwwxW+FVjX+ttlAxSI1hEvJ6TDWPhxjSt/RNwGjveZINR3x
krjjRL82z+p4gvmSYt7/7rODyGgxatiKVtZVXTb5D/Go5RviMElHyYPSNKoEC4mj
LPJPEFj7vsje4ZyftlSpdwNZewofiXLm04Wrp6iM7dRzAw2O4rGDr0hc8H48eVoX
0oWfar3ZqWLnw1rx5++keBVYCGvy5+eqPiZ+aRw5WxU3vY+Cobn3oyXeUFO/qc5P
Y/gxTM0jkkgxoShvInPGqhHyNa0+bo2NXMKe+2JCjSid7sShIIqPa43rS/gTXMcA
7flNhomDuel8pGNlf5kHIvyfe4dg0Wg9phW6rzbQnzR92rNE8ZLY6NmUXgKwLuER
k7hDCEg2Htl8g5wjgg7O+6Zm1dzUsFtqPWnBWjg2RP68oWK/To4iVHHa6eGBEeOq
iPGF8khw5nZWgjHxkmp1sU/e0qGDVvZoPTY7rbhwKqc5DeFqRcg8Yc10trI1QpPF
Dy+XcMnlMYituw1H6MheVY3E1rIp/FLt09nUbVtOchEB3QuEQDwDB5Iup/IPh7EW
KHle/Pd8ezY/Khda2I97Cl9CMvbmxDo8uBV7qIhtdqTTdavbeChRpLoMqYRjTe3i
yz1xKA5PZ8Ih3Mx+DsIoyfGIOZzrYvtlMaEowQHuXPhQZLNMYVtwOlNOKJkYPGtx
oZuI6GDpNjOI1tLXe+HGcCiPOBRxzgjY4Hn76ZizrL5mV1XcVaAEN5grnbTBUA3V
asuY0yWLBLIs0Sr2POy6bPUC8ePm566Vuc5I1M9aORvnVlIFUtShrdqNnC/WoZR1
zcDU5z+iNf5xn2SxE94ucMAH7V9ymN9CUWUyb5VwbpNorQWeOh3dU+WhDJ5KdL0V
wU/cB76rpu2SlGHebnm3xI64JfRZaECNDlOxQpI2QV6PCkcy/i/7u99+Wo4QuPJ2
C0RkvecjNG39PNssNg+CHJznyQBE/6oJJ3L3urNvgwEstm2gIRd2Fvp9YCSexsk4
uFlus+hrsVxqovWm+XAj4Sgi7fqETv+AUUzPFXVtGddYTuBFBjKNFtT96Bpm91cU
MnIIOUGNGXc5A74eNq8adROvYZLmP2yr5mRFZvjAz7zhQvPtb6IXyFgHpYswO8z8
mFnnpHZdhCw2K9ALZpbLLhd9KruJukoQ11pZy5oQ6vpCcFNVW06zoY62nAHYNATp
dZqPbIogSR/gCWNEhjWlpngFED4+AHEn6R/guyhkIEx0tZIGlPLB7Ct6XKr4fTp1
r3i41EM57f+ZOuvLUrO2sEhyX0IrCRQjoeg0wAFU33+cB6yLsY4QYfrSzJcXJPGd
NCuEF74ubTxlWzcBtnc1A+APM/hCat16aBmzR4NpLke9jB0aFsFn2ppsLvC5+E4H
ed+I3tvWT/NzxXaHyjrKK+FUWL42p3WBxj92pZopzSuJBAyUCShcA6tKEBrd5uuq
iD+CsqfjqnRLA20eFEkLm7A7HQ5EuWgbL7PSYBe+n/uV66KlUxTM6dBqiwy21ory
16PxtpADQtcEcLD/W2dOryoxyFfGf3VdAP1G6aA8XNMsw0iskWCsX+fxTUB+SNgw
AAnOM4Ro6ik6rxbk0qWtEaQtk7Z9Hh4ZY6mk0A6YDb0W8155NtJ3Ax961Yqr1Ng7
SBfDgR0bTiZen6ku3+s+x4yMh4BUc+T6ESHx5kW1z7ARnwYtgXt5/e6LhJU1czCc
qEB66OXBYYp/RlDOM/uC3MNmbYQhj46BZ8VlZB2sO9G/i4HygyKCizOfC5CWcIUQ
+c7fe93WUpyOBiTUxlUump6hKL8J4XmwnBLOnEnuq4YskxqJDPmOOyq1BGj4j2oB
xw4Di2nQAWXKDCFGNRddMrBwjO1RXZFfLF59uw1GA3yfZQCtXfjFUN2Wh9CawE62
FjPogheuPoruyaIFStxG+E479TwYetBwptgzJU5XHYvtH+qbwlz61x3mIK+QxoG4
AuWNvTAoKJm4CajqpqUN+Mu0E6MGEQ59M1/H5/oof3jsGjBFeeCk/xQmkcG9inGu
3OW/YmEE+VJqoW5eN7szfNjDtYLtzt0p7oIJBsewENMlO9SmqlBTzJQrrCsQwejE
Sf7qtzV2CoYto4w9dufvwjkhdsdC8qCqj2KwdZPTfNZNQ11VkrYPVh/+2F82ePPk
1ZswLMHoW7psGJm04hfzRIO8jQ70q0u3m5KOy1gJ0VdGjUM8L3CkWX3w9UmouO23
h7lMpiejTiPMRP9GZYeMhzmxDERJ7GHfjLsNNoIgZMB81FNdMVy8MWv/mm8f9aqa
HPSlHXl4XWfmgjVymKuG42vZte75j5RrbaLdBnJV7OeiBSBHR0XfTeenjtpsk0Sw
jYQNvv3yDYdaS++JBaJwAYRqS3zRdw49zR71OiTD46j/sg+9zzOuFjLXnNXIWqeR
LnzCUdQ0dAIqbiyMizwp4d4PRZPLepWmC5gyv6nGc5HhLBvgAow4UdqrX5/dTggH
s2g+4tzPLG6UeZPtnTVOEltN22gYXeGJ4airZ+BSBN1T6dGaGMMQmVRXvs5uxZxO
4535b7Kj8ESGPh/EnqwzoR3iSh1SzwHCg1WvbXSX0zXd+NqbvMXlhQcX9FWCJ9LE
lsfAHN7KdvEmVjkekvF2TzBScouIk2WVF0344+Lwu01QCbe5UOfZAm/yJ6IoAeG5
yCCK2gZ/Nrmhw7hJSNFpQn5fgtiGPJbj/i9X/Wvg4lFrBfymN0tW3Z9Y966yZtPX
8Jq+z1r26ui1u/7yhaVkcTQ8/Xhl1UXmmuIFRoiKAeMnYT+PV9p3RPQEoIMhP8Vr
3cGU7RUSQyBxiiigBhP9+u8z+psBSbdvFw+HBsSPYwG/QUmqx2BEO2iZu1oQDNdk
F+tCqOy8jI8wAn2OxdkdkgVCJrl7P0K4oSYhNvEp8zAtcIveSAYqeyKDrGAIlJAQ
pHiYEwt7+QCOldJgGTo0i4duS68lLN9k1cBx6FjbZhc8EzkJdg/xXUGA6k9Xe6HR
4fA2rJR/sAAXHPN9G6YGA3LDjSKYuBPhQopRsnVv1kaciYVsrL8ijURsduMdbJTY
AWtO61A76vl1S+2T/W649Npw2UoA8zOIa4QEiIcNA6j87xA2Lnzs/72A/ylc/XO+
2wUWuLHQH9UmW3YWuoeyU7J4FXQ3kMQSf5T52Q8zuUe3YAb9IapgH6CODOJd0GCE
E2nyBW1LhJXfdn1sOmrPuhEFkMOqmgPF9bCsKKaK0qw+/lxxUs+/JsDv81nP2h2l
CneYKGgnaMBV5sgzboRoppkK69sqDZ03iINgOfxQ0qVNyaXjA1D8QvF9vlNQNEK5
o4Am2aKtDfHLlEDm9hx11Y9tDHiW6u3JtEifSJDsN9lTA4RqYccBC8SyjK5mQ7Qd
ArTfyBkx2y88yx3zpTZ7zI5HsysbmpGT2JdjJxhngfjkS86s3IrDuboIGg5Mi3GC
38KXa5ieuTQ4Z1dFT7mJP7Kt9JQh8lGKgux8Oz8SV5AP5G5EGZadsUDrVsGVQsgA
zxyJx8/ZFc8Au8d2FwjSRdTwa2kLgCZ+3mdhjes8HOKI/sIL2Yn4gystZUCskBts
34hdpM4v7kv/x8TE2P+n2KBhPWEN73zYGP8T2/7pR5N2Lm2OF+JEWY5NErIJM4PA
NK8Bqab/1OBspnjQwvHO669yJBXRVDigwHJwVSOYrFySJKv/dRJIzbgpv2oWseiG
toMUJ9Cp4EQheN3yTOp7oan4ibMUFNrwNMQXct/d9C7oBS/xXT3TnjLKhdqBkf2O
qCCA2WSgr40/qa1hxwbnsy6qQ2fcgXjaitxB+ofDZj6baKt4d5Mk3J8JPsvp64bn
zGsxN8IBHliPdp+hYmfpk25T/Ym8dtC4XVc+ghpMNC2ou8SNIfCLqu7ED5ywE9nX
2SYUs+nDqrR7/1W5NajliNSRnhVG02R/Pe0fhd42Z1lVVtXwHj5eFCQDAvCvqm/t
eYYg2pafDy/5WbvZwTSYFyOMG2sSLEN30C079Od58X6n5tLkMxOeLwQfkxmKVQki
ksOP/b1z4Wd/ZWJrs4TsPdnez5t7FKq8yj95pNqIaBakLrYZpmM0kyVpcIRdJmFv
Ke5piVjguVDc8CZE6aQ/aHVLyn3mZesuECtGRLcnihSj1ppKyoPn6FobuCmNk6EK
+bzN52zsK2Ss+oAGvYwA2GBwIylO+74WkH/xUNbqhHukjZLB9kskWZ4qqTa/jcIc
NgumfxvpDRdNNkgt1URMfszzzFIxWoFzGWL/LYvIwksXLhba0DVfqJGZw9ykLFoK
ORraXo2jJgLzdP4PFE+IYJNWzTprZndDSAg+EFNelyIuNG2Wi1l50eQrjWNM3aTR
Btp+XPkXIbY1s8xZWTgDmHUTby37YyUaEPJ3qqEJku8bo5fY8CK0irxcXJmQ659v
ssHm4XNetNe8DJYMMvFfOwNyaECq8GoVCTvrHwVaxjkKD+1UXYo2AugVdO+ll9K3
T5+xZIt1YOC8aCzkCJguWAjY+DnTuQx0T0Mzu2oILEqG4R+m9R8SKQQJxJsXCB5Z
mozlVJhFqAmnk4xeoZy5gXFxKMmh2IKV6pnmpMHOdZih7/WxZoRqw7tAUu1nMXBR
0UvECOLwyQSv8H3dO2UScwqZExVoE2cDljIvZUL9mzT4xNzV32hzdu7IyWUysvnk
sdyoWiMjQAIRB0DhGz/SyQcym9m6WX80xjhPhEx9no9SeELRJcDSNMDOQ8E9/7Y5
FIbG4AQMg5EbaPhb+nUPn8CjY2z4of3p7QO3i4B5voruy1G047VMNCWBH5Q21qyZ
kN404jZX2QhDm+zruVpIeXoicrqeR83U3BeAjVXgeNBCWjnik/AYRQYsZSF+6iMl
k7nb07TyftGrM87kiecW+87Znoq13NifNks4RKZQELt5giux5CC8xwT6nel9lsnS
Ji7EqWIMhxVFbZWRj54DY7G4c91zSty4aTa9NIVQ/sRJClOAk0mHP1kOk61v1cHB
xOfhvODI+Pk5WEeZUB+iR/fyKlR4VD+o1as0yvHl0mu7TOZfnj//E1jpLKVivL8j
mr6hzC1zRTq+fqWCHeqRIO1v16ThaSpmLyDkd/JEjSQ4dlUI44neK9vKy5GSkfvJ
hEJkMJGhYJlH5LlV0vQyFUC9t82zMke53tum2yOQgWLPn5KL/sNKYy/DS0aNFmb4
6BYmMyuQxPvZirYiZP90w1NMnGnQ83DWTLqXuIhkjDIGI51M6bd9rDqZgUPks0xl
mLO4c0P3ANfyhLKaPszaQZlebrqqM9bD7/+Cs2QAlu6fHvFD3IOq1zGfKfXZK3SL
+InroM3v9RKISMPwPSUboTXaiQXK0ht/x3YwkbSwHmVlgsCAHOw+MSXj+MosGQbo
C2OvLiE/lmJTsqfo+8dXXOyBnFeI2+24djQEhQ4F+L7QEBsZRAWtsnhuD73c6B4C
YtrDduboTaH55zW2+Hx/+glB2DrVMVXZiYarsxKvJu9eVhbv/D7/IoewyrRzOHpl
2I6NvlGzR3VOAQGPrqYgaBC7ibCMPTFR0UgizHnaUnpj8sjZiMXxp9O89sotBLsv
QzcnIZQC9wuoi51cdg3P9TxGW0xWq6ISlBkr8PsJm10KSVNm4Wtbo87+wuFN1nXq
kXzxMePckw63Sj0kRG5cEHoYZJX4jnWax92EOLBaWLBQf2whxxrd5chBBNB7WQx+
BflFJPsxZdDo+7pEoT36Mw14f2kgjMtoTCgZ3BhPQCFqZ9ZMuhhGbCzga/mdKgLD
IC7hsLms61Pj18uiPvDubm5e2K7lP80jeVedSINdGJN0s4H5n7ZCw+QyxJWursaQ
iaiiknLxHN/0GZ7rLjJJ7Ol5gP2tFKMhu/xyVXe3IXqWu/t4G+quNiSvO6JIE6Jm
znXpvueCREnU9qX1kjY73LY5Aov86VVxRz8ycArSAB1Rv++ncZi3iG0YeEdogueS
2CZxsC5AgbYfy/C+Z98gaWWF1DNpYDTXXVsLtMHuKBIvLtq2h6vKmwbnHVGO+n64
WltDG+hUX/E51ZNuP1hALkTioL5imdo2U1G4i4wRrSJ9KNbxkyFUh9aeOnfFSkG7
qPn4cWs2awVHysafuKMAc4UQp6oWmSUSn1ipn9B+Xj70eL7pulkA69lYP0dM0iqc
3HtJDGbY71PKwlZNzBAS019oM604ACZTuikOH65LEwUheiRQp+0171FHHMlLst5t
RNWOvKhkZGgEP8wJDQU3TTTNRHqHn1zvE2KD+J/5znSo7uVsYWIK7Ve+LEMeQQ9r
rnHWQhe4AyDWbSFno/q3s9c5QczHarvzeRwuRE5E7ru+3HtgPil+jDz9abd+qjmc
s5Xhp4bWZTWhWYVQiyvewqa86ZyLODr3UXBTwkU/hGtMOyg14imN+zx7nu2Wiyys
5f5BzwuUD0a8GQsTznEafZtc/aknPWd1kvMa7JXTUNisruW99YTw8Qiy7jAkEslL
iCujr+k/zCfYhaDI9UqV66jDoqjTlRG+wa7oi0rn/j9QEHP7+f0h4LY65EuqSbQ0
kqjUZSgADs1q3rI3/xKey5KIJsXKgQrG2fNXaX8u9b/VsMsgbeKSmBZrohgCEpSN
ZHD0zQwqO2LFLumfDLZECIQwGuZR4Iges62IWIByyBWZP0FA9KUcpL2JLWcKO4M1
Sn3KAXPCtDc12HDk7geVQmYX6APsrXlckOZRKDdHH3cez5HpMdELBPWIxt+5tBIM
lyuTTHj7B4Kbh3WCl/nWdZJtQcUnO0Z9mWepRtI/Ps0Wa9p8CFV/mR3Uhf8HFYD6
MXFLH3PEuKa/p/palrspYo5BKN0m7qBRfbDEdRLmZ5SDXCbzuhZxNLZE2GD0YYqo
2Ft01Lm//AldgIW5obl/wbI7jpts76SGU0ugB84XCXXypFnDXaMdcZFUyKDBHQHw
OxQx/BvjGnjXg75i3cSaqJOZsNaxMbyK6GSiWUU/Q8CgXqoY5eeFlREgMQVH6sW5
289MXLwzB2+EKd2p9dUFpgTQDFUNMUDchjnzYtlS2O7p9anGL3PL66ut0oIW5Bro
vLm+sn71kaBbY1d4kD9AbxenLGdRS1l1DuXT5ZoT0bzxTn8COMPVV07SfwlInrO8
ho28GLoJRnRzgj+Q1GZHpjhU2rP28LribVwST2dsPedMSbHAz8GV8TU4NNZy4EJ1
VYj6pgzyvCjRxUXCpbIcvQFFCsNvpiO1VNALQw0JbmRpcsIwyY0JGHpR6pTP2h7U
M9dqfSCHt38KEBXdj/ElwSqslh4JWCKbk9OE5ScneoRmbTwpxU0AuLcenM3BNp65
sPBrSiFZ2OfabdxNyLiOUoa3sy7c3FYUbYbmWhQTEG1F7YmwGFDnQLVw3jJT2nuZ
8oiIXQ4NGhcfBAWkoqcI3VbkdzN82yrTpCbmgmbuilPVaHqp4XSx7+vJia5oiRuf
HxmoWEg8IaRD5B92WUndEC2rWz8tz57N+XZwINrZGiJ3jbBRFCxakaVLmDRl1Yhx
2qVtNTXmxZINduIFE0Rfdl8S8hS7/3kzPMZx8pRkOpNvrjr9zhSySZrLJiN0pZn9
RFR7ECSbHo5u1d3NJ279O0wlQfeRNHUsIXkpE4nJ9bjStcOXTpKYCSUDEdFc8lcY
6kwD4dNWDTOcVojkMRMupsY8760RGRzZWhEkA50FFmCSlqh/IiqykuW2o6HD6ufX
2K4ehahuCMEnrZ2PslumaxMvpiYV3Bz5ijZf5ee81BxoWehCHm6Q8iDPCRDHr/6k
1m7HQE/iO5JT1ykzT4ofOtDLuUZEImlakKRsHmrDALTDX30AXUD4v7kOJ+WUAeAg
mqA+2in7eEM2Z/7j+KqooT63t0sWL34yO1ZcHvJT8Wc4oQOcIbnF//NcjwQkxdMR
UiD9H+qfyoHOAFmWF5hQRoOO1TeBu7WXT4OFaoEfXwaHA+EwE4BVsMh9Fh2y0KQ2
EuJQvmXhHuZm/q5+vD9SEB4ahXB3WdAGMq73QWk4NtsBKWruI7oF3VHhafMrjQ+5
1scp3vweWRroLh6KOpNyPwLRmHcY6zC2FojhN7D+C4z2hNI+wngLhEizNbIS0mB3
fKEd0TMNTMjlN+PZT4nlPpSzCu+jZiTnW2MCOlUqCPicACLVsyHLbknyvL81cNsW
M93rRBT+FCDaG4heynz2JbqWgGVtOhKNCwfcrwok4yDfcvmRuvQGCuU96LuOi2TQ
KtlqEBfI1sCkJd52PKpaBwpGvmF1bEPNb8P8Vi1VxrVv8pbx/uLB4fYxcJfXXItn
7aucJnZP+7mVg+nGiULaqSnya2azGMJnrzQ/af//S3EVQj0Nq79kXbRdg34cEng/
nBCT1qbzluPMt3OnLGK1TtwjAeN7yO5f2Kl24zUOBODIOkqWStyU/2MFXGqBblz1
utMA0fXWZxxMrWmi5Q0fHvs4qAPRZXCfCmf/ftynnaJWVqc2jYRYkffMf7rFOvOI
TFnj0G8YgZXXdvM+GCQA6KWY+uPqUeCC+3Ya6ihzfjFuOlVtOrC8wG/rrjcRVht7
G1shm1YuQ85m2DwZHoJZ/DcRhiIgh4vbJtcLPXQJY3VtwwAkcL6UGBDuZnrvA3Ea
LPciShM6/d0NorGViGG6iHmpb7rdMOCvzWNuX+3Id9tX6SsmHFOhwFJtb9C3YBp+
LU8ITi1MEvM9NJLIGdoqiM9k2LaR9nrFVJ2qzgZKyAi0KX4Td/8AzNGVsWI80JvB
sbvuIFd1nuu9ulFhh112qjz2/ZDAs0G3Pw4M5F9ZSNvucLwCbfoAKTizfAEB/rKW
e4yf93Hd0xKf7Q+p5OYjj0TpQw5antfr7EFLkUVauwMJ0oaynXHemGmulcF5AQOR
x140as/OO0KyPn356jZE6ctigCd4m57T1d7TKO2N8eyqfzZCa3VK+e1E9fTIYRDa
xPhmqfswISjdA1uTzD23HPSncCxBij6J+9lFklEiVS+CRKEdgovLKRTKJyLEY0I/
K717SwYt9wpb8MA1Yk/e60aiq38Ab/zSzsZlrUvVffA2ExP0ZYP0Cx1s6xhn7bdO
zfIWAXuxMYUIwMow7FCWu/SU44TvDorU+DoX8kzqhR/jQl3I20Ohi70Rb6qBr5/x
B5mTIeldO+mkcEqTFYa4KuTlTMaZpleH7A93SVdoLYUNh/4E+PUD+ruAFWEbJE9v
PIioE6QxMWyKrTMB/YiZgDfpIYdgX6LN6HRoua5Ku5KCywKwNBC/QO4ezZZO9ilF
rybQXS5RgxGZiho4I9qMoxXOJzvU8w0qgsbXAOPJJaf5MEb5gp8HXjzF/5b6ZTSC
0iT/PU0DOp/sQ53C/YlwiwVO9KPOmlAhwizrT/v1Wk2uFUMo2bn6mImAVuGeSdEe
00c0ZIZHkhUVlbVqh/S+Ykn6dknMUJAvAJhe51/Hz70/Mi9lXtlAXjnLP8BQQMfY
ZQvLhqSpscG+fzSCKIL8M3HCwc8gBlKGva9asNveXkfB34PxKRm0vOKltJmjhhcj
rjRiWMoSSbKwWEMp0MNnRuBfnXDOvsxMG5wlxHVThh96aLa7R0u6+47AxXHorXi6
pUeezy4P0IE1uUPvQbn+frbIsyTvfRLQQJBSbulyifogbm9oF8rTobEf3rjFVnhA
q7P4ofPrYvvl0U0LPO5uE/YljKYhL70TAHVzil/39T58e66kneVvyYKMTF/yg2M9
52RQ9fMCnftg/ouOCjCNKucP4M3hNr3fB8MHr1tHrbISGVxy2MuGcdaT+2ozJh+Y
dWPCKeshG8bFtvTv+uRrxAPF7DAbtK7sQZMEFf4j9hjejqhQeKE6PHJzmCM9cVXv
kiwvj6Os3J7K1/UpN1oU9z4pt1wDTYqZcIsR7qY+mzRBXWKnaL0ip0F7CeWc0HMr
jGVtAReEuEMCmOcAttude8iv/Ze6rKdlQkNAxlKK4ddKTxwmLmvWxdJKfowTcbSs
XAvX/5VfeI0jPjlWt49R13MNvO1EN54lRVENNdzCpI59VU4WUTHp9oOrhwYSrDCR
A1du7o9/mUpL7q9uwgDiIqO8eBL9xJveRACanfaeGF+ibWydB03bebBhNRYqh7t8
3BtQdtQkh2z8BqcCkoaIojhEPm9y8jkzpythxfiYhniXXlVdAollCQvbWq8HGhxG
7rZBMzIz2dO9S22/xu1GSOAHr99/JOkNLB8EU6ZritSa+6bHZNdjs3XhpKDXiOlH
pwxetf4kCs/GlQ7bSI5xJAtT3nVh9K8F6TZsP0HVNp6g6N5fdn6qFcyE4X7lzWY9
HGnZQAqQcE+tQToOKjZpA/s6CTWgR5avwGCQo2Ke0RA6i735N5i/eCfS78DpZeX8
ysiDyhPYr32wlVPDRc/jX7gFf76FREYXotMC2YMEZzGRRMXnGqds5cXDR7POBAXl
Rwgc2grOIT5B8meoRZq4Dk8RGc0dhU4m5GAh9KupULcAsuiENZlUlVn/jvlYB7Dg
XmcjIqcEzgqSm7mIwT2eUmGXYhpYkmvrHyY5jJYVbFUj/hJofLgv+QM6uZ62jqJl
Sbszi9ZYeZYX56XD4lEaWduK49FJUegR8XXZ3f00WK0yL6AN7dYbCyKehAisDJa4
WUqEUcrFwsvE9z8PucQ2YcrsV4cUO+6JThF/mrrrH7rEW6stZmpe55OYu2KpO32f
7vuDoh+EnPWIRTiggasquydzx8eIemoMwIlLEaY7WrmS6NhmYHbwTbUGcRSXs0kp
MXYwUoXtQmsDH8D4hW2JapG3IBCisY46azlr9sKy8KebCL0JeCX/F22iluoa+gY8
az9hY4wBJhKqhLhOP2LAlxYHX/f5uAGAOQOrJi+hutyLkk1jKzISBHqYuW467awC
ng90Hk6FmOOQRPQa9DQ7RWRpZaT/BX02fnjIPuPiVT5MFNCtZ54pNqC559ExXBFs
xrRaDBarAr32HoVqIV71Sdkn4B18Z54H5INBgv/rfL8qW1ssoYJGi+voTezZFK5i
G/qqfcN0G3D8oa2NEzm/qfaGGH1Cju0vHP9pDsEE7B7xMd3JZfSfpZo6gcmU3aZ/
lpGudmILJzRgET7qahSCxuF9x05UlMV6aoPowt8jrePt84oxsD2HgzonNXLXK2w0
vRK7moi15+14NjKUIlRVhw6OIFk3wjnpdCpJfkIrSULx5lHprq47JbWTvV4A8Z5r
tJQspVsfIzzEKYsMlyKaYVNz9nH1UzWerwsuTJ2crQP26ZLcstB13GBXUR61OB96
WAJnJdK/FBfiB59gx+l2cf0K28ESwg+hsoNuH3EQUdauYkf6NqBGB12cK2pOaif6
Nvksz4/+RH8FbOwzKTJ+qwwfFUQ0gdE6KxKRiCsVxocv3Dyf0rFIeQ2HLka0b/RP
RBa6dCp43Yt5QK+axLnQne8M0A4DbqUxAIC2Hps2A5ovAai4OXsKcZUZv6eil+Ka
gi08C5zFMDFTqlt4JfKuQSHxFqoxPiIUavYCSk5UR6/bjoU7abwmBDNbI28lJfTc
w96zPp0xkvDWZRkFgE0zuIAxNGmjylr5FA8FadtA0jtHmVRCqinSokLQS7Vqnfia
jH8ueB+/7bRkFPjz3dg6WXcUWyrnApWeqom9PYS3Z3rCgUvH+nVPGRfVyGypB75z
yCuguwP7oHGxBGGaNigFJO5QML707iwbG2kSGljhcnwuFcfBi+R2cL6t63gYhpfC
XTbrIPVn7g7AZ6G4RgM0MTkE5yg2M+b0RzSuFzrTGHnGN5ac08MWOHijNKarUG9r
OsUl0El3MJZ9nX8goSy7cNZr1mo3qnExpg1Witl534NPNPgGu6OPHIpg1o3u0jYM
nforS34Zx7T/mZGsC/FI2n2v8fykT4IC9TTGnsHOxto7Oz5ze0S+8AZ96/V8NKN/
GkNRhLXqpkPkjKdi1Zxi+uqaoehQNi9W/AukW49DojpXp5WBrWrjBFWz2vdYti38
HDMEXZwUMYQFeZHbwUr9/lEd3TEjf9pBDkgOWY89hA1Wx7SnUKNz92gMIIR0uwvR
LZYQXKs+Kl/ruSVIKplf9potk4HlpAI3NiS7nq7TfcQUZmh/5Pkx9vWzeM7QwXm/
HRAdwtrQ198kx7C4I+x14+vIm1xQIIvKP7DdGWq1VX4mTl6kKugluudcVY43uWAR
uK8qjVldYeqiH3NnaOIj/Dvjwy1FSaNoWOUKsqgKXKWt85tUHFwPcsEU4x70FA+4
yWGtcC/w1WpjVA5dmjKCE4zSw16J329JdUOR21oVFS/jqNgqJAHFwvQRidTo0/y1
fbe/ApMDYz6xA/8lJGAriwsWAuRU+ibeExBfqTF5fVGFri7P3q1Wpl+olHJFmZ35
4PD1EID0oQKP0awhInrl4CrnDCAM4RlhczI6Z918lWaqAqBYY6LyQYKBHygJpDVZ
4qyNRT6FkCWEzqq8iTlG24iTZ612GL3uhhmZA8G5+QGVTalo1H/T4tVCtsUydRgJ
yf+EpMykE0OL+RnDQA3B8IcYQot6OsB7Nu7mCdahoJzfOF+pInZxuye7A7kELYzN
x1CacKFDJfKDLRMHennNVJuNo6Ubq1bI+imyRY2n5risKmgHA8SNuzMUy4dNsdBQ
PvWWpNfTNYsq+bahGbs9P2aNgyRz0Che7Qi4FKqJj00jooQzJUJUrApN1TME7uOZ
hCU8He88xV7mLCRu3seConMwkQmY+4b46dVcSII2AbvZWSdj9Kryr9EGQlOFMSrM
TXLm1+TeT3xvhmB8AXIbG0LfkAe/iOfjCNwEcVGcrcVNPvBy+Gs1QlhPE7LR6ZWr
C2U8iHhe5xyqfnon6QE90Xz0v62nqnJQsrKthWjjqMaWVW4Ngc985FKMXcp33PMt
TpwpyFg8rFIHY6Mh7BEpkW3VpVc2ux4EHPjIYCDR+67sPRFHF1ApQp+22UGeZywO
9tu1KxKTmNymYyRbdkavidvqrMjpspAVGD5/nx0ebO0v3DYndQZjQGtEYpc9LPow
Rj5ldqiv0FyWjApAReHFWK+/WkuOG9mtONV5bKppCV/hiiCk/GNs6Gk4VU+0zbvW
Nx8yRpBHql1ToTFvdGOXiK0seUr52FE+1t6vQBj4mFr1U5OMwtObW/o6jSoMtrK/
E2xCVF4yEr9V/C0jE0Vfx/tbAdGeutAp7IaQOJVoe8WSXwz8JPU+mCTdAm52QkNj
9E9b05eBOdmQzO7Pam7Kwheom+hOqMeZOPkY0g5eNT0d8MdUGdQZuNRA1RJBrbT3
onqEZ3n9arGIODL/pvyuRzLMvO89GedxRlyuF/9zqR5/P0qOcuxoYpeGiT8qou1M
QimGXUIoPKk6GMntV/p9Y/VIXzr3jJC89ArOacZuX7cdTThAS+Rz1cEN/HHOVuR8
dmjlHvZFxstyjdTfQSVsMVp6bu9zJFicJC2nd2SLy3EwzSXxo+iHPQJ/IQoB1jds
LtrcOmkM0Xr5r/Gnd/y68pMOs62iKWwOdMwx0qGE+BgTBr3zjG5O17rGZ336nAFQ
q6m+6Zk4EwhPZwiaZZCEBmqHrGHcfwxSxr8CKuqLTqjTeDZbOfhwJZLAisRyTeQU
yij7tVxDxgkG3+izqknOBPsUt6eDTd2CSEtjUcYjKNsgXwxzH/Pe0i9kpdjH2DmE
DzeOoHIGxIOFMaqlE7/zC0uBqUPpCC4Hdy8+c34za4qChSB0hnnkeKN+zWJMLlRg
G44ZhyKLhXUN7hWnKkKA54ujvxkIqIX4ETp0MH9BZ4Tmr3qLIOewiCklk3ndHqpu
3JjSu/vndD+C9BPRERyYVAuoptpjXbUE1BNHB/iwSUpiB37v5GyMKSs27/XYgc/4
1V8bRBlj/EEfRxGnWhkVCInrfKiXlxtlyrACcPvekP89UDNO5LZHARq9rtbn4Wa6
YLWqJ7vzMhX3bbjy/b7jcojhhhghCFRLa7h/COPu8iQLny7eKxTFtMuKWlwFWZ+t
I/dKXW9DVG1NkPFERcWRG04R1I3eR5za90Rlk03IId/7zvYFH0m5Hw0LfG1I5Lxc
81WWkEG5TDTEF1RC4BzJsP/ICqeXZZmyjFLmn0XW4W8fWxv9hTLmnwy2iEtfemu1
kUP8i/u9Cwz2hTCHHzTj2EVzQrKWxf6m1jxhxMdwdTd/Wh7ogz3m696M+q72lEio
wxx8h+UKbqjamQnk5gYPGoNmBhc/X24VbpEY/5inmUsOpGAUEO/Z4sOkFntpTzCQ
JenYE2Nk80HTGieY7CHt5QXSCzmY1NmgpAQ22kja005m+A5qoqi55TC+QK78ejrJ
wRwtH+oWmxzF0zOEVaMtbKRz22yh2LSYruiplAPHsgRm6V2TMdhOYJIShVWMQdcl
MspsdTPNNi+pdR5a04fXscjQ/WNH7Q+tx0w2pLf4gjVUG+xsIkTDTLSHX69dkcsN
CR0b0Y0txZD41mjDmuJSsmRAHzaBJbnY6GmkPplXbVjdxsam/kJbPOEUK8eYCFwj
+bk0UNy+DdIomCF+ML2VmepCwekpbGcXlSuolSCMYMUENw0nN8UyzRb7fgJXSaHm
iVMqg9OHjIhSTpCqNiFQA+Vs9XRcEbe0HyObQ9jreVyszKBBT4EctJgj5B0tdvqR
Que+9ublSL6vN5cpaZNy7+gpl1LeDIe3mMl2/0TRzhZLec+qmXptpPuRLld2A62r
Wuz0H/gF6AvesxeiSQhT3tV69mdmavlF6BGx9ZYO02V+YGqJdDL5lJZUbXr5cpf4
+2DpGI1igeAGE5GnLo2bpbIXPcxf0j8Y/xZxJ5z/Wq2qGRyx/vd+4tHKCUrdmSC2
LF2nuwOh89kqcA2f/7xi0Cxs7C4qW4AAI9b/AoBJKYdEFDK7GWmkS4mXZ+gLM+c4
IJIM3L6U+LMX4enZ6lVSrK0eSDcmEb9GppNxEPNuwG+gl4myrfN+EWQYEt7M4N/7
0FYDYH7TIXy4HllKQfljSppcl7s7wPZx8xb6UmJZp6hkMbSQWBer7MaQdVRaHxGJ
hu///wPOG1b2Qpdpb6mbpNklqzipEXEWMsepxlMJSAcu9s7/dEbO2p8vYVJQzHWh
/KzQTIrg3dMfN800eWq0jZXtbTfdvjHj2GdA++QOIHBeGYJmDmgOlqH73xoXdPvX
RSNi1T8cZaEntFNmAaxRR0wcVIxnt/+3DFSksF/yAtZBktratRU0eocHyoig3mg4
h6wfCfuztOHGdNUqWzT+5xCNfkrwxTdG9aCZdSCgMmAJ0CHfcV00xvPkbrWy6x34
oSycADRox6jqdD9n8iZDapNyRxGdMt9D1YBAzKTzS5mNiulTnE9K7e5C8zhkWrhd
dc61PcF0nTpKyS5kNho1/zVcPShOh2sRY96QjHRTXwYzfjcyIswWLDJjw6KxIIjD
x7mtlrI+9r80MEXMZRFVcZLZN2koBx5PuDin4BsZowhQKPmmv/brmeBRSFiRNr0I
0/EMI0Ha42UOZxloPkC+phdV1LrNjB6P7y4lER4GfeGPuliI1K07+SxfbVrjYuVQ
GZJVz8DGvhnbL8iLEcSIOoJ96oHlbyj1HG29uYUJ8O4OHDGzTFKQE10saxQT0KZE
IlvytHjhzBYQXhe0zSrXX12kEy5yH2+DqAiwBnzBu9lmTw5aAKt+RfHaxul3/sFE
Bbnh1pXe0Qu99jpVesYjjr3zfulgKwnroR9yFiqlWy9Lph1MUv1Rvk8PrgWqgDP5
v8lZnkMVo6vsMP1443sDZpkBBTFcJbKsuo0Edd6EWa6GOoVvOey4xxFE4vHaqlOE
bBO2kKw2hvgqrqCsYYrNr1R4wgVfifXK3hmjuStdG8hECGlOc37TNHoTLDIsRQaU
bI9WqXHtqSIAqdnz2V6+13Pe5Qqtnts8ViGxJrdU8Zg/uHfeGEmAWxnl8lUz4XUf
qGV5o5GHRRwZInHOqXaZwQWb0/FP4bbn00uixK4bWE2lbLQCSrRW5p3agPHAdhMF
gnMjZXtxPtc3El4JBaSZmdEdvNa55H7j4QioTDoyXm/5hJ9j3KRtAyjSiRS577uE
4uEX6sEwYKDWx1s1A8kiE2MwhqwSDHkp8GlhKo/J3xDFuC3Os/jGtsFOvKUh7XRe
IfpxjBJeGPSqKNIe+WrzISqF6FuiFw+Sb8dSd+9Q9LlZOLSMfAgMqa8ntqgMWdy2
Hdsc5lMfHnA4kXJw/xtcY2birD3UxGer6bHDgRx6z5H0MEKV++ElwzzKLPOKySyb
6ehWbbA/5QUFqfVeXQOsMPZxjk99zozFxWqI8E/KbG/agAkLTcqkOoos6kLr9H9C
D5joGlKB2NNd5uZG2nQACrZBApra9OI5M10Eo2FXaTu5KlQg9Ds+h1h83+WJ9Z+6
nrKdaq2b32+c8jsdcCo1fjtQpY/7Vsf/y38sGZxdApQB1AaLVxN2EDy7vbVw0iys
9/xIWEFgy1PfOmcVGrHLi/6AUX5ct+jbRriUAeRZRvDk5axXunSe5DGSDC/T1fcu
YHtgRIEDx1vUJbrrG5+aUsKRCk0neztLRW9Q7MYutUNgTmOYnSkZFuKmOT4LUyhb
feLUOFFKISoYwvYAPhs1DHQrZA3TLfkGXMzzorteyWh1n78uRpP6JQELhIuftVJs
FN2j917T34CuvgtYSYLCD6qIia+zpHlVkLRO7B52euN8uyTIGWiddT1P5DcIf+Cp
M/2OErROos2OI51iBsyn7XM9638GPElMHT47y4W4XPtD5GkYVk6BiPi33zv46hnb
JhoPraNBVVS9qrdoXiZEOpn6hUcw7DjA2Qk6SnG8VQIckm4YZNBD6JYeOK9rbMA9
sKslVcHs660kOmSIfUr/WGOT1DiRh0uoMPiZOCdGKh/QcRDpjmEk8SDIm4eLj1WG
MzAHeeEIXZJPBQ6v5RUUGW+kI9cAsUbq7TVWHrYJmG0oBVEaHKKID8RmVFXepHYY
uuYZC/YaReUSU3n0r4Q0N2rAEiKeIEPJU24M6azI4CicE3UK+ZxomTBcB3TlqiB/
8LXx9QsO38+glf/SHye1qbfVaSVetMSU0ZT3TLHWz3PEwO2l9Da0W+LUPhZt2YnW
f+mPWLn08uUYZe/HlXfIDL0KiR/hH5BdYoeAUg/u65ivuqhD7Ivyd5TVBzhctvRe
BeLyXfoYyTrPm50LvLEg66reOd4oOsjcBnILLLplVSl9lh4J9Y6ZE5S/G2TVDvTc
TtXDt9QAEfJiFXEc6xwbr5RRe3Y81eRuDj8ofLiiyxS0fvAtJsbPEAhBfhu6CNLc
gVsjmjU76OqbN1Fdr4OwBHiGyXdaUQSgsQiD1CQeLc+XBIbpeVIEbLJu6/PXOFR2
msMjgFw8UNG70EE+wQX4rFonMvc9WqLjDzGpVvqK9qAEry379y2cx6HVGIzAquuk
iefSlXPqjvz2D9m8txQ0DkWhAd33pt3VxPTchsiPhgGjBRVpXn/V5Y4cfU7156tW
uBXByt67d2eOM1jn8aE1iY1Bg66wHrqi4QBtO2esDIXlA9CSxQf0MmJsOBHJy0QB
lQaoySJW4k6oORjjRCkE3hLTzAUfrTWmISCgq2/Z+AZAfxs7G4q3v0E8+PDC0J6R
+IJVdh9ICxssfjSiw+OeUY1js49WJclnIjHilzSkpdb3igYkYYQN6lTdFxhXXiiq
3YMrA3HIodpFn46Cngj1lMlzBPw5kOhBsxLn4/5n2RFbYB9sdnzOhWSJHYIcYINT
ZhJky/nGxsrkZ5G+A1lpXWf/OyyptVukp6qObKB5APL1AQswqmioqkFE4O/Bdomi
DiMERQnw/qXU/5vT54z9ePhtG/bP1oZ+3BCyggJXHjjaw+2qSW+mpdo3MhFF8IDs
9rjNVT9y2Qztf3C+iohz1cS1xKZJHBZKJ37AC7K3WIfyvxyZY5YXTff2D4Oh/Elf
mEl+zgd3CNL8dBMxKwD+36mu7lz9Dh2a2kw3pTYD5v5MDGTjvQ5Gbe4aS94sqQzi
EhoXu9Y8MlazArT/fuw1WW/8F3eu8v86F5NQdDJz5u2+tcAHRfPMgn4lleFcr4ks
jdSDRAoDhhvki+53lxuu1tr8M1D+fBuReTSmKb1dT/I09cuL7hOJ3fh2RwJ9cQY9
y2/Tb6GYOkMcQA/1+zOedn2XiG0e8aDjWsy/rNZy85j6exu2uk3pDjnFL0uU+0h9
jUhwOyc+oz5ZcXxlR/E2bOhx81WVG6aLqJbcFvOPUkHpaLH2REpi2zr+TEgqXj/f
Yjfsc+eBHL5hYqkKEMrcC4fUmZ8SKLqpFG8eEZWMJE8x7n8jtbWZY3FHRy4DYkgn
PEtdIzVXytxWTu062YN7/crXHQSr3TZCwyyec+xUYKtTqTGi4B1YpIuYBoLc7629
sddchUFqHRDhEIKL5whQ1X54fgVJruBhCAozufYX1vESptVNVm4maHUS6wUVChcX
qs7h9XJKRL7nHzdhWNF7foGzbpBjHmxweyqn1X0ZPVgWIirPTrtjlHqUOe3D/NG6
pFjTR6QPf/hH9s3/OYpSSaqj1eFrlfiH2jwF2XXzBRMsVcepDxs2w5UMWolZn6Wq
153Sl2ijA9OaJqBCf8dUd63A3FfJIov++oiTx/lb0/9eftXEirWb1LIgOvPFnzie
3oqapgh81GaYgaFrBUagaiVEso4gHYth9JcdHjZxX959VNWIKp8HCmLXCx/Tk7z4
3CUckEUYcC2RMUHcfDELgnjYlSCDmBL8ciFbNIFZImap6ninlM2ZvCjjVJIzxNL1
AvY/ZgKaOIXNLixwt0xnTcmviKAFdt6k2Z4DnZaFsrrba19cIoiMiJBwB8QDwwpG
8NUqYAZZQE12iGX9X8qq2iUERElAiMejWFpcdrEy6wHNrPiOkdczKG8reUIkHWI1
lLSYR1p+O20qfxZthmcE8VJaxLa/x2YOJ0ZgMwrCWphmrnLMBLa/B9fLqD0Vy3fW
XwkLBosvqVM6sHTX5WaS9NUf2de36QYLT5gvwf9T6qzPtDbJ0WxpT4la+cupu90m
WgTVuK58Ml2ADTVGeRDzKc4/DeGDCuyQuAR8072lIV2ssP4agyz5dffFRN/BrswJ
ikdgjYwPNSolcDKzD3Rt/Sv1wxbDpR+eG6VRoYpa9/KChJE7IAxUPofXAKLOGjAv
XHN4saP09nJYuZ+BBFKvteFSG35TcHvmpDFqQ8DrCpntBnDWNtTYVb0uLweRV/Ve
O6UVGpXAsXoNRy9jEQqNdR50XBSAZ4cnHvxYW8KII97AuzrE7BPWzoMfRX3s0goA
Zk0WzqegRyfQ7vv0EI2kenqleLDZLl7PbISK9VA6vrLLsEoReRH9DtzIuDehKn8/
hWbH5zYaiFV5aNrgNyo4PcQwtMvlxQ8NxLwcp/lIRLtJVb7Q1urVNGBbThdZ52Q+
9I1n/Gg/R/ojtx1JxW6WHH3FBY57lX8y7dULaX61LIJLtnb7uN47Wy6y0UOIBq98
Ty8K2gomGYbPz6BEVkGqzDfw3t/QB6qQDABFNQy7C5+R9LNH8FLrcuaWSLWc71sy
eEkZUH53QlnIn42sQWcl2+SWya1UDhxxeTwhO/2pnxXiE+dE/rSPYw/TJHIUEc1W
Ysu+7zZEzdx7XZwYFrV/IMhVlqFsKNk5yN6qpMP8JNcHml9PZH2W5ta5kTuwayZC
xOyaTIf8vL+3V9t8CwKcq2r1/TuJoTJu1VJijBy2AUOcIL8rFSY8BQ0PcabPcXvK
geDBBKAuq6hVV5iNvGK8ej2wrKN/0pL9w15bsCVqM/60yi90rVYvp9yB4WzvYqHj
w7kEynWP1bXSwDG00egoYf3q46e3l7dNdXXTIF7VYiqsJfbcX1Tp7wp8EQzO311n
sEQh0hoxUwVs+jC0nt6xDgcNoUIkkD62wndKcBQgoEAC+gPE5s53j+XhAgOCRgmC
CEn0rGdp3fj5wAUAwyVjs5lPrQi+E+sTHHOr2Yaib/et4QTZEEp6GdttLdGifbQk
24Ja8OxTqHF2LcsARTzgVTZsuiLkkSZNm56H79NiGZ8CR0annnW8gJ7+K1rwbUVf
uBTjCFNnIshOv4Jn0bvtIoVMYNHgAox7rE1gMYpT0Woxf5tZ8DEKiLo6KgonVOjU
Sm2WT2C/0CCQfVWNWyv/imwAGKXMaoJcOuUryIw4eFF04JJYCw0AFaRG6hx4b+cd
2zdUN7862u/Lv7DO8oprYn72L0hVs4yJp5rNGjjBiMwf5UamB0kEDiRTHeclHNTX
VN5bHW/Q2NFBPf+wMt3sjR28dPuZJl5ihDC3wbfCxSw2nSYA6W5e+H3wd548HMCl
hkdup9UgZ4+x3MzRpYEL1xISb0WLQQr2yfVP3QEFt0kTwLqaQhPRAq7KwUvSHoVA
uKNnF3MgZSev8Dwc3QhTX3wh9eHm5CpLMLVhbXzdba0ISVrjuA63UgUw4ftGZfdz
TyWaObBQWN4kIXnDE/vD0J8Nl4rFCRknN7lLyRISV0/gR8dJiZ0xfqBbT1650z64
4jUMDhD0Q4rEsN3jMXjused2Yfmzac3PpRZDGK0dyHTrc12V7q0Egy9SmJESvWW/
WfJmFe3Wv+wMuDohq2QigJQAKc5gcrg8zI//TEjvJUQjWN1MYGsyBkEYQJBD80Zu
arImRPA/2FhvTi/MCKr3j/2kFNZbjuT87fQzwq23bhEBznQV47AYye9Y2BzZuJgQ
ys+vc6rd5TjrYSOJ4k6nlDaZ8Rote0MxaSDAx3xwf4S17PDREAGs23aeru23njpA
Is4lxe9Eeri8qEXu7eGgBVRNZPhEMNe/A1cFH7OCeaXtojBPyVyQnXyB4p9TRtrD
KPFFllSnETDakm6AIqG61980SwFzus/bF915OG2STr/v3mdxXBOlhmBUOawp1IhS
lr42QpLC0+kSXPc4urXPalCWpxh8rGtQnZRECF1Fc4OUcfuiX503SZR+LjlFdH1h
KoMFdu5HwhZ1cxn1vXba6HVedA8V7sXKzmc7Z2STrmaU6fsfbelOfWU3TaZqiRbz
atyEGsKnZaUzvvwpYDUh7c1v/drI+oz2pS7yOxR6ppCX/txg5ssHAuZzeslVuf0X
C16izPB7KjQqtpmPqLnbwZjBuifB273J/9cBZspzQDvCa95zpp/sirk1KLEXD+e1
KuW03FT/YZ8R0y7ICK5kgHr5oMex3Z9FZIAaGtq3xVDSi3RXc8JqsiR+U01GyEPu
Gd+h0k/S6j8KwOzJudaLzszOlTSIKls/G/aRFuKMdQ/JW89oidXToocAmT96TiWT
9bz57C3mhLu9OGWJS+tlNQ2M1RyWng74khWBXb1Mlh01F7Z/PuACJD/U5IgAJ8uT
2AK1jKRtbm1y0Jqup8uGlh+DnVdRMeA7COOjqSi5cBoUMLLrmNslIViKS9W7nJ6Q
hfn2AMcjufY5WoNjPP4UW64EVC+2JmB6X+7RWrHNtw626Ohf3kqReVMM10N/BMbQ
WznOhr0bTL4C4EjzvRqbVnJtRHsXPH5na14j4y7cAZliaihl6kfVghDycVtk/Pzo
4oHk7guRL2FuWX6yCkdnf3eQlPPxbI6AUdMp7PIXj2NxXSwmWPQkpdoWFndDnxum
nZDx+oYfptgZTrWcfMkXrr8ViWzMRU6FfdmaYO1J3Z1F+Zs4310pK0YDONw3K/Rw
RltEnCYIfDoi07zN3c1sqy91rnVPwopf0gWK2386Tdw/x+ziMPEadHS4Hr5ILfDf
ucYFMM5uHeNZRXLWnWOgq0Snza+He9TPbYSv6bYXgH9YzvFImQ5HKai5Azrw2UYC
sgnZ1w7WXk7791rec+vVzUGInd6pOcLbkU2YAH3KaxQAhrslE1+bUfKbl2ZQ7odr
Mv4zhl99UaWpNswI6353RSXudwn5N5EnSQAR2O8uHP0YEzSt9Ut24egZ1mFYhCaG
Vl4TJh2XEzufH3lQd3et06w8wVpiEw20ASM5BKNnwx14pEeno2nW2EHPM+3JjHmD
a/gbQnVgus1FMZyx9wx5aNbiHha7rfT99KJ1w3rGSvBsIVjgNiKXjlw7K89wddCe
mnJOySzMpNMaxcfBsgJhVfdA7L+Gl67tufJACQ0Y8binnmb6H0UTVuBoct6nWqW1
3MHnr9G6Zfwn2BdGnLuPsK9FJz11qAgRoYOIRuM41U8kAiY62plf8tQeFv9hXsar
2Lh0HDnc4Puv0wBLxm2VPr3ITDYQa2yyf9YbKTClIeX+S7QdbxRSfLNmui27qDtZ
gSl7k5Rpj6BrwW/l89EcTXy+NChvDCNX4Wi1gLLPiluB9Oj+jeWf1Yfsc7t8VVis
5vm6q1DS8+RnddLLB74O4s7IMNGnnBX4Caiy5qwUYD8c3LTqJ8gl9eAONq133w03
inXG4oo74xzaDNuqz6pNbpWD2hjM/QO9BNhjMGsc4WzX0/ASJ0pSv89nB5qkdw0j
+YCDu7zLY93aZvlOua1Wvm95UwRry8KK1KyMG0cgekn1lJ7IJ8aCyZU3WIKUT2ds
pNZNuE2Se59ZZ5zwH129g9/9pDZRPVoCx8vIZa63hgBShgKG6b6qi2JMS1AQfB4E
jKTZJ7gYPuzXnqSpNMGMmHmQ+ZIDRFJLLfmCGQNegBvLb1g0srytyWq9O+W5zdvu
aVVw46o1BTm4ZXCFRdMTidpjLevUvrMm40fJvXvJfLR6subqZWcFZXWBdu4WG5YF
twAcfAh2SsrBFUAokoTXLAu+V9k48L/MET4UbEB9/ZNDuXS08UK4saE8DDqRGfvS
ZvqGRWJfvAaGLCMeIhPENF9f0wQA45NMUA6ihXE78MGVPbtJOby9ZCrBzeUFa9wu
37T/aEaSTc+/U7l9odY/fEl4ZDB089Z+iyVTspdxn+BpvrtnvA+x840PqIMWvhQ+
8gh7mx8UObkAC0hJRl0ctlARr6ulG2VTjA5yyN4nXTPCZAv6N0uEiU1zRe5YlQ2p
ZXyEJxLsqXPZMxXcSsm23LO5/Yj3bedmCO7i2vex6F6iNHIsE7CarxxAjZntmnfo
mjg6pHsiLE12S0/qpm3+fioy7PnuqNruK+mHCR//4wmiKL7a/PlwdQC4OJfFmBxg
/Cbog9KlNk0nja5CuHkbBabpjDOeKkCjObECoX73VAhN0Ze40hMcv2ZbipItorzM
NRZYv2R86A+syRgliSweglC04+XF2L2GlX5fimZxotGsmhPmvHsS5BnDwcwXiMox
iH2HIH/tRtzsWECnh1ZaSma/wRj/jKEVdpTNaqfJRlwUCouoQdlAhIbbYPttib0W
GMz1vc8MxJji8oiVFSMRUjgTjONbDCZuzFIPlfKnq/uuD1bKU8uhaBjBDqMu/Qrq
cF4aLBEKV28Qk3njoEXMXgV5KgW7su+K3SNcVMcC2gV4X57h2UPwhf2NCG6sf0ru
iOeOnJguEPY1lBhjLz9AcNpQzFWPWcfhqltshtZ9vUPC4ArTLRvTqJYnEYdIwglF
jZuq/QsCgAzBT8KLOaFHAgDEavUjFERjpymZkGE7d/Ccr/ZGbEEDh2TVIislQprt
pcEyjLZSiL+U8mPM+NutzHkPoW+okh7h6AfvL115eL0B0nbuL4oGJJxviS91pm3o
pR/y6lnEfuDFx5ti1D2WQ8S6RSHjWCiPiC9heWMi8xCQz9GgL7GoeeWHiNyElEvB
TLA7E+goEaPbS3Qc+B1izxS7F8dK+IS4BmUVYsvEWqmUp+gd/0Uj83cv09LiGdka
Dp6+d+9n5Dzn60dYXdseTpumzY3xCw4qbeSw7zTSqQxTet7lUBHEEeQjQPI/G2UF
TTlqWCviJjK+zYDsXPHxVDokv+JOR08ljbwcSLerXrz4BEy/SpvUVVtkiPE1+Bko
BqkoeeOyRnNkMz2ho+D5TQbCxLqZfDsXAY2eygMvnDw5Ad+6nE5n6dVqYvVOgZVL
sI4sme2/zw4cN8RcIbTgHVKjviY3IrYl94dC88y+rqIG5vxCO8Vl1M8TTXaMFgp7
iE/Lo6kC/y5bLMVFZibtMYIi9TSUiKM6HGtChvw10kueCio0QlQ0dhug16AGFtUL
eH2Q5LI5gN5EE+5jZL0HoS/5FWKxYEoG3GjV6V8awmF91cgTw1ku2lkfbbqG4NHz
Cx1gomsoOj7PHYjBYN0N1NPabqRJssGxyALWhDB7+ENCUPADW74gagytAvhBsRoG
sTozU5jmnoOAoWP+Zkn0hMP/7apjsYC4o6poH79z1CcxrIa+/cmkhsVqllXq38mh
uhT0bP6JKLzPKB/KGSqnzCci1PgJ293Eb55BaZp2o/EN+B1QWq3AlDOd/MWP+u7K
SQHM0un+Et5H0KZeTVQCBSI6rzrvMihw/6KC3RCf5oZ/oTdWQ4NY5E4VCJ0XfY6f
T6fCjsRyxA2ffXw+V5+36CWZv3pBLXrjDBOTjjBIwCh3H77c73zlfAyZRfF1fY1q
k5461Ltr6LmTB9mA9deKVlgjHqWAwF/YNFpHDZxX1Wyo0MrkY4kX91YHpeOsmP7h
dwpxg4OeWyf41mOXiJGXDHXztcH39dpQgbkIV12Nut7zbJMnCc9M6dSTOZJIBRkR
G+ZvT/oEImK6NgfEcvddjHu4o4VJBRqahRAITLyzqbP5mOKGrmbE1lyvD+yNYp4y
XkcH6FLfKHKviKU+k+H8/KE5Pr25W+14l/MND6yC/MhDBgpvOXiZDyePCGGUSAXz
tw3uRNeM9UVNSsS6+jlvCAcXgaMMqp93LC9lHarhcEfb2QsAMmIWJBwGJ0yc/RHt
8+MScrKhBeB5YxFdzrmucuFObzpcev8U3EYRL+DOp4oSDRiNg7cYSht6dz9cEYgC
S+kV5SptitD41nUVolgzLz/6C/Nt3ulCTI/b90GDbxpv6M3aIyWZq6I+dGKQoY+J
OeiwxncQJZ+dyQeApAbtG+Hm7SR9QNZWcivv4056x7nxuDQ0mIzHJFIOJg13pRTu
w6AYxheZA6TEwrzy/FAgYw1QDtLoWmBGHgRVDMGy9N9Joud/+IGi1iobhba7hBRZ
5RVBqd2HiJ6AzQM08LNZLSO1ggGw5G4VFNNU07+skph3JP1q3hutPE/lD7Px+QAQ
b2BtHHQPVMDK9ohWm6Uu1L5Q6k8802fzhXUtoXgbkHLez795AqytfSqBFpu/Et19
45pQy6TLzaOa9L8xnREIq0fszD9JTGKS9z3Srocfy8KJ+COJr57u9sBJRGoPS3T8
jFp7B1BYvaKtSCJ0Zng08KkVlcZAAsc3FEXTW9Xsdxpidk47E7ETpfjH2EGZiDfk
GkT8z6W1HBkNuNeMrNWBzyyv9RfQA5dGRFR1F0B7RPfVIIjhcQ9TiADJQ3GrPbN8
DvfA09EnX5l+yK6JnGOYdvVhTsyR53NrpoS8GtB9uKQb2rPLquJywnDhOjYkDlLN
KYCLE2+JWanneiDxtoK+/SZvQ4Ncy6qcro/HePDyeSVxvzMJdabG/x6/a0rtN4h2
DHHzOmtPqP9bcvJjvyAWx4f0bgv1vV6yVPVn/+QlW/iXvecJVrEyf7lcFtJXuXcx
oQR+NBofYRbF/cLFoWygqeQEntmZ1wTQOBzzFhnjzLz1i5JY4rbEzYc/FbCdgnrT
w9XcJQkCYYrGj5D7/WqyGgc4tA0jTzZ4FHcpMShO+3r1RFUl8seF9Eeb5bJoDMFA
Fn2jKqToYue/4bF6W6uzXCmGNOefMUK0GBVtbUVcsDxIdnDpTnkswshJuIO49C1R
2/IhTFmJrUpkRcIbCR+Uhu7W+b1VDIbcObmIJ8h4hT0U3U6fEJ9qpOnTQLOEQo1L
TmyDOGs2FYy0HDGelkbG9d7cr+XETrUWeQyz6FSvBarhU2WIp877oDx8EKIe1JQC
0osy2PNgu0STV2RBkVpincGzItITnHE18dTmmtLBeYsfpELmkWKfdv2oIxZy/VBE
+iNBWiMXU8hJzb3CNDW2+42zjrriqnchb6oZB7Ul0EOOylM3sKmGyI4t+ZFoEQx3
5el2/4Tadno+8mxDWd5dxSHVySLWIjNMN0YIVTIaIwWbjT5K7dIqCcGDVEGzj6fZ
Ilc0VUtO3rbJO0wg1RpGgws63mirYRVYcScjpXS/qJVID0DT0ccSFZFQmMbNnYqv
nofW0BxviSltcyrj+McUKm1Zt3nqqQeM3Y305d905iB/5pAH5onKhurp8CL9O+7/
1u3mTywYNxON78fjCZkpxp1vSYVtoUOx7urxMWcUIijplPo1Q85oVfgYnj35BYXc
3zWWK/eaDMqYizuyU58DJChlpkMFD5DkTVXeMoLqfZ/dvO9VS9MvpPeQ6QOFnSlQ
ACXKCa9H2te9EWa4BvzSO/X9Odv9KUC1xieBDe0VxZlIolTU+gYWZZ7k5v1SWQ74
FkH+7xANijym/8oC0sgrSHV3ZfQY2WbGB6kaozMWLbQ1wU0eaXMCPlgUejzNvVuI
1r+E4oLXSCFJBLZtXXcj+efNZaCRth9M5orePegknTWTcFkjtFjeQUYbzl13Z1aq
K1OjFCAjDBPvP0mu/skZ2sVfkjaV68F+Mg/ZC9rzH9HRXUXpnmzfg0q+AJ3YP04I
BST6JMkEJ45m1QI2mqSAptz436k9BuaEf8Ffl99iVR+xUmoyQXdgp3oQHJewEP9G
TmpYcbk84Y8NB4MpRJQJWBNMpW+nHOKbQIeKQ7YvP45wuPmhBnDtO3qLtFPwhuD/
8Zt1tk2JXhlMlazbk4P3VizQaF+fy2MAn+VVYMjEWHptuGc4HpEexs6r63t4wtJr
LnHrB7VozRbIUlMuVq6KG8sssbbRQeDJHlDdZNli6IAJGtmOSKMvgSfLuuVzZ2qm
ndcaraIZSuJwSR+sRtGMlZnixV0gxn3AEi46LEJ88VDcpcUnKYxOkLcZ0yxZuqOz
sB1WQijAtYaCnGkF4ch5DINbfBbbk9g4E9x+W5CVEziffO0ipvCzpp+lMA4Vv00g
Xlc42DKbXgliL3CW+bk4qL3Ojl8vZW0ACX/UTFJfZBdSDt0u5SxV3KBuEiyGAKyY
sj+RXGce2scKaAaWs6KUwMp9oFvbD8AYYFrc23IzZ2B2jcbmvcbpJdyTFNylil5J
FmuDAYAT73oYxdMmbjZ4KrMGeDYgYP5W+mS+mlc+t/sc6eg4yWy60E6UCakpSQm4
DM8OfZjGp/xHa4je0E8XsuVHd1IZnfDImm1RhetEu1BufM82i7iVuPoxcJiLbKua
QLOjHIGwLBYPsmBdaNRr+5LhukXx/d4v8CHG8PT1mbZ3/PJAohw634KysLV9Ymrs
ypUhX2pMXVICqaVjKbtExx3hk9AHzisaVOyrI4TUCQtorQlHBLDjjwFQCsaTsSz/
Sx6ACsRY3mFbgwVJkmnxMKCNFxL/BxBO6UrijlkoyOFZU8hTDKPZ4h2FbsipgqJ/
3W7+yED8TszQqKVdEKQYksvTuX4BhKk2/VnPsGdUIu1Oc70YZOfvA7o36qvRVUs+
QHexWFwZQee6bXC0YAIINr+CdVh3DlF0TkgYZtukk59Hom7IJ8BWJI86zM+Tllfm
YL3FJ4mQCut4n2YMqFg2WEWqmtL12S+OslJ7Q2Lzm9bvUDYRQdWHKzOMq/f+Cbhl
r5IjtZOnfs7JdItdty8wz6at68C6STdgZR7nHlaUsajItvTpP4XParT9RJ12y/tJ
dRkTITLt+/TMsrhtUyNlTX/2cdfeOyvqO0/sMucZ+oc7R2gFgE0eBmi8bpy0sKkA
oZifS4HkGVtcbkuhRHaV8yNMwufPGNGTOAfzjXUeFa6Lms4LUkFXAnUBKNeywM7q
pB6ZmUQizK+u1patev57AMjebqZVRAg+w76AWV2SkkejENFQ4yAR909dyQOBw44z
nHQOkrRvuNjM62LH5tUZO6/VaGxQrgNmfLum5IKVq4IicCmGPAAf4/q2sjNImmh1
pgxZI9dqz0Z7CVOuwbyUMJCSfZuf1pNQBUnFd8Fz/tOYkwx0H4fI1+vnyZ8A5yZ+
epPxzY7eQqQzN5vaiUT7PrHspA3MSEowJHERt/JsQuCZHlN+GOZlXvXuSeguQcyT
rd+T4w7R99krcUBx8do5T6xqpIZwXsZLdG9Z/zAOJ5XBnCpt1LCaC8r9eYoA6gCw
LGUp/DUBQmD80iLTFw3/m2JvX73nDbxIddCfnO1j5pCKrNSx4gYttU8/vnjSO0NK
onubHf6aK4Ij9SNdjhwvGgUGji4DgQ9OCHt3fYZF+p7lnZUq/qd9WaWuxEeZyiM0
tNkypQI6200Gh/U3LTflLIdCjyScXvLK1wklmz/ic4lHYUX2TNk9pi0FOPQf/K+K
4R7kGHDUpS9BlcaAZxAu66/3dOvvkHgq9WFwTR6aKPqf9mKaBmIXJNZ196VPVDzu
r6y6gpAXdpVymlFbCHkgIcgqPAnlsy36ZhrAoqOsDD1839rJ/8zaHwi3LquqKEmk
9OaGbSVDNTm8qKZqVLzuh64Qc4z2iMkCw1tCN8N7ZaILIhPbByEA0aFoQ1s1UZ6x
YKXobY/MhFt4ZPbENpHX58az91EzifkdbGPFhnm0DWuHVZqiln1n6aj29Kmzq9PZ
X+iykwVn0i49AWHsPw7lSr/ti58Gpf1K73AmczFD56JipQf6WVHS1KJNs53AsO/W
ary9A+ajZl7EeqkAqr7tBkxIGL0lCjGYnJeK/3e1zqma5CrBzTzeScKWZ0P3amxc
dw5fF9kRtAGx2qhdpvNcVSIF8bYezBq2Oh1ZgKIWxL3jZeavfbuhiv2F02Ial2SG
veW8SXDksZm+lvBwirZZB42OjZ3P8Q+9RJVbsa4amIrwZcukpY9hMlB6OnTs6YMh
b9e2lnD+JkCERCqQGhpd3KiSQJhvP4IhHSVxURj32SjCbiL2Env3PeB8XFFtTa27
BneeByJKE3qpye/DTAprCgIRlY8qxWnxEMXlYh/IpGZYhFYEQCTK1HRj1ebw+v+w
M/S7ORcI40kRK7Khhk89ECAylgRllTC6XsIGQ5SVMX+0CndEmM8Q4bo6U0HPeuRK
3U+sDuBtAJw5NwnjT2bLYIbAFMHgatxZd/GIu6vaVMo1vye7mMt/atU9TMrcUwni
fFufZb0VvnS7eMj/r46GAprtmc42v4kP3YOU6t21gNntkfo1nhmxgGR3ezEWicv0
JwPxPEYXfv4zMnbfBd7fiz9dNaAUcqixTXKqgFC+mHtWKoIKJoOqHBVMEDxejv3P
D81NKaEb9cEWv9VOBH2iTgwWJxoCQaPBTnUYx6H6FzC+rPeF1ad4OsQkDDd6iSaQ
ovcndmJENFaLOcSP601Zj+mh5c3WDPFFJJ+DJranmYoueeaKnfNbjyqLRhK+sMXL
NmqN2HetPpKBc8DQ4LqmJKwcmv0p/SNBayU3zXDhqBqxb0k02s4th/0t2WaKCfU8
SP1Qp8uQLWCmRmKJMYiBgd3sbuppmcxfeMsv0vxbhN/CTyDaY5nV+26pByu8l8Ng
jfhqeS+yclGzoI9+T7TKHRckd4R+ig5Gt1Uk5lUWCuSesiNWiF25geIX2Rs5HQfT
2ufDuiuOWMbKHgqeLrOY1XRioxPlEstwfJ2AtVfsRy1Wn1GBnPHOWO5iExCu+Slc
hQ17Bqdoh6SAo0ouy38k1azMUxQ5S0X+55iSRo+ZMzKNrM25ZV4PjWl4YWdGz/k+
zbmP8+SMPJnbMz5F8JTqit9cNMgE9DwRrZwaDfV4cGYSZDRMn/aoiOOys1zZPC9+
hvN6N7tIck5WXit3vHsAbJYo8qTpUB7RufwFUgs+RisiWpe16kDIqWCDFwkLQNjf
WGAfs4mn6QIrC+ZrUHJkULASxatZAEmMoLJw0BZd8X5rS6+wzL7zsdI6By1pJIuC
CHdfohO8TWvWWAII2UaixpyEvDNPwi90jS0Bor9FwC3ldkVwYqKDinSbuBwElHfL
NcujnstvamvShUFkpdtmJx36L9hYERbANVy461e22XCZxEk59MzI2KNtH95ZOluR
LFOhSaGCCTL5A0dKEB3gZaOGl/m3bUiSKoC9cNT6Zeh2XGUwL676euiTK4OTzCE9
XNtHaiA4u5Rpp3qzfMEWXmQAOyVENe4WrV0YT9YJD9XRGaiibqi/+T513cA8Hwdo
UlyV0eGXIXUo/v+4TxHKLB+Akmw9IfY0eV5HFagubZh7VBdiAy6qOtwQVrcExpVw
Bk92UGqFlc7FORjXJtUmuqZppnzqLFo22sscrCYDnSWOyAAJv1sBJwhzuqU7nXfv
ILdnnDi4qo+RVxJmJAOMDnFTobgTHXICz2cjW2ClIqiZ9XAq9+1DQt3tjn3XXaWA
6SzV0/pBvqfbmhSv2khJJL+CE2FZEED0CZIflJPtt2317+949foIAIwm4DjHPHNq
DHnkToZYYEbJtekc2Y/h+urz/UXU7JC8HQhwUUG+Mw4QeWQSp68DSzzueCKy/sLP
Bph7AwCHgB9nNirr+5iykWSZa0QjjA3JMs0S7VyVoA09xui9c5ze17HNU/yQv92c
uDrY6vXx4lq77/U1XtFAuuWjLEuifrTWIeYfNEqyWc5hru9pG/nRf+wcp1euG6Ud
EolwXPDyT0d4BzRBjSPO3tZN3PD0/MTTIs+a/Wh+ly2iLd0IDXXlkcpXVJPGLLvG
mcCLeo4DZgs/k0muABGUbBej8nzF/pp/N0mFChcA5ZMq/Hkr77n936wRzsB08Ew8
uOHcCWtOSjz5S4N5qo86JAUZj59dRK8XcnVoobtf8RkxFZ2SAW/CTX8aWZWW1qKR
AfhAZI+ovbfdtzP1ZeUvS/I5nQimGIqrfCGC6X2ycn2V2I53xBgTqnjO2URafj1g
BdVcqMigiWC1YFnRAdWDfvJygGk33WGwXg/uQK0Sm7tKlrHbdxlotTKyptuvYQsw
fm+VzVeOAiHu6zzO5UJ8I6iO5PX4EmZgLFMI3Itzr836HBcU13r4lLaHuJra8IzD
NVlfxMNy3zwqyv4e7iPMLeoIIZHaFvYvdsCKcZbFJIgPJFe6LUCNSGi9l+G/dDh9
jagd8BVB0FlGeKGElce4WP/Gfx5hrtYpYIrMybk3jajalXqSK6vWeD1EQLPCm7of
Nt8jphwFpUwIYsThqJeSaQYh12e0MRnHarwTqYv6yEv5itOGyxy6JcD+TmZJUXTT
RUIby3VKa6NIzP+uXNXLZCC3IRMbuYlU26oB9TqwSrhozXg1UNdJMJQDZo6oZwHc
F4Jdhz7KIx7YybtNBMz4wfcdj3sKQ/alMBJn2IT+Jnr3c7mH/DU61egCEYZYWhrC
99+189QEd1iNMyfkmExroLzje1iesdXAL0AI6uvj9bL06Jm2X2eKhpskLzK168J9
6gsXwbJpnKJItJhHXprvFplS8cw9nS0o7WWcZySXKxWFO+btBU+IsX7K+bGyOTjz
kwlhii/FjEB34a+8dG/8tROWRcXM8hg+2oluCMujvV6/EssLLPEEK8PnnsOMa+Hg
/I/eAbq8K7yQgsc4eT5juwZJp7xxd2eJeBRYtiV8ZoV2Vw4SzIFv8UnlDe6J8gsn
t513MQ+CuhPGt1WZVFrhA4MMO4ov0lgUGKNLJ+aOxkG45lk0HOUWaSKppJtl3Trq
tiIWDqRx5lBk4zKwjZvTninSnqOmM/qilj0rO+zJ8fYOotDj3S7pq60f/EopiE4E
Ukr/3x8XP7GAmdvVstCRHPydiAQKLK9HoWs/IVHxvGT9WfJQYCpBS7HRpnhrACg3
n0Im5M57x73m6dFcxsgy+LMznBcyZ4O5pEmrxyKL3JQHuWHgG6S5+8lq2ktxtUWY
GKXplTSfXpNgfEO53eJEzcryOIjm1h48ktMwzg/ybRuh+aT1HFheB45KWI4A5Tdc
G0mjD9G6+EltX9l3rQ7YjW8QuD3NEdfVXr54eLq1ITE6R/mL9aT+7awT4Js66ZLT
5ZkHCZadYwqB8CrV2LoLbsAwsnrgze5Ifoir+OXH/FQaO0x9veXZYzPLUe6kGsr+
2/xxKmRZuioUDaFykzGVpU3KvVIDbI8f65ynzVlPkWYfCqJpXNk8faR9Dn1/7MEi
IpQ0ZDEBUGwF9zDEF0f9zq5zrUTzJrmRvW9H02J4klnWCmOjUAdkFe2eG9IrC1z2
/apE94FOuKzC9zjbTQ+8lHzQrJxHLNq2L8J3QstBED/kLhPJakUt3PE81ODB11UM
v3pBC3AuYOvc0OHR84mwtHHlBu/6GfjtaU939tipsunwL7CvFHRWfayVYc1+CsQW
LZHBn6B3um4FXa+cZ6wUq8g7hQSQRBvglMqTheE3FkO9kePMaelz9m3VU0tdkHh9
ikN/vbKBfMGHQyPbcOVTYwH9ycMGUs3hiIdbQSOkXucAOojMA+BmIIO4OK1FZDzI
kfAFKy44z5v4OpJZJob9fdJSLN24k10o06csaYXRVltVMLp3PrOG5alincfvUGHU
xK+w1NGnc/eaqzCZLVigtXTUtFtL/o6NZJgVd+QVZZfIq6pPV4mtqhbwrXeloWQ7
oZkv8W03wCqNFu4FTAJ+5DQqPTXEvR4ZcJBa/sMh/7BFMGLoZENC/rHmMzQYviAX
LS7dp8RPu4PXyUyeEbpe06R2GYVEwHhFihKCxQXLOxRgd64BcEmRyYGHQiKoz45G
4XOXubjXhbiuUDAqrfWFTQOMokmDsGOoJO1jew+cFXVHB/GMax+wTlo/Q+gjRMzC
tG0BM2gW8tSRJiHf7SpoTtV4lrWDUpZ4wt6HnqjISeICtFnyPESTg+DdrsqkOeNZ
Qli7+SSQuHIrKgRI211qAWmgnxRfaxVFvpMiE2soP0l9qK/GX74O0RoSDH0BwuRR
SI8wvs/OhC4O+2sj6GVyWv2i0lhWXZg8t647OfEpgc9btNQooZuuahaq6FgpxgU7
Uyy63xpMovC9q4vbOCe5FvHhjrcVvgZvCc/8Ka0mdemxXq6XOGVdAOUJZSAKjeT0
94gCchgfZPvFh/GM/DN5j/UimuZ24yvHXraEM8xQzg1FsR9PkMvngCm4WpsgXRcl
6R5smu17AdKwk5vI21QJ9Nu0lIjkJg770NAhFuajWnFEweQw7ROe7oerPkaQ1LnN
3aFOnpN1QX4rnf/SeiEOwkqkIuOH7WMh+6W1ggrSePO9653VrBkM0wS8HYB/XBev
1BXEuMfXdLlq187lWTtQRpNrsw1xbOfg2SSmacGYSI7jub9JghGW4i1eJLzzqza/
JnqoTGbQP7WN4ip0Ji9AfEZGdooip0Po0l4yavuW27gaXEFvIoaF36G6GlHyBnOi
Uw0TCBRcmpm6wmXBCBedbjplhSHm49IH0YNzXUmsvNvnhRKBJ9Ej4rpr2ElRhH9D
hgbg8Vo9wmwLmYeBnPJt0shw898HLXuVatHnjqVe0XPCUAQ5Pm/wG3q6m8gYxcMs
0BY0g41GZc+PZ4JMUbUbzKv8Q3xoogucBEzTNreaBw5JbVm1/Hk8r2yMFq8Zn9zU
/Y+04p54g9wbTwWTA7MI6ZeNrn33A1F9kDRNRfhP+2/UCqoPLEPb6rG3Jha3UdOI
i+KEr3NmI78NRtoV0kNeCBXtWNmulikNYpypClwdEwVzIsREl7oDQ7rTZlZS00v0
UapaBYumeplG2cT6TtSE/hmHQozR6gyXC5D6bgjqKFHX9Y4oYwY5g7rkuJoNw6Uk
Uepfc7ZngxXpAycwRTZqW9XILcLwL0+fmOZlicbYXdtIsyyhGFu+jLTh0MBPoxSD
aWNpsCfBgwe1CNkg5iCGAvj/1bH2qk02jQVw7VMuwm3IWXuf2tl1vly0SRsvSyI3
9x78iNESurfRB/ZrnWTrg9vVWMQFmM8pbQd/68Cmkn5fagA8lbtKteNeW+GT9HPu
50YUeIxKQx4pamQCysgN7VfTVYUP2yz7xwaIMvIV70ZlAqEbU1gm+bp+USecxmyR
JDA4+aqG7kNGMFUhK5lyByffQWRfgqXtRkurqHGrLkZfej55gxj9F76svhyjizch
PLhWywehqXhl2xYSFT91a+xPv1hhIq6hEhDvp5n9RILaRtvkbVu5iRsGGeGWW9gM
7hTxaLlDh1cj+S4dzz3t9BMEecluQIOsYzOVwe2X6c9GS4OyF3iYlJ6pqdpGoPRW
kklKVFzGf9EuU3YMHLTCrZjUUXQ7vGO/KN90cQ1kiiTdbNpGa8F9gIeY17C5wJA6
c4Bry8JJuV5XtqYOtVUEzAVZeNMxpDLacAbUSpEM/l0KQn6sYDhY87vXDGmYWNfc
1ZeOz8dRAAlcDCL89KAS/VyPaAN5phs6khLmSi9AsY8HJ+SWxigg81PALlFJovo1
mJCwDKy07IUUALL/JAZpjeDzPGU94QxTqFYwhcd/T/sLfa5bgtvGegaz/70bkmRP
peLcejLJAA5ksUYq3HbW1U9QSQ87xdwWYLHgnaUN49luebLHYkwJrSXwbOGWjDOv
382uFdfvluObHJHFQJYVt8JexFHZINOznVuKcpr5PkYRJjqa4ATudEmzMs8N200M
POYaWO1px0x+lW9DI2WZ1NzgEx/tPHE0uOsEZ8NxgoF1/q2+6p3yRtb52da5pRxG
6SI8j36PbhB9z6DGHUjAIX7qwum7mCEKCctfGMmYnlA/P3z6nLQLhQeodxHVMecK
AkDoZcQOlwvSeyskfY40ruxxq5XZKSUySk+ypFTqhJuqnX2yVClppbDJjPHXCDnW
8JmxyEcM5aWrSXcFroBDlN1pm3ns4ThepR8y7Xg4KqB2LaRkQCKGLhCXipuqUnO8
qmP72OXfiDkSMF/+mjK9UJFybor/jGSOUviZLo58kXbgw+Y70r0SRP5171Cz67Z3
ykKD2/VpPUA+JFmu7OfhmLlHOmpobwUz7sl3gJzn215awa44NBCeYXF7blie/cEX
PyYYKHpECVXn1sfoKqgUI9cC2D9MOaDQIdvofr2vL4JGDmYpnRVgHcxc0TZzELvZ
CAz4I7nMraRjwTCbvPECFbMnc333rTT8vZv6EqVCbW6EP2Cy6NXwaSc2b+lcnN4N
QDgwm+sqFY8Yzs8HO1VvcvXX/PuFIzuoVV9+yPOXMar6rFaxPIBcnofaokMGmohk
+ZW8rEqd4HlZxT6AcHg2QI6UzGl20bEbCNaocmfZu89v7p6q+NHKSDqtIaXiBhZX
e0VrnEsuWE3a85oYzyOTFKJdiKldfjxqeW6jtMP6c5R74+gZfTQCpBQ/kP5EMcu4
VTriS9VSOnK/s0CTxzzDhEZhfIzMZyuL8hbAY/OI3NZcvNinxSUDGUMjLudTsEpr
j+92IZX2IqBg8xw4z++VgOnF+77nfHuZ6WdzgIQELOLQFmP+Qquf4dHJZMgjRzdF
wlxClPWgEdVdBERUi/t1A2Ix6a+iB9ppZlELuZd/7yN+0cqnZFExqpRcKiZw+cbk
b9Wr+GgBsb7+nEDlJYUGIOb3si1A9JJ6zlns7JGqablo+NMYjsFMkr7ub/IvqKbi
oObjuEsAa+P0837G+cJYLhtOOF4LDP6WIRhlGc+4o9FdjRn1O4y5/zLCBZzM1KRY
FL2D/39KzWnYjmK/ZJtk24vb2XOuDpWFRWu9YvLLYHxcVXHMdBbdakggH2L3mIiE
ChfEfOo0+yNKKsqxIVUC/tNctWa4XwYTD6Xc+snBT+R0bVM6cMGvD5W7sZlmxgv4
9w+hTjwDTV3qQrYlDvu706PIXpwIQXNkz+WBnv0degSgxt2LHymVhsfHMVHlAPM1
q29tjpyxmQDMbzHSc0nih45ewwinj8BS7Or1f6qyuvwWNZSBseYMyr8zr1UJPMMB
IXxtLmStThrggaGB8+yBSQkDK4WGDj38pOyFU2xc5bBnr6Rc924lnBoadNLGKf7n
0BtsbHW3u561H1Fqxa+0z8Yq3OMhX9a+j2vUbiDVEZo83kWbO5A1BpkqqXXWWKhp
aqXqbmbTWjtyicwi/P1zux5SV9Qf3sBwnFfbLYOwTYg2fjuoRDP5sd+LYMF1+OpV
nUwukq98jNGlw6JmpfDjD/qbs4iJw5B+LmvMdJh1tLynuw/6SSMuLhL4+93Puj6v
8hFh60NN0pCbAGaBhpcR7yVscHEXFnqvnIla8oPkMiJNS+3i6BhpuFlAHZY1hC8U
nFEl4MfeZyT0ld35NL0J3JkH3LXGAsPzZT1E80NktXL/IyDsjJpnYudywniqDZ14
Wasc5Dvf8jR3w30njkJW73WzRKIKUCJ36m0M92dvuAZtdAZLbrHAzZG1OiWEkXyy
Sp4GxOQ3aaRIrBhtA7sCShCQVmEgXZVEVBYyD/LI6j2WQXUhowuTK0/zllBAuvj5
D8KTFqVk7KW1b1eLItcAGhQIa2mVUYFwyxbyAXK4KwV17bKDcFvNgq4ZXSVvhO1F
jcVAVLYi9QJlnp/2hhdeiJwPXoiYesaLE1S8F6TAVIWt5V+DraouARO+aFks7MPF
xYI3ZKsi95L7AwIv1MEBpiJXaYmvV4DWcgPB3e8Z7Utd5TJbK7ii2FDDW2OswbGc
S8e2cxDw+wKop9tyyqNYBrEw/fpxMkEpWAqr8q2LNXWwJto08JVcKDuQAQUssAt/
SLqQQdV7hYOXBgAgNd0u3cuv7rRN4oKLhgtmJh1GES3cn3XHh2JBWZ+5KOLnHlor
V5mGFAySONoYtdN+yPE4v/6i5NvtiqZyR9GK5dVYkVTSRhKHHUgLRpOwoSAAV5SZ
b3r2lVwgv4cchaXilc+btq3Jy1+YuBJZwu6fhqdawXCiySxK5zyVUSOtiChSeePm
ecCP1ZKyxiHdWUq6En6PAurGk/D8meov4pQGawlIGea+1qc9kjla4CH90PybdWYO
GQ0lFav862yi5CiwwbxFp3+SuYHr0bOjYheKJh4Qxt7vKeW3WYDOK/05Y2Ndi1LJ
1Z2QV6NNhCmAe+tV6kPUmHjPjDl7JQG9PpgLMThrstfZCp9AAAN/4/j6KCjBCbmr
2xbVW1jSbWLGK7fg1rpGxDVdsDvIBldVD3/7Tk97O740LKigXXdScCoaYMocZfBJ
5Ob0i2ZiK11nVdNb7fsr7YZ8P1r72hX39viMWiSEUxtU1WCYt6l30xgFkY2XAdY3
66BhZN92dlrdvhojCLulatazn5cPNksRuc5wiibo9E/+4r1Jyz7inIE3MujorpqL
DYsRK5s9WHu9xaQFiDz2YA2sILeHpZsoG5q4AeRW0FKCCJwHubE/EJ9Y40hbtiqJ
luC6vbzhpc9CdDGpMJ8HMOMq4dEt0D9g77gqlnNdJjbWbfv/adUtS9RLS44RpoBc
gp+kq2P23LTpet2WrYw0ECqfWCdDHpHfGsknkWFq25t+Qpo77Mocxk2SOEvkT80U
15QdSKiCxnGMRRO5gehV2TAF4XI9zF29HqrVZYyYlrXxzdUN18iqGOf292y+t3CY
m2qOapGaK+Ow3RGs4FAd9kUBfgReVTEKWVPkpkyHn5kqH7Ri1FqlTYdgiJqMie3A
ZIs9ChuuF7bnzTlgEma1SW6fCAxJwInrN1nybqzUU1X9NedWTNFIL6J1bhJtsCKT
R/P5VQRPbP3ea3gErfUBkVZA2leKATKROxt4gJ8jGzUctcNfmYv1f8p7yULUPp1V
nyWJ/CtzetL9NGVuX9Zy2jz7ZREg9fD/SPRqQRNML6K7582tQ+Vgd+IDG/4tApof
QdQ4IBGVA99qUMp2LJRNlaUsxN9jy7we//sEwkoLIUbzVn3W+zMrp7RrgYjTw5x2
vXmG5zliZmpmSWNUdrPdU51TPXmRQTxdTW1MqexMW2QaD24XVSBJd5m9vvcDVTCh
rWw7Jo2ANA13rRL5aQ6+enUQjC4L0GNkarigVx7BMDYnR/Ybxu5SFVRd1eWmBiFm
jNnaVebcQkwNG2SBOlUY0C2YqdFEbYKb1ryxRshvEORaB12hyv6eZ9ccMPizueps
jBlm3VBj1sxfDZ9IE+0aUYSQybSsyspdggS8H2h5DemO4e7tTDAZmQ66UuksSsV6
8YyYxixqzj0EKPuEfcVSlfxfcUU+6WwvnNdW9uYSouEpjn96E9UF4NTEeKnw/YHL
l/l6WKCwjcEnPoi+OiOvkggSvpEMb3oNkDUa+zPWYqshWx1UBgakngxzJqB70gaw
X1c/hRAB5a/IyHafyn5tcgGI2Jk05/EAuMWBpxuZjsGg8wOc+4S7vq+LfAcF9IxM
UZSyTcKf/DkXBJoTEM+yf0cLP2Lceb9kwUwYHLeHIQwklFi4s3G+JuXVwi593nPX
gKLpVEgCqwbOukkF22x8Y2Ln5nwrK+19e4kbl/xJGm3VFUon6EVjXqhv8x5RJfBS
alOMgI1zp7MfKCBxnR8joC9sNxE16ifl+fBAkQ/VkpC9MRBsbeZnNshf4h/MLJ7v
u4//NzKzpbzy8nCq5B5TgPh1V0FYQyAsHAuLSkQIrpMCe/mMSQyz+zU3mSfv6eRQ
3fQBY2dGZaRyia3+baycGslKoChjOYQ3s0rEhelGqPI1G7Rshmo0l4CSi9VWJD3r
UfkrgfgQozEvJenuF4A3ur0raf0iYhwa3kVKh69OXRbfp16TALrwa9kZrqe5WhpQ
rPplCRHi53dw/ARMi1RUZDFjvLYuusSsfOUmTz5js+0k35tF27mn9xupJtBav7Xo
IcykfquWJqla/NpAgPVdTHEt1KJDZGypdBCDdVB+zU8IdHOwW1pfMyH2r1jzVCi0
t3rrfP+8TUKSNQKTIBMjZAGpHcTDa/cdDbmUuEig7AaknbeYlFvUC0u1oet3e7mc
WdeEFnx+XPsDJ5VaqwTgFyUbKhmCxlM93C7hERtbRYr+rJS13FX2MGgLaitL5Zli
WZR9pAuTeuZ45Sw6BCsNB9UuVEdaBAvJuq2vyV41TtB1EMFynqi1Q6zdt09OgiNc
3tNV/JxLxiW8HYOALlhQpOo+AJZi144hYeehX74SjwIvrGyfZoLFBdZNWOIs7jLw
Badkrjj4VevlX6dIglh8TSODKgmkBdfu0sbfx/es9S4G1efxp8BiHxo7i3XqWHTc
ZGylwi9KdnfLjAx3tqIEX5f+sy8AGmCxMK8WSbeYgVS/zo60+3Lrlj03HGaqW4KC
WTX1Fzgwa9XuUP13zC50wiDP8l3eG0VosWGnveRJ94JrGADM8Y619iJU8RHqhpJv
G/QevKb8rUsX18LgLBxoOvman3wm+XRpunxWAimn3GyVAuHlFGLXW7aaueOYpRht
yXgrlnMwbI3EXjkP4PFYbUbR/wc3kcPuwg+1p7GDIDozEWQ9jaHY40KzFuyMeLrL
CzwP9Qc9vyUKMSNttN+TcqYnLudiMV5dIiAZuQ9ZopkB481lQ7T0E+I23/KNePau
BNwP7R/3CV/t4L/WXhH2ipWBtTzlypY0ogzqbspIIwcW78i0AaetlJt9DlUMu+vC
eS9leDevYVFcaB+t9+eLOUFEyjA9JJXd6ZyLVZG/RXHCEcW6MLHv46BWEzMcXCA0
nwL0dVq5ToRwUI8tHbwsf8FBU3UfFLfeZdeFajLuwcwb6q8PSCwBx0C533R621qZ
V7XRYrFtQXqJmUy36arWq6RjVvTxkVZZ6udWUoVEjnj+J8JqfA8MKzTaUtmuGVfH
O88Zb6cIQG9iFlGmOQRjJ0lwBNvf5EqaSuG/ehRhZblWQwCP3mBdvu1AdnXDKK8a
SRJA2rfPy3ifsbF7FItuI5UjNfgWMlN/qDeg/wMDJ7AorIc4TGZiEbTg/j7zjV4H
J6kAaM2WPso0QmlSLDcB298mTjcDdSFBzSphu7eEiztOyTTdG+CiJus55Xo1DrDa
XV1FtM1pf1gs2LZOy9+iIDGTMCy2xhkj4yb6P74Z0iYtRI9ChPlDsM779iryeK/w
0t7Y/DQOPVpclU4g/YZnfZzfSbafy8XrHaI7uLA1gk62N0kzr46Xkok7UztJd2Po
RVXasIqrLmzHKPDqMAVSj/BPQgH8G0FshTG6UCpKlbTfgISsqJuWBdua+bm7lxF+
QBgd8Zn7zxJ2Llk0EwDmuW4pIwxeYWjiq7k//8fd2wul4FRfcdHhCfbTNra+sy5o
3udTs3QVWn9QOM344plDoTbVWF4F+A1pfSTcgLlbagcKpb1DI5BaomnRnDgsjGbI
3Rd7fmVvNHESL/CCMtc30dpkxyJEd79Gn+brF3e5r20VCp3Y4NG6Dxcgd92QB0fF
yKumn3yQpOWUjKfcB20uA35hoD6Qz1ekQj5rEh+702Ism72ZgL8SBkJHcrctwf9e
4t6ysonDChE52tLN9HN2wd/sO8xmEePMp2R5OiD55sstJDFm+aPHkMYARacSfTPJ
rwSqoHdCv73gH9k3N9LzkEzu/x8EhCva9kd0XiHU0ci0Yay2oPKVlQSk0g/pJ/Dq
kk1ZP4BK1pAE20iJdAPj7QbnA/jp/9Hs8UK9/nuyDfzWxwVwvYMOheFPEd05+nuI
QCdpescYIxajv8efYUTK8j0DfN05YD8gU3sjil9UyJ/n9zd5p+tw5/eCgCeCGgQk
sY2ARewydhTEbUX259BuDTYsJZRQz1kKzB+dvUbTXpCJuj7Cy3buG3o/nvQAxJAs
xW8cO7ubG8kGGL0vrYo6fAdv74HBma+wnR3xYh0iC40vmRatLmFPC0uv/9JcldpR
a1f1eb44xlEFhY4hhUh6EpjYgL15SvEV7XzrIRpsiov+HNpwJ4+C9JwPtLV6XTe8
GevsMAME0G87UDnVxroG53V/IYP4X528ApEJOZqEDY1/nBfYtRr7HPz7sl3zQ0Lu
sWGzXtAeLnEnRJ3hlx3YCrXD5ykk2EAubMBzBlYg17vhA/7gtOcKTXRONXAZvUPA
tlmZbW7KsMNG/sxFa2srzvdIXxVFbRvIc9+ed5fAib7pANnvZRgUL+2xU2/Tb1RR
ZO7CZk38xphlAafSx2w4L5Wy1Zlj+F7+yeQnxSGDEgoPz4NDUXU45a8ACiwyHtFt
G8CeaYVQIQRvazCPf4bST6yzBYR+mZ/7lPWeHyZYgFstupLVerX57ufDCmOxMBBv
vTeHpPdRJs9FLkcTiQ1Zwy9OdVdKs2XNeXgWJiFTbGZeiSf8FXLwZzc4PJXzsDqG
rzPXno1GYb00BRW4RvAuB0cYjCOzfpl0f6WnQMvfKhGmKu1pBGJVaiMSKErP7jgP
kZ16NLvMGNcfVfXBMjCd3XZA6JPCEmMR8hBAepqMSDXMRSFccWw9RzMcO4qykd5l
EMB34WPmROVpACIRLPz/WuzX6T8DEAFLF3SCZ+lS3Ag9nqiSkP0tZ81PVT/mQp7g
jWoyYkQlDAkOO12VhygD2lUgsMf3ew23Rkjgy7ZG98YBEaLc3DCKbubxjVrf98t9
E4T4vBQb3XXKPsCln49SJDttVUlqmie66ffmDqI4hFw4q/JOPYBnwB1iE1ZjnTR3
vKJZ77a88LqNDWY9suIJynwP7pbl9Je0+c/GUGq2eF++/yASXDdcDl1+HPo/JX06
CLR4WaOVSGmMqVIdSEeu33Jvt46Dr9Obu8m/isrW8Pp+2nwZhVrW0HYNc5+VSjmi
YbGFK+Jty8qpsN6Oq5RO9gDfYhGqs5xd1hU82HWOOcQSKktMuGwi8Psa3IKkC5g7
PV+TsLuuE3/fh3TiRDVh6686uzbTIUAI54ihGmUANTOJaYqFPZitLz5zS2yelMTj
vOCWiZtlRciZqHSLfEbk5UWF0j16z7z+MAAfhATBGfZGhk6UAt0XXg7oBZSwceVI
NKjUFLfcLAtEo879Z3fSTzbvuVrQo9RGB4WRyvwaG8k64G+g5+rlOlPSmAjmoFiR
mWgRjT0muGQYh1iAtPZfmTj5Xj26I9WDAuWC/mLXYFSEzSBPQWrYNNXGHmXVVCMx
tkzRzA8EtEEM117EtE4Hyg9hLKE2itU7roBHkYMZT2WIK8UPnKK93m2G3j0xvnLn
cxUsD0SxDNGaH8zc+Shiyy9BhKXN/uvk2xdi3Y36odHLaKjotII6fBcAKUU9gFLy
1HCIAeVMxIuP/RMyKhpnay96YRMUIaDXjEPUhTrGkOKwf3uoMGBdu8vx6qt+qszu
ncracHo4RABmhXx6inGkSo48FWhDtG+3YReXgJBMSIx0G+Ggmg0msvnCK+zJkFiD
iQ1fL51hR7D0tY/OrKGprJx2vDbWq/zavaHm9DQgbAYoJRyQqsGBYo0Lw90co4Rx
faFqhniQzRaio42bjTK1KS2b4WAaaJv3DGw3RHXAwGs1i3R4/hW1adlnw2thTtg7
SzA3wSKHd2uXSRD8Hgqt5j8ES3arrXCsELpNN2HG80j+ooZC8pHIscJNTmIYUMrS
IGC5rnFXwZnnxsIpSDXyLxDO0ru8p2tGtL+FMcjVVipjn7s38DqshT4KT0lY+pv1
5/JyIqbLhKWomv0LD6ki3w8oy9qRYRca2i2sHkG6CiEAfamiqZhqx4xpxLXrZ2Rr
HpWk+eO6MEk2CnSMAVFU0mrJ7g/FA9v1OTnr+HSjekMOTx7/hlDzkWqq3GhvfNZQ
OZqC7MF5m8+GZT1Se5TOPT0klvFrFJk4l3Bg/Dhh5k+N0q9J1JG03pZjgZnI1GeV
Sz07hpl2G7DI15rj29L2i8EGFicYtDX4BUMw5YEoAPW4TkaN6tunNZOlBh+VvkUi
CR+1cpXvKeumZH4kaRH5Uslw3IqhbEqiXpgWE5Y+5E2NHvSgJB6lfK+aios3lkEx
c19qm4dijd0JFK2W+8UYAx4KaR7QBdJVI98bv3lhDUqyzCKEK7tmGShTfq3x7+3h
bqADmoRN5J9c2/t7Mq/kP2qydTershZz/HK35tslgfMr3wZ5/2Bj7NlpL3G3yL9i
laaHLB6iTyYpQ0tPyJIKGAA1JAb4s0nIxptbKqY4OArDvjrua3QfXJqf5XfQ1Wt0
gpSljhMeenRvf+tt0EEm6ClUjAyseuLKku++EipZAeBlzuNtrf3qKcwQbvstfC9J
+a3JW0pBCjKdB5SG86Mfo25qKy2VrOmlt0k8H2nbxjuTiy6Kge207h/pXkF2XQhI
kdppVj6wCaXUn+FEnZ2gSwmiwqBR6p/SkV4sE93eGjS1BsymRikjfDPabozKMoQ+
Ftgr3T86i/vd/T4EBbM+I1zzLAipvTpdK/gKkA49kXWrTiYw+H2QYr3LxQb1UCkN
8DbXPGOYwjgJCcpyn4sD2AMM5ab5wkDExaVkZU7D/M0YLpWz6As1fx2FKPa+Pi44
Qa+/M0V3ywD0L8JyxHuI+bAyB53FAr/hVMv3L/QjN1qrZkt72jAoapCYpBBeKFLv
qxKMAuV8sYIha0mVUUUvKmeq2r925F2GtFkBCTgNd5cB07mq237EjxJyG8POkzO9
hchk0K3i1h56D9QJ5KzJQwLIIXFEQ8yR5bHB2TgxI8cj4FMSc5tPyZ2C9MzcfG6M
KhtPvUhBXnLQJrXsgJMvXmJ8ACsNC3QCCQY8oQNU+Mj/I0wzM1vCsxSnm5iLgdmX
iHnFiYImraz0noX1yAlt7fK9iDBc8w6flshdSYwRASwelWG9782reDVzTDsWsPv1
zcOA8gQa1KfuLJa/+UjV1Vwh6/zFEbeoVLA4BzsCJM10PLYJMvkOFkvlVV2yBRT1
PoYTrHOUDchTIVOfFLstpH3CqU8zhQrTDdtgTf5uhWHZKmmU9VtmhJuQtKUuH64e
Cybe40/djLHNhnmM3lQpsiZZdZwnB6Iy4W81URvHxTXeLKRq9Ktp3qs2O5a3N6/N
YD2PvMwfbS9CDjAjGfatvguueUDfEizKHAMqe+BcMzTlSR/pbObMj1cweBtmcJVI
GN763zUSJcUormBxICGExxb14gClNds4hQopS1K1ftpq4Z3uvnBZlWbGwpF4wSG6
K6YB87i6roMrUXiP2tuRhDK3Y72B45qesuHfrf5ZoI3j6SyCKuVdVBGKJ8ZCL4Qk
8VBEc7phHmN4IXsgQJM/dFzJIW0dxHKkbXkivddYtSMpRzmTSy5WxNlCCLDUJmnO
UmUA++hrzbQ1R5kv+Vcy1Ma29WI2nSpfOKyONynqu7zFiiIkEeC+iJ0pv447LrNP
goZwdgO6yKQIpfbkz+m61DWskixq2CKEJtJ79SFBqhn0emGBrQInoqWzMBv1ypo3
F7TvyTJblFpFZ4y9vcHw9zYctYWmheqvUgwaSVWR3HA83c3MtpbzXe0SwIKl19wi
u0eFpfifgCPM5NNH5ntKzRn2bxraz2VzAFLyJM65Y/YwjdqNs7L3wJeqFWy802mV
o+Ekh06kWaNDquPom8mHtvYRlo8RfO5oEEUFfa07aijWfuTcsnZe68BywsXAlsQH
ubVw+ID+Kix0IPPGqVzn8xJHwCSebaPZVyz5SeoQsd0ohexmH9D8sxTfDGEoPYU+
IbsTR1WMPw28YkWtvdQvyNgXFseOFCHkJRcP1gJCa/MTm/mLpXssNEUjuWo7ap9Y
BkwX67ptw+gyOJiKiiAy0WfGMrNlU3GobBMOUlDpO3S7Ec6gt9GEAvSdtMcRU1hp
0MUb3r0owHbY3GwBmqq2FZy3xFCSQMWowQ5QwasD0mEWF/ed4srWwee0CydSlUro
zGWny4loFXbhTn9dWID9tyjpq9CSMhJsfjEJnDmArEGFUA7nbcHvvAsRLAKLx3TW
iKJ47LWJS2gBrgKR+1CdPBpbzKxtqjeVqP5w0MVl6XRnisGo2ObA4gQdlzhXSo7m
gMyFSO8F+VyPJ2A3ZMn4bxlyRnPiJSkpxL1wwkSPbRwVawUHoKaxuk7/sdl6iTjy
E9fA6YAlFIe2fRVtaRpOUvuJPXok7PbJfcDgBwDLO8CIF/nmUADihEd0CeJVNjv3
MPUyw2c35i1EvEO0QApRd/9fMotFeN4oBKYCZ2J7PsUMAOczMZoQRTHgiDLMNIlX
3t+35oICDBN7rGKDCcfM58hXL95yH28lMzrOUYyDMwYGLHsmcoOQF6qkTr1in1M0
Plhh5YiQXEkWgLDzS7FW7Nft+7GrHYO3Vj9PIjFQjRGJ9oIh6UgjzzmrFSHhrlly
t1Gm3KjMrz+UzUUwSBPSbH3TKyNmwYgO3CJ9Y2/eZ7hh1E5V9tyvMNwmuhm+Px02
itVWE8N0AkHlStIdXo8XHLCdHA13L15bFwCydVs7qQN9PCzr/Z2D0xtWuEuWRRue
VkthDp+kE+BOMxzbmxN0aoWj+I+s+I2fueL2FKC8/M4Zds9SYykxRGd00alGlnyu
4ubCwMC+XDQOdp/LfTDfdo6vcX6pXmqJ7vJ6wxNincgPthtrgFnnh2kgdbN+T3Ps
hB+UI757o5PhIsnD6sCEmkbcjICkiuK/kp2aLIWyak08KkdZEbb6KoAX9zaHnUYQ
JrK7HSniFwv/183mHHPHKB+c28zgwURlXfy5ujF4F4i4HRGeJn3lGHFr3KuEw57b
VlXxWSA1OjO3dOY4EX+iIPjqyEPaovDaT0VHzTSkm4yTYz20cnIODLLBXnGxkpbN
OdE0t7k/QKZ5WcZVAOBS2zwrMeZhLRkn78rDmYKTV19ZHppNd7yeoUWwgaE4Pv2J
iB6a5DY1KHjTPN77pLEZpePmVg5YMU7jiWThoM0HVL8uNum53uLhn9rbnqAGI+EE
S+fZw9FTzmcxcNM465mW6XV3pROwD4+ahHTdUQWTW8QZw9Z6VmxxZsXBtqdo/TOl
iC8t/J8KF71lYNwzeFPGcjprAX7zhTETd0PeczzKjOXExHnE0e00vDWdRTbvGY7o
2wGiwUcXrn8VU7ZWTDzD39QKmrDqdJDtoIv3IvkUf4Gv9rSiTvCX7Ut0AoqbXlb/
8tRfTH+cm/eR113XzcZpgRrRqjsOdHHBU/jZfmC3RtnOkRj32q8JjeaKxHUq+tF1
yo4SWhGlnHYm3IvNGM3Qdp7LTMNJcDGPOrv2B19r5qqoZDIT9WGSKJ0XvtaRHWc3
o5oVnksT5xFOveMFXkZMSIO1aBOCLRyDTdMhKCPbNRynSR3I0dAVOd3MCAeUr2Ho
WUA7MFEPoQcL3KCm9OwvBXfxmJeJGk1z6JMrUPgBNHcfW/tFQQO6UMFRuC8bBuyi
ynBkde2QUgOT1iuVOJ4PxFv+Gkqd6VQjTkoqw4rr5i7F8NXnm5NCRbhkZCSXb6XV
/YMLtsGFj3dqaa79DxbubgUBer0mpnn9BEAG6zMD0ypkcghhp0oxDnkiGzMDaRzq
exUZ6jvXkHG+x9aTf9DThuu8DEOb3r5p2H+INvHdhkdUfBx7Mbcs6GBEb6f4spFV
1OXg2ToiKHyg0zRacxZ1ssVcljsvbxLvXIoNPkHJCP1DcG4gVKPI0NV4QDyWg+eN
ib9b37bxGqjQOz16f/q95rMZyOI6TYwyAFHWqmNNQlT0SBlsCWsn+fzbAQXqVwt+
ZHqHfWOpDTf/j8ynh+GSSwWDUp/rrThIRw7Is8O++d7Aj8n0NK+H6KzJDcS5AVbu
CznSYxZ88fXzqnJgaPPeXxnV+KPcdlHrS+HXMN+UsTn4cWR0lIl1eSg66GjoAGCZ
2aqDAF4EBdYqrP1UKexqK2xQ5wSQJLUFqXd7e8jluoVMp6do0g9ncgnonkO0XHGU
ZsTnSQoQ8SDF6Z6xfjWjukQowyvH4exFBS/K5wYyR7p+IkH75+pCSgwE6ENUnMfD
2CzcctXPKgtcTVanoi7g5V76Q0tNbP6Yxrm4AnoeLrSGdQcMuHoi020eB4MurLyi
bD9XnnI5ZBNGTMyOpMBFApLZ/NqTeivBb9zvFgLUjaDsWQ76AwMZEWDFovSGI8dT
4WXvaLgLPlsgppLZjD9vYd4sEHcCFUKjsV6udHbO3LlELfEoYSju9FoeQC+7juG3
gEgTNUuJrQuOElhG0D6atBkOPNAXGigpGpa80GK31w9FnxbzN8VjuIhmWVUtU42h
nIgFDTP4dB8dMZTW89uO5HsVovMFITLvPde8bDSiqJSwQZg0p9CB4QP771wS6W9b
Ey4kJhbcZ4jmI3FKwyFNk1wiyV1g0IRIWNBH+aIRgnMfAf6XdLMvrm7CyfWlBcIS
WO57KsGQUcsFbCzNLcvTUIwap6TKnsIT3Z7piu1HTZ/0D1feSzlieGaTMXP+MZmm
X+IYN1ESI1cfi82ddKKgX1yzLBGRKxuSxBaBTJ6ofAlR/IB1FlAiyNdm2OfanXoP
BDzgWcBg8XuNRiCLFaDKsx8n1kwFf1UKg3S3vEM+0Odm4ChYZiKL4ZGQGk4184+5
6+4rjJuRTWJn8wpYJc2FgDzptqoOdXDcRoGrYlkEgtJSC0ZaMbN4LLHO3noT2Kmv
OKgDshEumuLwdtstKTTBcqbS5VUfLwM+tmixIh6tVr6S5b0NNa7Jzvif4pBSLnDe
JAFQY6C2Odoy1ihFc9NWlLH1bc1+3X+fEGp2sYDC5CnJTnb99XnyXPBftif0Oojw
QsDwN9tA0cmSTkgG3opfszKrQJKwjTf5l9R7VMocXIIz+CIq5mdGa8LP+JTQQBO1
JkSLgPq+p6QG+cOCKbJkfKaRD1OekZBYPMiLUmWvEppfYRfAyPsHV7PAh57oOUr6
3jdLB7Wg4BrAHQMS1cPNWbf3GXWSUov7B7+ZdcYizAoguYWFB5hUEJKJghXNQ/CZ
UmWKFX+CA5Z4r+T4v18JlBGLZ+N6Lln5lXx8O2AHEaiEBXBnWB8hm7qCM2HinJgK
TaJkszSp9Uin7xnxi95FPlr6k9gDf7fMP+pm6RocMM6UQhbnadj2k1r6tNn71qzH
RPJ6XARNo6R8vhwVb1PDCIBCvdVYSTXnxzLbLgqrU6GTTG5pjZLsrXnrUW3aS3qa
Lq29/sayV/DAxbMVbuyNNqbHEA+GsCzTw5BvVWLBng2OAvVTMqH6eonegerG5WRf
nZ9tkqTO12S1yWvuU+uLCJzyRu3LXyO+d0aJwLHy7JpjbHSCJq2Jvp6RA+Zrwbp6
K0iggniAy7YAm9Y9GdbU4MxRlv9L+ncnFd4PzxLDPUOD9i+saoG+WIspiSBZ7E3F
FsqDC39CM8pcNW4YtJSsGkJsK9LVeAzcEeHCd/63LbEJVL1KtRvZ/4FPKaNoNGIn
Paa6c/W8CuX0SKpR62cw/r8v69+bxxhT0zYkW57CFnM1TiIScEy0M9y0PAizI1ji
OMB6fqgNgIgT2IGEo5AH9VrvIFgDK3FBLG35fkZF3Kl1cSIoa0Ic81PAufO4EZA1
qc9/qL1OE9M1pHCWrfuXkIfajMP6kBSiDleFzgdAecuBSnhzFTsOhQfRQPcXsgm6
todkB1rpRYrDcbCg12qYc70Zx5lNe8yPWGQXfB6q9WLdafUzq5f4DdApa74CIEpu
Fzz+ZXW202vS1FGLO87V9mBvK9ABYpEV8g7yhmlXruGgWl3GCyrP1Y3lCxNRGoYM
oxeQ5bY9tJeYcL9iWqwpFoQDzERYlEtxLfoIE6+8fTnpp0cBHixUiYNu3Ib50Q0i
9iFlNcmdf92JO5ltt2pWYssPJby9Aag0XCzv5mOBx8sQJlVGzlYdFrFToPDaXIew
CumICpyY3QXslcdJQqOyiCobsoqvyEvmkbnazyAfb9Ih2L+J37jFfWNc9XpnQpKH
pR2nYnciVAcuwAlKKI3Dfi7L4jstKOazhOIAhjnb8S1vmbPcyyxer1Ybb6Ywmv03
Rijv5QE70m4RMmH6NiBpuO03X24WtxYs2sH1tffCYB61v4Sd0Xgmi7YyUWY4k2Cs
yA61TKks+MGB3EW2nbLL2dQ0II43x+10VlLxDtgaHd10BuGgcMg4So+64J0sGqjm
RWHMWnr529rNhYbf81Z0m/+ehWxCRdUoKCGzwmsNXjwC+gLkvmqoHRCpYofxHL1q
9nxIahPfdyQTt+gwEN8pcnlgvRzDLIIVhOh1pw1XOm1L7oh2xFCy6MOUkm08G2tb
MrSIDljk9UVVkJ0Nvq/gePUiHiwP2ZqxsfXTOTvnchSRkSnoa45KrnfsaJUWrrIo
fBkrrGGk7LwKuKqtJQ/RTSxH2KdW6ignfV86k0JlcgMe9Qnx9vbH/jVaNfA0zlq4
qu/7PtmdXgzv5aN6kl416zWQXsGXDIF4ZZW0mnc1vc7y5gobb3HYORmC4UDHKBsW
mlYw80LvRDXHZg+udnga0w0DTqX3b8uEssqw8dz16okBYdvL1H8htBadl0G9mDMp
tIO72qAMEfqghgpWuh4ZZqHLlmSNWzXI0SPSBwpuVMHhXKtQKKw2WxQELJ1iDVWw
WEGRQXDHAeJ/vFNj4ZqvzdXt0AW1J/pGu8P/TFXfoGuU65tZzXhDb9FU5vdV7j+J
R85UxiG6V5/MaqY8mXWPm/TadiXuDKpMiABxf3JR62YD6Yz4vcc7RjWgMElvBtnB
6hFoSyzHMU0yPHiCs2piuG/Ecp5INmuQdPyN0r/GuqSZtPKxuuXVPuA6CBJExj26
JUkfPn1nI0WR9WTqy2Z9TcQ0h4gMJO/PNXBzEx5rkmWjjRGUtNdPST0EEtpp+i52
y3WI/zlEJRrCrtBfLQ9gbgebMTzaasM39ZunwCWO9uPiond7DNYH2zLnoBBQFecO
+ND8ujt7geZVIPjOWwHzSUuwa+LG3Xob15efBei9qTtDDKN8cmbX3cFe8c7lQZ7n
3Et3gaBeP9STl3pHQWITtlh0MyDzvb0gLxSV7LmMSEfq0nP6XqrKZmcd1ORdagPr
bE3AlMsO9dibKZkZkrxPmYI4BNV9wPn0xKgeHVcRNmSc8c10zB81ymJ1udeeDiEE
y3GCOrwCyCzYHvDAKKqwcCcbBwCtPr6WaHO4TF5hZmJGjy2Ku8kS/FqP2XmQ7eBW
eNyXCCpDOehrRyDbfwde0vkGARlOH7oHlXKtlma36l8DFIv/faHqC/a43QXBjRjo
klXerRdL3Ts5nuN+emAFM1XUgjYli+2S9EFtCJ1iteMRseqJuAU5OH4iZGqIHq7H
4vo9XtH/CgRMjF2du7x5C7XDyOxKlSP6GN0kNXYa+1TUNtCnGXq+FwVeTt6ZnP7L
pF3aouNDOnAfxiKGFGW3pFpSR4bAMK0GSKLteZtLxNJHl6q1tOge4e/EU6zcFH7k
z995SpvtIZl0XYgCkjhS69bj/NsUxQSYFo7PcpdfiMbpvzjNF7zwXPogneIQL+K4
v2FtCcnji5csB+q0u5IbeUueqKNUD8bDFMgdRTwMM1FnmT7ykGrbAlEP99OYUKR2
82oEqsmRf1bFDdnksnT0pi5TqBi5Cu0iXYVCuwTqG9nFgQDMoP60m9Z91I4LmFl0
DXVA3d1WZ9rByne0NGS6+vqqbCXFvf0q+1wfsE8p/aJQinAnsFltBMIUW9CDOWE7
bcm/V8vRZFevqkphmfhf87F92+/Y5YLjh6NIqXoF6m8EBRYST/qJBwObglqHPqn/
SCQy6KA9JNktPFiI7OlCe7UIAQ6msGd4xQB5pxMSAEC/FXGhOPfCs6OkikyUNpGX
ev6Itc6Ij6epIh2Z9dNNNVvLuQxaN+9HG4rRkCVkrKzBTyLU3uVhs9vWSfO8FoWh
HuWZyShcnubcJ35U9lzOH/mGVY6oTBkBOOaEbgzOwPf1hLN/CVXcdTeNtuwUdSmO
lMBPtzrgCHPg3nMxqthXgRBgL9NQwoS4pTDFhV1AYFAuUbCJl4QCwkqbhkWbd27b
t9k0VXC6IY9/pd1h6Toc/aw1XAEkiwb0p+FGp48qX88B0MhEJ1CHpwkm7YsPpTwn
TpcoQTfXrDANfnleI+Et3X3/pCAiX7RaQvrN9K46ZRzXyRpli+WlxJvR/R9tab33
XMOpk9ajjHnzwBYlveHDBoxRejq0MhtSsHd06cVvkCR/GG8YRUfbhrCzDuwsPT1D
K3GvjOBQQhv6es4lUXAaUACF26fqn2BoWpkgDsFB4HVs8eDOHYMrP5W9wYCdKc2p
KCEMD1xp9cuZZfsYtgJaivlDG016qw76Emm/oya8+yiYvXnAOdH9otcr38ODjo22
PUakj2IJbAblz0gEmqinQRQwM2obORH3DmfePZObFrAgvWddO4Ozxp5WRp1JKu18
/hbCNo3ccl22t7lXQmyxk0ZyNmxcQ8YHyjYX4NndAXxi/QOG8BqzAqVdtRqCUnpv
ATKAPhtB7j/V+frFUaq/NzcDoByBYZpjtJqHB+WQjEDY3yHNnvpHgyNrisLoasp/
1u3xTSIf8m8MtGvazxGUWZuDHk65NNdRvHOSImo+i5Db4NFJ5juhMBSsL2Lj56Wn
woUcBM+x92TmSe+GvzLoOcYc8YIHW6Hsc9gHEEPceWVIwbIOmKUk8VTjv6uV1WRy
7lhIuBFDt7CO1aECXChvPQXaDt2sFjcI1D6E811TyKL5psS/CHFb1SWCoi3FJEit
CL0BvAtLF/k1/iADBZjUm52h1qOAaoqSo8ocJkVICJY8CYfF3CP89pI0hdIVgReG
Cn6jVVYb2qAd2EElfNaCpT+dW6nUkH8Gqq2DWdcusKK1m3UwxSfiF3QPFuYU9Rpw
5UBio7Sl7tvgOyNhNwseKWeNLwQXt86fKiJ/quSA6k2imOLrWVNd1+1IQsIj4pwD
5CnPQu64WSNugg1hUQO7ROW54OOjxJwNknRaHqMp/dPAq71HG6XmeAQLarvasaXE
BOczNeFQ7FzrnUw6djQw/o/aopHq45G7E9mfnbnFWzmaEnEjnma4q3gaIR3HxjiB
tWO88zxkHzPZxdEO8hl3G0fOZGct+aK6TiitF10oaTrAfxT2p2FFpmJGTExoS+4g
plONzIaofS4GppW8GLKKWV6EZ0N/kl998lU5G9ToIih8YbwB7N90R6ZnTJnhzPU0
DQNAXHsMIeaVZ6x9Ns8J7oQ97bhZW9Z+TmH3055viTeZudsZ/mv5MFKVmF8SKYkc
6aS0+aySvvONZwvaaiUcPyemq3VV+tpHKE5XUU1M2njsDlUjKMeuSidm1QpLtjIj
KILTK+KA33N6D1ITyUT1wdhOd6X8BzNJOEj4oyLZSTE0bVnjvo3dg74U0D1Djr4h
Nwt4eXIhUjnOxx8qFPVqhKKqr40BGtYnGDd71vPtmY+zNW52QtwzDb7v0tlk2ApM
p4QyuYL3XqjM7jjZ7bRJsvyALPfQEYkFN3GqLyy8B1rS3mkZN28ko+9HbQOqhrSR
24a4DZgNST4BEa4wfNCUTNq3PJGfHPbyWQ0eoC0g5KzT4/ffsSIph7GT+UMnZYFW
O70IPffEIb4qWl4XL0dpFM1tltLD1jQU5gqAZ+8vBLsghdRXkmoSpoD2uOVwm0VT
YFyG6rBOWfTo04CXlmItHsI41rAIGV3atYVXO3sOU1F+Wemcno42PiKGwT2MTBVX
mfv8Q6IU3pLn1fcR1QrWgD2Nj2FcQeB9XE9VaEnDC+Xb5Xnxib0jLEjrekQ+IMsv
F//3E0oL2kFIUgeqslEsAhJ7naFzITFbkishLK3gj2YOEGX61XUg8ETHwTVosFXU
o+vYV2mDdk4lEkDvSl6x0HqM9DZe7xTexbvopkSXUWc/FIFiC76EKnxMSt03cTmj
5MuMS9f1vXCG7ou6y3Njr1Tb0JkwGH0ZMNTbvP+EP3IPrYpcyJRGWoWT2O1VSBre
PgItVpBNRQNHi5HVwsz7UYQZnVea+Vh4fIOvk8Z2eNQpkmz0RQDQaqp3X3r07EAL
7iHTL/esQYLhbMwOn4hyMyuo/cMV5rJ6yeZwCeQkLJ5kLl9sQ4idDwB1dE2i7E91
33EAhvSF5Yhlzx/PS7x3EL/l8mnNhAPrrUrPcvazhnLaTYJc5VuVDUjfFJm7MRaB
2efSX59mOW10nMoeAvarrAjmUNhcAMJZk7x1C2zyyuuICv3/+juRCD7/ADzybOv2
O/8IePY50koNh6JSRfdcQIz9ut3DLahadv3wTN2NSC4K0WSpGwLbfOBrxkPwg9Nb
gsMFcQHqjbnwhRw6P4K1zFGqOZAyfrdkiMOuMXkkhVNU8+V0aGlw7urgjJGF0EzQ
NeXGvDuwuhpwLo5qnuCtKFndnq8qS6BUXZe5FVmoDJbb0WlQbUqecfZcX3CSk/Vs
30ve5kJ2UNO0KdJVGBngVaQ4XjEbgu6SCLub9IB7cJLTy508vP6m6Tuyb+nVUQSl
6ih6m/k91y+rLdIqY8IMHn2yE36aDNp+W6NXOYjnQpoY8HT643utKjBw1dUUAlje
pLPfkDeXLJZ1LusClStmYAi6uhpjNAqD/RtMxlCVHQJIxwe9jXY9OTV8v77nwdF6
q33G/aIZx/HdIHlanowEllOzdUGHPSL/lpTb1UlsaqiO5VKFw/7+ljhReZYqzgnf
+2kibuAJFxkK+hfPbquCtUmPrPG3Ex9we1FqMHZ+KMTgS7zBbLkOhbCq1a3igvgp
W9x9BoX9pMSsSEEyluSf0rbErSpt7ccIjm8vmtDdrPvNnjYCYJbXr68e29eNKuwA
lukH0+QvtTDjnF2CP8klzfQLGa92T/h7IyscXeVlfCNkOQg6I9Wf5Dk1p23IrolK
kroRHdQKTqfQ+MBaT2NyoB/nweCvSJKCyOQkrKTGUsvNh4qc8URvQJLsadngkTRl
e4DNrzE5/t/esYiK7lx4o+6+wm2oA+gxgThBr/YyE1s9wTLsMnIlQVBaKbpEI/Dn
K/AIIbo3I54VaxLZ5U/faGuLiCXHaHvgAJAgCmz0k4VgYQ8yfBmTmVXmRR6VT9DY
T4XO5/CTWCn5UZ68MgSnYvTQj2GUKah8CwgG5KD/3v22MmUdf04gFcqdqZJ/MEha
r2uhoOTQvTBCD/qza+PrV6SUgm2AJrKxICQilDMMaYkHCNItrCEzcMN9bb0B5Kx4
Bb8D0cmoEZFVZbneZXPLCY4pJE/EsFTHzCCbV82byjztwXJFDvoLSFy5BuTjZ7F7
et14uwbDEOul2VOA3bkpOoSGT5IdE9JQraoy9P391ri/xrfCX+j8Zu5BVFbrRfrt
A+CQmxwkUesJxSkK1mVQw3tqLH4xWewhEZ0bcp4iT1YEQYaOwNpctw5IvQFgVkqh
ZjaWFADDp/aK0W2OD23XcFmKpRZmkuGg307Fi8o6+KZ1fAmmEikT4VcKfNL3NAt1
fZ6OKfdShjYoiTUP7/aVCoeKm6C5cCT2LmIoIBdygxuJNpvOq1TfvbfBm71LnsVS
R5J7bHLWCpN3L5wpkD3MIG01021EXxwNPF0pGfQLcSZTqWR8gT8b5WbQpot4sQAU
8ROVTf5OX5VEEJoPINOdXrt8RfSJ6rfIUmYczvxDrWI9OIwOO/TaNJqVSDmqct0q
Pz4kJhrfY08Wg4HoseJL49NY/WBvYAwU0oHIuZsMp5UhoKqP55nraZ9JDnIetOYn
l9qohHinIf7n98it1+XF4g1hBUbFV1A0eD/v5u/d/M6I+5UURUWFIh+2hs1c0MyN
5Ew/b29Kr976M3bUgHgZC+LhZeR+c7IT+7FVEX5UEB6SBsTeYsRCZmXnzWF3COMD
kEgTvQUiWs2+91+5vra6n1wRydU/mAt8PDvTlkeq1toivsqk8T9yCrq+wgL4RDAB
+occyvxC6gcJvLEmBClWnETSLVWtC3wYmECcU8fKD0BxKp3YVncecvLDU5+dXvW0
7whcZUrV6j/GLHfavcPv9G5h+5or72y9Qe+HF6ii4/AUocpv0rM2DAM1G5A6v2/p
BhArTfruUjVE4R8TMhwSZvfdLgWQB0aqxxk2guez2TkkqeMblFnlvGwn1c+GY7nN
KiDbIViuksZ0Agcno9FyQc+Gq3yg6vEG1eGLt/zMQ6aQ/EAAADNMexReCN7yyZAO
JStzfZnkkSBhj1QIpih7+EfC5puxVOsi1aA3hSyVp+F0nAjbgE2DC0xc+1p6GLI0
68eZWTONV4whM1kS+ljHi5yiUVbcy6F/5v0nnE6q7p6hjL/6N9Xwx4xvie1NIBiJ
svhQconw6ANFM9TNmyTcDjWn8ozVF2hJ7ciOyLTayx4dpp2AwWSspM2LMs6xnGZ2
AUQm7wkZgyvXDAYgt3oPF4zg5uaNqvmygZSE0bv35LysOkPw7DLv9852GgGP4nAL
l8dVr23EqUsYAUJx5sSEJ2689nNaDOfmOIc6nDu4hdpI9rpHPggb/fMxRCqeSLCU
qihvViRjEjjN0s0FL+gsQh7PLVvMEM8Pp+1RMerAUwLydvYOGvt+ZE7jsEOtvhPs
7CrYxTcgBFO3QnIYdUfK6btzBJXYvag6rgpr58QEy1JZvA5dT3feCyR/VcUejePq
MYIrEOBE4htt1uJ8Qw7MOFD0yMUwe/P9w1EX4a399VrIt6Vg3Q2QzzdyU8EteBH0
bFh269aQiOuiT6KMZ/s+7mxEC5FypM56WKOrxi0gYn4zwORtvg0dcwAaHMZThOZQ
W9adOZEyryZtB46QS+QHFZuHeC0Yyn0fHFit8z5G3FWelspo1Z8RLWxv5Enj7vEG
0rmqsz48xNErFJ3FXfhATdWUx4GLGAp/YVUelgnFFzh+hyyL7wMbxqaJ+WKhGdlJ
B1UdQNYQbaGdLe2EseH/yVWGIifEJSypGZn6tiErEbQitBGYQ2wnHw05iXBFk72Y
7qtagyz5wEB9NH2nLiVxHwvUrMlLGc4WCmJUb0iXi5IZHWXiazeYCcPEtDc8+DH8
ybaWp2OSPPN7YWjjlI3x1dlVoYpMyJDPYltl6301sMRz9I0IZh3GRjTp1Z/VGkaU
TbLxQfgpybBn/yI7Jmhb07HE5xH1iTZKMHbGzECezF8BUw/FDWcXp8EIJAlpFB1m
Ay7ji+utTW+Y/DXT3D2k6bTC19R3Eca89MurJjBInAnS+LXHoeLNIwpnDPnGg7Bb
Wecg+rJ1tm/eJg75dhb/YRz2/czrT6eYxFxF/rjB6r1KkGF7WzBWC648YyNIpHn2
ws5eXFDjY8JeMPWP2csVqQedJ7lU/YkoR15ghkroayVvmpNdZoKAo/xmvRZQW3SK
9f57JXLromUTKYnI1DdT1kg6gys2hjveaKs1JbMIcriWhA4nwBewa8Z8nNEQpDoL
HwtWu89sbYJ0Ohz1McA1KTEN7jM2tjr0xKlJjbtkuXrXy8qB/LsTUkp66MNT+KkU
pvc6TYq4FeS2NDfdHNOfz0/o2U9t6HaylcG1o6CJBj8qIM7DKG93QImATpzn3zTv
Y4YAJh3PwQJZFeWZIQ3zYkqvLE/8y5mS+dLJL4hh1BSjuqeEWQfoSI85boyWHSo2
M6nTwESEoBpal2vEbV/YTzdOl4InpEwB+bkGTCJfkZqs9T8RHXm9817eeJljnRf2
GqgNf9rLGUzB5LPv9rJjVHJIUY8wi6OFCimkjLq9fqm+avpyLeCMLz1hHWjNxrn3
dfEEpqZI4HPo2pnAzaLwQjYlqgMHuO6enJ0395mQR+IjrX5Eyb3XTp4aEWeRC7PK
5cPWRPaQV8Ix2+0YTUkypby3skZM8GIloumwJB3GOs6ldTRvnW7n8KqdLU4mF+tL
cjtcGPqliHh91UHw9tK4cIJvJplFhuvGUGX3q7ml33w+hnolxuOYwe1xaMblgOoh
CIOG0GG36R3o5BzvyyiuzD9UX9LPpyyIp83iENH9zymq7/25rA/7aYaymQmKwLoY
Pg5pRLqAOkNdMFf56mJtUN0/NVHNalRm8xAKwYBcJ+wc+laV7jfRh5DCR1MMFzJu
NOIPHtsmYC3jgq/fal4uwCxJe5hS2Cjrlb2/dUKzwMa/bb7CUv1xuHmbtTH7jCze
p4Yf2QcnJJk+8AiTiAhFjhh5jA+jkF1NLM+akv0clSIWFx2x0Eyt7S1eSTVbVD4E
QkWpeKr7sddEm1QNgm3VBi5rAr/c65g1YFFzM5zsdkcuxnPryVvqsMs3ZsA0aP5N
Dtp+3IjSfEuNKche9i8P9IUdh2tiX9Z9hRjWEpavVnX1kBKaZffbsW5YIr4Dr98j
85LMc/xipJifvjtu9VqGNGPFyNFby8KW7rBPfyBqM2rLz1fMZhw/KKqvn3GbEmhN
HTcqetHC622kblRJskC9PZMlqXM5i9B5iYNx4lYUVpEPHeWojGp5Uj7MGfE0NDsr
C+2ugcB1XceqIYHOe7HcdOj91hNIJbDninMrGTJ2Cnjh4ILEvGLlN2Cv86GfBAxq
nl9ycfNnLoUsY285GGQzIBM7k793h2JcWo6bHtOEFrjm4VwcHxHB6uVzccxCqtNG
jn5QOk8yxiph24Ccm2Gz1hj6B7iOjg9P44iXrajb+kPlQFN6i2Sa5LrZ/YigomGr
SqeSHEcDhF8r6C7dcTz91vTK0W7EERxdml9tyrObtn0NR0XcyTlz8eClnaDvOzPF
t6akfu0DYULqRawVMnRdKnQQVY6+XgL1/b85HaiH4II43s4RmbcDQJ6wUgQUJKHA
ukoUtFcv2lAzayPM+vdMDT4mG9ILK/WJY2YEGH2bNSnfS40xjdzspMejXmAiekRI
ucTaGkxbJ/L8AbLo82emBE3mNzJYfzscgbn0Q0syV3eE3H/hekeVFk8H5J9GFXtQ
5VpPvEiWVm5xMS6LXV6TQ8beM0EY+mZQRLMSYps8E9s4D6CuksynRWoUrwkv5cdC
qrabj2MM4BiMsYdgdbuCXLz+HazlQWbGeM/NSI+plNQujT4Vom0euUqwc693+lZo
YYZyhsffsNCCJnfFYPYFQWGJKuQSPUJBKm4ZsTbuZAh9KpOkThKUxBA9pFNeSz5z
NtpvQuEJ6InzBK+3ZzIP15mD8h3Htlsp0m7P/OpmoXA92bA9Ue38WUz6XhX6jkLk
BOb4Mio7eK5qWZmkaS7wspW9spiVUxelNN9aq4rGw0vAEHAl6NJ+yTnqcYAFj71V
XDWsZinDxDNJyendFu69uABstr6eZACkL3LztdNiK1FMwhPm6OAbrE/MQsOJJmzv
mu5UeSP8UnE5e2wkEKzGp+XygwwKqu8IBfbAsxz+j11WFq92oDurg/uYId9DBiL4
qKhorbwJM2JhRi0GGq4x9lg4jivKZ39g42VT9TFyeHl/Xmpfnq8kst9UNJOWgxVN
Fck/ZIJFlHQD02ILxv2YhvKKghz88r3VSgYznVyzEEiXpYGBWDr1yLg+oNTdp5lp
BpJCc8aB54ONIrPHCDkUYshdwr7EsD3TbE1dp8oZKYMjFGIcp19auepy48IRzing
gjLUJVOTH817lBAzWMwSjoqrX1Xk9YI+fPW5rUoz4sudFaQekxhxVgDWAqz/b86V
kjKdtUHpCWlhuTVrEo5Gtk5fQzEpLInS+s1Y8TiWzXxtBOub962ee33aM5gk+EoC
Y46rFwpDHIr48rnQychFEbwA8gD6Z5ZPIiv5z+9ljG7eKJvU8MJFdUg30vY+iSrP
UByqVxqvNWBdg8R4iYMNEyqfWBvw9BlItK3ddjxt9+q3u5fEGE7zHndSQP6Zy26A
br5+9jubjSizpB32dnLjEr0plnjULf1nocvuqPsxFRkyjs6kO1whKH6gDjUjYymg
phCr/+AMjuNhCS/dbbuIRfSYpzTnWdLffFWFZYz1oy60KHkI731GB4+9RXwv7D1v
atS63RS9H8xW/JwvL2lG6op5mBa7xT6mrfCQxOo00NM0GYaRK6nV5hO5iAGSPPp7
GWST3x+BALrXvl1wghQIHE7ciSy1ULUsOIhX4dv+F53eR8s5a3mBkFAASj0q6r3k
TfFOxylUx/OW2qtp2rt+5DRlKPy7+6xCNxuGLThkI0e1mfl6mgo0qINQaKV91qDl
JVMAr21kRecDHAdzLK2F7+T9MvgWyUAezYrddHkHEdVbXT49VP5VvGXwq2jJef5B
L84ZSdw44b/wpT3EgOBfqjm0AQ58mCNbGpdNjkDtTGuHHusI2NnFTFqzJauTkdWb
141VOkEXg0vHTWSzmHsgdjJyP5CFh/TCB1DBTC2Eb3yeOH5rgSLf4OIdC/zx9wR+
t710mOeIrrwamK2ciYwpeZ58q2hieq/ZuWSX0cZaer2dHFV9DcHRBFgwc4QqoMPN
lTg1fNr+NuqdNxhFeuZ6U1/TT9tSVW0DiWocLXpMd8lvr1NLh+hmxXLJkcewpirw
B7HCMNZYqVhU9kP+zaHdmpuYNx1kNfQXHF3R+h2uM/1RMqDCULzaX0F/VUEuiWKE
lYFaJjxkIarIf7girjQk9U8wOR9fpxidUMo6CnvyVmmRL17ho+2hya5yNsate8o3
/LG/feSYhVmdz6Dn3RtcePcGIGn4+v7sNrGuS5AtIopTA6Muz2HOxK8GDh4F0u8C
tIpJpCokDbGYH/W8aGBBLvh8TsXuL9mRaeyazGIjNhmw7AAEHFLrWpwO17WmZiOU
yjn1BEpw/x3jTmXbkjHVCBFdwReWPLonmGDpkvUJWZUx+vL0BL9a4HetdAzLEBmx
r8rzv+8Lx+Qq3OdF5hi4Ohmo2Khy8X1mDHZWyRQqwu/DFDnLk+5caL9exRxxOOIg
1qkjg7wO0haXkqHIUHMCVShn2FKngDplBEGNYMTefMj9mhXsB2E2smMzoEDgYUCE
tgbTm7A3iU0y4GDeBq6AKaAEUA8pN3jMZw98ybRV1oeRX9GCbQN4aR11U2s8o4FX
ph99GdTS03NtiH/fzkWbmnElRhaOKqXG9dpBEHHRGWRQk5YwPm1GMNiDmGeexajN
FJNZTmfrm7c1ZAmeUeOn8+4aWYW+KqTMT6/+eGxzlS5eKFp48CnoKtpDjtiEAtPA
/2F/hUn3P4s9KgpL+o9sogaNpmmW301r91VBulZjrqloWZuStR3FsEqflq3k3+E9
QbUFqM/Qe5umydMsWMCs6YNm+HWJvGXrLdJNYQmpItArhmg88l6guQxD65tvCBvA
NM2O7OnpCrVUA1gOqlmeDIR3f78H4WANu/RuFGrwmV8hDqmL6ZetRR0ugRoxBa5g
xmhIZWvqUgN8xhYlqMDM7RwbKT5tOUdEs2Nen9z1PcM3IlpNpiHvdm3/OXhHYvSd
3aDsASgfFQ7nePytXuTpiZ/78LXGnIYNLwxocBAhvZNqceo1iPdn+CwAkYoPzMCF
nGjKVO8APmq9QSL+otuwGjqd7wdpxKh07P+GtWwROW+JzQ9g6v1TeL2wdj6PLWuo
ST4uK1dtGTojfg/kqIilBNNyDUQErYkfKG0yy5wbvuMZkJQ3K2yGn49zj0uQg7KP
eAVELR97WRryiElNgVpAZXpGyYC0xS6jqPhHc+lxUyq/9Pl6ixGwQzgl9uR0faUR
48bZ11RL8leLdRNQF/Zy2WiJm2VJmKQt9sCHWNYgcl3KSa4RomSmUovIz+tcrKIF
WQIC/ibI9wBBL+TBGWR2S6hZUpJ/iPu9gRhovO6Ak5bNPCND9BPXjog8kQMtD0oS
pIJSGp1CzdBPsNtMXG2X7z7zbTy08b8g43TS9FepLgYxx+MhoBq/tzsOjRSJ36+2
LTfm+9phRCpp25acea+mD+vxY/J7tVFhn1p02VYDxjzKIwVMWTZmTAL7F848dnYG
X31BC/PZFzOlskAmVtv+YIp0XSiqjGEVLao/Sp1fNVXcetRF2ePK7HG/Bz5FcVL4
gR+5XHEqtzyf0R8ZYRUDq/AnFOMFk23CUddi7Hq2uXOzybXkZ+sVtgyAG86IeTYf
CybF4E/bq/mYcoms7H551KMFMY5aM8FRUek7AwvN7crjetWKJKKsC/IY/12fq1Dd
7UkPG5ifW7LuV1xc/YbX/UbLB9ds3qGv/3ZY1+Y0t9c/pzZpz89yUDLcnwwO2T3p
QK6uDHdP7qb2yjAWY6SJeTIsZZE4yQQBqwPtXNcvmn4ConVxwBHEUFHFTUsPjNbv
GVD2R4nyBMuQCk26q3UbOd8hkwOJ1uQkmSbJHtBa4ijjIkD++bGUuE291AUtWgUO
W+ubiWhTJ7p4qzJ1bdhiWcIfQ3cNmL8FRXhSbeiasCh2esr6wsb/c1Bhh464iVZz
PSLHTwNjSYA5f9irr7MhZEW1DskM4T8Qc+1XW5IbVl9ODXPbUtiiSvjb60yCDbV1
WNzCJhnug24xt/hGfvdHpZhNY/o+lfqwt3K+rgZJkkec2ikSylt77IQMNyYTPSx+
2kMlcuZ78NasTcDwKY1vuewFmRxnldlTotBpsJJNSs71FICvji8tx1J5aPNko7ot
4SikVtX/YREMA0VgYdPN5zlQfNleIV/bsiDgl2UZFLP0OsB1lFbntTLMaP221qg8
/Avg14CGHE9mNRrwaK3iAiJUJYtUdm7W6vg1OMOkdwLAM5oSlFUPAXLSMOwM9T3E
d62/fwhoieVvMDRUi12iS1mJ1NlV1KZfZ7K4YFscKAjDdBxpcEol607gamyOMVo1
uNdjWltNsixteUhlLI3SfrlKsdhrO9U7FCbeiKNo54ckWCcZ5DLbC19l6L01/jKK
haFLn6YOMhMoKxdU1qGuxDC0r8va7pougHyDstVsQ1LOEilK6XYJzJJofrPRuZJo
NnqAq1PCahCzB6i9tx7b/eYPwekI3HCxo7dQ+jJU18Z0oAr03xPf1w7YTqFcrOIf
r6G+bVNvgXsb5OJpG+EVzlJNFIC/nT1fwbUtXD6p3lpujsrTU++XIZWseVtMQ3/H
QlAMF9w0GKvB/sTzwtUtSMu8z7Sycydru53/sDNx/2OSKYtmIW9eTUpuSkv5363C
73YOdKiTxbe3KfMF4Oo5qoiGO4ExrIVX6pVmZGKcPGifNiKJRhugf7bTI+kGlCKh
4eXJfAx7BQ71cCprROf50BUcwRkqQu3ItuzYB6yEfjeE0P3Lnk30950aslMn9cUN
ipyqdOrAFERSQg6AghssMREhDHU7ctZefhN5cFzmsks/S4A9K4uZXWBL0xkM+2UM
ytkZKVn8kvvlCU5/n07+024ktL/eHzFM7ckc2kaBGIgrP5nzN7WN6BZV32JM3+N1
2DUTiReFk4M7Gnsu3hD2dR/APu7YbvjHsYOV3Rqym3M5wJHFHl8gbMeqxRX1pqQs
X0HYRJ5V3j0ny1BpF0af+TPIY26KbYFu3d7KWNpK15Frpuqnj/U2/uAg3Jkyuy9Q
SVmfQSVJU56DOK0WpW+mkEk82jUcAn3bOMPa1HbU0eyonxoqqkdg1mKFP8JPn9W+
TgWYZ4+CcTaAi87owxvsa9Rp2CzeCAUK09mm/yOmZ603v4uf7ztXkqYRD1nfyWzu
bm4PilW+Y1ulD7oE2LAklMywBMYH6660Mu3XxnUP5AaOqzEcDsu1SfW3KQJzctci
mTKgnDXRPUVLUlZqeIK8yXvFzrQBwi6qKk8vSXlGChU3NeL994QQIGJ93/x3p4xZ
n8Zjwgywrzrdke3H9SVr1w/slT8A1Hi2MkA9gy3yPUz201ad/RSkXBFTcOt2hovz
kQVoUgUZmyvF5HvMeqBoQ+b2QeXQ+h56F+OnXwGIjprOpzOkjwptZtHOuRBivdBI
DLCyF04YAVw9TpEMVNAonloJtOoslZvgrKUDAW6BS35yD1EngdJ1yxrWEvsz43tI
8hnLrq3Sx7AeRbF/ltFRC0k4tHT9Qai2yRgssES3g4T7uQC2MRdGGoAu2ak5LXNC
QYs4v/5ilh+wLyh7QzjkBkLA3WZ+Y/TPifMRBtku26nTTz149b2vmLm7ah/JulNZ
R+WsrRgTuna3Pum4tkDnJsH6Aqu2d3zKCBQmFdjcXLu5lMF5qYUML3o4cGAZeAJR
9xV3heorJOpc1cbv0HcuoLnurX91VF4lORvYX4EGivqFNSMXAzU9Su+bvjSDbo1C
dQLtS5ZH5iyQJo0ghiX4ctxJtVpcwPsdG4g6FNL1BE5XIw1yftZnov5KM4N1gomX
uzOt+6Rm4RXck6TYkOV+yRGERC+bghwHfghlKBCf3wsL8cLw6woOfaE18eSlCjJH
xAlsme9ld5BHck/ff7GtjtLvQRdEQlmroyzt4d3fXpdfM47lcMUTimfffjKaN5ji
J7FtUGtxhn3srCw6McDrNFeW8sWvQK35LBrCC/nDfdG7Jb463SWhHOkMpH47ysT7
GDbMd4BGkSXPITLJo/TAx7bq8jYiIt0ixdVX51fQwjiv/naf99Ku8L1AEkJeG/+8
FpohJlE6bWNs9Xcz629oKE+KOfQ3CXowRw65r6hp9ZCuWKIFbVeusLpQYxxaLYTG
DzNcCZ8xM4wOGRv97xUNh13kgSPWGDDjXy2q8Cpp39aB9s60uzMH3sNSfULa5PvK
C5Gz/6fSo8esKUt/76lN6tLQVABrMrItjrUOkS5EFTGX7PNoA9OzoK1972mu8Upi
li8ahFIs7FZDM3LaKwPaZv9pdavZ6tfjUJnrw+DjgJC9SpAqxKTDLJ+lRCdL4xVq
B6Pv7NK9beW6hQF4ichaQjYsi6Y3d9gxhDbttriS0NmFOotITOzFo9LkZQ6HjXrs
S8ujtYSOPzInoRjC+wQbmBDTW11zzSL80Qqh9r/n4CUpvn2+tqxHd5dX4SG30OdP
EznqNv0+FupENUU4PkpYyZTUP16TtdG1wnG+ZndwA8L2v/MtgpJfo7k5xflY6y7J
3oQ/v+qjalEb2dbdC3g+HZlLfXK+Q3cBXHIQm3XpRbfsCNSGUUsHq8o5dO90gZwV
pIJ/M7M8qlDflUEhyjl+LAm8wCbPoch1pGUYETtXp6B0jJ6LemMkiDT9UQs68Mce
9g/9+nJvOYqEXD5C3t4gS31F8uCGCqhubnXmrRNtozTgbZ1AgY5HcKYCrPIwcbFb
X7/4eS16xJ89+FWLds3RhtCsv070b0qtGYBcmxIMo4cnHuWTfZwJBAdbLP5ywIfm
BJOJU4kNYhR638ZONJUnNnWx0+dhZQro6GZ4IPU3IJ5kucJ67Hk6UfWbC60KaUjQ
ncfrNyzX9xPMFJSJBp6yvDZCKgxKf/W+TGBhGwDVFreBtoqsgPiwjkK2LEOMkls6
/hRW/gkpa8w4+7QdSMk1iymiT7VT27Cvt5dD51qBpWoVCZGA18CGMEI2SdwgKcpW
qyNn7t2vRZ6SBEWnkOYKrho123K2RgdQA2NGbrsQle0HrYMm0qsdk/Vef0+PiTLF
I0DzpJXqwB1whHFZ+/ynOaMyn6cJsiRZ10K3PsBDTIH+0m/M0gC+tEmIMleYZyqC
kMVgwKpCvMiv4Ck34L+VPtYO58QNL26e6ksuH8OhYWNkmUhgCiyuhamsoZ9tlv+/
08GMWttdn/Qd3P4BmLs51Mx97+gUDnKm97Zsg08J0oLJP5RlXTDrT46WQALhxobP
tJggfuzUnDnA36VGiXhxelNrrASCatM1DCeh1PYz2AgFKhFRfhBl9kZfBNhr2qnk
n9RU9p9K5EE4JQ7GQ/npwY9CoI7OjxKnoO+O6U75gpZhztBzJBUr2WzBhYiiw6iB
Ianc7w0ukevbuXYje2T3sPs2TYTFC5BTsGcGtcpXhDPsUQ9W5l7AvbI+N4wJulpG
6RMnJy+on1+ILogGL+Fm+0bnybO5SkjhTM+drzoqppOVro6UJwaK4B3FXNBYgkFN
zgcLMF8L4OS3OCW8S9af6zzOw+OTMCCgD0NJnjqjiig03jry/khEPbEWXhqrpraH
eeNZvrkWAuDaPU6ORKWNBiWyG06BpTg1zYq9pnxkjnkFX0FcpHaERifhdTxjOCqW
xFRBML8A4LdwsncUiNKIZKQqJR3eFVmlpHcTXP6wCU8DDNFNpNahvmpLbwKxcIey
uofNy4GwCSyCsM1J4etNWPIEZDXksMp9StAgo9GFiEsjbE2Nn+CjU4oSUl7qWWMf
Ec8PZXJNmfIW0rqQQH6t6sXohVHiPactpIFk3uN+5xalefhyeeniNM4jAvfDwkQL
ZhWBhHdzS/YHjBtm/7HLe1Dy4emnaz44cTxMmEjhdYnKMG6V1+n4NoJnzyBOw0xg
S35PcjFLtMjbMQ8wOJvZVIloHRIOR9pBllPR9jsGmZbMd4XP0AhmglW65TcCZw2v
Mnw4E7mQrSwaLGcObM0R2usXIdOz95JehI12tHiWIJwP/1FLjtg7K9ZrG+tH96eL
VGAHEQSQtiF9CibS8flW9FjEEDbM2JohOLFDDQ9d79vqU9hrkbOyAIh0+S+mifv8
X9UygW9VmVD+cZzRmGVgOYnT8qBlaSk+1Yxhynk4Tpai7wmOfSGWVxMT8tZz8Fs1
M1G/uwbaanopBb7xQ0IHLfPD21QsRoGAKi6+Xna3IwaqoWCx45JgaIEKnIvWeYyj
Cq4LyeqBqunj2L3K9+n+T5XT39LS3sSaKAv3aeS9mH9jaNrBPwYifZxW/ZXt8HhF
PcvyZLlkdBNpLDDA9fGPwpxFd/b9d9cUAgNWMRdUeoyMuBHjpEezgDHccpVc0G27
aUh1+faGc/joT02SolJQadXUoiwX43fQJ3UhkemMctX35CCrdXnng75aYmHCJgQV
FBfsU5u7yRI/bQE7ICAF2tDSpef152reyhw/ZOievPu4wm85Q03yl9Ij64atBoYe
GRc+RDWilpZgdmvY3XNSbIT/uFnlVhIcgos9jg9rJnY3I8c8BZCabvmkOZF8Xgyf
MfzpZ/6AGgfyHOotdn1elzFnEupQ8BIq94ZfUBKcQ5C4IdzCs6LnP9O8/mccS56M
uDnjwzwE3NAV6WxJVnlwaDrASYpb7GEA6ip18+geAqQPWEZcuOO04RaKZ+THiNoK
2FQDV69USX+sr3MXN2iW0lBSlBIX5scHLqb20SNwM3HErQom+78PvDq7tpeiLoio
E4h7Ywz71fMglfSob0fKCQviXkb9fSnp7uaWZ9Mgwy8hK5ZuuGQazSOAtjdy5efv
nBFZeC6JgWP8qwm/kPZ8duCuzvwFw8UBS8/vtvOSYgnBMjmT1z8oI0lSxuqEsm9k
VaI76DmxVmuurvoSu33uqeAkc1WBYPo1u6NRPnMusTw53hBBekyKzHr0+DKNmNsv
+YIf3AK34MKTGrXF5tOjYiNnr1auKg4lcIIuPtXEV4VoubbBcy4IWuDwuvwA0mwB
GSEhethgY83cEgFCuOSUReT6MxksdUcbaTPHcxhjF24X/TvqxG8dzINOuxsvNAjB
ReWd/k9NbDYBhSwzWKJc+BZFpZBSbeO33eoGBet5gzm47gsGqZXAFtpLmrXM2znZ
bvsboNAJWJLXIWIR0MjAvFf7Cz0GDlRFrBiqeJgGxMxNBTzDWoKS4fyYZZrYgWBv
RRFWy2RuiBC4svfIJHa8EpYueWB6Qrd+mHtP4eX8fpvp2fLvn2S9qj9ONr5nKmbD
KurfyD4xx0hl11XSQ3esbNVzdfqv4GORJbFBpi+s5/LM9fwAnT8hjWEOyYbbC4g5
JPAffYB/R3r/jOqxCotmrdROyp39pUhTwjXDEnTbiOYGLYWmx5vaX22i+An5+VqU
20TrMS50HI/61G+NcSEiRAkydR5DJCzBuiq1uzSlHuVqVLZdi7FWwEKCusD8uNDd
GVraRYcDwaDJnZi49xlMPPV2d1mcxCog9ABP8NAVOJPTRJDwAzfJTYqPmtKV+S9D
+dqrrn1SaWCUOhmNvGUXGBGTNF7/27bzMVKmyYj+9O5CiCWwyHleWHFT3kugaWsZ
ZolgpZJKXqM1pjeruyNMQyxyVkcmFnHMFEvls7SEdpfqBRddCxG4aCFfAK37znmf
o325H2TCax6c1pVI0IieanBq4v0nq5VWB1j3Dupne7voC1Qr9sK2+nhzMpog1s5s
4gbQF+sIdcT9uV7uHMvLvUt5UeVfCtEI8yVRWvJyONI8fz8EISbQiztrhAORDHOW
1NerOWOEkXCT2WrgHUo73cZriviY+EGcqLunph+G/MzVA6iynLNWPEyNKvdPF7i3
yw0xsHNiTaqDtnHb0ddMneahh5u++8f0O1yBwTYHUK6MWhBtOZaOcYzo5Dt4rwYE
T704Bjjrr5gHUN/oOsFjCjTPmUzRKnEa4CsufOTyjUdLIhuX0g3ltJgmTQX8wq0+
qN/54Qneb8zgHR3oXM2Fp/fcDZ7sqe2ABJEt9TmyETbqL93jMzH0vPzYo5HufKtn
5rFELS5fsfXsWpRC4Ublk8dJNx3mBXZ5ncUi/7hsjw66XD7XlL+aosqkUHSB0VCs
rFF7S4K/EvOuc2vsntIq6XukOFB+0c9CgMPrsOpXF5G+fKyt1q8AXzJ054cFA0lc
I38uEl9C/IbfjWwnklXWDYjTrCb9+p0M9fjhBc5a4tAsG1MnZ5C1BE5IWejuy/1E
brICshMFpost6jUhAi/+T/aA/4iPPNz5QG7UnG/CHYryn/gX3SW9HtqtwjMj3Fn5
INlWovx1RA9Vgs7gQRPVHndhj1yJa892JAsanPBkS+xpg5WtQCuCZgZC0b1ezUw2
deHvj7crym4CCnTRzu1HjbkyyfPskEfr3WIVCd9TDeUpb9WSbDkB8vjsVCRKRwJL
591ajjDL23EHgy8mfajHBj+l/ylpSxL2/UTpcloLvL56lowPxjoecQmIDjPLkr2b
YdwduaAY6LYXF7yu0rH+S62bDyAWMlJmKHmxuCi8F2zdhle4ILsYu+NldKf9uT+I
EbxJrL9qhd7ru3kCcFDmVLOGAzDnfD5K5dnGOTxi894Sslp3aUExbzEqrNn9cTyr
q42/dLYhGzFE3mDWAQmsxAM/noa52+NGCHzUol2CBeuw9l+x6YEDeHzWjIr840uO
dn3fBS5Vzg6I3eWkznks4gKbRFKL28ib0Fx59Q+s/wROvrrdvmWuM+gqoWI2Wk+h
cMf7gXmsgc2DeKRk3RcOEkwf9mgAplaVfh28/4PFN2pDUERlbCMM6CyFcSo0B4xg
Df5AB+7zzURiIKzEdJU6/l0l5cXiiugUgpU5U7+6oRj645ALQLmQIC097RUJaEy+
D+iERfpNcHZyJ06u/krjonZ3R4WC6NC6qTnZjzOpyLPGv85Uy/eC2hC7Wf9yPDTL
AJpvhLx6URq/4lRpddxK5fiCLt20xpaizVSeEC+IlMcPF5X9Jf5b/vqR0iJJj+GQ
fBgGNkG3FzkxfkVgj6iRYht0aDYW7SFsaswgik+R5SzKuxRfU1TnFaTdJlKBu1T9
p+EnKFLJno7eWgDN65SBMPaLVicSCY2Mvr4gOTA7TLuQm5dNQky2wzCWeLXVa2mV
Wk5mTW/ajyIcGRWHvbp3WPVm3dW/yF6tWOsHre6edS8Hb48vL+L4lBO99+H10jnN
RQK2c1EzVnA0+5Z9bw5PY+wdhu1jokRHYIsjShaEeWpwn1ooxDTQ4R6CRnBlw0rK
TxiFMLWVjbWA/zHAs80tnpBgVprTnQF6mmMqVe6PU2UgpC8DHrF2cPpQSxnYqHKq
s2tmsytntHCfEZWh7QzmDuU5KbQaM2zFZkn91ty1OV7xFllu40J8sNjDU2SHfvLV
8K2fuma58fd8vwrMTSQJ4jUBM5mhMJAU1CRr/APK0O0TePiWNNL8/wS022LA+hpJ
dHhQ8oQdtWp9rGM7hVhdY/wERdm2hwN+qpPvl86STW9NYArxHpqcZDzwA1z5piU4
vdCIxC58EDqymW4AcEaw4spMwEa8GpSr9NNpnbeC7u485NtVAkHJ+2LI5HDC99aK
mhBg/Ux4hWI3OE1vNGCQZKFQykoTxGIEEmA1kVxPDps+vITopwgeySiGLsOfkKy8
ruf2TMn8tvr9NYmTUYdV/BZuhI1NFrPj55hWvCRJyHzmwEZDbEpa0umj8v/CyFqP
26rJVnHwhSEMSre+f79MDa47TkC4Ddc56MYznKtQQWV4d6180XS90Vqc97R3WnkN
5JWRLnM8kE8rScXxDvqe3uGVvs70Spas9HSC0UE3iI7arVUIbmD6dS5DrfrMavTq
wya+EqoIm/7Yv87anvuXZrsDhm28xcyTBUK3QivhEL8OtYJP0Pi3eyWPm3FyN5ps
bWvE1Kho/3ARc8eWKcab+qup3767CgVQGLZW2kVG7XsNHp3qZ2Yo2wt6U0qYr9N8
pV+CHqFyPqn/ToVxjUiQ+RPKl63oWmpEsL3Ax/w8OaRsHhYRUaT3q1VYw4S4cJSH
QDVnWY8epsGzjp1R/XdwMwgd9L6mqhyF3HCJKwiR7z/kdz0sGryZ7r/Ejam85Nz9
FNMq4Li0tikqK4NyzG+EdbKrjyrtNsHgQ11T7BcstkFd9PgxdItojuXiqc+/ZIGH
choewGKDSY5Aq3M0LKPnr9OYuSwtX2yrnejpQxEh/gIX8r22ihi5EYDa38xbpzFW
+yKdF3GC566qIHCG5p3IWwGo+xCFTKfj1rlytyed3hw2F13mwsvlP4YKUphBpzyk
clE2X1N6kwBc4NhXxaq2SltU68vRbj9o9O8SZtthFaceC4+ADLAPPfVXVZcUsEp0
yHyY9ydLCLZwQHXemgu1ZYnfGSktM4Hu0EUhIBnOjMA7pqfbP/soZANOXc3EPuEU
X4m+SyyeZ+HgPCTYptoyzLF6LKhHviQvL0Fqq0DPAP3+jt3EsqOS4MMQlsVnOBr8
CAkndaaW4dNQ55mgtOpN63YTPTmRKggFb0VNmsSTNjRdnZJED0QWD/9wIs3gT2As
2AwOSzzMukXiUylzr2nBNsPIiB9nSFPgabCPp84uV4dPxD/kY1A272zZtahseN7z
f3oOLJefADMFlH3uaKaXLItUaSX8MqoX5EuIF6lAZoqPH1bpELDm2Jxu1hOPAuwG
O4MzTnCs2RbbxFVxMt2ye0ia4kGCfRRbP1QSO1mLsZaoeFMn55B7tCtRSrTeDZ7l
GN9nYZFcsbPley7Vdkv1ETVDebk24btKqbgmepLanKAbtexwD5Q/dbkwdHXZlHMk
Whig4/CInJN0ljXJUMpehS6rAAdhXVd1pnA6BsdX7WrJeMAWTuJOLsxi2PmetZni
7g1j8oB5tP2zehbHKY6QRyTTw/KqePqQobXfut2dY7LsmcxpuSrib3Fhpoh0OkuT
e176PbpZ5EENMSuIZOEyAlw5Wx2vL1oJ2SsXAV0Rokmw0XU4tqtvrCHcR/VH4M+I
sV22bTZQSfAXVlSfqRqq6hF1UVoojg+ylQzDFwHrwpRu20YFrZYyEFmGkZOqRpXK
XDKZVD1Gbhd3Rt2qAogDyOCkwWrWio/c++jZlig8+DQMtTtfi5zsFQJQDYI5g0gA
uVChStCtSNY2h1B/65nDLFVseTW6dQJqLf9ZP58EuXRAlrwJ4rqYl34o801WjzEt
48T9IUFPuBGdNAwpj/aFNq9J0Zwwvoclyzd7rRHuDKcFOy5vnV6yny9BY0gnrvWa
y1d2X+eIn7EkfIUfZVtRCHavNxbc6MOfuos97ixO2nM1Nzo1RZUNNSCxyJ91tJdP
0r2OUdO2HmuZPDUhuoyWDnkVA8yS40NDj+h2OFt+GCj+FbyyOEHggirRp/8dm4zF
6qV+PtYQfEz5NLaRwN0dDULre4zICKfEi6rb89LW9ZYy6G90QL23MIDfhFtw3SF+
B15oAuKEdiUZItyGZUB0LrzuNCIZrvOvIDaTcewHimFMHqA9+WbE31OL0H6hnAQh
Diomrr/gWOGjjVr+kOqIi/SIFdyUW+ixlPjzmTPBncq1inzPJQKi8g+GK7CywscF
iAudkZS+v78svkrNWLlhucM6/3n78izmjaFOzvrLKYJ3eUT2nRG7MOQ3ovnsA6Nd
8/DKUhHVPazfVpPAQCxvD2D5FHlgW3HzOaxyXX/pV5bCZZ1pYXhM+SGKW5+90deR
7bO4YVcbZ+Q4me78WoJKm8i/jtbGWB4eq6yAm8+MEjtxSBSECjtpytx3/VRj+XVl
wDSkpWd/wEyy1dvEaXK7EZAOJJ/OoxFGd1mYgTiayE93Tolt/cDLT5awe8ZhjPnH
qAXoeHs/7dfYvefsu73V9aHop+/FsHdC8sYtbJUHzimhZN9DLGGb/v63ybIIhs9l
k+bH20Hs1fquEFm8kZ/y54FhsQW6TJmroFdxm9kzGo3AS0GZwhdBtpJqrBoIdSz1
P4hdH70jVymc+Fiz7ElSZW457cBDcciFF+M+qodv0niXyupN7AYWbf0DaQFCrKEM
fm85m0O1CqIsH0wXFx65gNs41IzQLi6NIgvg/PTjrVB587Bv5TZuTzRGjT+LtvT3
kS34HVl7LFcMMD6l3KQrN9rAfKfnvY92Fh3Y4VrmDbCMUweCxBgIPFracg5kBwW5
ESZgSVJRM8Qx8b2qk3mYK7l6n9ochiLho14ZAG/oXJCcC7yczJRDlTeMCtR9gBbe
P4O3NsEKmb8baJN21j8tkrdKA57zDLn6xUWEi07sQUcFWXBpPKptlK1DW3EiPtNU
SKTbCmTwk8PQG26R+k6u9cyP/6j1LxQDt1tARqb73bFFZKhOVAJ/II/toOFtlrUZ
ZBki5bNf5vl1NTkORCT/hhcAglGAWgkmDiYlEuDwiNCzMR4icK7DPaRvC6GuP9Wi
/EBmh4nEM9NYQgyDYDkm4oWl2G9W3ogt3jain9iCLVYKJ2ky0/yST8Z2tRo3MZu8
BzSGUhUZHEF3FuSKW2VXAId749MF5yZXJOrSyHDB1X6z56LH34dJDPeXjg6yIlfn
En5r3WFYxrgXGZUcF4mcpcUiCXEMUotnrX76/rb5nQirKLUqmr3SLVSxAhqqI7pR
yh3je9AOnFsRfng1pi75X4b8x0vBmtcy3V4/Hz0O7sBZS1lfcRBQm1/tKK5cREVi
LfKJYPYpZBziGo8D6oELZvTdMqTh7CkBTuvUdxdkohraSrXeqKg6Rrv/P+e+IyMJ
5KPyc+8Cx2h622tiq3seivGQxkm7NAOJHnAlu1PjaKcJ6a2S+phJTAM+zrF+PXuN
tiwu6eygRM+veEwSGzQZ7DiIlpn7uEMh7k5LB9SRtZQ7UQidzBfjjkHOocJkfkDY
GrTkN0tOsz8u9R2Za01AdASofo++KdEtZu6MUa6CUaRGZMjf+h14ZxAvDfEACrL+
rbw/S0/3Xac8IQuU239SQ+Nv5Nk4GjBLuTpwh0PMdYUgiU/HXMq88V8H1C24AVUK
X3yd8f6tBSp94PejAzk9ZVeBm21x6HLuDguUPzcF8PaD5XLusRD+ylBsZjT9QK9g
Kv48z4NYqio0RPvv/CIjKDCbwA7gLZH3TxtJwhOwO1ybXiQGVdFcKPXz+fNEj7o+
qq9nuXV6bZQYI/9MDnpVe8vI5z/8FSBszJcSOXtBXYmNpfn/e692WXI0FQhWSij5
ggvROHUZESA3+L7Q7fOUJPOjTWAe7LaFHZRAyj9tfVGX2wDTN48BYfDApJIBkbxJ
j/dg9Vl7pHDPHTfER8xgG09ivvgkpDqrP0CjWsIEMlV5HTOy3ICjFqI09LrlT7pI
M6a6ZRhxDdlhAm1qjxy/gtERbpqXtXQ7rvjITYro/pV/8zUKA/phht/2FqjTZw6k
SoAIjsuZXkE3eriGtH6ArNNeD2CgvXmF0wcstWuX5ATTsegoZ+nPK+w31W7nIyRP
WCZcMpGGQ4QBJAIG3UksAAplnGdrxrBqY0Q/O5G2sJTcLsiZ4FEUSFk9kejxReHX
lOu/unqVWsPHRy03n5fKeK7SzBq6NSxc/5bDCiQWcF7YEI/+jtAsGuc4Y5Zrps9B
bbedpqr7cBBTUmVxoIo0kybiVtX/bQ/ZY5WbzjVM5t/cU2dqKjCH4cnvOm1+heFE
iTkNelNyAev5B7VHD1apcIKThkmFao74Flk4sReF2G+uSuIF7iHt16UPqQJ2sQMy
QrjBLeHFo6++t2K8E5Jpf+eQZMKHuRQ56Fu24eXQxvI2ByIySpBmgnAACuxN8OwG
bNbgNWeyTSL76s4T9xAHjIQs57b3AtwMY6BeC+zmZ07QeION+MFmeuTGau1l2B8g
mi+/i7ajVR8hDMqYc38Pw6IuRpAps4N54uNyHlys8RBNAq38Vc+MtUG2Ka10AwJr
DrqQFVgvd3QzXRXzzJfiPOVMj8oyN9GSxaiw6WF/FjN+/r54BTRJiSNZ7F+7GuS3
5Doj2XTqpZr+idXjIwhdnDzyqoh7TPo1Nzs6McuDIthrf5oaV7hidHwcyS/XKcYY
kWfIiQzncDddeNEDdR+LZywuIJ4eB6FyYROrG4HmNfjD6yRjthFUQzpK+Q4g25VH
1TZUoY/aNi7HfZ/ajqW/Jub70sgThBB4W8aINOy73QbhXQJ2XGhD3OaBMICirUqr
An+h4Yn8EYvC2a9JrDcMWdo4vpoPQOXSpwqB0R3ZTys7adx3ZbMZR94daFdO0m49
Z6h6wgoOtgKL9g0Hp4yR2ZG31BY1RhEs3x8B2LcIhzB3/oDeeDqhYUQq3YqTCu1V
4qI6X2fu9JFA+6R2sBVr2M4rumQXMu6cujxfZSnlo18JTdUy5M/Ka5IjoQoe3EKt
fBTAA30MILr/HNWmnWVxdcA9FfdlDgo7IrE8HobQ6SXdgZLP1R+HCeluam9zo4rX
BNs4goSaw1oppRR99PUZePAfuC0rjT4DuUKjCebfL7Vx2eoLSE6JmA6JoduasdLH
p0btkVz+/sirhBL4wQBs43L4X18buO+WueI56ZKu/PvUrivam7vNImWaaSDLmpqb
6ZMkLkwgotMQUfHikd8AjCadDrhCzKt4EGxV7vTg9NmlaeEbZB+bALJA4/5yQV9A
15poU66XTbRXKAKDRcje6npsgREJTNRMIos2X67G7CE34mjXcYUnxbMuGHcI3/jB
mVSiWb35UBCNYI8zvHPryp0/CaYRjsWDJuRACQvd+e9oJ5YUVb50leF6iewRhc2l
Us5AvhtvAKbKtV68lHFrGlCU9elsinQKUxdDw++G+chUsIWR3jkEEN5yzydeXzwR
xNBlcC1ATF5lVtJYnxFoIsoO8xpd61gQTTdnYYjJhQbyZMmgKsGh5EXd0aZPo8w2
icy0mwP9Hk9LqS1Xg0EPnz4Dv6DhupX7YQ0jfUu8Q0kTnus3nvusPJA1+XurjHL9
7hcqIylh9fgfjvVGLlFvQuo6Pd8n5Ksuz5x3k9TvoX/EuvT3i0vtdwDEFGCKFldg
JjYdUjJ+8VOeFe/V9u5aW2KEv0yi0HppQKl41ia+xQw0ePe1NBWKULP+ZdWe2t3k
07/J3XsHA57kv25MrAdY3g8jTvhGRVZI+eJGWTNnB26w5MxuNd6ybcyZiYSjM6Ni
69cm6OdYRitOkrCUZ6Lqs4/jw376UOPEe8+2xpJ4+p4ao+vNfRn8I2PI17xnBc/7
k72hZT8Mi11yQfO4LwOLu+3LVCl1VDOu+Ssml9IVfqbEcpWzSu54w5UnSXZRCLn/
GN936SIalvmnBPM9fa38dH+zbfwIPQ6ciebMnPz1PtrsjnIU3OV3kf4Cn0y9c5zR
P+lLHRTh/7XB/6mk79Zwk2UHoEAamACXPYZK17VXab5tRGda8K+3gwAMcfZvC1fZ
JFLhO5BE3EQ3OTOaSfhnzyx0Ljz9pyVwZHzjTI+p9gGVYfl11ibrmyrz7uRfusQB
7RaJbR9t3CY1uL/Ynn41aTRyY422wkO5l3LmJNStfeUZrpHcQ/7Lc05G95RtBZl3
9hvQ+caB32XkMVEzWH40Pui8771PVkcXCEyRmPEWaQ5e9C2u7E6dTfLmfGYccYvI
KU9uSYfdaBGxzsuarWmp/5HEazfUeV5L5I801BO04lt+tuZWdeJCK4J9gRcx+ax5
KyRIUaydTq1MV0I2Pjf6ue74cLtvZD5Nv0jdsuX3QmscwtiCyVU4CzxtNUNNyTum
4tJKOwepwBZWA3lPL5E2cewVuuCesHmcrMO0wJRooCbYGjJ1Syu59cD5ct7ZOk59
8K3gDSniT5Z44TnRSQfZRmb8nKQg/NuIfDR+GQjpZqWxzMDdBAMtv2DfZtbIz/Qf
Tca6lXHyTaBwukwlvK35/tfB2gXbuc5Zrhj75rSsT9/ClgJnrdsIKqdBtsrhJwMn
G+lrUeqTm93Tz5ZpKiKdsK5lnZDDnGlI0XSR02iyk/tnqDlIeqCzHCBe+WD+oNJp
8Ay6VFwSZH9PgGtsceKIRw9EjvDvti67KntsfINWUBXtAgSsQ+TUZq6HfylyA96d
9wQk4JNtGVpA8Dhlq4mBC4hSX/Gq+Sw+bkI4fzO+eJw2OuiCz7D7ntyIqEa6Nm5Y
VSkMQ+tOMFOBp3Pd7pDFuai2Yitt6/g9JVQ7GHMx9yLfhzNyhzLTr8qGAPkxhIqQ
4dVTQLedYgJZiBbKbQmFAGmnQxIcuFBRz6RGrXbyIzCaTNebqBfgs9a9RWvXpVrn
C7SAaFwbf3XoECVa0eTPEQxlqa64VfnFK0ef0vzpczGX4iRr2fUCza06HlLLmaTA
h8GNw2rHTu2mQxhBfmkUn+JO5Ta7ls5x1E50ls5sNsX3lM+eQQ0egcrchX0HUWLq
ruHMkIf56NW7OQABDdyGMmQus+I+f+FUV/C8eedFLD/tYOjdUFigXdtXR61G41vV
cqUiXaZSwcz2p1+RCztXoeWPhrQ/3nxfyGya8PfKpdTOJjHPy4qKeg6NjBiRnn1F
BnK3LcexEcrrOG6gnd6MAquphv6EF4nyZxBISzi/ijKak5aPtkgsx0a30A4hn90D
u+7E8X8pJu0mAQ0WQUreHUHoLknwhRU1d5s7JSQMCjTUyLPkMYmIJT4p+RsSj+E4
DI4lhfJLXBggCcCUTEypb1H43dHiQ/l6H9yJ9fOgItzsyor4kVgRjuuaeV4Doukx
vcYH1zJscImCus83C7WEaJ7k7ttDJ/+iDq5onQYoKhAcgKQli+s9Jv/1D9b3umQp
zagY/eAqgnRcUALNyCKnICm5HDyLf6PNyCOrumRkZlnEm5bGJLUuH589ReqAS/KF
raJOoM2ekIYcYt2Oh3YkRJmCjJsErZAhof4a0XzfoCaifWwArTqSBCtdc1WhFvqD
6+memPOnAOgCLjCqrKup/cI9h5FHpPLvjqHbxLJxeSRADFI1b/Pq1OhDoLyZpuV2
KOqJTwwsROZTwzX/qIzMrZRfbIAV8HtKOQgrGPefW/RuOVF/HFWV5oMkuMzyYcsa
CSrgNCAlWTEgh/7xPv/0RfMB2Y6dYvU2a7fXms9F4YEW1Yi2HxBfKbdh6DdoMzs4
rPKfR03eBTS5Z1wW2QSmMJFw4igj50kck6Amifelyn2fnaS5Jl19VLVjcM7s/szr
M3TMuMSC/qsbyOdkz9ULnKe9YJAKL/tAhk+0ouu+nh+cOZsFEYByphk5b75zkmVI
7ZdLHQniB4IF11wsaNWQv/rPiqZzOhxAZdxqUidvkvEo6eYHzXQ/oc+Nh5JrzeXi
dbKVgTx5emPxftPqxD6N5G4m4y8Y4ZjI65pvbrtOH98qfhfhe4nKpcNaz+1qPjzS
AeDkiuaww0Te2CRCXhD9zpPdDC1LIaHJQfo3qrjIMbEun1UzBj50fVyaG0NRLZHD
0DKMnx81h2vparBfi2/NkQ3Z1YooUoJCZkSXyxEwIeaSuUprbNP6pkupKtL4TYH5
1r/V4RISw0hBv+a0SHEcl4ww0cn3QbbKisEP4BxFUwx3NoNfKjitiJ2v603LMTlC
EBJYDhraLfQi7OfInCY0B1mJ6vPY7FRZsBkVGJV6lcTYia8TJANi6dMUlzrLDbwh
lxfJcS2HDGnZhNZjBlO5cNAeqkhOVqLyEdbkADUfF7+tWOJYMRMlerAOtMj7YOZP
Un3c49ldntc0H80t+D/OCYGiWncUxAoI+PYvxVy3P2M0T7ZBJhX2TWHiFM2K6tsp
6EQUZoIM8l1hzPGT2p4NLetnAadKM8GbXWJ+WRdJ5cBqR08yvK3o8n94+QtjwgQ5
SLHkj9IhVSBe8kc834FSobabHTrlJjkBne7djtfHKn1WZLSkAzTQ3j4U6eze2khN
9seI4Ww/Mkr3BAmgaDhGXfCQV43axCFVQq2Ptg0FgJxONXbFn31WSfB5rPZrDLYv
UPeCr7So5waqt0xPs+4UU/ecOGMKfr9HqJTHdJFfZdf5Q5RwTYQPTVFXK/BFNBTw
MGMkdOnMxg8i7/qUFLChI7oO6pagJAGjVd9o1xo2UtgG/WazMKXycR/JOXNs62A8
uaDoGFqis8Qs+/3guYVaU3Rk4VZhh5DVGQ0ObKPK8wY5wO3+Ck2AawwvkOhHQ/xR
oZ5kF8ZXhFTX4dj1Spk+iN/ejtmZGcDzFH5i03NvC+jnC2gYLIA9IpzD2FEsf9J3
GiidJdpPdYv2XatoKrO1qNsMJWEJSNszPuAHU8Lof359pmKGuhYqDnBYE/dYgojK
jGI3fZQpdhz/H+ZK0I04Fbrs3O3rWEzSG6EcT/+jY7ztqmDpYMadVIg7Z/gD1ZtQ
zC76OXH/ejcJtZYQ2bH//mogE01LVhkvIRpSUoEewn6lAzMVo++YONPAwc/5GBmq
jV+niyZFl05usvrNNQU+RAhSe3RumR3fKfEgkVA6XOIsZ+goN+FcTPKtWCMFmKKi
/HwqWW+RIL2soPMx1/Dkv718sOfd/1VfWX0D9c72ZYNxsl1epH6uq7vqaS96cYG1
CxtTVrDA2m72z65MHHnMSt/yESbBxScMj3cZ5gbJKrzuLivdMQshpnYdCsbWzjap
5+jMNfGmcoq1dy+o5q8bhy6DcWNpRpcnGigEdYWqasCSJSlP1oZTHmePpAnLBPkQ
JApcff5scaVb88mcYPU7yMzaB9zp9EAp5r+AEP46cm3zS3dhPdTBKJr2nTlwlqqL
i8BisGgaGQV5N8BXnCCaKbYUv8NOXqeKbNLgjBTS8wKOtD7e5KYGlJ1krRC6TC5K
lcl8FeNwCMG1FSfa2pAfow2Ejw951V7pCpuwpR3aNWJwtYc7949IyPCRVg61GXO+
cZNj4bl6swa4zwKAE9r2HRm5AKVLkVoh94/muLcQrTVtoOlpiqy1HTrp8g8volx+
cgEgzJB6FvCCvUdH9i+v4+JU6N3vp6M+4+egZ5axESp6LsKAC7I8FFYC8Nu6ahSO
f6z09ImsvVFUYWVIB5ASvMJP0bQYg8Pey7lwCtBoZFMO1wOUL4ZnSY89er9b2L8v
gNc1ooY9ffbsmm5FDfUu6r2SLylzFSPwv/s072ayCLn2vbd/ExSNugcQse2k24rI
XbqT3873PhFcN10pdNeCLaEmUebv+DC4whVFnkMQtCJK1clz+Lt9WMkgxGkDDD49
HFd9k7xlYlPizqriAZoFg6dbvfRIxsr298YqiSVv7Pi1buKg9Rmnwvu8hEUiE6x7
kQ5xbOR7jG8eF12Tu4pooUODFi7hGQSrUP0VWS1ccxqPDypg2Bmur0ITVtnFfSxC
kVliv02h1IE4bGsYKKToHJ9ajbAZ9DlVmrsxdBY+sZdUBG/Q1hSBneRVZvXB9cli
C9sv8iJJFTbw/ainYymAEvm7816WbptYokqiFTcIjtuGx5WN5csS+kJd/ZiiQbxc
7d/8lv12W4iVaQsRAmJGqC5jTOrqXaRNxfSPIssjZvU+p9bCGXVtoRnZe1c22rYK
ZBHh433cz4qnXUkF1nu/QaIBnHpNPwxYVv1iMIiuzruCYaBzPcG+Piv+rDmHYs5K
ppLHgFyOXfUFND5QLEfJfx6tmyX5hNSzXxTSEH4gKHuZ1wzqtWuOQr1PUQORAVvM
4EGhPGgWMrxndLE2Cam6AcR6zx3LJWsNH9vdvgvgkRwo/ucCMMIgyiSFi5nXlPDz
5R1X7edaB8muMZ3FsO36w9gfBkQaczWUWGPoZOtS/I4RKiDI7Euk1H6ubXfSL3sJ
CsoLMTRVOteUh+3g9DDSmGNtE/Uf1kL5eeTUzaPuT/jz45CQEfFiwdyOE+AJTgc1
e8fYM2zf239x2tPF1C9tdlvcMVKkFNpAPkeSRSgMD/ciska/J1XpqYE1ulT8BlLu
AuicWChhlrj2bXP9av/2MiRZLHrJJSf0HGcbYy4FBbXfhZ8UY+T2p5/njXxpIb2z
y+eydOOCNIzEmt+5WJw2Kcgs+IycanSJW1NfslDUU6Z13+mGRRHS5xCXWmOvJNvu
v8Mq/i4z1ipt72xTKgbTijGTL2SDrv0dIIfMhP54n+U6SvuH34ZjxBfuEVbMxC/a
S3swaAt2RwSvJuyPJCYsP7cC2v+zoC/04MHDDL3GtS3NHiQ9/gqhhlL4S087kkbq
NXZVBq+gWClzCeTlIyJANVaKVFyM9pY/JC3nLIhd4wFAw9KZrRlGk/RoWdjnc4r2
kQj7zCE0sqqHkwIxoUvHu2jTTwkXNIUmcAfmATph3RqMC+/jSODzRjEIGtTmJa9I
8MyPHrls3RCqaRCMsI0Jgab3mcbGDbqPEp3NTYN7dtyjDHjLKKqJ0rxrxeAx7u4Y
jEOuIYPU7stXHCACgyCkPETeE60y75E5pzTcbNoITFoM4YUTGmDblrh2a81qvZyp
q/zfhGVsJV5JUBm4OQRLcf/LW6cywRq6CXPZwpNt3LROf9HOq70tFvGoYiBM9DHh
XR3yNEDW2OWmIgblxdqhMTEKfXFHYpN+n25kr3Fbg/Fn0rL07iGCqtAh0WFb94R0
k3tqmO8buahiE+/x1X6OffWNTkU+Apy9LxOzKA9uly9Zdqko6C1HxtJU3NZNcEJ8
vaSQ+F69pHvLA4XZpqmOXZ+VsnRYv8WWtE8I5OflAClU/ARW5g0SR3w3CYt/tBAE
Bl8PC3U7xmVBP81qK/LgFCyFj0nvAhNUEXIfZbpzrlNB30JnAzYJzcpIW6dP/Q9n
bACxDgrXm+BefomMvLXTq1ptSgjfoKuM3Z1HvoIehtrlrFBpc+nOIsmgg8b9VApu
qM/QQTTtNvSZnvk8UBDWxbUI/Q/3+TfRUxGMoCb5Hm/WvhWMG3/IZRfklSvC3eEl
keNUXGcRZpvTRLnxUU0BmFP/lsval/r7HZz/6YdfMkdi+wmct1b1IeP98TDKUGc2
skq7bZaFbEltR/Yn1djeZ5sCpo184Sy+0/bnMzhFfUnC5o7brASWff059ThGTiRQ
fXYjKjUULfi1X6ve2aWODKDHkuXkq8GYwc0LvQkTjsC7I8IwKbo1qiJ5Vgwgv5cF
Qsh07WLsXK81TF1krkiAuwGGRa0B8+IS0AFUsWYKs3G+snVHrWkGdJ3pP0m8xQk6
OJnIBrvV7DOjTe7N0z29kf6+gtnrq35awLoMnBW0G7vTwo0PCMh8t0VjxCf5mLWA
eKY6murEcQYYkjVQb99EhfA5t4tKmWtehKZrB3zLdFtosFTwWJUGW4CfiAsevUrJ
tVaKzYm0QJYV48Uim4LWN1RHprRnoGapUcMoZZp9ek9SvIgfTJkOIi/1XqdFAyAH
nUg36VifTEW+reuyqZ0sjXFhe2lJS2fHYcP5GBKkuKdfW7Equkmzj2H9Ba9CukIR
g1gEL04y6UnxoMD9mgNfYwyBswBaVAq4mEh1TXG1B5pg/KeapE6xzwMp0mS82CIy
V5PnPpJy1y6apjGIwLsY0v08657LNIIjmmSHu/LMxu9hJ54/hiYjp88D2zBi8uTf
WkFExKSkExV9hmi7goms9R2McpEU1xAq+w6OrwQBwyjAkDyRJaAQWdW/4eud+cwY
Npf9aWhahIGmILSkoDIbwL7i2SKgamQ8ZR1aPZschumtUoYoxCU46138MpAPD1oS
rQmsr4L0P/D/ZLn/msGMw1E/zWXvb1+u647K7IYIm7979h5ce8OUuZ8Ij+7/A05N
6iAgb7OwkdeQQvEQDSuFSFBDGitnTlfn7jL/mKuW3J9BcVmUQsMsZ1TN/Zi8M3TT
nmjL5RjnfZ5PYLaddxFxr7flAscB6jQf9w+nCp2mBtdoxiwiv2/ZQDxGvbtjj5TA
ccmgC6U3oDI9IXC3sEvaQ4lN4KSi6iNcJzusc/b7eWRNnJ2bBznQ0bVtMbvjISQL
+m2QIqax+iVN8W67WaWuOS4CO2I3LdKp6Gtg3MUaf0q/IsrEj/VuD+3Ia/tQIasa
ivM3vrOZt3fRK88xdCA8/znk7DxsI24i8wzBu1gTVUZqP1oK5t3TNGUMdatgXKsk
YQWtWqyBCeE8u+BSPJw4ZkByKZppPQrtjiHAIVNkEUlgvujlA0gVnX6GFgt9a79X
EjOZsdOd2mf0JRQGlKU2xP2ySiCCu+MD89gp2mSh7KWMZFh04rY2d1MRYhX82VGc
iBrvv7YYjT0EObtdZsVrLq5fDWVBCocGg0tCrRAIdWLawA/xcdhCGbGi0Cpe8/FV
DT3pyD26rB39/MLM9xSeCKzmEEIV7ukxN5jpfo1BeL7y05828EaEdwyNEFf+LIbc
fj6AZEYuf7XOT2364jCutuFqIkvqiaAxeBR37MlD3fLwWV8WRRH7DWsUsUGhPn2c
tmtxMwj8sW6Vj6OSfYiTfpY9rYB2wpEVWMoMkWjwlWnt7XDBikitHoN9sCCfnCHP
VQv0pt4kNAgrbmaCM4ZQEU6lStDrYbD4VMFNGHQ2jOcGwvdHMMXgAMXUl876kTZz
uBFDOPPI7RH3IwJGa5EXrCSRm8SL75sp95YWYm9/xzSfYfgcsqDZcCP+mIVnsIka
FPr7N6hUHCit2aQ8VcDRvX3yHYD+M1l6emBKc0sJTLrTGu40p5TgO5ZA5RVc7zZA
cwY/5hvVUwVJZoSJYg/vMmNJdQmFcSsjmYdEymkJ9B1ft6pNeQMhrUn7coF5nSXX
pHXM0HkjFxofpJhnGBsT3mzQrFUs3qdzVfG6D5BclkHKx7U8wZP0fCExpem/tEkY
+fjF/lJW1zvjxRzbVPXOKw1ZaYHTpGyZdB5VJTlHQS6R1pB3DAoYhiG8Kau6bBW5
FbwQxFVpDia+og8RosVV/1kynXuXSX70Z8piQcUUq8Cuxl+EnYiSzw1zlaQcMpUV
vgWmTH+r3TOYyR17OiapFa1O4oKnI4Tv1A1f/XH1r6HFNbE+8nJy7FirTr8F8SsE
A4mWURC6IArlcKWdGE8UnSjO0uQ5s07a2y7K4DYS6rzpeeeKbjnbFoa/O1CLpstq
cL241e6Ms/HCC8WHHeuVNXmNTBkegNg5FDjms1yttuvUfhGm1fCImK/KT31Mbeeb
l86KmJtFfyKJMQl006C+Q/wCeNgo7FHUInm1bt1o8wHlczwSwOpR1f8fyIc6CKFb
O+9yINhOnVorilhnTS17sn1fGTiwKKnVIq32Y2aVvgRz1HxfCn69p+wLLaa2KUvK
NEWMG/bQEhhA2gb0ZtqFNi8fObt3IG2vo4cW1nhShLro8mmT8N9Y7rj0fFZhmwa1
SNHW35PX4USFscXkMJ9Tozn1yn8ZBzK+9c+AZpFcCZ93m3/Hdqg7pNTBxAMqyyUI
hbSlZ2DptuhQMIKZG6jf779mUzLyl3PxzP4mdJlnNyz+BRDs4EcPR3MVPq7JLmao
J8L1DnWMWNyzYD2eC7V82sRTA2yLMyFA1IdSmaV4R+7lpgJWtKEfsvFbaeCgG5x3
NxQ0OgM/5VEFBPyBqtr82M+izHjRsG/h7Adqjqwap/0LFlFBRdisT9Qv402BberF
nk8nVbtIqeXsx4L1NvWbAaMHQiCwhsiAh4xQyRNH18CQ7dwzDHHBXhx3E9DRJx50
lrVK/BCiXuLiUzmmqnlbdDeHhYxISo2jSYiU8GDdZZ1LM0IqT28/5UQFb1+MqKzf
h/nwYLWAzhrlF1exx3unLIRw2k/HGjVWElrrdNlmFN/R37nOXNnJKhSW1ELCuLU+
5OCmzn//v5jNBrBPCpCjEgIVoGS6s9xsVO2x8ePsMI5rpmuLsNRi0DhEUqfem4UC
/iFuYfEEG8KsWyAos6KriqaXPJNrQ5k1vJNiEiu5Vk4t7XQhI1luGdqD/5DDdUj5
FWajsIzSyK37uUa3S90yYv5dr4Wx2CQKvxqsiEh1ipbh2tbU5/rUlot5XDF9H8pQ
wvivhfEcrq55RLGU5Gc45uopOBbTI73yxJ/fCVDQsWS4z6vOK4opTAzI/qv8iSb6
xf8uvEEWW3Xa5DgAq9C5fGdM0HOIHwlZJ+r0iKr4w6DaDpm8bSHmHejnST7bL73y
UtKwjdw+vlqhyiNlG9dX4NCF0S+D+7k7G2Fcf2llxKkaBE49A7TUOy4XDGLcCKmH
ijUpNfJv8H5jasrkjuQu/A1e72qGEwZv/iMqzJY7RPPkxdKnEr+QWgiIkXaOb+j1
HZRx319P8/WzTRuZ/MwUN6hOJg7vjGU7kumoGkJ1SYICilepUR7tX6UWudV/93By
pvoKofnCIuoeGL7/L7aAgEsncyOp2zl26FuKR20CeLvD9omV+PU6qPYVZ69CMq4m
zkm5OE0pKaDBTlEnyBwn4GauLLz35rcZ/RuJJEZnO/toX2akmIGuWxrTX9xhequD
eP6gImZUF2E1p/BmrWx8GcffIT9PGQDww8zKiURVofMVawrNSGmAHF5vvWLROIvO
bBLt0TyjJJfbWrIzcwrxFWumfKDkLlU8WJgR4UWgJUzpihGSqktIGKQkKTBE+Rhh
WXnljMVZQVGqUsIJnCWMH1qXl3t+Wi+OX7K3xJO1Z4gCtrM5dBfXR3QkR5IKd40E
QQrmQ5jcgg1EYqpOFc3u3bd/eDPMk3upWQS3UO9tHPp/UGSwFSb8restqCanzeZd
j10w/wFk/bzXkEqIRcToKNiYQTFNTXfRBmay1lycd48d3h0clpTDzfI3bU+DGHp8
Qh5i6Mr2aJJP0RxMgugQJySw2pjc6htxD6bDcsCxVgzWFBQCVbnZbD7TAMP1HeUk
b9hvp96Rpn4M93NIO7J69K0gfZRK+yNtci+7Te1M4nMEwECpRYdrhhi2Dm6z8Y6Y
aG2XpdaP6A6X83jmKxW/vSPhT9GV4h9mAHLUM5YpFSEPfpthPsqdYw3uAnEVbStC
WZl1bVjuChw12QQHtGt3s+ugH14nF+oXKYAcd2y2o7tq4Lhqm7WrebXqTMJ1nHBz
y5pgEX+cQAU0ltKsA6y3Aqsr+TviZtBkj3CHuh1ndON95FQaKrwYsgL0Pf2xeT6P
L6nZKZhuePYkQu2ItH/JlPVrvjryrYR1i2w0EuZ1yT3mdkqg2KhpNjN1UWu4CXE5
iHmCVRqH8ks4Jocif31wHEeVvJJDtVmDtB2J/U3sZNdWz2j6XnUSyZGUUopO6B5a
15ujaiyWwfuJf3yJ/icYUawkGt3QUVA+HblGwL1xxlMChmdzDLTW9PN2eiUZfeU7
Y3aMEra7Pd+4RPRjl+l4cdN2N+R+PnRljBmmAo7+skfQpaW7NkpgHUW8KEud6ZPv
453ZzeypC3Zxa8RBSsIddPagEpILjZbmgTMnaAANR0Tv3sohBorcgmvRWKeUMSQ4
iISsKooQ/kXF2jtN2jdFSErPKTwVgq6dBb77+YmZIPwAluQfQgZmXQjXyqZjkV89
BpK2HTPJRjHs9iYxG0sm0xcxoWci+1vkHBDxvkPxz7fiqsHn5e6vYl22qvzP0+7b
b2uk1RgeN0rUZN77m9srAZluuht/5Xh+gqCI3GkC2onoTQYQ9KzeQbNHZKkt/1mj
buSbyQIBhdWmfmvgpnculdEQ7aMt3xr7YTvS8mu4AYLycsLkjvgW58QeGladhSH9
F1MJb18Tn7co+xbH/8UhDJCv6beZ0sZmV3YdNoQLQyElsgejR33LbX1X6wSUHThs
eieteu16QEBPssWHQszuxjdC16WR6i8BP8dYikUrD/vd9vkS9CtjNoJ7RK4V4k34
BxrYpPhlhWE61aq/M+ClFOofcAnu4yeWeusFSpntyKbGQ1IiP26uRXS7vJEIuoT8
z/jxwSRSQglS/dVdfUfhxbo0prOMq0+l+X7E88mFv9ZZfIcjCBqpG9FvmFQrXKK7
4vT6FeJMuMrvcjLe0Dxhy0n1MRHSLJN2I7DaRQR/WIba9GpkrxJM8VkGE3XzbOjX
4Wyu257p8+opW7FbW/IPg5iDcJcjLj1pPTfqOxgqNcZwfhaB9PCfAx0DJjLEeo6/
JHW73Orqbr4LIZ02roUkKgyWnmZigfWfPS5FviBQND84s/F0b+whJPfiPAaxN0sQ
n0Do7FIxyLwC556fzptroXGHdp+h05CAJ3lZiQHCQMgHMb0MEvkXgch9ATIhG86i
3qQ3yEN06JmjgAkr1z5Wex1Hr4SvL1K4vxMVnv9KT79OjYjsMNjrH6IvtLNHqCEk
imZXH8DaLpdjeo1dFknCFE1ncPRmf5q23l3mu0M+jmgFTDgAGhdndfazcmCArDzp
BXfciVnP3cSSkhlBiJXgWm64JbTXy1Zt3Od0TN7r/p7LWsHiCFicQBq+IcQm1+f2
Tg6etafdkls4hATLhy8S5XjLXrf/q0KPQTJsuvfW+sCYfoiuCwobgQrH+Wpmu8YX
7tN7L7uSzmqu8pz/OuAHmI2yoSraRC39p+/7z8Kj09vMwy7GzadS5y0GPs5rshjk
TPpzgcI2NIQ33QAClLiiLdGDqpqJ1Rr77oZ1k48vu1S3swd+ZHd/xPUjXKbPV2f2
wvgjKuSedv6BIOdMxuSWIjWUFOoDSyrlYh7hTRJsFENzr2n6xfNcf8elpgWV841a
/cap0x3tOJyePjcwFXF8fL9My0J9o7v27IavO9sbW07Rt/2zETGD5LJvWtO7WhvI
jlTcgdBBLhy4GPGDhgaHIePbmrzn+vEwZXNIuRYZMKfQwI8OqdiTWDh7/BMhZ4yk
C7LiBwcufLbxb4yCr0zvb2H/R1gT0Js0TB6Uq9ZnVr4wPg4dLCq//3ZkvK/a4eE0
bkdvE4RjlcfFMkgvecejrthJK+TsE+qKTInWFymJhQbk7rg1jVgkA+43ni6ohUrp
UCcgmfTxjXy+ixHCGk6IV7+ABSICrHSDiNznEXybLFp3hbrbII0GCmdXmtOGc5e6
poAHK9MRVAKKpIYPGcR66Jfj0JWc93aX1nis1Le3/0e1pXQDx5p7rcf793tWZZw0
yGlDMc2kB3HYs84N53fNijdzjcJS+W+mZXDcJ5raXGKp2hcJsme6y6VzfOE0lmY9
J06KkUgrnQP8Shmj8obUPuJRGqjh2/Eabprer2znj48NXBFNDmKMlLVl80kG2wrZ
5HJMQoMXEUODHZOF5D6Cnvj26web/OFAL4uugAbwdAhktS6AyWQJkJbHjSviApo6
663VTDe0q8RLzevcZXDiLt2m8ss9oe0u6/cXF8Y+3bvKHqIjW8y1S0dgqcKFZZD9
euEyzEICTRYttqZMSZU4hZB0iI7s+SG7hqMWAZ9TWe1EWuy+jNMVvLvRkaqoZye0
FSoXLmLCaANwVwinADdLqBEqHHrjVZKVu24Xt8pTdCVYG11sDttZfVjOoCi3Jbm5
k3VPou2tvxUUpSo1jIrk3ec3ZKa5O7M6N8H0iXMa1vDxEgPukc9HmbL/wUzorZx2
1+i2GUL6NNDwHzMA27G6JKNXGwD0mK+G/7Thu1qv2qtXeQ319DA6MnlD24K0KRUx
sfRicmJ+8w7PqQ6MftCj/Y/+Yy18AnAYmBh05zb7DVHXzEBWG7vNYCaUmvJt1n/B
lVXVrxuV5EDdWF17XySO1Uzk4hnz0DLZtIzPqpr1bjytdEaBeIUlWTga0zZCh3nM
2hR4LxG/0am2ud0Z1FtEZcq/0xaz49/W7OmWIxImiOULtuHWEHCUNBJFqpuMunOi
eSzINo1HvIwFpjuJBPEWr2gqdtknqmIYed2ulT4kpWL0UJy25vRDiyXDksvNGfXu
E2gm0/Y3dmf2Z74J/neX2i4xb3sNIb9WBvB4eUoW8nGshocaTNSu54+GCn1DP5bz
hJu9eMEdWEM5m34KrP+I4sGvPh4bbonC4NlsgpaRPyGxcWDvw2iPvHu00T1mEfTR
TOrA/pe6bPAmMCMlBHFEapW/yG/UEk1L/gb5KfLkw5W8kVWhjhrkoUFxBZPb8lQb
r5IUvamF0hYbczgMUNn3wozqoAxr/SxS4trMgUcjr7cysZEAJKHBmrdaZ6jAeqYI
FQAELRUvufUiTV0oKC/NEQs8LwnzZBqr3QgTQRweh3ArYDlVApWnVIqRUUn2RrBs
3o3o3uX+mxvZ/2WpzrRWfprKXd2SRvbaiasinJNB5XkN4NujVvgFt+rh/lBH7ehN
w57Z+9a3ogi9isqEjOXLRb0sGtzXe+dNL5jO9FQwDzsfpmeHjXtj0M7jQG2hdNgY
E+m9uBsMV005AoNm6yO4b301xWEKAkCPHhgUZrmm/fSXiKy1DjnRSBfs+Htm1ZxF
aeLTBqUoh2bSaknQVzsr++gwFGKMVp2klDP1or9pMCyhX/IozuOEia+1B50s4zNq
5qzsDXLpqwmFmg2ug9fozIBioWBL82Vp3Q13EjABRqwh9HEAJmN6/cSfwKcz+JWF
xi0aSPc6Am0s/QTsZbi4RhgX6ZgSql5MmfDYplvi3ssWDPb90tt3sDbAxTWU7fy0
XYdq+6FAt54xbNhJUNB1qh2bxf0Pi1WF7rq4ymqbvBKp7T4SZTcLcHBE/SL+8eCY
eRldckQI5iCEV3ccFvBlMD5kJzEL1zs28E/GewxbYH9GvSuch/hZ5EC1xSa2187l
EDuxQwpsyoZlc7t02Jyf5bhQ2GKQJm95/wSVBFpoKnZ80PvUiUrW4E0A5MXJ0zzF
6EvqsSoswp7x5n4UvCB6hrfhTc6CGNmSFghr07P8A0b3fqVm2MhYfRHFLUS+jDgi
r0mdz7W5tS5gi+cwwLl8Eg9aWo9Zz1fTPojrfbrGL9ExoXWXaZUSNwqTiS6ZmRg4
MkLbHFVc17vlLad25F//wO3+Dwg8ROMSkduY0w3zS2cDjGWgDpgxH1oeW3JoG2vG
JDAIYO35GmQJsCTtv/gjKLkvULf8T3fbnab9x4tj+9OxCAB6ZqgZYQ+KihbRfw5A
pyNkvB9ovHM99wV2lmv2pnqLr/lRYJCff3RnsHxauV7klKrkKTNbhgKEOElnf/M6
pVVZvPIFJbXm/idDf7UInh1c2AUeU8blQkRGFthOzIR9nsWYlhQEnI463Ye/wf+K
34CAbYee+W8xg5I4+QwaNlf3Txjy6YasxGugREEmg8UVnTA/4sywYDOtjBR7fmFe
yImL6vQufT8ISXpLhlCIT4T9xcS3lwJZ+JzEP8yrp7H0KADaVj7+ccqIlZY7KMkR
02zYNOV9/72OxMx4yCURth805m5mOlSzCqrvQBktiQ0xHM3f0dfIhnxZCFwUK2Eu
0hP5r7pT8kKaEuggKjAHotpazqbCEwrhPz6hxkoZEEG4uAckkp6PTFu+2/nrI7vy
q5UJ+aWq2J8s3fT6VI4117D8i8K/p7dTBQ9HsbmUySKPZQ/F0a9/Hv0OD20QHOxe
EnAr2YPd9TRArlOlZYbSoRLtThcgBrhqDAJlgBaEiq3wBz7R8KDOc3GHbx2yrX1t
ItX5D2YprYabPj/K8PGw2zVB0VHtF35EkBJH8glY4+dwo5y4XT37QUtQRmeuw5wd
TiAXtpfgqlAooOfrGmYe0SLMTOfr8JUf1mjzR+A7nQj05ddayM4x3IBdIGfkkAUT
yxx+xvm8yHLNG+QGomOeWNvZID6NT5oaNyGYdK4iS4Bz0iv6EDGBrJvuSXm3+Y1d
tRowM7yEk5J+B0loOB5h36wFZmIH0JONf7au8Q5MAx/1lQBpTCBRFJvZ07ca1vli
381drjcPOl8t6QeC2A39wahl0X7vXgvAFwOoRUFvYc6BQB6X0cfl+GKsEKUXl9c4
usCHhNqnAQ1FJBhPNclkWxxaHM/OEJ32Rwqfp8GBZXlkYUwqHqTdTilePdSdataB
JgloKzNf0bItUIri3+oQPNd2130s/7nfTPFtz+/W9RBx7Pjg6sUO4MrBaPD3NGRC
vkMETCfI1MupjnxQhHoBYVkopt7bgWBp9VzL18nqTy9WPwZZ1AQ9mSTc4ydAC4YJ
DG4QrmBN/nyHef2TmsTbUgsRFfEE1Mbb9R21o/Xn01QCYgUS6qk2Jy8G9zfk5Hbs
rsFaKXzC/VmuZJicuNFHm04DhXXFMIrAoD1w9Mm3zfhzcbuBa5ZPmttR9iNqf84A
7b5pd8wpgGr5mqGv59S9jgpcYjgcfeOeLK70dsHK0B5VKFrPH2xz3i09bktmq+BF
adqCz3ovYKN8p3fcxyPL+DnsxlATOYkGtTDfZxoRP3b0BG1Zh+8PuYszdz6luBEl
4ZJjj32LEFyzUEJNz35s+5S+QKn4IcFuTq6qpBxsCY/PY5KDEXAlZ9RV5QsxQ0+3
txXLtFHPCsmB0U+AyRh2Vw3TpIZBS7rGQ10kVpPNKIwGOHSJAOiOnlo7RoyMm9Uy
Z0IBI6hovzshVEP1bduZlGNFhMU30WWzx7+Q7Z6eXnETZRYiF1KV7yJULNaCJFqR
0swQbi2kzJrvB53z/hNE635sHXa5zhX6ynsx4KomlwLKalgPz4mDFoXxXQYw21LX
HAgJs0xgCbN8m6pzZsCVaOeJBuEk5qbQdMHRv+dmPuyPgm9OYG+TqV+6z4GFjBh+
olMqWivLM8p4V9GOAffDz++YzoK3QpqvkgQAycT0Acrkcewkm8grDhhxThRGuLVp
AoXA6PfzmyTOkjUjxjRv8i+PXVcakDsRqbGQ9KFRvxQ1pCWI4hPPGxKSjwjT4XO2
cn3C0akp+Od9OXU/NBAebxwy+YnccUA4mn+v0iBxz6pM76SKRT+ANoN2HWHV2PTL
lsAMHyH9qihs+mN2L1n/NQc8/u9evtswuhCINmloOJaRForlGxQXgZ1VbExNNmDS
iXdpf+TcRvnYubwqN0hZX8kRi2NTPIdyR88H88Fv3Y7SWYVDh3yfF3En8NlGRZzN
DtAUR1cfVD3/rwW/InnhhJXeFgI8dkKGS5IhEgXB4i7jdX9g6hRKv2i5dGJeYL2a
cJ7baIZAF+Kl2aWo4gFxwdxqwaFI4F/KhyZKPTxdmxgTaRPxhJ8kjr5i8VJCb2lA
mXR10//mD5OneJdVeBSLQYLx6PotJl3FULFYGZNiLyXz+QaTlyWjjxGpbbOgKrAt
fVFsY9JM19c2rpB6zgr89V3yjenIV9lDgOsBHUBGrD9EreuS+3P/hRQmlySQO+mW
7P0Fb79O5Km3L0+7JZa6LkfXXVvpRoOTeBl63g3r9oLFQEnjmk/nOJ4UBxAi21og
pIkotDKX+37d4z3uY19ifhNTq9WeEBt2snplmP5r66WepLfaKlXmrq85YDJ/ahYh
D+DBC3Bh2U9Y62ag/e1mVdn5TXSa5fhUaX0D/zHRbqBRb/XsBCvTmdCdbwgQZXHS
hduZUEN78B8MlrHS5bOrJKCFO06ha03mtSG7+28Fb1ht7ksMN1wKcxiVoqq4AeEy
0OcVLRXaHNZspAPnUdHRelweC5ijCEKH10aUr0DcMUD6ep7ffwFUFwuOaFZIC4TR
GufwOGHpAp7nCxDFEbOI8/S0rsf81pmGjsF2CFKQYQ9XofYBL83CShD4EljvSLDa
Iknz28y65k7zoeJTnE0ttGA+nTaimM3CvJRl0JreOJg7CInrB5oeSiF6WeIPpKV4
W3MWmxTujDdb7i/RRqRc/s15evUxajuXLki5mLTio9KN/z6IUJ1OvW6G14hUuEwn
X7SdoPgq/g0m/zjKUndT3vpqVN2bsTR4BcjTWPELcPqvxEr+FOKjeXcQ0rsF5yW9
zoG98fPElZcPThoKbNZtbmxLUQprt9RsdmedhCU3tZ/lG/DogGq44hh8t/Wwq26M
G4lXwL8CswQZWcbRCIr4/cTmuHbYitBRCN+VW4xvi5lkFkZU/LjXPFBIcLeIbV7x
/lBdrffIa5ZBwardUkfu36S3QE5XvKHFRxIi5o4ojnZshBvB8TR5F7pxLSwW38LY
VqwyU2t+ZXxkAvUAecgOf+oqWSdvoKNMel1Ym2s17YAl10S7GTjKUCiL13hw54Ed
WGY78Fp+jNBHwwIMSy4PmgaWWmka7THdVAtyCdQXDi9RLSyEDfV0wo1UUpP3JZo6
MMpvFndhjFm2iMLirEYDQtC3Q/eAy/5CAF0U2ESczcoLlyKAod8RH6ti+fx9FLcG
8KIz1Nj6Cjb2faezJ9L/CFTIdQZjwLYRr9nF5bXpkjilRjCg23l6sEOCP0R0CwIz
6CnAXjuFiIvpBqS6gcPhUirb6bb7AIwxnz4XhJo42rvZKvfvU4d7q0HrHn5SlpNG
Xy51RP01lKy6aJ6zeRdJMzNrKmL80f5HaC1XCB9slHg5oU8upBcg5glZwt8b+Kt8
nvsFeRiJaNoT/k7lz0b38DJt5HzRvFMeE9N8wHp4gq4ZU/f+TLo/Ih/CBf3YxAQz
dwDOw/MNaf2cSySfM/qs1FCzqMF1NVTWWvt34sD89UjD+AsgXj76pqwI9RVdd8CU
SDwfDDlROQBadIZJl5wRLisnZvSBRtrtBPTJpOQc1uBny3QKu+NVugMzxD4IyLRp
MUGMgNmXZgCpQVptoxzztABoiC58ZqbZx0HXFXQCC6c1gACXbpJFMTqjtBvV+++7
TXSXS0B7Ir/j+MGclEdcC9vQSNNsRDIpoovPqlsSHQgG0fj13a8dAgLCIM+3qGvV
i1/zvdO7KX4Jv4ZVhaAb4YLN7QV14zWf0m2929/Z0fCa9D5NvrxRwdWYOUlfG/Vh
8kp4smFv29Yv5S8yprdHQzleIPjcsU7Vh8vxLJVpX52bCpPLOvpN6EC2v5240NsW
51rMPAU0UhE0Re5LNODY4DEd1n4ikYCg5Y4LzV+zVtdgLMBXmqbEzEZ9IdahLSxP
RX3e9XEN03ype5f1UE7mSVvKdpK+z+JciQDTU1y59FhMQ6cO3mM0RHk3d1tmzp84
tRFSxw27Nk7PSitMevuE4brbrZbPk0H0PaGAniitq+kKBivVO0UuKMFp2RPvyxxs
Rtk4n4gOlV6QrMOeW4h9hAtEeBEUp9MtysJGUKSFR+HUt6UXylSdWiSBXMbbpJ0h
kyKcXRgLymdmNz80CO4ZCORlsZUSj34a+5DpiOGkq7S+XDXBN3beRAgAkt/3eVkU
u4Or1S7peNKrERraXp4+IHwg1SahhZwjpLSs/OJVhwmi/JHq/BrheoWCZbeKlsmw
Gt9VhCA5g/L10GsUFADHQeDi0Y7KOyU3NK6YI3PoB56B3b4rM1ceXeu3jrbamID/
jzF2eFrCN77OeBLFFVDxWJp1fW4iPb612CS6kYLdCmahZv4KYPtD75Lqp4Kfnge9
9TYFNK8LcoZpJwSHXVgIjCgmqCokCHvnQP0rCegHHWeqOHZIbL66T5cEgHbDf65B
ykHT0ZYDyP2dsvN1E97qot7iNpktAEZfqSrOrgWyHrzx0Y0TcVoKF5Xf6l3RKMC6
UM1tseL4dKi5O++sPxK8umdNBYddEHPPp9WgaIN32x9kHY9OBLeIqehPt87dbd2w
SQa+hjic3c7uSX74+Q2L0FcZVknghmsmiFwJX0JpA0jYkaYvp43an6upJBq5bHzW
XrxsXX5KWce6rBfGKOrSSlaBiZ/suJ+H3QWtfe+JxWJvvQwO8Ov1ZsXPVuS6sMgj
p93OHjjjo9pK04niQiOZ6efE9cG2VI+VdUnDP4pBULa7i6QKNKjrpF7LVxBnuaW2
nhH3MggGI+g1Ie81pC6rcpLIbCViesjojoDUrn0FsYyoC+MVDlz5Wr1p6KEByPVF
MfsiOhN6f94mRcbwjq276W+7p1sUKtkF7/7vjIWCohRNVAI7XvaKFUNdjy/mYgil
HkALl+MhmRj1FwiiaIGh1n7DNfqrN9t69+1PNoLyrV+kTQWn1uaZQH+PL587qeQx
2kH4xxQp6EFfBOyMJdXboiXexLmQarkBZBgB3wKpF/eCU1mOBG8tDS0iVaRHFABw
5YHm29Fl14UfpAihzfcW2OuVX6ahjZl5BU15VjY/pAF6kKguKjx1+nABY5hxP4aE
Uc1JbgtoOlVLLOoD3RiHkGQQQ9lxHIwz/P2GmN4GtEyJBQJ7eLtyElMQxmlKYF5M
zo1lD5KMeXcla4gHQKb7epcOgLchtVvmTiiWQPwCGXC2PmxzwNpe1HiMCxkAlHHb
z9AV25toL5XiyopbB1x8uToYF1n8uSaAp0cVhlTwBQqecVj5jyxdWC1R1Izh2G18
XTe/xFnhkS1dEWLPZ1fGyS1tnuBG4AFPfTxjVwNO0auxajs5SFXIl0uj2FwM6+4G
J6Haus43LYCSgoyODZo0orT5OOmkBFvunsCBz4eTW/YFpFTafjxwZmar9j3ZcHDZ
N0i9+tLTrB/9KblfavuFZ5tiQuiEwgXp8tglDOp/n3Ja2KUU4L1x8slfGNb77aNi
CAZwKEvqXidk5qCUiItmqnbSQRk3UsA7aapG4VybQtQta44Rz+P35KOfrVIQ9zgX
p+YuS7ueW0jq6lRn2mj+sBdi4IbFO9k0/FEc66riSn8/W2PKcYJqGyjUzOQ6ypkw
jt2+mkJdlzywpejK+nPKAaQWPZ66vtdyLR5EjYYT5OP0NU2WaCrPX8thKaVxoGpt
YlsD1Ris6yQyVp+cXIOUygPX0UJfQcTD9KYdapgiyU3x6Pug2C2JwNAVw5stoddj
nC5daDcNuhCS8xDsjWI22sBSV6078tUT5OPfGB87A5h5JOfjsW30wc+6UTri3bSl
lUjuqrHx+LJEf56GUCwiVXAH3J55d0LgKuDpGK0kGD2Um+PC+0DEDfnEXhi0IySd
n4B5RpcTHN7r5Q7fDal2t4UfpPoSMIvqr3SI8AtZPj//RkaYUuFeg7hCmfJbwTT9
7CwRwTIKQbJOZnfd+NoYdyrijsCSedtiGjeqOt4Ux+Bxkt0DXwlsGOoFSmWoPFhJ
Fh+oF1RhrD9B1OGtcdLx1Mm69PJRNpwit+tm1WiFF69jnXLxiavobYBQ3TAfJh2x
Mq2SIE/NDe+47XYHoXo+2SK1Kzn8SvSjMHNt4pLeZGN1CB5iLKkE/ysUp+EUiMi3
Hp3lTT3ySLa0VwKZpP17IGb6BtlmKGpSr0brFowHYhLHJ960Q7ePXObCYyWvPRqZ
GSZ3M7GYLsnj+bE3BGrICPd/hV6mXV85MxKGQbp1Ha38swQ1Haxkal7DsBT55nDC
PCzJTmaHjwhCLU+a329WF7FeB1auHs04xg1GGjAf1PHn3lFu1JDkjp3QqkEhp7ze
iK0dhdcr+d44vN9MVbqUZMyW84zowh+XORk/bKbSNx0PlMaMVIfpvswStSnCvmRf
VWuxD5roKxoRXTrikwb2XDD2oUvclunrnGNNygTEWMg7BkOy2Iq5J1cXHaKwGH37
+/ShT4JdryZaQU6qG9QtgzUowpWpuZJC7kWnAArJZyW84bMrnN5rCNp1fxle+vFj
E8J2He2Gx+fGvz/QC/ylO38FOBB1nOsO8w9XB0IZ5TPl9OVkxanEe21u316DjKEQ
7hOXD4yWzZZs2W5O0kXG/ycwBXt8w0arNICNC1CG37Fb1bhcYZ5lIFO3YqnbI2WC
i934cYbzvPUMO9NrK4yAx0fPYmzLFzYkf8K4Dc6n/URwysWT20hdOOK+wIVavwb6
3uys+WPHzhwQpmvcmNKrexi0pIAFg6vfAfnZxZDAMq80K86SbQnGWep3QJFySWud
31rt6rvq83kn+5jHOM6rq+cqAQYw4sXPOedNMeH+Nq6g9w0yRlqnnK2i1qsRXJzS
pBkmpt+5WTsJ6u1PuaPBv0FYr4DksBnxcm2rfw7+LR4dI6Foed9F0cvxS1c+m8d+
VNQI1uTNf8XbsvwtohuGxI+M832XIsSEGVX4TuGGniQK2Q2UIKS+Pu2eEaLSFAxn
qWhAomv1VXUxCLuu+ty8mkMuG3kr8znbDwypXj1rBA5ENdRCbP3FaX4Vgv/GKpAP
c1u3c2Wr+ukSIqEx5QWw1M/qnA92F3sj70nW7MMFKAjesLr1H1xT/DakGmZKRbqk
1t5J6/NbiRqggQo7zVaoAqDMiicxXi93Diz+7mbA7667njw+EDF7IcraOIz4rvsm
vjs5DFuO1WYcLNNu9wTl6FfNVSIjo9Vh3tKPAzMoEtwdMch6ISYtfq+20SENWgw6
DkS//Nt0JJtCVUeCtXtB+Ugy/E8K4B+cvzA+M4HhonxsBwmkNA3el0Ysh+A4m81w
UDUKGd0E4kbiascdiP9giEaM8EoRZ44Dgj0oYky7XWE8RIHVLUl+axZS2a6s59L+
cg4YOeR5Ce1XNJ2jNGt/zHmVmT8hoLAUabe9eCI8blulB6uXiZgqEgoVPZcQ9Dk8
gEEZbUNoE0BYYpIBEnEDfoZY7j1TO6oJx8xUHm/PygKZCG9h1cYIQ0fbAbP985SI
MGgPtUsi7VgRIWMZVThu3IDC/4aP11XpaibsIKWnNvl6Z4YcDsqlcLfoPYurZ2lg
49F1eI//2vcSdAJWre1WYStBwR1Nmf8s5S+/K9g9GqMV1S8Er9qanrLhKeimrxIr
hocp2Xp/6eqiuRz/ocLjCbXu4nxVe0sif3JqSoa6lPES36cjZJ85CWjWquIrVlv5
TfDei0Yy4lBCsrUdmTrC95Q92A1QpGeQuqcwhyO8j9i+JpwILJpbuN3MPfWX5mUb
UtJvPmfHA8H55RV5OH1kOHFKT+uSXGAC2EZnySS3D60TfVo8iCPqp4yGmeLpWtke
NktA4SLM3Id4pIqFR6LsAXwskTIDsalQUepzC8E0tWEbeXE1vwapJ/xIZFy6l5dU
mSdWGT1FwZpeHBfhFHwsE6//Xssf/QmwVvQ5A48ceMFBtDHAzpB+GId+VYy8XNoR
I1dlZw8BsEu7OpLFi8E3KZS49U2yDY80ZKqVPp8xKurlTcmdV9wGhkocXIsv/c93
utDMzDJk//OOLs4WoZxOvzx8aJpxrHC8hB4Kh3Xr3ZuM8yvnfMfEmTuwmV7lwGVs
Fq3eVhgVRhXxBpH4zW9igzcxMeDOoMnsgXv3UPxXG3RfkQcXAfBLfGZtfrVi2uHI
PKW/Kv4Nep9QinYt4sbDH+bYSbN8n3FEZkw8y3EJx2Q4uoN5sAcx96/zmwv4wOIT
X5s9FoNEFEwqJ4DquBBvT5ng2OUCz4uAfVCbTi1qCOcda1FB7TJEzLGcFD9s5bKQ
/rJO5F3H5UYlFSJXI2lo9DDeoaTRl8r0c8uCwlGS9BvUVnSy0szhP7FIOnJz4U5y
x7Po3WyT16iyjLALQ0YHU+yhuXJQSZamHFIxA4mf7z3x9+P5MGBe3pSTguNpLwrN
7pfc5t62+lEB0kb/YvToh25FuJbdJkexbWsPQ7bNuLHRLRFcYONVLXz40+1/13Fx
p0QigdrKa7oV2LO+MTc4PUJXHfalwwo2FwQ4jp6Q+LGouz7ZtOcqbDMcZg0YeX0q
lihGLOpiYWYILFLxtWd1n0STuK5T6OFyQeDZCcZ1reCgFFnBUWmfURQ1bnIq6Dgh
akOymFSAKB9ifob8i/Z3dc0Ub6eVaQOL6KZEVvH/PgcXtpd/vPq+LAsqyOcHOk4e
31YmWLYGBbu379p6Mpa3M4HbFLwVJEaHFw3RKmiVjEyB6drVzp60hfFhDQSpRss+
SuKvi4ySdQryREw1+SPPUIc35mig+SmctV2GdVEefDRud67Z8DXutdWGmUxSc84v
uRO4r0aCiVltd2zUw1ph3mQchP3siSso5kji8ui3BCSp2EH3spK50zWKZU+AMN0k
TLzkWL6uvY+pLPHfHQ3WdApNdM7HrJtl2LZg+tKE8cF3YGbZMZtN6pTP8/loT5mz
WXiaAOgmve0GDDvp8hr8TaJcz0G++SnKmHTkmEs4HENo1+TarGCrZsFlZdZMnwZb
yQddmwoF3L366fO+6F3tZJhtm9cmCrH1JfGikDtuuz0oeSPflGRHEs4pr2+O5vHf
6B0PNV9/T6RnfsNeuQpQxTugIoQ8LqWYaq3J/kfz3HCogxENLP0Hz92q+i/wqqST
gxMLIt88tMdfSvVFRjdECqPUp4clR6+oUDsekytYnK/pzB4Ajw0pwNV8pj9ljRh7
D9cfRs/gf2rMteFO/P2zG3CBcZai40VREdBvY4bCECUoU21rgcSXS+/3EHpaWDe7
f23EBDmzd6KqApFALsQPRqrMqKpzpFmplPUfvD3DZF/clxqaltnVITmqZaQoOgnP
6JkzleKoMrihBlNvZf1/BVQwzWyT/tuAAtpN4067wivkKEKCCT8Qj58/1gEPMAa7
NDaaETAaJYdi1+dGjQ2tDneKKkyfu60PlrLPrg+c3tmcc62apcu45mfJKK0nWE7z
za7bu0kbD9B524QwhfvgCt+sqbpkmTeqm2vSxn+ZquSISrJlzUgaosOJVu2UH9Qv
zAkAWA0wBRWL4irmEhB85Jcd0ajTKC+0pkyYP02LVmprXOz4VhuqFVN9RQ30UOvA
+eAK7ongldsiDtQJTrHnBbTw3kFRPJ7IFVY5wEqF1vM8/4C7Fxts581vjW7bveUn
b1fk0uup9QknbmpGmBNOP8RkbR6g9Am8/JY9lf+DeSs1Y2FSNwv6K44tRvyF2Svq
sYftQaXKckajgOII6kRct7x3HVp665JrCDmW+kHvI16VfEg+xJ9e+2KRIKg2wkbR
gAaAewxbYJy2Nm3qshVZ8Y6y7x9VcY6vDMBI1kel8/G+jqKItujprV8FjrhwtQQZ
qBgz7KK5w+TIVrK4cZECHxqbT/m21EcHdgB7Y9Q2MQIAHpBMxOMMMErBT06ISryt
kGyuVcidsGAYI4nftK5FQSvl+0hYFP9lXBn+Ux/HDcYBAMcQ7gk7Ud7VnuzRCh2c
uNh19H9Vvut0Yz0HomyIAKKPboMf+FvBU3IHlJR3SqH8tKjB0GK3jbXTPPkFvP7P
3t/UJI282c6J9+mAfHTg2M+VFKVlVT6ExEo02MVNoSB/y0ZzOwiwfFCXgn1TNitN
rhkqev/CoNn9T+HUtYm4IrF9AEsFJepjJGgZmyswTE42wqBHTigBHCp5BHH3+Ak/
CB4q0tMHtRZv4KkAanQQ1Gt/BlL08+I1gdiHPx+5BdVBsG0hfvnenhUP912Z25R8
jTzQteIG3+E8Os8+O2CQMgwg00k+l0Jpin8IT/g7+lvjenmQLTMc/3OUZ4VPJZQx
c8EWLO9fM3oPD8CfXyRLOcVhBKdlw4ajX/pK6T/Flh+RS7LPFAvdwnV0E2lqk9uZ
UNI45vuZT4e4YaHHWgZSXSZQeWhhzYBYDHIxbI1taSDjUDmGC1IkmHOjTTjOMiY8
NJCXZx2pUSS717VW2961HBfiURTNK1d+4i87GxLg06V533M8DDeZ4VJvU+X5aXUm
1AukJq1DcSwhuQYhskIAyoTMU8qxQibkZE96TENnpfbgwd/Fo5joVCin8BDPOH+k
w2LzcE7aKfyv6AMYIKbweSxit5k83iBRbI6tBv5miJucKMXER1qKA4AUKIknirz0
it+CXzCLYAZma+H+v7CTIGnCEQynOS2UVPv+y/EjJYyrT9gQYRXhnktaiIS8CMIv
t+MSdQxttLMj4zo45CAsLAnuslS/vM7bKAbcDeiNOu10nX4ndMhFiXLdRRi23Ao4
fnuuMqEYuSSiM8CjFj7Sig4Q1whI1GAwMnlQIOnU/7zw+fziXMQnpA1XMdFHZm5F
OSVZBILsyWGmTaXqSgIh1nOiGcuCwB9YOANbymtl+FdZOZtGW7WqC3j0+zns7Kdc
F18rtyknPkn82RlvYbFjYBLO8kcVvvBTEarDEQL/c5cUEJ0kwtD8k6EtULpP4SZZ
hIh0L0VpkzRAfIjVxVOZmDlJxAN4g9RjT2munrxln+MxU0fups7RIn/EXAhKsAoG
KjNY7X1zsfdjW3VXspg2dsw1X+7aKxrUcV6yXllZjhI5c1iE//8R+7jxoWW0BWEJ
wGk6VfgJA5JoU3HfQgneaRoF3DDrgVpTDFFnmlueC0w0FQJNujtueXCbrmyQKXOM
Xlxi6ZKO2XGQNGtnJuG8ubtWAnpjDhJya8qavdPEcPmlUeDNnRjHiJcCFl8+D754
dYpNi8ix4e3elpsrY78rw3431BdrZ95xuc+golv5AGeWKMPQzP71ab64owWEeb8H
ZHJgR1qRuVXILSLGJ7btdBBuFTfm+rraBUxskRjs/+kb8ltxTOOCUs4/xqiIqdQd
E5LMQIfUyYoZ5P1vAUGYKi88pWeHwkh8SxpcPsUrkLu6wXWKzpqD7xyzDlvdwflg
zQU0eLBU7IrNX13jqlUdTpn3yedO4KBJtpiDsrPkX6gWEBco4M6pn8efrw/Z9KvY
g8UEnQrj6c+77USpteoKwFLZkJY8+DR1jYkDhuIOpppwac7FKQEpJOVCsezI9gnR
oaFn5uEUDrXSOrg2pzL2ufasXoQCSBktHmsc2hLyI0Joka3eeDiJ2dHK6N/PWM4s
xpEPhHiT+jIch6KeNdR1n44IxZGZZ6/xR0fZ1WmHD1BivdlrT/BbpXzM4SPP4Qvo
Jvqu6HX1GzsasJUwQl4Q0pku/WosQ/CiOJdx1ZM3b9ZaRJTt31bbD6Li4UeGRzsC
okJGYst8B//xZU0Ru6tEH4TwrozKjRNikwQR+Okbig5fqC9n7zCfQqPyLQ8n0aFX
XVbjE9+XLDvvkoLJCz6toNcuTFEQyQ/UtEee6gMHfyLmUp8Zr0GVpE/V8xh88VX1
LeFwZbYKAZCvaFssguD38xPz1eI7Kh5SbNz7blcAcb0YPHr9P01QwEpEXGA5VvXR
TY11VH5NALJZktijQbXivdHAUZINIr8VMLgRNlKHk/sat1AqFUZVtjYr3jov99J9
J0LXmBVau1CJ+msPrYPOrVbXq1Be+gMKy0BupGD10K4f9Yx/8uo3oKbQvunw5hcJ
vpWA3Gmk557D413sN3Lurj628++yT9ufbrl9K3a78SwYsDFUfq3AiARJ7tn+Kl7i
okzCtoFx4esigNzteZrULA0vUmibRm/HGvnEieqA0bt9i8wsth4jk/ENCzRA4I4b
qYM4euDyXZ5bi3guyeFH3FFHUoq3XgxywMiNbzbGVaZJjWE6M1zyaTVmxwjxTktY
9sIuzrfElJjV/ZUhmVUDXL5KcFp5okCOiJkB2DUWWXgK96ADNjXoFti0GdZvhmeq
kkEDNTR6KxabyWVBeUClbkWaWQBWNVlCBKXcU7NTKbh1hRBm1pBiiFE59ji1qBOX
b5+WLwZO58WXyjIIzkOUH9duwo7C71nMOxn++fHtQn+44+onqV+vBoXUTdETw9Jr
FabWkbjQCDfYk+uyR6hjs6GBt7WxBOBXh5x7bAgCzIfvHoa/oOZmuMzHGHq0ZOOv
DZ99Dd6WzqYiEqeyuBWGh8Xm0bZICP2l3HBqG6fcv7WDXUuJOg6VkFMAGxt81tqw
eiGO1pK65BcdKROD1K+agYjb48SUPsGU4UPozkNVNBBy+qUuWDUqfvVEd6l5qpUn
kn9w+c2US+6BOR4N+maCoPf3QGtkY/OwT/mYyjKDHXURfZ2BNXR1EYQW4C6XQdY0
320d7TbeNpDSGmaCZTBDKM41v5QmDYY05dLbCrm+dgxBAFMdepvs0t62qVmZjkOY
1YDGTHbxoJKDy5A7DOnV669SRgJBnVzEaB6rfstKp7bepjHFObxhPBNidnn6lwyt
nNOjzJnfqJQje1EGc/8RugpJ00ftNtq5HGnTucAenUTi62CVYDd8X+TOMcyrepUU
zlLZ6xRGyWndLWdDO8WF2KpxepGheeFU6dQRwLhH1F0p/42MYRhdDwdkGh2UZoEu
ZKsgJzUqOxAKIyTXbrmcmbzbMXlFbt56AdKETJ3SpPje6ryDI6HbbWIR4euYPjdB
Xbr6PNwpDzVceFWXEpZhKGHmywyuOIXpiSzXDVKNMShR2yN2jTkEZ0f35EooaQLW
scu2l3rDXNz5Hc4EZPydyncS7xzVdBS1AysU76tnGyHIdkA25J8kM31HyRgNUKLw
s+9wE9HTyj3g4AwpTeIWFQn+x3lHmGRUl+LGQ5N8FegfSK9RW1fiJt5rPc78R8Ei
XUJdlmwmM7Z5nv1rbQpsiBq8/MK+ZzZxXNS5di4v4AsUAwR58H7j7z/YHNYXFuMh
CW9V2/cuG+E7criWELlETOC2j7ph0pY9jJq3HhZAWeO9e4gHlFcN9VOgfPliT6ph
d7+WNlTTBckUWCVfB1gghVaDf3OfmqL9fsaUlFNKZ36MXKwyfoS1dd9ZTYxogf8C
bfYwl+OSp6DbIgJIb+zX4u1ABQNWPIgvxdxsZjiBQ5cEnE5TcrS/2amt/uIPuFLL
jthGgxquRpv7LJRWQHx+Js/XxdXfwzOtFjfgIVGTlTh/Pu1OCTCGk3DyewnZ2Sra
T5vDQ2zp7esNW5CzW/4zzFsO1FdgU4zdJYAG2ytvcRMC5hNSeAMU0iJC3BFWX9R3
kzrGB8bsY9iPf7R91HLpvORnO0cImtaqMYh8PpHahTcTK7jdmAJBBxKQVxzVsVuX
JVLkbgnfrbqAXuc/fETyt3yASxFN+kNCG4KLP5GYpBGUz+tBGkscAB7CbW8o9kWY
rnGzM8VfYKewNB4jKT4Og0+ZKTVUZbb6g6e1iD+AfKAYYT7GZGvDpgddW2SLZUqY
ltBDdmsJATtocvd4yobGiVO6q7WXOEKCFXpy29CL+wZCtcK5GrI37fFIX0Mqd6Fh
wWG8gerwrMFgrHq26oveUm/kelUNWf3Hl5Dg6Qg4t5gzVyzi12XmXu+LGH8P3mVa
qXmksDFc/PdBAsLw7lnWfs3HbAAZulzQojlMgldS9bKkTF39FriAA6Op/eiek28z
vGdLhW76cgosTisXdr8BYpjzeB9ruucXYnE+kL2LqetMEd0w+AS6FHqVEEbdGZPR
iXGa1xEzg/S4+qDLHYfGJwhFoCqIDMODz78zlif26kzAMlP+JS6JEJbMas5K0PMq
hfcpgMkb1UYCMyFvia7SjLMWB/MBzED/VS9DyBT9Jg53MY+2DUwj+jg4oQ/JMSrV
uUMyVYGwRRK5TuKBsJWkotN5cCUn9JPA5kVcyBdxGlPtcM31sA67BkXtVlTrxGM3
VchrSIZpRunv6S1ftQ8+bqYVDgXYpKVFkHkGvQjB5LSPZ0PL0Bkm5TZkBx5kacQP
wVxIXMWQOHSo5+SJ9ev6MV5wOIhAk5co2s79M5571jtI+1EKZDaqFjRbDqXY7cNJ
pm0opiWVP3XzOJLHCU/f2Ex30XNJVosu/8jjxFJ/rvBXShQjp0izTF4lIIdYuQqU
nX8WKTpdcoEf3hRGfVAzkHYeWQ8BmjdrlZYnK1KUEHHcmUVj6jum+Hs78mT8kLK8
8/ZF5lNZ51OGcDiOko5jF1t5HnsFP3C/zHdvjA5g81IWGblxN6Djhvpn6tvwYQN4
TapWO+m2KZLqFgBDe3Ug01Ll1Sol1hz8Bvkqn8pQKNZ8iYUUhjPKCxzFyYd52ICU
oaJzmeFCPp66gsveZwSImW4ONuYXSUHf3bY1W6I9DT/rD/AcCWWyU0vDxTYlwif8
DFOWWZC3REaZkC9sv3gIcTp8yR3QuiMhAG9UUQvBG0gd4VfaTkM2yIEJjodxzvi+
wxsEnis5f0W2+PZ0Ij5MzfGirTFbDFdKqnlE1eE1W+dSuiNDot+vPHZCPMk4F7bb
ViIXY2pgdXf5zCuWcks1EDqiOIAtA1R7MCbwYUOOezQXidRL/m3xdO5w5qGIQaEV
3NTzpkQRpQ/knU0A9q6spoPVzWcFBjW7dYTCoeUhIPR9qjwQO20pUQ2JxnJYSIsD
5gkhiAhlyWKfV/To3M/C2AqeduqysE31f0d5NcASBSlaqU60eMZN5lkHm3BONU5s
32m2CAY93XQLFU7za7dz2REUwg9mJWN7EE01wYDTerEQsqY+bwYoyZPygAVwLecH
gp7RPVkULgbsOsQN16sKDDLWS1bQ+4ypz7zjO4j5n39/CaqY64BUhrxIaolq0vjn
yjJbBDK+Mhv9yPeap29kurP2maYq3jkAeaQML0lFWsEm3EeIxpdIILZddeQUac15
E2z/InogKIwimaii48bNaieiE9GUyKBvUVa1bx39PNhPx+nMxbUV7JJ3A7aXsBNR
kd2yVUu5zEm0VQhYpWSOagnCWzvWz9QkGf0H5PL3pPKHiigHYNrytSZMDWjvI5Se
R+HdOO1xgtrbadFKSzi8m91w+yvoHg4vUlk6mIG5P7PqIdbRmqyh7Qavp8WOUfDR
lQ63nHauzFOM8OkZeWOOcrKqRasXgKzxkiHA69TXNcD37BMc34P2WHumbtve1sTB
gAI0g8bbWLi5f43FZyqxrlx7gI0Yxo8lSQP5bR5NnigsfFUjQq0KcGJ19kCYClYw
/xi1HLeqgAZwdhkKc5+yVOI2lDcBOuf+uYoE4mRlI/k/Xvbsvq5nOO5B2vsGzx5p
TVg/iJ7+eXdquXDb5Z3/2dnzYexFD9k06XPVeVajGAd4vYsBelmbN+SEuCjBPTfF
M7p139SD+6FM5AMbpgkKPxetipTTQzpza9TqFyBngCLiPsMo/SGOY6fdssbOWnxz
GrVs2d5kCaf6FOel/UjbPu4jodo4l9cvDNERchwV1dgzQVrSzT0pmpWApqhVlQ1c
y9E5mFXhy9Ggjqe4lokdlgAOhMpZdzs/fxh2T8eeaQwKeE/lIQO511E6pwToSxvJ
Fv9np9xjqLOTDtJQWf7z5TC0Fm5oMKuM/x/auzxvNw78XzgmtGKYa4hVKJvtlBSk
wsH25i3Ms2b5UX9ReCx7xQz7stlnp4NOApwL7VnY7xmLfsRKbObPixxJlRq74Ffa
KAkhoGv7TBMGmi0pU9pd9Q3A8hTMlm3eKzp/rHkHOw032dyBc90pOGf959xR8B0c
zyziE8VtH1z6ViOj4bhPaCddtsLLPawK+LfC87B9r671napyN18BgniF1YE6EXed
1mNSX5IFh1KZ0yxavM7Ihg9ldpBfEBOvlSXF3L1sKL0E/T9G1pY2CDLdBNhALQRA
6YWBLCTrivOzZRhZGPhiyVG0iqKC6hNvCYnAIgCjBoi14AYDRMZbA2980pXc+Ehu
pXcMGVHWyAdoAheaTJmIk4bMv4qWVxNElfrFUwANf5wqLiZJC/912gvJwCfiO+A0
smkfKBVCvodnmfPPGT3IC5As+cEQIDzs2WnlyLkzpITn9QzbdHl5YF7xGn987Kp3
al/GmokhDNE5YQyt+x/ta0iuvJ3YmN2qjY3YHvo22Rd5FLD3Fqcue2Slyt8uO78z
LZR6Np+/ZBLwVAYldTyRoXIzCtPWzt4UCPP35x2WqcbWSDdCSiLNWR2z86IAJPXU
pjcoTvssIxFyF4QYcsV95Z1haDCx2auXb9nfmzjipUGVNwo9GzpfZA7eG6JN+SPs
/rmLesLXpwlGDdSX1YF0WBhr0AkR8cJDtZJYs7c5bBnt8vK64iH0SdrDfjtQdJUl
HoyQWxzw+EM+wqwJRDkm2lHSjPVsgzBwUXZZrvkzoaHMVq0nS5bJqIeLdHfgtTry
JmsNtO++OtG7vnTRR2whhITiaRhf3vQ5eVNa3xZpXBrmqxZkBg5Nzv6c+AGn7HOD
OybpdSpjOmLsQca080Ntl6G6mLRTP7JW/S4jMs+ICETYn7I7fuFutDXxAcW1vjPt
lueZM/UdfXNToHi01Tl9PwtOZV2S8t3L8tAjMNko0DhwfdyQ+RFyY4npqyPj4w7i
G1FPbwd+NcCvSjEZ+d3iCbXS/cLWkzoMhHkb51lFxebwhnMBzsP8xiG02kbiO3Bs
sCHre0JBxmkZg0buRkIE3aeSHMvpK+r6HyLHM0uhN1QV2d9ltqH0iI1lTGlhxHCb
6e3o86XYJNsi7/fu1qaJODe95fXUE6V5C4m4eUCd/kk/xzExYTJ3xLKu9/lR70OC
t5Ci+Vn6sF/tyXhPIeoseL3M718Q1LFr9cSFLIRUA8a/LxjiahZWcGGBeWiMQlol
uFPmn92AeKpo7tNOyJtQbWR+Lh3LTUqVC1HWVTvsWMs3JyLv8kjcCfdc21RzHAlM
jo74Xh5DqTuDA1hDGKGqiSY2zMDzQVrniRwwUYfVKGf+92Jcv132ukNZnrgdDIve
JrA2K+nQEwkh1uVftyqPyiOtoXGwtToKQfqtSf1c8rYyp9Hdnogdb/tyik29KJqY
o5/1nx5NbPLH/IqVyNUSzesCXIOjIgbMR5TCCEpw6JHl6d3eYsmu7Xcv244SIkUN
yCtPAfrKxC3KzBQrBXH6RSHthOEoiTw1WZ0Gzwgob610MRcea4qVmRKEeTUv6SJN
Zdc77kUtBPRv8FcPlcX0ULotX4Y10ZhTRmErLZza0sog3rpDnmCYT/T6aJHKnJsA
hUHW2ECeGgwpdl3KCYr2/ooQ+BLKmSOtJFgzIS6M5F2pCF4x17apg7/LJk9O+GBl
Pv4KPO3jEJReglcaDbZwFeas2wuIW6Eo1RHjOa4xkYwM49reSk9s2r6vi3uruOf7
HPyQIrc1kwFRx2vwWKgahFxymMQwd4EPx02mj5GdsQv2tQ+PpYOnBav9NYis7asD
qgbvhJYEJmN/rQIQkWorxCfaF4Fgk0w2+Ya3zAzVExtu7i34MCDF/XsEBlgFlLoK
Jpvl9eQCXzDPiOdnWrubBYo7LakKaXpfc3fuOZfzwWMOzTHwxVWHM9jnr1+6Pgpr
Z+99gzZOEJQFXj88rMCET2i/sm6w5dLQcNvCgNvWBxaVe2uHrNY9xjS/ZIvNhCUA
LIpMre7RCtfMuZW+yi31rPbVCLalWKLxmGi0Zyv10oBOXgX3j1jb+wx0IzwB/xNy
+oofuTm55BCVv6XtXP8OszfhoyV+E5jjyjGte/WExcOQCwQQFLzFM16ygyx1itdB
+1Pyf3k4s1u2dN85/bEDO1TMZ/nHGTkwjJiYfkG/QTDpdaJqxbuSfNsBXLstm5jY
+xQAxxgHnM6fjr3WOpOOwaOGdkTASt7j0x2RnXF8lxLG6z7haDc2N9WYpLcj/eO1
rbd+04wi5ajpcMuThgqW98TXcHhdRoyGPHSHDc9iKmOMmKBiL/WY0DsluAMTPCpi
MSeCxanaoZvAxa1IE82OXXaktUZ/id6st0RL/sjWDFwLBIAti7yVofQ0SUT6z5PU
h5o2030sPRCIVt0XlyOd0I1t4WE0TiFxpvxFVHOJxjGTLBqkNijbsYHzeJqMA0I9
gTGkSVb09qvGS6CVnwSh/nhsdhJVnxeVmwFbcYDClZHrwmzjiFQH6WHt0DoPwpno
WLxW0WLISv/QyyEI59ER+6gwd+LsWndEpdQJIk1AGQiwCQmYqLYrn2trl0f4DbxO
WlWpMAyuKW8uPjpVEZr/172upelbQJS2YnSQyQaMEIM9HT8JQVWdC0wgsuF5LYdC
jJnOok1acufLBbF/kFrh/wXBv0DuRyoAifxy4iNZpwTvkAlRsNBRWpmmgIMfmyt2
uKMs3Krg6t6BtrGJoHeCKW9u7tDG17rLjBHEWgI2HRczKMZxb906luIDdJOoNp9s
X7yWz+Zsw+KU/gQ+VKNp5NudUk+yKRK9o4n6XwcFcPRoOEC4A1a0ez8pYaJ22922
uocfYDBu0c2HnZkDOHR09IXstOIRYeIEwG26h5fZFpI68+CMDBKKuVliVELB8+fx
7qJTs6oMWL8Tt1DoFIymno3y05HKzDIZDpTE786aAi+cNRCROQvIQA2zOZ4oWAqa
6WbLd7isoP+T0uFlP9Q6oV0l8DcBvq+vewMhBxjlNSjcPW6Ly77O7eSYHGkHLyg3
NfXvzsdLBvhlYZ1G0ydW1FpaliaeN4gIHfhixVFNBJ1S5orW1zhC+Rh/4vHPpgKs
fbwQjRuF9s7xRpJT07np24bDC6Ro5AF+A+qXZ7Rpqs8VAtK7ZxN3mfTg+QI5JwcM
iCDwdiHOZAybiWSACwObOPs1NvWDoeK1/GDVTjTCtm71na/Zk76zqZI27LYPhgF2
0gU2h3lp9Hw9VzlsZHEC4tg/mPw2TYTSNwQwpg+nuCxXzEukuKyH2TFA9k5KvHYX
QhokMSuOpCJCP+ObRbFRFws9tbqWavbN+LMJbBapX03VlTBE+D+86Laep+WvIGzH
0OSWxk/hjSJqxsc4V4Ul1PdGB6MYEXeBI/NackwK1TP94Yjm/29I04PwcSebGEpS
Bk++4BUjy5ThIZqy3oKbSpbDbf7nHTDwQ7CWZ6BYNAnpQvmgY+KL6AwkiBHN/ce5
olFeyLVQ76uemkh/rhLWMT7oXaYmt4ABVpvyYzcl4+42hLqZB0C6Ra09qZwtUStI
hOQSbL1i5BN6jiY1441lBdjkO8w+liA6F9LrtLJfq24VtjI36BLEmZwMKmCtjyM/
y5OtnwjxKBvLv1X1wyiF5cfSdIY+bTQNfQQ+6zuGCfeyaOmkzzJZoxOpJh0fZcZW
scUxCV+uz1vlEqH3cBDd3FJg8MCidGV+cqa30h0LFOSVBXUI6uL5hc0VhlRgdWa4
bteYaSi0qgsKPvf2a9488P1MJeebU4EZTjx4Zb2UZfFzdB9DY2nyz22w78QUHVaN
PXxkAZQfU6U6bxPewgEvD7RNO/yAYr9LHutic/jKT4vlNuHp8PzQqfErzXxmNSHz
fyGMTziCBgKnLi8XVf4ojcBfxDYD9NcCTqI9B+4crlVQnxAaTs9Md38Duw+i02n2
wsWE9ig3h6OPverGECHLrqpSCC4xS/XbBE2Wh4o8E+EkKK7wbK/Lv1+itDCDYxEw
dMYVjsZndA2RS6KoyEOYuwxTM4cV+ZuPm1tpeexo90VtQRgg4XtG/ZEc6ByTHh2O
NAW5f41yl5zcMlDl3UU4df6vwok3TFt0Pu7IngqJNVVZHBC82shy73dX+TOy+oRu
Zfvii0D8ULpt+pc/qP3q3auDFLlvbzm4egGB7D0mAOB3iSsCFAqtpfku9gt10iDd
izQYf+DVohq86l1dLKIfSWrbD8HNsC1Zzd3YKW0okMiW0WR/p7gmE+7H5KlUM305
fQAsu138v0yAih4FiPfPZKzSigfRnIC48CMTNCMehZQOJZAxllpPhQaw59H8c6j/
SLrfpzP+nhmxU06gHzm3ae183p49WhxVAyle/9BYjkFgqkpDpGOTxwePJ645z2Bo
iUFEO7/8vdIK3KbAUCVBNIeWcUjhZGqrc969cJjEYypjqcRf6mDFN0B/77H610Cr
lpd/3xpgYFlzDumwPpVi+hinpOrFb58OWHvFLK6QsXDqH0tzPwVkS/chCluZIPPw
qH+eyyPp7o5zUwVlSL/BRM4x5Oh7uEzHwxNzGC+AbAMoXKABYnq9LHK5wEJoRaOJ
4mvCpiZW/cvpol3cg9fgiiK9syRuKrwUvqaBYubH3lCqPW4o6iQACsJEtQVQbkNn
rpEBZegcN+uviHiPBQYI7Kmx92PelcZzM63ifmDZ03kTFTDqBCa9vdWRQLrIxDac
5euEcvayOZyMKC8keNCa1SZFEgHxJcBNMg7Vmu22cdloNTmAI8UTRPXjNKdKpt1A
4Q/p+zKK5rcREIfNiH8hKyFjcGo3ZAWaCAO+B8q0oVf4G7NnqpVjsipoDGRHrk8d
rv7L9mlo9gOjMBRpSqIAduvUmVrfUJKz8HXRjlT4a+Zhg3gYA0pQwDBL1O7W71Zh
zVNIXh5SlZFxiKnSNz07cAgWwN09deHDyPwEiPMY087R52LguoNB1vxIFHtMeAjW
IujsHfY7fEAvAaN+a83/2FvejTyCy4AMjaleFxYA83Zk9XK4LgvmqrRLT05DULHL
gooO+LNLvL3hXDvxX1sd2k22eNZI9wO8qILhMBNz4baze+Q0OigAbGTnWL3Vjul7
KF0BjmN/8XkO+cKsBd7L39rOBqmmvfPwbwZ1QYN1v1lgpqRHP5ASCQfNvsqlnd1D
CBujA2ZtJiFhwWrpeMOVFGaRnfV38V8XsRac12xZjm5W9/8yaGc4skBjDbmisqEt
HkH9hYT9Pe0xOHZxg4pofyyKFLSmqUt8kq+hsTJDD83jM5hEJ5sfjlnFteOof+q4
CyBEe5kNlJodxRMif/Ny5GENhwGqHxMwJZ2qWgs9kENsrVpFFxy1D+DgTXu1pyHF
9GVtZ++u7jYh4E74Iu7Yk2SBhbvkqBfCF1q5AWrt1UdGCJE99ze+O2/2mbe4jXD4
GlO2ZqLRJ/42+V/LwRCGjts0RxrE+QXTSgk83Fc/3ccV89fJugYW70kCZTDPmd5C
RWX8LOdOT0JcPEZnEBabQHVkhGNKhBAigqaG5D7MdMWGWudoNWnocVpXFQR9SvXi
yOrBE3ZL1d0B85YmaGDnNU8UakvWUdXic8ImF6YwkQT3f8WxWmOnHoLTVP/0vI9K
Bg2mxwLl5Ok4Z+QigRx6iJ8svpAX3oXN2BibXg1t6xUx/1IwYCRFnrAHXke3Pq8r
mh3N2mADkg+WfLR13o4pAy5nR5h29kMx/ExCc2YYiNloV5EVb7otsHeLld/jB1rl
Q7wUigAbq648BY+c1JJ6vafvwJxvafxhehx2Z4WPD66wYwhX4jhnDNh6MBmrhcgA
XPBgrVBxrosEMgJf5nTfSsAbZNZkgXUzU+MOCsrfXQaTaoddl/uEZws2+wK7FGOd
KAe4EC3rV1wNKL1bNCOMZ5T4f2nMxZEfAUwcKca+O9it2yqg9AsMElyndneGKe9U
7c6G5XKXGOx+TwwkunDDiJxzyii0xj7/YcgAXYCYOpYbMZD2pHUqABuGSjBGZwbI
rRc5FqeFtWQA1s+rDLqtYaApYOs05g+BAN5AD00TF+sYPwzzFhe86+mWtrcRsi68
RUOrU+9HW2HwQG7OUshdHKJ2UJkIgqsOOQ4xt4W9IwO9E2eQCSU5BpvFFA+sVVWw
4VuBrcMHymsxyCr5bFkaTNqezb22gwsTFROViWy/KS2/1QuKWrwMfdHXp2+KXzZi
GSX1fmiNAh0Lm6MVXZyNAcR/BMB+mQypcGipNTWeAPWVH2D278RhCyBHADMH8Qxn
yhQgHvWSR0dW4I3wVps+x4xZ6flhcz0W2wGEIiBbBsquYQ9PT03UlO1rTW9unypY
hhwkNszBzZVze4CLapz63fk96N+QM3nDrDGqjwmLkP5fKxzbtQtAitwo8AbrPgqs
CvoCcYjza9UecKAau2QsJmkKP72g1C6QLh8g2axLqg4W9eDQFsuWIZySiMjDJqn2
vEtGh0Ex6fcXKB9FQOZP1WX4EfZurtwcnU5MrSEgckSVC9xo3Pgvc4XByUKKYBS/
SCss38QzIUVbUv60isjBtgDiQQuvgy6W/1Cv9e25RA3snCHdYwHbQIC0UJwTjmXN
sy7VWDqySh0vTYHIGP8y/FnLbPX6SPy+bOIr34lYM4KKwzMTkDOckDZYPaeF+ano
hvIatw4HzfHXOrwBLqO2Tlc0p7GYEf5225rvXd1cDZQbqhokPrq0P9B3RI+NPooZ
IX/cC7oLhvfHw8qTaj7mIpbm9LAGYn1rfK/F32pglnCBFSIj61jEIJF00s0HtRJw
onrcuh8qMj4SEx7A+R12qxKLBmBjK2iKs8xAGc6zprVRV2zhx9fGjXriEsGoR1P2
iWRGVpKHmbj1osWNdKYDuP8+0UjZKf3RsIFyCZQ8w5sYJwjGOKJqf1n6lMlMT+Kg
3qM//6q9+HEENzGVRah1gAiCEkIVJpzj+aKxZqnxJUSreOzadwI/hyGI0j18CppR
a8UbC2lCco3rTNUrgkswAuKcG7f2bDKMJgNh7T9mQ6nRGLPJoyQSmwsnOrO2KpW3
dRWxIgJ9ocTS+dyGem0W7a3kIOJ7Fx1tNVTL6yy519mepdXkBUJ8y3+wrR46Ljhm
337PPBrQ6Lu+2tJdU/VPDBN3173UndO36B3hDfBRupbvPDEOromM+xEk0PaQ5lol
GVwT4sfXMAj/zQAD3IsvZhmanHTBz9Qk7Xtr1qj5+XgenXNlNnAwLSdxFcC7vBLT
RKxQ2mffrmDNfixDcO5iUEgPFDP4n5ML8aNm3bHUpNabHhrbeJ0DwcsYPzfh4+7E
R+E+jnuxIi3HC+GutzTvnhrIUWS+m8hdVvWezxvCo42bmPQ9/LlP8Oj8sn9SB5xp
5/8zisJRqlDz11Z9kwSb7fYHbhhv+aPsRyrpcJypoxucrhLOV6Sk/zIwZ/AiS5EC
LACM2e9epGVk97EO9GjJgEevZQ8Fl84dPiQyp5uSuvEc5Pr53tF/MPpzHAXEXOKn
DDlWRGFAlWs2zJmL/0IOqdUYY19Q9fIbmBgoL9iNRgkrz610P9MJSEkOTDusPWyf
z/MRHps3g0Y1vki43YsJJi5JPxGDt+oHuPC4ahTTXM7dqHzCUXdf9gYwQDte4Iuj
PwPSYns0TsxdOX+OovD2LW9wZfqqfob/eOngxLCm1rEppNlBM8A/McvuDDxRWMdJ
dBbSDpozgGQRFIhvhpFfW1JbeHwb1g02/ZjRW53E5wLcLkCAtwuwHHrgmgjjih3n
tJ/CfVf6tnyd9XnnTUBur6xlwZhtudguxUnOTxjk98J0HV256RwhLN9pTpEFO5gd
Ja2S2rhYXJax2cDhxP7ngpkPUASVQTx0epo6R01wlay2HOGf5MmkbIWMQ94kbF/t
MHYnDpinSbaHXHD8h1GJ84Y4unASe5XbGuw4Ye9g9XyxBWTnivjsDHANWKdHjR6n
OIQTFs7mv3HkN2tDDknOLAOelphZhjMCcDEE+S8q6WZrVaCngGzTHX7I4d7wt7UI
RlmVVBg8+7vePNLr4n3iAWr+YgFNr8ygaz4Y0TGGOtDf61gGBmFsECNVq9EUJG3s
oN6QBdyPoFhcYJlk90BAlMUWX+qpOFjysiLJpwTHF4NVrERvSrDpyeNuDNccfyiJ
7wzhJ9aKGwLoF+z1cbycOOzy9hLExTN9PdkdY4q+CGRVJIJhkBDk9lmmR83ehyq7
Hl7dSJi76m2+xH0zTSVrFgqXK4/agG8/czEl64gkixe/WeEuIxTDUe4yI7gBgZF8
NHKeB5UM9fxW1BvPBd3/Nkfylbbb15QWsfhZ3zhS0v4tit0oUIK/KJ+LNKVlBZpP
/yOiQIwha8COG/HEZQSGnxqRPmsRcye1NDvffS0FieyfgF73xSqbmu5K+wWSYd9y
Rjh/B8RsDlwZySxDv3aAjlDFd1qM3K0qL9q2OJemxUfD68vFXW6Z1pGPZBVjCfMj
x1ok9yjH6rIfj8L6irp+YSUz0jiuSPdF/XjDp/eUFRt6UB6kfhvN+AbhWmtgnpBK
lNnotqPbeOR/pbdcOGwJucNEOTCtM9Mc4MSiduGVapKzZTnZH/igX0hf4wtNwJIY
FprctiPqG3YuuhvbIE4LzyTY32kpgIYVdwWTJE2YKUPMpwqMp7Xy1x7/V1Gu9Z/l
HqcKwXZI1Lj3muAtYo+Yuk0VK7Iuq9kHlFka5MfJt0KWmrQGdw85DYea/GSGuN1i
++zQNXGOeY3mj3LMoHT+XUch/EuMEsG8Ex9QSxQE7Q1SsLr/QnwQiBbK7BOJ6PFM
xMdyf95ApI5GV3elV+QGa0ujZe8dZIx9yECtG4utpzoUNfly15dOL5MoFy+3Y3OA
3zSbZ1jy7lM8dhKS7qJUgs6CW+y4eWK7xFQsg8rkfjnd87RCf51ZKknreewGu389
qfQpAdSTqwZ++UCcd7xskRZGB3vbrN1EtsGrRxHsbaeJW22h/+ZLTYfqWchLz+gW
xnOOjKpuzGVkqvAigk1CM5bB7BkSZlVYNIYYC1QUUgGBuSNR18DeBNhdrtQf9kX8
WNcg/y/UVupdvk8leOjP1F33NwjoSHAL6vX7TP3AqodI2PD7S+YQ+ivyHqxeIxrG
p7APDJHCYXn9pkel6sDiEhshkuvDZxxY1s0INowHe50peTDhiP9e6dkLXmIR3fvQ
4pNcvvzPENL3yB52WKvP2+a8kYE/RcnqAcocvjwDzmh7ecLNhwAwexvWtxRo/8fm
Fi9Os4mTxBqNSbC1cyR/Cl7VlTPX88PPFzwCLsvEExh4biYqmzTxWqyVo0DpLt3S
CGiMN1puqMJFwgmYUiGWN1WuzlNOcOIbNnwnI+cpFNRIkF4nwouotvhi7/bER/s4
RoGrPR7nQmDt5ekAWKp2EWgio+G4snoHkDFy1Jo0ci+3vRrftuM+qVYJPixty//6
/YzBPt0xBbm1mhaWDI52QlUM9rmpi/i1my2Pj7vO4iVIgpCK40UNP5jGgKbmY/Zz
Kh09F43tAIpHONdMes59opulVKwOuAwPuHpqjus8mawU/Nos4lJ6LE8trWuhQ6W6
2qcz2aDXq4WtCIsaRBX47D7uQlSTZjnEiZ6V9SoO8iuu5lWKXf4OW5E9A1CRvm/6
dLH24DeZcszNQPhrE1YopACOOO7HgC1Ci8MaAhpBcB2A8SZqdLwYg0dROl9mzQ5W
kx5oOUJm/oPgD8p0W7xje00olnE/YCYPJrViYTVqo/ar9KpKZCHHr5Ytv4zMipt2
iDoaonxtky2e/fn58a2lpps5uJ4UW7/dcf1ReVM5SRUTJwgulD/6MJ7O+46soXHT
EXr+GplAbnOpp8+amr1cH2q5fespESx1y269yoblrmt5kUSs1rLs7xcmoV+Kjo5R
3RpVgagzl1ds5fkcxdaFjXq8nlyJqN1YjFMdmO7sefp4nUTtnre1TND3ihee65Ov
qbrF6L4wQ0Q6OxzQueFgpvQSnhwD91KPvz0nHiQHe2yaa82LjNG798wHdLWLQAcX
GQmwMb8h4pSlaffc6izny56uIcAi2JATNYQBLrs9F7yXPAnhWsSPX6Ew1TcENFn0
q1Af4KVgeIuRZdNSiLOvwcNUT702GuPtUjtzT+fVdcNAx1tFN6yWC94bRh1o5F5a
SLCAcv6hL9a1NExXMeWKAnGYm2QrrUiVds5mVlplP5KhqH55eejWL4wBP1l5Gmgg
jxQTlQT2fA6sHGenVfws3MhtCtASFqGWvfKAJc5cXY24oqPHEzI115EVtrU7oWuJ
cqt1JCE6I11r1Atk7jv00NswZ7WUEP8xnnH0t+q1R5Gfe3aDsasOXypodiNfKfUc
rYob8quveO5cDW/nk/sT2FNnjMe1h1ouq2DyxF1dAnVEC2hzhezgpzMbrY7zpUkz
cRfjFauKkBNhU9IY5e2RlbVKne+EjLYhLCYp45oIsCM788KuOBbL8I1T+WWAXyH4
wh3r5oq6BDDv7P9Y/B8BI1NhuLefhGvru8j1QjBFitZHcNHCIsU6JVsFPDeSM2dx
850zuvS0B3LdvggCiD9OPbBcLBjo3+XdnJk2JLYE6+8lPvWtsmRTSHPNzQZLWJEQ
7Vi4V8AK4CtLyHnCdu0jT/6YFdxyScACu2RltSasAAIapJxiCsXeE6dx+Ai5X6Os
iMu6QrQwGXh8K3VVRsfiF5l4ukv+71j3cIcr3nlZtSpZ9LyEPEK4p/KDs/3pqQip
7fGy6Ko6e5tn/W6fAmbLkY5hxzTMKlOiDwhNQ/C/9qFTBYrolLfpxSFXk+opMgmD
MtufwIwNLCMHC6noJBIBXei9HfL3O+6IUZgGdmVZleFId8tp51Kiw3rgw9ifwxNT
zi4+FpDI9MYe7jq8fABqy8FnhUfL/fkjDrg80KMX0qU8lm68NvwKWKKnDD0bXmYu
ksJKeLLFXJ+37jJpd+y0EovSwqTgeV4k9VadL6Wzg+L0W1tR5hbw9cigCTMBULpt
9lyY5E/N6M/QjKR+j/Jg+1+mwYBrZk4WnNTLSBzDIS5jgDqkvOjSRhnwD2OKK10E
rjsmrCR7dfB1R4DgCVe5644eAFBuRDeyh9PcFahzOmiNWsipC1+1pBywDpKnQLfW
g/Cu4EzQ1Ic+qaKpkJbb8+ESi55LIp/kSkIWJXYwvtR/Uu+bHvnMMvIuWPLP5teA
t34OaPA7imzfSik98lP/9c3XWqiyCbTHPVAHX96wtwkaVYsrPMgy/gXIIgE3CPMz
EAqr0mXSL/7DuiPdzMIgqOCwInYbAFiwilrqqpb7ZTaLbRW8SWT6PcoMd04Ch16P
OyV28N9/j0u1uZSGko/fTiYPyS3vvY2r0f4+oWpcdVPO0t9fXVFSLvWYhIAFMolU
Kqx+2TZzfgNea+yICjCwz3ZGkasfx+iC6Yr7hfCtfQBjytwJtykWF5YgSQ5lvFXa
Zx0LBhMDgPqtpI4ODF58S0O9xrdCWc9lIqkR9jg97Ihvi6t7D2JWSnuwJ8JfhS0b
2O1YFwmqoyBWD15jxc03p4G2pNJa6CQF1jLzNR9FgF99H6J8Fak+gvyWjpQaxrpO
tio1CuCTO+7DyqLhb1CSqgllpMSOVTPI6wf93awdaqtXqslCLfwhZI0ZLKm5HHiO
Pe+00bNY+w8zEtuBCwYjjvMy5qEmE/fRy73uVFN6WpRIuLGKp6bS42FVsbfuhKMG
O1R+sFfv1g2z75GGuqGv85Mn6NasOGxZVNCm4ri8iE6eTzX/lG9b8KAplAqELoF7
cy4qWRXGIBcWJsru9bYZ5VDTfIjhIQW3SJ0uLvX1gZDJrkiemXziXMVXhRhu5+jw
L2P9IDdTkUfnHyrkXA82XEt5X6oZZj3Cl3dN3iaorCsDMgeoX9Va6gYflHZL+3Ym
9Ac3kiEzIkIOtx1fPjzair4ULcNkAHvjy9kR0vEMAt52Rr3OiCN98iLAOCG7/XrN
900VK3C7dCFov8bIDSqttdp9Ffikr0Q6JTLFguxsH2Pwzyc3SPeio/puy4KIqxEB
mI//pKR4MwV3TSnWGGWkSbFjcmW6e9MjHNn1Q6lCt2PpDGJ20m9Cxp1bMwqoTegw
4QYxSso4j2Vzf1p2PLx0YL+WyfwcMpJlGCHy4wHRwyxDAX++k6Is8b+TIHuUc1fm
9vkkfeXBjsKkqp56rjF1f5bRtWJ/sP6fJUEEyuIRHAqJAumEJjHLG0InKBJWWWdO
OtRDjnWxN3jZEgo1JAfdOU2JKbbDLe5CfGjY5qgSUyK135J2TVDJ4pkY6M5r2KqC
AC6THRkIYgzZUTrn69yucxrSXMnZTbZ45fEIwx4M/mWLVRtpYu5C4B71kWZ5c18T
7RysZdT94aD+JOhnwpIsk2+hLfTXSuJOfQ5EMjlIJeSMQ5xu0F4yAK1yYklKu/xb
qRzwWfNLqNkaTSACkHt5p5NixAffIEmxgBxzBlDDHdjAw4lTypTMeTSATkFQTUB6
67t4iKZCuBADQ0TGZv4/8XQGVBJZYi0VSPRLgAOrd9HSxk4M5iVWLNSUYtnfP4+h
H+PBrUVoeowWbeIKucDOK5J2E+tIHtFPMD/gGkPHeQQJhVJvAAvJ5vjpaYbB5Q8h
PBFJAx+xwlyGkmtNq8K6j1vOhPynB20jKMJx1/ymsQfLaYj8Az9ah2fgYIYapiqJ
FdN+oT+w6/sX1b6bIKGbwO/PMc7LuOc11PGC6ZUs4b+FYMPMbaoKWjTlxvrbU5u6
czpa0jJWQKOxYVJziOOHDnWG6uC9gUqrm9XQeoJQUe8Is8evLFykJhewxNVyCruO
3ZfMtkUntY9zCciJg2VPaKtYbWCdXfuoTgQbdCW36dciAu85nG/fhUeSe4iXD0Ix
NUnAdFE9ZF8Nj28KHcPd86HCG1G1gL5/X5ymsUMfjm1ttW8Kjhagqyi96/XZNkuF
eQV2bfDZBDMxayfhKtueBwjGk4RRNda+T/w2h/VR79xhKC4HaZAt8Ej71uYWj9Bc
IrLYvH0ZcAbQCu59zU5TOb03q0k/Mn+ELP3byOkx2LHPUHOpsg16mC6lW7RbZBOf
r5QFWVkV941YuZ+KNq8agzVEIuUlgObsaENUwBt5VOXidD3IZR+lAm2v9/oASPgN
iAcKuY/jNsrx0q4gFZMh1G5CmbGhsAiIZEAVgLwsllJDvoMDCTIA8zyUUcAmiXlc
LZUvO+/eOktis4tBdv2YFrcipsOZ2Kc0zCQPN4yUpWBuiOoKjuWALqAdKG8M02F4
UwprjxYN/P5azq3TqCnoFDpTJuvuuSzURiUhtTNb2MdqeVXsqFzPdOgHCbsnqumQ
g9+BPkFJ9n7b7d0pn8bxEmPmKBcZsvW1VRBM6m+UHP7Jve/C+acgfA2yEtbbeopZ
YrXocVsUQ5eQsNUACPZu0I40iwfO0o27iJkC7o6KleoDyqvakyShDbfSMYCDhb1u
+5O+Wgegz0v66OQ26Kck4LyiMX5zrUnAN/uwr0yGrZu0PZVN2hjbZS+kCX/dzB93
ZXGJcpwfnUdhVZn7jpYRdBtlKQTKblSYD6T+CeAL8GrO/Nf3s8vjZdlSChSy2rn+
zCcEr7kNVkyAgpUFF5ztZow8t6qnVg9ICVO4hACPHuDX4st4nfG+ON6vS6tMt37W
gPmcrRg2nh5UR0dra0cOJ8ks37PUu80Ol6UnkUP2/BtocjgKviO0e8LMFwsj7q0/
PSScB2UYYM3LmaBJbbEdqwUp7C9p/eBPk2lP29/xAuwH3dZX1WHoD0ayyKevx8eu
LSftRzW5zOSCTpemZ+wsjRqhDz0vQOj9FyT0QAy0Oo9Dal3qdfAWvpPs8l4ma/xe
Xy57X/6kXGwT7v5ogM5vedoo5ZcJKboYGOPaEsmZ03+bxLB+m5zLP4/WhdNhyuV/
ygRbEW5qrM3Bf4a3pmzVRDAhs9mykMAwJ2xGVrRoJAxL611eTnBtSTx5FsLbVd4e
ItW/8W9GAmn8hm+VGKmUg0SdeXt5pJAnKHsPTHKgmEvkQYHfGfv5mxhOsO/xbPgc
0O3TMs0/iq4q23k0DfPPZG4VgbXUxgBMQFlwuFDQHFA/6MdEurNNpEFlnFX2rT5m
kDnGG02ysnTD233ZEcG9PccGY98Vv05z0Ti5emJx2K82BISgkSgzgVd6G2Hx1LWT
ipkm5nt3oL2ymd5WQBZpFTppuv/HjMZ7SUR5GjgefPt2mpTMHKCtMTv/OrZVVs0G
LomqceiiZVftn7iOgsDmcqZ4N+9NE3oDoF2Hms03aHNJvkvZKKWk/bhdvVY5ng3E
hQTkQYsdEesRLWdsZ35mal+8GUZ6jtWun7peUjoR5Qewc3nAqGWpgpzBOzOn770D
1i/K4SSUNhwwFOCevS2yqdem3vshgpfnDCmri8lm9UC6IgrDCawRFZIzxBhczk/K
Hkr49INmaHVUFn9XXgHPBER1BOwqIT77gV5jct45Lh3DTsPblVKms/yJb4VZ9Dbn
CxuZU1qopbExAcqPclMZp2wun/jBuygcXx6714oN4NkLmHD0wyyElD6/Bw5lzPWq
Xd7GlA9HBtO/zyrx1PhSyQdhjz5wCa4DEwZFjZ2lCdZE/36iRxQgu8r9Csyx3IMp
8Siojze3vb5g0L9um+sBvFkeq3egv9aMBiZRsIrLWMyn4Es7J4pCgNI/ETRu0Yov
AXJ0RgDOVRf157SDyq8yYj11YAkHJJARM7rRRuOLcbPL88KNG3Sf9qunx6xf3WMB
nRzTTKbq0C3kCX40aFEUDBDfU1223qeHPH5LmYbLjV6hIfyAJ8Ud5GVDXCVh/qF/
NfxDZoSKtxgzdTtpfJq7hkA6GRXe9UYeeNPSG49BYhZLtxocXwMS6DNQBOibUxDi
6W0lAAZrDJbAlYBCvjcj06owGldBicn3d4SvzbN0VLVSPlEAbcxyaxQirwJTt5E3
DthXbOhAAe5cPtO7CNNheZRRlv0j6VE7B+cONMUymz44/EiwE1vsjNReMtgXQ4qw
r/P+bxyj6RNwOqdPktR5RzmdnDy8ruw/4eTm7rA634oTVqg02Eue0/jtylLsRdYo
w6sVRt6dGKzCqh0sO+D+w1mVZ+ohoKBAh1sAaw3jmMdB+9KR8B5iZw+Hq2jBNHoe
CiqEY7wxoYVmrYv12Vrz15M2ORjRZQfmeiVIT+QuntvcSaAntHV9aATdUpeObH9t
ofbM5Xc+iu52Uo0Hv0gRd45PqThCwMHL2uMEUZ0rzPMa6FngtAlSZPVhGuch7Ip4
Ly3ruge2FvV5QnToAFglgXhwaT4KdUn+rPs1aAZkkT1qndHaqnOUC+k+Tbe0n4bS
nSGWvJLUWI4CeufC+HSbU2+Cqxr6OE40dA9hzdJzXW/JzG+b0mBG84xLUG/HUMdA
JFxT1lCf1L/We5YZ1YJJvQW+RzC9dJxBDjwLKkMGXPjcnU2Ju+QTuv5bYI3zxhgo
p4pCa/pW5kZd1JE5Old1SbH+T3Z/hAp+GUiHxEUB8qL5mlgAu3EFhprWzJjb9Y3G
vhsLTaOeMnBTEhoC4hj4cHZOLMo12owttlRk1RAPi5A1qiTzZKcsSkKwlHMGsVpI
QtMSRA62+EJIvLOcJLhLRlwR1ABHCSM2CRe30L6ukBbCjX3b6bJjEqSbvmgAkMtg
/EAr/Z2jcagt5e96bvOXYAIdlHDdw6VKmkPAb0Dt8b4ccD30C27RpaJawzLZgS4f
O+vR9hfUt0xjId/AZgyRNNZUyJDFVi6oMTknpOcEEsX3RW/3H7L4pDe2JfInI5Mf
BjEjK0cWQLIMeN3WfT48yM1tvepD9gkGHk5rGmcj0vYEPUqSJFsh3nB96nhH9y6D
tvSl92ZwHTNBmtsNOkP/GdIBWGEAiC6G+8eDB0d7032PGpP7egayjXTrMLXBEuBW
g+h8Paq+tYaxGWLJWdNFn45WKk5aTcOKD9fNCTHuAQyFJKPQ7ohu5m+VL2tX7PgW
1K0wltK/S++2GIoH0H3NWVckHTmrDCcCHIuoFzCBOMwuJmLxLFbkkWdsgFAdrYU0
GoDs4+IGU1Y26x7j/u/p+JgY8vmds+9M65QNkLOwjdOiP5CSG7WQ+1uayKoWLSRx
dzlRiJogsu5Q9lrfOWu5ap2NRDiqK2QdPCvMhXsHagd5LiqsKVF8h3+Erin+ze4X
LL78NUMtx7EqX5AKdJLkLJqSSwiHs+TtTNRdDPhphgVF/iHhM74mVpJs6Ra5Qke9
BGkQeEWZMmyVeDkpJrG/usue6y/Bw5Iy2rbmnccuw8Ey/ZMXfhps9xjsqrx701NH
DMsoAd93KEoRRyIomLPv3cB/32mNi9cNJ0ZaDEX00bUwH+EbR4PKLtFZC2ku5ur/
11r1rskh0Gd9ffHv88VHHGiPKRY1B99xAR0Vkb4NJR1AQNmEwxAf3eZM9LBWByUS
/5CJrvFyBQ9RSw1BX73G+3vlHRtyoUPzMbmI0k99rkMoyg7eX5iRG37bP5ZEx3mV
dhCF5atwYjbyKKKRVG5zMr+FsX23mOMv/FXRqXfV3Pax49fh2p8X48C8kL2ucyj6
G52p+S4PqwrRVBW4PWuldUgjO6JC0ma0JD6tINKfDmj+795U9IH4uYlQODcWnyFy
Z/xjkDqr+dB01VIoTMzA/WfTh/+o1qGe4v0udhLtTEanoUW+UgDukKGPbeM3tE2s
UK4xm9up+Omrk19Tr+Trv3I6T5TKHur1LMMerwKBBsqqA/EtArsGsF5kUK+5uCSz
+hSY9R8GttUS4d7/DT7NfE5y0l1/vgacNvrc2SypN7BBlGgsZgPu/xsqe2zjt+hf
+dHcg/ly+aFW9exG/YcyOns6LFa13bg97xkIuEbP726hh/VCKwKQAE5+4Gk+G+xC
d8qIlybcgEDasQG+BatA6nUUr6ZYZ3Uzw9WIn5ZQKhjD901TwUxGxvg8NKqYhnqn
3GTdeMF1Knuy2WMu/g7QBPb0orm7l5nfwUeHTvOWW62XAs5kwYZeVLdE+/rxF00/
L38eMlCHwx/eLv7XBOwffxECcgYm6VWh0vdpkJYz1Bg3ueIMk/OYz6W3oP9RyqXH
KsdhYlsds0RCMhtPKghikD8q07BYPYYfn3jsIsZc1u6pFKLYpre+ISCPrf+lgswi
qAzUi4Px8K9tQjLVACHO6DLyMGl3b+yUOndXw64PxNGr2cK2FH7ikiQwJElWcsta
PmrZeuo+G9PHp+sBnTg4fzK2Yb9FXGG+VsVuGVlM1qEihu3/VqkCrsIjDfrwcbb8
S0awk1ZfrNDQ3/1XUWewR7v7JjROKOHsmWhjT6b00TpM27ly/DDmUIOloti+I3e6
UA7qybI+jRmxxteKnuI6lU/xUFVdb+n45WDGZEQBWssDQp5g7c+un5CAgiIDjNlM
SBYKh2Ou+8d+zrYgnNy/zXUUcQzzulAP5chp0hZA0OcL/0fvA0SPYJNHyF+m0bja
Lo7kJxZcQA8lDxqHV8Zpu/v+UMDtYlBRnGY0iwIyAimh6eto3eMuhXoohEHmzOvJ
2vsDHbOEb8oKIrfQNbkJBgfgeN5uA7JESUL11pisciBokyc7DD0EYfo8gL+qrDUx
8terCOHMnHAaP+ZqxqOBmvBaKZtoui3CHLdHPSt9x+cZGcwEhpQNaZrmwazXSfWE
soFfv7zFGUYOYhdi3YQM/sDniHbEeCIVUmweRysevAE/Rlr+S3E1wBP2WEW84AmO
du3FHMaHzcGtvupZy2xuOXu0u8RW1LL+Lhr7PnHk1T/FcUUEVwiDst1Napzse+XU
yMisUSG9N7+17nLaE/Qvx4O84Tq6mq3UW0JG+jpo/yqEJhf7bwax2/D8wPZQV+is
vqVecnTuMqsM1h/WdApzVnNZNh6nfdr+2B28Y1z1VJl0U+D5pvkurb8j9knT3ixU
JGV1vBSFs6WXbcVHmIashAEuSUdrI6YlsY5hjDVvHXDfETRYNPTQkgaiOSQZmIG5
eWCzs3FibnfInnraSlFrEuNXpnsVxqZTeYmq8BmG39Oha5fD5fba3eTdgPGmpR6d
q25mFodCPl6tMbPfWy0G38x6FjCyMctY5aO/h8BCAzo3XW7URI9dIfrB1C0pkc5z
mmwmC1j+IWSktz3h8YW4WRtdZVX4vM11AbeyzSMlg9DzyAfVgkoDOvJ9hZvMACb8
q9XWIF5GGJDfzWaQB2+rvFDPyGW9xCxuUcU3Gy+kOWeBKxYAErthuBeBw0DjITL8
Kwp9NA+As5FArKM1Kej5C7v0MlBGR7n8lMwJN3Nneaj21Rpp3E1Pj4LHSq9OFekT
WJrWBOS8F2FOnTPYZ+TNELT2U2/EbuugqnbkX3vT9wXjnUrsQYPX2qsVJ47CV7y8
bwmtoY1GyxgSSLHxeZQrNgKiNwWUi8sGU8s39+pA1JNSUCOuaml0FDjztZzN18pR
eB/EZnVop9UZ7JMPfs9VBkkfBRgspT0KMmLDeUvelfgFolW2ow789eznuilNTGOO
PWpIGNSopOV5JZVitW6NX544tHyHYQw4LXyxxgYtB2gJ2D/DaK19wuWL1b8LfLs4
a7YxewM+rAqBkLGnvnhXc5O8izAqrr3RDBfG8la+hbzgpgnZFuBeB/hzCD5na+Vp
YBbCXKd4YcLYa2iV4tEUtnk+FSfzLYgmWTO6saHh0jpQPkq5e/e4Fh55kafh81xw
/EJxxY61vKKcLL3PFZr0XDdLCt1P94RYsc5SzDXtPpw0xlsEe94lmL+PSNgMpkJJ
SPWRZTyrIkXUvijOfdYP8MAEgV0JshuTimaYBgrwK4XX0FkVg6/ck8j6gg+PbIs1
v6W+suTSeeB0e2kkjF2j4IVaJXu5OnCIA9bw1SqNZLKQtHLmY8SUwzgUg4pwfZXb
sBpfYJ3CMtyvp5aAm4OZQ7O+1euid1LPw1+9/YoLpuGkGNGix+wwSw+R0vIRv15i
NUbFLqMEiUeWcEVdXkV2A7XB4Qyce3rC5SnQSs2eu/1MwxVPBy/qIu1+s1Wvt5Pd
0Abha9rqteqaArHHvE7VfGWa+hYwcoNEoVJ7AtQ3Y2PecK31xyJ2Ao9UooJ4qPnS
YKGeVqJ0Ebx5oUsy1OKzELGf8MXv7j3XHXKk5WE+fVe0x5/G6ayv1fvbpsJInrCJ
KJxnmTqYEmi/aBDN4/6xBHJEzRE3y4UGrrw4zbaWFo/oIS2Gpbw5KxefST2jCd7W
oLmAYtRyrAeCr8hgmhtA3cvwfhM4VGVjJUFRFPRiTg5p2M3ARC71bRojZ+qdzb3E
HkkAFm15up7TYCNcfoSYyDngkSBGhMav1hCnDLpapmXSaLArPrqw1/FHUsTRkAxq
Tw6h3yfPyDxpnRram+umDBE8C3ut0X1BcT2pdZtGhOp/KA9jYBriIAaJdXZ1ZQ/h
AbSZiMUEo9eG7m/ds7z2lRymB2+lpZy3aDczBefP1J1tREX16KSWjrbyBpEkBqLh
xiCP+K28KZY3sr/RfQSjITv9PA0eFNVHKFd2cuO1NQF4iW+0G2nnWmBs5rFjiQPf
K0g3kcn3/SCMSqgWAQSTOpblLMtNIfpT9VRSuOD1X+IIyn+mgDl1qnp/jtxwHRMA
S6mWo5xVvYns83k8sYpHrWNVglVdRhIRBxYlFRXm05Q0OXwK7LRg/PDV5gpdPOkb
hUdSXfVNT7p3i7FOFu8GkyncjF1YuuqUPYkr4cQXerNDJ1QA+hrBpM5kpIgEPTdI
zN40qS1klqftop8zcGYqO5Xe5BKAdwqDFKvSSKaUvuzqb8VBmRmiWJsB9kKw95jx
0vJaG4E7KJlg3ZNGEfTkshcg788wHsBGaxvUKzEWpJEotWDpK5+VOYVwowoAnmhu
esjy4cXfRNsBeCL1ggXdQcYcEfXfscvN+Iwsb+CBLR1q9lMHxPC62HB844Sn3yYx
IiuMj68CvwWE/rxEIriaF0Y7/PgwUO2nsOXkwTyJW6D7oDT6ZGRthint3KDWBuz5
wagFQNttiKLEuilJOENjguqLfuz0LLSM4P152JPM9Dpgk/kkHtJxSIOE43AL271j
zX8afJpvkGZLCjjfCbyhAr+eYj+D0VzrNGlQ61kk2O7t19xZGw7BgQ2Kx8jrpRVb
K2WwYM6c7MnXIyU48ijLWXJs4+HOHGilAhjGkr6AxTfMaGyniOJ0GhTfEw1RNxUN
KR2naPJQYJ4QKvt5ee7Rsdv3obS/NfVHfF1yjPJwCbA/LvodwjD0hcIwiYIxyXaB
g44ymQ7O6s7uhmtpi8K31Wo1k7u19j4YktNJMCFhU0EHL/pjP0Xb0iugCazmAPxM
okvYvK5hcOrc1F4iMt8z7dag277rmvm92roxTxjKOXvU6Y8OaA0+/r3DD9xG+HL4
3cWAfCuUmBCUMtaDYm3Xgs0fzvk6b3l+PrHHryXhGtCtJnqTORPCdhPeoD7hcyZr
BhSioASAaFKH6oQj4bhxNizlENXCeZICSAjFcnc3NE8hP/XuKyNZdUOYz5JdHGr4
AY2tHmHWCSqFM24G3AJdTzGUmVXoV3vLJRXfjflYPGoGvRv33s9vMVuEPuCFZoIx
K7X0vsFjjiJAR+sv6sfye6vVXScLbDAAFtfQY+oHjR8Dj0BpjC/idiYeBv1shUGD
lSzkNNLzjtY5phsVkFZoweX5jrOj3/5MJI34MYdF8IJxiaK01M6ZpAZ3becGYa+w
pw6qAhk9FWgk4uXyF4A/yGL7yQC5w+r8X89expRV0UP9gz2Wy1dBujD5DvsvDuKX
380URkfXjUhAyEycXLF90Z6WlIknkL2uPTTKR+fHC4cp8NOlpan8cfDEwV4adLDB
lymtRth1FkDOUtcOJvy0rCMH+rhOc+8de338nnFXIkLCv5Cot7D1MA0FYemVfJsW
Wo9SQvgxo3hrs/45xGXAwF7PHxL4wQlE7nrYgMx2CV7dxVCJLmU6NisAFliFVjKQ
IZWX5OOY0t1uJmzLHvDFenmGa8/UU+ulYRn//u4iSOxg3ydOlp7hyWD/3gwkZ8kq
MDy6q9/nQz2VSVOrOV+iMglcn7gk8ZqUsbJ1rSXxjrueH29jdUVc1K1KacGDbdk9
toff+gL86LKW8PV8Dvtg/6jh4lVv39imcWQZYQ8QFBYlibWRmow1yh65u6qibXFe
cuXLg70oqiZEzGt03dPS+QgBIvddSpzGu1E0xH72dneNtCl2pocZ59ihhCcFIPPz
D0QTnDsoP3u+KaH79kVxN/6BcLxbN7VLa+AgVMPeSdIBviKE2RRtWZJEhQKFJ04Q
7HnpQBhyuy72K1nV+IHLH9wGGvmOtTB3azxuA91/Kq3/fi9tMdyhK6Z1rNZR3A7H
hx5x83O0UtsY3v92mVCQTdte5S/nzhlb99BbNhJCsVn/6+HQgY+aIJj9hiw8Mj4P
rdZRFPv42bcEWNZklk9vM6+Xg3rCPnNtDW4aiSpR3jfwnUWaIxZVhhzCeTkl0xFR
iQ4RJsXBA1sIXqkV4s7wYfcvUN/Uf7GY9EAjl5sd0qzRZqRBB6YB8Izd/CukDXnE
ZgvJbUJuFdziC3TBcAJ32rmH+d3WWHxx2qbrbdkOGbKFkV65v66U+SF7il5K1+bn
6/mm75r31KYOxeBkdzQl4O9rig6wPW1noHsvXTbb/9jiVajs5eyMPmTmkToLtCGi
aGvgWjKhqH3eFWTo4+Z3rZUvRZyOpfRhKUCOi1bn6+Tj6WvTCE1gEeMJOiobJU70
C9NIjxF8ZuWt9P21bLfuYWcAN+XGwg2e7klhFHSneAr/7nSUcflDdChSmoowPojQ
Bn2YupogXMS8GDYCHCpKPpTiWoclh7UY5uDBFCOrQye+fAFew1ygQ+IuiqtWiTar
2CWmb9kv8EdOn5ZrXI+cwPMKtPq13XWoSoMJM68vR/Z2o4jH2V2InZjfxvheCtoX
p4wUcyim4xr4uoQQ5/6YG6IThHuWGRrMyteOw8smRbXC++EuTPCNpJRVSsBMrsLh
Ef5pme9VTYC92O6KH9w1C5QVdP8ZIeJ/R48g/lDN+riUJcdOP24XZE9tddR4i+zV
3lB1hmkQuP8M/vX1GwYNALL/uMzlbimHGxVilnEZIBHg6Pu7njAEPAFr6qN6oVgl
0PDzfxzUsfIwnuJrZK2D+f4fjiyYH5FNy2j2sJaoDDWZAMBzDfDxiM7sRIvdBBjT
oZsFPD1E8Wfy3yXIvfpz6Gh3ntsCGyjULrhyP3LOSunOfdi/JpoJ7UJ+Ur8SrFgr
rNZE/diVAgKqmYmBL5pJH2FtaxKEOwCvGwx8c2B60P8BbRab91xnzHtKpVMMlCPF
xJzEU7ieCCrl1sGsWdhCEvVNOoo9pzylNqU1fN4/h5bCJoIWo45XGGM0JX8tcqUH
UMDLhjNhyHJzsYYnanrn7ZfmVcTw6eKokWE4lu/poecSIETm9itGYU1IIxEXscgz
10lw2A4FKWU7+vFbvLkW545nHa9scnjazUd0RhTtU9p4qIt3dlL5a5svtxej29Ly
WsFKQU0pJtc9KzBGkjKThLM5dSM7HpuMP4MgyL8JW8qBPj2mH5w83Z1Gl9A7gN8O
Od5BQiW/sa48sTTNsXpMWociIxx5g0XbKETIsE6QWQXkE9kbziJ178BBii1gq+qI
QtQyQxPq1KVq2UN/qwZ6lVctT6IlokgASCDY67/QRyYCX4HKdsL3qi4e0HB/TxVW
sImztUXxbwROrBQh4zg+Kpfpp5Q0z5DP/24/MiJEyRxgrsLtZpBFdcG1azyEVCP8
IKxpXzAejZuBVXZuTeiwxNcEyuC5cgoraDAxXaoS5b4RMiKk37rYPUXVqzcPzicd
ivn+OQ3MGXdAVm9ma3pDvCREyN/irL4CKXN+rioidKLZcurgaSwbDQE62Q/iklFl
hBi9F7ITx/+b4Bel+gtUws3VgJHHJw1jlmITafB8dVopBQyP1OcpCY5DqD+HVdA5
FXIsyXrRVPcIFvD5tL3bBNpKp6KetRNTHlgcF3dlUGJ1lHpwTTTAg3PwtXthVOB8
CSFTJwFZy6vvsExgn/sX4jYurqsyMXCKmlwcsan4ez7pvMDafgwHcMOH0+H/ujBk
iwp3ryaOUNR3hIroVvLlpBTvUZ2xAnA1Ls8G0eqjtHp9p3yYpXVF3s0uZppg21bD
f//INhJacYRFte56WQPNKMTs8IUvEX1QIB/HJadAmQxGHMnutNvkHB4XAJOlEYKv
CPXMKw51x3+uCMf9hA+fRa+6Woujm1LnkicxE6Nmu2mPTv0/T0G9K3r7SamGlJgI
+1vUH1OT4t2Uwnl23ONfdv5lFrBiGuuzUUJNq1kxmDY637nbXZQCyEnGFXsgnpVf
6/vdU5TtDAwnFs/kSXGViU7bPNwWJjUVY8PChSdwa8jteRPubxTOiT8nauVTgvdL
ABdTmfKna6VNX3QadeabZRhDkh+TApLhrcty6jhOF3G2Tn/ujj1qGwdM17ZpMQys
Vmp0zKJuIjDi86u//UVHR6b00jLI8VVlSgCUNHZXo97HznyT/CeR7C+LxKb4Jo+0
YUrHPyGK6u0V5/paxstYejpbpvcBjYBjt4FcWd7KBHyqDWrusuwQigEVBqvEf+xL
cAbp5Cl/DuuOEblVluAl4GiGbfR+ohSV9jIREDd+LM1RazhyIDrlQk/SvoB/PgnR
qNJ5YegzwX2Tel3vAe3Q5P9GmLg6OXunaBdKRiqWFHM7e8d1FxgVORmG6ztuSRqw
LDM6qE+XFTCIiE2FBf9cTX440tPrpZUJwCpo37ApXp9TM4UmTJxQxOzA37mtW7L6
d1oj7U6aGwhrrH9ppljUBagsmVwI5BKllPZOutAIKz44Dw3toDXpu/D/OW6bIjO1
Y+7O43cX871VCKRRn3oPi786s/POij0uNsqC/uYDLi+Ex6Y/yV/R28KoLoDqiGmB
Hawx71YhmCKiQ1lZloYtwMZgRgoaO9/AxJVECc5qLmIFjudoW0gj8PtshaY+LW0K
JWrCX53iGXbIY0NUAlVA1/WcfpCM7iHyRJTdp5quDFzAWKtX16XQZ0UjM0z4u/K/
2q8AGnh9u92og3SINw00yrky9xwMX88ae46Y+EhWS3rkfwOHmq6z/ITj+/JqyPHc
XEs4Qr9AmrRyg9Uvz8C2froZAqAFK/I8VQUI9ZJsrVChGp4p1lHh4K7hL47Zr6GI
kEPc2WnMjgJBQAIHO4U6bPIV+ck0yn1m/F5BwD8dGyDiJsDkkO0/NMkw53tvgjkA
fySY/N4YR6VLZkHJeebBS7OjBgamAIOuFt4t09qnRwCGAz/kTaYy2Uj2DDUHma0s
5q+ipuVsfBRgyPNRfWTQVV/r631oqb7Gw19ys81AJn75Lh8N4gGBzRh3kyoi+U8c
fYOMgvGnClphtJY4csc6esMea9NCRqRp3a/EC1NHAoCaOB2ONKT2PHvyIHzf3byZ
Qft3m3gqo5jF1C7QMUiTO1NhA5M21rhV1ZSOIRcPKQP0Rg8tAVq6GjABc6FsxVqu
7xNu75pVgSNuPgv2o4e7RBf6NinrYYNv+1dIz4jefGoBtSsHUTQa9XMoEMYXvcXW
T8xN13sJ2VcJAC2rJexIlcPqZtVdl/h4Ogxb0LnuWJ7ODBWlmiPY4qh4DlPpeBT5
W+X3JQTqDwHor1ELAfVBtpJP/ReO3Tbh2la1hNBmHf/+fTLkEGngSrdZaKusLnrf
3/J5QH0TxSv3KCi0ut57o6dnkhmBKNVG06MCbEIa73JX1UvXrUa8PnFq+WglksiE
5Sy0gsT+WNuZLmB3YwfiKLeQ3Aqb6vLs9ykLwGjFo/jAj2AZ1cAOm44asXnA9MNg
YyYVHPrWUXOS6F3Y/h6tmLm7PMsnaAZv/lhihWnhPnl1qcAa0d7SWCpTGoJtpODE
SEfF+J4GLKb9oWiXlCdoKqqF5OkTqJl/OIKTb7pcS/K8YfV4mx7y7KOstNP54uZq
eE0KuEeI3Jm4YwSnLTSsE7pVzmGHB9H3sl3t7SIhh2Qryk9ySYgD0mEZq75hemHv
Iq+pJx8J7afujR/6gwkAB+V9M3qE0HUF2gP+AgkIrE0eLxwY1VMcOhU1J3+OOhzx
wQHU8auUT0RyrhTMmHSDMwlK+iSV9CrA42+wcEz2KKYfHKLv2EJqQovC12EI4I73
9RQQJBRDDFxD2RZ2VVgdgDH8o/7m4iTp5ZSoSMPDhrOn5iCoyZxnl0rc05W5YgRd
RhiF8WhGwLH/u6+DDjf+5rOmoD2jSzecrH9mVjpaK7ftOOTZLfXjoWxLEl07aLho
OAwe43P+DkoMiHboY2iLwqy9rF2/e6w+raPdEYXCSk+dL/vQq8sHnxItJXrXEUAU
JfR4qRHzcjLl/XpbISD6HxIoCVM90CJUSjts2Uxwfwm48hbE3ocX0SLt9mxe6LZF
HpkNtufIMIkEOkKRqB8IA3xI5ghMtA2s2v08ocI7d3pOnRSfO27NrV18kfvPQH3Y
PbsTiIiegngZfgAlSqvp+gYk6rVW9liDBPQFIIgm/gyukDwNbHfQKUopXGPi8lx8
cKkGxGO6TdtMeX0lHN9BvZUFcm0cy8w5xdKAWnobGwtMLVq87HsK+ZvLq2CEIe/s
8aTciFHb4EkGsY6Nly22anFL1YCJd6tQMgD1VlRmP9I0h8PTel4FYmqxe1VSCtnD
btdhpQaQuqi0CCZq1dbS+0N5akFQJwfTzXxFNjzuK0Kba2BoR/AsiJZUBWvQ5oEi
8iEUQyggfgGjP6NIooAs9Qk93FKB5qdIXTGv6MCuZqxmidC8dRYJxDk/dP4A9edd
fKC8YFXtzGQgn1RDgAIvigQGI3qURLGySF8osl/3BehY9n5u+JBDlIa+Hq8ZeQIR
9dfGRxv+DRtL1F1PXUnLB4OWcO9cn7pIHWhINS3SPXjFWYrHDgFDKD2X2jWHzJWL
dDxTGfKLYThpVWzkK7CF8WeJd2YJbZcj0/qyi8dLdIwTOp977Hs0r+Ly385Btm5l
galbgt3QXK0h53qgVRJ7Gl3LELVP2OFh3BTk2RBp2D0WxmKWI0szI/IA3H9FJNul
XtCRd3R4olmxIwX0TsOriho897CsGFsb8TPHMV7Rdz1KigjiAlEemgXEqxc/zj//
P+mXxQ7B8gPA7MSXkfggucMgPJ576hAEW1sLQsSF0vTM67sxPzzRY/c4A3EkdTiA
5zriUT9SR8H4wst1N/kcVLGilOlBskB0rexXMZcxGBlbp8/HqNLdBjvoAorP5RXy
NZra47DXyIoC/qq46td2xtLZIm6L+cHpyiiaQuYfXb/odP2CvnM7e2ALzwGwQ48u
rZNKvhjF/b7N9wEdC72+rj+rCdhNNZjJO8xD3EtBGWSjF3Zaf8YG6gMEJloLX+2A
mja2t1/Y6zKegb6+4VY1CVcrxLcXidiBUxgDEQjyc3FfZ9kvQcK5YqQAduHuz46D
+QERmEezCo7JxQbORQe718m8n+zMZmI7Ib1RuIBTUlsGYtid7aL65niwzDcndhjN
KZagOzwPpWWiYxfEDjn8yrfKy2kKFaRN+htILwDMcLqq4WWK+I4Xy+lmZ2XUkNG0
zTTrdY+c5qXLKuKrgOHtQia5u3OVDE0MHfYyxUGmT7J5g/8GMuHlk7IUH/FFJNdl
O+RQ6M9f3VCkuNq0iK/QP2pgHUsv4jedH+LUcSJTZqki+fTUeakWznALI+am3eHe
ClyoByMBe4uq6roC0nmMp/KQoRJx6lbNsIa1YI8I9soB6U77Goktnaq/LH/G10qj
oeUcbU9HCM2x7TyKx04B0TYlXyglDI81cESYGD+R2O7Ol9Ma7h10Z27JFcRR/d/9
dreilHVHyxW0zuBJYZiccx6OAZgRVS3leimfcv2A/+EzVDX/2oa3DFVLyKrsXql0
UVXbiNpYvPfEqaECXL1IsZuj/VRJi2wwO0dlV7s3I374tUF+Vu4H/Y8GArp26Y/U
hGWp+tGfzhnqX51II0yRTQ5FCjilD6xsT/nrk3NvC7YrefTeyQQDTLDjGnmbaD6k
7lKAQoOhfKIR5HwTbmsFZrzKB86PKv7iKVMSW3v6HftmlI4/6HbfdcdJXLpT2Rsg
5t11iEGrxq0Wcftn/9bom//eOWAy047T3NjGop0v7yVOAGMHeKBqYkrEem4Kgf6t
NmQQtQTvjq8t5TQhTNva7ZFrj8+u8cYUmNWzj4I6FxPl2jID4FVYb84z2DIJ2egm
LvWf2h5pAu/E+e/eN3tGgY7G6qmaKyOCxLWvzzvg6ksta/QP39yjWcQex6+v1nT2
noxh69QtfT2kPAHDrjz8EJ9vy4bgs3g/BnSNP6ttWmESfL6U5Vhmrr40ykgTmldR
dwY0HqdpDl0csS8qU8zYbO4vX9CIxrYSUFQQxM+8QIQHnDjAauLBqlXk53EE4vBI
1kVQY6Uzwi3uhRc8uRTdKNtJPRaJGVfU8h7uCN11VYhv8z0xWe8rX6cJRIXF2ans
G4LNHdIUs1USKiiqPaxtfXu4b8iIOoqsR0Y9kPSqF7okVyUbS/VFlqxTBk9UqHay
MG4WjgkPS71agw/d6gUB7I2hL+zhPCcuUwrfIFXtwruZMm7PN8m8vNq4PunEwnRa
ngPFuPC5nSj32MA0tN/CFMrHIGWOQelkRqb0m9lwdY4PgEATZYNHeTRTgENtASls
n44YVFFfh+0vfh2N6vkPgmajIq6qK1XhZ86xc0GCbgVcdzcnnMP/v3tM5LOT9cQJ
OpGl8xearOt/4zm0idq7hvnirWnlW21PlNeLdi31XVR6ve12DC0Yz2CaZ9M8nHLi
5tQ2fhBSjEk5+6Yrqd2mNsVE2Y99m6NR+qu2q1C9zqR08mBh1hB0DafeZE89LifY
FWJHJNmVJFdQjwl6MciYqmeCw5YBL2g36BNqkQUSxF6dfBZE01rzN31qw9XtickT
FjRTEDB3oeYIsIqRDFYfYzexnu2okVyVscVM3wmaYwS4a309mGAni1RllZ71sRuM
ZzCMjSIEI5IJlXKgRGXNTIludKjWzKVgc181++NEKpiNJFQXJAKMTLmozRkw61lZ
qq32VXBnTJrUI490POZTtJtq/EdqEZRdUaZfBL3D4E9lUDLcP6cB0fO+NW2hiI9Z
hpPkT+kq7UHxMjM7G8973fwxmgRQF12hEbEjvNCjQX/GiurHXriIoTeVdXtPf6YJ
xUKFIDe6esea+lBasIDVe9pb/+oDE9rnvxmw0OyDutpDbMydhnoc+krrAU1AdLG8
H/s2Aez/xI8wCK3XADjzBDE6NA7AERMa1bJMAbHA5qvGbmn8NQeOyBbFoLc6Lu3M
Ju6uLJpDc2AmbKoqDa+tEP6h2ZHcFH/6UeOlsw8RGvXCWo6JbrLpmi1RYtiK1GTp
Bdhnpl4shJZS1xk9+qr8hU88KM2MEvEQcwsc2cRFXw0HmVhZqlKjFwfWs5spZ5Da
Yt8fBJRYHcP6ioxTmmo5mu3hxxvzapFBHfiRtvKgDgu4/+CXlzo8Wj8XlVuUNQdl
Zs5X2O7VBRfSUZ1qCzg76WtXxbnjujrnCBnTRW+cb1ScWr26ycRaTD8gAIiL/Uyf
2A0uwzQI48FrJBSXc1vCRuZ54d1WLq6pZNwwr2vya9SeUYpUEIN1CpOITjvA9Uhw
fz0tJrejCrxuCDYDN8beUubDEWlbxkU7T3QgjyuiF3Rd0Fm8UX5BsdR5Fn/ecl08
8uru7maTk8V1gHhahkYjoEvhpTsQRlSzOLqixaVKRkgAtZICPrIYJU/JYL+Jvgg6
hx5cgbR4Sj+NygClaY7iSsZUOnHikDQoMA3/JSosOR4YKy8JoLUQg30QzE04krDk
T+cbUsdHy7l3QrmVDbooftbfjbEd11iz+GUAnf/SodPFuDL0bOjkeAQoIsZeLbRt
nSuLLoyo1a+aS2y3oonQBNqmltn6t5bZLwxUxAnywq5n2Cew/aX1fFsYCsIGs2Iu
EXqetPV4JQJluNZLm9KSWeKjJpdA1BbGcVlrTNocjcxWcbfM4SpL7962aXdaVZGO
6Av3cX2YUBc/8W3UHyTNe32mmQ5n/b9aOfNFmRZ/Ro1K/fSe1zp4TCLgK/6SBcp6
19x4BZyWS/lUw/KB9H+b7wynNh3U0ASB4xN2XD469JNHusNumV9b+FxiKzsfgj7x
YHvWwa4+gffr3cFVIZ+Qa0C7VGqOeLU5XTyQbtcZwRgjb85hyzcOqgnTFH/Drpoc
zPmAjaFJiEPDJmqCL/QFtV5w8s79pbk138j23CQoQnhIc30MhdveRpcJw01E2cqg
Qh9mctm7EUhy+7w3+LoKK1qJdwgrDiM3x9zUwipBlgUr32yDssJ3ueIyANtF/49/
jONXoI7qtM3y2IYfk+muru2GYPASe5CzgGBh0BUhngB1u8y2twpLchyWdJWrpsgX
ZKRXTXgvukt6JWkJah/ap77KYiZhUsAiQG6km5l6AemSOYprrOzsWtzt6bsmOEdQ
BVZqsQNeheE6whSAzMnkBLZr/QLTtKZoTjUzK8XPFXGeNkbDUeP9YJz5n6GPebbu
Ja0VcqsY+yGtEclUS7TD0uXLjvHP3H228YK1suUFdLUVS9bIKP9pHja3Gh+SkKzu
OYQJ+VmfaBQKEpYG54hE5jkBPRlVXdwWDCeb0+cw/gTP+X70B0P0U44wxVtCdnzR
aBufZ4EdDxDpm1uwXmydp1klMttb3St8RA/B3nTSJnfI4q2a22+U5ik7/cYLQZQP
07Eo5gz0StJXMhJv5J9/+GsS1peFQcyx2I434q9fA+VLvOo7PNq/KKm0dWh3XDZp
LFIQDUPi0677BFu2UoO5nKiNoq/m/3CVlgWH74eIM08CBB0p3307QrZ/+ivSYaOz
FKSor7pT5xubmqsvmyJQmhJKS1bO/TFhRNYz4OB2v/FQCgZn6pD9eUU1LV6xzozz
R4HzIdrbMVwA2GXJYa6uf6ajkJ2qn6DOkEThFN5IdEmvv2cpxPQwh5v52kUNz7TO
HUBrGeJxuRjdokcDiRdLttxPWVMKqH8Uv5nVOfEg/TiJMnp4wOtddaSr66TLkgV8
M0Q9tlbe6pocQoVVydKcsAddk0pgJgihw05265AggYCe2W0OvXz/6VV8fEAAc/a3
jmrtvpZuh0F4bGn8IciDxTKsbXpVZISHNFlKzFuZfQNnSFHSbrBqxHBPh8MkRx40
oHQVWNNiksmR7hREx7ubH9MXLOzmzDMsS3MbFl6UkEoEMl7djOb3IDh6f+2g7qXN
Gd0s8/t+f6sarT5Vl8TFpZyovx4k3sx900Gis043dYXnU0//23VlsBcdSXFs4+X0
uCtRqOq60QTG1vjiAQqSjLWDWkJaN7ZqaNs38BgFQnBJxwIoVPckK70s2eZ0aS6g
viO0HD5LkjoqW8xxt1j4YS5ygBJIaAtQvfA12roGaXNJs9pZe+i8Hemp1ZbngjWR
A/iLpzd0qx5rE6mXfiKI+FrAscKBFKg+1Su0BB5m0ALHQjsfkonSI/kywP77tXkI
G5ddWPncR+Z/m5cWYXFXgwQH0OkiKMtlEM/oxUo41NqqYggEH/5o4lyMKIjmMw9u
Mm3wTTGp3bTOi7Ja8SFsi8nJXPV50RsxV5RoHHqabEjDFUTUmGDC/f42OCRsZQuP
g7dYYFnkwjkCTmu4rt7aswG+x1H/ofQ8mqK8oTIJqNiWrbvJwsr+CF9etF97Q9H+
Abgu066ciK5lgsWaNi/Ga9O2YmL3/XLZwpYUcRIm7k3p8so5A26tPdxtoDBws1Nz
K4c6ly5KC8MgE5ZL2zaHDyV+sghyyaxzeJqnMNJbzAH5SNJCRWLoA1oiQv9lBVF1
u1bbNn3VT6TXPTVr4F0nfr1YiAl6r34Rxn4+mkbNIWacrSlbp8s/X9rWtDXevRxY
RgM6t2yITO/LmvKznmNl/MBk/2liCCHYFzPEspoGYCoZER3YfYaD9dZ4Wrh9aLNk
l4G2nuOfRBjz5Tpcdbdt0M1NGfSYri2JajMN4TczIuCoHHvpQPfa7j7ggUeuhrjn
YK+HQcvCVcLQ7ovGwH3YXKsbi5klx7JIJ61wNi5OBuKFzB7Nbvtwe/GXHNSg1k3P
HZ3Hdda8yFfMukhAvj4g3VJwtmpOj2jIek4QcUOasDrPs47581Ihb4X7LzrP05L8
XQWjfEPWdUiAb2/3z8BL6NewkkCwJD3QI1ae95jzLNqBLYdl7V3wMb1FXs+F01Fi
MxwzaNyu2s+OEgMSt8DkvADPLPFv2ajYIZh0vJ/LhEs/8HxXWpf96UIrxQbtKzN3
rfyrDDCFxj2RBI2GTeoW/+ixv/QRLtsg4ZJuK7vkc8WhAOl18gS0+7DROvdWwBng
dJIQ6EV85XrGwfjX8w9U8HF++uIWJd+U3lu+G+RdeQy0HgfJPRrXJFAHsxD8bkvw
q0l5NgsfGdSPn1rU1lBQ5PN1uTtTvcAbGP2Pp6B3MMqNV5ehHGarM9668X3ddkmY
sQ/P+agS9So17qL1d4NHOwhsOwTyCzIQce+FZ1Wu8Nodo4frFK27ztXJ6YLTD2SF
pAVRaQBG6/HB6YKmH4CB1IIUniIV9Qa0XVi66KUbjJNgiZP/O6Gi8HkQ/Nv+5097
n3m77o8ExPYsDjbLyo45DdNherARZ92UG+Fc9dI0jVziB6ErnqnqTdGZLwwwQgRA
aF7U19c/8ooUFtVFqUuzXa7T9uauqVis4l/LYd3TrEQFcfYjmqsvFIOYFl0czhVN
K9Rmh6FBEy7C9F6h5veWd/68zwJSUb0M6Cq+d3cMvkiYpzac3aADWeoeDGVHv6gs
/r5qwcIB1nWeLJTve06P5p/OZe4te6S18VvfhlolBDHA3px+YxtM7ZvWoj7h0Dh4
5uLREc5hPLXQR5WsCbeECBCCxti1KbqHtaIJ86DT4DlaQ0/qe+zni8huBBlEsPwc
8xaR+S1rg0OCUNlOf//Es6Kuj8EdHDsR2EoZjwZyWV7Z87ATLgGSsGivZx9KG5Em
W9C4TVVlwZufeLi1Y8yPIDEhfSm2l3rmYs2aeYD5sSESo7SWjsVpaOnLweyw4TJz
dW4p5EbmmExKfGC93mWfMYFhbkD0MA+tMb+M6MHKGlhwZRkiJ4FOfdbWi1kS8tpr
5qjNFB/Rbx5NsjXNNMTJ06k4mxWcc3AIeqC1HTTjbPmx58J+PUzSGoubhSv6gMjq
sgsn2zbKAeTbnmySjdLGW7Uc1NJCvxFNdRR4ykjrc+GJUm24YwNRNW0vZjP1F/Eo
b0vF4EXizAi1WOlstxL7VZvUZ+coJXxoNxQqbQ745vw6ciCp0EEVXoMEaXRa5YiH
D454+YCS0evFcSdV9Ox2QjHIHSt13q8I2zU9C7itEmGbq3brtEIED3887BMSs/rs
j8kR0vlfLwn206+S7baMmV3pJpzUzrFQo54CCLgoL2dfmcdMKOWjnmbp3ovDaWNC
cYTv7i7hloS8hzyKdZjaUFLD1DvhRerSS7TFS1sGlyquZVvnENjd5QOx/rrQWeJa
HoVKiYf7HYh5IcMS2UuIjRzIqqNP854Kz5uwbd5+lCax97Omk5xigFL6AHhSUa4h
Gw9V0LkIrQMiKzikdVB2pXZfCatBHAYYhcfWH+mtFV8ki8aPP8+gDRijqcMUApcW
X/ykhCE8CbftQByBCBW4FWb8irUfP2iRf6cp5+QYcSoPKuor91kUlu3w7+MKKQyE
x/7NM6m2cJ7gvvO7xXKRtKEdsTzOwx8vxB0oOgoza0ordCAYbUUl4o1ctafhLKQK
b+uC2AI0ehqBNAzkQH+aMemcM3+a3XMXb3U30gP+ykFmjGqlPlo50Swzeo4LXhrz
MBGuSerzT3caRafc4I410c93GNZ0Gd07/wcfg/l3aqm9R8aIaoCK2neaSQcmFalA
m5hfEGmK+htbhBe7AOPzBKBn+K7hCrS/ug6f5wcai5wyOYvwsCmQHliMXKpn8OTV
c1Wc8+jw6/B3ZoQMDVi2Ls4J1A+PAWd54iDRu3MksR9rH5MJ5ceyDH3isIvjoZTI
C5/M0g4nmmP68VT8GQwcF3wPIS3OHU7MpYDwvoYE2hinH1OsiVBwUj6h4yoAGkbx
ZE4kGLOOqpIuKCGlWC5N+3ivPx5/chb9bYCLQWRGfXegEYxdEWvVivMHULTbLmX+
26tKXai7Z72ujBLwOB96s0YZ7Ek8nBNf61eYqTMLeYfhX7rt4ZKxCkPlfcqY6pWu
+hb2P/bp7QPyvULtxTB6tB1qZ36jrHzFtBCijRslVX+lDYfp3B6yY4ayeo1N7j1I
/WoWivay9UtMcXngn2IUhfSpzzDsQ8wxVqE6jB5/XdFyONpyPFcIVj3O+pgD4z89
/1vFtxIeCw8D/z7legF9LXHDC6Kt6Thp/NzQ004T+gP7RccwbcvsDZ4Fjv/5fnXn
n7BhyM93vTRlZvAatwHwZ9l9bTNSA9ctboJdhyc+qpnvtQaWfKLSFfOn1E9/Tkq6
mQj8kGKg2/Ihl7im8M+xL5gk0of22vFYS/K+WIs9Csk2jQMyD30PLtkG/D2eN8j3
ASSGucB6/QR764tmADOxIir9WgepPneucUl8rZAIgEh2xbhhjW2Ms6eykMZMU2O9
A8jjXbXf6O8ADc+LFhuiBvAVNa/I8j7kTW3oczT9OXyeXdyTQpXS68zroKnCv4Gy
K5kz2gllwJAEgMWjH2PBvLksNqdvC8l1B3pEbzRs5udtNgzRI9+qb1zUb/nGinOk
C6QjMA51E2M4Yzpv3VpnFTlhbaTETtvYTuBvk3psifBQUZ9VdV4b4bF007ULBfxQ
Ez/2AGNdx833gNgJVIsuPU/64sNJmah0Mt9gQzIqxSUmHICHj/ehv2Sz4HcrHxqh
+INjXErk3Z98IBBugsPOzVoxt1IiKEizyDm458vHhN3G4rzDyLzD01cl6GbL8gjK
wE9Rl16uofm9YNAcb/+ZUdVDXxyaAVcNq+tU35d0dAcchoiSLlSat6huu9Op2sCI
Z7BibPUvEHNuYFlaXt83ld79SDDSVNtQtnzOmetFJrFevmERyF233rST/MZ22j0F
grj5o2JPsDr0eBKm3ZE//IwuWUuXxQeUg7jlG/RcSAAVARcK7aN0up23onoJ+9Tb
olqfAPG+6DPd7Hu+XpHA/qSs/dKC0+li3NmiGyX72eeILNHwmqYVSvYN5WGUwsOT
TK7GTSF0PNTzhBydCMisF/9bJmjg4KxbxDIuLGoQC66yhn5/oOtHEnesURoagHD0
oG1vTtcQRUOMA5MJ5dybCDrzXMyFRXRXPKjA3SpQJAmFsFSbU4PjPPCpyJv9YSmu
loSEoPHxlr9V9N0MVm5g+G+IfziLnIo/nSxDd1lyuasNLh4PU0XQCjOEJz8uafCU
DWKu7zqiDMYEpeOUpDeLiyTKVvpvrOzxYLwo/rSO8hAFqk4BBsgBuxZgRbPkoSp0
jPYL5HOHY8HwwIm5LcfQVYhsGJIl/dSP8ZNhIZqG+rZJpdZhBI+dzV5Qhr28zL5I
nk7HFe0Z2ivAXl8mAY27qOT5Mpba274NU+uRIKK0pL+QeBHYDZpRZxj0LP91BhTk
nC0LAclov6CnVh2a0rCH4dNfiV+PFhGt5uNIXUQr+ZnWCcbCiZSIwXnqC95+9qTe
5IiEZCGOSbiw53sZSlQ9T9VMzNoHiPsZ1duH0bmIhYfNaqGaz5cNMlyzAxVifva2
Qdia2Xpn1NFDIgnZEKi5m2ZGHD/ntZcylpTayT2r6irlJkC9TO3BX6jgQ7r0F/rz
b8R+7XT+dawRwD3QlpQ6XHzCcW2qd9AP07gRQKgJyzMpBZeQRbVyNgePFZkuBui2
m/MnKwloK/aN1ZXDNFQlePNbl//XhUz8ZU3kYiojLZrRpH/LQE6y6b/U0X5VEZhz
vhxseS29c4wfnE8ZerAbHLYdtUwuGbaetgoblydSwGNEw9m9g+KHUkGpdUAoEaWX
9uJ4MavXgUsfPL+8VlQADVmHucTvu7zSJo+dnqJ1lrPVu4VSCcbGv4zJvdlT21YT
75pDHQhaFlzUoS1zRndR0EwSzBYGKIB1ez6jTKy/jZpFtrYRSm1PU1AbjD65NVSL
lXT7M6t7wIYygIXQOkHuANHlzpJo4A46iu3ziwa1YLJYIoyEgmdu802/B5YYgTMq
QicA6hReX5GfBEEnQ/kMvppJGh+ddBe7toT4ODAIgHkkkueF7YtwsTuRaCrTBxMb
Smm3KG0Md5T+3u4aH2rCSX73IpFpLi4mCdAZAILPB2RKjsqG655XcJ58I4IGjjM7
BxKrAfgnFKCoQhmfNQ1vn03QHbbgyJ+INwOHJqKpARcnB5tXTsqliqI5Buwsf4R/
umpb2d/CCSpXfYaqpcFWXX09x9qBBu+oUobydX7Z37S7T07if8cQN3zk8CHo6Lxj
N+nvBaxg2aH73kAicWou5PQZxwDUDqnuR76cemOJmPrH6yX1Zpjo4ZKAy8x1uPCY
pWeA5Gr/kgj8uDnGiktLPIIyLPKefsdW/rq0nI5L2xO0TnXkPBproaKvgF/tlv6A
C6LD9V3hNZuKdrpiwrOMixWQfbH/8QaMom7Da3Pn77Lgg07hV8lEtPKKN5rARFQI
a36FAQnUTPwY6V4m6WXcv0AkuXORNtHZIO/yVyK/dJOalXjWY8UdlXn18qnMx1Ez
wK6kFEGENcYG+6dldgQkVOzGUWl8jRnJqg8Y/ZpF9gNTW71e6Cv5tmx1xH4SqnKV
kXDmt43TzM97Juu9w86WXJzvZAxkAALfDAAKNJO1ZVxDNR0M1dncXvtfvc41Eet8
HyRwvqZK1VBF2fytlBG/D8Xl825rwyKoTls9msWkWOTuWsz5WzigYmjfon2K8+Ve
r54WmgK1FwlXXQMu7sNNUN0xktgcHYsxMr5QkDWblXYx+tM2P2IKsiODG+yZvZP6
o7yzJutDENjrYZ3GluNSQfkIEBIv8pu/grQnqRNuydfCgfe2pkWZLrscsgYIIFS6
g1ju2fCaN6wK+NBvMZVSof0DIiCcgSzRasQUdW2aRWd9LrB2af8tBgTyh6BC/Q/h
nlHgVoK18gAOY1Tp+fLktO7dwbWrMqWw820Qso4L5B5uvmOKHd3az8SZ/4KxnZ4U
e8rEAK/4vlyIKhgiF9zfPuQBR7dwYoZYZ4Qrk9b2HLewOh5gjNP0qq4dTlxe3G8d
Oahu05uA/mw5Q09OikkZG0M6ycHeJTmvXQsMw+BG9485NF8PFPGRxQ+F0pRboxW4
YP1rTSc/9tyA+nuyyEtb5eH+FIb2exV70FqcDz8i79AxN+2jnPPV7kda1sqxJ+Qb
V7nufngqMISM8RJTCmvUTqy5kJsDmW06e72o0uotsjjDaO7yBCN7ivy4TdbbOHw6
fyMQoQ+SG252zQ3GtEW/SNjwLEh4VkJgcclQdII8hAHLMXgF7OJv+LEwMQYvsime
6GgUgO0zbmzpWvPxOKjukszOLikqi3N+FA6VSIrNMzXYiLXZFGQzwUAbOM5GhnTr
4d7sNMA2kbFx+Yx48L4eVT0O+Zilpuk8HwhfY9YlxjuISTsPs+irrPOiaQngej8Z
0LBH2Z2rEy/JIJJtXxN0zNSSIzyGbcK/7hAafOHbKqHrnqzDQ+urOFerq+cvrAQm
kd2tMGP+bx837BEj3yWKBN2z2nD4ItnW9sDcUrT3vrjpJUIM86CbvKJIUW+3ZLku
uJRW2pvRzayKbltGOIwXhOLpCi8D/SjDstDcpZCRIQ6oiA8iYtPFG9uOLrmQ+k6F
mUHml7N+ETLG5pbLzqi2cRqO6pr68+lDrTokbTF1jSY8YNgJ/bawjIXWUNze3RsV
mcW4MYdJUFbJ6gZxsVa+I8pQ5blHYlrfip7LsDng2NJC+3AD/TsvjM1269czZkeX
MKAIi3aLC7Vo1XXsVZ2FlzPaqTKz7jJsEo5oNt1OmCOFftfkfZWs2uWwjNLVR5ur
xruY87lEEo93CCpFb44v1FBrRveJXop6fYbNq4vePwGHJGStEICbXH+VdIwibReY
/VYGmAHYUqJcfHUDupy9LhgqZKX/m51+qtxGyNTqssZYpLyzPm6QuwcjVdX5w4pL
XGE1azStHn5W2MiMnpovcVFLEBcXagow/iqHew6F8GvsNeHsU9doVkfBuDosvdE/
dNMhj3cim+Hn/tOFavDdXXo1/8Ttc0r01+73+5xIPc1iYVkK8FZOLVhUwZEW20Ub
Waux0WFqJPFixK3m6Ve9l5bR40yeQUBDc3LXBC6jwiA1okj8cpNQp+prrbyUKqMg
nvw2AHn1BLgU0YjBfbjt0eKw7sEtNoPXyS0TQf/4NuKHxj9XgIBRkvf9Re16/nHL
sC9cvVaXg0ucupgB4qe0jZHt4QddrpGDAIi1XTVc2iRNvup2DK+XlX2r5QQDKGCv
Fy93AhFs+29QearHlkSt/FLp6WFFVUO8XAcRlbXLl1BbTX3uTyCKS8ssgQhtteJU
gt5MIx+1r33UB6RhH/EQ5q+p7oMLqH9II0XJeB4MRY81i621lfpOX1xhBUc68xIE
k+lSqyL21ALwmfnNceeshwDrZpI8qjlbvaR3aeZZhhL4UEW5pG0DVvRIzA854kFa
kLae+GfFXOPgnWROSlxpuRf+Y9Sst00Yh59ZiVQkERidp1T1TBLUZgQGlYOFF+Ib
azvMlwiBjyi81sG3jOoKSuSX1u4Qa2/dE9Ww7CeftFxqRph6VRtqdiUe51gVqLn8
nUkXmFIA5AngaQKeuzOgN7KGPgT3+lg7yyZUDX52322cXn4hyrAHlRzFeODhJKfS
5Ur5zbqnbE6QvrCJLysENtDipVqmzqCCpwvCEHVOEGCDJvdlgmHqrjCwMH1QfsTM
uoS5tGH1q9rsOEeQbFtRuq+Kf9cSsWxMYXxrpxmP8YBzH5slxp17xxEhz/4pZ0MB
VLdr72ANM4lUE5En1thsgkbiKzeBi5cOQMnzrN7uAHPxtQqhrCWLtBSA7GjpSEHp
AG26Y8HRreZsQpvXVWEM4QNL4EzTS3k7NrAXD5R4pHnSigSvBLVmvgps+hYzKKqa
FLBiEA6zDSbsJKfxKTLL064pC/GqQy2GPxX6VVUKylM2+Dhmk5Gx3uzDo1sAWLhK
yPHxCl2qiEPc5OPLDhDg3Wkozh5AwQt+GVHfheFX04EYY225az0jNW32Q4jpr8dK
8ef++Z3i0Jb6LF0/EmmNVEvKS4/n7d1uM9bLfugQ6LR6sfBBaWe5kENe5rPcDfFy
5a+ed5ELh1GF1Znu1YQqu39jhcKnnL2p97ifQq7jcOhaxkX5muaGm9Lt68oEItZf
iRnLwAihBm+Os0jQcck9J5ninQmuuY64SNv5RMecXywNfpyaLcvq/hxyuRb/5fW6
+ChZ08V+Q9z5qJJHl1kxKmqzcP55uefiS48mKEO5djZ49VNhIOK5IzkW9uHKKo2J
4GIkQdeA2wMTrx9qJJnY4spxJVvxhOZyW5yt6v5WBoNfGhPdg1pXeqs/djBmbIeA
sA7QuEA/PDsET955qY7M1zHwXT1aAY4r0M8/4Itaf85haQScXylHQ3q8Kp7aqFtL
Ym4R45UFkONNEGIizxap7wDBOHS0JuWwjHlJQ3Ogu2m/SKJnTcRn8JvjcI5OyPTu
s0BIw6OD975DANuXygmGbCSmFGVrPpqCVZvztZRhJcW8KAuYNOmGYmqDQctrE6gr
rm5qEBXMNpId3VhqdXR0sG9AQhspg92ARtB4PfNzEA/cv7/z3UEamIU3q3Gd5BMm
7jhwxQK25ycSSUMKaWdnPBJvR7XoYyebsnUzDJAFhQ4k0QpmfDPDqrRDDOPfFNu8
1DW+fYL4v9EQQVRy4YWa6RdGYnNJSBMMaUYNmPMPuXxlU4/5NCnr+JeOkk3byiAv
kvYqyNsts5Dmu0/v1stkdbMh/QIfmByy42fj1Dcf63+j1buyChgGpSbBQZlDTKNl
7dvXRnQFxKEI82j1cLU8SyrnZdXqQxQ54PZr6JudvAkOSgizykh8tnRnxlPs5YTs
TJlpaXltM46xFI2W2+lnUkczlZnSDt8DjiiR+rsONNhMpgCdCxLNnV9e9TFyTLLv
w0Wghd2Pjw8pAC6DT3n8E/qcVDkaKBZK/QuQ1vrJG16SJDUBg1jKBgYAisMzMn15
4f7t352vo+Ksq9Ifcd4CmKMBdMQlVcRJ5qMOiAODp2CPHizo1UYWpGjtXyq31wg/
FxDFWCyP+hctB5QN/vSDo3uDmGpsraJEc05DdZCeh2VYkN/omATMrFpIvVjeYSxi
+6+4KBomfwgVo/I6Ahz4i39Stgz0tH96DyfD2zgLPRVpX/tl9FEcKOiJXBbhvMGh
LLuw8tfWkEGjsT7g8tXv4tQApbsGt2/mUhoBn8Sf12czAXr2Hc4Y6K4nsG6oLoLM
sOkTPNcE0XcppLAYBi2ET9fyl7ZrOmHjzUPvFvb4xfBNRf2lFj3J7aJ9JdwCbmgO
lTrLAR34xnCgbLOy1LEppupAFtJUx5HjtG+Eo/Vzm54+Tb+dYiZ3ooKf5wRjs7GP
RWnCDHDOM2kd+07zjxcPHLRbGc5Nx/Sm61EhePkEdkzHTbEvvVtP0otuywtdqotc
0GsnAYIlnVIEPKOio+5omahtRXyKtu5X2THBZxKBKo8TQtWfdMZGcNVcZpWDW1n7
siwW9U8ww42di5kUN+A82U1NfA1+e/D0GgfH7eYJc6TCOqFwY4OZDTzQUO7MOsb3
raEm3wInwGk9JPfWdi1nRf6+rez6taDThLUWf5oMbkm5gzPWBnxJ5w5wYhaVy/K/
liK6w90CaYr/Rk02O8JthsNc0oWpTqw4VRV94xjMl3yQCmYjnStpbCqJKFscH21s
iMM1sH35Dtp60QZbEnYWIWuMzkYQfHeef4i4MVAuDlMUdPIL5+yROBHp0TggOcU8
z9MeJN7AMp2DFQDCIq9RWd13HiMhZC6HXQeS8pmjPKWvkYwhVuaMDKUP825GoB1k
CnGwOOF9XHijUGqFZVnVVThK+U0JEyjG3JgteTth753sa9Z1fg7Pn6AukdfYeZ77
nxORIPxvzMTcNIboPUQaYjSK/v8ZLXPwbSqyIZu5fYUdcdSC/00t86duE6j3APzC
etIDwP6d/Yv7J771xm82htzwvwrS20kCTgfAhHzCUiSUtGLcdE/Bd8Bh7yo3TIr6
61rIl491k5FPRXS24r9FobBe2VV3latpCmLq2gVYdQQIgtbOh0zR2HqO5+wX4R9L
gV7M+66nB5PchdyggoZiKNrhfkpDIoP2G6rIPyBxehL9zLOXAIkNBbo88yhjt3E+
eolPdXCYDOy1rMavUsAmT3ec2h9nKSl5sdx/P+mmpAOu7zC9wTaYFZqneZ1tkMJ6
86D/Q1aafCzFy4QSWame3Vwj3wyiWynzWF0lf+u2yfzqq3PgEKq+jqhx6B87x0Ui
yAtKlIcFFCtVXsO++sbEy0GuCwNreLWl54evVuOAV2yEVRRXD5Ka9US7DhTcRdL5
sItckZUY1Ql6SafG8SpsHfjEQwcrCPkB76v3wakJHB0J7Ru75Dai6vx9Z2VfXKqy
4s474jl9RRJunQdYyF4Mrb2+CNkCf1Ey/6i/yf48ZiJSNChLWqJClD90j44QWHCk
IKndV1FVGT/MdBqdV7Td4qs1M40Kn2PX16AZF36RCp2GaMvsiniEyQGQOTjOkmyI
iClmAYSQm/SHwhzyTdpxyIgpfwWEgnS+GKmxwZRPI2KC94tpA9cLYtUyx8S88UET
EEsiAP/uEnsfs0jevwuA8E1vfFyq9Lzizbg5p/kznyymK12kcek6ycXrlFEy8S9m
bT2iVY9zBbw7q5HD6zHWBiqBkjX02wyzsMbpImxf8x++Lzx8DD5gVC55KqDuyfwt
SjAJxJY6c267epQjQDzqjoCG5npTnaXNNDJtWDZ9rLrw/SDB0B+XCAoFua3mGSdS
I6kpiWknJwNOsn1kj+WXvPm1UEPfgN22P3vzhCr0XWundpTeEU0sOPSYw89GIWTR
9sOavfyilqYE/5d0Iz7ftyMCNquu9hwOAlYQEJ+ufMWhwH2mYbddEHbAgknYCqPw
6qSD50xufsnG0lIPIQ5nW2ILRyYvT3Slt+MNnPy0SUmNTMgP/vOvdZcBqLwwWIDl
oeYTNMvmNyHOZEnwk7OMjsnLvqTQuM8dcBEt63PKobJaX56Yq2fSPVnQgoTwmV4J
fLTN2cIUIXzLQ6PTLF/dam5clvZ/QxMCqXomCOj13cynxfDe9JgYPZGIbF0VLl4y
8hKku9DdcQoSXWvW2YcopJiDVk7PHoj7C9GpOCCVviLR4n4H8/lAQZ0xLMgl7J5j
GdeH8o6Fl4fbCqTrGyKRwdSyEaRNrURiFu9leIMsbPqziei0GG8nUhT75K9CQqoV
gPZ5DOuHd629exBhbve1PxKudUOG3zc+RR7C7p9EWzfXpastwwppfQO88wrPzioS
peJ+XjTHP8+L3d5xX6d0Z1mWDEuQjZqL37NTFkejy1geAF3UbRq9D7q/e4WxComR
JmGMSt6ifoAEjTPX5z7hjHccVRTmYmWd+/3gpnWme1n30j3E+VqXz+7fX8xeV1/M
IS0Yhfw9JG9tqOrKY0KComTbm5pG2+u6V2Rf2WZgU3xbhdIp8mCuFJMFr9549fd7
95Vgum9KRLiXR5C8BuMkf/fiQ2QsRRxrQ6sj9UvuyINHFmboivWIUwwdHbrQr659
lfgxHoX/EtDV+q6paVLUbbDX2x04ljbHK+XQ+MNUbaTaS+TB5KL2n6nYi8+fOjW6
dWRGJbS8eIcp0+2enFyaRwWnw7lfluFtIYOAGm/tEqkZMRO9Y2u4Re+CTE0TcltQ
jURpyULr7QD9nViE6/10WxjwYFwZS7K7WRYuZduvJBTJ0+Z7vKMjAAB/3qfsTMx6
UTpXw5QFORJ9UswOfNhMSnURGzAl9I9Btb+gwtUEYnYKVt6c6rDZRpfTXebeK35y
5XlFXzMws9M5xsr8XpOcPMwb9UwKWgMFwoV+OaosH2lDxIbvgFvawLgsCP22mcDO
Z6Tce52SXA1KGFRxfQt93gBtm7l8dNv0D6rt8YN8y9VJA0XEiyiNXcnmydKt/QRE
dqI5cFYuE6L7wT/mStUdyCgJn44A9FWNGMNFMJLUvjwFPhO620wsIPYOfsOnk+uG
FR3ustsnGGrACFxsH5UbeBaeIonS/Iayas0UtZR8zTmPUKqac5Z2kL1YKdsk4Am9
V0PaH/NqLNGE/ussxDS8aCj7DAJ7eG58WypuENHJF6PfStnI9OmGIDsBI1VVhq2y
8/jjrR/kM9WmRNJG5sg06qeHiBqraaFRBkSA2+GAIRcH0bCRxq3aa+bajKSUEf1d
GQNiYGJWwlCIzLIlluYzildeFWBC+lN6hXMx1lUs5HfG6OSnsGjcq4UxNWaBpvdE
OoCvjKvxQPCEaJ9T4jSrcdhU0yuhzyFmQh7YrzKRdRzTAYZ12OHDNMIGwXDDsXmP
a/Vsr7Zqm2Y1mTyx050MhNEvtKKPc4G4RbJLY8dAYXRAAPmX0znLZAHQP9cdQ3sT
g6jUBJf3sr+K6eAC34fnSG1bwPaBtxt5jthw0AavccA+1yHc8OywM9mZRBsB5KJ+
3m8UDHaIpxFOgdxUULGVWYWt7G7WLjvtjrliYaQnHrICXDq7sznsCMWBpiI+Q4fz
jkHjV/Ur/O5p/sCVs+rxqCHJSNMxXPnWugaDFp+aJjr7iiG1hoEcEil/38swsgGc
TuTPYm8MNJZ/0ccnKGbihzuNpxbtL+YwCwA5Qf79ayw/VP4t3CHIqK5cdMuM0mSz
UQTIB5FYfRKMOQxY4HIKJAJGF8pBn3ZP8+aBPQeD+ZMQe7m09k/tWMPE0t31RWl1
9B0AsKQU/u4ozWkqiVGCZR6zRS6rpjQ3Y6OKsqZLoYCOEgKaRIXhL2vyoNaDKfqN
U1nSaXL/jy+5Kxhh1/5mb/k5YKuLgqQ9xyekzjsQjEtqot6onAufUw9eRe4fGVuZ
Uo1oy681aP1kDaQaKI+Q4l7clFliOuC3DoLBXw76PuKMp5qOlGrjOfdO/MyhcWBS
KHepXZ5wx3chc5IYRVO2WhQSz+S5h4P509sZfot2lY4d0VhCVVQK7s+3DaJjzbaf
Ny+mqpcv4YP8iNEvFnZfFG9u+UUQgoyu5cAIDk9BEoRpG3x2W0rVuT5VnAeTU9ha
zwZZez5NOoWpxDHVnqqrQcqFR6p8Sfnq8G4kT4NCS2fFMBoIiEH3G5yJHBF+Fyd+
lc5lcPqkLPt1xhj90DMYWuUf8Ys6Uk7tUG5PyYM0e3FM4XP2hrPNrAjSY9nAwrv0
tir4uGc1uCp6FS5ycePVFrcQEr+6JVtz4gtuBskBNu7o84eA1ri2Be3vemUKeclF
x7mB4OnESNUdMj5exXMJ8RQkbdAvsHf4Rg+YjxnZ28owHNEFx/1zNpYGjkTM72jl
OpTKwC6838AEhS6JJc9giVn6G8siMIQ/KNXdSakUrVhdq5JTtnV+IE/3/rEVJdpt
tiReWzBMEnTnjO27XulHSDIauJOQlfzzZ3lh1Xf2qGXkbVbk9iOSpU84QtYUth/O
oNPuUiJhLOj81YIucqF4D6bm5kEjCaq71iHo881fg2BiLsgCvgKUNQZmntu5xNaf
EXGfSklHBLDVC9ZvWweDJeCxW7YdKToXNHO59XTzQcCnrNe6VxvaPh4GFCoYvljW
gGzxISrtvZK7qijmvEpfmjOzsEawdlRyfx9dx9qELP3r2JQ12ahvLZ53/BB0vY7D
ARXYe/FITNaPFeqXdNZDGLA3zTUoEbEg26992G2a8IhBIc9aaPdISoSKGyH7/AX2
KyJUIWksa/w6xomhZDe6D7f6ueMW5JEMmmFZf7hTiRwJrK18cL59eAMlqFgGsyyk
wxstctTZ5J59u1JAz3zbZlU4s96KY91n/BsAeHik28+UbJGWgLP721J6H6I/VuO0
PSmXXdjr0lbjyLTMcWxKGRdR8EUUrEDsyM+TAigOWIzJP4UmyXNtEGBQxMK5yJ+4
xJGyHJ/X6lcsnX/dzBtDByzu8xtw7H63bxdSmC6Ucbzb1YkyDSU10ii1nA4ESXnt
Vt4pVtiX5SgAwAPjzzc1J6Yzh7ilMr4z8z2cloAkqstNjUyvEgTx64XFo0ydJ4BY
RHstg47l2O7TizEclogCFlK9NcPaeEEq5TreX85bHQH6WaydY77nXr5reN+M0bfG
Mj94AgU37XhRPGn2uAQ50F9iqw3+7hqyLyb1Ph51elDt+4zvzmS4lBkDP2yjurJc
NzSH5GgZA7ZsApc36C9Mf40QrzHQ+zGt34qU4FYtXFChwkOWl+lKlgWX1sosOv4l
vvUWTxPX3J2HaxwBRJwCvXBavv2MPAVFFei/9VzLBl5hqsaJCqHYPJ25H0yJnNsI
4WJ7HpXQZYciJblyZ8r1X7HOh/xjOQWghIYuBS0bKyO9+S2hiKP7PwgOxN789SeH
kel+LalrL7i9PyHFWe5lVUcfgKFHA44zNxNtSmRIQ1Dx050QKWQLcLWeMSTdwjX1
oJBp6KhQklft/5PCzV8YxgZ2IThxb2K3hXhozHeh9LrCtioWGWDR1Y92X3NnUE7I
Omouwb66+7S+W9HAudoq05ZMKDeZ9GcF7/XM3X2oMAUw+aQgs9K+hXkwgpGWG3AE
5xfCiOFJA+NH6jDprHhBFcJY1avF0ygSd0STeWUSBHw7xIj20cPC2GTuwFvVAhfw
YpR4fzQqPS8wc6o3oXbNUnC5GyO7CLC+UJhnDh8PEsWZyPo2yynd+Zm3SzZIE/C6
e13/zgu8DwibaNm7UKP5263t3aGO18Lsr3QRfxDRQGpF3tFuuvcU4TC/9oHmxMzT
bQkKkj6wIxh9RJRHl8n8tDUDQwkjCtB3mlZSgNECUnvljW5sh1+/j03iFqqGpRB9
6FGdPb/tHdm9LGlQVKukG8aKcFXrPOWCoYFEjSLcpiL2fQdFg9BTuot63gGSklNj
KiwX2FlblabcADgT4KVoks9ThQK/tmepvRJ1uILZGUk6MVHp3BLQQ0VJcidHqTB8
4B2dZuh3YJMuAHlY85+W9F/dlCu3bDfm+P5C/WdpViAtN/TLGnqaj9uV0BqFow9X
7Liprt7hQW91rAq+mbZMA2UFwlhrN4qmHfR5SGyz/1oBaLf4TjjkzKTMXUq3hved
v5f1DIJ6nRW5bxugZ7RS6YFTek9FH7REp38Be+d0Q/h3efRCVv6SQJ9iyb1c027n
dc1PGLYABRXPHN2+EFg2MQQfuZZNh82f6Ch39IC2TO8oGHXDbgDnERbw7oaEaj9F
322au5LXU2g2r9tbqILA6v5F1cbRtR03jF6Oa8j33SJWbK9vhc5gNOUKFIWA/jj8
4TCyVBqyDrnlWq5/7lABjVvltMfsg1xcigmgslnyHa7Jl1Xm4CAflmmxSCfCeVC1
9zIpnR/ctzfqKpPb0slCJLik/++s15pUitFReelNs9N4w5GVB/JM8obFw8eLg3hh
1NKlSWguzEDFlHCL6dFYRfK5z7Uf9wzH/oW0eDi20awB2/YqC/YbximRz/PMEsB2
mmSJjwpl1F6JdDwgtPT/zqBGrI6v1j2Hc5MGQIGXawXBnH9AOa+IVVQfg54giw93
/iIamz3LyrEar/eQ3Z8qB5ggtt53O4JsW6cDhwVH0OxRDEBtrLP2/NPdz59oiGAT
xc0oXyOBy+Kn2i5yFdeUKliB8rOlWiDzbFIMHp62i768Kn6ECV0bEDbGHd9djBgd
+36mXXB7WKXmLFy0KxXxt3U5FA4cKJbyBzBKEbQuVQa8UXzTYto2LXisof5CKV+3
MPCF2OdT1jBoxiAy9jYAJ8ZX/Y4FMnyTOZIj+KUf4ho/QMiMADQEMmNLthhoZmd3
GyXBtcj/FgVEjTHEzPh+NZHkL8Y+ym6zITAhQr/T8jYIhCS0SwwXwQqlTnwlyeXs
+Vh34DvlHM6lDoha6FDfcxmefG1s44w99HeWS2QZbM05LDJhEOLmEWOuw0X2gqwU
SYYLYLlAbfgsN6yNmpr6rHJXmZ1BXKA3NhWLFDWSao6Mz5O3U1Y9NdWtoZJvi7tg
fjYsIX2emQR4vupfc4CRP5kj5vfx9cgfe9uxlfWo4kaQ7N6CkteNiIJ8hjyMQD/e
J7MU5rqgcn3U54YVUmp5HCSbmmur1lOb5M1gEpz2jQxcUzf3tifLGcJCyFQUW3PT
px4zfExNmciKsoHdFuz9R19dFAiKSmR07/oCMZcsj7/IPTVqtWOHluDS/ebjRIfs
FNjC9OALAdl3lZkcRAtn7hTRJz/31VFy5sZAYNjitSd2JUmfJxzczuk3mRbyisjE
1Ks1RSprg1Bnx83Kf4HXk8sfcf3FxEwKi/o3jI1HVGv5GdomhDMHPBoOVs1zLyli
W1HKY118CtiZei5IbmDenHY5XhJRvRS+GN0LGSFLcTeI/GWgQ0a/6+TPGWDlO+TD
pYY1dfwZYIbl6IoBeBBB8vpyh5TehQunPZtlQ//vW/CAJRHVbqpCZusXBT+qTlq6
U2agc3AmWnNObLWeFY4l/fbHgnTCSxM8w4VoUJ19s1bHj8af3x7mv13U23+K8kao
6K7x+i949I1C1idCB1Y+RKMyD64FLUAPABI7LvecwHxNLdWCx5V8TqTq9kJWzvE6
3jiWQVW/hP+Q6/Vk+z7tKYXcm2QZj1qgplfRMQtYtnyLA/AyTGiIMiSWjkHXTU78
Gr7TIt6sZHbs2lcgC0c2p8HSzVvG+a1jvh1a9DSUYVyU5YxVl26VcesQ9uavi9HC
dgCMro42jFvgdnUwD68vNo5ajlMgVRYRo5qmiGyVL1EBqCfQqzA90PGC5geAdfR5
3sfXXf2IjyIlRiDV3zrmJb8i5WMpV72nQbZ7fqy1AvXnuT1OeCm4xhei3SXI1OXs
ny+ZZyVRD8RLNLdtRIT9JoI6hBH74WRzMi6yxZZjN1CgHeZ+Er9Q15BLkbm7YqQx
Krbx/3ud9c6uvXvWu3ooOWNYhzhQbCKNq76GYhrUmnqIfGGTJw840feGJF4l3cY4
FCzrJ1MUJS5r6cSfquBS2/JnQqO7R9KVuv+ZAGUY5av483z5Pndz835tGZRGNpuL
4OtWddIoRdrOShjg+tjwuxFHkA4CuGbrkv0BinexrGY4OE7HkEdSh2jjsIhngGJr
VzXYf3zEyGsbapZuFhBBtCGsP07UCLG5vCjc/xJ4IZHOYxHUjeuXrDsXKE02s2AG
ipk20TZVrNZXevWCWJSRALcAb+yn3mHJikIsIkOIbeK/5k/U0u90v5ghuQKEPtqK
LuzDOgtjmNjPi84xo3t+0yNsZLFzpPqhOBa7IN2iB4fM5Bi7V/aQof1bYlKiJQ4Q
QqZbkyD2M6xC0HjAlR6IttXGWNJs0+eQKF45aSH+GT/RKNB8sLtkjT1On00Wsxry
rp+iqSN7qpM4XPe8JyMNbg2t8qdmhGHcqNxI1+dMx1v/hPQymowOwK+BIe8dMiJY
OCvzJjGQeQhzliexhVsOlJQD1nFOAKWbZ19R55Dk39QhxhcAUGe0r82vszFaODkn
6Z7S7/b7H2oKByV6ocZgHHYlt+Z/0x9hvhdEb82bOjDPLPED+vE/gdcbeceWkSJX
jwxpoei8ss8PlzbDr7wmbI+LiNyPAJxty95Y0Zop/Tu26+D6Kf3wY+dQLrUgKQH6
EyPSa//JdnJGeqBpsWHc2gHYpbNXBiQhxy1lX4lSvdkCkGRNwqHiF7iQz1IOs5iH
Ie4esOzMsEdXJnrM9w+ldHCRNoOCUMaUfzawi71zR2CHMDtwPcswBC9WzlMVK7DT
30bYlyaqGQ4Aw9xUFPNN+HgfSOBETtKu1jRxAHqK19OoILrX81kqvLmuBZJ8B0lV
dW+cpRVnrOfVnXUJe/Wn+44JcTHCAkeTxtWbPcLLsu2jR5C4I9LnCVT8ufllMOhx
uZlwdGQ4UvdDNm5AtxPNSdDXnVSgcCAGhhLhFJAtJygxarKq55oggL+XuZGsQ2OX
o2WszbtyLdBDldIdS6YOJoVnzDRzj6fkJHyITERz91c/41WVT0s692tRiTfTxvmi
yUzE/VkmtdZKhbOaQ2mYcxpazO7Zvvt/C11wUTml1ogqBQLllA7mZ4GuHSN5Xpm/
JanZrg+d6v6tYuh3gbOpgJplhi1xkIOyd0H1qXz2dMTPKSpqfSvx1hLz/+oxnqOx
DoeQ5uvkkeFA2WKj2q4LO06abzy+t+ZMktEURXSdRrTQnFG1d4rdTwXqQML1pucE
ZRWQQKFrzHETa6RW0NCnrjxGk7UDCRKczsIa06hII+Y3AZ6OnERgJFbwQm+XNM6a
YDf4RsuzCrOLnjEOABJ1bishy4pLGhqQth0AXHM+LvuFNKxuGwFkK0+wPi3KcIZb
i6dS5XaeRHLQqE/4G1WLZmXeGmj64u4jtsW2FjauHZkOZT8YgattlHE8qrR53sXO
Lnu4K6qg8k9THTrgrGCnB4PXJpFH74OqKfls8rrbKcKjlqFeFgM0bl1klHLfnyOT
VGD3+OfGTCMTZNNl1iHjiwjMe9cCDWmF2oyPxa5SBAs0CVec7IqlMMAHkUSCc5qF
AXKYTFAX7cf+hMB8eb7+5KNGyFuFjmXmaK2KkYt7fJFIcEzLbZu9e9/+1IywDDvq
go5xOTf2t6K4WbStt7JMo3DXVBADtucwQNPxauPow7nw9+j4ssG8ub0YK7x2i9Q5
Qq8n8bRVwwj0mpMe5FS7atZm0Ko/tj+7aC4oIfP+/V1OhSk2N6OckgpjjB+D6qjf
jGutq/hp56lcfz92lPQNUZqeOG1FtALq5cWjHgaX+tTDqtYyWSX9QzeBGGlb0AzR
H4K8uG3djCJwMkq/aSxiPQZYLCsSZbS7VOsX+EIKlOEDUPFInRt9vArmbR2zMGFz
nyXeKMKLjNSqn6Avb9Nn5olClMvVZ96x4WvH0u0FCwxN/O3lL6TXjaTutbI3itDw
Z09Fi6HkwmYSvXg9HASqvWXTYrt7wp9uAfBqVR1GcZBrPy9DgcltmrcGOIEwJK6w
wtVViLvUDv3CWfbEVxGxXofcxJyDkx2w8plWXvOUoqxii5Tr2oXZ7I5RQgHlEHmc
7BXPpdNgpyryHlMqKb1GwIVhIwI2hluqmoiEvZnPEhYxz4Fz/TOGc8ePH3zhuRQC
Q27XiLDz4NGZc445WvfxMtAeoLKYOh+LS01mfoFyhWC5bSTjMtWNFNxOMMLM9HsV
w+duDRbLNJzUKZyMbPpRMVQQ6gDcVlnPAYbIGxPPPXLEnBprylXPvTVHuGyEXK0a
ANn8g3FfP3508VnW2Gqgc25ti21L2NBWspPDmJd8ZKirTvTLREvZ3wK0T9iGOrYk
PBgPaGwbQ24TKs15pxJNkp/W4kB5D51uI9Vn6pRSjXLo51f5+ndrsVy8LwOOVrdg
wus1I+5yxYK7wW0vXxe4Xz8aKQoBPVtVMPDcSwcLVt7PJ+QIBv+SH5cnPk4bDCba
FEFVLqIzpfMb753xrVfLRMw1li4hMXPJqjGMc+QJmTdNNLhWTu/1XFG3HhlhwWHp
ZPjAnlbKfJkYxU45+kajbJowpaGO93v4LRpUggyExtVEnattjqVeptLr2uCmj/Rp
yZyoq+ZNYA+GxbCiBZc9/YiXY+WjUnHC3x0wAtNkA5CQcaP5JuYcVfLE1ee+PM8A
5+91hrgEMXL7M3BrS/BfpTxWQYIDYqFpswzqupRoVL4XdkhcAktblfHxmI/MTlrx
mrouvdpQRFQ4F6gTMo7wUSrRri7RamF3D92vyaHoaBMx4in4fMIJ2gN8+oiS0QPO
UZEqBmAlN0j0RjPWc9kRfyPtoMpNFOtK5kKTKKGvTZdzCwmpLAyx4ToYb5cna7aS
wXtJqD/igQRP5ZAmLo787WtaR5LqQZcdaD4KnJLqc1zH06bfuzWDiRdF8ZnybUUF
4yqFrTOFwhE2EZTntxYNJd6hfEnIqqk8n1dwnZeN3pprCx0GRVINd9QvG0pZRx4o
KAPNe3Lro76eNp9MNFCvV2WT6M32ZAJKxq44bWwQWKecwm736Egei1MnALrkBvMz
gPYgAEYNs8xZZPJCGE8Boi8ZrSPAHcvAXq72ANKC2eF+X9/DOkQlVYdmGhEp872O
kRAgDGO+PBiIHYV8odcinMztR0HRYbh+COlVNqhf6Ug5xeOFZ57sx6jy6vM+591s
Q0eB/hZNXbhwEZ48mXFiaq4bschR1BZmhvmbX2STnRGLGYpE2t7kaOnsiwlY1GTd
YCa5He0gPmoXb8rPNoJYVi5hNTwjX3Ops2XZFaCjBg2ems1YUmyUZsbUp/KwZxEG
Ewj++eQkxQD4/uElPg22E2Cty8fkPFdMTIqxA1uwbSoXBTogGtxD6xoR8ZBK14wk
sc41ShskHQYrI6sP2CAGl95xbXZMSvoueYg13mFH5cO4SGX/3zHoVgvSI84q7LzY
fj0rMtYe12FMuSlJugwMJITDQ+WR3SonwxqjmbBSSwEAv26uUWVWYOd0QznQQWDL
iwMLSaWwpywdFH5eDimYWSTkWy3dJcynQomOsBldkiLH77ryInrS0IvI/Wkl8LLx
XqZPUYzXpXHCHoqf9i4G+uFOfShiUjasnJNFKx4xennWhIOiejZD7t4v4wd18pmj
/q36PvvvElt2fXrAjotZ7RHgWEXBi2IqdmlDgXkQXxlRqgK8vamGLx+b2UL3JIb9
XWurvvldGWcSCtTMfnpA1JqD7Hg0D3fzT2oHGJuQXlQoCa/TXrqY+xtqJZRqg0NG
cb6xB6vM7BmMSVfkFNiAjSWGlzkgqz/JKrgfpejV9bfVyNr5Zyi18ansrCnTCaHF
MWmlZz+VxbxWRnD5LhusqH//j3GJYYvLCU8YzQ4v0CVnKM39jvXIxaU6+kmBxxOe
dqWwUH7fH1NakdQdWl3EIrvcsf/KZW0JNP6J5RbFZbEe6PajU59Lp9IOuOtDlEmr
wDYr86fPCbEKXAp3lo5zzeIeSSzx5hn4t7bcNWNkARfSzmrOJtzXfi9gnvs1Jxl8
cP92KrnrR3MCR06KNxIPn0Xx75aVQexOUn0joA0bzTt1Ym5VlrW7f2QDjoACOF14
nKIHSnG4ar3jAExrSJYkvAPWhSDHb+6Squ4uebBxwew/OkKGA6mFttn1NgoSQ0Gf
PVKquDl84WwpIMZHMkjRo0TIYjo7zgaelPxbENuoSxoDiGMfjTUTRQRIUkgCAw+b
i1MvLQl+Pfu0GsMqMltI27Qo9HLfkgbkFf4q17dSfubt3qqfTHIRp1j3MLpFuvZD
DWd/iD4ehDU9CGjSk7LeSPigenhWDvDz77cZoLEKXQZuimuT4HM+UFa8qltq89cT
rrx4Br1Kbi07grNGjZP3GGUJtYqJ9aYRCjGfuNMKKriPM/ZjQFiWC44VGVH/nOiu
fTGcPTZRWxwFb/6/bRhLgMVFO5/BhjiWQoptmkWHjsM3jz5LNSiyPXJQm7mO3fQs
BLd2rgBQn43pFPoNXkz0iXDfuWcpr08kraV6fxhhfOspDbKEINh5qn20Im4LkCty
/Ur/JcBXk1O3sFFsRhJ0FGw0IQL8ezRchJhSkmEZEP7knW8Fn/MbrcBxTWNqCSU9
CoY2+JoYnYZGInxgLQD7Ixdmnj2p1DQqkYTLKUkJjOYT72Mhq9Dz5jqEPkzdYRFA
MjKu86BStJj3v6w80in452WnNwFRCaPXOQoUGQyIO/w6q1J55FVx8t7s0Jud+ezF
es/yBSNXpZzaapSvdYVy6yMf9aextEw6Vk1VM3UMh1MDDxMvaCCtBGzvje+TZ1Xk
5IpojziCiXUnGGXjXwBf4HP2HXXP+3aP92lkWE6IY/d7jVV2KudESUQHN2Xk9kMG
HbdlVbuLbKlAaUex+doNmfUVVWGcG1iCLCD1kEwR4GFdZ7BdsN8iEQEZeamM3YD/
Y277ZwpNVH3bjQFVj3wPzChbufP98j/3j9QRKVLqcoAobXGU4DpzjV/qOg9Ob8bm
oiA0tDk24Uk2k95TkxlLLLd2+GZIUad0lQp/sGN70poyZffdaaN19p7JtWdx0Xxh
dDNEKAbRwehx7zu/WvvIPdAgNBBuXqcg4aCErH2Yc/w/u987i3/ZOSlFGVSOEZ0s
5vE7lnPaTg68YX3bdKfD9XsopbAA1SZuYXe2fpOYIQyHRDEF5rnoOJMU8t1hKK62
We+/kdAdRVVe3hnYFQjmv8hQCbGV675jBRg5FggupE7RWPCWf0EC9k4YIwh1YM1R
ME2vj+yTGUTo3oIOKM6dhWZl0RYTq1GL6s2dUfvVpjmRiE3SKPC7OH7CSP+QsGJ1
LwI7woOckTDwR5LnnrVgaYLtcNOS8DWMzZPKmlsaOw+DC/MRw6SjDyCjUsuTOEBc
SoQDzr6x3qRAsr0LZFjDL0D5wnJ34updOTSSYm0X/IQB9xdvFCgjzhfmesziPJ7y
hnWcZ32ew7xNvMCDSus4o5vV67oVpkzcyc8qKpnafKWMu5QnYM0HeZutYqkJpwYD
bdhCD5zGeC7a8SWg2tIJEXuMMimwOBRtZQGlRSeydvTAMGZujJwnGzPafJDDDLk4
kM3FWLuY07rP2PSSlCENUzssFGeLm0KVwXcyalqJu3uIi+HQFDFBBx7GfGrhs+N3
mFCIhXYXzPX+xBdaJZ4WzO+SV+SfJ5a6zo5wxgRHtoUvuAR92rvbhxgIxplTPs0N
XaILh/WdP5supyVwHA6xeUCHn0s+NAI16VJmQZ94k1kCVtzE7jy+8G6e+7fti2w3
XfiHbvKKHR4p5CIlsyAMfsKuLV2w5pPxemo17vjAHZ21P/2s6xNqmBfqCzHo/Y+j
gOsmVcaCr+GPpTOBQP8r2K5h6Xkxr/JHNQDc9viA+Hw97gm8WDRfsQDiYDhmluIB
5cHwUXRPvJ6EAI9P9/KR1F7XzoUQT5lC3WGMYmvX/KA9D4rIflWzoMS7wUP3Sbva
MGqD5SDKMJFkN7QHATOKj26oAT/tbBhSQBpjQedYAUm3sglYG3GSq3t30TbYtufA
Y0VPqZUZgNzyco6GZou2ZcZ2xLYTbMU+sPqlgEantqluLSCuY92Ph8PpJ8kbXrmv
8hJK8FtcSBNjJpHI0lTsQJX1yslcAy+Mw9xezV0dwc08Bz95vFI3axfpLKegnxu9
ftI7PGdL49X2IZTDSqUF6WWw2yYc36onuyUtxPgLHOaaIl5DWCst9CUkugVyFgd+
ngA52Z1tkvYvzQ09QqSgjRe7p0fRVNABIflJmkTQWSl0ncNgvW3+Ea+ZobmH3F+n
/HbLPeI531miLukDXQqUokqP/UbhfgLz/sAhWjFLC4epgRk9GWfTT4e6pW7/UPCb
88ORmarJi1DgpOXyoZtgltSgD7/knGSVAbjLxD32YI3SOKCpaX04MNpvT5n8jzLK
0e9h8iuOKBcM2bCoC9IdA30b1LRgFOkR6+sGyUYLaDtlscQrSvIYazjGdec76IKY
DNT9tUwwbya1HQANhizqtpuloG78H96v5vh2/DJMgxgawqeYTWFt0MGqiSs/RSdD
SbNXT2S6r8zkLtrSuGqM1+0DP1DwSyEXoAak89y92v9c8TmaEJqars03xlGB4CwD
g2jKs5I52z/hn27HaoxqBOvrm6IJmJi/MIh260aQkmRM7HPDzIqxcX8HaJEREczx
yxjJTCsLcOGArxfZScypaK4JeKowbvUSMqCATujzptRbY/fz8QZ4teSnQXM1B6h9
UGuu9GJcfYMmcBujTHcCaopCQV00SOO1rqg3G2Lvdr/ObWJ9nis9v1YYIiD4Ji+W
6T/aINOqlSeN1JBDQ9M6COq4OKV5TgyQn9pCt0FQC1npMEV2Pq6OMn47nIAWNryE
EFfXO1oOdLM53qXDpaG7Aqe9No/WR1QdxyoFdzwdJ1h2HpZEmvz0Qz08y4XoBT1t
PxAqlXQLBtIQFB1p+RGx6UObto33C/v3hgGQXPAXWJN6P97RI0UIpEJI9gvBUlQW
9UyBh/FcuibtsUHqpid7ZA9pRnO2+xqonMvRWexeqO+m4lluLLeYovO9oiTxR+SS
eXJ8ZPDKulDFfdSwPT0i9f3kQ8u9jM6CH/kgEK3GaPvB0IWBpz0cQ2UjmIDpHl8C
9Y7ovssXUcXH2jf1h7jt50wjsTB9uhr1i4XBwdxfw3nLeak1oHZmHMX/z/BqJpYv
BQmk7AsPu3O/XKsAZlC1B0HM6W6/mv0N5k1FeX8DHx/9slwVYV9p1CdU0I0IlCCn
TGr5SLj5yaWJGtHkI2pGkZkvAYA4J4IRmcywuSOqe9r/IHyzaYL24HOnT3sR88xN
lBd+c6T6mgDrBPsW03c4CBcVGUwuzJf53PKX0LyYdY1If1+t+kTDw5KALjgmVH6x
UQLCQDbi9nrndCfYmoGJWxe9JDUCiHi5CcmjVTHLQZRR4PzpVYUyX+yrU0vFH04o
kUnbh9mPvtzkTHQW4edAZrRJCVqZH4ieIETI0dJb5sIJDybqdtwvV0xVRMloRrl+
e7+fkMEalgXspdxjLnxve3y7WP5yrR9uB3jLIeYPRUaKal6RFQtku1RHeIRgKvhN
5gwnbFlmOX3qs2Sb8cnrFQ1DUkUFFcL4EsgtHrm/4mPEOS5XrqpgiCwCb99H4Lua
A9uahaYsxi7oZZ7rXWRTTScd7q8VRV1q8OkU7uXwPUPMH8iJWyfbYGRingwmEE+5
jh9tn+Lvg7mWNfV7v3JEdMeKMhhPKz71WRulxCeoIHaQYIMxEZfwP2Bj9ljenwNB
zJo+iwp6quH4SAAKgNC/AstQts4t1Wiuftlz1qY3vrlPEE8UI/byL++voDYV/pm9
DwAVWRUBc3K2JG+w4sKKYriSiWhgP7qJys5P9HSrSjJ+ZZu23YIldIMjy7bzROYT
rb2P9hPAtI6W8tN4xSznj23EaQmgUW4oulgdh6FnmTs1GDpX/QoHmSTL19uSXAJ5
imilkJtQAFDBiHqB2qmQiGvrS7wvGkahVD8SSxSOjEZsEjkUJIdutgDM74MI+tqL
xArcmUX64GZiJm8y7JZ8qiPYCYOdMWh9qdGG/kenWbdgDyrxj/5o4R8cGN0RFSAf
q9lassGQw/yHKye7kG3gp+PV9rFv8NHGpt6VvjsEBU+E1ReQ0BtFr3Mfi34A/eO3
Ol+MfRLkWgQvKy3Us7tvEUzrb41knvjyyEvPjzW/zbmv12AFxe4N6BNu1y1c2UBL
kT61NENNyBMkkUVDN+2iPBoWKiExlYPqCLV/3WAbE+LPxNTvX8ezaK8cGimxjmn1
ejEqtZVOq4botOEl+f2nffkfeYi/iDTtFypNEgng+cHNKcOHttmztqzqzLRpWebC
LQHPl08sqee7pgRppSZyGtd/AHcop+S7HmfZTCqX+y6znoPep1M6XYsF68rx6kkm
gnfgAcjdQ3bVu3LOLBa/Lt2C1oZd7EWhP0/yp5hH6mzJmPhAdQyk9HcYqDGdnSdI
88AHv4O0VufTRjLx8M7ucxl5D/WAKdq/EBQdtM4M2q4jBJffIvbhHLxOo6v2f8lh
IWHdQ/pACxW3T12dm98CVefc5+J0jZJb9NOAvJp1qmlopxgoseW8IM2fwNsqA2wu
Pd2nr/olfF22/Nodzvzrk6H3fJ8VC4wgY+rbo+amlIvY+FbGqVGi3qxOXrrW46C6
fJLWUJ5BnMpJQkIT2jLY8IYTlKn20F5rFuLUresNu0/aFK+fZ7cNltOJy7/RK2E+
OmsueaZmp38vvG48b7MwUj0nmy3doYxMsWyAkVRFwz1fjI9r4QiKAJvMxc13Wtjy
rtSde8W/gTvobTyAH5+LweBcDwW1+oV3+d4uZp3KlnHbG68ST/CFGgjEimz3252E
T+E8LD5jscAlp1Sa/cUtIYzyxTlbLDJybCQ4yLHryfQkxnKykN57T5ZZ/pdUQnMb
hUXqpIDczD9bIp6P5WfhOJj2WiS9EODMbqAtFepLca7RdSK0dZ+pKPWyP9DmLtF7
r757PGo+5gW6QGc0e1bx+HchAcQ6ke38k0jHwMu5OhZ2oz5yTb9aJJfPCmL/reqA
JHoV9GszZ/RDh/kebp4pPkL2aWt3HB7Psd+XkFm5NiBNaoYlsgjcxgi02HMDSOuu
Luunx9Y5AHCEgDLOvcNm29AmRxOdZWi8xCuvfEpGSfKgAp/y52cFURUGN2KcRcBv
nwU4Z/+F40HlkWcDB10LXRaMYX5jpnWxHtRHNpEEsPyaUXu3uEeS6KuHDpH528b4
yyog8AyMQTSzUlNyMC10I7zofWeHYyOvQGf53EpKRnjTj9VR+IEQ4qg9U+SMT8lv
N14RKVckgDzAS7+lPP1pbnKzPqZ5EbgPklZZ8ANbsBeyi48Efk+iz6LgOTrLwMCI
te82blqNwY08LPg8SLmuvyaYJrhn+47QiR6+AkGOYqg8ILHNhYVoukkgdVIiuQMn
MBwgfnu7CXlCV9S/hBm3AX26JR6CFdlAeboxHgwzL1V5c7lIknefADMxB/iZuEfT
QLGDKif01kJYk4TB9UP2fRvqAqX8I22s1dmLBeIzpLmyfrPoGVFP1mKv9NZNt9kz
wCnrB9xH0HS8wfucMcAJcgRbxKsJu+pUShdM56Ko+suc8KIfwIQ2PTr3LfKapoXG
To41Dtd+a5m+hVoQ5ynvECj7M8ARiVKO3duNvL4cOBDwCsyb49hXB48U0wbIexI3
DCx1adI3oY3DbmHLV1EO7/79EKJeGbel8vjucBr8BF5AJi6eUDZkUQ1g+mNStNk0
sbpYXKoVha4OJVjsy1XzpniL03q09xrwO25CgNU4kWPKhAwM7yx+mwOfaXaAlamZ
3W+6xxIKjDQJXJkFI0SvX+XxJly5hvTj7pAXwEANmJNRlCekZz8vFmVeVZjHg1DN
ysxHMwPa4/WQC8Zx0VQ1HSZfdoypBlSFpoAIxFOJT0QIfCnOYVyNEPqtAqqG7m55
r3QkVPXh4zViTCoWE3qxbCLdrCRw9OjgKk0bx23YcwlDEZ7gnsLUmF3I93+Klcgo
ytSy71P38JO2nTH2fXGjnko133Tngf4dtEW29YCaIDa17UKJ/kBdre5qq6BhGmch
yx0FmQeG6VprMsHHRPM1GIKk5yaBu54ueRMq/MkJo1sbNIeh+rBN+M1cldIuANhb
v8ObfwmP3hIQIHNVllKCCYm65Hlr6PAeSuPIBkw6nPUo6XUz1rv4nw8+E3ErVLa+
kNAQlFcfq58iDoSorKBMWUpPisFt/avLaG5DFQxbo9f/58s38r8ZzKZXk1JutNKG
oiKOPWNiA+CYDK33MrHJVmUWZnzjeKvtcFQAZyVPLO6Eju3cN7CQT+5wy+l2Nqd0
rzNTcDZNInSqUtVgdP6akCpI86FJM9Ehtpqc8oIVCQCmjFCMTtTlvTpkXR85O0e1
R2V7AGPIZ+BDd/a202v1A/FkbZGGl17U5fQDjE/qjE5xDKTNIcvPWpoHjrcjABL/
R58zusn0h87gdeqRqm3XE/TauVmeOUHbH/2trt16I57YZwhY6gp2vPbljDXOYqot
HeQjQ0HUuKcn9Lxoyu7qQlbjOi5We26WfYrSZVm98/kiWNkQdc0pf+v8b1Ii9QOg
qUH8XhDuEVuUvHF7YhfZnAcqOCNiVr225m0vKqTs8subRL61r0fALdYuxrboX7t9
6un7QjxxuBGsk0w/2jxxDrUCXoK0CB7fDEJ5LpRd7/RpQ8XpnqVsBII/fFYlJl8U
kZEFSOAiCfjSdhJLJ3aJlRQSdHFQD+AeXSN7x7n86+vjCGExwcNy5/2DpsM6xYqg
MFQORuefxSWvJadjYuZkObmZapCqjqLh4U9feHd9UWDPnD27wfNSVyyXqx5mi4qt
NY+SW7rV52cE42qG73zULXxVAlATYW2CHLk9CCpUhLJGqx2ih6b1sfQIMx495oVR
7kskafoGWFYcFh+/3tPILtMcgX08i0vQ9vzXNXfiroMuV1/Nm1ToPzWs2Eh/S0Yb
5bVV6ILteNq9XdMy+zhIWCtJ0bBKuFIKbkRGn/opktoNZQxPetCztaTFZdiu0Fbk
f3a1nzbdf2s0rxshl1iKw9tJ46mVQzec/e9Fkxsjlhy5u8+4P58ZMmdEZpy4U6Xx
ghLrhWN3bxlL2n8Hv67RnYRCNdohqyJFHt4Fej2dQ7+vT8qurvtFrmSgWcka+2Vz
DprU/sjFFUZNuK3IiM/2xTkK9Ir4JfnlAG0bC6ULEYqjO4mpk85fQ59jBcQVMG+m
6VAb4nD7TNZdWikdecJPBLlfBYa9pRPqqjPyPOeW7DwM2ofE3V/9JNd2RocvjeN5
xbUACsx/iqvYLexQcYdJ4rIxJNReLYdiqg55G1hy//s3woRgwZrt08/co8Y+H69c
6IUtdvEKgOzPkRPM9ZcMkOiBb+G6RZmW7rwSwRKx0W6JzU6h8T/1ENp37Rd438I5
OJmKmDF2ErSN0pBvFFlyVVe/WSr82qCd/x/5nSkTgWZW+UIsbUpq5omhVzcBQMib
PeSGA5W0WvagcKK24CwOWHkIJk1RLMuGwMnWMSaTLIb4sJixcgjTy8fbmUEkXt5t
/pga/Lufs81hltTWI5QOM+UU5VYNY5ZmiFIEp/SOOPGmjbwRBk9lQNrKddo3r+VB
cpnB94G6UW1UkE7hcq+Q21Pod95JGrMUUC8Iq0u0dodBpw8kDpzSLE6r6GL39H/j
PP7qOX12ZZoAo4k8276T/4/XZWUG+9LYYeDdiC2cwf626Slc5ww4bHOVf2iH+sNs
aiJiceWa8Y0msiVtKAXex666uoYjrlEhX9rHoH+p8Bpx6Tej/D92WANOOhGgMGf1
iGFFiXoL3NAqe+4hCPmr70YVhx02DiSHyFT4rj7rTYYNIILM6mY9RyKQJYHBOOeM
YaqycET3dAVbsvbNCnPZn/x96SQh2UbCRdudLKgGDNZuORkOyc5rJB0AecI2pbAv
tQ7we3iSa3YdiGTX8NSiYm+rT5k+dI4hoDBMrKiRnbcHLiwb0qnM5APqsvAbAFU6
7YXdYKMyXFSzAlfpqrbd4RbeENWz8Zk1iZ9+NK/yzGDPt1dYTyPwcq0qCUGyuk8Y
0K7G81tG/oEJEH0qz2bw6j4yq5ONruehBeHdb0gICJSFNGmu+eCSMcpm8VVGpcrE
NU2JmxPMJAWpY7EjwOE3OmK9tMwZGpnGrS07AZ24q4oTJHuSp8qzjJj94R4erz0H
k0TqypbrRuo8miBMyZRy+GbVNRckSN4Dxo8Dpjrlz4h4q06ISzmLm7se9Hi0AXE2
1qzZmlxY/Vdb9S27y9Dd9ei93Y4mbF/JVrao5N0ltsQo2RaRHw9zeuEk9DFJ3Xqg
WsMmi6A1bxhiueiI+TIj50K3Yuj70cGx/itG6Us69ugwF1H7uixl1yFLNy31HFsC
9b0Z3m/9kfeDvkmJA0bGlp77o6BSOQpIv45moQPaq2O+CchG6oizBIka6Yk2LQQB
lp/yYjhYMmkVXQfqnYdzLrDT/qH0AmBPmYDhTx13F36jozKzhOSUCQW+31MUh7+j
N+ZkgMNVJ6zEE6EQhiTnMdotSs5ioJTRzmJjEnm9M7LIJA2zoEOpIWjsTqSWXz9H
2yRw5vWANCwPoln6BLsZ3SYPf5lkQjrX17QzzYbAU2hxML3Yy9H7wt2UjlLMGNDW
BSHUwjVeaFPSlG5PFNq5dQS+xKKn9epnBJuJ6G3z7ykEe9qYaErDTIaPXsGyNCU5
iM3a4GPK/IltUEQA+eQEpvfXjKQYSVOdAsh1nYaSah5lU9ulf7ynq5LLqg6o1EG1
3H0UN1qk7SYG0nsNt9YahIJUJMsSa2fRoxJzxJFDgW/DAWTHL+yusOST/sF4WCP1
dip8CEI5J82c9imp0Ls8GYBMP0G+7F7vQSpMrmw+keyyl3kRfJMD1lmtfVnqMj7I
WXrGKVsidPdP725J6sz2HmflbnhOWKANL7A3ecmvojpZUfodK3Bqc1n+8DwcSYoe
QtRtJJKE7iV1dlj42zXZpnrKM7abXwbvh8WiueDunFGaUvNAW13mn8rTC7o28ODG
vceDRPs7NtNV2A0v4AIZv9vvtYFk7luZZB3ow7SmyccP2zYENhf5TJ8Xk8ULfUni
ktnIZZzzS83e3EdUzTcA5LTyln8JuJpN6/VJ9JSVe/LxJD73mHglekjm3WXYjpBs
bATlDoUKADS7GXc7uxlhLcEawVCmiwtnPNp/D8PjrDcvaugG2q215nvm+fPxiZI0
YbyS1/qEqD/LfGljs6Ao0vbUf+xNaljuZvdvZ2dFEbOXkm/plNfLjzNRS6xDxcx5
RzW1S5Vy7909oipqf2eBYCmEBRMtF9lq4w2L0dUeLDzoWMWwsxeQ77cqZBsZ4wOi
wmJm7D92C2LvhydEp34QrLKichQMOWvvePNFaeClCg+Kgu8GDVL3t6df96iG0Rve
zb9I5jotknRggcpGaulvaxiP8ov+tRjSQtagVtV1QBF8pWORiu3YmVonskg/6pAf
geXI1fHTK9kXChBlpphxAX8YJVuZJFmMfHtSvARqAsLprO0jjMLnl6MCFcuQ8/Pr
iulCEdDjcxmfjMChjQT4wacpRxAiN9i5+fHtj7uAej1+2k1aJNPXq+8ans2S36cj
BAst3B+TnNlhrK00expigXazF3X4qBafsG853/OfogmeQOJ3ucdLUCHTf3osDBhr
Bbh+QA9RlOnQ21mAM0+pXXwsK7S181MKTeQHJ3RDp3H8AaU2F6WNOsHHxheE3kGX
yNYO0raTvCMiNsYIApZ4euNAeBRhhEkevBAVbc9ATgRZTejl1XlX71bhBp/iQo5S
4Cdw5gF2bbPLGnUp04Zn+dC4Kzqbckk+TXTfbN47xzHcKVAjxgCyEDlwjD18Vnmm
bi8DjbEsTiuLuTBGMQG7ipO0SZxK/eZTwbnm/Jk0ZjpQlbLwjrkj3K07eXoUMZp3
SuzvTBRWY7gwDRIQnhzK8V0v6NqbL+viOojRplbTWl+0L12Om9/BHxUbWCpBwIbK
CPasvBh8mhL7pG79ScyJzN6hluVcrW1ylhWXP3DYgok0D9qeXD+D8q4taZ7oDxSa
ZBCdg5wtG8+kWYLGoA59MSPD3BdafudlGb5uUGVhIxYXkGHs7kUv0LKXZEoJ41fk
q3ilJDaaMzYdSyWAeN+3C9MsM7kBrq27pGnDbqo9FXGjnv68ORgNB9s4mlvnTf4g
ffRFqDAS2WEvYUnMlWQBozJ5td4aCN3/TLqIt88H9pWjfcqT5Erg+Q3yDQrSBZNe
mrUXvjSNKbsx8rSDdd8+hYYo2oIXGGmk8DYeFClFhEQf/mK+ze3vPZUQBdnzD564
MKqNk9KyaJlmSlDs/EQQNt1gDsO1q8HzudK8yFzleQkWyaN/tJQWPkLxdR9TMDYa
juIkar0n2IzHsYQ/N8lKQcwjiDtUTDCWIAflOxiqTeLlQiOczElBLK1w7NP2bsHw
Pg7Wnq+MYgY5G5haZS3X9zTY+cHC3ARksLN+dirBHZwkSpMWpTrJKaS8VIpnfSrH
kHVx94t0oaVIhCtyKQnh89mG8+rkTm/R869409gQPpyHNgvqc6XrzUwSFuMvtb5D
G5SRoRhhqbSSz46wHngfv+WOfS8VW280HJVeaJtnAUdLI8KbGASqzNY8BrbQb1Bk
0mIpPDaiiaDPywgi0Y2wJEREqhsazU6ptvH90EA5hFXNzSy5eK2Lgp/t+tbL0laJ
Ctp/ctKnw/Sq7kjuuUczId0CkzHlsmfNKZbvIg80guZJMKuvnQnEsuWPabqAajdw
CLtmMbMk+8zlcgiiebcNcxRe+nc3eC9PGnoiBYXnmuZmZXfNVFQv3mY2bxhgUWAJ
9r5Hgf58LWq3E420MBRw7JcXNEuyD5C77ltvD5b+/VmHN7Eko63IBaX02I5JB1KZ
iPSth2eYa4GmSr8PJLMrqx3UCWU5hOE26rVtrOLtDz2PPObkhvs+1m8dGIEi/5yM
3EMyz/iiuONBsuJGd1497xwxO+pJB2mES2XVK1WD1wpH671DdqjFIJ7phMzGUH1q
NuzY+HUX0FwZiMkbieJO/j8STY0rW8EMBt1xk+xPYzQWtgv6b5/5CkvJBDS5trDQ
xGwaxAUInD3QZv1VUtkX/mptf8tHVkcFNNLXEqsizhkufuViu/pu8shdbXGMFqLJ
/aljh7LRt4TG60mj9Ycd0/b1Q1XF0M8/DcyBbJlZB146jAwcNruyAamzy7Zgm4hP
3iUFWS4c0BjjCQXrap/Ti4BGh5H+m155LJPMFajjpaWzzxH2WDpEF9Imwv7a8hYo
xXIS4vALu2YcfeXCsyBIubjrIk0YP+jSqnwfYVI3e0TUAzWZzHn8BdO89AvWZthv
q0w84J6nPcQcqTLXnvy9Q+ufEqTge6msG2lBQ09IRmcoMPxiRpXt2AXjMu38pH8m
3o1/2bc5jV/zs5fToXGt2fc5jiUQgMtk39Drq0Dh0l4CRXr8/hz3a60EEyK3qrYU
iNA/+yWBM+Z8WDILnuZ1VaJ+5LwDTzLa6z7wGqhFHLmKT/KiPiTNbADgrt5zFh1x
/hJcGpVDmzDLGAiRfsb/RbjHxr/LV7mg5UpIqmkPnrA+mwIMHbLHfKo88mUzBTvp
+4AhbFTAktltpZDv2Xud12fToEPlkK3hrX7RHRS5T3CVUKONybaNIOIb5VkzXOiZ
0+P3vTUCtJoRz/PZ5fRTPCTpJWXWYt7J7iVLnz7yyVyEHKg2KhN0Ek5xeLo0XPCa
9iLpXDWDPtwFyi2LIxBbQWet/5oABK8mixdnlOizN2c6ZtgA/DHzCq316rVTQppQ
KNzrOtyCg3zECXyuM8TrP8Z1PdtyT1IKGGe32Cu2fr1kT9NYLBrINihat7hJZT9k
T0FDBMXFv/QGGBG4NETSr4l6ujhMXF78qclP6O3hjUwnEmP6JH7elwgJvY2Wg8Sj
cXbosXKGmU8oruyb3pIHqgllSWlAumlVuAVqbonT95hN4muRUyWwPIEaP0yk2iud
TJENlGy4YL3YUIt8fYq9evxNxvToBDRM2o8pU1HhcYypiTpRl9kckfDd0ubm/YAc
egMja0iLoI+eHQ039qHv/yiKRgVgap5j8orHHnykWqsaqTgFhlZWfD7fAHIt6vC/
5KCUHwMSPs1R8DY94i1D3VNFBfZYouBzRyLiIHx7Gad1204h6m77zD3gB/aaMKRY
EKDZLmKAHi9eMuee51OO0MAD92sJTYUpCENcYJRADoEMl1ZTcUCgPdoZa1MQmqCR
6ixl9gp8q8SYV7MpC70sTK5natgRPVw6ZcjdQLtvwg0ic4pHgA0okt8smq3XIH+A
bPM6uXfvCOrqpGwuaFPbBzVk0x2HkiJBIPfEQG7MJ0V13v9784g+vwUcaG+o8D8q
mHW/iGMvG2YWIap3oH2DbqCPFuC3PMehn9ArIx9nznWbeoYJ1LjShsQfhVYS22c8
0L02fLTuMUo80eY7+mC8HcNiW7eGPfwCZqwjVaQvu4BRTqFQdpNj5owtdhVuU/HW
bivQfxJyJXs+DlonHQApCoNYg79SFaS/FU3PtQ6Php1qcz5+7NhczLYEddfNDYH/
tOY/eoynpQuSzOU2x6O4eTtLT3w5AHqDVWkIZjQEZ7lPNxp/qey2aEh8753bIpXX
uWMRmtDnIj3GQFdUir78cuL/ScwUNkvi6ZIB4G7dxZ4pAFsgN1K9L9vRdKK6T/lX
ojvUZ2m6iTh8p63W4THdIeqwVIO0B8Wy+N6UV+Aqzqg4n4aHPCQLcUBjWxa6uTLc
isHLd9hH/J+NbI2s06O06mtn1d8/+05Pht6c0REM8rD5N2X78e0zHPIazfGDEn8x
P59S5E7y46nXIUeb9lFLZR2h12eb+FDpMuheAFO7eWvJbdfmucVBD0F6AmnXRdxD
vikQa7N0AdIKWOVPc/aKbir6k7EqfXf/KRtwb5FVJGzCTIcOlX7+8IA6wJMAH1Zj
MsEIlF5IAVAf00nkniglArXDWbl1x2hf2qpgjCcqKrCRUB/cRsLd5McC68Sfbysu
0l5RFv7+RNrTNlDhR8gVpuldIy8mFdmhcYaBxxqd0mbMwNXbRW7aqV0u2KlF4AEr
bum3POzHpV6+1mAFfKgnqLOyeBIRK1pF30zf5R50u7dpSs1mVbEnadITuGVzPIHh
h7CetOhZJnlMADOV72kT0Gy6tG/ASNSt4FoUKLNKicfgXEC5GTt/cOgXewjxPMVc
V0CHkAi2E+wHCNGJXJv0R+wfqbacxJpy0gIA/+JUOEPaELrXVIlU14WVJea8RGSO
9XGrXqjNrceC8xHbD1TM0UX6+WsSDLoEFlA2OxTiFUV8nxubLxXLvzlKzPrYyJls
RLvSIBn4ohKytAbdSwO0EF2R4Wz8XtWUhS/BpNmC+xY0kkkSUhigjKC5KZEzgb7c
KNZlAnxjhy0jThwLqqQLxreMyPrLjRjPMZKJFqX7ZnCDh5qRKSIcuouNx+66Soz7
nUnshZ0r5+Kz1G+AuVNB8Ai7orkSUF55D+vi/A77n/npjObXzjYCl12aNAFPjdDb
YkHXzlqHvQeHJdn11ShVuuFspI2NHmX5/L383yC/Il8S/7iXgwGFPw9pcXDw5gtU
yeTowJjKtBBD42bf5ysK5dJYn/xK218G33e+nMl5KGZakeVFUu6okX0ULjee/TfT
OOhhI80KtXjTwzBLhZrmdGmZzDjIhEbj+qllWm+rOgYcybXBprZ9r6nsI701DEI3
NkKzQVrFRxwL2gBg/Ivs8oHQ5UZax9abgODm4MUlPk8Q2OI9Ki1XkYEhqhkhrB0+
gp8bFlDady0RIjL63VR23FWcMt87r1h8+FXOpB/q0or79pBpW4QiJEd2IeAimbQA
Z+iImfL15O/EEjrLh+xB4uwVIdGFIBEbO4gYCFGqPDc9h0xYjLo7f9w4pzdxhtZP
EDHpBG6t8Cur9f8jljvLTj7LuvT3vaTkbnw9uJjTfwNJ/2R2KQSWrbadWZaDdsVX
Rqsc1wl26VSghbMVCUiF2PV2SWfTLFKaaNcO6gIncK9D/eB+CjVFFKVYCKsEU/YV
KOxq3EiNXWIOhKepgfKbhtfQj1r8hHxgHQQLmyPhMplDsB0Z6UFfYLqRedk8Dc3V
g8S88nqv3iroRirF1BUp8t9Amto84UwWxJ0971wyXzUamB2E7ESnRrqHbTT2b/dc
cwuUT/HEy3lw4L3Q9UpOWYZwz9S376tPwuLRxETqrAROtPY8JsN3ioUHDTxrFCy0
qVkTZoBNYByxULFv4Es+1iK+P21JprEV16B2f/uE4pTZ0s2sKvVzQUz+/D0bxdwk
cqwnlMpCchRV9dYVQMEo/YzWM3Q2iKhmhDSHOvGFodBZBozzMuTKrUpEqlHqZmCQ
tsdkkokvrLkcDOJUp0SguwXwm0Z3mYRxHzYGx7X6dCxsECLrJBi7E0F+1AtA7LdT
DJ8DoYjmfnijAr5VFs6aAgLxfpEAFGzKsZgEcLx9t0+/AVtHJ5kp45gskyY/DhtK
G0X2kPVLVmunEUzWu5TBANrJwkye5kCf98J4l8J68z/YkObd4vcVMm8fQMHqC4Nh
DW6lVr/mnahHiWTbVfppe/h4DDHFG5b0uv47Av4bng5vih32TeiqdwTtzZcrZE+7
+1C+BjL0Bso89VuoNF/Z+nAUbOU5gJY2o8j9251eEwcCG/j7WFQJprLGdpg9+QaT
WwXtdaLrkpPajWKywqOFTKlKDiSiNIaMzbEnxXG9VmR5Jgvix5ZeUjBVgLuPoXtQ
j2OBgKpzHLzZwJU094NwmAryc18ZJOSRSYExWKM7YulBaaFA995sT2oZ96k0eenV
GrKx7s7HtfWPRM2g2WalQxOb7F/ixYPX3on3svKUee6/4DZidPzBje2py4Qb92j7
iJ77JXkLGKfasnmxaC+KYJ/iF02qtmlMJSv48aiAZv4Vpl5jiyodWS76cIh8A8N6
/lknMm9TOxRqNPHy2ZZGrvozC7XO8oVvkpUfbKcFX+Onm3cta31pIOQRQ9hHAFiF
vh2uKRpYe/hGIIt1fh2nESbKfTRJUWgAQDJHgTGv7jj+45jf40L5Flmkc0cRCXRS
DafsEh8dYkN75xYHZlqwMRwlOKbXlKL4GZl5aKsKrUgaHVUJ4WJuwkPePsAt2PnD
VXBA+OQXd4o0fnfkqnEYZ+7wbcKq0skRS/DJbp2oBSXDlHwB6uc2PAncjGWOo8Pt
7wFmrGLYL2J84zp2FeJLRNvwBWm8Jw1cT04qqOzcd8ULN/iTcLb0odUPQwfj3MS/
1iPA1kIJMEtpgRodpadg/NEBTtDlnxRhwCkllKyVnMvmS0o5tl7q3PieXw+5JPRF
FFu+mieHHQVvRsYTcYI+mRTpEvF2ju65bmQcF1Ca88P8j7WfVG+c/YO41HYqS3ZO
vxi9ZOLnPzQ9AuFgGTFFHQNMGTx9GNHJ3zrvt6uykaQZQt7i5HdoabCLzUkJtud0
N4q60l040j6b4LQHuHHsMk0FPxUCqMeD3F2ssxu0dldFRwdA0ZcsHXwM/pRptE4J
fI2ptRHv+2gtn+RjXUifSTr4TOhErVK3SIcxa0l8qX1HFnCdoVFYs+GFLmDAkSjB
pcB+jmNcuPJR1FpSRfxcMXGyETvRPa1aMdXvSWKH8O2BHFcZQI1J/4xdtVDQ/8e+
5GNWI1Fo5/5urwpV1O6vdNsvN6bwYPFSjGCWBiCePyWavbI/a+6BmENVv7M1Cq8C
zSyqomT0N9LSI8nXnoXQFsQhVLhV456qMzutPV16AgqhWUrRHwUtllfR1NA9OxQ2
CFnAnxiDpNc/BhW8u0joj61iPQStQxhAenGX6VsaTYMQtHPzBb8J3Z03codPUb6s
rWZouZp9e5Bwdk1jXzor9riJpCgn++/oBkgD+UYcDMluXMCnyaLqKuMFyFl9Is2x
pvXNmiKfeVwOG4xhz+QGcAwCAlF/zAQZ8TKp0Yxy5w+hc112RQDTE1YhclAeAx/N
n3OwfqaCyWw2fUli2cwyPrY8UbW4eeqHixB05FZpqdN9p4ThovrVHEHKTEUjl7ZK
0+g1YT+/wmOIsn7MIcpvu8Oi3M7zGH6MZTx4zvpvRjhuA78Ey3rt8/o4FigG5MWe
1M4Plj+GJBVH5V+SWUT0OOqTH0GfKqsbYuEBSw6fR3fVUIUs+vXyv9jPIUa9Q5KK
i8M0zkbM126hwBK9YGkHNC6eVTJC2ZxJ8rfeoA/oOm+kXpzfMvFZNDH0/+a7ViUV
GmeZwohrgvg52BUqjhcNdG5UQvks1I2f6zi0ix059d92PUetFhImZpprssWkgft1
D5yQ07Z6yi438rfByQjSwHlOKsl0x5XE7166a5vjqa+xbAwqgW17ViufjeI61lc7
grUVdoJuPiRPg4TLhU8mXcrJxzSeDAbXR+VgvgfKTHqEALcHvj80khVGhQjy3Vg/
TQyiTaphgX2Xma1FVg+XM8i8859708SCliVOxFaYMMmcmEjW73jsRwGLLCjlj8nC
HIDRA5hbrX6bi5855g3tjY08DnC9Y2yD85lA5CdMZ+L1fASe4jiX+M0w+SGYgo7/
V6W19owOkbDVli7/lke+inTbmzO87iot7f0fSqWbatwrHj+Q20AwFg/ZboXGySyc
8baMb89w/s4EYYhK/cYiUBjEQD/nAecW0AZSsPXebNcsbEiidy7WbKLHvofuUkkh
IepisKkpPKl4CU/X8e1dDdZUpAI6rmBTaJVb8DlVy1RUCq5WpSayy5xXwaLH+XF2
DL+3KIH0WFs9f91mCK8x/2Ajn8pSnm/MiktomvCBexTfqmpdOzvbiLrG6BDisR8n
tf7jt8vNqDcfbc//f7b28p02BySHbaQOdslXK3bksnd8ONLdvp3ryRbzvkgDTMDI
VVTI8xYoDFBLBx4TI82i731ZARaGcn6Ci7ZvFbPJRXWQdSXwWymYJuieoP71xzK2
dRCbVuX0/PtSGcOk4eE4KoMJsytBx5GnqcPBC0pXLjYeYk3H8Syen5XSkuaS5X8a
zdOVFLE4QM4z5UK138Hz8LJ6mXCHrBDBBukurzJ8nBvp2itP6VTecUxqBsJ34u7J
JQlGfpCe3CpHEiyka5f596D1psbknMkd7XaQjmUWKqqX7ClGEHZ/6FOIcOY+Dkzh
KNDw40txiJpS6SGEe4wPmXXgnjufk/BCUbeaKlTFlQ7nnxEu0Wtdm8Qmz/BfNOIp
jgULLqn189IPmRYljl8uYQxFhzeHlh1eDBodJZCwGMgO/LkfkNIFhtcaAubMcFi4
wc/IgaVl3dBwFIHbRek+P+rmDltp+BCu7Ngj0otv/HJHBUlt6Z8eplzi9HxeAAyd
p6uMT8K3/CyCeUJNTYAhtfVo9AVavF8EPXF+gjFlmDOYNAgF4W8znprsDPGSdPPO
viySWYSJdDljnDyyz+PtN1xggrH5H1aGQbtx+++1BajmU6aeMr8XZHeaSOkj55Oj
ywwxj5yM1PIPRdVu9prbeZpmWjAQ7ahRwWE2Jqw0rY1dFQcWR0N6wgjGxgurQFjF
1g0jWSY6JngMygdJX7mttmvjDxFwb1jbvRZodM210p3ojvIdwznJNvB0zE7w0Di6
qSb7gKB/9Yef6ExFR83/iXDMhENxUyvia4KMlVvpuG3/TS6JL6ssApMhQkNUsX7y
F64O5DOHXj8oaHSkR35fZzzIPtfM0VwxC+urBDLSyKU/6kbxJVWiC9YlvB6W83pS
4TDUiTQiO5outuULa1Um1j4MMuYs3EOlqIxbhrqXe2k7p/27M4/zRV09SxPKEP7j
Q6+vNkX/EAiKuB5KYZ/0EhdZIcbc/VweqV71xVTLVbnyVKJl8uSc2nrMyGANpgtb
mMo6SG1bzY37c+rN10go1M52zvgmyOrMRUlI4d8sHsoJxKnhyyAPrfSDEcfsZieS
MJZVnJgFDVR9A2f/TV0bxlJd7b358jiPn4epvXHzXGND0A4Pnhm9c774OQC/oRxC
gFhyUb5LfYnyw0cshdE+sBQdgC/Vuw2sOp61tHn0Jx5obfTyTxAI8a2P4GbpuGsp
900qgPHBanKsYaRFk9pEgTttlvwR1n0DkxYNYlyJHa2Vago89jxcZTUQen+DtybN
Mbn5ec0AradVaFDDNyuvc34FF7y1hUfAPR20MNsvebzSo6sMDf0A6Ah83z+E0o8n
kxGqRkRp/of6w/znxvatmbaH1pEQpfZ70bKaSyffxBH7QZCHvxHTXTJUOPLRARe/
Ht+W350S0gS/Q1Bz0G0VIc3YUGIQH1cxkck62YUdeKX4NE3NTwUQn8MbfAlLXTq7
Fs7WV59fzhzk+tbzIFhTgEBbWMIvUXh/JDqhQj8aH7COvVRuH78gB6hb1brAfgrl
3fCRPwmTyqaEwYmNkQehrvis85E4IMK1xi8MR721TP+JGWJsPforR8tCsBLnyEoI
ymVzd0vYMqZ+6EfnSmf2saaiyP4O15Bm3ogmsnoaoGxUGVVfP2eqlZr2Xq4+TG98
XW62mwQayH2lzO3GKmhQUyP5oODCO6TRZsiyi3CseijkykBBIWMST0FO5ilOVhxE
ijxyPuXNGBIqb+Pr7X8rcvWncyo8nmd9e17a3863pLhZoz/Q+yfbUq+JZvLEptwJ
aubSjrSKWlSk/I3XLPHOhDneYvzrcb1wGqfjlHc8KwYlwOJwbW4Enn1ORGRF6hBv
pPRqmWC5Ak5H7djuEiwWR3lkXiLwqxzoJr1iKGFcCCNIJbiOc3vVGN5R73BR4dH4
IJIKxYXF4dUhpt0ycLEbGmtUhEdEIZdkZjC+cZ1+Yx327E62NjU9yaAy7DEghQ6k
QUwLx/+7knkKY483FfLRCW8qN0qqGQ1qrAwS1VG+Z3xlFgpkSljtyus1RbW5/vOK
9EmPQFcjzT2CjblzCwPIJe5KBu6xh6KZlZjBGX0LoOpouaySHcGrg3nIb0lBxprA
qHISrjk43AIARgUt+FIvN/FpteIioluBAvExvv0UQArQu747kLITErLgjZiWC/t/
eqZFb9Bc9vmJ89qDm+5S7bXPsHePfhxRx6pKUXtpp/wpd9gO6OEy2yNUriIMNiVh
asKwNZcDomQHPE4iW8H2puV7L31aAP6X8VQHFVadz4mu8nTGVuzfaU0sYGynAg0i
inxReBBoQpB7lxcOe22Qzk/s8a4t5GAwQJONE+8IlDg0paF5qE3Afb6Gd1NpV8yw
CrKgNbEqIAxTM65QjUAiWT1ExUhfoIMts6TdJwFx3jnzlMmSDyRdMcgE8P5K5iZP
LM2T0JMwPT4x7in1SoTFHbDaFTNS8/LSwtRABVLOYK6k27E1B4OZQgZLmiKgXwGu
nQdeJqPtzj+mKJaTjRshazgirQxxXFwCwEurxE06526stv+b8o+Qvu6rX7UhRYkn
BVU1jjv/p9LUZajQNHGs6lPxXdlH8QJqBPQmmPNfEyS8TX79WMIAmhiaYos5cWr3
UL0mZhjF3uGEjy5VhBtJF8OYyVHzBLfttC3tK3BdYSyLLuYie6YL591MQgrvcVCy
Y2A6cvcZYRSd/YCmW3jPKYjQEasVjcD8IidmiuWMwcjp9HL5UBlD1t54V+NmpS2e
LPrhPq1zR1ePre//LICmxqFgxiK+Z7R9IisY65ZNyxgm5gL0UqzewY3TE8uvba2E
Y2xF9R0bOXYrypjrFjRN4dzt628qxN9CR+2mQsdAfNzScGgk7xkPuBRCvtfzsHp2
xshdSYTB2Oq/iAiQMsburzo42Nw+/ddw4Sh2r5QCymFBaA7l7nfPy1cA08/awSuk
sPcRsoQwoMZD0V+c13fW+Fv9IhIGXAlRzM9EaXQ5IQMl3NL8GOBvnksHNsnfcSWx
wqeU+y2wbgCECfKgB2M9lwsN1jKYYE+Hg4CBJUXFgxzkfukemjr15Nh0hONhCRwk
SypYyenrdoiZwJ4U/rJqp22Fy1JWSrviusQslye1ytu7uJw82jmxhae7Jp62jyky
ZztDmBdlaWYUJ+i9fHW5X6Lnb6PFQbH3WBNUzvZk7WKYre2H9EbrR+D+qsOB0sSY
ixCYGjyP1cBmf8idOTyJ4RNUEyvlrDB4f9fnlOIM46fDQMNgEi6BimSvzfP+rPSA
f96v1PPPKMyP7in8qoiHVRSjAfgekJRS2zuypWxKZipC29U5hVmSU/eQ3f48Hmai
cLy14VCHKvk+UR4mGnlg8n8WrrazTVF0MDuLhNMetpjlIHXTqXBC/CF9aNS3e6GS
y2Di6nUSptBUtsXzdreMN10x/nBLWzUy2GLhSMkpKNSrZkIG8HV11X+VMsS0SrGT
KpJQgoNhDjzvIutDsHMXn/PNNdDDrnJv4b6TruOpgYszVmhyiBd/YYdeGj2N3cwl
ynk8TwyWzxEzqSluDl54gkdeSylkNBLZ1vQOvxGItW5c0/fJn6m51zw0fb1nShR3
o3metRNvuqEd2UMUjo6vKuaGJ36VIpKBkR6nv5iKxd2FAtNrpJVu0Q/9ND5RnhwX
LqxSrlWhrDG/2VakUgL97PJJOrjxtAtAb3CBoAwI3GWvHHwMLsWctARvyNOCzHZL
DadRC1Go5+E2CeHahmVK1c5dMZIe9aYk8VdZXlCfhRtgfXdgcBSyiisXMIgin09O
Dqh7bP0ljv0efGtxBx7WR9N4lheRwOCsFMxdP99D/sq7suLopLBD791YijfnsxhZ
20XnXmMns4HqYcARGu9Me/99qNK8ciIld9GWlTuuxPCcKwY6iOim6o9DivOAIdUg
fL0DWmluy2XL2lcU/j1zTFvAEPN248uXk+sDaFedTAc/BiVWEtEwWigwt9S4/Iih
Vz3MZznfFDbFmGL+aRkNylkGRLABiR6RwNZu/EbOR9UncZOMzXWGBcVtJS0v6hKM
E/1AXwhheFHH5MlhfP2AW87HUeflOysKrHr5GgZLXQX9pd63gKdd7xcOrNDrE7UZ
bcQJzAYKBw8bJVdR/rgGpMEVspRYt78fUKCyoQCbq+cKMS4VN4XVAz77KaR35WPG
oNLcxD9dazYUQ4sBssbaDiYNS1mrooI6ej7/jx3IbG6I/jXdfFJEHC5TEGKG2nNR
Wj6uKnncaJGIuBpPSjMu+uL8SzmiW7L/5b/5iKm3CQQ0M+K+CdReuCfrZNNKsHV3
ki53Quq++pJRY6PuwxY7p1apsGqq2Mt2qbPIjJ6hEZD49RSk/jXgEMJzzalSxlk3
nEq/jltQr2OSMrTRbes8Oj3EshZZ5al4YEG7xtlazGkGki2Go/iFaSyFFDiumBu0
/JSoY3zJu64eWrvA2ypCmZIMihKDwrmqUIxLjwGZzrs4V78Gyz63E7aE18/URYAL
NdNTFo9CCEKmwAExMAgKruVRNj4SAFSqCzR7SvpUf8Ut5NpAj798ofrFmLhdv5FF
W/qL5MBrgRKzOZL8GFmtfq82m7SRg4chTJik7fDQkfzWW4XrnV83AnsgPHlTVE69
8/6EwHCDpFf9n3Qa/oVRXs7ozUjKopgd+4x95iUb8XlryMAFsg7ZUfLLU+zQkXMR
x9/YuZYk44SrDJUYDAHVoPS7OEXv0E4cAEVFPBiSxRWy/gQ2BgQVM2RYL86upbJX
1M30GKrV49d+8deLVzmQNpK34ygKT7SZpvbwmTQ6JIVYFi9fyi/WoLz7YqiwafKW
YsdoukU89HRxIrGjVweWEpRx28bgWV7NrZuGbhDyaom7TNYEUIXyqV6jglTlaPeZ
49x/ezve2jdQ37JSg3MO0Q6zza8/HJloOjc0n4H8ggT6CehkHk6ygCQYwFyw8HpB
dQPr9izxERGwJpmMLO32AiMK5rFgPc+HBbXEVT+ZyXEhRDHaYhWIf9BVKmAH0p3+
W9I34yBz405/qXITraFNukdBjz5G4EirojiuecklJhi6O6E2J2XcN2MjebB1f+Mt
q/k2YfeQtNNMrWYrVZ2l9U0hV1TsGRoUrYTeskGmMvc3kaGR1GQIrQrZo3A2pbN6
VNMYO3KYvumGn65B4hOtJia5XijcXm5c/K7fUBCC7+cd4aHktyYYLQbBRRs5MgvQ
7pPTHvLfV8nk8nS/01ye1ScThKxr2qWNweQgiiZkvZN6g/6ugtlhPOoEt4XCqlJD
dbK6ZojKzl/bVEdkH0II5P3c8lDCSGoyudnKKducOJ1FiH2tdzDdWlLlXKgQ8tX9
KJuHD8LKFZ4TwOI7RukB+3Pwb8qNMK7OqVxHsHr/7ozeWXIe55kEhYBzvi/KjntX
PBTHtBptq+VJ0IYaXx+cka89gay5MZR3XSjDrhCqkqIbidcsBGnkDz5kM07A1xkB
r6yBEE+piA6UEKVkjfY3+8VJHSg5t1BSB+uIIUGuGDgM7XjXfkBlTqQPW7Cut3iJ
72stUe11E7UeqbNb8SgNALumYqgUNdr6pTMu26IsyDH6DXIW9CRBFXvMmPGQJfvn
9B3yavXjTBWaolvwKtNr1drXntL+fXcORXp8FuyhIrSI00/dJv5vwR5fisjAZYfF
ZZQzdXnPgBBfz64aLJOU6I8qqwfUVksuze6DJbN8pRchBiwNxdfUYp9XUOJ+YHrZ
Ol+b7xO6GdyBJqooQByIeq978wlUgDzAGavLwURgCIX4Ze5JqLQsFxIPAGvzUgPO
b4A1zEk34A1WAcxYBsINGIs359PifUZq6+2GPSY6RfmONy4RA9yIeWbmzwWQsy/R
AeD2stCX2f5b7TOcKmWE3ngYbI0q2w8kSbrLAtLOO8IzM8BeoU01Eu486sUcyCu7
8+jJvAjQWktEYAAVLrz2g2MWo4HaSWX+nXnzcxY+XaVLYb/5xSpeuTE1b07RLTDk
2U614dNhfPu7rokkWam5vmbxSyO/fckz4DZHXleWAC+oK6CFw30xtQcW2OBJstEw
L6Pm9XThKbotbSRQ80gWtLUQyutXC08Fu6vTEST9ph5zmv3jNHfIIr+f0o/4JuGt
jk3RdI4hwOfHNdQhYyq9+Y1Om5HzIynRAH8HC/nBWzKod8pUOwHmaTzFWlCB19ck
G4ixLOAMou0AZMlDkFvj3BSKG0qVPJDo/+CU1hkHgdIFoxOgAWFYE3hDWVIUYmxQ
yry/urAB9N77THzdJxxeJ5lA5U5ZRffoXH++ZHbcvMBZVJ4oNwsC+nFLW5aWK8Pt
0y9Yb8WxUW+QeOSH1syENGkItYSZvVR/8+8j/LQrKGeoq+8uy9dvtJkUkuuVgDek
qkNoRcXWDkMm+mcj7BFN+ZOjtNZLHU7oueyR0gpXtLb+ej8y6DkNTMmZTWn0rZXM
I015/JhGGCnRsfbk70WuWVlTjqZ19LS+/Xs0QV/z0mlYo7apz5tsdzjkiSNHMWcE
apQ3ChcKHP/qMjK7vpnUjCcwRdEPSIIV7Vvinv7m1grbe/JDFcqnITc4rkLLyGLR
6/x7bO3HLvprlhU48L+OWufGEaFdDUk4TxSBMeeRikDWuRVhG2chtrYTXxZ+2EZV
PDcUVAr0ZPSKPjeciMvKlkLP/N6gXxNyWLq1Ivmg1m5B0FDjwgY/Zpbt+NX84kWK
+aSNca1GuNqBSac8yXNAJbOe2GzK6OiDysYz2wUSjE5acHr4iMXwlA8iCC4e0KH2
yqfoRAmddzc6wLoM0kAA6Gaw046wqZwQ26Vovy71LOdB+oNYAksCedcCbOI5hQ8n
h4s5EL+A10iUGEYmWnuqXjNwG47k+zedHigX8EOP19vMoQ1h5KJhkZ/UF22MoV40
sk7P8qIqa9idijaZo/sR+O3WGnLNDJg6lME2WMQCHOfI+DzWpP34SG8Fkr07k00W
xacpOGyEsFWm7aGi+0xMvV1BTlNYNLX1Z6xKpNYKlZoZLzUcqYETiaLqbdqI2j14
1kKEWy3rwNmuBcG7anOQ6apBVqC0yoiYUPRAczkbCObAdBvApyxW7/nACn4v9yWQ
rSNHujZrgCGc12FPQX4gasFhmXpmCI9Xg6TRjWsiX4bZcrkDmypYJzP0SAl9Q+jP
FUSvXF0mTtI74EenjZcyNasMqBwkjhVsnPvkKz88tyOExNIg1q+jMwnrhvQZDFOk
XoawxZaYlKbHT9ubyxhNKPG/ZxcTh7+F+LhTM5ZWrAfDJ9G1pjg7VSAUyJmfHEzG
L6M9BJlkKrqU6NEv3LMpwqnQLfPGMfDHi9WW7m7yrFW1to1KpYpGFgcoCWjHK9QA
QoVPoKPGulxKMz9mBwuxBiYIr65/uDMrxcNAoN2H0JF/LCifhM/J/Y8M1p5QMmN/
q27Wt6bPeQ51jgP8+5OYxDB41gdDMpNwYid9om7+haGpvfusutRtZZCYsToRZ7oM
qSaoZ+C1lWOb8B6Qqqpn6ESXXaEXwt4HcpCdxzBgOTuqbGfG4mBZbwARLrLbiqI8
um/xy+9v1UOh+D7jL093hRXlndg44by2elawuuRN324oJAPwgYWJQcLWqQzH6Du9
TTM4x+bzpdhlvCTxmkqeiCTHHj9NpgmF2but54D5dxuH/CZ908PzofJwZitbjeSD
mcJruRggTG6crNFDMZboOeMZp/QMAn4GGVW57h00VJ74zuvs43ZEazGOqcDo0Z6Z
DtHaEiDNHesgPUiLm2U7XILAzeMT8dip1e7SeYQTuADkTEep8hNhFX3fRmFsy4VU
eR9Uw0XFLkEUG1hjbwD2QD6vwWSGNb4b0nVDG3BRXO7iqs6pZ4+avs6gAngPa3cb
KgUKbfriF0YaM2drKI1heU20qxwZWOvbiMLt+FZ/zb6xjaSbq8IKdTsvaK4hhSJm
fe0klZnob1jf8yCNlvCC/tdgdiRSnyZ+Te58yCJrXml1TIbhLhLhMRl7MLcyUg6E
er9rvsS2zZcdZwH7YGV0RtZu/mhbmkD7uryZvmw4FK/OxHT3tFoQIqJQA2knUOSl
wvP2YrkUVANAWYWCJpM6f0vrgRPf0w0Owg1Vc7P1F+OcNgBS/Vth/Geil29kgwWv
RF3pTmfZwbiTd3yTL0BJ2GuBm0LKGKNGyAvLtqE0Soeo1xi50mpryB7ns2SOPXAj
Rga000S27h0+NtB4L/VHD+e9VhDLv7o4CyD9bi3ogPY/OHh4PvjuGKWANNYh5IEK
iNNrtnAzwnqTh1E5syszxv0jycuygQkAIL2vyvmwIRFdKY2xMUS4H2U8AW80ffQI
JIX2QQM6guUp9koEiu2A8tkaGAzMcv0wzEQufKdOyMgmbxmpUNfr10jdAvoOseF6
IYTDgdLBPULR1gaGgLC/nyxBvWbMdIbtXGVvyfVJWS+QJcxvshDrcvtDzt/l0JA6
Ld/Rdvp0+FwsSyKiWWfi7IwpASwI0r/fp5V4JYGhDAc/+hxns4ZT5ZoEHJQSo82c
TGNuDasM7ieJ0e77yYuC0C1JfKnQtEtKHMdxWZ3RYm1wW3gNWUakOmZNILgsdVRA
tySR4GP2MNGmGQxtYmacc4PNyJQ5GeER3vS+UfZ0KVrpoGazFpaBx6U+SkKQ/n5A
2jR9dgRUoSdpthq1D5ww8eO13HFTs1bZwNvoLZ8o8QTGQfY34xx6lqHkHmlmtLRf
TQBG9b4I+ZSibgKkKO0Hzj6N3jL++QzidNHy0ni/HK0jQHo4DAbLwSQoIsNA9eLx
IyD1yixsoY/rgRNGBZexJxMGukR6yZhHPKmX0YnhN7ZPeQn4w0kpyWF2xKY8vBWM
XJORBnO0JwKKwmXI949hMYjN/QAaqiIIjVTvBIKQFksNs6M5QEaVgNANyntdavC7
mdsFrCIme14YWrP29//gN7724wxZ6XJUOATC00qFr4ZeYYwb7/UFmZomuVZzbkMD
R++ASb9f2KhDgMczdcsW9AzgvfuotvKgv4NRPnsxPuR9+FzAeyyHabipIwn4BWB6
QZewOu5npbwGTYcOqPF6/kP6pY2IDbZaGE3yolJjLqzVYVTKc3IlWIkMS2mZOe3j
0vu5u4Sv8CaABPlMEBDpXmiHEibbDdWxVk72FGTIWXaiY0+ByDUX39hddb0uL2tv
WNyZJ7BH+Kmnv2oz1F7SXXXmEk5jqylxNvKzNoEJ0CrnqS40rsWdLXcBz6v2fvbp
CZJ7nFrZeZrPfaKa91CCvPqZuZsDJcj1RmAEvtxvFsB+aA0q9PQQEAlTfYqpCTU+
ZFbWlmKp5wPSDZfEv9FX25TUsH0iZQrOKcGQotlf5+NKGeKWOgUH+thb7HUK8Dmr
Ub3i+lPHp1pUV8pCQJ0kXJlIQnasNnR8doVf9A69RzSm4+y0U3RIfR0w0s6YhOX8
qzmQ368xESes4B4WHHZm3Mz1km6zO37dOpvzj8xDdC8wLPKTwxNPkZnN0l0O+1sN
X5+DBQSSptfpZvmrjQCvmkTincJijSau63WMyc7ey/Mt4+8FI124IxlCOoWu38vs
h+vzOaZQ9CQuLU/JQb6uEyxkaLYdQLzSwP+GbGGGoPK2E3WCUFxSsG41PUfIAUus
iWtCSNoznGZcOIPnsJVL6ICfA8wBEDK6U3BJGCHJLxI2EUCUrN3egnPfXfdnysfQ
GGoLc0dgGKJsiF3hFRdmN4XD/J7dyUeJtpTzKw2JyugY1y8JC2LQN8laVUexc+jE
o1wVmqQlXCWSA2X9rBCuho/gBIRnZbQ0+rUN34aIg+c21JZdVY8opnkEZm5gCOn/
NdWPpGIjiQ3Co+LCQZ4W7nt+1zqKneYeT0+PZyKIQWD2/dFQTbMeWjTc4My1M4NN
2x852s/4W2jwB7/tFCOZnvln5XoUw5wpaKxKBUE2EXAInjaENd68gIiu2RaDGqOe
lNRYRDsKGbwC34NqaDAQQvBFQdv5IibIPRwa1oigSPLlvebJSQ8SOX6gnwPWfcMB
KyHqZF3pzg20NaC1ZPP15SbuIsg+lAEB4u0qUz+zbOf8CRA2xEY6xW6YQMt5W5ma
AajvRZrfdZH5r7DlPERfSzrh+oWqf7suDsnuxY8ubXZiumrqjKO/uw1F40+ivg4f
gyyMR5kE2jk3vr9UEoWbhMKffFK1WPRr/2NE1PTp5BxlDdtyR6c3VNKKFamzSI9U
sNf6TT1hNgTXuf5YTmOgZIZg579xUeQmHlxlHDjLme9piZj+ugw54PCKqlzngVLt
qJagiO7ZDLzCSVlSdYEJ/U5CPw1hBrXIxtJURJ/SCt1vwUPRsJPoEoQv7uqdxKtj
FQ+pQBCa72FQs1gDbUYv0WpOB0hsnpS5CRoxytd8SV4o5YllOqMxf0bJSd0D76de
IpOSr4Xw+JvUctcAZk+zH23OVFYco+fw40VieArF+FY9Y3mw0BV9PfDdOARQG4S5
fIZFUiYsUHo69scznzdY6sj9NaAjkif2PMkZVsGesw28d3k5r0wQDo0C0NELFAoG
xCl04V9PaVK72NfNqSoEPRJj3BxCnQ7xl/KceuERG4gdP3xUpSleYPTRuNLSJHhe
dxaXKdY+CcLcDbLn5ECPWOvk1bQ9grtSYtfEHcM16a8+F5W4XI43VXHKKIQSz6in
tTGHWvdEQV31mDiMqjZCFj5+tcCYEQCuAA03asSA+mncLmgpcCXRZ8uugbWxFfuz
o+63/G4biJ0uDxPDZk76uyVPJTN6jCQ6ep1uc8ZMnh3rVI6nMUlepTYVF391yp0M
465udyCy//siC5cMaxqvx7lNMvrArKvE6ysuBB7FNW0AfGqCZ5Ab1kCkSNvhPxwb
b3tPPiJuWwFUvT5x8VSrJV7pxsLdAVgC0JIghVVwqU7X9ndwDT3wuNsyiFE0J0eh
Xzcx/0KhzwZ5609v1QDh2bsjIovyInx6gkv88wYr3IQsmRCnV5I1E/A3oqP/0t9G
6xiaV4nxYjFIW6Nas6J9vjyDv8/v6HWSKEmP35SQV5y70X0+QO412vjrvH8u89JH
/c9shcKFZruCMJms3Av2QZRgy31Njh0N/X1h1/vFQMVT9yuggWGnj5rWw2jfCQS2
B+tPul4M337oqI+Hr2L65RXbNX8tqrPeUqJ7JTF5XVTZq/D4tWEBYRJIyqbRPdM+
yosxnCNiF9dqfIMcrW6+76MD8tu2b59zcqWvaUR30QfH5sYki6JRXLa9J6kDd6Oq
oA6lBwSHLY50sfXBdejbABhNCp17FmrwJ2lPjFQk4zbyUSaxZC5e/USHawVXROaL
aB2jkGEal4MEi+EJ7hC9mS6SwAeyn3oPs2ZWde0cVQ+mUKsVIKPAiX1IcuM9skyA
fi6bK3c8NeFCgmsnQT+uIZ6iJSNgmob9hWkVZhVashLOzP0fLCkgwyzoN8+vXL46
NM6Ukror8T3pUzzqsup/rw1oWl3xSgiJQpGlEz1z7ry/movlYNCPzZF12ILZ6fpB
vFGh9EAP/qcmzxzzMAfPaOX8JOA3SBhGvx00JK7UgSkrLLSbNsR8xOzyqm4edV/N
g0hg0QpJVKqpJHHQ8bV6QaAmMlh8CbeQJaNGRVOfuritcXJi3w3NYfl691BSMEqK
rwURqdxG1qz8svqROpKLns1yniKDA5BrlBT8CMsB5utDVkc43aK8lRNhBO4CxxEV
JJyQzeJ11dlusbwBJ/FgR7GFL9wOdYzRqjh9gWWlnryMQiw0Uf6e23KxCUn3t0AN
EB2m5WejuYUlz95PbOwERWJ04LKCjitXpiQu+HP7KQ+H9e4NR/ctg4fJINjoxz5M
9qCIolrvYFopu0inp3W/lIlMqylZIraV5Uj2hBFeePBHPSW119/QlL+NvdcbvhWE
7wS/kP1hnGu0B9MHEqmY92DclI0TquTyR2CHZ5SOXvNoKOelMxBUOVj8W+alTlVy
z8CKVCkGLieAnqLkeLVgzxVzI55ohU361FAFd7uCNPGBK3vQzb0xJmI2oZZ2Lb6f
TLeTgBwqOAJSDPQ+Ao1Vh0vozGNMv29uSEAc4Pq7sA3HnvrkyvMKkRD9V1QjYsg/
VqQlEUAlLzkyigxV31/bk8jDDS5ip3L8uhld5KkSwyY1osQXk1Qv360UdZSJW+E1
LEnvzEIAO5Tg6GUgvUPasOWT+W9q+TthDk9bFfmsKnzNTD8s5N+W9IpzL2bLmnYW
12Xy5arpO6/XrxKsu09eiDwgDYAThj1/wACKnaXI22S8VJh1xXL0X98cx9NE5sEK
JuAjQs6tQAqRAZjN/SO2K0mm20y3FgZ+peGueL2ur0kDG8SgNs0aGiZHVZdu1EpO
OCeNshHij+NgxG76j5xW2xx/GzzSMpxhe4pjZA9CfioX+T06CYlBzbqao96hgRcX
NjRqosHD+Tac5FC04hgpRdBT3DH4IfCM6lrrHKsWYjx2hm7418b9skmDeDdLOEST
UPq3sDGmBO3YHIDf7cHUo9vY/0q4gY0eGcZ7AfxQphR5RgNjM+GEQ93prI8i3fLG
aka7KSKIVzZ+gK7BbDr2DYTegLtFMiFsUw1wJfc6HzYhosEtEoFXOtgKEyCwfvyT
HUYSx+VK6+ijtHBo114dDhiMHkghQec1NWHmnUz+W/CWxnjAywFoP8wFUiWQKhno
TolSR8LHf6a8BpOy5SVoOrtArWTCQdu3tlmXah5yE95otFiwKvsMgeqWAMpFYDF5
7N/9cPUKyxU6gLFDD10S+/aIHvt0e2B0x6uge7OOhoF0CmE6X663dPqCKM54/OAW
NwcPMzJEMbLJe82DRcQ9CxN8ZtanBNnzO9wpLaDMabkNCLAIJkNZnD5ByUdgtS9T
cTHsYjva55JF0hJfgHzeAcy+7XKP2e/v7qnN9n5dP5LyHYzsRJwJYFrPZDy7/l0m
DeSSg4Jp4FRzdQkUERfVOxgcD0j2CqGssFqCzGpgO6J7d8RPldfFYdOXhGmYymcz
FU/Q1AUrdJ3NzcjebJhlcB7T/Rq81wRJwPpOm1jha23pqB1ydKRNMp+U8gzxUXs+
xYCfvZkwaBgWPdu25ZSiNiIKxgDaWZCzheh5q+XyLneV4NJQx7XmhhSnqtVmHrzi
79Dc37PejfH+SeMF8PkQwFq/E0GotcMU6fNYR3vQO58bon7Rw1wbcdbkrbO7YI1P
eXEL4MQgcYTO1mhAnbw57MkU3k79JEOsOSv4b63LpbPPSWoQwR1lJsH+J79y1msd
LN9bSdOTHoatXmPpDz6+fN0UzxI8B0knaboVBVoi6rrQ8MCaKLxYMnN9gBKkh8Io
kLQYhuNLnDWQdYHewmHOJXvhZAI0OQ+rwsuKhNDAr7tg61YMyHLnY6N1+D4r+f1A
hlp3ejnvkOfbgrSpJa+Atgq+yZu4MXLKXYidAiLNXXQxdeh4pyIqIKvRjrHC4WEU
xxDIBGMJu7mfnnN956zJBqcGEnWfWfUGhEDmBlc2VoLihTxikep6U3sUG8Ttv0Yd
nW4k8+mgWBhcik9X3TgGfSjd4ByXNLxMXSnRGOuOvbJeHOQ7XYdfiMI2vdkERLLq
Ai6FLMC99c59Q7Vho1HHnRBpD/rHZMoy4J6bWqSIBtpEDCF3BfRYt8BnigYBz0iy
lne823ZN9OzvcbnJFuFcSxXYPAKIX4Vb5mAsSlueXkUAdYGtitiVzsQokBn1eJgK
PlcX9h/jErlT/mvZYc4/NNB/tdf+30O8WDsuawS+jZ3qUJvD4zsIcOgBjbLzrqKQ
HJQC9/7sdhKZ1W3DRXLpzorzAhJIDmYTiHNb4HyB9vwPfoeG4e2UkpJoftfwG1Av
snWwPCl6xmKhAg2mFGIJ6Y72yZOu626Qjig3zmrt1csb5CBDsK9/u/iBbO8WR17g
KVdC+F+IQ8Um6zShlvyZL90V9K+PRRHry83I3pG1nFkqXCRkljzTUHtyBGT39WjL
3doFKDhmElJ8n8k2XDlQmrW5UFyzFl6ZwP8vz5sHwDUPUgmXNmgFGGz5Vu5jlOsk
/0uzrkqvSoGBVu4aZTrEFWndJ8TG+1PQhVZCwDxWxWuV5uXce6ElwaExdgT8DOsK
6B0/tdWMbQg6BGk6N8YkAxhfv27hMLomDrKJ0o5IpC1GrhCE0gXS3QMnJW6xEcSg
HaP3uhrlKWTKX5l7cU3MogLWBfnjqP0SEKsnLE+8hcscR/g5Jv+KjsAR4SbnqLOq
ntqwofXVS0WUlCcwAy7iDoup7KnmUlHFo2kq08iW7XGbK0ZEH0VKA/mO1bQFQIpt
Y0iAtsoutmZJrLbC3h3y+Q8Em5ybBeq4SgxMgpQ8b2iV4VwljfUVEHXuFCjPZcO+
UwYr8tu/CRw4jo4vAXpqLHtQhO3rxB8aFjQv9J6hSu8WyYbNUDLs8bdHUkHSVFR5
CiwlztMXTN0Uf/psynLsQNqt1ZFPqB2YWblAmVQqk0bTYWLueYCsiZ5WXp0z7Psm
WUZtsfmH9fN+8i7ti0OMlgS+A+hluTNfJtQNhpTkqMiJg+oX3WHWCpxcYFlzNwyO
JDMpkbG+ntJNjVh+ASy9VlE/kZJoVz9Uv4nFT6fR2j/NUtEnhn2sUkreuNLUGPzv
2HjhLvl7rriwrVSAwJFlSkYaZYdhzDnEAjyrl0O2WMYvr76qKNF0q3jflok/ag6T
yq1a6sueuT68GE4uwpKTV3j0HwQs2royc4kxt4oCmlftrFe9qz0bKw2LZpYK0kjD
rnXPvh1O8wQy5PiJVJi5ljPBkG5Xh9YpEFKk2id06IPNGkdkZ/dTXGfQ1gTAUCQp
bdnIRdZZCto6sGnoP9lP+Sup2NFH8zDtcsz7n91Lw9pHn3JH2Kt9pGSitlBBtN/1
NayocbWlqiAcbxwd7q4iODH91FYW2GxX2Qt+mP/K8xvYrXebYWO2PpASn5PDOzHU
8g2rKBdh6ZCqtKMoHgXPf5XTuDn4HPB9crtP9fRFJQYZEuN7AIKIUoyACt7Hf656
2eWfHLlj9Nh/+uhlhtLh9cBl81DEujW80lo4yNj1u8tRfpJ6sCtFE7wqDF8DfGwH
L71IB3Igg6JXmzLJpKcyNEWarlXMLEH4DOSDypYtL4RhQa+IWiq641dsOrA9yhtM
t5Bsm5kwuSAUjnAoOrJNxXHcWcoWf28JYjVv/ZOIVWPdUXMKLnepK8nzeF7sSJcO
qjrJyk11tPBOxrNE/lsJnoESSn+6TMKG1cGaWR0SU1yCcuiN0G1gj5iaEmDVQYnR
PtcYV88pngleRrhoJ33m9hoRsjsVokV+kGx4Nr9+iolBksoZMcCeKtQkHzdfNSnL
h+NdllurAvjmPj1CWT3fndSXAhHhxv752gtheuLLGw38tXMc6ayVBQ0HTkOXIaul
uxNP2WKAGmfaUO1LcqUQwFW9p8EN0NsKZRKdAk0NgddFv8cHsDgDBfSwGA804a5U
4QYrdgNfMaw9YsdWycncy8JgDorlpsG2szDALVF1S4UMloHGDkmdi38uG9OJOFbJ
XTjpImR6oKH5EnfoFpiXYB+pYiYdKsq536sFYCrJ8ECeADU/uRUaI5ZMyPOImMgU
dXFisGuQacKp8fvLZsHeg17aon6cWXBfotPitDTIwBTaDGCjueeINdiOGzYhPsFI
DVM4ZICq50p8Lv2oDbUl1gossnOsTvDClvezhp/u99Ck3TreU3BYG169icNL/kS1
kQI1eaeVtUdMpD4u/NG8gJnWhIvvLqZjSHroV6INchYjzXPGTbioxX77M2WoaL09
Px+pHqDw9MqKF4jtpZmli89mobWIr18TWVmDC+gG7dbC5Jm0C++6d+eqD6yeTjZW
4e6Q4ix7d19tAMfbvlmmKVuSy8wfDNRHgnOaQnh5bwE57lCHLCbl9G0XkDsrGy5x
U2Qur1fOHK+9bVtXZ7H+Hvig7CRQmDwEeL64zhz49HnmuNx39KugEdQz0ARQRYbW
zdHLVF1TQ2mIuEfeJP2wqFqPfXKmr+0azTliPD1YApTiwrjPaFYFUmNYxUb+Rl5O
yamNthvzF4h0YcREGdQ1dL1SmlqgK3gv1nttcjvpXPwdtPC1xI/gCGSH9UVYNGfT
jVshiLD05fjskpEBp44l+GLOFaAd8XJnqze4obh6HTZv1ZPpusErQgCrNDGKoTar
ZLJNckIi31LUK4afflp2ySGiwMFYjr9MFzKyllFhieJ0F+1DrPmY3zYaeiO+ZKQ8
k1rEkPKkXrXDfofy65/0t6Dbq8jp5UiaQuQaeqogIhBoIkaUdMGCgmC25C4UTmzy
vmPKDHzvFcUHR8Xa2BUbMJ8XHwvtfNcxu7LGdrZk+PePCd9xkpjcDDRRiXbg9Y7z
l6m2sQ5Tk1hTU56hRfABMkswJ6Yyv+ea3F4RqBdW8oYtG4dasH46Rc8FkkYh+xZb
icOrxnbq1n6zISp9ilDHCsTEycII4ghK+I/WwX9XY91ZKJHjw3RvyeuchaMOjczT
dgaKmPkEqyiYZw2Ic2FIflySwJlrfxXiYgI0TY9HprdeuTtFRqF+UqOMtiKcP3LP
eONi6/wSOKn8/ieBQndSotIJMXZ9KhcAElWOemsaJBehP8tQTcwubFRf7iL++qef
3/MSuW4HofuLRF6J/+pr5tU73rfvNhChbiWboZBiX5OZr++taSKZCBCsI1b6BHah
oOHTyftAm7PA8XE9+Iq5rrWzv5WNeUA8UgXRVqqufVNldce8u5EhY2YglJTrBwDw
sKXqbqM0aj39DHfw4HNicUKuczdgOLsBF6gbSAngP31kIP6iuo6FeDuR+SZYSJHz
MMVL6O38TVOkg7g8ItRVZb8DX6Z+gs7hzKC+2wCxw87ITqfD58emP2y+fgJpPazi
MxhpaORXNv736HMUW7d9RXPLAs8o1Z7saemOwXA0kVnHNuKlZzzX54U+LMaQh/Vp
ZG2tzVQOZf0wbombRAFXAprARKvWrJrH5QLzt7INZLO3UOqNy3/sek+lSb8O/hs7
O13Oup/fLFqOuLQ4234wqQcHt+C149Kt8fK89bsZLXm++ZaWlO0/eZQGSI7WSdxS
YhJh84Zbe4Q26pZCQtuYyWcfDgpKxvqz9TT32wiGmKwqoGIq93TtELYq+udGAvSp
VGiUBMq+lp17NOYrKtT0W6b3z5H476L7sOsDmj6XArztsR1sjGtYhmDX0J7NGq9T
FYFy0nVrxrIP51E0KJyZIgvRkfqWJDtnNj93if5myXBdAUQKUBSUmyegec9AHHUQ
bKKHfB6PgUhXJXMft+YOEnjwsPoVTXtQB2FBjJskPh1roZfUb0KcjTIrRK1J6MFI
Jsph8ISR+KyLVKN7LWjnWV9tMQZjLiEkPFJ4iszgL+paKYB4IfR5/+r3FvSSI8fF
s+0AMKrK7r76aU4LCTo8EkaDV9khs5DCvXjdOGdV58wWHUyvy8dergTi6x8R62SP
UtEwkVNPC0XrYHJtnaM/hNuyv/xcX/4s2tCjlu5WFk1Wf+ZY6TEUQesBJjeTm4fQ
cyaLZFRoWw1yRehWUplgjeck5Fb3yBKV/nydl91nvyPO+HWQHkMDwMyHt+F601q2
eYBZ50xXFxeJNcNMcJfCQ7zFrVDOnjnrgKAf9tEVgNFpt2ZIcQ9Trl0B92eUpqo0
OvZ4f8/Urq1hvV5+9b4/IoXVgq4Yhg3gWLEDsgQzsDyiGFHNXZe/S/k1AHGzi0B0
VKyIZjzScjUUmTL+SVb3VsEyF3++GQQJKCJlVo0JRWIR8ux84Cmx0MgEmkdPYpZv
U7Zpi4engomGULeNHncqJ6FhabKflHhRMg2yN0MgUgIhxGHu7A9iwqcOaFoVYtP3
xHrfKzu9ZUGrlaZ1/aZg435vEdXoiS4B0rU0rzwK3WpB9dMUfi+d78kx/Yi2A+Bl
sCrke6u96bAFiMUSg0nRb3yWCmjHsh60xesQZj+5NnrgfpW9vvRXvevOgiNUgYDO
H9ziG4eo8LW7oMim5+oPIYfSU6Qpm+g4NELmSF89ZMZKkbukbZGw2y7uFKCJ77qm
WU9YoItRW4MBpaD5KuqGPHoSk9uMafDZerlwsh6TziU7Fzy07I9K2p93WAe9H9hR
Cwtxq1a/pYV6vtDq6MOFGmTYd1qevAXoe2fzOf8uhNlVnFSucwnp9mPrZy40qYCD
cXNxPX7fkGeO354EJ5MTD3goChm+aYubODI4GZc9I66vE5Dab2lhkBsMgQ3eWBiM
DyEAfF77TI3WNt6wzHCs83O17Yxdv+Eilz8wQ7Tp5B7N6YZ26epgQ1PkOg/gqB7n
Vlr0uOi4OVGYT6Ts/fwsauKBzfIzpaqidqW0bpxdoJIuyKraSsKcwIfQvXaj03+N
3Ai26f3LJ51myWeaT5zENf3oYajG14ms4MEN6aSEAdegXLJp/HjQIInG8tauC6hf
0cUSSmhV/zHzqfqPrnSTHycQiezIRcNtcPJJoGuQDmTOFLy+LhpxC6kJNvdvg0mi
NwuqhJ5zea/Qxg/jxvhU5TAYJIAcg8PvndrxHQZmdpypetvQFLYk2mG/LICRtYh3
zrAkb/PpJKvNy71rxcRTaPfE3w/2OGam31RmmU3kZ/6clxIfxUleng4wwKmEN0s8
U5xVwLAXswjJ3d1OvnmOlE04+GzfvajDV/jeuhi3QeJfJ7JIieOV2SfZ9G/2/v5Z
HK5Fd0gNTqLvNIrqVcBXZGMV15iOUS2hYvARZFdxhCAx9CSSfXWszKODkAY27yD1
WGSP9BmQGOaQZG5gERhybvZ7+cGN1UN/qY4DxK9zEYjWH599BuJX0z/4Q+axMTfT
IWLzhptOzP5JlRB09ZF+i1t7sPtBoYk8KgM+bYzimRU+3WFIQRnv8p6vdf0LEpGb
IMmWy9hV9L9ml9O9ZyYJkw4kZFKEDtwGuIkzQfC6nOR4fQpYQQbL95sN5DgwwlNQ
R6OLwJ4GkHkUkmI6LTXx53FtIuGEdeTWBub2nZvqzyWUBGiuKzJ1V5EOwZ6ofiVb
lyklPbAUYwDwIiS/PXqcdQGJu161soPHFtB5bqMrztk500Nj8ySmPNDOSp5JbAgz
5cA4wFdilF2VkcScFka8eGc/pWYRhmSskmOgOmrjeEowFJoN17zsFXfvN1oSM4+4
vB1o/JVv3D9c5Ezsxcihn++JBNZuwSoLX01it6QqIUCXvysqK2SijB0ngG5+jm1N
ijYzhNv+kBSos0+svq1O7dGjUQcH3/3Ph/L3WdRu9YfDlcpHycimdHH+Bf+LwAhW
A7QnuQylBHIeh1ISRIIl8P1FYZOMYwZCm1F4WSLCK+RXLqJYrl9RC4TnEgpe6Q98
WQum6zgxKUBbnRdarnl8RnH3yNfOue2NF0+BGLK6IJ5gW/ipQCezvc9wJtI9yHXo
HlzaNa4C1QxNDUE86k7NO0v2njFfDRsp47HiCeF28vgM6cshThcBet85DG8uPt8G
fbnB3wMva4K3DokPGSBv68VzBoHE0ZwRaPyIddzhzIdJG340M3VloWBwPWNGBjV7
DO7ldP2ZTgu6uZB1lTFcVMkOQnJbDAPjRvMBnYAbxmEdUxknADs5e0gfjAUOmEG0
ZrKOiu6S6KimH0E6piA5xbHmSXFuZpqw2KMIXQqkzW3k2Jo/QI9xVVL5J9DjkFof
6zuVZsCSn2L6cTzmO76f0cXRk4Nx750QkZVpmM8YFdO+5V6srrGJIYdXnEivu9c0
aVwAnJt6jBtPZUwb2XREFvfS9wgonhGc8DKzoPWeB/QH48taDr97og55Wsvbt3w8
DDw5j4iZmiFWd0hFJP9Pp4KGgtdRUqv8K0QzX63LgSJUrhgI2ZwFJbmFBDMWLjro
EsAGLjUhVw/hFcykcbwHXr7XnaFkfENbICcv9ExLX/zAD/zx9BIZRzc+RThRffi/
Xx4UP7aIN7fhsSQs5OFpsLPSaW38T13sK1gnjlyNkQ9a5f8Vb+EENAbKyWh3rPnu
pbxR7up3EYyoOjpNTaGitB+kGKzEmVZIlML18/XlwXnqnyFU0qi3PX0QPdl82Cxg
8e6gJrg2Rgamb+2mQSzMQJ8j0j5Nn2wFNC3Zkh8ljNv0Wjf64JzlapceecpSqbYu
O5DfTBOSbKQ3H8wBbPLHWzO9A/afcc15B23SKOIcgEDm8FMdJZt70r3ANpYdUdps
ThZRkH+lNTKJexA0jttX2TYhYqxaI/SxAM6opFq0WUqFHdh03MVIb1H8TkvjGqZZ
iSn/YFT8sKfr7tn/Nc69O4iqsy8wH1CZr2YbQVR588nO5+4tPHKTUe1EEAR7HK+q
Z022mD/vnKvm0QNTfJg6MwJH+C+KmeT/OwDCAbFl7Y7moErRXEX/7+HhFXlyN50T
nZIE6znY1APKYbFWF6HPi09lRs0TgDVmDu2bFnJW/tkAaecubrcQwU3qDnYVwQ2G
SC/ey0mQJiVyOd0W8p2N5iLqeL6ZwtCeYe6/UENj24bojgeOErAcGu7dNAoKnUnT
aku2N+GFZGaBbPDuG4bzbm2fwTSP+O/f9qMS0zzQGNHD/MapDKEOnNaMbuJG55jQ
LEJlapjmJUECfJ/DyfhkbieqMXc5NdP9zomUpWthmS6R6btdZ0A22QW0/d7d4272
iufvEL6gB0PXK54f2wI6z480ExeZDfqDqRbl0pXUXcAkd4UfFFoqYrsqye2ljbyM
lhi8gPiSm0DZx4cyV9ifCNECvffSNyi3md02t/2RqcIUivtkXOpM7rsU2iUBLdW+
9FtaWx5AHPptjDiqX5HltDzCdqXtGLnJl2oZm+RTCW8mT+hvCN5fJpOTnn9Vktzk
6X6/nEuWT0QEfa5frUPImfJSSOAIouM531ZqHVad2MmHCuaazkJKvCjQ4BoMmYnf
itIMPxS4EydiPZvfee5favZlAILLpBX8c6YYOniSvhJearsChNVVSJLXv2a83B4F
r07TG2NE/syEH1+YwbBRtNPBm0uQnt8Jd5zGSdAT3BBvyr4h9GbpNXE/A4ULh36A
LC/QoxKgG4JZztuodyL9szGBvkj+br/CQDS3giGcwRMwey5k23SyhU3RnyevOln6
29+EbtvyJfSUVoHtm5v6TDP3J93IRnyIn28JfUYM6Cv5VYPmwOy0NrSY4IDFn5wZ
CeZuALQWelK8h2h1xBQ3vxEpCBXtwQZR27KXzDR06DeMqqzZ8noOWrh2Fd9JSulI
037Xono0798j4g5vBDIP5Nn55LtGRdmZerkef8QhrhQiFQP1YCmaWTNpfRQNOwdi
LJ7Q3Ecxr3iOzy9VWh7fM4NBKMfZzldkN9mnVmdZdlo/0fsxm/jU0ypupF8aiHIf
V2B3Em8184kjBeoqDM4uYPlYHwYbdWw8YKvOBEm2/m7eyicJzZcdOnX9oAAOObKr
XqjFMVgfXUJlMdjdqmVwqaSlt2MF8jlH1uiMYRbF4niSnKDEZzbdGQoWz0QGC3HO
UQvkHKrD8cqc/t8z3nCkUov5uSNMLTNVZ+4yfyU+B813MLe3xZagf4zeOhR+IBGI
Y3QpOc27rMfHWoaJUfxiCkatxiI+ZIbB8qZvnevjHE1P74MdIciNo6U5XfYJqpuQ
XcJ3coMcod84j6pyqpVm9OM8N/h5q92Z9/tJNVaaiD0YIg6eggEnnwiAgc+S8Bbw
44oUDTesVy+ZNKmuiziagdFnU3LFZ7G9Ckd+5QYxhBYYzKKFFw36b88FvqorYvj7
kmGRoZ7MFKXiCK6b5NpTgJU4zPvSzHPTgE7a2gfJ+2YFNo5MRKbq5XQ0l4O335H6
gYUn+k3OiIIVw6Guhekg0b5RXuw9vqTkiUXkfZ1V2TmpS8Wht7frQlbffWxDtVDx
o/cOIW1zcTMIhgWCqzcOKMCTjyb8CfuZhSG9lrIaGkowwvcRkMxQHs4R3zx9aPDf
HtNRh6OMNTPE++7+rsuXdjZXwb9Kn1k39YmLf0yNSG1tfSq8HSxqD5UNmKSG6e1K
gDAOk3CqgWXjsKVjnQRFEpvd/zdtqPkBiLPuBbKyQAWb+OmtULTfy5rswv4siUoi
YsmGqIgJhK6LvpVSyCpJaWFPHdtZ4fVJbpwW0tvlLiJz+Q1NzEYdiogKVldSxW6V
8lj2AgPOT5iJ3luRKDB7Qd74ID3w6c6BBhsr3hPHPOHJtF8IoKYW735L7OqSkPVV
7UvrmBd7cLJ2cRDf7snWrMqbXV67D2+WcTufRGrirucZj3sj5D8vS8mps3aR2msJ
HHCkbCJWtcZLvGuET6xybdL3YLYdwV12gVoEoThxf/4HbkfgcmruWeJputy4kkzO
I7Hq/CUAadM2yy7Qx2IjG6p87BW/9YAFajWXvP0ow6ki8XCHSgYdSu0/wFuJMyMg
J7CtN1ERJW7cX9ptPVWg27Ra5CciF6xZ3sZ9Z5Z3CB7+4GBYE48PjuFi5cCJFpuu
rTiITFSVTOLAdanyb3psrPrw7UdK44JiAwlHiJf+rkf6agjAmENb7Q8km2anCq5u
i1r3Cq47Mtdvg4usaU6Cf0evsZte+MmD5OnA71dbGlf1BS+XpvVO4Xi4uEELglPv
0q+M9PeqztlcSWYCJXmcr/h3EsIPmVpszueiGPRLGSIkvdJmMjkiY1bUMVq3Uoxq
nXGNCsypOYvZPcgKNv7R72Tc8qG51wiRHl7Lu82drlZMITX0cC8jIN8xRYAEv4al
emhFNYuJzQtNv9XcPnyxA8FM8eVbgEwZreUQhIJ5FSHRvDOpp2XYiIURPPz5Dssd
dAxfcTAweOWVkMIijlWz44PLAsxQXgjJDpUID6/R80OZSrnVbLHFX8kmpJd7mL7e
fkos3OTWMS74O7+tYP3kjoOfxnPyk7dfq65MbwbMC62myGSfPdvTQSfoN2XMhecb
/66A+ZW4/w920ZcgAXWKn9KkcfIYjZnR0HQXqWwNhHr6rdZDxmMkNtZgtTF8+Thg
55/cmofA/9rLUO5EWh7paEOsrTW/uWnzr5mjrqmA07iNEzAJZxlSQdP+AlUvMyqC
pI3vSaenXpORUdlc7fSMKbVceoXh5CVj5rD/SHgOv9i5HA2t2acVsON77LnQPzBg
/WRophLQyPm6MRDOz0FwcVFX+YfRSFnA0iZk6o85o6Tv1fE42ByuKjWrgyObfPrM
Lwb4ignv7Io3KqCwRYQopa/YL+qfkbu986+DlQNJTZnsQSCCdRHGeVkpe7LYoax/
QprwsmIPpV9TBVJDQXExFG//MyCblWfnNBO+32K2iR/lO/GByRtzbGtqtWNcNxlt
4enc/z9LJYv44dVx6huW7NIJbBHmc7tef50bw++w0+66166zoQQcNGICBAIcU7yw
H3EWiRTgKeaRSf/NQtXrkTeNisnTfyV81iddwGAkt5vgr0AIEqYNzRDmXmOEGcMc
YpD8dpOcDQfGU8FsBdR5o1XX4xcvgaXB0Yzub1TfAaxKJm0W1vq0XPqcD3zSvQ1B
d4o7yOlYPhGQjIA6yMPGRwFD34RstzbZyvxyirE3Y2oRiC86+WErPtvxsNa5aPY8
di5DiPQX06LOCyh+Z75o/lmRhztbeCGVMHPKf1R+2Tb2yzvUHXF+sUkbjBGBd7WK
5MUd9394s/5m3ddOBHyVlmX91NTBlX8G0ldQH0WviaE3Fb5JZ6XxhaZdsHYDRNpg
mQTbnf9Ukcim3NosgMgBlXMIPRurgozWtODJ2RpUimFPVbAsHO/SnpvCX2x2s9BP
Bb29tJL/zJjudfW4aV3UJelENNcg253SZ1jLvdmKNtuZ3n1h/gvA7YYX2gHbtxHT
L4Q1b3NWOK4TW/HGbzH3finyq/BYf+8P4xR/Zb73+/b4SkpSDdCf0NrwxERsrvWL
YvjemznHddc2z+HObotp8lxV4fRgVjqFIEt206tLkuDQg24EDRvfucV8DgrZ2eyN
NOKNUf1Say+gOybFZ5g6DcACH/kkZfweffu+QhH4M2gknso8YHWhgG5qtAYh8t/Y
+0UqW/QOnv4csyHB5bP84mZ4sV+NuSt5NIW4byc5sP8H0RxZ8QghW9ceFXvzh4wD
BYEl+0fReL8n8G+h3wTfA1HVjqVCCGptQ6wrmdMkEVcB54aNWYHFKvjvoXTjeMKH
OTorZdwvaQZAdxZ6PuvrxNjxVrEX8VGIkNYJ1VINtrwgMLhPSOCfOJgx4VjFFTyo
uIBPrXgdxakjitl0p63rEa/O4fqzFWEcr2cqEYElP8EgLMWXfSuj1qSrhtlIBYs5
30giXL0Jp0TXcHogXWNzCg1ThsfQ/1hYulkCVn/JVCu1VXI6ospffYZAsHb+pE+w
7VLCoKBoQ7OIz8SG/9O8rGzdunTREOO5BGHf6wPBzDrKJ4ApsSsCZuRkRgUqypwU
JUGpvin3gLCZA0Wg5Hp2s+Zx4wMZcLOjnQvKcEEIbL72L22Jv09G6QZhoBgH+13x
X8NfQcC4ZZNAaK4EMrHu2LYOae9u3z/X+oMOGUirackak0TvYgVuSRGQ2FWskZWi
HG/GLEtT8VMdI986Q2rfGtTLftYnGvdLAfSPmhl8IoY8Q8kWcp3ExH6dMHJzj+7b
VrP8zL6U/Zlc9Da9dEe5I8fe1HEGixU13KFzFsvdXhxt8VTbOS+E7tc/Naj+lrKX
eT/jKrC2c1CoS/MkuEXTOWfPBepAjTKeBLtpfFB0ObTf2LBIQohjrdJXBN8HNHsu
Mp4LYfmNxpYABT5JOth9/aMAmrE/1fPwa5czTpXgdJipEPNf1oeoxBnsInJpwpOP
T6v9x2zGARwbenVSVZTE9fCTsam3A4N/fFs1t0ietjkByO3cW2mTCySa24Z6Sdrl
VDgqR5ERN31hnJB1Qh16fjFpH3UBOrnkw5EfIr3g1BuTtS1sPCdCHIohSENH2rRw
NR4X8T9BYGgjL5C7Cp/gx401eL0RhbXDrXEc9G6kTyKNZWz4opQeZPdU8OTAYuQ4
hDCL7enSdto5+/uoVu2Hpd3h+cHmGVLperqi0WWqYroKi8bQJA5MmhgSN5u8+Ys8
LpOGVqHQt7PzEOqtRUrfmZ5gTtXF5gFRKx5hzbRFDPC3NO60BNSWIeUxwIsIGq6C
CdRvC4pYSMlPeaunUkzW7d1yDBtmjhR8L2fHp3ycHvAbESBxstgDACO41YFYlEDk
lP3Wh3zeFsFkPsUxFOCop8bqYsGR8iPvf/+F0GqzYSN9jaAQI1h1cgVu31ZrhPCK
NV1GRHBPv4EzaWoySSYKy+rfUpIwW1d/LndoCvQ4T1/5XMTa90+H+6lrrEKhVYaN
Um+ubpcvIeFWf5irpI9XZ4qTe9qfuvDmIiulerEo40SATMrECCMIWbrYkaMeqe1P
W/CEIBKUF7dbQh7cOw/wJxl1Ia8BVyJ6l3TE6F8mA0FJ5SCZ5LJrpS2pwVl3kkyo
i2hDsylJTih4zYCjcoof+JQSMt6YJhIySzeRni5aXT/YoZMxECUY1lTZwutZgkTs
FfB74+Fl9dgoHmXz6ULkh6SiIpkRdDm8YZ9pqvbMJ0wUHJfDgXZ5DDpzlUD92pMo
4/hbi9LlQ7M6tWL90j1KGfviHz8SKEZoKECyFcfPn9l05EIan6zoA8Dixdqk/Xmb
4IJ/CG/Hyl+jsQvE9hE8DwzjrMPUNB1op8URuynTbSqj9uAF3TJryzxyNWHMR2wE
p/Klk10JpUdHlngjGTNILr046zmkqElfcOC6QyDyfDzQQ3hKdtoQfQnALnpgm/1f
UooYUaT7EuIPVfX8iLnn1tm8FL8Urh2C6BpJy/lUNMy8WwoLNwdJxW+dufM9rf6o
+vmw3j23mZgGlpsvBahLZL/vebkCY4gXuoVc55o4PsPwAL0xMI5Wh+CVEcWTMAjm
6XNpqFd+YhgiM8t9eANCMgeqADvXG8ZjH1iCRPmhrKeTZAGS+kXw0/PCzGkPKm+3
7qJZRSaR0mimZLPwSlPRBWLxb1N0elDQMcN10p7dvUUKWQCu3Vcy2h8X+lcRiODW
Svd6GpbmCyoNVvL3n/+issxk8IXgnYq3G2M5gixaUGmYel+Sa3IRELfW904CxWSu
TMO2ri5nS0P/XiSbT9dwd37eNt6GVOPpx2HzV+rPx+lR29B/2UgWMAY8PlKu7mXm
+E18VIqP9LxCKkTdUBWL90Pgs0ZM91j7AtwLOrxs+6tD28c8TOs12yYRDT7oSHFw
c9fp9uPxT+kB3H7vwnyvDGH28y1ZJaqwQy0t53a6rlCvdIE0YrpZW2FpT2/XPl9T
tpcvU3OHJnwy4PN1SdZmdWMaxeW/NzsyoGfQPRIL8OlVfNUROkH2+F0zaaa7RzBj
v6kgqlS3FeGU/i2KzOBGe/5UzYs3Z97urfDRc9PyF34qu9tvmR0kzLenZQiLIuxi
KtZmUxVDWJJYyq1axL1pKZLj1Bp12Fb6Y6NY6rMUMRBa4DQ8lh1FHyyt8YIemlwK
azwxwy3kocUTcUfDAhHx6GKNGDhlIcQE6x8YsS/+Fyyt/GbCxxw/y31lJXSdubYk
R0uhI2GD21ouZVSkLY2ZEMkMsqjy0TAzwZtBXp+x3DKWmUSJNc3qIAKkUWbt2tRc
QRMYDQcIL/DZecM86JghosUP06/O5/jyNA6MvJVvdN0ft+RPe/TXf0faAuWIXQ7a
eY198bJBoYSPuo6vJNo0ufb0nWqppu6gVtzafk+gvjH6/6/1gG6pDlW4wIH2un3c
KRsMz4XEWPTBc7l0+p+Rwq7GAefcErUZ9yof67DGuIm7dc0+Q5nnOby5Rmisx6fs
jV8+7Y4cDF1pE4pAZ6DyB57PGf7JIHrhax23gtoE72W/PHG7nTTpzz/MII86Jt1r
uvxdIQsAem5o2OIeIn/k68by5dBj5VdoqQKaA7jaAGUt2PLZ0+fKa+8nZ75brPHo
nfpg37Es3OJeEmqZCd0+q4fjxP16p/wbdlZqh+4I1gI38vH4Hf6oVAXN4RYFd4al
+n1N77xXzjyXYu2EyEwReijOmxFtDHzwi3TW0Y0IcuB1YuMC/+LuAFECZ8cfQc4G
tqaLgKRzPOAWst8wn3GtkoZFXZI7ysF2RsFNn+W4fILm5dpPE1eNnqIbo2seOypM
PAW3fdUFqE1KrcvlpA9cauR2ZEyR9tUmjjaBzwhlF99/3NJUlyzsIActDlYukvmB
GCHbNqsYt1JEGKVtT2/Bizr5CIVwsb0wsOP9z8dUA1w0BTYlHLdEy7yhZrv0SIsF
wgVTHXod8nUvCjD0yMzvzsvCczEdLa4q8eqKQKSUTE6as4gmhdJYfpde23l9Ch7X
9TIxyFmQzo2OQ/Z5lhr5CDnLGQLEDKt6iTheepv0VM5VoDJdvd13v8QUT3qioEJ1
eweFAZZ0OGScV6EJ/uGLtvEXAnwaTGMGM3b5XconoRCtPindgAyLhddsmUYUyl+7
9OZW1z85uDTqpHGG1lN8lGqTLjAulVzAqVgZIchL7+tWMOJqE2e0tbIsDSsHjn4r
FpnNiZfrNdG7lz0oRo7ZTC6OEucwENBKWCU5+eQ+ILrCigfufsjanjdfgYabKxTI
2z2CRMY16ZLIGstlp8otzu604BCRbXb03iRo/ShzBsFHccmPD53RSVZcw5Mix9Pv
0AncNoUN2wcNS0P1cO1Untocsj6ZIBZqO2cKwsSW+2TBKs+2qNY4/oaPv3Q626wT
OFdclkkEmpOrzgT6HM1Kyk6aDXAUDfNW+LeUlP0DtH/aJ0sB3rzKFAvo2UeXzX2G
46/j+wGiG+hpDCH7GgLki2DJe83eBSAKiS+z/rbxuOeT5BhDO3TiU7Cs0ObEP5rJ
PN64ejnHlG5dMQYO7sLg0hCfQs3IA5/rlX/OlVzyMVcSRkyyZLNVUKkt6R4miE7D
soYYkmmcIna4/Aot03aM/DnP7XSW5v+FMWTPEK0Al4RZrx7/bjGoUh1WISi1pOBi
se3bBCNgUuAoYKR6w7tltieWBVQHFXRK9Ljmkg+IpWkweuy4+1rqyoNGaTYzFaYQ
cfM5w9k8B921za+P9R57wbsYPadMF38KsiYESIFb2mevkAR6lWlr5unYY3Am1viO
pQQAlTmGsYg/Dq8mUcljYSkpNd8I84pjnxrTs+dB0VFHfeK6kf61ASTuUZmwk03I
TlGBZASCM0f5AC6Ke3PllZxifXjAeC96BK62t55AoFkxWuYRmcUX1pGoV7P/Ytj2
5wWVMaxniVRoEqTIUzDfpCdQWbjR5dKnwRpy6wHKLMXSzc64OErZQcNRnDvCsYY/
7HVUIgECEtQRTeTIlSD5wMxKAKMOdCnzuTddrb1H95NpCWvFM+VjGWRDYVWSoEJQ
mtCRdzf3PIkNOj843UA3VUM+lv3uRBD3OZrk8DFiZTYAh4awa28829ueHmYyYt+H
nVvc436X3lNQKcd39lsE1Au36y9AUdwUnRLg3vTHRVqA60RjqrONz3Gwa5soMn4V
TIyoPzp7+XPKiPn/RborW7OVckc9Cr7uC95iFDJsIF3Ka6SUk8V6rGPXctWiww3M
5me/PJncPG/5mYFM6wnc0s1uUFyVCH1WjT/0hYT/vp50No8GTGGA+2zdBKDTEofD
VNcrs31kW591QobEB9VOrYlLWqskeIPOODA6r7tFMzXcM3zTww3JjaLQGn4ZDHiH
AOKjRs2zHAPKhmopj/qyph19KZfutRRrl7TVBeXWMwNiZhjqg/CKwkHowDvwJNBB
cHjVCoSCDnQMQnuzsNAWBWFE950p2NCAH2yxsdkr7lWQOe+b5LmeGq2iUioZ5jTL
FPdlaZJGW1IRdyYnmNkWCbb91sAAtfbIb860SK1UUFrvVF6jNukwm4hpDZPzTLw4
LqO9kato+/7URUBvU0Jv7fWIn11+ALJphXRa92XLgnOBNaYCIzKIqsVT+QNjijlU
irb7iXT7Y430ftrvhAOnCc0qLzikbgzUYkYmGs1tqTZ4akqmkMmoBDq33ZFHNtcp
kH7xZVuNRJ4TxiHSyc0B2qxU5OWgCqiPxONtcVJfT17mnKtGwi1qOg0rmQIh5E/J
EkMPhjue/zOLmUgvRSjjhx34WL3elkeYnkMthd3kQKZkssCYFxgBAyj4pSxW/z8+
gz4hO9yniplxJe9Xeq8iNQIusuO8LHEVkdORtEQQ2uSIZngbMAMtFM6CG1fhQFWb
yObD8doKkfE49IJq8S8oIDsq+pihPTCS/gca+1ZCpBaX8s+BYmTQ1L1t7KCXa8ir
dugRaaTLUnR1p+EZlPLK5+IlAclPPkCK+pLCt/SK6MRya6Pqn1fZ8s8o6KiPpYPe
+yW86EwaEXYj8+Jsixs5REefC1I0zZNm5NXNUKSO9kcRT9Isj/C8KesudO6bQ99A
Br7zHjMMAQTX1XmGjwnnDYfrWQUh/FXpfGZtdoGEfo7+a4woYC3uQf0NlhS/i+tc
qDGgbzJ21alrBT/xd8Wd4RteZvhLuhQH14UwKu1gFsEgNEjGxvbAK6cgBNne9AiN
vTcCSCjlLkIR1rPjNpS9EFU37L5Af355ybwxj9B3yJubOgEI2lEcf9v0RyO+xVdT
XFJc6Nx9LzFi7hMSgyWnfHVjbccJTAJnlziQNSZ3NMItg6dnQnZBLvw2BJLrJaN6
FleeYb5muOFTxJV3ruO/1nmLzWAdZ9gqeBklwAcbkWD/1EXvfJIcJllFgZN+f3ef
5adWRG3H06lMb+jhUxcbSvt4rbvwhGB5iZMHIgDowNqwMmSgkEaKLWxqc9vFxMZW
wPKidMbEteog5SSpTVeca+JQe/HYSnyKNKt7EJBWWBn5hSMqbuFfwDj0GbxqSxul
r50EMIicpA/AndNBCk2qi0YtlPoO1hcHRM8lKoixkqPQtxZWl/ThPO44OpaK0763
I9J8w9wi1l7ljTVwNQMoCbpwNal2kKV/+NHVoe32Ped4rjh77Tg24fUnJMIAuiGx
GvIK+d/3QIJt7+TcGxZVBTM11eNyTxd63p5AgxhEgdhWIMSykBk7bQsiVhYVzbzG
xxEQ2Gmzy+gX7pNsYbv+WII8+RKpDOIag+FMm1Y0QsJ1pfh2DibW4Z6+FD+mcKsP
L8v4gKgNDFsjyQ2iWk3Uc2kljAqK1cgdJk8XdklfvlnnpwbBcLvy6u5xN1Hw2IV/
wyKY1XnwwWLU4t+Eqid4GibdCytXaWNNiQKOZ/BXSbhQL3q90hqT2ky6irYKYJP3
AvJrsPkmpL9ywJel7yniz0oAWQUVQO77a2RTzCgWg3k4pPSpjwP6JZYDKQM+ohdU
McUSk4HMXhfKaS0gNoj78R8N4rQEMsBoLWOkzb6vMh8+xtHniplZqEz3BIZBf8o6
7qEhTTZfJXTqeeJfqu5eM6ohgP/tyxmYSKC+S3ItbVRwtaFp0m/34Pyo4oZK5IXn
DsNCLVyH5rs8jRUaT4YqPxk9BBqenf6361bW1y8kugca0k/YkHFDtaZg1ZHaUBRF
hY521hLRgLqdDOmeG7E+Tn4DzFqitBczn7CgXtEwdaQssbGahrYauxuNjr3mv17G
+wxay/96SuyPCmUm6PrdDEjn6sMxsCddOi+rn8wu584XKWBMElLC8aLC9/LXmQVT
PRpd7fBxdtRcTR4FB5iy08doraIrWPqvy8PPxjSMIgVJYNjVLD/Z+foEU1pBfc0u
ILalN0+t5rFDuW0jFa7fXRHSCSEQXfSxqd9oI2sapJzvxnB4nKp0O7uqRp0D5WTw
BDOGRszK7F1IF2TkZze4yahLS4VffYNQHlkZQsBzWSTVbwZVfj5204FBE/liX2dM
QapUphJoXrciVKQJZnXB3SJp6BOBqIEDQop7blbLPIIwrHpB3g80iS/4WTyFJNFq
SchgeT75ZlC2mphVdjU5R7bUUmjhA3iKkoMej0djeqycZdahB/t6U3jkh2YgJ1Lu
NxKbBNqrv7uw2j8td+qS1jDGTszdBlyuSqIFABbOqp/6G+80ymHR5ZgEsb/zmjyN
JMboPw3O+PaMlI1hSlIQtUJyAFbqDcik5aahirS2Rd/ZWmNuenNX4GkCpCrWQw4J
zXMkS+fVAbj909bWbnzaP928F7C6hL9ShqM4WirX8RWoWO617J9Heox1Gc4XqXuS
3sU3qPaAwxVdre3K7aPnfhqwCBjZxensaK+L/DM0W0d9lLNWBJqwHnG/gda+muSC
kCk5yOdJtSG2O6NHNB087ToNKapQ2hAATU01MXjq9IbzKXQ31vaVdOx26Als1eim
EhFLRDHf2eP57/FpbTqzwI0O0INYyV3Dwi8MJwLhVYYmtQFWr1cJQCHevVCran0t
T8UFgdCQxiq1wV95tf13+Tg4OGbCSDTsQu2DwJF1wSC9pxqutCT2aI7CjjgmDN8m
l9Q6r67R1Ii6Y8PEg11t4kZi5B7iQPKN2n41oPDc5EZg/yM7QA5e2rpzZNZRfaib
vPYl1DwXSWIW2dSlwudzZ6sO8Ip3qpXs15jf9VyxjDinM+knTwDl7yIO5GDdbuVg
r9Vi1tXVDdEjG4bHTmWDTrvEuthYaTQpfMHKslpx56eVyjdHUhHRxHTnKk88YnTk
1Nts2EWGVMFxrn9iCImSt969S5B58twIKdh00iBjrMRlTNoEM2A4ln0LASRYm8J2
NzP/ABtTS43alXa3ez40oTUJISJbBrvDA/yzyEUf4sk7W8xGPkO9vzcB2Tcvb5r2
Xv5ZnKzOulXGQVALrKFpKFo2Dwpvp4zCB7p8nAqsnrZv7tz50QLt/LunylFVIQh1
sUx5HIb8zpT6PWtmItmy8LHDSE4gFNLOsGTOHwvIGVxXJmG+cFbAljnTup7rk5I8
M85cHfGfsalMlv4tdJmbcazbOAHOYpq+zOPSdZsLT1Q14Gz9sZ+C9YY+xomQfHAk
m3NFXqSBlMrwLBX7I/l59Wiqw8wzNq6VJFUZQfk2i7kyGbJc9+vRM31JSEIQtxYi
qyH8rSUL2DPaa9NMVvhtyRn+XqfX6F6lnoOhqYT+VZeaFNcHT70qv00ZnVOBij6j
rGZMV4lzmb4MDrQNmyR3JtZa2S4/RdMlW9OCymovJ54L435dOsBFFdwLAzG/Ex7/
jqt+xpxXP2owcCYDgEJSp4lFafOceKQ+9aCPJYIUcrci8/EKQzRV5cENiz5CGSt/
ELl07qEFftDVzoJ6Gm794TViz47nYv5L0WL/4D21HjRR1JQbrfVmr9nfEHk/xjBh
idd7yLW/wwFlciF12ACqSjDIgYNfRAKCbST+araFp29kcf0xlKlW0eYrPzn5/ThD
GpErq9eXbP/flE43RjWry5QTyo6rWU92lknAPwfAMzXIaMNzv1MxLpAXSuwzcTsd
JQ3HHYu/qpCLi5R7TQtKxWtclw2y3YHDj95uVJAQP/Z7imI9XKbvXryH1UKtbovv
jd9HEv15rSsKJ6xRzY1q2jmu2ZV/wGOLujFMGRGuFlKYY8rg4XfUA8IA2eAboFsj
gsge+zDbYQc2pq5uutK7V/d6Cg+7m1jzDrl3bqf4ATwEO+y7cd9/nTbnI7cNab8A
Qz0G4nIjEXCC+rgXAEKpyxwHxvgpuyFlS9xO/IDECJ5JwobCjPaTxM0tcOMI0S61
5XZWad5Eu9yu6eyFCMywmmUIpG7KTOvAqzjT9JMhKdqYF5gRSSqQA5M8VerooF//
KaCsGWaRbAnlS3BQzTnDXPkusoqh1l0jRxOlmsu5VKxRl+Er1wQxNN7m3+oopBAM
5Br7QLwwKZDdTOnGkMClSkdGWQ7LrFg8hSco9UJXPD1kg8lKqZb46ZDLBOMFtIaT
6RKFYfE1lXBYU7bvniPccVbPiax38oq+V6YBC/CkUqrzARUv4KS/QzKf/tC2OVgI
4W0Y0K4roOjeNYYpCQ3kKfiqey3L+hq1EQPCMMa5rO0RN5e7JF4EnP72uVLm9Qgz
hiyW+qI8/XJognoDo5AAQ/PUSEXssUqi8DENox3asLVGYRAbT6ya4v+M5vhSVoQY
OJ54vMdlF/Uic+luiWjzZxGzIndOrFyshmeBf3+Nk7DarkaWAmgvOP9C7gwq4YDk
9AsYiTZ3yFwgS+pVNqaudl4CsoYC8um2BVGEMg/BAovgz07Jd8bS7OJ81JxMCAnQ
0HzadQItEuFo098bQrbTWj+Bb+BkgBf19qPmQUrBQaPpQ528MyOj2Dwp7e3Urp9m
86Z0DjupEVA2S0JrSGRjusdz3ng1DMlF9ywDJUIeWWXf5WUvbODJrzteWpkz80jl
Zal6x7R2O2pShg5RtoKggka1nlJu0eTd+OeRICkJ8M/YJye8xQiazBZ16TyQd8Wv
ZyuLMXRw/ANPQTZtn6NPBZ/sn9sRpVD9pORjx0U3X5bwj6sufb4mtnairE/XYVwl
RWPPqbWNDQjwMs/TTesNAqD+IS8/NgaOo3cX3a8MD0lYnd9NZDUvWwfIbHcMfdY5
d9C7+l+MLsU7leH4NnNpXG2V1J6gEBm1dSklsmv0da+TpOlKdza6jCtoQGN/ZtnW
Dve6zt6YBenutdV4TG+eFbtdsroLTlAawc/bnvKY5RB2xE4Ro3Obkig90yQrMqtp
Sfc4Y6S4X8Yr0uPX5AqpHhVDrK6QnK+JO+0Qfn/lyqm/UrrOPFBALUW56QDhKmIw
St/oDlTQdqhbb82oPvAs/nRm0SpZhEaqt2KaEMMcwFtx+1cFYAe4Pj9ZPEMbJa1x
rhSWxV4c/vkrkbuaeiil1ti2NZSjQD53jU4MDXe7V93K4ipWWm91K/rhuHO4ws3Y
kgd3ftzsHDGxU76YmybgH5L2EKaKAaa9x4ZoDU2fphTVuOAJ172NJFC/T+kdglri
95afqYRznj3cIdeheQ9INRUGHVcwbD3WUSmsJdIA8B4a7R58txMPgEoITZ/5LABC
vwZu2rFuiHDV62MUGjpqdvZEOmAqMIO76G6gsJyg78KPMypqjXQiRi+85c1n0+56
SeJIUInaR4RY5CZxL4ssx7zDOZmx0w6+onCmos6OxcuIjBKrnxpDpBG0jcXSe1iD
ku9tlR4WljP6N/6GOYMjCMkLmTu9yEWGRWoWT6FSeFzdMVoIUorOG/YOedR4X23B
V3gA8GRS3g2j1rIOypP6hZ9KYfeKecP9wDCnKc8mPmiADc5hZ1+Zx+2qdm6EJtVA
t1/QnOp1Q2/76DMJVuxmFRoo4TcCoIOHq9dw72BE2o7lz8d20SuOW5VWz43ISWjf
qK3Jsnm5aJ4AWx7atVzTlohIaHITE7DTH9Bz9XVFMHFMyvqFBy8deg/dmwoskexj
gDMpUxjlm9FcTI3VlfWk8QOiaSb6K6+Q4zGE7ylHP1Q17wCJcqpQzk/EFQoq5DWu
tODE0OpVM+cjAaiyQInm6Y0+saSAcjb/UY0w3x0WIBy4tHHqizmtLgRDWhix5/6F
QL10a7Pbj9ckhsFsPScrIsTcm7dniQz1RNDtu3xCo+3UafTVo8YVYQBZlT3GwEnZ
LGP2ThPp6ek4mpamHDGhyhJcSSaZYt8ZjkTvQXwv8y02Mdvpuo81IRJ1WYbh3awk
PVTT0ESYsunEFTZGxCW0d+Z8B+QwONU2WDquxF9qQkjXQIWuVthbJnDZiz6/EnuP
GMThlSkgaY/yMUqytK+qZBx9pHAm6awpnrtYO+Dc3UWYUKx9NVIUIWq0DTZX49Io
0HjAJvii9m9ZkM46ealqKczbhdHN+zE8syB1RDthJIanOhsq4XRHBiw5csdvPMDt
CxQEZtXFX3yi2GwN1hH7fHSnJK223Gzk01/I6TKr0EgF/aYZxmrfk+Q3/SN1oswt
FaE2jrhDsz+ofm4pP02wvuYoxF6Qy6hokN2CySA+igJ/5H5veHUnU87KAsxslLxL
Lsd13MkKU4mYKNmFVxT2lWNvIDPf3ygyYAUmKIY9MaX+PExX7fQZvmhxRF3dGRc1
chpCSL5iXIqc5wa48w2tODLd0438WPMvt9sjTfVVA5ONJBS/zobnCFzJQutlwuix
r5o6Ni2Vk+0o6ryix3i/GcLhvA0yBmS1bymEtC14bcuzjR11bfob3/g4sWFMUzKv
Z61oKpzmg8btH1krzKxsMm17AAvAThA6hUUHj8CpiC6+sj6q6ZMWJkzS3aU34PWJ
L5INPKLqgU+GynO+PSZ2nR1vkbI3LSU0ktFcHawYbypoMbsKiud1gURdviipaFBt
E4zqdTv/znJx2zS/i/DpcMQ17SZWdFarxz0YFez27MncEqXIb8Ze4BsMo6sQTUol
ulVoX1fPRoiMIibnKAkCdf7rSjT0C964QJyqQfKKCQ28P91Xl91uJJPgEUNDZnFC
+O8sqEWOL1faMeXrb/ivayOBUJ+A98p6W40igwhngcCOwfnSX09I8nDSakdqxBHl
pPk8vXTAfi5b/Kzfm6EIMVddsfs35m5+yaTkUUxXmjftC/11gzuuk4wVtxTj7jok
4IfvaBfFC17AjR1x8zPogrkYW1sdB34UqjfnDCG/obLVJ8CT69dGo+8hkn2cWnQH
SKJE+T+7Nl3PvS32crnc53Grs8jp4oiY041QonxcHqX+1hJLCKhkQ97quy7cJErV
CxppHJRA+gy2tcee7q1lomfDgfe5toQu9kyomV7+uIw5KbKBQMCGWTXxwj+hX8Hn
34GNEI6TuBw45gxxj2N1ivqGOwNboTIhWe95tDrbAViU7bDusm9JSz4VHqiKqm4u
TX/k3sYyf8VFFKevgim/OcG1a1iONDw2dcoezY0OVS9YFJ4t+90P2IM+FyKTAf0C
lRPW8K4e/Nzb2GrYSdN2TzTL9eL5YKeRXhEysPV4yPYdc0Ko+FqxTIYzmDDHc0i4
Du9poMyew+Ba2MdeTI6kIQocWQzOIOJOLp0sQzt+wtmNKSnITF3sc/N3PkZM4v2W
FTcoZn0WcaaMpDXD7ZFjGmdxxwAfBiCbGRzEUK1U8anwgsKUyHCj247jI/FSPFr4
1rLqnkWfVAWHi92V3hcD2uCYQ8NAjjcVLv85PeTXQ58flJwPtnJXTellXnpDbzm6
QU7lDVsrX41JbP2F/3bS6X21KGViH7qvVVvoBrHDfaovKoFxGl3vC+KVbdvWuFn6
WJFvEpjKw5zG2y/uGpXPfckASmer5gNe+eC5GuXTHSvXnf26E6tD9olWmAZk+RqB
3nU1O0ErDMVg0bMSPp1IeOoG51qOtUD09FtixIBjiW3jU1cc8Z6FPSsPJDK8cCBE
6W8B9B04p+1VjkAh5E0M88OH8vDa29Ak8tqhlk0HfujCjs0oT4K3VaRPfj+DCSnx
UiP66VVGaf/VvJxzutKxq56t5EWB574C/8EFdYZQTs+P09iUpuNAGssS5/vkmSf9
TL1adxpkLCyfbE9jRrDSsl46v1A5HcPEfzSn6iiiEMEpbLIm+JNquXamcqbB4E6a
r219Q8N5FeVUUMdtib4EF9ro3IYn2B1ZtSp71sgx2xAo8IFKGJvtQJjDHxXfwnie
nRkjSbj7NfzwKBax03I8UnigsWToG0yEoTRzpso/q/BFxjNqSPizcBCkp8BkMXo1
CSNTgfa0N/O2n5YWoCJHaQdlGR3fBriZcUeGxWaYPiv74PrsrWcAV7PeVee7fvpA
jrHi0n+DIXvoZyWhDd6r7M69qvD9t0Xb2ZHdV9TVLZwiVtRotvToobqV8nMGogXi
YVSBSKruliyO73lhf5jdkOpKQ9k2o8E98PCPKUStvE0hsCSw5vEVsIWq0ZF4DKYZ
Gbh7mar+PWdQSPd6PD57z7qYEshm9qjo+wVk8Gc5jijWMlS+XU0jKtZHVwO9x7xv
uD+ohSVI+4qXPK6okCnrTpNsjSmgV6/v1SrCzc5wrXsHoDSOUSXU+Aa1SCvcdfyv
6HDz/DTk4PdfGL1yeWn6VlBK44Aj0VqEkvGjl7onmCmPYxhUcXEn366Vvwg7GJnR
ieZ8FtjWMo3hLcpct9QHN8SmMPyUz4iDyASHBwdKz02n0PygCmlh+dtjcRynSOHv
ysBxT3A64d/FXtoJYtGGKXnpUlU7kNahLB+7s6I8FIiRWV2qVWx1+AxQeqP2srFK
G2K/DB65X++QXR1vFNeH9GrMoLLQSwLfy+g3AXXdkhA/ZI4eSpR7d52wF7rdzyNX
66t4z7VcqJs8tQ9TXL+upT2n3y1zypng7yKeLH5bthpe3gicxtxalfdWDPUY45u2
XQg2BZonc2xogmaLCFKM9lMBXKwlYWGsXlx6cumlcTE53+QHP1Wdib1No53njDTZ
Q6woBp2ZJ3yR7RkxmQuXm8wFo5LYCcaZUg+fFyR6AiieKBFa1FI/7E63ooGZao/c
HPS9AHLHf1pIOuiOEv9DA3E5UjUuntfiaN7p0qntas+ik2pFJI/5fs5J16LV0d4A
jOnY6/zVOJevBNPxA/SqOsHSOA6u6dr4l5VObH8XbQllReWPh/utqpKo3hq4b8gd
eSBEKbdYb4sQjKiLd6SEPNZaIt7KBfs6ftReo1CE00G2bzKS5hxZ14VDFa34a8GJ
iyU0to3isgBuDzTGr8clKFsu0KuoENNEobykF53T4ZffX9GQY/4W3+lc2IASyw2t
GQ8Cd3hJTx0wdKoCS6q/U1MSnQQqpHouQuvy4vUBo4ESveoc3KrMPgHA8y+VMa4Y
OQrwI+8HeVcrX0tPg0WqfHWqcj30X6jgABeTEkSzs5bGtzGA+f4rgyz/jtBaJO9p
qEULh5LDvhthSkIDQruJGEscDiKM8QYuFexTarNmD5oFN4dnQQyfkK0cZxbNnLRX
GeL4UFGiiuanlVbOyOFULvN47V7w/YgPjgCnXpc996dAfBhqH4RFSLgmyRXJDhXV
KKVakuBcVpfyK233c7YkBIF5sYJiDAD1c3q4AMDmi5rG2f5ImGcm/wRjUKpFvaCJ
suCfsB3efCeLm6+plYPJCfh5YzxbN8xq5ds0CJxtznmQFzodByYa3lt7TYHnUxVO
wOeLTu5s5Ol1HwUoT8n90r7v8lJ/u8XBxVP6Jxzz117VBT3/Ft/MrC0TbGVIVz02
nmQbnVMPLTfuM2/yr4zf419gTIDC+H9nycqELeNysRJ3o3oyts5EVjRQFGvk2wjG
VcWsZNRft3TYitF9pqAjtVYHTfH2VKtIAwqPWBrzVm5eaxYtfMMGW9eA9a+kn86X
D1eRHIsQUxaAa0p2q9yqZKE/D5PHY4fFoDqAi5jTUjV6OJ9kagjbstbcrR/S2/dV
tnGZov9uoQSlDa7i4pD7UuzNcXvGr7OyTTct/MoQpzNSB6KkMa5VrFhiyaWpOxXJ
wrpnrWloZQg6hDagXDVULt8gpXKjVMGxPyZwuolA/mIayjvMxf1qbFFDDNe+rkus
w6DT2MkeCV1LvuVeen4Ps+NF3a+effNN1G/AkTfQ1s0jt1vy5imvdY13Q8vs+a/B
zdk9+4ffLgEfW7qkiiJ/Ai+BDXNTRrhd08X0PAcaA2cvpqvusMOp71UPgFNL3sCz
aVQl4Z7G4FaB2CPD/PfZ/5n334piCi6/CVbrtPcSiPNbI3Ett4fGS9g+5s0vf3A9
vk16a5W5GdcfIuEKVYh040/VR1fwt7lkid+QK0m67eEu7Pw6C4tWEtjskeh9ON4b
ltU2S+bKus1X1QIKNVBprMYdcUm4V2JcUAPkxlRkl7JE87NWy//enAeaclsTcioo
eYwknRtqUtUd4PWKCUeNRKQmYScM9SPcT0zf2Gx0ZfHYNjsh+DC/NPbbdA6itm4s
Ki1hzpCmR0kg/7MiGl7ZUp5EIGRu9MdRdMOgy3k7ZTpRw+I2/8EIzNCvgYbOb7Gx
qiQpW4Q+quTfzragwcyVFcVqsc2TXhIntY4E50m2qfHDJIXGVOktaWN8IB7Kl+W3
Aqhke1UnfZC4Ot36Yo6DVVOk0jrHkX82GepEZKP4hmzou1BEXo3q3Z0fVI2X19A3
QU14yAgYt/adXy8EL+WZv5XIoiRddPGqo/t5KhIp/WvRB/h+3pzOBFPz/9E8Bmvj
8Qs07tNC3GA1XEae3XCF8VWO/wimlyo6hfrQqcuBrbgKDjFMpDG1+0UYIkCNH4xQ
Hgz+VgPVhoujcI64zF/PtOvySLuVl5Vwz7HUrKWrsj4124coTP5gbeGra7QKIx3z
RI85wz5r6ee2WPSNds4kuHe1RF6Urifom0d/YuBfePnCDxjSnXBTJQkXDCvAQJcj
wwyTEYIEwb3qCym6mEtbFMO6hZP3BXyxI46Xvf6I3wzk/gMlNqyoLjuEA2QUl6Mv
Gha5yPl34K99VCNZ5ol2mk7sqRn2lINgInIVHLIk5JHcHkqW1U3G6YW4Yy+Oy8W5
YwK3xIM6pmIb2AyNZa5DzuqG5LGdpdQZXC9V9sW5Z42DKHoMlQ98LY7jexqsS/RK
nxIUxOkJ9fjEfHgAcTmOWoTeJ3Z4kiQISqRxr37tT1xY0Ry6x5/eMtS1XtJXhia2
qi6wXYzqGOml4F/z1/k0q52zE+zoZjxxzDB8Xi4zTtnKFsD9luzRGfAbu5bOzO4+
riDpTBILbJUSqduKp3qZrnYQyIbM5EeUkGXmmok1M00iNwXlkK5qmkfvFQj3oyMc
aMxKA7LmrjuRXjbFFzLs+DcpLVN7nxEmfRZ8QH4kn0sTs5yT3LDPApLT6bq1fIp7
hsBqZxjCsEr0Tgsxakt8QIODIAqbKAazWzmfz6tTRrfKIMbQ/Zimv4FPF1+yeU0j
LnIKkeu2gGV5YyvEWmXmabVPqTNPVtrTGbNIn2DjNK5t0d5l3+wJrHhzeXRPuNFy
vfvBjvk+U4ceBu9RtkTUOYqiFvin1JQHXMOImBLVeu73P0Scdli7M0BQhCDirwGU
bc6RMoDEPQhDVeOhAO1hvn0l65aJ/dNiztfTQjeExMxQiorVjCZ2K3bSPNdzcm7I
/JC88TN/XwAmVk3jQeNCaSBg1MRm9EPIvjsiFufBrQpdy5ckWaMDZBklz84VFMIw
+RFnkjtEZ/fhJFG8KnWYxup8u1w6G1+UmqDtIobth9YL042smdcBu5AXQPb+MDNy
lZ6nN8BBbukVDHXcyE/j2UPrRHQ6JS4EwO8EdFn7oUo3nTtZzHqmxy4OFnYh72Sx
1IlErHo1j5xLm2yx0GBpzaYzQDLpmexCEDVdF8e4uMM4AnoilEnWAx4Q8tsMxW0X
ey3qTugMUuwHiDRx2biKzhWG7cpghLskJR83XLv3G9N7TyYO/0ngrDA5lPO/C5Dl
cTSM+tflEICfcL3YyOuDF6DV+YM/K8cbvGKZ0ivj00CTLMrUSt3Mbn/QjpiF/nHr
jnljz3DCWpuqYasmC7U5H0kSpC76ZEvrcmKSA9QfLDlor2eiQC7PmYzhkoFOOa8Z
vIV/NWuxi42Qo863UdWCMHZKN7R1u6nvjYwRA1A01NmqHoJ2t3kFktbruHCqg+uu
4e84W8txMuNKsvozrpswluzNnjmASzwfu4jeaAc+wW65VWVW43bSdw7Xr2Qe8lDv
tMWrBqmPcDPVpA7WHh4b7H9OfbSuKCAChieh753QwfoQc/Gkk5xTxkMXWoOdMTho
Vvit/axBXv7KdY+kP4f+zFpQQA6CoLeZe8utABCVVhdT1hM+jnYOssW7pE+2rnXx
pf489zK1DXz5Eqxdwdrzj7vzhcE96SouJmpIdzmeObigDpPij9s980YsefJvIfRB
ragbahPicRFkpj0hGGDOpfI8RLXYN7EbXDCJKTzt6HN4+qK5Tmco6eB0DD6DCbmG
6VTwomxl3k1778UpLbujmnWUoaSkyarqKqX9ffXQnwWnIRl/PqTdCG1VxsQk8Jz9
C6bk2u3g7/ufnuS+2da1MoKiVMLZmogCBkzRzda9TmOu8493NxkjlATMcQcTEm9o
wbwP2OmhyBf25vGyXItYriTOjcvJ2r5q3653ODdZw15DEEUfFRv+sLcpc41sIwHi
XyjUuugELlSNv2cRdYfoH9N7qX+mOFlXY5HAfG8uFWfoIpycZj8QJTXB8+Lf6jOf
58yARalcn0KH52mwO/NdVpShzIMXOtvtNX/rPM2QZT4jhN5Or1dXe+7wrbuykAQE
UGv9MgeYm44qCMsOyZ8adseVxMK9lpwZb/hmt1I+giPDBk68IkegQNkQezb9FlGv
BHbgLMiq2lRNT0ghYJoqfoYCdw5ZZw2sFnQnT+DD+3ri4cyMovxHajYzMU1cQvrQ
H2dVezE0v03Xqj2HZ6BggZ8vqhJMyXXS5wxQyfndVOxqQo0EEsyDKb4NJ5CZAzMq
O9lmrPLtq1vkpxgdK3905b81qqJSny4ATf9voLt3m31EZAyDph7LJXmThAcImKU3
kgbB3WRgMQYCv+8HCvgP7nKyV9j1lsMkyNV9qV3CJzwEnEE35ygka6zaKX0dINq0
zEB0tVEnWI2izBs6E5NRWrq1YCYuQwBjVMtTTY6BpOnioZ/lJ0CH8NBUL+LeCkgL
Qia8daWDkhDPsMUmVJObyOuNEciIkCO+b2eSXLijzyLDpNXPqfRx4fygPKi7LavK
Vy3pTfhMcs5OWZGmtD8P4jcHGhPKmsvJKGqDJEYDzg/GJfvF55IEFWwU/kGn0f+F
F0vDB1kEmhGslJotz34Kb0F59hfORIQN+uAg3UIGzC7RaC92IEJZKC88BDjFI6Pc
Cao1mQcq/Qx8trqswtDXt7d79VtN1KzY6LLFuqqU5ueUqXkF6/yjayS62KQzjeUR
FYVtF5p30m57w1iJprmoZLVhuGqjQywz79Gn6PhXBMGbJ8moa05ACPc5HhUi0DpF
0fueZm9Z1rlQZH5a7qhXImEJakvEs3fCEcTSAjzxo0S2trpw1i63a3Msy59GpcIY
JKZ2KJkWb/m4VQtgLgkS5pdZHxdwM9dTgyGK/SprPRErk24yVbBZtBFkcVMelFMm
e1wf82lauFExUnu5DGW9liVPRg9XS9CHAJk930LWzf0Nsd/ZjeZO181q/3QamK7+
aJo+Bx6DDjYTY7Mw15+wc20Ke+12fIbZLaLYkuzIgGpprEuZd7KxXcSqzLUATAtU
i43q8dULh9NR07KuB2ZBr4ZCv49xJmjvZXwd5gaYlMkYczGjPo01V/fdCxTr7Ads
q4MQiaa2Cg8SJu2urq9RwRE3RYWCEJm5uY7+yncOTu9G1ZLsnN7PJszYjLROC7hb
jr0BvViFIiO1PPz0ljDMfYe3OlP7ydMAlS7fngs4yozjchqwPY7kqR9tRFtwPU0W
uj5meuUIHOmwv+5DN1yd+0QDGS5LzAg5988H/Pd2uWPMgza4Hlc1EozSlBv+awsg
1kGBztYHaQ6jGjA8bFCXEQMyXLIJk4ONPSOLEHPU/ed/kqqHI783Ub2OQuIzUxEo
fOGs4t98jgRmcwruMLtFSpam+PXejNx8LFhNs/lFjOjE0fU7Z7TUfaHp7sxGpYes
U00V6gIGNFlZAw9Syvj2mgbxP0cKRuOco6HeKMYQu7XdcaQFXEWJw1Q+VvF1+/eV
U61ICrCd0eE+JvFF9ikTAFfOAaNf9f4RqF7zpUhD2hhXpGZlIsMF8V/NfM5D2Mu8
pWwiJttj8SISJioLAHxxdNzbUAaifIJx8bMaCA5jacR+YKWi6ygshM0svana4F1w
k1P+dq1SLSmHOBt4R5U79darDacXlSgd1vUjtTEMVVC8ZpC7OoYk/4FnvgLOBKiQ
x56OsV9GskGiOpRrnjI3nU/0gI7+MjiGlE11rJFMXy0J8p+XK6Lhcp8/qbh4JlNk
n+jZ385Ougc12Q+p6gFG7SQXRYOJFlAVQKtSygn3ev4UZac4DAt5K7cIUn0UIbGD
BCRNGofcs05ddgCS2iBzf0zwPeTrad3W0FJolaoadqseQaNoqKLcKMKW4pWLG4DZ
uxxKlv+MHngej3K7q9d0ySDS+/neh4H0Au6CaSd/HRy3XVG3nmNqZOtSOGDblDls
FqkG+2FcXpqlSriIMGTbFIoUn2Na/XJEO9SDOikMr8j8z7XlBasEPd9YodEmSbwx
bmtYL87/HcIP9j2BgnWR4s13Efrbdo+sI8wJodSjG+WjNBMJAfloyOif252m0O5N
8j2JcXSgXR8IPhc9iOGZaC/fhf4yALpsk7fpPKBmElGniUbxZZa4dNU9Wpyu/YuE
s4n8LFnFuu0RETftfPuoh4ZsejDTuYzljwN3CWI+rlEE7zLCiYFAbZfm+BxS15fN
w4c4pTRHa4AEq8TlEIZQvfo7Y4GEBY4EIPLCYMYjiIugkj6o4pqmM6yX7u45M4h9
q61nIXkeW6hJgLpja2uuucnoA6nfsagtCXlWBsxwUDvnazMJByxOrJTGbKPkdQJp
k7CEqwIarGwc1Z9WYXEYhcqG5Yszw0RErwD0rvzeNY2kON4Bst/wcj1j4hf0HhE0
tBY+76FbirmxHNiYR6EFhDyXtL52viSAvdnkhhLcOKpSiwV+z1aisi6nsTBOcX/V
MMHA+6Brv0W8zLaKsg0/kNmumLSnRl724YM4UT7oLbrNUE1aTn8T2ovDHiSzfR9H
QSxl5/0GxieneZE6Yb8OoHJwICLnEtcOTx0Xr2fH8VbgSHeRX19oMpWYfXdBbGUP
jCbGlsTWLnrHDm4e5KbkJrLrA+lCI8Nu8QY7NE/Op3JJMO9GJQqv3qdKaUlddHVu
//LitDNTaKtOChaNdrLP8sqkTjQggA0ZkO9TbFoxRUp3utm7wUUzFA/s6wE/CCff
sWHlg52E+bAONgQ1Lnng+EgEeX7mDFTxaZBoBQDCJt7DtL+fiYswnjZ8CEmHHSxY
l5G4ddcV9zkrkJSuwLOzHNtqLzpL3UjHYDo2TtWQd4ZAjpwBA6bbazoTcDb8/mzw
Q9+AA6T/Ztdenq4ma4yQcoyL0Fqotd/JYGc9co6OrAZ9QdU/vXbiXvjktElxQ89p
fgIhQ0WYoCKDwGXE+3WL24Iw8wri8UtX0Fw+DCECkjEh9GfcHwD0oFo8U4i+Nf0x
eJ/VovmA0BNi0XQ4xU9Yoj0gRixfX/QTGocqk1LZ3tjrYHDEe8aNJoGT8jwKUxDp
rv4+ZONGzqtincr8qAE2Rklep7nW/OhOXtCFN9Qfxerm+V4nZT23hM9eTdsrpSYN
CD8w1sAi13Ae3FFEJY8LLnoja8fCnl9SAlSu0OF2XOyM19wL8zxh31YcOyoefedZ
+32GtviNg1USX5Vlr7T7LMEYE+etg9Qxeg05asiWFedttWERP3aIM3a40hYAvYfl
q9BJoQCMdhRHod2wolb64MpWHBB/pEyAMaXK/ENrUNQDbUqAXOBhIv5yDAa6UyuC
JMk+QddxY2ptKACK5/0S0whTcx02LmcCxfZ0++mG2Lt0FPGFoE0ltjtbW0aw0shy
flfU/gucAiHPmqUR2hV04J7yFfMky5oM7nkPcFxTN73dUcFJ5pubqbzzjtcvgBDy
lKH7b+ikaxTpR16s5yRWoWdW5BOa+wf0ciiNMnZy9HRZgRtp+IR2SWUE25hN9puY
jlP8ZQoep8QvIb/Smaji03aSf5WEGaqcGOC83G0pHokbnQ6ukI8ROzQ3AqbtECyz
H3kGWMwnLYk8vEOnge7tAqYF6D5WdIR6lLKfgC+WXDxT0k88GS34V1ceZvlE37c+
3e/R0N0rv7o1x0IpitiDHEAHfP+keuyHsKhWN1ky6A1bW2cLBLA5dEG/2W2MRTVw
6bCyZJoWmf+O2Tu0cy/RoiK7CqhjIgxkhpqw079KoMyGKDfU1ihlu7HXTT5kOV4B
v1JybQf8MJS7mfrd15TGR3p4c+reYE75U6+7UdGZ95ae5T6vW/RHa4ccD9FovUUH
9tfM+7gmZ0lqj1h8oR8SIlzjlmOrB+k5NEITfFSCzjZtrbRaNI6XOc609bBRVaE9
CzcQlZQbusq6TJroVxpf29MFBc0nVfdj6Lkrl4N537+hFAATPpMzztnOtAUno6WN
FO5I4lLHOcoxV2XaFUFtp8h6oWFAlGeMhsri9eaJT/HS6QHdtQgzD+42zQsdjYhf
f34Zt/nvMxxOTTRICz35INn0yxt1O2tOyxPdZDonNQPfT8rLqb+7SNMl35CThS4q
tfuFqpYBPYaOqx/q2vms3zRg3C2sQH2OI/+YmJN8Bw1zDllN1ZXcO6UG11M2kFWJ
dtLhF1TFoL/KSz/zJhyneXPBwtdR/5NN8IRGkY7d6UI/No4hcYiziOCb3omczgvp
utxIOpyujW4iWCGknCBgo8eanoLGxhgpT+xax1Hm4dhwcgAwc+Y0SjKKQ4R0rxHi
qa4IEgBdhCCCrg68v1O7geqQPLwFYF2TFIeJdY2dm/v5CmgOeCdtDrDwyMoj551B
PjC19WI3cTtmnSEHqk7JKmP6rt+JypyR9faAUKLOwDRzHViKXoaicGTgU491E/Zn
YLITvZwIhvVcjg7upMH+l8FSXwIPvlO6MQryEf7zTIM6xkM1Z4+RPFrC28qjQ0Ki
nZrsoizZlq8kNbzOvZXyx1I0pZNJdOApkBCDk7wMYinrGBBy6vcnNs6iEQqQ4qx4
sY9TQG5ssF2+5GfO+7gdTQ6FPxN7wg8Kt+DlOm4r8EHLS32XghgicwY0NX5+rrUb
ssXsBdQgZOMca3KE2xjYYsTgo9WvswxP1zks4ukkyAVqVX14CHMUpPtHhdNzx4NJ
8L9j3i3Dd3xdXMttdcyLZrHUrus5hOfN6+IKdtBP1PEz01MXHf+GkAAHjXF1ciEJ
TYGqLJKJOPDM/1ao5cba2B0tCYy1nVjUHOgrFfgknwSIfIlu1djLI6U0kIz8UtN4
ZfxyWPt6m1G5NL9xud4bEgtr/K0RSdi4iuyjnk5NEaiCDKLGiOA57/Uy7S+lZNz7
AZGh77ykrkk9hCbzvLYsT6im8MQqe1u/VSEHq+CqBS3G1ao7ZCKZPPxgN4ekTWs9
faFVebA317lHMW19JfVdooa2btTGQKFDYIRrg29+7YsHzbk4XrebPgSZ/VbUy4f4
splRjT+OdWex4Yf7i814SxUTSfX5xkqj23RVeIozJSs1lWMrlaEPwgQ02bSxbGxY
nWdFX41FlkMN+3CzlR3MbibPTomoSWbgwmXmMUSxJpz073ZY9M/qVaqoXuPG9azj
u3uulwUH4QPAwNuPIHh3ZQdLTkFJleyRR28MaqeGb8INj4v89EqC7qFebXfc2oRy
/kkkh2ODn2fwzXcNaTjmYwQfwwll5SlKObB0GIlGNo3iERths3aG8N5AYAGFGA7t
sOJVRHYrbtk/J0MIjs1nswqqvR8ixIavPYI+qfGLOxnkVxxDK49TKVGmvhon5Acf
G4wPEnNHqHjM9Rz8uaGvMzf3kM9vNQ2Rhy/nQlNCWXw7tI5RvUwcohtKG1Q6z51g
Tyb1k7jAHpO0PcB4XwXBEwIgqd6fGGtV1OH6Dhaa/W1ffUhwastax/X4PfT/eTxp
QdnWpbM6dASz4cKY/x0lL6OABD6lgv35asAR4yTM0OB2ygcg2d9RjftmbvxhFe1U
v5ueG4M8Sme4TFzBXRjnxL47ZHrnlv0JQCqNnItNp2c+iWCENfutVhzS6YCg1y3m
QwLOJudF9reGHJ8U/HAHm7dzZk/6FcJzkh0nXfg/Z2VeWtM6z7szxIOC2CVdi5H5
8C9lqWYaWYSay2EI5rMlGo3WeSV7uD/C//DIh9Fba+IY5ECeLmjSOfUddzD6sMBg
XxkrOVkWB05B9raCYCvbc9LnmsEZVm27rCsxZu1M7+5AH4hT99e13pqU4/S5dDiQ
ENCs2uIvNgFYou9q95Y1UdAmpGOkWmFVP5JOCjsiO89CffLGGls0RmW/PHGWhBB/
yfmemvfj1tum7xjBKFFuNJVupHsBdPe/65P+Ab4tmXKirsD6czDrCuA9KwGdi0jo
Ryu/RCD4O3z4JBIZ76oEpHtD8TSffi+vupZW1ZJjTjkmH0iK8aIwMGu1m3agLVQ1
6XFp/RHkI+4meVpL6uMPdM5tJQDp6UyjuBcM7VeGzWYFx6IY+oymk6ooD83m79oC
4VzuSAsHPR/+cpM0Z1bvi3tnIRmZMoNZDvQqWQoaNaEX7gH2l/54WAoPrWBFy590
mlvgfE/Xp2azoy15T3mFlcUh8+BpeA4w0xtwndSD61saNtt5zJp7yc0Rw+zotRHt
oAQZwYGP4EOg+vF5QrXIdOBhmfm4/hhZFIoizkN16MQn53JuiCfnueqlXKMoikPW
5t4JKzKb9PFKYzrpVhISfE2tDKwMw/HkKB1RPHLbHSe7kQHzOjgvKYKJJYDkJNHa
VF+lnxTBYXr63496+eSEHPI6KfZxb1NY/gjJXe6DW2d/fdx+Btz/WsM6nfV+7FHw
KWdgmoFi5cBMYUGRTYP2QlgM409QGTznlPnikV+diu6ExMcCiPAGNrWUajVIH0v1
ynnDI5AlUwZbbW0mRBHcdb/E+b0wxYUYFlJVzhYkj0UjzGkfIUqGE6W5fkhyjD+W
gm7/cBrJKIznFmwVYphbPNfdi+ZdEvO1S5MII8OVIJ/O1uWVRARJ3wQA/MpteOzn
EfwVJfP4w7ONyb8zuYZ3WoTsGVIlM5Y3sybcD91lORJMS0qMk4AHJ4TSaQAayqt+
K4m6rNjY15L7j2Hj8rsHrf4rFmj3LukJr2yrXBxSJw06NCAVx42scpci82YCoyRH
rQw3MVADjVH9Y92/LeSNDiVwQxqnOyoYk29IJwv0J6VGtBYCQKrO5AX7Hn0i2lRz
7IgcPHHtRpAQIwbcIqmnO6w5umwusADdGGbjNnLul5PUdXm3OG8l7Wg92QBpNUuV
5Gkfb4zH8yv0yDEEStxCJDuPqvsIxRPV1AwXGKl/ywEs5OJalVgUzrNA7a0Bc8yf
1+qQU2V1aMiEpr8TLWlBvVkCHrdz54w/NtlXiVoXdU0zsioYU0Hmg3iws2TbNbBb
PlgfanAhcJtaAhSThU1aXWAg8XAUYBinV3jdEIdf4Wr6jAOewmNbFA0MDFyvPOoS
gfr7D8igyfUWdT5utXhPtbc5/YpUcwMZzShHKQr9OS5VIO+50lopHErQ1q+0WKQP
PRwVTV8Kh2aaImjn5NMkbzjPDZ+UqYJyfSnXFkk46zsCx7fmgur1AC0ZzkX7rjNq
2KNpnYBzQfDuhlzIZ0m1T5VNqJU0HAx5bysUz2pp0kn0HB1D2QDA6zjewOM8/54M
xBEJM/ZKTo9ugo2fFB+o6L+ws+9n44V1ByGGPkF9bac6mm2qA2fdfDwXyat6/Gj+
14UTyv6fheF/w+v3WIOpw6CEwNUaz3UBaipTtatbWWCjDJ1lRrqgBoqdf2iabHux
344o3H9aYOQ72fVo3AlnJXIYjr1fYN6SnnzlRnlNi87QAnoAs2T2BuH26cvFS7gs
qgayzTu1pIo5fsBL2K2lG6K1HCleDxBL+N5ulvOwQxGeeR35XscR4fmhxCrevAQD
ZbI1OOQw57sq8Q6RvBOwkm+TfjOQNKsXFc5Nu1M/JesC2gNXQUVdBSKT+CvOjMEs
MoUz9QgSbQIsm0+W3SyogVq4UEyF4Dw34kjclAJlbKeC8Nv4KbmkFybDNeICzsoz
kn2S/9YEXqj6TKWGX8QOLHHyGKftCdJ4j4vvVQKMdlUFyxNKyZMRHwAenHiJzy9a
PHop3igm1lHXQp/+om4OKPiH5MIPtYVw/MTmtU71DwWYORcmNMjeUCAThe+izBjl
fWiqsKFyHx+o+0G9lWYbcEc+bqjej2reHF0nOIljNZ33eCvS3yzCdusuA1g7RILM
C8nWciJL0uQHOul6iMSJOHagsxHdD9Od30LV29forD8/1iqpbH3OxEWMtSMSbtRb
P8KuQmHzomzmS9EkZ2dip8GsJQkIWdacYI55aPuH2rnE9tflrxmnkN+jQHjha0E+
uLxWC5P1mnmEETpleUzCrOgY2Z2zi+Bs+/4ewq29GnyjXbdJ0LMxwfOYiDueFuCH
gIZ+AAAnL2mFtvCquSHFUuUvdvvEghrItdKz22eWKOG2IJv571vx+DODmCciuCfn
kQV7gqbyzAEPydlr6+zr1MmaQnIi3Qr2uMAd6rDkTJxt7+A3rX6VE8TtgGOLvanA
xPMJJRGqdRn/EDqs4HeNMacxvlV9GDrDZgFs93eTqkOQJLzjpHXBUBLWKPsbTxkc
Ewl0Ro+oXj9sYs7Y70qCiJR2ykWIlFfFksSrAyd1aeG5HEbGgCzfc47/rkdiMNCl
R2Ac03UyGjXFOtde1P5dcy6uYRMCuTavi0iSQFQ5QN6GfdX9iNCQ8qPY/aj0qg2d
VT3sb0Tso/yu5hf+w+aomg+ylf7fAo8TYWKWVTZohViv6qXGoaDSzNu+KFb/ZMcc
wfxBvfTJdbk7BzLKHYHQxIp5bDmYc0/iiTV7+WBYBvGT7KKaqfhG+nyqENKbLmot
n6ZOoNNLcxAXmlGjAGguvK1DqOTlWsLp/I69/qrmiu8QqHER537SHzNEhL2GvNe0
7w37Q+AXnq3P8c9M2VMFZNsUrOcQDhgW/9p+fOvqKREe8F/Ci5/4jguSYAft8lMb
whf+LGs3yb46VeibTcM+4xVdH5RKNUX9jIIFPmnVcz4CzUxUZZh3MzQzzGjLLcax
5edMebDi4XdGxrP7Ctwh6Ub1qC7Ief9vBGfcjOVDiPioprd4Ptv+nuDEeOR9FcDE
ENIgfVKzcmEAKDrvvj6vAEF71+kWs2vHPytVbY9DAyFwuzwhfvWfC3veUC4ZkgMo
i1UacSQGCYpax0eFqKnOmBfSixBslSuAZEDabLXj3xOfN0jpYCMcDZGGu3M9WKy7
jmJ2zt/OM9XvRPLXfa/RSPChxKQ3T9sCBgtRfN2ALktvGni/Sl7Nzm8kw4kVqQHi
GhjFaQMH1KBLky716vUxWyw8KcdE5JZQh9NSf1Et1gqJjvhy/WmGcTWreQBFMupU
OzymGCpLRoJNvS0HxTeHCIYhljarS3yjo7IhxTwtwdSELfMY0zIwbvLNEed45cVu
mRlqCM8iGxsVi4/JPOXajoTpqFJRulcenzUThVmZf2Lf3EUISQtd7dhmwFSUea6b
Yx6EzoXputhotgv55/abukT8vnBDGIcrpLuTV96BkxunLxGJpkk96IuugxjtamyA
Kqc4Nt8M4Ebqr/GZG3sagHNeKZuPcrxxYvOtS+5fqBLj/vXp0zS1W14blkDhvd2o
4lgEzHaMRgvdagnQRkxYeTzslVoJmu9nhckv+kBM/ZflRsNUFm7MSfqaAZUQk3YT
N9ozI/btLAKN/57fLKXBtGgHR2Kh2Z/phtERvhZBRjXcoA8VanIDM7lKHS8NuKGT
7p8aZLcA2L+Okl3IE7UEzUX2xuakvzeTnFk47sjqutQ6FVbwg8wM2cZXQAFZZ3ik
BcGJHw+I1enpOxcrQHYTvOlRWLF6mb8+HRHU5fDaqFyVYJHPA0jpLLBvmtq6CS18
2r7V4r3aLGoM+X7GEo/J6cgcgxKj410H/wzJCUigh6jAYaV4q0uucIymHbL/egBH
T1wIpuw6+tMgDDLitj7IM5CS2N4lS1yQc0lDpl2YYZS0N031UJbZa4gmpzsAbUnl
msCbUE0sE3MhgZ0oCwCYf0sLan4dM5q//DBqdvNsLmFWPB2z87GocUCwgZ29dWiG
J5pmYtICKZyvUxlac2BmjO7UzflGKCwzaB+e2P5jkesWVAg+2yqWe51cX+5IbKf6
/7x1V9tbRA2qRwPoUevSBFxc3LKyEs4gD7QiaKwMpZs9EhfjvfkWJN4ot7ZN9av1
//V0VFWhdk/Xh30SwzvnpxP0mdDpUUIyynxv8sPHkdIHE7tYE0NuPe+Ksd8Jelsx
x6jJOEy1UBJirX+aNsu+CJL+yVvJg/vlY33WFrg3AvoNr2S9j4nEnZxlRAH/I+S0
lpNzWjrSCbEVYPJ3bCotfOwFiyh6BQINTuXH8ZYfCm/CSgVHz9BDNv7BDUayb2yY
rNhskOwRHKnv07I83iAGsejDluRtuQDVyNuNWXQYxKq1n6UwJ0slhg8nzJHVXCyA
yfHBwaeGNS8ZY6uOojer50icNVmuQYLqxrwuU5/PJEm3lyAuWn2drzqZ151GgC2R
S/fnUKauvo6Je2mWAsLpDbSNL73WNrULy0bWyEovJt5ypIph8xQup9aivk4izvAB
n9UfkkVzy13qJ8wEMHAf9iD2DDfH5gmC28vcqC+yBQcKjxTaPX5cSwW0BQnVNh+J
HyOmQL05O/weR/GU0hvqHjLxNJ58c04MasDOgY0D4zTOFQLaL3H07QFRZbs73hV+
g2gsF+Hus/p5HHUKwsCkMMG27hLFFwTcNMuOlZWeP+MqporWeaMYNy1JALubmBm5
TKSuB+yasf/p9cyqj6/46vCi31oFVyPC0SuGE+kt3Dt4Hz43kQ67Sukqtu6Ourib
7Gjpl9XGnRz30yJ8jb0kH3jn59xJMSqq33CBsKzavvGWdhP+DNZx+fIAxkAE9Vbf
C8KCm0bRyZ/3jIyW9pmISzcF9PK5WhirNEKcp5kbwn00N3+W/ai35Hzn3ddz/jDt
HE6pv1Qn6KuKAEy4YBJeKmWZp871NxgMbUscsh7M1AiQaTZNsKQWszpQ8+u5/kX6
iO018jMxYRyj7p13OMDjLWTSvR+4qsQTR0nz57uX91vaSgs9FcBjHlYzDNIrZe46
/BdmAuU4zRnDdKJL1oeEBbVela1gErlZg2l+QKBmFcOSHAQn1X+1vKWOsJj3h4tR
sTlcW7lGQk7ze6WQZ1Zs620sztpZoz71Siu79XBmSun/dHene1K/a1WLNQYYZGlq
Pm4Mu0zrDJFjkFTx9Q1b/k/s2iIa/uf6bxU5K95jWdX+mdaHGq14FOPctAWr8s1F
yrB1RIqKrwcco/I1Z1ZjFo77uJJijtfJtruz4J2ESh3z+kPwPBJYGC0BCoqs6RLr
2jrSSYVhLmDzQE+atN6WRSJ9T4eJfaKh6o0ywPu0bO578tNOXP+gP6/YAD+RquqR
SQskFZ74jrLDZZQf37T1310BxQEQrI7PSMBwoGa3oWtt3gQp/cqVhCF8tsLXUb9M
3Ml8hU1Bsx9zCqIEtPbv+930wUK4UDKpDPTq3iNzqdk5uwSj8YzEDEt/PQrmkicm
/4YT6gcOrV4H/tCOtWQiS+bbdByKPvAVoqBLWgidNvZXlH3Yr3fqUpj00SeQBkEo
ICkn1QZloEcaDUOydKvSqZROtPrLDLH0Le5y9DUlfx0ty6ioMBq2noKLJhvIGUg9
swVxFB3nC3Ryzkm/ISUkSOWMjT67VvmGfONB7gSJaw/gyc6WnHio7Y3WsEYCpNzK
LWry7ikc3c9NcLSVo0rOoCAJWeIYZPHRvQDRGxRcUv9+OkdcmHdZKWZ3uCXr7/rW
lm3N2GCtkoXQrTuyGsITKS2gnsYV3nzDPEaTNklM9EzF+C5RExlBhBIVqZUTJAjq
lljSksu1mKVqmS7JT54o0G5PqDJwflWbRV9xxOlaBhhxnMjVkQJ7ZHNtLMRUIC72
cplsHIwtvanoiUn1/cytEq06z/P1TyCjw60YahzlnbOpxfImIOSMCcL2odTliHVm
gFKHX6+M717TcmlHj35EOUm2zn1+ha6C3ArCvHr0nPJDjnik6KPDJVPVgaXE8Qpe
uoOAqVLIsf6q+NwaOLPfbm4Fcplbe6Nvw+tIySjl4EP8f9sijIJdNPDVxce3OqYX
/vXb7NUF23eNW+adgww6OisSYWTLLV3vp8Q55iu4f2zZ3zx74EJ7w9Nc5O891Q9I
6lgxHNhkJ4D7hyVmOH1KQKh/fGRkionThLZ6ghk/FDp4biCRffPHPcK4diPk7lXv
fnmEwESxR+xkStnwx3aIMG1H/jb9LlfFhPDGyzYy8p78gBco4hlzTIGe8yKuxBdS
9aOBlWBRukF7aTHhk4s7O+xicZBKMFqIXvqNdUxDbLPDYMt7hq4zhF86ifESRbjo
sSqHMlG8gGEIipIUfyJMhM50zb/erJmIoFAv9zF5LegReqlKq6mHgYElmBRQC6Sz
p2PgA7nEQv839n5aINQe9Img9q6rxrB7EsEQxM6BM4LtR45z4cqyOsZxv5nEpdb1
O/1U5YAvC1RU0weI3YXwscj6584juFmiMI5A4ZVf6Ysqt1zDEfE2/BzQBEYjYHkI
nvy/1qtEiYQemFIMg5tzLKyoSKKaD4JviF2QGGCFHufhPxp97GyOT1snBHHNKPte
ncECcWeV0TV6duTB9EsZCE58coCoZiSH7DshOApQtdVmcTksmBJTv2vg8CxgoWSv
cwZNbl7antVno0mkuWy3fTlZggfI6BtJLucl4LEeyv89rUlLKVw2JTF+xknMly9/
2+ZOQ5chcV1aLhSlCA8SnXZIdifJ/8xvSxWsN761RhytA5o1F05MvkTVEEfeq2o7
kjJliSbUZbzZDAve3yNNJgPqUA6kKENRyUDYEPOoj+HVNdebBnuTseAq07J9XxbW
2lLHMcrDLqEF0lLzGr2UboQDUsXh3wlCtrlQBCPXo6cDgcJgmH08nY+lAhqlphws
DAMyE77jdk6BLiCsHgMwmS6p4Z2vFBvxtSi3AFXAiz7aIoT5/TNQPFhHGogCBqEf
70b3PeJ1Yaq3Zy3UR907+wyewNpMCNYEUvmrJQxv7Duug8boPxhPzUXCF50rUWS1
hyBwVjDDnDh7jK7n6/Jf+EEvFIeiZdgPUg64zkzDBNiMWsnV5cK0E833y0jAAyvh
b2hGj4TH1srjD3ldsJ1vnikcLqrxrcOCzYmSKhLXcvFnJ1iia87b5D1i0ZA4cyfV
sfNsDz6Yy5AicX8BxZxCEgQf4TqwKFgp0U54rY8o9mdKlxmrPoTputVBkREibqzL
dDLiFnKwZXM+3r2dwG1e3GajXLCZSVgCCsrqtHsF2nsyNmHjROLDmarMpwFEjnrR
NpDzG0HLREG9xmrxuehMcvxu4NCs4cWC/M0THOYD1bHzP+OOjd2QncXQ3aFx0KXs
IHI377CK6jPJ4bpqGGXJ30NgRqkG4BNIHnmDEtLIKnJofY82ebcgSbbKZkbQdBDE
tczGTFL6I6loU91vKjmDL/BxEzjkrlZf7qr/6firrPhNYn/55xLaUcIewI3hiO3b
eZ+yGZhL3wZMlRzPxNW1X4FrUHULqvkkChFmXIK0rgDp269G5xL/9KN5B8sS7KXH
b4clART+8tpYl2Do69Yym9FPOxzqVb4Ai/4hYDfz4WLWsLf4gR8ebVFTWJr8V1Ty
+5Emb67OMJvAlvCxEsy0xGIs/5DRIzlOmB+vXiboWsZEnYio3h1A20SjxyOsKlK/
xIP9P7b4CoHoaKrBU6uF/Ta7CL9p7IfXTXta2B5Z7pleL5U6grPKP9R8bqpapTKF
qS3BtvH3dUeTs/i92/vVojwYlLBCUpU4Rd7Cx2PCM9L+t5ENw2M+8+1GyYGXnivV
veFpqJyMzRjCRYE2WGrsfwYAOdbow9jaejrDFUXx3vCny8Rlbx3+VT7i9nyoB9JO
CnBkL88uzIO8M/eJHxvAWA21MgUaBFdriYi2twNF8DmImEAiRepA3qA4HKT057xv
XXxNsBUBbrfknbFm2QZLhCncWyU2La/0eJ8jga+SfDjY/d5/EXvY+WrsKjz9lZaZ
OUdWHlxSwultJzSt95ve5gbNpgHYgZfYRGhxhl+u/wPya285hkZW/0C86lt5I8/J
eAO1vYLaM4bHbFNO7MkQ8jD1HhZFfCFk7kAoWGTz285Ht/UVl/Z8HNBkLccuZW4t
KrNSWWM8o6Em2a2H1CPO4cwUVkUFz1aQZT5WZad2L6OZ4Z85ABoAE6VZGo0vK8sf
+G7QD4NYZNpkYXuwxa1u4q+O4nwRl0NbRxuQ+M9plWzzhdZuFddya6emVccgONWf
Zla5k1WdSDpNvxhKz99hlXd0dMDJ0eLfFHU3Fue+sPBzWOiCe5U+RVE3q31yJuIt
36tFSfKVuWwSCK1//vvpI0koECzEgf/akcCiPEtPmp+aBwjceANsOv0oTPecX2RY
cIeLsGZMeUhcMYOqjEiZdz013niLF+O/h4gThjcKbgx6alEhaQy5QTQUpj6Ba0HB
q9ghyUIrwgRpFR2JNbHt7NVmtDTyRjaLFGuQkIkAnCcY2BpQFlyp9PuiorREYbES
i6qJOORlnV0MazIDZjUIo6Pv1yy0VUQS70Fj76L9KqxZWk65EAvP/cBZqY3Gt1r1
XQYxR6kXhGcB2HDTtoSlJd1mBQeBQK45L0vp+u23c7zfKiYTyZKnZn5vInofC4P2
Fahq+Dz6RAF2UqyhkgZXTl92y7EGuf4QDF3TRYThrmBGRrrxqJf9ahzQytl3CNU+
g2Q7pOTWtna8SgeQIcdYZB038ly6ItyCp0TUnjinfZZFJPl1ty/6j+Id8tnXLGIO
8H708B/VP2zDAYMOLkE/AuLtkVLxjUe8xXoeNo4qo70cEkSi2J9SsGZ3W9QNLjSM
OhTUWUi/d0xPgwa07SoedbT68WlTqcrQphMWr5EWkrNIFyNHjdM0tHJ5IVd9Xezf
v3NzUoysrFWnCNlLQGbGzY+qfH5nXv1m6SVkD3l5HugPo17ht1cg6CcdvnXmlraO
iqYaTTmRAIGHbXeDMjh1J2A63tlQ2hXfSZ7iUfjBLq4uxGF4BHs4h9VlL3rMXtGe
k98qWtqcPK8oc0eAo/mX/PRTqisSAsYc1d77TvJUOx3KduGiw0VF8I1B9+J4lsPN
QoiCI/IkIJtHrKlcVz24ug9zzpaFab/biLsFMzeQ5w5RsN4bS4KynVUZTtmsomyd
9J5lne5hWB/te1xxhvIjWym+34N3tdfF4YSYrQXD8mpQCTzrCxAf9CfqZLmMPFRG
70aWI8b/NIgbi5qKek/AZUvJZJfO6wgcD3HroPBoKwgd9pBF3y5ukmfavsT5m3sp
QVxO97twBISZ5UZTFJgRKqyRXoSOylJfNa4VTisHfLmBCC7pZh0CCuoRs+41FEZt
QAiiXn2sAJ/6dPFtoLDxvXxzTPIr6WmwkteKMKPm7dyRz6zreOfvH7L4kE4PDa9p
Qyss/bEdWpGH1SXwRLkAgz252yHHGnB4C0zZLLgMhwkCpBCU4L4cN0CUSjvBeD2X
1cJ4O3qm4krXOl7NRuKv8CHrqJZGp3GCOJPu32xXProsynmHbtvvsUpMTux8ig2K
zEnIMdkd8brcirp1KgxBldOIMj+fel067o2v/CieTl9VD71aDEx4BZyS+ZD1hRM7
mTBxdrLrv22z0GhTngZQVNoL15f/dce5o7ViBK8xVGN7aHK3YMUI1dzbjLCWrHI5
SAyN/mU4WZQZabetZuUpN/SFD+rJ0Q5spxTgGehE7YkbIRyIfP35WBKhs2j3xT26
ey4+VfSaAH1+W1NVR1vjuokDezlkOuj1a2mY/EWDBxtJ7yNWiGn4RAMzVLJztA5d
DltJ1kMV3LhPo0KWoZmJBUSrP32a2NCgNeNM/EqoLIjbQQ02Mc4ai+fVAxEOwXd1
Qs0jUIxZ831NQWPRBpqRs2V+A2/lzgQEnJu2XNVnxcZPGil9caKFStpbicazMy5z
pS4Xiv3hBr0JdBXThe2QZ8dkOOxqmQpnqdc8huYEmJJ6b1QQu72eremZe+2zuWKj
gfW4R2TmN6txvyvRQVVPj6YbdFhGaQwR810pAWs+kbtSEqAooz439ycS1VzkI9H/
IuctJmdpF7qe3ngCbzpiqlIKAi3yFYhD/1BRt+XcJIkLlR4YuSH0+F3FCgEBapn7
3gO6eNZOVMmDXCLpt7Z1FAKajWcQ1tT1IhRxF3Ht/piQy5zq/YhwWfTmBueE4dvc
RPTKylp0UlfLzj5r8nq2IE3+oWSeiqcrVUikjtmIgCUe4hZRKGlKjd9m0aHORK9Q
zabfXsdnIwAKC+HNo4bb9VYJ+KLij+qFJDZfvkh3+QKMcFYaypIJkNH//npDwF+k
YZnWaxLyFN9zW5uvX30mKh7oOOSPPfwzh7V24+Tld15LCCoBCwl0wgyszSKhDjSI
EufYL8V9jl81lfT3PXNgBsxQkfq35GwEgJDHtrOlM2SaeALoMENQvTjCuG0Ueshs
6dRJgkxAD1vcS7RHq6YAihRubzz0LHE5pZUgX0F0EqfR/1QvVi1HKEOjKfR9WlLK
ZZPZ73FunfRm6mmZ0ey7EYHMl5dhuniB5yLWhqaZKi0P7vKCdHlRreFdL6mS/cVU
4z4T8OlJpFmSAJnaubC2JAp6jpZHfYQ9+oXqb0SrlNEuh5N+ru+hyy67+KrH0Rl7
mTzMdIzzMU9z5GFYQIhQDXE+LhLY5b3KQPqI/OLBHikpU0uHk9EWNZwqnr873Shh
E5ijRy/wUmW3O17ZYVe7A42j3msM7lFtQk1LDvuFAYeF6+fpIAaX64qUE+Ms6oCb
g+joOCWOj/ckLrtUoPHLgcUhD1VfH4ON78Dj9ZXtqNzmdb7KoCOyIyc0fUTnNPi6
JHb6WbEaccG1GRlFeq28fk6wLWCKKQfZ73e6CY5VU4Bv5vdW0xXu5K1szcIfsvkz
JRGz7KkcDj7PmgVk6OVZQ7Zccu+KdjQk5FH1bOCe9CapARGRWvGXk3vvpeDLYyg9
niqNAXbF9LonMzQfRToQQl492sNXiNpNuobDqLAkOqD1i4g7p6taMx+Xd36ASWEs
+O4A6zMucImJOyOOZp+o7eHade2M61PZP1M+UDIM0j6BBMWOLBk1zDnHeLiHIZu+
pqFyz7WhQEfHWfA/qeu5Yqpg5I46j7aiDmhED7mAXcpr8wzO0D9KOBD5r+SFYmZL
/7JlzRwVk89DQJYVPb4eSR33T1PLpsVo77p894ZZTIctjjw8fog2nqLcrkwfUhYj
wjCGC9p+8pbFisE47yXCu2KoYhRrt3Xc5fXujGp8qbb7PXcWLUKQyTAK7u8iaFPz
Qe89+PDUMvHuagZsWH9dA1t+kPnellGdX9hUwk26NqHIuCug4E6qWaepGvK3+iKC
HwOlueBCA2DjMJIlOFNXco9NtZbWszci0JamuvjMgTCeLY9dHQ7mdyVQVG7yX5UI
7lEGW6DOFDNGBDAOrmBBVlKiZzXzH3RW1MWYE0sqUiPHRdX8CzhEKUZ0P+H6/ZDZ
8t+WYAvKfiGzioXVSOEgkz27QhX14CF8jeZqy1qRlD9wOkp3zVPCsx097vJwyGle
ITvAjj6lUAtTm89ebaYM6tmBozp7uPvL1+6Pe4J+JYW4cQHgKIRm4x1HPKAI2oyt
TEx/hu/NAFEtAzFOmdXxs4r+TT0O/Jaod2RKwIfzFvfI10SO7N4DJLx0/oVr4qsM
1e4c3NW0NxtrHb4lMhSQiybS2w/8j1X4gFXcTYRca1RtjXZ85Ro0kOYxG87BVtk5
AOZMdeMrCxDIoCNRmf3Armij5UKCHZkwtQ2e5FczNbIDfRpsq+9ODGF6CUAYqvtK
1ni0HZDNTeKvLl7EkN9OR1O8Zn0go1LMWCUVx3Kvsbe4kNuy6wR7QVi1wHmE5o7q
SpRkAClORErGWh9wOypwyqQy4BaJdMZ8ZvWqejZWYoffDYZNZdXaqFWDvQPSDO1v
Vh2CO+lvLDY/JoroFjr5ld+M4h3HWhP8mkSCR3YzHcAjzop8c7aSFiK4/lmAv7Tg
CW8uFKu70gndVkZMcYNp8kB+OJayh4DP44i9ErqBn30H4HZcTjxcdtRahYWoxQVp
iZw6Dbw8JcGiv3QfKkylSUsf57mEXU3QmHxTNGEQ0cwvKAggaHun5z2PWFu1xWgp
8opC63BtzW1NRiwbzfJbd7IJKSN2JDMO0IU11u8TyVtJAvrJW9QZK4ohi2CvwtJf
Hz7KNCa+WFCEG4d1DoDLeLzmmF37FTOi49IT8R6ltHG8Zj4V7hxwN4uQ6Q5pJCyu
hxD61YHi4ZkgjO52jeqy0OiJWx4FqJ9AnPRDz+8+mukxkpSKhqlYYkWn2PepQ3VV
swQQVepzevg7MPom19LkDRZgIbwT+DXlOlW9bT5E/KJ6qn8kwfAUCekGjZRTxH5S
eTKUhuOzTbpLC6TbfTT+RkkOVy6u7GPF/y3gnZM8kyN+lOXINNTIFhjQTs6MVQwB
K5H959O8deeCVjUi5LTHrQPgm8uEW8WG2JXH5PNGYaZecmMdcBjC2SYnYagQ5kQ+
JCEfcasN1TT4W2+FFBOvdm8EwRLDg6vmsxflsQVUuyJ25R3FDxqavx4FqpV6zC0K
pfOEvTMpXbUaM8Ks50hGXvo5QHK3vZwQfJIi8vN3ce57/QrJBledRnXTS3YxTnQ2
hkRG5mpbsykxAOyuwvgWovN3HO9Qc3mABOYS1oSSihLS9NT7cES1CMmsRgoy0PXi
6TreXrWLZwGEiTv1jjet0O+tp/X51W0kLYQGEYpd6irBSqLtKuVmv3JJVJUwAvvw
1F3kGyPN4qX6BAGFy4ALVse8OxCupT1+l3OuBhX9fWjHIUUWpAxRXAoxx8SFeXpP
YEFJyGmBjrhUl4qbnQlPPQfGBN2ThC3YuMzo2LyR+BbKM/KpQIaXgB5qzbsAJrd4
WhFKg78rmqmSLVfE7OvgKVyrJD55FF1vkRtP++HSFHS7MZCyYLaANHZJUPHa2Cwb
sI5Mqk9P/8EddZQJj3ZwRvfwJtU0Ff5h02gCgkZXp8wmZAbfOqNECOOczIwu7sQS
jJM0GCInHmDt53qRlB9FR/Zh+L3vEDxhsbDkYMyvtxoSts+lzEuS8xKDMnvzLJPu
N7BjplQVzC3+LITNwCYNd8vN1GRZrKdNe7BAAOja3R8RokgERsVpcMkE4ZYIjhoj
7e4DVPz1c+9FErZDY+vZIS+8hkF39SFK68lmQe+3nZQxLVtWrC9LY4z3HytTvBYV
B6m/EEHacX3psINF5uEZ7rqNrWmOmNZjgFGP2kvH0zeXK2BQlqZTw1euTeYqKaR1
+BbpQMcHM8F+Q5xpQji8S1ILto6r8HmwridVI7cmCqxBmfeN06Mc2WKFPp0ZD7ge
kK3CAw5dEeaP0NjMCJJNkLbGBooTCqTsiuNE2ijQ8NaCC9pvdTY6j/q+BFSmrAjk
rVyDrZRFdA3kgjvR+pFNip+bfZ65277D3KSxOQGkPvkdy0mhCuEMX30K7DWyA/tc
lX5L5z3gxU01/2SGpmadXzPw9s2SbYbmxS1dtXmLGv7ePFnKwodBedCR2QkjjyV9
tjfeotxvggZLmAsyayBvKHY1veTQ/bQ9oeM+Jdj1xCSlJOc2sKJY9F5uOIoHYBs/
w5ekHS89F+u2qtsVHPrlAzIQySxoKZaooK8M6zuvj6LWULyySZnfvrVIF+j6+MbI
PemLxI4eIVUUKp+v5fTSDy0DqAlIWtyMzEOmfR/Efc1yahh1uddY5Dao/mXoRZbJ
DdzfrXjkZxSuuYO56hvJ6j4XvZj06D5hneLNHwSb4U2LdoZZrXKJVmygF0KCRk7Z
Ny1VRZwrt45qoddUEakjIY3JYOx/vZSH19RBtnr66ZY3Wzz5GdmV1GkKqxzfjZOK
6CFby7cyq6+O5QifZAh7LWfuH/HujiY/aVQbWUUqRfW8w28hs49SuwTjtrqLH5pc
jnrCKNizORdtOeSke8zN0K+i5XPj/e2wl9cDALGUyGcNSiNyzqlBhRTb3FebRz0T
Yij6uTZl1dZEzm83qeIMCJtDUkdb8ZJTiP1lXigdb169qJbtxiZauByIfwOGLg/7
hIH1t/ivnYwd063Cm0Q603BNUI4h5r21ByV4WleOal6Ver1+UCCliCcOeRBH/6Zr
i+Ip7YyGgeKVRptUphrC1x9cHze1cU7rhJOVJmpzvqTp3UELI9aCaaF1LshfRcbd
vqyz2K+lDjYAAO/gWmbSJdsOQsA8HsETpY6yphqKnl3YV49r9ZEQMfdPOgoYnIK3
Tr+z48UVp1Hkp0kzd2QlJn4VdkX+xPeknY1EdVjBTGIDd8VV+IxIfqLQIvKiz1Tb
JPb2WYeUtF9eMUS74o9mcpdPOCLMzsVsfSB8FV59aTxL84NDrdN5gBbm8zhO6RBt
2lB98TgHFgwMFeDF1KPFMgkRXKzU2h9t8hiH6W4LR1XyqWGcrrksT2RePm5YyjcT
YU4/7Rm/fSmeBKKDgnvQl5bakMOG0nhW6ajvGS12XXHwkRKq+RcA0dHbrznbK26t
MVFxHJPQp5y5tgqvsmIQ/Rov3Kuu1vaWcBtxObQarsEHEc5jy5kC5jDjCSlqRZcY
O1gn4dZuSd8RGQ+WCwXbiRjjJruI19ib7wd/EKUrOx3xCbwQy0us5B1z2fG9v2PG
n+FZVZgV4ESKabTGgSvmmY+ygHMlS8fReelFxDCfJUDIx8hgTpY180jc3OU1GSms
XiW1saH4mxYVfckyPNVcev+tjCXmBu7SRdX46fBN7fYmHoH0UhiD4MVlxmLLW525
/9PlrsjaMszh7aeAOySRw5RQfo7et+0PHy6MH2b+yoRZ1ed1ujwqtz24bxawV6Js
iwdIWm6qisWgI68ToRaEL7NWdGsxKKCEbDp4pOc8pPTmyV69vN3lMHUP2vAIlfSM
28MrWvna4u8xMOlpHq1mtQv0ERElwkJuvJhq+5ANI09Mp3lC1ADERqkFbyIjr7/7
IN3L7ajWy0cxP9oA6BPs9d6yeYYDtH6QUWXXs8UL8ZVEllEa/Uv0RnslUhv2ANw2
anWiN3DWdrBQzdmjp993hVsPJK4BvwYHkAJnbzwIPAjEaDH+HXH8bE2iqSHJHUju
Peku3yOePqC02ru72IwpDAdCKG+wbYKGmP9KIhe29ugLdeaNZ4imUAI/gRgVdchA
mGmhF4G0UHSXWMwgLLpIEFXJuu9vi+Pf5HYuribaqiv7pPBne+TKVUiLi8jo9k9d
oTwEDdAOP3lBvAo3UD1eVqc0MbZijLxKHAjdLMW2Cfr5TGoU3pm8Yv8mBg9QHBB1
LmRS8twDnut61NsWV/+uzYcg4ZNVwibPTyEVUPQXcp+hS4o2p9iNmlf7esvk05Vf
ZnIsw4yhpIy+TbINxkUASCQf7W04JyZAKQbNiCKNzUez8QdbTeo/imcH2w498l2C
3XaqRswME+sk491NJtrbE23a2Pf8XrkffPu4z3eUsGDNFvTeocuOeF47hYhp6Cyu
5pIHyNtEk53Edhr6F5+ge6ZYjGNlyZhifqz95lGzvGQMYreAEP/ACQJruTrbhMmu
PFbGAzCohSFyYfrSM8iPTaCXivrPBP0xo92/RTodYuFs3ZguOcjXpVjfWdOJQVu0
9ssuDQpaBb7X8jpI8u0XSXTwJrMWMQ+/BY6uf1QusUecpl6YFm+i3Ue3e1yvU2Oj
R9L27VKAJV6KFUZheSSK7cSTlNxNeCEII8zfhBuZBCZDPF/d+0/MoR/xqeahBKr1
ZDtMlxO+C5OxJA4PmRwpF6q59HH9v7jyAV7RXdtlK6DJHylFEPUMOeEt2bK+MNwF
AYfe2JekeyAqu6zT7LbK/JVghTkjUlu2D4vbcpfcNPRVpx6xIp/euft4hQA939eb
A59a+r7LA47fH6eyc/NeMDXBziYa/0lu4u9ZbGJ/WgE7g/O2MDBC2NXPJtBWRNMB
r/MbgAK/xe5k1kPsMvfU0Kvgbt6/GTyRu63LeAPIrR5VckLyjel5cKztGJaAWfgr
epoijdRIXdgGUrTcgfMTxMr2EJ+xOAfl+v+BgkdxHFMp0WaDgvUZMvEyogx2jQUV
5nu4Gyzzp5bnVZrPO9eVL09dmqfOpNdfoD8v0at5ILsRVGmPXy7+2LDeyPqydeei
VWZKiKT5aLFN5zOg63xhO4/pvAUike/U8g8UEaX1jYkT/H/60OTex4TH74lvnMDu
ibJRBZ5USf+JUUcD1f5QIiFSzhV5s+ynt/8j4ORqcBXXekkbUW7z8Qmgq26qJroT
bQaP2qpx4lcXWJvfRWEHYE7SvXLUjmeFRAnbeyTPibG6J/lN5mMobzNNrkSOKAWN
HOGZRzRavdKDN22C20ptSvdShzPYnxhdf0dHpdqhgdCIvRy7sH0Y9YnDKuEBcZSc
74ah0ocSp1DPAY/mqPIA/PqQWnbs6wz82Qc5ojgSTu1guqArc5eRnpfQcR7zHVQM
x58a225MQDUFjGdh0hn/nbUswoC4taO4v1WCQLva3cv8GNNU6F6p/PLDMgRt0w7F
3yxhyFWuFhkFcTAP9zJyzHc6A4+g/ZHp4vW5qPci1CUB6CRps+dpfqVKrIfypNkK
4fX7HTnhMwuW5dcBQ2pXKOIPgnJI89bliVoMA9kiuayiYLOosC9tb9xrCJvhX4lZ
tPyL2fQJ78uQruetbtE+KteyJWih9psHc3L20CT85ZrnaEHqdZC6djpZ+5pecbGv
2tPyktFMcFPOfRctybeoDaCGOl1+jvw6JGLz2zDabFUe+t+MCfIkDch3tsiPEpPe
GX5+gY3601XgXoIG8okhleX1QkVS7dU0Adas4cT3BJ8SAbJsCGmBS5sA+h38SNzN
h6y5+5nA4aCagrJHii2+FL7Hl1HjU11iNMjvR8zzvWZPJtk456vKyiE35Qz8it8A
D87xEztYl4wFrZshZSqrClMJ8QGub+fSNVSWgzPj5h+eOSKXBWUPoXWLyjgoEQAC
btLc1quSjAm8JkpgYYAVRoDdf+aYt6qyQx4WYXB5LkNDTs2JA9IMWA7lGXljrJ0z
0yQRkrcXojbFI8k+qPhim62WOjtPVPjxCfnfITZPhiiUC3DbDRHEHguvncSaWcu8
aUONdEeIajCvn4Wbd7ixRjjPwtEqAH0fuC9tLZZD7mwAA5ZVOxhAmwDftoEdng7w
t9/PGGWEvsWvK3hqKR3U8Ansic00o1LJ21rVY1LInCsbMXe8pwooEEmAmfuVHfsf
+9e9tzyZ9j7nXoF07/c5eKLXcKC3Dfi3ItpfQf85WB0r7expLWenSD1zEVePbGor
+1J7e+ETnCZR8Cf8ufekzCH0CiXJ08+Xy46JsZhAUllS2hec0Ol5Setqz70S/rw6
MtGRtkD7XXmGgLQXR4rlxDMoYCZeni0k3mxTzRScBu+UjSJLFgdwAa21arCpmpTt
9sOkHOBw5WsD5aoBMp9Hi5tzVpPBU2bQj2Ll2glCYKI347D7t/64TePdXXNMdWBA
+JEPpsEu67sr3nE7+RGYM283Vi0mockBG8va0I2kj0FQUb4c/cGKuEceQN3nM9/T
1yG7mYEZkj2HgH1ytHUy8/DGOMNpQWe0hwsQqny+tQJNpEYrJn+SdhE/5zdCzfDU
Mq7INC0qGX1Aq6jn6ksb5b6hT2L985C7Myuo+mbBVVX3voC7l5Vu2E5GTf/X/1Au
u8GaEX+zN3mkP39JLJCibClge2R1YSMz38hPWRLhtJQYlrXtP1x48gsK6FRRN2yW
92UkSxaUP7jTAHNXiiJ4ryw10YEYkh5cpQVwOo9HLTGnwlF9ad5nwJUS1Blj45Wi
37Ntv4T4+nfBkqwDgLtDafsMyz1f/cqR7bJRfzqmegTgtrRfs3+og5CSEeGWg9wK
9wSw6dZTxBvpCucO7f9QAXOtCG6T3OFLTsWk+wSfehenIeQpzqywQpHIr5aYrAaN
0ieYg4kQ7iNcwb8msL/X/MwCDS9thLVn5RY/Z+Yo9LNw67DYHczwSTWyOs7AypX1
qNjaTuGRm23JuApPY5gBgzgUIxVW1hEFQc0shBg5VnvowyaIrSD8HM1njnEjJrMw
I75zcNx11UVUB//fSN9z9BUHZkBpqfQVuoh5At+oKjjJyXp+abOADamugbEUmXs3
ml7kkvTOH/dErg93vVDa/FqyJAZ8FnWKhHRE2W4Ek9MnK5tsExvpe7CWLv+QCtWe
n8xnxUdKcFe7XFq8BZhmN5JJReCwzPTWg5FZqzT54IQNahK4ggUbbTHEEynTka+v
2HTq9XPVOdIuZ8iwVP3VF6UaeEr/SRJ/N/2hutuJYPDiD0IJOYc6StbNec6h9/h+
blYn4ty02XOUUKucX1NjfS3ItGmh/1qIbfrINp60mmQpDAKnRRarkHl1CZSd5tDe
BMaAfcYgyKnH71DbPVpJ72wE9UiAwOyBZ417YAwND04Bp8QIh7r6eJ5zw6ULKvbA
8QLhxwItYW1iAKGtkasDrMZHwni3SkTj31vA2sGqLVFeUKW7onziku9o7qRfLIjv
5FdA1V4sZUSibCjQwq59vafM2OKrNIYoiw0UFCDxTu+dWYB2VykozOCpGjAEE8dS
oyvx97yNYStb7Sd16Ig+5ZpM78qkitSXsnSiB1RJCJYHHe9DWMjjoMWf+Ql13QM7
CHwltw+RM/7T7WY4ww8anj/UCTdXFperT9zen8JJjZpk/WbGs5EYtupuNW5X9VP1
RZO9NED2talDrlOSztd9v8TyiGT2b/UOwhVFpKkgtjFNT/h62G5NwFtrvfUJpMTS
d113roiCpbCIJU/V2klkCUKDwBfzKw46TQ3UOOl6vGHHYLZo6048pJDFCyOvNHCd
F15cCNLczFq/SVT9EwWSTJpby9IqQA/iCcs2iXcJ8qGVWRhxs/DemnouQv5Wh04E
p+dv2xXy6kvAYiIkpvrSphQOoE/qe228yNZxiqXuj6malCOJQG395NQ9Me6517R8
02gCYmvrbOvMZ9U+XxRXRNlxXTGECZIAtFRhbooA3pSFWApKMJA47MxTU/On5/ad
+rJ0Qf5Oq6cPmY0AJkQuJnZVtG1bX3RuvNDrTjdzX42TUeu0WujYLEE8igNgdrXV
V6GQaG562GiVYFmbiL/r+dNcofJUNry0opBxX8f5uRqs9GeNRxLLnOyzPewVTRkN
DbFBymVlIX/3DFkGMI44Wh0BnrDOkTOhY6mvUOxZcokJ3XB0t11h/gV54NqSZ0+G
G70JgUURnR2FltXMEejyFMCeVVF1yGljRvtEv5kHgM6uMKVxrwqiQDhMHYGKd5Th
OPigK6nipPuKWeAC1FduucGh6LDXVQNUCaZpW/FETEcAWXhMlsfFFa1LyjtLBYe8
znqLv1iJyaA9Ofbj8KtityNWsmq8hBPYfTWp5XuWZASv1yxBRLCMacjekUpzghhn
9wd1fuwJWNLF03hAvdumBnrCX1nCIVa9yHz6fYpo7rpGIgYgaqjZXRkXK4DtPXWy
EOk2r3adQ4EEtT/SKBcgrBnXE70xEWP3tuNIauEhH+fy8QIfwz6Fbp+nucrnr3P0
OIoQUArvwlUPvNOxIjvgtBTtcU7KTIY05MLMBdN97ciYTcSXMcbLbsaAU5lCEYkq
8bcQ1+sacUX+Il/+00buFbTSvF0E22e1XRdfP4BKidaPW9ONCeGFT+pcNXd97bZV
/mWdgkjMFkQOzQIRFbfnfqkKWD5B/WSmP/dtHXgn5AUIQ5Vo14RtyqSh0HRVnW3L
AYFqBIo/6XDFPU0c4udLEnNaRxzdnREID8Tq7fNDQn8bkjM0Dk3A1zE0L+0Gnyya
aRuUT+8ycs2ikhIxlwI5kFd6RYBr7oBjmqq/V/WzryuaTm/37BoA4GQic/jol8iR
/qVUsJ3SXakKgulPlWZMv9IUoLSfgnaRyfn2+UznaI9CtFs+AUTKT6uICByRtTb/
Jb7n190rTPNEchye1NJm+5wRQW3DE8OyFGa2AKqRaABWSD3imp4sRGUiXJkaCrm2
FIATwYivvaaPIHAIIgNwYELwua6uGL/yqWnGtjwhVGzngG/w0djikTGoreHzXQ5n
qSn/6xDa9gdrcW6D/mOLmeSWgTgx1dzSVxGEfKSB/05TomBUD+bwzfEhPluQIlan
RB9FKOrvU2BpOsECpcHoYf7nQKnq7gW1TFOGHkzaqv3yKh5AX7zajJu2jhZvM3R0
3NEy8TlNwVviJ0SqEYmSRQrHt6myFFACSrhXOCOggYRbm67kIILLvqkA29KY1vNz
Nupoa6IMAzoFAG+TGYBG2qoBWFqy8sadLKDg8l3VyP4X5LzvJWqN1TK5SJftELOE
PVm0bxHBd/wC33D5ZTkgfaybjHHiHpIDykNMt2JekUXvaBP1La5tuoSwOLA1vfCh
GZgMO3i7Mac6XnoUCqY5rr/Jry8EXpLB7YGUJVMO0rEneO9/5IH66xn/+qSKEJ9m
ietW8R/6gSvNSToK3QJRav3NomNOgtkuL0V7cUNHVYU2nxrbU0bOzEx4T7SpEQVe
yNVBp6SfNwKLOp70Bs0BpG1Yy8R6C3HzOdB38Ni9a5nEvrJ6eihtV0URJplcvfYp
vpRxfcQcvImirzxHyqzxmBIV/NRzxjGOXl853abYCDB+mF5/sWCnX4eLWta8l3By
5j3h73N8QAivrKJuVEsbvCHVixhfLyKn8l7BX5Wm1k+LZNk6sNse18Z6xXvc7ixX
+rTDtuoLVfTJpgJPAK9uur1jwW9tkBeZFWbeP6se27hRBIhnRjhKmxHwRJPu05s+
PahL57ldvL9EEsd4jIb+S2SVlXMMsRewomSgVzN2icg1g0k3S2a26Cd4xbLl74DA
dQbhzsQyHLRZo1FroocyrelVsKyHNMtfVVWLtrbey6F4Ya2FHbu3IKKAH1OJwx/O
gqAPOCQprlsQ1jCNeFjbXYQCUKs7QKxZHqgcXPRpku472hj38sC6WIaDmUBza2W0
2LYb3RKurspFkUh/hnovkFXctj2WECtDIatKk7kqIyMe0o3fJvqq1d/FntCrKV3H
CpMdq4a9pm5nczTRVKLsbYakeR2wLVscgVUR+DplLE92tt7igwcWtXTd6wiryG9K
xdm5274NvYPVBiolEFt/PGl0jT/P9hqCa53us4jzWgF2vlHPrS7k5QIk8ebPpkSN
gmkmq1S4FWdffGTRAIM3061rZs4lG+PxusR3PF570CNV1VDiCXaT2Ca15J6fDcsZ
Nfg5ukfmfMY0Zwf3tEO9VAsaqVVmPJAvxYAIVht0w0UlP1ncOveKvflNJqNMKuJN
HfWOsQJApdYltjQlRKlOPz9vcmh+4OEVcvyRI5wGGm50GnGuHYV2rNDgngy0Ne+F
9aOrHuKichvwm6m5yOymkyskazokYp7eHglvqhtBEA15NnG+IWwgP0fWlGPXZUUH
LlpRFdSw7ZLgH+gVLZwYqKp5d7REhQNKvB0fik+kSMf0MbhHgXpov0DFD/y8qoof
WNUnrog1xfri7MhJwyTnhUPooSEJtVz6TxUoCp10beTbnGnjM/tUMo99fZBCrQ6S
HwBg9HgzIN/CRhrIAt1lDu3hYmCT8AFA/F99B7NZUzBadah/kLPSV33B7ZRtK6JU
ptGduOBRzb1aNvXX3ebv8lA3nuVzdxRE9JCLGo0OOPo79j1OzeRczRyeiKgS9gti
9+eKFPAn/3/swbP/p/SwAyjlQdks0nJEgsynH8RdGlErQoTlPDn7IhAc0w8ZGTJe
XLWu2Ki31a96MyyynDRhei7Gc7pGfHd5hCztKHooj4iL9hPNoJ/iepnoGUnytICJ
vNKTSO31H3fnnbJboAvisjqn1LYZO1LyqdZ6sSpqwnzuENZKyQ+nL5KmkQQ9Rz85
a/B55ojRWCsZ58zbQMSClaaWr7tlXsALO+c2IqkhIt9SmjsXJIqC+yKou56Q+Dw5
qAF8I1BtvOLOD7un94ciur20wU5uhfrp7hYe696lK2ekn7RADIoyKWpInDfjIjQM
xTBUeXMs0lO5qeihvRxrCO4JKusravNQ028hrBoY2CeI8ji/eNthoaVd9yNB38OY
6LFi1rf0l2dkFIAeWggJKVDpve8IJKlZM1J2A9PfV27NXUYmdz9/uF9EvKHBBf//
bw8HrdEDI+wHAPWKz++ioSyLKsH0KUFUrnQ1Q9waUBiWrm6TD51i/wLOmof00nRK
cPZSWL3CH8JKG3bnVUxaLc3WEzC+6WIzm5ytPDwFVygBTQUhjwNEf2/7PhlaJU+K
Nt661zi1JO94Eif/NBCse4k1gTYFlf+UsA8VdbnqNlCTkS9gLn0uRWaamQ5XgEoj
W0dyLUPcU+PMvmzur5Pu+mTXzJqF1eGXavmGQXD3ETtjdBSlfrW6VBP/cZBNO3CF
gpwgIqyeqr5rqZMydNFIpEodmMQBBprnQ/zr7ELKAaZuA8F3C5Ts1KWPjgvGxC+3
RlujmirEBkJC2seTCS7jZG46clEKv65lHlVDpJZbu2oyhv7jdl0qd2C/7StBSyJj
V9KPMweFdkQTMDvxJTYkAcB9ACbhOYKGpEVxxwUUopl5WUDj7TUKtlvZVeZTVjtE
tb/oCA5a8iXqnYjPd2CoyqCN7qhzb7aYopbQTNPOm62Q/DP7ShoUA/Rv2fmCtlLp
KKGIxw6r1o7pXcUMPZUvHgY1wGlSYCZHYLelvXFgXyjSvy1CWIzG53NCsooxsxva
ig3BeJ1xFsEp0fzfSIZwtZCwnSUnxLMQvxfbVJltH6ZBvNVFoTrMidACunpeFtcZ
GWs49ntEnoIuOh/pYZDYF5X4Ab2/9xVoZg3OuvYHmFkJWYiYxj2cbHB5XJjgVigv
/U8RIiZCrKDH79b336YYEOxrUWQCctKWFc+q0MX8udDVWQYMxqNjJFq5bnlJdvq/
Ptch9EsxmMFnig1nlK7gB06sIZkm9ALKi2y2ycrv7txRp2XRJ9XBmOwCofP13obI
H+tJo3GAtlCX8FBYxIzJ7sW6JrBFX63rwNqeP8Lsx9hnhk+VV+dgZoCy7TkDwSwj
pVBIjHaKtQ1GkQ10sKuMVJLSVKtkIzPvnkJ3gHCi6G1VgEh4ohp3nXW/9b/A5JOP
CxkE5Em6solM7JZUD0egMNnR1r8YV0BOgpWybyCqFLcEpbbKzCd3Di0DcULFkQ89
KCJ+gt4XXwIuL3u1NW+H3DNdKFAb16ZNlRsKmMwUd6w7zxnmJliyC8/7bucXQNl9
4duglPuVMDvnwuKbthcDLWFrKLuHslIGKhppQ2cISFpWRuwQ+HpI81FkgCKGgfjI
p8EkHb0w0mahH7pbvHc7kmflfGcX/SC1WNCtIUoc8wt8892UvKYiDN7vDcAAGKZZ
5FPnucDvBjMNsphb6zYMz2ValCHVYYaPowBWw6LcPAbIPzyCtB3Seryle2bZs9BW
BZIBxe72PffCdSXbNXcVcy9iCGdM3p7QjT32P8oBF6wWBlvAbPRNHo8C5BWD6np1
1BUQNE6H3b+2zxGf+meG3NKnLN0cS4OjydOrHLB4hihwXsXjMCtbNQRo5tEnrypo
dynWuSPU271WH4l6BAU5UvS0liwvlmQwt/l7fOvCuvY7XeDmHsCTxOeDI9AXP4+2
gA63AftNjQ4R6R94hL7WaShjmBqOIssI9dlIhEcpxmaLxm+/IOJq0DCuPwPtKwHG
R3sVy2+yxzRHXCN1no7NCIDh7rzvnNsb2g7p8S++icZfWhdYG+x57A2VTsluYxml
E9pfEYdEXtEjMq3A26iFTqf33kXzRm0P0Azy1X2Jn3V0arjFj8ijqahEDokfGqzK
/jSSIQPQmaJvPEaDgv0jOVyW5IeqmcSRsrHz9widpJcW1pvi4czN9/eb5dTqqA+5
ecIZNnbSsX75CdEH1FTue2XTTCAj/6xuyvzDWtVLTHBx5+Vj6wgpWU9ZNcdmEKgg
EbQBLIm4TsDnlbZ4qoVmr3ckQslYB7CjTvL8MeH0Bd7IxXcLGx0tH9aPUQ//N41T
LKgMvrNUyIcOOSvfVo+rxJLnsbcREm6orcru8Urt9dW2Q/73pdhO1PA4ge/AIjPJ
CmMpOKNGYnHDBC4P/i5RA8CcJHH5OXsu2M3eMVbuJ2SNL4ofWbFipL7+9voA4Ds5
Ulns5gzpL7LI//vzXAzty24XYHn9QN1Zvo1gvmsjCVpTh70xwi2i/j78vCTm/Y72
YNhM1KdIrp/S+2RLsADPgSTpaWzOQtPcfu2lEOnrQKknOy/mm3SgKibBhZ4oyCcD
2XOH7/3xEoTvOUQYU1NhPSND7XWdUpf13m+6w9+6Yr5zMH9TI1vI7zABnA2nXW+b
hwnPR6j6xS/ZPbJofbZqNJdkUvIDbY5uA/COmuPiG03uTJby+ZkxewQokOMgn++z
NhdaVXLnqWX8HR6uUitsFqDuXz3ne/U7G603Saxft5UQlIpbUka3Xp9ENgFs+oBj
beaUKLUHtzW3V+C0RjWha/W7bspwO60NvBUQPEhqTnIPjoaevQEnZQ4lrfMXtqWU
hgm1Bj+NA0tcoPmY/4ldLh8OAZnH+NTMnxZp1en8ESPCHrv+JUUTV1GqysGImRay
PjbuuqpTeruHUbDDRAM0LFQJmSSfVh1Nw8QsO/YFhG3BmbkEad7kXZkPjjAMxkxU
Xiz83FsaaJjCS1weWrQwxAKLNDgCfh/9G+Nr9WbKZPjMCpJG9EvaABfywfLMyxIZ
wOdO3nofQVbRpzOHqaC56LERJT8YK6Am4DzwA5uszyT2IjB2YCT3mMFiMyLd0On6
XYK63I+iLEAI67gmOwyvZ6BScTruXYKaeiJ/C39DHCyqoYqbA+cXtklMUOR07mss
fVscyAQotwk0oZPAYXV/nNX+2LXlXNTnMsM2k7nS7zqtHaHj2604aPKAmjZeeWKy
Zf2O8QeN3D/sJ4I69bkXVh8QZg/X9QZkd1FLalgwgkrf0QRuIE9PiN4UC7cGHXhR
6Xh/t43af+MIndHmeX65P2trhalf61laUc1HXnxsrfbmcwUcJg4EhJW1jsF+MBE8
dUU4RCc6bGB06/T/b7b1RQ292arxRqJzicBJ3GbRnfVzZaH2n1Vnq9A3co8rBUJj
rp9gb2nlN4GeYbWUeQiOiJzYKHXApFEKdhOM/VHIM56lXcq5LcnDx60u2YdP+xCr
xWC9EqBsSpckPMYJNcmPd9yyCuriM7fPLnTM+KEX0+PxwctosoLcQISJdLRY4eM+
hkKiouc23bDfoG8rcLYmaigMdDw7kGDC8lkSuPCmc3cW/XC7Hl8AkuwmQPIS7aBG
9q9AEZ3Om7nSDJTAPz1Pvy25dae5fBJBfReqWA7QixEBQpWkOHFw4Xyso2k3ROx2
eNxBhkrvtatnZGyLpE23kesFkzJ3iLQpanmwVj2bjbn0EINx8X4S6jv0RFsxDr+/
yVa5yBnbtIIXyC7njFB96jknUm/nrG00Z6IVkt4+wXl/FGGLnHUzORZ17FN4FU5Q
zTZRx5OvAMkKjGCzXbAZGhwGeNcaxNL2nRWH+qU4a4A7Xg0rYj12ByLz1dj8T/Hl
YtrmvdE7nLANCBP7ic2zEW/DX8j2EgbDPKaDW2nr86x+Hc7t+COFN4Pko8Lfa4KN
neEFtMfyrf1yTEUR4IdMdJgeefh3Y9qs17OXsf4qtnsaSwM+XLPCBB5VWT5tAimP
Sf7po8akJi0x6kfMjZDWvFUvLYTIJde3J3cTgbjpkW9VZ9pEmllz6V8Fi9gmGltk
RJQoPt4TS8EPzB7m/WBDD+/Kz/ngOwZWzIzbwm15tw9EzAu1MFaizKpXVgdKD4hs
3KTJTPyIRjoQINTKJ1h2Uvtwbo8z+yzMT1g50FaSlXV/6tWJjdbnbqyThXZjH7lT
pu0Y7QWWrqBoXc3+g1X2qmHvjYouAZXD2F4ZsKtKwGGSob8CV4mRYbQDcm2gam9D
C5p3JLR4Bjx8vabnjRK5bXTAayNYPu3PkkS2/CZiI2oxUXqifK7EdlnhoZ4WbUBE
/LqZC9efAkB7zhTsLffwuyNjCm9Kmt/ta0c8aBUwmUHmZzI0Hx6z4Z8jvGi9TjaH
F7pE02TXn/HAaJCqc3jdcwQmY2hnT61pyzU+VDcBA3bnFbgYQrJ//X/jmVnnY11j
stW9fCI7VheI/QGI0RRoHTAqU2ATDjnfhup4HvNZ4lPXTSwXzq4ps6TcLwAoyYSr
52cUgARHBXYotohWc66R8Whk61WlmWZdHail64IFP0HUPSH3QBBlUbB5ciCQ9UZT
BVDxxsxII+SL3grMjJGvcT+hus1yPzqt3f5xdhXTd/ni0u6BiNn5xsUGyU7+X1Vi
zEMxNuohVyXsTgiocRvxJmaXV+ryOvA/dvj4rXaERO4JR/IBEi+SG6cNgyT2CG09
3sPhJORoYkubqh35GpQPkK/Vkor13vDuV+NACrzo+fjQwkswQJVGjh4isaMgNzsH
8KGzx3obJE3/BeIvj+YRi8JlGq9/3HZ/ExxJHH99GK8U1Tx1qtG6spoSnNeALNRW
3EQi3cqCdQ1em39biuBj1BhMR2h+Ryaaa/XaPekIMoyx6QgRgI0CnPf5ygOBlPuh
ZN4DOrE3o0E68/RjWXVcj5wXg/0AfMfKWVkxS/5WLm08AnGErBfu2HaMYPXuq5hn
swGwJKvLvavaRUUXQF5n3Lyyvfm+JK40lS70IB/N/CwIslPriTgl8+pqd7zGAhsS
AOD97XpnobTOoAw5XDIymuRM77eyi67t5EniX1evD2ivVsvaZGMkUZf2QiRzRGpz
tNfkGS5Mm7cCEI+6vt4jOy8eB9w1b0ybZye+yX9ZQyVqLWq2xm1S8AmAyc3ZPCRA
kqMLWZiuhXauckQ8ZeU2pZ3NMGl35NPKBqB3tIiMJQ1lmZgbJE3zZ+co7MY//t69
0rWDkkIPvrSMVIVYOVEDKtMFyCJUY0hr6FCaBbVjP5s5eZDPbYj9RiUazU5QndkZ
/S0iK8DWpVEd5thX02mLNIBLLdm4URd0NWoEDrvZb7k2dhZ8f0oqzKHNA0RT6vGU
FByROeYQrzhNm8tADJRELrqkJUoCjqmtUndyfv3kdpbjXJ5SpT/XsZR0KjBKkym6
RY04ZTGWAD/lFW7/PZsTWLhTPm6cibVe8nbUzPHEBc48FhBAYFNNYfNNbX2GQ7zx
7TWLdA+B8sIvFyMScnDVfXTvACGDg3KzF6vxsbu22IzxGXsHzpr1gKBPJmmIFO1E
tB9Ur32pqNjZiHdw0Q5IOsKyY8RqKJvcFch4qqPfAIIWIcHSd2+a4DEKnHB4ZsvC
dO8pkJUvvvN6HdOteC8AeFBKVIoqZes5+A6HKRYSqsHf300v4yKjDtVkQx9ieASu
lo4bvv5QlGNW9Zmr0yR2ihyCmC6T46w+VU/+OGeplaimTexPKDLIKRtWM/LR4pjF
zLpBQ9FxUrIR/hqRtd6/VnIQKEWpTQxNhARXWe1KZ4YlJeQ6aOijbQb1QLFjaJoT
LS+SqFAfrQgq3juDhzuq4RlJIbnPwcHDxA86+jjSU38zx8ccNXXxKGh2sC17y8fL
U7nYViiQrdABSkQgZDVOfl0hjCTNk2tNFGdT0pTj7jVw7gEK3DJJIFlkO33fPhKT
eh0lD+IOOvODoig8OGrhPtxp/0kpMkFPxX5PUtt1mzTGieWAl9//x4hTz/a9Ek8U
DIZWjw+q11yqe9kg0tmqxu17WTKwe9WXKA7otgzcMzkROEIma4WJUau1alIqKl82
QVCLTyG4gApdzL6qmQl1KjvAla3tcQgHJJWeyuryGvdx5LG64cGLETYlrABhqBdk
zvRHqjK7Wfo1YR+7xBtgQwuIV48mfRryDVcP0ipO0HUM7HsViFNmeiMBrGQGuaWv
XlixLZ7xcML5jlSG35zv34Y07sdTDeEdkNgSCKS8irWO7eRZKX00rgMY6GhHlmQz
IxBcnbn5YNY0FSnDqCCK+luEuCLrxQFTFVa2D3E45ryiV590IuGUR0LUOnvLTA3w
WYVUVI1XS/lYmrN0S66AuwdJcaasz+9dx1th4JmQeEwKPGI2Zr4PUF1LRcdAVdCv
tq2FAsBm6/HD8322EbPN6FcxDD5QCcS/R8jRzYYoYELWSKRnJXtlRSLLXx92Bx4z
RCPe5oqecwZUJh5ZoGPgWEO6hrMDwxge504mSGYlkmYs5LV3XRcAVlAxZA0valYm
6PPxnChsPx1vMdMdTrotfwL0rDyQsh28fK5Hg+oOiCMFzwSHzUiwDkPYqSNb4DGi
VL+p3V3z8se+ynH32YCuSyHCItSh2XE4WRs0odYQEzLWM11OKe9iZthJnBG1Ph7k
VVOjOLNmaTfIXLPE6sDsnxENsFxguI9ZhvDE9V2+ZXSKtKaWCAxi5qsTxkKoNfgE
XcFrxgeb8FCtKF9uOjQFPL6A5JVR9KLIGgwz9NzcpO/KxaMhnxe3bEOzMUSxvgMv
NcY8VLBXpPZCGecCZwRrfa0GRhHv6SQzXxuYF3XFdyeiluOoHbRQ8+uvvszQXvXz
y8HxGaZniTDdcpQacBULCViaf3e5Bmmn6bLcQ4VlgwORtt4oHWOXP9LkUmpG4rlm
2EsIrnEdvu7GJh7k4sI5Y6PyAcGNs0XwaMkGqOaA2Wh/T8h+3U9nA0wjLUitYbcT
xLYnd7OXookPp1SPvgn7eEeeJxSZxNBT+gXFe2ZS9qUDHpnBbZ/Md2oISvYuT9fs
et9+D4Z9YP1cM828UfM+1PrL6FX7MJZ6sJXXVMmizyP3Mp2BlHQWVqi3m1vunrKc
xi9gaeOhl+VHJj4o20A8Eba1FTzDI8Bb6/Zi7zYtZ7+b4Hlaz+AC/utt02w5XEV1
BCaj9urh6sThWlKzCrheaU5hO1Li5t1GQJ0ysiN8fXBrl0xLPyyylQR9/vHrCCc4
g2fxS2GeVbRGUNllUsirFpFmgwBr8dxw0mCL6y2BkSjArucjHXwHwHr71PrhnACT
WkNKWt+hOk4ISMyXW+35ZNkYLzDm9A4t4jMDvHaB3mX3u/uJpOM9bKBJgARHSKpX
prp2fUbydIMXOKzYkDjk0VX081+i20xmenc98s8Ajzs2qKfOZ7RWti95WVKgML/b
UcDXv3jMhRApxcCN+bTF83ccBrYDr3+7ByOrW1SwS2gbDHeZyfumcDwVv7Jz3ScX
FKOyH3axGxNGBD4g+tBINVwVmKjervDBv2veWNyc8NNkAL9G03uww1uUGHiBAnkN
0C781VRZ6TuuYstKjKUjYmLk/6q58KRUZ2T+F902qRpx3txgcnde37T24c8lzzfy
skg2f27dceCr5ZqoZWbedYt3smZkXMSx1s+vk2X/uTbHHGyuCAYHsG+B+i37mPgh
VzOMHlKIjDwQOSXGfaF+ox+LHvNzR0p5Q0HPFTb21kk6WJxphwGxvsCqA3IwnOl4
RIS51czW8JO8RUI13z5HWsUX2Zdac2Frt8ZzlS6rHBkf4RHfDntSzP7N5aLqUExL
GlJl5Fpb6KdHtD94nd2y4Iv6OTJOCX+S/Y6TAPlmmaiOUlM4QibtD0dJRCePiG4H
gDpRdL789n2vxUU0QWakndZQ1JRgqQl7No32cCwpKNVZ+QIKlPKDcMvsykH8texg
nNju9IfXos0HVFCVwujpXSM7uqT0zO+tDXsvyUtmjbp3CHH0u8Qcvxh1P6/2b2gr
DxVEyOWjeH+Bh9RQVkbVlAa9yJdRxkiajWq3lyy9NAsFMBEpvm1PJAxxlnNBwBNL
u+RYJvEuW/XiXXuNzmo9ilGuNYO+Fvf0LPJ9TKKwx28O0xI/vm35i6dvBeERX8mL
Dc+vdLWlrmsKWp/emyaGn7muluTDTO9sAmUrOx7ZWFF9W7dpgnWTEPk7RNn4wwxq
KOpNn37funF8n5iwH0yc2V3VF7oNoTsV54cR4wPgauypNNXQOG+EyWF0vhV7gaQq
NVwoU+zCtL1GH+GKGuZQSdiN1c9Y1Pr0DthDhS05FYqeNVz9lqX7HEqPfRqXIL4s
IFTdLUvFR906pmhTEw54VztNOyoHICM/7GV9KWwZuMmT3dtlN5jCCQECA1d8Kq58
GRaMQ9ynM/njY/4p768uaXxYIEUNYwY280q+wMGJminn9tBpzEZUcHav/L5r6DqD
ZjD4MztCgphmD5HljD+oB66iGNjNvb1HLkSFx1PvyVTtieWzfK+BNe4hzchvJggH
TfRe/NF4I/l6mI05o+wkHtUAKW/iRVIw+Thz0MW5iLCUgWNiHxbGhUDwHUlV7EPC
qWnf4cQFa3L2RCvgRyEjTrU+ttK7bVYaQ1bgkvW8PENekgv6eaN86tyL0UW/5jYO
uuT5joCrYl/d55f1UffC/TV4tiUirc9pKj2sp+LBq5nw94WHJkATcG9JFkIyvhxt
cna3f4MYr1UwaRR4bAR6BheY2wD2eSVGcxwS+nKbkYyzgMwKf+/a7eK5tdpx/dv2
vNFfpvmGc3iG0AVo+WWYSNgQZQE52rapFUn0nb9SYf/LxNKtP0h0daOcXrgxRihL
ShhtBXz342fGZT+fCfyG1vnwXhIfQPO91H9JJBKwgAhHTM6g0aYcA1Q8m2Qq5rxb
FnD/sbr8YKcgfItPB7QaE7pTHcmEliFvpi217xqN8/r47xLTiKdL7HWjvKqRjug2
pEuG5mPX2/m4xZwm3PaNaIqZ+qqtGOW5zVN6EGMIw1F7/e9JbnrKAl7MTXs6XXYm
av+U80KcjfuvLMnp0E2SLRDUMm5/LvavjWfhOGDPboyWeBEv7JrBRY18H18gPDi5
3GAI7yzePbcX4q986MgMK6z0UoYL96ThA3VSByNkz+85s+O4SVvAffi3KrNsPaY6
Ve7gBrb52Pu+MxPRhVm54J5Wwo9ktzjUCTcI0M1rpsYnZQkCaqikTUbJZKzx6aCU
xUN9CJdV4kR9o5YVT5Vcm4EDSxDP/fvdGTBO1oxFJDRhWh51zIOfsgopkBo/4Kmr
5VKaBAZb8OB+N5U+zFjEXMfzqY5r+TJ7/ZeJGvy0TTqmdJev4Z3cRLgzd5uqm4Cn
UjkGWp8SqL4MBLw30QgV8P7XR5FARfPqGRg0npxBapRU0IZS1vGZtR/c1SPpdjlf
lZxwab6GLIpxVXslysG7ROuy+cVkXGDYswUyYzEecnO9lzDHYFCOTjxx9cXUtH8D
nJ7JyD+VO/YVxVfn40+3gj+I/txn6giS3DrG73og/8Eq9uT1NF2ifSA9jslkHVYa
5w1WWDEYAmtJ+lR1yjyR6zZrsKSCBvCR3la1G6LiE8Vi7e+1Dv5t+t3BXYY7MDsd
4RkRAGgItCcEYZneYkhEnfH1LuGfGQ/qMQ/ujV3OC6CMUQ5HBGxO5rZAtREl1yDq
16R3fQIR5OLzl2N89blEGQmjK7LAGIy3+OMI5itQz4PKzUuaX0oEsMkK9xv4kBFe
L2HBAeAbyeO1rLBGcshYj7lqBV0n4qOVW+CCiY+6m23jl8jBjIBOfyHm8a44bvtL
OHQhrrmon233SeilvW3tMj3ndKh+NBQkw6GUhjowZlpx7Af5uIkNeisygg7FruYq
RbRYryQAFecy02NKoC9k2K7P2+BLJiv8WDCa2ka5eFhGqv9M87Ed6w7K7yH9mRuc
HoIW+1rAruksUUUgHXRi5ej+6uGI+N139fqThZBbn3md9JzypbxGpMYNDx3pzkLu
6BVuVLQoZA9kE3yOJqh1l8UZgpDRK5vhqQQ8L7FqlyZp1LjOqX9khHoCvUW/qfDY
b3cwpUNu7vL0PdStkzvOH983ERVj2zw2wkte7dIu0GRIZOqmp+ifkyEXWjM7LHJE
tKPgbOIV1fdgVDfrU56EjC4o3Ne/8PyBAWQT1X5RXZYXWpr2KeklK79ZInHujRoI
HU3C4RWfTEAfC3tDDpbpGqwyvx5rgJQDah03PKFihl6SclufUcokUp1LGtrnbrNM
tJf/UgKorj51VDw1I94XXWnPs9ftR8ftdk5q7itCVp+BiXmffDZx1/aORoeADs6b
a9zhJ1IRPVJ68dJDZOYKbmsktSndHA1zXS3YrCauqqfVdNkJ1PJg+iZmbabHHhlx
TkkfzmWB9vzrIgvVozE5kDQBdwIULtbLzn9rvQJu5lCXYf5w3Q610pVI6JJgZqdi
0vaS405OZ3XxjYliGTQnT//TOHBFfQyZRDjA3mbh/DWzH6okSbUBdEbIlqMzJP5n
0HzNEdljjbsLRWCGx2LC/4RqpbqPEFXZiuYyTFF7eQALT3TYC3eWPKBzELglBvr1
No8p84OZDZR3XdLgkOpNqhXPCaeV37d69MyKZnVQ9BaLb9sxiAeP0pBuDzfNyvzo
dhXDBj0zCeyttiayl62FCesRYb2dt1Nvk5fS5+6lAAV3BpO0/QgL3sAjqVceSUcC
poGTyQ4iL4+MnzamgtfM5NcwVCPQQctX+dhpFtlEbAl4bufz0VoEuUZWx5Nso1je
JH/icihY8ono3acbHQi65K5HtskN0eySjvYYztwK2vCkrAan1z43KD45+6jfEUha
mRsIE+Rw/gvphOPnc40PpjmET26RwJA0yT5bj8ezqEi1uCDI/mZqvFI+wLMQqojN
UnhULUmzn7EcOFCcIbTqiy7E74KrHIIwq5BvmH0NweDnxC6vvx/S7m6sXGsQuQ8n
XWNto5g4htWK38yylqMk0It0jrVGQMMURCzYdcDeAH6IbhmSTGYnQlD6iKZywqmc
huLF3PISm/2Ew7g9WhO+J9f3ZamC8Pn3HGnmSSRx70it55EfUoI6wWz20qmSFKgL
6Xm1Erx8BpFkIYE/BvAgSvmYDhgye0u0QnCSpKYlLm1AmMspRWpOPufR0JM4krXM
zKQ1ssvauta3El+WZBvDxwK8ucAer9LeowXah/3wl9zlpnK46vu9jL0PWg9CUw4x
zowXE1IoBUd/iALxbODM9sdzXjQXVEI788o67mlJHdGKdSfwGSp2t83TQZNqrLOb
J6lY8qLzl2vswGKoTG6D6DBaCgz0U+3FxoXUOtayzrnmFplaSj425wAjLYXMyr8x
cZTuaM3HMs+6BJxXaTy4lIVPwd1hgPTg6lsJYbmQLNng9v0Ozxou3sL81BWP28vh
7LBZHKY8aH0H+Az2e+IXyo23Cv0GqpLffxOGmNIenDxT3cGY3Yaae8llMC4jMEAi
Z/WApxAe07dkmO6OJRuR72Mzq4Ej3oNPWsXF8B1OYqv2edC/v2IWPVZHUHtKmW78
B3IqcqrnAWWIwvwuwuFmU/JjXnf+vweobYzPCS4RpqFk8DhEndEVoPskch6xDuqT
I9Uhlri3zEHBOCbO7EFKe1DAboYSYgoA74q2gyvuNQCSLqK9NFjnuRYa+LIpjm2+
emedezJty1NJhQgTZfgY1X5snEn7LNJVpu/w8ETAfX7tkNZsjbQ4YiGzeHvtNlaS
xrvnCMaZnVwJQ0Z1QBw/gI2+cwNkEYqjauYd9pr7xoCM7LjWiHfhiqyiwS14Y4+c
FPkN7tAWkuN8kQOVe7zhHBTg5kOFFjXBptbS0aRLFIGCYgMCWJWQ4BNr9N5BlUvu
O8FmqUW/7G5WR1qjxJHEEQLuaC+9ifXtPQ+3L9NInP1KsZ7pbfZ2iDQazVI5iqqT
/CmNa6T5zlhgyVV2yQNxxirJJNDTAdVPiLZYkEzuhcuemTZWGzZxMQMAnbauah+G
0MwV0zJFvJQQ8XwguciVYQmwS93wKMzrhvXbRCRfWNWtzXGlp4F0I+/dNkyoCnrP
Vot+pinxnVzZlOAtaJjqaFqRusFUH8jphZiCVBUxbvjKqp5aoB+sDUei1vTc3BAo
nP+TD+uKSVAGFewziQbG6Exu7zmvZKw/8YjXQNRSmSV29uV6GNUueV115R7gktae
2iaVQ0P5v7gf6GiYamdQfirdcQiTdkYhLBRXate/DJlkDH975bqTaRi0orxzTJZY
aHhRhfG9HrdUNbEeaobcDU/JXyYmbsU/jQTr8ZqaugsyfmFd6dvJ3yBU/aUZizch
hnrIO4lkJgMLEiDg0EQ2jrKdGhe5eaZWpJNkvO/cCn76BpErliop+hzA1Mivhin6
wDSd8+OK37cjysKRtct6quLB1qzjoRvPKiy8O47XsYWA2ar1Qz05ecbHLhcdT7Pj
7tRLflenLwAuA7PmBFCWGfxneXnQOF6SDKb47YDIX+j/hYlzpJHKxrXRZ8KRmn+a
CRhvTK1xfBarIq3NiMIcV3/sQzMCYPyzAxr7gjdtMYxCzUzoEotx1mRS01+jg7Uo
kIdQ0ZE3pyHtD8Q9lcywZ27FGYjUPi0YXpIs78a4lR8mxc5ESjTGszJeGk4Rj0bf
TeqtKmeXKQp/fQU48ayY/FNGotAcsvBbqTecoJTpAC9iLCpTJRbvXwBGEdvta7mW
/VcW/+WQnji+zSjC6LVib2iCj57zI0nb9/IViCQyJ9D1QRBz1B4U8MzjF9gUQVA7
JPu5GnCoGU6oc9C0CT5jIucwyfmRO+Eg+7dYhlOurJqnKkS3XGACLwVpN4jrqg+N
eJ+AtS2pXu4a3kpVGluvosx6AYOSWuZ/RCYtktVW2xe3nGJEzSHWDIrLZtgBIo1k
r7KWPcoUbVAw0Lb8J3Dsfzs5cBrVhqUuSQns29+LYdx0o1nuDuytFjN/sKyAYEsx
Bf5R/jVIrqeW9LFO+t3KSj/jru7wwCMLLi8WpYUzuHyT8q+AC/aNilD2k445mYfm
W4pUj1ktYi8lNVpur3hcgUQkvpiYv47FAt8Hwn2T8Q+hgEr4Ayx7Vt3z4bCOn97p
nUn8Wq5nl0Atc/aLXvALYGGwZ2DCMpJ2Ttxed5bwEPV0zal9unKz6rIvuJsBKnuB
3QUl65iurG/+L5fksAcxa+ze3Li+cbKm5btmw5Is2BSLcRhS2YYuqJzJHzSjGEAh
L7n917ZdX8V6TpWKyXYJIjlcSYVJmequdJFcgv0jm2JEuf8u8jsrITzIi9vaS56f
TSTFRyAX/DCSIzaglBq8Nyqc4BigtyKoRgPtC1P5VrVm7GLAxlWQBhAzTytEusZ0
60Q2D1Il3oWrjm+xiv5fLdT6rMR+WVOG1izRg0pJt+e4xGgW5lqHU/WABLLjCxgy
MnqeJFsx/xleZJiVRwxTCnhO4F8+PyUeBIW7jZHut+0zSwTcPjnF9IbJbYFgXtSP
wy43wbj9Yc0kqYFDJvE+1jzBLXiafSFVUdOLdD5R4yJsv6eIRaSAKyhyt0spUopW
ip1UUzoB3+yKLlrAagwTaeJQ+iuZOVhvJfggNV1HPWZFHN5poEOUdAN0dIx7fztL
Y4BZ3XFOvAm4CQwo6GL1s2KKeybKVkhS0Gi+ZDJncUBxaeLsagh2HNPFzqDJBpFN
BCJqfU6+dBhDe3fkrIRuMIc1f3vSNcIypJjYwEnyYL2XrzEVKF8nEu3JN2pi73yT
zEqp5kqDofKnWbWXbPmtwn10bZE3dSJb82HUKANzaSqei092ty0vpsQP2Kyey0PM
G4gLQ04SfDl6l/0/zEZQFO9vnxyGbjYOXOJbKATlByizIMbIlf1jQsBMGDJLFX1J
V+NQLFcw3xMIcgv/r/dFh+SAvlBaanJ60dIdzWU73uZIMMZ3zOC5xOTf9PXZo7HY
k/Isc92cGrbkeakXPJApFuPV3Y7Yzo7ZDyvltRUMpCfmPhmV3t+rfOA7s7w5mG8+
zQDgs4DCUN/zd4TUQWYeK718oUK3im63nIoyu6edFuMlwtRE/PpRZEkbTMV21W77
7NF0bG+I0x23HllQH6QNi9qz2QE5KQKM8kP2OWiL7rnRqmLtoSFAz10iJ90CsRrZ
sVmW3lyv4hj3cYDxcPGakdEyXEaWaS9mJ68GHj2COogljtwcikLr5soefrOGzqel
ZbeVpo8PX6FCq+ucpJvDJHCOzVOZlUoxED9sQxnWcZ9fXzH1O2Qdc85pvYe/kA11
pOezR1p7hfe9KcW1x99bF8kS39VKzUzNrEPZZJ2Tgzd0uunf5w+YL9NR5ykjKuGz
LSSMPwwpiqdCPTi+KVKA4jtYVDykRD1qnu12M+RoNkR9L9eBBYiCE0BnrPSdo8b6
Zw4mUo+N/258ISsyOSGMur4iQAXDQHCfa1lUdCKGvYq8OrMFkStNGaptRjXyk1pA
8enoMF0DNdavnJ2dHHHKSMdkhAykYpnbw7fjOSH/tv0e6+TUWWmJ0WMpfFfcrlDa
iqrxADjmqCEpSe+udVDq1zomQcuS6FwRgcR56qgUoSTPWSc32RoNtk/SaCayOznf
o5ESqmJ2aoutN4eZzujwjIhxGz4r2B3/Zq1QMQ62UtH7tXEb1w7LpoPWq3mr3ar2
gL9mq71sP35n0tMtBnS57HOo1Dg06z0ec/XVEqOs92OqY503K14zq88frKtJzxZH
kI2vovKxdnq6w6eIj5QSNlO0K52H0ZH658NGK8SbDcgrHrVNFVdrc4Qw/amNF7n0
NjxwODvQcHbhY7lvHtkEf6WP174HaBFEvZYKtKSNeAukXoTjzsJT4heQNDuoLV/Z
vTrZDqLDbumNPgZYtmw8YqFDyYkLCXTb5H3Mfs4U2iIyNYiOUL582FdMfrI/F5H0
1rZs4PmKec7PS2e8g3ilQjbZm033k+DeORixmAnPqcT8K/duzJqtqMCLj/Yk3xjy
SJFe3m2S1riJw4bKfeqS1bt/xHn3h55fnXROEvgzKOEk6mHxD6lkDu/BaKPXevZz
91IXuTcJxUZMVKqUtC1yDr3Sw1gI2CDjuYjCOlSP/KnL1JuP7ZazXau+hUQiOucy
Tf6TvdAxGouVRQoNyNBQjG+h8DyIdAlU9fGI0I/0SgbEjjsvZqaLr9M8hTIshk7G
80SDALLpBWhM6dPtaAwx37MGVKwHAM/ARXCCU7Gko2mj79exz6UX7bIh0XbkFKCj
uPBhMZDdiBQV99ys/mDXR6zhLUSsHujl3qtQizaQXVD6bAdnsHXGNNpJM1EW3KBn
rVJYHvrMqbqsAr1g3vZrzjegvRoSO6VhREQId0gBJgp0Z7U6Jk6firgEm4gpMhIu
uLK7s0/GwngtQyDScRtz15oWCKqUrPcoCt8OR6pNv8je/BZzRarqXFAbXlubv7S9
0iQHzcSxJ9WUL8qcCS/o+6DLQG7cc/F1TZPKHzxJbJTQZfl47iL579/7XG+7ErZ1
wRBHu2E8qAEy8BgdYdYeRa3gz/79A145mnlK+eX9TSDCn2KYpbq55oAWMje45/Ia
k8MjxfKUqGtt9NdvuSrHlsmwlw5qGIBd7YNY1fI0bYZYuc5BBN3rEyec0GfWVBy7
mCMuPd3KbNWf41+J68QH0XmcmpWIZ4sHN0VRRfgNZtcSQCdTvfvmN1yY0Ei2mDdw
dWVybBx0WaVpxmYF7QY5DFfoVeLCgh8BUyIZyPpyyMOdT7gYzYVeTwDkmVhCE/z1
E/WB0VaKvNsO1Ao0tX5wFGQ0nr0CgbU1FMlBW9Wlrf5gtl3JDp/yZgulw7xhUSB5
B69lHSn5aYfNJpg4l4YCk0xcpVxCTwVmmCU27itbQ9MdLRmpt3JyNKxLdVCc5A0v
ja15BdX9qlgrwrntvU4LJdjaiwe8bl+6y1n6+A+hY1lA6YK/3z/A5MWtVe4RMUm/
khJH7FmsGWT9hduXJa5gvFK7CBxQwQWzj98uCwX1iq6p9KZ7CpYXUWE/TYgYUJ3b
J5OPS2uPoC9ZkpzKbLbq1X5yQ4jg4YOVUdfZUrGpAJjPcZJuTrh7fug9TDenx9ed
8ewvytSx6jMv2ZoWyfwP9OrYS9awypXhnVfZWM7eVAVi12VTVgJjKlHlgTfBq1xT
rSrdcZbxLpwB8KuWakhQVrh/ybFsbL3OWdq9wMkMtDs1oInR1pj5jNNDXSGuPIae
KYzw0Xb/CDBLev6w6222IoK5/opsDBa61GEs7OjMwAGKjZlu3uZYUa5rZXkAIKQb
EP14eDGI4OHBpxqR55+wik4WAD7K3Exh7Lr4jt9Fl3xmAqtNO+11IgAzoNM1zB6A
YlvEWtPWH5tU4v6Z3//piT6KXimljOMhsNVygch0EUikJXRJXMBbVaDML8MfcDtE
jiN/ihVHn+3hPxdQuG9w4VYyj7/G3YXPErMZa+SzIkEQiB65kWzaG/p85FSXhjMu
8Ysrf4/B+nEHlMmIpUuctX1MEKNk//HSZZchQsQSoPE28BmNGx0x5bPjKJp0JG9C
J1JruMYUz/534lm/EejsZbxndkOADfQLxPDU10/9BXhUjIw+ic4j9AGZwePIPRoG
MCKa9patuJvJI3Nh6GJ83KSMsuWDQz2sN1HkjmlUgXS2cjRFJUFpc3c1FHIYGekJ
AXbkmxoXD3vuACDwdatJdetBM+3PYuzavNi5ifXbyB/j+Jz0jqdvtIHsfssCdhfn
fDOmjqj4Z5nN8s54eaSCcWadL/ghPa01U8zym7teQV7QCzX9u9W4DSMSSbXWd/p5
mxJlJJeN5dIXoY1yiiROABo8szRBpLruFAs7dAQ+Jb/aNnen/PP3U270IFtqaL0M
78nKcHZIYmiQDlX5YTC5CkMjkI6wLC2PuFIfPLrjTwqENqxj5QBqbI4EKDBVv4BI
ym7esmUAQQlRdIGa0hVhkgsISOXhwFkUjZt1Vr6PYLE80p5D+5/jjIaWoS/PQ1cq
b9JrbKAHA6EErs80GTlMsBjDCnEjNxHbNqMPx65xGAnrQpNK3v9bw+Zk5X9s5XX5
mfGkTjAKBRYK8nZjL3Mw796eqkG2vbRwA12uw/f3VA03lpqAYZsU6ukGlXeaUYsl
Y02BXtc2id1uJbvxo0JBx8voBZ23WuskZrutUpnXmc2oGJvq87qr3Uap0Z/GOw68
Vomqfj1BLO75GndfHzkvi7K1RVbEIago9QkSSd1T7d+Yk+OFGcqQMSn0f3wLfK2l
lBpoDEyRXrp6G/ihfEYsvDmgcLJbGFfuS8MI8dJTJF74fzJga7ZCgkh8pSR7CSEL
1I+kAsmAt9bEsxA9VbTuYY/6+zNH4r2N2OXFPB8g7nCRKZHYcQVIMxOKhGtuHldy
xy0AfqxrsIFcV3V6DhQuifAsNta4fAakF5e5OmVGupOzcJJi3SeNaC7Zen1LmMDo
AoTRt+GAQ4+nHeqZbTufr4TkOwqzq0WldMVlPBOstoxtbAduQ/OfXCI/plTF9als
NxMu45MORS125B4L193/AlYgTQrmSDGsER5IWl3h3wxIze7t/+shIQ37nPv+X/ZT
CrK6x7J4rH8VxB8UFdOgP2CZp4upmANQ1t0+NNNPKof76mmCccODgKibAERSD/fi
wij/wofGTbhsOXGKs9WzJ2TN1a3XW0PCQ1aF/v1NPId+r8Dka8W8evQ5xt3zfHRk
lDt8av79pclgMkxI8YBB5gIyE1W3so5l2sqvMjcb1+0RU4CImBKymzc+eRx5M5WR
7/6wrwGSoM9MI8tUuT80fbxApJE7n7l0+Vu5kmCnIH0pWbMYP9x+6Q44vkwNo+Ee
YQErUA3ifY+BpfSdzmAbnCLi5durbKLZdfk4n7zGcxymb4JZO4ALwRWRUy6nyesS
uh2cpJBQInLn9jVzRkjfqCveDfh250YgNuQSdE9G/hzvpp12QjZBmnYPp1+yAPnu
qCaSE/NeUdb3ezvVtdzfw+8aictTIVj+KbmaK5Z1RR5k+Pa2aYAbqYj3pyAWmTNb
VlE4L7P3ELI6D/1p32cRl5VLpBxdyqb+pwmf6lJcyrzxd7J5sK1mYJLMEKlBAg/s
gPXfFJ0HVAMoa3JfKLFlci7ps7CmuWqo5uol5Ul7eSVss6HG8mQ+okNKhJdrSSyO
E4fKfg/hjunSZKedd9yjSHGrJC2Y4HGRpPk44QfiEZscGCvKskESZII0QMaUxQ5/
pDMWGOPGPCNDsH7WhDOmw0cirYaa4R1Yr2BW3GRBP65RQjmfFoSHR1Lg0cTthWJj
KZMjo8zyo48sT5M36CuUBHe98fpUlCqBrmBT+aDbndYVjTFaBqjKQIbXeDxEEADE
JnuU9LSNtRRleSqN4NgJTR15YOwUcFFmGe0829gOVRXHgLNzz+Lj53nj9GONdYYq
7QtokfpF34xfjAyYSi5oKDA8clM1iO+UC+lMY6FcQ4Ij2kzIFdNOVy1hYQhaVt5H
q6Fgcu7nlyd46w6x5YWtpQJcHT+boerrjzkuzQKY4ADTRrHQbmCN/znGh2rXa7OX
e5U60J0Rk8Lb6m7OEIvZKmdwRkLrRnnv+2D3HuonrPD/dgKtRvQZkh+LxPQVtSyj
YSNxGL+D9HC2tC7h4m3ndWFIepginqBf52OvEBbJ49n1qC4SlmaCKA78ZDJUXYgN
VhQ3ZNjRXV5txJKiNeB5SC7m57lxR649XaNzC89z8yogTUpwceX3rbKI+bnmO64/
DrsOlEN+eQcTOp81gDDV76Xsh/0RZx6DKGUYlntZHsH9sGsCPl7OuL99yVNb4Vzh
UhvAwU+c77kN+bMo7mg6+EjKATDmiT+yskEiFiWrIr7v7nxDAPrIJACPKaWXt7Lz
pD1s+s6rxiIRTWwPsSS1uLZIUbQkjTjT0DAAcC60LEaoJL7a52c+420exFzclEEP
hteSg7v+EoTidllUkshhiTSa229PTRRPVZ8HyxLOv/kP5Yu3TVmLA+zz8WeJV6gR
EMQarHewIAf1UY3IUzx0v+ZyF3A+2P3Jm361KpC77yS93c9Sy0olpxdJBooH5Suh
3FVLF3DhAxjs8ok2xV949PacWY+Wr7HRw+qVYt+sWr9/ePhK4AMOOXfToamvObkr
H7wwYvwrhAI2hDCFJ/+f8oCVHu0n0R2apA1H/B1165Vtb75CqXOSU//SGbfRY+mB
kL728kGzti1YekNLuOJ2fwULYelBzwsiW0qm31wXgblMi8bEY3BAYCKuIcN3a1OP
dQl5LIyqUGl2KY9t0L16nc004229Zg+za0j758MmdsULXVrc5iXNRHoyYSEeHCuJ
1vv8UqN4TM8G6guGhDO74DKAGwR+YtPHo/i3GtqIR/QXe6Q1RNT8v3XV8JXfNmLW
McNoL9eTM/k3fzKnrCnbf40eDC7OAlA+R5czfUv7bV2JE+oM36rob7tCq33NgwA2
tqwqizgpyNgZHVvDtLU2fteq7pMcS3V1SnrSD0y72E8AU1R56ixw4m+pkODC0yJp
kvRnKgZLqWqUAYCiQVIN+oyo17aTOQq3lMcZ1XlUSYeOhiW/9LiMOoisX1Fofd+t
WtWeaYPZc21RbmU0KDRNVcuq6VNgNqtTVQZCAD4UngLP6S4TfMfa0pMVkxxsDuRl
cj36hCkFOFlHhVC9wj8yN98IPejtt9CvWVy/TGVMN61/Jy4uhgwf+6eKwD3J9hRw
gqu6wMdACnnn4Z7petBuZVSyFNAeC2WA27k2UWiHxRn0WNcVosW/lqKoYW9yKJav
V+MpQat7YfRgCTRcTDu2+HgBeQYoeXNDA9d//LmoOOFw0reo4EgEzh2Lyf5Mwp0w
9xnne2jAeNH/k2cBJNK9Sc1HRrSLzUAF+ZBlwslfr1fCCY18xCSMH/IuyRhPkLQV
K05WLEUwRNQDvdAY9Cq7z5dxKnEH8PtM1snm6nPQ+3CKc4YJMC64PhE3xFVXFSEI
vgK4cLuoGGo4EwgRqHrfQqgNtp1WMxv4yGtrRiAxwtNN1NRu3VBIW6c/MzTLfFFX
tCBDnU4rGkkPROwoA/tzyMsn3gr63QRAoN888bhw8HCY6WCN7FB6bcAwYgC4pKkG
MZ+cDVfic2+nWHuLAVoDQ3MQPkPn0iwqv6z/5NI8H7KLrjbH7pyyxuDNXlPDnwhV
3h666jUn9zUf1SWrUxAxcAVpGO44hNghy8QAOUkg5ZvVywL2GfhHhHkMWmDHpyfw
AoZSQ8XqhCRyhvlT5For3MSeojY2D6fimcfooBidtUCqarWx3BJAaUZUgeAZnV/Z
tgUlHThdhg1hmkGhbNPSK0sozPTUIawX0GAfVwHZgWsFrK/1GzCyL+fEbBzSgXOr
EgfDYjx2j3p+CWk1NFkbty3pS6qIiQpoEnsquLPwhJaz+DMFKND2CEAxFrt4lkqV
4ZMz8j/s7tXxofeSCrgnJvxWbn4VNli/L0n3KYhpyQKoVF31RxJRlZgtdBc3CWhn
Zr1rgucTj1fOvWbm4QYvvb3PvLxbyGZQNXxi1aquf1FoGM+v7kVHOU26yA2azSCq
LSOEd0JUYydm3yDg3DlldzDcAWxujsb1/j9lmLwCvxh6xjCRmU8EAiYlVrvIRjIS
WmTtTVP8HoO+aWaXzVUfut5/WQCQRisX+eHjvyJbJkxjJ8Yp/Pr+QeWM7po4q2la
z5ZCUUxjxDHxtVPnPvqE5pZRs/GQG8Sa5VavcB5GDW6OI/JCl7BszMSJYHI3rC5F
L6JguTkEt4GDWgpbM667hnpsTuL2OF7IiS7zb67g32IpWGE0cQ78FxwxTttPU2Hs
lZeMrQCGPX6mN2eJj93GIoAg7iBDLElwQQhLFHoXfq+0NgOGEt9VqMtJSCOQLjAG
jNzrbmDsHG/egXCZmyB2mkInAu9GHT4FMtb3CTFjgO3qmD9zXwdsYYEqVp35yZzR
TEeDaubB+b7b/US/UUWxs6tm7zCqUpLTdrU/KqfAiGQnkfVI67oe+0IG96wT06N1
RqWuwrQ8qLcZq30NeuAqRhERnRtAyvVsno9xbu4C7+E6I1P6AdylsHOoskgTflw1
dkmnaXLuWVxA6fTmsKS2qE4xEkbx0NAJQS2gky+4l6G5rWX4pJVH8otHVCqCA2Rw
5JU25waKHGfraymF/5jsrOfLlxbfbhwEvEhEKNwsCdVWtHUE6zfPZPFU/YDhBEM+
6fUYOG31BNeoeEGQJVJ+YPTMlZIpG3AAm2Yzr7ZDneyB9Qqhju682rn6tbSCpnbc
D4QUaBnPYwSoIPshRlWEMwO+r8AlWyBs167VxnJhg+yJymxvDWHIuHGUGjN1hu9T
b6xSREVoA0NVjy9vr0dJMSG8sijCeqrNdH9guIaFSLvfduZfamsp5UZqrhzRSM23
l5S9Gg7bReQkPu0NdH4zaCugRbZtIPwZHaz/qfJgqg9ftSCf804in/hF+F/UWpvd
yujHjoFoX4i/IoZm393h8scylMhXk+9pXMi1hdX/XmiFMBKo1rjjPutmNacezThz
m+X6bmST1gA4DpivMSIYn2eFLGeaq/s/ZgrpBFvhvlxwjN0K1w7DPvnJ+nPEVXJH
w4jc7TavxQSRLKmul+N8hOqeSh9sn5i+JR++KE3n+IiAywMf3gM8CCa3bRXMr9zF
YqwRuMOhkAkC+elhdK0HJyRWrxx6AvmxemyHhcWzLPzkXlNax1zFNOR2NNZQtNfl
gE1G6hXwvAJxJucATMOQGiJoI8I1JHP5XvN+d6G9u1m8XqaiisMGH2+22ffTNyAg
DOObtgS1MLEdegd/XDC9aPbP12YfzTUoyeXhULgZcJHJnMRZKFNpDd8NP6T4G0qu
s8ry7vd65gI85U0RMg8fo3mT4qespCzBZarxWVezw3+FWsqNJHxwD2eSDZKw4YdV
EVuN6ot78a/6ebYz9ztM8YHOV1xjnV3GPARbYSPfwA7y3abETk6hwIqUzQV/57HC
ubw2y2kKDDrn/VlcS+FauDt6z5N5AekgiynZiI+YD3kuQ9YDXjHL3gYdYqfP0rJN
fiwYfuhD9fAtWPBd8+e1fP4Tev34uWiNC4KjWH5SDql63dEK1CPR3BAcHHkZxBbU
ez9IIUNIe2m7I86/nxxf7eWxRlsmdp6PrWp7wEuzyP+xEyQtICL+17p5DzPpH9tN
LWF5ZH4MqSHaE9IxenmyU+vo+zogwCJafbnd/uL0NJjNWIP1RWwGX8wVEncRel+c
fdH0KhjCfFkwNiShrpjY0jlrOraji9Z3dbu8+9Gxl1UXr9eJyo83okyonxcSKOs9
8X5NmifrPEFCVh6dRehod0wUmCEOdowxYGL+O7j4TH9Ab50I3/BPgOAmn7Nl8l0r
7vJ27dsV+9Bg9AmqkxN+wSfuXoVeKwUxVe44QWHRFJbAbZ5JsYE/hQVfcHx8YEdx
vai4UgGzRV6k59kPRHa22iJC7h8Mk3Ys0bABam1opVRD4MrZMcZcXlUfzlYEYhNa
ywuX5WNcytQU/scMks6rMZJwT4dS75OuZcnpHKVMyF/jmBOMZyw1k9UW579CILab
0bvQs9eH85Ig8zCWIc6jnO9puNaX24bI85KJxWa4CIGAF7YYBdYt+2ZWWUxvOXCh
h9psJrEveZb9cYqfGaTQ4eEkoYmBaL9bO7ZzFV3rYz2FqmmmJ1RZexlqE3FrrPs2
Pto6FEp82ybFqqdpHeTc+XReQyWHnxtRg3bh91wc+X+vsuGyVTi7RCe292JeIDfJ
Wp/WSInrhIEq1WeicI+lC5nJXOrRnDHLLJQoZzEx8H1TOq11XkyOgilWksFEClry
B6wOWQ97+8gjB0HzEJOL90onUQkpj09AosZ/Nd8QakgDPSnh74BigvyC+SMfNLqG
sx5cjeiIBV7838IsACqvUEWzw62572TiLpT90lOt/Pe+g75TbZC0EqGT66QJ3z34
tEwYL3d7J6GbwfsQovxnUaUuP2CdV8OTe40V+jjPCqRQL4Sgj5qI/Z2w6DuCxF0x
46bcZBBZWIOueYnjZod3fi2j9eqoxI9/HfAAXwN2dsk3ALkYumhkXwteC/GBrU2L
dxmOzb2l+5IPr8Qd2Y+M+1gqQLKM7dhwto+IlsPXzzAPBYQFwkTHTpiFReO/n6hg
Ep9PYa6a3lE9rAwiu51ynahbEnrdgqChYLzTvrNiH8PJBWGRurL0U7ZeYgcDB0lS
i3EGfRV3t9f3ufVYSjs7vFH8d8oIUACkrzFY5GWbITLY3kp+J5056s2pksV+fZup
0OGIKWOBCPXPLlv/iz77+JMpQXr20XC2isr1uJu/Mkj7hsQaqPJ+As0Z6li/hb1x
+9jKa/GHwRj7RQSDYqitdut/h9I3h4qQssT8ZtNgf8GX5Zl01GTkmKt5kc9eRqVR
nP7sAEm8C4h8DUBVmdpDpNNm4IWuXsxYLTkRnkbzd9e+YsGPslt9BoGFu4V1umRw
IWfgGC5S64f27OHPK9gapEAnxWK57O57M33kt/DO6kLns6PYpnATb+IFz16YUffM
n9TDTlwE/TlbNHG5C1IpXSf8N0lifNYM6BVO1P9sRvK5rQusWz6Y2pLU/9kWftd9
jhgP0ONyYj/TmifOLHhJY/zXfHLJFOgD8dKUnkExWWpLZpo5luwr3JFMac31wy5y
L9xhMYtaT9gYavK0J6kPeDArJMxN4+FN2svVb5rKW8ECWyyYTyERbm0+Pg45hFyy
p4ETctW5DWqsairDpWqefgKz9KY2fVkVUmcjpVhmP/Ifxe39XAm0/Bo+pNTy7EG2
hI2Nu2unBVyZgLe67YzPdOZYcr4vzN3spAKICIIrVjMsBiGoUb1xuVhPtBZAxiMh
ZIbHwHwVZPfmH1/AlRl90smtLMPD9SmO3i+gg3L9n/4tKaHXS5KqupIi2CgZELVI
sLuEi1AajNf2nLNeZ8+KyWzMqpnE6RO1KPwuf5qvN8LbRKZVXSDqG34ZxbbUmNUl
FxqpiBVcNMpN7fv2SXGUya3SRl7+yqwqULff24mhL7qG9X7hWxewMrnl65hAxBom
uQHJ2yzOCWgKbEovQm0kGpeJGxm5FuYsN4lFFeEa3RC/N4ozvVK2ryXeaB3LMs8G
/b66ItzLzuJNAq+ny5F+h5c0REShE59C31PPUIqAGQoe4zKK0P+eqdcB3GvFomYu
m266ussuNb9/KWvNNlkKOgGao4wyPkTyqVE4n+QjO1iyPmr/L2n1iQNh5lTkhI0/
W48oCaRLlTYOqGkwveIxn0aNAsyEJnUG0rpJ8jmBfCj0iYvkLzzcHS0EQuWCETVl
eaU0mp+MQsXaIjrpL9XQ2pWotkUC4+0Am7whFuPfczFUoWZrbLs1iO0BRzdITdya
o58T7i69ZJrJ6MowP2foTrKE8CuRIuAJ6/bM2rS0YVBHkd9nZCK26ep70y4CDx1M
yr8yxbk+OALQFEhyVvKxaTYNmTr2UwHCu4VpkNN9/HncF0zUIM908HQPcvnhQ9zE
PHrenVJyutyenklafkU1So9oELzO2KZ/LOccUC9oDmlMjcc6oXryu/94saVHma/L
AwGAhstUrcSzcPerVkLKKJTZ7CQ78TpctwORIkigSdcAeTqjE3/LlyQLnHobTpDz
jg+771wFlXFpBuiwMcCqr7KWwg8HoFrnu8jnBvePJ4o2b5o5yfDFaE0dgmObVTbF
kx4VAsCmtXX9r9pY4TnZy7OSM2/XdOM66LlptYF/S2VaHGkzVcTlB+J89oOl5zWl
A5ECKOsyRYxmcienJIL12l+Xsf/hukMChTCgRZw8xACwqQtexFvz33QNKDKpgeuS
QJI61zNyrd8Vp3t7x9Tl1xGHF3w709ahurhdbBGgHuGWvcjzmJGPWmFmxV6riwPT
WzM8+Yp8Z9IJhhGHThBC9ueIyXIj+SG+3ilSqr0+d5CG7k/k9WVcrgM3W4xnRUV5
QSmYvkaGnmjyaddFswYJA6x3pWreqPgDdrW0kSSkveyNzUE/pOib85PHVMr4hJHO
oqJx9OJvEksZEmKGw514L2MwvtfsEfTNW3TkdGEycUn5u9HjuM3/VORrKhVWs/uP
bVhB59OdPM1UAYzq9t7X+wtucAOnE7wDLK0EEz0G19R5hA4Cl/620nK2GpuzB0qG
pSh3IDOc7y8xkg0mWAI7Pm0KOIy6QZoYXVbhD+f9zbyug+3NBrbLyi9V4+e3ayg8
rt5ojjVyTgVtIbMyQ2t1nBaWJCWep+sks2rEW7iyleeiBA7DlHvBEkF8xLde1DFi
ORV5erlcNpv892/c5bXgRq8F1zOBlhUt+jUTpGKpnpfl5j7boK2lPTUwefLoYIEp
gpHSe1wJqcD3tGKYmcthzFUm1S0bUfiMvP1Q47PpsJAbBzj/uYh/zXw5aByftEny
6y5FCZFrhVMfF4tsxBB2cf3wgVucMDeaoY6vdEi1FOoFE4xXYtO2yd+2VtF4VzFp
Fo6KK3Tr+AH3xlrGh8fTqxGFHCnmGQsim8JlDTwReYZgFGaDqiUh8oceEw7t9U1T
YDObCIwsJEmW3mX2veBGZlZ1pBd75TO4K8LDOAjylOKHRK6owNkNPyJIQJAsYlU/
cDmK3KmPPa+zz0SUcmJqqE9L4Y5dTF7A9SR3NkmFsMs4OBWlBJJIvsZrLgAEJ0ja
xF2MfVgcY9XtOGqCl/e8p6s/vGgTip7xfrLvzkn36K+TRrPxZPW3t3pGjJfmL0Pi
DweFT9KF5xa+/Rmu+j612X3D57Z/uf6Y4Ec1VgK37ggJWxONuzNQA+jwyDc8YI4t
IJMkdqJwqflEfPpBvvMc98rqOs8iIAF/Yjm81eYI1wlhNziMU5ed5xHVzNbnbdBW
IU0/5JIh6WB4UOQuoHsMESViP4dfx0To2HYki7mO6/bY+rKfFC27R3thLQNvJLmm
p4RDuKs9idaqZNpB6MagFYTLKdLreT8fmXkFawO3fVc0ukPClwqSsGRYOpix/e+8
Fu2Ev/aRqDuxho7GNew0CklDSnMFctM/rHC2pqLErIq4VAwDlZYELwBc5VPHcSEe
L1W16Oax7HOEAx5zH7iv/xvhCt+Mt3EFLx3XOERUd1lJfR5xo0cXv0TYkTvzAZNJ
upIq/Y3t+40OjrbeZMZawSMedci93pdkhRgfBhC1YdiY+08+p9fmWxew8J8n4eNh
OobuOzHiI2tS5eCYd3nEBHB+Wczwbm2XeVIrH0ckUgGeBAasTfA8u4CLVTsKUfcn
l+7g4ZTHCx2//wQQhbB4x1WqbW7yxleFOMcK+MqRch6bz5LOIkNfeUMQ3VmrzeZl
rhvcBf+vf9VVcksiz83iJb8nyBiU2YZpuuYLQRjaJ5KMwhN8f5acxI+XDp29cgIP
2jVNegkHkjLpI69vG5v0hNJrf4sQJ6L110CZ6o01hTil2rwWQorx+bUiQ0eNCiVl
P/GnJVD7ATMLwLFubePO34k8Rd+I7Do1fvOO8c0grjp3Q6zibtbU8GtmKZYKiQrd
BfUHooHCJ+bRuWdkflYGYWPYflyGDaaMNGcjvlIaDll+0/T5y3wyfYlhaIgXR7AA
ONA8xyRYc1ywxMMtDPqRyn5AuqM7bQujpbvMCod7lSYWYPT3kudS4sUfvfEsY8sB
hOIQb1qRNqiqZivJ0xXE4JiG8NgbgnybfjDlpUqStr62+f7Txb4yLWdCOJYD9zcO
Ri9oDkYAkinsYrxnrVjxZcDJd6iVflK19b6yBYUv/RktdYYFASs9kQmAPCLYIWl5
8ye3dFNDqlvfwiIHFrjOCqmPSnzuDBQbFHSg+GVfMBGSkzhn7/V2YhnihKQ9WPzo
ZqOx++0IcVAbK6JhnTE0x4av76FaIqQ2aJFBZgarttWnrmsTInzZbGlN/nuHUi09
+n4ANwB94K/c4ONEjltMVjsNAlRsgP/8tL+WkfAgxvJe2oENwnWpEwcw7BMLLIUK
rxSQqOn56cA43x7ukYxrlN/eyc9BiPvCVvkhnsieHRTDnSIP9MTrqMQWsjr+QbCD
dt6a9PdsB+YzE+A/K7J06AQfcrpf+WksWh4CqJzKaAWzDKJhSAAIs5/oFbKpkP0m
UgZ8l0ZIGhT5yoWiAXCx++umdbMEEZx5bEJg6qr0rl2iFIvtP81MeuxA8Wb75bx+
oNDpcxeLjgaGOKfPlasfWv5g9qz0O/6ap2gt7Vqo2Buy3HOHwJhTvYzC7k4XddUf
Xi0wJR9hx/QPS1vxdh3XWST/kPNVq+3NVHtrDN7VGlA2FkVPP11l0GAIzaCSX4vf
VRPxf/L9JM9rwcotH8VxHtgCgaPYgfi7d+CtUYl1pS/ZAIGz+GLiZluGxaNQHslU
1qzzlf2c2TlWbStS7iwjg02EzaGt6vPpN1qYun9QEACP0TtGgLtlafskkbg1DVRq
kAeySp0v9QMUFC6052d1MpLORwPPkCYxH/LuAXAK2pLd3hrXSrUfLeB//ZEKsoxD
BBt/hr5f9WMeTjoLmaTJsdUYgccYxBow7VoWXOJ0icuTWhsW0MDKc8cWupDfF1f+
0gs7kQbMaoVWozuDxGF25MGyw1d3utYtOy7hpeto8+5yxmbCLzqozQYYiiOjOmfA
own2i/2mtmj8pJC9myiuQPg9XN94hCDqhsUzZYGZsIeB5SFVklOBLFKDgwm6xN0r
znsMC2pG4s3a3lymvu5wwOEdfTVnWZsD9c/Ccihi+FHAGjA4C5MZmgcYrYYHL89s
raOTNeGIK18j0hfUJ4sSOgKHl4ChftWwSEb9bN/Aqku7s4a297QxG8zW3sriq2OA
SpJvnUXY+eJa/6/yIRezKOo5eKCyaq00vFkmh1c+lhLR7ek5OC8vt+npfCJso4Mp
H2eF1LlEVVER4U6qrX+SZmLr3WT+HDlESjMos/Nv5yERfb7Y6eviaykMQxxGKoIO
3UD2rwGpN0VkPCMHOA/r49SLhZN0HegfGq5W/wiBVpKrzY+d2TaajZ1SHv4wJHHO
Ku+/V+0BrqVlnsgPd12jTZHOvJrb7+2TueQxsy07RSxr8/xhd05/dI9UZ6s5ByJl
HwaKY3BjXzmjXvOd6xYqrOI44JF6iaJ1XaiZSNcbVZnbgmE7O0UEgCGdoCfmf+eu
SSrj513XkB7M79SUrOxctb5QP5W7R7eRDg6bzNIJVmMXJ0lnqxCQuFDcYSfxn5Qh
XaCyjsfyNtC5hkR78jHmK+w3a4obs/1UhXiJAUMaWiVfRWyU2DEOgk/edfoSuVnH
KESz3jxFxSZp/78TfXcZlZTx21FsybRvGVmnkhc1CnGAjDMcncPX33tHnocGrwvV
R2VaI2dNOkIHqe7QPZ1LdjNCByOZ9Vta9Yr6a+snhpmPmfBua01SIG4vY2R6aeZc
a9KVkxG1DY81ZnTgSrZx1oTRtln3Wv9aTSK+1RD9/p3WtxW+gdtCZ8uLqCX9S3sb
sPgfCfWJRtIALmsuiSjcXc/N+FME6WzpM4BoBHX3yGdPUv+2Yc4+YnqZHXxccUs3
ha4ejNg6VbG3r5hfK0ugU7oW7EjA+H9Vqqa/oP0W1tDXZxmGlrTN5LvrixK15U/E
GZMQ/wKTjOIJgu69W97qbcePju7Q87i0pHOEsMtpExhDjSjOAU/LZka3OjefG1Ep
yFFBhmg+JUky59a3Uh8I6i7pJSRPWYuLfzhTtrfSo4Z3qfA5EipaA+AJkyIoP8tD
8eepeWizeEucHK8PV1bB6qm7NnaaH4zHfWUQ9EsQR9O5FnbByBuKJT5+KQYtLJqZ
cZT3Ky0lGtwKog6FDfogXEQrs5Ev06IKuomeS2fxkbEdyERmJ9+H882ms+UhXBJc
tKtOdl3cfS16Fw+JlDthEEGzEZzmtEiH+0eCvgLeee4+12+sPdHAOnh/m+QIO4sI
kgZB0BYdoYOdfEM0sBqqNIoFqg5Yzc8W7V1hzroFR11auR8tkKLdPSlWDDHX2k5N
NdODLRhAMQONKNP6gkC7JSZist1j+XIrUS8NG+5YQCL9xOVhSV2o0K8efT2+fx7v
E6B66INMOTWsXR9FPjCtVm6AEgPjQA6syl19xaGrzceP8pWdqwC18jz2SsGFTa0L
ded6vW0Wwq+H9yEj6/QDprFnfp7oixW0unhQ7qbNQC4rPPgXhW+5GHSztgK6TefN
T9FmW2E67ibfpPm2Bt8rCrEeJgq9/eaRpWEoCCbwDV2c9Pxy7xTIV8uMNkLpoMYb
CGEg7aadkGhP4jDOR4dmfci1TXBvSWpjtExgSgnp4PGmnaTDMUxqep0LijdOOflw
U68AUhgRap3ZWQ+sEaOy06VpHJO/hrL9ZHhyTjywd1P6V7zJGwWx+Q43fp92LwZr
AMK4yLnarNnvvAF/B5+PlIMM8fP0Jou7Ws4nlqP5/kL/C79TwmTe0H/TQmup+nGu
VhnFRRoz4zqAXsh/DOT7C6tRSlOEGAr//4mqYhR4KvW+M1bvmeRLdtCEXjdefofE
S/CM3PnNCkuGZoN8qfSM5ao41ekGf3eYqJXFgorygwfT/UQbUeB1qbIa9M4rUtzw
RRvF2/ta+36xcuvyu95REB60O+1r6Yb3nu+FrbjQa28Cp0ID2lReB5Kxpmuo+xsJ
tj4dyJDx3EJKllqmwPKPrNvsa9CEJxBbFq11OGfmPqQzsbHK7JF01zCgWsoyv1ao
wP5tsG5Ovc0JOMRqQYAd4Xiwn0z9r0YU0q68WPHidQ3H1uQWcIRUeCjpa8MM4fyF
MkssQ4FTDipg08Xe3u07kNd8dfqrFaN5pArLri9TRpD6IpNGx2JC7jaT962VTGzQ
nMVG4iDd3fshuVEaB2+athZ/NFpO0bqk0tlj4nbGlhSAmPuLxnLh32k9yxdd64PF
kKCOxa52k5UjkbDdBJPkRpSUAR5k1LTl8W4zfhk0eR3nm9nJ4Ke6+GVT2+TppYqw
P4hQ4ZEY2NIJXeESgdkpH6btJjZTRPoaUu4ISGqQiJcD2c7fmtm4EFNUN8ZFEyiV
O2usGhExhUlIDftfqX2wqJRYA+wIpOzIwJ6q0oheeZyvc3kC4RNTEEiIrKQLj+wW
uJmaRaYFQbASA3he6/yrROL0JKycBBxImk5wk5xRvNSIn8uIuUPecIvDXE5iL45V
v9e/simP2VtcNjWnKS+5No3QstlP5t1O9N0gbJ5Ua/acsELE1OuM2TR6B7g6jpoR
32KjfOSLlWDEwSeHYFWXaMEpcHAVoLndb2RMpq+jS5w6hK8t+KJFP3nHFZdDyJos
jVlf95dTZufcHKji0HeqdNgq8/pekMVJTsoaffDRUyUKp98d6sa0YcFPEIfPhLrH
BoIql5PEWQVkmEpvZt1EwvSYs05C4XHwVm3E3A/f9oi2iOPK2zIoAQeHnHKWBoUo
yG9ETBhcFLgGFFHOQSotN/h2x/kduTP31KG8ViDFCpr7/flaH6Pq8KY5Lwh4U1Ii
y8FnnXnDtzF1T4T90rTbYFdZGWl2K2eANjwv8zS+8MdM77gDx2JU6hkoSOK9E8qG
MWsFyWIyhca+tP4QK+rOfFD94joIk425xJv6H13I3XxNeivBAoGQ6+yLXstfBJFV
lYxmwGnGOfiEAvExe7/lDH67p1LxIK12gCtAWPJkm5RUN1NusSPdLJ1e46E8RSTG
ff49LUM+7jfmaydijweMWyJdxabEm3+Rlhrm/tsHUk5ugOCZk84qoRJMHOUkpIyV
zZRthdlyLosO412DxG29+Y732AzJsikaZL00SA9wAfXTTBRtR77CYgb5Ajkyd/2h
klMfK123ezr+RqiuvKBwI+rO0tIyOQfPcY5fdCw9NaD8uoPrM1XrRZX+ox+gTYKF
p64s53JgjZ6/oXUMKfyXiEgZ84v4FEWD5Ko3gSnwxEL6CplKE74/mp4627OMiKRp
PwYrw174oFo+H1Ds0mGBT1buxtWOsiIBVGtZ1tWYbr3YEswAunK4HMeK+SuUwuSl
B7rktXCUhZsOHPpmjsBuOZTRXQp00eTVK92filgypMwcoA91G3Xl6ca13Cf6L5h5
pUSxgeplS5wcgOTZ9lvC01je2zsNOewkHYP28uPz4psJmJCqX2eHKaeBkNlA/5LM
Oxcoofi5DpB0kXXBH1HPku4GqQOoS5y09jsvsizbiBf10gOOetOtUM1rn11YXP9Z
LZdow52sVOXDHqMrHWXDM28lciC2A28dR0odFFWzZtcV0o8V2uGv8z0rKIUSh9GX
rqoOFHPnT/Uu0tFvVIXMTBnDs4Wt2NXUb0GrHMYRAbwxQB3hATI1zZsY+4KqKmre
2kAYKfAKu3foCphnvL5XPYe0wgg2wx4DpUjiptAVpqpZOjwHHBF7spEHC930gqkc
B1jM0coa4ugi8GFoIrssbzsg8jPVrR1ZIzGu0Lj3vDJAS0kGPK9qoiYigk7XQbcA
xpWX0FdjCTwVUSqMu70hMxySbDvTsVTLAAcOePCWi/TjocHhS81i9QKPWm+noUXJ
uRBtQEnqQ9a4PE8ORl//He9oo5yC+6N5jzSr0ruJLA9YQeRO+3J46HF8LLSCDeyB
L6su/ERAVj96qrLSfPWiARjByFeqq/3vA8r+Vwh57SGgTwr0wCGRHNy8bi1aXJ2k
sQFwGGr4owFS52qWjUGQdC5WoGWy8uOkwBVNrrbq0tlEk7PVG2G1mRyQ95r9sQd+
aturt+B2XNb7FPO1b+SqSqdmrntRrwdFvE3TH1H0zNAMxV6Ljf85PwRkHS7VJMzO
ECkUAa2QDxD3dsDOdbsRAHXxqQLAqMhsxwYJf1UER0Thk2YzMZ/cY5C+sov6/zLk
g33Zwf51j8NMgD1MJ+5LLpNeqMEh9gNUD7GL7DpOAlV1CebkLeURUNXpMP+nSQTH
u2Ir1V/hevVSQZ9e6JUdTn5btShOQAjnAtDAuWv+uzBKz9GUuliM+TWsxe8pOUnA
sz8abr+Krz7HLktQ5SnbqfAL7GpiItDMAa/TjhzUpgXDH1jNA7Fc4cd/3B3IOsAF
PC21jBeXr7ixvL9c6mmjSIzUVm+iy6g4TE6X0j/yVFeSJhPFyRcXftRHoGL1OfXq
RlB6y51td+2eC2bNFR6x7hjbFNg4YvpHXfrg+BMV35tXWTc3pmcLBYBYakQAf/sr
XZ+3PjPwDbkNHVIoTY2iXbHJnYXlVtnxTFCPnzvHreQMnIYvULRA654cHkhsnMhH
Pyls/NrE+M7NMPKSLoqBLHamvBYKQ/ixa62uquCrP6cIDF/yfB4vhNCPOCXFUphj
lv53hzsk70W37naGGmt+sdKoFUfABi3AyEe+WsPxPKAItyXBsuRW+1rcDPjeiUmb
QuZmZqotIZocG+BgIF1MfvWhsumRh4JI8FHegT8gT85r6eDQ5rbTjiwmdTqA9Vl/
zp2VF0yL7LGgj4jOyNywOQVb6Y9p6iiyR1GhksIOg/1K12hYDq2kYoYZajNUabxO
FlJTjuPcD6pmmxRZPfW7647cJl0ovM4SCccd+eBXickVMprDtyjB+GMWuWDd8vet
d65a1hxVsYuc7ZZcagPYZLtTTeiRzz7j+tgqo/azUqgQ3lvvGjGG3FUGLWnL6udT
LuLuCEVB1j96juG2wbil7YPO7OLagZ7/iP9IYvyGGYd/q+/X8YLOk+VFk57LleNh
La3NNeXhZ2K9unCgq5UPQdZSdhh8uoww+gf4M5PN1ARkL98zzpBBH76/LyMZBB90
J3gJ3e7VEog/u59nOkhyi4kF206PZoZFa5IhEF+I4pZSBc230opS7cN2Q+kaf4fs
2R9EmEjI12/zXiA7hvXhojKuX9WxVaEDApCBmGTDxhmZClZVRwYbHDfoSGnrRux0
SfOQNVz53XEzZwkOwzo295XuEoKWWvBFQ9woqa55BD7BLPUkVqIB9OAxcZErFuEV
+k+A+y39aT60jCXYgy25xwwSMRL3FSBYPv4EhwWakhLrh9ubBwlXkhDBl9lXvIcY
paMXoUpM8LPDexiB10kKdtlpWMNtsMIxvPdCup6/EIOqAEKWWl7xAxaVmGH6pEP+
Z1Z08LwnIzouyRSwe4A0SLXjpCQ/n75ixz7IQDAa4b6hI7ePyLEzhvDTy5Hbszv9
elhck7wSCpsXzXcnCQcLzaMIDm3QlJh8wVfnSNL8gPyqTqje6upRgfAAwFOeoPlR
M0EX+hcOYj27TYr3Em+lk8Nb0LptkG0tbiBDwanhrFh3buuOLHOQ8ZFeScFg4Ipv
6+HjKYl9QVnMcbWzACA7dj+ZatTtMr049SUTMrX8V/yZ8s0qiq2kf6InqPy+lmCH
98XSTqGtOR6wWZ7//rlQWPrr75NnRNQkuKlEozYEW+JxMGuoF9zUd5qBZWgl0VSd
y9NRn0u4lT3NQmXVK0PjrYNWwnEl3Y/kC0Mcpt6hI8OqJe42rB4884MjE0brvE//
EK3wdjLhM+7IqxIFcZadSQ/BDW9/jFwNXaDu3egEIwlEbdMsPDUnFgi12FX2isaS
B+E74KIbJWWC5OQzvNomQW2N8f32K69XARn1mxQ2ZimLnj4rSEfeEcxjUQ0wmH+8
PwefEAr42zwSatBGn2g3fqCOw9dIR0MHRn3sdqtu5WkMhZ5nlF543djXGfe3UKf7
pHH7GoQzCziMsXobDNHn1Q2o1MoYKvTgInYqnTff4yJEoO9iqAUYMgn23Gz7vLzc
QA48IaWDWjoMEMhVGIwnHFPkEhpKL5qyF2eHaT0AVc8LcqEO0IEqoQf1vxQe1e2f
i2XmC7SVNV7X2Gi3TP5V40secE7MMOiXSLYHWXi4rspbGMH74f1b4HHtDFltRw4D
4V/lkkLbY7twW7aurZakMJ/jhFSedqyONJpAI8kKx0CW7l6aio8qA0ji3jfLkrnH
rAhfMFJeeuQjVOUsnOBZOC9ebuKcBsx4U7AcA8eu3MdCp5z+KB2PmgAHfnhqb2dV
l9pjKa0Q16vO7GKfpoeml8zBekX3iiJidvzu5WLmxvCAoSmbB49+CzbVIaSw3T8a
C46E5rQYF1NmQ47HC/wIeef7dAW6U82mF1uWn2+qYJnYjVylEQJDMrGB2ox00G1m
xOIXG7E/bakIfMlua1wI/AO34nEKUjwnZ8KReft6BG40IDQEL8PvivxHwUx1pJAa
qZ6ebB3irhQTIz4uLC32L1ZTJvRbhl79S89OyKoV6AWe3TJ6Pr9U/zv40W1tTKLb
24SgsKABhY0xC9vBJzLvA1PryPtD0rCnylLjvLJRTZ8fxZZLlCYobYsXSiYOx2Ub
mwjc5FBNWshYyigERtxlBJOTSSUwUCt509LA+E9tjzeSjzkG1CQFDziHihe83ntM
kmKsnewgfeOOZJckVCdjhfweYrQETleREvBMRwBuEWNykxWCuMVfmlfKIEVRpRej
fMtrNmG7/PWc0+nty7iwlfmUnPGcjYIwFMI/jDZPAj7fXIU6ERPj0llYftYwdcnq
f/sYU64/vLGNLwjb3RYvxvaJ31GdBzzpjuNKApCoPBhUIzdzW0KcBTCASFAQGKbS
rvJFl4URNEhmOfIstfQvE7ykxx60sgHgPp6PBF8CDM6ahGk6RdvB8UilZSzSTufc
dxMWk08evs58CFdDQXoWB8TMtujMiNtKgwYzdq2Q5cwJFv4bJFS47Eulj+EegciI
KnAUDWSVpOeClz0bzpmePO86dBc7lEUpkW5SHei8T4o45aWdH76QroJtjoonEKsw
4Ou5Nz7PYz/A7XJcnIU34uWq+ZkAkRG6UunOnDncw+owmAQhIaYpzqNO8p7zBVSK
b1seCQHBm6r0X+R1vNHsvQCzuS5Vux4OE0Pz2pex+OR5pxSO+pX5nmXM+/cuyHsi
3YoqVq+c7BRCSoryxhD42FXkZj4ds+og+aQG82R9zBr+Jf4ySQtXcRzZrMMyOHM7
40JNOHW0y+cFydB7eWj11wGTVpn09+F4hd+H0/X+VMyCQNK+F6OQwOba1XT36Q0n
LJB6jFUQ9lTYHDpJZT7VrN/HkSf9rS3GZYNxw89HnkJsiSm3dKf5tOQH4cVirbED
iVN9zqeP6LGckxjzR2yjsqWB8+88pjmdggi+I6z5nHQV1eoactcCxdI1zUgndRou
nvQENt02SR2O9+rJiwzQ9/VUXNDB2Jz2F0OQZ92jsAHU0y+dAVPaYPEEMiMuC6+L
o/4/7G8bg2fFRgi8EMZnZVQF5HLMv5q91J+8SMuUIwdWXxFYayZdCWqPBUWPdsuE
RydiIaE3+4M5ZwqdZmylhHPfDmS8ICsBWlwtsnPCwlUBHertyOXFS+vLm9IOqwOE
eaqRWvm3Yt2u6oDXuMitf2X8OV2RNMvaxJYXydAypIlWNUke72dPA7ulSxFEF8gM
7MKpp8NLf/S3lG2Sr+Ot2KLk0HiRIfJsFs/5eVZ9Z3QxItVodrZP1757QLzdwArw
1ESSQaKWITLxkUASjlHHufK6Gqm0GKYOFLsWi5V8WpIMHTmQ7za0gfy4R4eOvTXR
CzyKgYITEwVtKwFWjAoKB/RDZB5K/MxC43Lo1MD0GOaFm0iQkckSnXaM6PqNwWNC
c0noilXgFF2qpoW0w6BFZecPmqYzD9u9i1GsuFJVjCk/VHus9qa9Ns8gzl3+7Zm3
JYhVVzNopRzMag7UV+EcACj6D27iYAGjdy+b3VDApfpzJaCBzBoJ9X6ADqJSqSaT
50HTotzyQDLbVrl1rHyliuEJd8gj483xuDtjB35tL5JMVtYNYfR3cZTlJnzVT1Ja
1OuebMV7ilZDXrskba4kgJslQgpG2BenEPevH505TiiA5PYcRbV1U0yW3sDsxnVd
XgZWYW//328uveNiArWWkF2FpztMfNoWyvkvNCoG51X4sm3+ptXlfmBCFZLY1eRq
cJ5PfJK7pCzcFkr+SSdD/8ck/OLLXUWrGLBiNKkuGm1S4wTVPQmsIyMNiH0FacfB
Dh+dXCpA8H1ZulqCeU6+r8T5RqEH30UaccRYcaKfWcXXW8YI+IOo0In2/Yaetk/5
jKR1H0FaVZNLts+LmapXaJrTy1uFwjYZwPauKACiD73VoE78DoFyxXBa0FfXBaSZ
FObvDuJEL86+0tlEeqZxUJA2sAF3mFRlQyw6wj/+6M82DJQ/dFyUdtgu29ojVQl9
3DKBrkult3zE2S5FCqDRZxNVdJS05fywkI2U05YisKiKMk1NEi4uA+SJWg34mZ3/
YnxpIMpl6oQri9xhuOi/HF9COr+/v9j/6wbhoxxP6dHkDPc9qZAtA+pavmud+Wl7
z4K/xY8UYOe7o5I+Fw0OfeTyza/pnNtShXIpOrEa0Uk2NtyaYWhkN54f4Z5WlzDT
P7aOY5ez5XHyl119X2dduZMG2nLWjTC7EYRPRXBey2HfFw0puRafpG5XSPL149So
syXtF7ngaTUDYNRoeDyWUo4PRKmQOy1AN3yFQaHkotbi0NL5LL8L6+pcLOy3WsFO
z+jEzyOqv2zHNaqOCjKtcRgt2Tc3Sfe8NRl+dhqYoUDGGrpwegwov5rHREfyRXLT
GbMJp5YuDOgh2nlBAi94T99HyfY9Og6aAsgleCWTiJSH5Q6ZSc/QDAiVl73wyKGM
oO9SYCb5uGBK79fUnh7ls5pcFEm7dKa/3aVHz5caD38XW/yLGjEgmFXNvlJBe9u4
mHjKKamf84yIXqwp1+yIaPwjGT4t+KJnQs1uq5pxCzTgkbvu2Ev+fNNLN2y0p56e
pX9e7vz3MbpF3sWjmNEDjeCTo/sBgsUH9INrevDZregxnrUu/oES9dxEaaTskUmV
zXSOOpuJWvuBbeoLzlJr0aKV6iwmpFk6ZH/LDjpQQ+Fwb2Urhr6T/Z9O/HyroYL/
taLQLBUB6pesPU322mTuuf1WzVCPStu4StIPWhlRf0VUagv7uzUZ2x5FHeU3vJ3y
qpl2VWE8y6HROuxuqy5Cllo0LLvJx0RCDbEVNGV/KYp8RWLW1je2dkSyWn2iWiG+
aOpcsnAmy3A4Om8MmoTxmu/lMWUU0YpsyGzBTCc2U4Xd4NjlIc8Fm/USwP7ffXcF
BxlTA+NJkRoDIs5On1A2Pqrb/zOuryrAJGwmo8o9njdwMMuMcYwrisgSe8c5LlHo
CuPYhwW2ogUglp9S6rhgb/3we1+J25mDsik37aoEhfoueoujgxXWUa6hekLREIlU
rEBypZlqc5XQuaaKZpbqP7J9lMGkJL1owy9hf3hN19nDdQLHRTyOFQlDBEIQmnoT
UQytfUFR3EeC5A/0IabbiKf3LQJAqQAygMaFEMqAPQq6L93TXw1p1PqI36IoCb9t
8rNA9vrJSFC4A+crFbR87vidGYd/GAU9PgwZVMUCvExwliyr7bGPRaJvldWDGUcj
OZcHIpD9DCOpWxGJf7mcbX+T47IKlTKAPpKmKwb3uA3vJqKtogDX3fM0SFmfUuKv
C5732CVZxWvMQqyi1xtADnbbSGkkboDuxC6QQd7BnHjrcZWZryQe2bkebLxH2c43
8F+6kfnIFwBCwy4PV47fk9SqtddRg43IevxAI/KLO2QHcJ0rXSQX8ZPPR/ta/JaL
NhW9ysaizytF7SwCZPmR5zfkoa4m7hq9rtAffbv9dw1W7ceFge3bxTWOkQy7IBDb
yybQ1K9WG3/tFoB7XdzGBqGsTr2BKWZ/yPLmQcaYdu6DX9MEjH3W1TH/rT5nVWvu
P/zUEMtiI90xIHAmQLCxyfuN9A/I9t6OLRpCAGyP0zWubyxk9u+X52pJvVcOKvN0
SkZgVIRzKlioitEXGP9j4HT4oEQbZEPVzha7G+m3CP9cjlSAPaRY1TcGGhp0HmLQ
uVrv2V88KRzWuo2cNbEBCR2ODL2f6fiIDmvLLbhDGVuR2+DIg7+Mnb7xIMTdyW5A
MphimPKTUiAp53mEAk2EUXDEU/ZYPdSea+IvndJoFP4d1Pvulyto0ftKHEPTf/aN
+NcyXWOyiSmkNw0dB8haHhgNxXNoYorokX0ixVeiDouQajUbiGLUq/LIWXaOUr5A
M5Xb+7Cn2qDMMdWRx/1tHULpuzRr/9aa+tdwrfIAnkSsgtDAGwxS2MamtLL5wQDO
cLNy0KXCUZfuP9InZQgLUuEki5DCK4a+c4QVp7TuCfG0J1YlfZP7qs9vl6L1HrZd
gK5clVNgFNAHEqut4bxyrF+RH972fL4a/BKPTRYQY+5meVtq5OtOmNq/FKZVaDII
KmtSzwxka9mFZ6gHU6ScLjjeMDGuGHFoM39LoJrBR/vrElO3E01pTOHFel8l3YGZ
zaEf72N7fSsHXvX5M2GFmxAzaFr8bN56udJz5lsa8jvTyKGdWUG1bW9CWVeoGjAy
OyyE+88T6xnoG5bSsmkbRmG96yjV2YhODIejbJM/vs2+69zd1MbzSguU1bWwJ9N6
i2mlsXQD3RqMAO3XjfimG9U051QWqlQRZzAsEwD+fPE/zX+YqIIu7yFYoVlfSjkF
Y/nQdB4hb9Kb402efZIuYx62q9NIwkQwgoI1BytC/MwaZp72k+H2bPK7djbdJEDG
aYOYqJ8QU/GQFwQhyjFl97216Df0CEymfSJELkD5w9Piv1Gnpxg688NPRWL/ZrL8
xsE9Kab8ISH11hDMj9JrAsnbXG34E6sKkWpR+JfX470O57f9SRO9ol3eJdjLfxZi
AY+lVBjDqRx3tYEyC8fUfDf8tHzfBmzXx3CCKmd+HhVceKaiPVdrQU+MsOF5JQU+
ivS0zcj3wYoIcj8kY/IQZN1LRv4HRv9WS1TlEeBetm15ZWjoTcnMIhzi5VxN3xgk
NxzyFQ88z9CfmsFv6c/TRipRG2bM+XMxnErg+p8ba6YgHl38iTfZCOtGKoV0du8F
/DXcppmFv/v3g8OTfjHS0hPQ+Skr5Z/8fzsSuirdPydDokUNWHNdcAXybgd9ehNJ
jE21713OP+t2gZgZGhKtkmqBTMINJJ5emUK3fJdfsFb2wLQ8oVBjLuajPVQIAoYg
bfPcG4HVJlFl9TTcWxE5C/hSglykMuwU66p0qXjVmi/qVeMaLBuyqu9qb6FH+7Q5
FXNNe5dbnpXShPDzJA2FrfqxT0syIw/iz2XaE3BhVJ6zbg4BHXcslVbLGOcj+DjU
ycI+YRecwMzakTF30myphESx/5k61+RXZMxlMMibJ4zzhxa8jeHDrWuYe6lQ8cVb
FimI6uCNe2Ad6cbGEbOw865fEWpWGdgtWkbY6xdWqYETJU8HzYmcYQdHemql9FJp
YRl3aCp3j3iTWvF3Rt+162DJIzozOt3mPknIb3mbTweYsY2oKbzPJG85/OA7vG/j
8Kp9VWxb/6eURZEdVGjXKDg1EYMPj4O6Btngt4eZfiCSwlSZs+2oASbrC54ESsu3
rWfTfDKSrGM/NQSS4l9VZbH/mUU7Sq5cEpWd2p6IqUUKNvkzLFBbOy8KO9Hq1M5H
ggS7J13yOZS/JTr2fMkHEAjNnMmVbJEtM7W/OwrnFi7la2Wr4HuqSaqlc4qvZLDH
myPqYSxQA502GQgj5I3ehUSCkFKnWvVzBe0BRs3hww/dOseCxbrQZWu7igM2eEYE
7DXaP/DVtcMh1XPncTl+0ietrR4Q5NWKmCGeFregWeiJDdZToOW4z23gF+6Nr52/
ljPh16FL23OjvNocEGsouBnglwLFQvmt4MgInjn8jRpjHufHhlneuN8F6KAV2aJM
O80vkPUNeDC8HenCNw6/6K5xAjnfV5KIzlrrylTWn0rkJA/uAkJAoN23/G5wjXp5
/7yqtSboq99p4foFlGZpARAsZ/ytsUBQeOrvJQVgsJxyWDPfRS3FC5DJ/mF8RX/x
e7Z4zGN1FrzIZ8HZLrHE3a0M2gRXWDBeV+oEOlNBYwNbXeiViw2apQ9RIj07nxZ0
+9oAPTxKLbPKcFJ7cDSnz1sXDs0f8EvVphQJJA9Ye31PoBv+yKtkVKlB7Pp61Svw
8CxeqL3k3b1Nm8W+4wTMFAtjyWClv814SnoCFdW1Qp/VM57+Jag99Aift5hvXJdP
EvKiRyuLlCMy7R5PEFWBQ21XZc73qYDgsefCfAaxoIabiBAUXwM8+uEvVnryisZO
WdGPIrwdfRAFGqsUis+4D0kc6oNHDMdUUgKNQ5saGV7tUPK6LxfaPubr55CvZxdW
gv/+vqkR7GqV3lfpQ2gitvHro1Qwem2SRY/IsLYxwzfmhAz7Wme+hJcR6Kw9Dgew
DTa+2APEqHu2DMQTDtIpZF4M1lzwtUa0zSyCYodP25BfWWo6uHsMC/y6Mgpwnwp4
aRqD8CLduXVCbkwAPhelIJfGn17o8S8p0JOUoIvGHIHYa2w2URtsgGDHBgXpHW5K
mQLV1nPQOofoY/cInjZ5SMJifDA6kM3pa94TZzgxChnCgrfhjuGFxVPnUbzzOdgP
aTvxLUSFGRel7V8O3Chyx/w/4LIBD3MMQGv1nUh4MC4LtFnrNf3cBYBoE5Q3IYIj
05THCbyrm9CCDxCp7TCpRU9pLIf0IIV8M3iSw3nqmFQRkE/wUpI1m1kDb1ga4F3U
tZJUZjstnR79OVwksCsKzT7ntErbVaAEiw8bjrCW03CsRQfJikD5hlhtPwX4seNf
4998RFuSbYrdXjudosYOu+PyMsewpIbc3mLgJ3BrTTgvIP0b+DgQ1JFqQrRQAKuq
T0b/XOnwfs7XodSG4BfcCPXcEEB6Rvg21jqe4mJAtTPk1eZMTCqsCbz6Wrb4FM2y
WPGKN+V2xSItK5PinxkZzbSPVTSOLwQ2li/H1wsVfnr+uTjt+CJPdKZYP4gtJssI
9kGfaF5qMurdgkarwP2xVL5VLiNkmO7lMnnDhz0YsmFw2/xTo5zG3bEByIGzl5V3
8Yl/GPgbmBIINS+iaNeiRwFiTDMCxPabU1loJoZlTj28PWGc+BAfAD616vkf/Lxt
YOIbd+8ZZ2HYsg5aWenyEp0RN0wC0zrtsVcRKBVzUAx9vB+wdpWDKyZp4Qjt94YA
4nPJ5pKcPLMoVMtFv9XjbAu1ea9OUoxyTKlgywLMrgbf1E3ayLO+C2yL2gh921iS
J5ershCvnK1iV/76c2IzY9VqIyQVPbg8fBXvue4Cl1P56Wwd0/PltRU5XZOtBa8x
ETKdNm/iaBihfP1RTxIiH06QtzUzcSLYiTPV9OBbqvt15xhKwZBfIBvrLIJUbhVE
vglUp+awngE1qpxa9v3g5z3zRW2PyAHUoY7ks62OItuNFsmSMIHtOs5emA92mQ9B
6L2H4QU++poDN2R/13IE6E+8kBKby+BkYh77owarP4kFuKcGQIU/y2Fa9FOx7b2M
SPJfd7n+/xJs3iRn2VZZK4JzqRi58eVCCpi3CWx3IerHqZVf19nVzYby8EwVQvZW
zPE7tomUya0u6xPm5pyvD3YJk1GA15+NEbTd7vger84B6Ny2rVWTyEGRKni2RR5y
caC4wWdXBIzRt2ZEGMB++z0irqBa4Lgu1nY+LC5VdPB14eJYLdXg005AObT1h+g9
VnLIZ11DJg/Psm5SMcK4TxY7HKFgppzPoeUozVnE3HNP4p2d2jTPIGNlHkdVao7U
LjK76RUN9i8hO8pXldYxxtTgi2/OItk0TIKsMu6Ebu8gnwNEBw3TkmmuomX+h5sD
dJ8/thOtozYHPQo3PL6DBQ8pgYhp2gTOkN2qFD8f/8XIsPBkmFz2ntgpSTZBRUfw
9xQxkOi+CWKfhSb8NfLdKgJDGegNaanKTt3JziVElurlOsLZo1cFTSVoQql6lJN2
8P2wCRJuNJ7b7Ic4HjueJ7Isjhc7nwkSn+XZTZuxfKTZmugfdTsTbUM37rMWidKQ
o6xR49B7ifu3tzDu97OoklcTLrbwdymrbGkLcsi+4Xn30N23th02F6gGmd0IbS+I
scrwG/yhTdzygZ7HyPG5+H+CDnRdaXJWtn1gtMt/n0+Vf8zNRxuyOXvXa03195oi
STRkrNO19YMUKc436hHzNJ5xCdOnAPcT2Zl1K9n7YWokfdt0qvlkn2G+z7Gho2E6
wnNpwA0PSPQX2SOgLgiGfRMFI/fIXPy+twktCivDl9MNuAV3pFWwb4j9MHP3bydh
F7xOqBiMsH5hOUgRpbgTCpg5tyRH7S50Nws86BmYUTigQDOpiGoSZ+ZeAnAJZqiX
oV6+Pp9F5sxJI0IExhYiOxKYM4KZETR/WWaM/LxqMsujNFYpP/QAYos/ThIrooDq
wAAY+XJRwIdqbmoXTmmR1s4ogoP1T5GjaSMRugWUXObVRvAoOHEppSg6+5s9stbk
r/PdJt00wTTQSW2+NB/3EqI/tExZ3mwHOn4cQT4tiZXnO+S2XhJvpe1/ENAmhgUv
XsX2jixjPvDpsIz7jjLfrRymf5XY5eWKXY3lc2VNZdEXutxZY/VrRUbE4dWUrxfP
9aZt3AR1m9qDJ+zdp0lJ9M38+OYlB1h7bfbR6y6R5ZIUv5JqhxJDPOYFw9TrSczM
vYauTqfY6Zun04ur0/hjBHrptFYhbe5tJ1cZSGO3DKL14uw8yYM5io5pMPyYG95l
lNUuK4jEZkmeYQ9F8t6e7DfputDu50s0c/KYbyrcqLB+yS2AEWoMl8pPx/SVW5q3
VXwxYYybuTwRXUcNsaQIbCxRjlP4l8/Z9QKHobrQRRUJGTLSDYh/CA17IelWhYxh
Nj6Qix9IvGhJcnBExlb2kwbT/V/VuhMjo62enpm3pZMYfOcFL+Wtf3POgtAkyhHu
S37tTO0NVn03hta0CrKDUILzkyppszNgbOJkrsqLjW9irQ7VHPKXoeIcn+XB0nLF
aCJ5vubywU2bjejYjis7xpweU//PniGPjZqGUkZvGORaC61BgtMFfgipVtrer4tv
yJRpZ6z3pxuRSIihKs2Rtwk/nKq5Wnlp6wf4IDEgRCk6Qp49QxS+aQkgaiXoJjjl
blGzDMm5wN6R2YQUHzdyZrhbKjAWkvLkIciIBYm3K/E0Cit8eHE9y+h/OaLiT1Nh
rUyLhd6cxACXdO+LA7w1uY5ODxSYt9sraZ+PjbhO+iQ7awINOyJ9BmHlGNQ7xZYe
3LaEOTNYjZfwqzvEgCr5y7J2oxiVrSf5jEyoYobt+iO1DDNEGYlj6v4U/dh5NJzg
MmSYRNei9dYcG3YYhAqapk99eSkA9M5SFPn1KQ45f3E3MJH1Mw6WiQUqf7loWkI2
USgMuRD6BuUWk+S7Z3fgIKWxir391CdaC6bApMF/GctwVz3H0kFuh6L+5mW63pS2
Sx0KxADm0/xowDY5rCd/T4BXbd6DhfA5U6AoJUdPFIfta0oCAAEQTVFPp3PkY5F8
6nWQbJcY0F7ddryXlh7RFUbIq7+wpGcaLX136CaH04Nq5/4iHvfpZftQpKDgDhYP
xXIiCIZ5WHW7Irv5Pa+7vewkQijIOkvuVWsKtgArFoZgktaauOTa6/Lxe5Gwv2pv
SWiqQGzIyRFGGJqSHcq7A3Cl1lgbqmMyk2m67snzZeKs3LPLnKGf/DaQNdT9/97V
yds6L1OdFjfFeX/3De9wlR+JlmXg4AyRZ+DGdVUJE76e6yS2G2ijbM1cjTNOkq1g
qMms/Tqq/TPUSha98WOb6chPuh/KdiER0MIGz3S48sQcZn3N3zRFJq55sd1E2SDF
IWituaB8kXmZFO3l+tdRu9qr1/XEEcBKhh9pSUn+O5TmfX1+mEspnsdyt13FIH/v
HuNPzkajMHtdEn17ukeJVu6SS1altg7o3oucLOtVrSDLSE4RjWB3du5f8XnoL0gP
im/MLhQdFJM1mnvEgdQvfuMrM0xssk5C8u/W8B/x30Y2wVOXC57m2rJIVcBFgEwZ
wrgcbjmFllF84eRS95zGbBDGmL+kOcZwQWbEi6JhQHdjw/FfnIugOfYc28OSmezT
un4gCAqEe/N+kx3fXVH4otYGZ7wQGBhrzvL7DRmiUQxl6MOiY02kwWhvEcKGSmWP
qbZVIS2ylyHzfudJ2nzmScDg6U8F0gH4GhJ25hVZeAXnw8ANdsAXMPx7Q0pFS7Ub
IBsQAwffTx2XdOkD/KY3A2ZW0rmzrMXpPdgfbR4Am80iLWWqeTQ0w6cm1yWO64Hy
luCTlzXs10X9afuLLQFUVJ5A6SVZ4TMMGF5jipY2gbXWwu1BDZ1QN9WHh5iVvLrv
Q3BYlA5z3lIhL75A+QCWT0CamjyOb0RivT4edx8k8AEBRSLw4uFYzG1Vz/F3VubI
FNnb6VaT5QF0bUT94Lh7gK6jAMxpeyqOEFGMiC42srl4BVNGJf5HIAV/HJQF2yHG
4aCju3Skx3eLi2hEKscHGRUDd5D5sZhhRosJPPjk6TRN1sUNOyg2SIxCt1oqcjX2
QNIhc0yAPm0hWt77i8Np6Ei6R+GIDzPG1I5EQZtSucQXgQXJMyu6MmZYfBc4DJy5
aKDlzTKRdJULQA7CIGTUNH2PFw9xr0mQQb3CRqy7mkDv4Ba0k1mxWyp2Ch5+ELfa
PMrVp1SwTRsUp2N7QXtSI1KILixRZ2ZWcURrCX1Sn04JZ99d45iHiAXgqK92e/CK
NKhLocZp0xpOoviMekx0J32yh8NMc0nlNJKNPVQvW0fdn24CCX2wRYfhGfSbehsZ
NY5ZALAj/PxDAESyrPrawLBDYi7jOFLI9Qap+9eEH8jQN3i/QwPgnSyMqroBSucI
6zRT3pfrvajttwt7JPWF+TDIIqEwT49fPTE4mXYWTm/Da9P5gvjTxN/4PUfu/meE
uM4lyl4GTeixOKGCMWfltY9ctV12+5oxtzzWS2tnplOW9UfwxoE5RHIXkUwnEplk
q0g4WNuLAMqilVQSLagq8T57O4bUM47d6F30bT4qBEt5W2KUsjRs1MElnmv8YLtx
kXi9rMUxUV9EMleESAJi6Vy2sJswE32NPGGynBMi3unbS9akr9a05NPOF41DVPDt
AgE/xwJ6vceF89/C/12RUjM+j+tORhsXrRaagvjjoPaO5BCNuc3X++/lN9Zz3nRE
CDCpUo/GZsf4v3O4hVCnEWAmYaI06SoWgJkQeVpAPHm9B53Gq+f1ShXdw0TcERPU
kf9uJns0Skx2sCQtsGoEV+R4dCN0gFnOsa/tyCyjoA+sETJoIZyY8T5FE4ddf6Kw
iatEonpSYj+vhZaVAsnsc0d8g9+//a0yLtKPADyY6o0neB5moUDLSSNr5gYxQ9dE
1nVG+d1lLoEdPNPEzZhaXF5DINdeckNFjAPMIAmuNQEnN6XNm5AFpmuRKhl06FUp
uj1GyS4GylP94Lz1SFTz3LZEiWEyYOIkZ85HsQQfRSz9O4UQ7xg4qEde6AIf+rLf
fAmUErvRILC4Ngnw25XrD0RAggSvzNGIlZ8lqkjx5F7//mdItLwhLGfl0LJUx+8C
09gbQmEzOg+5ofclObFCxG7VhPeJb03kYLBO6bAtfSTFe5DCDQAPpkrYuokOUc18
WThi+DyJC1g09e3WgMuMth2jDvwO4fl+wDcVP8ZNd20bik0MIWwAl2PfhHB04i0D
fJMzykNL6mLtypSIeHGOAWZf7K8zbMFeW15Nvq1CSh1sICfSjOzFuhyNL+Ch/elp
aRA/eiYVkuZ/Rb/i6zbnoWr5fnLnB7j8mCBbiqm2ius2pR0+quk3YWdV1ZQI/CU7
v7CPYh+zcsRsViObUlXHunjl6h6XCT64SRBBlCKiYK3mmIRmxRZ1jTEcbC9FsUF5
6GPRFx81BM+Qld8fqEV5GKT0cSlaYdyNeWR0/gEgY5gQZaF83o2D+3vKsMz1a6fJ
DQd2povNYXVPs/sjFs6nWxHfJF7DZZLcIlTb7PVjoLOWswDHsbBkm0XJXqpFw+YF
ytZoxHINopZvYqfKti/VxtLm/aAEzkJy14yn/1VrE6X6oAqh3O2QZdgq0rH5nSns
Ep/UKQe5fguNbwcXUwb8WLi/xodtvOkLswh8tEKoQlyRZnCmCbWYKRleYoJLjoas
DAMjikdP+CBrn8QsHzDgvJg1BUIhs3VOAt7DyPsKsPTlpR/HMS35Sc2UY8xoLhL9
7i8oi1YQY+qabUzHHRNYOdK1cmHSF7fgdBjvhE83QL6rCjBcH0VeOWHd8+b0sFTP
lSHuK3gkj+iANOK8iCCs4LEXoMAGAqDPhuv/R1uzmnlqsAti7kq+GutTS88gjoS9
sn5P4W4m9hMQyby106eOQKiMU8qR4WZGutUI7OdNkZC+56V1dZc+yqZ1ld3aWwKk
pBiSe+QG/fml3usByYnJOY2cWoRzhyt7BASRolg09LA75euUFO/Y76D+HqHttRfJ
Qus18jsg8kRQLjkjzADuWP3nXFgb5iXuhLAdTi7EXovCnZV9NGaMvoznuJX2pAv7
o7PBHCMven3tZC3Vjx5maIfHVkwdp2KU7AgYuatRhofuq/mbcDFyNeQlBOsDb24G
akO+WHWJfPms5P4XzkplN70bC18XltNd1aW8FbZaQDFR1yWZGk+3rJaw3yp2h5FB
wGgQWHCvdrWumlX0eixWdi5udv864AXkPvIFtVt1A18s62RLtbqRwH0qz6kRONpz
l8pN7ZfWEpxo0fN0tguLZB8dpO64mfIpgnhf+Sytzi2jvcNwUqsDW9cVJD7qkmWN
wTcUD+2vKMGvFn8xMG5fJtIaEPCIxu8DFLGzde6SqhR/V5jN8s6FlizlM7Xf5CJS
zGAVKP19ENLNG7iw01bIGdMAmplbXZlYoTnsrnwES5+Xb0N/j09QwqpZTNQMN2EL
kP9nDlsk8Gi02xnhcgSY+lEbi4vHRwpoSbRven+R42l3pEoLD+T9XYvcweih9VTj
BGei2UxtoSDiH0p9L4d+XM6dz3qLOG2lhbsPVgmQBX6VC4VbuodnK10h3/DojxCr
p56qCwhT6msCpBacWKSyyuVl2+6EZRx19CwLJAZnq+zWNukSUr3PrBMnmNqm08EN
0HYWPmGCkO1GLhaeSeSDNF+W5GR/mgZqxID3Ah5uCiJqgQ174oOjiYWkNSr+Om1B
Vc/FY8YOBnZgYanBqhMaSoTAPc8ULrLFkwUrNFs9pixKUop1sFKdoOnUQS+4ViuT
hieh3IPe8+/QQLQwrNymBohqn9L7xnXHWMe5rpK28ZwWfhUu2VFe42C3dE9o23aR
pf2w2UTQh4QdHmDeA3xta/UqlatrdP1LYoFAlxbeaOfgYv1+Wjfq2S6e7V5ONHiU
yR6hEgb7ct8ha83sFazRD4aCJrc3bG0ypnJRZ8a7oE7VwWatjwWDyUqXW24wJVSb
/7s1RZ5/rphCFfoWhxGt7e4Yz+G3mqPvPXkZd8TQjSBxBD5fSKyqk9MD6OtyKw97
XHhrczvympDdvhLfJ+DFH8CPp4k9s0Rp9dbGhQbSGZ7+efp2Gvp2XLWEB5GwNNif
13QTxM0Xm3ADqVewMGoOLPIX1eLl02Uev860AyJ3nr/cW5QEFo5DotFTGGKI4ZLp
Do+H11yCsiie+Ohp7HRUzD7pMJHfAnpy+0hU86pcPX7TwUudiZRgrb5CNaeO8pI4
f6ZK5MWq8VRC3xjAU8L/jTpH7kbJTckOiNHrjuLhF5f1pnY6pxZMyjpmiAFa1/aL
BvN+iGym3CWedEl7HXo1NvxyCxUM0fPIDAnW8OAs4+VZmYtI+DqJQoK7FjFPLv/l
chfp1ONRDF247lxngsK7Uku+qyA5iGvjkqdlyILwnZnVMPSILZ68oFLfSSq5dU8o
Tk4h77Rz+NBrvRbXHTLDXVS82QEiPHP61CVQXkCGqvdbOxvlZKghlVqY7C6DAF6y
I2X1bypL0qgTT1L868uq2pY7Uhz3ekA4Ng0k1N3siFcgBb2u8ZAv9jygLlMznGx4
o5o/hsRl4d+OZPjRMV9TOWR2HKmBVAE/2jW1qaQmrjBJx+xazr7yZhmufjFcdxdG
ynOLb93rPXS8zdV2tCQw6ck+gumG9eQFdnoyHhX9tNgGzEulAp3balb8/Fks1CgQ
XV6h5WbitvPfWXidH8YMGm0tDI9wyuSMGJgf/1CjYKBF9zl+AING2evET0RjRite
8Zgz0FV5MkUIhyNnfOEx+Prgm2xGSk4RfxcU0g/hPFU2x71EangcxUt7+FI/m1dI
Mx823CoWVNFOJL5hWXlv8l1setULlXvPz9SICIQl7syappvkK1E34Gdjt3vVU6xk
iO+R/qQWArk/es+mHkTfjWS7kd+2mQyzZO+nTRzHRV2lSa/VZBttFnEYayqvD5Qj
ZAvb8oqtACMJT664oSQ+yzQpPjkHZnY5ORZIUvX7l1dG5N1DPBpHTT72hB+kVpZh
503/fDeEA/qbDWYW13yUzWuPM7b9rJpoXEVZ3cr70yzJ/DWwmYDcEX+DLAn6yDTi
AD24wpqjUU5miM0umXielAAUQ4KuZ2tDNmuTfqQKYthhPdRIXRLN2GmwkWBFdx7c
ko2ZUfXIpXWCHqfH6DrJUOcT2f0m1NaXf2ZS2GicRfkvxB6TuyXD9q1X+qqnVIUj
Hj6zxFAndGSnvzVgVReMBqUgBDXYryNNb5g77EDiZTSwU6fkzxq5YcAasimU7U/5
lCX7+RhZCOvI061r2sTP02h9MUhYzm1iS32t0WOLMTzy06yCFCPjDp3Rn4tkGRN+
4WXafmo22fS/NxEEaHX1YJKO/yEiRSN4EA7ZkAQxHHudPLd6DVvk51mnXn7uYH09
DOXtlDzyLy2AMKYhSYPTUfYr5gqfAessFkN1GwLyABUVqAV96foEHimuIS+t6rMn
921XjYKSFgv7o6jRQf0cgWX8XudleWjXOze97s5aUou5Jz7xbtiNvL4/++1VfepJ
uBY8Y6MHceTS8e0hIljuyNgK08iG0PTtdrNbAO8oZ+V5Y9iX3ork9g/FFNW/3a8n
kO2EKcx40WITIOYsPzQtzynQbrWwb2sNzrjTQ9n1CkTejhnUAdvaJCG4rrN4j1tT
b3OOo9Je6KA+xT+S9Js8GCq2lgSR9ibTdTma1BtQLmHDZ1YQ8F0POI6ql4+0zZJ3
/vyHZIr8YBmu/ZI/uTNe1aY0TkJST6bSrwm7f+M3zqEzrv7yJMTfXOkPDF13Jud/
lmaTKoL471aTMR6thap3EpPudwIBpALXrZXU1baaq+F9klkRWYUgLv4kxlWlPXOq
C6kIVh8aOqBejTBSQaZbjTv0ITUoabr2yl3LnCd2T9g1uS5BB017Ou++0XvjNkLm
N3tncxB5DOERRt5C+ODBUPvGHPMLQi3ECt9KLsQvdvmneIhuiBqIi1/z++JbDqbE
hZBd3aKa4rXMW7NtPFEln8F14XHgmqvI4Al8gvt/lxoTXq/3gaHmRHAGbqXsoT98
UbawLiWNwN0UeVKgqPouyOGOelrOYYH9Saq72ClptguKhqF937dwqbPiT9UmEQTG
XFGAIhkVhLLcXdz7feBcpj2y/7heb4rmc7qQArvQC1NsfR3889svt71fzEBRwhrY
tbhjtnMpH5AMBO1gzWZCtwEa3gYD1fPLgshLC8ggW7pkK/4eqJaBvj/ZmaEVwFt/
ihtCCWxAmBIw75XiEjXCpN2o2ul+s7IdTyV5fbnSpOetHYI+G9rMk/LU/a0UqCPS
2UdqiJBB+aTPqAe9vTEdHt+6FnWzuUtD+VjwWRMHlc6bJV6+SxFnqpWgrj9r8rQg
tG1V2RfQbr+874jdi0sYQN8bOzDZzZ63Nr+2E0ik2P21pYFhuatkwWqbAD4UjwGW
H2h8e4KrpaQo9bbjjn/z3GZ3SHsmBZYtj6lfDkGNV0tqaC5JNaYjFUKb1WwuQyTa
PXq70ikL1wRdbqa35fMdFbV3SRkC1BsQsOp2V1tdqncNgkR4ID0+ny9WmvGxgpTL
I5+bn6rszo46sPq2PBzgM8sNJkU2WlpWs5X2UmR9TTVB6B5oXFjfGMXYzpZTTzbK
3egEV7OftV61MIcFENjgT/uygsjlOfxWJjc6fsQoTH7OzrwrnTlGXN79j0BPDdD/
NXq6EkqICJ4G5s1o0sDeSU0ZE/92wqdTQTgzQVX9IwpKNWdidayfxk7xAW7djQ+g
xZ1Y9UuIDnMamtUbpFjEfppWCS0ziX2vG/c3IpItrC9CIttLynx8QXRS580c7wI9
KUsJ/h+xM6PaFZ5ZekMKw+PP9vHG/6iE94GW3mGQ4no7RzWL9iUSqixGXVovDdL2
+UpKBwvovcYYcYi0bXKab+LCbGlppqJT/5M0ebBBB0i7G6cE6/cK0W0AJiB3CBQK
kc4itNv5uHC4vzq+dfI631vzROT2LkpcefZ/PnCCBem2Ce5n17fbDntzCeGHL78e
N/Gs9JPYEHomVQw49Q1pGhJslX28E+E19RTSOgaolTgNQ9lzmy4RJ2LBL5aEFunt
cvlXX8fg4Dl9/gKP1V6a3eKvmgz55hM1vlOpMkdZHdCQTzdreY5Moz9IKhrSKpgs
BhnFN2nChWAjjiYH41Jvb2O0vJmvXI1LwwrSrIQxUmFPrlh/VFvamIQaY7U1qkaq
fRM2h0/zNxKXqQUGfiMpzSow6spUyCkVub8t/FfULHHX21AHHBfDrX04BRxL8PtH
4Zl/60RAs8mJw9am2DU80+JsuKjjwVx2PE7HwYTD5gim+1g5fBU6/fOx6ghH1rNj
YWG71tj15zsYrAfpFXBIRcYIP70FPR+dzEoEIAicEdpcgMQQRKf3dC9Ahvs5X8y4
Csa11nRR3pSI9QhaJfyatPnl9kmEtn7+ttNWwQhmsOJDxBznY2FT3h2cIBMnHxOK
gBIjVpeeQTVWM/OXWX+hBh6iFgYlN/YTm9nEbszCWLuM/1uezrkRlWMfmrCDFClA
NzpPjPwemDINIQMk4ZlXadQo9q/GX5PgSyf41nO19FVjJPJ7pXvYW/g9DZusaeg1
G0XLThAg+31F57z0idOM6u+jQHlNE8b7POs0r1rk34iOPG3PNzkwsX95UHVgqziK
+ddhproAlTKhw9JFWK7djgWUJ2J49/RGwgtDnHPUWeKJA4jBCeuWLK9VjEsN+4GM
zNrACmTtX9wjelUTWyfB8U80KefH8oXj4Mv9U+oHZFex70J9f46HSaVjnkrjMxWz
oHqDiDH19VJ//6UGqNHtYBKQZjqxZipdNMUtneu0fZDnutRl6JYpDhykXHrZTVyZ
0QLqhkHdV545Zp0h/FIIzLLrLeVqh3c0XaVc7bY/h+F8RQocdFfHVXo5C/eBkZyL
/tAbbrNbRDYXj1mKr5fMaOmaxaQIZHs94nYXZfhKEw63XPYRgPmCuxNkiMBBuSlG
ovsM0eqWLSZCiu56jNT/eHe4G8j5UtLsfADuUiITrkgOoxGIpGMMbmySjwNBEk2o
vyuabrOKslCxqKv0r+spvCOfidKQ3af/GNGbxTXZo2k8Ws7gEIVG+V324HbzE7ba
PJWc6O8UdGppPqvhGd3seeYq0Ni39cJqlkVaSEuDIRnBR52oAN3oPMeJWQHo4zhe
+/DnC0eX25iQyjxTF/Rx7ZqQ2pgCjMy1sCtg44zbB7Og2jTAWS+LhcD/Yax3Tnig
HnG5GRj2nwb6N40exiDZT0G2kt6PiI3yZFgOjr5aTJ/aWtyVPRmXdLzt237TdVJk
nM/+PEAerFXd2yXatkycTYfq25W4MeEVR2+S5g8a2Ayk02IpP84MZKsFlWcqHYGQ
LlxmW5EKPlw23Tr6N63hDxDpGvjXgwHnYkDXnFt5UkMI9V3eQY3WoLc31cnxUxGe
t97xrW/UlmgtfwJ73F38k/lBIVzY+8VLkp+plsrqUftPOhsJocDwuUVxUQAaq6f5
ZC0az2oFktrsbVJ0d/HGQBtyhCgn3hpL84HYoRsmK+zhKXeFrrqwKbqcFDyrBOJ0
c8Dt8IsJFl0QqEdSV+QA0G2GY+MuMhZlGbvEl81lLRvY63r0gTiTNj5yGzSW3K4v
eGS6366o0qQ2DDdrg6metkBkN+O1nRnrhjy1Av1oMZDA8A1Nxi+7ao/YFiA33aMY
wOnB/1DZ4MKBupYle1wB7Q2BOOIdENMz2TtTKBcXINaK31S2vJkWgH6LOmcCCmf8
gxAG57pWz4gpNjX939c2j8CnuEeqjExnVU4ZCpviEIPflxkz5IvlzO5pUG1kG7uO
x0G/SkuW78q1ZxTLfTNXQdZeBtUtmGF9rTuBkRAQFxJ/PE5mFOLpP3DMPPYH3lBY
vPtPPbrT8Aqnk8FWokoz8FDWPClcAwiyfAgVy9Ou/lgLBd73e1zKg5uYV+8VY8DI
nwIQXn5jPXRuchbEvAq74iAp5bz02AgZRyJiZIfvkK8SK8XA6vSD4ZzjfWhfyUTZ
ECjrumXDg5PrOm07OfPhX+FuRFPLPQtMUrivqk0mxg3pwwifgDTiOHsQ9prViTRL
a0f+1ro1PGbDqitU8CL1m9jgz1ETO5p4rcZiPIYH50bZ22Z/bR5Nu+4G21VBqfib
CRbhboGFMG+z65dwlhpeMdfvKCAtP6iX3/SEJph4TuEkCVI8m9GEBn/BLOrulhK2
yprEk/Qh2yX53oNmhWQNXNL7HPPu/5zLF+QcPtXJjey6XN1EM6kBLGsK5vNNuRdl
Rm/iP5FDk8QUmJ48O9Q8V94td4H7YzBV2usQ+CYcGzxeKJiEluRay+Twod8ieH5u
GGDlsfkK4myJnz1U3ZIxRzX8V5aIt0Kl2Nh7FlREDG6MEUJTrolauAPGclqyXFju
Zqm9M/Dqli7kwUYVJwjh1kWYa4/xQTAJsMr5vo66AVT/Nz4SbuRsVcdMzLRQjeYc
0EOSaqrDn53rnCE7zc+OxgYG/kmzaHjKrbCjtNvh4hKCLowZK6w3bXETXIeE2bV4
DYqHnYUu78BIzAPirCuIVQgYrF/muAOL8JZqKzo8qr1oxoiOU+AWS3DQxsHmsIjJ
qKsV8CkV90O0E4b0Q8KvklhlCvkwSu6yslKNZUISsb1ZZL42AtlXUCgF7VH+3+jJ
bNNuXhrgxInU/lWHq6YgCpyUccYU1fbNvqvNt3k2G2/0PchZ3BwhozCK0oIh7pkS
smhz+SZ8D/ejWgb1xFbo1JK+8pksaz0krmYZv/B/73HzVaBSbZWO7jv2/LIpSe64
JDifh1JzQe8CeOeu+ikoAQ4ZlLOyvF5igkYO6nKdIFlZg71ziGjmwd9riX8J76aI
y2Ku/RsezCuGdweSNiykcQ+9Yid27TNf338zMpir1JcGWs+huYQTDzaf5KxZv9UQ
Gs+/AatHDjZFhqFX8BII9/h45A5yehdgpVGsu6Y12xuxmLtvzCeH437qZLjzHiMm
RfjNyx0r7lkHMxlvdUvvMWn3+/0SFSN2FbOFswMZ/p4zpiJ+gx11LFj7X4BIxsUK
n2c3EtAIpFZrb/8ZICVVLAG6rzDicXbYd8BH2TwTtbMWgR4mrhI6smFD/J8mkX/3
T6/uc3X4BGu98WHXf1jrqihKvOjkyVkJgr9vlKCyMglP70ksDpqb+8i46it0bpox
L702qEoCqhvYzJ53K6+zUJ4/z7n3FfIJD2CanP8cj32lXa46D22ZAnLdinvC5fz2
tax475LC2HlmbjMLWeBEjwaOMVH0PAEKd4H6A12Y0bqcHAV4NXXKuPW1nUlTCAZa
HacTMl4IOMdgjBNerRjSZTkK6vcITvlgyfPMAQ+ynfItk15Dm3ssLUAHKwQ1Y4lq
DdRmkBCQwETpRhtx3WYRwwxSy5YSM9MfG5dqVsVyvQs62RmSFS3I6q64W0c+NEp+
bQht6Ac9hXGIZXwrO7kbhQwM+NZJkLyb6aRZKc/p7KpsEhWaQQOyrj8kKAQ5fgWX
Ag1WFi1NB5GrgL8Kb1xBYNQXzuGBHBQJxtMpewYgfjye/vdHqjLhtZp4as34bazN
4eM8oJP+5tbs7TMIRMyy9fTovs97QY5vr/+Hns0hG4dZw9FJXBEX4DWnun3++OXr
BT1CgBNG3oqqEBjIfVZPgWMAW3dVQ87Rd87F67ZeAgBj7V3hzCLYJvpUsNVDttMo
/EKRUTZfodstjd3b0sCu9u8roHpmXu+gA3idvhgtxODgq0L4xzEKXDbdLWwydZdI
QbJTk2SUyR3snllXsR3UEJ8oR43XAe+7Gx+NQZMian/K3RQRkN5n9RvLmF/nuE6d
wPXb8SLP0CyWP4S16+AUQ9bC98uBql47ThN7aUbJAzNXmEVyinp5GN/wmRP6AL3X
7yIei+Kl3QACVJCLUn41+gSXBCMTOUr98rLcRUqzG7eFBtPA+9WpaNbt2NktYOsm
0o3sTRbNyit2RikCmflm/aHaq8sP62CF+yXWq30ZjQCrpMrqpqtO4tgSwB9FjhcS
MY9foOqBo1BQrGF4nSvXhY4Q9xZCf2Z9SnM7WvyVQmm/KsJU3SOrcKTsqv3y0wOQ
Zjj6389cegMAMmOD82jNSrm+6axh9v+oUXVYWjCHXZnafYsMeC3DC7ocaOLqdvRy
meK3k9KYoyYb0PMG8RlzS5zCiAoVbhyf/PEulgHRkR4RwtI/KlVGhBsG8LmQ6Mvq
RFISLVKgsY3l/Elgn8/mBclO6K/p5mGFRBDInnQzafHae9BNBvX8Lxv2ge44vme0
AojljgJnzeeeSb4Op06xyZQ+mZGVWD+6Gx1utJ9BucGKr2/RGhjkBae7QaKQojv0
o5JwQ9Wgcj+sMtGh8EoRKF2jLHrj2/ilf/kVJlAlQiOR/u91HXfzrb9MiwbqA53p
EDGpmzmOsf/LPB7VzxR77ss+8AGhHRGE64AoQzml4YyGHfdfIX0fdtbf/+eLHFMb
zTG5iPkxc4LESeIVzhqJg15Zw2C3+4UdwfLDPhbUk7eufrTh4TRlaYgqfr0CzhOC
ls9mNmGZYNTj70HvG4MCbQhxBQql3Gl2ZMx6TcQoLNS4UOv9HDfuT4VpJeelOvIr
bB3kWaAHKlYU0aJ0uufCer74rWJ8SsKdVxn0Rt60Vap9TURCp0fsC61RdS8s435R
4BbxtG/g0LpeFQWqRQUIdlbQ8OJwD4K+Mu4Z+V9/6JKuaSkr3xgvCdCgASZrDXMt
8NlIwROr2R92MVGTYf2dsXbwUhcd8H143rbzKR7aOULUvesQQ0Z1ulooWv7jSu+j
90jRPQOO3QAxh+W1GyPOzZc9tEr/u65goqkY8SOkIXZdbmawRefu+Qvk1sicCzml
fkfREhYiroR+30yxpOgBXGzZF0o3xnDPg3yb6uX0rkagzIDI3yQgb+hosROkE4Xe
5o5PkP6jnvBE3hsv71TDLIlOgQqOFvBJJOoLVBGkb2DWZQ+HR3BOEGlRBaHSYT4J
kP9+b/6fm1ni23HxXPMC/vKnNBjGfxPZLfik8ihmyFapEGSGXmYWVlu9ZN1cyFyV
JAtrpyhxx0VW5NDULr1CXxKYY6qOt/l8BOBwJdDLkXOGY57LRWX3S6Kfih/ibdhK
PNpQyApOkI1skwmRhEaCxD1l6eXYS58rmr5qNEP+so+xtnKAKQE+kI7bcpRTBo4P
0LWvZyn6+Y2loKj8KFk99wv48yxkRsRsypzS6fsNWWWu8uf4QGGyJiCf9womvjzF
pWMa7CX9+98jFHYqn0SEtsT6Oyo3I3tIeAoCui4Ed1BaGK9dgIFKEXxshj9wq2GD
W8n0OQUMNsnHA0Tcsi+ukns5244rfoW+I4hcU/hM1hRXKuEgGMW3mCWCirTvTzRp
3zQ3OZmKUq3yTvRMqU2qk6QgUBdjQeEh8DLpeH8bgZFAup+YTMprOafoAFX7oEfr
7CbC7mt5l6Wv0Bt3ZsKdWds2A7GzN1+GylOx81tyktNy3WlYlW6qgmzvAZzDByxJ
+YC8rCfiRL0uuqSPCpZrA/UBYdDyanWx2R/DkusBq64nDnXhhvH0aku3rtFKFS7p
r+2JCCutQNMeOSRrP+JI7VZkgxpBi6at1TLWyGbpuKYLCRrqgePLlzW8TbQsNOSc
A3ds/kgFPG8mflqzTLtHbo+ZVYE56FAWaN3O1QLBq9I02+nWmOZerDHI/yBs3NiW
tRKKidzsnmCCau33pajHfpO+QkEqh5LHFkuqFv1oG121Brq/eQL2DjGDpq7KUAeu
QD6/7R9jm+HH9M7B5txLl8d8Uh1JkvbZDj0V+ABt9QjBZxM7bEiDNTx4fMWohHYt
+DGWO9Zs17fTIPhr0qSUvkjm/oxLnzmpxC4gyaCCLY+SW6BACdsvpfd9gOmNG2AN
jkt17ve/5Nii7Iv/lnpcdud2xsDy1ruSY+9trZBwQHvhv3v++SWXRA7cGmN5GRXV
ycrrcAMezwVWl7Ry6WRqIP4XnGscVIqAGCyvLML6m7cEHWqtaXNJWJbzX0wpQBQ3
rAbI0DrWPVw3bpOXK+6ERkjn76NjBdQrbvNUBvyVEnnCnO0bP/+vL8hYS4GGLt/R
qygg+UDAWsJiYWtayv3uFvKC4E/r1fAyGEtrINoNolUqKPwn039LKK1oHDyPLmfF
tsfIrMtVpnJHN83xC97KPzknXzSogRiwAa9oJ6V8UUuwaia6CZjvdvHSvWPzO42Y
d/h3p2Wj8r0itfBVL5Jw/i1kXwMm4T7+QOhFt9+XFJnRbMcjE58YOXMwviQPSE3I
a2ED6TMzwRLK2GgwuNFXqGy2r0WqsnrRV+MiasyZLKBKl+Yr7zZYtr3ojaZlN3ne
BexzuZN8qodTn6qBIIYbu2jdbJGQE9LYVzHpxMJZ3Q8fShSmDqcSBphlyEjaBctn
SrYG5WQxMg6/bPJMAIL1Xm6FStiWzYPZKIYstXG+a3x0A0c7AymZQfkGOuTNJzOb
nIzDWtcFLc7AsOTlR0TSs2LsaIfmMrM378mlPPeb7+ciEEtgcbxkTDMgPgvIepNk
1E2bgJowvUecVLJfSUHJh1dlr2wyrbqmg/msgX+MruK54Z6jAq1P3OOUueGLEHOA
+VqKPcWn9CCVxS0Kg0X4MSOTgKPJ+gixai8iub8wZ+vjSAa7sVDkw0SrAUsUwcYI
TqHItxRWLJI2Gmj2NtsYyt/12FP2norSerwzscfc5ePMG5RoZDaNOHvcCxfnX/Ni
Fn6KYNfMvIJcA1kKsFahsfdamkTeF9BTNiGC25X9We30JykPCmf9xVaqBo4VZpad
TTTahLF75XDJ4KUYWqIjX3aYk27/2swo5aoqT7K87OxaR9zqt3IQCEXn1l/zbtPk
dQAiqjTQRShOg6pB8FSfyPc59Mjh50dGA5Yc+zNB2MlHu7XUuS/qD7K1yZKm7lbN
fdH5gvRlqryZXGK2EYLkrfxjegp5f9gKmeKQ9OFkwu9HcufOTJOuG1A/8LLAtRhM
u2G4gqox8RUs1xeHRjyIC4qhaT/Oo1iJqK2iN9aSOb9MmrOB5Uuk/y/QtyCjuXNJ
avElWyD/G66FfG9pEzqV7PGisSYv8A5ieqSOfShK6xZuOeWHGCKr2v9ncJeS+hv/
LPH5QRlQ/h6S4F3qr8ujBnE+KQHBMHTlg/mPD90fDUhYeTV1MKqnSsY32bVfV6DU
8k2BTxVvaUanM0fFgUJRaGz1kwVkFaPRkHWFX4sVTGWHi/QUkBnmHC7+dT8k46h8
1BWUX/+rzuYY3fFpf8oj0pzWBEgI6ya94UL4+ByUITpp9wRRc+UsPy2wD3Wa7TsP
Sc3x+6S5rNDPOTpPlTZ3rg+gGrCgTt2yey1BpEYloguk7xKwTshiZn8PzT3lA/mY
DAgOHbxrrzpWPZrW9AbOtpDR9/CSeagPwVCVXZ8K9tSPXNF5B9jwX6YzJzzU7UKo
P/V0jm5da9pCEfyshhZDSDqWn7kdRzhyDVnecp9TwWHW54cq2XaEtoZeKYs5NOo6
SHPpSeWCt+vDOR4fJFXYOIXXW9S7d0GotP53W5IbN5pUK7lZ4ewC0L5VVyg5lKx1
QTty1D2L4j9o++120jxGq/re5sPIrH77nsxGWo6Rj0p56mCyZdFOTv5FQpNBpQx2
n1znbxQAACIe1ALg9y+xMeaBe9wdk8nWJEbmES7Aemc1arEFIiXzLkK9cID0/CRa
dJoPgjtBpQImnBoQVlvP+hwKjXDbqxdDNl7dDxRSuzjbfENqm1OSLf3XVmzVkA6D
LQt1cOrjErNqo9Qg6jJDcmJnGAHMEYwAeWq3bpCo0FJYIzsjo5p702+/q3BCJo/u
vVjWezn9O4qHxAD5NDZ1mxMtrt1vqKECCAI2xgtVyD1N4mmDCRrAjx8q8KOlE3OW
+mBzMEWKPKlYnXhIb/RwigwKwIxHdIOZtDLZMCAf3nd03gUhv0IcPxepgb7sxF/H
g1Zam+Yvdb15kUofSx/d+8FOXujdPtHpuGumPncsyEVV8bDG6FtNdlSHGvggm3pe
a/6bYhIRf4cDIiHYy7QsN8KHwjy9Z1/mzQDgxuuWKq9MiBjamwoc/Nwpr0BoIq+J
LMPfwogFfB0UbB0vFVUup0oFKSeT7CMdbxBd7HBvPRnDVeXYIb+19jbA2iyn7Sn4
oXx8o6r3nhyij1Ad0Rw5Dyx+8YjC6/m7Xfu8WpvlmpRY9jN0Svs+7aL48OAldt5Y
jAPZ8Bhrx59tqL5t6oGgMTVvNjORwqDQNNS4ydd8qGKGNUnSpgcNVetug42tspXV
/tuSg/ZPgPN20iuUrDdqKB+PbezT1rJ57FsBk6WRAEsTia8UWCjVSaEjefYcxgqh
LoJNkBLQZ8GTsai3yHxAh59TZeRQKpXAWNZLfplFphLyV6RXvgk44lGkqxW0W/N8
Mfb1ZlPFCRY0vUf5YQbDok6CiKHxBMc2Tp0cnXgUgYUJzRLKhgeOLuWrNml6y8fd
sghPGmlP6hUCmeZsLz8oZX3b7w/cknYxckg5+HVTz1BzLoH32kypaS2wzKVF3+uI
Dmx4pOFa/c+zg8XnlFamMEyhJe/STljvBZHVUVz8CghAG1MB2coz3K8Hio2t3T0L
5qSfDbbhpaKaAzYcCHC88lNgi5bqUhMMxCzAHGi9+lSWMP+6ojqqo5LHfNwpIkze
LGxkAdENdjLOXRKDwgcwPsvio+lihJxk6E+5Vt7kCamk6AR2rOuTjhISJ+ZD0DrW
BgwVtNr9C1WRlAMSCfWdlhM8S09FmwlG4Fmqy7u82cAhEU2eLlkO68HyaRYDDxZU
rV/HDI/ejmSSXt5/US29Mah+2MgqocwfQz1zITlk82lfCxzY9botRHYvpAZeimrK
xtPZlb5VPDA1gJnf7isPBm2aLRTF2jarUYx6QOu7kT3AfeBk9AxHOtROu7GCfkjA
PvRlwML68EWQx/53auQr/tRQueDmjfwJidlK4XT/g9e0abH6Q3D9IbvTRtKoSyHf
kiViYq9N270mJuncif9Y5WBiEDl7/bbFQ+Z44bkR+iyKwKeYfgP1FDPzz2p+SHJW
JbRTkBx/QY2NhPSDXb7qgKAJ9FB+B0T73lKnmYFu4W9MO0/oTZiImmuioCU5Ugj7
5VfWIcQXJjMQxVXQ/IFCgKGRFNj966PHxRM0reB90/dc0+O4YzDsuNz8ATk6b0fk
szDqCTNypKP5u9vpJvGdsQBYflyFtGc43FMz9huynfuHO5QN8hGmL3G2ebOKQ8RS
CrQ+PvGW3g6TiE4QbplNLbsjPgxOz8cWORck0InPyU0/yWdeg7ADbWIcKbVIXluJ
NOwHSFs7fVNdxVibFgEARJFcX+2Cy98PgRWMgd9C1FZaDZxLh5pnQVtTOOHAYSpd
eru22rl/zFiiBxAG1P+QyxM/MMHyFgGfQ+SOHruPMRJeT2hzNzKoOZdm6NTP1bEC
4WXZmtpWOjtBljHY3GvtkkZiW6V7ZuF3LE2byDlPtSMUNBcyhCE19nHYOTd9Bz+t
WkXeEj5LXSLT7XRuQYVxSaBdOgSfHQ0atlHYvzXX7YfNVFAmxbjIFryeCm+c4uL2
C+5bwZr+0/kESKCvOppQYoHPCI4r5xFIdwNDsrClJI50sQI5FaSI+HSzexej63dN
yBt4Bh4KLdpelwovr8hzubvJVTVIXGbn5+t2YwMSvXTCsIMRxCa9YamYmu3VsDjJ
0QGHEbde4MyqMWyMUXIyH9IpHefWdYq6DwqGT2AEN1AipxVfGAn3ApUQnd9BFlvr
ZVBEo0BZ7bZJPikUb17vxqAv2LwtVxnOMTXQLOWqlAaTBDNqAT3kzYIb/SN5wMwP
jpOcQefEa+cN8SNo2iM6bMwdG8WCYXJCo8wIPmcW9RahMOpZJk9v0M5NXD8+b1KH
R2sYtFH38xOGtarO2tqnC6zh6Gv1MjPdbNQJ42xUKps03Y7BVQmXMmAbIcSCr8zi
MJa5ltux6R0ZagjYPVjBq5zxCj6G0OfOsRoHUk3mJnt3+SWwXUSgkt5ik1h4j1yJ
9uFEzmKgX2yd3pPU8gnW4+JBaVryH+P5ubY+eUjzvbHnj/ozMDH9sGpx3LzAAATH
tNwPW24YowBtWiPwTE8Si8Q1ucgr4TCz6wTlCXYmMKlVRlvuWxpPu5pUA00z0J1r
w1hJcrPl4JJNEcACgZYqp3wLWX1EkG9KaIet4pZN0VRqgy/eaaFC6DnArQMcWj7g
PSLHmMw3rWT1WtkcQ9vKnHkG1+cX+5kkZYXxZWpY9o8eLIUvBBHu7jLjHlwmI6iX
b0PEG6baCQV31w5HU9GiMiTUG9SP+rR/3pbmVVj56gTmff7GmyEB/Oiwsq0g8wm/
d/oKnUExZ0++Lu9F3wPAIhLyuYCxbTt+5HP9pTWUHEsieLWaw+nlGU4vIJc77wIr
+zoy41n8tNPBVvCL9KbDRyNdtMzDn5pyafUjSlUhkwv8PEdQrtqnOX/gpwB7Vkdl
5FXbHq9y38fWqpVPsFU0OeKpgnkCxSJza+ElMs3vEKp7ou+oeoVZn53xysTX3HTC
65Xi3LAwv5KaDUTtWS88gID5Wd19yRTuFpUc2OMJXVz8y4iZVIpdJWUN2U0v0GcO
Gu5b9wu6HIAePc/L+4P6hKJlmbiLYtZpTdvEVB/ltwqVbJnHSDr+RQ1C9IrSFeGb
1GzjNsl2d4WLTyccKZYMrA+oUMi+tYS9ExM1gPsWYXfTEQwJo6Ups0wskN1VQjuD
FVH2LnR+BRiLOxJ8HHW68wGBLGJROHHFFI/nxXVQduMOuYFQ/qinX+jZBdCB9mco
ZrMM5JofDVsnNW0khoB2L0iVfY5opL6raxHRhlerurkAEF6oXOlzz5eJr+UrRl0c
0s3rd7y9wmlayuYme/uvJ73HKC2TkQnMYA6Y9zOxNqsj9h2aHq54GP8OOSEJBXLf
8OuE0VySuf/vuQMjzDjxseQiH3RSmGher3PouC0wKQLBFnA9boxcmYK3u9/PW9+e
C/Sk6Jed6INBb6OsNoq1Zpm7vkX0w6dWyPWEM79S4wzMDth7rDn+yL7A97UqLl05
Gsub1sX6yJQdgHkqmWq8nd9i2TGq81ZYmAumrwIxo5V4R9EiQKxGTDDoPaNAXTZ7
hglBPI/OblAvlD4fM3PakzIl+y0wJCFHG6xlxAtAx+oM2QMMFvXRSzQtTpkKuaRt
kIhUXIYt4aAFv1mWAOOcW2Ta7N7y3M9D4/nKTRBOBD4aC+zEEkkKlrGFW/jxkkHv
Gt5JrThRxVNwkYusUPmnKMskgVIYnkz7V6cUVYhX+ZoOifobWf38q0Pziwd3wZvG
NLW2L7a8aQZwBG1kigsTffmhc8/a40JQo6sUkB2qmMfxPvN476aTyMeFtucWVHNR
/8sFtl+XODCSlEt0R/STjfe6oyD7uXksWAkQcN0NWgCOeI2FaE/2rbZVqVH4GTMf
15rCOEq9tlawD69Ywz1gchsNHbOMyPGi/Ry6lDlV1tXsOB+aciDGx3H0Pw0mpmxY
Es3Bbh1cJ0JHTOzikZyivSW6VLb0d/Sv9A4C3N4OG11K/rms/yYceH1WTLi5hwwM
92iTAT7xPTC3zWctRxiPIOaKxk6EUBoQi8PKnSwANPQ52cj0DB4PQkaoO0jKeAI3
00j4XrGGY83cyDhTEoY8AkhUSTy24ecGS5exQRc1BPxy4PMrI0dxKljaoWqH5fuu
VIP+TDNPq7YUmowwXccBlDRuA+SKW2BMWC102I3gK2r6jE6uCp1y5vnFfJ34uURk
BZHWi1oepkuUSdl/O4xLI0e27Xfvpix5LrUYvGniIizB3CxJ0IGmR0ojM5tWGbYC
erGBdnwQLRzUyOB44aTzWwmEvfnzL/sDAdx0Z0ZRuDmmkZKiWcDUv+mYT6VXgrsZ
vv9W0lq2xjo0jRX8HBhNgpumqRu8+W7WPK2aiHQVsSL27fFbWGkNC0n/5PlX85aa
EmATyzAmS7FEzqyEFDTncaPdAILpbsw9Fe620dvjWSr94xwkSVPTh7Wr6s0axHK1
HQB842OHA/2j32JHhOzJ5VqXOwb9ILeddByxuy5EAV4zoqEm+I0wsgFBHKaxzXSc
tXTtL+Q6jXw1u0eylOKhQhO3GenqCmpsYJFV4ECFDWeGpsaohntAdtV/VO7t/Yoc
3kPXPOSLTUc2dfNiu8N58TVERUT2Wm2nPsLOJbQxKWvoBJe/geQLGpAm0csqsRuK
h04DPOyUFLDE47kDrxEo1Z5ldyw4x4oXrRbMx7eASGyOnY9ZQrra8BrVwTlJ0q3E
LKwN7hORZAzr1oOsUpeC6bPKACnoQSU03CWVRjDXiS1duvPMnYqBx5mnBmm/HmZP
uYL6t+lQUUvQ8NdIqTRU86itQ7lgEhTgpQT8FCTkC9MGPVNa+ZAERQgLHYtraM7c
MJaiRWLAfACiuUBrm4DLtCj4Qob/TJrMKDSMuN5gihO0MhyVJpMjL25kmMdTV6Qx
nUpaXjE6SvwPCzMpXjsojcnTbcLEnxgi2lqedBFbrhWysGzl4DhSzKMSmQAb8CuK
3IGjIjccGZbNP3jLDARjj6Fcwjr8BwFOGJ4ll2NO+XxpTNxQQPpGyJtCGpdyW/tQ
n1SCtz1wOk4w1lJTO1X0YdELZYd/Wpb4tvLL7NJ41TW+GBKkiJnVxaN16HlY8ekO
VNyl/fYaDNdDR/DC1a9IiMsP+0bGmt02pnLTpqV1YVcE9IjFVyaXF/IbQwWM+wUq
9qNNLOzKHm2PGGReZ8bwNaIE2s/y7njIIyEa0/OXvnOpe4j1bgO0cmDEbC9Z1ICn
Gauq3AtS9nGSB1VXWX81GPiywwnPiB0nZ88IGiIG5rUP7KEHFw9g5YwXsHPoSbNz
aPo+JEgqYnteoxSSAygbC9/Wl8XEyTtleDskLfExKXdi8rttz6+rKv/QayYxDdp7
onsehCV7El/J+K34c3UtjWpWEemDYzE1wd26FJpg5eKqngCCr/slvUnh2QrXqle0
1zGGkuLb4dTaj9HHYVj1H8eJglieeRPajgFvJnUXbJVnW+i74HSW2I6lXxKIdsBv
oeyETEHxmf1GMwTfvrigB11QD3DpD8wKnxka+9XRhdlBcrDYI0OID6W1vjLgIlpd
HJb64g9tvgq1tnpv5lpdnuBr3tONcYwmt+EvVwEKf7Z89S5ad/qBZlk98GSI9Bez
koWTYC1xjwvFudNx8IQVerbALm+4SExd+kD7y1cZBgb4IiWd23dAFcBShmImjwk5
uOOipCW8xzzat8eUG0f+4KVkkdifhqweXfQYVMeqIHwc71Q9FH3PvRB4YwOguasZ
RJ8sER1X339yVxlJhVmlslvVQoR9jcQOvLLD0PirMkgu2NycBsyokYFAqEm1tprG
skgfB9tUSi/Zw9N+Ug544zNCeQJ79IGWq3ns3JwtfXUDXg2sXQAx8fzkZ9IDeUfR
vVB1ApPONDr2qTO9/4fwDgwlS07gTfbi+QAHzWReuVzcN5Jukq213Rj3Ed9bgCWy
Px9IVIrDb4jDu+cAv0O+kVS8jTSpqNlISmjOceKibYPwvOoJHzggHqxDzq+1E/pF
Dz/kW6HRxGbINEfVKLModX43njnpGUHiWMipmDn1HzzFc+5KIDuC+iY4xxcCfc2Y
OsEVbMABrnpnIqe4GdNDYmkhJ7ZzNBWIyMXatOoosn2iz9ux2TdwhYNJX0vj07Sq
Xc+w9lpPjP5/swuW9IL+vBNEh2Nhg55MVX1aOcQ4EZuREy/JF2QFNPqu+nIGIRQQ
E5Di/y5ZAamnnPSZDQla+l6hZKtCG1J3ZEgxvHOB0Oe23+eMvT+iq6GlsnjHFbuM
vG4PEhpl0L5Ji2nLJxrUPqtXXz/V2qnBa9VH5XM8BC4BKXuviet7O6fGlk/Md6Dq
WryHcaCtf7kdPQplRixTxbDRjrv8C3NeT9Vs969bfjFTYsQZSD7BvAcczPgz8Y93
EpwV8R0Dafr706tmtZnxDSmFfsd9/HDpHOQY/SP1u0AgdrxZmExv+vTPYCocNv6N
lCZo0nfrLWYNnKC3KwRiUKUW3MnLAZb6Fm0csDfzPnBDJx7FNXQ/qziss6Q4gHjD
z14P4uZj/SEWYtrXZ5cFdtdWZCK0IFO7LIBvt+i2QxTXCxrd/3U5Eqzlt8CO3J6K
Iq6yMEzTzQNgAMQJo3Uh0UlMfa5QcaUsrtu5yY34SSVVpD/6oV7ZMbj+Qby+jfd9
50kPIQDzC9rtJcHHDTw10CVEbLF0DORi/sCW1yPXds1K46y6oz8QsQLXpxIY63Dv
OryNNt2lIOy1gdkDyIHW6lyDPbsSkBM6qc+AU1g3S5QGMZ4ip4foLINrEuzjYkru
P1k6O/y8IGm/i0Iw/A4NizXM0kL8k3lawvyaDqilOfFWeLw81tR2vNMWqMQ5Bq11
+axBlfKjlrha+Tk4lnu9PvvPyHI2GKPkey3vSZYCnBUHykeb/Qs5Pnamm/ES72q/
mvCPClPe1KqJCXF3Vlfg+KCcgoybeAeCbUhYh9DPVHqTMXZEgoYqyxQOd9dDsUJ0
86y56izUsdjj71w4hPT27DsvUnCefHHbSGdN/OWgHEsYTSPKRwT15+oyXYi4sTJU
jiKXUsmP+WgF5ajCOmiBdbq3+7kjcGrZC9+mwLo0LHyNh+SZo6D8eYQcdHbhCWDu
WS53k88wsOVBGmPS7kkzkbb6c1eL7aWUVl3BjdngmGDPT8I1iyo/+NtvZV7BOge6
YUP1c5ACIa5CtrdjDyamAcrhHhbsB96zvlErW9bSOZfTUlzTENgJJhLoYZxL8qff
ipdwYBVM1SpTL5KOSmSsY3RBIFGSGaS4QSN1jOhgtrGGqYBV2XUu0yvthepRCSZE
bVvvE7G4ws3T7hYQ5sq8g+qkrK7rNrZ9GzmIoj13Jmf1A3pHjA2v4PrNZjuczz8o
qE5+5Rr1xbyukuLNth/40iCKaK1DXdHUM1g+tf4SqdGz4hfNbP2VX3u88/1NPZzI
wrP4/CiywL5+yN+leO3rP9TCYmXDQ/xNlq5N2aiph0QFy+eiHYjpGpJlqwgwlLRF
Z1K9KFPuY3Ev5MpGDr9xqJI58DNX38ko9RNSiKAlOult8wn4Si5SDvF2VkciuHlz
fkuGbmEKjhRm7J2blOzYxc9o1g774+cu25ubVBEnzK6ZNio2S+NvbCkT88ruJpnm
RSgnzNQvQwoWmqrea5Gk/CUNiq25qOsyeyUb0WxuN9teD0NVyZ1RQ1voOVA5ax2M
UGeP1fVE2VkJQDMs/cU7gTtN4O+OOGJ81TPxD9QtfIUXv/5Wt+PC/g1LnG2H03UB
euNOZsODT1dS7KEiQE2qZTCzRF2Jp8cySNCcvAspnepACviPhW8GjnJAWrMr1lKh
cUQff6z37tcUwYm+7GlmPnWEX4GYf1xdsjD9lebfy/gCwB3OwiB8U7kLOTzQc6Tz
/ma7+1c6ML9JwePoR5jTNRGzUGZtQG9keW7r0O2V7jeHF5X6NH3BDpDRCq/hvqeK
eIJxJ1/S16LN1+kKi9660x6OviLmZivfoTwClsEhIOaH+JYl6lo/7xhml7N96BOD
jX9LUu56ARWTV0qQDvtHA6a5wc0IsJganFOfm9YGvTzr6hpUA2RIRLNU01ezXpYg
AtgyoWkHtJIyNCObA/fXsGhYsom83I0zRjmm19f1eRZ31ViunjBjRwWT/jXVdRsU
dUDm0YHlqHwJGBaOrF9/IYbDYpAy5D4zROCD3TeoM+8zcUYf8OSaLQ73tocVJkGf
v0HURmpO70aiFwKr2yA7/UIZ2H4hJ/kefAiNoPkEAo36OFJ4CV5SBldxq2oo45Tr
HCVqoE+haA+xy7YyxG0YkF/siBVMJ2Jo1/0EG9SDjKMwI4rN8tJsLaLYUfudOs6S
aWredRfza6S7wwWqeNMLFOGfcbmNtasMKsjHdTd3Gm5+4V0DyKBqyOi2Ntl2l187
N505LKCE0jZG3HroM4/vm+ZiV7Vh5wxETGpgT1haUG0qfoLV2Un66UIAaQhojlrS
yZUl8x/SEyBcwHmYHgqPMR3OPdvVYGBaLSfZAebXQrSIZ22X1g7e/V/nReLt1G0b
I8zO7JsOrx6KxT0JmhBAXKq9HbpVnfMP/hhY/XuMDfgOou9jEU2aJCaZbth36HM0
daFz09Dh4ZAdSE7vH/edK+Wdv/5ZnabR7NeLZSsKfalo/L2l7hfmykAdxnez4+wy
//fdba0XH7KLoPP5frjFpBq3iML9iiUMSPxJCHG8pglSUif/wSZUHedgPF7JxY0o
UuVegf7NhEq27OdqhXe990ZMXAKSLri/0O71KGtldKQiBK2yCkGe3PXtTlA8TBhD
WUa3jsxzju4f46QF5mLa33Fh0lVx8EsVbGlxLxvjvyVJx1zrq1RnaG4DPyaxgg9P
mIH+UJ8GCGkd+JBju3xwyrPJ+petUombdge53/+NcwWeh7DtSQm8DOLuQZc0DuoA
IWXhw//pP0a+RxlaJUGXemmwiobJrXMRpzpnVFtq6iutEQONs/poRpe8EvXRmHqC
Ai/arCSxv8i2fYrcvWLIfHZabWIT4G1lsF1BdVNE8QM7JS0qIVZLErOFMVhkVhG0
I6enpMSKJCu4M9QtJpS9p2Y8FNxgrWjrH3rCw6bZJ/oStdePlFh1fctEMIxriHWM
dRQRyBofSgI3M1WG291HkEiv4E8Erg+PrlyMejSR9w43aOaJdVK9ZVB6RjtuThM+
2OlR7fw84V1AmXdPQr1YlH8kFmVqsmVjO+Kh7RA5+CuqBcSEM9MLv4xKVtlVV3Ec
/V0EUS+u7bZIeN2jewqIbZ6Text5ZqjiJ+yHBkAXDHr4GOsEH3dAcgExnUUlM/qM
J5xt6oZ5/+3+PnNUemd5A6Uab87dt3w9nOAoBI8JCbgV3SMHayotnKm5KMFw8iCz
j6GSm2YBWJriXcutTGcp5wTEguiNMZI08FnZk0r9eBqS24YigNwVed7emuvJc00a
4jcDa0J/TjA/DtkPYbQse+n2vBR4SVnYdxCLUbhNmpGFqn3wV9E8B/W1QwfUwHwy
FsY7NHh66JW3o7SUbgL0Aodgb7bPGseZXy2BdextllKasls6/TP6ouiVVKox8UYs
6RP0mrLhL5K0uPrpJzhY6psolzcB8JK8LxGmDRI9QnOYUdClDSkJrwb1pFa4YVr7
P9JyEUzBiZISBdbzJfNxtK4mpXSo6cp3OTP66DSC3i7QV7A7uW3kGrWDXCIUSbqs
3U+s+M4XmSG4HgIk9whWYkiDrrJ4QZXzfV9vB6U20llVyobwJtJCiygEIu0OX82x
wNrDsfeQf/YwnqumjsWPt4M9EApPkmjgO8ww8vcACvxIJt20rvu4bdxHOWUbKreT
WTv4+xRJSYUI8zOB9xxhbXKNMRtc60u+/AZVriiBjTy2G2h+cduDBVxlY1rCa0kc
Ygcuyyzz83nKYYOsHWSwD3l4NCgsUl3vo16JCapBuqMws9aeTt1UYQNHDuXeCPar
a9FRt73O0YWpay9DFztfYokVqTFvC/M/DlTonQ4fLBf4DRNq7RT/19+uv112B8qU
Uq/LBIeK96TRpHDLd2P/mSFDHPTmvYPwAjZpSkpZ9Zc8KefYUl6Xx31H2dYFxacY
WI2A3isND8c/fabtiq6ygvAw867xgUMSaH+WJZIClf7FL71wPQE5DeAk+G79O85j
KVT+qT3Pia0xkmsRuED1hk8GCKe9jWABwB+u2xQZUFgduARys+UEOQ1dFC4gKW0Q
b005iAvFLEMA7keCqbxQ6+WZTSqo4c1bOD5+g4Y+teW37C2LsJd9cjaRxQBYgu2I
dw9M8T9bC6nlPdfNHBk+DBClkSwAQQIqHS7/oKjRr+ymx4ds9mBpxYx5RlswKC/+
8iOyzv/4EAgd2TAPowrWfk/DHsaaJH2AQLHMXNQUSxdUwkMsosAPCwbwJRJfi2Va
huXOfAeecKiN25itW49Cx4VXE3JxT9lzqud9Y2vo3YxhEdHcUDCUUh8FIavwGBt4
uHitkBTk/IgVW/wQnT0nBCrbO7Yj1t/yRLlCwXKndYSdV8ju5HJf/7l+WiHFM94R
oOQfWtfFeQDxCqf29Qeut6EiHJpcppMzCVM/GYXok+kOu0OIVlfzyl2MehyIovQ/
79vpDxYxwJ3sQ4s1yZt0Lbcyq4vowYcNrRyEgNgrIQ2ufMLcxG1NArZZip5fb4zl
iJfqRASF1Vkw/JqPcD0Y5h0f56FFLAhSBUaBqzhiZ865/54kYji+sURwfW8WL21G
IvWI6ptOHfALoQQHhnsQEAIKxl+HWQA4JSBviyDcYJ3eDslco5q5HtBWaGsRzLCx
Ee8p+aMLA4fkMTUGFUEVkfRMhbKi/o8wne1+Wmu44WuWy63lHly5/4Zf1rH+S8Yv
wtvWVo+NIXxoSldb/HhAVs1I86XwfMstu/zf5wV2DBehHTm6FgGEiYBicH/yfzqN
FnHzITwc05Ikilnc77R56+zhhpD10rZOY3LfipJWsFrEHhlnMrpmAQ0tf2Yn5Y+Q
EPECbw1HQ5Y0J5SRLBuMDgSd/E+S2auhbdY4XLdGEFVpICilToYdIWziMlOxThyt
hJnzbGJX0GTrCc8s3IFYP9PDNY7tCsdh31Meyq6+TAtyfivqU6kxqpm16F1vLDzm
jwwoU4DQ2ioJQ3fOZR0PTRFAzRn41+WaWivEr/Zvf90qyEHTO2MfJ26IT62ybqTc
yvGGf/WzDvPo7mOVuoXpCzTykuXa61nePKiTFx2u2A/iHPhaiiJNAxzLil6sbjnj
R/6G4oC4+WrULisV49UGh2LuaRgk/NUA2+4L6zn2+QGkBTl5MnOazl4RkbdQajTU
9ZVOBmHbEji5HnMwnbKSZQ6wlnwypiUmZqUIQckonLj8y0CsAm/ey7rPtvO1dq+u
TdEfwiqg2+ydyLvT1Zj1TBKW3i6ga5TTlpyACwcshfpmVC/mGQDIDV9X3sRvKtEN
sAWzd+RdEc3wJhzA5rgqIEFOQddKdPh5F1h/1jLzHRY9iL00Xa4wWpdKPLU9sNju
mwGHnOC6Z56cWQ9ePgjiPunJXSfVsu6fViuVuGp4PCYwDgxrvVX2zKfng2ua81zr
dFm/2h80GNRCMu+3DupA3NP2D/4Nvk63RhwCvBWedtQvHf6OuL4gmQQ8fpTtuA7C
P3h3Jtr2u4/ZVpxrZL9JukcAUYz8Y6rlDyUkh+0UVlsMGy7z4tV+NTrx6MEYVdR+
q5NkSK1pYedlvbYtniC/8NjLOJ4W7hZclkH0Qxdbba253KLu2O4HikX58+arTQSf
VFdX4O8vkHnUNZI72YRWm9L3ts1x1BzCIygeOuLyBAfm7EdddWRpJ8nTceRklAUA
TZDLCFqpCB58kgfD6ZKfi5Z7IOG8q0IZdprn/1uSRl+WKzJbVb0AMawpTR96W+GL
h5q3oVI8OoadERyj9gj3K3DvZYHJshCKEhevNCyjHYaLJQKx1S/x/wOOu6aMyiqB
pRVSHU1GsBTz2W6yjZ3aLVVk1AipXS5kQViHv/ZI9qedwzqQas5hl13RjfQomSlA
EX6NeREzXA4KlC1mSWZqbU9S3viT677imsoy5UGVlZbiKHRpddZqFGdAzZ7wLKM/
At4IbYcBTUrAJiIgaXcXZx2vIPaLLXeUl6Kx4c2fzYgpX/kV+YdhB0IcUcIVzNok
NUePgpN9rm68T181SY/00FyOCDGsqoXpkmCA21WRHqG8acrnQqvwL12AplbLDHZU
1z7Z66CVHLmjSZ10lM0oWmwnGvu+NTrhH/xffp4HWVJp5R/QHQcVWq/xXOL3VqcZ
1Hjhan4Eogo4sKaJstOJg24J68NqTuiwVq/WffJz5dzl2YEJX8CTgn2kCGPJW/wT
sStkR5ToSnhgTVQQI3ro1ja2SiOXiBvhBlt5ZeIFLOtNrSBA6MXysHML6faT7dzn
a2UqzKVNlksmejweh8VG/b3rvQImRlT3t0KTa96henJfXNJzhM7s8QqPH+6bf6JQ
KatkewM/kUuKmUJzsWViEcmXoZl5t3t7+AFQaZCY2+XsVbGm9J9YCrWAuEwKeZrK
gy1+ZKaPxRObaBM88/agxXv46CGBFwLiPZPiE8CvfN5uJQaWo+FGXkiykUcENLIV
exEoggFvion2VRW5IGAkcSQmOnSYLLs/CUpaF1YVZaREyGv/5oLbbO+AKoKZt6ms
ZbSDtcMavkwczVxziJ59xIDy/rS0bOpAiGIWurXnblwCwHUg7kkpmS5Ql9/FV9GB
xJQqjfVbwhfevWLKqIJaoHRVGG1qAUEJsRzv5qIxVShCRq3HZe87wfpA2wI5O70R
1GKZwN5MKaeI4gGhTlYej8ZngoQosoWsV+06Jp5ROtL10KoPHsJmkU94HuPnWFWO
+zcCayB+oR6hS7uQp7fUREEZmW1v813S3rMF7QOUPmlam0IKXPHoIhbFTFRo3iIL
cTsfIkRwp9LtaABWsKriKwgV54WH6C/K7Z4a6vGOPPE3xr1BL5LDguejiQhMC3Bs
Wd5CSGveMJPfMlzSNQyWw/bkMYJp4YCJIreje3I1euUyiMXKQDuSIPJnYckZrNo0
R7QiDzDXE1l+2n8+Oz08x1wzoLvL4BALRWHPcvDFkYt0FT76lGjbO0lFn1+8TfP3
Uk0PRG8Fk8XvSSjvt2FVqLiAuQVoBWgrw/oqVMT3JFaYRy1I/gInKh5Y2oyKTaGn
V3pfUWwzii3Xug2Bi0i6pZTo3YhTGG4BaYtyNq2CV5q8nkDFTXNV8a3X2YTbZXvg
1s6zb/sVw+ukASZ09PwGihVolqRXltw0Yi3jWnZIhXK3vq2959Yg3y3103JVOhrR
L1awk0Q6oANPfsUylGxem+06HCwNLIjRNocJT5DAB06SgOo1gjXF1cwhRyBEVNmT
WRoeTV8xqcscPEEWYUcgS0qM2BW6I+3bKt0lD6F6mrR3fZEo4qPAGYcS5bqyan8j
BC73O7zVVnErqP0rT9H3XPShk64lnoW5bwKNt/itiMuMXzicgRhYGSoZxnUHkABk
d7hrKlFIDq2B/Taq+sOff5ROuKZ1jzk4ihInhBIQ/6ZUw0Pa10uwpn8aT162pCIU
ZjluGDPCrYwwT5ird1VLaMvQ5KiThs5/7NVFp+JXJL+UfxvLtIWxbEjb6zBQra8U
rA6nMEbjmzQpO67tUJ0ULe9y1yFpdRA9cQ6B+RIxS2HmCEoQJlvGGwZphadMBtRf
+uO424GVK+aerw3ttBCqzzeDX3CMnP/+GXvQyEmRPhgMz98mLz2DUPoLBEuDa6AG
swTAalhi4MTJkYlt7H+FrvJAPrdLKQhJu7aJVdwzyQQeQhRcrZZHVwdCNZWDIFzv
pnhJ6Y0v58OIVNuGRTWOgqOCU2Qa5fWH7lcT2nt/J++qR6gKw2Xgtbz1sCuyrxQB
v8fY7gBjXBwzMDcoK4HdoV5knwkQQ/EBxTXFlOM4zvxLADs9cFZiSEzoumXQ9Bg2
JpMJ1LbFcyW7NA9h5Tkz0r+Kqq4oXiusyT3nQfr+Gnss7M7WYlmPhPaMxev/7W6y
RkPCbWumCvcl7O+wJP0t4rsFScFH8kSpqR9s0Gi2SAdeseOXL5iNQs76QN7xy1PZ
IijdQDSWMr6jEYLGLqwDcAWZ9yWzn/M7KRLDDi2kAxm5DkmoiTLytk4dy4AtIWDo
VdZq9H3cF30xYL/xnIuH7cqPIopPDSRkS9rH6NvgQBwUsR1ciQiQVbSbHbUCYhol
EGuRx1G9CsJPHr5Ik3VXZc/jMFEEsTBIo34anTIS3Qfml42NOHgwnWVAQXm1YZNe
o8nbbZJCPIRcGoWx5gS6A0g6Ey8isKMpszzNS6FNGRYawtXh5Yy/J7P0mfGU34kS
A1dENu5nyCCkRalaBcCz46Ps5PX2Hc2YsBc9qSCNE8kBF9T/3wzJLRrzGdUld5sY
4Agw4SkP8/SQ4d+uskZ8FiA1KoNb7TKdvPWro+o64c3d03SwDhAo2aN4Lml3z/P9
wh5zp8YupvWpIerZpslebMBVUVwkyE+jPfb2rTZVg+W2GUkw8Ls2tW7e/bDk+rL3
Z3hg8zBZHRL54w6J5bVHTP7eJMf4h4sXk9B7bLPP7rW7kC+eiaG7/gl4mPoY9KGr
X5e6iiD0Nohg+1joHasI6/oreddBNVY6shFd4vzA9i7i8XiwQn6ySH9YdCQaFevs
MAhtfNfyoSZQDmy2uRSd3Nnm1OWU0g/p9F2ce96mr20kMcr3gX6IYwxxpNroDlvZ
lwPvQ5JQzIeRyVvMcS2wCicPGg3+vo2EfSoxCtQFswlUymiMbL6AEbhShfG67aEM
s1Edis8T5OxxolWmhWCKrJitrGQw3jl1fZFd54zilF+zQotS4q61QVSPx3Bc/lam
LxJFe0xCmN8R6w1D9St2qf8XYLsWWuYRiIW7hOMTP62f3tOJFy6D4upI4knTecW/
rAGsA6T5zVOek6r5FiIQ1IvRcK9q0e2FNj4SpoEtntdr/iPeM6OIgxcyaszQFM08
umWjyULjJNnMNaXMeQTg9YJS0NnSCGsqliZ9Ne2dtrIa/heTe/3TuptR5Ee84A3h
FQjHa1YYEcH/1EpOyvq5sKU0mceVAt14bkwquQYW/IsTADtT1XOZ2s9D5i5XwTSS
TdZq5+EcadKMx94cdp3zH2Oaw48HxBv8XfKgIitIWISevdMpmHSaAFOfd23w3eYM
BFWfq+HqxyxtzYW+2QX99Gu/vF+1Xe4A8rW4eYAMHp4E+6zOAuGhvHqB42d+6vY+
g6UsPLjM61YpqD/Zes49nukBSEmyrDWDdYAjqR7ZLFnVlrDK7kyPfb0MmSVP8YfB
KmJEqHrm2xS+ANmUWHJXzE9lT6ZYGvdsVQb1MZDqFKD2TmQx0LraiAMd7EbSb5Pl
gpJBh+kFbMHCytzlnlQbtAZRhcKz7H5QvIXu82cA2IooJ6a6i+HsMpvDCk+Q7d0s
mRif5ItqngEgofimvpg0hhupWQh3x6VX4et6hsZ0d8J4VBf9PifbbY+YtEHhduxR
c2ZXHR+0QAiFkBHsNJ6yEw4f7E0xCUzxG4fHUUtHnb71ROWMBN7oKOWrtV7UACNC
z2T9InhoJUF9YB8JB65E3Fx66ja1Ly+IpWzQTtzwRwpic1u3ERvqCxvGcr4FcmVY
+5zvvMDnalNAutg8W0qYjNve6I8cZS+NbYGqZgWj5Uuebp17MOYgLTb8Ih+3MQa/
2iRkHQF5lMeXDpJv7XZh6kAHQM17WfxtBdxJRgP4haN+XlovL6LwwwNW0IalL5aQ
isrB7TbUFcTspLIE2amMFOvCxfOO7ZiK8RAjA7RtKZRjGRz9evcyfMLQWxaFYEWH
8VBiSd05lQPFQ+zoCkV029PvF0GaqrqYOpal1cPLQ81eAKQTe0npBj41lWNaSLiF
kcYZe9txnfx23VNTE33rJVgQVc3/S3FH5TP+vfjbllwXVHjoVIg0g6wnkFdvK2Td
Z6vfxjUiuMzuWcbhqB0V+tRdwxQESj3MjCZR6TizrIv+OkBlj+ahnc8TXWeKam5M
sHJvSce9sT9qLtbC9ijkziyY2M7aZYmKLOKLVlBI48zdo5Ja0+xR82NAwRkaWhoe
fgTpqFCDBI/h4MARp2b1rZGhiJtgFPbkMja7whWz/myHN+PQoQwaAwWjtWb7Vu5I
OSOa4RvRqC98V82wmCY4lUh2TkZrPcUeqaX5hMELL+KpdVxBtqiM8wutVjRFjW7+
wEkPHtKka1XZ8Zy/SH3+JO8jO/S90q4O4PIBS46m89b2BgkQc0bRJ3psY2dOCkOe
nFIqwqzRhVDvTOuNUsPaRVd4Mdt1yao4MPPq1+MZ717X4ut0B/Yt4ZhA8uAah2HW
6BU9jvwNbmZA7qLluuW1sQ63My0Y6yUwZqoMj9vCa+ASVDwK3cn8JhyGvPi7RFy7
4G8wQVnfY77vlUP+0JHARw1sDYKxp6Zogr8LVF0ulcvOf8HwE3fduM3atU73pCcK
ZRIIcjuAkOBwwtcDXlPRWuqhdZLkwy+Ihk7/2y6vabc+fYjch/B/kb0ymgiq92p1
XP1+FpweCXSM6tZdI6aLeYsLzHTrAzfN83mDwqH4KQQ9mKMT7/vX51A5QvtWxqOR
lSv5+8ekzpv2ZAuU2JsD/cOdQQOKhMxPwWzKqfdEy1APq9dg+U9B1ehG+vsiMBvl
RNW/oLUkRHkSVcPRnjOHoQe40XLy89t9vdXAOzR33iuhr1mbFUkMcdXP7LdnciGO
ck6NU1jwjivBhVBKF50u7NDi/p2+zy/tWcL/Drnce37HdZomgKb5PCipUii/QY4i
qTQSYTcnqXydPN4fbaxIYIk0w27u7Oq+clDN0367Cirr7EEaBI4BNAs1yefopr8Z
SwJnFZtGaweI4B6pC1Ftndq+xm13v3XhYohOoEhMs984pivX9UvcpLffYIWqpRW0
AQSEDBU923kzEpwA4wUkkfzygiF5VgvgWJVlRvDmXs2KmqvS/WvEK4lyNRgX1Ewb
1x3HWI9zpLNhg10RG6wZ79C6DncN201DeI+x+Kd2R/Znke8yQSMJ5DredtS77CXq
Jq3wCEZIKBR3ZFD2xS+QKilY9pnIxEojlmE58JnH68bHq7vEt3zwslGvQ9l6uT6l
n89hNB8FYe7elehuQcfAIExR377OphK0XI4adiPC5hhrYAgxPZ5qZ9wZUhEFJ81K
Wo8OfXRIrRn7AOsCU42pl/gBkCZQ/WGtJXdRlL+Q+j+ZVDYAYELBY2TEaIOP/eKR
wn84aEEPSfQYSWsx7Yt0IE7aZ8txWO9FeI1DXBofEWxGsTc5G68t9mEcytyDEiB0
jnTdkFVyhtIAvVfoyoNuqS6h0D+ipRievSgpB71xyaSMoJiyc68KHFpzNQHqAH+Y
k2sEv+4fqyR0f15yg+1skGIK4CGbV+hnro9r0/O9OlJwJfWctP7VKOBzXUdVOKAD
rV0FejW7SG9b1KmNjzbIbifbtfO9MJCp1J6mnfe5x1a54VqYcO/bh/ASGYCWw6Yy
VF9+zm9rbmK7zwR/pYXzHdtz6I9dB8pPLlaAT0yrd7h2R8DNnLSM84B3HiCDWsv4
MJDFXu4+eXvfjNEjOiyEuQo85p+5flJOBag7FEGHwZSe/opdKyL7O7YlNBihtXcU
aCBtMr6x4bvM21Npt5QwgRq9Ut1EI0ChC1nh208PMsQNUnEFAxehuqudGQyTpZ0A
ClAQnKmLIkHlc51lyxB7vNlwug+qWyGxWyDCVP3Xea3BICIB9fniFKEE/EX+J83G
/fBy48zTamblMDHr0ojWExMWroxJUJxn57pyHpGTcd/IZS6J+TIM5OiYli1SgdCU
oWUHTeP/pKeAQYT7AZztFzhrzlVmalCi+/DsLqCBjRJHxjppVUcIDLdMk0JT4d4l
zmD6ipd3YmJx4XK193u/WkLNDMrfkLc3t/y4ZzRKGiH4C8UF/c9YBFx+AfIU4rs9
uslih4rRe/5JQkqqIq7MexscNNVYOBv/4KmHeG8+qeLv4jdd4f+hjNG9bNzRrY7c
VtxuZJy0vvdkji5kq2+uEBAcNQ5fDlasZ45aLyhw0QiRI4Zjz3SWszVVqnME0E6C
rwqo0kQh5a1JLOoK8Ls5eOg3hwFtvTyY6RIhD+j0vugNLqwZbaEt3qPq8xvqYipg
8hMy5k48NmeqfffLc+khISY9tdAhIh24NZsQfK+UZwaDrO2r/5KJzOBj3phJpIbU
b10JsF8WVyMj6mXWs1EC1nI1qiDZ9JXRCRUTFrXb0WmCbrunePAYTr7yprqsgad2
ztLF6DOeMoZ2QY09Ouien9jJRJcgvyfzraLOenGDUivt2itxOShZB4kqcfCflR2N
9xEvPR2ByK+V9yJe6EeW5Baq0Wm4MDSe2Dhz5MbygIaswMsF1v4tpBmBqBpNNzq2
nMq5AZKga9ArYXrBn0+89qInrv/uhTEKRqXU9RHkVAo2Gko652BuKsPhAQ107I1q
iOn/TzoyaPCiDFPjC4TnPguTqLz3+jefhbkXVnJGamiKEaJBTxDxL3djwUg5VUEI
ps5mQX1+guUnpDL9Mz3jE69TQ/exmmOTBM6JXtgjICvl8pWasZip2nKX3HomV6Uo
jDrUP5k2HYscsMLTVNZ2MTqpllC0EPFynt+/RstlsDPNHLEebVkr157S4GzActYj
Verw7E54hsKQl5GRKEqigAxOgG6EqEMgM82hCru4+OEICq8NZ0HVv3oqAi/yPlC+
i0MgEQy8c2B0eM2GrreeqcmY/RYWH87ygNEDxNSbiCYrrXljlkkVvITdCWYfh9wc
abxByv2CEf8nSaODYYG1AR0xExGXtZgmMvENWshJaLjIc5EfVJ6EiYLI646i1wJ5
Ebt3j0O5RBvr9LpOqpbE0jHFGdbTFlVwW0Y8/JaNDECiF3ulujWd1QAUQpcdQkRF
GhVi3lDBZOZb9z8+L+iTYOVRwWV1EDeUcFBKj5ZMKBZmtVI0B3a74VkDdMPkusg2
WXodagp+PaMYZY9JAgCLRQp2NZ+cdFjUc3E+wEESYkVBX5WNQ8tt/pr1j7SUYw2D
vZfQ784PFNhCOlTGIlDRQHdR+TAz3TCiLhtTBXCm1JgFbDW5PTjCT4YZ+CBn7V61
klS3u5zuGKINmTufiorNcPSc0fWDijg6DGgx+gW2hptf3RKkV4HyLByc7BKpCG84
x51/p1I8BbOxqhX1A83KgHbD64Qz7gpdYQZEIA1ZZMZ/Lg4MqKi7tlfwuHA4DLct
fmmb0WwhmOqwvHKaxnla9JcX/FNC117gkCINTnrJm71HeLHRv/jvmmMVYWe1yz00
yBNOQha/HNJioIJqif1zUwJVi7HdU5wppCWMxenI2eFviVTd6vYNcjoOrVxFKJ0u
IwWoUbUaZUin+28sXeBNCAWp1QmlNqhKGGsEXeO8dg7Y9SPezLYe3aHujsaEjgca
fn7f1kbsFdtuk0SaaYjxskvscXV4/dNYWuwQt4rR7rNKInoVvA/sUMvOCtlQwRub
VjRlZqgDWgxE/h/61Qv7CEasPvzKtW6qh+j+EeBRIcEfgPsvh7B0NDKZw7+yDYRd
hZUsHwQoysYoALl6gV28mt4YzGJiT2QPWMLcnWyNuVZYVC5/s90NBV4ScmfDAHTG
m6PwVGBbfJIvAs7i9HbrFEwlRn/XiWkSx40xzLEP+3Qq32oII6bXZ4TcXqnGXGht
3TPJm3sXFlzDiyZ+mF3Th0/pi9WYzXipIVmAaIZ+K7zbZtes8rCuV3I61uZlbRBC
03xemla0dFAHWrlPhQ9uEVV1/OqhyTvm8JbBDwH+p6Y0IGn3j3JHKn2S1eG9FSO6
LAoOyIv9poq0WLFE7Z8LN/Rik1rtn2rSjzyyd20UXWrjeTFDeq4SqPaYf8vL54dg
jxCpqNj8NDu/8IFuI16AjYV4ow1lWiSRniwqCMCVbyvRTwnaad+qkpX2knmX50Oa
l8XjfypoVaElUFwJBZka6fUsC45TjwvA2UsvL3NWryUIUmSslDSr20TMVGbazScl
04JRo2L5crQQfeYsSOStHx2Tkz90HsZ/OPRbklbMyANzBNSHlYZngCpJgoa4I74A
JF4dX+IG/N9+lrpVa50Z4p3FvYM/7QEsolPX+1LWvUqo9/UFgWAjTmE8kZ97SyUY
GI5DitM8wTubj1sgUFIidpdu0qf7znuQNLx/bE3G2OnpqS8xuEkYDo2eYD8Fr1kT
zDYgkjo/DtrIxE/NSqSACLhTf8EQWxeNhrbT/kB/d10P1xcN/Wf/7Zh8kO4ybSu+
bwNLml80Tc1hi4v/OQoTRIssGf6aHbCervSZuydOWDbwNqvgZhXiaeDA3vh7ddel
oJLrTXTVz9sFjik7LW7P2YQlJcoQglTvCU1OokhNYcpRsxQ+PBihUeYiFS/U37ca
qHv3Auvw4viiDVHZPEarJprXeyIOS4GwOOuS1xRL6kLG9yS1uL3tnC0tDmPTcTCV
nb6p0LQmdgh2u+eeltvi41uhG3iFVatOjJ8D9cGyqPHWVErQN4Gz1VHQjrd2pXCP
D3zyG3GN9rUnpYF9c15FpC5UYSjH8R8tJNo8fy/z/06Hzl59gFStdvRD6CBjDm/C
fFY6uzo9t4PryTpivvFuY6yAzeqah4rQSsOedek6gFMIatpiKpEfoE/jO3xgdnBt
np8akiBHx23qV1/bwYP8sVX55RTAI4YySnwuyatmTMVAHZi1lK0xDIr++WJsFZte
HsV3ahcw1DF/dq3Ds4nf1sDedZ+Hi4LHeC3ULhi4Y+dT2QYwD2UGi/77Tyegjax5
HltpE4vpJyjKlVoWU503ZeZh5z98UgntQmWPqvU8RX1NhDeqS821I+8CDghFlDWU
py2FYg2COFZB+R3nR+G3Ze3HMOxht2f7RfzdeyDlnrEZ3V5uixAyIRTHquMC7Skj
zrLy/W1zBwS06waOhRErhM5DGjDnDgSTJocxN2IjBgV4fg1uT/Sl7BiJIKBVgwdE
78qG++c/+wlnYZfqSRjJPohF2m1EI0iff4J0jxTuZdNivL8AynxBH0kZ3yjRPxEP
b6GJRuYplbZYbIuDXVOL2HvV2zP0fLHAlwmlOe4RJwfVXhr2SK+eOYFi2Bfyjeob
txqQ5odIcpMYXH0ODZJvUdkxE2r0lq81ZAvLoDeUz9rk77qBSTts9QSnumTt5QHm
E+49llfihOBrJCoSTk/K/mNvyet6KFj9/Qh2T0fExo0M9+jkKQTJJ9j23jcQpNCK
C/9FouYnQaiuuUCC07jLqsS3QD3l17fmg8G2Kfwro5p7Zqmg5kcYIbpHXQ0HwEfd
kubGohSq6uRIcBpteAwVkfJvlvdFL4dnFJFZhBEpNUJfPibyXK07i7gbYsCLcQag
LprKhTdacjswo5a6bYDQWSo/r1ueGzXFVt97fEgBWhjqw0uLKR50FQwX3WWFre4x
Detf2Sg1FzCgwPqoYLuIHEdMsIe86M0yHuBDddK/Ot4Pr9J+EkdDsi683ht6l9cm
oFrw0j4UGrOATroz1UPQPyLRdpCVdAZ6wsbTHDhSbLPGNiE0N/OAgTPosJZo9qff
yyRHaXfG1J1jJ32dJ5qAOmUvyD7Q4udT3/p3kD/u6d1w8XX3a76XrQ7p3SKA4C55
NowPdXZrPg2q3wy/qqcEUpoGfw8GiOr/EFh24tbSlDUEZlneSId7l9WlGbrfCz1N
OQA3jSQKkLuIhTD3z1mbx1uPx68Sny714APwJqHkOR6MHd67dyuKJjWGAYAkVc+4
7XKJhxQTGY3YokWz5ha8ScHuwEXP6wPgU65VJv7VU8qfb8pvxwhlWnva1ikRbBSW
XspbLfMEjiPicfSpIh4EaaRsyRD7b9SLGiO6WGQohY+PwWFRjnbZKAMaBzoIhKvh
RYz77KcylKax3bSMwcBR39iFEojB6LEsqoE0lN84af/eLtr2BQYbZ+gwvp8yRqvk
CWa2pmxzbNWViuYXZfKlKE6ZdIYew+znauEQgdbbMI5gkYRvJZM4p72NFT1E9t4i
hNxIvQQIBrb9pG88Bmu6wlvOpa9/WgSZJwwq3vX6iEff3kcbCF1V2vSCa/icveYq
kD89MQODtxGhQEyhtL7r3+14FgTE/Y0L/1BfDXeQMmYWWeo1OEd2EJyLdw3g4XUW
GxaDM0e7lUct6zYLFZw0kFxTcUCok+l7BnL1SLOVFlxfcbdVyDI/wcP50LJ/lKAl
Gmeo7ahZYAmzrRnTXDhlIDlBElTfGgldE3L7zep/Tq3paVJ0C5ZHiyJcljShHf5h
pg8ZaxAzFHE28sDhEVfiI/oxSe0uRJvsS/aIdTol83cIWGjH+C2KQsEBKHpInAMk
pmkArZxWSp5bTfeVFFB5qfYhXr570QcZvKjPGuGLouJY9Sf8nEjPLb0BuAFfQVnE
RxRNlJ0IdmWKmf/9RqnIcvFwflABXvhmVEozOXpNOJnY8vlLjn1uTscE6DAkALG9
JdVdgaopCg2eR6B2RxlVb/3ms85cPA9/tqSOzwBQxSFb+Ot55iQ1g4wNAbAFxp0K
x6CLJYO6FE5T3ZWN6zQ7SdaA3G8BSeqtinN4wf6vuDPgHxD1MQtTnE9GJNdI+Rj+
9HuggugjVHFqPV+LW34obcIMUa8sf0fHnL2iqq717brGZFXtA9/Q9ROSXKZseIIc
YK6vOg439P59Am5TNO0YcSkMZw7mqkkb9B+1mpUu/AJS3yHQmKeuFfuCgh2fuVd4
FXVXvTsW9o5OOCA725BoOWot2NgQUf4ZbzqyfAVJH6lf2q4tygi1wknS8iaqzLL7
hxXEsTk+X5QaCEGhHNfxvt47EvPhqIetV7PJBM6NO43RhhJkONOOvaX3SBd/Kuud
ejf+hnAnkYTnYn2vtkwJWi7dLo8Yj/W1A7xCKl6OYYraOKMAwwY3XTY9n1Tg40Ns
LofsC6OvagkQ4ZaFkq45CU9R50l+r1Uf3Dqf3upy0W8DvBGAojtHTfTW+ZcTz/E0
j36+jZE2uAJHLrXTm23lJwdcKkHThX6G339PajqfmLAeileZldbQArieA0RRtiDC
rYJoEZNw1OMJqFsu3NN0t85KMLXju/4vBk/meKiB6NqRFRV+zvK5GoZzFHM1l7my
g6NGmmgfoLdhFJY6p9skIqCgNqCvnbzWoBpL1w0O1yyvvyO7HWNa88s7JUEZclWT
0i6vFtfTbtk3wPAgrl1ng4DoTL9sJWGMxO9UYU5iMs4EzxODMr8e7+umJNr2RWp7
HkLgiBS+YcOyxF4SkKrlgvt962v88gMXE3pei+tTtaNjkJxj/wohnugBbtvmH6AH
d5iNPOBI8zxjPVqCJW7qEY4LdAltraZqr3aNOAhlCMEb1HsF50VBQzWcerD3jdQE
gUC5toRBA5XAcsawIpaxs+tHL7EDorkHi8pH2tGOAB69wxiXrQnkhVYKHHcMclcN
h+90wzKEEZk+IOLDkz9jocVN1exZyUHoQe6e4PK1W1pYJRf3oxuNuZrP+zPbdZJe
O+1Y6T5M8YG8iMp0rdmtfG5KCI5LxI3ZRVhmsXAUILF1e1rN4S+W52soE5cc8ZJs
3V14m/zJmXov/ngWY+LXKMCuncCX6K7R6BaDZyYfvFOfQMIEVfeqwcuIRNmYG/FY
ixhel0XKMuaXvOmNcBCxDYUcJo6vM4OJJpbAQuA5f4vtRMwbfAeLCqa1P5eZvaub
2wV5yk/1o1t5YGy3BeTmhZGWmufTd8/IWKXVJjyUef1JJmih3YVwVIbi0yHN+/6j
zFpdSjcTFlxH2dkNA3VZ4XkmtbHNWHeOE5PQ7nvi9G62izGUerpPhvdtTJ8qcp6Q
oEQI60wRqDL7JZG2hhnNrFEPKpFah40D3Tbm7TenOn6wy/uBaLrjT6n6lkVergAP
Ld1gsVSeLQx4cOhyuj41cEwtL1jpGpsxzbfShRvkDbtWOtciSBQAC2vPAEXq6O4W
11/9tOo190OUzmnrjX5L+up55VwOogjFHM2NqgyCtmTdq8PVYk9lndr5FYrijHf8
hyqmam/vgJc6QbyZTseAPnHS2HLkdpgMVrOmWyUwhYLcti1FJOevO23HuA9EsQtx
rJAp513KewmnLU7es2MW+ZnIpEYoftyijc5orJ1WVQKsymdJUVZLO1aC+GddlPrD
31BjJ0gL68I6CexnyVdr1/DlTgNUOqkgjiO8NkAHVWJR7QCJhtlGAAi2QuZTDcdX
HmPz90gY5+3Ez7+2jMG7yeYuuimAW4UMFe1sc2gD9z4s1mbkweA1UiSvnjUME60R
nJi7IIpkOB0jh8LRZwGZAcd7pu+lCF4k9ox/eOdPd+AL9jJnNZDIDmqh/buJCUD4
yFM69LFgcod6P2MIQ9ZDqgYMrCqeemtT//WlMNF8M4XQ5/i48BMYKnGPxVldpVrV
gnH+3niqhoR8PKD+PkYEkW7YjT6zr7A6Lq9X9Vr0t42lA0kEMypEZLYTR9tfUcOg
m3O32y1P7KRjdYy8fPOuec9YtpOezLQNMw4k9ACLhKnNG+IrrMqwLNf3beOEaRrf
iHEbzsDWxhLk97w16VkqTL9CtXOaTdvaei9TMDh7yrR7yK4/VcKKmv1POiUK2/1o
EtARbNKvAiX3C2gdo6eaw3yHJgYSugHC7aWz/MKC/1zdtKTNcDufkNXNiDCXJxlm
V9S8i4pdxr9aY6yJ8hO8v/SRSvASWZR2fIWkf3DSIppDbfOf937A+J05TOa5zNMH
AnSGGzlIpApQeCc5OFyLM569VeXotkIPzLqppqOAf1GYtR6n+eTLv7mhXxwUuhgF
tqwj+0fcIRMx1j6v6VJangA9twDf70Tgq4OddFSLIDKdjLOwxYikjQilNXPo/Nc8
qXOJibdQ1MMRUem8VVIlQPniKXgU8dqf2lFsdxymhDvlsJx3xcUARGRvQGldLJZ6
eSDeBlHYOv5om595LQG6BxBiaQ34e8EvE5UnzpTUvATQesgkiA2T1SGYsI/2Lbb6
i4rl6xcsEAQfqIJhzl7aokRvhWzHizbvRF99aIAQKYhEi/E9SfG0UDN5hOxomMRi
HyZKe+MN67c+cEb+Q0UlhGVT70RsKZ1kyi3oR5ff+gMO4a8lePtH6lgT0zckzfca
b3p8i2KK5w+pRIN5CwQEgfJ9MW+Ti+2Vz6LFQW+M+B+GPzFvgYzBJY/DiO846GQ3
lJoZe0SMavgAp6PDN5Xt9HToAn1hFdbi7eFLB2XIOnl4S2rA48+uvubHXypE6QoO
PMSz5vjOxsaaxY4mBQDRHSNe5wrmOHEe98mOM0CSSM8VFsgHjvn132HTHSvyuPYb
D9os+CPKgEi0Xa4aP5BSez0t4ecga0ui8ysqNPh522dLUNOz5yGPbT0f9rPEb8ov
4q0DEile4VSXms2fosEfuIpNouvNSrmVIhvGHvLc0aIW/vZiQodNPZ7ouokqYxUj
IarKdCVKlcexaQtoWyqjn9Rr7ung6EosZ8k2MozBTs7U4332ANtT5X9wAaJkgDnl
wAR8pkfJuLffU+d7TLAgVCXQgN4Ey5By6NMPRDEjia2sLyQEoVblzy0Cec/AGX7Z
dsgTPmXHx/GZ8P3o7vRDDurSSFlKROFwTl0TyBuzjJ8Sp/RzIA26wudhQVCN54ag
o2d9AewsIrEuYo/VH4ug3EYzOTr9IZXJWGYCuaiZvn4XHoRCoGgidSs0whD31MOC
jAtNVM9ZOg7iXLjfeOYzNDy3R9Xy2e7I+ROrIkIT9cMAV4/9zH6ryiXJEFmpwYLk
I2ZDYxYgkjonD+lb+EU/ZL9bkG+IvFZAuDjeIfXF4zA94dp/In4QoCvGvvK1rynB
03nHuQOWmOm0pbNn+n7u8j3C1ewG1zMY/zAqusIJ1lGpYKTMERkSyCAaalqEOmZ7
4rajqP6Ks+v2Zisze0dWwONoQUbwq8Xx1LvdJgqMHVV+iWGyY0GMq60wEH/LY5Uz
ZlaXUPA7JC+T9aMw+VriKAPPwFB+dNoaGuqEeqyf5W1DKQEMxVyfb+wdQq2ze2vw
N1PHClJ9ABW0Nw92F2NtWfkqsZkXI5le0msf6rNCBMJiKfMfpb/wYRU0QsNi0bx+
dXwTvWcTn4+MIDUSf/3kk0MR/FcH3lD4fMofy66R++nlKI1GVZ7ju6tTIpiAufHq
CvDov9zs252WDOY9zs1yUvvrjcf7eqVudhfPVVAPmRLeNg9OODHR/NirYnMGe5d/
ow/NE724W4qiB2ncJ/DCnHhYHQzlRBBRk7JyM2yt574naJzwt9GfEfWqo5EZJegZ
nK6jUjE8XTq95XQCQrcWDHtGGlJj8vzVeMP0f22gFQIcHtK6gt9OjBSFoNrVvynI
xl2g3cxTl5IWf17+Kkh7YkEHHMo73MjkLasS+UqL8R4ycBCQ/AKmlofT9i7fDwEa
As9myCuqMJ2KTWbNqzSV3bVB9u6EIUJ2nA419jLxXhlStbxi+K251WWFhdRrVvvz
tpVPFioSvRK1o0q3bwzXcb0Ht/3lGTovM3LFYlA8bWM6qwYdgxdmFCKLqVKuL+rU
X9lvqJk6WN1+tRFszT8JcoGTS5QZEoWSrcx4iUFXMPwfueVfIFk4VQ6en0xBbJ4y
SVZIuEYY8r/yhJp4m1r6tvPpc5EwKFWAI/buJHj1vRkJ2dsamrh0ywI3PelnOQa3
UG5UW6RYk0Oi1Y/w/WG/Hht++fhXcUPLsoZXrJvlH0OV8Ex8COg16wZyZZCZCJ+k
xREtz6P/BRQZYIqyQu4247O2Uj7fIp7z1uFZtlsYVynpbK/LrWL0QBqpLO2ghRqb
M6Tup/XnUrU6RMOVNuaUsvDaaoCjauBVEHnUDHxFqbepSG0gzhpj32hf8yBc7cDN
dAwYrho30g9Aekfkz6MR28B+evvrgwpozYRiCYJo21eQ24ii3xEejpKY5DzVbs/W
izTKXEApPBwfhMXuUA7ZzR/KfcOW4D3bPRKNZoOFmAG+eWnI1eTx388TvZUDAIsh
wO6WHh7ORNCCfOhcWbbrEqUPmBG8tsPzgJp2TT99w/ARbrRsMZco5/royxCHH1Ra
IJVF9EkSpiR140TfAheeEUioNfsSzERugDGJvEn9TjU13WrC0jT5eO7fQMh4N17m
Gll9y3Gap11rjQuHIC0xDn13Z8+M4DRwvapYy02SmUqT4Z6YAVzYLuMZxnMOxUq6
d/2mto0gwdoewUaL6gL97DxYITL+tQWzCIQDvDKLH718KNwbqcUii4Ctivm5f+V2
Z6RZ7BizqEob75ZtR7lmdUe4WzKmAjttC+w7/foT9Q3n8LVrXWuk4xt2WvWVu21x
rtPilUCjeRjTefU3lQBncS/jo6ZeL7z0K063fcJtnQF9AvmUInHJpnqNAQSXR5sx
4O9AblwjUgKXe+qtpeqYrcWbMyGkLxIbPJpNfC0VGw/T1NZLsBydMHQ4cp3nWQhd
WTxhymRcHGUYq9vuSyxke6apkeSUoCfj4Rg0rjBIITwJ9kLSiFpmk1j/TBT9Q92I
MRVrGGFojDpxJl8faFkLbxEkLdqruXFDacibaoAYBZUAiaFEgYApnAwRugpZEhrm
iPpk8JRIfjtGNs1DapgQRghRrvLnLsfIsA5XyodtUDznTcSnjg9UHMwiz3ktnzEF
bPy2XP8qgG+KHfeIBmjU8X6a/anuq1knel7J+9+BHkE73GHnEvSai0ya3/QRbDoD
05aDoU5k8QH2aXyDW3SANJbHLn0JWfgtH1nS9dRybi7pWRLY7hfTughORqxoDEwg
rIPbT049X0oVCfvaODZBFHT40ko+HMaGCWIXTitqUStBKa6x8FwZGM1ZlzCub01E
7XANkMLCAjEG2nqlxKeDHJBRcVWkHjGlDH4D/rnbK7glGV20UZ8VZU+zNNnBTRtk
ApoGDqnXmwP74sqS5Al+9NOJruDPlw1E/m01Ky46fxdYWTH1wcps3/zbJ8nu4pIp
38l61s5C4PD5Zguy6GrBlkCLGWLAdPTBZYriaK3xyDVKwm+DQoeTLip/fa173txs
PVyivpQ5ZcFtEZt64H5xFj4LCK01wF9YJ7p4FtCTUv2dKac2BCelbGT2HlnZZkCc
9WNCC13Wu2jcU91wsi+7eSm0hQ+XFhxdTHed7O4PZTLlMlBE+EYT9wMA0rQBZ3h7
MN4766Pz7AH4kOCffqxn7TlFcXHyA/FUJSSENux394Sx6YG4cQ5du97P9lzjqaTS
Ho1756iIefXcdVbjcPik7sSkSFzcNo4bevpGQNM9Eu2h3k0d1HZ4FZlN0idDp63E
ua8E1b/EeTRc9piiDP4xv4JtSJEcTI72rkHJy1sDOX1ypdi+V/xC7ELybLRutXdt
92d/lNnKaa/7RvPRPUkoN9q+PVDeChS/2caHbxY1vDxdPBq/MBtckq/7qUxxdkyp
wEYlH+XPktPeH80DhvQdIndq8fo4bx+fNd9Cm3bnhuxrFDFMA+dF0h2OMjtBFjI0
Mlgu/vd6S366Oe8g0RAAB5/AQfthDWsHXMRkr9v6T1aUAKEHpidHfqV5JAUqUXym
bdFXAzpkLZn3KOgIFvZBdd/FBFSe9+/G7RsENT6UYj9EmkhIVCW17ASZ0cQZNmIl
xpB66aq1ETRiqncuHPa0CXig9m0galOSMVk0YyEwaeklkdmwR40ywkFmVRDw4EOS
AYtxN6ZHDrC2TfcGcql/9PNoTlBQYfe6n8BsPxfVwBMnNaVcT0vpJ8JZcgP9ylPF
eQ0W81EQynwAWslcA0BfKoi+Q+Ndif+3c8u9DBKg5CtqLOXNV6B71L3Ld7XFaDkk
T4+t7RkyaBZIDC4HJaxe6sC18Ldsiv2epb/StWIdDz14912R/K3jrsJ1qE4MFOfE
mVlaUIy7aEA87WEmgLjy+8lUJbOCqqgHu8gV87swSjnHRNaHyw+bxR5ZxF+oMFtc
X3whXFtXTBvyr81eNHi2tvVYZPzCqWLYMp0rVaoQXyPB7aowG1+QVTm/1xgo+NH8
EhZuxF6W4lpEKo1V8UysLp74oatoV46se/qWLqododMiOfxKxvgt12i6JorNN1YX
j7Z2dwCMW0Lk40i0Fh33CjvQj15AKR/UnpxJwvAtn65sWwzPM9hE0rV6RieA4eN+
VNXwrQR4qSQ+IcfD85H5Apw630Rr1RihhWfovY9hJG0fdpF+RnP9aMCNJr6rbYk5
dczqNgnod4fu654PfU6jGpMuB7mOtIL+8ZJEkwDdOnnpVywC46+JBTP0mmN9Wpi9
4hJx7dBcXPjaquglutil0RMxMstPIDcZfvj3cFw7iazu3R1MtOs3ONtXF+D0wrTs
820G2uhoUlRSOrd2QnMk6p6lFOs9QEKv7m5P6jLIuDP85meGOYjzeNXI7f/L/iCj
6GszwO5lhAQSPQ6xqMM3r2mkZQPqsJmHsjr/QlZG6uO4PvB6A3Oiu2DcfxvU652n
Vwm0Sc2uFR1J0mc23g2d9CRV3o57iINbHujt2cku+eqYg4Yl/+7uYhmG5NDfJx7/
NGIjkZTNz8Kp3URW4EdMKFN89tT+rjRrjlYvZ1VBtdHKxKdFslQJbJXSL/g6onij
yeiBIgp8Q92vhBfivI6eNxFVXVJoJ9hWFjnamNugjJjinYySnPiIbjY8jdvKQsWy
wpSaCe8hJXe9xps4Q0MXpDOjtWgNgDuEqt0seZMoPOiF8srMGc3d+rU7omk5091V
MSkunranrYUGskZVmBOAVLJ7CcEN1EYmcpaL4qn1gfJsvGhQGWTgx2l9JS8KKZWM
FV46DigCXF88yZ0WJiENjDL2wN8S8upqvwXH3En6/TM5uh0HH8aKGTBYlfcZ68Gq
lAbubkgrKMNnTJ72rTu92yyvQsDC3tvXho0ctel6NKLUNFxDt/L+RsWsWVULw2Q1
tFChf3+xH03yWPPkmUN9TqWtNH4sr5xHxkQU6A1ADF4SUFrOcgYcVpJ5p0Qm/wQG
P3XRNqWqD1N7edUqyRSAmdG3qNLyPS5Fj8HOe/yLg1s6NXoZchEN5sbWHTzpFzNh
psWA42ib0iR6AhAH8CtJJ6BLILbS6Cu5TtqTxCiEo+ZTEjtS2Ti3gsIvdRbu2nhb
n0w9W+e0Rv8uSVR1cC1y5C3X6EoSMArOQHw7WNB85CIBDVFecItH5kcr43NxBkIM
+6m/YNRiLFn4AI1JM9nY/YgbjbO5WF/VSoKxJCMJ5qQb5Lbq3O4wjlF47jFiv92D
tuJ8qybVnLHjYlNcY+LhZZvTjGDELJCwvpXjfppPpJXJCtwlXJk+d2TTGrMXAkK0
3GEdX/PzL9RfbfFdlkTEcUx6ZsZqqps5LrKgKWVG21xboD8FS7fXSOsrV6LP3shD
EBjzSJ3AdlPIoQI+kQvI8y7x3IEKlQp/7WqdbzXCn/TZWhzJ+8JAjsypqIgtbiZg
uERQ76EiYyYSsQR0BdkWLdZ/6tATQe9Hj6nswVuuHcdeBg14S/YcWeORhb/fT6Cy
qSLqs6WGJWHPTiRVUwtP2P56KZXKpoc9hGRDQIEJZmPyms2HGa5IiXSW5aBuGKBe
r+i8Guk6QtEH9FL/SMnG/KlghJ+WhZltHPh5zrA3F1dWpfAKBQpSavIRYXTF87hX
u7PGPdUyC2csH0dHzVByW7YgPJneFs6eQghR8bngoBecVippdK4hRp6UV7fpdIHN
O8vwzXHwMJTrnpWukItqe2Zc9/1deBVq5yd2uCmJ9gdQe7CZ+BGQv/uaGBXn/elT
o64Zq94ngBmNl1/xr7JQda7qXeBZm5s1TAigUIro/UTFKamhKQzGbp4nSOpYXXjr
eIGaThb7GcnQ8KQ9nf6QkCivjz4ot9/odbEw9GLKOxPmned9jtFUDlRcPU6gIx79
daxk6qCz/MWLpvNjX8NsAQJ6+Dpb/XBV/9FY0UGGP4vSzomrwpIedZOGRqoAhVvC
nW46Fo5Wq6nDGvLZ1+XiZHo02g3gDJTDLOyxgItmXkq9qZl0keR8Xt16wAbSF8IB
GAUZf6tkEvvMBwfibrrhNyzncIxIVDS7erZbMBVEt/MsjONX//3UW2irKD+Aiufn
mPZ+rhv3VOe6Tca3bFGR2kx7tIOQCl+KWHQiR496MHhF2rF+aUJwJPDz0ZAfMcGe
bWmW/uj8P6PkVcf9QxDzTqJ62qzVHuLKMKLgd493Tq1YWpdKdEMRo/2VrDz0m0un
+O5v179xuR8GBoo7XZznW7kcCYLuhV2pBI19swwJcASid5Ma3S2vVlydKfb8Zymu
CAghF9SeluQjc9fyCiza6iPoTyDHabiGKRs+R9x2DKB1UQeNq/XkmdivSbD1eo3Q
s1n5Nfi9kZq8Gq+UcrbeReae7AzfQUQwEps1qBSXoNPW4dQPDHtthyg4R27LF8Eu
PH6teuRPn6u1JUl0evkdDXb4psU+NwCQj8M/xL0Rkr9VJZFbSJawcBrcrQpr8W25
zv0u+xszueFl2d9ulmLFmgWyWlY8V5pgis5r2CUFXNhx5Ornxsi2RlbShFTI1AoM
1EK/9i9W8zA3uNSFPZ8CnwdV8yscJI3HWCmELp08pD4Wu1C6WptGB8ESjLaOgsJ4
QSpFxtDPru+iHdR2bHCdQ8lmwCgm6aFZVtUWlhE5gq8Qi45nBsEdw9hidpZx0rNb
6Dkcm4p+cZAoEhXLVOkwd9xRDtXTTLK9TatlYHUSkbRnJmM6rB7vE35WSm69FXhz
gqzcV07x3W0dWTfXGl6+wDqf5Ns6VHV4MPeQZhoNDTMvky2TU/Un1JoMzH2M/NJZ
WVLGRDVng592IDlDHCAfD4tJDr3YHMuHDIze/IbhxtTL21+MSsHasiXp1NbmYKeE
iJEdERqFBuP3VJjwxl120drbnwxkRcil3lzKAJkr7zOpF7SPHZJhh+TJuCpeCFRN
GG7C/O508MC0LtA/M1oOl+L3vMqRYQGUrM6tOzfZdfsevfBrazhCjEWMUuUsbrqr
P1vOLlCvWRD9tOBBkIHoFy2gCvRsix1DMeAO8nl7/Y+3AZAffiRw91Oo3+4GfTYa
pqen2KMgIXT4Mv6vVpbtlc9Uh2iYFS/AXS+mAJB5E9wNgBjhOvOym8Oc3tTgNzj4
4wYBbTUm9tRQ9YvPTdj3CoBBxI1+CcG5iy2ZkDtkrEihgBvfty3+/jCxfBoYY0Sd
nRqRLZhnyjTANgpPReGAu9VjjR+7BZA3vX6mhilXdcA1rUZSDMPk9wNFf4Wgghnc
j66JdQKE2uY7iSlXvaL6Gsa2IlIoiUGfOdRWR9L1IIXdG5P5LAYlxfDQbuAl4qbR
Er0EtPfsZDef3fdYoSUG+tf9otLxge+YnmlhOOAImCDUpBInATDHalxjyrNoc/FI
DCMpRagX4n4l2IAAksMn/o7K+9673qbZAmlqeED9GuMOuGkpC1nomGTL9e2yshT8
B9LkjYB8pXamxtCWwS5xPEJrcw/T6y95XaNqlpIYGvu4uIftf/C52ndD6UM9/Yg+
ZhYEWJWeSUeZujC5SUZjw2GvYkGECGblNOF6drqkA/QKPXuyu2ldKz2n7PvKtjDd
fzxIYjbeN+/gQFa1WtS9a8Za7SFpRzwbyG1e6vM+XK1IX2bPeEdeJhO6X1TZ8l8A
fhulLsgJHqWJ4Gxj08fCsDd2Y/i5rojPlilSlYlIqtllX+C9QhJxbPuDr6tceIuK
hyVlOD5n53U0ODkiiy4xZ/XINipwCgO4KDlwBsT6D16Z0EhPOLczdwqoWN5TLZdc
a2raLafkO17lNRBMyVC9RINPzDZOU6S0Mt0RRKDPRSfxmXjHq+lHXO7GMz3CIUXJ
MHsOEl9S/+ViPobxmJRRzBo3QcaXYP9LkVTwdSUbmCdbQmBMVKSPgs2ed3SZ/nKY
YbHBtUU76iT4ehln/jxNTZMZQ7yzuaajmkPVBobkqolQrgvxgEyCT97iOSpy5NPS
HoAiSWob+4mkVtQ6u22+ISLAj+FwfdxaZKuApBTElaw75l9p9rXwT2Mr4excNKzV
KrVjHZ/jJ1uPIondf+5Y43KpRHTyGZutmDup0CbsR5JKmrqVaa/Qbf31cO0tu8Ov
vH4NXapGfaLM1p7ljVLs+bEvg1EWkPi0+HsetmTulNFUzMAzbVK5cBhh8oyodlhr
srKclA0X7XaI2EB4m0qtqu6pNxaJNBuFFf7keykCXNxJS6WNMC2kzxTKpldNvMbj
dkHaVdgMBDew+BtQzmP8asrnh8wV1etIN6ARGZvQJE+jntXANdKloV51M/CYOjAW
e0BwlUD9EV2kVp/CANkokIHLK/Goc0H8tJsU/dX/eURAiZvR7VMAGwo116f72aN5
uvsXZtJfkNpK10557gjn4O5iDbsgtnRvvq6ZwWSeTVseMf/b7VUHChExLwKFuCJ7
VsmNvgiG04vTIAgr7xLNRFJvksRh29RHk4DrbJWtdH08f5FZJDH9q4q8gPeL+aS7
DEWDmWGsuVGTsviRYW3HUgPICTtsjA9eFNYFZxeMSkAw9FbGmDmt9EQCA7z0osyt
edFaJ/ZIAaByCtiBmwUX5nEC0Yhkjf1N1zVh8P5BQdxp+5GvaP+RpQ7bCpb+XExj
BPISDMuMvx3oqNM7xUO3U1yKMmd4jrXmsfVeHpyhQ8cN18/aaHl+spMwOVB8G7Ju
cC9CcH2gcIzVGF81uzT6XkHMxJxTrJGntXrBJhTIMi63P1r2VN33whWGQcRkf7Yj
O0kXP26E+A2O6PPjyVpIMVRZUFFXWwxvA9hy9Ld2O47WekfrcE4WlOwh8dgjRQI2
h+64zJBmHW+6dsGwU/1P1eCul/oxnDv6Qqaa9vVuLSZClXJKKs0Xzy9PuIo+oAQo
Q43hQ+eUNjpS/AWUUDAeYWNCMemHPX3tDDrhCxsFpLWf5oggK67Ie3+u0GD6Ko0e
9eEylA8Fisu1i+mhQqshAunZs6hkpPr4K5X/6Ve/iiW7t1AczuZ7YSKsEfATUW8h
XgROAUXhpnq7WDwtsx5pEbPTHUnOs9UvAFEidjIKkYXXLLmhfu1HgVU+NeESx97D
cDcUrb9RwFiRE+MFftC/+ordEoFpsqkgvFfAo8zhsE35+mRVJnkAPYwfjfby8UVK
0SjNk9VKyfCjUorUQg/JTNW65WkpCy5o6iR2xNW4kHK27LcTtSJ28pLrV3Rc2sL8
aACWLpwGaQqYEZLBg3xpY/SN67ucsN1dbuURl2+7QJ7/uQpf47zkceTu+fgmGTM8
dZ8j1yoQSpyNxAqQfruNhs7m5HV0wHUdfBzcK74t+tQHVlcSo6JasRZWU7FoSYnB
Voe1VBioWh0nf+w01XAHzby5UsEF9PG0O2jVP6qQxz6HqqQdzqRg5enlKLG11CJ/
lN8lP0Qj6q4/t20ne1aVvxlwWKCtA/eICCbJvvu6MYNFHF5t94JnA3llL/oZMpAA
cK6QpuGZLjY9MtJj5xeemBVzK/ck9Pc9YOXouC/aNR6yg7hGNqagmuNFhcMFFYSt
cwo0U/5dQowizOe4AE4JvrQQ/aRje1PhzpidkYitiIvNs9CYCwo1TXzEJ6Oof4Wc
W4jXQyUj8WBHjdgo5kF7pfMajQyM9NqBsG94PdTvvls1SO6FOrWWQ9HfLz/pW8rW
P2ScsGtjbxPywsDklJ0rZeSjiwoj/wULlgT8KL8A64GBNKC4Aw+qvGSUdEHaOXug
QijFn65UVVR4Azp7a5nNhJ1q5sssoNzehAIt4VBSFhysZrHsmG5pJ5SslUZVoFnG
Yfa51yAu6R9fRd1vM8CGiAX9mJtQhnGJ/e3c1e9JrK3ZX18SLZrCCtc5YwQblOlx
GgcZgSw/mVJt3OYHTJMBsuG6WMwjHdQkhdeIFArHlufmTxZpFaDHGdRF6pZ1NbhT
hYXNViiPdbDIN18GBCh7WR3rsZDs8zLFXG0ybW129pioYAaTwganI7FmNhVcPxtI
uuPBWFS4sDtWGP+YXWpp0ltmpLS/gZK3qEZv+b5njtTGJ5IWcQGlSFelDvd+FwUD
sASWiZko238H5Fb+7us9WIEilg6oWRLyvgI6aIa+2ZA/a1NmqFJdvomWNx4LQ245
atrwm4IPNNU87q7iWo6cJGh0yiSfIDoa2AbDVEj7V2MGBlySTu9gperNnYk4XmwC
2X7TyJ8q/vlnv9QKrQb036vsQUZZiVVBLElBqSJ3SKDQ1jtvA49KgEl+796EYPot
sBRmdqr+XvTFvG8zUTz9peXAjILzeUBt2V1/l5ck07CJUpMLJGuNZV87OQ5M48y1
q8P9Cd7k9NFODCAt4hNlInqPXxZ2VMfnBc5VD1OA4ezkMXK05hxnBtEN48Rhlb0R
DxwCmKZIo2E1OGLXufIp1pgMr0ORF6kF4BBQKDHdGdezXL4eF2kYszkFuDHoTUkR
6IHHwwQukG9+L99c9F47q0Ya47zpKRGJnJOanrqtcBUSDWMmVPcugYggO2aCJhQn
rBJmDz9lSzOJZCgQVZtdOeAO3Iww3VQE1qf3OSUVV33jfAxeRSzCnTRm+xLYaD5A
Rblmyu7UdtWy+n6NkOt/QeS82x0PMMsWyxn7eCh5P+gaMHkpkQifqNV8wCgK6LPU
YtxQg6aFiZ1EbTe5bv9Q1euZFCIZ6lnzHM947SK1kokImeL1DsUAopedQDF8Wk8D
SdgsnpvS0u/jL1GMYa/Zj4D4qn/p2TUTcguxqWmzBUjYPgVjsaiUj6t8ekLGQS1e
bBsWe3M5UtLE89VNcYGnGhB9XQ6iRne/gTU/nfvkdHxMuROFsfC46hq1zgZ7KOel
4QsG5zLO9teVT2rp6UnFpkeDtSUgZQ4+xK6vyvbc1NwTLhgeC+4aRha7vzu514qz
JoHCwBCoXDafVHoSefFaiGQ8M1hirr+EUWWnTeY68aF4/Hw5LBJfn0S738Z9qRPq
KukPDpDUjQLoZ0Ub2WP301JFnLzsb6qgCv2G5zg59yyopD21yu6LoOsnkEbj+C9c
tG7Flf8h1WYtIAEjseFfaUwI9AcXNPA11duFKmwVTRjDoJsbvEsJ1tOTCMY//zmf
Mt+JaZ7bj7gLpVmiejJmPpVZWKF34mgDkTUartG7y1hN7nDFZNOUriFfP6KdxHEa
EPOuJTplKDPYHiVt2UMyxAPzcD1cCxOx2C39fUAGfk0TzYY0Myezj7MhsJkVIgaY
N2lO8aHSZZAAw3VGsVGLBvl3VJwvq10wu31NkMm3y7xSobbloAtkQa+EJDwCtgdm
q/ru+od+1UZv9Cjp0DaTLRo0Td+4GIvRTyN3/PSbx1bveedabeNqQENhIXtekqc0
f4Ou6APl6yaeFCSmZCUAmUFhfFShxlc0u1FJsmcDSMbLHCE16JK/xpo0HjUP1Xfa
gkLKPSbgzNeyaNAN4UJqKG21ONDV1qvjqtfNDqeWuxhZRNhYFFx5qUIUndc5Obq2
dMnDgNkMValzvYy6fOKvYybxTa0RSJWeQ/DNbsWFNNr9Uq6DZuSFHgws2ckNOiDZ
yJlROTtzJTdlXnnnemOgAVpIc+wwvK92UEdy4plZjdzBScUHIpumViDBC5KA9xsv
i1+D2dgNdn1cPc41KLWahrZdmYjh4/qOvlAMikikiqWob5xMbzDFHE8cqhIoST2X
zsP4xUby685iQqT1bETzK7O/axUZqPAGMJJwODe9ARq6lNlGpJXYTkS0YLefju00
DSxajVlhl6tnmxHXh3C8XsTD8lvwoyA1IrEXot5pIr5eApFFir4Z6inm8cav162t
bIK2n5u91+5ckUdwrPmeKj9weuCATLdWgcP4JVfH7uiTSTCXVVOOLR7R1TBRUPgg
LzH53dx++5hJlZZIVJ9qsGp9kJTvaxZatF1lwn8SkQ5NXGdpW3DeQqyJaczdUQSX
P7AE9+IcDeTFz9gsWE7F7yMYUlcUNlXbcQtTofUvE7h2ma+mDg9wJG665uKKo4gf
JLhLrm0kx2WBDCnoRHZpWHaQQXi7yU2ZN27VR/xVt0UwX9tMhVlXzTv83jVYk2nc
BaFDBbVx/IPHFiHEWVeYglMtI3ea+Wr7pBbVqcXfp2aC1jtF5q/2jvdVZ8GauO1h
FZSpa1Z1C0UzreMyVuSmpbmPcU26/hpp40rCgYAwmOh7Pjx2hp2PKUv2ELegy5oI
R2jjYT7EwU9oLeuQCeB9CL0Wrv2m446pw8CE0OXllpZBnuIk9BrO83GjxmntrZgr
x743A0kD/EHHP4dCCl6SYxR/mPkOhHq24mg6nVnhiQrZGEcDZb8s1I20iIWirmHd
d7yluCfHhBoiwjyOdmRL6fpmcR7JlJhewk6KBU6skeCHlvCjN5qokkiD5IRXeKOe
cIymgCTRFzipZQ7VVvP3n2toMaUfbblRn3uTi4Yf08/lHzI8wSrpWlVU7bfPWlM0
9STbVQWFosSt3WXrjKojuRVfb8ZOPhPxLp0TLaV5vlT46tDeYldhGvvCsneC4dFf
/3ganh1g5k2AN/7qE+vbJflQPFcpU2u78nzgZhv3qA+EFzp116kjsDN8lWZFubMC
zeWgooacPeHePXlmphtjuIYaMRxg+U3qZCjg1JylM/syHY5q8eVznKGr3i5MQ1H9
36tyRzFkQD1tRk5r4fkUwCBVI5fXIYi2ukRZon4IA1XS11pLHYXJilv87X5oxa+L
VMsrqy7sc7rWOED4DfEKovp8YpflrXgxmnrSA2v6OFMECd9siknRuUSnebKcJONs
76CpE/q3rBHpozI9F1n9a4KPNvQQQRQmlj5u4F+Si9Oo/GZc6A5TEPPRa87Wskdy
2VbFguFbOFReyyIkuaxbAKav+EaYzlpQ2adMdiOcG9wwsYXzCQROzz4OOSiymV9j
O/mFqCqnyOe8GYvGnAyfRFRLucBCn2fAcNwhIO1ga6iaTppwdcXGnEchRM/fp05Q
1DLFsIgfrtNMyo5vMzELr9DLv9Qdvz8xp6cKRCasWeKh4u/zh3OkLseyfrn2qrWU
J8Sjt8+SUAJ/Apc2ArS00s5W1/u+kmP3eNurJSo57XeKsC0jPgF7WOwFP4oEm3AJ
zjHJSHAmWSsfCvdijv4KyLw2DuIyRU9Mf/ecEeaWEBDDs+rUIZSkAPjRj4VlKL55
GTP387u59r3iMQuMKkVY18WImAWZYD9erGxzwPbfC6IUlxFxBb2/66NcIVOpc2X+
6fOi9TzZzv2UScAah2mBItbecqYMTzUeVIOqfba6PfPiMCGAGc5pq/0Oyey/sW70
a3oRmZdJuo7qVMqeFT6ib5YsnlU84eQ8rvezkOXspux2fy5UFWmdDZxwRNeOKCCF
xbPSEdXfY4gXBd8Y2cLIEnDzy6Y7yoxONCylXUlVUhM6LrHRQ32AhF2gA+pUCepm
w2YbAIlNMUxR6da3ey7y0SsideoZB4Ckd+/KZMK607xYbSaDyLFGAuDBBNCw1WfP
4/YELHuRunxjABc02TFQOjKklbEgHyzvzXeHua6YLqLVD9wCOL5/noVHzPhnCsPO
D7Ooj+8vQtgGgkbJHHatJUhvF5iydGzRqi819mu+6grxtUg9T5OeWJvY1LkYu1tN
kyZ2R1DJ62sK+G1J8vVHMl4gtNlSsfv1kEJQjueI3cBkQwzW4qm7526ITjUSIZJH
NvuDDElxvoQONU6mV8O+P7TI4gaxyiPYH2kD6WUAK6CYGtZA2wqtQxinkyJzhikb
wKY6plXc257WNXRMslQy1WGB6jABY2/JZW3QxGQAJpYDLlo0d5O075XD0SDBPRhH
W2wWGCSM6htT7UCbu5+KeorqskrV+u1+rPLDKe3pq07nu/mJAjObsXKtk/avdtzg
R5MQaxMkQyBqadrttpOcLLuAvSPA710tjYFr+3+jwr/fRb6+YjimWJUZDd5MGCAq
RQFaxLJM/c/GbvTSs98gGw34hozRb5MjLhWe5Ya6Lbu9hQ7qEHx37+lRSvCtxsKk
GF1lEdXBvTYT/8IQC/aUjXO2WGN7yXmsi2k1/fT/X/daHTub9XLLW4/8V447UOaj
4kfV91xaIHB4zt88XKQJXqRJPZIq/oP5u1UQ6yM+e5KvQ4/2ShU9E5A+R5qIiM1e
ptPMUFCiJBF400N34ZDwsnLXH1ANDVayNBP2S9XiOp+QsB7+qismcOq1SrdDsUWz
bLzN2JeOWW20XYTvrY9la+ftjmcabE9RQ67CS8CRhasikR8jBzj18eq/S5ruPPgj
FYzoZMLlpgczeJ1t69YAVLi/wv9bdutvh1O8t7waNOSbSiGARzUY6ju61v7ue9vV
JCGEns09QTzGM8kHwYcVVuA+RAqk23WdZMjBhowG9FiRkQiXtLTNOPBhkri2eyvB
7foW9eoDqIuDP7tEBHwSXRmZfoiwLoxAaoyMyEBj4uWNyJcDDOvaw9O4f6PsrxuI
vEn9mpBsLQIpUyBd8qnUYHFPp1yk177moA7b4Gj0eRGO5DkrNbNLDMhKsXGxo+pi
SGTeGYaREnO6nkMnRqFo5xwoZQI0TtAk+0ioCODqAra5PJRKmkQ4o0hy8gETTXCc
z5kXYh4HSiFZm0HiI19RS95AmwipXP7uRffeyDSe0h4zQiHJjLOUcdlunf2x9d/S
ZPJZV0+3P0d5h21jWDW6ikWkKCCoQeJ9Oqg2xgXpMuUdonSbucL/PLrJzYhUn/XR
1zFxT+fmKQaUP5/KqOm2pTpZj41wiLparccDKQnUc1AC7Tf97YWcAX+Z5Be0DhCs
FwgU0dOi31NSaLRyUmI35C2wH8IkqRvb2YsRLvVU+m/NtDtnwmNXqGJFCpE7Bxxc
AGp7aQj3BHDddxSrluGz7N8m4CVeH1V0mbCa2gAvcxpCNrOORJjc+F9/4j6LFVsh
bHA1HMGazJAWAQdGLpretIII1J7Uhm9zLhZcUcaVdJwJwaDheia+OJkHDmtHicC7
bmANNGd8wWtBmd1xhPB871efmTzvfXY1MreCWonI60r/p9v3VotFNiOLPiulMY33
AfC/jY/FKVg+GMW/yt/FkUazAHusxTqiy+o33/zbOgm8jLsCEevhrTsyrY+jwSQ9
Vcm1ExDWPXlkTQL75F3PcQfpXu3QbxVYKEJxGQsd5fvf6jUQss7x6v6z9kXomv8F
5y3MCV3M1Rv91Z8hj2JDpPRI+lY2WgcMDPGkqOJ+TICkoI+LYq2aw8MJvmYpBqJ3
gKjzTSov8r8YVeTTk1NaN+b2Lk3EbLJOEDXRgCRpwiJXCDDQ27PMFmGSFuuvdN7g
/aoZWevddq5ig0mYjY7k+Nafj2IMUvjmzR3Q+PBz8ErHKWrs7zSmrZQEpcnHW3g+
4unfjrtB9qbgxeAk7KR3GJR8oJAONWQaaYNG5XktVIdXxKAFSowJ5zHzHYS0MdPa
jLwdPXj5VA6l+XlEjT8rJ2WjzxL+z3B4pYDGZ4spjwIq1VKZDpeXS1gSHTNImAIp
A96VeruN4uvEyger5AYKfv/UGmqk1P78mOT7NHYShlK0J7fWwmISrrN2OB2zMiHB
m8RPlbNBvtMPE8+YqdyLRYROoXU+2CbjEkKrGDUyGcA5JWLX1l8T1JDPD+kGI9Mh
glQlelP3tHx6ta+bHH3Jqh83mzbUpdd2xIMZw0AhyJS6hIiLLOTdY6qqvhAxFMqd
92dOqcQxMAMrxInRkvagekNk4KBIYW1lOMBpkxGiFAbRD8jyyCp6nbTtaOJMO/tm
ImcxAyl40FryXaQd2S5C6rAhjYVEV/0D6zG4MK6lvbpI5X4+slxJUEt2DXz+93Wf
zc4jqivjCEiMOdFIxWDayUgds3pwnwcxdF9PPmmxYwxnLUxgPkUB684/LHZj1ieY
w4grHdq6dzgVeDDWy56069Cf+jPVd/KM6LNcrhjQ04y+6QJrhzTXFdVRS1aPzwYH
tgKwa41hGhZqKECDWefcs2RpgI8QfYvmdWs3B+4v5UDtLGcbOfaP9mct1DH7oaEi
+S5UapafZgIKehqBmEuVUcG7O48kcXvGmRCMTkvwpy7b2OGNBEDz+/pbRUApyaIh
hSAxByt9pCNJoKzMoJidhj+nJIPH9nOFJxi8eYxyFnYvzSAKUOimKdVYc5IGEWXs
lf/vGYXmRvZMB7IxgVT1mMKkca6OooUpL89hs5B6bUF9uB7KkBglrSlQb/jWAvPH
gek6TF42FvXy1nlZc/RO8uiYzxLRSKtIDonEk08wdzz9dwDPz9RZcudSC5nXgplS
fyXJDg2+PbB184mqTqcgUdRolTriGvywKK7XfzHwrsWKpTIkwasdkgXg1JFYUf8/
gwjEcClPnyJuv2wO25WrIt4RtCGakkTZFBPF2jWBG7Y40PHZrk/QmkRbVpgYwU6X
LnU+8sAvR7Ynzgmqyrmdkt81RUEnw1ZjpRebit3WzKt23c94jxHNJHcjXK54rZ2p
t6rSOv0jRkDXbLp0NI+hJSOijjFqmEK1A8X0ihc9hkJFmKs57K6PmvrsPMnfiHwr
CKJmpvwqxOUjF0TRkt0nTXljYFj5elG0gKWWSzXFLIUqRsfaXWgUsbpEbBoPpC5t
5K9pRuC+mJPEW8jraRORoIE/0a/3q7lRxHWvl8Z7YomePVYVfr2sFZ5bm+yL3zv2
ROhFsnphvFJ8ifqzfm96VZLDZClZNMHhenyPQDfCz2WC9ZNQIzXHvguV5A9WH0Ev
YRZzf/y6htryxNgjbmYfKKqCi/HBHNf49QMqLJ68/6gCxkaxi5P4jCtE5YJUktei
pNPyU7FZ7tePJT3A17qpAXhzSTjLOdF3WF3fnF5KPusYi354RDI8UGY8s5fwO5/h
GZekUmcyUSb3pQqOb24LH9tsUiZwP524+1C39iV8l1qzy6BqTJyIUxJrzywipjB8
g4iUp6dWaHLjOWQRtzbSX9/ey/ObsIt0JNWcbMuZuAw8AYqfXQiZ/tboTb8aY4D7
DYpUF9EUTh+zyx32n8INGIm22+sxXpsZmwu0GEjuELJnpbi5JjUBaWgVBkGEI99K
kJ7NIOM5H+MYQr0ZAvgiZDGe4UwlxJTKIbiqDikcu02UpMgNihu61uQU0MW+kbSZ
rFV26zlz+fo9cY6IwGi3eq+oOBkp1GrUNmpcwYoz2hPO2jDY13ZjwHA/hB0GOQwk
9VW64qXQwRR+M/KrlB9EG+GqH8Y93VL3VFdjklNJbslUnwczEZSyiJH9eJqMkGlP
4yUfXED/HppBkgMjwx0/zLYrhyNCZJc53tkFMT44cPDmqzrKj1wvdsSUNUMOPo6D
vnMuG7gC/RD08h1efqKQ8X5pWsdY9OewQ3AzBN7E15BzBifmG8qDio8iOBBp/3AI
i5fVFhN0mO3GVG0dCchTIhr5yQYvjJ0Q/TCau/ntPXZQle402pGcBf8rqVVOLBBG
HLiOpChkDciJr4cPqGuTGD8GgLWTixrWsa9Ei2Eiyh9EAOpa1u1jO8raEqqi+jCM
59vGbRqkRxk91AJkJ/LCQ2u31iRsZ+6ccvZnleIOtPablJ8DF3EYPqhtR0XdAfDv
ZdK0V5kMTVN1tJ8Ex8Rui0XvQP/PjuiPlKQKfSrSsqfaJ5qhEJ14aRFBS4LOx+NW
W5hCiJDmnR3sy8OX7LTQkPGd5zmYGWnYwzNMMpo3Cj5Ywrh0XKzcLgoT7OvnIR7V
d2YN1lCJjnOTfyGHjehnNuFF6qWledVb5/VbvPdXH3xZE3ICXosEK6OAkf0UTsAH
TRVcBIQwsMEsO47YA4Iu0BsdjfNAVpg8H9O9A5NwzRlnZmBxPReSN75DbOrDCPB+
tiF8yk6T3K6z+uYfypn82Kuk19XWrJgp09iPC75FhMWuad7VJkhscZh54Qs0lBtc
nGRmpm3x7+u7m0iFPwXS3K7RYPFjz0ajhn4k5uOgaan3//CmFd1vF7EbE7RRMNSe
TRPUejtfld88nvu2OCF4JhNfiOtIzWYCdzBBn/5hxxG5Nk351EEq/JLqKcz/8R0f
x9gHDySFb7SSQEph5L2z0RVmiz+rkwsOJ/X4cjP1ZwSFllz5Ip0V/lHDLvfoiCFw
n00wPhzQChmsDBsv00qu3bO/eXG2Y4tRpCHaV8YsMoRCJy7W6MncI8hZjby5sByX
K7+pMtzSkqFwQRmoVl2Of9VcctN14ohE1fOMChl1OxP7u1AI4y8NP2+ax+tQFxdr
SXKRZaM1OnBjcS066fiZVT+nid92ZRHJQDLJADR1a93qyGykJ48z9TXEg4dc5bLk
2+5KO/W9G8vyWJT2UdlbUEFPLuU8Cib4oDydSYziqIFRWMmTUCr5u1YaWC3tW0uh
a7IzeE+ve6XktE82mpaW+/dPCCEXBU0LOdlYQPjwQhgDrBh+W95WKdvDbeZxNy7C
0NCAnYucEom1zmm98JaojNx+ClcLRz+I6kX3NS5kBsjwd543xBIue0GYEHvdBkpJ
3sEK8DYnLeAEyomE7pPVT/GSJ/Qehrd5/0xZp1TKF99/Iw0nkPdElin95XwKRlGf
rwxVagMeyAeG+NIOKeduigJOgXXWeOwqQMs6Q2tJxxLqUBe+HeGy6uO23egIG6Pl
epCXIoIFs7J+cke74oDMx8D2xYo92uAE6VRogWXGhQZzPuuc5MQbecz0xjF+y4L4
3HxLZoSviG4N3GJ6vGvG5hjzirzUvbOynDtY8YfB7ruKNOBMbYW/PfSFjhzqTO1Q
fxBDHS/cICfSH2vQ86tTAdZVZffbySdWucYMiT/pbEaHCgYgjP32Fv8GTd2MpV3x
0w815UvHAVnK5znWcb/SEAyuN3pSi7uxNaBsM6hJFpSiVjZ+yYJfUjXg7sVaJkJc
snFoGpo3u5PJVijQKKcOjhuHikZveNucHVU+K8kuHDebDao8p96qqv0UrFVWGrKt
mV1WiKLT8Rv2l6tG3M/WM7jXikLco0opC02Rb12oO6Dm93XyZQQPM6lJiFUMhsk8
+fejOH3xxnAgpUMcbj9ntyNDSdipDDeM80sWIcnAlz3oiPX+zXd7AdcAYiddRk1Y
3EgJx51xv6Mb0XJ3RNd25GtyuQuXoTVpRF2sf8u/8zrKf72AtN7C+cxUuTwaVHC/
OEpXHBKbqzAk9yjOIP6oKSevZfqTDlv0d5NTtNXjA8zvIODssl1vwzAOGyJZi6GL
2xL1RPyNQCMaom4W14X8cbzIOQ9FbGUcHGqUNWGZ84XWtKPifBZyTdadY/eKAGPO
P6PtV1dKWvWkHmMHoVXPaiE1X9q4vX2k5na+3hka6tugRZbi55VK8aDptXM8Acjw
rNh7HPhCrgrHq+IsmVUFunIXRIKiD0mCzpycog49mTkrjmWK/ZM5Zj2f1pwHXELk
4ieGOnABWBBV+ctnnaClFNObcZtiKu+ilHlj4IcuN4PbmV2ryyyFh1M5dKXOvAVX
vVkunwicDB7hBLB0FJoAi7qw3A/nyTNUxBreY6qKHw+CAtjkIQq917HTEplzG+Nw
zK9eXvI2MTkmUl2t4bsi6MkZbk3YkEhEupL8KRM4bUHDneyzVPYSFi47U9D5DO8+
1ecavuJgb2tWcTTtQQ4o+F1SmGdDHoRQivTrAGtKEmOmKC3DZocRBXOL0T2O+9ev
icLFJVUytu7/XE3RmYp0Mln71+bGwmTR6ldjYjfHKGJbpAj3Yb1RzXQ9A1sgwN1v
jvhqzGKjUfSD9hjwPtYIg+04eI7vY+ESX8cdcsQOnZzvBrK8NIPkZFBOHgRbu4AN
GHyeBJOWQ4gXPhhML2WSqN+1FeqyHpbcofBVF8nL2uHrKRa7RBMaQ9S4vg8rqh7c
8FgfLuuhfoJbjz3tlADQkIXF2UlwaCP/eCEwPnBOHNbedNg6HlWzIEjKSqZyDmIz
WowWOVIW4SRcA7eaDr/hbod5AItpLIZDUX5gEHKdWTKlE8f1OLcmd5E80VxY1h/n
4UII8VrTbXfUrOygHdizB/Kdij4Bnz835qOhhD43Y8rZpJjc383/LHDixmJoS2ii
2pYauKD6LP24knTyg/zYAowiweTk1cZDuDkQafLg7S00Nl2rl5I3/VEZvdWyBtrH
78SHqOz4dHXHTObV7AZByDfgITMUZIC9UYPpfBHrel/5n2tcdO9uYi9y68GmzpWv
36vDE1ITnv9XwQ/yxq9SDClwqckk61cHiuq18I7VMtbwvH+4NLlaNPEqvoGPV4jT
ZfFd7mTKJjcqUOlBsZx+wjX/drhGP36sQUE0vs2m2ULoOZu48fJUeWzkvauGW4r8
XE6NYly6hNmmIaf++S9BvjA+NeqnP0eNLSkOO9/fe/h3ai9VuRvEpP/YMAHRnDZ1
sA+HhgfUa/poGNeS18vzZ/joiaibguepbCjyl06LPp9cQ+qvfX44Q4bpMjhy2deD
TgdpkMYrnPh+Crbf0KRT5HeTBS2SW7iGMQRnFyLxcn1kSnd2huoDs8/CIJD9TY62
ogThXBgO1rDG2QfbuZAocgD7lgWmXQYRraXt4bulnOGEQsVEIAtM+vUo6FONf8PG
ufLHJ0ZPHL+Ars4j2EVNCGYhhQBy6qYIwwLqfhO/nGe/pV0xmCdjnUQOKSmEjWCY
NfCvpZepA3vZfdrdecDhXVNJc/L4X05CZ/+Oe/CkVVw4GWw+KtYLDpaHqXnvLKSF
tHNpdaHEvPxqxAoyfyFIO9WVQjcpLN2wlTos7GM8Yd6AF9b648Mv2EIh2VffUn5x
3mA8tX6lrazY+utQ/AQHEPujgIiRBItwpQEssxCGF7RlVsJXUpfCOG8fb1zbTkcC
IruSNVoPVDLINPfZfGCd1jsYVgvW04wlBW3yVDdQxRx1DC3BGEOitE3hXrehwbFa
GaXT8jEiClptNkat+mEVrKXCuP3MFx7HvIKmz+VygypFuukV6xB8+BcK/JHoxbaZ
JTPd5MzSayza4X89tIcY/TyLPi12R5iHCHX9zR9us0q16onvMxSIIrbkbnb4RWg5
NNPudgDo5nWSwwBe0tvVpRvxdI3XCqn7xOaFOdPATrue0Ar4Eo9F83M6/v/hRXBL
1OJ4D2fJV46vfurOmZBYqG/n1qn5aXXdEqfik7cw3zxH0X9UuvWbNTaGz1EsdTEt
koVc2oMAOy/asv04TGk90V1xfg0H1zesEHaaxP+PM/WHfajiLRzUHg4epbxsD1Dz
/w6bZn57W0IzwgucMOdxQ5aKVuSpQWzh+40+hCtCDI8RETPk9xTL+TGcYJY7ed+o
qkwLcm3kLOhd64KCqX00N8LWnrmNIvazzlw/dTxDz5eWw5Mj2vFAzMnBz4ZwoBI/
yDW38CzIIKrgLdzWVPeM+DzJFnW3bV+07Ev8DS/olXQNkabIBoR4FSqhF6FHJWHT
LiQXIqBiBF3R0H788Ay6BDdbRN95mKuqyxjVdlx+gE1G0AgDZ7f6CZPdWmNjGNfg
PQuovgFSYThbnHIpM2p1rKDj17t4A0cZNVklxoIGvnldmd5FAkuJuC/pdUPjaYWH
UK0LCGx/6aVFl5Kba7eJEVx4Cm2iHmAOmQDhrlvmumF6Z1Cr8H4GHqfN+0zwmmzG
qjj2CRgWhKToAJrhjAN4ffNHJzBg7CLBH+9ntAu0NHXhvL+SN88ICs0BmIx36oT1
7T5QBVm7tRGM1rAdjwsPKptY6YhYrCJ03GLeE9klADkRMq7ZTOrmygpc3GD7TwOu
EXBND408Te0d6ooN3P5IZ4nRgnWyznWL5mn6hZyhEXv9ps30mD8qJ39dByBUgQ5G
vozLOVM9ZEV4Fe3HGtEBx23jfNGy0lWouKTOMUXJLXTg6kMX0BalOuugD5Iq4Xvh
Z9I6odj8dHOuQpA4GwFY/2LWY61BB8AzdOYs2xokMZZibQZP7F0GZhxrdphpwlTZ
1xO2QJ4WkXTPe7OWUzazBJpzgNOmbAiHV9iC6Z0e113YRfM7MOA7Vjp7KsN33p3r
58tE8YFJUzuYa58ikS/rKlUffrsvc/gkT8EY6s00JrVQbFsBObqzk1HaSxNw+yP+
VRd66a8GeUCah863J0MN/7LHOvUNq2R2BgS92d5RajLWoSim1lehUzMNeYMfDbmU
4HW+qSuzjrFhMYHfM6tAVK9kklVvWTOFOqtz9XkhKPJIBHUIr114A9TxQuHv0HjS
KEpU+X2CuXUvm7cG2daz7GlcKzLlmDVFNphnfKqD3W0xd0D8G6fOuHJiD4YZ6Xb1
2IaZd52Uwory5mW9cWNW9TdYOMoOEPk8mQ4E04Zw2m/syJIzd9pyHed/WRD3MMrc
kxra2GGP3eL1zpON4w9FnTKLVfq+SoDl432u9GG6ecn/hDCoKvte71NhlR2mVyNi
JvRgaU8KvobH0QkFivMn2f8bNj4TTZhEMtgtoqrBf0HIWI+NQas/2e6G4vDddCpH
N0QnuzolQWF0h+/YbcWlmZqyChd+d//ZrqrEpPcLb+vqK21qZR+ilidkQC8KMSwL
2+5MARioBH6KV7MTLg1M/1Qmnxb7xsAvEQbx2Gk/vPbKJa9IRpzq5/ncXC61U9WF
kdMyJ70DMv2nmc/9D5g1ED8UK3KK84Ef7RSfheNTt52Vme5/bH2sqmqq1ZXUtF2S
ftiMF/wYQRStuYJNTUCo2O3D9Q9N5S8kE+xl3B/UBRjkGHYAzrrgamQag8+Mi9CT
iSt6GEdqblkENXbgb5pPQHZKGeS5Uv9cDWxN8ITXSpZoLf0FpTTlruBhCZ+0m+Vz
PB6av2gtEfdPBKhfWgRd/PGfyqywQZVYrAKewbXvwA6LOvcN37AHS2onwBGNjlhR
XzuoB1+pAMLIg9CFpc6r56G5OH3SnmRtNc6LSzYSJ4wsAMxwuzs8XkMk2SYr5v7v
68C2dWm9uW5wNzNGiowM+2YT55VO9fYquWqfXbzCWZtiLRdT1Co2Wp6d4bg6GZ6F
jkKwRiGPm6+d4uMI9BtpQ/duScYYfDljQsa2pi4XZa9Yl1O/suz74gNmF0oIDjVm
TrIhsgTHlvCZBQ+9Rnd4q78T5FNA4Klz6uNOAdNO3FDAgcphDaOSWGVvHRuQS5NH
J4r914+YV+7XjdUgYA/Zruyxsa8//F20nEbwo2KKjmtogepymKK59ccAlyZtkZw3
839CcyikBetkc0K/Dwlk1vfh4AYTe4eg4vUmPse6yhdnxLQHnPdspw1eMEf7tzJl
tdkE9J/jQQc+FgVpDVKYN8umH8tc1M6vyqgoSZxRX7gJoTndGvKlEFC/eahQf3mI
O93LKIxNMf0UGWYN90HBU9p3sgFezxZDk58Rb+nxn7F6dFc63j+eb9iLCIaBVy41
7ybVStlFVHb17jzjMar9cBRM0avuhKgYaT5dQQBwcq4tQxDk/H4rOPsYLGKyQ8lr
z9kTkRyPiyFl8LgixOvVwiWXrBD0oOKE7srAneU9Oz7ec2Mw2ghqDjfI20Q1gNJb
ufLljhEXRIsn3wv/AfmMovDT3f50dvkwofKHGtj/+so+0a/1SiTP36tRtMZ8lmk3
29+qG5jj4dkjKl2CPDlOSevvVTrSGCIZ8JKn7aJ77ISdRSJbcH4SZTKmQ8LF6LAw
eNzxAPQBuYq3FowELw3gZR7Fatetz+/kcz42W1Kf6IbIbU4c+f0vjeNfdtLBqOTi
BmEiVfHjtKqMMn9C3k2DBnns5FU5UyHli0I+6hokHJNdryn/hNKPWr+fygqj22Ad
rpt9m7B1Ao99Ll8e/veC60F94P0cPJGAQlHH8eHnXOJZlDA5H17SMw519awIcth2
0vsLuGdqLMiO/PyPEjet3pEx4XYYyd+PCtLF6x7r31k7CwzpPOlYfcxNRUobqTpT
pH9bmO98r14FkgV6gtlX/xvXkCUqyAcDPtlyKWEoAkcALjuBTbmKZJ3wxedjom2y
6PC2hw5FD0av2GJNXbE4o0Ny77VOGeiRv0QOlODN9Vae7Bxya/qgFNmPY6u5104V
9I+x5lIwuaYU+Xpibcgns3DlNB09Xj/uen2s3DBS352qpiS6LsT61jV/Yy+7tm1B
/WMqV1w5dygyvr/qmFC9HLLlurCfwayWDcb2cnCF9cit2GyewJAQuC1wRX7XRjw4
XYXGEx/49fkmSjTkv0qFilhxzlwQ5l6d1MkM/aSm3cKzSWYdY7MS8bGryUk1VEdF
SoYLQgZWVWzZODG1Z3mVavDz3eEM7GN9pCb9hUIAjtcBxPqBWfV4l9fLssEXvGnu
m8/IdXfGpLZ4zDq0oNqtPwkkuYQc2jIi5mM/5lr4lUKnm/3WWTiqyqpOpHFZnBoX
/aFYSZWfflqdgnM065VoWDoGR7iZmnHEUe3eB58W3yfG6OBhCOCs+vf7DYGPyQMT
P7vuqGyOY3Mu7e+PWu3UA7O5mxPqkUorWTecnI4kiJc/3HotAj3VZRtFpYwWNJJF
GJJKIFad6ljOP5KTJkQsCn1LHlWxqAcjCfp+dS1vizRgbz1Luo9/eQYqU3J26h5L
2nE6PfgBffwnNC0PTSqkMv0GvmtKOTdhv5W20F47Kq2DZOY+XorBcTLjnoYG4wz2
ghAdc2hZXSugRE2lb2TKdu4cXsB8NmyPN+SzSXuONmNZ0+qyhVshqehNWddM/DvT
FWGOmzCr80VLCyZXJWQ8QwgBYEQdaqQSCJC9hvarSC8txr8b0CkTbcMwsQ1ZY4Gx
GTgv8G5BCgXfF+28H/u1o1PwPOfi7EPS3D741LU7r0noVgF12vY/eooj4aQSqSdH
Fwqkwqw4mbzSBfzWA6nu+tO/BN1GokqE+5iKu7ugmSRxcHNQ6z8HcSX1Cp1qTyD5
DAok5TFxaxceT7TsV6YQPaHax+7qYNHgDkNXSQOanHgjTi+oK/+k6A0i5N8PLw6U
LQM498zj68hnlhS2qMwHNelCBr7B7fKa7jykLqUhuqcrZ6d387ANRrCWQQdrfE0U
uKCiraQCqHPHjv/HExhQKvg76QHE6IUJGUUEi/wLxc2+bCnUbFrkylyDZQQ6X82I
v71Yc/G5NkcjIRedrq1sgyngVi49bfOjDQHoZfK4pt6rMV1xvKrsWNqHiqTGNpNz
uJKK9TPhnHBSR9anuFu6Q44io4Hr0+t0/jQDp7qCjqKUoDWNfiAIKv/IF+hTCBut
eABpYMuOKyDS2BD0ycbjeFsV6Pu9cO1PK1ibQmyoYKpjLzFRw3pf50MWCXbC7qx7
ws8RqE5jfWQU3isGrKreO2SmPFVef7tvtVak8RJ/gIobm8t682NNQzPIgtrpxGwj
zAyMh1/QVpEUdcvcMsKgYZBskx3tb1dlhrwOEibyoNX/P8tEWxEdcm7RiDJVrwNl
4NstwJzUY2Jc+N2VmdexZcIEJ5fvVBvh1MvoAF5xJK8ADSOUmG4ALwqtcQM6v+rN
pJVmwn7rqDtv3Lk6jXx8LFX5gVkn1E+wxvbun870PemxNZxZ+rsNB+BpImqnotuN
e6+wwzte85jomV8QiMrHhU/LoR0o3IJ2MyG+vBWRlaeuO6Bst28g5LHcs2ytxhzG
ydpTjPRN6/aW/X7DscKM8lkbWD8KvzlEQBOzG5W9F+Rx6OZXHO9lRirDbc/wN1Nr
4H3JHbHqydRnstzCK4CuAeoMMCOo20itx1crgAX3dFGKneX9h4y3t3yV++WdX+MO
0rARY30CZUc9f6Uo+uoBGpGAhDp21Wd8DF0cGA7GtepPI9pF5hiFNfPH4hFYQ8Jk
/pFWIFX6PYsS7kggBkCqK+QP1gNgBva3RZFpp25yoKeKWs4JqnNLKEL61/VF+dVl
1zmyOO6sUD7PakXYwn2+xEl7AiPrMa3f9+MEMACmwPboqp80/hRyL5WurHLAoAxf
7Mrubr53NbxjpnhAnQmynU6j9URQIqwZO5XONhd24eHjwNPYlu/u4J0bhuu+UOHl
LWM670abT1U6RoviIpOfYAN+T7kWC+ep1PGZpyHdr6iFtCkA37+YpdVyigb3pZLf
LNHSpfLbzb3y/VLNWBybHO4Ip87xLS7yx6qDKyJw01JVTn/2TsA/hj5PnB3/QpQI
RAs1gFuDDdS33rkl04oTfV9m2wpRcYVINorpA3w+xGO2QI9nBuPrSfw/vfoUtlXb
l/NXENhg43hz6kuYqw9AtRiG1QnQkavKLp993NjRpFqP4Nmbj3287/Lkxvf7Ryt4
Hhx1AbSx5aXSZCYyEEJx08al03/Zv802NnS7dlfvpT5JWfvxWNqbw1Q9zXq/Jm1e
1HeGn2Q9ar1yoLpObhDDNdUrvVt3M9twHkMAnDgJegHmxmzq8wJzWpi8hrLeM89H
cFiQPsCHyY2XnmHzvYISb94nQbu1hTaxk2bWh/jrHGbP9+f6xJLqqWc2WLbP+MUe
LsM1sHmjqxJvBeIAg5MQFcWRBXsZQg9r2+i0TrQ49cj68fXKrs/ybSDaBIX9BPjf
k1KNBKyMCALO+xrj4q+ehM8XdX+jS09tf5XUu/BzP7SSjwuKk2pn5GrO/jj4AIKk
N1E/coNo9iqtiqNAASkvGdpTAcPwB3iDRIJ/QW0o9jm6pIiy4K7m72wAwo/BX+ap
Bsh7yXD8MVgcQyFunUr3WPdGe+KcGUSr4bjD0wEi62STcsQPlpHbmwOq6EaiGfpH
hPyIMIJYAqYzN6IPaQzYbAQzy8JriyVYtvJaM4Z+OSSPUCAismiRzyVS865rQQj3
qdZ4t+RXm6oe2WBbnREKJ8pMw6/iO7ewMqntvN+rIuOuhXMrD+5VWc6WOc6xN1Lo
ZCIKv15M8tQj6lPfVwOcVPdLVhpMofv7P/f5EL48oC6+QPKS3PLlsRmDDM1WP3Sk
KK1p+8Sa3TtfO06PTnec2gXuxnbo87N6JuC327EgbKUwPZM6wStjWdYBVOt4o9F5
GDtc6ftoz8MgTNYbU8PYM7vhHv6K7u1O21yr919PCSGD8E3Hjhj9uU+zSzmt+NQb
TlTByqlVpEPR8tJRDRG7i0obbF6kR2N8Azb+hONBHStDd35mPe1tU/yc3G5HqNrK
whB6dvInvH1PsUEXe2ZWdrJgdezVvATyKRzEoQVKsAl3faARQ+Vre8XmLLFXoZXl
g72IyaBYTiulY8dW3mn5ImQLcJq+/CHi4fy8CqNFR/aBHgMkkEUR4m2nDEpvIw8V
EQQE39s8YdBCfRwvonwk5vF4f2bd/2Q322ZyCpO7977qAFxrDEso+HC7xkvjaVBf
rMpK0DYKZ2yEYBiAbRjiqVeo6AjL/TF/d49s9V/K8A9aTlS1d6TdWy7implecFXc
60tDMct261DuLDb9fbVExqKaFJL3m8Cl/0ksVGYonHBN1tyqLYMBEBTqHjdYjgh4
4OB4V94zw2kr8ZTfHW5h8YKc0iahEi1BXXcr75FTEPK7My1iz0NVZjix3P4Pbp3Q
SKWtcmIATFKhZPk3DKeIdD8HWh8Uhp0/zZ84SJGn4x/jMynniIvoz/4mxJvFVbYB
vxFzKbBYcsLJZX9dkfg6ydf++5zqH7GuMW389TvyxNyvHatLchSGiN1JyzFTBRho
vcVwVbPlCjgSQoW0Qu5Va2xfjJK6tL/EyMyCFOyIRTqdMflo8xSi7YVkVTkRkacb
60t6JZ6wraQQOyv+1QA8QoLTn1sL5O0ypyEceFrnWSyyRZ2zT7SD7Hrkglb8LPyR
1ErG0XwyH5xNyN2cCRKYqBpcMRwKIcWAoYjHGaBVbZoo0fsHgtskNjh28pPRJ3Xh
1IcR2DxMeuiDsfC+0COZNBikiEEF3EttmAG+HdHM4cs8XCv0QQ0Bfet8A95adPml
RUc9jBmJmE3eye/n66DnOzuJkVAKfIO5o55/if3pr1INNzFnpk3ya8vWBrlAtyZ9
Wqku10ksJv4RyfQNAAySGkLJtvPzspw49hovS1UM2Q/0HLoicCoQYQOwiasi3UDt
ylv4cUb0h0SeLz76vdV5ppkHEBORnwUUOqaktmSmr1HvFRaFtJBvcSyQGUDxjXkR
zK60vRqe4NbNPLpbWPrLAhyiO5UwFO8kDn+9YikRvY2+NuQnRli1e+IWD0cpTbDr
o/xrIeQmj8Y0JqdbW2QCFfjGFef+Y9lICedhLirEdICUh+xIx6o3p5EnlQPzjZ82
WNwd032UuzsapqDu4uudn7DazBCY3GWTY5MrA62euTF2Rman7hu9yI2DeIDYLbOY
YYDF8Rydh84tuIVQOZapVcF6KcKkB8Y6a/s9K753EWSnjIFv/f+/iacbFaxR5Q5E
Xn2arhMHiuunnbNC8SARa9vuENiACSySzIcNHG1nLmG9moGsVJP+Df5agd99/iXN
nK7Br/KeKndH7O2MJvz4na1dLu2nIIjkmMLD5XHJ/1589hHMM13tkW+FI0lNio45
/C6InHT8queImvc+mANcJD3IAbXqv3k3I6ZwUdcLqMlVZg+HKUuwx9K4hffBi4Wo
OfbZNY9pJA/KFp92ttWFy7pYEKJ8q80QvDT2yIm9uHCHNGJh+/UH1jPSFGckBz4b
mHpD+EbWABnVSQICWZFERw9CS43q9NRAuB+i/Cxr9Vv/mHgNSLHmVEjqQXta059H
OLT86t0AM7OdU6oQpWmLjtcMG6ibB2DdvtSSaNt8yXYv7nDDCMoYJS9WiqzOPrsF
lhuRAWBP0E00/sLesn8BlS1U4bNGEEQW6NOyZtPZ1Hr/DbwB57vGXNsfYFdS1xJ2
TentcFI1OxLoJ7xhhqm4vQRwXVd7POkA2CNHM3qQXVqX1djy8DdPBRfrayuAebVD
NEFX33b3g0g/wnIVjVLxsrkDMyVVUIHaSD8Bshn72gjZzSv4e7eYoRQj/a7J2RAx
QcpBesy1jGVamWj3yLWTtcHaf/IO+iCkuRTmKWHBrPqn/b1zP311KHzwb4ySLWxO
ir5imG5FDl1bkASI2oQBpmUZLezDGxslCCJEMJyv09y5D/TbmzR11ry/FTnuhGVp
jksUMX9+Q/bKveZm0Wb5mFG9ieBUg5VlN56aIuyVF7B1TSdudcmByif6LvJGe5D2
soZ1FH6SFQ9L1YSMBaupoN89Q8eJs31gI8YGzwI/lulTQEP/mpZgr+ZZYWIiAzY/
g/o1l3xp762oTFOHeHGE1wwxPBOif9lnedelVLM6DCS4cmg0qL8dHrY2m22HMgeO
Htjtz9jzGz0G/8e7m1wPD/krUupcA3ebF/zxVQwMnE8pD/lu5OXJzPmQJCfqYupe
z8WH6I5tl7qKapUMByrakfeRTqlEdB5D3eXIghgH14dyISTRQEK05t8ikSHSpkQP
JCqBmYjuwdPcyUgW8hUeksVy7fPnCZ5yZMpfHbXYflewnS+KFEjPWypeNpT562yR
sk0jnQyHafLdYISgGImzyJ27IU523KUbmDGXcNCsPBfv9nZmDmplvD/pKAVzQ4lf
njFfKc9Lemw8g24g1LCWHIDSJWh7t/YtQ5l1J4zqQ8jfx8feSSEyw8bcVESmw3xj
AD++yVHJ1SuUw/eZkRnze+WGc7ZxDf2eLYUk5JBVw1zAGuRttD3gE39xMy9V7tlp
b9nJHQKe8YYmam8xdIA0JQhpn4vtdjrCgZzLX9K4Fz6k2u9PlIIWznXXsUCM8hox
zr/Ln+z8X0/AIa13Jn8LJ0MJURwNRMCpSUtIzCKkDsn1EWRFxWk+l/0/Z0SGnewK
EiSl1A9/eU56q64b45xgWNDASAuZF6xZCOa68tgfimxjyO3pJHlOf6EHxAlgJEeQ
/uXobeiSWbZvtHPagMYNsgTFLHOl0dE1FBTVeALoPYCeG7Q6FtqE1L9y5di7QAld
nnTWKLksd5kjvIx8Bbm5OaKmP0R8Yj0cTtgUwDTCB1OM2EeAG215hgqIxZhMqbm9
Z+IrDeVB6mC7kqNIKWmrZ7V4ydjGgdxSHHJIJcZLvubiyQvjl+HQFc+eM/JtJlnM
eDALSiT02CMBiCzut0jlo9WH9NMJC6hCgBHlgZOw7FVyNQ4begOTtZ648FML/4nR
CJuvKYeNShuD02YumkgMW8F5fZAwKGPR6HBYEbTfX2dh91v4Y5skKxvveMm7z2qS
pFJeV049X2JnP+fJ10tpP0xhTYa38gOHMqHcl3wgKVLpIrrU/OuLCYGhaaY+iOZE
3qAOBhMbpkl0OMmYnHmU6ROGkjt73DFv3rUkw9O5q0G84braX32dQZ6zsFz+vPji
H4dQRTjS/E+fqJigToDc1FbskkmVLUZ5BlO6QeY+OhBEgMGoGhtOFJYlNfYOp9hU
yFDjT47LCumsqN/0A1/5hrT6HfDEJWtqB2ED1arvwKXphcpp/NKOnJIBYJqH8aUG
J0zcZwmLNz5L4ar5LGG1rZ/Pl6C7OzbwXydJ01OLIYTgurrvfaPVn5UeAOaX6vh+
Rs9m41YhPNue+kQk8JB5pvW5aoFyYaCEo3dT5eDDDgq55y68KQYVYgD3tumFaUYv
qfKKntOzrxbtJdqJt+B2/qPnCf/wSqKrg/TAC/SzhVftEMdxtJbz0r6N55/naY3X
ouhjwTirz0thBwdf3ZFbgLzri5xyB44vZxdIc6L0WobqFpk7lDOxlbnfwEzimAkB
+v5ILsUO9DxOVXBHAKgSIbP6wk5TV4FnyOKY6fEUvRell4j3oar6kopGikY9kTUi
23Plj/ipi8p5CITDp/B1ORoiETBTrXXaMBFTE0UgibzY9X941eMtlq1ZptxOAZnG
R5W3ZFfWhiJ/20u459024tuboPEoZ+JlK05gw8EA+ZOiAIPj9F/BSb5BHG1/Btvf
Dyn56UdJ06t+qOsSBbDEkq66sBOvPoYD0mjQQ+90YNNAM/XJtyn/b/EN6qQi6RTu
zpdZ58LIvkaybB3fAA8sGxn405Y5oL2kAUo8yClnn9GUaWdusx0YLhc2CVvpGOzL
gfk6mN/wUUJ1twi5LKWGIy9dMgGzd4dat0ZvMjgywHfPmDx0vXcFtYREeV01w2Y0
7lVXbBLiKeAgrPpwdojhUWobSHp+ekjMhmDRO2exAdZMzLzRSe8xUP42xTyjbaVk
7kKpbfKMqw9EYAhy9tiMOgjhL/c0kD3ci/AryA+ay7FRnFLWfUzzyRSMP9P6lwF0
izGYMoqwJ48iUH90v0E+rU5uoZFdS9HHIfPndvBQK+qZVZiky7qoweCOKULVv5ut
4GTRus1ayUPl+/oJn4+dYZHZU/i1JaWZqZ4JH9VVEa6k3BCSxEhWPrKe2R2O4e6b
Iryvhuo2ZJDYCmRsBy9b7Moy3aq36yGmf9BTVoN3tQjTLnEJ555EiXGvki87Fcwm
qBgX0Kzs2zE7tX3KMtFUuZcVIroPJoaHkZAz0c/DewhjoEesq0iO+ZMHNbRWWKI4
UKwYq9Fr6IhklSTw/CTB6ZJgZnVyfVpgY427U+E5jFf+SeeFeyNGSwjp11taQ83U
uHWFQtHvWm4zqqX1n0NAxpc3/B3HuVP3aY6het/S2l59E1oQ8uIBsZndIN8Ht+tm
tjLSBNXiuUsWloPbr3hGZW+tdWly0gSIH4PB1qAUhqH1q8qTY+xjoCjplaUBqcJT
QLCBZ4Sxld8ch4Phz35/5lDd43kb2JKnZmh0hfbBxDsFIcGZ3nBpFyYrzq/tVr9t
OPYZtyL5LTe2Yd6ysykLFvu6bCuRHZer+6sMvhstKESt9RfNresVwGg2+5kG63f9
cej7/R8y0Gy+aY+AYs0YlMo9ZDXmo6xoNYAIKYraQX25PdvoFUxaxnW1DzSSQoDO
m1GnZMy0QAu/lsGsgT2szOoqh5Z/D4phPhHL8pWXk0758kco4bYCXiKfnSnGIQac
YwYw0l6zAZQzk7F3d2afyT+l2XubW+FowzoTQmnFk4v0fHN71b8Y6P0fXt8m0rtF
LsAB5dgx1FZDzIJO4O1jlrJQIl8516R4KDRep3AtJ8lZPnhEaAaKeno+BkKMWY1P
t4mb/DnaJR24hQBndSQm10p+oQlV+optWP1mUp0aQrOJ07R8SZE/lkvOlAtf75wL
X7F41uy17ILabe6+IAB09EKNvfdecKQrbYLQVCj7CQmQy4VUCQFQBi2tUMUaQfi1
dAQ1Vvb1/l07DAMjVdUYnfXNceXBnPhAzvjIdhE8fv460XvvJmXcVzciHMTDhJRE
fyjhw9X8zRcaaTKEKgy26MBjWa4oBrljOe0kR+OM1a05J4HAZ2BdbzzjCDxI4MjN
gS3YJ533DirwX/1zo4GDnaFNpRPNj/SAqJE0DhEEACUtRDvn7cyg81sk6KANvixR
NR4YzFcJSbtPhay5aXAgtihwsiNSEv0/m/wZQjsEA9VZaKUuyWmUQruerlYlCdID
LgJzJ4lrhPG1fzZWqve+Vi842eVxGYOp39EZBghIce5DenmbhSUgFMle7m7Cft1H
FH7jkZpwOjKuzFoF3z8hgsNMGEFLd/Lu/ssFNbllDwYhEKK8lUy54uMg50PSW0lD
qdLmGY5TKea/lKA4p94XIWnaD279kU22Cz4jg07i6ebRYNBXllummUNvA3/4Lk22
9HeuCOJrQps5kx9/R1f7DVYFu/l0gzTkR+0zjY232ZcsOs/ZX/QBLW1cpnGqOfNs
pyP9fnjfW5bROXEnwghTzs1rN1s+Auu8A0BkQ9i62Ccl+NnKW+rLi1wgOMcV3yl+
bOMTmH4igEupE5OsPcXqQJsWisGe+dIMt1rmx3mIEQFw3kAEjs2LX2INP/cRi5IG
E8PCwyVHZYu2vYW1tl9RVeV50dqxr/l2Y0sQWOdgwY60/9GXBlyZMACkPfbCFI2W
1mOggw1HVHRJmjqLH6+ErW0gk2vy6JaVVnnP5o+8auRoCVlCLvSGqdgCVq2iFjBS
/PgPr+axOUS5bFkxra8Y69bLy6wipUVHmfR4tL1VCn+l5ZpjccHqjUleS0R3C/94
4KWLwO/tF83/1T6aQLmCwmOlcY6TE8CCb6ouixNVTdEVXXEz/0w1YDJz8CmRWDcY
WgKDomGA7atr/1zNvLiMGGF7NeTTeWrZ21KnjXfMvILOIAs+FpacYet0vDe3SQpJ
6UB9VcPaE8UkmTVkKz/hJuTf/VGP9uRP6j3Hrrb7FLUgwwH0sgOkB1IjUNpt74xD
1uXQGeVjTnIXZ2IVuiPkgIJuyAqhBntiogPpHqiut09p7fysCvBYACgCHrUHIx8t
8CJX18izeWq9dPuNknodLMn1Hlu/Z3XVthJsnxzOdLTdMLheFla5CZQk4W/sblkA
l+eIKAG4op3zG0m+k8+p6zUbI1heLDdhbg8VAhRWFJTROL6+dyYWCS+n5jLz/iVs
3gfmBtIO7s22LnGAw56VaBTvNyjnRGYB6XBdebSY3rsfM/ixevgU25r3GtgdKNUR
fZJ7NwcEuw8ZvxtMSXDxDr0qNwa0ulNdMoJAVhhf5iGs6egvYctV3Midhi4Ig0h0
y728vsQEWUHUm3C5lP9VoRHvedn5bdxNzBHoMFnGP10DQw1yUKv8FKWVDsaSJUf6
g7wO1NAU0T2YGz6Se4/0RDkaSHMhkpJEK3WyDix5wYlcubQDcsUFZ7qVC+54TWwX
MvI7KPUZse9LapCfeKPmmM+FjiYjdFtLtBOAIfUbTPxCUTJqbdBnxD6ZEDf8Ltb9
/SyQ3LrlXy6AWMX8brGp4viD+pgF1FOFSiTnAPWLvSbfaezpy1YAjk02GYQl0P3V
MN8FqM2N8z25zrvurUvTzcDSSc64rIiY1AANW2rOjvM8gO4K2VjbP3EDzM14ooNj
WJLC/MVJEgFmd/FzyqBfPMx8rJgm/fZrZhw7OP5eHWsypas8MQ7u0mMCUr1tmXle
Bpi4toxYLVib6jdozN69lD5UFU0Qq1RUZUqsk4ZRG826YZinXjGItw0GLaChI6ti
/3kfwDWkg/xFim23rrSbwm+mUDD+RdEQn0cbw5kxLwsFUU9XTDN3L2WsQZtLGCl9
XIYLULv3SsadYs0wzc3KJtvarF07RbWCg4odBQmkzCEtR2fYon6BSg55EXZNGRxb
PEgOlGJ/lvhewTey0M+XX4/XOUDTqVe/6yIGfspXAxJeuC3ouDdB6Ul8L6cTdb5x
K/slNiQeTk+ldTjO1jp2Opja1QarvW5pL9WQ9XtZvfbFcee+c/dbyTNCBLjKERep
Zc/LEbquU5ys52gVmKJCuOZJvCqMCdpqRo6+OMA0FOemQEG9d/DAkJ64okqs8D8q
vXL63SqvKk7KZMU8WnspsW/J2PTkDOgl2ZceWTpglZ4v0vMua7KH48BkJ8/D6DGr
V7jDcke1isdReW69u/j7AFQhsIoGqdDE+u3LX/a1kcaDftl7AZEYmCupClO38WQT
/9BTXjFuIWyyy4CGWKagYC4aSPnTjIqXimvnn0HVrKz1uPZpRMuUTlq0epz4g/EI
+YXJHooOwlPdGROFD+um0mz6Cq1nlgkQt6GdPECTws/EnxtN/oaqo55ETal5O8Tb
Fu2eWagZrlIyOtlzu91/U2ydZZE/cBqjvWNYCPzWurbYInJs7aALBrmntenPMG9S
SC6XE75Y3FQ8DWBtERypj/a+HrkvUlhtpvDD1MVV2vQF3HYGmqBRzgvSnTuAMeL7
ANDKBwRLeGWXFOEyIBH6TnLjwDXNCE/EHbYV8PzyYT1TVCgAFELysyKcHzWqMuSB
cYZyn/xUcWYgsqfZEQOnrMmVojVrPBqhbzjBgeaqgBJfqeWiRePjcrKnDUBN18Fq
zoKaBbij87/lMALMPDI8/aclWSgW2Ufwl7cGGuvYV+1Rilau05lJG3esZf/od+Bx
VYyKqY6/iVfkHVVoOWfHdY7R49vubpNh+cnru+Z9VXv4EGOsjmfPlKKBmBBkWbzC
Qb2qVPBEHGRlvaKnjtm5T9CyACpTDzvQqSGkGzUbvPcNH0nYCo55O1J7ow4iHY5t
nbK1aVcHn4heyPfthF0xbGrR3+j7RJBcAd6jtC+BpfztSeyw6dudg3Khe8nu2N1O
J6VWecow0vwAKRdiu/fb/UKpGr//nNNUfznb4UH28NhKIxTrnWBED07v/RWlBetL
erCPWs2/opWDpyKuVNbwaKnteh6uaWP08fLn7Qedzh0s/jzyX/2XafTNXG6IuA+P
TvroElOOlNRACZpJ98OL2Atf1c11BWpx007e49SW+yGWiRx0umYPELb7rANXSc08
Lktw1TN00IZaTEzVo+21xNaMuvhu876RNGHiP4JigK93yZE+MA8KRFK5fc1Pl/p2
g+ypk5Ak8rICVciLol2pnw82U7qlsuemXjBAj0zoV0j3JcUQaxEfosQLBGgRh9eM
tzwyOe+LXg1a+LuxIF5kBxeLIsBeHXiCk/sB8grw9t7CpQFfCxO63ubj5vuBwGMK
4nMWE21PjnwG1jpVOH7Qs/XzZnmmYsEr5hVbqBsTrDcGwK3b8Na2fxHI1tTInqZp
ogVl4zTxJervLANkc0Rdqzu0eGrfKtqFhUMK7TAuNpqlRHRHpELOlESoUuz0xydW
vulvB8BLfZHFV+jddkryqULKEESxS2HDYOehDfI5xORZxGh25fylvOm8a14MQ9YO
g4963HvUjdl48Bu6NscamEUtzq2rDzHml3J/4LVJFJDAjcoKh4n5CrWsUSEtIvzJ
C4/di8UrPtU0WZ1Oagi9kmcYKmkfqMDYN2C76khXwnk9dbP7hDY7abwgYmq5kNX/
Q3Kw6toBa3GLBIpDWddpkosiEAL2ApIQZWkGt6BcZZ0n07PNeSBpQzEhDvdsHgGb
oh8/ie1yc0eR1xu6Mz7B66UQ1j6fsoNAqnLbMAcJVtFypv5NGbGmSs0g92hjF9wK
ztCZsUcUTfLDkDoLt6NkUUJ54QyTjVgmrw6wVmna69YzwfyXfz/wixBBVl5TrKHD
Jq5TeWk817jMfQaMeuM4UfpcydXJrLD9WeIyaTplgikwTqv7LfnMGvm84hSEK9mC
+Dm2GF9liIS/lNa6lwqqcMZY71vH/nzoEaIwyepw0yU46TzpFHY0x0zjOPVWzvE9
NFoG9wG4HHCNdY5srspeAOyMDudVBFQuXZrUiCVW1pqS3lEDBj6KC6ujlunFm55X
X0zEn5gokR8X/2b25rawbbm3eqT7T+L/kgg79917I+flEwYbxDhsyc7DgsSUlibf
pNc2sP7sd5DPA8FdI63PCcagbGxF9YfBsxmh8w/imhn8nSGKOJX061ianUEOSiJZ
U5AD9ofEQ7NJqa/VpBswgD3awX/mARrpgB39Q+380Ryc5afCKuxm7Sd88cqeM+O/
6fdexvGRx1naRfyjwpNV7/S1hdpRJ2Y1b6FLqQSvC+jYPfWchHbsIxvpC1/nDJjT
TCPx2AzDvEz6V4B0Sq6+KNQLC0cq4qmkwJWshud7GgsiRjpL/dBYFiG1aI27PeLn
48UowWIXeKPfNu0F6z2bQXo4THvULHj35H8YlG35WKB42iUyrEeQaSaehzMuMJ+1
Wo69pBHULaj9ahol8btuo4aoZMiC/vGRqkLAr8s8stUF6li86B2eSTKuQNUIUXer
Xrky9rXhdrazZakmNKLhZyqPEcNd3kGu0l6zu+o+AJ0ZPelovo0j1Os/2fIJabXY
OSpnoQT91BHPL5NKuv0AROQKWlEJD/6THztsBH9UlLQGzH5VRPr4/IPId4LuM7lQ
yW19bWoaA06JgP8fr71k6bMdgcy30N0/wf6vWUs91m2rTdqvlu9fIkxBPnIBoNg8
VGpZdNPLavhKOAdjPb28ThtuU+Bl6OD6CIb+kfsVXydL3yLZLZ16NnGmjobLSYem
Y7M0vwq6HYKtSTl5Y0I4L8jS2QA6WlSZ+GKB8D1kv5WfL4C1KOft/T+ryhT1W5wl
G4BmiHY1lv5LVCurBEi3kos7ciM9DxdWwSJpiFcFvZaR23gUor/GKOwxdmPoxwvz
fE81g4CP6Jqq8FZua0z49C1Jyf+RMaVAVfK5S0Ouu9q9wiINddudeiZSYy/kfktP
mjER+rzbdyNCiruBfBBxZdEZRpIJxA/oqHt6IeSZcsntbnbwPlYIV/TXBdlEpoWY
nxam5P98VjzTvY9UMUZ+aBKDs9/eRALB1PRMhCcdMPkfOcIN+yN8R2j8Q0M/5m2W
e9cKvXGmqz4ZjvvweDtxykAi6X8lUQEGXkUhYuQibzQV5iB0tmzOTL6Y0yObGYat
9cS9FIEN2cWWaBm8NYYFYE3Pl1AvFHinh+JV1DZ+TjxE2XkPgQDsIKaUk5HPy2jt
PnUzvAcuNp0g4/aaio/zNJu2uIeEbBr6XMVY8c4Yxxr7grxOlGjQBWHqXnoucQ4K
Bvs9AsM0BiKnpIrEjJRMOQ0hJR+Aczg2AoiYzdZYW4mdNZoy15aN9xx/gnD5YGmB
Cq8x3GJf4LV+iTJ719Yafw5vQX7A0i+tK3cowHvbo/WlR+8Wu34H+j7m38d0nd/c
SA3JKCFrkED2meYP1S7VEaa2bPjdmReomxEPvj5nap9U3v9iHnY2DTjFQm+hf+rc
/J/H0IvIeomyZwpjlXAdD/1lagEqAZ0fc5XLK3Meppc33vIJj0YtL5wfT+N1TXyS
k5xK7Lnqyl7ckvrzLxZY6LCsL3Dun7TWgoRW0H2EIpvV2cIF1yELNzF3Pc1O9wWF
cQM7TmuC26zWcrJPOzDV7G9xT+UZ3IhmKDLvgO8YQUz2904yi1I2cJLxyEOVbNB4
CoSotXbABcJz58DnYcnjzqkW++Kl/qrFgW8wPxAXIfy50giMgxk/TEaoeD9FwAbg
Wa+FOy6b2RZdRoeCd/zNR54N4mMBla6IxeR6YlMZDA7KyhjGO2nK30n/1E+Widsw
55Mt2eLkGMq2FXKMZGtHGx7nj6EXNO8CyqJ9GXNqSgkV/VshVD2RUL2iawcjQ5s1
jpo7InQOBTnwo+a7ti9yldPN+KgFC39RC6PJuqZBJRLUJS1cCX+ofyC3Gmdl5QGE
FTgTU7ouBv3e1FoB2X19c85yQg3pEdeMft1Jt37f2xH12oE3zng6/pIkjma9nPt7
Pv8Vw55zbEjLczQB2mBrwWTNGg/ROqzVqQrKWapWtZQZW7esnY3OMJJ5rxTuN9vs
mMLoClrfcIb+z3BDXKAn+XJ0zs4HqNPvESK0O+Iea9I7s8oUR/JOKvlQads/GrBZ
BIXefobUAREadvfdo1THngD6RSn6h2pD9hod3aRsABSH8p5usNAcgzkzGBYuUyM4
lak6EQwy7fHoKniS78rtVuVGYJxC9BTYEwz89NqNzn6dENJth4CahORCxeIJPUUy
t+zh/yqy+vnMe68j9hlMJ3T5hJQ2GcIAfiF1xc+HPgFnyifwhwYsJ05kLZgG8AKK
4//BFCnlHPEic1xotn3ZfQq5gZaaAzZ2zAoeDxXSfS5urgS/a9H41PROJc92QiC+
8NjE9rBddxK1KEwh7/qmQlSOq+/viU7Ca2alcivciFBE4oIxrrIZBLF80hGKBU7U
eG8OfZ9mKVR3LeeA5DwCFgAmopHVvL8tJ0eHVTVgvEjHlwvxyrBmMrpJNCuOds4o
LZH0zIjBpseBIaRG0ZgwCl9yhyZCMiyvP0UtG+tJmJjDa8at7ERSZc1bTC/SU+3W
8MNHdXRGT2E0bh+MrU1Xvm3WSe8sefrKQott2KzMFUVUefy0NsMMhKHW6JvDFOq4
Ykane5XSokyUj1idpkamo5wllJ2zqX/vNSjNY8vhFBIQ9IgzfKkEoMjwEy3AyBla
TqpNUIY88Pxb5s8glRw7oTdqmPTU6VK8NGlyeI+mbtaULbYF3dPdAXgB+XQhM/1+
MpnmduaGFXaEhJFB09jISXahgG3JffJYMctke2ZcVMrRvAzTZYLU4mzZWWMG1YqT
XJhk4PRb7Cv7vtWGbixjZ6P4EBSvhcPT872T7RvK857laD/7Q21nnd23p+aPZeZ+
P23wuGfvJy54fxxVLWqeY2SZu1kw7X+BBHBS/2NLZ9lXcIF3rmDt34EnSisCS5ii
1pcNXyLITShl0PNrY/QC8gr12LuvT34eOBbgF110sl2a5EOHv/PNDsMy3pTfIwUc
3VCF3ZCbBAK8Ns9Xvw7DRZTGArNidecTOYcNs70zBxq/FXu3JHvrqQ5zMXMQHleE
o1lg35N0KMn7jG1uQAoqMKspG013gaaek2e/nfXmPvsx4rxpgMCXNqKaYYP5c2Ua
Vg4Icv+o0iWlWa5FKknHI56QAz7Gh6nqnwpD9pq7dd3Wuq9mZgXfDSLF72OHdt8s
sFF4oEcq225jpwK0gEFdwHkCTUsCeisPi5Layyz+k0auqZj+apCITh1OQ4dRCqGS
76KCyTUbdp695jtFKqiTtrSRE1m6GdEaot1hoHj4fmVZ5z3ws2Xlg6RxSyj7lgJt
coNo/yW3sQj+Qg7rO8e4L5BuzAjyn8yzoAbSpmel6kKJkR9UzKXuVNmvpyBRFBO3
IMwWdMiaoywsC+qhFSiUtDvXE83FgVK7IiYtWdxjnjD1eOck45Y6sYxVT0SogM7m
x4XuLczWdYZ1mA+cZI2m4QacTU69VJhVkq/0oRy9Y4m6VDVL3kGxSIKpoxg5FTLc
B2cEJGYOMMU3appPtWt+GYc1GM8mzf8woqoi8TIlg5lgc4Xw0fpwWcl2Xgt6t/mu
knnPJcCleA0Smiju6ISaZjSJUG9bgqFsRleVOQMbatV6+rcTdpOwPDlBPI9DC3zN
PF/DBuhr6xMs8lQj4dlBEtHAdhv/fje0/lf64idTDvco87KuXIbn8jwVoLROGiyw
SLC9Ecyf8BGed/M7KJKncIEzQF5cf6r9XcXS0q30DpNv6Bn/KVf+Tjo7FO9aNjTp
S7hUlKXWL9pPqgAR+kwyiux4LgVDg8m0RRKBAfPHjVgkICKJUr8slUsr8iKf6nvo
Z+tRSqa1257HBrhkeiZHcUvFOzvf+fbIY175nx2HrejB4i709JV40DYvJmcVOp/k
TxGpNeFnOJzHx7JQ9GO33XCvlWQPKlDqXobro4u9zKxM/aOmk02fbSzLHhliprXq
kVbCXO0PKbjCdz5Y5jqZc07b2vJCp5KhR1xqpUWAGPXvv7Us21yZQre1FslIYDY0
4iekTm2AESqfXblK2XOYNm33Q8e2SuGM9sb5YavkJNntMxXQ6bi4rxsyR59OYlsG
IDGbtVqhGy1X2/D6AClGMYwPDm43wDenjyJxXIzinRfoTWLrxb5W0c4zuda5TLGx
L/Z7U9PpG7SKy6F/IbEZPTe59U1KjpSZGmRtaF3DsQjTyT6D00JzmnoPDtcvbVjE
7ePAhV8tCw6ifS5hSTQEyIhMQsONYLPYvWEkZa39WtkE9McaF9ljf52tt7JYV3qg
RI7wBAzFZz6VOj52Xpx98Kn1W7R3GNO4fOWDJaVoPezBo4M/Oeqimww7eNSd/sqw
onUxJfuhCI76vI6iDTANWVFER3K7DqhAFzWoBqPiYMDenmLCsBiBeAOk7gSFoa1P
UVNANbPc0n5AzyxhkkTqcBpHsryR0FGaW+yxpAV8d6xQfNQiDeWkW5wB3ZpGzPyl
x+LgrKGIqN66XSA0+UfddaxydpFPNBycD0TO6unApMx6AxzCHK5p60hsR100Dc8e
Jgs+BCbShEQ/ac1bfm1LQda7fixtgteBbu+RcKym8qaHYUyLk0llqN20qchp4hZ+
aYDLhDGJoExfVW4Z17vkuTQfKJIy72/DHQEeO/38r4m1xtLmuWhB6/cAtL4eXDaj
HT6+FlLS8e/UDr1X8+63xVjky+vU29N04glxdxF+6vWF7vkuw13EcyHoc6Zo6Gz6
JUeScINRE30vrwVN+8+DAV0hrWwy8AERwZy9ZMpGiBnx6fkQClOeHvN6AeTeUr7s
9KCCm/B7iTyVTZU8C2gCJFq/fyTPubHUO+qe3mKVgx5dqpPKU8z3EFHTaGIMXodS
HP/o/taSFBxWoNJmfXvDGjwxc/YaeM9MJs8VmVIwn25R451/zNDZHLO1dhCgqQtK
mtoSeIqJARJDNUn2p8T9+pVbP1nDVU5LE5mpUb76FGJL2hve4OUORHhWzN+Nqy+r
RYDqi7/nlDLsDs2m7NwGezQjau1o61mFDu6YGAcFahQRUSWO0yTYzwvDKAfUKip0
T41IDoCKbjCF+5FdUwWA0qSh8Sj74WKY9GoAP/EpiWE8PwTme1BxoW8gM8AF57/F
XMY3d7NJvDOHwdOwUOIcGHtzqrwIyyCj8itsgDHXEe0tOEH4YC6RnEt951/yN3qQ
WCFOwf4bsWaA8HTdXyysn2kdoqclME9qSw7Q5EenbwfooPY/VN07FNidDDv8FQgc
9tZyu2dO7cXYx6zc9tLvOHqxAtYlrCtzfR4AaijkpDkstJ/9nViAt316/Uv2SQwK
bOUwcZzYoQU1RrlD57LWyGQT8VwBc+tOB/Mu8LZo78OhA7ifz8AztHGLJy8FBehD
yX6x11uoyQE3oFHYSMSbJIQe7VfBwBnZRjm+vQT4Wkx1YhYjloIhVxZMpYswfEBr
Nh7JhztpOVces3CHqgwU4x9HtZ0v3UrnyAAPZLG6Nhe/r0WPv3CB6uPUzjBaIqQn
gDBIArFZeursFj7XzRaPp0nnsL1cjNgTNCoOGxdzOXh3ko0zNWEK8kp9Io1Iog8L
QSrquJcrarR5XA6uqfxxQVTdw5OZSfbVoQC2jiwTAemVzIl303pogAcYAIlmhO+3
kw9/h+gWCyteZhxJBhPHLQcyiJebIl27movj54uUOLOTkfrKNuo1cgFbXYjecxLG
2A12PZBChDWAVefkdj6ot/ZyN1kTH7QkavD4ANiyqdGbQouJIJY7tgWvWA1i9DBZ
h5hzQZQMpvTpymAlqK8gm6M4IUpIwzDB3wbJuVxXLJcX4USlj1kuqcYJbhMzAkj+
o/ktQMAY5A3PAFBAd8wQczUmx8foU2n00khVNFKGke/dHH5O+lyzzFM2nrZm/5ix
TimA+sgu0+t/v081vJ63zPxg4cSxzHoaKXa6DtnQduSK6VkovdtsmX4tppT2ma6d
w/4MPUBTlihzoNFr20RmrA/KQDvCieVR2juKak20A8hnDvmMpewBk6cRBzeG97/4
VGzbpbYcS2Ju2mZz9TxyKhD/dknDTTUO8bREO8M3U3+iKDosa+vIr1XANg+vuThp
W+CjwCdu6FTJDvmSuael8+jUNEVMkvLbL9CwySSc6MtHW4BiHCzdWOiYoeyx64JN
4agc3ARZZo+vGSui9i75LQ6V05lAZArroacTqS6k8cvzfo/7OvSy7eG36Iy5APyU
SvTpOrD/unDkQewE1Atkbh6UiJQik/2WEnnEV/a72amKA50Xtct44nvuOB7JbtGs
z8XLqMkGaDfOJ8xmpFtQAIufGBu+YPy0w5j16Qdm5AfNbGKCSGML1426BDk6/wrv
43sJ/Mqi6XQ2kRNAp5E+QSMCbsu/XXqPB/x0ulqjPfYgJ8GYWLvFEpY1NhE+mCN6
DlMDXO0WIhdj3urTWX7TwFZPuE2ijq8DQucmvwdCsyWZX3pHldhimLv4ohVwUysg
84YYocfZyknObM1Djh7pxdBOfIz42jnAQjTb2+FyqLn8Ou91WsMPlbtmO03V8IS7
tSINNtPv59eJFak8q8sV+OzaTc6D2aGlFW7U2+kMtG6kW05DtjjMWVcBeGwPDyOw
cGiFazErc90QOK/89/U5HUWWwTdQaE7FzVPSv4W30HB2ha/kvrXgLhjEeiYkr9Jy
GfpzjzX8bPHzD46a7l5NFBzE6O2bzrhfO+ozFdcQzupAwt9vgYTCXUAJuhnKLzqu
A/ymfg9Ilrmq2ZR8gMBMtT5ytXj4K6EdjAjoKdI51Ch7io3DtM1adFpdlBdqXpVj
Ff9PVNud+inwqqviC1sc8AeimM8zR6Vax0DI7iQTmVLIHpmnR/uT+a3a07wIGW0j
NFrFqujKJwSXLZjZLN+joKkb2Cy6WCJ8gY4q9mjIbHMDiquDRk0H0xq5KpDoX2JS
kftbXfczJBUCwZJ8qkrv9MMvaZYgLwJfdZbkBfA4lglsHIngZLOyQD658VnnpDIC
2BJIrPeYlPNZl+1G1j6L9rvpHcimP/3lAD4eAmYdcsj8m/a0mmk9CA4Obog88kan
MGWQ7yAUZz0HdVo2B535EjyBrJ7l1hpiEVkBp8Ye2m8JNyjflIdasIPzIwQbLjK/
n/l3x710JEs6bJQ7TJ1ZkfGBeZ4VuuxpguPo9XDAaxFqWZR9FnatI5vRgve8/1dh
7W9LhDW85H77osg3ta3QPXQDoMdYoX8WY9j7upIKdMo/0FXBwoPeJJHQYyWF9Tlb
Xws5xQkSK0hvIVWWXEYtNVKg/7uj7rw+nGDX27VPLmy4BG8IJbsGxXYTuMXHPdnC
qieB9ayAgL6QcvwfXZ2zx8Xlvyuk78kwHCS/xcGUMRq45/jiWm8Cxt0B2eBZ4AhJ
RQTDpSIEv16owPW9w4jYKqChmQSd9egcqf8xkdfhpYyg3giBNHdMX0U3LIF5Asny
5G62iPRzmMwQeLcbGjor6acMrkjZ0CrOO/62cDg1ln9B6en6vyQumrZTGzV2OJ3S
B+Smlpmuc33XoTd3Brge1c0z7a9rNgWJAes90R2o9sLLi66nNOKeuf9SaGKPNHCm
NihTT4qiftRMoem+xzd8TyYR6mbbzHE7hBmYFqn7S+FYmwOqvSIUICfSLlEtC2cc
1QdGvN5YaOHapkL4hYXI1wwAJrXLiKkyPNF7GR/bUNr3WJGenOrqzsluIaL07v9r
21FOlq/zTPnNy7xOg6BInvNxMHvEJ/FTWUne5DcAiqbDj/cnpXee64JgiFVNZ0TX
vk0v5NqI7/MMCZdZEAyJ249Mc+eJxtDIyW5NMgFtVayuQFTslmBi6z05Re04ZXld
m2iEI4T0p4TM2xkAFgaQ5NweZtRzT5bByGH9gnbLRCcfs5gVqljVb3v+Zzbh7zhm
+ITrmOwiz5nfCL44lXQmBOxehQwYZSqpuqd0T0rObg6sX2I2MdN7A8f34EQe1R+q
8zXeyk+3B3b263ycNlvWONHC07jXw8jUuy3REcyJMsjonv0F6Qeklg7OMJ0HVU4z
L3tTguj87KrIBbUoo2QOalPtGv9qTw4dpfGdMSN1HlJTcw9JhM9sfpppuyERthK/
Y5RdwEmTP3qNtp5EFHGBdQH/W0fUJ9NaSL3iYc6FT4xTVc3YL1IDNKfSGxD39t1+
Xl6FM7VCeTYXEZSk4QI6Z8pyfO81cInKTmXxk8yWymwAY3CjJhZ7C/91oyn0HVHO
p+hPf89xcMZSFfFbu4iyOHuodNgHLiEvhQ8yV5//ymYJFeSF/KgOedvijWt58AH+
qX0TqxZixXUAATAw7olhXWcSo1tqlkFowFdaFiAvpChmVRd/1f+yOS+I5yoSjbox
VE5tCnJ746Z3565ZDDpd2YWIgtMc6lEWzV8y/hHmM/sVgbAEg0X6W7n2v2L6b/LX
jjDSpQiT/NWo3oOiTx0Z3GWlUyDM+xqGEr4A1+GR+hRoQ7YouOsATIhBuYw8ZVOG
Ly88RxM9/V7UWCmDgOdujhEqpopP1MHYVzL0nS5jeXG2qk7vJr+sx6e4dTChcwq2
hC+difL53GsQ6cvlLws1x8386b1/4pu65WxYz+2Fr7QXDDzGt+bfnVzGxYU1HB1v
wKSLz5/ennEB+1jqfU9/WHq5AIf/EUv02AAPzoAgJiJIlJx6ZVEF+MrTnxkKAc31
L5u3otHIJfOOjDa8TMfkGcevCUGRKKFkAbxO5mn91I2ZoPVaIKoHNNIRnq1mi3eC
thKs6elNC5k7Kl4aD14wqxttHo8/dXaP++qNn1prAesilfXXChCh6GlNfPofqAxd
jGFMeBk6kApx4E8hDPmYwCA8Sa9RPaRkd/rfhyWGq3dlWssBqdSyq0DRReGr8r1z
eD/CgYyhzUoxrtxZVdEdZvY0vCXpW+Uma/NMOLYZAC9CmhV8W9sXpb6qX9GDWbHN
oKTnnvjmJzqzJ0yeLKa/YSwCMuAG2hK4e93Pzg4yvZ3cmbRg72DbQIB0DJmb4Woe
+yUVHWATGtywIWVmIHzlJGUBCx8v6HLKgS0uqaIsv6BZOfIWprtPS5HtyR5E4Dkv
eYUEKtxH+6ozoHICmr5t7uXAJTZ8jHTcrHDg0wTbB7ZY4Gn75TqQVPXWEu4+JlG5
UP7PUuoZVOrHrNxosyhoue90gXBARHT6PLaTI6xgrddL1+WortXSMYlUX5ofT9fz
p9J7MgK2YhwspfJo736H0bLUJ4jAX7WhNkQsQqR6a0vPhAt8gqa0TQN/e5PLEoMS
+YplUj51jjKT2KU8kyL4O/7jncWo0+JdPvi90eick0QwKFuk1UTCR+wivVFbL+37
k2d7tbJUYPFqpK2HGISPCXih4/lM/jacUJ08b60D1v2zQnDNo8Eu5PoMeFXQylmK
I3B4GVG3pW0hLMd5BM/dI7qEu7vk1u3LE5s2xYCDkXUP120+IN1700RcK8wxjpiR
nNHclUl+es/xjiwFMPsym5vtX7LGPQ3lmyLAK9vO4jKF72vlCtb+usT/Q2/+Gqa1
Q9ZqhE+UPNYnyLzfcBjtILNeTOoj5X6zopo9dAxAPCRayKM5xQy/vAEjUGPK6ArU
TqPJpTIMIyS6ojuSevdsQ0zasl6fjU45bAR/w0aMo8IULQjv97dhDYqXdrhjfWfF
/ES2dfn6lS2gy02S5yk5itxPilhzA+f2uagjY9eGmlml1JLu2pwcZm2nX3VCk5nj
GE/SqzCQVJQk+RqXh9GtokY1FL+ciyaqMqTis/hNZz3AlZJA3UUmqvv28blWutyJ
5cW8OE0y17fJD5vLRGdF+dwhbJ9x/zo2q3sJCCcbecdR0ajO3VB+jPeoeaZ3xnbq
gdcmxEsh/VzH58UGwxqIhDcUxVNDl4zbFhcQ5mhHFdHh3RZgmTkComL04x/ofJJu
WU4zp7all1bDp6Wp8c3JwGhqfFiPg8Np7k+4Flp8iwWVvZ8BlJd+6ZuiYWr++EDT
IXqIMD9SKAOYAE3cpihc3dB2WOaEGeb1BQVkaO6DbmKomGolj6kH0F7jPAGphwKK
WAdzCxP771qYGZS48K0RWDf8CBxZuwgidhBjPG0Mup+zfQgNOzGJj8nOLEsya9Wn
XAwIQ0p06iIMxJhxSQ8BYXLIuCpjFmyheyrO8cuRc2tDdmgIOlI9rq8w91IlYYwB
kZ/PAPXbvYCkWQ37c6ofWS+KxzzbOvtn9rhe9biFU7LZh7B10z0xHlUhNLISNxvB
rhyVCIsTJV2WhJOHj23Q09zCPPUkKngeLtL7SaXMTIg/fH18mFykw0IRafdHgyv5
xYIgm/1SjeHzaD/MTEpBiW2o0edFo7E/Wc/irgSU3zRWcyYiOfB4yQDc3fXAyQzt
Vrtt4LDmfyzzzIZTNAl7jk6lHRXsEuaIcgHL8adNzUmhjm3s7TfydXen2+SYw/xD
lkxYkwOrCwKdMo2D3DnCn61nzlNHOrD4vRZmhsI2nqcrgG2XCJJrl6tbclaiZj+6
cASuWRkXj89fVveF/iaYLkeTtzof5h7TPOwLsEk08lju3cboJTFFtwvQxTmRtlCt
gy/HmoQfxGB9sDJ49iBUtQm4WEP1D48y/c1Fso7OcIF3oymtvkZXBBwFvTx1S6KS
o7bKucj4YJQWBK4QTlFVPj9YRjrbfuqPt1jAhZ6QJSwAIHpM6frxGqlFGu1reHwT
bg8LCrmR+yCNZdmlhOV/s05VfyFN0I+iOLpwGBwbyl2Q1tElsLZtSEyhIc3gVcv3
oNpD9KFsiLwzNNWTX/BDcddCIJrhXAngMn1lgdOhcFyutDewa8CiSvirLYUIzSSK
ppBj5VExZLJPUM1+wiHW+jjHQut6Mx5gvIy4Q0vIDpJw8CpnYI2Y8Yw/a0zg2JPw
DJwwNbQCPXBTWDEKsaa5wS5nUU4JUh6joS4IBFsjRa4yxby7s9Y3C6s7vzLG8X2/
MjxipP6oJ41pk1MpNwiDnzspGRM7Pkw1lZgNF7qC7P0NU1m4G0YX44C/XRSMrBIa
sRMuv2STjtYA1Dex0E6f4cZA1wY/aQBdMJn151Hadaq6vyhcjAwx9vTpEpMQUZoP
syx4JySqVMlfnADI3wQi6h5wYroc+NMbvxlECioOwtv+terTEwrlSftnSCqC9P0U
rNy7t4+6W0a8a0XgkVwwXLrwFovPtIaKnpAN8FOE+DW7T9QM0wnv2ARCXnK7W4br
qJS81g1ulCRlieFlsBI9ReYvrEGFVnh/t7dmln59ATDeB5wXPxYdm+pOFTLahUrC
j5Rr2z5uppJ0QUmrFHjR1jJIH8J2HDJdjRAaeLVhcPcggc0/x4NknlpVBQklJLyq
8gOY0ydZ7c0FF7rQClneg8mIpNmfKRMt5VvPX57n0+rjCjhG+YUVCzH9Hs1rq0JR
K35Bsh9+uw+skamrvZXY7KmEbvQhDS/ts/MOznSHtcEqw8d/NEhngb6xtKldOqVF
Z1L5CpgCzSvcG8MIHOW7wVx/SzEKItMAS3d/hQ8srZc9p983wcNu2Zt7VsO1K/aZ
GLugGjbX0hwNtD+E1gpqRE1fPpWg+zx0Xx2DuQCPpulU31NYmXm/QohSYEnp7W/y
oPcI5l9UA7OEkul9vogOBuukeTLLzKnDXumH3pcKooGlKxIpkSRpoxqgYtR+soLS
xc1FrUilSulk4samJjiGdT5GeLkok/CVv387H8cOoUWzi/l6qAPz982AAkU7B0Nr
2yR15UuvppUSJ44SayB/WQ32jCX4+NOanBtuXNpZbBuBf4ulBCz0P+Hw5vrMu+5F
ADWomhWCuAEmQlZ0ZAeup7qw93NZ6cALDokteTyvF/aFAFVGjzdp5qQer2pS6Zqx
2QLaiVEkQgd1mFC8xXaOTD8oja/ZGCpp7mTLjl8uwv1RapT5kdGaECcei7xxcz78
aDeYn63dXGTdfpcM9w7CNFTQ9StSFjqf86nYGFu5ZhKhjkJRZLQgCDb0DW7xZihv
U9SWFvbEb5Jbse2gQESPSbKUa6mlNRpuFyyvUlVJnXNEG+YQykjq6Iu9+fr6mkyc
Yo8mvIC0e2y0UEs1Zqkvx9QrvtuG2Ylcbl48hEOMiSpMmRXcWyMwNHmT18MqOWMR
Y2+6l+NB/MA5TxSd0p7PQ14iFWyAqzzTZKOX4Yl57kfIZ3Ii81da9QU0f9FEbzp6
Qjv1OX8v01uY1oAz5vaxbMnrNw6E26iLQtffDGeNwR48jOmdyKIKc5qC8w+Awa1g
sgIHteTDh8qdEPOgrEsQ62c2GldA4Xj5N9CV7yHUnulFam4OsLyrHRFpgPd+8Wft
nqPDM2Ke0hC1lyhGj94VHQFy3bQQk8/Rd56GFp0qevto+JFOGCG2F5KFY0wMqXjF
HWMU1tX3Z6IiHMTo7fI4akY0pkj1njDW1nBBvVPF6LmhYb0HZz7nOObsUliwWYH5
Vi+jAdAJh3V20BF3DfPTPkusX2cZiUcQ71B2pGgiuTVr/jFMeHg7EYWANffQbOrx
IQdhdsRKHGDcPjTwAC2wNioniDtsIUnX78x7W/vmjDho/yC9vewclPj8N0SYjGUC
hwvCpbwlLExJOd3DGk+AJ1zxYC9zc4hN8O9cXBbQkUCGuj7BaXwJRLYRqZzMCiCj
UAotxlm0R8APD8YSmStbNrf2A8oHnH/uPBzXR4ieloi05FmSBOqJuym8r66GgipL
xDVkWBf4JVu+zMT3Cocp+iU2cHZj3B4TdD2Arvw1J79Erz0U9W2PDiwErZxgNDqM
aWNnhlVlJ6uBBuDqfG7ydDxMdujEgD4xyvaIuhbZgi3AhRZmfQgZ3RjEotVYCh8v
vZYhKYy03Kjkkihaw+QJJIuwSihTB4aJ39d0w87MSrLnTbUvV+/bBN6OJIaWIiFs
vUPvi2Uipnn9/qTRZgq726Sw99qqNrIV4jxcERD0sjZrga44RbAArsB3YoVVxSP7
fSRyLdl8GW9aGBIzPrdNOXOmcct8JwvkrXvFzqibfoLpFuMWU/PiUbdQRwGTE4wI
MMYhPEtrKkGnBN/RsEjZ1ejTvgV4DZGbqQW0ITPx4wBZBQXWA3bvzKhOYCd1KtWN
kqevfg4lBKXEGFvtx+lREXQUjNIrHZdnwamTPk7d8hKPRyPVx3XicdV2h4Z9HI0X
GMSceSzH8ZX4+bxilAQjzIKAbGrtlTQoaGI02ejkleVebs8/8ozX9qPWo+2g6MHJ
77ZkxnrVMXVfwo1jiOYWLW1pPjIHOfaIweEjzWRpQVe7g7+3Rf1d4n3012quRAQe
rfX84bizPdw9+8osNA2PX3x4IxpwggerV+dLdFzZEDZLFOKGopU5W/xdytpEf9N8
yc7SH/gwzsCI+Y/BnFDlCdeXjt4raFmYdI3uONL4TENT8f4/+z/RfCquwEIcZIeZ
3ZBKEoKYTW+XQjfr1NErYwY5cv3qvJQl7w3uy13n0dwJq/5RzjIf519Jay02FNIK
1sRYjP8EcjIeTOto2Q5laKmuj/PgjlMOnVODRGvNxSoZtZLchal6I3oWOybAeMNp
f8Syx5FWFw8BcBUPG85Y20Tgc/LxSQLszgL/Ml6bzuB459TWfSB7w5A9nvk5uflY
yJ2ZCMn9z0o1pVUdYWBkSTXNY1nIPRfKDpnIqlpk4ZeYafUjpIBeMpOZ0tSP5FWI
A4g90datjTP5rZeRCXu+1Nqcn7iNNO8NSKO6KUWZvo5h8i3wN3gyzj50bx/5aOmc
zgi4lbouO97LQqH6OhxYFpW8ROzdqv99acSnT+3kH+6M9WMH7wvaIMJakr/MKw5X
uTB1uGYmHI6myRYViEe384zPfjU0S4v1XN8XP741YiB98FqubCzOTbPjVvc694Gv
jMUO9966HYq/zBrSD99u0F0X1j8Dg/B8Tb3KiMOof+cMPwsOl8zhn9JO6Dr2eS2n
wl7LU1j/OyPitPaWKGLwMAx0lXlH8bER90vIbGmgqOSzUSpHTW+ZCnoKLJcXxIAF
4LLEFbbsvehRCQZKeA9fq6typNJb4vWUmMHeP3tlrlG6iLdOSI4gwCbRhTMhZ6Nj
h6cVa7cvD83madLo8dtoRzxDiSSb6GssjhJIX8tt5RZLOt9B7jF/hay6Qdd1r0tX
4kSy0pqekNIY8t0Awt59wijHdb3rCuSXYbqMh9cCogUZklL7BTQJC+rKPoi9SNcz
QUc+U/XPBrjIDDDCG72KVqZHPU9JTvR0675/YT2sYimyccjfrUl+8BJMIvDIH/6u
/zaGoJLwrYMleiDMIeI5uLdZ485Ninn2uul8qjXApeR2bWzM5U/vG5v9t3q4uRgP
1KqmQ1oXqMPw7kU/R8sBjzM8h3Q9e+0XwAuBSIkrXZBqfl6KkrOdNmJ+a+VB28Ja
R0lf5fcKLZ1nPCyvY66BP4KfA6+r83bX7LOM9R2x3+YYwPN57KCox2eDupldnqwU
fi9AVgxaiMgLRsrAqDB/vROlqWIrUMCy0+JFbTqZGKfNUG3AW3J9NlJfBRpQYv/D
XV2dJqk2zX+gik0oXqbVtAJQZbXHq0lnewX3saFkvnpbsSvXVRo8eABG4fbbmskK
J0goCsqakmmOhN2/lQQO5EBLdbtJ5XXT74E/p7AWSveuhZwkAU+qCKVAEHIA+hC+
UO5WtfEgDowSH7QH3xu4eJWceWFY3IM4H7lR0Oirw9N6YJCrZWyoOQFeagH1Idgx
FOM+DYt6G69W/lNu/4gV3c/j8kN4YG8VCG3SPtFRxwSOIbsjmpWyl913D/GUiHoX
c/EsOKufhNe3EzNWxHgCD+TBYIttJMSQR2SyusEkvUPdg3MrLiW0dkk/BNrVrFQv
YQ8GzmH2vTdTcYY2n947uR5QO/1vbWCmAtoKeC2a/+xdlx4yafQhmii96Jv4/+4G
WF9h2rcbDPfPg6FaMRz86qDWNMtxl9186bYHkcLVXSw6B3SNQHYcfkvzMINPB+C8
DdNY2rMI3iOMKjmlx2R2Wis8+9g+/26Sf8gqa6mS7Ws3Mkt2RUaEW3g7XV/ZA3P2
xw/cL/7+omQ2saje9hm0ijiM5HcaCibpQASL9qBsZcnbf/5iUf11qUFOM+Wv3yQ2
QM4lCsWFpH7UFdfztFtor+IIs2BkLXnmw0ExUi5wjvpgqW//osfnKCKSj9TYJOWF
p7nRmgYH7pgZux0tgdLXIdRyStyokov/HewoKn0NNRzMkFwkS+wuoXnRqjwwcI0j
nfVhGcMTg8M7FwLApk7uHYuFRlGrfsKtt5boHjEDTV9jpnnzWxNcLa84h6GkwG9x
mj78S9QV/KQy/vzs7qgS+w70I8VDcjND0CnvOXwp5fgeIHaIk6m+CSQwskyBdi3u
yhgFJC9Aw3R2Ujy0obrDzkIEQDUw6d4VljLbVxrUFa6bgOyIW8deftznZ7dd3qYl
kiKB317LwFt6Bg95zoT6c6LLoGGEjCVM9K4sstrMBhKcg5lrAU6Gu08ZG3I7E42s
et9Xf+BlFH2p0NyIupupE9opXhkhByXYo39WVea1reGtEvf5H5yI+FyKAPxiJsPg
oQVYxDU3hvKYogD/Odxh3QH/FYc00lzu2Ra9n119wOsoUNnbfcUjCE2PYnz00Gkm
NSssBIXNHddGKPn1hrujjtqCL38CNkhNjV3rHWZcPoiXmRXHr/6k10d4dABjSD8i
BUYQcSgUIAokYqpng+HpXvnX3PDgtVqOZeEK6xNUMqldPGsZXcrBnWVyqf4ShzbE
NPQLeXZWDJQtqxo8FQ+Vc0uH+7NnF3BOspZlWvvt1zqsrjfGcDkB2NfGG5TRo5E3
MYkZpv2nZS8No9SpgFoJO89b0ATEQzkunT/c/ICrz54EHx5PJ3BJVSeLvG/FSNMi
I9RRboufd08IFdGq+U8waUY5SIANqj7rGx3HbzFlOAwTCfSPNkbEMB+SNjnzL6TR
A2OmhftubYi1uvOiVf8FC1JEMpDIWTAIhk42d5TTfOlP0XS3oPc/BzswMQrdwsys
yXxalsfMeuI9mvK5xkpPIc6cM2F3BZpzoTVXAzTKFHmpUKgzgF5dJmzVULkuJQCC
yFQnLwVQCCVskienlSRa7GsoPTdDfTJqEMK9sqHFdvMTxHSFnYGRxQfiqXOLs6vH
o2cEE/xPumGAxnFSC+DkznMOgtgCf079yrWj+i7f4lSoN0bnghSRxnI+C430gPo/
gjWeeaX8PkjIedutH9cblXorOkrIqTmcWx2rWM4f+rvHhpTbFL42jb2BJOdLTWY1
M0rSr9k2FTOh5tXRFFxGigiVOLoJgs21w9vBjGI+63JSDejNH3+oGHyzG8RFWj+3
S1/VYX8s+5xNWJ+mBFHbqXTC9XyvzXaAJDVjFRE3AtW2M6b5CMDt6v2tV+8WQWfG
M7fKoYPdZZl9Rx2DIdxClwLrCbnhk7X5ab9eDP7wqAlBF3LoQwynvQAEvwGHXTBx
hbReKcmT004b5lIqI3klGL8SiKqMfIfAnRDJCcTCo/UpQFomfbgVLblBoh5qqrKd
UAoiAKyJl50OMNgFRipZuyEVscQI2KGnHYg/4b6cxZHUibNosj0596GtwJLcNCP9
uAxycp9AIOi73AdxeSBafPYFHFeexpWVNQ6i/o4t4n/+gl+kEN5K7O3mvHOjp577
Z1fbKqQ+q8S/JzIfHJqibzSSsQwx1l96HD4CybSpsHNYZaX0Gqm/kckBCx4Hjff8
ZyBPAh/wJ4ZFHfMUA3PoNvvLtShSzZmNPkvQqwqcc5tznfvXc1HAEmKmtl2t6ZZP
Sgj0UTqmR8feoNKKmk9yKuI1Iqevvt9aOtbIlOR/80X0NUC7zsGuJTrXDQom81qH
e1DPfnvyqVL+MAmJrqjHh/BxDAANX/dTL0UmX0GPMvMvnNCo9YA5wCOAuWVQmFKD
95DQxfupX/xO0s7H6rpf6t+rwvsjjxTsBcaYb5gBC6H8N6nBYR9pX6a6CMtPHlgS
TI2CJtF7p3Jz8b4+vqUKWGXFyvJn3/mYEDATobAXRm0ZH8xeKkK0nTaCU18u45DT
YSoCU9GM9PrWnZBlkfWoWiEbhu7rRuN6q520cPmuGfgBkG3nyljtFppYKqfsn+67
2q/mxWH0ceno0rbt6jk5uUiEr6HpEXoKGJcE4cd0j5xRfDWVXRti150dyoFLb2Tj
LL/0DSyDeKfS1CXM2DtKZKfSk9Og7K+bBlWYjzkciuPgt8HSh30mcyeMacbBhqpb
rqwRMVruKGcbbv9f54d7Dh0orHizyhuA/HStZlCfLPZG3x578Gw8sbN7lXwQooyx
P6alHnfLEsIswXNL52JfTqF490V8EoTZ3FKfPd481dBRzYqBEpjSLgV9DPHI2mm/
/4R6rbdEbOsqG4lV/KSsqnp3XEWpd/MwnJ3IBAY5Gt2Jxdh1JEgAYK8xnxJ4+JCC
hZUWXUvCvZZWBwVQ30+uA/h7D7QwkElRo3P9oESX0ngSBluc7ExkYVAycxg+Xmcq
zcVHZW7ZaObJr49ION6s36jnxdDdSfT/w5lcLbHojSZgfKu93Ym6XXg2X8MdD1JY
jt0YA2ss3+fWFljYQ/55OPrKWZNFSo1vj1cBz/4VTdkKmxL/nOmQWiP+pMUQJsSJ
F3seMn7kSl3MVTHZ26p6QWYsYQI/XjhRqBj2vXokgAykNav4IIvxk2iMLCiHHvRo
WaqhGxEfK9ZDe0MglhGGeh/bKTbOzjwF8cVDUNniyyYnaPIV3eHXRzQC+JQe2sI1
1MlNDc3lg6J+UaNwWbcnjMmBCJBNMwrqqKx63adL0g3ROT+1lIXap5n2QjyudfUj
pjYcCh8FgJ1arSLsKY2h9wHr6nGYZ7RbFrwVYx3zjCG2rZJI9liX1C4XKIteudyl
dX+LZtr4vPBiutpT45S2GLc9m9/l2N1wv2nKNLCcYpYXs5CgXGttz7mZNot2Iapx
e+I/s5un94nsbAW8wCCN50x5i+PClLPwIm3YP5M1HpinDmWYCMmGCI4XMF1HMx7m
JnllfbztT4kj1+rG2E3t+UZXvoyskdMgue7vzNW8Oa/GWw/ijxJBU9MhQz1QKFsG
zYkq8Gcvtx4PeX+BXpFBRr51MbeLdWDp8a4yIO60NeasQ6lrz5L1btQOBGie61bD
e8q6dQ7guNpyD7YounJkSUhKL9sRbr5Tj9Y1oFpA8ZM12aFP2Bgpbd99/71nCyA2
34Dc1OdRbbljUJM971aSu/h/JnRie3uSiPHSp+6bb6BZdv+242sE7EJdEI1v/ZoT
NDyfAN8mEA6Uvaro6ROqSgOhGQeTFflLDqzr9ZT/KUPykMJWstPPUKlWvB5GxrJ5
ib/NzTepGF4/fLsbcKFpQ9iEnYZsB/HOQ5wcsscA58GRmjscXCxU9+HZcDi9Dd2X
WXYZeqMmyFzgMwmS8ijVHl7tNIREzCMWx5eluO8IDo7q1EgEXS4jnfUVcTDK9iTI
HyTM9yloPRrdiADyH9Dpu/RoDLeZjTKp+Aj83xIaB7LkQTuon3hrYrOKKItlOlH+
bJoh2h02nmHGZ4viQo1+5VfndbTfGYzEcDgxgjQdEG8RXzdWjZY7agnRMKCvCvSQ
RHsbklq864p6UUL17/uQcZUVgLhnIHIxHtImJ06jxI45cse6uyYQqYt3NTyg4mjC
jhlXET2OWCeX53g74+iIVPFsnfibyG96ZDzSMiKkytOZBFrDdCydRbN+Wd2EAF6a
4lIL4pz3rEOBsO0pGFqOlmkUrOfd9xo+CvLC9ZnxJbFO0X14apP6NcgGliVyC9MJ
baUMrRVGFf3cRVk2AvQKshysQsIEooiJrrLmqn5bJvEgPnrtIA8uvSeJAjgGcjFK
TQjSKn168h8OUp9YnJuFPOCog1W5hZE4gY/oWxevs0yW7TN6obRazpCMiFYSb6sU
mwyo4mjeV62uybEGViDEABvd2156B1U4/mwzp0SM3eomrn0PqzISzhTyDMkc4i92
VVSgj5GrERT1FgCs2yglakyZV0CRdlyqW2w25h5E7C+X38v4mt/0QbcJOO3nL/LK
9W02NBLh9o4Jr11yDIY3JoSyT/eURdhfWG2CrLzUwiw7uBiIJiwJ3lvdNWdpobD5
p2ZWIOgoaUeifrzkVPuAY7f+hdD/KOlhjVHOjyF45K2TgDDoNiuzUErF/dPZguxp
s6tXljjWNaQYk06cs5MFd2TP2tzc6lO1LqlfM115up9qYldduG7jTXZa/DBaBAhO
NTZECD9v23qrKQK7hvy265IC/obKqbfD89FBAPzPyxc3J06R6u/XpM9KoVfpK6er
MZSi7ZlvfPOoV04VpQ9ec3qYR9iDeHAiI+UnbgWlhPMc+5N+JVwKRStwn3VGH2iE
P2doRB4KNfWEMCp04MlsI/a685eADlK46O3NPfjRws0QJeZf6KwdhYVY3k9P9Mz2
fPrkYBpfuE/5H0TthoOpBEsILZpSmoxHJWtme4yLgXo8uSWF8VmIROC7eNwY5XHk
A7IJ2luhH6H9HVCHumEcAV+rgyWJrp69YoWdbbI7smCw9cqP/KBWcmYa5g4/AyWm
lrR84U4pbFjNq02qEoDKIn1U/LLW3REgCKyAxAha7sr/745bmacUuc5Dr+agK275
8BqtxsspmG/s1l3/WEfFuMyJtqsUmgxemMcgc7h9Pcy8kIX9VdfnSuapREMzWQ+i
6XvG+Frvk7QlPyg4BZMC4CQvPqeV7UmWfaCD08MDJMQeTK7XFWBB/ETVltcWINT4
POCWPQd1o34RkIanIPQmpAxCS01lxYjx4D7oVQcTe3ju+HUnHjmtx9mLSAIqW5of
TPWqWCYuwNoQ2b2J/1DLt40NyjeBuwmH61yaQ8OORIFeqY5S/tJsfif1ykLEeCUT
7jbZo3lsK/E8uDTrw6ucSNEj7RbyceeVBgGgY+daWXN+n9O7pO/XeejvIvWyTsa8
Bfbs57J34pI0vCvl7LVShu15T47mlTMUCl+xkHtifym8hHwNj1zJnc2aOFoMI3h1
12J51BenZKrMlP75e3QSxfgliDuh25lO9QsaifeWkOHlPS7BIcjeirpwsic1haSd
Kdj3AruCSm1ZhQwhl2XL5eyLml4A5tFlZRSf2uraWuWkx+tnKV658GrDTprwa/zr
SUDa8IKTHpYVnALQs2WLgwD+0U8+dMYJIeBzUQPyGLp2wuqU5nuQB/b0SGwesH+T
pBmcmygNANu3SR0HUQ9zKwKmtJk9kklOAuuppYokkBnl20nJ13iV2TwDgBFqn9ot
PmCFiaN1bT5/p87ovrAmvtlFiFuLKVnOWUdf9/kEWBaMuBRBOYAhqyPYa7HXUDtw
AhHKIIMfbAu3+O6H+0275sqL6eTJ0OMOy/m/NK7dkXSslWjcQrQfqcIGKZPSK7S1
pDcrAkR4sxxMb4cXVYH5F/KlxMI016q9yyH558pnmNfuM4LbpzuqCEwvA+lguCbC
v2WLqCatm8B4LIPKi3L8+bGfj4E6dVok94ahYr8c/aydwriU7N22bTTctqW8pj5M
SRTiXRw9lAMpg10jTDR/nAsJSQCJj7o4nRaotNBeudneFJhGPBhmxNCqUlcl/49M
O5Y5zBut2abob2vD9+kbB5HZt4pGtZkwiEZtMGld5eg8y2Qvfd8dzrCoWwV/Ihao
4Q4P9sU9bNNclT4nxebI+RMOyGv8+XiYgg3oUD3a/USTGnxWVZcbX+VEOVWGwxog
BEvwYn+K7JArohDUZ2w2E9PPF/590LvM4Ka/E7lnpZt8v78ND/JZudRLO9FOThfV
5jkMg73aOdzQYDL1LrObSwJFitGFgNs9MxhshsQ5DypculKwg8DDIFu1pI8XzS3A
4tQI/r7VdRzqQF+2PZiUvI9W7GWJktz7Xs1L1GQ/E3/AnbPulHZsFiD8nBc1SPFj
HbojE2n6cvlI0xUh3OhL9CIlFCpl2k0D60G8oVt6PVjigW+GVB1Z1eLfYHRjUXTp
KMYMlzt5gIPQWUbGg/uz12ZqsFY6yKdkB0rquNIxnfYAw7ruc1UceiDTmjB+UWAB
tzQPLvVPhwzcnTwUi86eiWLbVtNeOSukznC1/TCaqghatWHcKa47rDeyNjS/UjNN
PnvdLxEtUSWLP4Tp5Doxa1K/C6VCNd9yPKXFrzXEZeWGBf+XJHZvssVFRDvtcWLi
FTE8RHxwMjRZK9usJT/sq5/c1r1tYSstZkY/XPycbOCcICBX5GDhI8qUMh7XVY1D
cb6fOhHHerxl9FhNuQIfALMh/DAJNLnCn9LFnGo3Syc65gfoha1xfNsvPOXlgE1g
lqmsKvVLv+9iBKOapyq3xdSITZbgpsX94CfUzoGcoeKZxuWwbi2E0gYx/QSynLkr
dqLKUVKwwmUCSEEwcOezUlpmrf6Hw2JaaLAHoEr+yolvl3jrEYX9dpnAHYLAtSRy
PcRfnS2zTdPCgNWajkTs4T0ItnxFACXPrgyjlNzpcLiB6oQezsqel8tuIt1wmMCu
bX1o8n6M/xNqncNl8NbuyGe0jF9qAPv3uc4YKJrzykVKRqrDTEmYZ/8rVrFTvv84
Oxr/7hMgygZz2ISN/aQIYzS/0v+NrIkczmdpyjJk/1nUaDx+wUHZzp3N0xCxpuAb
CGgRaVSIFdULsb3664ijMerYSU4f/4HWlV90n+f/uu2ccY6MSGi6oPUekNI3i/DM
zkv/uXNI9DSM9UaDLPIYrSOL77qFAccN2U615FJDmQHjllhQuPnS4lysvFtzTB/o
8rEIaSRz8nZ1iRyAsvgUy+Eg2Md6gR6YUsul/brLm4IprCd+GMKWDKX1YzL5WKhY
QEN7Hqipp0rdqcITY5nRiwnNuX55ss2yGVDlelOrElJztcApkLc3scVTssvjP9z1
PHy4k5PCl96s2wcG4PD7OJoQtS9/D/gzhlZ1SY3fqB+4/VdZLEeY46l78s1Y+HBU
LXpCSIZ2+IeMN693/x/9j6RtgHnRJG4G8k6zOeQ1ga98VAo4Rwxz10wnFSoSUiVN
Z26mL4vD83Hoc84+pc/cM8Km6suWJpP/aoOeQz2DS/SGNmLnhnySrQhHISGWBvSX
jqQrdqvuGSSJhQ6QK8ddcH0pO3Mb6L8Gd2+RkBA2xCZN18SZu4gUkKltLcJbE/pO
Sj2S1100c6/Z2jAFWTTsDsstWin+vwreX9Jv7V50u8sLyl7wyaKbn63weA9x2pX1
bS9+j7VfXlZGw7LOu8pbog8LK6dYjMZtjI5qk8sej96Mus7lQrrlyPwuYpyln2gZ
Tlu+mtvWfeqW92iEu/QwQ98+S3avec1KA85IgQ4p4CpGsci01vsG4SjACAuTwRbN
LCuaWbR3PPM9y0ZPPazsGbDTsKxXobVisW5WTrGGnTiCiCy1pHOx91wGtBk6JXtT
/x7aqozRQu1UGXIGKsdIeHSelxTmQCf4kVwLv4pj386ULt/w1Kapx99fqFv1LKYB
nvwdERwNQoVVPfAkqvvPwa2/szV14wVCfNmJ19bbx9HhHSlXirC0IzeQLQPpcoX9
EDQmSHjoDS2wAhanxIab1PagcHKSFS7ram9ntPCMj5LN6OugRImfesIj8lvIJ28r
CBEciI/UzXxG/2Ai5G6xHj6iJey1fI17IqIqwQpQIg8cK38Tms0hdEDvPRYPsfsH
OKLShUBEM3r3Xp9p8j2SeJ2gDu9RXLWKRz8xn3ctNS2Z/GXeq7MbJ0Kl3GvYL6Jj
iD54Lq9gTw4I+i0f6mxIULaDuO3C6aVQ/vnSKMYs8XITCIgZNGs5rN0OeW0rZSe7
4wv3sa1rQk4K1m+FdzzGa05QLfh4xYHZR5p3yp3YutQ+ZVkvKUfJmiUEzTeNctbp
GEXDrfrWWl4fIT6Mcc0azi3HFMvqf1i8qByLLqBY5vtp6Ra6l8X5xq8GdRXaLzko
E1ByZGFaY0ZlCvXqsjub0EojsmJqbW0TdT5bwtxoODxoj3OkCfE79rZv6iafuJEQ
EtVNvfbLvTpFvUL6363bi04vJE8LoZ+sJwFdTycc57uQdntB3iydBnc6fqrLXhCM
2syE5TlUUqJVv0JUlUz3e6bpP8s1fZtYtbrA8FSM1wSIB3pEY6Zy1P4CCVFhW7wU
4B2/qphpgMw45t/wVCsNgeJT6cuVFUAFRekUTRdodOvdQW8Qt4HQsCLOHxdiFIZj
ciUn1pnm//t/ZlkT7c/43sTkAT7ztSov/OQ3j7X3FvAuizPlHNLFjM2vvE7cpBXU
AF6v3/44v4BJ03caUTP7XlDFEkCigU+d4TWk8AsMbk0qoTrIT65vLfo92KV8wRrQ
WgdKmt0wkE9hVMvbqwjXnrMvtCVvZAG8mljEiXolnFkDG1mjKN5UEMevuQVWr5wA
KZqjPMrGg7RBH+05lleLhVX79Q65EJ8n/EvjrwQCk+iO/qvpiwSffPwxq+KAiOKj
285EIgZj75NjX8FGsMUOYvrByjXlvGshWNjTcr1sJbsBfjQMW7qldxfLQz3OUdAr
5tDWWp37XsfZGjzDf9S5q5STjfXJ7/y079RcjBFrYnLZqbruZ5+1gmKpNBcRfxLq
kQftB5hsRWPI2nfJYyVQH8C3dIuycacpVTowuHwna8KrHIAUJBQYgyI3t+9YShzB
Mve85l45Pw6eYWG5h+GGKwMLzVlqPSi1KYar5lETJG+PIu5sXAht1RjqwDqC33Fw
bCuy9j9CnbHRnkZQHFx4/7Ye1Nf5MNX2mtdMiHCv0R6xETSzbWINtBQRojHdXSGF
bxv9QbJ15//m46jNL/tqjTbk4nrsMBEsRGQAzj2p1L9ALBX3QlZ/IpMCSQ4rUs0K
J5BuTq3hN0s6cRnnD9A4YhLaLgmL9kV9/ksj5XT9gEN+HfI3++1khEw5gW3FGEAc
+st/PfbL4NS4HXucAMDy8+Fq0maShXHrLKuo2JKMbIkUVYaqm/uEM3YLMvhLw+JR
ltnkom7berOKwwLEoZri+v9HT62c/cRCmr0nTscYedueaHaI2iI7fUV/Ce7p1vhI
h3uq7Q5ozUbacNd+zVO5m5YxbO/F4Ee22DHNqizTolNg3WuYw+xZH4+t1ceyF4gL
vvOpyoMOpbTBdKYJKnGSD3zXNQr6iZOrXxPpZNN4mmujEBJtqALSKDhCdSmduPn3
dRZginCFt3M9BN2DxrbAtYLmMT6VCbzObeqJmpIgfqS/1oajVMfoApaBZQ0jisYx
W31C8N7xII8T4+PBNTejn/nOG+AkOlMgobJWbhzTmn3LxBp41suqkA//355I6kaq
/C3CpzHpzgK6G2iQaC6kue5I/0iMI9avPpJixDa/kWiBwPAdjLc0PZMho04K5ECt
UKCkC8koPsTsZPOdrQnRBmuV8iI/lV/eiQDRtNUac9hLw8ogZhq/iyUvAeBUjcN6
tv5iuS2eO9kxcIBFw0qGq7JaRVCsf7BYPX6AKr0JUbeN0I84pHsrIA9FUySvy2o7
l5887QEP94AetmAVpvlWuz46BcdGeU0Ey52+42+Q77DGzyFTY/viiIXaOp/ina4Q
zAPxaz6OhCKzlRt8p1y/zvDzyQ7Faq1UPr1jbU3cFcdRpKWGwGn8nBkBiHsZf0xQ
XpXqMkOFnG2k0Nlp97wuEehbQHuNQlR4OA6klQLjTm8PhKGmYWmKgsbIQK+lJG5/
35KRtxSEmN65bM6xwpD29RYYqNyfHRF5ttB8BxJEEkasDjzitjP8rzrF1RFTfuS8
gFlfkNbqnu0oLkFskMm8He55jp+Nfs8A5GTXeubeySDQb2KoKecZNhtrcrTUQRPn
fXkP9Pl4b1jqS8Pp/YzN6OcwForgpzTKDHI5RrJXaBwH/Vm2pZ7LbAYcGL6pe7Zk
wtEObWeCkNgut5EQYCcZiCQH4oaROfOrdPmwFFZ3MCxTr4Go6ZcCR/lYgIN4K1BR
czyertCnqHeattwWILe2IyfYYbOKsZ+bF25uY7y0iOFsqH6mz/+6VDlMTMSkUjyJ
pIfjB03oM18Qkwj/k7SLlg0TGzlYMs1B2H0r9glgULJzHnR+NU70VsP0HAmlI2KW
8MywtBs47gzpILsmwY291sbnB/7UfNdGTmFp5/jD0lrak+3mSYRnThhMCMrv6TF5
vZSRG1rfSSWOWXjgEfGPK4V0zm3bnCkvfg0lIdHvyIX5NZfL3mWy+GunTNIi3sW4
TT2b7Iv9s0lNVK/jeYCsNkpcVJhtLvrDr9TI7cs0bIm1XJsL/GfJaEIyBmzGePSj
caRekNNjYCO4jgxGX1QxysK4Lxm8VNxfwlKCeFHAPj/vYuJTzVLn9ZB6mRTjHyBi
rAD6ruT/YH1Id9zsnTVX9+Dg7jQENsdvKlgjrBfwKUiKP6JiUHRVFYiCqncS2El8
uVsfvPnow/eQxneJcGVOxoo6HqUKdXlm9LOJ+/Yirv+zN5C6dE+Yi4baRajadVe9
aaiu50ZoF8hkprqVC0vSTxXVMpul8zG/1ArsxZUK2WRiGwqUruaHmJw6RmmPBl77
nwnIbFOSlLAZZDO2XvEqCSq0J7A11cikCGF3bIoT3LulKBEQFJgleo5nGXxbTxwY
5rUYCvFpBh00gsUzfWnP9Pl4VcJz/SmeC4NUmV2lXcxOv8oJp6W/WVkQQBPVI1WK
3ugAWyyzrg+baY5YHAsSew5hbXoHrx+nY7oNrPEkpGVcb7NY2vr4YHSzp0hqKRBY
luJtloEFUa0PYTjsy57l6i8VENdiUUlTGserKTpCWEwJYpUi+PISXqhnGj4PMn81
akTzaYg4GF0O28SPjSAU5k9Ffwy/RoOw5t7L3bQPYPeyqSvxKTK9ya0LwWl0kaI7
Q516UdHOQYsyrL6XOlpmQZzmws8CvFIN4U49sOy6hPngwlbdRCoIEmFNM0RCKLZI
EhcqByyW8m2c+4VHleL+lV8QH/D7kzfaDpe/KIHYX0LlgOrMz455BsVbwE2NWG6k
7NRUnC6S3uAeDXlCVYGxLJkvWdTqO9XBloAU5jFpUyMyy3OM9YQvWMon/WmqJDZa
FFqh+VKixSFvCKcwXf0ge+xvWM/r7G6ZRw52MW2U0q1qg06FhFCujjNcMdiJiqe3
VlmgvLyCGDkDFVf3l+EiQs6LTuXDRlb4cYC+/Q7ME+kJoOp3lvbRC8Dfh8CeDHIf
8ckzM4hdd6O4cRImv6+XPF+hqtsjI/bRwiVQQWfSVJ7idbIT7RUCRqcGdItY7Y45
btHn3fAUkyEvTJfcbvWbm8ueHd9zB5yo4kXOX/AjrHGa9vhRZJgBbi2aZ+QuADuQ
bkl0BY7ZvaeHHfBaGHuJWgF7P73rB2LWVmi6A0NlMyehPsp9sClP/2BhE2sMPnDl
hnzJTvJdita4FFPNz8bH+HH/E5nHOm9BX87YdnjbwrKoEWSS6isuqFZzv7TS/b32
f1ga6AGWsUqD2GKmEUCHsiekugJ5NCCejR9pXkuAYtksyWwx7hB29ezfTrh1IMd2
Noo0iXSHPUUdVT63cvALlJ9ycwxeIf8LAnEbVS/+xCxqpMrQg2Ia1k9g4HOnQJ+H
6HhP99t/Gy6wisvPvx105YwMS7hs12r9+iuI+XmBc4uPcvWbh+JrKPqSoAmwDMaS
wdeDqevBbTARzfYs40amsEo6Q76IgEfoaVTlL0jZG6k9iTOudKQNg0/ZiGGoIZGf
zMQ3NU1AEK2FnBC4vKhldOuHeWMI0igszfryQAXuq8vzYyZfvx9qmEeEow5S/Sgc
AM1/9AwrqUBDozqQ4TG2vTQGexhoHDU5WByYaI+nQpyGHxevLn8N3c0SWXeVViU9
a2ysGLVvw2f7O2/XIFXNU/srNpnUao7nPPFcyJdYe9JcEaeaocwmC74I8WJHmF7P
GKQGzAg1oB0X5HcMKlDXlJwky1qBYCHyElpR2M3OKsYTfyTryg6A2HJ75Vvz43cQ
Cn07CUmWVklfiLpK8/sEVO4l2LG/+wvEl9QpKxA0GiqycRAuDdI5tX3wo3wBVorc
1QrGCMCcCyO6TPbL57XBqsG4Qc3inpd8evanM+XVko7b1b4OZ/oJSp/UlgFB+8Kd
3yNFkfihoYF484EdF+iX6qtJbsLw8TMwtMezvhm5GWXfXaLaaCmhWS29E0B2JxmS
0heBw8yhpcV2v+6T5+mzyQNZcDR1uF+MeXW+CX7cxT1SXtF7FkPVe5hqNe5Ac26W
7EurTo5jVeNcPITYvyUi0DyxuKBh5P9KRTeqZINEzE+93VDSCo8tVJV8Na9L3SfB
5hROPCDE7JKyIJuZ52+Mx4BqeTwUOExathF45Jx4SpclG7dsdc4O7B5heHLuGKUv
HNt/QY7HGoZgSVQ+uS+e7Gki0KU9burIK8+jZ6V6wgyv4ZT4Frcqu3JA2BMGimWo
qnpyJbbnmohT0VYuv1I0cAlrzZWsoLoAVxTGBCLYXyjBg3a+zSULkEHUmrrTRmjd
lODAxcKWod3DzciLd846rYdW2jIFm0Rf0tFQQGywcejFlzGz7+IeKZFCRh4MUOIe
Ml63LQ9keVgEk3djGxtPZfwvbtAqACrHRNNXQYkKv7kwebTpZ5oF7gBc6CEQR9z7
P3ZE8zSEI5b7Hj/iPvnlxvE7j1YiweouTNPI80HeONvpWLeQ1+5TVIjqbRHR542u
yqLr9Nh6fYMJrblRECJWZ2ZwHm5CHfbVvbTIQsu8mNLEKsEtY1uw+xJnBi8Rlman
67bcACy4PnEe8Y/+Ne/i8znE9R5Z9j0uzCLjCt2IeFuWtT+KZEyi5797BTSOgwzN
h/l7y4BjiJLroO715+X5J4Bn85IzuR1DHpQc7/EZvW+EzUQ6+f4/U8fQowqncpzB
fIzqIhGde36bgdV9O9zKt6u977zqGvMuWnSLv3wg09p7n+KplsF0OLtkBEWk05T7
Afx+hJsSnwaBNeCyl/9R4ULDjRIs/89+nVMgaazmMxT1HPFAYOMaF0hQe72/BPCo
xCr2sJWiJYzfYXBUTDO7QZx2KU3uoBQB7KC9QxYkU87YNEjc64cOm6XfhIKtCvYW
BdsjvBso4uN79ey2cMMDmDy45OSdezW+2gR1nFnofH46hVaXK5Ru+KS5GyN2Fjft
pPJ1Wobfs5WH3dK8tsVYi8j/8/TDCeghY3HI4T3YnoDD/nM6sEeE2dsmAUS+vrGk
I3mov66N0PtGgW2yCXggAc+Gtrhtk/rV/+7uyjvHeTqhYSWWaYhGeMOjBL+WJT2R
Mn5ZXM8mIH3QMC1AqqCGHFb+TthQM8cL+9oI6thwYFYBJz3DyH0E6UPFsLPKUATk
X/TUVXEsuWxPXJi3iM/PBQ3e3pM3rArrTkjmPzUKIo3dK3ATf9I119uSz3MZUpn9
bbDbtMloTEHWDIHcy6t6ygiEd504Dh1dHULypTS3CpaQ5lHoSGeCsvYBuFKcmdRM
H/mZX7VydUHyeVAXLac9xqEyqtTFavd8Q6Hgzb/7UB3ksy3O7hzor+3um7MwHWEM
mw0FYTYM9SfdNqeZB3KDqF5LOyhEwunMSckBwszCB3paiUW8kKnlyc5imkFQ/e+j
VsPthj61uwXpLkzrSfHcpxOodhYcvtObwvfcfnABOxAcaV/iQMzQptx+MNoHWK/q
X6b+spoN3QBRzTma8K5EE1vN8J3vd98ShSDvzHrN6j1sp7xk2vuGly3JL8ZCrCMI
EBZEqOMbB/y/iWTMeFQi+PliaysR8lUrXe3XBA8nyI8XkWOp03YUDGJ2myy0On6j
BbtKjupzZCkJv0E7bceCzEG1XNw2xZA1jw45uCz+hIm4Z52AWPr6kXYS09DFZg7i
ZIW70cYnvCE418GbqPIY00o/6kQvYA2U3cEwtkIRGR63eO7Kl1CVL4uaWWQwyvX6
kMbunf+Dp2iPVE6z5HW+5bBcQ3LxLN4EsWq2XKkW/v7lfy5BWjnWydLkJOsjoBcZ
o/gSQslH1pahGjz88JhZQFU7iVS03oJ1+KYdS9dJ/iFXFwXqV8t+gf4XudcDwD8A
80SE24y9Ha0JvHNZQTNS0pfr6JbEDj9BaY72firqXJjMKdYlLqjnjQPZRy65awpn
xGGroh3HkSctkcLvriD4H/vE/ITjEEBNXtGUAs00bAkyvwqSMHxcY/Os9s6/Jkyd
RtW9LCwvtXXz86UfStUd3K3rTjWgsIWPAVR/Mfk5fZHYtxxqLcjaG6UOpT0sBFXv
duboDYYNW1pFFNXpryym0vPBQOks90i5qkHh1YJ9c1cSncC0EJvzt5ioYmKIEOf2
Mc+8XNbSgSMkuOindKl8DKk9pQufBxTKDh1abDancAXFxiOU8Op7HRIPndPhIwvl
jVMUNB9C2isf/MxdOQBzmqh76lRbKi7cGrsrF4V+earPrezOFKMqtfiE4lkFQF27
Sy45Hfq1HPExwfn9EC/MwLaqXN81/bnA9s7+KL6LC23Cjdx6MrsaOHzHHtJDkWF1
6JSimad0S3dHWkw5VfKN6xbEk8AVjEUs49gvkyXE9wf/F+uVWZkQthM2hHpjms5R
dDsfMLiZ0f1utHy8eL6PEde3r5oXRsef89Tqdod769aOedZinC4z11RplxBGY4Bs
ZTpVuqGCn2D6EZZq46DMudEgletNoW04zx/4QKA8UTib14rS2tfV8ikh9SjqW7yX
mMCEylMh4mb6QOok6KF0zag76cCkUJ9aQCwSf+ny3LvA1OyOEYJCVOX+iIHT37tN
BqvaKu0aLTZ747quhwYZjgJE6gov+JsKqu3uQPS3obvQTsDTTXgkzA0cygQ3ZV9J
EU3BRKPy/1tsistUQPCQ4hnItRCWkodIqCdi15xwd1kTSd1OmfD3lUhaDujM0qFv
eHBJu+6BqF/K8CIUAvnJHxxsaULZtkZ0rt4qckZ23mSAcitN+LCJsIXrXx5g4zZ6
eAVZYE2UPlcg9kh8NhrfCAnTlWNBicJ9wuNTO1AVi9GOOi5z0E5TpbSH5EkQhhqp
tDlv3HIwtqtSq0Rt80DGanGG71xhrxn0/02Z9l0xzIXUTQV1CZ+w9J2QprhLRx1E
7XE4xHNZ/dJ0l7DvK5+qQnSPJDGvCexIkAgixoQhpnS/ixgNXVVPEa15lBlEGJcq
IgM8zf8zBUiCyOxuyrt3TY4Ihghrh+pSRJqXvN7ZnXXbgyIkobo80HHxy9n+Q32p
rk0QHSl1Mgeit1+ofKrfBE3WEmKDiYUOX4XLHKgaBhPsY69Q/E2jPrUMNeK71G0m
q8iqg2exQEv0m07SP8teNt4Aoi1OGTopY6hV7fx+qB56eKhGpgDQomh81+snr46h
tiqhQamfd4h5qAJkORGFgwc7LrLbE8S9uXtKbHcNBokJs5Vvnyq1g9o5GrMaKLdd
fyvYiCa0kBFwLUdE6fLKJsPwyDzs3iSwMwlF/dV+xkAd4suE8LAoPLoy3WmnTBL8
hyqUfJ1d83a9+iCIUa1d/uYY0ZJ3CUk5Gzg8vKRpHSxwbcvGww53QIzS/yA5carl
jXDpilrKOum5dDSElxeAQSZb3TnICGbdmNoYJ9Eu21xynmKplarQVbyZ7YaD4dQy
jBPEKmILFgRh/N85BKZ/QuidLle66gfKiaCQVR1wtnBoal/gv39MPVdImA4ZWbbr
S53Z83QkNopwBaPcoQ8yiPVNaPCW0YmLmOWc+tKTgoZf3WgoJDzLrHBEzPyjeq5/
cdDbhEuzC/BESZAl5FnKps8tbQMHZ7gBR00jc9cbPQxS1PUnoDphgmnoN14nL88s
wfOEsPBm23W5UueZhJyf5RN3o7FsfyX7ddTNRuixkJa3JTnm9qMmvRHaVPD/fTC1
gEtJ+8ZNWmlJfCXoA5HHa1x8Z+VsZlpA5gqDYLrJ6Mn9wJaWTJoRwd2UloIloDqw
p1+uYs8HgoxVEsc6YRrMRTJWeasijEU7emijRp1o8EJnrNGDp8COHP5R2MqAWLov
FKkrKUINqIUjrZwmxJ2uuRxN2C+lVmGxGOMLkiDupFhCrYNlZJ2G2oPqgVKpCnTT
f9SsEjYSUH1LMDSAXBfq86MBW8dIJ/uyy1/q0+HcrdYJxfje5NhktmASe21bYMzO
q0C2NubSs5yLox4T8mNoSCF93VZK+jI9j6lIW+gL/p7aHPmeDxC+Pko+LXwi33SK
RRozaQOoK2kPX3gROptPhmaXA+Im0+1/ARZU+9v2/1bOUZNQ+KVFE5+37aDNYdpF
G5FpFyC4i/89G4hF0wzlh/wUfesE00WvUbg0Q4dbJwOdh3IIYvhiAcQf2s0bsl3f
vOiC6dYVKYVZoCRTVXZR2HmT7x4HLG+gQaoLN6neTgyxBRp8h0sjAXj186JFcxwr
iMkn9l/8wvj4URbfhzb5NQc2BDAIEu5hargIyscr7SorrjDIkQxsFMpJfhK0OHsX
773KtYbkZYYKD6tltTxOSejb5Y9za2z2EoTMhGEkhR44abwqC7KtlGryEZyCG7Sn
O0hNjQRY05fwa8pqyMQ0PYP2GByJUTtidfAD4KoqvlN2O3pzRrDtdeixn8OEJr/i
ozanaZD4mRjFBRSR9jUqAFweU+a66kO62QbgO/UGVUzfzyrJbLZzu49rYbX+yeJt
BBCdT6/czuRvS5KZJNLQFLdfOOyvKDw2FH6D20aectpcbQlpiYip4D9ESeQ4un07
rt3Xvy7st0WjkFago47+SESUkGA8Hv/uXjSfjTpd0htfQg5npx/PnsFFi9Umorn+
BlRkB+7203IeA++XY3uIGwu9h4TEivcx279TrKFdAtnMb7HIgTHOIo8WGCxJiTz/
pwSfIFJoMUIW6RVZrN47qs+i09nJMyEVnfq5xjGLPsdbozwnqTTN8yUZXLDTmyPw
HnWqBWktvgaPxfETtSxk/idSLrDItIHW6CayLoSv5TznQgYi/R1vmqP1mYX2aas1
t3HphKrMdBYIee+aWox3diEntMC3B9619RBro6n6Op8kH9MqMPJW40WQWRkfHU5Q
ApPKt3lERiY/Mvs+iWoS+0bo+7CX/9TCKU9riqC0CqQifVNQikgqSU19EW5NNP6S
e4yWrAR2yg3k7F1OuA374z/rCd6bO3MXSZS9kuShKGbwZJWzJkTWFzBwLOmfud9j
t0ZEvUh8rzhQSQGDzWegoY8qLu8Ud9yH9xJI9RKJxz/rkjOrD6R5ILd5jBzf7Kdt
KgcYpi7gLfwCQ3oBdHHx2FhsGQOwY2I/0lPccguIYvJCh0yS43E4Ax1cBpgpWEw4
noPupw48woXKDlR28mjazwcuBJzXlrcuNhbiP2XPErGt78PQ22rztEC5b5Hkg/b4
WVpsedGw6rivdmc/SPtthXZDYIhgKlJSg5w+m/8tMULgXq+AJHLWJ70u4IGb7DW/
1BrFDH0CnZHDSpmjglJY4LE5H2NA7QERHr2AftGz7VXbBUf20ANe/43vAlyzzWN+
KRGplhQe1DKHyS2VOssVA3eeW0nk7cDx7APjdBR2VZV6ouiBg5Tb7mUfjniMWc1K
3Is9UqjONA2MGAvwdPgFvlm6DtCS2VwMyYxzKK3VwrVwjPrL164ddIBcayLeFhm+
Hdy3vC2yov9mTLo8tJDbPkmPR4VPyw0CDo5dNbUuR+1vVMGPZoPU+0eMV3QwkulF
Hjnm4gJpBBxBDIGWN/RgzJ/Imd3psvkqFbHr9ZZaCkNbl+/GflgQiT+QBfmRW1vR
rMmuVEuHS8fGsa4YiPLbWCs2hM13va5L8RDQse4fykG9aw+e9gCxdVmtihVoDi0v
odggInNtdiikO/SwvDrjY3+qOieMMk1CV9Q9rIwJXdAyZReJ8gUtXJmh6z5sSdDO
R1w2x0YJv81DHAHyD0VTGnf5dmjDbAuPjCcNxJ4LvvMZKS7kc/rs/siHSlLOkJa8
TEkTs42cOchOkBAvCG0N2krUubN7vebqK/1JW8IRv5M1eqscze0YREELuN0kjOJ/
QeS4+fiC2Rf780cV8wEKgIXWI3BmvPRtZdF/IivjwQ9BrqafbGtuplEJeQCs7MYI
k8ZhW23s9nigRmbESJin2V67onrBrlGd1iEqanTr2EMSstHibq0xXh+yvQJDQw1Y
8z4x4xFDB8zbc93tMZFPu5eFk7OGunkMnrcpUL073ddkFMVGSEvHtVpnNspS3pLJ
j4CFqMS5Yv3+WMdLIOx6vb8EcAM8Lt3qXEo/oTPJinXIfZRpGEyowTD4jX9Wy3io
0/3frFkg3t0rJsVo9pIF3Ah2gGLGnYxqxY3Ng+QcTMkF0sign/KshEkX6evkijpX
IPGr+LKK6C3QNFdLrxseXPIESYSn5lp6I+E7dbTTUVqdCDULiwyNdt/zH6kfw3qZ
xMdoS9PTb/nWoMOPCMHSqiU/+SL9kb49GSWVVECtSE1sBZ9XxhKM0uhqmUH30ziz
GfRbPntJ98hNKUSpm9UTtdbIZwXF2QLpXU1EaoWrdOVoFOo6N9ddj3gzKIDn2KBI
lbCFP+tAumJBswN5DRwAn+hybZGdwTfgEsqM3AHgkr7I6aN+oGX4EzauXjTXmevN
HQBXKchtle2/bmxHO1Aq+qT/sUIKV3V/sf80y4mo0I6J8cv8bUX1x33rnezB9OqN
+EhvX3xxkiaVi47rdIMODAIDtRA/bWXka2YrxAO+/7fU1UGBjXPO9Lj/+I1L/Xq+
Q0y+/TBcS5rOs1cruDNLHJdpgld0PvP4PsIvRSbm1QyRoQS6SvKeEnYG2Xv9lA0U
zGgswOZGijND45mT2WRVrbclXuhwLQpNpfc0rZA7X525Hm9qDa+dJtmAr60KDmGE
cajhsfbXflv1YSJ3UBHwN1uRh8wLfDl5a6x22hfq3hKZ3Xxzc9J8ujKME5XWKs9b
wTh668KbSH+w8OZASy7V/cBCzUVTQTEPxLbJcoAGbk0wxuiU+/hbc3ws4Z1eOqte
g8xVz18K2Ilus1Yyaw9M3jSG1tlphFM6zFmxBWCv90kOJb4CruI67kRk+yWYeI8V
5F/ofZ7pbKZLdGx0vTr0YKxD0RnkETE6rB6Hd4604oj3iQ84sj7qiNn2ZD8cEqqQ
hqkP8C3HmJJYstyCyilcmtmcUXWAbxl8nbXG93QLIcWZs89+S1h90Y/WPJaSlO5b
yOWWJQKz/aqHEkyH+aoPemeH7c7siXmqyn5W2TPna/gKgPHVSSaEh9TH4SQCQZSf
Cl5nSaMMtfhYMgMhH9MVQZdwsmuaXK9QI/LAjwIarVsL9PPfM+m2xuJ6+4SrFkCE
8EDGs8ZZLntFdLwSBzJGdr54PraCClJ89LKHQhZAXSxko58+cWed/8vjnWz7Rarq
MC41JdeWRwIjx0qpLVYdWiyKgJjUUBEVS/luig15qcTNYcGAHoL2QlPAzo3sfa2L
ohi/WOqp8EoDjFJaevd6HTSv26fnFVn6Sctitg4bkIwfU2qlfjENc2UrT/E60MwK
Ir5bQ/C8NWR269mUXWrIf4BJuaWGKVZ/ezARtLYiRq2JAYSRcbjswESRZEixvt0o
r36F5ooUjqAtoFpBPUDKaDamXrpJa7dF6j0f7xk2bbCpMTxD3ZEcDNJlYmY7rqBr
KvosKEbWKB3xatPJv0PleIZVHMFmIOPW6XbT++d5KC9+TzU5lOvFcVy6s3N8aDbz
OE26hFRcUZG9Xf1mfmRpxIBvA+JsYKZfuCYAF9Mwk2YM9O4/ZpGw/VJ8k/1mdsC4
j/6S+7jlFAfW3T+IuLc3dugCYwTJI5cykvhcFtkUmukNwfMSKhf3Ypy5Jsi1hhVd
Pt5s0zsadu/1v2ltxQ/Fjdz+yScdmaqP2rVk8kiq3ok3S0oXcj3aQduoZigxApKW
VYenGRqbyod8elcfzLAwJRT8YxDcJEHyqI0kEezJM92osz8gqv+Ql6lrDlGplXY2
oz474119GsfhXcqgaWFDKf5Dzkh95dsr4XOpa4TRWUgkKpEJGnd3J48pC4kxLguZ
kTxyhxMRF0nwzDT26DbBciBptrZC/OD4OdelxYRe6SEMs+szs1RRIHdDdqA361wf
zwl+uNyqMeXr4PKcsDYzhzWx82uEo1MZIRFXHyIzJdc52oUBboXeN6zcSgb9NLLT
jqZ5gFsAlG+FRjTO6dPSdKJbfj9y+I+TACb0OhT1V/w4xdsbPbhTvpnX8p5L//9G
V/gM7hwExUwuBOfhFDMOwfixlYbIyKFY+3uR3UGGmkdTPS4WcQO0yeq7P4xRmRZ8
YbB2j6LVUneYMOIpwLsCwXLo1FM98w4Rs8cAwAqeZmmYomlrSBnC1nBI6lr9Fl3f
Kqr/mY6ceKdt6JJTu+Z/C0qd6SEpenf6e9SCF8pUwN/4SHUvd7z0OVumvuauI2PV
gU+3FRQAEZI3x67ONZz7E/1fx5LPVDLDTTi1kNVJ/W3AZNGnGHwCLr1FIgWJdD2d
gdKxMdYp/NcTCxvFA76z89v2dOGzM+JTVy7O40Z1+RX78oneckorW88zevrUBMyA
vneA53hq7qHzBeyt3Vvfx9MT1GqFaJG9s7ydCKyIDX9lkawM46+I5Mgirs6JocU8
RQsqcFdQDb/eQHbz4ZFLz4yXZZ93Vu80nnG4oJ1KCogzs1FqviLwxskF0JmkO5ot
MZ9obrQfAzsnJkwlBsIXVF+mF8TRl2TiDkOaa/pBgrN5wZgT4F9+OPIkoNGn2Rrh
C0Ijyyk4o+XaBMr2wSQ/yZULY7bkCa4HQdqjsRZbP1epIEqWbEHQJ9bgxFdV8r7x
9wO0H8rh0pyGyQAcaW2HvZliUUqeQaf2ulxykj6MPwfQ8TzrjM4lRe2XHS3OsZcw
TMD3q2EsKCsRUS3ypfzllnBkmbylKQkmssLpdiiMW3aXd+d6Rq61Vm6bHSg8REtl
yyZJN2zgcNkql0MrznQfI/UT/Urr0vwr8g4f6XxI7v5O8gt+Vq+y93rbSKUzTwOJ
5TvwjqDrnI/EabHEmgdY/8wF4h2GBRH4nBv7HgXMhgyQWTwOTxrI8cIyCNDOrGzP
UX0tfD8fWT+FByLd4T3IEdG13vKsNAguALNEyRW9/yGaK5S+n+GbawWI3AwL1vrS
PPZ/FBgeyYoJo01VDWWfGuP1PPuQcaZ2fSKp0HouqIMqBazBp/8v4J5ka/mX+Y4L
A8DwdKHvO0Lt+eK5a652p2p/raROWnsrQTwCdCUsupnavfixhmkQjqXkwknO13JX
jmWwYyetQcWAVtSFju5+DaH+CSqUPND78tnAzFylwaRSeHTkL4g/DoAlkk08/EIW
rUOzRoslxLawr58CegH0nTJeVm1KH0zxIvkoSMwHBWOVwKnU84Yf2IftE57q2G+V
fZxOPqx/Kfl3J5hEK1818/3TmXB1wmbvWsOoYw7Nr3GoPx5RIcfjZviVv4+9gSzY
TyttR7ShijeBbFR/NmMIRIlR9j/YHKskIyl94LwKeiqRvnoWZpxGE+HL8z+wSCDy
3zqr6DdqEY+KE9YSp0Jo2m+k9EAulFupyD9yk5qtnWAYSJgGAblKZMV6PVIg6wZy
G2lF7iLZYYcNAsL/DgnNltFS+rsECZ7rInVCJwCqoBbYfz1p/B5fFVbqgMlsRfLM
jsuA31VXAuLz1BOItQUwJLOZ+i1/ibnAgdufy6IzGIJ7c72F15N6Am1f0Q8yUNQW
ElJgbaMIJ2XfNvxBoc+YbyXBAaVoudwAZksbwignJlCjz24ORSMmrbTuzAQZ4gF4
RUrpyHm9oGeqxGKycKVibQE+dh1ka6Vr69cm2PR/FVKrBXP/l65yffojkYNyzGIT
ErP+GQYrbFqzebPnPuYexw9BSRiISqJWBoFnR1q65H8+LTcKswSNSgFNaEN3WvYw
jM/JfiWXSA77sElVyGjD0ohL3od0zMxkFzxZucGT9a+xQw5HP7FUyvI9vxWa2rni
6F24aK++ukv/j3ryJIgrGzsg0d93kkr4xZx2QPQ4t2RTeAmAHpgX94jnnofwogEV
4RId8lZ4604KxJh4Jb7jgUZ+wnA7Q5fL4VRSC5HwDpKzgXO3TpenmDOBYbsf+Url
2/DU9K6rKedZoB5dQzTTAXro8FKoRzS89NLuQrL2fGulMgT1TqEEjji0CvmgMwgb
2l5Kw7a6LCu1r0iw2wYjnKVIfTeLxITBgvC16pEQC5Wp0boWStY89/iGIOezxBxS
PpMUixa+FtuYZVDwgBW7h7XqwCtmoS4OuywqnOAcEdPmBpj+Y576UWd1ASTV1hbz
HDBe8STMOajbxSxFMwms4hkTRR1Io1D44lIXVxVQySpToPEKX0ny26I5NtMrh8eJ
7Va/3SPyRJw6yzcBwLAUO0rvjKAjb+rE6Y8EJerqBpNVgVkm77NXYs/1NjJnOa9U
csPLU3ATciqmtAA8TfMC938Vm8fbBd9XGf7pGtYzPiLpifOGrtaUsx7b7R6flDIp
HgLE0SRP/25rZ1Nw5ZddJgqW93e3a+mFExXVIFIPNNDbyt5bwPalZhjyStTKbhfV
0DOX8j+wBfbo/4SU6Unt/KxW+45PaswIn64zFFSgNo1nAIiJNNeFu1DeVxyZOWoe
wYnoQIcFQzw0MjA74AtfDV7Ov39ykJOIJFt8bwPPTpzjYyxqOZkraygeRjnjBfKx
cc7W2hxUpfo4aGcgFvqttkokp59PA6SMM4ToJR6nzZ+5/WxkJ+NkT0WZTpXWpUVB
KrgsZVV2idNF1WGYBpO/zDOGnZP6PMzOsc/tGNlEYIH4wPFQFhOsvL+oXsP7HpFz
i+GBLcGzBnUlZfwwtfyTr7mUw3GnJgE8FLtXF3r4vTDVn2RHLhDuiROh+uOR1Xm0
58QE8BzRQFLaB3ZXNf8zPgyIavVWh+JmWkWUQ8o+iQqjzut5LyYVo66jqaZkecGE
0/+SZaQc7YKzk5mtXg172J3mc8PuRvZYFmr8S+szT3InIx8W0rDrDA9LWqqN6/FT
2uVnBo548EGllPaS2Prm35s7pWJy2k8j8JmS7fIYnFNscTYT9GIpq2zYHGv0ICVx
8VYz0eYJrEJMtjMoNLWGXAxJk39f4kK7jdtP7AFuEXyNmBlYM999cAodrcQGka9z
eYRD2KV37pRbojBXo7TU6aMkOTR3oGwfLd7Jh9LB3OU5mqvct0lUp6wUylLzF6Y+
h8H5SOccZh8m4ZRBCdiLutjEkDtQs1CHPl+QvqLrT3AKeRrDRjxLI0eWpbYy48Fl
snmoS26r36fpHx1Rxlwcx0zx7uiVOTYi8wLjnpEvjZccRjpgl2VbSD1O43jpQ8HK
4Z1vJ6wwDjdRezf+2bJ+AoJjM0u4ejpRO9VzT/h7boASU2bxdURknBb8FHCFfEFF
dLXHWVR5b7kRsoTiTzDrVuibc1CCdoGdG7PnpvHIhn+SvdicT0j9aKAnDUwGYS6U
ydCrAS2M8PUZ+MqNwD6BeT2Ecysd8wT+nqaIQnvCnbMGQgKmCS65Z/U/nC5cLREe
jb+G3VgKfj/j0NnBECGan9y6BZqEAm6N9im+p6L6RbDQJWlnJuR+L284fhGzafPZ
ASPeX1uFnFKgKH0SOy/V1NWqdSgX+fiuizIe6KCdQNkiA6WBR3zJgxEuPLKNEimL
yrjB7NpE1g14+2qY9eG82IErAGm+bsPI6QDPt6o4xLBhtT1QOaZvYc9X/WtoIIHz
RH3yLHtqscZCsGabsNWn7VD0gdkboUG/s1bKgYZEvc7HmsVPqj7zPm3yGEWlCdKO
jT0kNPs3RHJdChg+fV4y21VEJQaXTQb918vTBUg7L/sz6mc6X+YCJCQJ9DX7RKkw
D+PwBkQ6ytQ2TuArGwxzsO8d1M/CVHGrTLE+ArU8ry2CrE8gt7TGkM5zrMH4ydJL
3lynF6YxTZKuHe07fKhP/Y/GC2Ifp7UKvFz/74xNzkH1alZe1ZiWu+RgJWUIFdqD
LrQ/NAsxUkyNqxneVFuKkJBEr0nqEzCJ6Qmf5gt0GrIEQZ+sCi+ASP+Kyxj/56tu
Ucytt90JOr/Q/BsJ1cCEQR5eaNgh+s5MJS00R7yv2R4ztKWhTqjEoRVex6XPKGc6
MBvzJ0xkKMp4Bp7pZ3rhUHb/GFh+dYPbQL4OwUdULf9rAkAD2H5FyFYKdCwIORvZ
iuOTZoFFis/zheomH/q2dEoYijZCX8TN25WDiZRZ/WQvSkxZmcmskHjtvYx1H8Mg
8yNOi6MThLygg09BSu209CoU2LgvoN5ISjjKSehoACwQOyreu83ZzNGMFMqBbO+o
tRWwUdmcb2KNtaYs6/HqOIfY7i3NQpVAlzHLw/bZ1+a/KMRLamLEDyANACaTU86U
RZBNCmrSSWq1hBJQNZjTdp7uAf9kmJoX5H7pfByzfV95v05vUlr2FDFADYzB42A+
0wlaDzHQq8fiL7UrwvKR7ed28eASQRtw5ZJ26bLXq9Q2txivl7rZfQhq1MrtPb5s
m8cOzx14jHlbbL8mjt8u52pvRP7ta1bn0ageEefMkFZ8dg3pgiZLEuJUZcOTxxiH
brxmFJ8/VD0PFeSOTc2L4lUrWiLeDBU6u7wqh8/8ltuWZDwBOwnis4jrVRRZ2pmG
jhX0BTUZ9ObVmT0+ZaoidRX2xBSj9hi5uoLcTK/akH7YmQXMqSfxCPKvnCMHZw7Y
Ury2ruxQoDlHw4hkozMuOV3Biyzv3RrM4ifcNJ4/66wAgMEO3qsYIX/JH7EHZ66G
oBP+dJl2g+HBwBvkgHQD35Ai6Z1+JJjS/Mr5YlQDiLGB4uRk8SbwFkIx8C0Oz9ms
GslZYGzCnh6ZZUzuXRZKbHAlWy9x2M/A70CA55KRlyE9pLqmu/HG6gAJ5Ol96dIk
q5cf9pN/vKhDbP6M/7s5wnJjgW6JawtsWA+miXpRHRZpCoK2zFSGvM3g8OtZ7ct/
ygLAFRk0rcKUEqz/q8Csh6sGSDmFIEnqw/wSbDUO0GwE/j0gMPEMgWl+9J/hOSSk
ldZMOCQZInUoMVuCzxU2Y89TYZyGMTiLd/xJA+7NerADSXdBa1dlgMuGW1DFgjDu
c3dgBDwqyPSnIj2ghBGLB6klhrcoVykGpFj0IGL8PTfwdtkGTwf0JYz06HmAZIAn
pdonezLnOg49S2LbpDKrl646+oME7zLs+rFsYtNN0j9ym5Y8ZG82CdRqRerxpKzv
EXSibGQ90Nuh8xX1LgKs4zRUfjr6ZCMtmsrEik1vuV6RRt4CcfMbLaxknHGsT7uj
sE8OiqKmEPT+ot43KA33A2za2u+e+Aw11V60GfDOFkwH6Tzyol3izyN3TgM/recx
CFV+BNdR3cKAdDnOK/9N57VViQg0FknBtqibw5E7b71VFvUdIObV8DqY7nfPBIQ9
0Uc602NG7VcTpzeNKIY4A3v+VbVY0K2P++aVyRxRfL8asRYmvPSFlexw7zNYJC1z
wreaNhTwR8M/wF2LOoMrUz1tGq74c81p43FbG98mVsirDGYjwiEJgk5wg4lZEPJs
xKrjJCGHdROumvksV1FDO8ByyjplWMr6jlAb8FW9AXAG3o1TRd3vBsylAi4/kaLF
BciPX+TP8Kui8vpB2pO4DpwfWogDYkhxNf8gvwdRg+idAlcYax++5UVZmmgoUJ10
REm8BfoHho/X8vhWChDaM3EIo4mP4lS0M573Bjov2t9UmC7rpdLUq5B12qgyWUcj
A5VlLbWmDpMxv/nDJWyREWkY8TBhbZovFiAidgtodFxrCNc02a5hhXuzWQV+Q2wa
2sI65kasajMImZCpsi+5KaYqY2w+yLJjRzs1FA0SSTbkgoLOJukVi4j4Fz3PF8sS
dK+/DZlygdohCww6Qybqo3fhi5Y4WRcswO4baP0Dj42yJdgOR6zJVsS7xp1zoUe/
zltIpvL8NL8pTiugUMXa/uz/MHh98mlvhFNt8UKGI2ZpTUxHy8M8yL0S/b2TOb48
XPPUDWeT1O8B0Xf5ZIdPWUUmyaD8h6/Js6R+L+Zmg8Sk71dmBDgO334vYSOTYKiB
36CuY+2h4J3UyY7lT+JXebjkg0yOP7oxhsP3UyfBgzhtPOJzoxZ6Z6767eWsdTZm
3FKgvp1jAEoIC1Q7OL5ETuqr+rJ3NAtJTpkAuf+TILondGdAcuQmK+npUlKbVNbc
3eSvDdWp5h8qVx+ki8PxoULNeXq8zR6jDgU5CnE4RpcGxummt/HNClsClR0M7aNa
2q6yTerXZxktCMZJaVWesgQItESowgZghUfwIugjuCUqspmi7xTMCi76+apq2LF2
fy5iUGsQCg4d+I8GDxQVlf0dYTW3cJ8un090JEhJcF0G2IwsfwyDbZilVmPhh2wH
E/cv6BUc4If/oUah7idX3c8LFSzXgKlaHG3Wm7QkqZYOjmVbzaN+B2buOLuiuSJt
67E0YWx12XNWZB+n9h9NFc4/d3rrvlXKcowfvtXqPbiuMg3bGwfeGO/bj/fqXTDn
XgM9xCDBMfEXuJe+PqiIN16dwsHy9dAHywmU739EqXTaRJ/6BxyoDiraXC1li6FB
83oSipyB1xFA8MVFNqnwueQovD1WvzzwTeiFyakCDzzCDpME/tYi13zw8fbGNpNS
Em2QomtqLwGH58EbQ50STOAxqvfbdt5b85XpiaFpC+91aDDAHvsxEE/y+GeGNyge
ra+HBNHF+rBbO4+kcbtJ6HXGzjERpx8wuBY2glzfHvu12HBi714DOKx/XRODdm1n
so74sQ7ZXwGRibkPpcbMJOSIzF8vsrl56FNTqqtJLMPdyAuYAQQMoONHGpOTfENG
KzrP/wrlW3i8NMbZdpZIXN1Rd0vsw4rw+Z6bxlxveZpP4gwXtV58v8K/WNIPOBwd
oynsiII2a3qhQQXad9ObNMseOn3K7ItQyHFVx9wlYZQg+0yn82AMsxueHAiFZL5g
GeXPk9+ZFC295uUPbfkWqDf9CNG3jhuGl+jtmzo25BcyRZmr80CGATHuuihRRupt
UbIZFI3X+QLoBkB3JIFItN8/pu8VQztY4n4pFoTKX33pXbnv8ZemOmzZJ7sO2tZ4
OjTt/7PHiWMpvyqpfUzrXGSi6WAePLytOzQ1nj6AYSOt3SvZ6//sPnmgoviFH3tA
IAJoL80cqmppPgJPzVEREZeXlK8aNeR9lrFmE5FnWn9oA/f1yai3psGoEeZEtq1n
VfPvXowHP8k1w9Cw1o/MJh6u51/UiJvLcI+i/RLFuAg8xLech7QYaey6RiSkzvwT
m/8NMvM3ouaAqIX0qgyqoaUP3TsuGBvdxk2BhToUI8aFPqKUk1DO5zN+n0mPX77w
/yDiG6xqPGq2z+WVsmhPArb4gJ0Sv/SNfsYbONpeaEc/TRqRhkViEKinppOQg/MV
WzRZ3C5g5VSCaiyv3Q9ErwG2JEK+NwTWyj7EIu8+J2B1irCdDKPXdrqM8OWd9J4+
6SKvlwl9c46NA3S9XojjDa05CZTKHLjR2yPxoC6e85u7waWJDdcAjaau3X7a2RxS
WwoqZDp0sAPGGpV2YotQJihxGmRk059M9Wdsl0HS1eGzCvD1WrbZ4YDtjshj2/0x
s7UoU4TrWB6tYZhQDGbQAtrUGW6HDaMChA0Pxbhn552XefkMU2lJWMs2XjZU42nO
SPYBtpXYpWrNmAvUe0HbKTtzzb9jS1Tjtwh8M2ZJpNnFcL3xbIAGE73PHzC5hwn9
psEngNI3OVm7qjhW6N+OTqLPW1IBmCNBV21WGQQMQ8xJdYsQWIJqZcxDN7zcmi5D
zfjadOOvIEutGD6bc1093s83qkZmh+nK/tG5tOb0hEBgnYqN6FMEOrcbAPTlmKt0
y7b5N1iXSpO/hhnCBTUr+gJ5f1D+wTcvKU4IOdM4BvGxPucBAygyNbE7+zuMk8Af
S6Jau+PSOESqBBmESYr+MIriYpYCunwORLNAJFZUI5Uj0AXI9xGiVUOuUv00ehpA
BiNC6eRhF6QHugL7SUiXNkBdqu9yzWKKXWcxy8lL/AtxUe3Oni6n3N0v4XrjJ7HI
SHiGDRU2s4rInkU+840pB2wjkh5agekC/xhiA+5tjSLvgpeF9a0sZpRYALUgJ2ij
My3t/brww9QYltpPI/RyJTJIWhsDxnR1JnUOpd7Y7VcVBilczHzFAtv266o6GahD
kGcYWY2NJtIB0xiqbW+NhG/xQtaAtjgQ/BASWCvGyZtu8LhNCou4rOwK9hABqFbH
qF3rahh+Z0CF7H36JQ7JfUkb15G3xK1XT29+bZO/rP6mRg5F3UBKLz2c0BibGZ1z
SCoNByystZU+9rpwcDfPiHmAOSZ0UgJiCDG+dds11FGrWtU75EKniVCTanFQh+qK
1qc6AA3da/6UatPbXKY4E3bnaNumcoTAsoPQvLeBssRzyW2WBZzL0RS/SnkMSGVd
tiGOGWSH72XAFTsy/OkrqYAFUF7IOM/hRbOySNIv2nLQhPLUoz2RuequrzwlfFqV
Z3pWum0/EBQZoXqvoGItHk7yfZhQNJsjq7PF0OyfcoYvcFqi3gvKqphV3IUMAk8K
aLnNAaycqWpY4Duvt9iqRAQCWq6ey+bYvWWh1pN17pESrG6N2kBTBhiK+jaxQkJA
/BkSxF8seZ4BDLc4Ozc7f2eDY/2+AzrFq3Q1x+ZbWL5MbieePlCpve/bRZOXpiyQ
qq0OgJanmBVcz2saTNx0p4LHejhcLY0KTYnXWXGSAoYbfQ4zOGSK+MLHCoNJ9xGJ
/svlxdkzr7TtOfU9C1nV3eYUC3s/TjKmS90Z4J3EihzwfsxOV6JYXqzRDxPNnGpL
SdhLXnlY+TYPpdAVzu+gK39nf10WKp0csWtVZ4gPNzWscdcB/7pLUB3M1UJ1AT3k
WRAO1OWCCwHDVYKq5a8VfU0FXXGJ5ef2bHr5mu9Mr7S3e6LMgcU/Rdrfa9KCtLgk
OdydOEYpIbb2x+REJpzvrtKHG7WXSmRO2fkbgKV2xijlAZN0oF9+VC1HgJBF8jiL
JKjJkiiQesOiurZlxbS4gINtMqq8JygC9CkOL21NNwGBE2THWqGL6tb0hLsh6O1y
gYZdeGwIPYBWpaSB7Zor9HNFhA+Mtvr4rnTpu2uKOMYcXDjGn6mXuFA06dZM3KQr
G5ZUFATjb3DgKvePeoKK8P4fOmMj1lDqwVkFLkoo2Q/oMpfPBR0Zw1fcys5sjRj4
Hl6W2bvFbeLOeXwjCZvWWVZwd1LZj51bSngMyMcFTIV57kLzY2VzdUuzTnqv7KoF
2MBhxZQyyyR3tYbchj20aDH3h5AoGgW187Bi7CE743HwNYvFWcJnGLb76z+rJynV
SChly9DCD/UdVD6Hnbyrjl9Ymo650Oqa0QZvXxsdHQXaQehE6ubRwKXoZ6tr5DOP
uu6AsHpcy6W5YLRFlIXX+pmqc+Azg0KCQlsl1gO2o35vKazy94yCwbXB8rM8RdXc
dCAnUhLquu6FJ3m643sUZIB5rCOPoFKPCn6HYbQFCFnNyu/9GS6WkPJPJNF+Qx/s
Vffti2hZCgnOiCwFrmVZtmbdCp06u4r9yRej4Z/L7ydF0UO8CH3e03X1Jj/e7mJG
7AGQq+/VGLcrlqe+lmrh8Aond4wMpc0u5v983lotEGGcfpyCuyEAf9g8Yh0tqNX7
8sr9GmpMB76mEXKYPBT7Ovd48Dg7P+kwav3ZUsCVOXXXkS5njFGut2IRee7jEfAi
0/W4++O7a+IVri+oMJVip+2fntq4TwubxfJI0PTJQmNSF4tXFK2ri3f5y8oI13wY
/W59/SCXsR3c1kYXVjx04wcNLQarG3ofINQQP+s5dXofuzvsObV3SpXtDVw3NsPD
qEI6cWbflp0hRIggPl05fl74TI9Qd9BBsrBwzJ/XnRIRSbCiXreyTs0Id1CdFVdk
k5zsHCth2UTEhVzu+B/ILYqCsQGctQoj7LLypT5MGRASFmxTlc+XC3pTTxAIGPmn
3w2hd2Hl6o7kyu/jtoRUpByQBiTIIFWDff6aDMHYqt6oDFqhzpUhcvOuohXmvU4+
5nsGZhaDLuzyWOCRyU+L0oUKV/l5Xsgp+w0UMYCZdSrVROpZWh19b1gPUrntNJnt
EFx0Fnukgi5K5VKElODiiOVr62JawOqbk1yiB1h8PC07QFk8Ot5++y4kjvKN6hup
R34LrgZXT5GZCdlRsWpc6GzP7PY1KU3sUZEjUP4Kt1Z7E8uZArXhAhM9jBE9conF
b5Onf+n0kt3vnKdpOJNxCKj0Fc1MCtBoG4CFru5YfQj2xjGOaYvFdruVCZaFGNTW
oM1vn9Kr+3LUIx+5lyj9tpxHuoiWvYy5LwA9UCd01pHqgO27hl+2zcFScZ4kXzKx
JdKsrI1dtAn1kroK1Y/C8L+wq1Ai6nDzxUE99EiNPAWUe2w8HbTTn1u00ltF+7KC
EFIK9kARpTSj+SNS72LPU3MX3LpqqmswBb2PBeU4rqcz/bhSBH3+FpcjJy1Yzxq5
+wgMp7ZJyuTe1lSR0LqSH19TsxnvBFeQeoxjx/BxiC7pN/YnZ62L4j+YdtbdO3NU
0+ZXR06UElDnLjmE7AG7ng88r/1U60jcpwX3w+nThefqEBNwMZunm4GwTiKbQjYt
KtBq67ANaRWNqIX2RC9Ks6pCqeyJChvcyi1Of4/srjAD15VC2WJO1GROYEnGo6sX
e1LX9GJkufGEgaENnRDUJlFUZ5Rr8nApiw+jjc65VxRxqk2jazbRv5urSllDwWq9
Jtjl3U+gJv9IRTH0Qcq1nREwoldAByqKH0yPtNaaZX5S52B165ikHsCdCyvrBjh0
frk5cEO0ePGfLVp7tF1s/yHStAO9Ai9xi1gUbSsLwDWZlrWHjrx1mPodO2d7IAxO
akOhe5MMClFA/qgcnaeDfJTlP53XXZV4YMav2pGJc27DUm7XnbYDurK874BR8Lob
pfdeTIjvBSDKWtn8DvgBfuP84pc/+jH3oNMHN3s2XwhddTqfIdDaYDFVDcfxCU8Z
yGX/fwrkNBNr+jGYN/JegcZnUIV9alzaPO5T7e5T9PL8HVpOdVzup/ZnkjZfD2BO
5kD7k8vcc/4fhZ1T8XjvIykLbz2/i1sK4HCJj+tSk1tDnsC6ikAzcru+NYdca0d4
4pjqpAI6T8yBEfpkvtJkN2SKZ9htF4W4XrHSzexUtwIjw7f8Uh+YrHFLGSPL+Mbq
VfBSkcEQvVffm57JQ4g8ZAqHRVKnd25NFOBQHZWt257vYxu2xxUVwVIRlaZv1O9A
e5lakN2ahUD+VuTgQ6FL9E2TuFsd90PsB+kIo/slZe7aT2hhBiZZBSUxIitxX7+2
sS/X+6s77sfwn+Oby3O4UPzKqMmX+4y+S9dscIUY3uvooxwCnG2XgzgvtdOS60LU
VTDVAG8qQdttfeB7Ysbb61/KPYzuTeEP3byRpLF7qo4WI5DrjlByqSWbEb0uJl9z
0QeWs57Bc7b2Ce9iuRN6R8vkxNmZJX9mEG+XmgU80D5cjiifFh0MhubqDmplEcDw
yRGiC5O7PCygFKIq7mE15WHTbbCWLcgMTujY0x+DkL2h2ulNQRnzD2JM8pMk6XJr
dUU2Wze+lGV9Z1fByUhRvepjX3bczum1Ab+88QIo8sDSRm6xq+K0/PA9qKKXFEBH
x30puj7WInq+lkd988eaf8BzmArkAlpG/FufFybuyyZ2vOwrKsHKwNDrk5yE/mXU
Pl49j4xYDO2IdbvucH6myi9IlVAzWXn40mjYdDyFl3wzyAQRvrE4SmB/cCtFEA3d
Si7wBHGwnMLL6aSs372msT/d0TbkQ9M/IEUmycqy2Kx6/xkoMr6BhnM3E7qWdprY
arTq2ZdRT3lh0oJtnXa41tP6px/uBbmhtnYjiY6jjMXR0v2/Tgr4DVFyzen78oMr
s2NWVnL0fPYmszMtLf59nl3l4+94xfKgdi5ONKT/pwe6QxLL0oWGTvfO62sH1rXo
MBZ8rxGsHMTaojA96Z7lCe2hubE695lfk/ODF4P5/qTmsK8ftz7L3EXbUbS+QBrU
tZaBFVqiuJ8X1nz51U30RjNzID1KtBedZIVeTuqTYLZkLco6FZ4+zggAVrTMxkIu
JBTHLmcRtSAEGlquaMp2OJgexV6P562ZRR2ipehAPyO0Yj1IbvrlxuCo20atRSFR
EE1bChMvhFfM41JRsrdp7+3FDH2OhxCz+GcEmiIJvFFb6zwmB0JS4Qt1aTBiWVe7
YDC6Q/YW6MtGjjbblmVKyD6r3lr7iJ+saNoENuE4vvWOh5i+c1w6ZnWeGg10mQ51
hpNeKP5sFTnoBwQIGLcNAHu+B44dmptmKYbCCljJUD6WFXCqVW2afoWktyYOfbaT
M2SRJJFgPjOI2WTFbs/zUb4PZWmt/tXKGeyJRTlsuTyrrn9XER7/wm70MvNGW17i
n5SIl8kd4tfuJOBU2tg4kT0CrI0DwZ99e1iB8mztG4cz60l4wO0S1kHrHne0ZoJ8
LaO6Z8qziKqpjD5jjliuf5NkyN+CDHdwTeSnhx01jnE/5zHExHyQLhieJ4KwLr7H
DVXY0R8fhEhgeztHWjKJZTL7rFke74tPccbm37CrpDcGqXOJUKdr8zRo71cIWDrT
QQjbjMouUzCxLn+TzWRoIX4Zz7QQssH+3Dsip+/ZfHM+pu+3P8bYMTB8uv4WAVck
CPEP9/1fCh5F/I6A4TuIKEgZCBIdoexjmu+xklysDq2AdTqvh/mJ1cQ7JjDs4Ik3
6xd8Xc05kxGG95HUkcOAPe3th5uYSGkf3pByPYcOwHgBygXzUUaPdxwy8GLQRRjV
wxLNvt6SJzPdiRWeRq7zOj9SNdTBy2+xP0SzVlOc5Bhp6Aq78PxFzhM2ZGfQNKXU
mMdms8zntYdV8IawgeuJzreu5W0n2EoVIIFWVVdpS53umBWt+Enq/qHFxeXO7IhK
XpxdyYo5BOA/kNJ8ORCrfI3gLmG4+mXcuD7gLMGh2CcnND+BJ9tQu4wBZj0UclhT
zW7iFLgJJRzXoTq/rHdfpb4A9tTHCDXfc70GmoF2aOL7EZyCATpP/I4TLHTrCu1j
1Xl2dLwgFXCxkGDtQmHElxiXTiGmyCeQN+y5OdCiCoDSK8XUScvn2W9iYetFN2yi
S02vvkmAXWAJ24YrwhYFnD0aR3BXgaUYa9Uc80egVpZMBrklPhOyCZpiAuTvZ6kc
jT0ZW1M/aektsiBIgo31U0FsAR4BE8PTav0aOHOahxumus8Onk95oZUVObPb+/tr
1YefMunMJakhAAFfb9QIVh4vgxQkCMnyvG/3DRwrnlZNVce229TK4p/lPoJDyJlG
Cp2H8Y+qZLL5W1dcefwu2vpint/yMSuwNXnP/I+wAh6PYQVD93Dzpfv7jcjtnZEn
zhVHdC4/WMw1J2b8qdT+suZJ+EPuRhyr92YWDR5F7L6G8nxCM48qM/K1ZT0+ZNi/
mKojwvuQWmuBZnJKGxMetncJ6rvUtgVhwgnCdyEBNQvMtVm+5ZCsA2U9gIGbgzf9
fIYEaWnavjZcOxGDPgiYYQOaoT1e9tTotUH/ceyBlm5eZjnWMu6Mzu3dEzzXkQyi
GM4xv17wzyaHKGtKui6CLZaVYdz8OvSp/snUMAs06zkFaiSPxTTJY+w0jDd4Tlq1
OlbDjj9fAO9JX6kop+wKd9qrLWdV1tN3s8P7IwPt79h1uhQXmv/jJMR48o+7ixR9
KH1Bv6WQbSFVTlNjMi2G6GTWpvY7fWSRTFzkv+N8NksJAFDS3/u/I+I3TbhvRXpj
VnQ44rqRPSG10htji5CHYfUn6UzLG08XL48mguBcT/aCry9+ooiq0V+/vjcoScme
hPirE0Cr6ezBrhLbozO9UoMTv+tdNpZnL1Pta2yy3YeMNIkcDxNl0JrZbjaA9pKV
yo2Iq0Gl7CE+5coLuLn3UIhvUhtYSfY8lJHBNV/DGttBEj2pcit+rV2B/ihPOMdL
SPJ99fsrt/tqMejGljK7IW/H95lLD5sBPZ2DFMrzLBhOxjjAAszpv/0kqm9TkLm2
n2tc5kmMCqDgKEFS+uiKNueceAx3WauyQTf2oyUOJF69mrAxCYii9kUlY41ocZJB
eaLJQJBGP9uS8X9U+bdC/oDru4caIItDaNlaAmyBE+DEyRUC6bbhqUhRFdx404V4
3vXlQrIhWeI3RdCLSHLHMnKQxwm3W+L027tEFLPPzVkdHRwIImjBOrla9X7bvZX+
Vnt0s+x90k9KYDSQ3q7reCgRj51cdrqD3WHEMgU9M0O3G0NyBrB+z/IovGKNpIak
3ZxgGS1Pkhq/MthdF1A57jfCuN5V93dRSxoaj4Q5pZ1tc7y1Ck8EcBp7JIafbMOe
RLaIyv8K7uMjXA7nWnzgszdcAibjjm9z9mx4b0YWkxXHVF8wKvdM3rCs6ZWBOIff
KqB2/VSLTZIz0HOiyrA2VrN7YIlGJ5PH0AFTRd1lwC9EERIOFf9mltUngCn2bE6i
eSZGFlx6vA+C5/kTqRoywU2jFjdGhGBujl1wCTL9tjH9LPr7ejelXpiTz4RbAcva
YJxEKP5Ym3fwYy/EvaoQvxclqZhz0Ju/m/leutnU1eWYAu01x7rdW+xcCHA8kj99
XrHyMlZ+0Weh2dtj16IXU8z2YY2nrog9rpiWQy8YtPob31wPMYi2M/51C2mMxspZ
Fx5WOiy1wlfwfkeQjj/06KeNjinPURisaJhRfeN/Xri5/18lO3lUt5ozDfzEA/O1
/ZwwdZ2S2GwxqWJDEc9qKgdooM/zr4FmnwqvpW2Tt9h2OQ/kTexTu9umwZW+YlLV
FQjEtEjAj0AcUDEJ4xzo+OX++XehtWi9L16Oo3mwmMTZnFBHMgmN9LVkt3f0e7CI
pN7CaG+xLRxIqiN9aVpde+6kWvAfhZm7EaAALFsdQCfrZBi4yk8nwjJdWICtg30/
jruOcAvTu5nnYtoZRa5wPFU9+S4MgQKblUiV0PHdule69m4G8fjcc+HaocWnU3lZ
8vbIjjfG2RugqrwX77fMWNtQtr3327WUKXrJcUSkeyPdZjYh1kUhKH8nr6OECaLd
3Er9VMNDOkWVcHDcLwCUclJHVerdo2m2hToMNQ7RvoONBMQV4U88zFrDTjz4OFCz
mvetHIYlXd6frpzueExqbxdEDUr+2Ae4PHixVXGKfpm/v2mSIwca+KL5iqnsobc+
9eJdDBTJliUWmZ9GDiUF6/4Dj3+1q/LPHijkJjbin4GHmd1snyQhmTNIF81DySta
IjWSBSvDsfKYl0OcvZyYwTJqBJ2VbotWW+630yXngWCDsRINbcUoPQPEkbnh3SIW
IqHPW8joZrF4DZSr3xx8eBxpx/dpgcBKsqGKIHRNmoSyU5FRykqRhsAvF1RWfIL3
Sg3bb4NqDUHvC82I2WvYwoCUOEabWLN0HKE6VConYJco8/GXpBRHWy5mgHP0R2yY
QyWZkOhqXsPit6DVM/xrdkXlfClk3MGf20KH+F4dctHgEs6AuoD02O/g2JHObuMM
xDgM19mtNXUkmWVb9irNF9+ag4XopVwclUUCi6oPPryIOkMy3oHpRitrQsy+RzXn
4wqxx0Cey6IDWFkU8InIg+zYu7IP4+2T0ufqvwnoUFTmNJ6szBdtilkJS+pDmITP
yw0yvbjmNOmHq7t9XyQJ09RzIxz2sSBB/U6zBzJRPwCJZzKUvmXr10TpU/eocTfo
BP+6tEcvo4buYCz1ZadLg1q3LM/tj0ASW5/VlQkCXukznRE/pUTXyf8B0Ob57JoX
+gWwP+ZGkevV96NSfHVJA+OGIB0VymqtCDQTpeSAZEU/teXIcjqDm63+IBZTQ3q7
mxDJnvsFJNqkBGlkaVvvI/iqYXSfaowBeBf4Sa6GyoqRXodpZ+TWLpC/udCVA5ca
FfcbsIp6v38qssfuxgUZ+6dSX/Ir/YdNVceStvDqv94IfOciualmencfpS6feCLl
I96sPh8PUUJXjjfLBOvEYQCAPuQIvnd0kqYKGNORuYqjThLP6zpdBKFABwndEgIs
XC0BE0uuSFTeynEEX/vjvBYAUOd465ZRRTHP/5NBHaXDm3ELK27VWd9JMvjMALvw
A/PMl+cF9vnDmuPt22c4Wa271Eq2eDmCKz8pnhjzhF8LMNNdShc97l2MmlucZfWr
f0WsRH3z5eonoC1HgT7/zm8FvIcXYrSxx8JTDmV2aoiO+DjsQBc+FBEn9+jyET/L
nMI4zX8r1BpW260mTguhHjKyjVJOAjymrOWI6299spQXcD5qDRG84DDT9EPxisv4
uq03rBt236AoL7MlDW8pboq/hmqu/zm8GV6o20eOfzGFCRZIx4oLiXtIoIvY75OE
if5miRxRT536u+GijlswuDaSBwsRfipO/8QzWof54Eyjm6e6EHDAM31yE69BltxG
YPhUA1obVqMAMNfbnKF/feyjmnmEnxKgRTrXscwOZldqHl0gAaw2T8mdHtmU04Te
V7IpTzVI/MjDjnhnkRNkJradpQNw5qgWI6KtK8dS2zUjKVB7dUSeeVvGFCYkPKJw
oa/0OiVnufObbR7/t6fo8ZJVF6nXb26aCKpmIp/0YVUtMPVZILw4R6V510piOeOF
dq4tYXBTkPZXj8/GuvO8S5J41avQW4zRjYGnNXz8bIvAXpcQLZ39CzhWB8Rog6al
zf06kB3czby3xwYrrAGmYRqi9vnpqgm/k+F4W8+cKQp+MEh9p8Fz6xugf2vXw2Ui
zbfjPzUANoX605mW7t7lAJuUG+8y/Ljwd8QSs1NnpVdiaOaGVAr9mKYGv5Jb6WMq
UO/+UoaiXslrAdBdJB0zPMMxY9111SfGmm8pEcTPIAX2jyAnj+V4JxL1NeQelCkk
O1Sn2uDbceMC4mEQ42JZxe8ObGG0bbYb2yhZJLTOF7ennsf5/cAygjzKEyU30yEl
TyKEU6UUMK4/a6JvpzkK5v37TErOakIZc3ElFRl8E3weeJRriFrDq4oP+rhQeYIm
hkj0oo0DYcYCnvM1j3J+T/CeRMUp/Ci0omjN59d1bMF6BEqr80E2PE1MFdE6co6T
OviHzdriyte4AlFil9ptb0TmaK85b87pBqiFoFs9O+Pa61efHkhHtrZkw9v/4OAD
4qrknF7Gn3vQ+/Aevkiw7cRoMEDk/NWCluLP1m/g7a7jvQW8FhBZOvrYLkmusOuR
P6Aysjiu2GeBGHW5NeyFgU+y+kZ3+31gBGJwthprVK+me4iiDuEqx7cqpTdoNcSX
FVGDT6bVCsTYjSrRQzQ/bhgdM1G8bMmsMvQjj1ISkxCoYxD/mZOmnXxMVEjDwJ+6
3SttvBD6U6xiCGA13LiX+l1LUK216wvAvkcpeWlBDdb8TpY9zOOisFICbNhzdP2k
nrU+1+zUS57pQTUPYMmjN2X/7EcJIiKHiLUhJuVueMcH00O0pGgyUznuM3K2NR3d
Sjsuqu3ghY0qSc+Yexs74KLavbuxWt/n/y/SmZVxFvKQEceiZmoEE75hN+eEU4YH
DUk88BCCJrNvRruYaMZViV7aIt9mhkg71OB1fFViOFBQkOzEwua8lT6PGRzNECTg
K8IQIU/e4IclRwQgO2T1ehQqBmnNWel+Mk/LiTiRM4tCf2EA2V5QrGhaq56biMhr
XjqZy1M7GVpLDzzTK3XXTbdslmYncniWooEsAW/ulmSgRHQeK7pG0Ye5+pxsiZ6S
lyoPKoOAe9pX1HZDYvXgdGTX89vwDp7d3giNzN94W3tGkgLhDp3jUapfsJaInJ1r
tTuQ/y5Q16d734FAa68sw6fC8xN5i51ZB0wZFHUzAMPljsrtEkrEP9YyqejOwSSD
5/i5jG82BZKDTDFiH2UJLr5+FZWOlpFcFWWk4rxQM+6//Ri7rBcya898WQYHhDJt
qjplTemFtBGLrVJ8wZrOWg+dipwE92TW3bIMsL743W7XvCTVNMwjHw8sOPmBW5hh
dBbdlXz9fNx+VjvS4KhxexiRe62in4KGB9HRWCoVpr8/Ou2GVaKYyx28CueojOgJ
MC9FKHPGpJ2M0IdUHp/5maUpNxDEXBWObrh395CyAa4dOLSFj9KbPolFj917wPUH
rd9zXdz8rs1IJ9iK0ltXbocmPmMSx0U6OmgXeVtj1wVxnrIUx/fXs6ol6kQYIrNg
xiJ6kaslmQuGrPwraJyQOKGzxzhwCcebTZq0O5KmXaDLnv1oOrTnQB2t2oKLm8Mj
+DqrF5btXhi4X85Ig2BMTkie+YeDKQRixd3+ycxx6cNnSXkdWfDGc/tK7alvf52m
r+kJ+hOavzBYfQW8SWOf7wuhdHKfB4EsqLVQpToKcZESZKIoWCADBbcNgafOpxQ4
pbQHQZ+BRhMR2fndzCPVR5aWQ7wiqPtiZpenx6kmsAU0rDV3V9wUuJh6Vnp9YSOT
OHclxI5wr30dfQYyZ17hsD3w7P803pjA7PnVHm11Aj95VkPyGuZ/WcwPXIe9Zwky
3Jx0tZQikg2gy+UuL3bp12WzQ6Zzd0WzlOuiPO5WYshpIpkz40r+yGuh+HkTpJRW
1Ay26FoQT4YY/edZqKDZ6pA+nu8Dx8Ih69VffMNt0iG9c1R4d30YcT6ULKPRngo8
N1C7f11gsdnMpiLqTwoZLE1QhV4uIRc3d/j1OkOLeSwmSqX4Ie5yCndhaSW6C5HO
GFSu7TR83YMpum8i1lCrC9F42MiNDI1XcQmG9UVbGh0ktWePJyp7MxKR5G+GgFnh
04tClHuUeXVcTuaYxN/hECXJsj1RPStqoG/fpm/qpFZzzdkwnolGlCX/uIY/8LQC
9t/Y4TYoUeVBzcJmvjPpADbTYZHQRgTZEHsvS//DG1frBGhFnXmyTpyN40pz1Zyr
0Vc1gS39qivFjAPVLlNYZOxkUp3TJX91Q3DRQYeG9rQMFo46mkcctUqRPLCnCbOC
jZ7rXmziP/6vKbc9oOxsXGVH4V9q0XgRifdOtfVzwsRJoLKTMYLFOBxoTsIh6Xpv
+jiA+hjqGsxUZ7Dh8N3EqsTWFZx7YdxyOEg48IW436Us9gCoHRVQjpXQJRVk2PvC
gH3HvLqAc5yfDiJ6VCxxa8z14eFo5zMjkZGnvvQ0aoTEzOFzh9H9pVLfd5tPGqki
1S6vRP6LKTj01rUw/jlfIbw6FpT9KQ93JGtQnxv5QGR5wPBqXNkUjk37tmn9Uoa8
RGv54qKGR1OUlIPiKm82+TnltY6MjH6fSy8ZpDLG/HzJVvGjRxYsXXGalD6Lav8m
KWYWtgG9Ep/jVz37+VUS8AYWhiVMLm6wlfB6gqKueNjOkJ8GGXJGAjNRKmYDT+I3
rSlkyTzh9KtAVmS15gvQ/3KPNTe3H/P423iEv0ZEMx8ojz5xj+Vyw/Gt1oL7Yziq
EousyWrOLeSz3XeP+cSLRA/SATrvz2AxBcr2cdgR45R+yyzLd2OFjQBBBrdLCPzQ
RiZGLgOUhlIUQWSAiiNGGnppa/mJsHyo/mBN+1FftrKm6aPrArjeY53rLRRzfSue
H0E5/UZinok/brdE5MDcppeMAoRQBNxC8li90WayGjpmvGQ2wJ1MSs7R6c3yhhS6
lpv6vQvXXSMxJ9eh32CITpCiAE4iaMduenb77H3rRvdlBdMFdQHvMpWPuEwK6zZu
+Vb/IWRXt5WlCKTRm3YzXhE6AtY8ZTBwBB6omh0Apx27kqqCftZkrF92zpxqTfA3
ByRVQIiW3S4Tcw6zhcgaiT2HPlGxfdxQcd60gd7Lv43gQ/y7WuohWS7k7kB3JYuk
40NLIgdccvrxNnNsBuYIBM03wXeM6TIlsoDAapreDxWlItdoFsPyZgezoNAATSyP
b3OZOV6jEzCy4h/WFQgrZJ0wZncnNi7FQm9FJwNM1h1ASid1VoQq2epliO8aZ+Ae
mm1aWK4zKr0S13tLSVsnK7qti4hTGPrrZGNy8P3IAT2bg1t5yd4ht1H/krIqUYpw
hXSZD3MT3U8fDGxY+ittUFl2k+/jyp96AuQR7AlktMBNBSh7qPAh16xNv7iPF8tI
D0hpfoX58/hOnDRWVFG8Qh+fY/zySVdptUVZKjdoKrXxyVJeiq6amhlN38uqgMGV
+nF2Es7FtsW6CUKCM5HoeU3SW9ONtLKTB3Sp3bgPVaYfOPJClPZik8rszIdRO0/d
m+HrWHX6OhRso4j8DUUBkSVwGTQub95t0iYXhl7AqNAVWWqFCa34e5YuvZEaFMff
5j5GbYfceg1hiRklh8gz7H4iLtPY5IEIKORavwifUuo6ptFH9lLwfwc2VoP4K0KT
YZUFlhybVeyyBnkjjdTy2UaWBeKPkZbtYoorb7nTo/RYWXI2gd9e+j60pTZNe3nk
BDbWIOnRzt1I28imSEfTEhcMSoZI89i3UBF5HQFGb2Mz+2ZLIqZSN51E9amyjZm+
A4K4Ul13H4KJRxWEMeS0d33g7pVQlZmVUyW2GzxWGuM9smbXKgkY7vEGKcvCAOsj
WtKdbykmL5KTbrG8QqiE8xHGmixP9QBSKYPcEsuB+YDRUKPLjjv52MegUXoLlIkp
MI3V1PQDpI2efleTlLCVGLn4WLD+lre36lckKGef48ox351t0SHOLUslp8PqQxEv
EzPI8SXWcyYj6z36s1ySoUq7Zq3VCF38t7a0YasZJt/5V+hnkAZp7td8M7dbsHEE
Lmb94dJPc7tWF7CwX7RFlIzZQeF5a0mdQc0qNMZ1vvPh+/KkwLNgTQohtVV52hgq
Bv8ypRdsePe/nzL1kO22/zlCL2kcbww6549CZt7sYiIMB2WEENi4g4/9hRp7Biwo
ZXLyYH6PvC1feetdOuWXOSH2b4jmFa/xjavOMLSe6WMwK0fRn8npKdk6xEoSkY43
QtjLCwagnnEgt7gMqY0LhOCLBbHRq8UdZtpw3pCAe6KzK2GM9aucmqdpUpc+CzP0
WVFktvYT42UyQJT+MBtnizyLhhJ70/7MKmZ7LlJCi2dljHVC6VQrn7TdvNYKK21I
F3UNTu1frXQw+hI9ZDMm0/9UN/B8qzEtsXsb8qOE80TdsBthMhEdwkUPgumwLSy7
SpzDvMhgc2kUQZIp0aHlkq6gngGbgYWV3zWE6WFoI7d7Z0UnAEfjGsU0RluEs2hG
54GeU7TmnS27kmwR+GUPjQVorbfqaF38/K/RXxsr/iakmpHyms+hJYzrNasJO6Bk
voGHstWEhvKml+SOJi0FuwEoG68P9OlCMAGW2QXCdWHhnpN31JaI3yNMXnkgE4l7
9st5rFj8FBlOt1fN5AfCCQmJAwTyZHGYuHx71IMiAoMVloYfkIcAI9v38KXqoREf
wzjpZmEN+qcqhzspUaG3an6KPFoHNUsU5vAAk4dUBoYYqIs4QWBNLsGCCa7aFR6P
JPvIP6pL6WodpVs5Rr+LOqOW4cJVNSuN+lHwrhJC6ArfMq4wUhVOzwfFM5Ci7BV0
VJfXinfSz7Kn1gIecbsBtMK8IC7jEmbT5U03XWiJuD6wwbmQERGBZ7t4TpkY+suu
CTh9YeKukX1h9X2fCRgLESJjP3Jv8ySZFFSxYuViVftG/QRS9hVxD+uvv9jKtzEw
NCagVDiEG7sxcUY/AzGDO0Tn7CrMDtKoO4stgT3AvOLg3C291s7S5ugj9oxEK3YF
D8sGyeG2oyVN3lyvCHQqM1ZhYU6Zf5czZwpiQ7m41vXQnYj+m+Ow/cCs5jyB8/X3
Fa0CoEY/ElqxGiLZWOfUKp9TFeZTlzhm2o20WiCQZnw3QGN7Z/JpOy+46A5TCdEQ
B1xRQPG+mPi5c9EgezwoLb7XHzCpE1bkOMK4BoBY/1j1iMbEN0muinsBjx7ibnm8
IONqzV/hA1rOphFlfBIBE7q4sB13/BYuUr3QleEOKSRslYZcGWxgwAdOncwQkKDB
KSuZx77xwKKiNrbv49UMvFuSV+ahqnCMt9VzgvggJFnNzVVHCcunNDQ/YXCgwV0o
gaHQl+E9FCzz+mUc90TQm3Bf0dBUrnD8FpP5OoTal456bROdACEjXUSAjKfcFW0u
L1WRURltgWcoisPeHZbCzum0fTX6AirfMJZs/DsuUlFpTXSGyYymV4pg9uPq+1Kw
LD13+sT3nsE3Iccns0NvpgzmqZ4Ibd5IGdMLJbsLc7KLX0Lm1F0rr6bjbRxnbo/2
5QJazkSh5gBG0Gd/Cw8xmw1K9Mt+EXY+zW7ja00pG6fQp6DCaJYYggDcjBhiJ/Iq
qVmCt1XGEvr6sqA0y8wHLNoWVRQejI8AD9s9It4qHaFmCgk67d48fZVpOwRMAWb1
JPoKdLdFYM37kobREZ+yNF6a2ER0vXdBkAgGSym4+ypNgSJjKoOgMqjqNWa0MnfH
N/lppKHk5Uewg1euDgNa1m9rOhFJC0QNQ5pBDkRde0BhCLpi8pkdY54NLkS8YZsD
YkTpy/PkxwoSTKF6aiD/yY4gmJKiMvel0Dil1lL+oSvDtUrEdnq+OSrzZyD5zFZv
HOicNKXOQnLJ/daJtRKyI1hVNKom0FHdIjpfwgpphS+QR0KVmvowpvReiG1qqH3c
2epTtebKrvUFIDrs1TOwOmNLYKXF29MzICgyhJocU8rDkVj0J/wVMZs3mw8kNh8X
+zQ757tZC+wlWjfmNSNzM9S79RpY9UuLr8R/gDya3bZTy2CWlOIAC2TCc9wTBZ06
lC5Wc0kOeqmFU5lwztIIrsnJdo3mmP5kXOQbeFVMu90BlAoFlhTd9Tx6KfMJLflq
1egaOlF6nv+bIA0U2aKzxR5AMGNWtckUunXTBLoXdOIf/4P1MucTtBjb3zpJj25b
suYIs7aG6dKXqRFzBBc1YTz2yZP0SeYQQHaMIZjQpZIzWA80+VC/a/6aKsiSyIQY
gwqbPnuo/SPI+qjiBg338FjUoh0duGU2d0P7ZpuCHXGxK7oz00a9Zx10Q0ew3moS
OtVXkf9a7TPw4D+rXAMLLulMCpH/5EhEhbcUeRphY/6bsDa05XBj/WPFtb7RJ27A
Ji3fjGEDiSa0MMkgHN6zy6xfaJqZ8CICuLlvhakPJwkvQS6aEhCDiAY/5lKhAOgY
FN6FqpcL3RP8q6lJm7fcQ5IHghGU6hPExSOAMMcYh9J+WycE0qmb/Np1ILiNuflW
KaOC9qtBks6sTXKvkUz6ggkWK0cX8EJgtbDuDUIAsXEqG1GMO/2wI7PCvOczLDFx
nAHzXyHTTyVUEDaOQeWTf9gB8a5RH57XTjFuFvMXVI/U2TeP5+jkhQ9OWS01yYmW
MCS7MtATAqZ1+dGz0j6RsGTs+toLuOw0GDtlsXdnrswjmnmke6It6h4wQdbTZ3Y3
uNt/mPavUlamq9vecUsPJe5T4rcQGHm/QkthfesAxeXW8CxTDaZQpCXhHVgKsf9C
kgHu5sOEKAG+JslsEmRl/vA2/cJnQ9j1ixIqreluiU8Q28jxYbZmDfDxqVmPDuvt
a/mKJBK9nxLhnJGieAcJh85IF+PjpweuZ/sxW+jdX4ctblbrMx+zxvY0xg6c6rwA
rRz5pHaZMgWNGu8hW2Ak2Iac+t8qRnaj+WxXhYVyffnxOGUBCMSWYHZCsbb83yyE
VH5k/U8ZHHlTFs3bnGYAMVbScshDj2iWunZH6pOaN21vaBVIFnXSZPCYRGcAv1xD
FJ4K7dEZYbzDNhI16pedsrNZ4lE56bREnVIzwnjDc9K7O/2TuTBIhdmHZAD9w6RP
9uO8gZBvYSLYKM4sFI8XNrgw/b8fo6jqWZYPu2bZcUGr6QPlZgteBpe037om0lUO
C4PlKdnsj9rlFR9rqkpzNwYq/timfgGAAVjh2zgT+MInEAb4gJvcxDxWWx03hktn
N55wCEpgMl3gB/nSefs7J4DtM2XJr3ZalWegjk8VENFevWmYPzOjjBFyB7JzZler
E0PjLg/6A3VBMzNE2kn/i3SioeNsk7bKLYuMB2w3AovxkOwGx7yJCRtNoI/Hmaza
m2KwunnWwqHEgTC21wu+cpZIdDOvBDSVw8EZ76MQVZEVRI+lI5bsKIK92XPrV4Nb
j7lFy0R5ki/qZYafy5fk+UvsGx+zukWt16OIS21LjIvG85IrFvLwOtraeflfr36l
FfW0925veXRqa63qUDJJW9Z9rgyhpRz4nV2GmMzzta/OXWLsLC79jxZepOvFKbB8
T2VY1scd/oRGMgLEPjKjsEgM2+hqKaFxRhgPrpYe9zlP3LKkCUzmN1JsfUJPNX0A
YbJBoWIQuqKQ8jkctx3XY+Ru47R9VvEUhtt0dYPi1vngu9qSFKY0kdQy7kUxzEFq
fhCzPK+T9V4nqMxWBGELYrIaIpN9G5NqVi3kFhjlT9hEMUlVb6yBm4aGzVQQnvHT
lReOMEI6lRGsvADLDdv7RQTCCbrB05Pwcp2CNfLJMhWIsVlSlaFxLI52LaH491ZC
KOGkRlfpoB24h/OxXmpG3WLeMrqVRS/EUUK2UxVFnbOvv4wt3YJcgZcWC6YdTHG7
6TL7SNh+ZM+4z3jBoQbU0hkaHYo89l3m8Qc97bnX4rXYYbk11J0NBXcKGxcDaxYV
b13Agp6823BfEFPqBG7kKNyZyMokPSc47DADSfSrdxf7Rrft3S5Ublboe+wkBRhg
SfcLiaJAaMDove89VwMxzPVmVvs+UqsmKKdejVvbpttdr6dCwJz0CYQYytFKQ3GN
rs5xIPElgZqZVEQWt4nxxZsWr0+8IYOOdelz7T4rWSC6kHPkM5XMP8nYcai8hxbn
8bAyeGU/8qBoq77mr0ZP+UZ8h10gqc6pvg+PK+Mx1WpitlwQJJrIwYzs3ABuawi5
9eanzLTv7D5uczFYYA4FKN4Tyht3kJZGhGCaJPy8qFUQeTPYHvrnRvZI27QKkqoE
YSTdIUUMjbwt5CFJq+nH8RoBJz+5UiSM4gGSHuO54UaMU0wypDDbWr76RbuF8Wei
oZwILOvLdfc1HceUnTadnaTu3WJ/1yenOezTKndcc7EwmoSr/cD1pZL1VH5AUqCo
LkQzV2WbpBF+Nvgepr2XxzRgJc4QSggSzGzal3G5WJbXUmz6wEyzEOAImewSqah6
T/MiqK1prPtJBv4bs4PiS1ToNF2BJ+lOutnNBtPCMcm7tw5EjAUK0Blq9CKyEC21
t0e50Owgd8TA/M7cZbm1EZGstoJ5HOWyoyIZNSv+weftOUPABoKfGq+m2gZDW2Ms
ntm0ITrNlqws5ky97w/DQXoJBk8C2ip+7GCpsPV68nzSFz1lRklYTDhddw063//M
nkEoLDrqIbtTKa5+wOofy0VEWhoWkAf7F/yFs4J56J36Ukvo29G+xGtGaTX7uXe/
jVRRiUNdysrh2URaYNcagYJqPCc8USXs5sZVTadc5Y4JCKD103YvKLXv1LEW+IRx
Uwhd7QesLCfYZk0o2WKKf9ZoQcFubCpZSj8JvpXLcAhNZYJyhwR42rcXl6gKMC96
HujSEG+S8AvELXsB+uaejMKlFNVi2Q/sJae8ybVILQSr+7QRAr5asVtRAE0fxfOn
ydD5IF1CrENJVWrCGsCkPWAi6/oZovPYJYtkYE/RdpqauiEXBUZ9guIhXRsOcZTf
NKu8Q0FTOQ4Lmxn6qRZ+vQWHEWhcy7HWlp5kM7gzutxfJWCSgzzmApx8E0t8iqKY
MDtS4s9tfKdiQ9THg1hI+F28697Lur1voSO3ohRcFPGxIDFeWCeJXumiyKX3Y5v6
e+rOun+GgeH7343ICozhG10YSwBYsIRC3SXJTZJx3zcwTtYSCSdvzbzow8+8cPKR
CP6Yg4mWFKm/aV6SqA+jXEk4ZPnY6aBAe4/QCQDnWrK0e8bbmYfccHOXl4UnMdee
3Rfpv9fNFOTFaRPkjIIxHF1C7hd13fYzCJqnMTA/MqYX0C51D9Hr9HwBK7/sATPk
rauhO5KCxI47kCUSQodYYtjWxEwbpNRzX071x0Mz0B7ogk2mnsfgs2GxZYp6E3BI
ri/o6UWgBhts0NI9yOc5CgmNxG6HAoJIxACC3b3vJ1k3nmgfQfz55jWhxpLfa4SX
DHnSi7D4IqSDAIGOvDQMyY1mydjk4/Ic1U8zpB4TIDmF4O6G0e5SxUeO60PJHPhN
u2+Od+/u/XxV5oIsN3UezFpRBC5I2ZrDHz9RtHRkF2eyZpu8BtKlEIfi6DED27Gj
+5OqiHsr5bLBUbnnj0IgDOSQZktnBPU+tnRHtIYxqOApv/m1Ab9/ya5KeSVawJzS
6ylr3m3zaEXUS38CSwfkg7p3X7je+QqTRTHQCkjziEzMXNbtE7TgqN0IYzyvbImh
Dl7ffxqnd07YLDMSEXdTNcM1H7mzKhPanqWsXB1PnGvbThrMBHqXBoeXqq+PhkJH
ObtCITsFrNI1oBO4jTMRlpmpJ9U9S1krzAGXXYM2M8BShbc/m0IcKhNgQAuVYzex
E8WOtYFgky/CUVjMqRBhxgapQf2EUrqJhKofKol7UjRwXUFMfBicQtGZt6/jtIBs
K4UCaZa1Bz2uBOOI8bzRRr/ssGwVi+8djuS7etWgydD9ol2LsP9FttL8wSmATfDQ
PVIBstSmPWM60OcfbO9DjEWurViw6Zh2nzK2dSjGOUvhhg3bRH+Ydvx07cod4AxT
IwAFBSVhg8Yx9fRPETxGjyY/t2krCYp53HEaxdkqvGcX7a6Cy5NUsbMQtg8yWzH5
rqNsPvBrJRxOkjiyO8I9i7XBAaBYnZovY1BbxomGkenuDl3pqcVZqR+67h3RjMQv
Z9ycxs6cJHnRD1FtIt+eaGyS71VmefF/B+DNIvaaA8LnDP3TY3MVsoDCmfjGW/wp
82gHFWL7pWg1Ld+Pvc4oaN08QHVyZ7+A9gWdNH4Tl/aYCoMg+MUwT6P+02tY1pzH
Dy+Y5t2/VChsZmx+2jnJu7nUGRb+miUgF6LOBZhnt+G1/G4IVSRFX5t73oNl0IY1
8tHBDNWbeP309inNy5Z7eXb8GBY4DTRlahoUWDWogZ298DFSVnwpSemXf76+2VkK
zpbxGABXlCHQn7BQPKBzAPoliAXNnrUpr+Vp0g/JUZ1umw1ih0c4Xxdn11WYyrDY
xTLABLJxcjMAeJud1Q5vEzKemRwNyqaXKzER2pd+AZKvCMGAKZj5JO4M/lSFGS6+
cxmLWgkuX4Twg97UlGNGS32A8cF6MwIxs1paU0G3BNk25U9YQ0H5XcRKQjFOnCxV
XV1iBJSv0FA7tMjRLMg5UoJk59VWnyC/V/IaR67OPr9hDj6/66wgzwrghzmqEjcU
/gCquLPwiX5Eq4eJIgDbMoDRNXgLoXYJAKkLzASHudO2gwjAhtpkPfKIhxOdlbdA
Y3F9yRP02L/BguUZ8w22oWkR9ExCItrWR4KKwA81V8/hijaUfGF7kAP4qcUKphMm
Zc7FIPdYLRdKyZci3AM8s+NiplDBB4yh560l9qFOdIJgYk13by8+LTiRnLx9KFIK
BscKXlUh8ySDX9judReUQ+9oaY9MZLw+1+rqBpxSk4NaOXHJNTFVigBrTv/Zx71i
vhePF9rLtFnIHFscl5hRgD+8FBciorH75CZtsDvRx2nNvf1dMmlY0ueeVqtaEAz6
m/+o5Fb8y5MS/lrldKzkXCoWa0scTd3G+lO33qD0hXqnaufnpaFHm5zyKlJeKD9v
FykqUeIdmmtetGCOoPmEMlBis3GS/lVOZPtNdhHIvyFCx0p9f9MPh3F0+0txKYme
aXloeHulBnMFPqvwap7UQ9RbLgqPbsAGUbUHWWPZVv3S4ho7rPo1aopM6j64C89K
U3OYKN4tv8vpgXTg1Qf8RvvOx0P3RvyPzY0dFDpd4pC/XitEq1mbYKq8VznscuoT
va1G1o9HV5upMELhgv9FhpMIjW5iJwJhAqPO+KmCa3A7JCv2VZ2GfHxkLzaTtbOH
dHFIw7P6hFwSxfV3iYbsjwtadG8gPX2th3oI5uhA/s5Ev81QqIgvNZA4MbYEuRu5
nbfQXsNSVk1HAggP/Jplj8XJYBHHnYbZCtSsSy6TgXblxFiDNy2lXYoN7KNzHvUS
k53CIIwo5YMGTAkqWA/1w9k0Fy+qCclZwzRuxttGgdCF8BE2eSg0WqxfWtXL/06r
SLqrVXMQb7BaLjgxitSRrS/rKP4Ifv/GQmvWUdUaUG10011WDh9lLolRr8E5pnp7
5MpChZeGQETBML0eev1w8wliSafUE12RIZdd1Ui3u8JhTTHSVdX0iYDvaI24Am+y
tzrrpof0jIEb7O+o4GiluOs2ZlvauV70UdtR9alW6gSF/4In7HUPDwJea1/I0qqj
Hqe/Nm7+iEGHXM0s2b+rwq+TDHdZd06zI1vXKfhf8c7pqngXmklWNdPE8a8sX71L
s2SZ4V/PY6o+UZKQIxxKsLJBT6walGfr8WVyrSqRExgt5vekV83PNYKVjADy5dFg
EiHNzg5DOPOyHaYqQ2UKtjf3iKJOpQ73zREgFybmnNU6iTlWXG+wLp9AF94iqVqf
SzoEvF6//jlJ/yg1g6vNaPb/lg4TS7QSIcMaMd3tD24Wi44qTj2LIyb6c7me6Lwt
dAQUiP6gDhJCIatPMOnPevCEN7TwC8oJwmFejlPLJXwyxy0nK5u/jccwNH2aG3gY
0UyxykLOpFcdoy1vJK5H67gH/zrYF+h7Q0z203wS/NoHNXIWKjFMfqgR12VqVdg+
etqMdyrptAjgTMMg3Nrbx7y5Xpd2r3uOY9dfo9OVYsQWqG/+ihcRBhQXT+seF2Lm
tk/o1sa+jG9nI/TU+qp6W4V0aWoOvwvf0z9cxcf49Vz7BNbIQ3c9RSDo710vrkIm
IYSv7C2/+ph+ZjD0U+lbGyfh08pY2KMCa1cFwEML8p4Lad9Tlk3S2IrDOWytFvKO
EGfUAvptDJ/7kprI/smjap4P+Wp17TnVIOdA66jzzTp4ZpwGvucwb4pU4cR+deHJ
bL6+1DcC77mFj5F3Z5w+JtuysOhnCCWf/0KnTfC004I5mxOrPacDLy3/qJymhdm8
QaL3xRZ8C5pnEjlLx7e+hqxg/1OSc2pBHPxjkxEEwKwjyhzX93uYNRwuKx2RkZJW
gfVGrQw1tIMN1uK9HDptn1Wpnut7bDef7ScVd+oAMDFWS0g6OXLrR7+al2wGnsvp
jEHt0clxm74qLFvgqRuznfF5x8OGrbMPFdCjQvnvHf5ddFk9qWn9RV4JV0KonEt4
86/aAg22rYjvNV1B/EsYPPqAHGmYscK2Cgzw/ItPfbkY+F+cp13Ib6tpmiRF36oK
22vgLATcow+BHNewQCNiQgNWGeE/UuYVmCVLSteEn0DEBS2MHs80UdDj9KgqQ1nW
p7i0tPk02w9Vt0uqhJ63tI3NbG9BpvvRJnBeapzr3lT4l72AgxBXEj2j5rUvx6El
ljBGWms6cj0Pj3TdN/aAUIQXyhijgUfH6jBWginYVrMEjSsJFyP/sr1nrIeOpXlR
7WhzHZVtRND3PyonrIkWS+o+g9oF82SzM9bpgugo8oYnwtJmNl4P5DroSF0co7kD
+1TB2/HcUg5Izls2eovLKP7EmBwRrEQ6JEVCBKATY7DuZqa3PicL00U/laQDoaja
48bjNL2Bu02B3OnoyyttPuUVp3FzeSdCMbW28q0gFnWDWPX7xgSw1Gwt5sEBWmqm
ebBFVK//Mj9pozJxIetO4k7VP8o+XH/SujlFw4iB0nNgpewkLrJRtdnVUQfQXWeH
qDNhJ0/EWsTGZVLV5nyKwLT55Av/lfj8+gQ2dVfbJg5HtrDNGwrMilwaqB2mqV8h
CQMBgIOHltDz9Rwv2b2xHbytSgZ0qFZlWVND0vqEDP3UVlolq3Xu8EDmxAdSR2mX
+/DBs9BaVFI/SCE/lmrIGy4PC6gFnKNFBSwvLs6TY79z65nEZ51m140NzoQWsmSD
RSzzOR0zdYv7ds3gNqOfUwJT19uFBgTiFhCik4h0KqXzPC0wUGOWzDzwORmKNUfF
3Wl3a+tRr/oFpBLlGBy3qz6qW0juwRpCKFZPVTEi7df4DX67ZerRzqCaqFGRc4AP
O/EwJThzFN0s054n3CH6/qiYJG/dvyU7jNinr7qDtBaRyT4k6o/nW86sCitwqOI+
wsRK4oTP0g0AET4ULxApkE7+wD/C2AhTU+L35FqGc77OTyKjxpD0qO74tiIYuZ5e
UexEEK7sd0FPwk7KPUbSrIfQGhXHJvcFh6OwlBwT8nzc4zjYwFbGorOXncgfoRaf
U3r2SB1fVHGyT1kC9ouUW42ePQaa6PWNxqgHTaeOLYIdl/Acl03/z+hM90su3FVh
dgR9EpK6EHNolGqCjkPwnghHLLxHGf4zjyNE/+Xf4xQIlNVXZYTGKhiHa6fJWcXK
BwCHpgi0TXcAKDfQDJCO0xVRtYA9PmOYwDa7QOLeCeXjC6L2WnGmlYpORL9WAAeO
BPtqSoF0zvI+NqAirj4sNuamKIw4w2fT0C1Me06adPvFbd6Nsr2MBJaKlb/79Cb2
zqLKy1KmbQbF+aIvm+8dAXJfN9LCejrUbKxcTBh2Jmg2rdUkSeMFxviwJKROLrPP
JAiu0qlkejVqbT1IH/SD2UmGf+qDFsiqrAmln4rKTIdOFYy565T+4/0d6fHGb29l
23+yaKbeDw8TE+q8H/kT6DAD+ZrIDA0j/xZbqkdRXiPikhJkDB0AmO8utIW1it+f
yuNmErImlEk0xZ9SEo9iRC/brHPxxYOqYYAXGPhXBGAa1AfYVOSlHx9vLcMOPHPH
5ntGEf/l4pBvlFLvVKqteFI5gQIHoEhdhWFg+ZiAUvfccBrSI0maWRSTCmnmagS/
hI+M2ROLKtW+KQqST3oGDuAXNpOiS8QnEg4Kg6EQNgYRucZiOXlbWZ4m3AC0VJ3g
oN0gqeCRwGlQQAequ+W/AwwEAc0OwCSV9Z8Fn4c4fAVaOH98sRazE+ITkYhi9K7t
yYVabVo37sZrVV8w8eLxXP/06Ys3HT1DNh4wRzV1DnoyHFbK2iQwgJWyJAHkLwM5
BJWMk3EJeHodZtoCUln4RcQHs/Kci9HW8AXSHB7+SDQdz+UTJe9HjYHhjPcmqDvt
dCTZw1WyuwfFcZO1fCaElQdb+bHMOFniLVFRjmFHmOAvhLj5hoIPae6+tnu4Y4lL
tSaZiaGUR7AQCsfKEcSoWEF5XvoLpbyrEVd/MM1WofZ5afeH+3ZDyZS8djgy/NOh
285novEkgLQszu+V6YF9X+R+N+UgZj7Yhzb+69epwmOmNpAJE07/atjM3PF/SQGG
f1rBmFdfmgpn6hMVz1YxZ4MNnHBwWINsS/5F26LNoyI/46mswCoPQXidqXmK/00u
XiftYfiK01OPwxfjEJLV/ixAc6yyUP+5fpMmqtz+lMLYTHZpdhoSrCIxHs6nt7uS
K4Mah1leUk62HrPoz/90+ewA4yXSNUdQSZBQQtsuEeJrtfDDKCNn4N184jQgwu4G
FGgp+6pU0g2GwTYQ3TfJp/Q+t0YfJDmImhja4Bo7lY7Xnj4Z2s67CHrgN60fnFMw
Sp3q/Pl7E92ifcIWPWSyCLBGgNg0bj5it9nQM9IzozxiDgqvG1qRXRk35rh9EkL1
OLL0HOAWQmpRlP0uWSYd3I7rveEl/NOztp1D0a4xigj/2451dVH3dQRYpvJ22ZYB
5haFVIij+HMzIsLsw0AIIXhF/9xiZguTQ2N1/MM1+p374xo9NYC/jxo8axV+nb8F
rCqtF84bMZPQKubZMOq1GnR1aympatUxzUsdVFF25Q29uNgYtT9DKQ/+zSX0P0m8
ep+jlKZfk/K/EEpRLewPCjxBP/KeGfpFINg2mFyfe7vBSMmn/59af4X6sfni5yRH
2sY3Zrppj6UmGOCERjUTWW0ckLzO3CY8bqhuCafKFT/8BFlnhzT0dIlxY9+l2TGc
ranhRXk8nXOy/xxBMUHKYQsqMdNHXTxnYX9nyRncgqXE9J1Kjf9D2QP61JA1cYmm
dTG9ztAOcdrWy8j88iAwopIgptIukS7knNMhfk9nXueONqyrhrVOkn/K9TNKz2eu
54d9FfTIhT66co84g3P//XZrMop1qOdPcKF+hcsTSDPA0f4/jNg2GKEZcB5yRU0o
R6RCX53aamjy6+qGghEtbbGMzlhlRfVTXyTHoyk5ob3f4u+zZLwVwRsdFSNyGO2C
ddBjuxKQSs70rXOPsVb94RcUmjK1OmD8t4gANmKa32PaAPjaRrA0t+AyrlHwnlGU
eybbdKCz2CCCHjNDA/8qt4X0TNEn0cfelUWoQL6hbwsmSmMA9lyFQIQXIwhfJm5t
Fq5OFh/yLHnMuSG0Tua/+6vMbiWqdwGACgNm7XLAAq89oy81MNMb4b9nQqNpMx5f
0Orp8C5ORspSnxWtS/TfaqHbDmwrMlnN4tM45C9foHFuVX5A77UFLwiLnZPYZ8zf
3jtRdrmO1bGQ/SRx5lXaGTIN4b6NRtRx3H702sOEZIvskQTx6tnvMDOCMg6CGkgL
HkpUIL83294r3TOS1pbyCSwd82XW3BKt+fIKzEMUoCdE1PDSiDbyvku4gUVhB02f
jM8gCYzZCCH6NSthAeHnqf6GWIUVvaYApItIvvPX7eQixYnl0JcehOsqFkVQK9ap
bas9ZqFO2zJlyAVL2K6b02sRgjnPN0fEYImQ2qvKjup8ntiTrot+3U+YV9GouRaX
rb/99O+okwmVsUh4NcuDsyV99j/5AQauYVnpQO96sCLj8XG1PPlJjILkFsZJDDdD
ISOjYhs4oshOsVnJOCTSWs3K4AqNRzZZ6iqHLMQw12s1j7bg2enfK3CyLdqPhr5W
Tz0HzWz2Wx0AQaPP92XJl1cQxxXzzUFATarbps8oVJ3PZ72xbXJT1anxTwueWgwE
wFYJe6HSY6SBbRsJidGl7xwuwF3jeDP6HPsf1QuJ7Wb3h+NZDU/KiP+Oz/phzOlW
WEwOe+jYVHyc2ck+PrlUw0hM4qQISwLZUpdShvLrN2d77ERomMIHXfQSu4ONechQ
wAoAseUMwWhJTBqz7bIMJvbR2Ibh4ftsCXz1Y2AAn2Ws9+FfSVD+dtJkwCNUXVBe
IGSlnPn4e7QBGSiIbC+uPmdqPIm0RY5Jg79ezFHNH6Jcwn9X+fFTP2AcHE6d1PD1
PAu0GPqZuwemNh8pRAS5qknVpHEFjicP5IVcvanEpi8bjPWFc1rqhbdhjPVe2VJg
mOR4bIQHucU5ZF9kKUXuM2Z//wQ0WOkSELfVycNPYJJ+amIAEtw9xcSQRfjn7j+5
aQfjylMFHCHW9Nt8jTeSWvS/RlOfkIFW3TCVE0ct8lYNFEV2ygABNvgb4JuI6P85
frtdbMwIgeGRG+8GlaiAmRfvSes9MeS2XqS+tGjByttPTSuz/MHV60Qdse0Flcsr
eRFIeQ/M2CPQ0SQYmzDcCBlZpqp36DnghHtZKOGx59cNeOAXQjqtY6PabMrJ3lBq
iCABup/Lkb+ANbQeHT/1JCUhmuupq9z8ab7p4YJwLpAoMz4waSbSWVmnCGvkIaOZ
N0SBqQ8JryONTKdIB3c5cJ3r/56TZe4LttG1YUqq8Cx2ccmo+LJRB9WXgmiOf7UX
y52p395MTCQwcKPyM0Q8EpN2biEhtCwQvVzFF5NlEDi/TOgAsQ2fgYBvaZUunIKT
KSTeCqq408DASQ3J4ik16URre9OpCrSHyKeKtnMnuerQ9JHgVED3YzGhk/GbNnK2
JUlaXmMVTOzxZMxRdRwRV72tkYd2Y0W5oEHtBDeq5Dcdcs2zSdw47p4p27VfTh46
aijaT8yDf6lJCPfQ7m7RrsuOJKl2p57gh7Io+KdMiX1T2jERqbiU+DgC2DSbftV8
bfrk5AVAnHUB1FA9oIM2ugzPIrwuZsH0ssJpQqUCbBYa/IvQiepf1gtpgBsQTPxa
VOqaWFR/ULMeQJylX7EjaQ57wEc4YHCLRyavRv9miuSigY4DsMIRTQUDB1smwCji
AlGz2dLEDPeJ7bdasSudwi53j7O2Z24+64Hl+BrrVHcost95O5L2UvAgb7U+/dGv
89Sdm0h/C6kD2pxyal5JtlgdYurbiCO6axOYU7Xjgp6zdalyAzxABUOszsfjCMvP
QSPgtvrhjQTBcvog8SlryO2nspIvhX0p0upMPplZRI4wFEwfhr+5nJW8nvPTq5hk
cowFnqeRe+j8O1eqWexa50ZCt135j2eKtxy1A5kUmvmmgMFB/NWGXdaWlDuaQTD8
3Ka9LzzgbsrwdT1deD3N+vPRAr/83KpvMDdev15N3HIsERmO0VdzhTYfDXDfQCeC
LaJBfDyEArL7mdYeYwKu1chArsNTNJ5Uy9E+jBUITWDvyOvB6xA1CoO/97bvHcGA
UU+FUopJF/zIAa9IPpRWWobrnNE91GoGd5w3OAh6zIK+yN9ojBooUjQ2oILqaeBS
NhfI35F0D8ydapRbyJYx2bZwQ3zmW35hms9nrwIBejdruuWsOKKHxF9LMDmhreya
/ZjboYwqJtEkVbnlYYJgszk7RQItkzcoWZRUfQ95+US4swPkBknZMG8nvYIHsbMA
jjDqRyw/z058ko1zO2fHvrxxhZBtlmSqfzGHphvgLtWxg+OHr3h0yhnfB2/TdzTH
GSA5BKDPrNVXKExwFCUXy5T+A7JIVK3t1Rq7kO4Ld4/XbztnFZZ8dR6BEaSeb/cz
g6z0+S1gQdikKnK6S3lw94XF+eX/KsX/hLmf6qrRqJbwOsi3e3clCYEHjhYTMV1y
Eh57op+yPp78L1kQJu9M0kXNAWbJeumozWxPNHaGTERtWFQ7YYa4BaWXKRJbdqiK
YJ1aLa+hN5N74+p8AtHGCzpSVpOfIHyLUs8E7E9PJBl5dLLe4SUQqLRrgr3zGbhl
9o53sKWAhK59SkTZi95pJSt6U8w0a4J5CtaR0kqgLJrgjLQAPUqjpN6UoPmgLQC1
qn7o3MjSEx+tGln/kkm7GX0KrcZukDBIdgby3hDgDUsDb3lbw+wqoZzZ2MJbZcgA
nGqepvpaVBB8OAQG+eUrc7teyNH9Iybz28dp23PX0qRvh3azBUFwCISYmDwN4ZPF
kRTNBr6JSIc3FKpjY78kIqs5M0bbOITwUt7hTnF+qtui62dAlKo8h3t/x9JF5puf
/O8EGbP4bJotFLIF6vNqb6xOVxNg8BdBslLqVh91nomNUQ9R2BvJcrjLqP45DTlm
9iZZuDiCZ6oHXmdPIBDVNDKc8dtam3upxN/scw8XHNOiG8NDXT0LkAnUMOpWgxxn
aXirXPB1mPh73JAgnjm8dx1uop5kOj+hm7MCiPNBJXTA2Q9LkWvF0/UXIpMv2y2l
DVwCnQHFli/hMkyNl2EOObQE2EJKFEK2/3kDdPaShcIu68L79sN43MysJFfz/OTQ
t7/GVjrDqz/9zNy26lczgmtjeGDPTBF0vR3BjpNpbdSgQy9yHui1vlDoz+059Mb7
btKo2VFrFB/IvS2Pa8jVcPZXL/Sv4Df3PxwG+JRpzoBjhmEZdozzHky1/LAMi6UZ
4jjOxZW1FsopDT8X2d6gzRDfW073hFTCEMLYywijsO0FKuWpLusjW3FyKjz+ScFv
zHSd1Emedd++Ah7wkXiGFdINBewQtJiGzlFTlsQvsjx/HcmD4dEwqKrvRi4Tfdae
/+9sGOPD5n1G2GzsLMwK61oaEjBqOAEPLzkycu5qKYvfePL5dnkNeVxKuhck3AN3
0z5of3AGkv736GIslczJsQfMCzXDq3v/iCkyhY/jUSTBIAj0Dv+Ggt+5odmtrDDF
yo+pk0I47G8ZMt5LnX7WoCZ35INHxNhX0ZH8k44Eu1ndwWv/zT1M9N3vjz7a3Z/u
FP025nEQ1AzBbMFbIajWMmKqra3IRx+co42+s79rZNiwQ8bO+2eEBPKYr+CH1+tY
/bf0yKpOi0A6OmzXZPK3V3UMnJtq6kwbESq77/YhTG08cD3KRPekwN/cKEuECyB8
RGUvWUDqXGppI3cQCln5fLxe7UDuRyiIQaKQ2EJr5zx0rofC+zlyRtHGzJESKDdC
/uD+IToMgxkOsh/Kaid9a4g0Bjxno2c14LE5R7/TVUbAgKsRu9WLCc3uRtSZM29N
A0bFIjs97aEGwwRLN2uZMl6mfTQL1WodMEJ3bjuhjI+x3D3a5lTuyIQZ+KWDncs/
SCGYRCP2YO7utwiX5ozDB35g4iskljkWodKT/slpQtDd0t6chLuCwoOr+WKzU4w3
F3EJLl2b9yVQcbkCwRMC0PLaB0LOv89/v8AeS+krOGbuImp238Mtz/V5O4+87n+2
KB/sbXXVgIDmmYeRJ2nFEOnWOneniulrr5LgVAAvsSHuw2kdkqQpOS3tgKqmKdU4
YxuRRBQpUkaEzM+wg6Y/bXQ330Ue58KU30nzSOMhzQza/q0PkMFfTBxveLcyXMzF
4aqXWWfLSuSBXOdTrxHXxhBPSlvMiPn+oqmrpPj5IvAfjmFndmzE4mKQMCIlBCAo
Vr+xDiUb09cJrWsndBOhunM7Ad8eOoKQhqlK9/oEDTGyWV0bsf7aXFdnCBvIXMv0
pdYRHdS/Se9Y8Xv8uqS/rNAI8FciytZqpTTBPzdA4t+EvWjKT+klroTMpeKi3nEF
b1Xhwfm+Y0eJX04Wn9XX5ecuVxMNrBnrDe2XthlDLN+Xnx99241LOjkXaaaAdM5K
LY7fIxfwJhJt6DoOkuR3EIzq+T40IGbm9CyGjc6ZNpTgyFDG+EeWESF2+VGm6Rpe
ka8Rk+sHUBOOy1gV54M4zdpOVHR0oJYgH7Ae+3739HJb/8bGmGVU28zxYJpxEtWI
/1Bw88bBkXsXii2svGIOptMnErlFvAyj/zsng1BRrPj2BBRuzy/SiuyYSkDHLDo2
znJuNMSLOKe7/XjWxMTOKT0EWNNJDV08XogqHflCa7gWl50jyT/0tMHpZMeDRPkj
LvHbXb2OHVy5n0cQVOummUt52ScbIWtBQ0qsOXZg+zYOmoX9RoyYHKvqnv+vqkjK
xBwmaIjnEghHjOh9ToTX+h+rxUl+QATc0BIQPeUxdPNuImUaDg/10isy5eOS76ZD
ESXiA8c1vbyr+r7FE43iS7Hz4vcp7EbIEUHDs5UEQ5/POizKADeJVUtQ3KxiEeAN
eTvwSbUQzfbIJETm7M/VIP91RizGv2yOV7V7HzR58FNhee4OCmqg/FAYvKrwmwCT
xcPLStl6SL+dVOK7px4bpUF13oqW/ThBPoryzVVDD+sl4lsuB4YopNWFUr3RKjvg
Pn+FokvS9apf79pa5zUi2Om2x1n97g7+HHtJPjKJZnNtU0j/+ltZ0UVySq3gPejV
jRSUD8uWYMDAoxq5sVTxT3FZpyldVuEXF8+giAUotY5vKXWR/bQSGY4kgYYXw15O
5ErbC5lYOv/8ZXkHOsy59O/+CRCBHtm8VYLr9RZ0xiD7YsXfrarq6iegj/x/U6HX
3fy1S/IJsfYoBf8s3NtZJxUe95PL0APYu+mlv0UM29wnNX/zarrfKFRJf6+BeX5F
4X0KuNZ9djaYhFMyXq0HqOOwz3v0o9KujIyfqjJ2Nj+uDklHBOvi2pB9JFRr/PuW
J9qZ//QYCG0p+5N5mliJcL6ZYk4gTStSVLWsvhAJCrG5vSt2nGQUa2rQhsHHwRuK
Q+v86PFJ5/qlWMZ74TSKvGMQJF5Kq0iKY3R3XJEgiYMAbi3tQrR+RKua1+42Zyoq
JxuDBS87JTvyeQSk/eOkeWczXbk7eltciAb8C3fJVnv0QOuY8/nZ5+JQwyVeL5cr
NkUYsTlh8gzYuQ1iTdXC2z91R1nI3mZE+9Euza7SFmByThzgMyhjFiv4SNrXp9vw
UM0lyZt4B4MCGV7xgnFUkyA0wjv+iJQg+ICmDCIekf4TnoeInX6mhMlGPDfN+b9l
NXqJGUSsb8dr3jvdSbaFkAmuFr+QFRjxS+xx3TzeQ+tN150Qa5gWoeBpdPfgzft0
hGRRV8/xOPUaWpv5wq+2wHbq/ZtGHB64u//eyVb2fHt7xvH/wnQVQLYHGJDFUy+C
0ReZqKSaES+Qcd8gyA3hrRv33KDHd3wVAA1jd2z6SxdRZcGmwNFwgUedXLrno5zk
hGNPJgH1kSlCt+WzlchuFVPD3V1FzkbgQo+SqGTm/1peHJ1YTWXbnmxxpRF8nGIX
Lwx3zJFQI/PUIuJL87Gg2L0cnSKvYS1rbQ2nBuqpwQy2iNZifo6fklkGvhHqS+0P
vdVpXeW+8x0wfpyeA0ccAwFfu1i/1Bl5TBM9E1QhQ192UUTdoGT4m5vMnIaxtzgR
soNmUNMVV5F7ucxJFHAO+kLVwKzEbRK3JDTDOai+WraJfPi/0QKMjQwqNWuqz3On
dIhx92JNMCOa1o3qL2WxyA5xfLikajoQm5CBXT51n3YWhKZk+lV9VpvBgzyk0I1G
n56HnmIBV7aALM8B+43EQkLxZX/76l+Jfi3T9UGHvfshzDj/rGWjKfaFRKqwnXbi
d9CJhvnEg+RcMmVkFK43lEMmSExXblSKaey3MrFXkQrzTyReE2p5IZ4MSMWicrLP
sLNMhohlUYhfqTIBDbvQYBbBLkhBi9hazxceD5BfXwJxTaguWCQd1/RfFmpT4C5+
lAN1vUYW9mjPKDMPWkZ8rrDF7WZXYWvVK5g6XBjSekZiPOTyWZXM//2wpfUyY+yF
QvYMsQhugYwa++YUIJh/I/4wfA8pr5X5tq5UFam7+Kzc0qjVLz0fbuAR2blVyT85
RV7nZS1KjKYFQ2UgGSncknhSUQ5CuNPwxPjw9gEYWQ+qd0GVRpT/Qu7waSzdIHlx
SEVyX7DN1BEJ3Bv4znaQ+Jgta9LDvP+szHxWazoJ1eHgiWTttZbHqgnSqGKVs/D7
Ws1GPP4XyazFV4D7cCN8VmoqGrlbjU+qs6npC7arQJm5+I+Q3AhqD3zwby7LWH7X
oP4ytSUzNvpd2eclJq7auP4XyZqocH6TENisGGSwrkunYqYtSTUs6YxL6CQaiOzc
oKscwyeiK3BHwLxpMaNtDozL/ypa1S6HgmCUPU4J0fegVQdjLSUKtHS3QhMFkfpA
SEtfLjvjkEVVPDIaJKPzhqA+pXKLln8kKZCSNxi+BETopMPB2TOA1ou6VnwDx92c
K/oZcP0XpP5ZD5+dkZ2Nj5+VQYAnYGdSkbfKx7d7uIBMlNR1Xe5l+oISZMFZNINX
JUPFQF/sMboNuAcUhufDJ8kB05TbYvhyeR+tK3wexc5tmX+rGHMk1/GV8rw1Nv/n
eruq9UQUqNJ+nScSmaASDvZxc0C10azpYqSRlMBqbLUrAc7wZgpcRtKKjNs1pHWa
4PuAFn62tyPUEH0f7Nbe2aUSUvI23G9WCetCqplPvj7z0/cCW9nHZSMTl1rvAXut
iXzqeXmgMPvgeZHomAThNasX8iNRSxUcWkWVsCsfA3MsLyQG2Tj5/+X4DdgpHuMG
f62tfucD1neE8aC/w2BfCCKi0BN1JOXiiE7CSjXajAgTdnL5RkMyTu7nw4IoaRVC
64bXnT0rP2a/SWJlJK2Bl8md0BK1GbIAkEE1C3rmqFwVrZIwDGyPu01XHKUJvnXq
Wi3XKFGF8gxKfzcBewECNOwuq3Mpdz1WERCvuCBQxzcCg71g/rjH79JFOI2T9PIA
JzAYEZbrl+qXE9Qc3wR8qPEQqwCBE3YR6OUq75iIwj1FqgPEC/x9+5bkRVE+nY6s
z7ppu5jgkdgBqnSk5ldVnRSwqC2Fifi9a0k0NSbtHX7fxbTIl9nqzhSmsBFvo/XI
jg1JBjp3M8zqqK1BksiCUXNi+MQcp67xpfHriAw/qSOiA5Rvbuobx6829wSuOjSr
UEsGqQItfsyqpUbvl7T4AVeHZ6JM+6P74uuH6IIojNBtasw5x+305newUlDhA6wd
E2bQwgsCPIs2dzShLMdCxsHjVCXFJPlx7V0nZ9vRrO4NaloUL0YPg5qsYibNuRwk
gYKeajvSksWxMABljJEYcLQwLHppWbkNF1RVXbV3qq1axZnmLDeqb2oemP9mj/Ku
nooMPP2dB55gl51Li3rpEgw4JSWzMceBScGO/MJN/XpZRbYev6iFe0gPRMB/Cegu
ZfUjFq6BxBXFpnhoM0yee3B9LLQWeGdjkkfq6KZog+3ymsaxiyoo6PIhc3v/jtHQ
oEh2KbxCmJOWGFpSO4rn3aIVUzU0ilYDCanMo51m1uJEaoHWH+Xzd9rWDTsqw6B+
unZYvFLG53iDH7jBAYvXDza3zrJuA/IwFmG7U+zh/xKXcBsLE6CK9WOEF1+ZIBVW
8fafKFG5da/bRyVVKNTkASDOVXyUxV9R9ZKaJNh4AV7d8uJEV3X9bFsZ1R25+Kf5
vcG7b1EdsCuVwroOwM6B2KStVuenfhI5lVI0T/MW+HojhI6RBA74y3lGdMev4fir
FGrNvCYOqkLJjb+QATcLgteiDtUYPmfyVltUmj/Yxg/qgNoeCEDzXvFcsWavgrmO
43LwojFmm25lHmhKpfduC5R7dz67oZvCwuwkD91SgHV7M3QGjuYdCCHrH10+gFd+
y7m3bbjvq7dmhMzIX9ddL6NXG+jghdShhQePpPbcopvdzgPDFqBuTkeu6y+7oZVP
BqxZDrGH0q2rTeh80MqdbjHYy9+XbwliC2Mc3uMP+JfiRiwZGRR0A4CxTYeWpgvk
j7iRvY7/v7OVq0PmT37Lhtkf1j6B1eibex9ibhYxezoPd5u1ub27VC6UUZ1LMzuP
WFI5wfrIAZWi71noPeuEHTG6rWeJ73TOGB5C6wGP1e+oeLSQsYel1CEwz2oNu820
Z8LIYYTsptI0ssInKSp048zR96HOLQF/fTEmR7+2+8q0kuBTnk6oIjZTVSD/Dx/d
auDh6Y6aTcEvAF9x5pcGJxeah8ez87dbOgh6IMV1ODNR47f+n8HGzXobRCpTCNlH
LmAqvnIw6i0fw5MCyQKHU1RVruoi9n4OWScHihxUjDQaJEcWDMIDHgfAc1husUod
sszAnVCkNAf0DC/VvKMOursyhcDsVSJYxWRJmEZa7H5vLujqkx6jxfJv1rpjWOiw
wIjyn/Xp0WEBFamfTKgrM4vwlza+sR153ChkRVTdaESxyAOUhC/5P0P0XfWmUm8+
AeTV9T+GQvzaL+N9PW8U/9eoeulTwziXSBxm3vluMEol35gjEGNzS5Q1p5tLna3S
yaf8qA2lQ4qDtwK72B6QImSim7PBgYFhgCE4Bivd3GeP0VQLZ8R9M1Hs+AdLh6dD
Sifa7aLG0L/9hSwvjhEPQoPv/5+3pUNMgK43YwyHz3fy/wHw5drZ605arVY+icEA
YNFMrikidTeoTsbelaybd9bSmGYkoUzypYCsBOLqpFvLL/mHIwl9mii6xquBULKh
pt/6tGZaA2nX1W7hyHnr16VDc2MQrZIJGNtGJD+WppaaCa64ZFLjifDZhvDI1FGF
h06t/9rEZj0N/ifiZpPUaG8v79Oe1n1bMzFCmA4WawgSFfTi3kVXQ1Vk9VBwLT6g
EZhsmipsSnPSJJL3clm4yyM6s6mFZHOKYW6cYkm+J8kPQKe3qfkxjJvPDYL+BxVF
kYun/NuGcU2MUnvM+7Y/DYiGGyZK/DAtD3QUntCsgv/XsyuaUDi0uz5fCp3ezzPL
IF+CrbdTixvLjWY7CLm5sCfMsdiazDeumHtRKUbAcrE4euJBWgoIV54hcXE8VifR
rUxgEFvpHHqEZmoT+yZ566FuWqinRu2YxxMwvf4KNJYJmFHWCAuL6vbKb/i4YH80
vWRaxuQAy/JvdTsq3sjINMkyqRIVqQp9RED5qrMnXyDw2+maNOvk03AdHNApDcMM
4c1XN08L9L1UPhAERPDHDEINKVZ8YEHwJHbZ+J2Ddk6Bz6ZifPsnPzYTEDImCOoE
++tXCbK8BCfwmfq75AbNQlMVH+uH8IQpASupiZTxGEiKE0fYf65J97cv5MLfnlMb
9bvaF1JIlRQm6HxEANmn5dudSkJmxeHmf5u6VobUEvgl4gWG0w5ri5KWLZ88mY5g
sMYnmCDjOrRYXw4ctWJXIXkeu4+v7un0ENABMtEtrFRZV5fsQZeu+ZfbcmwGLk2n
4sMbNuE8vG445EO+ojfYTHkg2iHNT45K2OAmKcoij4aOFoYgwDleDnkhuncfNgkh
+RtPpzF1k8TOvi8V4rrZPdeuR/AkQUzdf9Sfi9s43cAtbe4VvuP6dqYk2GgdlP2f
gBDPSAIigpmSRpEjJ3zuGzav9hvsOQs8p9ocnv50nRebKw6C/tj7wjYrbjBe9WP3
JkAVMVcC7wDtwAxwBf7NhmXZRTDVFNnP5btDA7AVb5VDMiQtwLLfQM90jt6kIk34
3s08jO62/KJsGJHgZhLPmGAVtjxNfie1bKsMv+yZDwLZRh1xr+h3YOpwqB5NQZKG
2P+OiqTrlW+qHHkLxBtouay6HDIRE9DC8Pp44ifSvfU0Np65nRW/xEaWood0zf7o
l77eiEhuSLZv5V8kyT7Z00+G6wordBlPn0bBVIjOvaqVouHpepF7JSxajXfueTmq
+lKjyB7dOydbGdubsUhMN8EFjnpX6IbgqNrW+qexKbNZX99JvhprvdZ5vZUB2mHT
YAxF6rh5qstdVdXAyf2KKVyPNKifPltFbeqAQNTVXzsMQphvAUDF2I4B6fVNmpN+
KbaqqzqxxwqhKoWsKhFzBd8vWTxdfGOzxmBJyPGTi25c+32C1GvLeJLOL8M+ABN+
yMHYleFeKi3XpSQ5I9rMRgDAUv0U7nbb3StR2VzdtEc2R/LREHJ7TsdHDcgqBRIT
79V8irOeSKcyqJ/sh1hpb0R5RWSEznE6L42549oaA3KBRlQe/0F2Tl0g5CPlfQ/t
Wu0WaIljxlAe36RO8YwnuClIT7g1tgs9XJM/RHULezGpAmDGZERfihutYbnSfTtj
AwM4Zvj/Ggo8uVLFMVwAPL9V9o1slojoh1qUio+XSIhWLUkDsO0BGkBcXPtrduWQ
atkwmKEkvWRh+1aqhIl4jqmDC35vGMkrawfiWo8YY045+6AbvV8xGHYgDXYwEBym
/jc/IkbS/aTQbcxKfOD3sx101tKADBxjhlYlsiZmFPgwk23OLWW6uNRWkibluN5C
28KAn8Mj+1ODsl4Gu+FuhCPoYK+z4LNbvaLEuTb1klkEN31ooQ/iFIBAbBq5+SAn
ylSMvK6lp6m6nvJlnbDNNJ83huYAzJivAxQQzQX8UL3OCMoa37rR1aW391D/jW6Y
5hrWkNUO4SV618k0M3KjofacVYbyHHdouwH3xACR30GlDk0A3lvGk+6Nfe2PGa3Y
kZaIPaYZDRYG8y/1xzwKc3JZZ/z9mtvqmjNWtHpa5iTNDotbOAS4kRTb2DCKJzQI
RuyZamSe42nNEUNFQJlZkJKqZuCE0axQmMS5pNXV+dkGjlOrjd34zJOyIa+yMVxE
vRfeEn/hMtzr5C2vWT8hUcgeN+P66W+UaMH0tAlSGU9DYf2B7XmhhIknUMdKkdxl
CHWjM+IbgyEqNjK5tW1rBXZQC2ea4uyTyPg6tSjXN6cCgexY+KIY8rW0jtArlEYj
pOvIckeoBuh21K/4L6nzG7gwRBUFm5l19YLIsd+hml8Q2PnOiBmDrH48j3FnlmBt
8ifVD5Ix15BCxS3qumfLzY0aU9S6688tU+/2jM/H2As2kHjylLqlSfsVnMII4SgG
FFlgFPAKILS92S5YNIQdhPnoiWrGdBi/aB0Pd4Vjx8mNZkIUl66OMd28+9w9TH8D
2XOVeXqLSP/FT+lavc+jEbLbhJ801Smpi2WevSXnUIbRX08aGg9YzjhKUs/o7eEY
SN/BV3VZBo/DPJhcFPG1TOGkOelXsHDkznaXeZt9eY0d2CtWKJ/KXGnyuhXcF7sf
LJGOEP8RKJQN7AT4vRtQtpfMRmDd6wvQk9xDCrs+mHx3LLscDB+Q8yci1PizKbw2
BAMZOKCORsQJNNzq0OPBGcawHHus3kfWsexBEDLHtaUq0xiCs/4AMrOWh1HDfcRz
U6frMH5TkBtWfd9W/8p6mKUo1vjoq4H195K/7kLoLBvmp/agWloDrBJOv5a1NRJO
zfMaUcR9NGp9NTVD01+8E70ief132wFGz+QUN+6ZEzkugX8Me/WS1ADej8J2y322
0YYj0sOH/yy4+kFkjlaFY2lI6lK5n8w0ryNf2uC6EpASVEeYS1wX4IKKmIGYD7Un
vMxztGPH2+4U7pRX4ra+IIdDwLpQItBBTNlmZwEsTM9lxnQRGmV4vU9tni39EcNi
MZS6Fzu0+TJEm3I7gEWBEe0bKbSPnRZcQq55OICocU+2DdRwO6svIPRbx6OyYIBj
iKP6lDa5u4fjRtiTQHvCGeHO2PbpBEOGBzcAJyuiQVruta/s69XrqtGjN9C4LSuZ
dBSYeLYSlNwJllyZ8oFB6x5NlhyL1DSb04opyOXvm//B9AhcpV3WleRKx4nCQ37x
Y4tq+Xy1ZxRYKkOcAZbpSzpr3LEgWfHNkm9sF5SLzMsH8LB4OMq0QU5PED+C13r5
V5cBj/XroNVdYkGnzLaDvG78pskX7ef+aDCfAAHIbPjyF1BS5YOyfV0iRrCQlZPa
zdz/r3KYy/NVqnoKrJH9MD1poCiSSmuO8maDCzn6JJ25Z+uMef5/30x+qQ4ogoqf
6s5yElWQGJd25cZnHWWz0nCLbiIrAVfPjhAWQPnGf5C6cLIeBHTFMe0aqjdphxYC
1NY5veJT3GLC4iu0jN6HH6Lxrd5X06KO7Jhn6cC9XnjhQFGQgfhAiqlxGhEN0kOK
u6byfCC72qa4TRvQcSEQczDBadHlKdRsgwRh5eR1rjJbcHT0gXz34qojjg/AqAEW
9q+pbsfWJB91GRY6sm4fxC5IEQy4jK1P2Jr8hkZSgU43clnELi2P1GdWlnwRFa1s
QiPLyTsRMTVHcd3c8A7/5idYaN+JO/djwg6A8khd/M9iO9h3PXdQ58hduOi+0gX5
hpA9S96upIuF1eQs3ZcBcv/qplNz4Edi245pXRc2PJWFBEWo5PPG3Czpp+N3vArA
Um0bbKBLOE+gbLJ8yk8ASVYR34GHE8KEOo2iq1if11FjRUMtIGDpbFPyLMpTD2lh
YqW1x5YQNvHxVORRC2tovGoHHw7oDwlNHo959SPPG9EpXQch/KwCnCApkuxqTN3N
Mmh2bW7DGs91a8/0k39hXKS7/74a+8weQDj8VMfMi5g0TGhUroQPGO2FKlgdpcws
z3UvCs8rzNxbzje/PmfYLkdVUHVcy22nG7vqyLenRcEQSu9QHfI53YBeaq0vLckq
0ggrMotEU0obDPEHNIG4o0R9UowMku66IacdQA2sVQeQC/1edUKjoSFTq2joQp7l
sIvLA82J2+J9uSGzuwyy8CXrw7FqM6CD9lSlET4nT9e7a6HYXbYQfP4TOH5qchD6
aJ9j4QxB2qGnNrEmtP7mfh7vsjsxSaqJYVIrkZAwZrG6ZJ5u6sTT/iNbZdXa6kcn
CQ/liCk06eOsrwH7ma7q4WmhKLq0b7UfUSazIQQaJxOfsJY5v9s4yZgf6eESaCqB
FuGPHdUJ4P2RkT+ge4ZA4nOy7ouWrlzrGWXczYnYgOx2gofMEd2TRgjOl538dF6L
oEUJaojwCwG4Sf8vWAU5TLCmaKFrdNINtIDZVQrwuqDTqbtGVvtAE98GJ7H4MhPb
tKbGTsNRErb9I0CPJ5jhn/uY9uDXae1wZVyTQCT9CAFk0F5VJ7g2fU5avzMrGBGD
eQUm1oVait1wX5uo+yHCRwN9DWhvmq+G35OhaKm1UqR50txitAxfsCud5wd4EDnz
zAB+pHpCPF7eTaFXMEaHb4l37M9CcupTN+pvSZp8NgD68wq3qhR73h5hCem6V9zk
IoBRWr7GP4Oobdp3HSQkc3RFyWIgV/xChtyBoGPicHdIoBrKKbG+lX9b5OLKHw9v
iLSeER1pCdFMna4p6e0G/6BPCr3fDsUNzcOS+NV/iwGcj8G0FU9hCm7HLE5/d+78
H7p5TKGAJt2Je6i2dP2VXKbR3dt9hXM1QUaSiYDP0DRn/dX9G0mzZR3uX1vP7oLC
PSOh69Ks1y2GencLUOjcj1dokvlYhoWPxEe/J12vCn7HiYY+O/MhXH6GgfokBTJ7
cWKrfTNus0PovFQEG9qBzz9VxiMyFRsqoWjDPEcImdyKcjuJtiaLFntAruPY3ugO
HjnwVeVO0qofeRbnJESvJBGm4y9aVJ+b2SbDNvrRRuhOT6c675EMHrpH4bkaRmpF
nKMEMOyigUHc5xJWhl7Sqopdv2f2PaMpSjEBdNgkLQ1KgfhPRHyypxVJ+BDwMn6+
djzLtZJWLBISi9J51AbQ7WKdYc7linhNpkRjfwylTALEXaN5uhjtl/SKb+q3GUnL
Y4J5x1gi82XC9SHF9Y20w5/4ABwhSS02ohkDWnqPWbw/qjr95jJjjMLus9hzCbsv
br3Of9nN7h+Amf8x/tuLtmhLPgFVx8sMvqe12N+ouxKNmuMMcW8zXo5DA1bRP2iM
aaLGVL6hL+UcdFoOekDt80RQfGYwi+y9jKGPB7MfEKVHSx6q+FT2A8BdXzSBZS7N
Nfk3jiqp1YFRrIqx8a5hzuPgQcYkxZzapL4owTnOFX00hV1r6SXzg8er/ZjHdO5j
bauLojD7XnuBb4PLLi8oVp/tRS+saI4cIwQOt6K94+ZulnLr8WGxQyt4GLk6VIcM
deraEjEc9WIlwJHiLMAXdnrF6woQ1vFkRb37fPD7fh/Kw7ik3D7CRngKw5uonyxu
Od+7k1sbXZE4N8qPnhIm5ycKJ+rWhGeOYE4YkGzBaozP/ywGPGZyqBjSsaMrZ/ON
kThcKD1DGPcbUNGnLvH430ZiiIFsZscpTa2UtckRMLC2bo84op6OdtZWT6cuwTQT
aCQ9bAwwDSrQbse8skqqeL2XTgELbxR8cCEz3uHBA09jt8Z1kRCCuJApK5HluFSt
PWN4RI8VLQKlXNLO0WU+dFdv6mxiHI93QnlNebED6GJzmhmxDMrHXuBDfarJzeKL
bykFuF9BWhBMQHKMqGRzVvcLyAaOXAglxdjX0DXxvtF4MeuCST1i8hSp/L6XTNME
m3NHJiGyniKIiZUvP2/GNYaUb0l5P5ypMIU75O9YWuSDj4b8234AdwCtUiMMQzvu
RA/Jd1rstejT/A5AUDVfBxKunzYh6L2oZqjgAXt9geoy487pg6zl6jaoEzIotbcV
jzCiodj3fv9qOpINpaLis41F3JMAxfKr2LA6dz1pEI6+pRn524T0iVihUXEMPWSI
78aHIk1tz9l3Gsvjwc9Ikn7/QagIW1p/P4S7a4x/V9iZu4yo1ryBMFIwkvwOBA8t
1Fcx09TyANJnt2gF/e3C+xgzepJUlMpoWBIuSw566cvDY8iDKy45/6vyNOIDIc3F
u8UruwYnHYq7RhuKyVcl9fOyTnElInvMpya4aOTHT7hYN4jW0KXUP+x6alBwkR5N
AfU7Bbh7pXrIT0w0s0rwKFxrsyHcqA3As8Tk/Y5jkND6ybLCG/5PJogvyFhPvqsK
Qc//1fQVZeWU1JxpjpeHIe0U+4Gl/goK+tJlKOAVyPs3bj9oZo39h7YDKqY3ccKo
VDHP/6KVeRT/kNVVImEiPCT7Cz6Qe61UW/euMrryubEO0WLedwy80tdUoVtjUztP
P2ZbIQFpfptwxo5VvFPZWcUcR6Qs9DGIWFEOBUwOoOybz8y0HXuGkrl7/kL9LJ5o
xQrcudi//lB9q2Ct3pKxFuZ/mFlXsltixKhrndTRUrkz1UG0ezsyfozpHXPEgRVl
IPpcNB9qW7FoV8xjbOKx2LLuuvpSXg2E8FFmc/c1A5iPRmwav9nTWuTojEMVBsfA
5E2g2gLvgKZZ55xpfwgHX+WgtSXzzcUo6uTZmeS8KQaH5/TTlE5FI4XbvwTHQvlr
K7lvnNNtL/8Dq5WO0egepzWirlHqy7LrWxpu6RTwEzRuqk8u8wwQo2o0SUvJqjNH
6l3S6z3O7SfVWxOIvt+/wR/DT3oCL8cp3giuhmz9h/VesXYH4huM+klj5H+XxDKO
L45p4ilsVfYmd7iOxXQt1EALOQPLpbkUmiEgEWt7jrwET0M7yqgJ8Y2X0lettn2x
CZ1nphVukNCon7NqwvwWBNNCfHUe3AZ2OfdOBRoev+MmxwHHsyci6D/stkxr3ukN
ej6McdFtutX10XeZ4dYytUiJ8/Vk2KURvw6XzDgJJovLHHRGlV/fQP10TDcaYTyB
5EY5vEtXFMUPzF3bZE0by9MNSXr76YYOEHpRttk+X5RBzUI4b2MOHHnDgz35wEak
fd9gak9perHyoPG5nR8VLh96tIHSHMJhUljUwOsbBjhBtAPLsyUjTchEb+mDPVKP
2GN+hSDAFx8PhpU+IQgKAprllnNfIQ/fC4Tuc2MvCrpzfSO9QTDhgYnITFH5HbDA
198YFPC/il+owaeuIA9r9MXA/T8r8VTQ5OLXx7PS+sm/JDdHRU/Q1mJKC+Le2Sy5
0Cj17Of3pdufU+VS5RMSclK/uDSPNRnj2FmEi4fCzyMHKovBax5rJJ8HQ6jhz0pH
8nvzo0MHcBbstjNoWqeDZdKP89NYWnnzoe3TIdBRQeFVJDrzFvRbNllANgDdL1iD
oQjjWx/y4O1/6xSFJ8GvldV9ukGa4o+CSf5rom/pUnMUxbS0EfjnlIVcdUGomCHU
hRQlJj9p4wt9cem5JZ/qgd71ev9PT+ow+Yk05mXyyE4RgQE3kE+IXTZ3Ilfsvi2h
MBdvTd9C8/g3ooPxOqLR2JwjnyFIMWRnA74sXy6cLFsfWkA1XUH5E1+5G1m1Sdj0
a9aDjII5D6r6N6SITRCxekqJHfpb1qEzfx5bQ3JkbqfJJjmU+dr5EpNMa8vcMJXT
kx+UqDBZR47tM9PIMletj4wNzmf/hDj0wnhjrInHhqu7lYcgEwPIWof+4tw8hyow
uXqXwtCHGq/i2iH/57u+rAyBgosU5nd21y84jQtdFExjntcO1s8Od0fqoEBCbsVE
CkiipekjEsi7Dg6Do8D9EkDSA3glMF5zwE5MBZtjeOHX+BpRZEdIruzWNhjBjbUo
o8gf1cj5Qv7nGgBnw5FLZhxV7zAtMyfFBPYOdqH5jpV27m3PpPV5PUHmJlezDUT3
Kw+hGNm91b02z0xmqLKIviheYoKo1i//0jqbZIrkqrcB3dyK56sPMQ6yunWjYYc2
eb9uBKShWVV+6NhTP33DyhJ/vQtvKfD30P9uyNYoVp0zwobpgNIIM3zAiN4D79kU
0WjFsM0UjkUUX7/A6Vlezbf0cH1+e/K5JJyBEOM3ZGzG0aCgTZHvwo6uWoQHC1ue
Kg+DZsBRgyHYkUSLrv0Jn5poxl2qwaxLE391rRbEVwlUmqSYSLVwiHUKJQxSnjSa
S66iNLJDPFFM4RDiMhBJwOrN55fCT3P62wkxfH387+fswqDsrJCDoipZ7dWyrruJ
cYt8sOxpHyMYqq1raH+iWocS/d84NKYRF65ROw8o1GEX6DOsqlyUHXxaROSB9EOW
4B9IAV6cmHMRvBfmdZkLKsOkqkND54jzU1oy67Z8DfOmwiueEQr7aDx96/t58VXR
kvE6+4o6UXIM6BNM/kMX+GuqyYeK5AUmLvqXoaBuM+595xyR+h8ajZAVMMcPVnLs
WnyvCA6YSMbnB9580jMiB19bHE2F79hq8pl8aVNzIKKhnLcql397SZguwo6gD4i0
xVGl1EI8iDRmrP1lulZCOfKvOEC5kgGBKntHxvYCO1fXBoPNkcfRxQHCNmQqK5Gv
YLSB4wxoTyhCJdaVC3qs9SP1OstYS9PmlSWdkYnnEY7922dREy0XkmgN9H7GrgaC
k7XkPQNEIuYMbdXem2yV+VJr1Qgd1xVolh1KED2oVJKfM4S3oX2xieY2r4GSgE4p
QaAtLaf1n1ChSma4xIGSzS5aJ44ZjubTrPp4i4jHObz4hlQZtKRLXfBfEurrMPMd
aerYf+w7Dg6Oi6RnTotSulPtEohUzcIBzV1YFSc1aPKYkvZTzfgZArvzYaPPGnJi
+NhLCWK2L9urB7hcq8a4ORaTEbmnyod6k+BGD12o9RksTZEgMB9aUYwW6WfTEFXl
HtOMLk1canVq4qD834uB6UkE5+U8TSVqLU890O9WwXjvdhFDc1HEDX8bWZT2Z0cb
otUWTfttp4ppCxCzJgPTED6tnXCpxKEZXdtV9cJorzN7JYihdh/0y+vL3y1aabGS
jt5WEJ5olyTJipqHlioH3y67dW+KTcZFu4IJcdWkerlAfRDPyKposkRNdCnEgM3B
lWNORMn3GQPAMJ54pF8HWK92xdtPlaIzrNn9+Pw7MiUO70c0hct8sUXm0Si2XZ4B
WUpkLSj7mM1S0ElH2+j6XoGS8OOSi4hi2j73ks2309BKfzt451mduIpYNATA4w/u
GsgcGIEPgsMvtzB6U7DcxWeEexIK+pygnSM37gxnuVZc3yF2Y8UJUagIAu2+H2LJ
2XEbpV03BHoVH86tC3hAgP5iWBUYEEnxS+8UMWuRXNDfjgmIv+36F1QH4Dn718gG
YeCBS9dL3jjl5aoVdCtBA0RNQxR6AQKgy8yyuB0cVAcjWbQC39bU3PEFKMUEOtz0
Cu5paTks05x6Zw5U5FcyWBMc6WTEJQ5Bd6DQhmvbLtqAhTDtj2x4IRwpGcO0GVVQ
PrJK1i/2mL/k4qpW7ATpK7/4H7lbpoA7Y1WDTjTis7Hd2Wdq92nbZNqrkx8Z2e3q
kMz0OVeuaeq15vctx4Oat+GypGJY0y0FkbdatyFIa02ykh8RuVYpszRt6QRyHWCh
oEyVcWecfeqj26xA3xJsrsAT7SP6fPTxvG7bjLLjPVgq4Zd2IDSe2SXwvwqmKfzR
0PrrOdyU5yi++AARAlRfXNFeloRVVayee7X67Apy2us/q/zRpEAYT3/EeQqVuYsX
Uj5FlQLTWOm6Xq3IWpRjejUFKKFvCbPHY0XCiEZVCqHtZRaVBX7OFVodvRP9mpww
qWHqN88UhcT36MvDY93+jNkk7zJ5bscHL7r41ePOMyWRD5XJEoRN2eFIePFExirt
fnG/NrTPrr/w/r3Dqp+h1pEjYrjuVBzlnwOvRwbudtquFPQI78xGmkNc/iu4soHA
a42hZZQbCVdNL6BEX1q3CbxtjPax54nD8BW5BSbHnOYRypZy0MORYzcsRMA5gh2y
pLx+Iw2QOepcWvrBHvno3r2DveI0aIjO36mRxkuYVF9uNh2sNKGVJmHDEQp0ZxbP
SjV135/uY8EESvG6wURjqocrGS2yBE90no2PgE7emknLg6TL1UAbgpv9JHgRl+d6
4uxBEDKpFDsVzXd7qY+GiZLIFSKqcnA+9se/0j2WGl207eg2F2eScuufo829PAQ7
kDlGc6f9/X+qkz61bJGsou3rnYgPmZoc9pZ054sUcpyznHxQuZkxtRYUkURnyooI
8lSigeo1IcprS9Q/CQixHmmP9k5XUpfIBmFBoz0vU9Ks0ek/9mZH05Fwv1enAPpq
6ZXtMHt4GAfLNzfMRDtr7jSmJF+ps6eypXb/tqDSgTBY4tLIp1jQ8tDABg63q4Mo
/YifaQVVTNQJwTc4QvlgN9vzi7ul+y1xIVT7MF5Kyw+N6R+V2q16j9rrFy0QnQ9d
h0bs6/8gtUpGNUIqgFPCXmFBtHo/lEb+qTbaTrbxbFSPhH0+AIvkwycD31FFXtYJ
vPZddD9V5JqCuhEgbMEQPUl5EkypEtj5EaTI7K3dTFP+gTqqSlorO2R0OUUnIb+o
bxxl7SCjoiiOKb0tgwtnAWptA+xpBWdFDi+rxuX8Ge0mEYUXp1eVWI2MTiZq9E7q
jDfde+4ZZLK8WOYok1OmvpzbjH0j6NMaBsj9wbCPQ1vX1ko+nPjb7nYbU4siI28x
3Fmfa/jAaEFmT8+zuuMT5UurI53z0cZNBUbz37bXNrhXtqYzh121xsElHq1JmmNQ
/LbRhTfNqwPoLxW5WFNi13DgU6Y0avlNs8zDODgER0CrIu6yAq4JYwigz95sqvbT
YVn9Hb/nopWgp0gjPQvsA1MAVYtVVu1umqYMfmhicfR8Br/bDravw5glNHiBCttH
4U1DqDfub79qTJYmVtmbxUkUQNhjerJJlA2KHxUvREOO/9M+md5tynC2Y89nrPir
0EQ5m62xXJktsky3p6CEJHbnQFv4ldyROJmOiqZWt3Fy5NWUiXwMYk+vUNMXj/XZ
DT9ksCroZoNANF80ES9FjScLxDRmJ6YXzUajiIDk/tSYFv6bmyIH9h3fRca+mpTw
iBsWzVk2YkLH4ZCePqcGFwHtNXrPM6UQInm8g6dcA1nBY/m0KBhOC+TZr9bCBIDe
a49TFj/7U8YWHvmUTMtuQ7Gmz+1bp/kO8N+66ShkA40gHJ2au/4JsDgN86+iKXlU
xLM4ZNK6Sj6MNSpdNfdSbMT69bDvDh2MBfS9eCEUdwHOArWU1vir5J7wXHNJ1JXN
Kd1eP6wpbpIvnnDw6ooGOfo2k5KrLjwjkAkVIrztT3urxZxIhGwbN9MRsyh+HVeJ
5cxH0PAtf6irQuyehYTeb99x0CKs+IMGow4uMEqfVwdfjKQ+EitFCG6raLd1vvJD
DgYtcy9VezvEbrLmX+yfrS+V7WN9+vITdkFAQznYmAPo/GWdDfxWHlpng0KgehfV
mMkC51LxfX1MDGhV1630S1sUGcq6oAjKpUwjaUUH+hKQANYP2fDmCzS8dIncv39y
0xGDvOPf3dSnmZKJ1nrI2YZDZNMjWRJWUvZbwGax5AQJ5wRoSNdQBkqWJPcO4Lm4
zaRKIeZw98b2I0HpmrHo4nAqj87QGXJ86m4NkEhoFp8asVl6eFrZiwhmooe5XTLD
WLeBFkLC+3Q0tG0P1qOcJto3VpIINc8rty5mcon/+30G0CzjeEI9N6pmWfYnntgn
d11CSlR3uQqL06GiANqCEATucLLTZUf/YYJV/aNgDRre4t8CFlb3EVLhXGCx21ck
Gc+Txw0+9ER4xqqdq59qbn/gpJr1dvMpleu5KeOaM+r8iFzmrM5XUvKmLwcsjEMo
g+3wDcR2cdf+QmvqKrEgggqUQo92SsjKeNjEA4hc8W2+qTca6PbOBcLMkYZ/nzkW
DZAMSIJOLIX/yLN3dAcrsRaYigUtOhAz4TNDxi3+0P5rsetU28VGqU9O+RwJgsb+
CaXAgvzGgUeWKeGOELcaCpH5u2n9W/blRQfNFRB2ed++S01SgK/irClaw3xlGL7N
zHwTz5whnrTOnoa3q0Z/4hLI54q9nPWRBRw7bGnA7rWEfHcsAdzPHZJg20KZmlK3
C0p4HuWbwykRjkTSM2tbenWi37ChKaAQlIqKL/1w65UjesG5OAs7Kayc69q8BTTU
QnxE8nNGOM8+49Oa9n1aLAfTs6chmR5e2Pe+PpmbTL7JCrwKu4qJPdZjWAOXQlxK
Ny1COZLOtK+/TVgEMbusK1HE6O/joMCbyvsYqLacLpfkRaAk/llwqIGrlEZJHZIT
FGnYumh3+kV/r+T+UFtQfY45p6jDbQpUP2DYjtFI0IVUC0Vkmlbm3xSDq9rAStBa
OtaPf9tbpAx6a7y7QMaMSOA4EkOma+GDDGsktCErSRLHsRCoV9c4rqn2xKmifP0J
3TzRrgCjIaWyMXS9fSsG3tuFCyPDwO6lxyB3C93YvjBdBhLln3r4rh4xKbA59UZv
vdGMBYeQGD54IIlHVKBymLUdn4fr6w0LfV8HNqILARKIfVKmS/klnStUl16ujkSP
Ixsh16ssKwS6n6D7kHco3S7Ir9UQHSHwdUhRvVYey2N7Fp6HN9laUlbZfcnG7mH2
NfY7jmoUnOjItNifZV3K14zf+I4mkYe5X6WxVm432wqHoXW8hqzf9eNDzfgu3kYn
1xma5yd6mal4nz8d9Uju38rors0JAWSUJfBBKmMVRFR/JtKAXfN+LDO0p/j/YjtX
we1PMqgxYsYCZr2r9jLLx9+j2qnQPebgkkAF61yx9zUiT/GWgTUaU9hWhMe4FrXQ
n90xLe6OcAGf4k9zYEYEBh1vd7TNyDakOpA7mRHaCymNLvzntGGqoggn+EIz14r8
+lEj5QZBIoCPN1tT9H46lu5FpV/XjBmK/l56lL/cHKY2+FeTe96JWxw6Axh/pGiM
XpXof0NStD4x3+UUGnWJElVCKyXKyc6t4h0odAUEd6uGnwelDgMo85EAE6LPPVyV
thPYAT/YvdxEQ9EmB9+Uh1tRm541Xm4/AqG6g1B5m4fUjmPFJBsH6qA/NjcDirjA
Vr8lmsC+kItaDFCQcGocvCxOxHyIXzWMrTVv+fSMPGS/Ec+atAaZLD6rmXyqS1ob
erWJoEZECvrrimsN0t0L74O0F6VmS3QVEpQ8EkdZMPSKRyOY/YZ/dF9NLReddMP/
6CvoFI/eUe0BosyRAYgflE0uDAmOj9mpH2QCSOJ8Y7pzexfcaUmRG233smC8bRFl
PEJOqEqT7VjCxqvMGbcXJiDdjL8X+dPrzkAn10wTMwp/vR2To957gdjLGOz2sjQO
UAvj2fz5aJ4/FlnjHhVRskKK1iRj6VJ/smImRNMOM8oZI3pc5QYCmwFBYjwDHJc+
iGLLL2/18yT7vdWwa3jazw9usFWg0IPQiwOXw8buhQtMTKExN9rNrmzCpnIscBSi
a555QLHULnmf2bWf0V+QI3vVh1fOdk/E0jxZbajyLrgH2E8WQ2SK28hlvimYUAjf
n+agAWCCTnwyRSL4EtlVzGfe0oGTHk0gJKoElouOmZwV1WSo7DXIG1Td2pwD48Q5
ngzBkq6fnN4zN1bFhS8Rmyswkq6Pkpr/0qODmC5miUH4ox8jW3l4hOi8QdV4YfIW
APYdtQqvskydbfuX3u6Ed70DHKUYSiwrjT2ZbpmIEWRrC6VJy6wM4i+AABUp1Zr/
dkj6s/vBJGKMkolrSqGaEb192uDKqPv0THQKfkxTP2qY1HZplrJf5NilNzQiHJ3G
NRIpJXa9kP+n5n0u/A5BrPrjVBRAcoChDohAi7ZCx8YMtkWYTsBDMFgPmk7g+p1H
LSt99xI39J1XZHUQRmJcdd2Etzbhtt6FGo1wnK+bYXoqnGr1d1/6rvt24Q8fGoac
Uwv7jZKgS46iwN739D7d/wqrgIneRvYoLjEz6vpacWebnqEpxWypaiKeHKy4unqR
KVi8yh1Qv+B18YE0QO0a5Bxww+lgd2Q1dPNFLTEx2ubQ3cC/Bum4sscuf0ukf8ff
TBzM78r2x3hjFjEg0rvD14YMVg0UTLUWptzPLbDPZU4AsV+B2fH5M1YRi7QFAWyW
XH59cnbxY2dczubSbEijDbu11qSYwjVhJlfxKZq+aYNjHd9Rik3G8vLbA2VZmOyG
5mtPVcTFQpVYxrwtWSPl/mU476CffQJxvIOC+SIpBB5OutoRllLTuRM38iX/VWRx
PKlKAslxpISudK66LUkAEUCFynX3KdaKTz3cuOYShMffIWkcqJS6XgAll/+3IdgA
MA9fuj7KMCST6U3ANWQdafseRVJzP4zxLVN+6ym1zuGwfUvneIQpDLnezJmBceiL
VHUYDdklaqNMg4Np7P7DEUOJzpVhADkmWrynUnNnePvR1JQAW2Jlfz2mUVthd7FZ
av1lCQKGke5BFleE1dHD124pZeUNVBmzOkkFFwEqFXU+gJrRIU2obrQpCq/IB9H4
PGd2YT/3z7tJSI6MkCfiHEzdliCb1FUn0Oi2Jd2rsEGeF30UM2eX+hw3BUWNQ4mR
9j1dobSdA+qpLiHLEuQLNJd97DtwR2A92KJlv1PrMwtQL0tYqeTWtc4X2EIxX9ZX
8GxxuySuMNxh/ARr0eORDmLp2c8sXNtVvSO1tPo+WcOzVAII4ZKQzTDQV4umtVYB
Dwh3L6dGV9RAfTVZfuZVGBGcTE+LinoNJvs/bclIeB0iCa6J6NSwfY4VL1yGJeXT
aJdfpFRtAZ1XtYzEUEk0Sk5oCECMmK1Jyo4Ls86b/nXr1qyP4Oj8VBGrwxiNpJOA
1H1FunTqd+Y55tjo039FBl+stGqFl6PjTOyOYhssrVp1BYLEMW3k7D67HT+QOH+O
+3hG4Oh4kSkX+HPuNu9d4De1A1OILpyuYxOKxpe8mdk/pE5Lo031J5yTqTWt9J8v
dkYs9VYXk8voN6ryiIfSV97c8ejPzXTSG8SoFmZqukvLrTkt1xQBIHTMcdJErrnO
vz3EPfhhFGc3/AzX5QIEsFYM09WUwUeNbCWNEY4JyYEyvOUq4a9SpH2Xxm9RTgyJ
Od+iOsWgSQJ02/bDwf8F93JqpZEznGzLZ/uMOOhfv1yO8O6mGOh6+G2ZoxghQB5S
U9zxECj0O50OVqpvaJV27v2hqNfHz6hDVD0grDBp0Z3YJtra8XE1On670PTc+fMt
6/4xCr8zVk/3ex3Rk3kTSCWqN0C9UQnStYvOBfFHQ9YEMrzHTI28uXdCm3PL5YLK
CqKLNdo8pTfU01NExbIEr+/UhlgCvV3JZLkvakwBFjrmrwnzwSmGtnRtcoO01MnB
8zH9mszmYruWoKhPnCGtz1TxntIbJW7mLIbqA+LXDtEBSYDw34AYiKTz84OuHctA
aI8xQwxu+JTH0pZfXgB8x2yOJPY/1EzK1iADLabOlLgETAPHfHFZLmc8xzSul2k4
+JPMvjtVimbDg1FGaBTr5R2wXJvkscUha5ArT++NulLWfb6apAA9uR3LebKU5AbH
1sfm8/PXS80mByO1CofcrIkRfrfSWvS+t8q17sIDk/NXdCgBlD952OvnyiUaPVNY
uvx3EjqnivqcAlAivg5P137WqYs0ti1tIwJ1XAFZ2nZ1qm5ld8Y/iGRrs1a4o681
yds4qpY4AQy1OloVIr5t6WlnIujIJPY0GxFHVjb7mEuMpI7b38YLNacyIUiqrjte
SheotM+GRMDhUc8uSiBf7dSt70p+6AtV5tEOzhURKRBDnFmaj9vxWyKqGjvhaQpk
8SpnDrYnPdNLvDmABodQE0e0ZTLSlKeOFOrtMHTuXIeK3natNMyOoe4zW24u7m1H
cCHFPppKZEFyQhVrbY9Dg82GeU/3hqtp5nnbNsaNZttY5ug8f+1UsHn6uvl6Ba9U
I0r69WYateSEKzESAQF1EGUlD8cbv3/6Li8rm0zmhMljP0BMA2R/n7YDzNt/O+GJ
PQeKWaI1LB66XjylHv3v8nJon84klYo4lAW0GaTnSYoN5o7BLBDnNCsiddALMdWT
Q5VJZl2in+oD1qEajQzb/Or7YebOFkS7o+/FmbDLHXdnERPxgJTp+nG1uuvoFbSP
v3cANssOIZk4OmsJg0EMjB/DQfatsrct0OVxfCiRLPyqPJkzsE0RKrADKkBpAxOK
NN5RCB1DhUtjy1mabyTU9C/L649EtNHNT3TRhgcjS8Ic5Geuq3nsQm3T9r5+6Yqr
tYWyTc8FuDpXEfC90eFHtVVV6uXCNl9ayjnhc9AqblzN/BhW2ZujuJoRT1ujXwMF
4EjeqVon9rYDhfF1v8XR79juy9o7jywhgTmMXAMP4Kfr+0GPZ39Od5ujV9NcUgRv
ljlIX5Q9zXJTflGS2vyjIjye3sV46qB9b4kBHmp5cjjg9eyXwSfh4PvBmziZi6lY
kk5O5WOWKduLihWI/YD0xFAwh2pRghtV5skZ+87bJHtCTn5sOUkd0lhBmwtQyPZx
BQC+oTMofUBZ1Shw32PTvWVOvJhLFLP+8p4a1HjDt/f1AtSOxAFNELreNEtQkv8u
dTA7ZGClx3ljeEqL2pc0yeJKwUDowiH4/+T2JafbSVYPpAGtoHlvpIItQCUaC/n9
9G2gKW6AJ1Ornpciy1PBOw4DVSNNHfvtz/WaGWlzEKOeeUTZP/+wPgR0m7dhqu7A
Q4nu+WF/fL9NpFiORPTnAcl1gOskVba8N9mZkNL2SOV5V1bnTM+S5B/ofdhO0kgU
Zlpuy3tmOCRiAZsz0T4aqZTyuCHWNMymLxSrHSDXuR7AdnOLXkKg6lpmGQqoxIzh
Jb0hsvyFVL1ww4UCY+vwI9jWDHRkqOqe56nKywBaqJ9mWjjt2bYEUEFZ0KulBcGu
ZtTiuOP5USqOdFeNhJ0zX6bdvMRCtFmBCGtMUKKKbGGKRo6xuVD44eK0FHpdz3X6
mN/sccqPh5/G/dtFKuemesznq4QZVLalsd5kFk39yO6zHMOoTQ5uFAb1mQ42jLmJ
Qk9meciZmAxS9vzb5bIUHTEVASnF1WjcuI3rqyFXEF5mTQoNDb+TYL/9HUw6lCQT
syGzKAxwq76ef62HMtnfJIRHnK3EKlcAvGQgN1ncYniXtBh137rxbDe5UfrC/WyY
yDNelHCPDI/xCiElZLemRjsp6uzeLrCi/ZzgiumrIUrtDYmWrOvNeIHBq8L9WFuo
2OufUMNfHNBUj/cZWDnGWuX1XVqz4C4r/nasCQ8KO+jqRy6f33GSjkrk8k4J1M74
fzHXKSLIQsmrP47N72B9vx9D14OGz9NOORkob/cwxetZDUuiWjPJpn1cTvgFzdhz
S1ABrMLUMgA5OE1dm7rAZvtck/QCTiJQT1MPK/V6/z8QENZm2ytIhROkoZqo5h1U
Fmu+xqT/3/pQGieicv9ydss3/LFyEkW3SidFaA81ooeyuzr99kinUBtIeF26wSbh
WGsmOE7dgLnEPjMnu4CptT04l5itSo4PYkdGMg2ZWTzD05QvOmamW3LOCJsNaAKo
Gvox6vcF1GDVy0gEzKuYAZDpi6sffCxe5GjiO9NiSw3OtkoY9KD3hCxDsOMTkOP6
j0B7/i8fFDdOoTDX/4gYY6S3cNApHmQitXaAR4sVJxd6r4TTZnVb2KJ9jfDXc6U4
9VNjNQTRPxPJ5daE6l3PJTqJmqQDvPbRHR2D9OygJHldU6ss9kAyfoopUxPDaOf7
RDQvvvHgf3zNBnVeSdR6g+TnPrQo+WfJ5PgEmVCbf4ou11H4QihXxx+t0Dr9EYrt
sWSGEIQk4hklgm8BiQdhHLtcWVFIH37SKBpq0DGm1vYS9bY6j8CfgIVHYsQH1b3I
JUEmHgXgWnX4oho6f09dn6Ybse9R2Ga4U4da1cZlhoYCxUNnUmNf6uf+LG8DorOj
xRezIouyxGilTaPlCOEP6stGYR/OeXNeqAQ4psNnq8sui66quR6JUtuW8Ba276Bd
5x8PjLATfewA0/YjsRjPNa/oi+Bim6ypOyeN9Rmm/7879EXLGJWdOIKBnwMPqz19
TGIn5dkaMrOAfRrPiS0VXKM+Iv16PELyuyZ/ncprBUcw3Rp66R/OiTpPpkP22xmX
LP9iAMY4UuDAimA62Opln8XzWrQp5AmzO6F0FqsB09IfQT5jjikgO/T3cKH/eflC
A9hLydI3tKFxVQuj9qN4rSiXta1VIyj7axTom4xAh2EROPic6DAwRpSW+cFHMFn8
1UrkfG2ui4+fiEUcz9Yjji8QddIM5nXgcO0Bq7AlCzbM1boT1B0nvqRZRoPjEc/T
vH9OtWrQlMib8sk0+SNeGLjQ47WSn0lLANZeGI7axKg3Roc5yUj/yRK59Lj+8Z6U
XV4GFKh0zHSGY2fi5CdaKfolEgNuaP73cvQYM3KPqSGQqleViJayKDS1pnY8ffH4
0QTdX6dAVmKnygConnv4Xsc4/XnuKhHsSUjui1KLAsoLZD05MGjagze/TGUiFpGX
RzNsrDT3SLszXgnW8egnQusiFLqJjWdCiFyZRhWU6NqxvKbo0VHkTwkmGWK7bXJ/
gx5fie/mry7tWWXrwb+R8gsrbVOH4n46M3sfQKEGDF47R4O1I1hQdULuIEGGY+kX
4VDIXeth2YQFka1+J3UGBFeWTonzMjQYJa2Npn357C2JEHLXnIyKVWP7EYHTIvdP
0/X5nt+B5CPYj/1d5uLnyaznLUxsDh10FkGZm0ePetvU0hJ7Qo4iPkXvZONeTKwz
MOY9R6WNDl4IBcnaJLQyVK/Rp+GXMOwfd4HC4WH9Et65mEUR9yeEuEdX2ozQWf5E
ZKSM4tW2gKxmU4xikxXvdq8f9p2Q2LtqUkMjAIbEu+jNtBMjNesoOua+Zra3L5nA
A4qvYnDYEDxz4n4bcxiXQPWsSZnXetN9w12ynhMvohFubmhD3EhI1Bk1K6/3NqPF
Ibrji/NytcRImNV4LAi1Y/ExcVPOvIIHZKWQnSfKd0FQRbN4Qt1oj5b747HmEBNn
fQjhum/TaQNWev9BvU8SUnwl3SFwhrf1AspDstgIKcldNKTiC8mE45IWoODFbBvl
LSyG7yHvjzmyVf3hyZ248V+FEMq/eIBdZtp6op236Cu46KPhVgy5c9K0IWxLfBxM
/R9k57vZ0t4p2MaIY3qu56ZPBwBksRltNskgtDJrE9xmpMX00GigK70YGx6QAoe/
XXfb4p8k+BK2WTVIXgHAvr0z+GQ/wPT2tPio3YsRbIy8ZGX5rJpSd9B5CfDGWjOC
aWx0FZ3i1Zo4nqzOe0WOEVi7gJ9ZbLRzegXIpc4CTvVpY85DlUZ10DOXWOOYyErf
OZPfwQ/J6Qtba04HP91gzi2CBBe6W9+3cCzE8+WP/8Bt2zHqpTv3mpd1UTk++5+s
DZkR6XdLN9aE9jcE2rRtyhWokgDvdCPLRsdNtUQOfOp3l+C6ekUOSZooCg6OZ7KI
wBj3QfZWVfzMhUqJxdSXETnJASiRZmQzcqm9kFBqgiiJoK5ds/1T3ozOrlYh/im8
J9sW8oRM1Xsk6M3iVwyvF4SknsfkehlvYHN0bLmjb/9pZajpIiA6IQ55u557Z8Pr
cmt5QfvtgaYkHOQ63TKD3zzmqyS4jWv/wHuiKYMjgaQvhurTHw+VsOqmVsSUreC3
f5ZKy7TtvQQZ4HOdxGpDCfYOJoEQpOBoGVQrHRDhz1Mq+VmfCYxDhpvWWZIkQXTi
JudWXk8nTejl8+GstCuHeC7P1g7s5lPpYSFfNQeui9uUDBhjMJhRO/wyEkMLxDmZ
vB0jFzcYaCZ/Q7ga/Q7KLoCPtmVXB897ikW8Z5HL33O/ZShtim/ijqkr+WoWHMZL
AjZZuzEsRhizn6zmxK8IFyjy6HBi+43N/yHzfFIyZfV6LRXXf0CreriswF+UkwHf
7m7MMauUEscGhwnvHlxwWMYIMyGQZIGFPbTdeSKAf+faDSL8gUS29dnVMwKWvNSp
BIaYAsXqPLtL0AaRE6VVPpJB5ARKefd+nRGTMI6b2pX4FnaElTW53uCuXLok0/m9
+rXvl8IXW1ZkXSQP6fiSnBNqFvcDV7C42/cKI63iT1j0gKQta5befu6rWhhYaaZC
13xWxX7n0fLFnYGXPiMk/RxdgD1Vfq7aPW/PKR47pXPEqn519VYSNKnaq137ReUX
nFrfOjvOpVTvuUyXyA/4vOw9vdGHrkV01a4NhTf2q/wZgDbNajeUq5xFAKW1a5Al
IA5lJ3LfLvPeGNDdInImWJKYYX+7sVd9D5Jx+fb33n3Xgt+V1Uemk7aKV6rs4QI+
vHIX5YaVAXkvUgTAWoBR6OEoAkiw1IGHjEPwnQY4+AgMZcqbeEe0RAQpJzblGECr
4Zc2MbUYbo+eamBFcBDWh060aRTkjntFRjoM/SS4twFYvrBIHn/1A99W1yBJr7aC
bvpi2HYLzGOqpN6cebs5WDwUNu3DMMRxcavXeKompziZI6lbnpJA0ltrKYHMzsSU
aXm5/8LFj17Yvr7v+GQa4g4drS7Ab10jxSUu96Dgxf80mkfWT8echedtO4CMnmim
x9QVhGK8N7GGL8IpGQvB866ryR6ejR9O3Cs+bAwu3RW3MNrAAUiQx82MVsLp67tX
tsaFAdAPi/WSHXtWk4cFuaAx5+RGKtDzA5JwyMkBKYz3/qdzuAHWyH/3clKP3Jhx
xRzhP5Yp6+rH0Kz44D1GGFjHKhHHGA/4GWCFhvtIH3X+efuM4UIIznHVfvyjGNcO
sZ1fN3GSKRhblEVO54oeTjEWEHAyB79p4Zb3l6cjp6+9RCwIvfrsak6rgtpTPhyD
TAN7cKHMQEfQ8yqhlZM5BO1TnCqOo37G84zD8WR26s2rme3+UutBmr40Jml43b3D
0K+65Yz+1At5LCDXrA4vR86ba2SzDJZVTODxdfZcnz/Zwym/xQuodw4m+fhZ0uiA
n7OVuGjWBCX9v+yGr1b91O5ja2GvY7F+2tRTWh7Nu4wMMEAHLEkK7n1FeZdfuuzE
gGQYXYY5fRBhJAQgBMwwTDOwESnmutXsTJSzjycgv2vAMn+4i39BZBqa6GrJoC2t
kn/pTmHyRvE/oWrRzEsmXMc5cJnPGBXwRhQNSkKGRi1zS5k3AZMgPdZiul5Ld0xi
ruUbgsdj4hnztmDpjUWF8ORFRooOW23sHCIjpmdvRwtCi5IiE4EYXLfdtA3RFoqT
WaH25F1z7rI54BIfcwTeNmpCRQxaF/1iWjHeRW5FuLq6ZSWdNmajidRWGCp7e1Lv
Lm/HESUinloWyrOK6vCjPUvu/J8/iMGNUH7pIgKS4f+8cTVTibd6VBhRzsVl0po1
UJtxN5IjxA7wWAAi/NdX1wkdBEEb3YVgYmaUky/FTltbdEpa3qW7Atw3DhkINAD/
8+fSYMy1K9cBwA0Ia7RDb6tEHLHWCi2afN9rlG2ulrrXmio2pr2/uEGpUtTlYz5N
2cFoBMC0sVWIIH4fK415Izw3mEfAYJKtvySjZhX1TswjGeVG9rDiM9YdDgHYv8jd
bWcXGB41o4ZHC1XVexm4Iy/kyb1CwvVNnaCWGfmY1VyUgeyjWs85w9jL7+JJjRZc
Obm4nqF+j2KYf5VxoZq+pLkkkIm6cgG8oOwzG2frXJ6jLf94IgYlLkSN0eLsJJCZ
bq0OUsk3jtFjtMbYOP00V1tePYE+IFQVSPRzRNFM561uv3KLcr/z1BQnL9+l1PHL
zCRHLTFWwlimy5fAcsSuYGfqTDnNM/hY2JzIhs5UEySk3k2IguvHVHQnZZF4qjcj
ZZODBCoNlBI/4iKdJXhaTRnXaH6TgZcL763EcvIyaC1QpFVgJJUankIofrKo4lEE
r8SuIbXksrb+gnv8xWEhyScn4X+w//UQ/Q0AecgJqr5HgmiBah1txXZrY1M9rbsr
yWAIUDCoNGtnhMNjk06mc945Mj3A3TtrKACTEBd83gSt19epljINcxc2h1dAFpmn
NYoTqyzEQTAqnYiFc7h+gTlHUl/EH7flNOq2QgS1Ca325hS5vfT/oRFWsMtoVP1b
1bVkpEjDV1ReQwH2g/5r0w4F1Q46D+UAeeTviak2GIXKPST+WZIAf5HoTDg3YhLu
RnPhe/Q0c/6hT/ivNNA8xPIs6qnxK68M24KmcnyvYtPosfu2z5eOAay5fcAuYX83
xXvd7WOHssCo330Apbj7ZufOjZ4yUMbyc0HlRWEmDznDb1P2P2H85/Y+ne5sXIra
lTCmV+npTNvOvO3Bbc4Fx8KoBEhXGI2toV42e0RCLVM3bTtvzwdx4VhBmh12Vm4d
3LGjXR8DASGu3/HdJlgwQm9aGCSmDGnB+Jy/nZ+O/MHqLDZbTA5JksA3Hocoip3f
dUyUzh/uvZJB0sBH4vD8mHydwTfrAUVgoB/Rvst4Lhun4XFec1oEE+bUxRb62Q7y
hBIVBn7L8CniCJ1XZPe/aqbqnSvqPjZLOPVtv9fxNZm8tsuDg5NUPiaB0urUGj6Z
UvLGMjGz7oXWrByO/0WhhgextVKcso0No8Fl3R0rM0n/w9ZZQhTfRKs4625RXEUX
mca3NLLhcHJdqTMb0I6VyIyNV9MXccK6JpwYnaQIPwUO815fbvljO7x19j/ssg7k
QPymFABG8spIZmNaEwOd68iLoaqrPMLkBW2z7PH+QdFyqqtU1ZP8gQ9zH0MJmO7M
BddbaMkej1M1EQuM2yJ2cahYc9MtggEju52ucrgTzo07NklA07G5JMehLRA7Vj/V
kKAmNM1Pa+EXr3JSTG64EqlFPFOhbxSQV0vAxZxfppqlQw/1lfB6TBJqGhToCtCI
Wj11RI9OcIrQ8/WdPyBRauBVI4DqQHdMzpNFXWCh5McUitvItGhkw9tsT0uLgSRs
kGxbzXTo8N7rGMzXXZOO189ql1aDoYCugR18UJGQpaOfsZv6ZgDW7m9eUHQJ6lxp
QBwq8FlrnlECD4vlg/oP5RA4pl1Ag+HChZu7k9rfzBr2uewLA7v1q61R9I25iKwc
ROOQ3/b14H9bbDMbyZGJbshjaAYPU4ob6UATto23mIC7EjHx6E164R4+nCfVV1wb
kn5xEHz/f4+tpYtK0uS4j+GhjtUkETA/b+8a9DdETBu7lecNxxiLUmqMGbdjSIMo
ha6XybcAHplRZD9xbTHgdUyZwBJUKdOqfo8Ql7Tk1jBxB9H+ygjE6g8bhP+cNrzp
izaGlneKNF1iWA+RWmiGKPywkpk0B92AD3OahUiuMCTAsmTYNf35W151uvbjooBx
iWcf4m7G05Z2bQwfVnFM+3DVXA0Xerc+k3JzVLJtC4F6xQ7wKlkgXmRQsMpnGRbS
hf3lsTR3xbhoQbzstxsy5P+n+2mcCnT1RfnsvNrafmd9hKsBjuRCpY0K5XKzR2yR
o983iwkddwZBHclmd1/zIry7rgZYgCM4omf+22ffjXNAVJCihSIMX1M2DCXtYu7f
yYdrndb8O+RuFyaDeqzE1nCbfFfoD9Tui6k2H1NTYq7i6PY0kJuQZlC+sqvvHCf7
gs8NpujIAEU1JhjNMhHVPaKDT3i3WUxhnGo+eT1tsU1QUAc0+B7AHyPlVRhlltnk
DVplKwHw8wEu2z+xyNXrmfcB9HdXASwA2xThBsIMO441LUOTE7xNq/U/8aGJODK5
KkDLt3EE7f4afZfew9k+fiRjj+YAp/2R11mzWtC+84hcEuRhtzHXVLYhlTpMXcUq
zF5fas9ud8QFyeLPl5dNK+VV7u5nF5O1rM4MsVa7ks29/P0B0DR08irqZQIGzp+R
LWq1w4I+OtBjZUCeuch+l5DAIhydwyHKQZW9/Nr2XpPqN+z7xDexBGwAccx9RjDv
QF7KZCg9cRSq+Ry7RivJYOBs8/+18+dTzIwo1S5rAnFJvCfrawzrtBSMgvmX0u0/
HDLytzBDhIePuJGPVSF3nXM2rD+BO96vzkaEHPMT4XvChE2kRJ3JsNaUdlCp+sX1
v7vkccm96ioxFyb82I4+4SqtGzFiu2EEUghES6qmPsknGAtlOQGTiJvD0zeGz2Qb
QZhjgnGU1PTVpPrsPyIt0gfDDitcW4kMbwdJJn/ds0Cyfiu/uGkFVD9wwUkuYVFm
17ExX3GuK/Tc4D8l7MomT3AHdy9ZL/ZQW/nF9eOdMz78d9TQvX4tQEilhhLtd5fl
xPEjJ+1SrXEsx3YQOJgvbqu77v+eUejKxaVcWe5Oa/sv0x6p+XYEgz9iFttSIIN/
csAFIsjYgV82Zrwr+2P80Ring3u+wAd8wHQSD9qg4JcR8GMGREOmpDBNRfjccdc1
TwKiLWKrV7qZE3+h9GU8MO8fgbgE0dBzJqarn2tBB8UNkEwK2+mfvNj2CBEY+LU7
KFHVV+uipoe5DkxWJlMBgUSUmOd9yN8Viwf48bOmSwhzYY72zkyBgygi9NB3oXki
+noWeS6hpqt0Ohr/0kQW5AjzW1tx8PvTqNnNZjJyFSsmF8MmmuKAkW0qw1HCIQqZ
sE6tCKaHMlQBGNqrzRE6UBGsYHxr1JWH2Wj5LWUhlyasw453hQLRvsLYLPFzxY48
QoDyw87QlhSXgiWaC1oGHVgw9lyt+X3417b7JFRBRmxV+ZTP/GvvnLR7BrB6keVW
g7oa2xPHI6KCV5hjJuXBJ7xWaOCbea5J79wqeSqPFaA7E0pSSYsJgpdjKNXpNVri
+JA6mVjym+S9UTkfBLfSSrhEZo7LGhDvRZGlyd069SGz3H1FNOwZyEjsW2tm8PG9
3asLajO+GTV4hU5hidCgPa/NMIxj9Xr5+B+eAu50w5FqsPILfuXpWcNzpvLP1WXI
p0bQCG7TqQNvjpVpbvo64pMWOOaovxfrRGGgQgHf/nzSELJzCWH4PBKYU8uiLNId
tc743o1gK8Kl74yEoi9u5oUJcfqJJG0TD9tiJv8pHOkkwrImRuxJnEn+uRbQMxSz
HLQ4lI9ukrJHguIqEoIl8vyVExmzkubBi59BlxRqoVypzVEJfUtqXYX1wDhTj/yz
EVxxM6XAmMilDkMcd/GkzSGNmgYQ7M5/hOQbtYEbL9akuwthz7VuzTgZG7X/RvPP
1u+AgrVcc4ySlvyRzmHQEZ4g7i8vvz7EqI60kXPNOuown/0b/jDwi2lN72FiCayc
3+GhHjkioXkiM4O4pJP5jRck1SJxQnnsVgFBj+uYo2qqOJTDlTOCqRvChOlwN6gW
3/8SU7TviLXtDcadc9TWR5OiF5hIBeOY6Xb7SVX8uhVgJdFIDQxESTZVKcRxv1BG
3NLJJyVFdybUhiiOdU+afeGKhATDkDn2bHzXlCt9mX3shmhWWr7vsbmfgpN1QMVH
00w7bx0F1rVBLi01GMVouKe0fJCeSE6qx3sR7e+/L7qkxZ41i5gg2d0eSzqzRoMg
Jvvyp6quG/00ULxl73fkE2tfLHPzeUuGT41zW/cSK3Dpf1oF7gT3vHAbtp+OvdCq
44XjKHS0S39v7phnbbTtS+DOmRwizHWukG0vXkKhk1TDCmwa8ZjERmBm29JkuesB
seM0mOzrmaWhrlKyWxMV7U1w1mY9G+pHF4BgD13/aQXdyLQF1q1jbqubG+so9KAw
HCIGMCv4l0mUD4QLvIuZ+BnmZ3wezUurTlqw5SCShtWc0DsoQIfDSqMHhsiVz78s
b0IXUC3lupcwbhrWdUxyzOBSscQfzjKEH9+NHInN0ZDhDz1+5PeM8n01+6zpUd9T
XAZnYZj9yLRNFFIC/Fy2CTyEGE/tfErBrc+XMcmF7VY3mi96FCikqBOEWYa5k35R
uI/Py6+Y3KCpKTD6RGZM0yiWgBwvoYbI0SUxbl3q4VvVoZP7bh7acI6s8mRNkMei
IrMCALdX/5eYmeKPLmxztqSwCboImVf43+35vbAiB3M9ssJLIO+F8utL52yhdDSQ
+NMR9uc+ZR8SEYpTPTfPylSWOxuc/bQTExrDRpdx+2NprDS9tjfvh9gtKcpJ2Xev
Ua12xOusfnXiYt0+K8JL7J1ED+P8yyoYaHl51m2zwGPrHwyRbloTt4pAXtxDT0E6
mBWpJoaFd+PguYr2SHo4A8kioBLKW0u5OTIhUKR8Z4tF906//PlKfaA+roGqaawL
RLRb7cyudRM9HdaMrGXKa6/1AuCZRhOpM2pWV+t4KUKt9niI4aCCksJsx1v/q/xS
0SW7jF+JVmAGLOulfnovlJ0CFDC6orHxRCQNjJiuoJ+FwFdriv78cGs+m/c4MYVL
0blDYufZ5rz/1QdDeST/y5Q+GeEOZaBiDu9F964yzKt0XRbFLKhAT9FMKyCWpIbR
cijJsHeKH8iP8MuQA5Glh5pA/HEErxxmLhj5G1tKXp0sX693fV74mV7RQ5myK7/i
BckhSuwi7ZgdODgmjOtyDsUbtKGAZXngC2rCypbdRP5gJI2UcpUPjqiloRaRRLS1
JLMVAyfoL3WAzNtpybRy09aY8ZDnIo7LmwqUro8dVf8GSZEvcVJ1gdP6r0fOqlte
/vqlIXdWqHCfm3Nd7G8daw7Yzi7SkNUpVw7tx5Kc0Jj4Kc683Tj6yPkju+6eyvGV
e46U+Cc1ms/uDDywj+sCJTjtFhye4YfjYAiQgG1sAraWhkgzMouNcyfdGEERcpcJ
GRcO8r/ptlBJPpepcJuUPocOoX0+1x20J9VQsyZgNnJ5oEWnKXWmAmPm6CV6wZUK
aCKcQNx/LQw0VyLOIBfEs/3IGRzunjygPocUDXWMW38l0JE1buvb3oRzqrAAxHiZ
3Pts9JpdBiBJTdbjIM+PKjLY/Lg7keChAs2uZ2LcAwFkFZn7L6MKY7cfsaUyEMJf
ScD3noPjqh8KtieQ6HICGGbCCkjJy0ncXn44sLOqkjL13IkDR/c02mBPA9jnHYHs
EQqfjfZ8vA4A6xHK/bhYmJVWH+4xjLu3iixuUNPLN5IxECaW4wV+GYsVofTjFghH
mSS5kSomAIkG0cfB0yQQ1A0n+N/iPRWABabh1B3Lb8dH/xDtwgYmoLqAOcT2kiYz
FsaGsqWGKQSIbMc+5e1qO6jDbhD/FFBSBXHHKPeDHbDH3lPm8dkl0gQ05xWz4Hlu
AdnDtbCuZGe6WrB1LVgnqxPyzYfMdzTHEIVYgAXklfowXb4cLh5C8SlfbWmJJ5gR
N04ndwdWfsb44cfcJg9URe9r3fm0HAo1xjhbnu55RHwPxHDAM0jPLPh2Keh4vmhP
tIFpsd9yvIsJ33mexWk8glxF0hsw/SmvJ251tPaOjEMLGBbhkp4JKtZ/sRSi7aGB
7G2bK11oEtwL5iKH/A22yXB9w+dpWhcjbhf0MiK1uyvxpw0EwOHggsHtKKrYw1+I
zZ7OSkmpQvHaR7VL56WEaarRxm7prtkiA8uOZSq0iWPydvxr5t7L91EImBudD+U4
p8PbVUXvngXRaRHz3wmQ9Bwe9mClAlGSxFW0lUgQ5wu5Ia3pcoqoDZN6S4dk6YYQ
YD9quZ3Kvy14hIj9lcWXi4eICjMzHWhkYDnxJytPaof2menPTjE4PVPoxdXdqvhZ
a9JtHpWR38rxSXIabOrdLi78YQlYe/aHpam0NcxmJdD1DNp5XBREtset478NOZlH
/FMy1mDp5hor6LuYjaogxFgDDrcMAjxu499PRNyRpMEMnH5xPLALv2h+tHaHhkK8
P2Qe46yMc6nSgpIdnE3Gu3vIPxBUCwsZX1V6LtsGZ6UiHyh5cWWM1FUktE1/WsEj
rsbVVbTC2K1N5XfPXyQeco0ocI65v4Dl1YQFEKBlgzBn9iiegtRSzfhWKOlqjZ+x
pGXkMcnAHLu7HRYTLqtZgbj6xvp4HHn84H2Y7+/eJ09k5RWWlIWWV4l4dbUcQPN1
3295KHWsBDZ+PBS3rfCCHgmznKQaFL0upywkSfIkjaWwUqKMuqEexyHrbJCUR0Z5
VvX5/bDCvtiCzu/428DBgo81TEmBn/F3luN9PrOJqJg+/qT9b36ZAUTq813hpyFY
LMKvLwwf81a5xx73wDUtuqPEGY+NJpkyd2nyPPdGFgPKRwubj98Y3VCE2InMDOez
V2G+JfqsFxYeix9jDsZyh1xciGdiEWF3dvNHD9uH21Hzf7h2MFUlo114af/asbeE
62cZH79SmmE1TUGWTDdXtn5bYvYkX00tL2smBSQ3f5vrrp8ThqI+uDMuZ3YiNnm7
2Znp8D8Nyo2ZzK9IxaE2j+hnMsjcsqo0JyyvDQj6K2jkkQJZyvY5b4RjNrlJ1xij
UHULDkVO0kyQ0nVl9seCUCEKiVMRT6YlkLpMJhOqO2oZX00lcFP5wo8F0LuBwYHs
ZojFf7pK+jksfgHYcX49QHbOlKH7qsi5qy54yPRXcK7aegLvDz994FUWV0AY167m
uCl23O/eYNUd7vdR6HohY5Ax7QI/TKqBkmAZRaZFwhTej2ZqVb0YX7xZ2JC/g30H
upzk3PnWc6ci0EnhWwWBZP61Y6CVEc3cpgRXqnxvp2Q8pO7FTOrIig44HzMH2JNf
Mb9jfFVUknWJFY3oufePr3vC/e1rgJFYqXWY8JQ857eBtIBHa3YUHyWeb/3Nd35t
wgbzWJEvMyeKTAcNe4o+lvKaSbOpur3twzG5H/3thJN9gI+TOjduxLlZDrdl+cJi
K3mPB+Zmnuoq9ubh7/oseRKRkRCWZrBVby6pwgLXPMZiHOd8zwIso4aeGMN3iapn
GE293zIpBFvNalGlpuu8HTXEbvqwU702QQt04dcRHx/SRp0ui/MbPGfLa8yASl/F
cqLhZsM8BwWl6nGjQUTQRcbW7v4PYnt52nxYqetQJYqwgY0NFGRsXh4HQqWvo0Wd
+OZqMzbcvihXHrq4ZWiAjKUTSJ2xRJqh5frDRrxcLrpmXXgx+ADghk+MW4vY5CPM
IUoyQbWLk0pCz8yqueePuNDRvMqjVK+bkWuAlSYTeb6ZM+2wwh0zXULa/jnfs7UC
uwbRF1Cns8MnN289pHgZX7v8I9gulBukDPZGhzfUg/BVFEprAJP82AuO3fnFaeIT
UmvYnZ3lYPGEsTDneDErxwXU9e+j632PLTexj8cNt0Qkcn7VpJHT6xqzUhABSb6X
oayO4i6aju9yWtCaHCfD/5U9oXSncNg+lHezeKiltMpxj57RzPFHpoH3yi9RLLj4
3MVjbCzLWBB9CQLjXxjetX2W0YIKIg8DhiUgyoQhnghDw/aY+Wy88YMc6Kj3Kkg+
8kTw7EPOBGi2JpgHteMrd1fgbidd7k3x4pyFXF6mddgyOQOzYcPHMmMaqKkk/86y
0eD1XXM4PKwppXvOlyyKEaNIv/qse8IOHTO4qvNmO9D9EQ9rjH/uGc0Lhp3vPNUq
Fv5uJ6ZbGwRqNfaw/xyryE+KA5TqYSKQGbROFw9ngo0dtkUhqQexurLVvYFUEIx6
4W5vAFOrCx5bvT/Ke6H0k2ItIyp83/APkixZBARK2y5uGtY60HsA2SY92DIDSNOw
Zzk9+FjzcDN6dglzQgy5S+9yDXnTUkQQ4+3Gg8nfBAv5XEDlTN8pNer5r1P3Qd9N
mIXGXG1fW3BKMLCAuptD36njUdqAOCfsokt6lbKzZnANZxySyiukCFzDRRk1aaiF
TfsCXfGSyEPYZGwVgYILeaGHtOgK0iQDNKyehUdoaiC7VF0FupDRYRZyzw3nF7UB
qjqhNHwn5hTL7Sur9cG6Y1R6JO/ynSl+VtoGjkGKYB2CyEOOxbCjC7WLyjL8PHOC
3XVqqzxXLdivVAJLUUyGze1638YsrFEeR2Zhyuzg6+8Gu4pglDTDihS1vlNUebFX
awDFaTozqfQHs/MOq8Mnzm50dwmlDxjyoPOk5eFBcEb0uI6e+LvTSKrbLC3qbFmk
9Vza+Vsrytb7GlGaeJNH9qpkTaQs1LHmE25hJp86c+KP35r574LZNxf15LIcMQ+1
tUOCuhZzhIHM3bocQBlbLHJVvL+hhWZgBaui9TFhG35jyb0i3w/ao7P+WatRl9Nx
PCgeGRYVR66WzQcSuxcNL6cYUAI4shxXoY75rKq0PzGlg5iwZPV0BMVcCi21GSPv
gh5s0YV0fdNFWU9eWTLJW1Lx7MIE+n7Ya4PdqkpbqNLC3LvI06ff0NQSDkzl8quW
q6k2WnIEI4SM+yLmzHkyt5bELhBZgW7hFooMjRcdwCVGGk1XO64YpLHqe+dmen7J
7/RDorFZsYfuR5vOHUs6RZCie1R300/f+4uCqKi/7qEO/I+oeRnCkuLlnREgkc0T
FYUcCSESAzTDUev4HsVPRle1aqjHl06bPcK/yXUIsU6AfBN38K0OxZFHTrjWavpm
PWK1seqnAcTH0K1p4sS3lUkUfmcUR2UCijIKin8q8Ut02+4e5mrkeFS8ixJCxfPf
rWcBVjJBwOj+4Ix505iNPlvX5KDpthLkiqbdACe+sAUS2UPQIsHXfZiqlbW+GayB
9HSqaHlNwZ5sJ/ju8sDa4ARpbpz6ri+KHkQei5kmZBtbnbpILkOOHbujjJCsDSxg
uawah35hqgtK7EEeuNwPKgNZs8XZhjTEzCTffB5hYA/zWphYYmH/51MfrxttvAW/
0W8AiWIZgmuEbUag8Fu2Df90VS8iqoOHvxoC4+H9SeTVKooPxKBv++fMuQv8xse9
lcg3pyzZzbc5CBgbG8r+LGVH/9LwpVi8vai7x0VvaRHN7jLpT2JzCmYe0Ehtef3P
GldQEwddEaTqFbC/oieXCiSrOgHLp07rEz08ETmAyMNeOr+zE/Mx2lRY/02jgqtc
QwMTa0hrFmsONba6Kk4czS4SpS+8XW8hS81xuf+j58ctfNp5DS3ABd8s7F1TL+4N
6OXaWlf66Z/cu8dqO+uF2/cjzx+RrTJM8OMSnO4ygkv/H3ZTmO51CZiDCadWWXGC
Uj9Jcfy0GU5d8FgXQPPRsTb37i8Dmoy5AMavWyFD6sbbU/Pdg1FRvkSU4tm2C7MT
ygAHmvJG0gnKTr1IhcxLmq6KVTpTbHvykYBqUmopUzDUdh06tEVw0MJulo6swt23
RgVUyOaAj7s3IbQvnyG91+2GP+7JwTLurMJPD83FL6lok0xO5sQCu/R2oNB/cp/y
fATEwTOSfm6dsdyVbIttkhA6TTsPjCwDEbRbOSmtcI++B8P13NLYKr4F+SP+S26Y
oZVUs/7AapPqildnBLkoUEpRbZX+nKo/ysTdQWitNr0bgyrZtVtIF0ILrJ59TEaA
GGidSB5ezFdEbTWD+e1vWYDgGgrtPjSw+gg+UGg3wj4SW7BFqT9GLsJJdqBxL2/B
Y7j2OKapYCHpwUJ6qt6zrL43S5wIcNuLZP6s9bU7H7V+DrMaKeE7EMYcc9ZDPf8r
1xXIpp8qQ6Mu+YoIVouqE6iZQMuFU83Hmd+8V64TscBoKQ4Oj7gN975ie+LaUmbZ
1vfODn3CZmKIGoEpiRQthyMw9f1b/byVLx+zmxg1HID0h7mMMVYr8JWWpeeemfgI
UhjUiQC2pyV/nzBVsyPvpANfnwVhgFyDTwaCFMqkSXayDO9mIRy/LnqzS29NDsOw
u/A53l1S/PGBthowRd7IEQN8DJuftKcgkzbOSphDuQu9JnGLKwriMKDElzkH03JH
3fZIRmV1y1eSCOUChAk+Ace3SFe7xVGcYpecOA5J68V23L0yp4ajAjoiKWRxpTFQ
jlpweJLYlS9pqrimdPGh+7bArY9FKpDFFQf9l1gF5sKheE7hLOKptJvbUBZaIc6M
9d/zt7eABHN6YKrEeclPjTTEGb/BlXK75I0MN9iNNirL+j2GCQ33Q3X8+9I4hmo1
l/NFruvB6xfOy7rIFrP4dSlSJYATM21TnQKCZbo/WZgDBDHqdLXQITIUE3qleEP8
JQ59HjXpFp5VCMZ+PCWBBEuvN8m6DxcEoVmRqH2HGqizqu1HQPrcEFXFGywoPv3O
wzudlV+nL6knCrUwbPb/X1OfeLJ3EIP1ot4LamBoqd+G7FK616cQaDQrU7gWLWGf
vlc3X4sDmZMN6ZOPfF1QsmsYnGEltrKwGNNx5KdslQvrXQvwF1SSKb+11mM6hs2Z
oTVS1OTOMmyGdOv6lpDXMzLZZJm0c1CrO9/PGkYUWjGLdUB6BvQJAwRqRQ2zW4/P
h8SIp2OD03KLvojFuO8QsRcVSpvLBOZBM7B7ssJGugPp/SEmmL2ZdBVwh7gxs6Ox
eMhjye6K4f9P9+1lZxHCPJ6WcFeaVawnvQqOHhK7RqZS99f6FIyUP6f5PV3TstOa
x/MrjbA2Zp9OaHI2Kki670a0pk2VKjmm+QX2MuvMqpJa8ifiXvARYI55qibQvq1V
Q3lXl4s1OFxPQ2ubyHvtfrSucmGGIKPxdzx/d6do0zaPFhktbGyj0zHFkiCeYRn/
0IORocuQOgET4sftxqqvQcfrnZ1z1+hH3M/U9wrq8eq49xbQOb8oa6DOK59Uybv1
Tfy07s3ddkduQxwYv3QIKVf0t8LRElpw7MEyq9RoYMahg8K+rYVh8VgfSF613u1l
LyjQDQF8KFCp1JL74ruc5/Xk7SHl24hupbk8tn6GR3AP15C0fR6HRhUvyGY4+Rj3
+fCFT9kHYsQakHF4766YjlQRImpOvwuPnBvChRpT8l60U1eg48STq1FAUUjk1rhg
RXpe8RTedeHX7kkx9SJnSDI2ptK3fMNaJQbtWAPcUHXJk/ZVvkzmb4VNUSMpA8i2
05zxfLkpY4wbvtm43Cp0k6mwkdQAB/tDL9C1KVnVWfICEYA5DwOqsfWES0HxIWNQ
dvEQArw6dyoARxiqtuhcqJA1JdTnqCaH5oO45Oiob83Bw4w7GBk7k9teFVzwXeEI
4AWOqIO8D5t8IU53Qv2UuMN/RyMShovKlwD9aJXMKOM8eXQk9Ur1gAbFDAGbWfNh
KxrPARsvWPvE2N2WHKfxxqlV+ZL2+DTzEuRLfRmseMHOOtR9qCPz5OGJpTMGhCMy
iHCmh5DsLPIxezECwM9QwJayZGWKurR+Yat65yPWtSKL3NO3UvCNSQtFGL+fCko+
wu0XL1MO3VcF6573n5VtfCw0VbQbT/ZddmFtRn6i1BxCArM8W/jYjFa1D64Bi5vG
aM/moeie4heYi0W9q10CxrI/ZH8So4w53XVbgsMJ5EdPK/7GeEucnMkc5iKnw+2i
j8ug7TwdS3azDpf/Y8NPT+jL7NvbGhSrSd1FnLv9KyzkdlrliQPLT0/9YTJAFpMK
57XVaPguH2oNA/34BRs7ZJAJ8dcq+Rj3h2dKQXyBT4ZibJhY8MPOGP8RCcCufWee
2cY4a7ZAu0Ws24EA0+FGBFMc5YLwBFpWFcukU0dXzaeXWB7Vc1Y20F4iW+6+8qQV
ZOQ1TnJjtGJ0jRppe2oau2wePOg4civSXUvD6/U43tZXyiFasiUVxRpSXHmm1xJm
R+/x+OvwREI7wphClfEI1Cvho6V2I2HZjAJGrUqn5RrukxU20xs8nZBmdPTE9FMP
dnjtpNJq1YnsuajyIM0bx9JbFOF1Uxy6ygBuRpveR5z2dFWfaHqUhjKkCTg/JAwQ
tJ4kYvIZ+k0mVPaGJ0/Fy/krz9O1XY2yo/zWrxt7xSwfuaXLFn0HaIMJtJV9JRum
7FQoScfaTdb+K4O0XjQxwS71AGZAhNe6pimWCmvt+5FxcZRCyllKr4joZ4B5s9vI
S/6ICvsxaco3eSlja3aixPX5Ug2Hm1fylbRXWV9EhWFQ+Xp3CbgMqrDm0RKC1sFc
P0bC1YxeZ/dL3oTsEAVm2QtQbW0ZeU/PXpaX9pjBX5K21Bm/tKySM1AlliMkn5tl
1UEevC29RTZafpXs7kwVzIrWFDTpBbCTl1XjiSyxkXqE1pnXNf3NAqBHm8E09OFh
fszv9wG1B8qwH377stKGQOuNFjENqdDjym+emL7iFuuGQxFPKp/zpNRxJT7qQNTx
kOkxKciNTMHKtEmI5bPw6zpdt+BA6ybksd0LfTGcNWOdWarSW69X8G6GwO8DpJBc
MxowZ4juFLKk5s+xZGLYdrKcjExL2NZIISluIiJJXU3ZVPj8g5nvTCG7ioOzV+N0
dORitti/7JZGwiDf2euex5dw+xlvWjnaTtt0WahtqXz638TYKzjhlOky9oHdk/Gm
YtzWZHDd2jPhBkj5vJMK/6Ks1ppe57PEDA0LI6BzQrkQf1eH/8w63Xhg0JPiqnjY
794+aJ4hDYpFzfIGRFeA7ARQFK+dGNZzkx20qC0k9bTSKsU0XLreRw83h4CG794y
0EqHE8L2SuThHhMmjGTGrBloJSamsveuZvY5Dq6D9qOJ7ZJOpdyIxBdHejE3zCv2
CLwMKf/KhXf6h+HQssMgx6v8qe7kLBf0/nPANrYOhNmoCSgt0YPSrT8YYqukObL3
rBZtfIkiRLW6occj/jJHCGSAU2K0GtE4zSj5KatSy9qN0KkjUDi9yhaIuoqF6bVU
iGdHQRZqY20QROUOuOnzoUP+rqfxXG/ZNKwlaUxawSh7qObIVVXGniWpLszAW9fF
+BFul2lmHSwr5trkVbPWpoxr4ZfBXfOLQg/XImz4DwhJyqeT7BzBax5n/jUOGUbW
TuAXV0lX00ZQiFPnA9l4j7JMbh5YlWOnPkiVS622JMa19XPk9xa0Vz9twm+XDSaX
X0BlRHxbS619MN+hkjtL3QytuTc/J7ijlv/P5PRH1n0LxERn/9PUm1rYKRtNzgdR
pReaKDUXNqJXLqXuJbP3hkEcZ6Z8GctxitF69QLG2UevPUm010TdVmMVJ9Z6Wpba
2j5w1WGdGhueUqJAoomLtt35fR79Ouz3rOPsJIrCdptC19YkCS65X8HaL1qjcfao
IxcWe3kgy2JduFCMU511ZjTBe1EJeuIbZjS5zs/GyPH23b/YE/Jbc/68BbTS3eww
eQQYvqjQkxWc7yEJ0QYUnm3bcck61EiO5hjdj66Cm/ycKpwE5mD7H0FN+WSqbQBx
+yRY9RFqWEqa/NVpyEcpGlWwoN+O+qcLESjXJva0wS9/9JBVWDo66e+rdWT6D67x
dTGaFvGf1FZ0f4dZYYtztZ/qWX5nUBqCiBTtIp5KVA93C/McsYK2kVKZOtWhfzix
1mgamBQX12tfbu3JZvhVcDnQv+wGQqNn43BwfAByKtGIiYZUkeifUsz+jnhIw9ZN
gzLNVsTyPU/mMUVW3awZxk3CHSLHHxXb0mGIZB9n3/nSLWFvzIDVQP6hexbpHGqu
Mi052mYNtqYsqKG2L4SzMurwIa4HGu7O2HX/gK97onZCCi/K1+LdglsmxIKXNlil
cF7kS38wGTt9zbRn7BuTKIbilgx9PXSIFJXQckFom543Z0xBq3uNHmp4Apca1yXJ
0Fzs28CP1JoNISLo0icKAjeVu3bPGl0Mf88cz70vHdS37YIwd6/jIQGmOgV7CibW
pdO3WOaJ2X2oLCmIn5Jh3ZQTRToVwSWVJDs6sXE0pTxuWrzAWA9E5W9rK2P/K3Mr
rLzaHDws8exPgpOy7vD4gsL1yGi6asytuMI60JgVfh/7/Wkjut/tqSd9p71/BwuP
eC+f6nKkbnzgl+zeCAdg3xl0WEgUNl2ozXxCMEJYgxp94xgaHnliVeaI6fQCox5Z
AQRk0h4AdpNvkCaerVIA24Ojym4sj+RHznwBgq5x+qwfNP75ExL/W05rD55cVo0T
2qSyvzuQso3d+/SLiniNA5LVsCq7QYzdvDy8YfxfRgMYqUwDgSn73ZSisd2xQ+5z
YoHiiUf/9ORb2tyy0It8jAMVK/YdTmowi0epZzAELmGA6ruwM+VLgjlVwHE/ZCEp
luStaBKb//fgLu435ynl6835W9xlyLb9O9alk/55Pd1oS64X5QBuXtibmVE2vbxH
bifjqgWiVOZx0Rd2p9g+vv51xNeDHevEuqgLG/c+6AWKBtlZVisUpfgSH8bIKfWb
8rDDd1QuOkID6/tu3EYRaNzIpiuDqCQqaPf6hSYQweXGd8P5a4VTdIWxWNEjT6oW
9EKAsaXsyXO0w7JIstFBsoh1LGea9Nn7ZaQKJ7BlhXvTT43OJ0aa1oKdzsQRRVAC
0PaGeF3R3E3zHh3jYkVbilJz81eIEi+msPpsGWR2ucwpMx9ZwsoBSVbX+MtfKX88
f8SewgFmgd2paLKaOgBhk5WCJYle7t6PXY6kzGolrN/KTvm8GpNQjnh3qZQEMxdt
BkPepzvTF08sw8UfLZ0TIZmgophavO1n8fiig9yE9RHG+VQDenYisAOm/bF2BEUn
IdqOhu0h275BAwSAMtJ67kKMurU8K+BimFub1oeruE80u0fFR5M1ia6iaVtcKxCJ
ZX/wSy0YeFS5IqpEvRu8eXlT32HhwpmW0hRSvYEXLp97BE6fENn3o1kvbsfEw/Jj
SD5KtmhKoQ1udov55h1db0YRsRfApyerIml/UDrbzmMBqGguIyjAMtZEf0+6Yhy/
h6YqNMtwF/rgS/sdNyGo5y2jzEWx6gnk6CJZ2gunp7r4tPQ9jPdL9pjC62ZQgd4j
cvz6ESYU5pfaApjtwamRI/fEt9v6krOMjaK94Rs0QhlPr7xS3u8el9cy2E9eupgm
vuLPWdVgkRtytbFt2ljeRZVtSavPOpOZGevgQFj4QH+4C7zWP3A1I4oBMRIeT0XL
Bdgla6hKboB1jM2pZPsHqoo+hygo4094GB1GyossN/10BTqnliVbaLp/zBM8odLI
gYH9r4DE2xq1PbuikfQts6wrOPZxs/0FKL60u3YyvhjB0hErYoiciWnSyuCvvSMJ
gd1if29T26hfLYynslLLjPCg68zUrVYNPw7IKdDAjnPV3ZAD5XE7koyrpYEmIK7Y
mwqEVVq1dk+Lxbkkz5oVCo7sXLSkAURXLeAD31cUlmH9CxxUU7M8PMvhfib5z+FJ
1lkpq4ERPxS7wuoASdUu52tFEHVCMjyBmCEmUi77A+WV1P9lkkcMrPmqJSGBCTk0
d2oWlMeMmSMaB6/Sqsf9MBvWW3+OKsEFZDDIyCXqKoqKPU4eM9FU+IP18ekUauR9
eCDCwTscfBWL46hlgwy9j7JfxyhO9fsec6TETSYq3KMl5w83r49MWdDUyAuFt0jc
mlN0swXvPd8EIfY5sxwCSg2r89b3VUWP9vIv/WxoElebJ0Qi7/AhQLF3we+q67F2
M0u/0uk29+6fQVHi+czfHOGxIJYQtVfpQ3gwrh9T2fbtKu1DNNGmITRt9kQqR0ra
Dtv6ndSaiTSdaVMj0bfrep3pYgjSJTyzhCp7DwWw8M7tlw3/cp/KIsuOa6K1iPKC
4uAU1+RSaRTJnXpiZb/8Su2PXMmDX0BM4XDs9oDd1Wto5ZbjhKrEOA4NtadKgHLK
7oRsMbsj7sUuCTf9rJvwg+b9FbIMhgSBSw5RuxLz2vLDi8UgaJZCVlZ9sE40Hgt8
8lHH9v2BfcYFOm5VWKzIQSvq+wNsp5tJb3sUq70RJq6UJKUBDIxFraxZLo52yyQN
Fyiq54G++u4M67xn/exM+e6lDNaeP2MFzwuf5Px8OGRaFrPpVVNdlM3IjKZyLBuP
veru7+JxgmMhbAmqtMw24PYWw1HPNQgEiKHnttxMzbkV+6ASV1Yr43lP4Mi0peIq
UYSPW+qGubCqlVtHDLDZLpzNUUOybC0SCUHaTXO9vqqZ3lerXc5h1phX4BNHXgxL
/8FbN2qIYBZVKlkNsn9chGcsUFUdgFP3DwT0rjOcGPcXiZ7BhTtrpeyGIMa11I3q
ID9hSLrJZg9pf6zQmSBndTAXlSJMyUsv311soYcKFrfUFuR6tvt8ogynytM9x2UN
AE5x6pz94h8fUPYCu05G2ejB5ginDD+mikPkmYSVXVaOjnP9Ha2j9r6lJMGNM/dn
Cy7BLbAqg2++UKDQIbIkmazkxQZVn8MouCvEVNcgkSyW8xGmZnyX9PMRR1OzPdT2
wUJ67D3s6j4Vxcu0cmAWeyS0B4JoeHgSIrnq6bEhVp2ZFZXha2OH7SzwMc3wg7lI
BQkXYWNe4BvCSrsSePGHy6bpilF9+LAGhoQIS93tQCL5O+XCZBqTYXsoWD6XVGkK
JyYJuor1Imn6n2FGF++/EgLh0xyH3xGpIVjgWfBeVL4vV4xDNos+x8IK98aba2oJ
91gugcu/BtUxPP0kKYtVCJtMKddERQwl8oQUIbmcG+BP0hLU+NHQjxHKAo0QHgsu
dquWN/ssyz+tZyjXiPfltWdox8q5kNnyFQ+WXhqcvzfxwKyL4Uy0LxQoERzt0j8/
lBDzRSUZYviWVkRa0D843SQ5lxD/Yrv/x4R1GBr+nQ59OBfx7gFDqUs3l3/kblm9
vD6eZfH3U6GqRJehg8iu9yQ43swGTXwi/Jhce4zuawumGmD5RrFUlLGAqKJMP2kn
jVBE8rZOYuTxjBy+DAT5EKUDh2kv+1HudtBRZ954cq1fD1yWNCpuHG7z/Wq21UC+
YtLjcyot1bRHtUQPu/aSAVO2mCM3yIVV29gVmG/XVXKNIRk+ixuUmgn7q+tjI0x7
NiEmtfJWX0wdUD41FXOTpnV322S2+5ehGx6i1gw6uQRoRgPeaJw9p/LPsRogBVJa
2tYetyUgJPhDBd3wY5+n8mhlgsXkJm7DNy0Aa6+3fJreNptqdyeCmvtkSj/bwZpq
hoRHHnM510lDad0QBd7DYRABq1WgNWRKejvDLVDnaRnx7NNpleXfAqT7lp1lT6IS
DfaiGgM7P2WLO5NJaOsgz4Iiq17C1ve/t+oQOdXmHI+klWMRE/99N5UW2vTH0DnQ
TvhkQuSYhH4xUiVG3+JTC3QfqaFBev5KkoQD5VWBwpzVsD7LZY7IzVdW8y8frgVz
5adrCk+0+cZjssGqxUMoPQWwSaptsj/MU5Yf0PFGkIBtN9BPT9mE3iOESLlhOGwJ
r3BUrkf5H37XlCIEYQcEUack0/dLIFHr99KTTI07q7poMCp6Cq24YOMURY1BitVU
SSMK610VBoMeY0HHDYC7Di9n6F5317bXdVi4qpUSgfbNuYX0qD2l2zvq5wMP1rE5
8ClDi8vvbM+cILRUvVHz/2/3W5sg/GNt+Xzd+RpPeVeq4G3TTX53d7afrnobTqhT
Fof0bpRdQlfsCWL5G86cN2cUnZn+590m5EzLtqA1oWR5/OD9vBRNQKcTbaV74vtZ
CSRgVSmBwAE+PPT0AUthihGFZOEgchdHQyu13tTp/ybZNHMzjSkO2uaX9DQRNudp
YG7ApUqSswMquSVN8FGTAajl2mV7rn2+yrT4EgfC2dekpi4KQIFqZiKqJt/86iZV
oGqFbYdzpqY2wGZJGmUMSLz5bTfN9FNb17szUplqNr0nVAktPGCtccqTEy3CpeBt
DTZLzebGWkT7G9P0TggBT5KvNgUE5miycen0fx7vZRs3FIyTjC0v5Ko8ujgqxl6C
34LJW6Gkuu024veW2hFr9FqepPHgYfxPLHOuBVHyPx9b7Lcjh4FlS4H2EjYjpKXz
AQ8bGAnqbI4SDIlWc8SFBhZtN1yMut1FZVtDyovRt+AcsH2jkRbLVvpp7LsXn0vZ
cbX52nSEqAYs4T1xYOZmDSrqucY1ONkNsKrBT1Ou+ZcqfJRKSau7kRrQxUCzo/ZM
Lh5+/N/Neax3dRE4CECoCd6P6HWGWXpz7P9FvvH7Qer5XGWwm47W8e9cqLKGKEAd
cwT5/jUXzzEfSNigT026V3ilXsQe50h0/TImnuM8k7W8eDNvEkJWPWfdc/OhbYq5
V5jgYlzGJkxguM+f45Lt/WsYWDj2OGSwYKAH2x4QF5amFz67PwZ4W951Ea5G1ld5
ADLYz+f0qy77+n8AKTWk8zjG8BQBjagcyIPw8hvHGJlcIpKjQOgHeNOgVUlupcKc
iiu8ApyH1eaj2z6tJDKyT5y3/1sZV1uQPzxVmZx56eb8mOw6pdJuzFZAAIcG5oYd
PAhW74SNwQlmwFz3B7hc+6GQUaceOKZ/MVeLInCLFf/Pc3fyKsjVvIWn+Bu3BbSj
dLpedRR+8C2q2y0jB8DvC0kZTVvK4mITAP7yccC2iGZFGe25aBlFG7xHsGWUBmEP
ZvgCYSwUpg07dWxfSOOJ3iva8Sah5imr1jQModBR919xBDHwaSij7z8JsBsCOHTH
pLhbKNd9BFWm7krlco8bqLnHRhMxz37rm6f1hISw+kA1mQBygqHlQUxmDUXZ5Dj0
XD2T/tpA4AnFYpXEuOc0rYr5pltqaeWMuhXtLtnKz0kTrratxlOBIj1D/beDq7YJ
CBtTJrNle2tvCwPOyP1BflhxgiWzuYYkjE9hf3MtlYTYXaV08y786Az13cl269T1
bpTIfpSYxJ2AhaqIC1KXSOebGQDlJInrAwC56V9lHrC1MPK21KD83NbefzGCpfhf
E6aFZ51vQQe8GWDQlZXaWDkTqRDFHivB+bsQqq9cB8CGbbqm6ssKxdKTFo4Xx+dI
AV2D4g4jm5iNCgPH7k4RL9cZMBvxlnL1Ye+pdhblBSUI2PeFQVR0xQE2XhPcF30p
F1B9+qCpITqMlYamro6EfYc71IsiWw/ftvUPcfacykkhkU8G9QLb1jpxs/pBJUB+
sWa25ICi1cGM+JNURcmeF9JmoaquTWKf/b7AQ4jdyeE4neRLQYLCQlZ4ATaGBXup
O+kjeZvg/C1tFZ6vxIKWxDx/J7xPdwwlPMDXUNGbmpjLbja1mIBGb8jbxnYP7wAs
C85ylhMpC7ONIaJPoPfjW/5vQpjC/NiAo6WZBsIsNqnFX0E2NGzTq/ViYXn0BUCL
R7kXrq60nunzcovAXUY1wek/qeVQqyACj+bL6JpMQDkTTWqGW8jnD7QFQq1pIbGI
PvW6/uoGGDD3VjC05+jc5hm0+g7InbmOT4fnGuSAcKTxTmatQskhvq6g/kit0Ztz
RvVokyxdieX57F6dmpL4ZrI74ZQ2gNww2KdC9Pc7luCSMM1lbv93mYp24Dnr0jtl
L78fddCeIYw2LpY1cE/qFv4vF2ac3YYBDRFt4gy/vceP+VFjP5Uz+8PKyW7tQbem
3dkOCcWJ+PmQliPa4uvsrTh1r4Z65en4b/hEVZ/q8x4yHEOeEWHYLQH4urEy2RIZ
u7QVc88wH5uWzZm+IfxcfRigNZVXBPTloH7omTpwOZ3lNq0psn073Bu90HP3l69r
p8PDxuQnaP+SiVEASFVGt4wO6IEXb8+Eh+aMb/YilBH51L+Aa0oah9fpORM4EWkx
k7v0sxJp2pw6HX3hlJNWrWry6uqA47lSU7w9J8XKMATFZCyulFzkIGPtQc2GM0k/
XyrdeusQHk0uBz8Pk/mP4CL56wauSG5E2/08n5tMGo++Uu2xc8RRRj0eVrm4H2X5
yHJpKbDKMkYqjCnHP8s3w/Dyzh/0Qqx8TIoVHldkIgb73UaJ3QPasHzr+kEJTWYz
Q9rpTje2teExJzCVcXTSQdjQuckLyNpFUZknzJ2VxREAbzZAdH1TKRxn25wo61WO
Mcajj0qajnNlxjcbx/ry6P0JwUDXZE9JamgQQvUE2OiXboki+wxKIERhLm9o3kv6
CRl5ijCg0rpXA7Xa7YqZb0wwUibm+pqOkzpGkm9DvdXftAk+S15pWJ0nTQ5XPZVS
AVMbBx5P66ybd+yAWxUTnruTLiB/pLtw8G5ZFpnvzbfy5mK9xAN03OriQqn1WCUa
1L6mRd9JzGuHasyrsJpeNXY3Ti1GcE9oyYWJE7T9cXXrdO6sniwv1nf0Skf9/lIQ
NLlWnqwyQJNvB9NIozVfRivJCawJ7cK3wmJNmrigXp03ZRtFwRsDe2Fm6LP5KPSD
C2e0nkYeVTk7hgYyVgQKqUl3auEaw5VAgWUew6LLpPLwKOYjFZvUrR40PbA9YeNn
EFnZQF40mjAxRhNjXnmnJIqEP6lYjHpMkrypMrL+NaeoFcNxDu9qWyUe9MUTRLt4
lZHj/lNR+zZAlTK340d7V8YZ2FRvWyhOJz80536FYbvaC8DGsMvpDp5HgvhJlyG2
GScXFrgPWOhbr8QKg8zbrBFdFLuQBgtFp8rihezALkUVrZ1Mg2OROQsKFuXcYaqC
T0q2q6TvLmwIFZYTmVeLMk/kTPItjbmu5pPGil77qNIzefaivsafAQ7cO8D7IZlf
R8OIIAH2NoNW7DLulc2TZlSq3mmekEetV9Inv/FgJRGft+p+jfboT97cpZ9up0Mx
Yzf+w0k1w5gGlr/Vb+WiiKfYxRJKm2J/EKhmc4ARyQx8DqF826ZmnqMp2WJ/BFmL
ixjSfdI5YBjFWOYaSZZv0Vj4wW+/XAl0Ztu5mJKR+i+ne1K0781oeVfca+QhE3nu
hBPEUGKTrwEakTl0BzbDrhonoHvMTZgkcQNG9x+/7/jxRf/EYqCO3/gJCoBBl7gF
AbQdWDffKeAFBitl9eE7wSb/0pAb1zSd4+bzfXHrWMxA4FJaxa8aR+PMk5AmC46n
qsclrkZpt4nTl3yW/gwJ5SfOCBMGmxugRi25GM0og7fLn2bQzGY9y//QmKtys5au
WYIw8KZylBNHzy7gfXSc/HIJrKQJitYsbn921AxBxQWGQZFuEmHkn3NZUv5eYYxN
TuXj86MofS+SW9QocQppEF5VcbIFp7QASxvdYAKrufryd/8fOJ45BLsn1gbBBtSg
03QnqMyoVYpf18Nv2J1QZv0WvfxCOf8j9grvWnHefkck/GhUk2sly/l+stZN1YgB
Ts7K36DgEiqg08tUh7cn2NBhY/B2omk58O4x7G6Yh+eQevDKnpXDcQ9wN+ICR/IB
jS24STVPs+JvI6aN8NDehGtAxrIPzJRGPG/8kvhR2Fi8oIy+ttgPD/OhoAm24dMS
9ZgrMEzw9LFjlhw8nstjvGPusC5hOYmOpFZoyb4b0hBrNUtlQ8Vg+UMmEqb9IxBq
wYpG1ExlS0s5AlDRcQyJuqx02BVCBqmP2BU6e3Cbrj5aoKJbUnwYH9IwpB8XUz4i
1cc17LuHbjCPkJzcrjdV5mppcLm7rBnZel2aKEcsYddzeux+rp8gMfmAy4Frw47F
vCBTdCGdhJgJko07YN2+dsXB2G9gAXtTdHtJJCLVc4+tZuNrgL1QZiNgiaFWNueM
jdfsfR0QA8+veW1mZVvswNnwi2kll7M92u7SsnXzx6eEcmMnXq3FahVxQYXfX5GJ
PxYzl49ACY1wWbcMVW6f72WpWq4iLemCwqq3g/34YTGqs2VewcmS4TxGSQWrFepu
2UQ0GrvNHRc7nZogJaAEHi3A2bVN0M8Zxf2IyM6a6RSuFEXaFBRRQ2rv7n7W5LEi
qOpb0PEdvPtkiIvqlLc4EIqOHEbtg8YzltZCZ+plzCshzoawJWP8k54FienjMGQ3
1fq7Zj1LB08bcyOOudiUZvWiEBAYAj3J+iOkxziNYcxDuGCK2/k7zhP8p4/uUmYu
pTnqYBGeJFhepvTOU32rLahd9neGkwq2fpyBMg3gvKq5DSgFJcEKUsQ3uU6EG4p3
uDKvFjE2mwDC8Vp/X+dxyUgWECNEl8T48mTo+QCNJrqlxrWaqPm+Ig+I41KJnfPv
G5XnJUVWAfohEVHEWYnrnMVLEPGdLaRmfxlMrmqJl7tLFy9IhJolJIwMymZOaWQb
tSshvcX4m+xFtk2Ky9AVLwJibdZrMPeb2UO3HNE7sxyve/zOkP8Yy/TrwjOBIBxU
xH0dANi1xYspAqGOwyYdW/RA3eiPX0sMKekHmgk6scgUiERC44Z5T911vyX+/8GJ
fNzmPT5psi/sjU/AnEG4y2BnPiiOOG6D47/LjAu+z8Pc5zK3uq2htxNLybbQq6on
84bFgtcBIJRQQhI4fiHElclikQPGB5pOKXVYCMjZQn2auL/J5Ra4h2hjPHo1dQKN
ZW0pLg3odIcQdpSZG5x3Sv/y5jGZHGGaaLHRGCQQetyL5QPdb8o3iymg93wTGHl5
Bg0LAhz+1PZcO5S6FABxKp6ijOCeLjlZ/ZzuMCcbECOeN+aZ/rlCqpFc8K9dWh84
Y1++4YdgpVqF/9VMopsforZ1ik4Dcly7qwpLkc8ddSRpkwHmUM1qq8Kx6g17Pw1d
4Lfd/JQ/0CM0UVA2yzf3Lj7/NZHOvI2USWEo8hedV+0bPM4N1CGmg6YgzEqAFKuC
vtTYWsd0WqbgjDgMilFx5YZhvcQY39I3JOr2IX4HnU+j2N8cjaQtV9LdyuLTKKd7
bHrZzB2lX7LMd8n/QT3acVyc5W/vCHTP+jBbEtolv1BXtqsD85L25wIlRhIFuCbg
SlTql8eD5TWoE1Jper+sJs1iRsOdDFrV9EVzrhp8jpqSoHE6YJ5tX0LU/7SXQpEJ
ZCf7eBrTyZLt4uQ2uYOljqm+0MeFq6uskeAmROr+SVL2k59he5hpQtVb0ojvFJKd
EZ08ZTgB1QHGYKx/KsUjwRVMg7PCb5iKcN6SFeTyRCg0VVxHUoGt04Zlrhmw3Bk/
/tul6Gc0GJLYrhya+uc0r/fzW/NjuN0K86C8ZSn5wKM2ey1ONTVZyZrgHU1+JWgN
iB5o4lg/fMuFNryjUOkwWKkxuG99JoIotyjFNpb5HNCo6nuv72shjFpnklABWmOg
zcAuye+p6Ga/8NtfcVEvju6YK/g9bFEEOtj9FE0f0TuVWt7wUXAzqzP2TRJbLN08
sniNwfBaAIfvnnmVBBn+c4OKOXxmkKyu9J67Dfy9+zkfSxeYcNpAZkwgoc3QvHKv
i4mBqB/PVNsyNNjPXvqpIdRIqGsddR1cgEBu5+7cJeKw9/+5uNYXims9YfxuQ8Y+
GKbJcE5ENOKjEMHLNLlBf4kqheyKCNeW3/V9rFJ1BDFJG/B0J/H+mCEqUTIjQxfY
Pd4HUaoHSi2KdgOaPxNXV5CFM5xZJaGrvEZLl9yRK6mKN3SYhLAXSPXhCWbj3uhX
Y9fvIgpSAeP0NL2huRMgxGsPoJG5wx6Q0QCdaR5ONpD6Y0knrHAleyiZtoam1ARl
eD/xceatiUGZ+PC+miI5Kmj4NTnuo9EmZxgsifu8C+STB8e7HAkD+QieFsfSQ1rr
qNF8jPxpfyrzubicQRU8At/lhvkOgY3YhgorjTWKM+YyPXMgS9nOpY7GMvKKxxmw
HNBVzPELedoaBEnnQIEq2A7FcKNzlpF/6rqapy8Vy7QuWa8Xd5oTeAlavnJB8pgB
a9nBW1XkGKVxKjGxX1Txvv4dDPB2n/1XazDcILVGQUJ1O285OQU+HXFa98mahk4O
wLbk4VGaQ8G8oFNBpf/m4V5WAbEX9wbsk8BAexs6BhUef5M+vNyOfmjjnlorffZD
HmLfNBnGbuhUcsgLF+wrm1r3RKE7rozoBB22vvzUAHxly8sFzSoR9Y8rTaCMAedR
Dpihy2+eDe1PRQqfzMODhQKHVUiNRfjMTyL9Vzc53gKccpvvkvAG7N5PVYLcNSRF
kYY6bRFCWzVdqnE/l1H8SFzMm97W8a7wNhZCI7V9i+msIbNFCQp9l2Lgp6cFJ+0H
Pdk4mMbK53jmQxWCTYAmzGgJjrP7cfN8EQwzbH/0+W5el5nimXS9mFHUYHjiLxAO
Ce6gcKvaoVrVDRmP9wiXmHx0fiFbFUL/dVgJDOK3+/G/5oyYDnZnAVkMTiVce5xX
g+z7EDOHTUAsMkLMIqAXJQYqoz+8FqY9ON0ZfHmekdU7wdeHCauFiDds6k99OY96
py8fEO2OLcYQIVg5DKSMLVAGGvdJpqA+0LF4gG3i/huM0p382NqhuylNxc3Epr8K
EPl0KHqN5oG0ySJNDTjoblWlpdPHEfl27nKNfutmjRi1vXz5/VdeRn/hHpEuDe52
hCfTQp2anOM5ww/zdPpwF17/MU47Wz5g+mVVr+8Vo7DuwaVAWMrq0uS4XY2jd1kk
DN3oNJh83LRQnAwpx2LHEb1UdZmV1wCkIWr3SQiSwLSxVuCfWAIgyPfywD6Gq2g8
7EvhMgCFgFT0Pw923mUg9pHfIZket1doWGFfoQs4KVBmuF+gEt3CnOu/hA7zcwG2
fi6qF9dEvoOnup9LFHATTcQVjTuH1eTGU3UZQmQdKYOaZLRBa4J8dpUVOCko1FEs
z63xEyfFfh9qvX/sR2qcdXs82Zs/e7K2Wkb8qmlgZOoe3xlZzWMu4VNnNEHR8FuF
qHpcxG2m6s7qiPF+7xpHdylIbGN4lMwMgDRhkwDK7PuDTqerdjGPWfUuk04UV6OY
ZP07QGJq6hu5AzmbkX9cEgGDJbtWB2duhA5RkEp1BA/HBzjuAFLkRAI6Ztm4TRDl
OBXWTCpTZK5lHaNKW301Nva0mdfUF4Aii6dzj1NO6j7OuDSa9atF5AcMOYz5AKyZ
Ql89BWgHcq0dyBa3pMxVfSg/V1WfL1X76ymTjXmc0XaPXU3ddUMi0qsFAQDRrHVH
7QcNpLc3clLL4bmq22GGzNPGYc8lhjMevHxDF91ByouXDAsooU+SyXsa0eQa7e4x
1zul9MiAVm8zGs9R3ztVmjZqOGcWoji7tIxiEA4w2dsp9bvDx6LZbkp+KE88BhA+
zF3YC3U7F5WHxMDSXREFJ82gUjqyD+hQL0N0oUaY+AGG3oo2M1vT+iaHKBbIKoEG
7EPu4OT4W5JWHsxBuqVVrUA5wF/w7OjLD+qxO+j2Is8/kt6e0Y7Jek+j7esjLl09
T6+7enbwW+id1Zug6iv23psN0+M+PIkUrOBNWTsaxiiJgG9a7TwJ84qQ1bmL79H1
jIL+9FU+MuYPeO3UAHtelEj5Y9TqZzAcg4nAsLEpQy0L/AXWNmhknUnnQGgUGDpV
0/78RWC/rEq3CM6wi3JgFe5b3J3Ya351vAUDxrNI/B5E4+XDXMOuh+EvE+VKIEuD
QW0EZ7DbQs+MJ9D92OMcaCvRVXLWXUj0sTH3ewfFjQgtE3Nn8eGM44HQyjHrGddK
QS0gnHe71rYJUXQRl9u3jdvuJa9kFp0d+3OG3ELGJXu7ndLOGtzx3uRlfoXAq1Qd
2BWytpCcygJQxRusTfqJ2sL5OZ4JxROsD9wy8Tijb3tZKfP2pdzyNGTtZxo2gQU8
7OxHil5VwqV10saPtQJ7xZ7PETSaJKnQKZdv03L5OSFhMbgOg1IYwGt9SJ2rwduH
cpgSa4l4UfgxMaHszEeCxTLcopXSRpL9kut/t2Fo3nZDmoa3rS2bKV0IQroaaonK
fHiIc7LD6cICxQf9wcFU1w9d0um1jptFdIQlOkdVwg6+2brWj7rUymmcLLk0a+D1
8Ez9VXP9zjwxK7n6ZTUhxsptFk7ojxfSpSeoBUTz+zZv+XwlZeO98drxaXCdFwuX
cKzaUPDSHHtlJZ9uNDQn8b+Z6cs5oB9489B24Ya7Ey5uwS+dYAA3DscQKPISLNeI
YhamKYrnZlodR41KG9B6KfmiYJuiVl4d+nlCour5AkDm2m6UX1evwkQ5fNP0RU8X
EqWS1X1bkVkdiltWy9nBkvtW4V83QISMLdFU0jMWzke+Ztx9d+6HGNhjVfFKkMLd
EqJ75qk0aKf4MqI3vyN2MO2Opxi045sqT8nr0LW6KfLLP8SnfjkT3fxgBgN0eMho
DlUPgJuAYAi9KW53STGmwYgIZxG9bg6nu6gxcCRNHcKWGN5MvRnk7DYXDDRstF3u
BztkU6kuDKAC956bZH2oqVnWtsnhRN6a4SZhPNWDJem/PoXJJQUf5UkvmA688m3A
wlXMC3vlYexN2yPX7BTdrxRhBCF7DDA4s7Jd5YXtsGWrK9dzCK44hRejTSOW+Fhk
8tSesOsyrPbRlxfC1q3O3ltUSxpsiGHCyiTUr7/rsB3X0Ux5fJ72aCitHKSmXWYa
yicJxKoDlV0MtRjrqSMMx8mndseCy+oeyMcTg0kfgLJxWS3L3KTJPx7RbGLHvgV9
mnIghbEEH8i5nGl4lo7sVFZUNIcEqupFtLGnKrTLU3MdWjLLYNxuvD/2kzMYUoKY
UNoy8ll8EFSdJuS/SnHCAVcZN4TAU8naOXvQvP6VpLJ1RaoP4cZkbyD0R05O+LQV
PQBPKl3j4Edb9opIzA3IdqZjx2WLCvcVfEgtmmHW8O12fLxfBXJI9yiZ8aJC26Ud
Od1qQFfKbRQf+s3JIu0SjSVjrl2KJ+LT4fvJP5gSwIEeasdHTupCj1jINGcCbUUp
r4zz2qNwHBKUI6VJonka+hqMZeGFkjpkgr6cNJT+v0MTrV1/2uHw/P8ByUdJw3RE
qn4NETVbKmh6vdwiaUydngAz2vyFXsNmJTfPIv3RVQznWesz+8hxhv2ZRfRbsDWX
ZFCP7AaDZN8csK7B8dM1KDQYsfW1eAhsZyFP2e/SNAXIgwJ0uXOhmffWCmviIQBY
wEuJhqQuZNfg5waR+g55wVITfky6A3z1HLysDsCYefDKkZR3sV1sTLeCaBPkuIJ6
ruyNMgddB34rtArzvB4FO3sa6r3yvSK00oLIRZz/B5Lh1Ov3xtlLsAzP02Dq2RVC
payfanWBCaC2XhrH4T2GbODWAoxlaPwxkHosHIJhPXhXZikwL1PYOU+YpuKQJ/x1
uluKwmwkx7jVcSbSUYxnxTRb72uLD42tPPhYmLqPCDhTLpEzvlqDt9J9ZARWWHu+
0XR+3zHofCmWwKVYuZWq3vXSlWY5xoFvXC1Op9wFO6kPqWbjxgYLms7WGPLQrZvH
CgVEqCXPgMworHetyULO1QcCb90b+PxqlpPXfdj+2f/mGVDYUarmt+Hc8yL/qM/I
trszPolL3iKDF0wxi2Zyoq84iUu7aJWuzPJ89lEPSk26R7fYoiJ9i1pJ6Zu5YIpe
LlVUR2RD25fiZ30stY2ONNW5KC7xK4lk7ZF40LDBZxWK+8L2tYLHiEH7NgkMV/u2
/JaSJr2TZTWUea1A7y3/eVGtqIIBkKjdm61fM133cFZfcV52WRhB2+eRZ+H/avcy
BN0DtSRBVHXhOgJhIVNY809p7k1Kp97IzYE9SG4faSCQjBFX7eVCbNkASELXMCvs
KXvzSkaAT3MO9Bay8mBtvO2XYF/IrgmYv0mcS3vaz5e9FNblV4qy6Xexes0bLZM/
3l38ALEn6o4z6zwWi/rQ2fpDHfWyHfvc8OMRfpJWzImjSSv7+TrTdQWtHweNe54r
SL6hIlwuHbR4UZm5vbYj0Ab5HsdeNk0Q0ZS7ubL2UGg9g2rhZvrbhnNMdaMiUrOp
APGxhEIz3OR8ZLqwGMUwe+Kn7bAM+L0jxeNyti82mnhlnXimMUO0bOjM4vr5mMJa
9noOr61gGfzUcykXyPA9vu7CTJvX34yPhDxSpz7FyNHj7zkAgm/m0iHjxQKsE2FS
wvSAK+AsHATL3yxcBe4/EJKjqgjk9GzPpbpq/N6sGYt7up4flfVaaN1nqqRwTpCQ
SuZ8P/SpWeen2AtqJmnacW0OfLS/19ehG2NNre58Borb8y12txGZwbXSRjYNf3z8
Hx6IlkQCorlqYYCAxB5E/7wq8PXqgjBj9R2JvLUXQRTTYFX5kTniO7VROVDwm4Uq
JmOZrgu4JAE/fM1lRVi6v/8iq74bvTLO7N4BzrCiEV0M9JBGL2GHMMfduMQ49ZSc
M3qf8mbiJ+VucC48O5E8FLmzW6ohGmYjLca7tcQFAMR6LxOVJ3qkkDf4VSQr3c2i
6RLJc6jeF7hy/JOy0I8cGUsNqvcC7Qrj9D+iRQTxCrUhDpdWNadcfQawVEMiqBN1
yvcRbLE55XZlKgeW39uqpGk+i9qQMQMvxJgGkUPxDAlGU+6ZcpAsHn9k0uVAYXmp
Jpljl2oNhEwJQfxOWpXZZUMB/TmWzzsLOzHpXth/FcTl1YTMqY2y7oY6clMtXAlu
1/ZqmiETAj8W3FuWHGvMtAVA5m0rHM1U/rH87ikTAHInkqbjqfVypBVCL9ZAJP4g
n8s0X5ejSi6hqAxoGarLcRRDI3JIVTXEzqWDsscD/ME7N21p1Sey2Q8q/ffVsSG3
7pa6Up4FrztTVtQnTMJfPPVSZ9/1eSvxWylwKyqEpiUq+HKazLdq8Okmzc2taLrj
JRowjCanhpM4LekMOgWcEqgD4Mr+yVFJ3bc8fr8FMTrlSoePZuNtDfMINqpiGous
+YF7tvDotEACvN4MUlXtRfwomxnUqtFfzzzrNY8XRRT0kUV3EGr+ieX9vwD8K2Ih
HvJh7gybmpPN9cuhAGFRLwdenqID9cHt2K+uOW0uC2SiHVKwEmthIA0H+P37jK2q
2/TiRh/v2hpSZrs6FT0YcVCRnUqH/wJn6RZ9pEEXWcjW9MgVg9560tRE7xtdjxCE
bcuEGl0g+dlh/5FB/IP4U0HC+yWDLLYIGmZTd3kDXrU8lJV5+CKOur/f/n1/BgZV
nX9pwlvmXaUErvk+Z7m+2XLIX79GFgXCRaA7Oei6BWE21mZ1L8TNkZoCao0TpOBs
wMmsG6GXxeoceZ6CObhFJFufGqD6Jk/d0U+XvzwPxvcbLAugDDU62bgCfTnDgVjd
wT6ErSdGZjoP29QUKueBwpPwK2OP0dgOJgi5zEelHCB38hyZ2AeDvaTG1sFkMjeK
E82srwdjYkcvHg9atQt6hpyoK4VMVllDU+GVfxshAsMK36qdLQ0J4lmmqZYMuIme
txBKX87+64CQlKBBTud9HOgY9AAH2qTpKALP9X0tra8hpZzZzYBb7EkveiS/TQEu
GCVMJOn32xZEFb2Po/UY8TgZeHxZgsOv1JaoePOj1sMr5TaHx8MOquk/pOQ+P/2M
JisOU6qbBTNfoLon6QkjgWFQRj+kT0/T3yPLd8jOQuClEqYLvzRKKPp2xKNRTfCH
vayEadTxjTNuR/ee+BYUPShGePWl0pvMFGSgkJY0AiHXybZtJ+YOOfvH9CVejCHa
+5EH7Fom6GwPfZz8dEixbwSUc2cXOpSgwYrxAW5UBPbbbhxbtwH2W9MsNOC/36di
rrsJOaSYtz3YiZvFVSmZFKO5Ip4mkRH7sGw4r/rKHfZeD8Dmh+Yqtd3V/CC8wa/T
SDu1HBcw0rxwr0/GzBthM8+98aZ84c7fLSkQPNRnOwUnjafmM+dzHf97Eu6aZyO9
ku6mZHyPloOl8xiZPiIITCqY2GkBCfLafLTOq2GXvGWx3k2wDd3885nFIGPtB/5u
T/CA0rPbXSIq+QSiMVmmYUuJz59HDTkQoMvv4wljkIU8FWD5RfYdmtiBHQtcf0X0
u/VWYxEYDqZ6e0KaCqrkv7mr4/tqQNFX/qTyx8ZoQFraLXTGd6euar0RYuAnLtON
QX+SeJ+mvIrxIZq6Lkp4szaRM9X/cBQFagZzSI9LCvR3Fr8bRSMngIM4X88gXeyY
UWGMwgCrgj2snXMJyNLA/PLXA+5p44ozTnoC0Fp71g/LL/Vl28ve+6gdL68xYPZB
ESsqoRMKqvD6cWH23EoR7k6RQVcbSOF07OdSwd0A7kyfHyn82JJyVia5JQ8Mc5qo
T9y4mHWf7bmrZTLBH6ogH0fwSv3xE7p5C0+E4XrdQBUcw5M6W7SXeJqJCWSXCSPV
4j0QkGLU+bxs7gwOrBIK32j26rxSNRZrYQWjBpMxDbr3DG1gsOHL3XSZJUPh0Hj7
34f8J8g+WiVr44tfwXXsvUeonkzIUWB1gijsK09OSN2z9tKmSV07jO/T8KPod2fW
c8MMFoL6pq5GTDoVMA+vjEv1+GDAloq8sIVkUPZ/zU5nvivF8gYTvptfl56i0l3J
2OcDI44j+Kh41GyoSzi8C8NhttNwapN0ADiDHMFAULmc+7GF1M/eYYR7ez5Lh7Hy
tJyBGN7s9wGFS3oZgMT8FXotmlJfJ9vNQkHegeyQ9t0ehJh1SNp4P+dyyJYBMSBT
4/TX3MFA+0sFQcPwVxb14hyHKAQAtEf23FWiPTatqjhUFVWvrk9NiShk+I0MPELB
vsljbQTzPii7LvPFHpC/pFmMDhksBjZo/VsEGsonIklAdjOPbwevQCjuTjofY1z9
UfHm//5NdUnOnlr44rjEXiSYVEdxMnR9cRYXWD9cq6lOMFGObwlEzsjDWw1GDljF
AE03rL425u2/c29+9DerJZEEhMHaJKC2RD2957lkZ5DZ2DmimxnTjtgeb4rC8kuV
TpsmhGUbRohQvyTXCTJydJVAeRGdzeGVHR86FjQk1osTFaKB1nk/cF56+eGxPdP5
YxxsGaRaEFDfdd/c8cR+XJ+PrTwGVmnv7UQ5JCE75O97L4ZHPJBU0z8BOEFGcaTZ
/d0fkF91R4Dyr16JJZrWANJqDNt3HeBaW6avHM/ntx3iYXgRhZHWXrO20DaOfIIm
W301PECIznyggZSnYQNiLZJBkYUELym8h6i6aCCkWyVHCC3kpYmtjsJXBBntnmG+
lVNJ2mQMYSoC+v+ZC3T2WOhBK6z8QK/lNpVXzQoTUYkMZqiJsL/V7eJXBR1tqYpv
WjG4t6TFFyPYx7bVWGAKwGfeb/JD4xYg/exhvDI6+p9cMjoSIU98JwybRyAp6qf9
Bi5i2diauq+CLzTxo4pLhihpik4gW8cEMzcx/usptuh+OtH8xwHrqhEmRrX74tiC
aooEk49+zusT5Gk4MwIQoeY5DOE0HBN9qyDkNQwv3oIsk17h6x21jPkx5v2i4w9S
OWjkkM9zWzB1tVzAsyvAQ5mtzcwADjm0D++RwjCGE0FqBIKYU6XesfptDvxe9IRQ
MkLwmM3veuz9v1Jg6DId8DO8WsmEaZx16YUjk+Mx3QdTd84SMH4Q9eS6ieOel/S9
dJEQ8WSuJ5P7W8DMRzqnPNWIlMPtviKrm1Pc75y5pZiWDqVQuqMMLMwmXKsJcPLq
GMqQjYeXL2xcJRn5Ca0qYBkNhfMGplgSuc9EwThF0bBZGtIXzaWC9VcC846ClzoW
9DSPPgAIqfOF8znE+H1IsndyKeOnbIuKCodkakcIY009ep7+fH2FdLEZGqFw2C5A
ECqySZo/AksoMCkNBguoDgeYKYhLr3tcZr11OjzPt90YLsSV6bZoAzSYKOGm6yqV
UrnSuUnVUchQcw/JTGEP05PhFTm5FnFXUhlS25qn3Gb2hepP3+Xy27UTbLliH2SW
NW4Z9M0nwcZwl3S1Y42gu/acGr5gtf/OfjYa30FbqRHKg2DrdaXKIw5e/qIqfuxd
wuR1k5OVgYnd7QKIxK2JXzsod92MloZv5iKIK8jPWNCXUecmaiGvxmBarY0ko5MI
fX1LPeQ+wBb5+b3ltmRUxtwxBWMmVZKBdNqAsgGyKvnho3ZdB0KRCZoLP8r2gRoF
IUxQSY1B1n1fQnHnvipLYaxqrYXYcQpKLvet9j0ZURWPgVKoObV1espKTdiud1p6
VMjog2KJZafuKLRNc6b5vBEKnfok0hrdV0AL4e8CRdW5bWXOymI91lDmSTS9jJ+A
S2MBY90vL5BXtQUyV3kGKjJAKBRpugN0AHmI4FdeEYaJJ+X7Vx2m/D133sfyHnY1
87oo75qnnkQ9M10cTCouvkgdxY2SlnkY8zOTSbI7zDlzOOHvg8+DlnMCGV9jRGiz
uhat84JBgnBb/ndwwkRwJihPULG87ts8dmmX9i7XPgAsUcZYkiTYmdw2K2n4EJzQ
+L8I53lRsc0wLWzExsnEDAyNz1NQGrGHAo2kgT5prXLLI3HTIkoEGfapRceytc1U
MN13bFY+hvz7P+prKxx9sMAw0w86wGYhRXUT+QENTX1jGFDFxAA7pGMBw979+z9e
2ypVp24CeVtGEFlkagO0vl/wNSpJCoHgewDqmQ+jkKW3CYN/3pVmuHfQF6ju0l6f
daoCjXtM+1Z7paK+lOtawY/c+xqy58jG9bYDBo4NHfsbimj4qYyRjcPjZR0YXZNt
wgQtsvCwmH0d2HiyPoAmNa06CVl1vm0EWNA7QUNJ0VXPKDrB3cWuP2RDhdy1AVYV
F0wXn40BohZ7bwhv0B2Fcoj+AY49RPPfDct6hbR9OTjfEeDrqNI4io/l5grf4epu
+OPvZ5/87Npfz3CAOa+QMqkZN19yr1xAQkK3OrMCCxP0HAli6hnvQclK9AubFUrx
Zy3xRAlHewgwvGzeFBnVxaUdXnI61sV+Q9TyF46zUqUmGiWq89vRokGVJuMHqxZU
dT4yN+UINIyfXuowfoGdsDAry0295LdqLoilvebZpjkAQyc+1zqlW3xrG+Xg2NyJ
lBySDyycNIv5kwZYKlLNFNNA8upkOuUYh99tRkCmBC3qxiXpcHvJgd97L1sRXrlu
U7JCl0uZaItuUhlsrjh1jN/8RE+52j4ef9b1fA6TfvZ5qvKIi4+4vm5hrXSZB8av
07dEn4bWDO4JyUdKZ7e4DFozya4JjRoPWn2G1XUJCfDGrIXJ4gfH9EkGLkMJTK3i
6qBXJs/MaW9AYCl5BOjegT7xzJPst84tOqKLpzyy/aMzfz+ACkeErcJo4nGVM63d
6zp1akQg0ZjFWNS2Fme2z1dSN4uEIjrnJAYEqqYWyFhOP0r2ytr3oo4ueNtEdgfM
3gwCJRCs5GXPFw8PYlrlI/wNsZGY8NeHtSpG6oDv/zG8MzN1p19x//QMfJTD6Ysp
IgI15x8SEHnvc7nWytD2LsV3mkORD+rFiZzyzL5cDTXdZ9HdWnxuP/irj/5U//jK
35XIV/ktpJE+lgwugfQdz4bhcYtEYJKF7nszhaUGEw3Oh++6NzpbHjORndRiJ+CF
QX8G0ljkFEHS8JbIRx+T3WBh3pG9Gf7FkFIsSD2AggMTnaoN9+dFPyTvJ5i2kodf
1yOjR+ETR2YfhP718Z0E7Logig1rCrkPcvn6kGkKDHBSGMFYerM5H/w16A+Pu77n
l5YIOMfZcQ27v5OYNvYII9DrDBu5yevlj5zab8X7iakYBCHcpVZiURCdrXMDZeUE
GXuoiBgYGypj5S3SglgK2/YOdQk3G3o/LNsr33/Hvo+EoZGA5+1ZdWU8SLD+MzhP
QMBukAVK2BjtQXAkHf2pBqYq/B/0rWcfxWdZLJDjeGojDcv/vyXau2zeIVpkndq6
dh/9QjWPLuf9sV2Uwiv1mSvEbkm8ZQzYILx263Zhs+MmI0uI+YDL4lv0bPr1gmr/
VN1y/tC2gqFAtB9mY7nyYdTUzfIAKcKJjhbvLcXjzs722eua7IEHAZNCR8sj+ZDK
s9/DGh5SW1vjBJi6LTgctT0fvnCfuLTOAeJ9wyNyKgRpDFSyW+oB+7i0FeXUb/yX
ztzViZxvVS2Dv1k2yLF8bwtcTfLWefpnHwGF4uEeM1SHUbw85q6flNgf3XCPf4am
3st77fIKZZN0UDgzjDx2R1TQkSe0+k0Wsy8pmd+/Zo0uwBIbvbHQN0VIwqxrZyPA
3D4d1XWVSNDHEmYFpAea34QJUrzlDdwX36ZLOfdJ6Tyn4c4E8VHiYVVIB6sd6Fu1
FS5jMJxTx3QEJWhcQ/cku9eBoEWittqX/9oRkjUTMVurYG4zw4N8GuaUTbOUj8T7
WTikWVKrCLYympgi5SvCTDcHbzaXu0TazjrJ5PC/Apr1X3Rnifohx1K7LF2lVCnb
48FJv1K25IgLxaDQBSNKO7tFCJtDkbO2b4UISOTTApesE+NUKl3O8rpQ9TeBuklU
h+0QXeUUCIBg9iAUT5X2zl9wfWGetd6V83Zf6FkQ9L5LhXiYIRWprP05YTlH6NXf
ihlu6H54ATCxwt5e/22foo5dvSdBXSDIaUUgt40LKZUOeKOX0pS/wp2UB+QKgJop
GPuljYTd+enWLE7RojLU/fDoK3kdWdvAHZcDxiopjty24shnI5AXy8RlUmY7AtWy
XH64v0ZEcHzqfG1j0ffgau7AK+wykNYsk47AwsQGRGnWvVjCa1pavO2LPCUyHSVw
zZpdVe+28kxSjHTIA212ycfCq2lFdJc248rtDTkHSp3iXzK2tuCjLIUcyeAp76uf
REU4reUCcjTx9yt919HoRDQoZo4X5hn99K5x3Dj0M3icbnVeTpenHsD0CMHYvnKu
XQNWNPx1qIQtHc2blo4Ju/9ARq2a6J4rz/SPb7DIEh++n9EmUqnJERSQjt4dXSM0
Y7TDQ/GIiDDwtVZhvUP49KwPMMIUpBgHGlxBaUu+LjiNzU6/PHMxhoelbHB+KNV1
IUfl7ScnpKxmqf4WJWz8E8CdjsTCH2e7MUoc0JRCjRl8MUxlwCbFpRyO1Yx29/P0
Vw7gv7yRQJui6iQ9Ml/xdKQ/vYkBnsmeGMN2IzXiX1A4MGBbIRZr+ChOoT2Zxit6
KcYMuZw4Gj9r3+5YT6GiFeLWscVezZ095G/bMSxxcm5RBIG4OIDFvAqocS7qOLn4
tQ1AtILx68zfpXwJlBKQ85Spdr6+UCxipeI0U0bWBD99KKimrjotyLqceZ4yBwlj
eg7PCTh5MtKpp6urYZDY4v2BMJQkNbfOwVmp1ScoI5VroYj5+H1qFWViuSawiIUv
od+fLs8BPmkfsgwJTyq22XmdFYSV6T/F1gs+j4aQlhp6XPyB3cAByRg89AOElPCc
F5vpsRWnP9LECRKfJPWIrgYT6t2BMeoHJ+nPLDyH4TWSZdVsrMqGM9pCF+IEy15e
UGQkzMHOYf1bOj3RkoSXD79PrWDegmF4bcsf8lRZPxgzaNHOLsYDfbBC7V+a75Vb
TYKY+SmbDnpGQe9Z5JHtQ+zHgsEPKwEBW2B4PLC2w7zKjriUYHYcfIvk3aMDRRtx
AcwtXK1xFjC37zGE1iXItXv0FxGJjbGbQu3+acoVj30k7aKMrnKLbJfwBFcBUoFb
KgdLDVhL6hgJ7wsGxaQoQxFxOEgfaakgeKOCxffMPrIdcDKig4wxcgYZCBS2ezqg
bivy4hsp6R8EtNClaJZO429iCNL39YrSCgr1lKytgfko94bRU2+ujlzqwzyiOm7U
RJ0TfgmmjWf0EeVDwwikFxy2o1VIaqLAprvJPJavopB5822UhztAzsOaA7Bvtk+M
0hcbqAh8F2AAs82I7OtUmCdHdhjsZm4VGknju4quXtpYecKyETgV1bMmyL0nutXe
7QrorOXaunqadf7HNUH+iCoEN2AvEG4UZn76FiqQpBHguqO5Vw/TXTlPcQqRafpS
ORoi0XqCQKd0odBDAaBluhSQYZmi3Wg4eahHF6oymiGoFE/UsqtalvuRU1J75bPi
NfnCVqnYQ2RhajmwxBN+THM4qNXWE8ACiVypIwbV2fGl+SxsV8UPSAmTIdztfzXp
fiRiyzVZlFOnu9eotiQbi9uyJMuQOJz3Ko8UOwtR+TLKXm7zHsXkFUhU1nLU/Uh6
IVQE6JR/0Pb7uzDs3sJTdnGR6PayvTUE0z8qypiXz5CpoJlUt60bnvUExcbmzMSv
8MIIn+hxsoEeMXmhNTTPD8rpshI9nhfk1+XbnkDF5XJTOxZLzGWZWSsJb8SJXTrN
qyumvK0VACEWvrMaUG16wIDk18QFVLZPJw7StJWEAZQd49hMvd2ot35E/pU/BC2s
pehRyJsNLk5+EHjDowO2VQ+TplZocYwjrU81HgqY49e+3UnpsWVzPRk9kBYA2/uC
WLupoye1Uocxuc4/UOP2XtH3Gu8z6Y1vdyWFENvLk3dpCrm4OuS4pfapyU052z/u
qI3M/s8RleBGzo6cXjg7WScF7KKtO95vXP8stLuBmtsH4eoXnl+El2X53tcDmPrj
Oi1SNdYLf8l4yCw4aXq9v7MFrPEQRGrNhsKAnJ7SPZSrhtsHvHY+hDwuc+Sn1QsV
8tpB9RFAv8C+aK8fTzIzs2o5gYrNJcmaHHVvAjRgIucloHTfnYbkjD0xT3oFN81O
cvMFT+ZHM3sxAndxFzhPGCIiG9PNKq45OOvm/3PH6HD/HqPNxzlq35R0dAHLc3yU
wwed8SVQTj34mKK4PDT1Qz1OSNTOa2mC/RFFRhcKyxLdxhCZyk+sCQFL7DaMeTPV
GI5d8yYwaXR6JXrgyNeKqNq4Qgvi3LFyu8/t+s9h2Ee+m0/9gN0PI+61xwQp+cgn
P12UQ9kvUjqXobBmhZWhzfk4CXCe/NY/0kAxt0kRmaN3kAmakrLKRvkdfSnIXkQT
KcJSl64tXFwvyn265km8qLhrHVFRXrThjWNj2OqEHW9FlUDwMuu3TIBKBFwvZ5FX
+Oj2SzB62od/1ge2thvQ3s46+J6SX4HoiM9vatmr28SeQRrcYVoMz2mE4zYzbw/d
Es79ce4SDDxdQA3v0hM9P2GRUyrnTYUwtC+2u+A8LpdyKynXx56PDEFAC6yGly4C
KqV9cjmqdoJv1iis91MajIGmfvL2oM8Cn54WIbxqiDlA7wdw6cs13woV1IjWbGgl
3UWCvxQaN0gqYppjDwYpH8nywv+Sxnfj36XZrqcWyw66HD/Ls2vN8IqJT4NiUXVl
bnxB+ESmS63marS0szVCQiETm1ffPRD17de8JX5zvoxA2PTN1CE5TyC9+0zg1XE/
Dazh84l36KgQLY04TguIZPkuI/3t9+vl2czqA6lv5/n2zwNgJPcaFPMecsLh6R/O
1Mm0qP6wjomg349tnfTet9g6GiE4AKAe7LlIFz7fW1/+M1OWbcomNYktutTMkYU3
cV4gennopsIYdJJcuXOAi7Sa0HeFbJJ9QgB6jApsFYn8qlliJoKT+39tkHz4/m/X
mvI6HY5Rm8GNN3Y3soTmCo6t4kl+v59OFExuwSrrT8p3S72/0kXB/6ngOG+n++x0
mY6S2ob9f0QGTwRA1TgOko+YaqDUIDuoAVrWsAOzhp9RSlbW0cIfeFla4UpRIqOf
jNaSRNFh+PxCJ9qKKJX8x7jGhE2pknwoEEx5wH8Jw+q+tLikLa0CRV8eQ/nur+z5
A/CxEaAiImMOkPANM4I6oRLaaIWnZ32rf0MBTmPd1h0aZ67xW+6YbBjYI/Zqa2MC
wKXYEFyoqgqwRqAilhxlueRpq6Rny4/eMHh/IhQL5sSaNobgJqaVVIPWebkNZrQC
K2Lc4Fxn1rqJPzN7kJtaSRTSlXKmH+IgQ7Vkl+N56OKsUS1pD+cawIU1rlZ80cBI
k0J+EU7Fkk212KyiOFFTxfqKUdeHDoUObEd8sj9F80sE8xsZpTpLf8ROS6PNlscA
mbAQ9ZolE8qziGECf1X68tEKqRYVkE665/Ph0o2NKUvub2YG34ATZ9D+MA+/9tyi
8+cbUmGvES3GXqGuxcKYdYY0AVCj2v6gr1JSDgIZEP5xmXxZ8Cn0ETGrJu0lBUxK
1aq5Xlt2GV4nkDPWEfjEtjAKfdIZXeDjtgwOfbOiyOGJjK6/u2FViLB6w7O1yde3
XlPyvwCuby7tUvt0WJGLU67pFglqFcSEvrJVU2UXlO4Sh7/SuzEnkhSUBQO9KX3U
Wu3Iy8+RbJhzNbzCbjGUgXLpB+TiybsfY6POPsXcNy0kqR5iCj0qdRp3sjz6NjuT
dUg1kphj9tviC2zW+Lhkja8AvNg1b0zd2T0B+tZ5AjfIGYE1ZIu0hNdXZzvMZQtj
aHT2pMeA3CkmUg0p0q+IChC1b9XRUnzkNpU0KoElFGrci3KVEAlFWg4WDWP4iv0L
8zxgZsVNIseQBvCESG4WtWNV724CjiypLRufCcZi0jNsz0m24krMz6sX+eBWEQNS
4/20blsnqbsJpeqN0QRDXpTe632WY8XkWg+1QCQPb3NvowCEGDj2PXYCqISHD3Tx
KBmR+WSaUHarJWVaTHz3JHdzjg5ifb69k8o4XTpbIj6y1xb8qlUBuQk3Yqq1vx6k
5xqjctOUdTKX3S7mwkp4ZHmYkpId780YMMiOLxUhUACFuiGeJWdbvMyPTDz9ryba
3gij7S9UODW7BJ5Gml5eTfoHncfF+4FIHK1qYm1F/NaanIevKuYo96w3IEwmlI4C
ZBGvMd7aJYrKJ2N7SDuKWs+cgm1UTf6fLn2+MgJVUE4uckpVza9GLBJcyFWHh2Cx
CUcpoMhB9ypivqoyFNVsGqJVpTCooAxkIJFMW1+77zE29ggA2a4wcEO5M1s7LpNE
lM9ekeEGCMnStVKW7k9YylGlLv2AIZFiaKi+ITTPfMB68lMmCXjfhf3ZM1B14UTF
05YmoxOSKcVHe0ttJB4lsvywnVUHnpN4EaNOkS3KWf/MJy23Nuc1kV03S6C/y/ze
WlNvqky9q+1vZCutqSFk2CORaeiBYPEhv3gSJHeOFD8E7Ij9MxUKk8S+DiuXWD/h
JB7JCjU8DkQR3GA3dRKUICf74zkWcpfhiSHRqZglpeBFnu2OOIVqHBa3EX5PlWZj
Sxr4elvhj/ANChFCEYEn+b1QZZz1XR/JrMjZXdpa2+ptMIXiowaPAvgGpdOP03Vt
Fx/OmY8gIwH9SWN4xQD7upPaJiVPTzA6fcnJ1JI4i53Pkp0GdPI9bNBXgTci6tuX
/+Dh1fT6TNEPGlpXFBPRcgbfgeppAUHG63owdgNDhElkDOWiQTGqnEdP5Cmp0Hmz
4zfywjFysMIDAA9Vo5guwLv1QvUimRuYjLm915FRZrJnQOakic9/fFY2ifEweoxq
0YCz4qK5FusHEoqoSDrT/LRzVbSrLBy9V1hRU7L+nSF1BEUFE5yZpT/yopgkQT+p
NWd+auc5FGyMt9K7TfJXYH+rEsU3QLbHF5b0pEcewvMlbnHZqDV/gOWtAIvBAO6y
nAVCYuQHbZ1Bh6VXZ7HlnuYtnwpr9ChgjOyuDfemsznUSfW91SFCd43h5QaOT+8/
voDOA5RRVz4aq9oZK6eRevDyJKfO4Itj9EzH9c05OOIhZ82Ws06sL8ypG61yJpVw
bCn5xBjYxmFStRL/Q5fpnzQEhhmh+v97FiCqlzNaEjkK8GZnlpZrhUn6XhjP0mDs
kCGJsEgGKEsnmrUGl8EpP7Gagl7ebkG/PQziy2M935/Y5jGOOFR2XunveeSyLC49
VOHZCpdwwNSuuOW6AxXJwV1wL57Ho+QDy+3E759axkWv6au/xlIOKvCunuax2cJY
/0LWZEvM2CpWQYH1/gYN9wclKVz7eBmUVg48OgSevE7DAx/6WWSyJRq27QYN19wZ
AZC0opIdsFV9AIxBG6uPGMLYT0hniarZmhzBaO5CiGhmtIwg4JloPWpzwBqluwRt
ICGP4Zs2HY30fO6LvmC9MN+TJdekrYHLyYrUlZzAe3Ej6HtEJwlHw2N720SIvvaI
47mDcmfBV2rIAMbpd3dM90vdM0V42pyqeG5bSUXeRgPOWHEWnNYciDBnK4jYqDQs
ImSbYQIUXhztGwKHoMeciSVYmIzbuFZk47nusIKvMD7uw2U+E9k2f9yL/ls4kriC
+IQXSylZ8Hdlo8Vaxo6Nvp+bq7/SGVfiOzxh0aBk/6Nx9Ge7aYxTIqb8RJtq8LgD
ffU4ZVMzn9iOW1TY7nV9x441ufyXr331r9mRn4GTlDCYf8GJ8kQDarx8cQlrUItQ
f7Nw0+zvudOnbhQRVYsZrfH8ZKx4toA/MsN//iHSZ97NUbgFuXbb/KR3JxkKeTN3
2+uZcgbw1b9IQqUuWriUNxIyzYye8TzSfV+qOpdJ9LqJPnZ9X9XnUjQQEOpr+u3b
UuXkivKQpJ9743z+AWpsuCTRg6E632awz9ZsFQjp5Ed1gfV+jGoAmlqvOntd7nif
Krnqqz8EqFTwE5a5FeKtcyBcBA1TQ0owh4Jx/3JQaNPMYmCnt4pZznjFWZ9QIn+f
8XOJdYHkSeb2FvDBGyFx+HkNXAvGvnEDwDsAmQ5RIvItubtANS0vIbO/ZCRcXE7r
dNrTwKhkyAqfstTzKqlDND182PFcgHKWDMj8SHBMf7R1HNtmBtlCCn1BJNaNCAQ1
V16afovcyHE6qveWYmOAwBY03f4lZDxzWWoQ1trpjtsXwZtTSus/cF7g5syjIy4V
KCDr8VqahFK0kYrtLeB4ebAHA2XLK1DO5wEYcoouzf1j7QANqnz4T7ExtnkWcbOl
BOhTEq8j5XWq4N2rOq/uEQCaYd8fxE6b2ZTTeFh2FxUupA2FdsisdjhlaUORUM34
0vEyZoswJdGBHg9oCZm0tLsvP6+k5aLfSQqe/5AXC9F4iux1EggpVEF//vn9StTp
Sbumhzn2zBzRR+i8/giDJ4bhSdyJs7YPOLV21LK6geTlkqYSz6GGf+A8YOxzvOiL
udnzW+uek7sd19x4bdUfhSYnqPuJrEzd4R0b0Sun2B07gbrvWOhrcWsgrrcfjb0X
jfeI38vVHIdS11xt4Ef9REwfSGBYVN1HG+ydYXBUHR2TSzsWeqo8nkB4YL1+BP5f
NP3680Ko5VVl+VNgp0ZCJbvalFXGJb0NbSt9kC5Aar3JMzc0FrcJ9PbHJlAYhYQV
PCbZ8NIjYB0Bh8X+fsOwkNhjpaLBYD93kccarh7He9RMgApFovB/EjEU9q8v8LrV
8NxYSa2XiL3Gn8ood26fimOgtFXGYsRPEcj5MfRYxQc8MbE9FONjj+AvI+HeoiEX
Fu/H/OWKW7/KIxQyooHXs9AdCvKIsZqpp2qkHBB7yCf2KxYjw6U5tGWYbqzux0oV
Mxw95U0khM11yotJ808wdRYrRs5GvnmtIjE14LJUMJS8RC15FoGyKE7PNGvWhynu
xi4hYQ6jA/1D9MRg+WtHoKn0/wWTOj05SyDDdSs4Is7s5Vl/bL+2KYHmahNJaq7o
fv8Z4a98sAsjb7F0ut2QQJ88RbdRI3XVNitKAkAcL64mgJFyDIRncfXbtQUgA+FL
f2n5iAz7H8RmaUInLI/zNVvri9+exPO1wOtsATJlZGwG4mvLfWQPPrmeGB6nfUJn
zROHB9r630JQlR+W6XOlk8RbMsoeElE/QPROSTNtltrxGqVAb3B0N88cuO2uEF64
Z5GK4nBgE9l+hOLuL+0qFe5gwzuIuzkCKe89CTGnTooq/GihRIHdKRz6h3bM+gI2
k8I0sp5YHDHVeKJ/j5p77P0ue/exxNFCpaXyLP+w0/sMS91YZsLs9qZFk7Q1Iugs
+OadXUIw/GpQToEDKHuqzlFO4yGxB2yRETkjPvV5RQmpTM56QKh0L5UZJZYlue30
snrz4IMEss80qx2F/HOhzoBh46N5FgmOPTl288eNHHhdqBYdmxvDPOJhQthf9pyv
sEhkv2mc4PCeJ12gGYDEPKvaxXPFXdvLLZZm0z6uaulwiPkbr2k4cnE1x72HXz0m
sg4KK2gxkEKscSXXDzTJBw7qCiSR6Ueo5khM3kWip1AhJIyRGWVSyCUYM5ygDDlY
c5MEeHb8KqLcF0mQOJ6UwbjSKtkkADmtn6vnbstLSri7FNhKSDpJhV/a8JsLEWTJ
6pmbJhKIMtcpGX6otfsUB52yFQjfkAzr5ky5640WRoW4ubS1I3Fl6jz0AwgZViG0
hTeis+/tvBMwMR2l2a6Ku9tQCsHRfXXo2suUcNQdGfgczLzU7bJRJlhcY4VRTJCp
LngxSbcqqjkyTVPUixDILjZqnVUcip3ovit8MK4YqRKi17Ur6CMooSmOcN5xwIRx
cJQxECakojA1s8+p0woJxlWSKFPvweycsABQtUeLCeVHuR49343bQ9T0VHkXqx6l
OiBozlJXpz5ihSBcabEI8jeI1VzJczHWtIIjVHYVLWT+CXLDKLP6tSnG3owUDN1B
pJXVNIB+Qt/KIgYg2eQNpXvAyWS7UsndzS8GvhYVvCKjWtdfT+kDVAlGk75mwanD
fRAAdd1um6RaBFXHhPsfkWpMfikHGgc7x5jFHsl7X7tj0lOYKeUISaLI+R3ssV3r
Bn9WgEZFvs5cMpuVnsCiFrksgvlrA6iWAnTQ6WIw8c/k59bcaQovBWqq5sXac7J7
tNaCuaGUGZyPIeFNMaJ71QLDkg5eSg/YClrDs/hp/LJprIjd1K4DgAtH5sseu7qe
TrBBcKZamS4MuArWRrib5A12j/HeWMU0KgnGqg+nkKUmmNE/0mTicPRZf6fBSgCm
BbpzSafogE6NuTHUgkGuY3EhjFFFj/QGL8kLPgSAUYe0uqNMrCkDoCX1JtomZMzr
xMAnGR5vIoIkcr06jqN8iP7BFB6Sbf2GUMPn1WEyvNVMw5ud5eh1NdKsXemzoCg7
svV2CvqYqUvgxDFGlKBxfr65v8qvtZQ7VE2+wG8CKPSbSAB4ryLcPgwblOmkB98O
7ksAE7ZSwVSyG/oNyC/6BTYudLL4bgIQUDriaDjzG/AUh53IeiY4d444LwBFk0VF
iBykZHW0ndxn11U+6fLtzXDS9d2Md8r4Ktn1mh8DYt467mR0uImgNaZNOuS/BP+d
xeYNdeHfQ58HguJzWR3cMTa9ZLRg90fzTic2d02oTNeHuZapyTTeOLLh2zvoLNdc
t6njMJC9+8Zi/CT10GVBNwiXr+u+A+CUv/6OMOoWrKiD9T69+a0x4/chEsMxsGir
vgT5e/1LNZ6djEDk42J4p/XqRSZgXVOcxEst7k+QD5CaASlWEgn2Kof0BUx5rRQQ
K+GTI/uSg35TlkMGHxgvPNMCAYVrzFOQONIOswi+5w9H3j0oHHk/m01i/a1cPJul
FTyoRSCB29IKQ5eZfy6fK9WsfcywxW1EJNGLRn1obNYdzAoHTLYgBog1j5J90PUb
bLtE+PBBqa8r41XPy1XI4ct4bgjqrft/GYSYU6l0kHpDPT6OBKPXc7n34RSpNVMr
YxnmL6DVtYb2L77aALPJhH6qg/5MePYc4uw6K1H91A15G+U7ZDlUe++eVmEAmQdo
2KQXOp7zXaAbuImIAMl3iX4VgB2Y4+9ureBImjHTChAmMCkNWEXCxw+C2Si43aCT
BmDvFDmo1XUoF5Dzz7xB683A1T5R+4ihxM51nu8i1B9VjiOcyWPXJAxdkYCu3noE
LtanuqEnOVaulUfeGIBXy95WHqUjRVCy205lg/79VjZk8MoXtv+wAdqX7OclXW0a
gycENC5/bu3qnviTZJicndDp0+0mA+tJFPdEJHmrN1BmhniMT3lnNvHB8LmiPvbL
SSaUSZ4UDtI54I+gyBZVvBQQL+rDOgteyA3t9l053ORWiJZ2hFy9UpMp4jBRyX8U
XenHtQOJpkrohkrG+bUsfzAIHpY4v7H3S+6Wi+sIzGCn+FEgRunw39Wu47Wi/Y3X
JxHdt+3KFdhxqMnzGdpTDVMaBZe+/DNqhqP1lP/31KeaTrFu7kxbFWDR2b2QbIlu
A43TweMb4OA7MCldH3BPaVcZ+QqRfIxi7H0fao+n3l893SJDy6s+WMLvkKk/9q5S
CdcRJ5PS6HIZgPBvp9eyepCavjqBkfHFKM7h4wetSafdAK2R189Tw6Hoe8BUdsXm
VJAtKjHoXSGfJvOZYnj1QepA+M1XP2iZMorCuK7mBXEse6n3HKnPNp2MKTOigt7R
m+8edazF99EDYNSpaJUwXsHw+X/bBAIMdxV8ElmcddQedlztnOU4IJ6+0EFVeayH
wC01dZ7Nk+uQDiHgrznSyRnqa3AZ7Q/5PS1qQQAU9l1rE9gfElRm/105YXDqH8CX
t7n0d8KLjjMc/XWh4P/TSs4f78zWA/+2FTc9TBPo3UgWSLAipYi119z/gbu+kO6X
zfiYvIONMTZ7ORSs6RJMIRxvNsAmTrtYNCSRBLlgsF5bedn06gyrDzvqT9KV/Ib/
YGu+AXTtv2lhYiWaubyE34eRrjuGIInetPQ0qN/yTSU977LuuiSB6ckSzm1MK2Ib
D4pTjHydrYBlBxrYQVFDhQyHRhllUhQg5FXH8U1fkiKg80QR7RPm8XLzFW78PlWt
OoWaRITEPDYsCdYXXjpGeo5Wbk/frb2fN5ny4H4U8X+x1mESjvgdXDRG1nAvrada
usmqfusVbfLnk5Mkm/5FDcDh2+ITU33Q678HSA6aQHjhuZZCf3JE9ydre1Cxijda
jEmOWF3TWJxy43sWUllI1KoohpLnrMCHAS0mN4vtCKJC5uUjhCm+gFlpIEhCee5a
1Fc66CitZqrPYUVOfgAgxs0Z7RC7BNEM1GNAKSDIMY8fgRd4F81aO5tMiFnR3BHf
4NTtgSKp135Y2YlEoS3nIhKClARJSnd/qXCdJga/TMHIYNhodaUjIfb+3GUeoyx8
3PyjTl21/wfmw3b9mxAFwuy2JtijjZf2gNNvlChDkzBsSklvD1dREyGFPKFMgLOY
yWKRdIBbpI5P6didqu70/ZkH0RBq+ulUgZ1et47pKrdyLhlp8gPc2dhvuibos+li
uZUPuI+rYdc6LbNy+TTMCjxby22wQy8uJdosA8JVtTXhXbXVdsGHM1r9Eszpsb+t
sKdQWDMZACloh63uf/Rn5TACATlzwm6q3mABO2hKJmN4wLRax8cwUi3iIJik+NMD
y4yjBRSliMTlIir//PzX+lougHPZJnv/F8PyRjIc95TlfcMlfDOXFHyT2qvHWufL
E1vV41G453sBsKu7rcp7iTTje3EFxSLQAKpqAJpAU5IF6lZEDSeXSclGDjEEwEkQ
/eQ4D9EKrCYJxl81LDWrE9o44jps+c35D6KkjbNmyPJK9zRFkJb5ReXsrxjyTxoU
fK/P/ccl0+tseF7H2W6Xo8avJpmmbNSXllIhpOagP/x5qnJPpS/BwkdUf5yIQ5ov
VXbD3W4n4Mbjg9NpcQuBQVXEEGHlChDa7+A/gwCXH6TjiX873zwCdkf2hBEHaIPH
VyOMyNCpK5dRMiaETWZbu4DqdlTg1eXcgX2hpH2k34MSm7vfuIio9nYYdZNawXck
8o+HjRqB53pdN/Ey3cwd3YAAFKxbvexXavOGksPaLp2+Mz6Bd3mrNhr5ggUXIT0B
iEcAS/C4PQM1tIhwpFsNeyzTq0jOw2Ov2yn+hjBRfAx24nNLiEVvbzsfR+Rmj5S6
221Ox+kpV8W8VvKYeYjHK7FW4vYUVsEO5Ghjy/wCfZphXklKqeLCeOH1o79xGEcP
s/T4wtGOZmoq3ZoJUAhMywJomg4siuLoYTUenWfe8BCqbLCSxUjMnXqwWUx9UBlE
m7LQa9Nn+ilbdBc6nt6ZmyHGAWknFLaoz9F4PK3QFg+jXFdsBf1f+cyxRZJZIaCT
aN3baiyt36437KrNPbHsqT73mB3y9Rpq/MS8nBl8DADLIvLiLylhpBREhLb8+Iz4
XgtEdyrQmyMfNS4Vni2f6T6Oxx+w7SqDi/AdBVhy8zIa1DXiVvgJEQKogX093pqB
7Ay13umd2rUbJ3+6QrnF9FCrOX4P4AbOoriK2stK1xfg2JpPA8y9ut+JYMhaJqgH
MaxbyvJMv3Dp9olioiqd+0sepJfauLQP779eSTL6R3h1jjStDLccYs9XSRL4hZdb
lr8+0E6Y5mb0nE59QX3KctRXIEB/4Hs9FotYPO4GduNxz8+Ns018Mxx0Z2BmER+J
7TWXNCkawdnvtXF50Of7sdiELlb9o5vQpoO4qdLeR+70T3wBTfXhS0NC2wOhKfVy
F3FTRMj5d5NYV/mi2Nef4RLeH8XWXSTOv3rozMUtvmnaza8ePJDAT6URyq/3wdXB
5No5F6/1GMBaVHS7lNHc1OY0IDnI/8zG7j4Kh2Kf4SSlwDB8TKSBdirbbsEqCDGI
TB8yJb/gEEwDisF6QIYdXLxe3MB6siOPmBiBS8KUbUmj7BMVwjaqSGB9St1GcWAq
84iCPfJ19GZf+kgjPyOrA4Dpk+p5KpWZyhnwmXyOn0Ji7BfjmDKvxmxwpYOqudz4
zquiznw4ub8Xqw/DlrJNH7Nq6ed8eJxrywzm6Evnko+1hjTM8Iv/r3jmo+s/rQlW
5wMABg+9u4Y1iodphJyvUmXYFXCw9L9BgikRg1gVW/2PdH6+KMcktIa+6efWqpob
BXLKlNsa0mxNsa1T+tb2zAcSjsaETZSFHlRAqcnQ7wPTia13zuHR6OeamGKFP6yr
HAnM+PQDUurGLilQdJxKvpAQZlzEoBNy7zpDesQsFm9L5lF1UNyOIIT1dw+WWSGH
e5YpPDr00e8n5r2Qcm0FFbrqk7A9TodjHjaWTWj417y7F6ZpIKtmWvjGcckmkxbX
qwENvRvEQNbeRH7QJLC34LXfTFwmXYjfRR2hsm+RWI1VDeRzfeV/1YBhf2niJ90J
5y1Zo4kwpNuW08Pm6B6pT6epOSDQWg6kuUoiTn2B1td3a3L3GPH+g6JjH4TXyVqv
oiMDWHf8k7WBDtBlsUGvbFDvl+9kPxs7aAfgSyLwNUmXRQgyfph4Rmxy1iptbINk
7NWc4PCVSY9B/8W0XAqZyJZgDhKlY1X98iJJgDG1o7pTRDkSc2/R7bMLJL7n15FM
qOekwSttj2cpLLkVrG3q1JJoogbRrT1I5J0AsV5oWn4Eb3Gr4i41J7ViXuzDz0Ut
1pO0L5eMe55PD+stExt7AmuxeTYzCZvqyoodCoMUUrc5WAIpewaLeS5NI6jlRpat
tRY05psp4x4Y6h9nFLJB1ct2ndLjsm+gL0dIzKTz3f9sdT/JqFR6BS0qBWbyn2mJ
KfO29Mj7gyXru1ITuR9ygGTN0L3vqqhm8Alqi+buwn4BWcpxiQXpkzucD6ONYmQX
mk1URGxgQPRjFpfW3YOYNm0whEUQXWafhq6DmxfZmBF2h8puuyYsS1B85ldzwJRK
fSAKPHwd+JMOsFAnw2MLr2JTjKnDTWighjjBLLGPmxfGrOnPw7+n3nIR2Y2E9RtZ
v5JuGnNVQNTJlLqh4XHuuM3H2beRDaVZkicngkt9meppqwYSlIjp6jNy8bck2eel
J51KLQonW9bP3S1P9cHeQTmLtSC20qZ7xqvkM2CXudWm4qO+nuSDJKtp71JTJGr5
5TP+eJd9jRv1HEk7Mje+tqy62sw7JignnfNf/tObyRM+OuwGaHaLpXbIdAoyUy7K
ahiYuHGqxfNZrlyOyZ0QT5xjB9nfGxUViN3IxlQkgGU6oJibOj4aO2ev1tSqseTI
WJ5n2DyQOsvG0syJfSf8SGtYGWhlA2LR7wYe0mAxPsgVcu+oCPBrk5ePzhpH+P97
Fyi4088a4B1YHKGQvI9RtrG8egZ3Yb8EX4nyfBrs5//ixo0Td0BEqrs+f6xDMToF
aeWwPXKYjOcpb4Nohjw3Sd6dOK4i3F/9LlA1VwNIg/vCJyV453o0llF0+QwI307i
0/rs9VVxlZbe2VmUJE5N5cxKRUvmhj1diBhY/WBSuteM1rgXW3DJ+gSbczSaM0vc
BVFCwekpjytAjVJwFzEOqVEFE22qjN3lhvCUWWGsXRhukGqc/waUJBioceXCgJON
cVYRscrxk0tCmvR0OM1Ut2VJthSvgZwMhDHOupBv0KwbicOw4ku3whJ88V21SNGt
POzg2/yLjJiiXyjWeMG8irEkGQRcSBYchbFpFFdxk2V2SeOfigSBm15AmiDAlIdH
LMEg/QZwP4YIGu1omcEEjEDnk0jSBKHCat7rOzwl19wTUWCIUi/cUekqdXVjYfti
kLekJZiEpxZpKYbd1h6ANZF3883Z2SKO6EsPIRQPkeMD8kCGcMDc7ySBQFECaqLf
iH+Oj4HwW53OhEIk4rAWMS1NM5bZ3fRTlaMKdOwKR1qjA6MjB5QTKf2LmdoJCl7t
xz8qIesrKk6y69RkCtM7vfWTlQAWMF6KOwYBjIRiVHGltpC4VUgxY/FTIiEKBYn9
7j2evXOWGojPAY4pF8/c61pKpVhuQ7OZkrTsZWXf72kMDmaIUXTE0rQ6P6Ml3+wJ
PWQT9JsSQFKLTZoSa9xCYQuAZyQ3C+eZnpXfzS6w6BR6H1thqgvGDkL77Hqyn5vC
96YhMAA7Hc37bw5usJBAR9QnuGM3ftMkmFloDUNqf7ter10p53wwdk1SUr7WHJkY
FfHpc4iXOk4hmNStosRhpQxak/AIlNQcljSmJGxL8USvYL4vhw/5rHUzf4wiFZwR
UgQFxrey34TPygy25lRJWEFjLDvzRTp2NswQU8eUKj4ynxpYrcXu5opPnl4GiHvu
U2tcFjGSfNglEdIs3+kuKVTD0p9YO7KniavLRNLbaXXqCWc1pq6WkSex1pgNbLj/
lDu2k9/T61wM2k7aXwjeLwPRiee+Qv/0eJJT1itfO675PdpLvDf5oZkdirHnesQz
bdqEJkoG5AkqM/SVxnIi9lxAIfr/9tFcA9WXK/HSm4pKjcOjsmYc2zSy20P6IruJ
CwpCeS7XkkBPBtp+bSjOHeVg4n401TAa4DXNTD7nph7VSw4TTCHX9PDLtmLgEi2T
9TunJsk9BqykmLsHY5K+DhUaChxd9yGJBaA0gsjBWoSfOBNzeWGjiqylasGv4l25
ntFGy2yuxaHeptY2brRUB/FwCfJmOv12nWdMP3IUnX7g6S5rwnDk4L7C1zQteVo/
8fEAu86M/g94A0NbjdVgs1/06m4KtH1fNYrONknkulNqtKzlJ1o/aeBv4s/uunB2
Rk0h++9ntU1krKdB4kg0aNvfa45yFYPmrSMErkyjR911cCWePV4QsjJQS3onMYg1
vSB5qTu/K9HjB3mHn//n/eAQuxnsidOGR6MEx2SHY0BFy7ipsjmu2jZd//Gpf7CL
hDmbRhBURZMUORNaswPeiAl9kt9qpb1dPcK86HEPQIOdid2GgaBkwP2vOjIMBp1i
Dnw13HM4lipW6wYV0XiRzdzeK39G6Cc/Ugc1P0kDyh+RC2pEDVKZvGrJaUG/CnGf
wC5iKdtgdG4TIjEZr5feb0Ny/wAhe20XKzCWlMOFDrG2aQ1P5qbZ/6kyvn/O4o+F
GpJz3zsOE5Xy0NV4x9CVSCYnb9tDLq4/y7IU8nLJZCaB2OTVbrCZot/MFaPGeVHe
C0BhR3KKG01M9pJtVVQYsbtcaBwkIeDfrKjBtKdqayiqOgy18MZgaAVOxIRw9h7e
IT93MLRujpx1SLTQJ4Vf2BOu7TS4AwdTQmErm52x32IURDVL2L0e1pvBtsylnquA
SQYu7RarcyFFZF9O+57va4p2DaowEW82Q1a7d+lyAyfahOk2P5b341l4PZpLhCXT
hDCFQx/BdxDuAJu91uG83FxTyMlaUeZrT5DPza1pYguBJBnahJmcJqumKEkx/52q
JpomNTbDB+ULHn5F6kIJc3aflKIa/25WD7GFrpbBA9ue+OLfuor5YE92JG61O24B
O8HLzrUhrE9H7JAyHR8ArxX4bWq3KuYc87Nau1JMbBhWl97CW7uVTF5qUedydlCa
OVF0U3IR+C1iHiYYA0jHx767ltllcDH8cOnNV4k5BzaOqjnRQdK1XRIu3vrImeEr
RsRSrQGKyrtWOIum5T8XowQe+UZCN1iaGUWwBS5FXscJEYUfwFomSR/SUsaWvRuX
YYpMpOZkJJedX8CpvHDx4TV915cS/RJl0DkYz3B/PZILiudLEtAenvm4eiitebns
W90DX49qbjNAASdpFuK+Re65Wsi5RShO9jnvy/gOpuTQIeS6tj257DjZSh1rkes8
CZywK4LnJ3UdNTFZgpWkozvF0gp2xg1jy42TdfWe9BVVNwxeCoIAo3TawkrZ3g7b
+DzbSRML9RcGtBBX3FcyJiANQxLiUC8FtnqGjukx2xbgy0vwiVGIEpqm/OHEe2+Q
fUJo5y7g4HzffgOhXhHuP6C3+ZpDr6RHLltjWGFRYApTYpXsGbHuoQXZZ9gJ4yGb
jExDS9BMH8XeeZ6ehDXGGT/YVe69dz9s/i8rQrL9vwFpUYw9fFtt6CUkZkm6Jr3S
HW7UyKftEz03M5GOBjnkRvA71dmvYAXP4xEnOe/lCaikoh3nnE5fiGoxSXDVvM94
wNkzl0nVmn39ei3oB8lTSykIn+iK5xq4YpBInd18xZsvoHYj2wuELmOJPmHxRLde
p/wYLLvlHIksTnWvdSFzX5tvVApv3o+Vzfy2+FP3FQzCLSCqQGLwnm4zv9LlFIm2
QaYByZXqcKFv3YdG3j+lXjKPaFNQDej7jxBbipmb1U7wce/+G/5ZkDHJ7xGdPb58
HlFuw+u+7QdeEAcTwn4ovR2REdFvneKENpeUol4I26xdiqnGWPkp7oTilTBxrbMc
gcLS3HXVUbniZQBCUzcoPBKr6oWDVhGDZcm+GmH8+wwzQuurY67tYy7ivNdeaDpu
pi4UTcXEbFD6fwyOwjpaL295gu62lj1c6fEqnXwHLLH10ER4/2xixCDZ7d3pzYAc
JysiQeJxGPxEbyAM/dY3pKIJk+Zzf2h7P1NXgOPj10A3W/H7jDxst1QJHG7//yQ7
D3/G8ETfzuQf5nCGGyrQ1DWcviKHJKL/sypJo+dMRXjthc4Tff3MCYc30hXr1Ozq
WP0NmPVRFLZuoFNjSEZnD706kwNDijTQoAM+FjB/L4ryJQFNoRtHAptuGh2OYn7W
5h9EbbBj6jX/gB7TbxuybnE3Eve6RNq5beyV/316ky1dWwGtxPgHwQsEI5KvT+vt
OIKAaj7cKyneT8+/Z/tx2Oda2s1F8c+1Py0g0hQMMk5G2surmNMq78eknBl0ry0p
vxqzOVj7lxc18YcqxYYCS3jFoLJFHgMBSNP9UU41mPl7SqHpN9115YC4kTCQ3V+o
tnEMYn8uKp4+rUCIO1sUJJTpJsdzb0/M5TWxibAJNxiEcpeh3cs0UWkjP4s4lFed
UiZYIYabkeiRTq5OORDS7MqV1+ADEybQ1t98okYeiCJI5O1JwPc0S4HzaPrKfNeW
/jeFe2ekCJuD3nTmWmp6bwGaBwTLo+26msItl2F72VQMBfjv48MOg/UEWI1hJzyI
WjgBYU3IcjN8VAL8Ny1MVgvzBvqRclAew2ko/bqExT3oFPig2cpuhKrp7IP9IFvt
HVbq4cuCx+4W8wq1R9nvcM+LDx34YWO2AuFAEx/4Iz9sfts3UcpqTJzCJwJCgp68
gw49K/szVD/GAsiJudGCXN9YXBydXfIhU0fed0mqCsVD1oMTLclwum3RPYds5b4V
bEBs1dBvvjkxBaS+PBa+IThrh0Sc/zZkpeuoXBN6KYUlIjuwrrRci0lAvqWPRnV3
XVgDEssJlj0ujtcWOv4YHbmT+lq/NE0ObESWmAULfncp4m/uy7yl/s1ygxMsStKO
2YNR9pihT7XGCYHPttA7MOfeHz6yJCdkqDK85aX/lWP9uYUZzrRt+sq3dpznWOR7
rcTbUAchZKObTWiR3u5T9gyDbLXOz0Ys2fWOaJScm64Y1cHQVH4x54ZalSTHJaiC
PHiDuosUqvCAZrTGjKR77jDkXU6QeP7yBQrcXXlNnPhtIczwN60JoEac0y264YDh
2YbV9ebk/9oPM5G66PzAu1XfLjcBPrRxd3jVXcAAAIUCR2zY9Yjqe0Wu2YmeelWT
/jcV9yH8wdqDbUi5evkAI+v46ijUScXqgk7BEvY7nUDWFOEn4E8mV7CbtXIkpMvf
QKp+1knFrxylKHhb8/tIHfguIM7eDl0I3Ujr8/rm5w1tF+n9WFzAawjX/ilZ8qF8
s7GwJpewNfkf2RbFjVlPV+Wb5S8RsHQ2xK6Fqvg0sLKTMuRqrNJIbMNqlDtaW1wU
lxOOvE6Uqjcx355O2Cij3JKsKTlVW9B6kN4g3luUwX14L5vMfyfKEe7eWX9uqFqb
loMgrRhw446OLvHwkjMnXbrIRvEbwvyTK5u6ie95peoYbKKWfz3NsWhU82s9C0g9
NAhXBSqjO1hovdySkAAs0umAsHN+gSmCYA7E1iuCpn7PuxyzI82oFSVBu6oRgccj
kjwc1IS0frBK69vlCGol03MDHmx5w4sXnq3fSJ4H5Dc01HpltNFra1fhBvw6p1A7
2CPZ2/l6Od1bCOTPu9c1UM0+t5cKqYSpmU+HDM198V5OqaTKKuQq+2z3slMhCoPC
ZRXgmdZ58gy9uUhzOyRLh4HgbpliVu0yygBfVcW8unSSq82vrVMNn11xvYuJfQIJ
q6NE46Qrxp0p2Vxcvia/e1qRtyRpHhsMZtHCyo7HMLz90uG5WBUnOVIoW6kbzN+a
WAoCH0ONpM4p8fMdEut8DTvGknp0Cqmi8gteFoQs4dEZBs/JU00doJskMhsxvS4y
2poi9AvkBUF19cl5uT9/Cz7VpPtq0DFtMF/BLoMMQtBEsHmjuirjlTm4jDGopd8S
/sb93HZf7NrIMZf2F21CQ8zAT9Y75kMGtlNjzEn9zNNs7eiRkoRKoFdmK+ToGEfZ
WDUSfxwIWVW7zzFmA0y9hCC4Qt705TVDYf/saBvIg/TlGOzu2V0IRf1SAdH9KJW8
ymaRJfIL/pzVOqhQe2jiYPsP/BH17TieL8rh+/hgRZWPpqQfAvq03DbyAMKktKsv
/aFfyQnuSELCEVG8v1yIlxM52eEu1Cgt6hEbYRHKFjkSOKt5RM3DekHm4H6HDSmy
AxbuUQ80TZWCyauhjh2E9000VYIydGvjLHjEAk9rGWpn6SZivQEqc2IuL+2IpfqN
HJUg4TZEnNtvlxekul5wrQBPgd7bNd9mGw782ohE7roJZRHS+0fscgP/vqWGS9Mk
SxKAwfJuPsdSZrtxYwJOB26gsKGZMUMITiGDGkwNa1Q4OcMG4DwiaAz3i0YFjKRH
DWvmlggpzFj2m26VFWykK4pplSu3YFm2sSIXTxLtz67TsbjiNgvtqTL3z6Xoyb/9
4Ac2BmWWOaa4aAnl1kTTl3ZTScvt3mNLG+nO7YX08/LIN/vPDu8a5NmwouUnKyqn
fNfYrWrIY6GN9MHJ58e2f5T+dZi5P/KYvW66omdP2CfnqhHNHoAQk9BK/PH156ev
yf9otmY7bbkNntAKFLA8YHxj5P14W7HSNtj7lwSZNEpHigDBYeW5CFvoDV1cSFaB
L+c7ZfpEhq89tCjpBsI4X0qn/4eVZ0MR8SEYIeqmUexScYyAvntp/77cSoKGqXYA
KAQgu1W0LyOo8nB5CJsegH0fsD6VBu6qxCfRrw/6FYPVOSYVjpqDhNiOLQ4OhvBy
e/d2xdxdygUuC5dsFsCfXIv0FeLexzQWcpkQdIoc6rDMeUgccDwD2WikhnOpFdaN
PLUklGiB2GS3fWYb+GHkEUCYrKvKSxImjhN0ZoLkfU2FQV/A0CZF3oMSDN0VAU7r
98cO0ytJyrWFzT/0CEjp0v1Zb3FDCgQe4FxK/Mq17sJ6i1uKYxdEMLXsgTEh5h4c
Obdf27wRiohHr8Udauh9ykg9D7/witZk/98nCH4tRDs1qoKH0f7hHELqvJMYZ/MD
9Q7ZYXJBOnVrK9k8bAuYTfqwgQbUuSJEprG5vnKdQXn0ydVsBN6fj/kJdNZtce3+
Ytl064xiS6rhZeTlGkcmTkM//Px5VihX48kO6xp5WTe6juRbhB4tWp5ql0CSBTp3
K8CKtjpQZzVxJRTeYOXYKDzUFc6toV17OhDLyLlTal+DqF6jELBdcGo8UWU3AXaM
y5Yx1IVo6bWy9/nEUx9HeLE2WNs2c2sP9PYULPBzU/BTY9E1SG04pdL86aUv6EL1
vsgOKmd0Rv622F+6voK8IE1H/farhWBcs+meBpl/AHiD7glrnlaXgfPlvSAFRPcj
WBmTrlLmgB7m0EOEv7hLwwWN+BZ/LbcyUqQRZV5SZBcP0pfBrg1S6xKDjbjec9JR
DB8AT3bYPtKb6G5IXGOhFW5xUfXRN1MpIlloFIov5DrXndYt+bqH2uoICgH1V87o
8QQN+O+oEkrUQlxwrHA5LnDhYNyIjsOWAXTBL6eEodx1/oMrMcxeRb/GhzlOaAqu
LnbAadZ4iUVhM8g4tFX2Tus8mbIu3Fzcpfkq4eo8v4mhc4GwSN6g7AzmDla8sIbp
Jk3BtXEzsdmvQSe66JBD/1YPMyFzdW48l6MqauTrjDeUKO8y/oXFt56iZ+l6no35
3beeoZPl9RI57soK/SjFB0yG72BOw7JK5W/xGH5FIp8AZFXnZqIMdwBRdjcFWw4z
inmxPprTx1LIvW0kBxfhPruvGwRiiykbVJzu7kpZJZVTA77Pq+YpkoxoaZsygaY3
HBWWlDxODF9X74idhGBX+VcofNPc/CO5BzDFFezLlLG8rvbK0Bio5vk1QdHFpjIQ
sWlfJnc/FWZeYfYETbU0OaL02MSRySz0foktpN50/GqIiTKtdaynJlwRsxAmpLq7
FBz0A7XIROiogv3huXfH3Y+w5w+uHfuqRpJKKPxI92ThT+p6TneO+RLzY1Hktirn
gbhebNPE9i+DOcx17Y+SPJ6Z1U8rDs7zedRBKr/YBM2/QYxRJEQ9hKHnk0ssH70T
9iDqHfLBcDh0mLfXPlLpj5QMbI0hByOtKSDFyJx2np+TJcIer4IkftsWvDy+ym9K
MBpXeAFl+8kzUfWnakm8eJVmcswY7hqYvI5Zs5nO2mQhPvGXyXKvp55YclOL1CzR
/FsIiUpqbAU7i7VKSCRy6RsITiWcEK3+xA8Yvx9u/2KYMe5Qhy8kNjy+VRSfs3VT
B5bSaP1qqmqK+jRg3ca91a9g1sQj/MklWKMVlMDV9XbUfHr3A9hwJ4lU5j/bL2cB
8N+9V3bSGa/3bqqSALegpHfb7XqQqL9I1Brd0MK0yCo/eU6YqF/rkYSNfQgCKU+F
lnZg1kwwYUN/IXyIQbcgcgGMdT3OSFhN9c1ArYtaLYDOYGS8cPqc0UDt/duHc2JR
b4PaIiFYdug0qOp9YISV2X9VbZMdMAB2hujS50gMDH/B+9P9NxmXheQjl+sfNrK1
SjgVCDHuxkjPAYGP2CxRzUK2E+/3tu8PnBxnjQtWeJp2wElF5NnCXm5SZ+VDYblc
BgRB9xMMAb68j2o52RkpSynEEDS/f84lRpPIxIEB80WAkKSUoP9Rh+JjbWJQtXZ+
qqKrlVNV+leZvrXkTTIWgWrw7y9p4pzDipSsQYp8HxQmGoHJigJmIHABxuxpZRhD
Z2E7GziJGC26zUz9DO2glWyN1+SI0MOzPp2hfeaww6cjCXw0FmCTxbkJTiJN6WPa
noP3Z/YU4BxD8B/31CaqlI4CGH7VUQMA03faTZw7nXtm7Nf1Xf2XTWbOOFPSW90y
8u0FAUlb2VdfvjgqjmqQQm+h21sbH6HOPYI3GSrnjbiCEE4VR5DkNDMBFA7bdmOo
b0kXFp79bPKQwvvi5WjXttJXwW41hlCqz+v3S7z8eRxi3mgvWxAvfSOn/GOzXkbM
vosWS2J7/mPLkSWJQ/eiLSC6XlpUkd48CVzekvjl15iXRcubEerJFKkdBrKGzOZe
BjjOUhMdPCo4v0O5N0RdLDgkf0goWbKsQqVkL3S4OFXRc0+Sy1YESU/OySJXL/qp
Kw1kE6K6Tg4d8jBQLwCiSKcgIigfv6A3QfzsZ6F/5cxr+we87DboaFdjSUHJ2/PW
Z/kP1Gzxnw63b8vYxFm33poYrsXh8Lu0L/Qb3Y18Fgq2L/TMf4f4i8Y4gL7EbNFY
HLhZiqAuXcJa0K4HvoIm22e6gUxFayslLzVnn3L86FsaM0tdgZw5oSTXBRh18cfZ
vpmgweuqrvgznuRymQetLg7fwbpGcsJkAP2Dyf13x3MPKhMad2OI4eN308KquWJ/
GFC06TO2EeRHL8OJTkoMMiRLkSh80L/OcqEr+jTXUxOwXoh0PfMY8trJGEA7yyyk
hHjp8ru57fS8zRts+IFxvBiDJSKw4z0Qvm21d3gdThP+mTp/I0uSROyo4gROfYQG
9WLCnOE8uD1EP6ArTDhRSRmL2IB9R/hXbM6rF1KgCs5ItCuxoeV9B3Otb3ZZBiWL
BYefMMZ9guMTANVl8iGSknAk7JJWOha7+RoeQxJRZKTRsl2uIOLPwM6PRcjmNPjP
yVaMuyB99G1knZgRt/FeESWwVu+kSQSd9yhQZJbazrlpmwl1pNlKiPP8inv+FRdn
ukV523taTIGYVhfAnwl0e//LWgkrQMhLIOvzpxCjIcoe6Ogowi5P6sUcLMPW1J5q
UyucBX1E3GbrAyHQE492ZjBslO9+a4CDIfwO1F21Qa9iJJnT09ALOwCH/CUpH4f1
VltCPGSWA7LpG+Vpv4KuT3qDIcZlQkZFP9ik0uu/1XrMa2l6OETp5geZUmBfSbOI
bXveuF0krTtC37QP3r1MGhbquQrZLUSBfRvztoav1cmtlYNvZC0p/ugzRCykgk9V
kqoMLdqs2htsyrIc0YHF7NOz4E4AmbnIa8DBgNJCmJdri/TCBnR03xqFCOSFZJJ3
nignaWQ6FISzqnX3YsunY9sP4m57lRMPX1SEmKxt+V6GqiysDrQ5yQdLtd7r4SxS
MzfOULwn0/ebcdrv6aMlEFAuwOegUC/cACxJfAX94fPjsDPMhmAgzyFXNWJbJLe4
XHW6AoWDVIve5h1Yr17SjSkUTrGCkaQAZdKrfiw8UegZxgmbJO+coiyIAqtGyFGr
AOdNbPgUKSM7iQRVthOAPfYXyQPwPS+yxrzPhxw5GCjNx9mrZ8PwnxwhpeWxLaXS
Bu3rdn62u8kh/JeG5GnGafLWsAp0p0h+vlz/2kUaKS5TuTRPF3daIThzRYb8w/F2
Vr81CQOhyS8IRaMFQ7kEz0DwzDq2bbY8phwZfHrcsWTjMhZLmjqVQYoQceJ2UaCV
cthszVpXA9iP9vs0RvP73wasxVuvcyJFye1R4+KrhnUMOiQaijYBrXpoHIzIBRRP
woUluoI+J6jd7Omffmao9fZpk6OioVx7vsKTHq4ZD2ZFnt+ISTzKUqLlHb2iOD7O
HkBJ41niXHFq2L5UV3LhMcwxx9PIT4YtWmCZzZ7OI/7ezTXOBtT/8ecg2fp8QJrD
KBakqK1EBq7Jc1TD4SATfokCNcRxUuqOgoJqp2WYD2J1Snh8/I/BoZBqjj+9U6su
7EwrrxaGFc6191/BecUHtvm9DEjayIOpOEMJ4j4BpxcS1WOyK4XFWAYHDXRFgS/K
ruV0UhMakjEsdoN8xhzZNdRSnTmWTCF7DTmHb9D9BQ3qg+pwbEiYWn2qdgZkw/9M
bB+OmNX2cpZFnePmK5OL6kSk5ss3ExeVw5zEQYTuPUMspllNR4iHK4Nl3os9OV2E
viCjrTOy3RKYUR3bdEvSQMCu3DqEsJVXmE/T/iMEm0Vblj9Xr11IpbMETgwAXTJ6
GDVSsUVveqq/ejB3Pv60YftEC5giQZtpzn3IEpN8JdGO25SOPQT8ddG9XeIL+zH/
OFVyW3e7gFPdg2+XgH4OOw2C1lEjH/SJmoOmRcrprqnBm4udrBOKmkDzMIaTyvrx
DTK4cqrONF/2KSmnlNPupZ/jK/TvWHb3euPvzoEVx5H7uneMZ/0VdIuQ4a1opDIl
vGCNa50JpNhr/jU5ykWdcr6zqowTgWCr+13qDR7yDUhTOXgyv1WsUgg/hjfE+VRE
HZ7cFDG9ck4xzacJMeIJAnhpBhWFluDmY399In9b8MmTsMz/08C6FDn1dBkF87Hp
Al8Ie8B9pd6Epku6j7jtYfAZ+cdAy/X/e7fgiH1sZj0Bcw6ZAHX/+c15RiAIWYgg
PIwktZJ015BP4xDWq7PrNRz1XaC0a+8UBFNBuBm04qKhxlEBt/fpwYopmq74Zjra
XlCcHzG2+LFN424wU+z2mYFwrCwRYZsQb4GGgBCX7xOKMZR+0f81mi9KxFiN6OOv
9oWOmf45LUZr1HGTX0nctdhwAZMVysueWxmJncSWtQ1YEtWUwIVSVLSk2L/hJXye
rc4bWmaRwzzvVZD57sPzS38GMt+r0s+yei+/POUUp7GFTZoDx+4tDghKzJ/GxD2i
3ZdfeMihtwPzzvUL0/YrMnZu4qfu3Kjf7T6hatLRG1B01m0OmdXrSgRK0S7gu0KD
icwTl86Ta199zgSprlGjxkQ75SmvUTHys2YMSeyDDt38a0EfbQk2v46N3hPHXT9S
D8l63EkK51WmEkNXAtCE2xJ40AhCvFvB8NKnQmBuYNamHLMDRz7J2F9xr0ZF/2zu
71dl6iSVbUOrS0fU1npFMGVI/kk3cYVHRHk2KgWYPI/2I4+8DaxhQM8SsHgf3t6q
yiVIiyycTz6+3QIhJPMRmmy7ajtMbKCqHHLlSI7qOfrizRS9suXraUQfZLvrOXd2
66m7AMqjznyrAAwihKg2eq2poWSa04PuoZck9jjJz9koEyW0mvBObChCs3rzH6FN
N9mNZTWVgZQaYnvyW18k7RxFQnyApweWu0fotVMW25Lro1Oa9Y+nkroldqMhyPCv
wi50VpfaH1LRMkuFpsC721DePcVo/BrUX4uk8TA4oR6atetwlLxL6Sbi9Tgl8PRi
v8niiSDEReaNMy9KyxsQ25eJUT6pQiVfOlGTHsAmKO46vYVJ0J+X0pZ9ZMeVmAUs
D5WM61XNGK/bYY1YOBmDYlWP2xO46lVrrPyLWO7n0n9GifweKNQRawP20rzcbqZK
hrecC83lTKHdZ3wd8DQvnE8YRGC5I9BEdPTL02hdofX3g8dRL7iQ8vcVhW8azPGD
2IYyJsgTsMTg5SR4KRt8MAZrRKKeJ2DkWmenZ5NnVEc6tUKLbPxXFfmZ8LhkNQ0R
9QQk+vOjoAFo17tqtvF+OdhiXFfpFfNmHOYChPPun583KSPG537P9RcmncOPcPu+
dbXfZ2DAQQxeAfiCx8h2foqEdy2fqcuoQV0yJjR6KxmB2/yuYPn+QfzoQaSi4bsI
2F/eWBIe5zjy2gor0UwKPbeRRrlgpQd3v6u5F2YA8laO2CMYwe7obVEfBlxyKquQ
brKviQltFppRdr2w0bUkiCVuin+HmSEJU9igoB46xqLqf1HP/7gG7Z/0/ZRvZzyp
dWs+dSyf1DXVpOBeLSdaVdfcsDexMHlCSW0SkNCC1Fygl5vjfZKY24ikPY8jz9iG
o6Ni6+hqJuyyPUth51DK5ZaMe3dX2wInn65+RP9Hql4xbNKbnBEkJDhCCaOIuhHA
B7tosxr+vQYn1FfumIPgIcYmmj8xXZxQJ+KOgNX1FUWm3CD3MBBuokGKtStPiEzF
DE4/QhRemly+h7WAt8dpCqF9qyIeu/rRlED2n85d3yPPVdI6TIuMot58uDMSClov
tRsptdHPnY9kg5hdjelFuatWC3xJ5SvXLzsW0HphmpnUbcu2Vj9uC1KIoEgkXXIy
eLBa58/8qFzb6KR6R1lISCzCxQGprKPMOgSyicFiusk4tfE0UhnGVmYACX0cSiUm
R1E0njq9TO0QWYPwKnBQqiBIO9ImWTIOHaP3qYBuwxL2NtYoR5fMC5F9UfMuMQ5n
hclnaNeRgsB7wridSA7E58niDJrijTnKG83uDqErLp0L1tl9/UzZQsorKfLBEkFi
hMGV47EULWLpnFs2WmJiJQ5HisLpIqEkDlPs+x7LU5MZi8XThf0AK/nVLLVBKj+j
DFBHeGUv+U8sMvJgLfI0pkNBNbR/IkxtnXy7lKi6YIeV32gaC4HuMvIso0u8Lyc5
Ds5yYgX+2kxy5/h8Yg2kIRBqbhIdbJXKWTyHI39Rxzq/W2bkheJUgSPynA2dOMof
NxPC9RF4F9N3/SN3+hH1ZLrrZoAkhUAe7CYo7QuwPtk1EeyPv6DNMq/xsCEXJZnd
Krv/fHygLQt15reu8f9brQqMtd3MhnrHoi4yvht4g7ucFWqrpZLJrHEUXzvXm82m
RHC5IYTFGsaYPtHqpNBbF/dkPUmLmCxTBM+TdakrgaN4wuwhsiWGrOdOWWlTDAmr
YW/opEQMLPbrGrW3HAwmvrDFlatv6Qzg/eG1zVA1iL4iyqksWGC5jZYOQ9cXxHSe
G25GKSP+7CyVzMD9MCo5zRVeZdnv+ara6ptZdRGyxHASCYUV8+p2JD5M6bEW484h
JVjDcYkoO/A8YmnYhNPo5n04UHEf8OsbQ74SWGvpPaSBkLQghk59U56lz6VVskWP
vymunp8BIA9OYI10ilyti/WXKx4vfVfSjCS2Lm+GZIa/L21gqUaAvYjIUEmLYgms
a2cHvw6ki2dI5dxFeXWWD5BSeii2/ocils8uv/UDiM6yneJuWD+e0LV3AWw3GJFm
0TdA57JpDYCFThOOAhkzOyuERWyJWCLAe20c+8gWfYNmkkczbaYf08/3cbh+mzgz
n1+sFC3Wmn2hob3YiSDruADUD/Hqc+ScpH+/Q6WOXgpv+YUEcNlEK1aHcmL9FKv4
cZTvN9jBXdwXlxEjR7m7iY5WRwkTWh+LUOObuOrLosnOsA/KLk9ewNX54Fx4bTUC
uU8DZKXj2XwbbHlM9b8xjuNxW/FsZymvH305ylgX5ARurOvD7fhWa89muPtZxiOb
ItSBDMpLUWt3esxoSJ9aOteIu3WV/GVz7H+ZzLYB+Bq0HWKxAI34RBNIa2/nVFa6
cNyMf2YVWa+TIHcqZdDVVM1cuEfbDYm3UPZ+lqFG/8ZriWoaQIQmEQDQER4GG0/3
1CkLpXombSSx0Xfb0KFH2je6FYIi4jHd9QQ/vJIs5pOw0h8lo6Z+w6jJxyNp2ywo
A+unqCddqFyk/GKhUwoNPnKUK+ILfERYlWLEfw7FN7TerLss+ifYT1u65w0+sp0A
BMtwweZOa1EY/NEJXbnUo8Ulznx7K25l+7bRzzNWObne0qvFle0CSYCaP8dxpkzJ
0eC35Qp6LfvbC037GN670nPvCJ3BMkQlhuiDi/xN5zcuVeoUX4sPHv3/vgekrK+F
Brj0rA6F00iSjv7b92LA5tAcvz+0DtjwNMwJ0gY9fHwbPqw5DQ/fRQqwyf5aGlE+
nGoTqOAD/1/J1Shz2JdRqCjo4qP9wff5TYAVNwY8ficK3fOFECNBVFy1PCcEmitw
wY3E1zL8Bnu5/sKbIAJskkZqzJaYYYFJmCcHLnWE/fd5eeIixUyWxh/pNsU8zeMp
5okV2baq5EFpBmvsdb7uHQp3SyuNmxSGclQdLPWeleN4fpzbMr+Ux2ARciOwixTF
IlVM6mPs4iDR6AVpkUQXSl2AbswN2Kjd5r9xUr9Hj/DMZLXDtrJmoA43qPhqB5H/
kUUjC4Tvf5xVJDTjwMJzhTOPIhRVa3PLcrIICz9xtyxUhrGFa4zv61MI9JFOjlqD
4NlKXYYUr6UQGohnhGz58VW7SDTuQbGmyQRg/tJ0pEy+OUCmOjEW/Pp5/AFlVn5M
uQt7Ioyjwmewm89U28w1GL5Ut3drzl4GvE+fUgTaJe1oAsafN+NsFzXicBcHQJCC
qM8V84XOfxY+JGDozkDwIHbM3QleEdcHaEbL7wEZUfXMkL3e19sncHmys8kyLcFB
DMxbAGZvIy1e+Rt/GXh/6wlo7aKoSwHTaAjwIS1xkPwJ/Bv3z147qvOAqkho4gMI
8G28LniOQytjKl1OHZ8R4qCExg80yBQYwioA6oQkzzXQ/xEmbblwiDUrrK2LxVPT
dZa2Qaa7ftontV/0+mtja53tbTlH8EGhxp/tVbEGAGMifLDADoiebDM1mBBVSbnC
tC5UfYkOr9sCVcLcQO9ZnrQqLgp5teDoYgTF+/LQxflkemPvaGTHQi4Dzh72lAPU
vDta+yNxSYqR5XHOUOyIi4Mw8FRo+wze54csgiOfawYPcYgOQSiRDQUDtoIZ8+mx
Yh6OnPOY8ycgKNhPM2W98S5+6V0FvhU1GP30REaFQd9QJYJLWHGnQ7dc/8ewsbfj
kL6hCDPPDcoGcehxCuhiYljRvC1ETD5CFQD+Pk5J1Rmly/lbva0KjZzCdYjDYJ+5
ys/HwjPw9aNmCUxrMfTGMw168Jj3LjhscdALPHZGwhpRaBkPlOifmKq+120pjUQW
A834kzp5kzMcQ+OEpEi3gkEs+DyI56+FyodP52lrjboZOMtThAjoQ/FNlRbtHtlE
hF+yegmBby9j5fJM3LQapCWi2RRQ4tk+PKtkubDu0vtmbsOGwMVyxJOu5soMYIjW
3wvenIda+oCSI+nvx06Lq/UyiDxg05YNp3eMfYrPDB3TCK9zB0r/jwudsCHwh6LW
ruAabl9R43Rl6UT0dHYEJ7eowIJuJPvRYHe6inEGqBXNNpatfbK2GTaL8g87Mh9J
sX/XoLqNbNDC3fQLB81dy7xQQXrKmhtKoHBavnu8/6L9SV57yzk66qAk2bIvE3t4
DC2/fAOufQz8k1bL1NchmPIct72X5+yCiRc/oRn1zlz6NzRmBZb0kR2SBBgWYeXl
al7eJZQsC2UAZkbkiECXj6rm7Oeg10sS6DfXt2Tdc4CYctq7Pj0CcyS1xB1528kj
bqXuNOoAzU+5uha020XAfNvpj4ZSz99hrx3QUz9A47Ka2v6V+HlY0VMy5cePjFmq
z+QmPrp0ClYV0B34FtqM6fF4s4U9sWF78xnRZl9lCGAjJzN5cvWZW7PyP1ZEjRph
dlJ8SK95a0yU7F7+VDpR/VuqWMTlEFaoh85orGCb6SSzNLrpki4Wraz/pT4YwodV
O+aqN5QK4qyzswrpmnVRcHKnn9GUZODlFYi5m0lxIGYBRnuOEuKTiCjlsfTe7EAI
cciUnr8T7ySXHb7ifzHYk2XMH/uaTedJiRXEPfcWqiUm3Vn5XPCnc/XOoaVHeaSQ
9YEzoYWj9b2Q/0H8HFnZUY0qM58oE414Z44ongm+kllDwib6n05c+DI1AKYyOR02
wYNcYKc6WiXakujbbduSYT0jP1Yr5qzgstJLxvhzJqrGxZ5kP2QozKtDqXdStV4I
4vV7hBFvAeO7O+evSYsCL+zdcuKOCdq0XBhOfRwEydJ0IgtQHz9LP/cMwNlWdIHJ
JGzUepJFjD3GH//PdL8Z8OcJYpgGxMSJAytqvAeOgQp3ZvvgsmUsI1SLPZKiLsg3
5S3g3tR+PutIS0fIOdufHHuZHYMUU/4hCKbDUqeWaEvRU8KAU3UvOrrB2aGUhEOh
aTeZLWSs05zvB7t9Gm0NT26GgbQh/RxcnX7LbfeEdsXHtw8YxkqvOATlwJ1dTbDI
LqJsEERne2etAr50vWAlC1BxtUIqAk3rTjFQNiJb51KpoMymrOgzIU+fL+XZs7eD
BXhF8W5jzElMIqVAvO/b7rKyBN7MQy13aGx9fScK4x4YsTUT9W4Ic2hqZezeAABW
38jIpuKYuGRpvmsyVqCfU3nUOKgb3/OTXjvskrSkdokmNpMw+CG48FajspTgjAAa
jz9Y9sx843cyOX/2gKNHTKScf1j4zEbl80Xv9w6Fy2QCxETctCcrE9SVk/YicWGR
ECBt8DVSrVK6w18wcr1N4jDhig/RB5s++bpVMBkBzmBB2WOL4BNYD7PJkNYKNW7L
QTBPmuxRSFhZWOn3Wz1rpeWswEJ1naGamlMitO0i6xhqFz7TMYSCCAKHf+iCMJQ0
nR4YcRJPMDPXEy9irMZ75nbYDkyFTxLkt4dXv0Lj78Kz848sH3xMMC9cgYqJUFCq
T0Y7+wQmPk1bSakSC6PqR2JZp5VLGb1whojwuHaTtSPzEjUeYyLLiuU/NhB9C5Xa
52x6928SNGubKKlQJL80o6NRwVGUGUojq1MypCV/gjgMbxFoMzWkhKMMrG22KqJb
jhAla7GVmKL5wljWjagL0GSkQGmfd6C+FvAl342/3/sZsRmyi8UI51DjaQQIbJ+T
bNRxr1N9moUVgoCCN03eCBc3TvjH2URWm0wHQ43p7Nvlk85uTFXJBy7P7AZGCTAD
xS9PtgjDv0u0Wut2u6x7chgHS6LVuS/O2FFYkVs3czcfFSmpJSC2T012htw294TH
/2yIi90GdM+UouUK15y16PkNt31Ru+qwzTkgsEQwNxFOnJrmtXgnQHIJe8T6XlqI
PSe/x/p+Q1IfPlhLtv813SOsmL9j3vzV/z45bFyN1x4tAr+XAf/mqOkYBBq67dBg
mXr8f1t+NuQneV0DjuRCWsnIu4yX6pjPHeUyS0hsTpjfGsp9AByKaDj4hnSwIViz
rDYVrAI+1I1BgvdO5en1hLzsvxXlo1wyMKrIBHA+V/LFGl7za1RMOAP7uXGUnWY6
kGNB+lI244j1KLfQKUalhV3UDFU9nBN5t0/22zWCfYv7Ot7TLk2z4EFV9A5T8F8j
nWDpah57+Rr74z8loYBfECT2SO/B+54WAI/cQaUYNxfM9UKOuR3lT6twhC55gNnA
kuUXARSkkkMrn0kfFLsnrX3/TMSUCv872arz6b7o9y+7eJOyCmevxplo8GiJgffW
yyl3R1gpj8vT5yLiivewGeabAAeBg0cRxSr/AXZwVbROOWwmZCDj4ENQFpskdYUR
xwiVlnlgw0b8Tw5tmtIiGnZPR3zxDrF9uhLqjDBOK+3maqE/14WJExp+szOLU7tA
SjukUeCOuFg439gsnadnE9l5RqIP6DSOC0InFf6f6gqeldtiEiLOq4mNxlXrNeo5
+8U1/tjgfTvKlqm7Ud0NZYIOKGKhPl8kNKzb3He/kZ9DCGTblDXFvAPhzUCsuGXz
/cST6QdX2M6XliyB5zDv0t5nk4wASxys2TSiOUgtGq7rHRs7AvaoYCXoeorJ6xMI
MSgpGohFzQh9hZyRDxuPGpzfBa2tie1QtLtqardbCgrnhW1vQR/3u9WgfP1g1ltt
T6MeZqKvG6e+bPSBROVrutlCgaobTEkh6X0tUlohniskFyMnu7prB6zTvvdlNahe
pYji6/DDfy06s6CzlwGlC+azjoFz6BnSRJaUCmLS1tubG9LR9D0FC8+/SQKKxmK1
3KOv1NI6xfx7HbxW6d5FwTDODT1ofKIjScblj1RO8VXzzNPbMlEkNRbE0WE7z2IB
+H+LGoQUSoUGTUGxIDX+i3nnYetQGiiC5c7fZlhocjH0Mh7Bd6X6NmMxOUVhfn/2
L93f6Msg3BXc7bj/18GmEJBVSa5i72uw2bGbWJV0SGQTbQklwqx2o4pvtrbEUbfO
+DaIqll2mlokRrLNWOlk8s5qDcAna3keL6an7A6MhTKk7FWTrweje1IIsFBi3S4u
onlN6yASdGPdh1bCiU6JgLV8xUJWb8mJJEJzWM8rNIws3x+kn+h0TvRo+QRBie+j
N5lQ5vQZM2/Cm0PWhi/u4NCS2vIka2YPO9KVmuAO7pMIWUU+8S3w8UPBs+3H5B5c
BPmoJHGcpb0uzlhIUA1KVwTI1hpMJJQfXfQMQ0cWkzeoQSYS/RM8NtR6Gvyt2OAO
jZCsc3yZZdIloM9BgoOjJBTxgf+wsiKBQoZt3z58DIO+QVbGfUweVpDm6unp1Sff
ABDUEyAJvbbeRySFQ1HRcuiGC+AEmsE073hEwpqm4bedpmVAT0ZcOS1x3weq9vnx
qGAuKZS01CRnJCvBEd/iSExTTk0OeGgUjqMjGUv600Gu5VEZD/yHtSwAMkRrFXkn
khXKFpNrpEn1pNXEf0YPbok4hzJ0NSbfRb9PNjzWhW43YxSCcUFG4LBugJXpW1mv
4gu2yaV19UvhB7okIwobvtoU9P6E7MykrvnL1Q4R6SsUY7bVg5XFW2Bx60PCCjIX
AtYuzHuPuKks1rADWZlo/gjdqAvv0cYKFQ/hlKveA3wFo4EZDUv/WmNRpJICuTA3
XVYnP3NS7RzPT81tytFqADk742e8qS2hRJAdUhR1yFgUZBsmtkWNmkY3oiV147Sf
UDAme8iTTMmHv7xCFdRSNCOr8LCM6nhn/oiSAylZduYl6Gif+VKukhvhIP0N2hn5
q+sVCAg4NxKN7kHyIYkKFA+gTjf04cG6NOp3lWo0FCxlVdjI0vHHGdayikYKIaSi
+4snZaJXfDmQSvr0Z3f+DONBc4TmTlFBs4IwlujpHtN6AQIe6p8ww6k90Oi0/P+K
90YWDAYa5OYEIYneVW6Qsix7F6CRTA/ePbP7Iz5zGOwgALFbOvOM2uCbp1y1TFsG
QQtyPVzvNmfQpBfFN6g48WQHniyAzv72+yHLkisHRJ9mrHMNne8LFCE5xd9xIOWV
pe1lmarU7D36z6ETiIkDZ5aL5W+RNNdB7AbKDNhGL4lS7OciZnJgvOEGY8Wg58ZC
CiCaQu0JVR0s86DZzfesd1AX8G7oo12SNVq9sqzEOZ0YhOIkpkzhKbhfWuYEaXx4
9pTXfmNAnkHoqlnm+tgYJcAcD1Js8cUENN9DDoE1+v9CrSIL0sn56Te0mnVl1tQq
B1hvSmpmtc1jcCADBnXEdXGIpNUwG0dmT6qd3DUYrXW353xJfaE+QSqQOtNtSOdZ
uYvTVETDv2JLrl0HquXx59RQB/OkFE4KshpjnSC38QyHUUEZOtIxWcVqEvvrCKN/
SH8rwKbl49u0RsSSXumU2IcxmXZ990KrQAbzq5sz12QPOPkBZ5Rp8wx0hOKouLfk
cRkSh9NTVvZMFovwIQTtFTERYAHQq8EcxldxFEe9Mn3bYL7arHE+83tZm7QcZ+Pn
NofKPTe5ftTKyu799RwwznXLLPITT2qGnWZVgSrSy+7FVfuYf+IwlzM8f/QdSPc2
U44h7jsmbNbZIkuTJsVy7bMsnNmv11ZCwwidlV6E7b1wM8R2fgb9yWeFOiU2ccR/
sZjjc11PrNCKKqXwQqUYIiLbsRL+ER2NyIfCKh6/KHrKMaanguQtHzdvnfKuYpPz
cfwsHKUMrMiyw1ozGFByaOZWshF1efbQepsEiQR18lCFfNEf9N8Qc/shLoTbJkJ6
n80UoIcgkXaDDbwb/LGnLWlnh8ddiZvNWA41AJf7z3qwW7IIBGsyGrPO8hSe6k6h
ChmlyaB9PxSE3FafeFMWdPATlNuqE8nOp/fsVBtJYV8w+3kCswgLz+cA1kC17YCi
67l2Gll5pKvNzrl7vgwB9V8RRRyDobMOpuBRAvDAkbDy9OqOmo927wCm+Clapcm0
UHBKS1Kala4MOveq2TNOAdFX3h0q1bzy0aPhuhmq4BoxcdMy4Ws3B5fxZJYtw+KT
aFdVUn13r/0u/bu3b1i1V5xU7RlATl1h8u8uo6YWL51prq1zaHkSWptVPlETsJrJ
ecAoXGf9AlMaIh/5gufGrQGOw7OtOxlKQguQmvh7AJpQKk4HqILhZSSzAndo4VnJ
uLMMLj5nk4bHdx5dhVJ3W9EzM0XBHyyqH+U1oXgi2nKuEcbK6wcEaw9SbhWvcKj3
B/X14WTDzZflfoSJ+IxAGv602nQ040iryQWP/GUWYv2ZZu3Xf69HXTW6sxA+Iesm
1SqlPzR9gF6AYuRGDWuxL7swNkqgImwhukukA6nz3KlclreAV09xXVQLo8XHQQtP
shXLtwMelE9mwUwfBNugDrOmkL8NyzBxoFzfvXBZj3kcMTSs5oJQbuof7bUXpGFK
9zNtp2wyTiUMnUxjH78CAZp28ua+X/zrj1oAuIbcWI4SXx41v6N3WDIIRQs7l+7u
pWfxC/T8tXOsH1iv/PP5/H4soHeYd6aewdjgxiYTJvYVKCWl0nphmDHymmH3io4y
k2HH+HnWZm+2g3hUyp6QmTe/Y3lPBcXDCj8B6jCaCg8PCCoGdnunElNWMLWxmSJn
OElmafmekqp3RhaCmk5YWBooTqEdFTorUf02aJsuf+nHyj0DcNrZ+uZnpDD5DaZC
imeboGW3HK7lQUlxiLHMy0lcVicNQHKCp/kbHomG/Dnqrb7ynkwKQ0peAEq+ySfx
FUhMRxKa0JStw+CQdujo+k5txu0K5o6Uf6051q2kJDPvm9//nIgD4q84Vh3JzDpk
uLKWVCXIy221ubTjkTppGxLZc/Nl/fAgA3/vtKQ6ofkp3MB2+LGdHPDW/oJV29gF
e/1fuBNh2T901DFuA4tY6nKbkS3foQbFDehZW+msNjBFHA33gq777NgrXh0hXi0P
GcPvD8kMWNdRypgV4sgKNm6MV9GEfEPOy2l1C2MMNVur7XiOV20bEvGRTjKhJ/t/
4aNSCc64/3FyXUxuw2ZXYmLmEJA3fZPGHL4rsD9po6L/L3yGGTJZRxHrzB8GT6Cn
tJR0/7rda2CHjrQeYGpCmMoXniaHSBf3L5fiOj1SVtApxtQI3yy8I/gERFGHKZuf
Al5/tZ/GGGZjC+jMTacgNx/mX0wmKM3E8LpQhJ7eS2lzxcnv21n8fezm0PlrCcNT
uuDMytKBlcCUzj1txHrQhRJb/GcU64sxfrWc99QrS9MisiFaqVdyWk1fNk389rkP
wEopiNod1PLD3OiRn0sDomuApDp/B4+tbv9aLEMkjX6njxi5Uoh9uMG3mqqsDP1C
VyWaUuGrZuruCfZZ5jxjbIneX9tEOMVC9L4YNrPpff5kWjdY26v15UZWhWs0dqO4
TvL3xNuEKtPTZa1CCJ0ERFOeHpYenKWQjOgtJWvYdamelR97OuiXZ9J1XfgG56nf
s9Dr2MIyXnuyQFed2urGJOuZb7KblbxRi8AbnWel1e7dag5zx1sMiI7S3Dm5kAiu
sHqszmtfBTexVXzRBxtG94sbVl72z7zSDJa9dJpWaL+Y3Zz3FfGJ10/OYQkGhzqI
DYaYr2tKG/vA6zff8b7rGyNMXP4RbOfNA9JeVsVjH8tvvR+UDDxGplFcoGQQRO0P
lWDG8jj4NNqikU1pV/R/6k0qLrrqbhX+SIic6RXgMD+vcO2MVijzqIIv2kOejdQz
JpIK2zEBjrMcYB4+6VReWTVSSBPymbieeD1rxyxhqMzCa3k9JFlVEUZB27XdliQ+
r05f8Xx5Kx1YKlTs1plZhQYt/3EUTQI3aRPAMB0R7t4FRWt97+IDo175wnrQafSv
aN+3fnhV+czIZ3kMyAvSCMhbhBN6U55Nmhvsoya6kpkI02gitgyOnKvVYwR/Qa/Z
RUdzg/V6qJ8aBMpsPvPi15xKpQiHmvF6CUU/fS1oFoixPNjuf1UfkfFqjk8EE176
0E0ykfa2bJHXZ1K6q5X0cN3wJxB8nBMcD2Kn0EcUKSAnLX7i8GcN3PLC310GeOJr
RMk59k5gtjFv+KJhbn736GF+NvYYdjPwBWq1+MyzQfkRQr05K9f8RLNP1Mtpbu2V
zsTA0OL1zcLOHf+VD0XlCitYMGuL6u4BFb1LodXb//ljAYxCUpqg7B+5edPfTRbj
i+xToqOdJojtoBXoSAhJL9tm+yZcG4zK3S+bB2IK2rGChjzJ7ViMqBvtFJnBEYBh
Kt6csycpWUYSdDOHopQGs5OJXQPacJFkb4x3zc934cISmxrhroJIinvMy99/Id2w
RMphx8bN7C/B6pG1VG5DWdepIFg+gEmaBUe73QNlPqrpjWtfqqak48CAmHzYZRdu
7NwEkjaO4EKrQpx8/kSs0f1Fa9QyEoS/DLtYPkQ/QZIoayvs14hhP1YxJEvIruQ0
grwqSaH/DOZDolRJGxgaHNFEabCzspu7Opior+FjsJ9d/i1eXF8xe3v8Vv+8x2C9
yWlPJzfisGn0Z2Pu0ibWg6TmDzCJGnF/Utxu7VdM88eJF8WUA8DJJLu43QoPm5Jp
lSTmILUcGUm+AVuY7N5hY4mgsZ7wHRy3Rvdxx42uGzu5+OLvdJPLCCKBAjlOz+oo
IanFawOjflBZ6V21soKAqS7qgo/j1+oTOg6nm6NKwsKB/UHsbHsI9mvGXI8kU1eZ
bQ/UkUW6ScODtudg4uoLS9QyP9kPyezUkRhuFuZyq61pU0ny44rR3JK/BQXvCF7P
gDuI3bqRlhxneet5FVnFLIbnBaICStb3bmCD3ieB1hKoQzfA0P8nNLWh50dV34Tv
QByhgOWjU3mFVTBOlKMljiFLhcYV213kPnyjk3BKT36sqJJ+TELPjJw/ASRzxOnQ
+jQ7B33rvylTstwIZJyV+auxy5B+8Gy+XFWQDq2/Y8uWAKQyVIizCi+lajwnjKb8
ZnEDnvPYp1A9IB1xQhuJ8MxO4chMZZkvi522LRrXFlRl5kWnUZL+TWxCsxv5SbsR
aYuXuFA1uQPdd9j1WVeppF8l0juZGdgHHwTVQE3PvhdXRy/8C+IHiY9i8/84bn2x
6gTxAz/31hwMwZ8XMZUtdF3SMXS3rnOfLbPtvEHYO542RQQJwpy94iF2Yle7lS4D
F8I10SvBK/O3vy0+12NT0gwCr7yYrErfbi+HPurz+m3d2Z2CCBPz8r4hIk55fUP6
akiOUDwDhEhZ4jlNYxpxcrPQ9X7KXPE+n8TVeA7MnmAoVRuQFMNhxdph6rI3JE/3
jheWhHRJAvdjp+Y7uEiwyGgZjfUyR46kvcURIgpjKeobVl32smqEYC84WThRlFQA
aCRFJxPoIAZzQWBmM5qGM1MWeqZ3H616gPJ8MFsswTNEugWwR21WiJ06gLmF5VCT
aiYP/hyKR9ZDmuEfW4OIvSBThr604sS6cNBzRnb0prwVwPXab+ExIJaPXtvKDE41
kExsuJmZNkpNnDKfvC2eu4HORSkPrD7dR5ibXmbJ0CUpOFo4KPDsHKWw+rORfQI8
EBTOk6ThabLo4MimoIUbxsVZW5oV7tupHghgCxaCULm6IAXkbgI4YbIfjnwq4PX0
TQ0B+inWWv0ujbZsOOweO1LI5Hc4A1p9lfRV0zCYoylxeoMqDtaBvhy4amtvXnp3
rzyfys/pzil6WH0Ecsuvd/qIOEVQr2q6EWixwdeXdYARJbHbdfrcCw5+Ep17AKNW
Ssat/cznc7933Zv+T0WKEmXHW7THTqgjd0rdAX4nOWDvNB8L8ZhEcPrtluRNtWvS
yCOsCU8TTvbZbzqB1YGdGBVzhIKKzr8k2ch8W6xlbQcbCOzqeID3IVOWoEmIddzD
loAIUxBhaGAEn1YV8zVJptwYoJOX5iOrnPHrOcwzn8yY26nf/07BXc6A3HOrYo8H
LWP9toMMKu0c0eoaY3hCqx7upxMi03k+LtyZ0Sqys480zeL9E6JxjylAt0G/MPjK
+Xgps3IhKZBsuND5UG/8sxw3igCcKwh5MHTbnC+Ob7lEHot+2tdtZewRJCmxfbXp
69vQcdflXkxUw2SRa8hMb2u15/um2g/AXKmAD/oVVm3S+3MsZ4M70Se4B1UucCOx
WmmEvF2XsozNgLtu3eNvfDFigWke9PMhg2k3s/QxIr2q+U1wJA6LRNDVIEEsoyR7
9SZLiCjCk6USW0aZ4eTbV8cDqKJ6ZzVJMqhUWVd0YtiDZ+nHPEGFVGGrkLvR5mSh
gT9cCCkKFi2ijpn5A5rTqblDjyJkw13G3wE1zTwIz2y8pwgkysENPR9wDKDn/dPi
stGbqJryKCc0mNIxh8f4cW+pwNzTK4VFSJDBnbN/6daXjV12gYZ26N/wEF0PLSdc
n7AG/59EAVuYdY3Aflb2KasUYMK4iFtGhmaPW/txMvIhF0PyWgEbGbIs2aquNtUn
sucUnasbOoc019kWJ62xv/CI4Zpc63OBVNVTK8+xaBjkw+A0H6ud9gFPzAFhvbxi
wXalp+1JL7PdkLGxz1k4couyY67JqVSkOs5qLy7f/J1dUz9iCWQPCANVAlt8Bft4
p16ATnZoHRGmmcflZaCUKpjf+SlrfA8GUMjtOpyfJhmM2A06NdF3gT1DuKsSjS0t
0kbExKf9vsFrAfrtot59VlIs6LKFWoeGMWeEBqaTghfzZvmRXBMm7xx3BCmxqDCu
2nwoWbVxBhGiVBPqLhM9SI71norbluvY3pfDjddQonjhJUuK1oF1rhcxIhGj5Z4G
Y7YPllT4kAfcIxNIeWb9KQWzeGcqdlbddgWvIJadhIcXuEpq2LwvRrFUUppi6lnv
7UCkESSHMQKRGJb3cK0QFNRseWLoFhxXrmSwnJwKtKGm64sdsC0QwPtjJUTYvCXD
0xA9NsrdXuiVYztGagsf6VohhFogD7ht3y5J330Zt/oEmaVR97AYOR+KxVok2Fx0
GipuKefwB7Ncf/vbrQpTwsZOhMSJjF+jtzI/FrkYd4uTdL82UUOwD7TUDefTKh9V
txephpAibmAs3p9c5n+OfYgWZJ3ILWuJIEr34jKjvqExsf6Ow5nDqhp//jd4pqc5
egfLY7Y6+eI4TjJB8y6AyXy9hy8SmPtZ1X/5CDV48m2c0Uv0aDRI4XjStJsP9MX7
EETWppw9CEJPzxUvPvMWbc8VHE9cphCcEClEI1ETzMSMiPldK9wsyFIn61vMeicH
DOo0Vqo9W4JglwVNV5/Grngw2HppaHqLo8GQI+VKnqSl/w+wCWpz5Em22jyP/6mW
Duaq4anlHDS5NtaNG7U3t/A9vDB6mkHL6JEJjC5PkYYhZSK3TvupWvhEZgazZgjp
p3T4nnWbsWXlSyv9yMkZW5VZ/6gZieQrUtUFfck0k6oOZ1h1BPlLjoYZbr02kfkf
kcyQESkB4xvU2qTizMl+KoOUOB4y19/dapxhaPWWmTZwNSqST1Q8Qxcgdf8s5r1G
YpTy6qKG0q7kFujfKfQmM/FB1nEU4lJRkNm9gPCqoA3ogwYkwBxhK1SJeikLAFl0
i3Jz5i2zEKo/SMmLFR2DGJRohAZX5VFJAaSQrRDIMj6RhjtKkZghZ6qfYNuAawtQ
VE/aumT0W/wnaUJMXO3OBqYMNqxvP3fE2hKhl5TCIvamhl6NvKziMivsw9fZmFLk
UfEUD9s9lqwYcc0N5zlcWE0xAikjthHPy9yuSvYJ4JJA8t01LM4Y9qingcctAL8P
JT3U6L6QMTrzoe9NlpQy0mx0K29NmWdQ16nQE7yNeCrVsryX9OAUtfHJvmVUKlYD
rsPJFx8O341nxCGY1xyO1aPsGnJ1mMoJ8p6OK+UJt0Bfh5yGBuDX0rgu0Isb2OUP
T9Nn+pCmSGnabtF7CeI+/Zc3T6dSJ60LKZReEbHiAoPlnKIgHO3elfDwzHcRktQU
wB98VjAuz6re/iB/vISyfzCGoIvCv8IVx24XWxDVZnwJhTXwKiDfUumky5yA9LnI
K17e+3ojv8WAHTgHh9YFx/1+lDaVOZcN10zUSdW0zCuuQvnQ5JDAcY/VSba1dzJB
XoCRF1WD15fKF/I8fRcLsLPGYmK9lYO55Sk52VbRsUSHEn6YqqymqhCK1Or7x7Ix
mxoeytVCquf9KK9ipZk+TTa0og4ZGUQBivB53oERgmcmivPqEbl9dcfldIon7CJ7
/M8lFSFB6mqI5nY01fz2gndGv6qeFXO3weAvuKNt4Z3A2vXcw166omdPqX0T3shX
XTSdEsXT5nBmmC3K+gyrarUETx1g985HzEq2yeiH8QU+YbZ5r/mzkVpAWVZxKhv2
y/6IliQK/ReKAG+NPKrhHAUYlv6rjfu0/aZI5zxgfXm1t+Tp9jXhD23HJ+xU2IJ1
Fpu6IIucOb+FmHmWddDXgXBQRHFxt25qj19Gn9MZ22e/0RPvD3nHHeb16RHGYkzZ
PtCNmaOfkyuvZvAHHpkK1j2MtCVRnTandXLCJW4eD2EEtYbzNjBLX4PT76IVDeHm
ykt+yo6j95E7PXex/xVrGjPwb39xYEUIOK+7uQjY1MWLceZOMkmlaqZo67JNq+lY
IlnkBZfK8Qabnl/rucNq39NBj4DsEA5AOzctNVif5sILLtjw6Sm08kc7CoAbqTfz
LvygG68suE8U5p/3nL9pXm4vDaFB4uvvaiGxOJZCIUFfdwdUUTbArQCfhIwo2R1a
rfv+LoTz2mg+q5SYkr6iWjrE/8ORPP6AiarSFAXjaQWaR43YoAjDBI9NK4fp7otw
QbhiXF2WKMpJDDBEkKd6RrbjFxY6TO9LFco9C3nK3qmcMcfBZ8yTWn3g6SwbQcpc
0gUoWnS+sVnhFMl1JXU0IxaqqTyhBLZAcP8rYlJbx3RHIm7C3MLMr4KfDI/OuteV
SGApmpugYw2n5BDqZ24hWDw+TrJY0NC/SJfLTMVczgD8FlxA/Ym1KZUHB6EvrPtJ
nEtwAbYkycLMam67L5OHjGhE40JcTnQ9RsT8QP5Mo/HP3Jlaz940wngTgtT6nod0
d3T5IYN/ZfZoJWXFT2rm50nkqIWHgW4C1zIC+KIDC1Y5jxE59wpzNqSagAhxQAJX
NxNrPQYDhW82y6BEVfmTVzMmcUZhm2VTYCiVKdKYnRmB4v0RgCDAFfSwFRKZwjfL
c4CwqGlsJK3wQ4BZrhqdwjJ5tA0mHi3AXE9JjqwXILvusY70JdjglTP8qpk/kBmC
UH/mxUamCMAQYl3APF4Fv/yflMmHEQKxWhuAzEzlOweYKcJiDVNlulegUWr0870x
fgJStFSCgDzHS5QezGsTq2DVL7Ka93gCkMLiiVsRWJxvWB6o0S4zeNBxms2h/8iX
wXhwscZKvLS5CNSNfwVV49dgyuRT7kQ8Nj2AsaMAVUohrlUIEB1QP/g1UDTtNT2k
TmnKVpDRZ2zt278r3cPop1Xw1n1P/5v+Qd7GVDLrKGXE0zwv9FMQf4QkynVDRQVB
cyqkwLsKUCTCniMatcfebiqAzO1bUCvHAdnA9bapX0aFmYpOw0KlOgUHXzWyK/fj
B3jcaBjYo8zU4wLzvTz4MrLdmvJAESW+Ea5T9Cpf1wFItmx6D034q83fo3eog05E
GqPCrRYAwCA+DfiC+91CS4sy4Fa0A9qgt/drTuO0KpEZkub01ZdHoY8ztWDF51FW
emiUDIjrQ1oSHxLpIOYj+f5CkoUhTXViOYQanUwj2tlp7CnwIlKuYJ5Bg2Wla4G7
oFaedB4qq0Q5Rn1Re3U0d900iXy7p9+a5GbFqKuPVVd4DV98CAPItnaB97CIEnhb
2HT5yYkTOFR55dtBnkJ/Q6npqi8bpf+1iSjuO0XEJ/zGFIFlqNn44qTGS08JQto3
dBgjags191rkU1kIZrpVrMF21edjxoWw3rB2gRijp68+hqoieObE+nEh+88etLLp
4Vydz+pOG5XnPPWc2uYV/BSwXWN6Ng4hmqcI34t8WT0bSepvlxwd8qp25REDCNSU
LbxtFpLmiN1ozr5wCEFYunP74y7EUkbp29ljG+2VsKs2rbixY65eV/X9L7JkNb8H
kxhg8BiFwmRtHAMR/oycfZLaK/hIR0qDSfeZ7QyvKVen2JFNEw7fJzYwnODPJRNK
34Woo+IFuB9ViQSTMVbiIDSxYqURWaEFiaOJkIB5YEGrx5DvyAV5IqpbYADoTJnt
xEsY8xpwYBGVrjHAwhg7FVwb46/cSuz/ZdldBzbisBIvKpjLbAvCfhdDtq+O3wcD
XuF8XtTFJIV84wtz6h89roeUR4070vAWF0baVDWah37WQLYgrdY0OzLm9FKfTcXd
8+QbQTkd7umqbF6Q/rqloQjhoXMJyNThA3N5UFFHXg0PD6KrHFgswVqCkA4FT8IS
rqh7OEjqccgoBkDyUPFVE4bKXaiKGbjCdT97qZwHFS8qd1vB5HfGVxo7mGwWR8jl
AW+O1QpZEhdgnVIMO1OlLjwYasBKR0rgYmAo9OrZFZAHAo6IlrXfwbc8yULDtRJg
k+Iu5uw+w+r04uE5rQxBWixwAStPhxErrx9NRG7Yh4FLjfXuK7rgGVCWZ1pBqLq6
K74ISO+za3Uuu1Km0VDNM/g07sNEVSyOMkeI0veFpJMUyuUxd1S6XEmzHqbYkn3k
21MCg3AnXWT1msjyEYSst+rJke3NGnNrx+7SFLSRVYiqjp7R3qIbnnk3XjFWjoEF
lcOIVAL+K5FVxKptjkCK8++Xu2oTfSXKVxGsG/soHOzk0gV/2MQkUz8+bqQEBG3E
slhmMENXI1so2+YDh1zoZ2+wxh4WAxJKjJDijW9dTs9WSfLAnCbEkt/k1nlWwPKG
/pv8U4KehvFrYva7HzNo/S5iEIeVWLvFSRGwmuN4h6hFb3eCXvdGDTOllph4ZbvH
7UZguXCxAnfRJrK2SSYNr85/5zlWNiPpCt6FxmWdWWw/JDLCVvu7P0uGd5r7JFbS
K2poJ4JHniox2hurOZ76CyndMNb0YkzkMCcPM511MOPVVmTZX1PHkMTc1voYuLEA
skdW9h+MbigR3yKR7MVD0N470TwdSgL0hfU6+SVpmvBpLywHEB8GecqCan7B29ld
FG69jv3j/xRGvyeWw1C0jigIXNS3OHg9QpXkmcmsyBDYya61JVfVuQVvwDEJIgaY
ZlUQP16yoETVSIpmKSg3CtAAODZSp9yAHxuIJEO65uC8kHD8SeB6nXA2mL+J4Cyn
KeAw5lvef04JG9wK6MkJMXYcksRlinfPBhJdPlwI634IS+ySPSejfD0VaeEgVxG6
nIdnklFDZ1n0082dZK9Oy7f6ZmlHppM0nGP2CyghR2UVMloLWIEpiHrdCJ+o7QHR
KD1aIhrPx5aWTs2Mp7gPqV95F3R+WWnqoO0ieXW82S7ObAezvlvLh1wZRCwGt6rQ
Se2nAz3iZSKq99JQ1pR1+WOeLj84btvAOdEU6YSMoHVlNc/UGCXpQkQVGtw6IEMO
F9YIxbQ5wxy1E2GagfEqGBHUyey0C609WUxlQNtJSJuf2xWMTP7nABwGWQQBYGW4
SvjFAyJ3XZkVdElUhh7ZROrn3YwCujvuDREubOJuiWQbjqbbb3yicFf32ZpJ3u41
hTj9kA3yqI6ZSeVdJalilIS/vIekDUBj6o1JtESuPNCQcw7ek1oGNtCN2Pr1a3pG
OKgIJQafQTLaMotEVyPHMBnCsUmkjO2Zc9MnLPKnT6/Wtv4XImNp5K6pBgbmkuvq
gL1glEvVNy8zN0xm9Zq5XILjRwNpENBXnW4ptpNjdz8vKvnY/udIG+986BH8m7Wz
J56ApqqGAv9gMTc9hc/GA98p/a5PSv0vsRdG7A9PJv0vOOtKpWKNxzq+BLnfJnZx
XXh7tjCOR5F7yWLEDbIQlaTJH/x4XU6U9/zMRiZD7EjoXVaxtqciieLMpd0bsUnX
MVWeyWUv+t4GZ74F2WAxp4uUKuIDp3kL1DeqsSOq4kBNwPoHhu7tNe7jNo/5WeBl
YFh3y+bTXlfL6kSpxXnY3OmQ0XezjQGS+nR+xIJ8UJqLSRipmUMonTO0tUy3TbZ3
V65mbkcExCX/E3HUj86Y9VTbotLsDsOhBH2520TGQdtJAp/ZwYbuMHTzfciFHbGa
Qh8i8Ks4hhEOnxZH7YMUf4xNusOd7w5kKmHclhFcccHO+iaDV0T7ghBXN5wlUjW+
nLHO049++zGvapgTAph8v+eAXYl8ySbEVvayUlXxbLghAh8j/R4AyxZ6wD+IfAH5
c0gSs6llg5C4rHBttHVjSJuZb25Gsvt04W3s27fy0fur+dDsIDWjAU2fEy/NiX7c
nTuh4LwdfnsLsGJ1e2Rrg5/JiORbb9CUc7IX+2ryQRaB1cI7ujy2nGxpa7ccIkiQ
epy+c/sJ2FziTK/P7/R57qDukrt1l6DfNLF7k0gyB/9ZdJv4Hm4dkVI52DMGAGjJ
Rh2CCpgUjL6JVqUmtlUctpU/psIZDXE9gatWJy5qYEBaZV8e8vrGLyt5oa+vyqMd
hFtev6dkbWzxBnp9i7B4DbFy1x1YUt1YOmq4mCo7xfPRL0rWjkPhh8zgVv/+aY3P
QlSSVs5iN/VGE8WNH3dhUnRRMlCYswIGi4UqDmik4KzTxVyv8Y1bgMrMCTBhADLK
0sVASyaAnVV51ib5mRNajSQWpYnjUyPNhH5RWnDY0teHC58kGCexEVoaDsr2K8/d
lYxvo9drN5A/KSkq8mu0scCfQgMCJ9Xs9fDehS2btlAKLNPha8yA/z0A8hT+d1tN
mSHDfa2g6H4NY+mvibCatRr14uRWMS5DYJHkmq7TbldT2gk3wQPoWgHGZDN/U5X1
5YU7mbdcnh7qx3Y748UoTa1RC8S7JC/5QA9JrcqFloq5l9xVwEQ3a5xMo5A2U7My
fqEsE3u5xSyi6UAmnr2rBlbYxy244ufejlNeyXSUjrr3BAzctL8hu21L8Q+SI6fg
TJ2jtbDYb6+bwwBTMMyOFiC9tY+/ZlDN5UikAdzbLcHN8ME0GrxLTdAWbD8iAUJy
Qzivl6wSBTclMlFtaYyHR8nFvI4rBKp1Y3AS9jBF2ZTzbJBSKZOwkmVqu+IO3m+J
+BkFEKfyF8BiM3J3DYU3rnoy5okRFTg3EftaDcrAPT+Nb6u8VMdyfzA+nlmZCOIZ
k6EU8iPtXGR67Q6nJo5OyBgFL3IHgs2jlj9D9t4F/BKv63DZ0of/pO+ftZWnYrHt
hZ8Nlj3qVWx3P8cXedKSxNnp9T53JOBBaoFW74SlDixB7kL4DzK1cAx1CDZdOcZx
SZ+8PG2/uFE0O6xmmLVfE7jls2Xx2YQlHkbIfPlfpnkBcFn0JwdIsMGBoNzwkhRG
BIBMd/4PkxD4zJmBcvTd9PWOpqkoWrUms+XkLE+kA2p1T7t25D/q/vzODzw/CG5L
P6OOtEUxepVx8po0zRnVXRI4sg7a2Qf0wnhLBmOjslFiYxjgZVerQtnhgGNe2Pwj
cqaWVjwtXrV488Xpx2dS3hec7vm9ekILJApiciOC+hFhDCgWcE8f2pPQFjMHlD0o
iJzyf8Stq3Rg5KON7XgbKfsRXi6KcvZrgi4TBpaZFpgctMZgRLmqPQBIe/eoxXVU
YZU2/Vb+LM/aSVxzQPOVKlR4Fmib+VCh66PCGFYdnXMLCMwYhTq4eGjuyX8iTYGq
PWO9xZ3xZB8cLZnHlfIQMWkbAFjL4yE+VkkUfBgkBGhgZqfy6zDxTujaO0VLf8OZ
c1nT6jgFBBHC3Yu2CrelMcLPEVBAsyKKaxc73fvKj8Y7JCFgQnsH7VETOIcELX1i
iOSeFQkqJz7b0cFMhzmaYrvv+gt99aKtkfvtNqAlXQA7tZ/OA5uWLI9IZE/T7QVO
o4PIHwxGCtjUel+lOB0hoRnx0nmqp/ppGqX+YzZdp4fGuWegaodL4mtRdKd5xiLj
v4CY0cSNFchtwnOwuFOk+KFFlsptQXk8n1ci8RmacQv3yCTxjUrvZXt2q59vMBbj
lciv4rjvr0ILfXtKZG+0Aq9q8ogPgJ5MuM0pDgjViFw6m/MTummFXkMYHavYlHpg
MawJhmQ8ML1mnDIV4PrvtCzkvZfGk7GFOQX2lfowrFezJ4bcCqrNNWWEDJlwE7iQ
slZnqql06WxgRfmq65qDcRnmFpPeSZ0wmQsT5QS9Q68BD9n41gNFot2AY9fCISLM
hme1DUh+YbXHw7Y8hxJcVbAaVb6Cvj7l+Har1fzyNxkyAXEzABdl5S7HM3lb0q5U
REL2xBb6dwaADtu1B83IQFX5bL1GHtlZ/C0JdssS8QOTh/eriC+iCsKgRwDHJzoo
AXK2UIsJlFNCJiTcudD9SkRXScc7qPG9PDhMeSFsHK+bra32XcQ+Q+V733r8Dt/Y
DsRGZ/SGIWuueyptSmwShPuMAvQs5QxqJ1tlo8fDVpUGh5ibAb2tZEU4VAvRhuh9
OYqh08aAv+NVWgWiY0M+grffNM7JPsDPz300+7zKVGzMCUK2JiuTSNluWA35FzKo
3AGlpSpt+Un2dKgkUH4FUVLor4M5NeJuLJndEf6+8TKBqCKHBQVu/NHNcdJR3mxk
uR4Ji7NLowk9Yh9W2nVy9NlrTV0xnABQ4Qcuaek/1NCY2vH9pCeGJCHutJpj4FVJ
YJcH/qO0BsTkU55r/GoK9MgvL2+AXIjeDq1MNEOymvuRAJIC4if/cxy8y/2CfMVJ
nvGhjT5EHcPlbOAWGwhfILpsRE/g5/oF5n56qxmzRCCL/cNghQuckvt/GGcHAmxW
K38Xl/idRzkt26HIKbZdtXdKlS8NtZ7gBjLfl3DDpwwTczgUR54q1IPqh272rvBd
JTL1K9LyeqlIoGCYexfduA47d7PfpAlxGy6yXIHLZI3yxMwRx7cdcJYFUIbMWhsk
ywICnyspmv7hIcS6CucNBge+c7U9rGYdDKNshUkqMLgYqEqnowPs8fmzErAkQxCC
C2HGO+YW8KyXo8Ilx9otPhyN5tH60J6DMC/WAlvWH//6DJ+SsE9fd/S6SMda9+FZ
8hMz73+U0pZmTYVVhlSJqE9yRZdRl7hQ1on8Hcys+H+G8KRmkeya0pPJviG+dl9g
IIG+EAAOvjI+FbSv83ZTgJg201B/hk3d93/831ow8v3DU2in/PRVShW51qF8GAS0
DfjJc+r4e0Kid55i+C9orKAOL26FKb8PmNbWdyXduePaZfZXMNsEmrHgsE8o7ZHR
d2WwFL7d0KL3xC/vkVoARMbVZkCuej0QP9znkAESRVNgMqs+6BZXWuoIcfZaKeYh
3idVUvvbyGPEFg3T/z6n1xeGkQ2Y815UDBPJckzGlqzB4UlM/HRXTfqcVJlZcTRp
sdnQVsOl5E6ifkgKwtrVVgwgfi8A2kvVCN5yGKnQpJa7n7sY/PP20FTuzeQSaave
z2IBOgzFHW4TBmc64FTw/2/j59F188vYDr8uR1DNpMs8ZXz5N+cexgA4SH9Pf4F7
oXbyDvVpJaoAFZInhVMfUCnTVKWA9ZUsbfqZRkxCEkdu1JHbtoSq2MzCoMadKokD
DUG86N0NCo3200stKK48VbSf6DYWI0yxiKJDJEKs0dq1i+NPhUdJaAppLjXMSGS/
Yb06OssEPKhgwejMlkkqOsjE9K9adNli3IZkprDAx4wH8d5QYcW3g1N4buh3JC1D
cbWEc3lp15Yeurv2C5TpHCDwwPmv0vZweoGRWVTg/qHW3p8MQG80Cqw5YKofXp0O
oyGQrKBxyhSr4rjdyTm4+tTJXoLiz0RU8PiTsdFBzgoqhGA8NXTWaQ9+dK9+g1Gi
hT5ADSUv8IQBiKsTqH60n+FV28hqangCIPjlym9H3XM8JeYc2HJ3wkHB6+c3f5s5
6tjJrRiX9K/eyOc9b2f6M6C4Q9R6Oa9LnVbfspuoITndkouobbHT2cfi5dKY2YJb
uUDpgmLmksM42veb5Kc3tNYqPUcktN+DYHy/eZ0wG7kMzFpAOQ/s/TZ5Df4oqzRx
YTSjkbpd7w3cnZ1cTxLCn75cPX9+lm2MOgmvm4rRks3U54VeNU1axiCiT6Y7RYLf
jpOP2S4FuM1mnTiBIb1FMA6dTmyTgCW4mgSguHScDBeTKKsPHtZOwexJKymbliag
SjUe8zhAUEuYf7v9gYPuWT/9NLerWhF0g5mu4204o/+cLiVqX8FULHdxFbWMfXL+
bM1+FsTm7ALSZBgH9s33iCMagEoIB74zd3NK+1cUOLBaSL5Z1BDIcWBo96kf0EKB
cu7XTayP+024mwyTo1So7+v/ckEAMTI/TFduON2GzwqylxuUrZ7xgjBimF5ECTtm
SElqCXXmZRxRtJuhvJap9Clqb787hRez0XNF4imqKZ1BmNWvkUenl4mwMX43yB1V
1lTXj/cr5OSlwCsggjafA2TX5mBvYaSIlQZCydcL3rIYVHtbfeXyAFAcPoQ0SXEf
Y71tQCyPOeGlfYDHZT4R/MxMkJsUMFN9pxBAHvgVdgD/JP/j5aedzWdABK/4uaFq
oZJRIzfuCcOYGJx+Yu8ChGH3ZZap2qWTRx3CmtvjHSlboLa0xA22EI/M9qWopNd4
elZF72J2MEqgoTym2t8yyn5GAENAn8X+hLCytWEOA3/DzVpshRauyEz1ee5j1CIe
o/1p63r7kyFmnoGs8FBed+SghcERKqcNbdZ2vNkza6OIyq7I08Xabcj0oP3rZWZU
HgTQ2JobYcupHA1eb1HcuLRbci9+QNReI9/hs3HH8N1CJzTShE0npTH8yQoIl2wc
M7jVG5V1bETM8gU04zLPhLHHoJeFxzLB7hfW7d00TdCe4Hv/JNdgz51+/7zW3MhD
LyQUfaDMFdzr7UFL/DQU6shk6mDdoCb+NSuPTq3j3ASqiG9MEnFqD1Qgm9uqoyY4
KwcOfAXFfQNyP4Vp8crcuEZreZnt2Qmjwfouj7vkbgp2+4ksarqAhkRUmHUykp0R
IAQF1gpCX0PuluD0IC8eyAxh9rtkNi5NxFTZrbDjGKhQIMyJQP5LeDSAzLO1jUFp
vgkBmHYeJX2QAVMs5IENuf9INZVh/6wZLhHwzZdBBMWntL6q2y++m1TyCJhTYfUh
ZqWZ634EZ99bHog0yIacAOR7T1Xndx+Jn9ab/1k5U2hwqy/25h+QoLSuHgNmJemj
Lrb+RggbJ4hIzX5DVUn4AjG93o/mKNWPiN+5Ibnan4FBb7pvvojWQ2U8F1TKA4Wo
6qH3cAIZxfJ0zWIT6RcyuHuumZ4+04y5VN4H3Gx9/eVvoeX4qr7+/vTc87gXw7Gl
/6A7lqry7LOMsfehfFP0+y6XQsqiFUrShTWQY3d2oRngxeei4eLrffVBnl1jexlL
a6gDAA0aimKDXQbE2dgUTNw9PFvkHhec3MJ+cDt5smYk9ULtBdGVt8QAeAwijI6E
Opf6t4pgM3yTXvDS1pUgecvv/0Y/BPnMZvChxJgvHdJHRAW2czXAFaKyWZ8CHJZV
9faBa10y92aiCpJ9AnJCDVCcRmX+2WXir7JItPEgCvAfJS6ybLb779D28CYEnjbd
UTBiYE7Y8e9+HMa/e1AmLhs17gDFDacB5cL6jjGphBgNpFdH2vcgImLIaiHS64NB
oKaPcuh66mFEfIYUq2RFPDgfnnLYJXE4elfTCgKbiDKPdW4ZSHMT7wA0i2oHo39I
L6tHE9qrPXZ8BqwX6ZT2fxfobv95haIxGbk1Se8yaKMVewDNf9tZheV4cgED6se+
v/doEBMuKDwbrE29Uw0kOx1Zd3c4ydvanE0Z4WAvSoVw8H1e9EhSw9/uC5tplcpM
jEgARDVaBkSwkNQvRjk+BjFBCJwezIZpmokJOwXOkEVXgfkCQoKa3BGW3Tla41vJ
0Dl8I24Y1ceTgKz9U08/yhKtlD0/fCshHXyeduqAtZX5YEmZ7+kFxEE2tEfVqnsG
T37v0qxBDFvY3E3KiLgZL9bvVMgRH4BhC+isborjocP1iy3g1aJ1A8rN0rMCmiqj
UG/ENZpTSwjN4Dmb7+uCEGM5WhuARXsguXvDOBiLhCqRv0NHD6stj/FQvxSCSKP7
duk6eenvUiFTlDFPRXAMWbmX0eo5Y0FYMZPZkne+BH6VPfxrUd+VOFFKUMc76e9B
78GQgAzUGIhsACVkZG3QU6JtidG2phYF2SXv45ltvOyWW/iZuR7GhEOzI4OF4RMA
LB/CfpWOQgCEttNndATdPRBOs0e0TZcV6ENTPHzf89251q+/rN/IquklU+lxl7Lr
iy4VfTh7IW47/9ZHkJ7jgUFwRZSjxvbw7BVfL+8GbzVWzJ9xNKQuNoP+VpVBDKJK
Tfy33lvVXI0OsNTf36kX/REBw62J8dUmcPZ1JxaDTT1EO60ki++ofdzccwSBw+W4
8Sm+1qccuNjdRM9KOUZdnwxZ9Qsu+oIAElefr7wLd9a0NWtXmmXlQCNeVITkEVMg
ECSRk4D/o89J0qtDR9LKPrRyhTWm24uV8pApTNnj8prLVPMlkUqSX0qGWGHeagjI
vgJkpux54voaSZXtNNZ+4YsFj5f0Xxh/hFh/E1fGgVaZCrZwxDe0Pl1J4+LZT1A+
MOMmEbns3/mHykYieZQTsh4XGhcjDGzW1QxOdqGMZJdoBaxORqtZ2OlEBJLz+NgS
GMkBnkU37BEs5U640YhBVanyu+oQ7I4NA1ogUkePemmjFSa/aezIRmZG2X0jzlSo
+VNRwleugUPc08dca4Kl+XnMI+omn2UplGU2QO0TgXMt8zY71arEkaofG5BLqL/b
gh61YHRkbMzjodylh31CGTM8Amm2d13U9LpwLAqxTigbkgVM1lib1idO7HcxBqDz
QATLb3ncV01OjYQqbeyYaRBMkLE/k+cZZFhTbUk3J8AY1HHh1kaWh4o01eK3V+PD
h6t19ks603HcDOfcvPVjx/qZUE5t/yVOsaXoIgkkJayIUxCekP6pA8CvawDsa5n1
mTOdMpYXquC2FIaJVGJ4NWfFe9mdecP0ZNUqESrBQairQwk95BNGE+5h5vIrgNMd
J2svXdKEROoE1tzyDqVziGbpH6OuxqnFnWaX3o+PzgJ7iRUQCSj5elnGeXk6aWnq
qiGEMj8l+wrbrHCVV7v28k6wd+TD1AcCDxKrcg80PD2kuokD4PjeQNncdd/JUfS0
G/W2lJY2/g1K6qe3+M25/9IwXd14Qeu6jlKnnc4k6n9z2Kfs/ngP8yaFHup7FYJd
pKG+wRHqUSUVe/pV5jUba7C02YCDK/GHnSLnDKx98dWTADCd/qP5K4SmzpcGpmY9
yhbK8rww8AUdMBPlq/cFuKXeGrd3bJT2bgBVeKrAjmn+K/BR9cUfdCY3CxvKjV02
wfzXS3Jr/PVnjXj4dYz6lASOhkxtwv9es6kh1eI2jYk+VXg+E0C1USbRfgKS1GiB
zbxJf3SPda7oLq33rM4DVnRsHtipXBjr9jNAq/yZ2Hpaq62FML98Ys67hmPjS3TX
Ocvw33SAopHsV+vzFQYzMnKyGCKLaPU0hwU6aHTj02n7c32ewY0izDNcPx5b0t8j
+b8B+9qEiX0bw2EXL/5nPAU/E/HHhMd5AIA1ttB0qA6pQIh+kQdY5jAiMYgc4WN1
y1CQMDNzaRfE8SKUOoEt1drfSPVgcCj9JLPxtLmCzUwlrg8Sd6Fep4dNF7hwoejF
JbQIGk7NDMalCgkl3ymXt7sWgJHJg9DTgwXue0jw61VgUD72XxWZRqhR8wwQi6Nl
L1qFdzCuD76+FI1kyTZAkem0ORHl2zdDklsaA4C00U25J2K6zI9EB0mgLCbg/Tgm
B9wO4/bhG98+ga0WRMpVLMCT81rn6Kgrw/neXbeG+81nSrLKv4QIc5aIiDORae+S
2lw8iXTwQ8vFS8QeiokfhAQgQ38BMbFa88DseiR9wo7/bNP0EKKRBbVvRKJcP5gQ
c0P78YFuwsvxL6+w1OM0MOdld+Fclxx/kOnjhLDElkjdt9++ztyE3IWoaO3zeS4s
gpm6ps8UOEXvkO+3rK+7PVz+zAw1A7bc4Vaa11G8qS8hGfiCzDve7TABOfL1tzBP
UnWDmUAR9SnVkodhiNhOqaexOprORHrmYGH2QexyjiE0jNzx/5XkbPfdqqwdLIl1
Kb6tnLXBHkxlSSiSt9dIRrgLb3UyGT+6fHy1X+oRCP329/ykAyQykocliNgfpUGe
oW77hRIYM3d3nVLGjVvhzr3XvqCyb0jcy22gGe0UZKJJqHM495xqJkc+5dckLqtx
IMD3UDv8hvKFl03uqZ4aNUdkODNst5+qXPeTHhrkgYOA4UM2m6ME+1fqZmS2OGdA
82tvL33ZsjhEAZ6H8u1ZNiqQNUk19IWaB+hL6F23gEdjnebsGbIYcpEhBPYalw6y
LEju2FFi7vij3FrHG03uPix2kaUPGKjlxvxLPpUW9arPviCvJ3ngdXFfw+CMxzlj
0FHsUyMlPgaCbvuOoDOdfNbLUhRZDA0AbqKFCdtjg+k8a31YMfSqi3U2h9r/TH2N
x576b1F0KObkg0InR8OCK3DFMg/WFCds4G+FetrKQqtUgfYqfpweC8wazvepLQem
V9/AgDilReMrVN406EmIB62WgR87/ujfNNZdYNCQ+nhq4l+Z/kyV7+3pW46G5Vok
HNpcKi9fyi7xXRlr4hjorogh8UaU7BkOWSrNjAqyyoM1v2cIQydD1eSK4yvzzjy7
yTK1YI2AYz0cTBnj5hFX/ZTqjr8JxHbX31xBtloKSTH+uBAsSb4lIoU2TEtwnCGW
zvNdFHlruakGhaU2shCsasBcKlCvDg8GBH1SEwt7Zc8y0dQkCDef/9vzo+U6/BwW
fgLmN/t35r1YLU9zy9Nzp3RuA41aG5HVx4np6EAz80VSGeZyTObcZdu6C4fbmUz6
lMUPri2QvIYCbpcO6uXDp0RKtg807KihCjP5Sya0NB0Qau0O1eYhj+IbsDX7+3Ge
xKDWaaiY/gH96pqzI7jJeg1XkNn5+iZnl0QbrJ9HHtlD4dKuhyEjJgXfCRSMmNU6
JN3C8JYULSNqWe5pOoQdttHvBb5ocs6HHz/zb/Z9ufNZFE6Te/7L1DEfZ+zsSdYl
FngOxhjmAqF4hXwyIF0E9rUpGt9qo5dGDvsiTA77cAN2qSSjGVDqYl/S/l+y9N1b
Zq2FWiuIjSynAk4neWobhXD2HgHwjXPNlYSbozm9m3+RSRQY0xFLwrFLtaoZLn+k
AbD6Lnbs9Wh4t+riwbe9SMaHdBkmGXJTkLoFvU8lmWS7UsTEBNb3ygnyVc4iH3dO
+P0AA1UIAqsqs2K7ij2UOlSPWCP+lhgJVDxLV5oLrQlghQdOwooBehBHcwNfN1X/
Tw+tM4fd5ghzNZlfuBhSvTHH2YU4NHO96UHwK2WSjWkZrPG8L5e4cOq3BTa747hv
DN79kyvC7knaAQQj3cdQ6pVx6pC4DkkkCJyoWxSBuoCkBZdjNRb0S9mhAbc8DD2v
CF+vseJLq2//6+Slf2s77BwFqivT2VwJIOhn3Zu+AiyWBzZfEN6IUGc64qO/V15W
BoW9HCE25hLkheB/FfixyVFb9yXJyhsqprnCK9q6k02j07iNrY+HhTzY2KGGnsPu
bu5ZYvHxmd7KFxOANllw4Y0gCfbtSxMStcOzPoTPmtYAsEZuqlS7zV4GtATCHK0M
d7hG6lJFv+kbUd/yfe8B0vhfr+HQsiM0W2fgrWG5q6/cz084WA7iqcy6uX7M52rx
9cCvPAzukw7dg/T3FRpOodeyFx/41+5lWo4TE0Z+fGbMB+Mx7bnKXCfKZ2VGILAh
udDjOn+4fQOMIVt9Npp144/I4kzJbGBZj77IQcHJDbdcSlDaYHTANl+rfIPwBOlk
dqNhTfCZgN62nz12vcGRrh+7/UfIZqjxHavHgENgGOw6NH8Kq7tZM5dZpStyyfLi
D3pmeLhAGmPe++lRCZ6H5W+0ydtwBPuXHE6tI+lkPq+ffplEFrf2Dp4Rts8n9lH2
Glm2My2Zjo2JqKxQtnEpnl4lU91CHIEM8LGo3sEdVc9KIRL8rBntkNtc2+hQImzx
B88hR2QXqAnRVflSOir4Jz8R4G3nE0puwKWYksxOELIvYkk1POBdTFPtNYwA5eM4
Onpz2hJVzUFiTCy7hboBTSrgOHPW2gn688dpXMGJ1wWjU/7prAvqIWsqSYb4EqFl
wbrX72S4ulzJbiYrgE29wCtUwOaKuFHCH9AY29Qn0UNNV7s4BiUuPb8/GxDvtef3
ldLY1rOrXZzAOTor1CvQcvDW/lSdwuJwLzPCkEnmUKO+KMe3VjN4JfA8tgc7d6qe
9poiDsa1bBqIC7N9ycR+PmV4SMBHC7IVoJcirMN/wEN0EeFuE2mhs+UoFDwIy1vp
NPCTMcKxhClYGI8oZxg+rLB3+30Z+vXXEpwPP9byATFM0Q+nm8EoYWuOqt45wN9h
PTT82NESuKdKuihwrhXmqryHhLN9h8u82G3At0oF+fStLl2CUTENsV2MpyLwqb6z
rhYIrROL7k7yfQHeleCrYtiK5dq2RDoGfxRUS75P615OneuKmOsB/7iL998opPLy
LpX2bpus/ftvxQ5w6Q0Y8qcvYionUXD5BIJg7MLQuqENIIFAaQP5NN9Kzlg76XlH
IZBTrqxOETygfS0IvhuH0uhCiawIoG/lkCIRgW0hIq4xM9aSsFcHXNERcF3We1h4
AeAqt462DqW3ZJOvDI2Z2mlm1GexWhl+N1yolQXet6ZLzNxJYBmhEUPP3qlFDWXZ
aOC1KOeunzToEyA40L1vgGsKjHcxmshhgAfb6ZM/rtQKklfnyHNIDEx3Toe3ETup
AgrsYlOHFOCgwgJs4U7hnDk5QZYrWgF4Cgp8r0dmJGVLUVB/9a7pJwJ2Jkde0JRV
P8kfXgkiFA+8pmTgl/ghc0tq9HjQjVw2kGuFz2+DUqwDXMvk1ctt2aU4xKU1NFFR
lXwNGFPB7QpR8qdDffvR0qBeCp44w3+6rRshtHRsUZlQpD/YZ1UqiSYI7U+U7azw
Aejxb80Om5BY13jVmhx7IV0n4+SO4RoUDrLVjl9TSLHX80vPOD+S7/mnc9PHZytj
u5vc3RlwZFaHzgF1ymS+6hlVfV346EX1yC/InIUQ+QGkyRLlI/FsLLCO0Ki3CNZP
YpbcZs0VvuPmcYmMnyS7rJMayVqfFh1u/d8G/v9aVIuu16co0ssxgrwzjguxx0xP
kY8dp0JnDMti+SFjHtul0P+av6twTyKv/Niphq0y9UrmWeU5hp9Eo4GoyuEu4MfT
sK1L0pqigIUy3NK6iEZx7fbkH1vFqOack7nuGMhKWKKYTERMK0Z6tFEoNZwGhP15
oUF+nv40AHdVJxlaVB7Q+lt/yUreue1yoHctSe+Ips7dl7lp+rNUHoB28xcW/0BU
OSmKWMmZptUb/xbH4DBwxVWgUPXsF7dX+MgjpBwksH5eBGb7E6R5JklAjb2RiDnv
7ZWLcRgsmbBI1KrAaXT+5KcFt6K98BtSX/ScqvCO1HLVcbqmQWfouzdCwV/4AUmg
eAIbNnAD9qRoK0WtUF5qZT3o5HDpraMHeknHXVAucJpya3teh8oiwCnZYenwlFU1
VO6PKR7FE73LbAKa4eCg5KtRMQF83ehNYQE/KEMwPRa4PpIb82ZplgyA7w+RcN1Y
R1Q9xaBnd4zuWZW60NbWuFWSsN1BgiYrsOsRebxBLAxE9ANMqHRJfjU5SUEEkX3w
ByLZ/fB6N8ECDuuEvvklvaEgz3xLTNZHYtbvf6xKLPl91iqvrBrz9lF0oN7zEF0U
/x2zk/aH2NzoiPgzGveTzmpomEu1ucm/sSpEW4RthvZ2XgtkskBkJMh11Bej4mY2
RR82E9XK6MxyrY7UUHry8QysFSh3BtDXNn7N8AAiWKJZW4BRNmPKZfqzeGglrKGB
rUHd/4uSyIIZjP5MqP0f9KW3HOAG3Ecwrl/lSD1wRQa6Dc89C1vkzRcna6Ar6Krq
NGx8GVb6Zw94LUjXZiH3M2xAf/zNFrlKG9A7vn83ZTKx29FYSiPbdOh6yMG9EaMW
1DSPrTuYe8256oD7zh7v6zOjQCUaFg7VLPQxo90P8MBErBjcFZrfJj64PfHpOMFi
mgCAWiCOI7gthuuPFviLTKFl5b347g1CcHg9SQUbxhYM5ICmmjQ95/YKlyia5+ew
ABIUzSMqXEgdsY1fOI6rny/xYjux25ITaTbH+Mxj6jAwVPo64QLfHKZiStoApSDF
JKeeuOWNRGsH69phxniXDYTUVpuCjEH3xDrvO3yf8YWxWWMz1VIcKkskKQ/wxcp0
g27vNqDzwIRfT/cG37WfcI1UjLZjz1GRcbpB4sx+8Nhae8Fkn2NYMiwl+mVE5XdS
cGguPTgaOuUx4HkzTRhXBNmu7k9J4wxAAQSe+dfvPhRQolZJc6XEkFHq13EX/quj
i9xcUMpkm6+D1d6lgfX61qnQ12BffJxv8BqywLUZYtokyMa1ySzdDPzKJHNHanov
8UQH3xdAI+icsSt5wSuxSmIRQ1qAtsC4PwVdN4fOsIlWlL5Bi5v36hAsv40bpMU1
/y6dWhUo9FsJisihMRN0iCUPG7HhRzQxi6V9gEaWQuyO1yJ4xIsCNlBz6dDCR2ZP
H4vrqlSFkz9874eB8QVAEZPnqj5Va36cI82GVqSQyURPhMMd3TbBDYxoF1oJS5hW
0+7k6CcLTe1qSavYtAY93qBglJJaNQd7Vj2g19wcto71aTGWwgXLyRT7z7b55UTO
lPp5GCrjzd76rBUypIYx6dJkFQ8O7aYIxZbqvJKiipS73DnRIhvf7aO3oh+jet/K
RmClOrZyfaabTJkPJuVYmxuzmZwCS48Lu5uczySMPtJBOh/rePBwoSpapmmp/9mn
dk1FLTNaVDUSvC+RUbNQ18hoNgliMnKy6+uIOrTC8lOjooxMHgdm4qMm7oq53mti
FUbq08pT5k7enX7jUjuGYCJ3ev6goosKaCNBSS+4MIRbTVh1fH8Jqtoaeo3JoEcb
Q7+MU1v2H2rS2oU6+xRqFKwBtydInZdJAaQDtdrfo0GsY9fDtl7iQdYGTPtzsP4r
fsgHfNqay5mwKPwntEU4E71/YR51INyy6euUmhGbeJTzwy1slhdJKcNnzwwYoyW/
7Fc2inHUw0E+gG2l3xSeLyx6j1fzniE94gum1Niyh5lGmwCjwZv0YMlgfnKjPXQQ
ltnb6CPCeNmdJ9DBGEoz6p+aojBGM6V5n8uHl5Wm/JC6LWhFCMu6FnE4ZioXjFjS
zHFSQCUmkhW8nrFoXXSFf6R8sRJx7j4RjnbFfStPY1IilGK3H5wsHhOGb5A7iijr
51dFxKS0f+xSpcSKUhexmCAplHbxZBT6k9DbOfAfxOgJAej6ByC/iinNcK56C1aY
s/DqD4Uux+EMQEuRQiuHfY5K1Ztb4vuIV0ZztPcsRG/AGoffBh0i8yHYXLf47qRc
SSSB3W0L4+dQ94Aat7lYpGsLQOnLsyGf/DuDVusAwZLq6MbjZ6Dp15+CyJ19259e
62T/6LMunRMOok0sL5T67Hp0Gsp3jp6Ba0Sbn1tkvENK2avS5M7YCcIiVx/mzTx5
q2cSwSO6Yh5A7Nk12XCD5kk2NKhB8jjB4pOabgmfvNScQrpYzqYo76PdpTEIGEjq
dLRo7/365D0GTr7P09kvzBIspTfwzfCDUMvtQPlmWBwoj2yj6n/rHVFzyGxd++FL
5isqQpv+/HW9CeHXP/VzHLFqcmnxL0940sj79Cut/aMLFMQwY/ttCUy6fOSyQGng
dosc/F/OqtOmMW0RamVXabmSJ7V8ii2YaX7iWFj8BxUXuHRGpMy2VMzNak7sv5p1
bh0Egpm95YumguS9byTDs3ifzU7heol3sRu/wlMU83WbtM5N9/Ywyq/k0DPc52Xu
hI/NbsahBd+P8FzvdO44SmF9Q1fzt2S6gK09+cwbHJuArMzkjibF+vRwDnQVlTZr
TpzCiJrbheFiQGzYZDoGkLyt/SrmAahNJkSUDqM5KJ6OvRqVKkHDj/WvzfDygvkt
4qPjbpWsruwEYJVnU2pUUMWF6Z3qmzRWWAsmtXvtPo7eWXNiaGz2w/Db0reN9QrS
3Adxm2QUYu9Dwv66kHuY6M0ReTX9jJKGs/znEShrQNYk7mWwDj7nJyMw8lbrDNOy
LtAfc9cCopKfTS5nwRVJGmQ/HaNfoKRHZ3WAPESgUdHXd6XzWr0Adf18rJAtqrhY
fjo4gem1F9b1aD78uwTXFHtDD5AhC/3BKXtbPbrKWzzkSFNLgfTglFPNpSEMB8k0
yU/q1d3cRDVde7GkJQ7dqRRGoa3lCR4rvF8k7wdovDVNN4V4s5orqGDRFL+IZmBH
hepwHxPBOrA0ke8hf6+kxd82DSkB6gd8W4mBhagP0i8fcqrdoz9oMrmgjXX3bW2R
RtNdcpsT3XmGRMaSDHHt1FO+GzK0y7hG+Og6kfvpGP0YQCmbwvB3iSvAkczaxZo1
NYi2Uktz8ZDqYwO3b5WunAWUI8Js0U7R5sK2JGN7qFF6C9dDZIrzBJRwXBlOlcP9
c+AuCQ3OzdBXkXY+Mmdkbv2xhvbJmAig8fWX+MWD3ES9+PC7CX8IUkxf9SCRlCoz
ZxkQacGPzwrYM74uxV7Bojbf67EEzrPPLDcG+kRhRZ/5YVFLkp0s6uK5GhxfiLag
Vx1xBMTI2bE9zCmecp7zVdgcX6C4/+z5JkN6Ch+y+GkBQ+gbLMNX/10wL92xALWa
BBHsh6YQElvmHvx/bzkxtcq/t6vLt0EiDl0xXYrUV8sLRAF3Fgjv3LNrc2NXILSl
9qg/Eqc0MYspPc7Hs5K7cBOF5Kq3jDAuj+MxyirtHAWzjAULIZzJ6cjFwOK0X/YD
SXYeufgxnuK0gv3iKTuaWhXsXzXqo0/cPx6TQ3UTI/0tM2JsPNcHI54YjkhmWA55
z2SfFD71qQoklyr7pxLHSkEk2Qr04iRE5q05Ml6nnno6jB/FlK55F+aAoPBiOTBC
6eRuVrHvKaRcduLmT86QhckNcFh48nNAX9NLyVc8tJgA5tZvB1zliKA/HTNJMz+j
zFRUIxDzwwyjYHT40zsslDkeu7JogZTmCkmm0D/FEP6eRs3Td7GgDFCsWEnM7LWG
OYOwOlQnTr31BYWqGxPePhB5HceWbWeM0W6KT8Fh0h7Wi4D8Mfy6b04E3KZWFlNv
BZmd5brOR83mZ1zcJt+oazigXKoLgMgo3KKQRrcZtQ13fsU5YJqhJXNjJrxee9IE
1hz8ExlfhcrKXp+kFR6KyDC0mXQiBAw34mZgL4NdD/bFqJu7YQ1wlhLp8xGOIuBk
9k9PgWGX6KYyjPkozLIkBxEMJMonZhkOmTcS2ixeUhvvf2mXKAhj3h0m4EcB0L3Q
cl+aZS0QoHn8WwfpqbIyQPIzlJ042yW/OmPi3A3/GLHWnOVdp2go9KI77ROHAReD
3t0hDuJ4DMXYiCQ/oL3p2iJS7KtuH1jPBcJl+Cr5x9INTO8Zg1IExKm7UJV5uC+f
00qhAGaJ3AgWWpS31ybIyDNbd1Wt4klVCfJa8e5yjq23LP3Zxbdl0gMRz/33+H1Q
Z0DYrjEyrk/OMqApgl2OTaHspae4U7LTsO2ppR9UwD39yobmvek9IerwvsG87YEN
U9g/wIBNv4tgPdrvT5u0yERx5fi9LDRVMnngIS5JS0WGp67kBJ8bbmn1qw3EQcGq
rxk8lCApuwtjJpr/YMYgbYpMnj9tQ7dnHuKSgPmyYd9Mr5FvrShMxEXPCSCu8n5v
Sn1lW7ZkimlcSNKM7675CvVCSbZlAvgr5Tj9OfbgPwXiHJ8Ng7kSdc2OuG61emHz
lJDyJoQECWbANnbgR0WNfHhkUTYPz6/IQ6/+P5K8id2hRrWMqmIhA0BIG2OPtxMw
j0+nf4Ba/Supog5T+WxGTbxPXaeIIyuVOHFGnxTtDOQyhLKicM9w+szzID7u/6LC
hK60ln0fLb37Jc8URUhbs4FlEShIwvKdms7YDBAd6jVVVUfQhvxWBbRk/2Z+guCf
ArTBU3/wR2p1+mZ83T3U/U6F5ItOmKgotpul1LISTa1oeOcoAUWX3XC/e19UXXuc
grRXqDjeKBjoVruJJDQYqcJ8n70SQxrMzXAR453BF1qpq00vOrewlCu8LpQhPWUk
8OZZZPjNp+bHGHM2F9DhY92tK27yvwRtI9Vv5sf93nQKll0xN5Kd5r89y/XFWb+K
celRJN/cotjxYk8ulhkaZ6pVrJKSbdnCT5uZuhwcTY1IUTp7JTVVj2mASyNftK6x
QWEYo8deHBaHKC68JycoQkH5aYRAtcNVb6qXvrdXHeM70s4TSpHLTnpQK1Q3Xjnx
klqS18HRHTBwvOcZ7YiINykRrvUhh0bT3t+rkqhVHp8NMcc1Okqp5Vv0u5JqDLuE
oSGNpCQOjKTvylmC6oa6NUzZNr4O8NKXhHOh3p5LoEwu8Ej8T75m4QQAw/T8p0HZ
+4vv4zSFRZFWLJ1gRFgrGap3sa1rxZkhTKDGJ9wAtgXMmUZLANlQRxTH6mpzBZLQ
OGH7ajKg+Hbgi7vYFfnuk9lzeVm7oYMJupTWaWOWz7lKjEHsFPYGR1DdnMgA8iKe
hC5QzipE0nvio540oonWXhnCiSw5y9+KBWTo4F5XqnjbNE6pHOYZV3O6fV0vh9jf
iwzb1r8s7k0+HuEFZkYA6aXDwqIZpuCAq0uHbrZvPL+YleYsgJuYeU1nraf6Oqa1
lJVBjcq6MYP0zrDZUIlZsVJLrR9fwTpiMCcyWuwE+qDLlySudATjTg6ZXmxb61CE
LK9a/TFN6w2v+EogwdZrSNaO7sGs3RubfqGu6o42sHngDi/8aAdyYO1MDWa3VL1d
BTeX1OcDTLa3RdJZTPch1m3BQrYVepylMvXzpxEsYqIQN1mBYxay4SXNwViO/TbO
ofWHhoex8x1UqPWRF3QK2XvstQhONrSUXwhLYnBmYEE2Gz8SttwwuvbojSg1WTwO
GjaUVnwb2CXh1jI87Jkxa/otlppC9hPxcX6T8Uhu9xBVE90bG/ArccppmiIK+vC2
9geMmSgiTXGrbY1tcEFyBkKVRU3qC6wA+lSFPY+6a79NpXhmKgcEJT2wV/Q3sxQ4
/S2Dx5T9CjB/IevI8w20+A7AUPv19q+eaY+KoBOe8kdP+LrTa0ThegAyi/HfZWgL
epqBi9b8Bjm99WIF3E2L/V8HUHJNcTHsj++9ya4C9CcSLmz+e4Wx7DxPq1EAovCB
EU3znN8oWodiiIiNxmGvoXMMe+oo5VTrR8ewdPicKyJnT1IRLHD2zF+Lq+jsvjYB
JB8LuJCIM3nv7bdj/3RgQfXL/SiumdbIEYcSJcJ1Um/yxmBpni1QnHzUgo30gmer
lif3n1fdY21YtKCKZNjgJBxABYRGGDiUGfbDE1Sz2GPqS75V/FUqAITPa7ZT+8gr
+djZnLu4Kobm5UTprX7saH5STceo4bWX8c4TjTdeLF8VMhsEYH5/nTN/0/Vj/Gtp
MPJopyBwsCMez7HKyLDcFhDZUbkBrkReZe7NqzCgDQDOEdYjlHBmYMN+nSwtrs0A
bwXLVW7OZRF4Cohjat1jLU/qn05KHCCIAbc+sYK3YaDrrvpW2TG/gbCcQolPs/yq
XM5olSemoPwj20Mm8olN6X0Dck8olLlcKnpPlVjHADozTZazW/kfiKAIEc38QofY
l7XAIvPlLO5QkwEpSJW6LM7k7zf7DOvvN64g1KfyAKukzRwzlAbyklEwUwSerqkC
T2J3XuGfjvE0gMZw/NRPZorzAqZfbYkGdBL4a/q2K2ahmonshqEMIVamPxPUfXA2
ShbE2jnOhC2lxWjco64dMTmlifgLqJ3LPbcLJb8GqITyglARL7wanCvViUs9FaHa
KmRhiWBSq1Iu8Oci19sDeS1tKj9r+0RuIN01C+ZMTDQBne7Nka9HKNMtUTg3ORpr
Ob9jHRjP/5SUdZU5vEYowhBD3/naSM/Pa2nogdBRvMr0nwVul/kq575O4ri2YfmY
u5y0VKoG9//KAPoqGTmExyFq3e5fg8K+gXmsrEsz9C5hHN4l+4URJtDI3gSQGFE6
rw5dsFMBrR0ebgF660KRdNjkv06yq8ccWQg2uMZYQcmk7b6TTOVvOKhv1Es83fsy
e8JmaNeKv8lVPUbhW1rUwbdf9z8+IRFZshrurL6F5BhiJfq8sNBCqChBVN+1oIOL
cNKz0GawDzjoLhT3/OcvFwMH/591m/UpmKnYVHP76mr88PMtmZSdN8QvMYis0GYI
cizkvgEho0NAhu5nBJbz580rcNEYG3VbbPzT5hSzeCkUaHBApe67YEzNKyguziUI
VE+9Mz+4jvOaUjYAw349tgdxspiN+Ym2HLh0e4H824T8mRfOZL92xTjg/mDBGwEN
wTpAXZY8PYuiXFiR/tQMNLriymyZ9PAQLeyXLVz83IkOCzMrvqTMCz2WiKxOLLC+
F5pXhZpKMAtcnHVZDVP0aFMBYUW9VfvmDTgjvsKB+WHtiwHhAC2PH7q1ZkCr1ftT
b5kF1MwSObc3aT+TPhfqBGrM62OITRArr3QIjY56eLffFQ5pwrfT0/eDsxEGIzsY
gBUaR10qmPBH09jaHXfjBvjb6jbsjg0HCEzpQeDMZC8jUpvEHWVULRsqCRcApVWc
LHDBWkbzhutMFO/dFlDF6BNVs2bB+1ujt+83Tq9PkyrUh7EI+AYFpPA6PYV/Phos
Rc5ndkiDTc4n3zRqroEqWMOuOVGUHDc75jpQRbUlxAgt9s9XBjXPSWM4I9+BSC2N
Z/+SVTFmdimOHBLGEeTpxB+udrCg1gDPo5TDgodRMCz2zj8Mku1+MUGW4+PloLXP
9UuW197/st9Vb0iLJJ9rD8CnBAWqQcNT0PUcF0G5cAmLG6o94tBpJOWnQC3oHPL1
kXabZIxKGPZMlgpFptTJphwA8PFG7vFiFM9fFsiXi+0MxfwiqvtoYRDKVA+7KI46
ePlaDN99qxbdZ1RXqCTgz3wl232BjLuO+1DEaRFsfXVRxzlqWTXAY/IiRcBWviwX
CvNPksWi5C+8eTa8aNs8Eoon3SfQmBLcDkaRrcYhKWpm2aT11blgEiH6I6v7VqHi
UMugnhCxEHh4OzTDQRjN0FZPCKGGGrXNh+lbJkMMzqaieO9mY8xFETy0boRERvRy
3ZA3NzZaHGbWd7/BT+8Tl86oymVV0CXp3pRFzhXxiT3RAkbxipBNUje3Z8g5G4UR
gZbKvfNd3czFWiq7i3aODesc39Q2SJ16Jbca+y8o50kRgnBLhWcpn5GgKmynk0sM
32bBce3wUoD2VKZqVY6S+YtHHLylJW4vfTuGnUK1vwirjEJM/N/yNiVoTGg595ya
RZ6JHJ2cboJYZo8UEGmwEM0BvgYrGTxtrGompbUy+l2h1437XshbuIRwUDG8r0oW
EjnE3CLgIQwLuP37NFvSHuerRxJN3BSrcTSSRWlkOj879jItxIqAp5jtX+JDaAbi
RiaAYeTf23/lSE5BS2lBzVX2toCDpLJz1ZMJC/VN4r2vpq5BidoWb3iTdOuoa3Yu
9v4AFTeDJieKhKKzmdmD+keWIv+UuUvB9+2Yj7pjReXd91i6KUr1cKWIJb/Qg5LP
k5rLSvaremSk3t9tYZIWs441Qty9ARG+uckoHMfWKsmsG6C6jbRbXymrYQMomxhA
a6s673+V7uSSSNNe0mJZO1/8jDJCSq9wZ8jJ/YEOfSSjJaBJH0XLEUpguwkJpCK2
AUXc9eVyhdEVYwOvOw9CbOfp+uCzytl0H0eBBedORGKszaWWlk6j2MuXmPVeCG8h
B3ea3n4K/22UnkIbd1E+BZZqZpT2BFA1atQgnYeHQWlZW15/GoLavmjPkco/ncHx
PkuW9uxJhfpj+77CRKe6DQU/qWUtXZlFFn+XftXnaQozeA20RTC9Ob1w7dIZSh3u
NJB0vwIjEoYdnWWSxnjMrdMpEF+fr5NF7siCS6KVxokSh3KfLip5ZoJAEiRabRkB
1kV7nJTlTgBfD3ebnlbTEdI7x5TIMWLpsRwohLmrg9RO4U38CCgeSGGDJ9ep+Lat
QRWfwzRGwmL2l0hY7ZXY1/3BQLqchaGPPi0XLCUtf1VUFqaaBJyic3ioO1IcOAox
QvED8T9Ca7NKMzRhDTBUSGYKiLvIRoUNYn1zsgu8Y7F7HqlvLEHV8kMv9oD0r9/2
O5dR3xSXpbCIeZQR02KwETYZ98sIKkHFNDoLPmp0gfX68CiFiACiUgbocTqb9Ou/
Wtd/9YMooVB5EV1+oAQrpqA01B4xd0WTTcaVCt3bZd1G+KpEU7p09dMe9TEyhafB
khxHDi672oQXg/r3JrDmxMgAvpaL+h+ixep8jmw02ULf6OzLbKpJ3VoTMdAR2Xbd
sjtUTJi2VudnlgLR14Lx+fnv/xCBZv6/NPQiaQBL0oyfT7XmsvhrcJzpr4ZRXvlZ
wtGHjKi9mMEtffMBJtr3/qdl0G17ferGhEaNXy9le+qrCyTG4TsPCZa8fNsPcQu3
bO1OFl+HzsiDHrYFyU5gJNmOstFqCFaNkQ9mzD5X+Nc/tmnipTZysaShdaVxYfad
iIvgNY3a+Mn5wingDx3VYNTxVQOGAwevu5trFTk2rYjU/TD/vTzSBfRRaNGIEcyU
Q42PBL2daYYr/nt+0eKkzVeGcC6CghopwXjPCjuxaDLWyrgJvXUAs8ZXXIArxCAG
kX5Ut58a26M20A1ujK8P0OwNoRJeUpmF+63XeWjSL0ywX3GYYQFeI2tNBAuMfzYD
IbgVt9o+IUYRbTwSFzjSidbVRLv3pOpP6m1vTfO4N7APw306wknWzYBWm2nYUH6W
hN/mU/gERSM0UI2Hl083wRqGYMrmwebIgUC5zmiEEtKz2PFtaEGXgQHeipXWPEQW
0yqBS9OFMf7G6mZa0TdFUJ9eEFRPE4Qdq9PYQIuKezj0Bpf+AspBokSkxqmqgMCe
GQK4aKzdMTLXRT5ghMJLfvGspPfgQSWWQAjt8JjzJZ+7kCcxpW8sB9qEgI0ilN3F
/PbyTJcIXj33hQeEBUECeWOhbzxWzh6Uw95fCZhMZKLJXPmMhx+LrZ8uTIOQTXZ7
in52w4bQrbdU8zNZxv+jPIynxTr9hhUKpYdlZwbSKarSUEORGVSt2B5CTKBl7esy
4PO4wQOXa3J6lyjoSFKf4v0lLHsdJcxcsIZPW5qYA36BI3w8kbzp4iBupwNwC6n/
d1OkLOCTNC6lKtzD2lVo63Bg+TFutXwpXP6NPDhWOY0baThP41y4O2ABKh4K8hmC
Tj8ZAc1xGTp6t5Jklgj5Bo0fLFg0yzFdXLAlwYwzirvmZVl0WgApLHujsH2MJeRB
7dNX1m1bMzxsWR7C97IfFUNF3s8HHD/3OjD1Dx5HyvGcho7KfT3IyqX5bqe4BFSn
KkdBfRuowUzk37YNWL9aVLSBChdkcR1j9dvXJv9tokIx5L4VuMZ85IQPsOMx53kM
4HpOUR9kO4VH8rlUFHMBnsfedSpfKi1CWTsxtgBruB7oKFciB663Jyw6wJ/wPKGA
/5yJuhmV9Gp57+2RjruUk+tDWW9HfzbQFLYLXzAgkC+utBODfCjB3M7d5y0XByVP
tB/pWW0wkNrpAAmZVBo3QFTrOCdmfnkNUYqNB/M5np42IPatdFwO+eaLrlmpVo5U
ZZ/pM2XFpIurdTgxnSHTDx/CE25OjQiVns+99fnPIiNgmeCBfS0kFRf6Dkm2aolt
3tkxRG9j/D/UTqoZKkdCRanEPyLhZ5ufz6t280t2drUeNvoJDZXz7wD6CIb7fZll
5ZHbSB9zgRBN81ydWvXBguITGIoRGY8q4M5aMrU9zDQRNIEZVHcgJSWVixWojSu2
swjBuupjkkDc1iwowxJZ86qgJUsM6RAFuvwh2hDYEpkM7oF8dgMBBxbtnVE9EW7K
9aAonX+FGGkwxjf/47wVn5y/U/VWf0zPpRLY8EE2Zd4iqNmpqPYXZ7blJ6rD8gPY
qgC0HvRSLj3cesDLveUk44vJvzp6MQPL1zwcA22Ees2/rBe9C+/uRfQU90eW5v7q
sPjVS4ph1hbgyqpNTpLO8TORIPaJaGdUW/m38bbSJf6RW+0sGwwAr7OF1GylokcS
xReSXlEEfcPKhVqzcnTmmY4+eSwKnEkR8R2fR3g5PyNLcWLwUfaaQ3vlJJWW7WAn
TGkEaPGt+mAegjsRtQV5GgD0gJNW7zd5EEWPmohTZddugj8SmhNm33Zc/I4oxd/r
GsLlk35d/qD3gr2BqJQm4XZX3rgYGycTZw9t79xKZfKTGxDMVsWHwBxXZp7hWM3R
Vt2Yz0IxEIdRsv50FsdoItvVT16CctQ8+VLpa20hqSxXwKfyMX4NpmJ/BQjepLFR
l5PUAJC5OhX0MKkcnMv7cRq7sShrVtMYne6J25SvMye/bozmFmbn6qJIrJ209G1i
FvXME4shud/vZqDYD/bF4NesSSmaUzVigEbZXsRmQl1rpR+ZW8HSUwTerKOfb5LL
4yjdQsgPsW2Z6lsjj68T2He2Rrxe6dXa8FEtjaEYRh+igZyLxAS4+MhwHFnrIphL
nQrHpBh1sYSIhlkZQ5VgX8gy/1cOyyBHpFiTLXcF08Lqz7EtewHWSt2++dZhVdVV
tIxDLvL6Jt8orzo8iaMW7Si6Gv5LqBbrjOdBThPeFV566TiaV9U9mC9+0ExKOkbb
NHEQp4c8Vm6kuJrzwZ+abrEPYiNx6n/JgoWboA8aIf1Av6EEHoABpEM1CXSckzup
zZ8qaeKx4FUCXARpYrLJd4gbLvFr9v8FSEZFw2qrRu0Laf4aAJgCwnsoGtqzGofE
edMhJcDuMWSYP2B8nJpzg1LR+HqOAVlyJ2iIKSDrqd7SLELhXdSxWMMLzgLzrQKS
pSUtXtMfUryFTmCEBMKEpFRy92Iuixr9HajTXr2R8J7MvCBjyCR/gjiuSaDiTnzP
R+KLyJh/2oGEmdNSeQrYEATvXKGXhdx/AJn5iXYSdZ1uzdVMCrqqK99Ch99eb8i/
p9lywV1qG23+su/d1feaqKc5FBllDYSlOyzw3Yxo4ulcXG2IgYFcVwJbawHgESub
qemPeMNUQ4ants1o+Mw/yX0ya2ePULEUeE4wmKhI4gplRQ7QkgOvrMV7lipoJvSp
MVCinG2ufAdum5r3tHH72s5s3KTvxM4riIVmmbVvZTz8fdzvic8WiGVtn+FG4ajf
RX+4y/bvKJ85wTtAGmTCH2hKz8Ix1TxuWG92hOhoDT197xlfCWj5zuWLeIj8XrdI
2DhrLedim+LqorXtNCANvMRaTM1sBULidoJHPl9TmrM4wrkNEdznJKkewTZma64I
C0XGp6qoO0/MWV0Q9CHhNZ+dm8rzKZ5SBWG8fKXOxnteMfWfxntH3gPXL961siE5
tekD6zKiXxPYBDgTKChAS6ZM4PuCs6UOtS5fLEPu11VptM5dJh5hOB9ad40Qr/3q
3Ft6oXznit46ZXw05YTcVBkPyy+yBSPbKY6DapVGLo4XnPAtF6jrk9irRqWJQkQy
G4EGwJZN2Iz8ITtyMon1hA/KnM1uOCLNSQJRS/Qd1YLAh2i8LekINwNpNEz9tdws
EFmwVH4opFE7qI5tnM4CHl60b7OZv3VQBhX+8TvZ1LZ6zTjzZDdRL7rFdtonSMil
8NGcyWvEsa3LLFf+Bc4w3FW/gOvuvb5MgFtwwDQ3MJigXHgCgC/Pw3P50lu9ejfb
1ejrVQ7L40SDJceWgUcA/qJp3D8Ah8B0XZaD8nmz+2fYSmkckwrBus/OAnweZeVI
oV3M6gnZxSKIRXWvEMF0p57auD+7M31DFSA5M1HP3X1c4dTxyxleer+EDy9Bxiek
vJDf2s2UaRZRShZvI/yVmwBRfMT7b6Xh2TxFYVfogb536vY0v5qWSgdDT87yNguK
1G/gMeViD8tLtTxIneBQ8eGLQ3T62BkT/6EjlHRMubfBrhD8uYfBR6sxjkh9Pbjk
z43Fgf+ENpTGzkZijlnqTuhPe/UE1K3C3y4yBBr8g0ALIGIwhrD/PK1nH/5Mvzqj
/ZoJkr9UNIKjQCzHy82eYOfu5msIpf8NY7VUTQ0ngwXY68j76wnW5KT0a9xpZQyz
zIRWN+j3Woh4NIlckXhOrnitgO+fdPetCG7F5754Y7AYiwo8nB2Ybfv2EtM09VA4
vqbvClHOP9AbrmhEIb81KGfoElCXK5+hBD5P6Hiu/znkHOqOJlQHd0pfasAH5K3H
laB47jJAePQxJDeTTUqZyz3VojvX5Kw/rAYCMoDan98M/b6cuhPlYkaq6Fx0/38A
oR22qBHIKTWMJsV+lpDcrqdZzVCA/6RtwW+0O7WveLm2hnOxJOPo91bK7wr1tY2e
ULrLgXn5vYzvuwV/XH16CievT46C5YsoT23CW6X7aG//buwD5iwF964ooxx9pwQc
GzO6W4x2otxpcolUAi7T3B/IIqP+oGgrQtpgBol1CZNp4hmiiqTa1V+gqQ60RYfi
ZZBb9lcsRo9GvAaBCvzV/FEe9DpHJart16GTTRwLPfNKv1JpuQHhAYmOHpsvPOBB
O0jDnFKv82ThPH4ufr/vkS8V8PI3GTanPq1P/l3oto9EtxGLOW9U/wIezXxpSyDS
sHwy5CSvEip34SIufNBiO+VaLmlDXJsMEgjS8eAJlJuSwQH3s4+OZCjQ7g8KQe/c
61jXehGXR6DJWpbKsrACSBjVsstWf1M+VWFpeSkXEAcINcb6kbBb/QJ4jbeUee11
A1ej30tdSrCDwCEuml2Iv6/yI2aAPsAD5bN64Lz+Zf5y9RBexDt/5vK8irS0UsfS
8nYRTlI8fY96Zpvb8Sg8Ijxz/7VmmEQYjh+6KMbUNjpes+kCVUznLbiZdcnRBF9x
+zxFVZRH7pIEtsb+BhhhMCI+smIb2N1jGEGPX/ahrOQv8OsyYD0eQeA5f4cYSp2o
+03iQIlYavy8hyqYFTEi6yS0QOHyIZZT2uNROLvbeCBOPsSzWQCCQSbjkh2xgHyH
PucZQGBLOqp6pb2YzM3uIxDDN/QC62XXnjNMBsTU5Eia8YEGMWbtFwxiZdELAZ8U
5qC4GezT+IJ1l9v1Oc101zAXeZi79a0G2Z44czdYG1CK/d32aqnJwpTLALuWikEV
pqFweuO51Mtri7F8Lx6M8vmomXSR7AmT8H/SsZ77hTJTihcuX7DeN9nIzREcSDAN
7rQZNTnqIv54j+p0sMXvMQLlvIETUL0xwyheltQiHcfsQpqieNBYV2gRIzd72WO0
gOgx1TVa5O3CnOkp7T/W5TTfbksaLwTKmU3GkVR06fCBf+nwsSEXhvdOjvtOOAkO
Hw4sLS8x8SwVdDTij1xzgdvOrQSAht5tOxLf1P3rP2wDFwvszxCDJFzyXM3EDu2Z
XAtOEecTn3/dlfO3QoJTHvMa741N00WHJ4VE4s1zVOtL8IXUX2BnsBpFHZ8QICuq
bD05D+PeldR5nKgAEiPqqApWfAOxVvDkXSBUYHwM8jsYp3PVWeKP0c7iT3Ps/xGH
yOWSj20/XfKQAw0LV+7JAtLfZ27rBbxEK7sUBq2EJ0BroKhOFIbMQsSGoc8974on
Cqa4JQOoY+GZBorautazERbaYbT5zyGgURGjXHD+yiaGB31tWI/l9bNclnO2zzgq
8ZpclPDNhhooCzjQP0fRygnlkHHhyaMcTyigYa0ZjhwdCQeYygUKnNtFHY9+JiNf
HRUQlEa8yh7GwZV0zo8DYsbzw9jY6NO6rm3IssEowsQmPDuLizHjvV1TtDqhllGt
lMye7GOijyWJpvewp0ewHJwvl+ICbvgF3zW58XfG0XhpY46CcqSpmLNlHhrnEE6/
j7/oNmo4/JVcmx1js1gPsJ950HyMLz9+tieXFclvNtMBE+8U1hM+z9rlw3usU2aT
3oUBiwxvj2dApHN4r7q/7tB4AxBEuS6kijj/wAqKeL9CfB6MFng4FTCGTReQNh8R
jkAIrmQHixixcS01kxIjQStLCK/FrOrN1I/aXbY9KBgWb1CGwLtL3jOjiAm8JY2Z
n5Fz04OO6gUXIcAF0yUSeo5Ss25U7bqEn/PxlraM0TZ0rpbk8BwLqINqg7oprDVx
uyJxLBI9i9Jcee67/V0oJvMlmHsj7EWYX35rEkVtjHeHvHmkF9zTlmuGbF6t1ht/
WD+AoA9h24Mil+m1QaxVWRbRVH+acIsLnNO/V6uK8JgrRebXg4uJRjlxIQzXx6jZ
cBFpGnGOa/slwkla+JRS1qTSnkbxDzWguusj58OV8PZLfw+C5ZXPCXqOFCXBOdRG
sXWfqhXcya5kX10oH4Z6ZsluXHdI9/OH1qWdis+g4JsmFRoaJu6vwq+03eNYpoqC
k9lfzVbugNKCkeakRxCuH8rzrnBZOGVJMjhbSP4H8dpIJGibdl53q6eyFfUHxpci
roR9tA9crZQrP1QIVRB0gZL8cgRDt0FmT1v8PrvZ+k9sg48baaDGENE2/oHNRD0B
PZ2zVrFfCJtetGWq/bk8u9OeHDz+E12ytMAXvTseYkMuaFeUM5SHd3ogT5KHc/BQ
SblLN19cGfUJbesgeIwaCqNJTuyxHUNpGhNyD8D+BZMBuzPLDOwEgFeMenxMDDN7
xpbauhKsaPIXefYo8qG1cbjAoP7VEVNnoSHlAbtDRO3J+wdpOHDKFn4S7vYnMQJi
iGQTE5vWgj8PhybJ4gbG/tCeV4ituMo8MBwk8kfRDQAXmJhYGYs6rek05HdY1oH2
XpPQC0QRpJXgTuJHyGx7arYmzdmvE3uV6azcwZOdX1DGD1W0GvQGrPNeKPXlRjwD
9Z/iHJXh9H0KvYLbIDqrdhlQmATQ6GkQipOw9IjtrQmXw1sirGtM04EAs3znrMj0
rB2nVUE5Yvlgg1rY6tc37uU40DsFyYl64uDnlCNN6Zo0ZJNNE5rlGkWxN0pZjyOR
todAtgkblO0BQBmOY10CF8k4f4DFNGkYjbhQHEp4j/ACPJOfkeswfEVS8/ajg6sY
chB45tZ9zgRxZbDNL+lbPS/qidMDdtx7jsCoptxxoCqzFTC2ih7dMT0yg8w5fJE0
p2GpYs+0EdpA+HxM8y8HrSUSCbkKKd3GY7LM+GYht2l9RC4zlPgg018MYNa2h+yT
yMV7jNjKPFBoRSk03lSrTw4PvGUSJ5jWlTtIlxaMjpN/idEvyk0ezAFcWZFD4+xa
t6AZcOsS1VmPj3gq5GgL+vs2b+WZOAuJ6H2RRZXnuL182CQQH9eBkNG3yV4bbOvm
V/qCwmP50xy61QHf6zZTUNV2yzvmx3YiLsGyfLK47OmWPNo2kZbr6n9yg+aKR5TJ
PsXdqj581aCLB66dz2cBXJPgEDNY00b6J6TIrVPHziS8fKPfLWogr8+EZknSNZKB
sjHSbNCiXPWC3G+908ACeUpa9pqX8NNYD4I4D9vIqSBgd6hK+52/TgQ0uC8rekzw
hbWScHztWOe9U6mymNN5+xJJb8L+28ReCx7GKXLh+0gs70d4e0y+RxQwBAYd4vbv
71RapFERhINHIn7G3nUJETnUcuIoZL8IRLU9ikso+gwbvgbw8qEpJJvhTHAiAjje
f0Wwxpg9+Ug2FBMOY7gEEaWwtybrQmbYlh3OVoS5gRi5DjMqPU89N9QAkTBMw4Gj
lzUqHWsaDkFIUD/cWKWmoTB0ep3vcv6ulmfWSxjVw3nZj/NxH96J2J3WaNePZnaB
MujT5nSGQhQ8PwImWexYv2+dzSbEA8+qx42aXU6xSIgnY464gly+0mhENjdg7Zjx
oY1h0R3VGK8iCaTFLj1R/TuK4FHqWXEMk2/pJtfwF9x4uE3Hw3s4akAVihrEJfQY
rXsHtTMSIwjQOr/IvTweV+8RRPDgXuOKuWTxY/JR3iQL9/owBGl6iMqRKKsfw4cc
veA+b6JybrFM68dioe5AjhZyzMZw6WWAou5XG3mt5EnwDujOjq8/CAFHhBiHYD1o
9n/q+MPyJGqDCOd0wDwKfUh51qLnCnshZn1B02qop1yD3otXlhddDdbui8uJFad8
6i1YGZKQUN1BTSI1pgxgBW8/teeDCNGrKcMS4JLHii/Sw1yjoGuXPtLZjQTXbrgZ
R2GP/EIpYpQk9K4MoL4AlGkbsgzg3ezowf7QgVuJiPhTx9Ek2aJ1Bvl8fnKPvfBm
V/qZQ4BlE7EwYqNSpws13N2EuPCMtvxl3R3aXLoYxq7+F3osVCpCZFzpKDhrBkl7
OYvFnkITfE17WGj0YOUs9U/e/nzEiYJu1ZoLiwqw6f9lgoUwu9N51TRocjG7QVQd
zRRN0LfXeYkHb2AH2pWii45dFgOfeeHqm42nGhV3ufsrVh6pBeTJlcZixN4OqKp3
k9QBG8fwvtlOzeJlFwo6vz3aFCICIMtH8qwwcxEepDN7MEnjTbjTH/qFlDxYf6EM
+VkOWE5v8/s5IBKbbsiQcD8u6L2zPwVAI9+gADNcvSzXom9xJIKK46SQhfX/+3R6
p8gkL/mJMP8fHi6OMXK2rE2vIfAKgoZBK+W0d+m7XG6UA3JlQfcbb6Pb79pG9IyR
P2FnDuZtl07YVnw4NOiVmI3rDRX7oKDck+SEbEN0a2+ovw7utwlngEOS4AAq4QJU
JhB9VXoO9m3S02k35yo3zWjeeFcZlWuHbmX+pxi0/jT0JESYYU78XO2PlJIBIMpd
G2K2T9Rc/ZLs/pQ17L0qqgANqd+qYFc9rE+EDQxCxxuzpMxI5wYqPOVkZtm9EKig
cdImD6zOX/YVIyY3zjHJRf26AsCqEnm9uLurMrGjIgrnMX42zZIf+JdOB3mP8TBe
yebQNXeeZMWMjfuTWhekDXRNGlHaRpiAlWqGCvQv64UHXry0E7nWV1zlUyGnp+P4
2UZlHelkzKNjCAr5vKPDGDaPU9qb/0KmfdLmGPtdgVYY3/RrKtJhbIgATTpesVJf
cP049YLX38Ieo8dNpwkUQexv9zxVrcopG2xp0yjSYmdswAsrKg/qf9IUjrcPT/pb
wp5tB6DgwXCZJ4az0nZtNXwpEQ1jeBUJXAGoEya9ME3YzCYyoavLxqKSITxYipCC
qW8eFw1L4GDMQSe6VcW6e7IIJWP7RRs8xSOCqRhfl5XMcumgzqtF1ReEuiWz5gju
C91U9BfqOoHKClRY4lpTMZHwV2UFxI4QhRIhP1Y/CfqFtMjRlrrawW91vupHdl9L
MFszuu5UglHNAiZKAOVv6yPfLUOOdcnyHEjhfilb4LkPU5rFndhWP5+LmCqUTCb4
sp5G+WWl7OB8JOi0p7hzeX7+GBkYYs1qKaKyXKDKf0Fi5yypZBVi92sbmUBnyBb0
uJUo1veINkWOoOEg8Sd9nm5eTrIwV6JyoEaYDiDsqgpE4A6OIdt58XE4jDo7aQhk
JNTOUeoLfFR87dfbVq/vfLTJ9DScQb2BANdGbxRoSoC3EgTCuWFIphRFBpqnPbYY
40fwfZDJQxoYeYcS2iT0rznMCDTrA765rw8fynhuQ0fxnG5jEaaw3WL/5VUa3P3t
fu9SNq4NecFzOwQriDoWY3x/oG8+vQ4M0hoxRvt8FCLUz4oxnDnOAduD8njc+TgO
W7DJX9OmQ3CZdj69HBbHN8KaIZ9uJCxbDcjnsiKaZpToR2EDQxYdVqgtRorJwbgt
bmDhU3CLIyAEK/aAOyqjGyGz0yr9LQJ4gd0GPwcTL49nERDWiws8JdPn2NIPnrJw
S4K7ktRGlBW56jaQ6YoJKkLDpoM30byK2IaXzNHBn6d+QHVU8G7D/6evxltVVBK6
g3m6k0GIoWIzR+gAwY2Fgsdvq6gCu6YCpdDnQMJaI+1OfRxbuNqZFuydDsO8fRCP
VWyI1mPMgv/VTYT3Z7cpmPqXSXB+gbBNenh92+UqdOWqNCaYFVTaEVqfj9uRvPWz
AISuro05DlV9J+hFtf3WUBavt74qlzDgZFFygGgBxP8H+AC4GW/ZPYejMKN2HGDd
tYIL7YVKeQqjmRTbXue+KZZmgvtFxqDF/GfI7nCdpasyDPLgKtp2u3+7fhEPa/7m
7weWyW0NUHyjvUI6aOkWbIUEl9cxTDZ/n/h4PqEMfkmKbkZEeoyvYSSavxYOR8hC
lVR4cDNRlcFcPOCicam8bDfcsc8D6GUnMNjEgo+8nJbImxTo329pR6szMXKrIWih
9WyYfdyF8aKX5EjfCEaExJbgBO+CI6QHRae1Vs/y/cbd8EXBHXGY0oWPKYmdv5N1
QuCwQYvtzA+fh2QE/HpiKDfDmLA3CS7h04vG6OgVAjQr40GMEz2Oyp9haGadH18o
BTK4Z8KvJGTYkOFelA2Iz7PrY0l23M0cmY+XumMWXOgzf0nVFGjyrGXATkTOghes
dTj1yKos3EMhUiV/NiknhGUaoENhnuaIcy/W1LIcB4l8tpsWGbvmWpDgf29tKod5
v9xfTvZnVDmeioHDAUlfkB/5SK9yZyllNwyM9utLF6uZ362odOypRQ0sBD7atlTQ
xBbpL7K+YwnO/J3AP4Jkr7rmddfOTCLEH/P/5dI2tDFW0f80lrk2E3n2iDH5WlgX
pKfeJq8bpafjrwZeCu6EKzvRRKGk60b+EWm/9bnV7NWZsFQkJFOSBkzEYmpb3Aq5
KZtDa6fR2WEbVE7+oCDlXDKZgClr8AeJpQem4wRLRXoukPATpp5I31tNaT+GrebP
2OkmmzEYAewylJxGZoGSq6MQNhhJ5MtoShvP7N3sea9TqKGQWPnvT8YST95z3+yH
fndUJxQzicNLrO1kR7Jz82pjc/eFi1Awn+TZqNJG6hkP9HpokkjRZDAS6Y++miMt
7MXFlIhDbXM26wqd8+DxkfevU4WPapC6/MGn0lSyOgGMyuFqsD8gGInxVQZAa1Hq
0JBfQOHgVMOAycUbCpwD3OXzNWjj+4HvSJx/Im5z/yG3HiX3argy1xp76kNrcDhe
nF1//dspDgk7VPSyPRmKCutBDEfMiZhONUuFXxHyxm6lZVWBM+C2VOsx6/Uqtc4v
pH+dCclHfobTV+Ag2l11zmzvTJMH3kq/yN0yyWeYj87RrsW+3M/oY2GR5jpBvKnI
v6TEZFfbonkDZFBlX3mONpRDzmBXRbB27fbmcAnUPV6T1N8DStxhV2wZMD9J0vJl
ucrmSjTWQW3gTiHSl5MZ9D0lBijDfj9Wz0O7ctGqc9yaJetlg8CYsQizL+s0pHtV
vAVbb47vs1Ag4IgpuoOThe2JgrVMpu3n/gheOND6JsdoWIxyUDnncSDWSWUtgq3g
r3dDYmJ618kCT2zWMlPCEIjG16zyDGp7dMrhtsCcJ/7CK09T89BXp92x2qabYzAt
DT7XyEskThDhb809CP0u+kwvV0sjjM+56Ybz9FZxWIx4zrj8QcBi2vkqHAij13Mo
+J+MckN8exEQbQvGltqqrVDL9QEZfTrla45UpriPn7fWeP5EeB9/Cv0qhoLiTOhI
elpIZt4NkSovRLGsL+eAt0PGMDiZQOOglsCwS8mtYc74zlRNtZazE2ZKUXDD+O4k
Ygnt9XFbgf8/kE6FTMn4jidSVNHF5N4LcEHnvMjaX1gZQU95mutEzo755UiAAvBj
5gjyhSjtyM3MGUpryH4aJtBVBjo30BEwhHIGR7LiF4sAqy/lXz1tYgirYj0MNFik
9W9pDnp2mAK3uqmFkKeizMaunQ9yckRR3esupMUCC6hpIM5rNea1AjbKRhVfrwv0
pysv9xNtIKVphNWc5vfVKQfbdtxPhgy8io+LEMi8K//5OHaAVoouVDaGf0dV+d3u
bGXb+RBt0E0e4Mfk91T1gt0QQIIc3A3f76cyhMMSJE/e3yO0AiW4zSxYYZcCzLKd
mMsbziN5wdMPzZZ1R+irzIt/zvd+3I1bVRkatahQNEmHw2uw2D9k8vCR82N/coOb
IOOf5DAkO/yq16VXvlvtsygbIt8+HTH9jYAYDhUN9bG+RdVl74xsiu6o6azNtiY5
e6AhCAkeJglqafp9vSvccTRiWTiBID7D16pJcf8D9MYUZNzN+SWwTrIvVBQlQrwb
uP6zOqcZbkC3eH28UZafdtTh8jDyaykGpNTRUhtR9EnNvWAO5oCUlD9+ZPwJAZfy
2n0yRNkgIfitJGbxrbmklUH0NyC4159CsbXMgTlEPF8jl1Ok/xsFDpLd5IdjlGOO
Bjjesv+qYhgWv98pNFUifoFM/QobzV+GSERqL5PHUHrT4yG5WkaCv2AikUjJ8fOW
nk1/9zqqWkZ1g6ow8Fr6tpWDq11FSjEhNeHl1GzUn1e7Z8uvTH+lp37GCB1RzYxX
eH8sqlvpXCqV2YwQXNm5Ym3vCV/pRFj6D0kM/dX/HWiMkbpzH5E/iZMB+IasOkUA
g7LFl/Dvc3Yv9li25hldIxb4sKLW53gFSPRBEQwxmrCwkvHzEe5w5ZVH+lsoJGMr
pO+KJvWpdSS1WTdvTFQgwHS3G/QIk5kOx7pAqt/d+3HMBFx+ld7czc7nnFNUEx7I
e7bN/eHhOLOHARpGxiCwXO3xoBQdnM2n0hUijIh/NcW3K0yAfJ/28MWqF0aH5+nm
+U05jmrZdtlzBODKv1oIcq4ww0LPgOM0/sYitEdhk+ZQk4+bAaY4vG9bKlo0Pq9G
OCgrTxgt9lVH14/8I3dMVsUI1X4CNFU+OXRBbGS6dyQx3tExbYn9uG5pviIiBmVk
WoofLzmbsSdQY9nPwu1cuf3xvhhBQzW+uOuNi4QAKD0S137oF/cVfTEyhO0D9WvR
WEtPyEFsj6CpFei4UmJF6yPapsPASdzn29IYvNFAgjJdagowMJctIAVardwNw3lA
l7PK+ygWx6r+uEVLN0DLwG4hjL4lvNVV0FKCohsqTZd/W2OYwyRtq4hWVu8sHjkD
PVIkZTbK7LQG5ICsBwt8xyu2edcduUXk4SwSwVsQtNIkDvfnoHNrE2t4unYLWxDS
ivxX7BGqbiMz4MRNPnN0yoJQDmtCzreuQnvFZ0wCh/VL5JOvofnAL9NbRU+HnS8T
QqnmOqF8UXXmXkKyL/W4sbS3WyI+YYxTU0qWf7zgvzyobk8hZKqGIvxyZgzkbbFV
EyRLIdcVgjkSPOiwziMRpKcTzaBPjI1l1L9SJNqPozbl221/i0CgO2HGxg5lPp6T
aCgkp3biI6kFdP/pyyWfIXoMLqBaAsAlmmVhaGQ/GemZNm97AOJFMeq1E5AupdFa
31rbzBqfSR+W9b0TattJki9U/TA2NbayDODmHQ+sNLxwFraTcVr1ih+8qZRr5ffy
yVgDdoU1+Wlo+IUTcZAZAP21R3h/KKkWqlQXdn74TWNFi6s5ecU0hZkF8dvh4nok
ZwC2LG19SwGNeMqQZz1Sp/GYou5jTW4rqMt0oTGqcBGrjrItHmlFR3TW5+mXpmDL
Er+wy5u5NO2Z9Yldcfi4fsDmCMOLR3FGRpcV9n8FSHiZjLOl2uuy26uGqcVxotfs
2Q2Fj8gwbjs7SnTwkxEZzBbQn3tyMsC5Hak9npb1m0WUpo4zDHNxt0cdZ7aG3/5w
m3A8SKMgSNd7V7Sf9jAH+cofN/GybiKWkN9leCROI4v9pAthihJEXIVbxkzhyOB6
It2fotkqqxBjKt+3U97G84Pa/ydSWw7PUDypssEcbF8RtZUExu1AhgZLw8T4qA0E
UX/uu7I9uT1M0NXqWXHpg47/GPPCWh2ju/Mhc4NSox7ox0hmjk48ibgUyWLa07Fu
f5ORxxkN9jh5ieoMfBkvCP/1l/qgmG9blAYp/dpKIkbv53ymYAVeGPaz+EZeGVP9
+ZXC9a/IenstF9McACJw0gAOoITNV1IObIquIV87b3ozCVDYg4jqrWmC+pexF0g2
yiYmzzz24eIsfhOBMzqv2EC7tSNWI1rUbIeNQgqmQ1yF+zCtVz7ALQ73sB/uE9eV
Ts3Y1BmNnZHXwdgCyJxKijUdlO1R20/JCw9O5slxRov9vFUEUdvMZNf1/1LKeQOt
Mq2dGuJRobmeHSC1pMrHI/ti6aZUqa1Dtnj4ONgvClZRBrn8BA7vgA7/Zv+p2Tvf
gt0yPduELIxxO20OhEOspX+oVRXmVRJNsEvTu69LhdM3bkeFqGzc19ww/pB7kJ0w
9MnmkkqYq2CT/31GJ7i4EvGHEKJNhgCZPzwCxUHmZMcsCmVcn8wYFsqYR2rqhY5m
j71V2nzWBFM2WZ/R4WyFyNe2bPZRL1QEs72PF20zECO02Lf67n08Icgj9x2heC6c
Q5clISLbTZA8GIiRua/VAQ4zubUXRgMb81zYqNNDBJxhftKr0OstmxE0Q8Cn4Pc8
m0uEDnJXNTiCmtDnjQkaXhB+tKWIcs9LOIM7Ax3DXgIBD1+dji1+KmEPeA6yis2W
zWmEtrC+RjrPSRBZQi+sKnsSIDozeFa7CnqMhRtpHqfsiBDIdhzb+kgh2zQsa1Gk
8XvOy47r3aX6vkXF5iKki3kxdZyNXI7z97GzHx+GbfsI3augqu3GtcM/Ip+Xz5OU
kagu06B0S3X7bKy0bwZhg96Xkx3/duTX28kKkZcb02gjgDT2ZWsdE+jgDIhSNHUx
6tvf+rvq9Z2cHI14ywdnxT3UvmoryOQmc+s79HTJ4Ls1ilfC3UvCHOSFfGxXBF2K
fPE+fZqNrImoVKwreSkSZ1hMvZTFlF+5yzLlzRKOMeRyMtXu+LMnbvQFhBKfgfop
NrJ0MUL5LLqETDuymdTt0e8MyBxmdT9//UGitDKFborZOMMYyoNqtvINGtVcFMPl
Z4IA/dUAxxY0AkvyvGnNwYY8o5aiA4W4Vvb+zpRFqYeB+vQAHU1znU048136s884
0bErlFUR8nhNpJRwS/2P8/YV24+IeXgsMlB0pS4vb6AFh1k2d8E3tnYhGaIw2i0E
39dg+Z6BPa0Ejg98h+F2IU7YcscnQN6NCxpfPr6XifxFOUC6x/aG/0XrzGizAJxx
02BsgRDDayn82zjsoLPUeeoh4yDRYQEF0hgAS4Q70W0bhjb4eQeQ/rTLAmXPdNG1
wwGU5zGiEUWLG/bjrI9XkMxgjImljK4qNuFKQXTwzCUCIFBCZiuHxC03J/LXWeOt
R7BiaFlYWlL92nblNmFaKeTQHHf8sF7jIehSijtcMm223ClR9T5BIU2tAGLHy3i8
ZHq0WSFcKMNjmXn03d/LV59IFvzzrDagYoe92ajljGAZ8BDBOrttAYv7etyAMAcl
u9+jFvYcQWbXLE20EFqKMbH9Ww9u7qaedwRd6j9/P9pThKUq+gtHwlt9HxNo+Gu7
d8BOJ3+8QB0jrBSrikIOmmJ6P0rCgrHFaZzYFYsfWWuanAHTx022WbwYd0owJkl4
tKHlC6s4OStCFjHCKHI0Up/KHX4lDkFRkzLm/NHYKx1zSRONxgvYRFEHJztVqlub
M/bsNePEeVWJ5xE8t6rUEz72C2/VP3CbNnkpzDOMVShDqaszh/AA1g/8cySCOmnx
88/kqbGwkAscqMIr4/ddSLe2kQ362CtPUBtoULq6k3rckT29wWp3OlY0+iltzgS0
TXdFZqLRftS3TjOLjm38nYMWXlRCxjnyYI7vgCN2vVo+CRgk4ufrpbJZDwjWgVRi
wZKniJWxfMZRp3DhekZ5zF8lhjuEKbiPnue9XlcO2N3NSpOsnv901G/0KHX1jIKQ
sBkqBhDxWXTXACj+HrUtXvMuXhu+ekbsi6lJfhE/hbpFOnW3bMQICHDpJmdLTyvH
gIlCqh5ct8y3TjcOxkowXR/C6eu7s7SU61D7iQT7KQqx6jadbHVwYiv3zMIn/OKF
jNFVu2pYEUbuWW9oAspVgfMwcexP4MRwIHJylJzP5w+1A/mLBkQEwbZcJoroPwFS
S9cgaNbb2pVDBSRs1RHj2rzZjSSwJSsfO/++khMGfvVXX+2wMF2UIRprhEzeuxDa
Bp6xXLBy7TbHK4ryccJzgA6K6K6nXy7rp5rDh3PCEEuuvETi8zW09DQDmVz1Smcz
35/TllFY5EryrJrBI+fIij4OKV/0Vr+r0OqWHUvKSR4B0sHqkJLYYcAVXFVF66Q6
20qLgv1pHibXoGu4SvPk3BfV1NTWDLoRKYI5msGMC5BudiLVfsPdARgqFSJp8wpY
jX8QBItNjzANXSvNrb0CD9rPWPBdQFkFyfqQHTxeUljcWREWXXlMLzdWmbivZ3Z6
lOqU1YRN4IQ2VQEB8dFvMSuxaVDcMFBrqFY6ZeCtsUg71Km5UfLgHAmW+5nS5s6L
Uzyjzhr/ioGWdSRypKQE9s6AW97ZAp+omw+sKqjyx7K39d6ipbEGQPp88GM0FcKB
dUJPJGhjHW+sciQAkmCKevWV/vSbHdXCoXtXP+z9DukyY2Og1SUMVq501ght6BiR
SCw0nqNJwcSJjNcfBgHDqK166Ywk9WgeaMyLosI2lzWPIH8leRxnVpxTOsL7Mx/z
uymPEKEaGjm5E0QsLWtgZ880LrYnCyyX27NbcbXy3Kjat642v0StQTEfP3+lhI+R
a+YN4KpvGMICvH8s/T84F92n8wKVvzv9PlV3sThhJ/+QFLeKlVZ5W8n4lm3NcBCU
pzLcrrnc0sAO0l0pgcu0fGkuQpL2524LjIFB+hQFUrrW15PDWVbf6eoRDnDl68rj
yUy1vQuiPFq+8LiDS+ACFraM62YM/mp7PxNPcd62iuuMHq3wa21Qvf/OzI09mad8
KcT+3wDSKkS8eJr+hEbCAoBK/IrpIsoRL7vvsyC+F4YrwmTXGil+oJJzjQVhmkqi
6nXYaq50e5efcKzfk7BrLMonAU56gd54TddjJuRltYmo4+3fq06vLBOyqCoCttzW
KLLj1zLsWYVyKbSAc1wLcuqv0XBpGLVidcD02Jlw0xqDi9iCGqyliDAZte7kipf5
0aNnuV9gOqPD86Y9AArHITk5GhjlGa1pkz75jL8zZJVYSba8SGl9fS85kPjsk0of
gBGhS7YCoB7jnRxgxrl/IJaYan/pA877Bvy3dFdXB11AyogaiZaZJz9nlFZBsh7B
C0U/EVFYX9Y07JLDGeHNom4GLtpuhh25EXjUPfw0IS9qZrNUKYiHPx2SRyzepyPk
Fh3xAzxl/vS1jL4R1pHisyvQc0I+C7Z1ENOmf7pbQe6w1LEhnDUaM29cWv7S0icw
Llhf+2wDASfJ01yRUbFpCiwd58ECuT7sS0MM4PIjIvN1/k8EBucjfBjkx4qc1j6d
zHXUOnH7Qt17Teqkv0WHdSoH7S2TV6Wrm18z2yKYLw62t1sGHKRgxIxYZAcqO3aa
d1Y4OL36m/kxW0wDlShlbLrYkFU1L6RM9tdkTIeOHafFE8FsucQzZ5HZ+r0Re2n6
oQeAY+J3XYA7Rhz4ciDpCSMHewWhRE1B/1rf6BHzjtZycnGBsDmPReSVTWI4Jp8v
3W4mL7rdBm7bJ50WAXebomnQaO7n9/BWKwvY6HFUiJqzZwrjOBl12ZCbYOgN1rUh
QOvi/eUVA7T8yZjsLiMmvPIkD3oCZXqDQTHn3L7f3ZP8zzccmc9BxVhCOj/ejGaJ
jfZ5poEJcbLi9e7SI+q4R4jpYJnQMUh+AqaKqUEHPqquQIyFOUybscYWnbpjipCM
Yvj+7SOy96su2iXNMja8EoZZMshXtjG521o/PsgT/nA7HUTQsSuPFg/w7+RfiItp
oBO+ggq4UFXKnfU4J9XtA6aGBRLPJMFdBs16GEGTyU4+omHbi9P2l9EKOUpbxCit
0PpShPl4IuCDx4lqCUhuveGdG8XzQ0A8nptxBzp3joz6tMfTAilVHAv7PAYRPkGC
AsKu08B8PnqydH8hWPK3yPCgLvB9ni1Nzar3YJRQGOFDuxszIVcPBOjiaZ4UdEcT
KbGgYZP2iQeL/Ii32iaIfTjRRQllfk/aTWKhtLMyT7XzZFoKD/fi5G53hKjRmfvC
n1dlXPNkyMVWCb0xy7/zo1a7G9IDzS65rkK3izrHIoDGEG7TUh0VqxH6Ett0rchG
O4U3AiVtJ8IM1FvqJveuUJLmjz0M1TCFXCB+7kOKYQlFb7/4aZoD6eX/PKFuFHXC
kTKWshq02lVQu++T0LuWrOBQeTRjHU11E4pFOqHiQy5vOey0Abc7Dn78ZyFn5y2i
xIOhKZmKc6iEYvDkF994qA83lnEI+/Og9FA8KMWT4RBb7slTfifZS0UUgVI6+pcB
Wh9qlS0wu8xCDGE2l8ZzrY+m63zHTufd33Qhk9NRQDTy0T0WXztGsmQCabe59bqA
+2jwcK5327CjLzGRqI4cwglRJVIu6tImpmc9PlDtGAQeUxrbQdP/i3Y2NH4ukpaH
h23NAN6APcqwtdTjSbWvDbtGOn3JsmZl0iXqXQhBBr36bzoLTuT267zKg0HgtUi3
hnE4qVUucTm13KQa2VEUNyu61YQdl0VypvoYV6Zs4zQ0B4jMkst+LrYCbHr27oGc
Vz+6K2ysGxxRKSM8FzVDJk9VmEdMrE3pj8VXD7I6MyrsmleoAjV6sPlNfwzO+cUQ
iGJwR2iwlv9V52G6WWH8mnbBSp2XlC/NOqbBgxWZWmda9ne/lpnF7icZI0m/1wb1
nhX6BKMr4MCf1SML7etgEDWJG6U1PTVK0ij9xAV4sq6qjqRn6AgGbCMtd2zFO1Ly
7cAlFAzr26RWgkB/bWaIch2ncZz4cPsx6TPUepSNIZTF2q24ZyJ9hywbwzoU/4hi
B0PUyiL2oIhYmw+n389oAIFmgPLDIoQ5CQOjqiJzzg2jdZuJKVx9EHUkkt1lbxzd
guQ9yg0kpqxDXpsKvDAKnxA9kY4VH+IOatfkAi6F8JW47bfh4Fg3Saj2qOj8QcDj
R0pFnFBxMoUdZZM3uZIDurjDFz0zbdvP3mbOifMvS/qpUkEmTYUUf0jcgk76yyhO
3nKf87bUUzPSpJWj9wPCvjlAuw+oWKRufoEowF+LldQG6j3Wa4f0idXB71kCpgdH
3NJiJsgibxT6nxw6rvRzpQvblZn8ybckZrB7xe4ptJB/Jw5xWrDcPYP/spBJZAa7
RKHkQ3+64wuSCjrA7Ea0kSZ8ZbhNLZLhruVNvshYDry2yNoR4to4AWLESfM8MfBR
+7dePCiyJOKhW9x2Rw59ZxILN2WIIWRhmwRxzeHJZ8BijPTa5c6ENzFn8CG9K8ty
D471laFZSHPD08+5qMNXgPh8dmM0Xl6PEPRVeQZNnBHOe/ZtiHaY/WzJC5YRK1DS
6Eqv0mC9wS5BmddsL82ES4FaSfUJPbK+DXkWzOuE6vlMEWpmbCOU74xGAzly2zeO
iSFpYjhZo+hL5+k+PKUZCnZb37hZnSjAUPHVq/NdB51+6fZVWdGrzSjHww2/VcGi
0RHw8oxQgAhia7bY/P4WYgODi25DIV8cwkhO5pcch6xCbINNAbbhM2tHSc9ld/PY
CSaOwD2bAWc6LtIW8Z5KSXzdxmz5X6dUwFEqVTj3xvHTCNlItk+ltIOE6ChZhPZN
KtouW3aY6055JF+b+wccGFpArppRqC1bEjD9/Rvh6o+goj2h9FjpyaqZWWqG9sE8
3/J+z3bPoJCRbV0lRdf5weQwv5kpPYzi+Tx1Dwy/ZOk8uIPsmwWJuhYuctNKQSWf
ybs1qGGomZI6zhhe39ExXFRMpu2ELJkpTUn7IwhF87QJ4/D0RShHHv0jjcwtDW1N
fY0vi3ypmh+27FLduVKlpfB2awhdxEE0tb5GSOwsTgvYSxSF36D2qajabcKPBBiD
nhJI7vviO9kRvL4Mkc0SSK4IzAyZV1TZJOv+qG5y1xU3f1aBxVSxhREMa82o+EQG
Pz3tl6MS8wkqMMu4LBl9FVjGjIkmaDv+M2MTPoYE2aEF700VCDH/wgdgU29+JSq1
dxfNN3ONR9BTl+7jwVWRzEfPxYOTxghbXFWLNZ/sYS555HxvmH5X+uwsUAaUEL1j
r1tl1BDmZPeSpQn0zExuEo4p81qaWde+qNPsbQ4pPUeK21R6IFfB/vOhp1fFN0S0
cEQPYsTuEGrl9xmebgjWgC6yBWdVINDahV91sT1MNPvWvGbuq08DJlzyqoQZmwmO
BMR6DftWzdk5+BPNOd6NyVliTpxVv687kQ47VdDJfCRp1iFIXn1pYvc2kz6q+ks8
y/DxsPl9FT+yMCRmUlY8aY4krqDXzjkU1mGpMRM04m4QHaTH26mMJi7dmgrcQUfF
43TDsPgkDz2kcSy9c7tTX8OL2X1egsFfcpjYD2on018rk9517zTNUvXZu76+21wh
QDisBcYkXFzkSOjEtOIsRnLcRsClMb4mSW7gUtnxrSRfGg6OpCmztLaAFcQ7MAPU
eX6huMgtVgAHj7T0leX6KBbzUqPOzkL1wQjHh7zMP7au7Skz/jK+eCBvIjXOWMNf
Nu0edygBavn0EYy8lRvnGUD/teydD6ElufnZy54/dsZKA689ZKwSwLnvffAKuA8n
nUXzkKXEFQOVz6t0vN0dZMuimdwDfNcy/QIP2Cm0KB4jDJOgBfskvSupPhY68OrW
85+Z+Gt4rXWexNjYE1G/vQ10fEMMijdqk9OkFiSq0Q3HMRFNRpbw0UC6A2CxGplE
Z8lAV1pQ7ZCJ0c8FcpLWvsDFDowAyHXNRN2Og4YAUZVLqhA0vn7oHJv3a/JG/zn4
S7VA07O3iHrfiw/PDTgNULK4MF/QnkRibTDkSW5jkoAQlE9ZW3pe1AiTg6J2BCOV
Lz2Y2VPXsChdie73/ETCk4LWuFHQjRkvO+9QiWNA3fSDtUqHRSKB5+PLs2o+MWYF
boufeg8VOOw3vpuCi6FP5D40if0BoEcHsqvZkg5Aqsqiyq+63Xia70A41BBL85qN
JHxqguhiZkGryow33JtwvDA8VR86RDlJvE2iJdyjAtQE6JpsPS3wCW1YCipn6Eyl
Kz+JMvBFUT5CJXUx0F1iTW0c4iSeWdI+qSvU63isH6OAN5zjjXl0dvgLEz0AGNep
Cobu0sroImE1gAJRdU/0FnXT/oTNntGjYvfTbv4yfCIME+il5Z+oCbdpyar1+w2j
mDXI76nZZYScUk60gW6GCELs8BGepRHTrjOSjHW8gdWQiFyVpcZVqhzhg56wuVSJ
nkrpfmSwOScWZP9b9Ip+YC3kJv/gPdYfr8pUNLm6fFUTBbBJ0jbY5QWaT+kjjtEe
N6yxsC9OrrA7HI0if4XXV3l+9DmQx0GiPE896HN9c75M9F5Acsj7RCj8x6X3CWyo
IvMyq2B4cG9T/5cOVn4Nw2Oht89QJxMoq+xWf5WCtQBb4S+QfyrN5DQmnnPMq19P
SBhl8ek4XIMSmA51ncjA4Xue+NxCZ4xvca7kd76Vh8WyMmHH/JUTxfAwruJF/9Wp
N/pr0LxEeHTwou4mMXDIrev/sxMQLOLT9s+0FcFRv6Ioq357kX3jVOmnVtOtp4TE
dX/LpKcTcyQ5pkO/pP7p+LZy3gzPs9doEuyygkfe7LiJtFFJZOci76id3D+UxNjX
190IUeZnskFOzL5Vy8po/R/Zes4RMbNxvlFIeW7NocS/YYP0mFD+CoFm3WrGMZvX
sCnHloiFgSmxzJ+nbwdCyZzQG67FdxT5ZXB5udvg9wIkbZ9mDawT85rB4W/vdteU
OhdXZ6ecBFyHMfgRJPAcyRaMJncaJHaDV4X92Gf4cGxWaGEq6bPEGvIBf+XLL7ad
3a6Yku5AOZwQ3HDOB5QMz/liNB1mi64TdF+GTE441b9tJ+6P3LZB9sAlmiBRDygb
1dpOsANLwd/ZgSLPf88b9fr6biP8Zp9t1ziwVy3lJNKKxVJ8i5dyxsXh1WmxxGLq
LbKZ7jVvWpW1vwcX+P9ka/qLy7NL2a7ycb1q7XJCqiTvVb7asU2sLUv0a/1g88EA
cO9LYCne8Q+YgWI1f3iGJ5pUBXvatMJvLyngQKL7ttN6iPFEaVB4GnV9YhSxCfvo
sWUZi9ogZhwua6PBVO4UM3IcEVrOHuuaii2roN98sNCvopbVCiZF8AZC5kPl3f+d
qbZDro6UtmXjqBPi6hi+yZ+BkAKG+HJVy586a2+Gjsp7nbvyBUo8FI2xn8rbVflw
mDI4p5wZyxQcI7Kwe1tj1Lwin18zFPiGX7yciUb5U1Ll3fibhXv2e71C0Ct6jc4J
emT9sQUZjVMMOhZQqAtHSopfT6I5Fgkya9MKQs8WM91UOH5ox9sTJ6ElRfCTQQeR
fGbsJ1oUzQl3zlEJsuU2FpQnRua2LaBuZmYxsSq2sgfUJ+WzCQMUvX5UAOw0oN3x
UPf2bWFjEgu6qkuZUwGOOnw4Fzkjveg/VP/3+up26Nky9f7OKRp9V2k+b6WwCAjr
tdFJ5tpI1VF6FQxBMKR+8lExyf+nvzMtBZMaxsWEyKSuyGmaB+PzWEElr4e0w9U0
Ff1nRM9vrxclAWmPfMTTO0xVRyl1SgKF48iIq4/v+2BR2nK0+A/sxWL5a2WzG+Wm
VsTW2O9nX5pYg0dBVz2KjrgQGzSJ2Jgw7RheNFyiqrp0GfEVPY58F9UrZ9xrL1dv
+qeAzBwqtngKiPymj316pftQuns1orAfwkrx8pqWX6LDWkEyxPDHMKpcswsr3CMo
TU3b2xwSGbCHcBwhPevQPm47pHpdI7VASH+jJPt824zwM7v1J/Bj+afhmbuL93AE
PGW0RDJLgcrQRhzkeczfbWJ1HjpgAJPkj2+aA+phzzR7+oFkss8CEwKcjA3Xn7a4
2G3nAs4E6Vd1jnAzZ6hzVLB0jrAdjTTWj0YKygXd9TmF5KYSb04f+iXejQ2r6qlv
vLlEVcTISCzCPN9goaVANKKJdc9tg7mM9pFIb7SaHzlS/JOWf1c7yyR6wCew6O1Z
xH0iRslAt6Yy8JW5hExqH5BQ81sd/Th6w/rozdmbSAyhcdiYDLmdkogKZ+4tKTv2
WFdoK3l+WiDxX0ETk+DeTBWe5z1QJjFt90T+woO871D6OyL8EAe9XvkDkFO0fqZk
b7EEZ2De0CFjnRLxiv+Egh1kpy3/c/iPQN3iz5uQ3QGQWzpL65kDQluZp6mRvp7f
aldPbk1IxvayP9Cp3W+kTTZwMqvqIciog2/xh1eJwxNXUSx3V5X5tkh90P/OzgPf
uoa/69gqJO0fg2vKMY21NBinKdXIju9co9/W1+ejrPiBg5isbrhlcVjKkMzdMzHS
dMT6X0W1BHGMdybLcqCxDaj8/iI0PpxDL7QqLlWn+yj/eRXDVXs91TvcrNpvl1F/
mKc5UGRp8NFo9HpLdL0ccry+ybG6EOOfGYoFqY+Wr2FJJtHt19qMqQbY7urgmuGy
CqqQ6HzxcgHiN6fssX2gKMNSZHFLiSPGwG0TenlMMtRL7yOmWUzNURyPxO65W9Y8
i1shbC87LL4QJ4hgCYUEFtGndVNYNQB4oEE2Wsel9JK00+DenhbsDzoWbZhap5GC
x6YsKQVVY6SomHrjAxmpiMHUY2FOZAeC9VN7vxM/j5Lj6VhqStQ7a0PWFy7irNC+
yTUOWkUH38ttNVIoHCltYUH3RQsymgXoDsA4qx0bBEWxJtWTRIW2FKMLY5IBHq/1
brcS1DGWWE3zCmmgwQxH4FyjNd1ewgIlwCYwwu8FbD0CGfbA+F3KSwvHrMdt6ZUN
TVfoDMfhAYmjLYL7gAzChcQAdSbLZjsSZhkXZypOyf/djbGep6l0+3jpet0//sWx
YbAqh+2MpoB/3rChk0s2m7j4yrfbZ7wTZoOoH0Hhfw4W8ZAfjVS1lo+tQhHsVC22
qtkvejO42V5r9KinGh8vvKMpa5GQczd+FWK2tq1+W8bFQK63VIBoynu5ET6TRCcP
/cejRoY+iicPdU1w0tjHvA1ot0opepKK6CV7bgm0P10o1S5YxVplkSCviCm96gOy
5Mr+zmfalL1lY44MViNq2CPwbJ/rPpvjwlkPmeEyE1u++7IkWyz45ct2oWv9d0KD
4bWHLjs7UVFHzcnpWjwCafzjZOHJi6MPJuCG2Zf6cUs4PGD368nFHOK8gK8AU/S3
39DdZEr0Ub31A9A8OgS7KlimAPoXpKuTIrJZ81VPWIJhd1BeveicCZ00YWd3NiMX
v+TOzBiLXCerGP9JrFhRl4k4BzXuF1nHnRHw09Tie5TDVjkspG4TAYBhWIXJZHe5
l0xa6V5olaePr0wpLKtnFgrRMOLmy+ifNMwb96Xx7fxETXfdseeoCiL9a3izuT8x
G+mW0YuS8LjcUiE/XZV5p+DPpQVE+o7GwSGi/tHiz+LcpilyuKW/J8rAiQm6rUdf
OremxUb4RRxjhqFh35w7ihTHWa5TJ/zcKMRyt2uucpdFqc94e7DX6v//FDGONMgS
rTBXGCs34PA7WKu20eY9IdvuAdLfTIsB4hphTcuoCG5XAMCzIw/kYatooaJrKf7C
mABetvzUOT4wdVJP6UpHibV1ilk1ufHqBvvMVZT6zwnJ4nLMUXTBW1cWF+V8Fmdk
cEjfjD2cBJnX2u+VxfzGzzCMdSbOsBCES6DZUFeyiyau39vCLYIrYJzCav1qNgTy
X6Ihus6/oyvnOWX5jE9lz4vVVlaQvHfl9xiZrJBN4Uxbs+BPqBVjxRrC9HlG7uw0
dKbMJJfwErYtI1xo9TuJ2i33nKCAJcX8jdJI0VqaAOL8KQuKpP8fbg4YBWV4UgXo
9y43qf74uYQ22KxfGjz/kso3IEdNlVn42ofx5qiFomjtSnIK8TURjK0M6FIPAoHa
bNVNu6xJyWySR5/RxyAT8W9W+35KlXpk9S1CS9quts8ZO4ZMGXIx2O6WcOHIpvw5
7jRC3TkgtCPagFVBM/fsQVbEsq3uI406tVkOy5Bo1EfdFm8+ODeTDsF0oxjqL7zC
7jR8uuRjrHW/Wm79yR/EA7pz4sRjoC5d9FkjvfqXusO+4vaP3xD9zclrA2/zEWoK
h4bcMOK9DHOvJ24enhX7et5dD7Dp7DmaPYwq8mdQfcRI05xeksgzLRNU1uVxXROa
S15tzJrPJrapNcw4TMP4VqHtkt98GSU4qH9QWNXbvszbYTLYOIRnQ8YNhltlO7jH
dwhdDJL84x0oXuEpzSlA0zEm5PX+/6YuRj1QwqIKI7VfYXaA5/3QRPd+WkqO84sG
Ts15qn6QhsykDDEjgSWw3T5/QoeIdot8hGMQflP/wJ9621Fgvvjy3wbzIrpWZrnP
vhKrBeUloVLK0cAhkEZiNNBGhUk1lId+CQYSgw31mtK8jaX9Z0+JCCO+yrQnZU1P
oZsII9uE5iZTyAeapwkVXLeiTUpnojBAkhgfDlndIuFKZWEfUybHh99FfN76a3Y9
Dswe9drR1v5MlXvjIRmgNQn+rppT0IBBOUqkwAkpoWTTnKLZgHTW51fNLzb174D3
RmgN5dvKxF7FGi1XfnlGTPFGHjlgUWUtBrMCNqfYbb70Cl0IcI/FdeAAdQLxFwNQ
SBwnG4yOhoVIJKvKwEdS+FlNnrfaJy8upi3GVueN7NC2Blo0SxIbeO9UWa37jdmY
/sMyqZqdCh4b2enT9NObJoCWqyosSqCE2QRD5USBWgu6Nam7GrnLmtdJHZPwx+cI
oh7r07wrQCIGnu8joBQwyKkqu705RwA5WVLZmlFFzqhtKyVNkYM1u9KKNiji4Geg
fCAToW5DJk4n5Uldkv8llUlrL0zd0HVpjzVjAm7zyHuiQhPs+gMGkwuvyviCPoFZ
gevJbV0zRGJLMyBFx6q2Cf5hzLbv/0kgORUfkJUdNTgy/JqUWzYMhuFWnLpzoL/u
kVIIK7VokxWTHU9wclr9KClJN3LcB3VWUHpCvPrNQOLXxeAPxMJVizFUCmEIblYG
8BzCUENjpUT5B49HM6gqOkcKTf27HRY35T5QkzkjLd1Ehw1M2pBrr/9JSZ5gO2Sp
wE4M1JAAjpEyKtyAC9X0xvKABUDu5IqH9z73p+U46nqAVjxicmoxuX4rZa1s3fZD
FK8XbxIDmNux0731zpUO2FKAQ8AirfOh0w6WjoLIkruUvUtwrnXCAXdQbHewCBeu
71Jz/tytTb3u0PxfdyNnbShsqv8bgeb75c+aoKVYRv6/FK+NUJAAUbJ8+4dr47d3
KYmJgLVMMsW2h/L/ks2CrZ2jBjc2pu6/Yo3lXD2eb/S/MD4eRSqITSHUdD5KSUxm
ijYatj/yOBumnxzlq+pilRY0UYZq1HmwHiXYehCFg+ACY2UVlVhBXCIh/BZmNq4w
+UZbWnNx1mMLJrKRaeHVImp50IMzvNdVCBijWYQTu44hsbx8DIV6Lgk+KNiItUBy
10bb3rVd0SY31ojpJTvuIQZMJUBaAQocOQb0lbMdkfZUrL7s4E51enDRo7o6M+gL
BKeegaIbrUOHxVnLPcjIhgITEHTXIGcOZBs3w3rY6X9/xOkYvfiu7PrP54lCUFUZ
+mpaetUW/zy//Dk2zHSh3XCK/3cIgqzTc6XQiAIBk4a/jPhoXTxnwz/LAVp3GdD2
5VGMEUvooAl8n/72D59isdu9gd0GU13T/jNLjoausLgQC1Jh9ROdnkmuNhcW2S0P
GMZxNWTJp8tJn1CXBaIQ7qfJcnY3Zw0BsRahYqAFdWNSPx1Qhu949skdE0QExeej
FH4xmL8+1Qb1Wyw9ER8Pp2BX1uDCQXwNglporIMASxFOtd+H/dlb7h6ocowBBdgc
6AX4YsS3f0gxFmxRZ1+HhXtUBY8gZQriJTy+D5f4/AJTUQoU2HU+C9RryoYa//EY
0wSlzvat4InJxdTkV1I6ZURZd7YBBpjWsBS79fX1bXQP/SM/N+ggGgopGxLsjRr/
NU1pLlefhTkLgMthff4LNnQwqjVVi5rKuJqICbURHfMkh3ZbrJJeJGFKxw3eTpwT
wwoSEfhn3KhIcxL+AR2ca7k2VQYKccWOzJtr8V1qafP12cAlFDSYZSm47X9PHNRf
JvmL3wmtzk7jtPVX34TRHMXq8DZuWIwnPudKIPHyG2DucnSovKjr8kUQlXwbqacN
U/t92IDFD+veCVVIAdT0xRdKVM8j0hwJJt3mmcGuPoXCPwPlydXLnXC42GR/ZMAI
tFOJapEd7J7+0M6HhhVVQ92HXstHswo/7qMgqdF/G759tO/FJovbqhZZpIk2kcAT
JSf9p+XUtMLEZziJcoTVRubSB07EVFI8XHqg/551xTXqXVQdjr21Ug8zluugHGvA
FdMyW2C8zBvQGgqnhHnA47eaCMwDf8+dBPs/NFTXKm4+o2TQq0gI3yY+IyA9oGjA
XC4tQrnov8MkxsQRCP43BNicW7vrNT/2zIbUtjfcBOtsP4AIO7VhVfsaS+9XHnKL
/g9UnRqFQpdkTsqZST4v1FgAZ0paPXKMEhEu3KOzrr7J/8A0qFO87GVrZ2Bg9pvw
k916w7PD/nJxoG6xq7knOH8xOyAVvLmwPUWXgRe0isEK3Exjv525YVPUsgkkIa3v
uKE8DJyPo6yxTPle6VK7NN+/ajgO+o2uQPCEu9zUOFi36NwiQMoTj1Do3ieJB1GM
Pnhdf+8X8SynQr35FnlWdZ9pAXGzR5BETsEmWENlVXouThK75OrTNOdXRpXLlX/Y
1nZ+LOPpvqjYGd1AuBpX/REOvBd9TUlgSsu/J6ylzimCiLZOv26SbqCUtg5BSJfb
zEsf3CQfYt1UHIV+RPNsRtF5FXsaaf7ntmakVSbtjeRPNkJCRynW8G5fSe//XH6E
1B/WmgvsbejNLUfqwr0k6NV7xDNyh20HYLmSp2PFlOWxTfnTJJFJeedNWgZ/qJbH
WzN8coixJFy77vNjObFn4FLdac7vv5mSKD2Z9zqmv2aWSPE7xudDioDBqc585eG7
/M0E53hsGMmu9vGNVLxtqsVm4pRU2DoJEmYPsxPVgfNKuUjqjjG52Pg/jFvxYgXt
h8zhCIXLln/3KZPn/sBVbBeBWL4kHcCqBSbz5xb360/6+8YUDOhCh0u1r7BcWkbn
v69qFCrfXNRTt12eO+SoGTlQ57wJxVP50Au8iNZ8/70AZP8BZopChA6gbZg3wld7
fOQ8XxX12PSrSbruYDfWnc/hjZApDqrVBN40Yey/ySEpk9JgzrdC6b9DHTRI+0u8
Dp3MY2uLsWMEOD/KNcyCfRk2HwqXlxMG1a2fQ/9DIjr+d4aVA/p/h6EyW+e1KKXw
Dg+sSfxDYTy1Z5kW/BU6AHgZOhtxA7FUcU8QI2E8PlJLWDO1Bnr9MXoRvdhvaos3
yQ3OQG9IWii00ncDAOSMxp05m2r27mbjyfaF+PpJscNv9dYnZ0p/02OU1WnNCEca
R6LuoqI7DNDCnbPlMngnIj/k74hiSmikoa1jZdwm2D1oQpdj7gwxrqBCpOYpGuU5
aQSmMPWmR4phCtreg6NhPWlxi5u70Z7+C6SDCxRpN8GQ7YuT4Z3jKjH3ziCM+jB/
V23qM/HQkPlR/C9p+btHCQpsNgctqWB7J9srEaS0XpeZahLm3m4MP2FzBsNncoUZ
mtlGAnZT75pet5EwZ6dETjJ9tfxETrQl7zZCc13JbdTfk6qxRqQ4+leMjk1QzKFE
JNZxSZGGVJDyBNH13TehTqovZpHWCfGZG0RcP7j0tvBx0nwHODBUpo49Ii4puq43
dEIZ+InTvT47Rg7fHNPsK0nJ7bTKiIAXKI5qh1yR2BG5oSoncZN5o1HjvvxCxG3K
L0vJMz2vBDPnyb+ao/bauj4rKifOlCQQvKyw8S5SWvfrtQPlDUkrjpvFrLAcoSsI
Crw/NwN0zzecB+9O8oQh81PD4NVd0jcytnZuBysEEmSlzP70uWWFV/GqV2kEE5gL
Y1R9M91KO6mFgfbNeDszrvTH+rYVCo6YsQyNQeNedvEyTI1TpdppWd9yupTzuY6Q
Nm01QXjGIIYSuUZwJyS7a+EGhzkpZznmN1TksO7yDXIv2HCKR7YFCmB/LMn5Eke0
324sQk7eLok0TCCruKBWRrw1N4KqIHc6RtKAgYsTK88hdrLxK2i0fUeRXlrOfFAK
hNZHrT8aCFSAg3GbsMzHO/+MbUBuKuDA9nduOGOQUMpQyawV34TOI0OVbh5VTvjv
U13Ojxa/DdhV8WU4jZkNP+etY5lWGDLYtrUWx67+af2cisr0cW+lgb1OlKfwbshh
mNhAsNPANsC6uCFoxm6R/jBZ4I9LXdTbFtTR++AK0RtZI0QGypa3A2LevxmgtQkd
zD5mpFCeY4U0QDav0MN8vCHOIJ2bKLX4kTMUjQksIzwNOeKWHRW6B2pgRxy1gd39
clHAx4H7WwLYy8q/088z2HnA+gB2ggNlc1GoMjVj6DLQo1mHmg8iICZ7VUFAcILj
IIgAQehyRsAbe8fLzWvAZAtVVLakcj2qf6SDfNJZgkGH1bOVGgYGafvcvjThqa/j
t+9pvqVOIXoe+EZju1ebJTI7WIaoUut7Sd/hn4YoTKBSvcTL7YgLLawfsG/EoeGn
dwgB45L3l6ddGnc2HOr6V2MwfNbPqhaBCFLTruYK7zj1qM6SIev/yHHltN1AUB8S
yYkTzO/58GB6ZqIVYTOwBfjXfGFPGEXe/B6eRjfVHX2K6aAdF0bPBQmYeKs59iXv
0oWjhMYzRddu9VTnqU5+H52Ic/HXMx2Cf9n7Ald/HSlvVVkLHkJd/itWkbhglXeI
lpTQoOmB77Hl2e2BVX8ByA0kEP1WCFtD5oO+StB/mbi/ASSEpUcvisrZcfojMhjk
NLwV+T4RIfClj3ti2VVgadAfO6VL9ONNcdOAEvViUZl5+hcDtsX+FLCy096h1JDy
PFHPh86GPcIdJU1rdthiUnCjvZ7xQXXBLtdIr4B52NJmzEon06FokHk38dhYewlh
CTJaTDY5vIP699zH4qDlJMig8b3RlqaKuZlkqduq7NE2gxYJJK9ta4sPm2EubYgu
oL+SMpBouYbhSA1AKC4udybpzfJCFM/5n5vMIhoJTQ/N+cR2LUdpT7qVw3Cp8fCj
TiuUf8wBSYpVeWnzB6eijGUilVmTeYwsoBegPkclC/cnyvAN0WSkZGOVQhAsizkH
UIewIW6NSQW1ac69kfTcyJeHuXuQKf0bE3h+gWyKwG+Z6OLkgXBTWjefa+tUHj25
cllAx+gPZOQWea6MV9BbtpHi9DTSVKiEh1TlNeOmNHU8XTLM1hQe9LXKyHxrM11n
Fs2sQEV6E1WOKdLaMXc2P/MgeXSjItEqFlrljMUkaltSSHsr+HQPZZI+lNX9OG8z
KEafwUJVr5SezkCfRXSvoMvTUn1nCZJskK5jeqrGWPllZsYOgz14CE0koU9bJA1f
pXfSeWJwtC7NL0ergOCYmgtwP/KQrgHG2zqFdP4lqwMUIAJHAqOtcHHHrtVd7kFx
DF/hmhw0WNpothkGWejSMh14Dls/9baifADWHrmBlTaCDwQhXqWixPn3wGh7ad8p
6cplIY/t4DVCKYj0RFHQlooUf4lcPtHxuE3y2uxFX+FpmQEQ7+HKV+tJ0lXQZgYO
cTla7Q0NijuaBId9ToAi5/b88s/NhT+GtzEoMKDBtg28YEQRK+B6stGPW4riXQKx
uSBY61pYFT6g3MJ++Texd10s2Ui0BKR2qxy09LesWZFsbN+zUEYOTgkplE9xGIvV
hTObnKRuuqgMOYz8ArW0npiQ3gNoc017grnF6tMFd2y5D4o/gf0tj2p+HZg84np3
XsA/cmSp9XFwj2LL4RweodRw7jyTR1vXIJV7g/RIH8dkUf2LWLeQsGKo06lbpL5o
erL+I/KkEodL31dPMCHBxCR+JJTENrLekyKcn0evsh8yzk1zD/FmOeEUrrtJS08+
R71bTn1oz/hE8qrGpPmAgZ17pW/06bSdFloMYBXyFaITM6XOoVOJNv+PdVk+jriX
hgR+8FgL/4tlrIvZeTKRSDgkXmfZMrsQRy2Pa5xUVgVez/da0DX/B6lWweI4WOn3
s6/3ktkIbQLn4+D7sKx9iGatLAhJ5UcCvWm/UWHpLjCO3BQhCtTguF+Jbwxhz54c
z5FC+gWY0K+n4JL87AqcuY81wubfagAVj53AbFfLmsBz8Spt3DeY/oixR3t5AVhA
leVGHvzTz9KuUNi8EJIwu0UXKVep47nympXNrW5EAWSQoBLMN+e73me4Qyf0gqa5
zNynr7fDNuzVZg41qpCDxRfqt9ZrA0gHLYZHTOds5ZiDUEr0MYibQDEVqRz27cqn
4jGpmVsUvlaJD6BpgwuwrA1SssAvgtwFhexbuwlHjYiRluDnKw7fnDokeyUdbPcp
eZ9BO2ieD+OTMUHibTF6vF0IbHYC2PFlgEUbwuMt1a07Kbp90PekEYixykkiBv+x
cqMkK7W0di/0h9kDYl8zpAYRDplSNuvM2+x6Y2ScPHWuaGpwo4anFVBmKYKt0EPh
blLoZACt5RX5AmG+LTYeh4xNaxOgkm/I/xZWsW7TUwQYB3e22quuQQCy2weJtaqv
I2LU4lN+rmF/1rrkz94IdhNhQ4RqqlBYM2P+UtdBpzf/iuRrDEeHDAcQtjdfHikR
z6Yge2ygeuPDBbE25nG8iG192AhQYnz3ZM7PWVNCMB5osCFmuJbEGU1TJ0i7qfAH
52shKlPU+vQ43QEaPZMudhllx/5AWmrqpSjOIdeoqk+v1K8zuBjrwHKmZfKO03Wn
Q/4SV521nU4p0uf6Mw22kSDUi+FJ57+U17ii6bo9fJS5wWwbMC36cAuub8X9c+H4
FPLmOINz5Qy5XUDlJR7qdzhB71h7GT/8EIdMhXM7dI9pFqZGnTJCEUqcZ4NgcdqV
JMkMaL0TPBZXwjmulDzXD8EwZ7j4auj5n4zG5gOQUwtzH3BDrTGaKsdLPZaJXnyX
OuLC26FD16rXxBlbV9bkII5ZPCIwaG7H9r4rb11pDgyLw8pyA4Q+ZkoHj2Ls3fOv
0WHl4uR70PuHS9/cQpvFVrB48uHcBbASR5nsmOu3T74KvbVdIpe5x4m9WTkGXT7l
Igu5UAWpPKFR7mHWkH+WibRziZpBXqSOFe5t5tLNG+XJT4aGUGoTHjlGiCJE35M0
zwngilnCn6YkMxkMWOgCTVRvBmSliM9wK1MAEkQgBLL1W1NqfLhNhpB1nCzKZbRg
XFY2e7at8PuIVodKgR9PENXnBaHoe//jbQPjCDIW3loDjTWv1jy2xHZxIuzjUKvM
rMYucjKd12b8K1oI6toZcDKVyauQI+aPCVklA1U7l0r9nAkr3iazJnbdsQsB4FIk
mWRQsO9Jfkei7Fu1jk5cFnAXtts9TJZ0G2I7NRx4FZWCuTHxgYPpMNNJExueHeU+
tvJSkgTJyFkhjZyl5DgkvOrKdj/xPzTi3FamzzuDG08Gtw/e3ns+aGWjkWABAksV
tsBSl252nx0fw6wbV3sAEWsQODE7jrT7HN+Q3zcQRHSZI7zfrirWvslhGm2I8hJy
ZzwHPDIvyvHbb13ny54Ecbq3k9MHwHIFDow1t0N2nexToOWEJvLJvVdxyWWK0czW
O9+K2lH8FlJR2L5eMXSb5khipYUiGYqr44kXHObfJJ+JQtE4XKDqHAhNGJSTr8z0
RkRcS8UBEZ5FZDShxjCFxEAFplwMh9ueBdfrLoSrEWlXPD2NtL43zEoqe5v4oCa9
2jmcPL5FBuwETSz1i3b0FWn4AG68BjmhfxpcDv0099s72yC4vB7UP0ZPWjoU4NvA
p0DBOByihFmhEk+11tVlnuIfw2bjMb4KesAJojjkNgc/SAQVzG2REkcY2pixnSne
qiNPgX3LEnNGznj1cr9igFGPoyyB02DJ9Gy74sGK25Sem+AaLZOGn25RXLaoiE1v
YcKlo3gSYMfKyGpw8ibLvfPVpxWmlAiEVkA3Q7JLgZftqtlrH5y2A5B36gNgBSbx
HhK9BOvyEpcQ/tSTE8rA/Y7NqJ2geMslJ3MBiSeloV0NSuBe1ygv0CFdm0K6uNgq
5/E5VSJKR89tgL+YIgv0XouZaWOGtOMqALmegh4lZ6qtXwIWYH+dpA1EpaPzoEr/
w4EjN/UsX/i3g+Yid4XnPKjgXhTnvRwTQWE9IESZ/jF9X5A+fu1uA3RGiOfeSoYb
Qjq6KSc4GYTkN+dUhnj6/aSSfd3i9xdXhwxk2s1kfl+AJ+iUdD5jCMwpD/ck9d/9
lmCTyjuM2eMClH3RwIjqWq3zhjdi2/tFYKW6Naip/hM3WXr/HFpiVlBPEB2Ns3WR
T0uh1Yg+I7D4a+Jw3z73HfLVPxhRyocOMEC1UMCIS7r05qfIxuqOH3VG0La13+ws
l//tNs1GzHd9xdmGszrMQ7Eh+JVifwXnDtXIe8P6v0Y09CmC3jHEFDGmSBbM6Ubz
xTUPrgnQ24UXENG9SyOwXPjId+tRVLPDy6ZXUsMcy5g9kS3CUbv5Z9Z3WeS1f3f8
PqpyYAkCa0qXffavZ3ODCvgWBPXOiA5K158ynhMLXPJj/MOIKLfHmJnCNed+kPUD
gYuSyLhYHjkJ/Qzs8v1DGOe1bUVUGtu23sFPef+hIiFXqjP7i6IQrRsd8qez7Bas
jyitbMHBxMVuROI3KKCgfS8HD/2HPXfRwQpvSuFF4WSMLj5JSv96UQjFDfgPHL2/
E5adVS2y3r0tfcmlM7rIo83QqS3EDk7Vwv6RnbsshktW4Kz/3WQsUMp5kIcIA4dG
b/9CzdOwyQ4tGQdKrjpgMN/SfxPbKjblDyGTbvsxr4yFV2RJ2KpU8P8EA+ZvGUug
IhWHyjqwAWDpl4qa1cjuFlm4t8bnHznt7Y72Lpbmj1n52EkUBC1VznCgBHG/XKES
OM2cvEdXN5etpDpt0tfwkTF1uDk7ioOj/I0E5V0UynHJJCErpC6tBy3YX9uGRxPR
4fIF/hlWfrxmrCS0av9nKgN89CiDCcqwd1+4ArSwDvp0BxDDK+wDQfsvVjMSwVRN
e1BqMFcrEWZVuYWTstNXcrQ/L/Py7UT3R/B7dBsJQ/dpbB0+B37N09RYZUXpdmzb
w+OOosPTIsDsMtz1CnwuDZNrhRWXkcwZktSdcW1rnuhGowIq9tgRJJ8at9Rtm+Ch
Fe8vMrFl04TeilruzmkAgmr/OF4naF49GwLA60K8alXor4CudhcYWygDMSvJbSLA
1YpWqRXCMeCuC5+9sxgTOWmAQ3y/FyszJvz1tZ7o2q7CPvE/W8vX44oSh2FjJOtq
HTo86uHUJq5PSoQ+mfN9OYJ1F6U0ZAbTQLbuW846iEWre61jUfEwmC+fs7ckAztx
VH6YEKNHCrii5YZdzCsRagFJWsCWb7+3AN/go6yCn+n7CwOUG84tlY5qjbF+bd+/
qz4lzSGyIZVyJKwvVhbzkp8JgjKZ0Rli++Ag34a/MtwitHH5lHBPvkO2jIXGnYIY
QFR4OtVAzfSG3vLg/GmqkZfGsvGwbZWHC6vQ5C3VYZxLimtros2D9fwsa/hRSZJG
tTnRRM//ddq4qPssc+82HDQOLvcADZiCWhBQ6yDjOogwui9s0tEJzGtCBh4qlVDi
UAw8SsDOKxDUG5HD+h1G9AF3VQgAbB+Vnn4OvGJQmIbGJaIDN1Jzo4u5k1jcWtij
zO4MdM6ntVoBT9+N8Trop8p2R08VJ7uEu7sjFAXitosiKsIYEaEJlD3kEDygXLFs
wIYFm1NRDCz8ybHr0Hnu+m8s2RZWQFwEceLaa6PRsELqggVdptbdIY8sLymGZG1C
wlpm3LkqBKoRJwCwIm2PAzwQA/+Qxqh7Yjcjr74F5+acxkcldRPjY/kviohuaUYZ
GrJ8nb3vBRdhCQtzvXhkTfGoH11MpWzX5L+18AHLgwEWwFsUb6ADPW0xFl2908Gj
AAo3MGi3mstoARkxIu3kJZWvO1zw2d8+vKSEyzrti2zyaPmCHVpjof1VqfHn4L0v
0eerv941gTbCMwuBYk6k4gbBGARXr3du4lEL2wppQq4OiKLL9N3q67ZHDEOBfWRX
yWU8D/47VXM3MT7YcUfvnSymHSGAMeNgxkrP1h2Lin51+0Oh1VBG8MWlGmvXjYvB
ve5i7BfNUcyx7GS4S5WY4Ces5C1Dj3hU+RsxqMYSDDXXUboJGOqIYWf5EX5WAxhb
9I6HEPZJDF/Clcyv1IuCBiX493OmD/es96hw+Swjmh2ZGVqHTpzKMp/3Ek/tQ6c0
glRF9Bl8zwAD/RiXfVyXJinyzPS6W4oT5taykqc1zZ7q8/Xja2XjrjXEl/nEdnK6
Jv76pL2LzYbkaV/Ho4LKFmNS7iG11DpqFkRC5kc2fVXOuFyGT3LBxZXCT/VWKuqL
jpA/H0hq3d8bADoONfN9blIAq/p7z2f6fpgTCqTjytoWbsqSDxb+D0iKt0wlpExa
sNKegu2efHfxVl7NHt9PibDF2r6UIYYYD9XLSP/A7EpWy28rAQuLkfCB7veGy7Pw
KVClU4i8AxoxAX+OoCGHB339l9Eey1+myNGaE1kdwrKF73ACcE9qZkxlWKK0A/84
GQk7tpTd2BKTo+Ey9z2l84CqgODOh7OZ8OselOL1e6GdItBybwvxGQ+Ke+dP66Fh
eaHjGZmFKATpbhG5TzfvBeQ8bZfv8FTov7wPDnATlt4vgPL0lGHUXDpnRiVY692/
/bpLvxiHKQUe21B1bfbIsstsujquucYB0Hi3aru27lq2H1MoRuQ2sPcM17WNk7xm
DDKDIdetwDeHpmcnNm5+bK9pb3ne076bNQOi5yH+0shPdeOCGH/frQG0dBBsSuSX
dsm0YRU2ga9co8UYFb4sN8FuiU+5thqIQNb/8QIugzMzrHvDF+KVMOuwlBMI2gep
gdiFSUI8y0VvjlUW2bGF8/6/JHG3O6of1sGHKUAw7tSM/NXmHs9YGNWtNRMtESSN
j0ydCVEnl+RuxTe4mSQ7PKAeot1Nm3IkIQjlrf2gSF0RK+2iut1fU3yyj0hvrUW4
oTNxHVBDmU47jYeHGuhVP/DfIK3ixSJiXcaxFGj1407lHV0XX/D1J5i6cMSjP7Ly
c/eCCmPBmM71XFW/1B1c2qcntEVVa789O3PgHxx2qbJzXktdECQWpAEw6/iiYdSp
Zct38r4UB/NqwhZl5NX2X9gXG4flhX27tNc8Wnml5MytPs1Hp1Ft/PpmOklh1ics
p8BhNlLSAg/pcmohuDCNMZTv9Uf0r8vAwx3/zbOuOrOwK6vftfuV7s/PqXIZO+UI
6kwEt9SBeMefYmcji/L+VrLBudgfySxUFOIAs/zZrNeE6wvwzMwMLURaxvoi5lll
uJ0ZTUIHCpA1rjHVU2D1n9bmPLxztIrbXMSpOQ0n+i/bEFlGTBO5d3EL/682tz/7
U89sCT5/FEOQHoA/kvlopVN9BDGDJp5JDlbVvpcZ8juU1JgrZBeedZTSe5tP+Wi3
xGw4UYpQePjG0cblbqLeoYs2efrQMMXUbPH1JJGD6ZW7muEzzZdtvHQZRhqUt6py
svDUJPA2SOMGdmtJUEaHQPgjGGIZKcrIHPIvr4TMljpO3E4UYZTp5huDWmt+8cgf
X4BBL7SteBahw1zKSEids2vbcB67QsFoCiYjamv4/0+h6hGdnb+duADs+FCj79J1
zUQD5Zw+37l37nrBE8sBY9/94DzmtcW5OuPjZvV1uC+805Kklcb7nvJxUbUz6xOA
akRNAKn4MhMWrxvrJvs47iPpl5X/+vPcR2Ya2GDfMK8uqQA6HEb7HL0aUJ5YrdWU
A+WPuYoYlFmGraEJmeSdgtMaIZBRfP0Z3zgjXE6aaj12EKOqDyiZR19WoT1JBj6q
S79gXxzg26te+9hhxI+qz/SXtC0M/GsToa/rQMJ9/qlSXpXSAJ06StNt1ReUw8rq
S2DbfJIJEdf2oSUea3grm3vMAZ5DwuxBusB06//wWvZKM5qiDyDkSJ0DJYEAleZs
PKDwbNJpijHBj02NP1RAhpNaH9dgSFbM3MXABlNiMu2PGCyWFi+UnKY6g0O97ZiH
aLlQ1PzeFZE/19QVuoR1hi0HofEs3Zbz4OljzGyhPjOpgApSuSLZOnA98MogCzHt
TnRU7UAmsxpB956MRMROn26eK60SQdqDqloXueU8JuA1roq1A+3Aph3jz60XNSwx
UBxbsJW6EUhmvkFTBMoPvYMfhJvRXcTynfKgo077fyCPwR1Bfm2HHEGQhnMrWmkP
kJtsz17vygt9iGuHrosuzJJDQj77dQphqVRyivHx32PmNmUWuDVLOeB4cN/CjK3Q
ahHSa32Qv9AkUUunuWSr3evGnO0kGgA/ZRqAfpNigHGViAwOp6pMUd1wmJMmcjT6
zbaBm7HGLJFk/UdoR6svkcxBezO8J83AnFW5d7Wzu+JinNxFslWFQrBVpYMR8c/b
WZJTGGQ+vN6yiKJ77QcaWWC1sPPEdHWDBBdszvPZ65YbfA/ZzdN7U4grOb6kMdLU
qGdF9l7p1sWHkWK3Eaqs8ThZH0WiCRWdBc1OMSRqEvCYhKG8K11A5r3q9S4ee2WD
NuVSb9nLVr3E8/5iAoNuQzM1++5TiJoOcvcnA++JJSlwqJTGjuPK23l51+OJgdOW
jgNAgNVP2qiX8ZP0TEpZ8u2koVR0m+Zm1FUBAuZmVU2UKZ2LLlo4gWs60tGid/ls
tSlINH3N5+e8igsVMB2+yLSQTuDFlpGDXtCmaYY6/034pMvwDMJqL1XleTB/1tCQ
dMzLQKubc5Aco8gWL/XgCpINpVVzjOk8iQIQEw4OA6m0EGNn/l2JenipwmnNdux2
hFahHYtaB8He38hLTGu2BSmK2JljNoawbjRXOCqu0eYtR6hYjQcv+jz8pXZSAEMr
w7eFKrgMtQfEA8cMNjXJy2NEKtZzgc5PSMlb2atQj/7dSr9E2xJHIiz1MB9U5H4Y
4KsCXeSuASjE0bUG9xIs+d586D5fJ9UfZAnjHM4I73nak7QMT/tMoDW+xb8r3Yzj
1MxXsGr0i4bWlVW5PrvvQVlC+/tn9cTXAX9StKJf1rfs3+PD3KVa0R7uvpBBZIhm
YLp+xA6wrj5T8bdFpa1x8zNwtTzpf9kK4i3J2Q37mB4Rn0K8DrjAzcwPD5ruOVJB
faIxPQArkyyJmPhObFtwnbXqsrLvIJwAvk5xRVAo+mQwVlSSn53XmB8Rs/0WUw68
Icv2c0Y4mr3y6+eIIrHAdtnPvxCICH8ur0NrFc9uK/W2kSiqZP4452onzWlLlm4v
YYogW3JY7l3t5suEsFOrqLfEZfXGuFov6LdRx2XSPcX2IUEVW9JtS+liwpln+wSk
J4P8bIzXWlAZzbw5b5xRaI/4NKtpI33lo7aUppbtVaQ3KMJkI0pLFtDT6q+F4Tuz
zKXiPQrew9ryaOLrBKcW/LZFbRjNC0XbXGQzdQpLxkHPEJXsVPpXkgZYTv9N8Ete
ApQ1klbZJ77EQvvQEu96SnhQZk1NY6dxSE/s6SGQWbHRgVzYy5/FtQGsHDU41VQs
0LOOKxHhd5kFGs+Y89u278/IrpdJGeIA2hYK5Qd7PP7xyOW4mvjvTEtPkcIwLv5W
rNTvvtCl7vnXX/EOs0JR2G+gi8DuTBe1qOcz1/YJOqvDodgPV2J91zIsg225NKnM
6E/jIaIVR+38TFDx+M5tMrr8dwRcghxKwm5ho5psXkclG5AgzBAWM9CQ3zg7Zxgq
OkahQXmw/wy7FdW6ElmZwmL9cPenDnunWMNnKXaFJ262ABse+J5zoGWcpwqNnsyR
xc3W92xXDYp4A6KYhgOE3jOSgz08g8UI1maDSXvpidcAt3JA2BiEw4Fivm6Y12Y8
khZVYVYOwZeqCqcWtdLdBdhuVT/Q3uuzmRB2weDBfolvbibljaNftcCKs/buRGsA
JtBGncyj3+Sbf2/a4hOKm3aTJ7nJrSvvZv2n9r7B9lKhn8crU5J+GB3qCUXkd/U5
2u7PfgY63yqbQdDj9dXp17eZN3h5iz7ryJ5ScUsU0o0oiwgI9znogtaFC4ko0Tra
VZ8TP3WFdtZ4bXWJMeko6jJ3rnh7D+jrdes5bp01WzYVaLr9v9vf4STscciZMsE3
cdnlT8KgcM4c6jbhlOm01hqzuJ9xzvo4tyzAuTKKRKkxO+MvywnybsM+EZoe9wVJ
LGGJ+NrPBROzjukl72Yd5uhT/HJW+Xj4VMv1c4GOGEZPlFV74ewwT+xycWFFI5ka
2BJksbgs4FYTLewKKBHZMi51js8fWWA3GuLiaeAlCvF0z03MOFqm+ghPfLzGL+Ij
md4TPTLlTZi4o1Syg88gKtgcsn3Zf2Suk+gv9LZNI18+TRkg2AESD2RKLgdGvyxU
c6avSZTJtYX1LGNjbiukxkgjixlnBQx8N08WqOHa4hnMtAGt7iKCJniK5gCOdC+U
Z7fxwrHqVV1TmRkr4U8YK8etpP91Xdc2FHIneBg7d+fusQRRnT2LP0lIrsRQY34O
qWWBt2vrbllzDvfn646oED0IQwIlnkUBABE8xwcGtiA10iLYkigvIyilgjY1DBTW
ac/4dMqFDmsHo3dUVqa/pgcnN56C2bRAnJP5UwlsBVxDfVtnB1zh2ORebvRwsPPa
TdhhC8Bx7UBSgrDXL8TZYOE3e3tq1mgNQnLU3gMQgx6XxhdJ055LbODSIvLimwX0
LZKnKfPGNjWGmP73fScVFFVLJfsvLuB/AJWT52D8BUivw6uJJGDiQ6/OG7Qju3lY
lChf34Gcfr36+HpJ4sj58zv3gKvY/e54onkq4b6gMfiwEZf7Clg1KKRNl9plw9IP
/tXR4ltId4Ug4F4MzYTboDrpZZbvFl3ySsSjeTQG8qoybQqUsrmTtpd1FzgqTj+P
bcXQ02T20wAZjyJfhUhN9aUgNXyG/ghpP8OwJCpbCAI0FdLIBpP/F60X7fJ1/+qi
pb/5bsw9OKSJhneAA/kQ/ujzqB9y6qFYhnXqjKu7aSlRWR2yRijt4HfxOz/ny5Pb
uDfDKZu2ccQb9KjIDcFOnS2FMPpMhV5cQ8xxve+WD3YZkssEnPLZTLckoZIe9D1z
WT6TVkbOiY00tGE3SGbCc8UWf1QIrsD7WYZK0SRi9DhBHErNIFyhkI9cV3kqLKKF
LtIpA9E+YyvB8pVtAnO11b8Lt1DhIzrwfS+/9YyRo5mZozmGk9XuskdOgNaqwV2s
t42QkNlQROGDGeZU1oBpsy5AlqQ3ptiS7ratXZtNDIsqrenudkL3RlctxJBfw7tb
tX+U13LWsXX20T4xW7I1wJoqh+LUq9ulgGhSLyBn4Yyh0Ti7jky72dY0vgxJMgEA
T+weC1VWefhwh9VS6g1mEmmRzUxNeyU5K8x8mhFU2NxLCXbofmbdUvt6+lrONglU
kofDHihdMTyTrcRDwp1BM5Idd3N/UgPeHEH40d1HVvwJO9yuAqsB+nNzFMgcQqO9
tqWpDsLjCe+te5z8SjjR6lClX7lXsuR2ZpE5GjVNDbixPR6bOKEz0e4xingrR/HD
wKMhYzXaQ8ANlqQfljLHo+8+F47ZdUHzCZliuEexsiv0FsV4dtA2yh87zmuTr1Q7
/GuynhVk+EHbLQ+LEOMTE8g9RFIDQjUAHC8LA71JxRgvPiZwMDHQz8C8xC/sYdTG
U3nq3ZsYZF7jhMg3Vv93HR3cDKGb3nIRio/lJZG59Bi5FCYp8lx5WdnE64krG2EL
wCXXXSSE/WyUSns4KqhQ1m6jkvCuM4ft92Yse8HnOlakOiFvZp6UYLe/DUyhviHX
9HdcKwUJ91TWWyVCqe9hbQwPh+xgUc2VeOtK1eHYdYSFEpgrxJG8RRPVOVuuRJGj
i1X+6JoGd2/zEm+w4XlbOaOZqlCcXmZhpik76KHU2V9zv2L+E6e7Zkl5Tg8jNfYW
UgZxYezYKDiDKpmHNN33gqIpccC3oItY9vJT9Z4CFiVHc1gIDyHfCvthHn9to5Cb
23kGhnyguIsv0r51sBg7difBdT44IUY46ZMKCaXWj+xzBz99AfMmryC6JINX67s8
o0xFZbqqFPpg222lLFCppnZLSylXQ+dKx4eUrqzpBLtEhZQdTNEBdVtLmQHEd+fl
UXZZXdiTINauD11DTdYTCgOAUO2wkKhxT89OACXp4LIg8Ghmim73q3ZiSeEiEI5i
Z+wkwh3ibgsX6tp9q3WfojpgbA3y1ZuDr9WJbNp2D+KDIiwPeWZV7KSWRg8m5F4J
baSmaf65DzUOvGJquK/KP2WwWpD4zXbW4So4GwXtpivSVgGDM/U4X4WqH9HPqVXW
32vVeMdTnk5/BSZlb29xEAra7nwMYxpVy9oJF4+qCFUIKTuqKNmw/tkLsQyKNfic
bIjNjGPdD/O4k3OQncTGljHdYHxPM9wNiMQ4RZBL0NCxobp5zC3Gr6X5+T6U4FZf
/Rmw1zX/8bthKE6+MiWbbigY7k3RtLh0LdSX+vXIZQaWBLfkUFq3Xrl8/4MnqvCA
Uzs9ikqCX9z9Ug9ug5Oqya/bFN1gdM/GKY2F2QgiIybAOgBRarBDEXOb4gwOb7dO
Nrw6Pyw6ocQNvs8lpaNLFkZnwgtpLaaRXJ3+hJDKjBYqzImZDVTIYBAQsPo6Rhi8
XbxVgURvPVJsEXtkopc01Rkuk5ZS+cp12oZIuTcnF8+sCawfO0m4C9PPAtKitalf
D0nmqCy4zbrvTD5tGia2Qcslv7VFIYaNfi49lv/JtWyhmAKoOOl/RYXf50cBuuhE
aPDQqaI/GbV0GL863om2tYaZgYK2W/v2bWporVfiVi05IQBVlCCcsRc4EbQLQVCb
Kv9uLAVKIfyksOfj3vFEAjnn0MlkyofLrSZ3qxwX5zzDIOg5UrfSV6IHZeYlLsVd
H8EGJz8+euT0a6HDeOGNyruUtQ5OnJETjvNVvoiz0+SORUABpFx8Lf5go2jcFM8W
rcEEDDyQAmpJTYXuMhECOykk99ecBTG3U2uAm9BcEPPQB/Ng/ZNcHrrHn0WWmn/3
O9e8w8LumFtF9YmNCNaN9e90Nz61WRiv6wt/0Rj2CcK/bS68A8BnBPm0imFzYguQ
kqYx6dbsz/+FtlQinOS8JNPcr1iDTQW78Ba2PfD7DmC0uEEvFMG2g8HQauF2UiZ5
dY2cxuJzwe3+ZdLX/ZBflqcmEORwpvkdmUxoekkJOFXv3EnNdyqRPDcCVRHC64pC
yRxgR1BjkO9GF4YwzIBFQMHssaPi68E9t+CxwkeI1tECahWhBR0MddRCMyyi8dyz
4IX0NRt7F3Gh/0EmPoy350ku2iSxQymIPbciKl0zgOcljdKuFgC6RZ1Ag3ZXcFnV
G0KnKnWjaaLyp1nYw6/VD4e3fI/4VRRMKapotmc8e83QbV2dbLI046xTDquWDhIC
r3PUyxUi22h6+OqhuPCppA6WOLXUtiz2cyNrm9J+aSFsnUFloWu7nP1W22uIgj4u
v+daMjJ9pCpW0tQSYTtOz13W5Zzv83xXbDD1BYzSvwOkCOA+y3zGab4oAnG76LSg
lJ7xYcmP/OLdqlhsCdg0s7m5OXe35mQ42rx3wM92W75uIhTY3S/ncvVZYijIC6ap
S1SoKQjj+VsfL21PLSck6apn7IyEvh/h2wsh4NeW7ZZ/01epJ6369CSS4/crwW0N
ORE1zxhsaoShtX4Bm7lflVuTvosY7al+Tn57ZCmlzfAi3kxqvkT2QddL3JK5FQON
XxM9/GzZij6glbMutCJN5rRJxbEsOEsnKsUbWPUMeZ2VPa2Iqa0a2Bh6nJeokMxc
+8NNhB9BJvrWjXAtc04iMNow+83+8NnjF0WenFjGZPHMDAls0RcETNgZLq2wdt64
ud9S5TaZVIza3tYUhWU/zdVbB5g+yxcHToi1vh83sz2Sag+Krnu2sVz0pZe0LmdR
CZ0nThpM5OmyXNpRbrcu5O5/ln3YXpOF7vyW52YLECw5807UQLo6gR11ce6rJU4Q
fXGeaReuUXFC9mYFC7Fqn41huP5cW1f6A40R71hh8prsDeNFxD18U2jN/AeLBqUj
YByt3+48NvFtRjwylm44DPOzkg68gJosC/EtwR/nsjDReAiTCZk4nhsL5uOAkXXz
FyG81i8XglVHPsoik8Wr/JTNqLFxmxgZJsduGjN+WZn4bsTREnVLollvu+fi31Ml
FXR8LG1ubR5xufl1VDicY/3mfc9snkWF0CQHjvv1f54ylzRvq4hw/bpty10NzQ8m
cQd69C2c431sfDZdON+dcN80sINQnejU0D91N2931c+RbKi3dlutfoK4bPTMVDbg
F0LGUtOvoVRymQjawsdGFaPl5lBF2dgU1TliXYbIucNMfbkUi34JOG8JdlC+9HPW
clpd2GXJr3e0Y/vLx6gX9KfQJm+5FwwcPrAdJEjz2LlxUg4sx2bOL0sF4OQM3TUo
VjCAlk82w0FZu4DpR+//ealBH2RxAGU2ds1R1L0jCz5lbEMkB55orFpcmze4kn9D
uuOB0pMjoCxuVnaiBEhxQpUlmKoR/RBYJvnyXxa111MDyv+ah4+bAhxm9hos+JvD
L6U8Iw4anfo8tgflhPeeqtqLrS1w0wrRv8K6XABrwhdwBJwRmecgJFpcDPtsHx1A
T9QKnrI4wv76C23Bbz5Yi8obCU0danA2aQRpQa7F3aXKq+SkXl7ocgGJdoS0Vp6s
d/Q+YeIeivt/wmDY0dRnFXrP4aU9U8kk8XYS3EhfSGqAtTd3FuvNjL4pMkUTRkXq
rjXppGd9rynEzKntLOUkfRQWEcMXD6flBOsFTsr7e4MLlbjxQKKsvNLLDjJy+UE8
prkVC1tA3f9XFSSDZoLH8Y3VMOxwsLH8/KgcHc5hEOKae5q0+ocpJAClwj/FSmJR
5ydeJ3GBViJ66RTG3wtr/52gcRvEfanGvp1x710cJ8IHPnxRIrtIEhcf9PJD+8vL
Z6yEiuVh0YaXwmdjMrhWfIC1SUpJw4eM+BxLl1zk8cnyzBuAL8wOwkwLryNWjOt7
WwHUBIDdP4i/2sQQqcom80cCUxKntvoqwJ2j3TxMJtuA2e/4GA9GQ7EZ7zjCUD1f
K6CTKx6mhzfOieU0KXKk2T1N6iVaP0yf09jbBJxg+QZdlO1mM/93r0PPvfXKMXQb
gwToabmSo6xqxB9hRRp9iZbzLp0h6e/FDGC290nBVLS1USq1gpnE9PfeBdcD8Mpu
r5yiLo023uDfrhVphpevarG7OJ/cQ1fOaB7gdKeZVTp+hSle776P30MlPJoy85PX
vO+EjjOPvruq2yDIJrXQxvLpBnteHryU+H4kSWBjx73p2dwzfSA7P4ZFJCWtFC+4
2VjvNm5s2VKgAwZc7LgqjKM8szOKMFYEXoV8mlzhl74vQxxWH1HooYqh2jl2Rhm5
s4sBTTVJjdeqhY67pqhJETOmUAWBVVv0vpiShXnW/pmoUPp0P9jKk2T5ZslCWE9l
fuJ7m7hGyGk6s7XhH9ExkzoTRHO6IQJgV4UQpyADYEkLyasZLSQpsShqIkPM1UAG
L9pPSsYwnrMYbtzQ7ZExLEGemi4jLe1ApX6j9ppLkLJVan455JkesAQCzthRvPzg
Yf35VdHCKpEATTcbwjHbQf1KBH6zKdcdKiyZdKo5trQ15Cn+dG7pSExrzTRDjUdJ
x0CWKLViAjQR3+yO8OHbYSyvLutcGdFZ7b7IlwQIx5vas9kMsPisJZiVK/9v+kd1
dKCcGFPSsobzYD8ueYrUoFBcSU6y7847nuMQv2PEa8ypAJAhvhwIuUxv2aGyYe6h
xq6RbbY2pFIjK7lOsWFq6+Nk9Hk4wBju4Y7IkkryHUAayCT40yY0wwURTG2Fb4J8
byMOVSKWB9miZahFHn8pLs+nu0TS/tgf4lF114iTFuh6154bF6HMbWX04W5pWGY3
4yPA/OF93DgxF+le6ux7Z6GRQPXgQwcwBlp7OX8S6rJossH3LjckCpy5OZEMT920
7qeB+yK3znMn/uosajzJjUzeBCu3IFw8oE2w3ff7qfz84f3o12HJitl79PS6fRrs
5T5AFNRzPxY7mRINdxo80xiDUYsTdOEcBSzVsMaAqd3T2lrItXVjHCxFCjlvQotY
yvL32UTb7tiyxeuKi+WNeXtDNFkO9zq9XJSz50nEFEmbaVh3rWc83fJfyiq75yPZ
Q0okLJHMSds29LqkZKtm1Q/lGn1Ar/QZGsccL+RLlUGd7k7fJJyufITcJY9ZI4pO
siBB+EB42T4wl+Z322zMLHdGtHesKryxGlifJ0T1msfvSRNuf0gXyD9pjunw/Iy7
xM9T84MVTpG8PmUNSZ7k5DrRLm3iEpRnGLydPe3csTN125qdJ2+wPI0R2jMGuWkV
q+arkisBwR9ffLlf6ituY+tehUm3ocU8r0AV8bbcvxvYI7AVYgl0Imz73KnevjVl
6jFzDA4O59ZpGTxoE6fAOQxsr81fjPof9S6r2PcaKSXPS2y6Vr1gWafE0DuRNH+W
OgCLtNhFS4ferQa4pRMOWZwbS1jKXu5RevDOBb1WCggSgry3La7/bK6UE12RNAFe
Uz2rLjLsdNGPXPZrzLTPizdt7fl2VCIK3LTh10FemvlFpYUQo/FHiT4XWQx+xK3C
rrVHhLPHYfQ21+RpthGOONoIK7572G+u3hrbhDzcA00yJF3udGSQqcsOwU0/ayD4
rGgYb3yb6EIBU+aZLwsdLSGWWn0ZbYjiSsJ5ob5AUIlKV2z6HzBWKhWD3PZO/fR0
UCFN5y4kmN1tsQWTrzobhtdZNOUjjs0lMB+OT9gbgcWFhxSbZ2qV/WlM9gyT9C7H
GTca0xs+PEh43Lnc4ekbGa+06DHfOLlaPUlRBbcpP8r3zuK/DG884/hfbW934NjT
3YxFXCtoKBbusLCRW4pfBnFL5dxjtLjI4GzpT0SoE+E/1SytnfrDZjX/JVYBITOQ
ygiIIjQ2f3HsYH0zZ8w0quawELAwu/VaXtz74ZAmwoLlf1r6n+jURl3v3hZr87uy
43AioIG/1xVRROGFaAuM50mqJYoO8lJdt1pbUFl2iWUN+9vgq9VU4QCNQNk7UytN
uJNfpkQVSO4m6xl0Wuc6546NUJxXcg5FsUHDprDEQR5EnPdu8cP0ur1jw2Ggs1PI
4fWiMlxDvms/j0eUvjd5HTMkO1wDiJyF0P/pL5SWSQe8SO8ivF728UvdDJPwOKKz
x1bTKS0+/N43m872X0fQkl7Ja6Lnv/exkKrnKPlz+OAZ14meKyXxodVlRuYB7Jui
sJx5zErKJfEdpM/l7EOv2xr68nyVcvuQxlUu8Ogv7lIGHVNFnrtmFM6aAhQTJhep
Xn6wJLhG6wck2uVuAy5vA5H1W/XrLOMLl6cVyHk4Mf3wXfaJPLeLMQBLPBFp8EP0
4aT5C7/AyyiaWjE837nhie3m+FzKVllURKy9AN+F8hDn52H+uad+d+GcRzwgGZZI
6V7e9kkatpY1j0hEElQ800mc1p9yuea9JYQF0iOcQXIfHniYTcQvQTcOCkvRS3lS
R0Pfm83UhMGvMr/8daJ8XYisetNRnlqOUSeTCLHu/chWrl8+Oh7G8x8hp03vrGd4
kPANJjlkUiiu/z6EuQxP5JOkz54WSm8n9IgHQ0OJ79YS2TqU7wVgO6w+opcm+fd9
jXox0pNDhOr4BJAHopyd7QxNhH++xC6VSEmCqlPQZcahmXuYx1niGgZqdWb3+JCL
/XKFonaKnpQdmgWcKoU7HdaTsaF7W7cH14z1kp72KiUSAPNmMt+4suRyA8gtRBfm
KmgBjwXX2nyWbt6B9ZhLe4ZGyNWZN8gBF/ZcelHNPb42UAenCLEqH/FC3OeRRPAY
qJYwo5UXfh3a9Xpv2mIXBRe1whWch602h6SXztk04NbKds7Ols+8eIE+NUopQudt
zm4VEVv6olzZPksqre8vVk4Gy0Hu2/igLq+Qv8UKrbSPp6ldWsNOcDIia0taUWfB
ph+MoZDPhK/j9nCmhRNfxohN/tplFk8or+OeeIwD3Str5YWp3naniuhTFyuXpAsz
2EsvF9ru08Hm68YY5t0VWW29uTLU4cwsUQY0qvbn5W/q9xgTHqSeFv09q2KypkiC
Pb5/R2ywSs8dchAuIwQ6HODryj7ZKIKrp94YhghWd2B/puqHAZmkh/2NDB2lMI+0
zHMysAKBoPJMBFG4G1BWdcJD5ThoNrENlX+wbhOzlU0RkCJt4c21PaPXRWiMoWWG
0WDK7PzjmF1SBPKV72dcIRYbJHzh0ywEpQgN9HtufhvOkNxY0EhC/L30stuSdiK+
qUKPYi62PGUryT+tn61AOfk0bOVdz9cOlB2XhSh9CWGzXIVYlfODjf7cWaqWRRPy
+k+kq6Pc+1dv09V29Gy1SiEW7xq7M5Ev/QzW7WewMHd1T9jNgrCudwurWuC8vyc5
mMbJx3uWDywkvm7KsFyswRlIBepurV/TiqHgcr/w/+FXA1aVAZIf52lVuvG84GyM
2mc98Ke/RL4Rje/OLXh9ACfg4q1v0cQThZwIc7LrJNL+B827X5v1qC9QpgrXJhIV
q8hB3TMOsj1/2Rol9UbflJTbV55leuQVlnMVwVBBHP3GBMlGypXD1Of7Lu9fyCC0
oR2+RKhaHnfhcmYXy71690COA8MTnbUwEevZfoMskcfnWL4wbXHuJqVcfLcelMW5
6DtgywpHXf5wlSgMGxGrbNpNZkH0G7Acnbe5hszOIgnEfd4Mgkg+T1w6PZj4eNpf
0EmXnGgINZhk2PGryJsQ+iZ/QlZrh3YojcFqoXVFxSMjgOskJNQ21eQcOk/RKacK
QJkOIPTfVbrKm9YXYFL5QkQ7s/d6n7rgtKMWWNJ53Ye6WRGrd6/+yWRYumffGKOt
p4QEGES4lB+bnGhymgdt5SSGVM5t18p6ROD2q1hmbWJMIsc1Nb7X2tj6aA+U6iEx
ndxMW8bXAmZpgRUyKxxxw/mQTr+oop8U5X/QAHY5dWLV3VW11zMLOXXnVXlbizkg
PpFVERjAKxXuc7bHXjXPfU9BmUj2RqKWNFd67PdB4GS+3LsmTi3RqglzZabZ8ood
b+SeG6n0dbbddHpLqwZo4iVtoFqsqnEotVwZftk6w8OrblJcWYxVkctQE23pqnf5
GX/hJ2vsVeXIMMVEluPo2qWWgxVjKOuR6U6n9DVtLYjotpchmsYqZJ66GOxg1GEP
8eZwDhWtoEm7GBEe2g9jA5PA0uIBroTuFKNlPi0cSOcw1k4PWwrb+TeKI4IcPALY
A4TK6OBbl8drEtKSzAroDMBfWGitrd9qbbW+PbZEwj2DamWF9l2UMQdGmpCkwVS1
MmMnmWa1C+qtAX5AznfQM7dZy4YDuX3ri7wpZ5tm/jOpFt+r1hkoJmBaImuJMY1h
p+Il8ffkfmgNJN0//C6mN9g+DMxnmsf/Fi5itKt68bu9ZhiIOdLQmROpHmeHr2Zr
7Ggjn08g9n+LFUf4G1LtEafXwS/KyXIn4qWdu/sMFT3sOHLWq93287UNoU/7jNhm
8jOboGV0kvXdyiG+gPHHdJ8GBVDvdtffb1Tl9pp7iw+fTB9oKXJThtHJyzM6+Ohj
9yo3yfUy4mzaEO1wb2RDedwlULQzZHHrUiReX6g/l5ajYN7IRl7/o/L9cUC6soCf
y/kBbQBV7KTetRSZYISBHSN1EgOeuIsMk+PwEu8TEyb/SmaAUev3IRHuhSVNpcK2
Nm1h/w+R0jEN7Df/9ORqULmPHNPXqXxUTki2OTAfVLm9ZtJm5Bnw2h98UFxqr+Qx
y5Ojn3lsfUDqPJGcss6wmP1M+DPAyi++hOC6R+aD+69Pjhba5PpiLH7O2nGImW5+
D9M4Z630VoNDmtK/7QDs+MZXP4D142WALTh3vRM/FS7O/Q7DdNABAAPpsLcN0LLf
NnYDkXuKWNUeCzprPm/akDPWNQPCbqPU7LO7eol8s/laXY/ZBWPXYRkwTzTjt9eP
YKXbX8o8vX3JzKtEUOY4Qh0MiIg/zp0T9LPJyG+q+UFClAm+86o6FUr4/5dYKGDY
dEiI79XX3be9RUM/febUWh9SRQQOp710Bs4bQOfVLr0ll9diKC9dTZCtgaKEfYYK
ZiEPkP83VRI8l69hThaiz9B+v945lqCADo1RWRaPdmGkFkXT5r6ry9acP3gGDdk8
feMnS5Q0UlT1Ah+bBoCxKEaG5fwgheCu2OaYNGdbAZsFxnSLVHW7FneLRFjadRyw
3weuO9ppvuCP5mZgIAbKfZKV0hFxVq0kWf5JkK2OHwmJPgwAjz8wrc+YDtwno8nI
5l8m5dU9gCiT4rUSgYaNbDv2uzYA0LpXJs5JGUCq8a4Dayo4dY0yE+YnIMiJ6Gzs
KDC+qS7TMN80eyLX0lrEvV7ZE1mQzR35kR/mROYv5ObiRcRWKIQAZZqp9HMGvuL8
CK+31Et1bV77hYB3vHKmK8audJN3YF8CCxJu0TPkuPD4zYtXxBW0/ARPYZrmFhiM
reehT2jvffqZxEkCpl+MH5JAxH9FYfFi2ASu0TjCdFG0XNr1x9bwGFdM3GYXCIhn
P6QX+Z2uJ6vH80XtAwxjn6ZMK+mDoRakipes1E7tEnsV8zwqSGhb1kZmD9RLzdfY
ifhpRtnMOpDCTzEZs4uSV3c9z0PDN9By0FnpeDBXJUwvLEzPQrkd0UYQufFTd8Rc
eviCKfYiECpHNh9Ksw75K4TMBQZN1QqgN9UriHYWNhUF1bI2l8CzfbWC51xDq4Dd
iCIjOXxgBaY4KJ6EBq6YvJhS3FHLTAEVE399jz1Tp95uexSbyjsGZDtB3uYZ5Dqa
TKrCvfAgIHcpC+dtPdU3sLg6YZYKqoQL+m6A3Zkirn+8FmS6g+UuKAsUzgHMj6LD
tVB+siPlynO5UvFBYAdFfEhI/XQ1XWLBT5FCXjcVrgkxcixAkEKN++VXGbTP/ntG
QMEF06GzsvJ2IimRs/IxqqdiJr7pmVcQiY1N9ZOAxh3f+9rzDYTpbbc+y6VZbgtF
zBzCusPgeT7+RxYfu6cHWUKg7Si4PxyROobHp/zC+D+qHQcSrcNkoYg6d3wuiazk
dj+iim7OVaoraMJXoDtFEPQOI/5IYAqtZ6yRsEdPN+m+48zEtwiSzre94TzC7Brq
xrdJTT1BxgmKmSLhv0jBEkGuxqmm2gczWB8wy3BAAPesVCJmre/omEh33R7Zb+YH
wieMkLE2xFa6Pm1oldFIxzN2CZoJmfvH00a89rQAmEUv+1lrfhNzrMrOq+rikCHO
a/o1ZP7xAdqRJxGBvcIRpG5iZ5e+s7YG5vzOs/JBg5HVEIrWyh3+fcfvc13UM47M
0vx3R1v94WjQ8VOkj5dW+gjsrB9NEPU3neiM7+AANZosja1S7yZOEpkLVXfgUsrG
YUGhq2zWQ6E/wVTgw8nWLfKdiGh+q9pxncTD/KT8F8nZ/dxr0QNQSTVELBgyAYqk
RLRqXiysgJlPARTQ9iXOlowRaS8ioKw8gz9phWqLIyvdCPAzOi7/CwA/j/1G8Jp7
GhBuFlfkZBOdMe3a847SvBOLcvAKtgAY2OlEEiF3O6ki5xvcLoM2EhkpND9rNSNy
Z4jHpTjH+0vl5SR4/t78YbquF9TBMwzqUHuRPWZOoktaXWMzJfw4G+Y082FXAiQ6
vF7SN5n7G5yW3rAY83J1MbEHDfrmQM96ujF+TaHpi0YbQiBTj+GjC4+wLn5aKoCS
IA6abPmSWnS4LBygXk4Ycde0gavZK7DWogkfoM/jqwR348gNUFtoXVXi+22H51D1
074/a4kMvEPhNM98Rye+mIrKd10842onPe63V8Z8pPOiquBVxb7VGqj0HXT2tjrq
0YkbE/mqHJqO1aeq3MnbarJ5IJBdF28DEEeCspUnBdUCPsv6KzslNKjBtHb2PVWV
jRuFhbBuvWy0jRLQpCcRE7oHTz+Gau62xDsL/w9bdbzez++4g78D+i4mJ82XywSp
5AXxGXe+dVMBXQ77yhHC52XsAGYjv/d5dZArLaVhPX0cPLxNa3RjFfiYXGph6XA/
zCa0EoIQSVQdidhH+z554nDVwfIxhM6kUfVtUwMR3+VisRBmD7QyypYQUu44h3y7
SJHcNYK46HTgFrz5T7+8FHloPazuLWhVi1GfZUsZ7VqHKo0yGZpLrUIEIyHIGgBI
GEtsD1mHB80IqIVzkP5aiGA8n6cl+7iHltWzjVMYVqvOOuMtvAmcL8LwEtc1qh3W
BCpFNR4dDWKSTSTK64jV7KvX7SY9UtymjLTSLttT8NGbpaRt0VBa663rQ9Uo3rOL
cAT7FhEGheLPRM1EtLwJJDL0MTuVrhhD2jGZXisQNHuWE4Eg9gvHUOpWxuT0jaFQ
dgLKMfqCiZGhTo8diodBbe7arXcBgPwKBfUsHNs0fGniw0Dckash/gGtqQezBawb
qXueyRu4wmkO9AGAVAhS2lkqrWN39aNHw0ejXbdJ96Ko+6bKoeqzsnyl25vUMsXN
smzkizL+ZGPYlTt7T+GhoKrxFw0ATOyC2cyv0WIznDVjnNb5Ajb0SQR1UK47C/nA
y9Wxv57glS1eIGuuyWTJSBx2MymitAdFC9MYWbgEtE9s+2vNvs/VwoL8MrNUz8Zk
GwaRGpPW8oYFzHnTMUqv8dhQUKEjXRJpAHonKMG4IFiLnt6zcp13WBZECdeTeRJV
ZYZJFC9PADaViT5hDJ8dnamLJWUqYSMWSyKjfUu+psAN7Wpe1Si6VFQhWGPw3WnS
3qrjNMvWty4xRf+RrbRkFtSIsAgzwZRFHrtMuqxWKIcNIrlj7O83VRB+42QUGgHu
YekXyROQ3B+aGWKrDOaa33nRLykz5dcy2O6ixKVkpDJTnYjeBckiuJw9s3vbdUt9
uc4wK+iU9/Qy14Zoo8bBfiNduFS/WiDfAdYIuEDheb0Tay5V7CNMBUyl6GBOm1Ne
NQxI1RFKqhYIh+3O/UDivxI+a4ltElY9jGu3NFHF3h29gnKV7VWpihVe4puxwYgm
+X6l90qF071RdFFPy/1AeSAMNeUPZjummQ236F0XSBSl6kzAlRGEmtgNk/H4re4O
xANOL8JFr8umavoPYtkibyOuBDLxcPJz5kZCnlR/ai/0xb8Ep2rmH9/hD4HzHhMW
0W5ypteovgrxK8iFPSNfbsboGqilY/eIVZDuh4eUTe6mMMsNcA6yHtOAlD4aFu30
Y7ItgSyg4LMIyjfSnjVh5lOzvpJlMqTpJbHG6BsX/e8AG2WygXT6VGeW4BuWtWQA
KmzZyG0LXZQwPKU63JJ4agQCKh1qJviI6fi0UDZSxuyWq8LdePIXlDyJdjJ6L6eq
B8JjySSSNoRRbRJ52liOYiZS7u/YJR5hsA2agsBiVAp2NhFzgkhdoiZR1OQ1TdYG
Uf1+vG2ohvAnI/yXgmP19BWOwc766f8kZ/J1+kJy74brjXDjO9QQSq1F+Dlfpq3f
rzCDu3euD4KxdGogkfx6hBadwZ+WgVArRSkdu9A1v571qvHokf5xEgmGye/Obsmr
dbbQqKzbOonDc/DBho+ElW7Uj1r8eh/LGwYSOTV4LV+leO1Hf45xQ74Cmxht91Ax
GjpzG3eoMlEPk4HRLaTUNVwPHMj34Az+L9TplVF3WHr0ebXpAoUsGkcuFZ3fc1hg
FQsIVJcBt2ciLbS+BV/SgDTRQxtEquqK7269U7xJW3cz92QtQsNe1tpL6jFAZSaA
kczoxKXhocxvp4eLeUhYL3kR9dQeqE0kqaF0Cw3BxGWJCsh32rKFwNC2lZ8H/Lyu
7buB7SDLxyVYrJ4j9IxxpWe8FbCT64r1Sn2UZGyPmY5V2mHxpkjahS6EqRWWatXp
849DFmNzEIUhSesPREGGB1oqyNxQf2y3Py4YCEM4bi2/Eirt3O5r4lvZ07PlcWJt
tA0oph6UMtI7mpuuMfgeHwNZlqTHeKyfQ8p+AHo761KKyzFX+NOYwbOnu82uGB07
s+HjNzfYmN69Ea7oSo6nrYeoHrfnyauEL2ZW477lT7lw6gQ/+qMKk8sfUc+W3KGt
0ju+JNr15LIIgbka1TmmA7XZQr/hmh8cfySp4BHGYlRokVg368OOOfVqYcLy2LuO
TGvKxR0BSp/Jda3lNGAzmY6zEErnyIkj1AGigpXFd3um73inRoP+UKEjH1HdjjEY
0GbKhXJFVRUHisOHoGSkBQNvCefB8MeeYYXvzWefoK6V4SD+1fLKFQiwfqBIq4c+
a8LYjuxz/arkyOs5BUJ+NX/ape47hddG8bFtg452GgfP1lKL3y4xjPpWZVSA8IhK
DTDne1XLDntVVSSSDlGB3lMDVkhEQa77VjhIB2tLDzsZIeilUp2tjji+6XdGl3rM
tuSQJgLNCsYSzi4wk3Uk/ep1JZrGS86Z9Fa/VE0zUYIZ2WoDVQLRYbASR3KvgeXx
v/+mx0VlSzSRomepEzjpHZ8zC0HEV8Kev7moHYAo4fUhaSe+A6XjCvkSowUV+wIr
re5IMyuIq6mpBkIvOqGAXj8tLOV4QWU7TlprjZ9bnuJhcKqgxGYNkcq97d/9uVVX
1c9ffsU2y877htzDDZv+VTW4E77V8J7wNBTqxwapSZKHYcd86+6oHbtmHkTI2YGb
YJg/mf/Bif3jEYrnF42b4vVDcPjwGv657xHJcyOV4LanJPmxoc7mXyo7+XgsY7ZC
/OBO78vWiXDSJZxnfVGk5TplsFuXuDZALO6fQGU+cBDqp8UkSBMhyOudBNkoJlcy
okz0z2C8Y9vlv+U3kkvZfPiONN/w/cwfhvPS2c4E6xsHhQuREim+axxklp3h+bqy
q55+7dJPQFDw4hCF+R1nPwNr3yYj6arfDnlp8mdH7OxcV6fNuwiTJnqbUpx+dbuv
iXlBYi06EX/5m38TbYTqy8PbwQ+4A/OKu1yYdGUyRML0m4BcE+c2HqaXPcrE5Ajk
GbM6vzOC85h8d9NsSOsQwxV/Fj0+CJ5Z/HObP72jHzrpGPsPb6CpV0RuSec07leI
913uabHkBxDbe3P9IfITN7beIHn+o4Eb0P3PUUSYe6Xg3Lv5mt+xKC11AWNu8yyw
Au8WGbAKqnjhas4GUfp/8zuXxMGOeKCtsM3CJ/PKEOvON5YRn59pD69rf5cUHoq9
laC6u7WDRjPquVICBd4cyVp/7zRLfpYoP/QeirWyaeFkeE/FZ6VbS2cyvgMa4XZ5
15tMO7/HWKNupp0U36FFRbIL+NFtZCaRQiHVNwYmyrg1EerE94YW3FJgd0ask6Dr
uhYaLPKUNbhJL8NC2jNjR0nOWUBwD+E9Fe1R1b+b+MRTcXKGsIWE+/dJ1hF+el+P
14InDByrCXHOO6R7Zou4NEx7BhdOg0YRtliHMuCW9vjLQQQLjIkPjf5yzqjycGnw
+bSKaigKsaMl1nleimxGZvAqJRhbWRmjgZZhtDQMoNd1ziHlGR1H6gijR4W7yR3f
whpzEvprhjERPO0VktGnV8WHPy9z/5UfnhiUxQ5dzKqEa2Ke3OwV05pg5DKBS57w
uf20ain+W4+SoW9SJTkd+oiQcmCMKl8MNBjyiviApqgOPygw1x+9TJsCdHeZ2+VZ
W04DSgJW2y0Bel0pIv625A2ghdzJJs9OYZ4MqkZq0J3oOYiBx0NzhzO+c9TA+Crw
O+06fmWGEqTWCbVLzTak9lJPZa5c+nTKFDMxeUY0RJ5uYBSNs1BFcwVh7GhPO6Gg
o5j2hVlN8CWEDdBq7F2YvQN6DPmtiXo8pLSBpNTays91GQHBZaJBfewXHTAIVhqM
a+x0txmwoG7gej1+3anWwAy6LswzvsFJdIULm2hMJURmwB5vkw0OcOJw9i8DviJH
7+BrgAPaIkQS9LpjQum4nxsRV5pwvlOcogU2wHMbWYIsZnU/ZlA8aSs6thMtPMEd
jzlTCE4Bj5UKvG7AkIsyHrXQo82PEUCKTWy2jIUp7YGEqa/t5MxZO7FT3pvoY2z5
6KkIM2ObiCVRr/8wJWBz30K/eWB1b1itv3hSW8jE04hz6sVx/M0aObZfA09Po7+J
HyPOXayELVxLMasorifmBYJ2/UudOseqTHmjUfrZ5P8GLeCEMxulpPBNCHKqHA3b
QIYDAbui4L0e9g/U64PwAtj/DOFEXJAKcVv81n4Gyge10I3bAUVepuZXsXW085xX
WCQRx7g3HMiPqD5Mvh7O3WtA8QqPsDoSi3fzGk1uPdTKU4W4tPRymv5Kf+N4VbZI
5S/rW6KlBCX89AfAlVvaGmkEt9tftMMrplw1OCyXO36vuAiwe86LqH56EFzi9RnH
gfRW2w3e5YJmgZoy1gIIaId9/RNZ9z9HosaTmmc32vRhC4l33FVpcstOiG7+dZGj
yDoh/nOdnaRpCpTEJvASAXvY3VQMdOI5TTwXrS7RJSBG9xTtpqh927DPvCL01QmP
mSeMaQlkkPlFfdessww26lMqgRz01wJGpH0fPlkptmoqJ1yEOi4s3/ox1bD6vPVg
o+6Xbi0TyxASYchAVZowkJ0jgbBHd0m3egv7JPfB8o63Kppr4BToSnvsDKfZUu49
FTP+hhD2ut16rzoVZl3ryhmKycciMhj27fa16jfvl0VVpB3i2gWYu8PDpAt1UrME
EO//lO9SJGbkBd6+khUS2gUM+pyUq9tyeISY1wvTAjM9dNDc0Ijpkvgshiq4MbqK
AyS0LbZipFYSOUXLtBovZa5zYZtVXrf70b/rDTF6iuxt+knImMhKbDoO18ryx2Q0
m3OCM2F+Lb9Agt0Bz8UIMmozZzEkVNiQBSUDvrNv5qTuGFgs6GPfAoBiOKy66U7s
XluwbiyawxOpQ2HBbHmCrtVWnaZ1FCs/Mw9ax1Qg4gB7AOIgX4SHQKmuzoqERRHM
NbMLRblMn/Y9WI+on8023qyMSid53lEqAWr2hdz9JlAt6R7m1KQ80n/7/UP1pUBv
Mz+pVZBFEiRqG5DoShp8vqo4XFvhaxmb1BQRy8ojMuJbD+wf1/p5Asn9l+MrA4U/
vrATRlm9W8xIldkFkKQYLL4eDfFkk1T6lOXmlE8fRMpo1xlwLVP3Jgrbk5sWf8L7
lGeYWqpCwmZU0rRHT9VTqb93Iu1BRZubYHZ8pIW4FwfzBSeNCQdxEiToDWK6J1HB
FgTDHCjANz0U+I5LSru+SZtv9If3cT0Mub/AS/1IheL1yFQDccMYftPOx/AVJ2c1
Tsyy0zlNKOYhkCivmLWQwWzEd6T3f1NXoD4QBfxprNZ5500daS5fUczOpGFXpkT9
U2GJZHjCgZxbP/NDwTBrvbI3LtYNc3RPFIQ4RRXnxEQsbvSASo6IkfXFXzgABQHD
uuedFSZJEKmToNOeW50uzJJwWVAQF+1sg2KhjCJsb2FIJuX1lXEVpj/b2XblCIo1
bRVQYlA2kyn0Yw6Q5D4S+Mg8mPWHtxnStSpbvXXJ84d789Y4bXAypM43USWZ2cSK
jPIlOq60ye2MHAc2XQhpZKw3vfMzH6w4VbkelnJ+ACHCsSYCjRJdRCbNh144U5Ft
HIqmqRsJb5ubzYw0XJm7LJ/EW95j/IFdIgyAqoKlongTdG8fOACHm3iVBx2WSSEM
a9nIoPBXghG7njrSs3tm/GvuV4GqhJPBF/qNxWKT1guIQRhq+HK2xTCokKbFoTv6
QkEME74LuEsL7q8Q5Tmi/wuNQ458SyeEJfoKUWpqGeEtoFqqD8d2PzidmEjMug15
GwCHM0nBwDdlL8D7YsKGixkZCY5OQN6kVqN1hBHV2kmm23ZmZ2w1lOLFueXI4mbP
bHQw8LtRpBxbwNAIzYS1bQFUvjlmYuTyXs4tmsxhkWxPoDD4g0tOuu9er7bMY5iJ
H59CZhwO0IU8B3VOjT6FGhLLBXe00Pd+ZYlsB2Z8AEVrOZUAHCaz1TECur/roKlM
3shaGuadtSljVxzRwoEaraDWH2526gbriQY9wJ9mdZ+6hB5qfyQttv0M4MHOq/bB
3f4Sv9G7P1TqyFJK2peYGBeLLVGZxwnwhJFdO0Rf70TTQuMCBpVGMTMSyfEyR1gk
84E9l+VHzYnYKQnkoXmPWbfOVbHDxnVAToesFu+QfAi985e/GDnQ5RyoNqIMNsAc
LFPhd5Geuna8Iz1DYAjDD9jziVDjxu9cRUdvUUp5qNBnhNo5i/piBHSTKwfPMM0L
SYGHFVEUAfUA9XZ6PNlgkaiAb/QjmdU6/bJvTQX8966R4saCzDT9fx6QI8gw0He0
lMqWyM1kX2oCFPPUOH9IdAZi675bdbzIeHRAF2akq/vvdOnoOk5ST3zw/3SW3Cpe
gqxwsXJxF5N52JlZoBQnhpFeNlhruv53uWPK2kctWNziv5Rebn97IuRXDua5H36z
Lk/ku7iajipX4tgtVligPa3ZP+4QXAhUopt6rD6ZERGxMvPrejnY1Dlzg6eUDqNF
85NROG0VrBt4pCb5hlLSlGdJaIeJtm7tMgUjsA/ucwkJKqpzsXXyzK2bg0jmvTxz
hwwoa00NHQcRvIS4dxnC9BG1RuFwTBDyTWzRV/BRzc5sTHCOZgS2PQFamwm6KYZb
N8NkwLXIw+WFZCVc3VkQfwWI2JvtxVsSKAxcy7Wc2g29qxlh0YYHptBCDR3ykVZV
1T3/DYj/47fnwUdPiWxIcWMce+hd5ZvFg9cpE2A6kCAJSbtNjXUlZE91TbcAH2iN
77Gxetu2aTatmB6BYFoVqNYZrsBpnFWY+iBLhAvobkV9/U2ORMQZ58qw8iCkgoWS
g3zvd6XfYBirMvWa90L85DlnRsjjD1Y60WXPIFjsxO2VzSwirr+Q9PoDuo8UTDU7
OfajwKbo6fQBLPDs6zHjNyNXM4iP7JzcRArNjS4S4ltYum1XkhCkszXcL9xD9Aj9
nKR3krIdUx5ofE7abEs9GLpIF/Tg32ZKvZMbRzXdiGp4PQGlHm/t4GM14SMzwXiz
3yb6/GJoBmCvwWmtwCBFgNg0n8nM0Qk4waUX7S1uWOprekVmxqKY7qcUm/qU+ybU
2wDd5ub+lQNsQl24BLOpBUSxWYZRu2I8jJyNbkzKrNplT2Q3EEjj9C/nYluc2cd7
EiOTxTbYhVlqpLm9KAf38OicmybNev3chZhY/sRK9iR+h54dPM4LAjsS4pqiC2pF
bZztozUiUnRArawZDwYjQ0i+Z8WKSD8bgp9coK4giw+jV3xgsxB1RHUef5MXc+k3
V0YN8LV6+ICepkJ4vmXpMWajvhcvFbxxAeslXh05PCT5GvkOCKp1+kuZSWhYeFTY
EzMOuxvabZTxRDwpv2Bv2Vl6+DjwqbHLkZ+AbckGZGgjhZAP7m1OehINTmzEB12b
e14O0xbxoCv/gMF2G+Vfj9QDxCXCVW2EWznMtpUP566ZNcbX8HGzUoSZX/Ta4IW2
0xgEK3x9WGgukHhAWOOUiV39+R1RYlku7/a4cNMwvnOdNd5YxNO3hmxsN03IfAZV
1wGhEL563lQZbDkvzEb1mfwcUdoBT+a5LjUU1JYcDHGrAs50vA5K8fMjMG01u29i
H3HTTEf4a8YYGmwKmr7DHkuWFF9VhbpDxwj2nQYy36B8+jqRgMVS4IFs6aBToqbP
kt5t8lShjAi3aTFg6Vt8loDQI9owH6v81Yu8pPnNJdvB3vgWXfIBvMa7dZUcaeWp
65/Jtd5PkgHXYQoo1EszJiXk0mjA5nlhwBHT9KxZm0jT/RzuQAXeLEMm3NAQrcm8
OhVwHCveUb/JgogM2QX/vEPxni+1EF/XjmDbIZjYrDmhPdti95HVRoHQJOoKT13l
bTGO4zznNYRJ65oJbdpUCXfRQZ3WXcGUH31MmTVTjaYDY8BoireFY2EbvaZB5QG1
oEBGOK3ix3yMfeGhHCbiirymks6j/q36QnME0OawHON6V57sxfqFTFttkkjuKYDH
Nj40D3hxmCFLzJkGwFGA3wVw3b7Z5XjlWa/GuTVu5oL7YA8fmf+x37CDT7HcCFo4
wBFlZUiOxOs2b/IWCx26HOjQ5QqPZmu9kGWRgmc8CbBK1ntY2QqwGmH0HZGHcu3n
31YQW+zMLJQcfOR+rHwpeww/OAawvdM3imHT0LptpIvUZTpxPZ2JCsVOf4iRrtdK
3zuhe7s+gExlwLEiGbMfH7illBD6RQ8e2SoVXoSQO6FxuCWzu6BC7dZOic2z1Alv
UiyqhqZS8XGDg40h/CuIvjZSPrE9AttW4c4omMR6uplHjas4ELmBSHENtMsLbYr6
hxgZinEnxcG4wJ7LihXgKmsQ4MxryTe0emidARbYxlcFNJ1KIaTpsbw3IRvDafm7
z7iZpzYieGejLLlLjKtIrWjblOolGnfpcc22Ujw+Irl5iz7eYdLk7aLfJyuWYFWY
I2wBnGKEnCULr+O5wEni6EUsrUH5Df2IxektZs3coda8S3WTpQ7bOPC9a+pU1hpC
wS4Z1EanZ1L13MZoNvJ0K+F1xGVuJCYbsuWT8mOR7y2HuUL49WA4jFkR2xvNQUxt
7umrbxzhao6IgkZPDKS65MZIzta4FDrULuTCTx0YPL8nFB3Q7VdJB3fucnRDH5mG
mU84wGq9SXeDz0eJr76Mao8NH1MjQCREz+K5kxr3Hf41TGdscJdv+S4CdmePVczR
ZWe+Rq4FJ5IfylLl4geWa/r69f1niYiqf8LyDIayC8Vu9FqlW3HXIHKW8NoVbrHL
KoSGIQ1NOFVgSOW3OiVrmjV4TBTOWW/qBHtaiNuz56aCYtOvypYMAXZwzm7bbQJW
NUHGTqjaz/Ef9jPH2Ob3U7MbNwNt962vwrtedyMLBK05Zma1V9w62bl6KGmbq/MS
JtFtAN43gI3bVTKDOHiJsbUIEKpt4rA2nDXNsArADSRGO820i249yRoPibHTl0M3
IKvzpeP7wxj++0648IK9ktlSJp5Z+cknNirWK7ZVjBq9v6IYDStgmzOfHvbr8Tly
Ev5Nn6Wt6Wi+6i1r57Dy7pRZ97iLFzzU+F3rBx0JknZC2O5JOCB8jEzlNm+AI3F9
tLA+MpRnXhb5qMtH2P1UoXzd1pcCM6NrA3L6tYHBnAI9nzUCRROapB4zCzY2Sobo
ZZV4EPwZRxcQX/46cYkyL9hjjnzIP54jFR0kOqTe9QvkNsmt5AJSv5iBngXVO6Fd
JMeBRIsHLPE5BoENmk8ZjXtp+3XJkASZsnoGrTOdv0CYvCZ6N9lZZ/CzzvPToRwy
PfHEfHLDPpIAbm5HPYN+JA+JNX4LNDRiw/K1m70Cwfc/mseWmZ8IXFe4l1EqLei3
5KPjk91BlO/G/2CHexNv3pZSgbAaDRNYXwkt4kT5rPN5U6XOJ/SVuflDmfg3DmQS
ktH7b603ZPcC4Dr84Q+SdrEaUnR8ITLYZmVLxT41ykkZGZAU9ka25TqyjeFdk5CS
QQIrdmUZbWGhUMnsRyc2Cfo8jBB6x+d7TEBnerPaGhvcgZ7q7dpc8xQS8w2wnoyG
UBQApB3MBLpxS5qZRlQKOx9Yc6ytiYQ5gGE0y2VzDm8K+qire7h2XXdLAZT+R9Wv
hVxgS18V9MaLW8dXcOncTU/esuwSXHRItr81Zf7l6mvmiLEtctZn7zh+mjGcXC6w
j9kA63n60Xj+kI526IB0aGW9o+xmzjS5AP9ZgPA7A56GBpONckp5NgbcOR0AQQ0z
zQtGYxOj5MtoBQpUYHLxuT+2xJEPHiqWQgcq7nNvGNQOqVOreVUQhGZktAUNw4Jk
9XwVDK8AFliozax3p6rSGvJJTpUaX3ert7sHLiaT+8fyuY9NStJ5VldwzEGh8Pyk
mTEYTu1Zls1eFWAz2NTLZhVWRPujVEPsxXmrp6zI1xBQUR6IehUk2EVHb2uz8KsS
QoBiL3YQWkB0rFXNVkjDIzgU90bXy3xJLhDPAHY+ErD4Ma+28xNmO1tJ5NrIf7Aj
+oK1OTBQYpairLQ8c1g7WaEhkwwM/piT4HgDk+W2Iqe6TC5NsM3oAHBHaAhA2QDo
Do9ntVovYI5PzGnwBeKnhHxnogxNHw07lsBR8crntjNTuqIu6nTaS87DedvrcGGr
sMhoY/6bfpFIPR7xreIVZSk80ybMyEU85zQi8IQYr+hyluSYQPKne4Rp0eQy7a3h
mV9qrpqIcx92Gtw6LaIu7P8f3gQ4k/jvc33Ao5s9FZFADtKAFH1m97d2mGCsv2S2
UMSYdK6dXmLqYKE49Fax2muF0TeYk5DxciQ6XqfD3H4y7/T2pFAZV0JHUfjFF1TV
U0lR1l8ke2nJUwhAG0svYH0PFAza1beGLv3c2zEVBHQK6noPidQoQZp6uudVWsvX
oEecicqw/D22+qTQk1eXKFsoTv0zE4LHke5P0NaaStu5BpDNE9cheMVaFCP5Q73F
Mx0Lbuyeghutzk7sH4TwzHivkQ1XuJ/OueNOeSfxukYf5jIf4MK4xFl7qBr+7XK6
bQbKxQNZDaYHGa0FKrZuxIFZv8tiSrEyVykfU4xDx7Q1ayna5s94jz4Dvxtv73zE
FxCtMPnnR6CKlW62FI//LtCoPm4SxjXENsfO2+3CoO8pKAQKl4v04aRRK+bnnuKg
xvVDAayEMLHrF0Eegc1td4uFdJzvkSBh1Fsf3ikB6z9+uZJICzwih5qmEa0s5j9L
V5wDgEcAorS/lOu1FsUb57oMnb5A9kX65c3rY7SIws1EXQa9Jzev+FgsDeGJ38GU
+KzvWJ2PsnZHfNDC7Ts6vj9FUdhlKHBU3RKimXDHF3mq0Io392sVhnw8sToNvKul
YrW9ILw9Nm0F3tKmkfH7hgGuq67bbT9V7m3X6KR3WePq+j0dw0bIMTQEBSFp0m8U
FWYi4XvskGKhexrgSMNYwmW/789ZfGbtMIJAisobe5yLXZid2Cw6nyDuqyxR8xeW
X67L8ZTssiB5SGrvyfcbRpHfBG/X2RVqLOlyTJpv76DbTTbh3GpxM3pCLIR+Hm85
zb9VYhIIXrdGoS7oQzWsLPtOJGE8VzXWus3xlTZ0rFz1w+PXQLwQtKLExd55WCGQ
Mj2JUppIL9r6nO4D1eAins0vok0qiGGjt2jJahci8iDY930y9j9vU1R41w4IS/Dz
GWvea8A0Kj6H/3JdMUPysDUNKZncGeL+vMt+RSNM0jwVcEX/SoELSjVOU0ctIWcK
IKEHASRcaVC75L5TMQEcOh9uXq0gT6YCjbT+Ji/QgRhoDpEFotNAPsf/Uyk6kjPS
0av8Ulf5JjYWwA4NTguaIzgEFhEWVQN6XNq4E6zmTAUlBA8VKpzJRNwUdpsJH2CO
JQcb9Uf7e5fVVmAiSXvyEl0fWtv1kARcvxLuyvihb3Z55us1mheueex6FE42WqHD
mRy4IXbbmbA97PA3pZGB1zRdKoeCNa4tZXLp0O1+AlEOUzGEjoANfS88WxHW4tln
uQ2dcwiOPvgMSJvxCbBO+o+5NqK8y6lFYUfu6OdRS0SK9NI2tWNUnhwQSjlvogTY
1KS2Ey2aVzpJY4JS6H52edXy6AF0kH2RxUfYbXq+Okl6iXasvIfsEjd51Mt3RHHt
p31Q6aXmJXu0o7fJbp+35iic0eZqvlMJnMW7Q0dpQ6J+fxZhvErcQ62/PYCXfLz7
piubAkUYWdaKlBs8HX1EtKCRkXIg/qfTAI7/N1GkCAux0IcJHzhDyp9nhVdjYylG
in71+9koVyBJxmROYw3tJBT84CjX6c/xmNqvi9ykF6NN0MlvQQ51/ocMLQ7XIbmI
iCRsw3heNrBomInK4KGRXLtsKYgRPDUVrnTrWqcafuZ8r908fKkc6Vo7e2419JJI
DtQ6WlllT4tfm5sYehq3EwWMK6iJs4MfJtNEdGP8pFVNuhXnTsGPmI6WSnqOcs5I
DPv56JCZFyonT8AmKWVivo5HPwnImgXXkSVg/s3tGpxo9fZcLRtF3Sw40Yu0sNtl
6NyaN9t3WcAX5xk/zskAhH5dYi37dOJaL2tnzbZjfj5yjhrcpzdpApEE0UiNH62c
H2jO6jv1GDByKJ5TXQP/Z3Pnru5cnSb8vYpi7qOBqKE2gYpgGJm3nLAzvET77RB9
GFV74GyGD4u+/hNs2mz5Ql9asplg6+DM4Z1GXud/5HFrWiKfja9PyG2+8rF0ZRh6
F56jZwbJwwlbDpFjxtO1KBIVPmiZAafJhT3Dp2cwy1Cz9LKNTFqF3dFHWUKCLfkU
1kB1R8hJLLhngiFg2gF29eOyG88w5zwShstsZYGivIjO08wSvCgPzEvEqVLvmH3G
IGxycaypn+ur/00sSDnlEVpUcNiMmb6ttQK2HTu0+aX42NS4MAO3s+8Oy+cwUjqN
JHhcUV6gaxyrDXQVYluT+0PtJkQikAj2FrYp/fRJ8w6U33nYTY9rmyItC6jZHGRL
Q+RsI4Npz1yRNJF2racMAPEsAQpB35W9Y+duI7ihRssSEDxy0yf2HqUC6gjcCU09
j9AMNGsfDiCkmcqRi9Us2ktDkH5Wp1zcmNpbVAiWR6vvqbHq7AC1P7a7UH6y4KmJ
x1oXmfm3Sdr5s0PFiIA1PpbAQCE7FHOXayl2YkYaUzi3AAVGT95ka9Uu4boJWeTX
Lkrcx4EXbm2YU25q5SYdcFzvD9HhCxTFzgnznp/dwE4W5DFOZ8BZhAb8yhrwX5ye
nY+YP51LkTN+vPChZ4O9GIQZNLe6FH+SqSk/VWakb8pHnOV+GjeWxRtwlkX/bGx+
9itUceJhcWqSuyCH6XFRLHKNP381P3qmmPhPXtrGKPX6NgBgFehB46jD71OKkFBW
oBdlYAchUhhgTSoanvQYlHlKlfdzif1uxpRxjr04d7fTTP2F5CWrOEiIlDzdAx0A
V3SjmJWxoxVh3vsKa9aNmkhIXIzvkHNjEdGzQlyuk29bCkd4Lvxm9E1uNXea5m5e
m8vWZEZ2W6dikzR5AaaHnhxfta45X+jcdMOEy/SeSPg72zAfjzbMD4h1iM1nKQVo
S/D9r9lUYOFILuArtCGl/YU1xjtRqh0dzgWaPn9Q721maD/Z55ZktkJ0JNp5n9M3
BffegqMqUJUJGzLtJBkdg2UFcb3zXf0gkoP3bObxwiKfIAWswgw0BkfhkaQzG4XI
Kofzb0/0aCqG0kRGAk3kM8X5DdfWvO2EUreJv8jCihJoY3A0X/3gE3W/en5uj3ZD
mGbiw/f1Ws3xwWImpIF1Fwe1FHcOq642eL0/rZojm1yHOaPKvX4oZp8VF7e5DQH+
Z+ADTZWeLmz/Z4ko0G3yOJzeL978KFNF3avyiVE32OoO2AXYWOA4CthExAdS3PbO
niQoAEY+FEp6DrHyuXOOcV9w71Z+Ndf4SjS4f4zpnXVja1B6rmcXbbid5dRifnmZ
ghneJg50w/S29dzhO+UODs3eqXvBaXM5O7yTY6rI835q2RXGnoaWEF4Mj3/P3idN
8smmwjt7zkDa5IAzRcrTxyiyckf87ZnYoDM3RxuKZCHIwnHHYvu2cCVWTUEDu49o
ZnYPaDsE0dd9HL8BxtfZ2KK9xsrJTJsuPecZd3toUu/eg12XqR1hdUSZRD1lJrFI
vTEnjZBfJPzoN2oyzvgXi8P0NupyoOONlIYwP5IV2phLvYh9oZIOTsjThOcyyOVt
oB7GqmdZ7n2xr7tNgfwlLKVgwfNZZOIUadKUbs0D2FvCWzCika9/ElT1vi7xmqnR
gkRp2ppUJdmf2Xt3MLW/iA4U9/TyIoDwa0z4J9i6CUKUQSX/ip+L/h6JIMahuiCy
zX+WSvFm6iHBNpUH83a9S5/nfnK5Rbp4j0m7RGPvxd31eS3VHPP05yvB4tb6sPEb
KahSnYZC5Kk3Ne/jxOUDRlit42mCzZAGTeshW2kwgbkuIwS9ClQ/8t9cI5nHsid+
oKtJlOMyP8c6knBObCz23MoJPR19L4Fhl9JR76SKxtmcTsEqmOGu6G2pVaxh5aFT
RmTAUd1pIvtUa3Ob0uY5Ope8H5lsGhokhIulkwZ6Z3GOqctplK4EY1pXzRCT9EAF
c1rzZqgv9u+/dj7MIlU38pvSxepJ2g0Rxk3a0TYavNzJtqJpNIv8sVlkZJDX/VZp
pK8Hw7gZFNNu2uHK0NypjSYyvEosebyeue/kge4GlW2VRiXVCWmwPfnbFSElD9pN
vgnLpYoPMS3Z35M0zutlEQyQn4d+VmPiREti1Nki59/nRfmA49UsbYmYzCi/ebY6
wJIKlnVYrtbHIBdfjHnbCp7kn8Q5QaO9pg/HhVlPn2GLESXq+L/KcK7W4Mo+IIJv
MVufKHqLxSBtKUXKkVSCVKdHVAx/O4uBfavbKBz5q5xlXOjG73IeYsrifufldLXz
l+U6F9Hbo4FlG4hr/DxisNjCkt/t/+C/F8mvoqye1sXvDPLDswl+ATj6bDQw/wm2
zFNPRvjeNJMdQqis4b/DvsLs/Btf/3QIqFUN5q4UFFnZXPTx8rwE8gycPNWzuSwG
XlRPjJb3edamvxvhXR8CywZXVqjO66fmDs/PJf4uAGC4A9mmeboR8awDz50d7byo
w8/UDBcoSqH2yjsU6UdstmNA3YT2qVDQX3+X9zXAOhguPA0qwbvJ/jZNTy56CNYH
F7CjBJf5zVbCWCBNQFJeqhu7Q/vRprwTi1Milbhy8bVGgGlYPpchi0HNwc1lieoy
1k11r7shGkx5/OTODbDnRE/dUdwG0edoJGvmlCWiKtYPzUtYdOU1IJDlcSmrEGEd
tEJwCjS7uAduZit7zmJ9mKSYLOCsce9Olc8dgdT4LQXvXGSnl/depQ/IqiqvCW4h
rm8e6E4h3yhuD66x2Je4hcsYubMAwxfcvm+3ROJEXRVER4bUVmgEcCpoMS1/tOw9
sDTSJMHzMBxZBpc6KCfbBzEjVoh3+uzsSpRIqaTUwxMKIiKhJZzvEsQgtbLwN1SI
t1fbkp482JAM7n2N/8a++2QnnWnbKtjhjdPPsQ8dNhpZlaFwwiUO3/KM7rujPIFS
sC2aNh2ShCx2Vdww77nDg8+lo4dl8q1eOsywhpKcuNZIJ/831dUp5gc+yUGnzxCD
iwl6txHLvowz+TuzbtQmNGMH9+wn1sZ7TwuPp08aZwW2J/qADCrs/FYGZEiRQHW5
BEBYgzkj3CiPOS/Uc7YKKv/Jvev50K6jGYohaIsPAQmNk4LQlG+tVMssZG2fWPY9
YcO+ctPQ9hrOEmhK5PsJFvx0zVtKOT+9Uck/86FgWjPPlOiz9JvQ2SynQgj048wh
NfQMh/5NDJX4RzJSmwREncrYtTSeG1WmRZ2gAEEn67Xx6EHpTDQK3TDKRi02+LFv
FMKove1P0bqDE+DDtvk4il3lfp+OqIaG5hdza6R7/eGzD6+Q6x/QcZzsyKq8QGsl
CgVYYaAOGCDxc8+31xAiKk8IGqZDmYpZLQ2z65LGY0RBIGHopL4xJHvQk+lgvXuc
+Tt38uoDhVgXoqY8eSXQ7BYIuONhcX4iKxUlCmHKMap7/lFEEI/s3sBTsg2w4VVH
Qn9IwsesXFL6S75uKWaq5ExlEv6Pbqb4tti+yIUSnlrJD24TmUx0AVAABM8Z5dTV
d0KtrrJALoNmrllyytJrrKY0ICAos1qwmiJbRvtpbW13j8q55JM+gJ9+ni2bCk5i
CJ61Tg4goqABxBpkl6uL2FxP3S1yb7wcPbt8Ivtx6NeaaVk9QFlBH/cvusFOy4YH
ll2vI/JVAiKm9LZL0EE0Gl+XsBR+W/17yS+hZBUS7oeJd02Pwase10lby7wJkeHs
BGenXHylTbixS5VdtP1gELclOTYCVLJ81uSbcd4H9teFJ6cWjYIO6ZozZWAMxT2d
oeinZTSX+XaWF/3Yy5D+7FeXiWkynSVqYjny2mihUeauUVu0vrDF+DvvQ5O3BBrS
Eh3tz7WnRIEWxEybt0uG380KS7g8Il/xuREydWGqHNZdY9oHKTgNw+Tgo5+JQduj
JWRbSTo94YQSAO+qdJ3J0YMioO1uvR2m8KFXKV55UAAqwbRnUUZ0JiAScR3rahSd
+91cZdnVp8QzbyfExg8T9R3Vam+0F8o9+ZwWkCc8TjAyPRhES46L47qAVw00uCZS
6HMWKO2H2PpJMGePpC1xfGMPns3Dzw5ZGHE6wGGLSqgcRkrUMfOzbV/zNCs+SzyY
f94L0ox/PJJzEMIRXQW1c73+cnTpisdm93SFNJXTCuiuyBzNYhQyN5B1hCDNz3CI
yS0GXH/57C9/iDfoE0BRzlGCbBk5aAJ2BccK3wUSFbxEsitm0mVAflSfimmj+pq2
uR5XKlRxGQactOWiLbtdbyn2tDyO9Fv8bkJEoHf0a2GvTiRV6U4Wk5wgTZNzjdQ1
kTtWAx80OFNoncS24o+BSOwLXXpUp+enKRS+P2ZNKbkBBUMdrfPpb0jPQijPPkdI
J9I1KZSgtItFc+uXONXwwziZGm+ttseNJqcC/iyTJlmnn86CZhBYMaXIbHFsShON
nL5Q4MRIqhOiESs2qi3TT8hEXZlNfeiUxNUGlwBhMSbS47kLzbHV50eRoQdjUYMM
B/MyxmwUfntBUubEyKjLNuRj5A7dzCKu24BtVWGKerek0yJUQzLfDlNqInEkUTkp
IdOYbbZS5xPk/kwfD/28YBW+xofq/AKMCk/b1SbyZHsk9M231teB8d3S7emu9Pe+
4scFFSwgHrzU3nY3I5VpYwQGwFHW6/Hxd/0GD/9jnlK5XBBxnoqzG5PkpIQeUqUA
pmO+TvJDwsBKHjWAwkWTgL90r1cs950yaIV5ZYnxG7Kw6jAph9g/mSaKzLZDoYIq
gC5VppTbPDzWYxzNKH5Ho6mU/wZeKL5AII7sOYqvj16yTfiuWYqZXy408vanjnFd
yBstMG8mrCybhLkBx4ZEm+FSB3Ndfuratv8FvtOyhCrsXM+stsADvBp9lh3tcV/y
/rHE/vc0doJXADZoM5pIh27oocp9B57q3LoV+RL8OMDgnvZ/+HBblmuw7vb5HODS
cFPExg5L8g2txnTDIQmXACBQKDXK+QKJUdBwhECW7i3T6/1sjx3uCOxNKJeRqgTN
F4E2eemEY0yZpb2Zg2NuNinS7BOEI2L18skKQIOze30UaLMUmPioUD4YnyCfonUK
mNy1Echd8/zRWIPFVmIsyd31jdGip1BgP811eTiWLb2LaSBsIHWJnM2ay8cn9GGE
qTc5C8ga4HkzlQtDNKNUhJ5gubBHQgSq1qfND7vTmuVAnvSAD3llDUgrpZDhJ/hx
sA+ZtYl5ncsxGWYK+xL6nq/11nkFvkowcHYYWgc99TgqfQVhH3MyNVZ3GpyCmteA
8/28PlwzvBImCF/7NISttma7d/TultKbxSfHWYAjLA8hEBbJgUOLw6DOVjJ/goFe
3/WchTuxUmqg0LReho2kPEya2DWTEfir0HuYHthpJA+KePgyBcywbTcxFwChO4lA
F3rvsb+2Jnse9vMo6x+pFrtU30Kiw5kA/Boo2wXsZkiJdxc8h0ZADdE0lqXzB3JP
I0RjuyGCEGj2uzfvS2a9/GJFxoI8hjnF1vw4QjYGI+gELiL93+/VCPYOTPIBlBh/
hBKo2AabmEdwcK2xuFJFEv46yy36HcotiO46C+k8vxQuFVMDtnNgdIUlvuybl9Wg
2RLY5QojzjAN3+yfccSfS6mKTuLb9PNgPnyXfoP0G9F6c5IDBb47uXsmfJo0kQbB
QIkgYhfZ7SHB4OvcI87KJIRYzVIfLv+81X39+qWI5DHO2JBVr1xkUWBmQs88u/ob
IdlGQHUFIoW3SH1Mo03Eo81tJjbEkkudC6BFXoFdVquqLnUo89lY0JUxQ3hCKRvN
HeADlhRHorSyMYH6OpsOqCzddSSqtrcy3/qWOSmI3koNdHHub/zDxRahFLKmvu+9
+meEFkPL1y6m3hqKvw2uNi0XJgK2xaUScXOEhtcOnn0bC8T+KXkBCs2gPQEnU145
RLfOqAyTmtU3SZAQ9iGfjRO3QirH+rAEItMTYUn4+n5RPae0T7YZ9ZhkpOWx/4b9
USOHRIfZ+i9l39Mi/GdiIRI8eh/sPX2mFS1HFAleMbP5Bd+iAqI003BTh2PXZoSI
uFooMItaijXAK3ob5MrqfyorXUOEkfNMHFrQINdf6Q9V86yTtjp6R9RYFQRBxGBL
VRZTPxsq84N30xJaXsfeBxDK4O0+mdX2qm646zvmeNgsuv4xsDdlOr2AI/eKeqaM
DUY17C+Tlr/b7nBDI+MUI0rApmwXWXXOm9qIdPOcKrp5UpvFQKf6Sw3ofLlY0YRs
3RO4Uo0+ukj8SZIZAhStajkAssgct9pn8yGYwxFaPKkilNRY9grJOUieke5JfOz2
4RLScT881FhED0bMmcIle47cNRn/NYXYvC6RTBvlPcHF74DUaiJI9GmtbLnRHyGI
HNbNamcszDWqkBQ1c1a+TCVZxLH0dDR1WqRXlxIr8TIRGw7a9nHM/xQsNBhV1RWd
A0xOaPjBrM2bPKgkVO5dQ8S3rptBiutUsMRZwB3IcxEW6BJTBDhFZ6kOCIDdIzQt
Zeddmyk1qusn+/MYphKiTM5XJKnfLMUgI/HZKMt3X6uVsxTJ/H8zz0/fGwzjsJXn
YglGDq8u/qoUFF42BVdjiwJDMx71Yl7UiYrSQcZCdzeV2aBvpjSjY3c8mXbfet5R
8WlOF/ZW4O3kRFuX0XNF3Sd2ecEFMRnL/lP52dHsgfCi5dxvbydDyx3zfC6xYjRV
V2EYicydSdd9sKQWN6oMtt3QQxwAy0t4Y21NoicjWvwY/1pU6WB/j1yJReuOBxRM
TeYqK3xs4apjGzfUceGyqzgqWiSsUyBSKcJWXpubekH6WrfcK9j6StJ9s6miiMKO
rel7CBglwftR3s0zyzGcbl2Fn4K3Ptjwf7wLAv4uqiKjtc5ozgWEhVDYVum688rU
VIXnNAEEvEOXwfiQwrhigV5Y9TUDy2J7FCh+YX36ozgFmmw1Gqo8Wg6lo12CX6ZI
eV5YhpKKqRqTb+mhbc2G2KDQcp2ziTLwMosRbTwWn8ovtj7EuASkmaD87cexkzWp
tnzyP4QKQRCmk2/4SBpkfaEaTb028hd4yjNCSRr0XybOMt7HTHO8TXg4Cab5AOLY
jA9VbM9rty3BGSVkpCyo9sS7wxdd0nW77JamYrEoP/dyywngJyUHYbfShgDopjEL
DTtRr0Z/qjmtn7n9Gai5HbIGMgZQN7AUEtaVOD5/6wgCl1KdIYhwLhIDHHQcYXHD
A5ARqg4CK3czoSwZ3r2rWn6Occy1sfqQCdrUehhuB9STN1ZMPwQjgcJjaZ/+DVgX
EzEwn41HcLzvoiao0RpQXmoZCl7397P8Ism2IYDC38zUD1NguYtRmzb2YdgWlpOy
Tq/s88Q7K/XgNLcHUz22MxpFfKG7Kk3bHIwQdLlUecfaWBZ2Vj5pUvUX4zpbFjUs
gyhB6XGxD650y5D2uWKVNvMHHHzNbnabCMgiWoIJB8vDDoQK18YKqsxtvFzox9Kl
Hl4SUkAJWCR0NACVtzFAcce0O1hnArmJAX/wF9/BfLmZ11wLIF6uwSlbk7Hp09nU
bXH+8yqPYOd/Qzq+msuSGYKQkoYYpeRgcOForfDAqZcdwQG1QfKE3IfRu127rn9Y
1oo96f5lIy6GjgrGseSikvcPmKTOXPNzveCGFoeuh6CVwzJkhSQJhg5j3YKmpUCR
CON9hhT4FfjDE3v7z2TKZijdG5Kgg1qyjzgNgo5NoubbvjH9QncYiFQq4lpYNVN9
jCfYf9X+K9lhvlarjH7H5Fgved4Kgs25CkWMKs+YjTxBDZc5p4IuDzsm8CzrYc/s
SV7Jj7wBYgF97zwXoIxdGb6Sg4gZ5Yj22nlT/mx+rSx9WiYwJArv7/ZImIwizr8E
KgV0RZCnsQEDBih+lZkNuM76dw+f4zDgkmFhpIUv62sGhqcq0OhWtyWahJo3SBxu
nsLUHe8Ji0svmaCFJUgDiZ8LtMFBQwKI0v8o01o3bJuFPzOwSpolLDeojRZy2emr
B4dSwOWe9XOokXFO4bI0bT0rMsVboCQokAvnfSsp64W+JQmAT9fmIMyNb17V2bxg
0T8t7bpaP1bZ7VsXjLzrtVajBOXZ0M1++2+6vubTG9j9O0eNVYjuToRCPhhzotDp
uOQU9CUvCqqtQGhnlMCne4YACV0UZslvr1NyDwv8LETFRuhpYCWWXfnwMYAEMoBE
LqJIpOBkNmhLMVrBDnv6mxfEkysg+NWfTm73EdBB+zvY8faxiRJcHMzMhaoGkwSS
FvB2i0qBi2IfgeYTyV+FtMwsYRIEAl+U1+z4wsPGwwC8vNlnVYn5R+Y54zPH7laz
iekjK4lipMCYFVDAdNTV3NIW+THtZ9Uf74Y2ntN/YTzgs1IYplKxmAjeuoHmEJm+
S/OzoSLxEZ2uWYfeLgYrHvsDk8JJYuO0lim71c/va3MusiVi5eYew1HhEK28UlgH
TsFAnfPhs2gKkauenK62allr8IlqUdA/LbcAp4ceQGg938c9BhmY3iAgjlFMzw5Q
Ia4zHOeJ/714+tjilQT5BnEEy9uKSsFKs5EF/o3vw+SLMSOjbgrvFEDg7qmxGelH
53vgqfn6Gezf3kL9ho1cSWkpM+jZEGcHH5NCz+hzsGP9v8MAa3a++MuxPbP/10Rl
jMaOh0Iqb9UguP5/s3UVzTC2DwcsAsRGMv5DDX5E38TQlZpgWbKxHU5EafihmZ79
0EdP/Yhg9zcVmuCFDd4sazX1i6l6kJ8u43jybp3TPlPfkTi4yO3TJYMM0pmbrXPk
EnrCMBh2rxpKGUjHXM44lwTXwSOxiqd3viiJANyneiouHjrPyPkMAkZx3Urv1Wum
h95Q6Ury2yRxmP0sBw5b5d1M7bfEx4pQbPgzM6avvnPNhGtOkcco+oAcW1og4DGX
tgEe2c4TDXHF9OyFDtQa1e5ADc7HiOdYfs7pX8vzFiQ64pAj1noBoHIjkf2YmLfS
8zlLPGMgCKhb3ceijlGbtcdKtJ+05RDkKAqi7R9PYqFrLlqFFBi5Cf+gn82AWkhJ
NPUxCzOIIL2rlscpXTIcqXWukTK43CPQGGhMWefwXsctsi3XM6VYrUWZKGpoKuvM
WZ7aEdVrA3p68W8HIrqj8KPo6Yz2BAmn7DYQmpUZXsobKyUJXLN04941O1lLn2d6
sNtOlwp+lQDSAUPv7EnawX1VnBSR/PtIticf2W+THcdTs/LnCb72uN7R/k9XOQPm
i/vXsyPCaI+2bkATQpbAvzDilzQmo93xtlNPGUEWidEm5ZLQz9Q9Ch3aR0QMxEAR
pW7/VzwqGLFqoUYpLURWK60iKgAOXXvPmLJjPL6pj4N/EHlVjFd6UhRzoLS9rNmg
vqf/kZINeQ0PCuciujAm86Abrca7GWN07kTh6S67mhboK1PUUIIp6WYoyuTIjNUB
qODqStFaZO9RYXg+bxFHyVL/vTYbmKaFiFzt1Qb4AoGhdAZ5CLHJL0OFbriR0HXe
DY/e3hjOqEH1Zjqz7s1qhphe8x8Xx2WUTsY2bpCUHXvfa9Cr1bQOEKMEQbLyWwpY
oLXrbANtbnwKAuYRWiUp7QcOCoump7LEd46WM5XNbBSDNYi14JTRKAePegT5XjZL
vTQGWm4HDQkYvHweTegnIKk0b4bU+2YWuYJWHJ9VEcLC2wSUCz9yxEINfkgV6XrB
RaD4jQ0w9Sw5v67mYwhNn+b1NbDuVutCs+gAeBm+ZlCKdentPQzToFdKawf2w7L2
66y+yiStJ5IBASp9Wzn/HlNuA4+RcsX7fVzTJAiOr9acPuqSQthkooJz68XRJd3l
jp0uwwP4WgxCubJ90z0b1ggkqXFsYbRwpWcYNAJ5yP9nQRkLxiLxkPTrNfj+Ej5Y
zPanqq9efJZwi9nJ/B01hJvUGnoeFLeJ5YkQeenMIhyjsjs6MIraZDareTPENHqq
bm9+UE6rURLukGWkFsW7pJXPG7YL1upbzFBOngTS95aiepI9Q3v44T3jykF4Ys3k
eL+ogIu1VwxMwq7qluE9SI836UIx3BoYUOeTlhPhbGiXSb2whbwjzsTeQVeF362V
+ddSKSL3mB/yqqjtirpImn7dQkqUavDZ2vdWcCwxBWIOX/NItzKKo74P7ziUVQKu
ukQhofnB5ck7XPsfL8X6wNmyl+67wYyJNQ4q2iazAnWD1lmJ9aCnFsU0ZY365ekp
ufldH/uJSOrU3OFnad0DRqncYKkQKJUqbNXvMUnVhyITCuKKpWTe42Fju82lZDUC
tnIoDWNuCI0G4gpwPwSU1nd4ym7IuiO4P3wMZmk0IVR3tvu4vSIiBvYwcAz0kiW0
UDqM8zHWeiNn5CVE8pjhHu1YiPw0FM0x1ikBvdpe+jLb9X2OE4kX7BiJ+yneVVSB
+FDVYVA0CpQsenOLpbqpDlZ4HaQSZ5T/A5kuVtJnHJ/hgOiGjMCkyeQ2DfAx+V+0
Rzy/lgknjCCKO5JQF8tQQ8u3IflX6XS3Z+ji0CVnUVrMGwix7tMFqx2VbS3oQb/F
aljzFr3h0kGCsXI4prUakR1YAcjnv7iI5MEN7nVpG1pv21WsBsbimUoWFtiVRsFI
iShwo7zo3H/0qxMvNLELHJHZl3B3hDaDP7f+V/XKyEn/10n73LI4dmndqX5F9utG
oIvn9TsgeFajYyA6aVM4/y/irASFlIsG9EVByaUrDWQPfuGMjXi0NNB7HL02Jts1
ET39WavAvKgcD32kLAx6Afl239cvv9bEVeMpOPdpMu3UCx4OAvkXokJ5uo6h5TgN
oyii4NUv0tm60Xb4La5bSZ+Zb6EiB+uaXVUIvcJ0eM3fSZqBg9FbtSLPTg5K2sjA
4llZAUnY6Oo3N4IXtCRkheUnTGos2m5PXmL7ghwymbPTdnbNjMsdahpFEw1jSkS8
gKASkB2NQqx9JtDptEMRStudzKxr7iv1EyS3p9SpoxNqXCwsLm5VUKr1tA5TFdRS
6rWlAAfB+1u2YaW1RQ1Bjumyp9HR3+wNMG94xHoIlizBDFgidlMMUmVZM7JEWTaK
dw+LRoIlf/iP/NptrWXfKLct8e7xweRc/JWqyRjzxyWivw73X4roYotuCtKaFdWI
F8ltofXujS3LrG5cIC1z8bzOJ4GziVInc1FTsSNCGlK3bFjn+ZeUgieZ0nPXGH03
nPV9uf2VbeuPioLNhTrrc56md1w2Pt9t1V9lpkIuTr5F1qCkq6oWEvR+ES6xw0rG
YgZQgYr5RqDJVTgfLJLRc2C44MAwrj0/0jHQLd3k4yVtMWtCVHmxnWNWNEUbHAWF
v052j/DBFeJy+PCIRRpCmqEFTbLH7NHF5iXIYbzhTdM8k3xhosH3+tDRPcKDydWU
vluWHPATArMPjHVfB0NC/Outh/GY7jKOTidaAQCXx0e5KwhIhoJDYpbvjXMbS0ER
VY7CsF9a/X9FhGV7davHtLBCSBb74XwVh61JSHSh/FtrrG8zN4XpRhHZ0FsII4MJ
IU35uU6zl6cKyPUCpONYv8s+ssjDFiavEKZodFpww64vTtNHklC6twMhOYcuGKxE
W/bPxfP4aEhE1VX80Ht7nTkptN0WC40r2uphSgHym7vV5+dzpmVSiUT/+CYojXcZ
eV6+cEyXpxdTEXnouVukv6qnYsyii3wsy73cKynJYvi41qrZdADkcpc3Pl00hV0E
npfQgzCLe6S1k+CbwNSA0ti/9j3uqMEpvRDJxkl/uOa2trWVaFKz2WRQ4nJwD1GD
p5JYA1X70NfrQvst/dSReDCQwee7Z5vT/H3g3rePrGsR6aKRI2WMSNqvpAn8HxD0
NUYhVaFPKShQxwdg9586RTdGoWlSoKwBrMlfu9OSt84RPYCdB9x4pBd0QSWZgJaI
DfbK5BYvChsYMl5DInQDhFYuVwIHuvuaYR1pWuA9ZGzcVYF8OMIbZ6O+FKV1CakX
gf8Aim/n39+d740Z7IV7l0sGb9ZWzQ1NjGa87BkmnZl76M40qZj48Jyl34QdG43D
jStQwvSWX9QZU0OxdQlfKHFmQ24fnEV/ltFIkn5sS3N4iUo3jzUkBTNr9Qc1+ufk
aQq84t4YI0/Cg0a4F7LEZSsQGb8BVgMrGqEE4Vxg3Lx1ucAoWrw0ySAG5ds+Owr/
ccP71EX7hreBpgq0rFxoBYnBP/lX9ffK7s98rOPrY++TiRVW282tBk0PcpVfAf3Z
qML6yYz1CpLs6emH0qzL5G33NxB47qKb2PX2v+kXAOzyBfArjEKpop7rFjxajxEo
E7wXB3v4x2Rr7o5VRWHl4PEEExngVhiyj3LpPEiUdgu7jDJpylXMs6vXamGxkdYC
XnvWo7jwUkP4IqJc1W7rOFJTKeG80Bc3k6xKvy5UImXyu4gyRdYgbyyowCzTCFrl
gGvD/2yFWAI9wctAbUSZXzUPf/uAJsWACePsRYk6JZmZBUsHNo5yIPnHNPsYnSrO
MKB5DNOpmA6gWAiJIAk2WFkAKpeCnC1UnICSCCrGV7iPF9K0m6jvFoKWh5tPpPUf
6UNegCC1G1gUzxO677g9WNMUkFsRaasRHRdMY+AhDauO1xAiSiwNvL14rWwoTGUD
FQCgjzRyAEilXRa+4crUXq7zyyINsn0a7L60jzGSYbU3xRLDP9Aa+GUzE8GSKOc3
0/dK0laDB06BULdRRQnGmzHNGPBFDExIgrGO06rgf8o8ku3CElt76yMy8z5FPD4h
l4IqP8HzXBsMmmjdfoIdF+uUfxkdkVlc4zJdoHzePBvckxC1K1P/B3rp4sgS4iBM
qyn7kfiz6lWnrizzqcCMrLpnIahvun+Dq5JBtRvQcUE3umNk0i5b1fRY74FL1ldR
pa+PFMtgIMpvAvB+LuSM3Dm3WGLwo/KYAwzONX7ht/1kglTp5oiL/uM2pm7/NUA6
W2p6cqC6hC5ry0fG7w8ElQkeQtnh2cVZZ9gwjwiV9Iqkhe93Imvm85gjHJ1/Yz9S
IZOb9QwSEEM15k51pJdEpAlbZpfloDItZnJJD9r3Dr0WYWZQ5DDu1L23K3oDWa2D
iCxynLvKQC0XC6I+XMdLcpyB/vXr8QQFm9Se48ocjfTfUU6jGVg9PtNHngFqkT+4
SNp6Nq90VXoC0otBvk7ts26QpyA50HjEcUHaw1+/csu3BbzWFE22mMKdzQGUe5lw
ZC/FqTQGdp9zbrXVAv09h136HpjWtfkrcmkcmyjDLJXxf/ib71f/txg1f2M2DgUb
Gtle6ZZk3r5DLHU3DkZxOjV3yEMOwxZ72IxGLGAVTq4+qq1xhjGDak7uTAt0FBy3
vzIDsVZErc3dbsZPozGNBEcjvlv/Au34s8bQVyGL3vr1yDcSWpKQx4Hb8FTeagb7
l3N7kaQBAdFg0crvqeTKZbla/+GQtbRCuQYCTXPTG9boPZaV1rbnkfvooouuFoET
RegR+9hbgPxi9O4Wl3Bfh0aIKvCg6/t7SU6m2Rq5scqVNvS9dBCHdkw6ofmtG2qR
h8x71WPvK4X59a8WscUMS3wHSfLqMEoUYwBsE2beTIHENZv4J88ucJzfc+akOIgg
HVFJmzu/0+i8cMsT4aidoNLnzZuKoph1Tkr5l7YEo8k/QduFadsJ9pNojyd2e9Q0
lsH2BBN7mWjrcd9tlPzY3T4/xm1Q3GeJwWwcz6bcekBPy+IU1Matt5hJbiA1JoKi
hxaGFe2fJQWNX+3vOv28IvirVnhrBgbBLZkqTC+WQ+bfjYkpwS8RhBfBhCjY7CZr
/PbdhIdf/2A8P712omRfQgb6EuRDDfB+oek0fq0FoZR7gw5Gxezx9LxD3QMbEoau
zrpuBB8Nc+MhEARHrV9BEE/8r9JwQEDrJFRPpBH/rJcDE/69V4VPqSCGN5ejlXBM
JxxcepqyLUiFeEyEFyd8f4SrTk1tlhmgH6bVnB3/t5Bq2o/3GoLzUGcnacbh276z
Yj/RNMFwtxATKyqFyrwOzO7gI632QqOZGazPQWHJq+kSxWr76SzBK6dzZDGAq1zK
g999SyhdQlC2O2r/DBADS1rN+XlA/+aJOiGax6eLeck6MxrND7S+pkBmtxyntD+H
L9LMcTKTcE+XgW/GRx5Wl/OJ3iXF8d+VZAB8WdScMWvulrr5YO7Uhj3hcMixr49a
c9MV70MLuLVtO/u09oHvOapWxC5UqzqLU+rndJt/EHwW27DM+wfTR8OdXc7TNFNe
117XUX5FYE5jt7QMFONaZM45kaZ4uYIhswHsc3ITp3rRhTH7vNqbmClL5SDJHOCN
L/aBiN/Fq7FZ1dq1xVbTS8VijAdtf1AxByrqNR/vSzPgiyVa7QLA0IsiScz/63EE
8ieZkn6FjR1r11zT+eoUjC5uaNkPtS2EHSE1cgzLeFfRRtY8oH0sVy7C1Rmsiyxn
un0MaDX3BH+xzKXYCqM9PY+WAW9hkqO06lSbIEi+dFLeNRsLAymYt2eVtiBm1BHO
ED3Lebvt6kpPctAX6Alic7SYU9DoIv5CW98M8mtJgUr6TbtOVDnu3MtUcigstGQc
GD0+7Ez8UvrbtsugIkbeMjMuXg8FBiWYqFrV13zprIxsx+cwB5UgdMNEWnYFtl1f
JPY3TJ7R9Kqf3bSj4l10IZlKKuQa9y98xz6yZfmhE4S01P0gPG4+vDrnhU2CeS9y
763pzKWYxDCduAUJ5ymBykhT24QZDiL2Mi64nFwwqX+usbc8P3hNDN+e/HgjceEH
PJWfAbiAkBfexJQFf5CInrrHdDIr3FubkzPhIJNpubSXoekNMUuZcjkb+A2P9JJM
NCSqPT9iBMZ0RTrDsg6TnxxCoRP9EmEIjgaxZI/Hokzl5s0/wZVcZFMoZlsoFx9G
yfFXiqbgEITFAvZnoVIytH6dEQcqZLS8dzkorwWn3QKufg1qc1l7vJh9AkyBEQgW
L/L4qndqibICvP/gmXdu9OBLHxiHEQfMau3SJtak42hNLTLwdBTWGf5hikQZIdc4
dUVakEhSll4JZleLdbyMfN+gfl9QcQ5EC1PFbVsRFHkIG5cXr6YG5fc6GJ4DDTf9
obv2zRAE8z4bft1bpxCEsmNVfvO16UWJEK76Bg2kSjY1jHU/rdDgy7+qS/KU4ByR
t8ssHmu4HNPewhvkAQXmCF9gyjwiwBA3nLChginMtGH+ZWN0NZb7fgCifzI4wG1m
+VYjdyjeSdHH3HQT0kiAxO+H+T8InBJsczba7Da8Esshun4H1DiLSGoH9MiPe9sT
cEqCWB33hTtoshgL6VxIht73gq+Hnw+XjWxzwehlTgE+IjjVxH7ApY8jAbcvPiMJ
6u7UjLly0T8WYXU1EGiRGFF1uvnec1Z+/JNcdhf3YyHqSqcgjdGBsyYj4O9IQdhS
mSzW2e9ELHlKDFAEQlP+QGA1JC/UpazLbHkPt635Twk22/v9yYe5ZlmioZk1Jomt
ngv6z8k/RfRVR7n+rv+V0VJdOlgFiz0EbE8sjKOO6Qpd0ZndX9MH4AG0q9HPFmYt
WzhAegqyjunBuzJwyM6CTtO4E3Kcol1ZrXmnAaZiARozLxIPbPUzFt2hbQiDvuzp
i9v6Pu651wCNhTQDyXfYSN0JsE81hCOhRgvPIXH/FEjGWnR2BwlNsN6CFKdO8WUv
vBvLwOmU7cQUNS8gw/dWhXIACdjpCFJ3d+XfOfptjihJp+a1/5yF3D6nvInjChfk
l3Z2zIAvoJrxsKE9sBsV9B3tL3lpoTe63yDpstGXCRxnTWs2t6EyVJ7+VfvSiC93
nIDmoON2vX0JS4weHQdXOyw6fS9i1pDRnGNNXAm113+39jx/eAtxj4iVNJDOFxOq
2UAt/iDq2y4UDKTiVBnoUh4E6uBBGjoUQW4sU333J4sE3S1ySmdrKIy5y797YzZ7
B1H+nv6EjVmRwpDc8p7y3mLi0vDCIfubCNKpRLNaJIr2SO8EcAutBhcE0oQ8H6fL
GplbMQOVaTULHuOTzwVdoFUWZtjU1yB0biTzIA7/SrTM3ELKURPOUBNHDm4wnTQ9
1UwbjCcZPJtWDr72g+me398tBPEkL3OMFPcC8T20U3bQFJmVex9IxLtOfoLZPQ8j
LYHbWquX1HIFKdWnsuK8SdR9gCNi7//Mv95dM3dj9spC/DZNb1Ng0CzhNqwzCCqS
N+INOnotB1BmK8o7kbkamXZP77uXaplC/OfBQRY7k++hzkmFEVV7GOQJ9T043HD4
QS2MoHEUqF+Q8z6NOhQ0Do5yJaXHwSaCkh7AYdXPb0vvrBubhCnEr/UPr1JSC8Ql
VLrSC3Y8GZyaXqDBz+uO2PYz7Xub7hx4BP8vJ3WH/L2tIeLFT6JG9PXSRZ/XM/mh
mbIOINgR6ckKAltzUFr/Uy+pLDmW3hLaHYH0DC8ilKmc0A7Lw3nkcTf3MfPXXIr4
el9uV0YnJB7ZcM6DvUmEWsXa/8rOxm/MXj1h6EIg6gjFcEWQv+JgvT/81CrhqZSi
n17q2FRsFda9leLsidO9/jW9SLHCwFH2kN2fa4BOLpoBb7bMpDpH9XNilI44XtO6
KEp3AtHtrjeoFbuNFV+YS+BASXGwjXHdLcbsdtFANvdPPTaGLs5pa/TWt84SQ+jK
U0qM1ljpuVkByoSmc6gk9j6fHqwAdxQsJX7IOGv5qdV/hfsflab04tQniuJyt6S/
7nt7siW5to2coI6SYmeJWVfT/sZcgdpmdYAwdZ1dqM5ey++6IDKQIxqXALhziSaL
dYKyLjVsXcAV74wAjA944vP9wmY5/zpquehyOPohYjMLekEi1pprxVJ2eRJUlmtG
VsGdbo4bme93Tdi29TmDOXXvPcG2fQpKofl5W7ev8FSbUPmr0BjaP44Xhkx2AXuF
6pNImdWb66XKgQpuHARgi8Z7/Ij83SrlUuHSAR7hbtMKTWzBUSgj+qfcM5rZGsVp
+EP5Ih5/e3qbYkNBfTmAAKPH8yRcM//7TvO5YuOVh0JIdF/ZL3eJ8bUhMY8kytgp
RRl69fOPw6xFxKoE9qHuvkE88TK3VhBvHU1kOu9SkuQAEg9SQxK938DWR7tUUmDs
utKRSxoO+/mILEAOVTHS/351BEUaVgvuvmO+U8wBRr0snebo+oYgoIS0OcNWQr8U
L9aDKlhtXS6rmywoPFhA7idK3nQaM8XjdnpZ6JMMz0q1dgVIU9VcUHVWVMnizZpb
wFeiptGk6QfL4p82c7rqn5r4Y7BHKF/8OBMIoMFmCDjSU/czYejpkX0bD6FaUX8K
t7rXy13jdpyG29LDZx8zedAvvaqFunlAN4GzmXRYzp2Qje0INh9bu2xgSkHET5dY
vgg+ShKeDNFfrFlPI7LLN4oG4tDzatAJDjMeWXo6MyBBdu2lnQh0D0ZAj4MaW2a2
hRLC2dTPEX7TpqOdt+0xr+MSWIiS3A9iNJgKqz/a4zph6ULvep042Ps3WOhMUhx3
dQiMtRWhdJZrv9Kd034Y8hdTvmdEQQ3KB35cRV2ffw/Lg4IY+L6ddJgCCaKLOYzM
p/lIq/QtO2sBKNHY89mbp519ZtuhQjKh4Lzfult0lYBYkwlULms77SEKLpjloG8I
/bgGpCh3xFVJO0JdWHs+fxueJLmQuYtSc0GtYdEPq0Xr+zplp/zomuRkmuCqCQLx
NrRP1IFdrenCRm7PP5v5g2CwYCgljjlYfj9UOyKu2lv6e2JHxAibCgkBMVJbhZBW
x+OjNTATbgmGGazauC06e+fgl32qHoXfGuP3R1VL8qczwsUmO7M7yp3W35Ri7bjH
qMGfQlE96vgFfLBoaGBV8L/qKX5jjWho48VFB6iTez2kJSUwVmi247A8+ZA5eo9Z
ZhAwp7PzCWtbXnXmuXmleYtw1hcUywrwichm3+KcMB0tLQot/7Aj2O9U4TAnU+p4
0Jhfl8Ba1gcARk4LrfqizLAIdQGNkTM/kiAL+0Xi7eHAuLjEdQKDuahlt6StBKGF
UIwK9EU+aWjVftjV6tRKq045K/7D4DsSqXnFyPUNL7ZhH6iewRvC+w3dEfC2LyTG
5pxKUDHhmnZmg190m2nrHQcs1YivacT4hIe2oZoX8FAXbl9w461k1s09kKDugo+3
YxoaLByrBlrk3MOppsO8ScDhZfhzfxfka7U5rvB+exld0+PHpnlARx/3aju/dR/5
w6GSewwssF01zTfX82ULzhiEcT8WUuyV6A8CXI9XN7PyBhAWgmMvi93iHUpDIdIQ
fPbyYxHYYWDH3QZmmgthBjr9E2XZQimnlV96typKvc17CiV+To1qsxy/BnRaYMDe
KHN4MH0syt23GvkjkoRWrzhsISy4wY7UnjeOiUmW6vmpl6RvGspu4cBxKK78mIz3
yHK/oZYAA3r6R6NDBim2vvberFIf7+BAjKZJf6iZuRDyzoeleI3gW+9u/hKlG/l1
kRQiuG6dLsGy3Y/XqrvoFvXee+zztE/St7FU0gItSw6Ilz3E4Bqut9hsT3yq+RIZ
Q9XKFxKoyw+4cuwiDdxEMasjJr82pg7PBswuLGGf2Lm+aNpnwh1FvGn3GRtcAnHM
9DTspS68ZI3pVygsqMlbPhGEr54Y92/O37EKnUMivnwPzEE2ZRTfs66AhOZSCdvt
MSo0BkEn5Bxmmfb8Uv1J35sme9L3fdlWkA4YVp+WoB18IQJRwot4FtbOU43tTv8X
fiHbuUP5sgNGBPTjMvvCD7NHXU/YnNXwgXu1jIb1wqwmDDKPafCPmQIkZElBSyyJ
9DSEVZMWG51/1MtLoF9rbN2dG7KRQ88999+Nff1u/d5hw7GoJdnYj5wnlHh2T38+
SNKsOV7m+T28AFtDpUtVTI+uvLPmu2pivrl9xC1evRGN5EeUnf3YtPqyDT+M6MoK
ZhG4CkHt3fa5EObvDvteddoDc6MfB+jyyh9bbm7yYkVvTEduukcakY143GJS1zRP
M3R/HCHGv3GS53TznP1UrOkhfbkO2qXHMUMzYTu97cwEtIDaCeNxGsvlp0KGak7N
+fx+GfBZ+zPn7LiuMvgH3qV9EfGQq+zYtemuYp1yRmHgyGE4B9Bf8ZPKP24FgwD/
cgjpbjL4yBeAHZ0+n5OIw/oZ0uIHIoB7nsgbczMj7v0ytN+QjBwIJSP8D9pHseP3
9C9TzOWVchuvmZHQXd5do5yMEyh4cg2m70wD12KquFFiAmkZkYEsjeY6psmywlpA
ENtJ8maYmpr9FAwNx2lmBm8pMRXxbX0AJFyF8NgUn4R/OeHgvIJ/IXWXQeOcLxRM
BVF/fnhkO6jkC6CFEAbeZWw3Saao7F8ZT4xo7ltwOyYD236Kr6Fmn7aVM5siwlDN
oFxIFf/LqwL5wI6NqHRXNY2YPtO62jFJ9fNLOXTckYdpyS+99SxrmGDMT7mljy0z
FsKJ403jqwRPswca6idcD+gIrLgdXWFF4ykpBnIcK0Ga6er587THQo9vGErweAJs
CeJWgXasP61zwignaBYzgxatdc+WJqZCXxvkDikyf6OwUw24+RycreIbeTXxblGB
e9fj+WGz1yG8R06aZPLyCAqqp1RVcdiAqCKCqiw4U+CXirDA8/0xY1Us68AC4e4X
dt6hNp8/idEreDwt7ABe2m+9dRaPYYfJpz+lvIebQv8O1g0pMhWY7qVvI8zoKuLL
02yrXWYHXh/pMRu6ltv7+fFk2vPkOWuw9zhRjhkSEx/KR7wgjMIQIKZC03EY2lqd
IbjHWSFOzqQJhzvrU9h9yr/1rNu2hEAeJ3Cy9U9nun/6uKntT2t7KtHAkigI7ljk
3yE7jCB96DMSNJnZqc0M/cqKpIsjbhN8WlHt52T1JyZXmpJU7xz8vG/Wir4IG5AK
feZaHlLy9hJ7I+fjlr5POaR6FhSiAWjD/BrSdFfx1Y1t4zwv82EZ9QoLu2PJnuWO
LnCbTZxbCzSsZZaONFazG5ZeNqsGUfbO1ISZCkemX0yQOAPmCuRmOVh8EttojQSt
fPgB3Jh4TyY8PkkH/Nc39l2u7+nUCT7RbTb5aT0Foddmki+ViSMxCU3INDesrS+0
yGcGnbefez2c4wd50VJkRjw0H8h5zHi61+Sd3yVCvWliUy2uSKX2n7lUTOwYViZ5
m5XEWamfjk5MOdEEbvcr8Q5dp/1lFPlTdSqHmkyn2xKl6+9kRXwUZieLqd4BmzCY
8a09zKnB31YKbMMDxlFoAATcuM/zCacZTTS2EDls+tokwHER9P6RAeoSX45G7ilb
JwAvsBt2rb22iLNKCoxz5kjA4ahnwEXoe0N2ETH1b8+bvybWlOf5/lvupaiBV4+r
9ZEpprypspbel0r9jxJAMcReYWKoqgBPOd0QPKm+Nvv4r6rQLDeLl8f+3jh2pMw9
2eN5L/ptHuTRVxgHKgKuRX7KYLAa0iwU+mt7gIcdLABucLt9HNjuQQ59Pw7SkKrN
g5uOogSNGyMe2DCxr4PSmGvBRypcGHKr2kD0GTMqZOoYIoYviieKtG6UtTv2/5ak
yuNCpIkRLJszRB1Wx5IVION/S2pSz44QaXdfGSOOk8iwl8ICxARMP2fvhULIWbSH
8Feqreeq1LThlYZItSMse0Mnpj+wOjD2CqNxmXCUlrFmqzkwwl8UKDzhNhIsC3rI
HBkV7i6FaVWJcZFn8wlhVOh/bhBd7ylK2BZFwCqtKvtRp9iZyWOyQ381CTevB6qW
Zor1o9l9YQ7jtQ6R3rTlgiC1uFfvLhJiraF7W0WjMcaKkW3YPUmTqXpQ/DHMbgFz
Y8Ap2/ViGFUORTg/s/XmWf4k3iNpwyVDRRxSdjogXlpHNqcVzfvC+Ye+VXwKBIHu
6IuNQnxrrng7j/6DCfwvL7xJXgJNgeGqk6olmn+vhAumOPF+zUa9BXnDqbFrN5oX
/M+jSW6jgtjODKwG13eTX75i/Sq6uxp/wPgSa5QnKTUAlYRDtpXZEkP5z1hetJaU
3tGYRf+VZwTMXhfSm5qKurZISpsTV+1U5XWLsg6peYcyhFHITyUfJ2ZU0x8ia2+u
rwEQxAQMxKKJGzq5/surFtN2yNxbbxYAyyowIeESwwDkoJQD1CuCluYAUXkpfBsI
1BDYSnuN3cS0UH6ZOEY4MmkCS+5h+c+b3Ipsma2zI0ZmbuAWkupUPZk1ImZ9+pAy
ZLPkOPFtAntowavxxH9U6/dnPNxwOLAQ91RLB24jC7PdSJD7+dx7piVzuyqFW8Je
z6ZniGMvqg9wug9QNcKJjbKQ4EUvZIEsh+OXEf6DzTOjRX7sVRGwOSRSQOgZiYRx
59bfAVIdJIlddXgdhq08JKzeBbfu3r/Psu4v6MGMonn7Dq9DzZYPnL06rYNglJgl
vCQnLjxNYGio+0xCDvbn18Ik1rALWtQ+xgzm69DQHQz0Rz65ssm7FWxYUOg99y5w
zQT0ekIyaWfnoFukLmOb3R633yvmSGylTsEH3A75WwzIWMW3dy40iKKp3phvXvkI
6KQrI79umjNzmkj+ImdOj34jwExaQHqRjsFRCzGJReu6gKGKq+XPcIskVd/4jD99
lrkXF0ztae/FAjFdLT400/c67/3DCYellbc+OIZhpO+HYmgoPGrEVIJTzxLJEDu1
ZGrYNUAucrUoltBfrfzlqKl/7pCeVFcmAyM70dk4i0QZO7MsVNqzPQ9f5kbZ/bB6
9IQG+IjtiQuelY8Kwawriuh+8Kw072tyiCA1whME78L/83CKj42NHIC6QR4DMidA
nb2cr44xhnNAgbFUpakJdXHFKf7/vWt9gyrT6OEzdKUIzjjwRDGi1qF9kqUd/vEJ
LNKpZnaebzmZXXPLJmYdKg1bICMKWYMeQ5TT+WjkOhCPyfaga7zDQ5zgjmqNBgSh
ujxNs0ClKd0puxHkEwr+QFyKSf6LuEmavTH3V87q1v2q2cheZdKEXhasItY86TIC
pPqjsMNUniV/4dbXtOQVsz8qJgCoMHWxb2xPHeamiQg8NG6iKQO2fwg1Ql0op1kg
gpByIwV7wLpSwAfsQHOI5p/7y1+T9U/P1i0+PIGmjD0zrOuf2ZAA/DS3XqDel/Ou
xHdP0QRhRKoHzQsmVqyQQz1/jIFdSRB6q5yxgr3kW99D84WxW4iY2tfLxMfYBlNA
bt8BIR8+wsNvJhkuuXcaSgMrymMuSahm9PA8/33eBqTjl+tdpa46/mwzo44YwMsb
cW7Y5FykE8kPzc0mOjRpboWD+5SnwLTHrb4K1saZX476d6NC80Xbw8ZvFhVgPxml
MH8ILmRV0BE5XBH2t8WB5wgXTn7T5ajyZ7zSFhnxJZdUo8CHDVjC4DNpqsx8uRQ2
xUq1eTP3Avvi9lJSsb2p+tC25AOOwBDWB1m20PZdx1gluLb8aPkji0FG2h1MfHSW
veaGMU7zijdkfQBXU2yCy1YkaOuGAPdw5fHDTgKRKltDop3sL3sKpqfz/5QDjuPG
yCDS7tSSx5EX9j4E6jv0OsgntBVI03mzSR0CmplYnlkcs2MBsg8menWEDFolHft8
nNIu+NDkLbzFuofrUIoH/GZ0dj4ThnYeH8KRB+P9QfJPuilkgMtNcOy2QNvROqQX
d3qvFv6yzKjIdNTJOQv233taWBbc6kE/eS9bZkHNKgsrh8dyl+iiMZS+zL1EZxl8
XUGt4zyBK5FSGnAXVapsmi3tnTs5WquB5h+n3x6eW2ed2TnyyOQRodg2BkjFr1k+
Bt0LoZv7r3/p043jJEmf0n4oCopQ6cfd27rZF52iEckdJFrEqfqWD94lcUp45LRT
N0wiVfvp5xgmMFy7EbXwPJxsQbEL+b3RQMPmLVbQ7yS1VykwcJSPl0JLKNFlFqiR
6R/ULcdbeI2pOadt3M4rm1rgqbD5bioC7fspnO3YmrjC3dPxE8h82EM1SOYcBS4j
BjmoY/oQruYBb9F8PDJuc6FYHTCel3O9o6qKHzNWRTvlHSbbQmzrM2AmN97fZSY3
7/8R9whDlytF4O3lsfisUT9gmEksSc6TJrpqqCKp3UfHAbb866BXf+N1ElexBo29
/T+llIIctdObjFgjdHQjweCe7/Ub288D+vA4L3cM72WFpA6mEUZMvgIMOdUalI76
FGqBoCVDBMkVY5lDCeXgRhWy4TwHsj4LzhbK1buBm4sWwFoIXtO38jOw5snXhKy1
/zRGbl2m3R+tH/hMd9miRe5oNm9TjQ1ujQPK25Z7pvvfrseQFSTiNG2vC3Zf19Q6
bvIVIFP06t80PwIDNg744IE8mtZpGvLKXRR7hKI8cIRFPavKtjy40o6Y4NaPI1NY
n67aS6kA938phuLd5ICfCODzRliVa4pSYl1goUEpn3Vm7wePWZhyy4LqDAW5oJee
hmaNsfGBuRh9VsbONMnzzfQHg7ex9JlMmBogmqTNXe7BL7fjVdT/gPIBvKG/8lto
aOyWQV8m/3XbG87B2Fg/6WjmNxz4GyKMB+DOn9YhzkmSBBPbiyLvRgky4a06ipCs
bf/GekQ0KAHcFVcMPNShQ7nLiYK9boH4/4xpm/Y1cKGhq6R7W7G1WrQGKBYt4R6N
xjWJVDfJtsA//k+ndQra1VudiXFyU3ZLYTE6yM4t2Ap1FSjwGxrcVRZJeebbtTph
bIImtf96UwheKGvncFkgBvu35fSpmeqs0TjuZH5mITR42lPqcQ91R6dXlqFT8Emh
V8uj4Te8dZxe3AXHtb6BeFW3+bUWLhF8xzvH5wZSlcVjOLgIvzO8JE+sO2f+3wmF
ClFMQLR+Mv4Ghy2d2QDPQOCmSnNMGw60zrieMswO4he4sq+MuvQjBlViXCuTyVlV
HlLau3YOO43s14gbvGOsS1LmmkM3Q7mWOcgCyqedG7rFaTyAfMiwGFwwVghKKFZg
m0q/1UPouZ15eaKzc8uZ2jBwWqns6NziTgBBwq1JkY/7hxvF8wC+oglTf+8rAgje
wRf3GxWDghq6N30rFpJjGEybLprhG54h0cU6xEZWFQxBrU1pt871OSmrH8qSZUFn
eTcgnrm1RWL+F/WqqlSGzU4TKaIVtp9K8qVeSCnSjkKQ13TuWGlhx60xhbMgkmgf
g74/VJpOr1Ddvn50lybRRf46yOKoIXhOVU5y/1lFQX6KvyZubyw/eCFnCvWYzHLT
wNPymVEYBxbLCtFT3NE08nnssiawMIc2aCCWdt6Ju9aMbsxyiZZt/J6dDKKkfS4m
XRneAfK7jEqA3C6nunSJTXccl3aiPxwa+qvvjOEfNdIyiLnvCL8/RLC/x4sM1LzK
XrN/kuGaGZGn65kNPoZTcxQhIp5W96OMpCeqFRyc/Lt1ceeIxi2B0D2gIUml9qxZ
PlwT1/iLRH72Vrg0BFcijVt9Ez5C7WcDNgUtZdzVm0Sj0rxAxpHZN2nIccSo5ta7
L1FwSEQLnhDeo1GnwjG3n7guaVNXqht4M/l8KDXJ0oPRdNHpVTJWMavfzX6qPVyC
TLJ1Z/64jd3N+EYvSN+LqAZcLBFEH8OAk2IWKpepOATv9Dy2WUudMLN2CfxYLXT8
1cT+M3Lw7pO59p4KN39AEbHhEeHAAS/AHRtBmmcJq9AIWENkx3eiY9npbk2KmQV3
z+ag9FUYMlsz6Ypx42xMOMISc5ZpcFlU+3HPe5RbSYMUQX16qI0e00JjNwK+4v2y
SMvcxU7cTihcPIPBcB7ELo9DGV+WinoGmrEck7DQjCjUNVy1pLfzkKXFxdbyJ2xH
l3wTiKTTEV518gM0UEd95zc2v8QJCr4a/bhLoxeKzUUnQLnCxpEkWoZP6J7XIRBy
o8nLAxeFl0q96PgWwtqs7cvIQCFcRkRQoR0XvkZCiR2eXDL6o5WEGCqMNUA780tF
r+36TXQ/L1lG9+1Sbl95cfsmeFOMjZkyl/lxeoghxuE8nye95HvsPLiA0Jd85GJE
+02qVVHryzLckCVkyKIyA/HZYGPpaZJmHhVwniKEhacWs54LxvDEaN2V3fr6E/QB
xO/oGOqj0J0tGkAJygelf+WXR5cyBKejyiYvFicM/AOeMyUxV4rT/nY67uMGsY7o
Jb9YPsNHsO/XK+XFjTH2xhRBzCzvSE+OzjYentBjH5bnGTnWggEvFJbcVgpYzK6i
hb0RVczKcWnLa4AfwPVxOmqYNnDFAqVQclX3XrRZQGdBIXdAYDbUVkqFzsGxGOOS
yhFwIP9jnmeNvptxiGy/hiCuIWGeFI3rSh1hQUmO7oiq6Axx/o5s/x2HT61Rl1Sj
W0YnbVcRXzk3anizgxLdyhSmvlIHGZrMHIWapAWp66y05Td58xL6LXemk8xw/pba
QX32gObqtn6SaV5mrZ/kESB0w80iuz62KZJJsRdx5zRoMasCW8npxHoBF12l9KzD
jTHE8cD8sHzdbvydV3gS3KHj3sYLzPhlb3dsXAIVUtlIfG3Lagc3mziGCXH0Z94Q
shQ4lRwL2B2CZRsO1CLdvZLaSVbNZzKSIW8vG24SMDT377QBhW+AV5XDFtB3xc1L
tS+7iaEh7IOiiNN8IwfxXCamnAoSQP/P0H4klQ32Vljb2c8eKe/NJWwkdSeB14qT
W2XhEZvo6ZsTwZnNqIxzY5nGP1mcjeG3XfeSY7iAIBenpm5WWnMv0baZGJvvjcmE
s2jLCI/CCECUB8+zUxxu/b26gQulV4IaljBIhSp+ks39PtTwg31NfUgdxsmb2Kzg
lgjjArezhPgJeyfTyIxhbX9P4P4swBEWHM1LDlFPOr32lHHn3CX+PiAN75XTe1SV
t0/TvzQfdw3fhwmte71G7FAhAyV/SgJhlVTEe+wlcz3qY1H2daeaDAWHPtmB4HGp
/CGfjuczyrLGdlfNooEsCyTqJ0V06d/V5jnVGwCicpXLJQuoiQ140HgaQe/8Sb0m
viRRm1j7J+s2G3LalLBDt5tWXxFjaJndm7e9hBP6OfNVcEWI6/l1GnFkP6X6QFL8
dWk+Y0fRjjrfNr+0U7ixmiBSzkxuNS5Izp3uVgJniMlA9LY83iyIuvnNRrcZ+UJC
H190VB2Wxng1Su9qhQQnXhA3IrWaoeCtg3ZJ8tSa0FAxHuD0K87C4oCgGLmcLYZq
34E/3KqHuRvxyl1mcENIXp8aOUi6BHfeb/dLWoLF29aouB7mInzxJmzYHPbipjoq
TU7fsmSwfhYjzCGDCDvtgbILeiAC9wREE2Ld2EGlEDfihSxGfbqU2hyKGGdTMU8g
CgzzysAN+m3eBlF5NygbQN3wS8iy5W4uMnFdzxZauw/+vyAjpQgKvpYjX693FDm/
fVuMarFJUOEnqM8qDBJH/skAYpGGOClNkpw/+gt2o5kmTz9L2x85yuKEDqn27Vhv
gYZkq3d9+4QMF2IXbOE6dsZIUZYg+ywsj7aOiny1Jy6kmX84v3oZkDmz9XDD9GKR
1HTmS1jxjFryZEitUwzpJXG5YelJB3bUxVwj0DCKz3Z3wpFn7r76evWMyw7W0jj8
2ZMzK6twAiF+vLhZqm0yX8gT/QqIg53uHt8Q0TiNXKofGN3ZqG7qY5pqb7LpDlEP
a+ulO/HPsxMDCkiMh4eNa0vqyiGmPuUVi2pf+V8qG8eFZzBWZTI5vqXX0mPDsiAE
g7s5hFO9osbgiudfog3PFQQ9HmCGBWRSkDrGbM3cXwO43gaGS/W9L8EULfyr7t4t
9+hNUzVcDRvptAj+kqheH13yjUTOsNlVE7tavP34CsVPA853PeawCQE5RYGeHvnH
3Fv/AHWUeMUPuaLvAdvZtX1mBrAixzpWJnjY7Bb0VWekqDo/MPh7hKNrvaXp7HF1
Y7EnUa0miRShShRdOpZ1dEpiUDPZb+j+JcO+H0U5dcmsPlh0fA1mlFgzZIJ0I2ib
GahrDu4mMtikT5knd+1h5GNQPO17pxqu9BSBcwXdIVzlhMy3XQlSJnJ8UGTRcSn+
fl2hPLjeWvF7bEIf/fb5OCuh90K0MuFMwx+1tkTJisCyl/F8mpXQTQM3ATJdr0FR
m3ioI0tQdP2XArbGapZ3TlPy2cq94d8KDaFrY+fic89kA0V3miuAAqtDC6kYUUHB
cigefwfL78ZCygMxrcyyajL56oFef4Rq60e06eL22Zub23Sq9OmnPFIWrb+vVjrG
ZqHsHc0PlBygfz9tFuFTnUXO8265cGqWxLSRgyZEzKtWrMglFmY94+tvddfo59vf
faZbqUj0IJwq/vAT57kmYfjbGRvGD77bK2cq1D0nZLJhlS0a6nGb2y7NZ+OlVgTS
XF8x/eBAgrCiUz9aAbfKCTEqNYRMBnkUhbyaOyZ2r0I5PS8gIyMwBoFPTBJ8pDgM
0K/DcaLKZ7SJk+4tSfV3hQycxNqZeWQdoFQzkQyexgYA/bVqOaLBhbGTX0cebvbP
ht3vReMirO1YBaMQxGP/bGQPhVjevxNun45uWJoStJpTuBQMHlaNVOToVCnwCPeq
qJS+g6/UT8Xsc+FE07r1OfNOgbA9xziOAtOFInWvn516o+cSR49Rz0XSEUpTEIeG
2Bq3ArXlKg53sYvfVvfeFFqdt1kALm2rgdAZ+I66sUQ7l0MJdVL6dY1hN3myyai4
zr3wKnTR0Rs09aoayfD3bI5v/58t+eaNVMNVAZly7xUh6RoPm/N3+r3U04etaQc4
8l0OpIafFjLCF9BS3IUetcg8+/l5eIW74ywOB0+t/tS7GK0Im+gPAtzqkqk9kHDE
MEXuPipDvHFZDndiCv36ufTGMzCFD2/uTOT6jd0E4u4X5Ax8hTdAY8EDRy4rblRd
/zfB55l7kNBDVT2chDXSFyia8qZXGdo/5RtHJt917VjN1yl5XfnLhzwApWkZ6ZqM
Trkfjro3Mt9TcsYtLQqL6ZpilODQY/6rV66PcS42nn0JaGCAOyh2SooFsMCzYAO4
BRy91fddlTYJkpylUVE3+bp4r6k8FeEZ22fqx+W8hu0PDX1N63nMca+U4I7rYpB0
YO/voiJ+ZKWeIxboxqIviZARiEVD+ObYJCtdkQa9d4ynxKip0bquWyBF7jdY6PMt
V/I6r/nVWxFiJESnq639X3CJXd0TZRIJsrKc6D6k7OzmVgSPKKSdMNwHFueo+cmr
zSqVMO4DTmvi5rplpPbDmqpNQ6xaNZq5lXnz8746tmPHs2kVraKh992vWd20C2eq
KlFKYfeUQsP8LZwHrYdZ2NPbIH6vy9VBixHWOoDcwq6zy1ZXpdt9F1q56WvC/Z/E
gvex8TtQ6BPwEup63CIQFgzeVuUOE0v8zU/E/hpDeGgcgumt8ZZDagENNp30OPsD
hhN7ib/Qi8TMvadwBxZZ7vLgcvdpaZCXvW3edA7GUOjH0nOH6y51iLZ1kTwgl/0X
7kgwR0J85vd4foXpD3hllBZNIOreqC7eubi1fmGREVcEWwLv+6nA7kIU2GbI4iQW
ngV7jqKannTtWr2GMOYfIa2rHKMchzV0skMWCbjrVlmaSy8y8slyf/dTYRamJMJS
L4B0aBr+q0zAVxs+X8ixR2T2jqF9gHUscHED9Q2tXmZu2UqF574/0F5xepv8YQ66
cCR0eEDMjgf4dNaMO6LEzXLk9lX5SImwjmTg/tTuyzU4708RMaKja5H3ABEeXxN0
3XYG6qdTP4U5vTOmSBQfZthY1o39avWsV3EUcsBKBt2RMAZu5IkcUd7qzYOu7B7c
E6qLzhDk02GZvXi3qyPjMf9MY3Pp6OTpzZpPBoqR7XwsN3bVLGmZWG9SK8qlL2Fk
GwFHCae5rX5CW+bvk81vASIfVjJC0YlsgM7yAUPH7AdY+pyqlbEO58L4+cFG5VFz
PsHbeBBwOyTDvCtvr2FN2eunl/ACWE8s320hO5ItlrCfMnxndSM8qa6/lkf59s9q
dk5/9rRV3HnJ/gua8wgJGi1UyOS09zf0fQKkmJ05vt1+UxOrdpggvLzJBcyWV5uY
EUZEog5mWwalsh8umjSo92wtgdwsYT6ygdBsQhf+2F2FeGmJYgjOx8ChMF5K74lV
jkpIenf644LCrk8yDvjaCf06dMHAHQgfPscOPXm+RobRgxiyDC98s4xSo9WvE5wk
t/mRoRz3ad5+yNUEP/dN0hxCSY0g/uLrFjnYxJBeqZNvb5FMzTltkJLu906J5vd8
1FIrfuJtzzbeHyUYHSQw+rmYPiQk9jGr9fZTROIIeT7vaTmP4d/A8A7xiK6UTV2g
AAjorrETSNg/tUMEzgO/pp6SNZQemG3ReCzrINyPNvcfUY9MKY90/ukUPHmIcBAk
K/SXv/xzYpf/tPLfmU+LVYsnp2zHHJmI22SGt4IPl+DkLY76kW0r0dJLOz+AFq8k
U/2WrOUKaWhXrwlKK3l3vsqbVTHvsO2BcjWZ/9/qMorBsPD/Ofe6bvEauW/U0lcN
VH6uofSpERmTHQnqtl/TOE2lpeT4JxMdUL1CmaBxvGMaKeHMsGpX81V3EyipP7oz
IVSQlC4hH9s5QkAZKSBwgYJEK19Edsg8PYYUomswppdGXHunCK0f9hBZT6Aexczk
iBpA5yeQrJxIc4eG7s9cfqw27VrWnLJeU2yWecJAaZja8c1va9zYBFP5CcbDfS/U
Svmhw7TjcbjjB8I3Yjc8w7GJDngGD9cKOcJtRtMwmB/kgl40pxSjJvupCY01sP1S
g9Qxj+XRO3iqfOjqYSMUHuuGvCbRlZqsinr4zOU5lE9DKvGIs+82+94II8KCmvE2
+uLS+ArmVEoem53ZeneWz/h0JNGOyTNFBFOUVXFWgd4aiEq3y4AVUT9bPhyY3uV/
XzQJdAQu/ie7+so76F60dX00+QRr5xWFMjs3A9UPVQh/ekPnUKbHSvDzczze8YcC
6F0DcIAHXKYcBqJMwu0ftRWUG+iYv0BsA8M0WdakDwo2OaGGwYcfb50Wgq/fEgVu
XglcFEnL0BLyEL9qr7gsfmY7ZVTC5arEjNLhNCqQDVD3GUaMmptTbxRpTlgutfVv
MIjJC2Agh6evtee1zigNrqY5WjvmRmZLPhrcrieWxF5EQpeZDzh3uDm9c+JqqLCb
HD70Rx01Bnaw+kDKWuKk8KAr8Xtwzp4ZsAxxeg0oD27ej4iiqjfRd1m9L5+75SaA
6i8tA/LNKiRtW2pSRndlz4h+eOlxBOLAJh51VxVLnnAo/aG4uaPWVvQRh4gkmmr6
O97SwnICkf5o+eIRG6FELWdcfjAqwcPh5otLj3luFwLewTQOn4DATN5Ob/GHfRjX
7hWjX3gKXw/H6mt59iMf+Lq3vLzX+cCM0Ol7IP1Ga+otEWqX87PBGiL59lIf2+9u
LEmkc9fFkoyz3RimYmLJ3O3D1jiElrQ9ZKfTnkPl272u31XgYeYdXS2fd3gXJORB
iMuS11uphJF4FYXMk68/TE5DJ3bnastyrh8xZBIhCX1K61Z9vgc1Lb9DKm0s2Ah9
ofibe5tIINew2ba9AmAD64ilkQA4AwZI7ZPfzPzhrkgiXhFFDqajGmwtpseuhuCc
NIkZ9HnjgKEN08YT2arBfcKNgYzK+aAIhDPYxQBg06xwQpnVec8n7l0EyUe3ykM6
yj5M9rNqkcxGcxDvMpti/uor7NKtExZeER+ih4DuPxmSap9Ax8wjGAHUVQdGh50m
2mRb/dAHgzLUn06qwkIrkhu/jQmxPBXytGzT3YHDc4Z9HT3e8X0v27JYHX51PMJE
sbaaaAVhcRTsAkjTdzMIQNr3WFQxrWkv034S9BOOywOjZuBBdWEfm67mFKvQSTu0
E1QzZw15q9KRgH/sK4m2PfatVH0sZBPsogjeLvLRJeIx/GSffmlrB7VYMn3BVimR
FURGfpK44LgQfLk16NA+nwQkZ1kcOvALvPMqzgg6Sl2Ic5iE//g5QO74cCdN1FZo
B1SVri9R62pkc5Mdc650xXYHFFzYH8abZRsFgcFUyaN1NLekgVSkM4RSP2HONQr0
R82QEJnC359NzjpHKp4SXDMzfcitUn/Blvl8me8/h7EplHGCmaYJFuW1ZVybaUDl
zULUpJvUnLvy/ZvFUSJAyFqI8YOLd/ZP4P3NYeiahNB6jpYk4p+JZ0im9tSeaysj
MVC1UckjWOKEkrGhCMhhXEPhcooifKHsoKWedIx2APHPYeFdVVdvEvN310FG4fTD
thiA/dcXLMRYxFZIwbN5J+K7lGSJQ1uu1NvtXoozGyuzVzVWP0LmZHFT5sp/llsJ
QUiONU/40+7bQchcNjErJITlBwIyJhXYee9zrkWErig3FuSUy8IH3UsvIJgsrWQh
nBWY3XgsH+lhH4xrqHrzMP9ht6O1nXFD85h+5wsPRgJB/zearWfUgzvevoDo9m75
CtFHw+wSXUkMYSPBJ2pH0nwU0wOpmK+y77hia+q3rTG3ectv9jmvQE02ssjiPF/b
oA3UN/fzuyka5Ymh/KAdlvgMQwwQoOvswcv1JiYILVbxtvF/WTjy/ZBHRhrcZvgU
2FmMY1UbDw6tCYJgkAqXjJBOQL917MkqgTYPLhEVc7kaNHNq3JKLn4m+MOziqlpk
dQy+PyWzq5zvUfatgcX9sRHlSCSFbYg7lwOtQnZJGZFtUUKpc58wJ/k2r14NkBtr
4uYYXvfAlBDGk3DhEg92oKKj39Tk6WlkacfQKNg2HFQAnug9O3WvC4QA04ppC6KE
3uh0jlHKZbSE5f/oLYkXCT4/zInaaoALQr7IhP5Al0nrwpUPiiLOISxw+HNL9h7a
TSE8sZDgHiLplV1DZ+onYd5ZNJRz0UUQE2icRMcjYqZzBEnhsgYp6EDQKYp60Rbb
qGXv8lzOxsXSOLRZLFt0W9Vq03Ojuxa9jLrhfWNYftJO6drm9wK/DMjlW8WkHuAN
B1T7fIPgs+gVXV/diQRH3bvkljVryenLGTyMZ8F2nikrnoT1lsvdrY2wNXRDqfY9
NsQR06e3Jr9HbAFgEdh8DKEcN14ivIIgf7sWN2Vnmm8W2Z+Q+1l/k1HV8W7nlG/X
vzKxxVrNiR3HuJHsPkO5t0amNmbwDn8RJraZpJEN6B7ENnAovqqZElTwL/9LDuVW
fCvv4WMKRmiGSTbkr35anIF2FWr9gsRDGaK4WY/GglvF5V1VkbAYlNnZxpMSmVP8
G1ZTQwEIVuvJ6dnEvGZTVCJsoLeN1f8gt8bXH0IY70QwgYc62xre5VG3gkyy/CGc
XYUC5ylYDGo1pAPlnJV1UBZzRP6GUagRCf0CZsjm9JPUIJSa+f5SgG6TrvAHvqj1
L6K9EP283dYC3IGZ6zt0tjCbZ4KjYc+Vqrs0EiMgqEZsEXn41wCM9+cLbjBuoRhN
2H3a+9TX61NkD+jimqvib9/o6wqBcPdQT1yIarLUlMki7ieRKzrlARA1D4StXuWn
EiHjT091Zd6n2CAmREXRdK3CRm7avwY4hDdY/tBcJgK3ed0YgHvPAHLIDXBsv/RC
A3vBSmY7csWq0mk3YY6Qo20fm2DTRba/IxiiG3vIER8nx23s7fb+P50edftWzmFT
hBfqyMV7yn2wD2q05Mixd4j+8o5hzp5S29Z5a1NRnzsfJjGWUUee5ZVcVpO9u0C+
Bxr6totHyBxjjtyfRK4cIoRwUbb68Ap3lnqpqVHtpDEeKSbqMOqKenHlSrYJM7VU
ghy4Mr2F3oK4R7eGot+P+qw2dX89D6D+7/tgcBkJIDvh3GLGyyZH4VigZ6PxwkT6
tzDiBGBogN09Z94GIbbIL6B09La4uCyTOUaxiJZC+Zc1GKhQ2GInWx5F+rJlwnWg
Z73u6mJCcioZlzGxO493QKHbs+JQ/ckXKr7Z3JQlLpn1px89rQ8iwbBz6/DCgsN/
t9gwhJncWoxjTt0scR18dlvTdAoejoy0GYS9dIlYn5vOpqLU1sGca+AIKnd9y2Ql
egR8Feuud0bQHtKkYfpZKoAJTBDRvXtyXx/LJHc1Xk0FNe8RqzWcnsgyLQl1SepG
KyKVCoUvYGP3x2UOPbwvpz4RngIcBsEigR6v3IKSGvvruUXyYdgyQc+vnfVpUykw
dte3+3ijH7CLiYCdptywf8fskcJmQp7s6hXbpRmDK4DZfvjEAe/OmvqpV7G+hFzH
7zTEnCUtp3B3tzrE/E32jgv4E/YM/yy4pwYtM4kD6XNpcK3mF/tCdVtwhqLO+B9I
pHBdlciZUPFZx+B3k0TtCbWVa5tU24vGExUxhxzkLiuQLEhF9v0Jme2wBujJ/u+S
GfnvHhuN+Yykpvft2c9TQ/xl6Q0KqEo4CM/wjwBEjXWEtyUJxFNy1LPq4Cdc8eVZ
n3crWu7cJyeSFzj5VyfowvOCCfdjLJsKul0FB9HKBOVUpv6H+H3mOk49LCt3drMv
tjXnSp2KLHJN5Fqb8sUPqeAQDJh5ha89AzqdTtlxsiqixsRSetYKg8nG8P7hk6IY
UtYEi/HAR2LQDOotwCUStlDxvdgraKwfgCe0gJXl/y+qlego82JkOM9PbFIJDj9p
WzlL1wcNsE1AucA4Zv4bdeHT5SWsaw3S+NpYdrRpgK2m0w++tKXkLphsVhv2o1Xa
czF+ZHB1/WgwCzMpBfo7gGVc8tNUfWaOYOLo5mFb+Twyrsa42GPlf9wc1MW0FhHu
6ULR88RRXwLUZYXgoMB224GplOxf/5+boAv6yg8NO1xTD4HqBHl6exkrDkNALMgm
s+e4+WIsl/eoVKIS2YhzEFZBGM3WH1wp0wAb0xjaYDHeHCbJAKgSGOpWaw/ItO4O
v5scID3w9KcdjH/UBuJYjsBtjC+uIxQIK8VYtDMBGrSURCQTCEPuO79egVVbFxFu
xzy4RXrHDGwvQ2VplYTmYCslj7Mvyz3Eu4qkZ9vEU9g20qo4PRKOqXL9qICR5JVo
NPRECQGDNj5r0j11W35pseKdMv2xCxrQqMJEqK6TYKWSLF4t3QeyyJI0jSRMUHnH
aC+Y66SqrRxus3+2TUOmXe7Xy09GUCWKMW8qekdxcrW3wYIB5JHhCvgaKMwxqVyz
X0K7m+gQGNAZibqheuJC4yTtqtCCzYu8yRMTMSaPTqgoOEyP/0XtOtW4bpZu+4mv
43w4vsNa2IF7MCU/S4x+Gy30XvJBUDj5b/OQ6r6SHzVRxSYPRDhZUQWkKtFyO+UD
zY5YV+VcTeA1NeK65WXisGNGb6swypSx74EiiE1n5zFcuIcRqiZ3h622EzrmHNwM
w6iIFbL3wERQIQQeL8EULySpJU216/93GnUrDhhxwXvKLVciSoSzQYPU33CyU8y3
dy/pEHNEPVbhmgNp3UV1+EEzONN5oH2yQkjjFkNC3lX7gCjuVd4BAHeTxt5dPu9c
1aF8GtE99ihD6Qfo4mukyU8neEhIscLfTnUhI4CmPlpc5OwbUsQycNDxOUrcnF6D
kZPW+EcLhO7K3z6Z+ch76rPdaHaau8raqwgLqwzktn7ESjycmRoUt2DdhNnU70CV
Tg26JCOgCf2muNUsj08bIZDqShUTFuGUE3iKKJ2Ki3H+K+yfUaeVB6ZWQhADOXtT
6LlaC451VrRu76ZPjoov84Ly8Y291EvVn0BLyl9GkWNzaO/Jp7sngiBxq3zJe/7A
aOMUpVne7+9Yzm3xHUgRrP7yWK+Q3rxgYg2Va2GkKiAAON2Zj4uHnFc3NiVy21OT
pF4G0hH3N2JqGozIXqa7qX7gFsJm2nyrkTZbQ+mBnRBVOnk+lOfkRHT3pMW4CwD7
yQwydAVyW+FshKu860w/R1KkvptGBPPVb5fIOnS/oFLdsZg0nBybcDopQOOJZFvS
kLVPN/T2HT5WPBTmq67pgueZOzZn9NXXaGMyrAATxr6SnxdUhfuNwivOYu3TTQBj
3q0VHVlzkpyx307twSgvsZtFQJCOWII6IibdjXuIqez/P7E/CprLQSDQiuf7vdK3
OuHFUF+F0URnpZhHOHCWmQHwMf7zlIauydZFthd+rb2hn/MgrqlwSMisAYYkaKLJ
yGSij1CcU+n9Kji8HRwL1GkDiIi7I22f9xhods90zUwkm8P9EVCl8bFLMWpXsH2B
GINmdCiKFJv7AJ1TwMuMRZBrxr7S+EHeWiTCKAy7yc85Y+96FxlU8ukszoMOZ2lH
jHat62Gms1x2LlqaPUpXi+kTxrV/r/Nukw4vhUNR9SYM5i6+o/b2irVB5fNQVZji
kLR5Np8r03OedlOxq2RvsEz2kr4gKog1Ew6bYDd6eZD+LaZWAkZXI3UKwrhpJzLM
DCJUNu1KcdyDIHgL+xhbVm5/aqphWP8vqJ0N6xbnRo5SD0oFYcB+1TjN76a3tnxB
uZDgPY24W1WYZpB8tsIwkvqgmhXvHB3sCApzauk+6ppd3Ka4gc6BSarVviuA3AxL
ofUrdMJeif6MKkyeEtXwGYI7f8obAwjV6v1C5+BkhzMVlEiP/PLQ2Ao5/RTuaeWH
Qgr3q8e7nLVF7TGQoZiRc2vzsrrpqelMR9TgqXdQJe8GmpRs+3xMuaOWZYWdfBxm
jlVn47IhTA4pufWoZsm6REFXfz3xWxC1tVC1g2PZ6+uZBbcZa/DE+XayQ95yqbYy
GJ0Q2yelaiUtosY+m6TnDhJb5Wn/iSBiD1kbCukPY3VwJCeQcgTaGoR8HXUGjAbC
ZlvmvpA54pozkFZteLFAFaSyRcgrJRwVbtj4XqUvqL05EbEZGfbFNr2oebbaZYMl
zw4eU1QspjQUgMaUVz0AgZZ7c9Rzw9HhaCs0xvfh5VRFwWXTQzRYjmMLOy+eq6Ug
FLTK+mITeBVRvZOye5XxknOOHOtC7RMogvqHG+vgzhUmnemsLo95i74CDLLtLvkW
uJxKOQlKnXb5guF7Ollsjx4/v8CzbwiKZ0/04h7PAaUUcPqmXoZgi0g2fmhv0PAo
XOxbTk775d0X8qP/HqpJMn6qHldm09HdHBOdinvc/ITfVbqOqJGVk7exFczXbK5G
OYKKf53yMTleG+M0cUXVTw1qck+J0CVFd9Q09WAOXcXEWRQleMDmZrvJx6cAIIW7
JCm3Xu7yh2Nfqp/7Nbm+Pixc63ElZZGnUwNMH5oSACE93L+1dkpNqrWl/evqBN0o
x7jZU084V1mBpnGuXhwNgIt41IhdKbkT3WhRje659ZOTwzAsBv9y9pMVsVny+4nQ
0lLBhccEOIQ2c0rcreCYeirp1pDAmth4v86Ej0uSWBZsPDVs0WbTvPOAV3yBC2U2
aZpUOri7cZ0KvMpo/W3ki31n7zNt1pT9c5dP88TpvhfO+0TaLO3yQPsyfYKoOEtC
RwGhP1f1zdMzVNTjhl8E4VOInOEuT47NYFi9MASNc1CIMmPlkux+2uWv0E2g7Ois
e29vxuYWWmP+6EAeDan+N0SNuPzfmBHsBXALzsnMTYvG9zmVi7bGiMUUM247Y6TG
wv7O15BciKKCnmfP9Eob/ZKpmT3fCYsDngzgPxTPyWY1tf0xzO5+vwQIsn8T794L
d9O/wr4ZGdhl8K6tAx6DDIhLeDSy1e9m1BZBHqyN/S9rBIBdL8LdGJ1OgJg86jVA
NekoZq99ssSCTIDRtGJGhgwBYzHkvN5jJVf4X7lhu4GaPC8QZUpRVbeLopp5lRB6
8OVCOI63QJE5Rbtibjfs+YBvyFTXBtWT54z6BbHMIJgN2yHhCHqj6h93Lp+ax2qz
Ku0+YRnYstkuqllPSZBy6W5caAdvcRq6GX/spTJ6PETP4NQb0OQRIIfUwDc9yQsx
e6VON6On42wZr8/rxF4+GY1EXcYSbDLzKxp/fC5f8jzXNR+BWNlWBijCyFlkyH0+
K/NW0mZTD7AYm+A1MFxU5KTRprUQXcojXSMmhzdXNxamFHtWjV3bTr8ssDrCVY/S
iyXg4lWVgW/iTLikrphTTNtBLb1X+stYJPggu4mMXsOE1Er/O8YWeNTYhUyQZS2s
ldGqvhOFHHneV0c1jlp/qQT93HJXUrBBC92irIwPjHNxE9SzzuiUKLAAuT7pW81V
2GlNSIt2PvCIGGne7mfFO/XKPuGnxIM6bC889tQ3s9V4gUStiN0UV5LZtNNMBc35
D+OPhCYvIz3m6mpGeatPf9TVOP7HPcH01MVPp7DegkK9ff8BuwshCM2AoE9MAglm
orYGGk6fG7bAM8aJWOBe2JUzVlz041gOehonksn7AKJAFGB3qKXzucYY9juonp2q
9105pDEM3kBe7Jm2wZZcJa4oJoJIvQ+xN4Ep7Y/y/8949PW3RNJZ939BZKcaSmdx
CEjWiyFcOcaLms7qJ7F0u3QblG3K31AVLztUQy3fS48ieZ3TbQssAPefA3nP5j8T
KxOZYIMiVjAtXoo+tL/VqfLgDRtTPbvCtK5cGCWvjnIjG1ZXJnQbuTzceAfMjVND
Qw7trHxqzlJ3myTPuZ40DfuUWRxnChuZCVYSFJOpjnfCSXJNYvO0T8j9VCTWwXjc
RwQ67KErfg//UOhzlxC5ndhxdgzMr1+VVsEhlUbTYpOTX5VmWdNp0nD21b4EyGBC
WZs4+r1ON9lfFwMcqRMpwREctP3kan+5nCL28KAex4IkC4xcsvazDDZw2EeZAEvA
AnF8lv16xgejK4hpNZx8HATurR12If7OCOZyLIGcSBXvVSHAnhUQ4LGzmdSdNfTh
pgsGl3W4hg3NhGwSOMi6MjBaP24oZaP6j7m8KhBlj3Zf9vh0JN6ISK9Zt442AmGD
jrcKLDXtam6bqaqXavlS3B939xTGK0Z4QHBcMb/8ACHztCqPhBb8BGNsE2NRNak3
aFRZ1LDQboI6VtPkfaIN2fIDdaFeQS587d+W922Mdxi2JLde+LwiDZ4fi3/T5RX2
sJNWEp7FsFctjraMKLa9ig7LoT9+goOgMIzBDrw372L391qbsgSWeS9danK3uS55
mSJWn4Afd0H8YGIXuI7fWFSc+L8lVwvnQmA5zh/9fFVy0DIBbNKsacda6TMDQuGQ
xVlpHqkKM6SEB8jh3cIx6HuhueAeukogVa10hhdXLobxMasAuogcf/Z2bElHLggD
1/4oi2CTIv3SSBDeO1XDI5A+Gx2tivkA8BeJ6JIIvEVeyASZL7FePiMt574iQJd3
639jdeChRfO5KVCMke1XQlpKiJfng/KPOkhqd2bO8BMPDMXU2Tf7Rdk+ryZSS8YA
Ritma7WmWJBSqyAof4GCV++C73ELtabMmAPouyoUlxvEfymMFXAmM7IcCF5IUhDV
d4IVPp5lhfPB0AY+lTuAS35Dtq4kqLjd9sOOG8F1QsQV2DgVgsLye5wmUJdIvin8
iDuFRwtuN7RSUB76MAeMWP7DAqv4RUX0lobQNxCa70kUUrpcK6Z6y43HuK2VGWIO
R0KHjhmiTd+S7D4fbxjXcm6/bb9Un8QQUt3JizzhOSAYv1+JmGm/7sjjPHMVpSF/
H6qOoRyJWy5i2nE/tDGUMjxSSJtBqFFPpDjAE78kH66G9VawwShIQOR1SgkC7+Y3
W4Dv6MBHloKSI8JkI56a/VjTFUIO/bRmf4Wmov6o2LJgusLDGjy2gwH3R2fYCZ2z
M8eboSHT3ssAncWT+Vhiq+vMxeNaOV9+Xr7L5eMDWFy/rblkaNwv9hqtACbLrrb+
H4+f8P8Eg4H9fUL8GjXY8/c2+HgDcbdfp1IMELzpgCMi1xRhK6EJIsDFpNNViqUp
7xMhQx0EiV8jbfFTvpaS45id0aIiT0N0capnybeoBnbNPkdrw7dWtk83KGK1E80m
V2Yfluv+rMK84GYykgDTQGSrUPm/s0aDgsILu64+RTL/EJk1krFCFV+dRxFdqjoo
5naClABuGS7AUfLxcimn4IoL+IzJLLFlYHgC2mJHJimea1ndWyFydUoAQ7OE8T0h
mT92KMZJdg6TphAnXF/vjGxUUB7i10bEDdZw6Cx7G5+QdclZK3sVXcoSs9ru1/QC
Xx9Tb8kiEbSxSYctmv6mnzEP9qGK8HubD7mCVdHu/zzoLs87np/1Gp2yMAJB9uph
bYWaLyonGCCuM8DabKmi1zZkXTWCbX/8LNCeUwex047JEsC/G/mnqRrPDix/cM1E
DxPoYxiSSRZmuKZSaKsvbPSeot12kS9hGT+mSQBENhlMMXUzv98a7PFrX+7ynjQl
QtbaJXLw8uQersA4UQRV/P5gHmiO63N+zPPsfH2Sysf//TtBnaV49MZqeM2euWYd
unPx9HdhQM+uLfG6M6/JYF2WPfP2wdJHCQDtqE1c+uL39W4FNzL42u7D3fNFtPui
Kra0e1CX5BDVGVxb587PZEgCdn7r91dBvpCOY9zGENcYzldbdIssCUUiAsU67vag
enGHR/M7pVVtNAMfN/Z2TD6KldzIKyDYREl8Kx8QFxsh7ejSN7GmpUMC4Z+zoCkl
WoUZRElaGr9P7gV/n3FxZ52g+S/y2ETaml3+11xFciq92tXaE/kNlrIKBYmQl7m2
8oUAIfnXBoJi86EB2sdXT5LHDTjY/y68KqicWsb3cJ/BcmYkh9Ar6TO23nkvhu7x
YnBs3zbfPKDdhd/+pr/7Dl3UL+IETp8TV6jsn+Ngh+3cTG9Zyb7nEI2zg6km7Xq6
DMMbGu8WNV8sx+OrV/C6lCK+NaFd5oZ54xeqbJ6SHnzbVDGZ6W4VcVEcNhZ3MJ0I
kRX7vLjrV0m0aWbXuTjeSA+TZFxGL6z1UieaHin5qUjnBBPp7LlpAeZeIw9whXJo
xya/UsHn/u/b9a9/8Ks9a0RBak60vbjcuCJ8xX1Qv/bBsiSDql9u/tVnN14uElEH
cug5zU43t/CSdH1qHpBctopKwD20tuIFD8h3vPGOaC4VC4XlbQWc8rlpxV2HhrE3
frP4FQeFtUIC/Llnn3hKhtfduAQO9dK2LA6odwWlX5+RysGzXY9/V2VRTNpCdVEN
wnka7ZTyUESy1ozcThFr9s8Hnu3vgMtOXLFwEuTTM++NPzLGiANZKjkiHv1jt/zz
5MLaelDzvLEmW1RU83Uj7Om2C6fmzaW1XApFaE9q2hNtenquNCJfZL2XkSkPe5uz
i4//QtgXVNoPUCWDSi7TS7I49O3zWf8WoMV5rtLfyzgMemk3cIWs0qNSpn6qbHiO
TjHFXcNAWSpBDLQ+FQs+anD9ZsbG71eVowuj7UvqjYb+ZQCjeepK1JdUTBHqhlJF
j2JN7D6JEjITohRk9p8x5Ha+8tADbApK0UmhsLR7QAuuz/nnWzAsLbkI5mvDAG5A
hFg03TsBDvWSQD9w9sI2XK2YfZUPXyFRSAVEBUcDo5KNBIXWFsnRiJ9Ir+jpize/
yU9ZEHDjKQ5Ln2EIicTzSCBTH7uCwzaYFobUmu0IRY8smt2Z9AR9Z/ns5TmpEa7L
PX4qwh96NB9oDwjE4eqBNYDq58kDjItIBbhMiFWkdooxlCZW1Nc0ZD6mBLL17pFV
q3RigWeoBCm5gEHYfqOTGzzAuLb8t7RkKzP/BVNt5Lghgqb1aSjWCmLQst/jLOCO
JQTeXy1zdswh4uyHVBv2K5SHlhTN2cbbsjb+RwjYzmEGYlHxMkyOSOgje6P6jvT0
YTXGBS0vtt+ar7FyAeVDRhtEthw1DKZls4GtLRFgt8FfMf3dufzm+KOBEI/uSJ9O
Gju/HLpvpd4CVX17XCRo0EwWVWpgyQ/131PDWu4stdtlaj+gZiwrvrwkqA0byCbN
RAiWTgqy01ztWIMowIFBvVp04LI96FjH9xyTIYYowMprwtx3NNx/nzjXvUBWv8C+
7M5jh44Q/iEEnUlPxOvyKoGISfUGZdcbjav/4rKO2RTpv8Q1B9tAyurce1FVXNVJ
VkWf1xICa6XYA8QZnTP/lsdgjYNWfozE6Z0mGibxe5GiiUx1WdVfE3ExgqLdlFk+
BZqZ0PdsqFFbKk1sJmXTsE6nP4NKEERt/g+nhhkf5cGmfgCYB5ttcYWb5+IkAO3O
MU9d9+RxIwL1lSjmTWNBiNuUx5L56FOWIthhORYVSZYrguIrzmu1JhgJEeHRabf/
KY7fgMdTdbUfvDO7z38HWkm8VQid62Je2AkvV6xRes96HIPtLFRiU5CogxG0iyuj
pSjplL2/LRHUdiZfMI53l4ij38fw60vnmqnmaxDsrBsmETsi9oWyAe1DKD+2GF1R
CooftJMUyICRLaoIFwOzYygznzp211wMYtSwzIVf499JQgpm1IfPCrqJTKIVAhVE
6PCENAAosfBc7izFC6hKi4ljZzv1CUtJ+61U0WxVeAtLBe/vsiAb/2bVUtiQmYXO
fjiP9PlCzSDZa0XhJrdhOvbS8NBDjTQWA9iBW0ee7QOHPyhwYKF22LBZouzaxkzV
puZAUuYbWnYFjsrQ4JsEVwi6c0wHwL3iHGRt3VSSU2Xc2zQEQrx7m16JbS6oFGAY
CW/51S0Yijw34G4v4kQ9tu8VVSP0PXAH9U4uWbil/JWOtTgR4b69PS1KLwYkRaI5
nx8pxngOktqAmeooRq76EIHnYw1xlxR0576aeA2sGF0xivUDg1CT24M6fRz35fW0
v7lB0anKgvHSx/caVM4B7FsQBpKOy3mL1a0guzt2siQZ/bGL+oP/KBbtClT6AadY
YwUsODUv6Q9wxHgsC6EjeHlwVNkC20kzYQhlssmBekEhn/1xAB6IpFlkZD3Gpy4i
XkiqQM/lW9dVNfEEXglV/Tn3eSn6FH5hsX9NiOKw3kOWH012PLYNzCMGz/kPowMg
2/aoeGyWq4Qe27ZEMiORUHQsAHVL0wVHtcJZEheOu15ZKrVV6TxlgTu2r2ZCGXPb
Mq25/rOvvndFwwTe2CETnenv09SOek1FDL6cyoD3WePVF3K8NeggrmOokl3e8VF8
KSontAplNW5mfuSMXpXtvZqvwenRgnANVqXbGrBN3Biz/QsT9hDwjVhJb6364Huz
rDocwGbcFLqvux1hlAxZfDTO2x9BFoTfQscfGIGp+kNKfsCpM3InsmthgrTbX/JW
iyWtyP3FNTOedL+pO3+eCPCD+JvKyRGzDSRFiZk+wvBQCVo4KfWekwrWXp/K50CX
o/1mZfWHxTG+Z7VXE8sdx89Bxq5qWm+HsWpzQzEkzdh8DjK0B0CFnz6xTeINt5/5
u7BLJBlgZIda8QnGY1wD3qsrYj7lCKX6pvecbYk85J5KdxNdfVDgk66/o7Qddp84
fQl6/+ak1pA5IBMPuPyWfzbSgPOPI6IZvvmt8k76jke+RezRwZb0F2ZxitwFbjpO
aVfKmuPxghpxf9zXa7YUZRc4tfqvsE+Pix9huAm5A66i8Hdb+4O6eSmSOAk29RrP
JBpxCQ6Vc8BWlwHcn5nEXwgIPaTxR0r6U/oRlTFC2Olkxqu2tx9Mc7yFVLLIzFK4
t964fH2ZV4GDcMov9GS4L0avcCsamUrEuJUSkxCNkHr1Yt2Yf52nz5aQr1pbidcW
GooFPy6pxQkkEFTshI06BtUA/mEwH6ayHzvNr1LMuDYPmOHC3nVKPBGfjpQgZi1k
zf188B5kyo/PcPFQvL6DtEifsY+ey/v27JSEQndTlCAzdauEcc8Dh/ropdmt9Tp5
alY8pvpK3hx/HtQu+Yh5ghy8lwrRtgPTxmZiiULdHer/aQTC3zyr0hwBTRXyr7+X
O+he3a3R6meRA2OBYc6L3u1msUph8wEq6Asy6dq003Ql6bxsve3JhQzXT5n2D8uZ
U0FO0DjUlt8pRZ9bDXZcIKtkhylgxd7+ICwnwkB5G0BESiYz9lWuea9JbJa6Ckvg
G+rOposNWuAerZu+Eau4Q+NFqQTSXAHl6Rgjbv737W1rK+U9KYKCA7G2mYkqYim8
LP2z1XawLAx1Qv48qJuBqEZziT4UsIotFrgxG+Ckh91I17SKHFsXgGVytGWY9nwA
TGWtYEcGN8zeA5XJZSnNXGGVrOYktICPtRHnAw0TZ++XpplA/RGo3eFeFYvPuIsD
0k4Vtkql6pzJCz5vkGepcQSXEQnD7nLmcedREIkXqAjYEwqEr0SVsmeY+hgshfUU
cZduspWH1LXnJHlwkl8PHErT2j2+7UH/3UmLjgqkIXZz2UOB14PKlTPftj2B/HDD
Z4IOSHwfXKLu117fXskfq2N0h0+wb8ykP6rMOH8Qk6YGmttb/8tLpAT7lI/yFFSa
fJJ36pBz1R+K9bYW27Dps7eUIDV5jCPBnwFWMsdYY4JxDYZuDlr9PTpCzR55AaAk
7xR0fCPxIpPglLd3fCWsV4DGAnvLxAhcJZWOCL8Sg5a3xLpywo61ZD1i5HjjgfkB
uCkBorTOoMYB8h2zsCj5ki86BzZkjUEg1CfbxYOIIk5g5eqd7wdkv2D/OkOEtQMh
1B2sbNKg0olpplwXg0o6ZLEzwUSmfAl9m9H76AXSb+mDqg/tObA3LxVD4K7c4KGn
MVB/RsF5Efq8ZsKFsnVYAVaFAUnJxQLiQrzAdoJWQ+QihKcN9RRLxD54biii3m+0
Q0Ig5rhFBvFTRxivjP1dQCRZ75nh0nBLWn8nv3kXwLPmtftvXhivQU8Tk5PVii/b
PzKwQhQcepcqzw92rGs5bcwoDlofHUsqpcjeZVvdL4Q1inLeWPgi8EDu/mm+N5uY
C4iqNzJCZa2HifZbdZAEjTTW271ZDh/uUayN0Wtmf3fcelWpn+A75aly4U5zH834
GnTq/TrpvlT/+ijYBuz3nUrBqDvo7fyWl1dcIcBifBn6XlabLpHkV6WmsoavCvo6
2jI9576TP6y0NRpePxHg/RBrgsOarQyhlQSHWHx6f87seXFLJl3ZfWvK396O/yLG
O392yyorv+9HXYgbOjUa62oa4TKtQQt1mseeYFzlBZUkmRqzeTtKF4r9HF4tJEfr
IwEOqki/Hgv5Z2dSxqZCY5fg1HFmYK1g1r0gcpYyayovLaU/5jpYeFw/y45S8svo
f6PBqDuHRJ1XWbHQL/+5lL58mloljtfdnquSEfQSKhfyLzFqxMN83A0W6rqfdTXL
Pm7zOmSW07S2qdCtZBEQKWzv/qWd5VJ7YUUFeZIYywpHe6BilrSJ+V6DG75KTFMF
FNaG/0K1pAedEwDxA3l7MLLqZO2PGommsPk/FeT0Sk0S92xVodZ4DpeZMTesuKAZ
A3eGoiqdIg7v5o4fIJzGYjRMnVnCsitQWW2QIHsPNljrsWVD20mEY3hKi1l1q0Wm
Jl4rYbprwUdsEDQls9Pf6Dr/+YYBfaZa9tia9Y8bAzJV/Q4GxqQg/f0Y5Lnc7g+V
3msMYrWGPVnZB3sqjc/8lQd8AWetbcBoIdDfyY5YK8MXz+67uZv3gelxRl1ko0Ot
4xjMdueBsoGzyja2IBRn19u1MfeI4s28S0jKWsZTRqG150n/xrcbOx1SYhMwiBsY
M41/ZjyyScIHDo7Tfjz8GzHTXFgxyPPed0wK2k1FjC2IpsgwLEY8+T/6rEDtw7vS
X3Tsz1jJaC71iC616/3E7H88Egkno3i2RRXUQCZa03S2+o7ce7blEG2XPulPhT3U
hgbizcULjrK5DHAFLx3DvXes4RJ3XX+ifXJkA+jqcLEZE1JEqMdi4OTeflPkvv7R
1kVbmp019aqWBORn1QsHvOfLA0UwdpV15RGASp8u8Si1KFh9cs/L3TeKErqVE1EA
VRA1TkoO9F3upq5b3od6XgIkGY8rzoMF8FdxF9uZpLunAE4808oA9icdL5agNnWI
ZiTc3/RPyYp/3Tom3FNSvNf0qsbmhiU0ytE3JNFm2NKYzNMrBiHL4l940ixEgXTy
3UQPHVOutSsWkAzbZ6lJd4tYqyjKOIQhM3GHaEfONjCouKG0A0ay4qhgbk044CwN
L9+BU0P/MeVtCVWYZ83np2lsSrd8i1LcOQlxmFxxFt8ui3P/L7l77ACb95FhrIEb
J6uNphA2fGU0TdRvMmBl3Chw3mygoGlDITzMgmY/gOK0k1+KOFK/BWICIPM/wrKZ
QVVDHqT+E+IPiqN6cFEVZOuVDIzX+MJs5FGpcKLuriNL1fvNct8baAEJCOBW7MTf
EQqUKTm/9ABFREYyZp01kw0Rv9R+pDb8OazKPJt8I3WJfUOb1JEX5ILDDU9uapde
Yr8ke4PFjhAKEJS7KYyd0GgOhqqQI2EES7TRb71LIF0X2zcnY7Xry/8VFgiFgU7G
cZNpO/YuhYxdhy/BQxQzAzJs49Nbezvl4JFGsZ3cqZv64xaIkQzT87fguMe3hdkB
xHeu9WHlphFpZbOZpHFE1AcvX8Gejh9E8wg5m/15fqc4qXfc0c1EUpuQf6IdDEQH
qCR4cWxNAJ67e4q5w59kMZQpxpdOgUp0ydOXZOCZSYN2Xh9UtuUr9hZB/mY5ACYj
P2zwx0SqlUMPXa1Ry5bLbFdWCKKyrVuDNOf4IN//WRi5+r6jLUjylxYrmQ+m/vhZ
hH7KyOhh3k22bq55ycZqtluPYi+e6xBhFnLJhnjGDIqOyQMw1WkzkNHYaToOEqB/
X4SBlDis1XdXJAaIGaCDkHhNVry5BIYU/zJcZcFYf7hpEayFCBfF0/pxFpi3hicJ
jxUyrHFNGo7HJfp/cT7Q1rzKJqf6uZwmgz6FImg9kjzwIOabeqPZV4ql7qLZdKq7
RY7NkPkuUtunyQOf7bHUGKYtVbGiuIfEENCkjGgZwXgDR4IU5xUxt6z+LCB7B1ab
2Hj+ksrdpKAg4OWsYlHFXYBsERd3f9HjnvASo6VUbhQHoroNDNkcEjpRRyXd1kU7
oiWVjj9QbV5qyQ+iR/CnL3AZKJa8b1H18Wy2NnUYfhEUaO/EXj3VLgKStWnZBu37
1RCn2el7x8ETfozFJwkfCOa5hyk0dizFVYtQ9pW7a8rC/bN240pPAXZ2kRIn2CC4
BOY1iQkmCy32qBL2mbZ+C8p0gP0hsCHVH1tImm7RLWPlICom5Wl7haFCvHVAMWFf
FY5kMlqmYVZTTjEiQN7+exPMteim15LpuFveScGm59p4ocNC8vwTIqo8tkDngvN2
500jGvtVQ8oVV0oQGFhx0eQ/REjbncHXfMqVrx7i/6vCFJrHOTgNHZWx/f+e+m91
N9OUJ5s5/rfVBylXcmh8YzWS8kllEyhX3WbIF7GbAatWre0GC/Wjreghj7L8lbNd
SlX1XKjagy5+YKybnXWxGfmKwsLM0AM5bDpu/6ty8v+ayQ7dKWwcaQCCzTwFQvhF
h3zCkiLd8CqfFutRiYdE5IPRPOeBvb2DvlZX7Ot/MYyhR35FcrJ9N09rLokaeD7M
A1gcc2n5s0Jvyw6aquJr1HlVCpGL2pOmPYOiCz/cDoPWBqv+aXWMf2Si0i2wTl3B
bJNszH4Y1S2384/kDnh9ukm42uddLVHjAvlMXYtiAPfYkRqjWidwOY7441W8/su/
5UyLy5XBZ3wH1S4vraPfj37vAJ0ZnbNQikvhdnQYQc/8B6wK/9Mdl9IeCVUi0OHZ
isGtUxAuAm7hRKyTV5/6pQgp97Z4Oqg50A0+FXxGg5rfkrfjwPKK/7Mnw3I/jXAT
i13Js6TFDvAVFYdq4t5e3vrpZtvIMWB5Ju0NTVaKPOHy5cq3J/9PyELYLebauULz
NmeJec+/dwIvurjxri3iFw/nINLIagqX5snaRVkVkYSjD4YgGbItWZlOeD/qWz9R
GN7eZyBcnpIBV2seNX1i0nuURN6htFQZn+QDKgDzVh7CnfOLB/XbPdlApMyKPe30
e3i8FWZMIXYeJLQlT3Q/mINlbGEQI7o/+cEAd2Ni0aUsIWEGp3Z7K7FbEK9eS0f5
qB4aKEnJ+iHfNCBMLMJ7+TOD5wAz3lDI9xnlLhTX2Sc54U1HxbgYQXg03bgt/GOf
SEcD+9BpfGinL80j99J6++kvc6sVz7MapOw1nHXR8sNwI4UrE1rmsep/rGsNrFaW
K7IWCz2plLe0tA5WfcDmjZQc64vhgRjAw0/rcBoVBTN4LN1O5IKk3gHk4BwyG4pz
V+85nFlPJ2gAmEmaT18unp0WkHQ7XXpq6AKshX7PEFyS2kdyJFcdqkYNsj4pcWFx
z9TWWApZ+dPm6qqrqpaBoaYUwxvg1jeVV2CnBfJ209Q1CqtvLMJsP5qbfQYTRwTp
CGCuu53n34Q1PcQRw1sG7dHjMGR1UUaRUFZdcsU++GdjqLRmHx1/Q0ACEIuNuHSH
3TmmZB5KwpstnlcWhy8MVA8gGUT4m9XtSevamVExx8pcyh75+CHFUZjf8bDE0wLb
aZlHYWcxyKiiBT9lgYuX/rVSsfUPk0XALLFK9NiEZyclPfg0+4GGKsYZ1B+on4L0
o/2A/8nF1s6FC2hCiU7xs+jdILXN8XkXrZLVafJFuhXJwG9CYOGevAQBev2Tjz2C
n4rshDOfH57bYeoWdMexN9rumT0HisYXP5UdmiYHGs5W5jvXui8WDPh7OUpgjSS8
V8AC9QeGgMy4ckXnO3QStSjki1BLW1M+6zT9WHiQE5W+bPaUzpd+jawovzSBokU3
Zt7/7MpQROZxpNf8u8jII9wKrl8zmLaOPBUa8LG4rXKh+sUBN8KyLA5mYLoOZVGB
kP+p6iw8y1oEgCXWytKxY8xr1pkOGEXT8JC0MrkktdCF/UkoU8HU4kxH3IvTBCyT
ENm2MNTrxDEL+5Uv2hPqlxsAqFNLQVl/bJoEIjRB4xGAstOTfj5EBXP+u451TEjo
X1eRpwH0huBC2O2Z/uokanqZRURgbV9W97yBGi53c3XSLBukdlTZlygLw9FleqQw
KRV/c2v3wGOt6QxF8boVLgSLnchYDrzWSQV0QIMHuexFlUAAHOh0BQqw8yHMZKpg
21NRAS6lwAkldBXmoVu5Q2K423pI0RPCbpjamZTkzmyiPex1xxlxt6Ih41yEu7To
M9GKuHiD7Vy5mSySQU84RxHWfIWE94+HbeQ/0Y+05LsiCIPrSz0KZ70O0hVpMg4Q
AUTmX420jMkByrwvMOFDheJV1BnXqMfhbADO/LGVCDRJ/+aclO1MbRODMg+smim/
xliBaTPucYPQH2NOfF3eXn/cOOnUuJLQOxF8EXTcD2YCX50MxMHmeIGC9YGNilRA
TGo4p9QwaM4iRqrgWEm9OYZm8etmk9NkjactDPdiFF2TGiT20ONHeP0BOi55EMQB
E8kv262AxhWTPyWdbjex6F4J81iHM5noA9wR0qlap+5vmN2N4BIwOgDtoTkt8BuQ
xlANYuU72/ifiEZK505TGTMIlWceaw/0HB3yZNioNuiiymtsDoEVJ5xaaerxH7A/
lwYZ9nvSslur1NPmtmHrPa3cW3SkNXGatb5PWxmmJ/eDfmZnLaGPR9AfbhcBaP4t
EtYwRg0uGq8D2DJb/+4meMMo2ZfH0qyrC+3135vsCzzBM90MoTLeU9j/997IMf9L
XzX7VtNwcmO9ztd/l2/vs0q5mzYovnTRTd55XdqddsjBdHYZvyWCkHvBlpAI9olw
wQYWLVkBmB0EUwFPa6P2WiNL9JtME3mo7V/TbH8LKZcc/VSQF9Vj5sC9lSNUfX6v
5r/8jbIN0OvgDnzgfhl9qtrt+Rrf1WgujVgM+v7tmj0fp4/HBwWvfc6/7WOUOCEL
hXNKVGhcmrCfXcJlT9+WYK4rYV5X/5XmpKKSKOhQ5tzZUtZfkU4yxmaVQWM3NEg8
whuC+nMdLsl+5PxNv6SjVbfamKWH0dXSEPH1T2XW46CJllnyi11t/V1blBVJPjET
VkHOAbytHmB4y7CscrkEreLmI/gKwSRJn36kxuHKG4t6CJAUHf8Zu/+UWmxYb1dQ
5YmCRJNw1JugoCJKpuoabhWjRd7AMzzNQg1vFHGiDxl9fMpcM2R5Ey0YXiZKJwa0
qzgKCb5p1bMVB9rwJtf8/iV+j7KIZJ+bpAAdcDw+Wbx7zrNJdxzqPYfjKjlBgoNw
ILeBmqC35yZtgL3FUTlMw0bV1yKX815fWrMUNAl7n1WOG+6yJ0HLvP4PZq1PzMa8
LL/lXlVqeabYCtnUA5Hv39v2dfX2tb0bQvCwCQSDk8XGbau2SdKZGr+n+9wKgCjn
gF2QQmbyTlyhhYUWZusb7n+7FjDKYpvVhbVy14tRX2LWyUDswu8/bCzU/Sc8WjHG
XSjGeoNu7wMKo19FgomVPBT7+DEHo7kTOr7d9YhcxfejPYopP1Mh85g2Tw3RJ2KY
e4rSUWRXsj3SNz88bdufrGOI+v6Lruo8/Dc3By47IyxoblNnSeaPZzOgIuSIqnZV
pwAlw5PJvpN7/Jia+5AOzcX4EAS4+6fqz2T4F4eAK4z9f0z2ANtQsUQYls92Mv7a
dn3KIZFM7TlC3HvecAbjgEh9AU5JBYcKFUMvgPx387N9u5fEQOqxw/AjKbWt5AN0
InUIlIanPph+mL/WFZBvZeQvQ64mmzCJu4tkkAfbasJSnXnU7hAZAH5L3cnu2X8V
QCgBfsOCI01vAiNQQAaZ6j8dYVdRSje/bLBx999yIHTKx7mUWo/4VCpZPtg0Z1t8
br1/9J4vwYMKzRDum6+DlkvSGQJZEmCFr4MFMqwxeBOdesVBn0dMi9F26tk/J9+V
zXgVReLH5ZC9rq6BMrd6NTgVjQtJ71zkLu9BRScH/4qJ2w/6Fm23q+LTP7zre3XD
p/ulBgrWvB7jiwvmokUyx7sAAinsbP8iEIlQHKTRs1RfBuiJljGIWDzbnsVjETg7
jpAhFNLdzCnyCrWShhrUNik/Hw9c6pySyrhuqPEtpEF51QE7mK5ef1jsQtNhQ7c9
wO+1PX5TWM7M5RgvbFeD1kXBB5SLl+0ZmhAHzYexzL2q7sbLfghubLwfAt9pzhYI
isFcKUQJMMZ9Hc+exsbZKRodXuORGSd9t6RjKVXG1A+ksCCWvW+QiYaX1HV1YTLU
d2D8VXzXLJvtulq6kZ7kvDh2Mdei73iKW+V0QwpAQPx0okiCE/EjpqFEPkZ4nBpo
BNCBJUZjtd3PGIZTuuKDAuynrWtWA+I74diKLkfJ/x6mRZAVFWZK8eHSaHj3skue
HdHKtbDt1PaHZkYGwkfsN6bLZ58gfMyix7GVh5SsUGIdRDT5iY74l3GOCZnMAFwj
YRkYmgtXjU5WWzib2MbUCZMbTZcVyyapdz03KqBxaVoAO8pqsERzGlsvIMJKeSbB
tu7O1CDCdzTfAppGjBf33t6a0wS5zoKGeQSUgq6eYRR3J72/GaZIsycoi4DQHjoS
cMj6GoU+NxPGig3wtLXheZ2KERMwTSKIbqlnLZPWUjVO4UX1WwV8RMmLqP0hg72t
hfQMY/HMuzl070AXYl47GaQRR/rwgtTCTJjHtMVf85dBTMG+3sagLXxjXDK63gu0
f45lQ6B51toc/CbvrIvKAio6hFjcrvS5J/joBIiEQc2qDkBpMb48y+CudftSJUDT
1TeTBK80PhHJ9OOS5VhGJyNNBDw5ne5zg6eceofYzoY9WSwl00dzudk4XVbGPvpm
7yfp4Cg0yM3Y+S9vMvIiPNsoOBaFNXbaPny64Ewoz+f6m7k/in4nVJyXZEILwdgj
plp3ujfWeVBxcVUvucAymo3vwi1+jvYKQner9QdNpo97GrnZx7vN+2npRPq4CU7B
DY//yoa1wpTLP8n1chO6lRXzwMet2IePmJQ/Oi68MaMeULWH6eGbPREoF+YVBdp7
cJRqerA3lRWV0XJm9wmelcvAqfRN/FQvQ/LH8vD1fvVS7x5mzOhMuUzGw1p165Ru
6c4VfhnsdtmFvfwSXzRv+RSG+f8RwDXXJvfi2KpzRn+lkVYvxUugO5tIq4wpnilQ
67ZUQQ7rOY8oa7ikdrYM2bNqu+DA57nIMct7tlpqUSnHs5NpYh7kaHeGYQWKanZo
7/jNrP6LKy4D6BEQPgavyXBM2Mg7OAF0vDGHDhq7VODaoh16dfSokorwlG+Drqva
Soje+kXMMYd27TTLILtsVfCiiMqkOr2w6ApmWuK57JxmG3/0MgQXGZ0w5uHmj5WU
JZdwhVrG+/HfFsqwGbcPI7Q2aVd002XcptZ+0FRWpmeMfo88ekL1PDjLG7EMAmp6
y5eIJOE0OtMF88j3aLqqCmyiyWkEOGE/7UIW/JJyNCQMlVJ93HCvoER2um1+NVrj
N0tbmQIgPyXVwT2CnnBocrZEcZutkBDvfdWpFVjNNeAIxLL/OguX4BIe3/vRYPUX
mowbbf3u2W0dCHc+7OhYaogcyNGJait4IRcIngtjfpm9xzlUdePQOswIEdA6SsA5
gsNBQAeZKXjP+eTyyohrrI+nVCKufcz37NmQtGP0ez1OBT/siki80eMU6FM+TuJh
z9D9cdwVGaGOAWrXGOAwjZx8j9eXo9EZcuXeD0Nvf44x5vZjR5G6guS3+kIFHZI2
RGknBrtaBRgo6X8wN84UEptEZuk7LWIHK3tRmVVYLNcgIq9GkLQSKBXguBgf5T1z
eaStGZTVKvRy4KS2pIit3yrXt+QfB4J92frHKfZAQg0ivOoUODafn2llqMlpL9HD
Jg6MUh6zJPvbuMeea1QOri1GvquEYiCcXJNPg/2yvg1UH7SRR53tfN7BHziL4E+c
BpapWFWxZE2hNO/U/52DfVHBLxmmWn593mC2fVrIB2FYnFVAtMxWfXUJQp7NtQCH
DYna4G4lBsw4IEZWVLt0ARoBHCsLqs0ZZ9ry6Y0/yT6aC7aaI7S+CZ449CoZQlJx
hty5EhWsuZd4lyxrYMINkYxXpKCMDuhtup9sP/DZQqux3a7rWIKjjKcYLTWPfK/U
JMSQbjU1usI1Ke5PeF7PJYLW/EO3ixPdJBG0xlK5KoUdCxQCubJJPcHu+2RYPSZC
7FYzwctsXJEJeyyMTD7FljUoHqZL/QYozijQFvB6vNIMO/WZFLcy3RN7TOHxhs8q
4mh5lQf2BFXFea43QKUwVUxnv0M0kY4E2lylhE6ogfk3APSQefUDG7ubebSgz47Y
iZ79wQd2jXqBPQmLeUoNiAbCTqSRfQjIGYP6xXHFdJ7B+8+FtCrXMB1D+R31/4Qi
VwvryVRg9vWlhOzPM0Lzrpx4kchY8EESnq4D002D07rq+vqdlLsFomz/DE4k0L5J
bWsaFFpnqjnPh3wf6NA1EvrIMZfe8zxE2LGX54DDzKmvEfNvhBlsA5B6gd4scVeo
AHe6EO0MBR5ZaNy66yVnoWYhTEQRQCISTJclsaabjb1GB7Z7/y6ypBDuvxq/8ZcJ
nOFn3HJCz2NrLZQ9+zmoPr/JV8VDjUT86gSFd4r4a+sddTKymvT/VCDFsJpFa4Id
tjViEEIWBF2p3DSAVibgVEttTpH1NFrp68wH7G9IuXNomO+Tz0nu5BaESuLi/AEZ
cob0i4OajQ1dv+8duwJM5Jo3DGyxDx+9l5zFzYCQjDDRtW4qTSYd4wd94WpF2FU+
f5+3TDeWC8sWTV2t1BSBzopmAMF0JH/9LTLBAl7K+0F35KiHCeajoipoIDZxGRw2
sThQo9kFa97M6bhMTM1HMaMA91/ay+I0DRhvT7XwkPq8/uzmfbgvACDN8s6glPSG
rYPQhlxdBLJEZQJK3N49yCW3kRJlxqp5pj3yVtISqIcMZCEKYHC3TytLfitA9VFf
997V4EekFWjMg9q+xjgHmHkjZOX2ikDmf04QzLTibhky/YhVdnTPuTFItcWhsz1M
lxDsM4whUAdt2EoliV26KM9Rofl9un0VI7bA7+66ECi40nSJiVHSa/SOlANV7aD3
2WqB5MwVgrRl6RX/x5Jc+bd5QmLQvn/bi52g2WOETQz76xQRZTKAvjQoeR8nvp58
knbfYnC0D0upKbJ13SDhNN+EswPVVQDRFdCeVc99s8vcdLY7w0HBwmGrWm42x4nb
y5bl87kcjnVFQjJYVuF6oUBqF9gGCAs4OAq3H9kpCtPwjuQJTQnmtK/C/Vk7nRdS
Exxud/uR/xvYYAw0y2xdzjJpDbCgyZLhvqWjQcenajOfM46z/pgwNbu8yXv4BsfK
hZbI9WFt4zAqdaNeaVOT4iiCa9UIxMyyBQzNmFSKTEn6T/XlKHykg11AF/LoUw7E
mmrNHZL3QYzY2RdKMDr49shlVxEkuj65SMRRLmNfDMWA9akkfPFge195sb81TYyy
JPr4kTKqzyz8QGHlY+hnHUNTaXKm4j5Q3MPGdOrki2khtBR1k8NODk/eeJz9owAs
p0uR2cPpBpvX4gYLnvs9RI6A0NWI5Qb//fRx9UUOZHe0F1BuLa7teIxlbkBMLHKG
GdVGp5J8aGB/hn0mBHXqQxEnIKa/QC2qRo0muOa6Et4bX5g3aWP2x2+3bV77oa2h
D9a9Sz40T5GRJHaXfXm/nf8PuFfyCPBSJDMnuHOZ40xAMSJ+r3aRwPz7lkJLwmWW
eLTbDIZApvoBhNvGFCefpIOYwkAm5WtRnP5uCFq+gQREGoFWu8dE4ed9dN95Np8z
4QrxBwPQfl+rBRw2ryjXgtYI53Q9sVuJgBH70esDEyGHjaZGjabJmlP0OEVvmeQV
MRNfz3xNUDWNNU1hrsxCNbZxvF6BPhFxDTznuUI8i9CmQS9/kobboIFNcrdxP6bT
l2/lij1kPx4rARhTtiQEtn1CJ/i83HfUl+0zy6Ki17ljiRV4E5L5530KYWwWbY55
3iM8EVByn1YbwpcOa59b0fxCDvUFqxeMFh22MsH7s6a6+GiVLYsCzvaiZtC3EUer
iuF+eAzsWhKu/IM0UhYreVIjjwanNdPTZuiNu9LIIy0P+gMKJzc2vpNvTFp2nqFM
IdbCL4NEKgmDiPddtQH4asLWvABU4lET9ur22cZ+27S/Yb8P0FG5DEkAH01MELHh
mfUX8+fib/BYRhqfNHUL9ix1OReDMH+QskknGbvQ//H20wH4ZY4MXRben+Vruo7O
jXJfR46n+9CW7f0+pc7Lf69GGq4ONUf0TkEoyxRCaPkBhreIUmudbj+iYakTjfv+
pzBDOhRHS9hu25719S01J7QdM4wBGXshzatyHA0os1BGo41dZ50TylZQtGX0Qg+2
xAk/y2ZFwUgud0doqa8kIQFLKevoXaHRSVULrSR6R6tM8IgVfcFmnsXy/ymd64+W
jPNVZadCblfH46wr1CGe+QwEkRw/GbFla+44EOJ1OcEEOROxOoBXY22C1fc5fpr2
XTWSZZwbcT1zrNOjLFoaTbTRwUw8vpkaFbQzmS2GxAUcPViaIg1tOTPV38EYL59z
XtPd9qmRGWwSGxYYX/aNNjpTyAveeSh5LIozJlakXzohZgquRy/BKHxaD+lr/ZwD
eE+A2JLG/hYAbFJt5fOQbxYxMvmb4ahfH/eRCy/aTbOcumyPxp/JYa10bbygnYvn
hRHMt7Jl8iOL6z+hVcF+2BbnF4lJoOr1PLthbJi075XD+aQVBl2UnSp5BYWwrnbI
jo9m8MkbL3Ni8mQr08X6F7uyAPpDSFA4udj9uErMxD12vkByK08MKIZ6WZCwOWOD
BOa+IvncMgQY01Tw3DRQ0i05RUdtub0ZT/bZiJanCRbbbvT09/ypbiUAjitdUXi8
DuVFgEG/Jc4z9Wh3yktVGS5GrnYobXA530BIQeEYdMYjVAOv27ymk3BdZEsctFAU
G6lsjubCajMdjYOOViGicgNk3sbJdjqks5ldaubPjMIbP2Mi3iZsfBuZD+vAibqJ
GHkM2YmyWLHErVTYPKLW3I//51iZO086ryoFMeJLegWgkwX2oYtfSCT8StlmKA9c
uaRJItPUE1hSTZuHVfaiMcFBO3f0c0KMbyGML7d8oo26HGkdhHNn+4AjbPhPdCOe
AKiiutCYu+nMVPr5BiMNjhxXrts3MBu6GUWah5TTyPMWu5pK5wo1DwvuohR/Kcyi
AcODnxAwMDdcbTPMka6MeWrAex2QP2RZgv3dtQAgP4vyb0Clvps2+vfFxfYt6pyr
VJzFWVKJZ8xfC8Qkbu3xIITBAoOK5j2cdGAYQtGOFCnfP5IzQ2H0pT10UV5t5gzz
vyVdWNfOVo5jThvcb058371oFEo9dKD3fjWygz6R5AoPLYtzTc7YaEvetSNsMHwe
qHFoIP4DXezyPDLPwhtXxxeeeERY4Fm1ZKZxKYXho8pL5jk8IFYJ3gJr94KDlSmc
784y9Z6gDymDtrIYUi0Q60wW2/BYy2gxPqvMSEGPbRUPlGTLZfbMORgyDqqGXvtE
frqvANSGIPBnl+ToOJ4MK4X9ER55sTUW+QGLn1G1wO33IO//2H+438EppOX87Ges
LMiQLObvx7B0l7Sd2NGNfquc1+P+7I9VR2hm+0kttp5/gYmWpq3BuD42Gf9Sz56p
Urks1bPFjaCVvStA8n/Ld+T9VmksP6gbLlGgBeEK7CJWop8kfoJhwmcHhxnParw9
SYP3S3I9fct1q7P5pe335JHhua0s/425s9H3ZZuEaJlmSk2KtsCUVsvi0ycJFkjd
d44FxvqEHO2qPfQev0FMFC5GQwXhHZaCiek9PvYxZC8wsOibq9DvvUa/HkQasoBC
9jj3XBZ0L0Gi86MD0ZzHKOzQhRyV0BN8uekOfTuPrEj9ttBujTHWR4gOIHS4VZUE
G3KSCjLl771EHpOBT3i3v4a8qJ7vdNS4H/487H2X6qiBdBy9BPtKzqMtOmLCvgtd
UsYl2gVvPV5wzzkWSGsaeL/AEr5jBU/NdqnSEoFcuXvOgCaQ795EFQEUfjycAgxN
1J1MABjT63Hep3Gln3C92fozSTO/++OIQTAWCtNKyjwmvpG4a94KtR645faoRvjk
mI2IVInRV3EZ0tl5Xd00DY32HRNHjJiWQ6WJcvG16FdR2BL4vvKdO2idLDWGmK+W
SXv2oCycRI1F+qJhGPhksVCoqCk142BUTX5Cg6vPKI8q8rike0RBkD/qFV6UG5Wy
w1+t0QpOsyQQYKN5GNXsJnW4/BbsmJC6Fr1yMgfZYRtXLuTj9nyx7BhBfCA2+iBb
G2blDoJmLLu2RrwD0fR/L4CMby+Z3V3ZNKVR/FWtrfAXWiHonCSgqjWOy0mIpNlc
vGl7zp8GBhcN6RzYJeuQ5u86UDXAMGhGpL8erKaRZzhWdbrOVm1JrntIgoIOKH23
YGg4AXuNrAM+ToqlcxMvkLrePtIjt+IEMyOpxQ7YOaVyystPHzp00ndx0ckY+QEJ
yiMGJay865skT1AmTAFO1SSMuwCgIrmzleIaAQy2ZciWxJTi6qMyKR/fZb6REYVl
vuGuHXMO93Wc5wr2OT0+0Dt73v4mbNlUzunAZW9JVn08m/ax5FAYTEi4GEmEbEXH
j7LtCSma3FQPZNsKCDCGeh7rhETOgKzjfWgcsPvuyaujdCCQwyWAbd20cOvSAJWf
wX9XK8zlotmvArl1QFnsklUVeByfgcFQF8jZT8bghBpVrCp/+5voOVW9w/P7flC8
gGTcLHG1+NEkhbYyPIJ3lEdIFBhmgOzj475lPz/UpcGxBX6nXJu9CWOS/8+6Hjnh
lU/Oo01a4qfiUlFPenq7LPWavRbbFiNG1mPfAzNV9qbUKRjhzqkR7qBUDX4l5yqr
U1INsAP2JL0WZG5JZwHwCheFV1OoVhBUUpHgiOQIwu/6j1j0cf9W3ida2dDueYBB
qblqnrycKpDsgMskER2lKWqmUMudwKPnEsShfYUH4BebMLVvteLx8onelQ/1ZElW
JVFETUfJn8u2Tx/D/v89krth4U90rMTk063iwPDiMaTxS+pWSgONc5gksniiXa1V
ZizlSfZ7zpV6XzunFMRrmtqJ8vlQQ262taCdBTbmWFhywcDNQnkBG23//9rMXl6P
7zWJdfmhnGbsO5oCfvH5zV7QxJdHv9XeW/QHDBZXzq5CRwNMA62owwS1KlDIq7Y4
tDdo+dBat1Ixr3OIf1TqST/LNeMYiXOhFDpMCCvv45La11iNVA5Y7C0sfQkVN6Bm
nbww/AA0WFZAsY6S89xdiXoObAegWnP9dKrzGbkb1nxviTOk0Uj5lhr2ot3dtq54
R+HnupU5Dvki195OkNqfaBMOju4PRth/yvPkQ0Lc6COF8+TiML4Xyqp86pTMf0fI
Mq4xd9JZGETkg1dKPmCyD50zImdT0EN3Mti5+IYUz5n/zviHyQGJ1uGoazRFSZdL
TUpwuRZe9ILObX3MIEAcYSkoFNUMhoqNwy5P+767dhkglaB6QyCIELyVK1JwSR6J
aArbAODGgW5XRdCIL6D++ceAfCdm81vF2IuAXEdkrt1UdaP3tsSmhFk+M5gTb/d6
LRZhRGmyUnGbpxACks5CLelPXeGBDKgNN0aOxOP4zBA+vQHd3Gg+fXU5Gkx0yWVo
SlyvvvZt1xCQR7oaILDBXIZ4bPzjIeYC8+2BHj7CO1baFjzjj0FBXFOk/fLEdJgP
5RYTGbz4yTlqbD2Z4Q7fCaOyDpIisgaHvIasuWl0khzOMi8E+Ou6KDqVLo+oNmkY
k/R/UnKR8DczLdyk2K1bupy8X6wum2JmFJBgOl8OajDbowemj42vTHbnfaxUtDe4
EC+geZCl3JzIj12xs/eRB7zr8zq8T4aSDTjW+UjHktz/UwVbUBYWyqxYBZgMXKbI
6+GC70bd6CiWqR+lr+mRayKvC6/VpL7Jil/pR+sjjZvceoi/T6VtVmLAI4di878o
t/ewUHhIP6tuzwMLZGX3ELnyGJwUfdjtv1TUwA4VGeT/OufSIvs3TPCutFqyDAXw
XGcN02cMEbrKkzWCDTPvAmc5Wtne5OMwudUzKQfBGzOhuPQaVloNWhrdciAtMgL6
kqycHo1BhuaRX2G91+reL/Yr6AJX6hvSqUvUBr27BbEdMjTRT3rvrZ/Yt7JO1TiQ
YAiTf2JbcQqKC2Mnt3PCWDswlj3srDb9QxKL5/oMPvsBetb7VUGxka2iFP6WeOR8
imjY0x9CVAjy+ub5bRGrniZPts0N1NlwFBIGQaL6PB1fgIG96PL+Xad+oulstLOL
fyZYVmOffi5GP5rxlmScjp9VMvN/slQWlSdhc7RPOX+fgzv+3jxCYk6EDWTgQ19G
TGY2PSdPbO9HfC9KhHSg8WItdZ1878iX2JM0rD9ST+Hs4BZJOWvc653n//10jggM
LOpSA+kZ5BIpOwXgTA3z1PwxXjbc8XH3QLd7x3QBfmDwoyFKgAxfxcwI4YucKG7X
IKgXtZVt8Kve2+QF/Qj09YroIUcJ4QDV3E63smmyL5KPeWI2KkR0MT40wjIDxZlI
V4Zlijn1jjwvI35ck/Ip6RBt/xLQwYt5stw33+5R04aQW1Z9siPqRCsAYx9Jbu3J
VAhITSuWB018cK9AOg1lrRenpnVLWIakpQrnoKR0GPwStTsDRfn42YkM0L3QhHUZ
rDmMzZHCIZhNNUMgd1PiIrd+shug7CWLou7uWnP2APud7VVgmkswbyoMVlwQBOpK
jX4Ms+wDNaKjGreAhZQTlTVne7/+Yzt7puce6tnRksKqPFpzdCu912Po28FxR0tX
xnf8Rk5PJGTO7idBM44hbbSWnpJKmYUFDPUe5gkmfhdKV3RmqcAKkL9Ab/sw8VU2
BJvwOmnIMfWd4D5uF9fbBraXB+ct6LT38KsCaYfj25b1s3297x2Cf9BXzJDFbk8a
B/d/QUvX65qOxCy//SnVjxnG019N6SaAsypyeE1Ub0yca2vtNNAoI8CcE1hhtbea
gOhhU1SP84ttZ1LKZ60LBqyqZX01/zRxbxvNh6oW7fnGtmYv930hcAwURl1b+qHO
QmuSnvsuYxvAdgtqry94rXE7tN6IYwf3wpp1VWYjousmI305wHNjJSVCJ2lxawUF
tfOBkqNfCBYAWmlorfBGhkSvKUz5CelN4TkbutBrv1UA8tiFcBW0wfiHFlDd+TVn
qmW2yn3i4v2q2IJ+yYSsSD2ZtEK5qzCJB1c0+aTGajH1+YH/3DbD7pD4iW1ROT+4
4ui//GH4FPAPJc2hOJ1QrUtqfvN+mSywjqEU/iM2441XfHUIU/L1wybaAd7i2Xgi
LLwgfBxnD4C/46JrgpUBrHU9vQTs4xFsQdBXYL3/lDIJBRp11XIEIUWYu9WYZgrE
07wonsDA6xmDYSrB/5SgyUCuP9PPfvQ5Gjk3ip3Pr+zOIpSeocyj5qPOpZuagh9N
6BA0+1QA2i/DXKxyg76kg+SHSD3+n7zG5NNKCaQ+elbEuXlbG3kOTA1/zJOjndtX
1LvtW6xkCo5S8EZAZQhk/EhykbKtyol8Ylzon/IPDetCs7aVGf/xEyoGaFbqnI2E
YPf1iHkBeB86KT2z2RmpSZb08UTenNpaZSNaV8/tc67lgTStITzUgj5xEfmhZP1+
VT0Hy66jFwreJ5rOKXgKAKaz0E4leYX7FUEqUVw3fzL9VxtjCxz1JhNxYtGpHZLy
aBvFEAJrkloogFFdkuSz8l3Mh4wgMzv0mZr8/JWtX2LO67/VWO9ooMnCYX2pC6QI
rWJKbwUZ77lwU291HIM9/kXakOAcpj+vWeRa/9OkOsc+UXyAnkdQMsIC1ttteagA
KulChxDnQpS9kNKXwNrwcrp0bB//edskSqQyRh2Ct/OSqzBDJAODTDZG4nenzD3l
BCSkD4+SA+s3sEkHwN9lzkC2jA8KJcdlBTlrjAdqrHeEvgHIjhWMSPDsJEqqBFYc
sDBR5scWSRN258jB7I49gJFSW9CB/5hsCUawLKN+ClIRxXx+cfXfeGnWQOtoM2++
6srsbYfp68L3PpDfzE6fkBvKTQm1BYHwzcK2FQowGOGahVs9jvJ2dr1DmkGID9Lz
lP2guq4MjzIBP7BhpBeWPofyuhRwNlcY2E05ydV/T02pFGQrnqYLVrfYIpAX+517
DXwRU4yqgIeVBiOpEqbUNo3QfM8dXMqIqJuKp2Pe/soeG3O+nNC4waqijTnnYYyW
zfeGAhjc8o+X8OXysNE+B/iYjr+FmpND+7LEsMlXSyVLiiW1RTZQfdQqz0qJGaUg
STL6qwRYG9+TXdlIXReJz7JxltlgUnuIfnTo32Uer2razaP0RUmd2z7XSGSp6S4i
KmCc+QkIvg+7DawM5rC81UNYO8EGbb9jjf2QUGKY/+xjq/4amCRePGtWgj9InlJh
Hqb0nkX13QeFuMlneuxI0WRja/Zs+uMEfl+jXY6r4MHgc/k/+ZVlCTWw4p+JjUXM
hzRvYhaYEWfPdGIQZ30D/kuWdlhAqV79ocHk8l2QgxGuMMf3wbCJL5M2961mCtrl
vcfxuZHqaHCwCF4kGKqMStmW1SVF3DKAoJ3r5OGvaQuHhdUcO36XCoJh74zDICYd
eCrV3l3usTwWtnGVs8H6Feg1eqc/RY4qP3jZ8M7581Nag2jP0nKXHZNvSVBxb9aJ
DIrCHTBTFECwws04p5s5BZWOQyM8SpZaZnrnjSXtcZRoUB4F35uuKmKCZKmvSOYG
kzXevyewSXwBxqR8T3DX20F++vIVWpk5zZaGtM7XAaqgw+TqBChmlq+q+ClZbh/f
Bqvntvpy63D5N9g3acn3hO1KwITWEPMI4ottBLdJC4RxgCBgqkWo7iaMmMrgTwSJ
EQpXdNCE8AHk9KGgjNrJ4W6bYOO1cZKHQH9fG4GQzzXLUPYvWa6OoEHZPFPPbxx/
2uW3B4fRWWl4jhHZ8Wbz+SqLbzEo01yw+/m3biB4/D6v5zAm8w90nys7O6Cgzgir
69C2f2k/r8gOagEcA724EtndSCxZE0hKTWBomlJ3EX3HN+eMZkaqL8s7WTqJ3ib5
DfZtsd7cxBOvCESOOW50LEEdteoNgDioXj2Lslazw5FF5ceq0JDLRjtrGzmXtiws
NxyoDnmdnr8DbarbOHfeLc5om7Dhkvlj8WoNrmWMY1vvspSlCcdZcLgtLUgezb76
ZyGzquSDo2QJ8ncloASLv+MAnlD80glfvhttn4BN+KKRhxEXLwiXDUS+2S+qjjXU
96SCWkKWa7Oz3jOiQ/hWqmNyUfEhLHjW4R6/A9j289dTnjzsFC+3srmoq51ztTPc
jiUC7oxNQvnx3F+pNCQAUpT0Iq+w0msOO/TD3977aZsbVSojErhaQjVIy/bYMgCD
bwY81It1ktF2hPeFrtJUtFfdlLx8nfAx4rpCJoRs8qDAqM6zVh7bh5oarQgrxZ0V
iNOPDHArX4XXpmKG2S3x5dY0WnVWPJdc05XdfJa9b3nsuBaZjmmLvLPx4rxtpcgs
ts+vlzBTRLjxjzXZbC5FlcIsyzelPTji0gwxSgxYEuiyRdy5cRWcGE381S64Q/xq
iNhEW8eAiB7unc48o5X6+m8BDoUDONIr19CNOCi1JnE9nqgO89/jw9lYKOsJbDRl
F5hXp6PdT9CiVhjXXW7RQiZu8Kq3s5o3XRAZMB4JC5py724VI1HYEf0DHh9IzqKy
zkUc31bewOt0KwFExEUBd5rC46waaQnmGfFwvacHlfxnrlwOOt1o1SvIusN643/p
dbWWZS6LyWBFmgAPT//OwHR49IV3p4GLTVPOdA8+Z0IHuhDUP/Zl6FtZZKy8QsYW
3FWW14T7dS5lgI1mNT7Ym7Y0M4DqxgfKY9hKUonHmR3i4C/itX6YG6Yy67aHuuTD
nF+87PWNLO/TzwrOSMoP9+qxnrW1PWJ2bBbyqEEK+v+YZ/7YsSx9nVhKlVZu6/Om
NEngAm9UwL5ce+n3T39/hAmPn86A1mY4rx61lqwixB7NuH7ws2CVBtUgls7l7Sxn
4SKJGI+qG+zb2b/xOJUoZs6aOh6HXql2RSUaMc3hp111DcGM045Dz9L+e6g+yru5
EFX4x0cKfx+NszbAEHYQZ2b5Omf8PzKZ11LkcFeprgvLR58Ox66/tAG2DFnAhgUA
OgZBx4U2EnW+GgycFdyAfyfmj5ASkBvpHKFCtaHN0MjRhK1LAvBg1Y4bVGZF0rBT
zRlBsq91dmdSwtDqqumU2PM74KY3fe2E4LOgu8zLa80A9NnUKQUu92dq7eTcQqNr
iA5uivJ33hiikBEkM0OGwXuWP7olqwHb/CC5lG239eZqIF5WtV8b4oRG2LaEYeSh
UayzTWGerxObcP1rOIX1NI4sR0od04kOsbV5gonfiiKS0+QGSWM0NnQMe5mZEZiA
55UWAfCLKDSnMcsBH+zWHpILXPE5vePDOAsRa7YFz6llCDoYHN4Mp38axbWP2h2i
IpYaltTVFBcDYaRCtPLWSlaSH7yzBbAmlQQT+IoSucXzEEmq91haOsTtOIBHHCoQ
Tw/2b0jpQDTHuaODuvBDruv5ycFLb8JNiHMuW2/R6jnZyQOJLjpNKHeWovjcrxe9
qx7cs3ParrLDoNVb0O2Y0dy++YOqW98gSbelJT42T6KAcfjF6Lb5bvAedZMwXKZ6
0R+pqAkj56QpfUg7wVAJBtsn8Y13GsenmfmzaM0o0el6C9HE9aqYF16ge6FFfAj4
G31C0eq43k6g3PRBL6ZiARo1J2PAECbYKrsSKoeIYGSEbWgKzOTcU5LEnGEJJwnp
YMvwU1TL2uX/b0HIDgZ90EV5n1WsfQLugMqkLW7MSfZYj8akG9otvq6/UmctqRto
Z9a/y5vgPNZ4x9LMdekIvXQHeDKAMBppKrmpIES2lg19eQ4eT0SxvplhNw/l+KGi
eqQrdhBOHHDHiBlFzIX/BoD0PU/1X1ue62LEk447EP3sv9PimOMnybLInHebAZuo
v94JPQeF6OkECViWMfLDYbZ2ba4L11cwNcs1wIhBHSvXKzkL9O9vmC4iW7geCeA3
Kn6sHApKjVC712aNSlVtc2iO7X9QJ6EJU63QD0vZJ5jxdaezztuhllGAj5lBa+Ep
WZ3qV7muMngysA96kznOzfHhVbXH9dcUkOIGnnjbHsMhjBJS8iFT5gWFkfdw+jy1
eLNfKgp+rCbaIb3i2uPD97BDd+6NUEyql0oZZK4EbQ2GFE9gI4RDkMVCEP3U9/IU
x45K40n53OLW3MRGFj/5zDecXh4QMSwnVPj5IYx/4Fw41tQooIq2kQXfHJYKE9CK
Zaq6CTWson4lvQrZkiJwQz4eBOGrzkq6KKDyLw3PXJYW/HqukN3gLKC+Lu0sJted
6QIhnpTTMbiSOh53PIWDrJzBClhwJZ9azuxTJ2p5TL+HTvNSSPYnOkT9H5TccnMY
Df+EHPbkahOldqb2GJizUsQ0Qd22I7fYxno3nxebnMlH//W4esYyypte92YaRijj
cC0ozoxhrROS6LuUigV7lUuDAj87+6WvkTLw+IDRhJ+IhIOWVpq0GH85WXUjVLGU
lWPL8hM3CvJlcQU7B7yiCirpMiux+3f3dY3kkMS9H9f/GUTKAPSmFYETK7EEelJz
C6au+HllWIlXqhQsg0MZgUNaFzRdRuGpe+Hs9kvqTANXGltLnTcDmRNZMbsN22rE
o/DZECiX8RJHq0tIUGvyHT3eJlZGgjoQEO4ODUjauQkFdL8A1zH0cutYTtfxVvG3
xDcfRmZbauEGyHQjQYgXKQBIAeoIsJuIfh9j9SXP2Yqpy8AlJxqv4CKyjWdsll5T
D3nuGXZel90UDhDZZJPofIxWRBVVemER6DYuWfjt+u5sEyRFD/jwt15TSoQEsvIq
O3csnCxswesmVLgm9F/2CxCorS/ztxET+f7H5o/Bw4KR6HRmfd+dUwelKoMsOWnk
KwaQ2/x/R4OY2yb32FFSr5QxXgR590sLdofvNVsPUw2my4a+kxOQKwnZGEuMgXLB
KG8BvpZPSqIVlpypGvk9ilVz28fzvprJir2j0fQmEghhsuSGqdbAxhGVCx3tszXS
pyYCMe/RGxJpcS7ILsy/AxOgWfWllVaYWoo4rtigpBxTEsZnW2AiynqsijKSjc6Q
MMhwnE022o5Fb2nULkdcI2v6LngBAh+iEHFFwWNYFybrZiiupBdeAUZDCt+MMbYY
0wW6urakzlb3nHT/1un8IWR1xPqiPdjUAzQlpUa3/k4SI9RXRfiuAPNFf28Cv3Rw
kXFKGogf+fvERvjFSZHl2Us5Gwogs2eaLBjcVJkyGiWXmK/nfWZ9BwWnwwoSYBeo
1ehro7XdDaZJFMBdeEOtHR95tVHaKAoikHXJZBeS+Gcg0ekeOAEl2aTVmrkGLXgb
9pcJTxtRIfnZcjr3k5qx/h8s+HndhTJgyGo5pVnpeCO9hXxNaydFMwr+uYrbSFke
CWP5x2v6LlzcN+jMAspt+JD2j1mHZRD+pxqqMWLp8iRzqkzMvorhpvzLK9LU27ZS
hvoxaJSpq7iUQbU2NalwysYTq0RKtrsRBOd/PEplamfyTVPiugAIn4pC5uwWVQ2R
TurLWJb2h7dwR3C2Zmc+wqhvgNSCwuDsEN8kLDRaoXxrUajBiaV3+h356Ve7HAJb
F7ifTIgbWlqQfv3ViphYJpbUGYqP0bxYCmaCnO2QKP44/MPmiHOgoDhooL4TjrFs
/B68ANZi49zmaj0S9XMI+uBUnvQ3l965h5Ds+5tf2RqXGoiR/M44AkVYsGA5bO0R
isHWBgwzqlnuXPkXq3spJpgyhp5ooATu31n/Vsr2tQy3rvT3/XTOHqEny8noyFQT
PQxDZJc6xv+KZAj4ZZVqGhrDI6ahK63tTm2ii3/C/dgsa8BTMf4AtNAVprsttHal
PUPJJGlIgIuWwaFMb0igUpKkb+TVBRu0Qb5gctbFEZ3Q8yznoAiIKv2Pp5Pnfqtg
iP9sWSRzh5Yfn528YffdEYgqfmMkRY6q6JlVi5hzLLK02H8XvvfL7jXzc+WjCN3K
RIsf76z65kr35k9h8pKb5CdccPQP/rpa9VPw5pjP0eAG7xBVHcRhw41FerzFdas0
EnaQgLZewfSRDTWYJsdGIPpPu4+X0iRx7UdE0yspuVRlk+3bPMCU8OMxM0EGfkZf
wjUIrdN9c/uH/OFPWBMU95Ppl2GRAGTVYtHJsA7i5NWptX4LF/xyG+w53wNF+tXx
MFbIbLCb4TPAk997gMBLLyR6xKBcMVxAb4ve6WXKKQXZoKEK4NjY+RIyXQLA9f8I
dKbfMgNk0G7Y21zR2aU2I3Q6O3JckX07Be8sPeD3SysFGjUUc0dKyKzq1mu+8coB
HtTBglqwBl3nBup8HVcKYRhHX7mWNHU669Y61h2oGBhpU0XwmvToKF5JtoWMpDoP
HxVLD3lUURSuH2euW5YWirTASpePxHWC2HSYZ2AbHsTDdawiW/OhFeph8N2G0Pbe
1w8ds8Sre88JrW4yqPcpynNpvj2AEO6dTdIfkR4uz7jNXlaAR6VPfsTdp7PHlb2l
HH8X9owMNNjSQnrN4aUA+LfghhCblM85hmuRb4V74z89joAV9MDk55EH/Y2aJKkh
o2WKJyeOE/5rs4VikKkctihpS2DMqBzjbtlRgSNm3BcUFe61vSriFWTqHml67iBS
x2T6mGD2QNmOLapld4ekbNLlkVKYibL+xO793KlWriY4W7bxtG/VMmCnv0ZODVlj
uuytDGWwqeLauwLZdJnq5j61ECnfnVk35sLgrTT6Uae+oTGj7GYLTX4K+08cTXS1
Yhk0WDxoNC1CGu4YtjJyPnCYyBINv/MDoH13iZVcvFPL8JnZ903yH4ltkEsFrrov
M1y6elvtDWXd7MqeH85x/iGmSKSQ2FBPblFbg/7ecbZ1+QSALBAkJ1Nv6myy+1dd
zaXqKdAgxAjTyc/qhV9lg+KhF4Ps+ZHUmMeFQ0W9667jWe8fph/QA+QiTTnDtnEg
aYIv9gtGRzLp3MQYiFUWcnvBWn/1Cd7nCYxwQkAhIdVKk6J6qCS6QHx5g3crB5z9
2tdktvXynUQxg5lFnYBJk6hVb6zY3DiohLWvtgZpp9zo7zd+F6s2w7zOIXSeoNUs
0kkR37zdVh74zwrLiDHnZu2RAPQ18tCOyb11eBpSKlUi0a3AcyJA5owh5TEG1VP7
iPBBd+0f9P06N8ECj1JlYlAO6uMxkdO97th+OVrMUq4jYyQBioUnjDHBvsWjq50e
yneRv5fuJP3uvlqgBzlfyUiH6Fd6XKQySYqtdDvxDC145m3uAUj+Y3Q7Ib0jVzKL
Z1jgwca7vnrKlbvfrgip3MvX6kqaCrLT5U3P50TnPCept0XTmLfVd8v7BjEfOU/e
B8vfEP8plc7v/+B2pnJlIKAEmd+vuX3wY7TbQMWuQJVCgMmj7Zy4jOF80c0a4PF1
AHyYocfhyzH2Dvz7fOaTM5nJ28lStcLlKV4pa1yabdEH0eXZHCOqzZFYObNMS1eU
IAof6g4Y/Apu5mXcvrfE9Qles3fTPZAQydj1926p0AT8wDJMe3q9ex28l6nh+dVr
jCcefnaaqiObGdkHsmNkbMcoxNFRWvWqPrAK3XKbv7Ex4MejyKma2pdr64OHfJ82
LkTq+md3bCSk9T3BGsEppc+9Hz5pc48a01OrI/lUgVCVeMK/r6OLwjhHRJSP9rxD
dWEVORxXTvUHPN31jp48rA7AMhqP3jyYzKX5QAxTSFH33wPKluycwY0K4rnh2ntr
6NzpAuoMbw+cIRJa12fXQNyx5aU0/qJ2Q+mDN+FCVdmx7Hy96iMFWUhrTty/cr8m
Qxe/lig6302doLghwBi1p3ckFhhONNM403ox4fsojSEFWAF0ds2JRuBBcfOYC2td
+03JYPZtG+Hr55krtjHIUKZRptFgb+KvvZVmQVsatUauJF/Hr/Xyzlfd3ePT0F+7
FVjVMy5Ik6mU9T1NFFWe36fOAxRFYMX2kXvYVC6Ia50WBKlBCVKv83Yv4MxK8aqy
prqsCIOXnO9qS9rwj1x11CX7M52AzPQGo4mAtrEBVJBh6+QyMd7SNmPRU96ChDow
n9mBfs8uutGVlBSCiToZDjgsmQxlS4oLz2+uGoXgw7JHlZrmEQc3KBbvmHfWAMr1
8lga7UY9hjvfK0+6U2IwXeH8fDaypmhapXp9n5wmyiaq322jcY4zPVVkMYfI8oD7
Jw9ZtKtYPflCaPk17LJLFudLRjnqwChNS0Eom7mwITfHA2Ph40CoPBuGZawMvDE1
wG+qfabSJFLu0xMDBquotcGH5evNyBNUI3VaPl6V9MwiyGYzUMy3eTgE2gKUqt1j
Kq4Em28SlNT86temeVXaaZDcudxKCQVRuNl4aV8oXve03MgoLFsYjKNZGo6mT5vG
Re8YsyPaFdZYaaAu4YRsxwgOvr86l9jOM53mKcr6mdCRErbkyv2MTBGdrXeo5XPJ
hSFJ8I8wK3vnmIZaGsChQFd6dQOYhPTc7ONdw8CZ5OD1BXs78dDjOQl0K73yZXpg
0DPN1TCkC1F/AdiXzdZw8vonAlCxA9v0QIYISNOXIjVkHKTqUcVvT7RoS59INrqi
E1V4fCyHVBW/Qvf+aEuLNpV73uS4MkwxaiBcg1nQH1fPoeapeJlciWCY+hXFjjj7
xKXGuBZdMj+tJk6AFLzm35wAlOnnenZpoW3cFPSVl/LKHb9jAkwoMzVkXx2azU0U
Z0ueH/cTH1qPWUAzJ05ZPKNtWldcn7vgZLECu6xmxD3x3LLLYsVyMQj2PozRwhvW
Fz1IA+UiBND9yEY/H5h8vnpJAZ2cIXJ3iZa9xcB36iDfdnY7VnsQeerOM3AAuHEI
InnMvzUfLe4sL7xGVRW3AfSTk2SvUqswz7yx+BjaImvQ8WQdRL07IgCVOnDhFFcj
d+jbla+3KmXncsQFNVIRbUdDboT6N7FSB3pmDzP3VE9Gm+KbLvI+ur4KYeT+sD5s
BLbpUAtpCKIqiDbCOkDJyZm/1jPGtcpvu33D82H+blGji0weh0iuXhBrwxy9GFYc
O68ja3oMlXY5US2Ex2kty67j0uWZzMAtGsDJnAXWs/CmYFrL0cWBl0A9KZIRSkah
99t2q6GyEb0JsglPY//HE+wIVaANJG5CzHg7Kyhqzg93sFxxf3N3EbSSoKmfgp78
lqJggEEmo9GPYBCb06i0YSoNy2dhBg9Ks+9Sd2qC93vopzk5CEdj/fpSKa1Y+4jM
WF/+nXANqq8zs5DG63A8rYm1A2HCUc9W7sABD0STkutfmdJBIiP9e0jRi0xdGbEn
DXiWV2nVFIHjfpDPmCyuyNKm8OcNVicMwuunOflchfOGditNtwpgkMmRtaGK1SLo
Q+sENUGYHWFUzGAXeuOnxZdDONkCEt5aJgp7QDAZYvHh8xyANgtVQHamjn+VfdbZ
XJOjPsyUz6l4bMeolJ8s9u9uRkgCk4BMIhFuttGYsZ4pILifbVq1+kR7fFo/Flkp
tjPqO1yzJ5ba42QRvhQoyohCzHukgrc2gEZ2YWs9MyjGsaQz+H3mM6255BuCz6zr
WKXek2bEoqwUn87IEjrpkjlLLum3OCOZ5F8fu5GWdYM2P7s6jVnV3dDgdY0mh1qy
jkl8owdddn93aq4EtOqeBJ0rbfzgRGVKfs5HrPDMTydLaKtPSX1QWLTl6+Wo2Dho
zihhA78569Npjd8ljw6ounZ5A7ogyMF0uNNyhzKUELmp2f2kMfrQLi5zYV1IRTIK
hGPtZavKGTwS6XcjDUhSVfocN/ulBw/YnpK/sYfSdnHVn3LhHtgvwkWX4usqV9Ln
uOFGavIWC9uZjvJJOICMsoHjaR9uG9YUvttkXRBugAiAzHdoVnNA25X3NNkIazzL
UMcKfOLoEkzmL6sAflfpg9XvKjvHkEndOgfNl9mh2FqhCu+5lT4OVwCmzikLczl+
n8aOREd3MqnQnG5bBdlbHpnBeyzrfGhhplyRdkGufkDto3QsvOLRzPYAUSKhhwzn
KH0YoC8nK8503S343wT1caUxsWfWRnI3v0SYGCj9kA6RVEZwVbjCf3Jd3YoOFwxd
OIO2P8fTufjhmkA2cKXO/jwC3Jd5XmadkGS9UrpeaFkyqY4SBOqYkCQ3Hcc94pNx
XA9SMo3fPtUiAviKbGs4RgInUnc1ScVMK0S8Gcm+MA2ewcvzPxu5AagypyTnpWJB
+b/j7Zl1GQoJWXE9j5z3GEM+ccGp2X4Uk3hcG7/sJER5zzsqJqYVfyuHo8O+Frwu
1SgicuSi3YyFrimxs6Jt+jUFhUfpnPeEPCp+kAD3Ol3U/fU/Ly4ScGLUF410bK3L
rUGunmBEnlWsOUH25Vh4EsQGf3sRlaSX9iq152L7FMRWaTgSfoFq1WZ22TSPcDNA
RnZeQYz8y7IfVH/qG5c8Zz3gRRUnmtkp/Ab8ETlrYyuPKZfLO+rafBZDJUkwdiTh
5J4YvuxuIctd98swJWed8I/Br+VRAcumMFiv8nD8SKvaK+BViiTnZzR9zRT1hFWI
OdZeSDiZj9afcoM/F6DaEFzIp9POskisPPtvZyY+04hXc//P8qg0CRiKJ34JH7Zg
/EGeLDcmoUCWgY1r7TepFAK3gaGU4zbgUNqvxAQB4g3bJviHFqLGK6uEI077VCwz
NgnZqb0apmG3nzdqDl5RVieqERxzIK2e7v6lxcKn9vghx7Ubcl4grdqNL4WCN3Su
VY5btIHWub6K/m0kSmCaKbFG7gu2sn8VwMVl0a34U5mNKXNpFqEw25xxwLmdQ+e0
vLpzdK0dXE9Y7C6gLSLbOIeTrxf8aUAiF3meKog6DXdbkqq/2xrJMnAXkgsMDQpG
2F4o6aR1jbc0wNaUbTseGAC6K5R2l9gUxOOh6lRuklibWS4MCQsj1ljqEYf6vkPw
JQcl5ib0Gg2ILsxEhMV5XgibVeVA5jIzcdD8STPzi8CVD5ck8Fj4Mwx5eYi8Kj1t
TEKPvOrK3BnGmRd4QDbOEpyIkdywYmjqEVHb/TIVhz1zj2V8TZDG4OJ/qRXArjSF
pkrrPFwFoCx1hhArKEu2mQr08+EjjSgw+Gs1E+hycnnvTwp7nRNJe1pmWTAgkols
OYzYzZU7ZG/kN5IRCnSDMLcNedV/vs/OQq/MczfmmdY7BP4s5vrnYpLsXgUXND0/
5g1G8eqweGGfQkmFJPHadsFEnW5gCzNSlwCygNXHnIMgMZkKwnInXPXazmEV2sC4
Nvm/CuYVbnoAmjAN54vv3CCV645pUzGZr1DySSST1gwzO6NCFAxr6oMFedaWwp2Z
cS3vwBlIB94xl6ozDEgTrYy6PIQSOYoYEDTYxQcvPPmAFfAwFrGwkTNE3HR8ne2t
9UIIi1wEK/UYd67/5xKisRbOazTRv4JMD6Nc5lp/Im7CU+llV84Ebpn9A+y6DURz
h+P2Tfprn3V4tnVBfpyndgfib8wmeiLLuEvWXiOl+xp80D/mWvQjplIdyssk4oXE
1XB38LtOeg0YLwWGfbqbm9jELsfCKRxamfbr3PtHosBm9YcxrRsf3iGT4WkFaxrf
OED0UowTAEvyvugZnpGL10V9x3aTU8c0tZGCehsznTv0sMX+afweVA3568n1LM2j
/gZJvOCilYXNhKragYqXnrmQE9NfC8JJB4AuOkalssqL9CQkexxV6a7yN0wMgyaS
6fsk3ysNkfAgUhzb/mUlQowA4bqmOm+FXHmrRH5UsSNQ/+C34b0JA4zFUvXsS6D2
zlLQCb3+gTTnV8DUbyjF/ZOgLzd4FCFvCMaHSQxzg5wqSbV+by90ckYQ2QDyJqkH
lTdV7BO2weD4edFNrmY9l7KrZunNq+EcUxVE9Zq9rUh+D1iOOV7vDrK2aMMVzcdQ
Rv4NvWX69IXjLb+58PS3O3rtbjk5JYXrtxvpvz+sN3dVdCZ/cTQsPwefyI9RgzuK
Jymu7/GUj4DPhczDrI0AcLrRZ2bruPb4GkVZRdklAa9n8CxkXSEnRHa2zOIBqJ7w
t1e+EGSBHb3C3yoZMIiDB7lJIO9i3Q+BVDuW5v4wxcrTB8n7W7oWfsB0jyo7bOp7
52DjPTG5vURL/tWn8Uz741au4UIavMGdMzKY6r6kyi5IWijwMsaP736xX0f8z4b8
E7ZyC8TNFOWSOJX7dNwuyc/r2cbDCrR8mez1dqyN2DCAPRiI0gtw487C7n23BhIW
FPdg85b7AjkIm9064EtXpcq2FDv607ZPBdeCz0q9cNKVcJzmtL5uc4wo3MBgDnh7
lJ29B+Gim+uF19AJd6GwBK5aAMY5GgEdqhAf9T6gFpkNVcS6c/widCXb9AhOd+5c
Y9M28stA1eS0Ev7NUeblVa1gpuvfzxb7ztmhwHVwW2LZbstcF6JEL7E58hFSH49z
nUEdGLiPmisN42ckkf1CIx6lfUeJlMZF8NploO/MZx4UE4iSYVQbASTEXnM6tFgg
bdBsb6Q0LXdivTaTRG61cKVGv6QSAvRvZ7xOywL/3gs2ufPWyON3HaGj48RrVfju
edAbSUY5bjmXRkXtW7o1QFxrGZth41U3JBoqySTbWUzT389p738toR1TOWaoiaw0
T7Apqi5WbUyAV0tEvAa+XLRjMZxb6Yrdhz3BEyU8HZRAVGPFZoj/es4/SQef82Ca
TYmXcuN75jTW7qayDQUdIiX5RNlUOxJiaU9m0zkh2iaAWFtqQ5z5qFHEjXgJEb8f
BZ2fHnqGWrf2QYtWo+ONKWtnk7wS3b8mmuBjN5vF/phAan/NiSA+ZKX4l6S4ltbX
kGSnNTmhiZ/eWFP2Mt/KybRwaAvccmlyR//pquCiOj6xQKD97KuyofsH6hKT+T1y
QYEW2GgIXcQuzxV28F8a1J5NpruSnI+bUgjHVQU+sw0gd8b58W7b2wDa5Qyqy9GJ
At6fzPQTb3SYSI3mDobF+HuhXG0YrORzmMXgPOiCRLJaR0pt1uXa0LaCxZUELpTg
OQinsxJ73RobSAZINQxQrDQU61+Zx0OVErn2NQ594xbnrnhFmwf+z7HJoEHEfrp8
vE/Y380xfffB3XqKUv3N3hpp582wgWrvCqbat7WGYE5rx2aeACMYNXMnbQeh+LH+
zxvag3AThWRJIi/He7l79mr9hvbDKetVuymApi8Y87w68aXcEQaXqRHquUM0tvGX
cflXgRjagO6oTjhspz/zt44gxsz+lTUy7UDJD2PAIMH2pn4hOWFbO/mahvMCogZ8
bdSkCml/wBfRVlo7LhlNzu8zywBhJVXmyGnWX343bnmoppos2eUpPuMy7vwv3Hct
E7ZedmbXeAzm0HyBTjJOojC1R2gJds5n5rPp/QaIfOy4X4BcIVZ9GOjKcHckQ8Xa
9ZBYlbfuGOLpH2s0eRetYuSjtPysNcNe7ksa1weeR+h/XVUR4CHGFIZTpnnLasZt
sjp1pDsChBJOHQ5qcMcqS7MNxYCKY9NydOCC8OMINlt59glhWT60/N9OLO7r7wCk
DkLbizfBzmwHYcl07Fgano7EWvV9E9dHWJDgzbQB3uQ7XZ2g2dvtoQfKARAn72Ke
AswMC/4Tizb1mjbfyfS2aoxYctGFEWKTTr6pTDp1f0ICzRb9VT+ggexxaaCBPNOK
GaY/jT00oPAgHUuiXw2BC+PzG2oifWu6Nl0jXzhE5k47gZ5mf8tgiwE8TwQPCLdv
zFATTTzWFNPdqbpIhslO3uNIq8LCIZczuYnjMu/M8Wz3qH1V4bhdADaZW06b8c9+
XFDaqL6fdw0g8ZkBUal2u4eP5Rf8dLIB9h6RKQxq2NWLUa5uU4OEw0FXMHZKwhlI
uqn2rBHQ8Z+Gkd68PWsfA4UDJhvIUyputMwQY7cvPyfmXgmsG5RncMG9x1LEgcyF
AvNIOb6UoxckeH6bkC3NajH2wOefR7E11eVHBnbpgYalBddf1JOG6yVc+y8Sjoo+
6FQ+Wb0wn42WzsFbWSyN3nC8WFE2JorsrX1F6+wzSasCWpLyZE4WPxG8gTU6htcG
fwZ70ziA+sqqH2hTMAZHg8E7/QXF/piRLWt7ylKcFEddxGqVmfmA0zD0FEmkNZNY
7ofzZ7Ng8EbAw7otXvaPCsymqTXDJq2TduZfi5OVA2/m9GqNMsmBwRqrIpFxTJOG
NBPnjSQBLpRdTAuur/FLc3IriOsExwpjR07WMaYr/CU7B9VAhZTTuRU65rxY0OHx
h0QXusyVBWgQlv0yGrDh5J4M/9M/e5VTrw5v6Z8qmNBX5RTxooquwB7mTO5RKJ5s
8oyuMLYqwtRIElmukPnHM8XFSvKyrEJzB4iQkoaXKpp6USfFT8bg6zVdGdF97vwp
eJznNLZmycbdY/Y8nCJW/vgdIaYZ03UdnUkgbldVMcSShw0rAq6t/eNjvdEKv9Dg
PdKtvC9nP2LKMsshVYKeOhyFfHdCsSccSZ7mBugpzVP0wPVFmn1ZZ4JO1OJStdaj
1Cll/rUTKKyyJuanMxcL1386MY8yGvDBK59yPVt1aCkjgAQvYdkZ4MeykRbABlkd
mEIxfCXUU4NiKzLG5KGPkHWEu8Q/055ZG3jRwu+RFuqm+Y3rAuJ7sIwXBez217Tm
2XP5UJmrwOxoifa8AyA5yJh6DXjbiR8PHK4s07SNVCvQ3gXtbNAreEaguoJjOqNo
biXiT5wvNbbLzbD3rdeM6AEkXe9t2cHxYu23Z1eHP+AXBY7rGFfPFFPjvK8KyGw6
vl2t2/mEHusLwlRHhmULnpd/EG0wbhgYssTyPWGuN1wjalnAdL32O7DMa+doltNo
UDR2k3pDqRn6SYcennsuF+OZftjgZqJTWkcNdPHkjFyDSDA+FTeZCuksKSNmDFEF
+b1UKh5zr/RQH1jEvYxH/vvBBkdx+BaniICNxRgZc3in7/1M8O+qD8DKt2Y8Rjm3
RnXh+wGdE6Cei5US/8aR7k+tk055JWgDbkRVUbYOOCRv7u0oW1OSRUXuN8O1bOqv
dDnz381fMU1jrpscDwRy1w+72J5aaqOWuVbXZhDAQ9MHJfjNGZEPJp1S0TT2Kl4C
6Moa9oPfc55hqj91rQ/hTwizL/E56lRKiA9Aa1PKkQzUjQ77qf/NDbJGvhtDU9F9
0221nEcgrcKHTjfw35GZI9qpjikPvjeErJkhKFGa24WH2E89+aNMGDUSMTI3+G/V
WZlOSMlwlocegAIMqu0eotQ7dyMb8H6MajIZDtfk83aSPQzxJSxNt6KVCTsgvAod
XBjME6g5Wo8nXEylJjGpIReT+aaifl86OEkLjRam4lU7JsVvz6r1YvaN6oSgM2jh
4KAwXiQMJvQ0JMheqLgE/tg3uoLu85aHTRk9pnlgTxzwomceUSzlkq8azHho0QgX
lYszGhUsDETQVxrsTAQh42XfMXPZMa9AhavIrbyDaFKQw5uJQuBf/tnKHPbtXfNT
S6LWAuc6jsPEYCFZnMI5jF5OVUMEEyQpnLGPRSCVzsDmbXzMyWMDQUL2ZSG+diEG
98fSAKX/JNc1H/SWAZhMgvM5rTUBPEXEfCu++A51K25yIopoZ4KXVuRnX8BdW6ZI
rl9VMXmWTJKFAHrzkEEltjlGB9v2VNayVwCAC5q2WLmOfJJ5PmN9B4u2Ouhur9O8
08KCH4q3fxeSJMNO0l/NDqgdPMa9EWMiCIlNIXDygoNjMub6vgbsM2A0YDOXvLbP
6h+poFCoPFSqODjiyqwfK8jw1s+4PFaTX6HsK2Xx/ZXDzPG8nzrnpc+4jUnMOw97
J+nCJb4jNRNBtWUOhyNhlJnC0Fepqn1ziY5LjB2HgUzeNcbIcVNUiaimi41TkoqK
mWl8bJe6FY7AnqEodniCa33Khg63NE9cl2vhbQoSLlePQkbH9VqpkbiJerYepmeb
NUFN7m2NnAJwrX6yHlNx2m38tQ3Z8WsbAPyetkzurNzN/9rkZP6oppjdTgGbzigF
OHStuaEmSt0MjUOh7Wr+fW8FYDDS+wftT1I+X3Uf3mJ+1tKgamLPxUtszvpewAM3
39umx3k31VOcdHE9xCCSiS4MVnxDFniZnXWgEYhpDtNXGm1U6ifEhMgfkjgQMed4
CJhsLitfAcDuW6ASDY5RDA9YShdRsGJYubf9yk928RM7ZX2tdpqVzJhctboBUY60
67pVL7St2kSutk5mZ5tNTFbSOjjoHJvfe05htdWy7ccLV/OqZZ68JpIswzeCX9/0
deJ6jggnlVHpzuCKR7GvDNQXEoKajkk1NIojAby1twWdxk5+y4cs9euJXkzlMiV0
4+mHBeZR2R3b0mZnphcHR8gPgxPv+btuTJGzY9aDQx+o3XUKaqZ33PKQ0dj4Y5F9
4eJHKJH8U5CLmgL9wmJ7q5p3q72OcfBAA/yZ/AzNR4yajzgRpw1CqM0yHMpLv+/C
Uhz/PfDQzAjDTZpdV497X7hMY/DCR6rp1ZNt6Wn+JtXMXbYWllRAeBsxgZZ0DgUj
JQp+MYvIdOyLnUvp12X9Oqg+Mu1mP4C5jScCCxknsxyj4ncgl+Hn+ZduIfdFblK7
ZzKcCSQ/xvGB8vJW6gqgCAL92JOWgNL3NYEYXXtZIMOMAlTDiABDZpgRNkx6Jv3i
iaYNPBrJ1O2WEwf9QryPYXqqnlEDeXb8/HzAyV4uzPZTcXfzb2Yw65+aj7EY++k9
5P/zi4WrQPQanLthMSFhgHG8OP+yT67N85UDG6GJCmZ+lGTcNX9eM/pgV/ULBTW7
zOCeRy2u0X0tAn61vpholsi5wyP61N+J7xKyolyox9auhj7NwH/K1tylDBQm9AMr
fUKKskrJT7fbM4VSJBf5lOcPPCE+N3LK865U4Hrhwe8Vm1VjoiqeSFmxqjrfH0mZ
K66/3SW/fiF+gQslsm9aPHhPtRjywQA95npLhQSUN6yHKCEt5os3FR0DGEm8iOKG
RWOyKt88X9a56Gpxe3yQs8j4yTYkVZh1+vKtkDnOXPvo2IVgc5FwVztI0CVs2Mxe
Si6D4mt90pGTzhcfaJsVC228Cf+1YT2FGe5Dkb90/g18oD+GPCOeCCddgB/brRgc
zcbSEVpAKuW8cO/C89MmxTkL9TE8yBZnfRrXdodi/Srd0ToWvmVK87wgIS7SLHgW
8QIgZlsOqGqJ2OlHrbHxbCm0XI2TRM5mtt0frXYKd8Nupy98G+8KmmtQAf4JWb3I
UrZR0u6gzCZfiOLQcTCXYhTqJ3daguECphziHmSHcWW41cL8OBiRwD+C9qah5vNN
ZWlSolOAta4vkGLDag7LJMGHyfS5rOD4NbRrzfNH83A+jUo2NiQxW5ukCCaZA9ER
eHnAlKpJHX1uxzJwfUGH/awUlD3vNX4RRzVGmo4hChVV9bIF4GSciHjcBhslVV3k
9D1NOenvOwBlyqanyNDkbMdqvyBYjS9eRZ5lHjx5mo5qptzrn3G+Vhy6J6Cpg9YE
khYUFeGDA+VnGvZoNKxgolLwcl4bGTTVsclRhFzeBjN7kClPVyWF/O4+jr7ZB+yJ
JCAYv+OermvO5OKFni8AP/2h1ugsyHxZdynQ3yhUk7RhEbXlFp9f5qwoHVW/mFBm
TNfbmHkB18hl09QLaOT8GtV1xn3QwBrAJK7WoLSKLt2py7f/xEhIA0azJIJ0A8P7
nrg46B+Ddr+wQJpNU2yYy872ggmLdzqkdk/UPpSfTFmo7Mzcds/xR85Vws/5qMsL
91SkoZD897aexOE2LSNVVpUS/DZzmOcS76rNkByjTpzlrO0ce+KAb/NjC0c1J3LA
hNuotOsgIs+7X+LALYIC2yltdn3CRvPeEzCHMP+s+aEttO320UR7rPWOR7rbeROj
f9EQJmw9E0bUW+nFZRKk0Qld4XaICxmyX2EhWGkXI/fam+pS8zisy2F0khqQcmSS
qcUv3gK/E6/P5aobtx0LGsT/2Psz7PDIX4AxapomfY3GuOaSo00ONQsLga5Oax8H
QBJoobq9Pa7YLe48sNv3LGStpiLpgyPvWGCY96E/E2aeu/lTg7QuyuzeqIRRpvIl
nvRbnUtVE0DehqsqE0kKpnddgiga3KWwhrgNZ4FN5QtwUanUB1Anva6GzH6c7wZJ
hkcsaWAurOvkZV1dG9iupAXnCIlFB3WibdUsiZjdUTCOkltJqXv2diWXBMXE3Lgg
fWQl9vM1jcZ5BfweO2uSkYK1uSryUwwU3PAuAiXbEwXuN8pjWeyU907czBdkXYaH
PMCm+w89tnmE9Chu+WvTVBZYePOpfsEJBvepneB2d3fy007F2KxC7oRXZfo8js0h
l4AacVj/nO1YI40n4RhanROBQqWOxkTdrzFJ7A36HwAd8dUmRmEEOBXKK+bZiPbJ
7RpWjBvtc2ZiabygWI0uLujdvpGQSVW+vcNbY3jZZqRYclWr0QmYXP6j6wdev3ij
nAK7yTW17BUGX22BC47a1Qw2n9gkAvh6KqgkDRqxfBx7wyEmByZQ01V2UFdDbZ+P
nEqJzV/Txi77cpZGAckEBJe4nY5D7WzW+2agMxertCrp/bH69S92IwIEB3qM41dI
ALbwIheCwGrYsRywxBLe+C0RX8FNJiQvjEOhznGbzQEDgalmJUQBgPrTzfaR3q/4
e2qR/9pt4S58PDADjxj2ZRpHFPBzCpF9iYgjAER2f79I8Lc/+jWAxOj8JHG+jXL7
viq+ZyBo7/KBsphGwqj1A+pvhNOMysHYA/YwzDHi/Tb55Y3/WKVhBMVlKNC9r2Jm
NthjNB61anHmh5jR6vW50rmEIkkg5rpcJRSD6mJ9qHoNb6+QgRSHCs+7H5wBkHOY
95x42dqus7f/YgJ86++hMc0Mld5hbfLfuB0WjsBeUg+TvMAYFzWn5BGTnXUGZgJ1
q/eCSgoHE/dRKqmw7Y331BUFr2vupJFSRDbIyarUXWBcAaooRAoWJUEbd9iYaMD/
pEdY+V755KQch99CtmanBLL9Jd+UFHgR4JB7Ru90b/U6MyvfI5eG1ULLuQt3ofiV
2HrOI2DiaAaYlCRmIyIRhKBoj7JoDRwOQc8Un12D86V7VJnfeVL80jLjlTSEN/c9
eSbXYFRyBmnsofVjDhxoovfGT51zuqQBGa0JLCE6T0lAhxcOfl625KZ/k+fTAyNJ
ce+f6kyHUKB7o1bJPPtFPmilJdh5jvDMvkVw6e3LrWZL4me09s7ZL5rTwhtTzpTk
69MuLRONyFE7vqS/6RDXM0zyGWq7skJwoXykVtzvlPaP3op7TYKnT5dHKMjg8EBr
5eV1vvK73EPTbMGwoS2D9I3qqO36EOB/ZPNvabRIHwNmaSL2m23h59s94JH46qsA
qBIbD/6LRqGdgiSLK13FKUujtuWOTxur9piuFsuXzc40cVllBeN66Ro8UhQ3hzpG
q41eaC8/9aFljyig+ZFpcDllU6WitgXgzfDNeX6ihxFtRmnWJJHE7//hFqLSA0Fh
8nxR53sPPNZMFzT5FgROht2AqbdfZ8RmgTIekRgUTC2Ki8CrfFlNqLMLz5vimzfj
zKVH1KyloO3/UmQMCVpISSGjxCBBEB3e6VlFnF13YiXwBTa77QSoX8c12jLOQvv+
XRhTEaHIN4OglLvLeHu9zqhejqQqmciTy2MUjK2CGeQBQDUbu4M+eNtx7j67GK7W
hFRek+PIBvW0S7VVXO8L6szzHSacg0FKiLE6yRqpJwQGTfEL7gwCDIyFW+BrZaQs
rklKBwuuNkOTe3+0hfg2vMJlPjxxGDzbDMRlcetQhsjLVqdQB5v5IGznzwWflazC
/iZHAThzKOU+b4Dz81nxAtx2CI4t1i2jOd1PaU3YlXQZZKYmaHO2/Ibaxr5csKQV
N4KjhYX1f2ZAoksJo8FXvUaaKFe2PlfQXRngSbnavXRe4NP39QhTYqOUfvfkIvtd
P6c+FZIFHT31hOkshEoTfUDPlukYBoTTVfUWOaAWmy3SxqrAk3c3urkJvmUQkUUQ
KP4JBYJuGnWfsOqk8IPS9gxJb2BQ/1LFgDomfrqEdParaEHxu4L4C9M8Qfbp2D/o
O0dLHnRoJz14gK+fCELLovHG/fViRU81Z5ZTQULS1OjDbi3KBI5og+ClfVAfNDP9
sCvLSFaIn/T4aDouYybxCuj7I6BM3pn6lo3XOFiNOBa2zEqtI7R3/6Rli73GiwG8
TT6j7LgCdBQHq+NozdoujdWQZaw6WydvP/UVFe54zqHgI4aDJA6vS4uBu05PGDeH
GTlvReUOHaPK2qP6zdEEXLiQd+hOBrsTsbCIv+ctXdMB24sD5u5oOWsYPLjJXaTo
703ugQWTDd+j93ny2SkJ/MKeYTrrv2iHFv2UXo96HSQqxe/elqLg0on01OJS5ewF
DkI40buUcd3LbE9a+GNNVoP7NlOTA922QLyChaY6TpvUWnB42A8dUFH1nX+mrAA4
Qqol0vL07WfCtM+STzJUs9taju/97ZpaMbj1AztBiHnukvwVVg60SVhxgAajvxWd
Qd3aMctdiGn9WbSHxvtWIKrDq1I9T661VmEnZvugEedVroiJ4FBhWZ5Iu2aPrNKs
qSXfjD0c8SRJoC4wcUkAdpiZKXButoDOlK6pZwya8b0OQFhMON0bOgjzRbL58f7A
CFGKZT4c6E0g8gc+dm3a1DJIeYBxNN4NkiyKlGP8MqqiWL9WIBNb2MBf3IqbLe5v
bRAGhvcHvYAnurLedCzd65zumAIn5C1NMpldqwMJtwfnWoJgIYWD23mEXemMbscu
o8FfON00xEq7miaRLSiVN0u/zDY7OIQJaE/c8UtORBdtllvPLCN2Gn4/Lv4/70Gu
FyCfZX8eDl5aOUXla3KdkcohDbA58xunvwndbcfMCAebdm2RMQQBPYSeTMWy3jZN
4AZVshiZ6+rNsv8nCjS4oxOXU4pU1OJOfqBpeZZaAmS3gT3VmU85dBENTPqqyMAV
yzfJu0TM7PIEIDabhgomRnKsr6jwLyVmthfVyS0VjL2S0RAMHM/9EYvPR6hKxIwf
evXBCn6KxwJAO1S89FLpCmNp7x+BlAsqX1JNrH32853ikLbVmEl+905pYVPg0jh4
pDrSs+Mkbin2VUMXnySkViJMYw+SGrbgXIAaVygbCAbr/bZxu2dDpiQfE3PNv8GQ
nn0ihIo16D67rTMnHuJG42cb8q7mBQZspWQc+qO+rB3yamywJ9yzrtt1TTo2EC8A
gcI19ckZWAZROZbESZ5kYgPBt+BE3TKZMwgs0BvxKJM9e/35RpRESYWa0WTeyEhz
mFawar2fqYD5ERaTn2x+w7tiSU3pCt+Km7nHle3P6/e/OYIdijz3W4MPaOfiqCRF
ybS3B5K1F/PC5oKAOBSK7jeqV/xInx+0gfcX5eq3g6V8GtHSqHDttqNxdmycpIm5
3ir0JddUcuXxEeDNJUKHzkJL08xpcLdzUlWU2DuS1SyTTjbryrYy26ecHMJCEKAI
FYVNbGHp+hB6rd0+2K1P4Tqj0quJgSJzwK31QD0u0MLsyPvAiDyke4QHxDtECTX9
4WJxxV4PZf4iwR6yRm/d/ljKxz2NwPU9BSXr+NgIygreMALJj3Panc1+4Ok/TGXP
SUD8nlOgEkF6xiVG72Hfc4Lb7O0RU0uYPKQzwvTPy9AahJR3Ja7caoJzmpt/i5p8
4VA2HIhdWPBy8IgG0LUuC8kqVln7Q2GSep5u0yU76eScCKqXQpJANi0XuQnU9XR0
KDR5D6zm0TxKXfk8/SMR197VrFex/HB5G3SunWwESTQzwCmm10FK1+gbtt/i4l4v
8ZzH2YLXR/bthYta0M8OzX5QLB1zR3gNBfA5YlTOcRlJRw9uIggMCU8cWA2WUZ+s
yC8Fn03qsv5ukSDYGR9tB6A1wYw2JVAAFSnlNLQvbgCpOxZho0oKdMtqLIzxotSn
iK1S2GQH0+PWQ7r9hkQhq+XHsAPrcc3h6lskRugUMmw2SK2B4jnareL0hIM5N338
TViEyl5u1LQ4h0MjJQqC4kfNAJ2VYHJD74cupujZz/eYRDnfVnFaBUnLy/JWmoAk
iJ9PJ6/fZNHtHs4dGahPDeziSxdz4v6zMsmsuocngPzcAn7Iq35x4O0oFzAtPAxF
Cbb/RmrvLZCx7j1H8RcSJzo9dZ9X9gXWw+VyFT0pQYMswiw/XruL6fgUedZ50qxD
rQFKe5zsxrLyih7Q7MM6hudAxlxsDIyW7m1pf1iIT5FQnRxRhJd4KNBkVNxnRxqj
sMnmv+y8zROINfEYWCGtQ4FfXyv62wU7eFRsD1VOH04WobBvzVhXtmnkYXYC962x
xjEejBhObSPl1tbgRM4g8YXJJcavs6K7hht23q57GZ4iUcmwiz1H0+5hnePfCOkS
fMYaRenZYRQaQvaDHRD0OmUJS7f3bcqcoe2/kkfbESH9avDk3QWEiKaaRqZWSu1y
kjlLbh0poWFMfhT1szCXx4HqZjx1gWsehgC8pU53BmH+ONv807C6BuVGPxyYO8RM
gzChatDqH4lpg3qLVveyuvMxrnZNIPbO65SZyZDMGfzKeVZ8jn78Lanz2ZqgYYL+
x3X4bljcm/YuAr4Mz4B8aDTlGGub6HpX668gZ6EFRAX4Cy+CwugtAMY/JqWZrJHz
GRNx0aqXNvIW2WRNersr2gU/HoEgW2TLTV3fXlJd4Axi96VrCDr3l0I9Aa79HtsE
YUysUkdgiv1CML3nvmy1BTpXfSQLeHF0OpTHm6s6S/jVz1th8Lpvxq0x8HgQXRTt
hAkXLR0cOaPmYUAS7zllS0hVU3mVB7KeQMwW4YSngV3IZyTMm4r4aW8Vttrvv7Rh
uYomDjQR/qlfwSG7bPJcLHEaE3ZsG/XS4GNhZwkYn3fnTxn3Vn+4Tmp2MIF8LbAF
vGz/AWrdiQ0kn0dUjj+8MwdnJEEB5ScKkdo8uFEHpE+q34Y+vCsekkMmkgirtaP9
KbZ8Iu/gVffrrzrPQbap7c0s3HxiX2IREEq9B4iRlcVQSrLL/UZgaGB54Y9b3Db1
3khIiRjMlNlCSWFGBXJwCDlEdtJCqzH7ZQOl5dtJGgSgPyYC0Si4tZpamXW70vzD
JgvGp3fz96hzzsTL6UkSL9lPBv0lYi8quW3ku7tzzVkhs5e6KVu8WV2qyOjeGR3i
H8HzKStzI1RGXpJJc/aVpsrZsvT5xCWqc63mmHMtZeyujndcZYa+pynDjM5NWyaL
NG+N/ylJ/WkAOp+VKXbgC/f+f86CO3V3QId+hkUjoMImk/VVqvrkJkOv8j2EiSJu
vnaEER5T8GjkPiRWWqAWbJSU6e2Fb6zqt0U2ZGiw+z6mIgsqolM8WEHHuQ/m++FV
8P2EZLUmqAGHHjpg8tLTOYPZMKM7Uatmr2Oz1SPKjbCZBkt7rQZFJgA8OeXCrHS+
HZkpARnp577VtTfnBymVXa5BvWowPMB7CTM1VZL97edWWL/RsYzQG6JQUQJH2aQ2
+pLyccA0QF7kTDLiOovrRkFAXsqdo9vKJnBhjT12RfPkiNJzbmwgCt+SUIAg5eYX
851Ez2aj5dWbtK+yAso7qbTODUAZ3o7KYrB8wiPoqKcK8UVxL9t9lK918HDZAX79
OAY9s5K86sZD2EOseQxzd5qEI5yZ+kMjQs4wnudrKPSGd9SYZbRmQnz1BMuRPw4p
8i4y83GA7gV2jkCSpbv8bgGRiUgT2IKIBXVXPI8dbfCpiN1N6GQ80SKpJ7POLmHQ
T+trriMJKeVv+98IS5YcFuTNkrDndNXWoqbogFSew0+F6ay+eqcOU2LOvI8Jzy+l
SiUKxJtLUcVkH+oltoGKt1oeh+ksgN5UYfMgFjWTK5HkCkBrYHHz1L3eXVQbLq0d
zrAGPNl/KCmBU072IJXpVyXYiAg7DN+M23KlXbYjiw8gDj0MK4haaykFVlPSSWl8
or1pciLNTpqarjDgsTYncQbWJYOuAro61gPadlnuesxhrlsS5n0SOwBuQztd00RY
rDdFKazV+C9flJcCIctmGJZBJvX27WgSarKNcpga74mC230tBP1QY5wb+Oyb0mFH
Xt3jrj5zMwS9X0ePgspxU7HMTNW6/Bdx3zimrO5qm4y7ZEF2IVKR8fLEkrlnVNuu
vv86INa6W1d0WCPoE7rnk0wDt8BcKsAnxifn8Gq/BQHZY1DgtUgQCXqgfR9U5qh6
+qfxyVVpDbzbihFpXUspmZ6HKDYXMHc9SghAkO9MNXA0TbJ+mLUtaKMhnPiDtscS
KfepIuYKKjyDR7yfVksfDgUjrwaW7wgFHGf2VLDpv5CFH1uHhL9jAMWeb7DZmRY5
rLj1sKIu52OcM08jmoQX3xc+L0mfS3OgAFu/nEpLKjWbOLWcA16+5aZj7lfAh50a
1/4xJktR/UkuTtLmSvD8Pk8ICVwENb3ZYSpR66OQghsG5zs/oIgrntPITJ/e0WyT
WnilVclvEfpmnz15xTSEqQIc6E+XsLbCOUnUP73OWmzLZgui+Cwe6xgmavmN7XzA
SDaRd5wc6Hzb9PEqAgpGWqZJEQJGWHOGfRDXhGtrGvIDuXyPqIgtHxAS9wL9ANwZ
7jV/5ioQe8mZEZHhhZGNktPwDpxub9ZKOaYBXH2KF1wGPsNNsBOgRyCLraPQ23IQ
YsiqhvWN87zqsdR55Ft2N+8AO/B5sCGReQZ5J6+UcR1liQvc8GIMssLiege+Sk1g
CEJgBHqOhGTqXoohhpdU81752kh96Kg+kGv5rJryjriQwPC7wIjfry/3udUwg8Xj
dVGZSb++Y+0YnZ94pGcUmZN0p1hbAqwbYAeWx3G5MyC1E/TccNukwgNUQuTaz3tD
i/DbbN/lEbl+bD8a+NzM5jlPLWFn3HHnWMtDwG+K3C62BQpDijMNgkZq5KVj6Yec
VVSBYn0TAEFeCMtj4uocoqUR3A7KsIr7+LK9shOe7VS3xH9R7kpOLZXDVnExDF5i
yfi9M+I2foaKv4+TWF3XShgtvzHYNF/wSr3/j9qtwN8Nbroty9Pd1I94p7ig7jvw
woXwDuqh+IKnBg6T2/5nDkrJ6XYqWcDT4FMOGfTaHjI9g1Xvh9lzgXYSkoUPO8+B
i8JX6R63Hf30QagevPrR6cEi1LdvHBzJsngt89eGKWAcwxZt4YDVoxFh7JFvU2nE
H4RYbktsV8ca1MJgfKOvzziU7h2hxfpvmNhchZXSgioifRjLRMQ/FaNkS68HqCco
jDVOvISZXENvWsUTlCUQCyto9UeGZGmpsDVaobT++wQ555OeiNi/ouf4EHO342Ls
Zrh/j4yPmckXr7klrgo2j73vokVjYTxeRObz8tGkLKLDw/OGMrA4SVXUZzPof0+F
Y0KqojUvVDtaRITejBXR7lpzHwDigmfX/o5MUZvrkcriygP9hMVzqhjGoqcz+frO
tx+tj1IDa5r2e4hAjVChZp+Volc3vOWwrENJiITWSK2iWxsoKzzH7T1i/733vDA2
jUFHlFAx0uJNEFbvglGPfXuT0SZrRkkVnDJaLAqkNoPUU6M/A8e5s+H7GMk3yFxg
0hB1joBYc/wm2WveLVeUEnNhkSQztTqGARnP6LEijIY1r/wAoxXlEHynPyIi1T57
V/vbDjp0stnHRA+3YsrBLHYGZWGM9eFmLPR+J3/eO2Zy06NDnJfQYR6DlaKdCx7M
+kULUSSrDDYy1a+a3pfJmfwkoaOtS2URGZNaZHP15QbTnsk/C6We3wnNOqAvkkTp
YdJTvpXOrV1F7g0wiFc3Bp8OpR7PFoHooLz6aZrvuIktiW5H1SHWpeF9PcN7LSyG
xYSi+2zwV273Ufqw1ed2l5VF0cK0PUOoZ3R0iiE5YbEVRITmW5VLG8tJWNZmAx+P
I/seurix23Y4UOEfbVQUcTsMOdkKPSLn4ydXGgLFloAJYe+65I1kbW7XwVvjxcRC
3M5A4+pkzVRDJQ3mcENfv7fGWnODqO2hOO9vH6o75FRaaG0mnc3JABGUen3WoELQ
mEhwubdg/s3C4ujcEBaHDTBGrSbnbcw8Curp+eSd/ttsPAcr4Fk5g/ZmXChFwOgV
5dq5syU44pBLyxNL19kfnBB+W+1qvvg/GxrMbaF2plWmjFkIG9uj+71uNH4zFru8
yGXKo/cYGFEBiTk7fznfdTPwchfi4+IJkiCDYgVXSbC0m70b63anLxCNPFOI2YFM
7+vQ2Z7u35aMVfynvyxstehZ7bwtbm1GgV6w2r72JAB1KrMEeOAt4Nh94t+o4Cq7
RjDldJDs9k4ucvKLYo6GNdY0xUy/n+EzDCj+pWJefwbJFZ1deBLGpyUEssQVBgdH
s+sfSnCiQ2nXnuO0KD92YhRGDIhpqQ5LPrrQXP487CaEFs+Kcdp3SsbrzwDIml2S
+kwxP89yUwosteq5nqmB/z02oin/NCtxQ0hobeUlClzKUGgNMzJ4yXLgSCyIWZnU
Iiz72gG1ASGDZjaTagq5xFPj/cqXwEoZh1uMDlDPeiVl18soTxwkK8tHHEGYhhDk
in+5T9NkGnZtW5UxxEr4Wr8G+SZwHFtsinWv2/U0DQeCls2z+fsriiAAJtPFLnMS
8RGIchmCZJqqgrQpWCiRjt5cenV8Da6MkXZN6EEhRezeEoo9urQX1TCzzI5JIMtE
ggz6VJG8akr3M7WI1llztBDd8erVItpw06ONkyeaZYyNJiJuQkOdRswUfW7zHjCo
djjMRX01vNyOa4Y6aSImHm8H+2xQmweZp1IJ9y5o0RpDU+/v76EBXtWB7jMm9Tz+
zaR+1NM4elpD6N+Lwg0w1IhkrgXVLvQKjW216MBWdwLhW8InFafjrWExY6qZ1hPF
aFh6llVgeP3M4Fn/U5ClBwpcMKchIB4h2ZHXtvnehH5+XQHdWjJM6RR1h7LN1mTV
K/iedMhGSK1NL1+iFCl18pV/BjrxMWPMtICMKG55tCCs7pYHKodq4JpAkT9K7J8u
x+WV6R9JXbLAsbWJgSZ+o/D8g6IGSwBukF1npAzuN9a639n0bNMBJk1j/oDbF37z
s9LWPxRbwPX+U9CiWNDZFb1v0nuW2Ajv2AuINFWjIxbf6kiV3aBVJDcbbuFPPi2g
Wa5O7A+toWSjlPwgRnl0WKKwLaySX9XQJgNCsc0gHgXjKChh6BCWMO4fEK9KF8kT
7iK5IJE1cCsoHheBNdnQlCQjv9u6LfGK7xQFvNCEddxoUww4GSBgfstSX+UG6hiq
7CE9O1onsxmrKGMWKOwsC+HrtR6yx5Hoq3l1dvuD/2bHVQ4TZ6vHueeyjyGXo/AJ
HB3oQ+Q0S8vJAEFYYxUElqsyOPkd8yX5l3amDjUgUzgwb0k1WObFXGJ0+TuTP9gh
B2HcYZ1mcY0PzscdHmI6w1oB6kFT6JlaEsd1Pr2ESjVmjJJC1kbHNfCyy5aCuWCB
QKgfVl5QNGDwKyVmH14GpT6cS6+N4ZRgAUbhAqK3aYW2CMkQBsbhTr3Xb/ACKJ7M
eeL/eLE211Hy15O8mqy2PoIC3KH5QU+PpcUz5e88wXVIE5MaaHgSSW44NEJ+jiyq
kKaFfvl9gUyHGtpMrn6vnsFTKmKlRSYHWwd256wLHmNJ1Gffsov6H225F9q0frR+
QUkAXxqvYxY68vxheBzS14aVtxRONffUPoczmmJQ67aJEXnARtgPr1FkDg28CNvb
P7MTP95bc8olxmgH8EtxmLHhj2cd8bN/R+aaPQG1Em2QH3qY18PQiU9J6sHJqFiq
bEdavhmsYADFOtFRYnrDszF3qCnIwGl49RIPhl03UAr/JYKNR+xgLoIdRzd+JPKo
kZMbo9Sazx+8r2kJZ+UoPhWgKbEcngyjR6EpCHqomMc1FiXgqZRtj6KuYoDFIrQO
yYmodtcJfeeZ3FWdpjgF1NrBhx9RVNXMxhPOK/1cgHZXU/u6MthZTTVgmjcgP4/D
BNXsOaeTxRYr4a8ScZov7MVf+cgkPAcTfKcz/L9SoLPlYctNNjmTYuz1U/XeNJYW
W4Pln1fAO8eaiqbu4yRnH4c57wY3sC0tPr/Y6e58A77M/O8tmW9NYBvGbb+9x7O6
BOCAIq3AFkkCNUZXkVQjQ+mrQGeIy9TXy2VgF1ZuuObWCwNoXdQnNcuLjS/wXfmo
jnYLA+5+NVLZII6MgQ38c7cbRjRMpnchVErl7Rlb0twHqL56/ZviCKb6ZPpH1rGl
1AF3MfKhVvtimuyPsgcdhnBDtgEZ+1+2GvuVex8jpmpv0n0PSjxSAK1Sq8R+4QMA
QXxAaumld/MNS7SZwKH8GGL0JnQncT7H63dayz4gA3yQA6iUvtlKFjq3+DS2+eO/
DdGZvDRhr7q/hTX1sUO2zhCjQa6v4RB3md+69fqKsFz/mwP6RGxyBfLoH4Ti7Y4w
MExJwKm6ZBljOoWPeEBZbJKtEYFltFksjAABngsj00icFFlfnCcGEjryxADV+2Pp
UdJh13YNKiCcY5bKP4RxMtvCXudVtXJIKEctV/yigvLGWNeu5LeVI90wiOj1ah/V
T9Q4YKc3vCQjuFJ4SHiC5cATNRJND771v5I66gsIlnKRL7fgS6S1rQwZQfVp2Zd0
J/JK7a5SgnIOElZENyvErzxrDkznrrPeNJhon8940HgK4cgbYY+vML5Rf/eFgYEX
28KITsah/eyPTaq72sy15py4pwq9kSAydGWXC7F/x6OJjCDEA+QTHAuCyKiLFV1t
qtDBjvJmu8YtXmeihMaDl22MxVNK06gXwQU1TjI75UGMsEBgYhkBaWwTFXAGVEkE
oejNbwUs/ijX+sd7SEGVGe0t/hLa41qQAwAJuwDWXdMveJyseAdk/sy/2MCn/JJp
2KX0iCE3Ux8lYkwODdB9JRiBcf8RQgCjbezyZbsuZyM9fflp22ABlLT3bAw89b2O
FqXi3pY4b+3dG8iw32EZg/fxjUJ9m7T8SCqH5ljOra2YI9DHxK/cxoNFP8czdL0P
5OXlwQXxUDRS1MvFhFO9lV3Kt4yn4u7X1zCir/XhmZ7ed2nyLn524Z6OFXG/6Knv
JbZvlSkFK0BBRnTB4z4OzuXG2RpZHEUHoemTLL4eDgRtleV01wteq/u5w9oJjR7j
vwv91FW5C8vCkp1tr/Dg566pAxkfaZTnIFrCo5Qi4VU0QRD+NvKS5UyrB5n+bFji
MYwHnuCvjk2+3nE5K/ZjOPCxUV1eKptSI1B0tj+7wbAm5Vp24DeVzZcrl2MK0IDH
4res0/HH8nZyWx7YOK+lmyROEgg6G0Xit8hW61QkZAcDo/rFJxQoR4qfBNo6uiMK
5aub+6ODCYg7T/HH0vYBKUu4K/qPuvoqqafePs01HnIBDTCYN1CKshj/MEEK0Bed
9kkMZY43hjyutGB2VUfuI+J9Wf7ELSURHm7izJQDRuooJoQUI6ek6FypulloQvZk
TLG2CsYOsOuT2POnFBM7gCaBFo0P0zS0spzbKjSHnGazFbIYJrZFDvI6SUPRGbEg
qtCv1komTXajqb8rMQLlZXNcdZy2cfgva41CkRIFv74LcigXId3ASHwb3+7Or2LH
d78gPOu+KY38ByRlObCL2U1pE5LaWxtr3Sq6yK25TcVOdyUA1vAn3UBjf3K9ZdqC
rP0eXEgDaQZSKK1kYIeiTcSa+iEcZ5VQW4vGfoVvtARXqk5eyhFNVFtY4w+Lvj+B
fn/I5WRva19/pP7XtrTL9Ei2Iw/t0Git4cYnP4vUz5IUzxH+kBpHG94skYzGyToF
BEfKl4yx6mA3DaZvb4pqTouYUtsY99yGN4YmiuzT9m1LFEOWGEoP1NRPPYbbtubc
+RZBtd3csodtzI664DxsnLjAUF3iuKyC9DUYQDppUSOD1wqly4BpPvi1BamPYby4
A7FtQ9WpkmpLOdrOwpb6Ux93A9CKTIlaxcRJ2Be/Je66YfgvNUkOeHSowqL9TKbS
cVtR/6Ux6cEp47aJRkPILVRP9vXwIRkHE/6r+Qt+hHkz4Z0jdgpef+8y9OSZImea
uvS9jOUKI4MyV4dVYp53nm7cvS9J320JQ81dV76UGsm735BLkhwKNffAx2QMvsW7
I3NVsz4HK/m2ftwhqI+aYaiTkmhXyDgb/4gAdD1GDiv98j9NDjfuGKkDCdfUw1J3
r7ifZYw2BNSRy62GcHNp8/PmVdRoJoGnG02LWXg5Tp4779dKKRLZjZa00o68W5tq
FnHUSDuC71NBngT2V0Lm5Pz1WUBvK4Hmh0YcaKGa1pO90+aRR5PucA5+vzOIPI5H
jngf9rUh0LTwgy+CJeb2H/JUEVU01hcH5REF1mV91G7UkBZ/P3vhMdsg5aDIPvgP
rCV+Js+jx6u+PT3S9ft0euDkI+Aiu3RaSwEqOT+FzvMtA90TDVjDUTWGIICVuoz3
VQ3TQRbHr1cTwVVVUiKz3zNLxAuY6buYzZ2ZvCs9Tv2Z9jeDsux0x03zZsmSs1+M
MflD2sLHSIVIRyS5834SOxaqFCoI/yHgUVaHF7Lvbjx1fbLYLPrXV4CSCkGu4ERt
XbdcyUHtnop1Y0hDmYOuhSRp9+2dp0jf42GU0ln+k8WAuuCiiciTdfMFW0NjvnfU
r8CTRyYcaxfeAn8NJbbP8xwKlLsfujE+QWsPRDeXtpnX6jNCu7HBCOBazgUMOLD2
EMkkBCE3GcuMq5Lyy5IVENIlIJuYXtEn1gPYG4QI3+YJMiEg4oHTJtSEqt3fuZuC
NZ/Ti5hH8jFVkljn5o0Eh84YUZxZqpbckvUaNj1s4UTDTztksd+sCTZfLCCU3a3m
hKAfIs44RywX68SV4LxZe1biiKGUAkQ3P1z26AfSvDS6sfvkQi8luSaRGIDK2WV+
8RNPwVIrpcqx++Uk0T/8LHk+Jjt68SIgDQf/86YnW3iK2mplyQpTyf7EqIVvT/td
NgkvrPr/2d/D3T+jCTViOuVqwPDYT53X6qSsGuPpwhNuMTMkrLA83eMG8tilH/Ls
IkaIXx8RHd4Gb1KoQlvUSApBx2NlJZ7QMi9l2KmRZ+YBLU6G+EPe+ZwZxEuFgcL9
qXGRmAMrPDitSX/eQoedHZ+5OVPK42tLjhifiNNO40bDTKkKx/DHmUplM2FkhGjj
r7oT4J8GxoFTKeOA/Et6Ntf0GR4n+lENeeyjSiEiStfCLieKmBqVjDFY+7wb3eFn
h8zEY6eUmOyMq60+m9UVpXsb94vvhPp9odqJRQx+tBtU3GjLloCMIkp4JqLmtO2o
8wxnLQbbCiN6d+DyoB+4Co8/J1ouv5aHah2u3REjovBx/Ze2ERxuHlvtaQNd4Z3a
VVNKmedNtqX65S4jL9WPIxtjwXuZk7K0hy2N5xEWPVP9e5Zq8r52rUfxEDTJy/3u
LrFd3EYzHG/R5+onFbkLTQ1uDZddYYtS1RrowUFzh7wQ1AFcBLFfSvotNegmjwPv
V95zwd1futjlf6Us33qx5f6aDM1YsXXQXQNoFO/ANkiiiX03STqfxN1pRxhQ4GOQ
t9Gx3Ld41SDjBeJVCakqA8M1rbdCKhbBrg+3KbMPblhaT3DolL1v1TL4jdqgIv5W
bKKiNekTASpdsIDkIPw4NmzdjMSxoAseug0I78BTQIdTvMJMxW5zGEqoE3UerDd7
OEhfvdJMSg78v2AKfTv4UB7JkPxIcG0YRvrpA6texVp7DSxRLsVn7ccwIA/YMvf7
/J+P6RdHk3lASHUyQt1PqkC9YGdVrjPAiQo+RaMHXiZYbAsov6baxcH9L0m1lQGt
7+h6VKiY+rxbOn0PYiiWfRm1TqidwPJG+H70O1A61e42Q7E0pKGOO8WDJj7S4lIh
Zn4DAL5ow9NMLr82+wz7J2l6m/OtP2DDvtqUL0TovZhL+i2TUsHunZpN71gi0YLK
8CS62wS8+an2ZZ3yD6SEdihkAVyVogPWG0ZeuIoVRvfKHcLTUVOz14IuQ6jpy612
vXpxz1m/W8EGddT0jDzdYSO/uPWUE/EIU5gZ97AR917p/GLmeJsGpgiK/yrH6aPj
w3EiKscPmSkO4tI/tgzlwE2ad3GSiUvEaib+cexVjvSvRLhZr7Zj88JQXQXOFi84
/krnEDmYr7j+4CGmHef5XNRGkc8tmsJ3sIDnT8fKyfDhoabnLyla3dXCPT6168mo
Pdt75Y6aL/yASoOjTwGipEbeGYazoC2qMRFv0E/y4Bk6c8d9F7tlH8Zrv9dKR9rT
wlKth66VMBsNDlGVM0qBnK9gycJ4r5uWlXOv/wdL4tOH+dkBig9ooj5h+6zZ+4Ff
vvx65KbCAEWSfnSu5H1R/K4/4xeWXB9DK/Gav5MI9WdKGCJtJpK7pqTtr4cTN7HM
ywFMDC80SaPFsTpGal4p90HuXtwBd8FhoID5j7zSM2yVWZfsayHUoKiRj/+N+xf4
XE1uo7uH2iHv/fMU1ubrMKKwvFVZpAMYrD8wwU8uwHlCjM9jB+Jb1itMSES0uteV
rjwpuexUnLXWbENx7YPyp1j82t0MCO1YEtmTB+mPZOoMyxbyCDndiZRe6Xk0NZKz
ehTqgXRcRjaEIZsk97hz3XoVjiYOAE4scLQREoPpHiWtt9sFabhPyA0FrsUv6uDz
pJ5YTGxOUn/QLY5eBk9ujHIAriFzL9qwRoxJ8qgxVY5Zp+yxVCHDZfxJ4mo5MnVC
yYGL+4QQ7CAyIrgqhMoL3D7SyLSDYFPo5Oq8YKemiJaarMBfI4zKnIQWSo1TICH/
JarMiT1Sgz0Ajs3IAqYfGoecT8mooaQiCBYZChQuuDJczF6H8aYgJ7ccYP7TpSNV
p1S4VhqIKCc/1pqqbbgQu7nyavpfx/kA7LlXPUbrsNcqVvPv7cue/6LkwZF+Ob1l
FbOG/yhR6/AA/wQKCaCk+LaE/Jtnx1BcrwY9TTy0HoXq4bI2z/KbrSQdf8qgPP+Q
eS0dblKQcHHORTBCPylKTpDYp5vD2hlFF8t1DhyhFojmxr7uZKQty7E6cBtRNG2B
6sBBu7o+PxwJTcfsHtHdUHoWcsysyA8ZVnF0khKFarO3ou9hcqlSQKLlA2pPi7J/
Ugzs1N/0/YNi/wx+r69acm0c9UVylpNaabqTVpLb0FZAK5j7eCadDCemYh2sLTUA
OMi+cQ5wEJDL4xmqmaFBnfspsYihyyOjQyXhOo1wBxkfx+BFY/oti34nCmYV+zlv
etemFkNh+t2hVyhJ9BhRYo7y2zZGgLTa8a5W6TkJ8jHwat9W7BU4prQnuc+j34WN
RO5uZQiZFUFSzy8lqrhvqORHlCxXkTN5okLz+c7oreE2wUu9PIZb2qEVtUFNjVK6
lo4JmwDsgCnJ2dpO24PE2KKZUt5ilj+pOcGPTYQeCjhJWX5VS+DWrSrH/gjebLg6
wzEsgQBfTs+ofy71SSXFdP+FmZXW84j3YXvIm/sqSbrYwMnTX141tAjAAgvzU2z4
foIyqpMmUHraHLD4b0BOauNwrNc+agJThvPFhUFCo1LGbUmwiAJRWPHQWQKLdwlU
PBGSsY2G9v5uk1me6bvcaSRNG/P9rTQgmFR+JBfLKSus3pOzPZdBF6E0B64jyMiA
lqf49kNJ/D1aOwKrUDmF9BurprAoQpRgI4SeGLtHKs5N9ShkiGpAG6/PdOI43LgL
AR1KeMXko/T9n9Mrem/h8Nyik2+AfDcAlY/sLWmMbO4vDoSfyypMeKPePhuNClEU
Dv8QUY70dUdK28D37Iumt6mM0CbaqtLmmMuP1xP3wQSApf/PZOgGC2iBxuyxXpz6
d9Sojr3fC9m2PW0LaoKUQ+swbMKEVLOnJ/BzVQCP58BkxJBm0ehzK4AW27hxcc2j
UWAX/53e3VQ3DycwNb7H7g3R/afJ4D8n4gjSSmApicCKfQLRAqLni0qtGMBNLZVL
r5Y4/syuMPAV3AFNSH+284ijKW7kEhKKvvBBcyzq9zJut4O6jfhT9mC1MC1giSta
I91ystbEUa41v4Pp8yXQgyVv3U1yAs37upgJcVwNhJ5Cg0fnLIBJoivxMxFUghAn
likTJh/2wzLL3TUamv5axuqDd8tqZQOQnJ3a4zcv3oA5pUxPFuOQ7WdMUtyJlTgH
HK5IQb/OpEo48EI844UOU6qzj2TlkQNxHTvEkZNQVT6OdD9T9YbZvMwkxJAfloFu
xlvUJRBMLtw28meMcp87GjNuonNYfbFUu0JeUk6FoXx56rmrcfnxyuJHpIoObsiw
mowpdCkefCGaCHfk6nAPuqDBgEZMFGzKFDXT8C3MyEVdKBNLhg2yaei2Mc6dP4Sh
qJJVSn3t3/xzY4rt80/TGJhG2y7MhkBaKgJ5o7MoUmrGOMv35luTCSUtMha4LPrZ
xEQ/mG+w6KX3BrEOC3O5izDjojgSzS/Q/0yqpT/EsduSQq0JV+VKbufn+QzgFkt1
4HSHyxqUj8WOSReLjVlfpGEJRPz7C15hVEnZQbPQc1GAa7XUm6srn+PUYIBUQBHC
NRGhec7GlCrF0+VOLoNgSS5l6y7j/k9dDqvlCPfu6mE/XW0gy8yWu2Jcq2Qz5nuL
4OMERUEEfQqfXqQQBOv8q2PrO2qUhmrwP04cY1pRj4FM37uMcNVU8jnmnfpt3dLZ
GyyM4twssvQYia4yAs1XqGooXTVtKEthYrXL1RWwmqktz3d6UenICqTyMWtKVZFo
uGg06d64TGq+l/H5J0XhkPzndYCvxcVyEuV6+xQnuDYmb867dfqTSTEpyVzzulIb
ScngTx++mBH3Cws9USZNKn14esIxFvQZ0JZqrRSB0gnujYpHIMwtkdcgK1fkzjmd
ZnJ+Ut1TIQVWl9jqd67fi7S5y4E+6S2wetJQ2plcQMNVGEU9ySXB2rrV+eMq136R
MenRn5eLrLaCi/xQMo7rFMRalpgvebSFgxHbLnB8InwebuTB16Gtd+uVysIg0hte
2tH8fb6jHATvRpBpgoz3TWm9V6BiQbzJ+2iITN/JldhYV31AHoReHsoNl26q/VXT
NBARAecJ7x6lnWVJeBuTBYUajbe1K5BqL5T+qgPXYBSpOJzF5yxDqgQOC+NOttBv
MYhIpuSsRbe9XIWe4rLmgx53UEXi9bqiyvRjpr+BLCe6Kp5qRxOqTOrEx597sbGj
QSpDWZdAXWpJML7pK89LGSIlb6O1/TB7egC+ftVfkHQjbJLg9O4Dpu8p1DQnB+AV
8WX2CF9PQCrN23FA/81dh0KppSXg9q8w5HE+Xp634oV2lnrWIlbKr7xYjr1lz/Lh
92qoiKUGtB//QMB8PPvVB7kV7VJuYnT4GCTw40mm2P/pKE+A6V2irLc7K0UgOsIw
4hJDrVAvymkDperB1MO+ph3DKeUbillabjfX3AWT66hWQ7BCcPuCNiAVN7O95HLz
PgNuQAtnam7YNDXiw0jOCT9iNB57Q3BDLSNG+bxmv4/C2Siu/o1nYaUJOl34DbT2
YSvBFHNLj5e/DGzu4Kc+pMzjeVJd8TFICRiUPDhN2Hp+QTFNtNWZX7NeTAUAsgPT
RnKbjvGbwNRHVCF01/5BwsGSo+yatx84R8Z7LmBUGsBE31lU1R+437pXzfNLmKuI
ElYQKbHOcbDW923HW7xn0xupH/UKeBN/aByWOdeC+EgsoigrPgY4mVzypmlt7OJx
B2QylaFDgGlkQAH+fPjyl6xlkAcBHZQK2HPAfxJMpajLR5ckOwlTCt4QxPdosgIA
WPcXVPzM4E/4ifHEJQgVEYwIY+XNCPMMMsiDM8rLnm60/JEs2R2KJnFD9lmzbdlT
Yri5S4yUQXPdRNHlTYHVowtZpP1koCQae269g5ivkXwviZsXeTH6eMR6j95EJV/i
w7ltTgasO0+tGVb+YZauU95OqEfz/xNbnJO2T1obMU0IJ/aVgrX1PvBkuVMZRCYx
D7CkoPryvHJY45hV43SX+IkhKRVSOSWs2mYRz5Fff04eiWzjqSBO2xe7V4bjBq3m
u1/epYMEdlGOglABxrmfU76a6zpg4NNrUTvLURclAKEdgHZ3EBtuXhMZXm7ZFxAR
E3S9CS/qbESyVBYNuCgIMhEezAdYlV0+TWH2KwW+UIV7Xj2hNb9SdPOQmV6jGQHR
s3Y/Ho4opcHuJWNGZ2XHCsIYwbh+ZeJI/5dwJDLMVqPTyPAQ7WNgtAbnuFrSal6w
H+KVqg16eDn8d2Hk6jTKTvomjQ75v3NCPnKktX22nOq+9T4B/dG5OZD1oYQ1JQMl
5LkbuWhhEkWESQmSJTQYmKUfL6hrH1u1HAZuf5GBYR/51eQA38w7mjvfBHWy6XrK
fB/uG/kN6EUFcuoB3K9vnz8qkXTdjVyaRnXOPcLEBALNfy0o16oG0jKhkiDnG8b1
ZbabTs8g9BuiP8AABEtrAKW3u2O5FFeN41UtYgOBM6+xybM7EO39xFlAc9orP23G
k+da4oaGmZJDEG8GchI6gKhj9n/XOkvsXBpXv3GoQ1d7RefPnl6eHQXIjTUMpCLT
azmx8ynDS8obgLr9u26ExP52jL2e03q3R5PXw7xu6YHZknrXpvIGq9SV+yATdhs5
B73dgljBKrHtFoWy1s5RI2+6RvqMEQry0LfjjihyChshGVoVzKuO8vsaGOMS46DU
QleJRV0701c2hvR2crYGzXMWGZhS6C3/l5AjK8eJySh1QlJlKpHZQ0VFtwnDEmhX
nrktgXZAMuEBNHnU2NtrzfNr4EMxfAxvV3tIBtSTMKLcB1BX8aVq7/QyS4zyj6Xj
mI6gbaxXregWp5seXjGqvM8bz2InpbGerHKKtUvjzHxYwG8vI/6VUd7dwRKKipKu
v5ouK3p2Wn0GUB+rJo9cdNELTRkfzj5bvGVABuLCs5+zHrYFsVMOFuU5YJJwpRCi
KOkpVrKQzqw/3QtL0PDce8eqJ8YGRFEGKg2ihX5slJtybWKO3kLbSqB7SvBpy7QO
IxO3lqQpU00MgaFvWclthAliEX3YubSViONlX2wBvQ9IGdTsW22dIMhBZf8CDLAj
GF1CfI4ttGvvSE7EWNo9GgYzhmK1X2Wh9yxqL8HvmQ24jpY33fSvfJU0vtdlC96E
QKp20KedbsMP0W1qNPm9Gj2hxemfGptFGTKDlIyUc48GYUcTFk3sJt9aeFOKkaWs
1wfsxA8bShcpE17c6csWzSKnk/sHXHPyFBVCsG4dZpa3Cv/7lk5pLV/cPHBSmsif
vdkeiEFiN7r2aW5Lu++T7rxdTNaDAPvVpbCmx1YfSPsMS3qV1tWYQNqTDc9Mles5
5iTxUoHAVKxwgFp+LCNBkJFYTncAbqm3TdiQtTGL0UqqGrLFMgzo6QJqs2LL/YFt
8JKF4RlkO2h6Rs1U1mmKL922m1XemBmunRGRQ2LNpjwspGcu4VKQIYavGGY3L/n8
oNpHg0xDCC6/dut2s1vfU8RsfNDiSUuXizFJyzXHSjlaX7nTrTF79pHB1FgaSXz9
5JPqIcJ79XtId2QvxMSyE46kCBvbmtJ3lK3irp8IzMaKcnQ9oYgJtwb6hF6RfFW5
dwpyEYqvaZW8J43wJpBj1+CGe7cMpvx6TEesXgKA93fTMe7e23r9kPeowlNlwWkc
4Oo+RnyI7p9bkJj7SGSQbqTewAJOK7A1eNZadQMa/rH0DPlyoiwiMIe3xM9cJoY6
h/2sD0I5NHfWzCWsE//GCJy9VeV8MienZ3Eh6oOjTZJLXa+uMBtHUm+t13vgRegL
XTBlUFDCdPcSxQNchVuSyLOOCAPp8u1qAs++AITn6reC/8jLCJzMA5KRVWarLJxM
5Izm15LNAZWjyRhkDpsU5KSWRSdGxkAi/jhNHSYWD7VADr1mkiuOuPWyHqwn46By
lqfgmUJFhNWO3QeHhNrnjEL8MXuKLoJucFgCW/BJgBdrAqnYXcvyIAyssQCZFAwX
y+tFlwo+mpJPgAusNhAA6EWLLiEvr+7OtQpbb4JM/ADa3e+xcbXXY+aGoqrfBM/9
4IItQXNyN+ZQZLUlmnFA1K0syiTa+ugPPMoT4BFFq9Rs58Ar+8zkXHSIYnbD7jCN
8Bgqt8VeSOGPUziJCVVEdxWQQfvtth3WkZUqPtHli392Wf0pCqX0yZltUcWgNRnf
3uX4kDOKuT5pOkmPy3uQ90KJMfUkxHNyRlZhtZTraK8KSMERkO65dxJV32gZHfmM
kke/Ob28e7Suz1O3sJV5FrQg1/l0zHEItZ+yXcU6t0LV5Pb9SSMv+VbVv9nwPXwZ
Kmuc5L2ekhMGYEmLaWZlbbJ4rhCKHjRsbw6gFLFdDeVoCuNu5n0YzIXGxNqjykmQ
GC9gLoCDkY/RqSzSh2xPMB3d2Foc6c4vsqKjeb/7JH+TRG/Gd6D4e706t8Y51Nvu
Mh6+O7tlqj2WCvq44oZDG/yFUnDvuB5AXxi+vXkhigmCqtzgD8ISPsGQw5/2yaf6
J0omx0UeaGD8Tvda1y7328CtYAnCHPaI47ycwy7oieWG0tmX9hqqJhj4JAm0nOYz
0ervCQCttkwfHOODybyOKNmRYwdMkQE9C6BPhd2jbQIxQE2GvYezZt1ZJwKmS3cL
+7m/7TbmD3hV8r0gB1O3DQ+Vcf59ByO+necSSJa0m426O6wbk/qXAzPqnkHiyB/P
RPo7cHdJmaqsUjH7ZI/iBV2Hi/fFUiaaT5eofcOl/D0IVCQGpEREwhYdfmHyXGwB
b0Lial5BqdaUFDJ9IjKCqopHU5sr3dIysu2SE1Q1OAeEOWddAcUzWNk/AgklBsxv
mx03H7FWqWbF0D5hLb6cJord0pfU1W508KYm0iQueRXtkakwhJPVWnFBK/D2VMLr
+AD/0PMLWr9HyNz1wLiO70JN9FvUW94Xoj+Ixidl38YGeO1x3iEAi7y41yMrf1iy
sTf82jZo6XmEnrh1vTsJC8qD3k7KKjn2K/sG8AQcMYb1AoLZUGuhsirS/FblhH8F
v8on4u7QgRHEkixpx4tEo9JBDH/55IVpCi9/I/RZHPHOO1le7P/S7ALGPG/Mwg5n
zj35ESITRHehiCFIP1dgCS+6OA2/sm/CdfmGM+b7IBCWcZsDKLzSnVKWCyu0gW6l
c6pXafVoIZIfg6lO+G0Tee6PQQzVB/lOxVYaFqJPNCgfy5mYQuC4GWFf/orNjPHL
dmv8J+CgF/AY7ovII65H3mNRHtBr6xnI5O37hNrTdHUQSCl8CTCCJ20w+72qMuJX
HmtFF7BdANmSM8MR5P80UacOJThQngAVAb+t5YT1I1tpo18HQe9nQLvxQPG8VI84
L0jW6u+IENClBg/QLdps0JQasJzDwEqLuoYTyai+/arCbMA9VK7ub3AqiHvgG5bK
oozuA+7oYfgOpjVBp3nzS6LOKVeb8MMeHUDIbczF9yNP4ce8QZfmySLaHouCzkIf
f2hxIZ+3vD/7m9SrUV/Uv56tAGFw2z62TX9fyRzx7BukC+pxXiGdD6IdvUIDJiuR
QiLmUq4GD/EPKKBrs5Dz4aMWG3XnKwrhssIel7Ruvo+Ms+A1dPVo5Dwdsr9QKhEe
sfNEMs0GqbyZ7PHZa/Dsfq0W+6adEqmnyqyY+e43qXiIQVjAxEqzrAFQ4cytqlXg
Dbu8f77g0OqQIlBe1LnOjPF4GnoKwVTEZ3reZK3hHmQjF7V09WL+PxU1n5HkYDbt
rcYj4eYw4NZGdWVLP2UycrJDk8xQOtVUglfJfGStQU6S3RM8815kP84Pke7U0jwV
hyC/gq1s0DEw8jzmojBneaqaHNtK7BNivw5Q7ru1wR5W3oAQSDC4p581oJBbJCSz
hwC/wgrbWDHDooUXUFGS9H0w+fUe5E6lKNNqfmeIM8N6DviABaEh/7ct8BI6LUQ7
AJALYd/fP2aOIALt1EyLPuKZcbLgHKNAcT8rmsCAVXwzq+aiYeibcV2+fhwEMteY
2m0WXxr6ui8sxmOkyJ36/U0qqnR6PbOJQoKGVd2OlmRT0WHVoUv6vz5fwbkoWA/C
DfHbcuNMAJFRyyBLdLgI58qKy53JyLzkA//OGtz3WoqbcSfqIGTSF6UsmIen8X2l
6kXTdpyn3wp8bSxr2V588P4pEHexxvjdOTikjj3D8ucHRY52Mc0qAzRj01xtiUJj
HipgkIwiY3F4bCYy+3jU1W/AY/T0ZnT+caPIviEU4eUudiNlEhSxctTEjuQM9sKk
jAUcuxhqUSxxdVQRg2jbNP5awvePMgLz1YIN/BKtpGRxvz5QwsRm5alGPYZJ6F+4
yTa0iMLZ9n+phoApcNG4773gZawE9JLXqS9A/9GfHXNqG1AzKlpRdjk60+upR4lT
ZlTnYOvvbhNND8zzjU/dRFuP2EVV8YzKf0zIckAge1uH+I5GoWdVx52QuXShdnqc
EaNALWKnlo4EqQOWt/nfMRTOm3/kPdxZEnqgp6n+7JerMTaYeLtUCj4nUqpJnZPN
/rDKdfKFubTc5bknMkxxvYfwFdY/VKDjNC5NKlob1FNkJdXJVvj/8jhnvcsGA9of
xKjmbj1sFwK+qX2cyMddYhZjYn8pGFkKPHgZ8TTiD2jNGG/M7drFksMTIBpm1qgd
VA/fYSH7I8l+x7NXFqno3qzWgbYL2vP9i3V5yLm7ii/2yKO3UAhlEueKIkqombmC
s1w6fbKznPsvGe+PBcVx+Y9oOIVLJML1rM1sFF/7qcx6f620fDKJUeNuVUz78Img
70cwCWrU2YWatPqaftIakqDMREOvADcOrNvExhHOds7L5JJCuDy4cwsMM4UhMXZQ
WLeRv7vt4Eq0uajvMzHRnI0XpxvNO4xKZdD5WU7DNgSazZe2QyAyQRaNzFQsGP0q
cuFdd34SvGDKrgMWmyqYtg/elrvCWif7YSXzi402dDxtt6hP+lywKRDj7JKgS9AU
CeuIHcA2Z7bJbQAGMpfOJ6+ITpDnPz8ZjlamfouZgl6Lyj7n68R2g96aTu1t4KVh
4gdJiVc/lgQWBOQc3FHdgWpzXaEFjlSHJKGEd2RegGzvUmSLYqjKYC+6Rb5ZYcMZ
qwvJDevAZCJ0EEziyxzfacL/agKlzkMQast2naujuwJ8Z1VoMkWwTFYIIHE4EX1z
+jrwwtiIBkY+O9czUEDV1xrmeBPqJFVps3xT/CIHmwIy4XCD3k6lq2kbZn4pc7NF
8zV49Zl7rt5k+TXj26xN6R3UBUizdmarWz6JW7Gg9aB9fnfALRgIjqVOPjJsp3qm
bFOsqgzkODndUqvBt53LmhDVIYO28CAD1Tbosb/AfKc4lEAXpUX6nz07V7tWqLqD
gbZ4q7sJweB8PyLCngyvDAIubZmyCjSklCwVGKO8ClHmgB7/QJmE1Uoac8q6qach
lO0xuLyHEwTU29RsQYYUWO1l+++a+vMzoSu1/k+8O5dRfdcY8TyzzqHyhsJJIDFM
OMgNMebWem4OWJ/GcZCkaLON5J00Y9y9XF0U6tFPtSk0ugX84rhCtyRwywJANeQy
gJ5bRFXYCE+Tfn9VzwGTwdjKSR7V4gtJ0tRafMqFfTQzKOYiLZuuzybUxdfHCdYW
CL48+NgQGqITWYCBEn7bKLr3tNsq+Zo8we4NXu4AGZG4Mj4Szr6/iClNmSd5gql5
p7MZTgpj9/em4pXJBKFvfApvE0QQJKzIcU6DVQDvxMco7X0T26PIiNtzGUP7hvFL
63a+HLOOzb1iWHuVlauSOf862dpNd4DNV9CR+/6oPGfTsNND2XP4D/biIsKOB5QD
K5+atnAeZs86z79fnlZ5aPbV7r8y1UaKUSSvh8YR3HELYWgxSVSg6bO2XqKoDAJq
xaFS72RGFUI00PsCFFNOWtbePSzuhEhGGCdGFFO1Oxd3OzgNSBJxTntx0YN6kNx5
kVQ0DkQOEGv6Fo2CEv/+CuEv898AxjyobQ3Rw9c/A895IFOPYv3E/NudTEC8unbD
qzRB6UxGqNnQLzMuTdPG4SSUa80k2ryP2o1PRFO5TeUchFdnBevDsnXSg260hshd
0Wn0iNPuWM+xRm7WdeJ/i2ZVKVRLWBsM4aSXrLww/qveDk0TcFtt2NPjcSvsUyaA
n3S6K+JUDOO83KQ3BATZXYsmnKWrR0Xvx1NGaNcF35z9Lx/XNBlB2Fq2LfxY8w1/
4O5r0um0dveFc3tsGOVSO7bgK5MVLjYxvkiGtPf9QApq4rCHaSbN2u2lakLfF3oX
4zFm3ft527I8jNzreQLZPEOAwQmDg7QEzVms6ic2bl8bu0oHcAvJ1+dMqK1r+3HF
JzzX7gs5i8ISO4dxHZUudhgzpyG4OYKTrYTMuE7+fUcjBEjgH+CnzbDyIhtCSSSi
qVV+MTwF+56bgPFRTQPgRc7vFnb/3oIzaNw35+B79vivIo1HhMRPq7YS/Hazcm1Z
rM16fh8NN6IgbNRkyzi3sXf+dNsQ4pVwGuJBJc6r/hw0JdJrkon0Ood1alMw0ypQ
mtstJgGVmJBOqQ8nZ9GwMBByJ5xEYbRYMA+L9wrHLVpOQQ+omw38jfrRRvWIGWB1
0/2rTWMKBikbyUqxZltxhwAET2hg2YprxsJfjoqBWkVRd78rLnj8JZqc51Fs6l3p
U2Juc2+NomywabUOkes8TGeEsnkylAHBjI3NpjI+1IXdKk1NcsNiaPneHVfCbOrl
AZy2VYlqTZ1Xw/7HwPmYHnB9VLSEbq78zxz2KW/fslGQdo5dgovbk/M2avndAPFt
7Ntoe1xmiVRIb9YBhjTNaI2ZQuqt3+gNwNmkYOu4nGMAe5TS4XgVC02oXoGIyzt7
Ij3DoIup4oh58U2MSXaqTPlRhHcxMv0R0O80DT3fhPEj5TWh2Gp38J7Yn/XZPew5
PAczFQclEpthBI4bXziTCcDaFspipjAxoFfdSD+8MvPPcRGA65iILygK97krgNDz
tihk/07qnNbG71nivjjdDjI8oThdAocXYbeQQU/sTbOp0Yqb9FR5ND+qurXOqt8q
+vnPPMytEeeFS0vPyTJ1puA9Os3md+Lhs1WibotxbHteL+DRJJCYqnbh8Re38Zg1
3I8oW+iaLci1BUI5fROhzbNHxoDJarrsgtjuDECuPbCKG3IwkHevqkbjK/Mwgn9D
QzlLAIWBUtHSNIhNqroMUKE0pPe4XTjhJldqZvD2YTG7LqS6Prp39Y3Veq44K/f2
qDW3u3KT7Iyh0OH1wPhaO3MkQh7qlaiOv6oZhei2z2TE9XeFVvl0oOqhcpJwvX14
ywF/Z/pKQY9hLE2JXu95rbGEdPV0Ev/h5QmqEmJxU4toANDWrSh0YkCojVpcMcZ7
FMgM+5xJrsz4R17OIdFP0kgYp5QHuqkb8c1Bzv0irluHNFdKbs8MCPgrZqiSrb5v
0z2JiY5ujm1gTzZ034Xp/zn+w0z8yiPsuuIqVYvSkK7TLiVZEmc5EtEuGcrUSQGR
0jI6omAnJn5ODGY21BJ+CNs7MxJsfvlmiHoJw6D+B8sIZ+ZRqIP8TG67KoplOikX
8DLbyHoJRJoGf5aYABTJkR+rDy1DWG45EJE5VUblk8xhjyl4ocs2IoD5jSmxcPlD
9L2ienVsHQIJFv+tjZBiSD/JkGJS5T6dmHTpjOmUbzRULtMCO9uZTKIpM4VSvF3n
OyaiVBrRi+cadFV+HNgufE2RKd5J0wybkZxpgAI9Z97H46TdBwn0NEk+UKo5YH49
6eaI3IE3ggjWIQLn+Tt/pWZUk+h97LBjihlmQuKcKEz3xD4HAGGNzuPeK6BqOqy+
AFX5WoC3NZVdbm4U7G8cJuJv5oEqbXPAFHZdKRZVHFZvMTXigEhYTiNEdZK5SLi2
7w7mINaMKj89/gxa/TxSJuMKu4b5flvSu9hfeX8as0A7VqKqXHHLMbKjeYgFcKKQ
MQ5A5vVaFZWJiqhffAj4t/gIG5VC42HowgSTXrUV1KNs97HBImqGhUrAaZ6GZS64
+ykQ6K0op8dd5Myi9vy4BKiyCg7gHs2AbCWMM+p2VuTd8B7Z/+G3D/8xd9tCaMZj
zJ9pFiaC2L0BjbhF4U9fORLEaDudmSIzPO5xGoi42wmkYhtwMUCIZlm04L5G0jrh
bXR6b9DDPp/e22n6L5IOQLV1GDp5uqO5WqBAN8TX23bcZa3dkjXfmQAchLb9UsXh
k9sJd+md/MH6LdQqFnyDZflkpmCMPGRauVCEfZrHu3Cqjox3ru8VaPtxmuq7KBYf
DJy7u7r6u54b2/3X3epiAh99aK91Pkyy3lvxLz8yf7MXlnUJVaSh+mM5ex0tX+ck
4srDYefYXc9Wr9+2IOIZKPG6f9UObATgKT/w8u/SyGYbnBmmgdovGeajhLyat+KQ
ozNr69pLs3d2vRvDO3BDZMHACUr4liaBprMkYVbqJrmcRadSNPtPHIghk19wYzv7
a3BLtUSdEuAuGeDLWosuoHWlGqNDYLKWaGTiViYbVwwYH0JCPELhfyk4DJ9aTan2
9/65ejmXIERewCtmXo57qg2Zd/8ulTY/6ComHAxy1ZkaBDWl3/+2tfzN/3tzf267
SQEDNHqgcW+EuuevgzdBIXlmQ+5Q+GYAhk6ln/jYRg0PiEspVtr1GwUMaABhBm20
spBc9jgTagnhAPquYZfAZZSWuL6Jwlu7NlKBXCDcpbhXghRYcb7eiVVaSrx7sDCI
P1dIsDPmqqXvjRrc+xyjoAuBXsxEiKNVSMloGV+AGIsPJOvZB+FrPq5aUG8JzrNx
ygjSQjhe6yVvAqTP62drsU5K2R5WSuRaUj1vJS+N0QLEcBbePmMs7Rk5VqjBnKNb
k2ul7eMre99fQ3xa8zijhMOjRbsvHv3KKJ9AXcUnx8DNY2QcGYBlHMQKHHxWUhdf
lLnp/zrDR+gNUTyZqM2JhbHlrT0HEUtjnlMZgu/o/wuFA909LoutAxFnJbjbGvk2
zXKs4Q0+WKtV5WjYEcHLlZY1knfRhIPG6qojsms3drtfU0WMcUBRe+ft27JhMmQl
B23AI+cxboFM/lbUSQzlNNP+GYoGjCz5aha+S1kp0/8ciHOoq1sclbZB74dDskO/
yr/4a6LzkWf8sCzJn/si0ozPQ55q4Uo1n8l6Oy41PLKKAq35v0wxFPNkI59nwvRp
kNbGx0chl7UV+ljtbPCF4mQBxq133xp4ORXgmM6pJRd63jBIsoZPjvWRsod3Nyvd
4iMsJRplvRifzckvyZrmBZz6YImL3f+7ly/nqLuoO+7NsYVEnrkXetz/LinqYbkG
lkY5er4xlEw4nxu8mEno//187RByYISLaJCLAihtJ/qUMnRzdlgMAHc833Vk/Bxo
btCkNYK19zraajySkBtVtuTJ/KPogIXs3q0KfP+NVhqRmpqX4EenhbEx0saMVSBB
/zDdNkcmogZZhRrDOLvBj5vvPJlEnppSsMLAxDol6tKCfkSf9Q0ZHU1nw14IDBBA
kFOU0+c4VFgzn5V/N1NF43ovt9Y2S/M3xFsnSP/YjrLkxhOswr2F5EEo+z5d0/+c
Yo+cJgIKzw+qyH3unz3m16KlP76JnVbsZlsl4ykiAt2hpLbL8+5TNMAx9nNF+Ab8
zLx1Ige+ZsL+ZRGMbfp8R6tJDQkZP85L3R72gRIKuIK71r+Y+26bCpz4FwokqbeE
z0nYOxf6ArioQ2HRYiSuQpvIzsBMs8Y+StQP3LGyFTULXVECotlcT+FLihXpB4qH
yEBycEnNHEru5RC3fWRbVWuvj2VIcXEDwckxSkghF6DN0oUeBR8FDOQKzR2Qk1Mb
nzodCdv0bQfApdOS+tmH+NIQELBRwnjUo+CYw29uymuomxSO1qq10wWx2vTjlN59
ehnM7iNlIHVM/EgVW/6Ldd1kFv6N1/gP4r4fMUcnhK4ca6LQomVu6nc6V7oe9HN6
iHhPbHjucz0LUHHOS8V8IIvuybfdpTe7QXW+KP4iC97BQPmfHWz9L2YGTrQhyHI+
zVQGxmUntVaQsK2aKda5TjX+Q7uahzbk9/P0m1zHx6xnb9bTwPOpYIHoXnTrGRkC
PGV1auUkfZFAyQ+mQL8tqkxURPkyGOSjq3oyHuaSjKpmmoYdAe1P9CNQmxb5RAiW
0C0N5H2Uz1xWik/DxW25qFPtYWPcCE3aN7lPGV4Meu5UsEHTFGrRtO9qHQdTb9nY
j4paMMJoxcLnuU0YeFVhrp838Vs33wU+uv3+Hhtv8BI6yJVc9XW12Rgw4LxuKSo/
BcUVd2NUeDQh2SPu5eS0nrcP3b+Gq6TRtJ4ZNdfdHxiRqg1D2ikGoaTBw31T4Lw1
16e5y40oZ5FKS+48eM9PVP7pogLeMocNJ6b/KcYf8UldyrVw9eRLGdqxsDGi3N1M
O/wGlEyiLnlQaJuLvT/6WRYOVirHWC2jpgy1TJoiVq6kC8FrIlvqFhuhEsg/EsVc
vSBHqzGrVEtUAEbwxlgJgrJpWmHgavHvPOT5tVYysi/NfKIGWA0uwi6co6AvT+8P
hLHlukNxtUEVky/KgOOwuAp1x3/GPEXBi8uBuHB7x3QAdMP8z6ki5NQMxwHkMB4q
gA5kqmV/fw74P40XQnMTo9NYyCA35fKz4PlMCR9y9YN0xSM+/570df3irGh6Hqz0
X4ZZtUYEmquBtlvbYdxcBWaCfh/DJ4m7+ttfD8Om9iT1mRUb3cEY/q0Wk3BQhl+j
Gg2opZK4N+lorVawHpJXcGb6dqfwhMMD6fiScISkUbEyaQRlfnYeU1TRoJaJU4Of
yxv0b42rzYwbXcv01DO9CHPLLK4cqGx6CiVKFnBmsd5YjKPpe5FGhir+gsJt6akn
hazsr/Qo37qcdhNIQvN0kvXnOcfaQVQBujPo96nB5Zr3ju71rpoGPLD2/lxcC4vm
djIu2oOs1WUziUt0GqKrw/+5CmwO7zEBHWQaoG+mLqFP/R004RWoHxX0NW7iSI84
xCrwGkrrFeFC0NnwyLB/UaPUzLAhRVr4jFg5QRPJxUaDOnwwCH7KZMxLkFsTiqER
e8EmzzABn+xSJ575PGZ7Ka9Mu7WB5Sy65BN1g73ys7yHz7JtZPCfuKNnek8FlqCg
f1auTrQzEg83NlwrSLJz++jLwKOWG3C/Pob+nUCjDdpjfDW7csK0M2u5K9Wn7ZO3
TC1lAmdPHFg4S3b+SKhXqDxogIVrfD/QFjskXG8vYo+mJ7jH+fJWgP+mSMRHUcN5
Y16wbFhSBBOa7x6LdgLggpMrhyfmxXqlLKitoDjo5Co3CulG1Pkp8Czfqw7COWUy
Yyc8g68D4PHfsV7nPayNfNbEXMfKqz2P1y9ZbF/lfT2tM80jcZHCpJbVhKGbj3/a
jNjMACytYqBuKUK9CC1rIHgYjCToC4jAgI2yNvNhGZ7+TQJQQfcySlYCNHxwKOuo
vW6odbMHCJZhgTeWgVKe9/wAxcFu++WWzu2QNZqqzlRzrBfsm/pUh5zwowZJXvjq
DV8Y381+gHP1WRmwiTqCi8akZ+XGQW7+jhpEOndOyb4/ntX8UVKbyrUrQXyOxESG
KVl0In3jJREtK9nmnSYvWlHe9L5BXdwmJx8CafJtLBhFcnJOa758kY9O40ngkDiV
krFHBDFFi3G0xvx96SmOZq5TpZDVLnX2wHvEI0GFYzVqciyFDPhi9b7D0aDzIXd7
mMdE24pCv6taAaNkmBMl5ZXhziOtrIIw7DdbHAAJ7zLfEB7PyCNptwLNP/+la4ks
boSgpGi7jZR+CmPJxHb+jlMRKcica9l2Kg/eNIsH3J7AMf7FA6IDPfO2Z8P/axb4
c2apxauAzqKbvh47oG6owffvLZmJoS5jVtRnwfyvKqcOQrOgO9p/eQAPcDzUhSdK
cXZf9Zl8sNpTsqihp5n+NPrFQaCnNbKiNHt7nhEmZ4n4i958Grhte/2NUUcsvh0K
H1W7HPQzqoCg82i8jEX3zlJRUsSuF02iLGMbVZ7J4kWK2kCXvJToxrOqNzQ8ZB5M
JeHiPxrY+hAttJCoGgjJtsxEpJ79SW5AIhwSI+fCcuMRz1NCf8R/p9osY2HQb6NB
gJJw7FrknuOV7XENePqMTw3+nWtA5gByP5hjnQz0DNlbQIjrtMBr7ohOnVC6X9LH
TGXE/T7+FKpZY8QA/Xe8MfTXTnwnEoUEyf1kv1zI4605jDcmBALaAC9AOCyP5+s3
W3J44DVMQkzUhWQBqtaT+dWkbCf/LRKEcKh21p8cQU/rRUApBn9fCKT9l2gJ8N3R
0/IPi+hfLU1jT+MUVSwZgT+0IoqD/ZJ+uYZRBAYsjjiNky8mH5YR/S76f1KS3r/3
2nH4O9+oQj221Tm3tFqTDH8iZwE4IqnVr/bGlw3JssygfLmkHNvDpJvkqKi3GPmv
1LSJLFTMlxapFy4hz2BdPcRa4GbCMy10GM2DeoQ2RG2HQWi797r6PWrOh9BTWHuc
od64G7qzq5+QStD2OFQaKc7wXg9sdokfkEfmepuwr51Tnf/z515qbmxGY6J4HCtl
QxMISXpmNr3mzItfPLFw9Apik3wnzM1iD7XmbRp966hJQsNvRUkv6Fpjp5Gjdgin
FuPp7pSuOzLj4eKpyHFkhexD08VtmpAAdhAlpM9u3cF1IHfw0HgF0/TDE1jzldlG
/ku/ZscN/+66+JoXSoxDcvNxfq9bKqFbgIFQs9MXVKcQQbRATmKMhH4Qwcwq8H88
0giPklIfxvjele/wNDy5XpnE7QfJWruvsMpR6VDwyrYzL4WN0TZatqs5paJXD5G6
BmQJssLZj9T/ccWbHoXCxXQskDXRsn5DVLbFYaDMM2zKAcLsxwGWS9zIbgk7dyNG
/ILqSzBuBm81MTkfc6qVXKQxSKQbbsCP1JAL+HBi1IUfWyOewkn/hmgLp3919MyO
Ok/rP1sHqKcW55Bp1CJdU2OpWYp5fuv8D8fphVML63uwC8R89ro67ZpqFtMaOVuO
mXxOuwE+cr0UDUGBpsSIA+mK6pMy6enBj58fvraIrnOeQMjLbvjHuP6JFpRoeBFB
B+xjKfBDUDDWYy0UxkvBRIDLfRJiuct/CW3BHvNhHgobrXd1yiXlAzVjsd3rtmgw
t47hqKAVY1XNW3DGex49kFEocs7AgGzidF8sjLorutDou8Fb3+PyOHTir8KY2nD8
ID0lJ+Y/LpdER4u00UsE5y0l4slG/+w6GYS4B10D0cgEBHmRJDczgquKZmguavYt
afWC05JDvExr8mxqg3no6SQ5jVrEssdHVB0Vili4TLoMkubsmbuwE7c0dKuLcLF+
7OjoyahBDvFibRlf9SWV8y2PDqDk8ceAPzhzThOgmp8LF24ERduJzt1DvMm8vlRe
MwsyXu91e2egYvheESZCtqCQk+VTlRNhWg4rLhBPST9hrIpZiXXOiOLvc+NoJ65E
7avXmldAVoe+ZqNuN70KbzIZCHObscbNu6Hgwal5TxHwhMTSbx4wlMNbXw3gkn0h
2AwOUCkInzBWuMkJfb3DLLnz0V/vny1hi2bVua8N6yksgepcNqTV7mmSzegPPxcb
izhoI7wL15H/Xb12aFya2k6qglwCxdNb3xUSvXjQBANsMXhmLHNrrC2LMnnXw12b
00DePWKo9DNk1Eu7UDrqpNwkHzRLE5Z69ExKwwqcQ6HQhIHaTRBDB66OoA7GsOeB
wUlnbTC+rsQlaF9IfILaROaRfXQY9wi0aPvQByckjsdNj6Ac8SLdTn1V0/MXmeCb
hncrOxT9Lgafxl7CwUICSfRykQZNCZnzFA6A6RoXj8BH0gFF+HhZ6egVODt/scJX
5gaJEfP/HUzuGbdPmceiTLsxM3DjrJm5np+s6vLDERk48bw9pPtx4m73yD0WJ7+h
+ArfxjFiCg1E3g7w8Bp3CmvwY4yEySyrGilO3Nuz4lA3gHCuCmWkZn8dDbfpcgRB
EEpi/tJ020yYNgZpHzAg81KGVbEtTMBMRrRC0DRwcE6/0+F3UkDyv0wNHww1DtgZ
DgdSq1ovpHNm7FemMMQrrmP6lJKOv6Ci/D2B1n/PYlUO7umPsworqkqO8E60R3Kt
FFDxj/+A1AmQvPBToYY+idoOQANRFbTTZoVdsmSoThwNML+0QedUgnCkSbE3tTVm
eCoWS0x5+eoLFIGfVxu+klq3KBZys6Ri41AlCCR/J8ig85iEAeV7JnRuOn02Qi37
d9edRT3f6qbwYtSVQZl4Ne32TzZx3akj3hwU8oWCGljx0FgC+8jUVqSv2h9yr4dR
xfGooIqven4Hqk55YnnUsAS1llEMyxs8C4VL8AdlRYtDIk1PjMZa/KcUGda6IseH
/pBh5VN4GCBytFI0MHf7shdKKw7dPjmA23mhTEgFka8SafxoLj8zR+cq2e74Upjk
LAuiUxNtqN+pmS7YIWvorzMHRHfPceHj33P/EK+hMV1vEtO4cLWy2C681JBlQIdF
+QeJzM2ZqNkTJue2jzm2QomARXSE6yfIbW0PW376hEzO8OAgGqwT6/nXR+TULY9m
FVK0U561yDt/uNsLIvU+BaX/agaSbzy+j20v7hksAmB5pAWcvhL9Jhd0IRUQeMJ8
/965qbP0FGP9v16RzaUHFbuMtXh99XLFE4RvrueGK4yGb6UTGTGjeAIK/T2A+KwI
nyQFd8iDEMbbAUrLaglbFOvSq33nNtMqoltuMJMmi93hzM9w9Ge+b81shx+s0Zeg
7hbOAYZgWKz6SLh13u7tppZRjPBg669JoY89CSMn4y+mXM/tqtziI5IXirA5Bsqt
/sGzIxh6UXTGIvzPYrX8D0l6KD1i+Ajr2n0lXn5wbaETw5d2RU559He+wsrgowJ5
emS3j5qOSVuw/tF68uMUCbdwL0IFkVt8WpD55wzZDEzaEbL67hrICWSoQ6a5cabb
HlQxsRd1BNhgSZFM1bQFHIfOum9uzT0w9nl5Fo2pMfZJoiw/gvHcoswAOiyJqZSq
47lUAOTeSQGZkzWeuheqLDXoREa5X+o2LnO1zbsBHB9DmZfMx3P/4UjspOLqEz6e
DTIbQEKKafyfSHagXcxYadQcJKKWAg0dx2oY/rIaaW/t58kHthAUkYbwExHgdfEH
U6JZCSTj4HuahdIHxeD/tXO25pU+wQBqNXR8LK4cl6kNlyGtP+R9/q/I7aPqokP0
SMRo04HqhjP93w9AtdJsmsPhnlLKINey+C4s3x4r+42fKy2c6+HqDCAzXrNbzkD4
Wxf2AVgCotq9Gw1tlPqab6krvQpJ8Kmvsv2gcLYSbCJa7qqq89eI7H2xTBUXYlOI
hvaHTSNMF3ydwJ4Xg992nI3n1tw9ol6I1ne57aEpLGktNf+KkrooGZr1geK5KYRn
pddrQ8pSwoBZfzH8u0PJ1b8ZsOZV+V6KqPcidKij+0UBcso9kEXyXe7tewMCBymU
YjmHkqFBsBxnvBhCJ5PLWbSYoyVmgi2O5WbcsPY1XGiDOub5Q63l8QsJ1mPyTtBa
uMsOwnBKyIqsxG9fWfcbqfnIznJ5Cl7ciqTQZyfukhRxglDfTfe3sEqPDcaKNwlw
l75Q26OtezVs3hgnf0R4mIT6TOPakCX5tmKfZlOgqTb/FL9PF4Qnpt5Bi/0rIgmQ
b7LWFMmgiXcEFa4EtKydjItJDH948EmKGbnl9o6aWBC+JyynK5QDybzP0/++axQV
0fXlxelV6Lkr4kG5Z/ImXUiBMyXmUCF3MOGSIX0MaPB1PGDhKgbgyAYFcz/Y3XHz
OK33/B0Hfbt+D3/innAHBoDcXO2l7vfeW9FFwCPeBYkheyg1NbVARS6geNo3UDm+
6YXf2d6dEV2GD2OQyFkuRZL3E9C7bb1qU9RgCfvcoGZuG8Yl4BGPZ8KqiRKmXCyL
xxH4E8Nk0eFqMhR+c+I5wT0E8d8Q8ZzSL+DfsZuTmXcMzUSD1Lojhe3ZRIOlzSc3
o4y8Qqieb/7PwNtXVpmSkgbPB4/nhyrDkd1rI6kDgvQFcKMttQ7Vt8VMGCCkEStI
005HHKGJjOjL/nDL1h2ECAijmc9qfVKq55F658oGcN5UucdwzXnRLAtql1CnS623
ChYkwd38ouKje3+FiRqVXmZzQ0vnnz1m1S3QCEvQMVw6BCsyBGoR0fn1fwn0++Fp
iq/Le5tWsPnxcIogpKFcLGJr1ZY+0/eY6b7ZoZf1uN8lwx0k8ybkIEz+5JGKif7f
qa+o1HlFRNWFRuHMf/JDAIt9thcwnBG9I8ssAvOszRuZ1QOETLyFqg+wtQXrTuS/
iHuoFh0i4VkyKTKXPtj+829Q/8sBRn7jGY0lGnTEjAETqtx5+8oyEI0W+kp966SC
04l5inmeP4jUxBwE4UYVP5Ww5n8XTWQ9s50hA0JioBRbOgJ9o/+3HyNakxZjpB/u
AXVsU1OytRVupcH3tx0k8XFZAgeEpGdZkUFVoiuLAChPvdBUKQTizJVnkqzKhawY
rDdqDYGFnZywWIFRda+nERNmZ0ScH0x0u/aBfhxO1QlSbxMQLvhmoqGk9clv1HWB
La91CrDrTbpbBb+8j5NfjJmznC8vqHgLPnaa0BsDyTVHOCMEtM6yFucVGapzXtlG
PZxU9iVsMP+hMarHgvDJWe+Dge7kcsYylzUZDBNEKL7l5Ys4cqDy4cIGJrVpFlZO
BPRYR8jubEZsOjnND559Dz0CcRj0iDV8w3JPjgW87ynRNtrR9SfgxHcrRr5gFxpX
God1/niJzp3k6EHjl0SBuRqM0QsXWMIJX9sfAcpGbp1OwYvEF6faW2nVHFxkEpe5
k0RTTvsqnQW1MNFuLvPOr+Ve2Poz/uGs6CLtUKHv9Q2uiGR/UMjzTGglG9/Fv8ty
zCX5xKrcg67nY87DtQ/Gd7C8+M4P8qU0RhirCMfmyb+806r8eIbDKRM8iozH8b5J
uaqQLFfICDJY+D6OIDs3ayf9mISWkaLIQrmuGfolR73+SK5Z7OF0BawLEKlWXpQ3
3t3/ccShgj9GEvgKtSCEtW2nCHGp/wdTrn6wLhcUrN01pCjGg5xuVLC92qfUOUEP
NSgAfn29BWOKimaETASuV0Qqne7UXyJtsx1f/Tyzjard3go+yYeqOhNtRl5aBNCx
L4vc7YS+IYgL6Ye7tIgcg54qDWmiZv3dQuTHCzLwNVHOUy2B63d5uCXyrhgTMe/k
p/i/8gl0ypqgyl3s1KqYoJMaaNCbeimlB14CTajVjXwBA743Q3nBRh4lw30AZllE
YzvsC+A6Cg+W0UQgtB3Y6myQT0T9p3jCVfKAVWUtJ4T2xJAfZnromodCA71ov0M0
zcFtFFo/9eqxGO5i/JNlaUPHm2PhX5SBvFEdtBvNiPAGpFvmS4XIvblI7QpKrgyV
qW/l9kO8/c2krgoqpXcsqrTuanKLTvqGIQNjh3aAueHW8rtIAFDT/Tyl30BnW3a1
ubOik5hauHfC86imjPDDQGMkVCZoZ60qtqN4qOKmiM2D72GVeLq7p5x2qqrvNMNI
ks7QDHApyCSUThU3K4Vn1XkGWeNPlf4rgB3bv5c7LLahfzomRRpfrEnpt9OL8ah3
K86Zu+G9lMjAalt/iVejPX9JyCqVJsmo0twSq6th8dMrijPDBKVzRdSW5xObzKWl
yN//7qNjtjx3tZ60t786x+lesT2hpTcVaNQzwOXK0JQ4g0P40moSU4h8PvqmnBzS
JC7q29tZ9rZh14MzUTWqX2tETHUEi3bCbApqhl5iaaAqwjTxsP2wRZfrek6sPyEm
UDdDGzx0VRPbMSvXihQE2xarTAaIOnuNV96yNZpJt9k3wBAbEAQ7ssYfGfzsOgh6
yDUppQZcq0ZDx+tGF6mS7DIHsLAlRbqVO4+W0WFyLW3thNpwG8D2eC5TCade8aS3
IicqJanJN1kGui9VKaNssGHlj6d8DF3PaXAeGDjoceanS5Ayf6xLADh0h88yTv1u
xDxQkznZat0prFohRdFcuhZVKQvzyGOirXjE2cl83/b+lJZt8EhRbMcX/V2GBtl9
uN3A7KsZ1CZtfBNVRrZsORT01xOfesQNzplDEbiOw5Mpxp/Zq8hkjKoHulDg2zsl
rRxRQU5QIVoN5p1pilaWybigPoa3NlSsYYK10d+5hzrLIIlDcDbm/ecPzkGIQ4GZ
33iXN+5X/Vh8+ELQ+F+SbLGplt0p9NiAlDii4X9DHfLurrDzQQDMAYhF3DE9MTKQ
ObCj7ZyvxrtM80qlDwng22T6ODflwuXOigJuR1UrEbZOPo5DvS9mEuimDBrSUNwW
FP9Rpb+ENWTY0ieWMabX8LnPWKzYMDGTiZKIJm4Vrc2Q/eGjocMkQUDXxpwNQzYO
PK/nZTCzVC4BqW/P4IurAvgrBILmgvcLUIe8lFa7CPq6dfyAp3+3MaD19pay7Mub
H94Op/976fmvMAMqnyXiD/v/HhCR0aJs3DvW+Z8vVGc0ojkXqIUykZxxkQQFKHCs
141CEbryZBTeN8HQBBtW43V+Ah2cZm+VKeei0ud7Somnk4IOxTEl4kDcuL9wKseQ
Qhe/pITrKwJIjbSGYH8ebv4VjhH5E/jHeiwX0vqJ4JB74sgn3mVcCV+j+eMvterw
WNkuR1TsJ/trxta7fRELT2NcyP51Cy+8bpp5nLlqWi8jnbVvxNb9u/gRJBQ3T9C9
QQT1En+3nCuNlvoUB5tuP23d8sphmci6PW44RqP68ECc4/+oHnBmo7zrmdKrwp8g
4d7cz48/8RLlsfLVh7C1MPX5WVkL+bc6ymtZaBlhz7191q2hHpMMmFNJyIRXPuJw
tA3crLXN2onsd1TcGs/2VWt02Yunj7NK2E2yHf7EPEZX+66mvInZ5PuXodq6EfJG
qvbjwu0tPKDN0ODsVOQfFsKE9wBoybcHYwGICm0HFJ8bV13iFSxo7icdSGarGOsW
EN+RKyRQUlkLVtHKO9v0Uev0Xpndxw9OPskjzjHh3/05V18CxaClhlrzF7ZSm1CF
0acdp5pygv14MBKL7retk/OqyH3PBja34Um+hglNarQvQh85KX3oQLbrFUgBh4nm
tEQ994OlP6mqA1VMlje2tvYFf5ftpBdcbN5NVrZqrUgOWpEeh/fTEWbIo6w5RAIL
G98mr3PKSUJKDeJH/TYspUt2QD2NZmYs6aQNmRijj8sGNaEh973VCXxnz+jMTBB3
fmk9jaGdPD2v3p8e5SZ+92cKCoOQdO4Aet8C9ibOFDO+i49mXrwO0Fpb5WkKcOFG
9Ki5mN6aoogex6o6oI3S2avcU6tKwHVwwZ2WhOr210sZ0jiYcJk9bm2OTWUD0+VH
WvZdyloo1p5lCcXVNtumH524VAPyR4XP3Q5Mc2yyobLadZ55QnPXGBlOEwvryG7Z
reLWYrSk+ODp3zplkaeOUCYfbfy7xWMnIWJpWc2gFy7hISzKxkXr9aG8n3k8N78t
w+uRVAGr85vATwchn0vAuqt+FtmInxKUm0ilx8mFk8/wp0Exf0TGuMCkc7Ts9Jot
XEwvmBP2bDJ6hDmKkwxZXNrFQ+SWQC4Xb8FW+/RZ9ZoraSRM2A7c59+1B7uF1cUb
uoLrTKuvwtFmjoLNswqtMeQ33Sjq5pL/fKT3HsDyDCEVHwZR4wId6t7YbX+v/fiC
BbA35rHQJYG40oHB2gCMlQVR/2S0+oHibzz2RDPj0LzRCO/6sbwZPoFWZN59pO+y
5uZFHANvDBZ0FumwxoXxh/oxC3ik5TBCFMWj11XbB2hibb6Hn6u7FbkBwf2vfEeZ
dn+kFwxnKRIalwGY3FK+RUBVco+EZa4xRI2i3UoaBMm9A3Z/fL5JVvaKElwfiG90
R2wRsYN+7aurjxWfwI0VsBVI84X84breD+ntUIriHe+iaFqzbyAOF3xZUDx+xOgk
FqPqMgR/auDQC+hS+rUyn0oevPd6lMMqnEDP+bwh3NxU9MM5QFqGXurjw3d6xLsn
NkD6TxwvrszrAQ+gDXlHKMm/IqVmi6xn5zyyqdcxDp3SCyBnt/y1Vw9clGYBiGxn
Z8tAWWlTwbBnkfeF/kcMov2YdapbrEZqgD44tQwV+GW0WCD8MF1wEFzcuN1XQVEc
X/R+X15rtHZNa7lLfxvex85hegw7tWLikIjHt1ZjcAhpRa+K+P1LR/7JOqlacRix
/ytJZnVQ2H1ub4x+3wRDoertu84vA7X2cBgW6u+cAC34DMwJl8R7ZdNP2N9Xmqmm
TTQh1UZPd+O++2K4mZQ1JLtBAQ4FrbEyUL2Yweq75yuMnnrk7ja0CU4sxj1RAuIb
i+a4PWNJlCIyhjCh0XaNpJocrZIwl2VytDlZuHz2mUkzia7OfrZ68NH5Nd8P/tfB
sG/RPRyUZCAHNuya1jqAhNy8il1l/o+0dLZBU3ges3tCFKtAxcBPwG2ATLtWC2Ef
f7bjmbQYPdM8+hJb3S/YkrzMGs1lvqqOz8fYZGAQRmAE8CaXPRlZPEvAcqPc+IPy
d8HxqX73EJx4Pnjox+Ej1UFmJIkA3Rwo3dsLPK136BsuxFMucNEG61RvuNGrGb68
sWvG/XifAqU2TprAWDWRD5y8VSaV7zfzJpqlRFt8zv1TKF/Q9oXflawlriFo/MsF
7Z5QferV92Zhkho7CAV1Tg/2Ltnx8JXDKOfggCPzuuE+SPu4g2uJePjadAw3eTyS
XpdSvAuVt/ItbeQ9EsgTpKy7HM8ANs3tibgOdYLZa+/yEZIJODcJNoBlmWgqGQVv
FtM2zjphLgbFLnOIADsZzWzy3JzKpRH1/FuE9V4iVoMO3UGz81IUvAQ5SC2gvX+D
mIjCLD2HHhfpkMJBVDuF6niC7zelgnc4EyCacWkFQGWmM/mZnACc4B5QztSnSMgi
97zFVUtr3HB08Apr8Crx/ukrPac0SS6Txj/Ow7uBWBXQsmoLlnp+jaDzCMrCnHQB
lJyvOZA2o4gjN2g8baW0pjnWVJYJJWSh0x7CqHSrydf6mgsrnYRVIGZNRKiSNX9L
3AMF6OO4fDFxF4Q7nvQ+J6D0cg7p5cbnLZIQY5jvRi+N4Xc4RnaQnBMrPFE3zMxd
QXMtb9H27BQ1fwcr9aUOhK2RF0TnkdoEEjWKrQ8r3aPv9vWmOEpt62WyVSDqFiYB
dcJ6SHIfOfKC0SVrnJFzjhNQfVxTmwX9yoWKgVWq2KlMdR4k/2DhzQo2ZwFaNBf6
5doLOiXH5AZYC+hqcsKKJs1xYwOBjbsbjyOWMLbns2OeG8t1XHK9japQ4mKa+/AU
2CvcVrrwDfSari3Q6HTgFGcKqnIz4BMvJQyJyZ/j2y2Yf8BHjw3fd6XR/oUVZJbf
kBy8g9u+p8lA9Vh+bbAlZq1HINCh0eYlWekk/r3ViH4oN+l31bbCpiuxXQ79Tw/v
DCZjM83qabHwsGZ/HufpJ9jdEWwQoaFR4fGaLdyHc15wEhhH8oXGsO6gDfPhJxPF
QD5AMcoUC7Ag13CLwrgnLLzaaTUJH8NSuDDQBqaUyRRATIWY9+t+sQ/WgmlC4fLh
HgNjSDxiNOTZ/MWrxcjuWkvgSkELziFijvqkvJSmASWCuzgeZA2PUMgYEQKlw+vr
T8p23+ngmeMAbqtl0dLFQ9LHuY7yaVYKECEigQQmE+iFJrqrjVs5DKKKYvLMUKN7
nnjy49kCCxQ7FNlw2nHjHUdhylKKxHGVBeCplWAwsFxCxgOFIbdXYHAv3mBetwba
0VczwVJTm9ouuLBENjxHYiS67DGKSM1qiYI4TwfC7lAKQy8AaDaB7xvLsx7jW76F
PcLePZVppnxEvkjAq0qqPi67U4bZBPjkv6xj5lIkYnW8bbF7gKBIU4xocKePAJCt
LlDgFUoYnwhJvDygLBEt7ICyIwfqcD13sutgLceoZ8naQ40GvYR4vsWg5v76ZEtJ
l7FQrPY0SUhr5sNrYHFYf5MQy6zv6uv7op49lgb2+cQDF9T02SqAcJgmXnjZUeBe
VrPGnkgBfYkTLyE9dgWrwL2/6ZaxUfxIp72s83dxptaTTiLJIAX7UpvL98QaPFdE
5OS/nO6NCFLt4iAivhJGwrUNQ8bUcgoO2NAKoFIZpKK2j5/cV9LbjtXWqoL2izyo
DsRZR/KY341K+E82HNUKy8OKt0bJMZQ1TKXEWC1s317HWYv3XK1zq71Hyke+Bgty
6HCGfY9sikSx7VckTHHgWxdvKI/O5eedDMhBNemBzvZwBqupPatwPVIpTXD8VgN5
mUTM5ec6dXZpqpTF6k78G1QNOaYnZBzjPdzjiDsMIkE2RwNTzF3sBe0S44DYoXMY
LDeqZVFApm/zeAi8EA0/dVezLGPMmhdEIsvW7hDSB5c53nGPxy5ANHLAse9fv2eJ
GPJB3OSog3GiF971y/AIttmXsUjOAyYpMDgSGaEB7PUgRc7kJS9HMq0a6Tw/5y9G
ij3UsZ5gPxgo7k0zhiKTFZR92i/7ppRJxg2OqZrPeObsteBy2mv7V97TvS5ZhG3y
zLK35DFcMABinGeAYbSwTF7hgUnXfihzrsM79mdipjUC+7XsETqy3Ho7srquQYfy
icG+NBqv9/xgtI2XTFA4T4A5VwhuE/1FLyIjmy+dYwOo2U+DCO+R0fNdbdMzB24v
AbeITZoOEoQWR6HyTI4gp/uXdO7d1SqgJxe7qDSsqFkFMR60X9mMiNmkgy2nF2vv
m2rqpOfWB4naRcGQq1JCPiSdPwkOtug8s/mT3rTVOG4Jx0SIbECUC3HVvgS8nMS+
W3J/Cnwm7iKGmbD4a/10kQ4n5nWEmGIu2T4kLqYURO4jrHZ3b0tVtqCdk7UwNlwE
lywgzszTSvJ3k486hLXcVuFCaSoARCjPD1ATQ2juyScArBaxkX64wSB3+QD8byOB
bZjQ3sIRCc2js3BxBRMJLfQNEofRUfIjbSdS6BeLDCI0m19l2Sc9YskemxB/dAle
mL9GNEgmb8suh77ad+dx1ww2K9Ce/pRu+qSzrNk4i+XCbTaNHqBNpN5+kBKuyrji
R66zhiw7dXV5LBDbAM5emxM2OQ3FKtxReem5jhJYzjntPZD4TUSdJsP/pOBcKfiG
dsWLCo/xL2LturrSjoU73dE0hLOjv98YnaAt2JFrM6P8BVaJlNM16ga75AatRPuX
GUyCSmRaLptJTI7A1JM/fDvBzAHEEUAMzvtv9anLVtI6JCDxCZPcoicZb0ud5DOr
gb50yBNk1l9FIcuDJ8Ycz4kjFayAvK5AcGs/HHFglrJfRffT7i9szwf2q/jU6njd
Z13/vZapKMMeRKncVmJWSH8GYpPGTuJLatybYXG1Ei+3uHsP0Y3UreNJvUvabP4B
M3AkE6on79mW5MLh7qQ+DQbnzWA8IjPwt7BkiZeOpPG767BHn3nlv3FsKqAcUrxu
+ZMfCscPy6saRQSVO5eoWP/C+6dnR3EV7G77cH2cRe+OUzdqrEoEaJnm9+U/CHa+
BKC3An4z93HsYdum0xJ3NMy1d8mogS5OjswRxP5dr0GW92VYhJLR0kjqv2JsPJb2
0hfcVTDv9yxn4fQ+6/dXSXROeyGIdKV2GLy14vRLD2fCEPbgcmwgkWTkCN/IfT2I
9mWkbzaRuHIwLc1iFLQQ4NwYqN3YzIKV1BIuXWlfkOAGva22WccZF0k2habTw5wH
LRcAmyn7tzNZiPMeJmyRkKZrUYJQcPjI2kpAMMlm6U5xoUnUgyUqfawGz267XlSX
SG47kSJRsMV/5uEUJG8udg51LotdVL9oqtDKeuVpfUd5QumBxS+FQNQRFcz9j166
CdYiRjz63407GDEkQeqVg+MZR+mpt/McTkXvLdXOGZUr9OuSZoFiuC56U/Q7wt1M
jlXpXzPhkeH5mWFyo03Xa9kxfbgAsQAm7BHQWoh23FoU60w95HewC4bcmvQvN5nl
XR7xAX9jRT8zqNtGI3DruOdVzgYX+NBB2N774n/Ij0MetjZL4lZc994Y0iySOZoZ
YbxpfjOitnX8dpUpy2q0cQy2oGM+Hhg/8bgBAPy+nm45kZ/EdHuFwER7eHZzEDTo
T4O2T2N54YOLda/HeF5OXLJwQwGZniUMS9xC9s/H50s9sQInbo9+EQBsOM67iv7p
g7LWsWSHin0kGCRslRG7Ayc+x/N/fX7MYaqfAYuu+XR+kLa5BPoUeLUGCkJ4gwJG
hl+FEISlDncUXLTv72UkELFf2OKZte9HhyjXm2rbgvDQCZLQe4PxJp2iUrlxpIa4
gWiRkR7mPyu4tZ1JVnzK1glZrjBrEngEsei4bXM/OqcibWSd0aljqihm/Z4Rp1RV
PwWqXJ+R5CqeCgma6LE4aPT+g0F5tmsRu/JuPumeTkZjYEO+cVbThKE2G66lwETg
fKyx5Wtl8r79wX2RlY0XWUWrxxPgHYhGmqgCHL+oKOXo3LiYnQUQHR+taacuS0bk
fw9UPep1kVFQlKxDhfWHZvGahPaO9XW9/kdvwXg9xa84m8w14wKR9DNesL+xxtZW
oI3jGhcjf75r7XxBqoFNRHZ5gngeYErmQxFvgqPJt/Fnh/aUemOELp0UguOcyftj
fmIlhNB56v8GZsIk9MpwK+OcZ+Tlv2n9n8jXjWMRW89r1DIy0asuX4K3y7u++teu
x4Rm17iBKonbiP5QJYiOmWhr89tG/S6Z0BIbtLInxNTwx0anW0EBsrebOgr0/CIi
vZQS04lp81Yb/3rjqveimnDhkRXnO3Xv2VC1Qfpf7hpTuYxCJ2IQBPnVt3cc+XBL
2ovtlMnw/svVw7IvYMfX4Euv0dSF3Uo+htxp/cRLLJ0F6pjfHr/sSUHUrYosklkc
D2sTaXDvAOAyjp1NmQ/sNaKWPwa89p8QL05nM2QQ7Ld3jvceZQkeNIRw6GDVcZxu
prmthFOiWh8yyBrumLqI7BQjz5rybXAfvNLXlado063tMsUxEu77aWw//z9ozEfK
Z8cJoI/6Ki3k4JRRG7j6H7/591JD1wmbierkDn2OjY7WztDiIk3N9L4ZpJRZkhGe
jSDFkujIIKHYzNnSPvaVVBqK3AHT/xi3GeGGJKu+QSxQ/vV4hd4sYeN8TPsdfL7N
78g5Q7eMMCL3PTdlFvX5VPPLO1DFM7NHZviA5DXNIsYDSMOIEbvKJpf0+oH4C+lc
GyGZ4wFjrBNvVlJxkVXjDfXxr5hDbR0YmDhmSNSEUyZY/7TL2axglT6Kl0JxrdEh
UfMmodPtOeO20+/n/F7pYl1mB7lqGKXxm2ljcia181LYwMZd3h1egKiB/XCboero
HC8bSXASI6JJZIHLxasLPOiFLmD6dMYfFsvxjXCxUigmy4gKwVhAoIUOACh8znt3
FzrEswomvsApgQRd6ThzLm6YREARZVD5mCKrghku+M594WQo1hxp3e8vnDUAE0v3
GRxE7jpKPj73ZYuYVoNy9JjuLKWNId5hgc4kUmxDiL9ljLnHNgR2Gi+mo53FsLiV
cJ9+qGvA4/m32iyk77qXzej8VL/4ys43o9pimnCIZ4wiyYIzD+wu6OfaDds1w5Q7
RRRStBtQkpgou0Ju3/tz7ViFmqiqK8Vpo9yiABfz+AW4upUdLNGo4i0ZdxtSD3s5
D0viZz+PXvNpK2nO6CW/0fo6ncy4fdWz+5USGVqX9rqfKCUAhiZ5rjgCYdH7UouC
O1AaXKGmGVRYmQrCIrb6mFhdoSqbV3mOt6YaArm6IWwBoDDBPxz/skZksf9CGBwI
tMJcW2NA6siHXRyj+mrcqbDKP7tWHcs87dDKnG1BDQT5FjNYXdZRyrEUQ1u1pEb2
l6bk/SnM/YA6xqcYzdLBM2RuHKEEMnA/uTdMAZ4x+LnhhDqDvDvaXfO1TXUIiqWp
PPSKqKIMMiklCBrERXsCzhdL6sdq/bevIzml98cKdARBXq1FQsVh9Qf0smpTvlWu
6QLxJ76VfISlN5X9uARdpey6gWJigBuw9RhZALm9D3YRcKS/wLInUt/KQvzWMWqq
QvaVWLR1iN88z8e9kuWwHJHTXtaTzCYGhDzXPlZJAzje4EM8oGZuFWQhQpVBTgZb
oVLmWSURlJMfORv8wag8tpa0aAtUVZCF4L154KneJJ59nyhSKVvs3RYeoMiMjOaN
cFjUv2WrNPoSB7r5lbpeRT5GsjMaFXTQVWPYwHh6U3VpsNK4YBjrK+hCoVYx4/1K
yGoWK9DPCdnB7jM21m57vgnN0+2/kQAADU37mXnN9Zoxzxg+xc3CVMbJwPis6qhA
evzP+CGTSp8t5/bzbYDPqm8TuL8svA9jjF5VG9ZRyPgXn8lGExaMnp6FbQwy4FQS
Tg+Dyo6lbGshg64wcCRAYaWLPpdeH5p2KG69PRUMMWZ5nPEPhx6rpUpQqKcjrIpv
a3RqbQPizLap9qtTAObt61SZM3c/j4vO+V44exXyAztP7TlnJ0cyZ6sK6iYNUl8c
wPbQWBpx2bG/CEdNuVIVoAI5EbxtQUDZOoJmmHennlnAl5gnszUqakJbPMdBaih4
NkdE2sz3b6ZwdHfY2XZd3tx2d/45jjXzOQrt/aUsJJdXhaWGIJtyu5IYAuqb0lH9
4KEZ6pM+yu0IHyOE2lCCv8ySvQLVqM9PfPNCxngGMqu/a00H6ll85ggVn2zxYTfS
nAlvOlP9ShxJ2pa+thzZrgsA4rc109tjNGSPFFU2dj1Czx9qz9RL6d85owv9xSkA
orNJT1lqtvf9YXfJ1jtBZr/FX8tzosSuTSUbDr8XD0WIRFn7RkkKbKpWRH+UdXhR
deRiSQEPtJ9ZMAN5qDe/iB/vElLDUM5byMQOfai1Lmtl7ZaCYNi4POKGUH5vspnt
CWOoDG1Eklg/Irk7nX3BJdiagc/KKkUhHHLKIwUHtYRFjqcRKjLtCxJqv8vaRZLN
XgyWYP5A8UuBUogRIJfBJINZFxZM2CCL6Fc0hGz4uy1Zsb8M+tAbtHX0/w4hoO8D
dhj6SchEguiPrfYxF6pXpGj7f1CLGWmeu7oeNXskF7yBu4yJDeklnu/rgB8kkUkw
tb2akX4LaSPYv3xyKR2IG71oZflfs9Cmv5ssTGv5bS6j7VGRF4qQ6UgSTi1z8mnc
e3bN1ONptoo1XpD4SqmrU8GBbvxIE+ED6AP6B1xVZcxhClpEdO3vmR1n9i5pmmL5
T/tVnqf9G6jAR/3NYMvbAlQEwVAs/ou6d7uJ3lVjFql/ITLW2Anp6u7LnKIYfNJF
TWYbHvV0X7ccyNyy5GDGg60IZFrtQq4DqJqMFprBCI283mc4JBpvs7jYytUsGw1N
G8qD7btVq2dlOn6qcKg2k7bQOHNdNI2bIZBPEOoZnXUoq9UKvZBmfN2iwatFMfJp
HHDnQXpyZW7afMGBtSSo6J2KB/sgDWCRY0WVOjzaFv3O380EHcSr0U56sDK8g6/5
VG7EbimyUC2Eotsvv6ATSz+z21kYDat1cNSC+kV5DyWdL4bgigBzzfj4VFZO2nMw
2QH7ev/sSs1Gik4XMPvlQnPhEZUBB7VsLIyw710WEn2W8qrcHxx99sX6TrYS3XaS
By1Usx7T+Apn+N2IYIqxvXrZpQeEuF2IMLwaADOM/PI8whgPk7PvzwVzUAJMkjNT
92KGAzsG0o+yjZ2MPoUSVP/P/RJ8ZCp6Vul1thGo9yVt9Yqr3nXNwn51zqiyPSs8
qxNcxO3B1wv8EBhFTXd29IHq2EmqaOGCnHNRbOkLNkxwRof5R0ytI4BJAgBiD/mz
HMxjBnvOF120mQAO6ROPza/4bX0M+gcX35G5AbsETIRLzruseaT4kHe080tNm/yC
m2tZpbs7Z5b3nYOlc4l86a7p8t4v4PC4xrbS+HvUZ1jgLK9mhZwibrDoUOFUPTJ9
5pQVY/DwlBsZSivdcfOoh0X7YoEU/sZdj0pSODqQW2Zx2BPRDpjwnAx0qON5A09Q
/L3r7cifQdUAeRAv1+bHv8I1QvApN9hTimE9N3Poz4HORxTPuYFaJ55+r/WzJ/Xy
K78jvyeW8aFy7Sbuw8SyJRnlAeZuSTuuz5aVSMy2dVhqe6qtRMADG4iDpEdecbJ4
tnE3vtgja+jsLd0QMI5D36C5bYbTk+Wj+ZcacOaSB3aTxEVDdGMeYb7PmV0LqQq2
iGTw3/51AKJEqa+fmRnNBQ+VqFw1gcDmVFMMYtKJSZndVk3iEH8YQOeo9U/4356T
IM42hVEea5AwPkK9kAzlyX3COU6ZGqGoeDbkZe1mi+gl4IBkPlbDB4wOu/ldxc1F
DrOYuqFrWDmTOaIy4MbAYsjoRojJDzSVyniSVQKvIUtEphkH1v2++OYwHx0dCIHe
52PGDHF9X6gRCGRxFAgpcZC3P7IFA3ll4/qF7oIAyhEYKHqjMNkJ/GXguxvwFBS7
ttDXAORj/q2bqWZxunJ2BFQ6o29bPfvGegRM8BQyQCQvNgeil0WdPZqL119G0l1x
R3192vu5JLGU/pyGF9lwdtfyhxCU0egvu3477VfXzYBleSCV5RgrdHsn/qTgqwGh
GGOMM6VR05ylPJZAGmAsjHZTu8Sgzkypz3muKYeqqpyNgOHHzMBxxDRJX2bOnEwp
fsLqy8JlQZvkegWg2Qjd7ztHilRnBkNdQWtyOj/U9FhWWrYC+UpLvG80OoMnx18t
PlbC719I8rkBrXw8suYVzbgl/VuAxXdAzdYKXsxkrtlrTUlR/Hvxv4lsunndduN2
us7XCrmo37vV64BwHf7yMO3ccyYInUCdhcXfyt+a5svG4Mce+o0V8K9OhvqClNBz
qJYBTz2uUvPrZswBLb+ba+HppMHDRuhsV43H0YETimEZLKZwyBtDiLyJS0TEjpsu
vJ7QAY1tID1f8Gg/mTuZ48jSGe6gY8I5UdpPvcyizFMD8SH3APLpTIPYI8+2O1Wn
U/CWIJm5yBb1nrM6ZNAraz6lI31rbQjL1UmwrQkJHXENAmZ7itgA24IA8wy6i+GN
u8p1v2dC2FfIyjzr1MAmci3y8y9kbnyDduGTgX6UFPZAFNvZ42JB6AsIr5SlE4iL
uHR4iEnkmjUMNAfLQOYlVflTsd8cGnM7wyZr/p47LvnbnUhvUIBrouSu+p18A/h7
9V7gH3Dm56WbbT2ZZug6WTunIfTQAsDIr1XFEd04ZIef1yE5RGOLAeV+ZF2giUq+
+hEo/SzTQRA1+wCRfpxyjMUhBMHBX0WHXn8vilro7FYPm/JveSQvgtFyv+UfTYtr
ZNzLZiasOsJK3csRjZzNLGVdS5EvEB9wWL8dB4bdJ+X1gV2JyFLo8HBDu0iDcRUG
CFmlVtNASSobM8aZyjQkzMgpMnzMrtYjnPTu9CybGIp5dKUx/9vjOP/h131C2FX/
so1F1jgElRSN+g7dm0FKpzA9aVrOxAB/exbANzNPVnH4HOIF0R4HiMUT5M2UJ9Kk
tcVFjKQTwnfTKqGCeEUSWm2vyR+srd+Zwfq9mSD3x1Tpq9K8fGybFVEMty0WNWRC
CXnycrq9mqkxkNdFJs33a+FhQ4gG0odjLvsFbXgF7L42LRLKbojGlnmT8kLGxiOj
RlY+36QhFBB0l7m2Vf+togAcLntx7Z1+I59v4e4ZRPDpKjMuonm59VxwN7QGX8Bo
drVntysM3eFNCOqSAtWt7sSlkS5u6ikzJVXYaEJJk1bzKtZ6CZCryIzZHkPWXHk0
v4xVm1hMTnSVXWPDxR0TXDZZb9k5I/pnJ/pVeG+IO64t/SdkOrwCclgeVDQcw2vY
c7gVp4G1SeihTRRLlMQAkrI4nnqGHQcwxgBgsunXcCyRaikRk3s8SE5F/LWXfmZN
tmGpu31O7tYTAjMIjMX3Y2f4sfuzKbkI4WzZ2baXKmGFzAoO3vObZot9daS0KQTO
N/Sabc34CB8Ga+Wnpp8t8r0il9nX3YZUI1/dbvfqujP1oMBomGqHNHrcyAemxu/R
9vLkozxcW+7MeH/5kmbNk/bZ4p2MQNeEzfEInkrNMAGPe9we+wCleH/xuTyDsxwW
oRXYUOtbYGmydwlEpczD9R0rzQgELqZeglMFyhfhMTVKRulixjwTRgoPz44d6DcE
U52H3WtoWqoZ+ZDLVryix1U9zBtcH17jWPng1cV7/NP1ZDALCeWYt08pAR9liEWr
0XAj+remrV6gKPtlszZReQ451sDM1hgEN1TSUZ5p1L+6mTj2fXrNHlemxnmPoi9E
0+GvPVt8NCuJQuCLuWj4O7QxEqr5J4Q0g9wDt5yErPqtuzuJN0/QGuoruSDlXDC9
Z45njyrDQuVGsu1tzhWjjZiAik9Q3JyHQlybr+CtbhLFKEgP8knBjF8ead2iEu50
0eaHi/uHPCjXUnt4tgK0J4Ib4qAwLO3UAOWFFhHObrTecHjpZiqJ7FzhGUevjgwc
R9xJKwSRlMMoPSzAiC8nuq+2Xrg0HS0dUPteOkhQ5CRNDb3/YH8Q7Mjr87PtVIwb
JPI2xA//DAYvPiDydE6mHup56jIRtEmm8zLx4wI+8ikiZNCTPWoKOsiWf1AOVlOu
wKmytVpfagG9YekbXTsYc61ZaLh58R3RncmgXZGuSXe3pJb3xcPZSyqsIo+p900Z
GrN6sWE7ErKYSd8aExhczIpBCtlRQ+Oy9oExt4FSArVRlh74qMhUacXJFVur+taU
oGBnsZdetIcrqmXWGPYQ2fQLikvoxfS9osB0F0X8xxA7vnoynd5OyFXyaIu85YkU
FVIRHZ6yksE947s4vDVExLar9Ti4NfhvWnAYGuSq3799qr73D1rgZtdt0pJxC8oN
YNEO6rWBDTrxvoYHr9/5qmAOqGhN/cChNsqvTO4iN4HzoRv1It7eh6hhLEVKA69Y
8HMEs6wMhfqBfZ22wffLPxbEzrv4tKdVeDcw/FIsrn9Nfwp1lkRTjyAyJQXk2ZV7
8moTfhokaIk56yME431rzSXULr2iPLCbTnJEuWzy1YGvlrq7SZUFMvQgyxk78hQC
crEc1LtVsVps3YdSPeTxscGR11UX1o1WHh/Nra0JCpS1AgId21ESrSUr8Pkv/X/g
UykXahbQU+4EW0HLgwVQa8dKWz21Vc71ZFZKMjm/x4sl/hw9erTetAlStcGaDo+B
Rzf337cOKyBudBy5QVKxbO1MqxJ209ylDZ96jkWoXTpPsk/iTaOfyXAxUbFx12kX
ck6NuR2Yo3E1rQq3wJ25TZnOJ9+g/cJcf/9uNeGDpEh4ml4NoB7HDa5UXKAyr/f2
5lZGU8VrPNMcqDk+pcHG/fCwypZhzJlxwLTFlFPyDIVuVpen4hbC1RIeTuwg0bCr
jJaEDvK6UAyNwId7NSg2hEW+wGxfneSKZNOj3fOuDuECkcrO0GezDgq6FrxsT+qG
9boU3gN1NDMzMAgNaDir7hIttHfdPZwSLzmMfiefBGbI/RpsAIE3+3WiwFOe5RzA
nwlKiBwLZ+KBR6ZS6Z8KfBoM0rs6RfvEC4IC+IPj1UOldf8Ar6wQ/NKvbWVIjL9d
I56SWxjO4jHF29dFtNpKvUDMi1czfnupublcEDgiXtpRZj5o1OVsfKYWE7v5zYt4
qzDAgzX5V+rE/fDzcKWBp4OhJC3V6Jouu4dCgn5py41nRWk+fgF35xGT6yaxcqoH
X/SA8m+VZ1/kAZ+fe/WJc/1+PpsyReKkTmSmErjWtsWyXqJ1aTmwjtQtifvoCEQa
z6tGf5BA//HnpFyAzlwfyHwHkt/tlar3I62UhL6rOH2BMivRq7ea94Ox8EbdoyUi
s/DXouPJknSIU/2w2LGBDbp6fas6HPRmh6SwdLuK3wdpQrmQN8F4Mz+iO9QJy5NM
8nLzI08eijDQtdPod0unkL9TjZME1rwxYSW6v3bloJBB/s8K9Ns7ZfYkG3rZ8OQE
+chwdbMRdQT1PiKvapC/4oURF7t7je3X1v/I4KnQZNuvi/3dSLBlW/rONETspwZW
cEjoI4XiKz4r3fw9bhn1/LHNV1bDLxEq6K8Q1xO4nRaGajMPCwiJ91AQP71JTy7U
16kI2/DPhdM956xZrg+Zl1zjZjGDozfGUYOcE5TKIWq4/UQ2DMpR7Yp0Cd3q9dkQ
gLzgDSC6GjcTaZBo+5K4PYd+JOTPbobYzAZhQkcRX90agJXCAdJ8OeVlkurGGvtl
MJsPeM94yn0yOSnxuyMkem2wUYxaedKph5xiS+XuTRWIHfu34XWkGnhZQh5PIcNA
ch8S0lym+RrhIQuJA1/8t5axJn03W6jJtAyLYGwdukONSpioDLCTTWVOacPOG94v
uESI6e0IglzD3FPZe6CEjz9WQuoZG1Zvl4folOpnYbY/mc/3qx24IlEnqbaGzkqw
Bfa/by44IWZz9MsdERe5hQ1tjREAgGyeKcPARDysjF0bEqpgxiMXM+/yRuIJcVup
y1U1BJD+shqzUNjOLEMInldvsRRQycPh7db/zwpa2l5trojR8j9yzTME6nWy5OEK
A2dK94WOFB+SXggn/sI9e09bSAOdJ1S26Io2lMIfdwPOSG0apljmMNezbE0Q5mQi
lSfm4ArylH4bJEhfltGrpkMR5YlscoVnjyTLzxeyX7hPLWfjLZ6qaAhGmDIs3JXg
4EcS8OsfdTrpM8cAsInT3TL2IJQD/Zc0cuW7XsfQ+2Tgex7HZzj2uaWK55gXNkLz
7cE+AAXDszjJPVduJ+iHtvbR/G+8VilOvXEZII0Y5M975IB3ZNLIxCKm+pkc1MW0
vj37pSaoLyfxRLZfq5kv260fTlV2849p/0OCTaGonYBDxe4wkZKQhGyR07Og6D1q
jRqstue0U4hofkqAIRlgtnuXuVGDjYdrFVWsnHLQfnYUYRhgm+BLo2Lx/gOMVXXg
D8nLPOcyoQFFZ51UBfdEtVOicHxqPwDnqSEMCn5fysXQn37swbsEELih0XbTLaLt
PYhDgso6odG0tKBMy3LKq0iMM7vLSZ0UyxtchsSwek7WlNIwOUio2Uz+PMhcEhbn
lFut53TwdPtXsLsIefx3RTUsoD0QtybFD3hKUfcd9qky+DEz0EkyAEuV1PgN5nPG
ZvF7JmZu6T0togRt8P/G8W7ZOPcauANecmijkNzTnE337U+21TWWoDse5ZqZQpaE
1TAWF7loX7WbLxngfYI3DwY5oTvvfpbcBuXtkzTDYECATgWmwMicQbofwMOaW+k4
lBTy+/yU/Mb2IjYUX0zfOXTe0Ds0KogGulJTlPRXIp3efjrS+qKO5P86y7PZFiKo
HHpWmKrcGcozsytMXl7YlRe1W99PEv1e8HDwkJnv7dUvzfPeNhhQxfNQDGphSrAQ
6p52OUTVBtL/ypNWn20SWoEaGnAjvkIOI4PdUOT4EF3bIg5KYt/z+a2Kz47xjSTw
0K/BAvkHRioWD+DBzTnMH450qANgJQBaJmvk0k+KOl69s/iDGBB6Q3IF3Ai1uSSM
t3WsJ0aX3CghSJDQm1hJ+SrbfEDL2huuk3gvC+be28FvDgJnhd3uub5PH9ymnuWf
1CCbVSdHAF7KdzlzpKQQLZPGhkn/uoXCvvWm5F5FwPLLrGAa64vlaVNPiLFFErjf
9s67xUoOC9sBlwo9PkWTUnWG0x71EgO8st6yqg5w3rysgVPQMvMQ660JoYFoquKG
beFL1U0Jq3tkptfcYj6dST0aswX09EHLyBcLC9IOOgF/y7w0APMUWw0CofA64xG+
QU8CF2/8TlH6hsqMDYIvPehAEiOyjsAxAGGWSpT5K6N5Kg1C92go3dxZooCxbyjR
0QnLTzZcrOEr+BaCcilu7yfoOnydGxYM92/7RfF/6xCZncP9qWlt7aTw8kBqreO3
1cpaMEKmHFXOORqq7V6eRBv4u5yVBT8AKA1U/qz3SIIhwHCi84be1Gmw0A55ghel
eyakqMjMi2ZHDkygvbIy2pp0Xzr3s9uRw2fuPZNbhIrRDBcTuiYRQAspIym9e9wX
He8UcL/Hc2T14IF7Ewj0hHwMpgzBud0aUTN80JMrwiZRmTc66p/nwJTyG8kgQ19A
Ut7omgxOWy5GWwCBA5MkoPlDKKLx+2sASe1mv+QpBgpMJqopm3ppNMDR4iAmbXsC
PQF+PYNnhMfSjjr++sKpM9q/Pe/ze3IJX+E1Bxx66q38HzYIFOVOv9hWsmC6QcBP
558W/2fpSRGNq/XxqL6TCYHj3TEWg1rfPkOemFikObwQVbndi74CaNx8Z3Wi5bh7
fb+gZtXSIanFmbpd9doZBhxp1n1jOlpyhbtr5RhchLRD/Q4ckgmKeNX2qG/34pFz
TocGSt9bMuMJdA1F8aX9FSLneivTAhotEuQbbw/LXGoHKtW1WBM/oCVNmKmQ0jT9
RtTnTYlKp1YS/+xoiMyiOGHw4R0eradbgCglBabYc9mntvlG6zJRuxQNvCyaJd3K
KDaQImMf6tWiJYhDLOlumDEUzjvePYbFE8owg5+KQny3WmnN1mlIsF1wcBBx6J2U
jiNjKsl1+5xG14zBom7EAUTkPGznbKKJzFvnZ09pEsnu+bGNknnqtt4+KA4DJP6R
IetKREFu0ZYxUkEgsekdDAQvcQXPLn1lI57ICWfgb6FWKZvYHwXzI38IMTHRlOnl
s332cUGCHyRWfCCHcKgnTTVKxTKVJ+aP2GYXihic4NbL/W7Zt5enc8EoE2LjQ1gn
Tt+D47flKGmLWmuFN2l0VlJfb2/8zypAL4MoO/2Bf27H2x7hPLKnYhNYi+oiGRo0
0mMY0a09GZ30BJaS40bHGPaDfoeTlfycXANBftrduvHafe68Bf3PEoohaPIaZJa8
AuPztvVeYH0BzBreO9+MNgYQ2kSR3cvOIZfca7x6eoxnVyOtbmUe12vl2/pc3viX
oLSKVFSi3vdHZM3lZV/1zH4Zno3h4f2It73QluFGCpZHBNsrYRd6qCiyQM2ftsVJ
MzLQkXcF8MrhkhJJy7eHXCQheC1V9F5g0o8J4exJk8ykdAkgC9kxaRiXFb8894h+
odi68KW+vtDzpCPb0BXGxD/+SwwIplqipYvHlNNjedKG7GAA/59jQ/BKOXXlKWEG
1Gp0VAPNO3CBFiRW6fOtuBZqnm6xTj1cw80WahtEIbYaslwB6Xx6Esko0mObH6HJ
qJNul5YTNXp90VGHkY6yBgHlZx/uibhckrIX9dK//xNP1d+AiSxQjhkfP8VkGWZF
e2ljQFSFVbwks1v4QgKA7G8lJOVGe5tLX4mhKedtOKqR4VlqzmGokGKp4mQ+LVsN
wKkiE7UzcX9Q8Zlgkz9gjWlnqJfsj/ZntGvAH4RojgTRzyT5jXe7MFOHEo1a6LVh
PCwaioNY0CD3qJ6ISNeRl03rid7uU7PwEMa5y0MY9oXLdh+yICPQcp6qohtULaXI
iwJwqFjxLhkuPH0TbcRS63/8Hb3frvinQsTYuRkoznZFYrW7g4/cEU1d9SQ+nC+e
FEelg4E2L8vLWyQ+aQdx/hz9hHlhmH+hhC3iNy54qFcawF9njxaYmlJj+gEp05rv
FB7mzs62fznqY5aaxGEv7u/j1p6XkrP0sncgIBqaCFw7iOSICpZLsbwpoYGqLiyo
DeNE8d343Id5a1oHGJuwQuW0M7KldydE7+Bi9/XRZluH3xrw+npqfBGLxln7mzQY
iZMhiV5tdGO/j87X4I25C7hNiKu+VkqD9GpUEx2yRP6i0EHGZzsQ3NOyndVlll/R
6aLf39+WIr2jQ1uFm/SWaEpKJ9PxPm5+VyJojqLvMdU+ct11gVI1lCe8PA+d/2jn
tWk8ZDWHJiXybPPyoENRFCq3oZivhjpYGbBalX+2R4jv2P6HJ7XV9KFE6SpaY1An
op0rhhdUAv/pxQkCYNDqI7/6YZpqebC3Ncc6sBtcfr5oMt2Rge60/qCgFVn9QqOx
QTP4C+96sTP1ggXx/AMb9lNPxQhvhnpvnHWaFWS7P3SoGWkC7Zx2cO7KEOpKlGAq
HlSjOGMqIurdUaV/kCw7D+zlaZUjLZsnodSu4WqXXXtCbZ1gNCyZHR84bzXiq5B4
Ms7wU1haVJVpihCMqnnRIvSnM53z2PUPAAG7abBMT2dkX+mkgUFEahF2H9s/sGpe
Bxqv/+3pmHExKRPMOpBw6hflHy4QTZJ4a3Ekpu1F+jm0V5QM2u1nBD0C1mAHpGaq
Fw+dG1RQl5MFvi2WB9LgK2vP950FSYiSj5N1NpoLpvzzobmVlYaYuqc+txyrHjUY
iDFOeCz31746NibggZf7pP4i7Gw+uJok/76nJtiwnrwFlr6JkC1zQwrgBzISOo4F
elloFcDpD96YCIMLnt8XyyCa/qrw4NIC/YJl7Et6soSn9pM3rhFOf9hY+51M1HY5
v5I8v77A2bcfSJFhO0wSz3UW5sUYlMVMu4Lwij8HkwLF5s1epzNu2r5lqOjcfYaV
JCnQPvvn8IXRQdSXyk4W3hLjoMZzPvj4w/9/OQ5vk78/RDSrhvpcrhmqReN2f17V
YzeTAkA6nj+lUntwJlKpy5VC3Koxa9sXL3T79vibLyM0fpCELgGMEyjjbGI+jFrs
dewjrgVDXXec9oqcOZU1NRugYZRe31MxYHdz9K0Eni1UlmBPcyMmf4dTuXj2+0BC
cCX56WPqggIcAqwwvqF5PxtjW/VChTpi4OVgyLAfrR7XEYG3hsQETf64dB8QD4zb
Ido9G8NBcDuGi/0g7noj/gSc4oVYrzLsZthTjySfaw2QzZ9FTVha6MZ4/br0daN+
zcVQieeXD7BKHCaoK9hHkEXlybzM/rX93fsPeNF7Yar+kwhc5KDbGtyU/hnRx1Az
IvX7RkuRFwhO6P2g0RnvC5xbWzzRg4nz6LE7DIAq7q0b26YRBt1EOx53Dm5YO8K+
n1buTt9nOBFzsPMHusdVeOY8pYElQckriMG8ipTAlIz7tXzZ0SRCCV8K6X4exp7w
Qtg8/d9yCNseMfbMufjKvBkpXV0f4WwHGbmnUl/Yvz3jO8JjUbJwK6L7+0B02Bc3
hB6JuCIYMlEVjqv7/vMULDFds1sQnePOkNaJ5E4ydxiiLMjLkl8aidVm8UP0a9tq
MYWFyMaEGBOkOxZnvxevQ09arSna4NWK4q+rnRyY4KR5g+R5ctEfRFYTzExyn9Mt
uSGUnMPbvHKEU4lO76jH8IwZINPlxdH2SIszw6+R19Q5I1dcrJZyjrqQx8jw3ccA
64YZ9S2ok7QIRkCetZtB+56PPYFm7U2PwxSUwakVZ8+No63YpuDsjLIzx4lpJQvj
+A40QSeSz6MxWQX9Xb4R74REW1FS16iON1QqPccq2rlYdDBRVtwN2PfF/B8j4Xk6
HLUlzHEVQolude0y3Fs6xFTdF4hLh/FpktvusHbr5WE5I70ceVOhnsQnvisy2jKY
rciAAhfEDlNxIAL40Qwjo6leWPRXnRXB2iMzJuxorU2uP+7SVWnpXJSJA/duzP7h
SGXqebEidH1nqJ28xU+zVyqQpIoT3jCmg5aD6A1vF4DL4c8fgm9KzLe/R0fBEbz0
Hj6QumljBoxOqgbvcPE+m4HC/U61leIKStCEko2HC4pJR8JFf6SD35ClJ6IIkoTG
eTMWGf+iesZEB+bCcid4B9by7jHBB2F3XjQSYbeHFSjGtO7GGyIjyqITumHdppua
q1hcQzJkaxrf2Wo7dsRH7ah6iXVuMTooNya7nxWtnO3ru7ZDCgAA9PtvvXYkI+4n
FOSWGnEgz4pBvn2cYWvEZRJTagBkYCXPWfYKeAckOq8sC1NamJNeDsHRuiKq9djp
LfIJt7550CL0/+Kvvqp1ZZxNmsTsJrRa1PBoByrJS1F9qp62uo69/YXBEQ3k3Vnm
hdRvtO0iSgqzA4UOdlwwIOhGIwyzbTV+wjbNXr+sDV14/RqizSfX+PQR+WVDYyWx
h43SYRUzL7aKZD3P7gjesqSLv+iAG1iw7NPJLuMQPXW69qdlgvs3GvH5did/vuRc
oWNQOGgPxk79mpvH8hu2pHw0jb2o7M98Gw3Tt/rTyaQTlXQfdrgt/mzJavp52Mdk
1+NNBAfO29phlPCzk7gwXWZhzhWNMU5SZnyojfY6Vsl02cdecqOweDQyejv8+Wsr
Lgq7RwTyvs4qX5XsgsK5akPHrQeJbnzD16/u2tSSh2VHmsbuqzFGMNHIAtTjrdyq
JJgNWKdzYUJV92lAADWM/Cg8m+jWzrW98KdEXdd9V/NqFnKl5JVXcikaqsWFnJCP
lHtvi77/TJgSJWiln1GjvErGXIczSDFqF4ksd2ycuN1lPdomfWi5wGb0GYlNokd6
0Kuc0DEg6g+xLnF3zQTk9Vg/dsbF3Cp2VlyYlUPt2TiLb8oGwEEGB45rIGflKOG1
LkxFcS+cKAln9sFoe34iLCgBXraFhK9DjmLe+fkorK/oJpRo8BgsOehejtCr5lP9
H74+MBEAiHJPyGLVe/hHrn62rw3ePhCxynbRf5/r8Bq0h+3BRwULGgfgJVlQYlU0
skjcRCUwhSPUssb0HVeJqGsHFbkRpyLz7YNXmLIVTIVH9AahN67yViWkp4vVKra1
mn8nW1IYWUSw7FvPM6klZHMVTjorwDuZOuU5YHjskzKjkGguEoY7VLDjkdpfk9Ik
nWZFLLhAwgWoKUEwq+xnCHUN3uv05n85kZUdHiTxcKHOEa9GcbYUp1i2F6+RQnJ6
qY698kFFQ4u7B3HH0nhKivFgAgxQZrkQ4HVifh/RNwbPu/v8CdpNBzi0bh2Zs12F
p9wpK2+Fl9s5nBqDFQgd0J1QNpu2q4ECf9ac0YFmTc9LwwVEv3YWU7d9rjAlEhVG
1wqeUm9NwsegVCFs2s5HAfe9fbbtEA5MUMKKb3USHFGxhEJEUGsWQ3wtZ2LEH2Qv
nSB1XiOn/MyjYoUgDPNYtv2MC6sNSjnEHq66QES0F4Qul+Z9hlloPJIj+qd1RyQU
J33yO4MSZBZuugRgZJ1KS4FaouPPUa7WWq0iSSrm505NsT0hy0f43vGflknGAfPi
gCgED7Ossuv/oi45+TyJGvLp6VJDrmDjaHRqNPIZ6iVrBkthFYf7kZmdBxVuJw3o
E8KkjdnK9EUchj/EjYycAnh2L5S4uJn8be9T0U6Fe3Gkfr8hHqRrSyooA9BTxm5P
1SpQhOyFJo5NT87xtytP3R5x7+OjbQQgCOCtBRJYGpvaQ/ufNjWwNsC6v4TgtMJ3
wy2cTporcYSPhGoptQAhPYOMdLodK9l79fvqIu2bdYbtfb9Y/sQeCE00dDaX/+Gd
i61maZoKUBxY4DvZ5TOgFYasFtR2Ha57Rik8I48KD/svsbbhzmk8LUZtaD0spld2
EJQQV4E8hDHaYRzyfHYJS4vMhhR25sXwptfrKbh59M39zRO9PDOEJ6jWv9Z2crKy
q67nvLc3GFvjn+8m5zcNSGXZmm5gUuvc/vuWYJuaIktDBIFHFkxsgdJE28w5p+Uq
xNUngfxMz5Oxr5+I3hxUj+ScfVHl97IJ9eAEHHAtPY/dBo30WAE3C6qw4o/GmY+S
bbEGB2HOo6AATq2yaqHyrTMagDXq9nqlpxR5+d6cze1o4MuS5Jr+6RGj/DgQ2e49
0miEoB3CZlCaZzro3OERJQRgnDq6nZQu0xSGgcMkvSnv7mHfVZYdy5j+4EObCH0A
yCDNItxqm7lzhvrApcQQxnv0qc0lWkEqFd43ePLEq6b+dUkHXbuRieDX+Au98i/j
Lnz1zYyCyDifNbgy0FCabehAZUmHOOTig3z2GCkuEjrGb+eRWXwmU8nH2kwp42jv
tjXZMvkzsSgpXIpSV6glu/jPoVqzsT9lQ3sbi5z+nxIjiinDP2wDPYLakgpmkG90
/3yd4GpwFopgfvdeyRr9QGOPiimpw9HoEJIOe0u6rzc9B6l1vRA/odONbHLftMam
Up2UmPAftUwoarwkCUSGS9W5VTMPVJgERZy+0RdI48hQJnKYMLiY4qVIUG3Vf5+d
+eLchEPYxYk79EcNJk0K31/fSNLF6lvEJlpEVSNYaMeH/UZkgepveUoUTYetdYpe
vltfLrtVhWboBPWn2Pott1itz6nvKdACjWSijBfntjE8TM6ztgG/mKEFGkaHJz9P
DvLwPfdwu+vZMw88pg8r8bZbO8Lrhp+z/r/uzn9VJhmXTqf5UhFEUY2pYMt2I+FV
i7XW4ecWhQPQUK4UFAV+J1thpQPMfZP+kO/Q8U6MeHoeEXZvi7gR3xaIq0nJkzfI
lmRohHh+1RGKpjc4Lgh7hF715EIGo0/hIAX68y5fpbAHhgFUE7PJkbTSFWsnvTlA
QSJXaOWmNe4KXujWeEzC6iRnHFSQj37Svqn67SscigKicnj7AInmB6arL/jY1ju/
lYF3BE2BMAzfZpVAKRzcdt2dZkfiq4/3YzLwEzgmJVwWjXuGie2Mcabah/90oxQ0
G8QW3IxBLl4gvy9X1aPm+tPRFghq3c25MMdRXarXj4NAIwRSvaE2zKacTGtONw1n
pX2vJgG/bXIGtj8jstKCELpBHYjLlrqr0ZhLWXBeDixI0jjR0nlKZENwTUmsjrHK
Sei+9k4Tfw3HTi8dF+a8EOpWEJTXmkMMhHobvRa2OyA4+fbY4H/MTUitTbE6c3zR
GLQjJ2+Ri52UTKPCcfyqlZCm5Ah0wcodFhsjO8xtPVO5XGjjc5Fw8+gWQOoeLAJz
x9WKtVSczMLDCkIBk++WzBHNXJ9qwLr0x34Dy8doTuG3XkDvgFSdXJsXGR48LOos
qgkgTRytj3cuVIlfRm12PKrxS+40rwfx4oFznUUsqdK3iwndlh/29OrFTM3bVIYy
SBR+sQqoQkTWoxZlB0cIJPTrL4CARlv5z7MRQq0u3YNjmzVhgaJZcf3YnQRsoK+b
v8OQnjfBH5gI9onugYEWGXKABvycKiBoZFMjM0BR9kz7Z9Q77H3u4nG0qiBZkAli
sW4MR67jLKnp70VJF3i8gvQcFyq1JCH0tomm/KbtKXeFgLqGDNic26164TUe1qvI
+ZqMPLxJS7tB/Zj7CX5jVNVdnlbr5K85oB52intEQ+gwPKz2xHcwO5Ct+B3j4fD0
dmSwvIsPKVnGELkPi4fz9GR6KKlUXsQQudk9SBDpTY38sI/xeK5ACa5RcgQT6cSO
KagpwH9cR+CTm00Jb+eDzfzLZTklTq+6JO7Ja3HwOOwDc6Fsnc/DIdOIGDGXPwAh
VHHjrnzopwymX3+BEJaeYheB9xfg57RS7lqqNNxEgl36gPsygZ9OGfNWMRXJNGu5
iihHnwW7j5RSG5Ll+vJDLZjGvQHq5HBNG2TTTkYS3jV0omJaKk5bVZ58uv/sVnjo
ZUzOqL7VcIEXTKaxbv4izhax/scbMh12rxqSeDW/zErISS4O/B5jjwkOxnsDD2CM
6Y22v7UGc7kq/fg5C082ktmlj3DJJG9/HxHNrwxMMnTwmheq4UpfojzQGMJyze5e
9JYYKUpVJbUdr6gKJI1MtMtFiRfV69FVFoqlGe3Rc4KJRj5FCxvNEumqCx9loigK
urPJ706J8JKfwZapJR0E5bDiKl/Fp81L66eqDtglQM96G1Y+4GXWG6PLBEtZGXyR
KLntWDI6ThF6Wb/vAlz54y7UdhFOiNReLsMzj44+tkovVRqP1P/NTXUu62uhrUfO
IeUChayI1NN/SjBMdkdrkUf2QOZ8zvZayCyRMm1hdZujHVPvQUBPXcmUFY9rHb/h
VXWpHELMOvXt98ofRg6VBQTpup/VZV+vx1MjV89d7rW359mqLUj61JYviAz5rb4Q
RLi5Cc9wPLXi5aB/Ct0pTQFuyr2gTR7X7TsHx7ktaeRqfJ3Gq9IpxdHGsHkMA1LL
HGPE03C4NQW7xfuV5eoZEHUZYJrXYIygAhNR+GNK/v+IuMK2AKoL8xAcTDa9uvt9
rbYVH25AB90/KsYtrRTWU2teLTYdYQogOHMHUTA0j4CLjwlQUoteTF8ONrc4qf4u
7oZ4nycy7BX1JRJHdy/bASohFDGVgpXVyCAX0rUw2ZXnn8SMoIZ10oF0GWCSS/zS
1x+rjGLbNz4mqr0ynGFzWcPFEDfIY+2oxvV66orBhlp9s8OlRxD+sgjGqiNG60kn
zyciA8xeT+WplzIcnxsMLf6Vt4BvbhcaWyd6vAFel/+qg7yqvVIwNDUK9jSSvabn
P3DPGtO0iO0MpKHLaZ5bFDpVsFxqTi2Z7yjMSSyqUum/nUGMwcAD5Q23Dmx6CKgp
pFmYiv+TumVqx7JJlnR8+tGSiSy8lgkKZc3+JnG9enil+eIdkl6ZC8JoAdyu2vwl
moVQMhSHg7L8dPf+bzzj+PZW9nrpzNsjH+nMRZyH04LSEMPqfXqiyO+i6+5ejb8x
2IHVlwkE5kYZRb7IG7xlxU1OIPPmUTPcVLuhQksyerVbsv4Q6yDQsPFJ31nfseZM
1wXhyGHXU7YH/GXZHvLT7r8+TsAFq2gTQG5ZC7OaKNs0Ny8+2OutnAFRo6raV9J/
Wb3SnqPbJvC6eseJqKNxXdEkTs+FSyP7tBYry2WUp+KylDUHgIFVHcqzD1dd5ooM
vrUDigZsDcBk6wlMbfEwVjduPtT+3MaQNnIS2CsfzGViNBvH12hczmYWo92C5FgO
EPQYzVd2p48uhJilFoMe696s7KM6wmvHlmcrG/dFYSmaB8kHFrdXJAKOPsSx9dm+
m9RxxeRjyFcpVgCQvYdOwQ0Gdoe6pj4l7I7mRAGp0tqX+Qt23TBHb4GfX7tXcN2B
67t2hUTSCQJVDU3s1bKIclBhOFSUMB//kbfcKFaV2RZ+CbxxAwkhkpi5/4pLV+Y+
YWZK/FNQu53aHCB31+YhT6IhcE2pIxa4r0AsAEFLBnVGzI3SGL4Ir8lxy6DxZ1bF
YM84WbgOVYmOLAwoWBQFFFutjFXZ7ueUafI+bnfPfC+ZkKr/IDObXFElPNNoiT9P
W82rRRHVIgiBzoVv/jYBb9Td/JeXE6CAduExsygI3wsWdHZMI7W8J1aIo6hadHC+
zk6PWfIc0YDkfUNJBFoqwlODBcZOizhjCLYBgWYwplEnktmtE/wpUYCrR2XZYLHq
T5JADsoPiZzrQh75fHF46Lbd2CE7zNdRblQZ0aK3QFuXfOnJXB2ilPdATKLtEh0Y
wJcpgSwAdJdXhsReNMHCZuj3eyXQjYl8RFPHgor4lUAOIau3PuDe8Wh6/erlJEmB
FxtpbSl8qlc0EP0jzVAQWZ+EYmqBGulDlgHm6XFYT8+WXeTI2XkLLJSfX/EtmuDC
J6nf8txSQ/uktDtUlsaxdlMZzje9PUrubH+ltSakjL3d7HC1PnBTL6T+7QcMgnOF
DiuEqg3/Yy5lk21PIo8AZvH4ykGeMV/S6DQR4QqiLbh8JlSTfQ6wVQQI7VIGNpnl
5HAV67YHTVt0KWT4j5ZTnBCOxmfYj/2fknJP7HEG/V9oW/XVoO8spGiiEGobPNri
eW+U592ypemw5f3L8rRdgl7veLerKyr32PeNIfJ6DROVwX5U8xEualVJkV22/Uv3
6HzqD8hZ07xnHg813Qt1G3QyTfrzZvllVet813JTiY3/lXzLG8cSPUNOKWfYnJOu
u8dSfmdDN0xIzFhYs0HyuFu2fcaXRpKMHOwAake8mWOxXbDAVQUn/2HkNey84Dk1
TbQRbWKDqnE82L/Jz8SYx2CSaqehfEEU4RU5962XFfq2jcCMR9V/Zl5vk/J3omjC
ZgXw//016ok8EA9XKqEvr0ki0ecQa2QExhWH7Xkh3AeolqywOnjynMXABYPe4yjG
W18L5zjZX5N3y4kLMgtT5YZ9FEPiFZc0Qk0vqscqENcVSb8J2S+7zE15CnVNUP2f
53YjLyI2INORn9bgHz2orwZbaPq2B5lSyY76taja1wjZYm6w4p3z/ROq2ajQsAc3
TQQ7CaHvJ0pXJmw4R+BQSpN2Pge+1BVYBiQJJfTQIDnoYbdsEdzUvYLww1NdO+Ml
AGI43suLY8FgD5Qea9g7QfORX3fZW2ov3XMWPusg+4SsWDEfGB7nKm5OyW+6c4SC
32l1BvXg9Qj2KV5rpVZuUedogcjUc18XMjX77rqt+Cs47zo7fPQwZ6AG207QYkFU
rH6r5GowwHfUGT54e3VuhuXsKACPum5yVUNNM3mKAQQ8juaK1VcxZEkzh5b11H7X
XSSlckcDBebe04IfwuoqBmnlK67n7+tPvLcS51bIn/GA7K/hdT5szWYLeLdLgvfC
Erj1707Fjnktv7azwSlx6yHxnau3rAdh2P6hg87beGdwiL1Smah2GTn+WlE61m5z
Pz5y7ysPqhOwzT5mMrvfSz5jQ62kFZr7hNCF3l6V1Mw9Y/YYu9dTIevcJtiah/qb
VagaDxRu9ROdvSGrYUPFM4pJRHv3t4bv3HK8NuzuJAGTsejyaa4Qm2ft8UAaGwfW
+y1hTSzTr4cbVioilNkTZmOQy2IKiepA5b3htiy3I78kFLQeqz/nDHSQVMuYC8Iw
mUvRc9FpKyDiJZlhxbTPfBlQ3EVpJOazOFc616XG1OXhauOwIqywqRbhWm5eEG3K
6+ttxxaO8rT++inqVfer/mwBozZIBAiefsTHEvyKovN/W71zZxuEuMe5xJrlB6ay
ndLzSwi7s2vZn983sdF4A0Aa1u79+CENY41Dkgvg0+XUZUOraEZxnOcgQTVvtZRr
H1uPCmnMkSdlhrs1RZ3DidKnGbXBvz1ilPudvZrCaR40Pl/aICQhAOTQFwqQ13mX
MEew4vvaQQYwOD54yhYb7DQipSUICP1T3vI5IzstglMzmrRjhsCWyN7/z8WnBU2r
yNI+Efzpx5nRDFySicnc72oqAxdiKpunLFALQ1KHQVR8XHG5M2uajeOgXl1dU9HM
ffVis8MA0mq8v+4O3tcGqoFq7rpQbFL2RB/U0kh0Qw9zCi1EXr2xdjyzQe7FBYMk
GJvLy1chNQ/6wiP2GLlwo4uz17vSyp3ZpobaS5YISQiNTU2g/aIZhex3y1mFDDNZ
fblyNoUtLtwm/Cot4XMMxlrmyR1c2yd9cQ1aGZFUc0mxlMGHZwZgcz4uN65W9neW
nGWDdt7iMPebWTuAQafGhTxpIo4NwJh6OGPEBRR/YQYpVcxG6hToxEOFe6gPNTl0
u8uC96xZ8Eev68MgIbBIYT1O6TjBXN03vXrChnrVUprzKkfkid6GlHvqDlCJ7j86
42WwjFbiQDWPrJCkWRKksfNeQfElJdicA+tYv+TZRBBKwbbqTqrSN8CixLXCEKpw
NFDZBzeXCm8pziEAxeM2GBegVvYn8FqhoNToDA+PrnO2cAJkpB4spRjakq+hBwXa
W0FqBQiIM21gvCbpoCtzAihoGFuuVKisMf1I8TRb9xiC/8qFlrKdLNROXvAraRbO
qG0H/7VH+H2nGW+IrR6hHc9A1yVCFbg0xopUEJzFewgRcftd31O90Y1t7dLLMeNu
4/YQ4W6pB5H+jkKV/h4ObpQL5Kpud9jp8JFUkl8XcjyIydI+yae3tcytyr3hLr2Y
q5X3GrEF+EkaCb0WbRRmhZKm+POfhjlHuhuEE4PyQczt+CEccF25AabbBxE1tnX+
y+aQFU4wqyqvghsDhnkwRv7H5JVQFGgqmIxjPSlM5zFPbAv3dfIGT0MhKmfNs5Qz
olUOF7jaLn+kYiPJjIgI1t0B2bQk9LPB16ESe1vHY7Y/ab55Dkxxb3SR7EdSQ5Nr
RNSqNogt4gBknuefP0V8XIC4HSxYUhFpObdE/yEEf4LdE+B9jL9qlzLjR6dqGPOJ
kHmc0ckjYyJj+QGRQElGBP0vmu8ul3gXgbIyNY3+50HfbtF/ao00lnv7JpS5zO9m
tk25zBujpOaqpaJ0VHVj2chnjz3NuMjv9sfAkfZ7Fmzs+mvQ/wfNmPRWwgKioJH1
YWw8ZG+NEmg9e0JTxXYtqXiTLtW0u1e1viZJu7JAcyP6DzwPt/e7BQkMTLvb2sj8
tN2kGlpPtdXrEf2tXIi+UGeFC5XOrlXTaB01xZ+1mVd2nqFhXO/7YW6Bd+604o/z
vhoVVFIaw5PzrT7Ms/77vJX7XFU/rCbOIvmOt7aaeg3GEcdPecipwhc9jENLIBUR
KvzvYNB5NRJeuRGLCwn/IpLrj33PoWPU8p79bA4yz7xbqoawq6oLNtFY+9+89ccp
DJla2va47tZLG+pK6UGbY4qkvFboNBPdc/GQHMxYe9ma6mhX5P8K0ZbwANH7b3YW
EC0X7NTsoz+aDX9mLo/qPRFNuS4cmpBe2HtwVFuZusbyCoylCxJSm+jRjqro42mg
WqKZlTwdbcZxH+jecG13QB19xd+i7gb3n8LUMgH6OJpzUzh04DE4hO3UYYJtYEbK
rohRPMBlS9MVZILw5X7Chr1IDGsqUD3MZwlXktNLRM7l+uHZaANARYoqgpBDUdoZ
p/gUfmXIpeAUUB7cYdgJQmmRZTGFp8n4WCxa2Tf3UH+QS/vHe3ONqJxuvGLxoeZE
07Ra7shjWMnCLmaF8DZ4BpUmiAE12QyqSm2+BKS/ke1Y3sTUzdo54rlh5OwjvfOe
D2tDnq4zRXNTRR/mind4sgJhguaE0kB8rtQFM+CTMyC+GJSDTPNAI4b8nX5ZKp2z
z4smHwvLueU7RDrU4aGPC5/re73ejUwxeDNAt1TZTOUpBJ3iTw2RG9u/rXaZF27+
npcb7P4z0Nd5orw9vD4ucCs/AjbjI6bzaCYT1yeQYydfQlyl/NygyB2Fwr7xTgvh
g4esw5Q6CDRZjmUPTxSgy9cw0aE6t5jxmzJsTW9+VgeHNlDEkKxz6wxVOyYfPH30
BGGqb+LEzS7V8cuQYJnQsfMVDz8WU9kJdm1sK1PLhNqlB++soD88t9DL63ifzVdF
TveKb+WNH6gqrIhS+hmTuoeOBq7LBiY/ustLqlgwFgHVh4EmsSgmHYSed4uIS7Az
NK5fv46+yCviP42XByBCqfjDEi8J3uaA4cS1ttGAxn5/7YxIFD0BKxZI397OlmKI
yKXzRfXDqumTRjnJLmPUE89cUQ6a6JR3RLyYO44RWlwBfGwPj/t26KaJ5o7KPcRX
BztuCYNCn2FMlCVmpyaLQY+2+x4ePhQM34VdgdkCr+EVioivRNXpgDpmf1EEW790
x/x6eWm9g1koUFztuu+OLfw0JS0tLDWCrnnKV/kKhOsMJx5ILtrneBfTo9LpWBE3
O6IR51YzVl+LM34KYqi4/YWMS47TWVvn0kVZ9mxGQgciUvCGaP/fRWe5UhY+m36x
rG17QmZ/4H1P1UZ8UVz+A5GpT9OnkRPlWDn+ts9wh0Rrm27mxjjoajKYh9g+Ttxf
0Sqe6hXxxqmSt/WmibKI35sNTosOrMabqHy+h+1A8AMrCUYFY61pvaUgDlI9K8hX
3tmjRyiu2FFvW4oy1ePaY/zSNZFqmNwC8W3QS6yhDlrNgMiLLjVYS57MbHuNcTT+
+pDge3dMOhCkaF5jiQIROAi6CrQRhlCVdiz2jgAY42wtE1bfpxkzlANmqXqNHoRh
nslL+9nreW/y/GzsBOWvILO5fXuxmWcNZvk1/vz3urWdSibAjUOXTPkoIM9i74sv
bV6W0SvPvVW3jsbFNP/q+hZygSd6ttby1WrNonn7nKfpUQDz5i1oH3GY/rJi9Sn7
Ry/oJLXvjuVFzb900businYdyZ/muMrneARNl+/L7tlOS1cakvvwCLYKkyAC8bTW
KH6Yws8yh+R2B0swoH05Q0AFlBr0z6j+ShMPPk5k9Qc+d/ejsq296Nt/dxAMzvnv
sfQMzNaWnFZDEZs9Odj4/FiHhyETCBpADC2qnVDqzSAD7Cq07jr7UJWMgwz8QCtO
X580FzVZV8YfzBxSPXrVECNVlfX+iymovNqbfm/fXyrWyETZvCItLw7sEx3jnjWt
KE5btN3Pt5xzSSxpNMScTAaAjxFkBxRhzKdCfnrgBUQYBoW8D4blmRc37ltXHbir
8bFR+F86nGKErjyzZBGS9cKrT/8col5l6Ed2hsZlJqaHpoRt3NXXGkL2F9V5BCli
Lrkyau3nNo/ibfDO4lhcRjp0A/TTWC+BqAohqbm9g1D0Fm8xePKszpHsReUSE7Eb
QsgTsh70sx9fx7YvlmtFZ7lyfP3o9JWazTccY8YVBDqUHZKkWTa/CApUN9BXCVlJ
cDFhM5gxCyHwDLW24LjpjEX3vZEpoBwTUOcp6ol39otiVUP7I2EobfCNesqpG6+B
mH3Koo99p+DTHE8Chdr8BPpHAtVUxMc7KUgAIU+1Cs8ri02JTUl2vOzOUJrWgWdf
wJRqPiDDSAr3wggOgqp+A/fcbmMUL6eIKGB0KHcVJpihcy9mirfMj/xwbgkcTfnB
CuxxPTPqeEN+fAFTEYHppZ4b4HRVcU0aWHYSHYv2zp4F2IcRK5fn7KsvU8opmLPQ
UAwtmdoWgrZ26Uwgi7x0OGkHbnkw2wmZ8tY+xsZzLzoEn7N0GNh5Hn+GGn8v0Onz
cWj0CmiqV1o62+iLnMOV02VCCmq7j1hg0Neve/YYoYRbnXBwGGqBNKZAf0MuCyTT
K6GeVvh8wnTAF5untjCvtqjI7pgeBqYpulqM89g7N/tZIujBQLx9SHMKoTboPxHO
JADtaW2ifgFfA/Iu2nUCAnHRYtOQXCQe/62J25zgiprpaMufI7SuRbtHh3mJYO+R
1Bomz3GIZXBbVw6R/ZcoeLja/DBlodOyntUQ2ZxgszLF1oIrzqmG3nImeFsvM+tL
WCoLSgRh+rhcaP5gHE6pAZpzDCERWJcgunwoN4/fdOhgthazGLlu3+8a8qwDE2Ua
+yNDbVH8XMyKdDTzZyKxBigGnusjK9vef0xboEzRbgk+1Tg9XrflKGaw/r2+Z12T
2dNDWHalnP8cz6xlHPJrMMBFmjqcbNcNvUCq5qMOhyUmXtTHqkkM0YBE0X+oUa1q
h3DWvgaDfjqv/WJmONgGu/ZmilicZ3PV76SemQk2FHEgxNGxEXMdn/uOEqLwuTHB
24vjhkfAlJsXTBcyQqNRK/4P8WpsHMCV8/iGGTrc7lJBi+Sj9IpUyCvc/H19G8HB
CaoSorLE3+SkBWdUfrWCQPGOpWzm76NLXnaJHuGJrt+b+3tMfi1JNntWoSSrBgqR
EfZ+lcseNZ5DKfngPrgElzHwDLIP6ZOTChAAJud+3/lTZM4nmRKQ506CILUwoGb2
103j4SbD8dNxceWSUBpkAqHeukseW6N245QLmk3MK/8CAIj7BvZPy5aLUL5n1GFg
+87cIp03Dout6otc7h2Y3+W/j80pDFJiZpnJWaCW2zs2mq/ZWP18Wzw/57MDA34G
vgyYCGx+5XQADHnEusT+P5O5Zm/zexYHXStMy3rijA8gUOpRV5POL05IEQwN7MIa
hvr7jy0tMpY/VYbsD/aDvf1qynLbEBjVQSXpP41VadVrg/eXHoUijXwXZKRF1NHI
vUwbxW93k3rEm9UzH129nXdO5x10kK9wWhEPBrTyNq947+51oIX4/gzhjZP39vDK
By6aqyCm/K+UdEoRuyRFGU3rli5asCoW1N5hBpMIVYmotnv0z90SKMMzM9S8Geqz
4YDK66rK8fLgyHL6ISVf2uYIDZl8lKt958yU20MFrENke4K1GvliClRGGXmvda45
wFAKZisPNIRxxI/COLo0nabJR9yut5gL/584UmGHzTcwr6Q3JRJuAH9dbvW2vX97
LiqHLqSvfv95pMH8wFs2yiswxBP3hy4foS+opMrmwSDMuYlfVXEVFCwrlCpSHaFF
MPcf+nvRlYmodDrwGNMxFTNtZQ4hTKswM7IcNm3t6aZQXnQG3Is2X6S10NRb11CF
/Rn6cZ0gvLypc7IvkU+7XDjDDPpFc0dW2Ds6g0ju0L7BmUvq475QZQLxpIhYb3fy
+3bhq9DBUb4bgV1clFcrSJHtirEjfauCSOCSu9pBGVI8m93yT4awCPiJA81zMEIh
wS82n/2trspdE2fByVZ5e+IjHm4At8pFJocoal7dLJnpA8cel4bSQsDX7BhGvpHK
DBreyVFGSEWakJA/AjWtmYD+BR1U3OTcViNkncTWRzpDTBhi88pBKqo2Ce4F2oNW
wmvYN3eIgaTvSL/GZRvKOEr664531M1mb5Tj9rBQwYQaKALt0wDwsRSFfHxr0jVv
vZNIYdF+PgGk3o+Qrb38Fegep2IxJu96cdvkT09haTycFyquEqgz7NCkXKMb03Cy
UISZNnyk21xDdAhXj/558pv8bki5oJ5CtKSvZc0CgzuWlQ8cVBSu0dBOBsC2PTD/
OxqsSeYNaiGA/P7IofzIyDLGuVIqvrKceQ9enEsGUiR4CHh0k4WXQXnfvlXR89sb
Q8ST58saI2kdaIJg5rjJQlWcP8e6XAetR0anUSm5S0IT5MLkWXVM6+8Fz/C1+ko6
iI6+g3BIh/+t9z+QwgVO6/ARpkGXBfEj52gvIpVIuBXHNrbYKv4JZKenF3kHNwN/
7GFkC/ClWz4a4oV5/+mawRJ+5b5SO6p+w2CipdgPLz0L6W0X9YWxTjR+uaUdK4S3
nCjZ5s2U4cx8GhI/wCE0gyNHH+qgVhwCqzrkLSRgFLsar5yt+74o8r4k5JF9yJfT
yrip+65c4xvqgJUKFUtqs4IRipDeKxdvUVfoaIFllpfDbzPwHMKy0k2lAspU/FTi
CWy9jh5ldXH8wRKfKpfgNz6el/0Ul9FhF00KYU/X4LNAMdbMTzn485GM5EQYGLsQ
VN5hG24peF1wB0P5R1Hp9FKOEPM2u3+lUO9nCbT13LA6Y60qkPJOdldnuRZAIKXu
e5PxqFblieG6l4U+hh2OqwxDKGOhBzkFv5xjo3pCIDgxqcZUBywErM+gBOrkaMGW
oNsp4nlbFgk/8UGpYn+4dGoeOI++18krLoFW3gh7TJWZGz34/57pzdvyl4J2KHNT
P2ms6FWHitAhFak7SsfsDcLvLIxJzh5T/pfHN9CZGz4WKnORJvoqRY+ZWgXBuAd8
IpzFZBZfkDBWZlSe67YYNxG/WpiDouc//Bp1UAKQFjRAU0vj4KNBMLIMoTG8SuVf
TaTm6kmFXVlG61H22UTfRqxOlYtF2lrkTofgfco9vMDLfgNR5lHN7QD7M96QvkQx
SZtjh70Gr6Fbe+dr2yY7XSa4tO2OhGDHYeDKbhqBwvfCwt+ziywwdmOwjKZJOPes
On/blA2miz4ioXDh34SYBriZN+ixTuMsV5ckImGvvRnmOpnjKJvMP4PrDHsQs4bJ
KMRxWyEugmkj6xv6H5mtjrTHlZxSldQGULeWk/nTYQ4aEKqh0aS9Z4/2+EUO+NI5
QyoCLGOQh8cwzVt6ygoRIntk1W373ZIHjeJ5jCaXBsvxR/xdJEbV2Q6B9ABTUJwd
9of/H1QifgJgCF3k9neIKX6KNGg6OlMnvDDWA8Nv/eVx1ENAW94CqYkVoLj8t0UA
jGjIbfoqMwaVhdBXSjEp31wz6XzJ1QGvasHEdcWkcsn5kDHv39uNv8220rGcrC0f
5xDc69lJ6Y5Kntdh3jnZ6atgSKuoEHi01aG7NCiYHncCtn0Hb9Kpe3SmSxVY1kpS
iyPekTGClCGnz42J5B1/WveVdH5AbvBv2qye36H9rsA3Imtjl1BUVRiHE7CKoYvm
wWqae70MK1cCkNAiCjUr9pxQe41buDduyRlQiHKtlVaSv4+fpVUQSSOGmZ3E2U+o
C5M2wuByz7RsIvZskRAPBr6paV2pVslNnyXtvRCi5EEgeyO3jCh5j+D5/e+zaMYA
NJHzBEw+gK+J8IZRGD84w4HeIyeAsYA19DLbUjQRPKPym/zXlYOwk82Lr9WhsXgW
2D8kIapG8kCHreB5Jzu4leKXDY+/BNHPzZnGvhVLxfws717qCfkejN6Zt+M7PL/t
GXQHv8SF9oJsEdD6HeV5c3QDZVgr7aJzp6s18too7cl8bTbDPR1/n7SZzm8j1YX6
whlFS9vGk5iYYNdIydEDPFXJ6c8cO76zWdVYJ2qomXB5WsLxYdc0FtIjm8O81UGW
Ta/xUx3Rjj0fibp/VcciHf33uIaQvVWuKnOcSE+aRZYyYlxmITvMMsHyOC3TMLo7
cVeHqNw8hTtgLKHMnxLKq4yETO5MMLU+4pfAjLQ+nXKP21R6M7f28pgvqHmx2Uiy
e722Rm1skzMlSJPtXCKcLoBuCPJiSb7bLJUodtgHGPTOz8LVg2gsstedsTi6vUcv
4qeqk2w8w5qoth+38iia/eUyI+FqtpcYSHyUEyLbw3o6cm3ccss/M9f1uYgT62uR
qYeo7gO7NZb5gtEfD+Rw2PGXenyU0rKhxi04t/4EQUZvRe3u9RAn0UTpnm3Wu0JL
C+fJxeLbAo3ipgYI1sr0uNPIp8+HjfVoiGqqga1ggD8OjGEc/TiM+Vmygnwj2vbW
TkedhnnazJTIcPBiGlxs4maSq1uWYy3oYbdb+vAChvYTjkJcIPQpIPTcYmTF79cq
7y0I8IeRCCSN5udM5xjreU+2BzCbv9lOeOam3hRV39Y7Nz2houIqUfl39klLBAAI
lFQjZ8Q6IsEb7Tj7UHTrjXuOt7KjSH7oB+5+mDh3QUxnnSI/u8MBad4AmKAGJA7K
A/hECyQzVA9zUxNbqRnMtxYIEDXHR/Fv5m4j9q7w5b09PK0n8nrYyPsx9jXxM9oS
snLtV9hE1NtWhqvyVHOnqR7wepjrCznVo7fRopZgTWGG53eqGuWMEvmspwyzjS1c
iCyrQ31qOUPWcX/HoA4mbWny+0u75/6Rz2QRCRP//n0E49n7hVawQ3bWrWfSbqNB
pG0ZCYy55i5bxyjyNPwjGTooNx4oG2GKSC6b5PNdA0kKX8JkIoSzmWIcvOfOHAbY
+waU7UwON0Pd9McSjufYvXl/N70BHkNbUzVMvR1fpRZw/xsYhB6AplaZWpUzbg38
1i3fK1oFH8iiwlD2CwF9CR45IQIyqXAE5yk1fXXYYLiT7u9YmlqrHlwZVdBY45Ly
USB9HWi0mkZVBH5vjjObEmpfF+uiw0E4kJMuPtu57oHhcB2M5miQLKQiJrghf3XP
/Y1t8zcTjUvRONyGuFRW/k6pbwgGkdpTC5KDES4Ryj92XCDSuxrLbZI5Ld98eZTE
7gTvNpkPjta5Cssy18altyNM/OK/Iv2i3PJUFJ0VzYQHA1ZUTe5a98lkxUnMfQFA
aLxV0E9s6XR4VHSABIfGoHt4UAboHn4/auHy1Q4t2Tv6grhtGRrSb2rYMrU7MeLn
n8olQUrg+btB5S5S7eJ4pSeaPJyU2D67hMkDWI8IyFNJ15wIEAOcV3TpACKQWz3U
ZDUpmr4yiUOod5pno1NkNvb5tGFNAIuqqE8ZnW0d2HqeG0S7XS+k3HHDzn4ia2QF
F0WS9d9Vr4TSZNJe/Z53HqmBZn+2aTiaEW5Blk28xuw5H6uXa3EKeXGlAUYYZtLa
HivqO4Irb1oCgoxBW6qucnu3nPY5fGLsR6J8mmQL6Qrdg0wfeKzzokV3cLiith8o
Hq1xBQjfpzb8tSrXtoR8cAK25K64bIEeaN8zbqk0e9Mls4dLKtHrYDFF5To4UKIu
+qxrqnorRFdaDonGRkBkmOQOy4HK/I4nNv4rcvNZfJyBBWEWF2mmjN6Q+GQbfNhQ
wlM/EV4dfxgdKrUSwpr1ZquPSTs/q0NqxPpZ+dcdmIaWvfzWnjv7jHBNKoYtMdur
osBNgopxQZp3MNx/Vucpjoyk0fetcJqarbMu9oO2TVLI62MaT/yYvJci1emY6zFx
NQxZov9qnG5LmMmGLNgbfo4OPAQDOPCuiF3nGpT3lvBWQF81Wvy0gaGCW96hNzxu
Aa746hmExvj29nWKjbGusWVSljA1N9F8x8m5bYHQSUkfAzuvALLGfINjrephynan
3T1R6IDQKOcwLAfJF5qA+VQZTbvCdDKT3Skya9HVOJ6qT3nm0uzEMxlctdWJtic0
MiAEQX0RWOJJjiuOCtBy74goYDf1PttoKK035emnS/wG6yKt1jqp2GF9BVe+5ENw
Zx6Y3D+UOQj9ttFvuQ9mlcYjE7iz7B/02HXErkNGn49aYTRZ+0LEAGgqgQmtAlE9
7p8i2rdRfLWx38wTOtoVKwHtfWhJK1WuPOLf7ezgqIEUsuFP3360RWoP59yT8a65
zNIs+I/x+Tj0dbC5P05ZjlMKZPFAvtKUtj7RPpCWwnvcG90FPjpohaN0XrKZnT1B
giMACrKb4OZTwReh058nXtcH9bBR4MtXvJg6RMXRW2nuRTfNRu8wA7SRnimnstsf
tY4Tp+tH8eFqdn88F4NOPfD6QEYjzwBqn0Vu3Cuz2/ZWc4a3NoglbSGLWFDdpjlw
m7St6DvkF020ZN6z6Juz5w35cje812XhVHJfOxH6EO1t3z5DjD3RZVBmIQMDwKbP
BI3RpzoxgiYWohBHLmssgS99/PuHZfC84Jk4XfKG9GED04HEQXM99PihrPdRi5Mp
cl5iA0km4iZQ6pvRF1zkpESMXkSON7qzcsbDiv1ApUcRopOx1wyfy2eoB3HDToVd
7Y7th2Lg2W7ZtFxNJKfnFUv2PmJZ8tNtXUhyFnUk9N57NmGqmHL2/uxdbepqM5A8
6hcoDfgyHt4HLf6MoAXQGFQQQ/yrmY3IlEGnZVJ2Qq1Z5E1MB8z2wYrtHtHrkLMu
9Nmw5KUDl31pC2rHqHw2hQesCstHlH8i/Ec6gj4lS5BI5XZ4Uh1RrOjHHWqHJ70M
istLmlP7QV+xSu4rrkBC/wHmUWBRguPWs0u2EMvbXfrjLFOJm09qodHy4SxgskTw
FkOjwOYHBeSbbGONE/rP2NrQuq5P9YycbfrkzNOgo5PM29QxEPOK8nQFgDCX6ksI
Q0QY7t0aHxcegNVPWm4HBV2msjxCr+R/nfJFk+ZPpIdUTs3pqcgtkV4/WxqknoX1
tg8tYL6ba/9Xb4HTwzX3vvfWN1gRiZJrrB8K6QHlOwoF8pfevoSYK9+zd80oR1MJ
1b5WB6AP+WZ3m3IJOEqx8kWYfcrJPZlptIV4+siHtQpDA6P9daSfuSnl9/WK+KYT
KnjhP/6wDSmJgBf6w1zWdg7cYC62mtYPXKeuNrtigUzL/gMv3EZfXfYexy/xxZqK
KvFe6EVuvyvWE7McYwPm0MR3/y6BUrcxEZKssWSDCdhxmVhi5vNAo63jtHuG/kDs
n8rsccuC728fib53Dk68oKYyZQf54FqdYafnRkV4wM46Z9EwZIHt6HNJ/nhT+z6p
BJzJhiCWIh6swYT6QKJqaRGjAi9Y6EmupVtsYPSYNZ5YHQ8IV0NbJE3DU81Rr1GY
qE/ZLKJpciBrZUbe1uv1eHC9DgYntoC8KU/rh2VYcmlWwjBMsoLhidEXfhw/U7l0
ZIka8iSpcwsmZ4V595FT3KOV/Yiu95sL+QvvrbfpYeyuB1IL4UnXCzC5Gq85nge2
F6TTVdgvlDpXxAfk3SOTW77MqtJlbZdzQn9jSAhi0tQrB0SL+knvUZ96CAMsvtzj
GTcjYZcCpRMMsUMSjRXfbpsAxCiBD248JXcO5EW4mikIVq4Nt1iCyjc+zUvu+r7i
wcyVBeb039yVf2FcEn9xyPVF4vi77uGYi0vLMBRhMf9c4Yl8Y4kvd+JRx5oXFHTn
aQKIbNmlmtP1YQhQu5z5ao0ylV5rgFl8FMhNTkW2vuMCus7j7pK6l82k0zJhbYYy
d2MpaYlTdIy+djXfQyg9uaDOMMWaykb23EeTfH8pmZd05lnLQmCgQSzmaZropwbZ
fdP6YTqL4rRzGzMoKierVQ+Ocr9+4SJw6NK3SXrc51HXlyD68J/52PbzB+pkuQqP
87iQNXqigSinbA9N3bvDrDOeY9jMWA9nLlAB1O7XyzfgGTiO6B2gjIAkDAlHy0Rf
RE+PK/aCffV7pc1kyj4kunyB428g/8Zo0F8nPbd4moXiF9nFuLk1RWErEkJIRSaF
pkvozV3vmMFqmT0fvb98qGQ1uMzn5g/f9SC7UJ+E+WU74ll1CI0X2ScSNAXFfKUN
dOG97C/bUZoWXCETNtbCNceMeJH/EL5gfxLQ4hcyOAlgM/m7jM0ZHGJ0bLYEo5yi
Jb8rv0R/UEu0TGlKzDAuBUPYSFKacTosjFMcgvukdmW/8SVeKdDOICyjosGekXNu
34z32ErHg4NEIvDXkQrbUEhDkRmoT0Z55E+M33U9FEAegxSrMefgbi9zCMR79cEi
SsvL6qPUBMnskyGBsVgRa9g/ZMzXbwZOVk97yBuHNL9GHgAOLQs/JQdgQ4yN7Uh1
Sm2rvICl4Mc+RekwZnkZG9SeXjm9/b0w2L9I+KE6dgiG9fvoZtewIv3B1dUitj1H
Hnu+w4MT5pPKlaWDDh0mu+Ise9FX588Neri2MTyVuoeJ9YrEgIiRGDhVaiHOf1JQ
NXwHWVGT5a2l0bgBj9qCFyOpsEdMhaGe+n9ErtvU4yH0tuj4nt5Cb3DsgMu0I4rm
i/+6T3+EP6JpsQh7vNZ0Kp1/HxO481HV/WkLQ781k7nu3AQ+qZLHunftqsVKDopm
fQ6/BnKH0+LMJtpJj+kw+4yH1bco+Rj3rvzHaM5rjA4hnls/+7hzlQiUc67XDfic
lNGWI+GpJqY//YMb+OUEnZLeqsDa5eMHVNiY1GeyfYBCeFVzAnYslRdxwl8ivzAn
wnIym1fJMmKqa6iIfh+mvCsfyvHM/qXRaGDYB7xJSuXL3JXNHJPuvJDCUz1BWuGg
okJnpzCZij6bd7eDVTgP0R479WlPoMcvqLWvuQK45YpbJYgCGehQLg0BTzosSVT8
J9fbRBwpjPi60Lp6QAb3uij55zYPT/vfq89jt6nFNBWnRy7OZf/p/y7MsuqpMaK9
jL+pRVTfKOz2O2MsLIQqjZWcRey+KWpSJNb1y5vmZQJ/MCh5TK9NfT/MguP7JKiP
qvr3kdS1YfAM3ogGktvx5uwK3q7qdbKu74yKwN//h67oxWPid/93NTtv1kDhUnD3
Y5X/Acixgm5N0Z86vkoKXHNtmJ/dzZV7gfhxWSNYA8Ma/8RMYjIGjbYuH3QwD3XI
MpB8hwPjtupIGWPw55q+FW5knjNNo3O6j/wfaB/YegpTqY4wRACWWcijDT3k2hXs
cPeYHf3v4DOhlmuE4cSBXCKsbO9+z36n5FJyyL75ROy2jmdqdPkMhLgkBweKXKfx
laRDJGvb/rGDkLkjASfTh4SpX3AEZZYt+3hrYDHZQXH5goe1X7lY1QNcBGxMrkLG
CL6vUrAjqjy2WLa2ClFFJu1bYDR1RK2H7lmRBlkqyrQBExG9iAUunt8/c5v1Nn4x
ljjJnN5pgXAvHJzupIebfgXyHYcFhZHLe0TyF3W/DhHPFAwC8WIu7mbzs3OzNaq0
QPLfkNGCdBwZf0kv34v2THiG0ybNbf9OxdHJQSVgkVAK3/hkizonFavvmOYPZS3Y
ozFi5QRwjj0QaYyCsE1hdv66aOXte0NeWV1rW3mTsQxslypycwfZVqE+TbeJyYIh
IySqahPfkvgAMpKxvEEgfSRawLdsBwYplep2sS2gfsjuRReBp4+2QGhLua9WkPjo
2ZR+Zf+Q3wSszoXCmioMUlajHyfxYYb5MuvCBDvBUepCUo342bUl4VNcgOgHgjBT
o1iTzQ/zZP+L/swK4q7M7npD/SrcsKk4nt1mJt672Tn1Qg4yj85vur/GoRl3nzk2
otKw43E9kirVKxgNIXDekHl/Do7httoMDKtl+YnbeYFIr/ro6koaLrP47hQ8ParD
1SJ7vXpxFRb/XjmCZ2cRIYlamwCwu+CCg9t5IpPt+cOCOEkQoeJnYbpk3fC2/ndZ
BRKmfDsUcDeDY3Ua14khr9e+UsCPc/O9xKGq21uPOZ3YMszTQBEMp43z+Bb1Sv7c
Ph7/vXCkmkzCwSfvsNBJgQfKvJd9BJfKtlubgsxtM3ysihuJAdFDWfj0cjxgloe5
Ek9tufoBokPOqbrts3aWkQ1uD/mugZhzSLe6bYy18xziCzDpzodGFn3W235Luvq4
pcTKCk89Z1K/1Wp/qZBOajfNmI1QbJctALYz1/WCocpC/DRnEcyTKxPjhHiwo5o4
+TgdLX18f+cB5IWssepe1E80CT4N+34/Dyj4P+pVyJQuHtoI0cM0+nVAaY9lw993
eN76lAdGi6r1otRi2C844Q0B0moQsMZMGIu/CBUKGMKRvTq8z6U7FMyQufRx2isJ
7JSC6/gbmLb/4HR1z08zG3zo6ocFNH+rWEMcdkOiQcV+7URuFHtzb4CyMkw7RmZG
ZA8PNTRZ9/OefOqYAs/2oLZrZB8Y9CvxUOu4D2yj2f0EzfyxKFabUYb+/iUCnz5e
ApkqufecF/voDGhngXg2Wy4EXKLZ+ocZXLlVWEcFSiwvJEIrTZymPFxcTt5Ccj4R
ZqQvv+YiOXHi5AkW69xWxRpcpYVmZG7XabERD6WaBJtpSxsw0lWkKZF22C13X3F2
vac+awuVFfxhm/Pid4Veg1xSjeE8DMV8FlTSAjjGNDvaECpm4pCQRT8Jv5wx1D+H
qds+SFOF7ZJDh8AJd8qTyXbq1FkngSU6nEX9gZqIJ9sPp5pMnbnC1wzKCjzx947N
fS8TnZrqB5yr9gTbel+ERGAjZJNKB6feUrTomA4FVtqDnRwSPpyhxjoJKh8zAKv4
ToNIpLAywCTs094R2CJBUe67MVlkjctAzkYaqTfLgZ5t6/w1YIFag1VIDQf9ZsUh
+27onWtJ/ggqgIzwC36kv0XFFGB3BQ1YF6HD8NjqJzk3vjnZq+qydB6fIimF8WAr
PNHE5fAVZrlB+pSSPivVCvChW6a2Cys8YmLIej6kQt/RU06Hz0H48B/4bYHYRDXO
PRpRXv4Wv+TXZBjHFTgPlh3vd0eGdI1xbZfVFkflHl+XaFRy4EJ7ggMl1eB5Te+m
IO/GGh1ltimQYAOTn/se7PCjz87O/2v+1QCIxfuLYzjdste1osSTI3X1YNx1Z1Pg
jGc92RJJ8fMCC6hSw3WTrsv/w+G1HSbzLovvv//mI3MnsrxlAROVvHUsDzw1BhRV
XiB2qR7+0OrljcWFSdi6kpA3+Qhce/nAnSOZ3qldKYX+s0dEJnAqhixVuVBrVFsl
2F2zErHSAShAtKFNv0MOyx3qroE+QqTDN4zypK2W7bKbyVET0bY0ECYyDGZ0ppcD
CXBw8vEETdldJlrOijLD7dkMdnulShhxT95/sJSxkvZptywfND7LRiwT3R6YyM0A
J8vNZPBji0sz9chIQkZEjkXdtPm9cT9D8YV9UxwmIXG+XJaDyE3Od6mXeNNukWSe
gTI+KcJARS6AtGPnn9EoQ4D9Sp3Jae9HFulv4frVr3GnET5gpbq5zrw51eJpAB6J
9g5GMVP4sj+dmnx8EX0nNRd45oZKGbEunqWt9vlaVVioFKHicMSwLFg8+ymNBcPU
d7slqBFfaiUUMhsMdWxGSbZqXa6BjS/RCw7r/Zw4nuxeZgsvVpasyrKQndFvL+yG
Sm7KIO6O35tgYgM3iNhetmNldTqFlHiA2jnbIQunfB8wCIrCc7RzPaSDDdWVkiau
Ja0K9hA2USSWTipjCXpSwRMVDSoEmfF1vrRtfLvHIpHPdah9GHKh68Q+jgIoBo3U
+uK4CqEx85kEYSK6wr70TPrO89oqgCJ2RIXuWBdlWW+yNnMrdk/clZGRbrCz9g+e
6kProS2yungFnwZF2/c0QlBaUs2udOYjAy4UOgfi/tBu5wN5jj+MUWIteJ2WvD80
Q2SoQ1rn64pxbx7/rtt3H72kjDEeBLuif8wQm56oBkv/MrC9mgVUevZP6ao04AC4
nUAPnEssILRzJcAqi/cB0MrGbuT5kXTgV72eho0myxX/dPvC0+bbnkX+GC7dzOiX
iQ8ikP/WzIzwyFP15n4L2i6zTiUQ5LSWfZrQlV7ZoUcbgOi6GCIU+4fmmQuMZXrX
B8ZQvlbZ5qtd1ln3AagySv/otIYA1NkONQh4+ZCODYp0AZXTHcFhOXYkdXSDHuxY
TMluYGI0kj5UU3FAudEGR3TcrYcY3Hjvp14VuztZmSFGL/GEXHetlxmAS19uP3r+
TC6cKUSDDxOTW/bZbl8BvzdyyBHBO0ZC7Joo97/VO8SDW3dbYq3YVnCDqked3Ekk
krnT3UU3SmfMBOGWInPuqNzNe6AmcT90y2gTY1mmRHaSa1+8vaP99bNYp8rOrILH
5FHKpEd+t+ApkgBO4QhD5wFHlQUXdzN3QL2UuCdwICHY+0JCaxB/9BHu7Ujwej6M
xkNWDuBIm+UC4BVJ3VEZgnxffs9W6G9oWSNt37HrucMmPZkpLty5NIBEAAzX9uBV
ahFuvox0d9d4t2iisy5UL2ErmTUJatcc5vDyeu68hKDHLKcLdKjeP1vPgxTy6ffq
MRN5s9qmEh183vYWh5/zf0M5AMVC+GgN3BtMeXU7WVrO5pvae/yZlieZ7BM+AwjQ
Xtui8QuHgBUUUpz1/zV9Luh7yYljg4vDWHoui5+QMLEnyH2wrfzoNNLevjoG0+K0
+dDa3DmOZ28Is7H89v27HU9RmJJrNvVBwMUdjO12JCIQaHHt9pn1thdGWGLUrulZ
QfOruK3Zl8NT3BNrDoqrUreb8tnm5yZtmdfTY4JcIRfUd8EuqJ8D39lYE4Bu+uvI
fG9U/GbwHRPjyNpup+ryzV6yvOd4UiucDyfx8HPtd3CTI19WgMbZX8p0DyS/lMP7
MdPEDwgACLveP0rPfTnT4bClpEkY3WJaWg4EX+MdOZIbfgYqJ/xD0G5aZE3TO6VM
9qlseR7kWJ5lGSsfAucoKPnai82NvydS++d3Jv7OxXTMcq8XKnsLfRpR33bKL6e+
1YvVPSFQjzW/4f6MBPYdsFM1ZMnF1X4lfWOrL34DuTDz/S5ZXk0pyuAkt4Y7Ptyj
TJRDY22D8cxZPYSq8hKF8fKpRuuhHLWjESgfU1vdfk0bqNtiUz5jeiOUcb27o+Wc
FBIebsJd3qGDh7Gc8L1YcU2OeN8FyEDh8xFQRP4xqQtZoLV1q/dNskFPufN588e1
8xcAAjwhjnyzw1xAs8/7pVuCGEw5EETuAzGhLatlUkjl83gQkgK7cShV1aK7lxAW
KFFY4lVD3hc6R8zNh0M+GtkQZg3Sl+EnLMzU0xTp/0yIESDNF9hMQaC+RBoHC/F9
yZ5+PdIF0QbFcwtszHVwGw0N7tRUczqtZ4qGR37rBW1Ocrvm7md5vujLoblJVKrs
YzUY4VG/IMLPbzOQBPhjWMToDsA6DQ4ERSLhlh20n3iNBuWNfDmuLY2W/5Cgb3jZ
y8XO9h15OJzwtJtPjHsE2e8caJ8DlQ9ECqTF6U0Tg20fY1PgAtDb5XaJJ3Wvl5gr
0oWe3WOwc/KIkIcqD41Bg2DBhnQjoSnUK/Y/POfLq6fPHr6JZ2o3WNyEpHwzPwMa
jeyuku1TrzW4EYybGXeeUhpOTObm69TAzWWkQMOihd2HZLmeHuGJCiJzPLUcj95d
a24Be2aDqwyGgLCKt2oJJMAqgNqW64fE141VCQ749KKUNlVqek/shu0bU6GWh2fX
40Sh9RGU38Z+bX0qFOKYYCQvqIggRe1BtOxhpkeB+lE30GZDuGmWmUCIGLpBbQ/Q
H77xLAeHWk8fnnuNT7lMGJZfMdOdVVj59dbnJXPhQzGIiNtqJDUZlyh7yJ9cC1e4
d/F2k/k5GhjRFPJ57hkU/hZ60NXKQbQIfr9S0UukxFLX8g6kD8uceD1cXWE2VBG8
eyzAvSne8FBSULyGxRPZRwcjmo+MnidSHOpau/hOCvYRhYZ1OrTin9vx4VIV/MBz
aJa9BdPbrc27wJDwRnY0TYVRVxj+sD+z3NEPrSNShwD6DAW3nb2Hx+mV6oGjSjcE
SAp62aX/JiA8seAYR6aORtIR8X7ujaVVr5ql6AdLw2aaYnRRl3vNvXnuRylF8rTW
OULUM6d7qDC+QxEEBvZqx18DMXexJR8kCEczcON48SNlj7LiiRI10HBqsggMfDFt
mSRH8lzFp4iG1NUyBoWiP+Zrl33jyTDMqSVmjKtIlJ0vqHjxMoA4ulQwvJgJz8Ca
fWvOPm6PLKp0NtHLLAdN6deUhk624O6BiLHOGkTbhwx3YXTaluF7jx+v8x6Vh9Md
l1rwPr+Av/orImbVbxX3coqkrQ6CArCfvN8tVVlsz3Ffib8/LunpZuXdbzrC2Rnw
N0rDmRDknHrzF4RpwVgR2RsfT81xmefy3cc3MGFtZ8R1IO+GGCJ9bpcDUhWugu/h
X3XJ/5ZwXR2tWubuQCzRAABWVIkJDHmAulTrijjEVYDxEFZ6vuzYx3yVJhsUNtDM
3r83wuRy2ta3BGfeOI40/tiB+jxDF2XgUc8AS500GnDZTJxIBaoKKJsfoUc0soJO
f1uY08TVzXCiMt2cYDVlWZtglcAfkCc6kh/4IfFNSBfpgck8LL4Ash8RUzPMTBzY
W7YMJLAmV+Cp5/aJn10PTwt9qYA5Tif27g9JP/9IzSGNFEm9WuN8p/HXLGgdxfsm
YpLoy51XMr4fFEuYGgK9AM0EcwEFIOCv3ZgoK/TUAZ6UcIe4kRN7Tk9lP1+kvhzj
77GaQOP6YCQP7ghAYJXdGm4aL7uvAtwkz8PLumAjU5jjulBlxCkEWFqjIl8hTS6j
iifKSi5XD8kqOIOe+NDJILy9uPkYWn/48iC17jPMroL58FEsjtlchcC5nwBF/KhQ
4mUUIV12pnFXghmM9h7CroxaZiUIopAO0Ilx7UtYWM9+qB5cyWe3Ys2vHM3Te/iX
iebgL58GohKGvHk29kwLmzacE3rMW8X6NE12cSnXtdnSRvPePBx7ouKpsN0GZzJt
ovfq0Zki4oq4Znn8bBs+FFRbHB29T3HnqYK7g8zXaiXwhWmL5FZk09bi5pcvMvsr
eVvvot2Aybs8E0A4UFl7O3oJSWlb9+IaIexEfpJWmSoYvrjkw211fsNa2d1yn2ss
dZABPcypTRVzXXcAS5rZGG0jwT+8vZ4O8k4GQDMDGW4ck78q8Q/ZfttINPbpKfXR
Is7kxTxqY8nEx2vfZoqD2mCJdi4xcHxclWR5EcB0tZl6kkqP60ozf8q3V0X6mCgi
kx3P+MYzfaEyHWMa3vWZLUKecW3yZsMuUqv6ISW4nNwYp3nRm+BRK3ZNN0qTJdsL
UjU+gn72RzuuPS/PIdR+O/goJly1A+PEN/qYgqhLgx/lRpWqP9iqJe7sXBjmlE7y
5K5PYWbTqb9Kmfwexy4U+4GqTb4wmqux8FaQkQ+GSoDFS/aEu2JVCzP8vjB3ou5E
BlDLKRAAgxhd/ruPMnnSdzzgQ66tNYYe1NNGUOn9i+WvPXTk7CwOr2aRGftZ+lGl
a9g2VyXKem9L4MqaG1arPfsTV1hskVB/py1YE7uTJ08bS6U/xS5Vu9Dy0KSbvpxA
VqAnNo/dIvY6B2htX9gwh8FhRduu8rFhr9aQQNmltgqXHk6LwQyYAJjLDVEPRJdh
vpaHuFQx+ynrvwwK74+/QC/uVjXnsP+/3WaFVqz2StTq3S8c0oDm0h2MuN4z3ZWU
GKq9bkW5GZ5ZkFoQhMurWfT7P7OvhBcyy/aTj1Gvr/KAMUkqqaGsx0sfHVhKpDbI
0E4jMlEyboByWgr1JKLNM2h/fznX87yJc+0sPrBGzhGW/Mj6jehWgQCXHRKuwKC8
FYslhTsqtJL1RlnrGp7FiRn4EIpdG8MtpnvY9Rwc52eOAj5jPlKVO6vwZh20l5Hp
S8Kaq2R5m6Irnl8YOLj6X96x1OQ6JmP1ZYKEralCYAHOsLWDVh6Bi0+gn9x9Ulwq
dJith6w26AusGWYChi0sfVuFzbXSkxdFk1jQ9CNqjkniAa8wXBP4Jc9tzowwn4DB
7m/edzMRy0VKpWQk33ycf98GalGb1Ne1Af7mVidgacKuV0J6jWzh0ihFZ4xaHjaq
koThQ2kBYfqfvGxNmTjKoNf2cPR9CJFw9t+tovk7HBg5nntAMVSSs+Es5DvtQj5F
DptaY1eQpLniIAQcN3baJlpO8RcSFefPhH6MLU++RQTsgYA1HO4esNtSms66SZ+4
918o5KltBY5U2uRWfOgkhLiuma4Ym0nzspN8rU7rXfGKnSXotwTE3B7li3lNskTe
dYACNax9k0o4spPt50Em8FWn9G1sc3q4N5FJhcRVkve6JzIYk1ksQALnt5MZvwds
tbG/DwFwNokrme9lqI4bFwW794tZuXR2tWlSrWXZpkqGZnyCgOSJcPzpvTYNL34U
nwB0c6OCEweSxi1sUmgHYVZchsAjf675ZBRGE8B+z8Qt2T5MELfZHpdqWwpdVee0
sZokYtYddJFegqdrAr+sJPVlHuYn3cIRqVRy9VpuNXO2ZGnrUI1eesKYjU/U+wX7
yQX5w1z/Df9mPRQzZx++6cITaJ767TADttVvTMKJI25VQK6F/rs7APnxRUK1xKQp
lUifCDaMhOwNrNTO9X5L2N6ZZXCNddOJsvfaMFAJW0MY5dMmzyZ5bzkoYPNIN3ZE
/bmc/Wft1JWWrGZQhStZyZIdTfJHSOSSKV7c0LJQa/EUgfeHKY5mGAcvrQWFg2AX
XjOYGl7cPuEXVj9ed0pkv+rjs697L+aLZcmbz74BVUYUsOi66azmXXHzzaqvEN0G
58G7la+VtM+CXd3j3YZG9hLxREX9p5T88ikIqE5JVrEYy1AZPqEPc855fw35A+No
rn0NFHzlh37ucr/WZpdZMX2JDuuQBzqoeEZXqulAD5woaS+65KdglI6Hybn7LkcN
6mBxpXYPPaCYzbQui/pyY6vR15TFrMsGRsa139HW/Uih+8PkuZrmiWpQoR7ZhSkE
YxUeOON6FgQNHZsn4M9oEF1/h0COfSV6Qv57lYb8nZEfUx7Vv4bh0WIN9jSVNouE
l2CfgQf1RYQYF2tBo0IGvO3ja+dwEnv7B4vISA+ympuPuNNp1/lx5LQr2D/kBUr4
iiZurJr/MIgxy2mQ9Oh/rsL/cuGT8MHDbuA4hB1JNf061Ng6w7ixzNWDN9yH/vjZ
c+owhd6svx9gDY5y3yO8CxFGk7LfhFI9b+hGl35/G7zqo6fx2NRIa20v3okrCDLK
+PjDJrUs5M2+dkCWYjmmj3TJr8btqzRVN8Vjb5hKbTe1vppnXuTiY+WgXUZSKhuJ
Q75wpBPuen8Sk5QZvKq1eFXOvRNnINi4/ubRAq/l/A/Fgge2lR/kVpLd/6HrLbez
QORy9xTGVFhs36PWKpTuGHjk+y7rj2yqxUrupwzXY5UPDBI9xgiK3jvglESBs2b8
4o6HrMeTA1o6VctX3hxhBcrvWQpWLBgiw+st7q6alrYRXRWEL1uGGXK2I9DxZI0z
pQzHC7K1vWRzTE5ZBFxKXNhGSXV3Fsd5QJjeokMMxy+TiaRBcs8frpVTg8qk6YYi
cK037MRahJ03R3cn3RrdeyweuvXbBbUekkz6RHL3hlHNOblHS2Q3g/WEn02kwwjE
e2ggLde7YBkb3mbSvWvQ5P53LTXAumbFycG+mYcUPdMg60LTur2YwIf4KVwsi4wb
JQp/60v/n6raGuQKW7+Ha1rQDrK+h5ifxNyto5PvRmZZaTM///6bB547vzV5XT/H
RMwVWnUk4rYOkns9URpVt9KZyIrsS+ohbKCGrgo1LlM3Qx7p12Beih0V9mWPfTK6
HVhy07rS786Zhpe2ap7BmhOZiA+NJHyYmhUAgMrZZmNcr9ozBh6qQ6DElkGmaNN6
job38Wh6Np9DLb++inQ0mjZEUqKdgaRrkjuxRegO370vnyVSdBaft+d8Y66wItWs
ilVwhn/uwkhjNrTgTbDzCmL9B/Q/oItiAYQMDyVQbP1KjIBQQLHU/mNBzypGRiMt
B8rCMZF3LWlIa9rSQDX+SHwejEylfFXCQ4wWtfVf2WMKd4gvz/9AZw4EX97eF20A
5uqMkPbpUP8eupihJYECFuO6NeEYzqu11gi6JtxNeQqwg2fGTg7zCIPuye81fMsc
tgkCi0+M19h0bdte46eK0ndbDykraA4l9kUEJHWlOTWaZwxCBpYv7nGVtHJcHSxd
49tZLnX3XIg+4RsYwPxO4Bnq8LUA2HH7MvYfufB8Z+wQeoBD3mIfTMdRum4y6Y5H
R7w9Esa2cUfHmw0ZbKv+gGLaXg/FnDZVDqB6NqkjKicWjPCks0vHPcxUGq2UpmH8
oTJbuY2YpOFXakxUWPzCf1asXcyrOwIWWRmuBJvoW00qcQh2UtMRmzmf65JBCpti
XfMIbn9Uo8jaP65PWqVsZhuXF1xUiN5XekWP42TdpOLvHeONaIxaIbM9wtAXrWmF
wuiM691edKZ760JWyElZtVrZS+6z/a47ScS3/g4XGrYPahxazYJNl0VYpL+Uxiw5
o8J6xqe6m+dlNkSQPl6BdiyH+DaCNDnLeFNduHDWZNMBXrLjV44UyniWn+SQ/BZE
9voRByaHaR+IoP5bIUi4L7lfN++rbxtQropIagg6NzXkg9LOp4eOvxKBcmJe/OMl
NTVe3MVbIEyyRjLHUCwgwg/GSNKqFb0N1XaTGV6newYipXWtuKzVhSbK8pG5f38k
yT7vSJpA7sVZn0GbhBrQm3UJCn6zsCKCUfbgaMXRKqKOFj3ByeveTd9jbwZmL5CB
ktkdGlbkw6P3A1KDaasnCDi+oXlA/7OI7ALM5WN3rsThJ5nSQ/dUbt63a+HZapMm
cZnCNNL5ceh4PJVq/er/f8oTlNNWMCgLQ9GuhRqLSf188Mx27Fu8THe01NXWY5Lv
0+fMfK7/ZpIJ4moub87cUd/XBq93BkYOMvE1LNqoJsDR55+U8dHu6mykVdipT8mm
cII1a/dsvI7W7qrNkLOi3DTODIa9eBnLc9MvVBFXxydtmT1nY9UST0oWzRd/8HHa
6LWcrJv/srM3Wtef/oxlvvReX345LeeLr2ReK6xUYHYRIl7LeIfOccMFS0XoX9Xz
4u60FvHoV50vtrY6JtClJgIL13sQgsfY0a333cruNHJUqn3XoRpkarMMD9HPZbwN
fpq4n6rT+S7HtlioQwHxylfEW8mC+9DL2114LQQvQ5iGuNxNpn9OYGPXuD//Nn3Y
pnPjupLHmRwHPGjcmJ4CcjMXz8q4u5JAel+5oaXcNmYy5+wdKpLwbR9I5FMn/ufy
gE9/aZvDLOnYp936w3uV84hzorLboUMzmuxQ/r6TrkbuwIK5EtheafpEuUjmlCWu
k3+zY7fqO3z4yPKPpRBLaw9jI3DOSOX/KoaWIkGNF1X+/S7hjZvSDHqPSxwPujl0
0XgAwnt17siYHYeJij+7YOnXD5yNj85lQlG0rqM5m+LQzdvecctVGwnBEsgqrHON
pcGqA3+RlD80NVlPiZ3nU3DTVfrszEYUyPkR1MUXrgq23LmYOiWI44vLHWGl1amF
lOH9SR/CcP3vME8NT4XrjPT5xP9nvGU0eMzWXDsIidDZwYYPTOd1Dl3ZczWO2zIr
mqvnR6BCQgq+Z3AINgY+lPpg0m6+WxIk2XSGIu2eUcBNKXtnyQhHWK8hh2KS6q6w
eGTppOMXwRZSn8kEIULyVhN7h6Bq0nzVKAWV4b5NfK7qwerzPDvpN+c6PO5XLvRA
O5LX//cEGdqdsXvemIg9idSnEVeItxv3GvvHFL/02IJvSNQKl+67JQ0W5A/Cb69y
PzdQO4MgJTQLbkhxmdA5RKWGxbzhbBQrBoyAqe+AAM93RBApBdfTwBjwAlcEQAea
M89uHbsNE8JjRynkpgybZo0XfrEBT2KxnnaVlIar/I9SwF6yuuaEpnhPyOuMLyET
9E/4DjdqLqXm9SyVMcveqdVjEcMo722UJ8GaxcDN5QAanXTeRVNc6KE8adMRMpXo
c/s6g07No2+uryF/kcf34scZEmwr0Ld51rPdF2MKJkpOXHXPnnq4HkMQ/zZAvydG
pHT+66cWmxzmOvnRuWYiMcNk3U9QmveCG1k6Q1cxrJ4F82z90BduYw2fH7ESEdc0
HxFdMwSYlKnGgY5I0JPjzDMcFZmNLG+GehlNb+5RwgLqVhZA2l8Hql7VTWQl8laW
VyQOVY2kHNF/qDHGn89IutgUI7HYUu5Cv5G4ljZasF1e/H3E0ApyLtpEBGnGPnlv
0emMHDDpYjBThFbF4B8k3K5IPoHTTbgLE2pcOSaIChUyH/jctUN0P/QbadM380df
zrnBEP9BpvA30HgBgn7bDxoztxeOX+5vj8Fh01BAwyDV8iDILK30nPngYkLkmzKl
j0ljLFxRzBkYr2UrxogW3FIR2r7r1LhfTSeJBEvzOdhyyjoKoR1+v3I5f9xlv5T5
HjPfIIBgZPPS2lZDOZeNcXpR2iDjQlxKejcRGv5FCfLS6k9NdPI3lvjREBGjQQyX
AOXpDnAbDX2cG7LbMCO1Mxth6AiPwqZY2ec8DYmV6U5yPKd96QAybdKaev8wsSfl
LBnvFXadAfULRe553oiNN3r+RyOBfkcvuDkmv0//zCenlHe9JOm3Fao9nlHs+Eag
u2nqwNLMgwn5LRIJtj8cjlzfjrtOlEDERrFnRwyGAtRxvxU+yzBm5y2XIMDST9dZ
vIKOt+PGdi7oPW0Jm4z5naPzP9wPLDtlM0zWj04e+PG0E3puUlEgzEs5zzFyjQPU
9RytU8ZUE/g86Ca55/YSvNetAR7ZicEd1OkjOwRinfmYfoF2nh/h+SEjtHeAeZTg
xgKCvC4SwF86QpnO7GTYN7ZKfnkB+Q3fI6gHHpQZKdzqb6f7Ai8MHKPxQNJkgBN+
qDCrWkTi4hqJA8whlq+VAjIVJOJVTpjzyWA5LEr95Cvx9YSb8dK9XaQ45J2vOayP
9Mg4/UAL+oVaDeB+o/fcVpwibgLaFStU/n9h4kzPoQGVEx46ysfm+uzMukaOM9b7
PPQ/cL07ghszgl7nI1pCDSfEayIMcF+uGKHkcIoGWmwBRlomukUyYoaapvaqG8j/
sb2Hv/FqzC5pH+FVIWWtCrf8etv+4COASkwV4Pblo3MnKAT3QmNn+uJsxVm/Bg+T
BUG8c9bhWT7ysO+xqD1xs9IZ5XKm0CJxt0LBCSK7RXgVAbKjErehiAZheT678Zc6
9NZPP/OmKgFF2pJWkJge7poWxgxdeOWOZWORtCJurRmKBhdTwIR4SYfMKpNP/HO9
Y85CjJirBQeNHYIb0cXjlExEIkhuvVzk5mAaBKtqk2J+Ac2s86TTCGuVqWBiDhd6
UTEatxXnWqK4LvTIQyHJ93E/yUNWYI7me+wTGpQcQxTk/B3gOQfdKDtxr7gK5Pfo
ncquy4F7CAcEsq07TFe6y4sks7XqBd1RsQ1+1VDFlHTUTqKGc+iNa0RilMaPwZAj
qNl8dxuyrCFN61DocwATpFhjcVe2Vn602V2tFiUS9bHWID0ylfPAwU+OGGUdVNjX
DcsBLg7xXQb8qbiY8JM9xEFf44HfKCBGxf3Y9698z0dR5FNuVbonsuc2/eJtR8QF
24RK/TME40cez10O0SW//tGgEpaU292p1/oRrDZf43iq9wXhyDcB1BmilPfVUfga
9WSqYyLtOSYoqRLqsD66zokr6vjTnp3+Yh9ulxdHttk4sH3IXrpG6LKeBbMESSw0
T0+LHSDe+3AMSwYZ++cAeMI4huRN/XbqMBPZ4sc6B+CKaGgLksHkoMI4qNMZf2yN
6Wd/KD9x+D7ALWfOeT17arW2xYHQ2/2V5AVLQDjFMdbT0nwY0UT/HwnxAH+oM95P
1Qi5J/YCmSPNLCap1LhNnxEAeIL0sevIqUJXOXuOlaqL+y2ucoVXHKHrAok7CdtA
WZmJ+/6McZSirNtGMUI3Z3vjTvxZGGtS8s06dqPohYvK+thdQWmJ0JeS2SImdYub
ndOzPAG4QPfoAOwdwT13FooqgIPFLG8X5xuoM7Q1NFS4MLDxUoy9XJXSfHmgEdNq
3Ga2dISUvp49ZbLGIqCj+sh/893dSUYgE7zCAdgA8H3KmPH/hbIscIbOevrWuw/1
suUMpldbcAm4m2qkwNIsMI2VF/jD4NxYKvUPY/37Z/vBe32XwKW00uXFs0q3D4qn
DpNLC4cHDAzv1sKF6tTkGyr7Qr6RDgFRYrME8wG/i/2JGHxr81O4zmGYxy4E3vhd
qJFsT2fhs2cy4kMCWuwnzZeIJ61Op+U71HVislGUzSdP4O1fwzXqywOlyC9i3Grd
5RYng6zN5mCzryqLHlY4wtZfoY+daalV6jF8D7FzFdWwOhj8+XJ04XcoVeZLLB4R
bmrWTuE/gzep2Z1ivsububpz2Ojwb/VAHHoB9amdQGiM7JceHGe5UAvPXgTnaXgd
2i+DRbtt2YhSgg0rHgqfFx4SOv0oHqkYBnxkZaXxw1LFFvMDkYI4VIJmiXTIY9Uy
Ed3Pfsd2h4VRcwGMI/wPaSEBTRG992aaduEjkd8NYeOesup/mOrB4ZOAiH6DLcd/
SipARijK+r0naIVuz3kZiwWLA22aNdu1dRdG6crJMcTVBnnCPsADijLsKsRyOKhY
7XNmJlDtCi2WpEztX112GYrMeLeFMxj3zZplIDVOvN1K2JHuG7KVYjR1lLTaZJGO
Iql9N/GIe/fQ6o+KIqsgl19oOnxl4uh+rbggMSJMozVDkq23L1Jte2+NJQ0YrmgA
OERNGYylyGaPpnLQc7gcFGs9YW5WXNpelMGGm7oF59OOj7XZnCYDSA38m5c4k+p5
b8Lj07pioaZD0EIjarValkwirnbzGjJRLLS5EIiivjP4mFpujSTXEA5iuzLoyFKS
JA4Fa015NMcsFVNud9wVLNY0LBSIeJjKi+AU6zveQpddfbIy5E/IBuFx/vqszuFe
9oBCgkLXG63w5hNm4669s2wyaxn5QKQ25pvJp3CR+ZjOdUJipxWDOpGDDFgF5Y6x
Q4EiH4bZg3Ris8/AparahXXeQWxEVcEfHt7t74UJwbVQWtr9qJhftBiQ3L8fc+eT
1CaQBQzU+caYioh0x+7CKWAhr/pF1oTIW8qAzSzLAJfBoeBlrqjf8CY3W7zFUJ2m
7WPcGpk9wdUJBePT1OcOdbqc4+8OBEtXjLEXD8VE6RNmigL+XcYRqT1h05QWVX8A
5Hz16oDqImUzw62wA2DP90jjKpXjClvjGaN452T42QqioZfqcdfHY06Sx4R82P/I
UpU0PHNKE0x9SCNEi14eLKMtO6MK0di95pjj735G05rBlf3iM9eukuiVnrszh1LN
o9HHl4IXr1t83EhicBRf2c2nrBCuMSNtJI9QSMVi2X5KR/LssGmyGW+YeLQFDzaD
3vwYAR/x5AXpLrSY0c+Ry3HBmi5LomQKKBSfl6jPGxt3lGGJm8Mp093tRf0v2y+Q
+QohGMIPHCr609qKSLEEb+IzarR7Wm0rrDNL6J4Rv9LdAgK8rb6OU3wMPyZ6yo9t
DxlfQxz+FDktU39ydCD1RsjKi7d8ius4g8GtS0/tnaQNqy6k0D7f9OasWzdPxcFe
cLMbJPretsAGGhDp1t3Apdwmz2hc6KrzUrjN50e4EIA339bAaLSsYQqmxog4oEt9
rBTRVyLyEnlzi9/F98idJa1WrbVFHPZGSZKpKEOmgLRmzAhLsb1iseu7qUSHKiKo
ejYHLulPy6snF9duCFzNHLudadnNivligvPb/RE2lnMt8AyvbnkBKHLPh6/dEozG
tqfI+bJWsLufMSr6fnZK6+h1SouUJoBXaE4jwnSmY5ybzwViIGA76sWmqyy/jTpI
SuMH4Trm0j8AuA8mtv4UZY6M7DlltGvfYY5S5i5fPEKbQ/DLXYVHYB62h+0vjLui
XFdpZEoYh+7YTdBUzCLBBy/jae0YcDS7MS829mOFRYnbNvvNtUrwqxB7M0bNV0Ek
l8Bb8AJ5XgUf9hYtyYNRc//NPdOpjJ9gQ2NtOuitCBaZUR5/mRya/nAWvIBxQ3uO
4MM6tc01gIP4q5u4iZwNdl04lZWICnXtZsDW7PaYFBxLMyaIM8JHnqpfdZ7jq0iG
6Wl3C9O+8c6h0In54e75YihWybuQh+oQQ4lb+HfLFqXFpAmfaDeusp++ri02Vm72
nOJuXRCfHiMYeKkWk98bUNEdHZudghkZbwyMAxHCtFazYfyr29Y85EYavJoHPCqy
kimt5ekB9n5kGYu4Cqc4IUc4enXIbXHpwAbiHS00AMKou9lqqyyEs1iR/pUcZaDO
tzC4P9vE8NdcfYlegfelwyRzP3VqiCNIYJztQTDGJ00HbJ+js6ZdhFourpwjZV0O
TbkOztW0wNuqEPb+9UgoTrzt+KywNWerIztNBvM84Ob/J19QUk/BN5qXWW+qyrTy
UYnm7gNMwtQEh50Kw2RyF9Vf+Ev8VCcQAEb/N37SNRTm5uj25drn6bSMndzSxEM1
sy7eb3M9QonHlgeMZs6xIfz3L1zzvOQkCK1uLuFc39cB6GvPsyW+7w/Nt8VKyDWW
/fE1V143AeIkZ+jMldjGlegv6le5YbNoMfRxg76pJUm5uLv6M0+9XozKBC4Hjwxv
04LanV/Jj2pOkoT0d/8xa+G9TZoE1KTxkHAgH8JoBd/xf+2zYYcRbPYN0zXOrWk6
dd8BekgVm4OveE5FMp71CoX0X4Zon1w8RmF/gcmfhMTxUCwLY64H7X2Vgx8O6rQE
Eou/MSaZG9Zabm1XOwW8GXZUbt2Xkz/lTztykZjIXWGBa/1FM65ifCN6jtiQX5W4
RlffnaO+mhXH845apIn3TaBEgQVY23leUx+bdmHS12yiLmoq+keA/DdYX62LLDSl
VRK/I9SwFFitPp3aVkgYAJmFknD+VxvY4LFtrBLLfgtZ+mX4BYdxXrn6PCHFb8FV
I/xdZ4c45KdxuDi2at0mcng/WT22qDe0jKVFJ9oQr8hnehb/RHmI5RcehjK7Vn+G
Ku9b2VERSgxYapnH4RbbkxpHV6iMR28QBmRfucZc0fpOJBlG3189lNrCCjZHo+L/
odvexr0UmtZ7d7SD98jD9a7Oeb/7+wxzxJalKlLuLxLFqu7dPagsVjxcBSWXotyU
wi0H6xgvjx7borLUg7XCp62iEOlu9YvyeFsJiRJhazt+rItRdL87+BtggWCCf1EX
APwDVFdWA9q+SDuv6r/MtJUSqmK0WpjlJdPbvj/LhPPe90ZYN1EgSZruwkOiPMCo
uBVeBYbqJF6Gf4R1FxAMctMIzpj1Sra20yo/+4wxWo1wAkqP72XjFz6mJcoT7JTK
LgTbDDD6QQHljy6rDR+8cNmFIVE3UZZ4M9SxZdOQsgCg1HcEDQZYHrg4Ze2ET9rq
tXSRyeQa/fZG2XLgrJEO8F70G38ICMQpYrmieKsD5kjaDWFtYcz+4GXrCj2ljugS
tMiCryRroWd8Sv/1/83cZLObiQKKgpBqdPLlKRDYgPeQQnzlNqvoyC24mWDCs42f
pvO+A/jWD/uG+oXM1/mCZHpvXsjmyb3eQnlQRGDlDprGlwpYacshQnfiKKKueywL
l/apJHRGIjrOZfAfWj3U7fXeYUFZk3H3kxoPqz2D8JpAK9vlEkMGPwvFQXX5EDsJ
MP+KjFzU0oSqvF337MI8/2jn8/0Xf68hLdjUo/IHQlLAo7u3CbEcMeNvnwsUPvI9
UGV2wmFEqi2DEHcQJPViVSCOZMW++HIClX51lBV19e4A8VWkCT/IQMuhrikntXlZ
4UUOh0idNIoGGevbm9wn3IwUpXcdUvji2UabrUnlIgZCMExm47B454bT8pTkY35J
YGRe8DrewqD9e5jYLF5almekra0mBohavbYYAweWFbj9nLkeuTf061stp7T1RabS
ceDIyDwYkS7H06MCtD6EMr09OMEfD4bOVhl4XzhKt78AQmdK25/t3DAJyy9ijSyk
mSMkFGxQzIuqwUalReTMwx30fLdJn41N1WYIdeio2EHN13TPpJFmCaKxMWY6WFyo
ZlUTw6UTO7zWZtK8c3YSpu8k4vrUpxDTXnM6Ipvqu2uoyYJipztKziyqYLZDOv2H
PUsA2W3KPe3qUVm46+bSeSumjvyWJyXnHVVvUdUx6C+o/oniW7sSqEwwz7pScRKu
SOXeh9102hwN2xkBNO16X4/in5/u5qfP6cqN1udjOskXw/h8DXD3wPii25lCgtNf
oM192RvL8khAqXHrp/U0G8qslGeqLpEBU4PVzx0IqabvM1YksdiOKndGrDN4vV2s
+RBT8AzmAwt5qmZil7m/Sw+cmT0mxebbGYN2Ejxfe0beVSo1n5ud3tE7jb/glMDW
XlQsl2uGomFDdyMTGYWdQ2uWZuydpT6O8ERR3lKWGClpm27A/fg5+5crgfYwX8Dw
Vfu+MV7EMHqqtpM/E7ZdE9uJkGFbau6ndtfEdV8icH6GjaAZc0DX5ZQO7XO7tPVy
6fmj6ZYG2Pyqx8c3+zCUfASxhSE8V1RiKrbljq74XILpHi7OpiO4IJiQ2VpO2uWa
a0CpeVkzLZfek2nghDUIDJJG67vbDYVO2YIY47Chbd2Cf5LPJNEy11BY95uYOiAO
WDvSN89vJDqXAlxoe9tEn1D1k+tvFqEZ5VBlmvEs30BFf/te9g8wMVSva5DceGe0
8XbtSZ52evhJEHhGGt8SlCRMok3YuQQ/s2Ov7G3+gl5F9jtjtRM0H1mai8drE83y
lqEys+E4UAamgm2PZPOsWpnhiZQiORK48ohcEVOZIffcQTsXrDbf3QHe9XJbMzCc
I9TYFq4JSPpRXz6csnWQyPOfmeXsW4MgbB0tpqel1XQZQm0eCw5cWiNMTzS3OTcL
F/2YFwx/v/SBpMokjJ0DQPUAp4Y+0r4wLBrerySmKvFoH6hQ+ZWfmJaMayjHaxj4
44p1k8ffBic7qskj4zxe/WjjNBpsDVIjh7iaJn6UgzlqlaCFo/AvJuL9I79rBslx
HZI7075D+sW4Cy11aUARzOnu2Wuee0MajfjUfuCQZdsGCcCLCjOpItT8toQjD/sV
wL74WrQ/FMHGgduGFdG2lL5vd0K61mRTlYHgh3wK0eYBecUH0Cd1COwvkJNK675q
sCMITBXuuNpBtkpAlW+O0LxoO9BOf9Fa1tUYmHXP/CfBQqmo+2nHJuNHGx1VyinU
ONdVwB7qJaW0laU0+s6qkNEV5GrKkwQcMFYwXNwEYxNCqOIyIEd9H7QgYG4WClJ2
Uc5chZNk3GrRrgue1kxplKITXlMHiUIobBIKlfC3lrQ8tYfSousnDZPfGvJm7qps
13PgGpvrPXZeqyzg0Nyjj2zFDk5eFohRyRkKxV1stm2rSNK2zz3cw0GaCrZM0tBq
s56dpqqKJOWquhj9Eg2g40KEF0tZMBzkvLcu6aXA1+l9CaHg3fQl0F0iiEykGGL6
HIVHrf1xN6j9iqjYYdJRetP4GHDA6Xwxth9+hm+VwH/2W7izLFKRIbgb2cEOFrhM
UQy53u6lUgOilRXFk6TrL3d5ipsn9j2TE8F6ZJflSo+X4KxQLpIzd3w2Vunyz8DH
K6/IE61g2NcBJyRRpnCGm9EFWhT6YE9Dx6GTuvKAkZX2NFcnRJxm+jP5qyQCpRyU
FMjQ01XzlsuJufwUAOR0TqWEsGTOHwcyDRZxxiVlqCxHesoxCHDbQ+9lZbBtK2Hf
qrkcmHBT5czMLbkRX0WFZc/EvuVwQYlnk6pEsdIlTQQb3Vjq18gHZgi4Ge4BoHfA
vYbLZdNzHS4rhgohf7UYxU5AsOnlQL/Kodc6AVqZXkSwPx6mF30pigNHPmcUIOdD
n59NvtNu/nR49u1EP81WDOnTr6q0WgQAuxK3Z8Z/DQh3g22hAdo9qPnrMkWwdeYo
DSUmpM4RyNOzCR5qvGTkSIcM+lUrM+8oafSXW1lXdj3oPG3HmLGTqvyDoG4UbNd/
GZPU1FjmsAFyfymYaVP/UDchuh2fgmVyLGIuVeAnqQibaen6hVOVtrM8C+z5Pkvz
gkOts0vuPQaorOgbKhVpjPVxMGCGZs3Y4kXbqUnw84F5BLPDZJBr26buqhtC9A4a
0fd0+ekVI1gdPgg6yxBz1Zmlxfqt1gvvkjEkvDZqxoUtu7s6xgKvFocXu1SjOJFP
NpWtR8aAx9aAmv5wJrhIU2mTBAcs0fyeYVy0Ipdj2PZlcfrpaqZUBsVmh6HoHKk0
vctqFUbpqE0GQWueGU3TibEoCXiYJhukqXbqmxRm+TT2VOB73JtwOVJj6Ov9WLxM
tv+RqUwRtJpjkIYjeOIzxN6I0zieXwVugN9Wb/d5CPeXT6wJUE0M9yAruBFxwaiv
bBk5iLg6rQTIyghg6SIw/MBt3/foqs6yQynnLOKnw/d4E7ImMokeUA4U7lxM+IVy
weY2ubIGxHPPhLlTVfgLea+ZPToTo1fDDblAehvqKBmeayfN2Cjg9mX4v/IhLWN+
rj5LB/+Um1bL4QXjgo6EhJBqXhwaNCWVEo/DpGuUZxWYw+l9ND6J3zMMN2Iwd1xs
fIO+uzPXE+v0rWDQKd0tnIvIA1R16uzLHD7eP8sjolEfb6g7XL5UjoagERi1ZOhu
cIo+69GowZgnxTA9u9RgiG9BIDPH86pfxDspDrth34eIV6uh3oZznb37RaCsu+Bo
HphDXlfhtZxsjn1k8dKL6lL3+ISQe3XVCfS5R0rhZFffr/xc0VzPJ1uZs5DrHzXY
pyn3LT24E0wT5pwJ05cP1aEJ8ufE94FGA2BQjjQvDnfrVz3HwTfiyVYjLwUi5P66
lnxwHtKQa1vCpa8wUkws/5blE/CFzOa3/m63V39E7b+qoxzgvjZUODXieiavseUM
mshRHAF4w1P339Wva7vbPz+5i/+dTjqFTRpFU2x83EGEjsi1UelIzFKyxqkNnAbG
W3wS1wtkW9KguJkKv7q+x52hZsJ6evqZFmuOAGYU/nfxU/hFVLV7Do+KVVrKSp1Q
0WiDt7B0xOls6nCdBZZENO5Iw9iu+cLe8GbFsiHrCURVMDQ8i89qquXtd5Ar+NpY
OJxwp9voEcRsxSWtTcAi5AYRhCyvHCy72efl9wBNQwR0XtfVu2Ka813LDx/DI+OK
L/74KCNKl3YsubUKgckj4PDpY4o+5LaMubwRguqzG9V85Vu26r4KsnugjVdfSD+Z
DGp7x+ncC+vy9Qa03Opa7b1C3I+1Kby/ZMEL/9morrKSU8fbZkxF+gVccNzqV5Ry
oUCse2DPRoHXu5L9lZQz8hGnz+ZunUu77fe7KPsG4SH8eDqcHB2C4jLF4uhmdVTz
wXvxKoEksz3WeorANwp9GNNnM4Mc+Bx5lW2dveXZgv+Mn/rN0hpWpOo9xgP1KRkZ
M+Fc8IO7/t3SoP5FFPjycwGLevWVUSvY6JTqhfcbff3zqmVJqxIrjXN6cl0xiMnO
OPtsYkAXmuaI7LoROhV3Fo6tTTfmEq+noMWoUc4ie5I+lZUjRMENiG72D+/VRuMH
oXObSrE/JI0Sj4tp460fPlVVmEEiYMsbFZiSHiqTOXmKqoJ2+yVptSKajy24iKmr
c9MR4lHgF8J9p+SnAxEA9afMffzEvA7UovLNKquEbdQX0L8J0zMUeS2FD+zd/kKb
S1BGO83y9hLbq5LwCDqkA6ygiP11ffN32D1BIlgPGh5qC/t+R2+XykIsJQlB1XeX
o6Mbd3OtXx1t9t6ufBd7bHm2I9A7EwljWG1XOUSXXQdtYtOfBFeGnl3sm7Re9jp1
PdjUR0EghPHrOBU/5oKDh2TKhgacY/nxghXYIEWYkT/VhAGyT/UagB9DUwb7y1Bo
oWo8OQI36M21xLrIrXR79B1gd6kq+Smm6euWEKI9U8K5B9K+vvL11edaPbDCdmB0
PuXppGXo6DH/XtVyDJP9RCVGH1PFQevi3Be5RNSLdUsMTPPzX4tAm8/SRPQ8oOjY
hKz9qcps6uQAcsgFhPQ9bUCT9zr/PYXedsjppHpk2fHLzYCWE4E4sm5pYu0HE4Xd
UpSltcsWFbtMzZ5WKt76tWNTSmg2i3rRbMg2Kbak7BGJYWIKGIsD+sK4tDngXNCJ
oAr3tWnsHMCuh2XuOOB2tHlLeAGt6zsdNV7SNwRAbtIlqsOl6YjCv9Z/vae5EYEs
+fOX36W6mPyb0R0vUzK2ht5Accw+hqZFLKB6DVzQBMZTukmu+ZQu7ek0kmQI0Dpb
01hJKX+dw59zsf9fXislHSK5HkresHyDV7pD0C5U2CTPdquECOVqlPLgVwX7Rtrk
YZKA8JeKu/aKv9VrmB9/3NXQuJYmHYdrLgIclcyyGlVxB2VWN94oC4csr0BMdsMn
vKFBFk2t1kDYEmNw7cpDrQuNk7+7+xiNhpbNtJY73eGk4WkNghANn7z8KlShHJka
6BZ6134xUSrw57EIbCiQwHn+Wflx7IH5PcSkbjF/UNxvVZbIIqqr2VOwXvr1gBrL
HLFl/DfeU/9byaLbGs8VF22u7t7ecE+IwbXZgL54cAIRwmDgr848v5Ta1gjuA0MF
hMGQEnR0QKkNLQMQtysgVUtuWWYIDDiMGTSczYHGDflJ7d/KfiFMLkjTMpRNOZ15
jg5t/of/xBlwhkiO+q49MFgPODgWjPlarN5XG2J2uaUtb2R8gm2dGeu8NPx41IYm
Px0j2z3uZeRyX7AOwU+WrDQAwVndjSsvQnfMX+HU1LFHhXubuEraKaA1xLB+sROx
mF9SCiltrYLMAC6Vb7oUsZ/8x1gKIe+MpcGdf/155IxNf+u29vDK+9LSChe9M9Xi
nBa7TjVj49NbsEXZIqINUIIUDZPBTbJ5u4JsxTjWcXbxeKUo1apqQrwzl6r83jY1
5jRLODjQq6xQLWiI/WY1/9fzDTBJGNH3qyrR/7hl+VoSsjMn/v38lAEEbp4oY63D
e8PDrEcTDoCnjWtl0+KXKu7MEVBvilHCIGf6feHMdQSspzHtzUu/WlY9mZNTzNNX
WV8VBGS5WAeC6vxrID+hD6nGAmUgfASki8gAYVXp8nvA1A/+OTBhpdc/O5CI7qhL
m+TkfIZDi0FnxXVloVrlh3/pT5ePeUQNfL2nQuRRcKIgBoP2FxlIzuT+rYzuPNOV
VMnCGK4/VBPluOegIh/FRwGTvkLG5jEFDlEqVMGCbTjNQ12KcF1HMDICV53pg0Im
bmqEfrPZcKj6HAuxuK9bqNgRXjqhX0bLsq7VT6FRyfb4m71qjLaK3ulQWf4aWKzx
8PZAQXOwKMcqDNGHJ/lXMT4YH4jc0CQE3jQ09YrJl7KKKt9XSiuJohPWTitAQc9a
4FRtc0tFRWN4/8pN7M/6H9REPcl4mZaQtkTejQOzGUjllcNjynjM7fpLhLmjh2uG
ad9OClcrx236oUZ4ToPLLOsHvBF6Vmmvm+P+9+s/Zi7sBBG7deQUFuwhR4+awkFS
WuLxtspwaUWfoxqNZKb9oZTeBfe4WihidyLH3IVfvhIi2pMiQpRb8M/EFXPtNQzC
OPCryeoTSLVFBKRO+tg5z0DKXY/mjUM99GNQAn7xgy19nQ1BO2PvzLa0zP7P+6AF
H5sX8Qzy0SHH3a2a+CjWYtI4zzz6y7Fr3PxfW7Bch1565dlfaxoyRswv8jbALX+4
sAiLg9eS2sV9LrfEZlHJFGtNGpP2bZRaNE4OCs82455Nj9FNJSBRfeEh5LIZ9quU
wEk5NMPy+QJmoHydHf4a1YRfm6uHubjSr6CcylUZ/tUhYk0gKoJ3aCo88MvuFiHT
bC5intDgCUrV3t3QwRfngm/4iuDUAdT9kTQB61+YKjBW5sY2eTWJCw+/yB4Ch+EE
XBeqJ6Uknc+iPgtxK4gzYHHYFhgPc/Jcw8Jo0hwjubYY7B1FdmzgVro8OjXR/cW1
fxxidCG33ze7WPEXong/w3ajV3C6vJ8Y+mMBBsq8WgVHAgXfvcNaomqOe+eCRVjF
60DxVv+FHvXZWpwq6vYQoEfSBbStOpDjbOGSFUI08ZZkx3YeDLzgONKkqCjnN8Qx
ETTQ6p2WQamDhaYY7hKWxvWY2idW6yBHNxJZ8m7uheGnVdc/2EotccQJo11c5Ya5
+7YQt9/2AFmuL9pf9EX7wYgEv87ZSmof36yyR+SMu0oe66LHwW8I7y7uKywB0Cya
+JzY++rxhGpmQRjaZn9CimJ9X/O0fbVo09D+ZJKMmS6dJIWU/Vlnfc4zOYI7tSBV
JHMnVzG/KXgVbWx7kSrUuCKbE1NZcwz2cEd9Rkqsd6BVvyS+/UH6nuNVQ9v5dxlZ
N3eksldvoEIRM3p+wKcFvSCIawFHn/jve7BNBzg8p5FwnxMmYzPJNSQN7OdLnr9B
RPv3EimsduBuv4OijRS329kC868zW4/5psMF0E59+vMunkB9PLK2QMBlDYeX8Y+d
FhWOSldWnNWT72Vlunhl6/icQxnUHNe7W7EDutztfmaoqsKiQtnzFvq6RMFu8Ihr
c90oGIOuwiIGiRkQdQ/f3nb8+NKI74H69RURgWPQDBZir2C+Z7lybLZQ80r06Y0j
pEtyym56ykBpJQLnf8LD4r6UHUpfxGnpLelIjpxdLyoDOwDyi1LIGCMeneyvA3V8
8FUTCs8xc30S6fxFXfKRHcPU1VLNn+0Tz23CbKUouFqHsEnZJkz65BDACyME2rVW
3ok+gqBdY5XzdIV7J2F35Pke18L8T4boR26bUTPY76z4WYKWGRL6b5cr6SEMRMK9
SmNqGHrOFUkOrYlDq7SVcCgfwP+0w1F3AM7L6XTOGy7tBTo9c5XyKc3gOn/0+uMB
udU9DRUle1O8S5zI4TcqUANjz9sxNHAmQktk8JQcFYmT3QqQXN6salECvsqPWAF+
6s7kYfoN6c7FT9vpQ1qDbgvzHzl3hPxNP+CdvdDHEvR4u+RSc77wxNQD9tD7/388
YQsFnWA0n6gYfst2AqteY4T4gyc1d6masc2UtM7Ryj2I+ibqXPFqBnIxZEMGQipG
8NT2jr0+fP/+Vc65XGybZIxkscIEsAHtxbYJ95M3j6FlsIi1u4qUZsULNunCXxRZ
p0AFASxA4ttIoyD8kEiY8vaTxMgGYICyGT39Mo4/Zw5SxeRir6oZoqLt6pfPCpDy
DugpBokoTt2G1x0RZvarX0A80I29UMagkU7xY45shPZI01IUypRdJbAOShbosn8a
6Qm6DGOa3QgkSjCz8aG0soDLosvZC9V3rL0cm0qFbTIbz06e5JS4x15RP7qhH4c/
/1ArOk6hCBPhyVn9XnwFmnoB2ZCja4pUQQ9gZF7d/gS3Dl47Elz/r7NkpgQ6zdxy
T29GMfczZOrWPxc5rxJWabLmw27GTHYoCmmaivjtnfn2PAvHKQ+ArRdVT3OuzIV/
YqNQMsi/pyo1MSTJJVPckivZR7S5Y4GGlT08+hXYzDT8rmY7UHWx1gPJA9j2qAKS
Dq239QRpKPOaGAaGOTFvfFcYyz7Mr+hIAVmrp+yBKLvHM6PZOCA+TAlkWDh9djTo
GhybVVqK3pXTqWxci3BLPSwL1407bw+hVuJFTIXBiiSVMKPMWVD5arfpHZeSTcks
6tqCZoJfCu9cuG7RY/w/XRtcoIF5OTlhfub2jzkpcCgAM6kFMgFTLdhvbxUI8d0l
yyI6/Ribt/1+N3GGQDHS1vjzWUeLDuVP1/75argFzs5vZVsu0qRx5gQ2Z5KFnQIm
qNkrCo97iMxqgg/YtbUK1FcieQ9FXSO54M5zZd+YFQuYBk2RD7hHvPnft03v57Db
yb+obPc5LKJxR1gOCj3RM2RJPt+tpGWYhfr/H57IhvtS80BNDmPAp38EeGFA95Dr
IQHaWV6/V04LywjZ4OY8mEsI2EgqpNxCi4Y7+4khnPHouRxzgvaRh2pRre5j7RJR
so1VHD9fA8MvDNzlfBlha7bdiY3KC4h7xkQNFQtwMsNYpsx+PH9TCbFn2AILBnZ/
WX6EcBd+7To7MpxVvW4lXc8g6EzgPWzoxyET1PNS3P2FXHDxkeTS05N3qIxn44bo
3weMU77TCqCE394sUTmLJRWwbRmY875F6za4WeiELGdXD3oQx973OL+A9lmD1Ex0
CGaMqXaHDKp4CIlveTuZc2IIRHCc3qgHmsghLVyknTYN7Nbb/awNpePSOMfCgJed
b3Lo5pCegBHNraQeITlJe3BVX8kaUKufrbaKGfpNJS0xolZVYZaAOlh2z+GNWwxr
BOdhwC81rWX4DwBgxTkicAeW/fLfMNbE9VfztYvLwtnvj6Ev9BYwxAKqdSD7S+td
3xSys3DCmiPwuyYwbK9TvbmG5oOM+35F1mhTg7peJBm5iubAXhusP0NXw59Du+Fj
4KjrRsMih6f8nJeQGwDff89MAOKxVMfAj+ehd46P9s2P3fJTwr3Jq3/Y3YGEphtb
+f/MsqqJd/mpLv/zpJ/BSwqh3Vllimam4lxikOgQVEciuS96Nu4lqeMBozYsmBVh
sp+EFucwEWbP6dhcjssx/b+zdBVp4OX+WLFDdu1VflX5eOzMOk1rl/10JhNiLDG4
VU9Btn51QlTRgIhrg3XWm86XvACqDhAk4sLa1SxZK7hShtSkCUV5Q3vZX7IDTmaY
34NF7CZnbtu0uRmVyMffgBX1qCVjmIraZkxRme6YeclOFuzMnxKasvaUmYcbD2PP
kv90P1IPtDy6IQGINzhkX6r1XEW5ULxjHLTA9UYf7ZaLH37A0DKOjIT+utDUfVll
0tibj9FDda1l447XPukPJv4ZH4Dh2TsLaXXqaeT2jIGbQlkZ10ZaBm2fOAOGvF8V
UhEmhJe4xN1ie2j59X2exi5q4p6CTBtqItWLl2b+1yT0ZOK6RnjuozUrZNdDCfuN
Cy2LuEJR8TGTTOrr7bIb5+g0sVv244Ax063c2U8E96XWJ7Unlv6lG010NvYPSgYN
680wTPjszT8nh5XQQH7klaNHk4f0d1PizeIFzhqBpHIGV+tgK5te83lIAg6ZXr3m
eHunfcso3xELuAAHCh8xaoljtdEGifUOWt1bDC6NxteJmrXGblwFXsMLkCSNZSnn
1pHlgJLl9+dekcBZfA6PH6zr/hNubmQML5Mqe4bxwZUllLh5/kjcVEu3/gG6ZEfM
NyxTnstg+EwqQO8fsssnMrpDNnt/XOWACPXF5jOCqJlUBGTMUcK1jBa4nUoWdDw4
TaYtPkCH8c2D0JTvWqzgFasp1/vtH3PGzKr04FUdm4ck4U8disJOqzbTiEd729h2
bWvO3q8O/eMNpdyP4phRIsAk3l8dNcb3/4UHNRckhW99tyUnRlswh0lq1ILmFgth
jwAVC/638ZncukvXOiPUSX35i7+esdWKd6Hg2TrQgtdCVGwbVB5QZzuMOStmKRkC
NKdAZi9fbBfDILd7Q9BcZtjP3/LIoLCeRK3eMtMFiXPLBkgAxWGbYaEVcPw4/dAU
TSToiTJR0GmHsRQ2UurZMJxnYaiqzIhqoKlwNwNl5j5TvHOpvYbE71kg9G+K/NBz
ZqMTloW3fSRu2IUPQGtOwKhspmbSpTdM39BXbZY73zaPFGuQOh8f/lqjfIrlmtla
yB8waLki+vSA0kB4uKC39N9NOa5b6gxrLBs6SWPnEEsc50ifaMxhuH0hzHfqncrE
z7TKbZgGJDyNgGX+Tax+L8NLCZUQfgsY/v7KMh4dxq7P00u86kEoj5hxJCqFb5ZI
HeuBvihzuKlt4NYL/j/8ATg6chGRAIaBKa7mrMmzDSTdzFAK/lA56hH2Z+RiTtwG
T5JtxpljI/Qu9KNQUWYbJDPRQQpUBbq15ztSY1G6gp58crIziiAvleWTtSg99DNm
GI1/MvICb2uC3W2rjNMZcbX0sOsgxDWHE6R0xzylY2ndXyWy7XD25YQMWjAj4Ec8
hmg21rHOxZkrV1OCmsfkcYzd5gxTyky9ZOQQOBGmqKdP2FBG0k4URZ9asN9DiL4F
DS93rDIIgsJKQb6KEuRSCBVESX/7mnw2L1VVlW2Ah3DmsaXRX6vBYn0BUI7/bbsG
qGryOaGhxFTedfPtPsSbWzrFIso82E0iSa5ZjE+O0Pl9drLxk9EAdDgjBf8myY/C
l/kHKi5Zt+KOKfPusn2Z77+mKusn/MbHA01tIVZAPfilNK4GpoRlZqyhiYys96a/
ifRrzFkoad03R71v3c2eYxmi2wCZ3pSdZWaVfRxhdCifub4r5hR2oL5KaojAQ/3B
v/ZiBuy43Gaubx7yczwG2TcgjTPXqHFJiiBG50G9TSVcuMHlthW30WJMlFy/Cj2u
gVP5SckfjO+fFMpbDunvtlcz4rLJppALD/C+WeVZ2Wxmq0eIqzoddjUKKkhs/vUo
iBURDpeTzdbY7d/KUVsiOgF5pBKicaA5GMlth60UaFnwGp5cf3rYZRIp68/z9gJk
Xid6A7debKYfq29rNaNNA5l7QciLiyA+ytMIWd/BnRGlqB3njuw9S0nZ+om44kpP
j2hDJOSCqNazrbzCR3Mu4Sc28kAoIHMDZ6mPCohPAAnIB/1cR7OxHWpIdcQxUwxW
FEC0smesr3yT++Q4iT47xgoBNLeeABH/wM3zBzm/qIhCsAmQq+2K4xV2V7K1WKFZ
szELFdNT5uAzCxIfTsVMYdkxGOEHRgnhvwjL/Ezyh3HByfhXdiQ7LVkE/pYsN9cM
mO+TNObqma4b2AhrM7neCV9XxFrh+dz2dZJ1+W71ojFV69LuTRd8TkEMSk8wfypS
InUmVeoFVyq7r6ZuKg5dkyHDW668K+7ka0Llim9ASUYMTfHxW87FYCFicjefCH99
TIZ/Ynjst4wTcWjuWDZNa3VrELGFQGv8JcllcWHG+SDk17P0/lfOIQdC04M1wUBY
o3+PRmiPr8/p+fBPAWOO8+utcq/fbI1OfylNK0PYSW+8Ap3pm9s+UgdtIQgwzuqd
RFI9AX7zVUDBVu35FOfNd9qiv1ok4ATPJoPtCZkMT/njleRp/u2SUvvzq03v2CdO
tXw4prLq/pV5jxynzJLxMt7hk/YoXM5Fuoqc0ivzuG2WFZQW1bg7T5ZYR5M54Llh
QE+ZqHELNNP1qWqWm5QCr+P1Z7ACIpYuN3jgdYVVp8qyD3WX+xFTw0Mpw8xV2lJg
h6k3Ob4ztrWiREQrSr3npPh7rRDg6CdQpxYTi5pFmEdTaIMVGbsVXgvbhjSG6pbB
NgR4yJYZ4Jn3xDVcHH3nUpBZlvU2PdIVIAa0pdgLZGEIQkLB+ftjhPN0KgvQnxRR
zvbbgTClWzPfh1jUZKjuB+xR9+PgLvml2cYh4FlTxIHR6ZC5eqB21/7R/RW4DR72
SvJRBCAj4wCEf43d32+nzd4kjRyLCu21IeUgIRLhA6IIWYQRIVmb5BMivPH7DhKA
uNm9AnabbzxBQGskNv5kI8IW7iNCLNpQAfOeJFb5oBlBrg8t3sNY8touScuZulKo
xgpRe+2/plfm4B3/ZuqbJh65gT90DKirroWpKC2Q8H+K6QdioVvaS4Q2WrjpuAP8
nbytMz1sD/hikxDTPqd56/M2HatLPrZqSriVBkXWyuQS8WY1W0h0iE1jMX1r2bkF
Zof/S+ExCMGqu4jPoFlRfSAIiBTOW8T2bWYWAgyf2+WZjxnaH2GB14HHDwKKFnzn
Aiofe80Mwku7SbNlIk9VczhHoNgyIKWEO4BoiU1T8l6Z9Jpd7aT4w3Ml5IPoRJpT
lVikjFAKpE/D+eEQqD5EES+VfkaM7ztYS//c7Uexe4XTslWQsEi6y8iC5+hhUiPH
ajLdrycV3Hsk7J4G8bFu95M59noY4P1r63TSoctgzy+lTvhj+p964T7iBW2cPfbA
iF+vbvFK/EOOXTO8r5emif9cpSTu+FaaGT6osA8kxaNb8W3U0jnMNNu4w0aN+J9S
XFkkr6ENUBeoyxieVKyua01PPFF5gmUpbm+Z3PX1Ygk6RbHiqtJUwQ2Zm9z1Qwu0
FUx0v1pzt0GAiAEH0p/RNSZlCMujY8Ypjb4ScqBLQxiREyy4x4F5W74RYuhwYl8K
kX3mMb6pTANb/JqcSSNbVBZtwmowARsTMZl11EABMoB4nKvqSZiMQ+hUW020Pd5g
BfQrtq3Z0tvqmWb7WcxLFUqCE1Ch5tXYil0Nt8hSMvpPQMPNjd6Xck9GwCLDVcZ+
px5kVf/xSWHscGQDOLzHIjI55FApAJONjzzsE5BZs+YQ30X4xOUeHUHJzJEb18Sm
ykpCakZCnWpqsDB9vL4ODIcmiTJFWh5MrzfUldPGyTIZdw9homMqOX1Za5EpXnA6
1LyRj475w93LuCErtnOo2TrDd61azPOfe6yeQhHfdxTUVC6+myxj8PjV+2zghuBG
0jvoWmxwokf++Mq5gV5cOsK7UrrW3KOgg+Lr3qa+g3EXUetnerWPOEdigjajitt4
TB8Te2aOep+9N6LKC92I1bYGvltnHF7HPD3Rf1P7RtkADxulZj9nfg1d6Hix/cBl
rm7oNysslm2YEBN+M4yb+yz2nqB+X6GWMSrY6BakZpdvciWqr6TCnPSOKljnQF/X
jX93DVaBKWhlYQCUC3cOSoS9UYUNk7KGR4m2hCjLiTZh2wsjA0mKhK4SNnHbohz9
8nfGuA4Pkplutm+ShmcRt6QYtM5Oli43NVCr0tIHeKDjOE/eKKXqQA51lahhQ6zV
4g0k1YETmGWfkc33UZRJQK26a5Aj+wsXvfQb2p/ZREYvgH+wBVKDYxD55hQOOnd3
l0N0KYOQVNgMFV3kEp10O5Gz5NQYHYS9LaMx5wNOhUrVtzi1hgCdoUdVgDIsw9Vj
VhQ1Q86OhhQsBUdNgIP6eap1l5iBi/bFgua+A1B5iaLZjwcPLOC2IFHq2yctvd68
JkGGLUdx2Vcu23go6oIWUjbgTWbqhuAMpNySqsw1ZUdPaFLvjP3zJt8QG/6IGK/P
CnxdcsAmQtHtD/k8XWp/6xTOAgZYAUoksC3rfmakWQHM4+NQslcsxgLMzwcXcdwn
iI+eZCsC4T1gnlc53nzk79xImZg+7cCApMEqFM7LKmWSmmZXnDE0dbhSlFSB2R7v
+ZaUI6nF9iwp9G5dZS0lhp3XQMIIfDpkKtErNCjVdYe0zBxVz38bBbmzBiZhjaMa
8yF1XST8mexgeP+/E1kJ3Doaho0aA4OxVGG8P/8dS0gT0ROahtoaQsZ4QcPhsyqU
ZBpL29y1eHlXoAXDOqKMwVPJj/o1W335shaRj+Z48c9UWekt38CbcBTT5fjBDe34
aIf7np2BRKNhWVwGKCFlSeBmFxJnuwHO5HOgU69akPTbSh5VSTauleDkjpK87rj8
5CtazctGm3p/KyIr1Zv0+TqdLJf6Q2ewFHqEnnaP1kZ5/vZr99OrHSA1Doyxj4UG
BrbkqCTxALXYONfpliYbjJ9uVQVbzmt9m1GAvO+Bu/OwVHTcXBsIsvCvdPUOmx5z
FOk5qO83K2OkdE4mJYrfwv4GtB2BNwiFbzJAY7tzVxkxyRf/USrQQHC2xNyl8zR2
yQ8fWkv20N/IBW4PbSbn3cY+pvMGEeGw8zxKnbM6Bzlc1w2jAYL3b8a5mcgbycUN
/HVZLJIybvzeuyqSfUxEHwbxHbbzHS0Hk3CZGzCZK57CEtHjdL/+iRyUCwuSPee5
i2pKNf/xvJqE8p4BAnpuhrcXjFlEwhLKwkvfgK0IwB0+TikpE/RSC7usFgJtg9gm
wM0iWns5awUTtKbYRy85yHGO1NB/Jz2L9CjJ+AN01ESUitzciow1eUi18n/pwk2Q
Di/0yYZ45WSwzhRAhoKwvwdejPwLEBr++kGoccZ5YaOzsZUDhdH2bWoOnre3lRH3
LblyHEkB5FDGWwFjkkNfqdFOnTrGYCrOe9E4+vYmMH9zMGTJsmIGOMoLSoEogzzO
WkblBtwySw87MmTlep0Mumjb4wlpK7/cDfi8dRdoZsDPRNWn0gCu3/1MWP87pr3j
kRwXzlSuxvnkNMuA+fKfJ2GwLMuDpCB+O09T37MmH+QOYT/1fm8KG7FilSf6bbez
bDNcUeQdnoxE0VHfjREsGgzeCzKa68fp9VnFJXOCgm1Qw64loD54PMr+pU1SZ9mM
TBuQKdDXk1qrppIBwMkmif4uFDUF23Vd0XRCmis/5nXgZy7URbRcNbLi+Ji9L11Q
ep0ZkJilCqtGkDhVDOUzU3kyUuU1z5JU8j03CF4xXv3a1EbA7WC5Fqql2HJrUsBn
KBbyaUXqdOGg+ucMQaOwX1YhqGVVKhSrjCtZimffPQ5yfnb4tpHb66lzxslATn8Q
dG0Sg9aFDekBz174VLeXsJ9/VgOmeuDD2VTwV7h9ogL7Va68bkcq24zoLAj84GUa
sp3ynrOVCUqY6CC3qykVd0fFiE41j/wObU3mHw1tOHXe1Zcu02N2PMn0Ehhif23a
ykMXV9tRehuP+mgU4oeqDMPz7ho7xnav7Y10o1zn1TYFEKuqLE7Vh47dEfD/CHEX
haUuLlqwa3R2piLUf2pOUBZU0b4Se98mY4FEz/CPeW19FAYLLEfrGMffpgve1DDT
cUk5lDzYW2aovEgZVPZsjK6k6bcYQjgnr8l23Z5ioZ3P+B+gPUt7q/sN6ovFeBqj
phE8jUFSx2gFtIjHESAqkgf/kfmXxJ668m6jkA7Qm6C5HNfwhQxK6A82S1DhDeF/
uubSMTWGeVkXU1ngiu/SwuPUCH4EkQ3ttC1ucQ8bLRxuOQWUAFhuuDznEUoYHosU
6EQ9PpN9fHfxaWDWm12544QsqPZd/TWBC2NzmhIwTX2TRmLJ1c17TiDhE9PMUFZk
RfNkyhckXXaavZnO8WxuByBbPA6KQxg+cEtQXrEWWThtQBxadRQVVCUSk26qJdYp
x0hv8uSBwhomFJXJv+V8fcLNYqO0nRaJSSPxg0pN9q1baWXBf7JCQfZwecouU2ny
DXe/74uA6KttDP6T/fQuoNqQLoq8vu9rMGdMfsxwIpvL4iTn7eSzTWXzKtpCobw8
4sewNhHN9zWyCQRLQjFgd9kyhgVzNEEIaQKD6WDHnY7CAMMOVQZDpkLcdpkPOavG
h1afm+xmo8l627ruOTMUroVHMKgjTA6aXvVFVLqDwXxN0XSvapMEOZkMwBsNI2DN
V1L2oj5tGxgpdAf4YLJiqXIWiEez9azvu/TXcV7sz6AEg86RcwaHPP8wLuX/dT/3
IbKTSb4jaiYqkcKfJjj97iQ4JLm7yjrB7yyPc2WT/3wEIwQuL0+FW8Ye1OlQ7a78
1qdm1kWOlImT9dZFeIvQjyUuLUuojbHWbf4ZQCnVZ6EhoZWLIuWhAzmJc1idtDnr
cyXLu5HvMqB2ttSwGAD8gZmzIIzYIEKz5ZQYGcHOmxN6p0dPoJYs6IrQSE4znXtp
3USk5sLdeo7nvIwCc06I1mIsXjXIYpN8n+J1Vtxngz9CWDH97eLkqdSov2Asl96j
Ee0OqIpBwpR+Re/rTmadBgxPRkBGQbtG9uGS+7Sutkr0fNz8zMe/4zPm77r0DS/8
7WaSAGSyKU3I4Lo6p5txsOdPinpOqHzkhEA082VInH4EoAjdwkI8i6CMzAbFtPNt
OIa9e5TzLYPJHZNSUcgCxTG8KQFHMopuab00U63U3ZZw+PWWfLZ7C+9/iVvuQlWm
+BmS9w+qulBy52zsIDs3PAmyIsRc9BpX7/NaukSusGECm1l14kpmlA5pZc9tX0FW
JWcSGUGSORfh/pgCNsAqDIShck220KiRhxQbb38sDPLof4MayWzS4kySXIp+FWDd
gG4JVgs/g/ZeQeo9rp1e8kNuDU5Q/h7iETaHTUpaK0Mflmn9cYBIwCkhF6UYdwQ+
VzKXlZhF0dglChTkycSct8fopA7NBYskVQU09LmrjBYV7dECVI+tHdgD37kpR21l
yooFqev1hTqj3QmXyA1p3DMkD5BDT1ugufNydeME2nJngviQmiAQ5Hx8TkqYAKDf
+dXLdZ3+Es14D6HDPLndE8z8x3vYWyPQBDqmmF88zRcy1dfn2UhhCsykAwsl72is
YVfvYz9E983UN+1dyZlX/o/LLZkvnlCJFRlSn8ro2NpiX6pd8UPfAwAd81ws2pvz
mMiitUqp9MQ7GKtBr3Aig8/9ArYUEUJZX2jhp8vuMOxYkF6FUUsn5Qm/csss1yPS
82C/u9gP9b5k2vP9nWYQ3fKwdFJP9gjY6Rl8LEluzJ0A2YmvGa0haE1C8zhHKPgk
hwHgdB+yQpZoQHz1PCLYbOpBLNXnE72pjCPWCOzXhNwLrIEtCA/ykROKG6dKsLlq
RJG+Pe1d6/R1RRvX2pOQokBixhVexCMIb7rC10BhtqLW9SreRZlXs2qygkYuz4Iz
Dbo7/Ec+/97MTZQbOsoYLarQqzrlfXGDEBjv/Q1lfPlHTozqkhjy6V02H9g+LgCN
dA/Fjey0Ko0weAnCxcXa5mNlgMXfjgAa98k+i0kZchkF5vJ4s1f8XTub1PhZ6GL+
Rk1vFh/TythIutJ4nt2xX29uop04AS4V/zYfDg2sDc351ckV1r7VQWHJ1Za69YdR
5X2oC06Ik2PrI4P8HCNCaBssffmaM7KhDXcU1/P+F0wx12dEiT0fHVVkymPbB6at
J1MrEDWuexVBli91MA57spukzepGrSo9vOQHrEuq7rQ5toGmwoDvrQSasKNLE20g
Kw7c34d3em3/7gdQ2QYismOTPpuyife41AxB/ebct4LZKUmzpGpOU0vicm7NxC98
9r7FsukZQVWQRXXkGkGpu/LHH6v5C5ShR4cYlQsA1g6xJsR1ZwSHWiKvI5I4o/q2
2S3cfR9wK8/0nk3KVR478ZgpLL9ESg9y201mM6uSCKQt0iVRclgaPz2EQKkBggPV
67EqThiH2cdinw8cmqsP1Oto13Yt/6xVtNBN3Y8UQAdoEY1OuR+iJq1Vd46OnoJf
ZfPpZ6YhYMN9A7o3ACvUDyspN3kvjSxRuFY0H0p0RJ3B/P6lY088EkLjIxuUNs1o
ka2UG3quu+7ivx6HxBfAv9eKAZo/AItTz3jENp2IWhajCzULIGI3+6EVus+eJ3N1
y+1WiZR7AOOZqUwUIh8lPF3rzOJTZSVkTQby2fEgcEOPHh2pvmpM7XlFmUV2heFd
j6lTRLQ0iUc8Jf1r8Uxaif2umYt/qjexKGQdGFQPcT7d8pYJio5yxSvqPSfikhsz
UOug8Gc+qo0tB1Ce2l7OTUtgalrP7Z94+evYsQqvjCDq6oplAudXOovWcu9tZUx0
ff8bnSELRqAJe1AdMGuFFextUUGiXyx2noTaqyQ9FcMxiJ3Ii7kp9eMhFGoX7/l3
VpgSHJxxyiAh4vAvu7y201MJu+SB8AuCHRFy9GhXaasauF6UdQkJGhbdL8fiZT58
hwIauAIjMN//xhqOxtaU0d+LQQF4NvD8dDGxSU6d53CDjWfWAczheJEqblGo69Cq
dY3FTqzhlz/QGjBZzm7c1AQgvNskA+4b3RKca7FShiUXl6NcLyCCEj3gwbMB6aTo
fsABEbkBQfcDg9bgTjK0L7WoZKicNVFuG0RaMHbmlT1qvJULSOpIyhK4E5E7rRe6
wrzWLuhqqgRfQRjQrS77ChhqzjtAu6YzWDoHWwQuLGK5hfc84Nps5hcmiCIDqaT6
1ZI/MRrluZcZtz3H/HN5QMNeTprrtICDLR0izOb6VfQCceSu7DP/71fNZoYFRzyt
RltoGguI6WcNqFg7UTlImEV7ZM249H0uQJr+dsBuB7zrnU8AY4A7kh+1tQ8RddlR
WJ3/Wv+cUtYe+0VjyWafAw4u1YsSOS8rEDcHqMFKwJQasdjy3gfeZbHDUZY9Evf4
f/H+jX5ariSigm8fqNdBnmwuzZ6KAOJKT247F44H9MZPjRMi1ERNV29Qp31nTbB1
KUsd31D4w/Fg3SHecfi1Ztl7jOJ5AOIHHjIbeNGIiL/KdWX5+u7T6YGUnLzSro5g
RaF/sNA4uPn5Kg0qMtRm4A6jVVTXKDX9XMxNddnJ4ls3LnHr9ELMZHOWBpesANyo
w1kScE/un60mQpXWsFJhvyIYQJSPc++8PaqM9cpBtm0OeJo98u3oAohvEBeVTj/h
43AE3cYzK532lXbee8WhpiT9Hnlg48ety6wOE+h6taliLZgCBVDZ/ws45WHB6TdT
Nis1FtHNfOw1Z21hKXW/Gkv9n8QTJiBew0mrlF5RFlWCji38h87bYjpWcEkjS7/n
TfSQBI0d2OSNH5y7xn/2xzv6Pe5DFApqmGVW6/BCmsxGivji4SaFldFCmBHFM5jA
jx/k3Y2xWHHoTn9ZTenj7ztKXNHjbajXIkSmkYXopx1FecsVs9n4X0Eha8sjsAIH
EpwTTW3fFDlqRV655BBl41+xA6yPbfjwTBC4O1CpilPVWwgbvKa/gCj0bUSIjxH9
Bgw/DP7yTytShAVQP0o3P7L4AHzA8//BvwmQzrE8KhGsh/HF2HZrK9d1w5XxaXLn
2t/99/5pQr86sF/iVBC1HQ1LR/zKJQvyKBMvJFFSf+Osm491Pxaz0TKhjQsWHwnG
maTLXUMkVIh42Kg1t3A6hXGL/s/F8JMmC+wx9GCkGz2w7HV1MaQ1SEbtwm5g13SD
vLV+oQuQZCyk66VXOk7mNOz8j7ItclmyG8uWvhsSNu6/Zd8qu7KelgkNTOoqg4ev
ZTo7o2qZE8TKvY0fQcwiqSYJb3jhQlmJ1QEgSobyYro+/NKklgMwIHeQRNCe884k
knasCacbL+DdsYgqoHSQG21brXVZdpPGP+KiTguH8lcsCpXvhO3Bq703T/xrrNCK
NRVk7QO6bb3mGRyXg/EDnTcKuPTZYGEw8vKVFHEigO6tB+mlp3rcttbZy9eL8OIB
WkiV8HmqKAb3OL1uTlx8y4RV+h8na6NF5fN5mSrNsm10+1jOkuzV4QEG3rH6pmNh
Tpy0JF9YBZjWL3wp6YDAjyiKlDKjnsZEPFhy+7uXlPcgRRbh8lzR1BZD1YZmp4v/
/Nf6agR/VAWvnlQu6Xu4hNoKHNhFuH2fER2suPad3H2amqflh8NHMTGSwbYp+CMP
FW+xExr9vmsHj1W0fU2E4vCS7bTaiBVbIn3X6UuztLvpsQLVZO66FP4vR+lOKQIk
gm/z81f8tkGdOCCUZkI8jYkBCZsAGcNeSc2RICL1UeQPdyORo4uXUJsUZrjzg3VD
jFSNV8SHZMbyCqJHvJFDJMuABYtGqqahZ+QExsFojDw8v0I3UAvzJJOS2JvcMOJp
siAHJCPwDEwMQaHurwSs2TabKlqfw1faSQ7puQlBQ6Pbahdy1trPrHAbIEwMwTXi
lFiApe2YqS7TEj9rXdPXNW5X366v9ymshSlwNJbhEDqvY3f/q2LmINFq2RgGw7V+
ueFof7/fKsmWO5WOD8CLPFo2T38tdFf1M6VYooCZSZ2nXBth/kSkodI91aZW19lD
X28tXz5Svn/M0tIkVrPEXfWOc7LuB4VHmyXSEaZK6bDkVXTGqdjwEHy8pNZ0kUVJ
oAuTsQtPThCgqA3yP/6bfCKe2km9rzsKYLtuwrr3+DdutO7HGzzMvRn79ZwVIs6W
YnIARfKZ2ApFj/2Gj+HaGmBCWhjAfM3iXRgunGL/VSTDpjWxu1n5yaMV4opRosO5
gtqV9w4+UejUKmFqPxtdVXtKZtToosIz2znXAGY5IBBdFZudHwJhGdCohf2pzd5N
1RR9hlkKiQD3sgjQUahPgOaVPxtZWJudf91zOuwBmTwu3lr4Jgdz6zjxW26vfjcQ
k8qrVZqpGnDv8m3ZKWTbR+KdHyILlBKn2p6Z/lO3NQZdz+2DEkjlWH0u+QvXOZxw
aVxZVUB1EXjiHYdmyn8VRjMFExuxmP/xuziFAF6NPuyp32QKYUyXAkv3yziqSO39
Jwh+0EAJ1kd6EQpxZhXewLvBT3XA4Ukbo31k8gYqf5XMmY5RS1t+N1VX13v9Ax2M
mrwdR1imGqQlAL2qPc7Tmbfe5tJxMT0STWNOH5/W3hmzEjQRcTyOZL4AGcsNbTkI
/JRS/ZXQgSJkHFAn2viLgf76jOx8JVnVj60Kc6jZWWg9JKP+BjHryB9R2ELEatul
xDFRdDV+x07XEfmKF7GGTJsFsNvtK0LjshQilCj26kXxiZoGgr2YVdRMTmNuJ21Q
HoJLrpzt8c3Xat8PrHiWuBCnkj3ABJg/MtDs9rwN512Qy0NI1OTr2Z1+Q+5KeW0N
QiJYTitPfg8pF5W2+NO/hKwRkpBGlB5SyhNriYCf1A9Y7x60MRTzKd+NMpfNMgUm
p8h0KglWpnxtSPVYxAmWx/HDmL2RECdJiSBFsadYrgwfAYIwv8sfZfQZWJZeMeSm
u9Bo0ghpLs5A/nSzM/hcj+CBvurwwFUEyjAacKpefaciDH4f8fKbS6Mdcdf8l4vk
Po7TS4INVxBYscPaXXvTO8zTJlYv1RSTqthTKuElGxGJ2zj7jOrg3UiKRCISdz00
F7DgmeYIl/jBkfGUUaDELXic3mRQ4Dgett7pL6wVkHWV1Yyob3zcAvqdxXi9ml01
W9nker6tNE1gBhvVIOkmc5tzgG9f+zrFTdyL6zEOzADQ3zeYE0pJqvpmvAGKIyyQ
PRdGvmXyjRoNCAOkehJJ5rVHEDpKc7v04l4ubOy+iHt7Zvmav17V6kRa+ZjT3q14
ZqRo3YhJjcG9IjC8JoJ70D6pxkP9bdof8YG4DpDPt575DwoMldeBTT8d3h/NEGt1
oqw+x4nblRJ7bvq3DLC+/P/0Vg65/9+9cNd9mnf/q+kMNC5PI6W9e73S/AyeaIKR
CepBYRSzspGRvTqwa/g0KjQH3/HfsVimtc2CRAQoBMOARJWYBlxWZVj4WsReYEjx
l5wceLa6rP+5jxzWhpL4m4ZO6hP9gfPiXXBzIbHCenK38BZf/B/qDQNF9mgSK8mT
wcMUMovfrcDx2BTmdvshGkqaGCBCNEYavEJAemWJwbG/zRkxSo2osZUyM48rrXYB
40JngEZCb1Fk9WZaEujeTE9JBc46qJYBOS6CKy9Xt2GvzaAZNRPftKe7ZujEsWge
O+5gnhV7jKa3CM+MMLKlgaWKFIpM08lKZvU1uDJvVkywxXxO12/Yws1prq4srH2J
FRRFXv8hOYHCvk6lMa4ru1bQAKzTdgodrUbaqQ6UUhS68tkPhM6vsyScBEeOWnFo
Lael5F0JB0g4qDWweEJLixMFcefBsNchdZBWZpTzqOE1TP5VjvT+E8du/TwUTT89
GflK+Ou9e8OhOWK4A1TgG86uUWi2Xaqtz3YjufFhyhc0NUGacYGDNUwbV8mrvYs1
1QkJQpxl3bZoBn+FGA8vbRECsU7tpDlVHe/cQmg2B/IjfrnOitMp+b7T3Dj3ApGE
OZjWhaTlBGs+GgKoOPwQVtj1Q2QkxTYiatS0AANZq5ntLvlmiL+C7ONSXsMhsvti
WpsflDnx3cvw8tNf2GuZm9yVl0R8YcP4a0Wn0duBKbVAE3Avk/Xth7+nIyRwQzS9
ssRqqRD1sSVx1ZBDhZCkGH6/B4rDkary8iidVrMq4UjIdcKAnzOIUi7r98oHUYkD
S3sGZPz6PVbBg8SHt/gXNtyvLq2zRAMEJUNrBVBtfbvAgIhdDBRkYrMZDKqm4yZP
hSSXmo+qlSTej+4BaQPp9Vw/Jvin5Hb3P/nljxRGJcsSm61GsnGzHXaHDb3IRfwu
PHnhxRWg0Y0zmfSr9mqBS9KOmKQYBX5G4UoWML36vBjnKFg4OaAEvlOf3flZZP69
usQkOJY46Aw1a3zMVoEE2gDye7NcY4Hzb4QWkfr15hwxO8C5c9epMUsaK7fIdfDA
74eadO+ZSMdhP2D9xXQT4fLamwVzQO5vARc1lewrpTajYKJCtmDXBMnX7//HAI9X
KWB+PKeawLiaLOT8YZjK7rNrcn/amh8fnlPOhpMgml9XpwyFKyi/iXwofxqgRLWz
vvaJ+fWd/9i6bAgUpIrb+meqPSCRMUmTLN34TrWiwt3S3UmPtPnDZ/UKjt+kB8x/
URbz1MRaFSDhn/oluIo//+yYr6yexJfogIzwm1eH+nkTY6f2UsmIimexXZFG22dt
mtihjgwFpppZ+UPM2rwzP/Xz8Ygc+qwpa+pvY/nWkkroioftZM4gTbF/fSwgRZVS
6Ss+zcSxiSqPoLWKXAR4hpgqeD3Cag6z/kN5pNapgnXUASyDLgesJKZj5MkxkOf9
eFSWmFrG0hBS81bbVqmZtFVMK7JdW50AkcwnuC9Tu+yVMIWIFmFkmThLjV2d7y2A
aDaLHkIl9TfrGPckZwuSrTh0QY15deB+nnu4Q2IBOXSAZ23zGBJoDNzgXLniN/3N
8FbdpVe/FQOO7+tO96mvoTLCkssSr6ugePBHhrTJfU/eIz4xC/KcdkMXIBJOaEIq
LmllTbEwnm8reqCgjFa05Y7LrU3YUqob2Tl9Ur9ZKGkXAm/CFhz7SKoqaHDxTMBW
BkqTVZ2IGhGwL6JWCxMTI4G4AkwI3VKMkov7LE+GDdglxrdCilJm9w5yRGReiheK
QtPzr0XRG6GUiJVXCzE5XLIQNbu4qR2/iQc60Fd5XWQX9DbP+LL7a9MhcVc8k3sQ
mMcmmKxn0GXKN3oNTrRFS1b7p6lpGTGUosxbxfvAl8yJ1bQD7wuIIDixj3hvAJzr
wAAayCetd1VkyfsRn/ZlxnMAHq8oodJBzApk70Sq62Pyow+VOvDcT8TZRrKYnruV
f6SPiFy1KkEO1sL2sqg0MahBd2GTVIYrAngTXGZ+m6YzYkwl1iT8B0b6zYvF77RX
aN/Z6E76xWIAiAJYKMim3QRMxKnR+RgxvNY5u7Vazje3lxXRVXeRuld5xHeKmnx8
MZO19OET/ai+vuUyo827ACK08YOKsWvt6ZW3OkSIaIqwzAsrfMqXi8bNTQMn+L+u
+c3duAIU6udx28YFEXrgiK6CTb0yhb2p+lrQPd29QRaQOZLr1LQit/J7GPcRoBRv
HI6s4QGVwSjNnX3THgLjz7qWe7n/xoWZZEueSyzcJOvSG6/t2/St0HkBp4QVlTUk
Rk3sUZkFIFiQbeKG3JdShWBgWVdgidsADDdCGbjHmE5tNNV7GWO95TgLzxpwbwqs
rVUr8LrJKlcMnEymaoR1siTJFdGAVgxFkFKjLDr3pCZA3gJ3/palkiGgKnXrc3KZ
vgBx0ofR9z+xIp5ReUZNUa58bSdAriU2uMMkYnLVr3TW0rfxGm/tKU3h9Rj/ybkk
5bXBIwNchDeTiJc0Tujx/Dnvc3zfa4gzFyrL30TWGs6EVFUT2TvD0n95Igo2XKNE
ORmisd6rGdn6coGd+UVjD7xuBiAYratFZM2staIWVnl81kYrWvXIpgCMniC78t3k
K/+Y5Lwkh9Coytl6NT5EIzs88sXpHmhqBnebEf23Or+qONCKQGH2HTeZ64cvkIBN
DjL3d8FGcEhT39KMRHq3OKFxNyJ8O74jPRcyIvUGpU3d8YXINQaBN/IGfkDuWd0b
1gmNTgix+S6FZlNacO7RdV+fyXlGWE1AAn2jKoEnmfl4HCmUKl2UGsSGvuhlLgeq
oS134g2z1oISSDQNlM9eQIxvRhFMJy7fjB/sn3aTfMYV5Ox5VJdyAFlqXceJtX93
4S4JqkeGAkY9QcIadOaQ5Msop4xCz/fqt6FD09ZqBbbJ0Rt9ifszdH9C6opBAPhA
hwOZTig+dpp9h/NuFkcPPvmEdHBuWagKlcloU0ciLEWLWqtjTNuOXxuJ6msa/qof
lwCnDTS2Eg5/jKB/IcmGzp4L9z4KbjX7z3YxE5pdIHe47+YjqoVy2zOPRWm743Mv
5saXJtmIEoZMbjO1p9Ni1def3xXn6P/qMFJxAJvzE3daXysbW7yc4TFpRJ2N7UAs
8sC4Sp2OeljSBycdjJQNaeVM84Fcbjclawt14TZxkh57GioDZP2B3LbaXMk/6TQu
Z89OFM5yvjMYjJ/I70JDLYuNGPfiBVTjdJhdKW6i+TmbgrQPgBRms7jxb1p6fgot
cLvRBWZV6GNwP2QnMxslfeOnXgzuiWHcR6cxABsecDvowMzzs55MaWLQ6JKvizyp
ow6kugUPCRb7MA/nFt5QcxUlkTYlx6SpUcbmSkWdp7N2BbbLiYmx17bT6PoQq+Fv
ODrFaYc9znlzPhFr0+T4/QHXdDhXu6MT0UgLW/LYmm8ErATMofM3DVtYIwKjOohH
rMCBZdq5yIdc09QncbPgi4IhWCLzG5Z5JOgzu4AECz8ngDYJV0FIBpQ9u0Jz9FLt
LqpIdU89Xr+FQyr5aHFpqybqx580yuXpF63e9bqbbbWjhL0EhhoB/y7xQo/xwON8
HYEWQqboVwQeFeIAIdHZ4wuFWbdhXKtL+Qc1xPVu5Sg8gANn62CZtrDXYFyzTu3x
7trNDMxy9TdC1KXHUOmXBnwizR+aPIxZDJ07mtVxn2+RNrVSoqko4TuB3Fe9G/RY
b/MbuwkbX9yB8myklXZ+NajV0Nh0b2lOuqjDnwwgrz8tZkPxelXhwaKLBcTDLdUB
+0TOC1SqrMg1yYgN9hJPgBXN8vZ62izSNgkFMblypEJKZ1lsbXnAi/IZxe4O+gxJ
3HMhVMsBuyF3Qo9twYqvu6V82aQu63FvyWphibO6GUuxgpW1kqAj5aCr/JrhrFBm
4qOx0H/INoTu+M8p2CqpT5nv5vHiAsRFMYUggkUhScF5OzbNCZWLTWnb6gae/Mxh
tynRBMuDTEkcCTE5ij0Ac4BF34jMkUXH3Y/S+P3xqcanj6wVLmJ2bbGeqL6wS7PZ
R4o2ltQOLim37K+RqtL2LT2d17dUTky3Pia8ydsAN3LgLZpChQgbXd8s4BLq2dtL
gkO167OcsrIitpm5IqMIFHwMNizNahnsGiBcBHVbDinWpA/PGX5rpfw+qhEfCJ77
V+lWG+J6MkGQ3H/9+CDWl7QzJvNUn1f5jtS61Mgj978aH5B/TJ+sO6FgYMvQXN/I
KKUdJElgPu9cVBav1gfVbWulK+jTM/eV3hV1dn6I23AzHeJaScpRB+lJynEM9jbq
Sk55K7/iY4gzBjnWGpMUdHQtN4nT7sP8RezKCpmtViEeWe615MCrHBL2RJiGQx6h
dLNjZ4qzDfCI3oUXW4gQLrQRnHKs3nex/jiVbfjlxX5grseatLAljMKBbxY4sgUK
2IdMhx5VJRizbsFpcAQfBIyEMp/67pPRfKbL1Urkw0wAzCl/5BIvcbI0teX1t8Q8
z7c1RsMWCEOIh1hFEJLL+KImyMlNr2RkI3NOrGVcO12all+lZ7zLTx8JZm83p9pP
cQ1ykyotFjDfT0Z5xgozB4EtnUtEFbisv+ubCo85uO/g/+ggIfuvqlpLA2mtXmB1
Nsgz0YmdJfbIwx3OgRhMps0cCCLOoH75E3SekJp/FxwDTEa5t2SzzHodxyMMv3aA
Gwi6kgbQ+TfDP16DxG9fYJerpJwykowBtncPrSnf4S4OiNdbECCE2vGz7exu/eHk
8NALXRy3jmNbUZ9F5sUzRSi8MJJKDQh/YiMy2lXU5+fV1BbngCa8gs+C5WkZqHkL
PjkRl5hH0UI4ogHk69mN35Hy3VPaUEI2oasEUgsNMUpWw8Q6IKoxIppzGqvsQToJ
9yYOweIW4VIRJVwyqU0HprBYFIni9AdhJuZwFclFjFPe8ME5i+tgPa/AQWBGKp2l
OpQabDIGe92KmeLevtQYZujUMUtn1PbeRqOJETLUWOgG+BMAsAFdzKhUk6Kqj2Ri
IWT9d6RNVI3RJyDSsrUc3yaOZd7PZpd3sT5xw6EY+eDqX7qFuwNkaT0nZRiyiuFn
bcEc3Y8xoFLl3O3/5lJge4ksW+RmAGQw2j7UFQb0VADbXqBCT7pEM3OjeWG+mnWn
bbsGc4/e8z/HffitSZSrijCzhpYohCdVIutmwSGO7+TyT56vcZrVna9NMC61W6Mt
Ffsoe8FSRFheDj1sJ9Sn8scTHlx1J5EM/v8Idpu+s1SZjsv0GMTVvzt8vv2EjO8T
ULAxHLiQ9cIc+yjCuUvvtKZGsz9mJwLr5+mdGnczhLVOvcoBKPe7tgI19C4WpVcD
CXP5Q6rG80pmZk4cmvJ//lvNTHI1nCvLLQGWXwP0/9ORxOH4yblHPcwwfUZKJZpi
oThYItNHTeQSLPWhpvYTHq9OttatGSWOp+c/+U33sSVdzluYkv/uKGWZzKmwJbFw
kYjxTPIrI+/w6F1NIB+q85acOcqg8Q04j/ZJreZBpT5hDnDCzLbhsGP3Sth+lTvX
AxNfsWMZ4Zj2fwSxbqlXTRg7yveVND8v+oKNCCOTSlA4a83fN+MOILI2pkLlxHQ2
Km3QSB4lzfdXy/AAK9F5SHtUk2G/4TwTigTk7w7B+FaCKC8fZfMHkU9gM9orGbPm
sWRvQk+M42zNhs2WbtscIVMe/oyx/1Tggr8fifTwAYj+X5gA/zek5/qX+K29TdDf
h75JctsQ2r06pHqlqMPr/uEntf0zIN6iGyHVx7wR4Xd+RVSjDIxk3dUKM0IAr0Vg
AKH3kUYThRwe5oM5P/fTfqY0d3BTJxr4dKP9QqEeeUtf9UDLx9dsynCWadAUuxPd
6E5qA2/6P7+3gq4B5Q+YEOqI5ptkmtk7ji8SaqorH0b1KHgtaTdPLEwsOjsvqdnf
lOCADK+gr3nTPvxRxf1qyjlaUGS3ji1ZreXOJfdS1ukpwt9tvdIlA5y4h1rbYWFa
W0aGbQux8i0shKTKkPv+fpyUx8N1k5S9AORIUxtrXnY9iAfs4dxh6VtPIF/rI59O
jBpoDZrCRm3fN2/sh4A9hT2k8S99EyOBysIX1MD4Cec7ylNy0aqGZ0qTauPLv5/c
6G4IPE0WS0kGCXHvyImfD3ffdXGGxTbe1/NIRT8J43pmCUW1QUqeh2RLkbvXEFuh
9pRZCghEJfH8xPbNxSvXz84Pdb13ZGYRf4Sqvk844do0PbrdEd9pTGxAnu3nfiiz
6xlCzklQR/GLRVA6wwVaH1+EqaAixhMDz+LfhdR51qbYSlrsgRqFMwFpale3hQAB
G+694eaH1957dckDpPrDyN+1j3VGmeMzes91/9NlL2e/w2ldb1pYFsfh17R3iqE+
cI6J1QVbsHvVYyRJ4UmeF+VOf1eM1fqrHxC+eeNjJWwgPgI2TCaHQt1ITr4hbmMP
Fl0YGWC6w5Dylua3uSOs/BqikmuFXe19vJGogejQsqo1Db4GZcIo8UjdHTw7nMku
WM+VTAhA7/7SYA1ZbhGRoI0wy5jhfOHSy+n//xlxiDbtHLpJR311r9xH5dv2PiR7
WAs1ro2eD6AC2/pOZFLqua7TfRMyPEuNe+Pw6fg7Il2Pk5oogQrY7Yqezp/FrSbo
S38r9/M1gBGXmYdcnRn1WD7yIVNN3QTImxtCjW1snJ0bAlralABJ3QkWK1fVWr8O
J1VlXnGnB0CGFAM8aU4LEbVasZRpSkps8cp6sX0cApAlfuSYCw5DZ6Y/j1otyWzR
T7mQFx+v3hpairjmrk2f88mWQvPImvSdfvMvjkQKQqqI8LfPj5nPV9ZA7aN3Engd
Rkgkj+F0XHKK6WqYUKl9yADWL3/An8CjNv1uDzAVugI9cqZFij5sQSNyXXi+qOPV
n7bAySxoU052SwCWbCCv5Wzk4Xzo7S+RSVuAX+tGmN9OPJgO4Rlyv2C6Zd7RQho0
bb5mWPC3C3wjQBa8nQwby4H6cncekfpTbTr6yLt4r2QHL/qqpGA8N/tI2PE9rAgo
H5q52xDha0/yq4COqHwSivicLA2NAp4RGkKK3qPsJ5rzghR0ZoGlxqdr/5vGBfPS
K+k0q+zfyr+cyx0Y1OTvpUxuKPb1iLfGyd069/SmylNqk/Cq9SD9On/K6lWwUkGR
YAye6CvJC8G4WGP8TeflqOuaVb/nmvu54KA+JEGJWAEtq82HfNBPkSEY0qRF3kfr
TBbSZjLp0pK09cDoZ6oIay+qNEqzKlv5A6wvS329674YPNfTJY1r6VDCLCvcs57l
xql9DLvjfs+SeRJR29GYgGt6hCLohVuv0V8tgI2afuPDaIoWfRBuRsF12s9VqKli
zFj4xNp2kjbPQ2qx9M4Py7oiTKAfkGZIvyUdlt/D1AFD9pjYGY+gd90GRgUTOdH5
vZ7a05iBLKzuGGWeMOGwlwiq5f/i6/yXBiIjrU4OrCOvC3o2zapiLLjT043B/Wf4
J1TQLxIV8HDVE3rD7D13hJQm9SEglIEnox/gH66IQ8GMtRFUxaCXPaiX/bTHS7eV
Ciut88/kdYsKk5pLaA1kNGq+t/bz74G44HaOeAJpy7tNQ9Cs1rmVpF75m2VZmBYE
Us+WgD6NipEbyazbGNNu2CJf3LMvl/aGv6XrvYKC37k+efXnMXQcA4MBQAueTiBX
uIsg8olVG5tZ4OoRZb2F92DqNrlGmweb3poKJlbVXJggQdsO8UCTqbjGT6a1lyRx
omAgN6Nd8LnP3k/6zDr27s26djDTwWBr2t+12i7CU1Xuti2WCUdW/Pz9Z+/xU7Lm
M6er18tN6BpPDQ/jFasiPnmASewMAgfjRCBGWrEmQ3e24ek/NyeYfluwbseEjwM0
1NGlebbTeEQioYOkUg4afHfktyZ6og3Q5R0vTF28TJKx55AWu0nY5DraI0wumsxl
ScMqORlf+l21k5dfb7kImoWxGA2AKESA309WCucOyAwt/ap/2nx1t4umnrV+Kd+4
tOa6OxLEYzM4cETchpHX4I9LQHzKcsIjuJgpWBGyv0DDThpW8brodtlqr1rwyZQN
TI+BwTqHocAH+JNIGENiztO+fm2joM71m3d6DzBz9eURG+2rGO99xOuwTYOzsfrj
+O9TOAeK+uRO6X9Urr8RSoT2/u99FQgAq9VEiK94dHjd/gjhI1cImu/qeLdvo74j
lLhmbfFz74UIfWCNO1RqztUB1c4vpwTsEyrbfIQMWo8q1bh4vcYsApbRhaQlo5+t
ZNO9xzbIerndAiifj/nq8ndTceDKUDVrBHLOl8k7HENXNVpumSGMZhVOIAhgufgB
Vll2OoycrwWRC/MDjhJeLqHfey8VtgrMhpL0nwTTUP/G/LVe+EV2BcjP1OUDVsUc
QghjHlx2V/Yks56DhJpGwWWiAPn9R1WjCZ5quSXerbK4cbJISemZeKArdTGu9r7b
oy8qlRKeaC1Ck7Idy2K+ZDYR+6kIMlaiie+s99Z+lhokZZvIDsgxKG6g/E/PSTCm
zG+MI8/xUTJ+S5nlooc5KzvsxuH3DKKOHyipZy1TfpXyc8QS5066YdihWNnuLzMy
csG3/INf9O0qKkfTOvHvszqLmpGF7RIb6+IYACtHqy9lJyBWdPJqrpvvT9i8k0B3
xzIRKu688R0X80A1Y7aRqJ/zpDjeiq2HfS7qw7+t5ja/mjPNRJCNnC1bt/W3x4jr
by2GPt8Q7ggGUZ8WdkgCVQxOFwtVm8EA4igp9XCKgLwKy+qR5SRt5mWW6rIhLW99
lBxej2O6JMlUfqKnBUEMKdlt+VSjjEfaFX7dfMf/WsElZoCzwgGLBSaZzsfoBKG5
vNIzTClXxeXkjttMnyFyPZNW9FXOAT9KN1RSidU/T9dow6L63n+bBCtsYkjYObAn
dJwJo8WKRKNmYtckyIHzs215MQhY/ZEtF5PF1ZWYkbw6nSmtVzlitVqj7P3FkwMU
ajBJmLiQH7S0symTioy4fnApjfvZuPvg2YekR5zR/IlzGeTIlfCsbTBB2MwRV5XJ
cGnY7J+/MygicbeSpMnrIswicM+0ixBv4ifBoLr6K5bzcbeVsDHdVITLwuGOky7v
ZRuKxcQ00hABMEXlNUD1DJATytENuWAnQl6b04Ym15nSwCxKwddjXfz4chbp8m+i
Gl6mQ8j7PMlqSHUQ1Lfx3Tb2fS0h3BvKImWHXnKCunUU93MRDOQL9LxgadaXAQZt
FdQ5CjFz6wOM/Ojch/OT29jAXbOOqiFuKlF5Qg8CHyq787mdfSYIPipGprId2BBZ
y6G/UFut24c7idmSMM9eJUKiB9hTPYrjWwGRbypsepAkKdZPbE+83tXDsttIvfTT
i+mBjz3MzlsYbuHLrJho0SaP6yIMJQ7aTds/78CE1TSLxxxwvE+Xzta+JcETNLm6
qZAeBaYPv8e1tAZkK3zysqU/6yQFWZcTkb2DIu6ePaCIiTGICtjmlMSPQYtJ+nqA
TDJfBCu2CSedvMff+KOp5tWuFmbbRILTK/1LE80bFRkIvjRE9eajdBI6TA3nElID
XiCcz1KjEWZ+cp3qZnZBk3GK3OOOmU1ascp0vF+rkjsfbZ70nO4Lhld+5Ch9iRCY
Uni1hyvnBvvaf+l9kOvktYPJzGR75rFk+50QNtBIki9hh2SoNLIYJwdansAd7k0j
q+E4apBYpSqun7hBo32VQ1ORzyjn59EgLy6I1iUrdxjA+NB1xqhNSMyh/t7O0eD4
VGfok68+0Lr9ET+9gQsQbdAbuo1lxl6xSxoEYOTbMkVeZgXuTEh8yjETb8nLwHd/
7jLcn7slXummnibUOE1Nqr2sZNBOhyehW7YLMhu3Ch+BzOxaAEgrxp2WmujZc069
ZvUqzKiBcsVP6UBs62NQouUKIawU9Cu/UHpWN7FVXL6rEWoRA6icrKxGUUEc83s+
UjwlXKb9cux6HHrBuU5ImMNOiilUfGovTqPoopwI1Ct+jPrDWpI33nyyJ2s6L+x5
OgyhuFaU38rIHvN/QjAkf1aYnL28O1U/P3N1n92B/ffsfV0TH09jbB/zqmIwOJPi
jAv/zCLCpMjZeSISodiLBlv0VLMtGk54FrLjtHhbnNmMDZ/hHlFef7jEWNMNMwye
Q0GcOcb05lDO2EsxFPRxnRqZ+kBVrDB9C5sz545GbeoU2Ct2CKkudZmVgPJQOybu
D4bLu7asfjIMoOMluw1cvr0P9SFQS0FtIpzAL2k3rj5tO7dUQyZV51cLU6X/CDeJ
HgCZ7SmG0XET+wztanLG3gYZ7lVNirMz6L81f26cPF2pFyXDhkMXyZM6UxXT7UY6
HyH7T66fr5YR0xG2oVthUqaavp/E+vLDsX4LkTZpZ6YErZyxEaqKt2yyDCzgRNKz
SEkY2s47PiPlSrsWPrxSeO8w2x1iTkvyNWL032xoupW8pAFPZ6IshBHSq+YTBp7R
BXbAGF0053YRNnO2f48Au8fwN/DBeYBRwQz/uyL9S6DxesGwwD9gRNou1aNBpxnV
ztErV01fqzEPKO/7Ky2PoATBwSGnC2tw4ol93NRvPdfRE5PGXyshS4UhjazQiJPx
HWO08VhAsLMrwqa2Q357XQ97KJlSsUeFGGDCzrNxRffkiN+IV+1+mLW/F/jFpokg
KEf88X16M9xUopqf1tlyoI3arZ++e7tm4GXiBUK28ufcwB4DJhl/IIbKnMwuCjmb
KN+AJLL7Uj9DBPpWCIfBuj0Pa2qNhz1FyePNohGT3syQv9T7MMDWg+H2IjXGQWD0
7jVXh7sPeo7ArxkzBf+3NK0iDR6gK09Lt/UVSY7dkglfMvlXXcmHcJOr3QMhE2rV
wNTGoaUgMcHgWmXal3H3sP//O6r8+zyKHZEE2JXMkLLcj0WUgBE6Pi7vbMzsgNK2
+YtxQy0gsELlNKR0StcX2NWmDz9N9rAnOWsKf/8tUKPG6npRNykXetgm70D1sDcv
kEUQZ6KYhPEz5vpUTpEdePhTiom1xiSiXEr6CsxgNaILRYCPnI+6cHCtyENzIWVo
+9vHWDLlE1cu5VKzLAUXCbhwnztP/elk3IQlHe1ujYO7elnjKqikIgNQn+CO2QCq
RrwAHxjW9q+7RcQtPGbPD4N/WTfwrZtOoKTkc0/YfUldj31jfHpM4b//VlpWTr7C
NjZXXI7rkFk/PfheWRfOZ2WcqG1n8cA0s183cIJQ7LjfJpwLxq57xf1JWJnLSK8/
fTm/zE6lBrhkC33xGv3P+cGEv12CFTXgwq7J5BiWacHy6o1crARrQ4pZlpkEfmVb
X0gxxcUFNjCcLopQU/wgacffXeKsl9VXk9kGzSUX4e5xDM7DbA/hopciZO2dolTY
vrWbiU5mCgaA267I0ffMdT/XjdOhRBtRFV0qIgOsKmf8uU1pRtzRgoIDtPsWgSXa
hjIlIHmSFfgzUvw+d9Z2Wb+Ul+sd+Qoa+z9U6OFBjeoiT27bcnQ3mh0Y0PYl0UYn
rCv/axN6Z0ze6rVkCwfkaPBOzZDHML6u/QDcdhZP6umgv81h6ZnLnjR5xfsoIdJA
2sIw195h8C8AjZxUk9nk8LfMqTKddZlMU/uZhlgun95KWZdgxtmI3/Dtg/9B0Kjr
da+ePTAj6xsqJjDcqSqVv0IMt50dut3f9Hnye6WtF1Rex+tXChI6l8Kv0W0pRjRV
4+TAeyhIZeBhw1goFFtNiokw8DvLFcDpzIrFzxB3vnchef1G8kO9U1Iw1Vat1pTL
ceIRT25r801Lekuo2nJ9sSllXqtEKeEZ7O2T0QeJDjtY8fRNOhin04hSf8OoN73g
+VzcE2iSitT6VPN3BfEfZ2z0bkF4IucsJo8x/bj/RYf69ulHr7hQ9BLy5IazDOod
tevoFzroCf4JAH87eYJknq3ymDRu/yVvZPNfWQqwRm5EvN6yyXbCKOME9GIvBi+C
jmB46FLkKieFqNLVymi23HiaRfQxywAP1mEHBvJ8UM/I7E4AFgihFQlOPgyeRXrv
0fZzP+P8mOtHcymTAP9RMPI9IzhashN+c0pIGjiEquGgNQaFyD75KKeGQUHUtYek
t4d0qcBLS1Rl1r2bqymv/db2eGnYGaDuQpxcVJteDltwMJ1la7lGYDrCrNt1yew0
CqyBFNRbj5VG+8Tqu0bsdd/fwL50cpHCFStZnni/uc0TNIMATI30Al+EvrltsHma
ByOIoCTAY4vofuW+zPxhns4Tc9dODszjska0VC7Ocr5Swjsuqcegk8gEV8qsvaBo
86EVRx46BQiQ5OFaDVzwS6uaf1PYrO0JKDG3Fdxk3XjHsDPuL4+0u12unOCSHvGx
OiV1Rjd5n52o6fokgYt3k+BAvLS9GfF+cnAjNrJKuU/wpSFNIR78GXibZiVx3aLc
bgUYhwnn022kIKBvZvdhckVEPUx1Kp990RlXIgA8Pjb6pIpn9ahK7qpFTvYuJvqO
li3qjPH//5oWedvPERGYqBQGBUpTrwQUQ655XVYNK4HJv50EU28h7W7Ow2PlDx9o
KSL1arma44IQk3TYLOgBzCHYNeUCbchMTKQzFO/9LPbbu39olY/Bd/o1x1Whi/SO
/HvZzubdpqW99eLVOp5Ccm1oU6wlfqXqxztbu/YTlfCLnjU+lcS5cUc6CkgCzuWc
0gLyk3H6zpGKzANFk6nlughDnh1W8cXJlcAkAeTs+/cj1czVl/2zL3XXFxdqkzqu
MltRaBe1Xyypey/XMlD3z2FUiXf4aKGfNZDENZqmNzmo33yP6iX0JJE+VHFzQd8/
H0c92GcsWClKukw4aY1JYquxcgjH4lHh9c5xFonRrQXWn56PseKlUOvv9RsSHE74
4xGZdDxu6uneCfJKLoIWN0EpZeIuvLVcGVuPEDJJ32moYhlMWSIICl6zJRzZKRWg
mpzv3JlF2LW7JLlpUes0e22yVUcyqglvn4/4BcBV3q6rWFVk4qIHMwkoQuroMh+m
snlRtMsA8QpIhBs6uJcFnbNcPucpaDjKjvpOEZK7sQEgNFqiUaJ/4blign6kOkl0
X/JA9aKq+BKL0ZfFUWHofKXdESBNpOevrNXhKh2xSpXiJWeT15L4yXQVD3AqnPV7
qMaUAuCmiHKv8F2Yvk4uV2F/qG5nTFqf78eBtU6ixvymO6ZpoVSlAOG3WjEp+8l1
Vz+Pc0w8et/Nu9ihw1oEmDdXcLGbSVHAVrg7UhhtpYCrI4mMO2Sc6RfSRcTueJv4
3bnqfTKsUmYu9o/yT1sk2xcYEBE+pFIGHmcmiWJd8EclXY8hEBz6DlUxEHeeL66n
hcAQkfpl4YMBoVSHROOdYv9/KkznNP+nc6f+L4MmR80Yi53hTmU5PbSziJ8i8inm
golN0Dm5jkFF0/8gEmL6GBO7oOyu+XZ86lewymN6NCk1T3ljOk4cofQ/DQDajDLQ
UZlQs6DwsTGwID23tXPMqOLF0OqGx9gaZvBDHIKZxvd1rd42dATe+b5u4zcSXy9v
2YrF1y3rDBkA2CtC2+UXYa13+xfEcmwEcbOQkXBH/2blPHqS2GqJWYED3sBpS00t
CsZyk/jgRUNA7fyuevFeWbaFPvycbYz5Z5yo8fPULpJTXXvKoplt7ubd91cvuGL4
3PUZdusy7IvZLr530XuW3R5jJZTwCRqhilhwhi7Vinmz5pSuLRJ2uJt4p444efpE
EHvZ5zDAyhfleJ8dpgk2GiHE3v1ZiYr2yck3Ds6KFHRIO08IU3oU87Koo5CFoZwV
+ZAq3nQBc2pCqdVoqtKlma5wMg8mw+UYcjXHfgxfKF0xJDTcvExwT2bGgyYW/2UN
4U5vThsnX+s/VwvBXCMPL7y8HMlR+a28chz7/SWJ0bLc3PyAMt0ndn0Ap+ukscub
t0CE1KuW//SO6L2QlNI0gk4Mcn4Nc1vdDdEz9diKgQ2w5ud9ku9HyocejAXZAt6J
PkeqHxJOh144XytWTuC2HPC7jQbtbFgzRH0/zXujte5M/3KKYK8nGg9bJzm3mE6B
4B0B/eMz9cI+kNzlk3RMvxA/PeR7dm8NLeiwl54718wgbt/Gs0gdFJvOS3tbZ2By
xOEJTYoDX54Es6Jbn8MQhx9c8BnUEy9jJsYTrUuZMIftJrSV22LxqgLsK1aJwBA9
xlJWqFoNiv2JY/qKqCUBNF4noqCbukANoPRIaUMuLrj+3gmCG0XRJVSC05352EzN
NsKRPEa1sjmUW71WlykfWxlfd+RDBiDd9hBmJzY/j+QY1HcCW3/rleOzBJvvdOeR
JWs3Ntu/t59F3dTbD19+AtBntgicgTkqGr+e3pHVF+0qPhLnS99zhjnrgBDYGmQm
GgUfC9+n8FufNO4f5uCsnvRGcVTvVInsY0Vy0Yq7PFs94Ylogczph5a0Ksv0FpYF
ntibBBm7njE/WLs1aBEabwYTjpe9biaoW/+rArxP+RFSyNUk+BUmY3jFqUhMzMsi
h319GK/PvloCejzo/Xg3TwdlVsh3mNUe0m3721RjaAnZhBC0o5z0zerSeTcugkUe
9+xk6Y1M9Wko0yHgaXDIelzV4DKzRW7ZwSuzlgNwB3it2pXDGH1H2MvbvfY6G9fe
moaAJM536enwGfl2t0iHB0OqhoMxk2pgjOwZkaDu9g0+ZDKL7VDEHEO5eHdv1G1x
S9i+IgY5v9uOJUVtqC2eP0qqD+oJtWp8RFvV6etyBNmcIJrHQRtr1s+/EGQVdm+H
8GR9AY+iWUqElcLYPlt5hCVv0JoawhR/WGUe9FwkKYlxysYZd7DqMU1gOYrbdYXs
ZOwNs2UBobVTECUqJpEWRXvtOS3xIoOXxhq0Xs+oyZZOP11kqdlZCuiFi2LR2KqU
D3lSHsnWClmAwe258XBia21fPxZL4/rilyfm26JA62qNzrq9oOLSx4hfb54/XYCl
3W2WHp2WLVhKt0ciozWcY/2xVRTrBaogJF4C68W1hHvnjEHYwLdvT87nYcY+T9iN
cSYNcA/XxRuQRhDulViC9VZYKS66QjjrEOE8ciNCrRpo06a2uGAJ/nOcCnrR5yR1
RT4OtAxe+tmmfpDwkOOo68glFomXQ1ScebwpVNZtuJInLxjN2rmS4bgH41e7Tc32
sG8lqweq4U5rxM/cqkK3Go7rYBRttQf2peamntq87srC88zngtfdZ3sdXbGdsZn5
DWdE5/+hvissJxFOlG+WaaRCl+s6mGJN3Qx9sv1MJyJEsBu1J45qJo8JswJHY1U6
BIBa4sTXzeN8RdniHI53T1iMkSR6ljltZN/73O+AodnNOquOAG/kYYVwyHfr3/VZ
t96ylJad+tX6r1CtzzS9IT5OWUA36zASwk3e2pVaygOz9qKm7Nr9poHW0v3pEBjs
1OChgcyi+Rxs+XhP+hH1T5RZTUbv/a/5JYOXoqNDNcpA10kHBHBmR5N84E/yg3m0
XDlTc7jONgFxoGYM6ODClOXYwolQlMpancpy2kM4oQ6YD8rd15RJvzg4KHRlSPfX
oPdIHgI8KwGkG4AnW8mlvihsrA2dFKrWdHp7je65r5ht3R6iUSMyFxAu+6P8HP7f
C5LFkfjjwKzVWFQQnnbsJ01pQBRFXWDrClpqoQxObykXQ9t8eKnJNdqgL5xH2dhc
/6FqFc6hmShdUOFSs3H0dKqaC6OFEpxwVwNaO75j+5y9waC2ACBxeWQjlizQIX4I
2p0funBvmWSli8OF2LMKYKntuoB2KedzEj6F4MQwQaldLTXNIJBiIAXjoMVS8y0O
u/7GCndXQDUnVQQKVeAUnHjmZFpFAPS6BFdXGrEKYMVx2c6yKPgCYJcYLzm9zgXe
kAiH2NDt9MvLXqNKd8LSp7urPaa4p9VWSWp3YSGlPNsZBeM5O2D90NO/uLjvenyi
zIa9Zl49NM/Srz3bLTdSHI6X4Hqa9e0//y79U5Nbj5Ib1/nRoWbtZUjs5qsTG8p+
7SC/EpcLgRdXHv0Da6AKkBPeN1K/AMlqT2MMauh4gBUkcO6WwacOiSK/lqrWt+mr
wf7Tb9ZG32yzNMfmNKzKPlFxJMnBYFTvpu9HrIq6Ab3dmgljCTmxZn23Kyw3ZgE6
07ug2yGYc2V9MMJf4Krkld3TQXpxQLOo6U+RxsIUd6Jo/1Joyo9ph1peFeqo9a/h
vz/ZPLKHUP1hXN3B6gnw6C1flLWis0Igx58P+B5O9nsnFhTWRscOTr8XAi/1c1an
VlOxzLQFS053P7jz4hwqvsJKcPMZqH3YJ5VLPGm5vlmKwuHorxKIw3qVVnvq++pj
GP+uk6FpvuI5aaFrKlbnRNkT8fjnC5xc+J77mR+dIp4ApZLoXsYfTwZnPVb0oVcq
q1nHO637+Ic3frFDnxAQmptAW2bccB+SOiO1PreKWGzFZiJXDklWVGTzRz+kpaS6
6kTHsovs64yqKDXLoL5TXkROpNtFYO90zfcXgV2wlxb9uFAXkb8+PNdrq89d5Nps
4f7XLu8QJqm1Z+3LhM38U5waLaUrXs3JL7SubsQuvDKDYYyNVkbTXWtJDayZSTNe
BTpM5zJVbhwxQm+a1L4sNLuAwVf3YoWjNOwHCy1Gjs5KDmekynhyZA2UbbwgaAMu
DIkAnNvpw9vK2zToO4Z5dA+IuYofkKFg0dlvclYtHwU3gSYFcAl23BgT6+nwoIc+
/Z5NaHI3L3aqqJjxbgflSFoOW9BRMpbtOBFS1ScyfkXI9xGJ4jCxrb70NGVXqs7n
C4l2eJj1h1zK9Yb8bs+BvhyMQCnifjwH8dN0njGG7AKsnvM89Dpi1h/nvU2closQ
5T5qsYx3OMrjJdq/6QX9XaEXUxB38CB4rCEaKsFYeIMA3ntdzAiv6IYnOEwUzowM
r/NWu1f98AdL32TwO6WY0LtgIq55PV135XoSkK+HYlOPd9YdYqO75nPEy1QiPNBI
NF6nK0BFEk5Q544Rk7R+d+Mt5+itZ9a6TvJvI6uC+ZI+7cgHxwy0z6+T+lsEGonD
UytlXixkNOSKVMyT5I5e93as+njLWuoAfC/1w6amFr0IaUHJ4sk1/i/DXq2maPel
BmonvSVFonK0fgxhXfcr6BgPxyU97xg7FURrMeFcUZ4JE0k/yaIGexyEUvWyK1qn
nrP+fOe+934JQKKo9cy6pY59MIhsYLicYdSLecTSdE6Dcx2+o79Lp3lp+IbG/lAx
j8K1EPa3C9FTNqobkH5W9lWlsIdCavMf7Waouij7OEMUYoZEjrPI/trDMv4MTill
l1gP+8FunFiuK3Jtyl2m3H0W1XAMveEmRh5Uwz+PRkgCSUQqV92gTGwztlvjUzNj
bFEtHoyqQYMG7Gdm5wNAGrxSWH5aIt027qoxOPWuEeMWsXrS28mPctqn5opyBb6q
lHicCUZIEWFoOcLbGS6e/1QHLKQEBy14Yp25MSBzUja7roFCA0Kd64b6wqmHcCBA
axTAoY9P5lgzl8ECoheY2n8/TCad/pNY9FjZzEvXgakI4vUNIO71sCFvDhg/zN0o
FXStd0hY20wzE1juRMY5U66WxLWUS4BPDgI3IQO2rOehDomGJjsxiSVfPcNxWiYa
LDkPMgp0JO6ERtUXTvwD18NqRsz+0POT8d2gm4ZELpQdY47Gu9KMgT66w5caBj14
Fc7reCFO50gUESGDZ3Fd4JbDGxMHfquLCons1RKjiX2517lnt/U8jvqrLqlIKbvW
4NClrePDwujk7i1dfIST4Sb+vpQmS+9d3F1jMykQt2kQ6vD8mgt/yRRm8yZ2470P
G83ToKGZcLR6Kl7EfwFU0b58Oz65eWSUvsbC/gRq+3bzWMPiS+I0FcvlkxnQqbXl
FeebEMEqdLcsiyVxdUUg3etme9xOytnEDVoXR3W4uyU2KHFTcuwQ72WvlymoK5Tl
HbYhDB5erNmPEZ40488ygjMitB7vrgXVEGfAX0P3nCIyPs7t5Xku3h1L+iFrwLby
z5Pq2JYNiFa3tKvMOvx6NZIX27H1rHWOkBPN6+LP9ywkxnYkRbr181g7hAETKI10
DVxk2WYzBKA32l9+qPI5Ym4Yz3mSbFIejBD6jxoITZaMlhuShyb8VUbkEWqM/s4R
eDXa4E3bKn/Bfk8/+OUKuQCZJEyOll2J/Wic/F8ipF5Wb+N6sKPGnhHLotfa+GuJ
1u5QN65cTk7zvCUMmo7lYXUQB35xHUL795guHWsZzwM8fPAe1Ks1lrL2cXjLzxlE
ZkMgJGXs51WI+rbxKDTGhEFH/4Q4wtDtSu6+0AIj7OQ5WgQrbBctsytP8e0JbrwS
0Z3MFPnbo6eoKZs9n+wQ+51zMf6N+KtPlY1FDVfSNjiwjBkfvmSYHqSwQxqlRaEG
nhl1/5O5VNyG9zR+IpyE2QEScRWbyqzUs2Di0rzhWKDeMVUoHss7JwAMzm9LytVe
fuTpc4qH9B89VPX+oD//Uam3FIFiUPhjGqGahgZhXLmclsbIJbLKq2j2PdROW6+V
EOee62RNPshIElChvmjjDdFPPRd7+8WqvX8Z3lpelGKmi+OG0HsA6jSDZpSGqFPj
UdCLnP2yFpbCx8f4LjzvxlwgE3Ma81I3j9IrPJYgU6QPRNfIg/hWsQTNPA8fn8gX
N84HhDnwA/5vFOyVEbL3ipACHh2YvAdZSW+d0OhwbF2d7MXCQcKzsnJvlbJbVRHP
OYvJ5Tm0C1/5qNPAIcsfSzs3jEM1ERoVQO7yZhrTgmBAkq746oFKjh8umzs5i3Eu
88IPBVntV/ifLB8DqPtl1wFbpboyuMBcbbAyzyiKvzw0pCbUGc5KoS/l4za+qOpF
3GDcWrMxrtDHsltlzuoOs7QmsRhNzLPTN6BJ6VmGle5QC5sE488V0fXdrQA/5MSp
I8h9HbJisxBmr82N2XUHJkT29DSYdO66OBlgbAc06cc+usDAAbvCeZyc8XcKWcs0
ByZPRTqUFjw8j4IK2jGeEzicTOKs/ip1+So6q0iweM1taoYjuL0AvBminp1WH4R8
dHWcP2KrB/4G/dWtxD939YM55iAdfg9jX7rHcQhnkxjgm2goklDuce7YweoaVe8E
VHYFQgag+W3mo1ad+J15e/75qb2iN+YVgH03//kUC0ssIIDGIbTvnBAOZ0Zl9iF4
lxqDxiBbq4VGUxg1besa5Po5+v3DKwv+bLH0ecgbXRng5hGA129d7Mgo5N/x0/yZ
K839WY0Tatt7CjxTCY5grGH8geGxgLtI2HlY/z3B2RRzRh9EcPItYewRkrW3bMLh
/y2lEi6ThriflQzcaEYjD3fLzKUd6zb886QdosEGDOLRzSSp8i5emM1K69Sf1qGy
STtbMyUt2I96E7EfVZM7ZeW6v8dGCkC/WjR6Jh99s0cgRj8Wz/NJtBypH50evEQM
JPG2dvWPE3vhuevGWrzoiyZoz/U0AUSPC1Zbh9GY0P6TP23Bf3riTwUjKrnZoaxM
55ZAbDOutXUlUT/G7+gaGBq4r0A05XvUWjTPqfsPhY4HFp5bIsf1gsG5d3U2/S5G
bH7RKJ8zkz1g1FjJLQZTgPQtSukjR9vkgP8cz3Rg4sqyrvd1UQFVecfZtffbQxOF
IIW0cHd85jlk+oOvEHZSSiDCpWlswzZAf+fANPCegxRaLDucquGyBiLvhDkD2536
fs6TWQgXfikHF287xkQGERZlferyefL6ZJQm/sEkIzJv0GNXpkDMKt4+GjQhVfxG
pqWjZIY6+FenzMKtm/xfna5HaixZn+dM3AxRNaX2bCA/B4zEN2C1ZzQZfuQpqmd3
GWIBprIGswCK19WQlS77vc4LrBldHeEzXT+mndxJ9Y51xOui5Mj3BScuUdQPfYmc
9YmcZkDfZt6illYkcyPAr+hfWaGQtZZPUW9PasyRF7WuwJk3YrQEzZUaVcpV1owA
Hg1HTbxrhdVJoB/iDlUu0UdqWo4eicH82yHgTnw0OtYlTqS8XzYzebIXn05OQTWx
g3D2inv5Jjmde5XNH+LYX6HlQJIYggMfwQOKfbhUzpoyUCKQQzdSTm41+nX4voYl
S1zKPRPXy2iHayBGvA/EjJG5g2yP83Z63VxdEpTKSy0ne7SQHn4wH6CMHY5OBDnu
dgC+EkZMlWpkk2tOFvlw3a1ZSy5HjrT68ICZNdaRnZ/BeLWtAYHmF6dLNapeFr/R
2uvr9p1RDJaHA5ZRAowh3isWW96K1Qs75z3M0gNXW2WHXW9gu6v0GrkLM9pNdeOK
JODyYKiiPgv7Tnb1GrKBlqPIxj42OChYVOirE+bqvpYFSYdiOWs2oQlpOCf10X7f
aHl4fe9buOhYXL7TdmfbCkMbhATD4nKn12FU/vQHCVGnq5X7NHZF227z4UIORZUl
/4ipu6FRrWaKYil1v9HtmmQ7JdivZy/5eSS9l+27zatorlbmNN+uiaDsPfyo4blp
WRNJokApGmh6vJ8yG403olHBWxPWFMJXPLDSIEeGvn13VYucXIbWQFBJ1LZjvttm
yC3YAAkb4m39zZCi6aqEU6RM0qalSPY8QEEO/CTigizTMnv2C9XCduD+cnw6CJrI
woqKSuICKDzmGuAB7vV4UrdA/L3XbU7TzhsqHmequnjVSRO90poWNrZTZOyFMJDO
V4NJUXRG1cZh6x6hdl4bQ8682OeTmvd1nLfAxvodxIpKXtUIhfBiTc2+CrQxSSet
FCj3bp/nkNDB+vg/N/U5WjmjU/mey1/3PJWDqH+evf2YLdqfwe6F7xgZI3/SPYxZ
tetTLPMcZDF7p67chfKJd/Ba3WN9zE8THm8B6jUlooxIUmqENLnqQOIaaApyMKRF
QyC1ryGxoAnkl3n8NT6JfozWmxGgSlhhv8LxynEfYNv2jWkjZtYbXv2W5hOTxCjh
54WSaskeVOwTdA6NPA0T9CyRJjgqh1Y1rwlV3dE7q+BQ41J3BEiu4d6M7MnVegX/
naWqxiMsZSgQL5Cy8+p69ugKn5CFmxiljaQNvSKi6RB+LIrINQdgV1+feJx7aoUe
7lCaElQ62/C225gNyz6geBEdHAiID8HvnwyV2lI0WJpCGx1U3sOl1nGLNDT+TSfZ
uFXUJem09cyOBuC3CmroaeJBiYD5NNCeU6YHF77wSctvDxUshPOEiWh1YEOo7CDg
qN5mDXjlP7PoVwqw7TqsiyMFq9XShygYekO32MdaCWH8zWvdk3OarzD9E4Jtk8wd
Ccb+M+7YfynWcm2P7u/yz+BOvWVW/Sz25M0Pph80ij8UlIYtkoMQ42uqf9rzcNk1
gJuqWtCCpqLngrSP1Pl+tORwTcatmyjkerNNzx89CzOlDjThCi9z9HhIYnrkbq8i
ewEIwrko0pkfIvHaY4iEqxBUUshpsPshx8QdwksN3cVanskIqwC3XOZKsRVFAnM0
J0v/OJnW9A4BKSeh7Cw+8IkUoxIWaqsTQgGVhnV2apb54FEdu3vq9XHE5wRyb4dI
nJTaRduY8SQqOzi01s+at1wwp4/RBirdJ8QvyRmAqXbgqCp3RLko6jmp0yYdaCZG
120kIYpywyE1t1VKlYZBOPMI12OFZrjSwVVARD/+vDkcWQORvUFaYpcDkv929YDl
WI+bHSc4mIWgkSF6o5IhoW+P/a1YW5b120bQoDSnuh0xKQzPCOboHc3VPU4PQIlP
PoEaCWSRt8Bh+V0AIPs3j2LVgNrfOFON/SB2Rn5zZeumatTlq9Uybe+1Jog2Vg+E
/KIpd3TxPg0r92Ww6dTzwf5v8HhtPHwUaxMdbtcWOU2qEgyYpy8RTD6xEGPbQuY+
3FfiFS0qxX/zOnCqhc1IhADR6lfx83jOXAQOHLga/xt6KPsa4WYHGwAiQ/LadARp
vwi5wS7c6Jt9mN6Xvlqv5V93umOwUNBxHXmTlVAWN8FE+mZWwbP+8uxJAY6U7ZKf
RVmqmSa4y8p+qIV/gGr9cryyemfao0AzTKSsTVDlJJ/XS73Iz9OXIMmtSRAkpdGD
SKgOK+7uwgl9nLtL1UwZe8Vx9bJp6f6EosE2egkBQY09zpEU2VlNTsAyfv3xX6pw
uFLNvn+5E5mzljN/Bl/+XrzPY4p2VrR0tDW3RdM8cGUk7PnlUEWNA8U+r+tTLeH5
lDBru26QSyE7QooX8wsLEE0wUcpN1oATkKFakqO6AdsmtAO4gjomcVhTrx8YaxsI
mui+2T5FE2Rsy4a/UGOCiXu6gSicFABdC2xpCLKy0OpA1XJAUuBL9ukyLeUCHAOX
LmxNDL9Hzh7+87D9UOcO6UWM9kZjm4ErA0KNYQXHmNFwcPX9FhgHkpePMOXuWaz2
WYIS4G0VfCI4HuoQbWYPGY0KHat2M6Eef7gWRDSmMBhze+iW8rQOBAEQ6VSskTOQ
Sl+Te2C5yrdxoCLugsiD8f7n7Rf83L+0gXdExaZJbPdR6yPppgkwu+zrnFPX44EH
dy3AjNm+kH1jgwrE2zFX1oPPRP5z7Q83d1ItX+SkMEicot8RkSaNcmwEf1Mqo4wn
MgVkli1ypR1PoGefJfs7iPf1rSGDigBFdDYwAk+7hXVtoKEPpjuZIo68IB6zNAAd
a6I0+LVQUQfLJrHQ1HZ+IKTlOxllS43GMJpGMvLq30oA4m0DCKwMXTmp90PFfApj
MatwDg/wjkhcsafTBuDDyVg7buVG5I9FJc4+cxLRyZfU/Ejthow5rtt9GjEDcsm/
MXFFZZ8YsUnjWomvc11X7Di9kzKl+3TMNUTh4kuOltc6NhgCwD7RRWFlIbXtb1Qu
Bnq/XRL3k2moPSjSpwheYIwRXzsrZyIp5qpqstKPb0h02QvYO3MNSu3Gh2yrAZWd
9krqlgNry5b98gok2ZSnotG2DZEVSUGHHnJSMI0W+Nj5LyqaK37aFZW2kOIo6+fz
hUxygL2k1wn//nvWHpJefDSfT/PNbTZ6BJd8LDahPsfOtZau7XmiF34Nir5gNPnL
juLJig0b6xmZxWfDFjU3OozFDkeyrzVlR+rAc8N/yxjcIIu5HQyF/dKiQYjkHtwV
yW50e03d8XtocHGZBQ1rrM8z9986KO/XIKg7aclp7USlhsZKyB8jlDZqsA1MTtxf
ptqcZWp/mtUNejioh1I1E9YQjSWgkJgzB9F7EFR5s1kdJ2w2x8tZ3uCkN9XaPwHs
vIIT6cuoYd9atXvHtIKGtW7or0MBE9JhONhOrVr4sk3JT9n10Rk8aFv+knTKLu7c
HpvRT6qlUG+2zDhsyHje36twtjl6XIfE5psKqDwuTH3XgxmhEXdFd5K3f6Yi9I5r
EY6Gnz6oRJhcBvgMhAl9BkX4y2OwzFtbsNKsNFBUMNwZS05BwG/KGr2H6o4/yx7Z
fSg6gBpTKB+7Ab3Q/W3gWHl46fVWVWpoe1qJOXxPEEGx0VZhwXvHiQNvFzBgP9sX
eMKat5fM5XJ72ZtDCGn41a4mze0BdscTsbiToDV67Ini+FAe85qkPeFrqxY/kXa+
yTA3rJVdnrKpEgM+TUzhDxrY8nNlLZauGwpqIN7fvYEOubkgPfgbYATGjg8zrI7c
J27VGUNjSLNKnGp/LU4qGO/jfFM/zkB07JY7iQyqvh5iLmVZ06wJ0iW1fbJ7np5w
uaJ98AfecIw0RBrssSklaTrDvkF3cO+MPcZJgNj5ZiKTtCh7uiQEdxYur5BWfxov
af8iAohWcl1z6BikDmEwnBzpwmdD6JyZiAgPf1SV1/fCsEUr79gMoUbW+PfY2pVk
nLS2g1ZgnLemNNOGDqJgMZqzq7cAWg1Czu562mIdun4JZ6ZqxYiSfTYgCrIEhSKj
0AubCH4isgUu9d2OhSvgCTmjtW42FG6FfPURPvMaFEi/rPlTzKWWZ9CF72kYi8oO
awxECcNueTHK1zcv2nQFwSYcG0xUCTwQsn0+HrpTOOGYJGu0SAVK85IICfLAVFvO
YIM1KHNgrdQb65iPKAS7lxdKXGajbMhY6xqToqCik2UYYgCDP5bAKdFRBz0U17U2
h9koEnjkHbqBl3qR2tf7WL35O6irBVxK73+yWZlBoG1QRM8iV3X1ETLUgj4eUYdB
zUwD1I7Vmq0XsWJUYWaAeTN4Nf/k91YXfiGVqGZoec9vzZx3IjFWagESQd5ZR7q9
UlTFEtO4iIfgm00oJnvLRPWbKd3mnBlgianws8Au+IoXrJmbAm7SwpBH0bmdUCYs
n94F1iT3VZKsm1Bc2nhXl867E5os6LhrQzpt2PRbulMvYjSJYZgAUqvuj37lR5Jt
mihQ8/4pxqnPZ/IamCtlC7nmJUC23ecnQZlk9XHON+hhAuzttZ5onIe1JTH5hcW+
D86b7bQHx+kkwPa3WZEKlIU82aqlTjKHR9u1wKm+CU8M9t+7IyjqlB3+FPOu1wCu
gsJK7cNNfzTzNokxc8n+/FT35t3Zqjyj4AyhJyzSFCG+/TkoWSSQ+YODOvY7RBzo
Bn21TpIsvYE2wkI+I/N3cP8oLj3gP64/eqZyIxsinq5ZTcsLXBqlCXnOWPen+kI9
PC0v3VbUcmPWpxzZ8cVopCFieeG11zrjJA98yrDZS96QE38DoGfJ8Xu0/pwbcZRa
BOT7lsLygebE+xHbvHAbLAZDu1/p9knk1rMrzE5LPtMdrx2Qe+RbgFUQ7ZPRKNPc
2dQuepA43oAwEmUp5pQTjugJ8KqQyfa17Lqulc5Y0fUz0hVNho6vFyqsUknsNVYV
cvmJS1qW/G2WNCSkJV0nAcNUlIKn9jUftQy/CRAK4jMfUBvfU7J9QlwRYCeOUIQv
KOYa9ha1U7kCFGgZ0558w60jpateYfaxjC83l6dyVebYQSC3Qb1M8rn/574otc7G
d9K81wweK1JrnMRNank6Fahpr5wFTzpt6KMvxPF8lEA4bmYwiMEmJlSjh4Ohfutg
RMiDuPMPugC6FKqpiIrrnwvOPXJbNWcw/EgETBa3mGDzhiAD2Xd+lR3WdhrUeCMz
1WxFLNNppqEfU5lftZblFdy9tRl5ATR8OV+Rkj/l9fMPS24848x3d42mlAXlPrH9
hBjR9JhsfSQC3W6PuOT9TJNHQVDI13Wt7KqxhTgOkf93DWZf/mcO68Zxu0qv2v6O
f68GCjiXzHkXOaC82IGpiGxJabXJRx885NyPJFjNgS8P3+MjDF04j0oSnC1oK0Ta
C9vRQIvrm3vaUaX6AVClNgNC2yC6aj/GRzmWnrUajUUsHW3rNgpVufmGUaJYgdQI
KY6MVsVteeaVZ+xlau/zCRCDK64XzXKKocbD6q458jhMQIVm7nIb2oKmAu6nbSq2
bqlocN7EazeUPKGmCrtqRaU8EoOFIiYYjaoDzw1uNDQJ5EL7A2JKK9bHaMWa4LUB
Y0+CZmoCDOGH8Zc5As35zbSfSMiFm/12drZIS3D/CGVO0QW2lDvrJU2iWhuuWXUk
Cmp7NPlavQYZp4e8Bx1Ve0OYqI/YzCzQO7qm+pAHg75v1n81b3R0KSUXTVOPnU3m
RFHZs4ddORBAo2nhyDSCrT2UDhNNdK0FuXiBdK9nwVrs3dCKyR++ehfJFpjG5HVI
EEasriAtgcSll/YIT5MS0D8Gssfya7P7yY3cDcMP7S9ZHjUsDin7iPtFrTNbx2hY
UK5vO35oruhrD1WsS8Gr2u8D4ibSB3lLSERbeaoWwPEPp8wUHkqJjGSBHyTQZDBN
JQm3lQbb8qB0KXtYghaPPky1CmZilibvw/40P/QGT0t6bm7fXhVsrPE3Qw6whZyE
J85ng9k3NqxXHJCAo2krr/W0b0gV0cnxRsNlUmj5cTVvVawXZUhFS5Wohpvlsfi8
2RZveKzj5xGaSeUG8P8TpplUtaxiDD09JlnayVc7T/3f51veFmAjKS+F8bn3zSWV
ZoUetpqGkm/juWjjrSk0BYl8/V4FBZhAdBaWk9JvtzVgWTl/0VPOuSRVmdRHUWG/
Tb8M31CDZGO4ThXVmTIWxFYNj+CHK6oVQSJ+2lQSuZp1zg7lFQ8lxbqiBdEaRWbF
lLiYwiru05a+CW+njWPc+TzwJuYJ35vukC5zp4t0ToQCMHlEEbQPOwUimmXhA+28
xKWFH7zKm1S3nhm0npcAQP7svRRPn2UV1Gcy4nqDND36TbGOze02MhQdVOa0Zi5p
lQmgkxJ7W0QSOzYnzzRgTVMImWgiVnzwso5D0t2Tt81Clk6Igq/Qfz7KyMwCElUj
l4jWQkHyvZzZ9WNUahNhvlP3MNUPBsJhx2E/qlE4kaP/Ihtyec1onbzs/ah2j6+p
zsDl7/cnX7vv6lllPmlNjfkVQmT+jRTbKHyKaMAYweUGXe0LSfyZBxeGRrRvAAba
M/eY1wuHrgTLmhbV5GLN0FcXmZ27VmMsWzPH4FkykQDvU95tkEEh5oZ3Y3yHo/fj
Krl7xEFshYcjrEF8Dx5HNqfK63Zl1/nC/Ldb+gCfT5E4gj6i/PV1SzYNwCPn+Sk8
LIesvzWPk/VOYrmXldUIzBh07hzydPp+9HnTHRaKF5MIpUXX6NWaPZYg2gPvOTLM
YObVEGXzKdSpgxNtYvrReE0/FlF8rVb2EtRzTkpoS+FzHrP80w1jv0mpwj9JOw9f
7x2L+gKm9d4MewRtNHjjvw/CDUS4HkPk3975nI+kNQJAKy2ECXiXw/m39gZRQtZU
a1p508swgzppV7crdh26SyrCfvzNmYLDhWwSKUrjiDaK17MyKG9SoOMAQbv5i7ZC
5Ajkdh4n4DuXpfyOrblSQ+Yo9a/sMx+T2A+W1uKz3GjSi8VJTpnk5346u+xNXkZb
hrQk7GHQIMbHoTNsHLogDiPEZLnR5JoX1kKYX8DmEnWhqxTqkheYNtYPpfGesg8U
ZwX2DEnvmULHnRSjNjEiyAi/jxY53lYMFBITE4eFWkeS8FfskMjtUGZWQR5zt6P2
B90jZ82sNgmAEY+R0x9KolgB5LcxqhEbn8s7E76lENBZN9vblj/DB+iaBBhnvhEs
SO84ysWsF9bW3Uyx+CNgBOs9+Q8VZ634+5oSHKBtyn9xvVtc0eepBmmRCeZ1gt7+
r2xCLNK70qCdIrh8VFXB8jbowgRoMaO+CWhouY0xLhaCXaA8Z7eq3s/wAroYlCr2
2ccAXD+j6blgXgtW/M3ePGBph92FSBt1KGybgDq8dkgSeCvG8yAJoPIqxuw9LCod
qffgI4AHHcRDa8IE+HFOeJ8wefN7+ySZWq2oGX6IIbS1uDD4tu/DGuROGMAWViSu
sAN4F0uh4smHA3XcL75r9xPzvj1QetXQ78WpwwcgfjeRfdfIdJKDldLCTXNiqHwX
057g/eouEuWIR+ZzLGqoRrFhlZOEvOGEm+zYRDZD35LGYrPBlEfukfKpX5gMvPaC
sUAEG15pNZ7IVSiYLf9h62zHPoM7T641Wy0/3uRKTAQgnDG5v+oGUz78lkctPjV1
WY64qKI/C/r4tTqnFrvJxGjsSDuJT4jkfeGo8NY1i8W7hDb55cbVW/dofuR00Z7G
49xgz+NOvz2erEA9z83zwZg3ID1x9ZwZQxO1yAoH/UHoRM2WBEGiYpEpP6Qunvin
oyGN5dp0z+7KubNhBlAqxs1W5EYRzI4pY8VGZadbG4Nb05SaFeIdStAfEIYD/Er/
SS/Uv0oxQVlWbO2UZT7Y95oejR2yVb38gwjZsnlhXMy4KVT58vYjmU5KbtyIyhbF
SR1Bw1JlvKiYQOsmaAvJto4qXcFF0VZxw+WiqjyplryQ3Mw05vj/CRRYouQJWfD4
d9z7fA/I7Equ3BX491DPtrLGCezxQ3a5TJH8HXy1hhQQoak+tTi0RYaiekkFl8q4
YeKo9tY3VYEHAcKlco0H0lhBsMuuwmYwzvS0Qo5RlW8k/HXolO5Cr2nTd4d2Su4X
W6t9UAKkoHoIw6cxyXMjEE2JrLkqk1/oiQKXctMNSiOVR5MFAJbNYw4rbfctoQmv
tcuy/h0Ozc0nOg2jfzF4lKVI7J6lKyLoFtXond+VPUbMEY5QxElDrMCT30ZwfSVr
LRoDccK1sGy4PLM1QumgMRSyxx8gfwc2xKVyBnG2eXDANtovg8sJJGxDAiiPejkl
iCiLdzDcgEmIgQ8Jo7GPZHzOrNYl52rYyAbZ5iMGyZDVtkHbP+b8/erJzNP+eKRm
9PYSxcYy1rnUOrJnvW3ZRxw66ILhsPklpmAFED3WzhBH+m80T1UPRHdaX2c9CgGt
IXGT9uzpOQQTCm8rzxkIBrkuxpAlqg9ra6PU7DBSWfRm/nvu4a5GIx6FA1ZAbqVb
knOyv4farkItamtBZFMAgrnt7JxRCC/GvLr42wzOJ2g+wkiOnvuZZ19ADh9YHGJ7
g1eAf3AMKJPOfFkB6SRkfFf/GkZ7PpAnAjsBx608r2aFLIM2K1d6Ucv9q6cIvW+1
VGF2domdDIwC+hPj816ERtHOZ8b79d9CwQnU4O3pthrma2NzkuvidABPt1GPwVIB
b50j1pxX9ncXggmzoVZ5tkwIAjF7pn+gI8l6K4iCkXYm0hiHEV7tigezc0vOTdrE
YgdYcPtl+T0MRrkOJYFpqTC/LMDHb+LQhQ6lcbSxFoaDoRINf012XMvfA/Xltbi7
Y7VSxM5zB2bSbNpKm6l9j0kQxpZKea1/kLfIHcuqg1TmxB5rJN5LUoqDzxFyL/9N
VLNj7w3l0XDkTcoeqg8IBh+y8bajmr6XXwVVTUXI2BBBB787exzpiiBKNWEUPPIo
WwQjnv1QzyzNXfGo162iaCys4mFhjekjtu+Ovho68hL91NjkC7daENQqYDW7h5eD
4IzdQLXxaaZjnQE8RxFV9h6SrejOYJ8zE1ae0rxoBcaB4uHU1AwYdpFKLhQGI6bG
fKeSTaoDUR+OoDQSSnPe+JHNg7fm54TJTYtvcgOqf+MBliyjJAxxNi5utT2fcN8M
sm+453ymnONyON3dk70wbUuKgvULc4AuTdlEPbRk/QiOmTtNMTDEBEMrKM8Y2gPy
u6LL8arHH8wtlwV8GKPm2OQZhJcJyP97UWJ8c/margKLuupcnQGUfxZ7+fr82inP
rqAhnDeIh8ke670vb0Jm1rGRLIhuqEVZ6FWJe9bZwgoRaCyY2y4JzTAqn3yEdihR
/fiS2dYAgI4g02MDdXrKi/7U1vHm2ZB1MZB5/RRUsZj/V0jkwDoP/UvskrmW/6BB
MbfvFCbWQs1KciEGoAGmHrPE+hZXZA2mRI8RLyO01LXQsf1/x3c9HkiNoctgzyQg
Q3iaAiPNoxPHZSc00yB9KSyxOU7vEcSc+k7v3mElTprNoQjy6OUdItyCvPLLvnle
HB+yz11l8Q2JA/xoCx6MwXpFMYbsRVpClB9N3kvmTA1dcusue2TZ4hHTTf50PDCV
/j+DieznHYyeY7ivUWJKZ8IbSbnVbPOI1X6sTieOkI52II6l+vQAi5U9P0+GIrWg
/4VMBr7Mk0mIrAGvp1RDgJWo4W+w+KgZM/Va7OHZXI0FKZDsGPegix+AiKEZc/FF
tEo1yCS+BjGeY6oerrDT7FSUQfe9xtyrAIOeZB7BDfy+89mBXdJeHL0CFz9ZNyoQ
lHclggm61FvVCE3m/wk+EDhFDn78VlOnap62NDPRjOItIqmDpHCYEBS18QCLUU0U
6v9pwijLw3/6KCsRMD6kP8zkt18dXk/V0riTCCbZC+qENMa5VIoYmnwmJdw3ok+X
iTWuUFUvNYv+LBSY+HbMJfEkfSyuzer3HVpQVtO88PTLRcdkeVTaDaRWtu8Idn/n
sDt9BioEMt3+XP/GhaWWSSOWI2p4qpe6iHJrhRXwEoN7/q6tLLs/CgSrZJ+R/s0E
Jeuiw7WwjhblbJagdAPAdpxhI405EnUhFzlowqxZmr8ekb/OtMQUNPWrY0NiISkB
LLQeJuw7/kwdUbwE5u/iRZ6fVXGvmetM0YTGvlSw7KQTFs4XOMwG3B/BNjk8tK0T
g7ey34dMcKU1us7hBDxwvaLaYEoPJ01k4s7M2bX6g93ubCc+fjwKlxbtckD2F2Ml
vyAl4JYqc0j0sC5gtNVjREzNHJdfnOgRo7N2HW9wsux7/Lst3Drwt0gw/1yQuzFk
2oZ+pIxJYrhn4knKhtBiHzQNLqaJb6E5yWFkjsjxS7gG3u6idjyOnWpfI63aJRtj
aRcnej/TleTtwwDyoc58yQcu7ph27d/uTvClbVBOQmYkqmhiCQVLHUfY6c3LkxWR
BVO5OSrDQVb3qgzX5P9p4hy6f6YuEKIS0VOJAldBhLxj/4uzIIJoXkuFdg81V3Xx
1cuJf4tdBJJpwHmh/uAHIsqZjywqFmUX463MACudjGh65e1ZREIZ7K7qk6M2wFt1
kSe/GVORJ2Erzgjiw7uB9HV/0iBQjkk6CChi1UA/y6qqdWvx0lhhgzg8highFVFK
27mmiqykqEWrX0hIZLhBWkEyid5o/SNj//J1YlgnW3GmX0v6zLCwSXmCZWJpsYBO
kCgdX1Bpv3Qqgv2MoVykL4gdtJK3lg3LGVSHteXTF0o+rUds5fFdIT8Id8jPQsCH
a5177ilHaG9+Ppw5VIaldJlVMk6cu0OAPDYQytr5wpnRVDXD7byHPNF8anOzruHR
IhCzGf2/equX9C/281rmPr48MWNiuMIUNCQKUsgHYw/RSHYdgo47UCvxPkuT03G1
GF46d7Aj3hzR1khpg4ZaM8uTdYbeUYiIjETpLSei9ZoVIkMq3tbW+/F87NkWrnJT
Is37huK44d7unPFoN8S9kNpgB3ucqjf30P4X4tUUbkMULv8Z11vCnQ7hyjL+iTo6
l/rf/8l4a2L4Z/OJV9H7rn3HirjPCWsGS9HsJk+Z8ij8dYEWLg0A/Oh/FVUXEEGU
MdKGPTIUhYnirjiCJiUTefIDvk9Qui0tlgMlvO4Xv7Qm/HmgyCHjw8//MklJpIWc
nex04KQOBlcXOEfQTyMV/379krDu4GB9zIfqxzcQpBCAbNzF8m3KbWH50im8IlJ5
FBD/cfZQImw/9V7TdsMb3FK3lOas7KvRduK3kl/ljJV9htPEveLPusmmEWE9bhj7
t0NTpnngmUH2VYA9mv6vMzIT5VM7K7qtTsZ0lfo+dB+yqgdrV+zjA6igSz1et3Ih
21OR3Fro2ut/Nd92TEr808c0FfWh0AUTu0ea9+ZKDXHXalY6NIZwvYK9YTWdCQCH
sThDrhJV44mPDgUx31dvm6qSqUkq/UfYsEP9Hu459wSDv6P6VrJIe+mxaqxrf3Py
V3tirbu5GgjWzVQklW5Xp62G2aH6xMrtLUXQXaIbpaD1+bERIJ2RY/lPQ2cz+RP4
D+0oWMudb3t1SxQxZ9ixDIplptbaRNFH5MujoLrkOOvlvSsGybMFz2vlEx7XiR0B
SEhiXPki+I9vCcVsqqbPfOfTTbCShosbriBXXH4X8LgEwxyhfCbrwr+PnsAu8Xgq
RGSC+1du9/amHs6LHjVMbFtYl72BxNSv8lKcwpD+jODWmCydbiEpzyqUcOVPFkZu
qcjJTFI9O1686+WxYcp1YDUxRB+oXKYTLbNxgLt2TB2rafbAtm7CGqZp77+iFYud
zXr28XigrwAGmEauTKy9HCNeQ1xaifsxdM9+w8YGI8/N9uubqAa/JQ9A2pIjjIDT
ikgzpVf2IQ87b10G7W5rk56yBIRAhASXLe6AsotlbWjBUjHCaLqj11X/QFgiJb8g
WnbwTn88VCvuv47+AgnhP9nCuywo3Nka3blGsyWsh7P0Ky4o/k1BDJ3m8owakUPY
IBu/jF3d6kdlVdYy+DzrJDC9DF3pBsUmMcnsoVEOT5uZ5IXfTj9irrx6pd5vqI4m
I0Z8JKfBtxYWpTyeyzZkj8DfH67WppwLHLrAw/ukszaEFUnZJEUbYk1F1xd33rxw
0XoKcniNX8tT5OcjEsqTx8gLwBMkcmzZZP+5/r+YpDSSYSGa3Ao2wkj9dlBtY13z
vuY6Gh4oH7Wn9d2+A29HkyXWfaAseVnUUBCLgxoCz1aEbwF98rLJYzBrFslFULOe
Sc9u8OXIb3cnVXUnXyAo/LsP29GXLTGDDEBov3h+Lj5SrC2q+1c31JlwNq6YA1w1
+O5LzgeY1qThGZfTwhIwZH3+lRwZ5A+7kNeJA0JGUFLQv6+QYZCmgSyLfJ2DfyvA
xZcFIvMhpoxmQozpsM3ee26bEikByNGCZqFccjjdIicMc8/dUdAVIfvpBhk6Uhy6
gLi8QxS17ysmWvplSrw8A4MicqnkYRZorScXxtVjX46wz7jLToG17MryeXt324mp
YnBQfS/o4iPxJqoWFJ4s/kAqhGKS4gYNwaJ7uPJVEGXo8R+ssD+yLX+rGO9KzCs4
+4VcWxkHI/vk9SN+HfV44fYrZRD05IjDxmCcQtvPan3D/mqj3UzsYSHF4ikKA8hI
iPlZ39EUxB8zKBSscUXT+ggv4HEvhBcqNXZUl48CraczR5mzFNVlWTcN9ZmfdUIs
Ck9s6+EdFlVPHxuTgB38NBUxs5iS4etRpMEM7B8rkEPzdl8u01PKOABq/HUA+MaK
6IJuNiEQjw4f5OMZU/Q/RvlPk/H8c/fp7vDv1+CsW82ktsgPGeMkd6bWNg0xq4j5
Rk2pCTHFnapOvYaV+IYV15iFrPk1E0x7sCVeFBdm8ig5LHwzMpuAkwkoKdo1qmOk
mPZZlB8bhpBhh5qZ8P/LaBfy+y0YH2CKG/vJt6nf0Fw3kWD2POjQqBdqmqDSEkKx
7X5W0xePuH1vtYKBZT01am/VeWC1mfvqD5f/sd834zr9NLVaWS1PzMBCINaQBvo7
uotrOofY3sWnBK/DIvq5swyzBlGfVSPJKdo9s23T+TGxd2G+Hr7U2rXOxdnz7zSt
QoVsQObOlzyTzfYbhLTsRcqiM9URjMR+kikop+jkQeXAjHXVSdxMUoRL35qtwgNF
GsxjXkgXe3FPaxAopnSuXXDnNqRxsa3isvNSwfe53zwF5cveqsQGdumRKUOGuSdS
kD3kvKGqZBoPypdXVq6PG0UCeqxbwDvj2eUTOSGcviawX4Ooz7b4XN9dFRlbhGcL
wPjvAhJV9wCCH1P2oOBmCHPhKmDxW4ctcapQAMX95W4LPI4J9u1sjQ6esi7aBaS6
Pl49yk57sOF5uTFnKkAOodiSt+qRECYF6P9c0kuLnNhHihqGWuDwgB9KkY+p0sMY
mggYm+NIyIYmsghtkVtqSLHzYd04BDLrje2JZ4munHT4hJenvDhqQSyHHVGNqwDu
7i7EeBlVKOKQz/Vhz3Evvvl8/JLDVwzAY3n+n/aNWlMBACtPPoOxTE4SsW5qj45q
6egvW09afY6eXbG5I450JyRAXMPQDfIKIKMZLJOPKyGlIzQlDCpEULeGhx9ZYMsA
xcaTJwwBhGY1FDZI8ilG3In7g8CL7KZm7he8wCvpryZZwmk1uystEG7a7lWpwBsH
PosC9v/ck2pmkPANIAvohm96SKzYwbw7a+1T4DSeA3glh9CrSu/K8s2Lba1y1JN3
+oPflW8ZqroXn/eqJG1Lfv2BEz8fc4ZGiwa5ewrzUx+sFuAAAnqTRWtmPO53EDhD
zGzoGs+gvvcVCYl6LJjmUgGlEIWY3RxVGIUbSoOsHXIyoCaZ0Wpot9pu1k4tCa6W
Yelf5fV6RbTjwRrLaAJIZLzW4I2vKxYnctwgtMHCfGqnNE69vUJSoG10YmQWy0/V
UsQR42hOn5W9PaekgQARj9Rpuc4rtx9OExPlwIh4PTL8ksIqJsGBN3G5OHw0t3T+
Dngc9SjwehGaVa4cS9JFDHZP+L3L75CBxhfMI2hw1ej0bMhKg76m45fbhJ7Ou3ly
tpqXbRBd+8rGEi0tjl1sZrpm2b4Gnv63LSNaPD1uAqcIY/KAw7wHds2Ymk9Genxt
QaILw8WyF0xdWaXpT9xEUmTnNrqmSQpKKBz2bJ7hvO37fKBQbeNL2jWR2CSA6Opt
XrZVlVufZvIpP9fie1mvgIfnxRq9uu73wVa8NEei/8emjdv0W+MHO9BITiEtbGnR
WfZZzDG7np22qszofdlmrMR2GX76dVShO3ydRxJ4MspqFRsDKo9gq+zeBSsY/Vpn
r2IeSrC4Juata/0cnT9QSiKfip8r9u+g7PLu78oJBzYU4WW/fFJszW9WIQEe3XSd
gtG+Q/qTD+pbVGyL7y7g2kAgbTpOxo8azI4k6mIIpDSobetW4U/8jqjJmXDiCpXN
PmJt4WCBwTwKvraBI2QV2J6CILmKVDkdm2/eIkWkFQ3cjQ94wt7XRIxMqN4gYK0e
WSocFmnVGiAOW2hjL3h45fIax12BKAXCmgrhlYRGyjOZmEALoIRgfPYhpirLIiZ1
XMAXexf+gTf1gK/YRzLzeQF2g6Vbp6InZ7jU/KqdcQCYFIxr5XUwyLLQVYeNfyh7
Wif6K6emgDLzU/2587SGAiA7qbTh7HioNYW3xBw51YSthDSQJgmyYZUl+rR8EKWG
bEkUuNDc+kFh8DlixiCrlmRLwiNBKS9yUskqAmkILIkftI4A7Nj9zDQlK5tigzUK
YaFKPPlwd7fj0Gw7nrC1KaOjgsSFPUJpgGLrRXLoeabS6EBxhH3O9FTwRWs+PcdZ
mtzYkrazddFjiCj6RPOvAOYmXSZjxbzBEhQ4Ys3EjuOlPAh0zWIxO43DcINEcsnP
sAsHMy3sxtGsIus8IBB/Tvp3tJNyhelKg8GdAtvTF4RSqYq95teiul7ICDc67wgi
gXSeC1IT+Kik6+S4W/AtE5SdQpeoum+btZDn4Qz6+g7OT6AS/1gdSr2iL8is+1rV
M6e2lDw6JCw+TcvuJNp55YF9e2kt1/S7MsoTLGkN5ulI0zrjA8U0XT/gXO//IwTz
yDjlzGE+V0ekug1cfkc9vWVoV58LQdFw1wT5JDc8f66/c2r06VuW+Gwl02L1VBHS
QGbVRWFljPG8ErNRQ3jZMKg1nGFeK3NP3kvQkVpmVqG1N15H++trNceXB5oNExq4
hQfP1vAYUBls+EzMAVLpnRlADQZOr3Pgy6g6wMx+1DDFT3N2nW4uDowbwzWX6VQe
7echdccKIcWMobxJM63tP0vg6AweMrVjttuaqap8fD+LejZuk/VMV+i/6uP86jY0
fXZtbxMgyxG4Th2paopl6s2fBeWnwV+4RadN/R9XY0f8yILy9o8XiYc8iDrV/Ct4
RzYpOxBm+yIf5jE1vkMHiQjP2R3rde6k7TzUZ1In0kA5hmpW2ZwLJ3Qb2/1hV7jt
5brGcI1wrlZA0hw+YWu6ZlXb1wuJ744HcjbCnrfHM3SZ3+ktLUi1B688JDf/VlfT
8P/N7LZ4i4rQBEMQGu4TtUcr9yw1/sccbVMpE5bBD4ZprZ6biQXT6xmhuH8ZwsUn
ALassFY8P+K56/mhBT8Xv2cK49vz9izwplAOA2A6uuHgeYK917Nj08ABub5vG+sJ
HlNOR+NcTZGWFKFdtZKqeG1dt8HXWoqtnVd4I3cIIZop7gOF3TcyL9yl/bW+90oy
XNf16RUrqk6B2vQUnwY4Sn3O4ia0Hi9hQvUewjZE23YOix2Jyqk3u8ThU1C7eOK2
29ZL82cIs0PTS5fkLMSKtk1qe8mg2LdtvxNrMgMfxaCUKroNOInk0gM6Hd8WgTEp
ucKfA2BQnt3JPYhNSeAcua8ZMbr/cgHIdD9GSbYawyilIdNGmVYiWe5P0Wm8VCCG
CII3uqJ362XBut/pRv0MK1xN3gSb2Hu/6pBaK4l4LEcoPzJggKcUH2uCIdqnOYll
KdohVrQY1C8o12ao/WUXlUV4738SafVYxax9by5tTV4XZJP7TNKZwTX/fep9LWgP
4ucOh/R/3kS3gtvOR4nFgVRqiAzUrEYcq8HgpqrJp3aw9MfpbpU2A4kQU8n905Ai
qX2bKzkRHspA63yumVPmCm/EAW3l2nuv/FuFWXdgHuIEag8Z0SBQ6lHTeIMjlKpr
x5K6GQtna9zhfCkh1LW2bTYOLmvr3DAPZyZKLpcccRbcKvbndqnhnkOipPUjUaZd
yIuWUx4J0HRO9/Tnfaf+Q54yz2FuIBI+IbFPDW048Fo76z5H7tYWUCy1e3ZaGyBE
C4+MjuY16Z5iZxnSuHvMGG5eYGb/eQctMHzCbXbYiKXp90KMoRxuaVn2uD/YphIx
FX0YS+Lxf8n46oIjb/qWPPrr3ZtY69390hkBb3Uk7jZuFGW4qZNOrLGHv/nLgQVO
wf32AMvAYZyoRo0HW+DlcXfV19HovhHmhORtEVjWvO9Hf3x/4V8emhhObL4x1Ip3
1wkNwHEhGYJeRSV9Mc613u4EfF2dDiHON8futxC4A5E7hGDZD3C5UAQH7vd0yhFH
bU4IHE52x7oo1A30I3fwfHy2n9KZcGx5xaQfr4r2Oo2f51coFAxDCyyJuZ+pQE5v
wZSRrfl7HaL67JR3y9YpW2R9RVILSyYihz4It1Amms+GUEObFl5dSSPS0lpkbwMA
sL8o9WBXV+FTLy3tqL5fgufNCADxcvBqEvWe7Js3crw83VcxVsCTZp11gExm8Sz1
FC7Q342Gf//KInoDMlcGcALyyQtYGfqhfHYSUvTYR9ayrnDUv8nZOS/AbZ9CK9Me
AKTEGNsUUwJow+uAmHVglruNfCIZI4LAvzVYFnDNJJ3CukYJsX5KCUtiFepxzWyd
sWNE4HJtYCeisxcpjrEh39qUL072aE3oLORLIUqoFEjCZJ0xQaii2f1xeQKoiuPO
7YdNPC0uv7N4iX8U3x9wf3FgVXwnGTYca9o0fb1322U4cXMnmUcKvqlve4Zrh2/i
0f/S7ubUOg/wCEMZUXHIiloBvdaNgxdLx+gTTa6WTzkPRVgxG24edYQz67uLz+QP
QM3yCywWDrQa/tRTRHlXASm79aienOV2APiRhP9or7IgJXQVrQ8Bi4jiBXl/vQvQ
Cv02LcBSIZpgMeE/LW/9pQxsvHYMTLHuysRztTi7tZau3uMl2Mf9zBuwZrTJLLNe
MoXTJcO72h9Ww+9/7n3peHBOpOUKl1l5wKodbDvORqwpLryp2VO69KyceclEW2oP
ib7h+GnMWaSAo8FQxI1uCcp3z9sSyPytPs2b/bmZHTFP01VGWgglW5MXyOElKsrv
rnILg11SWLn4BX0uYB4e+oAKjpsOWMgUnKIAd/uA0plVn8Vp6e9WCHSE8srlmJmA
+VShhquXHDL7hKPu6vgZtEup+kXmi0qGES/lexSk2JjlSFMuR04JgIzSsitkcNzc
5ZmRiRto7KtBIDej4wZdQrKxuhK7YFGrjfhgMam9rPdiIl2Zk7TPu+gmsFrHMFRY
Zg68Nfn9zCwa6ebYRf/mU+jV6dEDqhawi3WDO7Scl51If4wUjeEYHmCw/quhE8EF
RtcC76zj1E/R+dpx7ODXBQP/68P04wuCDcvWPLErMZZWbYjUewG0r1+IAgHg6yBN
NztGI42RgntOh9L6NBOYy5rGKzWbwfydD2GnOg1NfWeM61vnLq5vyg6Ab/6C1ASk
GUhMpUIPHl/oLFYxyCn87hhWdFYdWtXFtf6/1KvY/xVwrEqdKpohQQvWS4DCFCkN
RUe8iLMZph7JAwAozOT3S+9ZsUDNdgNUeqyDal3EZ6R4hCowcJJ0CAXW91E614XA
k7UTgs35QOK8ihG6Lacs0X+zQHjPjJfGMwN25bwaTDPDraWL/LNhZp/a0eJU3lI4
+X8se6FF3pLcWK3aSbz5JOwDJyvsjTo3pZft/bVkKJPnZiybYIEGkRMJP/5rvvXK
2Q94BmX1pOmQtQkPRs0aQlV13fYJHVkO+0VTy9UtBTrvykPX8V7QHsW3ApByI7P6
luetNK7UmvIaVRPAT50YF4P88f0sJhTG5dCeUex3TK89wwQF21nvnVWTgf/HBXkg
/9hPehLDFziyJ9Lif7lwArToz01xAQdJrxV1mjDJuUHPWBpiWmHW7whrJOlcRw9D
S5ngA+N0TJJE1liB1RnmFroqFBsNpTNFc2Mp++yi7PoNIlGfBBaMZv7LkSfwsLbl
mC14EwVDlL17QXaBZtzLrgGQJb70LTtHyg7y3d5PMvL5wWpdY03YVSIAnr+mVDf1
RpkyK0EK1JO0O1VOPxsWOb0gMkwz4EQUnPlZNCby9WFKI+RnIGuN6aoLMtTAhSGX
XmfECJJGTEendVzEAx//IMpzqkWpTstHm6rBnQDHRXbWLh4bbdq9kBLLfzuN3Gsh
H1IiIXxtapYcDLC3npr8gzFmVhZEi6iqHo7blWYpCkhP8TRzCdLQ6871ddnvmB3I
b1ldPd4F8CFV/FmBLKs3+luspvTuaZErb5bok17uGwrr5hKMMIuter31BjNaaKo0
6gzKnn154S05uBc2596wyby2VBvria9YMIFnLAcO2PzpCqtfFFD2D/SqU0Eo0Bl4
x86GQI+v628BBNvRWpWlD8/cDBZq0S7nqCNglFBmStOarVe+p+UmBhFTsB3n85Nt
qlz9U3o5Za0pLg9u6QsalVibZTRDb8v8VZQpHZE0VcH78NCo34hmZE6zXPpDsm9N
fNgStlxxFkt+P+rkg64FnUaVECeRIgB7nuTbrNQkqmXvAxCl3Phc9D65diLUc+7N
X0yW5in/4IH8UabX7mh3iv+RVeZY0RWkONWHQCEatxCN2LJkytHT0IWkaBXy2gI4
ZnSEvxHg/HtBJKfEpDZaUDGcIfNhWUtGi5Ad4ouDnUkQcIjSxinUvccqBCk0tHqJ
5dRevO8YAQNnH7sQX51OpIZPrevU0t176/O8QCd4n7StaQivCKoH7Q5rPBj1Y0pL
mZpi4Z/CqRzsQC5s+fTEmIshcJBkbiFmZQkBPeIRjb6ZCqlyNsm8bOowCMBSJP1o
oNpZXtuxqZdi+3ezHB6D1+sVteLhwtgjjJOkaXfZh5p0ej8LHP1c6LsxSsSOMwZc
MEmlc4YfHDanpFIg00qq5qVwgbMyAnM+88/kkA1TBQote83M8mC+XnxsT6iNIdlQ
NzEsMj4R0PcuDKIttrgD83y49G8VrzZasToJ9anRuw5uvvdbOzLhLp7zqglZe2vR
r/ix+PvVbood1MDEbwcHnPf46JH9MtVWLEQk2v2XVA/F+Dhfc/GfYyrJ7cRnE3RP
OK/ZHc1lo+MY2ID0lk4/gTDQT0yIjIuHExjho5nEqSNuHm5Qfj1RSMasvUZIDDFF
jsS1AaSK9hHaD5A+GygbkEGNdwKCu9ZNuQmeN4rKXDbQITyiLvpnE/Sh5b2dfXK8
Aq6oniYiet1KdEESwzRmx2QmurFrl1MHQZciB/3Fbwf2MrDLGk0qbXv3KveZotcX
GFror9Tb9fhTlI/xusXk8Z6MoVaIW6xQcz76YRu5ZwMcCP/agX3FOVcVU7PV0v3d
F3T7etwJZL5uENp749WYQNtpnf7R1/maiyrxNLfoTyn2IUd+7SWVQKQH52Wla6tF
+IZAn7vD5iLnwfWHQ84v4FuXhK0JTDnqyxpaIpVM06+VjEWuINufLaS5VX+X5/2t
zJ/SOF1pFCkBg11P/jT05tNw0bD+Iul5WnhVbXs+19BG/9Y+Oj1hzh7PtVF79uLS
M25lC5R0qEmdV5bwrSRt4Wg/oVF/4mPOktZ65NjFIbF9ZP46bIMbmTVgzknu5Ova
RsvNcceO+LVd0FTnqBf8gDI4yBkzXX0ZQu4BDNvPIv8SmrqMkCatljMNGLyssOUD
t9CFVjVjAvDlCTcOffVPpDiiO7yL2SwtFH4HKiyCSM8P6VDaeEvLUaans9eoVAEz
Qxcpsh2mnnkZDUDzAaq8vvLwSHcOsJpQYWDsDAYM6qud8Et6TJqqY5DEvfNnyoHp
Rn5z2/8UBnB5HDGZu0WHO+0Ou8aLvOeQ9jLvgU26UMVuL0vZsBcmW7gMliGvmOmE
8pnxry9wBmMnm24+6r+TRrEyW7El7qy1JPIk1Z58+HXoqMd+81+c3kUuRhO1N03b
4W2KM9U7oR5yD9LqGABSpR6Cd3C4C6Pu/widW7JyJGQ2xGyrgGaRB6H6ASLTtfOO
pgA/8oX0gMA2/iVYelqSVgOuwdCVwf6xScoKIQZdBXsB/nLXDDe0Clj+nKlKUBYu
a0B8839VCTHFUQuy1BNWxo0kwffLVR+XqmMYcyIisQR+lv82aiPj1ikBRA/DMLjV
Eib906F1id4k7F59Bz/ULAF2/Am8X4AyISU+zwKbw0YLt4Eswd/P1xuZXLAGXZ7b
NuMcc1g9oBa+tzINAaX43i5p8WbfhEH5IKovzrqWFQobsAIdDlT+oBF/Wmzk4CBq
segtcbzsmJWBKkaDxoN1vIV0w02L9eReTrpcjRsm3FInGM+vHvoXqSPqLhQwhXtD
DAfT7ClJlWJRqoKWBq/Rk4Dpq9udIKIPXJ4Eq9HKrBDskeDukvcQlmrwhzECytOh
w1cn7oBn+FPxLdGVeP0kWb6rLcUsk2AWApPWPm1hd5GVWRM92EuUxG8UvlGZ8l+L
Fm5qlHtpq7T4W7D7TdoiJ+zgD1xI2T+OUSLYPD2oDMhhns/6mQ4ggPCT2TdyHP/p
eHMLh67Drfe6oSg0vZfYvHI4y3H7suHE9zeIFcBoidC+TuRlFDHPaQ/x8VEEXP4m
q6y7G0gycwKGDXK18xUBWEWKiG98fBWhZTcXwZrtUo2TLbdr4yCdIB37h/sIFS2c
67kDUo6aKaABruG08FeuFlMPsMRWei6mspjJEfd1hWfpmqI/lAl3P9u3v+Moe5qi
zzIUaNIbjhUAvghHdNvRigsJTUXEFrRtZ6NtmOIKnRahmc2qL4UA5Lg79VqWvixU
31cl/pfcTT3zL7Uy76sqledlii04PPXf2aiNi/j8EGpkcZYLtFKkjzDxHSG5wpgP
IprL1dGg6XwXtriCiyEKa0lpd85odN+G/TDueWnKUR185eSph/BfL3G7eaR0hhl+
ODSCk87cW8hzHd6nFiomdSEahiRsKEbyBy1gIWL2noEhih0XCxdTjb3IQpFHl9A+
BCWhSa8Gtfjf8YI1aXnx2tx1EMGnul/dwzN/94VLlFmY0RRXPxB5FL+fAL90veTw
yAY2kgrWzqJPJEMG0ueVmZMP5oSSHqgZPFeLi5Ncx2yjd1pOjDNHtDxHa13T3bSp
pXYGIpAH2uejeSQTb00mk1xI9HVaJ3jC1RLtvKENx10R1qvdm9bDiihZiL35fZtC
98DnWj5v/LHxofnbIB/KJ5+6aIeB17+mcMh/oU1JCuu7qwyI6ImcYfwuAlxsQli9
c+O+uF/xtBMf931GdXZCa9ToOpbWjvbaPypgZ2mylcQPoWxtibe1raWpV3j+Pdvv
D61wEzk7miXaQO3hVaY8W8tCS2NjUosj0CHp+rtADwuwHV+hSiOqG5d6Jhu4nM0P
mEouBsOYoJ+P/HsOm3VIt/ydTpDvBbrXIeQTReqzlzk0rX836pRg9CxHOmFpiSjp
EpldjTvJzTU/aftjQvNLGCcNGDcY3qfIjG1ZBTL7SfY1IKcK2A6PMu745qi5rgRL
j72hQ6q0ra3Yr3pxOW/WR+413HUtmZCJwMyQebpaYRCRD+GA+x5jcieeuty0tucM
GbHSn3lhBj0cMr++KAh1D0/1HxjqkSNrM1UNiiJLUdvBHNoWuTBMucEywYIyiH3Q
QeAmDpBT6j4qmefUwPKK7C9oLg/FMBLWpmn/GiOnzw1NKedANPko25lAzzmXwLSx
jEttKlrws0BSA5Vjhxl5IqZOI9JyozOGHKgIJnWHGHadHTcYdf/vEN37jRY980OP
18MMpPXXF1gn6qyuDkhsNoNQCUsPVC4VSY+QDRWSX6RgGHcwzBM55Ig81chbNQLA
TZwcWpy3MTYmEiNChdk5H+WWwoDv1/+NSW/fIIEueww9z2EMPFQ/UpNMBEcn4Jt+
DJEQzNBioz9iUyzN6Jzu2otIKOfbYyU/sER82urpUzdrETydZfqG7mAymkStz6Cg
L2Jj5i4dU03trEaLMnq750PLeEwzXbufGwNO3VgHgcooHZ06SD7lnxZaCXiJQMFP
MvhN7TCxMgRqmOry2gW27IUJ/2eJWICwuEGsWGl8x+zDix3UlhbqgOjm9sOk6+ze
MrQIQms3dAK2+PbjnoWtzYPNH5eXly3J+axXl+WCEuB2eyGHoW+w/N1wJhflrhFG
aE8Ya2NLkKOawBz+FZ5jiB/NSvEQ1TxtsPC9iW+v9WZeNxI51qRmCPmEkWbC2cs8
+v4mSdfjqm89YiXcXLn32Okru/9MwMl60QYndylkbIsupTgJn5Wab/94PAqe6eBm
oK1Xcgb288dFUy6xozio2hsN8FLrdQlJgjnlWW3M5BVPmrCUbSIHPxsLuJ8RPfP5
M//v6UTqhbgcB0l0wnBxjNdCGw0u2JE7Rtk7UT6OOuR8mHw/KBjX1VRxfME8S3vE
k27caI6NBUBg6J5x2MwAjJ5ClbHGssOZDLTOoeSydAXdBriT0mavFeyldsxprx1j
5ttb4bUGdcrDKmRkMZAr+69iQTuQW4xjMbU2pjV3UfVtMFpOLXShxWqEHh3UBqxT
cMGIxlFKhKGyuFuBp7IDlVFps8eMW2q2PTWnpQ2Zcd6XrRBQOTQSDA6k3ozPIIW4
4luC2MZiCd538bwhlXh/v7DPYinTiK+24JoQ23ZiXH+9VZwsRCh6WzZBE9/TOlLH
7NZ3daEdO1lbvaxltYUv3C3InMs76xBGH60KoamYgDjg+N/vsE6T6kqb9Q0gg7Sr
tdrQnCYxDaPWU1VO9yaUvnaG1M+7tiojI3AuMC/0BnPU/mwSjBNKWey1wtOnrwmq
HpXmN3SN0WY0ualLaf/Z14y17ogKIluN7A63e6fUBcz+iOaLq0bfhSEws8L6f53w
U8mJ9bpbAEKcx04iXv/kBam1qllExaaQTD9m13a+IQeM187pbcC7ygkKub4leJjk
eBRw8U7ULF0Cz75zNyPZIoWTj3BmQ+1xxmmaNU+PoTUyPRxPzVq0hsCiVkuIveBu
5ksyRh/whxeepuQ8nLk/JMJCPq9YIbUH+FMvRoqzGyjhKOLIi9AqG5UAzGGJjkET
tSl+flE4th0hbb9+DJLFuYYGL/IyJTUls1g8R3fCxyuKLlte4ErRQpfeOb0XLH19
46WNKCrhLWRvelw58LzOC3IYUhlr3YiRNyyzzQABTPPAhzxpyiA6CoAk4SjwL+lN
NM63NZAq8DA9YB4g0RhTOJx4VXgg/cj9atzaOf8cyC0hfhaq1Ku7O/uijQs6SvEv
ZNaed9Uns7gnFmWrZ3bAHsTKHPEVyQSK0fE/+Bm/Jfsb9AbT9363ywNSsWr4QI5S
M9ZL089mLwYiu8Hc2lzyWNkWoGQetOzDv0HmytW1utXxrsono0BxBNofoPV305nH
njn9FI4mPn51RryHHIZ9SfYV4KgL+F5yoK+ClogiIcJPbLE9FCVa4ykx5++ljAj7
Pimr+/bkaTRw70gNIu1fvOM1xyxXApdNdTpiNTOCFhL2ay6sjJPw9deFbLb4ro2d
jvqNblXw82rNNelsiiKvIXUTKFDzN/8q9+FQWB3DiEt1685+JmbWv7og9lkYe+Zp
E9UZLKcXzKQItMX9QoPeRLXnTCJyMpKTpsXgPv8kpq374ByBVP4PoRCjv4s9cznJ
ggqqrzvlYhIOiaOqyDjsRzmTKaG+6Xu/boSRqsn41OLcqdhWnnDIJ6UiuYISUS6f
ufgB/TJkcL+nfLDGiqlqIDnlglDOdKwxT54jzd/E9Erh7Gs5lArMLSWPmY4PXrgi
GQr/A8dC1JXctVmlbRCZ8gh51qef/WUlKHOD2UqCmSs3MPAPP3Cw5NFZQZrKCZb6
+xxDxXDQ6XkJ2Sc0yiXdlyFPKA9ErzR3XYyDQC3ioDA4xmKt55wnu2o3OYh1msl8
0dTgDPH9eD/NtlFJMkFvJJNXQuDnOUealPMLuC5V+M/qRTL4s4fm6WHZwNmIX11h
l/SrNPRQwF4swvBMJJ2kYWwFFhfIWM/Mp+Do4fPhbTG8/ag6Cz9deF3PhxQ6YpS2
jwRaQ3eSt0Fg0Zg9h22e7uKHZJOF5tKinD0nuLGKirr/mSLd1vgckHJPm5G9QQIE
NBHEZrhEuJOcWP/CSIDHUgXqrQzd+FKr4J3FmaXpYUruQ+lsJXO9xUYVOS16jmo4
tt+oU92p49zP7ajb13U5iMbrNIBVYN0bCe4g97+ISm3+mrUGHyEWygOOeHbLg1qu
oYZ2jNbv73uhDF9BqcCTRczWpFsKFQxbd7SqU0d+3MhcusuDRoGWvJDOcfPyHtOJ
4UwaY4Pj7inkcuyaBlrMLgtUJ213aWdLcslHqPz8O6EajtIPQmugTqNxigOBd5x+
su3VGBSRSOpQn1iMxYGi/M6K/Qnb/9DvwIwmPEyPc+e6DiL5oGZMBBM4wOjpdOBP
oM/YB7hZWtcHxVq6hkoc/nTPOzmbgDyhgEbAmlpCY6E0O7chbJImH4qubWdk9b/e
kAW25Hobz30BJoCsCEBG/bBAOgUEx5WVOJisr1uIFx4ssPvV4ENImHs6Ab3zHmKM
Dho+oGb4VHXEcamPcgRKX0FRbdV7uhQs0FN6PN8eXmgY1ity98l2+yscyEORrULU
tPngKMdHd6anhTgVBWkJKUCv5L1Mpbon58F1/RZwSy/YcLyVzzZGHvTg8HWYBELi
aaHd6pC8LrKhCLZXeCMEvBZJWvFY2v2zyV22QMT1PzOLIYmvCYN/6BZywc+OgHSc
Ta0celfDKPYEzyfSl20ghSWAxOX3JqbBiFY+jl9FZ74LmfJkC34q7SySHIejZxJo
5/0U3DmE0bs3tkTpq0bT9Njc7TlNqbbn3OcxI8n3QYhxUh66himzAV4rowbvu/rR
ayDX/Y0LkaDuUbcIi+eSH9y74gA1y8tMZUdGhMnJcMcg9fKGr55TJ9rPCf6wgkmp
N3FzKc5Z5NqXMTMD7kiNlyJbCxsnjguJ/RKA++AqTY0XXpsE6HD1II9/kdekoClH
In+4nkrZgYsMSlGSN8Vppu1yVNjJK64pI1FQD2XyilEQ8kf8J5mXuAW/xzVu74PO
jdzviS8L60KikfdiixMiWDS+B4v0vTPupnjPzfG46ETfa7/JedoATNjd6ekKaOrf
e59z8j/NZZlDI/5IYT9eCDnpt0sHOBoC/EfSui/wP9m7Vwh3JFLNgUeEHIBqHh4A
OtRtyd3c5Ki0vDcAOtfAXRTLztAId+hJL8nnErjvXiH8n6d6YX3mtn/vW2GRLOoj
302OcjgJzg89kNhcZw1/gcLsPZy1yXFynjFq9S05d5NwONX+bXjb1Kc6FRxuQY9f
sn40/wunP4o78BHoY0rH8zRGTDguRRhJzoMLjC66HCb+TGBmX7OLC3WnqGQ9ISiT
GE65RyqWBBoyPw30dYva+GtXf+sWy2om6IWzDc5yZqBTSDVz4ULY4IUwGDMebYwd
ulb1K6lgIEDzUSSJw9MThmt+mw/tTWYY70SlJCwa3ZCenYzm3ol8X/eAMbBb6QS9
dSDVuPfRZvbnrih9BqdjMDz2KA4bTnhtRI/+2S/Zai1qsszLiVxZW2qPEYHBLDeK
rtt1OmK8XmTkG3bg1+UiuJh/Qh3aKLS8/gfcO8/f8gwXF3s6VF8BVw9mFG9DX3yt
A1w57VRLSYdwsLKXeeBq+txcB9WMipd60ydhY8g5DFzULSkwpv344r+8SPbZ/gxk
1HjJaW26Zdkvd6LxFOub993KRY7zW6mbbbU6ye241eMc7N0IBck6NnpynRP/XyEh
D/IaGEtJQk57Z+jvIp7wdQMDh3UKTZvgYCTPofC3kPrdsmz82yGs5swSHmdZ7b3I
iRQk6etHYRAGBE1+rdWolfCvsbX7kuuJ4yybTs3FyqnbYTzl6Ie1D8pt80WVYR6o
4KMX63sgVoe+/mhgRMgp6KP8ofW6ZhgvbaYsg+Tr+E+nq3XrSVSxQbhC2dswWL+V
FzCFLDR/HXOwRWsBpcSgbj+sXX+oVBt5tqZJOVXEEP0FxHmZnt/M4qnPB7BJWZKj
F0DuFVWeg9aDpt1KlFmvf0dS0Hg7+MzpK/EX+XWC0R/onDwaKcOI8Z/1sVfOztct
c7l95IYB8nMD7Gnm1L3yrallKXE+YWceOta2kYvpwE0i4Y1Lacom8eQiGjhkKEH/
ntJ1FS8OqtRXvgHs6D2R3nqWGIE2nUufSeSgO7rM9SCTPsHTaKjzu3LMyAItGtZe
ItyYPST97dcS3ylRldMxgqq4c0n9RXjJXg0YmTQ2rObWlhk31Ssuk3HBm75pxr7m
maiXKOeNAt/dJhIqvaMz9uv787CGm221TjBhXhfqHpdkb3jIaPUTaiYyuhsCgNn3
NWQUq8C4ntf72ISTlt8j4Wo9KzJILT5tjFMorSR5mNNRaq9N6coZXgTCyofzLhWH
XpQdwGQx6Rcjx48lw2Usg7Zhm5leWXZAp7fkFojr8On6uu7WSTHTIp/5RvBBiunh
bAah7QOl9utkMdDY7Fzq6qe+sU8w42No49JdX6OLFoOnzfL2xIYc/8dz3Zs6wSZi
d0nFPaVWZ524sm5vzLMAa3W7dipVBmE6ulKynklah1UJYUSgV+cSvi/ihMZa+Gcz
+xi+X+7mDbs8jNLzoEffBRisnO4SDYk2qS5a+lSq+srPPb4GmZWh0X+FwoBwKAj2
p9MSTPprVV2pB/swH810jgFckL08V933X3OlRYh1nx7QgcXq5bRdxywuiJKblnv+
2mbBXTS3MlWPyHlNMt5yJX5OEGIT5lwAHU4Y6B5kapTZTN0qTSFwMtWxNNjCOMMt
h6or8NxBgfdHMJ2XzSIOiBCbkbae+f4+iQfvJmAir8dSttBCjzG6xmSl96zTPv0b
IqV1xVjlSv8sxslrnJJhbt5sgiy/v3FZAYqYcFfSrU0oh/HsIAiyGkOAGU4r1mh/
jxJn6tCcv4vOTR+9E4oQk2k7PJiRoky1SrqbAq1mY8BnCcoObbk7AAvZHPx+KriC
rDyoC/tYacs0qIANFUPQNObAiH4rkfBmcRsGlRKMolblOjL6E/cWsXI1JSuHjz1C
NLUk+l6fIyLWwDC/rgpShWVr2m6ttlo71m/9i6IIQdlJxVoLRgiXQkifUcX6WfPK
cCZmapnmbxT858Z7XaRbRevJZdHBcHvbHqAb7A/7WNnx8MlCI4ztco2tFOApGtFF
+5YJN6O0v5ZCgXgmNj06LrDsuUaKiNs8v35YU4dLqQdBweIP6S2wsp0SalxIqzt3
lrzvrJG8aO1+Rv9QjoHGyPpHb8aFWTSQQdyEUKP7lVQ28whQZ5K0TKEMcZDezbxw
vx6i1Lf7LgtubLIf2NYSp0y9L14ELjeY+ezi76HKTJB5vyCp1jBRmfR5bOq13ZZg
2CRAIhEa2X+GtvbO+FATjB8yB9g4qJGjzkLAaiLYZcQT34XAqtsDK4xvMm/sAHfs
s/inSJj5Fd/dpVYFR+BdvZe4w5UMSbqIzGahFIXhlWA7Npuj3LG+Cf+Qdmw0nmkW
6DAtYxLioJ2SX2Ua9nKLaGVAhJqEHPzdn2nB6xC1bekzd9ULSX4TwFrmVxFG5jop
tvySVPACPbQRkQqC0A8c7w/jI6yBS3upowzl72duFma7sr3bhgS3fDre/sqD2Ply
Tow2psZuVxJTUNu4iB1kH3fFxjpsY8+czay5mUNHk1z2is5FDRwdLrTJS2EMxBrE
wqYACRWvctuKqsGYTdxkU0jl8t/ec30XLsvHmvNL+CIeQAQWo37E0wcIvwTDTFNy
hPKkT5CbwKBjKOBPY6zPrWAvAcIh30tYiBGSLtmQRVsM6WB4uUlH5J3Qe5DHtEHX
uCkyBY3KcwdjSnpiZnNZxQwZzHP18QHUc6gDI2dJZH4nU3nWQAjRK1tsg0y10f/z
gKxbk0f+etowmH+6xN/9VuNMBLCElAudcBN2TTKpvfEb/IjIE5PhhVNu13yukcYA
Zrzh66hD8eep87bsuJgceoU6W6Z68RtvVgODrK+MMNlti9ULV/Ya52ghj6AMdxL5
11RYmU02H+fsHsD/TQjXYnBgQZ1keWCGdQ7qm+2AmgXGZcQYTm2qKFMKiOg723eT
HrtggjLFiEobGf6PdliRuipTsclxpw7KGUCYEX9AGSP5wz8wWndndSPXN6rarIN7
vy3rF0fqsNixDZ4+z9dVIltF58NSPWVEswgLM76vqnIZ1j65+cKKmBNayu/zPkXm
xFrS+Ne+KYLYN4A47ampcITLxDHGCmJyPSGisT8XM4XJnjx6+iprrRKwlls4ahE8
/RATbZQraxpcGEQIw/rbC553FiMaMw1I0SdZ0DnS2wGdtp+HGavcYNrAB0Y+kHgK
APUr5u94sYM4ulB9DLtQDR6Vc0UVvJ7Bl5UxSTr2k3pW3EAt8JrPuuGmq4gQupDJ
JhgCSRexoXfszU/FmqjU7AunXUPACzRgD5uwboPr9XAkJhDMTk69WSqjuhm3rHTV
MOLzPIpnr/Pnr3QjQPe35B49fZMlOl2rr9LrHxZYEPQ/RPVvMPPdTU2Lehi9GObJ
QMCK1WOJxPmqa1KgI3WPZ81PkUxgY2jEzHlfMPioMdg51qy766ciK2juhCpB6aEt
GxiQ2sKVI+ek1n35MBUrmB728fNK3P1cXIYEhqsI3TtKmqK10U/7HmepSpbvuU54
9vfaVQseEZ2igLCtZ9oOezLJ1oi+jWi6+3dJwC573gqXbBrMtQiCD5nyAiYAm4EU
z3mxOsvkoZUCmwh0NAMlXACgxRswDPkMQDw0E4xPWRZTgFq7kEic+vzWU/gj75Sf
tmaGgo35YrmjGZVKRv+zGI4os/izuxf+cxDuhY5i5MKUADehR1a2sg1vdEXp2cxG
uG5n5YD8Xg4W7ZekLplOg+i0LBw9Z9UBGlz/qpURAjaWwP+VuBrgY0tbsisA8HEs
mH+EXe2ttbgyv844LNmBVz7JaPFHsb7WO+g7/ug0Pw/jHbbHwat/EPCSahPGK54q
1+fHxaFnkN88EJNXjx68O8xeOedZqjdjwvb9igjhgG0tNpuqzy+l0ZRojLHPM26h
mrrMNsTMPe/V+gNgfLloxn4QB+78ZNORAqubPMRwYNzO4hM2Rm7/mw2RRvio4BUL
DIgj6ad3Hu9TgMgvQw7Zng/tEZv8GKgxpeMzmXSF8FKYa9AUYQj1TYU3639mSiCy
ppj6vMDzX43emVoEGQzrCRRaMQhPF/9UUS9pjwbjwy7xqLrdz8dI4rPR6WWOE3vp
hFu/2JIKTgeOrDb/lAGjtNZzpstHbuiQ7zHRsJSzACfDHtngjEw7MypU880/zzPR
v/TyvRdkB1KHI1RTD+YHqpxxxcRLAA0Y6zJODxdZcrH949fngmry1bfNTj3/bbFa
tHaW9TXSQNGGV1BSoJxJzfmP6DFu/ExXrcQYocKv+jVA8BwY05oPO4yQT4EyyQeW
cIV9ACnjR1vOQr8dfMpDhyGizlLvUKC1s/EVp+jVItk4fOYT4YeFl0j/o8ZwAw1u
9BGX8Y0zrehvkJxvAMs+lU9RR8pmJDlyK3tlmNKbipGh7ikivz9CRDInhE78X/Ih
9EQoMBEryIVPsm+yrtW76qc/bGWwDpVV+1JiUTwa8hDNXNbaL3MLzmvCA6N45slw
Z02bn4AYe94LJ4p89uHm96FOInxH33z/4wz0/d5GFrAjThzEPaxiVFuPdudkvktz
t6YH1L8FvGaMDP71GfOZvcTLT2bd74goh/OtIv7oumig/DDnr2Gl6RnvcDAl/BI+
7BhKXPRD47Hhhp9rzgn2YaUDf3ph1Qe2HtmOMd8agYhEyIt5R4eDO6HjcwBE9F8W
hv+0J4Rm/minmczjZ6Ut+mC0x35tQfzYpBgD5dMpOZ1/r9WE2MOgHWHAdUwQg6tT
WPZvEJ3nJMQhD8pvBNcjMF/AWf9cTOERbhndSxoOXY8J/SB+OORMaQxYNTSLIdpk
NC7FUOoyBXO0SLEh074jFK7i/zvWNb4nGXyn8sLcizt0H2isRZzc7ieueD30kU3R
6/jEq2TsvJC+96n9gimAkA8JhE8n/z4BuRygnDlGl5REjgG07W1+iSV8H4lSxrBI
zaPRIqY5qf/5CwIIvM2e516eq8dqQZHaAau+tgPv86kJTVlTnblawgPfftuAdGzc
xwRknhGCdrm03oyjGrO7ylai/Z6Mtn1iwg2/uUL/oqKZQMmxpN/+qUiznwE+ISBq
veYqlYBQWhxarOSniezCa7ZPltieNJVHRM2XbusXHjkSm1H2RVFgdGXde8HB73nG
8kl+8FzNTWMyHh7eEFyGZ8rir/YJJ3TcPrOR+32aj5co1Z0BdOedsGWpp556nDPq
gTgewn4SFEBo7funqiNZGS5B7OGgW2CD+ypRwQkyzQsrFVLWPuQxyOyGpxnH0Xog
jLKeAOl+YzjouobUdQzzRQWMFd8Fe0LIEtXz+k4yOIBgWefMvlaQgTjepZn1vr+H
LXQaE9bnHxdrJmsvCZfq7XrcPbeipKab6nyS0ykOFTZ58fu3RAK66OAVUc/mPrZC
mfUpzBQt9AEI7GMmvseAlY+IEgAkaFijGMx9cDHjoWEH4CvgUIF4oj4oKODd/UxG
w0LhCzxNNRD6DPAisYkeOExm+CCyGXbXoN9ilMhBB14WC1bYEcyleWEWKZ8A+W6L
7T/XQoJj4g7YDvuQtupT+t0nN68SQgo9y9CvazPJf26drD9p25crkW0CjPTtHdzQ
AqnAD7TDjnwk9Mp6tzplWfDn4GlGMQrJThpGhQwQUN8ZFsexcmrXmrbPU38T7PtP
XYRbpgbRrM4MDZ7che/sDXj0mfFMxriQAMhaESd2RqCEPjaPzwYqx0/ltU+LxMcQ
2S0gajJd0ShfxFHFa2s0QXiNV6KAH1/tcY6GEG8hXhuJ3wZjZc4xVQLYbFgnbiwc
BtojOAoJayRnH8y+c/ABbrpyFKMoYelXWAUi6KmZIXR46cW0r/C0W6ve4j/I54Ma
McB3Z1nZSJiQ+P8XG/00NJQqUyP4t78A+LRrQX30GCINYPnrMXO5q24ZQNU935kv
U6twZeV4ytSrh77tFg78mVuAV2+FsHBlusTu5nmOCYNMaFNJBw/+n0MKIGAzyfyb
KdjCXEBOlRGLDhBvWpb/SdJRB1xIZdBrVsLrqzBCl/gkyOlMdfQ3QMh+bE5XuESK
L3PIB7pKi9PbQfEFzsoxFY8fr/XUL7dR4DhdXdEYkIhTZB4As6uYpPG7HI4yw2co
vHo7TnARUlpFHZcISICytkGHqhQXsWNlA0kOrnYwPIjUBIhvuZ0OYYdzAdaP4NEU
UsZQJRO7f1hA1w9p3Y/gUXPQVwgzodSDgJ2Tcz2a7JVygpDh22jSYjB9BcN3X47j
YaFLsOiuW02FKBwaSr8XPksC6l0FuDMBUeKW90PT2JkbSlmIf5WXlj5tcR67HSSR
Ttdm88EVcfvHiNQ1ibYwZteP7915TXeUuKhQdsJOfoMfmkjSTqM/vK4vvigSCin/
/rc/uQidl0xtOW1T2T59hNWTYGl8AYfYi2EHws3LA2P+b9g9OpW1ObSM0LXLn1fm
6s//R9k08rPdEhC0m7EczaGcXgX1Mddvd9sD0b7pJJansRwGU716pVcPQR6fvm5J
a46wdLCVCvIDS1CMUWY32koec8OFk9dcT5m7Sh+SsxYcrI3TShmABqo44Sxu0gh8
YjCAoFi1hGi5SACaKS49eeWN25eEwip6sgILwHhT257p4NU0PwNCBcj6frA2lLtQ
452Y7ziBw1vuZruc4Jqah8C0Sqz2HkfDqhqvYTtiYhkVo7MZKFLsg2qIzzlC48kf
c5RUet5pvNWdi62gr0ZyWtcQKJxEOj7EawxhBDufp/F9tGfzaZBWH1D7LeA0R+SL
Di+Xp8XlCb20QZYIkIpt0OOJnWMHy9qqx1LL3F/55RioxnnigN625kAGKFLEY0B1
7osgzzi0rDyilesd8Y5MIqfQlIF1NESp882jaUlvtk8EUpmUheFtV92QEJo9+lU8
QlmxBQe1HnhPu0jLfGdPbYtw0rxgQBU2oWuAsc750Pm+ZZ+dzNqFtrrb+7gmzV5Y
eu8xldGGNoQB5LzKpr6/oqxxlBq/+aRkAcJPc7oTSX4Y6CDEP/33uxdNnHvP11K4
HVupLkrxtwthljg+tspMrs2V+qRu0ugvlUBCXptV8JrBeFi0M8OhZxQuoZ9ykKRA
rW7oZthmZ7yrp8xJQUtcVBBEhJe2LbU32+RFw3viebZMCUDgZhjZdB4R+ACtM3GP
uSHoO4YZ1sCtP6jH06QE+JgIDW7tGHIgAcy4l/hWh6quJwK2vEXA9LdNFgSxZ9Qg
0urXhVCNF5ZVgejIAJlDWPSQpwsH0kdp1jFyV/fQKZXjHNfOC3o+EmJ5/vxFnXdG
T+eMPQf1n57oAGNJMPxPXuoRM08IEDLQ6cTxcFZP8383MqRS3CqFWDg8H4iMfZd2
uEpNdmEGTmKD7ziirZIIDZaWC+0dr4tl9yzC/Lw1jIx9AjL+N4fL6Z4HdzX7s0pb
yfJCCRDMalvJTxZE7NGEuwVNe9gGEw08S5PiSZXEscva28PvEHI+BInRM6oTkULg
ynYycgwHwrWfP7jbVF+Q+Uf24kfPm//s0uA0gvqY296770vlUtLqaED0dBR8KRQ6
VEoWI27XWD5SwoyerVTqP29KXztc5kw+vk6/K+P93gCQdTs0Vlo5+SWlevTMmrVT
nmlExeT5bd4iZKG0nvP+//1+Z33EHB69iruUx4fBVX4ai9i2Q0lAK7gxjGWjcej1
3OuV3rVbYo2g7NJIivIMBi4h78RNwHtDH5s9DrfPYfjAJsLtaa3YtEpDZfgsyGa1
aZOLLIuJBYKc1HSiJVh1lGJgRuplN3D7tb1eASoMuGChZ3aZnwrSPcpd+Rc5mmpv
j/dsmC/XSMYaDMvSWqr3eM3ZiQIAK1PKkjb+sp5AhG56Id+lFdUcjUScgPxpWeLT
h+hMStQvA6fj0hlITnjFAfk/DzSRs4eNjgzN38nZfkuj7nsg6L6jGB0t2K9E4jkA
u47bHGK55gzW1WdFW9YUMdVTcNP/x3PbhPT+8xRhtWD6Mr8DH+M8odJ2EHdHdjrg
RYFwFlPEnUzg9nfEiVJ/jQH8c4xaIpI+F7f7zSZa/nJcgyhFw4bJE09UTnho+CdE
NUqb9DRudp4sifp5UsTKXbe+cZnpgUeVMQrJY2vExl78qQz32vWWBLEFjSeXhMo0
ts8yF2Cpn0ZZ9Y8ww9UluDjtvbV/WO4DU8n7p5b+G51NDQo1p/5y5vgjoZgoppao
3yM4d9ZUQxz2KP3BCgnrRKQsRp2UIb168pH6H2smOZ2kvmpRj9a1rq2Inwc7vTrt
5gXIMzx6eJ+A3Ovh7+PYe4Ftvdc0WLfVCpL2StpJFS2OtBU0qHoYdfAlk9sZgfg5
lJObnsV+ftL6bU9kz64ltMsFYHjichUCMqeTvnH+ceHz46punNV/yigLSsjDz4EH
4ifcEd6oVwM6dVdYaBAdSb2zQqtzVaKHs3Auv0yykfduSQ5rAqHh0NWpVL/9HP2m
dLZr39zLZn4NhrHsN6/62k19l6P2qnP6qKGwivpxuKdTLX6kS1+UQEd6S9KjGpA7
jTriWGtrPOk8VkhRFO17lM6ijzWlmYZaEogCmzzcR2zaA4dTH3BR9noytHl5z1y5
zSHFWla1DnhmrTOHnPRX+wEANzXGoUyml+WKNRp+z4fpMPIOYuuf7cvILKChssfT
11T/RwsF2ItStjJlf8fXGZequphYV1uOzGmq098aP8fsw7Ez2i1BqVpv1ELMudrl
f5aqfJFxVNpbuf3Xci64zO9jl9wGxMEj22jnGbrSXhJXC1zCHUynN+CVPtC8qVot
bHfYTimGcZwW936EMPOu01i0NBJEP1kq/GXgIcajEMEuCnpebg2S5sa+W607ASH5
VpxHXX4KDGN+qLdas4FqQBJ3kCCe9O8Kz7R7jp3scNVStGPMM/WpQdt5XffU7RUw
4ZBWghMwlLEH1hSbvloCgu4X1NEKA2WhLeQnTh9lg6zNbwwo1YYdYpJxxYDup3oI
5wHtBMj/WTJTEfBoeFr1sWadlbZ/pjvcK5G4U4wkp3DGhYwjN0EdUTHoeWk7Mjh4
g7L/lKrKHFZJ+zCA0to0yQ83dUHy3toEvQ8OjpZ1V4IQnzYU+hT7X8uT3cpFTpgU
eCsM9W0DrirvT3HxOr7l6cmmviFcMP/XjufZW2CFnqtfJuRgMzIrGxb11LuEoLpH
V2f9RMJwhvuUgRi4rdVUCEYoDOnJFP+3SQ1iXiguoK6edLa41rfLhE00ztKyqlnM
CW6BXVf4IK8qNnGhsxMjjCYFhKCKHDj4OHnVV8TQskwCrAfG274gGQnlKBFZhTzn
YkulXDDrUgTjjU4xfsdKDklXPZfrGIlfRmCXQ/qWn0VlKsiks+UnX6SoFh0Mj3t5
fo5e2GkY9W6eHKBUIRma1Es+xX0Fq/HgFLjlehewToiw1/Z4bwfPBCibULHuoT7N
xjAivTl5pWbovKlHj8xC37Zmfm/Et+tgM5O73zFtBZxDG6Qyn0LKbgzDDl6XnD99
BCpJ5+1cKI0cxxkrYjcVK0Con+bBUG6m8CvUKfdiG7DfMRMnyRmrG+Z5DhkfAOag
3Cjtks57DjV/pgd0L2+xBv+Ryz14exbTrNDrMgJLgo+LQ8w1jXzoRUNZv/FylhCq
bN2pC1pgMl4bN3YVZEviV1ynRklxjYOL5exZbYF+S3j3v6OJ/3sMdSSiy7QBbFUx
/TyN51DT+mjvxMYRBrXxr16VJfih/OdjC9QQej/von3hTD4rdL99WYgviRdBH0Qs
5LTem5UUcMnY1UICqAdsCdmmYYHZvKM9+IZNTHlx4BJUOwTpBF+jyZy5l38PK4C4
kdmOIYh2TlcO36Bzg56KfqepfHV+12djCd5cZu2fUmZBzfT/puq75hudvx7HHzxZ
6UgmmT/D2hWU4KAZDorkx8ToUSYWiLPYVAFEoAwYPCCb3aGDyZYAwj6eTrKGtkQ+
84x/ccHjXrBHDMzAo26koCJ60cRfSBc3djzO4HWCcOsEtpq96mkJGMPcPJDQtjqp
0iHwTpjF5T136clhBKYcypjZXaJ8VGbGPxnQ0sYed0q6ZXfv4xR9plQsC0DVmLvu
hrMvHzaKeu+33JaJ5ljDrqplD4RbMzaXg4Y88gR1e0rzhNo8VcYsL2zNYQAmCuLy
3Swdy7WCt+zo0wiu+b2TsigQAML0t+gTRVl4aBxl/fwryjIQMoo8B4fY3FZI8A/X
BT6nTRNhGsccEYHI7ppLk0QM409SKOAeX4rZR+1sXBvylMg9Xvy/NvOEo2pt8kXR
k/GDXLtzO5BS9NlAK6yB7dfPzu50aXORnqKl43i4J77Mjhe8mmOH5B7/awx+yT/w
GPEeBoEFwwxbtPxSeaUmCkwbCoWucgCbVhY5vphjITwgZbAL2uXwWqmUCzQsRtUq
gG1CSUbOI4jZMezU6Rrwrs/09bN841OlUUPLRYNEAB/g+6yeLrQjx8FbSFRQap2v
DH6vWU3PAg8lruVOABxO/Z/DJG7DqCmQ5hz7mgoyIo6flA52ViPmObwcKh7qrpmz
28HbVnK2qvmKWilJeASHXQUPmQ4SzPOQPAWEC1ZwIbapdX9nsVD69wchavH8cV9U
yV6aVeOKnPpqq34kQMuItGwKmPNSExPhLP/hR4hDNjlx629+vyX6uFsYBdAxmO5U
oJOlR/urjgZLxbIr90iiugZJSP1Wrg+M0a4QeKxz2ILxl8UYaMj92a2DEWVlQDRn
jIKNHvwVMF6rfs2FRIPwBpSQ77KVH6yHlONSnW/rRRqgnUaSYnh6+E8aFbiBy8T8
i2X8IALpB0oAShHpDMq7vtEROAB9GIcTHN2N9HAuhSg0mrJlM2RHb+6iEMp0kXgx
foGak6Ms5PtPdjfQdQrPIDI8Yfh+Y/IbXKYQ95KN5kaGAcDNkUX55zK52qAIwurq
Fu1fVQVF4yVk3LiNr3t1lBBDyVsNKLFuBAXq28BG4/9x7v4jjkou4wAIhq9/BhMJ
DiVI3SmwLNhTbDKK5hSJ66qVMgMteNiQ0/rbdBBZuMVPVWtyslCP0vh7xkTuiXIU
He5u8dpX3ZN6MG1DHviSNsh9csTvpU+d7wPyUlfYcFpl8yG4fLfbPnBW527rqsDH
ua0HUI5/pK98gCYbAm64GkE7NG9KGxrN10QUqUKLJKKA1xmNXZ3PTOQZzXoyxolE
wFmVmdB1ta8lsqEautz1Dayrfgx+KNnMqfqXzqqtmK/cegXnZxz7QB3JriXDFpP3
+xp4HwM38idLmsoH3XHB2vnCpE4R588ZWYK8A5b25j+ZZezJrMJaqL/USqpaZxhD
5v9JJpcH5+LOI7FgIJuxJhtiqJi7LxNQhjcOuNZU7+2UbdoxWdb/tBeJkdJyHDUy
0r+ysth34F1L4KjhJWHJq5mMD1LGuftQ/odja+LCCGfB5pjp+K2Max5LQxiiydut
9m/2IsK0mfGk/8pNbv7l8oRjgFJ3LyEgfs+C1+L/z6d4CNlwRo7vpYxUV2KddSRq
zGKfZJzlB5obgWNDmbAlv5rtZjIweiM+IeqNXXppB83rdJWR8M68csTRb4wk8cMA
PO6FEoJKbz37+8PAA7FhwzNDfLz8b4sXciLfnENRQZ8MbC5Ur56YcoCtnEVRNXGP
IzgbWD6c0aEGmKeFeOCIIbAUjWqP2cFoBnTHWUUCtu0gkKb0vKizZ1E71uACkCQP
gjvaK5bQTUvaGhm4gQKf8sxUkvmr7r8nGIUynf10+awpInVMAhhphYYFQqOFoOdd
VGE3g7La6Vr9PUcXhAncVgWA64718R1CAYDFRiEfCV1QOoFrCNDhHiv710l1gEmj
FrSY4NusM4g43NwY45w/609VHPP4gvrZzK5h7H6PBR96G0sFnRymGxWjM9WDPSYE
9VyJqeN127y+gVE6gZvKyo/cwt25DOa2qqHc1HKiD9xv2vY7eEt1Ub0pcV6r9EOg
G9IbiN5dnu1BfBSfM2e0RxI8ptSC250V76gmsufMZGEksNhTrTVVPqSsovCxeMy0
zW68QEwls5dos0cBE/1uIbg2RYtzrdLMAz9kBwIKLQInnbQKIJwiE4uCGO+HCQ0+
aFKs9I13gOB/PcCQWoHcL92/REh7H/LRHxY+DZlsrn5C84Gsr03FFwL79JD8NzXY
7R8fbssDPmSU3k0w7HHxyUx2RFN4KTDx9UbUVcRvNq4zNRYqbx2wIv5G6VWFNRYu
eZY6wxjp0U/RdFEJ/js2rR/U/0rgU4YYn3kwpBg7t/c5/erMm4Amy1y0xobyOSdt
G6lE6Y10+p4jUXjp/M6qeOfy3WS6ak83zlj423Yp4ctQ/ydh5Uermp6FuT5dJkHT
M/6Johr3rlDzmlWCPTeSuMOtOFRe4tA1FOInh73dXtCNgOrLRZkOzb2nXjDN3SD8
aMLj7vYxKv6X6KkmZDsOSg4rJMeIIufVUSs3GAHsMGGp/iQrr5763+QWj4layZ4K
SAaiPMEEJyB4mif2ORinwMUvYtDkHzr86ZzB+FQEZk/CdzdKhp9+eLNQAkW20ElV
we6hEKhCdjGdjIyJzgv3efvyaWWw/06NcM4tVHRJButc5H7JW2I4QaPexW7SKoAt
JZNh2rJ8xacHOWKF+kKhGrafZdhavryuXEBwhZ+53gGNH7BzpqIqgpg4i9EPGjOS
NXJiULYnyGL9noCOMwQnAFUNwO8qC+TmFlbV4f/Ywp8UyK22lRH8+Ke8EaeIXr3t
g9VQ4GPGB/WSde1eKCg0i2NG32RRKbPlupmas2rdJBaqHpuDmxtsVYtukWlvCmpY
t0sA9vue6p7EkN6q8gbX6gP+FwiNXFLs+Z30GOTU+3xuE16L5aUK94IdqwJqKEFZ
26CudA0JPqgBwPXKZ9HMbVkEsRo7GGflRUSXAPjLDsEgBumuO8PTQ/SiO/4zBAoG
kPEwm46PaFE1xx1Dsyp06CmoMcrJ2HkHihmSN6+Cl7JySSLMh/zfcJBaOeZVoj2z
Q8/KQZf8JTQrzJsEjaYsFl69gpEyXNLUB2+W/1BAPAes/W27JJnWvhfXGX8JHXKA
DGY3t+MkAzJT+xH0RBJ+P6he+dsaSscOHbcCMYvyyXPLkFDPw+O3ClxM3JiR3kJE
Ij60cPW8z5vseGd+T3dTMA427VGFTSV3nnA424V9mwOD4quttmWDq/f/F1OCAeE/
3b28UQ60kDNmqK3k0oi5Tm/f2U2DlQm/+99RHTjUXgU8KVqqVJyBfpGw1g4PcbNg
SNKDgWsuaTkdjVnRRgeMyAOgJpkFRZ43c/H63rHa1BWVkecsU0f77pnj+RDQkwCE
nOiDgW+55KAFImQjbczZLbrSOkY1GPBzOZ5DZOOeD2PO3vbTXbfNglFw79qHutp8
jOZ7tHkaxehHUcKQNZWIK5GXIQ5pE7APgS3vXbWbb7hSEzrRsVbxgS6pOSiuRxQN
8ceRR4o828/yQO57eprym6ggz7ieMxiUiDkVl2VrLN5CI3jG7pEchnf7uKlg9h9s
2Csqz0tZhXOTmjfbDkGDyn2PY83kf61yDWz9KhQhC+hk0iu2gEmqpZVaqmToe3vA
8Yo0kNj9sRngR0dEZM1LRuhE8Zesurua6rTmoLi3DjxtjB9qOanLHR7boV3vLAme
a9wKneXw4LVQpre4Dg+ADgpHP18+h+f/Xu+0KnxRHZv1YsCH3dwBapceR0fLBmeG
PoBjzK0jSFa3v5BngjM9Md4OD0vR8BmSHaeG2cCELxxN04ZuvmBsrXbwv5Lhtuzs
IyvhwO1+GBMmrDf0+U9zQ2mUFZzpMxLMuZtjmoWX+Ze5EWafL1/RDcvHJ9kEmsE3
GFCzoq5urdvtelyNXGPLW9rsAfLYj0pKy7mwqYtS612ikHsXAVVlHOrESAY2qayb
66XEhYZ1l235SBgkPEC6DUhDTPuiz+RLN3IklVkvFy2r5VjTSEKJwkuNsIXV2q2z
Wrdov8HIdRfHqSHVvAjgU5wr7C4ainRoDlEfdbMjbzeqrzr8bnvOql0PF58YyuyO
BPEm/qZA5nMR/X317tJsBL979La4REU7+ZaJGtrYZ/ya6QekGS2gbmn1EyFUYicW
bjLFLrjiglrjZpmvnI7wFkxl+kXABUMq9dJZwB+yb7wFhd8wV2+4LfF/sETUbXrm
/KjH07G+SXLtsaQaq03kcEP4Ak32UwiFhTSPIazKzKmi0VRrDHRZQ+H0hulebCUO
jV9lhvdwnB18kjUQgZM+cftm7hO54lbyPzh5Xu8AoTtqAQTfrVoqLhp8zcPK3XHl
xb5w6PBQ66Ygbp+a3j13on3Oa6ONeqBmgJs7S5FAQjCPB8J9Z0x23cBYLsr/JV69
r9PbbwIPwH5qp1n0RtMrQWBsZytSQspmMOxj/9X9+EIgNZv/UWJpeazMKsmAPQDB
NpDXE350UWEgWwi1em1w4VKNfnOfSXQVIsyGsIVuDBMfQoF2P3fxCg/QGM1fCPOb
afIH5MtnRj1NslRqsJ/l8IfJX0sL52H2QoH29rp0NKCD5dHAbXoBMSg1yqo8TySg
FypIClsHLcJVILK77liFESJAJaG+9mUjrdkP1Jgc9jgXMK0L7TKp51+GdkOpn6TH
lU0OuVVcBW/e72m7DPYENSSJYBPcGe5e1e0Od9UolEapbLwQ/6UCg1TDwiqtrEPf
S0LjRlax/+dbaGDUy5mpekGovlt7vYVY06/gdPCF6widE/2zX40k4Qz9XyqxzfMT
b5zH/OcJRNgLGRQ3AAs34Uinfs8Rv6Vo13mtKBTWPSbf4lD67Jcmh3JCLaL0Lnmb
vBvHqZ+XsfslvoI3wvu7lt3VNBs4j2Kj1aj0CIZcI1DlLTIPkhjEkqfr8M4+2cvC
xR+GkWJavgZiH1NDih417G+AcPLhO+a5OhTtO6hRR4bHsqz1U4W9sQ7+keLPSvq4
CjQOZmny5FM/9QvbX5/BAzsuND5s9CdXmdiUOHUo2IoaF55g5ySc0Ov6ZCPFFRq8
IhU6TUtuJ8XaVKz98F34kxjbRYyi4n2cDwZAs8CCDyL6dUWgL3YLN0QdUA8PO/DS
KXZ74u6jPty57AXyk1987Gp6YZOd9ayNcBtZo76ZAxwFaLwxwymU4x5ZyyPfMEvf
NlGj/6IhmDn336aJPHb3OLNerAznKNHVKSuF/VgHHyCP0oyvt6AHbgTvbVVjAX6B
UlJTRHaAxrh1Dy0ioyehQTgcCNgwu49CSmuteE+4Bfj2/zY5NxQSqAc3cXxh9gJ4
qpnxu58jKaijK/s7p3vuVurvq7qlSxKJJTAepYg5RjKeJvWzoW5IzJndW6Gz9xEG
jeqWeiAUYzSegPxyGab8usxXQQVwrWx9xSYygjlI9BMttJ9OqzPV+de9Z1kt1mq9
3cjlD9mPe5tH6Ljsj0gE7oh+5hWbdcgqFUJSWQH0I9kabeFwpebtxJwqhjMJEtrh
00armuHYfMXRwKBIfvQGe9dMzgsZNrws+5Lxtw0opbR+x/IfYIDU5r6OYwdI0/U+
NPBqndMeHXpn+v3ogDVqzJwLTNpmgqRejKcZhTCpHz1GxD7mb7K2W/JMke59X84D
l3WSmREdUQoPCLUW8UPyUlOvL/dZekxPjSNQdX9ogLIBoFfPfpMf38tjWru1QU27
zp4OA3hGnrUVDEM8YOA3cAbwi6CLk7m1J24nLzhwq11vtPGBHvRVm64z5H5VFIiG
qshsF6jjgiGE45uUKNi5r+t/ECjPkxiefpAIJm/ST4JQQHwp/ORTOVbFbqS7bspM
yBSDHQQPWRx9bKJM/FY6fIgGNYZc6WsoHUcwNidw7kxd0EemikZfo6+6s6NU61Cb
ED9uu5/zAeRAi4aoz7uBBZOZ0x9vULaedFl4zw5CT2KGyj8xonuZC+wJXJ/IbKft
KPPYP6ahMMuRc8tiQkgNUJI3cBB2QxYEdMy19W+2nENReLCNf/yy/bDcX1kujkpt
Yv4+9rcSeMeDIaKSDmtW97Slg2oweuuM63mMdiAfB6qvRBLtz0Kcar6bTFv22Aue
VnK3nae1YBiReXF5NpQoWcG4mS3oe/ZGljeFt9IttRAch2zuz9RM+4RGMXJjvCoM
NDjTax9JJZJN6Ii3YTMx6YAO7TCfso2kZjprafjlgGvdlPMHocPbFIVabi9TE8FF
qqal1J80JdbXF+4NqQulzpqTXsGy6CckK1aCbCKZuUN5ZmFhqKiXPXHvMKE7VkK4
mVLlsq2qA8/G47yS2QE6HOuIUtWiSXUBwyyX4BYNKxHD8DfBr5iuXVBJqtMtMG9I
5JmHmOm1Nbk9yZMdyBJp14fuzFKLpdDIrhQVdxZjkFXec6CNZhePfYuWAqBVBLti
FNlnYCmuAzEJh1cGegS7HF5Fi8y1wrjKYBpMoDY4B4CavctEXdBnb86XIQvIcY54
E7Y5yoxt9NXXGKnVy/9esaQ/HIAIGMIvgdZSPwYrGabo/zeGY/8rQhZI7RfbO3uX
jXiaGa4NUo+Pucafs2hLWGW/2PVj9GaGhA/P9CGSYe9b5RshYVuCqcnTJHeirXsk
X+C+En2PmZ4Vqp7yCAh/qPwCwx1ciUZWGCak4phOK73leYrzM+1MyyLOzI5ZerWT
/8VgRlfc/tzkzI4djKgOXitnd9scdOrsDXLQy1RvtJeMhWyU6EAH5QYrOFEyWW0j
o/TELJNTAdiiONZT3HQLEH40NMXihjggAMSkjz3EPv/jOva+//djnf8zeVpKvsvv
qf9a9NNT7qStyTt6FQKi87hzptA7LptsSa+Xt31fYF5TE0zHsB7wtDxVkzmEDeKT
koiG9zNJFRt2ho/wkBOUqlWFMaFycd1Zn5E+xghsqA6XkS471MM+ygWiyofIKaZ6
iodHNItDvA2K3bOs98zGkjrjdt10tT5ChWzWCrICHUc2cWf/xMF2ClT4FYZBl9Bu
NNWhKeyOPk2cywbzo5hLZ2McPmWlKliE9zZce6L0pkMs8tF4lUCQ4BWKyB3R2o5n
U4NUa7H38wVfMMBhBQYAnh0nKEWW0nZNc1gZ2J9jxVkMwOuuO8rqAYCsAhUnER0m
LwWDhjnZPU6IBMqvteaTnUOL8/qcIRe2RSM2VPwHTVUpjPjXTErhW4PNW9G4jdB5
+u7IMZhz8y4s5guzXSshQ3s8sng87YKEYLOj4LY24sYcpBJx1J0OocePnJVX6k/B
A1lpqUCdrBV3GsTB5aQhFW1s6CLOgoQsgjzMq0JkN07UIMNWDvSRZsyH1LtadRlh
CXiIVxg2hVbOEmTccWJI9wOqNim5IhKGqoI6WBzU2uo9KJ7C8TyJaCWWefTW02t7
XUop5eQUJBBJF71fP9rvNlFcvBK69ZUhWhumhLM7XRAdHcZJUa3N/D5+zJ65qE8Y
pHDVtT03Nx7xfUDQuMzuOe+0jciE1/tFRTiIYPG5ImMXCcPeL0ZpcArvicc5kGB7
clvMZRutmysSvY3vkfNXgnYp8t3JKbPN5yoF30JLnTR8e8Qjo4YwSEQS7XjNun64
t/wbG3BmZHoOl3rYQeQTeEf5AMDR3u+oiu4YpCHFTM84UDBYWv4/DOFOBEfVHlr0
ClK3TCAw0Muzjwo4ECW7aQ1t97LZh6S3w8lEEtsY6vWvSyHGPxqmSUtnEI6ub5mm
aj5cl6plzZ7uX5wleWimxm7o6tnR9EuoEJKEu3gDgTcaOOyblbhBwI6Qbf36Eau0
Vi6ZviACDiaJJyulxwMjATmmA1yf0ymVQmC3aDFG8QeTWs7k3mpB85g8Bz9H1AHQ
nEk4Kx2uvn0LofvZEW8567tw+Y0fs59e5VAXBd1UWa05m2ao4Tziaxmg0BKijjrF
63ZGX5xx0sX9roehILdOlW/EcB2CFgAihCnYP3mqqhYO8tVCsRfN3a4TDXFvVVq8
IFNfuvmhPWsJkDpTLWFPevQTxGXn+5BSmPfT24wVvPucXudY/u9zhNdJtzlaQftd
75UJVYmgL0cN00RcIcEwPPNVtjvoAcQtd3suEZFoUYAFM6ooUowL41tGNc5dLIbM
X/K7UJ0cqyf+KkrjKYjKTBhUNsGL/YpjdCVOVRCz98AZ6gP2CC1JGYzMNqPny67r
SqZblyFu276h5XBMuwZzbVZd1gO0Sp1lQGKiTAoxmfmCXhtp30dsIHDIYQ1g7RKz
V+KEIdev9c3N881iBojdsTdpZ52zS2dHpBPIOoFYJBBloNKH4sGrv6TR7MT1hKmm
Hkh7bFi2u0CStQS1pjlNAXt7HnbAYVriXd3BUGKXwHQ6FNh8MWQCHFga7JCtRHgx
LA0pPpK6o3kOJpdSVJIRG7ZuWnNzgnjQPEOHmk4LilzPoaYQCu7kJAYDFMFvjlhl
tuBfbwDg3rltEf/CbwHsXsiMCY8LjMWrs5DKwPMgHjEu41oI/lnzglSnkS5c/CGi
w5P9X5tfKqgRr9YKDSYxg1BUk/NZEYIF4y/zCYf2egubQDel0jKtQwCXgEXEV94y
dH0ew3oe5j58AiS6vEjcxWbM6HO3/R4tKg3MrP528SC4q4PmAyBIJwPHTwArCQBw
reJ5Io9WkSnXwxX9kQoTNd3xqZQ8GfYToghvni2C93HNE7QcyVr8L5IwG+KIKKZa
bZ8PA7vmX6yzA2Yt/8YzjmNbhc49BM7RRz/bmKgFc35EUV1+ZY90KH/JORB71ZJd
obaXo/prfKgTuMIbEhWiKQQewfHWHrbZ+Ps1X3Zu51sAkmHX4oN/PvptkM7Hp9vx
HVF++pkyFlb9r0Lz0uyqGUI6e5GOXw36NRjj49EUuBpXz63VF/Dgv+VUYjyuuzBu
8V865hgFzwNNuEdtFp+wNSpTEUwyrOLb8/TIlavzuG/rFBqmQAKKTl0CBtjLO/mL
DgLd5lTya4emLG6wMHuiBw1tmfcAmG/lGkd+FArwJ3cDsPVefdKwBuuFy8zobVV1
By3qUr1STEgTphqPwR5XVfIkRIwjI3mrIxguF+Ck0um2MlXrHhOQ/trIDA1uKplO
GH8GJmG3w57GovGqMTvAEcM8akn+joYjYpQjbDqEX7zIENhEoKMpHk/oc2rcGcAp
2u+I84JeoqyaOYdudeQoPLtgs4YUvs94plpf4pxWq05TYLvhTsrCmwhpHAxc1xV+
di/50NJLf6oKR575QXWIJJPmydtSpgwqDzCS2XnzSKgjyovFtlkIdNNyrVtspukb
wVYurOPQPDzaIqkaYYG3aTBIxx7IsBQTS0S181Nl83rRVbMhXDT0N8ftMMe8r2ak
qnM+BQZjsLgKqJ6mb0IAqF8hJ5RYIrQQhu/sb6H+9Eu6tOVJ+RZK7NpsAqEcfBM/
yLNC98+xOvQMRdAFeRd9jMZ6pqvsoMKsYWbsm+MXHpWjxIoSVHM3PHFDRCIMe1VC
IQitKkBsR8krG076XVmKA7ENgh4nmgnyJy+OZfYG2sGKiVpOSxlHNq0/OC6lVzLH
2UEoPvPtYdRvDRyRQCCaK1XmFzMkpsIJYnZ8Fv6cF8khXT7x3d2hDKEmBBPuh9N3
rPtwoUz25YL0Ch7YARk7aaz9AdQxzn7iqDdIiHEDnlLdZgmm8R+V+l3lJHWWoF7h
lQXecatdTprjk+cUm+Gx+cASY0teBJC5WVHGKATTn35YTLad6JhHk+fX3N5PgwKJ
ikuoKAGkRz1cxFoCmj/lbbyIeYiphUMJfiTwTNTgoVMjEn4/11drg5rjf9Eyv8Qk
8meJ0u8kE8sdgpEPmgmDAyvYz3FAnehusFGGj/TS1KIjS3saSfno8wG2fNWjZ9zh
VAZ2jvYF9O6lQ+uZ5frY2mS25Xy96eWzXQlVY6UpIQgf21sX7Wkj5O+W5Oq1Xlpf
t/+4L/oFjoZazKxkHnHrINrv1UiLxZ3NvvpP0zbjddCBCccsK/qwxbNKv+1QCqxl
xStDLypiUfW4eQqdtw5p8BxavWRVNmWGNkcl3gQF0Q1BbHdLYQlHu+u/wFG0knBo
UHGj7EX1A4b9Nod9cF0PrWV7nufiWzwadwxI+tYh4arvIKVbh9DACXq+wL/d4fBt
mMb1G3bZi8CmncrYTwjLrA1mm2MhkKWkMf2EiLtbocHfV03J/iThG6wx6siXZA/W
tLrICfLIShyUBQ3kEs5ZSPhkzasS2xMdbkQNZaSrUxk2fO16mACNtXW418F2Ey1p
XWq43fijTwRtNZN6Z7/a8eoMS/bjwnz/BYMje5+8lsmFK2QM5NdNui8jdNPwZX2w
pIOvTwm9H2zeBcIMIA2HpllvE1JXwc1ppltIOhPxkGafW+u9uWiPnU1vX+07J3WN
S+oc7d4+UYZFVV/H59kwn/sqyJSZJHmmtDg/3AKCRJhe1EVPNsSPGGSfiztx/Atr
BVcQYWUuN/M7hZ0Gti8pUDmNCSA/kuPyvtHRlT8i42qNlb7MMY7piffNUJcS2wwo
Frn/M3FnBwX49XAdqAz51Hj50vdsoGnu3skpYP01V+TBRhmp7jsUrRQ+rIGUSg/h
RaAmH+rKSsNWrgmIeGD2yezihHDoat6Oys0IQtbZRVjpp1XOhBsR9uYsRo8Pcoxa
5UAgRhpgL/uKjk+SLKyAwl//yMOY7EUeYKr/h+FSzwfXYXzML5xyRdcLmMyjbRjQ
TEVGG/EP7iL9+EF5YZmOC9RDmZRQAmAl26XgvibrZw39jmUQ0gH9ZKOD2VP0hKY9
d1+SsivAvGr+D0+qq9m3ZpgSPb8H8H7Cz/ElluwPOdeNLUzasF8oBrXRv3y8BWEv
z1V0JhaYurXeBtZEE7EZyk9TEWtEGx5rAd6cDFMyYm4Zgi90Evv1ne+SHd1dnY/6
AYTqVL9hhjuAhc/fcK7QRSX7Ypwp4VyC78mVIF1IYYlMjazd4SW9n1xKDWR1NjFW
FOZ84XOn5gFfBcfxuN+z7+gu8L/IQTmTC17kYVXlgbSV5UiuOoMgSfpZc2ZaSXv/
sPxi28s8EXkKoYuul46ssfjKpnl1EvepZGDPSKRAMYJa7N+cYwOCVuxD4o8D9yT1
HP+NvArmK+ht7m/XpIcCWtqzUer5sjj5OnbMwSu3WQYonffBIDrkLy8YAOcrowH6
Q2ER0AXMVQrqD1SGkHF+8ABiDNGHA+1J/lQ+dfM81fCm5m+43t5k29TBw0HJgED6
y7bntExt2zpHTBgJgBsfa7oBrJ3uDqYbCDXoGGLhW6h5AZ/QClkNnyrfYO5H6VmK
gOODxVbdji7dEzQOWW1CyvbxhOM+zWlVzbkQV+dqxsR/NRwi+wamQWaOm25h619J
6+lANTWM7hQGNjR0E6Dz1DoH1PtqBxO/I9g0Ci2bc3KUirCNWSK+V2Aj+gx6EBj2
yBA8Q6eZ27I01YH0WZ7RM1AiLuTm6RTcwIyBC0jeAmWFQyFdFhy+vjXLir6mKtPZ
ALugIT2Ww+JLKIO2w85/Do6r4BRyXC+HWzohyyHNX0eEfMPpyvzpUa0Kaq7+od+k
1OhBIDeFPmGELVM0crmqw/iuxkbYnmicV7UcAY11rsBsQI7uSH+WYtF78UTYX8c3
SRFJE959kkxa9KGwmdjOcFPPyhohPDGuYSuRnEQApP1cmYadTK4k6wIIOzKxLaAY
j3hSZErTOj4t8SP0F92xjvwn9VYIZxZMpw/XjyV8uWEYKkeyUhxV4JEpn3HMHN88
GICsjulvKkwlI4j9bs2ZO0sLMB/Ct7X+aGRyobu2Ao19pzLFa0mbCCuSnLSCz3I9
Gxnuk1x3fTWSw9fCeLwm19ACK2NbhSCxuAPz9xZ0l9MtMUPnC/E7/Z7+axGuBzVl
oHDhhT6jxKpeHY4VNkIjYwDeozQ+B1JIsLO5NFa7LrE7TRPbhAHhCWlGq4QHagkJ
2pj3QP3GYXb49qexVWNka8ANkRaorljmmVkv72Y78IiyDQ84hrV4qb8Xff+vERmA
AXub3Hpue+mT2SnF8vCM6ecsJjzE4i2EH0tH/xOnLEvkpfMGxIMfpVtj4tGFO5B1
RntqElaEgjmjSBYXYFz41/4P9bzL5ZTllftxuPgf1eIycF15+cFrSYptasX8H1LF
BwhVdB/lyryst9N127bJnR3xBUV2f3ON0PrVKlE8fsRpjfxhWQVeW4X+JZkJDbD+
qsDZoXkrgUO/GsbegFpVuAeXb/8mTWBcy3QCAO7xQschH6UGrhMJmB2a2HUs3PyS
Zl8HvlZxKBzhuhhqaNazC82Fa1kFD9C3olKl5TCExNU3tDIKhlMpS+pERf6uKzgB
K7QNoRfMS6QuKaEYVQJuaV4/faq3jR54r9Ft3joS35jcz0h2SoNoEV2/nKCkKn3N
4Mk/+7PjhowgYCYBocvLYRpIxH6qokgAUXPMwFPbp3Wy/r0mJcGZDR+uSRBkuO+P
+bST8Mf1s5seLo7in2AH/lQR8T73//KRlbPtYt37OmMCWBYQFsBwMbvQ5sSCOiiI
DzNCo0p6aYwaiPXFvQty8rdCWMdqMBmutJ5ih6k35wvwGKa2csSbqFgaENlt37ES
LpziCRrhhZLm8bhQZigxx8mNrpZ6DOQHF2s5yCHz9yvZ/G+7sIqVkpYHnmKYwdQD
QZ8+ex0lj1WBDzFT2H6nBYT5+1zyR6gYqo2e49QVcrClZ8Ok4CkJGtIRAeo5+8Ml
2Eh/6eLGvuOYjZEANEWIO7vvx5iAytdRcOsUiXz8OjL0kdIhJFCAZ88MXHnmQike
XdUBExVa1nkYP53Ji7cNCameFy8hvIdDdp78Up/y2agRv0EvcxamAcscdC0pU4YN
aqTpj61Nj2h7IHl48GT7OPDvUF1+OgrDAW3LaUuUX40SV99Opj5ChQJdEGWN/sCo
Q/VtsOt1fKrfsT2lGBISaE/9OjBOSORFgrhmtgBuYl/k+Mq0VkzBDjPwuAmJgk6g
MjCYMUnMPJWLfCQK90Ev+WBFl6wtAxlzRONl9YBSS7O7k4EBn40ESVMTfuIsf0Ii
khCEx3ImyduCWsvvjO0bhLEujH+fVYjcrCqbVeCCm3B/SRVRipuuHknj/F3BqKVv
b/NSdRlexV1CpKpagGhVgN4cCkIE8kKx+hzSgCWsS1qKjMLaCCWtxTTn4WSYTx7w
XsBUMDcfsqhEGOpHPpioa6fLjojlWT/sT+fg5DXJc6/5W9f9+FaQSpB0BNcHR6DU
Pw58BSpDKKV+xKp3AVHKAowfNhq/QM7U8LtBcSyeHLzLxb7CQ7DoGQikWZTTZjjU
1KV7HrZT+QFD16HeEEi28BeSEgD/DLoX596ogHcA1uJE4msJuR4hYOiI6B05Ix2r
nONrg65G7lm9nVtvPQqVWTiIqL3IvA64EdZ3sh+GGygT+5P1H4gmpUpdE17JPUYz
hwnnGgmbGJu+XVxwUDUM4yNJmFnwPB0Hr4GHqlxN4I4mPuWTewsdTzTK48Kv+BhA
aydIfcpTjiERuBIfpO2elpcI7IkQ3rBFLODxvB88XlK6F/aIS71i0j8Cu13/AX59
AF71yv23gr5N6fesIJzDFAMDDS2DpPVJ4otVPwMyAJol9eXueZYjcNH6q/U906yo
LBlKB791ucwEGLHg5vIRqRpLUPHdVzBkHrmz0QQZUrti15ylUakEQY1wCbeTGF2K
w0Di/ItvMvFXWY+eL0lfzft5o0SWbnmhHFphplV4in/oPYofdq8ZqdxcSo3+Z9po
YTZ9mFAaLvU+blLMN6VPoFLELbsnKkAKT5YaWDfOy/4ly2AyDcRAXBSwlLuw3yM/
N+UmlEZkKFhhZYEBwzrxg+m+4b0+2i63LmMFrJ7bMSaQwGXEtimurrQjHlfMa+RB
Mw1rJSMNhz+CuCWUQ0vfCd73faGx2M3fBjgOjsKLzAra7MgjDVosCMy7VkFRBcpi
EON1Logrc4kRyeSGdtd+uNGcrtqf9VPbJhCRpoEVZ6peO4ozphZPT0yQ6DWjQv50
y7/3Og9HJPGGBEUKscOlVQxG0BY+eLI1W55NYKDPYqRFAjW88YLMQ5B3cint+K9s
FNNyPmQP0clSCRTbfLfazbz91cgxtz7Vg+SaTFnxwECLtSEDsX4Ix1YmoyA74pif
qYEId0ryCULQ+eHq8RkGPKEBIOpdgokD9BB8yhtTuX0S18X/9W/QHB+R+679pZyj
rfbHb2LmJ9Fu9ORTR3BODx7u5wZ8EFGn12aU1xbNhbfi1BQJ91KjlCTJx5iAsJ8L
vvpN30xL0mMmYJIJQFFqLQ47AURvEMsSudHk/6CJHKOM+3HWRqw+yobFJk+Mkct5
F8mlvA6XgIUIyF4I1HgsDgHZXIUlJ9EM7q9HxonrsbbxRoQxS8ZhyTBA8T+C0rYt
L9XWvAJaIcX13uS6SbJzy8yFZCxkYNiUfxkPWRJ1qiPF9HqXz+1/xaMIm4EgvMs4
qIGt9I957QJtq7JmlYtUqsHBiLwAO58HW6xF36fXh11gilFMALagRdVC1b+VAUK5
duKaD6DvhFqzdrqVLMib7hhXyaqNBkm6sfvshlTWh1JGfU32+da9sedGJUjtAmha
gvJGTKqVpm1qIH2my/VvuBhMjm6LnF+zsRFtijUCeJgeNQV9+2gRamG9NSQpo2ks
ir9vPhEixOFjE9tR4OL9cLCj8kPyu9H/5PAswcxyMXlkgztWnUCqja8fzQwA5n62
vjfRtBRLa/JZTBm5qWxdBoygm0c38vp9fcfX0RCgKccDumhG6c0KMJmpBjjrsG82
ScXsGLZ0hufUHSeZlnCH8/B21sQy9k/sx8Ht6tPtRBVQFY5BOvfUZ1dmXlPXJNh4
R/USrNfhnxbGr7o9d08uCKHdYQb8lMhXPe9B+3hHc5Bswu2f16xT168Vqv4eLr3l
AxtEgBxoWqxftY9yDxUfLppOF8haistZSzJ4vFIxxTFEIjKnxfVsLD/JAJfnGlvv
pa/jD3/U+sQsAWo8xfHhlVygbJaEWw87B7vJIlKkndteIlArWh0i3Kyq9HamKVk5
phjZ9fKuIR6BLgqJRz9ASKnN5ZGxDBS/z3X2oUpOT5JcDom2stWWgNQIBEo/fllh
1Xv8FlSXuXsMSMdVXOsdLLvVM+iO75UQ0VNj4TwgmJihfJblwE4HD4szKHf/kY1j
6LAJKftHo7FvJLGrqM9d53fjv0J9+wiccr9MleQutznLoArICJkcM2FSvY2xOqBY
Mo02VDIkNqJQCJwFS9cTbLCuSnct441+8da45umB/htoE5d5uxKxfSzJyvUDTWx1
M7bEd1fBWKE38/3jTnTUl801W2T7R0v7qZBKnFVWQFOJDrz2Ze1w11CjxCyTV+z2
EacTj41jmabwj6pjMglGkHXIMNMCxTY9Wo0Xzft+b/nQ0aZXMUncDYi1e8Gz34Kn
fLvtHXHcfvRIXb4wfvJij9eN3hYpNnmUYAH00FxqExd9UYGojoTJoayerOSuQ1TQ
LsfuoxoRtpP5YlnIy6YTtizSciLK3fM1CiOBV5pdwy6M1yi2FRySRPR26oxFHcTa
iBA3H2yR3BS0Ka1U5gq3pukxnEegpAC1K7Owc3Rk/yYXiF2jb9UOWvfpn3wdXJtj
+4q5CXkYqqa0VUiH3jqTmXgPjI/qzi9yl/1E+E1nYOxusz83IGvaXKHiUBHfI70q
gG3vs2SWtH1p9EdyvOpRbWqD97B2uJYt8F+SgyOt0m5bym2HYaf1UdHsNm5Q4bTM
BlxjCrj6JL2EehKiqEEVyiAuI17Yt8WdlsrHMnDgJF2HrzHW5GdpUJAd8pCgdmzW
6fXuYLxnq3x6suJayNytAQCIfFulil5VutzuJCHHN8zjPX/nMP/BnPFOqFuXvi4N
47eV1CsJcHYwlojGOhJRx5kIt/7enEBtvM+ybPVcGC2Vfriwv4Oy87qjZkONPBk/
iTBPw4BrwtBGhaoYYZS/oeYh2vt+qudZUpW3zKL+EM+OQDT6112h+k8yqxh1NfyH
yjvgg5BEkv58REYP0Q5MXQtrIDGwkV8ylr5kuD/DUSDs6kTETKHad6gmOMHsz4wm
i5TzR6GSyml50f5AiknHqPLOEgHPXsp93dmJuHTxe8wn3eJZtxGY/awkXz7Wcc//
1lNXn1xwiTn1S6duI4dVfPEr0+nIr1w1QpFrrJjfji/mRSChNSgA/B98UeIw+Nje
agAeFusxdqWMrkAsUrR4NcJnCh7iwpODGy8pZOMAnrWd35gYGGDTdzn8IjWOozgQ
O4k+ftQnyyALGD+SpzL7WGtDeKraNZDW+Gzncv3ByEORPAnZ3HAzVPE+FUFpqNJ0
5R8GscSyalzdRn65jJIAi7z2HbuKRXThGXsis+NWnG4YVr+FchZiT2chPHETYWcf
n5DqumG61V96p+kVqb3d2Uap3mO29vez7RJzDy12e8TvPgmod0xodW3ZY6WSNDUt
cMCFx+t6w0J/Ec9IdScQ9ZsKQvW2vofjFbpBBddjpi1B/un+nLmTDim0YW7EUEc2
Yzso1zOcHeMlO//tXCGREAzD/R93q8Uki4AWSt8dWd/7sqicGRkpDiXa1SE3kUtX
9IciHz5DBR3EWBMGecD0H2bVfKB7bzRbm95IHcWKp2VmloRmdUo4N/Gri6aQPV33
nEF3BJa7F3uVIkT5qoFSYhcDpITmE0QByNtkP/nrIXzj/DMR3Nt8uSzX3ofcqN9F
4Jj1Hm3aigI3852cyPQMelXQccsRsDBtdf6OxKLYbG6PhNnvhI4PGXV5i1qCCEmJ
d6Ti7w0S1wG7ILVR3PnmziMEsswAwZVeFLCWVJaNIgF/ODCOGSg7Dp5MLFx5hWzY
Fq0ABuznSsg0IqFd+R60dotyI+tTrIR95vuRS499FqPZzNApN97i8qjqYn8s9DUu
ORzWiSnPLvmHGBc9HcdS4iTnGjGBg7tpHADnnbrB2zLj7uhcct7Tv1SmSZm4Uyyi
cS61d/+IogbvmXt5e65JrZ4rV4gCqhQxedMBBd9EVOJ/VMqf9Pr3psoV34NxphIo
ieKkm8Ad0sscSP17Orf/lztjxQ8swQ77nzbMruGrdflp9pf43wzO57g+6dLfkaHz
3knSH8HFHxCoN8cDUtE40jReIO/Yu8oBPrKR2eClcnMA6hfcwnItiCQoQryaxFIC
RlPHb80Zwyl4fZBJHsT7VmI/LampDdw7OuANpkup9Orzgj+LKD22l+OhXBUEh9hF
dW3Njdg9+NoEjm9xuN1yhgSALrCuVukPG6iEjStfDBVPiUE4buamU5ggRhf1CSbn
VWlau/RX/OlnTkBYFtnJimUySrIEZX7lFOfiB2c4gp+3jT+O8QQLrkA50PouCL6I
Ykay6Q5gJBC4+huBboxEEE/8BmAJQiceNUN7w+5tx1Del5jsJ71KaBk1mlk9d+F4
XDyxI0CBy2pOBbqNzw6Xo7R737YJP0q1E7eUVyvJe+6AZ9/En4B2Yw+hR6fijq5X
UfhKaEYDYNnmq3Dx/RjDwcd5IeUMtfW9xAjn7dwMbd439JpMQ76NnFgco01RheXB
5KsUhAhzZwXMYFiJrz1vqa0LEsM4fK85r0Qzx51OJggl1mIuZr4RikSyrTyfdx0x
4qDeQNiYqo5WgeBwwD1CtMh3yo6UuulES9t+DCXPrktfG5roGMHk8+TE7iDuBX6u
/2osD1iCT0HbQMk4xFfbVV/USLBZ5fCh/z3XKu9r6EXS7iBxBtbqA5SlI2bNlzUe
1g4wQPlvLlQUhrCRwPmpBMZ6MiKjRFLlrVpbI2nTER8w2tHpjLkajReTi/6PzFfy
XTWATBYJA5+1wKRMYWwSapGCf+zcCqBXmnxp0MVN+x9mohOMYe6oPdbyt3Hd6vWi
0F/K3bOvOBwaL66heyXHiPviMwUqqtO91bJLEEnwXWkxINagBbFE9oo9BCJ+rv8X
/m7zuB+pzrMlM4B/6Ayaqu3ACpPuw7qFKSztdHG1nOHHKHfkGvEEd4p4+r624g+k
HsoQq34mDyG9rfGcYxwU0fBUZIhY5aXZZ7moYXigvvcxdz1Ha83pamY41QZsPPoQ
bJe/XrHiIO/L4CyYxivff7OFZZn6rxECS0dqVJqiFrV3uRIbCjXeWkRxxDlskVtx
FFTrGNtBdunOUW6fBbzbLtYrzCPdIdikT6lEU3n6et0aqOnktjz2ziMT5AlhZXfo
shmRjxt/zUTKJ2+BmBX/pw+DKPk5QRJYvUlFxFDK+ljkmYVVXAyzYeDLkRsfvURH
RUGOJDFsMjbo/Qoh+hbmaO8+fnUoY9umULk4DIxPWidwQbQl5YE+cY1rEygFDDVA
xSeLAns0kVRHS5fhRf+K4lPE3BfFnPVsTo9qwbVZjfR9XXvU85zosdRnCwmxXUOh
G0MAEtKLNciP0HjZAK3uvfNUbPet1SKqOVEoTXnxtpuNuxQDYAZjPeFbjW5XPGwC
7tqINLlhnMf5mEhAxe2tRI5nLMhEIIPHUgnLLi8cbiFLbSZvCIxQJYXf/0JNz7VE
+qYwQdzYza5HrFHJxl2YYyO0G7tibQK39b8PCk5iyDascvBuOSQnSvLlYaZcaDuv
gj8Y8A16+JeWBIy2KfPByhmYAjGULUgDdbFeSxTKy/+za2i90M9w59QBMmsSOX1y
X7q3g+9gsnbcku26aAvxN8B6HkJuOzVpdKJCKhm1PdIUjhW7zrNd+oZyxNf8caR0
MnPOXRbDwLM6rkVwXliVAeplTAAP6HTYK3rkmOwW8t955thEtboulhQ3aOEsfL74
BOZlP/9u8urHMyyX8P2choc3Gr6o/EDpN3ThbcSJat8H79UWPGMn0xlUp/QUjq0M
hFh9+ahL+PtvcwIgQtxezljAuSyhARNBc2VLhVevbtwbdNX4sR3gr0P63I1qW2QN
rkx5w5XFlTfZNi0LdcytB5cmzMkJhYfkeJDz2TsCqbZDjy4P29dIZK7iOG6GjlAc
9hmiKghRzaf96GSM8r36SaKUEIw/8NRJYO8sChBuQvi3zboL9+DYCEBtr5eT0pyv
GREkypoPQYN/Mu9fjnK+tqaHi5ZzmBLopO5fTrY5XC6HrtJZi9FwgISdrNPoizf1
ZdwBGC0YHaQnJVWmvNTrxnrQbrGK7I6SfKxRESnbBXg9QhY0je6FPxPqfYzWkOpc
7y8z8hpC0c8G0vxWqfEQG6By755gvrGBagZLWm6WhLnjd2qxujQZQYUvxnYqi34z
FI++MCqAx+3yldMyonHhyTmhQkPTezshrhU85ht5Fv3MkYvH2dMPjuOut81rtWDO
JMnN6edYZmAaCXSlzxmdj3/oQCGEonkA4ieKlVua2awdHMilIIHVkPTWPTSvFueZ
sCUMjCiyRqtRm5fld6qZp2Z6zwerIRMd+xwD8eK8oHN1KDxE+GFDIyBUYFZPEbWx
gpHk2dpBQ58yeeTLUolJbgsfpFKZe8c+HkMeirJJUkR86OXjd4fzxHJxpblYid6e
7zjZ6zquBCsnvOpGwZdjnuY0+hgg99yQWVZR6XCWq1tzFg2pu1petUKIXNu5KWQx
5gzjEZ8ypk+MEFxGo7q03yYvTs3PS+XjTO0Yqfzkz9SvMWKBZBPXtRleCd0d+WB1
sceJubnTM/7ZkQ4gyh8lMBRrPPQmiE1Xk26Ygda+0ihk+vQTmjLalai0B4jk5R7D
2nom0akf0J9CuvSQaBnEVAWyBIhMJXK3CpXs9qfFSjtBb71w9rnQTjuSxrb6Ftx3
NE/V1CJ/wPQmcKHleoUREwGt1rYqx1RQt0P9h74UjeCgYctkf3d0jv9Y51QbHf2M
9ZMB/L38jFryrnWCvb8HfgFwfzGTYa5Hm/Z8ZOFAaMhsW0WDgw2o/Q4kak9ROaYI
qt5SgNZWhkfuhcMrVyhfLp7VGI5PTJjq4rwTFORqTd3Jq9yJsDjLyEQC6F4FVuKn
07hZqxD5LloCXzcULfX6+FCfosv10n6mCh4kXTn3DaxfFQ2IGtViiaQMezlEQzdl
1TehxJjX8vovet0TMq7E+igskoEjDK2dCoKUTiot1U0Bzyh9kyvgdTmqoUYFspKJ
G2SACTV5C07Nd9eWCpZXtN8FZtKaOThbzd7iXBbUmGjuHBnCDxuYbWWMW/W7Me1u
/QF/6sl6b36JgzCgwAn5WSmWXRZHzJIn+H/2+zXpIFNKyMAusCgXaUN1zE3gpf2r
j0mj8VC8JnC6HT0EOUuAP05dDgXecGoK5viAP9Cur1m4ajRMcrzA5owehj1Q3ydw
GGeo38C3niE1yVpEIxuRP0HuT2u3f2gUv5KboKd8T6kFrz2K796cXhxwTsN8d0lU
6Z6C7jPZWRgJxAfTASP1XRd1Lde7KCfyVOK17W63oSc8RY+ascBjS2bmzNG0QFby
QmN3JGsATgEicld9lOAWzDNdJ1+4TLg0+bCcEFQ4AJxFh3Yb7I59h/pHsLKREjkz
Wr2G/iZRfXS7CJeSgAELWzLDnNs0Z7lkl/2by6b4teccK5GTUb/BVck+Jx8llulj
175zb8DnlUYQkd4AQ2VCU9N4vBov4jWWGxO0w98D732Uaosph6J5KutkkpEqeYDl
8wwlfBlNqxM4OGYH01xqj4s34vsun48rIQByxzqcwOCiPvV1l50C7w4WVJwtw/Vv
CYAxIwBGN9NbfVzLWSfjJXzgGe8EGJmnoAjYix40SN0lm18BC1QLPqw7aHZEojIi
BhS97xuuFGJhTwfempwj4pG4XGLMCGllfBzLjLm+yiniQRH001gCcazE5HC0VUST
QCloYoXsGfpLEH5oZzXFthagKdjR9Jm63m+1LBUyfqvvLXDNcpF5UWhZiXU32ABH
6k7X+ZhU++1u/DB7zACchfR6CitOGXZPCca2b333IFHnbkBk1rQHobgfZcGrQeS+
CrB+UgcGWCVKfMKaWHttMhEwZF4jZksiSHGRtW0Pt47AcLhcfrjI8+xw0L1o1if0
1cehyv8YRI72JWCDv1qL7EiRlgQOoO/WYb1UCzIpBoYi9ZH7GEXlZIqzSP2K3coz
/AvayJUBZPMilewx6sTeaHBVRKNj0P42iQWwc6S/si6XFTi3IBj5KiMAFkE7Bz/6
WdGkQAzqdiP0IvPhEFa9UIg7JJmm01KjBgKzx08bqCSwIg8neQ4dJtcmmA3u1SrD
paJ1lasiOwUqmu33xZhhStFb3uFgmony32EFdjkqilfMbzp2i0bkYGaQDwyNUzV4
8o3gN9rkl6w4KOwaVpBBNaPoeolHZBTTKNoR0Gjc42hrPembk/EU7ZGpJV9/9qIM
/TuiUinactjYGXRbHwdZQ4fzEi+JEJZL7n+bQvCnY5Q7DQ3Hye5X30pms9syP7hi
jYrBNZX9okPB84PM3gDjkJoHxHExeOx+O1FlTwFj3cikZD/yReXvaWezJl+zEqeZ
WpVB3ejcGJdqH3rAnNU34owzDnEO8fQV1FF5Z8nrSMXeI80T6+DGKHA6YqCVjmVR
42x4p4dE1ahox1i0fMGPz8xEOfxvcC7Co1VBWWblfPk7euMC4Yptaj9VbpryRwkx
7ICu9+DEaYVPP5HgMkTr+u6OVz77CAExkQOoSvnCXHowDE6UCLQGgwA6S4vjd5pi
bPD54+GmNqhHbQZo34+C0uj0QGFddshzPxoHjlc/yRrzhxLA2TI9JJmtRpK4GwRy
M2Ded2hJhgbTCCeFnhkVGaXD34oVs2EaVjH07NgXOlYm0RJXLWXcUVC6/OEwd2EG
8eq69c/ZzmqW5xNdRfToNzLWh1FSA9rc/NsKVnQ2k0c/lsOBsHo7+2qjl4lOfqI5
KX+8TJvvEnieR8gGhTwnLZ7BLx4IVSgO2yPmoDePT44Afqm4JZo1pzOmN4RRjaBv
PE5iZD6p/sOBUjNP+LNqY040yNEI18RQuQzhUOogCRhwBxsGVds3zFOt0lIpI48Q
MwB9hiokjvzG27gtpWVPmBLV6OKtHAMdKj06inGk+zK0NfcCPhBLPBTjBoZUIrnj
OpFRwI+v7s0MszaqKLnbm14sOMdk1qSW0FpNu2mRf1E=
`pragma protect end_protected
