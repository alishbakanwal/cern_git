// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 13:57:49 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Os0SupmBEc/kEWM0nJJvkokxub/rs5JWuHhG5RF9ES6yjhnZLv9cAZiRJDceAPVP
1RyrFyTGS/uHCfqhDMes4N80pEgYRnwiXErl3PBHzxeaUo0ykKu5z1zcoL3+ECYr
RTLPfLWhX7Qnryb410Vds/cAoIJxLlL+A+rdw5GIhzA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3056)
xgm+SMwlS9PMXH4l+cHqbdNm3AxAze+Lx6aWqeU1fFpDipWVafuEKWDS5CIbBgDq
2udrFCsHAGZLnxiCXH3b/sD+faMQ513bdZDwo5TI/2RoGdYyxJcT+5h+Lp6mSQRj
StA7PKgGpCHtIjGj5Tx/VRFaqy+sLMrg00ugmAGo3WpLf34aWxXFX5YqDoTyZLWL
siNXDKYOsXKiP0Zl+VLjbHxWmymxo7sPFrtbtZh5kYbX7cP/W8SA04MbN75t7yJG
Ft+qNr4ZKhZTMrdNpuxJdSHWGqvJVBLTmG7S/Cip27m/pOnLW22Ejy44H0frNs0Q
2zTW8VSXmL2Eu4zMcHpN6v3zhYAPUHPHcWVKsN+tYV9QFNK55g4f24BYK5VbcLAM
KQFEZK6f/SieA9SpOXSVkhYZzf+S4Q5xJf5FcRUYQxTuCvtkTMtH2MFQuzYD5meM
j2sViPQ0Z70ka3hZy8Eb5IymTQZ8s4CF9BDcGLL62ZRP1iFh+BCJ5Ryc5jiYLfhf
jMM1NReAl0IuiuoEekYV4uh49FcYaxC6DFhK8snF7GPv2DZBrw4dzM3xocT+UrNi
8u0C4TLkFE8oTdlxPTDzkeS5P/bT+/86BeLCet7z5ebu7rD2LSO+jOrYQzKqzCwW
jLRHlyApwgNnkfr2KRW7n+Gp20olZYjQblm0ENqRSPY7Dbi6FjN5RklrEMGaUt3G
GZVbz6PdHp9an1Stwp92h86AASo75qJZdErj9R1/QIiPELhnBGHA+aKVtCmXkyS3
NoyIpYmJ2ZBcK8F8X/WhzFiBnovikijaWK5HVF8UCz/ILQML+ApJ3rMdylN5Fi6o
Wg+oHila4OPHNpN25k/EGxrNOHir8yf80JVbmeSaTtYtzAAqEqmHGyJ1vZdi12SR
FCNrTgqEuqeQE6Le58b5gIxuJl3DQzLQKguYa3pfVUpGUadctTLcbkc4WzPky1qL
BNlZp1YlY3kTkoZ6i9gdOPCGkOJ4gyC5pUiq20T2YrI0lk9zLgZgrsbTv3uqMPmC
0t5kCvrdKMMH9SUiZLKrClyDTmTawxXFWw2on0I4xflnQaeJx09JMZOrageVKFMX
WJ+idblJcgc9QwRWp5wbrhy906SdDfF0Gnlzi3ouIuuRA8Pyqk4z7ZpVrNhAilza
TGFvZWi1O7OziN+Wxw8CHGEdHkhE7rplEvcGvfmnTnUwOJtROS4r7T8s9fj2ZQpW
h2Bc/3GVM48vSDkuxvr2+gEeuoMO02KjHjtxFHsldSmvHbGw/Cn6VVtlsVS66CqK
RXZF1954AUF2IjrBck1cIprQXr4csbYO4Zurve+z1+5tpEY7UBf8HZ2sIL3rHsxu
aipyVw/dTfURSq/awlbeUthu++dI1iSU7oToNB77GRwqSpAqTeuuu2+ZWMM2+i7K
wf53eVNtK6C3eCr+JYMMD21i/+Ei0xnvuvbzNaTH9kooo+8zDQ10hfTansYN/SMI
o1qtouUnyOe7Xi4zwGXCOz1MFhr2ln8C6OCLiaeBu6LPz33uFVA41u2AV8i7orJa
valleS3IRZkX0H8oZfjWQE16EhuI/qwskDdF9XqbCKC5+mpw6XqVihs/eHX301+x
XpoMHxPIxH+Nr6svWiRz1BlySsn1xc1riQC1BpfGmMCSkoMHx8UwQ/9HpH5fNmR2
Qx1sbGddeer6E6/+sDk/4Y/Ls4sDQ8SdEUHXN0URI7un8MwOY6Alw3nk2OFr3DWB
CUe26BhiDuyXRmuWUVtkO7/sQLswzJ0YFjPikUd8TWAs/JgbhYuk7ETSEO8ogg87
yHC+AyGBxsNHwY7FqtU98LZ4mJLyPDVq01vWeQruROZGf63oySAJeawyognwrWil
3w+xouPtY8FQVSMh3On3x9sZwHwTaY+pn6VD+phQpV9VK2hXWV8LyazBFPT3U2GH
ncsy+I/r7GdW7Pz7I5ROkgMXTMfM6Yk3/UMEejNVCN2sLa/nDwghwzv1iy5n7wZs
4rcb0F5xYvaqK/O+XSEKn5hdHR5eM1sZLpaL1RCJIL6+WbBRGdpHsXs+fsDdMB3Y
g5/8NIuBRjXCTCnd1cgvMNbtqOTCtPuaO1WMzFLd1H2iF/Aq7Wkqm5Q+Ozk1gkm9
vyFPz1EK5mW1hR8+4shfVbUgxV9B7ltkuT2bFka9KdqqRxNM9alBCoi9/fBsZglI
dLf6WP1xVFE08Zew0tjEcMso0empzeR0lU9U83rKPscLPJCHWYxyBXG2CsZvvJJN
TwKNqArqiC1qXZdRTJskxZJuqrozftPtRYkGssC6mBvCQGVIZosZP0dnu6q+/e3U
vVWMhs1g8Pr28wNdqvUl/TKjKo3oOIxQSx4bjRmsgJ/Wl70wbGlz4BtAZLNBrlEd
VukXWxlzp8S2yEMiBLRAALfnOhSMWLDDYEEgf7lEgDIj/ygVWtW5Le3IJ0IpCYBQ
VggmgPf9N+/kxo8iOyskCWWi83cLQ+exp/IOgeI9Se0hyFmCu5ZS3alVgCk3mipq
oNWyiHqPOLlHUhwiCe2yx7Z7KLGnXQ6kIhsfiU73IWSw+npQn8o2ruHmaYuvoZVU
QEPVSizjNJx4erK/IK+RkDzLnSHVgExooH8Du4C+e70jjo0KJM6/MXtYj1cy/RgL
i72TZHRy/UQINSa8POTy9825LzouqDyOwSV46yfiuQWqbM+5TAJsnZw+OMV4XDim
tN7diSfRxlsQjqLHrgzeD/cmMV7LwjdVbg/mmdCX1MHLIQFE0lT/Wvi0TsxbCqEQ
Od0BEdriUgHVvETQOizpohlLf/bMVkNCDY4ZPY8P9m31jkdD+/09nRSudhF8jgLP
EkI1LlZQSggm4CSalZoAXixg6URp3cOHbPHCCdcWRoMUOFda1NNbCPMS67udONZg
pRb+o+SWb5ShPR3YLykTLA9Na3m0IMDfFNpE36MIJCasUYDniddJoA4SX2z1+Km/
84HTmWieYF5vLNgQPmWiahbE63wqKpS5gI73S1zRS63AA6IKunaFBf27MrQmieGg
kc15abl4G+uixjZEiXwAsmRVuRBitEUg01uzF3DhXNqk1Km+JIXgtF0pA2s2gFbq
kCZ/NO+J7KgCuvAnAxiOHKQYbVtOjyrd12OTGD/oSPvXw40HYAKN1l7rktEpK3OC
/j806k76kEuerksRXwFiwnOZDREIuuFWQ1p50i8XP5FUIrttnJOLLqp/W5BipJxq
dQonuL2cKwYBCJ8bYOHK1pXmTEk2M2vvyV1PJvDPt6W5Sm3DGuR0YDtO9KsMewfF
VIJBW7N4im/1Xju+2ORTWiJk0qw0jn0v7+6q7NWmgvFDqhHWlX6A8Mo61FQgQf3D
uCu22TwyJS7x18Lx1ggt1UbUUlYgZsBBHXxHL8kpS4sFKzOtMIUWEOdWSw4Fv4ae
Jko6F+MECIEpdNckLWB64hHzdn3wzkTwQWjNfcfUppI9b9iyE4is4MhC183QzA8x
HH3oVv58TpDYVK0vlJ1Clsfbpg53q6XRYFIEYZqNO6iyTAJFBvNWRw0k5o9bb+KE
/aKPqVPZuB3IRDh+q7EAnnp28XDnpJ5bCsw5SSvangTDFxpgl6d5is2mIJQzQ4mu
fhx7V68PMGrMQmP23Xri81Dy7LKLCkidN7ocOqiHX6T/OPotcc0jIyxXLSruoK+Q
dtahHSh238ZHWtPqBQxMaObUIlzkTmg3P5DeBuZPpZFRwzoi2hNbUJS+CLNqQJfP
8ntk3FC72fS1AtqO5kawFPXyPni38Nx0AWQhVPF9QG9GYqRJtMyjbsarA+IBoFXc
W3nOFIqyvXwIbZT/9fRfK/g6detjfyvb5+TGSRhMZzq+58uONUkkrE6auUv6l/4W
m+lQUsSY05i+MX/h/T+FuJZEgqtOtcFbFR5u/rwruFbXWz9U2H7nJqM7AB0Q78ds
1jPqdYc8MVgoIvr2fxUGXaz6XT4wP+5hqak6xP9UEw6vqDbf+mf9AYGfJIgOnZi+
jf4CkOqvLmdI//fYYRsBt6p7XK4AzQiBIgu1noKQUwyN6t8xBdBkIa5KO7wrkDQE
Zv7/P4dzeYFtmoddNGw/07DvpXCYVm2BpJdOmcTYgz4=
`pragma protect end_protected
