// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BI0Rl/ZmIiDMOQklpeEf3RHXoxsZH93aIlZnenCQ5+TbzNwcvaSXbWLioFKRx6Wj
e5nWcYYwgAvWJjuG9xLc+s1F1ejURxS+t4DSl7bsy/gAzikHwKyz+3jK0xQd6KrD
0HMOZXyNE22YT7ukWSARah0h1xK0ayI9/Hdg/Y9QVm0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22272)
m27ADD+O65zh7Qma77HWX/cCxmwcdqMAzAn+ZnVCX/9NwrrKCKnpgLRXpsZCskts
glHoa2tzyrmvlYSuCezhRaE8EpddLFWNgXY8EDWxWe79Fttmjf8K7LpmC5e+vDci
IH+KXA/Ui1tdt4TZtlJPcOH3bw8UsRtUAe8Ig9mu+/2SFgWkxjnzxfoctRiqCiD1
54e59WmD6XqySO++rt3j9mhO4ivY0SMox8tTZANtftnRyhdRG/q6heFA7xKtQDyD
Vte1GuISenNC5C2b1+6wysJLSRa4PJ8ahAenadEv6qaNESqak5KYdKJxsoBgaL+p
1y66GRn4nEoCQ+o10J09D8sjXOjOFftub/pMibEs7yg/NogkHrej0axWzQJk3/qS
j8+iEcvpOoPF2p/JluaFlQQGGjKsXhvFm+muWu74H5XpYSTMij041XTl3lmu7fim
+q935yTugyQH1Tjxtn4hiikfjuZWqQxomzmpqdT2l/MTjeMwR/qjkpRrAlcqLFW5
h1dG+VmHxLFRrSy3rX99OtDpcYbe47W2v+dj1e/xLHjgrhKOOykZvYzZXpNGDxj2
ce0YLRL72yCIdOWfebnVHSH09EhbCouiK9ikCVAICXyR4hEGwEqh5HevKUNV0OAH
5rkoGl/p2jvZAc8AMP7Ik0K4B0nwu/ThcZ9JdkSFs5rP/uLJfMIp8pd3p5bVAlzx
cR2t+EcYA6rNlY/y/KYs+BFn1zNg3sRa/T5/hz2pYgyksO7T9kTnMtS2FMzT/9fD
vju98gR/Edtg/tF8IjtjuHaPhP20v3PbXsyr2fHP53g5X9kTVRU8p0DWAatvQX38
rBH5K6yzWuK88q1rhwdh56lrq4HA+6MLLrZI6eysxFW/kefAgmdH/vL+sFjCq2mQ
Ne4HOaSW08cB8ebFiRZSm9MoF1kcxFIpLkGBY8g2Y2kc0jmUHV85UiPurFtU7Jjw
b2gkjcKxn//O+23XC2bqZQrW52oEPsRJteERG04zz8fucMEfPRHScTPzTYeXBNN9
qjavNSpg3HG1nIO8lHqm7UJs2ig3aAM9dph3AW9TMIN/P5fUm0jXT+HbRU7tFZ3k
2aqqnkDV4IPyNxU/L6EWCe2yBH7C75i0WrUHkOqxtAoZDzmJQy/+jwxQ4XnJL2Ri
772XmwaVEGx0Q1Kg/QCo3VfH4F/liQxiwEGp0oy5Ta+LEPqCdVQFcelHrB0W5eL1
tCbKuvv6H+OhF8Qo/+GO2PE/NOGhaEqlQyZgZ7CDykp9JkeB39l+4z+xbfG+PyrU
hfqkILwQsnDS6ERBdYZdCmzQXQ84GNPCeNWLYJ5G5eXbQSt5qCvSC21Ea/rLVVkJ
+ZTvPpRCQez4VT1ABTWlVqPWSLqVi41v0YmCBkZVickWxZSPC4+bpijp8uV88RRj
XfT5URWwghYADQekb4mJXrhFfoaDF1abqaDNEc8Wq4WNprpkvpEYPW0/DG3V+eF7
xVy2lmM1hvrTzqX77CzN8B+g0N7IX9n0EyzSqbUJ9ZhJx6JyUfpEgy3ExaW1HFCw
3n2UpnnQzsUrTWie5JPYP2v8fuQrkOiieG8K6UYPszh2zT+oQragOsxzl/rL5vIN
bJtcLB+QVpdCaWVHkjKrRjz69SnZ7rJynjkL9hejM0Fod1/rkDtM4IpaLHkZS/d0
ZbhLRPcKLXQaG4oMpUdRNht5Qu6FF9eoysSjyLwlZ8I83Ir30DWqC8iyImSyKZ5o
ByAtEf2vrMtyFI3hGS+FcEt4yI4KqUv8XMIgY2diYGUKvwLJbSOiXG127OUafno/
SRXgPTV/kMzO8eNfh3xRuJGCI+DWiw1TMM3mrAf3/50wIHBRlQ03d4SatqU1Ilhm
k9jxNDtifJ8bWg62MpFF08JQYr05Q8vQITO/CD9HJISoHDLZE6dX/da6WdKbIZ6i
5twbpR5BuaXHUdbvb7HpNCfgAryXHzrL/fhHfp1UWuWdds7rwAjDnQ7PUV2x61Dv
qNv8EZglcbaFAgLXRP4/vAlpCPyCzzedCnjhbGBls85NwNs3IItq4z4xOjgiWpgF
V0m00lVF35Rnmat+E432Nn6iXsNftKUr6EcP6GgK6jdQjXJnyK4+GGyElmcGP+BK
bZmL8dlf+C6yd2nxA0sqjSYUAUkzxkrGMyooCN5ZpxXaRSIFGt9F/uZWVcoQGKx6
IvwmVOy8yRJO3IU+rxrlg3vBCf+g/jtZ6fmES7BUsggclw8+rEqC+AL2pcCczk2y
u+TvGYpzW0NAEWntiBPZ8izN1PcA/vtzIPAQu2cCGF5SnGl55/uFCJvDZWS6/YYR
FK76loFzZEFhhsWJ1V9jT6Xb9yQ/mIVNt8tOrn53f8P1XFBsSFSBU3FpsntC4YRJ
JIkoyM/n1wdgmH9dn5kEFK3XlNmnH6RSejX8+WFztiNLPSSlfEfrEBzsYuCtXbYf
6wnjN6vlAuG6E90a7OWyIb1kb5hgRYm+0SKRSyoBZtrpHYDntKuHBCg77MYOCUbx
pakhjW0mrQmo1Sbn7l86sc9u5LKoBY1lwsA8Cg87OYVctUck3re2qbGTx6hct6j6
ov0CNjCuAKiBvlltKcmQwRQTjx1MQvYqtYqkMv9ZUxoMbTwbc6RwZ5uJj8gGMc2K
fVieGtMb8dl95Fv5CrjBcEHmYgkWT4Td+9RqMyLXSsM9HmOD++oqz5JvgLjJ8uzc
W4b5scBk9b2eV6FaHs/eAlZI4K7h+sucilUHC70vQPT9MX8RxHhv8VCs8O7h/q1a
uoiATF4tgKqTOMx/WtuIDYbH/po8973gr0O1BSxV6EI4YENlAunM8wOHExBhRPYI
hy2kyY5UbcZJ0OsieUZV/tp5IJyRkJD1A8kmJHvpK8nCDRWWvSAz4ZLTSrvOw/yG
so8TYi58FVJvXQ7/yW5c9fX0+fVJZQNvVpzIfg4KXMP+V2HwA480wwgaYiNq0Szo
Vo+hWm7aPmnzu7w4l9ATXFXt/J3Az2yKdv+EVh8SjtNixQcnHg5WPRHu1k7Xb+ef
7XfmR6DRNhqv+fh2LbSOUe+5gSrGsrKfCOZA/gtqNdFCBKL07zSBINo8SC3aQwq/
u87JHGzg1TWJrTVy70fMzK/79TFtEQHQJqHjtbktV7laVQQj1v7jyoOatTVs1S4V
KLCRM04HXmjpH8+s652NALy+2z5LHGXKWjDRroIOgC5Tvn+s0GuQHjMlLHwSVjG/
2TiF6X1xbNnYWLibnwPVHZCxEER85V+fUfILs4Civ1AhOkCrYChywqn+tIZNW/Zg
T+v8LKTcz5lSmrCFqoAVebg+hDz6ySxsdlycj3TICeN4Q3Jt9QX0yGdDFhJCDuJg
1dT1HGBdkitLVikCyP4mvKeBJvcwwzMzJ7oXfknyBI0quywKvubLEaGwVsOORyeW
DJJHSlzqI5PnPVvcLsNRHzEbM+yG5AUKerMLTlnlgap5eYfQvxzcTQ+yfdXozP9H
GXkNyI3dEpSyURtSN/obRoxMAqZBTFO45pDRDDaj3JBEgevatEFuE1M62nsJFpP1
loz5V0rrQ5OvF1OqsUm9gIo4enHV+LyxvaRy4LWXF7dnKHan9X1NMmymGTpofByb
zoYTS1zdZ1YBNQO3iLauR0j/dtsXgin519SrJLsUmfkaAa/ozCO1lEwRrWOGm+gX
c1mEBP5HGBk/pnquQRowC32CIuMF6pOTuUFd5pNsA+q00TJUQR2od7c7R4cvMFWU
rlc95QEgEd1rQX4p7+233fijwIx4hpIrlOVyhl/oKrHUWIwJWymtMqkfMS+g+SoO
sFcW7BAZKFPUGOxU/Y49EXgObVbakNZQ8QQmkcTzz0MqAjU/GVYg7kcFyqM5NAsd
wQTRB5kYrASukKRykilt+pEKcLLQUHXOiukVxo/1um1WPBUR3aVM2YyrxEam74Jh
HfniyZ6F8Myu1y6XxaUhNoTAhXGDXM6JLxGXp/FzpTEoKYYe528u32t/wlIZ1Ytu
ZnTqZtrJ0+SrR9sxbq6oYZuDqb3B8qH9AEkSijiEtADtT+xh94sqOILsyE5zEW6x
ne/NlQVLxjxLRe44L0/ws4TIkddNbIDZ357tdugJVh4cYwpueGfhtPxlbZ8mf5lI
2v2HK2cL1jZaLfFIvSScJiw9kUB4e7ZaReOxyh5U1xmax09I95pEtODDKW7dP4I3
2Xacxe9Kynskqk8L49le88ikmgxE+ljBb6dywhbtC0YlY6NpWbCg9DBTLuWkn37i
KmedodP9/eJl9XeX/XltKxjE0h1TXCMuRRoHJMBE0c0SPBQUUn067WqINYZ8+LST
7ZkKNFd7tPwfwGqaagv60GqhTw4/9cLwNoxEhpYfRsCYrSvqNDr1ZlGl5dR0FmSp
7elrPW3KQVfZ7EYd8cNgVPMPy0vRl1g6Q/iaJPOOQCd65jeJvQ/ShxkwLJvAEkL2
ruW3b/lTvwuOCNQvFALD87vGVJaw8bHQJ/we1KEeGV6grm8Nutk04CIQXyYzM//G
WSnVTnJREh2pZxPDgCF5/MtMEsJ8aGF59B7XXVuRqasG67w1lFKKzAhdXlvsjKLM
JXQSIYE1J4f+LgNt5sriwcGZQ5ZABNrzyhFCz9Vb56B20CvjhsTLANXzNEFkeW9c
3+lWw0pogjVvzKXliSpAYtMWmWFst64lxOuDwPjPj+NU5aSMC5rt8mqgb2StOUE0
91ZQVyDELga4SJe0ONXnvkQ3DC5Vx6wKaWoSWvfhhQwtkQmEeLVrq7ZG0H4OCmpv
mzHWFGjfVOMGQbWOc9LF7zMxOAVZXcgMYtAGdupkDf5Ek4FudcFdcV68DHn5o6dr
HU9HNPs4M63KphPlJMnOu+yaL6pAEYlbveqM3wHCqwz/v8cbVZHenI8DTkssrkEM
ub/JXMM0H5dCD0Mxgvg+DyFjqUdxTXs37zo3N4MAcw0+oY29/8izWKB6jd2ioBNx
52xTB2CQMIPza6RgKG7fu9twWfrsHPyy/1ZTm8CVqf5ryTRAE1VQGmdDzuG8uOSa
ycCBbPfRzRIxEUwCmW4tryatX9xmi5uKpiUIJ8aEf37BvMGzdRR8cZ0DjLE3RBk/
sqC5Rmym5R6gt6cnDBzVVXVOuXMjh/4iLVh0bmy9FHmG1jhIj3s9UQ/cAPTZw9VY
WtFjWHCk9wMGS5IKknvosevm8i4T6T4f/vra4PwS8o1M+X89STRcJTJGfDEfLz4p
/Vn0cw6Gp2O48KQuNsamSgjze7R7rHILc3lpHH+PAg2zO+aWtQPsEYwJ00eNkpY6
l3+8xHwioIW5GPFn8+hMQf3lm/JmvwEPzu6SfreZakNKFtaOWadSdudPwOsRPYOp
H/waffGPKrxEcUXJ2iBYxJEVRhhRICbRH3C76GCC9vRQVVCay1tblCzdkCICXNOj
YO5qtRiLz9Ec/n+U3qVnlNKGfT8T6/q904JjlUZJPaITxi5qM9Q5O14bW8rwSq7q
RFrDGPCyN/q1deezgd/phVjHkxh8xWay3epGVGzXzaiGzuqCpIqKaYCvC62OCQ6t
oulHjLFEl6PV0GsN15fErI7RHayRezp+H88gf5RVveA/7v8OTwNtklU3XJWQp/q4
ABA7Hkw9/reGgs/N5vlPcOR6rfJFM3MaXojDP8BbKLFLF4g43hK9bl6niDl+G4Uf
xVqVI/rOR8rwOqURJBHLu/Ne5oh1D/IrcGPq6RCtUxyTaTTpSIGSH9H2IrSavTKA
eeZ3QiEB4lQTza+WdhbZhSPFDdiyybIh7Lb+XR+t+WCGXC0ltuLnjxnhA8OIY1n4
5tKUwAZPiwPzTPGvlmX5Xod6eHbQTEYOkCRTYy8wuIucbcCRnXIPlspVIeorX5zM
mIPPWultsmAEUkoSZVL5ZjvwOacy2S5X3jPC2zJWvW+iWewOHioMvl+lfx5b7fKH
W1eo0Idpy0eoLVDNlfHhRSEuKizkcKb+wjHL3ftBjinhh78UX2XCQilJe0EYQ4zF
6VtOu6AR4HW/CjWvw5KoageOHKEYISOMYFRO5VBb8TkweWAf37jFj+pmWyPT3mlF
Sg0VihuC+TdIMk7GcULLCtu2yFeOMhM+Er1TwVaAVMuBuBWNV3r1pGWNil8jRE2Y
/bR9mQtzrR/emtu80JpGnZP0PHZMYpffa4q0B0DcGa69cD4Wh0LocUE9BSlcjRp2
+QoOOb6s0DoQ62e6wcM454dokAOOS423wEJqnAateUYvPMeydu7OUWd0FLSkthTO
IqzzRxE0hQdR724rpAG4TvZBYaOtXW8A2QtztbNvD3Tkvdujkf2W/z7z5Xo5J4rx
jT8UYN1rFregbKTmQh60xaafq58B7iAk7oVLPvxLP4tGCzN/PoxKqzdkPhlUtfn7
1AapbpzjaUKaFaldHUZfhCfAIWkRKlYlfc36l+WJwRuijGgMCtPUmwov1H6MkZMs
MrX2wPAUsG8CmB3KByvmDPXNC3K3A8PrglTQLeHvHIB6w522LvglXp3S33Cu8fmZ
RViK6dp7KuxcxvecfiU3qxYPFv1SF6WVRc5RE9O1kcD8RWAtDsPIsLylqgr4LRXQ
QD9Jd2Ja3k70G839JD7h1BWi8XKq940biCG4LlGlZz18I4ELoSqqTbgI0jPVF6ZJ
S0b0Tic/5YKLxWRmm9Bq98lEVH7WYv6dYG4uYS8C4yfFDTNcDvoeGkxLO1latto3
jBbgEF0H8pOznEW5qgQDalfScK/qwvX/bn7bcFyrt1+irKQR0iEigvi8iqsjJ3oI
bNJFaCW/7OoRhSIfQ2b06uyWbBikAxqqkOpCaymzCuSXeLj6uSzLMMX14jEU8cBu
GU8XW5V+FTMTGUy6sDVyPx8dyNEEHmy2Yrgnd51ZXGnlCTT5AufG9OtHetmI7EHX
p4KurP5Hyz3k0RDI/KysV/2X4AawT1yoceMlxoVA9p/UAuUNdksaFQHI3Ls1dh0X
/mmkvz+1GPFYI5Bwbsnpr2ZM8INzUM5nl7uC5JeBlzIxlyl7indurEhuxPJ7HyXZ
2pHQaCk/hJ7tpcaXndcy5E5iFWUgvIJbJWaswiHrb4LunWROch4Pd9D72Yy6CWc8
hr+qx8EVukaSkoG/rRndZ+1rnj7fsZt3D8jATACn1GsQ2LXBsoGWXdF8C4Dr5rPC
ufzsS94kBjGQiwvKrCKE+fBF2o31VPPnq3hTxs3PGLLqkbwGVxS6wKy7L1PhDgNn
hPB2kU8glReYYcKX9ECFkcApdWY2M2ZWrBw2VJVcKbEInYXt/0os4QanU8d8lQaG
5FM69tUNVSpQg1vW6cewo+9HKGcUabOoukdy/9y1pi/wzMC2IkcyaR0+e+L2DYoi
emsUkUfaiNPDysqT7/Y2/bmRd0p+RSAwVutrFefILuZWTB5bH7cMj9Y16uoOV14X
b+YFX84SZtNxPB7lZB9KyWScYo52VCH8KHqi/wdblTQqGkermQRNYsk+OzoMo6TX
LEMdfxlZmUaPDj0uYvEAB6B07UTS0M/0c9rVy2rRqA0T/HOJRBvfZV3iLthBEN7Z
zTwBppIQepvGn5PcSA36+X/0J1fhTSkSFAP3ikj0PscJl9hViIXT+gVByEEblIKl
sAEXJOVrdKpnW7d60eEOD4UWezw0FzThWU9iOH6ycr6YCczLxGL3+IyBucmystaI
XVAXQADdfsRoZ/HzqiNmM3WVBjAlR+AU9EsETCagt+U6tMAZsVi3pQ73742HEIXO
Xz8YoUZaATOnfi3PO9/6zv1ybtvue8FLHG0mJXYcgxvO+cwOMjXW09o+X2/4Q1A8
Flm7SY0wvpikJv6HWdjZoLCmsiR/iGbX4OjTiksoUOIcJciaPzMxgm8U53W1ckC/
93KAOVVmZZP8s8m0LkEXLUhRA8pZomMsD5vA0B/wnPkFq9x34czzd/P25m5WlazZ
GFzQ5qtWcRHjrjPUqdydvSOUzY/YHYglaBe6hiOZdc+vw5kgX7MTplqfh5HKHZ8/
A4fjRlP8JwYvgfRc8vhYF2Pi/sYnKDOhHdiFH6jFafmk4CY7ZZzvNdsyHGPZKPZe
VoE2h1R5j7p5ANHM6LYLid8WK2oGt0JczKFrKRAs3ix26qCZGJRIE+aujDza3kbu
iokdkrlwnwg2xEwQ810p6JG9Tt7pyZXqVav4ZC46KI1VLFMrYZ3/o1EuHBZbe0wo
zp2Pf1mZAZIQ2eC/+2AbMdwXeSgYLcCB50KO5/zYyuuSV5n/erq/DpzmK7PzRAnq
UcJhPpqm+Og46msU9SeFE0EY+wk7aSqjBil8cHLq7KubgtjZXoBEItyuvXn/9OPV
s9tU2GcNVgwhXap/N6shdKJMlupzcJtLhRMfMimIl6MCVvyevt5m8jGFyM7VClJ0
kMxtPKUIdhTCBOaFZ7BgyU99oDJtooB17NKk0ptGSwp71qDdQ6IcMw5iS4UVNmV+
0K3YwVIbVP/4JE9NeJh2UShTY/7uPwdpRbZuKsjy83iNgaFzLzvlvouM0PLqjALf
bxY/z3ZVjGN+7H72PBHDGNfEc6PRS77XwQbNGdU8kRLFpfPON8imVwmcdyVDckjT
hsiBKK8Rb00wrIWNNxWobjDJX6p9vBr30DSDo2gSOnnYSr2JPUjX8CH32GtV2cj0
0GdCcGbwVLDfeWJsVFikUQ0VwwU/QqVgh6sovLp95ESqPId1+wiu5dj+WDJUQrhD
jv1ITaQeHiU2RROHf+vhEedal0Are49IWVQIH2cGwrrb6rXiP4MYozK4/t/1pRD2
fkr47SreRvdSWYxK6Um9dvmObvsHvykYArRh2s+MSpxUKvxcYeg6X5/+pJowtDfI
j6JJEiCmrfvkUOcBkxjY7flC5Kb31YZKaCN2RAcKkGQoFP3kIiwNkMQaY3smPJG8
y7CSLKgelNk1g/xd0c0aWC6WTkyNiPf3KZAy05U1RKIxUvYxFvKhV1EQk0Wf/buU
MAPrccApuh+toOo8/L1AG2D23hgrDyvrzMSQznJeN++dc9sGoYcEdxXnUFZV803N
o4ZU2H6s+V44TYVbxnKg8mv31nddXQoZaapObEwImUQQfYqvM7lI9wurtak1tCZV
3M5hWj7iHe15hkk8a6fn7ZlkNPnCOzrxDQtrqodfawtvrjIOUJwismeYZEBrdjH9
n9+N5d3pakkVzM/2BKLMIyNE43+69MZzgefCPlmH2kc8k4PpnEpDk06Vc68M9O5M
c8mPkKdxeA/Uk9CeJWwZ1+NJnqwF4f3AmI7AFJxNVK5+A02OUc2KM0Pda6WZrcml
yrjUBt0r+8LwkcFuX1ttXdD81/G5ij+n8t/NTI9drvhAYyrn2gHqJWIgRok0uV31
seHd1esblbzO7nWF2IWRV1CYSLSKjf/pbuQR8UcoBpddIZUoWG/uaaJtTxH82OYb
IGeAANE6WQQrH2sBawZtZSIGXCznmkoJKe9998tXXDSk2D9uhG+OFuqzIMafDWhe
5Tuo7mcuSUn/zubfjC7nl764HfYTX4G5WsDc5emY7TJShaTwcWLzZy4bqdHZX+DI
PGGNkbgBryNTzp3yg+WnFvVgrVYX9tSSahjhCJvkQM97J/jpwg5KcaZND7fmEzQO
hqRPelhsMX7pjMY8NKE1XOrQMTOy+gs1RQ5WftxepzxTH+8GsP+cFQDxi72dFi9Y
rEmn3gYzUl+sVK4mPFXJAajVLOxXQuWma3eshZJfCZ96TGraPGiS8TBWzuGN/uEo
dOPAH+4j049JI1q+//SPeuULPNd5ygxnsEslk4Ndjxlm4WnQHWmUIicdYwG+rDkY
oCrJTuKCfRoVg7fKj2CeEnqkq8lqhv7BARYt6AZ2yZbsB7lm0ce6pgemX8R1uU7L
+UJB0w2NVyn33qYGWCeLDs64KaL9ft/kCupw0qcCBBo0z1fKfIG/LNQBD90syX8D
KPxqOLaO6l17TpirC+K+Hj2+5nj4TlVP4FxSxFjy0j6VqfzVrM4xzm0+StH31VGc
uLuD37x/nLUb4RHeNKLKAPnvWhTorMvWjTS3cGk/fUvnH/MjRkIfViNVyOnsqist
MW+MJzOImgG6Z+XiP9dIx3azfXayrrop3sJSbI6Aq/soKx22o+lV7PAAH12vsJTe
Cu0KHYfOj8SeJPWzM4sxOndVMswKvMrCxK1t9JryzpnkUoEm02WVGMqmMzfOu/kC
q14iuRw8ttpQ9YotcOMUfOhWduX0y2ze5idg9XC6jZOteFZfGtGDRWn6gUQi20OO
6NQa1zzkCPB4XE/6hIjrPrvE/eMlUJ9Kojf5E8fwAsATqC/rFe+LycNtr0x30XaV
5HtEM/TjuYBsb735OYX3bTJ+EmBSuaGtGid/QLHnl0Ou/97uheeIcqCsoLCPXkZs
dPMqecs3he4wpurQxGdCQjOlF57OAIj/kJ88Kc84SDJUmIwZtXnXJp+CXw6PrXHS
DBSTO2WteYuMaZesQXshmHyh/WyyuxV61AMINGa1lvWnJ4FL5rIv9jYYMeUp4MPV
v4jbXhq/eBQlmmieNYG4x1zKXZysxWhsGqnR9Fw5VpoiQhijHTD/AaTsSV2myQC3
eDdpk/HNIoBb/Hb3S/G3iNsKLGsuEdIFZsas8QKGloF6axzhkoiEteGSOfVyU3NP
ir3UXc+OXc1ze3ZSoxATaNvx0Y1Bzjlm2UJkSG8gv+vrRtEgk28UuJ+1Ni2K1TIL
iS4jyg6ADX8QJ5BXXgDnTwXXgmNdO1H1NLR24M3vBQGvxZXwX0zygs+k7pauw3ft
UbimX+MBeqYnphqcqfTc8/YlcM+QQGDq125SUP5DObhz5+L8O0L2Gh2B/gND0tq0
NSwQ0tSoJc/UEZfWCpBbv8oXjxkjYq5j960bESjElZooV0nJLfaxC4igHu2RE3zP
Fi2cc8m+stLtp9Lx7IDidBcErJQMgeFZk1qClcME7sEXC5D5bX8uxzKlXRTctUu5
oSwSKhDz7EQE3KpKd7Vox49YFKf/kk+0ok3x9fgP7PUvoSz63kyZZUrZHasIIXHf
zRggYrzbpId0/PtO4eTc/IsBPU3Y7GlKK5f83IYoW0iT5sNeQu43NqNp+MO+z316
kmH/n2T5oSF7+PH2Eblt0UzzUP4zORnhU6hl4N2R+oIN+neCNCHJB+GarMLkfz+J
hoNwX9uUZFPC2JnwUNb1LU8+0DD1L1TFRtFA1H/dCXoYzKGStfpLC+Um0vDLCkTQ
9DT+ThGarDqcZe7zAfM/CNqu+pdZsjgeQQzitXLoNUknX277OG1AT9pX2jGUajw9
/5D67aLUxLGAjrNcp985kEJ5qACNzBMBJOHVUmgni2+WMgC0JjOx+2pupBk2iciA
lSwRcOZV08Se6iBjE0XJtyHroIKpvyTAVRA2Es1PhIcQzcsuwzx/UIi/ax+xAyvK
rtLOr7SINQrUvpTDl+RBA75at9743+msCsq9PKItqqDbkbCVXobiRZDeWVxVSA4f
eLfhiO0ac9mvF8mDu9RZc0oSauA7YmPDiTYzwyz2q6UYylZ0an3mAQUOD74qttUj
Oi65NbGEJcnHSZ0BtGRkXEas8ne1ZzE8fj+7/CE1Mh2pch+I1+IIguKp0VpPo4EV
LOXcBKuP5y4tPrzTJq+TxSGFgiNzuLtRYIAwksHaX3Lh5uVUv4mnZHe5hETelh4K
WyD4Q3AaiQXs7wxzwxHsud9nTqVwgtEzLOx5E42pE3v+XqCVTx8+jDMPQi266nEp
6bKVWoYNPdLXa7F759Z7JCi+3PYDcIx289NEgUVoFiLyuZAV8rv6nq6JEMN7EJRS
cEzh/kulOl5/6C9YULeiTwkf9JfY4yidEq00G/6slEGWCRnR/3tgm4KLl6Ei4tSz
mGcxBuvE/NOyFYQDTnieiAoV2pceS3DHRdo2opwjN3TufVZm/BUcTGtsuxu45Osy
dJjhZN4iu8LYfoILw7NGqgQuJXb57nqHCbIppWSZVGoh0DN12/67kVUWxNWQN6ln
QP99AWKcqItcM4TyT1ch3S+yB9u3yEqrxWeoFdTh+mUSx4WgyssyPTQ4PYPrcYMn
VYUMCXex+QKrVaijJM8zY8FHlcIirdfEh9eRAPH+X+5rraYzgi3FjbYN7qqP/K+y
bmHrmkYq5WtSLzlLp4hJwW2Ghl+hHRToHFlBobYV1CaobUwYpJibkEgkzBMFNw9i
Y6/VN+okJ380KjqvSFLBHuEOdAeMVSIoOyjMAAIgEXtN13NltwoHKPGixHCGmYMB
z7mq5CyOlSj9eRzIkTi9qr09WsmljueGacj5+1UZS0rGQCnNHnFc10uLPOBdHyAE
GbEWPJLQ0ogQqU3dbY9Jbpef6VE+faq2c7DYgH/EMXvoJ3Z0UXgWrw4g8HQH3s5A
47VteChHT4Z69iO/xm8rd9ZL77WcKjuzCAWA5r5H29MQIFSQ/stRJg9coPk9wAL9
PG03lTZSqgro6VlCQ20CTPkiGzfiqDQh9tMTbbemWK+TIvHHeu7+IWb4/PgfuPNy
UfcUCdmG+4UyNobTw1zbyfGk33Wj7D4rBlQ490rtP8rBwzKUcF1l98TzsRL97k4R
21tNX+9GI/5et40TBblu0FqFRaRgr5aOfEiuQM3fDsMRrQ1MJR7zQe2IsazTkzpd
Mhhx8+rG/StxWOUK3Kis/WRDmB3d1m/WMVegNbnrC3HUghNu4JD0ETO2I8Ao9Guc
auEVmZWeg2b//Gmq+Ha2DtGaiJ9WDrj6gCL0+QEnWs1JlxkqH34pLkhsvpxwDmO5
hPdDOWTmA0I4Z0SLJ6MUlz1fOVn1NblcWEDO0N7DxSOaztG9KBR505dQBzOfEdEa
NiBYfNzwcrbNuWe8LefZvVOjGmz1kEZsj4UTlSmbpwJRnBceFdg3GrHRexsvpHxM
ZNK30dUVRhxCPfA5KV6L4Cw4M1Xe5V9QpCeR7GhUTFRaWonhEOz17BJTWb2FNEfm
4Z4vN3WwRlHu3bs5q7neTq4gvQwAxN7a3xw1E/amCni8GixAztog/T7AZwCDXzPL
y6toq4lO9L8RvQblvsIXO9/3sZHnoS4553O6J5mAzYn8Akk7LR7iKC2x+Nlv/aXZ
VgD1VFMaWMAZMPw5/IzDsx8dOgQKBYHWlrHeuU6367h88x9eSoJEn2cw1y5Qrk5w
uB03J1RXwiesmLXkl36wow/T7whmt9urnCAmH6IKtX+P/PhPrvvzFm5JpH9npo92
vd8G7JDDjh6nrvtr5xQI9CxUaziEyTz/30wWKQMqL4mZv4l/TQmSuffRXR8uydYZ
vNFXGpQfLK2ahVn7QzpZXRCjcCkDHoaHiX21Doxn5+QS6YTu6SBAGNEzDO1EK8S4
4RC11c6Hvu0m8OCcEkBzLk7W+RmEXmeLcRur05SUbhuBHX2xCCs345ZbIGp+azky
PEvCFG7wud5eAeHLUCP/Rjh3/gJrUarItfY8YTXXAwl9oaVAsvoBdj4zgi9hNMYj
xm+gEkzFCzPwi9a9Nh+2RztxO3p2kGkDHNqBvNlLXbxae8EGkJz6SyJsdKSsey/T
kSTsZh4QWYM3ClYxnUYjy8UPMeP3RKhNWS/PDdtjfmwfX7s5Ys+kKKL9aYQgoWnM
qDJlw/yU0qH0sheDbv1dyjGzhmrgQrRBzL/hljlbWCH+bkUCkrvbB/ODVJrHHL9F
ozoFrb3NRt6TuqRC0lZZ7JPn3fUpV7UTf0z6XZC9ae1Go66UBhClwppZCH/3REIW
5ZXOAanEHtiTNF1tGxl7natYtDSQ2wXp7TQHtysv2lcYgZLPQHXprI+7KFIUNTZM
4LHxTeaXevb/OITcKnBoS5afNJQjkuheNLd6XvfjS6nMXqgNOLrFOVODmCukXp5k
QG5SIMpjXeCFxiN/vulvK0dgvhrBNTTt4rdP0HJVVfM04DdoKTFF94ffrfgdDbr8
na5KRhL2DxIeHsiFEN3u5saemTFJkd5OjEIk7dm6h8UM/4nb1Dt0rcvpX6nJm35Y
/mMmy0J0xWNP8EqRQShQzJ6YlgTJxUSO3dCYZikjyFRSj0IQwFZ/LLgg94RkEBX+
vaE3jJiAgU+Ifo3UAVqSS6KFeky0mjEJoCSL2wmkGqlZuLCVTgBhXCBPOptBrwNf
Y82WpUEGDciOrzn2CrB2QodZEVQjP+I/sHIgVFHDnFDkxNs/JxFhBhROdJmlkfAq
4V3XIjRmVJbj8KRnuF3th/t3rjtfhq71ZrdRsqGnwrXZk3bSqt2jE087dCZl58E2
soAGo0CpdXce9kube0iH+Z1GlO0tVIfPL1ayBOSiNhhP/lr9tuOtAUPreBDoJkpg
FJ/ZSIbxiAvxfxttg0d/rPl+afJeAiFUuAa1M2Qt+TlI7Rq5hj5A1Yh3NHu1kMIe
/ITHNVynALgdvxLDHS4IutW3VJng1NR6RV1RJdPWBqK5gdnee0OmbOYNuZ1ALTSZ
sFxLYAx3RnRXhcIoV2sDlsOx5NQlWfRLhIEa59un7uEk4lIB6m3EokeIdkkicS5n
rVKOwInmCaIlEIzjgfFS6H3+uCLJ+IE/xyqcjZv3521OzuNu/YokyQwMPe+CikGU
hSMKyQZ2oTIUkN6vJIeTre/gVj6YqnUMC0cOZZ+OxRAL9s38JKCs2jar/JUMDJco
ajkFScVwItIw5uaoA87bPfWDwc15atrQmjZqkyQ4hoXeqjUehNm8550F0obA91LG
ci7keng2r9sv5F1ekaKc7yY4McP0wVPbVvlN4xLA9+PU+ie4Jw/k0HU3CeBJTKth
kL5mDQz0tNiIh4HMIV96A0ycnPt3/8Y7OSXaJWKbEJy9Ap3gjur94JY19oRxVW2B
wSxdSz3/yMklYt/kyXTLxCP9fYy0ehukiF7+8UznN7xUfGSv74bxXBQNSfjmTxgi
+QNrzavE6zye9ZEd0m0IT1wmADz/e4X6OSkhGVCHGReTdPc3NSw7uVm30d85JQpY
DDPSYg2dfW9hQzwaQRH/lQuC9nC5D+e9cp6FsVSSnX24dzTpfnO629FT+gWs9iuk
qT8bDE4Vf0VKZx1mgcdY02iLMB2BtMg5T89lq+xRLH9rETh1x+zOSfh6IG77W7rr
s2pzpi3/RrhhzeWYcbYD3IBH8e67SLnVClfKPdOC/zGWuxVGKqP09OPS1emErbxI
Q4aP+h3dnT8hBxKPsMS4L9lFT0zGTgoW/PCWHGZOsT6n9QBlEDgfJAIlwCOvwebh
B7Ryo994MIbU9fWetyHAqWv72woc73tCpJrBqt+MmLKNQWCnVTXrUDS4553whqx9
ZiRoOahVVt6Mqm2V5rJsEB92GACKol8OcdVvC+K2xmLmfFgivrtr7PMK1hUt5Qtc
r9gVNeG8wfov/DnjPsQL2NCADkbI6VXxfcRcXdvYVMaXG/H8Zy8w6qxu8Pdk59ea
yS5huRsInadWLf1ZtrO8OULr5+yShv3fZWFZmOpyXuBzkUHQzdLMLcE5Rs6zCNSm
+AuTE6LwCg+QSxT1vhBG+/MCUYZAbVNt0siVy4f4yQuLLIdMA5Fdq07Awr/zh6Xt
k+S1HDns7wyS9Bs27OeQu70n7TrUFV0qW49bTbavp0SCVmlLpxVYlOMQrQ5bOZiF
sYhXTwRAcy5iutZU474wwlgzHylUOnTS9EiNMWk1lOFfwiQa/bUQUvtgTcFBkadH
zLiinopaj7sCpIX+qQvPGxhkUJzuLyW/AN3JdmK50TN1uwk5JFSScG2phMuqa3vk
PyhDVVXenrM/hiZuZQTjzyFHVR8bmqAYHmE7bL/M6doxPopgQ0nxF/ujftKA9Vc6
slwt44b47+uWYdN5Akqr5SKEBcnrsZc0xiVPY4JO6qoeDfxxwMqJy59JjYmap5y0
gz5tdDAgH6xX4IjlfOQDj32BWhy5t+h3ZlRa5Go9FEI1JzMkN9HY6p83xZnQtJE4
CZ0ek6ZOWnLzG/zNTLtRoAGM9GdW6XHDltsB7OrPjydHTpISxb8GSl/RKd+0bzz+
lNr3QvWeDDBdmI26dCioW7uGnTHCouz1mWNQuCbNUAp/e7B7vijOJvHt4Rztxcgg
9LyqHLI15GpNtfEGsS+GUVaZZpCl1baXOvHUXsssHqmdAOH5nnbA38AH7+azaxlR
2uSO6Oj1W7V5B6f85rev1XoIq1GZ1TDzuTOQ1Qw2vdX4XQwjcI1mPAO8Yh5QrQbw
8PuOG3wvtIxz9mstk1lQRo8SCepkJEhMlHniuAZpzEhMqgUS8L1h4qtr2Onp6xS1
BjzSOdTXY2R8q7nbAapLb7YOhQKWr1BmcTUKwZ6HvwkrbJ8l/htcFliPbfc3B3hg
rsvc97Nv7ZYtQDfEoc41EuPdtXAauPDMMPzTL9q+G1+R/mdZCCfYgr8Ws23tc0Ao
jWh0X9zmdz7jdMhMwVKSAtawXkD3hi2rVioWTh+pKRzraPNmpBTUwAnM8eEeuFYN
cMyxqy1HGIkzr/n/fpWcWwRM3E+ZFxJZ2/Pmkuvsq1gOekQA4CM5blVKXYP6URU7
mjLhByZXmUSafguene5wjPgGffMbX0nK65Sags/6RMeaAxrof10fMcTUav1CNP8N
3gOHW5j4PYEBx294J5kjAVqXIxDmIOt/NiOhpeLaVDsxpITPZ2syfrUzojpDSAXT
DIncgzmFoz3hT4e4gFIA7B91Vu606nMMuo7JmxGQwEKRFopPOWoEswmWzU5agwmH
ukAgLYSKBwBkfihIm01ZXEtxfYhdO8UaCldJNkzrFw3ND1icSN8vmRqDQx9BNqm5
FOcG2Hqb+o9DbnF5p5YCuQNFntBei17bFL4UjNPGf1aUeoXqciAk4mk9JWA17NqS
MBSLypm3z263VvQ70tjTFOEuVlla94EQCw0XaCZ1kzsVoH5Btc8gMOmAiq9Jclm/
rFCcrlZh2Hy7ESxm/6Z0RLHXOYBK5m/gOZo9bIX3e6606jwJGVbyAXzk0y6++4eu
09u0ZTme52wcjtWMg/LtqnXznMpMkP+1Zpef4U+dS5qYPZDtvc36UOd08fw8GYp8
6JeYbS8b/+c2JL7iI0f9hIyMNPMu5DrPiQ3PQslSjFwjyf4787HW+5RYVGMFV6fl
/bgd2c3FomYQtXVtmzMNdBLOLgLlTAr8mOIiN9E9PBmc9RkOEuRS53onG7zYdVQh
h6enu7+PJOscVtvmzHGIjdWk4rgD+oOQFZceMvR5Gy3opPbzXLZfTcje426DYiyO
JLC/ri+QbVrgefd57jjGrHx7yQtHEnW4fBwHu4u909o2XfKzd3fS3wM8FjLNURmk
cu1a9ULcwQRsaba5CI4DW6C3AS1wdmUzToIhv4iB1u8ofdDDAUHgEp7VjDfvrMK6
BS8eV20FiAGjXS0SQ6N3TPJFUtsztWgaj8m9UpaiSbg/IwJMBLauuI22j/KwtTKq
evMjz2mmBR++jdFZPV57nR94LgIn3CwkJ7EsRYLcFV9EmG+SJJSNlfqcHgocxm8z
/HBsbznA8kuloaYnXUxgqwjvNUS2Ad9sjDC3zuwILKrXh9hX2a4ErMp0xu0df7uZ
Jvp93ubFzs6dCOj4WZp8mUuVkQc8yZKIbK3pTXTPXA51+eL6M1O+uJ1extj3tbib
Bi5dUdMX1qsWnnFJb4jelMFq4yj6kqRONXjxsOFm0YI4gPXiTdKkqFdIdCirh1VP
HzH+KEIl6JgjLU+UMScYYf8pG4xMy1Pl1OfLqOiFiKrKZZtei1lENMJKjTn4P+6z
KZNB3+hk+PEOdCovIpmbmt4tmTnRngLVKlAhrtbkQMwFmHRqhv4JKWFPrXo7R/LM
yrUJQj00m+FMVuxc5erwqn/fi8GaXV42MNy9s7+ERSLYGPMOV5YGJr+F39dP62D4
VAyT2dDn9rWkTQBFjYXjjEaIgbwjQ0s4WgeznKVG1/pOkM/Wmv+RhNnqFKHv9gLA
JluGHJaUARr6v1bktP1Qz35Z9VX7QdbDSXT4Annddn9kqqQYpdG5iu56bdGaBYQq
OTRTV3Y3a7/3GWGKdnBRf63kV3CMKGw3T7JeWrWM4KOk75lXk37aC2VUVhaajr8/
O4HCBxkXDvXJXkD/6ngBPe6J4NO3V8Ijqz0rkfStocDZ7ehXIEt/zq4pxjMr/JCg
CgbIi0DOsR2yv/A1dqBXW+8D8tBJsGUr/5v1LGGTVDBRxO+abKw6ardreda3N7Is
+5zPaWp7JNeOSbDNAzSsHqaliv1yjWbMQ2oUrTXtvPEDKICrCT+b3EmUjthf0R/v
gIznU1zTshRtqRDHhX05oVIfwoKn5vbKsfKy2ElBHPFMTCqAFlWCev9p0lECvDSw
eNb0m72EPkfp51ChE5/Ei+N76tyiQTxO+DB9N3uW1dd0FwSTf3pduYfBooXf7ukC
21uPfQEgrI6in1nloYb3wQjxci0RFew2mWlkamhPsKzsYOAk1Bkm8BYI/m6So52O
dzDEQ36p0Y177c0lgz+q35U6LA8qfak4IwDyIgQKgvv9cg38dr6Bv/GikU6VNbPR
+sZOBj5fL674lDzUueVRgYnLEtzkjNugDetaYtlkGOPuOnhce1c3I+owpqGvnRun
h+GXjwElxWsXdKzl0LrxvCKNeYJn3kBziGUGZaJ7D9wQEbEPGdBm7TmHwzO0l4AB
OxNMliYpw6enps2BUROGsLZM2LBlREDtintZWyUwVfrqpz1HteFTIJ2Vwl9r1Fh6
2aHAkWKIEzjGei224ZTv7Ey2luvemYYqPp5nwQNh5EaGGCwxDF8Soz93IgbY98Hn
ZmgYN7Lu3jsHCHVHveDRCc5gvb5C8yWepTpgAhyNyHgr5Adwy5ohLuIPvND1lFV/
O0awxPG+LAsu4V/pNQ728+WoJoyCDZvfVK54i15+WBFduXACDLNNb4iH5EoXtbVj
eWQarBf85CMoaCn7rMRgupEBwn+lm6SqF5ekW1YTMJY+rQjg0HhuvOs3XUAC2flT
0vCayu4svnkea7yF0GAlq7T19geKUQgzjGMATcGdMXowVJLrfY1tF574jRILN9JP
ABkh2i8OGGs1uJC3wicQmmr4m6GEy/2yfLTZS7sXs50lCblAjjzv74fNT+Yd8KNo
MBx2I23rzyLl0bSRv71gSVlMrUoxjxQKzQj1ifReZhkoE3ouOsY8x8eh87AZ+6Dq
Fn/Y6huTk9LWCDpJMAEKrGIiuiflCQSrAXrClq0hvAcGaoUSuibi/YvNtmDFWGEE
Yzqx50HkMPL8wLFUzy3EcY6EdyecOEjudaqQpHUtGHJsqiBzun4KfgvFzi9yLhxA
UISoVlcj3psBRwT6ygECsW03F0dtPREPGjOq8UiDgaVZwA69JXA/tLiwE0TAnbsQ
iapZgICkcuA3WTWAAA/t8eB5Ei3sRmmUyQEllTGcg1mWLtVzdjP8IFAXBg2/oQcZ
aG0RxnfOIM+kv+wAuRKxuXlggmyYJ8ZFgVArJUIulAUEOWI661g+ovsUSp3qlSE4
KmLBZielZ3OrDZbOu9hIVyn+0LqEoyrvAJENFy5j6iFeoidf9qf1ldF1pbWrSCYB
W1oqGXQjl5f7ks1pyR0SvV2UJtG3kVsQOk+sVTxaWiBJ8ONO8dLBusSib0LHy5Nq
b6Wn653FN1BecWDmLyx7qDqczg7bf79cIamEsyVtpVcpeZXE+pv+F9Lw5uYPmjWq
oarCo2/DcLBDjDzvQj4zEKKUtLGnd+uEVbftz+eyslWyy0dFnY48qGhhBLZRikUG
/2hCvzXZ6AfWhYhmUeeGsF4H5J6LD3ucg+4wgCFJqf+6K302LhkQJM+X1I3mdvvY
MaqJ81iw0XeCX6rTFwtpTPymag47NrFQczptz2h337WVGDgtq8JN3C3ESJiGG/3w
M0+H5P6SQh0bnybx9QQbjvsz8W3fpz6Nf8TwDxLgNe/bNNARhEvD0eQSjfSxcySH
nFuTZ137ylyU/XfvU+Y2Jzf/WbxGM6xNz+aC669r3odYbGDxsSDlJ/S/fr7IwJdg
MoxHVZ8UEzKRau+uuWvgnNoVpgvfY2uiol/r5haimjTkeY7rvNvCbSxiBT6eeo5C
4Lg/cTSOTCneBt8HgiVC8PDh9PtzVUxP6ljDfBS36jr1AXGdBneeumFylWVIVCT0
XIGWRBT1yOQJe2c19UBm6cqaY12aJF1Mp0Hw7BxcL0qFpUbjxaP6KPqtmB+V9UX+
O4zoRjdUH6H1Wvz5H8FxX4TpvYmjjTh4pknyaT0Vs9FGxUex7yPYefOF+pl1gqLr
vD2rfla24fFcD6bLp0buYTt2RAnj9OcKivGI2HHU56wa8GQ58MB4lQoLD2yTNR4a
MMZXjllFMcuj6BiI1jyZLTg4RraWZKIB9JE4FZoxN1oOR9+NkVses1fyOcIC78dV
9jHtS2pKl5rg1k1VP2UZAl2L1xzHBUW4cgOk/KcXHYMzlENVIZckfPwYUEWjDjyJ
BHMKs8EX/JvX5dn3QiuJK+a9XPRIaOfTGWv1jNIjnYlr6wGxVyh6ZGVzTQ6YucM0
yUSTmi5vW0YQKiQShbK3OdPoMbR6DSYoKRfjFQ9+Qui4jMFXud6mBVe6riWJVS1O
yn/WxVc0Vr5flMOzxntwPVPHE8cEUgkeWjl+IWzB0JMNnhr4OdbMKDboJCbULvWB
d+bEeTGejs32lHmsUpYtuKor9ZLdarZ3p4fV2xzKIksqKXa25y2GrivWrRWMEu1D
pLDEUlYakPcO0ot2BJppyN1N+1YX/Th8RN6NeI25hsU42m/VS2Y5q8kLZTmw4Os8
AXFp/0UEYxyM7Sspd0zpzhhp89Dm++JZLzzcVpm75cg5ezdd8Ubo/IPDYelpLKLG
n+PMAlaT2DfClVpm2yz/didCE7NKPBD+q5KR27sD7BImoRFYsZ95qA6fqgEd1Roz
BMP7Db64YfgeuQ3kJ6MkbjLuyI7NDGCuZvtVL34M2iyyQkdHGYCr7NzmNtsAZdkD
9b3Eof2slSpYAvcPM88ocwIeLE1jgqEWh7MhMsaw0yhSfSAZjpW4agdHfYuxFPAY
wDFkyMDFXLmn+xQkAZmU7HBUu76Jb6+GcGH3XbfKR3dhA0DL7P8uC7glDnWWTgHa
7Px4eUjZtxfpXwvIEf+vfVQD4zjczpzVnW+DxNJoSybgyPAf0MhHJPNvY89uSvSy
F6KoupAhiug2ndXpYwRwDBOjn6Xa5mvzXZPBhnmGAZcSZR68bzrQRODYXAjB0RMe
tpNV18vWzTiHa4P5cMICI/K7OuMPXpqhbu0fTTEEhnehhpyVX26WAMIQgP2/sPa/
CzYi06MIKT3lbyt9qy/PkhlpDhBJoE7Pg6eaX/RiNCMmC7ujjIPqVfDmtxrZ1B/w
z0xCsOku9uGBkVRcTg97qSoRD6RmDmuimv/1knMnfyVOoesS4RDwtMsuRkueBeUM
uuyAkpvafCALj9g/Ik+wMZumVpc8qhssrjTmUgDAqOMzmJzBQtkQebD9M/bQL1qU
zXbxfRcqJ7K2FFR0aiqRZOiP89KVBmt8fLwVG12CFTguomro8BAkqdYskj17sABN
Ulm+uBXuwJb8f0RCpv7SJNBlCizxKcKOrtC97bFsj8xKegreYcnSeZT13u7v8bWp
nyrrFEuG5GMFR0/6dm+guMVIZJz3f0dg7ER0PnLqHZwyzMTgZYeLvdQV4ZrAlEYc
6TAwtYhzkT5i+8GNaut0bBmGKP2FLZR4BCmNbH+KaAvIDEXfPmzzq9E4GFaIRzY+
NUpSqXQPUxxB+a5rsM+HJgWaL7Ogm9Pp9Gi0tch0CMh9cfxDR69TSTusOsXZi6gi
HJAxne5HpS1dRvGnzlIjcp7ejzc2IAl+wr4woZ8xQgY2juUFeSE6Pl/8gKZDexB4
PA2PRlGIImEyc3M0HiALUy4OeIXa+LUewQQlGXZqlJ/m5E7f0lnrRUsk0tTJ+YUN
3907Yj0dl7yId5FgJo9cg5ho0I/j3iw00XMbFKnWvUvAhKEGxOMZFqzNHX27fZxQ
i0w+3bHpogDhCc+K8LDUJOEYcJOYv9IlndFpZR9vpKXuRkQ1qjIrHOXHqSmk2kS1
4IGy0VYa76SAFWPxHWUKqLHJ+iWVgU6zQLlu/p0mOpUTaz+eWOhmyc02OUseen9B
YnKKi04uaLbcpfKOlPyuZ156uku4aqMtVj3fYfOvIbzFD/Iqirrwe/XmfCcU/Lte
X3bcwHbh5Xiqr23inGf/WYhpoHAU2WOlWoPXFThjuu1dF3cwRmnQSAfs+uyI63WT
Uhv6djWQgtXmqyoAwYZ8oUYfCO0V91PkeMjtrxbqIb+zx8vORcnXIRau0XSb/IN6
BcKwUS/sCs9wwaao/JH7SSwJ9u8oNZheeWcnl4P0REU6DYYIyWn7nlXg87jg2YcE
MPIDkV5N5HELi3XIR5skTGz5anWLTxAzKq1du4YdwKQTEm4yiM+Jyhzd9BhSvkOS
Pio/UmqQcrqQyeFwvzpIrFYdyA+FWY0ecTYzurGq6O/iXiWdgaVfYG+vXkdbe7OO
JdCGmdq8/onB23rN6oNXF4GvfwzJIFN/Y/egRujwNp1TduRCsgNjW/NUp//zXDrI
HZoJ3NsgxJ0khq3f8Cace8NGKQwbES1g4922BJj0kuPWVszL+dREMad9KU4PAXyy
EGKC9JOZiRchSTuPguviY1grPN/ZhwINLVJxXpqybkW6jdjVYKFHxngKZNDmXifX
bbDOgckV53VCQq21BxsDWBIbGHm5NxbxgjvYzMVuYhxFykFkYCf1vA6C5V9AFeCx
vHkstRXVYxe9rP6Kcg/aI+Qg2YAy10pi5frpV/d3oqG7VOauR0RRaXq3i34x3O2z
NGcYU1nbDeVUzFX0+YmRdzDnF6aieJBnEZkjaWNcSqlT/2O4MG5D09J6+ZFJa71k
0FqDLzoaxCIAkcST7i17FwO9KWf6HNqvctV4vQr377pFHsc4eKdFJoYbGsGHOVEX
xqo8g0Yb/pOyjUB7qTDxxt/TumrLqEL8zsn2lmAB3xQl/0nSDf/ULFPKPsnJdTXJ
kfYvK3hYSYvLnlxkHxZ4HEEaxvGXvNwnWqfMxuhEO3vRqRa/LYaOTBDunxQd2Sf7
3BlcWGDp9baiad/q6Wwz2bx2iVORIia4pTVQ5Zc5orI63fsH/+puzVldsSTT+avA
pdiUKJdzW4gqgy4eFZXzAFbFXAAyxuZAuRoY8sEtG4IqOs6TMUQ//3vn+FpP8EDe
qUbKLfxXJfOrGuEV3xUWO5XHhbvQXE5T91xfFeIpM6wLzSV8zBvS3uBork7Rumv/
vNBftdvvDIuZuIfhgyJocLHMMmp5o+K5jq4rEuUn0/l2ym2zMCw34ppKVxnSuXk/
rEFEm+SbKhg+jgmEBMj7YMZ2EDl5LEXMA5Bol/6EcRfbTVncvzNZPLvYA4wOTPBZ
CqVnpbbc7VvUXIyr/ghV8cpfea/tdqWXTZY4PqoMtoHA/eR15H9sRwOJnbREZNic
AkUbeOHIoSQCgJad68Agf6u9amKVd9fM4/Ezg6PY1R8ysthxFvgxnAmn4VlpMsTz
E6x4gSl6aTiAY1iubWxaCGrY4bH5kH6jxSK9VcshKGUq7ehA3lkeecz+fK5PyHOc
b9QnDrOfBLJbpEdoNfQ9ctgdpGJd1/5nlvpEOMofF3kB3SDRRm080cehf8csONok
xG8TiHTBkEjV4+e3djitmQD2R4z3ExjbMnfFK6uYXK7HHfCOzq8VHSixm+0StoAj
kRb0YDBU7F5hJSvOAieIcAUXmq4AShPtxJk/Ppr20/Xm2YHxJSbFf7X391ZB1LKZ
AwoGVk7i/APoWrdzEXjf+Vgx5skmwVjLcWDokD1WW6UrNry5rYZfvcKYRq2n2mYB
2vBYFLlEqCxSKKrsrsqFC74d+hRJOa0iC3gyOv/V8qzqxBxZ7RpcQIEaHrN4pnIi
QG2Q5QnARmkWgv6HTCy79N1BdQseo1yHjSftK/in4kAoTONjh1cIx/mU6A9JQaz6
IAFMqpmPg2FujghI/ISPjJ86uxr0x+Ci66a/wATb3TUgrcGiOyBSmxs/9AnwPJhZ
S9lMrCVLrfQeVJcTGz05wK40xwErq1XtPtt8s1YR9VKcXrYXdQ1So7h43UxJbSDk
qGK3b5kBSskkZcvb9nnfx9L4rkGDXxX7dltixEJvGcrb8Euru+aa3mNtLCQFzDyF
/MsXppGkVg3v6KFLKhknNulmSSHjhGQLAu28ZEnMUdEt9KO14w9ylJD2ASMhCI9H
9bgxvzY9V7Wir7gfer62lrwxeXyk3Gu3RPttkLOAAobci/oR0oHZxapMu131f63L
fi8SpnbMuocD8YzvsTAB45//wsMszPDY8XV6aeuUg8sUS9Ooyu76kW8hUdVI6XKM
6XMVD5RfMBfdniodVfvO4kFOCGQkFHyYOuLVll+lGUV1qnb1NWiMXdp+DmaGVuJi
1M11PPAzfV0lfq8TzgNQzWD1hMSryapPP2JPtmW8yGQEFO3XP//vS+IsMZojz4/T
nY2IbcYTNI2f+a6E5r2oCLJTdblWNh6n9tiCxZRW1A2XqdIhnDbYZvParlr0rr4D
SMNNjWVSmHD7jHeYl75K6wvb+T0++tFllPv0ljt4KALKn7LhXitpeX84EDDysnC1
cnUJoyF4hQkFCRWPBLBEISc+tkDeklF4YEjiTBcz5rHNFl4cWskwbm6/h4kE/Hjx
J08pH2MnT4elqsqrh7sTqUq2IMr3eR58mS5peCIqhBm5t0YgGH1cs7cY4vftp7lp
SzZ2CTkuISc/B3xDgwlPzk/yAPh5H8vi/vmTRreduTk7so10cm3gl719eqfbyKxV
LPbGz8yMtApqHUZj2qJjYniD/XgdNEVQvPUJgm6eJ0KdVW42OtWO8rFxkO6YDDHJ
cKh4Q7Fxpskqul9vvtT58MlN7b4oQbXZN0XhbSdPSI0rMtBlLyJpci62xPFv9Xsq
EI7X+jZOGc7OVhskBE6dUk31SVDxukKxMTV0XsUC4Rg2QogNB9ogh+zQbcZLiRRa
9ygrAxOqMD8JAQtTFOtbkEU/z8ahH6V1mJG4xUNmWK0L9lx89sR3f9nb0qGckpqf
NzKcd7D73+UxWFLB4kiZwo8OwBYE4gJC/TIhXC/3CID2JutrPMN/1ecurGcLMpm/
grWqjOPIEGgt2XDOn9MX5D5PIZzcepYmiyf0Oi8mmSiBLVtrIqPiP31t0T6jP1C5
NkBEC5AZNzvSuSV9AXdxsjJ+9RHMzp1p+CUuR50HJDH6E7ZEo1GLpJMdIYbTZOZ7
fUdZzuVc1lifURnBukfxiQSt1pA4f4Kme35nwHUZ9jzhkZNLr0TmeSY3Ik7N4Vbd
ShHLOBHLPkS2HoOzcc+BRuAqgroUIteZUqO/ou3Z04NGGQpNu8942+1ieCTqHA8R
JdLtC/vJHKE7dWwiuCtOarsC9NQ1EWLDrh1UnWN1AqlW86GhDUkQtJetfqpEOlXg
HcQq+GWMRUqzf6Er84N4Q3lE4qB1L+4sdEsKlZNv+csiQzkt/tXKuA2gEcTmyAEb
3COFVqJ5xnWT1fR0iiUpEGVUvQ9GcowYFa1k29h6gC1xW8NOkfHCbvSZYNvHKolS
gAuYquhSxbwkgs9I23DMAieuYYrgSzp+tKwdmFWo/NW97j60GGZK27+iThgvveEK
jK7IYALtm12izXBHQWpP6Sn/Z7WRlbxxekD88nLXUKEfFhNDXewNlMZOjF50SSly
Yoq61kjouAQmG2/zlbCtJwYJ0HGh2Xjrv6ZyFdwqc3wTCBd6bcxdqjn2Gu6fI+2u
hu+NyjiL6Lb6exedcerZ3bTY3JAcJUgl3h/4p2kpVcHfYoLRtOh4GVGZqB8sFARv
8VyzBO0e+opgFwA6tm9PsiuU1fTTHcoCw5SJNwTh4bfgm+g928h1tpsduFOs+szU
fQIZyKsj8rVhmmy2PXVGc37Zi6VdthtvosuvaTzOtKQWAOy05U5u8sJXZ2eL6zR5
WBxsi9PN9/9vaJefyv5WOvd7Pi0/VCmKcUYVIHWgx7yutG1v6aZyCQ6QSRPrMxmm
UcRNtrdckFxRSkVV35oaxjcNWYK92xF01RpiZ5vYMdhmJnlVdjl6BVgCJZmO8U0L
dvBSFElGwRf1tzl+jragXUkaCJBsu2YHgj41yw+UDCa3i/wXpwNXEby6zFxxL0Lq
e4pyrMCT4tVEAoLpmQHLiVywOgyUqggQUksUVf2OgXELapMtjt9uqgDIl4l0g4D2
VCtivRU+k9r0sYs2AfMaP0LdAp3wCZBY7gez0/SubJHImhOp3nPodLxFK7Z8mF3J
7Cwvfr9agicXtrttAeOoao0tUNzq+WbiVXkeRXrOK7xjlHJRmkvUoMAgktyg8fBr
oMXBKDfS0vyLWCfA+Zf0sS8jEDNgIiruf8bPjaw/oZf8xkSBZcLXDsSRMqejCAk4
KfonkWQWo5Mu6MUgo7jwSUbzy3jkkByKpxHVKtTikRugDRTRggT4uN80nBl8m0WF
CEpKMpqnRWtblpB53FS+iEDieVRoIaFzg22/q2uD7eLkmZg09HyMS9UyhWoHK8Gf
sG/wQ5awjy/gBbPPxkGqnr/fo4dkNaphE9NCoInxve0WOEN7qj7j2t72iFrZD3Wb
/s/P/PNXir8w/KHyRqe2G80+/KD3jlq98zavW57fSvYrFmupKVQ2XuOWtyTGLf+J
d7Ez9iYsQc9406E6DeK//ZJutu+sxs6rikNaLLU+5t3lKn8NlepEQg/wLCnhAVfy
SocTBGgksU16N2/lvlyi4szNIV4NKCOMM88pqm6I4A1bi/nnMgFh68Lb9jTxdVeG
Gi99jU5DzWZbT6Zws17c9lzjlVzX1ioECkQ5dIPmVOFFk/K07ETyWn+kG76wQVGU
gF6GZHVT3QW+UlU9h5x4wnSrcAvORAlBQq+7sabJIxIvKl+g3xQOHOT8IacNt/Ep
oyb9gqq7zvusSEQHiRWiCi6/jq/ufDHOhrfxW5Wa43Ldmi7gWh3BsPapv8UDpFEM
AGsbHeGx/CJ2UXDV+FER/KbK/VoPwJ23NzL3RJ1g9cn0XKMNYNqC2dpNhwpxd7Yv
K/3O9U8hXqE0Pt3Sp0YxV6rpyhDqaz4Z03flGD5TV40Vtv+rW2tLGQ64XfuXwWzN
eId03q1na72FQbhZotsQCwyTWtiTOkEREv/alHjQWTce8FPUGo/pPenDzkqhUp/B
NBxMeybkGR6bhyImddP6FMyIDbatH+LH1T+kRELPaA/21TMyPyDouPy6QbRv9LYe
ezE/j/82WQh9ADaLqfTDx4uCDfCQ2QDkhEoWzNbAlc+Nn0VDTuWPa92IZqBCnYsD
1HP0E1kogCN6Xyqiso51Z9J8FFf+w8M2JFkjqO5sa+xw9XViRDjbTZV1ImV9Fh1w
kY/JcNDrmJeZx+RFjrDZCydeLZTBzCBqqOMdt5MY7Ur9/3F2uTC7k6lKXllhvk7p
NG34RSyjCZC3hvi7k8/Mp0Z4RXcOVmi5Vqhd7BE11PBtyQRv5tqepF8yfIpXDR8I
/8uRKit0R9D3OP+Frdkxa9U+5J5uQAfyuGGG32w68i2Kz0JOpr87wUGG74VnFgBh
gTsdxbJzZZOMdTHG7qfR938HhUQxMjuZEIDUMRURinedd9OXFOJ1o1bHkUrWs5az
Qq7e7t/A1wLOvwpaVQP5/3OQS6YtZeEUNlXs28wXmatUjqF9LzZoJMdKWRpkYh5F
bXdoM/ZWl0fK8lwM+rbUsGFpboS6COaHBxGALQt3mTWl8SOi0+rLe4DiQKM+oERD
78oF+xoP30aMD9D8mHK2qdplMxxqC+rPAspu4rUY1efXVkm0fFDGKnbJhfzsa6qM
/GgVb8aLcdkqtqytOj5pyaESBYxOfj/9pY3UoQ+RhHKWsc98Dv6iMloW8QYEe25+
cQg+tqglMFRZT7qnTo8oMub4Q0u9hGc+P+UaQdGH+EsWXdmC+cihSRNn3CC5IDGZ
pjlrTnyTMT+GbaUqCP/QwWPxHz6cG+zB3/MU8xadOIbpr17zGEfDloTs0YSxUbuR
E6TI7rkK+rEitAEc5g6PwWxnYyGveWyMaFvNmp3x+k2Uop1IMQU4AkoBqXJawgG4
croi5GVG9iJPcbO/YodFxy0EveVmRhequ2rtZC+lD5SVBadmaDEf3knT/wzYQX3g
8lGbffeSfqE4odFrRmmf+3idb0MQbtV1pdrJUMSOtkoJBRDdBT/qgc/21hwBs0Lg
6FKSI6ZQCGtLRUnEFROQtdN6utRq+7cazAGtZ7+csAwZC3iefadyY2oGtpN/+O8u
Q9lFjCPpGI3iWJw60EXYNhJtqJD5Vc1BAXFnalOURszKZA+MnUC3/lWordg+pACU
MwDEtxcFJR05LfoaxAdZ2WwAReIdhI0G7EMxkVzcgOJfChDAVPB30OrbVjgq+zox
GpGoNbP1e7caoOuKqMAupAgx+wcuZBCVme6tPhclqscDzrS+pnrFJ/7r285rig7v
FAmcK/Kl/VuusMTYeDbq2aF80oS/oNGuLKPm/CwbzMro5CTa66/i9GReOnLAg3hs
Je7hj+Z/oPDEI/0fQDU45M8oVRNELMBCgDJgV9HfbgUgjnB6UL1DVzVJrEd5ECHJ
SnjAJdG6Cwt5t/6axpgGSTJuQUnfzizX3qOeMEq3VOrneDkG+VJAAIZbe0VDoY7R
NfYSy9caibniU6lDJ5mhKgGAK93VyvCgjPg3HCzZWvBNrumZfgmpkvftL4U+qft0
7za3LCznc4N3gFOHm5toKJ57gj9jCxXiG/3ZldSDbWPXNau+AS2FThXUqNgsXUW5
UnrxXFclyqfHUHc8aAwsW/WxYb9R/o3pVAPDh0tF+V68O+Ng6vSmXUR10UpdfLyQ
Eik6b63B/ctzuJAp4jhN12YiVfznp5iSuU4kMpp7QwD2UqHPEZWVlYwsgeLwKnWO
ySCkQlADe39b0I6Ke37o9WGtxTrFGo8JOFDtr6TXn/5s+Yf1GB1P64k3zgyszAOA
BFaFMOwrNa+nKaEyrc+cHT3By3jwvCr4YVA9/GWIX6sDQu6eefY9o3ujgwa4/g7Y
NfyDaVsDnKFXO7nyRcdCbmjABpwzZYXcys1i20Nc9FKS0p3OZbbzppqTh+3P6kg3
Hs+4d69AmW+/AEU5D2DJSKVtHqg++jBJ/YkinhHnBj/pvyEnDZ4+aTP9K9bQd/rQ
ZanKcISHX9n4L6SPpZaomiT2A3qwmfvTGJ1OVXRnG5yClrAe6EuQRtQiFfKuZ6iN
c0/wXaOf4v8LKoOPkXGYA3H8XkStV2f+49owJuTwvZRdhl8afX1iJ4OTL1eyuPTY
ghfmuF4ezFSiHeg+czSob7kn5LfipQgSbNd4W9estwAGRkVX0MBOGufw1OM1wk/D
sD/NBMyy2QJeMKOLD//03V4rAGLXENCtCzyPeciPsE6HX2MZn5T3FuYj76+hemd3
jGm+IQ5/I1u+GEV7+hSOp4X1b9v76yO+YRraOf44HTQgiD91zpchPolJyqYszCKT
cLifNgEKHYkVPVG1rj2ovkzsdxo9KzpYGqwjflDl1E6/c0SeXci1LJKH+OuZz3YK
Oxb3VndKFzWybEPLFbOMZtNAPzc7lzoOrN+QcrwHmA3WCGvVPUhl0akvsLsv7nWF
C7nIQ1GM58BNykq2ZwkN5xVkSoJP88YuUqX/zzMR5iENPDP2JjI6SiIYOK++0FBp
gDkLTJnUOy852YLkFcuGOd0+oXaRwUkcaxYYUDfj06assbpU4eUvoMJazz4F6YUS
GtQwqtYy7sAivxUgd+d5/RL1//hbxIykQUtfGwnY1UVkcKVSiS4aE3ek6Cg22ZEL
+53o4jbHVuWQpWsetf8pw4AM1r9gClulTZBVnVzwK7aTx1YTUMyPonF7qdvs3FzN
`pragma protect end_protected
