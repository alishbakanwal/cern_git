// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:34 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
A2FwuoswACdWUU54rMLMW8Q26ARrhiMBXhBWDFIU6VZRnf3zoDc30jZ8y3IXoDme
BJDvQ5kadet4Jm08PzRuW9Hp7PvxD+z//3S27bVq88plVpzuqch3CGsbPF0Yg0Xf
ng49isr+DSIApKfGUwmvSN1WLVkg0/B63emojo00yYo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6544)
b/obdgr9yBSuLkaJQDvgV+DB+hU8RfFUo++BvI3i9kXLs+nzmUYQuW7B1USAclWP
U+poTA3hAVFHvquNBCp+yLS8PvDZzvjfLxzAG/hZ07fkGRHAM5U567uMb8WYNsud
kpynK7K8yf0JGvbh0fkyjStQbpAB4n8DSOPxFslvbKD9rbcUN70NW8LGkDXvNBW9
sTJDU0wR1A1nKtJEB+aF3+6xnpUiIc+znH5z+1bvPtVzTNFuMYy83NXF2/45nQww
/bGEhd0UKfz8Wpyz+oOuaelRi16PTf8luooHQe5zLOLSRdgJLnTxTI7m3edygrJO
KJFurNb2zj3jWYlWWHn7OWLvHWOrtfksov5blzLESUVTkTbObkSMZtbh/i7vJUIH
RfpijhxCyz/XAcImpkx1CcsafGs4bk2pYol3P0AjaEvpccvMIiwpmxlEej2nMYHj
JHfsq9FF2w1U4gt7Exk5wpWs2e6VZH1yQUAMII1fUUyKA40yZQFEMXzIYEhPcaax
LlieyWG79Ftl803x1scD4gwA+lY8QiFoXiK2fGjV3TWeqnr+NZ1WIWqA4vN5cl2D
RiGula5imMZQCGzoStyZHWoxBO+yP4DITrioNsXX7m2puaUydP9X4i1vTFBHV+nl
MUqh0xwGw4LJzHYURzfTfvRGRqpGZtmALAUuSTGJAUp4QhB2CmUffS4NnRLB+/FZ
NDlZCcOHirba6vycTZHP0IiPTDSSDnjx1X94KuQWbuvWTKCIN75tzgyLMcctFXTQ
2p39+QGysFx4iKyJzKps/MmS8GlrdOSpmeI1zdhM92iOn9gLt4pkPzEDHbYj5q7w
dff996KqJnCcYcX7G1LlEwhqwvrjTduAEcr9SWFGMU2WZ/jLvXsdAdvkzoMgTwn3
o/CK0tpKzH61HHOi5UStE8xKQj2GRf6nf88If19mavoKH9QdLt94kmjrlSHS+FYu
RcbHfe2Pp8Pg/u0SU0yJ1swZRJa4okU/nMMNcttoTr5Ll4bxRBUCkA79W9sjwPta
kWQIA7ZBLN3eREUfBa6EAPAXZ6YmfBIaU8jY/DAE/sXXZKYED8lHU1KS5mJ/wl6r
6U/fVrAC1bUkY94BafLh9Xw1rRibeY3t4brbry3lO5A1LMYVleR97gGwfQ59cfAD
JcJNWxGYoAAJ8lamHwM/gQPltF/kM4uIPKkMRGsEkoYccHUc2MhA1YYFsOEmsRPK
b7NpqDFMNn9kn/T2VoHP1YLEbaPvfcfxW9zDwD6EaJcNMTmZ2+yn6AOv1vz2pRqd
YgHLK4DWY+zmmHvjvIDRh6vamsyctB46m0C3hcFHHQOPnAOpC9eJ01Kd4ctqFvHe
8jsdJB/fUQCQuwMNZ3IJzE3j6AddhufDWOO+CsVM15H0H/o0QnPnVKbK6RA3KsRK
PWI/6tQTfuhnRbyBQA/x3ol0RQFBwUAtUJdynHX4axD3nXODlSdXT3xFwBOeDUd9
kuGmO054aanL0EputhxFWkMgJgIGZQjJvELc+trn7XthUwLPjRBBO0oAb8rJ8rX7
mWhDw3Fb9GhGlvexsVxjawkwyRJ4im/XgjAUhNVWtyEn/OhFd65l5TUZ352ldHbv
6G7k0yxuF2gArcWMdMEG9iepnDlEiBLKZ3ueV3Jrnn6yGun+ENVhF/rTyrupcaqS
wFeiqTnavyDAECMcwDFVcmGyAknTUJVryuk3WUh2DOnty9P+1eWt9QUm3p3ME5si
YEEE9gV1xPZ/sBkyJaf0WgNlmqOv0FSkgXD5pAqynu0nLPK+RP1FN0rvlA9mf6pt
cNgZBrRJ6O3BXEZNd2edFg6eqtvzS/j3CfQegzhtTmSeyBgai1TBIubQLAbfb1IE
xJW1h8AEVd4et6mY60XyFbeVbc6Kn7DGcx48ztPI1FkAGyDH8ELRQ4nIcdmVloJ3
G5FJrKRLGrg18b3VU6kMgSIyeU6A/QgRmlwNi/nfi9ppHhVzqA8cZYjhhFgwLlFl
6t5cTa5ZK0GsMRT79MWoHdODRzj1Ns1+06f0UocosulSG2Cj76GFOVmcwqbwjeIM
cTmDK6F/+oLC6ANQALjwXMoORAr7/r0xqlyXBk7AALTq0fGYtfXL3m33TEuXk/Rr
OrVi2I84iKMrmumaK/AKs1g2tVz/iYGZiAEsT6xQyNCC/PUeDrqUSN6cWml6ff9k
gJSXT6E9SVlZR1hVR69tPldADLzP9vLmPyGxKn3sRLRZYhk/cdepfcpmNngD4fig
xcbfzOxORD2m3ZnQ65yGRyCvB6qFwKmx4kFJn86vfWgOPTqbmGAhJdkrHCAtnq4c
ohs1Plfm8YhPC+Y4iZiBhj1cTk683vzA2rpenNukMJwwPAivqWIKnPLzZUyDMg2Z
yFDGOrNy3omK1ppv8i+S96p8LDvJPnWlGpCq1UvrOCR2Ysup78Xq6E62g8wd2w4w
DKCr94WTVLysQm2//9E3cqd5IFmhCdRpHnrFz5NiPrno3G/05n/nMRtuyWyEhgRB
XYHykBdwPq9oqkYWBn5+mpaNceTRLns32GHQ+LoloC55hqb42m/5FoE+Vc+1e3E4
r4nita96rusY6Z1UU8uapjOtX3bpSG0/xOj+2GdKUXFSPjvwglyvDVvOdwo3SPMK
8mJ+uYNw2arxzOD2vRwKACH+TfMci/ZWfqHOotzbs9qQhgza8qZglNPFUg9oNI8A
hEIl839cjDyYTzjY+0Ekgrl1nuC8rArKkKWG9mCHUR7sbO3UaMCftsnTHGNTEwn5
NWQiE+QzIpm+sLDjLFOVyHcxKRW4eAlWLd+kAjN5EamjL/T4uOFS1zQC8b5Odhzb
/SL4tc8WvTwho/LelbgbHFMwgE95e3UXVxuJQX7QSlgNyxL0yebSPl2vX4FP291n
SnA7e2+C/wIcVU+N0sp/xtyWVebpPUZoiIRR4NN6TOmN6t3Kh1KDQaSdQNptgzh+
DlJL8gb7HhzLMhIv0WaudkoWMWsbAa0sObFTGGA4unVrEeufwJxy7xvsNoygqj2z
feYIYryYU3DdxyQVf7NIG2M9k3wcEgvv/vwX326guK3AWC9bkK4ilGCR4mmFxB+n
G7EPrTLoff01CMYWzHy3IpQvMX57fJ93J1n9TaDDwxwn2f+vyoegX1bfJNy17Nez
BpTYbDSDVy0RDAqyfUm4LfhjsqXEbNT0QoxCRRc+nRwN5RO3aEzSmFSvOd+8TW60
Nt7vVpktht8kcMidzY3I9IObhwCS1dEU+vMW5qP7OZ90pLgQ1CJ4ZOtwAEyMJrJs
q44YFvSD1eslxKsXnipK+r05N+M+xoDDUFptICQi5VQ7DvMFVp3smbBQpq6k8c3O
nY9+7HGPxozENgXzodnjdWmPGOWvniILob2qH0qWRENJMS+ABnPJdHRDzDfzYKl+
tNQ3QdnvLmU9eQBRG7zI9gH6i0bkN+RBd5OHkFvBZ3K38nDQykvYRGdL77Hprfz4
1fZw/UOX6qVbOnfb1aCNE74CSlFgVoswdDrhANB1Xgd5ACh3HY7oHQQw/8P9rcva
QTr+H0HSp+gtMOxjo2yYJzq8LHhkVMbLnbRxiwiq4aQ9nUiS940yplFaGcPfyB1C
9ohk+ii98IB+OqezghUIcN+I1/oMpEA5PPD+0+vAPDtDzOodtr8zTNdAspy1pB5e
wqchQQyDWpSdC4gvH1faf6zQloaF1tdBQs6XrVtVJ7vKsx8VwNb55fhX60TVZpx+
DQJU7DE6595G/YsRHuTZKrRd6H88glIY7r0mbXBsXhpumM4CG4/ki42vtFB+K/Da
lgjNf2z0HCAMzNDOkHA6/KZ+xrWzNynfCuzkQQT0wMeoNXBwsovoZxIlfU2O076G
QKkUuh0w6FJn3IifSfSMg0DrmxBvk9AcedoAXX7nFw+xVJrrDkYO8vt+ERSgOep5
6frfaXwYasbFLPNr1p9o0w80PnBV9ciXJAlt3psaaSERTUg2qxPwQunN7GFTt1aI
dcdLuOzhsCKKGh6vwbjUSp50BiKoTd/v6WmPF/LvNZKeNYiRU7+bRwvCTNJs/JXI
83lLdFT9cd/uFxI3DpAftuPNygCLKW33UmTdvErzuWBuPsemJA6wQhyeibIjj8tZ
WIwWFOk9BeLoMhRV8rYX6pqF0Zl2b5K4aQBd2D/E3HbJN35JRozlEd4DjI9ZT3wH
Yoi5mJDSnzKSilGiJ/0bIsy0W/gL/Ls7keSVbgVl0XAYWlKagVaL5t+fHKYjImOl
n+TiJHu+fSxaiaFm3fn/JAILwbKqxMsJHLGcbpoZ54Ub/3As6Rvq5ughL4JPkKbb
BdlRelvWUFGBj/GvdB6VihlEmPckzUPiky/+TvFfMm5QLMtNmWz9HZSyn1v6hNTO
w/DJBLcAgXf1bubFs/22OKqrqN6fyQ4NBRsgqWWeluD7yOp7QjVM1Jk5Vq2VPzoY
UzC2FVsPaUasQGQ1XhkBVxpLKWk1mW0CTy44iaD6rNr1gAiOyta31fWlYa35eHTK
tXppvhlIMHgnmCVHpMHQltWssog4ltJi5yABf2NHiMCCzZwBdDTTLrk0UUfU8Fwb
b3qPem6MgcemScStAPahw2/pne3OTSRs9mfPrVAvUZZDuL0Kojiho0evZwNTjIfA
ecTSZwYXBqR1E6TlyP6ecSnlNvVmVxyhn37Z9IMzNAPXX/PkRTmKQ3i04M1boe5i
4JkftB6y9ybbzI3AKD8t3mVGmw3VuKGPSE6QS6j+J0k4522iEcEio7Qe0VL7WubR
pmEOkHm7MpO6+2RepzwUV4ZBmbImxtvt6AjcwPQFsTVXStHq1KzZfzcOhLehIB81
KzpXYzGODixNQrcOMt3xwnPCnqk3eh/0eZ2oPLS0on06EYRH5xL0vrDi3u9KVp6d
+dVMKn5Z4sTTQXOEmh9gNixMqbUIRYj6mIWdgZ4dk4miksd10IdVpS9L/xgoB1rB
sJRkWWcBdvqqwOqbuOJ6I10QamNmqr0DJU8nBXjNBIbn/qjO3qqz8bPlhosELkg4
lIJ2JM5cG5r4q+Is43FBSgK3YMPlgef3pqaQQwZVVoyt8azf+BFm50oO2w4i8OU2
wIVXwgFVEccbm3twykXXqerPqX0F05eyoVJA38uCH2J5miZSyRGJjTWUdTKgHFCQ
uszsMy2/ZKWvwYlVNlSaeylinMtGOZqmaeIo/93dAsTSJJnxK+YotaHW2Pfelq6T
vykRCVxKm4lnr0kpsLsIfVDlX1scOF0ydm6Z9u5VTEwy4/FimrGSZWkeDO7xj0Ar
VoC0ATMZTWH9/ZM44YzV82W98okKSUkc18/LRATcwQxjTHq7mHZESWmOejFOni5K
0wzFm/03a4fjjSpuiTfwAnrSKGTCwmDeAwt9ZGig4jp+bZOGucoBnnesSDoYm6Ff
z0ab3FAhZYTqEGtOrznFLYSVV1wFsVL9PWLfRP7UqU+8TIdAi2hmtFQFoFDHs4rY
cy5wblGvlzxokq6zPTPaxLyY2pqrey8EtG4/jVQMLHkCUJWUrqzmNBTH7+6mfe3Y
N3s9eN+vSLf5WNlG8tGzg7+Sx0gz8x3k0KsyZ/yPpenPVlJ7OMdMRdxnC+/5f4eq
oMSsjJuBhQnbISEJNFdisgRuPSbEHO18WzzzkY+VdLQkEouPofiRn+FpWIkqRmOF
XbjZtfYsnVAb/ZBI6TAH4Oq8PB7HT+PWlxr04XUoQRNCMPKUejaFjGKR/ApTus4/
aNV4wDbG8hYwgL3nlf9uxWuAKJeTxq4T3uCL89kU6Ap9fe6Brqly1XzlgzOsdcYi
dN29vHV36UPtJR/ccMEV7RrgwaWK7TwAvNtPFPbmveRjgxuUz8R5tYGUDy5VTyTb
d/aDXVWZ00PkL8nUhJLTrBn+r/iqsFv/IJl0pgMRbbEA5F15SalaGCR9mBueqJpV
O1Jcbta+3xT5DkKzE6juuSZmEV+sexxLTik784dEWIgOtLglgtcyDYkkbREIwkci
64hJF/K6bQWp0bEkF0mi8U81wvn/rUYsJAUZLQ7ISBRo2DXgjtUGzZdPeOVXGhuI
vmIJShiBhTiYbsLaGAsJj6yP5b3UyiN4SplohjckFOTRsgIYhtL66atCYpsTaozf
hfySIfS8Gy3PwdM+rmNjtOud63kww7o+sm9fAArUsUMsXZfRA5R4467MGrVlNggI
++Z21weMpDWDGxlGtOs3C/GwTmUOZMCjybRTNX0QZQdCsw3DvYGT5laP0/GBkYVb
OLauYRFbcMHzeBn26y7RatBIw4APq1TujeSaBO1kJPbZMCOkb/4ruzOdbfIRUX6L
I1s+vdWYF3VvbCbnIHrnYJ74onwBeD1AJJUpDc4c446DJKXp4kA9N1ZX+ExDs5F3
FU+/vHdo1MdCCkNCLz4RZvbMMhltzZsMgMVHqlA/7bWOwPixWY+lTY0t+l0rg9P9
Zn033/40+GiRVLr277c12B1+imISkL0nrdDt5nb5UyELJMeK2leV2/kedYAZhQ1S
+0vvPzZqcIYH3WqAHZawF077GuFo3Inexl8t+lTW0D60NXOh4Pc0pSd8G2Yzz26X
W7mLKm+cuPVC8FPdLyBy6qTXEB1mevqcYtaM4gdddtbWkdLb9XC15L71N4MBlDhD
UgXRHgOxHEkjfl8dJMI1tkWCBeHZkrWk837420GHXV3sGn7xTQFKPRki7tNP29qo
E2rojuONsmebvDLqEtrfEAnn8Q7QbQyNbXUmqBctwXupMdA0Cg2QZ6eWndMOGmM6
kWEnyr+rKIPYVGiPTc49eD1NbOzKplGLDt6r9OyD1O9MBlFNJfFfq41ie5+AC48O
L089n9e//RUf4FE3ZxoqDkmYZd8xt84bZhwD23rhJ5rSr1rBKpMW8ZhsMm6sXEWf
r9JXaSmQOC4ToFOQJohKbtulQQLx57+bHjpglWa6gWwVKLQ7XW3J2dDQiaPGacv2
syUWktf7HbzpNK5xsovs0uaZmtkma1RkagCDx19u0roagnH6AdbUvGwugrSftx5w
kB7zyEYe9OooJ259thfVrpmJP76nCzcT97WD17nj4MOtZ4oTvVJUutJ5worosRZa
WviAue7yBgxoCPo0QLirrxAfyn5wHr7+CbDoil70VjoJHYstAlXD32T3X8BW7/gE
MQZxq2HU27fZsj7sAktfIT2n0PdJCZaye1+WvxKgQOKG8f4HBtzniFEtU0VnLVi/
wem1cClny7SiQpVgiq08w6HiCjwycJPu7wDlpD++x8Czoep/4e1umHJ3zLIqfIaX
If2wAQFUxqHZPfks5sZJHDfNTuN80kD0bQOkxhAhCH7TZdLAYQEwSfsXHh480cqD
CgxdXcLEQ73F8xwPdi9pD1hIXD0DMDNfDoi5sFXimHeevbbBXkhuPYcQ6euszNcI
RovYs/upUwDjqcVqe42JyxuyAjy8McHAd48AntXasOIYKR7Z9hlcRdcEmwEYd/TV
B2oSr9z3FHyXYz6X2ZU0H8rvZsze/h3LSaXAb1sfC4u5zmjanntxW8SOz91ALDGE
kBv8J1PEKm8lawWyM+XxyRKUzBOOUImN7tBHt2l5J+vE25/9ZAjpQJU8Za/LKgTr
P2yA8HFt1WR/X0nDM2BwnNJFi21fM+SIduzjSeQZr0ReSDXJmOgOpfiDOJolFMtT
bieOPy65RvSDE6pp3pRA87/ubg4lgbHwa69MvZ1w/ggRXnR/PwhCRDBG22gS9lRp
3JCvUsTHKkSY/kSNodAF4Ssj4K6yM6Xmw7THBQasoH9vaWGar/BSQbaqIyvhKnLI
CqGAFxEn2p2No8R2UjnzBe5uixBgubq+3xte5gr7hD/w19XQcZZiDg1PFYEEz/El
jl7QWu5rqakWFVksAlM0Z3IHFMyWfMtpSi+TS6kwpaTwPY0QJGTvKzHNtM2GqSeC
EweAWBcyr9Q52ePiotBY69CinAA5tUtKSxmKlww+gZDu+u370HBYTDWSd7wkyA+8
WioD9g+a0D0TSK9kdxufnAnx3n6Ks3QtOJVtel7fYGoY0WYxebcKbUMBJOPMCy3F
kJm4QDjzw+8c7cgnNB4AW9n6AiCX+WcOcLGotpcPyy0ab05fq72kEluQQ1hhFMEV
fpBx8xdZsM37wBzmqXjDC2uMrErgtN1BI9UbLMsy2r3LZpFJLVkc12anQMuZiZMh
pyXgARtrhrFMKjkJ7yVlVwOEK5EmGIwZElDEBhJUPv6ulYwrreE4Np4mRsfwj8+X
XkewIBv8/RtGJFFazso0LKxdcbhivq//Ssb/50FMWvPJLYpw+ZaSLl+icdB+vq9s
HqVo4I8DYy0DSiu59hwzD0v+ixFnGCpWV1m4qwFHClU82m/07xNAAd4129TvyzZ+
a8igOb/3m3CM44wMDS4OD75UrenoyirKLmkfhD9azogdlcbgp8dm5KWT2zS/H9ny
648rXfWla+i203AW272Cmv7YMugewDqMf0mQ44kTD/uuRY0htG70d3xEn81ltf5f
XG06saQe89AN9H5oDnZZiUaPQGkvlt2eeIt2lJjPU+F0ZzeC94Q7FPSyh7F2lIjW
yhCsomiK8CESYWajGrpu6U7MaEFfGsWZvco8n0guGs/D+mSqx9vr8D8XK7gzfhKd
5tF6jVnECmp6+VLxpxIdQzvpb05myBhE18O8+XKLY61PcchgLHY24Qa05liNdybI
XJ/TP2NKq52dGPkVh1t/2kEH+XbR+e4ZdokIb4KxMiA8DO8/AMeuLH5+wHBF6ybn
GpqrMglPnA6OXGZmn8UQjA==
`pragma protect end_protected
