// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 13:57:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nVuPDqTUCLwQlmBIHpYN0FbPKNn35cndPftMeY889kwy+BWIsr645m6oLAimor5u
hcb085j1g9AM5MhUyCBu5LEyTVtvNGvz96iWIQvoFF/khzqJ6NKJQgn0jpO20n1O
dEL8c1JgsgHE+4CI6fedpBboxKNu+Aq+ErUpoxKGb1A=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19952)
2f6MI/mZuvbc3Uhcww3xzi4FwZxDMHhSUXhf3RXWAu9cq2r5HOGPCkrW38zLbB7i
FrlwiJEDh8zwBnWxuuWT1YBN0nKiJyqsiLH5SAeb9LicXs5+vj6JTxu8FaesyqOL
Mrb8sUCLvvfLwuJ936nGml7vIIL/C26+ExekphxKuJ1ppIDLgBEyWnfysqLH7EuA
3B9h9MM2gi9y4HV8rXSc9JPNf1B9y5KrOW3gHtDaLqYVY8aNrCrZXeYh00XLVYaE
Z/EtKgyAa8877TtaqC1yxpUTMVMBQfybOM5az1rlDNnLEG/stkW7KajVqS1InkX+
e+ZybYPQg7kn1/bgL6M0ctqNwif7jz5htuBPYyXoBVOV7FfIgyS4CKOOOhn5IM0A
4e9F0R7bX/LMfkIRBLzMs/v0iHIM/3K7PhfISrEK89oE5cRIHbjVtRH9+Xjlzd26
TCuW+y+YmjTmGYekOXosSiLwgisZ7xtFvpw6dGF85b1EkmGtZkY3l4LOEW4WQZF2
9Pw68qqXvoRLWnN7mOG3rNx5iV9IJxYhDLZAUfw03TRYgM6fn5zXa2fmmfR4/wrQ
TYnChREpV3vccqmF7eh8PcAK2g85P1+/kfBhhjHdKWUO5VwezUHKChtgWxvX2azH
/dN49niKYqnC84ZZYyEpH807aC7VXblfab0Dqw9o496d5Olg8UGFqSRN+6IhC6Pd
T6+4KW83MaIrP783kkdzUYT3jWTGQCQYJhGrz+dx2+n4g7NTYwiiLKlo3z7yBj4w
CRgquxWwdBvPjdiPQrwFuDeJvhD/JdYNPMk6Xx9R36Tz4rLLeWTKvR0YIdeDmphn
frpSZK1opiezROQxFQP2dKBlfxfjHC4tl33oQQ8J6YP/YR8SO+nrnHVsXpKpuk7Y
sNdBTX0s9e2hh+qWeNnvIAIB0nzVs9KP1cIkui7XMT4MOYXfSsMwwEnKGBnAyphM
a6mMAhcoZPZBCm9ArRwlN9lZC6K0n0NiDTGkro69HprTXpsLfWRSuwyNEC/SwRSc
KzPLqOnjQ33jAxCW70kltVG0zzOi1CoS5oBAR7xczXQ6siI5PECCz5rkpIE1BiSb
3UCH+WYsFqM4WSagm9v3q/KnyjaHcwbQbm1+WO8XosQaKS0Ae0gtHeihE0GVVSz+
C15l2rMh6kj3LX7/AWecfgpCY/jATX84aCu69JQ1Tz7rXDwwibvtCIY73/qMKGox
OUdISV3A6xo3fJFA3T9GZ9gRnQ8udNGuqGUXFNVcoocc495Jm/TxrPITLYP3r9qL
zGiZdSHXeIz6dQlRhbSMKtwjTJmdltRSgnM50JjHNFqk2mxtFGoVNhY+23zhvYo0
4kgC7m7ZG0BZ3wqseTyBeedK2pTWKEO2P+yZeFNgj76P6IA+5ImALBoqK/SvTDbF
1CxbWGldYYHWfxZDuWdTkfM+Fp7bIFCgQ6uoTCX7jzNBHNgmmXvG0ys80gOwTYi7
lt2wQoQGfo7XAVqlhg//rw66NcQsc5p1VG5to29yrmJIQ/mlEtCWVzAhrQ865vXB
NItI9UjtAe2TtTP28s/rt5/KlhkxOvZSC5lpUybTn+zz3a0Jy18aD33rnOSdGKWT
B0dpnWePVDTq5yJR9ZNF/2i+AsCFxi9IHmyvQloVBIDBZmgGRFHazRjeuFr6wgAh
lKn4CCb9vN4smIohcydkfbFz6D937wRAwsDd513R1cAMprbpmCkJAWfTD4p/mX58
656wmb1Bh6k4l9BXFTY6waGFkul4Uq7VZO9+3ycY2xU6cxqd0YBLz/StiWX5KDDt
3o4GcVsxx69z5kdVUVQm8gJrS6G4eMqaZqS9jp7v4Q+7VWp6IUZ8rSTTR53rhL60
WJx4WJyKvolM7wYtUHZO3myCpUiGn1zbN/Yp0Pf14MmFKWMfxk5lcdiSsfxPMLGK
AxPS2W3djWAo00O+3uShWsAw0576YrxUJB8UAq+qvMDEaJZVG09ORDAT7NFEKs7o
QAe5dTbYEdB0FPsGufdRYWLDEd3cEAttdI1Di2qyIgc6EhHg0X0Hg5Tao6U7R35C
JGbdUrPJ9FLhCJwCWxxYDrJKAvehnR82LkepYCLYmsqU1Xrul24C+QwzN5BxuhDp
6qNI4ZLFZ//td/05vQ4iNgws5v2Q6rduh+1saNMOR4BV7p7dNRluxPoICgf4YHOQ
zoJCihYxzgMj9k+ahWxh3MxjxQCjPkaC9boqszUTBLeXYFeRAUeN47GQ8kXTvLDX
QHgWqV1doY3fRwCwQymCDgNl+KaSkO5uNkAqzxPWrVwSGTiUvXlHh63YeJOeivYU
KlP27M5EIQXihm1g0Rd0B1p3A837vc1OqmoGp+/Ggvcjpwn+WzADQkR+qq/NmuEB
EGLkl7jJGizUJksNNla1k9/o1vuYmhg1XGD1VwjoITcssvy0eRFHqGser8MQria8
PXDE/pguvwEHfhZ1Np6GL9qf35eoVMgxOYduTZyye7jFbtJZeKhKmxZFOxrU5VQy
0UZo3yQ1NenN66uGvd30eOd2YvfkYfGuc86x3MUL0Rvi7PTSIW9TOftI173YDonk
lsTDZggzJa7ObdiloCPAC8/S/4XBBMF91Nq3jJ4O1rFL8O1se1hwfXross31WT3R
kYSKzfXHCHT51Y7OK2Zo2q6HNjV8gFi4HhpqzNtsd2DU/FCjCnXRa8kxNd2z+P6p
noXybTCVbPvKgMhflAfa4jrY92SOWKAlYBwztQbx0gyyX7xLJC9KP+m38sDCXs7R
TzuRlb1Xn08EDjCt4bZxK+2IX1VJuyDnlKX9jk98nVL+0H1enD59SRXu3rk6BKbr
yhxyfpmya2jA7DRWYKLi4MbkIN06MVRk/C+Jm3OubjoALzweSWQp6sZWtalxfTQj
eEJim3bh4mE8/BGFEIL+WWQ4YYS72TC1oFhjP3qyIj0YoiEHPgXDBLhGfcuqEo2N
iTiwzzpx8QAGdR+D/OWpg+XqDyWR9dE/t7nXJLgcfsMTR/jG386PRCthbQIS/fe3
JfEl0+VBj1+fE7bZH9134Ul9zhivU2waSvMpKS4elCGerc4hgxFCUt65WiB6XVuS
XHk6b73QgSOWdYOc9c40QI6D83xDlDYoLk7Tzzf5A7DYOWUjgJ9vY3IMAnGu7Mps
gYI24QrGBGNfhyiqOjLV1ZVk8KFZnI+VACo2O6iQ9zdSPA8It5qQvhoXviFdiRrC
OzhyNwxiWp7yDMc7goZGJUxFGtRUpcts11W33gRjsAAYaFQ/TsVbH/KaJUH0QxL7
heAOnn6daokqptj/bgmkZECzpuVnKMWMOmyo/UqZBrO1vSMqtGlovYAcf3Btkqjh
4a9xUTrc7Gpvr/jA2bfKloZqnmvC6FD89ZxyGaR8OBUdqDfjYTWunVePG/WeYyaD
GBbmqXyaWyj65Br6K2MQs9VihGVWdyanTW91yas65ny9+qlu6oMA6oQ+GBx1aNaT
R2cZVauihSoFAtYpUFp6aV1cj29JeIvW9rNPY0wUNt7TjfOd3eWq9SEuiHyeFE6c
IFnyCpgfkV8DyVq2KWU+DB0ebssI/vYAAs5r0TnFk/N+F/BziDeH8ZCRvON1i4U5
EKlVxHC3+gahhjnq3auDSqQBC57bGr24Lg3ZDKSis0XeRK5VEd9hcD1iUC5NJ55k
spmfGUz714gY+qBC2YlrSUWCe8QfqicOdbOC/HqthP1Q1AVIiTTD2bvIPiVU6PD3
3YypKlCSLIJGNQF4MA3+dctF3yKgDwFogP+TW10YdwOBfA2+EloZAmNV540JEhIr
215Cbew992Ph80Iarcin+aopUYthbF3TOiNQuEq/7nhp3t6+XTWXUQutpV2sbaYL
cEk06wKeN+ozo7qOTztj3IbrIqHEl3V2SfBGgjXSTJHu6ffS5J/n/bNUd90BYtsS
TwLFeGdGTfhZeEEOp6jMz19kbah22NpTDfc4Zf5/Td5LGlyblV6UhAjqVQ1SD/Bo
koFhDMoMpfy0HllbAx1Ix4r3GMWgujDBJ5Q0r6UKsdzkBP4qq2EmpjmwsAR2MBeF
8XBSdBTN8eFqcI9kunZlQwx+KvVZ1Oqmkuxb+EZpwgVCINTcVTdoAIz3ObL6BQmr
6n7PMDNNXudq7gjvTXX4qjGYUX7DTy5KeDoVAiePFFMIkCwJc40GZhQUub+ennr9
gMFhpx/5YPNvo6xOCcl9jn2rGs0c12JfFcd+ezCkf8iFSKFcEYgLpwnIxzJSgRw5
MgYhhva8mKEvwydAOLh6WNx9ANhwU6vCm3o9CTeBqg+xFRoLPomUAEqWjEFrDsK9
Ii1B7NzzmJ/6bR9zJMw+foHvKaoFkjovImZgyUZSY24fM+R7aAo9nB+jLBpUwdPV
8m9kZs7lLYC8fo9432DZgg5eGhK1Qp/mkgMPjuQL3LFLzXYdlbwtABtYJMYouXCz
BSdfAEiq1PfuxBvmsZqePQrZj35EH8YoOPL4IwcYaLUeOFuYRpNKdB3mhARpjwoF
+LyDICV5lhG48thfoo0IbYQ6TTBnGiCIEJHXSCDRYwyl4hOsbHlH3ZDR6JmgpdBy
8CIMWA/uxLPaDjAYn9cMKD5yhsrWiu9u+G+vVV3DfCdB7JYoqbvN8WE2EQuoo4mx
KMymMxbkzWo9mAx3jqJDFuwszSt9BjuLs2Rh8CRsZ0LT0VN/VfCZ5URKLGsgOKfK
ZkuMq9kYdG7ffZYQHOg9tSTTHhgaVz95I2T1oFTmUGTkQ5sAeitiWGrLcGpVterX
j/zVBTWkGkaxp5m5iDzyhGGgl22YmqWdVFzw7UbSH+epq+hB3ZSFEMzyeKQThl58
VMbeZHs+/bbb423yCk36OuoyzFfD0VeKd7kqmMelWUgcCYyj/DWZFykNgWgBfuGj
CIBe9XC48ZNfnmiMSPeHF3ve7vZZnRvxrYmZJTts8+EfrHwUiCyPC41F/tNka9fq
aVNJglgraDXLHUmioKVmr8ylHzBem3Ne40MmGTlhOpii9gXdagILI6lRPx2hkH80
DAPLiEk0a9osFXZ+cIt4wv7SU1fCS+gQLtsaZOqDD+4Ox/+TKNtPusidaXzUzuaq
EMHOwwb2rP21ddh4gh0TdvTNrtLGCjyJ9CZR9qL349gxcHXLlXTIDJ//gTVHtn4v
Vw/jKfBrMEjetZdXNTmWDRXL/6OETRcBTU+H4HnIQCwNyStKcEiyEm9fGFrWX2q6
UuboXKHhHvyp7I9NX/vgSWFDTUb1y6l+0ExBagcd3tNkfHvESduuQsVlk1wXKTtE
CQK2JMKXGlQ/hflvNqKOJJrmFtJYQMA7kPCclx8PPVkeVk5pa+f8OIiHCedOdpkH
Ig/EdYMhfjDuKXvV5pUea5ZfSNqbbhal1PN1mXNRMkQHadlM1ATImaCdoxBuVjjI
fesmfi2IEOi1Nye/XavZxryICF9vMuaN2Ytm6wkDtLPfV6z+nCzldHU4dhsbQ2rP
sCs4FroNtiDohErMP1qFNqilYWg9/CQm8axbySuOJLABuKwjp3kJmypXcawJD5qz
kUNJq1K4R95UQP6CcN+V1BlVMWwl/FBCLiBioCzcyY5Hpz90dwT3yosR+S00seiM
ETNHR1FK2ML06tXSj4fR74DMO3HJPSPvQvqbUrPj8FevN4esChG5K7ziW6G5hh+4
RaPUa/6EpurzrGBXPhSkA7asAWrlDL5UfOAm8l0E2AZr+DUV1J+A9tpHPjv3OrR1
4lQY9QxjOePaJTcAELHjEuz5N2VsZaLxln9ulV6dlTOTrWCMW8udfgJpGVXPS6FB
1heK4FNLvcCgVeU0PaepsJKCUgxAMwgXrsK8uNwn8DQqwWlYH+q7rXrZOlAu2sd8
Se0sHOtmCXT/DJkASH7rqpL9GqD8gazyo3r2x/qmcX/bM1Dr5EYhlv1LAFrlGNzQ
EHLcUNkhHW0EFUzZ0MCKpTXvLAlZpFdZVaiJ1WDE94PehnwDoiDN/Yt29ttKBHXW
s8OEJ3gZ45Nq2mAZ/smOyGHdRt6uW/Gt2kHdBapDR7c4v1l9qcDdtVYwSUBuZVxm
1hkiH9pLHluuR30AE2++Lk9jLmVl6uJ8x1VlT4ntYSKbztYd8Fo+ccHOPsq/wI7t
touNDwWFzoO8EhLbJyYzltD3fa2vNt9jR+Y19vOIYsWgxoDF7x1q0vUd15LV8FKu
uBOHCfprT+LmGTeWt7v49wDTIi6UL2u9lIXyB/sYgc2GvzsW95mWw2S62HAhZlue
HMYmBUn9BaH6QYRWrkf61SnEXR0DqW9O7N4Qlv8MOHa1PEmEhFcMNPxyS7JXKwFT
+B36Ljx21uIv0u7HehxBi5X7xQDu+s/f6CsdzlhkQZC7ZEEWAW0bJgaPM49x0adA
DNx8NoWUXRTbQHnQIm+x8mboWap3Y6r5jmW4fXEkgLXE5GYt8XV2rJ1wil6Y4gB4
3teaiA7nbbq4eDsjCzFpQjF65e3SHt4MBF7purRllkURJJj65TKjErwtZlO6R6OB
y/SAtubnqMUJL6Y7M7cogENblPwtSDEMapd+1aI8Or3Ara8GO+8HLkd2K4APJye/
nbBQKApK6M2IbsYeGUjkvN1eG7dQ+SLfB97FsOJ/bFQ4iwDQ+XYThPnU883F60z1
e3Asa3K+GHFkmOfX6oAug2LtKLDT1JhszWD3eNDCqqdxr8A7gqJ1FiD15FknRYy6
5kSzyu4JInrkfHSfIadSAYbuJz2u1AvB8pqnnuhzJMIQI4NpAaQg0j58e/sD8naI
AakUMjpUHzeGHOmlKCzoX5pPR4x8qyd0L4Tsjd7k4XdYowvxiAXKGoNtFzv5VOy4
Gtt5CoRnQSaDg//MQ56/qFjNo2MBOqxJI4ESuyciyjFZVaj8a0evJ1JhQ85+m1w9
y+bEe1R5OmRXnbpfmRsuRMbk1+JgwQXwCsTf93znx+Gz/YSen9pYOYXXHYPLxeVv
xAp79j2OoJKkCV0MN+L5UpeBWl/HPyxBA4RaVKaKYrhI/B+1/Y9nFJUhPFbYmdtR
KQc8b9RLrkKYM9oex9S+luMlHMlIDSdtK5f0XNuXttotjr0WX/4mJ0yKBzX6mnxn
JKrYIdRfBbfyWOjO0DPSxovQTntQCEg/O9fyH1btxikQSz8ScrdA4/e0HDtZk6U2
4O06dulYkW5mqltki0ZCFbYBS1HGyi2yku6iDoDg06cEVcWjn7MTkIs/jOVEndBt
l//r7wC2bECRss+iOOUfp+PLheVQrCBP60qUGc/lcGKDymdLyJCj+IwthhN1kAsK
G/C26ruRX7ZEg491H5cJ1LQGBidTO4axqohqV/xdbh9o8pNetN7tlhh0KrLVuVD4
bh9ssB/oxUWCsVcLKXZMkL+/8FGi0+C5/lZOwdruxsK8ZH9s1bW4T8+ElG9oJU6h
z8mquLATtycyD0Mm52QioRKqW11dGLAGNQ1vDeuFZXj3BMhJYa9rthbzPpZK6W6t
dYPozCSyjn4msGr7O7YQWLZctBWfTCikK6g1jFfiE8WCflwVzYvrOkl4cl+LUeBZ
HVEjR1QdA0zWk+KUwf0COu2Kx+7/BpqLgsLWjVzOB3ZJ7hg4yBY6h0VZWTVQvdV1
7CpP2SuQzPRR0R2JecVGHFPw6OO+OajfSTVKj5gp1WGuhd6fid/I4+5elk2uXYqe
YRYVo81ySPHTJTy1zTB9ReWMyYu9S9NCbE+R7HN/NqadDcdyz5+Qe98yeB/a3bFg
L81FTbSvVcMvQ+SpZY/JlHjy5+/vvmA/Agu5d4KAGfQWMRKDEAUQFW5+mLPH/7Ts
ICEo9nt1P62H0BgQaXLEr3fIW2AbmqUbksBKJRXYmXYSzCp7GMFD2Ht2esYWwQqa
VAP7i0hjnj/3cfEGmzxmFgMaE1kEL7gpx4R0l/pwc4vndy/xtQ9TCNqQlUA9vF/z
0xvgzGwC3+CLkLN2EOMNMRGkwcRHQmtBKtHCUKZBAC4oCiFm267e+h+3KNLhor8G
6ezX4yYT2jXptzI0bR1aZDmVUXEQHAjBF/mUvkqDvZ6JR2WMLdXKUW6P6VkuAoE6
FnEp4BtseI+n7M3GwDr3B9X5fZynbDsUkvnXp5DoGylY1zIfKcl8BAy771sGHL66
8rsuk6xirenQye8AsaZF1l/5zqo3vMEVGEtHkKf7BGVXnZQOqS8CNmHqVvfWedjz
zSiWJ96yamhtT8qojwoNCmU3EiN2CdBW7DVH8lTwya9HoCy4sNuYly/zKYv0vQpN
c/LpBPEjHAuLjCKZ3hkyzOq3p2/Ck+O9dPo6qJgdthk0Li3Y9bu2ZuP+2BkB+xSa
h7ieqF6s5odcVI2oPbm0Zo7reEpSjLjoY4OjbwE+6QXjNJMfLf0ZG+sGb2VYue1b
isnjxiOaCPNQ6NXdDq6RIOPJ6UUYPNCO86nlEfd0xwLtvVCuwZdjGtXseb4ri0xh
TI1OPfiNfdcVpOgVwE0JeZBcq9QVbUWBNzdw/e+m0g4Z19CEcsjL9xTx5Z0vW/fl
F4Q+MNn5r2nxKf+k4Y3xDAmqAgDvr2C/IGU0ShrFsLziKOnrChi19ar/p8avKbnA
VbYU3FHl6qqHZA3O8DTu3XAFEBY2GPaDjntX2BuUFGnixMB4Vr9zkRA2PoxBsXk+
/6xnvehhGByJpRwK2jH6SJCS6XnwiCbGpabUIER+Qzb0SJjtxckfJ82ej0xYuIWA
+n1SpH10rNILKLTpEn4FYRe+Y4mMn4w1TXRblU/oAre+G6D5bs7IQlI4rQqXatik
bFGMckQQcpLgRyVAzjPEIQXc8N1qfraBq9I7oxm8T8LA7KU/uU/1WgP1QNzJ9hJQ
dd8svbGGnFerqwW/YUrD5UksW/XXGrl+OaGOFC4D1IBgrX3F1BUAnwxnG1qJU+hY
0SBiZ5sdgOy9WvxRNaKTj65XsMt2uL/cB4SLbx5iDNZvIY1F/iKp4PFHioy09pGW
uROen7/+BnWxf5ARh38f/KcvPXIEvr5A3jr+3FgSggX7UwIs2ZXmIt1fJPDrV+UD
bXHnW0ZZe8+VjG7b4VI8vWvMSwthDpqEc2PFpGVRVLe7dLTtFQCkuux78oEON5Sy
q91m0pGqPaTSuCLEcLMlu+dU6JQVumVVwBYEU+uuh2SjpOhZmgBMXKen7mVMAhde
/y+9KQyZtUdrsUDLS3lvYAiZye4bGte+4/bQUzS7yCjJHKkJF3SlbPbY4qmPTwDz
5ePa/zCbjuxHuyXtdtwlVA6Tsg+eXFB0MEdeyiyUJ5Bqw+0tA37UIfBUj5KQn32r
U8YggyU25mTaJH6Ip9LF4RkVnl1b5hZfoWE2yW5y/bCt73kyRvYaibd3s7O1fxCu
oPu7BHqfsMp8d/87q5wSYWNE6TszjcIzQp2r8+88YtKZVJjrQmIJMlXoOSE4rcEq
GSscye1FAqg0/vw7xmANwp8Fj3hDZ9XY9D8JhZEgpQzLiSat7c5Kxnya6j5/Qw3R
EcAgCPjixKD2JsvXu2niS9CHWqA16ZsOt3C+0lY3DK7u30v1YltfgxWS896wsdcn
S/CqYPlJS5RCQUi+BuFgkMeXZ58fhBYG2YtUSO/zspqry77ugErfU5MdriY1S97V
oi9+0OAC9b9iCURwumli41HHKqB0Gux5u5pcn3ICY/4T9zhsd4KeFlkVrHpcI85t
ObFbYJ3/wZrfEgBEX63gk4DxrRb9rMXizPr/V8YdKXrUmf8rRd4wL1hCnyFObIxg
BSJIUUZAgkF9nELJ+pG2dJYgx8w6Iq4/KUVHZOwaTyrejd/MRgV4X2otxQqdB7A6
EAumzgdvTvy3i6MHoe1O9BkVM1JN19XMESHFeh1mVxvbg1w1p5j0jo8uARJMFHCv
GllH7fcSZOW7ciAurJEoIraeJV1goezsIxkLpnLUhks2auGuCyejq3/OuEYq1mqr
xttIP9SuN/z5ztU/vm7KhJaYd7j2N4UkvY2qy25PGpmLKb71vUf4OEp+C88xcti8
1ZmknlZA52K6/RRIzFEMtZPkOdbSnh+/sQgYEaU/jSzPAXZso+2XPpDbqn2Siu9H
QvUQv7ybOVvT7rF8D2cg0A/xYZckoL8j0xA4m8uKomMfRikaWQ9KISnpUzoJ6q89
bysVJkzJxm2VZZ1+z9e0WR+xeAMo0OE9IA4evIF8r1PPN1zAy6ey+U0gkI/H83Rf
PdozcAbMJ+xe9A/z6Zux/zHaOFsqjf6QbxznDxu5oPOhdUQggBXczeRN49mEpFTr
rUobsPhWlioTBkN2ogl9ZJSFtaLteek6ud0N78UzyYwsMoLlK7OoPTto0DcxcQzO
t9EfNQhspj93ZAWWpuqUeRnHtCj+SVPj6mq5rmKq23zEWN8+rRcL4nU12rSnGIrq
YMi/x3zPy/aF6WrwBZ2pnrnyFOWwe5Osdem3hsMc73SLrWqIOZBkQsNiaKQezFC9
XsEMHETR4GeWDxv5/JKY1zm1Nt0ConS5a4rXZfjlJ/wLqeI7u5Ks/WyE4MQYSF3W
+J42EbGn5BeW/T5h0leOY+P2TPqs6ehs+OvBWN94n/SBKyw6E+buQO9SzfvWsnx5
whxmqByFW3gRXNhW7XhJKa0uOMeY425wtBknRuccaskyfZVfrIAme+q3rgFa4sJ3
CH6RuSsTOZm2zj7TR0fjKjVYnL2sAtNz5dlOLthvACP6FZTJ+MUufDgsAzv9nt/4
L7Z4wJRnsymqz2UhdcnNEyWnsJ0Y3zGAYXj8sVjVk7ATKRDeIdqHqkBkzXuYgQmR
+2tvH6MfRutzkHLX8Los9tZOmvDsLBfsgXJq8ZTkP6bi4IHJfVLPdHAOFogxO2BZ
oBcuZvNbMeC+D7HtrK5uwLgb1PXNooLklVQq1ToLtjlKm6xO96t8k+h5cQZflOgE
6OYlkbB4mTofAfPUV5l3QU/cePHBtb5kqIfUloWM44skdznOh41gVftN969HoFQ5
GdGGvAdp4Jui9fUOuXkgZRv7N12hIKrzdIQJ8NGXimkMnQKxul+dobQoM96tD/RW
ruddj053RNaJffGr0iIdCU9xwgAw6T6LAoyII05cTx2TGnV9/3e8BI7LYua7AS+e
UzwtoMxIwuRXoDQRPWpYqlHSD9bHjVeGzADzzt6wr5zodZct5BaE1y57w38b7GTa
28sM9hkQ92aKx+iwHdgUA2dP5LsRH+JLsyzFZD94hzJ+iEU3BUAZB+1apRxzqFyO
p+3h1yyaQLaO8F/Z+6bNaX0PDhmV8vv3R7LllI0IBAhRtYbFaONJdWrS/Q0ucQi7
AX+lxUDbji6WR53oC06hYplOGhreTyOGsUt4fQs4kfLOGozb/UOF/CC7memQN/uy
KOWqE0mvhFmM59E21K+d9ojh/gON+Ak4Ps/wHdlKLGSDEaaO4AX51iECv0UdYv5j
yx5q7p05UJQDiaa4MAmIXQ20qTABC2PdH18lacl4B4TLZlIx9NgANwAmKXzoziXu
PZ7FumlqeUvOs2g/yJR29fH4rRWK7AbypE2Q+4duzEsy6EuC81DBNUYC9xzBQM8O
/0WPzapRZGL7y5sajVxYe9r/Y3e2fBXR+mC9Ot6WaG4Ci9AH8SHZZPKABiKhb7Ha
fvC+XpHlzd3vvRmwRoFXBv6ZjkylrejEwH2tS1t1UuesjVs2C2CRIA245l6Qut6x
m3TMPYYi8nDcuukmYKwMOM/+07xeuuLskU5WOo2JC9IAnbEwjWw9W6+wz6RbPtPc
H+M8wO2BM0b9rkll7BC3HzqA+7evkPWysbsTfxPVPklj6znB2bKnsM7sdt6qv8Ey
NGLYx0W8qBGXqw7MLkv+Rqxvtf44sIadg4w8nQC2xTQozOzX6OfEgeLOpK83Ba0w
y9jsuo+lBrL3ynr4KvOv0uO4MxmbOrXk+VSjKgkZoIG2SacpYDIFIivbvB8yate8
WxjMwegCEu0oR/o1yHxr+v1stDbBukWg+oGWvqKd7DpeaDbT9lDoOOBZXBSThoY9
cqmDbs/0wFcPYopL295sekKoSLoblEAMAbcjHfnYFH1SeWxP3F25MMK1dwlLaJ0o
7Zz9RV/LbfpR4TkqHRlzljrVaq7DmqeL7lFGuISdgUHwmhXmpmGac9R8yJxMneeA
PUn/9COuTj6CwWlX2l0aK1sVOk3N5lb4qyyHVco2N/5d5dhTEEtXmv8qJVbIcSGa
Ri9gip0krlC4agLtsoxXLGtAcxKV0SoaOTSDno4JCdjBuGj8ldBkZBIrOIdgcnhv
M6IZt8jjKeH0rUY9b9LRIQ0PTznuUbAiXocdtJ1FQrEIQVxgyyXoZZotJkNFRHIU
9TF1nymSL+OVKiI+ATSOahfxt/7hUbY0BYuWCHiBIS0PzT+Pcbexp4UsssH0s6J7
tvjoQ5cMkalIg/i3U1UNBFROhnF2+RjBSuvlhz9c8z8tVh0qtzGikJdu+kg8QEmi
6sUVwD0pmDgDHWbuo5vul45qQmENnndtUUYNjhfG/gRJn0STNpq3YAufwJahvF0h
KnstCCXKJ7F0d8k5fO/jFf5MURgx3hUXcYNG29dUM9Jz6TNNxJrDsJRJzIe/gnbt
M+15hylevXjOLKHzWDbky+GRdAHXg6oDv+/MFptTcn1hR1DjWV8sXhjIg6gb5xn5
bFdCiPa/QpvsyfMCkUPXYbhMa2t6BOl5DbIJ9zyakY8FX+fVpZMLRHfNy6P5Lcav
JucfcuwSc3koqJDB5F3gDJhiVEhEW4tyccUFD965eAKAoCzJdG0BbR+b4r9E169i
H/sw1FmRr7eDggpM1J27d9oRRHy4l3RaBm13abEKVtdc1bpr98QfhoJZqLykjMCJ
UGQhffpmwA1F9CKMaYq4JBuhTOwXcC950mz/bK13CpwmMF7jhNIIEWFPqC3LmDAv
+W/6jQHOGkrVO0oXUDzkVk7c9g8Va8ocBx7ciqxxKdubgr4uSVg2y98zrcBNWq0b
4jayMjoXJuvqB8GA1/TzWjQoyQQ1/lrqZhv4PzlVN9KwooPj+71971d1enwCFU6j
PuHbx5yMR1YSzkxHdUHW8kYWxrDbt5l67p8Q63tQ30eWYjLl3d+HUnLqIQFVJ1Vk
TobrfncaS3wThMN9IZpGrUjTWVnW3SZDmNNEOEYvFmufOZ9X6jBYL9IIQqhC2FUR
quXnDfTQxHXQzJOx5iRTEDaAMR8HUL/beHU1FPYLOmnx3WH9T1porOy0jeYiZYTV
epl+F/N0Uds7/nY6iOuSEcWC1wSqEf1BUGNffd02JXUyUgUdPDTi79EAdtoHLWzr
QpTvgJ2IH00dszYOsfDWKsbS9vaoP/UWBOHg/6J6oLNBTQpauUSW0sWH8aB7FOY+
8F0/9Sq53mtF3rHBl587Mbj0GImJo1zEwmgINerlCpvcX+V2M1j6CW8I0Ye0x3ap
JJe38tOztBw5xOrt62VV6wvue7+0a+iUkYfx0f0VTENumybW4jJLv29HwpJokuWU
b62tD9+sr02AlRqE7JT61W6xadsdxiLnGvYh5ig9zz+tT98rhhbUshOQUBbpDFZR
QBcnGIkjBblBGAl5Vdaz3A8jMWIXSK2W7iP0T8TMk1NILEQGhUqaEkXu6NaxGUCi
gug/WyDtHB7a0z8nYvsjlkwMuGzn95zJrfScwBLI32CM+y3cS/XNV6s5GjQH4Pnp
GflFcZA8nVX7LrXtlEUY0aiT1iNFtXwz+lVXsRyhagnVGiryQ0qcJOx1qBOS4zX4
cxTrLIlKBYOlfOfKPQJp9a4XwUXjd4F7VQRPMMyW22+9gmUdI8K0RKD/vbde4jE7
jmihF7ASycgKKASUzqyRnjYj7rvG9ZdA6ZXA64SUiZ6NUcHJ6mxLSZrJx8ked8dF
4JqrkC6o1WRXkFiZ7SL+j23aZ1hmtIADCfkJ/4WF/9rRLsIHtlp9E3aRads9iiI4
F0Nt+4ECCVUq8UbWDI2uuPjiKOdeMN/phcRzI6LimWPLJXOXy9ZC/fddxsP/dWHq
jgkK5OxtkXSoftpJmwowQLYf1UB4UBKwv1nMpNaN1FhxliWb+IhAvekMheHFEHc0
rvk3ultmlKvtWzux3gGyNCNPau7H2OFpSXGpq5beXQ1E5vsRi+xihGLuGGWPKnWS
Vr90/pKqWsOQva3txi2Txc4nwsKxyEc6ATBCSDSdZGDLvbJIXWjpHmXFdo+9an3g
vzwmP3BNPbW/S5foe8ATC378UO43pkswwb8JKlcWH3ZAiOG+KjXEF7W8BbMxytM8
DVXTZDkEqwPU+82QRaBrdAvkzADNrVPo+KNp5F44wsPyUxJMM+Z3pKNwrI6kFqSf
srfcKEFOTHFTDbxKNpXclaZ9XtV77cx0OJXtSBDnCVaiTt8s1hecCVIgqEVgEqMC
+slUpIZYtC9lm33DydCCTzrN85jBsXvrV/kFCRzEzn3a7mCU/c9sTY5P2As2JyWg
g/igsnUemuvXiqimnEz2IQ+4PtMTvdBDsl2FEqMHGi2o8DMO+7NYInwPp6V7FgNt
7ipvH3HWx7ohd90q+RbJRQbZ/5ObAL94mJokGJ7PAtNgI+gD5d77UsKu5nt13XIY
F0rPySkf0QD8KDYluqUGbIwd3i1yegw4e1wvaoV+ck1A1EwMaNpuU8iWEOv3u1dD
ApMaH0fNv3i7VWERSmAQYvPD5hYE2LYC0H2H9Fx70llJq2aZJuLIzfarLXzoWSCl
Yt3qIka5VKUF//NnZQje8EA4NFkVB6QxQh9+FYkWNmSjl0RrWTFIYhBM0VtEirdU
kXsyK0maMzWKb5OJRC0Hp8CqQUKJHRGnseZFJcEhQWH34VvBNCEnhDTD13CCLkRl
UOUd4fBn2t6xH9IStROdha/pPcZH0xcsthwu6uE824vXvklB6Isy+AlMBYyJl1Zk
cYKyRJ1u3+NTwozARnGEQ9sSdC7PslYskZ6a1f0sQc8KHtYPuH4ndZ3bFKsYCgUk
hkQh81nxYkHJiRqZU8mexNkHX0u3ksLR4ge6Ax0h5PkyPvneOhBvYSjwbd0o7Eaw
dU+cyAjpRSpIiJQmaLVw+z1F3oXDn+0Jw4/Y67djj2lQsjod3LiKInwlff6gGIpC
A1XHFyBUfxOu5bJoXk9ahDeciVM9Bz0SQYcAf4PgPnIT5+gedPSjfhtnfAGYOitI
d0ZRx3seTUPI4GN27VIGMI+6Tlzf4mshaXDzUXIK7i7eS8fC8itxGVpOolUNrlsb
XyYUmSvHrgWMtdQqqvZZGm9y1KYNJG7xiPz9UbJkWRm8a+xxB0OwPMn/XkFfPjGH
P0A02Wq8/WoIcK4lkRnwDmNXFRQq7uTFAwkD0H2RoXXvOsfeTXR8pH80b3TciiDs
Fj6D25yLK3XxlgE+acB8RYu3dMane0BYINLNBNVvkL4ElqxDyjwnqx6gMVB9loWw
PI4qf/i3oBYlB43+p72k1y/9ILC6OHjTdgcLHLBMcHPsvky49eZWcAAvSL5PwstQ
iYaVIQWBcMGn7ARFJ8jSfThx/bNJt0pRIzFw/vnVDm9uwNQPqffAmrt31yQBzV9K
2HywAHFUNRn8ukOYWHgSQsubCeeonmJFsv/lf00DQSxfgClwrzUN62asxMq98xEQ
3i9awOWunWHIDEF4igKgYAmBjTPR+ZXp3pTto0E2IEJoluQdnuwYPtJySymXKoyB
o3fQM2WUysCs1FngC0pfkAaFAT+0tt3Blo2mLgxCzmYBb2rWOhYQPCFdSMEcxmGa
8v8kp2QKyyN9gjYNWEED7QibR7yOXneIkbSFsvPYSTyaF+Ejx9MUYm/U0nBTiJTd
Y0iPoFd89ddXhUiMSZiR3vNwnwEA0JTHj8mIHIn3zsm7cRgN0QJThx5V/xvksdni
aYfnr/vunmWQ0JHF3qTGE1cePFUQf80dg0XHw81T5o856xZHF88gXbMzPU3t/BgM
OM+tyNeBqJBJjx/KL8Yeub5rvQ/1MWRZnpWCWo7IrtBm51O7O49lZ3FTeXyEmUTh
809ePO/3+8JqA8KjG2HT0NMjKL7AlyCW+hI1BgiPkVP3++Ewj/E2vOkYsNGZOntx
4kb7VKMO6xaxVt0LeAASL36jFNVl+DsWFt/AhSuorPPsgOs6R+B6FGbftzm3ku73
Ch03d/6fvb4dWtjQaw8dDN8/BPw1ByPrAZ5sahtGJscZuG94Fdzub9BDWfvlY0Pj
nQLvIspy6UTz6CEZC5/zmzzy08Epfis0+Q0vZ9z+E24//GFRDgpYkmkBeNnFZyp4
We7OpBdcccIoxg8qYSovZHY4Ede5WN+yr3BTCl1R13X2DQcbKL9Z2WU/NcPS0UeH
Xfu1f29yzx0mN3AQGH+gTLrYbotdISYbVFBtk0jrOWfIQKRj3QcCxwjh4TwtcXD3
x+2et1F3BdnvE4X6Xx6PIvd3Y5/3PFfuIgEpodozFNoVMh0qEj9JcqR/7s+UKiL2
NlAsoOpkL/oCIvsKDD5i8fHFXh9so8ankcXpzI8kbvE5VvoBTMIiki3HRyMupkSg
eVBfv99SWaHlwgdguhCKN5P2cdRcIhnL0//VGQFBtVN6C2ovdb/FiYAURk1n57gS
xgYHyGehkfuzd1NjsljkIRzzj/3rl3iwKUq9MVqjGdaswkFWF8DbWt1ILIUejrbt
jWF+pKiTqD48tbvSOOLuuONL2nGIkOKjbQXwR20DeOqgYxY9U6M7Ja4WI+PH7N7U
ULDeNHD44h2ajDD5zrPSeMktlZRwKGW0N+x8pXNSn8Cg16anvrj/Nh7OUZpH7gcl
8sg/olsOQBuLRgpRMeUfxrKykqCqF5Ql2amZ0QW9SUbwXNj2uQrwLnffd8KI9Z3r
d+AVpM0wm0HMv9gLmSqPR6hu3UyhTV2BAUgTeE7eNiIlvXdO1KM//z5DNaCbEeJC
Q9pVhUJcFUknd+yYfzwsZL4MpGqJfQNBmUIogqduPjvGa8qwnJ0rc04Cf/EsFvof
/iA9UxM9kbJQinGE88tTjatIj9cDU5CKk7bDWfNXExTGbWcow1i0pYxV57+FC/8e
1Pmd22c2TtCi3YEes0ikMATCa6CSmku5Rxwpa9naobDT7gsYuLyqCf5xfbORALbh
v6HpCPuZ6Cxn8CGb4xk8qtaYy65B30UwRrdsyB/Li2kEmkd0qwuiyJvIZrutNaKP
wh9chBn5qXAWFzSmgQ6fZM5e7dBoNf4gS82x2cQsUbTk3KzK0WkAoAOxUjxG65rC
nikllfV23nN8Zhd2m/3iOjDdMskvfbSxl6Jp2DSLJF4Y8boMHcbmfZnD7Bio88Pc
bkSlyHtBkVBf91vFqyHsl8F5Rs3GNKz+/BpGgCNu5tjNzXgzbSHbfYKid4IsvfXl
lHIhXhoFLZacBvUsfFu37fKf6GkEKDRCrytLlb+K1cgb6YXtREXpr6FqVTGShr5S
WTpEhZEPzvo9oQFmZmrhXCxS+itwms2wmbJ8RRCs++6bhuEtdTIXGYQDP3GgNLnK
5WSZPGLGeSBYWAlAFDbZffKQ/DZdn3UMwKh5vJBsJyqUGZ4F68yGxJqKntPzKY/a
AHDiNktrI3KQkSaIQCgLRHYOvuEeraZNR+nFMf7vvoMCIWzWymLWJNA6AWCPjX9i
r8HrFGTfyMmqpRn9oKvxn445MXrboVSZCwOdn+wNgn2aJstaN37ivuZdvwIlP2t+
Y7FgwJeCa0EXXlghqIHxvKbIFOwkg2CEjgHdPkFRkxask6/NkGzg1zhR+ykS1HTc
WEot9dEI5iUbksTjY+UvEVnJyVnkoydq1f+KNevBr3OZD9fkok1fbch+Jb3Rs+Od
hP06pnka0IrnmXrBvBvwvTOtlnsdZfN4sowJ09C8yEUKlBwWFfSdKqWI9CYvKYu8
fxhKUFrUcD/0VLrsXoqFYkPINr7KsUU7eLU2r55DZRFvyf2jveMV486KWzGdK3vv
dL7fGuJ0noR1RXpEZbCq+SKrLSeWVWYVRzgZrf+5OSQ8NqEr3B8jITfXgknZJeUS
RGB+T9FdqP5xUuBx4VlAZXA3v0kGEVyj9m/yZgNd81MJb3on0jFSrfUbRQKd5ypt
JvBzr2fzKyjq3Fqy7edzBZ4d2LL+l3hJ4IwqO2v08KAm8JPq9xclArVJ0lDoifOU
YxrD+O7axj3grD4ssZRmsEJHJby6HT3DQcP9v2XUVHPGpKXEYcsCOWymaqXTN/jX
j7thrXSsw7jHXAa19+p3fogcwCTLdD82fFHH3hIeE8SwdLDQfSt+4kAsjffYn/hm
DlFi6R1ija9fo4y3I85TOgLdsymj5J1ExGgbMqVQOGTt+PApzRKLsYfy+hTOqjum
PuTLrQF0MFYAkNO/XveiI9PDoAPror7nQvEaQIjbn986gdZNAP8Gn75hD7VQCCQh
STXZV1IJwxnPo8IxANKxwsxGu2XWo1gHbocuq/WUZ/TeniYnRqso4ssajLUdrmIs
z2OLXbGe8Cj3brN9atGlZ7685K44m30nB39q75M0I82ESLH+TBYWa4gVWs4xBJgc
c4IHGM8hT8v24tNTfoJvDvag0ISLhMGpHJXMTvjboAWII2FmqxvSRs+ocF3dUSBN
1MBnaQUUUC2PnSlD9PMeI7DEcU+WC8MZD5Dbjno+MvhrGIm4Sd2nMQzh0IzOCFkY
vtcU3N3rWdIZxPqaf7B7OYIdX0TJ7gUjvlnJ8TRfhyN/FDxfxR/Rw2tKmAFJjF5t
+IL8vFoyRrLfsKKxUeyBzsugJwWRwWlSB+JIWCmffIvGlnQZZQS40ByN/PUwcdJZ
N5EO5X21aZjcEbOLqm9mwtVgjgjcuV6YrjHTl++EJeuiB08QgimLo9Rn4sdeKLUb
CJLYUlMwU9/2xirMU9ZBsxozMzF7hDxQeRY+Y/FXg/TDWr/ycG/31h+c81Fs93bJ
YqCZqjuEJxnIrzukfv7GhVGRW0UtWPNh9CoiPxkiXFtY2+nyZzS1+xUJpGE2618w
bITXZw3ePcZx/2joikMfMlb3agOYmZutbo4LCAX9O/VRKjBfF7bDMBaJ+7uFdoIC
GKuyIh6pw3JwYg3xQfwDcs3EJeGy9phs8YAa27gXJyAyoRz+8HZBwR0FpCH4MXRc
umW5rbJU+5XbBbC5QgtMsZjJIgZtE++edT30PQR/3VsrEDnxmRro8bq3+n38XDWg
bp5ogLy5mJD0rC2g7gQNIM7fAnU4eecLoE2vp0BkRuTb20HjJ7gRrm0a2UJugQ1C
OF287C/fY6ha6xzxQdI7aFvsA3W4uBmY/nod95+o4azcE/TLeqjw7xE8ExvvaP3j
masR/uaRUnzf6O9l614U0bc4kNJCNQl2v8aFmDpH/vErw0ksEY7zzKJDQe8xOEwH
7vvPBktqiphHW1Swikedou0cOqDvqM7vJxJtQeple0ejHTuxJTZy1ktYYh1OdYJc
qHOGrARe+VNKczLuLD4OrKAqdxnD+LWqfD7PjjkYBkgAASbTEgYP24quAG7eHPln
PZvew2e8BBN3b5vg9qwvTPEaJa5U3w93KfiiUOo2LKg62ZxTrZpFTVVAc9J+CyxY
T8fre75IOFVqt0XwURXf+EqrfEiYrIgtn+BDFXbBK9r9RkC1ZcK9sVuHIGNM0K6X
VBKGIgL5NZVU+iCiWI4Hn5ZpPboaUzclNLfGiECJeuHIZACM6+hNtXlFO6gJGY1o
18lTt6puK1nfcYMLG8u9QTcdBtSWJK2POYADsCk40ldkUqrtWVKGRD1BqFHxnInd
zLgM73sp0GfYq8cZLuoCrR7ymq1mt17DKd8d56aoMoHmlDEvKFZOSIxGqvj6s+NY
G6YaS2EKqHyW8NOpLdktHePJmzeyh7RWS4OObHnTVcHn8vtIhORXPuyZrz/dRB3J
bk51WJY9L8DXWI5iNgu1tQGenRhqyFDfsBOX1c6V+H3X9xGhUk6DqKu42iPXt4Jz
loYFrvTrtOs1HB5XQk8LeojwSg11ld3dCgpLwejYYA0gWf2/d9a7vrCon5SFMNsO
x2kZAMQ4V8A9+5UblL1k1ZHNX5s+fiEBTebi3ECV3zpLQHPOIxUUoux6n7Qh0IBN
CWdKZl80P6HvFFfTBnvAw7cuJsxVKnvxxg8eHwAJYtpguhfuTKFvwPopdyb4C1rU
hcG3iAJN7/S/xszA7j2YGHKzphyvtfghQr/JrPFwGJ92fflDxdYrzPVsjR6P3cXu
8N7Wxie16VlAAYEgBK9k43Lkq5X78lpvim07rR+j2qjIlQ+jYWLV88tU4S2NYHnD
sD7bFt2XKU8UrCcw9/3vPPVbzTD7wc0AhkK+tZiZoRpOBrsy93iqe2vnIzuAeyDy
Co/9BoUo4KGXc6x111sLOAZtPyAlvtOI2EzxKX/MQiYS3wXX3zhHo2/3X99TRI1C
rL/rfkrmfng4ihl93/t/9kuCh9TYhwOgn9FKY5N7TaQ73oP3sobbFaXFlfdUKInf
a6t67tGUcIK/6aX7SYAcYaOX8Or7OnrjbmqieZnGcmLBbCPOfV2b6B9PoB+RDnpO
0tGs2NI77/We1Sj9GhfVYKet1pX0pef93HcWoeUk3h8oRw4IbtZSCOOfrUXm9VLB
hluj+bF+a4GQZuLg2lJsnslkkZrfECez8Kk9J05mrzzgjE5gB0aPVqavPKahk8lQ
TrqFCZbRlQsqgCTzqLg/GJoRpHazMcqbW4yjey+N3tFbgYF0+9YnDg0IsGWejgte
tqAHv28tmbrAxQ/e7X4u4I60NxSlbr1qCEXGA6bXnaoH3idnl+mW5AoOnWABSAjl
rmrkFtRiao/IDL5VjZ8N+FPJPneCJoL4ascux0BoJ4nNsqkUqbyx552r+jcMtI0h
oyxrq4XhGTLy4okvd9xUtOK/p8aE+BORmq0KP6a/NDrxTNde5xyFfEOP2qbxJNIV
QSTcWpkqu4CVJqCnjYsGqUA0d+ElqyEbIV61rJ2F6+bFuW3b2WaCCNYk665T4pFu
YtduZMZw+/83EpuQDzU459dXEQwUkuCjaZdYS27tshEX/lN56Zplj7qstpEqyw3Q
9OK3Lgd8oWJ7fer4rZiDLJcL8rm40BEZLNOMuTUlyT2g0fnp7v0bpb70uCpVr7PZ
oa+agySri5efkoaZtFZ0NZWg+FoAx5aHp7sABmzzmdQ/jggGwdcEFjttWPDYMpfm
2B7AbrsMm/azEhmUW8fGdaxAyoyqhunkFi9+a6rfEWjwOYDU1JK5UMAAc/NhncgK
USrmyXS2xb4FxBozK4ftAiY85t9Zfd9x1kO2J1sXEdjC4JWr0lQJ5xsoeFvrnxUR
ryiXAioHRrQ0kawtUYBRYLx2q9ZqGAoTESz/bFFJboiFR7Lb5iKx/m2gH2DR0O0/
one0gxYaSDKtE8ln1/yXLCZCGBSXTUwlgoEpBfOQBkHtk2YcBGS69vfxydYhJ4HW
m4kWgODzycS4J5PwRWKuhOBOZYRgoHQCq3/I2sAK1QM8G+gtV5QF9S1QjKf/QPOK
k8WlzoSKCZJAguw7RvoYu0zDbXfYIzZwPC5oEZ9eH8t5lriNCpyJ8Glbtuf4NFWJ
6yLSH/4nGYBVJ0dgvCA26d0SZGy9IiXmWOvuJ9+avX5d87XyWTYlShRqHBZMbhAH
9IGIcIlEd7DUld4Wz4TjtiiczXzTmNR4o191vcwiYwRCc+d3KaNhvqlSG6hw4BQd
us/HPuiiFBD4nBAt6QougR+e70e94knjGOuiwv5HL75CADPkn16xD6e3u/irPdQz
32FXrGhHb95OzGklZSbPmk5VJTX6wS6t1yhVMid1c7jF8kFqFrzzPGF3VPBPZSyI
0yBZVR1If393uhFnqjEmsmXNLa9Sj0WV5juYU5lpR5lDagz3jWu7u6IoIWls2Jv+
jnDuCy8WYETkQJ+WWMhzlQwGUg8/bG4hfsYWdOEx0A4fga0wVyfKk7VDmDmkvw30
xxvqQSdvn3g9///yMKe2tgf8QsV+Dh3ln2SoGPcnsXtJpdVzluzdE2t/0JS/BNDO
4dkoeaWsZL/L797XHtsyolZkELjEr3wb1cRSJkAya+L/VjBiqi8wxgH6G8PbMO4Y
hUTrZNQ0eVELUtcWoCyRN6iU+QjptpOZYsbBIRoQLNk33OmuD7dlO1bb7IyU/cLa
TvrHnlbkSprsai/1lJKYLZqRkRMXAH0g8x6jzwR04PjdrtNZcPnXXszkKPkJmQOJ
H7lIXRXl/SUz1+C6Ogw306TqWm0jYfV3Fww37zBFdpCOIJq8qR8XkzS2ioPSc92i
tnNhGhkhgDj/Fn7Wi4krYIOM5KHoJSkWxlBkTcgC+JphUPdiaTHuvl5ugEq5VevV
LM5QHW3TeSSOfKq8M+2cwiMlJNExudRCmoMig2brXL1rxIyLuhvJdFRWa5Ar2aZ/
Wh6RCVNlULhxHLJH/xsAy42/hJMANeqfrgz9stXtBosVZNtfJDQdY7ONTNTFExiE
IHV7dVLheuKzYxu+GBA6YkaPRYIwkQnf8Ep8OVhCgFWOdwDBb+dTB8pfOb24d7QW
N9N90HulYxmEC2bXA57eGGPiALBdUM7cvQ4GLxhrlhnFQChN0j3Hl84mfJlBCezG
eBq2pVHZmJwFBqCLOhWjXw9DS6JlCw6wDoHEvr4xyt+s3cAvi2zNGwrzv/3hoq/X
Dzzx894sCayxr+arckvmmWp4OvLYtmlRzjDd2OEUp4L1298efdl+NpAwgVDl/gow
FyX3N08HQ0gfiOPOaW+hHt0WF5YEqLeg+f87LWJEhJoqkGQfOE0ko/6gicinLLvy
NXublkPpUz72J+ddmIefifx7qKqUYLOPexFu+Sei9kLVYU6hzI2IlrWb8hnIO8NN
zL8so//AI8CUHwtUd0vqVQ0+BmtD0SqyqPqNx6Jx6OSplVkJ383DRg2ynCrfMmVs
mO/I2WvqM8Z35URL5ZnIiioLHciQUH5HXmw/RMFhE+E+co6p7QVPbicR0s5/xmoJ
jWkH+cXXLcm6/8bENRHhAXQkh4vhhNnDgY9Jx+KcwHNtTy2TF7AuHXkxUPLC9dy0
r81nkswrue18gKcS8B2FD6ZJs+gSiT6h1tr+T/cC+kUNp63BKmXevP6dPx9q1fU7
mcVI5+UEdEHAhuoBGPUxXi3GRzixVXp3Wr8XOWdNsPFZkf7lf80i0RmPMJ/+eaKe
grvwefJbd8vT4QdkDBc6FqyAK4lMqAMzU6DGP4miLEsn8IBMr5R8F8BBSHJsecQV
SWX+GJ4zZd8QWhYx8kUfpFENJQBbiUgIRB6zLLN2qmdSeZMdT4HuNI8UlMpkqVfk
yAMraGzuQPFc1Twp/I3m9zwCIdqJIEEBxPdfYH7HRIn/wE2ER8oQMNrPNVMpPyfy
KjSAkYLtxM7Zl1/JSHjivREgGUokJ02qTdn+kkiFXNy8zLYwUWLU5maA9MTUTG2J
rBFC6EFp/v91rf0dByTRfr9DOhCwdFtOzV2W0mhm9YyubHHEdxGy2j3t2LK5zOTl
E0VeIOO/yOYby1Yt2lGaDwneZM9Zy/q4dB0cM1D1DIQdSuxlJr3j21hJyJ25pSXZ
XGF2BWTIK0bwYsJuUjj8uhm7D0t5xYlw0I3cKZfjeT07TXE0FISSH29CrQbzzijQ
mSdsE9OzQyIg6+Vu9owZxBERuLCwlOxfX+i7HcZ6UsmAVa8GbTc681vLij7otWy9
hAqf5q43q+TwO5pV/7lOM/GNVJUkxvC2fPQJi+qp+bDGwzWT5f1GoZKVAHpn4Dap
H5sr2dr8e/agVwU+UONQpIUDv7azZifNEGPXGOqQAGgeeV1FzPKoNXShkGLjpqsz
bfbuF0YxmiK0AH3zASLrFhxF66sZZt1lATASDxqmb34yUyEf2GZZdTSRpIhtdG+J
5+Bzmmq2Q0TekyXbFYcxSuz27RnhFIqwVUjNMpavmhY9Jsu3QSnI9rVvRaUx2JTR
OtkhDsGEGAGNNKta9WqnQjeFJK3oYGAirHH/hJ4m/zoyxQQr/D36qduusI4oAtBy
HPTZOLEjaYgztikjAN6CBQbn6jcjOEnGYvnufDBvu8GqDOKy4nVB1YF2BzGdjJbx
hhfLixss8y1ZXKj9Qf4y5+RdwMOLFTSyfrd/nOkvIs6Jk7884AxD4Fbaf7CVEB7G
TDVB5uC9m0PDCYQe4lvAIVXU/WJNW3BBSsegvgaNipruudPShNgou8CUKYq17eRq
uck/tGkLMnl7DTtbau1zhOJukkd5F0XIi/mSoj9Rzv61siEdzqsjFRFDxZ0gueCS
c6cMgCrZ9kVhN3ZAvh2/vq6RK9nVGK7NXIWnS5vQToDsEGTox2mPcdOzhGwH8rFx
Nz1j2PrNAQEdQym7dCnhnztPvwX9Jb+g+SosvYOijTwjiISQLllDs697G3N8TCBX
YwV02VooqJ/zWbIm8JpLXL8vkGOgPI3Kvkbn+R1XMAiIGnKaCBNmeJfqf1wztoLY
ilWkBnq8GIWcX8hYZaz5ROYXTPX55bHjwLyQ1CGtiLKb4s2nLJCKQJfRpwBI2N9D
TqWHcDOLbwFf66mkvf77IzR7cM7dXqcAFibttqMkzmvP9747Bz5v/qU6DBRgiY2z
iFfKn+4UUeQhNawLgs64Fhio9azjrJwJtuSWwUriOzdaYKLbco5OFFZl8djlROh4
LC4ceWM8gRZyfqzm6KHqkCdJnzZON9u5HvcAUPh0pkPK/P0jot99cW75JmtCKm4S
kO7bUtvKvyueBrH8DOA3Vksry3VTMKpbyXh3SqX/eUd+s0s4AUYM2VSlnHQzvu3x
NffYVdUSE2MRwl2ORyJabc+oeXmqlxnYwDNL3Pr26Ha6xalBNB8BZauu72JPvPHg
cqLTB11vmZ6/ODRQvhxEOJEyYBTaKZVShyxiZH5tZGwrLVn9riUJqlwvHVSpkcyk
LtVYPn/S0BO/Dp4Ikg8I2TdcAdfU/kV3yBSy6Jp9CAKYk8e3XN4OsSSWRKat6RzF
q6UMRrsZjUQ2ZrTP2bLy2LtwCQm1ActzFcP7JCKu5FTS3ICun4cgXHUySemmvvny
8G5oXtSpQrGvRQSRz96UIQFeZ+JkYf4UFDlzsCgj2qK+xvTUnzGtH6MaQpXCsOUP
L7N1roJ+JiLz7CRbHKWsCLVNVAPM7eqoz+twJq8bIh9TAYO7/N1gga/5Co5Df3Q3
0CEMLzwEe96klE/S3mOqLzCHEnTrwVS3YWObtWACgXtDmKN+4/jHefO/hqKEr+sk
IcJPrmnnSPIkLxfGCmp3McpFss1IF9X/Zu30CJkT8D5oG+alfRVLlju5nI2dLe+K
ogQBs3NhXefJKoixSWfMT4jcSJLO1FS+YZOwxlV46XNpGPWftuk1VAgpEDCpHjs+
Lk9+czfEjaldaomdp3/u4NfMY57s/Ges1JujKBvTI4Wp7N4WFyb8cdz35cxN3ypX
j0yCMe4YfWXk60fCjlHqN/fr2qB7URmGSyhI6vGBJOMW6HOEfRXiNFkKtsPL1fke
UMn4e7VTuKb8zM7CfpzbQwlz5jrrQOxi4eUWlc579m4s/+6THtjLLH2IMxrQkcLO
Tpfxyih61BCigZXgcioleriL4hCvFi435O0XknIs4jU37dtN5Ssu+5EU9+tFGahD
oeM0L7bh+dxGByQjBhcvpPp9WII6E2VRjtah+P1eAeP9hqZqxOr4zk7hZtQ3Z7v4
4ngiWcnOfknxVHUp5lJwpUBWx/M3u0Qfmb/amejGEKJD+DmhbLyeUkRjbAQYcLY3
oCwhdT1bCfb0+Mwn4hjz20C1TtXIouE4skpTu7/V54YmYNcpXMD4K+iErQUr9wLm
rUmetF9LEjCk7ueRa2kPKa+VVMKkgzOEjoj4PeBdbGQHVeQjvSR4z9zy45ihgyzA
bc1OZ2cweNbsbYNHhvktbehrhZHW7UgDJtprnDeUj4NtLqapjKrVvZg13RoCO3SP
NMYRKFxVajpeC38kXabyHAin8pzljiSRg9SgE9+vFuwOeldUvsy0Rfr0t3AcCkgu
ZjI00lQHeqShwqiQSRLht1IdmEYvzYRSpKAgl4fk/eK6W61oF46Mz2aqT50J98SW
gwtItp3CWokNLzAJtkoH+8qZ8cx+9rhg/uMLsJXUFkjINUzOZU7B5ehjiJ5dAQfu
Ox2ZaxElOx2noRDT+bOhye1fPQ2bu7386Ncum0MKA51mQGOOHXHqRkMwipVzFIWR
BAbAPCLPHTE5Wb8I0pS8HAZgHXSdYj8hmmlUkqGLdGs14d+sGHVFxrDal9H3Oajj
O2wNNOsR9TLu+iW+NA7p7othq/qTt7smGY5y4LepAHl+ZXoP2QdIpCDenVAcbRJQ
OmgJ6IgaXaCxMzGr4VxB0jbsVVeHC+pRCd+nuwHWFHZcw1KNKKueKNIwVs6cfXcO
FacPGPz/3uxC6ELZyxxh+7+v81DOUBRh3cPHFkVSDJc/xfK38pGb04Go15nqpRU+
+roYJ/VgPySheTbh+oU4WJBn+Tm/uLBo17e+anxp/CzS77U6WIVkompoJbPNWZwI
Q3/yPejOzlEkL2ChtN+VgY/Kc5jhvIAvbmy5/S8nYR5CqedpZc+7p1mZ3+ygRQfU
wGbe2A9+3J8TFIziOq5adFcqokhd+we4Ly/zH2mB7FVo/vPkkjEHEHNZIw2FgyvS
HE+Z81vXG6eRYDlKrWbAJkEBgiYNgv9h083pG7b/dTJgkE5kInSP3CbvnhR94Ka/
n3O7fcvUD7XChUcASdoKNAp+4VSDFHsLFp2xCbdrLd0VA1IekkWNcXJpAzNeMWvY
JGqrxBxbhcFktfJu75mpNMdzPrOFvkCdFexGyppvS1M=
`pragma protect end_protected
