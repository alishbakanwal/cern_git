// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:38 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
eUe5zZsLBu+fuSzxibP4kgyz1p3UWgy1Zjb0ISwOqVtaTYjOv0pOFItP6wRS5uD3
Kd2LHhV7B7X05mxM1tvyXDK0wyzFPHKzqvs8qhJlq7GHUaDa1Rff8a3hB4TrhV+s
U1CbY2X0Sl0rEPHobqIPfuEd3ZKFldGGZg8Qwfrgyzs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8800)
E7jYVKjwNujEaZ4pJQ5b4Fi2pUCUjf46DLpwK6/tsIxCoi+2ZslPOgxgmPho7Mff
GOGrmvrWAS/p/skxoxTvlvdzzYQpymFox90ApYIvmrvXeYPv4QcBxlzJItcnJkVe
ja0Lr+2GT9B9xJoso/L3/fndm773nnHq0x76bp1CYYj1H/6fFaKw4vHejEhfpkaI
VaVlsOsKSYeHC4bILCk7DTKoFgI7JAKBUTzTM+EcgG/AciYc2L6IoXJZXNYfnv5C
IqTtRml4hEiF5typUgWy6fuPoct6P81WBpdRS08bpLeJ9GYGWD62feVD2jy/5KSj
GxyJQvrnw2txOmoGz4/7ed5+PP6NNVoTIJkvhEQ+zjQ7h8LB8f6r878EmvEfV8GX
C4g31L1tRj5oa0hGtCizp1UCbtLczeHwSLo7AOeneP6vzxTspaGeTg7/kg01tWaN
YQQUBuctZmtaFUfbMd7MLrqhyUOogZrELb1Gl3YTwNL5ehdnF+HDhDd+v/GNlcwb
yQESXyNCHOYx0iVCOkchdzQFdy120YOL6h23sXBV//X2tRdpMS2PlfR/PwAf4H+z
d8VX8vaYAA180MzxeqQ/S1ByGcJ6OzJrTKXQDaEtOve6jYQGLR+j2Wszr87cz0z0
3DzrkViVGWwuHSRD5jufUjhDj5MGXuYhHBi/r4YDUc9yPTs1LkE3gdy1c0x905PT
Vit4P1AO2Bpioeglc9yTIo2CoRRcvheRluxvCOit49KAwAuFsUVboxCuOzDWHPWS
rlEGtKbrHMvtJrXKdReROA9IZVGu3i14xRFsaIOB+Hpzya6Cj/K0WOmQDoG0bhuh
YiPFtQFjfuXfUSJU6Dsnkf1joA2IFXCwcNsehUQSuVOJBkgMqYlnZfm7kfeo7A+B
BG4zilMabeBNB8itKbmsI6QkroS4G2Mus9iRgp4IY47gvKZfz3Avn0if82jf8IYI
en/KnnzUoZG9gz3Q5370TY4PL1EMss7R2HfX5WCZ6TZk1zimikmD0rd3wdIUI4st
GC5894b0TK26u0DNAmvyFwkOkZNdVA0fzODkHOR/E3DoYAGdmslgcj+VayEpE0Lu
obXGoVacjMtt/6uwJsnSuaLNmesUILCf5JL91/1LQB5dyAMTFpik+hB+koqvABQX
JnEV2yUkyNRSspVXGD04LYK7mP9LuoK5tylgcDCEyzK2i2n+6wr4XQu5X3nI58wr
PQJf11uSBjkvzTLEqC7LMPqPvH3Enqf3+R3+HRIkfIy1KV5fWV8HZ6QEiBoEh4O/
TXRpmh6jdxKQ18mEwSvp38nYBc33dMOU+oKI+ms5SuBPszejjEXCHCXkb4csjM26
rMokZS2zM06u3stmhRBs5+ZvoMIUxYvsNHZLFdFUJRaRB6oMSUCwhsjaun1tXjYq
itqj2RHdaueJM6QGFszuj/89rajWnOlXlFIv0U+MV5epi9K9m7CscjTpqsJ3WJYA
XPR0JJAYWlyJCoXq/xTNu+zooybM0em/NWqmizqQ4I2H3FrVTRsygCTlwl0JVKn6
Sp35d3PYFGK8jPxGOZ1WyBEw/YU0K/vQEB/FW6HvO8LWc+x4puLLw0ZcMcUEHHSb
eqpB8n6i7JMnf7K5z2n72Admc+MHAHWolCJZGM3aH1KrW00RYrgsLe99UAShnfqC
8sO2jfjK2NRKXMQzYNODdgAOUiBF8AYxcgXRWGAhkggdGdq7gKMuaFV07yD1/ag+
6phx1IornhUw/ig4zTwe32IZRufHi9vUxPppRec3L1iK0FpU9uOwuAWfZLeBbPvP
IVG8gBizq+LaGj7GFGt3HTyk3kLb3zrhed/nhhYFy2gObAdLdPnW8wFwG16N2/VN
5zoCHqSmWyZbtAY+oYFJCprPoxbj47M9N8R1lZGz52KFfJU1wnMNeMi95FI82RPi
y4DrsicCuMBPj0I9MoqrVTslInbdsnzJut0BIB+f7FdHMmIAssWKU49LQRJlC5N0
VJxrUewYIh+iMVkDU6q1gJAH13Ctb3MrSnU1QC9Y8F/f1D+sET+EMMKTrnwSFYGh
PrGBxAESjPdrsUCXhyzM12oXCKtA6p4MPj/Nx2VLXGgifvj0A9k9cfWOoe1K7FLc
FZzbzIg4vx1uSp7yRG9zgMbF/KpykvREFJSWALED5uiw+yUpsKzh/8d72T5GpIYy
hnzEQGJXBN55BU0VjEfBvr0Xi2igDRTXPEsdgQljywEqCLzQnahshfhAPBntHsE9
TdRVBZo6A59bSfHgxDf8G8ievnn5tFDrgWywjQBht3GU5nNaqTOeJAdemDV1gMBI
OM0/Ppxx6gPKQeC4nNmhGIpRtgdCnZd3PQ8B7g4T/8FlPtxJijfQtELN20XV0rca
hAvGDKgrd3S3a6M3geU9baBPyXlHeSJUjGyLjl95n4zRnVAPalDPxBbK2HU0d/Cn
bL7NAAIjlqJitFI3sV0kfbWJqTNvdSVoehKLuLpWU0trPj6GPqgpNbWU+PCd6V2K
HAeC0QMjVoYL4UIsP/isYbWSj8NgRRZt5LZY14K0q1gsRAcWX0H9iM/8D4xJBSM+
NfmdrB6qFzczQdKFY19JdasGBwB+TrLDhqVGDHBN8GrNZobQGWaJK33f6iv+bvuG
qoOKuMX9FwhnMu0vUnNGYwkNCm3tD/FA0K86vNyaLHrSfnrFTQTybiTLMK2tQbI8
armjhFGkKNLCPLnNf1pFd8WfVGT73Y3LpFZ09ibYTmeMd6HHbkeC36j6IavrHZTP
VnNwQXqGgDZmEQi5oofUmuoHEtDMGIXdhoEC92Nm7tGsQQ2DZPYZQg85IP9q7yRy
A4TnQ+l010JEfMcGdTdZLgNS27n0Wv3HEch6SKGjz2NeIayqrRX0AnfQvJvOYi2d
1e8iJMTTWBzyFTr5jGcqVNHivK09rcV7wsOkHdndFHUsGKfCkEK1II14fjqWQDCg
vbeZsXb9ujalK165eeFOmpT2XWOr9k+5M0sVwSD8CveWX6BCKnogLTBedGP5z9tt
qni4ChVoRTnOobox2O534xh7JhMwt2rZym4i+T5O3SnrDR8YjmWPE8LbUm85lFI4
0QPSlztZHTIPDRjtJY6Xbsx+wIWj8K0S6cer9JdtiQV54LXqeziB5s6IU2d0r61x
XqFZEkeckuS3pnDYmvH1IKMOU7FlQ8gTMntBIYpOV+bpF4HN+20YcCbwuntKxAos
JUN4hloyMP+2R+ARS57Qs56oAezV/hUbz/xKa+r9ovgbYTO2hVVzCrGAssc6CI2h
EIVEEDA4O+/82JzHWik/Nz1mBu+JNN3RvIKjq6MQdPjS3eyPNpW3wbMY1lMYaH/d
cysiAKB2fNxRKBPrzjWMwdMHKdRxlESKZ94M8jwNWyZrj4q+zmfyZRdZPT/85udv
RVzhOQDt5OUE6qEQFEzNBklIb189S3ERqg1D99cjUFtyBDvisaCnHl9e/vvx+67Z
7L1NvScoBRfMQI4g5YTXhymJV4yRN6yXLlt6Iln7TAavS/YJ8Yy4FKbtwFv6IaL1
R6TQT/IPOw0LYA+Ydpb08cQPCBIC+kkWBcULmJywSIduftT6IkLdC93P4Y+mHHso
fm4XwYFKvnMB0yOwZZiKdU1GHBKQGRsnkQbq9FqotT+w1M1YkrLFVj8MfMad0iMY
cacHjizB6fXvVYTBuvyDEgaLH5AMVPSnwLYDJWJcmQOUQG5uepBkhKQVClkgFzXu
8nm3LjaSE/OUi0Ptt+f3ht3tdkRk5f2d07Fd3uWY2ZUFF9HqQJ/4cfaCXMQoEDNR
RIIL5kBhfVrTk4bRp0+ugUzKzh1kpopNhZSyRzduY3uGxvIJXenJ5F2OmIopq+dG
xsJsIR23cv2FqVFeAwWt5QCkLd3lRBT1nmCRNwo5u3V3Wu44aNqflhLr6esvr2f7
UO86Ddgu5ThPx/q0rWKnhXhwrRHzABKRiCTka9E7Pg4i8BFFvXsIZ8P6d9kwXLXg
dWqzBdRtsDhGdDWzwPvUPc/L9ylfKix5M2ZFPND7bB7lMbfHl4FfAFX3CFH40Qhe
xY/eZ1pyvgLrPdBGX+zMxz6roG6GMBLEv+KiX2xrZu8MzZfoq1nDhTsYUGTW1k1T
ivBpzOnZcEaRWYAIbpGJHgV85z04PcUM4Mg5/DPe9DbqZtjPm8YQl84Xk6MOf3Th
ef3dPZha8HzPIwUfCY+xFeot950FOJ9n8NI/8Ky9gH+w9hP2qMLrk/U+4/D9MpiQ
lXyLW7nzhKvufLSyoVPxR/ZIkji7f0AQJOPPp807dEeFA2j0EjeBkD01Sg4gOZmM
Vgme1cLAo5YyTaCJCLmueFjOs3XsjmZhFKEuNS4WXcN76IaIF0Ti+ZxbfFIK9vQ+
crnjGnRlW2b0T9Wet+yxp7AzxkfqFdJNkf8JSTzQ3XXjQqMGyjtPBHlecK176ykW
dHuZq37xehuE/WirsQFdJmbd/qYsBqoEuc27i3ib35Ga18tMBlPJHS7DuNWkvKTN
ZQjHI6P1awVgLCTtDMrdGM14L1VFdhq1LlHcRxTTEghBGcoyLMPzfXftC8uB8pid
9ZYPPmPIhVRvusW+bl534UqyF1X1IcEEArl18hYeaH9XaP20uQmFvrjT2L6G9HJC
LmFusxzj0BYdHbyLqF/kTR1lGi0uQ4GNdwYCw2Wjh2PfQAaXiru+hZo+yLJHWQAP
67Cea82LQSkPOsfsszIRWQ91mduM/2Yd5MQPUsqT5bJajliMOcMWmp0kxPE0pWCR
LjOjTyKsxjIB/C5YW1lA4Hl7tO2c+Z5hIvcZc21woUOgntYF3XQSS5iq03MEv3Bk
gJ9CBIq2fgyrMEGft+ssmBeVzEnaDWT/ltc6R4t3yI4Q6VB+AzjgKVTWXDjdNu24
HH+xXmT8JFDW19omvhaAgrMltkF6z12YybMSfcvI6GlSMTPLI4Zqxn4RL8dCXpSL
W+wSOkFk27n3WHkxuzPlnuE5dNgaQNDhnlfsAAXh6AFlELAusg6nxfqrMyNMwxbz
UUCSUNe+JY7Y85nGgo8PzdGM6VgGQFcfRhrXiAg/ymH5e59otUg6y0d81UOqIKqB
zNjbq/84t4yw2fljzzlUcVhm0BJ4VBIb7kuDkU7fHCvoZaLuNoGfQQzea9AeWnx1
xByXPXC9rJ5OVWA4XYWOwM/+tq6iYfwa62SdogmJ6tIPZPeKfFjn8pyaQyl1ekyy
MLYxYaoFkXlcZggvTJ080O0qir6PXHnVHGE/kJukLDADwf928ZwBauxWq/ls1/Zn
RezuorWJSGP0jkPO1jt2YwcHEfi/qhOsssZiPitkoshvU/EM2/uZxwt6eLF6Cb5O
a6sI9FtJy7rD7snBKMMPXVIzS4hjHGfNq8oB3GXAnqU41GBwlQpgVezjSoH1QjWc
qqHC1nWlV4xWVgOi5YvZ/X+vam6hCq4X9BPvqFjBe5xzq6KyhlphD2Dyt+mbW1xQ
9RheEC8bKfa12epCzz0o19RZAHsUoGZusNQAlPz8HZ7ItPig6xnnmn/7PXJEZetx
c4TgS8qUlJ1Jgu2yRY7O9nptAMq5CHK+kfoir1RwDXXZXJGf2BmBChfMJUL2Gp6t
cclO+cgrpiGqBGf5ln2GDc8M7OPsTMXACCz1ZMfFFyO4JxhuwZaD9nd3QDmC5m5R
msKdmCTCQmOedv/zDLnG24HO/UdZB5vmkTp+PwS8NrU116a+W/VwapRBv6qSQT0A
PxtL35FL/aTaJ3jRiE+xGUT7ogOXGYsmoCSUNxBn7BsApJHrtiKKOv5YwlnXFV87
cGXs0EqiN074fBpGZKSQjUriE/FwfC6T+r8YopLt6/aa+QSrZW+cOGfugcKOlbPK
b04knS6K0TXuAV+j/IQIZBXAKnZsb7s23jeCrHu29FJlNFhKc8FTYKtkNJDRwmkV
HRUxl6QtYt6nQ+6g/pK5+pPTuqtJZcG7tdg0JR3WqxnijoeGbWdZIHXEW1gA15y2
AhmkWiXyBYn8OJCZFumrwy3+D0ee15nJNSjQlYVumloHslqC69KZGj0f8yWsRyex
Flu3u5jfePUX5JpvFy6fIONQnJpIKWF4RUcQ6O9dL8DkubCdFTmbQ7Erx7Z8Ae9e
UKW9r5JlIUFERyEkT9BuuD8YsdTppO6W9mdgUlkma+F7Iu/YoAe2mJn5wLny+7lb
b3SekEToIILj4XoNryHYV4pnVFlExU4OKbvLR9l+QBTsMiVOEpWntCLjGop3RD8S
+UArKtFIR2funhcelBuIT/PX7JAWB9xBHX4BsMno9UJy7mDZrkDjsPiKnJ3P+jER
vJ7MvMVtVKd4+NwPw4l/LSOZVjoGnsH6XGGBnjb1y6p/B5aOhAQfNB8OihctNj67
inus8EsZEi2VQ+yoeJCHLHwkJK7lSSp43FFB2J1UDAdCjiPGJMApjzEzxqozrF9j
BMOcIj5AtDcfDKZ3meOHBgLAkkD2ZifDO2V+vP346RqogzDoWOL1gM+2PzYjj4vo
tEaC+rrGoX/tehgripKAuVdV6CXfgydDSfaqzbMiaVKGZIOMHGpOs8G5/oiGaHH8
ejjXp5LBCizx/lFBVvmkA4BVnHbEkb7uuRkkLsYowzrHpcMgABfFunQd7HS9gtJF
eZ1h/PwAJ9yBwhXKOP6KrJWG00Tksmp272LcX4GP26LUAlJg04WsuF4PoWNK8mJA
L4p4d5IUiKYPEA9VV4RUCmjVcFPlciVwOwYLbxXI2Dlk+qdLAr1rGTWvArNzHzas
wX42zFQdcy0bIB5zXaXTqsUODP3V7666sCGjS2JP9QtMBEuQJoq3wKCM4INUc1p8
mYOPzxWIsXaFK/wd2LPa96s+SeP0TpBt/m0I9YSD8vdOuwlGfPxyXiuZnUsk47wy
c/F+47UwdDid4mFanHNBM50kFQJyqGPwTjyFNZci0+H1Q9WYIE0fwS/FBS8L/LbN
E6C45jvsT9h41Ck49ZPNgtqbOR5uGuekSZeByE0fGG+1HzReLfsJx0upASm3ZKfz
Sh0PqCSRdtc0UqDNuMdK8UZudJL+rsRlzfRgOn2IkDdY0WfAq5qDSZH+OElbhajK
9olp9VtM9FZTGWyGGlPtlUvVntjRwJCiClje5XB1/FnZUIbbyN9v3d+XMry+W6nf
3yRM25sk45y2xN79d/ka8f5v5jDPkWlK9KRpkajb/HbNPHh/qyskpc9GP+xZAldA
J+ZkECwIGP/opPOTnvGVDMSwUTi6PGlJq7cdnLa3I/eZTW+1y+dmGMBBqPrCvvQO
UUUxZZ216EsNu6STfR+e5wDkvPSoQ8sVKuM2bX4faTnh/P1xOM0JLaNZU11rX8lW
CT8w9M0jRh9QVUEyPdoVKuQaaA05xlDKFzoH5vg8vxGCe1FcaZfZjZMbTp5JKGO4
LiXWSwbj+natwtRti2PSXTODnnzj2quYxiYOV5mXdcC/+UE+bhK8G2OX0Ssmlv1E
ikymxIscfEwGkbePjpa7CDW2vP4VKu/t7sFaZY5yLLD6KwsXnYxxPvCVutoSIWxO
m5b8bjK1TPHWVRwT/g5CPFdITLNVDs0DlxLEu1mSKTndFTCDBIHoJcyr3hqQKRN0
GO0oG39evFTS3yWTjCDA+SBTudbz/ep0PW0NUdqDhcMgFx+xeCcufYka8sJjn0uA
91I36QVaSEFGHgC6idLrN09CWpm7E0etgZhMI8ILBTHoFDGr9ZBE/xWLfxoiUfXQ
t1GRDyYRGnueyWVooYN8FsEZO8pmES6BdmVe4sB5JRNDb6tpJGO0i8JOaKmxk7pO
SSMZKeKvN7gSg+rS6QXxQraSZds1EKuT3weCyFN3curl1AXUs2ZVzekZJ7a+WilY
1nxnrLDfZ9TxQ6oJ2k0m80CHdpFYIbyll7KacwmBDcV9JmeTjhGZ1PJqqbjdrpDP
n3ojZ9SX7PsADEoOFJx9CGUQyOkudmGT8BqZok9w1zqP1wjSKCZqpoqCaUajPtQI
O2vlPk9T5e5pFY0xNk0QfGfwOOQRLmZaYt5NFYEOTjD9lIEdhTUTMV7Ow/uUzA0D
hcYUenrq6L3L9FRBIPpyOAm8DJ3nqKDaxFvPjlIJlTkPYgrlf+n56y2604hEosdZ
0edJcgaCYRa2WXo5o8Lc7v9fgOW2YotasT5UYfJgMEaDM7SJ+rWoaqVVNxxmc3T0
JSRT/4wZgQxgIQMaaMuTkNeHiIqepmcZGYc+ON2yiBKoOC3eolCQ1DxNTraQO4lI
MTnxTWfLjZpj6JMaHdRDUEJlnaxig3AG3Pgub/zrc4RMIMHiM1ju2okaCIcCA/kk
PNrPZzxSr147U0bR+wJKj6IQRmwtU7niz1nr2Y+1DYWdielxtXR8uHsdasjpso2X
T1cKpemrjmHKNXuo6G20oraqw2Bbfz1k40EOmwOaT89cHF91Z+pZYlkfmn1kcedy
AMN+EUi/BYMD0cwjctt35jNs/z3kes5pt3pKMCSwlTpqg5NvT/kyO/Zusjf3G+e5
CFEvgbBu07LR+hwnvKxU+DtDCpN9hRErNj+ipBzuOCli8UaimnSUL4ePgWXPm+ez
DDRzOfNK0pDPQ6B5lY9p32d2reMkGPMUWcFvXwCcLWoO4+qLgMFSI/h0FPJ/V4BG
DksTLboWoefm1wQu105HyVZF4xwIP7xFIeKe6loNVqu4+XZsTlAAYi7vBwfhse3+
EbxJe1W3IHu/xS18ImGmrinlArB1MqOvUs9T77A00tjAUd93GI33tYvurL0a7IPV
naBUPc7YlWkEiXX27r6SQ85lglp36GAPmvpcaYe2cHw2ywbgnW/4Mz9RMQosNENJ
ieSvZyU2iRaS/i/GiWCOY7BNpIIycybRFq0EODJECZalMR1ZN7NQSpp9ZpnxCFui
To5v1ypyuSGM/zYYmyBtlOVkN25D7WpDDdXNCqg5BYrygKkoedy9lJTGY7IJ6xOU
GiguRC54qryamhJjOY9fkmK2TSGwER/chNcZsHEVHx8mVnXPtuX30P6sNdXmCoYF
DRYdxqhOZO3OO5TGjCsGO751QktCLOmN4FTGpE1eJ/oQm9kk6/mNKyNwzF6h1Hi6
XA4BGQjUQ4cT/KjMD2eKzrVXnM2+bIEAbShMIa2kMzOAAPOkxFCQI3lNp6bBMbg9
SvUoMDA27PBTsb5Fv3UfDDqln8miQC2ZvtdgaJQXCOMi/dHv8ebOUS63kp6USJpz
cz55oVpgQRDE45/NF1LuKhEGzJlARlV5RWdVazr9Ax/GJKSsiSoM81qDHWuHX9/0
lref/6UAuFezzrXXbgMwWiEnokIj5QBEweSIrqdjCFUBCjI/sJDanDwdrheVzwWL
HvKejouXvp2dNmyOsJ+mEsw7Iuob2qzXdhzx2jwH24zxs3nWoue4DJ7TLtBbfwa2
rcqO7vW3otN+Y5jHgOpU04kfVYGSNLeXhFE4LJU9hSNS0YoGrSyRejIHQU5u6HiB
KEeckl5X4eAL5ngsdO/pbfGIHaUSsb5kd2DdTb6Qh1rQ5chOxUpPKsSVpdF5NPlN
zAUPseKmpRi+mPtdeUBOvpXHBaYcgAfbeHTtXqnfRkQ+ihDbKfeHC5uPx7zyu4qC
sSYb6XZYyipxAIyskuJHNQS68M6Yj+SPZ7QXTLNvDx9t8WeLaS+y1lavBjGRVIta
ENJbmi5BpcVtcoHJexHXAIR0d1MeHNwL2D530qs3yMq6fdUW1WpkWreNKgUxdSFF
zvlYwf6izKxr2ycrmWZEQize+q9qZHiLFvZ5A3hN+SKG5NXlQHRCJy5wGPKrxr95
UFr8c8qTcBdvQsxYRZVKnlj0kpEYgWhVF2IzFXAcJKMoxsP4Gh959BhzJASf9+WX
0UXSddGHdKyeNOJk61kw3QOMgx8JGs9bdu/ItUDc1rOptmnmkzCLzVVoR18hpuZa
cFAz1dgdsDWc+xIJB3puhF3jSxM6AhO6PuP25zk69n72RE0bhJhOkMNKveY4jMlx
3sCNljr51vVYnj+D/hXGE49wODKnUB86Q/HMbCnzS6U+U05DXpYDK5Qw5w5FtBqt
biszVltBo9CmLOltMn2u0lGRP+denp/zx/2paKUFK4JbTMlm53y9dUzaxxJ1lg4u
8qTN7Yrm5G85RunLA6Ar3ZMFe3cOAB3XaPmv0LJFNvLNlEgwERb4k8CzrMaBcfWP
ZK7mNNVgtezBDGQ1Ikb1ZhIajZA+JBYiQkkXsXUOVeo08/cNEGaCnsxnGGfkJ2/l
uKBxV5izUcg48Cvex2J8Q5QFbyxuNalF7OitATqFqfD6WriGZAmqza2WG/CEdxGs
FWwtX7VSsjgBzd6pX1KAvReJ5vtIeCdR97QWVsgNIEvVMIGQksiaiMQLzuGAouNB
GFQBSPGtZH9ObLd8W7xH3WCf1IsObeeZ/bvsUy3wU9mlS8HkjddadkZmUOux52uK
C+uIyZ2E8qY3ZsLICaH3DeiOS905LnDH0mVKQ9wBaccui6zY2l7JVSoUEflNPFoE
Ni37A0Pz7qSJoQPL4D2/JzBvtdc3xWrw/SF1uCO301nCbuiECDMmYBjbOEd5CLs9
827RWOF2ca9gSrLtUDxKoOxKs/TwMA8u2a1qVgH84YiszDUtHsxGJuQMQmBj8YGn
/Bp5YrDt08XbmW4iOlwYU4ZE8LwFJyImUs1xejNFX35csEvIZ9pZihv+dsqFuCPB
QXZRJR0cLHNxaMGfMHDDeIl4yJzndcUMNOS1MLln8okYvWsKQns3i7EzJnrR2ZM+
q3ctORCugtjEqx0ZMsexz1J9neeRqPvbnIiBoWxhSZ2KW/B6SLOSAKg9LhnDV77X
BXjmlSWmXSaFWTK7YvtFq0GA3QPGaPfFedz3Rx++C/evDkq405Ek01JD9Gxe3+ue
OFqEeQzyg8er8CEfqpFu1GlDDogU06gUjndVOofnOIBeWooUmoZioiIwyCmr46FX
BEIGJN5ROrzixOHiuBvhoha2a9Jo+DGM6gN4dRxh1E8zMHU+EOYPoEUyQhM+H/Ug
4CRv9OPa65Nd07dlGxX/hcJ5v6rgb9pFRZSzoGhg7WL7/je5pXoCHsv5YCP2dqYH
jUAgsGXVSVk8JRt5ryn1W2VYRBmMqVnbtmmS1s9vhzGqlJf3fjJ4U/hqkBiA7T2u
KxA/GenizFALKEBM/NrbTx6qghNBNW22QEA8p8GsQ0vHhiFEeFZxq8x+vfhjn9L5
+MDf3fsy1zdCjABsyVth07sRC5riE6tU6UoXsaG7POiFNE1qVjm71+4pfK+NuELh
K30GMhZ1O4O1utVT07/6eMkPDSNFsbMe90XYLrjU0r78WqPgrAUgxLSgWOk84hqI
PPaZnzDpXcnx07hWkPq6FmtnDvqyEjw0b6Bg25CIFb0Qq4wUC2xu2zsO+mLLvGrw
hqjtDRIstDjXfCjCXMeeUappiBJa1+jvYzXYLBn3vrARAPNEC4Hdg9UFv3d2djJb
sAnKe55Vm1YBSH1UgzAbrxw0guDq8jjy9XUqo4DNXzyzpmkcpckSdrBLnci2b1xP
8sgGUZscMEejETz2SUZVtnl7sazZ8iYyr3vAt4HybMBtJyny+xhieHWUVtq3QZNT
EPPu3OexLEOxcTRAzrrrVxZ1oorJIIUeXkHb6gJc9jZnIPPxk03Z2eDnOTj4qPMv
sgTgvcI+ZRNZzd3bpaC7sWjbTFIPauFJQuXI/VSKrOnvhe/yxgkp2ErLAe2DiP3a
lHbhpbCuzJ7pnAdgrmWwGU8G1j520aE3/hL2UiWwXkltBR8McIe7Lj8Tc4tTToUy
1+twxMHyvIBaYT/WYReMUg==
`pragma protect end_protected
