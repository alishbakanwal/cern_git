// frameclk_pll.v

// Generated using ACDS version 16.0 211

`timescale 1 ps / 1 ps
module frameclk_pll (
		input  wire [4:0] cntsel,           //           cntsel.cntsel
		output wire       locked,           //           locked.export
		input  wire [2:0] num_phase_shifts, // num_phase_shifts.num_phase_shifts
		output wire       outclk_0,         //          outclk0.clk
		output wire       phase_done,       //       phase_done.phase_done
		input  wire       phase_en,         //         phase_en.phase_en
		input  wire       refclk,           //           refclk.clk
		input  wire       rst,              //            reset.reset
		input  wire       scanclk,          //          scanclk.scanclk
		input  wire       updn              //             updn.updn
	);

	frameclk_pll_altera_iopll_160_tnwlaai iopll_0 (
		.rst              (rst),              //            reset.reset
		.refclk           (refclk),           //           refclk.clk
		.locked           (locked),           //           locked.export
		.scanclk          (scanclk),          //          scanclk.scanclk
		.phase_en         (phase_en),         //         phase_en.phase_en
		.updn             (updn),             //             updn.updn
		.cntsel           (cntsel),           //           cntsel.cntsel
		.phase_done       (phase_done),       //       phase_done.phase_done
		.num_phase_shifts (num_phase_shifts), // num_phase_shifts.num_phase_shifts
		.outclk_0         (outclk_0)          //          outclk0.clk
	);

endmodule
