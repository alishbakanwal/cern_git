// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:17 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Pj8ZhCUefOKAb6OzVgyt5/OrQrXuTq3MGYQxJnXVm0HmsM5romEZSp7EyJkEQZrd
qYQSASqIr0OToc/PQVz8EWyscKR8H2GoHXoVgqbHW/Gpa19Qx04HaZNESDKlzBIg
VGVOJA+f3TDBRn5NtOaQFZkaUYkFgH0yqsP6Oe8aFg0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 128304)
r6/vYGIR5wrYmTwOlo6sn0Ca6sCPZwXQ6H/xn9mZTsKswZmPg/sacEID7QZOxrx4
KRBohf3VEg2QtMEF4VsBpVkgsIsQkosnSWTxKD62XZOuX6YZQz/nQ6V04c0+9fXv
26YRKpYaDZxOgUFOY9SV45Co+ytrfUjhb3kNHP/jHiZ50BA7g2xIKALT0v+CwSeL
7HK26W1260UXaKEnlO7zerMYm4eTgSQAiAXDx3Rqm4+Q/uTOYLprHE0sFHSyidbR
sY3t31MV52dnIs67IGDS7KBS6BUV0WN5YHzL23OjG0iJOf9IDxFuF3dJg41xj3bC
oEWLBa393F9P+lVJ0Z7gbo+TPFmFTC2vKUYh5MSJDWlu9gmfsW4JLYsUXSRdA/4W
ygh9A39Vi7Noxo15/nWJooVJRLGU84Gy1EKN9nbchpDnY31Gjot9AEAUsjL3CDSd
hgG6Drv0ltCIMg2H93ZKaW9ra2jpiYczKKVtNWXKeRALXufIx99xBm3DVtXA4Y+5
G3uTjk6CV+WFi9QWqo7Zmno9PqJeT1YcXrYn2RTzDJpTjZQmP2A184hY25h/scGc
hyWs6pr2Sx/9QYOfdzPY3QB1pvjtXm6TPcghXlqntOM3eiVgKmYdt5Cyyp3/3pFW
eiVXOELmF/FmMyJqTAd9PLrBYj9IAfEW8X6mrtWnGQbufZAQXZCKoDjJaLoCMskf
b7fO9Qax/rtycTvR3chfqgSqZ+p1+FYkC57hHdSTpRYDxBGCkCf+hxO0P2ZDnnnH
yiRjYhWycUsUdgeBHrTyjMiP4V9Xf7zy7JCel34JGjkewA5mIWS9E+xIu5pmFltP
K3uVq4jBACOOO0QoyB1mK6dhuj+7lO+wD9gHZ8xUxCzMIrsxJ+gTZSCyKf62FMIT
vci+auH7JumhKxcmoTauiY5n4lyGWC1ph/2Kyi7OGC1Bwo6uxcjheA9vQiXtmrrN
f2pn0f4nYzIi3RFsswu3UMPytrQsMIUYthkyu2cUdYSbrgOrzGoSdhnZ1D8IZp1q
8Ff2UCCOzbz5TxQDcJA4+9jmyl8/wH8haWt0dLywvcjV3OAtGgeo6dj5/O86r1cS
m5EeB44dHRw8zNaSKYpWfH2eyy/6TcAekNw8XQo9dVQLbfXHrMnBo/msJZr/ohdp
JUDGaQEL0JsmRw2CG7rox/9fST+ae3PkLqzPXWzYIY06TCBfmOj5ljFNb28AUSjU
hXXapn8TpDr4HtLI5ZsP1hJGsVU4vfe/MFOczRbJJXdz2c1VnuaxvSCJ2CqqB0xy
+uSihoMQiEoNNifv7DxRO+VFvJdGPVkPtHgAtY2llu45AhOIrzPlQyEevpPIkFqI
iGArtBcWiyfpCowb46rGFQjUDr4JXpkLjQsB1X5TxVCz9dNOKp3myGY1OWc4emQ9
zlumPuSmigbdZfAwsx8O7l2FnFPPwVMwlB5fypoYVt1sLoMzHaYeA8K6qH0x1T5s
p7FoN5qV17KAdny7/8YCan12xCnlsHqSkAx4iv5ffGNoz/gwrtTFJJON3OgnFJ30
ZkBlD+xArlWEwc9d/qM5h4WhceIu4rLnh1yYXGBWYprkXj1dPqJW4/MqFOH9DO0f
ryczkESoQNhD8CiXYRe491ObQ2yxi3AXTgxnYXoi/DGUu4j6QOuOHNfiIyVhnHz+
ZqMnMikp0kXp8wz/KY/ILIBwK775eXOWlgqEuDqn7VHvrNe0saePBHdNi0yU4/s9
zCKcgZXezM4P1E6V1BUO2sr8Q72dQYyAg7ePlAmdAB+NfEVI8PQNOvudLxBRZkuN
kmxAJ0Lo6bRCIOQpNrAnXiSAa8qLmm9zwIdztOy3PWQvaT3V3Tu8+EUpYFd2hP4e
4RaGfnr5FJuui3kFMlq6n9wlBv0UgSgFvuar1rRlrnDPmtYmOYzplTUA9LqcS5Uw
gqHBCcUSDt424Y/hKn/ClX6OOprgpXMs9ot7DsuiASMeHExyKQnazi2+h0HzwxvL
fGL+jSPA1lnxGH0JGUJUIcCC3/C4oOz66d/oDgBaYDeWxJNvP4HtRN/mXiSDyLKd
R4+qNEIW2lTlQN1NEeEyX5TErkx3UTdEFtvEwJq2yoWprHhmeOZV+8qcM1xcJmAc
BEIQwzwv9f5I+fBwdT4fwo9QuFVwKFwxuc8PbAgnUfC0rTsYckVhdAJMDZ62GQMd
ArPoJQ1TDm/v5dNhlh+zg1wBHJV1k4d6776HoTzw99lRwXolFHyz1QidHGvczPps
idx/pbP0yt6J8z6MNdMz+owqa6c1nwwNHYqVCdSofVNuUyQoJjfc0ayMEiRCWXiq
4/IEKfBoxNDra81Mr/rr/LTHI7CKCaA9N6pEwcXXHt7sP1K6P9h+df7PNpUqpy96
WY052yNBgYTY3WAl2glrJcPFv8cQt0gTrEOGhmjywqQvWgkrBstkAXcae7ba/Svn
JXTmy27w8wW7z7Y4O6mRlnT9NWUD36OxlkDZEXGF2F0/nutJ55OPsO8nKuMxu13b
xF7eRTLa1RIzQ2269lfYmEdTzO/dB8LUo2Dc0IPk0KNumwanuRBpVYoJ7BLLz1/7
3eAcj93Si3vTMrRRbd1LvgACufd9El2cCapD/N5lTBkVApDsgCBEcit3zhUy0ISR
HBTY4yYp4g995fjEkGl/hJYpxDl44kntfXjV3fr0/+JIYDt29Mp0Xrf1y7F9m6Zn
SZ3C1KwyHOhY99UaKDAhu3EbEr2amGjE5792dD4Av0xkiPwAgjvXccnYhVYp/x/c
ouo7lvdQQ96MZD2IqElQmFprodnvdVpWJZTFbzWVTL2BGPiSSHXj+qA6pJNMFh0G
CNyHyixVv4zk8XTEHdR3N98lHx4OtcSYHs9N0ldm3wHUEeR4QnjAOgzr9hHsehUl
v7O/WaQlpfQWEqsPFS6pJJvixLt7/5MGk3eQgw34X6jJn+1XTVHd/6qkNAUmOhEr
nEM8SD52eoVWYPxmpJRtel3Lr0SGpU66L4K7J1ax4VFQFF4lekiC/x0rFVBLkCX4
+gj9sGI4WcALzNyENai6oqa21cNPSddVBMNCtiPSRGKceer6i7WqnR4CIG7hiQu1
IY4ccBMsNTSt+4yJXYnLQ+ZGXIiIDWpprXNfAa1JkIIypPz89uma0sfRFN7tz9z9
J8yxzHYOAVfVy8btLzleZUnM5ZRY5946vdKbaiLEfu51eQv7C4d6Uy+S9qjo5YHf
FG77bCNnY+IDtdRhmdQ/YVHAFV2Uitj4revQndN/LOPLA2o48QJMml2CR8xevB4O
G6nvrgrdzh5+5OtrY7nOVsDeKDdDJQDivkXLIix7FCFG0E4UJMOOJgslha9/dnVo
fVz7KDt+n59PY03vzgGnwvaD3iWLMrfMkg+z3hqpLVN20jM14X8e/7ERll23p6in
irLNhiAsjRKwG0vb2bFhxaEsEWMKh4VizpqK8eanLdXM36b9k9Sztoz28soIjvqU
0t5AG/9EnE2OqupakTABuElCTQzRYeIbrWxY/AbYzQC2DZA13aMDN4wwDh/MaAII
7FAEOju9xziecqOlW5NlY9W2wP2muAkC0s+XyRYif4fLnKVrNzOzWF7Epi2LIDke
u++6ecg1UXSk3zcSJyXmjRgWIBh4K3twzvDLNg6qA7G6ZyHTT2KcsBuXfKFFkBUz
ExBM6t7q4ajdnE6ExKJyB4GzWopDL2BrZibeK4JOQq7aShmrDWATf7x61WerYiDy
nepS3F376HAshrnMRjeTul2s2fTCKhlUmSY+HDdmTRvkSQw9Msy3gJbS+CzyerVT
uEq9AwUs9Gd6gPdPcCpg/4lw08cWYqZBd+1RSrLpkwFM5uEuN0rUWRrBubty5aYc
czH2SZi3HBBRrX3JwdXBRiFGFFj8GjHNx9AkGkxOQZeHwwYEbQnTyUztoFqDgB1E
NH2n8UF26ku43mjOTRtILuDOKsGnOGUKK+lCU1BbEPeV2w4dEPBjrvtdxL1uCyzV
AmNa6+7Z+hbFm/iG1m3oqz5jehLLlgb0iBsUhjYFWWyLiqMbN4dAzSb/h4HMIRQE
z33kBkRrmFVd+ym0W4qDmMa0yFzyb3OeD2Wvx1taHxA18H6GMaAR5ZpGFEDL0qpB
kwDT2xjBg6G5ThCkJUoCsNFP3ZM6Eee0SP/GV41kLFGcPlhsaaU/oyRhvZmZwhyh
+xiDgFls4V+UdPt+L8v/MB+t6EVgqwNFo3YU18lR18mZo3dL8HoNkQtM3+s5S+1o
DerM1EAakcY1knx+hKXqGKqab2SBi+y7NjgeAxsfGXOyd0z+TLPLP0enX+nS9spo
ox3/VBjXRcYSwWx7EBr6IB/ETt7zomEO9WDhgxyEYSJyEee/0BdUXlLZkGnHYIBW
PgWqBH2bnz7s3RIWSLW87dBmS/Oe5BsFjAkpRqd0uI1sYdUVzRvE/PTPHFRId/vP
TKDgbtdaQbw88/GN57eTMd4/xUBl5eWbzCW3d77X+e2JD+Fq600xtnwPJOWlV8SS
c2WKEcCQDHhugyiNyXtpeIv5LDqRrs+o0pUfzZdeONqqL7i8XqM2ekusSDzNcVGg
iHKuXveeJZWf3x5rvkgFmSv7ecIkboTIiI+CcD3BPjmH0x6R8c0eRD6N/Hd0ZlWt
zeHN1InzSb0o250fqvLibf/EmBcE1MzmqGCu7LszQ/myggGSDWA7ZQjTEe6Btuk1
UvzhvWsP3WaVsH7oG5nNj2ap32PdUB30UHBCkxvgezteehS+KMcDjLkum4J7fSUp
ITKKybtjDmfQwCU98ZTBEiT+zH14Ln/aPHSFjsdm6McFLxRzGF900neUMMk4IpT0
TTCTUQx7qnahhnmZ5azs7KSWThemM+KWJCCHOKl7gCJb7jgGkHnw+2yYLW9uE2Rw
/mRiNOQG3bVNg44sCwqpzWZISvsALfsnQhy9WxEAGBPrPA6NXhxC5hwdTZ/HRzVy
SH+b8E4u1Ok/8utWuofiIJwncg98oOkEOB5LkRIKK6Qikau7gsj5VovSbxyY+CGU
qEW+SoE/u7BzhA9IbVAR/4xwY+6pCVyi9v+iJYJwGaxEAFeEKt7gGSjF+pcI9m/E
cImJVvm9rsqYlAga/6aK66JIvwI3LpBmlATWbJ/UTdZh0926e2g1v3ZKC7/v0g3+
154+Xv2MmORyKGJ4xRKoUXe2FJQZPWBAhIu5nXLxwtQ47FHl7PTLgiThgAOgxHQO
cJZ5voe7l4dGpJXwar/zrSAxK2TPooABB85rIOVHoUSQdzN4vc5oL0oNpS6EaiYI
451QOdISpDWgE5ZCGbc7Cwy/4bX2BZfYOQhaNWs+DZF/nfp1IBoEZL897jERFKsO
hFvWKj+Ws1h4lhKW70AtKTm2UbONxvmp3ydoWUhGVFP0r1vxvkr1bTtL9SlD1kDl
ux4FvdHPqMT8AlkBzEbDrXeHQDZfVdDDIENsEreiVwQT+GKEkxUPW1tjWNJg8r4z
ZPY1FMFPw0qiCgHyyeITpMBEerg89Ad2gItKm4JUUOzu/0YMx72oWnVjQQZb7P/T
CLCbWoZfPc9cdB3Fm+hTYylhA4/HB5UukKOkBz09kXkTlLQ36L0BrxR7u4kpBrEp
TF67ycS2j4Pcx6X5eBsWFyjW0v26ompgJgXzXHjWRQb/lWkxjeKMSWj15dxvALvi
VsdsJdy6qiuG+n0nwCY28+P2SN3d+TjvH/ki8NPN6qHvkp9n2eV4hCwp6+xnKHs0
fyMgp5RqOgXNEs/wGugxxVfMe0E8MFlTC5H79DUk9+fQaod/AQ2AbgVsDGFAN4Br
gBrTb7zMZetoI/mT3QNSlcPezCsaDDqGLmxn2j4wf0cgQ02viR8kQx+mpGfPgCW6
k1IKzSC9lNgn2d62LBz89uAacmEFS+DnHDjEIQ2d4LsqA1/ZmIeyz/SbsT9oiZfH
jNPBkDbh4YCeAp8hnjWs4yUML9VC9PC47+OqC+G/iNiyBUiwpzJvyqymnx/4ZpmB
ufNEbL+P0QI88lblXV3X0WU5YFXVBj6twgFNkK/P3ObLPTNE9NyPvyXBT3ikymbv
K1fBZT/bjAxl7tukps/LwA5l8GJHkLv7ASr7oZuEmi2zvKSwRHc5EodD3AJoPJg9
oQo++J2cdZL3EQ0EW/wL6+yldgc3DfLW8GKuCvD+HT1NEqtBy0f2J+vIJ9YnfdE5
pRQ37hIoheF9QxrKt/V0pQfl9DVyluyj99qsuJbuwoGb7MD802LbVlYy7dqXuMld
5a6V+0zsZHNEZHFxArMXeRXW1Wc54dFcEGXyvFuY2CcqsRbt95a04HEu9huiUzq7
FgmxVt1tCISFTpTIDa1Frr6DH6y2agp+UssyZl5AszZkHW6nU3TQC928aDWLZXgz
z0ooUN5e/CETKge+sZE8j0lgRBjkwSgNtUjeOmnVMd4wcGNgC8ucPsiVvTaGobLZ
7NP4ZDjQHeUJI1iOsqxnoX1PUw27eomgkz70Lok5U7dJ4nTzqDl6AsdwyuANU1Ps
Gy9SgqHf+gLRvQ5F5LcEVL506boo3/WxsdTr0kt1trAlkxsVZ+y+AOsalWtXFXJc
dmFHMkPzMmmqt4lZ8rI3ymW/us+f+lgjLihVz7oeLYKEhawzd+fs9tGoP8F8RwBB
t4U/5+iOPW1fUtXwbVuWzmn5Xr2J69eY19QMxtmEpxjU+iLgq+cCnuHkwCNau/7U
Cm/DTeZ0luGgPf85e8lRAwBHMt5AiU3JzFbp77nYGQOaKJAmgpPozJ9lU4EREPz6
6x4MXBHervMwLR0hVKiP3oFywnMws4X2AJO1LbXfYCO1xAHNH2IPdagtd2SLtP2t
PZShM2bV82IrLK/F+/j3zyT4CbyNP5zeAgYnE60WJtKAS5jhJeLU/Yk6l3uSCPKl
aj1HdfIkKTW8oSBMSaJdzzDO2PtWSGCoFzlvfd49ECjCiXKbTJIGLvJW3pI6YxY6
o/LvI/QFj+sdDHeycuYnRK0qJpdx7ZaAAi3PddIOhkaeNpYfphidif7mSEDXr+MC
5R1meXyDOV5xwdDqdfvXhaG4k33lZ/LS7LB9fvaIrvTKeUjoBSPOogIiyCctA1CN
OFSz/yoHvtwgeOpYd9AX0C6Uw3vV8anIXYvQEhNyQ1bUUWEixGFPT9ZdytZiKhM6
KsQZ4NQHWauoil4n7StKs17yFzFa7IQ/V6BtPll8xVdIYHPJm0njnuXpmJU7NZC/
zxNtL4p78Wef8Sv4CCuIgPsDGxM2svsm8JCgZlzGd1XiDTm/zwK5GBeUCrOBcqQb
1ukHFcVw6Pqlb7eg5PTdUbxbIkorPRnTg8EMUihgd6+Hw2kWHblR+SAas+anrUXJ
24vW7o8a5XypzDXQxP4xiYi7HodjURqX8rU8Kj81t1vUn11N0vE4tLjcC2WjJBsk
NB6HuPUWtw0nSRFDi0P4vQTYefWfcbRraozMyjxp6Dw718ggrLDLH6q9Z7I8jncn
vXx6V/HVD36xKuLk2PJqDFlW4jbkwHbmO5dhFim1GUu2AwtRtanqd+jxqsWVTb+x
MlxZhezkcYHG2xVaxfObmzF0Z24cj4YUgTB2p+ejF4YZ3xurCxA6CDteyGN95Xzh
KzA6BexgIW0qEAqbn/b3OET4oqRaF3AoMqyNTyoSjddRpIfglzJ3g5DSGIwr0uzg
Ey9nQnMqOyu2xcaLGBfuiKKbuBh2xsvgMSWlH7q2/lmP7DovUTfbCpW2YVt1h2Z/
i0IHzzUh09L09zrCX+KCry6ujWobkWRqfxaSAybPNbtgd6fWJKQ0SD3PYRkrpy7D
h1UPb+tParwSTr9g6ppWPRVSsZf8gdu9s6U4md5BjIbMfzlsSzW6q0sseCY/oS2d
Q2J2/xAb1NuTNX6Gj2q93BsT0RYzn+2ZTd1nUcZIVo90Z02J0mFg0cYQA01OfD8i
JACAKF6FLJ60O5KWR9qioIBIDrxzJloOP/f7XYb+kItGM1FqwJWMRwxwTR6P8IJk
mwRsNpNIbk4lxNSMvVX9lSk+kWFXV8w0a0TMw6yhWi76U5fHcrEV/x4gzxXnfn4H
6LG6jY3/7Me0+KlYk/Zj8UYUbzrm50kcmh/ZG6PqVWuHYFzFw7NJnNNMupQx1b1y
GvY9ue/FAamfh968ZMdHROKgO8vyWryo/R8Kj3Dlhrpv8NnXcsiXxzDE88WOhpiU
F5YipJDrPiW/Ufh+5HM0g9FaegQoV+yeE6Fzu644tzpsPWcTNoWVX/LqASGlk/sr
F6MK/ykwRator/jlCAfUHsd71x/C4se55MOyzjXOUeiNtRBUyK7bkQ02VWoeBtW3
afTO/0gucHnfsnv65Fsa+Fiex22dpfu5YxTBnJTVOyYKvo4xtsdD9uugPEcy1cH1
Qj+D+wNww7VPgbBSBhlVnap6NwbZX6IY7ewk1Sao8HFXvBSL8l6JJy/1HfUo32xR
UgasynxDXXQc495rs92K7E2WRgVFS+egDY8t5tMRIMsib0YlBH/oLRC+0s2A9atS
LmN4Mr542UYSmMFINhLQTRXGX7E3lsjJ29yWv3RoBJnPmh8+KSWi9cwqEUv4lSSE
7vvOgskyCWAGbuLkaUPkNw0wso5oPkM/LuBFD3FZtKz4f0pUJ3Ja9wkKbgfgi0+2
Cuz0Y5y/H1QTlbwTCSrI5JYs27gTHGrkIPh8dwVW/thfWb2XuRX+46LGSaBurtaM
Xx/2DByK4F+LzAxk9tFE+iVxGUXYwcUwjJ35yf8q/5wOL2OiG6I7EzluXC93iuuF
M1wcrffhM7biiRU+LKZA52nigrTjjOGSokMg7SuYqNRK6j/lgkOZ4neyc0LAOfJC
jaFYlt8d+0bHmxcbookGZwVRlo2S9xlkVmS/JGtzzbSCkeIMbVZQYTgFf85Dp+uB
dQnmWoZzg6ppse8Ayx3V4hYkp2pjUIiTtFf60kkLNk1dUKeenkarS8sd7c6veDPh
klp34/6BHX2WlSgy9aRT/wZbiWbXJ0I3HHwVywqg+/YMtW+3x4Bt6r2UFpVBtu1t
ALNMdy5OwR9pho+wPP5kY8mDNGIBq9d5ZKvafp2QlYwao2/j/Ujq+pL4xfASrYJ0
tWF1hir2BqE+SHZsH9Nx3iRXhjNpQ9CS2+HlkOIeCxaSXClFvX5Fi83vzp9lhE5Z
8uVy93Luc7BzxjedWVhFD8BQhlRowAwFKtGJiLtZ0C6MnNRatvQp3lNDAAsmIytf
APu7ZWpsKhurVkKkQXhn27THm8aWWaDpA6ylbnZbm3UTHv7MdP1C6zNqkzCImM2z
sGUbCmz5EDvvvPLgLkhq4eP4XvltuWBMNIhk8IUcR4jIMZqzyjx5E7a/dC/OeYYS
UxEsdUF8b3lLsxQXCEa1L56IDlGaPuAQC9YV1rGqPQG5OCr1njbmExW+gX8agTKv
WvIqmOi5pcO8cGEovIpZROqSuaz2jhpz6pJ0J5JhFVU5QTJMQyQ/5cepzTa7ZSPD
nuEdZqh48uRqa3xYMuuhjaHNsRRQYfy+rXUlZLEPYVgYGEnYyrmeT8h4W5vxwe2q
xLwNgVANcWBMcYOpaEK8XpL+q1AXmhqiHmt/uNMdkZjCMBS7hTkjZf2fevWhgCRT
+V32lphEY1z21a5PabTHO5pb7acIIeZGddXM8Pskuq9ii7GX5T+mQ/3DT9efIv6H
ap01SGHdjdvHBkc4lzuZ5dcWbjoTFpPLQcrt9YCZWCqLYnQOIQhjmjdM+xrY6WsM
nPYL/q2NPiw9EGUmanAULtgUN57y8uP1JvbgEsFaD8oiwWMBYUzENDjbeN1cnq5T
NQUH4jPoChA02zEHzTY9DwkhoMWOs0UeImokW3OH8vpEJcq/iD/vbhKV+ycvQzr0
uraX2Igt9pHUfJSzfqD5YdQS38N4F+ZFjz/NZhqqC3+Kb2gQa7guOUP9NK8Mfi8E
dvbLykCimOpwIwBE06iNt6Y9LCrGURYNc7CUIhAhIhbA2C3aty8RxJ0FGCG43QYV
X99R9ZRbD10o3IdGpj0hoQYRtNYVWTH6JEWr8cF59GHLVz5PSsJ6w5Xqg6rZuYwe
2syJE6VOjlbl7Z2Hesg4GiV80VudflzSQhp96JB6l+g7mMxW0KAflJ+bzIP/E//K
lXR8rwlvaFmeW5TuIqjiFd8GnJBp0/JOuWqwIFoKRuBveY7CaQAKmb4WIMbGociH
Pc4ziUVP60xiK886Pd8iSuFanqGES7hjIIIbcbTzIMhZNCRJ2Rq10FegFlfZt06Z
fCiTXcMr7LHxRPOt2F2zkE9qFGzkrxGyTZ24DdRhbwFCxvGmflxz0ODaK2d1ZpVn
lz0wZnq96CWYrFXNFC61wIg2gOOyrm5noVH5882+ShHTty2ThN4RCA7irtjimUIi
DZ828PgyJwhIXcWCyPzS1ucsy58sy2xSDVyazqcu26JiDqtEEvA+fdnGMNyDIjuN
QPj1lunMqdaetBlkZ9BXCr2Mdrk20Ok1yAS82p2LDmHr14T5zz9pAUGT7JsiQ0fw
d3WbI5efLqi964tHFK3Nd2IcDocP/CFPfPoulYmy+fNCZkExv8U+OMsUzHHDr53Y
KiUOlT/SEz6yTUu0sHyCOZWUBIG71+hlGTutf/8cLTP61ZNDMi1GlZAJOxwz7LDn
V9gS7CC998LtsNoqusl5acKLmO7tbbNUwgAD3yC/QtOfH/I7H9E18T/yrPZ/ylkM
SKwx1tmp+82XDZ6SUZuSCErb5BxV92cABG0GRToTfRAkVR2RcgCIoQPrqbikMqCY
R/5uaWFaDJDT1mAawtOk5nRbW+kmZeuVkegYvCMULdQsknfnQz46oqijih54rMgA
RLM2l6G/6+Sub+6HZ5hii/8i5zqy0K8PBhnEKTHt/rp4iPA6kA19sYmpdNnGN3NB
ePl25zcd6lJ8K2vGaahUnKzgY3w3osLnLAJvzi7jpmvSWtegHxB6slKzbAuWqVeg
hSqMyICTH0GLp2rmcNWgahbZ5OFdLR+LtHeXA8MeHUYmIjunlhj4ZZjI+VbDmCi9
slR4iuBiEsRtV5olyOWu8rk7H7lT0tMSg7ruIaCrGzB8GPh48P1iPkWUGL4E/M7M
vijoGCn9d0pgvi6ZcW8BiU2OMFQnO5fZCNWGGHhr4BnI34bEAibeYoEn/kX4N4ez
dyrMRZozht5USyCvgfBucKomqBRdXsVS0Y/ipuev1ZfqBAMWwk+1oTPhIfO6tcO0
42I6PCTRJ4avlprOW/dCoAhgd2LJWXng4u4P8PDuK8TUikpKNFNQbMBJOWmdd11K
PQj9AyJYEOEvnrCB9t3BBOZ2b7Y7f9MT3HDIIEqtGPMC7sCf9o0U9O0pZJfdNiSn
ZjfqttjkcKf5/+C9vOeJ6t2F3/TRak8iW0KsfcXlDRFcsr9TG+6eQER5EH3vnauZ
AoinOY5+ToHzCPtZDSPGD0LLTWVRE5PXk784pf/nmvXSBe5NB2uoRnlsHy1icVdu
txJz/OzpZJauNVqjcGcckgFHWWntXs7HLGcVGJ23IQ/V26xISjDL58V1OpgfSdCD
6HMePR0y0ZSd1kIgJUJNpANehT50Wc1Filv2/iq2KeaCVZkeaz3RasruY3JU3QA3
u7Jno5jeTKexvu52sgxzHVHxmKKiaxJwtZQNmxAPNk+D0olmIOBcWgmQB610YO8N
Z2U4S3uB1E4A3KjHVrqSyAO/p0UOGOKjzAhbjQ4Lqva5FPjQBhAqi4PYXGJCIANh
0EU1ICvoKyQaju1flXL5FcVxiegdBPrkZEMk5IpS4rTKbQtnPjjncY3UxHwAKqu8
jvXM20rUE8fHz3AOHCbQmXS7lGBxZHSQuM5LygKmWG5DOul5I07ou44NPFGH11XT
yTUQsuGKtfLuBAXjtASUALn2VEKZdTccpQ5EkOsM/jFVV9JdjPya/6U7EZwFCgo4
cgCTu74ioAuxCZjAb4tq86RGSNVQPPeDrb1DXfEAAgpNHDQLTAn185B9Aq6s9POq
wSN4ZWHwHK17U8tHxj95IhrarbZ16J5rRKxJLNgmm1JHaYpfyS43sT0Z++OSYavp
i0JQ+rGx05mFPT0W9TyyrbEpCMRof/jbO5mjOtU2vM5oM21N8VpHARJo0mSFNyPH
yj175udlCTzuqr8m+jwCxWr+mgnoiihxiZgNNYkdmV2mEIY7ZAo/G4rYufl0B5sL
MSiOqWkaJqjdYH5qGakZfwzFnz0pNBFc2ZFqAW/0+EwDnp7put0TsGJMB1IyuQGp
M8bS0x2euDwV75em0dKxcVM8/n4C1fLVx4m/EWpTCndwFev+JGWrOQaK/dxMOFie
+5oVLp5xFeIAVF18F/fJcam1h/XK8iubG9sQrjXl+XtP8Jf7RuG8xiniQc/6zuRv
tQywSxJtpQgUH26WJSJMRIgbQntvfcgampV4rZ5dqT8qssxSTZhkmSj2W77W3rIi
nYpfYAGrxW+g6/sG0ZmSdUPsFmrSnopfoj+OY+Y5F5bW3Og8PWQUt72/eGRwpa0d
6it005cXcQdu/dux7PyCIxkV6hNWsSnm041MJFFVIXxOmxQK0fnwzhSgm9WwtVia
+6JRYdnDOPxvKsuM87WCgiI6eMbZicqFG9dMta66KJrrK9GngIDSrKHRIsqG/QM/
ibUszgGqNFmgoRMb5O2q/znwOdw7ziP/SdnP01rsriRu+ii3TV9wRqPc7S+hPZrV
QIWRtbZsJJfZFmxPMwtW9AEvTsCGQTa7DQv7D3nVWBhALKfKo2UDzGMpQrhxIEBP
B4IlVslFlUlHCkRYGg8knrbu1R5Tw3SRnDEfiDcQavXwAyDYcafb8tbf/5bftIeh
Se/nqCy7IZcZLS8YbCuoGD4Jw2dZ9IruNUlQDvvUT0TuoeMAtJMzEuOTpHzswdMj
8EHfXP8v81RrO++hYdA7M1v+M6KJT5bF1u0MW2AYMr6fmqGKURY5fJOb2BoG0Mwx
zoygTVmCmR1zpqf+YgABnkBHrMvqNbygEFGV1UR01pP9XLJl8OyZ/JcoxCl0elRL
o1uyUMf8i1ZMKFVA2PMODGJoLAzZmIV4cMCKapb9Ci8X/hDrTF/bF1pSVO0I4ONh
l9CdvtTBI2NBdpCSs7fNEakWZiNmp5yRDgoGCwho04McLJAmUx52kq5h3pwXW3/5
SO0Z8pfp6fcNO3MjcJGqcfhJsLWSpubt97oB9Elci0kv0LIE7ZwhGyUiPfxfdWr6
TsreaGbIQy8+CXHqcOWx+ClQAKWxgbAd/OfWRA/acytffi+6REewXHq6wbmtp49M
PPymeJYJmwise9W7pM7Grb0lmCy7zZ9nN8+vG0k0d9Y2BfDON+2Hb7l6v+CXg8dj
U6uYpR/9FFzWqMWgb8QrGXBHqQGOLLSuhZsC//y0YchDlDfXGpnzFTNK5obTelFu
1B9eHGuFLc7olRhb8GxhWE4w1+IfAZ2xh1GvUKaBcUTikVg7SlanWgMooc2Pj24w
z5Km2S3/LlB0+/8VMS5Q1WKIADVH/PXtOQHtmMpXI6lqeisCKj7rcQ4c3B/EY8MW
ODAnaHEO4cuwDcmzZ4oHTbRaJPJUtFc8lz6zlkq9TTuDFuSWBe89+MntEo6OODmy
HHekPT6tX6BIRiVhnhkNRT1yfz/ZybSYl1BCFQDxMunmSxPDLeXDkPvqP5mlHIi3
pJ0c9hvkZcucpe5jz/ieRgzlA5Kb9p4cqGpa7YQcI61Szt6fl9rnTZxZJDhgXxZ9
2Q0In6SR5lZj8Lgz45GggeveuZG5tjQ3CcM/VzEMcGICKtkvVLYhqN8/9NDsaefx
VJVwK4UNcUi136Hl3qfCWOTsyRg+P8xk0AzJIqyzT2tHhZVD8zN2X0hihYaIPdvw
nEFM/ZRqSZisQidazNH9h4EMfJ+Dld5vdbqoodRzeuoaMPpJ6BNavUp23h3piz/H
OwDMlo6l+Kvr227XeJBEccQqa1sG0hIlmPTSmwe7biXKxGzjEmK7shj+Jcv+L/Rt
3xpswKG+FKua8IDUeGrJOSq9ky9eiG+mqAhc8Clze2SL1Bu2ZsOJRY8kd1Y/SdzQ
/LD+ULGbZMvQQVLE+WGBysMMAv91andMqA5Kp8BOVFVXE1lmzgNWCi+OTos9BQDQ
Q9F7Us6hR8kkYs5n8TQTF8WqoPb3GrPUxafaVgL6dl+GhdfkbQQE8t3maLkyTcy5
mPi4dyeZax7uVPwwlEnsf/QapFFfLGYF0vLMiHAVQwqoW/hURvaJsCNTXeJHMAHk
O3iVPLxfKTJd/qGb9KXF/llS0yu6F8GQlzoOrekkd7gEfRT+3/uJzxId3zRd6frZ
h27QJthay+fRNDCDSr/GjiwJn503e505hJ7U0Q4pxj9DRQjjx1yFlT8OSbEXyCOH
0lun2+pMfARFtBw43S216AEdPbwP/KONzJ7pj//epSy+zvbC8NdGCrRDjunirwcm
o8bMXYPselZLuzzsKnKlUyO5MTActqTb1XjxGbkwgvSIHubSiqDhJKZ0DBOCKIyJ
MHyC5wszorFkDQtLdxGmctDTdvhmimPkPFIbBIL3NUBBZ4eTYyg5zbT7dqGG6+DG
ykazccna8/9EsbL6a2R6/qPTbISnNmxddEslvMw+qA8AoYs3zfbos2fpt/2grhBt
ILV/2pBdw8PDYPQ9G0sAXg3GSpgL1WnVc+L3/R+XlUb0Pr74w3M6xJG+tOFxzUtp
8BJP85e90iGOP89tMFfijPxk48N/UiLojUgZ06MzHlNIKcC8QsDpQfhBs6G7bKdx
1wA7nUo9J30dUzwo+EcczHSkbKFRZz2UGhLGFZfliaG05tYzbc1HAUzjOMIu1J9z
1h4HfE07/cewtrfxelFRHD1g2tKLmwYFt1YzHn+nOVIvhSSCSQOmcZaQwxRh9uwc
/qa5t/5Vjp/VA8U0fpsP4Uhhnbmh4T7Ekwtb1SzH7HJI3qy2cpx02swut7/2IZ1x
G8CiBmNto5OPN8jZM3rcKfFAow+e3OkOo3Q2HiOodQOcfSjAQr+xa+ypRUkUuiUo
9GWgMpgqwyCEf6KtLvZSZHFBdI8cWRLhG6F/U5fYetv3mivynTgO4PuDp+oYMWYR
UR2QhPxX2zfSQdieN/ivjykXdKMs1C2yxnUD457oxSMOrku6CTmIkObrSVanIZUK
g6zbMFIDYsT0hSN3kUKGMUBvlaSSVhzAajfKbCd9kEV+W6X0v24SMPV6+f4q9NLW
PePOD2Ef1+geGEScDp3hTUZm+/qzuOytO55z6G0o0SHUu1GVPQDh9xUVtI6BNebC
9C7WVWek/lO2qTAa6qvFZfIEGOC8lZ0nZ/+IqswU1C0yqdbygBzmayzF+6QzP6Zn
CF+biJolS8rkLoXcOz5AoC3heb3qTqygEjUDfKAkBOnTawydhaWp+p2vJCsRMncP
pfteSgIRlZFKQ0JiMgj0LNZd2klmmPtDaMRlwcn0D5WVRr0VSkBJ7Kl3c9WnURxh
DfuoDDlksmlulZpQiT6XisjuvpT38Lv+1dzB4vtq8Hpao0IbcMI5w/ax/MrItVw2
nEPpAar3ijlp7NQ/Sat5vwUCEW6voI1t3IKawOkUSGU641GliFjVF4ekUF7fFCK/
xQFdwaVwWJRrjGsoqpmTEpFQ9pG2f6d/8OT3oSzXtpzc2qmBKFq96at+EICKc8/5
Sa6zT1gefUdUb3+Q9V4niO8e9EN216FbVx5m2bc0S05x6siIYH0SU+9m+GVrx4s/
JE+sH0O03kq6Qs8ENjmALeQqSMSh6UGrYTCFF500mhfYCEHqH9V225dCchbop8JJ
G0T9zL0RP67rLK78yKAy1ncckUBQFAnyNTfSwYrCr5/MiDI1BFa7Wg2C6QFt2pH3
yYXWVRboAzcyZ/ZFIKWufGRDGD+KQykeCEPe7ZMPPV0wzypao1iAyW5vd/lI5EwM
IWwr0ZmUtvGOOnLfh5VhR7EIz6PSVaH6mnMpsASOAi7zpONvUnYKSCOtLHr2leCE
huOVHxxLAO32gMROFB7xGB9Ygc/f9Sr2+ZBlli5NB0O8OLSUSZD2oIBEAiNPZgFo
NbCqIhp/P0DV9DpZMobGch/BtTUGazGkaXyxJAwfTMYqHl9mSEzfnBjznmgbN9J/
+Z3KWwZD1DXhqbDbZtatB7HYIOO3N/Eut3oRfxf5XaZx3tPKZRorUw5oSMgJjfej
etn7bZUD7GKeI6g/yZaLhu/lxz3QlcpACjWucOE+4eGp3AYcjjUFWK1M/hVUlr4M
5GtCNaaecvexbGCy/qjnRZTtwb846/4daZPpSTB4Zxgj1tpGI+wGyczdIBD+vWpV
otEuBMXVGFTWJHyHDmaXI4ieY6Tj/LYV5yYJorSKzsUOT4VrAqKQBlvnKTGh87jX
wndSvJKv+o3SgSCV/rDtn/u+lk+fzihP4E6sjN2lz4YuPZmh+wFwHg3ZmQmr778G
t4MJpBH6/QIzjdRWJuhWp7HB6uOxrVTtk+7X4PKzDvykJ7Exb7SqYO0ejT3KjHWK
SC1wflj/IYlnmibLn2W1c2aMLVokpDswDI/A/QI1/zpsV0nToSA+CLsEexoCalqI
kBCl/uXP8jZr7Q77jn7NPVnKLJrJTbdQ3VG3tMTRQQRVddHFss9SFuYhNuP9YOai
5Pv8kXHVq2SRUUWAMDC+IxpM7W3EV6TiXD1sUDWLqdmk8f6RhD8WIBJM96ZIBW6A
B/RP/ntMmp6NJ6XbAiIayWsasRf2h+uO66AwxqQoKwDF2tZfiLzGGc/3dPVODv3E
TRuBB20cqCJrJjz6a9K1heRJdwl7zMMWntYpd4Bg7SgS+z9CNGTGUsOkzslI1n//
ccuSo5pUkNHs8TbF+0yKxr9GmLq0t1MTA2oGVhrnXPZh2hRkSS7e+n8aF+EMtRzR
6yXcAWjkbuTl+wTeyl5oJbfSwHBaZS2FRLGHr+hens7fChlrpkKCpZlZxz3hjytd
BQZ3lwzzmFn8DKUnNxXj0M4bOz10O/hcldQ5nq2HbHIts3UNhuAyanFD5R2+kXgV
00ADeD7Ybnw763o2kqAad4LfHgNgHE8+jeS0e+y+edG9jt86zv5q28r3X/psje0H
gIHteTPx7C6+zgE2zr6jGmJPdGIjPYBVb2k7JSTglIW6AL7PeFo9dWnKmRzsbjY6
Q4wba2gQeuTVy3LESLg77IoSpBQE68AJPte7LYFFd1Y6Xng9ue5A8i6TJ+qwffgx
lunefsy60T2f/4OkVlBbw0QJOXeRxu2LrpRfS3dFm+/8p6zD6P0L5SUD1Bn8vHAq
AA2aE0A3ecpDoAtBXbNboqewa1iTn4J6wpQoRX3BBA6j/AJ/z3wx+jHdo0XAjg35
PGcW6z3cntayp4n+fmbom743HBRnsSHv5FM36ON2gXTFdVXNom2RxJmiFBj1SfJf
oBgCklDfhkyT21TGmE/bP5+xcEMj1Yqtve2Uu+b1IG1SUh+le170DREqhOu+cNBL
fmeC+wVHzl57QoSJ0FL5igDIJta5DIsGdzbQm9t6xKJG9gWdHFdaFd85SsW4nfYJ
PzfxvcDyOI/t3OVFdEttwu7ZV7CCCQ28xP7iaQCB+gqyb6QMPKFev3lRjriSSAWL
17zvqQLjyFIqohzMS+nB1MolNXm/oApLd48KtiZaLHI2wL7cpjz5KnnGK5y/TWqf
YqPmd0ljRwGyuc+0CUD7vyXzWnE8F9Dh69loGqHxc1Q9QKuqSoXPmPGH3XsujnvV
27HM9iB23dEEhVaW9X0wdwFkjnYjD5wpn+4Ig8vdXEmi1jCeK8MXROumWZpZEk2q
elj6cqkKRXC3EpOLYIHVqMC/jjRW5g0uoIc3QxwkQkC5KE9ky4k8ne7EAeSmsQhT
Ss3GV1gV6tidnUCVM8FbXXmQtnLPvqpUhDN+Q0iWgie1MWCTMoZhU/p/0tYYyJxT
7yNH3QWd6z/uQ67qPvh4VXVWwSV4NqTVXz1bpNFogRYMGspxpcQx7CkydSziANrD
saOw7n4SlGXjGmI1WPzgKRHDnv7WBr5rn/uBF3xfJzIX+5JB58IlSOhXhOo71+Bl
EocHJBzaTHpgJl6hHLV2KZozKNOyCS97NANxbrF7PY+NNyZQ9ux3FnOy7K3Gi3iC
aYz95PyO48QrbU6dMKiA4tAuLOuXdrJwPIYs2kwZYmOLrt8IJxzUMcHmBSpYPfpH
MXPHFIQWd6hgFv4fGot2OdvFw+PhX7tS7Du5e8oIYshz8koAAp/bZHgU4C81G6n0
d1Vf8bD+ndlKHny4GIw/4G/KPyiYPWePAAybCyz5DOaefSSpRBm5+msgIp7dL33L
hEjhDdf56/n36nR8OP2TJ0MHa3oYr2aO9blfE3QaQuKe1hx/o20JFhh2pLbGWF+L
ESh//5R6Oin1SNSIMj4DyBiDBYaZx/u0dxxcEgn5QoTrCxp7+pLoj8TZm15hyxsA
E3UQk/+uTOJyTtODHBFoPjol3iCOkQpJnzxfXjBaQGHaDSvEVlxzlOo4JADaj3km
1mFwdlQO+S3O5QT5np93NjwDAhE8ecS/MNcux7LpFLyrBqZFKgns4WzuH3XHZ8R0
NYWwtazrmo3XYVobv/HJr7FCv3307D92fkwSEENqzHqTb6UDlvsSWaf3Fo1pi45w
A++Pj/ZTvQkd4h8R8zefIUwA0oPzJrE37oQJI1+wLsh/XLdk1LTQyzp80cptvvWS
3zqMPvQeULGggntGLTekBU2ahXb5XwP/6bjOXQ3IkzBdymHVWXr5rR+/SAKKDyZd
qriG7tx/KrJ98VJLopyM5v82j0zLyiwUhOK6WedKb3JOOa/r2XNp1wxWNV9YTM1W
o2lev0IzMq9eic3CJorujOdM5iGDYWrzYoOhqONgdMVfe70y5KF7eoJrLGX874AT
SHAMyPS2UctsCkpOuA7+UxavLbRexs92ZB4qpHg2Jh8/6Sm+2BkeUzh8xahc2cpj
rSZgYn71Bx/fbb+Vj8/kge8BI+/XReoDAZbUErryyKraas0+NAe2X7NJM+kxYkk3
Ro7dAf9NCx2cq8ns6Exv/Sl2V76CWWsgIRv3OmlCWZnZMqru6D/at/69aAPkjRTC
EqnUheq7Ce11U5MCypOptzwpMxNUsIvE044b1gsJUfk+ZMffGGZEU+ujmzNl5oLR
1FI6AvWWVtSgyXVgYRp3QG9u4DoUFMuoTgvxAD4TaxhnuZ2g5j71/0nP/TaedBBg
qXQZx5MtsxpsP824IBMnRJJdXb/yBs0B7CROH/GibzjiQBcGq2yWevQOwc5UHdQe
qnoSiMrtFgmGlp+8pUm59mZxzCOnffVBiSzFBL0DJg1OzMEcUzbj0Urj99wEwZpu
MmvodcUUDWSWGwTEXwnTQu5c87yV0aYXwSldk3KRmhGvbhC+mrUI2Nj2ba6Yi3QL
OG1YCnY1XKC4yM6hWxPV+RlLvaz/FpCGmpmnEipcGRLTkSTm+wEl6gC9WKK9y0dC
z8LS9OXn37kvMjckylpXYDae8EANm0Gl10l3jgCOTsysxpsuqr4fRiKseA0P6iDg
tWKVUDkRDCGhnhFESKf8k6IbMydQc83bMi4ewOhs4ePUVKui+l3z4XR5NeiTSIC8
LfAATi6gjT6cWs9Nl87SLRs+WslSYdVm/HzPaAztIV//M8zT2ajV/nTy2hsQauvt
6aKHKATdBfJ/MUArm2WMq8R5W8MA6m49FzMmR/FNw9o5XLGyH2+PeQisbn5lbud3
oj8lc3EI5A2z7ZFgFHjZmIfEBoBzn4hnNE4/VGhzGbbcAwQfNeVxYj4rzEXgK2mD
bFKWgry1uMfoPGlaQ+vImzG9irGUY7rmPs7LFe+KYOBzRrbcJVC8er8a+QvjrDDc
P+fv9KWhlasxsODt+mp1z2fL4jJXVM0T9qrZ4VdQQjlL03k9uG+doP1mQ6gk8cD+
JkhnbPIujntP+TFbPCmYubEDaTuXOV94oi/Fni3qNkAmTpHP5Y4VV6Av0jMaFvsC
tnU/d/W9ox/4B1yhwNcRdLbmOw/G1tgWevlUtKD6c04K3TK7t166FuiP7AqRxyKz
41m70daI3r1A73ntg83mu8xc0LOW6ooX7uAW1d/znBVsSFGIQrMAkaTtXhxA4rOs
KlUol9/NYVxSf/STIkEm3j4W95qZ311FiU68gdHEHzqOocT3EXTcHvtutUA+L7iA
ch6YDzalzHKiNIk2qhiL1PBjXbpkMKB8h+RG7T78ecV7Y25lNkGSXLSPdlxBPbUI
mEMFNVLbJvTl/0zKPXSv8zexOSnRaDa1z/lkY1vGBYHZJIVbC0zx32E6zMo9UNVx
X1/607LwsWT0jJ3zWmnxpoKtVjvicBJSuSzw6LFsjUhxjTkWif7ps89KH8ggNZPq
YJWTKWK8N+A/AYi/MzQhS7tjHAL3tHSb1Vcg1rtIx1u3RQ7OZFE1ihiKwH/RJ1Xd
OicFBJcAHp0Q+Q4qHW3A9JRrMQ/lPukAt/NJJhG9F1Gv0xTwtecU5hSnnvbfSdSe
o1j8uFzC30b8EhNZLbHZ0HFZ/XOzZzKbgWd2JcIHUFfmrUrLsq1EASoS33GYekUl
ERkCcMsUUDbHjHw2hecoRrZj0zrIss7e0X170Hoh7JAA4riWnjqaNPd4WIuhTIdO
UY8FEXxqDYOg1z+mlKIdnT4GVOKHplnV4eyzkIsIPBmnk3YWw7IoktVQELfyJubx
uB26Gllw4ePQGwRkTY7eQQsLkLJPuq71Sr3jikEtnr240WTxwb1UEdWUYkimmQL9
UUJ34j6OsvlTKsl1skdjH47WPiTNaxBtywuX7PrcoI+1+Ytpnvkv0SzRCujIEoeY
EV9qxjhzfH+lEm0Ne/zyGqAlGFGzW7rtRznjWyMxF55hP2r3ajrxZKRUKIWASDMC
Uk9TGDZtols69fUbbQ8eDfqqUO71h5C6pAQ2q8rkY0E+pY6VyEG+EC1CK1BrL/ld
+H/VdLYrPjvLO6tx2bwrphKLE/a0EwluYdHErC/ZZFUaM0wCZ9tDYRvVnufdwOv1
IlyuKUPboRinUH+yIFGzlT4lpUhuVv1VeNlD19s23NtZ5VU8LLCAMstUrFOirJRD
9pK/yLordp9YS0GolgSShoB0MmJ75gU+dsH7H/Efqvy5WRoCmj+t3gYJ4f8Ap5d5
80JhOSr7K97s+Q4BVgYaBLt8YqyVoqpuMD/LjFm/ZpV3oJuJn/Dj7AmDlCNSnHv4
OkI768U61PZQ+55CD5xp2NG3WValoIaDyTB72RxSFLEt9vb6bYZEYzv9ihDkW0Or
gXAJrLA3RmaceEfqo3k90REV4uoNgE8w0duHPELaTjExgd908PqcS/Ud/psqRtY1
dAQnMhLs7Uk58nhffQUowQcehAo9Mm1UC/mNkO2QhvZtEvick3pdNPp7XBC9A67t
gzypda3u6bd1rqnLNYO2C7k3wz3VBhDalvFY9Zd/J9I27NyaImL+tdEgFnV0rOdr
mtMDuxDErE0h01exEXXGvxZ/e84g2VPATelvAcXcKlX13xnBh6vWgRKYIrP+er6N
48WFyIIZH94KfvhS+XMFaOw3WL5EsIc23SgHJp5VRHQSEfQvlmNEg0JR3XPeLaQ0
5peyGm8uQgbI4liFIqLJjGdsR6qpIiktlMYZv7VivJZoO7UbnK2BaAnYyVTlvscy
XV8opeqHfsLzY02oOPhT5WdkXEzGktWYPuYW+fxVkIPeh7E320hCvUsTAy1mZlSB
+KtvCHAMF5Oh6wvZq0xyasf0FerIhKfwyEn9O15V6P+IMZpvQ/09oUQIKfWxafSu
XWrUzcvXc6NnR2kXlkLpyOnD96i4Fg6kDN1AJV99KJyK3eLMx4WclBGmRINhno/K
WJZso5P1fgPOEo1kUIR7fy1yEm/sdWtt7XcIsCZxGMOLJcCvTw8WTthCJ/9npTTN
J5GgLWU5mtbFgeJrWh59/tAOgZ4lBPMv/62ewR71U0uTNFHfpccPQlxM+hKLSSZf
oINKsQxPPQBTIwYY7A+ci/lwGaapKiLYgDoaTjSj4ZhHIYAhmUwu+UANwCeVbeN6
aZtyOrWd9Wpqr6mcc30lJJnURF8HVdsV0sKmqlhHjtC6nPkXh/SxvXJ0l5LtXs5X
u8tvSQdBhJ9en2SWH4xoIw1a5NB/ufKfRDFjiGLEeJKeZpoZqFDJyU9z9xcSDSmb
AyVl/mMy40/RX8vltf68R/Z1b1bERRWWSmy+I9JzVK3UKD/7DnKdj1gdm8OMasvC
y1cJjcbJrX0t4Mq7GtDTbvb9QY3i0OI8vBtC4KScgHWe8PzpI6AEvHKXDKSgNotz
yqrJyMcB5hV5XCMmEf1/8rp7KelH25bsYg7JPeO32TmgxO4Ml9t7SHoBaeQlymaz
uo+ZG+jUZevV67wVuUENV2YmaLeMN7l7xblSjr54H4IV0CwmQN/rVXZEAMxe2QvF
EMOxYhGETcM0QOgT2Pdts6fS9fNJCn2dzjJvxUyWK9GeO13KVxDx9dpRMiFPHV9U
U2UrWyemBRC1vOxEHt+ZkjQrTIofFebIquyfJyoyfeqoVzyu0Qv/GXc3hW7guGtl
DsdulAkE1a0LjXo0cRW0NFyL+TAjr0Lx+N+039S1Wq8OWoKofUTAsaO9GFN+u5e4
VUfGcKe03wTBVvXwHtvRQQW604/CNle7HCPAlMXdzJSCrdLvDbrR145Yd6Egvh3l
49MgSTMGHImK6ihrkzQxu+VqWfxIFbWbjRHbVDKgUitR31alIt7/V4ey6Wg7VNZ+
iwXAmT5N5feZm8c7IVrnA2lT02WWiTCG5yAaP8o+LXddHri/y4KleZSr5V/hiWfE
iUWxukkdaT9ijpDAgePH5BLvoIX6kQhtRin/nwGCQFqslwpXyWL1di3xA2KYcp6w
IL0bj1mDDrtRxiJX7Wem1137SrcIv9IxmfihdAa10nuK0djPqQLwGHZhDyBnKqYL
uV57odXU2yu9PkEYM1vmhiWUIlerFzRuBLvdulXo+fYKn7kTnrGUOFkUJLjFUOJV
6pU8/m10ieHndplU+EWfMYobWcFiO/hdkdY7/DbHN7/yB8vjE5jQyhsoU/jNJjZN
2nsN66s5jbsTJPmvMzD53Dl/0ppIJrgp2u+urauqQ+zyqPMMSUbjsWuTVVWBP8nd
kWO5WDDgr2vxKlNO69sA60N3WmjfMoBOWdZJ24dWh74eQzt383jmIw367O+exSeP
BI0AwpDxfaDIWJifj4rLyS4neFeGW7iOjXNkLNkfUoqnI0S8OuDnCc/T+IF5OdGe
BbgHtcKZcM+FufWUm0bCvdCGNekb3cbtSraqzrJcDZPAdQFIoTDBqpDyC7smy3q8
dOKayAVgj4P0FTRqWojdt4zjYEeHI2RWa0josm3wCI4CqdX7OAmdgM1Zil19aC9s
vJRcie2Wvil1PqNHclxqjV8nwC7CM+ga5SS/seI0IzZ+nIv1mUW7hIEr4S7PhL6d
eybtxmim7gAaiYZKBbBIydR4Scd9u8BuH6aLhpSkpreLlgL8Bz056tSiDEm0G0aj
zcJzo3keU1DVsOFiQ5Rw8MGV46fuwRZJPsPby8nmLy6UVC0q3o/dezS2rTdQqwcv
8AFvIPO3lYWKlHQC9PLEXGkWw3UD2ja041uAKYU0XoI07dSi/ImjJnHT0O8vuGzi
DHQRLJaRlnIwFY5mpAnRQ2c/FUgIC/huLl7j4Rg0fDednn/TN2fGF1Aq5xkGOhls
kBR2+ZgTnLinKa1obmfbsRhTlI9OmDeNm4yLo7LctaatBBzSzsD+YUJz4hReq86Z
2SzbHZ3OMtLjBL8Yn40d3b6pI7efId1CbMJJqkYa3H+I5hCNtzRt8ezveH6gzCuC
MJvDJ1mvKYvW5BmcC7TBx3IM2H6P4ADcVKIb5fHCVCLxIUZlRxU+B1+yZzAXSW2d
PeIzVfTE9LUe+Broz+0/DojQOVUT+t/lk2X9ffRCfxJqkz/5+FoI/QpYBacXT/CA
3LtRv7Tq0XBKvVfq2Hv1pPvQZgWscD/s/W0fjpgWN6vmdAKIXP/W0TfkqJNNHbj7
wVo3C+SJXSZJT2R/VBd2W1EfXBqwiAghtkMqLkNTLNahWaVxrq2fS2+jJiRRrUkw
j90Pg29RJVtj1El0/rfgcFiJwXqma2izDrs6O8X0cA83Lo6/FPxQwJMeCIGHEg0r
FoG+YiUr31Wv4WKMbK2JVUfglypmQ/WBv51yMVyQw2FxJgyFZjUg7n0uMhViEwLc
Kg06euA9gXO2Rm9B+lKSNGeQFbwIfpDJC305FsoOya3vYgONGsPbwd8syQp6jNqY
fmzis8TTNWwJzxLuNBp08pb7vjJO06lD4+2nPJWqzF3ef0xhDZA7gLSfAoi6jfS9
R3bX+4UAOd6KYzR/+0J0llSCBJWx5rBI5RZt99DHahc3VL///aP3qR7+kzoGS7Di
m5gJ88u394Ev+S+eSeEYxO7NQ4uHhHox6675/6PDZRB9c/eBoC+MDC5RuMpf1UNC
lM53t+NQLgq4f6Gfz6xqqXSbL8iyD7thVxp/En3F/oudrSLuB4G/PZslf9652Qqz
FiUUrfYe1xzW3qvHZnuEB1gSmMu/oCX6LwQMSyRZEyVYyFU/Ej/8W8FX2w84ZKfB
uAzEffAHTWdwBapCSfMwkasbOudR/LvmFlfkerqN5ljrIJO2vx33/5FCEn8QZrT1
cPt5yhuodOUYZVRhsvK7UcdIi00I1aGDSVjdFEozHguxILxg28T8Z3m0nGy53IAi
9SsFGTfXF2Frdg7+yDi17G4LYit6k8hBA3jmDWZdbt452pjN8Zbwo5uToZTbVerN
dmcidaW2HB6lPyASKUS22ZqxgxltGhx0Ei9R80d+6RYvKO5zvnfsVFDS2ve/nHiO
mDg8u/jJSAetw6QZtqYt1NR7WDZRcaaByXaPNvX16PRSHMsH8JNaqSylEv2BMBjZ
V4/e5fq8RT/JkO/JvcY+C+lznWDRPZRhab5uYMWIfOqXSRNUxIMdQcXHJYjOqVha
Fsp0UkwIxmeem+N40MZuDZZ7cc4cd+5WJ6E7op90lX/TloXt+BCzhAqxtWJnoSZp
9vJyPDvYYQLU9fcaECjLbCkQ+CFB+oyxoF8wLGbMhx5b8x1bUHtjPyijy+yG39Zq
62xh87QLP+Q0u+7NIWBBShVaVoQP4U6SehbdHZ/xVrWK38ZFJVbsOwhFzDvdCBr9
RJC1UNibmsX0rI+bOVwYcsYi5sRDFlO8sCA7mBxFJVbMIqIqsSfvsowAlnXHPWga
5j0MPyCAeTj8GQNcsqEfJQRQhn/AsXD9i4fnV7i0jGf2qmgCvWuD+rXLhTtlWAZZ
uamA7lA641gO52NKj9he1+Iaj7vwHd///DeixBacWit10qvkIChejmxhRo3z0Aym
qYJeyuST/tDpt0TViQ00u/NThtv9e9J4yC2+0IS9z5M0kXK4yyHEmUL2tTll00Tx
UsKgtB5OqvYIIkAh27AUfnWZJ4L+ojED8QG+k+7KHJ2AvdKcRt95h7zwf4PpTlcL
VZUkDl3rjbJ1pVU+K25zdH+q5833OD+IG6a5Ixq1RUR+FVFCpvCii83n1xfFowcO
ks61/HLCFJf20k8dnotXC7ADBH2zVWdiKzENW7yZhH29RG3ogwlbjnyIgmNCJle2
GAiQZOHKqYr1btybWnqmDQut2B1/sezqs0GwjU/o+FuqESDwF5t6evgk4twHj8J4
sNo6V0xtqAp0276PIg2Bqf2kTXdUxBfH+PD8ocZN3l72O7hr/oA00mZk13Pzyhjr
8+YOuJKBF9RSQ6wRzYZSj13fz+3MfCt6lpmdpAcodJ/lRBrmaaBraeudVCZNQHdq
Pd3+MGLYcVXNXDvtwvpjqaPDpjYtL4tElfZyd3t9dhEWaQciC19N1LigZ3tO/QVv
XHKnRVmNGRfQFxl+KaPue/FzV3kEVc2JaMsKiMXoULhdNsWo2ITca12Nnu28NpgF
KVltzzeHjW4t3K5rG7IWTKNf7qF5jkwMwek0lhN75yAV8gpYNylA49FTSwsvVjhM
L1Ne9fXustQFF/HvCJN7bgEpJ5wiTDVkE6SbZsXaWwcK6uvvMpkoNTABJBH0bV/B
OhbbnraTFE62wxaKw+0tG0E8rMjm4bUxQfoGK7OElxP6juAFKHmYY6q/b7zskeWe
lUBOTON4jfUTwHzLnpfeF6GzQ8FMZDFjLWtsnzOxaoguQiQiNEdNC6DnOsEfC9S5
cX2ToDDrxvjznBSoyrsrO5SR9n96URs44KiTiFgQwtsmVP7+dPvlF77m751HYGoo
t5Tc+HCnybaNh5e8zh0e1hqsBRQIH6TkS3FIaCsssAlh5BtGpILHI3MkFE75faIj
bqDDh60NuTxCr+Kfj68DHZ1y0XZhLrEQsSgFalSjjBYmlc/4ornLpbgbki4t5XQ5
tK2QAFjZwXXNag4PvwtKP6A21WVNT4o1kVOXOOQWAJiZbl5J6HiLSYpD90iMPfCW
ddIFGZrl9D9ldSX2+1SiX4xDEhSQEzWKIWquJ0t4fMGiudLbPotecMMiZfxgMk5u
wcoeisZSgvbSG0gfFt9nCZeNG+BxQCrzmuAVWFQWEl7unxaAIwzi5lgnYsYZ7WO1
I3hD5dyamEGvW7UghfXDZUGAR7Hf6Wdp9v1lya4EYclWU/Nv5x97700ih/xAJIgD
vpox0cCuIQvNb13NUDUL5Wufw0oMXY90oRNpsjyTmrmCWYD024Ij8TQ8vEQv7aBJ
ICo3oxxF6xrq6tunsB/GgSXRVOjQXREBzQ2yQlm07BIhATNdrGIeYGAtI00SS6Y5
BayRR1sys3dwIqKmCRINB79xRNhQ2uy4Ei+GEu9MHidf6buv606g0BCR5Bp8GHDb
hjPTUkNe9vxPIHPZKb1MpYh8Lq0si4nBIkaaO4usct/cVciTi7WwSJ1VqzMqwMKo
fwcQjZHvma9RavgG4XI1pAbnZozx03F5N2+qowsqg+RE0UlwDJl1GYI2Yye/Z8w2
KCbemLDUs0hVYIn2QaXkaLDXFB4xb/0pvVYNQofxMLtGFeBOAj0LDH5t4sVmF/8W
yabkZavodjbUGITVcyqzIlBL86N3oLQXqD1lRQdt/iubhujjScjhg54yShpcL5Mf
/5qn4ZbH7kaG/Cb1jvjMPJmjjGAKaS6g4tIAtly+23tIa7qRubD4L+XM0TvLt6Sb
K2EuCzpT1gOB7KfAFvAiaoSBQ4ww4srMR546MsIYn6hb3XHnRQ0T6Q7fOWgUwlxN
vdryMrzmk0xLMief3BMw8v5IvwOeLTW8Z17PdWLgur540LsvYUiVxITJ+5pYwa3i
QIPF7xcZALrBypAzpOM65ZEF14kv7oYnxwJqmWbisspunt/f3BjA8EH1Kz6dEw2s
aIFtqsGYXl0niEHPNMwNR3+gBhP06nSnm2ERNhrqreeJYspM+fDJAGG60CV+ITh6
rnAmWfvk/puJj3Ltl1WgeMcVV/5VDxmoYluaJ2XM+q8oo4c7ek/+LfVSmgHojwd5
ny/iEhdD0l0HfLtH0r5yR8mfazpY1Ko2MzdjIqGOQhQGK00X/NPTbhaUFA2hlmDC
oOg31UxAR+3neNtS4zuIUj14gXUVeQANg4A/sl+5/jh4Az9GsukiLAF0Yosr+KC2
YC/5kvHNbVug81f/cdUaiXXNFg4/EE0d+LNGJtgf2FlEzv1XDymAoNJzhAZ8q7n+
phCx4xj3KMCjwRaF8pa3voODsN4JtunTSA2GATvCrfBs67875d8uJdXMqQANKDCF
EYRa74D1t9+Qpz+hY+KD5OcfQMbt0xqLQEe0QYh/vnK50wroFolqE8DLHbokM1xq
KgofSMRqdDXKYUIuopGqUJ+Y6JsET7XMtllwCZ6vewfbUQsmzo9OWquIFT58fWp2
KTqu6PVOVKnafUybuYqx+1Z5ME7gS6UTSVeYX1q9Iyqomeq2uqV2HTfw7/eT+f8d
c4hP35yVouBU65tpsiQ7LP9oqnTBDtYSmxPm6K9hoOjmheZH3LEMe0mTP3Pm9ESD
B+XjBpjCPlB3Aek4sQt/8/Y6NGfwusLxC+OuCBSuHn6HDLdzSUs33nFeNwq6iDVJ
g4VN/qXStrtMRCL2tqGcAEA/dst1SSu/m2tZHROPhjq0SoyfBE+qA4PyrviAOR40
MQELywVqS6k+bCR2aSmL7E35PLtmzWDdunIMSobBYPhS+iMVkgi3+mRRGzIsme13
I19++WZOcyd95H5+r6hejn5J8LPNpUZ8ONMo1sDg2Q1bIQeCRTF94MSPJVbmPVrd
556mg+MUFRIvlNTFkvIuzzICT13Hf84bWjhwwY0KLEfas67ewlyuEwjJMIeS+Yex
QdUK/KVVrkca3JArTeydR/jdWhp9FLP/0POhD37IxWLruVpCLhUKdkYssnHmi7oL
lnGSacfClYAwXzAkW+gFBF9sy6/sFZKHFSd5OqTbLj86oXGnaOeUDNr/pSD7lkVB
ra8dSZbscPH3ZdYDCZGEPZ3KwXlaZqx/GvirBAwVLLq/SLbQeXsbiYB1O+QT5hgW
Z349QhmrfO6UdIf/EbBU/xHgz5Ch5UDIMMhS4VOOwX5pu8srud6r0r1MSEmlkQhx
m6PQlazbxmgoE/jzrrhI+DUcygPwamrCpJzh20N1lacgAURy7uasQ4dFLta3+Pu3
KSewvcfxujlFFx5IpX69/9eFUlQc9ldn2nerD92SthAfIW0gbW8CMuctf7myfxV/
ZoORl5mjVLPtfQuM/2BBWy9EYLtwzCb/v4SXCMxPxjyw0u0265XfxGyo9rQqCtWz
zWh/0KnQ0Nm/b6a8uaInl3MN+1kl5y91ytF1Ts6lKQLid2BuyWFJKehxORXhsP4Y
hJVeUdPSvDWwI9YuDtthTKfovWYH2QpTixHgxcjctMjtudB3ZaYoTwqzwQi1Y82o
Rh8XeifzAV0n730G7b2aVFstM3TkzVhHKdFDRMbP7YQhoMNq6ym5lyYbOKk3iNpY
suvxHfVd3gMo3DEn7zrB1Fs04+KEOVHnO2u/m2VQreKbHNvp+bamNi3jHQO8icwr
op38k8D5wCJPIZ1QNLzsW4YRoCGYq73CJvpvVRGsI2JRHHpSMHatEp5RWMHgTW0Q
ggKBHhtRhbrusJnhDvzM1o41t3ZN6ecLarHeJscKhPPg/TP6v5+ifgbJWmx+jlBR
zJ0cCk+tWYekh3DDgaiL3jyWdTLSpFJxUUr5mvtq67pjYD+f1pRjBo6XaH+eMggv
i+1k4jeNfKEvxDg59rMAUdWI3illtrsRWwg6mw/zqjdEOXLbgO5Brc1NSm0R3EQ4
KSWXE8LSwFcmhGCDczyKfL3RRwqpAjxUj0P/fdxzHMVJ7mYaKYT5sbx7qePVgEt4
KCP4BXuktJnrF+UY9GKugtn8GWtuy5LbpTHrOLoT4uE+jlA2wZpVa9R8aN9OA7C8
sZgRp2apELZLeaeAC8C/H9VVeU4BzSiira2hxGPUrj0qfOAbMT2lyknzTpZ2oDyC
vMDihaBA9AuCI5Zv9bOWVFy8qCXKs8mw78LoTu6HIBRCk+LCP8PvEq5VO45vaV9v
O/5srEdaduFugVaV8J1avEu3ZWO01A/vJ1hXwGcvHjJVsg/72eVQqduK7gPhG+T/
ymI3Dipey1/nRCS9QdEBp1eAvC7mNBiW3WgznsCjPIvWS5VVNpjqznHvAG3essuN
pp1quzqueVqRXuVd8+tT8BICtYQEf530ODZ8wzgvT1dfd8BSbWuJIYVtIPxhMrhz
NNBZRdbAjsGyR/akwBy2y8XFSBdM5fk29zL9kgV1WZe7EPg9RsOCTQZq5uTRsBCr
FW0qF8GIsxT1tiiQfwDID8UDp0JJvkLN4UzD2RgYI3DsPmJ54vvZ+lkpss+YXUXm
Sb/C18ATzbtj4wiLjkUKyHg0OtptZnzXkPdbV3DzRuS4cQqISBGBk4iGpq+ySzdi
ZcRLUQlFtqnbSx8quqAj4P++8X3RlfYQVbhmiclbQ/CH5vW9bMky/AEnvpbF+Um1
Gk24izWbbRy9lXaS9H7tVDp5y/HWBUUJ8LmfUOMkvQ7I1AhR3pYTr8r6OJ3r5osZ
7n0ysi6MBG/iRiXytnaGPC3vdTKUT+shyLli4pUZwi58nHhQbITDhrbhGq4hft9g
2iW54KlvyDECII3c+dQWn+KzFlE+XKceOYlaSoIQ74Bgx210ZoxZD1y4re/X3XNF
jxtrLlKQ2lEPRNqtTVZ8JFTP92bBekHCPtrwIzHCW3S/8oIax6Oj/KuTgJWN7Cu9
7DxlvwqvvkJ48zRuHWnQ3KDQrS9OiEFuFkxX15uC8O9CPvfETFbuzTO8BsIOFLgx
7z5YGhbBiGpC/ngCCpHWTN0tL5TAkTmnaIWHCjGcC74EO6AiJWKKLJuD4iuBt1on
4ueEvP1Fl5xFDUTpmqasBxltZEA+tdVGKpFPiy01k9Hx6FGt2hXNxzr5nJkjui4v
iA+iMRWjcD0aQtABi7jVhmyft3FU9tUfiekPMS4LzL/+cUcGnXklM5SnZb/cSrcY
xKaVxJe6Wo2fIoSXS3VyjMuxUA9/AJESMLe8hL+I2Ed6eaCmwYnpJdA3jXx5g052
DmeN9GMl8vUcvKdvLdoblsmYW07fr6gB1w+hynK8ahAPpwRXPsbjU8D4/TK6KBtx
AWCtYP0IRy6Oj/3KBhh7KTHrGuepY9xKCkNgAQ3kh4MMl1m74ZFwhCjcJ70MigM8
TEtffkzCnozjdVKUqT0wP87UC5dFOt9MLNSLqoJe1s/+r8+8GFoufLR7ImbA/Xvg
NLfp4NEwTBemPHIaf2rW9HrJIQeLvGo9MX/ULg2lJ/xTCJ0bk1Wf8jx/f2gXR7tL
UChxvpytXxR/DN5uxYs9nsAjyuPFbMHIsOWb9RuJYzQAIYaTghz6fksy1sWloXrY
pZJ73eDFJDftPnjyEt0VTCgRfn7LxH913fv22tDST8Jmdysas76WPXqYHMjkawKg
cjLox+ZZm1xZg5H3Fklh6PQuGHwjky5SoJwaX3yZZjf9COkoV++1hunTIoAWnkS2
1yagkCGn6vQK8jndtsjwNdpSeb4emZ1G2Az6Wub4tEnD7qhV7Ez7hSWE+CLbSHXI
NAf+AO54M+ZkHjVtYI3+YO5AX+i1e6QyLJau9oj8mRPivUiFQrbdXm6RzBdQqvuW
Py/omlKZZuDZrJWDtkSEqOAkAF+cF+QiLreLvcQz6G2xFJjdxUqDWgod0W72Pspe
/JR4WfuaQUxS/zEith2TCiUbLcbKIvmMBKyDybNB8b62PAzxcJE/jBTnipH+/ipd
bsIu2qB24k9gkGr0dY5X07EtVpS7w+ohn1ZOjW4SeRl0sgz/6nDhH9NiPxXzz8kW
BQfmdLZAGx0bNOHzQxwzRgK0v7KkO1WMRbAGaRseWjcgEQYXn9/xHsrV0WTmcgUw
yD0fLQ5ltNroqMcO6T7tGnXJSmlRVupwUy3Me3W+W9nv6pDn3QbKIB6aXTGzxPLp
eUHm0U9aoIXPVgDZV6TBXLjniW/APMPuHzFqJqhQFlTQWjVl+Y2EK8VCi4W9DMoZ
echALkZIKK7N/9FiEYY7WCPTQ7/eeRaEmG5rZyu/D5FmbEfY858nuYz3Ahd6Gj8D
0U2SRxWEZvN8EflfMrADOQBRhMceWZuRCwG0Z7/rdOwsIjdeNCSa3R3F1k8HoI8+
wvHcFfMxwuA1/OG3sI9TXxAlI7CrIFNyRF0bbIyIpvapOXyqeDZrrJ325pkQOazh
TmL64z35h9EyI2QfjTKWREkUVb6oW/RJIc8gHsDFJgwSRnZ1aXtcHbhsETUXsvu/
oXZSdRS034enGKhZOJqusr3mUmURKzl4P1061Ooa40aVs6fOej3+c0RSKfZaJXLK
cMUlSdePLBIad1obUVFYyHSqeD89yTDVDdsC3i6r+uRI20G+SeLlNejk/hSadFhK
pu0dtY/3cZgeZ+bfF8GdDXVnrZF1KblTZY+BSIOWg3hCzT4XupFn5sx+02qFya9A
153Ud3owL88mvs9IdWyVtClUb0gz+UpxL5M0ywHEt3ZvlKGcgi0QTYxDyF/Gtybg
4ghJ8ty6pHpIfmccRMEQQO4pxWfz7afUfgQ0VQEaoJozzgzFV5I866ptPzRTaHHQ
P4R7a08SM7/+oYDrWrpSV0fKlSwAaVZkuy0QcY2y1klVR6V7dxTfjs1YSyG08+t4
XP28/lAxmS1bLm7c0ihOdCHeaXKbt6vSh0UgpuLS5qE5qNY2zjB9twmT3xFqsVv3
HKaFGk43/jRTBDsK+RBZM3B/whUHM0yM4YYZyYSPZZwRqvXTYPxLPyugQlf0PsKM
lO6UdN4BJn2ydQjV/XfNSNGFNVqE51tG9rgO5I0bi6ZmJ8QvK9QVsaEbFDnidwM2
y3NW7nB6aKME9afABW0A/2muvrhxGWhRmpbqyvdTIxABkYjF6SVTQzBfkEgxqSXz
UDwYOrUDjJCFDpPCWIt7JXP2KhoHCUlvjXWKQ2T8m3JeVutKUtFhDrabq5bjjFN9
/uCX+Li1ZA/9neC158OopZ+FdeglQssp+i7UX1iUpz5pSDayf7rZtyyhfSir/8Oa
UhLNRu1P6RyikQ+zWQBf5NfXLYPys8SueZAabopfY01r8yycNc+UhqJ5aOR4Fzvv
k0CG5Cd6vTnJn2XgkK5kWO1hujXDLCQw9isSOZSg5UqWUKLknd/5WedCXY/ZKfvK
gTiTjl34DbCgF5rzDhCZBinR5tMfW0ENvDTUvbqrCf52d3FDlJtWkbYCROGK3Xre
ijGYkCxs3Uz80EaTu3UPAdRruz2z4gpm/fFNJ2ZpTZrDSbDDoqyuTMPfHn4RgSbt
mulLi+dwFedFdjmsONn8CgYssQBnLaO9Hn3Bc9JCu35BCydPJ2YsYZRr2/NfiZ0Y
dF+Wcn63HO7CsPveSFoBAtyx97YeevHYNujPkLzJiynye/9mv2Yn0oOVekuF2g5S
d4fjEkB55NqWbHv68UUmSPLEAyXCnSmEkOjVMIG1Cm6nzyqLZb3s8n8uQRg0ISej
dq278lq/ZL5bH3zBN2B1C/sFwPgmQNz9+D54L75j5gKNz1nBG+llvzD2RuoSn+Ay
m0hreu4h/qXGIwR8xb1ryzG/BrUXpxmMfn4NehoAN+pSJnaUvHVRTwxYo3PFFqjA
Y2ktxyYlyYAqpLmBVAuKXsA6G8pah3uLzOZ/eKF3vNTJGX+Kqi2GGZM0fz5/HeaE
NlndcveXxl7dBCoOHqj0aczgct5st3E9B5U6kA454isz2XrVDNVtxHEV3iUVgFHt
b4ZyVZWguy4MTLzRWyp3OT3F5a9ehhhGLmHab1M6jSCRrhLrrPWvocudg2TsXdve
PGhpBXd6rJk/iFgndHE819RtP34LWwZoeWKxhweq+3C/2PKei44qmR3V56VY0086
3h8F8t1FLqu2ZFJ9ag8wwjTR5iKhoY608LQWTDFG/O1NiTUlLOiyxI5GpdamIFRk
B2RrljmyBdB1IvnqmgYvOii+4DpYtA8E/15Ct8+4bi3TE+BiQvejboxvO/GeWYTZ
jiqOt7gWyJYC3y+qOkMSCI/pyxoHLhNDrlMfDUk22MEoy1LXix+SrlMoAviIF5ND
Tvbdj6YXk3hna+MzHY9u7XhxkuyPH0YiyvPzOuUnh5KxsUi+iPt2DizFeQX0HWvH
UiHA5x0oielvOW6TwSIeDIQsaOSNIAvg2N32q1YN5+dc8gCEr0fELIer+eFjei04
UTd4AQFhHilXI/UZG/YlS+pB3CF3Q1dAVgzFEVddBvkBRap+xh8v6YwzH3v8DZh1
6VklvF3YLrz6/rqndPmrp/QB0NL1ZQqIinNHGAfndXRTqhpikLB7kYEMAPBMjgHr
SA9ug8uECN1zoYegIBr9J4CqayGqvaMtOnWzKZA63rs8jdzZ/Zeer9q+MmcgMtUv
VJ24DHFg5AqkTvULMdvtF9Z7fHiiGiP8wtv+rdHIZe8G7h2FMTdTaQoIQuiNA1Ir
lkI9EUnJp4F0ISE33QlrX6P2yLGRVJFmHGptUyrLvCFPiK8qKMNih09Su7USeiQN
b3P9boKV7c3ayUeWqR0av26rbEnPm9E4VKKQ0JF9aTu5cEGhabevhPUiABeOLqtG
n8NeFOW0sCOhqe7PDLpD/dl/s9rDRJw/uekyy9HFldVWtmvwD3y/JW4nbEoQbkbt
mtNVQR4EFhaB8EJEM5xCOYXZp6hfgHhHms4fIrHYvHFoi3WNvIGi2BsdlBMlRytv
kZEIHFNmY4aNaK5rJnmTdKZc1qW3Btf/RxExjVABsOffYftTeag6JlGxQpAptOgx
1fpnsKSO8M7A3DEXxMxMRbJmmoV0Bfg5/W8tv1aLisgxKBRYp9FXZLYRRHsoJHZc
1C/kPNIjcVR2aTV4sp6oBs+ypX+mcsNj+w417MqL5xZrnd+SQkZGe4MwXNLa/8vn
BKIr3oxZRfd5zGcrD3BiDjlcDXPlnZahvPxS79slxFeQfc8puQ1RHDAnWzQGlvDq
aPOzW64FSTa3kc79C+0+tNvikjLWCrajOoSNFczcDXl+JfSr0F0uumdnduIN6oAP
d4oJPGVEv0bbqhOFSFDrAEaxHPcooYrmAURw/KXo7gn7Tdjvm3AnL6GSNazMNDAN
WOG+4VIAX94v49rQhEMKMgdJGdnh9mSFJ/CBooDZv+qT5PoG57Z+HNpW1ZrbjdMx
1cUrBr2f3aGGVk1NV7Ldo7HHNCKcbgQed4ag1mblVbmRmlwimw1Rspng3aOJjJl7
NxfBj41PISM/M+IgYbF53/K9LcLGdrvAPzjDaQwFUNmU3sGf8AAq9bLQQsDEljcW
h7LSHKIYnbkgEN99hW5JNWE5CoOk3kAog+/AfIyLQb/0okugPFa3xgNoIaX3tPb4
zLuQvb1qAmE/Gj0oXD8WjuIlE4mySzgfS/BZdpxW/7AgeGKfXnX3IXsOS9spIYrJ
xtkhrILgpBHWVChrvTVtvYnnD9wztSJZ9JqCfmv5cWQeDHEh5wdnykDHUL1lPXNL
ZvQS/035SmE0Wp5zfeVRA1pnjb6MtwAKpLrmhbSlojwD1zFgIqRM0RhNI1i1tfA7
Fxui3Dq4zH976TLZ2l7pWbIbyYubYuAMUaOF6MmWTms+WpaBD7FaNYkTZ8GHi3K3
1TwN/unYQ3ej4aMhJh6paPlD08jLTggBKDp8uk6Z1WjjFKh9QfCQNXmZX7ZcxCOb
pmmjWYBmvW/5MHQpYAluYmP5xQdJFQ5nDoxWnXItn7652tBGL1jXrBG5KQ7uKSAg
isrBr4SF/mwGbPeayVnKYsUXF23xs014IrmFE/UbWVCDo12Hl19wJz4CcRDOOXHw
MMPb2F6g1lRPxuyH4l+6w8q9wZcibwhFt+N5T5gVCqRsi2vZ219wI7KSKb4vLA65
IGGXbL9ssEOgCARI8Nv8u9oDT517e+Uc6zbeAprdEt/tZxFY7fm7R7SDaGhArl2n
1nY1WJd65t7IWJQTlMlEr4qUeRIl/FC1wMgE8mtMBgrKkiiB4JY6Q3Oc4qdCATyJ
4rczLoFg6wpu4uk84AUFgiJjLaW1Rd9H0DX28ZKcOc+BGb64AECuhDNeKA5WIygv
HuL8+RqFWxQNlW227jr2YKBfs2qlhX7tuVWmvz9OqxGNT6wbVWoyabVK14KytBhx
e18o5zFBml+dI1zaIkwTpWFUzE0ywqo95jTkjYYKzu4qZ5JGTTqoAn+7xNB5ZdGy
3rv9EJndsgxuG0I8+UygFLZ9v2rI+UXd3NIibAY197fwi0hwlSk4xWsPhQhtDNop
m2w3GvkxKaFnvrU+X3NqoHAfPn93fPhGyCAYPgRPeqwNwH4Y2gtQvGWcY7qbvmiQ
nNO1ImfMwZBZXyR8uSLX4iwn/AS6A3aXVXo2qgC9Xu6VUlRO0DGsPSTotDJdixhB
2HIbTHZh51MCK2Ci3KnMK6ZRi+saLcpYR9xiTweHRSKzS7dp+uxsEQrbl/8Mm8xz
yt8ULsO3/4KAffEOh54ZCOQ4QMqL0sOTavLqa5OtbRRstoZ7qIftTyRUFaDGoKqZ
tZVJ7CRHcBtLPFCiatb2ZS416zA2NIleSKJ5zJbl/awBR0nqcWudfB3c8u2ktreW
HmCBYuePmEMhBLUv3UQzw8Em52AZCooWvOXwr1VLuNI92Owg7HsW1ioS7IsS6aZt
8Jc8P3016iGf1cKbt2q5ejwdq6tRrKinb8CLTfvm96iLNmvLuFgMLYLQHK302sNA
EdMftL3u3srAVB0NhtD44gAxntdNGvf/cQxYfAK6dlJi6SPWL0YGFKzK1ZQt2vqE
DhCd7WZpx3yuHm4+BccUICvbz2sWc59SS3R3VI+AAgRAQkDE9Eyq1gFJW5GYBmbs
T5heoGRruNJExGf2x3I95wXT6+huqRrwd0lu+28mhIOajBxck0rZWb/SNXJUDD0G
g3MCWuaMSL589W79Qbo2dNRa0JNDcdlHDtQPi9D0FX64jFPVamVMr11t1TiA3Z8c
Yargf0S2cLmcgvVY0jKqOknruYnhcTN5kY7c3lcfMqBnOpfBSOJ1SJvvyBm0NTIv
rgSWJo/6DqIArVj80vpzh4WgznbgONhwCdZDyDuPHMWtTDTgRe86oEFmKCOWOuVJ
Dl3uEQYqm04CCbvgDQkUDjHWMlcaB7ZeDKoOwaLsADperCJf9pjtUPxmc3tqQ0q1
1gpIBowOOXZWFZaCiMdM2g2W3T4gjPPqDBaU6X/1iwf6r+EuSoe0F0xf8JFQdCcg
iFEFYNWJmX+ZDrfXVdi0ASEDZ4Gh3OxmQcWYbDnX2cE41s6Uf8rzWkb+Lrh1/QoA
RSKNGPaBG5UwbaMw8w+u+/pYVu3Uu0ReWfNT4pynAqt/Jer+Y74qWSm3Zvu+7s6B
P41vVr+ofz+MNKklPx0gTmNmCgXffivEFkoITTkrP3+gLypWlJpurUdqCJpDggCw
r6pc8CzVQD6Qus2sd2CPyPk+ywQNbftgh+5kSfDcHsOPF76laR6xcphhVpYiNnqs
E2xUT9piSfJMl5Y0pbz2rrDdipQzrPc6bEw5nm9CCgg2cUNGlvQsNln1ju2CxyPC
tyh8ggs/ojmWvggvCiGIw0EGltep2lCtZYBvfOZiYfFFzL2lHySAW1xC5d/sPr+J
Tzr6goR0QFf4WU4PzbBXL61b61Jz1ydVX85bQmShaJm6eihAPZajft51F6YhMxRh
jdqRwwcCG79gnC1+w6BqL2Y56vP6QSmj5qXzo01drkiKN5EPq9ioqnkmu4kOijjE
mbo6LbdSOdmN77/vCPX2arFay682QO0cAnwk+h0i8NdIRZi7/GnUITJ6OTP0hbFo
RXtaK0FQ4/kKBuvhybjDTyuyLY+A45rC2NO6Jt8VVxMGaCj6AUI2n54KLnWHLSRa
SWIHkLkxcPM2I4KNPdxjIcfCB3msYM9I1GjksVDw39lDLLx5aORY7WnIIPFIq1hX
33LdD/14JW/sJUSYjWwLxRnOIXMjILVufwiCM7GkCg9WkncYLVwK+yGL93yHR7/d
9ZiYJ39U4WjpXcbPvmzMCINr12gfG5+2h7FYh3bJDoZtQpQY/vLfH1Lgp3fp1Sja
pyLZussl3YgnH2WLY0AtDAf7AkSOnjP7WC02u58hdyCRn6KKOihgLo0dqWpRnEd6
/TJh4G6jHETxM8YYcQ3cithm6fZIOyCJuwS8/xEYywfrk2+VoFHXXKBLDTpOSXnp
SOjwGgxNALoPcyD5X2tTSnWTNdeSJS6xgEmOvYo+u+ITXSWo+r95Swl9ioploQ8Z
SH2rQaSa7r4aDC7VlSulCZo3YF9N6fO+RcIXwj8FaNI4k1BJgT/acxpfEdEHUO5A
vgkFUwT65aICLS8ntBDYr2EGFNDPirFylqRdfCaYiA6iYRUw/f8MdgCr9sB6FEFd
VtajrsdeHwnpBQHi3gcvCPYLGHT2l4fo0jbWQl9qUFz0BXefBsdyXXpATneYJbui
Lg1Vc9DIGxXAiizuTDQo08421zw4gHPmkZrSPkHwUl4z6jg+z4m/KHVBpvBs7BCL
zUve2+EE4Yoc7rbGCKjPdw2i2CM6Zuwf5ps9SS/ugLmyu4W6inGIokP/8d8O+PEc
V23sjlBD63ELuyNw2h/N68khqddoziHS1+3cGjPUPOkJYE5Hs6QWjoRxpsOJ/Is8
vvsj4xXYx16zvtUKFhE3x7gMcDPz9DaRagSy6BqGsFLfeAt5/TCzEy6y1h2CIxtJ
Yw8Zrd9Puc7uWp76nsDiqeJng4SvNCyERUjLf1TIfRZujE4gh+o4nCBKISw683i6
E+kYlVTFSCLQZivqQdz0aX0eo7LY+YhX5Eo5N7ywqwIYEVu9uEPUwFnr9yDZx5cM
ff/DyHVglcv+ngQO58pyWA3UXJ/65EZy1AycTDpNcg59g39SKlrvRDUnirstZpbN
n0iBoszubDv1vPezjLoy42XY7YPbopVz5QFMSFFGhcPcBEq87CvQ3S8GFPaLly06
IUH9pXe6aQcwD8zT9D5mzHPYIImkT8AeZ8npgoEM5vYPMPKeDygekhY7aCPVs3xX
1kJBGRaUnVDV2hzKgmQdRnFW8g6r0Env6xaCQqStBj2WP98i9mSXlI/fWBN19V28
7iANvuPwpwYXyvP4EjzWBR2HVVlpCSFBVw0bi5dMh0+oG+nuKs8Vx973DkKEnCPA
36ELrH6+CoM/XUkR6gFK6nQNZAiweDWohGIAzLXYcT8a0qbN1Non00gvwEho8T7C
YKO9WnmAGSQizG0b1pRqsh2dmhlb2Xls+dZAuUCjMukP4tXv5XhZrqKL6rV7JjZG
NcQ6Bm58I+okejU+mntnR3RoTWR4v7Pmtu82vYh6irwZv3SWnX1RvsgZeOyC1iCW
vI1SKi4VFPPK3n7nhskEEl13GEZ3qyOtN1+zcQetmoGC9LZpxNujG2icIE7cNaJj
1kyR4KdkXCeEj46H9Pl9blPvMVWzhpRFJ4ziyPvl70z8PmX0ZWuZSpvxtXNNRMQe
Jl4FCpg3xm16wAVwKDAjH2+1bs2yyFQUrG+e2lMN/NO7j0//8++m7kAhZqKSPTXg
m6+OBV0NcuuxakIURllz3cQKdqkTp9eWqPuIDVhr2TBgLDIlCYMNo2jdOOxkKsA/
qgUhw60+gdpcdPETlP8zYARWNzc6ndMF8ZLSo19X9i584cNaBff72iMoSPEtS4CU
1BicG39VpyS/sA3T/f4jAf9R8JGEUvPnp5jqj69UvgtpWzYSi96wG4rEhI54PsWe
2XT+qXsKyQUfTkQiVnC0AxCJKLan7VWNAPJ4GE7/Vp/QARXzPMIaIUzTCN5lON7R
ls5H6GMPBv907ZquUcHnAIyGTMJERz16kDT5Jq25Vixo7R/6ZwIrl1b2fvyZVgXX
32Re7AyxlyZgH5besG9bkJSpLmuZGdnpokGpj765phQGGPfFk6SMcCf/6ysg/WW/
XwxvQzrroYAYBtUdRzOXdIjB+dL/7T9otNAOjJHPAuHzNh3B2iIuBfaESqX1Db+m
fOicwWOX/0kiio/fWXlZkndsUcGU/2bhwtjbTQjjGkP/3fkrTxUw3MPzxZrzSkaL
TxDbLpojdQLeKNisM8mUrq37HVcUNCT7GsJHfhFV8PhbIRmGVbTSxWUABbFY9uWF
kDIYKi4xXXdQj2p5iYiA8QK8f13F9/cSF+nN4/8ErxTcTWiQK808JuC4QJPDCbK5
DkG3TEGwfzIp51GZG3XoKtj5nO68E59NrPAWPP+MGHTNcuvqXXzhXNTcbUdPnHs+
7hjn0TmRdrzdvmJgSV5mw9x8c5STrikSnGyVuJmp98JfiLa4vigTcZzMHou3kx+o
BBWm5aFrppE+eZl7ccZExE8OS63DaEzXtZaAkwx9eYWj/MMguBABkHx4wENKfAnP
Oq9PoNRy+ydkUH827jZsJj/WWR17qWypgiqM16KVkB8I3/dfebjBsMGW3TxkD6tA
JcbFd+Paz8eVGk2Imv34moZmOPjYjMgNpOHyO8cIwNcW6rRv0vxgvEm9fgsOb41Z
vdfIksLPpXZ55dZ+coAiKS2KJyrJZiKCN8g+/DnnB5LSBUwlVHFMAdvpvQUb4HXy
A/kw5JRpG+Ia8woKAf8ZN3L7C9BLI9MiKkOvVvhDepwhOYblDSNaZfT53OQew1op
DhNbuwiIrF/hQN/46NcN1I39NYKf7RbtAerW1bZROqGq2cB9yvQ4AlJCb1UdKvOo
jIUFgJkz+PmGOFiP/ta8xLkO2SO2L4ONchHSppFIqflqWtGJ/wFPrqPZMJnx5IjV
4ZxnCUtS+0SfgwJ9ZV2jaA8IH8meLVD5IdWyHvy+BTx50SuCbh35NpPzFC1rsUWI
/Zm6YN4c25jzBzPK/zY4+jdQU/btm1eBpZMHCeRB/EOilXKeIZ20xPN4VRFP7Y7l
CvVdHnWfAU/P7ckuXZD4lHYD1aBf6dAxmt9D5LxNFYfBbnf1MmM2lVMxhMX3wi/s
bCgHSk8aAwwUxJsuLdlpiZ4519ZcBbf35STR9369WrsFS4v3tBfSNk/nXMjdcb7R
f+jhkIXJ5D7gqQKnrhOsiLBaZjLAUajk/8pyzWpXGBgCERiCnExIIbUF0j/LwxD9
TmVD47wCo4ARjPSSZqwFqC25mrV8mbSIWs3q7gIRk7qQErFIIbl3Xb/BNQIKT0qQ
VTyTjAquTExMa0md+ZzIa7BHpEb8vo78SicWYF7ZLmAcp2/5oCWOXx/tmLmwjbOi
6sHEZeLF5NuWHsaAIKXbYnkroM9zqBoRXTrHsZiqxz73P8uziUwBPcUdkcsqKxJ4
UE/gG00m48mMlPrezd1Efby6Ao1Skfm4ftpWDOXSCVCrHFrOqWdP5JnePyZX8wxH
6UNqD3w9uSjJE8AS5mFSHKDgGecwKPr+dqHVNq3nYyPPBTAm4CmObxwvDrZx82z0
iyxWH1+h9jfF8y8B8QE1Dc0Ir7DH2W5qLgMRVRB6PLlbb2zQ8cdXIopgQi42pZ7E
D//YSKJLEsbYMFC8ny+cduaFj5+QYum826rp2gS4/UB6fFAxoQMO3XE2QICYf4jx
nZKdVlQ1kBpGxsryl1r0wmXQQsogzip3xa6keCM22adaUryYE3dlh28HrDuX5nlp
hKfFG6+oi4iDvmLmjDWzCOlKhQRjXO8isv0N+k9fK0kVd3Z4c2SGZaxK6aGGmDNM
FqSBTvHtDs/7BoxKgmKohGoPyEexgnkchlT8chi66eiFAl+Zqq/t24lEWt4JvQb3
JATZFedlJxgDM82OPQTgoWZXaq1MAtwASjHkRGDvfhY0CFueh4ZhssRBzgi9O/Qk
SQ9VG2ZyShzh9sT2TUYOGvCgK9Pyt9gsKEl4iHtm5qKgIHhNcRigvF6ho2kOsgR7
2T99luAg+Pp1kgWIab7TE5XuJc0Tsunu3BExl+14R/YPc2vSD2Diuj+KYkltOgCK
JsDUjNlCKMCZioKcYt+uLqpGPvWkROb9pg6zO5WSLRIHwSJIkerMhlh96tWHcTM4
l8X9FTE7NwKHJCJ2LlPw0FHIEOWb6iC4ZMjMo3hr0+p8TnJdGy7EbvQimQQNQcFq
cToiYEqRUb97+uXPwNb2iZa3Rb1mZoz88SdSoZJQr6APPorZTZxhHEW1EpAJFwwu
BT0PRUQzSiL0i6cU+bYvssKLdZnn02OOAOgaFrUcu+4nfHR/J+GKwg+1jv5palN6
XCEC1F8NCIoVd9u2YlyFjX20sSXg29+BKQq7eZC2vC2lT0DCET7m++Ks8thFCCms
YiCUJFsbS1JliXRRtx6tr/NeRzy9MJKEmxcPiIzF0k3MhKLh+sMkHZHtaaiaPCRs
9/3rGRnKJ+lsCj9zSoFtEybcsbT6GkUBOqjUWido1bkzuP+FyE2wsTXy+LHvl4D/
MRyn4o2P0nyKBBTz1wVSeX1A0geTCuUmNda/pp/WlXWkwFXWwdCeMSZAHw8LLMq2
Uqs3U+WMBboOrQpUQgNIfzrJPFgTNV8fM2svQjN440mMGqm/zT3OGSHt/Ha/kIE8
VXpvb+TqCYMBz6JjGRyVpuOvtz8Ina6WkjKcnQVVgLGio2o33++mxkflpvOLo4cd
sY7HtIZcAkybjMBMxxJz8lTPzivrR164bleKR6AonbvpsmXf98J6md9JPS0DT4fL
owfmIPcYIkzxa7f/5FA4OLMvjPScFSQboQ+n9wyCX6Cqz1jJgMgvaiMdND3bV7x6
eddWqiLvLrRMrLpQbgEF9iMUGROs+L4F8pmzLhlaHu8Xy+avMhHeT0wrhxpQkyfT
mHPc6lD7WEvNeQvtepAI6BLOuDu3vU8+kzLZ6Dml51FBJdi3fiLddsFOH26Peg7o
I0pNxTghYUwqjzm6yMGaNGkocifLhXT4k6v8UOGLk0mFFheGNcAJNkh3DoI+ucEi
FzOOm9Q5d1kMs88CbFopXhnImIxu+wDz3BCv6MNB7v+dsG2liUeT5L9K78aoosoh
NWkFz6wwlh3KWEeZmsAIbzJk3TPKb7mEC5vYqwZg1+b6r5CFgq/mY3HFzVSQDyxb
+RYI6Q65d4wwtFrdN+ZJ+6LGG6lg6sWEGFnMmDga6fD7Mbxb8ViFDuJA6XNdw200
AIjrhQ5rGYDFqYIWOrYaHDyjsSMDC31L3x0qhv7lAiwLwa7mB7e1rnbNM60EyJT3
u3N9kz69QY2WhdOuGMsBw609hE/X/2FG/ifWjoH4z07GVsllPT0ai46pyenybYfA
qFsKu1vg7Fd8R9dd1EvnkggPLIkzx/O+uYqhnKswU+NpVO+AK5jHMZP/6rDR0+DW
VCELIIcIYOTmgLnRdsFwiPvIifBXfUbuQOvskFF8ibsalbYytuY/eEff11GgKj6l
gxRE49EBMI0qIwG7xgGb1xHZs8My2TvYMaCnNQE4U+63rrBwyAf9F0CkU6MBrK0A
QpHgaJ9gIeOjInbZdfP1CmcqiW1BHFrn62wz88kdv8t7TxVLWCwi/7U6bcnb5gXO
6/9Jh1AwJzZloyobs77uzqyydfxscDXseT9TSeWGy8o7dyeY3PvIPPhxotPgT3A5
gHm2jZ7Ksk3+6vGuRtgjw5R73ZmjOg4Pwd+P5fl6wIVmWWe028L5FNZUAwGf3QJD
Vyg1BSSQcE/JBvKgmKEZL9PCESltELIok2s2ox/GL4Iy8w1I4HciNxsASoSmgNJN
W0mJxHBk6+xmGUShJ1O9/zkaAXjvjFC48hnoUlvLvzeJuDVrKV6FycoKHlgMjB4d
pF2V5aRnOJUEsMYp/h9jRowXeZfA7vr9R68ZAdtl+JGtVFIYAXHpsehwE5/NK74K
VY6cShdgjlJpIHdV5NAscCB8z1YwcYE0sd8eWpbV7apnCt+snp8VhdfKTsRWDHuP
I/IVVBFduuk3k6RVOThTQQrcPxV0mouMBVnhUdg/0BO9aX17kQNGGTsG9Bm3sB4u
irrTeqDU78TepKBr4vLtw2Hpg7+w+u5Kg1F1s5H3XpI2tOoJNf4IWCAG5RXwZ5S9
TTcDhrHHVTJwFE8hhI3ZQW8jw1wDaCQBr3ksQulC0OYleDItQA5fo3SyYRKB7FAq
2OkQrVwQ6G3JTYvkQIbBlW/Bu5ZX3WC8Mmo/GDCvv7JK3i5YcqJ3GBVRsvbi+LuO
OXsG69hDSUpzHQ/c3nTo5kZv/QchgKP4P9mcOCEkCRkW4ydbJNQMwGKqLLHJRDq9
KAFwKC3J+Sm9Dp117IPiOBiBC8r6ZJn2H6EHcKoBIKhJVOG6t7gjFwJgWERUt0p0
e5nHxnYXRBxTM5a1gd+je9u09NiaSjgFQbEAUXYIAQZn/tv3RrumNUnpxkcckkzn
EIHL8PPdWfldjq8SKKrmRmmRQBaU3c1FknUPUk0fQlhcTyEQSUax3qoVEc1kj4V4
ljlPDiaADhFH93L2cphPNt9GuPMeEomqRbryWliltD+nNNhk91/28N+2cyMFy9RE
8Xc2xbG5FlWiP6f245JyZVEZi/PUHn4su41Pn+3C+UAutOGtfpqU0gstxcqrlNfT
krCsrHut/dS7l8O0DhmFM4VfwPhVpgznsvzwTQ+H8mL8ypR/HjudJ7WUnd9UOjsH
WsJBZo8P51ad1ZJfAbfHXNcvf75/EYH1g4LcGGlO8bCRpjbiNJj1bgEuExZWw6ph
QSDNJKlHC9IojH+BoGbw14aeVCThhC+623cnS7+d7oIyArW9HaCBxWl+Lo2kG9hF
wLilu53CkwBbdsP/I+RFHPfuTRDWO/K+KDMImdqM7/okA2lsT3SRZcdJQdRt3tJ+
cK88pQmlVFSEup02tfqxfNjHAqiFY4jtCE8juUdOq5TvuVUw5tYck5eVGIufHGGe
sNNuTJIRP2pF6l6KJOmzWqoQgAkW9SxKdE5XMwvfGmAfPbmY5+F3MHE0/5lxeoqG
5gvwgxqyuLCU9ZOaO54AZaQxrnCr9sKR4vDrjkMSYys05dU+XYsmbCvKLWb7Ih7z
vheY4ri3oK/K8f31bKjKMkKA5zOHjzdsCf1H7OeB8W25lJdTWqAl2bVEOosDCZMh
tgfKJCxiqo66pcI/TIM2NLhF6EI1lmS3JzAWy7jB4O+vrZisTYGDDOM8F9Whq2DE
2cvqgQ3rI7JjCHShQWVyWVyqtSaahaZDociuMAawl3H2yL9BddVVb3XasnivkINJ
N3kgLJeJmDKSkvQd/xwBKDWRU+eHIgMxH/tHRCuaPF/M0UJmtssFep++vtdquenF
2uKqS4GfnKJHTC1eXFOjbtmqNWH+7tNuhoCz++QrQwg4EFCQJZ8ExyLozTNoHDLb
3PY2Qqnm3jEMX1Fc8pwIzIBV/NxOP5jVyoTcqSIo+Yf1kNbOOWVTxVkoCPvlQ8iA
bY1TaL8gyXdOLKJoOvcpJ0AXphVcm1zG7Zm49fE24Eoq3upUqLrMqV1/VDuQkHUo
HSyvq0/DIbhT+SsndvwpbeX6pkSHxVM3azgJsp+4+2h2GY7OE7oxFaGakd901lmp
B+Z1ZMGiqAEq72e0q4rPaeqnCKF8Zdx6JTiLTbQ6pfprjAffLx1tKcRL7l9CCov7
VQzd50CXNokPcHInwBoo8XSYetYN8PxeOTJEZdc9GzCmNhOcLSprSzNYi6kFXeFH
xaGiK1lKDTodiWO4jVTcPxwHv5pRshLe0/zbpP23aaMlOI0TmKeZlr+OUxdgYfyW
KEXiyMcnEGLJQIkIc2I1c9yEQ67g3LlSxPnvFAfi0YtnJdyZdYn/sRAvlqrua7uN
AEk2yJA8HVnBBt1wpZFBCcH1KCgz3rC6L5jiVQKNEpLd9VVM5yfXHMgph9j8MRNI
Ij3KPS5MLXXYjf5grzhPc5/hSUeInteEholKxEC+ExSCCAAeFATPJnyilKpB6SB1
KOTCK89zyrmTnVFfQ364nLxoKDSV1qmQEEQHe2vcJ4sCLQcPGrg1xCvPLaeyWB8w
MjncdVp8GOFBTkKcowHC9l8tNVOkWenTgUnpyTD4F07ZauBi4CemhcLZpWbqqCbt
olMmSI3e2SpJYsinWWFHmMJmrxiq3I6twt5J0VKHzBTW2XZ9CFRKdmGKKGlgE2ql
4kEmdUn6rY+2bLDugw/0iGKwuWxWyl7Wh7LYYvUF8hstYDyQSvzOcuBe5gTdVGzD
ffrjTagmxfc5V+0EASAsvW5mbKODAwjJxeejsWNbiFAFx4eq2TCf0ap0kDI2MYJD
PiAR+9laJgYJaeFlE+YGaUOxHaQPmLJcy3tTpbjYvxUZ/lBEow8h2qaTu5/HVyVy
a/lkcosQsiv5VVHlM1L8qhOgh2zgYj9m2/0qVpC/KbpM26s9730GVImZ025Dhuv0
KWxB41FK6+ameZr4+ZvVECRkn60u5s+0/GXtzbx9ln0q7AfhhJYTJ9yNy+5rgCAo
8Ta8JhLQrjiA4176ycm+ezLoSfJPe5A++PQ8ThqBDk7xFWyX4+n/GlgS6Rz0YYwf
4d0pQlxTybtinyKa0uKVLm5NJs/l8bgS0HkZUV1qfzC89sdvob3uhaanhZdgyUtU
zBwNbrzE0dUke+iK9DfKoyryMddC8xAZiTBPa5YUoWQoCAAr6QSxQhwLVDeCzkm0
tDQ1EwxdcTszJ8zPAMy0jirxnTgHSZ5IOqC6tlQltM+LYjJpH46gwIHZrZDlEU5c
nGdHd0Yc7JvOm6eIBytAB5Np1utAJem/mqVRq+RdTl585igHFumpi2ikuGe69i76
Y6e63ll80wke14ckEROUsM0Ch1JgEj22JQTQvHlxXCPHVjAPOeuZZiTYy6Pbi7qb
BZcYzKDkpebZVe9JzLhy03kEnBB7eDX+dMbtStbOUUZ+uUsEjLS0F3otAV+qe2Vn
Ib1aq9CFtctUK6ceb5uETae+8w0fiiQqSYk7kHd6R0DntTJLcFG49yV1vWhQv54/
IUadzGvn9AbeM59ylOiiCa+0abgd5Xdawv5PsGgZ90f9cY5NFok8aOtfPb5dzDsk
owR98MUkCYLRNjLaN25RrbRLrBWIbtGFdq8Y4tVT6R9QSTApuuHMdpXdsqUQx8+a
qYuTC1ZFYSXbcCCtor09RiDD4HHlTUICU9z+XYceGwfwT8VGXea6TI6LLWyxDw8H
5A7AyinIOR3khiXd+QA2JV6Wp7Q7gZwxHyfBA2ABcqajz+zT2Gb9CK3jsu9Rl21+
SB15nur1vUpM6UGViXJwDLSlW2rCSd1ATiCuJfF8sbsgLS3vEMbzSw9+wWF8ROp+
1GJiOBvEVW5InZ9RnpLoeSlx4FunfD8szv9wONa/43UIVpfT1QZT3OymdS7Bmbca
9k3pu08qa8no1W9t4Cw9/5w4Zd7E68kgvJ+lwkE6mAvWTFUmQMxNi+2Yexhadjuj
zcsqb6njNt5DdXKNrM0mHXG1TMUpbsND1i0rOSZvkIgKrvKum81uPntAxpQf9Ubv
OBrErkwk+s/1gvyEdykHV5pYy/H5zMPTE+6376SNuZdJuB0HRfONX4XAia/r+aXI
pKUDlfndYX7YCk7v+crM75pX+wSOjnQhikYpBqQUM86J3BuIKURG/Z4jbYiPJeJi
U1rox4KJFN2S5h+cwIesL7J7CmgDigr4hj5FL7FlDk4xUmXsCLhS58RU5/BXl6yx
bz6hE+oipm3c+S5JNh5oxm3BmqyZ5UUvp5kSDvkEXFXJSBSN+qrg7HbeGJSt1z/s
fyofuLxMYBJpZbEthduNr2h9dc/YIy/WF5a1AYc5FBODFu6cwosTFyyb7Rfvkh9J
qcT2Fg+Jh6/cVWRvVLshlzcJhZXBdy396qT363wzOm31Fk+e8IsexJPlf90mKLuR
DvumxAGN4ujv14uLpiYgMxxX8rojyH8GyqPc6GMTonWOJB0VYGMfQV8lZb2UuVm0
jcSdN9MAlvsn7nIzyGkkxUEmWnWmJoRiBMBfM4aUzvi+GM74/e5D+aVlOZMelJGw
mrLAtXjbicEOH/2L6fqkvvbm/9r9F+1KbLHV4pcRyf5a5ejJLZcZ3IupC26KnS6x
Ubl8+HpThjF7BaKgTuZpnpD/kRcBZ5yIIaUxDGivfI8sMUmJ8pBIrsE4kBOe2WTY
Haco3AtA3aI4PCOcAPzZnRKM1KA8wYgRSCITIujyT3kABQuGkIa2q2rzVxb9BQk4
LH1tx+mDKPf8QU0yxVoXofL9RLHrM0rQoZ/VYi6nSWxfopA6jt+ebzVm1llrvD+y
y7Lnt4i2QpZW+vq0vxCiLKtBHMiwxNWgbRfuAyTZSZ7FQigLmlawFeUItEgFr2Fw
ew15OJVDBLlOTmpyWz4mnSdn5j9wjRgxVON8LfVGBfcqGogX7wKJDFhRYIrmF3Jt
arbTc3JHNf8ApdjSpt3pS+yyKPvDzxf2vwasBXOckfEGbuSIldoDTevJnZZsO69V
nXAX7OlKccW4VuXK7V6ZfkrKOEP07T/AXPaocE/LaNA+MjqFgaQMjzt6+HL6u5GR
k34ZHX89h4Gj3u9b0sgXeyl0ABE0v6IBCXbbPtuSY6ZhDgV2UlVFaMBIwjBz6U1t
mKsLSwItPYiTmy4AvTpFAc64YlSlWhDwaRGM9w0l0guN9ubtqYRHcirMo2AMfr1r
OMtcuy4Ep+2WOccIPlOLBl849JtC9MZODsnTJlCZ7iZVPd+MflfnuU5Z63z70A8I
SOl0DIpHvw4ufO76hRAz3j1bzkh44j3fC+JUduFWkHz+ODcuc5X7hdz+CFblSJDy
1fZ3R2w+QyUI/zRTMP0nO/E0sVS1ke4L9XdQ1za40LD2FF9dAfRmoDoYtUU+4KeC
ziFaUi8BxHtFOxPIqVzRH9KUNE+RYlDSbPtK9LaMsgsp2nL/od3MskTguRxNQ/Tu
l8D7k4Zb3qxgRAK+y67qI2TmpiovEprFBhWIlCn/prxXde4tx2IJKFNUnq3zftH4
HHudQX9CMUu3/ngWk2V6D237RiWfAxtnPC4pS0TvXb0XPgzNM+C9c/uRURV/WHap
ypHv/B/kH7Au8RwId6kNadqogOlv/ixThIKbFVMG95KtD3jU1bjKRbwjkseU/JnT
imnxeVb3l1N6ADbG/8EB3of4Fcje9pLjI35Ar5a3MzStHX7A+Rgi9TAN1jQiDbtK
e4rkCbeyp7sjNRWjuftKWhEFtCJEJSlCUGRb7jTRQX3hzzLsBwbKPGy04Xm22IGQ
QqjYcWaesC1SEKoVkyz8YXxsQ1SZjmiSiUcaWTR2xpgrL7kSox8Ya2tjyouTT4g2
joUclfd2I1tUl9KiKLfmtAMM8QtgoHt4Eb6D+Z1PsZO5CA5LqVPtGI1pKnbw20tz
VbFWQN1mERY3jQgdWTq5Chd3VNLEn+A9XPtGm2M3Oo71OKB/Y6eb77rUauMDiA66
w3Y1grGy4tLPwfq9POJ8r3mkFcSvEtGzzc+8I5/R9jnqWh3MuE/p2yot50vLi4PW
rseJZ7Ce+CG09F/aEoZCZBMMLtTg2MlufX2IlA2SY8RocvmhjQSfa+GjLUFtC8Cz
Ul0FVbR1SDalPyzhDxo4hiAwSJUVMtYFxUKEWbq16v+woyCuw1/CI7hdPDUST23s
ZDbYoDS1FafheKTiaPOfP4N99mB1Hr8ZhkHdbgl/QAXy6VpiJX7c3C0INSO9U2L2
n1Sw5++NcZyHtLSmwBuatQkyGZl9bGpY0YGWUwu+XCC/xAGRfzSGjxB4m2pbqdN5
ODrHI8bGSbvQ9sdmFF76/UkK6mBDxL8cNMpTuUbtGFUNewRiETKkNZtP4cg99R+H
jOP5nerQKn+HuHEjrmHDJUg3JHCN8hDCVtjCV8sTVy8ag12nSHXgY+mcLQ0HrOyd
upvagdKC1FE2OariKBX4bzQpcAohgRDsZ1/6OXXPtHMayc+7erMP6vyL0Yn6rZe6
/f1mpzyMM2VI6eAJjtrHn9tZVI9BaQXs9Xx/yQVAFLkXheRPvkguAqpwcxX0BojI
S+ej0oqsCLL8aXlbIE7kxQ64xu0P5VgNOHF3jKMkJhW1xDJQpA9fXw6rSaguWKq5
FJnMlc5CI2suoo6jbrrYbTQToK+f6UExwb9/F2jeWz527upnrcgMYlm3w+U9xfMe
fDnsGt6IG1PZTy9P1Uk+8L/vK/DxBDRKCLhdjunwu6kMSuprASP44piefHRikz0/
SDaHmx4c3oGWJu6jSXk1gVpLZJwWHcN+uFYtsqUZNmdAKgCw243fSSCMNS6l6a1s
gd9Ua2/haUTKKP2NTUWY8J+CyznbjfAvaIx7I3ERbTgWKadCKm+yqagPg9W59nTP
J7MvMjQBi4VmJg5HS1vt/PJwhQCDzOkFpLCMvdgqb3bqCTpUR0Raoj7s1v9bJiGm
Gn4fUUK5Tjg8FNHP1OYYuWZP/tvQsAGsZhUivOHQQpgkvu6tnp7TJc1aWr3d38tb
7JnNG5oFMLuVxaWswVXeX5ZEKC+3Dt//fBVjJ39FF/EJdXGj3EzqRu9DKKKBeirU
IFKCKYBupHyMC2aR53YXLQKz5v7oQdbaHmatbDrstn77DJg8EEf9jn4KvCASOI3g
x34BnkfT0X3B/XuP8KFPD6oHNsqSV32FQiySx8WIBtqiN7euQuo3Xb2bNZzwRVVr
sqA06E2GAtLUreomBQNud/KBCfrLKsy38XXXGm7UCJOdNytfa/Uk+60GLZI8h6KN
+bLquSbU0Uqkq6e6XqSimmRjI7Ncvet/Igyyscv8wFpiEW0yZz+7YJ4/JJUzTllO
l9BCZEfbOUMuHVOmgjFx+aTYSoFah3/NFczZ0WQf8Vivc8w5G4OsHE4x5qVn/5u1
V0KRUn4/IUL3eBQLhNJrSgQXoFQzaCrqcn/vsWgOkFTQ6lfWinIVnMoA8iNbJXt8
QmYze2hZe+RH1xJZ5SQSV9i5lDPjFr3YUxuLtLZrQBBJV/JU+5JWW6cbt5l8Tx65
MMRwoQxbtNjf3wM/+WmHeRL4yOvCd8wdw5zfGbP00J0xSNfOsrJiVzQZFPSFutHH
jW1QnEWjgf0j0+pqCML1N73Z45b8u9H1iVlB0rKQ5cLvL6/6bdq+dxfl8IfYulVm
aOJD4jzi9K8Gtz+B64nkjGbBCzS+6j/a247G/lJfC+FQ5G05IMCyJG6AFqbAY7/6
j77s3jay1zdLlXlO+j8HU7KhLu7aOClZtegawAPL3BIAs9V/Fhl5G9dSoQ4kCfoa
GbqgwqZI1s1kj6PZ8gdQq0ldZTSX5CxfMWHyN6KPXr/JRQDTJ3xix+SWtPi5PTG3
uwJjROUcNwNzp/asHH4LplL8laOksIcVb5KNgVwRY3W1pQrTKZKNw7vsiE94RD8k
nCHAdOsOPNQMbs8qv/uPUlkcFHDSktTr/a1kXfbXdP+N1besqvmXzemnphTeFU/R
uVAhyoYodJ2lZW3/CJ6yjcGwTit5BVA0sKEYTPBiVPK2EjA119Q/z+bwF0Adodeg
EHx9gse7dxUsKv0a3YTiZSFVTVLNc4647iMTOYvnrSN2GLu661pIV/hqHNI+VCqj
XmnRcZOKU09YDJ45lQFLfimlmuiT8dCpeO1hz/THhoQzDhJ8D8Fr98+cMkmGiLPu
QfOcU/m81hUpHZK1Xi79ZCjenqzfdjiY7ptQkarx6k9EmRdNO+NU48DssRxMzJCS
YUTWKWTPJHM5w1DOPr0fMHtmdoOQH/OrkbJa5y26hYGRrOhW4oUQlIeqhfPxAugx
0DZILH8egDY8sFu5jA/bjdgjLiM8WKgZvoUw7uV9OJDsnf2uUhXW3bfIa2jzqfjT
qr14T+n/vvntw/QEIXDUzbHv43+SHtHoYewP0XKKKw1n4o05H1VcqK7MP/vv+5w1
MM6MBmyFngiB4uiPM6nzJFYE/4HmSP1PYkPHX1KpnsNVp9IBX9ALmp3MKjDJyf4g
up7wnXIl0dH/RshVKB97Hb00N8Qoni/ftOSDw+ARJBVKMvRV9UDr3jX/B9+a2OCE
yD2ZnC21MmWUXA5OwhUfKh2qSWxMi5+qVMrmBQl3TXQR1oj7wI2kl218MFZQvoWG
YxKVrMQBFXDbar3cdfLM+5SqGzIudszhecF+Sf1B1yDT9kPqgSAEli42wDzTrerp
pseH7loo0LIZiyyJDtPVAH66BraTlOKj6RRXA1MzfIUkDZziLE4CPI3qVGIk7zRI
g3lbWChHgmjVZEfI8wunEG/QDsdLwNTyoJqFzlYkiRV53v+MPAwLJj41CRvgHJSX
ijo332LkTXLorxkn7dsFqQ0NsfywczhaQUD+y8DyWo8JZIE4wHYpjglbCr6XOPgd
AfnR5Y2I938EiT7SrWRiCEa4HHmNEUGX4qlgtclOiG24YqgRrB1dk1B8yytaZ/MU
Lye2ha4IamqPyR8faLy2VvReLBrYdYMqtEiCES2xCb2+BgFiINaRIgBA4ajcIM0d
gzGhp2GzaNAFehmc24i6ZmtsIP2IfuBebQQhSXRM5VhAe5wCE2ZA26k1ayujqNOt
c/C8EdIW1P4Gyi2TZ6PY3HfXbK/C+BSRRAPpJppA7ldAtBijWjNIISssY64C/3Ko
3SuizWbPAuNTd/H/B11+YAb1SCcKfJJsU6pQOEqm3ACFZTJvGQHJflT0oiFSSEr5
Vc4tRXDMVs+ym3Tk2+hDKebNFA6ULDWKNhOI9L5z4JnuUExcsYffHGH9nhUopQrL
i5y2Fu1Ga9Tpzxl9RvsUQVkb4CndGoFBnazk6YGcKSZ8RyYEXkAc9GLAQJtDnVx5
wwzBJK1yD9M/NO0re/jx7Q9nhzASkIPiUtvurwuDP5ldN7aMcn7BZUUnXJtjugDY
sZCL7F18+37M6ch2kGXbNu5YoFob8NerzSksi6aNbSQCARMleqtnBcwo1DzKmpVv
Z8y4d3IltFOiS/BncWqe0Oy/Mxs5qWqMb+DOjbVTqFAJza3Wty54XIYeU/m9EUty
ukxId5s2UaWx5R7ydsymBJRhR7ZMAb9nCQUgKSrphx4FbSqhFIm9vbEZqg6Sv/C9
lHZwVoCsRVLLOH6WH5eZ03kXeLl65NQM0ylM6eLo/oeAPlgo+vI4mKaP0HdxCsfU
/NH+nchAlapRpS2yTRJ9H+six2fR3Nz42U+QeTP+NILMGGSk7qpoOVl25ce/jccc
ks5rPcIsREosLlA1lZYq/h1zargVSqGtgT79rKtP+eP41icpH/24LSt8EWb61Me8
jny4xudn/TPsmb+ZHYDaq9Msq5J8eAUh4bmntJ0a278VSZ6Rako/CuBdd+e8wWVx
OEKbl8p3Uduyb0ZLLdPbagVeLVi/ukTaBMNR7cRr+2UGxbDzVtyC73ThPYM4uxdj
+04Qwjai9WSQehW3jTeH/1AmvM8mhhyBl2IoCtEH1eH04kzgaSkukEjoYFZ3eaBq
DRi1CIEhhE1lEdcsJjBuTfIY/d6CixVfojN30VR6efr8tcnphQO1LHeNalyZ3fs5
3n7bhK7NerGwKt1VjaZmhU/lzCaHQGjTsGAJLu7QgOAyM86P10R8qdNOVgqg23eq
2gz5f6Li9zISuBj8geUTVKon6GxHXMgZJ22SKewNwSI+CoSHlqI6YLxdRxmagyjq
pcDXHS0laZv80pSJUIDK9XCBelUrXy3ug/3rAQWABSELAP96ol0pkrgcRwlyPBsY
L5oBBVI++S0v4loMNSrqejPr37Eg2q+Iwl10gb89d26Pi8xRJ5s7S6fZQbS/xRkj
QdgHlmLgiZF0FgWBK9lf/EYE+gVlaim+Q8Aqrga/WHJEAzYNGlVy1lrcOOiJJprA
VdxT1G0P+oj0N6m6c8lDTWO2NEVZB+p7bcLCsqaXky7r3B62YxeNER7Gb2Utr+Eq
h6XJ2U48rgdk4vOWQuT7JLEqKkS7cio2hh9bCbMh9I9hPzWREnxFSbq9EvLy2klw
lMbW4MheZ86mucm0G2chVcApgyb8l10BjJmZ2B/yRpkHTA9HdSt5557SOL+eFjQ+
xcEqty2130kRVxQhnpr/Sp756eUjYoZTqKfyExELIFGpkltz8/O9U4GfdmlprIQn
GV+hOkFX+6FKC3wLnlkE7yNsN+Evb+FPRfHBvszwmKohbYFzK27WVcwLfCpLrnSy
ELoolcycBKBa/rlx4TueWOnwg9gvJmfeLnjmZ76jg+webBZPvFHQQeajh8IcCqcv
J9OuMkf3oRf9YxTC8FV6sOplrCVbPmV10/e0i4O30MFSpyRdoAwm9s1yYI+bzQgp
yAyQSfLRjVNprVqFFtWgKnesJ57s5z2FyVHEmy3RoikKaoA0TPw9Q8kY7k3jLMC7
XQt/kNtTfZZgyM+oqreVu3d/CO5AJWl847LHlQckrLBCJbqj+0lzx5ONulE6IrVL
olUHgcgtDEDE8mQLfqgUqu7EK/brkqJTd+PL9LYQoce0UZG9CB6ex2ahwS1V+Spp
7pmvCfIk73qiHcZ0jHMLkPQR2PtQ7fXx5p98U3MmDJu+/W6vzTxpSey49LChx83l
1GS7vzfjMcLB+IPoUKTld9BQugKkUQblGtRvclg+luJYaLAA48ScU2YDsq2LAQ8c
lC4AGcP9AEu3mr+8hg7abukodqaKU0mxKXVy4zHMUJM6p4gx4fieHBiV31hule3a
1MlvHPNfZIDvARFq2H8dl/UqC+QxiUFvhcV557FSt/KIYW/+a0FGfnlQQ2Qfk+G5
SEuvuZWdeqyOK3+gVsoUTXUATd8pw54SjxfqoMFps7O0OqHh++3QsDKPl9FKkUwS
b+zQ0hNUjvfXPl7aXXig/fH0zbjJXWMMe77B/AnDuxxN298mqOJg4jco82d5+2/4
lGRhYOHqItb4G6hwIxN/Udqn5ICvLFf5aPKY2ek4T93lP0GMPWnPXY13U6UkDjvO
wUK9XQcPljlRvuDQIc2pJ2oxxV0COD8EF6j/OCHzzEPM0sMq8diqdxRY6BFsv/DE
Qble32gcFPEeXVM1IGr0euKEDRglGmudEkKgbjQIUsXivpUmolPC8iWTPeVoUemw
dzVMp7Q4h6R7mGHlwAkR4e6lJQauYsmmHtO+Zu9pdOpvOlsnkTC6PmUlSto/RjCc
fVFZ/ln/FFkvuvvkH6YzMk/K7F/zHPlud3PGEyYYcHxnFV2J6nfUXEe7zxR5mubA
08OtdubYMVyI8zJaPgu9k9kyf60Wq6nUF+CzTHhNqlwFRKKN6YO5gUHyn7gdc/Lu
iUxk2Jaj2lbCKRe7ahsrtl7HmG/AnZLsvooKTRjKQ6VJd7RCxWwdFHga1WzFKfHp
Efij5X6HLkk7HDa3RFnT79Z7OPP4Uan9r4objhY+nniUgztODTluA8BFL7Hc8Ihg
rRs3iGCoazV6ruls3+4uxTxHqwY/df5wBkaMKg4NVDykT+RFFK0M7oZ+C0OX7kQy
Ug6lC6pLZLG8yoSPCiSySjcYw06XXY5BdkHVLuxjhDIZrd3bgcf/r//ar8i6n58i
Sd3MTIC6PNYu6oK3f0tr7o5bBHPfnLdHAYG15LsMQ9v8BDZ5S2JblPppQTtka8+C
5nE393JWgXoDOtczEBtytZslvvvwcx0CwQsPl0veCCx+d00OHkQdUhq4jKqwPs7t
v2PuZ9VGgOkLJ1Ys5qXY/ej7ibeFhEc4KJIhsBPV3hqU6oNIfK8WJqg9Q1KdAOlL
IfgFor10i91R6edV086Xq+EanDhtL9ULaGr7WDqynw30E08rXaDG+plo+lRgFwNi
xpQ0S3UXPgo11daFpCDl2/lmbmM2qRvUtJ2fmnH69+9Xeu2W7jxRi4h4VilaWKXz
Tr6DHBCl+0N5DXA+r4GaF139ooeYhzb+oQEOV3QNP91FU6iVZ7579z4wai09kx5Y
IUx+hDjQmaGQZfYmm9rd6js69AjJOSEO0fNL/HyRQMbYsLbxZNGMMtyFvcUFFOwO
TlNvWlFbJcrX/Ah1JBz00aNvR2dPlui60DyrYccMfe41ZeZOTVzuFd6gKXDkpoFv
v5ZoRf420/f2GUQzaFc3P6t9/ybMsrA8elETA3l/s05G5F9JiXEaDzmN6/ncIKZE
Ye1rm/52upx+A7+Kiv/JmfZC7Ul2S1WGsX8u4AlOERi8uLGXfKHLAp5Ve8jHiyEq
MjTyCwXnhpciNlRDB0ltM2KL7aY2aHIszS+ZhyZjy+6jzYEiWJ1MAwNiYopSLOHu
2xTUfnCB9JIgNPmgo2xw6QgAfFZvWdprcZsehhWiJXjY9zAwXaeLVragmAmli3sn
yMeGnNXK5gfsmegWYt5FUg0ypr+D4Bd8UyQAQJN92lCpAJ8jbepvYO+LFTQjU0GQ
/TAq0NYLYZzqVNiKoWmGqRI6dgyZCcZaGz9vSW65Yw1CY3FcK1YVtZFCy5bg8QNa
VkgilIk4D4gWbbcHzgFkfvfuZujWXSchAvzDkJWOUXsjIeBqbfaK7h4nPrKRcium
hMrwXObyZ4/NuGXc5ddikEUFcZnMFbYtJT0BNZDrHX0w1v/Z7BYM0XRRD5RCnp7I
qb6B+iq9H5ZvDZB9DwkfYSWcHdAGIgduQODfYYSFfNDC57t4jQ9hx5A9roO22bkc
QsKgrhHrRlyFcdOmbgQd2EUBAFGQP5k0fk/WuDmOK+DJUjJShQQTcchyDnVfC+vB
XkEwBUmWK9SrOBczDnK+ddcNkE99G95YP9dIneIc2tf1iIkLDfNMUDGwDrMQQ0M2
Qq+tltsQhFDjA0Fmu6hg3NOmJxiSJhcht+beJ502laXhsRDLmBWB4GKYBCwUe9ts
q9h4Y0fhhKjxOsGjVDuS++CCmK2MsO1BmZHUFmUC8seNPq2Jkmn4ttFXdnqer/6M
8AhNc7FVnjvTi8QcccrtpnK+6rUBPJzsL78unupyynf4YVGxcd/bLTFotd8CzGvR
Z4eq+eEqU89MrzGUYoNpzb5rYiIpQ+GF11nURXAs0OjWSL2BbIXjZdQZa+WEbe/z
W08m8jv3DdY1GJMc0Gw9XO+KOyZnyIY0wBEICtVpwSZcmpW2vXk9v8Kei/Lnnfxz
+NprlfJ2fIdm6hDhnaBaWF8hUtMdBLZ2XyzS+Eyxg57nKtwgDlBWhPixdtBQFLwl
GbodM4qvsA8dU2nz6a932S5MRaq1Um6oyUEYYbcHYuz5Ea+hPgVQW1fnvvTY/WpN
rj4uSdUc45foFmKoUutDLE3IruympqfAZdua6fa6jnN3iNUQT6k+lUw1trZoLQDV
sSIHKbEOm7ZxY5AOlL2dG/PW1hCXRURFbZhLDKKVCzdtZTB1L2mof+k6BZLHnmLK
zXjA3l2BWuLAHDu/7UOiu+joIBCRyrI/ZZxlro2lMCHWfnZPTvjnqpIz94SV7LQw
CSDuxbnKHlPRhCSUypa3ofaMDnwRAlria3hloB1GyojavE1prsb7ShFqYWoJUhss
s9RBT0bEh4DwRsC9M18Qpfj2Q0WgcT1B5HvwZ3sfb7mjfBM0KAG3eu8GFRji1KIC
wn1CH84tA7O9zduuOWregKoNTrDeR6SAPDIfuKT6wxGLEe8Srg5Yyg0FqPp0vvud
sr/6k4URScyGBK9MGCrPNcLcyWwBaJ40WF1p12BC3LB6Z0OlPgKg+k3swQdozxjx
RGylDn2hW+hYhDSII+TFJQsL1LFFh+8xPiPkRAEaQrzaQdXRhGImXSG7JlTJRBgp
M57bnC/UBrrE/7DvasGVKhe6s7HJzYJOmCAegXKJkoNHKPCxazQUWsN2h91LoYJX
KsHZe2h6bmYd32Btw4CX6jPEmAdAQ3t6WGOOwvAy+Z0AOOIeSBgVtAG6i4toRaVP
ZJBdGbV9leWqcHTFG+jDuzKyLx5sKvNdbWiYlkLBX8Vsqt/JwuzOuVNGzC9fafJw
I3fpnyK87t6kBA3K0nckxlR1ycAGoNctA+6uc9xjwLlCLLsN2fvHzRpfhj1raBBF
w8+PCljovUnzPDs7JyeQzKZgF/tHOf2ytL9o0FMYtd3W/uZ3NcVJ60mHrEJl0YPI
VFk2yj3K81ofzNL5KvLZHEOu0buGzsRbxzzgvW6SfUp4YCFcANFNAsST1hzG0UR9
Xu/AcUI5CmHQIIVEPB4JipxbpQslvFi94KI8h3hw/zwgp+BBCHQT7BfMgENKn4c9
K1u0kG0uS/w2rlwADjQje2fwJta5Vpi/YY3vt7FulIq6EcsyDEaey3uKI0IDgllm
8COnsPGuKnUfkNnan15EO2YT8d9s0nVMLb8TtbZpqrjUzWhQhCceecQRxAzlk94c
prdo13dvgVdAKqAzXrnMgjzZE9kJ9EPigYLgcwTPwa16d1vNRaDqbbgSw04dbESH
taT2Om+akInb6THfBItdyOB8FJ/GxeUrr3rD8lBrZmOSfMhBciCjeEupdmBIcUUj
eXqwAS93wUKkx5WhKEkFr2NcCEBr2JxVJseLOsiMnoeLrv5pgFeJaPJ4XF6FxpgS
IONieVihZzfeGgg5eIArxuU23PZ6dg3d5vIWhtUImfAkf56K7Ts0TxvYB4rUYa39
gjDZmIpPqAp+F386z8DfIypTvUVz84MhNhwkJOoB4ZkOhBTxEzd8iAO2FRi2xhi2
iHmieQsLXkGsVWzcYmfpW1+Mf+6tP1HJdJRj3AIn9u+fb97hnxcohyFrWgISI6/O
shu2wLfBpLzDGgtQoz3Kvu2C9dliZavcOAiq5mZV9v2jDK+dtq0h3UQnrQli7VxR
awA5vdjstBIJ0boapeomRQ3Hn7L8Obk+XkG6IgqUZPfbG6YK7zB0WJv3E9ZmKJpA
xY+TONs0EhBtFDmgSXUqoA2KbmKuEpHuIiaqc9ZEFQSwllsHha6odNdMxlzC5NZr
Q6BqX2p0c3Bo6+6J2vEZ0KmKA83yQdkARg2o4Ve5IctT0Rx0+0zQpVpQMZxCksUT
px2dUyQ9qorN1aLqhRlwbLE6fioO/IWHy/YqUIBS7brgv1EZCLHO10OK9dUwiE8y
LybxkRqo43638+3Zqwd9xMeXMMyX0PZMObQjyuuJCCGgWdsv1Mfo1liXyxnMMk/H
ey9w5vUdN24awz03nGgQF1OzpQpYlE7K1vn8FFOfA8sLE875nCiFRQL1OGKslwAL
Wfr+OyJz9Q7pgG1x9Fk//6plb35JCX/nmy6lI9ni9Y2KAY+Z4fWMQe51LkpazyvR
XMsxV7l4BfLbhLLc/Fiug1ebVQSQAv+L1agTlKaKlpQpiId3gzT051cN0t+UgVIP
Y1mXFGVC9MO0Z8+VEugWdGUQjDTO78Y3/zmD7sUZT04T6/Oa2ScBdGRMpTLlKtru
JmEm1X3dQioKAh5C3os61Ekrxd4jtm9QyXseJMUDsYTxFL60ZKzT5EHft5gMSZte
Q/nd9hQxgjWViuucnYHRbDpcOjIak3Sa3qUEJakyW1umEWvYIc2JUEB2uv8guc+w
HJv3EkWy9CQ2WY0GS/KUzcZLAambq1ncfoTe+RadhDzs6LNNtnO5A5fxbKfFxUH4
31YuehFvpCsujNJt77w43yk1XSJdQ8gZQJ4uCKofS71r+vqS7JjS3rGKyfjZE4PH
qemqWlPV3ugQMacsRYCLeMGnYZLnNr03r6BdsSMa+y4LMIr6Y5up6+HTZq31Dcvg
DeCDFS+WrDyyioEV7w1q7TNpVYvv/WACLIlqB2M+PSBME4NVFntgH3CgaMXrTLmx
gp/YEk/jx9ygcx/ePIuLk3umaoNZOU1JMKzBOQNiek2bxe0tSbHp+wbri17rBiav
F0jrFYHPo01uwFjM9KlQXPK0g4s+xDytFmY9BAxfEZWuBf6AB0gVBEnH3F/OXokN
GMVsEwmy85loLjfhMILk2FeGUO/AkKnst7xVOeqmPcpW4IclWW4Gkxc6Zt0l6jv+
mXZuJyHraEEHULbxSVkO/GJrbEWzpPZM+o6jLHu98IGdbtj2r1J5WXniWy0Z1bzf
obsHT7ji57AfhrcOghsP8J5u4Wkte9AFseSU7Z1cysPid0f064oHJB3AA9kZyPuo
aK40enBtpYDKAzy8hts5b0r8O7zHWl9G/2Zi5Y0OyMtUWpolzAm7Fw5nN+4BXDb7
mNShfdRxfn2ujWzm2j3qC8qsPsdybIEZ1uUTvWkrZWF0bExmA5An9lQvrdidmgwk
etRBDu9bh6YFGsHnMp4axzg8a7vFF+EvhgaiKyGc/xZGs1Xdd9t1+Qq8E8lToDz+
u3zHLkxz8dRcxyBqqWypj07AUj5kIXliklLgnEKbbWaAlwLzJvq2dhhIb6a3NfDh
gSo/jf2V8f9NVebrMlembaQktCJrIvSAVLrd9eb/bcMpkJs4tlRY4Cp5RjQ2zYyp
6OrgaYGfJnWaXXieeOjEH05neP7v9ad8VDPIIFmcRwXHmIPR48gK6c3g3vVWGkyV
u1vt11urQQWAWQhV9QUIe+tJe7e9sMSw9jJIIElpD/69MLRJTEcvnzkcKXkkGkye
Qw9x598oCXDuFfsNwfYvQQgQq/nXfSluiUKDFy/63t1hd8uNT42f0jSqbSa/e0Sg
HzUi/GIAInTN7l1HlIzYHazsprqojwfuvNjgoJkUL09RfyYWyD8Dz+IoQodXmCDD
jzYf2eeubARYUdXHpI3UCdE6MsKa8GxrIDcjFWJlMWZPnZpc9vmF82x6+Ox9NLHy
gCtigefCqRGzqSyYHR/RIZnUx3qjp5Z2OdaUMyPM361CFa7yhgBmtiE+HN/fd1Zu
VJD4AUAv88c6xkru1/FTefv17PgXQ+MWjcx2x7GVHTLZbYKX3k3vwWWEZ8nDNUpo
/kcfB1AQaN+/Q2GLZIE4xp40Fdf2utXN86l84VT8Hu2uNPFMasfemPsNAaVq03Cq
kPTkG/y1mUg2i5/6yIYvhQqCddYo+j2GHiVHXaE8NJsA1PVG7FSbJeR0q4Unr5VC
bVFq2osbUvpcFR0CKEs344FnXUa2+ZaVl3YKUvlPaL4fU4eoUrmCeLqu4znaDulR
7S+elPNhjRIU9UpwCKNE5HWS2kQBqjNvN/3K1ncpxnOHx3WjqPJTpo1ZmFKqESlp
7WA33Z5vAr7d2yX6GW5uAGktJZcwaM97bIvxFzhGNbO4Zc9MV0iLT4bzg/5Ghb17
O8r8/2Q3Jr3mD6g+scRNish55BMd5Glq4ikAn6GgdCNHzxOp1nfzYR/YfrFTi1yH
MQgC3+fWgP0hBBIp9HfmuAGxnzCTcFkcOrmqFkvUewBQHwU4suhCxkk3rO1vjq7o
eA2n0rXrseLsU1CGZLqcbJmXZaXTS0Vc209yg8yFhUDyaTbpQMkjVA6quqBXDRTz
KbJPHH2rujD/XJoYCUWlBtSum4slRTIqJa6xfoX5GXlwQ/uh5LBjVY5L/UQa0kgw
r7RqqofpYlhU9aPgxmV2Lnj00OZrU1qqMzBFalO/1+24M6dbPKn1P9FWSVUTRkPU
WTZtKQcthx60AFmDLLC86jGLp1dzIGHYGZvkF1yhUAMs0C40m5pd2clTuJ43Ljik
UfAnRnFVMvkcvUg1SgIUgzk/zabxifPMH4BisulSWbnxI5NqIdJzjT5mp3T+0vD7
qM7bccAXNdLNT87ejgDs6ofbArIwg8M6+UxX+Zjd5OI0W93y/tqh3HDHHu4k3sF/
8BqO6XWnX+jtBdhbVEdBBiMNNg6cYpmIT55sGnXH6Fo+a7n7wwNefJRwHZfIvUPr
8rXNAr4MvN9yKPwNPNRn7M7hwcJ259rsbijV+xBo7iGrz/psLL4wuhI6IYUy9pYk
5rU/FVio5Vxrv3hFuDgMYJg2Rceoug0oS2z0UZ/syMGuYnnQkXxBOaeUGbwIHALF
nUzUYdFaFjatNP0PdOHHt1cYuTAXtgRmQ71k8JLSl2jVADNxayk8A1T5572/LgLQ
Mty42OShXtqh1tJO+3jfqryDv8rk4o9eX4TVrY/WKjW6U5i/QKDfWV//MJJzQkbu
AL1IMBHVqE2/+PXyzXcFR6Wgy3bUDMVFkXGTqBXRfOrxQmltZLj0NT/hGe+UsDGV
JQwNFQX3loamcNtTIXqzi6N+99G9FEzP1VFDDDR9xC6dKsrn/XWksEdXpM2baeY6
esbH0WxaDgcagwtLofi/fi3DFcxOnthTIffgQdd/qy40iHsK5OtEQGQR+8And/PO
QmrRoWkkBWSBUre5KAtG6IKzK3kkRftGvR2669bL3AaN71RSBDQjLzhCuaDe5TXa
8I4pCq2g1L9NAbnz107einOZ4zKjTVaO47nFDFk0hPKIpv4zc3/ZmVGfR0fLeSJp
DmMmX4z1b42IDRKjA1mYrmtP77uNvzRqwKX3PN05YZ8sLM1vFvFVIVwiOYthviI/
Ivtd6XJevNcAhnSAGpR4/uLdUZWLI7s1T/0itZ0Vbe3kE8Ye7zeTDlaGAW0nr+Iy
Q6E2AeMrmgQ9kzMPCnE4hl4LIckpIZucyYJ7Mbzopfd3l6I07d4+4WV1TsoehzHr
f3Gh2d6btXKZHQXNShDgHh/uuMSPfA437KDypNpaKcXmDH0dNQeO6NB24kXtGxj6
di3AP/8UTzxKAXiXe1Rfn8UXkQIRR7MJXbBdfEHFgVZHjLzHJXxVfM8cVSH8Ejni
fXgZ5oosKWo+zNBrrF9/QCrP5pkYaT9rSf0PQ8xF2Ioeuk98SlcbdTFhLhiUgIkE
wNpnGepJGV9DKtMez85NzOmFORwylsxqfJWHhh4XF5F/ygjL6nlI04LZr6BSNcsg
U7WYWubFnqkkaXAmEX6ZlNOOFJ1CWzkisa2dFTzl+PMP1OH5xy/Z9q1ye+uiRBer
DlPGV81ATzozPghgKyis7+tm5M/FWK+ZtZRNM0Z+A5FAJei3DfKzQkGwA54g34bP
IufK0oNc/+94Tbzoh9hWGIhvpOIttSQ6ZFj7vRwarfEsaBWsHW2EfWscCtK4t0B7
1nvh7ZV80oaMgypS1p4nA4wO8LNXPWtLwl+qxiea9MNiSC3vNC6U+k1fpbTML2OE
G3VeXCzNnJXeUu+wOHfn/XmlJ2mXZq6w08XfZigfWnjvjnVSIJhWjnjuplr/F8Ze
r1teEOvCUTn3gZXUOY12oKR3AhPK23A8/vbt8ZF0xwpN6B3bL3+WPtaKRyTuD+5d
jNrbttlTtFV0n8/RvNSN9+nna8wR9uJtbhaSik/PCors3c3+z9bpsZtM5MPCP6wp
u1yeUQOruceu3Z+pU43X/hdlgMAUuKHar29Gaw1M8oDmRIYW7ULdogduh8Gu21Jj
GOmx7k7dxWQqadnx4fkbEeKiq+qOUtQfcfgqr6iyzCvTi6LlvpyDlgl5YN6jzqJm
Wrpi8W6iYNJmX4O6595N2VtP+S2YMIZxiWAau1cI0Hx7j0ZoSmVl9UqOceQWivD2
ZtYc9G0QGKgrpXyHOyWDlJi0V0FwQkenitvoHY5lKVSZPFTF3qoyjserdkQnUErf
z0hAc/ffpJX3GELqX0k7KqBl0A0u2GIa8FRj7pDSCe/PpecSeLiGckS3ujyNBbHZ
A1lPG1OFLezFk9l3ROoa24oW9k1lZhXB/n9ogAvcvIkdz4gcLTuGKdj8R7Z3IHg3
H4IZ4X1wcmfXLX3qCt4YbPTWfY1UR6EkVr65xase/FEfCHIjN8Fsj7AY2nRGsLP4
sZx1yRo1r5ezvv1KwiE8GKmh4X5IYv5cSapBcx1ROS9oxxoGjRhXJtc/kLzhoH39
eORDzthG4mkc8yPbFtwO1x9PJFLGXqxRmt4WbwcvMhxZdJyBed4SUUYTLGpUVH6G
pG5LIE05fA0zrwFGYB23ABQtq2MZ2Z3xRETHBMcyLe0j1RM8waCp9DHLgRFcl+bD
9FsY3gCZClw9qdqbavJ0p+2E91cs1p7lJ+tIm+OMaJ/ZnYrCBEUPQqH7VAuVfPdT
mW+EJ4xDCLPjNWzTe8QRDNzVtaF25ESbfi/Fn/EPc4h7hIuf3KoeRe87J3ogy7hh
SYJ1Hp1/67v2kLQCLl3j6epa24D27XYg+JQrl0MdaXbby6JlAotvV6L8O/iCdSST
uth/PnPHxUii/KgDqCzZhxdZ+NDsGv6/aJ3aHGZVV0WdLujH/K0uxWi+cn8pvzr9
4QZ8B650er3FHtSaOTSlwdWGb4+xNYwWE5ywjNyVfXIHvFlyr0o9nH0zclxA3y+h
RPaFg1OqdfSpLSGOLzsAU8xcd1WRO0/smR0QPSorBmjq4fvJ3Vot4gBBdzWILJv+
cEzTMEduyGHLYsrGRrsw50o1VxXKm89vDOogqdbbhmGYW35LRi+5gxZDsHWK0veq
6SS8IZMiRA4Skdp6U3JonL6tIj60+0eJW9HtmiO4twU8Shvz1rz77Jt31mEWdVy1
e7kDyTItn+M+keXHCpmI089AEWvYHyrg4pgOF/yWoPeOZznYj17y2rkWNHybkKsX
ExeRMQKsFj1XVx1Eb5H//Oil4R/R/9PNaGksO0Wjjb+wiL49sTf9lduDeoLNDFaq
WjpmVd8zQgKAZibZPJ8s8+LBbfcFWddWrZQTNMAF0cLfpns8J5gWeZEe69kM9O2W
KJY65sE5Ammz5wdSJM3g9nMFwmCV5woC1oI587qgGmJE9Tlop84qrqCsxEOoEBUU
f+oE4PCmozgTKTJUSX+BcAfIMomQipkbnJLTg2sWYAib8fqDwsfmqjqRUQ/A1RSv
oKmyL0N6yVtdhZjwagANZp/xECjbE8puz9xcuNStr9hzRZkPVymGA2Aexu53HAUu
D2xKCxXqkhW9oqG2QseZ6NoTFM6XBL3C47n1oTRNFWVa3nk0vX90J64o+XaflZu9
woQHc6tZ2bKaOauAeKGA53QQwtH6M64mSXsa23MLBQVyU3TI5+Q9fQjxXGbcrKUr
kuPRHSE4NjpPQEvqWAb6Pg2KzIFTOCfdy5L5OWVmi7t66KyNDlD4XpFgqcj30SFL
PZui1YdsHKZGosK3I8Xr8Do3GNyR4JsUa+AROU4RcEo90pJtZfrD7ycd8eQPV7DB
vNzrXBA2oEFgW1aecR2rNBDAvIxRhqQYXqE98Rj445d1ghGt31WQ/3wemHKHtuiF
UMNnSIWPMHGNeHDsTqSdgIlLxBrLNeNA5G7N7L1fav4RsSMBXtvL8CABrpAiZfqz
Xr3DDgzOJsoMGFEexUSdG+lBNQcmRAuPX2aPIf8lJz+SCKfeEGgTqPoRcfGCaZhp
8BgBFXMWuCoy8+mx4qhicwdrXx54Cv+V0drfl3W4GE1MCXT4k6nAQwcu/k9aVFqq
yns5S2NKrQHfijhZ+c4PdXO2myqZJEbRJ5CdH9ldlHbCg2ZJMegbNELiTJep2fxC
63kzYS/2uvEempOBGAFtKvD8hOev58tvBSZu96tnjPuXw0TzQeX7OuqvHMIvWYwe
9pgwXw83XJNGR2Gn55MhlkKi1+7oma20dCesxmx/ASqcylDco9fkaxRPgvmwc2gw
KMPLObFa1qnQOSm0L92uCf5mU5qICw/YPGD/z9NjlfqYxdsVE3FBVh7A0bUKjaxu
CLzJy1Sdxv+rd9PoYpRntLYGx7eQ7nwQcKpi3507Aq67x1bGefZQlW9hYwMZBKqo
b8Q5noXIkU4ubucg3yweIS/OrXiWfnvN9dsSG4Rde80OU5XZDSqhMbIseeV3O+PC
GLjFs+ObdjYHHVSygVBmDi6Pg8C2FKv2FYJAkuikZcuqFLKI306QK0BuRREb4pvv
bFHpkcQjrF8kxqjYErOzjZOZIWcAKvB1btRWhjJZ/v/eDJIifuJAAyg+L8Wi6y3M
5yTIjQa/IEiY0fMbCAjZxFuIygsYyNhnMTryrcIqvlwqNmoBNZR1RHYl7GxCZvS7
qCneNndypuGMaZq+EeBluWY2/IT6aey3H70rPoU31sH7jeRf4+rscly41QfFEHmP
+qC24RsoCOoKbG+uDdEu1BSSBWhD27O5MWkoZbTUgFmEPnGzNKqZVBIEDyE3X+Oq
J/hDWew3EbyoQ5LaZhBQALxAdDfbvrwZyL/YKaprzfjfHaISQ1a9OyDjTeNO9UDU
voUvNhgbLZ+G0PXNg/23MWogQmfpO4OWMIOWrcyzZGK3hV6zN+idwjTrk0bMmYSS
M+QnFveqeEAD/dKOIcT+hNojWHoXayGwNHGj9LuOFvoF9VvsGOIVrpuvyO9+bXzH
95vJu0J5DYor1L7VQ8+kBYCTgoDTQEy8kXY+Gx2CHrJOO3UCOWwqrJpTYtdiRAvo
gLpPhVMLzB8ii8vaMgKfKVhrLPK7I0OV3COEL4tu+GsfYux6zHHciGXcEw0nmIM6
VwMNCV0hSPs+pT8VKwWL5EsRdqtnifGJI01sR4r3vAYYQvWqATtSuV/51gO/N+3Y
ZfXThIjiQTf8/cDZkxmj+dqQ4wzZ/4vtUPTDkl50+fC7u8hgw/aZwh/gZqO6JWR1
EpL0mcDsGgRG9PTruFWp2Q5OU34SrzwbNVtHiSYrqunSTI7lh3RGMnf40xQHqB0f
c3C7rbUpwLC3g4jpTtkgaERlNAuytSnBMIRwcT+LyjTlw8eChVXic36ceSGCvt4H
+DOpDE022Yb8Zt1v24gzBp3wM7+n5KdTeAPDp2b7FJJyxMqYVbE+3ZvW/UhGIh9Z
hOVBIRAkjvI4/FFqXWhC4EoiC3KRx1GgRq0c9FnpIKkin6BRmPalHoHibGzYNaX5
5xTM+a95XtCh7hWJnWdT+h9KEu7cEbw9hypQdxanHPlqcuPsyVSX7ebvlohjvA3L
TlaU+WN7X8xZdGuNmxXJ49COv3okY26qj33fE7p7arizvIPbpWM7MqTi9S5ZVKoE
UiJ86sfawVzW4HJYSsGcBH8TucHCeWvGJl6+9dz3PM0BCA6AkXlUSPUC5PgQdHs4
Pzu6BDovcILkOZr04VX7Pqe3VkwOOA/bFp7VaQIdmXGL2cSzV6SS3fZ75Qw3i6aV
HdM9nq94itJ2SG0w2Cv8sQTjMKXiKDHuTvd3Hxh5yzc6O5lU6bXWd0J4icDBFzEF
C48igXHrMFM/QdN323HLzIAhTNDbHtXD8MnfZ0WV0+9AatO8KrBP9uHEtcov2YZ9
kifY3TEva7fpWFVsRlIJIfku7rLf5w3FZufGhVHuIqIAVq/vY5B4gzBmzhVChyAV
BtrqEnE0e2EPCcUHyJTCbvuqG5p22dpD8ZoTZQqRV8LS8zE9qteq45QB1qgL556l
C+cmssCiYPoHvoVBsmhsEI1hhY+ITZhBX6X3hlz+ajf/iYUPiCUdKH/9I3O/7GSP
Ifw5j/gj7cV5Jjf9Nuu4d7Ta5F5R0IKTN1oAQJBJpxbA2ALdKHZohOTLj7SnC+D2
tL/gRVfrdTgsYKFzXPwNjN2pXutnINsKygfXyBcCODD5dlrVNyluPQCK0ZEN98+D
QG6NV26hHgy0uBamdGkIGlI5AmYxvNVPPoqZ/E2JCOxzzdyYRn56whByWnW4u2HJ
ryeFw9PbDjk69jNTiPAuPjbGMd99u0OhJ85m8Mg3do7YkmJ16HKpTsQbxWx46qp7
ijleYAiAw9RAVqlNCzS6+Nfwn3PJwUaQ+XQ3qKhK+BkfQCZORKBgZ3NUuUJGk0uT
ytuTAQBX+ML1e+ez4TboW2VSYndeSgGhM5NOXlnxk05vowtmcO5wrVS0oLpXyC2K
U70Mttx/DT9mU7/ya0dY1b9HYtdoaGTdJICGh/PxlHJxvLjN2s4KnZNJTRjVqrt+
xc1teYknrP1mlG71FVIdQUDtB8nDwpLzahZZeZgSDATIDivdE+6GhNDLEYysIXeW
K30SJsIQdmk78X8ZXI3uCBXHo8pA1617Vp7bq3SnhFSTUbHMI8ik5WtU0jU+qDnM
bpIHlCXYKF/zfZtGSKf4m6zX6lNOCEGmT0I3tplPnwBlQERnVdbDWadrKIXsGs2F
cA0eE7pAXXOtUO2uT9hLhmNDOmBGo23gpD4R9j3Fpsl+QgdE5gRrWTPOjysJNQt4
tGFCw1pg97fBIA2ptLbufg/AxXKbqPH09OX0kcfyNyPT8I5A4SqMt8HwGW/4UDF1
6do0Ufe3PWQqfGtmHP3MivPPwwDVY8AQVJtfKDvgO6IDh3s+NhgYJHRgh7q0Kxgc
EPxaa+xYmMotACc3A+Dq3RvblGExJjLpdGZS3PmiyBSbSItyRGywhvg7kE5RVKnM
cyf5SCsQmFmNJevdRVeIhpIw7y/1Lc/yit8NnwdD4BYtxL7edfG0VY2IIKC3FSjS
vRWZlCPvES7saOAZyF9DUNXPRMiXLPY7Df0XKeloLPaYzaZ7sKXYIQ7S6SiVry40
XaHWX+eMAB364jm1QMsaozDpahI6Rmn+FQKb9Zicn6/dvqwyXkF0seWnXRZxE3wi
yVlHHoB3H8itYLIJRtuXts4kqu1RG5P5V4okqeAe5VZEAceaslDCf1fak0iR19Py
JLuNXb5rznuYNCMRWaCwwJI01ZxEuc/hLwYc4r5z6rLhc4aR4hty1V9mHw2dvv+X
aYaV5RaJPte4r41phPqCftVKeTogQZYHwzZ9xauhrDkuW7WJbnSQYgmdRmCTCi/y
70oFO2EngQmvNdh8IG7MN6ln8aCWv4zf8Uauc4Cb17OzyFygxscxeiPOdVrWIr+d
nS2W3AtX/ZnLbOyyoNZqC0PeEElEatH94LLYvog7OOdQ7jZQasBmZGQbIMgcdXEB
+6DHkUgq3rDlwVtwSvCHPg/i0Dw0ZGYdOwfvIYTRchfI8n9cb9Zh6FKsSkonvQ9H
eX2zAb9pOYPWu3RSYsT6Yt25mgcU7a5Toix9Nh9ZNbrgKPEiwM8aojaDeu+qatnG
DCWxc2zyXkL3gxP+bF2BECI7TBlh6sbdJKTdnkCHPsRfsidAHY1NUqrK0O0zG5TY
/eUF9savbVJbIH1WMVeSJysLV3T5elJZgOogKaJc8fYVr9x12mUBVbfc/e8uMi3+
GVgVTEbwOxAho7aFq2qYNEox83QwfkJTzMGl8HfQSsm2NysuiVydxwabAI4QY/gx
J4OWQFrtUqn2nv29K01vDUq0nx7Tv5DB58p5V924GRFaEnGG9/m/6L8MU5PU94IS
oD1L7QHTIH7zS8mJ1WupK4wxLNo2SEf+84KXySdqXLK3kDw0BTQjlge/WPK+CSLf
TCgpBXv7LC4+gafzwTpXMV2ruejiZKDlDo1mko+76sOdMAgiY1Jc/AlCaMhvlZ9i
YWkq9IpTledRIw208Kxk5u5KFEfAN1sOjiJ2Qg4Ah+3/9hxwxuepJI9eIrTXkSLa
eLh13bFWlHl+UjyoZwbjcGg2+5umkBMc98zQO62k7Z4l7bYIos2fnI26/0t0GQpR
3aEWvG5WNJXcqRu/2E+9gyZJHtnjahEaUzVG55Fw0vhE/A8SM/q9COzzsyzv09vC
z6nIgCPgphp4C3mznVdDM8NJsxpIogqbPfYr9aASU+zQaWNoOt2yeN7CT3VL4Uhr
RGIZSitTENhAtsD/HFhiUQ+m6PXtkfxC+cfT6R70aA+ZgjFnzV94AriFMnhAX+wa
rSP/tqeMN53JXIUqreLwQv48D4FnTdHc5vPFe5zV3968r1TzS+nbrhPyJnn6xpg0
saNzB1dH4GXslbNzoKpMalmNXGWB7XFdWI5LmuGrKDOa9J5Wfda5w2AXlJRw6xUZ
VUZEaiIxoT/IRnq4AhS2DwGR53/zSMCdh3Sk4sRCmB/FLCDTFQtfyhOQiLFezik+
1ri+6i3DXO7yYrFxonEp7CgSd3og3mvu6/SRAXe6vYu+elu4T9mEpNlMIEUn2X7h
gqpD/uMshGT6FIgfALHjdfQudKsS3240jDAWB+7qekzPtz3I8T6oRhSBtzxtV5Bb
8/J6dCga2+stW2C0l4T8xH/3Xff8ops1VGZTWjkKoOBj64rz1EfgarSfxsDGXDo4
INeUyBVqhGgRb2lFEDGTz9pvL7fivLN447gvEghhY6GqXQjy4ds4LpG13HPiFJQ8
vvbt+Px9PUkFryMyFkGQlw38CYEygZahAX5JrfXOZ5b74eiHICTdEJe/V2v/xTw+
beSxPIcClGybJhkn8ifs6aHRkMcU8KM1WiSo8fIFuqCwYLRQpS5OgD4caNQ49iCT
av7nTTnw02/9dBlBb8wf8ep4xmuOvD2ZKj11tP5n2Gu1MqcsRLZovFBhGYWJBd15
dDiBOQyFvYaobn31gnSUOrkCj+hlhHOsiPap0ZVvr2Nlsx8ZH8X/vI30/d/hOejj
D/P1BefkEJkJRY5bHFo76CAZxvNFcKeA56+W4Y2a9NhUNfaq5G/nRJG7UJCTC7NB
TZhjCIzb9GP1VQlt8U7J4I7atCNBpWxFNgp5P9TySnMLjDHLAH4sjPeeLREbETkU
/axdEdXt16UOvMpSRMX/r5bnmWTnhRd2FWau4UWIDOigkO1MqeK4k5GAvA/Fp/qU
Ni+EKjz+2dKal2/C8Y9Kah14e8VI6h03r1gLmzoOb856nFH2L/aWP6Aoxz0zH7X8
InagEZax5oCQVi/CW+qnPuZPu2mx9CHaLaRYQQ+gdFoepIlH5Y/MBHjZ88nJkULK
ePFVLClhOAHQowYufNIU594RAxV2QUw8O2VB6REKwQ+IVGawBT2qKeO7D+CxxoJg
k+Gl6qJJ29OjAEWlIbNMez/SD9mcmfWBfVIoqQ02zYPgEy5REsmvJzlrhiUZKQlE
+NZ6zHOnHLraHB9LbQB8ESKdtFDnXOyAqcKyRTkelr9PDXxv1MfcjkfwEqfrO9Kk
mabiiO95KhdQtjtcntFLiS86XtC+SMgKow02dNQHXcCIh/4VWHK9HjC68274x7+o
YVvs8oiX0TUuyz2c17cFSmhc7rkiiYvFNXD3e+r8t1pTDyxQ7kTLkxp1ZUeN6U1O
J++l+FfKWZjAglJ3xWW58qJH9I7dT0vDuXVSW/+R8FMek1hNRfkXW6fRRqFjb7IP
xQhsx2h9tR4sIdQHcnQIriJpPbLnWrlAG8SGVBWVQ/sx9txiFa8+gK4+br56TIts
A/2P90ToQhrfmsDigsI7QbQpvE3DEVNLwQKMyU7iarNCl0s3wL+aJXCM7/NGjioz
PSYnKQZirOv2V1PFVpQEjR0vyCbAYsTphgkj5ukxJ11AN4UjwfUyuN2Fj6RJ+rP8
FtHLJ3sgjaBEcNJj1cLdm6LMqXSllJ6gms5M5W7Cnd83Q/HMo/xCrg0aSB+laMsg
94QYTZkFrIuVAJ6EWrd4A4bYy95Ym0+MLl0GwiXdaDEw32U9UatXn42N6agWQ+OX
tGHSZWFgrmZSLBO9d7lqYpWhAHUa55MiVOI6vrvp1ZyaVudu59FdELQBin7F7hPJ
GyJ18kawSnLO5A6QP6W+Bkrboe6Whh+a1F5X0YkBdTkLgIsnsyjQl9dGnhj83j95
CoG+Ra83KnXQKDQEll6dAmwJWDGd9x5+X/aSvKtu6uOvPrUZ0wYVQ8oQbOhFaClj
GpYRdbDD34vB72YIYfFwwkdfla2s+1W2oy620aJk8zSfJz7gdbWMKNNFJfT4z6P5
zzCassSFd+zcwxasfDG6aS58BpbV41OmaWsbZztz2M7/2VN0M2ilLLQ7yoSSgdtj
r1YJI9vvVO1fm019X0QTDKZVexPYRUf69cDcTXCtZ59YeyD0FMnj9Zw4AJknzDCb
kKfRQ0VC8sWdK8hxV1VN6GXOgXjyEgtveRdihq5aRVM/HFT3G28tXM8Q9GcNwbek
Fc3eay80L4SHrnIl17YxSEGADuUrXWzUdIfHtGbAiIwYzXKskwS3+MXqLynmTA8Q
rTDah1faAfGhENBUl15qjmGXyX8pzWEVkIgKZmVnChueJUuWl2N0tkDtNUBEgito
NU5617L0vv4rs2nptKmnqxCxVulZpcKjzQeB4S37/M54WbJGtzCeTIJ8vE5vIJu0
QWqvzgRlq+kmln9F33xbHjkbN/tPTa2LE8D2UA9H6qST4XV4H8qXDgpbYl037xvJ
aMsXa/Er90dpmuw1AQC/O881bYrVc51pgIhwXlBvS/lGSpy/sKYdbrVuooULSYQ8
u3BbMiPenf5Mr55VgQoO0eJ5wjtcAornWqPzeC3Pqud5MAU7AXN8vbZmgVk8iRIA
lTgNmk5zjKHMVD+Ttqk7C4SY38Af7LnuzsIy2evH1sJwNewQQs92g51A4INgTvDY
qC0kR8DWgj1pmGODng5cg8tjE5rnVFq9SW2swLgGgl9LJeaRPZB/6BRQZGkt52jN
vMUmcuvM9XVci7rCjXXPlitJaBuOyPf8yDWICvjdixlo3frjvmGWoHEKeRd0iKA2
LNPTLtykg9ElnEEA72qn44k60Kv1ciCEX6rrtzjZ4AY/TLN7slycR189BZ2sDcsv
i4yTqFfx7PlEevTmigXGzr8cLSKArk49QWiggfY+ePUm/gqcjx8Qydbif78evh6R
plhImLZZ3NF7Dtnql6dbYIROhKnqMA8FIglcik3RcchVqu7DI5RGN54H+3Tm709T
jTKObErIGOaOh+VsKOGyMD0iZaifnAn5WCNegD0BP7wTf/efHX/AS7407UC+YXal
B/1zED90HtEsLyhgsV2xv9kI6HhIagE7fc/3LwZxGrBv9P6BhoIeY4wrawcd7Av8
z7fMPRdbtJ03+k3g8HSVKdt7An8FWDJSPdZFcrcR7plbEpaXEcO/vsh4dqfbOsnZ
sa91GcezxGYWxM81RlvCAg2aGZQC+iwFmnT/qEbN20f+61+M9Xt6+21I10qpfNQ+
dKMn4cLvOxXBPQWInt5b//SQYCK0jS1+/ewP6fSZT/oXu8coCTUpgYB7WEi1HsQa
II0WwquUQCHu4j9FP0LhRJTVCu4Oh6VLFSFQCFveQR9iKI+OkvZHCNXZeyvbkV0s
6cyaVXU6zD52GBRWqsvxtRqd1zF6JbxFubOxMwRqTXg3pXbBhUg8sK3EpUZ8AX3T
UdgdR1q4FdHy42OYERucUltfK0tHPhjyicMw08+xeAs2PpEgMtgpNQJBYokgQNnd
vLhj3RxnmmPXGDlSfk+Ikaq7RTBw0iE+wBPVVXWVatO9Uj1IoUww9g7VVHxSxL2w
zlXBJhE/KD6R1jdwF3JO7t7IRBhSWWPqoDAQmjprqTqAvTb3LnL1w3Prrutbjhyo
JyPOCZ86WIFVI/lsVRuzvEyHyrMF+J8uolLoa4ftdLehYAfH0kndO3QFTgSnnV9g
Mqyuxnp4r2NtDIkCwUEafByNC9tQM9VPUUjJZefO7vA0nnnBN+CHs8z/MNJKfsL0
FH3EB7RMlHUriu2A3iS3bL8uAeQpjW0dCAKJIWm8qQ1C819HvY5nmvTUuEgivP5l
/gqhOjzKD3ecgyXBvRFHwbcgxeWbmZNKvaqWk2F8Oxlf6yJ8hJOQzqiPq9tlHyU3
EnDoGNEyYYfGOJK9ezR/iEG+lVGn4GijSXtmJz8rPwdEdE1wJAFt1BQHgX+PBUkU
bkF1Z2p5YCNwaiDrC1YL7OhzEKdDaO/clSqkJehF8k+AD3UA33BDz1JH9JFxSCkS
mqfm2ppJ6BLY3yBjBp07CzFLJLfey1w/+YfQfCmcF/p4FD3MI3NDktsDhzO9G3QI
+ejvTtL74FIxcwjHK2ltd0AUOi1dqPeLU099CHZ/Sv3qrhIvnZ5hueg3k0xuunrf
ivWsd77ucXF/DfOFUy8R9nxp6XKJLnGfGa2ti7aHH6boEAQAVsPqQ7y+OUG6I31L
nzeOZ01mrv3tUul7SU5BdnyvQwLE4RQTaxPk8FWPYWPHozOr1SlrCc7HLyimk5Ii
6mzYqXMeVai4aAW6tdNnIWk7Jz8gXqlouOaX/U311Lfmo1ZN6v60yZceJ/PsC+91
93KxHRhrAcxMYaCp5n9YZSmGRNBXNRIDcSGyKrp2NfH2183gujKdJzyMNbmHEHPI
/8E8qWaWaRd3t01ME3xxaICAwKq27kAwAZjNBl8LNmdG2zYd8VYEUfcnhEH3pOhi
d+aAEJUx/M22zUnzlM2CdwdREm99d/BG0gbTz/FoDXo/4LmQNOjZO7JJwhul5Wgh
NOEmyVjEaPyo2iCRBHvQF6lR46F9JoJOWHvUxb5fyeXAe3EuHkO1dJxkOby9L7my
L+N63Yib9JkDal6ox7m449g75b+ZXataY1G88MAHQNEKJKGlrct30oFrfCqxV0pO
EMNtLvbKDHdPZuX/295j2+WMx5fbNg99KWUJohDT+P3oNC60PKZqnfKVyzTtqY24
CWDwmIWzAyjBO1I+lgiFqNrgri7ZJICIjeso1EZsjhp1+N31TzKUT2NaYp1M3JgH
MEv3+EKq0aH3BNzZ5gjo5XylHPHsjilVlI2V9spy6ghylwMdIPrvDzaHwOVvdSW8
KZKOF33XOSsTkXyB+qlCrpP06tNfsqc/9EBXT0w+EPk81wNnNRlETF5tqC1aPWVF
4VOclzWaz1yqs0wGQoi/H/5XbgyHMv/Z9EIjMkkul/bHmnJ1YAJSG8XlwhJSCk96
7dPS2TqhOt3yi61FZTiQ8opmlYrqOj4f/qKlisagTA1tLB7epCRoAinxyIpBXxHn
brZebE6pAtL8HtOttcdEHP+VaJfaEQGC3GX4rcaJsVjHHEjlPVmNWhAXvBn3ZdvB
pRkmJ0srlkZW2Yqy/OAihfdQ0mMs+Pza/KXzl1iAb2Xzj65PGZRn+tUNNNVyjV/c
gisQQV9ICIe80tFNDSk2uc9JXktRcf/0Rab7ruQBFtlrfWqdQW09aLTi95QBP9Vp
MKHq97X9thu2FghKvmxduKNMErcFGJ5fouDixgYXh/cVK3zRn5E+1ykiGVU0CYb9
p5wLGdNPPPN2z4Z61gVTseDbWtgTvVNWhhdHBEnGSiMkKh1mX08JiVriqmwVYtjg
7lNBU5NrnUlJ8SoQxOdmqMoNS+8hYEB8m0V+d2cqSF6qs/iZThCc7Rcx74xvPGH9
uarggZwIJcDFbMG3ZOr36S+aYI0RdeYSBG/RMv1WdZmcYomWzaqWZlpdmruQsBT/
m1/Bz5LmXkRop7sU8Z5JZ05WpugxVFcj1oleNCcfLVXIGOY4t/WpAgrl5xoTplsM
iVIrB7XLqc4Xdz0BQCYEqg0KSkeOVSgFax2qhLvnDHkthymPk+dIe7a5RKb6gWVp
co7+oGV7XUt4HM0c1y8i/+PNRNufBpuPEp5YfDug+NHEh0zUhS4cA8nTntTtannl
cJjmDfkGBgKlsUheLqrLxDMfrxUb8mCY1e0bbyTXcuJTX4WQPqnG0ghkaYVSp8Fn
P376HAyfLT1TwkWgN5QpfqzsPwxAMxu5A3/uhkXEbG0wc7tXDwmsTC9OttK6Z2Ng
IXLnXb25QhtwAkPNgzvit9qJD0liUsN3S+Ksuq0JR/WMkWZJcnngWcpk9F/1AfXn
EbFKx34AOaqvc3yXqP+4EgMT39gN+B6qrHcfEJlMxd+oXOmISnPDri/4Q4MbaeN6
lX8+AcjIPbaILFX0tq/RmQiQ0rDxGQ4dkkci0WgS1e938GL86N0bBJWN+0TvZI1w
EygJo2Qq97VIDwDcSSRHoha4Eqwue1u13fiqqa9i5dA0M9SKYvS+VT5S+VxnXAgl
N42ad7ftKtRn/vPFgpbS+PwmEycyT/BY/Xpiyv2s0NaO+OLSidY/5Qat0ra3X2HJ
BudrAVIsVJL3koBahppUr3p7IsnfjJQk9saLe1ZZgFvAHC7Ps+qlhehEjfyeaC29
PIW4JaIqQ9cs1jdYTwYQLcqjnPF8L3+SDpjlZ+OFqYB7xJ25V7OmoGJgt9Db04P0
gZkdUPPUst28L6BHrLQHj4RN0J5njWohNFPfh+Er2C7MrukkAriPRtcCyNHUHyhU
LHrZLFhqFctf2CT3trHSZqHdkRvyhhIWnnVb/fab+8C/UMNSSHxV5q/5dxyEGchx
gWFxe7qR3Za1SplNrzk0znz8LTl0nmmcuvlplFyKGzS1Yv05ndN8NE8qmDzcI1/X
HwPSc2KP2D97U3oZD/CdWBcgK3tVg9NWTqPXkcuUx/8Bhg4+JvNAh36Rr4QOkA8l
Mjb1a1vkrrQ/il11QhwP9pT+IHkwFA4TUhhZ96nnCAkK4NvDp21rkh4XE0xdyMtD
6NvY+gIA7uCDB7J3qKUkQhfImZdzi32SIB3Q6qCasHQay/fkxYlO/WpPhc1t0BY0
pZojMOThIGsbuM/pgfrERZF/5r56W/nZzLYQqIn2/QxknlxOPS9hbAGGdudODQRJ
XeSGbMoTBXjcdsd0Ta4dnczR/zFjxuAlD7Tu/lmOsjSTD1reQLPGEwjTn7HKCd+p
EfEIvg/dl0VlIYmaqUuE83JhNmb+AzEgrirYz2ykrG4GcAz8FYTpHfjwVDQwzvFb
snaSzTDHHkhZqLHHnbpi3rqVuHkD/pAS4uffXbFaPJqkZi8SiihmROyGP5F5UuxH
uLJYf+FW3zAZgXZZ2Ioq3xB8Zlwh8LlbxrrMEtPC+ZU+UXKG+mOQw8ASf233fCV2
ogK/k4ing6JJDG0MZOBF7NrRu2pFvueAC47FMOFgB9R4VmY1bjeo7TT2e00Q4Hzj
wJhB/sg325owoIRN373LdgT9+jXszn6aoVhr6LZM0S1fGvl6MMahmo+1YUBTpcUh
b6J3RddG/pMohdLTpykPLuaJUv4BwCvNs9Hu7og4I7hqNFG8897CgvGkvA+uEwJj
2m3G5Gst4EcchWMkuyZT9TquySwKuBZYyrtGB8uHVuJYpqkGpUrWbmQbrOeTjDXr
cx8CIGSoVazSyJWuivtClbiOWgxrY0Mi2KZp2SP+xwapjibZmrrGef4x2VzJJT3c
QtQ4He/TKe18mpzl3D2ArgubbgUjY/zIixMd3DdEHZKkpB3uah1ezBV1boeZ1H9S
BJBy/joiWzl84SUl/FTaRBhzMTVi5XP0f51radY6RXSHElgYN/unjej0ORjp8M11
kRWJomVVyMGFzzsz1WNDZZdc92YyjSttAyxrnBjKnCvwPXkF14F8xuNm3uaduW9N
s8MFxDdA3Tnjsh3kzIIAKppsH2gNCwgg0T4HfbL4gLtxkZLHColiUgjGMLjVgaBb
6+/1OtTrY6PMqYnu/Qfd51rOVwcdKb++RQvA8auVpOniA32GV6t6u67FnOm/qADq
4KnqZ2RD6o6lyMW4UlPeL3AeAI4fUsQ8wPidel4jgwxnXcskL9UrkNPNlOfhtiMQ
OiOp87SXUZp2JGPao0J2U9rRn5quaXNSWBsgAS/Ggai5Wh97Iv5KYpXnTNxK/2yz
O7fgABjlXLYV15eElkiWeYJentjcHsDYcGO0F+RjXZ59m414dSIqTMVdV6HwKsLx
HC/Lr+hb5uGyblYWkOuGKtJDbeUvgBBjnDCzvFGo2XXG6NoUfHZlydPLbC1AdAFc
vu7iz61ihO6eJUfBL0ga4Epj3Hj7ZCfwuSR6aSuBzhpDqEl8SVqjRC0sLaZXoHJb
cK0ISZzRPcmvQjG6ThhG5gs33HFWqnl1it8iLKRhbf9E25ROVly8lz9lCQIPaLiz
Fyn/V5biOS8WiPE3ghtVGpEFWrryNz6LvUH5FD0u4ZrJfTjoIMUdh4iuncYBS7xw
xdiZVrN9WaxKR6nSoa17N4NTdAsBvk1KEVQ/lHaMneAHO8bQZXDQpJjcYTN0y6PQ
tyhJRp74cVT5haUylk+YB39XdW+0uv+buHmQycG4wGCd+h0kSZ2Q4ZA1rt2hoDuY
z0StsnDgNcD3D9cgMe4/E3YiDbzbm2xX1RnpFKSsC0UrOKXx2QCtrMUyLE55aeIn
sskHlsGhnZpdSpbs6BEV1VVYSMIVkI7GEoWos0v1I+BQfG2RNmA1EjLRA6easKlO
xGLMh6TgNskK58zd6qmA2hHlLjIsDLaqSTTs94VdAp9QqzLS2Y6VwXt63iqpJVSv
VsWKgd9V7xyP56iuVfply8TZ1j4casqRHThlpuIBeQz2b7TV36/a8d1yKKduUN4t
w0ABlEhrzaIfHsSEsTOR01bSkeR1zXZUFWidQaYmzouY5t83+TfNliyDx3rFo8Bp
Jhj18e6CRshG3GahBVChqMmAnr7ht2oBeVDkMCkHLYgXJ3b4uR0aBH8tdtK5kD89
X1dVk2jpOVSCVjZRH74kgMUNlL1tyZXqe3RyD5fOH2XTXXtoFJNNWiw6kkOM3j1a
v5gAAzE6uVwwzDtuAng+oXXD+5CMxY1foN85hD++e54GlVkWsHmQyHB3P0JLTEG5
5pP6c0MiZBr8kvL5mXaQP6OQUgAlAdohsZ1LNY737tlh6zknzE/laF97I2ZMw3g7
6YNx+SlG8M2yllp61C4JzJLJwZCqdD4JuMibyrjK1USlRTUdcwB3PUGWtMQpnL07
Tk74dyUFsgimodWjQIYHVmDnl/+EPmtuMzM5NJX/fQ79QUNWLF4qT1CMJ9fCVQx+
Wtm8B4521xvW9bI3NcpSjq9whMWyZUkAtMNVcpE232aEc5mswPnYNBpoOk1FuzHl
0kQtVwqo+Ss8qwDbHhoYYW1R0H8zisCCjxmDu3YKU+6IZXa/SDaSd9ZKUTSARwRx
s/PjWHshyKUFIV3KgQf4mmOtRUcC8fdyb/jSMzNskfulFrrXWEXqpqgGxr8aFSww
CB62GKNxk2T6vpbSgaz6vXQjHs80CqIW8PVhp6K9c/1N37jS5PYwnp+/+5NgQ3Aw
ihPK35uyq7OwKkALLjmTPJF/3t3tntlBWNnpVYo/CJlgZ4Oy0KM4oRgE/rHLs4Pm
3LIk5uU8y206itlpZYMvt4a3lGUyHCQgqcWhkfopsGZpgApqKhVQkr5f+jDZOiZw
Rx/e0LKOOga40Pe5XHP7QXgSx4T5xYb43ut2PQAU/593Xe+/K0sHYCmFuEd+b+s9
WtSku2S8FoFZ1nb/VfXKo/L9ojU4bodrC/ISo3JQ6JOlv6ZfrvYmI0IITVHKn6P5
jhtWm9w04V5/3vhVOkFpDOf0oGCyfKB3s/f4X/tZpqfUzzjz0ru98a4Mf+M7k9bM
AVMKn1hsBBOD4I72QfCpzSFaAIKj70OM367fs7LkBTN1f5nvv5UbvWQeA60ftyns
lCxxohdvWnD0egOJ48vGKjAM+pQuJxT5b4n1D18iGkhJF+UXIpGvtwS+hVpDeRwu
y6+VRvvWLVUFvbp0DHUIny3HYHN3g/WX4ZsRD1wXaFccYtCdHu7kqCakJiPYGoNE
nr2pl9qSHDICYN3ek576sGXFXrXLDD8GVUaBIHNy32g/NdUbV+yGx/rNs7Q+v909
eyDgTTdYEYrLh9fHn+BJd3P+flcMZJ/j3QTdc3CBdTIqrCkq+76NvS8KyWudqi6Y
/AC8ofG6oZZMTrhYeqZpbK5QkQzel9ysQpV0PCaVWpmZ5RkXtRp5d4hb4qRZnHA/
d0Lnc8fK+ZYe6rckKXRceEScBx8egZehQ77LpsyBk3gLMeMjpHw+Hg9ScNtDTlQm
YOe60GLFx5y1+kJEQn6Lo51Fv4j1TBFEnZ4tplf3qaJ34qt4NzMnHeakoCPdODpx
sL9EgDSoz6wOBKmQ0teytfE7M/tOMonsQmQonWscHg8g0cRLRCGpxgeMKqT2MEE6
1jjvo3wq5JUerBnFCZtPrYbIgLQMDMOXY5IghGRYHZ3PtqJf9KEJIKr8g+iGMrQu
g6RIyZRtlZ5xiwNSx/ps3+tMaQT+60Fw2x5oKjVq10jMFniwK5U3WmmUwtEYAOp1
gfmTba1DzwZz+pqaJ1my0puLmrD+gm8IlvpEY0DDSaqzW7SmXIEGS8Zjxnid2oP3
Kf5WZluRlaWPBIHagmidFzu6rPly/FPSGS9Eyf9TdVbnng4gFAjFTIM6cUZImnwz
ntI4Eyq6C6wLZ2BFLBdmUctMJopgEJUCsO/+J3vLEJ0OBfikh8AN9HQtKe9eORUr
zGR/yxzmmkcdzWb/qwciOrxt1ESqf50lE+x3Jk+afTPJHEq9t+ELxHtMyonzTVGW
GXttUPFkwtpiidP7O/6KR3M7iakc5o8uxMKBeRXJEHhMKyxwp/XrZWoYqtmQxe3W
DdQmB/oKtJ1rfzBmfH7IvSGAvpyumUDUXFeItgriysTa8AGJ2gm+465qo4oaFE+c
PfMAuajovknSCL6itp7USCKTZOVDbjZxpfxzM172VRIFCWKRWYEiMPrRLWEEce9d
bKblDUOfdz/4gLAq9Zw6cCIrZ/lpVmuCUfpYGONukQZED1WhOeWIxNmJYGuZdHJR
Wnr9lMJ+AxmOwPwAUzQonZHye8HS9b15q+SFL4v0KabGQGnbvfPPKGvS92cKoIPe
hr82kzu8FPJBhDfaV0YcvK/nrQw1VfQFbzgLJojWrM7PbQZU4YsgXdMtt3S1Yg1p
nkLPEd44IxTMOe3Xbpp0ls7UmUHe+wzVGUty5/3WwcDS8gItFRINEFrKBxtg4TBJ
4qXuhnFOw9B6BX4M59lfkxIoH1OrEqyb5ADh/K9CVYy/sg2w49AF3guk2DtaWOB7
ld6sieveEzV5RTxnPyDf5Uuf7sFkax+RoZyyolW52/e9GR4VYCVpwQkny3auiVlP
vwalSrOZfIrHoGU7u83RV6/AsS2grxOVykjzTPlBzRQQOmuzIAQsT+vjteLbMYHR
WcMKj7kBhfjz88954Sw2TjKIvJZq3PTsoQI7Nfv+N43UxzAFl4GP0NllOJJQGWa/
MCzZGPsLJLkeU/8wL0BCtn/ltsPKJ3Ha0i8EORwHzJf4EuKNe57DNcmYpRLzPy6v
JocDMUxXVrH6aWt+wMEAmaxka4wcbqBxXCMu3vAP4gQQTGfVfWbdvGi3EU/TJ/UR
KkNLZ+ck49wsW24EKBsC8h4kzDgpJd0bFVq8d1zUD7I08R2IrmNDdUuhyWZNd0oW
1oUUQKklsN1IiCQdpkRszWuWoFZFkdijIjozFirBxqK6e4ExJardAJNUwcxsob+X
5o+jRH0BIDQc3DVRRs0+Vk1muG2SItIh5QzyO08cd2jbfI1DXf+iL/Eb5h0JBBkp
5KVsVIc2vwBPcvugHWv2jkKChdl3XwLHPDfSeiYOGRMIHLj2m25urBRSc46bLQsP
gfBsGc/xMpFUMV0epHxCSk81f+e5KBvLIi6Z+++KSL/wHcyLQ0QYE12+B5EZX6qN
MV/Mg9fozz9IAbejgxRjIO8ECu+9EifRit4jsX/VoLukeR+7ocfNzMK/B9nf4y+k
gz3lToJTsjl62g8Ta7hygrHRiIwyugMejrLMcZWJLybAjBLhH5G55tSXEsL0KUza
tm3Ucg4c96sZyz51o/BB0PhIv2CUJnJwbf0HvyQtPZVob3Q6Y6k+7wK79HXi8Oip
dUAz3BsAuMcFR4Pcd1Gj7V6p+W1mWPDlU9JiP8XNWCL73n4vAgSOupFwCNP31byu
4an+a5Oyk8mdbTUU+T63qIxnuNkj1tiHsaQ9hLHF3FlEDnNngnxDah1+N/W0ZYw6
hWk49FOlhk9i9RZktBFktYb6f8TIR3Z3rCgKAEMc2ZZLlB+PIqk3uv8WOLLVLRh/
FZeLWstYixzOKmSxthgfQhl4dBb3nkpbOQKfaaXKdhDIVXVUraU0CeFK6Zn1Ld3Q
n8jHWri29FP6wHK3jubRq8Vhr+TctsZ+3kQ+BHzdIR3jRtkaHuUTpnv8YJOat9bf
S/wyoCMhWTzTiVGXdHQgJ0k+LuGYe2B4tQVsleN9VrVFiXQQSMqBChiBvSkpvNPE
Li8Xd2QQzntgsnqS9rNGkTriAhAlkZo6xhVz5ZYPujJB9cWL6jqxMHrN/B1y5GqE
WUEJhVJD+wELpy9t2z+nSJh5sHARH3QQXk6P3/eq3gUsbc6Or+AOpxPoN0Q/uWZN
/qKohOjBC62nYHCF6EFvWAj274WKHTj30UelUFtRSS1mYX6of911nGHaVb/KT0mQ
8rS0hLjMq4ZQKRMopQUJbvKqUI3dC+WouX7XPgPk9Gp15ZEor7GXl6gQbgFfiWMP
nCpu0cS6k7UasQ2uPht3ozROaem/B9H/7XxhQii73eHM+eUa2O3sedI8XKwSOjPB
nXo0L+K4mrkcJfmZ9kJlmHCZ9g3Kc/oaN1mBVylbPOnE4K9Eoo47eHg6BjYtIYPn
DR/IlPhiu/EkbPoDmItDh+IwkS44p4ByuG/vOp/nrTy2XFbGSMnFQ1/ARH86T+7l
1sOOxA4hjhovXtN30GvD11dFF0NWewn0uoVJ2brFqfFAzpnXPMXF68vHpOGNh84l
1r7ZKfSj96CUeCn+2E5IaQ5AgbFbGxZm8afTBZS0N99LICNa4oGTZjpEbOqRziJ4
jQunap3XkG77eEAfRs7QEmZVzXvL8kS9mPlw+BDiuzhv8mm8ak4PG4w3dGuzBl2R
Yu1HvEO7zGyfH8y4oGf7SfD6VyruEg+m8hMAYskG/+BQwkZWBw8erHdLrrT6QU7C
uWt3/nfS6Sznzmus0UtMh1bmA3GP0M4m3bCVDRtcnwtC5Wwo2oeKs6mNv2dbZEYw
pMtpQyKssAQO+BwsV1isThTX5CF5xu/j5nungUrByNxtkqZAnhTW9EpXr9bSPcOQ
OwKV0YT9vcxSlmwVpOaz+ZYSqzAoEoNwiqq3jjuDPkXxcWUgFOAAk/6dZwYxe58m
dTKgowWgNqQAw2vDTVvEEwmpj/GLHPXNdBryJaRYCoq9bomNAR7jzoyj+7KPlpEq
slUfaoClO/7ea8m05W0zjAdjKPoj8eQbc4iKVD3L3u9susDhWqdlRxOevyV20oS7
sn9NHJQTrU7Hyg/zl/tA1BjyaSKxDb1wHDj51yzfxW4z7bFweXUtXENHExqkIjin
t2dgJ/v2s1DINcYCQ6Qy+1DO63y12P3X6L7lh9QYIqEWzLvRKg2YBxIrAloPm3/G
1wL9QKaVThdM166UaMe1wcuuPLugh48lPrJXCKXuJ5kggC6+jXDOZ03C/m4bidLa
2J4Vbzg5vm+yH2DGCmuSrACNuTlMcNTIqkiIQG1SlfVOFyfLCgLdBf5daqeRS641
Lhsqi7C3K0eUHbNbM7x7IjnuISE4OAj3t+D8Kcrz5WtkAC2/A9Kn5HrfbhR0qZ1p
+nWk11lkHwgfsR6/VWXkj4ro1q4ctS2B+bZXZEwMcGh3glSMEfBYYGOZ+xKaFcXP
t3hXDmU5di1SnP65OJ5KykTBM44gZTCY8jLyBxfKoc5WfJlM+hBqY5SEK9QsjluI
vmG1rJFT76Hc3lGNSLT6VTRQEXslgrI4RSHzo+M3GKgkcdVr0k2ln+63iwJ9/1ri
KmPw2ugn2r7dIW1P13v2sVrm1uwOlEbcSENWRCpHn4pPbNAY3MUJQLW+2w3a94vG
btLsI+YfdblS7x2m+EuX2FbgA3RDUmQmhw7Pf3sVTk+DnMqLXDlqc3iw+VfKPn9E
cvmyGQUua0I9epIT1IWfGiRafmk4YfqF1YJzQHJtmzDQpQjRyIys0DEuc8FWVnAh
z4iq8qBc3FY5nOEhmUts4TlYVKNbPILE+q8kFRyPJoZ/voYtoSGEiI22YKxPKu0Y
SqGcgRl0vh7snd1ZNfkv9+3cN7efo+wiDxGvlHLQ93USXnQaUB8PbVtsX+NQcqRz
qa/bAZhqX7FzU1ySabyrapklLLp61fgRMhcWRHfx+zGPb2qqiXTIu3V1VXtMhQus
4BYlrP5otwTlJa3FT7BJb221NwPxO3tJ1wmULlYZNhPCAY17URpnNCToqgJO0AjB
6VL7FojwRPMMcdP91GYC5Eb4C3um4i2I4yViNOtndzJiXwCos4gbF4ucd1O1/Sda
9+ZmZEYJZej7AWkpvXwS/ObFqPjRPcaBjMxtpBi+OCmPaUqIqqrB6bDJUXqPUjkP
Ozq1epn5ZzpUU5uktUYhzCiBdRaz4StTqw4kYhNsYMyVyRh9V/OzLrdqyP22EmtB
7b+hnLP9qZhTvdTv6qwjFylPn0sqJRNfrJUxBapdfZZjMREXhwUUDvYddq2GDkHq
6Hz9dSK3gkoVcnXB8y4ikgk8xPpoSEkuW6Q+gbOkX04Ex2Rayge4j2o+lr+EyDTG
dJ8U2zNakd5xNV50PHIuYyHQEtXpRkx9QPYgLC5hFLCPm6sFL9adIchOec60Hmul
ILTv32x2HAxpaw+vss6iN3xBn4txbXnWKw1kjBg5kXoAMbypQ2P5FGlOLqGq5vEI
Z7pqkN8IB0uSzAtZF3cuIXi0zLSJrdqS8Sn7YrfGDKQpKUWEKfXpdI0+n4BBglSd
/0UPsvtXHFz+c6BgFxGHvv8x5D8cFZWjSfOlNlN06U8LHfB9ZBvAzCptbqyhtqlQ
AP+0TnccV6iD+tnojutesk0Sw3DcfsfFq+MYx22OB5/jhzrY6M6ulscHDRnZKw2I
2sAjKv/qMBJH6v315aI9fNCf/40LrulBrYb8LPtrYnJPBXYwCOVxC/VT+aZGtMDU
c6Hc1iwPLpkngEiTRaVpRshY0G7L4QwukPtTq3pt2dodm3zUDxghAgZ+ZvE6PdG3
2OVSxP46NN3B8wM2an/SMruU++XZRHIdNzWYux0BelzeRMmpCa0h3wwULMzQgOyF
BBq44wmKLQ/gWl9CgHXZjwixDyhJgfjzcXsW9j6rpLK6G3SNqc1M1EdeKSvqzt2/
1u39VJl82h+RUA/9BRuYSzpOSeIt+xskXoAiX6LhGKp39Ovf+IX+8lzVAAU6AKex
1N1+8MUK3Lq5TvMaVk7E3+tVHqnH49B84Yz5epJrdA5iIDtGFnsNFES090rdwkyS
rWlYNSC+kt6UnI0Rq971OnJwmmcfLsAr884d9j2n5wlPC8u1NdbW3OJjfQ4L5NTJ
hcQ+YWdq/amhRxVAfXAhkKSes3m0ymQzwmfD34282t4gRgyFWLMPSIxn+DFq2GFU
mCv8Acn2kSpdr3ncpq8c5zXl/V0JLtjTW1yZfhCult6epcoy+d7zeXC60nBxKi6j
oSiyi1BYES8eSUeWyJCZqbDb2kWEuTcwvx5IE1gvapFaJ9uYbjAU+G0sbzA+ZqzS
QRm7qF4NB5JXm5mAj01j4jwQLjF+Rw3m8ih9HITpPD0UK0fUV77qtrYh+kPgGWSL
5bFtPgPXT3TLkLCEYypHgGCAAJkA8zHZbv/SPpdSWSYF9FDcsLe6uuBC+s66kfJB
tDglw0LomznuAXvPPjUNaOJnhl7sOqoxx03R5aNXltiWQKYphrY15w8wetKLrZMe
guQMlkXzY27uSxr2IegSY2Ke02IV4hNxgt3v1HGMXX3joDzWrAYtlflF+WVQIMlV
vouuY7rZtrBQEx+/JxIoNy1iRwICMi2rdMt7IoiKVVsPpZuAm6vcu0Z4Uglswz5e
+mngawRtXNWqlrmVOM1pgmOR6XyVVymVboXZ3nG18XBthsRbbQ1mF2nruy7UNIWy
AS6D0Uo9bWV1kUIE0+4WUDd8e2N+ACwg/V1TdI0Meup3O1hgRSkkdXq+rUSUtYwt
FhEuPTV18Z357qEwkeFau7qxwOEsTnzNSzGDFQiJ2dP6pLac6la20HBFyZ5tUkka
W0FTFOLX/pF2SMIp4hDgC5puRZG74Z0GjWL/+8c+tM8DBZ7C2x8XV2+CuwWbm2VI
mrAdiHlyvcd26m7lymKuCB/Iaa42DyemL7GbnlWZCfhNWZRg4Aes+iixNprhgGCj
hTxYwnIRflL78gem7FgLPKt4fATqldzt8w8kHyv7C9iakOMJr1aSLIMvILhIJiZ3
/J33Bk0T9sm5IpWtgCNhaxnKzvcnRY52HpZpjdLVBzzAr+QOwfsdHhZKdVik8Apy
hwvKfCzbMHThmVQ6Mdpq5OPsEzGbsxvP69qnH8H3dTpPN6NCvcP8wxdJU6zbBdXC
+8BSM7RnlD7J9YDnHqld3pLezk8iQhY3F1Lfcr4mW1XaL/zwqEkALCZWpUSOVGBC
jiV16jMh21AThKSqSfZmAPXvLFmlZArZX+Sn8rbmsoIgrJdyvJW9Pdfc/KAtK0pn
2YHM1YRDcKsM1EZotJQdYuO70SwKt1Dp3+XYJPkMkffdVmdj7Yio5n9mPG5SbXMl
/oJtMdUgZ/BWnUmIBUmoW/9m0T4ieVN+lOQMgsF9yqXIRLDTJaTL3BWMpK3O4j9F
R3spB3ZfJA2OnXkl4+Itjie7EDY4RheYSCNWm/hOcJGKT7AyKhYhzXsrzux7OjQN
B/irI/EfQ4Rs1A9Y2Fw7MVsjWAq+shnNAppqUmln/aVg7qkJzoXu3Vrb33Se40T/
oWxjT33ZxBmgIpHgyxhVpoexS6oLIpK/ynJGCsotzsolsaTKFR/JM/HDRzWpOlir
tS9APAVU9ZU28/lGZeZVJhqUA9EPjnfitRdXC/bD7kCyEf3X+bJQrEYmrZ0ZKNY8
ZrfrwSYgS0futGumYRY5xz6DftiA9ogHMpv+Dmfypb9Eaam3tRPi+qbpkiScP0IZ
XpKHJQIJtL6LG41y87PityV6iRtbvtPAjrYlmJQI857eQGtctW77rPA/rslf1JPT
aTW4Oeo3fHgMWp7wzYzE9UeIgrSc2sysIgXFGIl15u4/wdlX3+kqBc5VqQzCUlrq
rLYGUZ6LnshrmH5Px9Sne6BrqX0O26wPGFpMS9KfFEoU7eOdsF1BjVLkzzVnT+Ld
xzPcawuyUP+csrrc9cHg7mrfd3T5AGbVK7bbvrv3TDjZYzLd6/Gj7zy5ziHk6niq
2gGQq7nedLUMqF3jIIjO7RPGn21W+P+a8m/Y58WNVBTZclnabFMRPWrJ+kC5UkgF
tdO+uwjAnWk6L3HH5GMJnyW7SFjRWqm3I5kSIvO80n1dPm4Y/Xu0WWJmnu1OkyZZ
mB1GYm+yWuYhSJSWMWRDqZxr9rHZ7yJRGhpoxzibT/m79PMXvbHe8iUsXNvrKoGn
2cDsIO5WWORTVtKOr0sGm8ohxdz6MAvqZsOAgAIp1IcxvvApp2VeAJPxGqu5MJdW
c6ckYWP2X6UMCqsL7JpPJg3k60E7mPHD+7xPNTdc8Z+rneu8EFiEAm7x9XWNpIzR
Bnkx8sW1ayjW/7Fn5bsxDXVuNnfIfG2sARavbwOvkHj2MGoVKgYbDKea2bdWKJPw
mq37XH6TT2PnICELGTLBsm+Cq638jHl0YIlwOEFB4CpRFw1ih7wVkxpH+54Ux6uq
6PsxpXB7u6tw0VrAkOZc4WnzKTub0OMV8EfCiVy/UqZMapDXkQsCynpDkuKUm9iQ
+aKT4ZQw58+Cw5tabeA1t8kENwlRkrSTl92gWV4NRX1W7XaIo6Age03lPXLas9K1
P5b1X/cz5GuORwroWK7z2ZIBa9hIg5jqk1JRIGVqLKTJQN60nVTT0FMutAWJs7ah
shRQKsj8JiDNBXOrxmVFIYaWpCypyjg7sJRWxj7wLwLUkneNO4kA4tpOf7vklMro
7a/pAI6KrayVjt/xzdta0mRSTiiuaGU9c6bFFc6Nj5Hwu7l//qTItEACRI3HoAco
dzduEOqGZHgGUfHw7qnk2Dw0n+d6vBlgZ6K42uYUEl6XvYw1ZbWlYYwLOKyRY3ys
IaK0iutuLEdY8VY3sG/g4GCk5kOB+I59ox2qcDIWm6CAu3mPvoFze8Kc+JY+gD9s
7SlCCP63e6Mb+ZziPKPWe4HRlTD8ckz2VY4EliSzabKH6xyiRyA3AFjtbkIIZreN
Vq6a6lYHknzWBXoz4ujvkb0+jkrdC9xUArbZ69FJklGj1qHZyjMbW3zRFfWdNAhA
I2PQDKEiD8dAvLoD5JQraOOamnDAZj9DBQxCcWXsaZfgQpdu6t/zw6yV4wAbNd/G
SuPrkwf1lOF9vyfHN4K1e91WeYmbQuAxzPDipz92Au14cf6dGvQpTWjJ3wGvsi0+
glLtYgPYckb6bayHjqy/IgaUyz/6CMfEnRkzUJ9XiGkihn8VwR+5WK846R4dMbu2
DiwE8DyICW1N5adx/S4yZcT6zxstuM6wv6LZUe2Qz1qEIW8ZzyeCOxPgwz8uyxMg
GWfFI0mep3naJiNqtzioYMkTVszcxAHqX4wWfPn020MPIiBDqk49gBnfssvMaixz
cBc73Lm9RTvCbbTN/RBo/JY0vjg3qlMMIvUABKdxn7XrPtYU/s50+R01hAlm9HSU
/3UcGHKY9NTBYuwU2jg5GDmtRt6pzbyV4Oq/3Yzp0sGQlyczZzsw1Z0h3wxVTuvg
Zt9fAIy0PqdxJwV92TQUufy7XTFLLCnbNgc7d0MlFv0d+Wc+7QjBAFErEf6qqrVb
dQp6bP2joGUGtZz9CI/H2V8d7x2Xy3D03owxOLF3knUHu2IXxXBKlTRaBFOB8wqC
w5aq9xJSJtg5xyNu/O2i2DY8rD5ttqn60kpf8lvIpPWut3B3aENA4PvlFx8k0Xha
AcRJLAAHKJtXKjqpQytXeA7dxAzwvi+pPCx/1FtkiylsYEbXEONjkwd4sN7tyCsJ
Ar+DLU4r9C3GmeqzWuWJGPUotBg+GyZ7j5EpuDwZZ8xErO7nCmi2/csZQVWtUoMG
/bkfjSrfYfDY+/g98AS+SNQSjH80uMQE4vdu6pMOFxj/DftkahgHhOHwDsg2SRd8
hCTAa7T4RKGa1/QMGN5Xecp0Gr5Lv7MIcYXlWv7WFtl5c+kE9W4QZfSxvLiInBbx
9eWbQSPe4oe+YLaXkjn6YlbVGr6Y44GksD22UN/8RCW3Fg4/41C7mN0l/H3w24Vd
LAx7S2mWjTfykHpuW+CTTNojb54eG8DQDZw/tMqp2mmz4N8x1pcf1I0wF8ObhuKw
Bb25CgLNA0mIEHbl6lnOhiugCu8UN1H3EoYWrstGYnEpYhL73ABpvI+JjRu0+EfQ
OydLSYClINKjQ3QVGq4KpRKMZt98zHVMw1Xjpbp91TDfa2xYw2rUtGJfQnIc3lTf
+rcW1x/nzk//DWac5QLDBMBcjr4T+R7GWeoEZY9sQfpdvZRmiLp1+jHFGZZAmmAX
AkvdwTz7oN1tNLLiN8XISb20epOIB1pAPQSGHt3Gnq+/udN8jS9UuKT3nViqS0Xu
yOquQNXJlGkMuDUWrUZ4Xitul40n6BIjwoTYWd0Wwpk+Km+RYGQWK7/MqOdmb6cp
hJbodrfci81mNhHgO+RGyjl04kj79jCVeIcp54YLfWJgv9XVLnxMCOl0LgFVd4NF
FTAUCtN2r6ipz9qxM3LjMA6g5nJlv8a6NjoJq7VeA/A23Qv7BVlb/yMcDJ8Ipk55
8ue1PMynBohv9nOZJoprlct5Vj2jiMjFxNz8POTy+fAcXKIq3UUTTp59+HYg4WBi
BS07eQ4BNbpCxCWtXzEy3Ymhw1W7sVQorsMe1oHSgAnP7U6esOdI8OQX9KfB2ZoR
Hp8gnMMi4AsdF0FdUz1VVbdyQzQN7vZ57nMaLbfMGhvk5DN6G5uE0wZ1yyQkWmtF
WRJKcssL14p+GW/5rqhkvincrrOH2Oia8u8VCuZjese9pZGYhtpgeIvS+7EMEPxN
WclI0KmMqNOSDW9jadoRiBUB1TCiPZ9hFJ3ur4ZOk9fU8atsvRG1TD2R0wC5+sra
Eiaiw2TlC/HiNY4aNZojdwAeeOMlO+nMk1hdJewqngtLGu0isfJxlOM3Zbc8+LHA
iSrgi8NpAZyZofKjtMo8xOZyPU4Ftn0tmF4L/ROoVZtTVrCnICLTpJI4eu2K76IF
2mYKVnN7185l3/ZGXAZN8GYIhIUTo6PKwZ3l/SrjUquaIbwzMixtZri2+JRJWgqd
i45sHoiZqXPy/5yyHYIzk5usZe8opFXwAmH0nMhohdczqfRrcxuuwfYnG0IQQ8BW
VHfT8ba+ozC1zykPomB8Rku/dCR8oANDka9EunTQpvc1pb/X9spWmCEyyKv1zgao
HanQ6HTUt6wfn0Uz9oc/ZDYGiMt4xFmZFgFcj1g2QTuFSCZsPolxHDkh8Fcg15yJ
bs2OZGF9OYdB4WlRxIJCS8rwb8x9UBM9x6Fr0QYyqH7RkbWDwOmXNKmoMgv7v0s0
lb0EgeFpbQ5FFn7cxkvuQRrW+lm5NttpDWdWdAfOJzkYlM6RxKLd7uuMIeNIkBqc
kNSUMOuWJxKojnvulAriMY06XVAhqxvXjUutede2a/Loq6Kpm7J1MI7cVT+0G1BY
dDkqbMBAu6JCSMbf7O+OT2MBRMSEH4yBYr2ZpSwV3B7Ba6KdORKufm0kpb7Bner0
TrSEIt7OkrI54HaHo1i0hWfkn4RQEBtqVcWTUQSlO9I+GgHU2Nv0jq9dOH+40aUA
BNFDdJ1s2KFPKulrbckPxl9I489IOblPOnh5uzwQg8ykZy2HnO7qSe+hrooxBHNU
hYiOfEMv/LboR3pC806wvPClMSnD+aCMGipV6rfuhKFHI9Ei9YDf4tuZw/T6zBQq
NmoQxNKOrWYKGTWTK9XF4iSI+GndNnHlJApUUfc1vmpoqxtk6zAgHUacz2u/x7f/
GKfE06BxnQVZZG+yblAUa4DZZSWHOCFyZYu3BOrq0YBHLDaQJW4zdpZN5Dboj2tU
ne37VdtkC29Dng15QHOuPY5cr4RE7e+udKt3fHAASqffvE8Zy+lJ6VYWiDqXwnAF
76+FdQ45Gb5z1X4rEFvkgxpMXTD5n/FOUF53+YfULpGvc9BYNQmMK7jG2T0xysbL
FHKSKSaXv5iRHpPoqSOo5OGkcn8IiBb3+BESiUr4OcCwBzlWq/hCSbLLkfvMso9F
YDtjBaQEgTzaQoby6vV8MzdGqMtbVyKU0rp9/i/4MEWA7e1lc6lFAP3a6VIzPINt
KFseijd4ARsmqQdpcoxkPfyppZ5ulP7v0Q3f33GBe4TxgjZcAC+qwwTR27MLP3hA
BJdVXDbfKyG+O4QfJoTmui1fS5FL50ZJNt94gY5gdojRH7AYzP3ll5Vg+RnNh4K9
gbqkzzZggnJVDbZbetzx33J3IEfRRXaltg9zgAWAZD8esswFPauNgZqyl3PDT2f3
C/5oQQ61CEmoQrihxAG+Z1F/cLEdgi0arK2IGjR92mefrdECufWkSS7iRGcFAho0
1oEN6dw4GT7hUU1xh6C4Nn8rgs4bd1vFDoZPfsNT+fpd5UUXE9kJzcm4XptHpaLH
XdPeLsnzGwmzgskqpLpM7zQ9oyFg6xKoNQhTueHM3e8gNAl0Uq8WDBEJk+9QH4Ab
OBB2RKnqw04+4imKsptw3aQSRO8rTPxFT5bQYwCfVE7K/nDwa5uNlIrxzyg2dlBx
QcM596m/Jhk/1p9HOnMXYyCVAzXAk8A/LVV2XNBllOn/yev7vai2PQABcBWB8wnv
oR5s9B7UsurAN9igeoAcoTsfdlCCsU7o3E4NhO2Z7t8XTIDKdTKK/EF0uhu70z+l
dUMssyFo1xCV5awaWmL5FfaYsH7DicVd1AP8vUNTNTcUJ2fsq78yEXRG0buJveAF
VIlMAmsNw/sFGsgUsMyEqlWRHJW2nH1PTyMNX4PCxjd3nQM3X1OCxURpDFSC63CM
sXzNu4oVD7S0THHIyYIiUx459HB6I7gqzSVpZa3Ipec6H0cUsb7MuhWoqVGtZqSE
wqy2QCpsQNQC25G0nUkHm3ZPYh4soTV0OvQSfjA5eemUjcwSxOT7Q934686sPKox
nPnI2ejeAEx9ed838kyRjEYvKMr531QUumzdqaeq31kmgDT2f58Wli9b7X1iwm2q
0SixjeJqOzW+Io38o4P0E+vr7gyf1M3Kiu0ta0617JX7Q+BCODgZkp/D2brylU0B
C/1/ekWp/R966WFLPjxYI7TAQ1hIdrB/7KQc7KL13+0GxXh5OvKkFXqQ24Mc9YEA
xKbWs/vCkiGL5Harp3bIhfk6MWWbVBwcCo5RyC3/cFAaik+KkCte9zhxRwDmYYJr
4nR+WgD/bilHoDYsAiRtVMri9w3jcnF2xlHttKfgv8UUxh/1ovxpRxWX6DRcWgXz
4iDQg5GrZk/zVQSO0wtfaIKK7p0FhETu/zCQrplrAi9pCAASHZNBnVgG+ARgWrJm
wzLhaOomvpnsnqZiIDPUWxWec+Wny+/M9mi5Ahjvi9/8bSkq3nB7CFHKS0wY7RXT
pLLcHRJGiHi4wteFSo8N8XCUtcHkiKP2DbFZJjky9Uh5h22CUiH06FnfE4zakfLs
s9bTJcRSopYAmpMcrpxC9mdIDG+wWE2JsRasBwSjVxqbZSk0Lnwgvf03TW+RCJyu
VBBysOSLqCkJLopQdFsAoTi+SYMKdwUYD5PelkzRYP1c5o3JV4BqplonmzGHJFzP
PO7ntkqhqL4bYpkRIUyCkOJNG0BveSHWqJ5UAs3AqyLkW4hq+a5c6TWU6yKoCuCJ
NIi9jtFtcJAIPa6A4KUihvSVrnoZZgtHqZeF5uyO36xCbcMUdoQ5Qv84nzGLhiVR
AtSmm+wJb67EyIn6MY45FUFVcHTUHlcLwRIy2xkcP52DIjIKdOgyKbu7N0V66lbS
nVzlbP7jWms0LjVPlaGT8BX0qppg/iFx66Eip4MVUkzsFO2JazvlsI9mcwfas8TK
fJPohhqNwkpTphmpzCs+JxqCzawZCrBXCcmGX8vcRfQQ9ytLIokxTrAKDcCXxomR
tYb0s/jsmRmqWR0QF0noAiLScal0lCSJQQQU3A/7sVSYHgb1fooUX0P8UdixuCdX
TSCsD1Y3WtHq3wuq1b0vTn//y5yDS0FcIcqo6qYcBAbHoB/uvJ43FlhJFFn2R808
wKJ5W36Yyfsm9qgIyBaqIliA+wCpA4MOhzeSxYovg7BkwCbsjT37WE9lnFEwUe95
DE0yBxSHfyfWUkwyC89PpaePGjKvik5OMbMuXv7WZ/7Oy9/v7D9TxXcffDhaEmmk
7uHCoNJyZg/rmpXLO6DDyykclYMmizbnmZ894kZdDKO1SLFdk+Hdt3yK2DH9wAJR
YyOAC1MfPjjUJqX35o/aAgXHL5PEvLo0uXzOQVz71fJmj3+zyeo2UzRvqlf69dZ3
b3VDo78s7Xz4pWjaJ0PFW5p4Yj2/BSjCpMqVsLNf2HQgquPowZo0KaiNm+5rhPol
zbZiP+iAwUjC5KjH4F9+gBMrxfvn8MkJNGahl3J3lct6m1dTiDPE1SeE/EqiqmYh
EqzYwTs+rGylXnUnxPXzIIO07edX2rdsgVdXFBbYXw8ZO49wNEuBqCbs/41amSsG
3dw4zUifV2VDynqg7joG3oUERU3qbSDPSFzBOigsy2EAsC8chTwFgkfUVrgTjZpL
Z5uuaZhOvjh0nAbnQ+XUX8hak2JtVThwzJ2FFaTRDv1nx2KDmYcLb24cNc6vcPKA
USLGOBRSGVRecNw7t1HJ8eTR8YCKoxz+1LbV/biSOUFyMVNJLpTo29d+/JEJCtKM
EPPdCuBLu4dmjRELbW3qy3ObdL24cKqnANnkRRRLN3xz//I6jumsf6RwxzFd4f8P
LLFKhKgY8miEZiRWj+h08ZDrZYMpHquSOSE0cZklA/tNIDzZUZMbOpQfoa3c+OJy
L49oy5/m4OaxZqhHkyZVvrzvL387ryj5qu3hZeR7lbm0MPDqZab0FUuOTC7rD7FW
yGs08Tzqq4xaqPdk01YwnJt2qTp6JqfENqlgh/U3awUaECFsnIWw3gJc+Od1QoF0
psTiFJsSPSJwYkDIMpcelp8gU1OG2Qwfh+eDk+JnHmeQ2E9StKlRiakGFnHy+wzU
E2oxJRbhTCmR7BbooCo8xtCuXnweZRLarseF7NHd2tWHRxwlo8P7nUSOnUCxeK7R
Aog9APqRr9sYvr/sJbx7mVO3manKBQKU1pk4i8LYOsIr8vaHi4nvg9ZNHIKpNH1m
ZgkgEr50IdkUag0SGYGenTtKG8IPfXZPeXQMfJdjtswLgqo2FtYp5rlM2bXrX1BA
5ZVxYSmv1sjJKWt9dWnCpArMb73T1L05tNvCu0GrOGrzPz3ZXb+hP2LKwf1MreiX
1HgQrdhtylwrOzp02b/65SBqUGfbq0riAC8l3XnyJAX6DBO8WG0lzczwTXyLIdP3
fEpTB65xcDuhD5sj0wol3ykeIFpQOPMSDuAy72cYCQrhNy+RjcYgaT5xc0dxKvQf
3SGklbkuWF6yab+RaiPqKvrKCJsS7ZYFba+wlOgIsyxx/47+3k4S9302cTT9hZ/L
1H9iqYiM7/Q60jaF6FU0uqzpk8JpRnxN9kZDrvsds3N9mS78lPxWw3qq3FseJAmG
NrGOFSQfLkjkLJ5YCuLuN3sQ7OK1ejN1rryMipwLFY1exe39YtdqUSvWXzJbT974
cj79DtPjbsefcd6R8e/6ExWsHr3p/Wqn0JlJf6A1BA9/PhhmpCpvI4Npxg2nCq9V
YZtOxmLg6vkd/742veCXRD2JTf6F3RGPNqtM9IWAzZ0Ruc94ntYcVaGAI52rPdm2
cChlDiSNV26WRSJ86MmOJ56iRnlslZf4KlbpVyCkJX+cd9ZnUwvLJ0e4Y2K7s4AY
xhiFiC96/3BG31turG+sbUmHM+tsfIIPqJHt3QqasA+dvJZ6ZGsd11+qtLIsKkWo
BWQOHgWfbcfQ1NsRLEkXeyC9Z8+xAA1hsf2Q1JOfGtHtdHRqX6uYu+VTXTQ6xcGa
/bIaUJUnbaevPB+Zrrz/HoJl4AS0dmKQE8opl14YMGuT1xEL2olICt1TWrg7qaU8
HBSUZKU8D6rzvyd28sepajomaM5e5oy2Unvrbi6z7GaOgYptScz9/WIe7M1a7Lzt
ZRKrtEd6PCgoeTawRLBr11+3VD3rSMOFM6pizjYvyFVyXGtWvmpCV6PF+ZshEyun
Sg49AMcMAcNytolB3+Q+E6TCx4POqOt2F/RfmBSyBCIfBOY5VqaZe+NwRN1lhkDL
47oFVRRXbH0zM8rUWz/AyE9L07yhGphtyP4F4hL/LiYOU9oAGVX1dxNUnqR7++pG
LaNuRtbQqAZj8fVGNA7xx/VbBbqXLIGZk26B1LUW6e+l0xtBux11im1VVH6OJJ4a
XnzkvzgLLOCfT0ojuG5pzgxT+7NuYX5/xXZEAlXlh3vb6vqlC5FyCjLwI4549VXb
KLQMq3Ke33jOG5EkZmAb/A4LRPS8DenGWvQKD3rk/i18UY7ZhZwvEI/HjFr7U6Pz
qPJAle7JFMiiNE+GtbAovpMF3iqbf/JyLdZgTj9dXJmGXQC+pKTK+9Rx4I27T7yj
+hV/bGoSmM5s2L9MtAo3KJVpxs4wNjYvcdadku5WiPb7NGE1FoOPSAHew21hYFKd
miuhM3gD1C8jNz/G4BFCqlbJ2KkIKpLyPTRvrLYGZt714uX++iQnxMF0XBMkTMZF
9rAV2St+h7vo93l7nDPY1fjim4ha4qJjO51MTPDLSyoQID6wx7p738g9S1uXNnoe
/Px6VO2RtcVbYsPcpJsW8cQV0rD9G0zGsdE/m4Rn3xGoSKJYDcpII9dtqvE3EJvo
d7eqlAa1FcR2dNm5ce/CU+uPfKlf4FzdpF8fSQiR7V+Zvg5RJcPmfp9iUnFVFpXx
BgYzUdE+WJdb0B6Iq0yeRnhrpHt0lwp8I/oekVPqdqSdXdkL4sK16E9unITMgDgB
RM4UnEEYKNOMO42vhMx2Yw9cF5PtbJAuV4dd5HTYR9Ogjlkx9NKTSWBgEih7j7F7
GX3uupm8IGCSfqEstE4Pjcykhy0eRdL306bJt5VaAmfMf2DVtuJoSp49PSV0a1XH
FBG+rvQbUZEgd2OWS3/TcqqAhd0Nb4eynsZ2j8DKwAip78dQ6j5KddogvCNhFGcY
MjxunTUT19SPffpofiqz7eTGII4ifw8MBLf4LfiaCeP0WNoiFZLyDKEZyBFaN9J2
p7DRdERcP24dGk3reDFb4aAKugg4fQoVYDCl0W+nk0YaayCAFjKUAsdjgX4jQY4X
+hilKP8SNvZUv19vj9I+XOqg/4Pr8dFsInPWwhyESlKI6uY8TuMsO+GhZb+ozGEe
DHVWur7uMLWpaYz4scikWCr9zLi6WPcn2nFkjD0c1eRfxFEklUR840YP+FE2h9jO
GnQaytk7skR5WB9EzbwAnOtleUytthfpDJEBs1WvpODqzBtcZALxBQxnICkwxwGj
B63ZFhfJM5sCyG9w+EOzemLm8Abx5pQf5vNnbUSD1Z1Z2Gx4/D9W7LEuPRURfOhx
bhvuLuOisSS15I8GndDAUU4jvBuBwrAJip8U+1iGgz5EIowL1rMIry5m6NtlREJS
CRTQyv18lNPk+QFOfUnx9q4H66k+yK/N8NY6O0ywxO4+TnQLol2s0aWS9VFTzk9Z
9/g9+bLIDU+rF63wQIaIRY5JImtl1Rn2uXQeLME/EisuE84DLItKco/H2AajW95L
QCDXImW9xP4uXbLc3AQ4hXtAhxNU/+Vuuf852WsgFgZdTrLXdLDRZGqhBK3kgpqi
agHN6KADvAve9Gux7IV8pk3c5SpaGt7QNL/RfSuE/k9BE55zyeECS9YZ/FCCBEzV
un9ZQU9HnMZ83cXUe0tZAQzViqGLk2eL6JUIv5R0NFeb/5UZBPGHoI6JwFf5RH8L
O/QwRowNr3a+wSu8woFZ5xb5PRPTog03zDGMpIwP0RW/9YOVhka8kXg22dveMVk6
183DQcMEuefbanJBa6wC1PsTY6Jkb72m41UfYawLtXwH4YL0Xi2xvwLphRqwLyE7
FJdKvD/YkKP1kYZg8wd7xvQS9chKr93fW6V27AjuFAiQWotco6fptemtF1ccrp0q
ZJjAmhFgCBCdk2E/HjG8BPS8UiHZx5UfG6bDRrx1CqJVp7n2sFZYnk9wK1XEirrp
ao8SNoKf2UXL/cwpt/OEwIGgjOaHq7/28YFaxCutnLrcDKA3/1brArQCSZCeJX4W
5ISZ/xYoc+UH89Oq8ADqvzCxY08I3jfJzR4XhjjB2DhmTR5NT02U5eR41KzLeMyS
KPy+wJElPFj5teHjpvnj67SWRrO7Pb9cnxRofdCv21RzlsQ5RbmvQIxiubv575gp
RzfmDWH4qCA7Y8NhF8njlbCmEntHTfd4N+U6+SVkcanwszpAUnf5K8F1qzE0nJTE
W0hvK14ox9ysIZ8BVH3tm6QRkD3COJ92DZ6Fq4sm7CkrCo2f9wdamDQKd5Qy4/bi
fvgPXtHi5ya++2e58WmLlmqjNUssR7deYfe9YAEZUPHUA/++zXPinKmfa1dIdH96
gn2X3Y1DTEcYYxYkfAwLC54Rjo29ScQwbG/kejLV8/DLgck1QQDqFftdCXOuzflC
4gd9+oGqWvSQvLoALlkI4IMryQmWaO8H9pJfJo0dEgHiKkEFxnhPimzT/QAXpjPu
btWLY6rdPlkjirXNvJJzrqK68X7FTEM7bmnJ1jR1QdtoqZ0Rqik4VN4yUB+Vc/4q
J2WpasgtKR8i8zmslR1pSwr4lFA1kXsIdfLO/IFKLg8iL4I+gmEPh7ozgwT1NLmq
dxJGcGuKmw7dFIjMCxZq37zmpoTeOuk7QeSNeBqnHR3t0Kdh0cxff5Cowkjz1oSo
hDIvcOdO/NqJUzk+ScSFPvfbH8byeE3dVFwG1K5wDB/r7DXIgOr65JRAl1zKqLak
QkDRXpx2RDWjh4ANSahfZ7MslSR6KC8qqqtguhMy8267wXmp9j49k4HcNlVNO58a
pb1UDeXvjnzrfRm5EJVPOUoF6EG5hZhu78F+dJtb4YvAo+43hJwIgTu+te839H7T
2G7AcusNWgqKW20wkXwI1Ot6dWxRWkZIAUi69cRMbPS5v8+VZF7va9YZAXnGtxT1
M6BE8/qZ976RHfdNAF3lM5QWV2WOXyKGLTDHpeDeb0Cs6uNm1nBZFwpkkj7KnmEc
1z0zxfHhdbsDSazMUufd3qJL/ODMcdrQhcM/FEQK3nYfOJzGfmgVVFL0SkBXt2Gz
qnIdgnt3tU0CcvHwqQpmml+Kcl/gcsPWJ5KAUJULk5upAr87m0HWS/oBUsK1CDl0
UtlHge7ypF/3SJEUYElycSgYohO5c5m70Hbr3HimFGdfm1UqXBu9WLKjb+gA5/x3
SJLUbHHFBlisTzxGfYEH7qoMuiTmV3e07sUmjUkqKB9YLePvrdnBBEoqYKEh1CO1
Bq9uF3jQ2OD2ai5FcfTwSEK7pj/uWiabww/I34PlfeeHoD4sTwUj5NPtYGHu12WZ
jR0D37a7TbN00F527QmCrOroBpw0B/NUed5Tg0PpLHdTr/n+MRjIVR0mEBU13kM5
NvJKnZmfngHZuheC5QpJcW9x4CDMb3j4APqjEFo5XAPSQ+YNsKjuzPGfUH/r2ryT
h0cQ2hgVC9OKbq5PIeEkHSoXN5sCHdVsWn+1r2am9HaWSLqKqbzcEkUXD5+roDYB
QX/B2qoFu/Tqx+1mEnVe/RnN1VsQXajfEUZ0SrrhppvfFwNgpYQprQjAg5KuRAg3
PscDyTy3hVpYbXyTeH3lk8HhF3GnoPXF3vpHFkLLOCHmoMdUnYQUcJFiJRgoC3/W
SvRNS3usH8/tDtqKZipkVfjvNoRPATXguQPa0hxTpSxhf+w8dh8vsPjRZDvI1mhH
/V7QGYDmAMfJeeb3vTbsuCTr0zmCz+PoQp4cuWPOrui6+HPck3zEIpH/EosHF/xE
dL13pUSnvuTEhYRKvSpyVH1DrT/TdSJFT1VGpckyZvontAswTlSVKGb4gxVhtSJw
DSdSWI+ObpqGKeyySstmm6KSC3Br70LPw19sMmk2P/hJ9Kp6H/gpFcXVwPXffgM5
KH/1WAWzKX+lHAIPhOGHsvweqx990Ye8OGpPErJmVqESnog8S/p9NqfL7FdKLLpp
81cQHGoWbkG9thR4JHAGVQB77tabiL0Ii5Tihb8nyYZZX3JqOBf0r2/X8g8i3wVi
d238XPr845Ani9VoXT3d7WXQeHj79nAQONHUVN6NCUsUPCpXQ4N92Lkhkltvv96b
P+C4gyuwcbh5MmpvPW/+s0Aj23K2XCZRSl3fJasU4asT+txlz3CjeQITtKrBTXks
FTE04FakjH3Ip0XDX5/XuFutcojtShNMfg5dGB2Qi7myEir0che8N365UjTYKKs5
zRnCLkm9IpmHaRJvxjQKenDnP2bn2SdfnSXVZtD+bdvzw+gd4g95uRdkbhn/Rj3C
dS3ttL+ohz4elBIF2bnnQJ0IiZIOkRy9Ytg1Emd7b64wRzOOULrJe+ZkftqaImEj
M3kjfAgenkrz9sZ3MpRFFO/AlRAW+c9CcOIyYt/tmo/PdD0qrf3cvyHEVHTy/9xb
8JaCHmdYDsJjTBW3S7sYsaFHCBYbWiYuITb5WwTuTwewuqSshNBsGAC2O227vgSC
HhyVyNFUB689Ls/f8a8kxeo/5+8UvSxNbPRNUyJVSZWRDx3ZYRdfcdeBw/XvmP48
QJ+MTJ0wZGqhhEX+RUC79PaA/CsI/Cw5eRy9GHNm6Ozno0qwvjDTZaPDz6L+lHjd
9v3Gv6YuMhCUKmKti9Tj1I+1E+O4HHzFpuXjny5LvevO1xOuUttsKNFCLyln71R4
WYENa3GjkeaC0V55pxJgIUz7NC+7Up6AWKf+kSAIGXCrfrxieEqSFCcpMLp337qZ
cxnVCK8zuINM0FD42kWj4Tgt3/3CHrgMrF8lS4+mdHzfOkKl28LBZE9/K/3KNrj1
p0IFFnmcfS2CdzraeR3BALR5s/JsWt2VEMbyX/TuSHYfOQxR6LO+OUEjwjRRdBxv
dpX3lvddF/EIQ1zKOcNovjJB+8VmihTyE4jFsJO8Gr4Cltg3apT8+sTgfB/z0P7u
6KkT9PhzxtzXhWLefYsQWGAxkkIwyxbbHBgYjjmM2FJ4iLfxOlfLP8WKvDIGwzt1
R5Yw9YAE6S+CrZI35iajAFt90PFoc1vweu+gEoeT6y1RGlMsO72yAk34A/bkEElO
A9iGIj1e2qFhQ/ApdjCI3RbeExuux7WFtPnac0KAAs8b4UWq1tHEXfGLQnsNidVF
YyMunIlBbbe4ABMZV3TSaknb+fjztiALliY6FMhzGcuD9+NJ0xyhOBD4RgwVnX28
VayArwWbyzokbPL+XbvabkJ4Nb2yid3LuWPybd3UBXavnevPvukQQZTpZzFZCc25
+4BWmCbGFtqqoXiuzmK7YLuNzmHyU6nzCRphmJx5xhRdzb3P80IktEmJd1nRmOic
zmnB5jFdYabVI5k3Jw5PCfapMKxcazzUYQmJn43uycs5FQbx1WVQLH+HdZYUYoDi
4dTedfePE1DNdyyB5xpRQ7SPwJ6Sl8TDsz3VacK7XppDB8zwZJ6kSPHvesF5lO0+
yITmvYBJrJKR79ph5n97QkatkB/kDJ5Q0UtzRWWDT+p+KcWuLJRp3EnJ/K9eITaI
CUDO4JpAsaMCjCQ/FuBMyLm8QN6OEBDtrhIHg8sVzDXgPZ35Dafx+B1Keh1UZARe
K3TYzioiuUAiIlg3a4pl9hLyPB6/EPgDMrY4roV7Osyj+znXYdvZHfPuIRGL9cPn
mY0iLgK3hrW6e3kZ5sPCOZ3chhPc3Ks61+h8xlC/EcKIeTRIuU+Gne4D5sno4HxW
FdTI4JyMz0S0FkuZ6tsbAZh+gxtmCc0DGmZ3ZFDc8Q30fJYKffjoOCbOD9TXtqLh
9OypupWhdPlye3k7grhZa2ws4Q1EMOxM/0y7TZyxwVzkncfiU4d4E9dfpVGv4ipx
C6n+Npc/wBb1sWbFQx5jR+/t1Wpbq/84gpniUdGrmAmQaaD/B6AzLI/yQyZvnf9n
XqlbdVK8toJVv7JR6Psafsno2phkGXkcIjZOtsE4aIfp99bgH/5Kc+GoGNuAvR6W
q0m2w7Y3pGx2FGssIqc22N4juVFXNRZmKRUsEaB64OZBCvmXFYKMFPonYSTCLudZ
uNW8Sh4wT/PLZXM4p2zWCXYa8B4EVQhUXSs9KUNKCB0P0dJTswaAwJ7MRni0gkjw
tlanLk/B9Yl3WGQYhifE5AhqxvUgjHdj+0BjbmcsqpTAVfjXXY41/A3wUL0ivXqE
mIwAvcRCTG0Nmsg0ejZKo40Lj+dFAuj3BMwnBIuofwAQ6Fk3Rgoei/sFl819ASFQ
RsScU/DES7WP/jUzoXolSDRKCxEbpIa5gIGEBbMcE1s70p7Hjax/373u4CgbL+CY
iVAyAuJ3QNWx5aE4GERpbn/7IbDRm2aNwFdSW3zoPYteFIRxvlF3qjpZYQsHsBOa
Ec4izDyAs9/JuH2AVt4KZtDF5guNu5TydRdbWc1pe/Jpylrd9uz7m2bszp+iWDiW
sjI7s6ZpxDaYOXOzxRJ5U5Dy75lbc+YkzarYI/ZdXdhe51eFNK8Run4xF3B1KRm0
Nt2Drpudfc58V4rz7US/MqX2070+2jybAMxK7SfsAsid6l60YTdWzPweABaONq0F
wRxbyb6293BsubLMNd3Aq/isKAclwef7eqD/5hcekcMUcukQMmaQGveGhgAw7Xj9
sAZBxz6oujaoKHRAqFLf6TAaSl1TrKeFEKL/rIL7c2uNUfGc6209N7+QwudkKXZx
acCRfd5bz+GLaZ1QIs8INnEaOpYzXS7KbwMf/uLiGjURzp7NHwePQyWNNBGb26bt
TExuJSD1QoSevqNysrt+NizACkxqUUJfJir4brkdxvKlnXWlII6QHXVVceFzLtrX
jponKamQsrtu1ITiBYaTrdg5NiBRDoeSXfy6kM2RbHn5DyswXtGFn2hooX7UuZFW
ZKGtJ/7Ynld1w96Qwn3RlwpJrzS3GtS6xFmijOCVMegKQFugdCG3nVeXbMemlPjK
MkzMQp3sve4zjrEQkUkOGc/6OjZ2/Z6WyMFpByTTcErjgL9eMh9g3qaCYlNFMfOV
L2W0d9VnhNvVD/t0BlCKv7oEs1xqzsvcHQTtklsaASKCD69ZSURuj7CH1jiuD9k8
YOPWr1cVAwkoUfF6v1G9QtVPLoNaY5YVzQefeyaZbDGdwGO4K92cAVajM5gzu4Cm
yAqKhZKVk9T90dfMHI8sS0NmrT4PRFNklFr0Eie42ysu1ttQVCKb/WQCs93zEmzW
HAww/OJEeDiIateHupz/P1l8c8g7MZEP7SXwOyPeneTVxnU4vsUprHGNejVZzJ6t
LmVu9g7Wxzcj8DtB1sKNAgUg/UGHsSyibkN1Kwgs5RgUqNtZlc8uDpLFhK8+E8Ps
qOty7qBBaJMQcb/mTZx67MzTxJy+gXEDUOrBx+eyHbBUxAlssciMi9cUefdxcO+R
mjqcp9xsIpz5yNC6jUAwwhvcww+vgZl/wxa9+Miq+Dc8VD5RGkhfJLe0Kwz2a91A
+sglrQbJ1vQDB8rFKejqiRlXmTg0+EEI4RPFYksAdZ7OPRWrTcUPpZAUr8SUdf6H
q3z1ilAs2yk9WgiSUkuK+f2ARzzPqDL2uDfcb0Jaz2J1Qbad3y3XYbo8GocSLXdw
BzPWF52IU5jmCEjzyBP//gCgU1FV3sTzl/i2ameO//aHyQjtZ28Ca+YS3Kw+MWsh
x8LmZpyIpz9iy7SgjNDiNuK+hogNjVORwvzsCQwazszR/T5FUNHkt43zoTDy8WES
rvicUFsDer+voYiuwlA1ZzHMaq4hx0KBZBJAdTAV9MNnNQUPCHlODek9X2y56TRB
oeD4iq3JjvQfs7ojPnLrpAI8/MNh/RpR9ebeETORM7sNyXfHEHM/p4CUG3AM2H7b
XV0CkhIVWo4BWj+P1jwJemCQqWrk9or8U/sV6QWe1mtWNHnMnrTeoOxoDBxUWGaD
xC18a5vjSWZ1+MLD01nHFXw1LZHS/VzjFq0Vva/PkFnsKBUvR7oer5zYWRR+6rpr
fwhs71HY1KFFJ8v2mN6U123Ghpf8r3zaht/IGGBgYrk2hthoOG9yk6IKZ7kOziSV
cJtgJxtJXVkHVK2l6Te7GYqZmEMRi6vPZ8s/p6ipC/WcY6BXlv6qRfZ458c/56Q9
zvGpVThEy7eaXvT7aW3AamXKPNYAiszkzpbsu/6nYBNYlYrU+WAzQlNBeLLq9irw
47cx4XCSytPePPPO2ueGUXy0wZp8JvFXOyyW9EeBuHYPNv2atQBfntC28UcdJvY9
KQTnVq0FmwAtqRILgojco0T71RFjtkRYVQSoIydhKfyvMHwR2zPn929pohwPPw/a
gV3uwHicOcqsjjyeo0qgqf2vBtpOSlTRCbo6KHINMAsPOdIX2IDJjEWsFlenp3yD
y4on9YlOPzhgXZ9OpLWadFM3tQEIBofxI09+gt2jRZyRaOkI6GcRMem1KoI8fQgS
TEpQD48XWglEYk5P/8khVQ7CWJ1/01qjrOh3xQVLUm4zgpkqR2tTkUV00bwjmL07
WkNm5FU7gUaCc7Pz0Jpx3w4GgQfa0S5OpszUoM0Ot02dqFY2BukNBCIhuHyg2FH+
Fg9tpTDq/cNIZ7DeAM1XEUtyLwoGuscQic/9tiZlfNczH/8TdEiyMSM3oUlPx2wX
wVXaQuauQg1sz2NMlqz9lJbnAGvPjtdYsHy2HNpIugG3N4d8XCW2jLgVqPiwdxlC
o3ziES6A9bnDWKYF2k8OPiDZrbDnwXs2KGTFf+3R7C1hvmshb4EtsjZ+jG45CYQB
Y1KDUdmeqdaAi4z2qgx6cR48rPBLJZJBPlH1sk2Wdg69WPOaS6UNFIqaljf9RfYw
q9gj1+Baym3UOWqsRFf1dvSQCsGpB/QBAumsYmNxtoF5obz0sLaZ4nPvk5zVKnyQ
FoZwH1p/34xFWUCR/OsfSXWyWfxq3CV13fR1sQHh3ywzJpah6FJ8GU4kbQsGeYKS
rQ0siK1rXy9DnknxtAfiiRtrwFV60eXVnwLGPso5fmH+iKYv8KYmX2AYpVMcz09A
ArBHsJL2QCJU72GiKXfXtJATTND8VEiDTguUNG5WSxJLG7Y7RuyQ4GQRnEVVsmjq
kwWaIQ7gHhTB3/F8deM62WcrldvhG3+uSs58wvQ85GGmWi+uWW9wNuYL4qCPHeKQ
fEzeDVnkaoSmgZVgaI1iz/ESPa84mC4ZHV9Ft6hKSqZ/qaAiio0zwjNgfyxJyT+N
wgKBb8LEsXcfOPtu3pdNyiQUKPp+2KyG2aoFWfOi/EW2xwEzMxBM/CM7i5MZ44VD
B64tXAdAHq0XiuLDJYTHD8CW4E0yTdFwdorgc6GH2XgbJEHVH/gCkaF44EAecyP9
6RArA5vlXUC5eEhwE8lSnjxfUzz8pxjDt5tsd0XDdi1WfNz1HQ4B2MDlZ2zPwMwc
PeoKWCDFPYcxrKk4aL15HozlxjjCby0e9gKgn9HTgb6x8DJODRE861yP4gBnii6N
2iypvGTEzh+WggMoXFaME9Itnw0MNzjSyneyk+Wu953JnV96fz/wOHgwD212IfvX
f0vTzygPqNXbWQrd68KZRoSF1ozCCo20pKr7R1pt2JWHcu9kS7VJ5mtSGjXWi3BN
fa/Yd7aGHf41RDh98f6NlnEA74XiyVihVnpIhseuqZAP6B2DLvPuBXPqTWVnzQG1
OLypjX+VIdT1e82qscdlWZLn5eo0rznQ5iFsYMV237vKoU4bVTvixyj9hh+GT/zq
HataEermYAPaMHlj2SiWrDLnMOYe10m0kqGB6yTFJI5qM2rTF4PI+nbK9gLrN2l9
j95YXCLXH4fPqHHjDoO5js8OHpPONUKRmBMtaWBOwOqZ9X4stKsO9SzjCnHskbQz
noW9dShfmuha0zMYb6oIj7axBvvvSPSxMDFa9qnt42kKErFrXHKW5qJaSCt6hbXh
MvMjopb1QZrJS6QAZZuDTT0EE0dx5KGE3VOtiZjng1UyHMU9eXCyjF+xZgeHZfEB
HaWyWtxPAUuOXgEu6njDFLGEW10ktfSNQ4BdiZRLNn8eQxKjUJcivFSOxlVnqDok
HtwJpiTIPYvlSDT60a03/EkGlVXEZxNIiZ/8AQA8hjlGKEf0i7sxc1dXpY1FCsTN
f+xTRpnDJNzzrVjP8z3o3rlxCwCwysga5/xRxVzVLUsv76OP+5e5gxY/y1yCNFGC
fEPFZ++xZKqbpyrMKRSDo3g6EZJwnvv+niM6r22yCFOsHeaU5qL/M076Jxsz25WA
Ks9H+NYHq/KZvJdFatJTTcu6IKWrAE4/sRNRJWvU3+A2nSbBNJniiwUMF45gCE6U
wo8ptwzP2vLzBt/0I495anmmG6GYFte01fTW1QEpzsSxCOXDMG8m608jTLpdsH6s
30bKClBs2eVnglIegvP20UzicfoJp3UhW4g8/If+9XOfKYu3bKy8D7ViIsyTaYQF
dfCwzIuYh5wxgiZZEGzGatR6DXjzkVERDNcExd93fPVeE4y+EcNjoRqC9/+cgeSI
ttL87AHWMWNWRuHzPlcvE7XIG6/DXofVQWNYCLyED68ut4mHzY1j7eGlBb1KaA/H
d2+TsOWmqW+DJReGHpBQ5KvSOiVOev/OM6wnLgVZmj0X7sVSoWhPl9azRmZlwWjV
t/7E1wVdS1OcZcS7PWWXudXapSUjo5d+uiXyUEMKb3bdrRjR6ffOO4oeUFup2Bav
lxDOEpXWOy0yWvMDk4chQXBC2ISW+hMEp4QqvahaWF+beqm/eA4j1J7Tbhp3EHR0
T2W+QQUoDiQ7kaQvlDWDQgcSTIbkXNVJwtQyN20fQERD1LCng5nejq8eXKC8X3X8
nSSndm+JyVRgNzTjLjeefEzjMfJZPRamoGZ7Qn/9AfcFlHdvLh0DOL5/YuNEdroL
w6c+j+x7a3SAHDe5yxOqPn9FVTW3/vs6e61oDidboWRddQfOc7HPJ0+8yu/HjO3q
Lls+UQgBfBQODKJ7Eiwd3clfF9s2OaTeTwhVomzWF2MsLaUA6mhl02zAEbvHzBZ5
8JMFu5VulAVroSuW8A560UgP+S3aILk94IUhmnkVzoV4MIWjG4XjVa8vKrXB5o6Z
asQgFohLebVg8RL83tBuAISnFpxQLpW/mkAriKaM9mREVksOLrPTSzDveRbXuvoH
QanFK1QsnCnfzzGW51V+nsuc3wF5JGIj9CyHd/ei77ObfilMxTHNXMSOv+tIi7Zw
jV/xW5gMPsFt9TzdxvaXLrxvPLVdGqCgUtbcLTzKfbPyjjcaK/Zz4KGNbyICIaUY
+ty/QxMUr7Kw0ZbyYD5Fz2QW5LgQagbMuYGCBLNJ7yszf8PCBFC/fdm+QXjL3dcu
N5DBilvYRcYfPqp+dT7aB4kAPYqbJ+Q8tjPEnrTzpKO/9c45X7XOXI2kA50BnpQn
38Y8z2l1O7xN/zEG585K7VrvRLqcA1LN3auYOx5x7qvaNeUZOiK3yaF2OWvITBuO
veK3JIdnv4QrhDMGBsxBT3/uKAl/ZAKJDvbUVaamyE2WQbTHAepyFqLmu05P46Q8
bsn1FuuMef00ea6fgZwtLyvfS1FcerK12jqQ6oUn5R1bPns3K1ay8TXS/VQCQ2D0
IP0MEzy+XpeVOKSmkFlixQh/tG02EBFUv1OKqQKh8pQx4iL7ebyhOgTuuill6ArX
efIQoL1vsyrisuw6sYVVgkD+PksRERMxhl/SpqKMJEyoSKnngm0QNiBHY7lzn2G1
+X1xWaMdvZQSz3LDNUdmyZqIiNWqXCIdlhN7y51RfNxr48NHGK3/2DakXlJ5DeTN
afOFMBwgx202z1RLK+Ew14MEm2g8peut7cszxhjXf3tjqjPFj+KFJOU/dxJkojlr
pCHd7EdcBrQXQD27n0n6j7bjSZlRIZYXMFaS742QLu7XqGH9K0mDnAHj1FirqoEv
cVd065mGzhJQx3vryWlPxd7gdH3gAcwciRHFby+5d99sjJhg1v00JxMtXnRqjhu7
hTugwf3paDszmzKkK+y5cm8l6TVWbdIKb7vaN3dRV7gpEDINey9ZwGTLoX+3LhRC
FSJgXgv4tZWkYj/EsvUOIdfCjb2omkk9gkYWQfpMLxfrupI1RQBvAfmVreivqRbV
HqwhBNQCOcYldFH/TF7lwlL59H181c7tgb+Dri5JRxwB0KMLif68iPWADEunMW6t
jLSIFFaT8x9tYaJsAGTDcL0aBIiRzVtrcmGdwUnhSXIU/dO7R5l0B7Zga5jIfHmo
HlK8BVZXx9L4qGDqWFLMltG3W9nAmkwlkrUyX5BiHkAokajuMQUClXCV4AlxwnRj
7p62Zuw89voTgUSbSztADGrTmsMP2s6tmOwEz6RBWp4dszdong4NWedMCvmu5Ub4
+0E2/2/+IYChICJMKgxLElQWKaPBGeN8oilgM33Tm6FFD2W9wNcIfMPB0aBTSrlj
OSkgiBXJvnY6e9GzrLU00ukE6g6e8fgif7B6PB9D7EtVgzAM4WTFkxkQsh9BhXMh
ysTk7/ZdeCQp7xbhvA06yNY45In5HsbTQWG3v1dWIWOpwX2QeTDT55sE2coHajx+
U/nVvPWKcxr6xZjZk5L9hWVrPCFYNCQMdWwQUDepsETz/neYMvKWzBuQ3JuH0Pun
ZYA6PNFATB0DXlKv+ldNGvgyb12vSwoXvZbIGE5AaoisPhT+BJWv5Bb/WsDVDUzP
BdAH+A45gnGUqFghCoNKX56L0tMYW6GpdyW+Ubi5bi/d212atXRKheYuAUp9WSKW
87ShijyZyjQuHCcvj764m+D6rG8KhIfNhgnmNLOrGFtsYHX1L7mZ41898Rjy+SAg
nsYYAjEaPhysTTXGIKlixLifjD7hNFYz4notKbmm1sAZ6CvHVXkeoJB4Cydrvzhh
n9ozl6VhjHEORxaBKCKDCcpOKB49rEMYMtJWGf7qW3TgNEjKrkpmhuruFkALbPcl
bMuHC3yz5byfCDUWPS2vrvYd0pjvpmzPC9N2BeN9NnRIriSTuACXSsDO9VSEgQEU
VfeZjt9fzlyZzK6x9oUSUO9m1i2Lp2YrHbwKFTRk01JJ2Hmm8Hkhc0xsomlVSdx7
R2nlHnNqcb/3lC95OvBuB7JbYiDZwAaYRTZQS1grmzZg+sDNdZd8ozX7ENQOOod3
UmlSfKLMjcvP2RTgDkIkPTOLRMn+IVulDY2MB6gikqj69OYjlS2C02x1Fbyy6FRq
M4uKom7uP41SsWrC+WeHtZ6OS6hYxy7unpiM/RsvY+24I2F3UpiSPVox1F10k0c+
Aum/Vv4bbAivuEMw4DaBqDxVWfBL/VEZ4LbPB+a0qfUDELiDeYyp2m7hDxVMthfo
NZv4+Sg8TEk8jsAEomeKi9NFwq3Sv4ko1ZdoIj7T6S73UfP/U73emr/urcaLWKLh
sRpQFC5X9ipFfswUVWxPiICEdd/00Q10zNEHx95Yugtk4SI31gnfpENRJJv0pqvu
gDmQTW35t1nSjSjqYB1fQl6p8DzCfDdNXf5r7BWt4YyVyyqaPbmr8pp90QUo34Yh
T4sakTByFiV9GPbLfwiAu+o2f+YXLxTgWZL0T1Te/Njyz7Z5MU9McMH4T1sQtKr+
ggXUZcOYdYXzScKata2YBkwwsvc6wAsf0sJVLnT/3mZL1N1ueSGXnMHioR2Nwjgb
Z1SxlSDG4gFlcqDfwdMKeodHMaxy9DxGalbs3MI5dJR9qWwo0crXhhTbWYv27GP4
VQRiDDndlXOhw7rBoYQTuRDFM1Wq8/qid6F1wd3xv4x84bZSUeJaZL5vWCvmtp/k
9ggqEYhEv+K73dUR62ySFxNS02GFeKecjHirGmWHxhptkfMh1IdjvC2/Q3TQWy5V
7OID6DM3xSEzbgQfEGADQkDXrw0Kw142hWajDWVv68+evRaODk4o92DXamOl1OGa
E1ugg7VxCC3Pa6s20RTqwPDhdF5gzCnqqZtph+I7sCW1Sqo0jL2yf+4eojlBEko+
MEd1GGNGU1ybuqMkkjHS74/uw078vUWUnbmIfsc5T83G3Co+A0y2yWZp8p6v/exw
6fwkFm8cRhdFZ9OB4ByvELjV1cSWTB+qOTCcVidJe4LTVHejJjBysieddTrpMUM/
krsA3Qlk8AmLaglh9TPqpeGamCND+Z4BJHDSOHg6txHzM/NErLfgy8joqVrccu6p
jTgZKsa9H8eLOxqgaNTEg0WNQ4D0n11V8C9R7k7+ON4PhTMmuCkYTX8N4O3W9JZB
gybCRWColcCi/8/4O17fvYbQ7Sv1zeHqI5PbBLrPI5eCDAVKAHxcJqzccuUcGzv1
cCIEkUxPQixahG5VIoLwyc9xtUeLvkD6VykyepNNHFYwtjbJxlgiK66tMyg9GlC2
mbcw1SVbozMgOmtvDBykhyzJQtmZQf/3SsiqFRa9Zr+wHDq5yyqjO+f7M+yWa9Xy
Bci6Q6Q+RTJiDp2D9TWQ6qSBwADfUyc966MqCuIc01OBObDSsxubMNDHMwkpRe0s
WttzOsONHwnSbuOouIAK9xybuarfFUaE33vCMBOxqCPQBoFar3bVEzMmJ7X10BV2
MwqPGOurmsC/KBrlzGc6n9k4dpotU5XB/FxIEY1M0KLa9fBxAEK5MjplakA+BsDI
DkhUw927hdvKjLqH3VAg48Jr4bXi9YrcxcjZXFQQGya8Si3ktukmtRrVlFA/Lm4W
SLF3lL/aKIlK3Fs7laKqZud5S3qBxUA9nKSKQLLGB+BU2WjmNejIgBrqMBEu8fQv
BiqIwCH6gyCEw3Og8sAoP08MJboA76dgGdMux0ol0yxm1K8Qtj880RUvApwqwrec
LfpvBrQQLqxO8/FIB+MZO+EEsqaZ6C4aGCgYFPtH/YjNWmfkG0cgSKmpgVs2ZE0O
ZGSN+TYGzO1z40lwL6P5g8bsr88xOSN11LpuQwGjjP7mXhciXekfwBooxCwtE/lr
qHI8XJRzPh3XgBWvOOTzrpiLvXwCjMHyFBMYfWEgK0Kdh3hY69LwLT1Kp1Dt1TII
2B4m3uKs3Ul3SBgfQ5zNToWXrPAJh1aSXtHzq+xnm787eR5DoohlQLRWhkVWCygD
FhN4LG59uiybg8QbhDn04FDC1psDFjEBEf5wMxnvWVZqJPjzh0fhjFLCmJSWLPtJ
kFyyPpoPeFkqLSi3ayxcBWljpaXCCG8BvT4IOKcxFLytbp7TMw0vuE3MbkA/v7/E
q12JOy2eKKRlgQGv7Tn0qqFqqtXCu2GmatjNT8VpXbbryELdky+t9XzsjOXz/oaX
b+RWAxJ9LOl+yC/zVMy2V/7U+TFvwRjKviR1AtwWQsq9aR6IM0gr+zb7rL6u7sVj
OSsjQtFEyEIs+S0dFL0e7X8bfroMAHOZgq+83f63UItfzTvQ4IBbCWrYAbr/v5yk
P5HWORu5prLZhaSxu8mmdfso2ZycCu4bNSbFPdx/j/isjFyVj9YULZzCnbdGgT3H
jSHjMM+2I/aqwP/iNite/uNwDpj6o9wG1JiL4OlkBD8W5Lc6XyYIvtGz2HR1vI45
zBeQ3KBpMVZs7KcS+GY9B92nJ0W5taoW+cY0Stfn5p0UHxnPrKXgTooYq6YhNFAe
eAloEf22EywrTtoW2a8sCPoK89nv0U3xFi2m4rzk2pLYeBw5JPHWV83A0nDPvRCD
V2naDJnSUlD5/N222bZWa0KbVaSEQwMlFi6oosDAykJk1UYS7wUReJj8DWPAqj+U
twdFhQ5RtL4uKd+mTK4316/9AVXbyVuBnCdEHk1uposKErqBHbMRl1SQwBWd8qkB
rv38JH+dAAnZUhIO0jbaNYTTGp+JTsMmy8p7Awku9AB8FPBMOc/w2SIcgRUOeDim
g1NcvSD606HvfNDjUijdJMUrgh+yMalQcXeV/4gCLM5gjPwdFOTAWDRZjqa+6biN
hoISM95EGPptJPXCQSpCvPa+730mAv0IGC75s0gZ2yjjrAP4cquLJP5OMoWtg+Lt
BTxNBRNooLcWU/VbQ1xOJfKmyw7X/lFbODdsRwGug4KNRbUktXPjt6w+zFnc+2kA
LLJGBKovqOlOkdMl3uN7I1EXDy6JBOi86K8gO2/VfX1PwI4pm17xMHGHU0vzxZcf
HbLwbkLzK6Vu2sfRABIOBt7iW9tZaYoTu9nxPy1bmlPQKG7XQQx/ic6f4bxm7mwy
RElqpgrBFVkA6J3O3T2kqoaso7mxBGXc3vtvCC0vQst0NMbLO9LZ5Xis5EJfEfIF
MiaExTjr8yMbv+09oDyM7w/SzTZduWbKL3sydoG4AasZRL4HwFMjXGJlg0dfdqlr
j3IP1GIYec3YDBUgJfbKvXWSF5c5e8rdrc93fXKhW6hZuZXx/vim3bnC6tVfRnsH
6YezuZiM1T1p0bqOfAS8t70zmlsapDOHPGScM+iWB5ndPULWfkXNrAlI56vdBl+X
Z6K/wVorlcPwmPTm9uhFljI0BJo6rdMaf4Bq7TZntP1EbRXoYKkGX8qqHiXD3ZFx
D3SrhFiENMUGi7EwqxxyeHLwhUkDWXxQUVaptIrdT+pdei8+JCv7wwHMSuvLExBl
nwga5ZKWj4u1JucqUNR7KJKqCKj8F/jnFuLaXeMqyN+UFWtBjrVNWqMDByjSkafS
CdMvzeJWkuefpvO5gc+m46QyzMgos7tU/sfeM2zGQUsqZ8CtJTBmYQGgL3n0AriX
TtHcBlKERoVcb36PY59RU5T/scYE1QjaOKd3BMAJhMYEdnKHaeKXqWmm8J0q1p2B
dYdGCELWMqqQmPYUCk0TrCNwb2c0JDYesNSMVXtYSLcmORR7I79hysYU/PF+1wzk
msH2aqIoFkFN4A6MvmyzIQ/X2xMwMp0Zpgo4Cn8rPwv7uyfE1GIz5euLsvnZ7gNF
pDLK5Q4swsX3d9P5d/ncgWZERx4gNbdtLoPhbFrvCjCfyOYYMj3IhvpXLcnOiwQ2
p/w75j08lrbA+Oc+BOtI9dG44I2hq1vyGRvjZR/MmlQGJzWdM+MAXu8dTZ/HD7UK
Ad+0jiBSHrw8uGG2W+BKyh3bRbcjZzdLsb/4U5JCQW3D23RT8/Hbp+VdwxDwf/Kl
47brJXI5FuPdtfaE8Q5ONJ8rngv13SDIThBRfDKJGceShnwhHoUc0E6yFJNNfKHV
DBQDqHEyn7FuUdXRg6VsxPq3wnVLh7TrYvihP2AOC8ctyyn9umEuHk1U0Epu7xR0
N6ObIdfMcjjZZPe8Uuf01hAwZ+9W1TiUeXqKVfY4HMRZnw5WCCssORCda1JSK6VB
Mz50tsPi5rmt1QLGiTD0VPIWkP++XPo9Yt8vGZe20jfafTNxDpeA2GZQSDB5zeaQ
Lcnjam2zAqPZmtYNMTEbtBLvLyAMVNdZ7JtJLgVpHddCZwewGKNBL19qk4+oXscJ
wjBsB2u6AQgRI0+/I1NqCIQdAvSG4LdKEM7XJjrTtrnvFyC7WJyNGsB9omU4Kbxb
dDQ84P95ikENCrB0K1druIclUZpCasHpgdtb7trTRkGNplyaBtcwbmn9r5ivDeha
3vPZr9/o8oVqGCuUKgWlLA8T4mKZe92LUBe1DBFLL19Z9dSmgOFvP8QjqlNSZMiI
dHZoR2kjNgGMXKBSiGIoCjZo2lgmnshvp/PrPq+6moOMDZX+zyuMwVZ1Smm7JGDC
RPZNmz9gTYqFfGY3oulG5nTZ66tWbypxlxOclAlWFzRDUVP5uIC15JG/I0lU38sV
OBR1X4AGYDSd6Pgl7qew8stuk3z9MgrhbjhD+fV+LUEuJM240x2VZlfLrIqRn8+5
2YjvJ0J2uMh8VXCP6KspVfbU5KkLTv2kx7kh/5ktbgEreYDbWoJL/nF/gLHUuAH1
mBPZmbArHN8PCYuaVV8EttQjsDqQ3z+1zVitGZxzhvKXJhOLSOs55AT3h5ia8i99
aLBN+Gl5Ijgej89UV1xdX46fUhM0CgQ1U32HjjtWLRhk1IFSp8vJXRMhs8DxLSEQ
vfJr6WSRQsXu2ZC7F7bNLVUp7xmnI4pUdEosykKsxG4aGb91jm0NBI462axR7gwA
UqfTWB2vK2XRgtJSTUUWYjiCnxUI4NOBonk28NEJUupPdu9FBNAsPfCJS/6Hbz20
VImpe1jPHOk05Gdd4a7YxFOFrn8MhKFRb/3g9hAfZ6nPXE7YwlmLynvWnDRWxoWe
IqNfWLoRSN4TWhpci+7C8P32kklsy2MWmixPJDs2BQyNQBhND+Mkq7eZ64VUTbD+
HChsqC/mXrg+S1xi38/omXSHN5TD0FCVABNUSCqNxZ2Nf27ihykFBVCm+sf/UzFg
rCHLmcBBWSV5rPg8XAe4MpmE/TFZjGXjlIOTIaf3J1sh1fUCWcINVsD+sxsQKp1C
MOzxBR7hCaHISS4t8fDFoNAxYmaBXiuoznjOM8s631wkarY5l54ejtFyrtHprZld
xtILKy/sQKdfBHSy8QspQz+0sE2E8BePc2cnAdOLCZa5ADsI0N39FVyvVg4KO6Lq
+kUigBs6/BqNeH+dfiF9mzxApKz5mbQf/jIsj5fYwXkEJ6jUDty9Z4qhNMDJCBoU
fGJ+c5kJKtphamdLQwa5HzFEh8UEBMKlz2prs6bUASICSPAE2FaAj7CY22i+3FV4
SATGpalEx2xI/f/X+A5Mp+6PjZ+tLCWv9P+UN0jegpTdxrUSQeqixlaQr1aLv2c6
Ygl3kj7h1M/OthOAh9erSMJImZXc7whdLX/7d74LDSOtJNzKoGnHea/6z5kxStPp
6u2SzlSHFAlkrooGuTJAel0RzkM0s7St7OXOdEk+6uKn2OxZu8rmNACsI3hstwXU
mLl4sbIzYYxTC/xUglJ/OHvs1Q+ZLe+FGX1DWMrD9wqvmCTzHoq67jmeCLwKIj6T
2Lbk9Ekmoy3hijdP4/tmHjGViPYp9O9aIT7+fLMmMSmvQVl6+rmdULf0sN+Oqaf6
2hWFnAD0/xIYA2pUWbipehHTSTb+pjbHBGu7YlB0fUPbrAjkad+rHFqkBuw72L93
XoOc7opeZvh1tZ6G4rYF9le1rrI86LJuoG0JsAIZVEPXKgaFf5/DsZMDWLx+oaNy
HKY3QVGshyjR0j0p7SGsz3c5+F4J25vR3EjMv73XjdBp7hfjIp0pG1lZLflnkvBE
pt8TWFNx23Cp7PXzF7NqUcH27gwHCyCtdVOhP4SQ2fiac1/o6bR37FK7++EQxLVF
we4shPfycL0loYgomKLulvD5JQBdru5ccMZ/2EBiF/r+c/7gFUoAKECgLcy0Oh+I
dS8u4+DLm12DvK20W8SQZ75f3FXVW4hi2ziJ7yHmCKv4iyq5QdpD0D+OSKelkoid
Ubw9o3C33tMAnoY/ABAnsqlwBOVyrbNvBULDs/wEP5U14k2uZPP5J5UQVjvlwxUC
4KBp6n7N2+8W5VWzTvfp0n41Ok+k2q7Z4pT1AfqZbrWyGNwq95S1QCwPYPjhj8kK
qhgwDSRNNc/jFHEDfhqzcUqPGXdTsrWBGOZo2mnXerlQ9+127AxTkJjpRaCJX4yl
O1LV+1pkNQx/hgjuDGcaB8xPj6KUg9AyJkwA4lQ8hbSkbgNJj36m5WtmYPiY7ebB
weRYJbrOsSLktcrRkEF4/03udAVtMyPs8EgltsDk2lfK2attWzL0U9liIOxmMU3x
ecyL1WL+jxapInDw23zgczm9Zd1ol2KHfBZuJe9zaKse2xbzrwXbweFCWtRI6QtX
aeqZDve6sVxmla22BLbFUum8s86ClN3GH+BJ9y7ZzUavUs7iTscxuAXp8I0011Q0
0W9KW9iRW62pWR+6vQovNEbfPmVf2RnDYOw+neURDkslo2TsKQU8KU0j8fRSMYPK
ZtSh7+p3Ui6NfxtzlnNCoIxOFv+ZuYknwYqyQgCxsJ2lWF5wR70bL2KAC8oHDBNz
aWQ510nLPd7pZZinAo55CheC1AAzy2Gn0/BDMauU/tOolhTdBNkbpmj9Ooy5TcBF
6tN+sPD9bHW34B4Z35TZoUpnsSGuQnt6+VM/x3/1ptJUC2YoIsNQQqBu6uXSi/QW
xJ0w2Bnd9C+JLIG84qL58zcDDj3E3h3tsx8R0AGM7cMfiFZ1TG83xXyTCUal12FQ
nRXcHDJX4VHUzDGK2tViQSXqiqvDNJdpIzxEbUPWqRwEZmmGfvVLVjCWAipgttin
AMqQnViOjGMIlDzbZP5OKSI51PUbg9PKNAWekGg4+1ptgksq5YsBP+iN5bHGRw3k
Gnsx3hMKDACIb1emVlQ/Q8CT4S3hPoXsRnV6zbJJXAabUeXDSlSix+ydZc1V1eSP
Fe25Ax95eC3Tk5fYH4WtqaC6536demLmn9C0OAehOFkU+G0Cgq2J39ByYGU9TGb7
WUnPNkQ1yh7gEEGQCjBDqhcNQaOaOUCONpXWTq1mt2DvTIzNG7LPtA7CLHxuhq/e
evhNj42njtpXBkRfsSWq8LNWHTToXpnjI9ZSIk85Z0Bl8fiOyZJ/sXUmL94/rsp4
vwEI2VOuDsvXjW1bx5+iCjgTyG9NAK5rzfMcZG8FIl7Qo/F1/rEyUM4j/Bmw7BGm
x6Par1/F01WmJ56OjCwnjl9FbruEB6+Umr1FvC1h+DqW5j9E2NyYSYVl+JV8R+uP
xqIMgJCuMudsf1FKNJTo0S7xR9DNgWcexiPpXs3BFccQLhV+1X0XZcoGk20GIBX7
EMyOxMmqZyaC4AzocnAl5YGlLH0BCnlKSUheHxOHHbA3ZOK8aAFQNBFua0Vd5F59
jZ7jhQq9NY8T2w0P4N44uG8HgL599yKEL10o1jgELRI2QueNfZsPfoV27n74mRc7
3BjnIyIdHlzYBvSNTLV5ORWj2bn13MK5ntmbakk7s7aYSSlp9sQKOBdDmC5VkrZZ
ZgbA1jEI1M+J9VpFqgUgAYc15b9w2DsTpj5gFRWiGSBNZBkwHRS8VzQ/iqC6EQ2D
r2ZiJkMKVhAc+4I+SOuOUOs1yT0pgYLxlUHlB9L0GrwsAgYaonxF7byE2n/w9Yge
7JajsZqoeRqmbjB5qZy9M+b1M3qqOwsCdbduk/enbxSnHaDItAov5HizWg6p54lx
gkVFCzV3t5+aPlxhAzsm01CAlLx+eUhZzW2SATdXVCfIvf0PTxoHXflint29c4DD
EELvvJcZf/Do1c9vAHLy2i2e0cyMEwAy8nadeb4Lqgi5G9wobwLeNA2OyR6etMx8
hcmg8pLw7TupE2S1pviKALOIL5iWGo+qYTgum1wHjos2hQCzbYMeyPVqxCaEr+CL
UKXnMM+4OeOoS4H0ykdG7nmLf+k/G535RGUsJEAtRV5EdN3gkweVpPQr5TafJ/WI
GvmhmYhY+AwiOJ28pjECsuPNCWpH3r6/An+J/cVsb+dUvWAukf1P/LPz3NEAL5GY
vsShgi5zUOPvvz8+QEA+Esubrf9M8K3iXSmssPt5bylbDJMIp2b1zMHLo38t3Toj
b7VKf4yBfy+aF45M4YBYPeAGJF5FmE3OUUt+MFx2SK2XvMrYNcpMZQgI5xUAC5/C
d6gyS/LXMZwVYOCqHvQ+2VqbDDqCvgwEkcAw4MJz3mGMkf2GR+PgH4+rLzXTP9CS
ouZIVAS/CTUcKpLkrvHEGkc5UfF0vL20K5kS7x50eg8txJu5+H21NZGor7crvNbx
iFax1zI0HBLZQ/u+SzvZzjZAVTa5bX0wZ6wv8GVdRBe1sI5iYK27hvzYRWg4xHlW
TwoVG4ezsOxuLRKXKL6mx7jMrAFq/AA4FSlE9PcfOwPwk3KXvHjqh+9i9zfZVs2z
bPn1IhnbagfSMZj2WxSMx1TtPtQULHzz5zsIalhqoDJ07SeYaNfZQgybQMaHx7wx
nZ+XAOd0wgpZqVte1rohOq53M8UPJcLP0PExxWKutmBwHzXh6l2DA2ahoFnng2OX
FDtRNiBT4ktYCySV+HpS8gs15fKjBvHWgsif0XC93utkWGO1nIBmpX5MXId5reX0
XSB5kAkcQ38epcCcAsSCsVQoVSIGGKDArMbpLytlIEFihzoaxzORuQUSSfNO+jp/
0PG8KX6ekvOcG76AXCHq0uVHJ49i06EyoeaIe+2IRJV3ZnF71rfh9pcIPF+QDR/h
fe8cUYM6IIaSu5buIEAyDcoVTQeJHlkGrK439n0DwWrRDe2ie1WeHLdHx4+EwiJN
MTsqJtrW6hbvl49MNizJCbNLRmwpEVAHXHO8YkAJwRH/qdkHTR3ZDQ/iFqAxNdwG
5myYe0Fqt0RVDH5KubdduP2O8jKfVIM8eiNe+JBEG/EUyrkdrBSDvtv+lDJw92QM
K5DblCIJgQU0pMIUm4wKXVhZGP0n+CITsCYX7d6IXIFdL0sgSO1AaFnTdWxQOBlU
U747tGIDD+GckdHy10RXWNtw19/bYF0IrjJitI4txcXtQjvVKM5pX2XsfofAgjaA
wecEQy488McPRriyo92rCzjwO9z5HaF/7ryI38AEcqcTFXHSUnvpwPRh6gxfzlHH
O5qPHIZqH34da427FjGYiXiY3+VwaLbtlQuLxfncHWggNNbws6YlDH7l5nJibmUw
dFaZnyZ6xQaWK5u32Bk7URvdBTaSEstUP50lyffsdP5rxeLy1NWMr415CAi4NH6X
B7eBiC95Mmxa+Kqivt1F9+SoeeVEm4AEKvIbHdT75g+dpSMaFQolStMk84dqfmAI
6BmCDVp3P+W7QZ6kEMTk1XzbUzno2K+m8yHsSQLAh1CnrJ/p6oMSj6iS/uHhLZcm
y2y6+QjYRMAtXZ6Hs7GQ3EvMxT/qgAEZVyR4F3vbuQnBwTtm7mDG934TBUU8mNgh
OjmrKVLOyc9/agbqwGWzIgkTyooJqQlPNzEBvjYO2NCkuG64GmbscoeO9Rnz+cPd
V9OY5aylla8RK0DlIyLX3lS1PjpkbMzK9gpYJlgDW5aNn0waBCYHtGO2w+IJ8Lsy
UjL8YV8CuWvz9Ra1wDp7o1OM1HcPntAmJmi0AlOzGtvPkplTxnrHQZiLikoamtnS
C08A+L6pBC74257BFmiiT32n5QNoST+EfjO4h3VXmjcy/urc62xnmxO2CLN534U7
HDoDb7+vF0Txo975KUJiiufeaBku4bwWbUnqavcalJ8yT+vqiMyI2HnRWJAIsjai
nCEOfWcghwKB5Wh6i7sylDl655qjZMSU7QBMCB6UllrNeR5BCHXgcl5PMY8CjPXT
KjW1sBkFnH65KQDnTj4CkeAES0zy9h8/0iFaFEohdK3EvIoRoGRrfmwxzldjD0n5
3K3nxcVHnDlHzfwqx9JnWo+aQ8X34d0cvdZzEEe2zNwNCuFRfcA5NfTaSB9gUl1s
7zmckUvz7E2U8Qe4vrusmv8HcMyRyHJyK3ZrafFsjIHtErTy/KKKQkviRqpr9Qia
TZEYII8fiitPfURjNrLSEWOYzwzhadyqerTJhQgjhw3Bhdit7xTxqzgfkrIZ/TjH
tnNxNNwY4Y0lAGEdvM3EY+tequCqHu+BgTMtgENQrLxpHv3ayRhb4PJO6vZEewGC
PzEhKHkjFFBPo7SOi4ho+o82XlFuC5gk2jih/ucw2PJ83Yg6OSDPTtX2yngwNnNa
ZxSRehhGhGVAuEsZMbBjP0pIZZ1ohpjitxfv+7mNKyUCJ12T9MbuzGtnIndYDMUF
73b870IvKkDT+TB8mmAcYphmiF3/c0hhT7LGgdNClukHRvkpOOt5pKGoPs3XzvUs
lN+Ha87fXB01dqeDgkx0vrLqy9N6zy8pwbLpz9qZ9KKTc1qKUo8+MK79DR3wMqQ7
YOL0GBLtHCb7PsDIuqgpbRS0jPtdB8q9lEWkxjHSof1cPBFH+M+gjECc5hm+jQXe
2wbjg1zlxjKWkvYcOaX/j8m7Qz5r0qH3i+iKMyEuf3xdDKHOY2YzAWsFnk5Ts7Dh
zBT1JfEltQBwy/jvBU+Z0n6tZHc1B39w266kIfi/zKoDc9czFiDbasIBZ5nKJVQL
8gkGaweF2pOAr3g2onLBBVLGjuvPVOzOnJUdFkglomnzHYDANOZSuGdhF2HTsITO
XUpfTz0AwB0hUSuInXG2mMUbO6aMgG+Vs54qCOwRtkiGGRwwxoeZ42ZND4Do0z0e
WALb9NF1pyokmKXcJAkPbY7fPDoaEqktkeBzpg2dqCSchDj3+gY2Ywe5Exs88/Zm
Soj8Xw6l3snbHKaMXx4tX2Vsjn0luKfLMdhWjy1qd5efOBA22Xn1SR00NYVDQL9j
fN2iP7uswgHewfWjyKpzWeU0iCEjqXVxksnbrfdf4Mx8WEDjQt+oKqxIbs/T9w+4
l3emvZbPA3opcTuqpnEGJ/T8Wx88t+IU1Nvg2v7crA4jMNOTY4TlbOVCBGlQ7Iew
mCkms1Sdc3XRv48d2QgUkzpm7FKsdUwFZvdWgGJDyaXk518jQp5uitjkQoZyExcN
TinDU2PrXyJRGZ0GRJlAp49mqlsnhRt6lLqDxmDfdsMQ3ajhD4pRv7CvZ4vAQBnW
U+4X+iuh4ElLes8qE8lllUMPNqxj4ltwJdV0yAMx62ANrHU0QqMvlo+Gls60SgOR
bYDWa4aoqrsLqeJzKMrVr0Yr2EMeYk4f0KO1Dec5eg+YT0nFZhhj3IVeeqChsTGW
7OeQriz/vnIZYAB7VzuJMw4q+FPSEHe4rtK69/5ztWvigK4KAd6QHgcbLLh9OmtP
4xUXPwbaYL6bU3wfekwBOoo29qZVLAFdiPU6rxEyojBWADEXA1C1P23MnnT5QH0y
2xcl7vOOAsxcRHPHPnJCLoxWl/8/KKaDG09ZOPuvhRy7hg5hTlgsg2qr4VsZp03p
Mj+n/8woh8lYpyLACV2w3R6bvquJb9BeeD8dRFpEHrfn9t6+8k6PfhZRjnrkgIEC
OaoPcuf702iqRE6ObOyKverJSYdNVMfatodPSbDGIdUbk4tEaCkgN1ccMNfN77gn
J333R9ky43QngHOVFguKdSnmbRyqbsvxe+OGe0WYHRkUy55IjqD5vz6PJfNg9HBV
tg2YBWCAv1xcqAVAvLXRQbp405H3+pQtK5wOiewQ+MzpclLl7zeP8y8CtXas0a9K
/YDEZMJB7GuJvEjgFAGkFxbmriGRUH8qpvY10sf+vHIFDt1lbdqXa1ZICw53tPBr
HggD+O+aKshL2TNFkr6ebskO0sX4XKod13PVRfopVkstxi8HxBgk06b4mUTSGu7z
fI7TcyiXhG1E996eApIrcLSUYynmudyhJerl9420L0Td8lecgjTaw29lj4NGuxAX
3+37aQyCjot/24yVLczWQHnX1IukHecGjQ0xjA88ZaaiIs1Gj2u+myJ22yceOedV
UovQN6KeNW7UMeOoBk5DTv3oq61D6/LQXlZN35PoQJaeSlXgLUPDN4ZmQq3o5Dg+
bRLJWoHlq93Y4v9MKq3pWM6HS8oEO7Rzy3PukaqUIZX5k8ez1gGRTrIA6sc+/xMf
0ptmIWmfeq1NE07Lm4ZwRcKlJKzOw2NaNLNk7tG/mHy7ikETMWeHHE5+kUupDXy9
wROktntLdsjDv+uV/FXoN17G3v9EOsFzGT91FklbWrvUZBKNy9qrwEPb23abHAWg
bjMFc6mG+lO33BaqjFDjVi3Lq2crYFC2dfgOCM2/dBSgc22leBkMn4BWqfbbrpfP
a/36HUXiqqc70OlzqdvlDxP15GG9p0Aayhm/fW4T6CCwZ/TeH92naxAW0xMXZsqu
ZWujxxxJQh/8XTcr3WcRXGPfTwFLkN659cFdFdg74m3D6hcZi8Jp+fYl402W75xB
mTiyx+YbA1N2BILALhP7s7OJq3f6Bo63Vpk9JjPS1ChAfl3AVHcRkquR15FixjWP
mHrjPeSlBDbSwxkKuWwBmXagXN0/Ec4+qpNMuWWct7HzkHR39DnIUnzjWpLtpTdZ
jN/0rJ2kFZLfGG+4k35R6Aixo3QO8c70HTuAhJ/y5Xc7iiYtqT/0T6bi5vT6PoXF
Q8nJMMXW7tS/EYiXB5TYWMGHvQWtKrEezT/U/i3nNRX3D6sXW/5VLoUuIJNfkDtO
IOH8P54T/t6WTMDVPE2ql7yYn/2FA5l4L4CWY5KErEbLDn7aR/Otyz9DK0KUKbGn
m8PnBukRjdeU0AefN/yug8Agk7TaR6qxN3bNv8Em5N9+zu8gnt2WgxBc3640O44o
7kpndik3aViIDqALSOzRfhcZHntmm3OL57Lg/4S9UGsyvtcEBoR4XShv8udlrZel
cpNCvbFls9bAw+xcAmct/e6PaiJ2DbyUfFx3dIByRz3q7PZHz5HVLzQz3OP2Pd6k
5l53LIgI+c+8nZ8Ukj14MUxpA/YKEMF3Yp349zbBDzbXXfrsr1Ov/j2rSnKqQeu1
rjsd9PjZz5vCMJl8IYh/Tu/W0i4npbiCyl8qKh52EDf/PkZuz4j6dXV036QY0mWc
geiw8BqozMeTt6of7afT0MULezd5SJTGAt0Gw3UZJCDWLbwcsNJq2fvLK9gmyS1/
uqZtivMg/Vs4AWhH097+bloVG2fbRIDpSB/621d4tOZUmdOybKOcQjGUnolV3+1N
ezvWuwY3vZckEx/rpdl8MnR5zWiQXmyeExMNBSglqyKvcTCByiQpvKLvCYQbNtlu
K7GFPlPT6GJfSzgyr6y30hVXoO3JtKMXtws8R3uCEFindeDqtVVwtYN2jUtHCG6L
CkBHf2QCMAUb1Rz//UfZopctwPvc6++T0719xY6+vNW4R2+HTKtMKstTUoLu/0pU
7xqGm7bndkmEZzjZwsVeQ8VutwhXxvC9OcZPJ+snLZNCma2e6dr8AmDHeBGlnfFO
ZaP1qTJJXttbejlrT+BqbjExthNUTTn8+dSH9JRMZv5z4yVir9sSRmGOZUJelq+/
ndGr7WTPZfTs3lN1KUm6ooY2U6cLo0IFmaMwKsXodaIKCFwD6Zots7nU/KhnNa0e
aY9zRylh5tm5j1yUBdIu430pAlJqZ6i5Eynrxnb5og+XkjtQJLGm/mNm6DWA2PRi
7ndhMOa6i+Z3CMQvHphm8TqpuoEH2QkvB5XuUkXDMXS/fd4W1EuYjvNchXmMEvwu
dTNB8FKNFEq0oQ+qBSIsnG47unq31WCgJleFFEAMP9i+16+ECIsp28kgwdBkAMjl
OkeOodlIONb6S1OorgguhDGOLeh04Z9PGzPfL5pui5lBkuT+udsUdMPyuy0AWWkf
NNEVMQf41yw91iIccNCuwRQtPJqGG1a/omIVwYt3jNgNzsD4ZA83G4OJ7+C7haMd
wOhiU1vJiEj+j/6TpR169ss4uNZ36+lrDqv/WBliLZ9ECq3m1CE6dtnfCJQiewYl
yNVqzCRn6DbKP8OxVeJ/Bj0bcDr63/TG1Xvea7MPtZmpJTanI/p7g+NoVEX8FpJS
JX5O/KMEF4x9zz7vsx9x9wJlAzeVuYKGObtMu9gL6/QK7jX+cOV28Fer69329TaZ
f79/pCV0rTgkPeSQegi6QWkXHdSKaZUkS4b/4FrtIW+T3QdxVIaacYswGAr1aRr6
xL3ejKdxFBk9RSjSmmh0pIcz14qwRCyxA3wuEixRSxqZPLWUlBblPJ9A3RnnkuWq
3yUMLE7YStsz/14jdIGAM4wzPXzHd/1xdmAMEE14xpg9zFsZZ4QS9VqcBcgGtgnX
eIWJsc5h4G/VYMriXY2fC/YpEO5nyRk9E5DYu/poc0EY/3yJeO8lFt5FBE+iILto
pJEqYMqIvCncGs1snYHas/hJp3YRN5EEd6ljx6X6JuScbL13bGB4GPSiQ6HbnmDb
XfEtDV3EwLI9AreTUGXH1dS/GMixWP8cFQI0ajLDWnfUFiOr0PwAmBvn+8dc/DEE
V1i0+53+kKtQ0obLrDykrulruV4qfiW9YFbMO8KBAcIHKO+77XPDlpV9BE92jGXk
JvBE+nZzMoJW9yus4Cb7u+5kLW4dC9ZmcP/QWSDqkyEteJNp8TPCV47Z8/Ett7oH
PWVmHAWnk+VJKTHj/G8Timx1xFRl0AvWQOM+GpLJsOp8yn8poiNQC+gJMkQzjzK4
oVxm800o1MLO9wRSBcoOVZCM4V0+q7fuy6sDKwun0EL7c8RIooA8yO5LwssriR3L
7et3hqSsSfJWggMLmR+pHzBB7SpDjv/hvISqyNP1zF5e68rlMyViAc0zRLq4FF/T
vFeeKX0mRhYwCEbY+tstSyKdAKDqm6DC90EeLYB3jVGJL6bcS/MhYcmQQ5CgqOl6
ScYsHIq9/4r+U+QlZXd+XSy0oeTGabfXLSHHa6RKRWSRvtgeimL0LJPTzGh5CHpH
GgMJTBFpfVy1XPdIj/fFnWLuhHdzhNCwIv4/2D/4Tr1RSbgmm+DsFM3aKtP2z+D4
w+4KRNDl6VEPAoFnJbR8/fHKaTdi3rDuWEBQyjyJTJwmttdbGrOZXqJIvwdu2mUL
fPXLaRSpZwt6bAnKXmGdqVCkL9H8lNVME0mqwZxpiMnipk5qeiddF4Y8S7jjIcA7
WN4ummkovryn4PeiWY3e58vKJx+XQsaBronf4BkkYp9CZnrUZLdDnZaXBci8/9KH
6J8+jQCq3I1UazQKYBqrnkWIHPjl018Wy6NB0UzKl9Pqv/8dm/aGUFckD+Lx3bfd
WY1aacrkORL3fv2MXtf/TWjUyn9f3RYin5MyGvT1NsaXG1lUVRyp4aIsQ78QpnZg
innyeDMuII92GZDHa6+KETtRrSAUTyBaKkkaEKFHF4+TzzivwiRKKBJYI/m2fG4x
7aUQhHQOHH219u0dkXpOLEZlfzdreixWl8jGRqgHFIOeOoclqoiU7wcuKNz0bgPS
guJS9koGvaxPiY6S/ML78OQjsTnrqeZlPSitsNmJtuvg6PTiyUIL5fCfaXBC/AHm
GLrBsWAFVT5szHXoJehkx8NjCuwNKtT4t67f6I/ddWiWsaAr7M6JOFStHJOcRJLC
4IE+T9ttzLeAhO308cf8CRY3f607+XmlRswYoazc5bhP8TpSx/DFbnXznokTb0mp
Wv8ViNbdzh2Ef96tReeXS3gie/o7KHDpNwDdLQaqOv5SwO0h1EyDGDo2pNm5iWVK
z55g/slH+lZQjFeNfq5ZuPVaQhxyrP9z7hEWTMdmJhilxb+ah11t+jJI9gPXpWnl
3aZg5LXAyWwahlebmGK7sJbBlDFSVqdJ24OerxzCGfzB0RtQq9P+TlTbOJL3IYwY
kmRyCAlz/bEUYWuNVBipOKT3AK66L8u3qzQ12LZOsJlzyECgENASl2niDEEbQlbC
XaVhb/nrCv4e96e6FTN9Pe4qstkL+HyNK5kmKWDEcq6vNzGKFyPVy/CJz/oIALBn
47R3jXRx1VqkuejCTIstVkaq5q8e8rL/CnPyvFPxJFUSeTebXdniGi8ebU4yA9Bt
nWM1x+/SLQWa/iYyOewaLE6NT6wMm8gAhHej4f+kILFHh0REd2q8UrS4p4RzPdSO
4LsbNKIPzkzxNVdb7YvbHUvblGM/KbaDJ/Mqv+Ly4stS5iTdZVMwPl8DEW9VAvt4
SGJHp+XUQSkoe0G8k8IGTCW/0pLVX3goRrFoX4DcIMCuZX904X5M5UobRjxsdTcx
LgYyS552PVTUa0/5Sl6NxEpk+KMThoBeSQT3WWDsLlmAHKBW0zHaT1hZNPGwdqUU
CUvG31zxLFgKOatPTp0xBBu4iKsnQBkSN5qLdDsr4lKpjj+iVPdPxkA/BcRV5J3a
ZFBKdOScpnZNMNsvsYXuxGDvlsvsdhFDdRDnKkZzjLDcJrkj14AwlzU4RB8q5MJx
ryizlVgL5ErzF1y1itZsSV30asB3Ai81Qq35BbpZtpE3v/0yWdsKg69Q+fLJMARP
Fj9n8fZCmypemy5RIKVe3vrA1+ShOY5KYA1iloTyxWIgL7hqz55aPP7Hu8kRZu/n
XTc+8kswu0yUu5Z/gaGKeCMt3Z2T634z4UkdYNqSlMF6k9kFPZt/8JDKn86lrsjW
kgx3XIAoRVGvqFr7W0x1EGtc0AEQgJYGPV5+Q9oAiTfr4Z025B5gZRfDnVHTCYA1
6B0lLbG5w3Bq6bcNF06l8dObWJ9Jp5X08SsG9g4Y3NP0zHAPGg0SvxKrSKMjkGzD
uAwnA0oKi7nDp3oy0RX05II8T2MsAMAQ6CbA8yy9/LdGEqpLJ9Uzj0gtCxz0XDwK
5R9Z+ey+Fv2RzocxRu2KG/XGZS/JI9H8aJWy0bHf7oNNYQOYRl1MaC9jJZQwI1Wy
MClTJ6VVICRmCfym54chEBp5RfvSGkZe1Cwa7aOlEaiu/N0MlE58htHUW81io6lK
dH7IgoYVGsxf9RhZM5tit2vSG8X3y2jgYDxt/3ZtQ1ztIRwIpYIyLVcKktyJK8u4
HK4xge9p2UCwjIJY07XOyY4w4w7vIrwCaORZ+nzjW5OB1Sbo1yMb0uUHdru/hzES
7Wn/NNleIjw+ddPR+FeygSM+2b++LG+ripn2fCKEZdOMRqFf9z49+1Ibn7BDbAZR
gaHY1wlplW6ds3eLJ56KL6ZKvLsd2Pu8IBo6/+am27riQ03EE5EtQPcshCztbvsr
86lnh76TEWXyzDC2FxrkSC8/Xu+m5Ha8tYBcImhvtu2QuOOqru64Vm5xYR1sgHPm
joewpBRXu7Yljso482JEtX/BGaMPPyKwFF6DGYX5erdTknkb97pV8B2Ox3R76c/3
ixVep8dcC6xK+UX9amaNfYPKQtkiNBtSIex8b41X7vT35FpfmYi0GNcJqUYSVSuW
+8p4jHFARoqtmLuTYLTWfIFXKyj3rPxbpBw9cWWa8V2488yVgLGEl3pCJKWpjdHJ
h7yS3zKtnNBFVzMHJ6pXdCv5052a6mczPSJYtLGlcm+SCjffLFJYDQ4H6f8tDtsh
P56oFuEw95O6NmscQmjQZuJQ25ufXhPWP7qUuKu4L8jKXaB+fAy1SQhuSeA83mNt
hoPuocqVfAjUSoQKvcO39st+IdYYPRGU1ZAon+xsO7a9QBxxYx4ZDklMNZedZSlc
jPJGegj0Pe0Gak0Rh0Fb9N6yqntvZW4V98CQIkgxA1BJGhKOCRBMhjINELPhwWNZ
EG6TEzhBpfRrIF6FwMeeARs6ZjqoaxKijRyWI1OdXapHEjFco20sZsV0E4Pe55dO
/Ei/5Gjxx14dllAWoSFoFNkQ8369I8tqOQ+989D4DoxKTswcaHHObUIkY1sXc+mR
h8/kuEZJam/cwfFTKi3tw9/CtHEHpMRft/RvbnICcTJgnClL5eTqSNDFBkHGCN02
1vt+7BTPZxy5tk6cxfVfVicBjFE5Lf+21xzbmD3oPLiCCJN0a9FdEpFWRjUgMukc
d2nfKLAI2EAmxm6qtCqUQUSsu1HIyscAcSwDX4IL1A8thO9qrSe1nMbeC3BtP0qy
vr/tqe655X6B2A74A0D6KIta9T2h8lWw8/yrQ8jja1psp6qiDyWzkg93pUXzPesp
Td+7xyGAaEROaRSK7tP8LGRkw/FKmphZu+ySsyT86gZrwWIRW7MOtrF9NlZsLpB6
EsgRP+3ZmBAFDdKSzS+GJX4CuwlsMaZHa2s/B0x5IWgAiQey8ScaMcClBeNryNAW
DoIPToV20pvGs3OyfN2B59Da8CQHGHzFBWnp7Jcve57mpH8wl8ZoOVHlLaU+KlWE
XMG/kjQlutRpeYKst4FuBQ8mT+1O3mohGLlBsSwQGgKqvuNbZOggKIfduN9GebYm
+M3SK2cjmNL3sAIhpOeP5YF8SvAxTahXGzSr1Cswmjdnrvhq2WORp5yl5hJFtKRB
x8oRwgSt24CmJVvVARXjwohiI/PTlhQmNP4cZFTV9lNFmyFiI1HPTcryOpQOFKgI
FtAeX6Dxgt1FNDBwRP9WOp81wcE7bkkfj3vXNWcUyLUH8K04Z+WKDL2OpCbGMlWU
6RNet1EThmzZzmUzPyjyGjbAM1Jc4yXpw4S888YVwCIWT88lQUsVUWARMFmuIVVv
8HpqVUnJMcvT9yS/VfdYygCFTwT828lOB5peP001Jf+bZn4ABJbQVBBnB56hjKeC
l/ccbRPsUpoyEej697uf3IW0eLnXgdRDTdKaxNNSiQWzJzeNeJiaSd3eSRK/Fpcq
lTh7IMtzTOcCLVheQzuaKseZ0P7S6ipcASlVU9XRuIGkysiCgB8NE1F483aDOcbL
H0ADxmuC5XT34v2xpIPiOOU2r9Za7yJLwEWwklvfxV/DtksfwFFU7zwmQEUB2QBb
OlQ6NFrFt1Bip4FkPUHA3XrGQxJwYXD+IfLd6btz0i6T2m+85pOVm3cSJ2X6RWcd
kvC25uSCB8E3XJIjWYHWavPlkg5uCDDSmCL3jHxqlUsK6al2tery/w9bVpgp4m2T
wN+aQbOQGbrxR6w2RQTeVv32zGzan0wqt4U7NAF8/DwA3JnuQWTbQyjbCOyC57Wk
pugWGqZwDrMN8aJ5AQFpCRHw1KnNBIxvLfJhGIR08ejXinnCTgJqX8N2tMeV02ty
Fqg+Nf03KkM+vWhrUFOEnvfyE6j/lhfKL3B+V/ubDuPPQ7XioxvpqMRYaj+HVdY8
WHYo8BnMyHgR8qHQlkTqWWwL019iscoqX2veiJU6knNnvYc5MuPQ/36XDJ6YnNkX
yItvqKutWyJuRpw8O14FbCUtqMjCpL6Mf+feRvbJCmvWF7ksAp28KOxFo9rpqjXN
X7SaRTZkrh5ToPTLmaC8DJ+zzWsMobN8cWqm9Q3dvCpiefv1/JhIBff+e5j5Z1Sg
FsBLErAl0rs3g6mK0Y2hL8B4k1p6cqxsJuzO9eJOctuoV/ffrO8lyw4KfQr5WfrN
KcPAFy3gaQjYskt6k/yGdi94ocedFDz8Ei5QYPgEazgsXxStf666TLSdJqb6R8w/
PFrMSacRJZiYjFeVvlfgM880mM3MUZs9/SYEWnM3DXCXuoOdFKc14RDVGnwGqPYH
Gyf1QhzB3xhPr4trb4DqQucCyMuTR7W6xKRyOFSYJ1OYuqjEeoU1wdPbPWQXKEBn
LipVbjDAUs7oDbK2usn+j0guQvegz5ihI9W0JnTG9bh4Q3TJmdrxe1ABkGEpeKru
2MdKx7utu30qcxGaJZMNFuaUNlNdALduGntJkR4Zf3apwwrd6YM2N2pcZVPyiITF
t0GE9wydIsEtN/lk2X7WR6RfaZIyguRd7/1KI6CHE2yAZztQ36AfaMsxJXooRM0e
laohMrBQe2iy2i1EiTlSUUgAfocq9V2t23BYuNO/muQX5TWCcMdxCdS7ccudY1Uv
E4dTmg7LIBnnOgDeu2mFcGT9H0jQ3+vWVA3CF2qFKXPf7pJqTaJCki3EqNbKIn77
hcEYY3i8IVtDRZ9FtxURBx97ycqsdAT8aQUgWxyZPw1d3i7svbxrMIWEED7Ssgug
qBDCZfS2RZqQQmNzZmnA3PdoX+AlYFNH+twg434r2MGcTIw65nQigEfHPE/rzvkj
KkYOZif5MRW2IJTDmzWvvWkfM4qPr9S1B3ePpwit786F+3WegKMWEWmh//7vBj8Z
6Nqag397BXUuZFFUMs948hCmzBnSe5GwWV1GlhBaIZxQOT7mT7AqXv4GbTQuUanJ
rGoxre8DgOEF+qkm7jWPLYFu9NUvI3JyFHJ/ceHKr4tntYkhraoEbItI6eM23pc2
nKaBILKHQNQGzOXbYWVFQfY9Xacmi7JimfUBHT+xKllI14q8W3qoVqUittDuWrp/
sKjurE20/W0CzhdRA8NWVPMVyJZLNTOiJoL7cT6h39wcsvEtSElQM/rwIqhK+R6E
vHrp7E0o/mwIGluT0o/eg/v4YwNS3qzXKLfWrLZy60bFmrqUSLanMFgk1hVP5xXM
jFfBMprXnYshNhqDfKCEloa63Cf0W0SYiNlWtu3N3xmQATfZoOy5+7ftwqIKDjnq
VU3Fcb7vQLE0R3LuyPYOju99tboismCZJvaqnJPS5TS7A9aZ3gYWXvPY/1XXoWiX
853+cmfTBdiRXR0DDxdOZws0h6z4cUvJjpdEJYcx96MLagmDVsK2kGHAQqE5wN3x
pC0cPF+4bsa0qsDi7/bzP5r3ZfzXOCkX5V2wPFPGFp3R8aBs/aHX87s2lPYOPtti
xz2VUDXnLLMSHvdtyJSxNdb9juOIdNw8xTNDwEUKnaeUZsbpdPTTrCwviSIzrOIb
3tDo6/3MsgWydO4xwbmyyeibydQum3ujoTHOlZ6O8jdWiYy3Pra/LRO+xnlDtjMw
mYwg2e0Z+f1nrqZMnP3m4HS6xjw1EKO1f5pO5nMz4zanwytTFd3j5dC4Vil1zGv+
0jqSSM15P0TxmDmp9EQa2siluTaMeTlvsRW7/uvFha4ypOQgZY1qERF79QnbH3e2
Ih+DbKh2OnwxM3nEA7DVD4QRsvRosHaGuMVsIkLmaTYU74H3h/tcG/9TVSDamj+o
zzaa+u6BNthyH9qQoP9F5c5XH1YOyAwru5qzVxyRMsVFNlKPeL0pMSiR90SM3YpO
YFV8Fah//L7n71+7VNKiRaVKGI5bNAntZ11vR2B8DyJxq5vy2ZMbDeIn1aSK92Y9
XNWJhvJq6sFg6QpwcQquVBPojYf7pIYqiJt9FKzhObb/1wRYkj2d9l+GxaZj/vLH
n4kzDt1KcJLEmg9JGiQarBDB4pa6yZteK1Lg9a8Up280qJwssI7MYKkJ0cmubLAG
C5b+8jA9GLAIwAzOl6n1IKvoF5CV6mVc1F8ZS6PncQ2eviczpi2SMdUpVkN7aH2I
XZ1eSu73DppF1bBpDm4MJswNKTRnLKHWgghr3JJpZFfBrsfm0nNObMtts5RhcpgZ
c/bXrUgSYMT666PZELOZ4fuqeeeVWgQIzbXqL/dr0YvnhytIBvYl5jSc0hQaMabb
vG4i5noVgSOIottK7zWxzTZXDKSSgKYaYrabT9CNO4xcs/S1IcY16jcQYH9WV7EK
JsZb7vwj7zHycBQNnGMTN/KglOTCneM/wj4IcgIbkX/euRk+FxHrMJEAtGmCD3Lv
10zfaaordw+GZ2qGA2c81k5zQKgHCu6hgJjlJup1qwn6Ff01kQAtBUApqi3HHl55
U0iejBxSUI2kEQNnxBXmwfNRny0mrBjN/Civlz/gvmeTS3sbsLKjEB9VAljN8M7N
2HjT2RqrSi7HPsYbOOv8w7MyGo1Q+NuDz0FdyqTiOqPS9R5y6LZ6RIsYroR/1hsv
WArvwdxeICdqrP71jTry2VxBxTOMDKHzZGYfU90ZkgVh5qCOus1QwwQida4fuM8t
NvqFP6SpPanE3uwPKsXVT3eRN19sndLPT6Wi1Gclt4L9EJq06PJvXesp9MuNCUlE
HTNlUKyTT8nMCNiZ1VXC8ZLGfPKLUecwqKLT0RTvCwEbrGeLnkDh19Q4iSiAh1hy
USpCl2wOwmZczb9AtAVVo3OXs2XDpuMcC7ZQYxi2Wa3DNFDLjSMasPHc0gdDbaJJ
3JCPD27mSD6SRaHQFwjX6v9k4WmStNqioHMvHQ/b6dplgtKHYZYHuKDmLt1qbXO2
SGiJy5pEtaeJtRmDdu6r27HNC1L7EdXhCaUNxnxkcGowXTgfuQ5n1zgBOhIlCr0i
xbESfdFIrzEnUPUuq1O8DZWymiPBtL4R4xsRwqgfcaTtOcshk7xwlj7wfLy9DTWD
NZWn87n4eYLyhGTMjLHILJWrNIoTg7ymQY2+JgcmcyAlp6Jt+z/a/Z1yHkzwUuXi
qa4dh44dec9JvGCmzA+B8ShsWIugN9OpR+OJbSINbGOMIi4sND0cgCq7bA1O9TSJ
84Rb2+Qj1d0DFAeq9grB7wt3dDAtoqtere/n1zPWlJ2a50kqLO8dpXQVwgCSJ0m2
S3DTFfc5vwhE/ECO89h9S2fBgnFJ4M7pza0CK7/NsQLAVEZh2M87zd/lGymby3Dq
kaJ4dfnPl9QVinSwHpRRNg6JT7qJyXvx4LyCYcyTEWkREtgatSS3O/NvfkGjFBtR
tmbgJ8oxX4vGS1fRD0yZkcSRynb0QeamPqVPrCmzifvNuaWVjE+8CAFx0YnkGuuA
nRrKxmAmY255oij6+XCVqbXjLWw0EUkNKOqnUb3Klh2JTV6NAkoQHrxzzRKq9Spk
NMjaEjbEOg11q3Rd1hsn6WCdMo2u2xjEgDoy42wZtqivWbzYUJYmUEHgRZ41wvMq
BwAcwihHfsahkF5m+DwlDiMLEn6XOXM40PqzT4vBhSwO8Eb3TR1iCUqLHKhoUZa7
Uvm4x85HwhDiWlGEx+kjxL7b036aMkSRWRyt/g1eKw/8UVbzQngNZuUTzAbaJ/7d
UeCRrw/9lb8j17oqz5Kyjtegc4UDjWrMeI717C9l9p17t1TNQb2d11CDaHz7Q+9o
VTWG1//PT85QzVDL7QP1orHuJaXR1yvw+T3fVqzo4VaWauTSb4Ff8TU2Vj4NRDaZ
Ub/1P7vMxoQtZNYBTlHc7BXReyPifkANFJKn6V3eEYXQNFCvO5YaJvc58tn1q4Yw
FgVStKNLO4NAfJjf9X+hDSeZC78Xid5zoGZ3JT7wokaP6gFrLQmX7l/TNPAhuyw2
SUAVuJCKMTK+j5hiX+dYIXwFHTGewNeMZppmP3NsD1sFio8MQwMgb1KXuaPijnq9
7+TtDDxCOLjvIbIJceQXLgAW6lp4N23AqmelaZMbGlAQK2+LU6gKrFObmZBrYDWA
9O3sp1ak4r/3Tk/eRWVd4jOgHLMA3wJ9e+CXn1GcL08yEGFdZH8li7r8Z0Hghh81
RFl/j7v9q3k65yTrig1IkS94TjOFsBcI89B0CwCSaZHOOiJi9nwRpwL188x0di30
s4aD958XgCaCNAhZf5nRL5SB/W9L50v9OPT+5BFXWFlNleX35Doe16MXIsx5NB6X
h+83ULIokQa5VMuwO9Xg8Prkz4CD1YKpbuRdw0PZqQXBFEQmQ93/eXa4BVylVK5g
tEFr8YIvnMN3YKQVVyv6YPJLZASMU8rA7zZPJW4VSlESTtsiNTdQkIHcd09L3vnG
loIZn/8Gs59v98zMcRujXnOBdifsbnhfiHAVsCsyOgRqFyiJ1gGbrRZNYdtVtgBI
HBaGXJAMFsMsIIWnxtNVVhZo4xFmPbRbGIuApv8bMKi52KrOXU/dLnkSLyeIx6Kv
t/i76QvVgMVh1fA/340yYQ1DOD67Od7mEacV/2i6gBo0Bphxl6y0ATVLPNMN1Mei
hfso+N8xeACt8xPWtW8d6HyIFV44sDIcWFgWVJY19hVNe5Y27LQ4Dm3VIfgQDFAd
QPQIeQ+NqxW7sT2Rt4d5ngyvUVYvQP4cbYqDZOEK149UM69ybOmRcWOd9zZPtJgg
GI61vq8lx8CY7yo5xzpjVZzqx0fn9pWV0YUoc9LOlwiMmo4QTZ02DYI9tSgHSXZv
034V/41zoVZ2QwiaD1px0w/JulZSB2gEM6VqiBZ2RE25RVoJQG37zizQG9ts4WPl
R7cSsTVMEbRO9ngXL/rwhExl0QtUS01qlDM6MHENGzCmJwf6ADWyBf2MFemMhDQD
YiiKJsRu0MukFCeCHk1jHVEyQ5e8qILTnVde/DEkMq4y2T1HUO/Wlk4S1HxWZR47
a+qpVoww9LEenOr2CmuE1nzqFQU7/dZYxay29PiynkbzBG/N/b5he4mWtRAygaim
PRzXXsZ4vlrB8120a26RX4t/We6J9z2NxC2LVQy3fYrWppxFtgtNPdvhqEf4tE80
DJiCDEeof5O8Jc0aoyvFIQADf5CAc6SH9pgIM8SeMOHCCpIkR52YCpKHO8EVU7G7
F31bRYwhFr4SekT/bdMR7NGtRz2QvzFbzKVpfyn4mcf2lY86qxAOT/tTQRRTTpbk
6liqhoAilPXlD6bNoxYmXcDzif/kWXEeXCkFqiWl52SvW1f90bE8L+ly27G82vaO
fi/ofDoeN1Fp8hSs19+RR3soX/SB/aW6VsbKoMfP1mzbJU8iTqdEMBrpLtjEJAwz
x5Hh9p+IKfSADKolbT5how7TO71Sx7a38co5ME25r8ij4hF2mjpOgN/11OJZ9eoa
VgC0aWtXfk3BhwK+h7BxIMW7q1LIt2Me1sVr+O9BYSu0xroV8Ge+QGAYBq38BmMu
wMWpk2S1tvfKoy5XvvzwIHxl8o1pDyPMPWsVIiPsfypnhlHKNLWbak1f6qZ07mnF
QWNuk9uq9BzEQEwDNHnvyAUEAvfU4pgysSS83FuK+kvYJ54QeVxZAdHv3SL5Ek0h
HIIGl4w+UK23rt8QMxVm8dwwhems4tRJhLdEbOIAAz04OyFE5M2ArbhP1dn7F4K7
WEup5l8sYpW3XDjJPQcbInbCFGVC/3czFPnnhBHEHcMAZzDJwcuwahmlBAKd9o3Z
Gu8NwY7AsYrgPyo6dz0MY+Ea9L7HkzHfwS1I0lq36uZXj3M0aPZpFBr9dQcpzDnY
h9T300y7lcwQP/GFdGwv/fx+ESMDXg55wkRz5ZSVkn46AxrS6QBc55TeApLD2JNc
0nubqCd+aOlHkfiieE9EFJ+rZCmFLe2dhfjL6A+4JO+nUaq+GEgIkonllNr8fzUN
3u2362d7v+6HUESI84M5CyDn7Bo21TAsAEyveKk+qrwemhdDxtn6UjuVwZhmjNdK
Yxrv3FGTFdL6+71J+aATa5dm78bdUXANPqOb0emaAzjARglhMSp8KvGVpFs1/QNp
SVvdg7e6kDlAwSmHF/VePbde1AhZa/YUaWFxjFGRlyBTSyrrDISD2iOrMlDNdxBh
mT++yDNN6tAh+FtkdVOVfuPLPhVlmB09CtA2JS9yfr2+lZ22j9nwt5VmnarEpsyN
zuH/dyqt9JuoK9+2YqvJZN53evqUf0nwlvmse3vDaaiQuW5Y2Z6C9Tb6UITddUrZ
ID9wmbrXCYB7T4vBjK07rI7aAy8fTL6ONAjj6lRBJuxnL0iAfnUBcfDJhwVtbUQw
PS6PHPx9tBYABod6ei8UUz63NzZ96wLOlSRezXSkFQHr5t8kJhUkdh/BIO7zDzP/
4uX4I20nZvcS8obks0nX2Kj3p/wOLa+aKI0g7WvzthdT7AGxVMO+d2h+B2Cis+RB
13G3Nko8/S23xkm09OoQsCIxZPXb48Q49cCT81/GpEVvXp8GZVrLhrwqHmi0s2Oc
xydxt20+2FfRJxgJcetEbLL+xwCAxxmR/Z/LO+552mVMCF7dKLT4baw6ai2CMFYx
Ffa06bAC5q90N+qsJP8yhdOtvUEuKLNsuAVuf/hXHjutwaC6WQ0Enrq0t+MQpowt
BcT0mxVB6nZWuuT3+PoTYJDmUpzFQ/1u/0GxtzKz/E1d55wYHJ6PLBYvelK7ZvYY
vk1L+a3EKegGwJB5dsFCk/QwcYf+mGCq5xaKM0YutxUu0qV4mahboQpjMd0kXONM
jK509VjBQ1s3IFHOPcr4qbiarvQWBDosmSI6tRf+MNQbZPqMEAXxaWJkJLp8Le82
fDCH6KQ21jiLD2++sREXKNUvBQdzU7QoP2QowItrSCjLpHnZmNrND8kXGBc0DDtt
YWv8MATVzI7AJUAwo0/x0Geq5lY0zqgaOqzFYip48h816gImxtZfWeQcR1Wgtdru
/W0nNRf35C8XS/L1AgCirS614bP/1YAIsnelF85mdZ8DzJmL1QEX7AesMMDLA3MB
wh8SHq6rl4E7CY8RzqvELB/flZ0MXlwM1sYZDrDH4m/e/UYUQV98UumVtMz7vtNU
PTNfbZTDAC9QOihkD/97tn6EXHiVqMPwcRz5l71nh41AgTOnryPYTDRraPwpR7ZJ
NU2UzUrsvjSdiSLnK4dvy6g8zttaLQ1ErLKcp6th2/HuR8r2qFZ6hLJ4ULaOTcQf
wNld2JvGHvLGI+w7m9NxSnAkwnGnIpE0EHqKPL+/JFXnyiAIYPearHYrTMBVoX88
v3axCY9dtrdN6jo2d+gh+enFFi3Y+NwpWGX5vGTGsLrSgr7WCiRSL3CuYlw2MouS
WjkGJgxPJhf879P3UXLji6tVDjlc6rTKVt2MeRd97t6f9l18hNONkz+sBRqmePtf
fU9L7N5greKCYzMpIPoSGcK17VgNI9VSOBK1KwgrxQ2yex9z3BsnCY6es0MVpv43
MwnGhd3K7rltdRgItdA4Qtj3Glt5mgj3RhtM3h4TEUJES0lBobIr6t8JdoCN3/iK
IieSbWI+b8XGCFVIHrq2p49rLCp/cdrT+ZTIh6WSM6CpoRTxj/kROLfIFoqt3fBi
f6X47rXuQAyObzXvh/LCakdVCBm5O8fzWqNGw8p+D+jK3IXGgXL7POhsnuJM9Bwl
wpzrCr+jRuM69VMx5HH1BQJuyfNVmTonhftIvmmzu7tY8DJ/SM/CBKQxyrl2Idjk
ey1WoyQ1URvWKFifMB9f8lVNrxVMv1MSrxbfOpRmP/1fsJeZs7DFJzh/irKe7bbI
EUVqUcF/j2NZGwdM4iGunbGeFAjMnU1xf2pDnxA16d2WT0b3lj3m1v7UEcaFFaHX
rj0L+9nUGmFI1/xi/k8QxoR1f5lh+xnoECASH57M8+lHOb72Pm4S2vj8hog9mR29
oNxM+wZ69Aq+MDeEWD+YYW+ybDzjHd82uKlkzCxsGmfXEEgzRnXD8nE6ydqj/aBx
CQ5UMB14JJ3NtjDU/K1w0vjRYSlcOMIvK3mSXAjRMq2oAQ7NAMBEVvsLNOTCMJ/f
S7SMPBB/fLQoGh/yXLw9RGfJ3PrTH/gCzhUDTShNO1m7fTbxsaczZas5Mz+9sLgR
3BUgcBM+t0pdCBQgrmgXQAaaVfA1TztsnZIXoXucfgbs3CysgvxkXd6P+sq7PGUk
m8jVqVlOhrQ2oWNmZ1JJlu5W4/8p6VePVVMPIQZpx8flbfPsOVSQYs35Mlqz7FAk
NfSh+DhtLtpvdEMbja+3ChfTWXSkcY4BwmAmgJM9tJxvWA6F3LJPIZm3OVdCMgCd
tcHGGWaysgSqxUIMgFHyc/WIb8Pah9pC5FyloSj8hVjiB+WxUAm5dabraSahROfy
qYaWCKB2lYUuF1t1/GiOxTUmGLdxIabMhP9IRJTJDGoXl5qAKLy890eAhGNIoLaO
FfYXIfsMaGD+zrTRjPb7RO2gRu4kw3g5S/tAIT0MU/nTOWknAhRfnuk1ynTvqSlF
HJDFhaxZfIAdA9NkjeZ7fLNS/4j1h5DMKgCwP17TMu+WPZH7tzF32gXaSqJHzbrC
spnTVJIM+4gVZwIuJEIb6xWA+iFEKDqPlQ/4uP0GLfEzx+b/DAOXnUQkBHGe+Roo
1rul0FFbjMylmB+bfkS6Y7msSy9nOMYAZs5wIbUSptKSD38SGo40blLB4NFbQFiF
ogA23wgA/1wvjNe0E6rGO3/6jaTNyYSWFoEO2QoY1foQNp4Pn7Uohn0NuojKbGZI
OI1eT9ANZTLrhnSKZn56IThPxyZsR+MCaBFirvDmR/red44M904a72uFAe8gxVsD
ZeY1rOmmolfn64/XCIHZWpdKXlS0yOZb7i6LtkpmW8jup3RTMiComRVbh1w8q+72
XOa606zMNPavnmZYeg1RSpxzo6bzcN+xsVHzatrVxanYopclfhGdnZ5UPlIAWq7o
Q7eeIC+RlGNgS+Ryl8OzYy1yrax+IhqH65Y4j7mZKzXjcx26CC3iZasKXtVaqF49
5sCNIPY5SeOdGSeokn7oJriPmpqBXc/yUawXiEHac1/ff49Cl3VQRGNM9u1mgyEv
qDfQJGtXtpRPpBq/WO3EG23jCWXTUS/a1SXMOlFbzF8wnVSL4kAMfSTstOZUWuaQ
i/BUBJXfkBEP6YAXRWCxGjnneX2q9w2bGiQYAXvETAXpmgJ6EW0F7mYbUCcDfPtj
c8lyiBeX/IsxOo/jMcVecCjahfi/Q7RoDtjC/mflgXwqlpYQNjB4hHjzPeQnbuHi
m3sdeWM/nerG1PP/26tupTP2ysOnYr6Ib0eWOCn6xXnn6ifKhmm2nh0jo3hHG92O
WoAOsJpN8R/wyqNgemmsxxNXHl2CBBiQ4orhvWQYfUh+GRkCDfNq/2ZUzVYoTidS
Jz34iNthh/QbyyxQtqgwRwwxNXDaBL94Jy4lH/UuY4i7Fw8uk2qg4JIB8sDvHU1i
HZdYCisvMqVXDea1INYAvDlNk8ppyAP7Z/ZcGj/BsQemJskfr75QOVdygdbOnf2E
65ZOUng2t5NI8b7xjkRPIKYmudDOLeLJlaMfdnWE79DU23+aGOcZHB1WVj+Lvs+1
6MAYn8i9YnwGzrUNI4peRJBurrO0Xi1OmJgFuV1+mCgzLMUwirl9CU14LdWFBv4T
e/2UCxlZgzeSCXfInVJxiOdy7o969EE0k1tn6OMi9YTQ64N0JCmOFqUhLoMCG9Co
VfMeEJ8ReU3ITk5msX0L3FkZf2ZF423GHf9Jj7XlchbeTG8/V2oIjPhvK8x5hsxR
aTJMfaH2uW/yvLh5dLrsotlxaF18sCKAqaVp3KAdUJEz9UiVXYDqBiDHdwr7y/O+
BXKRY6k8mzL/0iXgkirkiUx40hfjSt+jRCy/tCL9ugKzQjTgW35m9xd37zfhgoD0
rEk0x3MuyB0/asmMov1TLFNRGRCsr7fB+gCD1aYnIdVch7QU5B7GzAkZKfTctGIC
Rola60K1ic4RZ9Gt15cAYKG0HgYG42F09DvW1UIeBdsPWIj7xQuNRopZp/0zW6M4
n1gVSQgwXzGjEM77/5gzdoC6NWDamlmpssJfkbkipfL24hSnj81i57CetBDgVtdM
ZY2JQXzmPcR+dAdUdaJ7oILLEcGGQJpYRO26XpEKfROpXGKb+Vd2JHjDD0pHWs+N
7KxlFACMF16pTSoG4VWC1JUbxGVFG13k0WOz6jfaBAMT4PK+vsuI+nPWbaOp+wP1
6k0dWnwT11hLJKaixtJn0hlAnebhylkkO78i5LrPKQSy4nyZtdIaUIkuElP5wPhO
ehWyAfPs0xjATMWQHeGOUSna9iK3a6F1WawCGihISHmaezAe6oj7w9hegpn4wNNk
apMqldYljLZXgiAyrbXsOJh/vQqsMNOG/W/wKC7KZeeG47SYzTJ9M5KmIWSq+tsa
wqJjuCXd2WvBLDCJs7v2rgAUa6m5Pf1RMA1iZyS46Sig6KTsmcorfWw6F1pBsb77
G9cj9qckpKf4qBFGngF9Nm/PTlU2APHfKJCVEzOn2+RsWgFxok6oecNqc2/fWD8u
VsVwWfmaAqE0Ju1tMJEzGfep3iO/0y1Fo4CSG1MErqnNv/EmKUQPhx6x4q6iiyc8
G4z9zRaxg7PmNK6pRaPQu5UgU07UbwRfW/Q6ub4hPF1ttlXQuZ5sLAb8HUCSwdf7
oBGVRX/lO+4vSxElbZi4rS3V0rfjIYHtYIH4DFDNfHExsqD6w3cAoKGv+z/swpYh
mBm02jMaHIjAizbljXUK5+IarbsB+RLDk8y6Pbybm0a5Yujbtcgi7hNKCQ4HbTxm
2arbpHMhEYxPgEx1ay/RCxyYCYcZseuFVFRDNasTGc90ECbDBRQAq4VfVOa934A6
rAE/lTOkTD4klr7yx+8D4/xpsIwEruzEbaUwWNvZouZWgx10nKNAEr+j2PZ05VSq
PDODls4vQMqqA1ViV7PGIOq3jJFCCn/8CtEip7S9nX8MEdY1DIgMDJEoFtTcV6Gp
ntBQHWP/sLxYJGdhAO2GeqRIIBhMGSERKj76colvW1MvW5sdhJs9N7rZ/HhVMt8A
0bZAqh/+SpW9KOInwIhUj8CpKNQDG38Jkb0tlLOhj+eVHR44SbiHYQWcUmgah2Sb
Lq6K6Tw5OqFcWJZsuGk8PRmQeRRX4SzIfXNjyjfHgeKMEIdFNL+nNkcCPuesZwZy
DHh0IIQZ4Ek5LWq18pQuwUCrm8TOT1h8zwBuTOgzXeYM2KLIGTLKD1cZmsQbg9b4
Sd54CWAPhZhmInSl6UWHVGvMF0UZb6+YtnNQ84TcBhXncV0BVUlZML9EV/MYeEiP
OGfQcEe4bzvKrmOQ3iXQeqlR1YqRv5OFNU2lJTB7vc1zl2Y1RXMNBd8URNxE45OF
bRFpp/ijEciXUxfoBmuTHntinioRy8ND1NNoPHfzh/ljttZe2AAgxOzWtJMrE0/9
Y/NSgz+tOendlxiLz9A7/RmH34GXEosX34L5VVEG5gNf0mToS2NF94xibE2yUega
lki20ZKH3qOi9O5siiJ0+xAwUlYJYN2lFzpKSL4lT4hsH3uy2qvlob/hpCwnHTLD
4FzxkHyNJvrqfDOv/kxTu4GZwK//Y3iOwnMI6uoj4hAkkaf/QsT2dGBKS7THfLbu
nqQfnCHGYN9i68DDS1MH0eT4+d3gUgDWlWx4klSmwfHV4D1AAK114WQMPzB8dXhN
4rm1GV3QwIOp1m2qZOnyrh3ACaG+HpIb9D2LR57z4D/pmyCgT1tCNV3jNRxzjApd
bvuem5cQvdrZH42U9OPNVaaiFmSjypSOaDnhIbE6V0jPshsRzpB4Jq53C4s47+x4
ObW1Dioigl1giu3AINUA5PRbyKgQLQUlLovC+1KwIFq979IgDdPLpIeLTjs31wiF
QC1P2KyUfFbBX8mdSCzn1AOoiih9gowXSLNMJtQhHHscix2JeRuRIeFm+P5ZrCod
v25IVolJKGDqza23Nwu5ckhT3SN+8RJsiwruXobat9r1K7HTlrWiIzUuC2QDhz/k
1vuQ+0mQYXBTJwkalx2M5VlXdty11+TtR3GJWRcmaLb+n8/uegLtoYJc0e03MuI7
KrMeDYZxBgRy2p6lr29Gmq8hbKv9YhAnguh0ONwniHDi7pqNtA3oBMi5cBLYxrzg
rovwUlCcYYM+yvHBiUe1W5dM2IXl9h86szYgge2SA4fsTTaBTDRFEeh6UXdg5zLe
JrDOu96+J0Tc9885PcWuvrhm9ROPxT5tBWYxYp06VK/8iT9hFMJ99UGf3CoCDsze
pE6GRxyZdtE8nZl8Ny4z0hJpHarsi3CdpTtaguFo3GC49iUtgwh8r5kqeL+gybtd
2JIFDmg7mtGrUoCtWjc2JvWinKITaPjdjLAVRQ77j4AU/v0/4Km8aJhuot/9KS28
5pRQ0MFMxRjH+LwRN3wS4uZXBnwqSG1Ra2Fy47OctL+4G/C2S6PRATer0iBNyc38
TFaHI5he0XaJA/+7Z0t3RC687X0Thy/POpw9OUtClMFyBDtvNjNjY+Z5aUje+Ve3
jE+Mjo2kra5VGan+kw46CxOVTH87JlsHN+smgvnV3UwFzglmFknM+qe/39U0Xr1c
cb2RGmxEHuyVXN+InLFGJyL/ddRxllLcIdcu4/WUmP7+FESYn8apnKA5/FJLiqsT
f95b5YtWaiLLlZSN8W8wPCEcUUM9SV1+eq6wm+lsytMl4RYPb7Ar/bivXkIrXypG
RgDrS+J/aY+AsJ1NVSkUebHQ2nX0iGUrNBEv1n7qEAdh+ZHszQszTfDhA8SaJ8+/
YHpSH0kNvxDkkMEbCcxCE88HXWmgYu1NWZ8+SBhGoeKdE4X7H4TYlldx7XCxCU03
1e7B7u9Lbswq0FuUX6yRMq9BsY6C7+bdYIWpA5ByoCVzoHCSyZdX7YgV2LZLF420
J1P8FSFP20M9lzsGxA9NJg1y0P/nnfI7hUkaPPbT6ux9JCFtRPismFCw9W8ByL2B
4rdHLaAin6raN9MdkS63TBsfW7tg7hlkD03gmHpRpcxkdAtjxsre3SMaXMxyY53U
PwHsHa6rIhjKBO5RqbHJAWiqyofStsQqrdWivtCIT9zU+yd8zU2nKEQ0tQo6Afo0
FC9xn8JJRhXMZp+ri6snq7YR378ewdAgfsYOQjdVj9WbYRi3NHFk6KXxtGlUGq/W
TKoRhutKq0TqB6uy8fv6JFS6F6vdAhzcxpU+rypyv2wgr1jbt0u3rE/suWXb4/m4
ZBnL1qkQ/51Bia2NCrAZy+Y3+Z+Ol3jCe5rt77NmbYYyqTwW9p8KRra3PEw+HVXU
qnbnguDycUQHAz9L6RQXXqfHj+zJP+l4A51uDw5fqC82KTSU/mMnFA7NX+Aibu3V
FelXaoMaNawHI6vvDz9kZOM+2k7A8rGZfX0gQciyFRvzNqbHdhCkY+yBmqRt6Dux
3Xz5GnbsdMH+CpYCBuJNA9L9hohptH4lbfInilUem21/EAWmg6EVOuikVTToda28
yj50iLQLq8niguzRIXNb+E74AqRAPFMUK8Md7q2P7XOTW08F26JAUkXR5GCLsEf0
M4SJa8thXmgdeIy8qKdl+bmVEggqqXpV7JbpCA1UTKiyrXcGdRCMpHleClvtHUjg
K1H3Py71evRYs1pKuqsXcJzevmrAV368EK2dAnilp/01UQWww4B7CC+2edYeImtk
vNSNCRdCoATa3R1g9iGpt7fGdeUhRGeNZqx/CG/X8JD/jTkzs46z6cpdLF603TsV
kpjlz0UTKOWOXD7zsJyeukeaTEmjLYkU7Xgx5qsQElA3gUgf+POPx4/927G2Xt89
040vB4+IhwyuQIuu8MsxvNQxFG/nLUQxZu+kEKCYwZw6MAOzDfqNIMTGS9uYcFc9
pD5OY58iUpcx++bUpZhM5bDRlDoHelPD4MvRhypYTK6BeYjNouZKqQcAn1bSiyl8
s2K39dZS25zMrepDXapaEeTKHQh3B101D38oYHS/O+LDdiQQz5tRouVKFhleW65t
BoIxs06sOzVSpX85s/HYHoo6aIFix/xFDvXJdlPhwaXRvKnNcsMTBPx8iTzxQRHF
8nS9X0l9QXXLQ8soaAiB0rdvnbl32XcRQWtyAPY/tX95ijmbBp7JDF7poxS9RNNG
3pYM/xZtboIHhYZ3sLto4/x5vjg0xuqWi/06Z77wziVjPBiDjqg3ceFgfZ6FDK6B
5vDPmO+GFWKwqRFimUnaXT5+CP9mx5W0orZmV5/HesypxfDIQJXdI48oqj8Rb7Mv
S5yhkOrhxJSnxCHWHJbedT9gouRAdcwyko9GrFBbnbvq2+LEuIdKcGd1aII4X1uB
QSh28CdnDDFcya/WUgjuaxc23x6WympGmyk16kJiurKhl6tm4lkQg8HnDTFtloAw
qgxmO9xY3sdX9hHgizOwcrRu/7c+bJno55RKSds/DBwTTxV3FIBis84beWQ8y/Vn
X/1x3Cd9U1BdM1y1yTrvmiYX+q5prf6n3EgFZmk3danJWF6BczpslXdPGkDV63TB
TlzuZ88tN80SbD4LoPoKPKpQGVjoAL/KD0vS5uibaSz8N5bXirnDAInrKhfBbjec
g2jtfEKYyqJcyAvLGAP4lCTVNv8YiaVmiI4LVdHJzEenQ1NwlMtWr2nieAWE85ah
5gXzEq5TsM3R1gK7G7parWd0w0T0cCBkK359/GXsdrTa4oa+2EEk0qFoaL1N78i5
AixmreTlXwuP/H316GGwt8wcsZzzOR79HpNLPG3ePO9d35TTVvYzwFM8Nu6jQ+BK
duroEu5ch7HYSOYDBxhJTwomE99GQ/TFdm+mPliGdCWespx91MRWZptUUCJ6FWF0
yg1Marlviy/teMJkUJRuw8co+Z0bRvmwpShF7swpgNs9Jf23OksK904EIzc2g9Yb
H2RcCCwGwQCHN9zaaMKWidPwI41DmIzNqDhkjwYZk3Hj369xaywXeH5sxLPXGCNX
BqIEMY0j2N/XMjSvEGtmXIGV7RNYrYh6UI8L6Y0OO5pHjMPOUsChGQloRl+Qrxno
Eec/ArQyv2eYoVpUzALfsQCv23Kjfswhi2DqWlCJklGc6BMJ9pw03NT+Rt5KJN9x
Rt3WkdmAlG9B5chZrgmRMMe/OlSD2Oiwr4l/Rt7QEjOuR1/59LGr2xucsrB3mLuA
qQ2QQWhY7e5OwGUaGCr1kYMMPzxjBiFAMdd/BU0Z/vyVi3Kl1lCPWDgtjSXmrzKH
zgveEyPjerM6yH2cIvnbqLUeCP7HjbNMz72bdL+6XANYSDc0n++RH9gKmWw5HgQV
uKfkHKpcRJdr1m+BAWmG2QWRixzzcw8dLZR5lTndS6oppByFhbkjlBmrtpqt4MOv
vUGrDZDHLx2sAIydZxLFrTMw9y00dJoRHc6RFOGDzN+N5Zf0zfaY8x/Qa6DVq48Y
d3O9qKiNKqieuguD4FnJ72Ob27oeIk4cGO8TCUQqovYefevwKkuOTRe4mL/sX/mx
KOH8h5dSHG0Q3V5hG4AeIwge9/9QJsj95+f7+Jmd/pK5JsAqASPlJWhJMGpXSP2l
HsYaygeAEwRu4WtBw120mPVRdurFz31mKHDCV7gJBcPEbbEt7JjlJFz3BQ6MGNWo
/UgNkN66CZ3+LLwTjZH9FVidlC4sbpjdHdbafxp8718TAs6TqniNV+h7qaHDtJ0X
cZCneO+pwLG7wu9n+M0rznU0LJtDHq6dJF0t1xsA9PLHM3CTjGd0Od+XNmBFuDRW
CC1UveIF2RBIdfPoo0Nbr8ycyBoa2rjDnpGoe0bvVQW3xlzco5/LXvoeC4NjDx8g
nRzKH6lK8UiEYBWOwXqdKU4S9EdhP5v5cg99Cq7ftnFgtB5dF6tg2OvNPiwU98IW
3foJaJxAflaeV3gzf8JRes3U8pvZy9m1ZdItYeCVBj1/Pr4QKy/M5zqFu3Kk5lyT
M8gC9ORryrfssExGjxOMTiWO98Q6FDiJXyoSDvmVTmi67HikK92mrUtlxKihvFRB
q+77n+gpz1lkrPd/gz4i0164f67tpRJLDgS5XLiBRt+jRGZIR/zbWyAVgTtS/k7r
plTp09XzzscAelOwSQAs90+ci3wGJ/A8Bkcc142PgRWnZg/O3fkgIGSTgvE86iMw
TU//eHFjCmkmeGP8PYjxkJ7uBeYmTglM2rAg2uMgAXdEogRS8BjXQ5/nywk56RJz
AlQlwlcFww8a2/33uq7d9hPfjHBRG01qRFgNqOZLzmrmEFS/QMHKKet2vQbXEsiT
B/B2qP9BJ2AHbA0kdaa9JKfOQt66eLDmBG2kOax4OOdLq6WNVKSSHf4FKTVMaeoe
MdAB+fKtvU8f/cPtdurorvC3yrR+kgqdXhmdAhXR1VtbqyoS+MBml6FwxEHtAHsi
ugc3j2HCNSDMVcrYe9BM5s2fuV0+XQDpl4MjX5PcXE2Zj7C2EupT13+0acayefzf
p4dS7+8ZWN+iPnHsqKObqT2n1JJwLcfFzdRezXMoeiMSSTxphOB4NQPK84RUefW5
VWtKABxz0yNFDMeV8BlBNxs5P/C0TuE1lk9Dhxff1bkSTdIEDk/srUsbbSlo/qVF
dAj6aGcycGC27x0TJQfCOhAgsQ3WcUooWe5EMif58/s+DUK1qjZ000Ftszj19quh
GsH+1fMXpGfNEXA0q4c9Y30QTIcLJIBEoQYoszdLFp0nZ4dtySZGtbAAgA6oM32J
Q7pmtlU0XnYoOo3ZwV+xdQ9Bt4NF/XNT9oLYu6sr70qw/g+aeDX/wAYVWznzWuM3
5mFu1wcKkGS4tDpA3EJZHNiDOq/G1X4wXsCMCtra/8OAUP6ECnAl6BF6Q3Z7EXuu
vY1YG7Xpilaa3QZj8dSNGR9/1TQXlz92ChUJe6+K0eDRZlq34BXOAsWkkPVDQyJr
Aqb5VE/ObnW2eFf6tp4kv+TkYIZAz8fMcnLNNZ3wnkY35whVUAmqvZLLfgN8mZy6
m42etG7vYIl3GEyhgo6UEniycgypvK8HZcnhdERUFYcs69+YLZ4jIsjG1Yydspsp
CjRgcUBDk4wWdwFTfLTJGJUXs6x36YwMRDHN9QGyIbJXFCHPHEgrwflYty8F/ruV
z6oIHUll9M1+dzE+/CCHlMTczxs499ePmftgfkgil/063LHf9F+DjzamgTmjOluu
8Aq1budlGfX2Vqcm2rb20Pbe5sCEbfxWYS5m/bQIRoTGtTr2EI5MYyJg2q7RLEu9
DAL07/LCCNwr14Dn3HrlKGZYoM3VdtRcghws1+QWHMw577PoPYUTWVVJtlsNo9+j
bydRAowgsgc5ANKeFYdk7MaiD8PsUbXcRpZA7+WBNADSu4YJPYn3iX6A51+4DVrk
Fc9oN0rjPYho1FmsQ6C5UZLMAqDJUZbqTW5eLUJQSfV5rbJ3WgzKtjKlu58tZd9e
ZPv71sYa0fRmvTiyZiXo2/uZBsaI16e7ZzSTYfdUGhAD7Z+8Hl6kwDyYB/42zyhA
y4W3pALAIxD/M43BdffLOmzKhIoAPaLansrEgZvJbUPF5wOxuziseoimwiOeZu+0
pkuzEBdKLVFqnh6M7tr2rGZRE1hgXMdQ9joP7xSgb3kTZI6w0ayjnybJ/ocvjNMj
vMAXys7fngYiaSbW+vi+4t4w66vbqzbywA1tJH+pkGtFAWFdIXAKZyj/n3PhdvsI
sNegawzMqrhN+pdFyDkA7Elvb2YwrTcF5rcM7QSfukUmWBYhuCvNanRbTNWf6i7u
CD1xs4gMfMMfgHXxi1WnCPiVG2buBAt0qDkIPzfYDhJP9cwRL0LA2NwmPJB28Usv
Wq/errSuh9gQDYOiumliR1OX5lNhcbGDFH4ULHH3bmHAd7k5k4hjomZYcOjTisQh
vWZxyaR6PrYk4AKhLWVb7+jDHL70tAD2i3zZzNR1l5+QsjlrjOI3TTdCGgCyeZ6A
k4zESWR73AVs3GBQbW+JiGT2khOXiU49geYKGo9uJjuEeL4O1JODpimhNdZt80oQ
jfDMxoSv5jBoiU3PeE25mpR7Wn7g/rLbUAw4W5DQmyIHw5JSIDBlJOZ/PXL2syM7
4yK6BADEmDDRdDG05ipxjfbZW/3l+DdWBMiyN42g3+PX9uJXjgEJcphtbrgPH2Ci
gIga+ReOtWQz1d8ueV48ll3dIr0uQZ2ukOOBxsxxaZk+xXzof93SGDEtTPSK4knZ
GK2FTVy1TOv8HNKHeTDIbIUPcorCwYNTko+/RjDdo1aqb8Fu24B1IyKZt40d3Kfx
E9O5C0EmQ1/llW5L9inYByzcXYWkyw+LlIfqFnC+EWG8DYKtfW9RLLHJYwWp4BV9
k+xC47X7x9FQC3mk2Bc2S99Nn1S+LoL26r17af5ZyunzeXvsuTJxB0a1oD2JVFK2
4zFXTwXTn0LM77Ed2v0993OodhngUvm4K8xxZdq+YJ9pnTOnb5Me3MuTVz7f+wan
/iHINnxJ/AVt2WLwCRA/KV6dU+bmFlWb80noDd3GG/6YOWZFoHNZw/vxvzCuyABC
Bo6YIxw6Gw8TNPFMe2xPSYQSn8O3YqpNpGDOzc1vM3KUMAS9xM1KdWdEIxLSFgvg
S0NuWdYYA6hPBjSyJAqaDMnXEg4GuBM22989PoAUBf1MlozaTHp456LQVt+QLWpI
5YgHBW+nl8RAwwv8nQJ1aCkmuZmUVgbAReQvNSElLbfL6c7Zoa7ws5mYmGwrkvj0
Z6jX/rh3MF5f60R7i2XuKkPcqFC5takDK9ab2S055EKeyFd780UPv9oJJ/MIj6EB
QoykpwTsAUiRX+epziqF/e3FH41m24hBvPKUDIuRH+vogqyTuoJtMCkJ2Nw0rJpX
vkF8RYAPmIUj4zeYi5hUBWhmtWHZYOsi9mGiGKqWeirS67oLLfwu1HkuYdkrRNtK
U0RblR0pim+tk/nWRjKklrXbjTsKt8kwogFHEtJ4z1eNPZCzxzE7AJYb0pTpmN1Z
g21iM3MPSUHf8b1TKoc8msyvKF+Ek0NSar3SsFFZFi1D9ws+lgq8k+QLAbYfhvvy
9TrcGqP0fdIV0/qCs3pvTa47PJm7faXtVhI1mwuW9XnoLtKYD2YCS2MPCY3L9+Ms
Cdy7DFVBbiuMOMcyvC6/iPAM9QxbCyM0zB1QXTP9OIgZK7QiJBGwuPdWOvx+7hrV
s2BcLkdoPwI8BiXy1XPmjOWq7ckWu1LeUYyy6hvWMSdxODG+HmGB9oVRynz6ZPZy
3wlVIR33OUgc5/wS4MAW9TkjdRInARz3s+DmOALjLOYylpstv/xqKypiV5bWxi/K
lBGCsxoNODIYVcYWgJzN3Y5DjDCd5YnN/k2ZjAzxKUqlRVd5J4iWGia9WdkLuY88
SQwjJhNv64ZzvzClIslYaMYmLOJ64HMzI1seIvh/M+uOdbPlKWnA3GFcaRY0/wLD
MgHGtL1I5j+UocNS6PPhPzTXQzaCEeu3n5wzEkSvjw57WSW2FywLr0UKhIofhJxu
UAtByhNLzHbqZLiWFvG0+ieryP3AnvY2MX+JoWdn52IVUMmr2f/I6K+3ZJXzXgvZ
N3UvWLbdcKf8gLBJqZzoPVqR44Vh0x3LZ7x5cEatCuzcJNtXbj/k0QVV+SBTv79v
lwDGqNWLM5F4ZtBj1+/CSlded4RWMIyq5u/2Roi/k2dL7Ztfmoww92nSFTBI8NNq
3/AjYa8sdE3oExA3NwzmH1fEUcH4LluKZkBdo4afybQ8IwsWbw89lfjP7MXckcZb
YfExQNzA2T4dSlhK3aU+Ix0weOL7xx0F9uTwIU+Qwhm/i2cKolVDzKavouU9zPcg
zF0K9fzrJFhbPxP/rTScxP5q9hcembnNoViZvAeKr9PXsfRVY5C/4nWU5vKOtrK8
q5HJMcs5+GqXe7eOPmAfYOPhaGlfm0LUwFUhS0OolTQJxomXr3Tk9MVvC8XjMQWT
K0lF2FNtVeXGnY/n9XPmx6h6THfhaV8Kul2msrfTkATmag+fv0lA5vQqmQJKSlVT
OxiPGyw3UDhYKNsPYFMUdE4PO4Ye5dFJG69C+O0p0WglUBC1z4VDprUIx7ZnLWTD
7BemCMw2Q9j7kX9WWdA/uSNgpgas3hBXwRKDLCGFw3D46JIaFHLa0cBp9fHX7tkk
9lOrsJQo8gYkrlQ1dzjKLajW6wdBfy14+VYWrzwqSkYoOiBX2OEdHOgcMMBK79Sl
DazrUI2j0VrPb8w+nMvLyx9oJjkxfwc0A0oY0IpZamRZxoa9rTKqaxbe2mM3adEr
Edm8fbyKcVCShxGhbX7litbWNXkb5Vrg4hup/T8+1R+/IKqdvNuxmsUJJBefya8e
lKonm8g6OWEv5VDGuLGGwSMh7vkFhafqooBVlyOmi93g8ByRUAUAH6bjlx4eHwua
QFRJruz+CqMhPwulWPJId2TjIQPU4FNJF6j65+aaXA80AJuATvxxzV7ZRrGdAJV/
FqrDU0douWAvYrPerPuYvuV6q6AolAEUPbXf/P7hkKwiPbR5QpYHlUfO+I6lyuGL
CJPVzGAxZX70AyEy4mfSqPCgXuVK9iz3yXW12Fy3DWn+lXz5A9kMHKdIR+NPzi0T
QhWBkKHk0dU3Lkfw3TfNlnqILwk7t9bjk+rDGTwtgl5M1KqvuIu//JVWECSmtzR1
EM+f7YaJP4nDs+C68diRZNiXvqZIW4zKfM5WHdwJb62NcAF3FpSPs1gOyQgqhoGY
OVLtLcZN1CKVIseZECLel4SzG7wYpRDSLLzWMUc0G/8o13sNvKPCN6NkzMUv2HiM
xb9fbcaUlf7aY2aHYIZTIyt9mE6hZJKAYi/XcWrbMHq/77SVrbw5S5sLWxEJErvR
X2IWRv2y3z7nfaJi4LXryxa55SghVCsvi0gK/Bm0TsaufX4GEn0ZE7TVreciyie2
0xbTm6eFe54het4CLh97E6khuur94Aj5esrLyaeVehR4GHY0hqn/hW0wQD9I4/W5
R5pYcz2Yw7U1OMAuc7lSZBRMKPtPyX6MoMSZJuvqSmKie7G482LG4TNMVnsJmAmZ
w4za/Rm04PKzswamrOb+wgF7yE2j0k4C+FRF7Z2/+bb4P/LgSGImSI4t1JJg5ZCz
x4AfujXGctz3HYhQjRoiVo5UZUt6sU++jkfBBPGrqgy7dOQOKoqYpXrityKLc0Vb
jBKDqDbn22Zd4Tz8d1jHeR7Ce5+pwLGtEKaX/8uZH6nFUbSrY1LE3IR6MRziOH6x
GOqdNoYrtMJSop+5A9Z8S61jWWO7ctRtkPXd2xiwk11CHe4tIO+Y1pNEhZmJg0xj
pl4PJIjcf8FR7OwtEgyH8QWLsEr+8Nyy6AMSrqCJcCoADOom6LanNKwUF8wdLq4B
bSW6nSQDZzd/glM2LCm8SZKVcGa6c8oUOskP8NOpmKYujZbFH10UyBBvCLfa68fT
JFyLVe90d/pcLq8oE5J4acTjmrDYAfFOFp5pgnsyGRNJ7/VGKw/4bLmxVPVctlTb
r/6Sl6Z2RHJ0PHt3GXOcSbmNp4N/LdgRzoI/iRu/N4mrstIHymjsHCK/hlfKlQAM
8EN4Xenl9/tTHRWOYQTTh28uJUJj1EhbR3qrFQ8Yx3urU9/1LaUe16ySL8NCn6FT
a69XCFn7g0f2lKCc/s7oDQzBOuqFSVUkFblquNeKWqZevm8kOHcMc5Rri/0RMvIi
Iq84AjtfRd4gYrYX+kRZYQdd0H8KSBokvge1ksh74q/OVdOtHaQqTjDAhua5Kx9+
qoP3nNxQBllmUORxXszuKEbPKurbbsxFuJy+4YnJ5Y7H4+hAoIZl1KsM/GhzEo4R
QYLSYKxG1yPtk4CYn8kNYWTC5eWW7QhZMslKfOlg4sdAunowqd9pl6HYp1I52EOE
MPC41d7JhbjzjE+3xRRGxJgxvNofPLU/kPC7vQfhutBrlaJdjX8qn/5X2mFfhzgH
MvOp990cR9yxOzs+otu1fiiLL0fc9rMyYswa6cyLpuwEuXw3efD4+fUudInJn8HI
AS8E6w/rJHhbzxxECOkLG394+YQLLjboF/7b/1ur/KjqD+7XAF95B0Dx5p36VOAw
fwcrxK6ptYShbUAZzcgyGBmXAGFz+iy07Q02ktmmet17RDSPUsK8tfmlQJIGStOj
kLptFZkXfXUWdC5dzpKMigKzJtHxSL/4Ln9wFA/JSzbQAb9n3KhFvR6JSAffnZWS
+k5NlZ+TJXwTXQgE+lJ1+How/X3viopaXBZ3rFvEYLmReXuahvDxBq/6wMVUARUR
vIsmrQ8YB5ua6FntbhBZl4nSJD356Pm/GG47uV2CCxNJFe48L3ZLkfAYCXPg2Vsp
FFTe0jP1WpU/4ryPfB1Fv3KDj5yM6MQlALRkPP1MYJPpHALxraBf7DnPL5xdMLO6
XKnBGO/lTb+/qejkpboBA/FPualkIHyVIwamQ256wMb8RfhXf0/3WzOyBKgUwLDN
W+EaY9JH+ArQ42z13St1Qz288ymMRwpl1Mnl/TsP38o5NXYTpzAoZu+snvcbFJMh
141KyYJtGTqRtOpqjf42HwZFSyXUWFl5RPC7Ry6QO5w0jm6O+9hULESS3Dplm2z+
i4NSBKulwAB3Y6r/B3hGpsnnu/rTkIQ+ZPPSKyOME0Q3HOENQsnO7sc8RcGtwLk8
Q6xNirqPAPixV0Oif7/yMAAmmn3yB2mM0QgGkNRDHzoRjC+ZF7zCSyW25nRkqYxH
QOF82pV4upESCn19RmkY6B6537z4JVwzN9jzDhMiTOR8oV6Eb51Kv6XgHc86XQcI
SOn0uSAI+KE8lxxvBfyLcY31UJlRvPGNTF0K1S0UpngOVcKaoqsoSjbm0yblKFrE
3paquetD+rCTtsGIGuSI25FdPu08wztobBIitcjOwi1x0uAe7UVnDogeRG2zCeB0
gdg4/ByS+s1wDNiMV4snWB/VXOGlt7EEz488zmMrk1rj5V4Y8s8KQUMpcJmpmJVq
fH6NzQramGhWFnB1oNM6aoLqgIeWSBnHjOIZkNASGtVlsxqmZ1WHPRC2tvHnz6u+
yshIGdrU2Mot17VF5/crCD87imAvJxBFXErYzxCkR6hpugvWHB/jmtiONQ5jNmjR
vJbMtdIdd4mqjXJv5OvROWsIYOOP+BhL9dbt7rKlD9MNK8hOD1b1CUwU7/Gr5B13
dUthfDkbRsWEmgxqn1IcsgJHMHuYTuBhO3yDM+t/Ht+qi7z1Z6C32K5ONHELrgDM
bM+g3X59QaLqZt4PO5YaaMjiDRdWkKSm4xl6FG4msQTa9R/cY7oTg4iMaECU0ZZp
E/UcfzgUZhU3pshwokGimxdqahOQq7STsznN5+ODnBIVBwmM04iSqMXDzcyqjQZ6
gI+Q9cpTS2hLsPZfa6Ds28zcghTgo0+FprBVXQVj8nq1yMKAz9F1Rknbj9grQic5
ncy8rU3/iehsOb4/0zDS4Pe+w821tIUKi8bUiKtpBeQHkfT9Es3c0x/gNpIF5LbZ
O/boBCQirGgAgNX3N381wNJf1IXYybqxw17ZMRMPJ6VMsW1NEpvE9yBufX/pCsT9
/x7Zsm0kfeD9sCNJGJxlveZ1LDHv07ZBl9QbX2I/rb5sE6eCpMsdDLdLSpG8lEP2
eotpkxYJURWpbRiUQ+H5M1W5/1Yr9VSteGvz1Dl+9xD/Rjr055fVRuCtqQhQI++M
VkEiqedNcyFKSPA78S2OGDslEoPzl7Vz4Gj2/DDOZWJ+sy8QaXv+SUMPvPa2vDid
ec6nHayy8mvKpS5uCViSTJV+6XTjTZNoLm01uXzKrz5uSaaEq4bKKQ0edsRkGHtD
cRvbYqDdfCsqDvmY7w3mLv4+KoJl9gfWRYDRmh5Dlo6g5Cy5UabMPVH6nvF0f/p5
/xY/8qZG6uGmQCklop0IY3iMkaKPPQv7F/s5jTzoT6SzlcrnTPrAcgIJiALA52tx
U5JfttcirzbPLEwxbRVnjyxdH43lye2R8+P1JQqIgenGRrDNPl80tGYtmyt2QtBT
tV7JhOSsuoZqD3yLbBVWS/Tl15XX4mTA7f4DQZ4Iv/ENxgLgNFT1yXrL562evFGU
Q0DS6CShm8q5+8GSF0+YE2aBdz2TqqUV+3WtfTfASOX/yGdBxupR4SDxI+UqUgw/
GbfpcZVIepmNUNPXTB5rR2Cpld7VyRr4lvxgP4syGcgbeEjsxMu2Et7vjLTeNO/r
YgQnqDfMiY/YtT+ICQ/hlCPqxi9gMFvnjCE+YJ79zu6vkw+DjnOExxZVu1+zYf58
RD+65zj7rQ8lYl2clE107rTApGe+w2sAal7jRWryl5v81qS1FsSx94Mnj/+pbwNG
AC7BJkSVF3kgEZteaKSJpB1zo1JA4L9i2Qgq58seONNoMBLRGbPI4QEUSwqvF0lH
3gdX3qn+yAi2HTZF4XQTAm9V4uBUEMbABvCd+zDx/0sOQEymSWm3adOHhp5zJ5E/
Orun76sS8zcdhrlN+dJA7bzECk7gUEJ15ESVVCiujrvm+l6P7HlgT4WhLqburXPL
IpUfYwuGrElKjyEnxtOKLwO3/x7ZP21AVCE+fsMmUi4JvAFXjryD2C4wtdw03erZ
Nwa86uztcwPzD8Yuseme7u51vO+kEzwJViufW4L++TB0O8hVbc25glMrsK8eoE9W
xKKa8RoKWpWSOUtHm/5thlhn4wB4bzJOAftq+k2DZVrHgI6aUROg6fbamZwmmgCg
tsXVL+xHqd5NB6k6VjabM8rgNJPBTvSU1lU+dAVebXTuhwdpUYVlxRhGD8P/iuzv
u0CzA124YwLVklD6X8ysOeTJLbPzdVkXduc4qEztGrV10S5SoHgxEdBnbr8bn0AD
4nKGkIZqRC/JqY1dc5Jz3WrZsHkdXbzWHO99FlBxyWSVqmqGS9Z8s2N6ZLpGZ43o
pdO6WUxckZTm18ASNojnAFiwgbvjfOCj5Zd4CPSoTud69zFhnWwxaHeQ0a19uKg+
HQTcKngRuZWyQBXBR4TNL+yIuRRg6HxQqZJeSDIls9a+hMaKKGREeLPQQXQnKQup
yqAdeg+2Lqavmw/RWtVTQQUHnCwMM5SLCPUZDwWArfIpz8VNZO8DOLvLCnaPwTZ6
iBteWXkDLmjtXyu7AlFk9WjnHQEzl00Rb9aLQZMWOW/4zIM/u0tkft0QpMrS4W87
mD/u+XbWnWWRDhqa/0kAz9tpgYgvaKpwDB/eZAp+KCpHrVK9CsYg6/2JXsUmq/3c
ObsaxKWjnFmEKKIQzlCznVwVUS0Mo5BJWTfwm8er0VqTo3jgNR8vX811oClkH3S0
yWqI7UBW7d0bPowKQMP4EcBUFRaB3Q80E1v4cXnxLIioQvsmJtRiL7R66rvr28C7
qJWl7O+7EE32QtubL7OlnnLCwE8cqZXmAyOIvGTT8QTvCgkeyHH2BvHNY5p4632Z
znihX8jkSIVqpS2GMVu1aPyVIwUUNtUTGDfACSVq3jh2Y66w3JnS/xaa6CFYlmUQ
6FWbpW46onM7C9zHf+VZQzEp9yyniV81m7OutcxcJhAzuGzBbXikY4hudvU2V5Kx
N2QLCMuODKFzXYPmvmR9Oz2VEm+0cKZjdAzb1OxZhtUssnZuUtVO7/RU6f8F/hXz
w/eDbStFXAgaZ8O6b8raG36H6wmGW3o0utvOFL6DxtOYIoXpPFO3itzU35XBIXim
h9ZvaL8ZjlORfRUVRIyS8QMMEJmnGeHPGUw9Dm8i659C23neVsJxaK/lN9j6k1bu
pdSfi3B7Unp2Sae2ac895cqEy7/0Mf5H2bErKXl9Z0EIjUymWdYUIMJiepAhLAO0
ZlpTfqBc6Y8oa6iYZTBPqRCRc649LPxufYz3V3nSRL/lJj67xr8VhxLO9ZhiPc1q
tDMXaf8tRBtnhkoYKgR2SwN3ClabjHrvbr2nFxEtslO0dS8tNqteFopIffaDF20+
1RGui9wAPluB4WHgeLSXsArXzsKp5SOWQZI0hOjxosWD5cgUGTPPL9D+5KsNf7/k
CBKp7RYBE9e7Amh8kodD1zVmuV0FCCIGq80jkijTYP5kXC4m9Mb7sQ9v1IkuVw71
EhBUSpgJtGDpb199YageqTjUOvnfOEtjIGxdnxDxkjlOQCsBiyU6dwuoBAmguXmB
8FUX7OHWPQq4IAJyVXk5gyRnr/1GJJIDv+AM86Y+lBj7YmubG54RU9W6x1SMs+Ol
zf/R1vWAmBRmOWcJ6Sq/q+6FJuevXGYUNy4Oci5HfqQQYZbfMEAInOgFWTiuqfVK
FpSsyMzQpyFDZoRUOTWRTZ6xzzLZ+1UtQCpx1nMNJX71sU13q7hvlgUzn5GabrR9
GMHVuMh/uPF6xFfTxxE2jn7i4v6ew+2Gd+Vaf97W1KJSrbzwYUO1EOHnBG7fzpYi
HHFj/yekySGNZvd6UHl+LitspfThsHBVHprqWXnQK6Xeyw8P4VzL9KppDWQUtsQG
e3kd/NMWR0BnMmIaMkQ/gAmdPJYM9Aj9ULNz38LyWHPTT+ezZNx9gWAoHmCbl37d
Yc1nFdQe2O0opEvNt4UJx2WpeRz1oSpjEOmO35AZXgzJ+2mN5erBBYfNfT93KDZi
d2QreEovZu79Ut7vIQ9GrMBBdagJ+fHGfQOLMBQ+SYRECDV6oLkphTz+3aJlEk3F
TGxJm7/RIMV5UnNlzkW4M3cZ6UzuLMwpM3b3XZ2cHJwe7T4LIfqpni/BAKapBoUY
GAG9IdSXZUk6tvIo9WD0SAa+AFrd1luElf2NQ/OwcjgF/+wSf6gNnHR/6PwCNKwa
6XK6madSNi4D2ReCnrG+gVlG8xbTK2mGJ6DtX2aGCzzv/y76VzHlPT6EwJihtqKN
mpNMNPlbtq0aREOQNxCokMuma3Wq8QxUJyCGJdD3I3TJFRI9zWxXwwRxLdQMOddw
mA7mYr51oBz5khlgKEkktb1yPg5sn9Y+SeEv3Z4kodJsJ4S4UaRxX30ZF5AnBsJY
N7/D0HmqaXGlLHuKkIo0yWJG3EzckDPDO/rLXYwgbzou3Evi6k0kUovPnwVBAkAG
MLONOk0Wm0WkdDOVuQTvy1WKVe0rtHVmG/S51STgVvR8CID/0cfrBD9Txbmr814w
hiwckGzq/xgJnq88yVCbCTHLF3XBIZmqK5wo/LmX9wHCVbyYNMpuvWNqsqYbpfEo
EkWaGT7+rif0lIRxy83iksF5/wFboxo8zgTRL3bG/VGmJd3WcQBmNtEDuULYedyA
mvriSx/W6CgYFDeBiPpJOLvql9AhWckcTuFs2Z//LVvpgoQWaDWDj8kKCIGEL9/2
jWieGVV3Qs0urAz/Stfv5QAmWg8Qotod4fMR2Qc+P5zJF/9CqvesNdD5SAGDl+ak
wlBFik3AkODsRtQmfK3aAUt5Bd3jrEdrBLBVNUPNGcASY8sfQp/jU9PjZ0IS/tUk
bmmXYTnOsaNQ04FQ/Izz0PxW0ltq9PPbGVYd2za85gKqMeM/xCsaa50rKbaVTpNl
6COgpeafQ0HtqHACzHN914tOmyGXqiCFNfedu4tXzHJJVycJTvq3AOSpR+3F8BMj
gFPa8/VmXaG40lnBbpM5YSL/zqv1Vb6F0kSTmf1qUy6zPM4+tlgX0AyFcUBTDcFl
6lwufDr0lkdyvYe64Rn/aIOzQ71R06rJ4lp/yRbs0Mjz5XSon+9YUnkSdvKsMRgA
nqGCOn7Cq0ARQtwTupFIRJTMAXYepc2UgZEMPiHtGB7RGON1s01GD0OK1N/csnef
GtgF/c2PNt/0+ZMfcRVYUgD7x52qloeKXetWdpJrIUga2Zbzq2/N8JgaYdxmhZp6
ly8RG4h+5BbNclaEFA6UqhvCBnyo5U+7A6voUuPIV4KLdM8UJeuYL4ab95upi2D6
rmOweZ/1YJDwoDYEH9xsVDQcrj+hwozhVqNXFIrjT7QU9BD8kaFJ/QJnHl66fAoD
etxwpF4gmc+h2/NOhIf2joGdtPxdmxBz1BI47gk0r82yQm5uMPZcnpgEsYbqtalk
ehVBH8Y+95xHoxF/FRm62Hew9jnz6YepaoYunBhG01TgDOf2x8uNHkpu2CNrA/WI
iq3L90JDI3Fi1NNQzHDY6v7eSmascY1GJUxEs3ZvlF1GZrbWQEJ2V1bVKqJyq8az
cBVo/mnYkvOg29ProRKTEQ2aOKanLtYIe9EHf8IDdPtE4CdX5CdtWzuehiJSFY03
2VX43ptuB5xCjnolriO++qsw3yiP3hpe3rh76+6QmVHHQ7op9NeSzipxJIvD/rmD
TsgcoDErqxKoJuRvpmPHEy5I8+JDWTwX2Z4UvRreboacOh40JiJ48IbDCmQJsZRP
rJKs8bZF7YJuLDm9aTiCZJS9Rr9htEnyaBRqd58JLt4qqU7S26U517XZ5aaGkbFG
pKUlO4nQv65gdhH9fmVe2lEK3RhyEeSlvjjqDyZ5FneClrvRLErl3HZ1S7px2VJV
cjDqW9RtgCnbynXmLXzuMEmeJrs5TXTtmYPIm3x2lYffva7ZcgYZ126LZQGE0mjr
LgDeD/v0S1wmJfcc6GCjX2xIyZXsg4jJ7Sm6glUxQH93kaoSQG2gUaHkqvRqOk0G
e9oaypoo5JFFRFtTx3Rw3ViWIA8h/uGFSI4TCXzMgmWG65xmi5tfeR736laX+PJD
/oLyxj8k3HHF1bQG2pALhB/yP6P1D3+d6EPxrwW4mw3IBp39cOjNq+SyracjbUzk
uTxZkqwGdZijiWHqM4/eTTZU1F9ftXuMr+d93DPWTKFmUSPAp+67OBWpIOmmMdVK
eVzesf26fg+itdELYmbBZViWN1COvNr6uEBYiZYHxsKb7ufg5Z9XztG6pQObkMi+
sbMLtd8bgQzFiHgWfoMbhChYjNtY/93UCOADh5Dd7NSuO5cmtVNOlIFn+0c+wWrE
HeIZ86lmDnukBiOjHABnQGqRTU4H7B6C1bUt/5pKvfg1tpNYrXTMUOviEK5hljS3
AqpyQ4lNDvgiAC/ptzIEwBRfnSA19XjGbm/lB8IF3G3oaUySrp9MvUS4n5v4n+MA
eYjsCYrIW1lL3hWYW43KqkYwfuvwdX+5grzf11g7ssxnXPkqvRQgsZW/2OALjuxG
YCrFPxbGlY2sKBVLp1GNO4qQZ4CWFLgQmKGhWpQ3anv334IfAHz29ToWDYBKJAnx
QydS/AWyyDdlul5OlQLvDJJXvbWf6sw2989MVdalRNm8l2bgtN4Va82ARayLyrq+
L1BrseY0xj1eiEokRmsXkgHkyefzRE71AH7o42qPv5SJjVjMSRsqBjFqrSkP5Yei
P6V5m1zEchu2KPjjpvWpkqye9+hNRVnyHP/C2GQUOxD4ueqoUfmu/vnq9QuYf8Ru
0ZGdNWFcPdB1rl/7JLOFx2l/gR567rINIg37i4e1F2KJ0CQrx+OrfekNIJiZRum8
oomEDLg6gwUVbuHYBEKe21ENOd5eriI0wkPDF7uiP5ANvDP9XeRw+tg4rB0wjr3X
+CMnDPWRpLq58ZqeWeYHk3AZkh4HZ/2sO99ks28pF3i6OpLUIiHHSRhxC9TcPCH1
8hKgX/DSmjnxVn8VcASrXryAXuc5YLhWPZTs/q2NnyXGGA8RtuuPKsKH1h5v7r9k
xOqiXem8CREmZA2yYiPWkvL+WKowHuxIeg0aF4jSB/HVxt2+rGVPBOk9+9zM2Qga
f+ncZll3zRUJ2bgw2wb4ti75aAdqARseYIv9H3f4w99i8Im+C3S9rbB4D2geElbs
PQ0U1fBef1EBo19goyIAR7iKgf/W82IqWpF4grO9w/0YRrm+V3ocZtS6tihiA5Nn
Gm/DM85iCfhfr7jXlP7seVZc2QsLJixbR9HidHCVoRof+VpcM06PLcz6vPmb0adX
h00l6r+cL9eH3UmP0ETgN450xMlwh8iRHh1kaTjCBlYxjUfLmHLU0+OfBVVEvJPj
GuIYpJdigAeNLM1BBqdVDsfyKHVpq0MIvY1ceFjU/3kYkz8jqZ8hxlOsm8Y/aB7U
2G3J9Nveg75Gq/VVSY+b5NitktKJe0wmQC0SsKBjkDPlpiLxJZs35KmUgZqGlgdy
guDGLZ7Ja8XfDvTYtWtNCiyEVaOqSJaKY7ETS+YHh+W9U8edaqFQG1eXF+fD+zLy
R+ONFfpZCgnAD+2JIV4UPW9+3bt5018jvxIEVaMG2PGfBWruzTATs8YjFQNsNAdR
v8E9/YJSZCNizuyDtQ65kieK1zUb6N/tBgo5ZE+Vs3hGLzksrO/duWjGlFqUsFYJ
9HnWXM2VAyn0uVt6bYFshGxfSN1b6FqegNV9bJriytGCe4IV5du7nk/X9gipEZvm
yTKfaFETLzSK9XBpH3N6ntkKTePzjiIHwJ8dWZH0Xx54OYONo0TFIqUoruJL/waz
D4GaIvnKottD7ZzedbNWsR+2lijOmVXhm0he7wiHqgvpAEay5ty685c8xRNjgCMk
8z9AE69rH2zTnEdAdKnzMewNS74Uzl/BWeFDRVHCejxgDq2rvHiD951kcdqGSHvs
PSc4RpmVj5bg11j5DZFvO12UjvBFHMWiFq+jIJbPNZ0Mih9t16f+pTyUSuP5HxSO
82KeL4uBO8yhJlqN06IDemtyLgPqxGmcXWqs4/8bf4EtYNM4R56y5Zg2CMpEON+v
SnsqNQRW196i8FAr2jDvD4s+UQuRYvB16js24KDgC0BIF/WzghG2bbh2eAC3lqSO
ltyBLm8mUN/st60OZ6Ltz0gtyhTB3OZy93gzksgYulGyyPn0vPF7IY0u0ahVb/iy
oQ+XNp4ZInS5Xj4Qk9u/WPiCsTcKwddJDQ+rN408VFqUAIMerWjeCusEOuWqO8Mx
mSYqpIB664BHd3aBkebGOSPORceKUqiIackfI+b99/VpJz4JyE2rrzAFr9WfZ8wu
wk9oD1J9In9fRYaBdLAcjRYTqWmR4yjUlBTbonDuHH7nVTLCUEZIG4VCbpztDaOq
GhzHREt9BbcFLQR8GIoecUDpLuAcZyCWN5kzoX76DyZFIkmL1q7wOoJ/AQ2SZ269
ssSY5YtCq8UHP/Ljx5tpLfNEacfyv/8ed+FjIpvYFkTOz4lHm39WhGcRbr3QawSG
vW9LVDteOW5nXCdKigIB+OXo8Ye163wQuF3qVak4itGuBu8jN/mf85cwmz00siZw
OPnvwjz+oJ1/cO2ym6MMgBLVGkgkJvwyRxNbLomeHTFI2FY9c/dR7cYeE4RKCSD4
BZor39ycIoMPtABkIZX+b8KVK0IoQ/UNhjYPuznJ2v5JxyzU30mYDEQrB7Plddva
KJXL/i+ihNhXNqddSDMQfF3BYgZG3f4+YhLMuyO0naXseE/gQFwToH3AHwup942P
Lk1LpxIyw6hw5j22hbp8SEeZ1hFafyfWeaoUdbqD4w86c9cY5aA+Kwq2h/DBg6dw
PLPj5OHnmjnPlc+gjdi2zaF8Z1LnaOhCQ2lCl28JWdTNZOTywVsqr76VuejSKbpR
BN/EdPfY+kXDX50A8KJvCTZ1S9sKlB6DfAoauKzUE6fNcjfUHtuoTQ8PyM+xvJKZ
GTQhE1Ei+NJWIJmAFp1qc9lm/NiBFdE8kw01pCSUp3i3Jg++8j2lQ6va/sQTEpdN
Mb4Xy6PVs+e2k6jYALZy3fvjBVYB7ox16FFAjs5n/UxkTbSNpd3xFCJLoPSDyAav
Hi3VOpjBAJqCGOLZwyq78OCSikURe6shYvp0qb0+YsuiuCzWTEQJ+mj3PsX9pgW7
NO8Bg4/t6tphRycLjDNoaGnZ9HlbRZkXTyugOC4o4jM11oqUXqoXhBpA9VqTAyNE
0YulB2DsK/bXtjyw+03NAS87bnm0EgKCEZSIF7bIVQBin3Y8F+n+aLvPFGIWC+P/
8XVSZo/bolrrISuezmY/O31NvTMv6LZ9BKcmBfC+hg2M5rYvSmor8yGAvy/GNzeB
/r4AsuMAPSxyAvvd+RLYEdkjhLx7AiuxqAME7eBrIrzMKC0eVcqhlUmeH0PA2D03
G2jvUeVCkhzsBIVzPuBsuhEZCtrP3uenRjIU6k4hBJgYWvC95CzDaxZIuEO4hRuu
rlKZ+owpofCfElQ1Wa4O034kYSTkUClnJwOg+7AEH1YrK/o2qPcE4evlj4o1Rd5z
Wm6mRZo4IcEhfGLh9G4nCKMViJxcH9VaqHAULWZL4WdJ+ZEuXdCgFl3DxPDztzTN
Bvxs6Zw0BwxwoPg6lB/aFSPW+1T0g9hUXPKXzveBBZtAxyOcYbpFal7hTeyWE1aa
fjZ/afsc3wwRcVCt1KQ4+cGSl6AoZ0nLGYnkn8g8lAmSTQgZ59uzMmjaz/jWeNkq
gYw9q8u+xcs6Qe6ZKCa1VlX/utsn4lislRtz96vG8xEXpS8erW7jGSvvALtzA1fx
PMaoeVDzmmxjYUn2PdR/rrDCf4Z5A98C/lyj2LI8hALtvo0HzsPpJL9NLdPMgYyX
nrJ74HqLryMcQCF4ruaJ/H5rK6sTPE/xOQ7HLcuQ8/KmXL6LcWeRVqxHzstDR1MT
9NKv3t6PuW5KJVDa6kn9N/Me3U87uCnTq98xLMUOVX+O/EiXoCQqmPExwfv+kpS3
4u5ZXdlzZ6H/7mLo/CBOrplQibP06Afx17XfNDAqAhlcWfE8UEBpj+K8pcHRg5PC
eVn0aY1jocrJrVQu9D2ZWXS5WXID8fGz3EnJ8Qbn3xcEzPXsjnRJcd1be7orSL0m
9MnufAN/dVyp56djOdZo4zzs+wXTm/KFOSvf2UpZ0BoRrbT+BMLdcim+5ehRLxoP
km2qwFRclU117q1gS29X/3TyjRhzG3h8BXcP+BQmE6pzIcTeDRYzWN5GuAY4qufz
cPULI04+g7Oyi75aVCwc6ZLGOLXDzoxXiGwzuoD6k7Z8H+HooR5EGqEdEmTMZYrg
toQRDWkX0Tz+uSoHTX3gI2JAKpPaoFqa+gIKY0hknitiQj/Vh5BhB42Pl26fHyju
UWwm27SM/wKrD8wxRl2kyqxWvz0c85hSwFKMU8GnJM4kKYYPws51zy+17/Ma3a6G
295zyHzUIMmcyTMZEMULNcKpd3SiWmsLnEsE7q5KKpHOLAP+/AEpkCBe/+JQ5TBV
vSHpSm26TqIuIAP/sCaV1zS0tdc/hre3FdQxp7Ya/r8yFZH1N08glFuf5l4C44s5
3p0O6XShFjRLlbIeD3m5vAd8kN6xjRx8W6l68rp1CtrFs9oGqQmC1NxvdP6bhlhb
oXNqeSygkEhvUim0JVunuPmtmOnc8YcPt+GS8u1n2oCVfMRjU4K80Gg8yMgmat7h
j/YgTVpfkS4WFOL2z8qtzz2cXrxVR4j3RhBI/cwvFolCnkiIVD520bfU6Lwebhwq
qS7svB7wUtSIDlLM4UGygXK5SiI8wWh7bWrDJ+WMs0roO+qEN3n1tUXEZuaV1rBb
025fyH28w0GSwwqz8gE4YD5giu40kini7dDw2mlNPTRZwAM1jC6RPF8v5+S4gTkU
2mS8s94Zy6NNHE/6pnZ7Ap+S0KIyZV0ie7ilABLn+4TzQj5bnmndNc2tU3u8vWWs
uG7aJW4WojXyR+GWgc/KWAiB4Fx8WGW4rBb8m5W4SzjDGgh5YmVVddZwaZBzwa1k
DzjEjPoUFE/62IlpBNzMU1xTHV804u3CdSzjdkiF5yJ5vPR3uX/gL7aTjlkylw3n
kIR2unTONqzDkFkzxnj+WVwDxreXBJP5vzABf278i0BBFO2FpcEQA2U6f8AXMeRE
OWIAFfdg7H1OQaFN/1r0sK9LTtPMygnTjuFHYJZnYEutaScEDdKzXbiTVVfOy0rH
Obk8Ick6sYHk3m2IJ++v9+00eU6kCzOSvu6PFV1wihSR8XZiB2l7u8+IdfkJpe1l
pPAN4bXvMb+SiqM3Kr/rmOtlGYfZUT9Y+GKRze7kMThEorOaNj6iU1JN5jqTTdJP
YdHIj/6hzFB3ryr1nxtHfVdFVVklIGMS7wtY0hucXwgfvxdutPJf0g5HBhIlFp3Y
aV39cXPnntypbm6q7AiKpPTakU3YsXnklFvRKDyECoW4/Zp5F470/z3z7lnREc5i
P8lNqhwskNctMuhMnBf20wubV5d10XbE+jlCD53URZ2rBSnrPYDwAJM35rbSeQzt
x/bLtPRE7WHweWVpSzitBd9gpEqXEOqVr2oRkDukS63rLGSI8cvwndihit4tA+a4
lpxuuxpgGWBUqWypsyQszUNjrks0F/PcDfO4ktUdlSSlYksKzks2fEXIr3D+lrqG
IxCtUMnQF4PIqrrF1nsINzZqc/ln3/uFL1pNbgowzCuzl6bdnaPlJojqr3WL5sRj
2qdWiIh3J9pGRns0I0+RzG87SJGzHmsZRhN3Ekcj1zjkXn2hwk1O9MvXi3a/hiJu
hvtANYgpa+fGVIvvUNj1WU4N/89oGztO8nHWs9+mKXi8ScjavIufICNnrT1ca6JJ
Ezan4PVBQi87krTBjSH8TkzGhQmtvDTVvZTne+cVzJM1AmdajCEDJHf81pLvWiZh
I3hcDUlTEAdWl92XukGHN2RslPD290HvBpT7hW9P9nYXLi01m0/mppeDy8VLrjHQ
lP178zrPUXZ3eQb2erC0yOPIa5S0kcXc3uKopYnuLo7/f7lmfkXyj7sEAodIgU15
yqSus3e8GfGyqjdOEu1KslPo6b6RHP3OBkkt8NaVyfm7JDn6vzbC+q0xmjc3DMjF
SKfsVFVHsDIYrkz2SjvJP+5cyQMB67MZzJMqNloY85tVsZWqXQoXlSnuJByrYMFS
hnlVRETWpl6aM9Q7ufii+s2XgPJNlpOa0JnuYtgVTDhb5L3w3Dr3c3GjTV/VoOtD
9ZldExDIy0DR0J/nQvMT0B+hPqB3j4pR9ryuYHPHt5FZcyfiAibJHxvOVsUlFQbo
yqZrjt240jTh37mObAkXZLwt4lQGO0kUj3o6YQvVIwc7O/yAUbwahZQBaAs/g5Qa
v8Znsz+Q4kKX8Tbw945S2LYK5D5kDVDPxbI/ICT/OkM5FJKbtziOaBzveVgbipro
KVPVis4GvhoWsJDTuzwJ3iQi6dRGUjEKJdFJAQ+lj4ddUCOJBsJq9OopVM+dGjKp
jsEZC2dcZcsuhbuD/LMbTbVn5F/9ZTwHsJpHF7V2FU5TuKRKNn2dS/vEJDzMZV6F
rSFwMnpml6f/eBmOo64kyRQrG3YkfpChTz2PDxthhd5gbfzFoRkHF61C5s0v/wx6
sHNhStrnroQXCJvddKOUZ0hqAcAtgdwkGSXnWIG7gM/azIaSm6Nf3QQzo3k23HmL
gzErZS8Xkw/AqdcaqwaxZS01rYU3gsfDFmN53JDCJLg0SLT6Ij2OLOvDUbIlbqSp
UmniII1GRfhtguFAXPwHdnP004qu/c0GpnirAiquP/AVQoxg7ixH076LYnIGt8Sf
0lSgcJbnTwTt6uXi1Oxh8bdBD7kUkpLBy0V3w9BdUV2fEHuKB8owLkxcqOuwGdbw
Cz4Nt0gqAOob99gWs2YMiCJam82g+tIGvjC9U2uKqRCxXGUfoF8C3IZ6aKW1HRx7
g2YtdFYbRd1rc6idFSHASn/qxLTkeFRml5ja5nXXLTkZw9KsgIq+5PDr7KSWM6Hn
Cl9Jh0H8MA6zThxY4qxABeKYI2+LlWNsXoXfnmCIbSf4/H4CZJzZPNHIq3Cabm01
BaZJ15yk8Z9y/QzpiyxdAR96aoWVI+r/F8QoheFh0uKTQbJ1ucScryiho6q1RkGM
2uZV3CknVG2v+ynuJ2LLfNIHm0OYKZU7PAbKnqbsi7t7HPVjKZQcLmNPy00ad+DM
obX+fDEdDN3GZu1qysxL5cyjI3XNyN2l6o79KbnIqYiXrLPnzX9/X9qVMvQJyzub
GEBnAu06ASxNQER9wn0d2mQgRpSSvYGwj4T1NgcrCtCOCjnn4Zo9I+s66WyBYN+Q
ycSU39m3x4QIbd2rWVWvqAy9J137y/8YVBNE8unWVhF4AlUWHjfyDqvP2hKw4xMm
jiUyutV1vAxwcVhTuRvLxSV1m/yldZSC5bUcK8ISjIoWlh9hUHaXh+B3fNdc8KQq
Bm7sy39v537Q0jyOATqe/0Q9aCsh1D1XaR/gEpwvIGkWN8UtYaG/d5PrHvdZElKX
OGSumdHtntXnnQRrmi8MNio6c25jZ80WntYzuRwizM7A+EZoDK89/QbqICKbf5C3
bUmje1rfClL+tHqcKYIzekrAUD0CpwAotjFHcMhwZQ2fDV2EjMuMmKlPOaYfVXkH
8FxIcW2W6rpcTbfLCTEKAcFj8XzlVishmGN4T/UMARRVVGIRhQGOxTrvLXiPQwOt
yY40catbCBySQ70wggJ5mCCWF5sQXVSdWU2gBR15HUMWQU0JzreLXsyAnohMMDfb
0sAknrmrRAziaO/Og3V29slXRQZBXcxcJSyQUvQz0Cx2e6vWzy4cv/fZap1OzvE1
ofVhp1xVqYNyK342KBxXKJr+xETcdqLUTEXW78Q5opUv11pRdX384UEifEGX8I6c
py5/D7AOVJtiOBrCuN2EfgE6AJ5r7PhfREHcMuPsEEPxb+3Q8LSUFngeMqQIXFHH
gKno3yk8rouZ5vd1vE7ecA+CsUJ87n3ON2vloOjPYzMGSpY+fh6WKxDtPr6a/3ry
EP2y8u9H9L1d9JyTzG4kvUIlHGAj+lvMtckpH4KBp2yaiJcX9T+usIxykqiyrnMI
qtcjDHaTqbkKFzJP9PB2EooX5tygOi3VL02XQHmIVe+oWoq/6dAPUr97uzb/bJAg
TfqnpbTs+3KPN56KLLCnDaMMBzt/PyZjtI/gf0XckTW9veUeTg5pCk41jylwJ9aq
5Ciy9p81R9zOZxHdnihAZIn9TLDQF+my1vCZPfwjTTK/bOwF11o96MrGiCAMsqum
bwdDFkBr4kohC/HWX9AYWet3FHxSeZvsLeRj6Z58ZGn3urPbze+xZxO6RloKAxEF
h9+w26pWYG/yQWD4pq6XJnOYkoEgesKtKJNYZV3K6dNFF+FXMBtaGlozJwaesY8K
r3U5Y+P/iLlNho+3bAKE7qvU1QO4y7+eclQ9TCzDviPsWdPImjSR8cl3cSePUSRe
4/bMzhdCzO3Ike/is2Ngs97js2c+QNaleqxShyU3YHnQ3zf1WkQ20JkEUNB+i6ug
GeMeOqJd+K7kNY52dnyrj2JGVZB0zJH37wITCNth4j2rYBJ4QDpq4lgHuj0QdqEC
2fxlhNIpizAUb5w3/X28DmMcul3Ep6NtaioBJaf/L6RubjJvEmjkNTwP3wMebBLh
9Pl4iILcE8Gs16/aFBfiZji0olj9evBALhPZrEZTCuo08OgmWWnDmotFfpZV0LE2
ri5uuBdLFYkB2S4cuyGg8rImzEsYzRDhQo9g1tR78x1uZJgELMuz3IupuF9e4Cz7
ubxj6KNDPkQcqo3lIPY63pJpDutE1cPhjLjLtbKdSi2eUotthk9E6bFFEvSAXl+K
K2lCVs8Vkjyb7eQeBcsSd2kYc1sQwHpx7a3rRF9mKYONgG2opPfJDdzpBSySD6sZ
IMRWcFh5jt9rfYVj6wkgGofP8vPkLvZf7oEYpI22zfFjys7JhMGYUUu2o6+FpH7q
X3XcFWMyNfGgISl1DgU9mhewbbPpbw65upXFKaQWBYKScoNF7zmYIXkDZFgUNa5N
KPRus7uURKHdP8A/3eN6hwoHMsZ4nB9XhUk+vNZP3hu8jN2WSv+SymiiXrt47/Yt
bOcT27Jlu4SgABVcMzYWg0Tr26svmHuMI8lXHSyEFIPBcjw6VsWG0o/Haq8ljPA2
No1+9P1Hp7Xywla0s/l8BHhtpWl/JNg/ZaJ2/IYqVu08gq3jrEp/9A84f+xEiZqi
Ou5NZVIk2jPGZ3tz/xyMggc9m6PG2eLchMd4wZpfKBm9awelWX4OaFOWwpquUQUH
prW292ymR7CTbc972NiTaz55swiMWy/GBmNptt7p2+uCvnK+H8erk5MFqwHvofF/
v8q948imaKAFtaemxzfHP5nBPZ2hsvexuXikvBS3jIPTxqriRfNh9k0rMIlzJbqt
Fsn9fjdPc7TiTCFpLfQm04clck3dRIwTuop7ASXuRxN2bU/Xjz8Ks9TfaxiOmXmj
zK2NxNbPAybJIlOvii7hCMtlWPGo71/Zdq5lqFF8tH33tJaDATgbm1xFdg3nfOCG
X+1STtmuX5CIsHNfgwn6JswoL7figSaf8R7c2Lvd2qS9PYBrubc2b7L6VxDon82a
XI3X05mrcLuPKAfvLW1Bv+N6sNYHXYhSuBJfpomuUP0bvuwxQ5VYV1eHqOMQlzBy
EmNd0Wogb4NImViHoqOi5qjkG01xtku25szVgVyxevNLFhP2HQfu2uHZDKBgqYdy
e0G/L2QYwrCniZLVAFAKaBojlLPzgjZ8B84V9htMNRx7k5umY7IRxSG56BIe3Qsd
1fIIiGTVACvMC5nmN+zPsIinAsdROSerbfIQDdBm/qKhaxaBVfN/NYHPf4gTVAyE
mSldZz+quKnPtGTWV6aKx9vRDvB9Rw0/sSg90RG4PK4C6xVopGtBj4nHAce9kTPx
meyEUmcvM9vy3i7Bh15r9brb436MjWIA91qp7r3Grm6ZeMVCaPcVBrU+T80Bgxmo
pDpmp6TKUs5yCLOYRMf4lYGT571qUOuA65lEcypkJW5YcGtec8Ecrxz5lJ1ax0ia
dJrbG4iPRoBTEFCB6dlP6hndfoRx7tVQYKJ45kjgbyhNieLarjncBAPPcWdnrZEr
A5EvpLXY1ZZHzawOZlsrnx3GdCk3X9OpWcHjhKUhCkXg+bb45TF9XWLw0wh3uccJ
ti4BbAgwVcn5SEA8m0yVpGCLRcFagCyDvEPZ1UqpDftrDajYPHiog3VzsRPjt1zr
VXfCfdj3C+0oOVyfGrgZsw5zjtr2l8Xklk9Pa6KW1O4XuK9UbvKx4yfqB90gvn7F
H79dW4lDm4UpfAJFPhhmJY/JrO+qya5XmxwstXGHHfUMvcpqY7dcB9Qzn+VOFVNQ
L/pG2bw4JJYshCLV7Gb/2r9IzVGmOa17hqk/Dck4CRB8+TadsCOyNOGVZmHZ2S05
VTHilUeeDIAm7gwvu9M8Ool82ItOOPRSgZk2MqmWBW6kCoR1v9ar4nj/XOch/Cez
XqUn9jfKOhkba6079BHZw377P74d5Ue8lQBbhSfg0LA+pZmGFunG7Jw+yKjQBUCW
OeKvULd4g0NqzeT6jy5ZYcLM3rIpEuuVPM3gQoyMH3vqd5zfhMtjzY8cymt1NJyg
FyT/S0uZgexFWal40bfvuDX5hqwtxy+2UCBgf4vg3RSE3wR+nkiMI0aPHniE5Nz4
D/Koh6rYRQbKJhzl++Nt0bps4OVcUBALRS0lHD2acL87fn/FKjCu4K2yrnBYi0B/
+/HrCbSyX3f5x+8LvgpCOiDT2XM2mqo4t1ioBJ0s4fsGxNyV6Yjd6Hl/Ew0iQ55V
WimNUn3g8DkbtMJFeSCcMungL17s+9s/Uz0eoCCIPbFdZamyLpYMtTB0wFmi7VeO
HRsaKhRHC/EeaczxEierFQTZ+KOJtTr/B06pYipPc26gY8jLsFWtUp/fUmKkw6Z/
51aCCiI/JIDoNkJw5tRh7RTIkiQ3tOcZQchQqjbZVBRFClPtk+A681Ip2Ab7wyLh
QpsSdVcfoujzKuBcgSCtG2plVCTQWJYe5cAdyY5DJDHVmlEJvki9aLdw2JXihwBB
eyg5gtgQPte5ML6BbYx/+xwQhl+rTkw/+q79yehf9VcFZULHT2gMnJvBTIqRT0zA
6RsRqLWz25ViEs+nBDJ6OedVin7REuCM/r79lYRGlLfUdU8AjPCgwteG7zd+K28N
BSs7A8KXLUuGs9ibHuoPjT3WtJAiYlapNpv1qvwIRN7adFNTPoDZihV43pcJRYNO
KhQ4amENYdchivtzw3k01x/3xIQzrtGT662MTxpp8Mq45y4oG/9DNA9qGeZdkayC
W0X3d5k0GyG9TvXVkbvRu6dg+yy5wiSA1apoNmn+XxTT4EqdHxulNtTMW5rpaIq5
GK+Mld/+bQbvkcOfxFbkHMMP3Z2Nw6ekAu/TC/+WgVFZO4T7+t8lXo4W33DInwYm
DFVwJjQolWldAa0qbf/DbkT0WfttEejUMXPhFIpWed/Nv4DwQNjMq9YYqQWORruL
6vvNU25aoFgPSEwbjYBihbYPaFKaF8NFuc3eKXdYYapkWVSksqmSpkt2k5Dw1UhG
ElJ00sC2t/777fpW71StQvuPkyweCL8PwOFRKcj7P7DrBo8dAVWRAlgjePArs228
T/bkLqP88APwBG04VekvNmwTqlnyCARyMqHZphN4/QOiPv+VFMbWynxQ4siKbOub
d4VpGuZN1imf6Dz8hCrqZb+sRL7xsBfO9IKQk43uFHudUzJ/Y2zNsRlo/+A3SMBw
Yj5PjwaVAKgt+jhaVxnYQeMWZh8tK76XU2Gb74MddmYHXLBBcIpsnx+iWr5VqgOO
PhIUt+N94z1Apzpq+x2kExBD8vVXLrzF9se3Bq++U4YmBozIfZClDCIM9E6ktmeK
l2nFzTSEkl3FepvaRUPJxlBNeMBuSb4xqr9llh5vOyFcgogtghHsattiMAwOHI9c
JsBUbw0myD/mDBpGWHUnxSU2UDGXxY/psWN9uI+PASvRAxxZ59SDjoEb9JG59u/F
UsLM+eiufvVUvPpT73mUTA7B0mFfyx9+R+Awt4DP/UDwZZ0worSwh1HSQEHuZYHd
O/m1fzmpwSUL2+YEGPdltFV2k8SVkU1POkEtI8y5SLDqPyhed4gaBTaww5kdjyNu
a7M+5PcwqGSnUcbX/W7fwCS/bvhABB7Ea8sFMRqLIU0cOKsDesEe4L0Ni/8VXCsG
kDuQhUlElpo4lHbEUGFKkZSd/U6JS1grCcIgeLMsAR6RuopPViYF6QtwApbeGrwl
v3yi5nohVnF1dCVTPWyPmnuFNmAp9qQR3L1CGsk4faR7qO0EMD57MYOztFa21ZDg
T9jE3sZ8OFJcZsMGI5R9GBvrrtsMszu4eY5gVzNLAbd+LWJeQdvxSPm7+RzM5mxn
toqbKXgLZLzRs8y9ZUYtsWoGzytxUXjSBWAcHMuoQAPKgue2EMLRc5UzwfmpTEIR
sS+daw9Ofq4IJ8cc4M1Ue0lsnkg3TwzOlTiiCPfBGaHFMZe/TLKA4CSZipJUlRDk
K1IqxXLWMXIqyXst7GdM7sQcMQzmmSxB5NS50KMFX5fMsjy/eRy9AwhuJJiRMU2x
oonXugDeMxQD4MIBmSSBodvDOueps4Pz9YbLrZ/PvRGIQKhFu71NvdLALlCNakmM
hpxoVa3x9nQHHf0zl/OKmFOOBFGySNZG/L0wbm8pe/BUpLdfUT0Vox4hmdtbYBhm
FjDmvpArKRAVrhcOaxHJcFLSj3HTY6Iy/MPxRiPlw5lI8/JtSDv7SerIvJeIUTWN
btoWVv8FgM6hEJ15FOCxtCYihOxiNlspq7GRoKBQeNOJpuWZ4hom0TnmhJb+Fkcq
q/GBYLfsh9hwUfe6PDEccTIYvFb1KxAi8a/1o5bUqWvT4gEEPbp5hhd3M8LwnOIp
LUZbgztv0r99w1lQwlEfKtHuizIf3LskOvVFDs6ziF4Kt0WJgj9N7DUvHvOOzGYf
2n/cXQagrKGQe6F7PxLsgUgUDdknZAgGay6SXJwUhPKf3wUQqCT/rAvWcO3teh+j
TI6EJbaFAr6ApQGWHaMgukyIv+vKrUe2xSVEMKuCkXcMMBC3dMEScPPLC8Qt8YEh
6P9z4KSMRgDsXJF5mvV53IJplK26dmUF7p5QId7BN2nuVmPZ47V/Z/sEe12fapKM
ZWG6UEEvZhlKOx1SqfwcKtdh5IJe2OdgWoZu2jkupRZjzUMyH5HnLiKsNDcscQSW
49QbUWHWuAp+29xbKBsLNl5AFrOMG40am/vvS1a/w38WvsQtHfsXTrExup+VHOXS
ibOlFvatk9xJm/yKeHkpfJ9O7ry79ZFwsCCg7/AbOOwBSqH15XghX0/CuF4zX+Tm
Rf7sn5WvFVS/tYiQ+jWkWdJ7S6L2bb1CoX8rgEsFrZhrPFl1O5m7FvbmZCeWU/mo
Kx/4H1ozd3SNOd2R/n2dEWo3TRsr4v0ETb29PoLd7f6MLw5O1H49Oyn7jyM0SXDj
0Vrtsf0gOo/wHUGTRUG+iOlEu7F1MtZVcOJboWGp+EXc+h4hlouQn3Jm1gyvo0sj
J20d5+NTqIsA03kn1ijkVO6ynTKc/CnX1KXHWmQpmJK0NqcjcCyEnSXtGwSh72d5
qIe3LS9Dy7+tX1OeBTmEIwmBMDakE6J6SyKLFnCZkTa4PjvxwpvzdIQ74nZ3uE/+
mJYFaiyTnsQ3foNPTMAoKw6AzN9tMXLUUsbCj5J+sNFdp3Do81KrFjX5yrbxxHmb
+fFimSDWC9yh60oU26SSHyvoKKB74OnMe9merj3mTVi/P66/rfp1vyySdtp4glnt
Qkg1iWL8XomWaSiNieVn7MuSofTj6K1JyMZWV7z92RoaqZpAa4if87aRCA/HUd4J
0j9Nq0+LkQAVn4at7EM/zj5CinA7UukrVn8TBsiDfLfT7h3663I735WJQ3hsmMj5
6Fro86s3PePOzZJt3hAHpeEvu0mUTcT2PknVJApkPB6wI/2d9RO9YtQtnfC2/IMt
SaYY/pTlJ76T2VYKPPIsGkxp5tKyFUd3vIGv2nFNTyUmx/dT6YUVf9S10Q9Airhi
owlvK8v+EFm8SZ5KdNL6hvKrnWftyagPkOrSB/aACEv1/A2dr6v49o87lqZUplcX
ZHajh65KhzIMdq2lPNlK4njSV5G47ihKiZfw6kaEw6dUU5atqrGLi8b0S4JLhvVr
ndsULsyk/iNNTY/3yh3cfjlM4OiBI0mzcEmKugOQioQksC8KSPCEuVclXlWiTS1F
Wzd/z+c2Rrlm/+igZnZd//ICtxyv8OSgxpxDIsoozXXHgIFjebiv6CuIp2X/MA44
hV6Ju2XZbRfvklLRUnGROMtuhn205lsNAcvNy1QvSfV0V3NrQrFdiTHcB8kU+CmX
atJV09jpC+lTewrfuDiedsMUSmzYArUi3EI3WNvubrpgVl9ivuzNFNkjOAoRMXnF
SrrGJmn6qgxktauebkSNXkCdBshZyfuRnT+6oQbAOI6FdgLz09bvgmXM0T5W/JEU
eM0E2a624bNkWUy2zBOw+mW2HDzQSTMjsg1A1DZ06kZK7jNzZFJGV1huiA+O5jFb
GRvPtoefDD12ryXIYPTdn8Xr16qcqrySsBpZgY+aYtZtcXMf5HP7xd/dY9rBGWJf
RoGMfiBgotkTvy8YbEBqSUjlluSwm7wZSDSD3lFvUw4+dOKNCHUoEKfa1wJ98o1b
wOfUvj4LpGmRWzBmoRN+fCVK0wxF4MzjrpxYS/HSD7BAqGqRunNDoZjGH/jFQL81
LwiygsnXPSXfy33q3jbhX/yQPBjBe2QrlFTEVzoX4c/akTigK43qKw/OcxF+Lgkh
afVaBjN3XR5ezgZbGr1yPlMY1gXr7p5XvfoZdZMeERGGUEKWgjRAqsp4eh7ZfKF8
HmGBXM9UtTN80jE1kzjYJaI4O1x0pZWKECxGRr3ikxdnGojc6zIcyaKy2Vza3T9a
0binJJsT5DTXJtyw5GInFkgX41w5ipwaRoB6mqmxWl2/eFRo0SetCHKcNttxw3rD
iEBFwSReZ4DLx2b06OUJqCkxeN1Tas9XeNyR61qOZ4LWiJmOy85gAPoPjY2/mU7j
Y4gXUth9gCVDqnGT8K4h6fl0tfpORDiKTmbSzb4jv0tuSHeMLdn+Nay7diTDIJxK
zGLHi2fefoHMu4JIo93+xWpHCZJmjCOLS7DlFkimuyPryxwmOXF2qII0U6YZ0h33
/zbLnWgbscAeHnEGJFO0VOLr1f27KBGJ9rs+xnEmSL1gUki1wm/iiLLkGDOn7+SP
2tz128Ms0R0G4wEVVFhMVHDNoi5JpI8wxRP6BS2VI0DeRDAQCy6D/uYtd7vnXJJX
aCNc+QoLPOXJipiLLA99U+4GX8kdN4Q1/7r+WTM3dqyGZniOVhUBckEmErjBJmPj
g9yB+7sxR1OXa3lLpQwkdaDx05kiwSy6F7w5QS6eT3JWI4xX8x0em8f62toW8K12
DSnXEdRzKuHYC/mHUT0t/zxX0XqwKsOxz1QtWsV7W0qpzWp29iGbVvVMzWUSMHSn
CLrZq8ooYqh7Mx16g47ngUYTuThhG/U8BofD061dGvj/afxaqb/u7tHwQOHSN0lb
Y6rzq0ioTDTn7sd0IRbvCPLTnEAsU+oXRpJu4ND6KcBYVbmnj4Wve8E21y8ezMLX
5k8fBkTAR0MStiAxC9AxpjyeQvrnr6TvIRQTeztrkOnnYYq1blRs2NJ9UBVbiF+1
/ovXuCgDx/o0etAz3DEMGNCzvbpuXXhnOHH9VW/WGBStY6cv+FUHWPAW3/JmIisZ
llrJieMBNxrNeSVpRFxvCjFQHsXCLaKPrZMg6fNCfkSJtOE0VL3JP7/z/XzHqZK0
2qZQ1s2jhXrAhIHkx3/DYG49xRs7ESDCN8BdFMeVSCpAKAPpAKmFB/6/lPyIlFeY
MOA9756WFNwJLdcM9pxRTmFHxvNTjUpxX9yuPT6/mw3K48WsAAuVoHqiqeZpKjef
PicG+M4f+qK6qYMMcP3S7gI5lCytErTUWsMiGth02odbfnfpRfz333eRDolJwMjR
FzvxlnpEvyMCH13k7fKpKSMBcmdsrqi1FCLa9DhDes28TzUQixb6Dy7jsLm9wiwF
eVFqTtpxcuW2vl10P3swhR4aULfDx2A9aBWmrVvBQtLmqVGRLpzdduIKn48FuZBD
/SJY+MKCyUGulbm/umnodVJ1Nomvjru/VcvkIPZUAkSWodB1D5L4HArL4Qt40We5
omjUZ7OhOYmwmOZbZmnnGXxKQqrO6nZXl5LsSbSEE8/4j4y1BXD6O5aZBHWRxbBm
LrTxy/VrQ+hSaXmdXlHn4P/V6iq2qVjZudxN2K2Gm6Xo6tOwSPickMZovBmxSvyZ
HX4Q7rGGaIeQrcMiHtDfTJBHbLBnr4OGBL/b9gLwAE0YZCO7iDY/xCfN9HokIwH1
HSg1HYGPt/tuObs5rNmoEZL3Bd2a9GQcqF/ZkINDknKUjWu7y/1nyuv5hOldoG94
fgETa4CrN/oaR17v8kp+b4W06jOV5T0F2dXA/S0o40whrvatmf3cTRejgA3fGpEV
eFFMutV0TM22PHyMADKuC9IFCV3499oAiq013wKTPrs17ZHYv2U/o3UdEPxnFkHo
bIpeej5PONy8iG6GznR43us2u7LJy5ysYarNMiSWtS7KM//SwXVxEsQlogYPrCZh
jimWBvhp6WwvWSsPXoJzheP0wxA4cDnfN+6J6CJ74/zjYOa/HLQ6WtYjanHPJo5a
`pragma protect end_protected
