// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:16 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ImKtP5LTLog7N+eg54bjQgjSbUK9Ps7+zn+/pGOCw9jD2IaXTkkmF+BWtXdA+skL
SKC2si03+tJqjU1spR0QWhaewxCUXNHKxKAYtR52I2whFsv8+Oj580H4AW8276oS
LpBsAn3ujDANgjCV2XiFqvQq6WePFe62wHjcMCe/YdU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29744)
MGWHVRFYihY5B0WUgPxMvSzZSppBfuX+/pRixMrFM/fLra4VB2V82eEEShLPOZnH
AazcSqcILam1OFITEhcU8T2SHn/NLNVn+ChP4DUN6zXYP26U+XoypF+GaJkUT8rc
Ifp9X4ktcHLHM10TNe7NEOsp6eYgMhWOkdbDQ/ij+XhgiTBQ764P8BjIyHEOIgiQ
+JtDIs8csHv3fVujLVKqRb/Paq1HI8tmLTTBdgAeOA8AtDa/vHtAWT55QwYqAIQb
IJR4NLt45w47yeUnW/9NhXHEUfbvmvfKgW3+qqay8VEEgLVKwzp2zg0CYI5+017b
Zkt6GsPzMkbO1UO9Ru3VFYj0xbGjNWtL6opwIvN3v00C/SwK4FzyFRVR+p2vOede
KqEX9m9CZ0A9P5fsFiLfUqZE2eIyewfgNwHsOpuhebxz/GGRIFP/O3yrbosw12oS
Uy9qsySN+ftpr470TfF9iXdTp10z3n3gAZERyL45U/Q23CJxc27zR71W0NhMHRSl
qhLWIC+ADv5CLR+iKblxE4D2TDxmA8rvAA4jNnGEAWYo9rdlXFuiYAluhzU4mLA9
tFyaz7MpYOFIzWgvCjXehzgjTFwhBgAZ7Mwn/oBuqSN6eSp0ElxjefQNMvRWm3i+
ydJ6oyne6K/LF76wWhLqwJmrvkHj/A1WjCYElYa5uCbQDBy3NVg3uiY1MaYYbXhp
NcNbdMUtkr1BuxxUwuh1x+6QlKpIkzNkdi9iiX76E1sby8ADfXUCzi5NZup70TLd
vqOVvq8cQaTBOvqbityRPHkeBy0mZG33ljDIh3LdyPWuI1KSumAE8VEVM5I9khIy
aBYPgecfTxsqzrS8BLgFARNnosaE658UB5UlCgTFU7/8EUsDJoCmHWG7P2gpia1L
PqIQkw5Npkucnaac83XWlNVaGQTw5ZmGFq0w7SV5CSiUIYdC/fBZ4LakPqeXzTfS
8yr5O3/yF9CogIMNJ8mvlY9faYDvVqWm1cpzVuoBK4w4RrqcoPYQlXtn/x87MgMh
DMGfZaFQ0csbxXr8942SXyrL/jSLEQy0+a2bQQR3Jkl1PN/OhgMvO/ipEVjlYH78
n1hYsFEdgVpjMWvKLL+CKvVjVMgm75tUk+j0myl5oSF9ctP/pWnsDZVj6hCmYPAA
WxQIjvD9gmbzOCoN0jEMqT7oH8GepfXk35/AWg9KUmR68yOXxIyLqHgWnrHbc82k
2USTl3FwrlX8yK7O6JsYmzUpHvJX6Th2GeAcQX9JT5wXaJduA1GPITAHsEH9wPMa
FtcRGw4c5E/OKHXsPTbAq0q4tplo8EQHuI3EXM6eSQzFxh+QKWCRsWT9JZIE3bzb
jKom38q5DIOSNBmOfsYJvtS6G4iT2SQzdckrURVggMnq53Jh0vb1ecNlB/20bHHE
TLJ1LdTwGUoIUFqYjRiYCFYt/yxxTewf9mh0Er2H96391yHMJ9VBGJsEKNtThJJj
q38oHRnxFG/DY+hSI6SGdPa/os1PrPViiwxcTX3hhvN5Jc0DlsAeO/1iHL6muPGR
iL1OG4bgoZYJvGDPR2lIRyB/G30cqmbTuHwqRD5d6piUQaZTY5seekKB00RXwUAs
wBgfFRTpvkQ2l1LABseiw0MQQeH2a+bJzeiryNn/0v9NG0/sXtv2ERFZ4il/jPqo
Y/qZ//wn0dRpm7elmoqGPXq8AIMIHAvSnTjVi+EJnwgxxwYSzMnrkdBZX4iOUS8b
OMgf3LsYiJG6hVU582dq724fW6V+B4UsTOj1HQpJEhWJr3w3/e2V/Bigu5sqZyfM
s5FokSWyUTTPoRJZqSpprK5Qj+XcWC62AY3QWTTTkHVnp/D/X0PKN1KPBaEzK2xi
J+lI1k4fiM4eD7ece/QZAWNd6Jm7gzWk3Xjju0UL9Pl7sgWqf28o/PAv3R9rxLLY
lme5BI0+3UWDg7aP4PcSDq9YZN2BvVjlDl28WCtmmpxdIbZ4I45j78S6d9X0ejor
EdZqI/MFVYMk2pHmitvkAPZ61OQmOMhzs1BrBheFDSgDO4oUjaYQ4eWABBVjC9dl
0069ALiCtR1naqy2GFvKrn3cyz9sM58z5x3Fdp6gXwFHE4mcJynqHbDkdZVxM5WW
Gs3JH/Q4lf6drDLXh0YP4iEtk8xzE6zysRYmolHSZRb6fN7GZ6lziJT2vEC4YP5m
xLN+hG7YYjpVZ01KFnFZPl69IZEyLV7Zvl5Qw9mFJdOeoJ9vdCpL9FCjF2tOXHMn
ioW6UgtCTWKPZyBXUIkRDruRj2RxB4A94MGNoK2BxlHJe7l1Jtgas53aDvM+67+8
bcL4omB33qFCXDSbZzSm5y+UMs2+ncrUZugy51Ex/SPjvN2Wrb8dz9gCKfl0Byek
KSdRS0ZM9TCtJGlNaqREMZZEf35USA3AX6LjdZVIjEDpNPK0JnYLA4Rz8hXQufou
+OFb1ozhaXUlxUi9xRIuHTSG1G9pOyVqlbT9xs645tSZl5wKfKbf98WsRXkEe3zh
6E/Uff08+AvhojQ9o2q+JWh6okS5Yhy2RjImM7CheKcOqItsm6az/ZFPpIWN9X/p
QnSlzVZzh7it8ArKaaCAnvvNzijZSTsF9VHM9GoRJZVd39ts2DI+Pkn0TwlHdZXw
kgJrfdahERJKVXLwQXCKRPdwz55IkSk4u9g2gVFlGFT7ryoKAwd/4HGmy9YAjqGP
FlY2voKD/Es+hM9jm1BzjbSkwV96kKC/eETqP5bO5gSmGXzBY7fjJ899bofT49oh
8/lAZkSqFbSsmIswt38OK7NZ3ylaSwbug1Pt6k0VmpFWdUNOrEEGgdF7TPTN1Vf2
HAaOqPzvmHG2/vbw+XyBxtrB+Y9vBh4Kq13Uw89pTN1MtiaLaYRBspXngscTldOL
qBbxuA6W8m7eASjKsXzDfsi1go7d8eF+KFf5jQ9ZLDR/ErrE0jpl4zS39u4QV1SG
n684NO/QH4YV7sPKCfOjJNVBsIrSTZtFC0BhXPp5yR73QT5sHY0/cVx32/3e0slo
JDhf5Noc18LA5fcqYYxVkbPMdZeB7SL6F5aTn69Cg68nkuzEou/QYh5pK/UWBwd+
KTeU+hye9rrMnUk+IceYb4YkV5k5gIbA/TNjvHtX1qrGqweDZz7d6oL5u0CroPfo
1xtlrxZUPa2PICYUxIEJikZbieUtMKx3zrSxsuz+kbKjcdn5mEpCyXeATMACpH+p
+OI+oey8g4WHP9+yzUh9H5Vn3YcfDLlOh7OTKDSbsb4/icXfMnFTFx0e+fm14zW9
wMg/r+2o3oToCyMqA4ANDn8yXtVlmpwFYVotORL1nXCrDCDM5UbnKi5gAozb0j94
b/wW46zjygJ8yT7RzD6RBHgRDKndTy/+fNJHIIazXlwPvvB8lvm7EyhhgDnTQgm8
iINUSTSoQ6TqE3ICMr00zgUxERDNrwnwnwTj8ujxONZ6V1R/Qy3B8t9c/yBOab/P
QEvdeXqdYlzRvXghmXZCc0nX0KsN2vUEEGLyMK9XNByMQ7Gexs4+y3/aLXdEZD8C
NUeVauhz7OuTDdsMIXFG31mfxJD/sTaB2z8JazqAVIIAyLkTLkPm3LPoEmZDPqp+
uTIM9RcHLV2A+uswIotLqS5GJ780tF/Wv+Cq8mfqqU91YpImMO40Thv+hNaNuJEV
ij/BoaJHiRRrXQ20zT8QQSMS7T1DOeFnXo7RlMyz4uxnSz9dY37eX/7sET6/sapK
Mc+wPN1R3AYImoTpqjpUj9a2dTmtO2eCX4Vmg1/EI/nCAWPGFbbokV0Wcvix3GVQ
RjxQWhXtwO+au6C+/4SunIZDSRTGQW1o9yFHa7+v+VCC2GTFU5m3dA+uARCg79Jn
j94lil2/FRiAmTKz0uLk2RGN3+4qgBuzPBnlJt7ZY7vJfoKfqSPPd/45fcB4bCtF
TK7/ZyN5/EHZV05jn+b8lnHwOsKPfW1DdOwkmsm1zCrGVdDiur9NbSsy3Ru2ESto
PL4EcglJBPH46hda0dLlLCEzpDAtfvddzAKR0fTDpMGlzJGobU4WBy5tGlAQ1Z1F
pLobCjfI3m3q2oMpdyFT62XAaj8XDo2SJm27Qa8HBf26xiij6edfGeeM6bFD6xsq
vjgucIYwQ6te+lALqcKTEeT0CPBxCulfBvbx3r55YNbW2m4zMyX8guveoU6AvBL9
wEuf2/SHCHamzJX+6pJalx7oRGD0Z5lEZ0VEPer8dvLcxYBESBG4wMKAnamV0+6G
s+crr222I/KSlvUaNz6to8O9VFiCXQTagEVX9OZg7oL3tV2AhjLGboiSOTfUjOF2
WL+YaytseuEwXNZ+sTSR5Ziat5UiPFtzXkQgGTUMOi8OKclh2kK3iuP8Ujuny+Hw
et2LF7+dQQe0KA3Ojub63oEnLVqExz0ftgjsrKKtddl6xp5PWXvJo945ByEu6qXO
v7DDhcW6/4mAaECjdUdaNDKsri3G3GfWM3DhVy9Tm+6pwUB5TcWPm/afN5VigFDG
v86Oqdzssjl0P4pOj1bQzaldqgKG29K9Ts/Swa3n9ZyXOHyFh2GmWy+gEcb59DIj
Ttousy5AIPi4shJrTyPyBOJQyS41yx7xBGqJJNjZzNiZMQiviUEz9G82osrJezVg
NWcRgGG2HFWZfHIv9kMPCByEoE6rORAwMdflUpUeCrgrfcT0ra1kafD3X30gu51t
iPIU7u0aZWfQsGrsHSnIOFyULakDF+wjbPfLX/qOuRTAVcj/yxwtfFL1cYw3RbUl
/1rMUt0NiZqELkGJC4b3omo+cFO4NKdJwCq8IYmDauOr/tITphrLUGb0nXOiCkAI
kZtVd/sUX0RqCCFykv0UzWGypBMpRfdx7XmMkGbGH4x5NTf9/ICgWRL5qv5FXbmR
KVJiSkWIP1uLjKJ0dwOA6hLbq0pketZZyChKNctoT52VMyHd2sQSTJWdnYifYacQ
u9+1B82mwTr2227PwJqQUXIJpl5G681AvZJGrUhbMsemjYZyBtBbja4kSi8JKCHP
V5UlF2vwOCUJkQ6K11erLUEO7y6nQfOPpER7zpSvV6DEw4V3fnM5rECuWNPTopr7
51dxEJINbanKzCG2VSs92EqhfoTZyCEkvYKL5tItUn97Ck8en6kRR4nvegAU4hMc
qhM0eBQs9wRtaJyuumliggaVtXMlB6AuVEBC9Xy/WjhTQ2Cp4Gqb23yoxutKfTWv
cDSp3cBznbhVshRrbddEgYK4+sWtOkI+TGigw1g8lrmNmidVdTblnxmVzwHX1CJu
7Oh4MVAfrAAjBV5aIEr9y9cJAW0WiSzBeZFSNPu6QSV6++PVmdyEi8lZJMlPOfYg
/UkEHkO5iv8CEjtHVS4+pMWAC6iTQnrd/hg4M2/6FjWXrs0PfcmK0msfhciqFBNd
iYZ23PLAsZKhgStX6f+OCOyEg9aTE4/ufvpzMcket+yHY1x0X6ia1saQYq4PXCyK
kJkwuv4rG2li7vC7Kuk/OrjMHwzndpVIqr65WgTRq2ey7kGjsNjpMJa6oLnFGxmH
BJITEw9zVAz9kem+k2O6C68mTskkXKBOzvMcRrCQ5t+ITviNsq24xu8F/uCJooEp
RvqzJdhHTDu7WBAKM21VwazUjnyhKGZp/fUuJ5x9Rnu15wJuwK90yoaOanyHXfIe
4YrPwxOLz8yOc+9A2iX4swAcV3J45tyPvb38Vg6sS6okFqz9he78JhUQrENRdYmt
ispwMZMhEL2frHNeQVztXkEp7I1Mqrew68UhXuPe0889jz/4QQOG8CwEFhRZFxm8
wv7zYbNuYxtBnXKWYnxVz3JXwpd+Sd3stYLNwCXImebBmprEkAhtpojX3qLDD2Me
OF7aaJjq8PeKbnBbGZrvmR/Q4YKayrkPzaT9taKV6IS4OL8l+A87gNPCgQ4i9V8P
IfnwcrCPM1NyELCaRUZ4e+kFBJ+lLHgtsEc7UKs9ne2B1AGhMBjRGBB8JF1h+39q
AYKqpCVQRFBzqp8RqkdIFG0DuGVHVfKIRb0zGasYw1f0pWFDrc+A+R/vGdQjxk4m
5w3k6fYkfhMMnnTXevJO1CP81qvwQUOeDU8/+Aj54f10QZfgXAbzArTrY5Lr/kOv
2h0YEtaTKpblQYlha7aHSymTCJe9dv0TL4CUYQKUlDKKyA5a0++hl1Us7NSLtKuZ
1p9d1z2kbJkIuDmAZHFI1gub28F2ELiiUU8+vVS6rZLRn8o8Uupjitris4v0Gi7L
YTWzDDqJP5Ri5b0m62gju3STO1aiuu+GAuiphF1rqZZHBvSIq9dZgcaevP7zhxpI
1hO3T9xKZtz9Sq/Ea1G2MvfDKRsTQVu7IvvnE6RSpjHy6dVa8a0nXUrdXVe9nNjc
EOxy7So4GPNMLAQk2sM0r6utSv5gqAtOCtS0C9lqmu00YP+WSI70zqh51cCXdMdz
jWHyu4+IwOoehfkU+cuOs2dSnm0vWRjRWlC1yfa/UCz7IstpDwmolkyWYDsMWTfW
W7dTWEaHishlm6OsyYoVcHOQJuFm/83kgJDIoX7br7tdshRwVgK/8dRH1MQJynpW
05bCDpHXQy8xX5eURx8wp0ayzD09yBFdGAwUGJLYplzT0YKtUnyHgiw2Sol01IPp
9bk9CsUPeZVjyl2joa56/RNdsO/LCD4sy09+AMIuIzpv34yIHwqtnDEs95a9Db9F
XHiyLzslVJqnwBKiobYTWJVAMaUobpfyKk1DR2bO5yrWkIAf9dQ1/OW2Vdv3Uitn
HfjNEjtor2h0eFG4uUo9XTUxl+AEG++J4Pcngr2OTQVJvE4tOrmVr1pGtz8o37yS
v3PzrbSOubf1q3rBfSjIk5uVLzjw0ni0QVlv3q7qUT/xpMvvF09yTTrnq0q0insG
62sCoTlm6xiz2Kii//hIo+Kv4jXlUW4X6nvi68HB6tul2w4VbexBnyCoCEVIZn+h
Iard4Ad4bLy5Fpy54u99+qOxVZ9+280HVr7KLErM9ZiprpnkPSg5pidd1f4kdbCr
wGAmmyOVb3TDkxNn/sNx3T2gEmZrHdfYtaNrnXjovfI6LEGcoPySf4M13U0RdmWe
BlMnIuE0obzVdxVfUt9WfkP3/cqxkPnzKco7lvCXu9QkBa9q+8z4ss3uMvEKHuIb
kmmFFaVmWSdOIpShvr+3ZCFB15LS3aF20QFliBCJ/9OOdxyePVxShSSX9hUW5uiB
mEInWCkmR3kBZVBgwfL3vS6J3pZlTK4i5S6Ll84mM5KoXl52tvlzbZyEr89miK0A
2hN4mBrE8V0Uz7K1ALEHZQWFbTdd11tpD2kXfYYEqOgOaXYWM161+sj3lW8AKpA2
YhiZIz8cHICy/raSz2TeAEEcnKUhYopXtCLv/GCC8A76Os2a1Xfbwww+PiUP0Es/
NZU4ACnUU18m+luIb1PvRYEPjarSFiYsSfA8nYfk4HWFw889ojOXDukC3bVpMxWi
EYZTkCBYCY6d922vvjIomjxrhQThXhGJ4R9fGI7RSEdzTrZJXhyjrUAAFLvzb8CE
YTc+Dxysz8tKxeQRAlxPApyjbTMa1l/IPxMhOpZ6uuddCXNQqdCGmW/o7T3zwVtz
/QhPm/ehjmpl6G10EpvVXwopTVzcp5hb7A+qe/adn0q+afX4+2fO0EDhH8UfAOyr
GRwrnV8tVqBJ3IIEPpMQFaWOl86mSXtqWUeGPNULDVmX8Y3ldeRvjY6kR5oaj5l3
Ews9Txniv/LAzMknBE3RkjkBMRACofEWfW58yBPIqrqufNsqkcL6bzkCd0DkZEkB
a+LtTEaGgkeKDet50G/WR2jMdwdHgEI2Ya/CoW6zbY6CDMNWDWMv/GwcvZddnlVX
xFE3Y1GTMAoFGEbJ7qlRzD2BphVXG/bcYYyrKUK1EzTREQNP5ZmYY8bq3cwfNo7z
txHTSv0xPXDdnT63h4O5xUmQmp2cxCxe1LB+vjevpCLl1EmHnCeSfIG278gVM1FD
6dq7NIpS2VFwV9hhcnLyI0Lv4Se9HsHtcYEIS0Vl6sEJ0WxI6QnB0/cpkZHnE9lA
F9yrbXu4pWLb1Pckd3fMSPAgS5cWodPJWN2tVqyYmZ2QU4853jqyuoHj3lUaSCwK
pRiXM+yUnGHtbwAVpxsvWg02uggOHvqrNu8uO86WAvxLGuZSxgXMbxHbUBW8fA82
juIKtkmU0/vYUV48Revw3xhC5Td75pvSmE60PmKE0oCxWHzIqsOD4yvZVAKyBpEd
z6v3LJP8HYmYcYUTg3U3qyEUpUZUAQ1zMaDL6ZALvS89xDWCDK4yjyhacF1lj39L
1QbUwBfa2otS4TPVw57DGbhwIXQghdQb33Y0j6KAFyFodoaQHkwCfOs7cg/tprAQ
6suzuPqiP1YBuYJ8fpeBKlnR/F+hTnlEW4HSYn+mXm7hQV3AuHPh7xJXPE+hSa+0
7BFSk3inzysqpIxCnADJEns8DzJuoMDPSKsb98I4QfWQjv4rCJ/cMLyccmDSwT+O
nKoDAW2w3N7sqF+Or+PMUHEs2MW5Bufm87YSyTW9GvGsuiRzrF1uNff/VQJ+N9/B
kHCE0rdpq3g+Eb52BnQazPGmyX4mrNBwZ/Q1cG4TgoGjpaO5Pg/KKvPxX6SoD7xl
UaUjw7K2s1JBVcwTAqSVPkMkYkj2rEkxjuF0EOEMA7LWh4nwtDkqdzWFrtZGCKuh
hhHi6LIsLPT+/+0A2U1GOLTAxJs40G+Q4+ys3ghbHx2fJBpvoTvTU2OuJ4T44VjY
iy+uVs3b5DxRWLQPPX0HVBuQcIzizGV8eY7bAvSMHFPuL4cAOXSlkaSjFesdHwZB
6fLajSKXO0T3Xm9vZHaWNeJsyeICFLq1MHx8VsSjSZiOgRupX4s0SA/+qAFtGZaP
sCd2u6ciDd2d2fV2fwydM7mY+FAqBeekUmpt66h4GJ/KTmXQTnBm0L1cYUmxEqWy
3Ri22xcGwWv9McnAbqJMY6bjrbnyjGAVeLexv8JjEXXJMd3CidOwbjdqguN1+TZ5
9jbsRq/daSEFXwSgCdMoHdeNq+wc12y0UI8c+MgSu2ybIWUajpOZF4gdXWAP7LzR
V6uCCJYpWLrczr1GuMsip5UOLf7LVF+bUIEqG9jA5eEpnAtG+RZVMVIYc1rHEyQZ
23dDih2o4h2a7ngVzqZBRSHscXTX+wG1FzX4FO+JXBvRWhk2jY7Ko2aF3bTeNK3c
WbIzsHcK41SrKLBGeDgJn07Ij10lyLX7Y8sCNxwU/frF7CG9GUiyyl4ST9V+lRuR
vGVAkHX97g6M4n3GLpCH4X0xzvVLB/SXuYFNlOofkKW1uJa/mVP+8Zng8HvP5sx7
6fzVythON3aWsrtF7xow1lrX74ejnelzElKbd0iXAdvaf8XSSEQ3R0k3Z3/DGNQG
8zfDaoi2pSOhnc3hixrdge2/fhRfSLAycuhrY6xAXKDfMsKTMoZTfxDwe1VXTPqB
o9r87yXKtvtQ8mdTuRVB8K1neZy2hjM5ZKNxhfFr8Ci0+R+2Q7fYHURy8MNASDXo
urmnZEfuwK1p8zOzaXzeopd27QGZaRkoTXv2N3YMawy7psmzDrJkp1y7oUO1c5DO
d98sT5fm4PGHKFQFHRb/0ZCuH50B2JCo+G9JMCBzPpQEEB3DcTSwubk6Cdt0sGg1
dA0jyxVJvIvFj5miPq8VAOxuA9kvQr8BXvf/jyx+dyNla6iuSPZ7AMHR3RpsIQSC
uCKrDl+3kvx9hLz7A54+CbTV/3zj8fSazHxunIv3bX9pWbPw1HyOvFNW3Fwiwqgk
uCVa6/cXlB4s61m+9QuBLUZ7G6DwWLpTHT3IoVZpFJYZzBPpl+N4Xfm547vt+zc1
XmI5u4e0nWD27zU8186WdbA3OAJC8F9IHH8WgOC04SlwRx5zeEp58LzaEzHFeoFG
bBexhfa5LYPbqtsGLIryXLJYmOrWATEmwSrZ+va+UguEviQyR58U8j1e+R1Lac1V
SmEKrEYrtbbUwC9w3g6AP9JWddMpGaoZyVkt8nGQJBsa8j2AwUr6Ynr93CFqbzJ6
eC/HBhU2hM69hNFELtJjygMNStK7RqfVUkv6hMWeUvnKTUgK12Ib1Ntf31nAi9AS
nBoAocrAZTpAguGsVtkLDBOP8R79XqAXJHsXA30H1PqFhwk6TEplsf5wD5VWoCIb
BN/3ftjXIvmGRa1BdVGO3HjdybsrUMyLlYSjjz31KrCIDZRoDvG50kTLrPxWLkF+
yoN6Ripxy4iOcavq3SJK2PvPctj16G8tjOT/MtVkco3RBSs2dt0EYQ5BJ9TLOwa+
L27COveoXUD2jc6UFlP4b286I6Ry7+YCH/vlt8Ua39C0eFleawWuKiFsd5GGCV2+
Re7yYAkn+129bGKZYYJqM3z388jaqW49xStCf/i4gYabVjgyORhjCOG+2JPVrpNq
x6EOMPieVYYV16UbHCYnb/rbO7sP4YHPHngpPL77kNv61J+VoTqza8VxaDhALHIo
y2D0dEvNZvF2NyEDY5EcdfgPQVpzYbqr77TV2d2EbJTzEOcVXCqt9AHiXgiE23l4
+YyTuJwL4s8iipwXEOLJK004EclE9Ci7Vs4VAj87r2EsoPZC65+0qJzBNjWT1dyI
arrQc8nri/M1pdKbaVtKkga83wbPA5t1MmG0QHonU/v+mhsypZaOgIP1LZi8L5m2
UezynkE3bMlyzwkUbzi24k16YmxqIyFNMMujWKeFvkuRQWPL7c+b3xf7jr5S4VG0
59gE4HmirR8aKx5NrPvGmS59V4FZRakmIzY1VT2lwoTq38Ak+5HFDbVtrC2AaTwd
UcYgQ+dWYlZgrnUs/GgWuG3tSkpzny+OZC2Hpp/Bbtf0rwz3XyZXevGbJqAryoie
r78Gcximm4XbLbT0b4EKnY1VR0XJvU0QLbChgSDX2Y8zvccraweuLgwTPSh0MdWY
b7I54Yh3W4YdEcyBiWKIPDrLxx0sokeLXquO7ZhGQZ5tUmifvraND4RtyK1Ds5NN
Su/7dGa1sEngElQVDOFdxuY2yYkT6npljdeJbhuEqI2Y5ohvdwjT9RTz6RAnBekl
LxO0+X4GhizNUxQD0n8nal9KGDijV/fgV3l63HgN/ZxeaLjygdtJQ5ysR6hwrn7g
7+jWE46/5fyayEOW65zhyEU/HvBn5f+eic6mzRTcEuHcLANxF0fsSDV8GGw5NPqC
+zDt1zPNH9W/HR8oJpCe+dwvi70rAVeZQvWDN7RdAQFNeLFy9JmcdXNWy7U8yMUC
3F4TqGHQ2Pc1ohAZwML4myCij8Ajax6utIYp9jNKNYNNWqxdD1hUymQwnWq+6OVR
4KpV5uWrN5uPwvVuqcS4elvs3x7M6MwQCSrS/K4PTGd3FsA1YZ0L363z5QyfQf87
Dst8HY1Evo0fQuy7OifnArPIz/A973xhbTcG0ZKhZPhQRqHulTY9ycNpsX5uu5JC
gcoxv30rGCq6x0UlALUSxvp0HT/kFU/QpM+SEgz3bzJ+sJY01IOmt+GHdc1J+4mN
7OOuIFdSafJbl1XTjKnvw3uIdE/LjBvrbd7ZrUQ3nLDMA1/PIPT8+e1CMjowXf+W
i33E3CH+dwLnaeLrQv335Qxp2kKbvf8gcpbzR++nqkgwzVU1ASUX1y/PEkdrYv8G
0Q6GOoVaGOzkxaMoOrJdshVdho8EzlzBILJmF3xwWaAAtXLkT7unkIX7HuBZ7Qbw
TrwHNqPlPL78bb3H7A117Q9pDNTmEXaMisuVJdBZLjm60bR8zfGqrEW+yB6GX0Nq
BBEMzGQrKSAH0E8iDY5Bdf1jagGuqbFVda5NhypGEzdkomEwJrt8QHX8TmHUdKQf
Bp+fNLpshvEhLNJysIoT0uBJNv1gCiuX+j92RKZ9PUNhrdM6D94/i3Q0wTHqDRhB
AIrBsUPo+E5UOIUVoq+eeS0TZ49/YSRjIdPO/VogbHm5a227HKUxrIxGPijPKdzw
EDzy3D0n+elUCtg2thehkBAcPMk8Bjgpf+hK+OOMXgqJe1FdNwtiL7LQewoTi12b
Y2WUum70HHVgEYk4wNueMNdGsAqwEa/BUCF5w6imSj7Kl0iA7wfaTZ0SicW8IyzS
qP9OLM9oZ2layhoeeTDww6tPYNiwALQuBIc5A3Z2TrevqmcgM94C/YFF4l9CTPPB
gwyiFRLRUckIx1J/YkHN0xUBWmEhir4Glrs7QGmUVCCyHNblwlhpjR/Ds7wT3S+h
BfYOV7c3LpsRZx/YAtaqCLQV+DBV+cx9k0MdBS3PKFlXW8mhdPf3eaaU0OffQsiD
FNOlHUt4gOkTFjYs4cTUe+HardbjrSaJrVT3KjLsb+ABlCJanZ2L5BklOqsN5BpJ
UmzzyGuC24uSLCjwuCzn6REK4V8yW9wpMG4WL7XqQ7Fldw7p6L0g8lU4VwcSZbZ9
GswWdR5PKUDKQ2vGI2Ay+1FLOSzSRzcL0MbYBxKWzqEo2EFIH7MElAQHKCoEk+Nv
blSOYVxcvlsjH/EzIvB+F7GNZ4joIaqxBJgeKvZY3TO8dRlUmoI17H8IY4uuTG6q
u/r4u5CqWx/gsbl4zlyqgNdp6Aid3Uxg60/GBt4p2U6if4uKtKRJl6WAWSOTaoMv
GoxqvR36EVDWVUtx7JIiQo/yML55no/hqwRfK287TZsdIwBxwovFNFI9sfLB5I0+
mbKJShWZX4eHRMsUbMJ0DIRU2DCKGUvnwKhGGMsGKWC3Iul/gwQdu+0cME/CsT/Z
KajWWQVzGSHn3v5s/pTlFAOJycvokAGeJ9w+W1lOJccQr5Ef7ZvQmIeNqKRjTlWE
IqnI/FGi5q8hJxxq/jQeyuLxVRfTZ5OfWsl4hatQHYTzHUpxrS1AN4gtID2BbRJ8
akf2Lg1QQd+WTwGiAmx8XTzv/0y50EJaNbWRjGmlmOHEtSMgAEettWzyt8rPVnCj
c8agpc01mauW4ELLXGBou+B18LAQZN439HlmbIs12PTUcGvr5LEJqGS/M0JLL1WU
4tw8+o3ODireV9iHOkUyUzraotZ3DFj7IHLmx6vOtDdrZtsIcPQPfts+ExJSu98F
muegfemKX5iwcTQMHc2mrYar+3y0yMTrAhFPwJYC0bZ5B382nHeUdfxZnQFcNw5i
LR6sXGps4S+37wq485aa2WeT9bh+AmJ0ZnoSiOQ4m5+Eox7Z687QP1fGjIh9ff5/
jUfWy1fkmWyux4wD+o3o090A4lhvQlVKoEfczO5pV/utwXiAt/4dUZrf9uiRjwo7
W6f2FEmlg3jp956ykjFDoKbGlBmDNPztJZLyz44+tj2551C7BRlBKc+gTkd5AkaA
KHkg5oaOWwP6GNtF2vUF8fd5y0uYV/dY2lA2ik263leWNtJ+WtdnaxPvk6LPCU3U
+kFlYKClImGqsM4Jd1ujgAy882fQGNpIOGfq7WYlR7SfW9DAWzGnYCepHZrQEbw8
hjhdk8mCYQtI1TFlfETnB+WuPoWhGtPyqs16oW6WLJ+JDYLJD3ToEUCNdA3P45/j
1ap9DFnGPZOvDw45CMCb5/H8oPmIH7GvzRptcvIui7wPbnMfNXqiEH+igBBuUFB1
9IQ4Zqgn02sHLfMB9S19BnB/bJT+xmgqBD1M+UFbf5cP/ey6m7xWSdTDhQNU7j6o
885azWX+y3sC12m0vD+EqBD8XrjzqzTRePBhTIGrz+qcCOxOpoTUhTP+1rnLq+lF
aMxd45uya5A+zUuMRPYt9UPmg+OpEMxJLyDDfahCVpTmwCTJxnpEZkr3FsDoXUsf
5q87j8awmnKIFVNTw+dtraLS2j2S8glxHezgmgfrPCH2dlJQgvxH/6QWW6A11Vcw
fF3af+iWQCggt/SOCssyB3K8Bgoi5kwAF3JwRw9JRy3H34a9sb7Azagowz/Znuxo
HyZSKSFHKqPUGw8W2de672mSZpr8/nyhxQVS/ClB+f8TSI+PXTm/mQqtYJ3aW7qM
QvKNfHjrM0hsG0qADZ6APkwbujxPIgbNhULrh+3QIg0L3dC4o7TK85Y+rxSDq3se
ROmpIZvM28fGHhYLAljWPqkLEaYpdw/73PBjYmxdAmu7LN/2ceL9craSdksTI9tq
zVKBeVaYyzkQAEPEeDBrwQAYisV/SMOv343VucuaNRCDDL6cO88pYSviuSUqC04K
P2m2l+StEn/YW5TbHX7t5RCXXGDv4QOhJDsyST33wMuBFzNij4nR0vGLZ/70Nfz/
qkVD6cFakMe4ddKi2VsHAhlE7G+teiNmlYdAH44Q5ApFRPAX1JD7tYcR+4oioD39
/D7kN9JHYVe8aHmKQlAbbbkxtZCs2gnGEiuSrl/1mZKXZ47OQ5z9Hf6pZ4B7vw4Y
OILkVlYHlEQgsqyAfVLn1m250m5Jk9NZFdqErm5501pZLXu5t/mTGB1wJFTez2F3
aeKTqLMWi933ME+kjHZfrs51icV7Xx1eCkovsswVGGxpvpzrGyr5wMpZLJL+UoCX
NBjXzqd/wy/wGLkfPNKfs7ay+mfT9AxWKWu56TgFD9+my5m6pvoOe2e23/ix+JPw
QqlGmU4ZHz1uIDMIyLRtERzFkC0yCw1J4kDD17re7rHRLfGALaVgti1oQHlz0YYz
ldZ4FxECblTIzmZ2ReSU0a9P+NGUDAlmd1rE+022OaxyvSL7jZSuYDcxYzGvMlch
9bORwuoD2Q8wtlX+BzFA5LPvCfTIUWFwCm6aY6rkgIwlDr2+11gC0xkGjwQTzhA1
+a5VqsQkrWWksS1Gfcva5hjpBi1RN5gDUYojXeHegOfsJxXHMPVIgs9jyyZ5PeRX
TUSVM2UU2Aov/aoVV74MLnWnNMaVtEl2pzMBkQDIVyi87undvD5S43GDU4MKWry4
DCcjX/2Eg7MQR2gAYU8vqPD14asFi04NHDbsw8r6fm3NqSsHPOdKpzNLJnNN3Apq
oscQ9PFQOUTt7YViu/K4SXdapwJIkwv06wyxNaSkXZaNh8lb5TCD8bD1d9/qn+5I
u/4o/QN6dS4RmDUBKx6dvEdsxXhlZ+GCu4ynqH08Z3cYxNUmH6zMPnjDCs7chXkH
Q06aJ0buYxOUzrXB0tiwyHes4Y4ilfuusPlxPRWx9NFxxhDsmM1Mp91CMdBZ7DW+
orgzHuqwLUpZuPvFMwktlApHiu7BbDPyrKIM4Fm9ABXCVIqfxqDtwzrzJ0cM2B2u
B+lI2fyqK2kuJVEvs/O6bHoQUYe3gRticI7l46hKPRq49XpAo3diA0Gm/blJFZss
Zndf9a62qSIuUQ02YZfsffWQUalbKhwe5O7/FFLahIP/xq0+Q0grMAwPPOv1oap3
V9APUMehlSIFwSOdTb+RaionehFDOIv5zjQvPJHvPYb+tLS5xdpshv6WG9pc4erM
ShoT9dIJLP0JT+igjELNPVY+dj3i4aDdNIiAmdo6q0zImNV3MrnfHb7hoeA+2hub
3oNLwlFip0g4rRGR0PIilBmxu+qjBNTjHK4ANM1lohavBGPl2qFSuSCDqNybxyK7
zlYjzVlKuRkglkKPFlbTYxRN6cq6MVESG0aWgDmus1KQRYn27uyX7dkJuK8ZYwhV
zpojzMzbsq9j5qSrZa6KPWYWdLJOwMFHTO0cJgpck13vaL1Fna4xMl6SuQZDLx5d
5aZ5S+Q40+cY2RUdRtGN/gHvmw5TKmruya+iOh7EqIOpQCpxm3TUQhNKOyipJl1x
RdKfpmJyX1Xg125K/aEqYpy+HmTHG5AVSk9WLqMxsTsLcjVfFIqwtjdUltS0M84e
nJvP25B7RMF/6W/rfTTqp4cNkCFd+1z9IunZJYnrFMIQyrgza0r3WPSILX5ZFkTh
Ol78cTpX3GQk6CEI4Sn8I2PCIji4PEVHC/tvMRWjZVfpOkItHUVOdgrJ8e95GwZ6
oxMf7eAYChTxTGuqVHu21HXGhWws1o0czPKLw7WXKZDJ0Dkr2GpIZIVgldjBD7WI
8qZxOdHuZBFDxy7p6+X8HeBTj/+5qtZwbGcoWqx0zYuE4zqVhtlXPFdcAIB9vMtk
+byjHJyIlMYEkozB5z/7F3AjG/oEDVX+OhMxB3w9pwOWy5ArsBs2ECteeS6tkGMe
5rHHLoZq013HSoOLRQ6iztLxjewxz+xna2ZjYIAUlLZ3mW8GKM1Fr4ISSAk8BnGl
fqH9/SrppE9HhqjE2KBOOI5NOWqoRvWY9WqHa5fR2m4Xd28FogsvEanTYENWHJiB
q3FEcOzhMrgn/AyH4kYLZoJ03lT5yV6XwoQHehEk0NVRuUTavhJwoHk/fViTksHR
7KFvCgkrPBK+ZroBV9h+bRoKVslN0QJLgfbtMdTTXK0Sn+Y0KoN6xosRdcpOD+3I
W0X2jOFrXcKiTyTiukBaEZ696/xNDqXVDNaLRFRwbhCSICF0KS/6wCQNeNBVrn9n
2+qHq6WCBbjVURW/8u+vfayyDBMj13VDgZz4SJwokJvGOKjwnIYtw77tE2Tjypt+
x+Vql1gXxzomGEtbxLbwMxvfW7N5h4UGlNmfaPq7yNYp9AOA1oIyRNSnIYQghmDs
TWBCMB+QSyDm74i3V/GzOTXZqsXRRNZjjkyTPVOXD3MDbeeQcLMVUtXDCpgiBH1a
P1wQjUTIw8hYivjtOMyvDNLnCfI2nmeUnZOMT8nJ1T19N378172rdZR09firPFBo
UH0c2auNhORlYHBchmWjnGZaUg9dHdVUrh0zluTeb8t08h4qSs27htH+SFNLfrV8
nTPsnGDlsIjAVMFJkeiG6NbQ7EwDWeOIaVOFUTE/4/Q+bWXeeYupBWTwFCtTqtNF
zFEO0KLp201UOb7aJvMjGZsQYxW0i6gDsRwauLthZLRn9862GL6WUSgu8Ci+C3nG
x0mV664er16muRutlh+x/SzrZVHvXJxhibQB2B+AtBnPRQaoM3w94GH10XsYk/mz
Iy3wbxI1ctPHfqBuoE70g9rkAI+2OuqveLfW9XtfiJiFU30Dp/ixbFKT4LwurW0W
2q0ytCh2GoD1gKMRiTm8Mp2uBsR2IAPUrZu7IhIKo1sK1BGBGwvdlc9mtSX2RM6h
jcwVFOmy8wMpBbgs4pOXC6ZDPsq8/FgFmQw3+VMS+qpfWKLVRmN+tZau3n7iJgpa
WsmFfi3cf6QHzlJhSWdapXp3iiiOFui7I4o5oHyos6SoF0S3/NmqsdUZQznDaWpK
ksGBKN1vh45fgev/7S1oBowJyiVOVt4m8Lf6/VuonTGEkkN6fRuQfGp1UHN5yMVv
xMs8ui5GvxlW6eUWCGCcgFvJ9hd/+sKADeUf4TFSUji+DsFoHO3U4ohIqL4GP8Cd
xssszsHa9AZOAkWUvyK04HvnUVOnL8I+z0oJa1fgeEtmwd+QMMkO84q7nCCwX5Oi
clCp+iVrU3ZCGpJmzwQxRvGfKhupNMW4kEL7Ke4fZ8SG0DfMtYWAMYSYdTflKsDh
SShbCqXXQx4MomZAhNSj+KU453koCaoexV02QJcc2ey55JtdgNS+RUm/Oh7gcXel
ERDebxYK3Zhvs+cmxOqrGxJluMNZUSibZofOmbjT/SMFwxfg9GTT0o0IJ8ei/yMK
DxN4mYVjRRO3tVNg4t4BfyqFYYRxNvFxcQTl30M6wzulTSsWiW88z6WA1QvN7xrP
2U/+zoIofnD2u3sxjIpxpzENySY/lnAMterSxuJyE2ffF92EMPRur7fC9sesz/7f
N0hFUINDkxKCTcuGW2tTaYaI8D9afeEkSVC4nF6MtxJLgCzdd5ZILLUgMhv7lT4D
uBPJQQD6/8Fsj71YZAhCyrX52dSBw3+cIsIjcChYSJK8lEfdRQLL4z5TFxDmwn0x
FYoOlyITPtn1P04cTNudalwIvcr6PG50TUfVaGAK0R8TZaxK55Yzwr8AeSkct0TG
c71kFsi7KjbOmaitnje8l1hqoufb687XShXw2fFwyq56uo86NQhVWW2VxpALOzb+
nFoAeWaVoNaPatBu5GJHMMXjRXGaa8tCedFHZGx267T6FsrxQZ3xpBS1tVWvT+h7
PrlP7+oWlpB1xYS2AFsYAM0bTUt63RoTRixJ8KzaEjs0oY6snoAIAHdUDtExX2Tr
wq/gG8LDRdctqhXaFsLeVW7ZS8fb9NrHJQoVRBOe4iKd+h5XBb1JSVvZlC5zTf92
UfXOWZVctuaLFOG38f/F1TXIuFvKbAMzTWHXm93Stqbo4p9VDTHpFp5cq9DmIakn
bdegFqHAn18+WUccVaWkDKC+RX8kR0i5WCi1Bz6acnUH6uwWljp9N+JMCzIaGR5v
oUKKVQE9+4tNdL+vhoPp7h968yVnnR0cZ2TxXStNyipqr+HN52peJbXBS8knheMQ
hX8ANwfpSezEx/bzO+k79RSyjEGzcPMrj7FhTaMiA01yGS7DIW4WHDy3r7xs4lUz
Cr/5lQM8EOanZYZX/42/vNyAtDxL+wu7tEeh+6USJ7OqxQkIhE2JmT3hu74i4N9j
KRlEJ7LcgR/UrKZtwmIro4JlOMsQSH+dTNOJQZ3jUBVRMM2n5SXzDGWstLfeAhc0
AX3IpkoWuJfbrsdr0MQMLYZcg84iVwKQojbnCdiF3mtxITpxtwQ9wqwcHPQlUMo3
UEGKcJmJRMEzr0tM2KZs/DYYvMKzsd2M/0qcO+VzEaAJJej2AzOERUjSVLFiWQyR
Ednw/+RmThoUEIleEhAeteppda7c1jIhJZqBoI0+gxmlYWqSvXn0LkfnMIOOrsnz
izThXcN2BubZZKTfUFESouBTOWQBH9elAzEu76j4QVlrqiwZT59Ux899wTFECCwS
fPIjmSl08gmTI0uyxo3mRHwFTVk0en/nD3DU8MAolzPGEiajAOHL9H8a4iJ/9u7R
0taesLiUgD/vdeiVHLuIJQbRRqPFhDQ3bYCJ6JRGD0G23sMTVXujIKRAl16gw8u0
GEm/etVTrXuoaiq23CPX44se3IRpJ9xZzIwHWQBmeB2l6jMe83iXlARodDLGsWiK
VwlqGcWhCLppYxrmHTwTlktV/Gk1qwXTD4vOQZ/bcO9m+06onXpbDhsheeg01zUN
ZfDU0McAR+sd3vgmo9BBxEjK4VmrleKzM1FGVP75JRGHR8s0EEhsRVN8idGXKBiy
JdSFV4EyXyAZsbzVMB8S8dl1u5rum/2imNLdPQDUniquWY0ff6u/aV3bszNApsyQ
Mc6luyJdZ0jGkrE6Zk6beLgBMEM79IorPid8nY0RZm/X5e0rmuk3F5W4jdJikrNF
HgPLewD47YOXp9RxMdN3Mwj+3p60jF4TkoZZvCtt0iN+M0gK4f2WrMOE3Fj+Hdst
TKYl7LSK4a7a4a89tCzd7CyKbXBzaF6b4+hIcVPVHrGTOrPNvkDyMqhPwoClFATg
2rGA38NK/wW/EZEZeiO3hbhkMRtW1Ya09u+vjznmWRvlGM1Jut1nay9+owXMgkWP
XBCHbguEozFkWl4TBzijn2/k9a8EpZdcs8m0Qcre9cqM6eMzAynZmXskM1d3+TBu
L0BYpRge0q48iXJ2d4sQ7Aw8JkZ5kKZiTH7GDLnipW08ZhyGX0v38nHeu0haUqPE
TGp2uoaqGsvQDFT+Fs/Znr/w/jtGfaAUi19daBaGRCLNCbM5GHCLQPiUGppM58vZ
w1nFf7JnxfrvXRd2XFtVJW2clv446ug2AaV8p5VB5ZnxpxpR6hNUTwerGY9UBFrG
P1meYwYv/03xzjKdD6J2+wdnYK+66XrR+AX7oaEXooHV+JxBo6ESDUgTyeIC6TFm
eP35KBmG77d333GDFFLFeEn5G5SKOzP6XGo2VIsBqnl5fFOKflVnCT3CxsMNE9XY
mz7VNQ4bpM2vCWfWJmFd0Q9VA7kePn2O1+OQJumuxQwW7UgafhFeOjY+rI0pHNOK
lKF9aJEJTDtOUJJLNBu7bNNnRD50qtrrm0ltpyV49IMegfMA5wgVs4WqGzXvp88T
yogQO8E+4X3TlQ6m4BK1LdpWRu+2XkA/4Ezt++3xeUyZamfPeZ9PYt+AqsKWKoko
0rjG1AVyvRtkWvL5GGpw4pC7+A/FxC3wghorDu0osMjJRoPrdtOFSjc3Urg/zCSm
GOCyOOOyLalSFl7I8nC33rBM+cV8BeO8fHKUqxGO8V3I7743qm1dmwPji/uFdcIw
bzDQ0V8beuQtjoW7JsYq0eYUBOR0Nqfy/euBWEYL7bEz+jRrjA2W4qnghrpGfK5T
DykVLtFoAo4Iw/8tmjq2wnKJRKA1rsDFm9WQ8RAXQQq0ISWrHP/gOZqRVlYYe8lJ
UVK6zDDhgAatzj+TfD7uHA/mZpM+RNIejw85+Yg57+LjOPHf5tTeQ0x0OYeN9Yr3
rFJjLLr7Bd/qtSEwvxaYiWUGW2NGcIZ1n2YJgUsmw2j8eWfc7YwFmrSGAe4PPf7F
Su0kihsrwoPa3cIrKtWyOSIwCI8OPqK5pjvwLFC2mkiqDYgfngf/91bCBbq9jx+I
CnKhAiFJMWKiI/3EYZun+h6sicdeopgHRpQudXc7s4uIfVoWNvpft/wp4SdylN7Z
AyRz4MdHvPvjQvrvl8vJHCBj2fBuQ8wPiIoQe3O/Y/bkVS3YpJ52EJuuScyU86ZK
lgLcWg1e9UnEnuvraP93haAUjjE9Y4tGME5SH0etCz8b+ZZlV1tGv0XyPMJkzzNn
Uat+WIQ/RdSWK3/3o2ibJ6LJ5Mzn324d5gM2qxO3Sxqv5E83qh7VBNVnCOUdtWhT
pWLtqvp2j5vF36cNAa+Gz3MOJrVQ3raulTdA0nT1bVmOlQELoYNQmTs024rDFaEg
19woZf8XtLwCAmCjQNjgDyzVxj1TKTpj6pVGMUPFDEDzE71Llq3NN6DKIyzTEw6g
HTXzBV8i01GP5X1B/cV/RSQ61Wv8Ye1nsuYo097DHW/CjaADH/Wz8Ioef08yC4Cx
I6hf+bf4kj4N3XapyWDju7tY2fdNvFaNZ/Hx/rz4chXmMTcSgiRmVR0h6d5cR7E/
N66WY2JUgLgmpnTFDFHXg652jJvlOo0INKtim0RGb/nW3W8fWBzWJhyMqnrWpmXD
K4C+O58VJZKKiinuyL2c5Tau6e0f5ZTyLL5/FVp0/RcLAgH0lk+fOi42HQWg/c3d
/KZM+bdZkoNJIuvevg6fVK29Bgq9+MZcyKhoFOqLhxCd+YZsDLcspldwjtS2hiRm
ixHJumwmOSSHBIuGvLzG5rUNRATE5Gs0b0jUInoJe/28iq8LsMiDebqWVxlRsa/n
ikjROdBMFT1SAJPIUrSM57LOkxMneD8By3iyxW90LnC4YtRYY3TwraBenf6HBBNi
qFDS/f0nEcSP82WcJARNzUxVj4i1tNy/wGniqMIVkZ0vjH6nftxA4iXVULE8xp88
vskcLRto00Pye021CPXQHOQgOh6yF0np2Iv4E3snTiiBfzZwEBL9190ImcDimsTi
xAshqoOQGwcWewEYg9KsOAsZJ3yuP1+hVC3HKs1OgF9XFQZQ22QbblFmmtb27dfc
otbgYvJ7tSjxvb018k533tnKE1kiA7lN3/J7pgC/XKd1dPeu1m/cMunhWGeRCgqp
eB6lofH4lqV07G5dYTaXbgA/1i9DSPGC1dr+CD4JmdZvgGYPyDEXpLx+5vHXkeSw
7gvtlKYKlCuQi1gKEiRVRBs9ncOLqge0kvbgkJ1vMsAPLz1whhmGtYkj0YGgIwrq
dlNwv664FMp07yPRn3ERkgBbZVXUBgjxIHswoxvkmWSLDS7GsS1nsLhC9wpVcWI6
xK3DIPOZwZHqJSBRTTP3p/m0N4cCtRZOAXlBe9JXXEp5su5I73xP9WkE47T0WAEQ
CtAK+w8+EV4l6Ax9aF/gIyxq4vyqcmawLJv0Te0AbOesdS8U7CptTJivnViEg8b2
ZM8o9ppEZfFDICTuKNrl6TKNZJyPA3SmSKZJr8Yo2pWWbebss5M7ktA2E099dgbk
uP1t/rrYGYSQbigEFIKZDOjARatXS6njYWS6OqqKiMcoBw1baVd4vE0i+yO83ZYl
DgiaurZSzx0BB0gb4QEIc3pf/d/4YOcy9h7CC60zALWHX67Ls4UCL8MzKAmNpUkj
TEtTx0F0XFvY/cu+zG4miqVz1p2LOXt8sFFtSTCGpzysvAKbOvf1X10nmgDHZRxo
pGpvPuhEpsdQWBVGMMDWN4hPim0knDmFPgA3CDaqQi8AiqiVlH9/3l3rcCzouZ/o
IO3rHi6l5qbD3x0sjDU5LRmwjgaOIbW080nWlrPZ47YLpVTWVu7RM+mn4ESpTAjK
+SFuNYrm+KA5MxSPsz3/Eg7624eHpHbbe2gRM7/6ir9pzO3/oWGD2YJUAutWq48X
57vRCHm9HQ2tcJQWbbwMDKdo8MJnnDN4TACyv0EoLjQ/bOAfqamacYV4eGz7wGFn
WWt64Gc+t75FSIKCw2EdsuAcbLcTHDC+SkctD9mURcin8rXiUPXQ6QcToM+9ppZ+
MW9eTE6jh1ecdtFAL2V8Fu5Pdi2JP940WhQzgkFQ5cpRPLKQ+dKQEvro+DaJK9sk
8wZvv60WcF65J1BNl+2t1pbgbVwH5FYnqyEqREBPjd2Ouq6yZqF9iEH9r79M5lUj
v4mC+bnhHU2qpYnY/uqxYtI1flN74Fi2NjFSpA0O61jpNBsmChUg5ixRK48PkvgD
Mwd7oIboVRtwFx+QHL/Ak9/5PZZHTErSIX93nYX27Yo5fsKbfShfHLEz8ogaGHO1
8+KiQCCdYM52VSRLmwaQsDylxiGymZIyEPFSdDKd1LfECW3uCWIN4y6ogxjjoqSS
cfhnSxcA9T+e5MVBR+dx62WfU8P5FPaOjI6/82w4BOppse9ZRZjS+FU+WlEWQpca
xhEIVO5b5br+mB8r46guCAu/PpLT3qrgasX3g7XddBDFIKr5l/AihYXLafnbXzwP
h+CXxxJefd3JXLa2cn1x++0qsKWAbAO6mZEsaiAcY1FsGCJ1duPSKtyZd3j2sXxk
G18zogX1Ml0jPtFGP4KUryBXNCoAlmObTnM1zdHGTeHVlC85AtlQdRCYvpofHNSz
l78IFbx9htLI2yd/HeqehTIZrNE4V99FEa37Zftvkf2ydLFG6/GiPnlqHtNNu6Hj
ZnYRNZAmewH0SURSXU1pHgzHTjQGJEaSljaA5GvFzKajUfDsTIyCKwWQ84dCFNTv
gVs+N3Co3PTYQP9XZvSSLrT30V0QEPIpls5iKWEbmV9L7YlPFdn54H/ga6EAZClr
Mcvo5I27qcq7POTOIHOz6maiuHsxeSY6o1crNwDs+pXFMpNN5Hmus/KnpYTOSJOO
sYSVrBLHO5N4SOz1dz0DsyxiOlAUfYb+N2z3mei4JmmWDYD4Ge6OIyNITKO/Qr2v
TYRQxx4Sbkj8fXSXUhbQk96VtCBhpMcdTdEDRTiruPgl/UmcITNyXm228UtIPunj
VlJkv20ieKDVM/BDylYh3WVHfJL8PX0Ov9xVAZRhF64SVWgLhN+5VRyHorOInIW3
Cw9mrNLa2Twn/gh9Wq3/yPsFyLVGRNCnQygnRvWbRMDQApc768ERGNjYmJR2xM2l
3SvXmYzerp2rFix0HVBC8pzmgGCRjDlgGJly47QQjvX7EgPVxhakl2x4Ai7QRJpj
7/fr//RdeVvMipco47Q29ULQsCqowxl33mwvvztNoQGoLrWJxdCAZMn9jnkca1Dz
4QAtcxeSkj0hOJH0FQl3F2LyA7EDNm91/meztjRb9ZipVdLqhczD81kluQfPLoLG
25MH+1lTE0F80AfOU73z7V8bArEoNxMI27rQJjstPambvL++xQ1pPvZsMfiggTc7
yO96YbF5p1yyXlveZCHtOH0wwYguKTRqjn2sDl06fLuwAmLePX7vkpgGDH7NS2p8
7JG7QFcXhwMtnGqzvv2dSKqIlPRh5TxOzqPPhcVjtpfTVHYoPYUkxT7BmbGpwA01
0vb4VPyyOpqz4EaStDKVz4rdZ0IJ/lmnyeD3d0t0FVEJyp0B3XwL/g7VZNF7dZgT
ULUBeNidz3XAf1Rt6QN28WQfn5KkP39v0Ys7dEU/koZMmnWwaqYUtcylUhHcxhWQ
t+0vEIS3BS3VZ9u3KG5pQJbB+Ba242N/M3jNelBs8VYXHbc6mUfuoGtDASHW2EUQ
yB4IkXvyHD+PztOI/xyuqqVhxHe/kTQIYj5uStsdzPeAZCUFlc6faXg865JXasB1
B1RaBJCLxaSBtJw8YH+YuaWFiAZrfMWqDnruu7R0Bxm035bRsoRvuE0bR/W3IGae
JXVojOA7v3RcGHJ8GZd+VYs8NToazbaD9ETOQmCePwu2Fl+K1FOUIPgKoSSQ+m4s
EJJlLRtA5ts0pzYQM0F4bEYV9jJpsvBWltfOPPko4RI2wviDTJhFn0huRWpUgadm
D0AClwzHUsmcGoWKb3mrDC5kMiv0YslvCzV1DZuAGZYJLprRvBAo0hTNJdFxhhZ4
S1zKr2riX7oKFnkiDY2/YqxW4K3yEaE35l95Lk2ih5RAC23O64Cd0pDnDQ3hF8fh
4VRabhb2mTYSoNjR84+FI8TNOyFHjyCteab6a1+u/Avk+WyrgxJItQcO0fz24I6E
BNFPa4OS29H2uPMPUbklZzBdq1tN8M9/iz1ZCkt+qohYFit0AjUPQerLsGA9FSAR
R5neLFd7QMwKAdiAbD8KM3m5H4PMPtdc0Y74LjJpjIe2FGIOsysrOfFLSSPlGxfJ
9quMYrvvDJrZEEWCH9w8V5L/wSAt6T9/VMdR9prtmGEUbLLX9Sl788IfdmwXpXt1
Y07VqzTaXk35IgCgRSzOCX2S9bUn1eCKYLc2SrTCkGP18Li3CLANHFMRLmCeqgJN
oXFRxefFUVbR43/dUvO9S0/fbVn2J58HYy5AZ/LtjJzIbx1bdqfx9MveFg/5fEDo
LiLfC3VFGu2yKHSBd9BNbDRhp9lsdsAoMRDoFXmKGNU5Vx6oN41F2EXxKybuB104
oQ0EMYFtVKZ1Vil6EaEPoAU44y9en+AMohVTfL4lFsBEl5Qp+3RuJuchJjjnb4/S
UaxBFAghg4kSpunbP92oKSbkqxtMEWiBmgz4dQM/BBCb8ycR+4ULo5kW/PCwl2oo
apHi9UaLjX3vNAuHhnZFR6JMKraoi/Q3ekbxcM+sag17n/RYE5STa3f3qDjlrd9f
5Mlfl2DoMoNahZjRX9n5xPUEsGOy+LD99TpFQHI5SHc2GvUFbSHiRLqh1234zK6f
n4r50IlV8wm1VHVc3xT9jtaXjIrpUd0cUuLGFGjRmBn+Qljwo6/lYMrSsKlKSKln
Xn4a/gNQ41fsPEP5X7EyLk1sfBTGg1LjJpJ+BSyWxU1yuVv5QWT/A/tKjW9DTq/3
Yzw/BUV7ZLw308RJCWBP5neDlX8OIp2qzwNwFJI9eUjc53gnwqTRMR6UA7FWdAQ6
9RHJNnsP76WykJhmwXOqXaMeAuS3Xp7oY0CO6zqnWwSQKkX1js9nmyWXpnu8vXsx
0YjtgLFULZOqffJzJ+EsJ41nUtYoRFQZPqzXZWdCQ7QwXpXkOwt6nZWvVPY9Fg6/
emclnBIvMYoJIn4mckdfliaHCKh32wnuVcjCjCDXNhuPCSC35L9hRF+xNvzMIUIX
QBX9Ar2pIdEi97KHDiPKlyaVGt5UUBxiVEL7coElEaZOeliCM8V0P3A9gj3a6QXW
TOg8xQLgdcrmwK7zK/yeYCOdL9Hn9kH2PrgIkdb5tuLq9K5ZgVpZGLGXo/bZrgVo
31rmHZRcG1fzObZ73gLWHBlH21CHeQ8OgX/OCmXgFsGgdg5SjgIvYpbn1iQK7fRP
3OGsyPMOSmSNoMXzyb/Iaapzh4FQfGB+W+kcWPbmGcFXeRo0/1Wd7bphC/M2iB/u
Ggm02D6i0vw8By7+/wMcBtFk5CPQW2TYGXXduqAAztCjAzu3E1rjoPg93uIH/FI2
y5tSq3qGFpM+566c3QF1CfyQtXQKmJ/tSbry5pF71g1bgQiM+MNA6bMwo1Y7sQ+G
E4lk2R2xcaB6kF4ok6lIaEwSgYa2xEZ0dMTbhL/e9OlYXHBYNbw+xK6Aq2eoyaQ1
KdqhupgB6QbjID4jqv0hnch+cITkgCMO065FcemE+m5hiBs6BxRcEoD7KPcWFKv9
FiX5hjqQyBIndh1dKHt1p698VVkSlp/i3GXYvZet5TTXaoGTwGG6wD1dQexr4bn6
hk3yZD7sFGI6yvA+t4MN213qIUF39643m/5a3Nz0A5mqw/tf3IiyTMQTFO9Kt4DF
yHzNVGdCshY9DaoOuh9QFs2rCZjdaFHWFh4tgc8Wy+xIUSikbDj704ObB2wkt5yF
q2Dg3H3uZVRBK6k+qSXLPPVxEvY/tV8n2h+vu0QGGRd3kOug77fuS6ucDKp7abb6
5p+gDuCG2Z9nBm3WTWuXfAbkbX9y/axSeAAaYgtut35RPvexYNlNuue0aKjI0Q2A
SuFvdhaYROjW24SgjejCZ8zoyteQ8k6qrK2Gs/DhBYGwOMQEwta2kN6yCrR2yjDW
pOw2ofJsT+kM4/mqfj077/XDCdAT4L9T2u1qveDAO7V9DLalK4PE81X0GTkXMrMC
j/scCR6wEDuSMRRTV9lgEHUNpjnnE6rfQbSLKRvvsKQ3jI24gjlI9U39qtRGviPN
xgJceZ+V4gr4GU1Z7vqlJNna8Pk02x4IPgKNimtpyHlq1j8XXidfEbo2tQljsFb6
EfPYA+CZ29b7TBFYYmSY3GUHDnHXJ3NmbB0X+LLM8EuXVlEwSGoNjQMih5NAXD5o
4zzOdimYFdBISWiqFyS1qFw1A1TBYNcN94YXfzaM3vxWo44hcDnvBZG7ZrF5wLRy
HTcQlPg8TV9FpRy/5LbQVSYj83UzUmlTg46SOxry8kokxdUHR0KXgjKHlOdBZNtP
aJP7trYKjsywMpK2AOzd2IIm5DVlTa3EJGxWtOL+YdqennG0XfZilUucUu3U9MEm
VH+U+4TLzSmDGJQsZrqpzlwNZQZHPDC59Heorqt4ofYuaaUmm5IORuWOD3HDf4iG
ZDHgObQ2+lh4NRi4k5nvFHxNyC66IEGUqPMkoblGtBf+2nYP0vpCjhwU+6Gpmb5j
SGtbjxBGBnff19loPLLD9YHrCELffgDWtoZrwDpiXYvfGdqHiWN4zyn61lHBf28j
FuDeNfIUpNUfQX11ZpczIkbcV2Uxbwoo6mghSRzuZIlDi9b7Ruz0gCeNsVZwUfAR
HAAFvvLUjy0l4G5Kdsece2kdeby1dREXK3CWgLKsz0sBAz4/jYQIYsyy99HGPVj6
/3fRgP8Z+n3z2MD1Sncozytmm1Xv3xDGUCI+Hzv7cK9ZXNgbJ/Vr0h39LVz2eBTC
VbbihhnMstY4tGzcTzHXfWHBtzVhpuGPReJEKUvZo+GOWRDZ9b/OVj5Zntjo6rPJ
IUjiaAncNMskfMLOUFroVRAJeEZFwJuPwHirZdXmF9GQNtCIN5CKTQacIKnqSoCo
jfhct4xw2Ab/ElxtGbwc9Px6n0tXPjStMMM0MNJB2WwY/R3F6Jdk08uOIwVwPTwE
qXKWslNaG1NVKFrvn78pms+92HP8GD47Lk+b5gvP9Lje+ZYzNrTWPkQC1zfqlsx/
P9uq3/qritjCZ69ik/tM7+3Al+arvl7vb8YqDjFiF2iR7V8s2slTQ86iEHt7bVp0
L+6lycXxDrl4x3sjh2zDQjwsZFB3M9BMuA3iBZe1ZBJIaeNIjVUiKG5LvvatVcC1
qBiry7l8MFUVkFe23fTXbeyiGXwEKkApngkOVtd6F5APuhQPbabA/FlHQJt8nU2C
0TbfWH9dApIYRPvIYuNlbyLofocf/vAj8MQzxYt5rIc0PKlO7etXXBap2F+t7t7z
uBW05cedViJAB68HuRzk1KmXQuF3xW+j9cF+InEY7zLYH/z5oQACW8Fb3ofr7Ami
OJ1tld2khEfYp62/AHeuyYxLF5MDymwWa9T5dkDwg5pAMoungI3BEsl/tlVXaLXY
8iIjNDYN49nZTlMaEnjSn4WBglwmEl7jBTsPVGtNBIgZTVYxuOI49B8f/S2oiwcZ
rC2FgepSbxmYcc6i/+MmLigM+sPOx1cjZeZkb+3Qb5SU6IyGQGnC3ZM42UFpdVds
noZ4JcM1MmvPg6O5gWi/7+5Tsffz6ZfGZlqzWkU/W/QMHclsPyo/JXvo030GjKlp
VqqNrPlhZ+g0B9SEEe8lgAbxDcSc6fwDIyxo91//Ab8DIuMTHchECgr3mmwZGwvb
erxKI4y6FeeVreYXBm2n6acJLKhm0bCigAoBhKxbfLced3eEvEedxT0p0MY5ai0m
QVwVbEVzgENolpsi1gnjj8U3YsC9342PG4mcZIElE9hfiRM0Q/cZ/Gr1rT7VrGx9
hsFzBNMNHjvYkh8y0jT0udXpGqD+laPESwSe8UjaZF5lAW8CxczBFgakCjUaZRjR
HaO0kfMrNG8d49gz2h6XORsd5kmxrPpbilzIAM40OJs/fIHtzrH+vhfSt/MLI4IZ
LxcturBt9sjgFYvpH1fgxqGJqf7RDg60giqbn167xW3MEn/Fe3e82gd2UwrMcC69
TfoFOax0I6r+uz2+Sbcs6/EM/oFyIgteNmIohgxLzuzYUl35Y+fI59UrtaZtzttP
ahHW72pmDkd9r/r/mGblZDasgVOMa+gzAoyDbcObPA013/wsOAgjNzbGRohEzvsd
7OoD7lAaPhMta616ClVNBCgTZg945wAPd1bndIqC0r/BK+1q87CxAzPZ3DCS3tWc
9b00O8JHZ1GeffTV69HvPW4SmgDro+kS1rujGB2o4+pw0cIct4kRqyYy8srsqXoC
Cutpt3APyOS18ZWCyKFJjmW4rgKasAwJ+IzSv01xa4zniKNRmtgs/Bma8uWJp82m
Wm7WwwvNuaWD+NlFgXIHtxtPUmrzdlkjGvT7zzyFTi/5jn80vVgXcbdD9L9ChKow
gEQGAFHipvdzs8jYps2a5bV+IoNAVoqKDiwFNDRBLln8wrZhvvlY7eSXg1jAda1T
Z9/CN8++rjXetjYPE5g7kw95b2fi4/bVJzIrd7i0qOyn660aL6XndwX4TuhC/7qx
vzwc/3z45MO2nPxLSEpkDg0/r4LExhKR6ji8fKvroxNnWFsNNVth0rzDuhOltVNI
YZ1dyUmCzbUQ7ILwrhIS7hbsT5p4qoVjjLn13t99KSdfcd+8tmRy3LblzXDaM06o
UbSIDbIsO2ppKCliRaBCc7IMziKgp+z3n78VSGWkuZD/7vogzVZYEC3x5prmckYV
vnWANzAidd+MESk8t3QV9wpCS53g0DYIh9yYvAj0Hvx3bSGVXE3f3nLejpofD+dZ
YIC9lYGMqEL9N+eYXgWf5slZPMUFSBAMrFn1bSipNFmFwwThYWz4gSlAcFITAD3i
uoxA4jqfE+9QFds3YFetCsxgsb5/E90JL9EWxBir/iQlef0AfAxIRgQXTx4ZcY6d
havgmNk5qO2wRpRMRPsAJijegvuYVn68PaHe94pD7AKJCb4vbdrxO6T7UzFmaXCL
F31l+rvBukxa5yr/YiQU4uqlgJrRrAHiJYzwlVHpRLVK1YnevHZOgjrJGXlvAeA+
pEFaYfbK7HrIO0mgY5h5hNlFJBB3HaTsQRrHtR9D4mQtiIonCpKS78z72Tgzmqc2
z330P2LGBZPbPjZG46jZX0mKeVT4MecB6nCJ4cZEUmZZ6KyfT2Ko8Qbx4Uc7KByM
t2BA6ldyqDhdLkS5HKODyHb+JzlzaKqChPkySTPez4JfCD6ZmicSjg29Mz2qOzuN
/7ZEj+QoNwQNKTX2E3FrjfCtyRITt9jjmThyHoMOYksj4055tNsvxxgF+kOD11q9
kyXkgXddjdlViPBqNaAEwMzyMDLlNwE91rGqJ9xoxfTCs6nM91bnXL3upzZlOzhH
GqVa6Lk0w4/zrSef3qtSMfdz2XkilUdamlt8MTdo3+bmRO6nA8e8zu6BnlGVL1+4
32aFcXzgtD2mDaZCj99otObOsL0XRgEnjwLcZ29OTY8anEnd1V6t1MnJQElF3qdD
Ke+syqszYUpwNl8pTIWPDOLjQB0z+2jPHuneXts8FlPd/GRsmgxG57N5q9UrQ2qs
0J71LMwqvEZMqMtJOs4G4LmSnqLO0517dfyAj6yoWaSSr/FicTpLOouRWtMkasfo
pwFIaA+Z65xlAoO7v68K0u5ldWvRg5v5q9IjBVb46f0EyFXXrBzllcyu1c4qrzrc
+sA0qz0oRnwwGlk/7CDjuz1mI3CX30iLgFXhOOoQc1O9+TH1SWZA/dmYdQmQQvaZ
JOhNfme1QG21wfxCziGk8xP2x1flh4xwcRqvUOCch8Yav1gFSMCa3ZbUhdyIFsPh
+CYLDijIsgBJ4sqM7s3KtLrpbep75ks/TlV11cb0std+z0WDofMSrIM71kMEsWZf
F1SP13NtBMZDXms4mCKxoVdGNKwLlwea4riAiut3X8kOe0DQi+cB9W+riXc6n93u
hMP0qBhP8EV75aRGXKwab1nMwxeV3U1QW51SdurKEi7CrF4OVWW5H4t17Z+X0/CS
SgH8HZ53Thz1ghveuBpmVd4qLUB8Yd7q52EZu0Qe51+0OUwTKrvBj+7Xgi2A6vO9
x2+cN+BuVrVzIEMQDXGhTi6p8y8CYmDL8kFi++aU5N9LoaAFKmQGoZtfCBDqa/E/
JaKSTE2znOd9E1WteuG0TOslJWYRoQRrbAb7/MLXBEIV88N9z0yaU/NSzQFTx1ru
1ToskQwegPLLgOJ4HcIMdix+GB2h/pK/iwzP3yXFBvyNkQIU3c0rLkB+2in58Lso
n4o4r0ywgkK2qSmW57UwWrapILRroDs4N5WcqkXxdELcEJ/Mwn7V9DtnXfOLGyBR
mtXcL/qOd9Ib57ytcOx/S4tcUB4iwd6MAkbxVMgiZfrL32uPGeSb8TIBWUbqFrYN
+G6lIVt3Cz3dR0QiImAubIvp4LSF9piaNRsJxbknxJ6dQcX7GuJK7uRusCiiIXNO
j2mDlZoiXw8uHf0RlrxX//t2YDTzNXXi1k0fRsX5SJYW2FWSpHt9pvhuCA/BCTSa
0n09lJiYy9GsKtNsywN/Ci5ridvsUz91tptnVqgxyFsmu+bthUqvzlm8itzMZY5A
wihukKrGaipTpa64GbYgDW9Townu142grUEcOZMK/8wwERw4u+1+xVAlOqcu5iGu
DibN2YUfRvFsLpMp1MUyd+B15B3X+tPP4Z8GIYuwVXG8jaWLBa5RMoA/nn8ymhAl
B/Obql2V+vfIVabjMjOOxSbU7RuORC0UswBrMCo9vPW/9+LoQl5OJw6dCJYK7cXc
zP0fvqnu7vgMIUEbfXjWjMXOmBW1oUVjnXeeQrz1c7GHsXPw+MJUc2ETwJpWMQ0M
Z/OoyV2zJNFk5OSf66VvIQOeigaUatRNfThAUVQuj6L4YXn0YNlPiW2e8+j9ezf5
Fqb43ntZVQhiIY60Cjod2qOwkTOVyjQ1Wg+2oJx0g+HEpyoc9cYPErntxhFTlk2X
VhsEXf/D0etATqDW/uNrNxSecIJXRuidO7Jo/E9+CjTo1kqTZwECkRw2oTTJPwe5
Szb6L8UsN2oKqMuCrTmJxyZUZ8rdjOTD1kG9sycLk2tnvfDNp0EnHvQ1+fCWeohx
ZuPEUf5JOLBaBg+fOWeIZic6YyEd+UoFqf/AI2QYb6wGGDjBpofFkcYcLDaUJmMm
R23MmA6GNjICViLd1dE63VsKiDQct9l3Luu/9hJJS4NYSZruVSge5gkl823TUuxf
vPnzFHOC1/I+8iYavtsGaMSxrShG1Jwzd559TosRzSxVacy8f/F2dk51klCtGKhN
ES/q/elzm4QXHroV4zQ/nMdgSxAXnHvoGQ9KPrKtFPU+83Qsr/ywnpDpLFPsopS2
wYuCiY3iXyRcFHuj2Bi4wa7tncads9VVLbfWKkB2Rmo3A38zOaHuG0tLPe4NKMux
oh1ny9vil6N9aSX5G8+HoC1hpuLKk8sK3mWaa7tsE69wTQ2kyKE/ozlJkFvrYJ2U
j8beF3CmhJxIn9Pqkuk8VlpoTJZnqh7AIX31V6k3Cepcz5PyGSJ49qv8iQZ7h6vA
TUnNCX3nxG3t6ss9rk/J9Pm4DBHqdDFOsyAYNuPHXka9WzEgc5zKMsitwPoEbF2t
XrIf5R5xpCMH0kIt8ZZ9JQhhfQggTGN9TwdgZ04ApdlmUx/QMDFVtiluEdWVlQXL
0LzRixzkH4ufjwrSY/hJQ8yJ8CEtJNhYY7QlOUMAC1hRMzNah5ww37YDYsyVQMU+
FLupvyV8EdIBg+X1SM5OZpUX6SLmSbGIFLUGjzZrB4sX20VijNp235OPX9LQKD+0
dXad+2WA8ogAwj+jWuIWccCXSxSaA5J4cAfgskRa8P55vMEU25VygNGEjxlGyssY
2gWe5gmOKg6+O0EOP9aAJ0SgaUebmo3+3FshX6KJnZjLIzDuEtqG2kNTnir/vHIU
RhuV83cO1hE97qtp8+3B4IbSr3SoTdL5Rb17TKisHxRye6iOLoAUwWcXz8cIA7Mb
LhZE9NzYgdtoa37ithkbBOP65iWBX4M2afFy2BL76I2zYWGjM+YO+PDKpkNSMa5V
P9SsWijbv9BuGKJCpdfgaJG4EPTNHdZZ/6YjA3R2eUpf6EVp1k8BFFJaInd4JGVb
2Uo3PNYF1411aSM/OjlNuivPgOofn1sXhhq3dbUhDo5ofXccsk5AoBkBsp+HHX3z
/0rOO83aotBIBL376oJDfobB/z0XcwsQMdwnKwyrloyKZR4MOF1Vu6fAjayCTonP
2g2gG3dEEIq7hB81mhcTBXGH/pMUee0LjSRz646Lr9jnmb23NYq6EEjtJPST/m9F
wBJe2XH7UheAOoJf+Jlw1eJ0VUccsiC9/fCh5BP5P+iStMHIQNBpOGt7aeKt8+1v
7/+pok/0nRIQnVCut8pmLJFmclPGDMfNd6wGWo+4OHrlJFiaCVfoDSrMrQseTnmb
2LZmNflEUHfvdaf63jchCXGEsJAqsFDPkygj4qZnpJE5BDWMVn/Hz+BMIeoY7mrb
OTGIIn82Hl4lJldQ0cFXyKM+xwMo0oMLzE796f0WYmIMyT0vsC3L9dD6c2+v0xlN
Nnzn4PDDjd2GkLOlHdO9IhhHpz6OFDlYnJ6yHOskAVQGB5vF//CdMhp2u0oI5rkY
Yn6z4uSYm28IRU5LuI9v5CeT7h5flvnR3DwHpYpJJ22eR/n8AxerrltOVFQTAZvc
V0BgQSucbk8GSggL5cx6IrVAfKIvWvMCM5JDbhubX1IAd1uZNqB2LseqczeTkCIv
bk48/41NgQlY5c6geJ8wNF3vOJuZ28MrOe/dDv6TOmGIGQva7ScyygiJTCM4gQQQ
fR3vTbme0/5/dIhev3ofLeUAm+5d6WKbF9DBBLbLunKpwiVrrCsw/eYM50IMTcnN
lZkRxinpU7WJfKQ5voK6f0sgrjk6Id1rmssW2sMM21EDHw1rknRL0G7QV+hPeoek
k7Vwf5O7WKh15egYqSXevcUFN/NKZnOkoBznb4cAA2SdMFMwCfGw3KRLF7adxh0p
YW1Ki4BvAgIcuRq8VrdLkKFxjaYyie/M797+nPpx77VCI33P/jQ9NFTbG9wz10tK
dDHxDn9jTMyjBeVCjIaemd4l+8+Bg59iF4awRuMf1nTzkKpSMUtr8+8j/2Vz8JO8
8krDlrLfrT+ho1b5IqIf5AOsjp3gRr2Rqd5rmhxdquu553pXtZ7dybIGtIxdy+C/
8iHjRuuRYBRI0QOobUcBz2spvAvTrI3wl0ZSziQvXuY/8LenzTXOWpwXGFOFt2LQ
t85GGaPnL3HAhZtCw/fvsnfzM0v24OkdidV6ixxV7ardo5YbhaKq6kEUOXYrhMpr
PviGqUAPXsd492RhyTjRJxTEfqN1pQaU4H6WBIKe+6r5Dlg8h3AeOkJPhCCDIK64
YjBstSFZG0x8Y4iBKnwnhmY0CcsPafMZnjxRT7FfJAdUdGNowghPDJVaO/2CLAHn
B6Ze9Lqr58MftWQHwoqc70FLBU+fCVFzFruhP8xnZqLPV7esylfodp8iWNrXSdzk
8zT4xP7ctYmFYTpDgmiunRsWd82ERNbINW1BSeV1hHY2hcvYWtpSQzxlKPb7EV1G
e6wofGUW/ub0TNXSYjd48UfgcPvfd+LbSAb1nP5OzbejlpZQIqLX6Va6psZg8nvb
uunl5mvdq7lf/qJRfjl7pZ7I2rb3h50Rl5fQNYVDBnE4NLOWtpdyrxuGfRXx7hol
YBDuu5SQIKD3xft7EWZ0a8puClTlEFWS24Xpclio6ZBsY2LPjUtN9kiBe1+wRFIY
69tP19lX52A8s4pbDpSVlgLx0ZdUHSE16IyJwMFrM84o7rB8ClUq4r99+C4EYHmi
KD0qTbbyAElAtIgAqHqWRtaNybP9fj2+QZKnDg0m/JUdD46UwmmpDA22qQdCrB6V
6RfllIKnEqSBYPQFjVcygBP9r0cywwEoMQAkJt9qr5sI7o6LnKwkDNPQqi+zLAMV
/f4x4eeT+klOL75GiGsJGCAWhXlMUWb2giG47Dy/52aEh6ijBuUVWUP2lq9cl0Y+
mAM0tOp8KniIa5PembFeaDuVPiusEkZVTND3fII5dyr8zerV0iMxWDvzTPxGYpMd
UnhJ1P1PO2QhCXUW1r7NlWF3PIaFa8/ci50eCny/oF4rlOFUe+32cNN0VfMQBZ3K
HmSRxrZK6R7k5PNd1O6jUkaG5U4Cj8FKoxODuIwiSKWFH3Nevv/OARySf0n2mvga
bryREqg92+GRZLfQJTUB1CV+KOQH4j3Llgi5XoGOdP3uwEdy0xDxK/R8RyUXGTYo
TopeEkqVFyg/5bN1C0q4WqnrTqjAMCJXqXHe1me0q3tTPrv8yVY7y6PS1XvY9wnq
tlGJYFJ/wokUOtVk2dpqWO/D34nydhwuuQKuyG9VL80f5kFrKDH3mzX/M9kjyg+z
zX5hq5+6LOlKJDTywyNi0H4cLo+hDtZZ4YVlbJ93VAeqnb7tNGktuVDDSPWE/49E
5COHFpe0aCGg+NWjsyLFXw+85eLEyX1pW6uZNsyBSrdPpfEjksazrXe5UCfis+tw
HJQ5rumeNCiz45NdaIyHjOGjTz4GcfAw/6jlKuR8/LB677NuuE4Bbx/THi/ov4JW
qT1dJl9U/4o2Bok3CO1YUJPeMnR5Lftm0PIYIPl2Tmv3/Mgw1U0WmQ/8NmRzZ884
CKGouKzdlLnAfdD1qBg/X0gHpD4wd+zZTgBkOt3HYvsl1nIBMukOliv9qm8V7tFC
CMvtNA8nAoGz4FU44fTd2LAFIfmJTQuoC5xH50jWuC6Rli0uvS9bFG5b/a1ta2Da
lwDx51KOEsFGbRNhD4LLWH8WBNDo/aYj8eRJH3XLXo2l3xn7H+3SfMliAFFtegaD
gV3wDgks8PYhqLeEbesHnTzt3APWQGprEhS6fOug1qDqTZZyP7S/nzFn8mPKxDlV
TqZ+Bgabp+JenEQCaaJIBRhi6eWL5OxXGt4wCw/tnW5Z6mSGpYD8y3tGSlipwdIi
7LTkziOmwfrwtZA0VSElPkyfy2ws9+mbxbuus65ItTHeQ0UfyJyS/I8Rru+daQFT
R5WvObzz6s4iJ4X8BRwD0ezdECmUeeYXo6jZ3cVy/ilR3dvERHZ+6H+QAITQsVEE
UuPoJ4EQjnL6zqJFqi9cPVJhPopL3leW4jH1bvNf6unDv8RmAjoifZLbKyO2fiKM
Ssh6tEHdddcQhY4nI7vtTYalkleFFDX19QT+Zk8914Pgc5+/FGUh3Kt8W01HK1Vw
pjxBFaGvDOjAezqbEtOpmcFrOVk7fba+3y2rKtBXelDNWhbzyKupYn6yRdLwOvNz
7Z8XDzNfowoMVE+gPwLjfJuMNIi8GlPFE8YdzUY30ZvNkUVU56e6HqNz5TPnSXE1
ylNph9PJ5k7y83S2RcwI1/UDD4dvbVE5swYFdrF/7U3yqMMnCiMhFiN08yzksgc+
zZRZXxj6bFwfiqpb+u3xDBpAdeoPr/aTHNdrs5Uknvepr+MR5wKItamSPiqWlOmn
tFHXJbKv060w0tT/h+AdthLMxRLIDPfYQ47ZKZDTnxo9UayDbHj3hYQhOJJzVQoA
JEIvMsECNzrJH2wY4wWO6ej38nm3DAzmeHyvL7DoagLN+rhu42d3owF3GM+waG8c
3Unp/vCqxx9vz7fzed0IEeGbVBdPGxEzQc5AoGnl8I8tYSHTKvAa/a8081n+e/uX
pNFtt3eD0y6Cza4gJExJK76BGpCHP7g/KQpF2KDZzHWsR/JMyAfD6glZMxNJCAZB
I5u67pedYzfO/qsd8eCEt5NS+QvvaXE4p1XfAlyqliduNfYBd2lJVQGi9vdNp3An
reRsaV957UzRdCzjs4chxIcm6xGPgLt1GYKcdbR9J0VImmWnrA+EbcHDTsuFqsdw
RNt+ULmA9zm9/K6RthOOBBm8beh6FQxAZ+noJOn8xbi14QRqJF1w3tNESX/q2Mvs
csFvAM6LYRW5z3fC0PpMWv+j1d8Dc38od0xdm1ZXrXWYnsaJH6DPQhtNS259t0AB
stvwohIhHbCveyIS6WtIiMNpCB0KPWlxJrJQIc7lzGDirNOjT0Z+eoD0cL3Nemor
zVYF7qHv9NAtToqR28NsNAq7MCAGBuGhsheVgfZVkMloAQVBr/5w40aRpjPBx6/5
E426LVAmByB3SivniRA0x4MbSLLlm9gFxjFDKInk1yfad8Jdc0ko8zhM6bR2OqUb
5dkdj/2ZRJqo18yzPe6foartH1A8MSGlj5mtGSAEpmjLM/meCiBuI4wAVXP2aseM
osJJaAm10pUnBuOxGNZQvt0EHvZu42VWe2rl8RcJWzaMLkioxepCbuJTXmDtZe8q
MotPVTvWYrFjTPb9L/50Alr+iGoz3yvTCKEIlBLGkVTHwf4BQ73lcKIl7d6QU1WM
4MJFFCcR8nFIHimwEBgzZWGi59GlLHYowvjITM3m+5uJV5iuGmXSkBQRocFeMf/Y
7DWIa1tCC0DLHXcVP0Azr1q8O5Y37rZUh4PDiquoGaaiJw2lW1R3pn34BkZq1uw0
XBxNdIn6gIwGheyFgP7hiiUA6cC9XaX0BmrJmFNtpVLSj9pz5B1Wp6eU3PvlPULf
ttA3to9x/yQvLHFKwpZzsfi6saEl/VkkN30bZJlZLJ3S6SuGOOAHKzeYoZ5XacaZ
QATCEan6ICa1l3V9mcdotBBut92JAlw161B8oTScQVfiGVtWEBUxTZVWpc8SL/Sn
s1YVMKl5OxDpxbgIfEeKmOAoHGZRGVL1GJS/Nb+pihT7mkrXvS+P4ckZPgRT3LCT
ve3VprPEVUOQJDqn3fN4LTYvWpov6s/lHZpTfokTL+4XHIIpl7LzaOvRshymh2kB
fvJ/gW9fKizNzFPsZyi6Ib3MCcFpQyfo1uPB3FLxEaQTWWsUug6WNjK6GNx+IKlF
aVTr8djp0xouYH87cAqhY4xPJhy8/gZpaOzo5gJn0eqrqnLQLLw961M0FSwnrG01
TGwz6L+9O70h9N7TcM/75ynkeDHp2vw0hM1Qv/Rl/xQi9+GS2mF23dCRr4bDpRXk
KxWPHeqsJcRrdOxqmszVjIhN1QSEz6DjpYwuH6bnflTdPw5bQqshpxCBrXtR23wK
D02V0mMYHAncQYRaMdWNrwbHP0YOsFtZq1bQzuULVUyVubimYujaQDNRZpGXu6WC
X8c4ngFV8EVgtjDjiDjKkdjyGJAZvHhHkBS9ZV61cgVsAaUA2zzSxKPceFrrHXEt
G91u45qvjcDjPwHmgT1OuhJEsdpCItW0MGvWuC59Z6p2nHbvgltzTgc3p17q4Onc
LNvmtCBag7VwdqzFO90/JN4etgaTu17HzcFdgLuE27oFDQgc+JcichACEEAK1nV4
mfkoShoaKA4AkSdl43QPIOUwEdDF+P1wueOvQKWNoJVoK5xSQdZvUOMq+qnag6Dd
0zeKDl+LqpE0nsXla9otm/zKiLfAdVQm017yKzGzDPTF6rQMcTIo5p1sVYMrchy2
t/y2H97WaL2b2025eId+3Nkjubxumb/++Owbu4fHAR4umrq3dojCDkjbrG6cM9t6
R1TtJgD1LAb0pZHoopnTMSwWUt1d9kCdSw55DEL9CHTRb6SlE1qOdALa6/pOtDTZ
Wq6lpp6JmCWwaWddlpWp8PW1MgBZOavZP5yBoinXjOUTLenrrQTJZjwUbQZjJ2c0
i0qn50CdT6oSI2SH6nDEUHqSsdAKrqv5ja45DJaw/sZEu8aGq7gilF7E5hmdUJm5
Qc/8rh7pOowNEEq73mAKoac0RCmjYoLTDOeYuwRW8eirgX//D38mZ9Lh9A48OWLO
zmxFLE4Hxj8m86BohqRu0wbpnW52P+5LSfjPrussUIIsMvw0RzQSXbMDZxEtbVR7
ug8QUSEty/qZlKodI5Vn9SKqSeG/T412rQsoREVm98PGk8Hl3fz4hsN9Kjqf+e6n
FlGFTqXu15twB3+d5qNntqpf0pBk9Cgb+bkqrW2Ui3Sjj+Ryjj/d85slTslQ+dvN
1wDCWrgBLwhtlbpxLH7mVgV/yU6StZKkSwy1m7Yfu5PYYTziVxwEtdCcZEssnydm
S7C242SMY8ow3rXEmuZ9QykIHtXbxtFYQxxy9zHFfLG8DuvVVUXvBK5ZPeN2w54N
QzupFyD7jsfNOfjGXX32TrTbD+CMmrna2dhTI3hGROzTUY0i3FrMaH5YIPujRiJy
f/iF10rx2EeQDq9buJSPrI01umerrTgVxFFPTZirMFC6U+IpaYUxsnZp6KHH7oAc
BfB9U02Lcw8LM5JAfNKIzc9mFvA0TftWYA1YCb7C/uvP5fDD4J6qW0GRkBMIsDjI
jiq/Xkk1Y61KAbRbqo/RQgBZIAJd9q8jq9JvPxwILd8Q1ALOi/7jnsx/+OPoRs3s
kjqi5ogWpi5qAw87KidGNhe1sMbjHOFtp78ysCks4EiFCEYj4QDHYVSNUGdcLhWx
lCz8vdKjpv9RWHe/nrOH8I9hUMdK58f1NIYOzTbYY8uNuUuOubO9wzrFldRrwrnw
6yB5WDQGm3mgbsAFDKiUPuxCVtHz8Q/5/k0diAUwL/hs7IB/2aKbb0kDXPbXc5Kz
m9N87hQu7QD/rF/wT0aGFpdEgnwQlv4MiNYq8wu5l0rOxQijxZIlYaFpR7KaM+yR
dU3k/wpfcbQ4yXd5aiSs4I8E2rACWG0LL8diWpgexbqVN54cZQ9WCXCn0suGb1um
Jro9zc+cj1HqqO2eezYRAAUWBM4/F0tbx3wxNZaF44pebmm8SSpKu3kYXY13X/rj
pwV96cmSGlObR+lyPlwNKTy8952StIKRwCloLGGBlLXmF06AaW4c2jkVErT2nV9N
3228Q5El9hQBuur7jQp/jQDrWgM9aI56ulHXZC//as/ZheroHJ/whiGZcypIb/8d
99DJbVjmxz1wttFsz3gUzSCDI3AvzbMZq8SDaIGV2a35Kaz75hk0E5Vfc1WpOCff
7SeYPuoUqZJVyOkP30rpFpVe0puMNCQw2Uk87y12V1IgcrWIKnY45ShRWc31ZtNt
YAS8yQWQL6QhcYwBRAwbCxPLjkqSq+GJQfNOle01nPS/ivnHeDDYbiAuOKIKY/vb
KR6FJPgkJBvZAgKUf3LVN8RG/IN4t3nISylJQEsD7pKZCRiEB9WhgXIGeRjaGHTr
03h2zHzZsoytze8mi0qiIu96gyc4HXFCDv4onqlAKEv1UC7BY4VI08S9QL5Kvrfi
n+LmvPcAJJRrnXSJU6cX6csN/rzOj4GBpCxpdEN24yk=
`pragma protect end_protected
