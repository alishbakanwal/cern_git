// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:11 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
H93uvmT3bTxaOOota3MWesSP6FDKZJGqq9IuHc8XOVCGiEItWsySf/gApMq2cW3k
ZIzdG+6jBNaNm4YAy1podRjVT/r1ZZa/m+wWS73/1c8jv1tQbp0oRamEaMps1pUM
qvzTL23s2MWpvbP6wSbR9NevwqTrWpHvfBQt91jkKAI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18368)
Tx8ib38hMegcsKMOi/qaUrjMDgcVQySYP2RJbQI2JXQpvSI4+s8/gnYi3ulegZGD
QLjUgJ4BJ1St98uF2Brya+lWOzKOf9ZOI7a0PDzg4ScchZPcN2eGoxwzIjQ/9HpG
21l8r+X4ksrvHRqCqFjI605kqhBfAsgyZ52GwA0Ru0RKzPwfTDMDUf0ELEE+8fap
dFxgHiGLddIeeDRxGhenF8oSlapC4+2Xzi2h+X7qYoSd+go3xy0KS8/P/Ou94gEF
UBHg5qvj6rJReYCq5t6LG74TqRXtU7+TtAm9Axc57dZG+SgbseTmM8jsSLVigA1S
Q0WY8LaEooYujIXcfRKQM6WHUmooBXMB3ENUrd37wkRBlKHNKLIyhpITlUQiBnAp
WNgX+7kI4evvVVFNO/UyVW06tPMMmE8adTZOHtikCtM7dWCV5z/4yvLlzSnQmWEA
hiIaSgB9K4kdRcwiTuLeTPxnaixmUMtbkVnRbEGshwhT+8yWFS+y9+gO6Q7+tOKS
mluCee7J6QfiDuh+UPau9LvYd76O6Ejl9Z4lT0k8ug3qswrT1nKeJEyBZt3roAsa
D08BguYVt91CocsyPCuQQOKmyqRJVpCV99gjwlt3JdWmuEs/Y2xFZ63pBRu0Ojyt
rjwgoiHBZJntPYSoOgjwYw3mkow4j47gXEziUZgSCbis1cXYRLDdRfT7FSvCALjm
uELGkVdFa6gT3QweC/OVMjLE1b6qmyKzHFi83KXuS/96IMsdMtlRz6SbQexWO3En
80C4SBqlMRablzERCqOcHFfDX232nd0x0wo8yQotPHzo4+aZXlioCyAuRpmmzzpG
RScRuXctN3wbKWyzrzdiINcIXB0z6rZ/rH+iywT4nYr7YrqOrA2KQnLYQZXf2Hm8
CQ2cKW7XwRv08EDJEMUzaemSE7W8ONqrmMe4C97c8zHqnQTfr3ROBirwEDOzhqth
hFY1ponckoHEhJJR5lPGS5I9sRe2WWD1Htq6RymcnysyBIlr09K/F62eX3VOuihZ
QYnSTbL2aekNsDxZI7z6kLxcveltJorDE1IPtCc4ZYajnBLGQsoIWTMutfsQ+loa
MUh+ZJ7VhzliI7VhFWLUQGxRqGsLmvFUbeF3vU1DRRKYWELzYwGwVfI7GwDU3nbH
UNQRl0FXA4mAepeQkmSh4VFvcSC1q+qEU6hC26b5HF7RLxCgi1bC/V5xrzX2nr/X
GnMhh4EJ3lJyNTN07GavlNU5ktnBikjDo3l0xFv5q7+251JNeqbUOK2+GehjJuLK
D4eGycxVrCxZk1KmF4MPm5b4YyYYm6uEmvP2HuH1eviIzskrmlSk9ZMCSjEwwI+l
hmd0KKXxhkz+BQlxnMirmIKYb1m2kDJKyjnUrlRFCVIGhucUR7SM5/RhYe1L67SB
A3dWWPIG3N6LpkcoQOhrU1pY2yCVYcouVaEDZ3A7+/2474iVYqhfsfLCV7ONBNaH
Qvn1UyMn2GPWF7Te+fjIgTNzK0Iz9mmhA5DI5OIn4dCQuS/CqaOITvJDRu0cxWK2
wBMcAiUe7nSpD8X1Af2uPBtqM+BZXr27VO02BwuwIfaC4F25DaOELGRAAwk01P0z
vPjXBMkH31vWln6NdTZOyPaMuS83CtzZfYf062Rfe8V/BLyTZycHfSzOEO3Lstsu
DAikRG3t7D/6751V0wKMGhINl8YT3l5mJIGdtdcKtMlMjbfESCI3a4PTe3svfwbO
kquWcAVbhZnyAFjC4dG2TZDUB1MGKSiXfKdubHLE/SpjvQrjB7RjYfLBo/xLA0WH
MWPhDpL2zCWrFFUs1oqlS/uzNiXCr9cRJJPJag6ZvXsQvQlZMAbajg5VCBkb6+ts
m2omrnL+rgVsHz2BAkjxIuaXFcNaMGHiIgT5LrtdKFo1VHHnIVi1B4cyk1Xgvvqp
bMSsB6dsiQctLcu4cvXN6gCZsodye3Wt7k06NxgOTiqbVvt+okh6ePMjH9RbSeJY
LB0/XItgf7I7ziB94Qtn8g12NjICTxH0oat/K2hEHpen9xqGInUPuREYjOoHD92c
ZBS3tH798K1ptw0RraE0VYzZhgipYqe7qpJc7yM+/wS7eAai1573TnyT7wOMhhgh
0NjUKtkywxZQXC+vREKCJd8SD7KBFJdQaW4MBUiN0hrpXAYo4dQTcVTGvtNI29v6
wG8IdXizv2En7wfJB0x2ycxw+etxTPSo9oaEcUiNWPxKI4qm1WiG98H2Y5yLFo8b
hc9XrP0Ry/UxqnRA11Dh2/RvBHNNfZ48Py60NnPONC5zfBWrhkWGAvzNuQkFUZv2
yRFPQe7X4avz91ZIw1HqB9/wfr+dY/9DnD4bShGpxuVoCFBOkTeMVY5gOFYlqqo2
6sCBRTBdXbi9uxIt/SL1bWcocUmM3gPgjaVIR0rH6sFiNYMQfpbsp/71N3V8XlRC
gNsw9MA9yRG05crVXQt1DSX3xKWd5Kxw5FFYZ5373AHvN+DmRC2x1mN/v21N7i1/
fAq7NfYSg3ojKo9KBRKeVhPdsHsDFPXavxNAFDvELw5UBPJTS7QzvgZ6CmK40X/D
cDTUjqGHtJndHF2YY+38tYsYmgzsWmVp8OYOXmVBLEUkL2FRdSj3EE3YCAMGMLLI
NtUSy1K/muH9nzNiiYrtlZdvi8DTL9zJzrZLLBeaKEJCCT17TeqZ5EFH83R5F80n
3Iv7Ojb7vRykqBompWIORhCgnLl41NC1lrKdaZJcvEA/QVCyrU0P3mzBq7l9czun
5aWodbZl3n0+BKEDzYDiwN1UVzwpaYltxSdpDdGv20cCzSklXulRU4TBHX+HsQSl
odyI7rdxK1NPQS51LoP5qL2m/41RWEFoZSSbNe+hsWosVQeFOxhcO2mGUsZfuRsS
/AbvxszMP1R0yk8LUhpbLp+P9kKb3XqT54TvPsBAKnkqBSrtveV+1BIqg4g7NoRK
ASViKqlIMzinZTtXiCKfYPOWs3JA4MgtWPQhswoCM6x61ypEmNKcwL4C9hR8H4g8
EE/iguxNI/mgpOK5NdipsI1ThUt0kplvjnaddWh3WAP3z0aSjWGx0RVChTHD8rRA
4MQc2NJvT/j7nRgP3i6MvEpsdV+B4dSYm/GDyfTUsEuSmwnxArH1vNhcT0wabvFR
dFLKHVcmrFuyAe/BLbSeG7uOIgUpJzDrtCplXikakF3xHRBI94MJOpR+24v3ylCV
XA7ucfar11ycWdqGcVqNkFzkF+oOSM3+cEhwUt/Eab098XvmAfP6Q6u+W9cQG17c
3kuSREkObh/MO/L+DBXQTCn6lXGwdp2oyto2ctNpbJddv0Al+tvi9qaWUoWEHGNI
QnbyFiPWf1NmcaQ0umiWwV4dDF0544TLozBcGi9XzKiX4r23Os1PbqtPjuksnWON
kTw4oZABQN52yOunPGU9WNJOXABNfKstaDgSqmQAgoieN+ohLJtZH+XDcXJ7dzFH
/oZ4YPxMfnbMdUBB4bGa4j1JdPkDfZi/EKPDmH804OCFX1GrXBt4t4wip8X1JWEq
jNpMyiZsPx5Ce8vZnotn5I+wCNxW+A0cRin7WbyaJnvZ4+Ui/BFoieDQUvXGdWm0
FPkkJ+/oMfgz2DMl7h7gxHLI7rirgB4028aF3p8C5lPQ0lOgrKBicDv33SV2tes7
14/PVzsGf4pmmgO2l7+7NJwgDYGN8SDHKhwkXMenoBbSyNZuTgTqQyVwnbvTMhAA
L1qlTG/xt6mcCq3vbnvP7XHy5fScMJxciQUoisBZmHo1eTx8dLxj9OJi/klEcafa
Q9qGPnZcLHLFWSUQQYizyXivEjweqn3/Zs5/xlkgZT+NOBkW+9BPxQfLLgiZO01x
R17ymCeruiWlH+R256cgKA5nB+htFUMthLvQ9saJmqR5/LTbm5XI9qTb/c+phZte
4qKBxcS85vzD4ED6cXW9K8ATrmuo2Fxp9E7U8bE8Ajejde1fTdliD9VNlUrCtZU5
1oOeXgxAyX5QChi/9o5zGr6ysAK9Jm218HD4dtP4oElmERBQl0iqR9uu+2vmwKZF
KFfrdwo07sRYB1MHorngeJwtsaoEi1aNgW0YI6U133/G6iE4VsjAngn8N/aEB6DR
UvOTRK2eaRSUAS/SZQJYxekzjVHAtdd9w+IySUOVkqANJbY/ys51DQmv410NsMQv
yBvHeZR37UB4rvIDabt12WztmZJHzkTEHEBR0vQYnu2nlbZltpLGxp2lPuBDR0YV
nMXDnDN/1PjaCP3l5GfhgB70E9LvYfiiIfbHA1ESGGy3EQVbvbDcqo6+FJRHZvn+
tf4084+ANhUBFw463lDfnRCUpddDqEyFdTNWdrjRw9KbvnBmPBZ49C/0YbXVDyu0
CZP4HRlwgCaghFpbkncG82xpkqkw81qnA0pbDYEe5+ri/HvuzAD2I2wGLMVM/1WW
hIeVh3mThkxJ2oDyWKtcAUO+KdD3MVhZ6Az2YQtHgnsrZY2zW2fS0puJvOzOi+81
SkW01mc2fHfV7/wCQtQLN4dP8sdmGrcxOKRIM9DZTyElwjrLLIbB0CfxHEl9uIR/
UZQGXWgaPOXBSXcxpbsC+Wh91MV2+/oI+/QFCAZSIfok5dKP4o/UKgmmDu6Q/Raw
PEwGIrpfRsP3txJZPxic2qn38dM34Cdd2ft8YHh7VTRa4B6smFI1HeeSwdR2T6TI
SRpuat+5y84f/xAtEDYUAYpC8UqcXVHdjQhreehSDaoyGjzV48fg2m4KUnVbwvfZ
UWFa69j1nk0n2p8X5blpZ4tPT1o+OUoJy+pvoueILxuecN5gc0CH1ayZYou6TLiz
AK62gNaxA58bnBnCCttwSSTWODZrfh0ejfS8bus6P/jNFOrojhI3LTZP0zxc/b4m
waCOrNLvFEEW/Vk6I+4uGFWveY/4KdSXjJUhTCURIR/No1qu49+3jgT3l0id34YN
pm8nYYVPx2rxJa/Utlx2UqN8gay32RRhFFbkThne9ffuplFtJqsGxiscOmwcw/Wy
g2zASer5Kj87g/QFbaVhkNzK+AV6pkNPasigs9Ff6/s0K/oOB41NgimY5OK2khrX
TEgHUOuK2f/ONwfl/Ui89H2KJt5O68DlsYGAZRwk1fGv9eYeDc4NUeOMZvo7msFB
WidlwneAXKlqVGJ9yKk+Km6UGnw9563UDhQ9ZN2Ry4btH12ceDysR+PgWuU8rUA+
t0MP3j7NJkSX+H0oy7o1CJXtS02z2BTVQa49vbWGq5i3vCjuR/YO88WPRM0T/K88
05IxrfWZ9FemtCxpllUN6bL5U9UZ+KerBQ2AI+yeuYVaHVXjeyqv8auu66U4LDNP
F4dfPKBp99om4Q+rYCn7Ay5A1ZnscHt3daZUIMIz53irCUuoj1u151Xr2eru2+OY
IaqMjSSr36wezXw3cMoyxirOeuZPshh86FibOYq3TaxcUReK4cXAI59sH0HVy4Re
NTVqX70ufQ3sGf7pjtp0mctfT/SmHHOfZx34Rk/Iawr2gKwfvk4YAVodhFZUs3w5
7RGku+jmZF4EgwAHxW0y4u4Y4Zmc6ohhz07gsVQfKPxvlZalpGVm6Ce4EUoO1iO5
VgzMZDhJlHI1Cw8H5XktaP2W+oPZBTp3b6K5ZnZZopxBPEK7mKJEqrWWmpJhEqg+
z7PMz7O12hunELNRFBQQTAUoenmo/97WAv6FmKMTrxIkc6m1l9py7DkrsAy82mni
BbL97MOreGeMSVFdPElS9yvsAly2fEqNbb5kq57s+xbB6cxceD5+icjdQi6ikUyW
ORNOoZx9ondAW5S3igf7CE6DTuC7RtDkzrwz7jZXdHrnnfRzhNCRKEKN57oVU9Aj
aJcowjnypCvNlVJQPka9Cbz91faqeTFdeUeZHJqBnUYnen6DGlHRQ6XoSqtVY5D1
djpobGxHWmxZ2PXMkkyuyUjhWO+HvBXRsPZ1xVlR9lvPLhAlvu+KAWmuGFmtuD10
EjkkvDaZD/1xPueYiFrtDhI5FWoEffCkEKKRlt7qhQ5qxxaiXSHyh7J9fGAMeIyX
IkEXT0cHywkziKoFrNL5R+fX5KVpKmwRdX8HLyLGHtR3GJ36mlU+UgqFpZYKKaES
BJ4fRMmQ0612j50K4vl23w0+tA0z8zZsyxdlXVr5OALJyWf42w7DIfXZ0SEtzBHd
i2gSwW7AyJblN0ECJ1Nz9j/Ra0/WUrVdf+AAMFpW+VR/kExCEyH0G6dKXEPfoChK
MghskMoWph3t1pcyu+ErMIHOtvQd0rtFE0Q3jkm1bBbTxGZMhZlHNm95h9RtD2x8
4/wJb+HwPgk3ZbqgMpi8G09m8kClqNC3M3quUcdcZ7Zj70lsZPHr1DIbQiPW5CoY
udjJfe96sR5z8VZ8wfN3RQzXEBZEfYnfX4zgyhjEASRWm9vppEzTUpe3P0GI3Lem
LO3D7kdNNg2RI4QTHzvM/hkHGUJs6FmqmkwkySQwkvJN9Sxld92HTA8bWW5dc/Si
p36SwLekNjesUfm/iKhYs/SCPpjyHZynWZ7HIHsXZrN8P7j/wGzLtaTgbu1vT6A7
mGJdE8A8a0H/ZCagND2/oNnTyay1+KUiWFBdb/KEz4KFq31lghz9HhsCVXaMX3EH
bl3vBjamNnxT/G9ucghkB1ofH860BWzIr4anww2evwNcMMl9Du3HSkQogdf6tOyw
Wcrjy3WNtnrHyi4AjXGQwCcalW/7zEcTTtGmGaJ0mwlK2NnfUfSD4lYeHdvbYoKM
Kr2BfNpL7XHwZagaG8zdoHpi3Mlj6G0Xd0m1s9OOWMUdmIZ3gQ1YCK+QdRyfLppU
kbNd5rTQfWmxI6G6tc6vy7Tb6mlG6dnXibPZgR2594IOSKLk7HpnBj6hjEbgESra
ayUhb3w0Y7e601/6VFbac8JvqQ2q/7m2AZ220hLXaVdRg1Q7sIWl6abUP0TQMXkn
LYnuJJjbkdwEUFnKoKGz/YSNXxpcqd+oJGg4mZ/MgENwLjePrCJtSBxFxm45EQyX
QfHhxksbmixqPqMHF1SQ4k8wIFgnjqrBfNCcxbiOlTOi9vNYZvmlEA0jT+I+gzRy
Ri7nhxJWefLH2R2xbDmU+wjCjhCJwgjczU6ppSD2bgbvWMMhaCf+UmiBaGHabL+v
Tk/XLLFPfaZiMd1TOcJBCrezlHB9J5Z0zE1dHf5m/8qUnuk2VMovHoDNi0z998Ly
vn0hI/n9qn+FRRcB+IKY5/7lu4On4k35FhU45gqkAwkPZzfe5BRhfI9ETK+z4/zv
naKBK9+lKlAKTNNw0bH1B76dlGlc8+0Fq7ic+19erNKdAbZ5OuHQ4eZ0AtW+5o2Q
kZseiHNFggDEwsJKGD/NqHFdT7ZNLVBK4lUhzjJBV2U0MK4cIWxFximHyxaQIOuS
c69ywypmupWyTQDGZdGeFamdheiGt3S0Ad+ilVhXbxLC8FiYgZVOS65u0oAWqeoX
hcEOhpABDo7Rfpx/VE7C7AYu/6FXgWSuyY554rIaqFSpxg2U4dGAyZ+RHGun0Hh5
2MC+lcuzA9ocpQqVIT2GMlhQFi4yox8nqGwCR0wHc+gKm8GygRh7tdzA7LFc5XEM
AJNXbAkikdSszJMlSg7sP2wEv9Pqsx7OaIkAVWgeD3P8t1+Nr2Gu+9D6PJMQ/Wf1
uQ+K7ariE7VhlrUhmXUcxz2aGhFkxIbbcohXyLxPFY+GxFPrd41xVE88XhaVtJ0l
fx5UYo6swuiPgnRxwugfpnN/WvcdnKdTllaZ9fL/Bg1k/DwFCSSSxDYKbq0+Xor1
TwVW/PQV4V9YEV6lf9h+2fqIvPLw9AqtwWvDKomcsLMEuI4e6FzWOvHzHCwyztLE
tvu5vkRhBgO0DJegxlUXDgontJgEMLR8f3U//M37EuiVSTwXRJKfOlzl3wQe5vLo
iDus62zGrvwKbvLSlgVVCjS1Ep8kHlLtFFaO0r+j6bAKyMSS5WpkotU2YTKZVxKu
IMkk6We+ClO4x3mX1NkcqBB0WaqGVaeUAhhk/dyhSRu/dPT+PWC9zHqknUshT9iz
PM/3FWx48tgFtGXuoWCnaVmKOt6T0AyZjim28SAJole2mXzAveyr7GytVzsURlzD
WkRr5MMI25foVEJzO/PuDTiQ4PmPMBKLq64+nIZj42fJyxpwTnww5D4YOwbPUyCb
Zi7NIQLXwet9Ax65OJ3TCGHonbdisOVRpeceJDd9EcPYHguNKOymjpHQ2m77RTJJ
yQ0fyBmkEI3mwXGt1sASqsamGQrs1t9bWwrW4biHdyt8e3izcQA0rqr5+U9Lm2m0
raftx4tqxNFe3S8MgwsVJL18zP/bgbvJ6/K/R55/ImgrXtyyBY6HPG8CDAe3hHQI
EmDNsnbvUS4zwN1oGuIboBCs+DJrjlaDlEOOhW02IVJTPyHgq0BjBC9+P9CbUpHh
ejJ567bup+jtyK1RQxnif5+dU4PIp1PW2mCgDbiY1l0xfKZBX4zaPqB3XEj6FuMx
n7JO+YNesTDYMfG24wr8tJwfBqGP7ksTLU05zaDFSIiCCDiEiwcjSeVpQ4w1RNEK
IrSJ0eFnVqcZrw4HanGRyF0FkmtUo/f4S6ZbQCnUjn3K0vF063vgNfv8LK91ksSb
ll/ncjQupGQGIGmhJrMMbvau8F+EHWVxHvHONKI94L+jCHneug+QCXU8ibIw0PO/
ZuXAYEv7ngHb3b8iij4L0BVN7BdnC7tWbDhBhVhQ2zcXKGtZx1qFanh0H5r2Sk/2
ytimrvJU8xYfgYz296ND2LwfK5LOGHmimdQqeK1XYxBy0All6u8HwX+hzB7+WT6d
Osbe8F73vNOkp+RLG1rFJhLFrDwWVAG8pTNa4vAsQSLza2J/atvDrZr/hyUzF4sf
FCGlCLC9zXBCUDiK0IfRD8gVlmqWi8Fdj+EOoSGgqGncaMANgOK03+lcncJgmGMh
eqkb7S1+GL5zhC4yhainuxJiuBvhdjWjDziFbzNE3Dw+mXty4XUpBiS58Fl56STK
NVFkGPsICxs0Ndf/AeaMz28J/33I//yHWZJce+ph44sxgzLAwNQJwn53BClYrmgl
43mltI1XZrwHJYTt1JiuVbn93gDGkO9urITaBeIcu84ypjClyOOAfDXuCAZat28t
XRf0RdAHwyqjBxf87CXfKilyxcxxSKX6S5cmfE5ltAaQ5kj+4eJz6pPdxjz10HGL
scrMi+I+r5ENwNH1QDk7gP8nOlqAJ/q1cAJTaQsZ72rIvlvoO4I4efBf8IeWpUrM
ohIJkaS7eb+vo91Agrf/VBYdBhuV+nKEZuM1ZR0Ot+KQXJBqlUqv8ItBR15QrEB7
nG8P3nQUP5052vOWZSA8lTpkdIF3rjYrIrRrfnhMGtVqnK9ltN+bryIn4bNjEdnf
EP5dWqP5ZxaHSTf5cUYYg5nwsoJLqKyi4KbzuecaQVUfSwHoXgx1c5n4r3HsIbiD
gfDeb3nx6IH3vbRy/MUIV0AVBzIOJ4TM3wvnf8OYQA+WOrWeW2mqQlIWXUmyfDuF
GVooDecuQAmeAgWk10QqVcrHNtWauTaQMMKmttT7B4tmm6mVE8j32LGFi0mP1ofG
prH1rtN8WOYuOq2aaQ9mqmgWLIDpvxOEg4Fzz3BOFHLgMoiV7pHPw8k74OlaWuZ+
VU7w762kuZsRBRukRFk+ZyCoJd/ouuKLerhfqrVaf88+gex9+F9klIAK9ejrdbL5
uPz+JZY5T93nNxyNODW5QgxItxEix9p4LF3LzAkIMgRKPXlrTZx3Rj0N05F7WDMZ
FMIgmqpt2dkpBqJfknG8XMtX+sJbMYLGgJGVqATimokIYf2wwzTlkeeX/+I4O3w5
0W9Rz/0DD+aGnrli0zgddCiRNzi2XRX2du5nQoBkE6EQzt03wbqQ9kdzKsZpq8ea
MfEYVK3/7u7/3FJDo4STdAWJEPMBi/m5hi4jScpJieqmgFjNXf8wx5zPI/h+TvnK
XeHYD3nLBLbyn0jAzBjjRJm+rmQBCHfj+hlNP4e2510OwRzJ4D2X8WmZ8fii8Mkb
0bWqzwPr2S+Mw3vgegicfGMmRwglNSfpKLxY67cSiifQoD46497zfN7+LHwbrkjb
ycLrU0JhfN77lGcX44zTFuAljps5vUG1hambMhMyL/btnMEzh1g3Mm86EYd13n1C
nYhGDvDvbgbAQ6m+xqHa+O2hI38tUs/vn3zRsMjC4axQuCRM0PlZhh80mn60R9C4
J/LB9pLjy7o1ZCQonG9rsAimygrNH/5F5tqY2Uk8sgOCrJnYzhbrk7oK+FN9XTo3
BR5O6qsKw8d5EBNlGoVvcJ8S1NsmASEyDD7sO2gsWGenwytKm0S3TqpCeukauJD8
fMF5zCItvEF/Bnac4Cm5QppFNs0MLCRIaDgq8m9vmNZ3o2ocYcTneOTPErwuWuoX
jJZ027Myje+kgfhq3aOFEoqg5IQh6fS4/53r008IFyhxXDSCkmW4plVCzcz874PZ
WkvQgWtK3vT9QCa0oJE9w30pKAoHdOBqgNR0euP6eRS7ZHkI2ra2X5+i0XbIS90k
xTpDq9LeHHC8yqa0NoyccqJrNpt1qTPsfBF3fg1frPAIiazKMEpYye225SktiNV3
CDImZ6kgEbBD7eOgizsA/I7X5EZyJqIBUQM7POGD9gVLyRKXYx3AQBiiFsZsvZWx
X5KpcVMzUMTUfYnCIXEBMQgz5w9GER1DF2jd5JQJDrR3RdYhZPArCOk5DO25ofEi
7veTf30lWBi64oDBImPjnKFzTW68701qhKHrP/zUFrEF9TDzgIOp+f7mdnIHaLdD
P5rh5R2IAOLw1ppuaIRaJZ6SNtbUNqDKCcpAv9hf/xwMtMekna834aQCFKrUwgta
S5ksrtmmxiR1zZsdfZ5VGqqC76p+G9EYFmbO+V70wrW4CpnXd1KktFolU5hYfxJB
3Wj10Mp+AHS5KRS0hWoa98qxwSTGsenJgumPbyHYnAlRAkH/I7ahP5dK0HHUXGW6
8dZrZIHrHJYHwZjhvSfXHGApY/RDbBMQuwzRk1x8N9A2cJQDlFtUwZ/AuVZOnmdH
eOdoJOIc0yVEdpV5YwYnO6DD+GNkmhXbrlb4SDrcm7dEnXM4hEdX3gm4Et/HFJ2h
jn/IUKtMv6JcdpPdyjizjlpja/ns9XpEBuIYQ8iHxWj2UN0LwsUu4U9n42NEpp4Y
YclE+WezUKhN1l/jF/N25BmEnHtzpXpPj8NYTsgwNh3/fF32ZrCCm+hbtVi9VHze
0UiCSZOOQBvFYwOQcwrvp8yKj5GYYpYQTwNYuFISOEj2uorYL3dSnWSNerrUpBRk
yxLehu+jkE2iaCgYE0a1iWjG1wzPcaid7MrOi7ysTfXNt7+aLcKRBlFxgAlyGd0x
xrlQs81QtSl+U/wQiCrpz9Cgo4iUrrYbv0PQgxeQ1ev4mnI1oLvDq3dJhiLWLHxU
Z+o5YcnyncEgv1BCPOtoLwbRSZE+6l7kwhj3qv008GTOcm+57XdJyVYX4uJ/rv85
L5V+szgEdZ68QKzVT9xtDlkTlaFs8cxrvlqL1uJISOd1SvSkC2WVMcztamHAohAL
OqttHQJ2BDreDkNtalcfYNI1hIGpYpbfjGL1wbbOnkCaOgl0NjPLHmqo4CB9LIDr
NQmkGJx8x0bxBk0UtxrpiY24uW4Wx4jES1SR2sr/eL9p9PThJpgWQNrQrTcrRXXE
EmqZKf/dvg4OvWIZKrcRnrdIErgmRvWA50AW62DGyPwJym+DBe+Kq7EHs+E8PDKy
Drdg/wUK+Uq/sCe6RFAlHNSEZVLZ9CmJRfRnyDfqvakN4tokctA5OCRIz9nXjfkl
HduCKK4/dqRYJn6kiS68CWOmD0+S+Y66MPh0P7wkMnFPDvh0HiyMMPECoAuySxZ4
aBQza7sBlA0Mw1i0hR5gNERgHY9lEfj9YODsAHO1LnVqY+aD2+3f/Ad73Okp7N/b
zapDiDh9V8e00nEt4cBQizucf7votF0X3lk7sRj4Fz4tcJ9A0LarSEItkeBpnv6V
ObnYXK1vOpJaG9dEmvaGZfgNFziH/nOyVy0Ks51YOoTvnjx9gjjfKAs1TvAc3kH4
ib3K20OfJLbrOKkpS1jQebyGYr1TxrJ/BVfThZmvNgTV3fAqWQu32ZG9HLLOPDJD
YVXpjjRNtTwFrdO1CBmZUkl2PheDg9GtUo3NTCIxS3b+IG5BVlYrkpwXJsL03Qq2
+p6KcdZFOzzPDSz30jxo8N3OJYBdtEfWEb6BArpP4g2lmhFcQ3kmyLRrxYcd4R7U
dK469dVE0N4fEk3npzIOmO7PrGR6jUcM0OUlKrluN11GVufx10TXoe8d3i8+bjjL
ApMVYlKVLbq+PhDavUYMfTiJtzmcohKcvZdT/G9acg1BJAw0PbfTDiwUHi/N+K1+
sJ+rxZNdiuQNQQ3Aw7SbpNqYuYLtjIBttPYNxCG9atZbkIDqax4t/mM/VDGPDlQc
7IofkntisU+rTBYXuNT4NdKEAJlq026Jhyws+sQ6M1LOuwTZ/kaqTWs6SA+A401W
Q4qDVZJ/mW9oyjYDaAAxKor0qlrAgvZz0yR7q+xn01s/FIhyBcn5abNOYnNa27aR
DFQmUYdpmEyXtxlyurm1F4o9qiMgv74Fnp9adqqdb8OqZlSufdO0oqdLrUpIr/8F
jhVWifSEaSw1hXDi6msizRoML1guG7/1O3tOoph9iIH7AF58ZHkXnmrFsGgeOcgl
jnIqVc8nMsl3v0a2v9CzOMQD4NwsCrAwIoM4iM98qVeYWMfx6spB71/I6ZQNA2Ia
kEwlqD2fzf+Vw4DLKDqa0tR1Uyn/Fj7lpjSns8+7atswHzID3VNylE8jpbytUG5P
0Zqz/O2KijkXY/BkBFA1Q7s+aL0fY8UFoQZKhz5zf7mha9dGiWArqZELU/Nkb/Iw
76ac5esHgeUtqxafL7CNcNIV4tzyDONce8BKLrAWNKHW1AlrN9MOVRfh6lCqIByO
ASY6BtqpLtYlwNjr7ac7i7oV+GloqKAOlaTL5m3KWmAlbgtsccCVGNm2tUZsnZxH
wHWN1Z82Sr7qPXX5SlT4D8kMDXfqUjUOrWf+9b6TsUGGroUgv1w1sKkEGQ9K1hW4
7dBGyF6G9Bkm0vpkYrzoZ8VM/Ih4Scf9PCWY4jUIet8iWCZcsMmqGJnqM7QvBrP7
14ah32/Ei3N8s4hQhSB56dnR1sSZLnknooElfwctOC+bgBkZWe7seT/2YLAaLrm4
p9lkSGmuNRsFXczVqYH45AO4EFd7wuHNSYrClPV0911tXI+LCYrOUJvk/nX04rlC
G1dE4gZEZT6zvohnvlOvWcsbE88tfhYcvUQ9DRUOksh4D2WBiqidgyBIGz8ReaZw
TAMOfXGH03CfgkuSkt4HKN4NBxXpL7owunCVkkcDkR4ddzIE3UrnwflFfQMIqnEG
+bE6gV++wlj69JIF9gA8Ng3JbTlLz3M+PMgjjbgh93IGk/QcKXpB6+rKPO4169Ih
p4mLZ3XOSILgWh81q8MKGcGJVPO+By78S78A0dAoIn+7bS/07thRHWK3sHAqczYq
KrpdpdDPZbJqvH2sV7ChrXokVqf/2DV30rTIXKs9n098mDnHfgvST4mXA/504nSp
Xy+H9PDrOUYk0jHg5pCaQtRDkBJhYap4Mfc7FnBCtkZ5aZ4qU1G6F3WIEq+3uDlJ
V2McIHNlzoird0DZdDoVMYPgIxN+UQEhxiEt3AnirAraTA67nKQ7uell6xJonw3v
OVX6c/b31sazWm55DxN7XBOO1TsHtcwDHot0UmpA25l0iP+fXDoMEmTr+wTTHkxJ
iyPEPlFZr2bvKM+c4X6Fr836yhguJvgNYLrSys+6X16SCm/BkeCpwg7EDfg6j5rL
ItJqpfXfoHiFI8pBYGNrsj6TPJXQV6XscgOYzKmgoefpxQSDw/ePO97Vp7zyQ4E+
7GroqTCdsuxHRB35nqidyO0nELOX5hRGZOA1fVUYJAO/2lKnJZZYvx6c7z3aFrc7
rDJNx1y68KqsXCtLrmPOk5fYFdGz8rVG3JlCSMsz1dPWIDPpSoxZ1l4XfmapLCQa
F/kPKFjlD8v3/xZ8myESx4YczbEQBttIejc+A/rnwt6yCMcRf3htI78qmuWFNN58
c559BtnJelsD562Dza+DYX7hHr8Yb4EWvgnxmF6wMO5u/YCDL8fZSq/GQy4Z9AWi
CV3Mp/JUEGPk0HQ4oGnQTJ8cGVOcWr2QLrHQ+nDY9V/idRfa/xtGUniNLwzeEtWn
P7onTuVpvkWghE/aqqHUKyLfARTvQD/YYiJJih17SwItz6tLo3b4VAgR7udL6C1i
JqIKTt1eQGRz4nP5Z8w6rhjABUZcCmQ8S4LqEptihFmRBg7adaMA7iLEFiBj6PdB
gUccQi6LmCMBN23ds2zit4e7ojl1PgtPISL0sVdwgLZaWOmfr0cbipH7YdnBxx1U
x99GaJ7a9frAYY/rJwVKTMa06DPPrt3Tbv3pIrmUKYSUrhzF1xU3tyk4MVa86XC8
08zdUJDJU/mSlyYwmzuFT3FV6Iuefd3+VKVo+tIjvFAbG04hQQw2j3XNQ9nxy/R+
TNc0oueG7ySeSmAYz+71J6Vf8oBXsAINKWYWIyajRxxGT32CVJvWY9Ttn0J4fHiD
BSu4YUUiFimhEj+299cq2wuTvHbecUAzwqiXx6bc5lMHLzR/sIZtEMjrgG1f0dyv
4n3O2eg+K5TCTuKsueUXzaVXMYa6n5MpQvaBsGmKYFZu0HvOIUAnRNsiAOUqYZ2u
O4tyOo60mnC/lvamT15D7SmRMhnKP0j+ngpe41+ZyAi2sTHQw4uSbR9E1WAv32tS
+ZTgDHMfDAhJxiy9nru6AU232qkHzdmBGE+K4vEVKqFATnWCBgAPmwVtLl4VQxsg
DE2KpqL6q1NhycVR9l8LQxzLQpleH1ldPQNFQmtLsDIp4wHpifrJE8ilAS88irS6
nnAARjvzt8EcyFYhinr/QUfpNbQ9mM9VEDKQGQzpJAp5TTocWS0/nqs7N/mfImZO
TgSFIFk++X1q2g+al1J74jzBe8od4cbbQzyFRB4vpJjuqUlarVv73ZtEtDyoAJVZ
wMG5Yn56A6pIgLVFfUPoFbgU7ST8AoeWwg9JsaalWT2uxhxILKuYKUZFomUWdA/U
uiVUNvNfGbUn4E+7W7JvR10imc+hsCDnGj2A7kjtnM/6r0IhOEk93OzNvAjcDOUr
9oR3wxLYkZ0TNMwWdk8JkliAd7A8lhyJNtT0/WiVCeBhhDAXrIuvENBrrzE89Isg
QZYS+KsHC6cnW9erIbj/uKFJmJX56KIGmMTHoDPya2akMyhv/TcjgQuYTRLFFwMt
4Gwl8K3CY8lz7ulL1AcfMro6yMkKTtaV7QQdjzrJs8c9YTXdAfPXhoGB3VAX12g+
C1140Pzakal+f+0qewv6/5D1wD2CvouT8ejoW/faDwuq7rxJ7yAltOt3TCr4Kmni
TSj4Poycf56WjrfivkKURTTu+MlsISUKy4MO7izpd7A3BhIjqIrahqnFt8FaJI7A
0xMe/8CPTaf6N8dEyeyq3lpNWVNRs8A9AKSQeJqBuoFf6/6zeNzQo2YXuVj7zJet
ffSnBLIJaStUyyN6SxJptT62mdU80EsL28l4JQWpF2ZvSi2QEEGLCzq4aT/IK7qW
pJ226HUWVR5Ig+44kw5bMzUYBD9qHYB7owbGBRnyv1tHIwdKa6r8O/gU0tYBU1ti
DUZwPF6A3vr/SscIET9CERSvZEqpbDzzJfjq3MFcnJ8lfmGJ9bXf+L4KF8MhHM8E
vzIl/AMITe7Xu2WjesiXmzhGUdpi6hYcxA6DmatQ12iGZ/mP3nMXo8yFT1Yb/W82
kjElG/dTPbHbA1na3He+URo7p8ecG/8+7jmsvuX2ICD/5OWsn8YSD6D5KNfMIWF7
OAD2QJtcrD2Vr40mHNqFht/soPnx6t9VZkULtgtxz45oA1DmEDrBBMM/DfZhd/cv
ARlRgV7Twsw2MOesGFGHwrin0ZS2p/oFsKNWt9gE2cmhAjhWtqxAIimjf6z+da2r
5al+z5RnSjV/F93yYGvDqIzfHJlBO9GQDXYhqjM2l6y25+KDW1YzZwv2J3NSIoVt
V3rTTYYnv4t1xK78KjoKOWxSEGf334VpatKs6LqtJeKBrl4TNaAQMzLijKdq+euS
cGk7VzHWO7bQMw6+rYNKHShqUJytAteCJ9+NMfdFaKNQkAbCtan2iIxbQHsDypbT
UGwayzYkQPltNbb1qTAw3kNxh3FJtN+Golr8qqYk/tgMlC/LowanEbr6tyz3juVx
QjA4NZ70hl1IG0VXPCrXKgFo9j0LYk3H0Re7V9wVYIqJ3ncxsmJW7eqzI6EFCBc2
WOjOm6hh45nJzo9TZZfXBVbOnB++MLFs2RcOEyqYDt9CT4iY0PTsbsVXiKuM2HX6
DoLNa7/yJvY/14bbnFOrAKtiuAHc0ie6CQEumep0odLzhI+UL2Sd5lwr36ckzh2+
CIM1opmYzR+i1Ah+zjXugTuNz904u7hL3Rb6oJAGy3KcrbBEWYzMwQei2LOaRd6X
k61boVaxIMntmgUNycVf/6/NI+B9g3cgG8g8rK35YyBgvldyXFYyDWvoGdPXF0mj
3pJc96sgFGAjdb7rK+FO9++CoWEML1vTwS/CTSsZa7nG8aNas5GqklvANaEmT8Ga
FklJsX4dVR7fYKG0AkTXkS6W14HQ2LwsVLrCLlcNnzWM9+1LmFwZK8BOLR0Q6sLl
jHMyrTILtWIZn+Fy2BOgf+HHYAaMqRxfIiGGjhgYOW9PapDtsmoyeATWZ9wIeY+k
/Uo+zHJproN3fknL/iGib+XyuOPynyKIQV0Ef3YWYGLIVNUekh2LiZYsvgBZVKfH
0FND0sNf8H5zdnudibAzYTwcwgyaLrMGCG442X56iIjDThuKa6t1IPJ3RgwKTTbq
aS4YA/pbIMIwYIzxvMdEPnDLJQHhBUYfI6bvu8WjXJHm/LoMW+OzkQAYUnIHj2Qa
RlLYML7TkuAJUIVoQFO07Ow9IqCovu8QuApjmQDZWzp0MF4mFeCfu4VxHDm7ZKvq
lMUpAMykDsUtqaykBIXC6Am9f9cmUPIiGIQFXKgVI+nEaTocDobIuXntX5y8Vfvt
FAjFeAGmNGeOoY/OX3dTuhHb7sOyFMFd3Z3OrfNvpn9JitU4VXo+n55/2gQGWU5v
Z4xN2UKZ01YsRswrUWNGuUd3CANKNAcxVpFL+0FEQu83oJ52WojOscEmDNHenpHl
/KQPlAxSPPLyGTcuAsBYVJgngbviHV3my06l/wD0mr2ibiy3YEXsrvjOWLBZAe87
A9DuYldIjFWoRwyR0FBMiW6lFSb90k/39ij1LzbRlzq1j9QJMKQjr+jQ6mjiCw3r
P7br6g1HgADjrk9I4EMndhmJ1JQnjM0qD/bEwrdq9D94ttVU5hr6VWjs+cRMtrtN
wsyngegiIKIwuEUbMfZvkwKICh40V30LufOjHXZsqIg45B2GWmqSBoI5TsXzucad
CPzIdnV5hBGQElZ4C7D1pgK4WHM3HGKCxg31w1HGoAh7PLSG8MX7/tyYQteM6Umb
TQW8Q/2b36SwUU4B9z+J2LKgFxQIINCnax4nUbBlwshOfGySplsLQjLBEgnCwn2a
pci35AFawscGV1X59MzC3EKwwmiXBJet1hvRkU3aZlt3aVHYVYNGJyPh+7bw3I6/
WT9NBnQLo/tQaEPOX+x6Fkm8AHDp31U3UUR6AvyOpU+XRF10bKG+wyC3Dc1g34u5
EmzNxfDRk9oSVOesplgidvfso/h1bwEmbdftvZiYAuL/7FYUYu53S53kAHnuwnB/
y2K7y00cq1YMkMvPo8QjvBn1xpaahoLZJPWSpNx7xT0sRkD4+YHwoSyBsiEOZMTb
ef3KFSbOqdNipm3CXdVyzCie9GPEGgtFLq+hMPLC65/uS1VPjXZVPqseMdTMg07c
gtEovWbt6icXKcTq0iOPwmJFhiAfXh6DND4oGm/kq31Ng+yacY4OmHhPLRpLBhL+
oYfe10kIt3JXpRzmelrIvmjjLA2saXwVofnRjfucEkxFz989YkxXOE0UC9RnvS3E
TzzQyWXxv3s+lROSuZO7AWsRCz52SXyugDIHV0KhHKIzT02sO1n2gGDVykEuHxD0
hftSGZqeSvCby4yjsqDhvOpVZDwS9/PWF808cK+G/CdyQnFmKcLIt7H0krexz3gr
kENxRM8vR7KmK8aXYXVweRhOWnDeZvXSXgUU1vdd7QwJhwwgSkBO9pP1mRkZOVyk
CfhAJxz7+aObE0IlRs6M4aGvsZfIzOpAr+bPvU0VFgubxWWGqM/pIILEf92+NvtV
bRSiSrKeJAWdkuHJtdUBGeLMC1KImnZoBr57dHIxBl4BvspRZu0JolFazvXwhxZo
IGHXyqbIPb7s+QjoLLHdNHOyKAIbAb8vfiXu5lUltWHwxUuHsi0Id31gsRuCp0i9
nFo/6xceV98w7KLEueGWFk8tEXhEOBU012d0WW8dUgCk1GTW72b2BIFgvAlrQGRb
NWloagoGokn0Uc1vkt08Ha3w2NFFfLCA3oGAVBu1c+mvQ0V+euDTPOIiaVjmziyZ
W1mVGcFnQQYRCAync/YLn0ftbghR1ZQtMRyDhboWymn65/mY+TnXhJDMCrOb4xwr
tCMeMJ19JukE33fnomXAPI0k3Ne5PBnJpvnRFTBOVQKIQoFSqGK45ZbQWMXHZ5aD
tzd/ybvyKF83yHI0/XZfd3f1jeoAsJ9R/vMAFFQA/HNp5vtWE5dJT2QkDmgibwje
RvAiqGAixgHkF0eNjpcaPT2hguF/ufZQuPwhM4fUjZoxJnrUUWseZA58W7uxuTgx
JyD2XxN/ZD2dE4oqHA4lU7GoWa89b4D+Bt+T5lZeZbIGgbLo6m03zDVgXT8UxfuZ
j8/V8DizHn8cJyW2P7WZHwjL4Y5NVjjXS5YAmBZYg2eG5mg7sHUo3Zsf1wvPoJVw
f58qmOd7Gf0V1h/XPV7tmZPYXRfA8f9B6gPPw56jp7bcJBI1UQ0k9mwaUhV7cFIN
UNSpxBG+GFFFkv4gJ6Bu2YorVuPICyOiKaTKcKmzuoS1x+IttF1en75/K0mV5kmg
VwzBn/7KwOJWJVdJ0cs/d591b0Z29gR5lInj+uMKshTZcZP1VpnRJzGEU8wXvCvX
uji51hMI7Dhj/M3iufeoqS7RZtC4DtRteUzSspqhYJFpr+ItVu+rLeguAAMYyGp4
cahoCgsBiAEEU2XzKm5wH+oDxKPZb9d9gp6cHqzutLl3eCkqMM7Jgb2PSQuOjw/o
1Y2qcmy7ZonC+A74kZao+6lwXeihTNSfoDGp4EnJeSk3VL6cYEGDBRHNkr40NQ+p
9V43rGny+cLxMrURgSTgVUbQP3Dj+dgClUCbXRDqkB5KvL7umEELOgv/53B2FkUx
GFY6m+Wb78y7BepfCtn+sGpfjko6i9WLG2xV7WGSPIs1C+bSPZlUt9phI7OjvdDa
jz5vswyXMy4iiZT+JAmS1nGiVtOc7+i4dqRnvvYz3GPY4LqwxKpkCNrFwpo9GcmK
J2TrBAOUvCMBulsaILnLuRx0THZAp4rGKo7eoYyPdGGeIsQR6Dgh5EnPth5BIB6g
Ie+A/fh6OteW4PNLJMuPRdFd9zuN6Y7ZXcfqrmYeZN1DeVEzgO/M5j8TrWPGkrII
S2S0820xiWMA30BYso/N69qVC2j0RfXcRaK+/McSNOF56AlXVjxW8wF8seToBWTW
SxEXBLEiXZEQtopwrxhXOyyKR9t3YQHJxRsGDjW3VylpLRmdSvK4GZeEa51Y0LU+
OVEyzDRkmfd0LACAFTWUfC42MMsNGnibomWekKIhlcIDOzOf1oas59RFTD29QcWy
86eSnYHMCUmp28guW7WRZeioG0MBXNmrgnMN+x+nAtUd9LKelc7AqXhFLqFrwim4
1aaFlOyzaBcWKCp1uJbjmsZNDqSssKLiyDJg2Mgpg31rtoRaB1xzQ+R0gNdTjyQh
DXPHzDpJ7mnM3ZHuMkxkxx2RWfqOu04OOhwbyjkRd+tbpP9h3NIZWmcXD5dPo56K
2ZJ6vSLAIx8z53+WNO6BY3x9r/mDEKBXhNx6JPCnLxHaCZQB8z/DvxWhvdW9HSJv
T8QxkCgHGfN+BVOYk1A14qAc8FZFxLlVa2/Ah4lXumuO3oy3W/XhOhdv4nC/oPAS
pbRyWmKl74XmLpVlhNnGTRCwzlwxPYx8/AXt0UJh3YpHbPk8TS7f0TAeotK7VQBj
4fbGCsiHmRj4LMQ8t5y+JjumeE/y6u9EeMup0qYK8D46MGa8zkshINaDPYQ/X3Uw
LW44GiH1OslPHnlTBmEpnEcKd5tpPglYbBpB/Iu3O8v2+cPdK89PpoBfg3AXyBfK
1GhUm8rI0tvvQ11TtHFw7LiKeJm/gXTA0oUIYxtXdbtm+m8HnMcZklrfXM2VmJ61
16OsDrT/496wKdWzCHZRw2SJneUpCIfcbeCtYOFILTZp9L6OUoDi30QwOIWo7kFa
YTGdvMCmqtzZRVxEvVs/M5lYPYYAuSKv8FhVPp5iEQX7KJwRFc4MFGwrjCKXDlPj
GwOBbWQV3VWwDF0Pin9X7FOVPkYZP00OEwc05+XWol4ulvcG494/cQeJatJIoCZz
AGzYG49A7JPhWgBaKfij7WprUaHr9vGCZooHOpiqXWZiMZpWTP/L/m8B1HMxk9lZ
L7ugdV80ZyzUBLXdeUeyGRT1xegP2htyn25doBBjO6B6Gfo9Em5kEx5gSa+YOHHN
Q5GJTNS8cfamn6my+sT8J79P92VZH2o1oAt1H76sYdn1A1Lw+m/oVjp+sPGiHUbX
nLfxGiOhN3wW4A43iRb3ICH1Evfyxbi6q5LEMHXLUBijl4BoJS3IOYIMf/wn5WGk
bIiQAZ1j7LYJamWHhsrC6jBe6Lrdr/lIYMKTxdvn8c4mZnyrVg2KzZ4YHOSKqUGn
RUIbmZVZSSMfE8kRe+LZoEgG+jY7MeQxVKjvdlbETdJLFkeGXV+dkV4f+u10UIcc
TSwvYo+GOnuGH6VUqZXlqoA2ee0hrPG5qQ+9YwHye5ETR6glWZzeajhCWc6KPKkj
j800iuxPIacNbo4CGguOnj28OaNgfXMFQvFSiXnLxpTsfPHEcf9NOXBdZWw3ovAI
IrI2lP89MekfovlZcnRBdiSndp5W2fT35Cq+6g66NJUEFUpcUKgUFNoymvysdfkz
gOx/5n56txvu6myaKhzbS5I9qsfQ7iWcXTDCqKCmRraLG5YZkqCa3s9O8hvRDtL4
tk/GwQB8G08B38ZLpL4EZCp66/25IHOJS7VbicD3RNEhBuC01OpEqrDQefxkuAlA
Nd3QV851NndmqqEFXCgyl3cHeSZd1n7dH2b+2QP5xz94gtlTUjrhmoQTjFY2NlYd
FTYieQFZIVnRJoP9HqfsvEyZMgZ+DQ6eQUYWlGQL6Bdx7xkr11cA9qd/xFG5j391
H8O3arwVzl0jXjlgz3TDPNAH3M9WdyApDQaHaq2Fvfy5qj/cJ9B4r0oVvL1K/ayX
G1ZxGBo+gz8+YhNlF3hxctWzBOv34+rNZUlQqOFoNyfkZIYQijvqsd/ImHEQTYNv
VK0hNRDV6yu8YZLWHIrtQHh+shQq9JFq84lzTCUvDw4bRjDCeoQm8vut1Hic9RoD
MlD/GYkHQpQT6mH3hoBOeWV/1mVqbQRCOKsY51Hjv5ZFAs+coSaWbA3P5hsjpQBg
fjrPuoywJPJoTabtxVNq4LToCm8/P0wWEO3pwsJXS+bfKB5fvuGE0lEEZ1zqNqFd
Oc1apaKaVOzzlIkl7CkU4Zq7WRcwoyWP+u9fIGOUIPUhnQDOnYerQsFQqXNUOSC1
9tRLBh8QETChiUdCEdCOwMrIKx0K/SDab/WzO1KH0CRkX0uFpH9HlJSVhKHalFFm
3yMn07a5VBYlQrIzIudyiqyb0tdApZG2drTKy5NwhCvOxcQ2k5KYMY1ytckoLdZN
pJ9X4RSbWFQUMol0pgTI02SXexEjwwf3lvTdT3MWsq9wybIS8vmxBozqMxJpjwZy
FEdeLOeUoAdK3DU9yDCcC0LqPc5inea293d1k5ptjWdY1Fdecwd+GQJGk/Wb9t19
3iMWMDjaWElHqiGE47FRgwM+xqrf2/FYJm3JsNArwTFo1zs8ZifZKzsxQGntRdEj
ft+K5sSdYMERaXJAuHNprVoELZVjIErEr3z6bH9uGvPh9fzKFZ6gNFRuwLMnfB23
neBzrhmFaTVUOJWEnO19pV4n13OXpqZeQq/+Nxk7bQhLaynSAjRfl8nQrLEZC3Qp
+2K/PakQMk2WdTKFnjFJ35OnAYjgI1cFkuabdNd5cjASK++cccA5xcCa91st3FLZ
Q/B0oRVkuA8RuzPA1ha8dN2Z4txV8/QTOE7sOhTcNd7xSBuVuvT8jtjwDImtyjeA
lHfbCgwOeR91VkjtPSzGLq8bZfgqGeW2qqzduYFv52onHvTMiAMUIUa8xrFw0n/n
aWDWWHqVqDOSk/62zGdsOMUw9XOYzNsUGMSQ1pvi81bo4vsN0VteKlx2eeuXGZwH
vk2r5Fq19JZ5RQdt/okVqzvloLuasEIaaZbsLgnZXnGS7+oAXS5PInHUsuOAbzUp
XyppKlxzl9C+8uCth4R4qF4UViihcIGccPwtCKKjPdlRzwVsPqU/wDOUm5jyMbwa
fKEy3a1HbNuJKLxqM2oJ1si5EZvUf7qXPY2YuzxHJnY2lN4JYJiogLwfR6ZtlRF7
Dqd6ho9fIqbK9LC7hBCjHSjF5W1pdZJt5FWxTC+8xh+oa+mtJIlrB36aY+CG3Jd1
dzsBXbc8Cz/8Z0y2l6GcjfFFgq1bDVlbseL8lFz6vPGnSo0cm+A79hTGOvJTnJsZ
782BR/uYvOgXW2n6UxChB3RQtKJ1eGKy5zW6lKuAybbS8USRgeO7MLd+H3QyaEsv
xgtpsw+4LqmAuprYMKGugL9SEH9Wrg8GviWVvpxL+zP2ZMj0KaQoC5Oc64GsvEp2
GL7gFFJ98BIsnUrg0B3QJYWF1VCcq/XO04UHry7Pfe4BJWuI0ADg74yPHkF/R4Nw
JoAYzkNPzpJAfDQ/MtzkMdONOlLv0pskuOSr+CqVfe4sGI0+iDyQXZnvMS3civg3
YObllE8MJ7M7HNoNbGvULYPC+2j3pusgSie7LGks3RAAnIhg6hUlYzzbWrXUBnX3
MND9t26m1k/Q6irC0DgD9hH9/uabjmxgGAKOfaojf+GEJQ55HiKoOX+3dStjrSl2
nLtH9Lvrel6LNq8WD+PY6mNOEKHJdnOMH2wlbUQuWsJuyQnEj5z+VG07FXAB5gRx
3bBwCuEgo8srhbYBPcTa8WThAkX1DqywFDlVcIplaxeH8mkbXpRcfDth+iKFgjb1
6U/ntaAKJ+0m2x7fx6sdRGl0eJIUUwBemgsHjSydY5CXPxz/+toUnbwK2uUaaRSO
RwjophQkbllDxzWESznZZuyjr0ZSH2eYGrgOJP1tLKEnnMqS5ogIROrIxsUkGa1X
pdYABeuG27RoSVoM/iVSeMpgJc4p1gV9YwxaU1g7/e+tZ6ywYQPVugMJ6c1D/RAb
ODudR/XbMobRsD6+0/XUuKoTSpatuPQOEwCGJ6o2x4Q0oTBC1X7VDPHn0VlGVUxY
qjFJb8lCEBgm0B3eo1VX5+XlUQRePwkC70lOU4O6mGX4E8LoV5u25latYwlL/9NY
F0WyJ0PIWL2e2IaJlTBaOnKizDcgltM2MbLT5U4GPGW9GVQ3+MCKTHscgSXQK7mJ
RQpnve2CXwQCtl4kZBVwtIe+6xJb2KErZwBP4NFjDr/MPYOsG9VnNjLpoSox8oGA
I48NmpezdEyJ8hhQGvatXwyFxEpoIIYMMJmYUcPh5R1bbJnFajJMtrb81sBnQl8W
isrtfPKve9dTGxRaamvk7zy1b+7xgXelLbuZUqclCjDS32o+wH1B5DlTK19L8K9D
KeV9SABIldhR6vZQos5Ohmflat1VgUqCKPi/3XvXa1hQFSEYN8bY9fbjgf7a4j53
uHlxpSZg1yxY0l3JWRcXm4KaP8nVfFJTqU1vCwbkvuNWA1bLyec3DPVROFxcS4Kl
gPRuL9YT4AB84SmYjsD4q1Ngw2+H/79sTErFfeLL/Ou4sLjtlOjErkE6b2lonTC3
7L9jyoQ+ksToZylWmdfxfjyMcxQgnDUQiX2xbBKbLY9dKKiwnMgqH37CQdlDI9xE
sDHrAugcqX/RHhLagbtonGVGb6/QNV1pXfGGJRf+kTPPHL3pXQdHXRAww81ykWg3
DAf2KtIkT7nRTk/wYRxGe/SMCtxAxJA3HvsbZOBftOAg5/6vE7R+Bjg/qw1TNMNm
EsnRPjamf4XCmyPWB9Oq7UAf03nDW70WaWUKSNvJvRAlADSMkRki6VjBp6yx5iZY
Y0lCT2NRPLaDupw7E8qG2e8o8UkEMhG/cSxemKMUJEfZgQ2vmRpUdE2bTrtidNUw
eCkmBJxPtt9cNk4aMFu7BIrxEmz6XzKNQ7DRa2+kWMA=
`pragma protect end_protected
