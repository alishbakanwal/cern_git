// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:40 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
eyzh0UaOEvezEpB25BYKAqtu/Nvtkc6X1ASKkJee/Lsk3A2PdEalGoX9fa9eJoXl
Zx1xq+fuXKvqSwl6lb2PyHvB6VBDiIQwCFFLcRtxeGgCcfhjHExW+RDJ00kHQrms
Z3QwDGd9nuir3SVD1Ct+98ZvsBXAZeTV4xloeqS1LfI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30640)
ykEahzQa7gvNMZt/H7tQFtnBpzu2kJcnfXwHHjX+GH/1vFmpoZVX6vIUiohU8QHO
crBoyXr02s9/qSISKcuUigvZUdS73+JNpvBbV7kZgPLK/s78DZvulOkfdxWIPtnU
2SdMHlErvfAlkiegCeEwZO2OOPb9yQiA/0IciHj0pDmm6i6MfdS5xucOgC5byzzK
uUvdRN0kPkK9KLeCCqy19BLa6MxPCKQ0q/2Ivb7v99xfP9rDx3oMljfPhGUMnjag
2hFmOozA8mp7RScjvib7mXc1In3QEArxNvjTNbW1yNoO1Gbr8dg+WOv+/xIIZs9o
ljQt/KCXqih8uz8zbTVDE+3yl+W0fiVBXtCre+enfIa4n5X4cs3Q88RGKqQy8A3w
aHuC8Wc/7l/trI++lwGIk3jzBT0lrt6ovHXnPaZru5W6+I8kWeUXbcWLt1fEVJNd
WMy4fQrQ+6ZozjEdgsZaFapGjuXHrjJfoT3i6HrAOr7ArInTak9a3coXB8Jni/F0
bMAo0TI9XAeqC8RtHD1f2j1pOsU7phisgrYml9MjYaRt2EtbGd/mN3BOi3nwOH9T
hCcTk2ARQXLXo7X9PEDvz4KtIx+t71p2LQqHVM6nOUfkVc8KcdlXjQ2AhADEdpCL
f0D9IpPJ0//1izpSrIkCBk1L12mbZ6taltczXN369lUcIry5HVdBezvIJHXhvfLR
3LWZxUyOs9e5jBj6n34JZa20vdKD5/dGoeEZaBk2i72Xi1hPCJcHVD6yoFXCNbWE
hYA6Tf4s/rBdSKl8BCebnxrxI4kbl039NZqIQX5vEU3ELMXI6Zo/NvA9lwfMbxcw
LNIVnE5k9j4LDvt86D51T6glA4FVt8phDKjZwp2mKKbHCrYjRBNbxPfZD42t9BFX
S0zh+flPCYI7otbhUtLC2eb8lVGlqbaUvBSjpHUIiV91GZDXD5SXP7DtyPRnOB4k
Fb7SbNuEtLBx+imadowh16wD2WLNfURpn+vRFbVZEy2Gvpt8OHI27kM0e2bBXqbO
ewkUgs3Ni8rHKJsMgSNOhXpxIGXVfW+s0Iu2zXdN/NsU8uimxQdo3uGy+t5fRX58
9SjkENCahSfC66R7ukXNOHFybhb09wCec0paY87fSLMON7F/ZN5i75Wy+O+yYh6G
xzCXrEBq5fbVuoZkf6rbNBei7qXJDaz9ptwvd5gMeJhiYcOEGTMxBgi7VEsBfbpN
t0jPxXuEhjqtv5WxG8Ljq7Z084wdYfxr9JuBdBt3YqDCClR285iuULtQ1SVwJumN
zDiL0zht7DUnVvtBtRDqqCZXgOy7ZKdXIJp+T5PA/OltKo93bql/CQbPrjvi49Lw
ZpU3RwjGE3glBn1nwK6RyUT0BNLZw7Iiw6Z9ZAsJq/R7kHb86HA/1MuE6o81+vsr
gZruy0Gf9LQS40TYPjJ8KmCtLsmug/NQD/7WZQfC8WTQL2gkMgBrjJki5bCyQo60
fN0tl3EXjz8zPu28P0EQ3v/RQnr0cNdsDc3ZsDvGAO+i2mSyq+1dGYklm576EgeN
99Gixy41QyEpiLEx03sELM8qCLSt0MImIFrABDEWFah9t/udYq5WmLhXXw+bcBrA
Ei3Cr2HmEAXUg3ol9uKy5p3c8b6CNiVfKcSYmxHHlWJ7sGXvZ/xhnteWRTwzUX2O
n22n+cI4hxXkP2/ixgcf+iDrFC/n50BQ2wit0at6sV2DcieWw/9LLoip14cS0Tf2
kDmJwVcu3FUrnwQR6qN42nZVvDvJostQKVZ8blFlNX2S+jLAH3w4WjuSbCeCfYHM
HRrxuySu41MmGNJui1JuvMgNxNB+umqPP3Xhz2M5flmdokECj20V1pfY01X+mFEc
l+hY+iaO7i8hVrli9h/LheE1oTTrdY+f3reyjD7KG5VEXMvla9i2vbbgmmeuLXZf
g1KcyoaBSF1uA303pqNRqvCBFWjQSxV1EUj3sIPdFAvXKCqo7VkYSqCk6jq7/9aX
fvwSCoLM7lI06fVzLo5TfAqQZqHkE6BFlb9ucES/A95msdJGJRhfTjdEL8oMWS2V
f9bQR82TkxqTtVsaylvPa05WAqe9/tB5C9719RGIEXriwKvfxaGdxrVC/afu9RsB
XWLXbFuQ3dZW/x4YnzriG/MCcugS7dZ6olUZY/zraerp+fHj6k7E7Ly51s3e0dnV
zbGFqXkW0gNadErhqLkgfuwIAUBIPIpIDwnQnhZ4ZWCN9ogNvUfuuvhs1RKKK6SU
/KIVs9qQ+b9pCaaLCGdcrGa+tIgLpNED9iGsLzMXSrt6yfDA5BgJWRkgm06pc+4/
5mFjctB2jVlwxk4xZvhbahAAm7xxIj37lXKrwFskRuyvUCkVGDrh28yn2gkdbMaF
QRdUIdBq/oq0IYoJWv6FZvRlh3XVH6zQNgo/LznUahVSKVu/ZJwVFDvtzZxWQPmk
YnKrQEkQJBR3I0AGEz024mDCSxsqtcAulYmAKh2KApQYXKXyNko4Nfw1PCqjNq4+
Z6bL/omz0dy+uRQGl6i/WggZV5WH5ErxyZ3qzogs3nf4cr84C9Arp2Z2ns6mebvk
ycNxwvP1TlOzj3O7VMTdBN6xx4Q+IKXqAFB0CoKj81p2JxCx7SnmN4z3t/dPFWqY
LFUW6om45hALaufXTLhEAwFYUrguIV+D1UpcHF5qN/7zYg+4PycofV01tReYieK2
h3Sb8pyAdaWUYXGjAPJlQ3yaxrfZHP3Ax40ktNEDNTKXv24OyMixi8JuwL+37oCP
QKvlHKVrjyvsaAGP2UGqPDSyfeV6jwmdetqurwatlVJ3YONUP6ZU1rT2qVeOfLfa
3QRdjBrmojaNJxoUlCtI3VI5jkGMQJq6vwks1mxxcF37cFyMxubP2d4IiDO400f/
a48vDmAGZ1XqyZkWXs9qfWfzWjDPi6BWE33OPpF0xvC/he97XFSqd0QAGMLggY2C
lCBos6QUkbnAZA3Gfk9peaM/C9hO3Upgi6JDgv7GPIIqZLxrZybLlcDNfHGcoAQt
DLJUzR2sEOlqhFYNv5g+dKWF5EOMrg6ZCyHxXSEouChedCKfQwlGusVKGEhNF5ai
0GCPlfOh7i0jVClEL4Bafmb8GzquJ84VWO8bXHTwfSi3UFWy0ld/ymHfyM7JBazU
IRAbO5lyjSU1w9cSfhveXCpTgVgsTQGbJvg3uImIUF3zUY6qo5Ff7m9K4IyqVXHw
yTCW4zx6C7Ate2phMvyaC6aORRRCR4Y4DT6KE/5WC/5gY9UQ9/3qw1Wg9afKUOUs
ZHyi9SX+/f+bhYD2XuUoOyixpTJo9rAaNFIBeXfYdCBZ9XiHHf2huzKXWxH+tlWy
XbHlbE2AVlWsQjq3WpJTV7z7MPomSBn/BoPVPVGEhf9cLBP6Ta8qNBKrMeeaOUXd
EsEwaa4Obl2lXuWctIwCAPg6P5psMewh9QjvhyBcGzHSD5LL/EiwxnHJMSUPoeUX
d/8IbEzQJQxxz8qNKgpFu7pAqsSBkaOrHADld6rh0twY/muQhTAOH7N7AUBTeAEO
etS1YwHSSvJe0AHrya4hCrLZPMBsNrFaUO72d+qtKjS9Z8RfBKruJzLcpUaJhtlR
gYSWZHdDBCkYFfWdpN2IqeBeoAV3jO/qsb0Erxwv6cZ5YZF5KAwHyb7HlefmmeVv
4YLs4+/lLP7Uh6MK8cT2aKuPIv6lzg1/jcjDV6i5PETSYoGZNr4RTm6TJ6pPfkb/
ZKa8wbu+mMFcUkzuLH4/CpMl7+ng4SkMHgaUu2OEWULPYzFc3nVeR1BLwqp4Vl0e
s7GKo8oRSWtyPWKQrSrffyu752lf/nY638pBJ1sp0BXgGdHtF5+aMt2rXicIvNKp
UXLbBgOxL0QXfw0xLjzsv2xtP71EmHIJ23lyyI9ckYxExzyuivS9AV+Ik2TfV69d
Ycave0kzZcAJiBMp2zPv8Lys8SO2Mw1s1wetiHBkeaAErafiu4yX7kzDxtAdj6QF
OxsgcMVje1DmLBtYTUelmAU2zPapqv8ahH/3IrKJZ8Xd3ENW7hjN0zREcKrio2JE
2sPgSh1F4kqSEG2sFBPFgmC/ey8vEjy2vg5X4jFOfAWAK7nw7WWWUlFdTwXnv9Qt
yl5/N0Q0WYbr2GHxV8EtT/XiHo4hjfXBge24+HMf3tgoYGt80w2K2KYS5wWOS+xK
28lVnPyNnIuzeiZ01kVdxdHiKKSzRtj6dyxWP5iX1L6oWZLsA18te4hzd35+27Mw
W+j73SyP6hpCgq/BM6EnA8boMDQU5vz9OI8EoY/66GPHAn4yMZK4jJ+ZiWIh2yWp
Em/G7ZJcfXV2uPEKrNGEeMo+jHdBzB8iTNmmQjm62nuRcquwY/pGlQ80MtTnCUAE
+wcs+3fX1q/p6H0SjWOs4UYZs/WtzcbVLiEBwbnIhOdmp/fnxTJlqiBkqh9J0HXh
Ad93SZRofTjmTbkIcVxjMOqwNvOl7urJvpBezhlTT2P5cbvZFIsarH6RFPy425I4
iZePm56QeO59M0BbLKlEvvVXvW4iLxraUSB/LLlRkJJvw+6zGZcPadYw/NnvIesc
62ESJf2zg1Eu5ETf0GhYewuzynfyu9Z0+OiB7+2ZLXUD8iVbxvY2KpirNtIt7OfO
0P99SIThshY+bPvfChVwvOI/X+R58qgyYiraYKax076D2AZC13vChPip/AGmLP8D
U9jV9egwmjyHOoLAQvhSdxUTnr1Mo7Zk9M3iekJr8JcP+OfFQyPqbC91Vmo8Opcq
zajQwpLdFrZRJkEH3GBWPy/1oHGcJZdQtvbxzTelIXyCNnlv5r1GwDYZ5iKSM63+
yO8rJgqEa8tZahIVbhIW51I1SVhd8WHR543JX7h2kvaoxHhHS7UozbiCETuU/cIj
lE9R0b3Ct1fQEs7vZYfhre8K0oNOSCQEcCMQP5zhZU0Imcpq0DpbXlV/1/aevdGU
BoX67JObyxrs42Ex1gQe065VjS74XLVgVDWGG5HlCMSYMu1E/rM85hzP4DLdTuAU
/ZGuTUIqJMGAsZsgIr0l0hr3cluo5U+gRIhqfYVtr3PP7C5JkCe69achB27HsAS/
vBjxLnkFYImPWoE3NWue/Kx8zTT1RSccwZQeXWUs30TgjJ1w9Esx31Hn+z3vz+RV
vDhDFrk7TODgDwLzX5Aia5IVjMFev3Cp94K96gtXnhhJdvnV4P47gRoapNSYDsbo
06/Xzae1Cj33gAlDaM1iBRJbQ/69c4tIlq/eFkGs230TyWzG+6phDiYfcugsowqu
TzMDIA7W7cen+uUFM5myrkcFW1kINZecKc/vBvugRO0W/EEyZfQFafbwR+tP3hvj
/vjojqHo8cN1+M8QVZd7H7Ji5oknZiuvNO5pVHP2MmzIfV3+smN8xflrbZyGrAI6
EV8MDKrPC/XpGIalPD9AygAMaoJhteMkiaqHY9fRpCUbt3e+KTAIna1FBhvXHpZ3
hAxARJG/4kiQ8H+XUYrzve7FvYf2mo3eMOhcQkQWPDrXJYTjFDddIWtcegvtsA5k
MqAKEwzBA+sfdp0EqL7YcxpQMXrOf1qT3Pgk0LMpaKNqVCmKz1kR8g50KnaGgyfg
+zCsiTxsQX4IqL9aPyFrZiPTbEr1MszRd3eC4JLHUFx/D7FcEjo6jL8+Dd+206VO
jyqlX/fsB/fjumCCA1fgoFMljmOyv+nhoRMLz5ikU1Ac/QnrVfl1ImaaDTYmz1+O
0CIp16YoOFw8X2bOFRk6pJ/q/PGkFKNiYwkhFgvA5I4kweQ2/QVQtaqUosDxvT94
0v6NBhHPeCvMQ4D+3Bixy4EvueX4NeE4oshVzc2+QWxGxfyktemmlfRSeTSaIrIa
XSEqxzcrCN6ZLAWusDfrFbgivf9uFPK1mGyI4WoZ1wQ2yWgday9mte3naLigoxQy
oF+0GRWn/Nk71uzzJCBex6rxXRJ4qs/FNMldEFHYPC2Oz7NiOKSY3fy/i3fxaELG
Z1ocRh7lWmJSt2be+roqBSY7OhhEcspNPhLrAqZrk415Fu0C0oqO37eqMTrWAIhq
kXYTRxWWun196hyRmvTRE21gSV1nLfRejyGh2mpOIzbdqBQ01Ue9TxDFM7pG+vPd
gmel9+zjKoQkvASCXSc9yh9pNbiUTjgnPo/26xdLDtDW00Ps8alhC6oarrojoCcc
alF+5bjMrG2BY1iO53Mh/G2xWnwXsKpHcycZXLrVDsBIoVU59T7mf/9gCZkXa3OL
MFaW3utrf57mtzK40TEmZnrwjJ3CMVvWjjzoNfKD6M6CaB803t2TEYuC2a11G1ce
6fQfDHhpDW0DsE8l/Ml4kF2EQhLDodkiP/iiTp6ctCgw3Hsj5N+ChUfYyseuMEAu
5ijrE4HG9e81xduZfDqjg9C+exlvRtiqV6Q9WWoYxUsRLRucYWoGHKsJcYE8LC5H
oiurorkMxJtVuM88+5ZdbTFXCFfSYv1j9Nl2OWgaydlxetOWbQEI9Au1nODvqrbu
pXjXHQbMFVtLutwLiHJR8cachldnZEmI6a5ol//RFWi8N9CDGLrS80Df/ikLE/+p
RMRJR/Xdvzkk5PNMfZpRpIyE2NgAHvNCIQBp2NgkWdhtIl/zgwAvKHuowLRDEEVv
Pq4zB45V7qTAqXDP759+PKmAiIZ1XOghXheS2tlFYVwux7MKfFlJbRoeSnfLQ8P8
eBlsEiesNVTVm0lOVBrqBWL5WxQwWd5w1HLiqiBi2KHxIRlJf5/tioMSoC4wPcva
Ed5UhRre9rzEG2xqLh2U3ROd6oXr86kbTqHRwXVS/E/PQUPaHWX/lEUwHuOYpdn6
4WK/w+62jCx8SeG73xM+WFPKZLPJpZLtyN+M5ZcRZti+aSd61kXl8M1M69A3LTll
QaFS11VK4+qurynpxN+goiqdnujMBCFf+Gfu4LFyAeCSxYxdQaTgBh76abvxjK6y
LT2G9YylZK4I/9ZjwCJuCKVYbYwsc27GAjhFG6/rht2UDTF21Qju4g1Rkx3YyP1s
HiRb81i6FzK9+je7gwotdsRpn71ZAFISF7b1VHGwXdS0EBErqAxkunL8pDybBfJY
MKg7pth1esYrTOyrkxx+eorLVnqxAys4KjK0/Fs2ykm999eJNjsx1FqIdhdebBkB
WgmORhBrBnvEsi+VgCi1Cmdk4QNXoVqt0kaz0xYn0XuHzY7maUG5bEpaQSSYLldt
hngRaASkmL6lAK56PvFJnK6mLe0V38x507YcnktYQTt1zyc/+s3djS5+QpbbGTKI
eveCyfDnemMDyfcasn9egMREh0ge1cLoQ+X3JH3Q0bi4qXLqR4jD+LbmO3HMDiRo
2q0PIoGTOOEyvw4k/Rka9sG0V0HI4kDr5yQ3fLuIKCHpgX0NN+K8lsZINoaQS99j
aZmQ+TrIqIGEvUrkMLgPGxluITOzyfpejMURGE6EZxowR2srQmUAiGFpXexbmqlE
LV6+Pm9dG2Vp+amqmxSP/Akw3ITFrt79Gb526SRmlNPEOQZhHLrNN0rc85u3Njzw
81+5rRNTZac+3HA4BKfqvxOs8VggMSeoZwat+/kvIaqNzvdrG97rc9jwoX8yEoSk
DI3TiXBfQ9jjn7P79Bxw9jyLDvKzu6vtuSOAGRURNWYxSeHPwkhIobe4KYPKUcml
OUPDtGmL5SpYp/Xh8YrvQo5+Me1lsm1en/M839VtCGYucI8Mfnw0T9bpCVgj43ax
P/1ikPSQrnC3f5Sh68CLlNgZVl9udq+hP1tI2vMLtiJLPnXOAm14o0lbRctXz7gi
jZncUN1bfg3cuLaEV/hA7hDHv48f4IK1TgsQJuzISLQ93icyp6jDFvxIkJ+a6CAw
GOxRxM4nsIKrv304bkYR6Wc6rY67rSjoExNw4OkcctpHrC0VXzXXbuLBtkdx2A47
tXxtOyJXZOLcAUuSIgftPZi9Xa5b+8FKnSL9mAdGjVaPMaGETorOopc9DdddfcNR
QN4kKhG5SgWWzsyhVLSAvWC+GdrmR12+ktb/0Eg2+MCJidHcfonHEl4BcUSaql7+
4p+Mmek6F6bez/BFYwWILQtnhT56s7ktYoRjkiwZe1gBi1dlkC++G9+NBtK4RQEq
aDBHwHD0b319RtoXb3fwwKrJXsEJ/M+T8uj4krUSawktdsHTiuzr+7IxSjKhZlEa
0ZqTdMZ2Cnl3CmtVXtU+6EO6jkgEcso7+9ZAK5ja2rbUTC874M+CbLeCy4qPQel0
CpF3KA9BvFDPiTbhyqtFbaAozyzkXbOsTjKxq9QA+y8CDFNzlTsN3Q1VLCF0w0YY
E2MoLXKsAOWuymM7vvrHEqaM3eQDCDaeELnssSRHG9aqVAvNMjgW12AXeySTH/84
kLW+hl9VZ6aJcEnv0KrCV+WHYyVtwITrFH1uNp7ykRe3mQmo9iFyHE6vPQJQP9qp
6DCq0XzQXXlKxV3nR9Y+rCePaTXYOHuxzixHzxTAWFB/6m41bXOkgwNIYh6GmPB/
vdZkhdbp/21oaL/rHLkQhudQm95o8DWaVSZIPEojmjOwQQyFhPAVDFFCtrjY3I1W
hic4lrLTi6hK0/4KnFW3wIDKRocjx+GNzzsQFbtNIYZIyfnb3MOklRwYdlJrULxI
weFDILnZI98RZUUqzz2hEaAC9OrwzrPRRr24Id95hUJR5ft7uKmnqQZT/U6gROnG
WMAl0AFYInqhhVA1Ze7h3Kmc2mIv2XUY8nPTPovMk75a5Peq6Mnf1cX/FlP5qthf
8F1ioT9Gg6S4o6giMul0sPSLiVLLNF3Qhc8+xc1OoTrDI73cbvnjxhQ2W+lxEhv+
Fgif9dmf/ZxaHJUgcm02sy362Axgk6gyMv5Jis06Qd1wYNKM7OpHGvrzTiBtv7fb
dXeJjXwnX82LRxjxFRsk9C4xaKo9+/ThIuM4przxNr2bHsf9dgv86iMpfuH7J5Rg
J1Kw9m2LCcGU+yoRkwJut/ERPUgDwtX0/+dKYUx1M0SctwHoqK3rcYp5bTSu7v/n
fR3bjmkvkLeXZD4s1zR68Yn5V7hmI5An7iXIRSHUQ0GE3kEbq+GZNC1bfAQbYe4r
IBw5oykZgnzBY3HMzsItJIHf4gBsmMhcjz7DddGZVdAHOu2dnHo/FbInqMRObdhc
K72FAyrfe/a6d94SE6KvKnHLQKuF4ULj1xFTe1FGSiC/Z17DuGtxkVqrSpgG0be8
XUrX5FPr9l7nzVZ8BM05Rz7Dl4r6U0iFHqJcBI5X1/jOTp584bUrTfUywiPADlR+
Ep6o2axQYdSG/I788MpC8fUT/adZ2zYmP+DROBgv26uhS5msI5OwlonwW0taeeA/
pItx+2Jy79nIY0xJjFveU1gXtgBuZA/Ts5rtm5ezcVjY+mDs8vhmLjra8P6pm94J
3ELszCEXL6PvLxxHlS+8G3uwAnf+zYhlFJyjuNct+co0SMG3dDWvzV0Ap33fl7jp
YWEJgU7Pb6MyUVizhCBmOFqjQna56vqv48M/MyMlxdGoHsj/u17fllcaVRxN6H7M
sFG71YJExrIV6kP7+QQGmDpvmu7CrK9FLi/gOoH6Mw9wUpEUsINYsCOSIiGwH7Zn
MgvEBdfoOh3CIH/zg+IvLQp+WrfGsdeKGB781LUj9ajXeq75nFWFeuhmajItvz7K
YMmLGRY3NpnDyJFR3INP6qmVlqgSBFHsR3LqWN/lWQUDIUtUw0YIXE5XEqxyqlA+
NE4Un504203hVk058MfRpANMH56r49K20gJfsDV/Hzk6iiJ6z8sJSYCN6SbyAwD+
k7//dTGcO4hgAoDQTokbqEfF77mJwybD1ebLJm5YfZZdVuAtSl/9Mjd0jUgH1M6H
6u2pGWbUD7z+fjBfXA4oHTlOSaiRdJ1UdZOeTZx2S1iujxigiJJT352bC3Jr92CL
OqGwzTctK/Fz3GXhIgJX+TqvORkMTSvZzXKPtmIH75uB0pmCs21Mn0FY/IeNkf+m
tyHnOKTEeB9uuhb8e+RImH1UNUXSAi8nNidOAKK1INRwG331B74pNVRBzQlFp8J3
whN1Q1tmSFMLgP/eVuwAgZ84aRlFNwk+5nTPQefI3Yh2qux/jByLdgvAtItVAhXP
Ty4ra04uHSxbJ2lbi0yGAjU39RSlLmMUdYGkex4I98ErpJOtY24g57C75QbNvWRJ
Xm5Z7pzowydNZSLLcH5sPXN56EhIl5VlDqNeCQLtt/8jU0NuIUCQZOE3VlMQ6LIj
aI+HfOhGMgbjuUbiOtoZpeVJcXCMuD/KwZciRhNsE2PB5LXQHGe+Cbp9Yah6A30T
f7TxT1ZpmqerY0r2htCmAVbUZrP+ffdTvPIltIethSPObbnmUsmmTbqOa/E9PPyq
dD1m9MxFTqJMV1Zy0KK2+Ls9Cmn8yGtOTjQDgTL+w5b0IxqcC6HDijNi1GB+LiO2
g+V9cOKkbdnNNocZEKklCt3RXSOUfqbJbyHpR4Tj8Cy0kpt0vrFJfaKUw/ixmIPo
66gGhYKigoo6XWw3Qt4tqTCc/d1FnbdsnZSAVXBrhxnQURvk+K5c2Q81/ZFE0TdG
wQaDPZlaNAFCmEv/Y0ut0LwZU2fll72svyco19GfLl7b2jwT4agpHPLK/FPomR1K
URyWbTsswn6qTQHC7Rh7II3hnAp39JK0xU/yaXzKnWDZEzn9777J5k6rgSfKtlCB
0CwnDy2mnoGbaQAcTbnEMoGG1DoM4oa68iltaaB8Lpwc/QiNk5O2ZsASvd+tVWrL
QXzldObnmJThGd9XMvug5y7rBHlb7kg2gq+A25roJ65//IJX4U4pDqESDj5dA/eh
Ku00W5OJIo6oLiNw37RzjUxFuqNYn1M1REl+aiew/h8CBuAojlTVnV3Yg9gG+kI9
3rX1IogGbwja/U9EiRSsK+fPQs+abueiin8CfjFEgoQ3Si/0HG982kkdT4pUuuGX
UJIa90Ky28iGOuYOUvkInetVR7RhsJOVnXahFKttfPbId3Sg+7wzPtz0UbdoujfU
2+O3FJJfnb2pWHuY5RRDQbWiupEIx2E1FuIRbxJxbdrHJs4hCjMX1xFjdo3v8MmU
+ka5E3lyflWT1WFCGlSMOAPhPtmPejit+J4TbiccAEAZ0xyJ2nxtuCkrVH3JXToj
k4KEMrqgepXsGxtm6uZkeoYp4yD8wePiVObQXi3cLBFx//341rCo9r152kWhO0ph
O1zNNMLzC2vL29OqLqVFzitzIDIb497DAekq2r2zi8KXczXxvam346mz50O4hwMK
4PQ39PXR+TakBQLTbMxW8eewPrmLTLAa1Xm1ePmXSCXBfnWkwV7DtbSjEm0XBzGz
Hln89vcbvelMroOZLnMKAnqgqv4VCGFsQsTDa8BqvmMnroY1JdMjiQDLrhNejp0k
Q360Tncq+XnB+3J679QkDDJg7rM7xmyY1WYKN8wquluRlhYNVuoSdece/MEQ/bQ2
xdRbeoPBjw9BbAFuwrzJzA8mCcprMj18Z9cLC0Pw7U+1IXoZZLEYM3DnR9sWd+Wa
Zf7Xu3zUi9brdG88aRFiBN4zITyl6tuQrPAp8Dn0vDQK1ccJg+xu7FyNgfAtzAr9
d4kFprW49evv9W89hblrOkO5mtd/Gmx8x6tgfnl/LxqeLaoEBsxxJo6ygSOOfWr7
dVtueMFLmZniAQ+LQsfglZiJfPOjmswqYui8ySlCxVDXLvYRX3CnZNaOGzfS1uvp
nGUXiPdftPlW9Md8i5ATZFMgCH238oZcLXSDdRxYRKkDL8V7yU01wHlivWpLNwj5
offHC88vfW4t5DIqp8xuRPxWez9NFlaworpoSf05KWreI4Uk5Ppxm3zvUp3Bg3LK
w3dWTDZu68i2UnyKFD/M7z4jAl0r/ioIGx4V1E7HSNql0cR/tE3FaBXVByF7V2ia
QWK4b6M8oSznhKXLQa349LuvLyckmT7Q7BY8F8ZvP1EsBSpUuDHMl/59OHma3JRf
hQM9yleV498TjcUfyMtGcCCqwj6b0F0aFQ+nYfGnu6N070BGmjm8l1BMb9h/wCG6
8zaQRVBMiUFgHWCPzgtcxk+UXRZvoFn8nigDz2YSSQlb+9fWPNm8PztMowJt5gHW
l2VaXWnWUaHoGYGcpadT64YhZdDMIsMHPGpYVTLOEbkgeAyqAB6rDADHet0xuhUg
YDqfu1TFDDiz3jFRSv8GkZ4gYnXXJxp199cHgaVCjU69WaCtfzn1dsLy/Ibl3rY1
P8uVNbfHP9W+PIGkOa5ejHgxA3KNsx+3HdFpA0LJ8HurseRErh6FUtCHdeU35tBq
yf+zhk8bMGj+M+1+JPORDxZ80IEn1YDJsig4YQBfuJdPO22+r/MOZoXN0JvsScd5
Gt65mQagCAW1F/F2WbfX8Pc26dYXFNGuSw9PXXskkmVCqfqR9/zfnTLaq3m8nCPD
hE+p6BHviHwktds737mGv/1TZ6p9CzB+h0VgDvxhuuH8O/fmMWda2LU6XbfHSVkB
VpdSxI3pyQGpqRYR74FoG0b2j5D56c8E2vLGj63eyB/XDn2Me5yYKOIUeiBKGKNM
lENhzCXuBReC6wPngP0qzKJFCrnIWT+7VqvPBpL9U9KoVe5ftXxjpiY75f4K3F7C
RUVfobIr7niuRTE6dvuk/7C3lXkplYvkpnbLiEoZofQbgIQsMz5/23nSUAms0HpO
oCLejIMEBdKa8vflZ0L3dkgDxbekdMGguCEdPFujl9YcDnaT+Jaei7u+MVetYxTy
5tAeFOKOFQLufSoYhJ7sOC8Cak2w4nIludkMjt2E+NJtGB1mkks8HdwsfBAoRpWQ
4HE/rb7dw/u/c0c43VnK8QCcAGkhbl4ZNPzl3zQ8A/7bl/vR9W5r7O5O6SouLCsY
ocZUoDhSeldXsgKT44NM5yIOfkq9SUmNkTVLQI4OcZAHWzgKW6UGta0NpnpkTqHV
aCVGTOEiaSpy16AUj4j5iUdObuirFP5z7LQZTT0BOFbCm6h7vFddtcSUSzjvQzts
hhk46FBeQ/UmLG9uS/4qYGBYMJese2tB8BnsKQo4glnTOCvxNJSgtpcscBsByibB
OPNQpSPiyqHlEcrDUoQRHYUzTj5u/II2Xv7HycPIpluIrVrd1Qibwqwrb+z9gJ7A
1KjlYf73yJGYBAaRDYPwzEYLWRPJLF2mJAomUO/k0AXPNU0PTjBNHDdNDNZTWQ6U
72/ckRhk7teRDIyinj780xF1BGre5oT2q/8/AJMPIIieeOfjcfkvSaW8JH20c1Qc
3z3Lqg6srijkKWuUCP3//fidTxp8zScPH1AhZ3osU37DLFDYU+ZP2kBSKrzLvh+d
Ml+iHRYiKZAmijyGpunxW+geZLKjMFAZEP/YMmECnhA7X+ATIbR28lgw8fjCoktG
ge9LzfCHAnJlSAI5ylP6OsoY9/LHz/1ubNT0C8V+onG4M/TRZxl9fQ5DxR/o/5dq
MHG5LcCu3zwddGbwnd+xNE0yq1Ik8y4wzDKy5Aqz/BExswiGTIDdFI4+O6h7CLEQ
3kipJvR74eGeQsgv77sbKXzXbWmbFwB7ME+HziBUj8Z/qoHsSVTD/TruW+YI6o75
V9ATT3Po1YvwG1qHC87r+TM8rUgYJmrVwa/8RX3JW+rE61eJcqqqB3qGPYdZQtEV
8eH59EqqTp7lNjmdQEZUh24MfMhko+KMJPEIONnmMSAHfpTGrvFsPDuNjWGgMNCP
ScEMDmE5CdBgFyJ1e9lnBmic+xXozT1iAjLcVZ7hfQFPNRVTdSPblnhZE8EXqzFp
ZOJ9C+7kp0HPZllrR8bBSdcHxOa7OgUbeKml0vTL3FgLgqLru6UzS3hTIKnb3sPd
N/ReH1w3odJ8ZXg6QPCTg4naGwxBZxdSJXJnX1mRDIwiuWIis0W4hWh7P13mPNmF
I7cuxcSt5OaSZtJW68tmEEj5OQxveuNO47VJ/uP2xX0o0gKUMZbYtBuM0YDrI0+9
Ip9+7vi6ABftPmWjDOR5roI/AtoYhiR8Q+rSz3gyLZ1fbht1kqlvN4nCGqd17Og8
GUWZJAlLBmfk7Qms6Ym26A89xlD6sfpPAB8wZARf3SD5SwdGrgs8lt/mRofXvRw7
Cu7R0TN3u8dfJJChyKQQTHshkdZLkq30ita0Qj6TZ+smsGuP7D/u/Er5erqX9YOj
J7rLPIcnE97Gh5ckWpaijLwY3T5YhrJk4yQltPVztKJayVj/alyUat//ZKpqgoJ6
tXmpHOOdOlg5u7+ck90BAa14F+XPQM2bWrvNq87huukeZaWnjESBQDZrDxdPlEZF
aZR4GNcK42sVnDioM4eHnhOH2k4Tz8zdoTzlJtdHC+VaK/M0xq5eYaRHyDZGYirB
gmIcZD2cVwiUE+gWIsGWmql5A/bGJDJKYVXQeWAu1DrE7jl0zom+Z7LRivlLj+t8
XyPoe8Rf9G4QP17ako3DrtS+iByZ/zkokoz0ZtGa6FLBrIJgxVBc95t/AHGEDUT6
If8jwlN9SDZo/uwst0xxUbnByB/Xf7y/9upKa+O83OLDMB5USa+jSUVi1FMxdHM4
7UKhZcoJwgNEYvNIYVAJxpq/5zjSnNq+iyDoHDue4ooq4a78mHf4GIC4zjjiQ0Gb
+kWBlqOpez0ew/eE/2fCxBL/eIpa//+0xTdyVzZCwvCby8sHwCo5rMFyDVF5Y2zZ
y3QVWggYaT8Wj1SCvz0HUMnZfnv4Smwu4T3oRxHGVJKdooQVWkCJIdlgPXkLTxYm
8OuVKnClrETcW6AD81BlwRw1x0orHv4Gb1BwaVUEWF5k2zzLEiHGZVN4CnGeBibI
4dRM35zrdxwQpF3tZY3DSV40SWvm/86giI10ndrYS9M+Nv0hJ7duw1SeWgGwfjy1
nwYuqDVSSTmOAT1uueEAL/fCnJ6Z7hOCtSL/DQ9ecqDNxnn6oAiLgvkCKyVC8Qfl
Kr3aloYWub4V7vqTJXRD6cn8i95/be3aKoAs6t2LydYfKlegf4oIaC51KBYXMSf3
C9CEjsg7ECYgMbcltcC8Ev9hR13238b1osmymJRqUMkbZa+fuorfdRzXsMq1H1N7
P8KSXmPFy75hrgPOohUeH6TXDsjlT/KGlmsv6tll7mjCHnl2O8RNRYLu1HzaF3C2
91VwF6pwu2ar+lElk6FwWJ3JqmNf5mF8Z1xhPRytQLDHFTR29icFqFEiLsRj+//z
5C0SxLGoM3r8XAaSk9c9l3ZXxD6proym3V8c5E3yturgFg663VticOkN07gFr8H8
F0/KznSL2x8Dtf2ZN4bM9u/9ZkszMh5dKU+eq6pSZ4MvZDqUMripcQ1thh/HtYoY
fckeanSCGkJGT5wtwsPQ3pymwg6jfSiD96X6NOIo4xkBNsgL6kUQjCK1ifpO5VLZ
qtbB1s0h4O/gZbHSNJJQfR65c7T3L6RrjHRrcgVlnamwjjc0ot1NETgBHZW32Wfu
/258BX0R0WgeHvDpDtYi/LGtdZHv0DYOdjeg+LlZMXRwcxIXubnVUndVzSSn/+JM
TEDwWjg+Ks4W8/pn1idROUsdE5KeA13vV8QGlsRcdNVeYhghFyt0Q5Qnte36nClU
bY+ztuBJfgZjupRYrM6gND8Lp7Umu7STArvuxJ8HXdIK1qQqqWQ6fNLBUJYDmUle
MAszgyDRm9IkyQ1xoow7RXGNuTDAZTrrsonL0PAPryXuEOoC9m1qJuAFFCnOb1Zo
svAoaKmIE5NrEarYViLhHwYEIQyq5VzE1hvHW7ZdCTQse1AIVGivClGVRmisCltd
ZyyHsZ+61rF6IwfSysKRlPAsOYU0QQRCKrvthRF8hyoMqhDLhJplvkhDAKb3N1e6
anv0M5URkgEYpLlC21JOZYBFBSX5Y0S4t8lKkEiK5prEe4RVIinLLlZYTX7uicVX
YQ0sjAuH5fQjBPJV5j5xFHGqkI3p3W4u/ucH5YES6oQExkxvUWKYMXg+BjIZI0UY
ZwxDRwFHXYR/IsR3X9dh5Nu9pazX+DjkDT50dMX1X3lRp18Ty0Y6f4Zef+nMW/je
gx3QUQITU9StAhMc37sdC+vvHWy0EnMFBiyFQVN1m5hjZqZ87OFBbVVNolw42bOG
uAaKZyx0N+RtPY//x22n96TGbp+ctTkxx5PsVCdhSAIM3hAhV9CIm8Tsn15mBE6M
TZRkJfEXYlBdaCGaussXPfFlImZ4PI/gR5kOuFVf0EFrc/0lp5wJ0yqy6dGSrlB4
PRw5uh6zqFEjgJr4EAC8cZSlS14O22P0RQoQ+CW7f4W9RhcHJInWOiQ6dLaAwGh7
hDKl1yxKLTak9HVOeBR7fdJk7yxVSHi9cexqpWgZaNefm0wedcSjr/cPiaCgqlFP
DoC40sCa0Hpl8pL5xRV5UQihyhqWJE7rSJBwK1Jbhw8kIhrarwe5guSwsdi3RygP
otT2hEwtH4cmd+fa2Udb6NqgMw6fYmOjTMltUIzPPbCGmXGabBnguqR9aY+82Gvt
UiwfZHn/EGrBgNBqL/o4LwE1RcLFkOe/M0ZH1tmxACmQ/GeD5P2dnCjhn513/wkd
ZHqMdX+/ayQYTnvUi8+vO7TeoUZDfTuMlijgZ/FGlLl7fRY6cNpCMs6U8W4RZooy
bPeKDcBHQ6dWvynVp7vS1B1SUJZzyKdM3GD8/Qn6jt2UNguiZLkj8cHNfUuzzlx1
LZIF0C+7J4H0hIx4v4FXCXQBE/WHqQwMPL8xKgPWq7yqNlcuaU88JcH5Xc7BMUw7
IIGyao/bk3NS7GMFwyKr1vvWxV0u9/JHRhhx+yyRU6kFwBQXcVmxQL0On5Cb/AvF
tuMTDlFvD6treMcA9q/fF9Vlz7D76ZpxAwmpu1az83phXuiTFJpXfJy4WsCvz3hL
dk29UkYGjZXJMOJ5T9KYmZHhqSrobdzdec/2Iz1hrO4d0FJRMdPqcRPZrCqefwdD
sHFH6LcopmwWHtO9iVCYxufUJOWSdMEqTQlGUoG/S8a5uk7u+dn3ltPTx+DZN9vJ
Rr72LHJnY+LyWxhL1lTGGeFBpFembSWj24PL7BYGmRdcuJjPVFoeDpPQV4p8ogFF
H1Vl6Y6NRDXIOxbdz81g6gHg3Ng2iEzMMsW0yP8eYKR7gC/nWJtmUW3OkksdZGmG
GuSWb3PxuqF7HMvJ9nC0TojMkEyx/HbzC+Rls3rxffWMPib6rgstqbFrcAq6XOoS
GPgXNv8/EptzlNd+cA5lDohMzePKlNFFpw7Rd4Q1m8oVQ4c5IqgIvHHDXsn0hhZe
/16z9PZTdfFMNEyhdkoVDq0Niyb18NWcm0W7uW2GTmGI/CZ//hfI8ikCOIhvJI1Q
8PBW9ZoiuzpAvRla3GJGv+BdR8DrP7CAgwBf8wR9/2ovvrc2krXW59pA28DNrHG6
g+WOi5y0sPX/d8zNGJix8qsS3RLtXpzqEZu9E8d+TEtFl2cBIo1TMRfyywGVaqna
WqEAQ8D/tcyZPdw439EAra3eI3Ne6cTGQf0qvBkGmp+mmFTEBOkcf6fXyZDqg2A7
THU3OSBnqBClgfqn8BK3ZfKGbT5jpIeKJx9TduC3fFafrtkqYl+DWnY2mYDiWLN9
5eodeiEMpfsh0mswgaSMrI/sTGu6qPQ24epj26mNYNnMoAVWzqC00nx8dGFeT3hw
ZSQpU0B2ToGJrUCPhDbK1OmtMgm9LI7z6SDKJgjyVLcCVsYuPAJSfq9Fmf1XEc9J
ZUdBuLDE1l1o8fqUN35W6Kp2IC7NVj/nniEDnupEVcOUEgH/hryz2gfLztpCYy8h
UDwIc8laT+m6iuPb+BMVM65UTGmTC4H5WuGfzkvcqRGidUofkm84hWNy5jB4SrV6
T98fSHrEqkMNL0/vCn05fKDgGkC1NU6kebFOTiZV8ZgmZYb02h4eynmr6+bN0nql
WlGIVlOw0YP1uRVMjeIxZFFXNuh4XCu1NFbsaY7IvfSrZ/Cw/AKAH2A0CRBRKSbn
TmioTpVemi/WWq2Rom1BsnkGXelyxJGjclE/PMHHFFcc4W5+C4IWPMXiACk6Qmwx
jrm2MTkLDiqbAOdGddVAnYiEuFGSq9qwH4ZRU/fDuCmJuliOZ612EmV2SJt/3EtK
JD8atpPLEe9GZWkewZ9bNUICxK+AzVJoFHLM6WNuyMRhiLiM9FlP+AAxwNz6GrOv
3hd/mFF7Gs8f3SVtPJqpl70TZ9fao+POmqbrAOefR0Zxyqbu1zNey5ogDA/AALrg
SIhER/tSL3wbzaysFDgygnJsNc/L052wWZtQrr/0+arM+APtbth4ruW8/WhISrBR
zpo5Qzf5DnNDH7zYeythmQmEjFkc01N0UgkrzbOFoi36XYv+ETMgMRYTuibMbP1k
uhvF5+ibcSbbPjGs9aDc/yRRVpcK5VC0Xg9kJhcjca9hiq+BFE0QW4snbg6+jTAH
fS5+dQvA9MpMTRXU46VtG+X6xtjSnNSDUyEWlbZV68mShfCglDkRGm2lcjjJfP1h
H420SKqmu05AGLeJTk/S56i9T4FNY3l1acuK8iYN4jg1L8ECGgJAPnwZBgRZ+H4S
0qDSQEY5oS2v0wjPka1cN4Z3g09BfP8xCGvyrL2Koi8hD7nuVdPu+OghqITv43lU
Z31C13HfsKR61gBENxNez8z0BSj6uTF3n0ToyH0qfn8rk3IM3kA9kwmwuqr/6lKg
D92l65JBRYOioR1iLBSwiEEceqHg0vS++PTMqDTPkP+CEiOofiWM/hjoUDyMjZlr
LzUVjvIdPQEyIdEqWLa33qb4buV6wRyPza1podnGMdD7GBtnwiaBGY8zsunKff9U
Lie6y6RXTim5SdNyPXjUOxUG6DG6g7ZbImrVE8pz132mJ99NnBjOpc1UE+dNp1Kc
u9SfTvRigCcemxlds6jvY9upmmX18Y8zSZdR07DXCVqhMPJMscvObS3LMM6CMifM
VcN8cAPMICW3gKalRmrSe1PX22v2WGXp71wu6LwQETdef3dRAnlN50CqX26Ik5Vx
8OFAGsx7c2JyVPFDwW2KIQbJWW0ziInA7t53trasG1w1bUl0/EJEx8/qraSVd/YQ
tScZb2lsUoFCpUcf6uof4aCE7NQVaUoN3pd/5gmogE8RdHDxolsjl26FR+gwGIp+
1pvSST0nQhOmlgOCc7hPL/COotKYq2oJeTB8yODPYRDU2orYlzOcH+tqFSgXZHAK
01I4cnFMxiYLBXXquZ83LRcgn6UDm9t0bIvA4hARWfgebj2AB+jBZ2dlCylj9CQv
iD1pBq2pTNYGP0b/OWaTa22S1J5Ag7+je4GaBKAArJh4Ux0x6yGIZO/WUG+UNiJa
jkSLsXcz3dm23g6wWEZz89CxMcLPACgGWIRyoRO7roavrcaEo3tkXiL0EGRpkmns
pR+TczzVz1EOEzuG042pGfqf8ST8UP/oOXpT2eL4IkYpTb42wIp1u+9XIk8YUUN6
c1Btj8bqOKDhXgOli3HkGb5vfSpi7uUSMdsrcbsYKEO4pCcF1mD+8sw1xNRY++Yi
mSc+6FHCdAtdtbp0HqnvLRI4iSnTg4Hl+p5agm3BgDxaZEU/Cp7Qk1Bhz87N0ZP4
BFDVTLOl02lRawM9I9m4s9wvFqRc69DJXArjs9zdf0n6+jsoJe7Qul+jK3XZPj+j
9G1uNGoLlj4buJNG5X6yKTnUy6eAQT32tdEB2VQif8/i8fuORQtvpf9cNC+CuUw+
WxVHIOdS6kOFJhYOMDwT+KvPVzISyBBJtLrP3//+8O/myvlXaryA88h4bHwn7beC
IlSmZa2zTq8zjSUallneBuiEuk81YL1KvMfbngq79V6qaHnB7OajvcYV28YVd8gI
/p5J2cjJ4aZOl42zr8rvLvtaDnSk7u1SLdoOGwEWWtgV+0gu+S6T0Jx4ot5I7rYW
rFdB0HIV9HDFHoW49DQakFoU0rDfTPVNSFs4J5AHXmnw7E0sBNOyYb9T5zhPXBxd
41WXnPPe30WbKzq+3XrJRile58VyXv9fKLhdeN0p6h1s4B75Xlfp6gVg5X9F8f/1
rpRkmTGb/R2xE5q4G4pezEDnxbuafQyPqVlF3Krw7YqBwGSp5oRZujHcmdpPB40u
h3Y51LAH+tL1B561fRStXDOv91PwZPhmNxU1qFAfXAEAo0cKxCPI/TQofjMl3/cJ
DmaK+ub4hhGef9jVRhns0IaodMNj8YmUAk97LC1F3bBi7ituzpiYdqlh6aiGrGT7
pclLMAE7vgN39Brs+Ltf1f3SNrYhafzmzX7sI81zQDtfKm3xpoBhbgzL6nBgdpJ4
EdBlk/N9TFsdM8wb7I9Q8C1D1m+HXf/158PT/KD4dLKB7jexFJZhq9fkjhzq+tM3
gR6TbqYl0X8ae7ZzGKmS+moVDJaRer535AWmlcoMjPOQVgKrz86/PYfkr+8zJ2pP
yHCM4piW+rtLCxsAMBvWCrZX7P3oUaVo2f6hZuaKKZCWJJtiPpGrDuO+IO3CKKzt
Mg7ekukU7LjoFXvgGxHavtmOV8HJxHvRoRJ+AD9vbKBHLU4CTfr2J++FPC8OUPqe
9jv7LLXCr0EuOjB86mDaPPeRURA9fsuXAavwroiB7zg22NY3c3rBXhX8seu2qVww
sdAFuT94dqfHqJifKu9NvCHwpfW1ezYbPfijP7UQT6ZAe7+nae7AqRgazUB7CIbB
TQOkmQ8g2MGPHGEG46kgK+Q6iaqV9xbvo6dhf3VZUfsNjCnJWAqqc4Mu1xG6T9pB
hhA615Yk7JoLo+vAWUE7Yv6warj0hW99kk+oAlal1Hs1C6prQ8ke0DUkGlAYIubZ
/4buSzG2vPshWEfow++HAS39YWDPZdLMeyfVXBSWPePzXvvjrJubKWNX1KmIxU6G
8m3p0MbJGBeovoELtk1CfvN0RSH0Jng9vL2APXM/4S+4P2lBcUNKvJrQOf7Walzn
dYooHWt0HVzJ9Ni2vXBi2Y2eDv7+ShkFr87Idtn6wPWlOB1efa74EVnWq6cx6qTf
Pu7005NkDlZxynwaSJJQ6qAIZ4gbT0HJQRxzRu8DNEbrn8+FVSNwNcaQK01Ww0ro
IRikyTm70jjINE3fdT+AQPwNS3xyWIV0qGXPZKR5DTAnPCqrsB1DQZFKGkl8Uqdj
6Xar7DHSs2RMkdyBoMat6msJjoZTRevlArTxwBAhqWsOFIfpaBapWeCPTJKnMvAq
/2tUWGa9WuLOyGVlV7t5p22Z/neTtjuY0uqbJJbD0ClW9DI/reXag2mW6TWrX0wY
ec8/Ce2E2SgwCi02wh78yCDcMG/bR7pKOJeKHCdN/A1EClKDU9Joq+UVOIN322pp
n1qgpko4GMI5PDvS2UtuOyd3s7QzJS0BNTvsf29bFC7irswW2I7E2MeKplK05Abm
NWW82gj+kkbtmoiDEQ+ZVv2VhwvxC3LZMhdXoZ1Pofujx6p2zDVmh9R9Ojxovril
KICYoQjiCqJA51Hu6S4YIOza1R946jP9lCZjt4qyF3Rdk8i7vln7bWmDnvD9yweC
YeRka3/soQksvVirXAiYb8Xe+bybKRgeo1NhtgZnboM/zk+cGRPopfXjB+VKCiNL
pwKqbwhDHL9sv/ARY8fSFBQmG08pTwJs9VzTqsiCp3TDty4d8We9KgyeVswst1z6
rw29hTrdii1skiIEELvvefJsQbO2ncf7tJfZKu+USVkWUi7tIJVYx5Z9T6HXMXKB
cTlFhWGrYUCUuKqWA7TKOCdoE9Ox1iX0RpRLchI8KZIlVFi0byD5L6bZIi3JSNCD
vh5+HRBS8JLYLX79Qf+6vHoUQesJDy6N8yhpDj0KbNDDj0kxpxDpu0zNOUe+yABa
HJOhMakzrbWJRn2U/cuGoWHOcwHIVuE/krdtiBjiEbZkZ7gMq0yiJuc45Ufbq3sR
msWMeSxuDie2eOqHCv9dm06mYbMZS5seasDZCoOJp+1eHiMhDWuKvQzGGvSTKu5x
CepxtYcll3EFizIm9hkCmcF3Vb/z/AmmB0GP4t/Wqv1NrEfwJiqGttFqHRYMsR2v
+xAt+R2dQ26H3onQRnpagtg/vYD5XLR82rw4Uam9AQzeazPJYhhRfhxMtKdTZ8/F
mrRRm6IVvg4Wg9s+E9cxrGxDyIBovhGo6tQQp3OHlqu0kRQpS2ABW1NclTvCxBOG
i+5NdBGORCQXPyeTFH6TRtb5a/CSUrJ0w7IAqgXrXFkfiGOCkS1WT/aAExT7jYhw
33gcmHXPIAdAM9bFXjCO2Gpk38Al9at3XskfURMiL9KZ6tKzLe4XuDuCJJsS6CAb
9vSMuHp94I0hzKUwW+9jSpJkHc3MDmBfncHcku0MTpbhWysqCjPFz5Zo4+n29NVf
fF1123fqjB5sREBCUFrjvaDZ6j/oojKTWEFhfX9Sz53dqEZn2MMV9D78sJcTMFJd
ecHkFxxcvMnOKa6q0rqgsuQ5OqqFIwWqGJ0gGxn4RqHBQifmOHBwT2YPpozq7ZtT
LWiHjbt76jKDd7fOKkFz5jbxDYMWzc+qI2NN7rBjw84DtiEcw2DNE0DkpzZMmpKK
GXjn9hAVWuOZzvbbggHLzbkkYlphae5A9FF7psDm2OQKfweFBQFIYm8nImgXlC4l
UeZoc/lfd9OP1hfWLvn9J3OJWUhUWYaOM4IHXLeqpTisC+qa5PahZzq9QVQ0tpeX
MwpgVrkGOcbMs/xhJ7otrDehb1qT5cVz9suXUUGABZSOlosn9pf3FqO5ZiNnmuCa
ehj6IYegjINQfx/HENBpDIEY/meKvC1CEMzqf9dobPQ8ViaZ8afYYrNmmWVDGHK2
7Uug8yY/2JfCS8QFf3lOIg+5Be1W9oJjxA1+AQxVSmE5mktx71hCHtHfCU4M89eC
bM/v6durUXISCiVw+9WoNXvme1eDn9+IzxReEs2/REEOzzdUQt/0cF0MZoaJAfUQ
GdacA3WArk4gc4EMnkkMJdTFDn1l6KnWnIzvOZT7bNLTa8ps4J9eRa97fcLuHf3k
KAo5NhZJZv8D31B5R/pkKtIN9lrTYMiyFPiDvLJ2MBexfGoPkvB4s7KU4iACnIJV
peeyYMcRNJFdpYQo2XzXbtPOLHtf8QFI4dx9VFk/QEYscDhQ96oqnX8gz4eB8GXc
RuWB8Gw/4sitJzoKtgBLtqY3pVuyTT4JJNmP/Bp2a4GN/wrOYpab7qxYJ8cumyPG
wgKdvtCAsAzowKoYKy68iWqnhAeGab60tpk6ay3jl1kCPaEp3gd0DgH8lgfauwmI
uA9tkgIXxWG9LBQALLkgR7TmU7sBfUBUN/Ya0lkXge+adOGM6iw39yRUiUXe4KjL
Y4EZ6NxPajJxYnUtBgBLsgMnefMidLlEyN6taS9/d24Ap+7NTL/zUCie4cp4P+dd
82UfDbRJCcgln9g/IQATjKG6wlqVMeRzBtjcm7bNnmZnBUtgf6/5fxaUsZTjwCRL
0um02lRKVQ4Cg7gDTlIqY7coh3kHPjYJxh04DvmPcLlKq89nDEddTn1mele9qb+N
NMuGQSQ4Ei+aLeQGJO8f5/axiosOqgN+nzaUvZ2qeeYR8ZF/M1oLwmuQnXNISLFR
mslwfQBou4BGCTYwAwhUHYzaGatucSAfALQjgL7bIJZaMzOPeTX/q9iojd0zeu5w
ukomcsgEostGoovIkbBvkxPST4yOvBAaWPfh02r5mxpfqJMSNOdAYqVr5D2KDbas
7QoT6SEwskmXxJ9suJK1XS7Hji0xBy4jlGmutN9PhP4ShLNe6VDjc2KAT7p73KGj
TBJMIdw3BZmEVThJxUtHdVM5Yu4limoheKs0MGsRiQZKRZll1X9EqG1+xQX3Rsqv
thnQUoPLVwhR8LpVkLlOBt4A3i7zAqblDq49UuDSdbCruC7/5zjsA2/W3oqFCqSY
Veox+cFph4dzG+NgYK7OV3E3yLG36u396WC17AMk0xeaMYmcnWugludaInYCWxTH
HRLc+Yl8py8zIfTJoj+I6XEH2kwUBoXriLabnKvuJqzaAeQL6zkLc0MLV5H0GP4c
4jGqLSQNJ+iOhV9sXJt63eGPTcj05mLJFFhP4AVQVOMEvMOqaOPnaAQKU3EJ3Jmg
rdBuTv63iAu16pfK7j4RwvW71MBpvFt8X+uffJveJI2ypIE5lfLP3m5ADKF3B0vM
k8KImZihFMvrUpvkhAOFEPNovhxCmYjW6IdchSMoTDft9+Djc9e2zgD9reOuOPkO
CJXjC8uHlOaTBlNlZfxD4JiHFRD4Ep8gvZ3HDrY8/OG0Xm4nUTL+brt7cbS1Eb8t
LMPJS9tt14vFqpl3ZoEOWwh6diDAXcq/YO5u+PZV//pBcvIHfKF9aizMFERGVd8b
7A0QTQJftvEfiapv/wUlA6M5jV+5cByWVjhIb1BzeVcyt2VjOqpeuT+BphMjovR4
pfcWJxi8uf5WsGl5hkCJzFQTyJ5Zok+s0pT2loCdq9HMt/FUzpb3aMPreRIXeCk9
cFAswmYvRZBZTUzsE69L9Izt9L5KjglWQbxddX7PHyEphPY5GcloI7ef7BunZNUL
aMJ+olXTKckYQsiQp9xB4lX3tRizpYm3GQVgjy3IJev5aMzmMBd99n6/1pIwYzrQ
8bWcuUoohih/w9KOxpI1rLZ9MHt5d9nQpCCJrDYCOgLLyof7Oq9l9r4izvBK5GEX
/hbAO90HzcT1HieVVFKBrCkB0qb+eaXtJalzjk1drdtV9b35RtyQAiXGOPsL8b1r
JmsdxnMp5pV8gL+eRXCovOhciFeZrP8KdKE6nMZfD2qswK7wpdzZ/dFZnX61RWs0
KyFYsAeSifmzJxG0n90knII2tnxhgmAQN/VpiMmxYT7SwbY9oXaZKfXP9xJFpRN3
0opoP2wA30xeOLWSHSuVXwEDyuDRxumJw3hk30VKK0957KKVA8JD/S7U4ofYuTCz
BFT9wahrlXlU2O9qseqV2sUD/4XApds91jr5RygrLJFv0CrMtZCi8H+lc8y+oSeX
fHIgCz4wcI/EYQNGLNDwnGmtEpeKWnkg9lsEqS3Rp4Ub18FHeV2jZr6PNVa0jDh9
JuZ8mWHaROxInWOcIGE6pcjExlj9qLQKq20iby/RGmD1Hnbj0fcafiNot4FUDDMo
CFhCXurl40lRqr/4dONzSgHjZSRcyxncQdX4G9RK60itDOIUu99EJxAY1BvLQAzm
7nPrdZzkM1mV2pfLYQwDuQEFfG0BePYl7lRXwGlcXNy80CsRilNrqprpZoKi/zPY
gayjbbt3owVOpLqyKvurdGqwF8JeuEZ9bOBnrWKNTuKR4f5eHMWNRcgvsaqqyweu
UIvdjBW6jCYESAFwfH2OiJ3C7xqbx3lCvwUAVEIzK6yhG65I1EywZcij28XJSiCO
YPjK97IojmvOrHSFO4fdEMGv2/Bvdr4e2qxceb0Vtz3NpqzZmPotcurzmPPfFQSq
oi1EjgAYs8+OrhRkAsx2ZfOW4I6zVTl3LxlIAtnZnVVsSHpjBx91PUwd4NGjkls5
OBMyJ3JU2YcyjBTrMJmf1jR5RkFmgRO3GK539TDYZyThz/Ox3OLFH+biMnBzQ7g0
BlRJJE6zPWjZGuNDfOxqElIBu9m9CyWMHO0FQTeD4hv24ca6TmF+w3llrDPcVDAl
VlEkos0MVfJWvj9trOAr0Hs4LB04TJ9ECCS0Hez7ryA29B2tsV0EajJgvnWYkLKw
nT+t6Dao25pwUxe5+Kf0oN3IwYrJQ698/HOaPOXot13lIMr/K8of5+VJGbwwoWXi
5b0gA6gvodUkcnoh9tuuYXvRwCRafQkn3D2QFVeF0UlFh1YwpxymPee6sQJEGUWm
YNpFB+3+NVlQD1GeqB/k1YkBMuJmVlyPkIPD4W/h2uM3KWXrjyRaV9A91NcOL3yI
y/GV+3IxIEDa2djlMsdIn1365auQv1VEwKkKd40PPms6yjnEfgA5Z65dRGQoAm3H
mia3RCD0GEVuNdoNScX1te9j+TR91VNqB9zkXVM6mrSOtwVrrF9o1SKtuxyLXC7M
t3sxKIjkhuNSGDK4hlWeb+h6Aj1Az68/gHGzPQqDDaltgXnNlKF6OSA+uJLzhSo7
cz/UzRePccR4BYE3SKEBPKvMYlkHfkXKTxBS+wR6odes74uQUxAGD7FEy8Sz/q2/
GDxVyG5LjXw/unpxKN6f8f43yajyULXLTw3B0yh8Zm1hMLDfuuLuA4kRchCSNKAx
8tZ33E6uxaNYuWh4xzvg847MoeMbbcj4WdDVs+UVom4p13EYVMTOhM5oTDvOpiix
9aJcxSfkkX1rv/n8Dzox4qyfMp+yl1Ku6YIa0vKRuE4fKj3W/ib1y6YDwFJrhizk
3Mxxcl23sTV8Hdbow5MG5r/vuZm1gTmgzyp506ytAY3VkM/rwa04VfSOYIjcYLNe
0v97eaJwdyuH7kR6tSlunhNIn//Mk+PYhI7TIy93Znub58tKgJaHcuz22rOobPDw
3BKZpR2eSaxHKbRKTKXVp6YW0ye+AQW5DB2z6gYhGoMFjb1t0mmKwwLGnXYdSNhO
b5yemGuwX1iuduB3B2AT6YR1h5n4Q6ivsZV1E59eWe17EaxHkXhjGhnlQgfgKCFJ
WK0CYbNmzrdRQ7FBbvsrb5FZiwEEoBMfGsI8f+pa1a12jlYaykRkQpyw1TD8H6co
ERZeY7VH1jzrLBn0sKDfrFFUy+aGg1+zAGoXpVsZ7k2a/O1YS6amt9b76WjoFE0R
ML+Mx3PjwqtEmrWYMI60KRaK2ppyTwPMsiwK0fhOuQ77EGqGxlTQIEBfILpBR9/g
+WUI6tKe7pMKsHnx46d47jX9Ssx5mEPD8fqXtwv33YFARLtLNgaODG9DpCx9/SYG
jpVPD362mPBNoPe+gFvJlXtHoZJmuJm90eirliR1jnxd5tiGSFtjEI+rwZ9M2S7c
n71OVq234cw7L0t0/Bkt9Wi3PweXv2bGjPuXUn9IVc1Y66rdw/207u5268pa73J7
PUSSksUXRRU1nqEGd2l7gzdrl9mlp2Pshr75lptJBa64RwyuXKxixNfG3CRoXr05
5BtJCdx6yZ/6hCrUwyLo5s2biJfojy7PmjMJEHh728rYzO7MEBh9l60Plj9LlYKd
VfgVTqkuKx+pTBX0fcNmTab25M9HvDbS1I2Mmc7GiV/bxTXajd/01CXTTxVSjRGG
Jj7x+1Pze6v/nlfCNu1UO0b1ye7TURKlqCenMSACYYci8Ub9I8Ts4a26KdgCUfOl
4Ak8wcPi5FqgddwwciqPFkYB4I99KDDLAY5gdoOTyu0rBSWcArBX6N1caj0zsUI7
Ko0EUJFBxaJ0EhG5S7RvGK6c4JJX2IpaGSYVSVLgQ1JHZa/PdJ9ldwrU6hgz71M1
6mc6vyt3v7Qluxnj4qjsOqxfQfX6DIVvYReEShu2aEsCeM7rMlfGEnhF2T+kbWkl
n5MdrKM1iarxvQlvFDrrJlGPtkJvaabLoQJDqPflfm0TgtOxi86Z6toN9Vlz1/lW
IDShUNVz1r3UmHUcqtoX5sg1UyBStVbjSYD13sW7Nb/ZFgYzEZYxptQsFVeBB7O0
TGn8NMuvIBVZ1lFpkZ1fS57DV7s70LuzCysglnmh9DtyDDPt9oJaRbinfzIZn0qr
B/lFUnEpOj2fjwlw+2lSJdnl015k7O2uZ/ahlSVlp2XGDGzbEZHIQBb8EK0xX59T
vRv8I/+fwwfIqXcWtN/guJgHFC7lh8kNPZxi63f3VxWGplf5s2F16r+hLDmnZRZy
ncQDxtVT4fdHXYLOxR/sVdyp5+ZgKzAyMKGqjrtPaL5+Ap0tQjEc7Swwqcg7zzez
cIm2i3YvPXSOqEO4Yye+Agho26B65WsqQ+Y0mkxEmIWBghJEnltRTYwgLD9CUn+7
Zv6KSf/NWunxzOJMHqkmeiWljC1e0gCY64mucIV+FNwOB0wW97ohpg5/w+zx7cHw
JmxE4gm0WbsccSmA7NOnvoWBFegGU9ITFlZVGtmQC7S14mQK3Tu/f5NKt3RtXaLH
b59jX3IBjIqOPFTe+m/u2IkSC/7pKQkLXqyVY+ZsiOiuZKwlqu1NBzr5sRaRMuod
ifES+ADGThrbg5ApNGk53XhqlCxE2AdiZfYFP6zk1nuJ6fSs3oQn9YaCr3nG5z74
DPf2qR9jkIV4aVTCmNFU6TmtqTVyUURRNF4f27GsCZsnvsWDmcTrIAp/Sl7LubxQ
LLOgvrDs6DxwKTQ0zwwYUYbTTogPkJspSHLcQbAqM+vVzBfdOzsXe1zCTXSwXuzu
aBBw2rJbW9Asl0Hr5Jk2QEvfIAsZS7oK32km/0RmE6L+cwRO4GrFveEIMwqkbRQt
xNa8BM7oxGRcVKUnQ82crbjzfRNw5vb2NZws0JYD/ydk3vYxmFbidsBlxP2GwNlr
YQcIrpnEjCKn/A1r/3hoWvdQjfVTD2cuaykFS5T5/1VKQCdVY57mLx7jOjEXYgF6
ixEkH6gybjuUaDC5Tt1PUyTR2Mrc0ot1RzpUYT9mkJhpg7MknfrbcpYH4QTiJ34k
rkjSpJTcGG/bHyWbmrFzGBNCE6UJH0crMreljPJ/wv6BKE9DUcf0yUi0conrXnyP
GUVzP0KNjRJRLzt6n/ywnTm3zXQQXSqpRTpzwC+aTXpLN4gyjceNNSVrVZwkAKqp
v3shhEag/WfuWxmLoCWRazurZpcdsETF5A5MKDcP0SelLdumce7ScJQe1HRB++bO
gimYklCtWFY2g6O8UZEb9jAsQFpSeMTrrIM4BOd1CrLIjvCWJmvCOJhnakyGEuwH
SvyIMpI2pruls9VgRkZpM9c0EewFNYzP1lWDAjyJakfzA8cYp2F2jbv3I4a3kERQ
OIvFi+3J5RdqXX/dlPRftctG+wLAOsHdWInHD/VibhGXFCJDpKogWaJz0kJZWFD2
ZJlxxY9QmoufTJf+3NwJsyZIuNViKjBylGCUcx1PuUZq8oqhsbbgwLi5USi56RI3
BGJ3zqrOk/qwbiOLNBhJPBH/uuwnqg0Ld7V47VOPlz8S/4xJIlPH7QUrl1ygzfA3
mi9dbvH2lMi7fYyh4flQR+3UHSbss7Ufh7LvSGndRY1c7z/n7Ow0J54qJrtJQ8Nr
64CnDQ+NssHFjXiswrAm03wP6fcflSR1PkrM2O9gXizeUw9g3ffx52HM+UzF2zJQ
WSgzoHfcHJ8RkB123FM1pSjRA3B2/jSu0Ts/hn6+R2k3FjvDrhJwDlhHkI5t7nE0
gk+aS0RNrv3U6ZY9ny0G41vDHTTN4f6n8Fs06hmZ1dWkcqURUa0AZnVpGqk9/VKZ
TGZepwvaE2Pz7Vov3Eeve3Vmgilu0qp+sHMQtaF7VB5PuDg7/ZNnhQlTHKtElm74
KuCGwdcfSzfcz9RcMpOG/I7YOZztLnByUepdJ+NpYc4axhDR7+XJr/3hNvnm/Ph6
EFJpBzt3gjf6DoZCVDAgpUZkEDp65ljDCtzq1wrKlQgjszcmpn5AY59ha+qutIj6
MM51RQIqZMrWroXT2NrbllVbBbvzKgKuzcCbUaRuUXPDDPhaNE2a6soPCO8nuVqt
VRBB8AmvKZcTphmdKcWz5SvyJNFUHtyNg7K6WKvV2eDp2u87/29J2pytBFsj28C0
xycqnVPhFmahpx16p+SHrTXPQpjenIJ402UPmcG6yTP3cKSdmd69hr6o0lmgh3XH
1GBcrL0YSHTKjsujb6ktA3YfDtbcFhnRGiLookKi0IjkTosltOAHByjU0oOcfPaF
TBRzviA28OqL+vxDB2QKFoq+FKroD0AQp5Osj3ewU7e6XnRtGM+w+AJ6xjMPrPny
zpk0jJXnfePu/b5rrSISsVCuc/jo3dn6qmmMG70w9Yd1gdMgz0EY0DzSvj9gCkni
IobveRj/wFlPrW+Uv8suGM66mO+dYqWD4uLNqsUuS8ds5opoWmXAJeGYID3WkyAm
soq9KQPR8+35oYe8gOlm73t5ePyvO9ZQlvOqnY31AAqW/90fzd0/LDX29dACA0Wv
+OJTKNhdXIOV/44AqOTGyCGm5E1XajN8p65/cCHdcFmGJ/mN+0VgfQ81gEmexl4R
wq6m92Of2wpBgz52yACU7mO3n5MYjLsQS4KQyGhILqFzFZRMe7ay+TtfRvj5f5Uj
pNoanS12zuPMSiXk0UalxbHTgNeYhzOM5bgRLI42J+JDxRL80Ugk110jZJ3KWTp6
k9390o7uZ6OeSzSUmzCvOLCFUaySeJoIhUw8o2qD7hT8BM8ReSXNtMJi7tKHemHM
nMOZe6DKgTMxlwPW93fLediIXeDxMWVWOWx0H8JIMAznTEis7WDWeXrb6YUcTRSv
zLIWbCteR8JKmreY5QR5k+2gy8VMhZ/ocdTlmbYl0Hq0HtiFzaNROvWW2d1Gyhjt
JWQRoe8Eyq1Zm9+uxDsowR0rUzN6nygsTX/EdLi8iZqYGDoBHWMTrvdCNDbQkMfk
W98DMDV1kybcs/UtSrbcwAS0g9LYySiSRokD9AKkgWlVDkf66ICAINsM5Lwwzde8
PSvsUoO9y3QzTAfP+0ouOzc+jxpxtftFt6vj763ZDgUpgQxQr4QtKeuK/4agLJXE
ASL5XZFnsS3ZR8Gser4i7f1/fNMTjvfFHAWewhAd6nmUs5oPrWoToOAuWid+AKEm
OBuOOEIO37QtDmTBNR5NBtD3cql1rk9O2U6OQs2//r3shJqU8Vu3fg6x5v6tyskC
/Zl2k+5hHneDk7baM3rD3EhjcT6afwQF86Rct+GZ4gAXNqKBeCms1Nf6rtFV7T/x
Ez3RieBXMaGXD9hvkkh3CMM9T/LPUSJyTGXVvaXtnDTpLGRca9WH0kZgdn/hFxuP
mZNC4158PPhBm3emsCOPMH5FXNkImjLVWKzvOVds67maCjAvMDFgh0JfqdWXcM84
s5jc62owxkBHYfMCDmYWkFCTxlXpYZGNcdNIFx4tyF6gAyf7y5fEl51lJwZZNTxG
rD3qMpEvmQqJcSuVn7U6++g+DoQAYQcURp1snPiNQc8p/AL2MRFomwwyqz/wHaP+
wRkf8+X/FuVoGmyR9/pKg+g8jyh1v01wEY+MGnmBsarDbFAooq6qnUv4h2JDtm69
knBZ8w05B7B1yJ2DGJ5B3xROk5gNzUHfjiPfys37iQ2QATTkmeJ2nBouqpYFx/Kq
fk+t+4QihYySIOBp84qy/5/bRvIDBTgq+BtSMhBtDr/skroR9SBqcPENlKHd2n0Q
pKtDnv0a3VwUmh8qyRTswQQjsr8E7i5Di8bv7eE1ubBqmbwngZLdW9W13mcETMR3
MN3RzdM0fPGKIlhi+1gO+B4GClWyv5KShMh6FzagUIPKdHOqgKkEegTLSlg67IZh
P5Ek/NSW5F2q0WVDEh1z7sxbOckzS4CZ6d6kFYO01hBHosXK8raBIvZwEu3XR4Jh
MpDtvWAn58KB3VLvkQRgu+ddZqxQabwyRoZwzHGJRry+3C+L37gJb3PwWWeU3wDL
YSNQPHEtAsaizXM8fkypvCnGCXKIBumhC/vDZUiCb+2MAWrhPd39Jb7GYFV7MayH
puHw44iqWm5WOT29EWQJqCnJfpJVOBMTGI3q6S6wPJiG+2oqkSxP5oMcto8Chv8m
d0dKCD9FHjNISvNyGit1SQEzBTAXS5rWOUI3+IjB8/FZXDV3PaKMayTBNXs2LaBh
9M9sSja2FgMTJaS6Q3Wfu2nZG9npQ5QeQFZ7YcGCsP3Tn5cHcjOXzl9957907vn2
QXVJt8YlV+ug+UiZWuGCovoMVi2sqO1mK1LFevSIEwceZ+s5FxtWQrL2KbF02I40
R7huO491cKNahwwPEi4qfskbfRqPkSgjl4Ql/Nb7ReifMByb/HBkMKVrS/HXA/dz
eeSWDsG5B/Z1je0rpaqfP3rWsSb1c8A7KfLqgId/obPcpapbeymBMgV7hI3aTriJ
mQOrro4SeLZESXEaOmrqqGv+5MURmXF6XRMpJkk6UwCVZXRQZMCvuU/q23qRzO7i
7twbO+ahaA91KGyd9CqT8qP9QX8+ckGERbJhVdnR/S/CPKz/ez2fWC6klpQeCRqi
0HUOVg6QkyCvjJs3WuGPbgRLHbiw8Ge5DrbqbssukEu5fD57cXdvdqKEX9bgrcFW
HETlHsdBzyVillwFyY4Bis0gfLzP0KKs5caActjXcDcxgfW6OVWVkCLK9l1J5BRh
ETfGGlMdk094FJxmo0GEmfsorxEYmd39C5kVjnNqfciRSeg22KMsXw4jB8yNTm8J
ZKXcvLaEPl0no6ZnfhDcaTEWiCXr17GyORyIbxC0rJpNwUDK/eMTJpDc+uuBGFud
26yyZVHJG6mpqlrzy10xBWlBEHas2daVomVDwDOB4O57hr7tVvT8TvrY7GKWpKIP
m/+b3fH361G8/G4JLl9Sk1Gi/rZ0hwhs5tR/XTfF0Cs0XttuwR55sPX6kxXSJt5x
N5VG1Hz3ZISummvgBGPmfnTxilPS/kHVFOf9Qnx2wA/65e26T6RfYqegDxQVARg+
IpuWMAVg/HSKQlWCuiDyClrqayMFfr32Q/R0wpik43OJJaqCCf9e0nSYUrqjOsuU
9G+QATQYXkICwA95sQ2Wsse/TXVwuF5XVBncpeFA5OQ1POl/c8FtHcXqu+Vystea
xVnDKJwFf2J0m7CWY3rJQztDyjadrPX6VThisycPgFJcDb1DiYCtf+i7l4G3LjTy
4c10CFR6ofLeUejugNr1P0JOcoFsdQTaxT6o99hInlx3K2NKZAd1dv49A2YBRGbd
E2yLNq3rKBS1yrZuVvslRsdj4EbApu8eXpRcV20sAA77sgm8HedMVxLQLUBtQX4v
Ipkt7m1IKFDWe6tEEnVhkY+c8jNhMF0sXnXFCAAU+7cUhvrhxl4zwl2aHsGGaKDx
z+dUzfEZWB+CYQb+GJPQHB6ED4YoqjGTFlFN8LWYiplVRHsLHOW1hBhv9mZjpvL1
rrT2wWMJtJNIDs68OHc5T+6MxtwYfCt/gpA/pC9lnVqUx+ani20mei8SJvDePin/
hwm2I7V/jXxTrb30/kDcxtl3w6AvcUlIGAYV1uGYJ9tBEeihZtJoqrIPfuPLiOju
BolM/0uHPiFkIXnoDNk4uV0cumaA7/9XRKh4OPg9ZcEwrwZDIHSsWFt3QBjY0oFe
XdtWfH2o8IC4x7V103iZQZ/3ezN82Vkrm1xxoOjlxSMyYqLCJnItOv1xzghhU7EO
Rb8aJveNj0ujzHRS6w2b231a0hCtJDUF7MA6bTdRTbVSKo8nvIl2BKBbZw0YCndx
90lKKAlerS6sAQiwSOp+CV4IIasGatDDIifVA8WmGBRcOtaQuJJqEtK5htedn+Qr
iUHOrMMVvWxCNIBaa5np5lkQiT8ZOT3ZvNR0Qnh7QswkQ0nf3HLlY5SUiQ8QOfgb
doF1hFnbsGuEgCKzbJzzNNeetUFdH6/j25GYE8bNZ92asFnvssNXtqxYxxccb2Eh
BD+VGk8TYSNapv5/6Yx3woL0gC2j8/6zcrQ3iZBPz58u09Nd+Vs914CsQXyPXH/B
+FgiHxkMw5ltc5mvfgGMSkeARGQGTEVaROmqiPasURdEtj4klujOhkfjdCB2gdBh
4G7F3XbfDflsaKj1dVNX01zDwmT1Q7BZk0aGt4ZzEa8BdRdbc7fZ9WBXo+ukMCOq
IYtxwu912UbKNZj+TXbMYl2nNdzsXwQT9UFKzi494FfEz+CfvuwbZxBdBC/oHAiM
jvY/4mF8r9ZwYQRcJ02mDU1GqmolcSlrXk8ebD0fputfp4/GnF3+mRjBgEGfJWX2
yRAgtEwiS6qGv0/0/v9cvjn8APPlUuJFeOKdP1YpCHFGd3Ex18v/qa3CjhQubgKs
mooqZQxvIK9ZA097MfHbwG4FgQMJWX8cT7QSFNntXBw5INDGNCp8aiCZmV68zeZL
8bYEeLT+v4/lZj007FakOe/K9Ua4azJIog7XEbaBRB31lCYlgTAWzDxEIQ044hf7
5NlqebHi+mwFBtYUUDIM9ghNhyZlrYYCErVe9nEjIKvGv4ZOfmywOnoJrPryWsnF
3QeB1U5reCxudbJlrhoGjSllRBRpBc6MUcSYOugImsl5uGkTYeJ3sv5w5nZgwl5Y
mSpTHx4zZlXrJqS9pc7yNPFplNI6QNxG3nSkR0+DOpKdo6Q/ym0umfPZt/c0gub7
/HfXaY36xx0cGXsfiN30QlRFH4lFNsEXCVHoKPs4EHp+MAWOxv/Ta7eQtv8MdCuG
lfm1AUlOJli/LsBJvsht9ZqRvCI4Hl/W19B/n3p/5ztphckiKrM/3mgjKcLgd2xX
ThjUJv2PV7XE2LKrAyIZAdlqhTeub4adkBSgiTR5MCO7mQcewTYQL3hXPHqUdBA5
KgRcj11maa1IS7rQiGofQpr7/s3kZsDD3RD1cb7Enx6N7mxuCiURFkPriIlRqKhZ
L4jtUpPd5i80lWnnd7kafq5UFi5IS3pUg7Z2WVeUyVQMQ5rGrSsZm8UE2efen+W4
rV5OPcFs90DEhaIBLYay63iCc9l9hS2rw0nXoR6ybjHIVPx04cxWjdfW++BeE9P+
zGDu6z/hVtEad25c/Cpp0GpgljJS6N3SXjwxbBHUWGBlp0+q8wfIlcTMNTItJ0ue
TJaa+lBMvRfMgI4IMiGWZv8a+lURp69Ku3gyoiJ4GO7R5THrbZa7nfPmjas2bcpK
WLpSKPV3uLICwSK45lwOYz1OOxjlSMozfpQ+SqlqFY0yPNXDI/0evwMRXZgFeXQ/
rCgOgvLRHv/lMk1W5/dsmzw9j0isAi/aw9SGTzvzBhCNTextdjjC3OYvQuap2dvH
ZLfYeeIFle/ogGz7WOPZlWcQaRhgdSnC/s5UV07MpannhWOuhsQl83t9QMW1/7gu
uTrABtdrUvuCvNDZFxU/ioauckOblC6cmo6ARgTAxrCCBji72dfRCakoDCok01GS
97oeTJshUC68cEiWGYAsGoW/V94c2SjqNOxxj4CStdcXQKFLCs0hNNYGe6etS9/Y
Q5T4IGWjX8dmRPrjUYwwUzhD/q6KJ8JNCLvbTS+DwsSikOopeQbXC6uSAuh0D+nA
2xm086qw+DUuneJqwWzXxLTMoP8nFFmiSfJqrP3ciETA6Jr/oDLMk1obv5UVr0am
VoA89LrPkuPOZZN6vow2XH8pKip/xIrk4V8HxV8dopoQVe38PgHyHtJYpTio8Slh
6WVRgeLj7CJxzLKlAimx7ZFdwahBxJhRqb2hLRYHN/nyfYH+V+sQOEuPmn0cnxAt
jDIkgvYvG7iHQ3KuV1e4mpQmAjBsPG0HmqpFdv+uvtVLi1GLD2VKP9hH7C6kFmoS
1qMW/bpTOp6SbNAcPz2LqLHr3goQwGTNiUayEUx3PzYuswg8R/6YuhA6qeuA5RC6
edjeTruvItpl5Ry7y3gB8Xfk2pYGBaqCX+mkyNgVjbQo/x+C6jyTTmzqJO3XGkdF
oWVgDKGGNKZF7UKau/6EOhOWjGPforve70EYUfVUFEcpvKXccnByrUG2JgFyOjIr
FbCmlePoVouhmbIRxpm5OsC6RJjM8fHO7zs3XSBljNUdufRJjNDnarOp37msoqfF
3pFwTUXBxGQ/3osF2ZjtXsPHByYkflO2WLiuLMTa4Si/kBdAEGhOuaAT8b/bsJdW
S5Twp4w+Jf41nNfTvexSqYmheWwc6jzWqUxGm6vL6+Qn8wu5aREzcuiwNMOFQhDW
kX3S3KtyPoU5i4ukVwTx4nvJ9VAjwfkCICT4EehjvElVxa8imiyU4Ez5+nFfafC5
soSyeSlMYvWpyMMf8p6Tu9iSwEpdDAmWz3sRTfcCsdG5l0y6JnL08NZuwYV0pI+g
glYRlGfRxh9ut+cQHRZB5lxeY6OBdpLMWxb5zrEY09ysHSa9HFSEUis4/GKHi+/W
QrRDD1GfzzWx79hZzz1lt0mqw/XnFZ5qVm28U+1EPTcxqtP5qJiMnG6LYQoh//d+
VTBkmd2RJeiNbwnVdmPAaHhVpzCV8CACldCaf8uGxYrwiritki6NyvTb8LS+02iZ
gjP0Aaks7OJXWMOjbvm7ulI3n/aaV18+v+40uPK7ju15WePSvzujtjC2W2d9eMwS
A5V0hxATl4A9wQjx8g7eEIUAPBzr9NF9j7E/N6eV66cRsqYVWUoNvxyNsDfy70RO
oWa/WoS5bA1Tka2OE4X/cblNMgUjuBG2zd+G7nFc84u9V1935juwU5fYmkbtr5J/
BHfCvyuPqjpIaVpaTTIGpAjoeaz6JsWTt6zVjgGTOyp8jHuDS1BnIarksOHFrcAd
iLrR7o1WllP0gWsW708AP7Nyz0h7zkoxOvPmMNprI6MlTJYkk9oNtX2PvfcPqavf
RDfGT5KRuZr/B5KVQysLnf351Mk0cGV7fc68NbRDuT+KNHbtLBbKVZQmpTOHZLpT
YZJN+bwO/HaFCgB+2RGirfmOAMdL03EH+SLTpX9ZCDDUdCJBBwEI3SW/7ZrknH4c
W0Cxtm6t1O8bjm+g9jqhAmZmxSlCGYWJ221O+AvICHX3rnr+UlbIghy4XTagiqo3
x5p6mVHeQNvtX1qRnHLgoroBdRInm3uSi3TU+SPq1WFunlhB6pwZ3FegxJS/9QTC
40BVyliTNCOVqjliiMvBHcQNwOJ2/NARp5V+SefnDlxj0mbtVYFIppkcrRy0Cgej
1g5lg2uDSCsIorx3ngDJ6Ny4qDn9EaWBsxCIyTRGi7ULdIsNeUuHTWovcxDYB7eI
lewXg0ZNb8nDLFZ68vTXXNCzK4wMm2sWAwWBFUEPh77pY+o57/ZdBGkk74DfF+FK
x59eUPYu8fDvZrf05dg4vUR40368TMLHKaC+jdrtHF+WsPcp7yaOqjVyFXwIeb7j
SJ1qDg7mjX9h8yjTZbDJn7Vonfk5/GBlSs5iF5hiAS105RNse3Ai7zzo3JnDw5gB
cihqO7zxzuSDOAA4AmjqaYJNwWZkvEWzw17X/7gCqhUqAabphWGdZn91Wglm3A+p
IKlQMzoYci77DWt7e2JbpN6lmEa0fWLl4NkfVNalPDcudCHaB3F/CIdYGgRe5gYq
JTq9XEpjU0ssLyRHw08xFJg+IAzbQDG6LMWnRRByjvm/47eEPsYGEZYx3ZoDPqze
pAPZMFvckiiaoSqbZS2Yllx1edCcSYFmFbRPZDKm0EdfhhInvsfdzW2WyuUpprJE
RyLoQX/kINKBtHjKdnyrYZJK4tzmqGN1C/wvF2HZTnLOES1BAOF7tORLN4G1GJuC
2pAcoL+ujW6Mhy+LRB9iO/rVpw8stg8g+UCam0p2MLCnQo7wMZqNSN2KwgDMHnn6
f4E/2Awj/d05KY/PmeZdCXAVjK/yNdTwwew7PnJPDMqm7FWDAN3jTFumMTofv/pF
YPno2ii7S7lO7k5fdoEaP76V6stfpnCWKCS0OJu3IFAS10rqP3P88rBK3fzCrt8y
kQPy/wHBosXgPySCpmRhpqlymOdGL8EGsUi2tE34OQ5A2tvYlC5j4AjsV+8Kw8ug
ZW4o93QXL/8pfdaU16BDbarve4my08sSep5afJTM7sFipfmsFjUubT+kr2A/r891
cvdz2qlGglq0EGuBeqF6J26bnD+mVRj+ZwH1Mj/9XW0sedtizCL+oS72GmRyTVb9
SeK6LodwEkPRGgU7Z7T2rQ13ZOmVS6tSjO7csMoAisw08L2B6UoB+aBXJ1LikgIb
zgVPpgmXWn7p4FapEp3JPVaZwb1WtiJ9FXE4eIvlT7tczZPLTipb/f+v51ZHa6i2
edCZZWVc2kNfZVfir0CohHpgDUw8g9odhZy8zhnO6G0NUuC0/y21hB7T9uoEl791
PgUA5hEGwjV+z2LjOh3pAoRDCsoSr7ZosYo1WCAJoi/z6ZpoT00uNBYAWoWmopZr
Y3uSLsZCL0C72LfBWNmiCk67id9FHp1yTfTWNkA8GSNp452wHf63mO4L5H7jg+2l
d4UbN5cfB/5go5FoblC4AyKArqnXzb8S+qcBWig681G1LaGATVCWKsm1gBJnKgEP
m3WKpPq5Iwb/4qjKgzjgk9uU3YyPV+WpuaaztZKSt2aw1b9hvbJiTSZbaQu30Yyg
9zesoDsZWWpYPEpxnD1SVJozHaDTPxv1yf4xL5yGJPg96oa6O3M2oRJb8ZElFCf2
TDMc2e8niSLuEYV3rhJf6kq9nUYicbCfethAuoo7yTPYSHiQs/xwuvk7V2MjuqJz
d2rstUh15fmAaRoMFpA/BDvJfi0YCFtT8FqJ8bJDk1DoDjNahMl1bR50VzNDSHkx
3562Q/XMOZbJnsTqqmRGBMhr0HLtV84L+oS1RiymD1Pc/gTLh0dZKZsC/2scRVeL
eIyjG6LRGQ/XUN0OCqJ8TfE0UPqcKT0OyC4hQHpBZM2yBe5VN4uxlQI9ahHzQKpp
Unbgk2J7uiEYF8JTtrLUYTRGL3HpMOTlAE6qY4y53k4HEHO3uw6DlcEVXVqULsTn
9YvUgjhm+Knf4JPsr9VeSDBn8REX+xlvO+HsHRnH567BcWFmYDqOl95h1+942wO5
/CwYvhsNT5wi28x3mCkdiVpEpO9zsvnkyFdEHLvDVafcOStBfi2oFWVqzPsbM4JC
G0E6eIqgTohGXPBqXMBK5KDtRzlARWVSfqij6b5jQ9PBKHTcyh74o8As+7jrla90
CuDKdraU4BXoPKanmxEWWUlaPaWjVd0Nyxha2UDsXCHnY36SL/lNXyTcROCgBHAf
qN/VZls9apshrrc5cXBzsKZ4JFesw9uruIFLZ/OSmFaakNqX2STLqrHewSj9IoA/
xl0CJ78cxDSzFgw7MxBYAZTjU39hS8mPgNks+RthbUhva2molqkFdnXMKjlS8zAO
bnOowvY1NM4LF9h5qjsly75YHWzXou7GwJRi2tIKsSPOmxpqA/ydudKHZab8wxxl
ZN0paac6aaLRahGUA7zoqiizVkZMCEqGSFxCrbp5mP/p19iGbVSvACCBry4kHpY4
LJkqzR2wtOFbIidTgZJVJrEiBRoj1HN40WqyAdbW62Zc8QFHDpwvjdMjJOfd3JUz
xW73yA0GaX2iELAd2TTxxOTnIKNTK9AAMI9r0rSHJuklPzg5yzgzVbp0ZYm/DS+c
Nf9wncKh2u5K+0dbIAWOtckGa0JGhCl+AXJlv5vE7CmUoS9/L59HXJk+Bj4oP0Kp
7pPAgwAK2Gv/MCya63ytq2MkigpgB/sDT0+QIxJbBTH04yIjIKMeyTQtS+a9d1O8
zWdS44YGVuL5t13qqAfAuFN5rpPdo7aPRHde2wuU/YbMsy6wJvu5dpCHK/J038aw
r+6xt6q7AfgoggY9iJVEPK6VnYAOaPwoKyJOVl4agnuAY8ODIlTmTl0i1Mfq8+u9
+E9wl5Erj0h2zzAqdC/+rjnbzhb6mw64xy9goDuyhVR8lyZFdxN18zWK+7YOOOB5
XjySCdrYto8mY/yg9mwAEERv+TWmPFAUXPXxyIu+9uyMpL+gBPvj4OqdUX0RvjmR
M7mgdVt9tWlRxSVG67Ez2h8rwFwP2Ozpxq5p0JrGlMw5EkymZx6lgKv1+veLrLV7
SUDkmrlXlGcb+dFA/ouJyiNE5UrWfrS96YOLYb8xYp9qm3MvQDhH5qCu6kXxslF+
0s+MiHXElzigh1BoYWK8K2PVJBw/WvRUsSyk3/16aK1TERF6xFCcRUqbeRT7IGeo
GfCPPvljyxUOWXKqvL6R35S851x+2Y63aUl2leT8qaVm8pRAIwcrSHX+cKcmPlzd
3eNAzjeuxbOI6yW1hu0Qy7hObXVQSimCPyHAxDAPrJbpSnfs/53Qm0Do5Z3q1pZ7
PYv/qpy5Y3PXfPWiFRXGfkfvo76MUPrNDfw8ybPb7/zDplfth/KYNCqRSD66T8FH
BnT8Ay3/10BhP7kHzBKwVa3HUB72Mz9DV3gcaqKMjJ+uW96Glc4A0MaaFFr9QXFZ
LC4YKqaXM0iHI2g/6+ABTFTGh+paVhJoZggcu7Kwggin02EBvxRAHmP9arU8X4XC
EedI9xbNU/oQTpXSawDs53fsm91S2GfEKB+rVFheS0cM7j8TZkrXBMMuF7tWjxlu
keWLZQhpmpiYVqUGLgdM61SirbF18uwiWnzMGCBlGX7dR/fQdglRGUOiojCf2LHL
Lr3NeONfqIQ+nIzNfJF318ZlhNJLWpAajiU/IC/+ckRhWBc9fA8+GCWlxfBgZakc
PjiNjsSHsjrxh8XQlrFMb5TbxFRG19BrNTnEx+kVQ1oWW6ykmLJLA8OR/yC9EPWo
dCLTbwagehhKXJzfLXyNYRG7yYfA6BU/e+UnxWJ18/3UtzW4+LuXmKRHtVOBhEdy
/8Fj/oWnSI50ZertfLKbHyUuhSZ7SZWrHjepyjy58p7x4OiSwTDOb1ul+ttshbx+
41+epUUx6Kro1qb1soKBlWQSqAmv7E+1PUDRsV/9/0175MkwU4UxI0xeOGfSAZaG
SqFJTOVKytDNJ+xU3kIGWeNy9uJTpv9sy4DghPOxSfy1NiS9xDS9brzw5ATFozoA
fThfjJnJe/ScwJ+74pOJsKq48lrhZkU7R0Lj01vzG8bz88wLtf64loTTJGzfsr6Y
YbXKe4GFKdPwCr6Z99X7iJ51Iih0lxXyE0Z7qUSTl1u5SY3t8+lata2XlrcI385J
cMjyPmyniTwmZGgNCyJB4lZ4m167Nl8EtMO6jjcoWJwBy7hOccWNXq3aFwLAJUgn
sz8MLXmze0gpaPDepC08UTI1LI5u9OWrRwSIFvj5+tINj5SEcy8aOnJyduRPsMyt
0GYWNRjgru+855e093ap1Oq3mcPqR41LATrgq0uMjX/r8dxnTSBer4YLTatthDxB
i/JYQwDj4oI17UaW1Ts6OHAfjkESrj5Qswzw5f4lJOaUAF8nfuIqRo7P4g3sJ5/o
ppkNXIHUqQ5Vxfeqm6gpu29wpXC1pp68WzK5KOOEzE9inhUSZg8k7BLLM8M3X6Pq
kCDrKUcYbRf26rF0dtYdwxwyPeFUFdH12X1oCskJPZLCgCY+imoNp/TavhVwCbDh
0VS/VVb3ze/t/wy3vasSBg==
`pragma protect end_protected
