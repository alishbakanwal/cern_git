// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:42 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QUBDExyjkjNJUm6oGrY5BOpIL4gxBr7v4mpD2VoFR5zlvPOaHYr2kv5TiUz/Bnbt
c8jaL8hh3UEAq694extQD56V6HwF0GC2NUWDJ6YgS5lxocKi41fvktiVxb9I6VKZ
Ad69BWoUHFcPVe4J24Yy1hzdkgf7jgcDShZlqWv/7sM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20992)
tZGP4g3nuPaclemqf0dMPt8pea1EITg2O9hL3cU1U2YWYfn6L4/nDIz8oJUdQ6WS
uINie0f7Humo2L2KQJkItjg04dzerVltL7MTIzGCt4F/ecMwKqit4Hb11XC9sbz6
8PdvTgDyiQRTlprRiDVAChjqlNcF/E12OpH8s2TE5ZLc0Lfq7JszaIWFNng07to6
sG75jX4ZYh9t7yY6wGKOCq70CjlMwA3PZl7hY4b1M0wIcO4+K5gNXROBcB7iES+F
N0y0BK8WSadMj9f8BxEbhBr5xLTuoLa7iBdkSfu0b3ddRB3QnASochCWeT+Oz8rp
CqorDBpVIvEsVqRKMyBFjwSzFg7ShAf2taflupr8Y+zTY6wa1fjMpz4o5MVzz6Ym
hPBlF65p4oN59d6FcX4K6adtaYf+W321SjTpfjN8b6Jm2HwSYet/eUecsa98icbo
yGoPBEIZ4aXtu/ii5FKq/UzNvDzBuztKVv3bJZS/FN/Smliw966EC+vh3H54MIn2
GlFoIR7x81ehFxLrJujoKxNAoGAvDI5LdAxixxQ9UjxKuSNiLHbC0f8+G3Y8AJVS
5L+vi5GaL/YDGLnrMKV6iPUAnb5bFikUZ6AzHerEv19L8zC7bWYU1rqBxe9rBUzr
JsTRvMIxzPu09wwh6z/SlVoNeDEvUba8gbYMj5FKo6kktco33rtPIcdQ7LZaEagX
Zo0JH4GqktQ6i3AJcWHL4M8H8/p2PjxNfpAXkwTNxCcJMYt0kYFj/hxPJsvKM0R1
5373QJ0OWxDNPaBwxGIVb4D/078BRNfbRXD2hhV/OKEKAfSPS7Zv6z2SFoYr6O4P
MgllooEiVKHK9IuQE4QJGGZykHWdoNzOMZ1slp5juBOhsgr+mY6/9IYWbPe4Hvmm
A2dKF00bthrFdDDT+Hx9Wbea/JSABJy1x7b89tDgJ8j2fAmJFprujtCzJUfij5fz
Pq8uiKRWbFvo4qxQIGMZ3VubQ2jVRMntk6/IvBOXtX/OHuZSpo05i0xMcBKp1fVV
BHd3I/TPBVGWVYBTDqMLULv7Z+MgNzpAIwBHWK8F4TrRgwV92pHU1cxEXrJlcxjG
el7VaxN1ipEZAdfrFH2eRyBmS75UX9S8hi+eQfzXzksNT4sgPG72l59aO9c4CfbM
PSmL3NbG6yu+M86AkcHT+fA95CjE+P7v4z7G7RZV9dLSf/dEtd92I6ywZbaDzNtB
ZUHMXauDgLCCf+n84A3J7FMBrG0ANjQdfklUCqHKioPCjbL5MOY42bXVJEr9urHx
BRyVlOAw/kLPI287sBPPGgVFolFOHrhnVDdJXCkPuRXR7BGriIZbi0ZRc9v9aXMO
fCz0EpfyjlZ37GpmjLhwNbRfUOiZ3vt/fH/Hju5m7cSOZzOp1goQKHj9QhyYINuT
T3Hc2sc+H/T5QNnsR4LovvGAdp1sPGYN6/tclDvDOFFYY0lhHOQLzUPyFw8mtiw9
W7JimOM8ie/qowSfhLtP5fj9O1XFnM7trseL6plQre4pY60qOI+F6vaDZbRT3PiV
yqjfzIUNIkUM4X2ik0pePMLNNWntl76YnoQpSiqtFoEF4Nz354tCMFLck2qs8M/k
nuoEKNmVmd7HtGlBc9dR78+CPmloGdGLlI7hj0ig+Do7MaNbJKEsRiKmYMBTVCtM
BBneUrvvo7LMHk67XrbdT8IzBlw5HmftLaWCzJCrY6kGKiMNKk3Sb+BLphXeBD6j
cv696Y9IrlZQj/Fqg/15y8MxVuJNpKBL+vDvDdoXVK3QOIjzaULSCftUxKxfn2n3
n9IQeuFXwer59gqi/fxj7gVf0ccOZ0w4g9BjfuwKwHbgt8J7Ra7ytZl7I6fwhx76
vM2XT8xgl8FpfB+M5XXi2gTChVaWfQvCV/nM4SC6DPajXlK97BsHJWkVk0bHnYT+
gZSD7sRlz5Q4QZtv2rkuAuYoLGTO+vXeXqr6sGQ7FsDrQ0ybavTAz9diYFgWEy78
UgifbVqyO8h6YUw2sFlee6WyasGQ4q8ox3ymInRerx9CvcmXiPcgIDaSoXnSNusw
2VxnBfEwc81R+mnD2rdx4/bpjQQyaYyFUWYjz2lk9VyIeI6FkI4qJSURsp9czVzk
bYw/r7Fh8GC76tGRkG4BD9++NahtrHrgYc7I94o3oj/LZ0k15hh2hp5wWz+qT9NL
NRBjlvL51BXqfmcZqouJnP7Zel31RKh9AVuPB0fCnHz/fgjlDxWUz4OEDGY1y42G
XDEkp1mt1aQGO43dJwuSUGEYB38IZIaMVT3SdprfI37ejOr8lkw1HbiZJWzBWtiE
Ypf+B0f7pbVxsUVxNj/LjaWp5WykF3+ZN9+1jm8yaEWAcr9n/wKWMtwYwaBODoD7
t2Hik7ouSNwTv0QTSah3Doi9vV+Jg/y6non3VyjFAQYwmdwhKMygcwVLG/DILKZF
XuoJ143JxTfxCWEWRJRjfKGt98YRVLZaKO+vR7yxRsmOB9eeiHoWGrYVuAnJXyFe
FHneTDnqaxm9+RdG9E7HlFEwX97cCImgKBxbgN9Ppoh1w4qTFLWYr9Iud39WUuVQ
nOnm4mW7iYTkMt2Q1JP3NVPk2Kcn4MoOtsTaUzLjJN/syq4BsalRXtukrPI7bd44
tYLpXQWkxbX8c4MSQtza2K04oOOyxC2gF+P2zelbcL5+VLSITI8KrfR968vNA3bg
OLGjLp4W8JDfyPbSs/b4mlbVPQ4KzTgyZOnLAcAYObY7Cenpn7AXBIQiAUGF4jdf
7eUAx+x++Xx5wbdmpzLeJrHFyU2laZCnlcIrppbVZJli3DVufym8d2PpuCr2j3RJ
hq8Nozt7LQW0WAZXs+sFzl91MEP9UlS//9yxNahLi2eInqAf1FsiLTn+rKxCb6Jy
ZVUlmiCD5r5dvAEJncM06PpvZw8q3KN3ZleF0FTKucb62C3THD95rm4NL10ny13Y
IsIn4slQBKsOeG9Zt6DTvF95y7EV3hwaU9iM2lxtHqOz0kz4QrdEGMbNUrZdB/rT
HrXj9LRbyJnAvN7hIj/L5zHhTSK5aiBY/zjpc/9NgGxcT/TltB6cIhdtPTYiZF2o
xO4pQ/wh/8XWv/CxNfYvlvGUXG4ttL2YuDAaEJsNrB345V8UZnYSv9kdGS/JjTtz
Re9oGWfkB39xKQ5T32h7W9rF2IXGWAUfMB9yKMGBaP/XKrRoG/04pte9AEKR02DN
tB7ksokzxXPZkzk6wXkCOwSVoNJkLPBzac5p3RWkQTJsylaCgzGZP0qg45+VEp8O
sDQT4awTep2lqPI/Bs1cDINtdMStvBIjOz0mZDNJy37Cb1PYO7VOaGMX+NHAqBgR
oKBaVODHz/Sxi19YawkA68nf8Zwki07lsrE6inNP4rNMPhKuX/aL0Yc8VsKmchyS
gvVkNskRwDQDbeqmI3xIo7pjAcniPOFhnJTMbDcSwfm8o6/9qgc0/BodgRWESRsu
c0fm3kA2y/QZ/e7aNl34z9Z4oettZrPm3H7Xf/ICWArvaeS2Vp/wYy/ZUx2E3KPC
//1+qOxq4O83kGdWyPae7mUxUXAYuyI/HDCIQvhB+zEGVhgNEut9SGjDDQ882ecn
gPmZkMcCKUC+5+jbn52RtpN1t1RxBOOh/eN8JzHHzSZtF3msQhE5uwA2qhLYfqod
s4rZgcKbEkBpu4V3yVN4u6KZDVe0BL8mEKRhC8S6oKKVHI1Rsa1N4IFPXFBlS9hH
tcLsY9n2uD1fh/GrOYxVFE3icHfrOEtQLW8NlgsAIDOS+hD5LlF0mFA4MwWmzX0I
dj6zNgYRxV62Z/1BYwP7Ea9TXrHECmrQHoMEVm4ZT3v86Q0ZksCaQ5oH3u5xFa7r
OF54rg80+E3w1mnBEGJgoAZqIvInR2Evo45fWqDi9r3xbIQi1eGBonoM0VtXOOgp
1m2tH/DKL0h0aCRxmt8IkqH0bKagbhHStg3YjiXrVoo3lEs4qIFSiI8caqRjTotw
PJ30ETDqXNPowVf6C+MVVNpnynocWAuKuD82sLWOdYz0zn9pzQ09hCqAcFApy7YF
3VqoH9sJ5/HqDVY7n9bvKGfcvfO9/6lXR66i0eP/pzy2Tikcst3yD4s5AnLFV1D4
NhJrBGd3dDQEdBMPDaMFO7coKXzLPDMaFe/cHGTKk6gJpgPuAQVUSHPuwGwOHiWw
sdKV/phHchdh0h3IDYHTXROa8rsxdAdlR/4WBSxZojWn8J55NOBbjk5g5QNd4p5A
IKkzJ1F7hEtX104r6KW3FQdrpQUuv2MsscmzWNWYq9PHknwBw+e7RKo/L+rncfmx
55rS1MfHhe4QNGeJU4I2ibgsSWa5OZH0GaUFfETRbYTayzm2xAUB4h5AElzRAfs4
cjU6w6YZI5TG4xkDJyXZ3QuwOu9KFvQZ2uGCvkBk+DtfGLWbObDjo7ynclQEL8FL
dTgeHhMrAJcH8nA7dfqOWJHx8buWXdLmsL2rHFrC04ParZHmUGrmuBQt0BWzMhIU
blTwURCtj5+ZcCoSLoBF3TI8px9w0PxU542Ee8tbToiGk9N65M7RkfmjXe6cp9GS
n38goplcUenLiMs6jN2WoBxk2HoD91g2hxf9jDr/MlO7/2QK7uy6n6P/If4ooyhf
dXrhv7MDvcSeUOtnIM9JfSITXWBLwQ8ZYXQLcuE/9EydS4+ktGJzqgzpkTKKYfZR
/D4R73/PYwoJH7vichJlKfRjxYHv3t6KpQC1i9YeeWqe6gd7q6ZG+4yqr1j8SRrF
84PQf2nTRJLFOTM90eg7sdUayOketTI1yaVfv3F9UROETAWAPZCcjQ6o+sfZE+xb
vsKcgxOWPeiQ8Z70I2m9MJdVIZ8tYcfwQj0qfG++MxBmCqvYy4OtIjuiHx98MsAY
pizfRK9Ogto1rt3coNgP7WmijIxi21jfo0+w4eP0Wb8vRwz7TOc8z3l7iR/AhqcB
ucJeR5xzP84JzTb9fYL5oFO3NQ+1vL7jGIjXlJiLtqG3UmXRjvyszN5+U6clW/BM
xdbFwZ4tGAT3c4qs/iGsREG+LXFZo+XcguzpJkYbeuDKxQ8dCc3Baa+XaFNLDgTZ
EFLunj0gc4KA95xKu0C/ZxqzKC4bn9Y5ZfaJMKJpbUrNUtYjSuoYBCeTz62DxXd/
zIzmmjxPCYkwi8eaquGBBuAoy3u1H5GfbpqJD5UjcmPN92fhOn6uIKTgvk8UoE1w
9fM3owD3Oea1lwVDKmisb8HblxjNpjUawrkv9/TatF47LQqj/Do6VbtjW1k1OFsq
Ud+kxRHCLGkpch23xFPCjRfKUfO7o07+xnnJpQ0dLMId3K04DqYew00qbWQOvZaE
s/WpeUppBTLgi/5DLzqE/dd3kuvdOVc+oVH4Wbx1edFQ/iXkVMCe6TfabHFo5nmd
DqDYN//9PY0l50fCpP8wHuW+Kg7yt5lNv1LWJLnmd6AYITZnYzzDjC6BRQ/WdJaS
eXsNPVmVfn7hjb3sIxWEWxmzPnJ9bpLGQ4y8RtMw8ATmI0Z8MbF/Cx+biBpGtQLt
a+yPqUKMwBEr5+N4KJz3HkiUWRkJj4t37QBGJjGcJLkjokzydwPU8kagiDesk+IX
GPzpNM8VfbfAe5nQyOTreL9ofRb0K/xU2sCxM+revHXShQlHkutxlETjFwq0uZ5p
4e5CWE+gvBqYTCE/0CxoiOD01o9F2L0ZmvQUCO8NI/VlkWpjsvdiaIPRrt5uoICn
BvTp4mlORD36uvFzQpQkBYSIdQDWbweMWDuJpKU0HfXMitVfe6e0UVykMGCrxGWz
HTsbL94wOEzn9/9/I/dfPkxciTCKCi0oOLDc/9g15OK98Ccf5TlTgbWSlKWx7SD5
q9x2inAEvpPc+jaGcgTDtRA+VgJ3/BNOm8YRq6ut4piOQzUSSeAPLmSy6O4PCCm2
60TcUqRnDcAk7R1L/lzUmdD5qJ7F7ieJXp4qnWhshTL1dq7vD9ajf1CXVq42sfL2
UthtDfsHtMI38wia3I2s6qmIUeMOh8wkLvoA2wfxd9Zy8RlCA5YQsW8+mp+3j0ox
ulz6UD7yk7bjpzIi3a0UwCWgF9X0s3J/UHyvyCIeoZb68XKgxx+IZB9CC+VmQA/2
T9KtReLWNaFOPTqQQGaAWRWUfsX+v93sJZ7VACeP0jzQlAOKTvPNyrvP2l9OoOh8
bH3lnu80EiZBfy9jgMDCkP9Ey+ds8wcyrqvtGGhuoLLFlqC14u6niCM5jrarGcpL
fi4gcXQfKtOlDsPWPaMJtxuQIU1x8ef3VcL4QUzlXcQqq0jqw+cnBU7lMzP6xoTe
4Snbgh/yvneP9a5SegI+dCYWt3ZikOTQJOO146/z2tR04DjMl7KAybppA8npJDHv
uUF+vs9d3zT4dcK/gUoaoIWmcrU0Kb8F/ILYfW3v2lNAMA7MQCHHHrWnD099NXrR
Gdf5RjUy3Xm6aUe0JtfRQHYlQhCe2lIRGoCUdGIEFkJdzwcWONJ73MsalLooUN6/
PMxSz+4wPqoVfmd4npFXN9q4XGsO8geRgiyOoWGqAj1f97ky0kjYkpIL3RHf0Q2n
nmqXqDBP24KBbzlRKBMIPWWCIbvTZwhl6F/AwqHouYGigYKDBwgjCwT06otNYBfm
ufFGxbKALrqd6ml8s9irQLcc3y/9/XckIef+xcc1qxCqZkKgBEAaF3aM6HacRCdq
p7BLdLeYImgflqbFY7otNw9vvxJ+LufI7YHnUwoR2zs8xCFQZqjzrlHc9HjlGay9
E6hk8cZLMk5vZmZ3WZuXZtr6XUBnTUZ+wCxqdtIWehNVEG0zODsuW+1EDGR8Sajs
aShMLakgBviC+CZ7g1gcjDwaSCrybxAQAGSkq3gs16xmzz6fJxgB7TKdjqwEEE61
npD8JEih4psNbq65KbYu1zTHAnbLmQq92ZEMhKJWrfVonF8d8zn9znWdPveBm9Er
J1xw1OZY84lYGOt1VXlN0X9zkrf1eTtoVlrOHKCqncFQF17ga6IQfqvyrXf3A/3A
ndfEUJ45g7ZVIUxK/acYwRSUiXARZbtJecDvjQAsu6WifFDTz5bbvvPkMUJQe0oc
kn41uhlkrc6/bPZ5/vlRfznHC3h38yNUZN+eEujpNQyVa4Yq7frs9AFzYvXByQ56
grFEXgl+hARSTxZuzq8SIxlc7dZ6Qak0VAswmmclN1ZLY3KXoIeHehMxdzlzxbNi
Z47WwZihf8Fjafg56VpXPMKZQgAMlilIzOOi4fERe5OiM6vFVozONAwt+WI7s4mF
XTOj8zyt2oONolyozoqM+bGRnNt843ZVYObgF3oXXj5u1FXnvH2V3orb0dwcUsdA
z2soOgcbA7UJNQGMQWfZCtwDP/FSTIUbMcZbY8KMtTOG8YcIdvsz6ziSfkTEvJ6p
n2z2DK3zWSpw38FvpjeoVskzYE5aBUMWvZVY9s17d4KcxK41j8tGQ5gm2THB6zrQ
ciwLAi1alMqNo7cxolnQoM9p5uc8dNh9p+aUMAJ5KcRgLe1sF6J7VP5s8dUO577Z
JTc3ie5+IP+tGNHGzmdfVLkMrFaiZP+09B0NQkqaRDe0UU3Odj7TbeAkaSmoo6UM
rBqFL9V1ZqdbKWiYV52YnHeb8ezSocGw9bSKcWHcTBCwM5Zlc4Vh+S19z/KAlY4+
qstxQNHxJe5vxPP/zCYh6lBIlpAH3CN5PdNeiyf2VPb3kdcy2MYiOrtkhrASnyqo
r4UMkYIEx0H4xVRPnF5zpBsAZNk95O4yj+WUKofRjFihJ5MMyKWXQ6DWWbAUHSUM
UPsYYLf6mLmUJNc+++ArfEM1pfRMfpJPwyq2kjpehlunkbDbRTd/vZt/8OvxhJrR
upZRktUnRIj7PjUgz+7SmYmqiZJGqSX4aNKxb7eNpGvjelNuuyIywUeHB0exazD8
IiiOHI2jhsr2i8+IHJV0pDONyG3+2EKh5fSJnjWQVaHX99OKZ7qw+cbGdOXppx7D
0O8fWqE51G6Fa+gpov2yfIFaZnosKCHTWokA9iclAyy+/Ijpk7+tkYerP6SJShpb
ws2NUkQv1dch4aZh9JpUf2Llz75AiErvP+bhQGAZSlKJ/OinOFlOtDAFH7tGPfQr
UllWaVg4UGYrD+dIywj7OeGiHpaVX7bBBhSdHTLY/a7tsB8iE/Dk96UAwUUNF0sl
IOAC4wobfqzZt8N6Q2VelftWSCytrfEAuwPJR/JByRRru7amITMx+DsDpCURIewE
p6gVBmdBUvL2qpMvFVrelMFottDqsTCD0LKPDKSPySuT/eSkxBQClbXT1poRNMGX
6D+XCk0FgojzTzkFCQ7unvMXIWfLcY76WRG5QDNtIqNvzAdUNRKU5rWScWIQRTz6
eWjkir0eWNsSOxhE/ByByr3eLQs8p3xiHEqZUQHfSCwyda2ouT+FcnvDvQZ40sBD
pzaAnOhfhkCFSKQYs+u5ac2qV3pwOQ0bqBnCVGERQb/mG1/j13uwS0SSyVp9AetJ
FU1IaErQBLeFsFZRAwdOS8drI8m+k9l7OAJW2phM+dlNfW7uzP+RUFs0kiZJasgr
57YhDBZRX5a8mwaWT3/hq4QkesRq0MM7ft4PuIiQxOdIpm/vkKDUY6pJWQ1M+Iey
KXLIoCGRBge2llSFqs/EdrrAai31JP8fDAi4oK3Kt7TbkvSfrqz+TLy/Ux2ISjI0
B9sUG6D6mDG+HOrO4r6BCDzdClvBgxGCL+C6JZNzzrFU2B+wed+IUtIfqrblcZsJ
1kDfXB1vEpxCgcD0BKApfO6bfvk1l1PGnlGQq6wjhYZCRRmJcIS81GrWC352iryk
X6SuTlV4asXOuutIEmU9ythyCA3FO/NHZHWXnV0uKZnFLQdvWSFtnbareT41pl8J
OlM2z7psZ3BEN36c81nWutJ/2Cf85bSJbR/xaOZz9xnf4mqo0D/0CT7BP26QLwnX
h05paufdh6d37zdI+nLQTvrKR+xjcECCE7UGaHUvVWasiFE9weachJ0eRes7YRxv
pHx4sVvuDg2BfoM7BZhBMKI3SCjGxe9cpiy90mqUYm57xIoqCIO7D30CTTsVvyYH
ZYaupINFRx6993O0bv/USzCAipLlNIDlgtrq3MqFmTmC679XFn5fcxgzEPruNe7D
hOAaOIYiUbLFdjifr++MCRnWCmHtYfk10XFsZ2eCyp7KvVBqbNek/ypLPv4Vu8Xp
fdATUA8jReEDFLHMClJDJIwfhjfbz01FNQyj1TcRODGV9b4l0M1NG8pBJOeKbPgl
83+l0Giw3I4ec9l8fLEvjJ0e+oKX839Q5fK9HD4zMU80/fRPoViJqoVglYlOXh/X
8kXC/ddUIhcmxRLqiNlbpQ5D8rzsv02sBva+DGymen1eC0/CgUuo9idw/PyYUX8M
Y/j4R6SYJvMYz8owsB6z42IIeSv+ZkKHGR+Drkd0NOEQd3Pf9p8SmpBDPosU6KYS
2Cr4Vlj/GFUJQ0gPEoFLX0nWs56DyzCX/CzRUSmuQLXD/8l3aiOiECkxhqFb+W4D
zlX8f3r+XNPy0CITEV1WQgjhTKO7uOzb2DckCzAsU5Op6R5c0ta64hy2a4JtesPX
q57KM+RaqibIAo1NpeBQ+cZmHgwvG5h1T0azzn9nxxwByrOpg3h9pYzKCyTnb2M7
/5Un9JXxPab1VU9I99IBjXllLbUIaaj1ywIjPlRoQxHzw82Xp4sC5Lrt1vm3D+eK
jB51E8vZrQGGkA7f9f+Ocp1bt7/NIJGnAzS9QIotkrD3YyQVfrAS0O3Gxl/hkdP/
uN+IetygIoiL0lJWMW1gJ1p7in7lQteP6+23N0uot0dcYySADimHhTJIF0jJsQn8
wPlyg3L9M09gqcBBt6G/blZRW9035HRHqIA9LnCrRHsLrIPJ1emF8J0ey1hpQMVx
4LC2s+N7zjpBxoGKcNc+PzGPmdTU0C9iH8BvTrHqWCmWYT/LvpNO1xcwr4WsNZ3b
tkWMS+9TH/YsIp1keuCIvH6NTqnj6X4jyX72MpfO/M2gfwtrwpLzkPdsX7l8df9d
XFJCHqIHLPtu0awl4JcghLI5g4g0GiB8ai6IgbC60SgwSxYGMC3sIzaUE3yxsEUP
cHVsHm45gmycJ7g4hmyK9QyltYy/2k1Eb3p/ooqd1ZGnlX2pnvfRHvl2a+iZW58i
NfJbSX6A1ZfowikyVxKnXZj9j1VHnvldi/SbqSm2MogTLHVO9K6q9OcyR9jLVKEE
l5zv66o5mICgeJb92pd4OSAY31CETHiNFPMP+TPpx6AiI1yctRJVNnL/gGECUWI4
xBV0W4AO0EDHApEPUPWWv4rHs86RvuSsnn1r22Xnmd9bGOhJtwzsQ/VOuGdFLG/P
d5G0Xmb1KoGb6L7N3zQmjKW1INi5n4esf3Gb7pl+lfLRU+nWPHXdjWFT+8IX1wTr
hX2JzRT9S0hqh4Ek4Q1sY5C7Kw1d6/aH6NEPSBK6Ap3OoP6e5mdCaCBmo+9y7q+x
512m/rgeNhFcIWN8hzd1PzXkqLk9yy3FgGx3S4IwP+OjxzVv9PW4ecoRuUm9UtQn
LcepwgwZoyo6HRGxBD9APsPaFtSXGNySouHpdxyx5s3ZsoclWc25CjO8YaKGoKuJ
0BsmGT4NO5gN4CWk2l2b5v7IgcX8cUWO/FyUE5AGUMWw/J0kNAQlWua6+nDuz9vl
Go38Np9MOyDuoXxeoz/0IU+aLhdDcIpFynFYGnLupeUw1ELB7qCB4GoEVfCNaYfI
NwwrAsiltiypG3lgz24RhJcRu1nglHi9h62i6uR5Co7QAsKfPfqgsAgo5vDBO0j6
DGRudjijISQrtfkdJWSeFJjMJehuT6LeUR2BAX6R7TN6tEEnE/WuSAZKONEbkNaX
LgOjAG7h/xlQ6AXWdD3bQHgfvGce7r4Qe0fE/obo9JG2eKyJ6vMKIz+9s2BxDNpZ
v0wtiXxVYMBPkjMeQ601oLiHqnxZhqC0jjrJgnfAXAKj2XzKyWJNQGfvtQHQqW4f
vlqXbpiFT+pEjLozP35XudVlOASnPABsja+fL/YsY3BTLGfzf4ETtFhDz2fjVLNS
h7koftKO/c+t/7SBCHEGVBPq0E90n/NysgjyVAjdIu/T/3PT+QgiQi73bjiBriYR
h5y4NY2UCr/kJaHHnTeGgRi6O2soqvJch4xc+Vnl0KvSvp4xA18iuCzuxkz14kkO
3TX2PWYqUcfwsLLa8QQfvuJ6QIY8Hl6tmR5hgKmh+JOz12rja0+5GqITDzSnxv16
QVcRogAZsN4yHr7c5rGKhB5biAgWdICWIqoTEZZI+FC1ef1WOwhZeCQBoJ0Kkqjs
/ri/kg1RuM7FPcDhtfJ3W5493zJHIb8K7TKkG/ED+81RUDGB1iJwWOUInyM5tXsl
q/NhB4YCHMt7odwTUS9ovamhGpjZ7ffFbtM73RagmoCJcZ+iupLAunBYFpSEYlZT
TcSDJvVv++ygoce0AzWagKoWmed5xtpePEyFEU0vfGFCvYw0S3zLWjJk1L1I472B
FlC+XKriUx1WwQplz+EaD812WvITzROoOMSJwPC9f41OKsdh/hgsk7kD0r1CiE2i
q1Xfn5SvofJRBHvi/6s42OEftN00hDO1rk1WG5nA+NvNUGKFMYeA6/ADdvI/RWn6
dEe1RWu9Db4hSSIlPBFyx8qZRL7iwj3aSCPh+G3VPH+62hJ5BRFpGiLnrg5iKN1A
jVYi/+GpE0d0aZJlfd8kUl2g+Hla/UvgAkLeF9CmFEW9ICFS1ID5tojI5PGGjy93
2xImtbWOdUtH810HJe4WkVHGTG2w5FdAI1rh0NXn6yY+lyTRINibxQVVOB5ixft6
pD+t/+9VcKR13KMtCn0X/8neisESHdNbtpJPxKiY5Ibs1YeiVqBpjYUhVgqzkP7A
GAatlJFK7QSY+JU2xt1BkxLYT2zAANUtBng288kLtLgPuep+tHPmxrEEBuP12x43
6lYBttoK+xEYAQGjlDcWMqm9A3GqrI/7gAHgvviDQTqJTleQWdEvm5LtdHvb8SsB
vkCTqwCfqIT1nej5/GDGe01qnmnkhxDkQgkp7gYVJXIunEi1USp/mmfgmzj+O3vv
opJPDfRejnwsdyuF2i9frP36XxaalaabTKgjP6+RBb2JQMe6QfXj1w7DX9bYd8Pz
K8U93lg45NAZGR0WFiSSiNYZ6ZsZWVyjJS+gSrrfA8wJOKBOeQY9CDjy2ZwWWEGF
2SunPdESiEribV8cd0g45Y9IWcn10xOEV5g9DmjbjX8q4L6mBP93r6q5tY3wQvdG
TKMGTsQD79VxdIKvtMDDdMdxODiShvDkxZvgy2QioTZjm4LPro4PzQ76vQ8Fnk9f
2XlIcDWhz/GawHi9pmzOwa3dF5HaQZ091hR1MF5T/fes/90G55O1lNRoc91xbGDt
ktXsxUWETBURYyck5P9RA8nNJrA4VMLraHbLUaf83wYUhqa4ZoS+so9M2TEcPnRq
Z+Qv6cJsgCPAdB0SYRlueyNTzO7OP2I1BXjoKn7fMJ4b7roC2UWqdjnFd1OpCP0R
2sPTI76X8zWGw210D65KfIzH5pn0QNmRL97eIH55paPY5WKCV76Hjbq1h93eISkh
/mK8xVcWP4Odott+5UmsVKjdVit1KUAkVZjfO5nJ3GmL3IQ/WOvsgpSDiy9nuW0+
ZXO4Us19jGMTFiuenj1zyJcbXoGC72dZ7B85YXEivPRz5jF0qmxM1BhF4uIaySli
WfuxjjHvJ4ypZdHoBDHoKirOt2NPl96UMbImMUMJocvxcs6CVQW6iSo8rUTt4m5v
ez+UvDh1DYQmPnUgNu/e6HxK5tmavgfAfEqD9wFKndB4IypBnqsl9IRuVlO6Y7WV
Za38kbVh2zyHlrXYvpOceOq/D15e0urFQWraNL56Vjprn+mrablXqNOgfL91/vdE
E+TzohNzCN597dZKv4MfARXixWluSn+nCkz5Z5QR6zZ9KUqvdjsm1onijJJrJkey
H1AKrE4xMBCSv6ScxYlSm0eTymISGmvjPrFb1yOjEay0QZGPtjYz8Q5L5+6IoDvF
9T1qPeik/1zCHH2qspxTkr29P0qlSBoThjIuj4Jpd2ojRtRHboVXmdmfVlmX7411
ycEpkaAcUuYXR9uKvK9668l1PYfGBG7hgk1HQ0XgDQqxo5bp2MtKYow9daaeJCkt
NozagNkgmWcItSs8GAznBQcALc6xRJkdjokuA3x2H9iZSZ3SvHnPMWKSKK9UgHfw
mwYc0QQ5JvlcQp3PTzGur/xxWfx/K9724U+xyiQiioQTkBQJN/t8X9gJZbwjsqZq
T2FJ3H0OgHWJrrI9ZbDO7ZD7obOjsx7B7larYpZg9Kb+wriZcNrHM2PUpWjHSc1w
6FO154yYo0Dm0GQVbCY6cJ8Mti0DztzyWiu9ev+DyIMmrGRUyIT7iw/aTvqTO6L7
VpfldlzDlmpyez7GqNLx602w6IIPmfV1G0aJAehbiU7fNwPp9sHeqXj9qzN12VIj
cuHSAnaMexq5yQP4CyFG5052RiuVuc4TtFJQZc1oc/NjHljaE/4NUQSYLLk2Mp1v
qcDKa5ESjRcT4gEZOQ+mwMbI6ZD1aL9tQM7sghPmzxkeakhu9fuTTmwXeQsphYx5
Fmx7yudyqiC8YhRGY6C96XQ0w1y7ss5RdJ9gthAiPAsh6UpJlbIZ4YwTYsMhFwqz
8jS74qnil8yWg5mjladEKGckiuAFEW2QZCmWfdQd5jbc7CXgQNQBFpEN9ZtiCrW1
ujlzG5ymqIau55oxsHhXk/rInuu/H5RnpjvuwZt/Bkzi0Oj+nkECUuyzxxQ7dmuu
3r0FIAYbwifQs6ljypip6SoVROV92C1iNkGPSrwVVx09BleCIqn6Hht10HLOi7D8
UgEsdQSdW5c3oKdd2O5nXTvhAyyJ5bcptcM9JHCMDBIZnY2inpqZEgCLQj0FT5ne
WpvnzkzKRrLSvItYxz+VfpYN8tzRpk7jFiYyg1WBXyBfactjcquWSNjKsdGMeO/Z
/+6DWko7nVGUp4uv8Lb1pP8DXsPP9GVOUKtMhDKD1lA9fRRELNLzkyoH9bzjxDHG
uBy7uNMHVM/FLuY9cu1JcSJ+wn1goHx2yAtAafk+BEp4P6nBgHVTor/CKnSqyX3J
+vB18gKt2zhynBvLi+gW70ULARkFS0FNGI255a4qFh41XE79mEQMFL5MVJ/ox1Ij
3UFZhDLq/9IT+e+Hiro1Tscd9ZvM9zSu/n/LxLBW2mv5khCryq651YN+IaRBVuay
iASUwvmrdp9EL6zuWEuAmtcqCOep2ltamMpvBdtE+dFJjqdoZWl9QCwNZXKm9dCf
tilUfAE3/jWXypxIZuFWSuuQXKg+DOX6pb9gi32HJcYZvilIbKlztY2gyGPiWkT3
OezAVwyqOy02HSiN8XSXlXgd4+1LQYtV8dPkBmv6hnZnnVzOyMidXMCWcl1ApJgn
Vx55tg0LbZVXuHH9P/qYhcaIS6+yWz901lh7uLXsrRqH+l6yAroBqTZ96hFttf9T
mq6i47ZZIZ3rRK6E8kndllQBhYJ121sJNHkRMrsKKX650WYsVv2K9NlZu71QQ5em
TuiT1gBdia2+07j7X8uO9BP0/mjpJc5ASnhxpfX807szKs0W9Gc00lVf0ZpCN9HD
oSiWjJDZ04UUYAEkfm3Pkz44HDmDZY5uY11Fz3UeLaNaxvJ2VqKnYkIizBxp8ZkY
kNZ+kHLnA2pbvz4EiLUhvNzkg+8gNQsRP6ozbIIY7mgC6pxKhS5u0zFN0LYH0V/j
3SWSiJnbO86iVZrHyUZNm0+Fkjb4FCPreXk/frwQNgwjfU+h/hjNS/jfZgmNh1JX
vPxcfjuieJplsiHhbOrvVfS1P3DH15x64QAKpLMuPdaVuDa3WWteUsvhfqxv4XIC
fBJ+jiQ5ov5p3sc+UOnSeupDH51y5BBMt8fXRpALiQZa2QoSaP9pWilLDFPhGz3h
O66vbcOYt25usU4ibCR09qJnxVRdin3QaKxTvBHZGt3oK/oSYxsBSgsCSAMiHdj/
agDVkvNLErn/jOYLHNlRC4vhnweLoU9313ww6sPAM/877rIGbUFOda0oAz/7XsMK
J37pn/C82NTPHgD2WBDfUmIyRgOja0AmcyBdZ1FPTZ8SltwllfTqU0QZFJKiqisc
vt30HGcz6PbF6Yy8lZ6B7a1juw1FpOUNl220ICiHVMmag1F+xxFQJfCwRrhgV1O5
ERZhKCLeTBocXfvLu3VOsQmGNco+U82xlQmHnKi/ln6Iq/mp4bDcN+MUZj2/kylx
Ouk50bgDhIU5OvLzafFa/COVFS/041sKDq3T2fhoSFulK79pxP3v2ghL/Cl8nRy5
RW5YCROAHkQUk1jPpqQmmDy+qcAPZwz5x/Lk6IScr42gw1IKy+Hwld6RO/ska+Lo
7XslIOoRyGtTuR2rGNRNYjDayYMxA946T9lGxWVXsPCOy5FuS2gFy+dE9QRp4qiF
y9uamk41wRfkoqvo0fIKBRmw7lMGeSAT6a5znU0Fhp8oi7KfBRRUNg1ZrjsRxjZK
L/LLt2/gcz/ZqkXmmJeF5y+K/6R7OlaAXkHtwYFMnw9CP8oTGPDrfKumNVL2bs9F
hZDQB6+K1FHUxHcFtFpPSzhYeMT6X6pqtoOGKabL4JW2bfvr2OwgkMeUzae7hQMi
eRAyWeluVzwC7OqxIcmxA89FRGcBom9ud65RlYX4H8VYd08OY/LPLgLwmaio0uc/
XiUDEfDi6gQi55hOE9ZN4u1vWSvrHDGpdR4fIghfvUKAJdKiftZaD1sWG7ckcCd4
/dkF0mFmGkwO3caknF4SUsTX413LcXOYql3ZYLz7NqhUKrVneXGxp2gkNpcfOrir
MkrwPp2FK2+yKlYoO7HWT61xiENMzUmcpX7T+7j5Bm3peDQFWZz6fAZl1pSYt2fE
Nq+rUHdGs7HkBjDRtv7nA8VDNb1leDP/8zCueQO6Tdn8gx8WuQt2AVhbvYHEiRpd
EGiKe2FuA29BujqLgBrRpCnbdY8wMHXbsS+/4heW9fjajMV8UFjP7y0xqD0qcQC2
M/yNDqhAkKYX5bixOn9dZqfwU5DVZ7VkOKzq6otpFxrup7CAbz44bgWSPJQN063+
NnwggKPoi1/aV+G1ceD4VUybOg/5NwarPwHBw2ZvcJ2+SNxg/zEglH5uU0iigBqE
gq0u0C2COARsCGmK5wGI1Y9UY0631pwmZiybRLtKB1xtvVrfzKph2nj7nf66C+zu
jshebThCOU3CdtanPO1C6H7OeuxSsQ0zM0fQ1mnmNSrOfUWVfLxwiqkNsawvbXsE
2j5EiXe6dLXUGkqJTeLkX461bpe5SNIa9qCLHTKat+bG7ZZHKr17lytDZ10no9Hx
tOIzWuC5vuV/S1fKr2cgQl2ZzxoqxDZ9ZcfqWWDG9pyWpcHGDj3XMu+Gveok5muP
2BOU3Pu9HWE8ZisuSh90TbX9C5gig/9YQ/pRiQuDyg2WUdzQ4gXo7G38AoVm8gt2
qUri8rJcM20ZqZahyGKmhU/Drq1Gi/tKr2Qc6fPabtzWa5sjCPL7BaJyMogMKaVF
Anc11B9Ay4ywrWmEQII/31jetKt6qutZqrdYJaq9Zx+tkQ9KtzkHC9M5dOAdNcJE
cn6ADup4rWVTCf0BXeL/E3gvQMYPnOB/MFUYeVvVxWsUIUGmoJM7xFibIaMP4OKC
ltd2qZ6VEHskOHvvcR2lP5PdfEEc8GBWxnyoHD2+AcRKxpx2yjQnXZxnln++qMB1
xpc2U2vpCITOP8gOOglyITeykZmbsCscBOfHLpLPtd2kdmLOYlOsPOSHm4GxAtzY
d16LlHiCJhkUqAUa4J0gZ46ueyTxhM8wxOwFucLKT6S7nlW48s5zkDxYTw8J8hnv
TTkfDF4PIJLhcr5ULr3dxSDewd8kHymjEOO2LIglRuzz5z9Xc/94NGK1JGK8LGn7
P9jHrTn5aF84XApwjh/DB7cnqz5xR5R8013mA/SMEjsAK3DEd4uIsroWbxVk9Tkk
rXxo3XMETwl0iY/JPSA7noIRHBIbCtpbH+AoL51ztlbczS1Qo4kQHBl8fAmnkbCJ
hZ0MxgkSwF6U3LiOiM2Qz8UgKhqR68X4rOf5TB9x5nyB8/oXyUBgH+TVBy9xuy5r
FvPBpy4k+IpB3LaF+1/cLjgIdDzEoaec/ALluPtx/4Y9Sesm2SemVDUUPYxjE1RU
hBCCvsplAGL6UNbxwhLMpLqiy/8XnPwGdmFnGeWcwP9lig+5n0GMLllUVu0Jz9Zu
2eLgqHM6Zicnz8nrL6HuzEvxDTaVb/2uMICqn5IlRWHisqlH0QLC6K8PUw7TCMOC
o/dS2M6JLG0gzh6dcnPXQGE5O1PMMr5E5Ee6zN1uihZoi5SaUzZ8q6ynY8A6CyUk
ZSc5p5+7PWs7HzepGiqTPv0gqXegIcW36S2Qg656NMy33H/QzdkbG2cl2pViOiT2
NIVJw8JAYNkBhHKM+fRHTLZgQYI7mBLfsYvXldQHIPi3WkfE2sYNsMBTUGIa+dhG
AMLONvvq9i6JBRUGpjDczZWD9XLI7Ovgzrjh6aMJezuRNQlCpRtKp7baSx3M7o04
h8lSQ+CYEbFrrpmEQJ6vs4IQ7Q97xfc2t7pN9QlXNQXnjffpYLGF4cb5UilyMX63
SH0DeWhbWag2W2JGHwPsUu9PpxHHj7BwS7NwyM951s57ULhTAuPsdtUugSu1av72
Vi2IbSVce0UDZRFEycUefSn5IIVItYTLUxNXBSLfaxxm954pzBXvS6Cs9mNyJ0Of
tjqAr/XywRfCMx76rU9IoEWt+UySsn76NIE/ZYA2UxV0w93+f/NARzJWe5nBJQrX
mM5gokdxcM9lgtx1O8oRA4+BVgDZn/7pZ8N78c1I+QGrfiaR3POoQ/xNFRzrsyhx
4eysY4eQxcoRA9D4h+fGJH3WSC67kaaNuPM93HGIk+GSfVlm0ZnNyDs34y2atold
L5vbBS5RHW4kDDc5Heo2RsS6xfV99aCKlrxCoMBI8qD4dJ8kiAJNRQ0G9EZLI0UH
RS+WPT779u/i5iNlr0XAULqlkhkgc/JcM/IWlQ1Wv6nSroCh23sVTiG46TjX43SI
W1i4LGYKl6dYBoA3A5DRZ/i6K2YE3P6OaOL35BQ3P8NSTQnRwnxYCe0sGbKl/kN1
eBHDmhq37H5yUBoMRjcF/HKCdN+K9j48+fKp6Pweqg8BR2Mj7e/Ri2eIxLVZXMmb
xTWSMzBqSqOez3KWjAmv+uQAQoHOLg6DkPqdwCrXhH7tBqqaCo6O5Mh0VHDZtQoC
+9r3IZ8Jgn9Cp3zYyrUfHFA7V4hD3TvCj9aAcEnbRgPcVp2CLdtfxyoPzsO0zoTN
uBb8jDUrU/++Z8zcjDqz22gvR33OfFrdIy+YTOT7mPvYA3cK23kXMdar+8sBdkhS
G/hDexsMk5NUxie4Jd+FKts47jQ2n+uXqSSvOkrcTYx5VL/udj3FjyrUe/SIp9Y8
LiI0pl5N11hmPRmUmbpol/VNQOl63D+0ZbDT2fqDCu11FK+MIgXdsIyPawET5482
5ER32brkmMu0zM89SvwxoQ9cVG7lsGZZ/sJOoyyrrgEjeKlOrEwVp5SHJVsFs0Bj
yp4GcCSs2Kj/qFXeBXLnN0wrIRO8pt6NQfQc0fiWwFoI/09qWNq9Xj3c0NbOaAxN
VGbM6IohVDDX6O5B+1iRBE2sirjrGS1Hz3ZBTmS82X8fHKxfKdadF38YyC4dzU7V
EGWn1zPbY3EhZzqbBSp01d4Asj/OXGhFXS7FBtz5oTrT1tC4yBa2s5YxNoqvv7ED
iAPdHxEkL1K/rZLj24E32QHIWVoJ/8fGSUHUfxgIsrpLn4TjAYRvG3cLp5c5Pnvc
3gj9W04B1m1q/dnWvRkiWOM/W/8qMKO07h0g9KDIFeVoTCAVO0ej/GGs/0erEY6h
nxxFtjagMGDgU7KYAc3nyAr1914F6nk1rJqUDGN1esTVzsfeKfZ59H4XDXruQ9RQ
3pLk6tjlqKPc+fGKgMiZPiEv6vQpHSpqIuXzbVC5aPkPNOfoU8IwkJAQBV2fR41r
2LjaEkhx0kOLd657aQDBecRZ6I77BHxq7mVCnKZv/LTrGq7WZBKy9XzRXWIymkcG
9dgFJAwdZdNAG9V8jfXqYc5N//V1n1IybneYG/T2Crwiz7xYBHEiHiWqIZcWdL0s
0HERqJC5TkSSwhRvKTCZnwY8pfv4yX39ryrDQM0+B4n0yhJnZTN6WeZRHxm7nhnK
iOMCqnQ5Aw3FyC7+6xBIV8ErGHFodYbZuyr4tEZpfsGmhWG40375h/peg65pKG02
LnLsKfiOjApxsJKYszKd8G9sxUz6ylkjta/t3Bqcg9ZQBUpBWvFictNunNpLoVVZ
Rlo++a0UvhIH3lDWVbuCahH6aV+60VKaFPwdXK3esUZeT9O2aq7+qj7pGRqL6deH
TFhNDUt1C+KCAYsWtG9xqFBNVSQnuyVpvFewC14abOINQ560y3cY9CHwJlVX9upo
OXUo8bZUS+a/OWDsQt4Nqxw8JW1NtAqzeeV4Rtb4e0/oej9xD37eJ5jitC5Z0588
vtfiI0iuLQc4Vr/UTUiw9mrMu+qZH6mV0Sit4ETM+K1KjDmvfFY7MiUGRTL7sWkp
SL+i1AFs7PIkvEiRORsB2gHoD8QubgCrXuazUU9POKQjm4AZAIvIMSBG28BVmdDs
qmrfqZULeLOnlT5lyiprYW2b474nNyxRyDdcwTYig9gSi8oyswhItMEkYnoiWlwN
JskU9QmGHFb2c8HBjY/dNlujdb8WXTEXkbaICG3ZpJBgyXWG+Qcv/rISsy6n+sbV
eDOKPbycxY+pKoC/XfTEB3i6pNeadiZ9MZKFwTxRZgotDdTyc4zTWun5LglsoyM/
fo+1QnXNrR4iFJG50kT9M2QiWlLOOb3zvUXyFUg7lgq41RmYR1L4aUzmwumgDlnJ
vwzhqVuCS4yogT9bs3QEXWNB3LEGuei4jH+Z4JeoFuTgD8nTJXJP/kNbvaHVVcRX
2jdx5QKY23GIQjOm2Ud+NlIQOX5DYpJlfFY2n1MVo7B88F4LEJ3h+ZDwXnfPbIEL
axfvx2nthWHW4nwtj5CUslVWt2eiMEjTD87trYf4pmJ32R/kH5e6w1RXePaJ6Q64
5lf5MkKlbkaTjxHXr7CDQJyLVZ0/HXn11Fiw8520uZJKXCyu3UpJApqcMxvx++f2
zRWb5L4x8d6+jr0lmpyZ5X80Se+obh6ITgG/ePuLpDtN518XYGuDeKgGo5x6TEaV
IQjupk/0sUTlY76qMVNmauacjX+8gWSIO6xzDt/D3lv/M0UCSJ3lS0olk+UAkN2k
qdlAlz6Tz7jLftghwlcbYmBiUP8DRVa+gPLMc/FedKc2eR6UL9pdpIiw+a8IVsK1
vsZvBoqPkmF276F1BDrpAD7VjGXP9RKwTtjb8/zcCHbLySS2ut1MF/EdyXa0LnqB
rBsHLuPPXZgusNJG4rnRdtDuMQpBtc65yVxWBXZLUvsqNkfp7FG0Ea1UHkOWw/Er
64atyfGcWYqSbSTu23nmlYvbG4V12YlimwYhlTpQfEw2R+Y2/BBFsx7hGLX6qAKe
rJSaYfldhIXE9+6bZKjzVZpf7WAyilAyFd14tmL7oHwr9wyVq/Ixx56yg8IW45kj
biduioNtCFxRI108jvimxNOZiDu0kKWfUTYr+Xdc/pxeBxo9RRKwb9TrV2/3+TK7
QYKxRe9mTdEIHL0UHDarhc1pJPalKQliBflJgT0Hhp51Ouc0LK/u/6T6PkL2CQaP
vEM6IjXsBqgEPI+mgpv97X5+Hjy/hvWiZPuVZujBWsfO1HKjRBE11F0OJ+Iu2uPp
w+0bdWUhC//7TCbkCK4T/pJVpSj+/lNEw37lDWJkQLOtUgaXUXqhm+NemzCLSLbw
7NudkuPAyrH2iU+BWx1i3APV+E9mqhyQW1FrnaPEPTKVf1aMLXCVGFXBwgnj+UKs
RHo+9vTaGZwEzCK8s+lCD7HgbtVvwTifJboAMRanF+vNVaJepqQobrl4fewH0MsX
c1i0W6nR9/9JeqMQY4vJo/q3o9fDlBygUMAnytRI+vmtBWS7DzgYD8iOkfLIk/9M
sa40FVEBSgi8VmWTM4HqKGoDWcwxEv2fpuhN3OXbUuZSjelhLmtwAfUJzvl2AOHN
GLXmELTJaAMoba/7mFdcZGIHh7scN4y0WvKTVVRvUX6kSrGGIx4UaxtavnHwpYUV
R+8bIJcah6UV3GKDWWnEfybhOYIDJL2DPyVCmjKwy2eBNSAqVhDAFK1WEa+pLyJ7
z2/0l4IF6BkFZfD5DSEd+6AA7zC2UcactSyeTU0//v63Rz49YQcdEJYDLQiefNGc
GnAYzDrj5xtVTePdF7wBskRaMC8+TCMWW14VxuZBahgMsMJinzB34LWBQo7UiOx8
/gewR4W/J+Z8XwrH4/cWzPRUBUv/dYBXLfx77PgZIey0LcoN7VOb5Gtnk8zNXRwf
shMqvPz4EPACSHhQY6yQW10Oa73kWsB8p3PzJCRmJG4Yqo0bFKiN1yYzgW79XP9m
cwWS/KoiOTF9ws5gu2JE82nTwC9Ji9eXtGZqAJtzkDo4NjQ3Yf7IphfclH6LCKVe
rBGQa4ZFa7LFSobIhTf2m9bDMWOjA8VvHaLlZkgRp3cVZztIR6LViR5Wct7h0r1N
PrT+sBUitgLL5z/jJXk4vhRlrOOghzhwqCr58bkMAC65o8tS2Etm98X9Br/rrIje
mFUadLUZXP8vUwg5MX37WqlHILAuNvR6AmQ+YU+HEejoIiZv6uyrvhoaJeN2qKUg
AvnmIB5orWpgs32Nzb736S8rTXnIIHHBhOKJn4uZX7m6kVU5EFqBgSP/GRBjOoWd
iSUbdGutzQfYKlqKVfsr8aC0OsltILpKfxaULIgtn0rPoXgSjRl40mXJnGKZihgp
vdf7/R3MSyVD5cq+c9A7ZNE5ubJn6MY+LyiM5pQ5Sqm+Y9P6kon+/V3u/fKyO+7d
zYHQerUtRpx9MCnOSJeSqzOXKqg6JbOhZQZoycIlX3UV8YD5Yh4SCqpNkRFyr4M3
2ddMVuJB4xL5aHZXVJsqAMNmDS0pQAPY8vV+2PRQWLjYEjMVIkepAou6MrjJPfTV
jJzZkpaVpq7b/MPeatmvDCNSNIf7nCefTilB4FDVwoztnfb654Kc4v9lhX85MWvA
r3SoVDS0/Y0FEfdwUmk7rYRQ6upXrXs6Fh2v3j01R9Yw1F74dSQvAkuFoyWxwk8A
owHt0zsmR/ZqtUAEqyp7e+Wl674CT7cp2bDmvjvbbOQG0RSsCMOBnyV+uwW8fDTj
qqvckkMY4ejSdpyF2vruq9ebP1I0kpmlqVC+r6g+0bHxYaC2Hym7aZ/63g8uM3wP
Ha+ZVLdv0PkgmCNPr7Cxabk0rEFSXNhUwjMbK0IZ7BWSAPMSMTpxZZOWr8w8AG5C
guUBkjFup8fubYTqenQ8AMCQ9xLxOqk3NvqUw+7Nd+32bY19wVu7Dt/sZziksjCC
8OPiUWJYvuSh2Hga+FXC+bV8ekiMMAh1fQZ6gUBSsedXTa+6USz3lI/EZSuexDCc
lE0NShtjSkJ36pkj1la2RvzkB7Qj5Ylbyl+x1t5PG93jdLO9rc0t98E21U/udDh7
Uhd2viC0W9RGzUIY3u4Sgz6kFuTNZR/ag/SXcnwmTsKib/ZuHen4NZVUnGWYMhXG
r86T+F0Zf8pqKT5KN+HaGQEO8QUWmiSLiUyFEKSBvYgB9QI3gR0f8XACnFDPCa3/
Dwy3K34K+vAuSUn3BeMeSHSB93BL2GU+F9TH1MEVtJIgGiCXeRLNzF1YrSH1Yg9v
BUBrl4Ez0FmTwpgrCwURp3TCz25/5uyYsZtxTVsTzX6ttDIjEiZ5mpjEVWr8/AZF
IBknWUSWcVZMjmGays6E7BRSAaqT6Ym4Oj3udOojK8ZrPNuuZEnwKcU3Uzv/vDue
kjUSWF1iKrCIVSflhDjU7Gytqqu1KAait93Dd5YjgJ9Q0hDX7miGhUfTn8v4m/5p
QnAtRvQQvqBJB8qQOdSaw9fXoB2W0Y8lpbyngGdzHjsDcbQHfQIOrGrkdD0cjkUF
qiVYIG8I5IGMj8aWLPpmEUj23W0VyCtglV/wOyA1330l+YNXncX5sjW5pUGDlhnZ
Nwl1JEmw/00UvKjvlBDNavVTlMa9/yu/F8+xYicRF0x5Cx798soK25dBD6G97D0i
D2JdnfGd6awJfU7uEdSfOSekWZhQITqDMal6R67SKM6AVzSd1GcaGM63sg6jDCF8
c7VgQVVHgG5Ku9VtuNVII1hjdj1Coyc9+PTpgKu9/qfbN7w5Df9tV0NJrGT3hK1x
KQhbsyDv75dnFEmVOEAqxRR2ZZmR0XMaoRi0qzdH6IjHiNbL+DRhTga1Y26IKCSl
S5ULyh3osCDmkFruAGEtRSzDgswDVvbEdczvD78Qvzxv0Qaba1JpkDY8Wg2sixyh
VGp3K7xJST/SsESBlT8XAneGW3U9seBfTIDDgWHmUvCnwvVLVbV6P/KoJEpLHuRu
Xy5eTO058exY0nAt5lRzr09peuM+dUbzTquQNI4RYc7VwXTfPfmFzk5a5gZRDTMl
2uApW312qVM7ag9o5w1bT1JxsCN8ngd8/DdvBazHMWL4Cp50vYsE5mM4DjQOXi8L
yQH1otcVkkbEOD+SUJJqHNROVbzrzV5KIXlFvtQlTAUtU4un51Ql9OdH6cF6kzZE
QLHRhUcfPFklDfJbhLmFr+gH0F0vL4WZBKnwVhC6kGrUiIGk0NAKjZaz3Y9C8QAX
PZke8g3PPXjiYelpLR7UXxfEPdyvYFKTaY1tN/AuXzdltI19vsy9nPLMIoDcarxQ
p3BbXrBwY/0s5NYLW44ZkMRyQEV/lPwN2XEYwGfJlVjT8ADCWJHJ9bQEeutPzUYv
yjpgFPCZK7SkYgEno3AS80agr4hTBqwXm9GE3KEzPFCZIzQ+oR7amVioybas3ecR
vnrnKfBiymYtEb1BK+7/SgjCaVyu8WACKla3QUOviXiB1nE7ynSW6caYN2ADpaS4
gXwcczYiZxKq0GPTlDh+5HWsIUrBMK8xM2Pv1LF5rL7jivDTMnHvkEMyUZPrYwFh
+J5G7nB5HliZQEUtZmc9tUAKlc0XApEFZDEmXauouYPqjgk1JFZD6EvVLNEmtxMN
T6fLdHRf2VUdaqy305MaRMxtRb4+zLFnIqiga4iK1hzhxPAjdYlneeQvaa6yh9dH
lDWP0JxgdJJMILQb46MLRTEOxS9W4tXiDZ4P/gqfw2dkfHuY9mSPd3JOhI6/riK6
aYe1wl3xo+rkmZb7HHG8615N66+CR8TKlcV+9wIw1l+6o+tNdIrccocYPdSqQAV9
ecs77HGn/3HwXOPWfBIWsFAM+ao4o9JwLdKQPf6HoIEw78kzCVihB1ppiovO0LGK
5lCH+a/+FxgaCrTPueSALQwUSfrvlf+fI19tHUx/tjsZYTwe6wtnairqpQnN/gMy
KwwKDudrDds0gFQmzHst31HHazbCDEo9Lq6DpK2BRDBrzQn6E7Ir1qybM3aWhxBP
CHJdAnsXq5sQgSDRSavJJaUK7DBBXRkld3y9WbjpV6IeGEDBehQjnZqhDw2mz8UI
XEf9xPsSNqh+/43UxtlfKV/GB1c2akpGlWsqhw1obILElypLGu9bB8Bc9WTXm0Yl
1z+MhyhIZNC+3DXg8do+s5G/ieqKKn6fP4PTRWxkxuZtMSVj6Bne3MlCQIK4bfAH
pj2AIxJawd++A6ene07i6oIazln/2RDaSgVKh0H2xVioEaB9b1meSz03o16x9BjY
F4AjHFzXyi0dfgdu2v+PmCT8PG0xFIVZJTPy5aKczj0nhCdyZLGMC4AIXclKvfCD
YX+N7ignGH2FrwMNlvm8XbdbOsVbS5E5TOgw56akyrLTAP41lOieZYkm6JE74VIU
unUMsK8iRgyO9YVNUrrJN1JoxfUXQUos+AU67DhD+wvRnhXZyEFgNfbvk+4OSnXE
/DdE1ZGyJsHkkFU91BuUqyE49C8PBwbPGsmF8DSgKV2gcXiCA10RxTj4t7ter05i
RT7EHZQ6s1PgqFnrgrzi7pB5MCyDkhy8EqSfIjS2KHONOBuvqyq5Bu1qjjLIhYOE
35Qykazz+Bjvmx/cShy5rNZDIXYg6hreV/KnnMthm4w5tplzCX9UVA2Y2iINcDY1
Rol3FZhftrAPAr68Q5lHeD6nuv1Ut7i3DH5MORgGE8NJjAjQtFO1VUHOp25m/m9j
GJbwau+j6SEEJRUKVTLbFS/Ym+k5mPTJvL0fTqqJQ34TtNmJBZgqenJ07fMsH2DH
I+HcHS3hGkAe+tL+fam84JhSUTiStV+5Ey+urAd/eIOoM926UeDGrx6HHBaUNizJ
naRigwQrW+iNNs8QzT1hiVxmYqAJ4I1L81O4QtVFPzr+xiRtTmJ0NqJ4ltFGhyLd
Nwdm1s2PY9BU67ilBxgeTrTaQWW8NT9kZPKWV3Ouj5lWGqvDnlTCXymA46Ys+l0y
dwFOZ1WVk3sgQyGtH2lU6AtmI9GA1Yji+fwqSWBj7Vz3FLYgwzJp2a7c86AYHXem
yJB+XS2rX26wLw8gd3i/Lb08jBP+synzbGev97U0xbh4hyVZ3/6RmbyTRl9HmRiZ
O93k4k8QXr2VcWnyyLsTKZNdVmLgxXOPSwifkS4CXS+Cipez+YfCH72eWqYbo9D8
8E9n8EV7rCvIWRJFo4ftiqUWTxOWf6TC3FBMjmFSu2Sewei1dPCFj3iuIWHKqtsS
MfI3tam39iBK9gx6nnh2r3AIfnVt8dRcKXVViMWpAs0sxEDw6zAyIzAbypibkz/W
6BnEU9GY86ve4q2Cpiqv9Q8h352/onf2wZ2YoMudtMycdxz9tcGRTmf3ADbLTeUk
nHaBRXYUotqy5ZYSp6RSz7r3hi8v/D60O3Risuj2mSW1x3LuuXWGAgvranranXjA
7hxXe9/qIxsgiUg44y6XEnVmrNnMkjdWtEioQiGW+uWjMr5lX7KHA8czh+gaGobe
YBFq7aQLIMusm+rDJbGK8OXRAT8WvLoa6ctQslzPFX4SHv+uEEQs6oF9YWGfcVPT
eEl+4Sc4AVKJbIRTWfRzjQaX/HBozrVVYViPVI2f/Vi1GmH+U2xh9VqE3AK7jP3T
HOBCrK1d8mX5/HSWNBD4cdZST2vLMh/oAHjZ/kWo7X8aBP+wA5l/pkjuy22ZYuYg
hx2ekp3J+VrCAPyVlM4fCltUW5Eryzk6wOKswzKR0TJgQRZEezvER9dBHZ2VUpcZ
HJuMLS4SdGfp/587akFmyP2d843io0ByTyKoOkPgCiFd57p76mIjy9hMhM+2Vt2R
XLLJ6Lf2jMRh2ioMJodAe96czfKtRXnhYQXVweYKVGJ9FA5XcZVvbgxGOUhID4AZ
CK8h7yi4QJURZeB5p76gBe/GyW+Qoo+nLSjQUl4q+1U4znJTJC1XjKfZ3XHvyOcZ
NewjvWuZZ+64M6F+2t0MZyojRb18THrHJBcLaYZeMVR31qZQnq2HLnFswgAtPCA+
G3erkcYC42U+avfRAo8Y0f6trs8d29O8SXjUbYLVOjSYvC9+d0JnZcQBuW4YbJcN
4kncwkmSubPzD/6n8FYIoDuYwWcpGmyTiyZ/QoWVw3/SP2ek3gMXcocClVHjGTSb
XSL9oxjJ6V52PFpups3bqMsmt46IB34/9xkCzjA7/BtUIMmjeYAL/d4B0R4/OK/f
/8gm/K4ZeTFJN2G5Cfk9ioSOJiGAP5iJ/EmUgr6q2zKdpWDdUIfkFruftKZCqWMI
JZf72IXuqWpk+cDDzlCIIUu8L5GcqonwHux5CgU7A7oxeGKyZbvxUUn9hN3tDw0y
tJ12B3W5F2Cl8vVCwQDAWyv6zjboxY5uoE/B+4L0c4km+QJdVSkZJYkAtj+5qsGH
bBSz8tBFRxrwedNhFnkG3MX2iV/A0hUpZi6GstaS1C5ewTlI/ZFhpg4798vcgMGP
XD8H37BRjVxizA8evA//RB4G1jXn3jXItrFKfxSkwL6rnTrXM7sPlAX26LO+sXbs
7A/OtnPqnof8Ak1Sei5BODi2NCoeuIVZVhuX5kyhpMhritv0QMlR4YRHn4c4W10a
1EoRvagnY0SXgyAzIplt3vcboomu5Obi4/LhnaIpyn7ua+33YnxOAFlEWj/AmWt1
lankIj2ye9d6WmAcgh8qQyuoFu3tAGrkdv5Vlu67+CLGIUWhDbss1wZt6M/2Tfvr
rHKA1N4ynAiKHgrbkqyAImWd95smrt0Y+EcYc8Dp5eaRGRdoBRUNsiROXrEMCofb
UHtDEZclsEBHb3ddCbkBXFy9H/A4YODw8suMNRtHeC4lvzg5idU2uBlInll1zLHy
Znk8EW2wR7FhHwJmOFzD1ul2764q/JVxt9HuVbmXOBb90oDobJyF8OTSF7T5rjmc
4vT2U6+qOy8C/kTSDINke3vPj7hN0shle8jHxRYN54SXcm1b/frOCWvBZK8iuwUt
Fn9kM8JEhiDlEQNpmaLylxArSZPuxn1pE48OM97MZx7WXFewsUu+tJy08163FsS0
4HzxfI+Sq2c2+GKDxNcn4T/nTvWVSQdXa8C4b6AWPvcbzn0tgvpEXu/uUvfhHKDL
8yEfcDuWT9H4hrOdhPoELLMtwP+Qd3AyTTOprO3CTswltMMld83Y1PHfIdC4XYyc
UDRK9qyME05Xy+3lJZ/K/cN30v88X2EIVCmATpE1LrIionw7bWNhBWYZ+ynTdQXd
pvD4uJaS7BuafqTYAS1iCWqj/w96Qd16M4asaJZ+S6530XKU0EKWqc1uICNRGP9i
zK6la1fYpUeruIsk1eiKonu2DDTXNcg/qWCVgR+0U9tKtBfYXkGtE4nG+bA14/I+
rYrStG7pC1G7AmEZmBVFxEG+eFfhpdX5ZqhuZrJZRvqNXkNZ5Hj5vT6OTWWQvMsS
PXOMZhAvPG68Pk+leSreN7zp9L/7rIhatgMoRX+wweJgWJJxfmYepSpm6RuW6ELe
f6IJZ1Dh31n4n/uRaXMMeQ==
`pragma protect end_protected
