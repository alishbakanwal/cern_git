// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:41 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kqNe1geTqjULX6TJv+YPiCGesOheNng3hkVNStaov8YgjDD3AFt4VqGGKh7GtkrR
ku4L3DNBKXgLpj4Rmy8r4Gmaz2rCli9CPNOAqp8YxEhLGpJoa61troRRg+Hnpkni
qCk+H3riJnvmtJxSrVkblu24OzDxeSMTwE1iIHUofJk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7312)
r3nylgHpuv22ATp8uj6TGXPKIhaS8MwX0piN1a2iJhX0H37VzIYtREuLFOvOfnA0
uKSkyf7NRlzZT4+vF9HBCaGudISKJFwLaNCyB4wfBciCT1z8RWyKG6HbnU98Ivus
xzNY29xqoLE//W9P+HtwRYVQ5HdE2J+FUd5xXdaAGAmlqTXC7H38304LYif+qZZ/
44tEzhnwvheOcTrqyGNHixZxt/aWceKi1IOAleszSM8lYBtMfd6yxuXKSO5nWn7d
XvPqOfy06CwR4gYJhyi5sjxNrNpNII0IFv0QTdqJbS8IDAm3Z2tv283p/gVb9b8r
3z6xs9ztBVNoouqkxiuwvTSqluF/S7HI1xyj6w9iW8rw1QBE+X75ttzxZ5M9d9fK
seiOAaL3uSLve8ZOEki+7qXFMa4/zcN9pB982ri3BpB3fpaJpN74APAzAdYkkMjr
Byoe8v6qaY2wWJ5Qzq8uKfnCiNIzag3le2M6E6MTS8vCXCJVcAMUhVV7yuP1rEu4
xzZl7MEK8Rwy9wLpWK4FqTN093jk2VST6zwJVGNN6YiP8pht9nQ7rJjMRDGdzgFf
zF3BTXC3xAqvSnEwFBic+hw5mGyUaF7q9cjXN3R0k8iyHyAkxGSxIWTuRcf+koL/
n9mYWyhh6OaH13tyQ7i3OK7tVjAu66ylah/scQqC8A5qDAOZqjMv8fAQ3tW46hth
kDWMeoYFhhfRuSH7fQU/etcyNdKtUVYKJDGthZgyMNJJJB91tmo9HyRqDVm+fh4u
6Bi/Ri1nyz/GpvwAmWLWCb4SP4aubJDMzhKtvBG4CMGsyYo9CkfF4wqX34V6bOsR
aYJdCJSjpBm7NOlwoiODa/7S4kTvHLfAycRFTvAwUHH53zBADr1r+okdN86Wv80v
ekvgDCHzkc+zjUJd8G//rGiIPOBXxYfoQ/AV/kQvT2Nli3opvYszCq7p4PaSnWQh
AfW/ub1WNraowkaAgwf/Y30Vu8fmxjsAuOiAGfLluX2556MOY3tRiAmBkd0epJs+
1ZRahuFX6I5ThDX47cwh2+FV0W4cAJTN/zKw5WN+wfT6WofUjcu1hyu9SmS3zbO8
bO25J56j6wqhstp4gI3u1Hid6gRsHNUDDf9NHZb3RcWQxk2SmFrBuCoYWgJeYdG9
bn8QYxNTh6SkPD3rAhepRJtNRn5AjCFhOGbgpc3uZNhvnlFRWnduoc/oqrje8v03
gJTmiRs9fYBzUlqQD4UUIcZf29XQpOWqxcFs2unF4M6NTzThXwD9omFK1MyLI4/Q
vWrOIl5+iASTbW8+G8f9o35Dn4mW1BRrNM2qy+BwTPQ2FziqUD9HTHwsiVsKH4Hu
/O+EiaczSNhcpnEaQTM2l8I019ad3YC+aBOBwnKcqz5Xd7Jizi6bLbYWucI2RF2m
J40R4PI3JLNBQl5741ZNRHxte/T9hmHKSu5KXuS04S+1SLH4ZJ4yzPsUoumB8EiF
pxQW/kpzTz+1PNYBDK2ovRGIWaE4TYe2ko+Y1yghx0LWQMEqP8gYmhXEdjEz3IAW
RV9Ti4OX8X7Vmv1YR0FUjK/y1522WCC/5GP8pgldlXphrluVLmwXp/YsNydB4fcC
j+PIc2X9TKwWRpaHKQzs6luHpFpYEA6snaRwSsqMh6YYH2+KT8XK1mzdlKh1bSuQ
+ROUQdIjh6oxpebEzRDn3hBAR5j4h5JXcs5u6WkjTZdJvSqhF74nOr5hfjeHeTEj
nO+bTfae2cMOTAPAvXR0JFnElPZqbUPzdi6+IpNxrEngJZqn8DTQEDVxBNzSCwM1
PlwdT/7QeMZLSx41HkqC5zVH6cPeO3C40Ni/rY34fWwNQs1wwCtVKITLJpZPUTUG
LcLkKIGW53LSmLpbc8k25rgUs321wi1YVDdeD3Bb6C5GQV4WWDttLFuu+noqmnsL
bUhcNj70+spB1nYUbn+1LlPWkeb6kViaulwirXicTI+++tePOZuuUsQh75Zb5Axd
+pcTsgmYWUaWDh5hw2xverGPkQ2b+KmCJXUHUzAwQBEox7VdzHdIa6zoyboEmnhs
cTg08XArjK5U0IShAwIPmEYoWuRYE9TgLaiJ9BZg6i4HGQ/Nczoj837Q6bRq/s/7
2GkuVwB6mRRGzygN2mnMqjTKOdGN7hTEyTrDTshUVHQRir718mQtEcl2QyRFYiiO
6IzFVNMT8N/IGsbG0QuXJQNFFIxrXQUDu7fI8xITbBk+oonQG4lAhNF7ukugI3cz
7cyrrRbkt3w8Rkd52UXAbaQ5I7x0aSw6Eu6uKQllzXZ3eOKPaAUSzRJFoIisyPk0
S/ZaATfHNTQ74KEhTbOSMnOGtz8srVuQL9s336yh5C9Xw4QltUWOXk3nM9ZdpWfG
uHwJKi0Nd+JmbgrBS6EilNBIvRSHPShJvYCWqsPHmZYotdG0FXar3scWiS02fl4w
dj3ocUX0iDYgdeaFuyTsMvUSHGmMry48TAp/PlmXpZMQvQQuB8xhYdAm/88ImNK9
ksctd2zh07HJE3VTTTfFekQ5BfjrjMvw7RpC8N6DkzC+9W9KFrSGwOeKYG4zbj2X
PJxUmRvKFmcS6y/kBWmb7ploeQwzX4eYqay3TBJlNgTotfKs6pfoXZxsrR6o6fAB
lX8xH3/4TrkDemI4dQXXJDMvu9plbRhYWMQ6Po9t2tH1lQbswnpN2l3yyb3ZvQlW
6Jd4lp01Yq4o96NqaV0627tgiXGokHP8OXP2Yfci3rQ3Fkp1Xfg2OellDPrm9u46
X68hzIdOyO1MEG1XYdSOvnIFbm8Muj3Di9n/KQ2+WaPCMVYLCfO2lttL7h9HkBwl
HioaxCx1x7+YDN2qGFSorxYPPi7DeU/sHQACeEREpZeSChBHEpKtlj6lnZVryT8+
MX6gEwdYquZneitzRxbsKZ3wLg8ACWSJewxzi6oalgCQOpyw1C0cTaQracE0wkat
i9eoQxXkU861FYwYEOh5/7gu9Oa6Bz/iNtHiUtXTIl2ZIXC2mADWTlq1+i/L8kZR
25e/9PX0H3+JK5vUv+NBK9qolbrtVr70iUTaSNEu+A+BvQ0jt/JVBPD8Fi4kOKJ+
6vKarbEjVB4DLKK4EJWDruDq6dbOfDs6yrzaKYduc4blNN7zvg347TuTY/gWaVkN
fFkNmmGZc1BXDhs9HrX/aLZOrFCemG9bvjAi/lxeFok248repS4BLw67EqgqXAHg
zelFW62Ed6V2vNr29w0k7q46QLbcE0EBJ3WHWUWtRJqNOCGaRkbgZxObm1oEDEN1
r5DfhRpu6PsQ53W7q8O4k/QHcOmSC1cxLqCOvMbq31Ku/BQ+hhN3DM/iLubn94iv
T3MZVXMgxmqtwcg2mXzATe1uLYiCV263zM7hog6L4Xy/8gsXxr806NvZDHH0PEgc
KflE6FMssahhMIUDyrx5hTu9e0k5wgONt5+Ne9yD6+DFbZSd5KX4/qWAxT/upprx
+itg/MDRWSUEX3CpCWmlf/kGR1vtcWP9zlMidoLwsjD9yixRqUckQuET6ix+/2Vu
5Oqfhilzy/boF4UeilrGlE6wt9YD/PvrYbb01CZyruTiLcFjtLNs/ApG4VBe7LI2
D7sNvqBMGkkq14v+CzveqmmjN6Ck9Crgdi40ZCtsMs6aULy4tvTZFJfhH02ObQg5
e/yajuqAnkZZaTTb5HRtJLlxbbLl/znHm8Y+sQ2vf2CHZxziDEbja61ZK7ePcg4j
oIAcgJSrF5XHM6Uw+F3hNCd5edp7EQrDDc3DCu+OD9K+vGPsFq+imgmQhia85Vkl
lgZBwjcTAg8UazcdKZ0OpST3tGuA5XINnNd6qdE6zVArPCQsl+sB6bSPN0GYcNY/
dSeZHHdPBLYwPD5eAANzlMYjOJrfKHJ+IRj1giYYZ0aSDXHpIZsl/CxEfImtU4gO
IuNsoCZlZ+YO1icrZLSfwhFyb0csiPwJWz6+N/sFNqMDHIqfeFFJMyTrPVIWb7YP
H91qwHpOeGBYtoa9BnYSpzVL1glcu12sp9p11uAca1SnUN+1OGA30XzfuCRA9wpk
DQPB6e6BiQYJibFB6oLbxmysJZQYG0Yx/wdDbOn36dIA6YkrYlLXkl9Xxlci4KgJ
bfzRedYHbX8vCsjsgMnYK38ovCv/xPKQ7Ckxz7VeUkEL5Q6SbYo6LsqlQrOsE0AT
HMnFdh9gemVtZdUMw31adfyJvNO5HyoyflfBAjP92huGt5/NDqPsoKX/bWlucom2
G0JNHD8R0Ct/qqxig/72aKyZ/hfT73G8AsOtvzIMSQ8ex8xisPxIneRChPtlBFkP
tE33lrIqwOgnkTp/5bOp0Eqrh2PT4wxha2O1FcYHidcy9qIkp1NaAlm2riGzWfZT
w2bTbNXiTJWgXNGRhkPRSu3e3BUbv9ASqUFcWxocSHIPVG7efjUxF14c47hYCLBc
uJnfAFfU5yl7UOnXtFIy3bxlmHB09UuD3jHlHsja/78LA2wqY0mGnnMXmojPiWqs
5k4/iB4lOvq/7bjv8fttqDyZN/naEC3iP2jE4oa1PQhwqkEsKfxvcjjwpKACYWFX
txTXRz1z1Z6ZeuKFovMfKzI3qbnJidm0chS2ljyvWDStR/4R6bTwI+DztjHNLBlN
ikS5gxa4U8A6rbWmBkojgP8oWVD3oXKYuI7TT5jyo/97s6JSInqEWZjNoHphy/0p
hT0pIOeekAIsGstNajskDeBZ6StPaAVjF36j4gRzwMta+TzA0mgSp8jv+8OXOmXC
dxuSGy1UUV9EEPuWTrJqNRrrblVoe4Hj7VzFlTB0YRNOnSt8XQO0gwl3gSFHLUYQ
wanzW1zgucNv8iFldGADkqy3C6WymqXB6ATfbkkTFlddcFilmBjXHRDE+2NJz7gq
KzZHT5qOFBO8HFyDh8ft1I4Qk9BeBByQACN6g5IjYL1fDqU/afc74i13MxKuEsmM
wGl3YhlaMKIKoPIeOoEXkM71Qjztfe0Ns9+CvpeGhOpkLR0fsANq6L3JseGkWid2
NBbcGrQdVeADUIkh9dA+njeVDhbQ6Go6BVVt8AVl7h/Al6ZDtbsFr1+PC3N7XBdF
rfwykFtbRY7CgfgBBIK0jLJW0TJlX0smOWnForqrEl6pyZzBr47gmweKcYy1i30v
R0MBf9P0ZRx4fKIdlIC5o2Cb5wprbk/HyLelBfsvUQxeOc7KfrupYYvBSIR5Xeyc
4tKvExRITHXzvY/AJAX+DZ7mBrw+ffuhrAAuJsZdZoT2UhM2Aqa7FxoNojpJB1kL
r/oI3K80U9/Rh3MCTDEEinU2MMcvO4SCzTpB9S57fi8jL2QbGniQYt1EU1UlVZRe
tD8UOGaM/ucaY8jQfE0DvUMEsTo/A321KdbhGSS1+Sewmifn3zxQm/+VKETRB7Io
72CZSY7EPEunWqXL13XYg1igaHdpKQRDuRFEj7X3PBPBcXTUeSyX1iaIFMOVQwQh
jY37pSKPxKzdzmTHPDyoajGPvjLbBW39ZBmDITnE6TXgXGmgAligRWPRua/EmoAi
d/iL3cQZisSSMGda2Z9q4OCp/ALMIUUEXxkPexF65lbCG+bM9i/loVItrmDUGOEQ
Euv+8Tf5k+EsVRfzWHl+TNCDLFTmvQ2MEIRfRRPPN+mJJxLv5+2v69t1bzYV7hIL
8OmLOO1JIZs7yhASd/ravu1EmZ1E9GGT9in66shmPMViKoOupmm4gCCqbuFKyHbx
FINsgumN4dLFHGV8lWGDq1c1WsSWJP3yPMw2UgMMjfWvU+D6dLoKAu71h2vZ2hPn
IC6/ZfjDfc40yiBFPg6q7Kwfo57PbOa9PQIPiWAgWDCD38DU9lBZaYo7ZqNmBxPd
vCPPh7tIEqnWMND+DsEcPBAEqXl8fr4r83EO7mq2G/JDGdvain4q/xY9LnVS2tm1
V0zIw4a7XWBl2okBXDfh2A/mLFsLr0tAioEDQsUAOBG3kYjm6/o6WW0TqAn5QUFH
mwl8YHgMm+41WeEgqY1qfqtlaNhWrBzbfbh0Y/pFpD3FzyVGiN9Zps1MJWKzPaRw
FRSHRv+8ppylHrdQzw+wNFqK8FJF1wBe+C0AZQWhJNgrzVhk3gFaI8klpH1uvMdM
JU+NILGncO4Eukjfl5DZ0TlPx8FK4copmsNt1DBWzcwH8nWbS+T5DNlzJFBAXpTx
JsSICYikGtbsWgH76e/WMwb20dnvIV6sjAf1oGH4xosXIt09GV2WJLV7rMJpaRFN
DNFwlZSkC1SZyHl+DhHIUZpPwuz1FKaOdAbbXgvLW85pdxJbguYgLlf/dHSmnyDB
ZUtbqfOwC8CMZm3P/7jDe9Z1AXl8rXIh/w2bUly5DcRf5VZJvOKLwzCQ0dSPja7K
ZFdmxRHzKfuRbi94DF6trHi3DSXrgh3crVqyk+iSkzzdyx/XUIZo9bc3cJdUaSTU
QQjt/M/xdt24PomUXOGoxMrDGPk0k66+1OLksIZTzGpNaSI8nLckOpml2wO5Huv3
JrPeWLOXua1eKWt4J2jxLfAo7nP12kaBdu2zAv86VjvUjMCQ2APCb5XfOuAoEm4l
plsKl8NbmoS5jGuRODATMne8vy06/t/Z1zxblvtbYz9r+7oj/csUnj2Zk6suKVEL
/musp99pAyXIfqI4VaSM7Esiuj8xBABC7Zd2KAMfC62FEuYAA4z8vIkGc5tRR2R9
w79FGODeMNe4IGF+dYnly9tEVHQL532s7BbnckHOR2k1pB6YyQTzOsY2Zm4qBLj7
zNVYfHcsak3jtNMPIngoePVjkXq5zP3SGiGYWO2FhxF3PU63mcROFU0vgtwvHqqt
4c3TgDC8xTfVovnK37Q2piEVTJjVnRo4StybJ77X45lRyIBYmFgzfhExpSQ0vW3Y
FadPQmqfsyP2K+7RJS/4jRxuiBmVQvN/dDLeQJIv0HOJbt40ff0AJTPW2YckoBDl
etd0Cnw7nRYp98p2DQwsgeqB0/RcYND88wwt8LFqgfBDLKyKZrtA0ns55I8SR/bt
3WvwNOFDA9RQVXiUTjkWk7sTzOLv4Pp0OKw9XyFXrWaeb491Pc3P3PuzvCjX4AOu
rlsGG82W+VbgQKP2wlkTGXm8i+Edwrk827kd5Hx7KPGofisnEpWB47lRWA4apmxY
r/HIN22ugvf0IcF4tseXH5msAC0hR/F1APiE1boi7jNrkJlxM87QudNIfLLU/6vh
vH1NOG9L0Tq2oMV3UR42BghS+GWkts1fh0IBcdA1js3vidWTqaBrJmt+g0CH9cwD
jt7qLFqzZUGrrZ4dYjLndyogHdAYmvJVsOLvGDjqx3wn8bH3lidJ/lN6Q402EYRi
Qfd2NmaFcWX83WNv/5bPGwuJ1079VrsLDzZnNqZFGuRUKWrn/2vQ6GMdfWSBPHC8
pC/XbSPLn8IiqYZwtCJ+tTNEhcebVzmA22t7lk6BmyR9y+dnPfiMqr/77+sQDUwN
rNLzmdLnso8rmyg0WLe47mvFU1s9bUaYQl13t5cayOjHOC3eNgP7HD9TQEj1+TUA
XyZefEixHMe1CzYgsQyYhCmdNGBB9BAyKVTflcXfYTMtv4eGvSwNVcxsDT4npJAU
82bQEYlk5scBLosTH8CnxtG9rCvoWWzNVaDzCZIAkAZ0Q7hSEOvkyLQrwr8uMdO3
4QfNL7kjkA8Le5O+/5rLVx9xuChfPltsDHGziVeLmP5JWwZGDrpHcoqq6TkuYMyI
myEsKm+JKEob16oM1LCpns/YRjVxncazdk8nvN1lvenu8FJ3bTkQ8ZVApeTIR7zK
eWbtb2L3Gk9JjlFayQ81EWDXHxeRNdkjL8/nU/kek9Nxdyay5eQN6qX+6VnK9HXo
5osjhsbwRqlyQOQXqSJrO2Jz9N8KihgoblHJGA1EneF3J7KQn7wjbL0WcGTQo6C0
yRyyRRdTFn9T3ehPKpd9kVgjwmSVMSm+LV88r5SX6WdfaG+Zus0v9Lqa0S4dibKD
my8MLi1eA2aelhPrdpDLTBhnqMSC64HkrLaY/1y3xhOYID2JFI46aqjyL6DZEi4C
B+fKgPSMNUkmoPY6PPFwHmvZqiyO4GJD+oSFxvW5j5Z6u+lqRlUfNGpCE3Z4B7v0
WZzMlG516tm+daN/PWWRv9KOggR4LsOdp/WIvBtvlR8HIBqq8r+CIy2enoijaLzJ
S9KOfMjR2OKM3bCXUNyoctVWZcuIF3HUSuHq4vnN2pRt57Q950uVmjdAFYcT+LMR
cZyn7DlpABUXaBBvEl1uVAYbGIU+XDuX2y7urwrX1htBRS2i+eFf+hfiW6VaDSZU
ANf25ZpJKQ+0Y+iKsXHsucf/xMAEBeZzw8hLBrxwwTNO4bQPWy4vjeqIVRSwM1Q/
5F7pW6MvDHCv5+pK73S4+fC0FejjC5XaEHx73zLZpK0khp4CO/I/M7Cy+1v6SSPL
K7AW7BFTe881wbQZc34InNYCBDRMVzyRxW/BetvULhX6kaq1sAjXPFTyt1WnGl0o
QNa57gTBzXYPJE16PubC4pn+x6uL8l5vXtx2liMG257MQTFS2YUwnXOG5kHI8swZ
DFv79dZ8rJ2ko3acY3OuijgsUKLpB4GNvWZWRecVoeqY5gqnXkOyx+t2a9gnLjxE
DvkMI58Wl8vYdYQbSwD/UVji2kHk9dE91AVbBtPTeaJb+301GTSn4iKQbkakoax/
ZbZ0RW+BhjCrTxASXO15En7IP4luGsuxN0DmAAgT+WnyMGTyjNwcxb+WDk2LgdV+
n0Xew3WHU5f9egt/nGSXX/RIZnsn9kWEAM6egeymXLjT/AbajL8bxB2asbGGM04m
xFBUVKkv1Q3+i8i7hP7m0vnxa8UIrKlre54cQorqHY/Ngk4jlyp3ng0wJmsZGzRF
u1WN+5L/lWsGLgUOizu566q9IrNzmVP9tsMLK8mWE5zzdeinoLgQPYBNH9rRobh5
51IOdCh8jYZnzzmV2/nIJAdB5B41sQHV8iWG/CkZuzG7bh7bCx/sF0e6uDPKR3g0
JX7aiHa/5sKvkooUQqQPMflr8DkNvcK7PTZ3vsQn27cSTMUtBWaruTygGTT8pGne
du0XCXrLs7Uzzw+qF40qOhx+3RUZ9WgZcH+IkLF26KX36RnPcfIWODx01zCQxdUm
vPk8nE2HxZy69sXOsGACUvp/KxQo0kjjrNIXJhWzheiW2kyVB19ImKu5d8rTTCrI
2WnXdSaMrfBjtRbVi5eL85eftvfOpArZ0nYg/4xMWWvrkhrlWFgJWo/Bj7ygsnLX
GoDR18CajpMkl/3ysHeC1j2iP6/rJ+nd8vyOhPgsy02jMxdNLBN41mg/I8SqCUry
r1TslXDAnsUhqshBGbEJ0N0xI7LkQhd+trlzaW2Y9z+M4KNMZaRXIwA/pJiSWRLp
6jK4qjhFmbcS/bl+wNUVxYbmT8t+7IHqxWmLxMAjDPwk+VcDk4mWy4eiW5o5Dqd5
vQicLMgaIFFFYwC2rNi73rE2eTc+b/Sd5czNnwdYqh28dBURP+SU4A491t+KARPI
GAY2AVvVABk2YEnr+Eub8G1qHoWohkLj26uZpTs33za3S4DSfwIyFHr40SHgin/3
AwbxD57a98/uqjITyMkl7pu0Xc4yLrh2IUrnZgOjfxjAZ8zfL6E7m/OHe6M2U4Xa
9O7wQOxXQJPWr5lVXdLNMv7VKAV2CHGUW85nkulo9tl3zcAm083Vh6cZM5Z0p/DP
MnnA+aiI1E/8HTTz8EEkaYwWQyBOpL7HW3G4MWijuMv9bxve7a9Wi5A10DXYW+lC
tCqmjejB3NYxJh0+MQ2gZA==
`pragma protect end_protected
