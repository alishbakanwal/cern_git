// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:39 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PXrDRVc/3yRdSTFFem9kyieW1aruMFDWPGcFUESxSfazWw/gsgOPJEpXUOUHIXcn
8WdmFTtDoOhZDzikI6Ahzfz6Ex3inrWoaKThhCKsCRhiRKHXJd1cmMQrjytqoSJ1
a/3Xy0dCNdyAm3JEPDINii2JSgstrb5Jkb52Mo9jZHU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 23824)
BKyttsepciQE7dlRTUSeNnCfR+8dnsE8s1id2I7JtjVibv6xD1Ih5DFiy3xc6TG2
71qN7WVDsQaNIx1QruptIhazbVNfGC6yCj3Gd83MSyKXe2I96F5lL9VIBZMvw3uc
J6VjnD7pLdUeSHgq+97C62ejWu0cL/svogqJwUllUYP0o3X/Vgzh4+uDi80/bLgq
dCFNDowJ9bp6xOzwiapSCqQdq1+Y/z53F3jh8ApDvlejU78/uyAF7eJ33UI+mJnQ
NA+9hI+/GGCvpUk5YCMxWfo8bWkQ1XgCH/b0+5qlmuAh5JLhZdJ/XWUh1+VLx1SK
0sfa1sAx/pNg9dcGbfChnaq1jd74D5UB+VPpacppTHxo8mzkY4XCr6pH2AyYJ/6Q
58Ip9ISEx87lwndiFVFnIdzKgNIIhuV2LPZLcEF+oL849pqaBjS1ThmqKwfOLV0/
c+ZZEQ/tRD82vDwKacEawjUfJ/q3Xlg5iiTJrlxuvsjIP933l5rlxvdtuCk9nrvt
lniIZiBOhTe3vTFgS5JvZWjqkucfHb05TRt3hj20ZA4MZT/XPxEpTu9+OnzaJ+1z
AKyKmOD13E7gT+Oer+55iVtBBpgNWaTLCN1Nc4MalMvOjT7aKHlwRO9pS3Q8ecj/
2V1Dahlo8wQuszXnB+ueR3lgBkxOHEMAFJAIR+DhysTBrNzeWwPsAfXR5ARK3kA/
gZ5AIk36IyRiXVeXVctMUQe9GmqnlKtj+JyvrglG7jC1vGErpPxqrC6JwfkVrU7N
XjYDQOn2f8jOcbWhgZf08jC+qYlsTVs4kg5WZK/wvd55r/kr/R3KJpkipOG6h+ib
mdE+70Np1uQehrsO9emPYsaV+bOHqzbhOKTUk79cVUlAzK8NGadBk28AMLxVrHd3
xxNMmeIEvU1NEs7Z3vJW+ogcZGsDLUn6RORxCBx8y5INr2foNs930CQTJTExVe/y
6lJ3ciEzRRnOlcq875ZEgYinh08GSv2QvG28SFJO1NqmTpd2ezrnXDktjIh/aVTI
pATYlwVNiMtY4OdbfWSUAoZGizuBNmwkoD8hKOHOfUGSIOEZGKWrSk7YBNTA+cu5
d86PI/oxDkg/yCNi6VvnSBuJALG8SonrJUnISrix18q/zCz0ozM0XUTk8GdPMS2D
V7hxCLF4aCQdf57FCGBJ024yYoo4SZowv4Des98vbFm5+A5wXLHzccWqGu3VyX9h
EmBin0LOr7KlXRDkuSIXblExcMUwpFzjes4Atb0ndwqsOk9+rJ5JgE61dfsqJb8Q
VBMmH8G1riqObXnH1BZisdit5X5tUeKyY2Ey1MEHgl+K1Gl4n9h3W+fKQh4mKuqp
U1xW4cHOcMSI40zt8dwAe95+ffb/7OYwOVcoubOXbviMX6ah8aI6Si3zsSFhntdd
MSPJBMb874NtidXLpd7UwkJQAYr83kmW2z6ToYGRhwVsaim5ceefsGb0q/Ue3oND
Hr7gkrWFpV2npYwlSBInC5kfomrT2w1f+Ln8rJSJOjJ8zPqDK7CIa2PXWR/+pVfO
aKhYRnqTvcBco4i+IgsiQNtBTFud6vri5NtYLNvIpzOchgp8WGWvOxU0u3GwXq5Y
zNSp7IXMpO+Vb+Bdkcxu2NcTck4dFzkB16POL2bY7ImxUMCLXw4zPzoKOtyACd8i
zAoYHioeKOCbh00lmxgTGotl5z/kEmdCtaNqXC3SxQYiibraPLirS49gSNvI4Q17
EWcGWOJ6nDAy1tf8Zz7ZH0Te3HKnFfNPTOvzIN9jL8/u3AxKZjlA9JlBFZp6+qjX
1pmHKjFCDuGr/HtJ4sREXZDpENffOb6/NNMLpW6dkv/JMQCw/BVWEDg3QY5Ytdw9
rh6+mqCB4UW+wPnbvcu8H0EdXDFPNX+lHZYCAdCqjIVl3EbiME81+ADx8IM8WsBe
K7ZDAyHm9bkt4FlNyJJUsh/hCIFU4ova3xaq6fySzZd/5C4REioo+yV48ofIN80o
GpQRi0LexRDujhyDrZ44Rtm/D3XZtNH9URLmTac2KPZPUbYqh/43QDshj5j5Z1+D
gXkgNldrmvdIVMswE7FC2d3Pt2QD7FSfxyVSW3xaTvbdOYOU0DPe1+PQSzYPFr8z
W2pSEg5jhgRuAFj7WUN+kNdi82wShL9xmIxCtekdUCF5UoY9qVCgWtvQJriStg6E
s4CYKb63CkKtVNo7yzlohOKkqLRt9/HSze4pzHihzL3lI5SQmfksb9/KYF7dcCVl
2mEYngfrrDQKAkyvgyXBVG2KUjRckwRoWxdnVxNE0JDeAV7Rty8MEhjk5ADIKRnR
PUV99miMkCY69bCePIltk6UNH2FIIE1HMwZYXcfjykNC2s9wYnFG4NK3iJ6Iw8r0
2YTVn8VfRuGueeDBCon0/ITv56zKb6vcPh4Z1N4dms73agckD6LBJvuYmXPbO2/I
+AsYK+4CkKIzOmMwNYnbZ+bjxMk9XXTwg9C+N9Z3CpEdwP943iRB1jLV/oPKizrs
ZYhI6DOdFN5QHy4ITDJS6nUZWHt/X7s3QExQalFKA+TAzii0ncDvJv4QCfhJVVti
qyWtVXW2SGs934R1wunhLne2ENCzq3httjT00cdZ91eeyX9zUvQ9WUbtQ7olYYkU
6sRzxqyzftQ4ra773oCWj0jRIlOIgOQTJijPRDj5uFAOMO1Jv1w7vuAtf30Em5iq
vgPC//5cvqngGJrIC9ENCkzxBDTM9OJTq+lZvCIiXImdzLZUSvmwy3TfiN5j/bzN
BeMF1bVpcBy3MOL/iI5dvhq/zbF9dL6Ps1wEga/ulQ2mcOTVXKmz5gGg/ea9X5qu
S4znnKfEOIRsUDs4A5LbeBVc3V670pesmZMSbqAfu2znXohVmzwwcW+IwR8IBcPi
nTLzEuhqEfOMK5LJ42xwqsormUZrSyPOJXoFjquhbJ+1MvoaLa3OU2XDeOcSr2va
o75x68nRs9cSNFeK0GQ5Yhw9k2O/TgXlvBUWiXgSidfuX2guYLOUWt8RMjytipor
KzRNAO9PkVqb8HUKitwHoQ21+9J7Liv0L+FadMBe5jEDcWPXhk9c5/n3VSgPRnDo
E80orVXNcYeVY9S+7TyIxktPIdK3YEm/Dbjt/vFmgT4MAkChSWDcCCbQ5uCF03sb
zk67AZ3mNprF17zgMjmKs5+jS/ygKdfbYzOlRNMeyF0aHAotlCi46YP2holcn4mm
iL+s74x3aZjIbsbELO3Ikruvf1K7bHEsa5DZVrt24yxAnt5AXQO2/hMPRGolh9L/
b+hUnycbDOear/IelQdczQbdtnTIIaOpWep9tSBqmjCIyjh75OM1QHgNg/6q8Oax
1l65TtdodIAwfGEl2sNPz534AJynQKc2liLmSv6Lghr6JhA86sGki+vUEw/wKnYF
7Mi6+DZxRXwz0RRAM6h6RqmyurGSf3RKMErQHTF1ukWg7ITk0TqqUT8JgQg5ypWM
ivhnFGNmx8mgYb9W7jXGfh9W7lJMwrxl38+F6oaEbLDnaMpyWqZaZxywuBBETWLj
1cgqKfA1QD2I5hxCoWPOO84NyoZhAGb3jsmrpIwuuMXkNnIXgax9jlgAP2TTgk92
Q5LKiAbPLAASNf3XpG9sLS6GmzwsB2/xuWm5kHFtrvprADrLVzERSvEOvIetJbWZ
3JjdScBkbpeuFsWO9l57aZhX2NO1fQVAt6h2CV5UjF+WdAb4/ctqLNcWdWH2t81k
knkVyDqM5pRUIW91yellI5XyWtgmdtvtqv8gc7wL/n1/MNvAh61tD0sIMjN4wWUv
0E4i4hwEX1int9FMTjxQeVW0m6ajUkqan857xu+x9K4D+QWGhmUyUT3njHxCsf4J
ydGjjV87MJJO02fb3A7Gnwk368qux9AVp38XtA/wR3vE7czlzjwdclElVvxyDEUz
tGglHYHzrRAlacadu5Ixi0FfX71Ur1170yjl2u4aRRJmnvWEJTG5dccSxUkqf4gw
vcXnDR/kK8g0CruOuQxtm/jJv6B1/739VV/sX4Jvv8nfQeYrUQ9dPWfUPzA6wr+u
MAp/x4421zDfdUbLxi0owV93uOYozX4H7+GnljP4n+wT+XOWjsDPpTw+/I7OzM29
zD53LUhf3B/bPe6otQ+GbU5HMsqbmX8Z5d9zcdNurTsicYAW1Ylw1ipkbGpzFdkf
t2ktlEEcASljlw20VSdks/8LyQnGCrccsLCBtvNkUqwDYe4CDW5/BB3bAZWcqN0O
+hKkI5rPm9sq8tZwZKLU7eXwFPSZzQFCF4nQLWT7T+gUIMGD4rc3M3sGnnKbv7oC
YWWBEpQQJ62KanvQXZABM/FAU8JjtDavtxfR+zsNHBHZ3vCdmvm4FNdouNTobPk2
CmgP5FHxEKuBGA/ma4rtXlg4Ij+P2Q7LQulEXCN+fm/u0mYZGNXKNuRG2MkBH/xX
cgdcdOkNhzLsEyGYQgBJgUY976FWn57n3iRDndCDYG6Z2XZzJ+auVGkL19qLplOY
6yRBg7tDs4crOw6J72o2WOmxO2//fC5DLqTrhclPtFFL7UzzrcIruLM5AZoPGjTW
5I21QrtcSM3Fghoj5bYyTZY63fOaXC7M5jJFJQCEFY5JaPGwGGVYq2cS6wPRiWe7
oE3R28kUYDVGaojSVGGMcmi4njo/xRUPI78Z/to8l+QdhwWqsAVWWLlzPrjCvdST
pthMC+VVkAQiNnJswFYUhFxlfj6mQmzjKam8w+aDENZ/YmAwOwYgZrQ4ZvcDg5Rc
VL3d5vQZqFxX3kKuWg8kiIPrINV/6i5sDGchozqjElZ+uEpuxUp+zHRVgqk78NKO
Gcf9zx+d4SCdw9buKH8lLHcF18whdf2pSROJjkw1BiiSYI2lEaBH9MkehLEbvzJT
i66fEsEHLhpmgNrpjXgf3RKRqLlepxCKgwJZKdTtDCBZ9pS/sGWLYZgQs4NFg3rN
PwlOoF0Mc87uJGFg8AcccWjBURa0gNxO1M6FGEzPQngdSBGScBot62W8/UYeBisD
oDiT3vmeeTDYcVJx6JPevVt8jllaRzDCZsMx9bVC1fK7XMpriUA6CkTs62rGmHvu
6ad7j6XTukxfj9X4Q51DZvWKZE+yZTZgSf6kO39C5PrHnNAbvZ/9MeNUpjnTXVQR
/hWiegadUGZnQ619NKE0EfViAtQkbrIrETEgPke0Rk7TeN2UUvllmYUM7vmJ3LFK
5oYUsv3YM9IXzTg8r9cACfoBKOtCtKrR35B2IyskadrMLb/hxbobnTCoemddTI2P
5qKLPcPNAr+njwb2MvPCzpekhGYiw1t1z+tTZWFbWgwOXOtWgmdQ9ZqoilrxcL2h
rkbA9ebF7uNLthBm1K8dPkviEwIxW0muwDbqDX9ANka4ecNOKKY/6lIdCMlpWW1q
Mg6M2SJBfk6RmuyLvRGQABgysNPjEi4WAlXQsfcI+ndRFVzvNx0iHh+c9zp/V9I2
9VIPcZTa1lGHjaXYnFp5QD3xSbHwtZnNRESuxD8IS1MRitoWwZ5o0a9h0BGoR0TS
ghNArIbVq4Rf3Nmn95ArbXkALM39pfdAyXqn3OFDT+sEylMqvUq7bgCTnEyHOgyX
PhCMKVFKkHLTRXMbbYs13pwwgwhwwIxya8shlHjOjKtexgX2o5y59CiAgp0u+6Bl
/KiP//ZH47Zfj9/H3zsTSP9wNEEnyPiOn3+EbHZQREBBWsDQ7dpnO/is7ZNXwaAK
x0x2tTUD3bDcv6ZBY75Q9VldC5CPPXk4a3tVcr0arua+n7nB/paUpfs/06qhNZoF
2ieg2B7tjPx9RhHmOya4QEum5Mavg6fK8yfkNeqXMMezYXM/SC7RSTroLMLOf4XH
2B8CeQXWGRRP73fQCeGb23RzLsLxBDAnS32In3A8UMBFcMX4Z9sxIkbx0tC6VvHh
TwJH9fUFA/PBKJeTUwC8SeyKmdzURurqOymhS46vR4RYaiWHtH8KjsPOP7+mB71q
i7jvyplo1G++JsNPFvLURgvoTp49diR3PO3eun4J8WJEUcHPZj8ht5cOfMqzBwM5
XP7sMTZJx2EqSPPLHHIqSRfrhVGHZl8aj4gUutupn1yKs+5irpO3E1BkaIKkljqD
Qt/XzWv1CduYuh5Lb9Ht3Ck9EqTFlV+hXP2KoZHVbbqZBcd6sV2AjyC1ZtRdMF7o
8O7mpbn2tCQUFsXFMLavA6qUa2iFdnsEVV336pgFqYeOWHlXTwN7FxB2j3zuegbp
7lQ0sX61NG1qcGQKaUuNhuqroZTJ2vWNHgpPj0nk5DA/MBua3RsOLdnecgQ8WXPW
knYyCR5fykeKA70hprrOhrDfMnkkYrNkkmWtZc5f2oGvoYDmT5bEnAXwz7NjRJ3B
7GHs8zriI0+ny+1Wof3WbZDHcAjQZWhCHmV/LeyFUiWwhdlhOT0Z5JHikLAjHmpJ
DnahRJYIxcnyxT4sNuNuR0yvEo17/WUXm0pUczFvQ08fKDyh9Sq+E7rwWuZVfd8j
omZGhsQFzALiLB9eMXWzufREKbacH5fyTdsZ80GimsorxUmDh4vhtokcTfOsRHGE
5wiTD18IXutIsCA3HzYWkBgJCGT2AEoRUIDWsNsLfxjRr65yYmZutuIRYyqpaVCN
7coy2whEunJ/nUlY17M2GWzFRFr8KH0rEXhxDJCdK+B5HBP4UQYMaLvHxVBeDhR/
X4/92TSmPlR8Xegfx+2PbfWcr41qgaUI0ki13PWT0GmQXjtjGiB38P5wNWg1bnQR
6PlXnlcjOro8n1PBMB7+DTmS3TiVJHUZYXXz6locaQt75hGgU5ejGELY76B5484e
0ef9L2BD4WHwZWc0GOBDhkngfASWrvYE5qd0CU6g9Do2ia1kwhehHdCdCo8IjMn3
cyU5oSZ5iRaGJwGwbTPPu3yxO2I+yIwpB47Nxsqffzn/jPP093+Ut+OMmNJYpJ8n
xljZJf5Z+M6sBTQG4CVK1S0V2k2m6ghDZZU7D8CLkmzjY59WfGUPyWjNEEzc+xvE
1K4EwHUYd7DJqx0Lims/bKiqlemD+hhuZcZ2oQEdqryvmQb2FI08OEEjwS6L2Nyh
+9cKVYrN6opRLXS8ZfqZhoT2/gP5On1psDsEXGq80JPLa+NP8zXJ5XyzLOEBbZUW
TLUfEpGBTtDpNFb1Z7yLi4stnw3P9gAIK4UPHOkoJMo2qksAnK9WHQpcBwKxQa2g
kTL11EtBdayvu8Nea1Lzf2XeXdku0cSK6isHi6V2X1mKBiNCY/6ceEVJ55JJ3DBX
u/tp5H6Bgju6SCtDJ7eDjG0/BnH6fte5ZGlKeDoKpJKNb6v/2iIculTwoR8eXIec
ghAINBhCmmPgpa1DhF1K5xodCveL6XaX2fhYcnew9l7YwMPAXC+Fox5l7AOIbQz7
HVPYsfjDQoomslPF5UzM6mTOr98aJvOdZc/QXjudTECXfKSrjrGXq4OG0tOC2DfD
GBKllA4aD5jhVy265G7rKAwfwS+fkBOYHLSEkZjtbpywB8AMmQkmCfscOEU8g7WL
EHj6BnrQSKcQxV6jRPx+Mfx8n34D7wBqiUli7cA/HHaBqv4NOa3UpxXUJK11gQ2Q
y7aeCJw6XSIVV9aLX1Os8lTOW1E9rXzjjwBoj494nl5pg+RWmfPWb16fvQs2AubW
6+LsHobQGK7poFMr3B4RQ259JOWeCcsHBFl3AzrNjziyiqUrph9pAFvypuRJhc00
cojaiFKW2fV2yY5LUzxiYBcenYFpKvYQiBx7f2/3YPy0Q1DPbHncICRZGNzRjtyj
ZS/j7RPwBS3KtNGIGmSCp0ANAbYFLL4553YSQDDLmQs+EVNjoIEV0ku9siby3N01
5jnFCo31b7iECbtNGGquiuSaCeIAg+LZovyGVmVafmGArTm61NjmcNf71f/gi20s
G9NCu3hL9LIxi2qbheOGc9PwqEP1/ls72lEEBv9cxaxr2pFIR34tJ28Ffcwd8Vvc
2Xf3JMCZ2Bvnw768SIUTgNRTaxa6tVxn1ACGk3PpMV06XdE341U06BcuxfsBgh7z
KO29bxRBwvrTJo1aqTDMbKO5k3BalQ0mDDfJI66k2K5Rf4usTUReURqB+DXY+CKO
+ulRLN9Pe2aoKRqwyBz/WZcmUaIg4IOlGTsVwdY9d9T/3/faCfyhPOqlDfN7OETS
fN2p/jCdhzk0f4en3BvnU0jEpxDhHT8EfqrManaW9gAMMKrAETzJx/HlhJkfImHg
5tparbLjbWqTqJAaZrpHoZ13YDLCNWGzQUgjHDXhMHEfuZC05x2el/X4VRCCJjj6
fxsxeQ0Ok/6w4js/0jXwjN+lAsqsNjv4hR83kJ5yqIYQIa+awjXrijwatkDF6bcc
Tn1c5VzEIJdp8attDEQzhIAmGTapWxVavHJIx//JADKTV/jLM/D2zTXNo4iICg65
WwIQtuBCq0IwmptzsX8NnWxlbirXVCIXeZxIzvDNVW2M6wqrPLF9WmO7y/w+LiBo
6JfMA75jvFsQYjhyjdc8ZSvONOJxFM+ohkNeh2K3L5hRjDvsndfKnPAb2joLwWpP
lBMRdnF4L3J01kh4BRcMj0iGOZ1Cg78idAOULqQHBNt1yfp4W03olyxjouwuvkhN
fCGSh42d75m7sBHfs8sr8OPVNm/x5qPFSH3dklsjyYGC+HH/sPWwxzjVnkmo+kYe
BQTWYLtJC0on1Z8RqErErk9kawEAGEOFU+4pVImMVMGBmureVf+pYUy6rOEyqjkX
H0D6weTvvJbZUq6IrGya7EKf2iRQ4M1iwx8TV+COiWAtcRJqstF+oCwpZfbkEI5m
gK8ggubgmcPENjWl1Dd3Fnp+8PlTL4f+WYXEr/zBgujLnHK/1DX12Cs3TNW1W7U2
YQZFJsNmJRwQCNw2ZhGipUItx89Nx3MA5zfEw+gvGWLUFq1VGaOd5f7opWQCaq41
2buKNqmFpXmE5GuKUBy47tNYJtaSv+g3NU4XYpxCWtWOP2O6WSH597HZCRGPMT1X
K0Ua/h6FeHx8lYUTo12jRxsThckR0ms4NQUbaIldGVTVxoxY46lLiJKMPKZbXL3m
FMAhm48+yza31i7Qb1vLRHuk5b0BjLdiz/074u0cbSLmIEKIoeENTfxMSkTBMOmA
zgBxEqelO56xT5JioCLAC6ZhZRYYL1bAzu51KI0NMWMrPFqim7P17xM5OVD9YmHb
iqCSPa6Av/ke83TKnrMIKqIKoFKXfgiHMZHSpmmHbp5fT7gnbWzGaLiajYoOltBA
8jNX2pmSI2ktiSspJNELrIZ6+bvwDWsIQ8IMOOM6PK540Hxk0XuFjoZUQvbNUA6H
IWeDUzimDQWyAhqEPV+V40RbUf7RRbGD4r5dUIPr92oWGcMcwrwSGEWK75sksosf
kAKNKAjbq+o9m36fbIMH3fDMswn/vAVMxy6Cyv/0AgHno/di/zmBoDMbr23R3/KJ
BCDX0nWLTowMiOYSYwkhAsGtW8Gw9N9niRHbZTlmSV6/BnhIJB3oYzwH0W0Y/Dbm
aWBGApkg51emuZ8xD3HTWmUuQwy9KsSi5wybXPblxqsWY4f7TSTBHH3C+5tkM9KQ
XcnLdnGgBtX5POb0TXxsNHa80fZTUPuATuh4aKSE7FcWRN780FTlgZ02Y/lhTA/S
jvgvyKLTO294NGpH1Oogy1KSRx/QLNXwL7e5JyfxqFQcsTniYpvsfDTtD6989vG6
tV9OM0UhWbY8Gyzv+IhzzULGUBR+u1c6AEeaS6NRq7Uw0Y1xMTLcK3Zxa739b8y5
atZF/6XYWtZWhsjEJafzVdM8zdBcPhibYS8XBgu7gMqwjmlpKQx+YlGBynQM+ZO4
ZiXh3uwnv2IZbSEH4JGG4dMjoa+1i2j5DQuFfS0g7MZfrxOve+JLwSsKRlqegyNy
AZ7o0XBQzb0g75Dp+e2jHd8kdCSoHr7p1spc9WH7ad56IK7KnqqiPJxGXOdpObXE
0CPHIMVExL/HMIFMunSmrLzOHiftFxurDh1DcFHvTQapGnMf4uslITEUqpOmW2zl
3cBb5JNoiYIxE2f4CX8rYlvBdPrBTkKvAhBOvckHbNCiXX9oTOCCEfibALXnD+aa
ih5pNxeIo6Dd+LbsnS2X3bO52gi3HBIS8xaCCpioy5U809kjc00k9v8vNEZwGfd5
TxMRl5TEPGY2BF+8NvRRKuAGFORJeavnMrl0d7XUNK/YxvvfqUiZneDM2agDLbIw
mK1T1bP2o7jTUQ+vjZvv5d1rhIcLNyQvb5jiuqTRVvAl8G8TOct7YMqw+Io2wQEv
xbD3M6Z1pouvalSFDKjswuMjPyybYM3ECsd466WGsOXiCyGgBwB3RDVV6/FaULaR
eBSR4dIleuljCE7dV1lwmq4rpgauw684QqJb7wO5IHPGbK3ujr5y/ThtRlv9VNUl
cIcdhdnOtewHjYCRJIYPMeOQOJirWH8d0G+YwNZj5pESMJ3MIfa0XuORk4Cx0VQI
K+q5S/czoib50K0xVX24KMoMG10g7jFYwVZy236lTuuOU2vGtqzkvJGWYMMPwOKc
d1ZR3ghnNXKfIDFcDMPMFNUo+XHlaeuQEXfwEirhTonPaE1q6nykMU7GEM1HP/LT
fjwLudT+IPiVxHj0caH1ekTf9WSePdPCbaN6xEIHPxW4EuoECxIyjC/B4UZQlzqb
WTK16DcssURnPfIDneUW5PQxOED35W3p+qNiLpTTOopbskq2gBzE07EWpI4W6Itx
4ZzDL3+ErHMdmm24PYHrSWaLxo5PKMS34IU7tY6yXuavbzDN4I5ySAiFF9utalt5
j8UXmWJ15xucjN+pREFBCxuG7nYz5OCXoY5AFmA97cjSF/JMf514jncpKCq1KI3k
3SKimPb1SxzwUHWcnny9a23hWdb/JJqlFysM3Jd30splasTVlEn9/WVW+VeuRomN
7g/UXFiyvmThX9RbeUPZ5j1oL0B3EiAb4qjCc+mokz7SHJOHyxY/YiyP35Q7+cuO
dHo5jQb/jI03lqZh0ixfCWmQlllJeEIOvzRMAt7jJGOzGaEnXZuyJtmHBJRHspGh
cSeLdSMAoSOHgwuXuRuAhyo2S8XUYjU3VJXqx1i+o7iZMM/1XWV42v7Zvj/vr8Tq
ch6tE3bSgb+xYA14y0VyH+l34+j25BMK/vkT0bXCvC4tzfJy6GVfPWGWMaQX22xZ
LBSMWq2A7pIZxT6SXYLc7CJeCz975vDeNcSwj68O9yRBYJSwz2LCb3wipqlPRTFL
lzvfj3q6EOkCm0NxAzC+ZDQJqJIb34voQcB86bf1wfU35RJvCCrAQDpVVDoiXP6V
P/llHvt9nyWLWIKvio+oifgVQmZXI7piExZ2ZD6+FrdN2XvJwhgY+nLqtHokL2Hz
F0tzCtBH1FFSqFfbWVcjzHzahC8rEbvTCYphWFJ0kLhECwxalIYYepK9FNN03UMl
ReFWpVQPHw8wkLJl68xOv94vTf2XL4Dsu6PXEcLzQmf2w7bBksNy2HBVnGgosxaw
Y+IKcbXugm38Lrj+I8AqEvPP4dCHn9Wsbmm2W2jO/1siz6g04UfBNoFy9GrtaaS+
U60Ft+U9QpGg9iEg3Dlrn37bIH3JQ9y0aiKOI+OslHEfSBqn69xn9BF6ZoRJ9/cb
U36UlKUkYyG32P/gxf076d5YKMCIH+6+9VoJVr0zq7+U20y16g1v3Ezx1h0Gc15i
wzLcv5AS3rKfFyEk7Ie77NMDEp8YCdY4JlC9+ak28bSKCGFIyMLpXnWTRpt6oWmB
xIaz34PBP3cTepKfRiV48kgY7fthtM2sxnAhVMGpQiAHmlSAgtDNaxNd51SSMW38
bmvOfg8NScorEismf1QULIa8UvFiq4V0JFLYvZ4FSY3qRmY0ELnfpTrVeX5ANJWB
00GMlU33A199CZFgOx1HySvDEe0K/wP31peZNev4Pty5ugoCmAm3i+8pC3ZufPif
uClPmiRXtFDd0oibTHO9EBHKzwxvek+btuWU6dGXZ+icZweDeD7HiFG6352aImnY
1dZe+TatF/yQMIuJrzKO11K2z4CSyRWW2tvQwytWk5C84/b1qap3zeRY+ngHnygB
1UL/KUXyZ0Mb/zRxoO8ab3nmGPsYrKg0CbfPRNPM97eS9fZeGP0Dua2rJnZm+1lF
KLp4Yu4PdALzauyYUqMu/ThYhMpkSrqMuEFBEx24qCTU4qZC/IfiDom2+LNe5rnY
BNtvynheM7c5dt5r/3W5CeNMqdItzspZVbIHlMJEfE69jpJK8M6yJcss+OitwA1p
AHSeFVKt+w25jy3kkttJPJGLAx3jL7/7+8+wpEL7dC3yLzno7HH4ksPn1zRk21Fb
cDjUEH7DSg85jCiaxLPJCdOL7CvVhmKktP57g9ofM2riVFhaW+bf1XecCS/lwXQa
I5o4+fdAhI3RPEaRzxlgFXatntgT2YcSU79nQtEaOrPyRF+UgKMobZvy/5Ad/n8j
1YcHK9taJDJSX0fFT9a7JP5itp9AAy6Q6jgwEfby5bf0n/e1iCbADTwtD8se4Xqj
Hue3gr4yUZdrf4KMVhfBCZ1OBQ1FF3KcKWXchJ3aUQSKYZ+px7UAgiVxfoNqbwYn
mcE2UAVcziqBaPcYyQYO68fKD5Ttr8a4iLVY+o/dUd0C43fhRAvtB0c4QNLWBO54
pmqyuWbw8yDBRgKxmsBO+aLJdbHTfqx4PIvT91w4RPr8V8B1RRNh+S14vE0AvkPa
ISTJRgUpUcZUQt+dwFv4YL71fVyXgfDnYMLj3YzHN7alEPWkCybyH7XRuDgcnmy4
QWoTplCP9Y6cQskjyJRnE8jngYRLSufnfpBFbemYMB2vITgrQb4IibSVxHyd//a0
NIWQzIQ3xNZRxv1ZCIugG0UU87o2uOwlP/aXPDKcIQJZB72jbT5E8+p0XLCvD9jj
fdSJv2UE+Dzt4bf0ODboHUSyvoD3jfIMF8c1sEJTZiIZz6ynHFxAJTqNBlrK95AH
lUW+uNQYB1uX0D44x+v1zIjXgcMJEfWqHpKwVt9Vmg1FQ/fZwSevdo+pDCXDsnqP
w5i3/NQ6cvfQUJHlCI1rsexnzeFFTICEROCRiYkZCFjWOSXqpEg8XhkO8A1yGx1Z
NcWLLe6sfE2/MEOMzRTFK0oin/4u+9tiT435nH2ypKiEElqC0V+QpgEA0gS6pxrE
ba3fZWkAC3BL+HHjwc8kLMiK3HpPx6GgprkyT13ABHUlJlJQ4KFICi9VbWx4bXW0
uG7E1rPo0bwLnNvywHfq4qf8VNo8gmI+J0O3SXU25tTTMIbszyQnGPX9hhPX4Fpb
605iCiuEygRPhdH9Tw1o0Cf8vPOn8Zc+LfJq/oYezXXDb42HF9CEIV8QJuyzXIKP
BEg8iGMmJJUEXKgYOz4TT03WZJcRdnaJzc9S+17E3vdH6HVP/G5gsVqBT9cR3lA8
/7Cx0Tb8BTrhUsR08ZwzVeoZF/M7G+NhGxUHThn/3ZXqjYFKEORSFJ8WmqI78AJA
yEYipEI23p7jFqazYKMlLbE3Lu0zUed7TFMM/+DRLUvB0FBf4TmRKx4RbQ5hUo1Q
3VVIx39PUEHf6Jlo0cfbU9Zgmk8oIHYqFVluyZFKhvbbDSCwnpuEzF5eR0mzfzLV
cx8vixL0xqaZZLX/mbYkR8/PEkZMIlnKCB0He2zCQ4cV8xfya9ud8Ml0nsq8agbv
kgXVwJl+uonDTh/JKY6+QknQoor6q5H8QBir3b3xx8LaBzQP2A00gg1vn+N2BLZw
zM+EqGvzZTMvNfBinqw4tmZicmAyAuCxu+55gqxAzddcZOijdaUU25N9L/Sr5pT/
CYYu0WKc1w/RVXNuhhmGybtHXi8VDv09H1haL95Yoveuc/bOxzIdjh2Pm6YsPkwc
eK6V1W+miT/huS6g4tcm7Bnag5t95tET0s9Rd4hWrzB17X+fIDGCrCW5srQ3L7nH
gjn+/KMmOpIK4TKdLildTuoWuFqvhws2dFHRUDYZclNcJKg6x7Gqg4M+ZEiXDB6c
+5kN08yc1AFy2ftFRP/bJwLfbmGfZAKK3vCqPy3A3RiHVYdbBw9jkRhnZv77Zwv9
HlqBLxYKTFe3O3n9aZ1ER6ivSPhCxsDx7ExozFccswJAIrF6zxGF/11B1o7cYczn
Lb4k2gcA9xRKfr0HdZsLEhlzGvlepoIkfuxwheUUYFCjtrnlNEOeiGv/8JfhFjFY
WYcd2pbmn+igS1lfgH1vPfJJTtNzAV/B6kwOJQW1EvNRZd9qkmrkSM0xqo1BBJ9m
wiDWOALX+OkZNT9N+GJy58kIUiZwV24PZK0qNy0Pdtbqn5oLEPL6RKTp5s7slv5U
l916dskriLoPMv83569+zBabOVSzNoMV8+LTlD4Ddx1HqcG0Dn8pEsIkhqxnLCem
r2xnKW8c8zlxpWRb6FPzX0EY4OiJPpeMmNxzcS9Mf2BX4mpHloISqdIoZ9cakQ2L
BCjgMJ+hMWRzu/qwWT9amy+tzEjaR/qTlJRdVs39Hpmi9i4sz5WY3NSxjAPh6aMy
8SxrlncuslYaK14DPrZ2+Vq21GIjjq0A9/2NCKkvL/tz/JnKvAx2bXG4IhNCPbkk
H6ce2RKf1UnlAf6mLwiGBOI5XBZ51oLYQfYM3LvtvrMhfuHtNFce9RQPrkR2jb96
bmDp6qEUa3c91P5YkCcifcegz30RiJ/EsgG8fLxlHn9jdztI9knnRhC/24GHDxI8
SQV1stQyUnzU3345b/WI0allAwuee0hRFz1z0iu76BOXJ2qkq11Du5Y0Cf/wSGPN
l9ZVIH7sliQTSfpTF7pC6lHZ2Ll4z30onJHDHo6Ovt46y78poUMu4A+hj98gnUBd
jqJqxcyTDhK0+XS/yA3EA9RuSJW+CtxDUF5fF6Rae+jAL/buFq8O7z0aVMyM4IZ+
AsK7yA0vyRnjRbmd+1oZ8PBgfKbeKB8/U6bRs4C9l8sWBulIS7Kpad3jyvIQD8d6
8vBYfv3/yd0TmdMB2Pb5WNtNeJZPAyTayQUpA7tnLYUxvYq9PwJhyMU7rijACK9u
24PX9yev/CJSOef26qGOJqqCANZKEwEFFyv/6tMAU30hezCofmnp+S00W8+6ARFv
qlbQER+If6XgSAIg3wCQV7g+MJeBP61Ytq5JpbKgFCrmdG/SbfGX5WwrnUhXwnzg
3KlYuoPMjvC9lt23SGwGi8SdWSxWafJgYu6F6RUFVztx91j1uJC0RQAPXuymTEXq
TDhRIHA0JprLJjkWNnEX/rcGcRgHsG6qvuVIaJ3jsvr2sZZb0m8DpME+mGrLR3NV
kqbl/I7e1XBiGNkwPS0Z0iFoTuL948Ew6ZoVEh306RvzsDH64A7Y9/khd9BKKIJX
L48VFGCYUKSlrN2GNS3BP7jehvxIInefaxux6pMdwmsVUPQW64bq9qypS//wWYld
3T3H/o9uOWJvAyeHjNAGIEyGC6CT9s9RjhJ3k1e5+CGyWfpL4a8f1tCthzihswZ3
Ea1ESmm7zfZksZPAYznf3snM3Qm6ZrkuPJ/jbN4W8nekTHRHXGHb0wSlgx3ATD0y
2FEMqj6a3m3N6O9/LaQXPAngK9oseJKmW8vl1HZeAvMAl8XNOEX+zvIrdu2gHhuV
noQwhd1vaW5KuknvNxhZz+eo6A+UJAUEiM8UoSeiJ3oB59cLu0SK6XhO2nBOTpR1
pnk0Pz99NLsxWF0qAkayp2bFjjJnflF6NW9cAkguKVBUKpiR2jiGO/RYV2zqpl7A
9fQEoiMMa2B2lVJq0lYvcf3lhl5VntPnUst3tJyAjuNPPPqhoNykSFWoe6XAkac2
8ixUFjz6fshqoKIl7viTKJzC4j0pD84vLeTRckUNutzdsdZ9IP70WvggAshaoWBl
OXPNKuJgOX1uJRCmWLiolx2/c118HXF2dpDTmOQHTKWQcdrmTFnIWw68fu/FgeGH
dp7psZ4La2cPVGTcTU/5BWQ7PuQwcieYI7qNJw1OsGIRCOjo8NbNoHYslJcZm/qt
SpPPF1GFNjHYd8MBsjmq1axg6gh2Iwb21EmaqWBRewrndA95aKbfYsNzX70WsyyP
NyGoAymz0jdYMKZRxna1mAXD4v95thuqwoYSiVLs7eBY9HFxI8BI5ULLNVWixepM
S2ucmq4nJaHgMApAI77s0Hv5ub0LUa+4Vgy6gHuC6ub1CJhdA66w9bsenxpoVoxq
hRevwQgS8Pt3PsD55X70M9wIHLLRWIxPep3IHvzgHjicppf0oWy72wiziuAq7yOo
yjrpVTmy7ZhobeuUR+qFJSgc8YnZwDWDF+hHucjoVK9WrmyH6TULZFWoAeIdOiGW
BTOhCSmQ2cyfWRndQQt3uEuMMKXD3OXqUMuPTs/zO0/y2WhgYOV3jeNLM+/p8dq3
GM+XQleIc3bXed8xsCDfkalvau07pqv3DU2zXl9V1suZ5/Qb7IswCg+VW0RGIVj3
glrLwEAvFhUCWYpFHnwPplKCWty4jvQJWfgSPHvY5Z92U0paVT05n1Lcf8ZjoySW
29CaKMpg1iXr/y1k7+fl+DSuOlsjb2qe3J9f5fgJ0tWua/TPqtHNzRiLDa1tJsDx
fP7dUe/3BepW/2c5Gka/aEcvcm4h+tR8MaWD6q4LLQuADEWE7VIEVsg7onfQGnkm
uwUfALwYi4cNWkhf5MLx5aDtU7e8fL4tWFPCcm1SOppHaMol83H15qt7KNe9X2Jb
jgNlKoOMRsvu0t6CzL3dZEk8vpD5cY+WFXpq1+bAF0GMgw2zWsTyEurZKB/mQEAx
QqYPUx5OgO8tRbzGzQ8JQ0OjaocgRYlpQgxySiXRQRYCySMII8k0+qiohEciOf4r
5EjuJ8RmZ3de+CONSjX0RiXnGdidXAD0sdUGwhPm+KNAhfvq8/KjNNZ3CHOut1lx
sxo+SYyZbjEulNa1e+y69EyxhU/TK8ZHXADwzrCvfnKiu31v84xMDqQzfKCOc9Tv
Kbj9APg4m82VXCdpMPBd2VqpXRA9gZvMu/frhUTW4b2CplvVDSAuUYW/aYSsXwqO
oyOHV5L2aHVtlBk9xtfyt2SbDNEVctTiwevZItdMGjyIkTjFW+aae22X/nxNS6gK
5vj2OHIcorVY+fECFfBADXC1vFKHTH6pP1aND0kdfH/9alK4mrssl2DoX7pQt/sC
c1lWlwoBx7yClSD3YvDEmg4GC3jgRubIGpyHOOqkYigJv1YhABnGFjPhWyLyZGbm
JbTSGrj9bv9aFhO+h72NvXmfIJHeAR1V5hurXvX/ZVHpzt7/0c6AEwebdyABsu4W
pQtQ7Kk+nftjIWk6altkcizulrS0BrHCBLsE4xmFteHoBBv4ONFQMKdqluEbmHjr
RDAJz46K+TgdOc+AfbyLezBmJoJEJIAt7OGsh5Qq2qhp4fykL7J0gMv9VhCBouJT
Fk6s9/ahIwkgOvFLjVPPr1A0DbeIQD9YDFksFrISuY6RZM3XiIV57aXheA3yOEOe
oTWsl+jFwHy3lR8JLDwNb2bigGpNXKhJpMN+h95qt7TelwWlQb6PMFrh7rwAH4IZ
UfqfwS2aBRKGdAC3sYRRM9z5zSvCI4oz9une+v+Xph8bim01xQMu5gVWiMNDAdXa
0qXNWwJ2GPQuu8HeUCNuyCQZiWt5wCNrWNytqe+ZsntyNK7tHUWaUMdD7REyZIPS
PMV0kP6twCyHf3Vm93DmIWcIjCCUBFWrjBNosQ9RUM68ihBAoZw+pkVXLFB8Go0z
zQlUFPCv1n8A5X52TRsYESVOGYPo1xLaPpnQ3tzjCRtrm2kVD02K4+1AJjo+9DWO
EL0PnoiXO50HS8O0BvItbJDSnPGlVg9LfjdVTQzlDVqrPcf34qb8jZnkxNKxVZDR
jKFmZ2iZcJzkrOBDrrw32L3i3Yupq1G51OBcWflmfD9kkOeqy/2FAN8fViVbEVhG
w0jqTIAW1LB1+ELxDgLGq7zKP7QNefPTRrlgDiYqqjYM8SuvzrFNE+ufXHuCuer3
EGWSiBgnFopSlA66aNk+Wd4FmrwDV1qBSIafu8+acPn4YeNVFO2A8lCqppWYU50v
ByUeNefMf1sb7bjg5bydswAWhx33KaNmYkm2neTRRtuTJcCsIkMY6E1w6JH4+mmo
E3LCLVDhDoao/c9izSi7yy5xRQ097i8xVY8RGAdKSzFLxI2gvK1a6Wzy7OFvdPdR
u0im6etXcetUCDGEvWvLo2ztdjj5GqBsvHhi6b3F8UJ1pO7ljav9gJUemgIAGJZf
sP7QDbSGDGjdJNjjmrZYvkoylO8EWDAKOOE/jny1ZAm/KIPXX4qVE0zaK5p2lcw5
izoxGEM54rZcmRtjvpTZtP7tUoXGCuneYxnsUgO7mI5cSHw3Ro+OFVRrjIkaQ2q7
J2gbeoIMkXwMrxjc1DCQ678llc1g+l3HQxY65tZ6vQrIJxjB4xbK/2DkLlCfMMtB
lEJT5HFiw8YVXpa9qPIRtE/EXU5k5UE4xVwQueDLzNPgBqarV2ShoRhMGVeuoI1y
CBQbRwG0AqiJiMR5DikDy8yVTtoFW3PwIbMsYtU0xS5rii8CEmJ+B+AJExC3y7be
BptfbHsYYk5kXdgUEb5qlVrB1A3x2LOSs8a45dh+MmwGIWQtDmyCPhfk9kpBwHOs
xj4L8pgSbNOTvcAY0W3GjHuUNfObenz5qcgBLwmCjkIhzzKU0QLTrWP+HKdxksOU
hAVUcXAbaStQfsYMM2fr2/I4NnXVq2I3ZKYUoTC0poOaI8Y/jt1iGnWSgh9TgHsj
H60sZ/xOi3fmqIdnLIPoWP5DFVd5o8oQpWIMw19+D/bxJ5FI8IM1BfoGRDBbcRfH
qcfJppw7aKL374b6fCo8dbmkDrtnnXHl0So8LwVxZca5MSGmAYFUUdOu9xiyrWn6
AJkePVY23HOZIq/QYCogtCGYuruhsUVijy0FYXXwSMMa132NxT82ZPugTegWcsbM
yacBB8oX8ow59hLfYAzqHV8CM6e8l8ZtqB4hf4DiVSxOUoNNI/FzdOCJAvpkp+b4
2x5uqqh8AZGgdTKV1dQmASa0yrbrxTmkCrVVWIu9+cDL+b+LvjQlGN/x6t24D+2Z
LXl7oyE9BrT38TOI3qyjy0m+KaQS73jkFoagZdVo23prBPGIT6GNrRMb6Nmdbp+v
Hx60XEkALurfyd0oRrtm12UGkI6UcLejggJZiU68vEfn+SgZjXM/7I/y3XszUr3m
izK6Ih4wbeePCTPEk0PlIRtwQGicjte3zSJ2qB4h+LryZrvcZzz/FGFwG0Iso62T
uipJzShd5yJBPZd+BPvTQQz8pYYJ8qzcLhsEV/yW86wZ39AsLbRN5HiWYy6SmAlq
rL8KwyzyKXRPttzQfFgjRk0lR/1A4/quPblEeSHWXNU/bfg8j5EM2CZmSiet2pwk
lvnIMFNSBB4ywJY4rXVZyzaHrZajGMhMNkp7mCagaXE12T/2RoY/UFHlIM/NBe7W
9ub3S9JtlIuJD3GDiI7bg2jx6fMN8Hco8H+TMranP9U25N9n0k6pQe0/sR7Nyidd
eMhmAyjDwHlvW83z/Xw+RIPxuPxVVljV67Le6vAdQac1v0w2uzjzI9TSW27ILiQt
StRPq3stACLmOYRWNM9dc3LiOYyvAqYAAuWB3b9M1J7SFVfuK/RVFI7xscBtVMfq
KeEGImP6E9TfAQ6OGO3NRyCXPxNEX5H5RtC6rD3Gu1e9R5LkMXDUih9iaoDSp+Fo
XsOmqPL4ghflMqQzHRpdrmgivTwMkUQDkWE37cCxs78rzA1GzfinsJMl1pxgBOji
u7QzI9FSVKVc07tr+Q7lEofxiYO5SlSSBd3qAHmJOTD41acA59cFXCTuXBi9lEtl
QySuYu2mSnu/jWzsE3TW1KOdr0aNbBcc9PZFpNGj38xGu2K2mgh9YQTPfrbMj/OB
5haLQkN5SrbHoS4ItdFc2NSQCuyRfZQWbEr30bQzYRalTd6AUzYhragnNNZogefU
jwi3yuS37maClneubvDdspMpz7I3ooo6WFc++1LV9v1YxY2ABAetGPrU66QtyDWu
r9NGCzfQ8CgSJqkHnU8NS82XsZysW6F6IzOBp1uKZqEnaPVgfrHJsue2sFa2ZDDX
NOFG43GP/xwwRKdbAdYmW/K81dPhspyGTQJmCm5jf0paLNIypWQwj4aajI+/kQAM
vO7cdsaVCurIacygirS3uSMv5VWE/EkMUqH2G2olHml0vaBcLYFiSg6T0jKLpa8Q
Op66/eaW50UQTjo11ZAOy1r7TZEFZlAZIoWlCHsycKghnECIoGTtfXdZReRS1Tsy
bOqIQ2Txd47htCGQHuO3Ep26hCv9FjoVeUzhBaivyjFLmntum5CSuT1XlycHrqcq
lSv5RjDhzoYveqNZs6KUi6cL8BIh5qpkibS+bmcvaHhNLXexNmHcsaktr77fre69
2TBWLbYTXbiDByTMPP0SibDYrKy2O9XeuDO37bPG2nPXaROhwsE5Hxdenvkohcoj
lpJYaxw6cuHsqmPZoci5GP8n1Pz+jJdCHJgLt37J1wZV3cOIrtrIZKHLhW3AjOCW
clTCscznWjktDZBk+JAaHynOlQzuIuzzlz56CMiVwGyIkEeYEdAFcIayo5t9Ie62
fTwTR5I00jxFVGhj8FejpVapBp+e/97Jy4Xozxcw5FMnwndBQLbIUw5Gs17iDj7/
10PAyapMo6NsudgPi8Hfp/zRpGLn3hgS9mv6ZMvOJEKOoTGzP8SQK3G0BtkSVvJ+
194ts4Dh/dK6M0PhzLe8oM/bYRjCSIab4THgLWdGHGmh9XU2cgqSA91CV99WU7eC
Q1l5b+hLkRP/OkwmoP/EB7lndduyzgOHLRmsro+WR56zsjptTxKuCDvV6S6aMu2F
ZOrImM82/Ln/2oCZ+pkHSvB3xziHOAFTSUIEV62tssbCcSrVs1AER05iVmAVnpt1
rsbCBKujj6/SL9HRPlvq4qxixH0o8ILuqWeWbK4eCT1I5e+I0NNrrV2/B65KGQR2
uGKQL1fgmIF8Oy+YwLLyoJwBMsbkgl4Q8NRfS0lWwr0H20yqjp6w3k4kplBPNFC5
pU7ZV6HtZREju9ZsEowz09zTMX4iEGy/+Lb/g0PZS+DL+KZ1F6oWd4weNm7nGg50
seBG2P2JooepPEFUhugEjfMONkTLfi9cz35ARXiGLPhDpue0xM1zr2SExILYOr+0
MVDIp7xDtNFfR0NvC37xhHEGKKMTPDvHAOqhMFi96QuU/gI9JIYHAX8gSwPFU0HM
ncZqSjiIgeU4HSozOQAxNxZr5RmXAg/nwJEKZtf/EB7ZdJy+VjJCi9D2c6EJEEWb
hHqgy31kHZaqlIIDpVlEhyNd4OOBoDWgBLiQfERjMihmAY29pUTe9yDpOEnEw3MM
nnGEXw2itiu5GrDCqwmicAyQ+PMMZ1oyBeNZEkM9ptXbnlkBRFGcWDctcRD43T1m
WRx+6+OErSkxGH/yTL3uPh5FXylLHq2tb+NDHeHX6xYEohB2BcuEmNjh6Iuk1pIw
5vJduVElzhVAE76m+YrGqqM0vODQ1bUzj+Km56kIvwnnt0A5tR5qvLSgOdllS3Rc
3EOBtXwVlE30+2r5rHfGpp4MMozEn7FUsdlaoZqvfjBzjQF1+BFSfLYUtj/xIG3T
UEIA51UnMsi+u4yegp7SSrvXclCh5QzffzHOsbLf6Dus0WO9MUHCjSNeJ0Rbuo7n
YuHcM4gJG+12HWS1fPXODndcUPVMEPFplMA2HTO6QQvmWx12cstv1OSFncUiG4nv
W+mqfXidSiIOlAGeTxBk3WxJ3m+M20pC03VEdX2oV9kHLWcEMAds8ishBnPMyJh+
lbs1BK1MOSqZUx4+917StHko5IWxEhBRepnGK9CKoCQl7eA6W0kyVjN+SO+uxpAb
Z9y82FpQg8X3sS7qPl1yHMFC4h8Tb7hyTdZwvSLYTeZctf1zMOJpY03dkO8EeBl7
zuMX6bDyvD8qJgeWTAioIgMbrU8rVgee0REs8jkb6EdqYUGndSrnR5gCrDOYCXVb
n5AQ7tW7eXBCW9bMXZ1E5Egn1YmtX2nBSDj5ufZRTUvImyPSJHt+mqyvqJrDJsFo
vOPx1aDtllzvjXpe+uI/7bLWBS8TAlZQU/4GO93+nnAqw/4FaKEYOyZQLmwwRcrS
ym8JQMjNv8qU/m2WLBSAqk1VUSwNy/GG89M1h9veW0EAhDaTWKpihkQ2sZ1WgvMq
GvCzFdsii2eCy15LLShnIVwR6wRGAq+qhYxw5zIuMY4YDGg5iHPOgmEVRMZ9Ch3n
IRwCvX9d0vvLnc5kuXAI4920XaTlNU3Ckw6jQRhna2ktEiFDoI67c1kdrD9WGSsE
UPQ3o4es6mSmVaaA9YMql2s1gYUTsqVFk0iKfsGPkKhhJg+jF4HK3QcPoAwYryGv
sHXb6K6hPYmK9TrLtKfhbuBFeqlCpJzkghs+wRXUQZUD6WqhY9WWhdHCFTK4tGqG
t2PByERqBul2ydVQf6vW16lAlnMD7IuIKiaobyBRtb9mUTi0FmRof7FGXddBUxn5
UsFSjj2nkxIE2RZaeEHHG7XH0S+EAwzlUf1orAVSSJlLc3bT2jWXbwJp6UVYrjZY
EEcW88NBwP415+TkOeG6COhjS/osF9C6v7wBltWMwsOStLpIQTkiBrrq98pqgK2j
QJ8G0qb9XoYChJXNcKcMnTdcmZDdsRFCdpkOtCy9khzXpiDGL5J4BgZP7lOAFVvT
ESRQmzqJr4dfHmqwuitlE85ZuhUAmLnbE4rv7jTYa7faT2XrqTzMrzdBI9Nbe67Q
NqZZ0BntWOCm/f1aEBAfM1rlZB0S0SWb8wJ8NAAx0i6DOpOcJ0D/E2Mq99Vig3Uj
LoQpPHyRfmGE7n2fPTfG+5sJXwSR+11hlmU6jSuvwfzgp6iDd4v+CO9C9t9v+rKV
kuF/RH6TXX8yWEkG9Q7NHuPB59RBE0V1syBbbhIg9cF61HHwzhBNybjnF1szGAHK
wylx4Qf5nByqfonthTj2HwO1A09C0M+sCJ4xpWg/E7X5faOLKcz8MYOZQ4EZmc8k
hMM8onzhLhOYNoAt4v9xIQrbaxzxcidIYOWd2iU/ZonuAjt38kt8ZsAhpB9ibNm+
Ohkpz2t7gN+LdBM/YdGMituyzI0Sj/ezgaYMdBE9nTYLADGod3COHKxHsko0S9Zk
DebNzLCvqMD5/NjX6TMr/UlOuoV/7ryUD393vFUCDwp80WD18XXNjBQ1BJdvVXTI
1rn9OsTa1VU3e9zSwwrkNIEpX34quKLEO2dI2LSbH6xuvbL6GZfc1K4vROi0T5R8
3T2qL+QoFl6+JO9cp/qb4marlTSOGSIt0Jp6zzH/Flo9Cx6JFdHKt9GTFyMgzU3L
IY9KqONWMUF8rz2+++aCoBVqKjwYJoqH3NoyDu7gwsMnkq5EgFNeEYO4HKPHoAjh
0/Uc35nWZRDrUuWDKey1EHPo1bbuTDlH9096NcHydZO//vsEPtH3ennZ7QbLKC4W
z+xKDlGTSuvDCXBFJyhK5KacZaKmzJfb/RbTLwLE1A4rp3NKperJ9+uL+2X8hlzc
Cjs51Nt7TQR+3LSCjH0MjhTvBQiTLucujFmr5gojdrGno5K6YZbErZbDEYdNt9HY
N0mEoXdquSob5b3kUhIcsToJLMsZ1VjhbD2nUQpWfIkmUEixp0ELzgOsAyceCFiK
mpP1wD/E7TnjnyIVUas8Q4qzt6Ks16eu/Opl3eHQwK98NO8WW7n1WnMzCePFWLnw
VLu7p985/sOLptiylN0/wwKHwrL7MiVfaXfybd3akPT198jeaW6t+PUw33z5UvpP
fjEngY8I5c4gfAbvgpHndoukf8c4wxYpQaCmo39aqxSyEpUzefaOK0MJPMPIDrmS
IZCj49IcyQP6i3ehNy23p/yF3iW63ccGd2SMjQo3cQmkmlg9DmJEKI7lSEsaRUS6
JNdDqnI/QnEBHRfvE1yXh6nuqa3VVBkoFHHZC6FCe81x9lN4WvlVsBsA9Q4LCnsb
1/SSn1D9rMuJufreN5IYK4UgLZRNx6KtQwzRzeg9wL3VD5upR76z9/YbnbvWMyT1
5b5YLLHE4p+i57hDydjXMKL9PcRjhytJrZsrMa28kQ9pW9lTYTyYAjmStF2xXTSA
e1VdN1Ysi0pUx8yzHxStKppXukNS+vuIu+spieK2u3YCkt+gdr4YlVKD/GWF3YpS
Ipzi6Vjkvdm4bXU+koeeNoq2tSWYNwsPdnmQL/W7d+vbLd8oUndhbn5mmIrPuxlR
C6wc8/txczLtBUt7YOfZrLRq2HSp2CtLZgl4tPXeF45R01l9mvzL3lGyjTKMFNof
rNl1n55rgX1XV7HWchwvxpuoDXGZ/y8yqgJpWsVwdJ1U/TkIPoU9TPveH8bcJbfS
0Dyx6pNBF4bFZrW6sVloJdoTzR95QpJ38ra13kJYvW/M1rP+9HiyhOIPVZw+pD5M
HAl5sgh014HbPf1L+Pj6DC8RYM0qe6x/96ej39H4ya5qvu7MWBejvlkWV9GBEwVx
0fX1AB0yIyAZUPgQK7kU1eU0vJ/fvtR8QFTyQhLWpzP7PDTZ2QlQW5Pki019jOl2
Sqy1i4Q3YlAOsBFe/IQgXnJiULtkL2KkLGTDDegrX2qi+wS4QrX9VkItF4XoDDK/
Y8ZjA2LAp7tl+6uQZ0Q3fGtD/3NG1jZGtByEYLHdyoZmmf0jIWHPgQtfZfIVyaiV
qRAcOTzk1YU54MsGjGpWHEjbGdccOsfbcDM89hVncaLhRLwhcaj6y9OxW9/M7CYd
bwrS/y2FaF18Pg6J+Lswc97Yl2WTRwmzkpgPQn80M9I69f/Lh8oHmo9Dm5WPu7Uv
aUbOsih/e2o3DWfSfpA5eOmmhAQlhoA7B+aHYgSAkwIvzl997FGtgic2bUq4x93i
r1H6we/t3z3vfdQxKbhhcG0eE1ezS6N+xtbQ5mOajHiw+Swgf6tWsiXTIdvBhxcm
C+/oYzTFVAFc8eZoyuCetOcRGv5PmYpK5L/sPWYhYrj0ra/OUufVoYuDJg4JeB+I
VvV+hCWdo3i5W8u3XLE/t6tBP5jamCFK5k0GP4aVzrMQjYYS9IXW2ywnlGJGcEtR
3uNRy6Sd73YzqUjRpBJ6Xf9VDha4MBsSX/X2wJvNHa9Rqpzxe1rbiT2mmFUXaUfG
mpTHlQf5ZDL+JtSSoRV2hoTgO7moPxAnfeZXDrI5EiVZYsgMooybMeQygqUggBoF
SrdXDodIDxWl7wTPTtZK8ysRSP9nd7M7V2HgUJNnHbYiIDKAWwdV91ZtukTM/3fq
ResAFTSlNmqWdHB5Rzr7aJQBEu3sfD20spqfnE9CPVcm+2PE1SPExfXVgblXoWBR
1rcjIZS1UOTdRn3QM6E8q+PjIZ46b8nKSkro4m01bkjtqxhm24yj0tYBg3UcQqXS
M+wAKap5bv0L7ZNxK98btLOQ9Ls8pt34ugXtTzT+s+2gypnDoWwJh7OKBt7Hj4Q7
a+rtGAEAzyBkKLOvh3yoLe7Ur6x82+5W/uoRx67jG6LtYTNB/nbo3EukUykaYLRD
tUuVH1Np0/4FKkv4fill6XaoiysI+OswZBRrhzYP01nJBXUPmace8uKyS2fOyFsi
SCbo2BqaZz4UjZ4Hob2mIV8CHirk9LuZI6L+cN/swzuAzjh+9/XTacmr1B3vpXeR
1fyrLPGd3xwUft6HxVkifzNyY32/lmHg7ieO/wKAE24L1WEKIJ2hiD4QhCXm+nBM
HQEQQPZyz0JgczRe86IJLrAURAQSgeMUPhtpyQhXxQfQoTIAXom8W/Z3lYglimwl
6DUBy5QxDZd7OG07C7PmoWsMFqVy03Auxc0Vid/TLXRlSkb+smzrku32PA7uB+cG
ADrFXD/QfJRp1MWeGGi67D288VgYWULwgMH7MQ1hkzpzXQoeRss7hSdVjpSNuMQX
WSwRZe1wztjOdUpWGrdLQ6TgfjZodzljqEtfQhGe77YjkAotpwCGunAOCsn+PpY2
bj4GuEQsLeSSp5IOYF1U6d6FB6vCKgZpBZ33Rp+zTwkMn7M268A29xd/NpQ4Es32
AI7E2s2SGqj8isI+UVR57BNdbAU+POuzwpmh7I1WcCAe/uUBFVBP1nbo3KWaXB4R
eAaSbguLS45EHAcTukvWv60h26CSYluWvaz/rPx7qt5wnMwq4RPHSZHazemHi9d9
emwJOGtSydDXZr/WntqKx64T8gzVqxByljZbGOPsHZ02LMeTuUCx1lck8yI/ItI3
0ZX7IVd4d4HE4L4SZRJ0Jka5I2Ttrw0mfK1AIOCJvMLinXGnGRMBCIV3LSAUN7YY
GHaJP/eIIj1FLkhE9Wovk+2urO0bJzkn4fphnYhnrIvVbuPMJsuRnKb3I+ewZbAD
HL9hZ1hOUExVnj9tAwGG0fOMQQmG5p0K+EenyvPA5I8N9P8qgGqaWSZhnlvkt86s
ndhC5b6vCzv81mZxTZJZDvQRiN27CJnukj8E/hxoslqv9oCCcKDc/9G8JGumUq0x
O2QEKiKvA67YfMx1NCm0g3QO/tWu6FIpSq+Mnvzr3tdH4EKHBxvEMEKDf/7uut9v
l/ECkkU8ULc/KGe52lT8EUzcEdX2cbuLzoUA6rRSe/A6HL4PaDzs35/HciUBOuBK
qp7gPcOHFJUHGYSDVOfLXOtfFnk4nQ0ydQR68gC26ZDMurvfP5yuDB4xhSAhU9og
PUBjZmmnkGhWe+ejNB35N0Pd+BSLgmYswVW+pRFll+CS8mOJIDdf7g67XxCEQAba
5paFCAKsQ7Uw6xk7OYKk18uHfP6pyRUlsLdFwNlQiGoDlm1FNqLWuqWs78DTI+u5
qq+nTsbLyS1IqHrdcVNSZD6M5y8/QijTrYf6tasMO0G86cGDRy46oQ6YpyRIR4zW
mkeB0w7oa6mDldOGishzbQ0jFMz1LitvJd2TRe6gFYZQ7Gt7L9/101uAqjFuoLuJ
W/xHgKQ9lNzoQL9WISxAFsl6FxBiPLxAlHCFH5vHPm7mpaZ+dqSrSihxitBQhBLd
LNcMsGEImEO8L4JJdSyt8IVycwZnWDbrLwJmi7x04glX5JakZPQXIWsmepuzoIHX
kTDYvnw+exIkot+d+jogZUk4bWxPLgvlypEFMBVa2pZuh4/zKF8Zhu3CTiOpM1yw
iUw04O1X4q5cw1OuxW3OqxAkb+dIm9LINswPMmGhPh94mn9Ou0mZX8VouX9SnJVh
nCeC6o2MYIvj0U8MGIztB1f1veSqswA+OkS9Rmxrlwu2GU6E45Q3zQmTqOd08f/k
ERvHto0359WxvqPAP3Yt9Gbv+ay6QfmfUQR5KJRIbhu4djYsrjJS1kyPKhlsZerq
nlwhwlPjrInAMGxwD6CubmolZDS8gmwwW7+EwjbHxQcXB7GI9CElO1IaAwQ0jiMA
qOxMK37rBwBKhoC4VTkyGpg0Sea/+1hGrEiSN6X9X9DARL+RYbHuKnsNLOKLHIvz
qeTpqpEeMFC0T7duYTFNeD1gHqJPN+EARyo1jU1AWdkHUCYZakdz4uKU/EA7H0vd
3ZAuenYbIc1718EflFiEBN5wBnjGPQbt8sb7bPRIZUvhQuLTriUWnV+qxHdE9Kl+
Fsut1fzqNj6avfUTypzOu0gnFe+yh7YWbcVmRW5OvAuAa+gyYh18CxMvB7/2n6gq
USPjTfZ1LGlwxoAzdEHUhIjRh1dnFQulWWNaGwhZSNFy+hWBnoeN/uFwXERRZeav
HF4ilqUGiPGdq+GxmDv1wKRw+/L4dnPowoPLpYg//QM3Unj1lT3zbLrTcGnYc5j+
ZOEuy0l9wkGbYMvvRTKSlNjPuWm3H3TnIBc6qHHS/bBqgfFUsQPur4sXVQrEc0oo
TuAhuJd+H4yAdyyw1k/aiQaz8KBM1FpDxu834AaigxnHzE2tc4JHX/72SpSU/yob
bryHT4tMluZOBYyQXB/AhIdmrdSOB1cGhD2hdk0YWYcRkadDhWylpSYQ8MntQEvh
hz4Zoa8/lE0AZ3zl9DqTa99WGcJR8hQo9m6QOD9Y+55nQC5bk6TeP/BjB4sa5qbC
Ta2D/AJCawYC67hwZ0sV63Xxzdh+VRsZtAyyiypHOE3uTUoxFvXLfHQHzpf0Crbn
6TaABtLCkViAtVFF2zOxjjzagDV8ReZWmPEdJVf+cG7iv08EOG6fikyMDGpZCgHK
zyAP7r1ry9w688xlbxLSGx++dVA9AmBmJwkpaWdQAA73gYVdfh9EuZX6J+agXlM6
oRA/3aqkU7EopxoQPDirwzSgPn4baJk148NbVQdGYLSk/DEX5mkzs2/GduOC2/+C
43/fTYJdGXdCfZ2UptoTUJrScV8u08oZew3r8kgvrud4PAyNbK6DywMHKRqO2xgd
Tqczri74H5aaj3wXG5+qwF0PnWH4fAjrOJ1ZG4eK5uT8CvVZ2ZE98QLGlDHSj4U6
3KnPmejewTbB4aJXAb01er/DdFqAn9HhPYRdq/Llrcl68oESG4XlJHxfOBDMDOVZ
upaJSNh8u5QlPTyXgF7Be6cavto/2sk84SulEOd9FWzkdsJRWGxG1YXEPh+EgSKL
CkTct2SLjR52J5K8NMnc1PXyHwHyAQvnq9fPdSalfsVAxaHg9bOdMoPpmdZLeyqh
JSJ0f2BBj2BKIEeEgVDnnYZ8Y4KGPglCvd0YvoRrYEerZmEmxHr4HzxohwEZ5rOs
aw8uoPItKrdyzcM4RQq02LcNVA89c7FTkX6/Q1wPXIhxHJm6itZJjw/s0N/ttCTQ
VJ9iAwNgKcx5os9BkmlgoIiVjFOSruJK1IQ2ZeqwFjrlBvL5rJpB92LIuxpGdxHD
kRsA9z+s7+xx8ikvserPJr2SZFvPYyhdAtpdI2YNlRH/SI7XniS5myTykcwkYRoS
4S7utQZbVxWz//1g8Yz++C3wcIlg6Ey/lMaj0kALVHLF/92DI8FJB2xvqHknUrkA
9WcrdRf5JDo3+Ia2ajru5QnS5y8KO/GYfFIf6rLxYlLzIFTKDj4dP51gERCca/Ud
0piLVdCOH8jFoyDjkXSyVSYKjgajs9QA33XNvxGxMRFM3hYMNrC1G2PDMms69O1+
gCDNvBHQf7gA8QK3kp3KKYhmFbe7R7K7VrCtN+QV9F0LeItyPWCGUqE4X+SFnjlL
GfJ7OZk+45gMZLlYpAkI1VHyC1qwr1Ufm+JbJIMFUFlsBTZybv9Y3rLI5ILBZDN/
PxNU6SSRw3VsDaDYYYeHqed6PVgq3/2Dh9w9s61LVVDFWMc7dHcK1oTlh5uRH7xd
FdvABxUt1JC65pBATzsnPSUzCcE9+labFjBIzS5ykrpQQlosdBJgZerm6k2I+T7z
ZCFmBru9cCVt2Tj7PyTEkyyvJ03+x8G7FmnhfpUCBpFae0v/dufMDwiYNf8xYURN
SqVmEeNH1MBy2UsqmJ7vgfsomgwIXYVX+c4IU10sNXvmmavl7dtsnbgSvw5SO2tg
MJzEdaa8VGufLNoIcylPNO2JeiTFdafyklvDDu+KwNQbOunbYPvjRv6pYmo9snMF
/54SbKzrWPBs7CeS3JKQPh6LglHWtKVWumPPZD5BAQi0Je40ep9fd7vo+Rs4Ok0Z
ekahPhM9sXoMJ8tHTP0ewIi7kgGOADiB4EPtuQIburgcOrGPHPXHxkT6Gxg+xa5P
LycJLRSig2RvFLEqsvz1/983q7joq/6F+1q338f5inoWyyQP4LVmQxOgb5U8rPDn
qFfaQz5sZdvSkdx+NcJSMHZTD8N77JoWYPNElrpIUchokEc46bksis1WChiaEgwi
nsIZVBenWWsidhGTyj58ga8IghDKiGer5SS/3TlR2xLwvFDXHAknr3OYluW3O26r
9pFd+VqaMHmgELQ+WwWLC1Ob5RLV1DZPM9aegbi1ENno8yw06kBZ8rXnNiEaOsXb
8xWpwaxFeUWxVmnMGOEvbSYjXQBcC6ZQkZOZbHexAc4T3O2movTXliVD4dUjXLYT
DRv+rZN4SnoeBaXxZMaIkLHSTUYG/WIIVGIN989pFa2JagOzKDvLbBTZDpZZTCid
RmYloLhJQHWpMDWXR2aZReT6Mz9I7z8LrrQjB6vS/V4KI4gjXrPZVS1QIm4ex+vh
QThn5kY88oA7dwnB3CHiBEayD2QgdMDr7W796/bvw+aZzNVrqghThJ7B2MfAc63q
tL/Nif65CRCQYl1ic2yQzGIjEYzBeeLYyOq+0c9nVO1TqqwRTpACBURJ70KA/jdQ
ybAXaGg3oZZZw/zDeIzDHYgS+7NcWT49KBAqhdL6scyZ0D1UamXbYWT3DHbeUKR4
9d6umaGGFCrhrhRR+agSRH8hb5dc0mN0dOQDg5HiA2BszLd2VMsaji23u5pblDZe
p11E7x/iO9H2+NkiJ//arKXdo4qIrWCex8/ogsEny4dyl04T25IXVceBNe9jaSiA
At1PSJ8iuznKIxJS+QTtLeH83cfhIhJPfmJeUnJFOKXGtK1XbCUzGGMSM1t8rsUx
uVjNxm4spTj25JMJ/+xPnuOWtJUbGwTkyQzJrSOfstKEVQzcDrGnm93sl4JA3jdx
MpDYDNQ5WTBgopSEtwTEErWjf/Z/BGIvpMugslZ43GjkWkJ6Rw5lw/t9B9wJ9LG5
2BXkc9XdlKstNlNoeyA+rV6wbWCT58nFX6dVQ6nPS8B4cV/9SfHmfUvL3oufBpqe
yZtA2W7H6gYhB2iC4IpWaVEvmZ/xuB3DO/ttUasbx9Becbpno7feLPYaJ7kqk4RA
QtcQ4VKVKA5DtNasuk4Eu+AWhOcR5rDby7vaVZlxUSp+tDcX8gwyiVjO7Knuhil+
8VtuFC2VYNStZdU/zxeCutjeAFDlKf63py5rEtaL5wQRnE32/cW3UTL5pfA65PGw
mfJk4p+tz1FONWhtNFR3Ng3OYFfbjHZYBT2xL7Nw7gdHLmhzkgQaac0jPxFS549R
OzMNu1FDSA5pUcbcOU1I6FfQcvuBZxBmzR37qhdUkvQ3fH79IvK2W4nfrwAQzm66
7KtM/EhzvIW8kK7faYiqG42qT4f72kfHpmc2a/BSi5Z2B6xvOZFh3to7OIk641Jf
T8QSSp/tPxSULPxB0f1rjAXzmRveMMjnAa/dmLmOUOZxQCTRbfsr4siaIma8cyln
bnjIk+rlxX8zwsLcqju4kXcQLpCar8Ife4RE8qt83/FcBVRiXnahH8sooswXtPxh
g/OJ/PRcq+gCDKWfk0aAA870EvfpD1c6ft2mZ8NWYW5Q6X5O4OUwt1Cj9u/KbFsd
HngpgQPyiBYZDMqZHwuIsWtJOWjMDf0g5mlw2I8J4AhjzV71zh3CjWLloG2gd9QS
CmUcfp729HNjsyQ3wnmzst4DV5DThWvZBrzBBTizbM0OnXs5Ns3JYAz0XGyrH0G6
g76zC3h9SCv/2NRDX7Eavk50YTRwwz2KQQLA2AwgHYPwuC70Td/u/6muMWcKVAiu
fdkPdcwJYYNbR8c3FORa2G9KLoS+i83tVNJ+X2qpOrWdNWHbsPgNutsAgSI6dATp
42Vi1fGmuejDxC1y9k0N0Xc3YxRctpoz9aceKFE0imuJ1QXbFB8HBNEs3qby5LKF
ggQUGROt4KmIv7HCtjGY+OQPQve4D2TTkYDfptJPuRg5olDqJEvy/k8vGInDkbY8
XOxTy9DGjMCpJlxbawAVp1imghzndcj2xv8heq0Wvd3Hq0kXkg9IcVomFoKeA3Ur
tFIvhxR7lSHyW1csDV1+eG2WIUUCC1+CZ9ZkDqHGU8RRIQlYmDabfge3IudETj8A
pH7WKlft2nRYdFReySDpB9UNgK71fhPUS5uaOmaEyG3crhXh2Gg/aXnBrFRxK/Du
lWYTQVlIhQp29zj8Ov+4Vg==
`pragma protect end_protected
