// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:36 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Db8+w7194OV84dqrM0RL8k+JT4MDkAdZM9ezmrnH4p6sfe59T/PvUYdY5vzCLU+k
gDi1CjDY205g9hFVDFJM7GJ4qqVCHVMU1JnLlAj4YFCagPHferMf00Eb6qtrYerI
tsn7+1sR6XeuwY8xXmmLl0ximgamVyLmL1hH9Q2HK5s=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11328)
ib7ZsxhaiYJDBV3cJc2iITmKaNYViOB87Ag6vr0UIPKt5mt+Hl3jFIhVN1t19kwR
Q+O6hBT6CUjpRNsBTEmbYxMis4abAdp01bW1dqH2rQ2z4SIF2bUTS4vL322+w8+0
bcvphqN9lMkLONgtrkuLRNY2GnhoIOjbxQLbWRgG59D+LDCCBroiZbKA/R6Voe15
gO3pQZHNrwIonwKq28es5Z8Vl7SQaUMn+mJG+tfcW/0IZUSxpDOI2g4jDJzCdstj
JhOFd2CEDPCV/mpSWYoh8Oz7NYkiGr3OOHliNev7HvXlR/PwTi8jJY39j2znfSjD
v4lWa1XOM+xh0TGy+BSRx0MkYbAe2B0XTZYKSsJp1677mLW4flbUAkmBVy0alIDV
ZVRYkvyuy+5qbNCvKL2hz99wX+DRqtCTYylKoZv3nrvcSwzFX3r3tgLJQ5bVM8UI
lWHTtfAWmiqioujf2Upkl0BMgg6nWke/2oB5+2RicMHnIK81YdL9vTnP+BDctaEK
qJk0thTnjBL0L9hcl8xUsM/y2I79+rpCPHxNxNbbrwyO3qUemxa3Ofu0sy+HmJs/
L3foyAapf2PPltWL5QH+y9oVOUICwyguC4nVG1yJOo8BJ+38AsqSLNPCNzweMwDO
PafQ8heGV9FmLjp+AX5jyn18cqxkzfY5hB8WWaJLMOmuJ1NVzsTTv2kcwJ3VldaO
5NGA04u43WMQo07grYm95DDZuFczT3c3NZ4oCSsDhN/j4lBJBfz5ZFriuTsSRoTy
J1gePWgck+JvjF5MBdHk2MZeXsAoIE7J8IPIG1O0ufyIbKMBWzs2nkCAmrgVl+XU
M2Ml3TjA10OXNGBmjvG1A+VCVudRRahUjcvLvCtypoIada18tZAkPP0+ci35UXM6
acDLq2Qe9jvZCgcOUrLZ//aLsoaF3/9S2cAtTWNG90bc+nptnoXDJrGEd9Vkzpyi
5R1Opf8f7WvGOlSRV5HmYpOdQyH+6eynCQfkYGqER23ftFhyLbhHB09oOVLVctlm
LU6C4tQTj2jYmNMJhjcCiAsM5+KD9crdNr55C+9d2qk8z5C/pIbsogVAsxBXCa/s
YrSpCVqXZfWma1xIfyXRUxuYxRTWazfSWBR6Q7pDWt/Sbx8d2CL/jixLjw1MY4Sn
0PdLij8lgSswQYkmzfP6GYO0f0ISjc2nTATDhz9Gp/X1D3sKMbDNyaAOAuhe7EtE
u9tj4dTYEGS5IFIniM49YEVS48SjdJiWDf6O0FbaLqyrLtC3vRZSFZm6NF1TCwuK
2EG3dtTOUKiPMauyTJGyxO0V5JgCcI+99sOe9vtj+kOX17hI9maVV3kAnkaZr7qk
7LtEj5YhlJT8q7m6z17U7a3EebLyweG7/S0eIPUCNbriN3lH46rmTv8rweBroXMj
RbQWUbJLMcZB5JXXVnSPUfaWZftvPk3MQdY35zZB1GSQ/h4f6paIc3jDNNGMn2xY
xAq+nVBynnCscnu1Wh1A+CQeakv64IHy2EnE4eh1kIt4zmk8fhGtwQ76v13evyeB
S3z9aPut9TBYMf32q9TNRkWWtu2Cjc0cqJMcO1DjiDoxks8ENUkilFAxbp+vNJp0
l1XLsKP4dgtwy8RHhbAW7xT40+YgTbfUz32y7YxLi/HWFq170wdUJSwgVL0tiDUt
ALBpoCSsioUIILwDLLgTGI/fslmM+aHUo5T0oET7+HuNuvZGn0HdLJl+8x2Kp1KP
CJLEsU9QaT/GeAQUVJR8Pyf8RQ/dDE8/oun3U8/Brh896BKz8tfEIA9VpNSiVBZY
D9G11PHATNKbpoWNX0Wp86lRAP14O+6fcpkGyI5Ain4MvluTLyOr2zai+Wi1R8qf
FXC9k/91eH0IS+isaoXHc5iwpBZ1avhQ1v/qrGfgeRyFW8JToM2tT7GvO25IJBfI
81invHD3ZsgbYQQFgW9eo3XZIGILDHfrRoINM8iojTV9WK7ghvrdkXKVzQvXEfOW
uo0DekIJsN66lcH9GtAwHwCEuU0yLbBfe4Cdej/TsN34fV0di//QahuOkF22Fyzk
GEyX2RemJa/8lTXIWzuVnBQ/oTrOd5DhPO0UTl1zeFWW9C6CECZqVmD8q2R5v+sk
bT10qJxj5jzaFl961hshJ/SVGSwMVzYi8TvIT9B+YyEHOFP4X/ZVLrg6spWPTyBM
Y7c4QeVBJ/H+nXlebc9w5EqMfG+xvFFXyOjVDAemld5mvikgSksqdDh/n04myB63
cFcYnJg5m5fkEPdKdrveJnWGwpGASuDC9ptLThMr7RIef4BRZbvO2obVQxiFxoKa
1rJa6jSsS0L388Yjg+4d/G00kdWBt0G+jEVL0P7729ZvZZMGBHFNxgbGotyEyTI1
pLPWtM99KuMuaf19upAKS40/B7imROq87PzTONAqVp3Ks+OLGDjQA3l4+APAnRqP
FlO4nVDb8/o8y7SoUUF0n9yLagO9iSaN9H0S3DplLoOTkD0mCIgUojhUmYWNPFOt
LEw7qSI965jl9fY3VBZ2zgxIGYadwrOd398EVjWwigH0Z0KeW/D9TqTMvkM7p0vy
sNJ9loVRKE5MRKStA2cJ3IrWBGl/FBivt0qtTragxwzmZE3Xgmx2TjuIHnimj7N8
DMxVluN6ujk8fEhhnz+UAEg8wu3IoFrxg6wHC2DkmWMfA6kUFtWlobIThC6spqIZ
+u4ur8j2V2GdTK7fzP8OQJxM8uWGGIMzunCurrmJawHoTaT0gzX8OcTrLlKp9k1t
Y/Ecvo/jQ4iYOUpaKAGVD03Vt9YBZSICY0ptmyK41lHpoF1dMmuOrcT7nwnUwXVe
1HYPKyzkiZB74vfq4LliGyeh/yS4z97M4YVmwXelIfply04w4pWZK7/4zRaPlUna
DVJPrJ3tm755w34x+apRq1Nk3GqXgyA8dNtdMHh8LP5NiMVzFUUnkDzsWAPKRD/o
3FojB/MTrHaBD5FhJVRqeZOCxbD1AfLr3+ZxTqdcixVnSwKyB2vtAgnkhgYDJuhP
g/vszrbPwH7N+TJT+bTrPAmCNiY1G9iseyyxcmHs+Agr5vvERjs7o76+gs4aRpXM
erisH4XH+qspC/OMYKuyht29+6IJUspoQpg/fid84ShaRB0Xiv69FN3pIDOhlp8i
ae602fcddcdK4l16iCHWzXPuRggcfM6XFnjMlLo3ahMbCzsDGvWMjZjRYphBxXV6
AjvAwgohpBytW6l2B0SDBHloiy8j7fVO0XiQA6HUNeB6T84khOExPsnsB8pwIRnC
1lGccORr7NVCdLHfOjr+auxeva4sZY55QIRlHT9Ge6qJTneAUCBFGaCqcxIB1+tN
GnJR6yzjIpHuaeMV1ptfJEWrlgiAIwossoeMMtMfqtJEkdK+Q1bX3CmK4Jy7ONyE
r4ICAWQZ7PT5GTxCfm7yWOXZr+nqPUXWrAffHahngFA0dzjrY6jeZNdBXSsrqz2b
TdG3p+L/Hc0GNw6sL3YMnJN0Pivytq+Cw7ez7/yarr/x4cEstZ8M5+coWs5VrOV/
fYv3OyTLLXKonNMjkBrXs7qXiisgZ5w7B1nRRPSA0RZx7UynWZQzE88dn6OVxKXE
e0CuLAgiJMeZn1pIMtmDk4zQ5VDCTmaDqLQlTrP3Ja+QF0MSBcmnfkAjgV0B1tih
jGtXQMAGKnREa0gjuon7rH/yLkbS40PCwilqbQY7h3xjOEqa78DQgYTCjYmhxvmm
Zw/OToHtykA7sGKnzHLqPyGkhnJcDj8AjYQZtOzKGqmnF0tICd/WRQTaQwdw21CJ
X4cDdW5v6NJhLIdgxMDEtVpFcKKhOWxmm8e6MLCMFONrgp3KQNS4+cDsascdb5W2
6Uz9si9WVtej0ZBbXKi8H/ZF8+YI4UlgMBxq935LqjmRhRb5Rp/s5rwt7QtdBffN
/o4ebMiFxgqYi5xO11Te+veH9gjveoHAaYuRvqgNGPqP7zg0S0DDso4qQJ3GKph6
+xRJVtHjLA2ZxP14OTgFqMBvsoHPuEd/hCZIx0Pv8hQO/y8NEKxVaABOuSPt2Rfd
yhroBmcnNBHX3mNV5QANrm5j6PM+eeNINGatxU2x32nV8rwJakY+sCeAt+i++CfM
njLzmXzbnQETA0JkJQfTeuEcWc1SCFGFXyk8UAZsqCOJkp6KdCr4cp6N6jR07rRu
OWyEXBHPISm1R7qye4ug4fmhcadtLoem7T5aULIcH0GHHWFJS5P036e+qpFZZWpx
qTT86pNTSp7iRDkgxMGThHmr/gKUrRYxGtUbODWM9eWtZfM7afNW9ahEJwCrnVR2
s5m/JutgmtVaR8Oz/JFrzI9kSQEl4TE+SLcO7M8l/jGxoiBOeRZLMHeSy1g4hetL
ugON+JoZfVgM9KPnp8uptJW8q6Bwm/Vvq72juLhzXoKZi/5ebW77jVZr+Obwofzc
GZAuAFOuTruXusd++wcwicPB0Wef6qq07HnQkicRGEBADeTC9pXod4lkOhEa8K16
KRfiBBxsKEfIlBKCCLC00rP/xxU2cgYVaTMF1kLba0Me/BASD4wVfXxMYy1m9Go9
aDPRFG8oHAzDgBf9it55wKDuzc8iqnRtjNpnhrX5Y7SMH1FJrLnzshq7QMFix0g8
LGeuN6eUWDslUx5q0tP0R/cqgowsMriPOTCZGCZywuIo6LLjfk0pte1XcgVtbC0Y
TEgifkpuKb6rYsPAK7k0eZycQo8emNGCapsCXZOanDc2yz2IB8G0bdFfEq3VZwB7
IgCXtkDaDYBJegT7miXN8wMC8+jC1oNBnZPLoVL+TzJnExVyi/GF7wLZikfFZPil
rlyZt0iugcnG+gFUNAgx8/sq7jsl6jAjmhHzPvdniHXbaoi30ivImhaquaFLSYnf
zq+wrbSraRBYmMpdeSEopMfgK123lY3A/RP2NOPOPCszq4R5buSJPJp2luPoTvir
KbBl6YuZjFnW2MOqKUwGD4SiRQioOJViAk85ZnOKutNSwr3p1X2pPAQy/OO1abey
8D9tLOcnHN5gyB9MHabNf4QSYzddDle47fAcn9P2CIF6iH571+27JKuQzFsDVRVs
RTxMtbH7gexrvZyXI3lIhkRuE4oTy5o11QBpMOi1TbQ9OIoSMbnA7KWT9/looaxR
OC9Qd6NwHiW+fr9/3xgzALrNbGdb/EtShHNj7mXncfWxuZ/x17uYNVcO/1G2wa1f
HTVCei92SyqjGW+ZVybybTdQtXoeag0Uqal2+YSaWBtFbFTyxgltp9PZ2eEqwxyh
hFfmLqJKmt23yhe6Ns6wM8lqaKZBvKVM2OSCMLiT/FMJVfRmPsFEem60dy6K5GH0
QANppdsT/hqxp/QUddFFm0d1Au6oOLn7NrAeBfhSGuKHlL+5cScrsxSNepjF8+p5
9SWMfSgBKEe7lKF5LEyG9ttc7ICggGlidD7jtUHTfy1mD1W0D23Fj1+kIGqy5hdt
knsr5Aogvv2hav8dmlyRXGFIx139BzslBfMbzkN4xxvkLCadFszpz8uDzQ50RJvO
uZqKy3hxaPQsIGdlZh5PJD7Mo7sH7zMQIkTDrfBoV/V/u0PDdK8U5tfmbZokop4H
7moXq0RAFXBViFUCzRXU2HqosTk2f6B3tCpXJFmZk3/M+NAiSZixsyPuZ9mnwc+j
s3olSmKTqdGm78/YGp3OG8O6rTc1ikzZLGBKSvJ9nevTHtVUT+YbEgG74Eh8WHUM
ybKVcs4/v7GR4RVsMAQxqN5yAki9kjR3CDAKJBt3Qq0M+N920MI5vVaQ1G4uOcol
Dd3kfWVo6D7fuYQa35YKKlNkmNFH5nk2h2lkJcSlupiNVPFLJR8pEUQ6kAf2ZkEV
JfPrmSMfOUHknYvQjohK7oKt1e4IgjmjQ7EvfS/GqKVmwRQzGNph8FGb0FcWV30L
3gBJQ0J4zJG4xuFeSV4dKszfNEowthwC8VkxIHtH0TFFlk+b9noyHzJCWvnXbJFG
nYiLQG1Xlk2utO+CfBWD1JbnI4LjNWRjoirgc7NRAUkrHqxVlbDqpm5DZBjvoney
nj8rfbyl1W60YH5G4dDz8VFQCqm8FRFKMgHXmWq+FiR6hqAqMd9gUyx529jV9hkZ
+/Ly1L0wZjiPt/tl8EJXDKcjVF4OTCwYK0AYyZjL621AIPCJeSKuJxRA+UBApA6i
rlyjaEGL9nkX+CjXVN8hWYqEjAl62CGv8QseqMa3tfEbGRBcyimO59ZQRe46qPAC
yT4NW5ZJU6Mf4gtrKE2OdyaStX9OJXvSNcHttX48L+4ZTHrHwVUrluvA0tDKTl9u
3GiHFwZtoS1Hz/Oa6gPOj8+p41CTu33VYp5Kf/HII3p4e9VnW+kYCymER8XQrtVI
a8p2F5vVEnYspyoMqqUtwGx9DoGdVuouf81o35hK2JzbwTLERad4Auqgvx+0OKtt
j6cgFbc07APYSbNEf0GHKMOpNi0qS1rGxOXxJvVT4xNg5uDkYNmePCAXeu3Wg9dH
p2iMPwaMPeloRgaaY3q8/+AXr28qkdYDzu6yYqE5s8ODeYd6HiyvgfjKGT9idZXi
f/eet8zbqJbom90xL+LzMZuinOaklYE1ELo9uzzyj33aPjCql8uBfZtJUh1OKiO3
31x638EVt6CcTo7fFYJWIPM3P9T1z/YHj1qe/QBoOpezPCVSjantOAY2ui6kONp8
oahMnVzgVVTKUzjE0j6LugRqniQd5t6KPS5qjD5IFB8IkXZrrt3JLGj7V3q/7xiZ
nk7nWcaddLWyfenOklr3GV/Y7u8NI3yc5/uupvXDFiyNaH0FqvjwT2zP58vO6NO7
f9wT9JPAiQ+YntOfEXnUWIgffmETjDaYP8R9uqCfr437vrU0UeryX9W1gUltiLFU
7xkzF3uDU/E+rSyFfXWGlsDQF7PLj3SNNfNUWkLZQIbAX9xQ9es55wYgTJpQApLP
HzVn1gONOvr5nOxwH6MvdAiHUpFA822b0EFbcvGDzogpPBx+JfsNR5KF7cvIPfi0
6w1Je59Qh+uju0db8KGybTUGJqos9FAVSeFfMkeXyOhZdOX6brXFeKuZKrR6CDjo
cpFLBqGkr2hEZE8mgCVp+rzsfsxUYqVbw3Gt8ZiK54G4rnHfMxNoOMsGzmfZzdNv
loP1nTPDolRw8NaSNVNCQk85fuL02YkLLmlSb1wLAfhwtMbKL3lxH9TY99ydtke8
90WfZCLE1HgLINp8IPzov1AdEIdXePnX+HSnaOgMwy6RTNZ1GfMmZM5JVlqPOd9R
Fmrvq1Pu0SsYYpsAJB//gNr+GLbgkcAH+r4jv55ZQgIOlQmmc+LaSJqM/lz+F/z3
i94gXaI9M7ABsCU6ku0PS4zCycwYn1A5yy6BTzBsLbfPGio/rP6sQPe4EZzXb6bA
p9TPxNjwFAYkw8/gVLQR5sP4VTGkRSYXm/oSIc/4xkSziixsLXtMbnDcYt2tX4d5
jnvVlqF8tUwjJgcsAvReCaiVobn1qXpWNpp3xhcZklK3yAbS6Qp9kcvrstd2ZytN
FhQ4XU8KJ+q+q0hmyvXZebELQyv4jFbHxUcFyT8093MTWqSK7nzC9zkd/iUAiaak
x3QwVARmDiAap3P60WiDhegIQ9/ixThUnRAEATd+kJMC3dJEz1sjjGsBzG67T5LW
Qk1EOTtRAlpF+5Rhr58ElmMMmYPoZruPxUafifmvAIToA8PuSSddjm1FOxXllRE9
a+zRk76ojrDL2Rbc2AZB2vOOiEXYe6aB6LrthGNy4tn4O0MQ8a9cqSRuO9lCERfZ
pWZPFUsQ+0xPJLL0iiooqr2fSW2/ftD5zuZmKPXdT9gxcVm0tEKaG0uC5+wJsbyJ
H9JURKP1ym3Zw9Ym38wEw7W2VmKKLyrnct5YJIyF0qr+DJlfFp7uYIgYFj7nimjD
7aD6R1886zEYE7EOfCaEUhJLqoYwKxbTxzYkroYhmSI0Z6qYjDGkncsrn7zUxMyV
SMBvghw9HDMN7OHnqaT3sabqtR2fzWWXxgfQSDjHFNFgtj7t2r/lRLERGQ8flQID
cZWGMLP7rhtCSqIZ2UhcpMoHxRbLBisnkrsmSD10B26cxOEiz74A5xicKB6i19Bi
4XrleI5ITkoeqapdA028RbNRKliyqUr1sw8ZqT+/Z6uCOZp7BPOyubsuN8e6mmrU
dlg10FVr36GWoI0+34y4YO5koeNIeL3ElipW0OQJrofiliI53im9V0/g3aV6yFJA
ACsx4tzNHMBlT/2X9xafC/9CyMoRqh9zVCZMVMA0y23KP5fgyMVZ7caCK2Mctovy
4sQK27iWfVdg0F5eSBcnS5WwAhStZTJdA18cXU1Jc301P1UtrOlETE780TF1LyuG
Cwns4saezWolKMeiNqIOJrTUwbkUYLq2utoHGBQ2e5bNPfuKYkwuiqJBsba+PLso
BiTEtu6aDK0C6f8AU/y5PTZ5YFkx0xi8JC39giBGI8t34OUMQl/l5QeugHLlJw23
UHOJgkjLjaZ9f0tNYGsedcOHfDJbL+aNeikn+6Cib9gtfJMwPM69JpCCRSKTp1GN
iee5sHnTDZ7yN2vPg3100am2YGGiIUuvABcLFlUzLfV+Iz+QMEsFSLEenFx3twvg
B9M8C+8WJJun4F8MXRt1hwi+oGC6KFvmuo6sXEXQaeNm0tvjyI77fhEYuWwoea8E
xyQ3ivQcICWu+FsUPqAJJnaG5MZK1Nbt30D92/Ku8i7cYPgm/ficHByP4XRHIitI
qvWwSefBBu8FO0mieWmES7hIHjgbzkMnKcQGkDeD7nqqz/M4mwWRInEddGH1wXv4
HPjO4IyTGIWz7MmqEY3IvK/qa5UzV64kU5DXhqhsT+E98rMbHMH6+KtL2c4vd67T
6M+4jtLsWGHvbSrdQ/ZTMRYPmuZNSFPCrzPIkM9HPmk7VxoFSMe6f0amuNkSf2u+
4QmsjbCi5StRqySsbfgoYFUNJOzjzT9gGVVgP1VXZ0Km3Mr7Jm1dTGbGyDJlT2qx
DIA+dguSDPCCtxNaKlCTIPouRYz4yGXouKGZsB1GQ0VKP1tvAF4yzbaIf95k5jNr
unk2fquEqLEC/UCd/6ocQ4SeHw46O+ex1sQMHeDjRKhLNV0hSh/0a/2WjdXCPrVY
2xYo7fZiRxjaUKj1dts0Riq5DZz+z9j8HQEP2iBTxKgxo20s2OOOUpVaHAtpV4wX
I0eGBjNHesTDXMtB0jyhaCicOnGSntJkQiyE5xLfv/0hwYf7yjf5tHs++1FZilAw
EynfSxrA4ahstzKVSZTbsqs5Eip3B5FeNBx72Kwja5Cl62k81GIwNbRxH0gf9uK9
BPpf0VllOMPW1I96/hcrX2+QZtzY0VrxDmAxAoWh2wDRzlCWzlFPAdbl+/WLsuZn
/vku0U5stTyeKA4+3uE1QHfQqsZnLSu1SX0ANx6eUN3rknDyw8kRekzQ334nIitA
h2pZ2N34hE3EN7y3xX+VJHLcc8Ad3QsXfMnNSTcRGv8IYPEh3HPB+MpJPkEVKhsi
8Jl5Cr9yXzc+1T6UyME6dKFOmnIA4Vsvu5KcUzxxaJhJbf2UtfgOPI/m7HrpSwNv
Jy0QTK/qp/LsJSoz8zejla1z+XiEg9O0LFEp+M7K5qfEDOl7/5CV4AYXQBO3iuBf
Kq7b0i4jLH9ILw6oBBSnxIVAVSUmCATA8GmLXMOAEeGbzntiuApxJE6fM7mdQqcJ
qoePztIWb30rqmzVnv4env6DjiZSvPUxB+Zy9uPcozo6UJPikHLnqZO7LzdT/iGA
R0LSDBiVIJfHb36MMcq5YYHlfvcEjz2mupEH0QHEm4vlmAQTWlZHkkYB4QPTn8lC
ecfGq2yaOTQkRu40GI/WXbBnxl0zOmUf1ao6KLVFPUw61Cyv9oziZt/2jrVSejOc
S760pkKnCsE4EfLkcR5bzfmYBJPPI2WeMkXFq4iWiqakeYORWmrvihj/eiPcf1Xk
bzcq0/Fae5FsWxTDfr5O0Y7t0fZRwtDJG+h9VE6S7LcoRTV+prNhHYGANPM4bdAG
IXEWzeD/07Er78Sni8KNNYEoZk0b+giy6wOLY9QxItE5/y7U6Fm34m7KyWy5n5H7
mzmTUE0HOVvlyEU2BIhjlHKUwZIYvsOgpEMjHgQiGBBACQxcuM6BEqgnxMkrUfeU
4p50UQhrqgTGdM1I4CE+zHeZPZCh6acl6zYoFQ0vHm6WFMvstj4akImWqIaxE9oa
DKN9rZfE4MuiAf2x/7pFM9exLmcrdy2AyK99bjSPPndGN4MbjFupBCchrPQbxNTz
kke5c4+h1EieIKfixXhJuucl+N2KNL6Iy8TCmklo8eIt8PE4t+02tyDje6LULYIG
xdxF7Glgqu1zAJWDY8+z1miwlZVy5vBInJ9AGGElMJbZ4XTkxIXbSPIBJSfXDlXU
tjdzoitlSIsEHMsTd5SJT4iySASV8D12yhtPAa0L7GzhNNkX8ZwoMjH7jIdn28FN
OmtqimiltkaYvcs/KVBRzOoqft9aaiEu2A8Yxq+PX1tIqELBStpSAJS2zA5JQ2Ni
8sS+YjiOSdqwBRIoMJ0bJpOuiRJ+tOv2BEba3wCcuFOcSeIiYV7524qSxLhZCfd6
X7iSYxIi6yIjDRgP9Lm+scOku+N4nXsKW5nbgRvaOWTtzjiqikvPJK8t1DmhYZ4u
GhSbO4w5hHHrQu2palzyxRdwaYgHm3WcFLlWrr9xu6/aP2u3O+RhIoasuNZZJDLP
noMEhJyHqopoZe/T1K0rn+WBevxsIz0xjift2Z/CaRGPEXRPEU6QQh1fjl6OJhfq
lgnnzfYxRqpYfYC8BkA0TLaYyfBCGy/sktHpPqk2JjmgEhodVYa+Kctab96+Xr20
8ncT30sk+R43UAEw/9cz7wbS9eKJolHf0k5c2ngcKZIrzXXqlM7E1n0dxOjpNoml
ungRglmxhP/QuPRNJnYKRECkFZD45rqfMApYkcLhiIlA3M4qEuwzWfDOo91F5d65
B7g/zedrild5Ooy2riZp8HFtJrjcVxMCJ/PYhlqcmf0+awqL03VNdaWS6OkNI8si
GuM78pJ5ClcbwQvYMtPjUathBB/KrFhmeVdTzsEWFtH90lMjXkCZz3T9fdWefmIi
acISkLjYbpetPFwzk5IY9Dr/SW3lLAXBM2V5FNgrHZuG7D7zKyA6eCquUye1fSqO
GT2Gl/PCyxp9zLKb7uczlPze9gRLOI3lrKdaJShBarK85z06Cl8W10Rbnr48lY/C
EREGIK4PH4EL4Y5j76AAtMHxI4uhTptY9/hLpgNSU6WzDZ+BmUuCj7J3Ya8jmrTN
P14Ze5XFEYc4EQK7edsMfQF/+HYX4/Qubtk+/ljyhd8UVgoSzrdtqwN292u7Iabp
2UiwaXLBC4jJjywctsNCoxQxFmqrojBnbkrGCw11GjtwoKialkVKlDudsS6oj6gU
EVePSr2EdATPcCZKxATDAfhUdU4DbQFhR5qkVlCUVtPyKpjnykp3TBJRiCzgAvSl
FIRlS5m5oKYoxjces04dZ6KivOkIC+UK0raaoIsgvbYsPtqWpKFXGyLC2xN2r4bx
sNpV1ugHsdrCLXxBpbyT5aOXx5sN6Cyt81OIv5doiAV8NEVzk3DnNNffEBFfeq/k
uum8ILa21TF+lr3XiHMDV0mlGUMTSgVparL6pI1G1wiT3XC/kWtJ9PPSwyIBJbrU
5RV0XKU3mlG2lYAQ4gKcAQTu9BpgmGnznYHHGUvDMsWw1OtALuwF6NQw8ERpSliS
70ao4aFn3b34tL//AHWWVA8kOAOA71u7sqeF5W1e8GDUSdXEQof/Js6ed2GvwcXd
m0E9ROm7YZqVyTtYm/XJ8nEEIAoWcc5U7tLGgQtfvPAkVE6a9GeGY1qGNjA1cvHA
oEKhfwa+tDZDFhmn5Mgc8ToaXaY7QwzxzKp+yjXjGgSRoiHfy5fyXfMdNl5Kr1MC
Tcy+/FltLleDxfDZ+Nyive2GYTNL0doIHEWq/KT/fGEFbM8RFIU4LX9T03+3WodM
wbPOPMETEnzBsSybuYajtDiUZVW0FbMPXTr0g4BFLPqVwimrFkrXABGEbT/QllOC
JB24u66qQQfwfyBZdjUSDKkceHswpAEbkW2M07w/RhpzNgLXX0/2o+FODMnq5uO+
nBR3IfOE+7wp59I7WaUvFLJluavBOlUVWk1K7yIJ2QLR5t6pP/jloK4ahjM0dvMk
cjZwhkd4SuNcKEpZIE31V1H09TsKUCugpCxwpLE2uBt0jqQ6QR9O0NYn/4l8Qr7p
Lz9iaS+M1EsDUOuVcYmTnACnusib/EhneskFgu9+po+35u0eoaIVoHfcSLIPGxKV
YxLzuXgj8XREl56WQ7bU8czwiL7LaP6bW/Eu2mMXC/syri/zQT/B1LVazhJy1pkF
1N7ZbCFaOp+d36HBBKrIicQBNBlbv6oQ872XOS5hkZLDJJM3QWo5VlmnL2Yx8Fwz
2vU9G3T9ppl81oxDJLgKrCs5JPRZPG3luwawlnb5yHxeIPRAwXhc/5QIl/kC+DqE
kPu++UL0zS9KIzg2z/c+c26yrDB/zGgO8bqgAFAAQjJWnY2Dw8TRr7tbDYFt9Ac5
qENQrZxhYauBOs+qGLUAAeHpLuydwIVoR8kEdsNoZAz6VWIFgsxI55U9+Y3i7tfl
prd9Ru5iOxxSsj1MVLbzSltnjzqGJ6AZiaQrgRa38AnONzm6fyOKv9uW94X7V1Fy
Fz/flBq6W196WMj09nhSrCyYxVGZnQ/fUTb1B5FQYxpD6sjhTYq7fbsr3O4F1KcF
HlAxZ4PnCr+PLGzWuKXiddG0RC8yxIu5D74efiwQb8JBNKShWNdsTJrdENGwsAuc
6H6n9UiLQi1xblwfyOYeK5+KarvjBvO9WuC2bumHOHCMmqyMJB5LjD0DqUO6oTok
H1U5iS5x7mJPiAe+QhwBx64Mu3hyDwvzQJnBUtlIa7S056jbj6E7Xdk5gnmbS+pf
xNRXBKFSF0ApCVai9cZrOuOGykzJgJ2VYrRp0pA5vjSOVxgK0cqC+FeDODFxmk/q
U3RS7GW8PlU7Y+RVbqFJ9Ma6q/jHm09piKuUZAyne0px8hA7Nen+AaeSizRfVKAQ
MRwCdeFbUCHjzkdWkddcPUU73xG4sY4uMrneJvsaQVtKakqYR+41Xo57djlEaPBu
V+I3WMA1flQ5/VZk/ZW2kDj8/5YlDckwjtdPN7o0VEqhDGXith4lu5U/7CCAGKlT
Oqk7/AYcvJ6J9wquApBvt0VViLd0dLTPUwWW8tLXLk4Ayah9nZcqzLSFu24a1x7g
pGhDtOHrJwze5HxW0XueXi1WHlCI/CKN+bhwYnAvS21T6YzjWCgYTgeX6T3xMODa
d6fl9Nb5O0Q74bpjxgFTG4396tF1wKdC5lGN72jZgi7SefjFwwc6F6tdfEXiWSfX
6t8qv4Ifgi68ppbnli2BitjvQGglTvQ8wNnAcGyBF9X+9MLe1LHdk7MU4xRk20kl
B5IohGgSqn5SNpqRyjIrbAL9NrRek5FOTlJUF6beZcIdrnNScx01FYpwz9wEp6O8
SL9jKdxynEJz5KLQmIx9oUx/QS4G04jjy3lXfEM/SAG07HuCQ2oTQVZxCBI1ShdP
zxp4cqaKiERikIGTmr9FV0c7DPGkJiPREm+41UqGYJUYt72fRQdBZtBymr/hnVXe
7XjFUPzmvXQ86WqMG9jKIYIL/ky/i71ekINOOdSGJGZIs3/GoTTdzrpRHCtSA/5E
kcyHeBXaSRantogUh6GuMiuGN8biJnAZhvn5WLeUbD5KgOu1KMUyipSlLtQfdSW+
DtsNI/C0cwqedApll9YO2I5UzbGw4HjTBKFe9qmjCLzHxyw+9moaV4QpC08zjgso
OMnDkQZDeaUy8P7SRsV2Zye4VTwgIIQhfiYbTyCRUrDfPHXSwdkWWG+q2o3woF7A
MYRlVDpjA3n6rVZX4ZaK7H3JBuaZLrZpcCF5PmCP5LM3UXpQlAzMGxc4r479wGIn
oMk1ILxZbRPV/Ft5z1VG1CNWqzR7rjyfQUmI5lFAdQzP0vG7gmfAMzlLT+BbRTRV
Lgu+DN4VNcWwf7fKZGffpIFRcxoL+8R/CUZ8pLC/0jb1vyi0jcA63m1L4UYM05ba
ZSVDAdDS7My6dPPztOAQ3WmtPsX9Xtt2AZnIsf8+e0rWPy8ASDkxONSD4vuw4i82
elnUx7pCuX7G3dEvnoxPSR12KNWzMtR0TMQhxkRGNMHzTZSTYIzEpdDDw37uJoQO
Af2BRsd8gGF9rEW4qMQvIaX8nTioAUvtQ/RwyNG2FNJYdv1UmFc0UiS3ynaooTQq
W5BMwrlLKZbQsG5m1oyDZIX5FAQwDii3DwNODnRupdfzCZt8CAAwINvQiJRe8xPw
tIqR+TjTV8Z+DjD0Shn1GZvLq5Eotd5eFPipbQ9P7k12ADf92Kkecv4jYr/MWOof
EWHfza9eGizW19AmvFrcnGltqfhDbALRdJqRpVT/G8VkuJf+WbNdXFo2TtnGkRUl
+EN45DqpA+/AiURKy3nvt4g0fLfKImLLiixeNKx0wHdjzNrH0P2Bqcf8OtfQ7HbC
eTjPKqR41glSyNhf2V4JBv/iVxIthxIgBwL1ao0OKBo5kAZuQ7C5jrkCyZChlsBt
40tQ/yfKKz0zjbzKBHw19TdPKNhnKSSOerU7XxyVIhSTs6LSdxMDGTWAvG8zopxk
8RkbGq5JkwzGtUIA7fZXfYyUowDfN/l2prWfVrMe/EgvPq9XXh/t63GOLB8FW1Ya
zlSAXtzidW99+YcVpTXomu/xJkDpdaMwUboKi4y43OK7eOF1bE8QpKL3jYzcEYGO
ff7PZX+dgsybQBsbf/gGR2jyH/c3eTYGrlX5b+z9aGhbVUvrX/7d+WDa1XZrP1wK
CbgPzBkEBKrp71aW8YMXcZJO9kepp4Mc1K99rPihwhhligloqFkXiFWSOKZfKQZ6
wRpvkU7guDlPaGr3gD/gU2Y4Q58WI6e89LVIfByh2Wjm089GhD4qtd1MdTqoqMCp
4LmXctLOC7Vka7zwWMBigp0pLOIF+ck+LgxIZFLEH2tRVFfekV8jhPJtwltf8wvj
fhaeQW9HqP/TcIhBK3dNOQuZrEH/Rrh20N6dAtviPSLFbFuDLSEwafMTQWetcuHf
`pragma protect end_protected
