// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:29 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
S0xor4dPB2gHCjXEHUHx46z2ZZ3y1o9RwiKYCDP7iia2qYBi8UtI15VAVHF0orHg
m4ficXLinKZNju+V68OT7tEMmO7x6YFGFEG738a0bT/RbqWOopoSJ7da1YVazAzV
llL/C2KRlqZFjzYgKXnH4aw4AL2KQ2Th79Frgkl5wV4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17280)
K+xiKZUuZkwgUqh/CEXc+Zx9weZPKJWjIfFZ7d6t/tTueXEDE0DOCOqhsylkArpv
3Mv/HV7qhgRMHxKPG+lcVKmRKRVhhkQOnZLdmPVweoXHFy/7xQHVj22C2geTAzAI
0ri8F1J54J2wlRmcO+srzvetapvN9rfW9ejezlx3qW0z55FQ/oZLByGBE4s71BAA
HUaD1VulW8OCn1iIdn2/+wYELz5itf9WnJNvyqRn10rWAh5cYAW9FfV7tbZ665Xc
okNYxkAT9F6NZbAFtiDNiKCwyfd09bvdg2uxF0mjR2Ph+z7Cd22WZEfs5mT5pgxi
x4PIkwlN3Dd7SJrCDc48v6XLlMHW8qBYeq8diJfNTMs/cpc5QlKM6yHW89uwB42s
sgnJ1fqdFYDOXcBgwavZqVNjWi+X7cQm7fKnjlmSDocR2fwosAcKFNAdHcNg9wTV
Q7Eblcw7Bc9Whx7iipP9VfU4bvGfKXCvvjs3GQikrc17yt7HKIBSH3HLfFAPRO8k
P8aE7bZFYnBHzTu+VLoGSJ/nsYekgPWiFrZVv2T51ul6mr72sQafs20gLmoLXJ+5
eLqf+KqJvbXpT64mfsffa4olhnEevdmFVfOiTAZT+z9pGps6vwSVNwRldY+QJg+X
wLgUVE4yvvcjwN35+1uBrxPw4oNDJ/YRIiF2mbSBFaLnIxE9hDppHRwCpJZEIMVp
sPqBRJXz2lZAEwlVRXz2iLOiZDoBaGTVwZ6cuqyURnWet9+BAIGgjVGBGjAGmV86
a4Djv3p+jiYK9fFkTOwS6xqbmr4adB9aKx7tEPkrGWgSe28mDBGgwtWeqrJOzUlS
wuyUwPi8m4HCA1T/UAoglgL/ELKJi0uMF4jC6Gr7ER27ZcxOnR9vSu/xZwGvBSrW
AsD+lB2gvvrC0ujlyfTBUFvQmutSXkZp1rt5alOthkRbH2Kur40043ssB0rKgvGS
YVjmnqpsLIzGyCDY1rQF2HB9h+1mWLe7BskgQ2QTDdqfpKQDIXmCMnz/XgjTNwsS
3Zq9UVdMTV6LlRNZI0ivXbXGWVsYEc/LxxlQG+CkOduO/I14DucV7pUMlJ9QeN69
D4DiyhxZ5nQixb7VCmqXMHfdWn5Y/EPmFgavOc511mMAHcUJj3fabtrl3zlNYh3s
Pl9ZSRn+gyGdonJRrZ9dc2tK30HdGVKYvd50QazfHOAowvKSC22tisnu6e3QHFdx
Bd9yZjBV2vv1bsjax+zOXauCqlhJBPEW5fWOKsf0rZKFDBq1wZKfsOqK/wThzAky
X+N3IebRdF6eMHxV4isqyWG0jSm06LCqZ0XiN5mcZrchi4iaAoP9d9pCqrvK4vzQ
72BSJsDgPy2lxHT3alOP563+x0YJ86GOu/Jjv+xI1QfUYJ3eA0AByn/vw7ISFZSz
hQHDOltetoUxeS1vTTU61YqGYyiNWyA3GNEihMI1i0MD5ARgM985gcledzjvJndM
TIgmTv/MK+fm1CGb/sUZnxywaofomAvhlvGmn1POMJSm5wdgctAgHLQHGf8MOcOo
FxEyDOhrOoa5ZattS0SajWJQ332pdwDoVnFePUS2aTJB+dg0/cp52ucmwULsIUmc
p2JPMP+vemkxDweH1VrT2OtFbhMYm7NudUV7pHZjDipYPR0Bqr68skmkFwQ9ctew
9DPHcC3JVQL+si3mTNQIm0rYKzKBXBZY6pmpyr93qx13VDve0I9oouxmv3mapbS2
DlnNsqrrg7I308/YN8aotjm4Lpw8f+rHsbnKTm84ev4ldG9TrQHmLDDCT5T0m5Y0
cftf1vTCOOuWh620I0xJpvrsXnMrW9/jZebpNL4FPW0GHnmBRpYeS6WufemHgmip
sJnE949TTkM/94oveItIh5pRxc3GC6fdMPBvBDDuMq5OoeJcumMz0LwOxmbg4Rbm
qkdpbX5zsGZbsoROr2spGeWJJ1ME+rDwqhG4VAxnfWKQ2M0S0fxuGsE1ItHJaOtH
xm9tb31ZzgXaoaF8ZlMk3SYdQGMSqGv5fUSNsupow82/kFjC3eVSw2pYE4o7BuOj
uWFTH1D5h2yBesgIB95uBDKYNx65eT8DehW9PPbWUGTmmiQaWnwLu3SaT1xX0OxV
duVrZj9wa+KT0iOR18FcS9L3tD0gHFYaPzdcvBGD6P/sdhl48YOyyl5ZC/jUD9XB
asc4SHD9PJAfonXM1jCpGJ4GxScLGRe9VVmxUCHoJaxWeB2zxczBShF/mStdpnZO
azy6FOQJhY5Dqlq6Y3gM/TLwBEcBXbeCJ353o8xU+vqy1r+bF5T0tTsxRgdz/XNj
UwhJ0rzcjMQm1bILq6cw3sApL0Vk0pmNqKVJ40pBEeq13bWs/0+VHSTB6UoniOZF
GKLay5MGjh96w8ciBDbYDRZa/TkVYOD1JpO7hzsP8XDqkkBh+8I4PI+4cwD/de92
1BNiJPyWU2EhzR1DELY/VOw9nnYxhhN9HXTNcA8HKnL1fLi2o1zj2dX/7eJxX6ni
2afOItuvepSDZ6j6vE+wxxyVb+Yv+U86j2tYgPqb/KcxS9ZZ9MBT9JpRNiLKAgeH
9dnirWDQJ5OUGYYGcXSxekYfS4ghbh/i83nQMgtqZVOjZ4meBodmSBB+WuwVvNFp
pPdciMs+NxHZDiybgIpSnW/u62C1dTuXe/WdqpGjACKBMGLrdhShBDW7TlEJiM+y
p8Glf5tqEMATmHnKZ5dkv/TYYelhVN2zCNK/JvXC4xF26yDCjcpdKbydx4w/sHMD
txjaV/9xiK0Ke5fm+MyeFOULlCLIWQ59N39oX9GfxJudzM1hkBkYmQZ5aSr6oo1S
OWO7saL0pvKB6quN1igNJ4BzhuZ7Hep0NX8LimnehwSEmZJVYQVgxPqVl60h0vAy
PmZ0R2ZPS3DVd3/UGz0lT7uYEyRrLXdCm2IzH9thwVzvU+9lWkVVlmcNYcMM5aVy
uTR1772NLL/qeVaPKDJtA/qb5NuQtyZKg92vZjXVWz24M3Wq54KxIq+VrdmVI15i
zcm9Zqz9xT6/pVu7bpFVnddHk5iVMpVucF3Qjm+k+YEnZX515cfaXI779iULzqFq
lpFhJv0DIoHIcpEXvwXXiy7S7iQ0Wo4nLZyVLDaCG9xwsQtMI+FeBw0SD6EmKxJo
Orz4vnGxEy4ihnfl3t9cgiMDpnXMVbZCzRxZAShWqd0B0jawTkXH78UWDZ0DHGNI
XoZ7lc9VTmUNUvodeYmEgjzY5cWmRn2QqA++dxUSE7X+51TKs9pYHcawCZ/nXuzq
L5Ay3aKkrWrFq0NibKXhvuM4ZnUcLfi/ZUIrKLbd8fLzAwZeAFjX1NKss6woqVBy
BbLajK+tcXAUIb8URxHAkFHRk/ZU3Ba9rfuWQHIn7fHE2tvBRGO9de14dmEt4RI5
hyOVx3QXCzdgQzopv86pKWVQf8rBhDW+bqbeAH7iOPbchaDGQp1LSF0wC25hkXav
2lM/TU21HrXhoUqdtx1Xy4k1TubqyFynD/mtFOt2oUcdiOEJPh+Y/S9mANaNvH80
BCqsdXbHN/uXFl0+wh6eUMSdHgtunL/txINPPHdWAEVzZ2EzTRgTkBEQjT9Me1+R
8iHmunl8sBh38dOa/EaYxpomCQYjkEGihmbw8cik/jT+Dlo0Yf4197cs2tmaCDp7
Z1lAtYDUoBCRjgJvCE+kmPMDVWJx24LllUcQ/68LQKmMdo7a/J4pI2H7cj4F85z8
q7LdNoGPoKWJMRkpJ6/AUVQNceaxqMVPwDwNjJB9rqcT4DgGntLc7SgZB87+S2Fp
kU+iTUK7qYGDU28uv35q/PXQfGGhANEE+ljc+Ij6bwYTVGaoHzmWrdfxkmglL8Xb
laIAzhmqa9fu7cA8K8KWOCC236VfHlxEXqEFEjcFJ/FvyP24zUJYkPEy2g4adpJg
UOlbmh9oQbElB28LkD6jwe8vX6kA9Hj4VNwAqbQLhADi69wCKQZQNKutTUsMynNR
rU5VT0jxoRq044A1in1l+xH6ldh6PGF8T2TFtGe05AkPUkC1qGiHJTPiLwpaSau7
bCq+zaFJVYDxPaeOqmSHVi1h+Njv/L9EF22m+j4KM40fFhH9as6vPrwmtDmbifXQ
RtmEQUietdk24L2gqphoCi75KWrYZY4K+AKHv0fY2yI8UfxEUsIY6HKjSpCRV+oR
YMIYq2UzcjuzPbKctxzuL9oQcHvVm81FDzYhNQHOoz2oi/6HVjHsl6WoacGIfVr3
ideDh0jdQWwamSsE25xmQ71hMkr7vschyOBAG6qG6VimTS1JsvlvxSRCItYdTeoi
ETGIYMsJa8HKxkkfOKg3/PsN9ld+PL4xDINlAx5tZuPnR+FqyhU4w+SeiYRJCrXk
pHjvOp+JFfjYOETzh31fXr9TfNCxwFezX7ir5cjkmPe/v4I47gJZCRYfLknW+bUd
Ii1JuSS9kYaeJ1JvFjRz/8qOrHfrzMTPJiii93nCto0LmS7HoVbxQQ6zcFVhDVwO
TvFgrxMtL0vxj9+E8XNFE2pIPrl6ZAkhdKPBA0X5rCQj6gWjEa9HwVFeg3fqNsh2
V0TEsBjpX+XPQ//ZPR+qWmqlv6/MilleUXBZ+efHwSR6zkl4Su/5/PaG0fEgyxGI
du7T/xcc4CYfUOhC9FrXgBqKPJP8KoLVqltvK3DNuzSh0knB/1P6DDMNpY8xCtSp
22AXIKHk4pEv7JOoMGJHEygZsXykhGTC6Dn53+SFbGDsacF2a0aG2jQnKC4Z8O9o
9ADPYELdtJx0TfFMJQYGqb1qAmr+o9IVv1hjdy2c3WJkw2bZMbf23SENRYUFt5t4
GJZvrfdl4Bmcyu1p1h8QoV2lrFyh4g5iBDZajftGVnVwCUAiRNNni9OnkuF/cbHk
SV5cVJEkaDRS+4mU0P5h/40hMHaYS0uxsW8RcewLJMudlCp8v/sIbFPx4DffT96x
et29yMPjpz6FVwA5XdzsaE3izYToxkHBQu/Hi0geeKn7nr6+xvkhGqBrm8K7l8zK
9VXvzed3BqdYIKaiGiAVC+b8Ft5j09dIo/rlZhgFxYIeZqWtbjia/jKLMD5WVM0D
r30uHaZUk1TDyOm5K9rHmKszZ+N4XUJBlGWGOC/S//FwrBVYY1YcOap1GH2eN343
qy7MnIfmd8PGJoJuKYmdH15hMqRFAnVVZ5N4A5Ti3XlRtriIzuhxgPEwNLt+gPiK
/cXd0tY5JbJJKMx3uN82eF3dfri+ZSQN3UkyXY2OInvmTaCX4dL+F1ymsrb35SHT
XRFrSqFMnP4aMETy1F3AVqwK71N9q55SZyfCVlhmJwOZv/vSNVWXGr3tEiIhY5c6
POMvh5bYw89fAPlFCnIpAimr0d10wsTSoXxtZLHuoDB3ikcHoNeshXrylLiyjEML
YrwGpLCWdTYISKE+0+Ixd41VfJUn5WHTdhrSjiDCf4FXkfbKeCLWiJN56Sd3TfXC
g+J2NadQhdrXHl0N6E7VL01edQ1z/2262bgpNUYPvU+Mdw1x+70pCKIL4KVBIEOJ
EMX3XrqBBpPfopgNDU17bHHihg3Hewz4etUtXAESgzbn0PA13HljRFytSk7mXcHG
BHnTEnIEmvFJgmWbqESWHqc+IvJJM91sVcprtoWriXh0tzCieOj23r8kF1S3jZCy
nqwSdCgXFh6QGhHuEnb46gOdHge8HYO5fLCAJvxv7q/SdgzO4IJTEr+pr1dUsxay
aiDSDQJw/lv/F22uYSJAuturc9O6rWcyJklK6jq+QA7/JEUnNAVHsmJpaLWIWCpP
O6IRzgGNZZ57ntetbhhqXSr4WloxmTtC/5EvKkggussLWMhqT8VddMZ6ReWp9hRc
2Id24kGP9D6cc6/ItBmvNxzf7R3mxAbHMy9oYlOcMPylYkceRkQLrlZHJg7N2IdC
DDZvmtg0dNTfvfJskR5NhKjHbttUbsHQm6/PSaf2TT7n0o4xcKOrd5A9pUJ7SKN/
WznFq32J/NBKWcvmEkbVxxWGYUQ8Tc2H2agSDqu2VLM0J0/i+d1JSOokf9qSSiXa
xpDXVTnng7Gy3MM4r2vACudz9xdHXw0P8UY1gNGCwfM4x60QMk/N9d9el9pB/I6F
PgXCsva8IhoYa3os7yP9L58jVjghirS8JoBLkjZ1yAshN6ID2vhNaLGsuuR+4PsC
TL7R6noOBM6LYtTp+kTPNi7GlQschk4Fw32tTPzcOQpyHuT9HjhUMvTHdhQ/jUWd
8+laIK4c/38TQbHvw98rWJJGk8L9oxXsbMAANkwLQbRYjPjBjNm+MaQSh5bhGTbY
ZYA0mGKLWHrHCZDQbH2aZ5hzZgwTsckTRtb/UmX8GVLuGjw8AGQnc/Q9KpSKzlvp
yuXk3+L4uhSaXdDvpigMhJPu+ccPqS3KQcgRRulWqeiO9yp3dpZlSIAmBNe8xW29
P+QiES6ZEimaaQCyLNwec2vDw3bjVcj0DWyuMLO1CrioNGdH5rhS50H0161d8M5f
vXW/9WnMD41/osbiFctAddjAQT0a1PlVK07NR2hnPKb+ZBB8WdzOsBKWGKmnyVWY
rUyrVBHZxqs9b0erMIn0OOSfmqdYYn3BzLxwf5Hlo5N8T/JSRSa0VPCzyrCGa9HJ
aRm8G/rf5Ye7a1Wch3cmEvM1cOF4pzox4/dUCAh1xaaR+MmW3l9BCuwDGMM1aehO
5EbuYM31VdMNQTfXZPVlr+R5IUZ1CCzM/eefObdiUhLuq319tPrVM/cEO7p++7gn
c0kp0hE2gWxwqzrqlnHbbLLO4suDsVFLJog1n4zGaGK5ISAM8idUIx/CGF/3xRCe
cNNnl1Mkgv/xn7ZW082gECZAli/lQqlICapkQw3pngDpF83sHNdBpX8cKhWnL3nF
30v3/pIUWlzqFQyBx3zPNiCOAS1hP9HniFwyBAyyq5EeQIyuEEvvJhWmf32XItiT
7amiKA4KYSxVgfC5m31gKHqDqQFITgArM90Kk0fiU64ONRDimHBcHn4QYAti6cH3
CX55rIxmS7WZUp6lVXO1K7h5r6h/VSKrQkT1nzjjV+gF8BAtOHJEFqcGMf+oOUjF
8Wn2Q2Ybwmgz5ipVX89/vqARe57ShkGZYMMjLfQC7OovYGTHhVGBEUnIAJhNdg2v
FIkdyouX/RDQt14JWuJU6vhujvjW3B4cGnPnCQH1dAur7wMGdSpKBiTz+dfX8jcv
bLIG0bc5hoDkAe2b98rw96U8ALmHsyh3Bqr0d9J5nztCke79X6NsbZMq5aWqYt2Z
6XxGYl/NTD3YK1xb17yluHYzwKzNKGuSlvkXruAhN5nz4i/d11xtwxpzymjUQEzj
szcJsZ72qqyj5W+G8Epc7z3Q948DnstAJo5CkA2ihSsLjbJeDvSG6JMLLrDU4IZO
scT9MeHQtTvIZ+RC+ssS2+FNbEKoqE09ZGIC8YQfwsdTvJCkAkIIlwr8ZeW3CcvK
S4SCCrSPBScWhFwaogaNqT5HbQZtiGp8j30x7x1CEGZWXRjW5Kofu9XrBmv3TaaX
tPJkwPES+pAHz0HUhEkr/yhkWb79nZVjWHK4e33CkGli2Cq374AoCXuzEHY2oI2Q
hNhCT6MIfNngVpccw157EAKbgIFfbOiQ831uxIfvdDP4STRQMMdaapA/fEcEFlXZ
bMyirspwhJE10eT+Tsqc88WQ5EQzgSCN75YK2NfT4Lvic+IgwXGVotNlmiuMaO0U
kTZ6dOCbbrBcwP/tebvUbVU0Ojvwdt1g9FL1u/W2JrJav7/DSXq3h11f4l3Cx+c/
v6pnPCfzqg3GFzwWJrF6TEaA2MzrNZFoZv1WeUmukywspfOUrgPHr8CL9Qa2ZAbP
W5i3lM+LcPjarmN+FdqwbqCNd+0Yb+P2++ldRBs/2ncGD9uNx+nNzgFLlsDuDupL
LzlX0cga5feAmu702HptdCY7yGNr+W81pRB2a47DpMIeRAzOqnBcX5ch+xjY2Uzz
opsVeeVGNSAr9tXez9SmFMeyCGcgy1Z7otc2vdgUyMdzyLRVWmPLZbY6VK/XOfxd
mmEpGrR5FZ73LqC294JcKyojHWsAP9TS8/71wXb5UxtyS+xYSb3XBdneLM2r4a+R
PIUVDns/3aZsN99Lj96iNeWyA3Gg1QW0lItXWa6AhcWRrmkKuxsGQQSsYE3cONlL
QtP1981VSBCab4hSV0QlWJZSZYOOCRsdxYRjb29/ht27VKa0foOR6kMqijmUwDWT
I1azGr1D1LH/t29qSUDQ8hR+7BxUHjK+JilyTQwTxkLSwB1JcpdKIrlpMV/mQY5f
VjKd41vxEEB7WDIaDqpTJayXuC7v1fL76tx+RW0YbwJl+TU2o/9Gt5QtqPWg9Iqb
h4RefUdAKh1LK+K1Kg/NM8TxaCYcZuYUrV2acIE6fgXB5sKkrQTBURX+CRRqQTz4
Oiloqka5jn+YL7YJTE6H6d5eZWLs6jB71TRWQIpwovdRUPNtSXdfbtLzn9zuxjXc
ljbnKxkC7280Iyz/Zm1pUBTngsDVEcIvpl8Hj7WH92UXnGoASFjmf352uoNOtdp4
RIjxGGBsuIsQSrI45KUVeEv5jsEm38haYrVEofNwkGC2wME4X6MfY30BVPF2QIUS
q2EESCFUhiLzleOxTWWi9LlktFL+Kf5O+3iOaRQC3jdTbSoPbzD25gb9m8j+qJW0
1v4Rpwgj3D7TCeJ1JdeujyD6ph7Vl5OTGcMlEs+vjtPthxshLWfqh91/CCEcUNCj
qssXE1L+C0ORQ8ALfz4/s9dswG6M6Xf1flxR5Agm1gjih2JkGHuviFXNIr9wraMe
W97L7mmzfh7lBCxCLgsOw93M6vyDpr9O7jRRC9s4Tfm21xDXvMQtlaGrakFv7YBP
ckBEVLdi18+xNDzqAgaIy+aA767+2UzEcHFoZCy4Dt/GUc8xLYc2h9PzpobiFVe7
ZvdEueK37F5JshPFvKshmROzMuMqyst7+TFNHXXGLdT4b9aj4sSOxaWonHaveaTY
/ijUdloCPq7zrO4HdALLfYVDAuEAdAuzT2CtwKRCM/nGx3kuzHGbPjBTmQbKbFN9
1x3puuwP2ebF3c6sHuudBfX+iHW4SqRp12qTgW3lP6/bM5oMJAXw+yDb1xREA3Pa
D+uUowwIjUQLzZS1yhcKR23NpqWgDsf5rECrAWr+iuYpX0Y5YlWVokUF0k4/UgRo
CNTYwYH9O+HkMavbyA1KgXBFbu+YY8uXZRSci9vDvhUNhELEqPnVGam2YsL8/eUD
+oUU9k2o2mNkhSK+ZbOYaoEQfJHpWHJtVlW+5bXHdCuGHIIXgCPsdzTraI10Lkhm
L8NqrJOR9devMWSt0nM00OnzPTKb8gCQmLySE5n3ir6BBpQz0wLOqyEENq8wld0u
GwhEcpGCb5qRh5vMMFpAMKjwl/7zxDosAm8wpVvIrN9dhZ0hqkgboFdjLryd9Mo/
pYPttrYYFvR24jVaSzgjI1T1e2pIAynadDthlcv/oMXlSEicISgEOgCU2v0LfDva
NEbJ7QQHXD/eGogymYQ25wBOFA3IDXuf2FdD/QERpypmERNbzXFTdvZv4fpy9y1b
AcrTAkJxiGV+HujXIbjG0Y6/8iMiEnKZiC5Ahon9y6gsZR72gYlf113lGbq3T2PG
zk751bKtNolLo3RYpstr7w7wtq7R0xeDCgy4m1FNpI8oDMRJezbE/MFu+wK8cxpP
t2jQzJCJYACVk/OHzNsVMXTI+2q1Aypx2sDVoG/OtxJTW3IJxa/1h+FJVWWwY8t1
t96UmeL0lXgu2kBJWyYLJXzZcRILrzcf91A7EiNOewpsLNb9OWJTnnyjYwWz2yI0
mKECKYojRD/rbpxF2Rw9B0NDTBYHbFMjDpaVMgmk6hvswAdT0QgYb5XA0k/jCWiM
E9j8cnxavxhduuMD5gX3WnoZsldVFDJCTYzYsSqWOpvn8MyUGquj45Ttk58s9paV
oZEpTOOms7NkUreE8t1K5Wk9ScN4O3yDijb3Cwq6+g+9CiCX6FfA3q/F7F8BiI2Y
rDQJa0769HP3HjL5we7YokqPcia6zRtrvP8kE6Q/lkDlia3oF+6NlJPpr/l1SOv9
aK4flza8fXbpN81EF/KLe8Kh4o36oUXWAZXCyJyLknEMNjZk+GfUoVEu0MZrtO4X
wFwbZRXNdsgl/UbWhgx4bdZ0ZUKphxkt5y1EcC0mHoy6RW/beFJH87EY7X8YwTmh
lh2L8VpF/g+7jBM1WHxMGKNQuBEeSCSPzkKKpqjcr6VZ32HWPYn/37j2K0bik1oj
mqgHBujH4vzznxAYnroY0cJH/8DTdBALQi5+dnCSmc0HJxPJYjV0i7D6l3Ee6nre
fyIZXmMN0oeAprxgSGTBitsUEqXQBO0MuuVSaYj6v06cjk4JpV/ohERRKGI9rxZA
My0NicypClN++xMzcYoB2q2dGchY9QNJxr1DVM3zZgSaXV2tDSSPgwp9XT6xxkQH
xxUF3Ab+4Rv2uPnPWjXas4UKI2Xi1MSM3+2Ls7c6Rv8xu6D2uOW8d7/aLhTnGkDQ
c7zLB1NC9tn3R6W1gy/qG8/6i4I2UxLkEolPPCYeA7LSQ9s4O6li36/yi8E9mZpg
Y2OB/Xq4PO2FrTl3cffP69zAiJ3VdzfchHMg0zBj5s5VkP6jiRZAGakSZFqNN9PP
mr1A6kzgo7u1Uh33Djmlm7GT8ht996eIWQwvXz5gChmQwLPZ5N/yUaABUO3kNSIK
76+HZf/iy1Wm9ADmikR+gtSD3AhmbIRErBszhNO7T97aDPYQImBGiOOC4GneNE99
7NXu4OD2GLpFFbo1nF1ZDx+v04WxjZadWkUKzEdPNx9R/BfblLC7J+lJxnPQIOD+
TSemFY7c9EdHQIgUMaDeGe1F4qw8iSRhyX1aXzk/vpM1f/j6alBvpxkUedBoW7Cl
vQ4dSvqmVXYB5L5YDxv115NK+gz4lWQQazp5kaSkUlwuVOyeQVesWSsfThKk5LJ4
S19/ci0PyzHoZsOp/cr+cpnsNlvwjsGGleP9fpq/uN2kbvy3zLb56NzWEioyXQhe
YSWYzeBplh0oKk034ejCOHpWvD7njUNlWoSve0nEzYyyXT+MNlfhGi2cTYzvNBzg
YAoNRD90hf2WfXnfQPAoKhtGwoteCTpD6En8zEDG+fz4zk1LXnf/+rzKL8SaRLsr
MQPywAryRyXURpfEbavv/hmEu3JaPUfeJ03gVSY0eo1ZeupXkhJPDZjjJJ8xvVNw
r5iqrGWu8aOlVMHGWvewoTDIf+zuGbhfbcMBXKWvGnvya8lOzjwgBImWqueudjim
6GPrBxvfyLOar1aaXKy5m+k7qP8BWeqZ3EjvEnwDTQMLtPqfQdCQHJNm0D0McZmP
alhg7GwlAJ8Z96YO7R9MOICzfqlgryDObDBEJGYseL8XH0FA5gnuKamFb8vtJsjX
eJnrxhpU8s5Ps5ZQdtUP6HPGJPjgyji+j7oZnpq0vtbueTwFsbzhHmD0z56Nqc8E
RIJQFQa6jIMwMFB8VDa/APvJO+wxvUJWbDV6d4buhc0l5eZMVHNJV3SbgNG5iBsi
nOoz4jMmiz8KX0J0gOiidFi5aj5Y8VM8zBIlQPOwLGyfcxp04pvRPMQQ5+D6H406
K4knSQx/JdXG+1BcskoICxJ8iRMfdyIGk18Sj5gNO5lmwTgjUQcfYuWP4j9UYL9t
Ceu9gyoDGD2duTRZBPqhrjsU88kZ5qJgFvXn0lRnUFa2xfqiigVHWCvF8RUqKmyU
6MKKf+kSj+A3BQW+dFg/PFZledkHN6UTBhxrMa/SOi4uj0ZDAAuNulsiJpPMBD62
aT9h/YAVh6lwRLQUTNtE2/wFJvsmiHazLa8PffZsMhMQ1F/bSzMBI62DWM1jbqMP
XVPf6t7NVmBwvCuUMfOAXnSn8szNsKo+j1Aw9vFzNqYnmqUhGV7eeURt/hbYrxBZ
+cvXc2p+AIv6VbPJk6ts4YC1vLKB+eP9ExCo0MIPro4m9il/sk5cbSC/wvjfw9d8
UGZ4D/047usfyKL5/6r2gfuOSH2oCnJ97NMfsljSA3PWY8CIug6+jHN93u+xh1Zl
3BJJt1aYYrIoxHuu8br81aVTYXTnK+sQ4BqVIShCvbuP3VZOc3Sf50me4PzV56dz
XgI41WRjrOczHck9Kyhdk7eC+KyDj9VndARTu3AL2ViQg+TXLmykcbufQJ0O/XgL
e/pzHb+lAvx0EYWbdVTx6ztG0Ukz6HGkwkarhlGD1hx2r/3glhCvqT3tgB5DMh92
KS7ss/BcxnrSSZfurYq4tmbbox5CuTveQN+SFUbQ/8ZzLLXIOc4xwBFG9gCRa5Hb
PV0DGDnXa0w8xJpb02GtfpASi8GkJ8bFgQpz5GvaBqDypHLF27XYFEtx0JT6wkoq
mop7QvwvEXwek7Gp3wsrsJ5Hk528QG0AtED3sAf6bEt3/az8HfAs6Z73jozIm6mW
nGx9xoJYpgOElGnZpEom1jD8fpXAzHDoxyK0MXtUu9nbYt07UvMEtWwi3IfjY70K
O8HGnGBGGG5BDrgZcG3x4PlJkOB1yhT5UUD6zixTYMaWIlOy336+2IecypD1VPl7
RnSedhpTBzwAkrnCrURGr5bNUack/F74PUoR5whOFV/dQPAcrIAjrdd947Zf3dTi
zjGm2Yr25YOjlHHJO+S+aZ+W2fEp8/c9nJqLgX2Iy2dsVNggYNfqMvJJKiBRb4p5
cOtrflMuiyP4Up25lOZC4Dmn1V9NSMAcdC/Lmc4qeGkThT0p7L4fcQbhJJKxQpic
AHb32qngQznsP/drhFTdYPDyvMICRYtjNgKqfv/U5R11QbBsPd+o36Iesx6k3SC/
8ryuOFz7n7hqEFKb+e5CTnDBjJUi6ifyjBeeFuNbaKDKntnNS7u1aVnrPJeQBtxA
CQOfqA2gNFnnrJAxdBxN3eopoqzwaqykgME8KA+HR58VsVTHUd4AqlhvuskElr7G
5eCRkisypFLWh6o+fOn1RInaxYBONZPs1P1MIwtbI/ycWIMMEVUfSt/eGlsZ+qpO
vOJ99XyPICZp+CvhGsEuM3EQWfA0VOjABJBg9EJvRqG9iXSi3gj3ues1znlTEtRM
HnCzx7me5dunK1C9PEmigfZ5r/9OobhpdqmDmPKFdHOM6zraGMxfvH9cJmgz5APO
dU6ij2XlYFxvqX02QHdn0kAUwG0hru+renQEXMXt00ZKipv4Bbrixq46LhqZu6Eu
OsT1u/+aJGCeWaXuVztjpzE17rKqIZJifEHmvGpS56JswyyPuFNhU7KLZs6bJJ30
8onRh8aUVdiJfH4wNIc0oIyIQqSYoz2b5dOVWdQgFbNRa2MtMqSFEHSQTk3Xk0SJ
gEmcRWo98h5uSF6TPWBd4H2XQyr9rWXnBrJ19fkcGgP1NC6o20lprV9X4ltnYXy/
Ncv3vgGj6ARvxRBUnnDk/krftj9z+yNpdio2SRe/2vYxLefU5DKWqlmXpoSoG4Ba
7XREm4a5IXrzdOmbDWVxeks8FxtH6W1KOMNEAK6rucp6GXZX+71zRD/fEwiUnYI4
eSIvFdoIgC2sjXR6AHHkazt7kvf+33ffHjH2dE6AEfZ12ld4uA6kj/NlXe7tORM6
14O15SN+mrRX/LMKF8PnxAi5LJ4u+e0TZhRHAIHQ9glJD+xCPSfonKQIwrROIsax
uFmRuYWjqRcnPHJ9whOT5S28+e1fmOUUxwhrOna/nd0lG/JyQIYv+FDXGDU6kBCt
MJJAOpDH/sLFPrNlkvxdJUXst38KTFIxqP+kf31ct+yx8fPzqlLxwmXd8HUHqvZt
DMScJwanB6Y6rVwl2PrBYe0KA9aTnvuP6YZiNhTekPeKJ+cLx/yDsYhMSSEUcysc
/UdwnT/EEJ8Z+cHrJIoUxZaDDIUrMeeBDHcbZNK51VY5X8NSQBXC0DaKqIszbROS
mzI8qnvpoK/UDFyOOp9sdf6/YtvqaLEEhCc5pB/RQ7OdJ3gmN4hKv/iorbkV/iqD
pJbGwQlgMYvNJWJ309fGj5towNXzLezJ6+VMs5OLOQi36GkNoyExeKmnyE/qLR0T
MEUvo2N8781AL3F/aSgIwb/E4JHRRMWqJap54HLhEVjQUXxurtyZn2LSbAtUFRAS
L3baAmYcTM6t/4e3hThR2BnwwhWUb5MfU2gDmRJ2phBtw6GvDNVt4lyiynjPuWOx
u8kHO239kdfxWDPwYglYI8sXJFXzIKwXGkF8VhfazlzPcy1FYgAQ6JPbMOKpM2IV
BG4qmmvAT90JysSZ12hB4S9XJ1W+5QRdM8wjX3SrIkL26cumr6RAeh7mgeI1R856
gyplvyA5kdyHpaKgzbcCZctudYcfjRKXR2W2cmXdMYIj16CTDNfJ7MQuNTFzbRms
YKChw0XJB9aucoDt/XrnXrBenJlwyoQJbWK7W5v3eY+s9F+LdVoNy0CTUK8A+CWY
1r2Fey1Lw0A0Qceq+0bEikGQozIppKGMz6jsnCac6K0CGg0qO7Ewl2BVwmz/RsTl
cQAW880yOukF/VOvfI/WlorQ+IrOwAxym/ujXjy4n/EnjmYFtreeyALMSySx6ygF
HUsNju4Aa+dQr66l7iSafJf4FvkhHZSPPnnL5gYuWF9RvCHf8FXp+1Pb5ShMcozJ
cH/N0iq2SYgJVXwuDrmX6l8IzjOGPZQOC0zg26hYRTK+GjL8SLePCAQvAuxLAyP+
JBYjZzeuZSziLf9NVQdiDKJZUwIZkaM06cAv0+OU9BaL4Oa074htmuAI2epqtLHC
Rt4ukxrl03vmVnXbj29iYFziPU0rkKJVOAHCN9ZV1BR9R8BI0/+frlJ1r9QFWyV7
HHstUJRoP02ShDcxNcnKdVhfQxnyLUEL1N4FO2vmPYyyhSmZvCiwBWlEuMl67pF5
y4rbgtewcU5iOX9siNu0Kqe5dJqEB6g9Tb6qyodpxHDtYcMOrjj8nJxCdWLpTSiH
ki6hUirTWft/H9nuNovxOzOl8bBvDUWPlagpZhTdUEIZNpZtelzj7motznCw9JSw
Zm1yP1CGEl2hu7vNYn2wqLgBI1FB6pKhcsC4UtJeAU8QKnSj/+M6bg8NIxp6TOUK
/hKL48vi/c+Fl6ig0w5fo8SnlSOFBsGqAViw8uAjfpMmM4TDGkNZj/RP1mkbzSJK
9PQLa5XyjXncxk23wujLaeIny4G2RKZ7R27ubi4aZpLng120UBwmDGh8BTChdLhW
nMVlyb3RJOap5SN8oDBsFBuWQx7Iq1NGfPsvt8km4hz3uha0G8ufPgaUIlLB9NaO
pLFp+gmFtIUnJvOzIgRcbkTZnkanD5GM+PKDdpn+1mXHFDYtXid3KuKN+BVrRhAC
TINAT80BOdbV9g2ZLnNpOFHbRDvXYjQYKiY4dKEzAR7ylE7gk66NWrX+pGijygvt
5ujGUev0Lk7GpYwYuROPRZMoPvCYYnVYZcOd+/AEbOQ3Vd8VrLP5VzEBlGj0Ug7H
k99i4tdRiuNXKtsW7EbCBkusUnUHN5Fx6/gSu7vM7kEuwfqcoF4IIMlnVex5hp4u
4ZTmMXeFoZTUcXFkvBLoJWRTbUDVcvjpZvb/y74CxNcu1NE9mfMFrxI8ZFctdHXr
lAQCmeCmkiSGfbEDYkF0/Yyv9jT//NWbxbUEZnTTHinggGU6cnFXv/IiBGWcroCi
M0FYclS5SXwBP+NyCAQPqPGld76ieADdLjCXEjqod8+7MFN22i1GmL9i3a2fS2kK
GwdhesqDuDVbvyGSVoO7OHfz4enJpxml5LZyijUdlgvwL0miIB0bKneF5RnW7Y5L
SNjLwSIfdk3L5EVkvFfnw2DP30E6vmLTlWQgwPSDpss2OhkoL0eMXZDrkaxL2bgO
zaQdYAMMEvUtB0e2K6hwnU6w9TTItLqSYvfAzQPwrm0eFN9cT4qzupdOFh8Ell7I
2a7U7I/WskC0j5izvvEdd0XIDS1tslIDIS/n3rP8jKPleyGGL+jmU/exiR6P9Gu2
sikg5J080tX2NnbvBMtIWjH5juUMvklVMPTz1TYV5/a4aWZLFMYkk1pxt4XjH7E4
7EOcvTnv+1jz/aljf0R3u47RrPbpPLcRmBDLMxERXhVSc3pSG5fbR5UELTYxQe+3
psbeMxgXBUan5Ao8ClWRjuW390an/TqMQmLzXAa6snxgnqVKUek2w3P+NHww/GKv
+Gg9DuNrRb/02wU/dzNsVC6Pq1+6jBvAyyLzIqmITFkT7X70P6RP98qRS5WpK3V5
em+GDP7e3OWRD0ylJ932i2xuc9o7e1+nFjslMpzH629DyjJxefqEh5Vjqqj+xIgP
JgwPGEmzglPe1tDJLjgjmN7pLXL9mExOsLcnwY3x6DtN4PYaVgK+YfDE4WUEOML1
Th65ncnWp/Kugx2ZP6eMCFvWJGQVbLTGb7hdGJubtmyhIBj7euAlg3yi74NaPri5
IWIz5anNi28F6/PPuSD0ml8VBfDbw0wsnD/S5YxXkjb+nKS0qTJW79oCzjG/318v
oqxdZ2SpM6je8Jikl40ekoGVa/3ogY6hxi0qzNSpOSY8cYYJ7LHMjgBvkX7FnKkF
ek/OcXp5xcTqKJe3LgEEQgAPADzjZgOfnyPnhPj+eChxvGR22mjuI2GGNy1BbTyP
wcwCO/mU0oHtxQczYnYe065RHW7jdld/xuVWg8+MyCVp5ftLzqwh/MdVGBq5h+P/
rogqALIvlRzBLs2Jg4/YqRNRWM4LOg2gNqrDh0E/OtgqsTJ1xNN1v0calulh2V0I
X4PRw5muf11rzux8RssKZo5R1uvL1wWQMFi3h9B0Ggl4wVrv+cEQ69QmlGG2UofV
K4DLYKG9J2jgJ6q47DYKVqlDIrtZt5QVS0zj1cVc3hx4JhWfnMxowA2QnxELcfg7
ZFny1spJdW6NQmt+dC3pzommdtfOOFLuKArlbm6/AClhfO9l22zw5nxfFCC1pIE/
AqM+Hq324qlEyf3iF0zQ849W1eEkVI1bmG+rKFbCte9eNd1RgC20q/LAqH1tJfwH
PDaDPduCYZeUlBz8TNLQe0EhBkipotGDDbg9ajkZSFg55E73ZL31p81a5M5NInnl
TsHnrNSUWvBRBjtTeBdA9chT4xIkQoNJUfYYJQxAMLCEAXxL6C+jqNeY+p5H7UQa
Q4stLyJyPt2JxIoq4pOJrVIZqrVk2elEB4yMHlSD8BI6ycHIuEjCwWeQJTudYLP6
nwEbxEEiP1K4oZuPj51uFCJekhm0IQoxF1bimEumvobYWGVBSeS9+snczOVCzb2g
MCPgfuYTK5TMS84QqzxP3H+f2a7b6pVfqAsdFMeTlSpjpRGyQCkDkK6BPL4lIGJx
XnFFYjz4uuN21GQJRKuV9OS4Zu+jELWZET0LJAjHdM3CvCMyGJF6ZxcRMLHyqB7Z
3xjv8b9Hm8RWDMo0hS3fHxhEk/y0qWIxwS6FAAZOfSHXJ+3sj79HkzPzgoaUWeKR
laJ8RllLooC1J0VEh4mJYm72voRA+KjNV2X0W7lpXsMwZeFOu4vNavlh/Sdzw8dv
/VUjK2ni40lTcfymL5dwFebcTL3PiQeuMozFZwoKecB91KcH/E85jgXz/D4eqXfi
qQXTUp4llGYAsOJptx17silKnTw2H8LurSaAcBJUTUVW2ljqjT7ieLFEUDQKRzUA
BFp+uQeVar2Mi1++y4wCc89g+HBlQAxeahj5ZPrFoCGkmBTen5URRTwyXA6zKfuu
OsmghrJDID5J1McP85k+Bywdzyc3JSsxytsVCA4WPG52H4QF3t9911iIMWTPrZlb
QUqmfiYt8QracfDV7qw8U9B8Kem/bMWB5uUhhDJO/YXYwVdql8wRpbmXC427jBti
WErXXmDff5L8otlbuas+X2MmovrMUGoV1Cm2DfahjmFlZmS5WhmeBRfLxFfz5xfY
hbOwWeC9+gBs5Wf02tvRNTPHo7DiOeypT8CXWpvtW6y03v/cJKrC3l8/ydvW5Yve
qg3INre3sxyLH7RG6RpYhzoXbFZImNpHWlTKGB2V3CcyYOMkVyEIzeQgQCiJ6KJW
yCnRKpiQyZU2TAzEP76DXE4jvS97kZcNYdqmgitJ048Tav6ccoTt7nZp7obzo3XK
0iNZ2NpabX6RtAfNZCacwaf9WVE4bAqOrMGF8rN58OULnOoN9yDNkGoReiWQChwn
veAYQWGOXNypnW3xLiZ39o1phV0oQjLXFBspzyskLGVmAP1kvqBlfp0M04uQch/C
8mlNSL7yOxfwjckbRKheWDmIb4p3FVe+hPq4eKuFNK50eqjtdyVWsDrfp7ezoNv4
bT+02hszy1eLD0V0dxMGjtJ2sjaqyhkhdISD84p7zxeDvD0KSrFvUyHbgvEyX7KK
jMC9hoCZXfWK6aGdDBWig8PiuMKoHbUKHertFCL8DgZDMmwVviRyOTKUfpqtdmyi
2FBUTCZoZ7I0LvQR13QlSbIinHk96qxzXTtZN2RNbe7xyxhNr8k0q7g5ZXTfGcUB
6G54sw+d9ie8Twwkdfrnq22vrYYE/7gnN4SJXCATr1zo7IUIih7gTdlUy1oxR0Sh
qqv08hbzNL8foG8FSqyG0OYSgTIOFZbshg9BMqtCJ7K8OJ287RNBbwJEYTlgOkDs
yffrX9A9UXlF0uilYJyJHvWJOVk2J+wILWbqy6MQCSSoru3eDk3VBhmsVFr6+xIu
ZY/YMtFtnAWknRK6sebARaTEiBvnC9Fs3CUBLFGVJ+QAc1y9ubEdxi9hPDnXJapM
+iL31z63yBQb9LRQOlyuwSk9cgBY7u/x4d5QWOrBVIq/nsOPhENzqztfla208FSo
R/Wm5hemf9ERj9oUHEL9rteDDVpk3xEAQTIeEHAEpiTzEj7GnHUkpBLmkSOXrNuF
KO+UWiyrMBmJ0SxMe7uA4MX5JscBEWc0xPm9u3t/c9jqQ+UcpqQhV/PPQRedkyeK
kiPCVgTu6ah50EmbAcgMRtYnOVjWNUBGsyii4EQ/6ukhWvu6ze8qTGJmTLWvgo5d
9ELwsQO9awLoejDFJy1PUlD2SaTe5hXservphBzJz76e1QGqyf5gJ+k3uSM7vWMU
698WTdbAu7pmuZZh45r17TsDVBhfwi97sZ5SNxVKCd3dNvsON+6rlN7YoO6mecC6
hPE+xCTTUhZPY6/8uofee94Hrqu+C7YacHfaiLSvdfzsIrVxcjs3+7Yzot29pKnb
FrQBzuvcnfUSe1HVhkLF2s6JcFVpcM8WP58Z4Dhhvs5NjIaHoVOfyo8L7IvieTkj
ryDVhCY/QHB2yPskjfWubrEaQe5s2WPBS/ZRl+jIeWs3mNZqP0A1+eakSFWE2ePy
6eBxmX/t+GtmmXrGkx+v6OGZHFjKJWMEeHKM07MK07qPUCy5j35Y1JQ+EuwBID/5
l/mDCbAv0jQNmVfat2UabBpR12j+VE7qpXQgnfDQU8KmWjzAN25vnuLxDFby39hE
aRO8B35BU7+8IXUMA18VVBQ3MvFuDLpH7MjYoEyx+kC6fm0O9NI2xElzYa92uWaW
WwjM+2PR7x547Qt7Po4vo4+N6W4nkyeQEL+JyUFg5Uy8r3V5mwlAGWgW/6bMj0wN
3QHhgDpY7vTUyyX9/kMLjl+OndVk0tnxp6QQdJgqTbqw7Zwsqos7CHl11SRUpZe+
yuKLxQmqqd7vjlDDiya93SVIqyN7/jO7ZZmWmU5Z1/OeblS7cKugUH4sDr5hGOW8
eDOAQqe++vsgD3TwLLT16TRIItZanRWwfRDwsL2z8uZ9g68sRZf4jAFpzBLDH2WV
eFl62IDXE1Dcgh2pY/zOy2CBklJMqVlNZykhvSNXMOKRKmS3zYbvyH4Z98noXtma
RSNcl6MQekj7STnTRO9J3l0hWG0AaUMfeJXsX3Y3NIZirrGeaOZasyzxiH2ABLLe
7Wbrm0DMymh4t1YcjFSjbJbeoBqDG7v7lKRk0VbCYopGqyzd3qNp7Nt7Br+KPyCL
AH95uhfxu/yegRzVz/RDwFh8RSI7KHMZYX3bnt7qTSKDMFMkWyai3b1b5f8QRiVD
mL6tLk3TJ21XiukIh8ttuwaeQt2nrRvIHOuqIDju876AZrwgyU5b4wdOMbgMT+pl
urBNfe3/fI/2FX+Dal2D3ANh0En14I5MstTmMqthni1MBnu/FdcwmNMzm5+ka9bt
HqVuJlmR9LCMfr8+9WfJvFKopu5FzXKsqvnE0vzt5R9tWvp9NrPqXDr0EqpwAE1J
7v5qrRyDnox8rPJTPt8eZA3qyD3z7npV3S7a2aiUpD3u3/D3hwApZzQEJLWn6L0E
fA4t4mWKaFhBBft1HMIjEraKXHKodvSNe7Ehi0xnxn+DOSe+C4hG8DfoJi1zWlk4
zxDPkuUlmrPiNsZVTjhxixe76Ifl8e4Tj2kuJ0Fj/O8PBe7Ps+J2QvW8Z1UuNc4g
INX6QWwxQSwqpxfVnE6bXN2/8glNuycp3ErNlxaBHI/ZX6Qemv6RV5NHLICqTN8I
ARmvNWt8UMI4mFnYbfNksxxhWnsfc2geQbGA98tcZPvPuPVTmYYmOG8ln+G+F98n
FQbDSKBkZjY81VWT+4pnFO1251BLfZa8pDcqAAq4lyAOTlUx+a281SgQkKd+940x
6RAV4sVIwRezRBNAdXreWbNHGhoNvKkq3Dv2ai0AuOLBnzlvPclcqOK90xN8ayem
ODwmwuMhdEKrgTQcor5W2HlK/gdRyffatYjKllNrgHh9WOWopj6W3F7exx5+ELgj
GfF54U76cnTrbpsGHTuQTpf+fuxtesBUlDpzsKWLql1pcp22v2eeE9xbAOmsv3jE
aOiEiUqci8y1CRhUURs3ICZe/0fIllkmR9R/atffuuza+ZcuVeIwMSmxKRef9qpO
BGRwjcwVbZPC9RrOVmg1sC6CVvEPnlE5ELxrCvil71ueXavXKfuPIPQLDQulvS8j
zb4+aj66mZCDPSrvGhgf1LptOl+jzzLD7h4MiTbOJ+Brh1styMQ79eAGMVzKc9x2
SphJc3DmVaTuonIghe1xcFNIAx1v02ELq+QPLwgxHURhkwUzOEhzzdPJnmhptfmJ
clGSfnrcqtf8srNH4PFOu0RLsVLBhAWaBMYH8HtUqlxWIpuf7N2R7VcXUYOaioJj
g6Uo7rezAwySEeNrDjRxXsxCkL6v1Et/j0P4WTY0SxNNySs0n+bp0uuTdG31K++x
P+wQN0+dd8Ipf6e3NXW/2Ux+6u4EGHC6HOWIyPIKSxXcl8hE2S1P9nqryWRmpcix
JjapqlkgMVyXTEw5CP1srU8eGKRcJX21k5DRikRRdLY6ed5zjvgvP/+Xy9sleYHm
ypX7ctN4Ts9V9XgJM50UCx3y5Xy/sVaiIMs+oLRD9n6+QP4NYcNKMlTkiZXzbVX1
BoZjDhipv97+UY32Nw3c693w3GmhavK+MNghpO7advFaMrXBVkMqpDcEmyleylkx
wPXuirJNAPMY7JTwH0yRLYT7+PoT9in+c3Zg2vXaz6Fq7g9PNTNpMeJKI3jXw41x
6YoAPc2UliFe6UuV5Nbvn+3Sv1oDcszi4c4hJL06rr3YA7MeQd19gTCJdxANxgvB
Yq4sVEoTGHonlOUTdBeXVD+FF+LsOIGkjfBZSQgm2mJM5ttqYi7lQeWcYFf4+4su
auEum71hdXdIwTZ5lv1qwENd6shL4VWtUSPM39pRd05dlUGLtIq+kjknIe13XFn9
Ph/872VV3zmsgCHD0qqCygYrM5cjm97O4lut0YmW19Rgf9bgZ9lE9KFJ/lwd3SHf
1Eu08U0AxguM/IAPECwkYsjbLe7ytqPVdyvuZ/q2TmTGwxi+c05GGrfMU1ESif6K
pFW4vk7afufoacxgE7Yfnfhe2NHaFBrl7dBU5Dqh+9evNKOKPj7hgUAPawlByqU2
xqYeC2aI+4XMtMhcA5D5Lh0tydS5pWxtYegZc89XxFUZbclYYswyChWTqgp0FwHc
Fmz52J4wlOWds52l73XwZZAbsFT/INEuvlS+hV3iP1oGwXFIRpmfbrre0+7m4qU+
Ee0HnpV6XFkxIQead7ItzmH+EIEBlFZoMROXICek9GxIo52fp3roamWqDegpNW5B
lQjBEUdRrOx4ckTTIbXQsVh8dpqcrjkQtxndKborFbtsWlACUlrdjW4peBnUy7vx
P8vG13tdkAmdsSB3JxoHHBcQ5fASVbK+v6962e1m4df+HLy329x2YevjBw85yQ5C
pN9f/3VPDs1wXS6tlz2mWiibsvwVVGkqzN81Ts0jTci/EzrE1jggxm47jRh0sBlX
xSL55tjPnliaVzppxVzmDVePAb95RHnQlKMs05r9eVDNp2mSmd+2H1LiYw/0s3yl
2pvqctyflaLei9xlUWvJkY3Rdy3JUhcPalsL71xVxs5B0WJEnqmYKsA619lNMjnA
6bilVgLM/QqarGUkZ2iX8FEGHs6OSSeKGbixU8ETiKLoo2K4veq+BKFXl86pBVsE
0cCaHl4uFWBUDvwzw6TYRIlb+sgLQZa8pYwg0zQ0huaTJstxqE2lNMoKJElXUrKU
UDgNoeMlfnIMqgamCiFjrgMlxrSI2Dm78BhLC4kzxdDqjwTjj7vIDe8mCw2lu0Wi
kpQ8pBMrpvvXzPA0uAuzRzQOqL5BFWvve1jmq15RNeVhZbhhdpQx45mlqXM/N00R
bhv7hpYw2Cp5MVa6ksoxVl22i3e17FizmA3eYfA7b4d+5e5y1VyNh8b5+l9YG2Z4
BGo5o2xY7VRXRavazQyba4ePrYVIu65oD3HjAdkakKKx2EuPO23W2fdsti4xh/KJ
pl4IMBM5CcCr4xDsrFTnHT8YHgVqJhsbh688Pi2UGVPGJnycdyXignDfsicyWv/D
SuTNWv/52q/lxORo+pdbCRUSlVzQiR4HgvAPYJ0/tAbaJWjSS5534j5C8zDkaR2x
7N0W7ron0gVSafNR2V4tXCitM/wDPC3mJjC0SP5k0CIn08x3iKskWd+3d89CBU10
TUEphOHfpMXfCNwBX3aFUnb7oUl5bZXeVkkyBrwE6agPMcsiBNOctCNnxB/TV7w6
nFgI1+XwlUA6W5xwH707C6HUekRrafiy9ViH3/EsYUk4SPp9JUSWxMmLdm62P7o8
`pragma protect end_protected
