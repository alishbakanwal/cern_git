// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:32 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
smbzoloivWcA4pq/5ip9D7Fw0ej4ntIIPkVmPr3WzzOIzZUeCGkDsLGicJVFWBxD
3RfBZjweOy4vko7kUm1N7M3CZSvvf/M53DXD7Ec1FoEikjAT4etj+JZcFeq6jcOl
8jk2wFmx39ADxmvqtk36SqYBWr19+eu4b1Fhvgu+3b0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2836896)
usF9Q3wvlTyzm9Wk9GVhCU+yXHLSj1MncsiWrboDcgqnCxICQYQBLvUH8va47o83
Zbwk1hC6pz5j3NFM5jGB56tEe2KtVGdR+hoMmhgvZ8+z5heWVE5YgZcZk2Kf8TrF
eKlUc1irrZs5U0SlIqcAHtvEL0U+/407csc+rQ7RFx66r9kKQNNp8GXYv7O8e/bB
zj62UXIJDq7JkKXYVZMtb7M6g0/zuR1KH3JaYM1ElAfRYcojGqHt3xvm4B98fI/4
vyVanKv1hlVnpIxGNtl9oU/g+LE0AkApONNNKqnG+ur4JLhEq43ihOfC9KfzNrkY
227GeLa97yfdRgAif/P4C6RLbKBc6Tb5YtlknhIU9IITNb8X7GkpITPDXRllTea1
luf6Up1EhnEsbLApFx3QY8+jOfCIFy4HhOZZTMERXH8VesvCOo32myU5AA8OEY5A
tpPn5ID395/V0xTIzD5HMJX6mGcWheDSB4ib8smkP05EqFv3blun5OuBBhU/tWgQ
R4tJzykkqswuNHKQazAABbUDuw8hUi6zYaXiKCPQFyUAZG9pLnxJqZSU+YJb9KFe
hhFu/kXCBQAm3TRcPMcWL7O6xwL3BxO0t71QDHcWtz+EUckDWbWmnVS2Nno1V1Bs
MJJ0gM5fXSDmtqFNYpD5keDzsTFuwI8LvORlXUHaHoPbWrIXmFxp7VNBjYgsm8qQ
7DR49G2BoQEgw8PbpSOU9yEPC7CCUpeTcfPsvD9XXbYBqHaziJ555A4UzqLie88z
m0YFPAV0/gK2W8V8th4fQyKC/d/S4Ip/9FnMxCaeEMcQFeKVsviszg0EVaovYAYV
xjZXNugfOwODEPxIoy4AIP5232ylte5WKKRF72LaFFM+rPKLDPp6n9aBpEv0xFlB
f7PZKnNVxrh57ZI93C/hM+6fVWi+ixjnDkzwZ4dAbkA37isWRwKXzkgt9CYdtQ4r
BmZdr6p6xquIwfK4MlUunbqCZ3IyFmWmmIwI/AM4hA9485vmDiw8KQOmLJOvaFG7
MqOYTYbkXRd2VPzidJ2VxB8AweaIvr8aaBZODe9oP19HtZU+3V2moRFVh85XmkDm
F4Qv0Pz9UAmMQSm7kSAF11G5ijQ2BDzpHJslF3K7ZmghNK3e7YxNqzywlojabuwu
s+MRAFYmAVTYYa6CyuJvThVJIwWAZwIoA966lcLkrxONdBzVvgrKdOsW7lLcYjoT
iQpcxCGCTJ5om2Gy+7LH0AurDv2KVGkuTM7EpvC6dsd2z9O6y32NJ5EQpsInO6uf
a8NjChdE3h5O8gI0HkLk8TnXCtxehffTllTYAbo2LVS2AbyVpEwBfi3sO5FGJGp9
ON4KPvHr9jlOpJtnmUDS9qXhnqGvIAXgLFF2gt+/RdvEHIuk4my+1HYx9HwGYirY
OYmAIuExclqrfM9wxruo33rxG+87GR1r9INmreiwK1mu7j38B6booUEt4FwCaRXH
oZpX/MADyRk1JGcffU/OkNRCIjwReHewtBnT16+PgvqcQUnjQw4ZphdI8nPTBkK+
iSdJgwz4zHPz2drS6KU9QLmkieTU1LhbltAIrAgsJ6nw2J17KHxfwu6yEYkybULR
z/W3DeEeAY9ybgOmaG9gQu3Vc9CLyKNYkF1EUpVqNjlPEGX3w7oraqH0UWFdpzQl
PCkVwULrM7Yx+br5Ns9c+CMux5gAbkAfUquKFtrQ1heD4tyhglV3A8GnKPGqv/h9
AVyw1PBv3P7HZBVsogWhfGJZR4X8Tx9EauBKGLijyzr+3ZeBFRD0ufiwqYu9d3x8
go4zUnS+tsg11lTulcogPjOJav5spO6ldtFLBdeWAMrZlbrwl+u8pCtklrHyaYLy
zFcW03bP+Np7ERs7rjJgB+Ci1Z2eX2gR4GDqmN54Dfvf0XZ8kAzyBsLkPR5lQS4h
/Nj3DovTvqqOh8yTyqoNJ9RgH4AfOgNqJrY+kFrYBfjQGzW3iySl9rE2nAD4NkY/
4pulBR+HNxxQSF3ZUWxESoN0JUiLuvJ1w21YSqY2yTEHv1DHnCAnGy1Rde0le932
fCKPFNnmvrx9rAlzYq5pDqWmE0rBSySDsqNAFBTUY+MSeVYMbRVBRP18eZBl6OIU
VeFz0oCT1HJPmZZY1spIf01AQmRkYgm5kGzxMrFSsINAPZT34WfapWz1hEGURTT0
JAZKBeZoEIWxi0xesNL9QD6QF2wKR2nvFF0DIUx3Zg6BlkcZzyA9FUmzVtSUmhZm
wySXUa7mXVMms+RUDXU9ffEJ/hw0tp2bQ5fpJCKEYDwrZFz7Ox3q0LnUAzxFiO0s
X5KyPWxB7nK55UKRWu4iU3+QZqwXgDz4sE/O1Hz9ReI7cFh1xNIB50AZkvBBT4tW
DY5rtW559qLX5m9rjwe/8d92UyFX2mW8RK0rQAk/35wJlqq60bJNAt/UtSBWUt/h
uyG+aU7Z5/xFVs0rFFD8l0Lj2iOS6X+bYyhh4qq68OdHagc/fdO4TludHuB7AkEA
Bkd2toeGlpEBu3Vg1C2OAJOs/RUAc1r5ijb2JAqAxZDguGjATJjdz4W22cDJNsqu
gUisJBZKjrglvWRhLpVDMiAUom8gkiyL1IMtRqNZPuvWCb3G77/tsP+PsEsyWu1n
o8+gyTWugFsqx86cFDflp3CWIIz1Tb1O1L94PgeglOV5aVAz5f7RYpbJtHdIHT0E
F5tXNW4lcrOjQ+bWapl4ggmFqja5gLkC2DcA0qVWr9Ei+zCs3yQA790vzgeCE+eP
thTy2PvxkaoqBENe8q2ni2D09hdbYDB51vnAQe79bEB8aSsit0AyKqu/STW6kvx2
fjt+ZctoAvcLZKdiAqM0sPlVgBrrTG3AVgYAQZrho20Kh8pfcL5CRkpmYzlMw5/+
jumovp+CT49rxF7ClRnOYqT3aGYWgOaM088fzMGTHSr6IyDDlRdovQFBY3aCOENJ
etIHt6WrLp/KeIS9raBEudbCsN4S/oP+VF+oMrLG8nGUYU8VM2zII6nE07Gbx5AC
hZQG5RqsYa+wBR3TE3CwXmMZilcdEhtJOL/AZV1KzpnMppxXyz3evd3scb0ENVx/
b1I8ZfD3Vest+INi59dBI2Ppp7Whc7BJhT12GFHmCVZ31EEZ6XCZGF4Wx4mQP+sG
zwv2ZuboMplndAA2BD9hZXtrDJ7iGNpqXtfW7zGtxdfYMmktaB13FSJiASDcoF9N
lNI7mOGhquxfs9xWEYf0Xg33aWtKGuynpg/G0jXLk8usqiBWbfzCZTa3VVBOOY9e
a9TPzwFobY/7MXy6XkJ0y+XYyzgWBnO7JkCiirUong3sshbJLoN7Ec0yf76Ry7O3
q+z2cyzXbr7ZBT6tjlhi7aeruLOmWiDqQ1xQzfh4uXV470iXYbJ2Sl06krUnmYou
wj8bvbrCi4+Wnz3M4jpPi0jWZ7yVoItfHQzyBaEaLrR4vxFCJxgD7yitOJs3f6h6
nxXG8hy0A4i6k4I1dzDmjkMNH5H+b49s7Z6WoEt3Sbi/tdrZ2cwhoi6B8fylypGK
KXLkjJW3a3I6gYauefF8x0wrb1KAW8Af5ESYvO80sZ8pViPM4LZ7RE1wZshvWLgC
e7WJjqRQlSsJB/k1FPBco1QDCExcJKIrWEO1g8GmoF/JJ8vi+XQP7DrmC74AjQuL
PbvgcW6RXYHekB5GOAnorOxYmGygd/waycjWG/gsvAxtiJfhVYvbxOp8H5BoDHQz
+l6plnDJMCZ3TgxrVF7mZZdsIC2KbWZ0P44K+jHv2PVSDN7cZe/jiqR6zlr7Leq4
wrSVCFMkLmoFUsIIT8cxC0tzrGgdGvaa2k6PGTKM7oS++px7vCNZ+brThb/h8p2v
g/jT5QFoeO3C1NJcM4uUtt0ucfFFdM5AE1FoAEotU8LS0Ruke1qIysSRsDnwiqwb
NlfchRd70iYfA3RO+QXpI36n/UJeeoQQTcmLLczIFOZ+LtCr1/gz6Q1DmTxuGfGE
Xe54skH8iWzA8QVTVVxSKVMzhwp42fP3U9KDfcYeUu/WJhOrIxtDdh0eW6VJhMhT
n8hXuwCm+9lwIJX/3MCJeUKLxU/Rkau4IIzSg6GWpU20bMWrorNOk0AdSWllrYRD
hgWypejdUl0J+4+uxnUPi43KMfbQPIiDV36TS2aNwspJZ1UhKdINLlBJotuLilcz
k7xUUk1wDSIGsSgeC1BzXLuHKWpGq3/0ATVzS0kwgC+uWmTW8YxxHfyFD5lBHYRn
gaANg5xWJXaK+z3KrEr/Irf0pQ4tVakSZPmYaBpayQ/bUox2AY/sXTXNqWuCTuVe
rMEe5069cxOd3jrL0jiTh6n7/j8/MlssNxZJKLVCG5pdPlgkWzP6JdLOGqgZQ1Ed
HC4UczqjudkU/k7WU4Vr+WYwOyPCWayU03P05zGDPwnnwcpwZO29lcUrxgQ4Szez
DFR3c3TeEv6Hq7FqGa2HjBcjap+Zq1V8d/GDNyoaxEi9kop6MVoZ1ZHXZBET9ni7
waWRSvlj0tkqWCE1Lxw4h8d6wTJT/v6NOaV/pMKSql4uGUSbdgFIEV7zb+bVnWe2
F0DMKGbTaM9WxVcDiigJcst8bqk5RTAggsAUiYM1MzQrersq8AM9DqwXEJ+tYIFi
8tDkcRTnOhDrUUtmBlrWBkM4DiGYHrFr3hfrv5IfiOivgZWkBzQEiBlMQNNSTD7D
Mv0PY25nQZA+k4PEYVjZi7MDwe3aSfGLn3IsdwD2BKiPUZb+KnGQXSXXR67tJYAd
O9guyqqZddyCC10HjO/bnKh4cjohY4SFfCae2yucZzlDdRwsRnZZIY16dV02JVE/
kiS76joB9xnoKmIYit1ZXhyWGW1sv/D/UEYcO0vr9fCyi6dRqOfrpgYKmTfjGmAE
EPyfZ2luaaqTy/s0RpAqVnle+YpoZWcy2Ih6ZVLMz5qwtx/fKwrZjNzp5Z3HuYQU
h00C5S0k1xZFpwhT1Akio78V/qxOz2/taKbzF6HfUgVkDzzQhlkpuK4h1/VgUvtJ
zSBmr+pPtHj7hQr1oal8RZe4huTR3B0iBlcohrURv0njNOqJKAVBRt2vmSudBPLd
SWkUkgJDcyeoOFOPmg/V1g1BfU6K6ef/Yi7NJ3vfuJEB3gZbZXpyN3w4sFvaKhWM
RyUBWGTQzjEdPdN7pbDzbrQc1Z+qePIOGONAv2ewS9goWjzDnu87VR6JAX01QIdT
I1wxmejHVVOsM34N3+HSYsBQ6osFqSxbcfLMa/Hcobag6/2kBCxsb9qlcL7+0Lti
lYeWB03nwhWYWll/q8JeDAMhSMPvK4P4tuYRDEeQzGJbdq05DFceVQ79kYrldV8L
l/tfi2zY1DWlWVPfRkpr9sugR+JdiqZoEWzix4OL403rbj9QXNP5ZngEu8S+c12d
yYdkPf1B1xuhtITxgB0j3KjHvcqSJ7oDSm3NjUQ0YSkrZaacn2TQ7KEkBiSQvMbW
GIIJZDnCNR207Nt2/nU85sUdbTSn52SaVROy0N7Wb+2hMzfQwMpdQDZkrcuPdUlO
pg98+qRmDcOzQ0DSoA1Fkf+mh/YbO6EhF4z1dxpj5oamgTjRfuvGIN6y4l9RKVXu
Mnjo9O2/Ph8FKIyarP0Nk2VE6CP69D/bVPX8FGPF7BfWRRZW3L9wI+IN+7vtVAi5
icjHg6JYUQqfJSx/Dq16LoQq0RCUVXZP5NydBi7V3GtF0mwOR2pIoCwbnL8QYLoM
muLPpkeFvYwAGsdiT8FjPPxsu5G2bIHqp35uW0x09VXADEeUq0tQrB2X3Aw6ZwY1
x1qJNmeTKUohKNOXpEcPOah9wwLWobzJMzHtXIQdoYUEqdTS+S61qvXsnFlq73UC
yljQ+nXs3CCB1icoASMaRNB8l51EetDbAVMmIy127EidwVjlMq0cIOgVXDTscTHM
qON2WTLHpr9DIDqttZQpiX4d0ZdF9/tbmlrG/D5rBsyFMwDuyX2GvIMaSrOP07A5
hIkKAg5owjGiJWqk+rqgBuM3zWNZwf7EzKd9UzfQxvC5+0Im4IYQjU3wSPpQfr5I
AYwMyVA0EkbMMKJ0k5d3NmYtTUXay/aEV8XqLjvQS2fxo4RsMK85MnRBxy3FQwY2
9aIm8zTxGO0HkVclJTML2qToEKxKeHA/MKKIE83AVC7zALRmCZi5SIPTTpoMzlhb
0/9DygK7zVMG8NIqeDjCU23AphWNLrmACPIkdIYtKoaHNaq/S1IGiFeAsvlDzTYM
OzrcYbArCLU8dVuMNgRMXcKuao/Usc6xrcjNN3eNlCR1Nqr5EQEgp4XTD4Hv8W9d
Ne9IUKASXFznGq5HMp/cU7Eh4EHkV7k3Vn9rqCYHDZNbKavYlFYADHZJFJDD9t/X
zOC8QBmn8h1kSdPPhzvIK7ISJO4UN29TvIiu3gyls6c74b4AAcZ+UB0JXzl/x2FE
3Cb6Drcbn1f9zf1TmTcpeARkmnO1qRfWlJxyYChn0358Rr8Y8c6geDJ8NXxMuQgD
HFqrepKA9fjAVJYi81ZA5IsaNj14Yzgkh+g3qpPPXrWhMB4pMwGxC3Qlh/99cnvw
yRzFnmbyyM+WZz1JkEnA/Ts7FanHbBN10wgYj3ru1tu68L6QC4XLyZ5IO6La4xGj
nSV+tpotIUcpycB7aAXZh3kOH1bmH+3qU8ryoGXCodLWGZ0t3T6SjMJXNvlHUKRj
nEqnt6KQVIbkHn7YFjoGIzkl6gld91PEssO7q1RAbM0lbDy1EB1izPPo/rVXflZC
o+Qwt8yUuhl0HFfhHJUPW02yCOfYacGE8W2JT234fIbxOrb2ggMOo0gfNfcUZm3G
Zv1NZaoxjyfLz77gl2Z5jxB6heKZ6TDN+QYqbdYTlBfPJXlEHm5Lpbe1tewYV5rN
qZY1gC5lcQQ/qVSc1Ps68B+p62XaCj0N9jfg/1FcpUClQTawA5VLuC1ZaWdphKiQ
n1bODgjoXdCtdDBWGnCUHtJPjiJoC3Cso7qbnvx1D+iOi0CABU73HgVbwUJMR2D1
2R0Is1f+zCPiRGsLjTBNxwj3zlO6Jm6EEvcA++6DyCA+HcIwhpSCcwLLj/tZdgSj
1w+vGAiFjlJTwQ4n0bpE5vVG+SeGZl+ZVVvgyNJ3B1TPynYh6IDjpXFMEhojMv72
oyYa8lf/ZUeMW3FQW1Bt7osRCH4yPch+qeJVAgLebt28+SZbjizHXLcgQCe+xfAM
SN/5imh7P5bSkDAJzHH/k95d50bpItfaHZgK19nAClo8erjZ76j7MW8ssn7+V4cl
czXEtxD95rMHC0DxvQOQtfq4HnNsm3tw0E2YE24CbxTni4XFCl92DKssp8BRt/jE
8xZYJrvgDmNefJk/3WrGyj1QU6pAIvPvDXSDCMwZoV/Gk3GtN2luyCaM4mf9HDBh
lWNWQY4qKepDk1J7KSKYWYM0jaxeQ1z8LIkLqo6er3yy+l6Je6Z9YooaYXalz2Uv
4OwLDiVLS/Y3Y5xO8L9Nfb3yHg13MLwplzfG340voXmnKxzDwMq1D/W+oN8YVg2t
C6g//ZMhSn0R5t/3NVxu9j5lKbAgMhdvbpv174MhKx7tuTr1YJwwZw4bry5t956Q
30jolzy6OacGVBBPk67Twx2mF9bMY/fS71JIXNFTOTD+iLEhm0d1+T/UWC35kA5n
GjMt4EzGUyieOARfoyx9QwdlZVnYWHBzIAfVl5Tsu6CX/1RSJ7lAjhD/IYcc5nG2
CKszgWOhW8kSdq+JNSXeHjI3V+Ya7TN6XSgWjrr/eck7pP6mNUsrDpCPWhHUm9yF
E3kv6BBVczk2lDiIPazamy1DdnuJsWjSS8NBJZFm37bzLRhK086x0RqmHCSs9HGd
SxU4zduE/TZiOL2ZGaWhEJntFjA+E1EXb+JTUfpEw/dgi9DgZmgxRSOlSWVQg8zM
7A4mCegwR7lHoI6Af6IyHDccwFWeA+an3hzEJlXvUuWNSRRC/3cuo5U3UawithL2
OP4gEV2DT4OkZj2SlxdaHv28sP5FrSpwnhO0jLji+7ebaJ8fU7eQK0XwYRDsJ+Nd
ujk11AeGmZt5+izDHuenJuQjixsV1N/jGLsbj86cGjWErdu6Dedf3eX2ZpCiCQNS
EiM60R7cuMLP7vxoBMxGaE5LT3GnLIzYhJnuFs5xN0M13GRGg7MRC7mveanMuixn
pD3EWPjtC5jGlomKe1OnqtRJSoPBD3ZoHvHI8fR6jB9GgGxNkr77/OSVFNLQpWO0
BBOSeWgX1JN5PJBIlL2t2hFBYL+Mw6KgJEgPhaDWi8X0S24CqYgrpQOOsqD/hP2N
/B7Zzo074JfX6rca+ELvhoC6v6MjBUaNVGjh+hlz7jO6Ij5VbBqUGBR9Xw+/Y4Ml
IOnToopnRZ0pSpit7Lkj3fWRPLi8DLnPusZsCQBW6+1210DSxm1BW+UQzxPc/VuE
r15IuyqQnq6Ajhenpae6uBg5JnMsSJabwOGx71EF6hsrldqcKpfL9gpjVNqh1Jkf
kM+KfMyZc5FOXtXLQOhVapYO1DS59qWIQZALHKQPm/QCw2opMogCw1gZYXaG2qtZ
tpq5Qpibkplgv7h7hhsK1QyvK02b0QQLFAAcWm96N0x7PYPWbJDg05O2eW6X/ALH
Jf9eqLFc+mCBwzTjPGDJOrt57bWC4WGd8L5VNe1GiKqeg3tZxclWLW6Z5EsRnbmV
33DadZ6r7aZr/tXB2aH6Z+MC78NjfrSPIgkSowNIwGoR77vmY72+LFoOc3uiYf81
ZIsbzWsB39tXXnC5N70/qTNXGlSmIn4wc258Y0MAbkbdjt0XGfC2HW3lsA8E9Xe3
vjFPkRAt7Tby9WFfsRU58s53cSWHpMVz88hIEOB5IOdLXoxRZDrj2dfXz/BnwF7k
Zqe4Og01TvvQ/3wQLedTwg0Pck6PVuPn4NM3thSMD+gUh21zkaxC1U8CZYKqa4O0
i5wxAI8sFlm6plK0r5AQQf0ixpuJX2WsBVKjZjrr5NJ3eeLTshgv+Ngo6CD55+SC
T31+tym/SorsWBTwlOSkF2La3qgGZhadbD7Q6I7oPXzwE8MTUpXyAqVxpRytKTR8
G/9tOrHeaTSGVdaS1ItT730vGeFpgmkk6jy8LvJ/5isLqJUcdhrpPKzJGerp3656
hb4BAdbJZbAxDA6UlshU6V3weg9HjxjBj3qYJJKxMZ0hh4X1kvx2k1C4iHiwWrIs
tGLvLqrzCjqQMEL6Q9g+2UfUkh1H5hvdAznewB6PdrsStpdWHb+Kf7ZQwFdc/utf
vDlxD9aHvnTaBz2OWkZTP5NtSZssL5+xsrQI0NDh+X8MRsQL6OKd48thb6/B+Vyp
U6OHgieOzB6lxB9SZ6UDl6vT4JZdBhuPPu41l4eKsgeeSjFdy5MKaiK7yu/p6r+U
SjbVQYkz+vAuAD7BzHh7oyBUWbvXZRYTcS/fvGVwdoMooNUDnbsPmERmomTLYNYH
c+4LXaJSyNSR0VqnGx/C39ToPdS08aCP0nsOfMO07YCYkhy+H9D9ZqHrzyPCrctZ
1ONlZWe3/LCYayQFnslUnFxYNGByDN7dxaeMrOdKf5LN36BVNrzPRiliJczhS7JC
LkjlhIiEvimDviD/WWXB6UBdlRdZJHX/oCWnvXVj8Ktl2Ce8MH5oSNDN0qgDcXaP
6KV1M0ALPHU/H0uakL20HM3qaBCZX9PpwMNZvneI313988O0fUmp7wn5J94FuHEm
5ouAclbIEuNjRhLUmeOHxe0IYGT7X22VUsAqJutwgky6qbB2cjno2WzQHtbyNTqn
HVhj6iyJp045XU59Eva7hA1z7mIG5HM+yiP7OfkQapUXk7FYxxrDU7sZAXQA7tXL
xZujqEOtuqkeLxmRP7I1Bpx8OOubPu69dZMLJfs6WqKiC7staZfRzifqc2vz7Pbq
VG5eouefDM/ZQlOK3R2hzmdR1u+ua6UuI7EiVUc1vngXrPSe4uWaYtpT/GsfSDgX
2v/hyBrRZ825P3TyYPdrJlwMR48LbMQbu4ADYAy6+wAb/vo4u1zojrtu6HFxhbfe
qm6uJGzcn644LVBXQQI0kNKDpMk2VCR+1cNcHnmNNJMMEEQUcAv9J7uLbbP3hWJ6
omsnLrm7JkuwWA7IHTtrSZyC8MLVYU0mYh6mR629ugKBXxH87872VJlNQd4xifF8
m2J1ASyoBwhE2HsvSeOtgM486H+TLL23CfY8cR1VSmZidGPtxATpiV3iQ98Nxn7H
24DDHPcP2kLhXIM+UM6ehW8+MEcWCPVru1eAWqUoIgzKNv6nucrZx7LRgQqOAL7O
ZlXwjjbMQgqqh8suvnn+Sc4Xc9LPLL6BUtyhxhJxQ2+Bu20VD/IDWYdt+1QVwrgu
7qt0wSsVKcjfKsJ39DL9h3HOxUrOj5WVOVFYBiLiYLzpzGSddIjYw/CobO157dXx
zu5R19FV06ItFKUYwsb31jwiOz8ZY3Wn4jfShopogaei8Ri2QqoKIBRpyhxfHueE
pd544ToQEH7joa2T1r3W8geLVgzqIV/PfHbvEtI1NRo/isIW4yvBmgDeyEn38uUd
nJSvVbmYCBKxbFBy+v195HtfGEPXVq/L+n56Znblypl69F+N22oFJmOvO8DDJUgc
lvz0EaqC1yCMxAkY0OUZa/KXpU/gLWtMw3qCaPlR0WAdDofkW58mxAmbqt03qHbB
FovJRmx/yWKTf5oQPlEUxeEV1Xtxh6M0VB2Z49VO7IYs8N4moLPFK0YJPNRuECm7
ucUMbEo4lxmi6WSstCNSb4LMIbMvBHNqi1nGxPnpLro+tYcH4f/knW/Ud97GIXMN
rGNgSV4GejeyJUCTouhcLdKPDY3Fuemg4pEVrSqAuFHXBNS1bb/TtAdby11E9LV1
RKg0iWL3QqS2I72moNpcv2YVczXFgbhY0FjPOA6A/rTKrUyPoW5q5DlSKokSFBGd
j0hKGk1DyV2nlv1JYTuUG9IMErT1dkCpUc5gXTPezzuJpk+nFb7d4+c7PbePBVXK
vfIXzCpR/4IhPo5CMZyIJl5qcp5W51BFROpYGfNA9QzjNMGsGmAOR3oRDzI43CC7
EDrYsy76GX13V2zGt+FDqIovku1g6cBvLzRw6QZdGoFsZjLvqwB46xuLxWL5lHns
YrGPgIzH5e3v+avmHcKGNa707OWDWHXeNcncLgQlsDBB5p6X+di0Guzq46TG8i2q
sCa1Y46GeU1dxkw7N+lNRpjioczQnad+HhGTHqeWv8fM7SGdEpmFDmnsNICXUcuO
qS6MWkFGCEzPQgJinT8THiQQHpBwrb8Z8BPhg8j/G/NRrr9m9MLPIylCtENltJ0H
fNN/AnExdYWKmqOIEl4mD37/2jpL3l7UIxtcAUdyJNTWY+jvZsy6HaBiZhiVWxjl
swscoEH4DG584jVh2+DW/ytGpCDLc3xuTLDV08PM+FQ4HcLiePx3cyFSSHmLWp10
W+ZLy2k6zPUWh64Hk/qKeF4EMc8wc9QAbK/Ts6WEZVLv6dsOZNEexd1Ax+OebUX0
UgyWtbeYQtdTglJCY+SR7NklhlDiLm+T+9MfJPtUkQNeCLW/V7K9A884+YwzLGDc
x9YmepXvaoN2Tcg9nNVotWNnSx3F53//Wl72w774KyHVdOQKHjvF1eh++fa5l9hX
kr+Bq2yndqDTlasclEiQCaDE1PjmGt7D81vCmRP297tFt9XW75/JSUdhFiaB2Ctr
ijTtrDtyEGRse33dZ1L8t/kA1ojgjP7w7rdIKwL17m900L4UUnlqGljG+1b4rIvd
JCY9phhqI8hC+p9FA9AL8tilY9aqJWUoEIEgc7+QD8oW5UdzcmU7EROiPK+F0amV
G8UAYs/Fyx9bKkysFw5XwxYzlfoCf/dxn2aKKL4myJeu+1rKzG6r4nKB+mn5TOss
ku8SqpuLyELgPTtpiXGu2t7Ctecj6OL6maIh0Azs9xjaN0cjOmP+t1l0mlgPTZMO
IeMozSuChkdnoG3IKt245cHRe/KCeAHVZTTSfsDpVvZryuPFhJHocmwX5Zoi5Eak
YK3z6tyE4Ka4Uw+BDO9aMKd1mNljwzO0NGa5XC3ZsTtCqtaFolVHEJnlMVkbbMpd
wKl5laBkkZE+HrtTxpX8/+pS2iW1NKXTOtR0oylX3+2pPZgvVmagMSiCO9b4xxHa
zsmD9q8T3Ts1o0sWV8nTndyg06KUAExP/rCkgYQQpwVrCafNAlcslnLSmBN1/LyW
7dHfpGKoBECProaxZkivKGRlwCppmJYUua8QhZdT+ReVAITY/yWEOusjwvTc4BqX
sgI4UyIqEbXQXfPHXTTGhpjnS3RvjZa9wwwpzCdBdgen69I+SOtEz4cqI5WuPfJx
TVo/uvCCIxJ+GMh2IY8tufCD5XEUBN4qtC8cN7udJzvoK+hcB3VjxsTGQK/ouUjj
BGtRYQvspVNU0U/27ovPA9eDT9EinJh52t9KcOMwnOws2C6nzZVVUKvGuZb+PoE1
wRr9R5c+2XRypyEDDslac8TnHMKJOMe0T4KDyMHOhENtbGxnfdV5V4E60z1sgLid
mt9KlZqZYCnBbgZL+x7eMG52CRK+NCglUo+ESKnrOKKgy0pqzbM9Uc7RqszKa5ta
Cs5xGihKP6m9yIPMlWxnaLnLbxuN0jRC7fH5O8WLtvfJg/shlao48HenOPA/ECcY
vaZ86qs11qvw2sy3qZf1YRKPWpOnFYOEjGkVE2Dripgu3wiAGbuHEvE+gTeG2J6E
65ANTtOw3UR/vRAsHm7JY5R4R1zzuj1g8BbKvFCxJuNJIaA34Vy4PyfT6pv3h1ln
o1Virjl2uCNrh7Z1hVRVJryhBEFpyVWbd9qJHdmG5Kjzl275n5rcuLXAAu9DWJ8l
3c83t20SsMgWImVhT8n+Xp3qcMcO2gDX3zynrp+hu1B87tPkHCSZnmulOIb58zG8
FSl/by91BgDuk2eUifedirxYjAbhXv3E+bKqGxGpu2ocAKJ6VFqRHlQYF412fD0b
6Ijhhx+FT9KiX1I57kdNT9q4FbdK/LmpSQwbQ/zh7CKjacdI2Mi3uJwf8xiV8544
Cw+66mCGvssOcAktElgiGpPjVt4OYcU3shvwgin1Zu/UTTUW7H4orKgLc0LT1dTW
yzXphn02ijBRGzray9owbWRvA4a/Z32fxvU/fbn0Vn1Jyi//Hu8kwpC4N1U4IKYu
oUmrKqlTfxIffum0sf3S4zYy9zeFH0/A1RyqWLiERxn4Lmre8Yyf44UBReP2L6DZ
+2kTJsdj5QBdmDWEpGAYfqnXGWhoNQJ8FUBnjF3yJI+Sn6+NMXOclHkiAtELBIQ6
PkNDDUARba+MNN8jxr6eA5MoHqxtJf4LyO0GoG6lQBbhkwL72CQdx1ME+lqPmrDm
jzmfq6BKT+lGWkwqWJ7myGvmhjCiTRXCHeXTX8XCKXdh9Yf5zfQORjijjcL2sp+n
xMCh3Oxwn136SiRSMQgv1pz1u7iUVHEC8lBG0j2r5uZT6ZQCYI9rU4IS7yrnVH/B
D9y6jLBws/5ft9Am288E36Ftpdu7afTP60e4iYj3zztqQxElftugTPXrP3mJhwCl
OlnAETpP8PeRYzFvYXXruyL5iO5zbaWpAomQ66OEm6wofUBcdN0tiBtJqvMHmn4R
ZOZO7voAR3VdnjhzLhzugRNQIA+qVAdqRPEk7JAx3d1IEP7EdBGgarnb8F5LWy4x
uEd6AXndN9sfTK7YrSNjhoQhrQYikoZ4BUu3bggv/nWMlUFbQ32n/kFAzFKvdJ2B
zplUSwMT6c/roIVYv66arExn6IH7ODlAroyNnN2zyCHpaevwp/znXWcP7eKFCgCn
8CmhHYaAuiHrDGJzhGr6tgxCCCdTtgH3mSpZAdgxwWLTo4EPHBPhX94V+61IWaaA
+O6yO0LWxqzrkfc3IqSA/jFpyeDTg3FM/b8raFOJ+NtAGPlGd1LX7u9f6xgOaqiB
OPDwshFaONwpO8ZJ+GYprHYfzM5TGACsWcZ5fG+VftDAu6hZoGyfyb/VroR8W/7w
COxcfnf8Iku6qCU67BaQiDyzmhezjhCwU6eCUaWfHB801ygVoQYvTiFIc/yZBZ/4
reUFX7I8loUqsisMc9Qp9cBiJDF6dL2U54ZUAKHvsmN92mWbM3chISU3eX01ZNM5
pFtuXwjj2HpT33oMESH/Z4Creb1e45ZFaX1F54uMfKw/2BL4J4DrjX9wtHDUOJjZ
gmLO9xhNh2lciAf8c+F3a6DaVC1MudcqQS/cDneu4c+zWmlMtDLqZODcC1jsTVpQ
5ITl/5azQwS2ZTFtfsvWmVRAPacd5wTaKcn7WYWW3x6h0ME0hxsKOc5TFMNtpKP3
UI/QX+kxnuYfCXuWI2y/3e+QKiNEnVagevKw9/b1Ob6m5DFsQAn1MbpHPl17AKf9
k/squzofa4BSc26VXxnx7me9cnn/Ej76+9SZs73d3buNp+Ia/1b+BE6RMWmEnh9c
cVDmxFMmuTgyJHFp5HVOvJ4ZB+rCqdY7uWxOH2QG8cJoAO8EyiN/lPBd6NRzQOjS
go368BkCHGJHaJMN2rdOhPw6H95Am0bEr0ugqipDOj+zvIlUkBqNpdd9dkIbi5a4
FeB07gubfQpubZlfmIfViCPmv6OmQiTsUKCe6/GoVVx7rqmWQVaeJi2A9SUlpPCy
4EypG3EdbCz89t++XcxWQKLAHvgKKtZNH53Yzrs2sIz9R9h20kO5HZ3taAlgltC6
JRj34YhIa8quL1D1sYugMGLIzmKmQtD8x/WlcoiQzlsE4c2hl2qBkmro6pf8d0Nr
MLbKZg3TZMeVal8vkFcSIl+8fdmDWTF3CkIbe3legQsoZc6RfccqTUxlxmAuK51g
rKNPjbTuWZBj8IJsQd9q1VYmuh6z9wWcI+znSQ/vJ5RDba+KaWSG54Pmq2qQ/a65
O5okHZdGKgNfTAfWo9Fn6Y6t37DMiVWxixaXicI4UazCV/vWX+nj6B6hZk0g//bu
60EJbL13mAWXKBfrAoymsDw4iXpgBOqc7jaOAHNjtq0rnTMtohO1dwBev5ZK97ZH
5L46tIFqI0lYyM1guSE/eRnhmer1XY23JdPI91qyevzckvtrhKuowBPs++dHeCmJ
p0Rq64Ov6wuWvQWTAcNIMJeRFY90RJtTio1jqDeVy2E9Y5io3VbbjOGp5Y9XX6Vb
PRg2J9U53hYJNmePsJS5ImmgKn7AjUkxiY8+lLYQqXfVJ/SpCdweFK0S+3Cb+ySc
JLqW0QPKKuRpQAaT4ZbTfUxKDR6QTTZAzsI6tjYimHSJjmioD2+3AnTRSHzYZKED
Nh9F4HF2V9sU1FMDdH6rOtfGlP51KLjCTmKSiEbw/Cva9pSrhADORqOeqrs8JhTd
Vy+9XrVWx3PlpRCXoXpE6HgAu8C4t0ORLz8Swio/ZX4rMFFTTTehjUNeCocohvl4
COcSsXo9XsZgdTRH8XLraeXORpZX2XGklzmoEYlADBDxdHjn7Gpg0t5fMm6UcynL
ozY7GNrsfSuRH5MuxW1dYb1NL0b0lcRtoQ98cK6eG0eaHD4HYfa1byLBBnD59Wws
g3Dpk03GM6wYw9uWn/0w2ivD7zBfPBsy+EIQB1MF826xAodle9HNEoAQ81xxDelt
1lOZCXxYzdX1/+zIetbg/61+M9OIWrhuwXdm6To19spg1r5H8U8+oO5woyMaPRKL
CeOOZyhAX+tXpBDSqS2mqvxiz8xc176WwKZvQMAygefDAy+LAkyyIwvsS2ZdEjsC
S2Hv2TuKsLPw45c3M9FBtYaQ9jqyJrF5Rzt6F+3s5NKXLd52GKRGdrs1OdfUJtWy
DUwwJoSw+rd/ECwnXY4zTXvo2JD+WKNENf7O9hHBKP86hfpyQiPNnOMj0TfXWjAV
pA4xrWw2+Lqz0eRzblg0btEtwsKRI2OTwDtZLzoXolKhdkzUYZWxxqXUB01hjH8j
euE4q5mwAep1Yja5oYdxcyffMqF8ldQHsozRVqvy48GdplbwvIIlxQ/teIImLa0Q
6ZpSnXjXMb8l8TVyplvpS2zNVu8ZqS0RIBer6V2tV7uSbuiQY+H3BDlaN4AjuPy8
pb42h90NVm+aQ1ZKPTFxw4hVy90epYOdGspOaRld5osc9I+KBZC+Swwf/7pUik8W
oK9oIaAi+GiMX8f+GzTh/amcSKjgLaUeRL21HTsr0efVM/dLNlyscd2X3oYy508I
uu9GW+o6yU+ipMX85XpNMgSKXmlFiHSkv6ip66PHXHRUur+yXNsNqK091r8LsEy1
xXFefTzbW5/NXCudW/9LE8jG26JoEQ3eEndeckbsm8l3uQidAzUMdBRqAnJ7iYPH
9h4qjJzsVOnMIH/QTXOkgL6oMw9W34UXZxmZEwFOgPaNOEGi66ThIEb6mNHV1qRy
URpE75hvPmqVA+vKKOue6wX1YIQxcLTfpOWikVBddTcCyF3PeSo751XIHU1V+c69
qjicEA8jwQvfEQTZpixk61GonlBJad4x0iH2JE6zX0zr52Kcfwzk4wOIVdfGhDTp
EHE4pEE14g48iMS0Tkm9qI9bMWJ0eQuXqAYRhuK1S8IyXjbGZgfAOU490WSPsRV4
uRMQoWbV21wWbuJk/3SczsqrzF4F/F/5Kb6HrcKUNfYjGUL3a6jdM0ud74KSEaHv
3S5KeXPCgZoDpUoPNaMDc2mJYSVvLzg7MLAucJWB3CkogGykFQFP1mZ0L/YCGfCx
yF/NQnfzKrjKQclvY2aYL7b7un4JEI3nB8G3WsaFkiPpspR93UKgTNDRS61eKRjX
T9pWvVCAYMrPkVw4BdRuKDrWPu8XhR5HDtoAyC3esIeu/g+r7qTP34phps6CgpuB
ZmmGKYaS6ckdjbuoTaBLEK4wPWYfhWwUva1lGEx8mFHcHMSpiseyEwHkXaRXxVOC
GIU2/0P8z0IMCkfbTXOKWWWuQok1B0qZ5Di6ayl2fDDqBh2bkg8sguHnlVniEpsT
CE6cwlNMaJ1n71aZXNWekdk2APJ7N14b1snifS8p06BUJdoYA7R3vNXQzHACJtbd
9YvRAc3kpUVMFuhoM9Wu7YVZ/QBpq7Gh7LzznScaQYAaxHRjMbarAEUMkEjoNK7o
MZqIXTXBfvMrf9JsPz/hSgBgD/sQUoJIUiMD+rafGbt7/eGRc+fQIukzQ8L6PnZo
F5dDuhJcJW2bf6C4bRBqrhua57uYKBHjfazS+K//sQQVZgfJjdMMkkgIlBNGwWZL
UwCY9ynP6EoxYTgHqDqmZL78bpmjyI+Tpi+bxcZ24lMsNhv/CNQFcfe7Wmj2Q5Yd
Yp1K84EVQr0xDSSkRxX5iRvKWsB7CBzSd0OtaoPTwrzuoD+vMrZEDykz6rybdbXD
J/UH4JnIM5zNf05r1PYyZluVaGXOUwSKhMy48wKRWt8vXKIaPaNnW4VfxC3M+gK4
y3xBjQnj/kuOkqF9EeX9kZ8Cds7nz/Y/SruUR1PkK20eH1wxepi9ds/bPoUzo672
VwaZEtkiFIVVDOdMYwq4lqms6VHBd4/DhKqmyjW5f+EtDQ/zHweVgZTCFRZsITfu
xx3Dfz1GmGIU/PWH0EGl1o5CGA4/B2hbBSySACo4v6ysTwOpzVsi2FhCcpxYKeAd
+7PMIkQYXL86onY5zm55gWjm1CMn8DDtFOwsmIrpq1CTzwjSz1KfUrNQrHk3K4JZ
mXtBawPhYEWS3f619fEIl9ZErRv6vPcrp9KxtZPQvlR2QxG9imFSedrh957TYana
f1KMCoKVVf8fRhz2ITD9NESJhSGCoLrm8BbUdg0eHUF7y4sId+vUReulZ00rBW+M
RDtEBbx0QMFxNg0KID/dtY1G3ws2BeUk6imFjzOyPegLaAe9dhKKMOSAC7mkrm4h
7hOEl75u22s1AGSgBOuJ3THzR6XoAE4IjLy65JNxAy4orKspdUnZVOy7YJGc5ktD
LA7TEb/NwH7WJYuftvXggE3qY3zQXR9coTO5OTh0YUOdqT9MwI9Xjh3NX86OK/n1
XIn7hW7me+mDehrjN/JnnkxP0SYf1Y/Bgi29mzfAZ5T335aT9VNnXzm1qwWSHIhu
O6stGRraU0mIsuWGhR/I6uGKcW6LJ7VsQFjhl1UpOEi1yoZ6Y5MeGFI7nzahfVrq
sRz2WlsjH0+CvKQg+7/xkzEWwf+Onm/XPnbJdNPb8tLwj+10OcHi/saPf+WibAtC
GC8iXtv1B/PdB0TEebZ2spuxvgJjJJtlQgjhk+PvA3nz8QtDUCBmXRGxeeCkvn+v
MQM8KEL4DPfj0F8Jqu2uKA+3e2Do/SGL5naB8xw+eopez1Izi70jB3SCKAyBcf34
GakgWdlUhBdrugoBhk4GkglXt+J9nSiiogIPg6fOeHIWdURXzS7x2gO2yCWLGTgt
deNgjnNdNBN6klGpkng25ZaSBR1mJkIjkSzu34UMkBg9ueZzhl4+jfKuNkP/AJJZ
LVU8OEX0S+jLJXd4v0B8b0efeuZYjCBRO43fG1oPfURwwUOpog2jJ9y6q2S0U2i/
KE+b6N/CbqZ+lXmIOcnt5ctls27ihc5sbm5f7akrmluIVeUPwUlwWrIDYZ3ZfMKH
LSWSoPc18gTK8wfY9SVNT9IJYCt73fvL77bwHpkiUkee0O7Dc7RZGEFK5oP77P0u
HpDmrF9NRyxOQ0Zx7s552fq2I3AoUkEyOJnfPvYySJxTQ56mSfoZvRwveFj4K99R
XPQ4XkbJtNXVsziaVG77ujt16EXBbRTWcRewzC1037QHk/QUeXi5W0Se5S+jKj3j
nYXhYInxxKRvz8NChfpd6oNzYxLEjn58injC0m8338Fd9Wk6X7vDs5pLLPqdPGrq
bmj7Fd5dE8ggo8loNmQE9qIWucR25ekiGhLHPuJoF8ei167xG/8mLNRftJNbkG8F
Gmy3gW83Hc2C+SFFUFUQdf5hz0JdqKlZ7PH4/oagbGc4zboVMjKh6rDK+HrCYVjg
TyGfgGGyW/H7ucIkKZ80Y9VGDm4R+dMvmRlM6UKWXecLPuVvMinMqvJVnjdP8bLg
Am5yr53iPQGmDpsjNKFdW9wCwZG+bFtS2ElMF9CQyq1W8CPokp+qQZsmBCFiH+NN
FVMgaMXk7lhpATx93xrNvK+O0ZExB/23PY2qOa56OP11g/iWcNphPOpH4UPYWJtE
M2MKHW3AG9K8P+rROfV2QiiRvxndWpAlrYGyeRYHO4WjU/gmW+JDUGzwpzPEH/+Q
MqREtN7kPpjO3WxA2f8a8ID5PDLNBlSx2sftnW933JHfJV620spo3T5bhZkLHRB7
4c4ruv7nNMewYUFWAKbKARLIUtzHXOtRwqR9h4/QPZm2TZ7nhC5CbtLjJN8I7+ij
iMjHgY2wyHuRwd2Afu/qTXEASom+vCbQt8JIx05dBkbJVNrSw0jbzOXtfuCePuBv
pVwpK8yVI8r820P3PgNiusozE+FwfRXNB/rDWxZzRrvQmQ5fMIjlfwKCDJBgPgUu
Obe6Hs69HWCp2fRS6Hws+LZMGugtj/nVPw1zYyo2OJDhDOzviZ0YSwyutH8X8fRE
tarZ3L0yui7b5Z26a0w+5uZQJABGZB7yH46pk/+hfhe6167gt5RJ78uIz7cZdayV
uQknJ7YwGaWaebnSPkXxJVfF2HzyfTMho4Yf2noIAWaXrlQuzXGD1288V49J9rZW
/5MtUKuUHrCsgwnrP+Upo4Zd1jcG9xSLurFtZtkbtzlkj47KwVUbxRdwaN3hooXh
ZKYnW3I5qKNF/TuLxu+thZt163DrbwTUnHS1pi/6qNlj75NwNfh9fnOPwyR6y7SQ
sSatuvWh5nd/YQst12kn6bXyd97w5L3AHELCQ+ycbvu24t2ezc0wlORsqW2ktSaH
5z5a5BPz69t2DX5EhZ9o24SU0Wce9lA71CByQSLSt7XQIA9/IPD493DkOzXm+bR7
LGT1Y1Cb140jG3pS0IKxG2mh6mNwn0gcINiV9XQl1W9pg55Q8wQ1VHcDyi82IbOf
DVvXBzhv/vsfiz/DPWRamoV1KngvpcjO8NUr89TxwvuCEcfYrgDk3dbLsD+i4RoW
riMo64FYAg9DGiigtx8xJ+0My8mOzxx6koqHaSLJlnQLICXB2kMCkyYE753muZ9x
jaJq79d/JY7jJ07w7LiM+azqIACoCOC9WHSQqJZ95EGihgtvZYwRA6X7mqH8W6kB
NpyM5U8PHrd98NZzo7A/6Dc5YrOKmrHvvwcH3WtXMc/8yc5svTV2E4gOsiPJ5pTP
wwUx60v7KnhxxmVqycDpRz5h1l6K4K+N+o8SMuqfdL9Iectio3hT3Du5tZeUhTnA
oO5iFw15SB1pfUI+Gw4PkSTYvU2Wm3xvIwLH1SaynHQsMtfGchAyWujCK914Tnc8
/61Ljc+dvJlZk6rXyFxuk1s/EV/3Oh/nYVPBC1S6QPjLvRuft5yGWUeLrZIzExsM
3QG3Gyei4o9rH/UQmkX0eG9nLE86mbnKdNuxACtUVu+jOXFmsYqnfO6rMnZgScji
B3Crf6Y9CdImVPEAJ9N6tMk9bab6zBcEDTkgJbq62k9+FBNaMfgDwk/NLFESL5qM
fgrXRGybW6U137apiAA3o77ZOZLvThcEej92CRqzxW25I+OqQwPCFqMsIg1QsktJ
1KHik/UYr8NdgLHg3JzagQz5eVISOJ18+NSUJoQGG7lB6fAUhYOTnZvXtwXvPMNA
q2/Ci4VM5sdJ1qHd9jtpEhiZprr6bhgPsGfYET6uY2jQXhBY4dFT0RBx31miuSWC
n8CPh0mf5K1GvAr9WYP1wHSAwWyGbGDtzRhAkg2Ld1BbScduUZzbNMpS4Biiq9Ho
Z47I/v+u22p7HHT1secSIuXifmfJDOcbf4def1HxS3eCfNimI0hhZDDyiDNfGPJ9
Nli2arVZ9UtFzdDjDcStmOIRXps0nqGEA/ztypQtF6+7jG/KXR0ZfI3C+JkMy1gz
oI/UsCadUQj3j4Yp/aqorKNDLWS7Qh/UQZes4QNddvJbwyNXmM5xZKfjZEk80qZ+
wv6u6Sqn1L1VBEZNXFZTxqSaENodDHbOwkYgp79QKFcCEr8S2eMo5K+eTkWmdkWH
sZxhFzW7t42Bu+EiZSKqWp2NO+iRgJDUVB4k2ZLQGZAk99d/UXY5FBz3Yq+1QvkI
EuviykzEa9pLsjDWkO6/WhJ40PrCP7pMmsqYm+0mFjYjGPNa0/Tf9CnfS2oMHYxK
k/t+VLHhvlhLf8pqIpyNZpUZhxJ46j2Bi/ovsU4g4tRaRxPiLyCbXWN/NpDL+OXL
tDasWPoDkc2+egsDmokENNDFhXd0LrFbklvxa9thbUH4Fi6erHvTJ+WsBb3MSzsy
f7167JMwNvZ1qh+/DMQazfF9l0UY6NK5CpJe7tvowih+RpcCdK0NOGHTTQ2Ai/SD
dsfM0IUhzKHqX4Thnq8FI47c305RISjmVzxAYGqfj10fV3U2aYP74T8izqy65it4
vXh232ZJ6votjOfSKQOt5q7qcHLXGBDDWdO3hxMuzf0zjQJfERpGcUPWTP0wUir8
GQZaGPOWEevAXpdwP7a4ar9hQP1PRYU3ROWTokWGQQyH4yQWsBwK1FrcDspZDkuA
e4nrFRBxvvwvd8O1ma/fvjd4bGltyUr/EHo3PZN4nPCVrLgh4swFo0n9wA6CT3Il
vkv6nCejAQYRcHZgmTchyPnYKTlPj/ZWpVm4DL424A4dYHJyj0RzWfgUmVgNYUnf
/SFgYZdyqYhTcWRz5Tljzt3K1BFTA7TX311ktmvx8WSM0UsYSMnQ1QnyqFmQs3S8
yK85fICVNLR4BQDcvyVEM5N9T52dDYhZ+0wqmphIlum0ydL740eLhg/DdU8lhVSJ
1NxwCycm5Vej0DaqqQgbSlapN9u7ppT8+2ZCSP9+8mUUrcuZlW7RRocKYnTKZ5jL
UMjju2PlE9efAH/C8wkVm8V94ZJs7f4XtjuswdH47d2TAJH4b0uPqBw1kxMT6zlA
zd/Ko9qBZ0uyLDjC7SMZv3Xr1Qz6BirLD7CVflhVGhxzVtG+ci19UnzS7QjOz76H
Oz46MZwcQRyxFQdAFMa6oy86L3cBp4unrut2yv/FkLWNYRe4rPtDoTzVmyWXdL0x
FE0rV649ZZRhKHMpZvn4ozQoBJy5k3AG8zGYopjp/twM14RbIcLyHo1E1f2pGLis
+3dWnvqOWFL2FMCHNsohYsHN31ZjwYKLz0bk31VELIcBKR0uE5EQusc/VI2+a2qD
UpLLqFtoAgzXZrUOjtwgPckWReEGMzEuIJUVzNl0zXzgPljthsZY6xHG13FJa5W5
dG8vgmS98DZ34nGX6BJL5KyXZ/lTFxPf4nqY2Acf92FgShuAvoW6Z/HKnql0ALcM
Ehi4eMcQBVergFWlp+WbJMUbhLc+DTwClLv1hMjZvsxjmMAy5OpSQL+dwAnSxkkc
TES/sRtdbG7kMmLnfUYXFHM+5Yrjp5r40zoRf0Cqcy7r4l+tmHw1C5icFTM0ESPd
EgiDF3cNyt9LKMmZxvcxtw7zwAUkCaWFz4lULkfA6ntareCWeRejmE4IK91dX0cz
Fgbw0aXvfCNbKQ1gV2ZyJj/z7bg2IF1YlHxwCGb+eNOoFmDRBsmb5xMG/AOcXZBf
U2AOpOt6rxvM5teYcVbddwMQQyv1vHDU0oNGxhMj7YPdFd9zDAjnaToq1eklMLHk
G7oE/Dbch62JqRM8bP6DT0pFla1Wees3g9F2F/WOP6+TX9sXyuTZlOWTw08wp6Ns
YjvWsmmiXbtt0/XxpLEfiRixcwqq4AHE1MpyO5DApPNZpzvGjT1E5C//8pT1XZKO
7ZaALRAj28G6dLmXoCuHCZOb70lk1u++GMWisvwSe/pDnpOMS7Sj+lmm4jrlnVNM
9xpywCRirM5NUKaShhd3ihZ3xwl8pISD9qouPXTjV0IqbnqmUO0dY3cvWMkyO5vU
UD8LHEN7ZMxOT7sRqiVPnnqLDPidXDKaxM/hmUCLG+FYZSlW1VbX/XFhYkWJMsWU
XHTdxuLhSftH45OeWrJYW6LQinfVmwaW+LfiV8zQQv6A6zJd9vWL6nZdWDm35VLT
qjKk72IvGfipeivKRcJ1YiSw3k1mr/gGcgfWG2gBRua/Z/aOS3KAhXTAOAI3KSNq
0Dn7C5o1To4MMXbR5TRNL0vNOtFfGDu7SBtqhCSJ1ewMX0Q0ly1hx1vp16iRKjVC
1Xs28gAk+iaPR6Sdog6P+7a7V92Ee5jNXw2H3VhQOBLl2VFca+p587EiRECAoQzW
niBjINBpkSoRHnh8jO1nJxnlQxQYfvoPPljDV3qkPrbEukL3npPHqiy32kLIs2lX
gMfiTqYQzs39sOnXMw5/1PdOgFgT0bmQHdFcdQzInV2kRUAX+EKJP5OWBnJhyvUV
BJXywB693rtJXha2ooq7+ZIn0vH6Z+RVXlNeJPQoRTGdezVSG595DkxpAvMUoJES
3ne1bWTE6j19pnsNc9uKNO/ZarpQnDY6a1OdPgP9d7xMAes+xiWtH7zI40ELiAC+
WnLS6ZCBrzLRCH0aZpmnBg5pfoBKFBP09RSG8t8U4mosfilvEVtHaf/WIm+Iuzx/
iuSJraM9UAMNtVXYuyFd4HvtyCA/IiwlisJfdrK6cOL4fdMH43Nx0EcyfEkLtm9J
D8frNaYu9kqhZcm8dQAIYdJww8coH0u9oePgeSkSzdx9ppDmxpgp9D1ys5D0G43f
dEjPLiW8tvLtTlJn6WlC2kdBUqKp+UuOWW4s1VqKj8R60fRIKvSxtMKSFlyBig9B
GocDS6knY9zbmeZmMKZI1qBScKBDmeDzbmUDRgnr8wGm2xyoJTB9S7MX04ACqrTU
hi70cGKths2uCQ50KBtVxERVNuxTyskZeOOIMZKmwpUnfKzY5h6TrCZEAhVaCsn2
nxg2VZfnilUkRMSYTwxHu14x4zj+vSMs7PfwF5e76Mq7tzjwIZIJQDEsCIqSrvm2
8n7qd8IKwEO7hkrOtbPbMeXoC5T6by3DC7lcQS4wtt+mXD58CDeOsPFcN+hvhSeZ
3bopkKaEQI5osGf7olDOvDkFR0efkdc1Ma/6PJVUdXu81GAI2YwaurqYZxlKbv+t
LwIv3eDviOQChtfd7gpCZCupFfcLplX1fFRAfpyuShF4Jr0/n5GUctgX3FPfkV1a
gSC9UfHXQnX3/dZ9pI6dNVaIPWHzQWWdKjiQDX8Y13xU1BiCqfukuW5mYDQq8gIr
wywapRZw9fphOd9LjvLP98HIIfjVeCvVikdCzPz9zqZtm0q9SfqMPGNnRtk/9YKk
DMJjm1xmQ2OUiVElEz5YhX53x4jUwLFIwSWd+x9iGr1BzN/f3lieOyOImGKfUwPN
e6uFZ6d4zm3kt6E492TluGdkFs6Sb5O9M4iM2kmt4BcUNKljtw9UyZnpTZZ+RLSG
b+N7cItQhLojOrQnhJrtGPirvoDavNj1M/1GKikJtqxfYiJBWSBDhxZNdlMDnZg0
hhhvvuNNEjP79Weehf8rhxAeGxkaoOJSIB3XAAitAQme0n4WRxZ0/Wxdkc4UAsrs
Z7xaQAPDaJE31gWhGeWzVedHBXmGYeahDCifHnBAj+XELdz72lMbU34fGWRH/KmI
xdEMZesD1dZ5xmN7vc4uJ1u2morgTXZMDHhwM/HFhNEG08vIHYh/q2dNs5aLBXsC
2z/Bp9Vx54s/QFh+aNWtc+U8dw44oxAFBZDUzoA6xfC34RwH6IyYqc7cE8OmNNSS
g6wd/BW09iZgiVzyjjFPhbH7x90aKnyLW/WVaugn9iKNZEoQ62lx6j5CXXvpf54O
tcKi7Lu248yo8FtnWzfG8MoOoOGIu4nHt0Km0LREsZ5ZLY+8SiwhZ4quw2EDszOn
S/c/ZnxPmdW6kd/htUGIJJPzBVtCAccJLXvw0qEg/RVj/Qpkl6MA94e1ScdcJtRc
UgJBSANiv5mvBZbY9gaExz0SRrIUW6zksQApJ4bhKxVgxLgu7vjL9e5iMD/OY8gD
GMzkz5w9gaY1r6p6yfeL4ROo0utWL9UGbOT6Wi0dOSdbS4Xq94qMgPpY+E+BmHn0
KpBfeQ0MX/teT4pQUnNyAtmerddXdnBaO+NRiAbc5Iw8ldCSOOgqyIaNqi+X10FC
+EXQcd2Dwtx83eO07dPVP6/aRnG+kXaGFYNX1/P6bb80dO34WNEwH9gcxT3ajDLa
dCw7kfhwHmTdsTJL+ad5I/cz9kKM4+LIDTMeWMt1+ShnFzg6PCSnCDOd2mXPxkmO
WqbmnAJJTJuvZVAUpGWUMeh/PsjjtgIeCv6mY3mgclUvYo7OXgvWU8Zq9OCIfgFF
22zohmEB9TK2uLSFQprJSwdqwFF0+MYUhiZ5X0K7r+Vs9+FXnktKrDfzldY3vWbX
ysFzxbmHW7voWHSIxypCES5j7PzM7bO9NOu8tH5CBZts8PCaQqP9OopXutfE9qVC
OUB4LoG9IODCp6FQp89ZjHgVkRCcD1Hd8qq2VA6x+SRg6jgqN46XsXDiYrJTxnPd
ItViQLF2hko/Qu3XEWqtyPWJ8pPWQco9/kqEYE6MrMwTgN4Zxy4kn9U4JGU6S/yt
bs9sQ3wvW7lfaNT1VLlfzeOaH5ao0Js8XtOc7GmT+iIQ08hXuQOdVhtLl1ACdU3G
0DvFqSXvbE4zP6mjbkVMsO6HlaQG7rxeQgx7lprre8JiejdiUT7uPGrOvxxh7ful
ouFkXBiOQwFUC0sOqWtf4hns0Mru9PfL9LL15UcYzppPro/8m6TFXbZ8dYtYvKd+
ugferh8RRKXvNEbLRUaA88kZ8m6LPstioFdM0M6SRc78CpXFypzzyVD05lpa0mXD
i20i46U71z9Av0EMKrYahDEeaMBkT2QIBWeu3BDYhpXn5h8o5aDLAAkAGrewHJZm
DCCH59Y+OtLAqWNNDOoYhS82Mf7m8qDb8Oi793FjPrzDovu61aBbzMnL8ABO31hb
hh8jnVLls5piULiYByLnvCbLLW9L1QXxKfksCwq1OB1cboXn6exruft2pvPi2OHT
2/r83Pqh4UZooiSBW8xgeRFg2hYaWcTye/0aq97qeHlIyx+YGfUP9IKmLQhEt5i3
QsvVsaQXYLzhMF0T4feTzVA7Phvd6fgUvMEJlnBh53goFfBJyqdORzVI75xArHIB
kWiCspucNjYzVdRjfo98sT6zdVid9GoXRxFNih7/zrsR5aALzR2VgVhOr3WzP947
N5ZWqGk7fvHNnR56IedezRao+l4MrVURD17FR9hS7ikuZpfAwAQbnalWhGkc1dfU
1YrSDXwTtvRaGzvsAZ1QNyrdYNwXDep+mwcG2EOasIjwMrSyMV2Hmo4RO8L7ol/o
ng259lFs1mLyEe9wMLj3yxv9KjbceDNb+rrhJIKYGLETdw3xZ+eLNanBlayjPjUu
0NKY9FP7nVTqZ134ZSeM09kDmd1uX2bz19kzHvEITWPc9bbeGmYIkCBY9sdzzzDo
H2i4vpQA2S1E4yv2fHJF0+GT920jFfWyNxVKawpseaP4OFrMfOHz5Nyo+jAEaDUE
tTibjO9v4h99W2boNPb182IgVhenVHqEeEyfs3EcBTgr/tORWxSgguT6li/6vqbD
zZNAyrD8iBoi3j+C+oxqN3/UN+m5VuFMtfwfHT1uupv4RyASy8n2IPxPdp3Q6CqR
J65xYfREHqaoCx2bun2uctahBBt5rRNRga23EtspvRn++Rx4Mvx2rLOWGp6Mrvbs
ag69ir0sysZFJmB2kGMdN50XLE93n3/PhImrcZZ0hzMfzWnciLDqoVBldyasZCVR
fb4+QmyV588svHkechAWEB+i5Orpp4ITDVR0c1BiJJAdBqpFL8elv0v9rW1FtU9O
XdnC5qn8fVTgKt6CWuBg6R1TpZ7zz/WWl6rM54FliUafQ2rqDjJKHTPrtmiXFBge
EIzuZqJw+wZJZKRtlSXP8uF5BzsHw1H+q1O2N5WLeQNdGyDdRvkrc8FhHoMte4rA
juBKS09O250tp2tMfbA0u8X/ZvgvCOzNX40Yo5ceLat8YoaKZUD/ZEeqeHbAPKLb
D/VwWsrRliCBOHQEzfdB60Qa8SSuBMYanQ9f+kKoDoRYtyhFEJIKTn49Oc3050lh
jcCvtVnlFFxnfitgJ8MHPYSPA56DIpXpS0UdAby+RWhsbzhR5eg4xDLDcaEH8pKy
i19FHvd6vLJSlRgUkLqAhPqeu9fjZATMz+VanWwpFAK7NlUWWNCJvNtXo+rNYLB7
G7nWTixeecgEHfYc2l+fcwJeg03/5jja8FlJ7O4W2ofIQHDY8JecWJsTV6Jyz0St
vD9ce3712OPppV8hnKYk1wH07RgrCaQiD68KUdSZQ2+FVejJXpYpmLR+Er6haKpG
gDhB2JMmRyxcFfWOGC58ZXMoW01JLUi6l+hohXD6eSkf5ZYIN7rxrmxOiPYPLQHZ
1+JprQHPFwyxoKVEoN+GrqiaQ8afTbJxWocVS2y0c7ug6G9kYfausBeQ75hm3zJN
SMer6UHpsTX2GTyRUhyQKgK+m3isW0sm2wsltdw0pRwjZsnT/s1OZPpoHxS7TcmK
TNokrkQ+aukbvNqL1xLnfVU4P2Wuj+IEJ+HBp4f/gFG5smEjehla9mGylHsWGS3k
l0zE0I5PHB81P+lPB31G+EMAoJiGk5zGLfHbWu+3DrzB65vfADDRHK6WAvoeHQEn
+iVDrxj7/4QLaw6u2s+DTZRMAjvxsYJD6QQWQtf2ZxNMDjaiJHyQIjGX1V8aH5nP
XMy8IBdxdynIjG03Lms7n8O90sxVlog3CXDYEbqjFPKtRp4FMr7z+RRgGSmBSZwh
n8v2PXoQfM+RKLcQ8GWanvW4PDnmg3M89E8Oy8i3xQY7w0yv3vW+4fvMnRDXqHIs
dPNjGBt+zq9j/Q9171lM5x6tj9osvIQ/Aw/MF4SoH1KubvG2wHETYnQ1dbZS+SUn
8WkL20NShxaZGfhnAagD9n9beIPCxTvqt8HyWGtj1/jgvuiAGevuYV89SPdUt+Ea
abkfDCK0hnDeG2f98o+wU3BU5pLeV3RZaRhzRqgqyhIz3uzyrxNG+22u4FSznOm9
UdJtt+O/w99gjN4AHGOTltw+cuT9m2bsGNNCJQ5JssrG5hPU2ul0wrua++LxWN/a
EJDpN8cGEbmHdsJ/1ta0S0BSqLp8QS1IoNBahcc0OQZBjtwAol0QxQb0jbJm/Tmj
1ooW+fTb1IeH5kNE3t+PlretIn6SYeaFVrApKJVz5M1hakFSDWKKCn+m2gFs3YZH
m4mz9kB5iKtj/P7xOuoAK1d1FuNp1yaeu+XnugPH3hjmL7hpaAWaVt4krCpZuz0N
jGPYHkkP9RqZ4vAwaP8WTAmVFF3GyYNSXRPl9LKGhz+DGUZS+F6YnL7GHVCHjjaG
6tGk50u3WWgn3vztKvh4/1mjPxq7ch0vjThGBb68Lo54lPlpZqRTNUjZZjDWZMYK
d9EYM0Rwa2fMq5eBNM9ZWgw9UsgE/+d5xxQFIkJrMX37tK6uMt1DjMvuWtpSv0+2
A0mgP92LKaNBFFerkEaOWyQxXs3gJZKGCBtXHSDxm9cl3DzwxIER2qE6CaAw/Aa+
ErFZJy8rQfzM5Bh/3SPaa0GcBCR8+RA1X4YBH9P1uwhksUAJT8Feb5NfifhveH4T
BcleUztkn3TtLowcP/RG1bqAeHoRj6jHy6ZTtBL0cbfnh1srAqhS3jGpfA+kdNxM
0T+DvLtWzp+ec/ZsdvZaWDAZKn5waEUG4ujFgD1sQfjyD+WdNeiuCM0gxfbpVpIT
kU+8VXrGuSlb01E+xK3aTGWVDpMBnckqCnWR0/hzRipwxmMoqdDsx28WpGR+MsM4
P306N9QCkOOMnLkj2X47U7MFqJfPMejt33hn+1vwq2oqBSDh/2AcG0yJXh14V+3C
elf+U08V2FfIUKBYxzCjHIZ8GccPUp/XdFvAHppvLdz/CBc/8v90WnkrUVuLdcH/
GiFdoSHRTqPQC3WTx1zpoBodCebhfgtBV4EY9WabN98jx9bCFBDbsf+EYI1N7NlB
jR3xTTUfnKGLCAdn72ENIGHNjMFAuKkunHTknunjo6u7y6PFdZvY7zfy5ta7zdQy
K8/4f4Br747U8ulHGguP+zu4Kuxplr6B6c32gVkzJRS05AHvRkGkrbChdcJEKpQG
vKHSUUlGymcy/NHnhxrN16m+sk3U91szjTWqByhxquhuNqOyOX52hwMDlJv+shcZ
Qlf32Fb2LmdY3sNuejoZkCA3LaMXskb//Nym6ox7sFwcpN08G0an8pu1dDJxPlMa
JQbzNnvHsXi2QsRqdMz9JKDPzB0kClnZmls6DDNthuaKrDppKeKPhxKd1ehexJxJ
Mc2tQuw98TclscZHvJCexL9lHnEAdUsPee7CZcrQAfo0NRrUAg2H3vVSaQSDkJyr
g7CXdNAbTwNUM1ZlrsGxbpDyKoc7rlWw3SdJJqvSV8GKw/YCP4faQJ4k/AUGBybQ
uFmx4+mgYaGrdENx3TT3c4yxklhRsbmOp8sWAkkEqn8HmrkJon8Rlebq8839i5o0
iHDJOR+96adUNwFuBMBhRk9tYSTi5ZJbri3TUKLrr2//BCGwaMyDiN30oW215E2C
xBpj1LwPmCRhQVQpcvIx5X2lfdQ/K7HvyLoduCqZsCZelggf23TKk36GDGr9mn+E
uUR1mczmnOIlaRqWstzHHsdieoB0BcGgI3BK6PDHq/qHh/96SSXOXBMszmiDNhCF
DpwY0ua6qDFEj/gVzWrWP4ws1jkdwfHICn7r63oHD2bugnfxbubsGErlpX898s3Z
PLZy2liuhBRrrQ6ACsZAJj30uhDRLYNkXrFQ/yO82qxleza3PxxkEDXLb5DvDKGm
l6pGuOo/whQfYQ7co1Najft4KQiexnCmb+68obvMdTroPmD9BQcAl6X+05MuJmGm
9DMEWIeueH/Q+g7SXk2kSf0x4oBq5j2i25rZksXt96Xfk/WiLEpRk9db41xE3/V9
RHDwHuJQw1ZtNn8H8dcv29HhszNJqQH4fJ31f3R98XIaLy1C7TK+XlJUn1HYbZ6Z
RiNkqDAyiLd7lnvjHmqdnVE0q6Xug96qJFOLxBLsj/s2gQHME7a3Q2MDg3NeTYMj
wWmC/yTUYIPZyFzuOxaWzJ4aysTHJygpIQtoPrdws5TUDGXoXa8bvE5FL/XrmtKN
LcGeC1bbcYLOrfiSJLEUOOaOV2VDq0XgERWMJFYTHMW9mlsheuymmDiI3hT3IE+n
jBR6dfsf+/9HwzS0Rj9H+oftuvsNMTXIVXefJ5anE6prMAvn8pkoNkOPpQ9Zn9Uj
d1XQXbRyhvrVtlOiRsBP4F+RakH8TmzLkFA78Tj8U25mOVrsoo00davaN4/XAHXX
F2+jIbwruId29MC64Ty8ehZ1hNW+JMoZ0GXzia59gWa+4QTkEqBDUufohg+ET7td
6d+VrN9WZ7mBhqcUUaEPv0lt8fI256rdyUoAofdoYuK/rKAqz1XzUFefb8D1KRSk
TBPsirkaJHE15PaF3QIZ+sQtM0ak4fSBtL0HgSG0WxGmAn6bvXqBpqFrh7jaHhMg
yRQ/XncuPGs3A3HGUFM9PY5eQxsQMA94u3ChD5E43ymO5ziA8lpUI7cC9bO4KcOv
wMW1/hCB2zQRdHQZnsuzXd9Uss2rwvuXEgTDbq7cwBKrBKAhiYnCH4N19iGTNB0W
BMI3D5c2c/pwHfG5eu6tZuSB3UEDvI7X9uBgxavzsJvBz37svCSOo9r+6AAVRx6+
/hYic5DMGYitdEpj2IAI4hXIIjoBFbEK4lNCNLBb4S9z7zTOjcMG+7h8UOW5K/Qa
Rd8DqLe9Qdi0uH3y3tMiCzaJfXzoaTOO3HUDpbd4jjRxX5SqgvwAeWTj41cimxUu
51JJGNMvwQq8ujY6xZ8vab2Xfygj5hkYmpowSsCRURrC3bNkrW2XykOoi7ArDIhq
PZQgq/CbMQIhdI0U7v6Zs0P6qsvYe0aiBj7aYSqf0p2zVAaOaFcWqQs01NWtikz7
+oyAEUXv9xJyhm8wOqTPxPeS0GshBqY/3NHINxi2Gje2gqJMo3w8vBYrccVyBite
UkkHGri5GC9Y3vhBT8p0Bxbrvvtg7Ex7Ek1bFEHxw3k7aWLC288LIeYXRkPGlkWr
uf6R8KpGYaFEr2SsAxYKx1G70uU0up+uGCxJrJP5Mbu8qZbX0U/K3t1cK8t4uL/p
OEgp8f+/bZf+aPlBP4H2tl2m6T6cvFy1d5/v4atQ5YmfFqOjNY2UVrsgQi4aEmf+
vl077FmhLQty6ZpdIVqKE6DmzJBM9F8eIYo++mIOF7WJPi2cSotoDEDxNUj7MxCL
MCfo4Ad3htw3xVig9jZHb2C7iXEDfvNADjBQN9FecIfnJuYRgl7uIjH5LHCoXLgT
GhCZaZGDxBZB4/Czo5sSblJgrxb9SNMcj+RPdzXQtVGzAujgpZBWCAPUDSyV+Kcr
VmwO8S6unXu+0qo1Yigs3RWj6qKQzP5q6I4GetMdi2f9X5bs9LJn3Pj/8ltbz0kA
oijgk4n5hT/C0SzgblheEWgohJr/QcnVbBVX8aTLeE/10v04YrCUJds/5/uJWnCn
9R0k5r6cf0VBU5D3sMX1Ug8Ohh7kuuAMRxwYZ+MCagSt4wkvw/suxVHFsAjOCqYQ
31g7gevAiLxSnVqBnG8MsQoPW3qY14Dxyuhdr248Zl8mvBUxIMHZI6T+NRuJxNT6
0WrMGi8TN1X/K53w+Lv1GwyrMbKK4xg3kVxdlhOI2lLryU9v8X0VWAjWvGua2eG9
JWS+VwICBW5hrWX5GtKYRT5m91wRUIqs7Mvpne57Oan4jJ3VeeTDEqSJ4Ony51YL
pRpergq94Dubsa5aKqi0jrOLxfEatLH//ONZukC8kRz8b5T/zAk9vwmSxxY7dLQB
DMupGcWZeo1c1h5AZR8Ym4JzuQ5vOabWZ5zTeCufU2mKa5tB+q9kXGmIwygwGn6R
FtNpvuk2Ac1d5NeEYYGkRY4JjDp7Ba8k3wtdamGRgnIcZaaWZ4n2hiLNOHzvMBJw
ZNFKI1DqCz9GibC757P/P3MEIb+R9lcE6HlWd1hex+Bkk+RvSVO1AS9gR2DJ/FYi
U3OB8ynJ0kmybNnrC6MF2Hu/BjsSkUqXJdfH1xGR3/mUKWi+r2KmHNp+iqhgVpeC
vwLn0RnS1R4cQHMAY1mxgOaqGKwBnyWnqkK8al5h7BXGjwdqsOw970V66OoiWlsc
OA1G0qbge1/1vU+7e2GTtPucJmKV0YtYl91wW7cMPjS0NCJHiO1V8eqtn0BoMDQ0
vFyl/gphxllNvc+I5A/b02GahIEvwEHNY3ggPVbml39/rrlbyprM39tiv9dn0Nic
A9acIQrMWnPIejbWU9roWs05AuImW3BVZAVxwa4jO1j6wqsnISlU/S/lUItQTTyL
oRMKmunUA7pDK3Qi+CNe0RXep/ygmsJE3xGPW1Wdy2a9nvLfD84HX8Ctys2mJ1dq
+FDyxIM/Zj41UK4zXGyPYlOM2moPqin/gsKixlYRVvTJuD8vL9gbhIRXZblzEDL3
eBCpmR/WHlApfGt6u7Lk4se/j2lVhOvAxo6/0plBfs8OFh03BOR4B+YS1Nt2utln
9kFoq1zXr2NTxQ05bZBgO2BShoEo6SKgdky29rCb4NV3NKhy6vyd0RbG0IDvz2Sh
af+TlSksjiMybOm6yaJKISGjPrF7MUh2oCxf5WAzhFyfZ7XFWSVZlzHt0iesY8Vc
g43BlaaXKCZuW2sfB3DeoaUTNZN/CKj5dCCtQHrIgZcjSo1iG7zs4esBVZBwpoRY
BtpLM+LNIGrdEvEw+sVgOON0AjiKIxs4dJGpkkHhIY2yc8nIKMy4KYzjwaAUg8NU
sEXIcDnG9XJcVaVui5vaw+/fPRC9CHEyIzLIbJ/GOK+fK9sdOyYSVVmJZPdkhq4v
KOS0vB43vP108aY1+GDC3Kz0Yt0BoejUS8TtPGoJ+frLzbr3hoiSaImfmg0pcT6G
mM9qaGmPF3sEFvUbGUU7UO553xpPMGEzDr7rM0z7XOF0PELIwK0CDBPiMmLes7jP
38BJOaFxMDRU2eErCstg1ksaDmO4CDqAP0Q4vhjFDC9yT1kSBvRUDlyEODyW55U4
5zvYQ9EcL++wISsD4CtCb+mkMruNSpbVPWYjaE3WF/dvGjDPUpyNfUHGN3CUhybH
vujv1SFuNzWg+Xt734KOWdVYKbNiHJqDXKSh5+bAep4otWi+pnA6KKgkTqJdEjks
4BUKn6jQEgYyR94bPOrJHUqGndfSlOsFxYyyWz1ptXEXjztgNwU1Eu/0UfhP3rEb
iypWxCz5jMpIrQZtAMS07vQxvo41qW2VjUUnJy6BsWTiYtdqqzdB0ln9XcFgSwXK
nzZVZJmrFENm5YdnD9sQXKottMpdEOlPnVVyFW6tJmSVPX60REUffAzFbL5YJX0p
PBLKoD6vHBVNsPGBYaGg4jwwqK9C7eFek8J1QTpckHG2/8/YMhEfG2yFZ7TMeuME
Zr4lbirAVXg4R8mYILNw4Bb+HEbl946dY7dWIeJaqpnbiVZVcqMuvy1ihRuc9J8K
AP+3gsabmZsxsDrwf68JRwpihA8nJBFHqOIb5dmhKrtnYcrk2VvBtqK5e1DgsfjD
Qnml+OR5tInGUvDBHZDkxd9WtXnxQG7CLOJ35rMEwtVjg+YEFbL+cTP112wEfGjo
oTh2vOCR+7hU+qNuHOvykSQ6FRcBKRJ0ejJUN5teMGDqTqaA4deaMt5rJYqEP27F
emkMGhMCN/8cv+zHB0loWhz8o8FDd1SzIO8B8QSpuy0IGtohvm4VwHv1lY8vu+cW
TrRSiV5vz5xKh1O/BepHfNpF+bLp6V7Pp//MbtO6jgO2lsNwvpA4vL3e1jKrGFlZ
gzkFfICvU5+gy/Rwcrgzpn7HNqPjWRm/tFtu5ZaIKlgKaFpAYFQwhEhHjwaFcPkD
r75fZM4EJrYfY57+DfL/k+brNk+B1dVtRd1PNHa/+KBq8NRrmywkMq7XiAZ+gi0V
hfPWeSNHtFryLjT5x58YYXHEOhYQQdu+uM5gR13Ra5p0CZfeFtbIrrAZ0R4iy8aJ
ymNBfpK4Q2Y3Gbp1K3gO3JOL8en5bJiSeHXTl2Gp8p2eZYvOVoKItRzp0Ih83qyK
1ApFYsyypyETGD4gs2zby1JYrRvg+F05+oG7vQS46y9DVRwiRW4LGExpQayK8G6u
9lvONbN2hkRcjnLC0r29sj2N3R2uKWK5csBsFg3xVYHVioEziVvbz4bXcRDwMDWZ
0mFWZ/EorhFjXtRWHI0ih0Gq4zVAqHK3Z9+T+R8QPxh9MRXygleWL3UQIrqExV5s
DNZ0ZKcCK4C1r3rRVwQlOC0oPshJSJs+hRPlVhTOymvZQ0vI25s/YnZGfpgjKab+
l6OiGqB88JJ3uTtWSp7WNFy5efxEu8piLGBLQwBDfpFGHy+MeVi/PAk+V3kxHiJs
9vpWoFyrzy0BK4rnVybYSZj9k3lsEzndOPdXeL2g9Q6eiQHj/wydSspFOZfRb3HR
rnop/81cQGEuk3XAdROmTQIJINTO47AbupLcexRw0TFJ1ceqwtE/olZidAMK3wrk
tJM6rpShSkcsxkZKPeJYg0BtywrtcCkZ8dYgmMkhqO4LmBhGPUyf45cauOSG54eO
XNkGYu1fTF+8NAvCa4geWs0lIvzyTsyAmLwr6V93pYNd+03/8a1mv6KILDPkdXnP
AxJbN6yEPApNDp2ATTeEbFxhbDvAj44NREGsvgME12ChFYCQ58SaBA81DpGQIuLB
KTWACF94UEDUlRced73Z+hKmkIW5CpyCH1V6Kgyyhj/oea1D4hBBnegyxiLx9Ids
nnmpgiMXITbVbPWDrug5su2lh74QpiJJt0kxRfDrl2kt86ch50P9sA/RH6YJNmOy
+muDAQchyB9pFmnTdTPJItCZr9/RZXxzs9iYvs1+zQN+zQMf6uFvwEGyaLmXrNjm
CSwN7CPde9n4teJXPZc8v+3qZF2FCBnwAGlrTa6UD6fhWT7YjhmphsA+B/99uc0u
ZKiCMXpwnuy6sKL9/AD3Mx/+Av6wJHFsvz4FoEy0V2odV7d5almFlm7e5PzQ/ShU
qGwd6PPtcEo5DQdXljKK/gOtxhgxr/Y6GbyLgtN7kL6vkWZnjGdREb2JOllxwnRq
ZjdXXwXePhyDuJVnHWwqdhMYM2AECRY87iyzg+M7wRB5hiNEQG1Usj4W4I9n0dRJ
9YGC87oOxnufD1vjgNwXHbCRwuxILMZtgDH+sS0Xa2+otzBU6jDiZmjoP4eXQyF4
5zBBIBy6ITUfkJvwTkzz93Z2AWuz3p63lBJnpmHMKlgeno0DrSAGPuDbNRY+xRot
wJyU8fxIen41bWxUnuhriwhVZ+nh4KEd0M5pPnkd1fZN1qE35P1NAWYiDirM+dO+
OnMqJRute8nZFIWn13O5JMw2Ns50QcKv5RPudQQxxxEMoifdELjZwLkwTpKlnVLN
EbohQsLCRU7mPXnuzw++/qUhEbO9AoF1k9bOusZ79xWjnZm19HCMhIt0/d3sAstF
heVLXuae+jm2yVAQ+/HMwLMSNMBfdiLN1OYEhRFoJEKCXcLcUz4Q7u+an79IJXQV
daxMSICFx8GcOqZ8apOrHwqicjVZyWh7guiqf4RxHLMHUkOuNCDhq0ayIpK3ma+M
BsFmSsT3JfT/3rZBAqKgcMEnftYwVdX88NFwHTbSQR2ftiozOxpLVWq7W8O5YTKA
nwHwl0wgbUUVSlNbVFrHWCL3MZC4BSRUuGddEDyYKtzW/PnYizm8mkuHkD3lakfa
Z71mxxUE/jAdAmNCo4qkfLVF1gF9VP3tjWooTKeTTq+s7FK1FNog5De2QXKVNpTq
1c0oNvhapi73YGkk/uHM0JwruisA++rerXTb07z+tmkFM/sYRwEg9LPOozU2Z1pv
W3n9yte8LyE7e6Luxg2scTo/jYvkkwFKBsZvnoMyLHb6TziGislHENrwuDwhh1iz
5nhfRMT2dBSF4PUJfjLB6qVt20WRBHS63YXEDfDl49h5RG3CSQ0O49zTukywjV3y
ahFDF/vHl0AACuklyik8uwnoFjVNY5ddzyEUhUSwMjw3GZqafu0rVJVh5y7zPjUy
1rgVCG+qk8yr1qQp1jx1vOZs8j43MrT6busOVwkUX6sO4EsJFdAqNRh8uA3yKk2U
cWSigREihQ8MJgSWqNiWe/9OUbYyTIsQ96mr6aqQlU0KyvNQaI+SVwUiTGEHXXzG
MJWGjXHT9drISyQwpbOzY85nZ1EiyRBEfyxMiC1TOXglUg42cRmAclg4cEYj+Txw
gesRzjlZQgMaYkJ4EVwko7mqP4beVi97bRIWjPi+9RrkxvOkZkHYRuPgG8J8SDgh
BgszCf1VfvgoHuPO4PHDOlOmGAiCIvcJbb5j9rgAjpYSZTjOqCNXJeBLXn1KY9zY
KmVyzAgR4HJcijpmyz4cKvYFopNIJ+6MthecuouWcG/8Rvwv14RIJSedt1DDJctF
S5EPqPEKsRcit1ngr2ZOqHb/wSRCMI5ddOTFVNicvSiF7jLOzRgUfAdFtoZAKOXE
RCMdU3ToroUXBHgxFA1vQWr+jrpc7C9V8WcObKufeNTIz1VfGUZfvpNDJ5ha6qJK
4IoYmJv5QEts8mQiR3bJXwR7+vODJ6VKsMXatHH34JNsROqLNGDgg34WGBR3zecg
cac96PIVc2Qz29QWo1VIaS2zF9pWzbRBHENmBUNcwgobBf7tSNHrAFwwc3PuzSKJ
jOOUAtxqdQqCswJJQKOkdOOZCEmVHeOyGoTVUdSGnN9Sn2at2L3Dz318h+BnLL3n
AdLnCsVKWDRHTJCFJ4jXGwjAoWi9oPGqC91V0W6U8QT1QSuaBZ3Exl8w6LR1gPzF
QxuDQdA1BAp7qpOvj+0k+SAeJEHYFrQVqvIU7lVJYAfxHzbpqzA+AbrNFZON4Hrh
uiMKqYvbGN1kmdAZk9N6mFmN2cDZti0hUVHY5E9HsCSAJvq8H2ChoT+RDd6z3x3G
8VhU9wO7+tx4Ah6CsOUSvBEjRgDCEdiOAFJUZ0qouou3Em0dAhucxR5IMzR13PV2
a9L5Z8ebo8LNLMk/msfLEKU+im9k4DZm1R97FDLO4c1KLWiiFHrJcmZ7TQM9PhGy
NOrdzsVEdC7oU7SmNrMGMHJPCKpxe8E/sKzVifzOyPAH0zs5lrREmBUo3EVbDw3w
00Kh5wz9895HlY2iMxyI2k0mls4jvlW/fRutK8Li8q8N5zRFDV+I+y+IB6p9exhP
PJ8TObDeUHqnhWsdx68SFCO0TQ7HVv/eY9zNWYmNAtBvNBmbRn4EfQRdOuoHkl/B
Y8EmG+uyCyhZRmzfZ6y5zkCm7zIouDEWdB9LeHQlokwtmTmWYqLTqAGmMMStkIIf
8p/RiUc+Z1g6AB9ZiR6lSmBSO8g2sC+BU6bFQ2ID0hLYTKwfrF2JkS/S4fly9pvn
cjTV9AhfRVQo9imf6RQ0pMg/kc8c5p+/Bc6DMKEDSxNRqQ5gNApICyErD3NkW4dY
0JqdDxIE5zIrBSn1b1lPGRNoKn0spj57Q/aOaLJqUrqhLoLIFbADbZJqSLHuyDSM
GNQDwnRmQ+4ZBjrMLIQZmeGRTzSOxAGbdf+Bdz/tMRGRaczErW8A0/VGlsu1vpLO
QA9bhpuudsBcGVNRdSNtF9044rRHy3BE14GmTMESKFcBMNnrt11/kKUC0WH0D0Kr
xkyvG5b+ta/qkKiRre0nX0Nl/XvwDPrIVL+/uNpLDV05ibmjZoP2XLhH6/TPgbNV
kNi9WwjlBc1k0sc09+5U86CNnxXtSendFZqJNeGR8fLk2qF+CyilAfg4/8uo7owu
7PpBP11f4Bq4wJiEFHs/Qj1f7U5VXJds7FhtOUxeZuYUg1d3j6oYE7na1vl5j4rF
4/29Mk/di2qYGW6dopfwKHcScyIzHHH+TmA7+cM3GA9BkJeMDkJ3trX1IcqFJXmu
AHBktCC0b1KVT4Iwll0lgbNxTW54ocVS/p1OsUQM42/H7nUFfE5LPuahtRGqCWmr
y5sn4sEOcdTO3lKGFy5KdKP7yxrTl4PilrpXNoVziwErlaQJRnW+rbZHAyhgZhGk
wEdVNDI9gKnEyVcXG6sZmOgU02SaearkFRxFb+vcoJpFfE9XitCyjt7YkeA9I82S
HSiJORsSAUZ7LFe8CmcGWYDDbuLTonCB7OiXYo1LcBD4MTVhl7Pdd05pT+iBFQDs
yJkxQfZAxfp8SOso6NDrK8uBxBDIP0e+cupweNLeq+FOMiLv4ckuU420PrAEvdqJ
winlpojGL8Eda4Tkyug9HFRoPDOvXRJBhuMhtInk1O7wwlpxGtDubeG0J3CfRcS/
8Qr80uuf48Oa14CqjJjIexSOv2ZIQZIUnSXdkB/z/U3FM2TJrAVOMy9Nbr5Jpwn5
Iapspfjxzetzu7bSLhOyh3g6VvzAvOr3zodeMivwD2wtLPkvK6ViAK4T27C4oilG
L3X54muxv9UJ7xQcYeMjG1+bg7OpWmWACPDaK8APEEWxl+MSsCtZq2K5zZClBngT
kmxVjgx5/Yuo3S8w/oHsTO3yfLYQJD/b28Jt/rH3h14KMnxDJxnCYSJtkGxqNT2y
zXeePug7oHoNloZTlIH/Td2ohO2GFgenT2JiIyAM8yuxfbibZmRcQPL9i1HIrfvo
uFJlaamzVuXbl/02BgPwQ8M8C1dwMrTUAFOJSrqQkA6UgwHDfOPlbtjOdnabSyf6
Gv4/6F3zOrqhRHVBziKRa9Y8BuPBqUa3leXR6z/4R7TKejwWVqczm83OSAgR65PK
qJtR2hw18bVFhD0FaaNJ9/FGK5dMIlRfwaNn2fYcWWynkTpxVizlbm6zd4VAUYGj
AtzhXgczylwEteWPJ5gsUwKC2cn9gMN6NkmRjKGRk4qrayVtesKVzd8jTs8gQ4+Q
PkfQsAtEKuixY9U4nDBD2EzNapyVYwB+gh6rV2wsJkRgXVguEtYC0WK0r0TVGDjB
m0vdw9xByam+MrBYMI5B5ARTH6pP+HB9WDfFYOiUJ0Wmu8zvF+pXFHvUNEuhP6nT
7kVIR/ixV25NvYj8lEFiSIa0F2J6/8F7IeKUCqnkxrW5bA0qgPgoTIZEMzvqAj0W
DjfMHs/6mPvKDyLfbk/42ASqOEl72EL3ewLiwgurszPreL+sWWC/7dtdCPlELQGT
Esb6Aarq6tErxFiKiCrkXJQFlH+qEdkJVnmMH+dJezWu7UdaoTobkHSHjvVPQgWl
dvNPa0ws9PvF7vRqJUd1yDxgmh8jfTYP8aCbpcLHAbC5LfS10bYtkHelNq/tyiB9
E93xGsJsuzWpv/uqwaRHv/CKPqGBkis+5Y0Buj/Q9Ls7lPN4TWfqwOQzC8LfPzQr
89eMorg8+AZnp1Lk7LleuDO7YNh4DUYZQdhFQEb2WyrQGBJ0MXOBXr4aL0sFRAr1
f1CyREkjimY9uLF2vmzyChMNRoR//xP7BG9BbyybWXPAZeW4uly2fHuUNXaMTiil
nAYo9b9MJFEXKPFwHmbCOI/shC78Q2muWMHfe9bxDQxh88YYTuWgkCToJ1CPPdGU
wuIyyH/EjNDCSxbaWvvufnlaiK4Ek+8S7OzimvAe9C67qmI3XyHBh7eXuHOD6xnX
Uzh8FUx7ALLwr42TJRfq80ntLzGnWeVCJoqKavwCDSmCD2Rp9Wip3a5UAlWmwqya
WNIiiPzF9lWnAhdHVAJ19gdoGezuKQQlIt/dN7VqKitcI2NjAeHfeqvBJjdJg/wM
zPgmCTb4l+WZyVTf3Ck1Z3DpciMSmtMSq6N528NlHsylH1dNhtRh0W+IFI9eqgsD
bX992MZvlH3qXdSa3PV3uFwqbCicFj4PgCnaCl7UnQB+jSEtIcN4nZnHNWEvWvX0
5rTY7v+TwbWaXMIVKFzLjAqB7DYwRRj82Wt2mgK0FLLLNXh0rwqRc2xZOLcjhKx2
uINnM+Rc6mliIJpuLXji2Oq9Dt4hEy8q5Xgjo2mV7zVEen8WkCbJm21G6vTMjzAv
5t4vYNTAISTJ+Mx9s8PN+QVJ3OxcLQ6FcLYheZKQoW2djqMcFZ1CWQ1zR1AiBh4h
3LxaSJ2IwsbUpfHPydJxaznTQR8pMDk7D5on2uQFEthCXyOaU9Q37W50bywaMyJO
WpuYNocarLCS0l+Ozi0NVhNTTfMUakPfHeRlZWTfl8iUT+q53hMTNsCbYjP/R+w/
ePSJ2YBA86oWQmS5vCimI6b7yoW7aBbXlbVFBpoQg2QrR9LUCAWGDJPRKesNS8k+
AXqPc2lpEo7MOUOlOKumGfM7hccawhbL8Myf9dASKb8p6N1qDOvoaUBoK0L1vKRv
A28Jc9QrBf+sfnAXXBz2DSGrjuiEI8FlnrDJS0ws/kU/fs+LT5N56sAMF5C5Rysl
3cEourVtMEhcrPeaqxf4rnfjbZ4nuN9qoxYAGUaPArPZN668K/QzwuBdqolwiEdH
5CKCJUv054JXj3t2vTnCaBQPMAmDGTXMadvYZVtjXBqLRbqHM8ae4OIYD13t0itt
1XgRaAbkeyeBJsmZ7DwrIXnWSTQyXulDW5kTkxP+/TW1vEfDIb5RbWngoXUmdvQE
k86rb1d3kWvtYf5uJNx/iPqQOz4/vb0Mob7IIOAYeMmIMBRuWTrU89MePg0Byx7B
sDlnFJUlPWvJlJED2hGKpZA+lX9BSuGBo2yupzEHV/lqYFvCoNAnsr3wHmyltRsk
AZ1Qe/ACmxfetnC836fZNY+EoXbKmjxGlWpt9fWGf5fJizhURw9ZidaD4XUTO3yP
tAOjhroy9/I3M34rwL1QMHbIbG/K6FOduss2aRVOGZ4Yj5NeE7MZtFmvBF7fC4d3
dX06/RvwEOEAwVBVQAD0WNKb8npoNrWs/uD0zB9x0GkSe5JDpLfoqkuv0Ke4jmUW
wDqY+zm40umY55bZzkPOImfKhneYABBh6wevdPNKLKdS7MFEL0AsQFgGj7nBMVF2
AkaF0w8wxDVNMjLvkXhKaBdjOYsCQlOswlf62qi3QHfvHRDgEQ/E4jCsyyX2vJTY
2zmtcklqZ1ZLNxDJbPUlcuohpinVPmd7pnSKtdcLbibMHe4WWjJfgRRwE73QZ/MH
sh7hnEoROtdobySKm03Oeeq2kfCxx/nyWcpVMxSb6tLnsVswXc729iT1bamcsoho
Qbh0xOXuXmvgVLpuclw+LV2QFHsgdXCynqqZ/ScuYJ9Z4njEbkYtTyX1Fd+GRvfs
si3pJp5ERpOMqalALAbwh28eS8jdZmuxU5e1uf0TcJpwrLzneMu6HnFjVR8oCS74
04Qt1S4LFKXZ3e0sLe9EOqKuGcAi5NSvscbLOGqpFfJOIWXyzxl2EQa6sLX/sMkS
IYDfBDhy3ajVQlJGBnO11MjZGH6yI8N9yPx61M5cbcYYTsTBs4V6hmS6ggCJXZ+0
tAW2ky4oUUR1lTG5tvGZUN+5AJQ/qQAwd/1foSlOXANYoVBYFGXzxDPDAiLzX+mz
EjkzsbtDSOzO9dI/O1qamv3RslBOebCQjaHSYyjK/9/Tvr/kEQuXj8HhnD1xTjZh
0TfLletxkpYf1nopEd/dFNy5ZEZnbkGQHLu4hvlETfzvpHZqKkwKk9TKbuA1xnzm
cOydrA1cupDYIGN5/6WxUA1zm2QBSlCiSfp1gqa5zfsMJqxyMLi7HAT03SEfbOdS
v/XtbbGlfkYyiPxpAfJnlSFriWhAMUxKYEB0KHB9z3tfSIkmMOXLb/8nDyrGPPrb
T3s6DaG1LO6IPtp49GYFRD1OP+Dt3jofcZ3/ZczM7y1v1xrbHE61sWGKu/aJaV1c
+IXW+cc/yCr0+ULPgeL0F79eK9pj+4qlvYO55q9xc7IUSAK2wb7elJ/Nxhzk6SSQ
6o9fMFNXtrKO84h0rQG+UDQPETGsogpJWLedge0OpbZc099AXbJz+/0TiSPw5ZnL
0BakKO5bG+xXZi5quWju/lCB5vSOpa9KGotlEZNCajO0/8MqSh/24KF1wjtBO2e0
icQ7cOpcx82+c3oIUBz2rVUEF4loAGQJjKS6P7vjpFVbm/ulVEVcPon9tzYNdrDS
O/XUHwUR4xClPS+A6ZQc04EwiZHZM4tadEBiIblNHwAHHoqoL5x+I8KVkTAwcXTM
ONOATp08YkK/U9+TMF9xRCujDskPxhjk1tIo1x/j86Ar1roz18XLRBNg39uE+0V/
FZSbT6j2yHZ7LJB5SHJIiVn7Fowrbp2xAKUuQQBzaPUQwAzFgoGw0HGQu2nyaOaz
NtkAnuhEaJrKjWHi6vmMBOBUVzmjXWwzaAeTQLLYA1vsQVdaDxf4HWxHlJxRu3ag
Ypqhf46oTR75P/kQN3fdBTrVVbaL/GuBbVMTW1LThsyV5xrcYFL8cFAmwZxI+IQx
lPl0ok1tzr2ZkZ1AohlpJqWEdOEHThDdSL0kpwaC+cfpvkm+6WrqSAGT4nXN5QMB
0tszHtDU92FwJMAA3tdDD/aivBcK+q+zjwc1iDAkCbq0wHmYuFSdL01KR61NUdB2
RrIGuYVmODc0AiYrjBGcslxwj1FbnRg5610EENdnpHMsF30TsJNmw5wxE5QN4tK7
VRdfQIKYZ0DWrd3THkZyvrwEql5jpPTZeO5+AMxryGgRSJTFTXidetCe827K1Ak0
IfRO1EJk1yHLxjW02MWk2Gg+9jH+37XjlDUfkeAhU+to2t0mxE3WMn5v5rJADBeq
ip5M4gHXD5gjmNaL0QEHG0u6gUJnnloI4yhyFFUP4Vf9rFTSf4SHbR6frW4zgfpP
uAWnGpnYD24FnsdWjACYvkRKICoddEfn6yKiVFwzUqlI7kRGgTNnA55LT8LVD5Ia
F6DSGiMKchKkGZcmEbSAlBaG8gCDOlm5rSvihcGBepNeymqjxUG+aNA4KdPajvbQ
2LHMdk3dv06L18mH03tfdCeLXnGtVCQZ3hxG+LbgpZUKCnP2x4HATlMrcWe9kqrp
OaE/aYacm10H9T1SKWxRSLtcTgR+bCMfGeADZ45fFa9fdD0asuXZ8NE7h+qzR6Zw
cBuiHiIJzYzusWr7a1QpxChHCWko5AoVNgP+4MCrsHdVyPmDCt3NgCyofzlqCR8f
nc0TkwvK0bTKykN+F2vvfqWHBlrOImlZ+0IVUhvcFN1ReqVF3GdewiPfe8cVtOus
s8m2H49eQEblAxENAVKEwZcJGk+F4XRB17NBYCx2P3WKBu/5GClHzj2EIyHLMFZ4
wa5XUXRjWyVLYHWILUD5PH4ZIe8FMBVzL7Ei6t9rwSJ+gw00FGBkZJtjunX5Fug8
Ty845WxTVftoNvEtOWQuTxfWHUGa3TraVEp/CYHEF88mBKxiDleKyYA3tSlkmFzY
GW4IQwbeM/HLY7moPcWvI0iWOG4F7BpiectSyEM0BjFSNtKkSCaIMRKSdExMCj4i
+dwP3OEoiXv0/ySa6MDNQNjsjd14mUOkur+/ZK2q5x6BaHkRSSdk+cYQg14tJvv3
0rXF5h0g9anF1/5hyHQ4ycohf4t86sawlAxFj6cN0RabkfC9zrxcxvbaumwKbZNB
6/KCzvQHPE0a3vivBKkZTECKpLuVUBk4oFNeMIcpUzoDiuSf7BLix6/eIJy5k5gV
86tYbzwRawZCWGCzGs0BmXEnHXwaXzd4D7Wnm/RgmRx2v12BCmZEFpWXOhqMxrBr
t1d9r3smH3xTRNwqTO1cW1IckDv0FG9uRZt5J+nxN2YakIe1jlMfHbbFOJgpCMdJ
YI1N0SOo1hiSdFiGo0oQJjkf9KLZtbsvOWiGfVm9UUN9yN/IXFW+MbEc2nx1+p5v
D8UYmPkgvve4XZ0JRp/BiD7Pa99MkOnWgHsvnajSGW6LGqhfsvI/DPnAOnPB8/Hg
gU1nqLMMQAhuGiTqFEWdQq9FweidS8t2nETHaMP/ZPUwRilgeIIPXbp/Xq8rD1Sl
YyFXyKBPIb+5WSc4ttPA0iGd90UjLk3neMwfhzhxejNHpaYq+sJXOcjlvaMPIKVU
t73yr+bC4ihzbU6Iw6Cm5e7uqNJumCdi+QNM+UdrPpI6bmqy5I/H8teY2j0myNoX
MVVBI+P/9sOWA5WgoIVGoSkbsm0rFL1HEucO8FzU5iTQPsWJ3sfkaszJ/9nH4k2p
dekOKvoPyN0n1W9w+vNk95jGU/zfmp5IBWyWuwsxAzMvu0rAA8Tzj+di3a45rBs6
JHmz+cx0Fhyf8YPfPJs5W9eeQ5l/PU80LWB12mJwk+hZ3MbpLHZklKlbqkVd2pyS
tzaVZ/wDpbXaHpjxL7qfiuyXAg5tAqR0Oz6iFhLl3uLsnvFp5scEkS+lTL4FNaad
BAiphtL2D/cqER3P4ZZARZcrflVBhICthY48RPRsknNuj6fzIKsyz2p2S1uWBxKn
ZhAj0eo/MbzueiJYugLE2FOd6Tm09G3VEmRMMXNUvwYcpJfwaMzRXqPW1NbahmZ2
7pNEJn9Rlhj+t0dChKC8utxGlmOxpX7uY4tGNNy/ePMw7xG6XJghQ/lZ952Kxs9y
o3kdWuEI7Ev1OPiKu6emvGhPdTtD0haHr6Xzgkiv8opln1+0yekHtUYED8I2vz0S
9WwD6y8hmPZ9IoQ7QNu2IRDMZv+Hl6hGoEu4Iecd81OMXtlsjZco+ieEMbLFf4vx
Ij+LES/CAYzyC6gbiUT712PZUeGGiVoRqdlgWqsS+DVa3DSPVrrL+K3f2+E/kc1h
lBWpVaSMPQntjTaeOeOKVtTWdqFRwOSefPU/6v0ffUbJlTzwSomT1nuDbZ5bZxIj
umhpGLyBvzwzS/ZcObz0gptc48M1khOnMspSz9H28kfAA/6Z2vqhCVRHOE7+EvKz
hCBN6eOWvFBGg6d9+0qNCFakNsj6FnLERmM8tNR/20KlLDRRMwQn98i2DZYYOnWI
tDipHELjKKVJoQSrCYSccoTxOSHPXacrQFBZYI91HOmTAt/408VAZ4BzLXChLNcZ
aqXUJogBcLPiYUI2ulrnGPCA1WN+Ar+g5xBQxs0IhwaGs+H9YpmgVF5vp0U/mG36
kdMkgkkMDbgVPWkkTGxKiffLf6fxC01OZ46MfKZzzOeU0FrKb75EHCXLjjkShXcH
6c3m9H9qrgtm/vUrRdtN4P4/gz8YxVl+1HmcRIbwDg+POUq4nCX/LL9hGdZYCR9c
kxl0qW6G/MLugmWM+NmYzuOI5zri6YZb8MohkiP1zleDEKHWMvUca9RFoZs3CAke
ZkDag0mP9j/DCNLhmG9ClLQZVRpbiZ9bkKvu7eNxHrtqk1vFOCp1m3/RcDow/Dmi
aHAYGHhbEbeD+AXgx2Ue2VIsDAj413EqzysdX+xUXw7wX3mJeMTKwL82wHOMbPBa
f1Fpp7afE3iyFwn41XFBXsjBBpbx07CAlYM5xgHgelVTqAMG0f+aqQZ5G/RJF+tQ
qShP0ANwCMIQQF2wRhGwgKa9wt3F7BYOZeCLJZ37dGzBVwMcXnhgw7aadQ5W4oYT
hdJ86ihHrYxJVJ4szf6tyu318r1VbH21E6oqXYKSwlWAQUz4uQJsfHvXhbk/eZu9
KtbY5+twoJXETHWeR0UKUL/65an62ABuT2G8ijeKaRu2QaorA0prMZLCrXP8os1w
sfplgjqXmWtE0an50JyHx9VMU9WBIqy981aSEMU9YMAKdgsC/aSNc45NGD/VMa8B
s5xhjZzdzKFGeWMSez8mBDC9tLidDEM5Bv1ASbok8siqBwo+iCcTdem3ewehBa/a
luA1c4pzxa6p2QoLIAxfih0fjUdHweTOUAMLuMg4YuNbc38DDmcIJjyn1KeKRdW6
XrhvSP2V5M9jE/VciSGMuwgLSNIBWeCxZwdyPEg5yfzjlum3iuCom65guOITfdYx
SC7M2gSTlpac0N/FA7m6Jg1xIPwZEgOF6J0KYpG119Wum0qChmzCWNvAxF7MmsAr
tnQ+Li+U37l+12OtnzAgW3iENpJJ1YJlWgUIE8t6cd6/4piuzwNY6WDyVbeQ2VW1
1UrKL/ZJBwKLJ18I9OlTqVRNC+qRGIqf1oBdnT+dPFIxAdorGWGvCHQywM+WWPwC
8rO3MEhSbbp/3Pd+HX+LB+/bP4qq7XVVJ/t6R+jITFc/gL98AGoqMjKDH1JS0EwO
wZz6Euy91pVs6nBzrD1pjmVvob3/+BXGRIrnUEEgYUJZK1qOJKW/U1pV6kST7o7d
opc6/Q/xP+e/KVBZma8iDK9uwt3y6m5zmS/E+ozPkzQ2zgiIJ7Q31u7vCACNAv/q
zkTTcS0qbvzT0ODPoOTNHAEizKw1YTrerht1vfRX02wfHcallA4QhxNHy30gjqsM
bcKDpOjWvXr2P2xTPoKtj8ge5AjYK2u2CDIXPEGly1RRxBR+sKDZ3bQwP3YJx8Lz
mgaUb9jssbBh7ZYY0yWN57acAk6HTPlPW9OCDA2zByfr9pI/ZYgY1NYYymhfPxt7
8E4QewSVp52VHBbk9piSZ7ugZACr/HawpeExpPbRl2CN3uizl+zNcBXaBH70kLMJ
9FYIGF2rwahWlP5PedVaBjU1v7S83uBTwFWBCfBIuZvrglBneEeYskLlQu0ZOngx
g0CaCxzR0ICZ6GfKXr0jqKwN8VGPz7ZiWsbRuZfWfb4uIk3aOzEf/NxhLX8Y4O4b
oPSXUYMy1h/wtZoV95ykkrsk2UdRRSHVqKs+KALuMXI3Hni3aDGku1ZFs5ZJw7Qe
T6rMd6VFoQSf99venumI5li/AqY5hyaAX29warnvHPg8iHpVhCD7uirtPB48SfBt
DobppSg2cpO8AphWZQ1aBfIfiANqSnrJSbwO5EZ8XzxsPvuN8yScaExL6xnm4n0L
24gbR00sSkaos+W2Dq7dJtk9oIOLbq/OlO8WzxfoK5b3CWy63E2TCHLQuIevGcGJ
vUmAbdLTHPxArG63fDqygFQngrBVQTRPKpTAnZQO9miKv9ExOlVuCM/ZoQuEPbGr
ccvlHAUzRP5Li/KGUuy77YiMe3yLF4GqJTmYI2LM/xqNmh5oDZL+D0Uk90zRqFWn
nG9kf6WHhv+Ap1LauONIUg7K9b2KyAh3EJrxxpPxuJWVjd+va9uJbsn6wP3BbjJm
DFPWtDiN4nVnE340OkcBRz4hyFssYDzjmVgAsMmmBeWk7KvKXLpBRjeWrbU7Dxoe
18BrjEtNLcE03R8vg4pioVR9lXuPqE3zh0yaV/oNoMQHKhvwY5yx3k/tbO7FpF8R
wysEmQyNYDanlqy0hU2RSRTFUF6mWuythJdIobl+97jfwINcubgiVXfTokOK9OwA
IWDmDDu3is7fp1zVjj7Y+Tl6NA97CKXAKWvjjtaHn0/EPVpNVD2mSACCZdQfRQGO
gSy/soPMJNv/C28dy/IkaZwikiAwzQ/MVepdzS7LiQkFP5ol/x9Ff2vZEkJA1/Th
WDgkUur/rX+wrCiAOYZmbW/z2/wBWd9KlA5WHyDPPziulBLr6oXaMxITcibhNF9o
/v6biNY4iTWZ9/UVQj8Q6JyaoOz4tQ9TrFvSMleymaWCXcI0VFKyqpG9nFICd29i
5nVvGTCcx6uRc46Bezl7ymg4U7KUulwh/YVgp0zFSHMieqV6ek7FDtTdVu1m/D2I
wqCLYz5r+vo4dJU89qpLw7IMyUq0CsSFk6NOem8iJi33g9GtQR3xOICa2U1VsCZC
hmMIiP6S22yzUDo331oreuSyflJP4o6LE3bT6FA5B7lVyrqisbTxfgWU6OOtp0Ni
D3Xlpgd1hq2sGymL2Te9pxS5GSmeonKvikwYE5WphF2FiNslXeOGv3rEZ3fLyfKF
MF0bk4j7nHTI98P3vVR5G2NIFuaWt9fIO+BTJSlRp1iFROv8ICFH64AKr9ackUGW
+Nz3QARQSEmBmZnBqqUe5ugRXlbur4XOsquhhwIvZ1/O8PRA6UEd0gETs/H3GnFx
c8K/eXIyq7bQtpHgNVbH3Rv979xoQrcW7NluEiI/ZC+K5jTEiHPlOhGMQfbgHFTv
vBhrmCDm9/T8tpx87IpwjY3GGbiWGki53T4SNJuyjuhUFz3bmtKMEteAtq/BNR0s
r1ok6u2Zy/oTTTNyzMOr0wRm9qGmZZ81v3QDZSY29pVU8avFyVS5Iq8ZRVXI2h2p
woNm9d3Z7IBRHQz2eZcGlaJphowpO5Mue2M9qqDPLZ6C1FaWSCzZD5l2pwXUFq5C
N3zKQQjv+B7uRVZ7WrUaRb2pJSj2jiKYpn9NWwGI8VA3+H1IleKlunxdI7eRkVdk
AKwezNZw7UJo54WvuINmmjkBmFGwtJ993iPE4K0x/iwljh6/3tQNizuxU1DucOcK
xxKYxgqS1girddbdjk6LLb8IpiNRxrfHqYsb5AeXKpsgJGgGGCCalvrqHGseTtuw
M3WfP3U9ryI8nzcEIUbb30qHppayU7ha2Q9k8qMUbl6fgCr8vjBeXAtqHR+BcXlk
Ixl1AKuUyyk5spATbhdHTOFliE8FdTXW2Pamq8KmHiQ3XBvTIL/2n/d+mY98AYws
X97EKB7WhU2QetTcaLOAAr62pSl752hVRhtHbFK4aQARQPzIYhl4v2kL0nePv+N+
3Ccr5NtNM24s7Qiu8lxfXBAZDSMyPtdbrZvj+DSfXQ1DGGRV5CP5u27Paz5WlIlY
reGvD5xRw2JBz/+vdwW7nTksN8Nym1VsNIegKCuy9F131o4kLqk5A9UccWdx4DQU
ZdAkXSjMIh5SrehXzbo1foLhTgBoR8g103VTlfFg5ZkvYfo4fpmP2OFheXO+YJXx
t8eqVVCYohMvFKbhaSqGk6Mc8FWSqUtY4U6c/y8kNQYXAT2Lb53H7rxr4qGMMWlB
Jp2ymMIavu44XFvE8igMUONMq39fyXqZMprOIk4YP/C6nkxhQsvbLns2RiTMcdYX
7efMhoeZrxD387TO3NOwZhWrtdzCM4xjvWThsEDK7ocEowB+dUHqxRzdmWI/h7xE
CnrxXrh+QkTBm1M2j/9ov9JEPO4Z79+uz0EDd3RbDUuaK29yGCzI9DFVndAlcEzh
WjO4jOsfpUaGgWXhhtSCKNrfOGDd4NOEQqzpmt+GqRseSUpWEevgdKfdJq1oLUfo
5n4LoqhJMDKp3QCGMrfwIaM9KJhAdXMmRtaZowB0aN4K9twvdjbtKJjiiKyzaEx8
HQ+iloc/RqdhJ+SdMOTcFYXKlAJ/v3egAM2PYGqKei0UijCt9VM2d6tJaYvti0vr
k9tJBP1OfrZantwgEholhtD7CkuEY4q8HESk7Ntpzsw/Oz8CgmhkqbIDtT8Ar+5m
vOoYTbc+8Tm28kKFoIpp1QUrXINsYvxrZI0dWoqmvaqfeAMSPABwch/YTtmS+PmT
2HWXd/x4ImT1E1BLqBZ/ALWzWrk8ugegPbeuPlkuOLSFcV0g3408/SgWbbfLhog2
7PovsDSyOtAp0ZvQKFRSTNjUW3oF3W4OEcErP/yPo9Pwc9FbF5KvjuIHg/7hu4rg
5u0ZHcQ5GYCEnei/p16YX99LkKAUEjLNTaNrCwe9ly0dXz0ga3aDjhL82OuMlLoT
C4MjXA3sEgpUseZXiQ1O3nMZT/f52dhNPM8XxkuqFHyh8FIbbuSPxsdWqZ+NfRQB
DWrAnJnKl5RV2KwSyq6XcnG30BL0Vvi63aBWJsfcgvVTn/Qfmvv81K6BfpZ7g7wc
EFi6z29GXm2E5CYcM9fn1lQD0GfcquS+b7USdD7RvCzyl+WKCEfnMxzGzi7z71RH
kHk8NhBJE+IjQ5vJsgGWjXTMMUrqOyzKTwKY9xEXJZBtUXRfdsTumx+1DzbjTi84
j2AWIWf3eAW+eaodKeVJ0n56HfcnsZEyj94TL/vmbKMx0vPEGPWj4ou5YwKdpRli
jPlfp04K7kNW6I2gTZ01qAD47osm0gfkxCQwSjlBfdzaCAl/ejvQJRUilNZ4NWun
wp6wrQ3J9/Qa78lMYMXLv00aY4TpDqBAlPFDXJOAx9KqYJQCIojMtVlHL2Zfp/E8
V4VOzV5M9niVmvxZdaNRKa9E9CMtYTGQL/JtUaOgzeTxBgl6oL5mbMX2cQFcdPtl
jT7vOHIXbp76NuGUOyFyU2imSXgnmwFzWnHu9/zmqNYLZTP12b9lp5CmZJvctcUa
gQL1NMHgA4vCrWksxuz4UaOz0hOi0Wz0ddUkB61sDwvrNtscosyg3HFV/Nq5Q8dc
tpTAeJ9ZXTlDE1Ixw2PhsQh3DWL3I9MxrPD+nLkPoDGUDRQh9QMP+0URqK4+lGpK
iRBhlyyhDC/VhX4pJzinzyL/7C/yKU1e3owVpuuAGMW+yaiXII5Z2t+OMgvg6vKR
if+nJdfFd3sg5XDuiRDB/F2fZdCgw6QBj3JHYlXQpTFmJMqUXtTeEP0DZgeYamfv
k6wyUZnkZNGQWlv0shE5zkC7OkRFB291B+HReId7a4MUOKVa64VYe5Ls5CGbPYCZ
EOZjvDdfMESJanvbfeMbMxMlpWgB46hKV3X2rap5LZbJ2wV43jTBcmW3YCPWkj25
1LqVziNwfkADk3Z3lJLxnR3vjmWUxf9Sl4MLuPFARPwj3FJGbo1e2RAOZgZKvwHE
EaiMlLC6zrdl+jGWaSBa6TgcrAHlpMPYVXSWAJGJxs3/UV1iaWbIuACNlHZFSFSV
OQcPvK8SDnfvi3LfgkMse0O51G70/oE5c2ypc0HJaNJHjyMBSi3eF9CngXsk99i5
U6+voa5A70cCA3tzaTheoFoRPN5ubqaf9JBEM7OGMrXPfAII/pxSp88wV7Vp8w8w
sH6+c9d/Dn4zCJqKmjTbIQRn4ImYCwJyI1IO/yejsGXteyaIWX00VK+pBUNuGjO4
khWanWc8A/GDOSMo6kBezmSL9ah9LAiJgi8sw6tIfUaubb8reblYmsszrhrBwYAO
IpL3tWxW0ysSVq8bmfXjWctdpK7YuC6sY42z3IM5KJsFA+OmT5daWwrh8vJl1eEA
DSAXoLVMFNGBZvOUPzTf/gIbfbhf3gHX5NwoaHvnQ+D0XxYLnX5IbmBB17r2kdNk
vhhelXLBgJCHYZe1TnoPidh/Uvzullk5YjxBpGyb8OYdTjLYk1hta2AqdST5f+fd
zQBMPg/cmga04KhlmaqSqlJUdDkLcoe76a+xArltWnb370wCXJUufb8BYE9oyTpF
uszkxwlSgo++olFHQIlO4EPfSwnMR0j9hMcKOElVJZ8I5PUdKWNhxYzveYUZX9iK
cpnq1kYkomJzhLoLUX8cSyg2CNFIZkuc5PmidU7l2irdcCpC7PBshRS57DxVWB12
9vExDRKkaPnJwS/bt4gTxSY586+jc6wy1sz6NzsLiHaDYz8n++dKT+dHUlHvy6Oy
oVYn+6qYGcXlxcnH46oH3ZfuEtq/qJqiL0gNbmVtZdMZbw8TWG9C9LU8EPN4j5yk
NGV7ibApGzOXsBMbzlSB5vnh33pCeu2HXaxBxFKtH2LQmQHjiybZSBnVT1rUWNsj
z/56SR6UV+Iw6/CyS7QuDbYFNMZ6xbLF4vGPn3w3/tp326oOA5KRrYYy5iyJPgy0
XWFXfqb0jCJTAC4g6BCU7c3aw2oJ+vdgs+7D6k/PkfVUh1GQj5+K1jXYNTiSVhMx
T5hmZEz49ud26UPLkg7917v9N+iF1KgAkLkveHJ6NNfOuFx9pmhxyI2JkxpfqEz4
RAuXd3Q/RoWIpQblhWg68HivZXSJHB5qQtx+CgGtHIQxNSRovcj9eD5QP/wsRY6u
HPOJ6MltcQmp/WfJN+j31ccuDtdmq1n4r5VLMBuc8BXe0wU0J18TCKW7M+q7BK3r
8nVjGTR+qYG6UDMWp4YpsopDbCoiNn6dZGm1Fa4Nce5qFZuqebFPdK+mIJJiKbJE
/HPpEc0d/vEiD48UtlBJUju137F22dC+3jrVhIZBzceoqzXge9LwHcUEE7Oy3Hpm
TAxfgzQTxk5wAxkeKb/To9+Akpr4rpQODz5uG1PArwam5BeBHlc8gl+rnrmZFBfI
NJdfoSDuySSqxkEogSSH59+N366AQ0GKdcoAp/Z2e405C9xetvt4vtdZBIW8qiPW
zwo+BPvUA1X0UoYCE+5NrIN5rdWhXkeOLYXVu97PGg0QGmTvKdcV7dX0Feg8c8Ud
hC0GVfbuXRAvYYiXCX2kD25zUmMefSlTGYm0aMkriLsqXRunSzOBBeYcwBbuv0xE
8zyF5U/lp8JXBQoLU39bWOe2+/hIDVgB3NmX2PX26HLP05CodqpTyEk41q/UP/gx
0lZHzVQ01Q5MxvSkUAw8mHpCBvd8J3Po3V7TJuFiwmxG6fuA3bJbfIaPO7t8ILAT
V7/jJDT14bhjT6uRLktS0C/JRvI6Tgdf0D+KHvE0Kh+H1SYbZ+lJZZsOoc7AoeI/
SaU5XvzMcaCF/Q1hPVbPzx5+tKj6zOkxbcl0f5iwcu9VopbxoZLAWgJ0t3XjN9s0
C3Gsc1seQxmwI7qCTwKw3BG7dqUZC4kfnePmL9l6ojCrtE3ESPMD2kIR+6g1TLkY
NkEvdpyIRxmhAWf6waezjLQTfy6gFuMUIitpasDuUG6aYOjqwtgDBqGJBN/EiogB
YyQfLHbprdt6lcsurPuEe91hr44FSGCRDTcQCKSDnx7RvQMM5Qx6ZgkZJYyvDmZf
cBeuX7wTM4JbBdVe+po9nj1cXXGGv5TwoaLMBACl7K2osgmYrpUKydkI46bcG0M4
DXFL/RpRV4e4lJoSeL/xQ4rfozq/n7VQnfRN0Ib57hhDX5sNny0Q6131KJfddSOb
3PGkqm7iVeJFpklQC1tS2uLx/hqtCplbNVGIhqwipsyjbjo5knaspqlzChfXrfCv
PvspARW1pKIvoLv8wnopPIKxutVOXaqTLkdj+rPA2wN9Lg6+moeRTt5Sw4K2OXz8
lqK6dvlWMSIMVDJXFDA9VdSEpsrFeqt9Q3u78CN4AoFTh6LfUMD51bvz3jPyfQ2K
GvWQM2Q3fNZj8Q7lbrq1XIEtikvTVgxI+gry1/e2/XfS9Bwk/lEIhespjKqzDfUZ
eo1TZfQZCML3uq0smS1wozJ6pH216tfhwISEggMlTb8EktOZdnFmFBcBU07tjvzO
78nC+SN4pMUc0uGNm7XOOb/VJV1wWhVsCm+LTNReBgl0oInxGNNa20ZPDloEImw2
JKNfE1Mu+sojNn+lw/hiV+nQBu35S8ugW+W9VxPuW0riACG5xuheaheH6f4M/iBW
frAf6hzDp/Se+E9RJCoUtAI+vTXiTIvhsuvVmjcqkNcEDYCsmwGoHz1CfQ4wPCQP
mwZPh/fA2ogWmzFXRBtsmbnFm1pm3gZeg0bV3tjeNFVFU/3EsyYvttgpdYSOyzEU
QDb9pfG38XRYYKuGsX4K1FyFo/AXE/Bw0Rr0WMjNQLS6WesuD2XH1ZrWen+qX21L
Ew1I3a9eiLalczWHDKtKBslrkJVKOjDe20Jw2RLz/zPRcovVKVXULGnndNY0W7D4
Z3COuo8J/4BpcpTzYg4hYmXgGKFxN2tWM+XmMZVbHwvnyJyUndG+hy+SankbZ28y
drlOhRNdeRfB8eqWcZe4idQ8NobweWKaYWCz859Rwn0mafwbBubq7Sy5Km1G4y51
IqQT1MNc9dXawayJggul6Z8lxyYL2z/7lGV0j644D9s30kZfqFV0JUJsSfNHjfF1
5y8pgr+F66KaLM5TzM2yfl1Apz6Vzhlqnqxre3Y4xWepOnIg4YasJKYOcY+sziHt
xXemDbwO4cPws9uY/e47mpVrttjj5ChunSbK8wJ0WLrZmIz1n8vO51Xq3yXBVqqO
u0rwEIinuw9ydNNltgFMK8Ix/BgDbWPEJBSOAJTJCdFTAX2fi1/7aEIcyUfRK/2l
+03t6B+UTnncGrixVDyFOEDL7qacJKNoZLlY8fQM5+O+9x+odh8HZmY+vXJumNN5
TpMoHK0lHay8YTxd3BKqHec6O6J/m3e2w0p8Il0DNi1K7fX6206F7n10Zq2UCkBC
kTnB70X5hB/PVgZlq/oXjOExGLebiwHHVIv+WyIVa91YNWpJVtGWdhPoHYZufEO4
SNR3V23q+04fcjP/JpSJ2b0sY+lko0uxvd4JiNcUTw4SzCEh47YJL4obQGmVCs5B
5UBk5wyHBxQf8H4A9byw28jCzWUFdrCj6xHfoS4IZ8UwKwARCyl4YuwQWwtZy7Na
KcYjHkKXU6GJ0pSlgyr+4myxCQOsRW8pxHuNgh9G1fOYO4rSZzTxElK3UFrFWNfU
kJ55xIeBYhG/OC3JwYTOsbyvl9LJE8AEW5r8i07hAw43BvnHbM7Zs8nmefaiNzGN
UesGL+j4vdaqfG+5ZD/pIpVPReNHqTS2Z6iTI+kRE1ZD2PdevpGkyiv6lg9KDn1c
f+a64OSZBfzIum93wVosd0NDIMNILWqvhqrqL0+Dzpqa03Jx8ZN2gf94Ey+hMbK2
I6WWe+BOsUHakplSIpaqyDmD4Y29GBA2QG49erVU1G/Y2ilZNdRGsNRTSpQUSHth
kwNezrJRJoD0I3V3iF9V88pPszVHsu5ACk+sJG+of18w7u3BNTcxPlhcBWJnlwrU
JqgcP/+K8DTl2R27a4rUjKOz18CHcKl11jWFaoQtG2elLjeDiBYQSbXk8eVYWuWK
vkAbVzB+PIid6dmPshrjV6tbGw9iJg+CfpqjY26MFiYLZGubEuFJ64RpXkCvtNli
QkiEeyyNSO5ozC0GsZJ0vTuM8LKM9+/CL0KgsA42etwQdtFIF9MCjHx9DtdIgtN2
qxKW3ZD1nBqk+uV53Cgz4+pghK5/jRKRDohmVr2sv0N7qk+R/W8CRdzwPlu3+3H0
GHqDWkDj7pfDwon5idxj0bqi8LSommlhita9D0n6gtnRj4H7KMocLSlrOMmGbpAe
K0bqxhOQRMmJ6poNJ4IWJ2w9udZEUyB9Ib7G3tRFGbj9PtWYY6FIX1E/9cpDgOU6
yqwu2YMLqSS+PnGne0oUwIqwNUQLc/W/E2j/kVx0MMnyXg1288/DxMElXt2QV3S6
VbPyQfgiE2WTfWjFcTqKfp4rWrie6bIjSm9OeZ8ZLkwuoO2UzW6kuBs6S+D73gu8
Cmojuf9p0ODwUikg8W5rVN2Zu9cYwo0XUsDtExZDJvSYzFHkLt3Ss3YhcgHMyCte
Eq/efK92vZPX1DChHrQUZ+EDkpSNM7VgrB64u2zeI7Tri4R8I8qV8OkrkNNNg9FD
Y6hho93xdO9diZSwX2BN/Qpqpqcb4tS4nANLGmR9TslSEEJtjSDxE075jMSkGS4f
g0OlgYkGfXHz6gpDp4AOJY+StXZFhFqi4qsbH1hMY3tjaciH0zeCzKXx8CGkuMLc
skTdcUpxppi3AdARb3jL/sDC2TzAToHymDmaQuV97lQwYssiFJ+6yjRHSux+DlxI
qk4jEMKNRKaJv0Vfq3BQHBoXc8Rw5JQdtZONvM1nWNCtimQR5H0iobzxh8TXZu6A
fxLEg9NKGtDA9Xuvj4+bNf7omEOAOSOGzDB3WMDrqOyKxq1yf83LBfszl9Q/d08O
fDI72cqoQzS0h1cRgfUw847MwQ0bFIzusHNsX4Rrfm7vWSTKcELMKPZrL6fue7WL
+8p1UZ9kuxP5dYx4+Tqbm4tyYx3sFYCqejILnxb5AmifHT44SPWT4E/8k5hUyWpM
d4nj0FmUJpfRDkW2IMYGhf84jlV/zOAOECnuQbErsNBarCKiwUP2tanQySIQv+OX
jZsZ6slambvrLnyHe6m9NMpnHlicpW1R9wlRIszZ+vTtNTF/QW/HAR/WSJ5NwR0Y
THzkS3D5WmG8INtxymDsnT+Jb3Ru6hBG0USH2aHkpRAX52UHRZug18Gd4qzehAWr
lkKd4S2LBpDnnJlxjYxQWZKy6SiDMp6yJmixGS8prPMKvmaouZh8nL3//Gqg2nyE
CM0um8hkn2N+OTiptxJJiI2kV8Iv5Vy4z7jKP/NeyexSXGO2IKePpjts98/xEXT7
Xpwig8iHqjvPWDuAD+PBYvWRFgMgI470uV7Eq1cM9TuWjXGhy0U/l0BcSrMVMtEE
4anaL7ziHW3kEUjuR2qln6Ykq1UmNGH0i8ucA9FOyR/iHcdKD6U9g2awfRANGGPe
TgoCPcH6zdVXSc/7qhypCvgmoSfrJlFEn0tKqM+3XEXQocnbpyxCBIL9efzprNFh
aMcDjkq4o3Z8bAjFsmR/A63PeNrdkpqq6Gb+9FEk6h9/gC8q9OcE9yTUUZfm4AS/
gya8O+cuXvlZcySrnr/7SWbWJLLZNmLDAxZxZMI3jOo5/pXgaDeSrzevHzHHA3uF
iPwf9i7Cjl9tNNcPFN2TioxTUK4y4W+ft3s1AMNuZ69eE5+yEbaMhMcCa4Q9lpOP
S0PiMLdOAou9lWS85GkIoLTUmijpqmKNWj8q6FGS/ooD/Q9beuf3xriqwF4lh6+/
dKMoiH9fGls9E/rX5S/DWuzyCWwkC2LNpXMGX1FOppZhskSqTLC8AWXzkFAzOu/O
fG340G0S77+2VpqKcw8QZkNvDARii/yqhemWUaMddd3OALmWr/DyEUZhh566L8Eb
986gut4ilCwAK52jCT8VytzSHWp+7Hwz6a4jgVY+aXtb2GMJE4bM3IMaUFbHinDe
V9PgD4oj1v6M0EP4akKRsCIP0ZEqJJSlc+Jyf8D3YkD0n/k/wemZMAF2ITeGAEE7
KUsUUuY71gO/T7Y5brHjx59hlf/rAOZtzZHy3c3pTyMvfhrpYFniXiE2VhRlb6Od
V2pvqvS+xSEOA5Mb85GWSN3Obm9C/gX5HkvuDlzh5NGXGuqaCybmh6cDr7T5H/Xg
UOihchWh0QHLGb5Tq+8XRqBRUegjtalkNyU/WkMJdjXbVf2vrpRAAbOMlFSv9gtA
N+pzqSUaNekqglAx7JcV6kO9dXLrbUb6h+ePaVbCgu/c99psZgLs9zjXVRWAqfS3
WM+Bi8RKEqqHyXxuimeoJuuUoCIyjTx/dZ+/dWgDI4nk4LOAkAqMLywQNdLYLtvR
VduXjI2bH+ukYLXLPoSfv0ACWP+Py52gpuo27DTN+vWIGk1XWhxAooq/JfA0DfWY
MXTsRd+C0lcifX582FVJOlbQJPb/CI9YO81022uXguZ052QocvGPUJsnbJagARNx
8Heq0x5DnLGCotLO15H6Q3ktVmdANr2BqmlNlRI2mueK5y5AJkOMFpMyfGHenqjF
3AJht55jN76CC1jplJBvJJVPuXODdbAqRHhIBeMLziWUPfSvI0I0jMlLeZB3/Rqu
fNNySlYYvvXTksc4xjDLUtBfHL5QgmsC/5iQbYpDDpxSjVMBrVY78r3c5riGnzUG
ilfuUvB559aLYiRC5S2qiU0o2bAKq6vAA517fSiXWEoydfmr37w7pQMMO8coowQY
I8l+CfTfQjhebzZjROhDByPiA26Szr5vV+9Ak+OEHa0QK3gf9g0qyT1tNPiRrmRk
Z1vjSbzcGMBe+lkDIgYlmlvxoKkqa2/lyCV/Se+O5H09qSsQnWoTtJUArH4lVu2q
bbRYLEe4OCLHeDKiPHChb6xNwe0r84nmXGjgjkF5kg6ZwC5HrFfrkN3AQRgEg5TR
dgYrP0WvNF5G45QThBDHKsbNYaDTFO1M1bEbl+VwBjmWU5+uGe7P+n10JMGXLXw/
jTOdZ2Q6XgNJqZyztCxHwxX5NAsch8pWhfTeqUcRz6W0DjSMb7Guc7AmvjVqLQT0
rkqxR6K/AxC8Cj8PvwBbr5FmvtQCV/MraGQSLdJZmwbKLXm9Mg9LglSEMPsh3/J1
YQLiN+phAzUj/HeSXztE8HqDP3BpD7XubBZlwJrFAiITLTPgkFliBP+mCJ6mzeB8
vK8jkWriNNBUtU60kGtatLeYnmkQDgTg3zeGzYuBY1QlScoyRr0y7th0Wy81DF0c
w2f3clo26vrz7cLYmziW4cFYHDwqVWk7u7m1DIGijXEhWyU8tckThY93mW0IeLjZ
0XfvnHY2JF7Xaijyo65DS2JKLh1tlyucWuqfxMltO2SNg87+HVdypjpXMgYt5mB7
WBZeU2vtOtFh4ztEOm5TjzMCLENsnXtr6AtGnEoqApQEYTBZ0H4dCay2xzH9Mocr
Qnfgie2Pth5pHhe9kW5rmvOgJH3+AGnbPlYcGInT2BtPSP+vphpvLJ3glWV5SG3l
+iBwqjT8B4ARJNiJR6gDwM17tphxq+ZvKsjDyXYlBLwA9JvEqiBRSX0g9F1prtbK
rBc4ZngFis7XLHcelmT5qYhOoFrfXFSMYjUhuJ9PwfDW1MhP8jtVArJC0c0vTJ/G
sQIXcEtdvn0zWC0VSgrspKmXIQ6f+c6Ph7Qb6M/rM6VpFPYF/qRFxOzF2iax02Cq
InIJwP/XcOzjtd//S1rtJSH9K9zg0m4r5CubIkbwL1rY4+MxvTseqj6eQSQaFou/
MOHpOhpAtdJxIps7/IvjVejixmsCxXZ0TTRMPaOSu/VimpUfJvZ7SSbhvrWkp8lw
lpOF1M+0Ie6I/5B8i3ElGRxU0YRefVwNDCZbkcnBXf3oFpa1xDI8EA3OIrfUclF+
YqE0RC6k9xvu4Vh4S9VLO1XJ39YWNMSJvwX6k5ToaMPUmMkK2lehPdjqqXQZANtP
UayiiIJpl+GTtpz+o10l18534/DYvSXjQz65QjTEZUpL+ld4IIBrfZRHIBb3bI6P
63/zim2C01WmCWVLa5IgDvBHaPKCgsxlN6lSN36l/bCUXHtxOm8TyS0BNxQX7W2+
IFr4Y+HBnvi3Qkuz1+Xg+BS0tLAY2YLnaSzdQ5ObkE3tfCe74GCSJaMnThhBR7g1
97mj5FafMFMurTJUtngC6w1wIKGc75x8pRyIM/CUAeVMS52fq23JOP9B2FGgcxAC
K9j0S9yNC6Th8qvtklOqKmggF61ivKkGN4Ah9HhVXs7Xtu8vfYs2xxXsB1I728Q1
wpG60YNSjEj3SOXH0KUqH0rKsY+LIcUAcaWL54ok+AE4j79fGaowV2Seym2kjGTx
bI8r8cbpmMtrfDROddYB29Kq6Bh7SwHZHzo2NMOQDrrorgRg4amCB0lZ1KJSx9Fs
8MCTzgTrQkvbx0hDZFIuXmxnRo0eDw9eK7gokpKzVehwOxPX4TMT+amYFuZxXqjY
k1HeAxmNbbvhSeONuN07IdrPrpxKaCZBKw+OHpjmMfghuxQFPti/A9kfrmgbzyEJ
WcAR0ei8xQPrEfqEoJdBZSqPvXVJWfN3LWf+TWjrBp5OQ0wlVqbGzEW+ukw66yg6
vhnnk74nQ33bhTrCfoE8/QN041qOsh5/ngx+lqEjaeBmYjwdboOFMxNmsADMvHdQ
R7Rfma3C2QiRYWkiH06l82XmL3KLuNZ2cM4/zXmFmFl+SwYYxUDYn8nLkhMj0sLo
hRzb+4iXcEiWflTjNQIVTao0m9hZl4xoP43bdfJIBWDO0K41Wn8tp3j648OIyjib
aK0BoDHHMGaju7CjK2K0A34Jpb4CYPmi4aAy6Vr0/FednyHTk9nY1C9Nt542nDwG
Re9gvuAGF4kqTzYHmSG6wR6gylsuqBFwap1sr5MsTq6Tdj3k5uxG1/C2ahvO0MJY
Oq8GFJbZniSQvbo71O6F9rSAQJu15c/6DbzvOA2NgUiN3Q35jrKfCB6TbXR65XrN
3hfBICMvULGEJc6/jqNGs6YaLy1akj7WEmadp/3rkluUDNNBVwrgU7gaSUKht4Q1
SDhb83JCUHPx6AU9Q3XT3lb5ZBCegye/S5ucygfwXL8XbJgmZSZH8GeTsVsY7nxG
erJWwcYajEnw4ITV9ux5ZH6k9OdNVDIts0xgpau2F9DQlcD56pff+oTlIRm7hfpY
/De429m3d8QMD/3LZy/n9BVmhPNh6z6eHfRO2QfuIsubESBBr4/gdJGs5Y/O3cov
fEngksiEvQ4HzRj2NuSNz/M+OyaMOwWrL/hb7CZ38oH+9FXewmUzTT2LxU78nZgl
aK1pv8mk5XIizgKJO0DMA1LvnD1xWQRh3Cv7OVw/qCDxiRZbXFjfCa1jv5g8afai
Ynhce8vhCZKdBkRVBfiNWVGPH9DuJsTTrsmT0OdvrZzhub0SXpcC7egqr/j8Tn7y
H9G+DK7F/KrO7RNFMA0cFXcqrsOYqi6BL/HzIw+u/Z614BoCJcGB+8AhvNpRoFcm
HCub+QpG0qQvA7GM2p9vfDqvujVcZ+OtnM9wzQl7hii9UdI3hYRNL0i67BQR0oQF
jrxhlxzKA634g9ubhJMtuIk21hBEqwZOAD2e3MJUduL1QXaWTZby4JcdSivT+M4D
Xaf5Ob/pA55BcwZTWjosHWPReN8MP+PUVH3TPkPaSpoqq3PC4pSkVXjYfoGUZO+a
EUpfwElgmYozCAgZZ+t+NYIZ1I7hyu6kCpEcsu+pjHlEyubJIDRrlSdnhytxn6Ze
MttvEwlXC3tJplgpPmty3aX5kpJu849+2HMcjutnJ200xiLLod1ny3i3J5Gpa0jD
EvfD78lgxjquda/BnA1e0ZO9EByTkO7bUbI3Pwj0VQiVTj/oAB2z0N3Z9d4P5rBA
oxXfVyjuo7DKsy5FXyx5oibhpbzr8fXfwpAQIAqPPe5afx/00w3wCA0L/uzB4BM0
Zn3GMzpSb86gfqdbe9U51WqrgM6WO383lg8NDiTAX4o17Dw2NsURSKUFB6XN5WNV
qnYQYnzLL//bm0hz125WhSbQXpGt+BQmlPTj9Q+dLUmOzSQy6fwM4abJdP2xuahw
jPQx9EWUr3eXoGEe3sxFyfijBxnBAppO4tPVpFvcequB8t8q4PykV/5wRh3waqCO
Zdq4bPinzYAVvy05jb8kp/y4qQsHQLgP566ypz+ZiJJgI2hGGxZw3Pze73NLxjae
IYbvHxalql/yAfEqzYxvL/e1ry5mGxnl4v0YZj5gTi5nDk6+QvhaNvlxou0cS501
Z1DcMAuu6mvg2r7VcUP7+DCADlmPqfGyLkpxjztzbDqqKbKJVsl5HK/D8AOIM3fl
fraT4krnqEtjJJdhEEqWmB1XVUeXVSVSI73UN0qvOykLVrpsZIFLLJltFQ7HJTvb
CyjLn5B9lq9o6nbKNMLaWnvMu3XvKQ+ldEkVPil9YN9pwFiD61YqDY2kMVm+4ZI+
u9bcYUAsDymsZAfeUJl6/fwElVC559gEs6H6GBoHz4gRfZKnpCK0Kc8oZMvLdSxy
Rl7/PlRXUoPvutbI1d5IJf5aEzIk4QxACpfkhv+gTHu9vGEKQk8SOBz4MlnQfRxX
VF3/Al317cHXlrhPlBjIu3l6aAm8OXLOd2cNRDdwVFdexc/9v98lV+z8yqAzoZ7C
Qhntg/zOpTdnLT9GPm2qVQ/vc9j+QvE8zQ4mt7e9WfcMub9O6RiVhBM0/eqaE+JU
arrDcwwsVTaxXJCYXXdzIu4XsZfTwWeVcUdOxGO5Zspw/aOsQDTeJ5x2reVmlPUF
kks+tmDDPb1lqAbbpfLS5GlzPI2XU7b97kjaTpUaljtTsl2llGb8AYGndUIhxnkM
xfiGu8j5oj03ykFTG5pRCh92K5O8KodBOmH+qXHsESPuJ24xxppG51qqwoE2oj6F
B2rhbz1yytAD3oxmUNO9YnfzfLtptfQOEA0Lwd0DDOorqZW8rJyyFd3GiRApioWy
2rdrROQSSoH3/He3bpc8PEJRJzoLd3rLvP4mXFq7xcEz80jo9FuqK5FKD02JKIyF
+aazXe0+5t+lAPPIwD4v7MF+3r93oaVQnO25vPfz6Pi6cbDCDwhTdyEmJmVS9IRl
GGTsz35SvdS9lyFp0bLaL1GaHrlBcFRFjBC/7oAIN50xYK7eqXMQdCk0KY0K9bg5
3E264WXNyZqBHEJWqYfpzrMc/LcBJs64bjcJ4mNIippWip6exFIFn9XfIThmI+Zx
qhrLDeHQ8A4whaaUStEaZR/+1VQR2c2yZWE71EdmQrh2/5340Gr0hcPofJ+zxVH2
mL6q748nvRUragAyCZ8sEgjkFlLK4DT1/TuI62rj8i7YsOp5l1xWIvfYLGd9Jnxf
jlrkg3Ty5bkd7SWty94wYD0wq2HiXWAErVzeKbORCqhYjL/ACvAAPGlRNzz5sH0U
kabjHiN+OiR4n4Ep7kJT6I1jOxXlhn6IxecPW4QgbukOcygx3UGe9e3Ls0n8b3xg
V61vzBT9rbytwHfZneQNuxFvvmKFTF3ZU1EWdIgb6rdQhEPxHm9+PDsyAqd0dGEg
PiRPARwZaWE1lyXzzOn2Zlm99W4mk8VaGlZlhfe0E8UdXxhuASW4Uut8V6lZyqBn
KfffWcTrV8Pa6OnPoIcJnyBZb4nSsGbZDZ0ydqCcGtmW7NaM26NLEjldksE940Qi
wq+9z/bUfN6rDc0yJI3a8fMFHaX8oRJ+xbjlg1S4wRFz9+sLFwRFxxyclRyy1oCt
2KI4qZlUk6trY5tTpiCoIxU+U0ihZDCkFSS4a5HUZF1SjpQxJGFLweTEN+TJSB8s
uThr8LvB3++MSQUvfRwmTe8I8S8K1TdB6if1BtBBUno0PMJCShtW2T4GWHSbalxE
d5SwhyPJG+YU9IV/kFevfPtM5Z+uluhhsyeZESgQ9jPeauz+4/ffxbe05sx1k1/g
oIsYbMX2+n8Bll8RWqLST2y0ztry13Lhl4R1mutbcJfODXLxEgUbkEk0Hs2E3cJk
euLU1E3g7tw01/5Z+5e0NdQTewWLY9ekS5hSbvH9nOfkgKFqh9GCAGnJR2mexZ4j
axQX90L6D1Cy1Nqadj6IGBZ8DksXg6MhwZYrIAciiBqB7eO9RHo9p943Bo7KRO6J
k+PjajZnXt3BosV0kZMV5NE21qsv0bb/L98JVSIc3hRTEMTNv8L4ULtmvREjjOhe
tZ7W7p7oOIuz4N6PrCEOnZX6oWxffs0MLFKXNniTevmtM9nFscuW+Aah1q7mkZzZ
rQZlM9P98Rx9SBtMfT/Hka2UmVl60FhVTH5HGqGD9zdNyhcB4TtDZAes7lrLAioV
H7DKpwQFSv7ztz2PM/nkBbw04aE5dPHRA9kNqZLypH5ZroT9m1u8zP4svQV5ACPv
95O7iSR97Cl8UFZiPz70CDaZFKEhZUM1wUH533/AwHRDM0Le/spNzGkwOwF0f0sU
VTQYeMeE2j9/vzMsTj5HhVBd94qiqWmh78w7XEToI/KJOceD2vt/2ZkclD7aTO6u
RBDFJoBlOj5B39rgdTanpQsV5YACF6k6vgs7zMrX2lnSSpoTJn0AYhMNGmNqRq5e
RPH52zXE31QY9xcX9YxjVJWTn000LOKEYxyK6dZsSNa9qSAWXfwLW89tld9gu1g7
+DgQhjLRQJcIfQtdHBTqEfZQepA8jK9XQOb5bEsTP34DXbqzlBlP6QzWa+7ca9Yf
sGtLVF0H9VoRKz+NJfeFIZKyfvEZzyiz4Cou1m7SxiDyB8xmGegsOhi2P9I8dnb7
vChUGprOd+w5Lue04aXIbobiej3zMmcLJDS32tfQuzEfjvJau0bSYjjHXlH1Mbyl
E84lBtmWvCkunyRfbHY9SVe5AF2qq+abKlOHBBr0+7zjmigh7NloEZ3sL8UMceyl
I8RMtnOQzhoq5rzq+EvWr2IfPKqiewTs+kgCGIm9XQlB0YE3jKrFFcdzCjTLAfY0
h0LR99kROGKleubEK3KXCq9LGc48K+KpK/rFOqMfIhLRPIFhkUt8y+Oh1pfGBPS+
1qboV8NEZBymPwM1VTOEWvu9heWRTGhfwy/F7lBwI4kggBeVKYmGLrnfNlV3HhDf
z8Gthg6n3W8JOscS8xtbphHqLoHnTQQnzrOBdD4hxmeidrYMkwyPwPHhEFcQ70Mw
oyDII3TjiSxO29K4eBCAviR9NEcLh/XatqWvsdmmmWJnmYU8fKkoYYufFqIcXUdj
ybp6DBnJDfF8RM6DysD9rQLlDMH5bnocPAMMC8/zyC1dgmcfN5ewDpIddCcdJvIT
XyhZ3Q7c8ZkBJxGmo6U8pM9sDF/Q6FjNiEXqSwtwgWjNdUDC1tGoevVoMXdT+JPh
ZtMMoAYbv3l+wc2IRy0bSQhi5WYM3Zjys5YdXrd/RgHjgFYFm7mkXjJ2UxgOVK8z
I7180oHjNI5YKL3sEIM0j3ZegY8513SFNSvht4yLvpzzARfsNsoN0F8ECIEsT35T
bkpk69SSng6WR480TxaP43pnaaGxMYg/pQWyOdcubnXcKeP7nfqQSVIpuZDPjxxq
dfooLB5vXXHjmleXmmJRoaPdHL+iCWcC84AjMfoNG1v3T2e5aHcubw1tzl3dWqPD
RImdNxjH7iL3dtNtCq8M4OTj4vUYY7eOg6Xp1fYRKNWUluHJN3cuo0gwNcD7h8AX
pJ8tIebsWpugl2hfy4euvdjcPhRiCtr0E5r/fuelJSEXPpOW7el7acDOnR+AObdH
l/RRNzBrRbSMeheh6d90lF1FYh05Ev+c6iblCDQ9ykxxyF9mYK74JSxLTbC3R/hX
WyZh87kwb1qr2QJTMRwRhbs7eget6ZT2xqI6OShL4yR2a2FDD8cYAfOXpH8sqwdP
7c3fknoQ3x6UcSps6yBlwyErzFWi6bq6atZ/IPFVZK7ctoeWz2c4ioPsrEfZ6KGQ
Nm4niDmPn7a6y61RKyu3dKnmf1fT8RlZHCSkisqhlOqkFGSKOdEPuaK9bkVPIlHt
cnOQNGzpQSlS6Z6biK1nIFQ3rra0djfQVM/cnPHg2VY35eIA3LSqzxqyk6y13p2Z
dfCDIDdGx1JiBHimPdj5Ae2WzwmMkHuQ/JSRTrusjK3EzmfwL69b91bPyAlylMwe
JPTH8bPViuv4a2NsXkKGOM9l664Rasg+anbeTVjyAiTF+ib5A3EZlVBSu0CXAW2r
uoXO8VcwiCLGo2eWsJhzqoBppcE0p1R8IyrBrmUFgzmrf36yb5F1ducWEqRW0knI
GHLy/K+2ZMcuj2KlR5Ax5hwgpTVa+n91l1IXkoOH5cc+GhSx8tnfH6LdZbt6EOeP
ouTTat6WJnwWTe1Z+R3WWtmcjcbmWHLF9xs3MJMk4bYUC20wJ1x6KH2mscaJPz/M
ZmkdwkaFVOMPE/X+d+WaAE9SeCf+rrCYJp9kpmQsfmFUuAVkV9vCWL3SBcHGAoSO
WDT0nHbIICK+AkxCceEF8wqcWbE3hx7Sc0eHhavkgoRXx1nusSxd5MxCfvn+ZhQL
Mcl+aL+uEL2R/VigXKh6WLbL9oLAF5GD+E+x+wgoqGNskfkYqbIrMvDx4GnHUhsW
Kdubrnoi1wx17yuKF0gRjvgvenW/KnWtzurhdv4IWUiz7UAZ4t4cIiKC+fMWaCIk
6oSccUtLjeENH+m8ue+cmxml4/cR7KqW8pCRNyA7JUhSKFhSlmcwvhLtqFgo6RgA
El8q9NfXp+Ni39y2+hJ7B6KZc6o61NZx5u7azuKoYrrUBYaa31A/UaxqPbYvcm6m
2WKWQjKym51pW9aoLZYOKBE8MlKS5tjBN9r4XCInTSdhNxMqB1b8NXOFN0TT8npP
fuVFo7yvCHFBLSah7oWJ3nWglqF/HhM6jduX7WP6W7Cm4BtyQPofdZX7NgBJE4Zp
AxlqDGoavdXJPzSnJs722iyQRWLiC2gQOQAh7dw0LSSRo6PasqpAZu9AUOBS8DPE
qEI9ufWJoYbcA4/OvIH0W4L/p2Mj+6TfwU3vhrf04H2eEzQwG12aVNDTXQkS9uzT
uls8grYvoWOe33Ux40mHxuv9omFW9f8ItFGSWqyjV/rxLR69urinje/x6jHw9wQJ
mYTZJubTIx0Es8VgJtursrVy1CqmzoVoRP9RllaR5/bj13DAAcsoZCDyH4GNp19e
hyAVdoreeXMkhcsG5bn0IsASXRTQp/8zfp0AQRp8apxBHgAN/jGOrGKpgK9//fPg
T2KWRvvNtnx04zOfkOibIMrjltvU+m5spky1hDX6XhVGvJDPGymaaixGWPajNFNH
us1hO2iOo3SdGMwGYO6L721IyIo8mgWKeiKMX3dqskPxA06T9KkBb5A+Ztnv7Yop
3IZLVRIninj19Vr8h+dr+GHKk4BtwncDXVd80IFAnvG6LsxAKK3/H8EDE/TypMjl
TsVj4aD4YgSNBMmSN/VoDy7i+B/9m7QQ6ZKynB3Wk5gxpEpQq9IKLXajGR3U1ImW
ck4Q56DNvbs1l0TaKlYBQMHaxKfK0F6D01l+fzXhKXHIvyjU3SbrSk3bettDqA+B
UW0Y1EVSkXOuCBNOHi3kKDLkhDjOzDeBKzNlvHTJ5WhuFmSi29B1WxH2wc/zWfqN
hcYWLeBxqvap2L8DngXImLTeGxx2Xt1V9Zd7fGmHBG2+n/36gBdLcGzSle3KKlsn
uDoZDNl4sek9PpwoquBPHXq3Q/JGwZLSAeAKbFCq+89BJzNDC6MxNxA/m9wsws44
WQt3m5qT1hvStwp1BbWzLKu731IXhLzo9sJGHzWefbeWuTnlOo3om1/C3zqbofUb
1meAbUoyap11XmG2S2zCguJ/IhLJNaT+vacMBI3LIdbnc6EV9Uz1HEK36hAVhY00
54DHtaxR5yEsqWAcQ32lKstb8M5SM9FkavjVvW2wu1PP6gDLhkkCGPT84LQIX2TF
BL31X/DAlZE0CCqPwfjQYRkLvcy/4ye5Wf28pRozpQ+28lqT9g2OrqaZ5OchkW3M
YBbOHCHUb2ys1j98VrmCE1tCYF7HFGt1+W+5DTMQba+DPhpkUfBp47BGCPtZp9/n
Fm61inwOASr+/4pXlYrJAIjTcwr4uDz4KlPAJkhagOflMqc8ldr+9lwCaeVEdmoU
yKUfI5SSQWrpimgVC1T+AjP79S6uN26uJtfn96zirWU836Ofmy8Uo5EXiCh8dbKa
mJrLl/YfrS5/kRUgEKDu1Mvm1wL6eW31QiZm4vZJdhqHK+gKC9VKEgoILZbf9xQ/
WO9SLLEk1h4JJcL+zkiI+G65629cuuKkF2LPYPWXRZKBJaM9PeD33ZbXS0KRDSVm
LW46TRF/gr+w49cUDZR+APbS+QqDHjURHI8Ph9EgcIWRhxBrOP3jAM4q5Bqs6Sy0
tCFOTln0kQqvIJOGaiKJxF/vKRJrlQG0uel5RJr7uJBNAHpGDi5MulDqNOv4g/vO
emoclydoEIc7LgKRxYPFqfFIBfCj6VE0NWQy+L7xRSAbqJmI07WMvCL3r5ttMVZE
NzHOC58mR2hkZCb6mw5Y3tjCMTNZUnhCJy1Kg6sMF2apNpw9oTdwmVBXq53aenJX
qhh9L7HsX1touaY8vF7N+2iPNNJQluXi6qJ3fl/c/5NdAaZGogchp/z3xnH64hNO
9nGdkQowwra1y7w2SPAmsOsQ2kyTfxrZO07+h77IL8tlK24TzfCelOvO/UcGdzi+
OWST8inBDreuVMOmVhwQ+zcwBfJXVQea0/X5wtwnCiR1TyIn4DY0PvL/UERDZPJ7
VyTN7YFNQXU7t3I05X/iBtorLBbgy8iC+xaSs7sQTeun2Qq8tOFBwq7Lsc1gGP+M
Hyblb+d9AJTsg/bEPu2kA4bF36/PWoFFZPIm8Pat2ztr0906BdgirYdAj+pj02ix
PKAdE3r4oK7CMc0shxN0Xlpe+tENPkYEMruR63l8US5q5cA3zUgUIfL2HmLiXNYn
vBSoHzAAh/e35dIfiTU4ykp9AWpFvhhhWvAGPDtPPP+D+mLVlgfT3lqIY2yK088e
uqkNJz7RSmgMLiCHO6fsc3h3dqn4UYNR9phwhVZNZpCsC81BI7XLX3MuIquwdV3l
/77OrGxg1XfcJ7OPOuV99pYiXfN+yyl1zTe3HwFTHOTH3Q9D6jpEVGUc3zNu7Xu6
mFM/byweMAT40nszI/054HjYa/6jAocj8EjvKRg8XxAm9l+QgPchxnUDrauMYCdp
zkH8D4UYiiUxr8sOcuQaplJs6bigOEavs5Pn1AFXyfkAzf5xhK8gxS89pHRoHyZ2
OKxYgSRENjtafHtfPyEkzfCSYOqFYoWul1IGg5H78+kZ7oSB3XlmjyioCu7eIDje
fZl/2yOT0eK+SjowFhzjCFCG8of9TH8sGcMLKqoTFMiXHJ135fSjigzx7+bFlrbV
VJIGFQopElxjukgyS5RXJTE4/L/soQ3EDJXog+uR+OS97R2zTHaFJ6AJ9mywT/3I
r+DZtyjAVDGoeRv1pBzWXWyUom9Zfje2ovimeZHd3R08yFgY84oxlVmZVkROc5bb
2PNCQauOMCCPChCzA/dfKd+AhMsTUiHEsYIOTbMcliV57GacFeieYyifetI2i9iw
pnWrvTUPRqscjMyyxyEMkeVlJFMhNV9MDL9MAAGANe0L8Ns0MhkFk0rEk4rchY02
gtDmRkOa3BDbMEd2Q6oY0g4RaOKxaxXPL8VJ9rwLJt6Jsfvs41df+6X5k4zjI1QG
lyN4nFxXCoLIsqzorVO4HYKYdGNVZk1ZUnYPTj12B6cRykjHXFFeLUc1CQ86DCGG
xpqxAhUacupzo9FgxL8XB2agT91CjQKUxoGO8xF8h6nbb9wckrJmks0cTW8fEPTn
+DHdCkr2UZb+r0x9ap+NFD5khS8gURrZJAS4lBvJOwBHjibOfnawNGPvS9LgCeK2
/XgHw+Q2XgU+wfWOOJpIekYVMO+TEVmpCERwwt6ynX8xkr2/AYBpv+1YQMRR2QI0
RNfgTeKk+Aj55tmrumnVxsZP5Xl8L47yFm5WpjJ6s5VB7rmY9AJYcAdHn/uAqkGU
TOXKXDrx7QNj7uraeVrJNVkIFPPdGCgGkCcceBZH/7cNhEANwvDucsPLar1Qrn2H
5a8jPnehMiDeVN5DMy4dwoWNlQxCUwO1/g26gxEBijlMc9FCnQmRosJurA7hsgkG
2PWzkCiLCpuvT9J85rgeCFrIgDMbZVRTL2jJ0mUb8WyKcaGYWZ44QK5oHjnb9LIr
exXUBRkhnjLqJ8HXY8df/PYPEFhfV2283glWO4o1pWk0wihjW/50BZGk+rM1kzfe
K/VWGb6mJ6NBKg8yk6NU48D8AbdT87oyvqf+s4BMJJ9mts1sgcgT5mXHqBttKlOU
64wDviibybJdHCE+TLhnM4vxQmwBPxe4pOZrbGEi8O9hd/OrpkeVmXO6qVe2EMQp
LpzVy8DrRadPftSzxHG8TYfE3vJKyvr/9nCCrIu94B7tyxWCF6yGsSr409dcLb7l
TCYZ7skRklbacwXnYrA59rtrEGNgPyzL+MjJYss8CGvyVBlqRSTgs2nQNwg94nBM
spjUgplqgak/GZpBXTYo1ddNhQ8HrlRBIHzkW1TLhmUwzTBdKiGz/n/hQ8kt9TGm
qKFwHr+fq3ciLol2DqROynXVoQypwKAOw69zpywmigo4LJ87vDBlnXa/+m00NMId
ypaqaJrluFG1o5UWtEWbCvKAbVVYmk+7bm13C5Ow7c/OEiYMdxfSacNJAUikUb0U
xvRLFoovjSnNq705EgQAKFVzmPlAZLOZX6wTtArkfbCbpzm9PgxH+CjnnHgkitni
xSgd+mI1lfqUzzm9czQAIsFV+syFpJXoQD6zNZiJNJ9XwIkxqXPVN5BkRZL9z2sy
sSRq3ffRy3rfsaDRi2YBluj31JrSka4ja/lBGx2JDX1xA468jCc91TJtxBl4Tl+1
MiK2wvaqs+22f8w65IJ2c3aluLmCEPjjmZgo/99UiBa0+ZwXADR1pKQds0ox0czB
jvXuGCaAZOszf76fSR78ZXYT+sjESyCv3SDDshAnfgHers2TO5XZKHXWP+RYlwFw
wbLpZ3z2+TRStm5ncNENgdStkUNCQA4HdcCehrdACTRW09A+slEUXkWt22xk/Df/
T7kg173x92Yw11KxKfQJ+qXcNupPp55YPdij5/BieOBosrnUihg21WGD/fdsDDsO
XSWSyhbalQoZrPQJYnuK8nnplGDKaob2eG6bHpy53y/X7qh9D9+mdJkE7QL7OKtW
kEFm8WoxAY4W9xwRgVnJXrfvYKIf/WnIplGxTC/jyMThn81yCNiiknWBu9CnPFqW
PIeJV+FR9Bh3PB2uga2tb9DADmL1sZu3mkJVYkyWzBXXmO3yT3YRfbvoZ2kp05rJ
5hdN5M8E2PXUqZP+Jh36od97pReaZkA6j7lcUCDVsMU9NbTgTELPZbjUu/PXuf2r
73PPuiKsM+IpnhxUj5uz0KFKebIWZh3DlS6TBuaVs3R8jQEXRi1Q/24/vGe/hUHo
QqzhADoNZrDh0UCn1x5TiqnOqFuRitF4Q1ujg6hgTRweEJYsI2SZbAvshCY2E6Lz
ECU4tM+IBJ7tdLkkupPcdsSCQIfQNsJ0UcOHNDnLpgLXuOZN3uyXWxAeWn0tgDfb
D4Qsb+EOxW4CqKVLY+4GD4kzK2Cvlx3MjHQtB68HeF0q6Y8gfCQGCul+m7EllAAe
SQNQzJ9hKxUlnU6X7Ska9VB6vFui+yHPfvnjFs5xzdkYvzvsqkjxRj5+OkwR7P6p
EA8RyQXq+2mLh/Wu8hU5R6EYgNm7xpT/33plbEtxO/6qYJTu155sw6xrdeluQhFs
JaIZw06F5+1TH80fFW2V5/PDzkbrRgISnmmj0u6sbhCv8X1aThNkFhdBltBiMu1h
SavnyN+cntiv2Nl09AH11e1s7/hTuKUbxkjvW6qwlyzxBl94DVJ0EaPqZB+9TASR
mA/qxIAa6rleFnDwJTX2+7ZOU35Tdwb4opPNGPggcdtIOgH3FRGovsP2Zyp8/ACq
TyPmTVyKg2DDBqwn2+k8jZYFJyQ9E99W2fNNSEXqX4G9c3+kuWuQtPJZUfJ+7nXJ
Xoxpp3WHoVQ4bhUdDq8PnXzFvwJ2a0Ma7VfuV0aRJP7u3QjDeX6jMjEDlLxktEdt
zA6nnLl2IWbrp54IGWS33EZ8WUwMPVv3rAi2Wi6h+d+B900kKnjNRxZNg4nHvrrf
b/BG83rhwKXLivsYlp/icgwY823Pgkcg4pEejKcsWG3nTX+sVzvI78T0jSXlw/Kq
TnB/0OFzrlflqttAAGx49Zqc7I4FnSDdWeawCjA0XHEBiOA3/4p9d3JIdOBaiemn
RJEP9Ae1oVUh6siSBE2GM9pTCtU1ClchqG5obmjKB7x07U/Cl2ilQkRZHy7TeU/X
5WAV1nNmR5CsnVBo4RDB458gTouGVK8FjF9kyFleBxH4TTtRlS3etcvAtn74NQ+F
IBVnzXD+uosMaEcH5EhTV2K8O8nQ8A05ppFsf0AWmkIUfpST9K+qjQ4LtKb/A3Ur
KqcJPpHKBH1Gt8oxPH9khsS2E2CVG7TwrDmdmeo29gaGHC9Gjb+YWt9dC9BEt3ri
PXOOiveysXIVXb6azAgG8l9mLSV3Z9umbZLdKhBamy/5bd8tKU359qnlGd35geUX
7VHKjSr2jGaB02N7jQi86drsHiEkVS6tXT1IexeIsYHeulE5oSKLWOUFlPZ3x0uL
jriVmXAapjnLyD3DadnlLep0jnHtTanrCfQsM/0cUb2bp7dJ2PQefSell33fX9uH
k/zSqn0CxFqiMzPe47ezAKyFwe8YgAIes15P0ynDqeXW6JLcnRsE5A5iedHs2v5u
olR/FFUEJhYz+iwFxui/K88zV/zFVd/LKT1IawNm3LGvYHKpEZH153BFlIIMzdKV
1wmOg/F6dKJ2ADOEC7shJ1mmYKjYvO5yzB0YjTAfp9ok/DyQVOJHvkQDrLiZMm9S
FDmpC6i3UyhneI7JMLoqFjQrUPnl3rDjRWE0OCgyMTXqnL4gGDkyWlWtHME4bMfl
TtVClrfTCUamrlDP+dRPWvyJIeYECHkAf9ibClgkxGrMSEjAZki9Ij9PML4dILzA
FthbxKzkDEWCaXVaoKHBPd+FwpStkspSvFMb4Xb2rdPhXghlFeUj5xQ/WOaEmWev
4AtQCyq+KZndRL8NZTPeWtO9318rJ1Ul47WpDukECGsGsusYSqliLB5Ij309hoHG
h25xfQYsIkN1gRGveKBg8SUnF9lnGuSQ9bwEe8ei72VILtE0eX5JaICZqBj9fafM
jXYEk598XYLQwP7iZ5yrlg7v7YqWdXnD0AWTqRhAELmY5nRX68nTiCz7uaW/7u3J
YLmKXcXCR0mq+uFtUNUD/kZlvpCvjDp4DLhm1n7V4FOgyY23vayyjjYAj3c8GxmJ
Pjo1QWLiR01HpITZcBfJrxo807UzUuGQURcVvctrCjD9qbu1nf5eww39Ng/Np/6n
nyzsNVMb6lyDBFA9qRZxF6IezgmmgZ+SSnpK/799dB17VzryEmF854LFdEiotR6O
UmljjHvP+gBzc/uiuclRoGd9qBTnGf7agZjIk/tEOsK+vAXdxfH3ond3qt0FRxj/
T9Oj1bpPHTzHSNY9l9RV7coGOIqyXHpv6ASa5JdJd56/lWXXrsl/DrIG0oFNuKlp
BfeRaM1n5GtiZsS3Bf8QGOe6uSAtT5/rCdCTj24lc509LNkrIasI0txd14hEd9vK
0GVpwAitioDIBxsR8eTV7pb1xztZQ4j5atDkiRVjKJSigPdRBhD65VTCvyykk+Wt
khAxjrQZsjyiQDZwR7/BJhCKbZvNS7mKtOmafF61sPLkpiw+svmn0qF+2Txfrids
w7dKaIMXh+rcTPTsoKS5KomnGWBgQmkT/lvXMJG1i7Lzg5KpuBneBTbKqPkoflCw
8zgteXAiPQGYQoAC+HMuN4JcvN8fCe9gJEKu6iR3OKp9IFmQemsjTmpyg8D7JF7s
BqjU530X605kWPtn8YUno24i9z/uW9QtBQn/HGgL8tRr168856jPHOV8ECGuyCas
ZQ0iS2/7QSfWkpQIJo/5e8KH6NqzkPKJZ85XbyQ2q9rIWDVwPI4taMtdmGycpK7K
RT82m1cEfpiPYSjeixkHpyW4vmpA5OVOsptgh8vE1N0EZFMktl73XEBkESiETCFM
DKIKdSJyiwElWAmgLtgshDjgXBm2M1ZGPHudeEBPkCzxZRrppHk4VV18Ir5KRG0i
nI7K70plyKQELlxckhyjLvf/AvjLDgObcKQoS1PYNqo8OSNbFc26pbSU6zlXyVms
vXKSjxO5njhoutg/sNmpz3LqDiCwvyhijpeUs48DAqJXtC8YDE//fEfomoZmNePy
VujoXHZTGhhcmw2EEIp6Sf8kI+BbhlYhOmUPa8dcuwwykTXIaISUsUj/Q4fuFHR3
BMS1V1rPvqkkJOloAgvHNgciJTtcXjXeIoo+l0md9NQfBeSM6IiT3bfxosoO6km7
XrYl7p7Hc189GeWdIy+TPtFvwE4JDwI31vAiUPhko4k6MRydoO8yTWJEjoC36hJv
bg0rf8pk9f/0rQVVgbMHcMnpsuHKswhf5+M0VebFofvkWndD82H0oxxIi+0r/yBD
4TCglxInVkJuUYOhwqIhD13Dpv56CACUwhKOCSsKrsLbjce5rULZ/hrnxiQUj7Rt
Lxl0LThN9Y2vqk5kn/mBfc5vfwO/cgDPBKxW6XO8I+21DE4MBgLSMVPDvQsfE1Tx
41XQLpZbdmn9O1gTmPBz2i/V1enJh9k5eAiOa1v6JMnOVgxgEZDnUd00Izu43DM1
9NNtB7uLkBgFCxfyfZP40HHkqLnYxOX9rTlvQ5TrftvIjH1e4pUzszRSRtoSBQX1
F+a9ozEGHpUk0A2jiDZez+6CB6Mhf7+eUbYsMSR9iYX7HN7/yo9HF0sLcHv+t6au
YuZTJpPJftBGitK+oZdg0X56xwYi9fclJ9GXjlZR3bxk6U0SvESHGe7+G0588IrP
ABbNfzhEK4d9zSEZNvB0zxp4M6CqQfyAM9qdOJu/DlDMTZryXoqkSNYq0+3U0gug
s0rMibLsnTAstXSuTd9yXCmRpwWWTyBiPnFblsOwdtuxWG922noDmeLHlav323sp
jSgmHs+87C/QazeDmnA8ZbkXp1zuDX5oKOS9UJ6rM2hHM1OOMYUnaHLY8+wIK2q6
CKClmHnbwTidGq37/Cx0o/PzAJmKzrnGOpZpY82yb4+/fk6e1uS7pxxWMA4nmXFq
IRlREN8oWjfNrDnoHm6aBonrw1zqLgRNgUw52QLH+SD5ItY15BAB5/YbtrW9ZFlZ
2byjMXJ7lsQhGtw/FsuoF9mSErgGRJ/Rt4hnjTCXEVD3mObtB1Tdt+e+J5Y8ufMv
8Dn4nrnRPVrU7Eq75kfW6L0cECgqQkREbd71UlB2hhBvBHtKQ/rwvenjkRUX424I
Dqf+3G6hrIh1jpdSCopboWN9NCdN2857E0TN13KcBrpHvBTyYcjBvi6/kzSvOvFm
fttMsVc2tEPzbuZq63JhDN062LkteMAgGI71yOS2JlJmckXsJtX8bDVvEdGn17UU
a65z7scklXVYXrz7Au3GfwhWfsCrIdB5yJW+J+UzVvDsiHRUFi5GLUnLH/u33TPA
S/Yq16DPh7uAMMq7IEjIQwQqqJcOyqB2P0fou3cgyTFF8sm+WFNg7fhUpJ9LZGH/
iAKk3KO+FZ6p/5JwejN9+frKZg6K4p18boGuoRAqZoTDjkmlzGW6GNcH3zCF2/6g
Y/aw2ul6dIGIJaYF7kIGUYNoLFmXAldKquC2eNvhfdWuEhI22TnEucBNQhgalOpM
23vF+HzzPiRD1FdsaON2O6jgtGAJPjNzgnjHRmDZ5sfjWPX/2biWjGl0zteZLz73
fb04wQi6wcoQvxWJFuiwu9g1ryKJ2BfgSHXN/aYIWmG+HesLlc+YcI8w4ErzsBPN
eckPQMmX5XTj/L2Lt75RPcReXji/H0rJDNZ6nXV1gxFAlxu8SKHmFQDKfZhs4TB3
9JTKU644B8TQwC07d8EIw80S3QyFb8lEnGMPeVFxNS5HlYXfUdxd4zMgA7PoOWdt
698kFxLFuduDIg9rUQnhBNbU5+jDQ/5mTZ64TuK7dfHpIDDUDeRWeZC4YcNIkAEe
+OXObMlNRb0yZKKzb3VgjUrhOBUDFYCeM0EDsfsc74kktajhC3Qe2TcZIYKKKGU6
Y3rkjE6RADhq7zQZ1znaXtrrU0V3lDAdyOFRYcC5rf8mD1Gjh2nW8qRenKs6+Ic/
xkpHEBhYtPP1QVCzSu8ZM7P/Yy2Zv3mSvODDwVihFv+2ClATiftNz0qWQNlOyQRL
WBYi8jwd29tX6GOMo8g1rgkmT/xSZ7hA6fjWI6HCg+f4whdzaxGBi67+pkbzYn83
m4u/AAtTBuG8oJ8JUJ520J8cT+RGrP1/JPibbtPxoLoOEYFsVvH33T/baP3eEMZH
D4Qf9G7PbT+oPrMu837YlrxQmCeTy7fWuJBCFaaWkKxaa6ZqNMA2cJrskES0aRr3
wLLCCChnOXBcDMMAZPE73AtDRhv0PJPSNEwt5CIH8Yk8qD6zpVqldLmtgHqh1sSJ
Tb5QJNDHzDRalUcE1MMDSrXfkx3PlxWkPQ4Ndc5hW0bD2v5X4kS0ClqUJ/TWoBL/
x1By5AHxWtFz4A5ZuukOz6D8S36pWpokquubJW1yWsw9eRh0LA/jTCjHCLrVdiea
+cfwEHxeFUUvfQld+IOi8b0tW73klOTSZtt2T7fqwStCSWsBoShdml5BHFa4/cV/
zunRwFJpjdwmYY0VvIopbAQUbZKSPhZ8ar2nbEEvXuveBI4BhexqgP7GzvAzNMyl
jaB3cl0902ulYfWW8LZi7E+DImnrpFFwxM4YKsRx8/wPSlOOnkekkx8+3ELliv5W
om7uU3zTcl4KiezAgPTjjQW9K3DU7SoZ8jwxZW0YCAao47bAXvufg1RP/htecw6V
8FWeKMoxWnWpDNiKzN1RLas5AvI7vZeaYpDFIvmEAR29iAhJ6MLOZ0Ibzjg053Ub
QXfPURO5NPcCPrbgXify35sX10uDrSYjgIEHyfjSSXiqbfrq+zHo6Bik05+HyOKu
tMVBbsh/aPqY5LlcVeVXBVlqDmFfogJj7AOvs4NbKJG9joGjGyh3ghXxXc4koAzl
3ipYIPbvhF7W8/lOZhyicPIof9v2h+jK3X1HxyD+zrtH7AXs70I/tCbpq6RNjNuU
qFK+2LokIt+r30TTtEGK2lxI8Ltva6+iADf7n7OjEi+ugNQTgnyLZz4oGmB8hP58
M3XoZoyYdSh6mHJuTwh5nN6cq3OU+oOO+Y4amTkTuEbVGR/OuyZuosg7AckuCn20
luh0jwUDapi9A2gJwiy44NfZZE6rJWfSO+xfjqQtR+mC3jHiUgfXeMmIo0xnTZKC
Ss8Hy2X7qzXrhaC18yZwlGCqBegcy03C8mdFjg+xaKdE8WdOcpgeouMl2rITyLic
zB7eXAxhPxj/QO3Yp4nu40BeeXvTZa9XBDgPDrL3JjH+rCbcgiA18dhWDUZlixh5
VCCRdgsdyYad9BbLUHWI+JOi3sQcklD8F7J/PIKRu7H/Cri6ODSsu5zoe2R+MR/5
lkb7hkkUpYL8K0w7KXAxUUoP0W18ZvhcmF0zJFPFrBD2UDbDJMG4sIOTJEb6uBE+
yAdpdXjM5E1cZM1EA3bSuFMSGjEIf800X4y5ouTcV1p7ux03mXDPe/gvQ+3rA17U
Y2qri5qg1UDMMuRuPb+bX05iuFUPHcIuWBlGXpVPGI3knGAULbu+bPsi753XswEb
OfZjTLvLr+oJ8AEA1GlDyVBzeO+TTY3cahJzdg70oOt9CLBJEljneJyOyB72mmfP
SyUXTKa7tnLrYgWs8u6s3vl3BEgwD6PnPA4vgbazCDLAU3x6rJdmqyqkL0kckBCG
xs+ZY1nRqs6W9CVLUNm+CwVFfd53b341CSVCaEM+GA10fxrHt3tkiHARiaH/kNHL
CyA9bAM/VBBMzZ9Prph26AZa61hB0tRQEl9lBlNomKylgjvKwtL/tbNizTzuoOAL
pZigH0zt1eby/1KFq+AQh6CIWTTcO3k94TZe8oI3OkkENoaZdqrvdb+BnB4EIuJH
+BUkE/uDBVTcGgxa/cqJEWMoqtx5iJBxuNBZ5jR9EHlOeP0BAZRXHGJWwlBxZho7
iSVRkuLwfdTPn17ti9WknDYTm/ZNu/zhRrg+AJAcbqpE10BJOwuJQH6hNl7ejoUH
SUVAxO6xXfap0F62Fof8D+aGzVbqfiK29943/Hh6AlI+kWdNBBLKGGhQD576pneX
1SzOpsaszl+npIap38jB59e1QsNY3h8oX19j1y7aIoGzI7Buwpt8YD/g2sSpDEzV
wafPvc66N6hfe2m46l+psNS9nWnmu83PCFrqBhpEDpbFuKdNx6i8QSz2EEXTvqtd
RGjykRDoB7+5QwRVDKS2QoXdqsqWy4FVhfQ+/l1834gOcuijCoQqzH6ZllcnNe0i
0L6S5v0RPzI1hAY6CsF7tOiKsxx9fRIEyOv/gxscaamRALED6FCaa26tqYDvoM0l
D0pD/dox3NmBiKlhG/T7IFhg5MGT8uCXrxUhD+qzl2MPXJMev+Yy9kC9qOEMK1UW
fMhVYgoco0YI2mIiIAOJWfxEkLcGdnMkqKW3PAZA6DmBbE8I6+v1G5EBWZrSU1Dr
4QTAfbB3z1VN6x93Mt2K0lzM7mrndrWAObqeIGyU32nc+xJt9ycExgOfTZ++jFBL
8itOmCHyNZR5oRXx7NLmZ8e58imAi1/zMk+RZyft8AVoGML7/i23m9zCtzLtKR8b
E60OrTHtNxOMW4YmyfKWHLJAzAtW+pGu6dAAAtVJNO8f2GqnbbP46PNxGPKMFrbk
gm9b3LTU6ahHmYsGFeRZNaEUvf/qfXsaYLGahgO8yQl/OeiZx4Q73u0ZDgbsEzIt
72TMfGwXqSAdWhTu5q1ef7md8qKbUHmA23At2wYIHlGfsPMqpWMm3epERLNObpzo
EORXxTMQmPK9fbADCrn9iB69lNYsNssr6hfq0cH2qSsDJfC6EglQB2R4vm7dxzjR
Pm1WU0DxM9drRbyJ0Y/SeryQUQe7yvPmCOxA9C/TwKKtHwHSe8G+7qobxH2zouFl
4/RZeHULyxthQQPo/HmlR+fNsj8r4cFcALHGydAU4QQcy21i+jk/yB1rsq+CWWlZ
5ynAlOjg1lq8B7HmgYGEBHzAGmC/dZCnTu66rDNBCqziGsE+aszZAN59eWzDhX41
WWx1CeG/35dv5jYVUvzaW9/3yuBNfqYfzVKGjfGniHAiNKvTWKpp3NIK67BUa+o/
eZLplG77mdVHPGsz4bjWCUlLE7TPyZdEMx7pGs7IsJ2G/sKjoeT98DOvc4xxvtcV
4WQWs/2nnQ9Z7ayIMp8OAa3vqUk9Fye5p86EVNMWlvQRnMK5R4+BXVRv5wQGTbZE
eKFx5kIjorrxB2iCmUzuQ+t03890hlJBtoSFBCqXyhjHWpzN76pgs9FfRUSXb8no
C7EcMTYV4ETllQrATLmvVy/WK4v2j1yBKp967fG57YBlvYYtTPA+qguUGLnadMmT
k/loID6ZiHUBdm0vyq6UIWA9VI3XizlP76KDpE5wnZRZCvxNo4fz0GcAw+tfvqnc
Ab7FyuLO6CeFbKcXsDWeMWv7oed2RGJDBEHhE1l1sgEUjd9ldDxlbfeTQugCrg7a
3nQ+rMCci4HhX9cGYtEDX6ZmmfpNa8Q0H/9B7sfwFhfwlCspKea7lOwyCkJWX7Ez
VsNb2zGZuVZ8zDRDUjkTl2m/binu0WMJCiJ9ZGtyQtjgzOVVtFmbOfE3rKLZzZxZ
Fd2ZBYPC1nP/QVk85JqZNEsl4hASBTwx4MKF5+AtoXizJuXE3gMtTfQbNlaWqPJg
hApY9xlBiNtaa9hT+4OKls6ZvvTQyx2ikgF8YNAHhO3wZRngn3NTEEZU/isoebwU
I/fD2b/rtUBknb86Hy7Di+P99KyFnxoRS7Ot3pQiDJnDvWAxMiTeZfJ/A4aIbSBF
8vQisvrXhvVWiRFf26KsqDC7DCBO+eGKvIPnL584BgbJSa4CfVPPoPveHwI8Nqee
BMieL6YzpKtwwAfjtbr65YTYEbTc++x9EzDMD3s2x9SnHKJb+ux7QUoykEyuxsIv
AGv0f020F49HeMcjQPJI4s3db/E4fxTxb30KvXbW36GCosQJOKZBqn8+AK1LiVrz
Fv5xsCpFaqYlzwZvgBM//CXppf+G6A6MxfowfYRpnLfH8LgirYpWl2iu2nUKpL3C
EmR0tVOgVE3+MnpFNWJDq15fK8Itasodl+jnTAfwd0LKLmmkZB4QaHwz2J/16k33
Fby1viSNgaBidtVlq0MPMsmUol5kGmlg6ma/GFLTKNNCp2RjEguogJRFUQ88BjyF
wHMVyhHhxGSVzjLU97CyYjCYAV+VHg2Qbav4s3RKmIl31EfZQSf4ZILhWMpy/i7d
QRNc81VigFz/hriumuRpYLD9BsoOFWEKCD0ByPna025uvVcA+iE9bks+uUMdgXri
R0Nm4STcVgj4T/K7AQoQvbbP+fuc2NkH+Wzt8Zs1upvX+BVg8HpZoWEMqK1bFslA
y8I5aLFrr5wYQXJy2KXrStJQ/KqCjtFhrFCri2ryNFdITH1w6DyObRYUOVGxf6B8
dxV6+MTYKOKMEouWzZSr6Mcbnhm2lScn7dpkW2eEDVXEbUzxKOoqhpUrQZg1v4rv
C6kS8BfHqqIB1DL+FOn+NBU8Lj6EXyaJkVEU/f93puyXJvGZsTPJIAUdLE9xr3l5
En8WHlZ11FEIHlc/C0+VMC6+OQY7oPMWLrfMM4VQFCHp6x5noUYSkMkK7t3vasXg
WHzRzsYnz19EAYBIMgiuzcG137ioMqX8Cvnt3JTbOLPqJ5M2HBVekDe+k36jZnsA
cdYxTveKSXm5Px+KED/2H8Eapme2qks5X0wZdEuAVOgn++REvjmrWvmy45jpndbt
yhocjBeYTrEgN//FpzyEv0IkD6MU9Xpo3MP7aZ4jZI3AOvMuioaD7hbAIrXd2/Tp
LxHdg9BcDFTdZcQWojIOfoYsSqqiJR1GNmQeYVIu1/npkr4VRmnyCQttD5z1LHMc
sYY3F7ZRSOSWYLwuSTuAFlOdVljlNoZoukMF4KBSVDXnGXffXFWMrqp1zJ7ilivN
eRMXgaaW2PgsJ6tGJO3YaegYjxGEjy6tQEkkMe1JCzh1UQah1SFe0EE5yNwkz8um
fnuKzTMS+dmGAafwWeMAdvFuHxmgWzRjSSJ8B8wULEf/ErydSHvGb8l95IYNj5XC
p4sZio8GIL0yGdxCYUuhnpV3fw/NRHYXMQXkMiojdjs5UvAorVypJOoDdCWzIDsK
Rnh3C9ywhctwA7jyRMJe0NLEfLXxJf+gBZ+Mzvu3eALyJ+B4dweDUSqCPtbpCDJE
WX3Jx0hNTAPkti1M+eeHDysokvoij0nZIy7D4YryCQX2crOgWstEt1S3ZlUsGBfT
KcJCQBidn0ag15ioQDsC61zvc0GUyvys94YIGWawMoiz665nXEZsrwFNb6sddOyn
21hKzubQ/5kLskeCwYnlW7H61KByVJKn7RmW5Qr4WriRBlEpsAyN+KX+P+xdNPZ9
lF5B22fg2Uf1O4i+DrJhWm6GTICKSqKrmfEMr7lwdlpkXdmhDcJroDlCls0dbLTF
hWbSsLb3y2epuNbFImj56jQtMztU8gev22KAabfYvdPg8Rsgnq6/E2VxridoLhMn
ahoW2uXfMpNdV3ThgwSfBJHkbad4Dj2Fw3gRnJgncm/uFxUHirwNQPKs1DQt3p4n
5eFAb8OD+FL6Lm8B4yZaOnu4wC4zXo7GioeEIWsHDInNMh7RHJNQn4iDevRtuy6E
njcPKxyNIJIJbYcou+75U+bMmtU8/Zlw9NAdSBjLiLTdo6fxPc9icaNE7UyI7bpK
Tq6yM9jUKKgeY1a09R7Jr1l1NlBHTGk/VDaI10nsi3cOTobS9V7U6GZ/Afj4r5z1
1jRtO3paAbMc4OGDB3sb4KDP+hzqIGgt8ahIUVLf7s1z2QqfjPTzPf72V/4isHXr
HK6W5+z5OoZEpRFMsVqjvq1A/cq4eFmeaBaKT5sE5vZDJXJNgQeBr2T9sckRJmZA
wBMPN2ChiAUTK83AeIQC0jNmTU12cOJHragIB/zbfdVlmehsqOWf+QZ6qiH/m+Nr
nymAVdwRF8eeRrh3mSiDqodZJtFK2WtTgs9ATWG8IErLkyvIrZwmGs3zfMAMhuiN
yAzidl7F/LWbxAgVZdjkEp85BTUT4SelXGkQXDbDz89Py4VF2nNfzwOHDI8csmLv
rJdRx3SanVX+vOMrKLC226wqPuN8sY5ssT/9SAhQLw/UpAoK646G+T4zW+HVXXgS
KkWH28gjpDUqyZLpqnhhN/IlgXx28R0ZbHZQxfpIBNo+s0ptFwoD9lLoWS6va8HJ
YjUs2cKjERSbwzEITtrFAjD34w7RWqd2RFiFCSDFLDdwnzC3e5Hr7gaSLbeN+pen
I8GIa6oMQ770crWHKcV5embEuhAfxyxqEd6/7qBjPjIjbGaQ2MBD3e9KolMDQWgI
V6iUHKfwK9o9EBGVIsJqCpOhVI3uo8lDQAab43hKYNVvHCNsx7shl4got1+yjyyv
b+JoAL0uj67UsEBQtLA1ZB9tcjmY5/gkKG9JuUnSXkUfvNYgP9mLGruqNDHtuSGN
WIvglYJnfyJsFagq8c9lQjn2iyZAsWmrWi0D6qZO2j08MIt03Ew3ebvdOJ304xUh
2flcE9WHAwXKCp0Rv1cQwEmTTFwzeZPdr2QhWM8sq0IzyP0nTW6VG2izQzhcSCoP
w0u1c9PghoxbSJpL5SNLTC8Sl0ohCyqBdzmiiniJru00h03JllTVZ2uhO9Kv7uT/
SG3DyrY24BgPNV6kbiw19234D+Vq4od5kCytmiEznWnGXz7tp50uVxjByhHhhFvc
mVDVlf4vcTVNHWiL4y3OVQ+J4nuun7/dc7CpiZZXDk4LGoElyhJDGyX8TgGX0B3l
BiHtaGTZIVwVBLsvnd2DxYKPJ/SFtR2Dz+wSCKfK/58C6TOHcj9pDxwhFrRwxcYU
KBcnfeR4VNo7o5Ai7BpiHmRYQLAiv91QX7Bj8VNP9NTau9R6b271icwvd1iWpXNx
ErzQCUUzGFM69hVsHS+U8nHCQeEvWZ8l9eBIb3kFr+g9DB8o2OjrhxhxET/DP9QF
SM7AiVun9/VMT/CC2T7g5yjgznrrSw7qj+SC+ellan9v6km80jGYgXIvl8CuhxxE
vH0hFngXjLUaGW87FQYUmUCNUwwbfW1/6QUvqjyczfeU0ILhsSwo/LwaoIzptweS
rulHmo+4q5HsJqxhd6bVHdLI6uNcn4uNtpRSZxBbWoUEVCtA6vJ/VdkKU//nEa3S
q1cP4wA6RRskYkgrcYD0iwCWTe0HwLpAAHrkZFYgLI7C87pxtxWMIx28P2mBABAs
xpqgmoW5/SDanvxl9927FRbhZBEbp7QBS0U30VsBC/tpf8M2liYxL4s6aBTVRnOT
O+8lCsi6YVLajALZ1vPV7T0ICnDgcLkasylnssl9SDkipvIzwtmEO6/SIooB6N5/
sxVtf6BxEVFOx/YFivfZkYymsBxw1nyMPER8Rs+JMbboHVYqwKVWbnscLHa3Shlj
NbsLo9DwNXZbwMEn78zWjZtjzQXPE4EAF4CU79ntx8xKaSyhN77z0vGugxDFdpKP
j2JH1W4CtXu9mDi4VA9alGAv2oh2b0XgfRxEaSmkD0Oi7+pWSUrFC5MlGmGNNXph
FF2tiaWj1Ue9JTLTWIQLtoj6KPllVQ2UxjNUy1S+npQIpaoe9K81eEMzUo4pJCyT
N4s9BKrp++nT4W5DwjsdFZU+Vrh77CpXQFt1y3rmT5mNxFFoX5X68nwuOipAs00n
/Xi8HRqCe2VaXFztJ6sP2e3snKqI6378D+q1N+VYMHjgcYu3ZWYsHHU7Ab0TQrxB
/Qy0zEicCVrbjWBjin0IKHZUiYQbPt1Dmu5urvSLZ3hQZDbHa4JKh3Q1u2EZfnO8
+1wjeZmQfenSFhYWGZsor87vn023pG7jrLss8L7O/GxZxrpkEg0oB7lBQdRe+LWU
UOwZuyGwIQ8IMVT6Fi3srT4iVVKeZL4l0dW4UxzxHcNkb+5cnxIU6Opyu10CH/9U
9vGBpyh/bMJFbHWVKniG5FRujMTQ02XmeIVueIhOpW6PkbmKFUt5nm9OdLmfRniQ
MWek/o7EnViiGazNHGaJPJRYJy2VHEer5FV05Kdcf+e6Vve7yrlZV7H6lAJp8+74
CNDiV92EpZKkjJrfzKjVwjYnBmKIVbcHQ6Q4L/1Q4MDwropXeFw6E/De0MI1/qU6
VvDX0xx9DWkf2GGAZ/9EN1tWNf1oxXiyWxitG3V+pNWpOs+/VWyi7eg94r/UroTD
dbeJ2kKaoMvWLmih8FF8Y8ndJSpuMjKskeRC/vwriWhLzO/360gKHu9h1HvYPiuf
wj7nIBU9ux5b/j1Dv3lck1FTrFHMBDP6X9zD3zsrjC8pWd9WJeIu9T8CS1H0YZ/N
ndQ3T/QjknyTOZwDmws6nFSCMLgKev0emnNuJbGueBphVAL+gA8CfIqKt3sodHis
waGTnZq22VLOQOLuHiGG5mc5+OMvypagtgcf51F9Ivgw7z6qQJRmai2sWI/zZVpZ
ym6z7Ya0kvUkWlywU5ze5m2amICitvEm+PVXtWzR6SwCwyuhXpUWjZWSYwkY2K8Y
mkQSrfcYhhRfSKQ9QXjWAd+ofZ62Q/NOZ6ksr8d3gt1Ki+HGroCLd5S1r2SBOAkZ
QUmJyjlIneTi6zDzETjxDLid0hIGq9a9h5tnGC87hA0ZUQiyD+1ookvMmq+S26IN
/fuel7dEJwyhOwmLAH2T6B6KtDGTGEROHUMf3Zh5xq8qDMJYpef/ZQ+HZOZyH5ec
+rHKYYHvZbNkeC5LvnmbQUbD/Pqc6wuMfEBSB9X2uhs7dQehS5SPiERqX5+q/egj
ZZFSmdzj1EG3j2a4/UfuEpDn1Xnc5S2RvCvtgimRbXCaI/ksy0ILRSsgPr80ruOD
6EStEJV9ZkkerIymJpoZjY2b5PRkXuainRXbVGQeN1CqLhfQnrhwswp+xhobsb+i
xe1kgOntHpZJQGUrvEoLASDnHHR8Psn1TpPuc1DgyOvsu3hiWCF74ZnUf7CLfi+O
rPSBv8B6JT1gCt48P8wJFJC8f1IQc1fJaGaH7yiZKWlBxOB7DCHvSrzdzLL4Bqdm
LtCgLOByisxHFaG8IN0ovhtjhNQcYbhD9iXzhCdipWhB43agiarBs2+E7xDzJF+z
FqMS8Vud/XFkaZ44Qiqsb5kzjDA/WikqSBZQ7bPg+wzQR0JX00QnU9/20sbTRzO/
/kVES/apnvy8eMJGUTuKh/8riuFuN2FKUZhcyjRlVElXOejdyWC6RXbBgqn6B4eF
xcSdiCeNECFhQ2l43H1kXCKiXbvGkhyxvftWeAfOhVptL6FLf6Yxu4rRygyaSz28
QbJx66pZPt0Nd9ZCFhQwV9jX9y6C8VZ65x72cGxmHTyNG+eprRnTQHzwO0vEgcIG
LriRsXL5zDdVYm1MgNnyI3VHOyaptTiKSDatqLmUNUmmu6uWTHQJ6r1q4BxBq+Bt
l1scjJNYS+CPgjxOP//xj7nZVK71iNNk6S3NcUxbYQgSdlO4F/PE3xwST7PsvhJq
TBk6difTQVqwPBHmxUP3MJWKosOhQffzxUmjSZr5kw5jn++E39vJ+Lz+xhkIxioN
Nkv0FWRG1vGJUQcSXdL3k86NBX8/t/TqU47ABXIS3m2yM44cmhSdh6ZpXRW0CeG3
OZGcaoxmba2DJ1tVi4PqOmOITPXEN56JEV/BHqFP9MJxJCigqDYOZWlhhl05gwco
gXGLrlbTtd7wATlh22jWPzFzsrXRVt58WzXR7kajJX3wMYUE5UCZiTs+H1A9D33p
T0pJVJmzjHxfS1GCIoD4UZvzZYiLyehcfpxUSn4Nl/4pUuel7nnWtN3JZ8gvjnha
7DjAVoo4Lb/2zaWsHJ9Jt2piokhHDm9kGqQgnv+Pwdzqdq4KnGV63Sj62Zdcf4u5
OCYJAqXfuFi3RUuh/sZHgTOcOw13TYyRuMtbKAK6ld/oIpZTUJsT9EsNB35QLvQ+
/HF4un+7FHleuhz+JDV4XMZkBHVOX1bMRccqJZ75JKMl6z5mziIYXXzrrN9cdWaG
KEIiQ92JEEYEPCJsRBrxMEf4PerH8jJMG2u5RYbnWyAabQKH259oTHJsnkeZTrI8
kCXxCG6GR5P6OztNRVuauFOVSERll8YGw8u5MT6H7ofRyh1ltIlgG68cHp4YW2oA
uHgU2FBdfBt9rC+NIXHdRQv/UTXTPMb/JZ/SsuymagCykoMTzfYVNqVkXnrx0OCR
Qt6yakJ23LoG2kc/kidjocSjLaDb+1vPRNt2xaU8GTtSwnkVcP/zWaI+fKUHrPcN
Qcf3aoXqjFvl6LZzYg5M/DwhEnJtLaUet4HH0+u6dq0u9M+GH3aAlVe4u9elhQyB
lPi22umbOBaVlsIJvIyPARqsODVGJ8OOfYz4ee494qGQJFmDWmw3BbYg+rL7YMk/
2smPJtU4vTvSZQzFZPPQcK5ZKVuB7sR/Mq10BdG1n4eo+fCWiNkva809GpdC3E+H
iFwFVmKqKtoMPbk6oX8iJt2dx13cIl8ex1YEEFZaojy1rTazlhiTQsYydOIcvGwe
fxSQSgNBy2mVlRowSkb/hwsZIbC8B6eGPNENXwPYENPsGF3/JWkL+Mg6orWjfR92
t7wIBtDD8WA/IhPfr7HVpD325m4sZr8ccGIMr7loMaZf1lKE9IuDBpyeX2DZPYYh
Fx6rpVYm5KH4A8ljqLlFPpF8k1IgUwhob2UxzUqqxQpiwB7nVX3ujoxjlyjmrHix
TSVRcP+SfIX7EDzVb99kZyZaE+g/6ZZma7SgTodQPeBsi6HvCzhJQ6Lshkvi3wmE
R2OfHavivdKJzXVUUywrVim6AyqEAVrQ92rIkX9V72OOASqerEqy9r6GcOkc94tV
O/k7c4tbTiv56n/o2yTKMuQUpxSIjV26ByPm4xcrHETiuyjRAIWtV2vYlzTjhrcW
1YHptPeD+SThyR4CWATXP1T6UT96B0BJESfyI0hQaxrr2tyh4uEMPBRINuFSEuI7
2mZ84X3NXXlEKyVWC3Ry8GCwsAljeuHeC2uTssEtuAvUX0JIIUPXstzJKwkChAoC
csAZ0usXADsIxI8kpTAmKzMu0A/YdX7Bvgz6seYn5gyWGdEyLgPuce/hBaFbgGCG
73SqmdSp5Hk4dBaGEh2Av7mk+nJtXvr8eljlXlmOkeVNPYptt0n0HTb5CvZyLAXP
Mjt55JRzEH+yC0SUzUKZ9Lwp0NLe3z9BlJcTW0VfKqqF6dcvAjE//GPIYd8gzJ03
6b3QrlbsyAIRaXCnnl9LUoLXgg0p/GOE0j9RuGsoK2szLvnrKklHjO07b/79wsmg
m32HI9tnIX75iICedXr2qXDyCPsxzGihS+6JzCqyO/xM9XFH7X9vqOdLwQJ+m1dN
xaqYAmof8Wmgf9taKXt3Mx55Hi6NrfOha2f1MUet4lMrUvhO5aUuZs/FyYSsE3FE
F8bGAeBrpDBnAfXT7frMq3Qcd7SRsGVo/PkoO/Sy5YZKDsGJoknMo0eZHKC7f6li
83G6X6rf9GQ16gO/8vDHKoqSXqUP8At0X/9rwdTTGgKY3Ev3fRSACZhua1MyHIXb
evmwd4iuGNqUDT+yjeXtF39o7Hwbz1iUxONMhny+MovXwLE2wdh7ibXOVKgmNmY4
jVEOfL8gxEqw95OACNh0if3Bqp0pR8IHJdsOmXKTPVnB9wcCzd+qAD2rojnf4CCy
oC9820xxLBQXHJc/SLEtyr+SMNp6nMnJyKjkiJMpIoYalhabXtEnhbO23O25hz+x
EaUrJtQFBskBXDx6kTRXXmaM0ZuGicWWAZWYpOGrGSHzapFzBaoxDca9uAMeTLcr
KA/VK00CrE1gEkPneBQS2tOzPFWVFYawo+s3hA2cvmUbmSFlDgQqOJQH5hbw0Am5
3FP5ysU0JW7VfGT5QnrsVQSaeHm1HhxkyBpghubYcXqe0rhmV6w86vkSjtFrGpBm
JAixphTBt9EaNnP3+EjjDTM1irYFD/QrGb0iujSm2SntXHCeQRWMTiUvbNeFRTFM
x4dfhSZQqNHj6RXtmjdF9IMYFdRllVh/GJpEqIbkyOHcBez6fdkbGhigjMqZkXv4
3klAqw2ookLcVPDw0fVgv+67QoIqPiGuWYH/Z/nG61fxHacgnsTmdUMZqBRI4k9F
F5+d2MkpmvBZm8Vchs/cYqRrWEGRAxLBRl2ikxkDlaHJn9+SHVkkA3nfVOQuoOk0
IQ/Hg8DZvaYFQBIbx0eAzdVCjU5acQWIvb+dBcQKN9e2rVZgMwXirpOUwJ7slHfI
m8v4M4ohYFJ2j/kkY9uksQYyA+4ui+pyq0DdrFE/vZnnQXvm51Tr/kX7NodqUwEz
ZR8qwzMeZKvwst7OGXhIKo19oZdXdzCn/OnfgzlLYmFypm0Xij0T5gDCrCFzpdh3
I05u5tXdhjtc6+jXkx0T8Cy5dCWHwdlymKsHV2N95fa47VfovhqQTmHoQd7E4apR
2OEWUziZD+h17Idmy/eG3VCmXEyf5c7yus9MW4KLXvL+gr2tBnIRb6ZLt7kEKfC+
xiC+OYeY6kxuIkbFWZRqrO9Cfa4+7/QUsyvkCcjStN0ovz3KjEHbbGypHYXQYeC0
HKD9ZKIGa/Mv0UbQ45sRQyNXP/ITMfc4F8U+9RBrkq/zbzsSvxI8SUjpINc1qkMd
O2IHS4YSDVilWm4K8TXiXPlHdXYTUaOBC/VXDyNEPvm7FbqRz0tzOv5jrmYDZ8/Q
tOdXGGW3U0xk5gRfC+aPrycvGnHkA3iKXKKk9f2tvoUgYCHVh7/MKptb4LjyhhLb
25veWiiCYvbh9ZWtworRzz55Yq8SlPiYiamSAnj9Ed7S2Rtm9AQx9HTxsHVKYovJ
8N9+XUW7vIKukCbvD4vyU6zdCxU82c7jrG4r46J7dt8Nhwq8/PPdKoJ/a+SEaQeT
QcoEWSKql3i1QVDqs3NmnFev5p2brHoHVjor3vkd8wPy5YLKXctz8qZxnNk8/7Gl
0sylC21mScGcmp33e6O38yyYO2RepfpDf/SBVWzW4EmiUflLL8c37PAWadryK2kf
AFpqbIvLW03SHGl1wqur7kfQ0tNqyXmznJZb8xh34BiC+iRWH9LVYzRKhKGTXp46
9MGEQhlOje5ICa1DVUJH3ngnWNZnL1dqUR7kRfpRL9wLeD6eJHrd5DdAAcE5Mfax
LV4QqGQEODYgRy7EUq1S24DWSdOv4O0JBwF4HMKwRqKdRkrmt7f9gNOK0yLS553T
APkD33RWkUkNnN2U/364DxfEqfSc/iawzm+gbQsgULdtOgChIQWnNvi9wed1pMNt
5QbnbwJkFnlvmK/y0g8WW5NlKIQpNJsNH9ooFd1BfdvAL7coQK7l+vBRiZDjoJPy
l9gix/j0WwJDjpi+ozhT457i71G3rFhmrMyZ/YvWhWW09v4S6i2+aP4j1tereGeU
mvckl8eYlPmse58s8HsWG16YDuCJliioR5SekY9HO55CigeGoiKM7Q3/7ajaFlR3
pwslFvMbSWiMAQqqvtINTjWHlf/jEoZhKoizMVOEYCVWfiwUO/6M6cNKiqcJdvn8
3AIRBJS+z/NdbGIZlG01MAEn/WmQO4ePQ8UYTNFJ+VCjFqcSg/38zDVHRAYJMXc9
TuFDGirtjAg1N/UYIuj/xlvL6akLPR8AVBuaqshAlt90HdONZENbczDPPMPaxWjc
nk7YfX5H+OF9D9Q4Il8ozT0kxBlGXbEL71/1MtXOuNAQ3AH/VJrBdu6zO6R95sVN
UqGvIYvcv/LrE9rjQE7TKKgtBogKehul95fh6SPViJ2d+DMR+CWPXb4a0HKK9FIY
f1Yy+HuA1fux3NxvMrmOZEFiRRFbW5RzeZ+j7PXLYe35bYXGpw3S1w345leC63MT
WxUXfcpO7YD46hCXJImCY/6Sn0Qvvv5kp2RjK43S1jkjbyiE0RmS59sRxAdPxNdz
SqyrWogDY+plGAU1eAHvjrGRbNWOG0z4XJEOqzxpLs9gYK6VFfiO8+kKFaid+NhS
0wo/XTbs3BziNzVsuHXlcem+6aQAuFI95FRWDXHprF5qPr55rWMIf0WCG1g0Pu/+
xkDSYY/yzK8ACgaNvCl4/aydQU+CtIU86xHShJcXHAZSLfuWhyguvTrZIfXlHK4E
pqPLjMt4dOZx0+EmHe/nmfxJPJPqWdQX9LeUu+d5HfefFdTVwpKqKRpPY8aIFAjD
h5pO0/HNju+JJIh+oxid8TP0CNGvKD+gUeveSFB1+0RJU9IYldHkBWlcQbhUmfKy
jKJ9I8g9JipKkv/gU9S5l9KBfCYh6FRXtfX1q0E97ybGcW5UrWv0hEEs0Joga44l
Dm3In0lSXg/Tqmo9dkpRXnPaua82M6AgicAQeTnZbm3gDeO17O4h5OwOzli/i8Cd
22kqyCL9HF0eaPvUWlYYNz/VTVbSU2AClT+rOx49s/+v7crMsf2XT4HyaWMwvD2h
SMzST0q2+LwptW5Q+0+OH09f3kYUKkXhC1MLeQKNSh7RTW7wAy4akfTrmP1skT30
Wcei/JoHUkEeTdoeNGlgL8pOwO54e5l30BwAcBigmLfPtmvD046bdz6NIz6b4y/R
33ws9XEw1k+/WUuaCP8zXOo1Ao2xzv2MpmEtZeTSd+0i6T+5b5nOQRtDIOqNojlm
FOF5Igo2m7MyzfCjQXbAmNcq4c72EZEOh4TQx7tmisTvdYI4m4SweGsBlIsZDdyL
rCVR7vKcW/+hUBzlDy4nWaZ+e/t1AImfzreNwtxM/Y1hW4sdFSsoC4PAZiE8iclG
3YEYF/SL5EB6haj25qxtYa6c5W37bgNQnLLUIc7tWoH5xKbyo3OmnjRwBLKtR1T7
sbxiNUAN4eZ9Td4s1MiMqHfFslcVyntFIpGroW4C9DkDNKySM/rpoWjm6SG09+0K
Bzt6JOiuGG/fbTYAq70IjahuYx1r7vuxYazaqfxckK5pz/xOZNmxrScVkTkEh3gT
jc+++zRtbZm/V4wVTPz3ZTSJPJrTYyXlouS+fXE0TrEBjUuDzBHquB/bCFOkPKQp
jcHQsJczo8QcEb8ncGYulPXPNdqArc/1gbo+pgCkm+Pmw3L/l9NGXeflmzRh+U39
jl0uFEs4KzzqOPhUBa9qcyVnzfA99a66ldDw5Qo7eFXrp6UqDiwKxQPPmhSp4Yme
Bk8Ev1BEgYh+spsno3ykOUeCNLig6ePH07c0B46UnPqu9tHV8arVL3iDhTm1u+kz
T+ktZ35v5H3x7Kzclhn5ajbM14ukXq2EbyUc1iZPEOcNUEB5/tq73roNPt+wFlSY
EFOBxELHfBkxqf0k7texCUgnvosuhfmuMKcTXPyYkwWCE9Cw9u42hQkeZVjufuFJ
os4/dQeO0JBiKNlIBc7M4gWOViAktQjY2PZ/fUQqAx15ReBQCdo4JGgGqyKFl5Or
Mo5NFqlmcDPKukTLTTBW1uasBrr8Y03iq6XgItuPJepyBlBwXzGU58bujp68THqa
BRX7iWxEoNnpVI+HuSTPo1S2Hr4Fk2Ja58P/1isyEibIGFxKNlgpXcG/GYBmEuJb
qGo433DrtaheVHRjbt2tM4xQQmNpijEnO9r+1TIsZbdIokvhVKbVakHQ0y8WAWPf
L8oR86beBV3YTP+aLC5DGhEu9lqEh7NkcrpX5w/1xVnzEHi/M5KYNrAbOeCZtiFW
bBMtIVUJsOgLNIUeyKOsmafSJ16NhYEY9RFH6ozTLSRSo7D5gj6A7ixtm+9341LR
7Ztk2F5RjypxKbJbH3nJi/uMcZRBXMGK3zKjlX+G6lbrcAwte8CmCD7wuncTxPLJ
nZNUYdwkBOS4/jStzNR+v0zKPUVp1bW4oJWPfDlEN7A0nztVlKRT6kSxhobZId5x
dEXYWEO0KOwvgIVhUOfJDP4CgUTjCd2H4KMzOCNr0ZOM9q1VnsxnfwgvQPd7JQiR
6qyf954+tMK8eJmie5B5PD/99JtS0PMVWRszPTWTpBPhJWcuyeNkH+Qj3ZexV1Xo
dJKTGjRMX39Ai3o8So7X0eVuRdi8Kx2J4ES/sldmXEa0OeUmS76lzLAANhj9MOl4
a0JzD+93CsGc8jHtIHaTy720XcD6UbKNTptHZECGvj6gpAxOxwaQVCZpwnaTs2nd
Upip6SAy+09AoKzq84D3o9RmW0kEpR57RaGlrQLO2yH1Qel9JW1qvKTCU7FJQPyV
CHT9dZrPg8ZL6UeDRdFABrRknf9VJG/9v7lXAdNKz/gDlkQT9B4RJl++SvIV08W9
LLqDMS243LjlTQdlUlJUlSMalAKcyFSO46eUf29HOO18iPy2cKhebzNku3TwshRi
Gwta6/V0nLx3FQIm5b1pbvpF0MF3zBvEywHRWKOexFZbYX5h4BNEdYWWcvPuBL/8
eUN6HFDmPvitoQvQxTTJTSsaVzlC1xk5IX6Oi7OENaxp78GCo0+b6xxLzkWFRpkx
UXNxQEUkLlCd9VE822MGg1X0L1kSJGKLqBGQ5Ek7TVRhMSNqvy5qd2Dx+Pwljn2n
iLGpeSaRV+MA15g2TV2/2Wi17jfkNWs9iMhESyG7XcCHY7oHCpDrPult0yG4+n2K
ySzSlX0SeAYyKtMxxb9AHZyFplS8HTq2CFBUgZOfnBod8y3Jl4B4H5ORHtKmR5yz
0nvu/U1ZeiVdFdiQWGMIz75+u6cDcAvcYXWTlOj1ofIPPx8TeNqIYr7K47JeBHTu
zvEHP73WTFbRr9x/yeqxz6e4iK6NMG9iexLi1Yl7ch9tnf/Ad9MRZjWPnBDTm9/N
+NP1l//CvAoAUYfE45dyc8cLvZnZFYSVtualiOXqeZ2AdbNb9E1OlMPvpzJTj7F8
fUCpLuS76u7gW78dgXiNWhX+/4sSIrBiDxKbGormAs7dVAnbiltRr+tf6JnywIo7
RZFiz2OlZfeJ83/Vr0DayooDMIKx9rfwZ/NfL1JBfIc2SDvzqu/tRezxjNdVgIQk
8pJBSeqTNsqV1v/vhD0trV4RkkcrHuqUI4pe0AMo/8rb21MdRrnFwaDwYm5n2KPU
mV4gNPGBiqcSWOYaoJizF8Zl6Nh5RC1LSjt7SJAQV1DzbqOv+i239tinkFVwUXy9
XwGfMaYbpR3J2QH9bbWa9PnasOSya+rCYJoiLAPbOBgIw5PmHbej8XyKNF1Xo00/
RiENn5O/+KzUwRDOOSeYqK8jlNZ1np1H4soL6dDIoU+e4dosAi9wlgdPshvahShJ
nN5MKUzEzwo1jeGER6AIBMuOT6MCxVL7QgPqvpTl9aVv8HT8f3OKXqyAhE2OcioB
KZeIgRSTDv7z1doIYC/SWxgVBrw0k9OXSokZ4VE92cyWP23xCU+pVTIKCTf+NSk7
w/8bxcWeyM+EpThhGEi/b+xJVZNHYeI+joJcgd7eEu5k4aQlacMs/6UH5pS+1MEB
LnCOHPVCH8Jv5rSR0dAeo4K2G8gqLXwOSbkq7HPvv5YxyPAMuN5bLJc88vjjOmNs
8Se3nu+nPz25UV1xT/7mRzJpeSCcdEpv1KhIQPg+zh+HqL1I1+eGDvFfyiMO5f3r
30pBI6JWgEl/6syrNXKnoVbukYBAa7bqHmn20d7X+5p01R+24/KL+ST/qXgIfl/y
OzLdv6tcFVqCVuUz3iGn6v5ZHCf3CpXLTRbqf99RwzsZkUwTOEpu8Rb7s5wF5cfZ
cZJLGio5wniexT7JxyrQee8CSBZTgyBCi2V5PFk5uNFmqMdESjWyqyB9SJsHVTPo
QymmMa+hU3EOgncxYefvX/o0kcGd2mkh8fTGjPgqxat9g3ESREX3DwbV5DMmPk/3
5bw+I7ISSMkM9MB601+hBWEfSbmLHN6a01jOIaGZMIoIe6URQTDa1qX5ItGkX8Mn
L1NYwoVz0l1LQYMXRSZLoiLTniSNCy4sZFU2+1Njmae3NUjKn4aChkLGG9LXcgHW
1HjjmM1h8s/NelQdTpjxxCFqYrLjKFpxQ2M6YmxhsrDPzVfyOfVIcYiW7gE+IME1
0Y4w5apMMIaabdO/xIY4SEuaKRBfiZo2FGvPC7EU9gatgJQd+g8EDGYly4w2xXF4
rFEyO9PiNXmqIV9VR/d7/SFwUKtMQjFlGJ5d7ZhP/yv/9P0TNW9JPg1Uq9tSrs9x
wcVo0t38V7esNMwIn4Woo+KjMGbqV7Kn4PFfivJ+Fk7KRbKylBYBId6NbKnY8cOg
gN92/a5fB3DHqmtMPPrwIz/krdskUacvnQujKtztcsA2YhvSNCpJT+BOpIRPD8ZB
FwtZzqEup6zLJKHcTKhcOau7e5X2LPRA6BBwgZv8IcaKzDlpBCmzB+tZKckR3/9h
Wg0aWa7rcVBoqFVlh4OxZcy4QqSnCl2QmirqA4T5fgK258jUfwcHpY2KpgTldPL8
pYFbI+UF9ewLvxpYmy5kmfOJ/DoECt5hq2mlcCWdVr1y6ovjmhhPYM1rSUP7ZAfD
rGMypriAo7g3Dfo/N0fBk02lLJHQ7PtAXBJHqmNhUSe180Yjwht+RO1g7FGQlVjh
Gcz4t5tia1dLi1CLgrmUBKWqAdZjKnYOUPVq0v0xwg3Ft8Hq//IPM25UWp3GBoDA
8TS+2XCWsLKvi+puh3SPt54kfb8EGjtaW50bK1QOpanNY+4GwyAvgisHnhcqvM2d
Jkd5GnAiWCf7yLQYLOimwBCZCnwKjCifE9jkCDahOSgeSuQkwL3NUWVsu6jSX68U
BOUVF6HZKtJCh1cfr2TMK+VdGKocH8u9dB/PZ8303SM4TktOECX6KOd+TmKVDJb6
j3rDKnl2u2ju3iDyJuyO04EVpyxfLz81Nu/btCbd8b8H7ra447RlcJHtmbHe0mVs
UFjtJVciy29VjjwbYltKZ5cSZB5onrTCdTbboitu4PO5wqXuBZZojhWr5ErIm2cg
cZfpQA9FQyGBvUbaRt+LEkVntBmryY25w0qqrnDQYHl5JLYtuc2MJVXAE5dVxs4h
9Hcnr8KY9KZhbzZE6o5q2CDxJhYiaOrF55CFzXhX3lyh33m0GSms02YnKFO9tC8V
DXXzJdfeulsYGeetqzXXEWcVgE8GQHsPvxIWVCRtoSMALuKQzZL8RrzTpclp0Jgy
dWWUoGJfzpA1QWua6pomiKQn31uDznOAjGyVfDwz+7+kfO7fPrq4iT4XgetoBv90
09c+Zldxn6uaMGn718IWU+1h7Q3Y2ysKG9UOrZLtABm4vYC+CRxf6yVE+EA1YuR7
MH0m5GjXijChyvoB4nb7JoHsHtPblLBIQrPLHbZ+mZZeQiYnMW1me4wAVtTnNppN
wW8YEBJH5TrcqcRLxIde5xFpPH0ascGotCKbcwdQrSO2lP5RVc6pj5uZfUcAYSMN
haFt1BJ/skVSWrvZQ9UDrvQQIY/B+WTB9Ai6Jn+Cf5o/eRwkqa2N/13ImJHh49fd
BRtdVts10wF0y+CR43xDQrhKirtczzITqsixZb/BG1ey6TMILKGYYa+m49zDx72v
MPfglTT0TkgDi+ePRXH5BtDu+zmj17mobG0h9WX9xBu05k1affYp7LanpPxqRJKQ
VMGLeC5BaUpmO+sg/HZSoQUGNsxjUX7/4rh8NpSE/aKnkneodMvWkZWmHT57w3Fk
yM4NfibDHh05fdxbsjauf4wUF1EbUcFIuyHwyFG+NH2kUJEdSIm9TXbZLWsDwSk2
zj35bk4FTSK549LgUfGFw3gxyTvIx5urDiy6s8OvaB18dYG56E3/to0yGLYAc3fW
vCljCiUe048r87PNoCvYnpVAkYfcn7USdPb1yUKM86fQ33BXPIpeieJoPTwRLbfD
vw8pwgvDQgPuyaYVfyfBu+/lrj0LcERuVL0FgoHhcJmrUyozruGmPx7kMmqCD3Hr
IE2EOP5QdSuCYsa+fHoYJSp7bhn2tvpFfU3dDZz0QqJ7V1x7SBPL6wpmDY3fx8/H
1rfOZD2flCIQnh2rfaNUpA7NMBkEp6CeQ96yQwfDZ+Nq6FEjKUbWD0+xp89DSZBH
W+whgHmp5yxo9mW1J/EZyDL98GgsFWHECQmlzYOs77U/wXpZwVEKVaeygEDld0XG
eZH1w3X4zvJe8tNLub6keCKrmHEk6d8PUbvT+Cnka8XqL8w5fClFua/R9qofqDWV
qAwh16wVnnHoOPbg05X5UB5iB9ZGuzMC9AP4JquNfi2A1BkllhuGMtVUF27eljac
nH69/jNA4DgMv2tQY2KWqTkQ7IXnqA45cn4ZNuJXxckJVd3RjNUFLu7KJ8ALgdqx
D/37IKblia7Q53SsFd1IRQf0Xkw4zsFZRKPargEr1N967wNjiRhKhKm/+wJicub+
k62o8yP0QtHOLm+6Fbe6t+heZpVPuTnea4thG+JLQQSoVc5qzyt5wpbQYAeloWQE
yrL1Gx+djJOo/k3T4bNd9TSmVPZ/ZDRlpt+U6nCE8lBXwXknWkAvozJs9pDFKrdL
u1nPmZ9LenJqj7aoRs6a4EnLj+bX+UuSGJ+Mysm3RE3S54y1sphCGB4XnLd7D0js
j1/ZnQkERn+1dRp+M2HInhd49CRd48ohlFF9Qw2VgwzHW0y3zPrzy7FWtGGpYyeK
hycUedsp3zD8K2qn+Qk7rgHPxkO6joEYUBUrN4h1r4WeXSPuu47e26Z/03vEULq6
rBzpcnTmyuhbjaIgSz5me2kBOqNCdcR24MFq2k4DbnH/j6m/m2VcTKFbAAYF3+ne
uBn2v4bdL7bm33Ub0ncHqeQt8L7j3Q0/ZBNYNi3CbK5e1piM129GXPsXfBy931p3
ceCeyNZQM+gLAkJ2+bP6vVTB6T9qGnBlUJcetFjgaYM0m2eeqE2IhgSJ9DtipLo/
tX5ffdDXM+vsHfWOg2FiDrlPGJKNvAFd/hql1aH57gzUDMG3yvsHxdiIXili1Xqt
9yQdK0wegVoutTm5wDYYQZsGRmW6sLKOtsKdb647rB2fMmYW//3g6OaAqhYQzCNY
vQd1tNGSRBz/WHsKyW6h7TrQCdf1fKtqZizH9XzLifq6p5fJMx+5mfoAZ9gzel5c
0qj14f2ppz26zkTC4UQgrlGMLIPZv2lI9q61PV/y+aNa130nDyNXEptRnPHjpJEF
6HBNTG5uCX11qaM6NZVINtzlp19rduVEzwDqc3hF8D1LqjV0HP8s4hGy+Vrgx86G
lMA+tbhrEwAaA0sObURPF0CTfGqNB5Opj8HaJvTxTbKYdpdjLgLtvHKXSgR+O5uX
LxLLYrzCV9VE1ZQlAbjJjWNlX/K0V7pWEgfeTrfUTzm5bTxlVYoIu25wNi8xmyIo
knSGV4zuMhlV9OemHBDGRzQ/TUFiJ+hr7rw92+xvpyB0EqQZOzMvsbNuCmIKqel1
5ANm1BTS64BpeEFnpYF1vQrDjF+yG1L5NgplxImp3lJXBLNCEbJeOpVqpICCVkfO
nEpVz8x+JNT1/amRlDsSexeZnHizQPFStE4Zhwc0BeFtqq6mhTPtVepVIH0Yb0UP
nww5XLzGdwowaVpX7+umiZvOftV3DYsLBA8QtwAqyigp1QS4pTBShYwjtpt9khzx
zQU6xX2Txa0VKhj4AJdqmSFN6jtg4UEKBtU7xo3Bnwmmo8Z0K2QnIFEzBYMbxTZi
1Z3/C/xFxaTdEism627IfNaFqQjKPQa7wPNkt3doulMdpFecWjDbqfULHvz6u5q5
QhaKEqXbWdm0yw+W0kxKPHFrH4HyRwPTOqMn6XEoURfJQTZ2scoqHVLZY6zm60Xp
7eG/SU1UGQnIeUIKrrl1PRtjSirjLb2tlMe26n9Cy1oTbvi90fgnhdLnfKhmoQwo
vOeAOgQbQo7WqNGKkoe5m3YFFwyqK/xm/7kUzebnP51sIWBtsDSo/AWHoNLyA57r
m5osRG3Z8z2o8KfXy7cfxDriEwXBlenhcc7JuLpmjq/DqOl3Y1MAcQhtyi48F1EJ
qVUse4mlbKO1x/KZsVtnlCck0Z5k6bFNTS+a1kB8+HBNAb8bQ/qKmaUdtLGpTcCE
W4Hnl6QH95gZKBvPaZH14AM+VcufacFSbz7+hIC5HNAdvoTqjARDlOV3p4bO4oBS
/1PVf/FgwphjDtjvfaQmm9f1uYc8G2pcaMT4XDGoI9lT+TJzLEuza+ZdoPWMMlW2
AfE55V0dtKFNSQE/wRborg736S+0oiCsoBj9RQv8izrMwMruPRSN8cfXZxGRkVdC
N20+bOO4dGsQmoH8d0fv/vTTwVL/ZfGdvo0vVpm+IBsMkTPdcCbxCrDMrEnN7YTd
8Pm03j5dWIxXex5BInztN1GkThPAHISfzgCF70kgyzp1GwjlwImy2zSFjCOEW16D
TVMUk0S8CP/7lHJ2PaFzE0d+bpv2lCl2ZbN7Nczbm7Wqu62M3fhFnWb9IEQoY6E9
PyOOgdLpOhGiSXB1fFX8xj6navQ15/UdohLv+eGcE3TEUWA0283gvJmCmO4T28PU
cXCkBdlOSL5XwkrvUMn/QSEg2FwWzrOOF9yIVAP48sJqG4o63MYousKkyAdyzRhF
N2oUzaAV0vShn9pKGR6vJAZTjz3LL+o7pvT1b/5wkFIEWbmwXRmp+p2MLKRB2ryf
d34SjjMhclmLhfmvLH6JehRNa7/cB22LCFd1Gun9DVObXL6DutYNmS5xdQQejJBD
iU9mVC9y6BwFuWIMJDRrhMln66hc/JjfVEYJNvLfV3kZgBuzzr2xDgPyeZN41Xt4
1BxoWravJJ2Exjzl9KAo2o09MViJJd5liYtK3SWdE9MgfmDbIhixLHy85pnJjZBF
I4t7FH7GVVUiojwwWFIUhFNrdCwu2pNywXGTf1vsK9mUuL5aaS42ra3O6P1ngKTh
/I4Vq/lxTpzkG9AtWXHxKP2ECkCyfgavnB2kEEn9sFdKCucpq7mHGV6vI6liyeRV
WLQYHlIzIzrw3wr2KXCwahyFIYc4EcsVZwdJQo1VajJnz4slnQtLSRp3mK2zxA84
GNBisIgDrokqhNget8RJuc0gYYci104oTfdYq6oI/AFgW6ZS+NEZt0iz2aslV6ag
vFcTuZAo55b8YlOyl8YprMltf+6m1MR5QmyFOZ8+TEEKaoaVqB2lIZUSc5hkzQIL
krBjtfgVYck4Y3XEUdUMaHA4bbzKjlWqYrJFisxE9hiPEcPPSr3wlMbR2yjhvpJi
6CJV3Qf+M6EKfZ+ZVjNpIlOqjfrd7GdNd8P2pYSa/BOkv6CiiqXFrq+Fz+goYq5v
EGuMYoaLx/vNCSIgUiNum/8sNb0FzBf+2IYcO8lmYC3v8kRgIDEJRczNlgEm0qlH
tdVQiYYWCBkXQbWT222QOR3YtFjYs3f9BoOFZSzBT9qQPGfqtZss6WPUabsHKbXY
8xw7ZQub0pi8OCo4IowUyVMBRSeyztEjrohvwilv9q9TuEmgupEbUPOD73Q9NIL7
FoLq3nQkG+6wi7zQzzLy1mc832b34kuBtL3rmC+4K5c+myg5qCL0OsY4wC0cq9Sx
/YSSvY2t4egCDZM0cpDed0EYK3VSl3zTEL92hoZlyN7Sxf5UKGLj0ARY/v72/Shv
oL9Fq7FVThCQFCPEzc5+KC8XQ2eY1qRA/KuG4dfpIGdEIeIgkoP1AbwPa5LtKFDO
+ahscLgA2y6YDk36uEctW4xCRSjhS/XcTPgGPOT4ldk19tkTREbdtlERHB9K0svh
aYAD31wHbvTcUq+EkPl7GtLXnxmEkXjlm6+tzHtSvdZbiBU0CB2BfSPmUCQalNAd
t7C7402/AmMYhJx8G1A4FnBuSnhz8X0Gkza7SEXoC+jdw59xR78/wbE4r73QxGMG
jljTXLNqPVolWZmrXigYVdpEsI3u01RnIVGOYuLFU+5HnmbVJu/ST7cN6vyffVh9
rJ+n2sYmmXu7EEj/VPYSupRIkU9KTdv84kyXkOjlU6Ss29hvDYqQxGM7ovtpraKZ
sOpleSGvNugTMd3H7gcXBbk8yqd8QgK7janzKwVZV17SKEKR5y8jDQemZJUk1d8K
dOl7mtbH8cakad07QC6oWrJmFHxq8Sa57tAL2xmED2kF5ufSI8J9xY3xnWc72b1t
eAegWOoU1DBvia7MIuJ+Tt/imA+PdEo8+XEB9sBPmGZG4eYVoFaMby3Z1L22PTC9
FDZmFHvONxwpYgmMf0q849ihzCxGRV3AVv79uGkzDhGMYMFGB6yFHrmuPiyfGK6d
bFLIAbrmQqsPILU/MNLaaSnPRnj70wXhU+oddsRssIztMiIS+jMNldQf9O+cNHTH
eDqX/bVIY8GjAC9qM7XjtevbtEFn1sHeznWoniIi4n6C+rHEnwJwCmWl9+fxlU7K
nRLJGRG83QurgwNu0fPgL9YGluN/0jeIHWnPC4B5drR0AhUmenJlk0zNCUVEtwQD
qZOGKRmXpMioupk9oi0o1bPyHIy2gZrZRMhGajNWh2U79bE2G50w/XWk8fWP6fsH
7YKyevOeqS2Ylv0jkuWfY4IxsA8mAaQZRdNEqrtdzN40sKuSTLTDj4PvNLmBPpLO
K91eDJMto/L112HPHp4dNkp4bapAg+FcqXpD/JFsta7fbtdoRc3sP5PPQMnzFMuW
SXx1oqzQbi083NjgSmO3QNsT0giIyfzzOqerO4Wqp7rjffbB/+oxr6vHW9/Ke4Js
NdknUtjja3CA5AjmJrRx+YxkJFjIbmnu5UWEjshz9hOtCPIo38GXWKvb++ca4s+R
0TI4JDxHb/V0QhuCSkcG7ca7jjkDaH4ORgJA1lO5ywFh29LrgU1Umg2mLPyxSgXn
a8Q8fpRpqgGkURi0vFt/HofVRSrfzUg/tm3Fqx3KMbezVUrxWTbFjz6PI5Dl6NPr
JzFhttstNKgj1D0ooUMCamHVrcORfI36UV48Hyk/6ZebARk/WRliuJUacCMCOBLO
xk2/8htwz/lABJWu7rRLyDtFzLa+4i2DGT/kmB7dqUXCdMRBX6YrojuvJNVJ+Vhg
3mAjg3OF6ChLk883ICi74A0LLBD0D4WKbd3nN8vkQSWfl1zJl9yCFPaU+4zKC7VD
1q3ux2oJsgkciaYe92Y93G1Wp4ou2QZ4WVBu/ZuqCn7F/HJLY2NRp5FYqDbOBmKQ
9tV5WBgYS7SXNrmapEm7+xb66mus9M5Gl/D+T7Mo+bFJKIf10efL6OJbjHLl64XM
vV2+7Mn/khydDyIvcQEFkMNj6FcPKql1eQOl/GdtvqODD15/lHOncYVY0c7wcMl9
j+c+uqAAjYjaZf8PrA0VzFmv++DT3nUdGXlVmRlPTgDx8k90BoZlOzM0kywSFm1S
mXgBK6+OSc+OX9T1Td5zHanOw5HKKoE9kKwu7/51+EaC53l+q83U1IdAqMwkmQ8F
M3pktRZuT8ccW9a4znUX5GG9HYcEW+slB/sP+fkLx8IMzEAdosHnJ/Lgqmi/jBTC
EHNB/vP4r5ey6VbRkgh6pQfGIlPMmb6WGYpiuGl5RMPQWF89EEN7smjjtN0+qbIP
A2BXYhZ3MRr/DyxmZmKQZAB808eY9hd1Q5bTSDz0DHr7tI5qiSu7x+bMWhdBZAJ4
evL2YCYhZ5KkEWnziCklO2YOW6fQCTQHgUuFhyw6Mt5XojMv3RrGt6dGsjkndpoV
/qzTgBfZKPfTwfAfDK4//XLhWh2UNK5WbVVJwnfEcplmls0yOPzNOEXGaxTnFE7L
ytd/8ZHeZT+GG0biOEaXDJqe8PF7CUTdRQ4hq34mGj2gBSXVeWi4Ilw+QZFS53O+
Q7ADYNvkap/gJCo7tj3SFgeKaP7gIJrRIaGEUPKrxGrr+xZmZ4M5jAAYZVn+k5oi
6mtoSuC9v2sJDd4L0oj6DWNqxZJQ6ae7TkoRNxuyYPnKsorU38j4tVkSzEgxJfsG
63NOzcpBnoMM7USvcopqnZyXi7uZ8Kv4qQr5D51SbJz0G3XxxHCRujXa70Iexnee
JCouHBBoFTIWfmSUy3oEncrD2PiDxN4jf9HuQ29WWTlXnu4kZx7CTQibDm7LFI7H
dH0coq7/Xatali4oWveBQuEocIotMPUt92AIENGGgtk/vnyPROKghZ6Y14Mh4mdF
ONsJGLL9y9W56zIRrKuyNLyTuLop1LZ9QFShbEF45b6CC4jHirKDmmJjBUj5WLPo
2g2MJjPBqqJw9rZqkyB+UsxOwH5B6N86k2iiE6PD5FDSNn6RRxxfpl4XOK0VpE+Y
quhCA2Mdt1/csj72nNVEkFgDdP3iKd6uWZv1pE8fCLhGF8zUFdO/kUTNTSgvTa+0
BOSA2yELM5X9XH4vFC0DcVK2xP5XXNesZ4DRxAQ/B5rMU5kADH2b79DvOdUBpv3T
SNmWp7G3uFyOP/aL1w9JhW/VKyR5poVFc/sLAaESdFDGNqirLmmWwSNLgw+/zN9S
qybkorL+Q2iqWqf3sXP+71fRejP12To9cMXsRlDLjuOSTdSynyS0gL3TZt85YklB
Ca97xk1J0ZUWFipcY36jTjoFGKxAt1Mn5IKLThMqXXmoMrdnKFtkmAkTQrS8ZBPI
RhTxpmagbKaYYsW89xyw7drH7cA/h1G0KeGzINj8MtnsDdzLMpb2pK1h7uChOBir
eYpq3WtV7ijys6feUzgzbPvFaZCyr25Jd5Bx4w+aFL8MacY994oMCtGr23niLCM7
GQfcw80jXDoIlW0ep48Md3Ywg+QEfXVcAXNI4bqijNWZ9A7WrfvwlzdsKNjo5UbT
E9simzWLIsprbdMTwDfB2y4fyBy5BwTJO1tFnT1elgYw3ci+vPev04kwcMofnh7C
wlKrNc+vyunQZCXRgS5FuLQtscRFKjuoOITUWukJ3XEZzfHtap9/JCwzT1BeXHK8
Yt/z1n1ghwx3wtrm8Xw4fyv7izKyRjayeHqFbxP1dLENkaJ3lZcB2Di/zDpMaCr+
sOEy74X23YpDZn/lyIKYlCE7u5KDDQSRJBsOx/GYJ1fjr/Fo9dgmOnaCO7sNXIyb
ppoFa1bpFreYbamcTb9Tux5yq8d/dfGJ9kYek/4vfYdgthSkCkpAmJBQ1N/Yk4Ng
TkWx+uSST/YYNKSVKTtYd61Yb8BWkJ5/Nn1aGhnqactmCu1OsKT41/8EvMYeUOP5
E2MTXygRTliTy49RkqGiydNMifjy1mTHk4LFf5Hp2ggfM/jxSRX3qcgu1v5ydM8X
kjovsQqHr3wGtSZG2t/3pmCyWK+c7XCdKVAyvStJe+5s+tLXczwTDvR/eyXxFdQq
r3TOMy3f+0UKWNd/0YWr4+NXx95QbKxY8Zi5RWWjDmeTTNB1+NviebRJSD69mthp
8PIxx+GnNkSgeQ04QZ9h9FVxGJrk4lmw9DfQj4TMU6ntLA9E0BKCNyEBXSs5sHKn
GaXqr7klYD2tsDhHDxUtKru9mYmj4+i9RJlYqileCk1GXEqDnOBK8Xz8E5P87mlH
8tATafcUjSGoRGSaQaWZFtFJTB45GgUmgVpgz+DpOB5guMz63lCx5XvLsrbU1gEH
+RUtx9BPYkJnhrY7gOl884tnEnVHMKZlURQE4dHbzfBcZtAM2H5z2UOS5tmMH6Iv
n0YkL+ATLznwu94Is/W+lrqG0PEq7CZYF7hsTOZ3nxYlLDFXH5cognJq/MotzI0d
EXdU/y3gRsw+DqjASFprNTUBWNbe+8ExCBAJW8DKXS/Dnh7bOzST1oBB47zcED/S
osIudS7vPb+t6FQU4+1hN4b9TXzsj0b9nedUQzCOD+n+naO6AgK0xq3dZMr313Uq
NiqAe399sZXWAXdayeiRGKkopAHvFm3AEwRKY11p5OwhJ9Tx/fAEnS+eO0/BeVfb
9/6AEyyIOcOT0gqwoLfTBHeHRNu1eChFXoGO2xfhcj99kJn6r83Oe43mpTuZ1wN1
sRLbE/S9PCz2+60KeywY+f4ElDM9Ib08My7UzxKyiQjiDaa/M4D4Ke17dopKmrne
1KoEnbGA2ZeXHC05XJk1+niVRss63ru+H5oShudiZaqvRUIX+hQ6UGzClSNZQeZz
UrhMeWLO6an2RzyqIYKT7EX+u/RCZt5gyIzH3tAuk7jRY6scipxhkTH+sK2YyawU
yVY1QWFUPHaiwWcUlp4F6T9nJC6lABRskGgPSUrWgpsi7BDPrYA19DU8y3kzIbQv
sX6KhYc1jy8yJflSI+1gSiycae9lag9Hn1CBSrR3P3FTofWMeqHQsyq9KQDhvE+p
8TwwggIEZznuU/QkIPuYbF37oyZm+Hqp0nl4EYFVfR1F0XdI+GCSjC2XktkJRQcX
kZ+inccOCwtyYYBr4hNwwjkGwUsA1uGDEt/nr2ePLnQ9JV+jcSoJ7CNmA6QlG0jl
2e1/KWSIq3wmzX1VmmyLrskbNEuOmUvtgcB5d3bORtrTVEChYpCeldAeNh9+sjjP
C6v6cgbRjjBuO4SYjfC7O+Wrg+kVH7ndKrLo8LXetAE99q1ksgTqPex8K56QE+zc
13OGpru7jl1a0wA88OFH1Bz7kDJdkZK/Z+JRJF40rFzqEZTLqZTR1AxOPzl/aRpP
3kjRNJkqH7/tNtl7z1IKmLMKy3KZQTtywMxjeUoLODdTcda24ECLi5rxh/6QTDoI
aNus3sqkO0kt/Duhljo8kt+ONtQTRwTOJdDChcT1rpLLGvnGrmMPA3CiHHSAYqsc
s+yhUSl+434pZhfw8Gxtz9JjtFv1ixoHqQPxgzUX9+yGkd1bqZfQqsCXdY1jfx6Y
f1fp8xs6scIVP3+h6YTwAhxj+JeQNtivuvHWgobYg50lTowqBeTqhoB0udUIbsU/
mDbzpvuaAiQnLduaUnu2rdfQ38e6wTcfmkokpJy+N98z90ZJhNPP2DySeEsnrRre
4U5vzdt6UpKVm7BmDj80aQlJ1LJhv5utXuAwzGe/roSV3HO8JYSEFf4fdzzMAYUE
aFZKqJ+pIp94Idy7+NAFW6vHaNJOn71fTDOazqZ0chvjCquWICiT85T3i9S75nZd
Yr9yYMIcLglaeycDgidkrmLGU/9CxqFhz2a11FTl0LKAg5N7s3OazH0QuC/c7KOp
UIaIqWKEuSJU2QDh6u4SHi1jGEUjkTxL5nGc5mLflMnYso8vV/Slgs+PHkbX3OIn
W+MpdzQSJ4FoodkAmJhzKs+s/6TlC+K58+tvuhFlMUGfBiZOyrCc79FpLmKijXTY
oqsZjti4aWG6zJ3cUJqbjTQO+CCNIDihycwI4Vl0ZNIQKXEruO96OrEikPACG+n6
sYUdWAsJI72UateIyDPUrtJPalDGYjUqudFzKtJoUgWfH/YtJLFJ9+yKRXl88NWA
8oIHNRg1MZEAgHdH0vb6baSmqfHiz7x2QUOMuB+UfY3CuBrt4XOxHOwu/b2B5Nyj
iatUtxPx8cDJhGGuopHZE3XzO28fqvSx0ZUyZvybetbVAL/PVZAi7lEJLMOxVxWy
EYtbwBMNBKbdf338+ceoQOixibtRF1SFHmWEE6yDHcPjjYnAsG0qMkdsuYY83ldE
IjsikpHdHA8dvQUgKR2PT9EqQvYW6FXQvJdUdRpz4KexyZaxillJlHuupg8uDsRU
ZLC974B84EZGxJYmnU6lt1fbn38WDHSu8RUVYWpvUKyoWaFNTUVKpaSms6uP+kQL
T9F4wQH+SZOgAqR8VdcmNS7tsogrNLcjL6oUHbyiezksMNeID/r+IRmY82ttSrtz
7muG11UdydtTr+nhTA7ziYy8+dvm1aqaADu4p/tlp2ZmNWXppGKXPDiToTvrU2Jf
vTOEFlx2O3qdQ1id6piArrFGtLBIHkAG0PWNx6HWPI4mYNWrzcWuETSSakChvcw4
tx1rAmu77gjv/Dh6UVdn1qSqtUTdcNcp4tt98G7e5o+LUoQApD3SKBvDi5mF58t9
VMffIjvKa+inuvkjgPX8Ul1bHzaOqBwpCWBFnqxXR1Wyi3MRixhm5maV/acyTiOY
D8OoucxKe1EnoHWpe9Hhn6efa30mS1LqsQpDiBS2IzgqzEQSVfpkjEMQyHuYqIfG
Yz6qq9LTqWQLHHYNLCtLhzgbauQu0PIah5MGhGOLoTvtpPoc0wIlChmrUEflynwi
K//mfVWAr/HML/Q3UJB5QBwZkx0v1AtW6Y/yUYs11Cow7OoTpFWIuO40S8E942Q5
4IfjeX1mPpyOh8C590zWUaXMfDH5m+iyqebGGM8Nsu9vDZUHyoHkat6RGZkVapYr
RJICufr5Rg0s59aslleuEgYx9hU0m0LtGPxBTlcN7noK7awUqBzrbWH1TuSIcM53
H3AebQRXENJg3xYG3OyMJqIEFN/v+vRbUNYFbgXMLSKCb8R41JRU9leyjR+iongE
QYheKCouGbP9lorW2BpyBkCTyLGVg73gYEKkqC84CRpMHd9omQGuJRPCiuDOdgCW
PsXBolqWb7wqY0EnvpiuVJOhR68xBn9TrsFwlxw4IYUaNUFJ53mNKUr9CivMC6gX
0rCovmktFcHusYz2+UceDh/SMXf6gYMu4R7Qdv0Y7zna540gv3vhv+WN+TXC9Rba
wWcyHr1u2vfjWL0ZcDBkYtoISGqRKwT1smtiYvWUQd75myMXYwiCuNtJR8qadHys
4u/ayRqUHpP+ggppaMVIXOccAGR4E3QJ+v7BDhdSVf4kldgJ5UDktbuMk4fWLlZ2
FQssGrOiKy/84wElySt7p94MIycvQw/2hqeP3OiggSb436WVS3TkSkuGyZYyDDfu
DmGt0QMSx3j0ALXOOA5ioSbwo6TrjkCSexX9V8DiV8bRoNMTBCgW6noAE87drgrd
mrQZrqqGKmFLjx2DEBnerVi9htnoEycd0g/otninV+5gQJRttYUmY+Kki1CvYbyQ
oAcD6w19a3Ek1eKkC8XgTZ+OegyMJCaM89/BuyiZLjYxwvW2a4oODY01bGZoL1an
8ON7W13gOo2WJdkS9O/oxinvTIT5NXpZrxDp72drLmybipxPmkmickWZ0RoIjFp+
haTVUhKa4o7NiUoQF2hrmvr74SmfQhSiGLTw8m1moSGZ6sUI4vkNKazBwHkqBTs+
gYUPBALvv/1iM+i4KApRdLchzaUwQguEAC13fRp1DHMIgQPZ7VnP1Lui8xX7X6WV
y/KWRn478EDIAHmBu+9vPZaJhD8V0r+oZbC8gkT3o65SiUikHV1IvAU6kuVEf42D
EvJQWrX8Y0SCJm2JGivJKMjENHG1fzLhb3z03tVBMzBvH72cjOL/9twB7PJFwXx9
znuFK/G7mMYBXZALfycsMmm0RtLKzv5DuhFgYwN9uANBL0VkzvKMiggYl6t4iMPH
jTq4AgV7NbzoQgxQha+mPo1i8/eBt9mwnr55zLylsUgcmQEs7IYnlTtV7ZdAWd6n
PxcH7wlYghH+LThe2vuBM6qkEga7AvMxyaQCjIgEgK0ls9MCIqqVEeW61zKQ4a1I
fKTWy4/UoPDDSx7aN8WMGPWfpU5mJpcbWmRMR11DZIl+H04N8lmbwIDawjWJUSKo
LxWs77DB0wIn9dOULUG8O0kBoJyqbrGVPMvGz/jiPCQCsAjhtlL3rT8SpnnLgdjC
XdJYv3KLdzEy+zEuwBHD1xPhezdXcxjQDPWe/cydjfhjWj9gy4LdLUvm97IrsNXs
66/Yr9rTRT6zFvbuM+WE8/T0VmrWorsbUuPDeEsTyXSg/0EcCcISuLH9GIY7hdjV
/MatueLEU7TyR9tapuTSD+8xd0QWS1oPPWYx4hF6AYinGo8u8LAUbkxf7f3kSRWq
MzQ+jED9KXDv4WNCGvjhjuwdtrIlJkNGWtMLbfiOdB297MBb4Cmp+5Xt+hqo6ZCS
TDk5SAi/T19Pw44Iu880OH9BmtXqZwT1Sn9TQbwnXIi20IkMLQ/47f4o2didrg6h
xMOWpihsZLcVmQWdL1/7mxdLRQOpzAtk/PFLzMzEt1lF+Z6ioYE20THuregVZgsn
+b0Cm2rUU1LPPRNlGT5A+ezIQxTaJGDMCtPzrJBDlf7LOxjAc/5heP+BSjK6++2j
c5NjHmvaSWntqDHTShb2dui6rFMU/A+dWH7iiMKd+3HJZ1QHB7ICBn+QtDzLGJlj
9HWLhbA7N6xTX9HiO+xgQydROEuo//VC8WHkbvXCXtciR15s26zizpae7YDnaYPY
bn2jaRFvgLsbv8xhyRDnO87VOqhkH4XAz0LjQtgvzojGhnp8anpCtT/1rLk71E7Z
LhIaNTuGOUq4fTJlg/S+wiU8x77Tz63kbzTuDkqEoZbJ3sCAvX94NnH/vcE02+mp
KN5naePIqpwqVpMmPxT0MbOJtrZe/jvFBKX9ClIK6dlG//th//ao+N+l4SOFCdRt
u4G8Bp7FEfc3JMC5/jUdtYjKIbzk5mm3u2kj09zMxoH1urEDsiPPgk7Wo5fs6Jp5
Dlw3+XmVpCCLT9fsNTluTHY3N2MSvIGIH/JVAw9+RsaVVx03rNvgFH0pbXAnY7GD
UMBGMutxyC1KZzDeMRipvZMlGBXtJt1jaL3waBwasaiIZ616UfVZsvpoP0Cd7/LN
WVxIUr1TimAQLX6/g+blNdu8tIPksb088puMNU5AiVAZrE93TEKidwR9sD1B5UQe
IoO8z1Y73qFeqxwp46qKFpY1qHnwrr/I2GM/W3Z9MvdepwT3YqLdPtvFHO8rXx0V
lrFtIkpAVupO2uel8xT+30gDN5jmjI86UcJp00TAWohdIT2sg/b6Sn7/hZh4MHRm
vW6z57+cAK9cw7Bu+jDKTYFnvI91vlpHQtn+n8c7WsQn8oEWo3bOZtd6biBhIl51
jZkVXOALtC6sc3ePWV27S+Zj7mhYYFAT9vVK43pq5Xvf/8mNjuuhe+c7BLJX7y4f
/+agzwWLRiZBqFcrONnL1YDoqo7qzTII23ES8ByWayXITxNnmV9l4Lr4nENH97OZ
vpzSKWXdiZJTyDsn3JaTwbEE+sxZ4IZJaSzJ6AdrRC4RKcWjKUYETuDVD633QwTE
ASn1LITnGWB3kRcibH+s76OClK8/2VO2wdKUF5z8bhFp10trrXp2pLAeK+BVPL04
YJJcoYdyeei884egWi4OlRshMfqyFaek2CjIXQJ/TVg+S5fjr8YshuY6qmnh6Csr
Nh3WCc/v3FZJn+DzmfJ4fm8397b+7k5PnFSoxwns4Ao9ksKHd4+CBHdx7RhOQSur
6HZi03Jd1KHp6gT/0hZzTkEXtqBDgJVTDpXVtEBBAhGt5MGHMw9WUJsHJjlGc+xR
N/iKpKMc6Pgu7YGtNj1B+XLF29pb5grHFaGBGWNIJQnu+FVLxxLXMx3nSBqk8DzI
ftGn/H0mUw/qzFBZOUPJZi0ZbM4XIuSPQo/46uD4A51mmhythtEh5mrXFGCsnTSr
LiMxvvidfGsKcmJtHzfofny/XDwAmPMh35gWlR7dsC5Dp8vvJgPze68jwnXviqkq
07UbJh3T4bZ/WWpxft0FOYy2yrgAZzix29Pi18q1QfYNqgDwOlUMBOZ4SRkjB+za
74PlcqHYzRmP0Fyno0Yamv//+VFAzI0l864cbcsPTFhb0Z4VGCPejVyFjjG2nVWZ
KZYXAt5hz1IXw2uMBXStXR4pwgbcyQSwmUZeHwQASxMIhU+SrS07AbqKDhUXiR9O
3cF5XxrUzZLmAybLXegUe3Wwrsj7tZHpx7Q5GomF6EvQpUiNs5+zwwDAtRcRbFG7
3y6WarOisi3SDvbb5eHTtyqyiXFRXczBG5khBBhBwpSLID0GyyyJZlKvoOwA6Y08
AURY8Y3k+gXhs9Vc8J7pXnRe7yRhQ04rNc0dcUU/uATmlGbX2Ze3I188wqtUwiq1
osdML7eubhoVxbOGWvy3zKhXJIhpDkbAeTh6YECWJ39Ge++YiLaVeglM8Q1XcePy
atm4Xj/mz+thW0k0I2pYw/TPpJQ/lJPbGrk0SYzLkaafSL668x5SXMhAsJjY2km1
Q/YqtKjSfNYEwcbbbFmHiVkGmZVMctjnR+QKQYwJxaqtfmeXYjUDkyl0F5nLP5WK
582bYLdWN8+A/c/jzjrIZaGyz6nUFx5hX5d+AjO5UbCV0VQgG4t+76MK35++fiKN
eD4/X+g7UO8XPRB+3s5TYHk3OPiUZxXJ+XUj483l6IjpElbLrAB0weaSoShLlJOA
sa4ad8US3mnyH/puJlOS17qmUwl1907KGvznqdxQMOuGrDEZT7RBLUl7k/QjpWBW
Z9MRazeElVAuIx0iiOja0MIr9n4KVhNXKmL65k4apJN51RsnUIkvTYwt4ofhxch0
KGBl2G4y2tYRrQVg6L5cndLeglWOtj1zY/ftlE3Tmd2YvEHYbB8DpW7TLll2WmyK
2AdFVZ1urqHBeAFrikKBJz5Wj14Gkwye3+4N42fLvI/lYkGblLCpQ+fPlXHubfIZ
7N4rkSZa/YBB/4ri2ruRMNOsHOsxVeriD2d3b27kpev+yfIZ0x458wVglWEW1gvT
h2LUZKyBVGVweAVb6n9qnuncY3ykV8Uhnt9DMlXlceBMtziMMBk7FBKD/HYD+zVd
YrwpQeOvkp1GPJN7rD/4/yHSRw1UuGz6g5tIDMsffGIrTqk7KHaSEATEKZcf2Bk4
LVOQ8pY63DC+p3Ib6LELmWnbllLSM5AxlUVSWvxWG9LqSjOPiBhHR43X/6+AAbBZ
7RP1xfmxhPIIzjukJWx27lJaaNLKhnXMGbCI4G9g9piBGUutQAfJefPUJZMgk6et
z+ArXSp7qrFDouvJeY+yD3chDS7tgplTed2qk7nWdsUzj+pIBzVaDGpB+KKI+Zbj
G5Q+QuAA4AX1Fd5o4zabAT8NA+tvSvS1bE1miRIcuxFmIjysV/McXfo+Q9piibvD
jA4MLLI/6yBILHoedENpLKZ0LzroXoO9ngbPqbbivD0uvmIeMwOdYnQ+pJfthYdE
x49nDlhUeUhDE2H3DnvidSPX3PJEFRC27L2026qGXKgdnukc8cZEAFcr/V2WWF8h
YKLa5yzIHQ+A4l5UnhPf80K+bMn+kTL2noi0PQch9hIiF7DEB96pDeeK7AF5Xerb
VIuVD58S6D7ipAPVqO1n4D50APnsL/GeOn4QDIN+NZxqy5h8LNv/oPRgtuIM9G74
1BzjgM+6aDNGtKtI5UbyP2+BQCaeBXmkSVLs4fBnHsLJGUQd9YIQAOGSDhWs+mLJ
Wzpi+wBgT9K8CNH08NHq08glEVQLgdwY1nHM5sbXv9DeFDjWRwx+xu67AFeS8QCc
kr6u74Ul1hwl8xAmWdyfMOYTu4D+dqI2Uum9MlokSX82/tRoP4MXccTDqBXncKWY
4P1lm1OUulYCFsHv8PKnAc5ohww9LyPAznE86Ss2CQFXRT/5o+rjy+Z05J9veZf0
Wsg7jq7DIIvxQotPbYgRYEPuD5uLGmrvbxMojn4RozBI8F9I6g1oPwAmSD07nS7H
4GRrQHonCUFgna8sOsX0yPVcYpZwC17jetawbDqBi7z9aVH6rT5gONk+JCreUbB7
yQ813Y6t4qgXX4Rl0zysWw9+R6sr5K24cYvyZ8UOq9JgAGv4liHf9gwxQ8cgl6bO
r4tXc3RTPHLSPwS7ZG5kwcYv324vzcvgmhJuvrY+ccef02pLWYqr0LLjNQHXCMEY
23yGAogTFTfqK5MvQaf1GQO7y3HgD+GZye91MM2qpiqCLURJmIBsA9BWGMXm/PAd
C9T4wKZlCvJybtUDQt8C1y9WhxL1XSzwt01di+UkLtCwAtLb4UX2S+0jps3KnUpv
iDTt1LpUdkDxHHOleEJMwuk4Z8Q9EyUqaDpmn7O5Y/ES/xDu1oZObtEQ5mQ1YUbt
00y7BD2avzEHsI3AR7beP5xg0Y+G0iDY7kAgh3l26pkBh8ZoKjQ0rCn6Go6oWmx5
qHHN6DicWrdOU87zNuDCgumlqjEFho89ktscWs6lIdraVpJyzwx+2YW8qoIiRKyE
WVxnGRngu52xSkMg3Q7IYJGh/ND53TR7Voj5KvsIpWt4SAFaCz0bwB2hFZZCJIEv
2EmgHWI6ir0YtAslyN/tEBxMuCBDj0mkAC6sKcse8jGTuSPDIWMt7jyY0fwgGtmJ
lniQLmgrs694VNUqP536frXOp7KhzehSXOjLdZ26Hcax7IfowmiKQQeOsjky2zbK
gPwGaX2l8c1wRstlaSYOBZM+LQ+qStXIDZL2cNliWBJlo1S97QqxxTAlI9TKjjXp
yos1b5jRrN87Eh4fp69XLWklyOhYmYjAuKBFUZnqdRsRPWSwH2hC+uEEdTzk00AN
016nm7rHZ5QoZxYiTnmvjCW75hYc/ToliixZL/s+syBNX+wtAa3ea9zWD/ul82f3
dzUC/QdpkEeV4/1m+rl5T73Hx/2azUeHLPUu45Gj08Qhl6AIawXd4mXi8yZU+F/9
V+x0J0AsnGQhM2XVkQmREYux9YjPyzGAGI7u+aQw9fiO2eyPhtUtbj0RGJh55gDt
cvO6ecwDeMzcesJdkuLGGxgOdUPREADDRVJIYrhtm+1Q0EdHFsKhxcGaMRPp1lKB
TRJlMS29k9MYhBWao2l1m9FtGP19OFgi/HRmO+tBX7zIJQWVs1d93bpnFFT2TanK
Ts/8mpajSz0f5l1hFAlwbEG9RUhmMyYGlnNpgdinXWIJQ3TDmhgiAGWeZKPDcUUG
ytBIvvDeMeC8hciDSsNVPZp+kYyaJJBC09sQra8VFxZPftolwQcOT/6ii2LWHOlz
Jb4tBcDS87GLnEbZ44tNx7d5slK9Jd5+AxHFxPyq7zmttlQcuf4Hc2qqJ1ufKvFb
pB1jeO8uCFHv82tkRbMiohO6qwWrmW3JFU6AYbyVlV3URtun0W+LqEiEJPCP7B4C
9SgpFTonTicoxdxT5tWKA1vwERoVxpwf+QCMOPZ8aaFDCogQ+DAD39Cv9GqKBB+B
yIOcpasxejTeqHMIEUya/DupHOuGqRN4bmLHINAA7zrGBFztiuXa+cptIAPM7yHK
ShAXUnq7CtrV+DwtxBkfO3M10CJenFJ3VvvFoM49+UMcxlOFOCqMR3MUmL15Q//R
SRq1frGiuL8EELQ045aAVAf2nWPD2D7trREkM31qZUWu/iX4tT9vmZaLKRuNmJ2A
SwF93siNTc+nd0cx+SxXkZoqAoVik5+PqNQ9DpsFIvCd43e36CXIRvbLJmdczDCB
0vmkWeeZl+62Rz4mieq9yXR80exc14w6+8pu58hos0wd9T+csoNiJVOMSgNRgpK0
e5KJYZyLKV1tcG2ta9zi8/10tzU28Ye944WdaiCebHKsp+XT0pmUAbz3PEms7pj/
9r1H9llAB3v6iB4BmCzfYJSj4u8ai6YBt4ZQTMSEGkX+oZ3qg6XuercHtjdKM4KD
BT9DHEca9jEGvYWL13oBBbvPtxY31d6nKXUEahlfJoT/6GwtMIWx8hIPBogQgLoW
4O8LxudOi5Q1YUeWIeRUIooVvogsYz9Esuvgz/mX9KbiT48SQcXn4Z5VvsXyzIpT
x7VLLLY6FJdpwc5cSdQf4pAyMtA6gwN/fSEEgsGxXdVgjME2DJq5XX+g0C91+AkK
M2es+M5GVCa78fjIjIufGe0mLb7RcwaZKGNtHTUaCyZ7jTRTe7VJV2P3TmHyZmFn
cPUsJ7gX0iSTetIPm+g512HgzBBKWdnEGbdcK8TkxB3fejFE7CF59AiwkceVMYpq
Rg+Ubufyqb0PT+t4Btw36HjNsjOpxIjPpI64TSMY/h4hWJ93H+2zEEDT+8kmo/y3
d5QK0FBqBbSEbXmzCD9FIHCzHNt/79ZcC4ma0XGNR1C9uqR4IpbaCHoFqaRiy3EJ
LpC/QaianVqex6xo4xc/jIsXC57JJKzzJvGwdT3hNdQNfWnlqZlc9IUo5BBbBzzV
azDXNeQqWav3zujneUbcVnf1N3ygdTs3excgZNW55wXA7Q0y2vFnkChSSsyhBGC3
kC+XjMmVs7X2GeN0H421uKm2tE1NMdzaJR5642lIffHFx//7orl0PWtlPmuvYJMd
dOUqSeLpt00lPxGmRRIsLYgtMnzO/lRMzMb0P18+gUUFQBlJPMjANGtJFRdofGTL
gYNXdtYDtlStf5jbQePlpGrUDOBlhcqs1bjncBPjbwm1p9aGU95seIAzDjNZSAqM
2wgPm1iBPO4yGThLq/25KyQ99lLS+ifes0JOgtr1XXNsrPhaGD4isrxF4o5XQ9m0
3yvKTsjaBIcmupLRWm2Xx6zRtZqOvlErjZkUB5RUAU01Qhar3zxytyVBMt7djKlJ
l6Eo+kFktm9WmuhdQp3EfwkTUBpIEwbKXC0Osc3PHk59R+PuW+y66CLvXx1yFaQZ
QVt8VZHu0yTXBGGdkz6/NRB8+s3ZFhLLpxnynCGaMacmQz2NR11zxh2lf9yQLvot
UjdfdbIGeLH3H0hAapiRFk/PEaTvarC7J/lKaWjJca2NhaKOogr5m7vsWDQGo/Ab
CkyfCm77E+jXOTUxRCC2AUKbTO1djFrgSxl0vr4knMu8wP8oSf7Y1SVkxlY8/wjc
cRBTCl+uliH9cn/jePMs/ERKWlN/Vc6TgK3r5rny2xYTFJm8xk0cLbHWnIKsKpG4
0JLC3uxwhUuY4w0prRZ8/dAgU7pX1aBKHXKHYXwhz2s8yRCkGjtSP1KmR1283vBc
VKHEJ0VN7fwnfT7RRV1cLjRjWIdc4RQAvtGWcInPtV8yeX3Z1Y2x/gKofBMbMEyJ
Cj+k/cq1tq0kPsa48rcuYIkib5gG1B/kLEVogJkz3h4XJpvtwVGqaF0fOu8LPNTV
6HPgmR0BsYcG+S+Rws2keuAX2Hx+m1sH/1UTKsN6KTvEhVRY4mZFF7kW/Ig6xUCs
DMLdfdQDRUGpF2Mb+oO3D6LbfraU2vZ51ch5wtG/0mO4CBCAU9rmIy196OqPZVa4
T+GkEhtVD0xd5mnmO9V/hpWTs7nfiHK+yLW6/YacM7ByVdyrP2+mabdVeR/aX0Wz
WwNyx++9HoIRgoYTszbSkwCUABS1t/7ys4LRjYX4WWCnz7EwCfMw2CbcSrApsNjh
D0/Ik8JPj28Q33xYb+jVfgXLcyxAFGChMF89vzBeCvjAONH5dr7c1fJZm8IoaVwd
SYEm85oh7Rn15beZ7/tH7ga/nxSFc+yHWue0utblcODwAM+dxfk6Vl0acv1DwSnK
UJdjoxfufAGsHH/eQ8lyKrZ3VjujIu8vQDQHE9p//7j8c8iuF1rNCHmB1GodsbB9
b1uvIkpm2sEvNG4fgPcfqUb6/S+EZtfMLoQXWEjq7ibnbUgeO0FYbMGZHJxdfGdD
zHVyS9frIvckE03CCucP9iBNh3KdTnKzezCPfpnElyXAMjRbjW+oXoLyXUniWZXE
N2+syD0Cfqh/GliqOTjdXtnzlaE8CEvEUfqfB69TSjvg8hy7i4VtfT8RFdAlGaue
xfPlX1ApalYIUS1SYTTNnPY9RGlpkwH4csjOkrlmK2ffuavbUwkQ6Dh29M1x9Am/
kK0dKouMH3bXt/ijwm9vGLmYdAYDKqZAmBxdE8MTKgSSiTnJH6vyPV0w9BrTgIfe
ADnDb+vd9snKKOW93u8LSKTzLd90hnOXHCd2/O5yX8W+9J9obUDGW0DHv78qsdch
7khtL0KG9za/tv/OERPe5L507Zd7dHkVNOciik7f8AX6LHnSs8r8JvCpMW9aH0eS
mGiUqqDdzoMO+fCkH6lZEWHtmI5C8e6fl8OZYhpVx5nCykRp2AjUAdUCQZrNXRlA
WwbccNhGBALo55H3f6YeqV79NdulmQgjlo3Bp3tKEiJAb35KAbiaaxiByqdDMMNv
rFsfIXyyl4ggWSBEh0A3XcIXAKbkUDhVEygEchkD8mr8pcCyXllA2vx1RLt6cU5/
KpVr52n+WkhCSUpW8f+xMznJk0Z2kk475bxN6JRb1zLOGKKvyIHexQP0tnS1SN7k
GUWFdLUL/Dg4LkJE6VdI/aRN+aV9cj7vzPjkrGe8Bf0+hdgoAuNqyyi3M7DttEpY
vJYjnBtMFtZYgiJuziBo1CAuh/KQ26Gras7H4QkmjE0epBdFpwGlibWNYJVROQQt
XOiyYdXq2QDkNxDu3GrrVZc4oCvZg4e0buF0lGI8KbqGf+kx7urfYjERx3Kjkatn
7XUfBhYnORODRsRk0sxUtso0ZQgw2b25sUCQRI68zMoFcAheluTyqiKsBos75bqJ
0YRSwIUzOj9bHwIzanfFz2XXdKOITgxbYXlm0gSW4HNku5ydbEvCLGFKvTkoAQWI
nYJ8nzQ6ttlWYIn+M+Df+oEsKktJfIF/Gb0bdulSZvwUtEolwzNheMWPTs2KlQGb
I0Z+O73srevozJJCf/2i7UOkCVuKY+LbzTIFFeRTv5ZMXnuqr4WsEKOBvi3BNUji
Ku2TgfCdnQfLcehY8PFQoZQTvd9wZcybj/V/P4+vs8uTOSJazD0htBkOJfyzSD1i
+vsa9axrPEJztnHbFBQ4i/r5bde2QewhIVzNQiAxioylbn3azYZGRt8RlU0Oqfd4
5qncexHBaiw5NtXuzslCYvcEKDXy/2sV+iKW6bxxqHDsydooKZglvlow+MJw56VB
qoxpAm79e7jsmOukKRLu9iw8PSqXibYRv9oZJt+y0qu2RB3JFUNhtMeM31Fsp1c2
z5r9l0pgjZlHAtpefpIjY1hWBdOr0OFn9PeVl9ClcvkqxmttMOHXife9gsxx4Hjy
4fCghVGsyGk7v44IBj/YNLUjGfUQ27aYHwKWHdH6JjhkVAcPGwUBEX5WIidkHmwj
6/WOB/kpM+zFTcJpaIo3ShT7/tgDgtAsZUR7c7SyuSn1oLDWGsfBZYlJBrUYgdqV
AQAgaJdaYssMR4Ok7R0DtmX155oOAR6WGK3wBCGebQSnoo5e+IQQxGdaKF5QmZ/d
fhJ5rkcBbOqQHby6cOZDLkSEkOSJGEproszNrr69Wz7+ZezatzhAbFRzOsl6Cr2e
OHX2d/3VPlUHdzSB3dus6EBz54jhq3IIa7KW5g3qWqIRvh82lphhCpSRF5dtqiMc
D+Sz40awcEeTclq0WlPtGvPS3PE2fMOWSQyEiaozZcNeUrQ2R2AFh+owBzWMyz58
RwlmISwct2qCd5FA59OxwzXxvHO8mH3+7dldd8lhzCUyDT7TrqT4oWCAoTxuyGAS
hf/uZeNqPy2/wxDJ9uM87y3Gq814To7AiazVMWaU1EWZCu8JNdTL0V0aOSncWfj/
l9O5O4v/5BCuSJvzP7k+JBR3GA4b5FuWGrqE82rjwDmi883TVTBP2EMhKk3pfkTh
LmE613AWYUI3pHxIYbAXGrf99O61+rIwmONY0bBJHeskocpXurJ1Oz97Ptrsv268
Em5BKQ/6ISdrvzUb18vL8Iu1DC7QYhPPJlQQMnx1iC1MBKD2JUD5sqwXd0SNMDbe
3VP2maGDA2O4sdzVZZ0a0qI08arMwmn4QyA8h5ucSOvymnall7uidP7sPsQrtv71
5kP5a1pnnkx6rObZ2C9y8mVI4sJoVj4KiqjkMo/wy5WLRNnGwJLTgPv3r5xWmSQq
CWwuAKxf9cxNNO+mqd59U3b2bVkFa453adUZJcqzghC0lMaDX4cAIcvwBzWtoShM
TiAdvEf1fnzSJ5fKmsowAiCZgKxQjE5Kfdf0msavVMx9q2I5NCgy4dVtV8WHJoVp
gzBl6CdCP2YSUhHollvdNb7cZ5MjT20abtwqLkNKN5HN+T3r/p4XGDhMD4OBV633
ccCvmX5Ye3HNrRuj5WDiRvYRkaCPQfJueyXE7Das6rKmJ5q/iZron2flTHmfP+Yw
EKHdpXCB08C+njsVHAAn2Ap0XtQq6vmVMWkajS/AJ0fnDjd4e50HKqi9G85Y4lfq
3R2PufI8BkdVsLpW8144c1JTnDxqGlyjsYxRPfLJ0OmXAXkJ+xMP6y/ZW6hij7qN
f5SHdqZhi2Eww0wK3HEioIAmafEXHyidWWacXXTxPR+tLKj1UJ6RLeqjDCsGGOd1
YwyKye/Og+AdB5ZWFcvMIqdY73ttWlgGK3noAHJy/mpoSssjwaFsj9Z9x/03puNp
jpRiIsgJnWx/loQHwbKtOmWV5ci8FSE0Ehvuj7ra2thZBj8q4VX8wLMbXb97KTx1
WL7AIqSuSLrJZNgco083jjmI1moTV2EqJuuvwRFa8ODfH0Ly2LwxQovaNfmPnqb8
97Pc3duYtgQ8SQeu4iPev5YFbRzKT2k4hvRT5QXkqKxAeql3QIz5eO5OM7snrzaO
hF5PSCU78vvair/V8lC88iUkJNgIlWpKSPDGrIckIHcX/B4UsIEeV+r+ahQf5WPM
V8AbSXItRUuHGtf5LbecUiHppet3KTK2ETXyCjvuGTZmWzSGaPhGayyGQLPhoj6L
9tJWxrIbMk/2h/NPLmAfmWhqajRqVghr5ymmgEos7YVPUnd+G6t+V5NEjLZfvb6b
jdCEaMSX7oLiZYSm8W7sB8+EUJNZTBHwrPRCJ0ToY/d9rZj8tXD0O3gJwHRJQMjT
d8HY2sHroQ3oCQhi2+N1NIiW0lvQ+wH039YIxiDoc75OEcb/wB/U1FJb5nRrqn3P
6vzvEXCQuMn3tPkbhCZVcDxno9dKSAatJFYuVIuDpXOjhhQrFMIF0mhMLDU6UbE9
+JJUrMbLCUJmO5Lkazxs028PyaFu2jpfb1EKXsDO3PGaIjYMjpMBCtk4vCsSkRgM
rebiqrz6eTgkzgE6bzdFxv9NZQCYTEcbhMoqRXxJkHNY/4sPBKp0hvTnt+8y5zDZ
fTFaaij+X0K2WKHMV//3DZF0he7Oz5s5+IrYjkS1TB1tAIQMUzvHGGJnw38D0hYO
2YREwNrs22ga3Pf3qRF+5tMyXWtx270R47jddXsod3s0HCc3g04MaZIBSQE8QVKp
FioBIkD4Pl8PBtMvNVQwPjjR6nV/+9n/D8nISbRDShlbUG0qmKIIv88HAiKcvKqJ
yclR4JZo6NzNORJPjqFB3yXLAO8a4/a7f9MosVxSeuZ/a7ZWqGqf6KVnk/geHYeE
WRn+YMKYNwzQGHwMMIg+FZIPtySjFUfGJa/CFpcv7EBd8Z5GOwsYYHsf1pITJuPS
h0Ms3cWk5qH8wVhKSBNCG3sR9xZRsKLYtcSUpzw71Fap1PXX6n9QxU1brxTxSC9i
OgVwGu60hMaDpbPpCsD5KlpM9EjsAnpVg6fh+5f466Y36nk+29Quu5Q3WJW4CYJx
nAmH2+6iCTYSInsrcGcaDw1WXmKCvDjSmbNZzhLoLTb8ShCLptu2/LFo79BFu4+B
BIrC+uGNzNvkLSUPvUsbHGBOcDQ82AwEPvkYJyJcZJr20KiTNibi6AbgFQQNWgnz
KNtHbXMw1SYev/KC0oUUXXpUku+tZuFVeGN8b5wD7EJ33hVlwXZ1gh0zEueLzKGN
r3SuJTDpJhzTm4KRjy9IYZOfMYeSBVOuJYINWyCwRTsQ2JLIyNSlQtD2frze+XNX
x+Ej3bi08ZNjg847iWYyEby0A+F2KNSuBMr6WDu+4Nu0zfd7liW/BJSJfWUfmapp
Mo5G4Zroa6foBrHeLJ42IzeXNyXCd5RzTdKwUu6K3/W9UI+/+lAiqV72uAzcf/0A
sjcAvLosV/hgzh7BpMaYoTWUv25fMeByCBLpzvbkvlrLT1nRc3CrFgpK8zPJH7sU
NOD8tbHGmXzw3W4snmyrYQfpjeSRsI+ufTvwgoph7XNBqKx96TmsFhC4JP9q52Y0
2oKkxG3y5qkl4aJ4xNZGaLExx7vlhcA7ocw9iE/Nf4Xst5qe453OYp1QIZXk7Zi0
yKlXwvIlRFbxr4Lo45iiPXnectJqTkwGSvFEd3cWOKQre+lUEss0ERcNie4saOvK
3UWiXRxBKle33x+yfFTCTFkDCYBRnrq+s8u5f9FY2eVqlL4+pxRYkDZXtS978dUp
GufBOviFyRvxTo8J247KTlwYbyrhXinUiDfaXmGAOwcEk4yAr2PvVRAoW3Q3QkzO
D6s5ROjrbx0Irpd4rJ/TLH5fjdZ8gzyejetVDssovNV1v5OQDrrtuw86tuURzo3f
ursTOsTi0ZcbNWVyMtWk4i/owIhoh8UvNqWauWeTjfvEPgGHVavuKhVVArLOs9mD
w+hLgZbiOYDJOMDlT7l12WIyM3IZIrUVRHMFls1/OvJ+5KGfkbhE+D+c1Q+WzIWZ
otfH64dXPvwIjcEkTTQk26sXYBvhzk6NgkenuzLrVCPGq/BrRhTVp974FbrZnC4d
n6isglZ0+H0CZtSdU7FHNpRVLtzNI9qgvgik3QdQM8abxUt0XCKfyN32aO82d2MX
7YAE8w4qrMJb82GFa5x/DzPEsuh12xim+6px0jS8MCunYKLlHobgEl8nv9BxH9J5
vRwdoB+eWYhENDJBMY3e97cl8cafi6/Z/DvXOGNPRNC5Qg5Jfq1/thQKYgYWHkgE
9DChk2eC4lq1Bs67dViGSL3atr/LSkhxtiUZZMV2Bs8+4JuObwu+jlRTHtZ4bEjl
6mSxudaxYsDw41TtEUwOWEeclxXtIfyU4/3lXDlbgU4deqQYdDAFCosPQIn1NnJL
/AJFN2m9Hc/FfsCT5i8UkQmaO8bUsR/9PVfFU24RySrPpFddacnJSvrnh5bdldOm
MQQJUoADPR1eXpf/DIughwSxkFeaN8Un8wRLKJnjzu9unTcVjr09FiD/wL1PksQu
iQgEpiBD7/Pt1u/9IjkXR8dr9TxB3u3tZR0pinF7Pwdof0pzm0mM1QJc5B0oG9X4
rLBzAt4aBT9z8QwJdtdMUtwFR4giCVhP4Br0CjayBuqk2rkbmhBHTWnUog/kh5dx
a6CbpYn2yHyuDh1lnC/Mstco3CamW22wLC3oBgCYKWgs4ViSq6Z+eh6KpDLY7e1r
BXx28RNYo5qlRbLOvhW7ENaeC3jrVtz3BFZwAY5mXpTtvxYhq8ZM1iToku1U0NNH
k360I1aUN8k2cCiLpcRPBwKOgPdgfnWmvqLJcQRxy4p1+w7/C+U5yHf2rrpLjib7
fFCWvGJ4B+CqtnLF/5PgkfRsts+4cPoKVXZ/vMJ1HyJZr1SDQAAl/Lub60yIjhd6
ifOPOZCx+d+CIXwAOtMtbeQCkpaUBWEzVwD0mUbGmRKm0Yy/S2RXZ4FPegGW7Mql
3T+BwuN24PGqOA9ncaWnkDJydUPaFtTwEWCvQHAXx2VkyY4mGZFV8XGLHEzVV8vc
LghN/XdKuCY1Omq4gqMrlxJ9GzqVgICcSxW3c2tgYU2NgGSN8oa9JrWoUYukLKLa
ASkZ9RshLkwKcEg2pjkOVhtDCLbuEyl+uHOlaov3Nf0NKs20OGF8lfnB04fm7y/X
dMVLczy7AG37YqlAlEYx1nptIR8ehre69DgdNE6lI6m/v9pISbZOyVR/28LjfxhF
t9ydKt2d7Con+MBHvGfAqL2PJ4LM67EyT4xzBG5NwqqmycAZ3hDZX5eKmIgI5uO0
aUQ/+b88TLr1B8X/5qaG52F+5MahfTN6MTlJI4ptl/gpwV3ov/4vd4dO5r47+W+z
bu8ESFLeXIMj5sqVGjOO2VMl77wO6//749d/7QY0Hhh7YloDcR1Fux84UdGT44Dy
tbgQ1J8mGiR4TKuppbze+9HgWRXXIz6ex87hnHlCGqqbmAB0xbF5HVZAMt8bRdGm
ANwmkVdRCb80+KitU78wRUMiCsX9rIpKjTIFfCwWdsEE0fqpcRiTAlqlVuMCGOYK
X+jJErS7mop1GDjevm0voiYWilq3mVRYcNUR9Apyfnk1Qa6oUjSGz71oB4TDSbRH
CbWBazcq5Ondj6EOVI0bhHHgxF82gDFRMMvv+1lQLteiP6hkWAC2KeChVqohdESt
WCYdsAAJj1BpP1WaS4PlgHA80jNifPQRAFfwqJbpYHcAQr7lbR7okIhlgBnJCqac
e+LkB+gtFehPFWu21CghO+qc81eyzHpx3RgAY1RJieZWRpsLXW6NcW/TPdbq0wr4
ZEyXV1T5rMie0sXv4YjkXdXJiHPJ1/xPD4Lz26F1hYxRLVVnFLYaW0OI3/cdDF3/
IXJUZF183m8I0Qc1MGr70ifsL3leYzVjRpuoxZ7OpTNFoE53dvI9pEawPuNhBQXx
p+fTccxR/dAIheWJmO3UH33B17x8yLZKJlG7Q1LbZc0A3xdnVyMHXzoq5g9BYF7m
cLqEK6/Hai0ZOhq9LM+Cz1eTNPdMWYg+55m1jiNUWR+bigUZuB/Dd/mLjcyyJfxg
oBEGmF0Mb4h5ywUx2XNPIub1L7bajCEtETwhyO1oRsjcz0u3loOSJkQR3QfQ/xPZ
KTXavJXQiEfb7ztZdbAvIIRWt6olJZaTkoxvV5JUPwc/pS0wkQU7eD+0nyWgX2Rb
NVAN/Pzsg2Tsx+7XyVAp11SQamw6FgHTIYBMRPt/5aleUniPo8ksvd4Y4ulQEm0M
jawCrlvszs2fJ50HC89TfJPysMfTQKM16j9SU0zs3p02nHNvg9klntI/eGaCaWeB
oqUOdfbuRhtJ0SZBDo/ngDAFA5061M/CNg+PRewjSOXUi+iEeLMEP6ryHG/9brFR
gPnDpECpoFmYUhPpp2kUxQeD1WjRZf5a/llvW0JzxnYb9ZkjZMwIH1Z/B99KRDUa
gO2fu/mG5pNx5GUpUQ2Eercb/Zt/vX76RMIVK/VoJIeeY5UfSP6kJ06RfobSDqWY
gSmi25Za8FNeLkU2c7gv+aMRTkhIx+VKwtfaaPgBlZOu6X7VzDrU5YKcmSmr3bt8
Sht7kfJPZnDEOFZEJ1KI7eSzIgJUsUnLlqk/wTNGJaq8xru3YGmkbeVNR0IPcWhR
OZgiJhAQrI1D/6/pphYZYl0vBKw8WQp2WrCqHWV0ceI0Km9X/Ajxz1TYW2St66ea
cCyIOuADHOj8Y6IiCGnuDPsAb1C9loZshVge+FrrtBMqCoFoppqGjIKd04hE1ZZe
iId0ryN54+QLWQZc8pQzj7I56a5UN/BVhz5JgE/ZReWfPhkMO1TqTt5nXvbiIMm3
uLetrfTjRFASGV/XaVXpLI0OIRkt0n5cpCs9v5s1zhaGOxepZ1v96pJtsCRaLuP3
a6plQI8jibzm4el5zEFQCNcXVOia3G3n6ZZRjpxKbePZ7H9wpilvQ2SbFF04e0fD
pnXKSacrcHKA9pKXpALMT+rrZgAt3DK0xcCmQ6xHgK9dbWI9ia7QUNQTb9Fj7pW7
FpAK9Kr4uWGQtUEuEgV6oIU3fDPM5c6SHmf+PbhKf+60f3VNwMaUQtTcMvCglo2y
vUJDMYBrl140UgHmD4U7yx3R3CDzmvdO1MBQs2XzbXFZdlSjpbbJfYVoNpmK98KD
9Ms0zGY6FXpM47ijRXOs5wI8vl7L4/ZLL1D8qpEpJEflobZAqls9XbC1M/VBXLST
kKJFlKx0+Apzytzha8KwRpcVL3Hrh+jJa+M6X4uCqXUuTSNw1Gw0A+qvpXeMOv2a
PQUhoKIazMM8fTwNMYibKfbtfFBwd9rOHw1GKjvoRTAs49pfXSmvavaT9BHRP8WG
v7bXmX36w+qf7M01FnQFB69iCwnlPRLvBSlEK0sKL/8/fPlv8GhyL/yA5JDEFUIN
mXQmGQAZxRglhXtvtmS/vJfavJDuey1UiWm1Q3Ft5LQKo3kyA43ZA6Cg7iKKIIge
kxw37gPiQ9GFIAtL8UhHas9ofhg2L9ALAVgkse6Xr8Q9FbLbnwvWbcpfa0QJcZm6
9t5sICwyzp1HP9tCsGrJG3AFWMg04/itrgd0WYBqos4Zn6VQgjbZ/Y0xRkHx18tO
UFY6fIvd36ON53Xrbr9rOTcNTjq+EiorPn3Y6Ety/fJtylcWTSjq2jAUARCg3+qE
1ZFVKq/LrZAYUnXaldo5g87XNMdFu730jbaSdLFkhTYNMINgr/dfsmUkTlIDJY5y
LUMK2SRLsiLTnUVFzx8JAdSsWXaGnmeDIv8okukr5r2+DazqbLft/eYcMwrk9GZY
9ms8oDGo1ljCMfJawbvcwxGKPtwMbxC6Yx4b/AJpxFKatqE0aYC91owBmFICah/W
MpykxV7XBWbvidjdNms/We6MR4LphmfJn8wxy5a3IxbDE+iPhy965Ww4Wlb6K2St
BZ4rOIt+Ukrw7iDA+2NpWEXhBOTcEvv3CPIxuGICL1bAxNoIm4WtjU/ilT1jVrg0
jeqTvuZh7yc7MjO0LnzRFIsmABBb2zpxrStVjF1a7liDvH2JGE/PTnU/2nfQHqIb
GvkSw3ldOD5JFADmgiMvJMLLPHvyBdc/yFLvqUV45f0iYC2I0zFZOx9FSHttELEv
zHhjpdsSYmbHKecpS64pFxmaSOOc08wTDDUeKxTdYTQu86q+ftbdlFyVyhAigUxl
miz/2GeAVLOwmUnY+Sj31Q2qyUzHlnWtcubv40WGekLWeTrGAwv2Qqrz9qPzlsad
LW5BoCgzzj4CtmjIH2kF2vCjjEewcwfbjJsI0zJx7aIHUekbPYPI+48XTPhiEVzB
4hK16gGaOXmV0yoWgGxLKOHNLaD6MXNSCvA822IFClJivRLSmYGPFqS6Rlkey1Kw
0Hr5dB1xMT3ZFwyVfyw6IcoUXO8ahnH35PBmCrOHhNgkdiovIWaG8aDaG+RNQ4ix
fUJiISM2elv5tjPh77D+9gvopozi77G0/bgUFyS6r9XZQ66b96OeIcIeLKJeAUW3
Zd8wW9p0bUnKgYXiqmdI9sILZDlc+fUD5KAffQoyzKs4bB1iKwr4LlDalXTsf0XI
kpuymFNGcJVMS2cWxkSW6AvK+KgZQTkDgPCIMshdTUNT3PLoi7WjgLlHpRL4Trju
2S3wZ3Co61pM8wJgroinj6Wdwo6enaTRtRUw7dktq8rmWGmbRiQ2u4pd4mExxFE2
fZF8Qx61hwG00OmhdgIBshBS/Sfxg0ZvCEqIHSE3TtzUQ4fTCvJFDcDJoVvuSCwp
EfIaQ+Q76akbkCSZRIFZRg/0szCVPw9VvlPooQho5IcCQgh90m+PweMgorTSW06q
M6/9BldPl39B1MbGw/A8qmYkaScsxwoOZ8xM3AUNnx1OcFLDI/hBdKYsEsfPk60Y
4YGZaT4IFNS918bDgdH3AlIRpLVnlEOdmrDQIl7r309HuwJGwmtn6xL4WQffHXqi
oKSIgfe84kGvffYq9VPjsJZerQIgTxhIkTCHFGQjrTesjBWWN80D5eo0nx6dwElr
cmqhptCmHUh/E9XVTPCs5OwpMF4dZiM5i06PBj21s0ltyVof1IjYNj77KAXSF50H
LMSpiI8W0TEpaLBvHoCYffC2sAE2T9akQT2Q2EDpHNd4mFA8f0a9VLfP/ChcDbGs
SO232ft2LYCGtkvxNXchs0s5JSzhwVhcaBKaagY1wL3PWNpNfmehMQxEZtm4A+tw
3n1KmQ7Smst61t+fAHRs1p10ipxVn6qWSyA5X7YJFnPdzDN9b+5TJcrPbAjMTUbZ
N6KVX3duydMN7bUameBgFhbyhK7Hs4ElcIlsvMogrokVH32ATnpWy8mIh6x2yQYU
w45Od8naSpmDJiffBOd80uRZA3Yjw4MGkespqFGhzcX+oFik1P5NTN/7YIrmCvDr
QvtSoHC053TZmnhYZ/4RotVjyXMc/xTVHjJxJ4PBDnaK74Hi0d9GJ4cA17axXnFK
0xfRkYrn/q4jS5MY5x4wd8KWCK55LZ1lPvKBevormxxYtSF26FPc5slGst/4Kai1
91SSCqBYmXM+i4q7nZBUqpgi2Fm1IoxiRX9e5vkYj8RNWo3oBFnv4J06KLDpr7PF
vXw9xVWFxOABNs2F640NCgVtgTOUzSwvKoRwKBVqn+810ZUAlhypYY14V4uopnv0
f+l98IFg7DEbREVlVp6JyrU8GCn6JxdfBDQ6Tgeh6zC+r9cw4Un7xDN5P8PsNqNt
RAmL6Vye5WuYR7jmy128g6LO0QmyoIr3yy+p9PGMXLgjV0rJFR/IzQ1tm1rE0QhQ
JdYhS+R+ARx6jvYkJ/AyQjGs4YaSg3+TUSz4nkVj/7z5cftLd3sH9Ihf3zGGV/GG
PWnABU8ujDh6lzxuDqKy9Ixp6sf59Xf7zQz0Te1Hv36Zj5IkxSygF5t0UnQuBSAx
VAbitAeR0seEW8GA5FVNY4nZ05yvOyEPJrvZcKWxeiePVPpGDkiqfY5Es6oU7nAl
McLflv9nSiiSAA49TTE+/4tYX0EdSTQSrvwo3HjkzUAMetkbSWGEYD8JLU3PXIqy
EOrNHb+3y1nKmAfVwA8tpM28Cllbklmd17saZaX9QvzvyYRqGnDBcW0Px3ddWmCc
PoKxt3LWOKzl2iT9+O0f5zGSiOcHq/q5zkbobWU1bgvzLwe37XnwZp0hcQLPWzcw
bRIdD6G/DxEERJWhtYu96EPKFI5uz0onc1PCTe8kUUetvYp/7k82W/QIQPbKg3U5
LJzWW+8hmhnefKudabX6Hph+sfrwgqSPCBbzMf/l7kyaPz6umzxVsl8UU2et4mRn
qvOj+9e+JHI+oZjzV7EArXeWCNz13Sry6n5ksrdd2jQQ7gBmQcvXA9lHf1J2JvME
X0i8n5DqjjPIAqwYKy+MAtFGiNjfysZNQs4b00XXmy3YetAK6cr+ExATf+k85QT3
os5821ekLzyT5239YlxCN6f+e0kquMDa6gr7QX0MWjCM7PV4JHsp74dfYSavdV7Z
o6cDL15XYUrepJ4wKhZrBYZrG05KaEvZC1XAEPk65WeRVe7F9DVkcaAvN+n8v0y6
FJeMpnTNGjvfR9icO51IAgufTHhkFbcwomsHKUfOm5LZr1Mun3zmMcGC19Dfs5cV
fEL+wzpqlH0ETyk5o2jpb6kX1/f2I0yc1282ZUhoIIuuljQI+hBzuV+po31GtZF9
S9/B5oyoVPcdgBgrYoJbL+effx9qbcCsBZdgrtZLvUpJM4LRKaVbGexegIS5pqQ8
WHQGpNSJ1WuI+bl69LscTpZcVsjPM685jfAqJBAVkv2c6U1i4pPVBEhl/vijkiGs
5AQM1FBgod2PvZ7Y73rIapnvoMVWXbqWENb6iH0h2hj0noWNXUbrQA7P/jZYfrCd
DQ7eamKfZ5qGEzk6vfNVRC3/0fHRk37u0CseD+uAU30qKZ9M2T4yXLsfxsdXKGbp
+0dhLropajPOAEkg5iZ31aWzqKbK/qpfvth8xQSuYwtql+F621Tx/ebsv3M+tr5u
A5thDt2MHn1IqlkqO2nlEgP1gvnZNEwtrHLvudxaxFkxYevpIzaPT+SP1i6JVjKD
bTuSyAHHl1csHCGyz0LsMi40GiAgp7F1ntP8gBf4GMYS1Hv8ghrX1MqwXhE0OB9N
ReP6pLv5QWs6TPjGe4omyOCTnz2N3AXfPi3vDgZ6+nSSlZLvhJ5CDxClWdQHbiLW
0A5uDpICbYA41Ve8KabuvvCGvhO3LSbMaNZz7pWF+e3ExNomf7yYWi8vVb/aPBda
7NgnXEVbtR5w5G9ztom74cn1ILbk6j1nk0Mh664AW3w+ODJ1veLVPAYG+PLP0Pfx
uM++9KVpRK0a3I8JM7oxJPF+2WHYulEBOqhteXP9mddaW+TmeCf+X5UXVF4Zo8nY
NXqjuad7FC74xZRRsYar0rr0Sio19+E+g8Lv51Ri16I+/HUuYF9BOpH+g19Vr7jB
9LiiW7qSU7wtcP5kRyc8bGVLDmiWQBA5hHwq4d9SaRVUeGkRdJ3ew2KbfQ8wjc8I
xwnj7fb+BgzoykH40F6n0fIgshi8OPCdT6cObRLhB+URLd9nXqSQUiJ88hvF5yn5
jYtklibzhuF8mefOXhdedS35XB9CmIeFARMkPPp2OA+lPGmgG03YQkhqzxWA8c2F
r3+WekoIL2WzeRhs4ljzyHragJecXGncnkM+8Vg669TqDD0IhhbIQbfqaaUDowZe
aWQhCFsyuz32CnvfAUcJzS4xSI3wKv30C/pPCkp5PExt2bTiSlcLbxdb8yiCqRfI
F1fhj2Rjy9Azx3ZUVYAJBYxKPo1jtZk6/jYPuszyMikrs/8abYXsqWEPKgPCUhiW
ErcZFeZdbWi8fXdR+v0eyxV4sVYFneZisQJ+gLOgQvf8vuAnCBj0SuH/m7lIx7Kr
l+T7sqMTTtZi7RrMw6z2MzEe8nQj5U0oRjd+AqmQPIkl9j0N4z2p7k4ujGw57Iwg
m/LF7ZNkatPa7jAWY/3mSn7d9HVJNYJlZulOk2NYBjNxQqAwU88pVhxyMZ5o5AAv
N11Po7H762SdoDFMppBwgBgFCQX56vfSWk8laZUzpZK+SJqFuetGoNpuFUU0RCNL
4TZx8utMgaoIuitVh+zLFz3tJUeIu5lJSD3fIksAiuOOVR+tpUfJqThZjVZNQ/YC
0C4YxvRBgU4Mnr3RGjGqowWpKbZQsXOGpu4eJlHBw19moXJQvc9Ch4UcoKaz6Y3N
LcSXMepM79zvTc5QtaINxC50ku2XX/sVXId5S+BlyRDThzlu1zIMZEmlB408J9mO
o8EPUvXT567DFH5B/apUmHsr8pgqY6IJ7wBXxkY4tGURuJkiu7WfrAtcsVIaVMh0
dQr/OQ1GC8LQMi5i5BUzQFaL0gN5+7Ybo2FvrjqT0cYnJ3C72wo1SUXK4WY4y4x4
L7YYGLuQ9VS70MHIVnsL2AGpWN7LAsyPsFfAJbmWaqe4jBwwK44LR+xeMOJYPwoW
07JCJqXpOHOr3697tBmv7/AtJz8aHxhqYe2NsryReVsawP0Bm+LZvkpq2PDvD23C
lun+ln3+tiU+oqBTWo14g6vdzzaGsYakkcKEVNjFeJ+sJQ+ykHTMY1qDGveJY246
I1FcNFSirqfuXvcZUMrlN4U4LbzMYO+lVOGysWcNJ0g+s+JtKgmKMFTR/qP0MFKo
r8uvtEc4IP8rQm1T6WgqDQiaTJO6iDfu4ghWh1dMR6dSSgGqr9zto8Kki0AZttkV
8mw0qpXjGyfAK9KVDwQ/1b8fqStKsohta6C6fcmQQQj1RmbZWskTADPP/PG7tEy7
LB2VzVaz3ZGbxp+xalIn7RzkDjQ+/04zX8u0HVRE10peptx2uVYhzbXkr8/dJ8pi
4Cp2Js+UkThadIHj2AUp64CYtTuO3mArTVWE/muzOHsWY8imLN7nb/PD55oHz+0f
uyNxqoy+TtT0PRfAx66lyRrT5Djgc9ArKF/HN6HXWpMyVZk5CX6QvXhOeWzC9+S9
VeVEpsA5eWDIxs9RXAxwM44LM5o2b18aYqj4hnLOQ2fTtx9HbgR7E4ec4l/AALue
6jnMjVvEGIQSs00sVV3KWqxJ6ubls2U8zBJA5aaZmeDNfovnKxSZoZNQtfPKoRHV
5le2mfbCsTK4vdCAKEITqYK++vlkssMSaAh4FUYZ2FqqHGSDDHDZEor9BEVxuIgd
i3jZ4DIgfR6DwaaEFbNbUZ6f+iNC5CQ2befAp4asgWi723V4lrsLhFfetGcTm0N+
UtNs9r5p+cFlDM0KhPZ2+MVjcZOFzJkNPqeK0SmWm7/x3r0ojxhB4IYlujUSIop5
bnP4vteI3HNVEjUH0WLQMjGnWq8rUp7zw1tEJF1DEyqMWy5Bes0abXQuWV1L1jXa
RUtKS1IqGXhojCRta54uImHSo1Hl1tbOdOzigfENoLME5buUgUzyMx6F6pLpshVJ
tIyQwKc37S3UzaK7+z+IVEq8krw3uP571+5J9mBzD4LCHStn4dTEwiNddFKSW1FF
K0tG4x2rfWTlQHSnmaGDKdmkm7nCmJp2J5pR6d6uP23PpnQlcfEDUR4itB0/HuaP
UhKwN/Eio5DMlTHX+J2iJ2HjT9iq15DushdCtX0Sp9F8l7/7+IQKkApXgqEUYm/h
yvazr4hFtFiHyQ/AjyBB5kRV5mBz6nFYcQQc2pdjxmUFpusXTAxIm3bJeaCuwpQ1
7KNqH+XdWfftBK5G53R11J3k0954hOkGZP69MP4Mv2M7JfFiB4BV9ean/gC467JS
+mTFwexOUGaasFTBmVRYxvblt9Ool6YELbmvDsQpstoSo8FsOXetpD3fJBroQrIu
RPSxJ4Hx2ThHuFZgEFYklNvagdq/siT+l21b/9OXeVHfLjyAMMX5UnoFLGfnY296
zxuEVJDYnO9KuPcdJY002pRn0AJg9rW1d02rF1JAh9QxFsIKpx09AZSkKh5NVZqP
RFT3bHOsAKzYlwF/cSmghY768aA1sszG6VN/ZpSR7ze7a7WSt3Ik04tuTPyAS45m
VB9bxmiFvO2FzLfGitU6yYLcrAZiSP0suOiIJxPcd3WXZSij0BgjznwcC7/8m1js
IGSdylSM3LTY9BkwbjdSzQYGmxVe+9S6RuXzrY70Pb3UxqKH/HbM5qUULQb6+nfh
3sXRQzeW5n3e/e28eucj/l1DF3MatyTL3vWVli2kte6spFM6auDtKIMNIkd9nlXp
YLLrxe21R/0pmaitzrrs2Y1m4hZyntmkpbQ6ZJAkKx5WFxx96+EEcsdv0MXBeJD7
ERI7W70572770xOVzGMNgDKxFasjhvJRtx1P8e3NdLa6aoYO6SrwA19iMh1vW87S
MM6G1kGdyidaGXUsviWkhQCPQgLSyisyz6joLvwEJ7CL/TxlOfrGXLMNdkWXvgH6
opIdJittGJGJJ5vgllTPFUcP/hIwE5IdaAqPWaBRZDYhvx0BpV8TYy4Gk6EOrBhf
eiEgDXrOrL3kz4w/DRELYwohejGfZSVrgJFUDaWM6ychWxYzHmq4JwCfyO1r98YT
UcI0Gynxj+JTLzbJpyu4EMpkcO6yt+49YUXKixd++AmlSeW7pQCUX2sc8ZA0QBPO
CBhXCKg7eUO79A4Gmi2FUr6nnGrm38oSQ97Hvu+QlANE2V7tF8U2ESudF7JIFdfI
2sjydL5pb6i24R2TUhjHhSCtJcHE76vbi5D269N62ZOSI8/z6iE885xdC+VIVnV1
MHyPKu9oGgZxoV/X1+S5XQ8y5HO4Beot8mRsXwEZLUOFFZfAhsaw6hmm5gMvtrjM
Xm/TBiS11MmkTkhDnSNARzBYjIo2ftyOq9u1O1gO9u0AHw687F4L5j+1tgSH3f2m
2vbmBRgXdiabEtV/AXya8NPKPUV46Kpz0u1eb677IFmvzKia8qTlT4FCLqmwd4tz
TE2147rj87hzwqBl28rBEQnvpx0VMuCIYezIKqVQGEOWLeBwWTxxpztdSVEzpn5D
Ad71zhjzWSKRjS2NI2tb47Fa/U5gkmsjJKqZvbh8hPqVzxmKSbgC82fFz+7TTF29
1s0EtweE4xnxiRqOupjgVSTwdLP/wBpWTVL2AlZ4N4rb5IqZzIG9R1iwVjMSg4io
uKsu7oTAGrbMLXrwtnvGHxtpySmNoX/MxETKnNvQptux08M99B0oJvCKxZ6dU7dV
1F1ND59k0qk12wney8obLd/7lE7Iga+iQ9Ad5gZgqqM2HPTXN9QETPG7Jb2rL2vn
dGpErd43CenGhzLHfCMesSzIe/wwEmNLdC3W3O9JeK7zejxoeOJnXg7Z63XBy6A6
OXIWDGcNhvmopShPUCl0IChAoNenSbF+brQe/IqL5tdZdImA3ly+w+UWkwkbJZkx
2WpviZUBhQQEpB3TluFlRLdHugguzFS8A8gbINbxI0ZeW3QH+KELH8OIb3oUg7pV
t1yQPohtG6heBsjS6kNi/+8btMUmpBlNguApmD/dhKXhAPUlGkSCQgiSFiZEk+rE
ccEAOhItilDJjoXeaJYLMyCLDwDtNLNUI6CBtUJ4cW//A4vcBCgfY+SI6VQp5mKq
sG17ib9MJmTeqNIwLiN8PlFhJu5xsg6uKGqf+TsM3olBMl7uJMjMLrGtvxTmcFQ+
QbQmDeY1iraRkSrPj16Pko46e32/U2dOnSC1wNXJMw5vJXXzOxZdbue5QJLi0wBw
ya64GG8waZAjPiXHz0O+3COe10DW5WYyzmZ5S14/qI7eW4JbPCndUOKm5La1Kliz
tRYId6ca7nkOgwZGz4f7LeHX3KV8SKf0kzcLITrwdVsaTDtGXuL93Dwbvp+N+jX9
Hvle57/rxp7Gl3eOiM3HrQ52m0i6QQoLyhD1X1LU7tGtqmrqpP+VSBt81E2coQkW
nzMXVSIg+SW95Cg5NIdSgU453OKatsbonnQr91Qf5ocLZvFyHVVALLn5uabWLOVl
j5mQ1rU8a3YbgctUyP9HCnsKmhkhTSF99vjah6V4cxTyTQwK+ljEGDnNSI1e63yj
M1ndFNQvQ1ioIi5X5cCw7ghj8uu1kajPlaemY+UOLJSxTYCrY3xO+ziKSDehx7QX
TTwvXlMN67/mvzAJZVCAkyTz2mWQbtBd4YAfQHgubYgSnrzzqJsqBEcfBoRF12uY
XoBKhg7Z5Jfpxb6J1311o8xZ9LpRVP00LNyKIDATF1Yoedc4YJ3p/vVp5b89eYvU
nziALsznMcY+RM9YBXQZeBcJU0XftUbDrS7AT6kKEI636iQpwiXAKGKKDeo8AOQS
eOiscE/0y0LsiYgNZl9m5txHnqMU7ndEtNQDqFRwBxWJBztWwsHi57AcqTumLoEp
YvO5WGMmZCTYH0E7E6vQT+bXpaT7UJkaLpqx6C2jytxwqrryzaTPNka22ZCnQRsg
k/w8KkM4U9Elzeg/2FGn3aztS/mh+7KeW329lIcQx70SERJ9qjKnv4hy/79vzzoW
hH5DQJoFqY8ooUg/yZdeM9TeVkJIP3OCeKsKBoHS7+QE1PJnOkKsR5bCL7LwVmgc
quQbSBenhKPxoiQ81nVmGRnePVVWT8+U1StGUaMhG5cz1aclsY5ox7SZQsGC1Xhq
tk8PDqWI6rNnzT4XwMAuhTLt+3tc7cIVQvkJswX8R8vGPyf7OBS0TRt8bFLX+3fU
pLWJWNSvQ0qRgb6efMKPBTKGnWzo5fOA6tPCIgKzVMHwWvgpfGV/eF8rJlEpfvoI
EOMlCoUD7e7qTsEpWpvC8Xwzvl5pa6XbUldajWxoCW3MtQn7YL3ppLSHbkRC3Y7R
IFP55QhzVJQXTZWnYXTqPsWE+Cu1HyFzjjLD9K9zEVrCDFcH5oPVDlMQzsbVaF3J
Mh0tUyTrp+HR3/ye81JxL50Nh5p+kmPicJaA+4L9z76X/PBbka5rnKwBGEsL57Lr
wua00+/88G/nZh+U1W3WXEeXzws6Uaczonb7SfO1UxlAnL2S/ghXKxTUvTbA6MZt
t3NaXgfzf3rYxWU4mR2pfb4ewfdar22by5Qa9TAEi347IEyKgVEKuq78Dmo+Y23V
YZvGtzxxuLlc5hcW6rh9Egw/uKjQGsJoCDOx8Q5amI2b0xKmNWF29yO5qhETaNwA
Ckw1hBaalKArh7YxbBtaisw/9kPTlyBi+YsuSBrLWyCEBGgEz9266/wKnKI+Z6ct
D/HKggeLELBWS1V5WuEIVfjHZbjhktkuPq4bzlO1FhMFzAGfFRnLduhBXP42GUL1
m8b4ul3D65HvOGSwyH0PhN4SDXnPOOudT6l5aeoQuAeTWYehLpP7pWPXFY2q0QHV
8j9EuoSaWXda0ixOZkQAunLm325DEikD9h03E5rISuVHh99j8eUgUoRswgjINysr
VUmCiPtmNlwWoIIFCr92Z3QxGEu9rLNRLlArT3JOkeGwApqiXeNILQVhBlcQqRvf
SKU1cduKvV6rC3yO7/Yj7rK8i10S7aKpqKbT9lhLJsvZGRCV/J3mZvNW6MSCA1IL
bPIDlbB0lmrqz6egIQgrmc9xdQxFWiZddpOyvTq+xwjXySuKR1roc+HAHb8Qntdi
QiAYL4vvu7JncMgHJe6dFZPQOGbw4swTlZLl+40VaBZGCAjZYLefpAMDjSvEVGRG
1aO2kk/8hNs0SY0kH+5efIZEYKYZg1srMt7ybdC9FHVLio+M+fLmoc3eIGdc4HQY
YiS1+w1k1ZDlY3G9SHI6LmLSQfJH4jjYMwZI6wJ3Ru5kzcKEV1FNGqYtVpGsaYzX
kton67c+YtexO7oIsOCNXVsD74U+v4cK0hnnufTC+rIOVnjOuM7bGgtYh2Cy2bA8
i+3VP5VkvLVFQCcR+X3YNuC4fzfmbq69K4iX1kRD5IUyJ5grjChizyF/B9bdurg9
GNdAvxu+/tznbC+EOH4+Km5JDmIKt4G2VSvkFu4RYL9m20VQOJ+vVRse63+Fq6VT
IsGzNJTfrNRUijriZltrM+IQGyW/5A5ab+b9a2YncyVb1s2zZfakQoh65PFqp77H
wsft0h1ddmP4Xph/7wuVtM755g3rdWSE6NfGuGSZYMsP8VPQiMIxBN3zd+/TiFyE
feJdaVQ9riELl8Hpv13tCLyjI0K4KztC/3Oe/pwC7FcvHa8mSJa/9qSHDF6pBBaZ
SHpIJuChSeLp4OSObp5Kix52ARzyL+FvgLhrkU0674Gdd7eyytjt35YVvYXmWBFX
HDGhFWspqfD5htd0nvanEemRsK+e2lGy3FZdGdCSFDdH0ocmJp5MP3uJfRnYRvam
HZmJwB30XBT6C92+8ucEpYkOve+tb9+4LWokkTZVaWy/r8Fn6e4ROczHfzZA8brE
64Yx0ShytGWyB9dkqclO3j8navI6OTc9M/poSfB5wpLtl3+IEOdrNx48rHoOBo17
yH+xafx6yeHHHv8pJ9xRPUi6MLRAG5YKorw96Qdt5UKr4KNwbqP/9HTIYO1eW4S+
cDGjYas/Jhq47NtJ4SiYJMJMGV/8e5EfvvdyPkFdJ2yPxWPSDFwjXFA2deK4YeKc
7MyeQN/4zhv2wSrLMeNcfG+yhuSVtlS7uXHi+6a1JsgLD1+hXXZ3yIZsgFwcMOYW
eN8J6gkOeY03SYmY1iocaBMZgKAg16/aK2nKaFR2Y8l9LTSs2ou4vJFJlC/wJSW0
6C73IBl4L6LI8cI7NkqWGjYYjX3tkvsw3DAwSNFHMrZixJJJpZQ0XS6RJfdZDs6a
cI+cwP4jNqoxy60jdVo6FFElWTv6VDGb9ZI0PafwwJshq8L78OApU/UDZQqQlJ7Z
V+nkttyy+Nx1AEtD+k8u+vDCDTDesZD4lXoOSWXCQH5DWWbjYl6858jTYHJYB28S
M5z599vuaURnG8I7A/vXu/4rNQuZUQ3xW/1Y9PKUfilzsCTaSfQs4KjSmVBk2Pom
wPu2FQapMyNeb+E9erPDmKtdGJ8+Cx8x2YVpqJh1CgmHMN22otFfya39N+9o6ain
uwKfaj6TMQlRepaVA7GIxcjnztCiPdherfYMH7xzYkuRsAyfnTx/jw9aGmzQfVB9
JczklmgVHSMH2S143JP8WHi8Ed9dywReGzpA1tM0aA35VCLCYunupNUrTSQAma0J
kQ6ry6/jxbBGA/d8fs9J+812c0YjnOI1qFU44rl0hVRtMiiikrLODlEGAtOEtJff
YT6QDtSGEF0dJd3gqV/EeDOdjBjeT7jejs7/v2DGhYOpzA6kHHSioThA7pLQQvC5
Bwdy5VgST+BXLQllxZBXFhWOIeebQfyKWRd3f8ppXaIADpWo9MfLXKW/b6xBygKZ
AuknsGGudJcpDULyfDucEpJKXvikjAZq9PNfMHf9wYPj0Z5bo8WwYZStCY4XuLzS
GET0AnCcF4WM2QlaAXaIbnrDiB+/C1ajXl7K8Z/44pFGgA8HmTh/LpwYWdgaPEy1
mFhtrWoZ6ngsgsuSLnpBjyk8znxLBZOil7IYVsxVZq6nFc/TCwtekyzeEKPst87z
OlwMPnS+qG7SiDCNkGXPBFsaok0jg1ze0/BSms7mIIMwOyr9HFjpYQ6236WWwdoN
CllVNMnuo6bFX3QJGpOZqI2ZAitmjaQa+SOjvDFOJXwgjD3Bt2g/R0c27apbA0DE
pM/SKLQ0aC++IPmeZ5O6sAZ1LTtPyZ0yzMpIXam8+cXtmjW9Gx35auB+GRM4Mdb8
5YuH3G2aGbktPIr7i5aVFLrkiLsyXCcCo3N5koeYWGO9HrR2E5fKzM5y/+BVcJMt
IZ+WtLxPXyEvisIW1usokVSmq/LcKhWZ6C2o2xPgp3YOFVIy0tRnOYe/iTuFFkP8
roRRS6obcHWy2W/uKuQM1qoxlT+RmKIKgnItrA9GuGxrf4URN3mo7iPuS7qsm1V0
1yyaAwOF02f0mHSQH3rQRKoT7V6Aj7jo+fYR756dkSbvfY9WfBPGNg6/j9jxEvDc
oME7oDIiE/2fhQx9fWk99IR9+u2UhdZ2f40GyaGeazSGwDC1ir4d/D8yYVUhngvV
BlYSydXOU6POInqSqvP6z3xz3581si+2cahE8wno20viWT4x/Pp9Pfl7UZj8v1TY
2WjlpzrkNkSrQm0FJfpwu3JvN7WHf8jSP8D5OzJjBPXeNxykHFPnL7fLL/ilpoXl
6AoW3zc2s3JHIj1PAqIC8fSRuStMaPa++voglQoVbUCUJQK8M2CBzWIAz5jNlkrX
G2gBFNuFUOoxPzaCAhHx6XVKlU9a1onHZvlIc3J/a4JRgXSior9iJ1jpRJqs/EkA
Ht2HKZwEHtbqwY5oK4d5uGhxXJr2KE+hikZ2Sg372K1303JBkaxfs8E1GVQuwCBo
Y+yD/oNZKqtupnOiqpGpxo1+1oUkrpF/xZzOaagXGYepRHT22YX5yMck9+z1R9P5
uaoHX0+xBOkRZRV1b4I5pHxs7q+3YRzctB3bMEre5HSAGVbaWH4M+lOR6qXM06tz
YUUjUkL0rKNWgxpx+fjj3+IIAkir7vQVI2Y0ZF7nHtYh37ZIjTyfgAl52s/RlZvZ
t1E37ZLiUUhiQQlKEoivj5D6mGVRzhaArsbMF60LYxuczRAJ4EQBEOJY5PkxnZ+E
6qNgbfYUWo3u39TXfCx8UoMlpD5cOR3ZeN+qIwZ8ynKWENkIU/l9VUKR5uvLF+Jh
LYoSBbRj98kCQEJYmymgc1VpnXHAOOyYrj6N9tauQmMe6uVSA6FLrLfM3MlRyxKO
rhPpOUONuBLKHNUD9BNQXTAwhfUKIZhmdcBp2OSv/UKLVyQniC5vWddkg9qAgAFR
Fvn6n3yNMaCqbaAioszW+GzBEPaSZ2E3vxqoKk8nVT8suID3XzQGPsW+N67keu8A
j7eo/s9uOafdSD4I7lHh7JHT6w5MoNq+MDyzIZCTzhCm9C/7cXi1E8UtXm8A52Yn
Bhhd8BKktnQqvqGnN2zLabZdysoHNVZzzz2mIGBAuee8k8FaMJUbdN7kQqBNHC92
roQHaCmDzuHeZi/avXLEtlePQk2979baEPadNyrDGgrE77sFat0aI4B/xRG+ztYB
boe5Lz1A2/0xAbI+r3bjqd6PCD1rTpAvAiDy2FU9reJzBj0fyobmY0GZgt8syn+9
D3e5NSpPu8VcjxAbSIk5Xpn4gu1JktQBx80N7gkvNbnfYk245s+NG4tsfr1iF1sB
ZKqaPuGzwKs5pj30Za85lmNQ/aM8tiEApLaCYdHLuEM5FryfiYC47iDT72RJRnfy
m4kNYjhEOniRH8fqzsdX3osmvrJZgHrPxroecF2ZwybTqISprhHm0D4PmO40ohbM
nfZYVvnpHiMV4KbimTav2jiI9PE7D1owSOeWKIoNw9Ajd+AcstUmj+AlugpnhnY/
y73BXfUrcmojLfpIVtRxssRb7YCTx0Jse/pxBNV/4BeeVbnCZGWjAO4mSCUUfPcM
7tepT9TLswhkyn0l6gnejHczPBMmvS01QhHWgMScv49RtrS1JFjXkYjxNvdRdTIt
HyS7I/9DTN2/wQn90fdsPgKTuFr/vWkOOxgXwKtbt0Pps1EJLsITlvNIJv7jC6ff
aPSpLj5AaluGpRQaZyfrearS5/Acrhk7wzgj3cwiFXsh590IBt3Wd1A6/IRGaKCl
DRtXjG2nnG9lwjm1TnQrr9FS5Cs6W583Olo+sc/j2GIh85DDhA6t+/r6wGF75QgC
dI8h6SwmPacXj6yG4AYoaFnq/l5Mv7pM1eGGuZXc8n3EOQfD/38tB/UxZQXbyTjG
esdksXw/tk9yjrnJRXCwDTAmDmJ6rDP4Tcd/Z0PrmjBkvt+U4W44pdEC5NUhnA7X
UFymogB3BQvy7sTOjm8lwccv5KqRW0j/gKCmpAJHZqry9sYg6FvCuJuLAfmSOsHF
QUM2t5+M2SqVCoclpTdH2V/q2UFzrurEjEhyL3RXNkdSZLlC6+alVohYm2yq6gxC
Pmmqdsj8wUNITmbnMLUgPgTy6Nxpz4Mxczpx9le8w9VK8iOxrA2CdqmNEXBpuk2G
8iFFL17O2TJwAubs3b9T+nnyGpajDNw9/o3fgEnnSKPhqEyPiZ8Sd+UZmhHY2SlH
l8Afv6pX+86Tzb4beecO9w0pCL8K1xEZMhIigFaFgcjGQ+aFYnZtMFgwzCrDoiyJ
6jM/kKQHGPLSldhbvPugietY0SucN4iRcs1ltfXKKXxHVGqU7OLFIBtK7vdVoVws
kGutVp7KV8yK2rQVqbiDItwVBt2cr9sLbOP0XsWYPy+Cno2Qh1PSljMCWSVGVAJ2
/MImeU1rFqQma4a271V5+WnzDnfN0MEYPcgRriAdnwgM0/tqjxY7RTUCtZaFkq5Q
JqqEXKt9Wx8lwEvk34yKSNG1560ALv2fT2a2r/K6EZRasZfDTDMI3jt9o6P7Lyei
iAx5IMOUvrunmy3u+8AmOrISND5WZyQwhd3VaJJJ/qUAmlGA7BT3FBLMlF881uVL
0cpD8JfhadlGm+/k7BzlDder4RiRMQ3lc+t5++lkCgGpX1L3j+lx5AlcbmMbmqE1
BpnUo5vlDkOUis/AA5VR/KFxMYan4crpIistUeVhMqeZLay15V24jG7oq8ce/OBf
gDTFTQs28HiLsyV2dGcRSbDnf2con3niVomZBHxvIIsJk10WEdZdk5Bint5x/E70
2oNwPXAsr2jck/DPWDNqSUb3CEzh+o8TlB4qlx7dAimGUMLTfTwu3Y6qa1w8WlWc
TYlQ9TvQc6nAY3r5H0L7q3NZ2GND6LbdTVWFD4fOX5fSQco9z08i6SvTANin+iYz
TZDbLWHytsjxch7iYb+7vONOJv9Cf9HiCZql1LSpkAcTPgqgeFwYeoAgODUYSM51
UbuCyGEfSaOIExkTwURob6eu2avvBK5A4s7oYthkivl0erxaB63LpFugC2t0F/MG
vzi022llMtAaqR5aTHYvzo4jBUE5rip5qL09wVAF1219QTbFt5Ov1OTYl0YyWzpL
awar8rzcYTjcs6yC/XggYscGXnIxOa9iO6XnvNus+Ake5lMdjmoQX2rm2uNAyClH
XP9VoaJOZqRokAnkPcY+25P92RBC8f9QmMKlFurHRoukHk9HynXwIaLrkt2cjU37
jSroV0HXAXyjx38jv3nQR9kvxUi2RQgr6OM3SSKabfDgOvdFsbeO0ubJ11jkRI8p
Vv7EWpiAAVDRNqtjecXiUKV+F+5NjlUWl1cDdTuT9Tf4mLiTysuXx5AJ4LniN1WU
kpnMZ/T7pj11g50TGl3z60k3V+7FFLzDNLJMXwG8EZoXdVruycVihawhNuy70dQk
7f0tdircKyHCaUvXc5z0+8qyrgFlUjw0DC4qzp6QbDHlVs11yNzNa+rHoyiS0nb4
JWuoyD9KpS0+wpaXsuF3Gdsi5kClCAKlGnJd8bGxutSfY7CWYPsqJ1Wo2gbkyh6l
4E5TaXuTtuS63MvyOcz+MslxckrGM/E2hdAMDUqlJtFW6iJ7nB4MWwcLrzilHt8T
ikaHqlUtWpNKdIKX+0JfK6v2NpvO5pQMJ/dJI0FTozEOtgt9NWjyLF2JVHLIPrCQ
1/mWzjJrst5Gvt9wmZxfi0KiR8aJyQG1lP0yqLJLix1lV0+b1T4nnLitcl6uWdM4
E67DTjX3iyHmTPXIGMVE+34bwocUdqu8gyp8rfy/uP6OoiP9yU3yOgqaGGQ1Mcc0
dlzvO63zj/WKs5un52I5GDqLE9Z3IFNQgGQ/wXVkdKdELOS5GtT9uhvVcmv/q4+M
Cs+nDgwWjtZ7pe5g3TpEnlZJQwKFrzCxGETR3Zp/dqmqeQzOkr1hafcK4UMic7mE
qcw5uYfjMMCP6EwQbeOiD3NTlILa0A3fi6ID3SFcFMWQHoHLiR+0mCwrj5NSgF51
qCgRmApAiLhwlPaoDl5x5uaqxWLiwtYs+blCCuQ18AyD725EnX9AzuzQHeix1x0E
rewkidZ9jCcfUrprwR72OzQVRn2SrLMccSp/udTXv4el8IF44wqG8pPI1MdNAohP
fAG11LqMrGkqX2TylnjUCRBXbDNxuv+D8crs2c4XWcmyV4PbzTaguI6nAvSNSRLe
EEZKsD8mHaRMY6QMSujhlP9FqdMlhWbhU58lxUudgkfzq6vm1ePQDJURMqD/Mx8q
FTfIduJKHeFdAFkf3zDPOc9fLA4b7EqcrBt8gZ/0fmlUPUmIzTBH42JeoBuOPFIb
mGwKYd9l2DthPekIRa/v33xEjzYpGWebMe7F6YG/o/44UOsNRlOF/N9JSz/quhg5
HBKQspZeAmJGPYoK5dScuWjKpwhK6EOyeAA8mrYPBUTlJoZKQ4ar1GKXfkmgeplT
5klYmJcrvDcegzMhRVl+SBPeZzIa4DfzqSXk/nLB3AaBK21EY8VZm3q6LER9+mU1
omL+nbwMIefMCeDMe5Zl5LmpEVyoqj2X4dERpyvqcX5yifAgsMSpC5FFWFsIk9qT
jC73gHzeCtkOcj4pS6j40lOgxu5MThrcbveLGAoMEAWC1KcLFk3QZuhZ3grkfRyU
qca6d2nN8uQ+aOzba3yjktIKYCgH78tsoFX4TtmEWP4FUWvKje5+Ta2p4INa/yE1
JNLBnscyD9gc2pDTiQH56UR1isV6WyyBZInuAL/3HapvG6qKtqq1HUQx6BoGE+Nh
OYO9seekAemJ+WwkyV8o4V4QvDc0/ReF/AEYZItFEJJ6QCk+QsEhi5SJYeusV90T
d89HqsHSdQAfAw1wQLFLLyjhRKj2AoayxN/QXYuYW+S0ZeHHJTNlyEKi/3Et6lw/
OuGpaFxRPRLMjyvUA0esGsKNPrPgvn4Xfm+HQlDVE0KenxfUhA0yrPDMUbX5x9fB
nF0n3G/3gKJ771gCX49lpJjDxj59eyOlmBsGh6rln+pPb6mCzXUETLs8+5kKhmYX
9Xhls54GVT8u4ibRXnMZjUc8GZygd0tXOLCE7waGYpzDAY8m/i2iQDRJ5t0BAqJv
xR2a2ih+RyBVXZAmvcRt+Bct62cJ3X6y9/fqNB1hr8Vr+8xybajcq4MkG6O6TycD
gYoG9V+WAPfRMQpZN1Wf+61N0PQfp6xVT9S4+I6Cy7Wis4ltLBuhwc0umd+e++oz
PQp3kOQJFI/mzw+Webl7Lo1HetZVPMpQpb9Rd8gi6BrRByaW/XXQYTVTtkY/MNoO
BeYTbHPEtSlSU92THwbr70L1UkTa17N51HROYaM8I4NFl7P5W7oYiaO6YS3edo5k
QJnNQNdJW+Uu67dt80LG7f4kwmyHCFnDmvPPIfzROmRrwjGyS0wD04R73z+fKx+j
s/IA4UDW8wWvKfZzBkK4MfrbKO4nLV7uT4NP1QJw62KMRezv2Gd+qLgkHakcexhT
zSj3QVB4GD3wjhg7Z2Ijvq3NoZJlHfvHmYQIx3MZukJ2pHyHfslwKCITMyB2rBH3
+zj1FUJG4Xa0MSizjMafW7wYX6dZMFjpThhxX3S8QJcCaLEJqkZKyw5oWVOPnUyV
1NXIWpd4MGfs4WAT/U786AMVqagcv+cRxLbUi0MmpwVZrjcpSqUcMoQ02YywlzN3
+2PE1POvZ5wiUbLzEWmRK0ZXXPXczeHYtff+Om8T1+sMgNPs3IlUNgv1Gkt5Y0xY
P8nntwEAVcSxOHWzl6D9hl+p2veo+6KrS6GuoM1ZLZYJOXHHN64W7guu2t7l/ijd
Vd0X4RURRI/w4c6ya9kM2K5MecfRfz7e83ICtZ/JOPINWmYSFK0HPBhxorufQ/SZ
VhDOigYEX8oHWhJlxo1aqJMqjPQcBCpl36YCTg/ocp20KDHpLDhrK/7zelh8buG0
AKEH3783Lk93U/xGoAXjPRc8bj6tGYWFjYEXp6zqFLwFDJy4/0dR8bUVWDSs42Ni
93oN2U2pEsfKUoDt2hpCfvJV21xPHUdvHxCMkzQHtp7/EfYgUXkshGs47vnPGUUs
J4BSHBdd9wla8G2md8dhGQkBv5rm2I1zkuIygJnfjRQRg+mE279cFD8GDl+qPElx
8TvrUBfvq808ESjWdub9y1sYfqJPsZEiViMSxktgpHe9LJd/ebw+jYxqD5SkuspT
GQ5V8ihpoQeAF9mMmcLm7nEhb4jJv6BQJaZgHH3k2J0AD4si0EGoaoMlC6HswEO9
M4a0VPWEPslhuzB7YvrJ6ZHmrhp5DlFZ8h9bMp6JojZ/jQfDcw4kFaF6C21v+roB
XnmyGJ0xxdhpgpJpavsZRDp8/owqpmNKSFFZD07Pa6F1CRX7Tyibs0r8xszzzJZU
xgmRpSE4g+Z8ZtmSanTqOyThsh3mApbPOGYK88nW/TDppmuVBYJrE/F68sAuNY6d
aJW32o3qODysTnvCAikvsdSj/3GXtzoOzn8xCbvn60/LPVcdC+tp6Lc2D2gfEVFr
pX9wRcryDbLeGd1MoiLvDwXELA75ay4JuzR4iEtA8dTk9VnXCCNcp6JNcBSMBWOz
JxRuFxicqBv3koxnEhoYvJF6c6up5srpvcfF2xbLZSwi5NB1xfdo0f73J8r3xCL2
+z0r9Lzzapehlcbf2lSMRHJNvvIE9zVrqT5pJb6l2SevC4lYGrnKvMNybkrkSXjf
5TYGIOimvDr3d0otWHm+51C87VmVsfEVd3x0WiOhpSRtHi3U/B6R4HzAXhReCk/3
hrl+fixbqKr1qrKdhoZ8GOeh1tYC/7gzitgDUWOYbjGdJgu64wiohqvjA0uMqQXL
jSgEE9kesZZH56QUB/QqxH21buBu7SGS074ann+b6WiXcyPe81Q4tbSaMTP0xNGV
EZbepM6WL9imRjnYxNhPUakvVoR6seaGJDVX3jJnwRu1R1KOpIJ5EagnrwVsTDed
5lDNDNsSy7/+pX3urFVu+TT0Awq5/tRsfVMImSa5mKEAgGMnEnxMdv27dECs8vY5
NUad5OKqdKr4SlEB0A9whhwaPWe5OXCTHP0fiZjqGd2B+4sSoayOkc4i4DFrLPG6
CmvftYtdj0x3159zMWkdoMvx/8rMfeRf1VOm2VvByMVLCCFC4XWb7TykCBbKVGlR
pgM1BBIFXiM7CQ5+fFuLpoD7PsKkwOcet7SD8BUs8V90XqxNNb85zVgIgIt+laih
0fBoJ9lSYspBDdUg0mpnmPnM0iVqH4JLZMXmE4cv6/PMbpnUuffK5xJyqzcShjUE
XycKiTCLOnC9D62rqJ0QmNTnc/5fzLvlc6Z7gnJ5nzvBYaBctZ9OztjpmyG7CvpD
UeL+/dYmo7ozY4mZPtPInLZj+hRwb1hlpE/we26OIe3N3m0WigCx0ysn1sGirt+T
u4sxXTZZlXZYXu0uRqPhxbanvRdlP4w3KqeBoRYGdx4HVI4bKA38C5xA+/u5nD0T
19x4uo+obu8kGwseo5oG6LIfUwgFqL3gCq1VkaWTToElfa6vAqF5JStB08jnMy/O
jKD3UpwqWPjXBqtEw0TyvtBGeiyqAKtYrpFw4B3uG6P9HujlyjFfLKghbfvuOAOb
bYK6XwzY9RaP2TGKDIB49PLdvDQZ9LIstKcJONAwfGUNvO7KWhVIGG/JlcZ2BtfY
6uTyeVzuWtJeA1iB9Le+Yn+iM7eFTLA2AdE/zlPzFA2OA6/EwnTiS5lwm3vNi6sU
K392XnzXSNRe+yFOPka/kpsoB3HcVwLcMk/1r65x2rSU9XegJ1+a78taCu/TbIAU
Va3VLxiuJdPISiziOUb/8LhzrdOR9poJaELu1pV7cE8pQTVWyhUmZ10YVGqTe41/
LTzSCQ+z6FCNiaMPqoYKNcb3/S2wVuCZYveWzmASYBGL8fTxF+sZhKyFZNHgE4Uz
2VTQfuEOzCeyapNCvaVp89FWycdUwehjyn1LW+Vfz2ogeMRTmctDyTSnehOfuau4
Z+uzNJ025bbDE3Tarn35SC1XKd+qer6s0wlMbLdKgj05VsjWx100O/RbQlxUVkPJ
iulH+jmpHMu8d5lXROrh3GlhCd7y0Jfgdv1mgMLmGXL1xjIzwRUuNZBVRQ/nsbxb
zPkCKTtHhjP74i+b8PiLc2+Zl3xCyR/acAWHdN4mTRHY1fHfwhyzQY+L6deSoPHB
FD6G94hJQljYKjD2mb/urTLS7moB1cdRIxAj6r+q7X5Lhsh8Chl3x5X/nclQlRjo
xxP5UhZz1dgtZvczg5pHhn/M4aO9BIi6lavt2JycFrnBgM6Gwhp6yQQdyY72Iw6J
Cq/YKxXbmN4zSvd2EAFWeqVgFLx0TExgwuTcId6Lq0N41ETECnqrR4DcG7szQXeh
f/OPajKqgJ+GNiunCj4rAUHwAuvX6uQxO5K9kbOJJlbyqQbQHBGxm531OX052p+8
NGgs6Wowg5eztY4iWSUH4pA96vSKnfZpfKGsl6QDaDrTrUClysSZ7nymXGYa+vk0
ln/24pS0LotDq1UKOsLxWKo7fXDOofygb/DeUHQDggw5W5BAMp+ln8v5EjxRnSvP
1pQRtLlOyX6uetjHRN4xGURrzJR5IBl+Y6G5zfi8bf6UONpFAKCsKExkhR1i0OL/
MTUOaqxyu/xMCU1TeQHuAW1jJMSYjTnFwe0undfrSKRrHodUj5lmIOtHHaHWUj1t
fV2jzSYDh/+aVbJSbbAQ4Sqk2ExPVQ1vu3IYlozX3BU47tdLiHMUsTF1ISHKshhA
NBey1pAfnqw/Aavwp8uW9Ml85EOWOU0FSe627VEOY7xufU0nnBUdTVVfUwzAAO01
r8LRXTYdPiASjwFZoLBDRKD+wtYi4SsTuAYP1eumEO5ma6nH+kUzui/rfmtfxBYS
cT1cH6ASUTTfAvHlsXrAoIG0WsLbRlEP2+y1uobYiY0mZ/KOujGfRjMHj+GCRppY
/azPYWYhWgSro/zQZU5Rpmvo8zH0ijNAkS0ga0Gx8tFEqycUMLsATN62OJo3hrPF
xT90no/OQIZvF7CkBdVzBvSIFWiHVvd7i1qTVJBEMm14ici6ORwocmFi0XmOM6vT
9XuuFDJh7ai8hyO5ywFUL4lRQskNZlgHK0Cdov43e8Mw8pWWaa9zKDG61AluZaSA
ef7DYxx3A0O4Dm5WL1boVQFMbVxw468KhI8HmxfN0UwmC/L0ANM+b5jmPpuH47C8
/HkmGxobMUn8vxg9zQDf+5IYe/W6PXhKQjuy6dG0yZt07VLgqu4q7Z3GhIkeQ2r4
AaCtRVNM47IbN967Z6hUXNv8PcyR5qBsrTAUsn5kJHAYBDOI0S9RIAA7hfXGeBgK
NYqDRAi82AMVEfHuv4ikxdJ+xIC6Z+znBdrX63ZBPKB934QzQNjph92xnFJMZbj5
wc+pI1bpSfuDajcpbaUvv8wZqHo3NaMkgmuLdrxDCTwDTLntAbVOnxFiMyIA1Frz
KVrrTqgLBXvsBwN+shre+6YmtWBtfGT9VJpxlr+CM8W9GJYaRpIukKgtNp+yOhWA
9I4OpZsZ2rayE+8XqAn0eh9tfhPuq6NH6LVI/6wszXhiN1VeQYSC78Ud7rN+yPZV
sLfd0uQkmPGmJdfgC240dCxSgqKm7KOO/FUtDzo82XrCRGOKSw/I2NkBSFjjesUA
7M+Q1Po3+FT8XPZcavIziXO865WJNvWx4xsC1F67VCFr3og/z/JLBACiieIuI8eC
15jjJ0BV6JqNt0VDLvu4pixt5EeMAJ4eLk2lJJuB/P3DtDGx080HSxnEZZ7Vb9gj
WbzdTW+7kHBqH5ajQC5NF274V+0gpXyZRgSusPxEPYkVFLz05m7LmHMZKpfzU6UB
GwlttiNJbU1C2uk/TZJdUe8e+QBprCSRjGrNcpl1r9HHcg5Yqh9F/VHu2OWIlGgl
0qx5kB+6lDpdHKD2NnQJPdXIakmpF27MxmxuADq/AQQxaNI2lNcJiyQ2MzGQbOzg
z+OLxi1Im79/9cHr9s9CoPrsTkiJO+TWFTp4smSIHK2g9+QQbaTXN/XJtuudfdEH
V3sm7Y35wyNraR/P4mzaqfyKu5q72amYtYAbU96ukBArsN9bYqPH3srm4X1y683o
iuzZq/v9LDEkIxB7/9VPUaEM20QJyzm9OWpU7J0XYxkQJGfEudQejJqWXOlVhh1d
E/K/I905QixN1Ja6Hu5BI0RnSRCefUueEJxI2KmRIEElXUAVq0NOsOB/T/LKTzEM
8Yas+9qF2Lr+3Y1ZOz82b2s76sjg64xf6GqUeMFj4jxrb7gsG1TImWbSPuOXYxBV
UHakO9VHguTFQynvBlc4HSbqJK7ZkH6BeH4MwRCAXkIjKSD778mAH7Vyhuvys1ki
+9hPs5RrCspVRhcoRf4CX3YAm20gRVtf+Y9c8fU3pfKbtpTvposPK4jFN/XNltad
pxb6V8X+KF5G1TpUZqv2lF9sbaN7Xf+LfBAJnLrHTryLmtbMkvHgu8TkxYnjBPfw
A0YIswsui5YszejwgGDKSOP/ZVko+Zdi6vMX3Y1e6SJ3nSs8lSl1+QlyRWvXB6Hn
rwuSmLmleOWS68Q9+IWU9ZzemOTfeBrBGIN2sZPyjW3Ku1iCnaUB4vX5BBMZHV+H
GnxpFRT0XWoeqtG1GfyJY5HQOp8jg1hhlwATySujro5ucVLCnTEqsJUmc8HtP5hC
qcQ74mRddccaUZoJeJfVdanM2zeZtMb0bD10tehnHzYEB+FVNsE+0DxJNcXmo88+
oJwqkw7u7SkZH16GWCCl34r84UP9L6A+Qpk3PnddsLgW3MZTXevDWF5tssOed0Yh
R4dHjU+GjljINAOhLBzfiycXDc/VBr+nlsSRwEqm4wUDQ3fNoKvabyMhuzqJ1S8M
zNyKjk1K0yuJjIK36DYNkFB9COpjTXgYGqAkD/hdMBHh+eLlS9GjZCn8zDvFhHWZ
y0STzr2zlTxYg1i81HNdVEIX4jgRIh8ed23I3rHKgVjTXY/qfNjXrcGj4GZqfrR1
6lvkVIfwGHJdK+r/B977xD39nalxJ0DK5UU4zgD8T/T9m4l37s153HtkyrFCtITD
w7VuSZkyevoRuVxTBLPSGFy2YWWT22ndzHoii+Ur8fXwvrUIqYotuSBrggdzt1Uj
C55Dbs8jm+VuzMY4kl1WRSkMD/fgfFnZ6oh3hkvzSDDpVq/3A+nNr5AENJPCxtzc
pvnGdia9R2uk0lheBYu2PO4oP/YdM+7b9MdzCXalvohMoJ6FcRa5TEwZYSg6xEgM
qxxOOcSFgllpted40xrTNwIVkWeEbxu3sOHdcq+kwk/vwKaLXhTYVaoH04H6tpzw
+QuEmSCydQATVyz+3+937DNKvn4jDtCRY0ExB8V8AQQUi+mbCTMSvKlGOhtVxzCj
R4JG9swokBM0V8C9jnGoKXvYZIiH8ApagmjtfxuACnFicvntjDEAzYKHW11Soxph
jgg2gB5eTjKtRbtwfXCnUxyIDocHLKY3T2ybeGJvx1Iwzlk3dDTFL9XpUj8GZIWj
BMCDB5Z6KRaxGWj3os+tAt1b/Z6DI3UQtks/Yaiz63Z/A0Nw6D8+zNume9UY4Ck9
d1viImRw99YNaDTIJXzyzl/ylCvyLDlm+BNlS7k6BiNS3XK8xgHBtHlZPT3F9e+M
yeTdYAVPYWlriqAvAZFVaZtVAg//Mo8P1sOshBOUW+ELM186x4HQlQHtAtFQajFO
VU6GXA27OzoSCX6Y7wr8D/t6mQwrUSBia2J6ubJBahRzshm2OFDD7gUl8s/H0Spj
hBCQhqf+aHcUVJZCIDRJTgkmsBgLFScaDMC7BS3EFIdwwkQBS3Yhp5upuWfsLOx3
h0O2GlgjUsJTROIiwnbdwKyJW9WCYdfiwseQcQSogmqsvTyn6djk/FoFTYZNM0nP
ucUBL7FQSv9Rbn4c/BP7pyVpYi3TgywKr6VSIlTb0KlAajctXAbxNfQVbasBr/hi
WZSdl1U+OqvILZdyOhg37RyPHIUIeV0ArX7PspkjblT8qV9ugNgwSp3H0nILJHzT
K89ZRQQmB8vc9sdyMCuqe8DjVTL75ZgtSl5BO32axmTZBCztDlLVVp+b/kXlWgv8
1TZooFg2ylZE5VGmL9aRFnDgRb9ZUdpx3VFakKiqSCccpI7wcRKoNLInCIJfCRUL
AZM0H7oWw2iBiW97cwWgWqvIRwG6a9EYmdkKs37jy//LdRClm+oyti5K7mTvaLr4
S7b4moXefh9sGGC4qgcyFZREwT+Cbz0GNmkrw+KjvmMyH9RjV6aJtTxWlsBp/EqR
/j1sH5WU2YU5kKzocTtFeZhFqEik2Zr/4RoAKC5l6j8LB3b8Sg2ohJ9DU6xs1Ltd
XroV12Ob9ponb6FgVrdGBLFS9BUFbSeMxUqdbfvU5buoMqrAKpytV8qp9T+wk/Lx
P0+hffTuwgYmCw/3s8Fj5z1KMVqzHT/qR07+lIiZMZFGfOWklAOEb58C63Rf5KYv
OT+UMS+mXrWU5tb6aar7boseKP5nm3eifstCXtZ7tvc6XS65Xj8iz/JzDDRZPTA3
fyAsQBozCxFPuwf12RwPlCiV8wUOGlECOFf8lFO6lOkqfLKgaPcSxuf1+/yPNziP
dfN08Zg6dwc4yIIwfJlZ52bvL8B6cijGksd53e2MWwLsAQvMDoGjLQ+qCPAUnk1k
lQRDbLTNESYKUx9zmEl1cr+TVSTnCJVvM0a95N1aZQ280ImxtivesdMnALB6EYjZ
mt47/uEEYcGMWFvkYLoudLqcIWNBzQ/yqzdg5h1MofAAgNb9Tx0o+GdDddHjKKuI
JCXWNJw+l67YTs1ZDdeaomEJgoCDGsCGTVnTX8HJIfIC++Ys7mPoe7YPBFjLGsmr
iySSx3h9hp3FtL3mOf8bl/n09/HE1oO6/7itrkK0Q3kJ0ffNI5lIh2qWlikyJc4v
YTsg0alFPCLwNF1qJ5DZh2ZhQIQzdKVsNCG/ddlvU3ImTvoXg3wcWyyQjRBdsNWp
pw/wwPN6tQOEEAHNe5nva0rCuOLwKnpSO+G+3H3qLstCvukxXl6AaKnLBi8XfQSA
OKgpwCt8zGG56HNdSNCT3MWu9SEkNryIHwObni2dLHHgPoviqGBFVsqDzEsRIljL
VCjdS0k2ynErnIeTfcA1QGscYk7ViOjj3iwcwbnHgTuREM926+lD2wZX8aO7yYpK
yVlDXF1QufEZ7aLbd2gNqs8zpQGGglPNbUWUSJlwKFw5jWmtFmCgI6rgzde+xh8L
5PLTysOKfVATwCPInzrHmroXo1gOphnB/4gCN6agmDNe5RS7lqc+ksPeSgJOlkRf
bdKk2ljRgYl3cCy57UTmkIE0ymhpECE3+Fgw+7v9gENc9YTNZTGtcA9CVRW1oLYp
otLzdG1QGy/C8brY0cfXdQsdVxRQ1QmTbqspEOonQh6zSJOudTMd5o+OU5bLCRpi
yts9SudcX/BrvaaM+xwSsRG3dRW5wNa+/qUmJRTBXlflQU3aOzVXiYPKG5uuV16d
aHT7hpLXOMpmwz7KZu94zkqBciH/XVtJeT+/xeunMJOMh4FB/YNUh9YczR07V/WL
AHkidumRDmlABQfmmHdwGt8gcVMYWv5DSbN0hg5c8+wqKTzNjG49+bfTGfoV6MxR
RCrE93LBuJ/zwGPtjDBSK3seLljvp2ShvE/9CjQkHeTpWBiseC26O7OKpCk/djpo
7DCnmpOCp2bCqZRi2z12R1phzxijGALwVaEr248Ks7P+Y3kDFGWlX9+YjHXeeIX2
dWfYe+XzTp+IpFPgexhKJWoJxvQKZwuL8mKkNsfwq9T4pb+fQqEk4CkQfmwCCI/R
VWorV3+tK65xhFhZIHSi988koo60lyprhPARU9jJulD13SO2PGqniwq4oebANumf
uCd1a8ck0vtoP40k2IO4JXN1WMr9mSmo6+0RFKJprDJNgJ4F4DGhMkEVdHRWKVgM
PWqDquUhYlOMg4NT5vkM21bOb1rubpx6YEChQPxYqRS22jWiMvseyfVlTSozIBIY
AmFDsKEbMEuuwfyEL96ezVxO+RzeADm1lcWzd758OO9LwnZrf1qHyzCS43v4d0k2
7u6NC/sjBbvFUI6pMvyJJkP4w8Wh0HQJaOWOoZRVQyF/d8OqZ8pfWVK3XFUCEIay
rTUg8nIzdXNM3dSTeWclJoxosLOte9tYP0COiY/yH9aeIOQhvBChKoBx73chkDhY
TX31wFGqQ35BvzfacwDah6y7yKg+2DzmrZK3ow3Zf2+YA34BzZ4XewMJkAFZyLgM
ydoxJH9s7WBbWJFaIW6TixrgbX9BUOW4ZSxDPCfUy8XVzwryGQ5gxH0LTKB8SI3u
J3D8BKb1TttJzwgjmnZUyKkZSqMtYT3dFOwTDy4IJ1UpDw5TdT9+QWLC/hRLJ0PV
QPPNqUBfMeoSVbwWyazAqNsdJl/YYx+tKYgUZfhEHTv1kpE41V2Ehivk6WJ2EZKP
M1Os1Jc7jvq9evX+dDq3YpNFCh/rgtOuh2sxOu6W/zvRtDEemIb6uJ88om4ZeZnn
IprBxaSCX6vzVDMq2gMGLhYYzkoEBKJov8OuyGAXxGoB+hRGd8ZAGYeN3xO9umIX
mnKDiCDMRHrFPIdRo9nRl4Da6DlXMDyKLCh4iECW3joDvhQMGAaMgfnqUUgPqvKW
4F8sh5ZPwPJ0malnmM1kWZzQz2nBU+aojEJ1H+qywxmpa5+BgJSCv+BDbd5khi68
LDDVRaFM4HUIktDqa1lWOwTpVBrIDS2e6l6z2O7TbZUdzK8m75rNwgkhuQ46a/iH
iTdOuaX5a8Wuq7OBj0CCIpTgAWqjG9Ep8K77nyaH4DPjYmNFE83acwy5sVoThf78
x7Ch+K8VwBOuwLIOAx/R5NUvnDG+s2Mjdey4prZs4jxnARihLxCXAB2Ug+SyFmho
fuJysi/w5T15SMiKjJhkSsmejLeIMpG3m51DALzS+jXY19qLd+Ied0LpGtemOmYi
0EjG94tiBg8DZDOYEGjojSh4Z2wX0y4CKgYSyTjeeZCt+XfDRxLcq5xj+w2UtQMg
YNlQR/MtShJca92oo1KUeLg+yV7hY5+32DE8wWCPMMOfZw+nfFcwNQTnO2aIMWDj
HF7Mqnh5QUOMj6SwCr/1tXEc4CoNrYIeK4EVB3gf9paVGFdSVTGMC2enw30c6hIi
sCsAo1CrAQ6+a+ecj4PplB22T0FW+2zN0Z+O+IJjhY4aplzd4E865W1i979RJGq6
fqvxy8tc5+fUeUbyqTZj3HKWoKwV0cVHfl2FVAbDIEPnNQiDXxCrTS421OtUT221
zFw6ROs6hdlzP/AYpaqwg3cgDcxi2USDQ173YHQEcd17D6LUvHpFs+zqxLCRtVrl
RZ8IBKRQ8/QT0EKWZoXRFYVyuOP/zXLVNP0pCHXLhlqwRMfRzhAfQlbLckM4TRGq
WYmAmjwAWeVogD7ZVEyQmdGEoaLisSKjTH1we6FQ0IFuwwCm6CxaRKFgiX/PVRmI
dW8afK3qVsd7aUSyvhcSyRotrIcKTe8VMmOmF8xnsAD+6KLthqr7KyilfGTh7JxT
sQscfv/avMphuV5+hMeqpO3peL54fbUD6l0ROzbUv+6XoFnyjqzIc9NddBYyYLom
IeYEbOe5X3q9b+obrXw+ALl5Irq00JgcWDK4c7d/RdlhWbWPVq1x3Wh73y2IQ26U
5YzyA0uXJl0mCL4tR01GXzWL2bhqCUTgM54bmS6rr3YLHgnDNcrXOmcFguTiiaun
ds5FHeRh79999b3U6Dm4cULLHLJBH6etQTBTnANbt3NZHkXXrv5i9wgXawPJvsp2
5gVAs0GOP5nHMtKgrbIZZONok8NAha4B0E+hKOOHk7DAHvTCvYNQH6i8H2vPTj0x
EfqG7RdV+U4ESVYhC0Pi1jpJZzUKUTQGMKDhI00ER0N8fP/XjApOLGgnGUcp5w+j
vQpSc+WwbizbqGnpHrzAP7BkcAPcR8xE9ruQqj2Ebj3S6PIYC3qJK75zlHEuF+m2
gcTOWSmWOCNsrTQkizYDUwxdm2lSDhZBSQMdE22qY+uE5rZCJqlItu5trD61alx9
A03ZGOoIXuNu9Y6aeatXuwgeE2wUAweB3Bd/q0BxDU/na4/LN4sIKMKYYG2P1i/Z
Wu3BadkDk5NygY7R6aj3hHLn57/3bdd3lSVKhKCuCQzJxG2vvQtjWEFIaM/rVgWZ
WjjPyq6p5FPn8MZgc8eXm0xNcpeSno6q1jyPNamJ+DCYGL9hKOvshD2AsxoOIanG
L++LeorV4EZjv0V2hpMCq4q6Vjt4uCy3257mrjaGG+gHY/QtoD0qFigJLcO/Khl5
n7OAgrMg9onqX317t/Z7CnFwy4ks6bPhMsmYQf7S5yID1Qm9nvBvJpqJVaNBiegG
eqFrwl2dpv0ZMSuDLBTpdzKg5gK5Q7BRRln9Z8sxttUdr6nUGwPkycth1x/vYS8Q
pXJvoX7MgfeKsTRiVYikyWdowe7aM+b4VlrcFqsSBBj1/+meA6cigH9Ysw+hmPdn
NjKGm9XFkDHrpJaG3maDTJpPuT3od1HlYm11Uet8T7DsDT4TGMXw3XrAjlIhYz7j
lkbziQ/0UpNaCzrHdVR3rxg7Rdd5RtrFOm1C6qpVYWi4+B6kbqOxAXpn+FKM5YOv
h83Q2Y1Oc/kg3bGeH57LeYmlb5DcJeziYZjKgtCAoClg8CBIvYIDb/9IWY9GOxc3
mpHT7ZHansrIaU5g2uGMmLCWEaCcq8Fl4bxOLvY/P8T46EGN+1e9H5cR2pJxiuM5
7RWe3LluaGVUp2bOHnR1RtNhOOJXPkduOMxzpa1Rpm3LcYTXAevpbS3Tyc2e0Jx1
BKFa9OH/vKfqgPmApVFqMKWw+UEE/jrNc6qzyNnQWaq4Y0BzFb6TzEic84O9ea9V
qJe6tj98cvkiJ/8CpXqIUTiP3L63GxeiHAfzXxDHT2c9VlaO7E5soyx1i0Itzhk5
qHPmTd7DvR2HF38MN6VThDSSVsDUuiUfv2TVBvqQKve3l56YeAMVvIQRgxuNVfRa
YhUkYGx69oGuF9yJ7NuAzdFPeBSRWukzNxv2kwlOxFVF2ZJfio5Rn1J1F7sIbSgf
b5/wL1g9mg4LYOjVERkv5JOBEkqJlS7oL3s++ufXowMSsxvY8OcI/AT7vMoJLt9L
P4h5QRxpNmVCIGw22X/YZVHu7WKFEvzbzJVfgcNYWAHnybkbtIdQT/9+QJg8vTqc
HhJDI99pPzb9Us4N/wQ26lPjtjtDok8v1D+yfTsUFoDRbHAtXTDrKNzBOCF7EMEV
ej9Iri7rugxTB9GHVXn84yPU6i0tsyy3LP5ukRltSAsf61QckavgFEe7bJJ40zB+
qoSQREYTaO9XaLpAfaHXb5ioshorkpBJ9G0myvpFiZV5yhJ6157kkk4NLOnX3KfG
L9FmJS7YZ0/oG49ijJhO3pFHzXvVA1YO/f7IR8pkrCUn2ALeLNOBVJ/QkaYCgT+F
d8zK4t042j9pv9b72oz1g4vnZHqzszFkud8K6Z/nEYhrNp+ju+7oElyjK2BeQNyt
45uCU9AKSTOQOw+C3sLqC0VcagFuPCrxTRbDOKm27PWkDtWvzXqDUa1HlKt/NO7O
DjH6FNQixbLGbydmrueITZkKjb9iKFKYkOv1FmhKtIptNA/WoIntuz+JDZEBJtgp
yU4sk/a4yj7sf/l23lvse1VBi2aPFkH7K9FRG8e5BUegrsAR7vIVywox1OzKc5HG
fHfkqhMi3HF7jD5uPZnDd80EMpC9qMJX4jaN2rDu/isAudMGpqOrz9MzWE77pKLY
b+UD2+0YIVb0T3q9F6LdmcYUL3auFOl7Ht+bwTyXTkzLO/LWs0sA3df4O9Mmq0wI
S7qYIWfG1fZWBM85LOztRvWbBmgzeULuu0b4/X/15+zznOWJnMtqORgzyre3fUAO
UIZVY05/6ecY6LrnwWnxLM3UmzLo2FOuEWTa1u6EsFOG7/r+xht0DpQXN+N1FFQ9
SX9NzPwWPUUPI2tccX3fFEjOiobANqjxCjQ++tbnGmyltIpvMIjUQYC5tw3L1IhU
PMej45Xivsshbp94Svku2iyQ51mBwugzHzFPzHHst6dDg6/IYNgaZzx5609cw8vW
eZ4ZwhKovFbxUOCi0x/QyUMgOGRnurod3ObvXxQ7Uk9351NfOacgyvPEHCFSR+WL
KBoGzd+83o94RekQqYb7Hg2MG+gIWVkEmb/m56fxjVV3YiYcTpHu7687zGVZqY+L
zwuqAIH2AqwWE80ivHzJZJcy6omyQix9tl+S4MGCjppXDzJ1WrpP4ABlYHQzId4h
Vg3v/Sc6HjQWpaQMzgDFO20wN18456qlFtwoG4pQ2LhmemPRHeKKBcao8ZLoqt5/
ojX/BZLveWzzAkuP72Zt2jaZa1LuDI7ECMUQFqldUse+5zvoCTKywDc5rcgNylYk
UntIJZXQc83FsV/fxZucOrgVgndE1GgIj3xZGBtHawa87RF5LWUeaITsg0jVxXdt
Tkyc6lSXhVkoEPhxHIaZEZJs1rex+i8VuoNdwZKL2rgHzUOjEywl07ia/krjNZ4z
3lmdxVgvF0QAuHoNk8k2HmVBTfgPi1aU70/BOeze+fjKMenJSd/R/wQkRJZ1J9ZE
wLSyAI5R25Z4NbJE4sFik7np7Uom37DTc2cQhXp2FoX+Vosquzv20WL3XebMEfoM
R+xDzr7qdow0x+JvSoHU0/RGVz831iVrI2x7kvUxY1jhBH6YA/CEIj5NqE1mg8PF
rTP2TLOhCOg1A9zm9nFsvNlo3O+2dlvZsH7JvVuOerRV8eGyOeOzH4o4kp+/5sPV
9B/Og+Jj8di4ydaRty3KWDs2WYIimH1jZq+Y7z6FoDQnHpBvlOnxuGk2Mjw1lPtc
82rEXBTkW8y3Y3CHWIvyltTFevtPdIfksY7i6SQ7spNZm7gnQH3qNF26ucQXAp7g
EPZls2y4Ceul6zcD6dvbR/f9iNT5pn2qwGhiH3wKLg0RcZWIhAt4nWUCY3bvMxuU
gHS8QA9HwT80elWAo82PrLCuYyb+RB+CctFjaMVyykMxqgAAF9NwJrCOVlUvR22u
OTlGxqVZZMaG4VxtSCcW5A8LfGOmhGQ1txOEUduOaa6oi+Alv+6kRwj6++eMNF9J
b3qXsIQF/dPjIc52N8kpYPjSO7zoQwNzSDL4CkKG6709h08rgXcfZa5psnREAsHq
eEGre74pJngVzuWMl7wCsFx+JD2NT1Z82GtAjjJpH2elwq02oYwi4DewcrsaDLHs
WEKCXWzGabEqHqRQ3yCkfVDVDR1hK+A575iwED2LFxRUl4w6wQZDyv3ITrEt1jvv
b8B+NgBSK0MgUsQ0GCNZs870yKfFAXWwSmZdf/7dwRJunDM7y5niYjIfCqmxecI/
pxRkiBoSQyTqjYdkzf0iioXcfdXhHZMmUEWngdG95SUjY2i0HuklXTzBZn0aUE3N
geu7qi+DUgsciC/dkgTSmR1eh1y6lo6QzwLz4HXhr9oGQhHTO2LiRNN758xnNNWH
8fRj1dp+3ff4fOOtCGFYx9zWbqLPqkNGIys7tPPDn2dBxTIEhmjiUHTbNrjMiq2F
CIIfGwOZBPNeRdOxthkh4QBavEWeA/tFKp/8xLRuHTaGEsWjrQJalLuK+COKRagL
XhG+N/sU0G2UEg895fzhgUf1uC0HmAsSi8iPasUO66WAu6mdNKDXkEFHCiyM/e9M
gbOgjcPXDUX85RW8bvua1R2QfxakQXTxw9UiTKfxxx81ikuDRrb/Tgwsq/QYHIW3
9bJFhhVOB53e4HUdAYJMDwj2JiyLVWc90G/p7zVAh+31wDyvPE/4+CxtZ/O9do8w
CE7BMtax6oKhM4a8JPR/G/uEoOAyBwpoivAJksC0SD6rwCm6+AK2F9O+O2vruj/e
N0uQqvQfRXDJdydsykdrdOThDlZrEu1ei6JGEtogxO+wXkJ0vUKq13mXY04xTTBg
io6G4hOiVk+CUTEzh8IVRuL/6AJIkQB/9UzseMzbQd1LnNXOMdTr9qqbsckrmw95
93R7pRNRj4K0CS84ywBb0gGtJb5s1br6DrdR+EgUwKAWjnZvqmxLHbGtU/LLM0M4
nGtEIdce31C6BCtgHr4xivXaRCnkFGt+3IZJiJLO0iil6Yr/0mpiQFdQYnhLEegd
8jsmgbvpH0uBqSNuYCVaxwqDDCDGKhqDUTfL+TLexFbHtL89VQ/6X4I4GGvH2B/k
whbr2cjMchonnxWpw3tE+EXS+gLAmaPki6XGHcFc8a5dhoJfnSFiceGqhlJzcYpJ
eTjnqnDNNB+lUxmUExRoR9g945N0WbzAVay12eY/24c3580p8paB4a8yJcPtf2gF
H7EGm+AGhlzcAGyIzYq3mUnvNPFgf3/dO/vaQp/PzhSg7dA5BZlPlvyPzOpDgIMp
cnTCYslznsyeJeAATTLUZJeKEAdmWKpTym6mD5NGDtVlTSnuoFUmPgWRX6KA90xX
lhUDhlX6LMbAH+X+chI460PcwWvekO92ZNs4WuK8OVEL6MPwUDCKI2zEtdiBDg3C
N1Qqk6c9gjYnYBdsJRqcdr7HDELGSjSxd68lEBtwxg/vY9yL4GXkOSCyoOUFq7Gu
G6pjY/8qW9r5kBWiHSaHymOqLre8Glpiw4k3BNYL1qiohEG01g6SZpmCldYpNRFa
GKTIf4oH45YKr3pO5QJ82qkWGZUJb6/r6VqALIhuOmVyKc4KgD2xTgXy6F3kKCeD
efxextKm8eOs7vGmDT1I6VKTt2anxdMKcl4ddtGqhwCuAhBhNF8+UuK4KoKAm4u3
LK+V30Yq1ixqVwi7h1HBIpp3bTTGfV8OyEyAtj3HWfrzjSWkd85MQvbdcwFXJZ5d
e5gan/DsvpXmMVgIqQYpieaWcxLqBbGgbdwCGJE+xwwWJnbhwTJ4I7yN1BCleQN1
1vxhgOZ4Ba1qmZI8vOiV74qyyGDLwTBfwAfQo3zqtlnwf4nlH/rkc8mqXzqHZFvm
b1zSGI5xTtvGZdE4WzUJ/2YDcKiKeIWT/mMkmuEVeIxZhH5v4ebZP9HppML0rLbV
3NtQfxye2mfj8H/q5zhuFxecmls3b7tPoxeQVPuGHEnvqubKok89t8yfK6B9PT72
p+M9+9qq7/XeTl/9KqXiVQlavpaiOfP1VhVki9D0XuwQ3X/zYKCYqfOXb+Ta2zjr
OS/MGuYzFgl1mhhAKuUyifxMbiCo6RrgnayjtpO1DR6YMIj4yCwCVNwpnBBpVpEk
hJN+w0sk7hvepoRwbFheClhkuWzb2ugRejV7LoImIYYPhExkPeX0m00KH3YKho9T
YdtRAF2ObmYEo9+wihIZfnJ7OLK5j5eQfOxUa2v3Mt8mqHa/uGIhcSRoCn1VIZS7
oTzI9DHAoFAz6o5KR7v+LjAApiYLEiOirP86m3fhhdNnu1iCpMlVLy6omeXtG5Te
S8ZTkAepsGVBZxtm3+bPy8M9QqpWOIasQCgAhplh+yAkP92Xr0JWFGaQvFfa9SMi
n0JxYP+pNeclsVnawjrOahn0nGS9oEmICn8+qtbgJB3PS4tsRYe7A4f4yJPwwzE2
Lnh46Il+sqyUdY9Ne8MTTgcJ57s2m7S644/2cdQ9HTcFDLXrEN6CMRnZKcoNOj9A
5ADIsK57+UzEa1FtIPQkH7uySl+G8K1P8W+SrSKIDvKAoykOJbG3HPnuNyPRW/Az
DoIXq+OFP/+poJxQsWPk6uevru8Hi99g91nBd6+kbifE5tpaw06Gr2Qlbdb2jbjq
eqPSQEbRx6Vgnk3AfF1gsdmD3nIDQg1C2f60kDLme/j+kkJLPL2SmPGYOac2C1Wm
T9sX05RmNI3hRFrjqfM68YeDCIAgrl/OoxygHqbAU/MfMkiQ8zjE0JsWvT2Kigpp
XuDOf/2Lv9hD5uvvp+9GnaE+baHCCOKbql2wFO2UCIamFLs2yQynNJiXs3OAAFXx
e1I8Z7AqL1vDqMiuUXMVXmu46aHXSOMb8dXHQokoMgVmTWIk0YafPZ+EBTLOn7ay
l690Pzt/XO70lykJacrLp6IQnEriIqcybnaeHodlFFiRJD6v6/OxZDpDd4RDGgU9
kD123x6mf81RfOu35RTGoy0XVq1QxMTvD9Skjv0vZ1+LB3iAcTeLcdfF4MIz+Sgq
R9fhz/kh9nFFEpjQtIN8EwJbXs8xvhbMPKhvkt6lG+XG4CjRnYIxYZXTX0tZ34ZZ
PPh5MkOiHx2js+nFlXKjhFt0oTKeg5KUZK7G42FLMZfAvA59CD5095f2Y+5qMVGd
4XL8o7EjRi0c9dpZoznmpFLSZU23lO7PopH4RTfdLySC+YYezzo4o+MpjI0f665k
K4UzE+Y86q3ZjIaCa2NKeIKaoBAuREaJvw87RLxfXkcfnxpMJnsoBqZ/f27+rb1F
1hCCwk5ieSCtugcYC7yeZsvoz+HbxbUpte+GYaGoB2dYkHWwovBNO+b+JrWkjanU
7/pkgT1fBSdEh8GAvaPK8hmgs69ycDgID8tiYkZSpN98Vy/iqaGWyRsYr01n2UEm
QL4clI7NKwCFmiT3BVhVdWd+zOyoPARYl/tzVcTNjwxsCKD86hzwubk9OMVCp+ec
gTWsw2FDxf9fVw71p+UaO5A7OZoPLiJNQXnpsRkye01xQQzOLKa5z7Ic1rk3sfwz
6uvz5KgXMqLkNm4HEuVXcRRUGldHo4kVaSSmfqDO99k5CPa39LgaeK+l4ROgpoQW
8jrZcq5IQvT9819ImzdoM+gYaa9LkEGwHS+vz37qojaO0socDVm2t7nSmj174rW1
rR9b6hiYrgv69q0eV/qC6r3jjC0vm4S1P8piNT/+HP+Gp/VIaDND9+vCIGQckaHY
5wy2rPVzByvXXRxihRxxSf0upLxN6YEmVR68i/srOBcT7QkhWqSchwLSxBh1tu5G
y6nRLBqfC8T64P+g6Tn5QKvp4ZbYGgGNoqObvm9yr2utP1cVjnNUvpY7Fyk+14jv
hUvVZ2/tdKCB0Cwirt8kloN6tsTE9jZspFxk823MzKeln0+qtqO3Ip0u16l5aPFG
87b23Lsxu757lcaQEFExnY3uGJA62HbgkxX4KnJRTaB8HODRGNQu84tyaQcQGm2k
pZzwB/RR0bIROGoSdTD5f3RS/dmjFk6MVOIyoptZld5zbyl9GqKgeUOmSd15SwFa
GmhtdtRVpJ+522V9QbO3zrsYzCwCXOpOVgT4U7pk1xqm0Hs+Jo7w1kp7SCLUL9li
qH7EFXKWmPCRE0/DNFa51komXLMeDznC4c04I/VGbt71bmvAP9GT+Wx8z6S5S3BS
prV7xz6wLAnzOl6xQ72fSA/lT2zmX7ZvQuRSixefXrvt7KwnyyjrRRdwmkSMdYkn
GuI6q9PoWJjdrA1hK3WXXqUnWoGWpkwEAIpRHcY/agfESKIqxq3b05okiDkC2g1K
MPK1TZMC02pj6xXFCN5W5xkzPMIpTJBstjcyO14j8rhR4aNp6ohYzbXWPNfrHEbA
gWsCB4ss2P/Gs5R30owSaSP8tg4O97VFkbD6zOGas6aVNfa5LIYnXK4BLvlTptOo
n/aXycEKK2lhnAGdr2K3ORHiSDaRWH9lv/IlT2Ji2GUyJmFAR55X7lnwULxvyLDM
0tKJaQqhXSpbG86U7TYl0tLtHuyk6tI0C2KQNQ3VqiMdThb3TSSe5jvkOLhDNVZA
vxzSL2CRQolgif/a4yoDuS3i1rn+ctD0DcqYOiwVUtigFV7nm1KHSBJjL65Nz0HC
mGXPrF5xtvjGfLuqAjUL0xYP8Ly1smlqFqXtvgJVxacqs2NLfzEM72vU0TeuuBmz
wBlqel0N67pYv4LpZD3TSEFPnmxvrXVwzxaMDy4+sdh8K6bdA2S50W2u6d5mDZmP
lRY0wfvOyPnSZb0I8AaOfGuzloyeuMecP1Fis3YpA+LX5GSZ7W/h4yU16TwrgML6
0QXREoAiUrBQ5sMgM5IiE5F/7G4mUVRZDv+kATMH4A9Wjgv/9+j2WAwlItlF2uBa
Kd9mK/AiEsq99j6Zgx+nr+VgPmGdqwJWFaQkqvp0gRflZeJbWhZJ/l3f4EH9pXJb
juxGK2zm6wdAiCDND4ZrQa3azjROYrMbj9I8XZhGCde0CXAfaxqcUhlixwVCHmXg
TeZESrJ4tVZUek7UcAKywjZFOP3fNrDaz4wv1Zy7Kc0SOoL6X+IX8t8oKKdHv0WF
1LytbvDWCB/Q7VpGWxdTmL71NSpnXY4PRg7n3Y//4AVjNmGz6ZHbV9Q+2J6skMal
SVRSUCb2FBGCIiVWNOuuPUWs+H2Q3WyoXcGyqHOqbr/yfwZx2QnkwKuz+WAqnjQy
zCpXIjF+/7hR7pXms/FTJMDV0NWCNQhRHFAPpXE0J0eOTn7Kk8r1Nc8LUE6isRS/
RrDzmHQtdz3oUG2Ab6OHtaOFxUq+Am9xj4kDBC/ub7AMFp5WviPHxJIVxdBy9p1N
kBHhapXpbI/T7Fr4MMqEczDJVtmZwyNZzS24O3QHJpqPlmXdDv6gmXrvEC8QeI4D
5BhSEUNB2/svqAXyD0XtTev4qI46SwCEdlCQRFEep/6VIVNbQNz/gvyKGnsp1z/z
smBrtbq4lFo+3TI/GwOccrIYSWCBNMf2mIXdc24QLx8yYyeryz5Znt81obDVH0HS
F000nhpgRsRLrwnNRPDy30hq+Gh2Qtxai+FWSVgh08zyJZRPPCM71Nm63JemAVde
ATHUnw1PYm+2I2d+0ia4BNGtSrrDIdcpONL/Fc9HqBwZyMXL8ZbxPtuignZP1su+
24nr4381zT8fPlJ6MPBUsCNNuUpTA0S9I4dLRZ4THT/Hm5p8bHDQmXLpwqwztqq4
Cs6e3GQDkUIrVZwlgyFgIah9vIaN8A667uJOuNnUD2pS5a42bHp2tfz+9dBR7tsm
V0h3ap8dA1eIHEWx085ZDNiz2/96j5i3RC0meDKrqgG7r35Fdtg+AQGq5+mh53wr
G3dqjnORcHCTC4K15y6YCxgY0EhctS/SiLw3+1SuD0+HeC5rGoTCg1F7z9JhPIY/
rRa1x05fFEU9DgVEMp3Y4wlR8kP7uOvNpfnjtM3D3xzmuBOA09kin1L72WDPBiv4
PdwNie1qOKeCgSC416gFxHVf1l/SMjro/M8M8/aH5YqQSaK6oSOU/C/51dz6haJ+
UHMsK2CrD9g42avzUlFELzi3GUJB8QpGXLrw5xMbpbU6sf5rpFikmcQN0GQBWOav
yJJ/l4CSWw1tCuKl00ROzCUXLZMgiDIVnBEYRKbvXFkuQ957IJ63psPYcMAA8a+n
+u06R6qcj+7PNaM8froTBTcQT85hsKiocoTeXzoZr9WN+qaC3NOTkTCVNkmWPHLo
tcs/4bGwsQVG/c1TwJ19nk/cdDBPWSJgsndUe7ws/2rSls4leYvZ6hTSYGBMtUq1
da3Plv4vtvNMly5qP0bIjEadnpOSmI8hka+zEigwa67RQr6EswybI7sHPK8QIFFU
Ad8IHeKPIIPKFHJjQ8FGsTo5FvCzRCuEyutZCWzAnntPx5Rhlz2l2D7IV0mODJll
UQ1Rg1KR7f3Ebd/TWyBKVBGpYjlC1pssw0RmGvjEC0t4fhcomXY4c2H+jAHCe6YK
jVsYqo5QSwBRJlVIjlAH1s6idWVQ0igC6NpNKWD20cWxG6dBirUhdM4/imJA+tDp
CtO95ly2hmEPrNcbxwJ8UunC03pfu5fQJMW7i+MSDyjefWeB6HbbsiVnxtlbuWvn
KPdymb178a1Rpwo2Ghdc3vgLlil5oR89VffEzdos6t5DFjLBFZ3wlpX2gzvqQwgv
0rFGBNFutepCLm718Ro/8zgWzwVPw/kmpyNMGqFA6n5GBg5vD2KkuGxOujfiApXW
xCEF5O9zNAxXtaKO3cf6CbAFLeg7yITS76LeZHTvTAUBsaVH3Kht4//pyjjjfLom
ZTTgOEK7RrS5x/3bBLCHFRmthFzZGwye6g4XA5aQkfXotiYVmo2x3q35x1psBW8p
0O3yE4XRgJ4mVdwHqvNaCPgqhGOTZMVaCUCpouwPErfYDXxql32JixJl42Hfn9Zv
fhdfCgHwtc4SK+ThATZo7ttEl3eGdc05mYFL7jn/eXbufTeiCsgs2V+8cl6qQjHQ
wPq1Tu948ZykHqlIRi5j8bfqiFeaIxXv2+qY7U8HShIYDb1F9SbQUw9Q8x5LqEy5
eHTKZkPXm3J/P69xwpH21/RhvF9d9kMG0J1ZtOUgb1XFC5hQ3OfIYePmDxF7pa1W
qIfMVIH67L16RK0M+3bUsEQ+/mTiUSSFTEyZAQN87ilE+hgj++H7HPg52yvxhucN
oUnzv61Ra3bT0DSiYhxh5qbhrCjHLl6EdGw4HUlaJPc3qJNuSR04x08t9VPQk8/7
dnx6tAJbSF3sX9KLX7zS3zM1k61c4HuaNl6cmhnhrgDUePM2CCMlLVa1UgJ/RhZG
fq+pG6npjTyMafNA6v0kv8YdYVaR1SPGVxIN1vFIwpU8bwzTr7dO9el27vyGfRW3
umli2kHNTvU0UH09nn3aYL2BfS2UCeV++3j610Yy4hXC5r6xJB1R+qR6+lvXt/zL
NRNc+oRZohOCuPZT8VadDSgWSo5rHcwEplQpI/98diQyxna243/vCcwl/GwFQr7J
okA12PRI+g85mlA3OsVKwg2rQkCfsqj5kQDigjzRwbjQ3GUbeZ0HweX39wiLqtpX
sqfOAaDN6sgCNfOs5I9NZh0qe8pGjgdbmUG7hxzR06v0t2fjlB/9NERxlV8Mev/J
nqb8RKCWlaejjwBW8xBWnf65Gh6S/mkYHsevR/oxZ2g5FbMefHFqB1j9DUOHA2TJ
fJfd3ipDRmU4q40/NhM2CCSJMliF7ptaOrtFzaMQB2N0qRE2GD7+iyUz01eZg8RM
YfiH9+pQawYbK+0br1/aV1VLevAq8VGRR0PZdHO8XR+rW1QOudi2W72ynRfOEcxZ
jnzKMGkscG0ZP0Qs06A8mHNH0uzsjcyDJjnAKPHTxFTdoy2qUF3gUAm4ZOUwvdhb
8SBfUxsdwtgdDZ/io3xj77rFLVUFOHX51zUkMsDTj7Gq9Loo63JT5GIOaMQxCZAL
G6h9CdPEJrcIL1Zug05IPNBZSASyCVCZa9q88Rv8lvOfWSwQt8+NK0hN4FbMAjnB
U96vpHYZAB2RzT43/0YFZiT6IuoYQ089WfBrPMXOLZUt01KIH/u6iYLAK20pLkUG
yFikOB3bWgxFvdBUIXgy2juGTt5ECeeYNPu1y4C3ZSKlAUzptmskFpGEfYg7j7MJ
tT5krwAQi2L2W763c28xlA3jigIJhRdoCiQVuzROCbyJ0qrgzsquylitetUfnoDP
6x84czPNFzn1kGOcORXxlbvFOEvAKTVS/522svIFNilEGq9ycqfU0zHzrizgVBPA
QtTNNtP6O0EWdU/pepyKhVxV8waw4gAiBz4p0oTbw9e+W0I7cJifaqg11yUvntEr
sMe4bOLoyV1dSbVfC1hSvrChkutxW7FCUcPDQ5njMdPu8WIE7VJf60TVaZk0gK6Z
ppRZIG007a0GgvxXn3kQWaCWLeGzMZSp1KSIOmyzhHdd3BeS8/BJDZDZEbj1RlF7
IzYjp2m4QSX6WbvLIcag6nMvg1FXt/sg4cZKYADigMuF5wGJHUnoctXEKh36xEbl
iS1fgh+9GbfQ4UUbJcwugR+CdW7FaYLrGiFqriN3JcDFEwmTABI4RHwZZPJJ/JDH
d588IGDm0gmsoY5LqFl0Z1QbA6DxhXEmzPqG68l9nxmXA0/G6k9lMmWkiEzcVwXb
svC38JFhBxmZqiR511jr0xuMl3hg74r8H+U67Ekp8jsNqoCwWwNzPdAx1Rh2v5Y1
QetWEMigQBQ1WQFHY6P2Njn+ToGp/FSLaMH5MCWUXp9p5S4H/VLN1AWFDhOF9WCX
HZuBecrnMRZ+3j+dEyo87En6IOIQ2z5Lgo1eeCb3aqoOMs30gRwi5ax+7KymGr2B
0is/D9VQApRKGWahUG7FJ994sUT42uXQ7uPnAWsrqrTzJGpPFq6ilqJoW/lQRvSh
jxy5IdyvjDzbfVvEW2obDhir3v9lY1pedEs35QBzoaBCVzuFLc0ZUlSViCyNkJQG
eewKt74gXuGd0jTP25NeZGHYfK75ma6pMkwt/3kNdGhFbWIWB8z8FlQm+CSEShkm
lkyDwEMWfgrE+EAN9R2ARe76B4vgulq2JIIPQ+Tj/vzEu+zlkM6/o7GU5b0pCHPT
hub0dkLWpJtAekSn7O9OSKbXDl+SOmxxab0Tk9e3ZIdfFXEZHuJIjTrI0kuJPzkC
e5d6PSnwYRXW4JySJVx+uAHVdLLT04OVRvamwyKo7pahsh09rD2wbc33DMeFXld3
kS5tNT1OjloLawtiHDiFUqQZzeYsDhAQxsm9qKFoVEGvNjRtIB7n1xSjdAA++4UR
aWDOrDdS8qGgT6mCUhurf7UB3d/HFc4wKWiAgNdjMIttV8DTJONl25Zn3HszBAI8
a0+7Fnog1qa4sxV8K43qDP9sJc2+IxmK58wR0ACd5eDp7s6wdA3fcpzBK+rdqfLP
r4gbILK5v3smfuI9GTTAycYWqQ/8bGviy7VrOWuzcHtBjgULQGgcN5/bRH7Pi0tA
BtLo47IxkQ+Fs4s+MqUyl5c74Lw71v3LxnJPAEqBoBsraaHIjruqK0QehF3b1M2Z
/ZPcvjp6b0sU64RDscWqIyanyU9nvxWXUWJASUDC14mmimYVKHgqjlvxzRcQvUqm
lon8Usu4eAzTdOWGK1PLIBnRCeiYSN8ZgteZu7lM7fa8PfEUodNFp3o9Wd6H4I4t
nbIQ1/IOFn0NO9phDDdU+Qww5o0VmC7WfkVe9pD1nzW/YtwCkJmvamsv3D/kivZc
NJJct4s43NP98GwTjVpngUNmCTofWaKEJuh1e6Saek9DaZchLJcTrogyAkoynD88
zHJ3ZJm5i3o61iUolduku5MseF9iyt+VLzTmWAZZIj+F8nvIFvBcxMZ60zPx37Ni
bbTssT6I+v6kAwqekjM29GibXXhmVSrtPbFJgcQX3HgvJqPmGdsQDnXlX1xc7+LO
LQq7hzxiDt35SQye/BkqASc7Izxx++JgvuKFpQM+kXmQzQd/Ia7EFnjYhtVQ9v60
C30Y1rHpGcej/tIT/BVWq9uhPGO6XmndRXfKeSiWF9JWoDa6crWwK/HaDRu3VYcC
dEbnPY+USWE3fYc7tS2QqcNGYteCRr7o9Srccunixpt/plPk5A8O9c2g5LNmiVYE
i3TjUiv4x2luvI8bFlNcylmbzI6tmb0AcBGgEPiHVOKIODJEkalug3b/x+fqIrHm
UxIEVjmRn74PrVlLGijUx8OHeI6FN3+7WA18ajKdRF+iAZliCTqaDF6Qc4uHT7kp
bGyCpA/d6QWYz060zq3/VcGzhY9kNZwDbPC/mVVPJb37JwXouyCOIGx1C2RPzSLh
Ei1o0aapLfEdQ1oZdd9utTVN/ouw9DvyzhDFc4mTJiSdy8KohrH5KCnmVehiuzqI
KvQIslNyeWUseSoubB36ryjDXVpm5tS4ndtLHxN8UD2oGm0OHEYYlMO85nM4kIDc
nKlyNYDPGZGQB1CefI2yoqptaf0IeR7w4ieJvCg1hK24FL5VhvhGBttwMmRiE/0P
FKLUlxDgA3WCjGhW6HbhplzDKGbNwVL3haXFrEoMI45vkReOhBg621Ps5c3YNHlK
QlappCYn/rzCi098iE9md33r5hlX8Yh2zSbgCcXBhXSoD2vxA0U3H3VzrHqdh9Xa
mVtVGj6sWb23y7Tv8su5tVZWPo0Hp+rJk8bOBm2PFiB7NSY4CD6mZKAtgEuvT4qA
D2MMGXvkKoJGg7q+hJBVlCcQbh+sFxUEsHODGOF7QE/66wl8jlwpqTCxvb9IHoDX
u7Qzg74xVBEnMSVssTgBL9ORE0dPMJYNUtiU3osK4TqZvOtLkB+uz/FgLolUz8pP
Wcs5DG3eWn6RBvzomKwKV0I0tAg6LigOjxcrmuIbzDpfR1D63fy9aN5yGezW9Xic
1uRJzPOAA4VuNQQmS4k4B2v+XvspdffG7PjKbZewObBqGPycPiIPqJLYYdGd/eZo
T5k2kKavTKCAh1wnd7pSI28EaP/ni+v2ivy3vPZQhYJUJ1wqel/lt0EUwA1hv0No
xDO8Y4heZJ5M3spEPTVGhRBVE1PuBOeUWhlF0SvwhTp9DlxoxkYIJ45C+MYxnbGB
Owy0SesQaJnTfXH5E2iN+URrwQev4j59JoguQJrmLHKuoUoFB4XP2POC3cXG5a6z
hBV9+2jRrRLTOxxjmkpEyczWVE6x31yuiy/dMWV6ixqm7372D1NHQF5TBgSaYhQ/
xwFD6iSb5UCgj3XNJXu0jNSIzALsbplxCdztdVaJu2SDHbX+jBiSBvY5MI/eWmDC
tD9udXhfwKDCSjYIX7oLoIPU8v/BsTRLUtkIm+r9QjKQx0ewLtYuUgczk6kX0Qg/
AleUsvBfFHV2bBxDFlrXnFedsVsT/Zy3OPEQd5y2LDEQ9n+9cr9pK29/LzZYiiFL
sSxiqSQpWOeVvwDwecVfmTk5gMA4SOUcWh1xuD/R2sq4PPK+nam0bNTH6w7tkh/X
4K/wNn2TKzlvtJqsnVeAUlTRdYgjhTbu7gQxvsVn2l2MVZVi5lymDJD6FiTIPunc
+5p3BjKqbrIkgUEKmELDwtKa9lMs/g2q0YBNEyDhnw5xMW0AdL81SNTSSag9fU4Y
QeqokmnQafzVvBv8Ihg2i+ifDubnX9xn7QDy0wM4wsU8MHQ9apd3s3Agqj7vqk7h
B3u6xx4ACz+fPyoXtlXvqNiugTMe4ha/tpVrD9854G8eRs5LnC0lT51ac2GjN67g
M/qJOOFwkR72wWm4fAglVbTmF7h65aEwZbAcMgKFmBDdo0YXYdr3uJlvibqIg6Ua
k7WPWL+s6KlPql9xWohOpnoLOIHCzh4ZxKq1em2ZK7BJ1UWvuxz8DMGewk7mqHox
x4ymsIi7FSoM8qAOG2uIkP0jgGES3Np4f5AGABjnqByAzfPho8xAj6sPdyW8eqU2
vYy79C4WyQqbEKqvKdmQLR6cXRJE6BWTIZl4bKUkog4W3z6kpNdFVfEBnjeY2agc
ZHNAITGNhMa4dSCwuYjYtX5h0VwrEhqxOAVLyXhRreEUEBlTjYIBP2fIRhgp3U0Z
peamYLotbANBzfOhFjxJ3tc+8Ib5hYjpapBXHHIQTAXhEJ4LngERizhSBfE1fg39
yJ+PVWek+WIF5JMcL8H9A1nohG0cUjuYHHiP8Ecngu22NynfMyg3v+rpJ+S8LBIU
MWhw1JBBfYVSlKQDZ0uxfdRdgznbbrxxbn1R/JoQjFKKRpGMK1cWfyA4Nduz7Fg/
yAoluHzMsIDQmv/fAbz2d+H6NFADuWyZrHTxaQGZYOWkBJkobOxsdh/IWj/B927G
tYHcdFFhH0y+h4t52zQy2qj9qf3hpJCz4jBrtb3VoM3c1Hm/ZtTUxlBSnRZEOgjN
pNU3NSBXdf99Dtom9CN0ZhYZQYaXVW0pA3F8vUEvuYM7qqW2Uw487gr733EcBLFS
IVRzGamDi18nJGgnIch/CBSdo0fTouKR1KdZNm1xsj/vxwRqoctgplgOT52MmPfs
CIERyhpjAz7XaUgm4tn5vQqLqBrKdoO0mpVsuu/vZPuLgG13EhQVRkdE37/0adjD
JKV56O3kK4PV4C3HikqMk88r/3d6NytyKzPktc/OEvMXEa3zL/vQdZws7ZbQQtzG
EpuJoNh+qI47WUQ/wAcnepSm6Cz69C4libJdFQdeUFtJOQz2TIQgOa7lH6lu12uU
eqe3Yk7bSdnPWyosp8j6CCwrrSqnMyKpGtrTonKVHKZfL1KhXIaZkkmniFoYphVo
MemksUn0hxCEM+7AqhoKz6q/BXjZMXAE6W2HgFy4OHX/fwUABfYGmecYh0vxbszC
OsR7Wc72fgz6OeXo12a9pRGFBpI65JARHRmv69Ez7aSEnMKDxJad9gVOKuumXHxY
g+jJqKwban9GvBSGRfwviNW59w8c9bAZxxWQgGHhu9/bW1v4pk5F9vKvTcaSe02w
R65sNQWlJET9SfpODvCQyXUbLRgls2ZE0inN7nRd2EfwW33NbwE5mx00szkvQCsv
iAEoNt//QJXrWettiUaDkEbky88THYXwo2IQjjhaHeXPbdZz4+2RqsDayg/Pvgtg
wQALwI43sBAoUrzWl+SIbh/e0gT1rbN3MKxRkTjI15ILQJwwv+HUPmVQVh92fMc2
ZeBYKyPDZKN3k6OdinNY2Rb7UpgjhmgOOLtp5X5GMiX0xsZFXhKp1zMd1i1olaKV
ltOl9vCDmR5/USf/G6E93+mhjmnDj6MRw8N8LCZqoWPj+phXk9v1qO+hWh0/rsra
dozIA55s8VFWJ5NZ8JulolmWS5WNVyNWtrakHPwE7ol6G63ru9U9Pm1HdIEGkF6q
FuK/woiE4tnd57Cbjn36HnLwrzbv8o9NdFdjK+m1xeAsaYAqHYqQMgiyOABCbL9w
F38wMwhiRdk5YHoUmSVuJBgl53tPToqdmjUYPKwtr/XGoz0aLqksmp13Y9tWYuy1
pgp2jZhm3JcuC8OKC88Cm5hE8MFe9WwVE6tntdJzbE/zHrju1RPyBn9CR+Mx7YX0
zkMBchVtUTda3l1Z0gPLcLBBR8kv9EMOHJLZTyD+beVVKciX8MfYfQKoWsuPJp5x
IoYX9B0Et2Tp6wIyZa5C1RitffNmYHd/9XyHH+27PDn4xr4a2OxbO0FKRqsHTUf8
SHR8YRukurzSIXT8lMe55te+ss2PsIevtGVBTQJaSNlP2KHQaYnHNRnAok7MiMvr
mh77X6NUCJXgSXp5GoBUbtk8wp0d2YdBLeP2yIue7xcenToAXQFtyD0P2r1xHBsA
swUjOvV+CJaCuzec7wXUDHxNoeF0b8xfK84V7aqZrmYd7I6NjCPaP4tMZJRzU084
eiZod/czclWOtQXYlVd38zXBcx9bytVXYzFA3m8tiVEYdzxOXuSRmdHEv5KjmnRj
u2uSG+QTvlfsXkni4gFMyLn6ROS6UfE/+fPhVTIIUmFBleUTEgpBNOzeHKD7xWym
WCVsFYdULbPefyf4CUNOrhzOxHKExifn45J0wsQSKCYI8shGPcZ9eA3JSnte1l41
H9L1ju7S69RZOmTJ0knKIzd7jnSMUhKi7fo0vdHb4rCGc7QPTdur0KhZpVO+dRZm
Sea+rKl3aXfRZpjUpBsIyuSGlUv2Fzxsrg2Dqwkiukah07ocXHhGj/hZ4gF0jgEl
3QQBYpEHxedrbAi+eTSko0zCEXCi2vhjUxB6YK68+r2FlXDrnmYDQaZ57/4ygnHi
8xXzYReAMHML1lAbpG+M7g5MJsqMI9Ak+HDbBZWFKyU6X6NjGvTgpMW1inFPu0Iu
aDP707f6YFq3BAwZ7b3ZE2zNOJfLxV0d+Y84qHbA6/q8Q+tS+1md4egyXv88gDCz
gRkLkaA36ZKqpCZ7Po8AFO0XKcZsZ+rMiFVtZiKL+UuQjvZq/5V4CbR4PTGK53K8
lgfhPfUAzicAm/SedpVc4hkOP12aj4NCvKuCfdOC3CcfnalJc064nd7F/DxwCrga
byipz7G8vL4sFDtWzeneHuhS/pxpkM9UxLd4KL35pe8tedCI2gLBP5xtzMk52yiv
5mVoaRGjzA2Oz+djU+bVQ45AEUiapnbIZ7dzKGU8Xybw57hRE362WPf5/Bt/fzD3
Sv23UvqhwbQWu5YHGmU1zqIQuKavicYLy3s7dhBOOONC+RZ6+jUNsEpe7x88pgoT
h2MZUj277yTZzM0OEEA4WmFIADZj/99TWXcVXoj3xlwMaXG/Hkb2ZgAyzXEBdhCV
IoPa1ApgnK7uHTjlta4II1kojol9dnHt5xemsJwdtEHdiPgR6ZM2i5pw8XE1x5LU
Pi9FMAyEhifD+wRzhhnAK3fWYtuSZLQvpzJnMuzXfDDdl2fbCSuqoqbwdELzOq8b
IGZQkJA9kxlyW9p27Q9sGZWYV1eHYmhg6i6frZyD+ZTjiCh4cFIkRO+N3444PaU0
qzbqFRliCBQbfNIo387Otb8lI64qcB/8cAicY/SWusfjZoNhYCnJ7Nk2H+z8NvrN
XBSuBminGaZLhO3C4HgFxG/F4+TAXYhOd+Nitp0m7UVe3XYngiflLZmNQym5+UFz
Q1tQ0DBGvjQkQJZPLgo4JuhAsuy7sBti9TEa7WbrGN7uDR7jfgsup7B8xSrmsQS0
gqiHlHNfjUmOD8QmtjXl99leWQCIVyGI8V0hX74NYvLDaXB99Sd53kmjbEO8couD
CscmI+/KGZC3P788cq49IHR/YUZ6EuosYILUw/8p7ufzxzKIsJGujKZkwTbwclQl
xpda703ROuaXucLv518JgMd2jl0U9/WIRjBEibz9SNiY5jo5Qe1rAkbEcuJGCge5
4XJhbGxnPKPPyz1c3xyuv8+PTyvxHEwRqdNZzj+jXZV9OKBW5OOdj8+LNYjDoL8d
zXsLpQnTXRZsGxXpb7WyB9tTkf06x+P15PY5HTMl9tN3TfAl7Kl4fYT8SP/ACLQj
hCIokt9pXGZsYIMOgdkv4tDg+UDZoE4u9CnUkz/1hq/abhPzCEL+iqiOj+i6apSI
hkP+qP/ap+tig52TNoutAvEj7TIvNNaVnkzd8t1nOIRahzqPAO65VMuNqmlvuWBy
MvACmLQTOjDx/GY/A8D0k82u7FiklGnFWDPOMkO9HsvjTmlC+of1mls7l2gOmrm1
U5nF4XRpuQin3DweOGonmBV8OM3s62dv+PohGTQa4YNO8usq2XIHiVTB2NDjDZna
DjTINYiEEe+Z9ksBuvpyUHpKYZVzaLpxjEQobKyFd6pbG0L4FdyMMmhgWJBB7TE3
hFlLWtH9Uz1KFWmab7mAorA7ZJODRCdrH6xLL2JeXDVz0QFjfk2rOZv1oYFB8kS6
daoWTh3E6W+lQXC8w3p9j3xnE8FFVQw6bFfbEgkL9B60UPPPlBNBoJctyftTJijy
5CMXTDq/98pHs70gSaH9xR5EC61wRBQyP4v24VS0vQ7gATwnR2yOQM92EuKlhZae
1rI6MoOmvve19Wl7sa1RDATLfCmLG3hUywrQWJT/TEtBcSo4gwGE++/OM0tym44u
0SghnCZPwr77/ntSGfSeBe/jRmSAzNiGinQ0/bbY8zz+BnGiyppXeIIiUYbGJzHw
OvP9FhvMkbQ1hu/m4Lnl9LOl9FzbcDyFAXfqulvRcGISwgSIIugTMB8inPwMkuCH
FjsTESdyIyCY2tRItTs2aUyrF8r0H+cOZwMS3BEpUUw7PKuo0rQkeJSD4YJ76CjB
b1xhV50B45TPmvIR/Zn8ZpRX4K6f8nuEKeJTDTorfFzz9gTBdjLXny+v+SUO5req
cwHKvj402ksdElo4YoXHGa9lQTTwjpLFumhhSkBdemxPUJDYs4x0jE6rwsWVFf16
cfucwUTzhYzT12QEDmkmQVnYu8cZ5811He2+QESP8jMYLV5EaOKcZ1qaQkuAYQzn
PhaJ6P5lR3ip6r8HRavLwRL7dj7ATo8jZx/1HkhV8+ny6DqPgUcFYgrHXyNEeE4o
i2pB3DomsAsPttlxxvvLKH2uEspW6rZwJF5w8nkwGBRCD0/GWy7hsu9HMKsGKDfc
i37EF44bMKzsPVTwA80fi8U5ZMfvD9ttiT4MxjR5R1R0vPLSMOGfNYvOOMIBCocK
2NnXrFJCE2fsoNDEft/RWkGpDPKdJ2TNon/2Rxlzz53+P/vzkxzpz5Dvc+1aiFmi
pxoNGS968zikDUuoimphEpP5KmWg7QZOSPaAPo6vaXSa2x53pl4GQMubKVP1W5lO
D2Wj+bFWPye3FYSiqyfQLO/oo/W1lPnOUprjDp6Dq8YqgnsORotO8EkqVy1RSBmp
Di74yOcfa8Y7VVpsuy/btemA5IwQ/837kwgqVYwQE1ivBZX2ZXVp4SP49Ff1edYF
1WG04ssYXxV8TQCFFmkdTFMin3G0tHpEWvrNX/9T9FBqwAC2i75NaC8MNLUM87dF
MXn7YWQQYmYeInAsg4TEoxVQwGsWc1pkCM/kNr5M8V3I76KmBMD2XVHbPX3ALug1
gxUVu/amUMObVyabbYO/kTJq2mciYmnAdipb3ZAKy8MYzHFhQchovyeHiryKRrEm
DlszzYscaXbV63zbVklUmpaneDtgzX6aop1jnjMc2fUb0w89e+xjNFXtJqo61FCp
spzyOgMLiNzvd7+4qiQuxT66JIn47H/8sXLTwp7NqwBYtU8xOlGs/ZCve95rK/4T
uvDM4tU415utOBlL8Gm1/F3/Xs7GzFmFXH/NAwnlnEkjjma8/HGmdsv7KYQ1aCXF
2SubpLFQ6NhnZAyBqgtLYBOh+bG659JvGd9vYYbkLfTcHKOJ5qkD0TIaX+/FfDvU
m8RWkzaoK6QB/p4Vpbx+9E9md/0Oz3T2fLrw3FNfxqOUB+rxP5hUtlJKlsMlfrTJ
9Kz9RU5FRvEKgzr5osMZUuozLyW/GMsPebH1Ct/W+Oq2TMFp6sXAfXNygCOOywH+
rvFapPr4nb6J88gXq2UunwvbXqc1oY1FTf/bEYwq12KmQZcsg9ft9tRWPANHLOzi
XOOl2CWFLp1yN5Mb7hUFkyqC75jPNPMc4I1KEQyd63rp2+XuyHQbVuxoamzHw5lT
JEC0VOULeAmSG70onoekUMuwGeBX1pMSgP5qEmsyqCi5zSlgoGsMxWNAIpFUu7PI
uifPdTKMbbq9t4tDxbvzFssWVGR6rKLhVTxE80SVAsFjL+Lfq/foEIANLrJ1WJgF
mfX+kBrv58pRExq6uK3N4J2HDrgQBTpSufhEnsaEAN4VWzyqVVSZ3xzkkV3FdrP9
5ct2N4S8o9PqfawF4TGlrk6KemZsg9S4vTaQVkU3oxvltXb29h5x3CkL3eszm2/k
U0VWkDgVHsXFlzLg2vhIjTWn1aXzKA00P6Opj7vC9lA1QchCJE8BlTs/mrWX7wza
nsVHRKyYiHlCloI53J8NJ792v09jFrb9cxDGfXsTKrBNfNTNjSpMxJuVBUyRN3Uf
WFzx/91Rsl1nW5P/4JKhqj6/HQhNJxCnHi6zs3bDG9hWYIC7+c73aaIz/EOhge4d
B0LbfOlV18NW6onRxRcZOdeDQMSZh66BdgArUCwAo5h0Ukqk7i2orbulVBXTex4T
8xto+aDuYUBYbY5/Uy+bk6KEfl1kBSSwfCUCLM+dL8K02kr+NnDbRQuSIXMnOAEv
4zjEcevx6QiIvM7HRP5KLGA0zSZ6Fi7qaRpUQdwNnnQjt5nMO7t0updZ+quKxVvu
7VKGm4eMAAvLRDOHkiyteEEQOB/TMqzUioaVTLNUzjVLm4mYMDhMm5MNLUa/TeyG
w7xaXiFF2gIqn4DrlQoF71N0WBPd+vfTKPjyKoOn30l+IyA+QdwY6h+YFTNJExZS
oStVTiWOfeRNknXVgAYVcStCt5t0jZvvAB30ZhohODEZmPMYN0/J8T+vBiom8PKX
KmeFbCwLtQncIZY/joOxeWeDkR/4VXR5i3bbQEuXNvuNkSrN/djbvLtUBkfDotZ2
DFP/2EcQYtfnuRli5Zrku7a5ZGm9Wm4s8IUcrfbCOsaDnIqoOFQVpppdNv9+xYVs
r6K3jX/lgDKjGMUlDhAiy0FyXo+H4lOBvf+6KnP/oulC0FQeRpwdBLZXAfjSxd/o
0zVNTDX/ayH/bWXsy6bbA4ljRjvc9mn+ACsyULDSbQ4pWW3AEeoAIKCs24SlHOT/
UUGlVVFtiSm+EX8K8Akyeq5xOyn4G18SCQVgjrdSGxB8+/Mz/DDxO9dNmRByPUup
onNubetLhR6KSSh2NCIz601CVQBYZP89PzdvEJMhoqficbFUOtTuL3SEp5GJ+BFk
6XWKq9HKF86IV1LkBeOLjipXBWHt8nOGmW1zuhi1FQKAlT/2Mvp1xDa7Yq074vMi
cyvWPEAE3ZcDtF+Dan182yT+eK54pMu412DwTEUrjKO0xPSZYimql3VnA6LBKw1P
UKz2yockJtKUZ/7+ruBRsDwzyGp3iuf9fEqT/8z2+mcoQRQBEJfPNv+ACCzh7g6x
42jblbeympLbHiwx7ynq8DFUZcYqc/zyRL90hF97x1O+yEZ2yHze5gJ/Uxc+9lwo
9y4iAzzC6bA8ITOiWs79GchmRYmegm+muxH3KVnH+a7Le996lz6xkLDY3zasKOTh
wftxqa9b90pge1aPXUGZRrZO5oAy3rfpzRFvgh5vplEo76SgpkS5Ybq/BIDlMhYK
TMXtaar7PzqZhgTgwYdw28S9S2poXe8eEhHZdfY5xqpv4c/yx15OHWBY94NwiBCZ
+Z4rlEfPF8DEibVhsfEJlSUkKdRh4QokYVw8xEDsrDuYRRSjMHhJ9rw6h7ZKjnp9
QDmAHhoQXONpiN2JpU0itZO6tfHN80CwrTDj1NXWiR/O3874HnuoTNoqE8HdUX5C
+PZpI9c6MZEx8qP1RvFzGcTMPTZvpL76vOWlDL8UpML6nUxghsETxagU4CVT5sM9
AQqfhgpgErkFHRgCPZdjihr5y6VzfgPe2oQawO4RKUbZCBbVrSOa8oWqQzXHlkbj
KC8B2wv1CS2bBudIC9p4BIaxUcwrNWqZED90RbEkI2P71FApDVIq+mF0OuSUqEiZ
6kL7rsYjRTYYvPaIwFHmfGTiuagEvLPm0bfo2K+Nkecj7faIu0gN0YY9QM/81G5w
OVA7ChqcztJaw6bwKskm2xTnIOkUyZGGtkUDtTpQOlYNmbdhr7ZsPW2BuesGY3nD
hKv62ycycbBVH6nA9XUy9hglcLFdp0/dTIKFcJbKhN17BhesVgq8XcaNYxK21ur+
QCC50N1r0lpgLNM8OXgSq+Gn13KA53MRnzV+dhw1i9rBGmhAJj21zwNzRKFNULEy
CdsIuK0ypyhclGowWHgMyMWl+vsc28wbfRQwOe7OfqVFpWX6Pr0qE0i8vawxnbN+
A5cCt6LUxd8UsJRg+MWZcD7NdBr+j7uSwhszCN0rPfjRQ4ohORo9mU90fOglDl8X
kudfZRz8DviIz5oR/+STDtam9V8WxQRV9c+tR3U7I3mq4hWsQLOiSAvMJJOoJCYD
6iknQdqJxhiQannIhyM8u8g3dbqbNaMMohJJx5hBWgyDr/x4fH+v12o7ooQD8m6v
OHoEFzX2bE2ES+bQkskIXsXZleJS1uLkzW1Gb4wriRETRGcknI7uiynDz6g8iRPe
hLNBm0X7UjFalle1i1ce9yJT9Im4ancEp7lFevO/wTOqemgXQ/pvtirgEIORAtXb
hfQa6HuhJT8WmwkWdHiQBhQCVHY+jCvZ+adwCvABGAqzNvJwuYH2dy/MXtf9Wgy+
+2sK4FNX1kmdKFfFLRp1g1R2ObYYdtKqaFHa7Nl9ZBrWOFYjRhlSJpkqaayKzdlv
4K61G720DeUvXTerhpJ6n5QcRO5Od782S4fYIgjmLiOe8YV5abvgl1b7GyHIN5vn
hKzlxgYGj8JeoadYW0WfKQfP53nzEDylR74UX8Gdf1gE7ijz5XWVutIPasjdhXhb
BD57QaP6I0+xyZ3VUOkAsN8M5D8p4FCR2wO5WF0v5FmXpRH3dxDLP3iV7YJ5hJa3
jAa04IF6ND8WZPgK5HTZ2gCLgF5ebxZi8AF4HHAaj7IhvTOpjQHTFdmGWsBA9yFz
OL6YXAODB6nOgOev7Jk35OPDTwdYg4Xxw3SdC4gQEFn+QQC83XiSSc1ErmCvn0w6
WfadWyTpaAPKLRX02ZNsuYIOEUGrtCVhUPamIcxWrPi+TMsqNphlvR539Pql+eCi
kP/40gT53BMcXSl1KkQ88cDt5ixUsMgNRC08Owbd7/A029UQdZh3Rt92Q+PqLeB4
trVU83CGq63NLiGr40pgJZKt2xitgbHFGl2PnX+c9zteWLwVchm2B7e8QLZvPCd8
M4hTAu1L6ZsLMp1i/jL6OLRDaohBZ+N8JhL5GWIdz400CB0tWOGCiXd8Y9r6kkJ/
d97kJNKWP4+1pnSE5gZ/45slpSHgSlxIUWnqnurKNEuiNlFnrK+2SlIUWH3un3eP
V5Hzq65pII0DYaezcnhm6mEXWJ+7bvJ6y3EH9ramDK0WWt1+gplULEdXvMiLG/CG
+dKMxtpS8UwoyKFQF4glKsmNU8oh3M3kP2yLEMxmhKw3TB9iAIP6OjvVljbeCrHn
OMTXlA2saL+McMInVWXbs/jfDOn2NzJr5Uq04Pm/HAtMrwquInMMFrAZPm8iIJyD
JmA0/ixGgFCVBMN4OubBVUBOl2W0x/ddoDdGD8HisDFVpZL0KnsC8nQe0J3jBTgw
Ri3moN86np6bcccdJhhK7OOkoO8L5StM56incQOR//9tY+fWqYCOGwPLT6BHUUCC
4fL0PCqBYqRwykbTFFEfPq7dzxB499eA/prrqT1sijxOJAfprXjyyO9QmYw/YNkO
UuzAfP607BL+b35xNzMg2ywQHAGCbv/zbMurvA9l9s4GQRT8JTrvUAwdabMLytU9
KoFdPC3FCF1n5vQjqkBqMWMJeYqzOzujXG7F/jhWupdCP++rTRuFywBaHXkEbpKs
TUZkqY4omox8yzk/HLXMc+y80sazwIzFojNm87AXnQPjHsWPv8qHep/6s5Qpf2aM
KfWssKLK2yJFAfxzmTxKUXNo8QU5RGSRE9LgNiGZ1Sb5A2CZR8AWoumD+h0Gsjmy
ntDFt+izhHtPJfgy/W11S50xwtiYHDvtBZRKKSdBQFwKzROMyuu+o4AwD0ZF2wQ4
xp0BjP9VS55kuCph0ZtpgMvNyFv5qBgPEw3B/4TAOSI6m77tdNNfXxq2/huz6WDf
n2ViHHNHHU0hQKssStvfoVqQ7Q+DM/HrnFV7rKjS5u6N0GyRCpM5cvm2idKEy8fp
MaSsuEZf5yo9gUIGA0KB5hF9cdg3INdLzDgOgDWeKCehTLAjwT7lnnCjRPOeBA5G
PmE6hQUw7/LYDl6W+OTkVO29aKnBbVxAzbYAaPdxe0Z7EP00hEYW0C8Ff6YqxrW8
LO5+mO0Um69MIwfsuN12iWJwpzf++51Kdxo9Y95m9KG9RE264xxGegiiCTb35vrD
KVyA/MkaBsd1kbcN9SbMQIOmwnuYM/eXoN8dBnSqOIQ1c1RYCsg4REae9OXmI4Ok
1z8uI9gap4yb7VFVJIRVbmeXJKDJA/anm91gwm0fgVxLcbhP/BoHMlSweAxX79Kq
LeDHVvkFRgPlmIgVNq3rjahteuPL66mNgZiNVIaZ1COyqyFT21JQ2n9j3cfwQhqJ
m4NgmFlHPaGtgTuu1nK7BSc3kztXXQyA4/xWgjiOCOduBDcYzwawP6STOPz7B37+
/NQTUTMGr0UaF16IxlL8MsFR1FRWzFUFtW5+y06ZA1+gVOASsXskSCxcPxm36j7S
mlbIR0Se5Z5lWJEfk1zCQE1matsolOFb5s04SohjBTsOOw/Ew5v79hxqHl7VmyU3
8Iz59t+zUTv7VfnsYcsmAScI4JMqi6q5f8Vj2s84/cYPHU2YSTb2lPoABmZOE0Iu
fGQXBrpv6wMCMOqM24Q0XkJf4VZozj6r89Q4X8WApN9NjfTfS+mkLEyoSpUx45pP
gNtAGHjyah98lD9gegMmjU3BALWx8IL3m3jF950oit1GuY9r0OCbPgGlWzRjoXPJ
6YXFxcsgQVlPGcgAGOYwLyc6WXzl5CU5XjNMJV+Da4HkIoZIV2y8K49fI6yIw4LZ
PFn4GESEfYi0DG6yCH/mUZkqFyifxtmj+JCCYG3aBL9ZFwoFKImdbZiYBNMdWykE
lGa7aGojXyn8eCSfozywY2p1akSsBOUaYArtzmT1o5+5WImkl743J8kiFhj1yhJi
JvZ4puGb4IypYPRGJ2HrZN03uLVZ8NcKEZcCo6mtVHIt0r2JCcUYA1TK7HWxzp7u
iTVHyDSfvPDIfMcsYoygAl4G5rrhJKJBU0Im7kOyv28K7u5g4XXOBYtWD0Sz/DGG
nZFg/E5aFav/vp63BvZ7YQNmx7Gk036qCKFUckyYtvyLZEM5aWmEOYt5wHRDy7M4
T62pwrIC88rIbhQiRNbc0kkqdPSPQw1qkwYm9Z5DBvBxuQbC2z93n1FU9T+ZC2oT
Ks3O5MId4f1F7SmJ74T+48C+C3gblWnox8JkRI4DqCNvZuIzCoKXzJ91BcNJeFit
dyBBVCzlzYvXzjB4dxj/DzpprPPcdiAZtdTPOAnmkgyTP8QTFuTg/tVTGs7UzT4J
87KZ1mzPn0tdnQU4BfFxKoq+7WmCuN0WR1JiHpQ3+7OChBxJktunlXEv3gzdIMNR
eydwbZdbm+/BfBHb7YLL7+ZMghzdGPWELOuUAib7TFInmS074iP4R0AtRfFEsX6P
kU0MjPW+X9VSaeN9stUF13/VfmMOlF0LR0zScv3f/oaMC6OPUSut/dSo2eJceqZB
9xNZ4yqWr13NzKgcxqzTPPbHq7n/0K+CYbH0eHaOVJwBecrG98q67jlyzuGR6kJB
zsfkXltu1iMrZMu9owDRtTap4FopOSW5yNuDpBhkE158k0JpUBV4Ip6G7OEB4Sgw
G/93cohFvvgqOS7WgplfpPZguBQB1wCYdW3KYO5+RlhcIXWCOBLiaHFYW8fhYW/b
UXW5m2deSIqRKpeDMxP6FGCppIuV6nQBKVW8RXvGOyygRtfBY4o8C8oBwhHXXjM1
te64kiq30tEzg0EbVdKRM6sz9z5CNJnutHCnj01lOO1XvPjP8JRJcP6eVo1z+WDx
KaAEIJoJRw1EXuFtqdsKkWHuslTLCiFB6sonSLQBM6b2ZAZOPQfglQ+CFIPApvb5
hT4XFea6TSRtp+5HJHhRJ4MUE8o/4bOFurD5pJ1i/G3vyZfL9Ne8r5SexTsQP48O
wXi6KRwvmQnyZ4faH56WAvuoWtTRphvHJMUWk7ACWqhlNl+FVa6jU8GdBbChFqT/
vcICEqALD73C12HpsD3M01b4wWsvRsTGPgOzspPCJFfSXR95XCw3EHy0sAK9ZeoN
qRpzRNXARK2JsIzYew0ov993hK0yDn1xc8VukNmxvmS3WA0FvZnEFby9zNmz6uZ5
jgAHkJQ1yU/JIh23iTkJjhWKCddacNmbJosf/rKN2e5L1aXwe6S44FUqEQ3/Jblk
30sn9ahffwR5FqZkgYkzhI/3jwrEM+/x91bULsmUbeiZ8XmY93qC/LpM5sb2G26V
EKZrnQnvo5rgkO5rUHZ04zQgQVzVrruqmUYq5PFQ6oqoaXtgv2oX+uB6GO5QXwy9
q857cIgUpjrg7KWyND/btyFf4zASOCv4h5SeNhFX2OtB2FXX2/7Dynua1OAv+BSO
es8KcLlKncfF9C3lkoIixZwKEQ+qH1tdNpvUaAis6z0aRnVMH9NZok/WA4o8+6yh
fAZ9v+uAgphLTYrXXFO1vL1VSG4ea5czJK6GnysIBEdd31l/FUiZU5eyoKoFbMR1
IV6qQ3yPJzvHmMh0BtyDiPQfDAPhhUZ6u9eBFyGMNoQpcYpKNZn1OJJ7tgclfMrq
os10A3KL410KpZx+rECE9wvHIJjQu7+aEZQDOFdvzcJjirpzzrf0SMRWU7kihBV9
wwneT5voYh3sGa0qLqeeItempPC5kuvfx2Ylafrj0RTEQKccdGjO+68yVTszIa1C
58xrDa+8uF7psVYsq5Wdi2RFlt/ZmOuDI3kAIwcbiewLohfhfMQJx4umYp20x+ib
TW5ORSgVP+wI8pQv/x3yK1hnFiqBqlNZEVUSbkCf6KQGxeUV1Hdo2dgmIjWFr462
HanJYG+Tv2pcryyOg2hemxn+TznFIxAxLdaTv04Je5vgW//AkjYkf98WcA8+ZRxJ
BGb9gPWFbRiUFHl6Q8qWqxMANRmr70ObCkmDlxdBpPzwxsJFv4B8TEiFjQSsKXdM
3h6cCB1KajxT/pVca6KAtsReSKaUO1gX6xr8kOiCQb9y++04M87hKrxLY/7Mxbtw
7sMvFbi8bneMVuBd8/DbKvORL4gMQwJ+XfReaBeZoQKn6v3p/5aCUrwRe8mPCRwq
YnfUaKlQvIsJ2olQ4U5eZzR+5pVNx54HAdgyyHGzzupNoFeFRZvQQTLWumKbYwAr
md6avzIgiGfapICDLG0eUTtaduLHQ962AKnMiEuCVC4Y/+U1+q0JSs3iggDwa3s7
tCVgExK4GZvVdeqnwVkmqIu3QEt8bYvG9LLfo5K05Li6ILc9GolILWklDM9jUXrg
kxYzGba6meGIF06J3Id/lLMYLFoUiF8PhwYUcDQ3f0LgotoeSXoiSxN50HvSJBSi
YVBWcKckBqqpAjvCEIKfJjZVJf1xMvlE7rlp43J+rNI+rXdNFtkOaHwYCFw9uOxA
0Pe4oALj+BdOwwqR9IM5s1/1PjfJnz6NHfZi570WqbOHN6uSc8qe+fkc+MH8Zztm
FHZP/dDIAlDziUuAXYp19NcFJChf+dWYtZaXGT8hiRUBrSPW3tikFx6YyGyqzvAl
mj+wbY/DKdesYhegCH1MuNGqLTF3ZnmpETXsdxkwpvFI92MIpfrSAx6Hc7SsZOyb
tis1Q1fy5GuT5SHv7xhxyDn21TXlfaSFCCZujSU42EZUItfNTb2WSGTTi+h2gy8I
mos03VeV5McuZ7LaCL5KVIo9itXeKckofthfSqvwpvIt+d/SylgVJPUHV4JBF2Hg
/JLx3LZ/Tin3LjruYv9g8VG4sgKvg0QvtVwmzHpt81YNvnw2l7xsoH7fP/739Db7
nEF5kVKHj2r1OHki+Lzje21SHHLODy0rwEhk1JL42TJpnOuqnL7rtqJPYEvnABmU
gHrfsx+PxWte95Pejhhd/ipD0hWFs8rdyveIKORINLlcJ9c1Uu7bkJXGjSzAE5cQ
QhNXuJShoaUTIM6cMCluxzojdU9gWPlggKREGcqPE9itIR+C6dGAWJwieWKkCAtF
gjUKGgCgZjBFQfOxP4FC5e+vjNtoINIcgEZGB19zZ2Of0v4GJ8pHte1q7qW60I75
/MvHAOX5Y1ygdwWCcz4cSMTZI6VZKovV+UlEJpSqX6kY2sxShU7DXoK3uPNz521S
fPmJDG8UmHtc03faX1HqGaO6obnpg+jLz26Qn+5dWtdnaPwg2SiHJJacZNmcXqNx
IXsrADXdADf3qJi6FOGKQGnriwB4R1DIL71RH806f0bc5E9zlF4am31w9rDV97kU
dSTX/XBfS+UC2sslI6P+KW6UMlO+Y+AeHThF37Z+7pkGCUWkIvZjz8EcI5o9zm6J
3YEPVd/JxT2j5wGYkvYfMsq6k2dWK6YM7nLlfglyBuFu103e/JeCV5Fb54Kl19Yt
7GF6jncc9BF321B6JpYkK3fPr/lN1mrycO4GTq/IEpFxciGV9Ug9/FLunAoP4z+Q
A0g9pdeC0noDq4BIO0sB1OMwGxMjC4b+C6l11sBBFeJ7nGEtbcggyJW1/Lbmk4pf
7xXhQ1zo2SIytvJ3Ja3b7R8aZ7/jkLGnWXLY4b91RkO01p0evzOa29b7ajkJ+yW0
wsUZTGBGVpiI47+52HeJ4U6iCEdZpnA20YlRvvsS3+967okwq9xhnSuQQ/Hza+nO
4AOPp0jm10Qd6JwQhyxJ8/UuRoaK5eW588tDa7VUhdN1NnL/OCSEZQrYxX2tLkZq
JE6OPkZqobnQ+3UeBf+Q4fOfkInHKraTZHyfaGCc9JeUKeVUe/hLQM2KlIBONbS3
zi7s8H341G5qKB/OKxM20RD78OkiFxu25VgETmJpJS7LYL/XN+UuK/J8UkaHEWDO
F3xkCAYo4gi5e/eipUbCR22kW5BJzrLYdP0I8wyZwvWPjrr5YhwRo9Rb6qxQvgVu
I089q2mgbQxUt13kvNC1fhWfKrGnUeeRtY7I7TaEOLdJhlOGzL9DFc5lsagE4+7J
vON17fukgYSo5EHuhM+hQ9uGVEekNDP7Fk2lywURiBXd/AX8Olr3FZ7BflPaZzEQ
Pz2bV0RC3UYxyFeZ3M/CC2U5tYZvXe08UxSJbJrQ6NqqhjCMR1iaL6azRXLgDeP5
RjlBQeWOGhQQoWNY6IIyYaQ1PZn7jZmmnj5/a480hP06ee5hhpAXkZ95nj9FkvBH
msKRyKKMzTJ/w7uo+7IheEk99nNaa4cbBUYlEyxsY1rgzWamtJOWlPNQ2Y9y3Fdg
wmGzXzfDp2Y0llmoalwpHeJZzaZbktMGGGfigwpTAr+D9/eXPHBq9D3Vpjke0Foy
1xR86aKxzpy8P0hRZVQJ3BYbZTfInNge9O5Qx/HMEjCgUvlhZkkT5c8kLe/fT89t
oRuiANz+S2KGk5WExqazyEKX0zqfpiqxS6dot2H699dznmWlMo3ysRY/C/KaTGoa
VcsSWAU6DZfgXG2IxacOqWCKkIjqSf0axSj3rg6XN72ccpRVKn4/lnMjaH1J12oy
MKwnK8O6AwrJxkwJN9Um9DEE6zSgfv4TYAnm3osi7NYLUuVf4bZ67fKX8EaVvulE
rcBlB00IX58c4vqKK5EqOxDITc3ZQxmQBhVhcx3/1sU6vSZLS+iTQ0aMSDpBk/PB
Og4ifflGGsJ8F37QTd65uon2vWr+xtnGF5yf56VVb+ERL0Yg5BIGP3EfAh61j38r
jQ3vVy4Q0QsUzogMKUxOWnWh2g0Vbh9g7R22k/UbDU91YjqIJ6VxnSL7+f3G8q3x
xC+/NGfRTL8yq9b+mKKt5Qs6kYQaiiPFr1JAOz6uN1/3l+s7ok0MMWT9trA6Z1PZ
SyGgseVArsHvMPhTxdzosWilIUcDxz/fvCyfP4I+E5KvWvDlTMXu5ti+FqThheLd
4NstODUrX3NDaXm50Hhzaqw2gurxCr9nrYeCpRTcxYgwJfcD/bI9oO08SnhGy/9m
RcKWjd9Vwwje5nJ0mUykRnGpykfDwTQLQz5LuuF7o/cLqvGXCfgQXmvcPqFu5oA4
EzhTU/+0luq6RSAPwHqOFn+LUDkusQ3xu9WC5SgQJRgufHx7tCCQT+IFlFO5c00B
ti88skJ1CansRGi2v2JvYGydIqQrqZS4y8fXnWgHR8vBisu9607hrzjlE6JKWLgV
AzPtY4Szb9mZCMDXzz47uKF2J+T118QuJi/9MAq915na//jkx6McyGwXWIYS6oWS
4BW/xkZmwBJtEjGrCozRLrQ5JQ55UUj8R+Lf5V7kAnyGld9Ron0BG/1O/IBPLCG1
G71DRW3JmmUBm6mGt4Ta379saTT2fp4SyFY1/Vsc1IICOl7bzruzFtvvoWTUVw+K
hF/wV7Ovmz504PvY7JVljTJz7AouImEqN96tX25/Z5bu5eBXnqhWlWzhcC9WMrT9
Dk0BLH18vXacna/v646KLiNXIqnY9xJe/pyi1RG1NNcOABCsA6ZxnClkMHsTAmbp
MklNT3lBsQrjZ9I10+LInrTr0D6oWuwS9fcTeEM5dSKC6dCd0DoMxDkl3FLUVkz3
6qUY3DZyNngRXs/f/F4NRnuCe7amT1m7m05kREgdMvN5G85gvN14Il0Twpr+8wZ3
lG99JNAx9h34IV5veNcQehqblHiz86eS8tNnjyQemhuRHQiwEVh8XiJlR/fLEGZk
JJT6jQrgKZA6inTYuArNAJj3Wm9f2FOdycujiO1VZXEj8zPonpIB8MX0y9spOXjn
Hye7Iki4E/lBCrYDM0vHNjzHN8GDCM52+unXoK28T1A1RPyBJW+mNgoOel1aVR+/
6SiZBuBfUY8WWcjOhk5rL9ZsrN+HpyYxR2WoxsViWTYO7ZN9jim/9Kbp8cUD1IJ8
lwvScyIbW+hrsmRc6qIuHl6RJNEaUe/W6DtKlfS+0bomWsu1IkoSlplIN1MtCkQX
8J2VwFFy8NZEuVocZYZbe8KkgaP66N+ip7Qy4zx5y5lX5+VXIEvcPtgelhA7Auce
aNRYEP/7OnURDUjn3MhVgLmi+yMr4IulxiF2RMtw+StPGPBLzoCR6fVhIy+GTzKj
i8OShjrf1wwTG4qWUv98J4JHG0CQiOLt3v/fiTeK0RhOjHU78zhZjkMKKlrIXK0p
nai0mWgq7TWsa9xqQq5JpO4vXzKzRXHDjp8cVWzNA8FA8vrtUIRONwdiuSN53S+4
ObWBMIM+MB8Hpwd6D9jMBOiKJLFGvJE1Wh21YCrmuhP5g0qYoZaMdIbARow3lch3
J/XR2PX0R6MVdlZAmlTm9k13oiUf6CZwP1Lf49M1YO28IdAaDKFXulqnC4Jh6Ukx
8XxslUb1EXIucd+PXG94VwaZjJ5tID1IECH8y7bF1B8ZQB+Jeyk3rU1sXuVhCSlC
UUpxd9Q8jmP7Gy2yxjcn3AY+EXvWXkaWhfLnzrhG3YKsbiemVVRqMb/Zehomwb+0
WD5rgl9mrklz0XeIuZt+oOpArqgZV8Dz2md7yI82enqKVxIAQuB0k92lIfA2TL1T
a24t5M5ozR2YCXbZo0xQ1smY+Vq3xtV72mzd/Q9cva4y6HC6yYb3gHlXI+9r6Gt+
b0P5Q42RkADt3cbtMQLftdKv2qU90eLx42ehyAESfranILzGjATsEZe+rx5EgQqS
YMkEdwsJIJeEHBFdwfB+u2wQuK5XmGjg+J/gTDHsqoT+1UOgyFk58xMWmBlSHeDo
iNfCgxbAheb3rir9+RIBsZNJES9XTl2Hr5lMvDPFL51Y2GxY2oEGmnGjAiGS7OVI
UuMioOqrLzRoBCQg7LVzpIiCNdC0BoL1GpcW2tU6D8NWP0iJP1DD/XiKlHHPjIiy
FomZxz1x1XIRRP1CtE1yi+tp3ZX7OtXW2jk4+oHTc87iNeiYdt1MTGcOlsTNpfYO
XkvbxUIala3uSV7W0639eQ5VjGuBrH4lvmuN/1/IoYMTPvDb1e0G80K1NId3zOFx
7nQUn7AO3EbLxYui5rKZ3AC8TDffM73P7lnLjl6HSYSPEh7zQKwnsM7nsFUHy/cy
lX289tY32JYCjLaLYjUNtZ8kKt1i0WP3BpHrUeyPP+ZfCIicgaAkzn6fL1IBt7Ut
8jwtWUwV5Ix94Ag5ybqCysbdOvLWZGtb9zuBn8GNM1RJH6q6UUO1iznxI5HAuxue
N2HsNaiCCMbkhbEYOWMwLMWAn8PVqXKyYsv7Xe/l2SB85W6aNqJR9ZIxcleDrxYm
SVR2xErsd748PHyFoGnNq+tHTGi/NdujGLnHXB1Fp0or3DAZlniH+mwdfYNgGXO2
CN9HNpYtQf4irq9V/Ur7FJX9yTmPqr0dXdHD/JZivvJa77LhgkJfIo1roY0QgHzX
aosz1WV9u1/jw6DF1xXkAXMjrqWvVJcteilmxBaiYKVWDMSiruAUs+KGIxO6Wc3P
ZRGrSHYeUrn+xVDrkTfd/RLEM0SlTI5aBTQfK8yBHsoItYEtas6gXE/rATL+pxeH
ZTg2iUfXfComosU5znEcUdeVirAcB953NlrDevrQtLdZJXPvvWavcaTEon8zwZoO
w6XsfTBJOYmj2a6Q/Kn14YXfNIkhmrkEVG0Z/KXR24arThZLNdES7X3eN4ZVnzSg
K8PqpVAmbw+MFUcs9ju9DbQLjY3YrOEsjuaosDS9BvK2+00vckpeng6BvQJ25HOK
YRrgH4MKqQJvykeIXyAKkKAcIKW1HEJo143AysiZmTFbz4SaSNOxPctUcsUcU34k
5fFNvD4N1rWXs4bZ9MBkwncwIbFqCX4f2/0yAZI0KksNECIMyzvHZbGy9+qGnCfq
tC1jIZBxF3S/7Dkbs1skzGHZNKhJi7zLK6qcENfDjvz0IVRt2whJzR2gt+QPvvgd
YAUKSRcXzQvivPM3Ku589DEe/GN+YQmeGMjuLPtsFNChgCOT9Rxux+RjaxvoNLBJ
47h4bMYXEGB45TC17i9WfVAxHdMdFZUfXwjocYmIEDTD4HoWdlAt8BISerJVPrN1
Fh0vLZg7qBnBThiQjJh44gDJG35rmYLOYU7/d0uJj82vMvI6ASP+/yNCXiaadoTF
hT4lsbX4Q6TfI1HZHnuWs2/FtXK3I5Z567p+wIvshROyp0iY5KOfA1SO3DnHJUQi
b4GeSpeDvtXhNNxdgFjOSGtLByxM8gmQD5JyS1AUkZ0saPK35opaVNCsyYnbNafH
aicNrPY31qfnvNNZV3gww51+AfXj5WgyMrbwMVK1wK3HhyZat9ZegHKULATX17Cm
2G5dX744ktF3Ql9nH11udpapzXSqkSj8gXMNNJQ3OAe4ryECvkwVefzfvm+1tmxb
UQ9sgFXbJM5wTtzQA8hHZdr74Q7YFiyj+lBnV08+h12q9Hd3wanwsuFKS0PcOtUY
uA9T/BM3kSMQtFNb7+hZh2g4DSFnmc/bhN3TBY2gYnND+hlultVHjsM9RcnrAzdq
lushorW9JGDM/+6koPjiwOaHnDs0RCKt6ydkXWEBaGiYwPm9LFwn8956J7CQcAiq
ODRp3XPOpyLh9gzgovAnLfsRcEr79FnzJJPX+xjxX2W5OFysAJsFJnkMB8oFjZqe
tTge0c3S8u6bley11pODIfBktBcMFXsgw379WDkECav6JSgPbSp10/xuslBpsDfO
B75yQHSuaqkDsFAx1yq9ADrOCSRIKqbyBFGPi8FLTZOd7OW3yZzHz++5kS6hIC5e
x3hdCpEMCriw/UZkf5Tx0eCf9XE3U7Wl8p4tdutJgfCgRJ6OQhz70exUamQyusrh
Om7UexOYlAtksz6i4L/vtVIKb6/UzWm9k90AGkbEkkBbEV/drqFo2dG4hM7KYwiw
mAnvoBDPAEcYKjNa0gt6MDNlmVEg6yzBozLcnEnYdSwDUOVNoA5/Rbmb4JV+/HS4
+SZUBrwwWGhxkgkYJMHlhzqROmDMXIA8phOT+pm0zZpskMEad2XaUkjKll1Xg+FW
GLa22BT38OBy9l0gwd7LyZubrGwqT9uN5hZc7qD0oMzkHV1wmstpDzdSZr+bXCpq
bpAn4ZP0KyH0ytQvkAZVOdlJ4GT+j3PtyrVjHFwUNx9rAZoXlRlj318rdeJzit6A
Cf3rhTQX+nNPkSNxzWyNDVvrD8GQWvM1klrebuRkTe7DHRyEywXzZMSl2PAoLdpA
nU2KL/Pfd0HH+RanDBXt66GgcmTli/mZBEyRucTz1yPXe+nJlLy8AST32b6XM+1k
MBXE2fQKOV33JULQaXfwdLeNItOYV3x9RR9Jajlh/Bqw8q9oUYfgMJvzmPgNYeWk
GybBcCurCSoXyZFda/O5Y4ITKEiCMVaF+YanUgYPylgH2wr7bCGquuMcVHG6Dtl3
Od8r0q83YClIsNd1mgJl4cieeal5u3kp2CnwWUVQgVRgTUBep8YLcE5mpBLDAOMN
0Y6096QTLKOFtE5Jvxezc0kHskOdM+dd5qQ6jKbLDFtZJnjDsyNt4oAgt4pd00MB
k9SXC2EaUFESyEq5RKMhy7GnmONAREho4j2gUq1Y6Q2P7+KLlziU08I5PLwvvj9j
H4XKN3D9SRQisM29ONEQcnPMOmmu5jNZu2u6PDqZ5OOsMHjwBVk261UuMaY7+iz6
MKdMjotPSVpBgiWxODz5Dv+O3SPozJEkqgnWYB4lZwVB1w1XW3TfVFDC/mjwKtz7
V4iY1PT+OCcaB0Nd77DM0SnL+x9+TrEMJ7907OG9tXDyVsVG9x4aN2SVCi0qArGj
dHv5zUqtmi5AufcCogUSsRdmBKrNXVzVCz+IZTJWJytbQzOw9AkLD1aN3y/H6K1m
OJhp7R1wBOMbWT5XiVOEs6KOC/hdO+cNFPTeOGGu6RWSKPJ2+mZLT+Pq6Nyf1BSX
V0PBfgCxGKgHG5zUifLFnhHXeZheAHJ5ShLspQSJ/QYvjT0oSyJAxmqcFqiqXuhW
fnLra+QMyAMAYhNwTz76gfD9002VLENNkqg/7cHlMyYSSFxOLefGMF1zMmcCPL3x
kPmDT7DO+OqGDLjjNVIUGC6yyFZ/6o3CmTE6aR9BFJnvhdUZsDeWYBShG2Vw3upu
PaMvfIAoLQOK5kAzph0pe5xLGPzP4C/7VBDYYPyXosDjSSGHVcdfMSa8oUpM/c0O
6hO42h8H6idTW+YDkKyyuocdRbWccKzEUAiUWfVoIF2H6kDjpW7UFbPv5wpxWKsw
B6M5kE/p7qIN1I28jlOB+F7mMrbt9CTSvt6hvcizSTQW4pAbnMoIXtOQO/mR457R
K/R25l8V5DQ3SNK2KS22vtWsuvVjEpa0+h/qRITPFtmoRV70GfBQ0uaPlILNhI9N
c3x6Ja+eh/TA+1NZqWE0qCfI6Z7PW5gRU6gNXKjdZL0cGP0abN1fVtwIifasWJ6H
5X/KD90VbgT+Geb+4sDhseyBH/S6DHt33U+8JYlTiW9eNw3J/oLDTN54zp3Y+nss
f36YHT385dBzk5OMAl/jkO/KVwJB5WItQnXdQGnRN3NGKXuhTLB9vHWGTMnNoNkn
VBqzuRQvq4OIbzmEAGcAkjImyoiAPwbC1DAMR5WMHchk/KppVDQamGkc6f5H/0S2
T6qvYJbJZ+ZFIkHSynGK5bJuxhu2NFBF9v5YmVrCuZ/Rt2tVQaDbUBotOEUw9HuB
Ea1BNQZjL9TWzjUCz35oSwvSPKqcq3kU8LecLL+OIMTpfAhD9rrzTIJAn2Ng74BU
jz9nTO4MJf97eCHbvQp5qbTz2oODDr4EbBS0pGfnS2FODO3XvrFX73soyynuUZxy
6de/Bdn1nmxsZqQIVgcJLZ6CPut7ijLMbWSLGmEZyUiGxGFFm2mE7U0S6DBd3lkt
BFJCGLUYyceBCk8FToYIW3vv+QHwXYxTWnAb9ZQDfMkwjc+MLuwgs81+ofmyeuUp
PDDGIi+I4Ls1TiUYAaQrJZX+kR0VdgjZWgmlohr53bO4hy/86jHBFHw15hp7llVq
2nOja2KIj3RLJe339tBAtq9x+iNpE7ABgYdjgONt97RYUD2nbXVQYtQ8/AzrtMNh
8kMVsUE/1MnpPaZCtLfh8M/T1hF97Ree/Y23SoWnIwpmsykGMXPwyFxkCyx7vlHV
A6SJ9QcK/VNPawznOrf8sd2z4V6UC0yi7snnFia24Z3+qFHPWvK3xK8R18m3r+I2
WYl2tyQWq/WaBbzdDGOBaHbMM6fLYDfzS4JSv3STuHwnhv92+5w1b+HVG/mJtkEY
h0RdRDI06iKAlpS2P3p7OSnH08GosWw9Eztk+mvC0L4ApwET2BU5PRUZY9Op8QVh
8E77YNqyJLCMRvhOOiREKr9qlHBUM+TUn2fMbyvT2DtSpPJiQ96GkOY4su1+xD2A
Wc0uqKEMZG+9/ktd93X47fGtDXVHgopVf6Olfsh8ztS3s9nk0hLm3+kry+ySp3AW
yJRGlVyyZeqhrRGnipXVOLsssFeSr/LM1WV/TnOfvwvkTgeoN8d0nbShpt94E9DZ
+Sd+UIuENqRRKEQZxUtvSh1zd6g75IuY89dXXQHbvPaQuJFElhAg+KbyXuh2+SwE
7N2KTmqgf9PI0tNSNQXeFD3QQCc7kSx/aJyiY3/npGSOmmCtAiwGw9oRUUWR9dcu
MmGWZJPSOSLmzttlaBeCKb24dpAUY9rBVt+4jBpLZh5UwYuMF3aroTiB4ZP2wqw7
z6XtR8ul0H7lK6nUyjNCJRBIKkX4+GbcoMV4EuObl0lBbtYXTDNagJpIVIzyD+3O
qPm4DkBV3GHXMqwlkwpdoJjf70TElqQ+InOw6C84sX4dhu4clpoRVacyLN87hAF8
Wx04IG3PBnpK9ATNylhMJPeQjT685tf20nAreWebSuAYklcmV7JIM5n63q/Dv1ji
VOaoPl0WcvcIJqagNp9z5NbpSmsYnPRNpnNfgbQLVxdiGsVzEFCa+UiUglkCoeve
9WvjzmEMwvwdD2/oJjQo6PZiep07jL8GNgG6fhwYFcLagxa35J/4CFounR7BHhUU
PKGttpfOGamIdiRgEENq0vfbVDOSkWhfFNreBJjhBwIgDcO7G9lYsMMOAKdUlikF
9jj3wI4VWbKC3IYogPg2/xdbvlRQ+xrvINPOP0bOnedU5lI2K3nRN+wMkGhQ9gWY
pcJQb5v8sdKkqmxPyyO5Ze5+ySQli8cTZo5OUOoqpKs0DtdiTDuSirDHqK/Eu4ut
lByfMY/HdJ9r3EBEMUK4WshnILlydumv0WASMmgwiwvk/TmNey04k/r1j1JeV73C
x2lhHy5Us1ZV3Jy4Up+TquXb0WzYs0c3MvGDBW4RryI4XxpitqJ3fOzADd9g/wAn
QPuzjx1AvnBLV3X/iR2TmTCt+Iu0xd2WLMHIKOubqWQlIuFgujA0MZRRfyKlmY/a
p/jFiW3Uo2nW0bNESC1HDhqeJLMmqomBUXqENgs5EIqdUzFMgQbWCm0eH6PZDTH3
EmJknU2UbsKlP+slrwonTSaqKEPTxuOUKEbU7kfxmVa59bwZ1rDllcZ/iZufcutT
46UopVkmaQJ1Tyv0oGU9F/We3prIClMyQAdHNGO4ZcRhZ9dERWaSnq2qMbiZR7yJ
vCByy36geCYBwPFzd1NGjDVWrVbQChKzE+p84rOLDNd8KC/kqLS8LQBwwGAHRhvf
jxth8YT20s0d/Yhn8I17K4hW/tVtE6b/ZuIg7Cx/KecAVXIEQrK3jGmrnR/fD1Tv
8c731hr8rJydsZzzJsBWyjJ+Ml5ZiOsDIx9v/nymeHD6rgYh4PaCxI0kHjk+jV0L
D3brllXzDuokzaz2J3CL3Ddb6QZNoqqxz7/U9V2FRTTemb64j9ahJfq4g7TVLFGt
+G70habLig6tlBrvhVLPLdXF7ySZ7k6cH7oO4JyxOuSpUMFFugRVjrHKmctHorzv
n4WAV9+FHt+DF0LEfVekHArGWwCsdy7gY9yoC16tLIwGpFKeiyIZudBpxQXFyc6e
SXUgR6+FspMSKmAI+ae45gqNqzYw/F7AcvcySCoqaf9RO20M4zXWGC9bjA4+sn8p
F98HAS8PPN/fxF9ITZCifStqBmH+hM7+ZsM9uYs+y2TR8enbPuCMlYIm5j5fRv2u
i5QSkeU1mG6/hOIDM9xOWvHhW5o/UnQememVbBzRDWStKZuL8Lfe1t5Cv3Vs+WT2
8ttjeXA81GwQVIX7+ubjTz5U7jWx59WF2LoVaot9QXGtLVboJYUuWCN02DUaa8rA
j+S7ChZoEvEQFBFApjpsqw/QL6SuFcMRL4lzSmOCsU58Nfyxznuw2E3l29qk3GUq
CV1jLeMu/mqkkIAFeDK8rDUkbDqyRGXROgYFa70mJ2ZCut1Gwm17b+M/UFB3H32W
jjl2E5NY6gbe9W6j902N7+XK6DqlM6MQnpWZMGBNpNKR1Ttxqpd+czyBDUvNzx5n
zzjf1Uf4QbDjF07j5M1u6HhCq36+1ikyOtgyREXODhjMhbaQ1U+uk22/wn8/z9+V
lpjQMKzWta3sEqf0O3+9+xvYTuZZHmMuDqrw7WKl8ZJyhgzROE8quF4GurKHCnbK
l/hArk6qqKfZ7hu6z6wi82hnfxvYlj9hzMPnRKShMLrBi0SlWRzqL/IBFYHS1u2u
BEo81QXGcYRFkX2muF3S3g+2tWvBKLRwarjXeicW1W2yvVm0y+DAby3oSexCCIan
3UUl9ZlnwZh7XKBZKkgSuCGNLXPnOC/dOXUCmLtVaA0wVDfrsgk5scqQ8VgleKvB
KCEAqjKjd5fYLuNKFATsUomeEphhwFflah1LIsrFTSk/chvipXNJVpzUirgQqZ54
stg5fAedJzEBzODVadHIh5M2tzX7KRgAfQiYUeWypKnf+pQ5wRyABdxNNkV+gDCD
PHVBaLQCH+aifjCR5rnLeSBdON9q14FmSQ3H/FRrQUcKbYWqcwspZQg22Zujz7kb
nSQYWk32QHyLPT+/a46FeVPvx0rW1/I3ryioIuxOr+DVieExlFDVOyi53Xdes90A
sSBg3uaV/0IYrxWYL3iGSujTOwc8pptgshSchTR8TR+I7MtX/pIy6zbcqMvn3yCb
4uRvbZdg+qnYCpc0dv3VQtTXLE+zZeYnHx5PItsowhqw6bz28HMjuQul3aCCqYKx
1mXMV0oHO9IeOmrcM8vdWy8MHsQjX9YJF17HTVngZRNlpKsVyA8ZTr/roMjVaAIG
YF8pwMxBS7yoNZ4DtASgsmjsDTjYyrvzKBXYgn67b0206fPy/dmEqGQZlAejluG0
xrmMqDQE6exffj09ZFHzHFkF7JLkePk8BlmQso5yjR7T2AkzPyimr3QNsDwd068H
ViYNAtg4xR0pHcRchHy6L8gQutk0DqfLWYBgWBEmhbntgpcVDpeHcBVe4Q6NSA7B
JgTtKFtmpDMP+qtN5tziErMrPdTF5TApmEHBo34QwNuDZkbfQVg8/C8y96JmaJuZ
1W9oyVIDiyDFTPos1Vxy8I4TRdXWCi7ZxgFCf6oOw+aMZ1ZoV43BzoIsIm/clS5K
IoGmI5elST49h9Wi4SHvj14rvkzxu5wZa09hNhxBUFORN99F9DWnLlGR1bSrdmUX
UG69l+hTgUJp0BeWCP0XjAFA2Y3nKzkZYU5swa7E3SVAf7FTPuDYJ6qnYdPbCx+g
IAAyCcLFvPBP2/zNq6qxvgGsIpghBnf0MmB9kvCNMkBy8f8bni0xoujZEbakdNOe
xAzjxB82YvOzDIEsxisE98+nz7dHS1s6OVsQIypXZeD1fF+RtAgAk1rAh9pqDhmB
FvbjNLIOf7dx6X6R7oR9BbTxsNPpiOpnSqIo2JtLgqFeLjms+1t2LV4MsoUxpOcC
Si21wbrdi7MwiDUVqVPhTDK6yCYnLNZ7NrYn8xVXB28ZMT9/Gy6U1RW1GsOcf+bV
BLHAPLFJyjWG/ps7wFLzBa9aBz+XhtzOZR12ZPSOxXnmu2qkA+mOuWL0r/HE3w2s
pLdHjl/2NzYq8vAPRjDlnzEQK1sMBKVIFTYFdswKNLV7WPj9DXmULSotFdBZq8Og
AxXnLcwpo8opZSVrdVs2ncfSr51LlM472R5RY1Q5ve9gKUMpgunDxaZZD33A8F7o
58RCxBynSvgmXZiTjAHqqgDrTfyM/S9vWdLt+5cI35oWHNbSGJ/0urKkusIbzDQq
Bel5dc5H5++rsv+Vi8UgzBvli50j/eGbZsA9vVz3segDVRIC+JUipKsagm4ApahQ
btF+OI4Q+zfA9NYkc9PNSe/hIckY6uUojuhIytOeWcoqTZgyQ8LyQTOi/7N6xO/6
6M8+37uRconSB5PdrxFbHu67zajZ24NpEqHQAM6K16p/1xekdNzmtTucvnZEUCcf
Yau4tPEVTciiaN4XaXWfhbA+Ug6xyjLAFG9ib0IqLkNPhJOQc4vy1BOsu38NLiU4
uk4FiD9+vgvmaU6X4gE/k1ezb01grNWYONeGEXbzM+kVpJrlBgDaE+nnHRarlzyi
Cf7TqnKoh3HK7fuH4kc+mr8wTU0RPrEWYyLhD9qFejVMW5G5aZN4S/+vvNQWpEWY
CBN9wvsHpaNj7Dk6EkNVH9PPBKN249XSEVeT9+gM1RhbFtjUmledWnGJZJqx7oaM
WsQv80NlApZuwVoOXaTADiwU/GoC3uNSDBbpLJih4qbTG2Np+FoWBgloGcRoW6US
Qp7cFvmpDKwdWE1FjXX1sIar0HMHU6FRnmv4p+ugSO84gsprmpyL0yYP1flxw1Rb
tQjEtisMxCZH7k46WojtlpBiE7Y28HGbnlx+gQuMZfRH67yvpzJlEs3HX9LH4B0K
tH94FtxKa95EaJFDg665Pjb20QZjOYEpd9KbHs7davcFHiMdsHolin7sNnEuSN03
u5lIthi0s6aZ3ZjEojJI+kOsoW8khqDen/izdsIpn6Vx2a62mo6wxlAHcY/Ku+pq
379TZMJEESbo4ZSbkLvvk8+ANSAxaA4COtfqYqTPp8sKnkXSqvpX7Kjcbj7bbF88
FCv9I9LQYLc75N9a7QJisYKa6y1fYopd3yvLVZy3reMaizktp6dJSzBPf0akROpB
LatLyUM1TUi92V/1ytB/Fjtu8LIsZIkWOVeyCY1CgxI5iuEjJlDW3PgWrKW4cKFh
btBG+ArP502wPic0A9bZzVmtedI8X31HjXC1NJvmHYpNDo/UAwIDfjTTN5I/krzQ
RjipkNwLRWj7NTtwQkRDBRzXmL9uhVbMKk+csIyC38q7451et6C4qnksEF6eqKMn
3q1grfJ/COnQZq7kPskSroblLcc2fS704AavYZRef+7iEApVz9El/41yYIeOtW4h
i99aK6KT1u9MsJYR/va4xfFCNXPrN6XWEvQtsrKF0Y0kVYWNhMcemkNtpO1FYIlT
utUR8v6/rq/9CTCu5QU3z00s3BJSP28wlty+cXeulyKOn6Dhdx5+EbNI+5Xpiv/J
OUJd4Bq4ZruETzLcCvz9l6tHZkhHmQwDNeG/iXW7qQULLpXzIbji+281L28hZTEt
ua+BfkxXFb/Neo9zUJ5B142Aab+a+GMsdfD5HPMFSPYxUe/S6FonXZGwAX/2rkwm
acphRZvTCeHPc0M9Xv+4xy9cC3zlF3/hZ8139uKRXci4AKkh6ZWSyzP5/IJnp4vn
iDoxCDuXBZKhomyep3vqkXYD6smqPm+f+fMpqIesmbf189mLlC4Hfyouqtq5JFrq
2KvbX0GSfS4L1QKC1N3dX3dAhwUGFAi9kZwiPpq0d4+xhnqf9uf/wz9vD20zxkdH
IwRvOvn2AooyokaZhvxZJl+nSJ4fUwIfc92X+YhccGym9qunp9oW2SCNjOGzHOwc
0ozWwQFMcHJwaWp40+baA9wuuHwJyqtCbhOykJdlkQG43mo+8wxmso4XCz7Wfk/K
Ik/LaNeJkShE16NIiqPYPHN4hg0vWuWbgMocB7f5+it9ix/qDRExjgRTbpiJKS9w
+DJx+OotIInKM9TtDxRBhXnX4K9zoCWI/oE4HB76FC7q7q9X+Yn+Of5Lpq+0rrJp
+ZB+Hq0p6UUPBSPX6323njnIb5BpKgzIl9yj2Hl2i5Qp4+YJiVu6lOMsTnFzzu43
YP2H+7HtANCodkcy9o/fwYysK9lNhFJzxBHsheo9oCZcQM7PxtgiS4c5vpN7vXx3
oOGf6yNCXHd1wsAulbc9ZbGvaTon62gV5fODLAlnALLF/Mse9wE0L6vvqEkV0Ey4
72prLCnf7Hp/00Jm+a5Ija7um+hLS9vXNLDBp6llP36tb06LEOy+KUugp/72HUoV
c7dLOZo9sHKVS4fweUzvvIiV1VgVXRNhjun1zAC/yg+N1SErO+7aPBdjb1ayXWx+
tPsqLwVHSGxRW+ou1yLDxQ7I/cnT7GpvWXPcqPRccYqmLlkwb6u+a9idLemhPZcu
aA8DHgJ65fgyz/h5MCzLoA7f3sADS3/kcQarrE8sVpOci5LM4bZ4i4DDpwLcWwAk
JnIS58VFuP0EryyXw1KaqrJ4D/HEcacZWaBW15oJeeRY8C4sIIFhFVxS+TLs+SSl
LTqLJNmKwpHF/6Nayx2kkZqCgcgUvPx1pRwE/lVnBLk6LtJFACEI57qVOUz2zTwC
SNrMIXHeepR1Y7NjpUuD7tMEIgTfUvbfj4Bjyc4HWttglCzIAkh/FlZfAh0Fd6Z0
Bx8R1sQOipkw1ZmvS97LPWA+KS0EnXxOSIgNDp1ZwWlvHY0dAbw2AxZ7hNkhSRt5
5+fX0lIGYNs8r5H4U7XqqeKFoN98jYEAgy2yWbbU+18cS06INjNDIyFXPRE9JKel
6soo/+pOnkb5bR2ZCL+NGsyIhEMlornyXIbXBA2NStlnOy9pfDbGFqVDk/LvCGq+
SlB/PMC2PwHpUFUQT6EKz41HrWbUwEAtKLHE57V/ZDwLvzomOv0xDEOXTPJtyXQq
/HCo/6lhBcf5cCXhZTaDJqSIi5l4Zg2IhkfpfbOpsQNpMNshRjFIUz7DchCbubuk
AzyaqRNxmm0wR5dytYxXi7aqOQ5EIzlu0nWmmFQh6jcLmvtHceR/qO1Q3eRlFWCa
mDE0XXzzkdg8FwnjLMfkAGhpR4okUZGUxcVd4rJwr+vKIr/m6PRrydNXyJaXzrsh
uHlA37EdlywFmXOxUQFhO8hSmKQmKRBEQYpynEqTlSc5VUWDzrR6rSCfwSn8206E
g1iGdJ+a4tT5xgZG/CDntGMk9DS/RE5OJBSfDnw9/yEWXXwRcVPrQDJJgUCl6okZ
Xtl1vfv9xkxA14EG3di7WU3QUmh+gZODDHVyRVjSikBXokWaPzdp06HDNT1bES/q
WOSa0G5akejqMwVs8yVxEsYE4ED7/3BrRzieW1gGG3OV2te/pTKhyD3FfPzXMhJT
QRRa6GmCCYoRmu9v8/1nOdRQ511rX6vdnUkg+b/h5OvSf6heaAdmkkwiczfFbFfG
+hAGAmj31ewKO4egZpaEFDlIi7CnlLskc/iI8puRl1NGBR9GxhATvjwfuJhbh0kN
KktOrDuxoLw2RM7nR5oHliN0OMeX00079mfhUcOXlJc8EaclxOj3FrmgMA4NDtTp
D2j7Ziw3yYhrcbPVtb9mNaGPmskMjfFpVggKh9JixsvbuES8B+ep5CtzVBFfY/i1
fj9piimqq3k2OouhGaYtEaLeGL6pMMQYYRZAzi1CNYuzzdo0OY8EWeGCWPzMR4a4
+mKknR/2T88seMxrQZgAKrbs6S/3w+4PsHjqRj8Iwuwejb4D6xQJVCUr+aQrPvds
lDriFrvLGGyXxI92BvbGC0iALlISXVCdTYIxc9LogJre8655rQU5wvSm3lcgMFEF
z71/La0edoeWZLDJmR2+Kdqs5vTWytQux1QNB3x68CXMgxfSOsyeFQZ9CbwFuyfQ
0D2hDUe57qz9qDEPzK5ivu1JbVIJkuvbS4OGxwhJc64Li80kDW3K3Zr646j8SPEf
Fnd23mBcbxcKV2GqEaIeFpKzXLEdWF6/8tIFzhYdZ8KYMBXNcGLexkd2PmaLqg3A
qsTiXuwhf7cGmqlOwsGn2IX/ni1f+maplGYayytxoEKIhH/+PPuFVWvEJovMB+S+
Zet1ecvI9Bj7oF4I6UtVgl8NZzj1iQmZvH4eCcGltXNiOJuVIn7n2fQc/KWXds19
n1XJtDyTbbOxmFh9D1TGjKvfSbKOjatb/fnXf6tVDx/42HKfqF2tGjuaghB4dyEn
Yi/ipP/PHicUry6+tGoj7zPBfJ3pWXmHwyfM6tn5VF4IEXSeMDoHLQe8aBMFZPbw
ZXh+GNLhEdtthBRDHDNb0URrdD/AbCyPC+3It7Wk1CWnirD6eFEHcJe0nJyxMi+H
KadO03CvnCUP2FrCL9sFt74OZO3nSX4nzZauLt4SXYYHLeLjraJ0Q0NiZ5wsGHdJ
DRrbD9sWy1FDL8GKvl7n/XhUanXij0nFwgSB8FuD52j4loFxNfRlKxZOqN5ek03r
umVyGp+6MutmlQXgWUh6PFD+eu//kvtoRY0AoKMY8yEC3YBACNSKmRQ5PpaO2W3v
kzWhRi+40XHFUmZHfDVOfREXuxBlOz0L6iIo5zP/0ebQx7HSscSRXV1Mbwu2rS7h
8O1I+7xvLBAIIemrUhcj98leEV/9B+20wro5Pkk81Dn3qi4zwZgMLnq6Zu0FbnIi
blQwHtlNEZA+anPEULg84DYRWq+3nso3a8PVkmznb1oLw08jRNvABka/ISzFcByt
95jsAUvvVQIqB5HbnDDZMnTxrRePYHvm9XpE72KH+bvrS7skecFuidI9R1DD62zc
8mFL9eiUSLnyZaHGWMRjLe5JvNqWh3qe1dpBkmhglj77MjQP51Mrkx2opJmfDVhe
J4PrgvMkvDyuI3X/iou4RhyyTCdvzYRnFCQHwgUQGCJljsGzX+IQ9/+70ZDpM9WG
YmTpyzeBGo8iuKW2K9T6SvmsGiZbk5ZgGiD8jOeWp6ia/DKeUSPwT2huLivkfyq3
NcRGDPkqW4fI2ZKCJuF6z2EnX61hVMIJk1v6T/hC162qq8jsZ7M2yiFNri7o9SkL
53GYNd14lf9M67qVOaJPyxU9i6pn324rE91+46Yl4s7b1L7MScatwQuwWV6qThAm
xG6tlSsNAm7anfvcfU77+h8U9VY3SbaoI+LqGPkbV2RVjHs4jXnbR3Si6vZ7YBgf
ugzxhN85uA9lO0TF1J9uiccljITIHQt6fn+rKQ1zzrCYgwf4r1KYwIXaM4RvzVSP
GgrrRuUB0RVjRynS7M2S79I92bKZ72r0WSxGS958OTtPw61BfbN4cd3mdqIGWdoa
E6jJHygIgGTiLGoYrAp/4Mj5B8FwUqreAxKLu5wicTzVJnKsgLjIhrKJDng8OJvl
78eKZVOnDYMxZzhmwtDJmRmruVeJwcJkRU7TPheq1dWBydAAlzq7cmzQmo/Ht3g5
GMGQ2op1SqLHhpSnY42WB/lDMPf7919OJHXosFf+oq/jWk7XpR2/b3J19C4ENZAl
9fvGTvo2n3qjc1QjfDAysy4q6vju/n1hhZnaOvezXfQ2eqyN+f5YBx+iPkalonVM
E9CBnG5mfuAFF4BfNJ4FJnV0CyNv1JThx2ef3jumPX15PFZcqY/G+aSi7GWDGl92
XcPdRqPbPWSYxkPt+js0goiSSXkmRv+Rgf5nX6n4nljjggXdzKlWVSGVXG5rHqTG
72pyz7aPL6pbYYYSAw9EnArs0Bu23xDkcHuPEutFGiNxZ7qcU2ZFF8kWMf1JYv+L
DKaTpSyGAFo2wmiRcZlKhItiUedAaNEkjvMTK0UEWKLBR1Ul1zh8OvJ5fECuH697
0Cpbwx9MJdpirZX8bhcpUb1YyWSMf5JOGFrmCOY1ZTC37kNXXgtmQeGs4z61AdWe
QVP/4quB/IrQIUwvLQeF5uRGxW2lmzgvdVUuUyFESxaCrI+io1CArHvw8VLxjf8y
8FnRzX6BccbEzQ/nAFIBN+GghpNkB4fv19NiWV7qFheMpHtz899e18zz8suMVZzm
IphoU07GNW48wFo3XfV1ckWfmt70hRhffYMRXm6qhyLjCnFZ4UB/IfuEIiPhK4O7
Nvhjul0o5I/IMG23uC1JBWlCxwckKh2cwZdnYFlTXiqTC5fFVjUavUpqy+MCgoZa
YdkHxmt4n/chGTkoAiX3gNugB2+cquUUYBboBsuK689nvBQgyVX1AFDlOLx6kcz4
GNjf9FGOqhablsYETo1FFigcy304Hh1c+derKqElBY9CbJpCl1T3OqNw1zBo9Q0h
UCSf8GC8yzB2Bb5xCbzAzAg6wbwNSLRvvtPlwZs6UwFiG3yTKyQ7ou83oPjn4o3Q
a0EkipBAFcEPqXVOeszNc2ss9C80d7FuHsJt8mkq7K/MocGSbDvdMVy57yf9c99A
+3oKfvsMvgckA6m48OhMDrXUKOLU9QcA/KjsEdEt8hsdjOuemTIHh+Xh4vCeSuh+
Eq1VCNr49dxmQFcTC1r5ghRMH0c2lc+BeIJK8pAZwRykazmx5iz/DjDXuCiCPlZA
jtMHO5g883ab1dqQ9GqyXiYZe3I/SIeB5Ep8CvXdPN/uHWk03/HgVn36+YewcvAl
5irPRGQwCQk0347RdhQUyoyLMikVj6Z6WQOtCH3bzvN4/8jh/519l+/6KcIHDUUp
IlGkXUEzv0S5MhyDLwDO7F5uGD30R06IvFveAJrkfwJ1qadbPZNIutHoEf0yIVz+
coMyLvp+EAA9RLnmai0sRtepgtV+rRO527EfmxTlHhCW4g5t5y8tt1bVYpaylnA4
2UEcCgsCOVtrKcW/FF2BkWjw/t/HwN2OLesVB+Ivk89YUyrXtJ5IARYWrBg8wMHe
yzZ1oqO0c6LNyWXEueqGUd8Mb2wFiomGQ/iC65nH7dTdr0t18+DygHmlA1ULV3Rp
Noq99FxQRXSiw/nAFJJQm0vQdg2dYol+INaIhdYicGF4qRYBmU224oPQSowXNVoF
EclDqoqibqgyyeBlVolmFJm/MOkPt622gxb87phjyvT/P9HtCFf4h6d5fgtJsrhM
ROTEFTWdA/9oeMJwPV17fmau+aevhNCyBy1pieusXANMh8fdxHu6kU/WRxZHT5xl
bOzSGPL6os8VJ/eiLstNSaaoDlof10ruP5bCI65ZWk2I6FJMNkIE6MtWEaS+7EF/
YtPi+0wMcqf4WsvLGuID9q2YLztwXbVC2UAiE0MGADLowz2at7w2KzhfXDQP+oJf
1HmCKXex5qb2W1QYhkXLbisSPmdPXOe3Z1g0W2sWqyT03RGbm3sM3tuQH5uzGh8X
KIdcFdq1X8d2iuTaMayBrjFJ+3+KEZUAfsMTywFpIuBGpuRqX5a66nqu9nOeWvN/
NNXjuiZY9k9RrIS3cKw1UDKSxYR1cCdCJH+qI3IIYJm9jYt9u5CM6QXBTH0Xw21L
14ccjFGNcS1UIjr2R7mbu8HqfZ8wtfwew4r4mYT+FYiDrsKiJnMvejbEbJB8j8rD
QzWkp47octZgsCgj75LUmxCO2MB8TUKsMZB6Z7Id4tWEgKk1pVaHlmAXj1m+f2sT
5/49EKjZDNYAHSVWVN3vptWe0V37v0NSaswGFq6eeQFA50x/yyNeZbtu1da5fEF8
FvPAgnN3AE7VTpdVjFyuqgZBX+XoIE84Q+O1LXAlKO0DAerMWOcSIEXDIwcL1JyM
Z69F0pgG0kdyRdbLqN48VlYMATAOUSgHKIJV0ff2gx4Z8IvNda+P7y80xQM3kr03
MXF4u5EIknJqrw1EwLkz/6SPF9udLLfeKdDuLfFSHaJ3IcpRB7O6bB/GnRxl+kTA
SYjN2LHy1hw7k17AjZ05QVosdAveD5ggoju9t/g2r/5TvfACb/XR4Da0ig0cRZQ5
WcPrbi7gnJEAYS94Kw6E1XEgahCbOt358qRCr0CQvD0/CuRfTL7o0WU8vqst+w5f
pX2xKQ0z86CrVEX4ACntok8FWvfZmNMaPklxRxA5jICgX7hNtUUJcyWnwo4WQCCd
y3mBLBVqPJuyg3jlKuj+OkLyZ0IZNnFTXUWn/qT8mD8g9ZrW9ukh9Dp970CgQya0
gfORiR+jrdDaPeXgQBMByypZgcuTxH2up50Rvhw7tHw90tPcllIagvg24xTdEXeS
dq1J6QETQhEKA5m/jk7l57DOa71m4zmRq+YUzU7T1rLQMf7fKzxysogFEp7GFUiQ
vKrvu3x17/YZW1YRY2qAdaj+xDLF25ZaW9W4h4smJSlHVGIZ8k+kK1dBhqgO1FlK
mRdLmz0zgmCdmgTK9ZHTb6qXL2V+ZT5Uz1RxludR/JqamveD44ndAKvN4qywKDwl
zmNV/Esbr90aNieb26U9oxRlEk/yBnbhIXDncFZEVjJsbqg69WNelmO+fi0uE7oY
8n6xUnnoykPJkAP5afdm89Hn9WtUJFSDAh6rRjG8+xEloiSWLRr+TQXF89gLO9pZ
c0N+u2xlcKZDkj66H/fSNByL08UHUkc69vqAm5QP7FrYVhG0HnW4gjehgKvL8Kx/
M21fpzhsHZ48ok4xdSJbjvCV9LbddhdtSL45Bl0m1LKVZCysd9fOQOtLADGYyqvv
sDRITdzFwQ3WFzq1xL+Oo8TVII0Sd4s0BX1dN0MsQYyLDiaHNqCrGUoXdB9/pGv5
3sjnT+xVtFl5j6LwoIszPAAs4nIv0An9keVHbThbmX/77SIyMhXQnPZzHGhX+noN
LYDAqAcFQHua7bPd1/F7T5CVfIn2m0bFHvPrvs6jSkW2SFuHfZ0lbodURrx7qvzp
JUGLvdrGtXXP0E/du/mJGG++WQWnueLUHzcgXvhNGxcg6SLNVwZlVgX4yNjQuX+D
T3r1EadN5aWq0xVOA1q9a29IbHpOl7zq8ZvxBktQNKW9jV3jo/rTzyIXQ8cD/7JA
YKUsyUEn+bJEUmLl6AqHPrd7YHpXrCnLwsygdyCxPDRXHwp9VRX3LERivFIKpO9v
sV9NMVFJpkijx0oXFxQUfA6eluKS52avfj8xbBGT6Mc6k+vbAgcN8Euu2Ur1vT5B
jHQ9kiLztcgDzk/77Hm1EHTHaX1Z6oVao+T+9zg/yz61rab3J+7C6xRNt1PvVntl
tuYer9MNLy65EGr102XuJWs/9vYclmiCgEp7zPdZUO3XblAYOdKPKB1pX8jW8ICT
oFf7ydy4q9lhuzGRfk18iulWT1s5cJy93QpvcMPjbUoEtEKmSTOkLFNwd4DAGa3d
/Uhg1W5GrUiuFdz1o5DB8OO0dyOOmVe2Eyp71zLtSukXruYXzUYgpXeQVetj07EE
doaRfh+Qml3eijLQzGsNAA1JC9+8i/WuqeMUjCh8X5ZHBNzXXkA/DC0GxbI2J+UN
IMtLYjsfThxj4kRt7kW7a5K+Gmn3YSnQ3zfdRSRKqQYAoKokPsVmTLLc5Kg/QBuQ
D89uFDwAcShXS6Ko3nscj9uxa0yKfRaaqRSr4CXAbGqjKcy0Nt1zpC5Uu2F9J3hO
KgcazJbD/pVQ9imsK8B8Z61JMQPP6LrQ+hSRl1UdXABTB2Z5nTwDQW0qWq25JMTd
VsnhIDGWeigu0aDu8QAiNuAmyyF4u/6OoWrMvmZFnPHccFG14Fy2AKQZ5GwU0Gw9
FlGB0e7Jgs4LajViRCahrF0cFNOe+KPOyOmsZFucocfHKWjCO2e+UzN+b5qf/SVj
pzjMWQaEXke1+1H71QvUsfvOzP3SHjOJXZvfXXbV25dirALNljKt/4UzylFfcgwY
p+07s0rQ0E/SQGUH5r0uKylA7kNRRtRFr6EBIONiHhRW6RQdffLETSUUcUUbk6kH
25mOyRd6DGFR9Z2ai55jnG72CTVUKinml4t0VywfYmWLxvf85hWzibKY1PyDiDaT
WMaOHHbsI35ylfWgoeRAR5gCOXqpoEe4jnYFn9A/6jNSXpXUHAVuFiuwywiue/zB
9bt4jFSNLGS9u/OC5li9a1OFSxjUzPnqzfw32eNhohu634UUlMAsJhzZ8ERTz6rh
mMJdHFgqD72yADBY0+7PuJjK/3rEQPWBTcQuz6ohXrntoZ+/RgrKPBGxQ2sMbXOq
eeNX0uyn1eZfE2muGbBXYYHNOjEVmKo0hY3kHHaE2ptf+yZQxAEHGzOZ1gapzFuw
frGKe/84IVkxkcq8sElMGAkBwQChpj4pd0ok3OLL1OaAw8YvktIU89/4RsbBoJCM
pNERrT8Bpu1ica2FiWFCyIgLuqLCB+mAqemEIJl4syyIW/46TsO4syrzj1VsLVIp
bfPDaKlbdlsbL3XgNnmZcmpATPBGl669fyjkuWArWtSHgUyvVmyiaDGbIK66IzD4
t5aP52n2X5vT0EsWwlijnkZR43A5hmQboJINlNtaAPrD+0hYsUmxmUc0tF6T4pRl
HoytjdPLU4FVU87KdyrJMGgqj+lqBS5gfuL6ChasKvzOtr6t3okAi/fPV272EjLy
tM6m/qSUtuuNiNeCwo68dPjtzMYamhcGQy+bcDI4ObJlpqdnKaqC4RLhwCG71y5Y
fgktyU4ddJzWXC9h91zZ/bmKFsrwzhSk76K4QMfjle+MSaVj6jczM1PaKwGFOPzW
pCCnq0d3fzLceeotxR1sIeJCimZqi6mcvKjz04/vLPgEY6Ij1f3UaS2A1OxMHMzz
ttLDVFbQ2dAPWiu6im56tYWzhmoO5IErJ6XLGIhOBPEsQvOI5bJ9YbD0nxxsMKh6
cfKrv+skOv+O4644fYEWTMf/RAwT57ZC2aygHDbr7ekvRTCTjEmSH5ZvkJstlEU7
GAkpsj2UElp/Gst2beczqhVYWotfr9/FGDxZ55Gz/8lo7Vb7kEZtF8+/nOorGISK
mVMkcAN090kW4nc3s2m9zekTb6kX8hP4zSSeOF6GCe6d7js6OgAg0osih/Oysb6o
+6zyFuoG3Y6+CBxHolvD0Oaf7ESjrNA3K3wi+0mCDG08EyxW9/eL56bhHM+PXplJ
9Y4ZEnTN94VyMNnq9OIwssP/eqC+MGZPMv/zxGBEgAk4R4scQIs00acw61Y7cPAE
+y/iGFEa86zTqadx6hoUJEy9fI6cP0Dsv6QtUblO++ia4tOrYVjhR4OFapDd5lAr
kBqzXpy5THLLJsNicG72So2lLjB5jUuU9VSXkJo6bOe5djJNQoq3KGpNAFRz1O01
tYcKl6/6fbwduS+gNNw8MXBPT3s3OadZpr1cGciA6R1svFP5u+BNqxaxvN4zut6U
GWafaRV04rK86JKBy4yuKOsSBS3kKi+80AxM0h9bo7DLyNBTbeXCiAh/vGmEb5ha
lbdqajbgAChcIeAYvGK+Y8WkHDawXp90ZFowSD4ck46mACYGgp1+tvbWhin5MEog
2r/MaIUtV5wDZ0UCDlKpMsg4O9qtf5ZkIDIu8GgH1GIc6au4AvxfrjsVvhJziiIN
/5FbeZ45c0lBZuSgZ9ltbf1PNWoMnwPdBc8qWdjq6HuHE3Jss1VkxU///5fs+lq9
tGInVGPCLeHpvzRIHHhQtKu+t2lM/hRAKtGml+Tep/ktBfQZuv7ur3zfWnXaaZh2
WsJhcrCcCquDinPbAclTFKCUte2Dk0ipiPZ8Z0XR26wz1hUJ2OEtIaCAR+F4VzJz
cyiIeUt/MugA76grQdPD2RpWxz8kRh0n8OCf1qllsWCyrUyTw65wzU0bXG2fHLd9
vDzdOOJMbjz51CiWotqn7goHhgSopYIA7k7fFxgfvtnK7Mdb5IIhOUp+58QttYAF
S7AyhFW2ghxhjo4F9/tZCtLYyup0+oq1Ln6FyD20hGcPm4ziIzT3aOSVmx4Aj1p0
ziAhGYIGrZYUfDLVIe50vhW5+Ow75X2mgzlciLod1Lm+Q+V9PKuT48QEpX+wegsx
x/ZAeSvvzVW2fCMWYAE59dJmOkFCOs02QRqQ/TheXe6rpYRCalMsGpL3n0ab9iw4
y6iept5L7Z8Vys7VmwQU4X1079n45yOlnpVeOP3PsebGtYlnOKsMkudGgv6m5Hr9
M4Gep6HUZUHr5mZ7/9I89/oibdfRoYJswwtoa7Khph8N/d+9iadNapLeKbzSSQ29
JP3Nhzkgp5BQsu12/t8gk22u+1rHA3lXkL3b2TlZY6hgZei6djaEYxVpWynlZRPT
7y3f+UbjAL+WLhKVQi2EUhiAGHeSVbsypirxf4lHyyuO43H+BMauBLv6YJOYjWmt
Z8eg1VaONBJ6XL6Ua3FGbcw3pK9mc6cZmeJXkicoZm4tQavRArNk02iZHWQFg3PY
+KwakK6Umr/BhbSMkV1JGDIB/aRF3mk3BtKLdyV3ulICqdQBQ3AgBqkrzVShi9s2
x1c2iEF9GTvxUFazMGTGF9WPd6QjZLhSCp2P8VVlXaeMDxCorXUClXM3+zMiIV+Y
GLFz7QSyD4KplRL500he5EjbqwezQsgCAWeVk28joolknBm3gyGq8YGL5WNk9gZO
0fkorbWmSqkexRLR4EQvBMj6ETT8rMJDEv9hzboOodTDT4U20RIdBHl6Xvj5tlkH
cjMhtg9DMq8b32wIZ5iqpWnVxd9kuNoS2mxEHfrZZL7olf3TNevNIzYjK3uotDPe
1jaPVMfbtJHrG4NA+cBJ1X29j7DUGp40dDRk9e6MERIT70GclFDRT5xCK/Df5vM7
o6br66tbLUXn5KSklFLiZ34q+DuG48G8+FdgqFJXBTdf9UeD+WxMEM35G7p/H+AM
nSWqyeDBG3MVnoPmqXke0AHKil019UKCmjmF8NtUGGbgWYarGSXW1trCecuQqI8J
EpZk7DUCnfuJG10yz3Y80uB5ZXt4f2hljItC7mNfCbKYVA49WUGPD3c5HfZ6USRI
FD49A8kbkW43L1/lTThvbx06MUPYRT4jDG+NZpaeNCL7vQq6gDl/y5+6xFOJDymP
cDlWt4Pt4G9PuTu8grP3GwkavLrKgG8dfp0+HnP5YLJmp4RdgZrqsu9/RXvIyGPi
K8/3YqcIR4AXNes8qmM68tjaVg3aMxCICnIWrNT07bhoeAATRJuGce3lnhCUyzvV
lTClwTmI816g0OLx3SLqdcsx+JVUGxtUz7Rw7mZuxjLS5YAHm/E4hzdzI0XTofT7
G5gADsbNUz9HV6uq0lWJ/K0LaL6+Wvvh0bZwfR54dmZ+1sXRU2GuEM15GL7XLF6B
T/AAXbJvE0pxjg5mJupS/FHSZm0XddqejA2i08Doh0Pa/9Kceg9gwjssxjEQ6/0y
UiOsvxdEeA77EUXtafzpUX+PSt1gWCVVDCwrZYQ7UmDQizaJw7abJFvLyTsFbAGM
Y+gkWz/C7O61wgZYfQtTJE1Zglgzxvxy2C4amnU2CW0NVav3WYzElb14TcalFZ+5
IRlRxR3T3eRJXaBnVGjx9xL+RkdiHQ3M4oTugGggH/1NT/5r7vhD8OiMcPKE0Uje
K1BZwR4ozm2Vr/CqKv1OKUkvUuT94spwoiEJjpEwNaTXvlc14lICs+5yPCLz4FHf
mXj0SdsUA+A19P3yEDF/WJdeOApLl0PSGxDN/brD1h4Dkn97EvL3Sh9GaI+lrIcP
FnvHN2RQtfizMoGg6jHTzEoG0rTTKcEHxZ1OaoVffZyS9F2TrPIHPXw7w3poTO9I
jpbPgkIVx4zVy7abZONfBsWfr/d7Fvg85Cf7LCgiN3x3BPOJblS+HEZFsqL0pTmU
Puu5IV2ZI5oWNQWP892S441XwBqPFQMn5ElepNpt+PcjXyZ2Fyf9T8dxPLHLDbNt
AQvbtycdZAlcUCDoIOpIgeUNU25RVsLlxbafd0b4HMIqUcPnIiZhIrEiGeMYB6Qj
6qwxR+s7hTVDjbVCKzdQF7wD27/t9Yw2zcprzoCqaSW7rYsWM8UFhCjasOL/asKH
540J4NEWXm/dvKCk1rcE78YaNU4hyBVX+SlcGcN79S9TOWHmpNRJRaSmkAek85Jj
ZZhJi8zjQsmTmNrrMobOvup+BE6cj1ac7unYgzlqBiOlmu8cP4zRut9GtK/QoHvS
erN4V+usG0c5Lcpm1sHLjdfw/lH6S4Kf+U+jGPeGkrdfS/BvE3qu6a9YlxhQ0xEk
MCdBon0/WbJyZ2zKrmMKjEKAwhWt7P9JmxX9d0NU4ATJBqlDiXbd6bLTLWW11/Zp
8NHl2HkMbM+sSuhpnyj1uz9emmO3H/2y6WHpsKBx7xf5k6Lwl4ZddpQj5mUq+I5q
VUtAMonsfp7IMpqHnSx9I23ZSZBpe2M9kmendgHxHxYnShVXfeWZbqikOVriA/IN
mAlPSzGrpZe6hjB2rEM7oAiKyhTI31akLn7lYtSNg1Ol0tp+pGplMbIdZ0ujDrv1
mtMWa0rfG/lo0HdLpb7/2xbtp4W93UGsKvZp1E8U3wXPsSuRQlwxOUuePZTg9Qwz
jvKhch7GsCfXfGm8Zyvy6Snpa/wyCE/XQg/nsuqjtdY/oFbiP73+mc/zllTQR7D8
EMwkiKRzk8pq7IlnBBu9gX1CP8MZwY2dBSj1TwdK0mMeiwrXJKgN3k3Z0Smnwjdf
kmJaxepI1WS5JeQ9Q++gPPXvAY5qAiyICKFL9Dyj5gCvUwf7Wa5duQAYqirwPlO4
oadrL1zVDbl0a3RgFDpvA/BuDuThJhZs5Sl0uw2AJi7f8wpZGK9IgIRoIbG39rx0
fVyPFIk/L/YGw5p+Vew1zIFCeiteXCAJdclF+tllkdm2u1Oq4X6nIyG7zeeC1ADA
6FkgCn6Y3ZIceW7pEpnt3iRcYJO4FdHJuzwFVwxxN46XPtM06N1N/f5FLmtFnkXq
KFdiBT2GnN1ckS/2uCTC5viOkk3or6CWC9QzL74RHbIkR6Jhqfy7NeT7h+/KL0Gs
QeSrIfrVkSTjZ9DH9CiCkqgiEJ6lLMNd7MQ7b7ZIOSFBgpiCyUErVb0YtxC8d5Rr
yqX5bVNqWmIpOKfCTaB+1+nwjKvT6SZvo9CjfTcUv6czLZlv6BZEaJqY8LIRqQX/
K4cpKfnGVKva/zGOAP3SJ2veM8Gmq5+tASIeUsv1lzvOnnhoj+3Vj8WrnAZSfh+l
S67AIxq2GMXOwCEC62Tu8riRLncriuE/kKj+CQt2OGAiaL4HO6E7GkvjToZnSi/c
CJirm1tjrkZLzPj1snycVdSWzlM0jkXnK3hp52Hj5WabR7jPfIvby5cigg3deWhW
+f81Zri5B0cSYnDTIBXXSuT9dX52YAIL0GhtPQezF4LkuyPx0P+sSXjrh+ZmgTOa
KAsJcoESxAd6nuEo5DHOz3JNtl0W6GUu6YLdjIb4tPJNvRo4z8I9t5PSfu5vNXuj
TPvPe7ARf6p2dTw6sN1pfzdAn6hOyXuAVhOOBIm4t0U3Ns+iGr6UQK7DS25tOlsW
lxpFWUb1J7YBn87q/Mk+YQEKA+8GIpiNZ1XkrbClkZUPp4ecm6LWj/QQJo7Kg41s
CiXacH1rqXp4vMnrsXssoZSR5pFtTxYmufqp/MOB43AZ6Czfy/h0189mMbKgnO48
EY1Z8z4BmbPKUzfCnPOgP0ktpFAuMGXqAFrjXAtDu75n3lylAA5g6tYXhXcclcD8
2TCmX9vJq4PJ4x+MpvwLXdvij5JIauzXUFvoxWmUp4VccsMI9un3HY4LD5ylNkkC
88y0b4K8ksni1IgjSNVPsxVuoGGhdmOjz09ub5d51BQ0GFTiwT2wVTEDCB34BVrb
z9FEWRo1M51BK9En1AryZP8osyhCWrFQS2BDWKTO+uy8KifNGOE9vtC6+/LVZ2IC
TJQR9J6GnYjD+Eqr9ZCJStPHlW3wHibKGhgRuxbJenCy8W90bLChUPelAuLGyCVB
cgkLaQACI4mzCrQxFS/p6guwYxymaaC5hvYuZ/TSke0VJ5d97a6v5cJTrzxksaTN
S0LN8hrdXxPrrcfebP1kN29wYKDjzt2pssG6LcvqMZzkXoj7cv63DsUl8+YwkuCD
+LvmID4H2VRHnZ7/yA97RqlcHTWvifxKwMgQB2OMvEIGdflhJlEVAINtBusgerBk
RbxapTIeJJKHjvclL57dUOeNp1itRaxdBxH2dhJ9e/rb5p2SBUc5fwJpQQOHTmGA
oiKFKxSJumdtvEVoM8OMyWzDNbmvEmgiimpKPdb9zJMg0rLJfAKVpSmFA38tEbIs
80URn22JxaR2jJM86hZ8Y2/1a/lk+WCgViZC1DQpbcWXHgdGf9y7NpizbHirD7vK
AaD5Jse05Xt7yqAuRIzauxD17R84pI2OVYV8PY/aauaj94QYW3LM5Oxo2zxltYQl
VYDY68ald0MO7uSDcU3heQPizhNz96/CMCgCGU/H6L5EqHbyR0juFJNAaEwHd2ac
//xIexCJPex/EMyjS8cKki4os+ndRYjNRpz/woYSj+9SIQ2sUlCSVjVpv2Ra+C26
DVCuho/vhaOJtG1auYCdSbnmyCZ/C3W0Gpw2ZlPmphWjTkrBa5V5yp9TG62G0WBC
/fnSKbgVGQg7gcGlbuggr4ge37Hih1zKTxo2lGvTAcNhdDoFS+mFzKVa+tYdUpbG
EO/NyH2Ku5ZveN3MUMe/8FsYFjtAA+LmooneIFz8d4YSR45T+AHRJ3N5loKf8Oka
z1rIgY+82TpV4A2GMddC1e05EbSUZsCyF/0BSIitkejnD1IhX4E1QFqm7I3GPXpL
jdMWZTB0nXGrLUuagkGvkwyUnBC8r1UDk0tOhEvTubNzvDzO19ZnfEuyeCHwDYXR
LYtyLWFdFD4VsCWhr0dV/2JF5PEf40o1clORl+MGXpVIgWihKly6ftDTcqW/ejxS
rzYOpkQrqJFbNibPY1YcTh12ds63SJ75g6z8OxfX4seFhW985UVuZPSSVp9P7KLh
Roq2L/ixE2S+y1hoFWPXTwMPLCcb+804JWHDU3O4+qIAj16xs5/zT/mZqOhd1OYb
5F28VbN2oVRIFCl76ZBFzKqx8RdW2OIbuL6c0EpL4mIMiJMlXbiGLVJGFSaqznCt
tidNaIjTFGhROwpPC81Q67eNpuu7zKtfN/pioSh4QHWnpO6BYww0w6vqGWQfjsPS
sVgDmn/p4ktsM7RXts1bKNI2wkxRGQ/Y8fPolEhO8xHaXoYj1Yw/hZ/sBwG4SkVO
bBS4LGOEmPdOufPpl0yLZf7tV76rphKEDbjx2VvA0o1LPwJKTjaztVkcZC34qJpw
+3rL2XJBemcLem0jbi5mtBn8XZHqompWIAA5WBi2sXEhlChOA8zZL6xxyh/rcGSW
xEDDZQXLDrJHYC0QQ8u4iwmZLRgjII9N1mMfM0AHRXQcW7pYcInbiugJ6XWeO5FW
/Ljr5aBbctPvLBroE0H9QRXrh6YeiSd+uBYcjwz/RAsqChFIqJza1I164TqNaqlY
T31g4hP8cFMvaUTJAiOSlUp74o5EUMtUqABSDPJsZ3fDYMI2Mem5pMGnOfE6OXhN
Tw9yhn45uwzg056acJBX2jui+lDU9iFxnAI2U5Zpmdyyi5tG7GnJh8lj9Jrjyj8U
5JpnuuKGZYQtgkseea7Kw6AO4binh+5pLRaiey2BGZhq8Ec/Zt/c95EUSXNkWOjZ
LUHRYfhxUQFWF+e3OCHdjFL+trBHL29BWvrDBf1POUxxKpYiLkK8ZCylLLOAkAYR
uZRMkRQbDpm5XnkMc9NqQ+CEAl1j5fB5tqmTvt/f2echIe0mdGKX0mS9+y1OuZ5x
ixMBMEMOgXfvqhf7pIuKcdDIPdeMzSisyuBixid6B4kw58zwMBscc3+iwGW66GOg
ZKv46naqODioeidBrpN0P4FFlzqoWlwkdzBN8/cXkF+mgkCUeNeii9cwKp3mtrEB
ahAaGS9Fvq39D1yk7h0czo0e/+gT0eUaalWgGiTrwFCgecyfkqtyLNR1KgBOlpcL
GJC6I1nyV7hud2dFZ0O51BJBFgl3W4mcnTd4C2MawVzT1Wp/fWP9dgbyo1EY2hD+
B+LIf6oZuvOGsNxwCTfzuEzBovO/E0Jn/pF7cbbDUJvb150cgCShy6F42eBk1/0D
CU9xOzOgpKdungMay5g123op+SwTDPB0Yuo/y6R9bXKgTS02QafTj0HYzQaJxHXC
SEuLzSPyHUBCkRdj1p4z2Mg4WicRzaKtS5N3T6kS95jPLeoA4J7ULDtmAPiybShF
88b1Hku/4Hbg6AjEUdyNqF17JxB0VO83M84t7KSrA4aoCyLPT0SqIxIbeRyUAhxM
3ly4H/QCbWykZuzfrdSaEPImtSXh84hZ0cbEZBQ1cQSabxG/v2SIxVAu6ncc5a5R
HIDc1zMp8Tm4Dl08ItUXl6xtBAWaRcpz2iFG0yKfX3D6mUxjH1Gr8NTsOgNKaA/Z
9XgfJpgJkzcwqHs+rvsBf5Ihu+NK3ISbM9HIjrR1DBsX3CAbb3Sm6u48df9w98a/
ZV2jyCiS3frs+qhPTIrg+RtT3r9wTdZsDiKp8uxJVzrCOIC+FRcEGYJud0XzHvTA
x/YIPHM8DWb8Jz49/TmY8cbHXN3qndMy2w2o4fd0iQTF185IMmmIflxSAXLVVC/A
1G6/bL9GCEXuQ0t6SP5rAiuZeCgy4PQA9iNlSfm6BFtbZ4aBf8ECTs151Nf5gi7L
GpTph/thf0erQcWQiBPVPLazHUF2j6BupTOB4u3P5cBJZiP8dZI3amH9m+LeczN+
vLLyyebz9R9YIBAkJA6Vd1/gmYEY2but0l6UZO7JH/FePxXVwdhAySBRwgfuN0pt
+Httd48X9g9K5EmI4LVI629ZE2kBqqoubgrMCv2V1646E/SghlTcADSc7HWRvcTZ
z2i5WM/Kuz9gGIpDQDoa98JtXrO0sH1fb4PQoPHcyu0SWP+MEsD2LX9s/1MXdQGr
f60cEWGI1d+QLJ2ur+SSPfgF5Iwm1Tz/WfQWRyaFMSlStkGdJLRC9NPPig2Y/6Or
vyMAZACwGXHfHyajj4rXox+6qjiWrXo1KK/fo2IM4BFpIv60le9Qva0Eo6IeQ70H
l6V5d+Bgy8Ql80xI+x94uHKpex0//RQZb2DiHZbwSMYiyBKeHDlWgmuLBNlrkBkX
6QUKeBNRi1BdRunFdXNlKxQCDS/b7e7miIS54FoNWuRM1mv4MDn7S7zUQZHXDeIQ
Ajy6KpBvJ5V5sNHnJX28ZgUOTkAazSZCkZqtp6DfnDXINEilj6yb3pY14iB0VA+N
Vyi0pP+vnxnEmDbqRa1nWqbiRJzJl5FSiEyCz9E3HOvGGaqL9B7zjJFqSaz8zaZB
+gCPSi88ExGhyhSLYEVnOiByB/YTay6j1nTynh/vlpKKSVjzEoI2dUXySZNR6lM4
GZ98kmv11mygvEGRdif2ECXqSapMhAjALUW6odfMTA7JHPSYIqUzT5YBVFwJNZur
JkxdbImde/gvZFrFEYrmF/NOBuds/CIWQAS2/TyAMDmWInD3h0hOtv3zYIlbbebJ
z2k8evlUmgogYtkDYxjKLF2H5vMF17PzXCdw0vBRGNXuR97q/82n+8ZtYMY2mvVm
ZGtD+ZCTS0fAABHbIMoIlC7EnAwrIZXe1Yrs57ZTZlE6E9ZygKVk7hTVOb/6EzYx
z6k9oEiZIhFlPKm/dxLQHl0vJYxz7LwIQzdmtTy3GhEgjc2Zrvai3lI4aSCvembu
gqjnhmRVONdStp/HnDRBU+ZQ7LKlQ6WH9LEdAukqXCaUOg+ovDR9X4gX4O9GuhJk
G0WyljDaY1KJZf+HNPEY2ZhNbF1l4trIonh1r0Zy8I00nbSbTfgnlttQ7R2Jz67A
hxrtdxONt7b28LmePhEkAEMcFpo0KIvrDKr8MNKckk/dhLrKD0ktxsGeljpSTBq6
m5aUEYfliK0PD2nIQ5FLy/Y7TnZ2I3b7PW0MsFMe47ewPAzJyskfcaRt0Crc/tvd
SLqJajlLEqUkUm+1SeXb0JwrsTB1o4DXEdxwgCZq/Tc6vUZtWIxGOMIFeJgnYfP6
8tpPszhjDauSpQKfOAtyHTAnqLdPwMa059bnhdLLT2KzxAnXrmUOye8RrPL8+Utu
DOLyAPfwNzAUg6q7+ZAqHS7y2aA/k174eOskEWOe6+4z/fiQtb3Py+yOPw7obrvY
WNxWnF3HJbnQYXKAfaj8Jsj34Q9LRnhK+H7Oi7HCMXyNSqzKaa7hSifOl+xdiDoQ
igYG1wzoSN63lsv43J3K32SgcPSJtBf6Z5/ziI0MEroyCEGKV0Yhuf9vH/yfw5T/
l3MeWzpAc6nmMbu+w83bvj2nnv4f7o8CFLerzYSDyO9cTv9m2/6RRt1jLmydGHZG
7XHUtMwtCu8QI02SEJNj9oaNXJTEr70Jso0xpsyqL9x8S2Hv8GWqDbJBtnnEnueA
gML50iyLjARngFH6u/QK2ZTy2yyPjTvJVXpq1ENVZE8VF/5W6mzGtSQZHaqomCza
D8H1dGyiRJrydO5cVYhD9D4vkOX94XAotkUFVauCpszQAwqS8WoX1CNMa1enQfFT
Vd17mcWebYoD7+Mx/vZf2FRraIeTSKcQDaEaDZdwZQnnUVO43pAzewsEYOdfm+wv
WIBZEHqKkJvs5gEbKEqz3MtXMMg/5QvoApBz4vTOGv/0HWWkRPDm8z6oNhqch2Oc
le3j+3euhz6tii/kri7FudahDNtqHRTBUSJr6fuxE1Ko9bsa4fL2f+fiIsSHLTrL
B2afXemDRjSTNrWULsNcVzvj8X/l4La+jYp7YO3jcOOK34rHIIBEPFLjL3nLVYS2
BhjBrRm5r6yyWtWj4BKbZ/79IGVZ02ByjnwnAbFPnGatnq0UPp7kCfqUA3qcagp3
L+ldPv1ytU3V1eHCdBjkseXd91r5qfSod1nzm8wEo5vjEzVECz6JfPrOP5O2HBn1
zzIfRJsGs5GwknwWtZdJLHnm7WhzTlNxrhLUWNRnR8tdGimwYzkQjLrOBI3Q9rCv
Vo3enyGWXMoH9ta4cp83W5HBCBMuQ72PMxFTkRpPetCIhUveiTXy3+Zsq8ANaUhC
pEYrAYkvWuozGdSSUeyzz6WQ6t3+m79dORyJ64MLepGuADCPor31yaPYvTl243JD
3/77iKQfl0KHDmladGWbFT6i+x2fKprz1LZyaUlDwFeMjDmXSimg2ZIX6HQSnv62
JlpmbxUjec1P1ZSDgSHgFO5gYhlLL48WzCp9nT4QxsZVYSOyuoAo8KU14tx447XE
TUvJfFU3jGEZGm1wo2uu1RZJdklNS18ueBM/7+4PfBoYBDurJPGFwGcR11VqV2N+
2h9hl0dHlj7CHgbaBoolOP+jejql4CaC0Y/uR/uXZkQzEKCry3wZ93vq+QcRJhQV
9FitbhZ3gT0gXZ25ygqplT6k2q12cTm1c9oS4OR4rEg1W6atx9ggnag0k1chU2hV
JARq05o0As2NKWNAu8O5QfTzr/pB0w5a+icjiAhV4Dx47GU6poXCpwyxYwOs9vIY
A+vBQ368Y7nOmdhuKKEHhVYmp83Rx879FlWNpAKQgJ+BLrroUzpqnaZwIrLUEMST
pbmIpSUMeAPdQG5NnLW++3xtw1wMJubYRsHcTYfzYZu0i/jaDyGXmio/q78xK06A
edFtws/bOpr7DY/G8LxE4FS22KAgtG8zxaszcKzm1bVEeZWs34q9q0G5txLy3QSi
iZ3hHBZgxO0OrUPmt/rArg9zMOYtximcD/fnfS88/FX5OTspzLk7QFroS8LT7Ic+
ArzaYuYQXO8jspUv+Bv36kI45SrT7Ra/O1sYd6TyIT8AWN9q+xW9e1MLdjlAImah
bIpkl9/XJNWShmM1hu2Gdyci6toMMT58Jusm2v2twupQn7IFTtp1SXWAShvPVPLk
Pxw/wuObeHiERXLpBuxy19g9ekFtplzaqdcQ1+EDd0dlsMNu49+j8pYAItltvFQ7
ySBjSAF/kr8hRKmAmavYjFonp/r1O/t2tH64aJ4CbNKldw8lw2mbRv+w8A9pQBte
ocH+zgBt2/F/JOA9W1PNmkhBppOyb5QqxR3pPKkoKT6FzGAnI+CeMQYgcwFfbs2B
2oXOvgcpleTqjzxOwa0GcoGRcD1q9mmUkB8xO59UtixsCjpA8FWtbnxa+rIgEhK+
uz4efL4TwJAPpxz/UIEcZW+pP4n8laoESPwYJTfisnBTVrN0jXim2XrsnLBfg14N
9S+oM9+ZcZvbTIdfgWjhS8MB4KJxFca5ERKpWjCwPKaRWmk+e6uzDNqecmgCBaVr
e2zwis4XVGJlPcdIEbLpGllNPtvwQrehmaX8F85CWUOnGvOH/K0w8LvUvm28VG56
NBTaYJPWsVtQ3F6SYLdi4TRdAE/9IJYBu9uHKKzR0CincOmOIPAHM/vxjWAGUCUR
B4g+nX9+SMjA1luyEFroaobrICXF511W+pgXVtB1syxTq7o5c4nQJC+zVQFrUZfr
pLwUfK71PzFrlEh46DhSE9w4x21YzD/AzFsEU6PHCQsw9tw86nwVcgbeaJuvLhBi
gwibZBrzs4zB8s4HNHzENj6Di109wknHar4JeiTJmsnXTKUISUS5UhNN4hFEUMgL
JXG5aslQt+eKiwdK8E9E3c4IhdgCNkuxgpM/vHNZnNbs7N/mH42vP24N56PqvL7B
ID+AgwrlexvBQ4WC84P2mlag39MXKmGk6dJh6XwlKltn4xwYaLCz9/9SCk5wyEHT
tjRh/+OPVs7E34RjTYi6+6m8rpzcipQwlQwCExjx3Yn4rbsewVKrUgibaLLTAElJ
3ILJdSrQNNywn00T2oZO3L0HW/rR5NqDToE8Pc3JOBqvAU2aBWleLyQAspVUUkV5
KhNmBKIll3A/mhQJ9CApiuxRX5MFzstiJwm/qbyewd5auG7IXJV1P3QbsE/Nj9Fm
IJ9b/S3unfhQ2ZcRxaf6rAg6gfrHxUGDPqY0i+atUCKEBnsdhMIknN5IX80ef6XE
ss430nWRen22KQDiLCiE/1fDdNAgLF+TZALlfaijtiJggYph+DUSScDD3k6p1037
iX7bGlhWmUPKDu9usXygMazv7oMude+70HGAeJaVH1WsZ1JAmuRIP4T3wbWji45u
2t6OWMDZ5weBUONJFPk7HYccdUtNdvi7D6JUSGPrNCIMGPLtOtX8Plpla1tb3NGv
WgwFHsTkulvpSWm6vSPVyZcAkzG67VwO/E46uWFj8A9Urmr6lsjNmCx753We0IQC
zqTbLmfPoTSDkaTfbuRlqvo+UzXYjnRWQrSu0RbagZy3njFwuniK0mFFpXK5e495
fF8ezBFV53xz6obzcmtZdayauYZkrub0z4Qc2Z+lILVsOvZJeO5vpcLdwUgN8K+W
w7fuIPZbzV7AsGjgb0rnQbkeVZhDtJnrzhOAzHrpgBRyH1J6VuhY0gY6a67n+GS0
8aki6NTaCtiYaszOiQ7pzahbNLv5acCti4QCuuduyUzVo86Fop12bfdMAEZ1yBYw
9y6JEC+Z/QdyFz7M999O0e7L7a6Z1dB76Mnx26gnIgTlA3gVQoCbYhOpR29/pcbu
pD+SjzN1qtzYjf4m27qk2bOJDunLr7toLpL60Cq7YIngJ/OPvGbSD0Fvfk5LJ+ov
rR3VwlgyFD+H4V7SJ1myXIjGlh8ArA+YysnNBWTmD5kopaXBEa0askimXbruqyjp
9ZaWjGJJ5C2AxApSlpJ305uGi16+MB9ImT936k7dZFjBhzew+aQcYQ2I4uywdTNx
Zo6QNloFL0F5eqDaHpD5UIUC9dpnNWdxVa/9yJ1X5JKOPfu50bLQhc+f0NTrQ8sH
f07Mml4E0/hib4tuX9CdsTbwfgL2Y3xxBjVshMYDNqkrzcRB8Zwsnx6d4Q+ZIKT2
YY3Ctyh/pwG0xywbKqtdpqGVDhmXcoS9PB4uClb9c0NVO+hSZTr4qsqJEm71KPYq
oLs8+b7ZWmFGx3LGpTw/LlnH61taTXfvz0MS9AeKse6iVdK8e2saauvfaJE9KKez
Uz+2fc/8ZcImyh51+9L22dBb4gpdHGZ1JHy+rxHpVOENNlgOGmEMV2iD4M3bAx86
VslfjeMF3GsyFaX7GmlMDSy2WmOa1Q8Lk6weV3t8VbBr9+4Far8V59kzH/CUTNEt
q2w4F5ocbODe1p3Mj9eWj7Mc1591qPXr9QhQfVMFO4byR/nAkxoqqd8V6zGn2X0v
CluudQVnlQhXlF5m75nBFfOsO2XqatVh9ykeGZySrthaxvHgQSKSKOgW1DH3NE6m
ucTEk8feREJY6Fb8CgIQ/7W/HYuvw+5k0UI3H578qiBGWrjHuAKxlwg+NQsI+BVA
dHEPEFv7qDgCLYP45j92nYx68ACo4xR4rqUUitvtZA6/Wm6++mTKMjkZMYtrEcZo
E5tjzV+jlZJkLp4C/L74hcOREwwtsT1FAu/UrH6YsGPWhHr/1XTS9ax8AIqT+wwZ
dPL8LT8kVaojy7RWmx7Z2TIskLxkplPUh2Z7mqsc10E3xRLIGHCk/rtZZo7ZRzIa
qmh0qa+SnpXAstFJhON/kRHq4mcdwIk8WJdFqEF6olbmPSCm8Qs2sL9WAgcCg5f6
qnU9/bcCY+tuVqzDHdoXOxsCBQ9me6kFvvDezX4E7XO0LimmPC3qBtNahOYhAusw
w1v4VxvD6ZuIsXVqZBjqH0LBc4NUgiEkUVr0KGrsb6cPuNj23JfA9+n8On/B34RE
0H2oaxPq7IQxDS9v3WRKsGi6WCCEbEO/9yEzqlbV2rVqowQM1vxNPczZ7KurJ37D
KS2UaSfzirP6kXtxhsl3OeRMUOnCM1fLopcaOV3YcJTB+bpPilCuKfGUencTumts
ZMqkdaYLjGGNL4CJOzm/xI/8KXTQ8puzZriffgGcFMnpq6wplTmKIssXZfdIyTUE
CgXRfg6AGSV89RoV6xP2MGXm3nAa/sTU2VdYAW7Hdy+DXMDPGO+XUriaqfEg80Xp
C73pOY+NmF2ygGkYHmk6QtaPqrQcEitBwTHUVJDaHID31mnAOVL5ndtc1t3Nx2ET
dqa5df3TZvBPX4OKWBRwkjWG5sXwQ5GNZ5uUc8l8R8JWmx4qxnTuZ7ByrOe02DKZ
CwX0Hi4usAeNsv3nDJSDOLbqVU1phFwjkDwm9F1llczSLm5NHB7NRbkMSQyA5Hxb
AoPbmpanapkPee5tWKxCu8JhkzMDOrELdAKVc7/cyxPd6ptkXwd5ihdaAgTtNqQ+
C8Ssfs6yKG0fDYh07Y8NV5Ozm5hzUcndEzQVzPx3ddScJYICsu2bC9ABTMwSKBkT
RiuKPTKyWFwhHUvANQJs5SjNATfAN6Kaq/l8SM+z6YrbLwyEzsFEGmhk6i1eHKqp
BUzbATg76jgN6QUBtb2bkRG+w2OWYBg6swBiyb1PgA+Zy8RK0lxD/x6WIxcGH5dS
ifL/I/XeYVlRtiwi7wuFGylu+GFSj/JhkJlr5+I6Mjwwrn+Z2c3BFILtmhhhVcz7
lZfXBf6AOSP7pnHkh65SKo4D01/ZPXbday+ZuPKC5K+oJyIlZpUgGCZ70RvKS3cp
eAvSywzbiPQDcw93bSl8iDWEcYLRVwrc3QknCg3mjUnljG+baGDUGj1/RKN4Xzxb
uGqZulGraLFDKxJcwtj1ZnjB2Mit8dxA52qa25UzAx1Y1HhLnoE2nOf6QLOtRrkj
MUrXfOJDrYx1GyqC/yNmfgXu8yI/RIeodros06hWfEe0eeu3RTlQ2/xXH3+rtQsi
aur9YwKJyz9SZf8P2r9YYs1jpTB6DLopNlkj+prDaeLUUgNbMroeIvYwgib38/HS
Zc2pHKZrwJxRdUHo0QMwF4aVC+35vcM1GrsEtSB0JI23xVR6oHwYY6Lv4PZ5Vz1L
48dljjbw/7uCaZwev824tO7DnXywV+zqIrpeW+QCnEGuLXzPccl9OkBI7DymcSfn
KFlwsP4nWsFFyXKJwlxh1eB1WLrH4mO7CtBUQWQEgytGwTPjnfUYcEcFAD6yIQgM
qIwoliu5luanNYbcRdLSECEZEDiTOMBP+C2VDLQcE836g8uvXXHZ7MSnxPtYIm+x
6v6NnsXOTlJMmjOdKZq4LIaHwrJtQvgb9oqNeHRLGMx9MaffpxECYIPVwnvyn/T7
GrmYezIIzpZo/AYlt0y22tdE1mqBz/T3zI41XDFQKFlOhSHZ8gVm0gHBQOncqERp
18LVJbUaNVyWsCZKoQxU4YGFg2mzNlaoVvZi2fbf38L+7JoC16q2FbTfqQpOJvp7
ZDJRfXCz4Ho2tH0rtqFN0XK3Jc6RLBAuK5vKzCD6E6n/XSCKfOsCCoVFH0mXY0bE
cCnUbyOgBQtEWDZCCvc8pFPzDhPTeZUZUCBGO+/CPW15m+5fOE3flMiuM7da16RG
PgCPkX2TzM5KujAGtwFl/hwzvtG4Np5CESsw0ZpKFKjeOFepAVIzzAcrqZ2jxpsM
Ok35mbX0bSD/ZzwWKGRxFcxBr6oP982TNJyPzi4NvkeA09GmdQBJmpKImxb01Kn5
krJjKUrRNE/hbF4Hnd3tqOvQHuHGQjI/bFurMQKlgpVUD7lsaAD/cjE+bdVuDIRS
f2MgsT3BShLoegozf9aNY9J0/SJPZGE/gi7XniK4q3Bf4grv/ULPZUHKpEnYwCgw
pTJIHDKfqbL1bQp8x+7aX6GNJlbEptNJl6NtDYglZ8Y4iVFZ4a4qjndq6vGk3WuL
dpgDLo8T3wrF4b6V8ugCoIPA5265BcTPfwGaYyWhPu6udZOUrjgThs5450d9s+Ex
ZrzNVB4LmKv4vHhGO3ZL0lTe6mxRmKa4nAZLQeZ3P7v1bC+G+jsc/VwG130v735i
99lVxDTf/GvmKoRQj6Fd72mKmSUjn+pdBZ+S3EmHxTbKi7RLyNuNZorzVFbkHKLH
68iWG2by5y9Z2iBOhDdRiAjUxZoVXeCnfilJFXiZdBJG+m9Y7PgeREqaEKAztb8M
lLU/aYReX7+5erdQ55Yt04lsde8MX30VG+vZiFuQtDDSaIfaFCalCgm6i7vbr6UW
41KliSEfu6gY9+BCk1NCiMDXZbVPHH1Qazil3XMY9jg52rDl7uh78MCd41ZSD63/
pL3fwfIEqtztx3lg6wYsaawzK8tbAjKwwSt8necQdLD3WeFhFOg0IregJrHyx02L
Ho4fhT/LBRogleYUSwoFBJlJKZOpTAYt/sgRz3STdyND9fBscQ8137RMwHnBiF5A
PLLrr/ou85VGHQvsr7A0NIk1ecAKKt6PPMBf8AtdTPawxAGK+VMzoH+7SkUToMYZ
C347X4FEQIE+YIZeMTZwUA1hqF9Qcps/E/LdsaVorsRjqwMg1TgPxrjqnZIkg327
7lFQhnyrQNA3QdmN0mZ4jhU+wchonNhuhRbxhPHbO5bRwYEZ71qe5eiGjimB6gQC
ipW4uTSqbZWESjsuVwoYC9VvSbygYMJFRfdYDfUM9AgE05sioFNYHQpncVDvP0Gh
UUFvvBg6DNeZe9vceVRM+xzwP97lSaJiKJpAoJpNXszyOkU7Em5S0WF13ZRhj5ju
A5tyOYGciGyAcmbYp3+SeRHG5/d+4sRM3Frb2luj0NxuBv7bCJ4jKYeKZgcGeyWg
hTc3j4wsjAPnAy5gradG/A3PvaDhEcTnYcSvjTXadPOejBw1mW3dQb7HkaHj4fYl
JGML6IYrSgw1olsfQ3N4ve6H+VxX0wTJFn+5R7l4/iVEUK73gd+aj2ThMcHEiSrl
2N+xzAmtyWg9h36Nz1eWC6aiVCqzxTboA5zz/WM6IFvnEWt823BKTbwOOkvgzqR7
PqPgwEZGvhiBh4fVB1OfDXoRatuRBXLeM2glOTOCAh4ZJTi+6CePb8T3ml6x3ZZw
64ywuvwsyImiQwDeD3pgYYp8XwWApBrU+CYIlklh7ZJDd3SpBEE5FCsoXBm6uQzS
Iz40eakFw499vJfCjKxXOH+32nkL2aEs8gmCIC9Wr0lgxzX1ZKXzUcZ7QmXtg9VY
AfHGXYAkJ7QFYBrFxYXpEGEEOTifVCE0HFlOxj6INwQB56UwVlLf9lMBOprhwef/
vRpKwGLwB/xcnhHB/ZUMgG/DdstK/6ScaO4rEObfVwMEtgyLwgGW/jVxlbzGaySg
+wssOVFVKmyXteMp13DNWr90dYllUpsy/K8vYsJZOWIuEpJXJcBBjaStB7wDHjlg
uqU/zbds/JHSIm2WbMD4vaTUtZH+GNdCIb5gyD2LtjE7uszvRvXuAej9rpMPSgyV
Axvu6hXug0LZcTJslZcbx83TceYrKqK8rfjEvQ8OnayqeXPU5hN5nWMEp/cNx5+p
L47KhCLfETbKgVAURRXG307SBYukx1E8DJLYPsJwOk2E28DQQfGKvKzdIzBk80oj
EGiW/KJYz55x2zk1ECb1ij4r5bRqWhaiK/HMN9911hAEVT6uE/FZDidBy91kE+Ss
zXDwIg9HaIZnpkRneNNe/XnNjnBCCRvfD+dOuZ7fJZKNaMa1WURlGw56oLa51Lt4
p6nIxMczgeL0uTzadTZ/ZPcRZcRi5cuEVOe8tCLECd/Apwc3sZ9wFzYornM/IA0A
R+T0NYVM0JNx6EVn5pl0MKK8gL1xXVnGLDscmGa39n/mQppZiBLYL7LlFmHttQKO
XUZX2vs2pVFFMuaAZb1/Acerc8G216ieHu9nZUFx0AIqTHY2bWADut0qDarUtZD0
uua9qzUBLAc0JA/IXHytvks3/FqGuSA7445laD4P7FbIVTkNomFAGbP3ya572vg5
FLHWic4mxwHUBbj7NUlsuD11dsCbPTrPF71PWf4CO1ZCHSmz+gdFJLAyOPu4H17I
Z2d3n418I4hBz75fxT9sDfqT/3OjQgiOAS2cug/xOjOOpSPm3F7qLLoVZs3HcLuj
IWa86f2F3isJUQehADkudnaIA5hPc2viltOWMqm0OP1WL673L7VCKqnBCdz7VYCB
7aYTGr7rkCJUHuozNlwt6cLevRJIpK6HPCX/oWopWYOzWh5GQ1cnaEecA7ao7OFe
R/8eNNPLNj6Xdkl8BKoCEDw+st6rymoSXWA53ptxiGIKNgXF2ou/oaEa3AQ9QVjK
WQLqdYQZoEnnyjQtam0DJ/J9Hi9TpmBtvj/pTpeGRbYhDQzfeuK4q/l57FmPeuvu
W67WDG3N1o10DdmUPgWaeeGncmYCNgA98/2QD7WbrozXM5EuBfrPK3KXYL1GqQj7
OlNtM7FrKSQMWO/gDGEddf3mR58z2WffUJXnyqaNF/7EuO0DoWh7TPmWLJXpaCS0
wW+v6SiWJAFiEZqzed0RBdJZzRubwgyPa2990YDXHNfH0dZDnubGQ5zibyj6r5m5
J/Hln72laJi1gx9Na2J5AfYmeJ6IXKVYZo3QMe5MVUhbUS0hgVNvGjxf2YMHxm0M
2YWMenpNYw/zMf/iUjP+Ypc9hZNO9q6okBo5WMtNQ6ERfuF9D28EgjF1qMMaCoVR
f9tLVDBHjIyKo2/I7Ol35A85nxdbFHa/LZSU1MpO0aXumm6wIpdR7O5Ev4AtT1Uc
GYb38jvSUB2tX2R8W5zdMgR7NedXFyk0CEKGyAToHnpw3OdPNjDL7Q1cmwZm5xcx
SA5ehF8qIDfxBxd5zpIEZBRlg4Hwc3FSOWyQ6Hlpl/8TiMwbo+S7i1tiCt3PElmf
18q9rD/YDzK36uCuO6w3Dr7rSlUQhE5Zln6wIIqpuq4ydLDKBF/OBzW1fYg2APWI
P1u+OwKMl/v0MZ9Umtdrt8SgkGYCDiTj16DkE/OORTPwUbCIHbvu/4x9dB/UYNXN
JjEViD3j77Q/tDtgVko/yGkwUUcfYM+GukcrdpOfcqv4ePNa4mgd1MuJIL4EOpE4
m4ZFB0LXmbdTKC3O/3gCPXCNL+UxjOuHfPPHcts03K8F94x7N1SgQ5g8ddC4LW1z
CD2sQnrGj2L2hQQi5iawsRhVomsKpc900olCqPGnSO5gSHNNu5f/GPwU9wUuBoNq
ggkXjfCsIV4bGGdudMU0I87BhX3/Gqecg/H6wKrgK92yJ0Hkcyvkdx66S4jbwdQ0
zd9d1sMHz1dGGUoeDQB8KHtLJI0YjEoXAvMPuDlulPg2r6lLyja9GcugY9cGrFG0
szdVzbT7jdg1S6CfWN+h8LgRnU5hcUv8sKvrPxhIzhSD4aybt2/DCdUZu30ZwXAM
hegIBBgjt2Q8HUboL1UdJYAsBKtrphOz/4K1wHO51xUM8752pkOsHZEY01eEPnj+
qV7wvF7KXeSlZVRJRuUjBwpxU3X6qsnWX/qO/2se+jK47xrFfiv1td0pAbUtXr4W
y/xAWH61cEfW6zHGd7OMAyCgcpck6DgPotrkFolx9VIReEfc54ZfsgrIlcFvNAb/
QzWsVuC5XRGe45CD+syfk6CjetlurTmoUkxibZ0CLc9dLIa9C0TzazqoNZ2w/TB1
uF0OLmM8rlqZChVhNv55yPgqdRJ2zu6o/lQdLjXRC5tZDj2+/mk9JfvRO7U5d1uj
PFOej5HVSy+03lrZkbdXhqNH8mYgD+bocXodbP6oGSyrysb3CXHIs1iqQHZVdDn+
hQWOsoPAaUX9tYn9Giz3w1q5EGFtjYstSWveskcAVm0mF5EoODMwr59oh8fR+5PX
cEElofkJPDQUWumgyChf7PxfO5qPxMEjLp514lYC7xowvbQjDFNkYkf7q/W5Hmam
gygHRkS6hIdv97NYekmqw0u/JHlKigjC1RwpNRS1LgP/TIW7OYj91pSylAYWdGFs
YRYuTvi/nTya/Xdt1QkA7992XM97Wd7XILpRP+VmoPShs9t8ybsYI/SLLDeGq0jp
t0ZSAL1WQG1B+yUIbzruFsoogCsUmp+TJSZJ09UW/zEIYVA3RrXkq/vzihAq2zKs
Yma1qDA6WvEaYcciD4KibAhZtwH9TqYMU8Kl/kPk0cKU4vPegdp/CEn+guN/+UKb
822Xfpo7AvMMbLDSxjSk/dH0ykOcmUzBe3K0MCtWlvFEA+UCi1/gR+HeYI0djgwl
VkOe30VMLjvGMTC0kqL+XriAFV94JI26pp4XrliUM8gX4Ry2Mal1hX1yBfyhZ9Z+
aHDJZMFbHJKxhsI7R/FQ7uEICWZaqzyaLjOkGwPikKlR4hZFpNWhESOSDjMjMk3v
wGVPuqP0jfx6V0QpUjYdqacigjqZ5NhEXpjnb0dxKf2FP37nDd/6KOUpT9CJM04k
Hdi7EOiOYYj+/KSLu9qMPhC6c6/jnYnpP5hpuWtjOirN3wrwZeKZpJvo01ZuQmim
Yjm+Hs+IqQiNqckAigad2+AOqnJs++WNDSwahpSO1o20OFXBAyp3hCOvTwyjQAtn
YyQXuQun6STIuER56UNx19D9Sxbgnf38QfB7z98Huc3pU5kPdxfap8RbZUYNeRvS
TqmygPyphxvXl4s18WKF7TbLp8daPERCuVvW7itVTTM8ED4gJwg9HFwXL/PTmaIN
fWNFI8p1sUThsGr6qI8/IYOlssClLdg1ExaWzXKm8yb8zr0Lc17SSaQmClKVKkN0
Pw4MJ9aITZJl3n/MDqX9/i3G6ea3OXJuXXoqWLPVC0vBCTNNxI4fJI5m+FuH2tnT
Qzdji+JtlQ94H4ijX2QaPsB6RRJMVSo//kfE3NQmqmoGiO2mwP8VR+T63B2Q2RM7
LiJtVV+DxjCRplse8YDWNLe30q2D/A+m8jz9SYF1YWmM4tsSYE4+1cA04QkiWS+H
s8M6j9MvE+SEAyrxF2qCUHkBVTel8ii7Tp5p5Z4sxgNxMGD3T5P3wK8607wRWluQ
yTzCdMiloiShSFU1C/qNGFAKBOSVVtr+EO17xZKFivhgVmXcI/Gfcag0CXeh3/Wr
ow7vjDo3Tq0zP6D0HuVhOWPPZSt0S7gc6OzaPEG/LibApmeXm4WUDvvw8ZLs5o7J
MraKclY9vHPt1B9k8zfkUIhGoxlEaFgg29qTzac2mT3Vjr290eeDegkPKTcGnwyR
2Sl72DbZD2O2J7eAfMYMZ9w4Q+vp8N8+N6b81PJZdpb/MuDvRCaxqeP4G4hEqztW
mjqHYg9bNpkJyZgJljWP4mlfumYUZ6qFGUVTeSFoevI8ZgQGkxCWMFZMUr9bfEoW
OqxyVvbOTPnmHVHhA6mtwlD8GnUvWeP2GoxbinQYwHwvhlUjQXqXaMa/pqBeG+Mk
3JWk9P8OxbTzUSbAaJqzLdQXhASK1IVjE2pBSoP4hRldF0oiUwsjWe0+Mqa6JwB/
OgWyO0KadIalLPJoOCRquRg23n3zDJwZdXVAO7C+6sxC9etMUGWrRqUQqR8lndHy
nbVz60mJrnjTYSdUUA8W3MvDYyGlJ3aCgt8sVh41lkMpkLkaJ2Q/tIvO/AGQJvtH
FZanCdhD7z3YffXWHO4cYbHBeUj6iYrwD9gjyV0sl/k9lZShXma3svtUMAf97QP/
SITcvre7qccol2v8fAYdn63vu0t7cxXX9M1HAOEMI4FBqFUOvGM5XgExpH7b0wXp
m4d3M2a0jEiIwX60dcz6UknVUb85nbXSC2z2nZm0M3yv8T+qxnC2EpR8ofvbRizW
xrjKIatzofeSCaCH2efMKn3WjwIk3Mlx4C7qnhBDXCJMEUQcATHi1YGd4hIlSDl0
HsGhlzmGYH93hb1Hr/YhyYdYfjc4m6FQhlae5T2/ft2eR1hyhBY7sgfUHfI5E8ZA
ii8aitk6tWv2WHgCvl73gihJb39XlTi7h8GFrD5KYTxN2cC+LImiNdzEa1f0UZw7
x69nTneBH+QVaAvgnDBvHeKztEA2qEfv3NHdljeWQmQ4ONIDAV+4gMiVTUdOc73z
V+L+pn4HN08t5opAvfg/Q8hDcn1+DoDPTVSl4VC4t6/9xcbzEPhxstJyxI77sGxs
CQuY6yqI7exu/08tX0srX1xMgVjanPnCS+MrJMIl2XXRmQ3OPpj4YILCe9c5UxuB
Fa3T08P/J/ZLIGSDxQxhzi5N/Bk+FFhnguzpua4F5mRjU2ErZaQ+kFEUclt74oM5
yRqpjWRO8syO4ZoTG9WlndfpgU0VVcrjMZZJGRgFHB4Z3tqVuEyo545LjLAhGnkb
TCEaeA+SaDXox4gGXlC0FRzF39Cr2xPMTdqXKWtDZjK7XSM1dM5/wCAf/b/RV6dc
RbnVkVwhGsVkCN62ag5/fgT71Zj9a/hNJo0KKOa8cakXmEjlnJvRLkDuiOdW4AVt
m8G4F521fObjkfzCHx7ojMem8jufBVpEyZzFUnHuPdvZGKoIpm0XuN9za2hAKZph
ODC84FlwONkjoPfsHiaVNyS2krLdiBB3SSvZCNVhWdSd/9CXQhOMle5FEmOv1V/u
wdyXImdsz70rtT2SKhAc3eA8AxevGlFNX9UEHRf67sLHavXWC31su6keXHnMi7Y3
ZFNtSja7KHQtPdjYGpjzpMl8FVs60DGRhOQ/76rGs70VbHOzz++waYWfRuaDWT+Y
4cJqyMRK9JdINdZekvAl86/hl3kU7e0XSUjw8xCczqpAkq7hD/03jzdlLIH/2Bns
3hnTpfLrcK8DXcnHIoPPG/HFmlLJUMwmOkx9RN3lKdWcPAatsDjLgPdqiLyzC1Lp
08rc+t2fZULsDHggzS9bXIwe86G9xJuQYbsRU33AKoSKKubnea1kdE036o2WS0cS
T6Am8LqNNPV8X/uTs5hQ2/Ubkc8xeCgyZ+1D9tea9olOm3FZbrWwwQIWk7LH8qBr
8bhElq9KCBN5hNCvP9dJVjR85IuK34+9noIK5LBGI1tUNvxcnIvnAlXYOEKOjGMB
gRti4Ba3S9vDgEcSuYmyUmTUUbhbx4+EKaDuS9illCWHpKYtCekP4Ep4agVouHxX
y8WGp9InbnswHM9gUXO1hxGOYetKJThi0YkkMk9nz8JwphmLzdAzzOg0cjcNkgEw
kt01atWXJURJpMI0tkpbDjBC/mRPUokYrmzLAmDcy9Wln2DVHm/PsPO16xbBzys+
77jvuLZ2Kjnn8fAS9sCSiZqF7txxAUUU2S1YUhHB/h0NW/EilLwMEzmlCBtjZocF
rtcz2eFmovzKvAw85cJc3OM866vVVRVJd6L1pazcQxbxdP8XA4W2tYikyOfVA5XM
dRQ+Q69KTEDTZ8NqakvLJUe2s1uf46uvDhYathow+lQojrZ0Kjc5uKGQa0jwTYA6
mqtKfda62fewkm/vPiBnvmCoC0mlYqan1a+j9G7GyAMNhacZwQeMTKAPOt8zNQ4X
F6JTzhwAfMC4T2mxtjMwefIJXyjbsIiL8rjKmsJ1yxy+yGVasB6tAe1k1GnZk3iY
oQc1gzF51oDv8TpghXfjrlYmPOZuN5oJTXODqFIeRz36dZDBo0lsP+2Hby8Zo7NJ
0C/L/Qj3QMYz1v5HhPcNTWPuwfQrI6u1vN+RgnBejCrq0MhPG1QfCn61dnHxHPGt
D8ADfmO6lmbZ0nDidU/fmAFsdglYsRTeqMaeXXwv+O8BjC6b2GE1oytAOXA7qKdS
yeZtvVmhjp3uczdO0TOihn4jBxs6nMZqi6yqviy3RlvEXreLu+TxhVJ0Ue/Mq0sP
prCtLHEvLR1ORadhf8wjhUiScyYUEH0ikze+fExnb7VkhVl5axyotDY33Sq+UaV6
4tEi8gxWK63NhDC9NvDG1GZvy5Va8mfwMaon/fOF+CzvMSSpyaNVEFIf6Kr2i56k
vDSAvk1E6v0X6nyZWMTiXOliW0FFkQBYh8hTPC8csArTiR5RzCTF3HHWbdh4lgnt
GTukNr8OF0qPx64cttKMhB33JGySeRPqtYyLJiGhJszgSkhVKEPVtj4VWsxiBjAf
1ZiBBjGScJP1Pseq3qdu8h5kaJtkb0HpXrgY5clanxVJHrCYhihtBHneidVv502w
zfgyLd/gE5NDVltJqJdc19wXjEB5iqk/IFmUJpbTh4cBlCWds/mp5cZ36at1cTyH
IccaaDc6cuCt7rdfMEwFudo9MWbLY19fSRQZo+ZKRaIxMZl0nwWvwsOrWY67l90a
J+fQ2f5791Jdf77Em3Ards1jmpcttV7sZaYKCYfGuyODWpo4UvAGNvbpg6jsBZ32
gH7S0196pPs99uoDtsw+Qut/eQpfumw3Dybmv1iq+PgejRCXR0IxGCu+Qugu2RJ9
fXDRVpgSvVY3opqdDwNyG241USBvvuQwRzitIa5ZjcoKDaYX3qtzbH58OHS3Paq2
ZN0Z1/FdwuVDO2YEt+ed6zl6e5JveA7QblZPah/Kb6cmIJia1oJAiigy1Z2ja4te
gNzcToU4haC6ZilqWSb99Os5VNmMQsDHOqSS5cFq8XnN7VmmoU2htdfGTzNu5qMm
Yq2Tx12VN+kE8tbdOgqDbbIJlZ+LZo1mmUzAFlfQ3uUpts9QGRA2B9X5dAg11MoF
MSQgPuyBuzjFLxeBidshp9hYReCus6Z/TUnq0I2xwLnYyeTcmfQdwH40qrmQk6E6
mRn+/5KoNBysOuf/e8c9pQHdL+FEkRsR8KlfpBbfSMUzc21PjYFdLInCZZo16p1j
g4HKqoKj76NtocT7osifgUNtI8RKZGGyctpXs/v4fIiz2vGSyIaMsrgmj6DdwY23
XW3X32LTI+YG+7+oofJHhcKQTvbY4izze0J5qWQ/JKIwFaNyXtOZue3ooBQFq51J
Ta2FgdEZ4YHZGmO9tjRQqvMOPWDsH3VAvEzkfa/n/N7q2zZdNiNlJXEnY5ZDlJnD
lG1DgRFP+zx+U+Pq9zmifpQA2tdgjwPDMOttNu+Ey+s4HKyDY8PwqGoNzT2STVjd
U1yFcM3/bo6RhQ7l0GunHkoQ/eHdwoOgJfBTOkNTdDJSfPhSIKKmeYvOVfGGNRnl
fCI4yDIQnD2ZFCjrHV9DAzthk1YUtyoHp+9dQP/tx/1pInrMqNdUbFsLb6mxSDIL
khka9R+2hkbaFodvkxHYXZ7BkEjEWYDyn2nN4GaOX6pmfj0k01gm9urqzY9oIeiP
vSQKpcUHD0D40f2xg1WVodTCTSJeT1SO38yqVcl7BeUgtlgFVeeyUaNo5Q5MAUKL
QaKZIG6gabEj5R9h3GhwfWHnX6zdqV0hdQ3Z+ePIx3fSlEYLUULvp5HF79Rr8475
yE0VgJsNVYQXKn0Vb17GataDVWF0+++SxilahTGwN1PVx8rTK7F3WOaeEPEYziz2
kZCCvebS8ExLF2Sl1vQ5OyqStYqOcga39btWCk9hlRRL9dpozaukTBZwQAFDCTG1
yWTKvcO0jGSsHoSFuiaI8XFFZbG56RweibStrNKnHJj/gk+2hyhIZYVtzstWub/y
d6DBrC/LU8qz07ODi2rbmoNnwmtMT7MpiAIkN84OWdevtPmb2Gs+YuWb7jb27x6G
nPrjMU263ukgzFKRdpuASfwyYz43oukv8b7qO5FA7O22Rukd8s3Fm3tuhkcNBHNI
uOvBHs2OXE/tT7a9oc1gbHv2RMiHqCkQ3ltPrYnHpjTb1l2yUogjZMTwQ26R6ikd
sxi+/Ho97SA69tjaQS97T/J1ZGIlEdMfPm2vXK7aMdwWLZG47VfeiZ/ZrK59ihXR
diCDq5BdnyZad+4RMEdhbA+/uE3k1sua+xfomY47zkXC6++6U4a0CFEVZUIseZ2E
+69de7oHZcpKRmXbsQSPip17RsFvEnNXilBHtd4P5fuRyuxZvp80oFxBiXBVih1D
mz/0i4E4wNgdOMXyxFragVsFjcC0sBuncgAXCmT9y1updh/w06eYronguUUAsnhD
3kNuzOmoLhtxzL9N2M/nqN3tAyQseHH6vgix200s4FYUw7EKp2sngNiTuwB9q/tb
KcHxi4CylIvDMzaJq9vNAT/2zuAkRt5vB9B5w50SnO1y6z4CAm/7uULF/9MQGr0N
1Xzvv1tWuiBmymJ1AG1/OHbBf7Dtl/ZV3iCc3qbWIWna760FY7XUAGxGXGTGYUcf
tv6V2PKEyjB3ar7VhdevIha+72PLposTQfd0SFky2Q5Medu+47P/Ti9pVVj49p3y
66cXZgxEhm+i+GGhFgsxu83sbxnWfrrutCAISue0YwVgQtSFMIzQdkpmp8gpaa/T
fmojY80Pk7o6Ja7AY0U3Z9mqPWHsT2QgzUmhbbJ4OY1qPy1xJby3P4TnZ9V9x5dR
zvDmR/LnsIxsIJd5cpcxCFnV1A1TuEevnOkmcn9IquJ49letExd4wmk8a66E20+W
k3puq4RZnQSYZsea9CgkdykIpHys9Yu4s0WkVar4ADhYQnOb1yB/TdO6i/wbxBCy
ExZNudqVeHPrlZKY/lejaOee5eyvB9iiOxulirGAnUpULRGzj9NnIH5HTdCcUnJM
Z9wzJh/Pv3Vf0/yqRMhmUK3rIgzpx3JKO5JHL02gP7qmHpAw/QDbQ/fo41lXlN3P
dsGyZK9dtLmPqKndo/wFEgQVl0xqrJopOoXrRRy4Z82oE8CzChw32K3PIxi5lhOl
9/k/WbirvSgusu0v/HITujwlAl6oq+bLKfcwXPbwpqfO5rFQdm/vSOElPI35b6u7
TVVxNvXKKvcFyo1HIz9NYRZ5s0W38QhsKKc2psKfKJU+GZL121YhgefSg8N+kpNH
8QWFIiV0FfF/Qa9UMU+Cy+YwHyRVcq6TE5uRHo9tlMhwta0WkG7x9/qZWo9hyhAi
wJSCActicS1sl6tRK+23HNoTQqhP9dwl0QJRCii4722yTqZRbNcp9lsA9N/1+EFl
D2pqdNF9szPhEF9BA5XUetrjj0fw36/7wsdhGZr347gg0ga97MYEBzGorVn+/VY2
CKVwd6brxr1tec+C6GX730JYTsOK/JJaALmrfghU6u+8fJ2lNj3m/8s0SnGp8pZe
8vuF6ojW3rhCNKHpqDUYEDLciwGkTIjC3Nv0pk3J/MsE+sHyWrbOum7ol4k3gnra
2F23LJDPoVayeucp6mlQlDzI9hckU7uqA3gzsGlVRiXQPY6AqzEi8TRugbY9sjGB
iOYDzMxDIEXl9jgnI5zwNXU5eZsI+BFwo7teDPwNLAUHx+3PrUMz58iQHVQQRElk
vH+Kg13vKh+10f3VJioJ0XFlyiglWbSEwcYUinagYLQ3ta/2VlwmbJoXNRxcqYpo
Dg9e4l+0Di4QZBBI30Pn/OyPlxaBp9hQLbG6Fq98R02to9zrWLQuUjs0su+U0t3O
PoACFCFfTdyXVxiGtuqu42cfPbc3pIZn0Y8dmuX+/D5345ZNZnVB3MsQ8h7xPQ/j
eq48hDPNe6uH0b2xV+utUWxxE7S0jiLi1hk4HuhVp95ys5LvSeJpIZCl/Td8nq3/
5jbAvkPS1Ti4sa1xj/nXfR7TsWgIctyET7r8Pu141OG4aEVuIUrtUsowoZtzPwqj
IbYnwWm57NMC9RS+AHOE/cpMmP3E/OWDELDAY9LOZOlql1ZvcSRBiF7qEPdCIoLF
UwrsBTqcJsZu1Mwg78Ck7dahW7FWNE2fHkvQ9EOp2hvqtNGPui+txFFk1XPUQszv
hHHW1qO4b31+OFGYuFoa3wds71ex0qs0VTRLGrViBg8oKIt6g+focsi9gXcIXv3o
9DaQhMp5MKGZ4mdr/Lyp6gSd2PhbaBJ1JnThyqy4Pc+PJErUOgTAKCSjCEpV+Ah4
ZgVSIwg+mpHiwhoYUReAA3ZDWT+js7uhZwbmHnE2GmKGG9yx6KCpFtgrxsG95dl6
RlIhOiL5YnnWHQQ8/vM4YP/ePkIx2Ebxv6rLaaCyh4+5rledsJ/jACQWxkxCfsfL
tWvPsYLm7MsRlH/Y65nNYfHFugfinMnvgum2rp6nLBvzBE52msy7rqS8UkTDo6u2
la/C6X3zUkCAT8DRlI8MWTlg6+SIv+J6nOHowXg5c4/JgyWsvxrNkgkgNlgyUtri
B30cdXfbEcSVIYWoyXWnY4HEPLSkr88JSYd+FxFdGgA6nC8AFK7FpuNZ8TsFVyZM
QyHltw5nflsPN1EXgfj2mMUyN16ZSnSi+fMA+J/Id0GuIg5zG0mmaY7mWoUojmg5
ur1qJyy4cEpoLk21HuFgNGkm6vhe/3OtxDr7uWbZXQ8TV5KWswBbamBt4hO00aKl
Qn7aVWZ1jvsLo2O+M75Eykzfrw+JR0vpCW8hm7cFe/FPqCqrfyhYeojieyjWSHD3
2E0xUzal1oDt0OVLZOG/nO/A7fYf3l6iscvlgf48KtflO8YWIgPDknEzpBWePfdk
vrNufYiG44gj6sUYO0hvsQ/gMvmlmYN/YKySVlwONA7h5C8vnfjkW20SmUizkN1e
70J2fyhmiJMV4UebFY88JaLyLLzwoovM12clqLSYWa0rgXk74hoHasAnLQCYjgzu
MTRWfGtQ54r6CHjzZbr3Kw14F0hPoruv2QqTbzL9IAuDIQnTTxsGNj6eF/TjBKIU
9ILLC/3yD2FsNhSvSRb3tV9hBKBV/AcgKMWdDmSUpricxzfQ9uZCzIaJ6Du8qmNo
+eoP8cLwrAZYiSuZVXGggs1Y3lXMl2fAeQceADoLvwC60rgfP4bR3nJKBh07/2xX
sqDRG2cOeLCFOpjpife+oMFhAkA2mtK8dMKUrvu80SMXoTHx2sC2EV3MwlIqwAEc
c79jD0N8hlLEuJElYK81NA50LYzaz0H9nhp1kwb9R4neCFCC+PO6zCvFz2RQ/4rb
xawiMe//8LWwTyUnmMxQ3JNCi2XCxBiL6c79vOUxl+tdB/0calaOlX5q+zgUNw+s
SZ6l5QaY4/CLE3hL6LaDSQ0zDiXOnrDSkVteGfRkzi4E5t1YMivQvh3hGVohd9Bg
0ts4e4FU/c9M3VMknqn9fRN3xiZSsmXLqJZbCk63ft91K0cKNABWbQVnUOCdXpWx
z5eQh4L4p1R4go5dzkW+8pkZfO2ln3TRwVX/22M+3BHuKKOGUQmUK1A+3cWrorgd
7zV3wv4eoUs4k0yiIg7ra7aX/bACfW9HaoZw3S3ieyJXJnvz10S1xuSvL3nL2t7B
kF05qZhBR4asGqfB+6cfmHlazesASVOOhTw+MBh0OWb+4ktUf6Amz+tGriul0vX8
Wyj8jzZ90CWlHyhx5Zf5Cbtrzi06Iz0FP+9kQLJ1YBiEXwRh+9nh6uRgfDPtJFvQ
l2+WZJRHJZHVEBwkCn30MK+/M0H2sV8ipeHKLRtUf/cdKh+72fV+VEkH5aAtcSEj
mqgeu9aPBGOEf4TvxOozTCopXyJzQZi0gkoH/5cD9YcgQSrNffK7R2rGfI2v3UP+
Rhb/qj8I9/xCzyfYEmIoi4S94yEIn8zWzPGsEBYVa1ZEdC0TlU501qdH1xK9TMtq
H95VaWmjIbaFM48modPezNHHlN4bL9pHXUfeUc9H658sL3iFK7swUwnhlnG46fiB
7ePfLBXhiPpsPVxUZhoG/VtuDfOg0dTeIdEapPmL6NTXhEmz8kVfC3JsI7svx0nN
cbSrvZ1TajRb3aQ1EjEnFN1ClI1Ju7vZAfh0UMhc7QY2EzrAwlPQEEu59pG+UZwO
zwz4WUHdzZeDEdaRecV/1X6pdqqfl9/Nvha08cLX9j9mf1GmMZs1peV2jzrkHNq+
4dqYPNYkmWVqY+E4OwBYbUTAQ0Q7U2Tk3iAcGVjnFBellrpZROwTdzFEiyoe//EC
Fsqge273EW+K4jz9lKOAEeR5jWXwaV/Stje9GQHKNMP9fFY9P1kxlECDZCkF3tlO
f8LrHrMoVkfNUIcdkLKn+A7XiICO/2lDJuKY0IeLbFF1dIP+Hq+LkmCNq1z80wh/
qRykIS9fq1dVWd1GD+EvTHmi7BDwBf/BcNDmzI0farpkgN8T7txBIewnUMhm7fK8
PY9r/ebXoAFZvefW11GKxyUrfNKuse1xO0nyy9MtFUYkAdSywTCS0++7CjpTtyex
4MX+lLqEVExd+8OTMMrbmC1AJy06IP3/tjhpG7n7eeqwGu+OhlT6nJzcwA7DM9/a
UywVlG1shiJ6UN4ictCdZ1NNZKq8t7GKaomdzcDlBo59KdwPX5b+rJLilzC0ffn5
dWIs7Vw/tAj9B/08QPmL7wEpapoER36ueE0diMDENade8wvbhaDQRC4OEaUyKdwc
JFoycnAebwHn0wYDG3Mg02OzO6bm12lbCKjOiR735HuKSQefRFiEwgWsEEnaXhdM
BkuIFTIljhGPvS2QqpX29lwqZgHXfUkuI0lTvTA9NXD1oA3W90RzCSzFGXPTztrN
62jlAqbNdnUKo35D3RzrJfXkm4ijqCtsbzMDvkt6FXQNopdYZBxod0FhBVtyrbkE
M48vC5btbJOvpnHkZO0os4tz7uMJvMgrWPkrjeK/6mrDcXqblN2EWq6BfEGycw08
76cmVTqwtkLxW9Dp1lMv9HAtK+PkUJRf2SMux3pdkQ0Beu30lyQgew6unX/l/7yO
+/0K9ZTh39BWdC++KYuiGkWknzBngI7r5vtoBR8Fnsgz0rvkQibmSePhJu/jfEly
Ilq588P09VZDGiLIJen4C/ZZpqo23ENiacHzHV8Km/rhjfq8HW9dzfeUY41a0Mru
wSttpAz81l+KQny8Hz8xFTROmFj7yzZJ0sAoVMKppqtctzfQsR/TEcBYVkxW3ULh
Utm7//uMzLUUoA76JXSMypDHwpPTXaWneEK+6AQd8YpyFV4s/jok2EBNWwbNgBOC
TCXW1R+Pq9CzArc4m3LPByIO44PDub26XgC6QGIQSHHe/smQOM4Oy3VPNYk/XSzt
mbfco1xD2dFWagUbstH6nMZmEFlEPefhwzCGIrTJc1J7gfQNPbJg02GQHGMeVUuV
hqLtczrBTaE/f+hto1k6aPvvD8KNB0N+MKV3Cp/GwKMpnR5KNb0X4XC+KZ1N8t8X
PFj/lHhdO7BmS1igMF0HhfeNoNI7nEnCjjgMSfSshtlddiRNGCS/ybMbnx0YuKge
9mxoo4kuqeyqWgPkxsev22IzoLZ3bAz0NB8eAYxKtFAcCIdYmyAkhDQYEVl4E595
a5nbFrAkNAvUhiNT0hgXjmCxl1Od/UnLwZSwRh8hC9OI5z6TjLiruKKR1bL4RbJz
a3mCQgNnF6pcYhR+sfD3P4b0f6tUqc71QNaq66EeZzApQ03ZRGEIttssus0mtxqp
KS5VS/MbtIpXxXWzsQN4SRKDNQCGEVFc+WVnI505eG1H/6xaG95ukhBdPbymwKMZ
x5xSuhu0Yr6AgL8GrSXgbq7ldIlYIBRa7RXhKSpjMlcJVYJAb9o95NXsuXxviZbM
QTCpSLgj+fZhDe7tOeM0nT9Bn0HBS8thFWh9cGpuou9AsdPikSIi1jv3ykLFBca5
9JRMrUoWkGaOKFWV/GmKb0uhNjEj7O00NKWx7TD9b0dIPi0HADPQQxhscMmA9cer
fZC3HnTG1sDzdxtHvC8HSZRBs2Jd7g/vG+UMPbvWgPFCyuvXLYvtkg8lrHjU5FOb
tNjw8CtKVXW3r5sVBKCAMlGSOzkd9KUMACkgNEmyZXJU+k+n68rT50pKrxyi0L5e
GIiDZdnQJQx+IAQhgGwYO888RqdAv3TzA9iEynlDevRsZZ+l6pnDN64DtT4OHO3s
QyYS344nItgQaO4Kf+i4rHHOhKPJWazwULRx+gpmmCOFS1lO7ikrRCD7mF3HSMFK
PlIavmiMM6JGXSXEqLxATMN4hOR//oMl3gpBBOtyNejI3eSPZbqLS82p4SetJoLr
Io1/bPU5r3u539EXR1z7fOPkpqGy1LQ6/hG04cfc1Pg0RI5yzEVOaOxwo5Yo+UCZ
HAMCvAE1Ladzedd5f+vAxZPzT5zrHoaM9i0dZRbsoxtP3WGeYkZjGGZlfLBvnaQJ
iIsEvY9WfxOsiuPBDuXtjBmyOa4fQZ5aOx8s/Ukadjx/GU9V7Lp/NMU5prKqHXn7
IdGsGhjUq9e3AnKgjK8ViJITlbJE5ije3f+Z369AVgSgfVgetf1Z/4fRkbYzBNwz
ENAO+rsHY9zXegagqEcONsEv+qnfHJf7T2CxyJY9HY483x3nVdzSQZBUkLDx7RM5
gJf9jdRuEWWdO0w4/d8OW6UBGOBZ2F/JC1Ar446QXjld7tFs957SGp5LiDH3eIw/
TmBPpngsj1aMRl1wGGNcYtTp4ysB8ryDGV+Yrx58YXZ6ttbSRv1gIMRtUVYBq0cm
JSh4yqxhFzqUmKsFfW7CeSHDqcj1Ay/ryKtetA7LuaVMbHsAOwdf5BLieslBZE7k
UTZjL3zSViXP9OgaMZ6iITHiDLPrT7YFBQq+En/LKNHOZYk1Cm9IeRtdUy4fSa71
32E01yPxtbv91Ku7lB0t0JjoG+WX+nSzWIuWekUKkqC8aA+6fxwoqBpcY4e9uyhN
yp7/X6mdFhfZdnDTTLUSM+UE2+jMsrwythAVM0h0Hmf8dcspQO0Sbi303g6npf4Z
5Prxd2nDmsSlc4MruYVLiWEUfs5wKCGf/EJ2arInRReRUM8LFP0NJ88kZ+ftQlUh
Sw8r6xi9SSKH2yCPbv54A4w4MwsVwiAuMsJ0CuMBGtRsb+EQXe0c3eLKmTSO2jjp
gqvqpX7WrGYl7qzkT8MvbDu/LUy9w3wtIM5zJ0w/oN1baoDtZDIzgMX3/huxqh4D
zKBeR85N55qFG2oUNKGiB2+rc5mT/5BX0QUZoCzQJXKjlEUEs9NkQ8KdX+mReuHG
AAGCgxB0rDSeQBob8WYHPudifJOv3tXtkEtm7R1+V05EHUKy9yUWHakm2kzUGjlo
nwdrtRD4O9ofGcyPsUULfWqLpzvuMjJv5jSoxjAJp5fCXBL9kaZSIcLAYALLQ8RD
me6u3MwGTvBspK8TV+Y2jXi13CTD92tL+wdZwx/RlLhEd9OTI9UFr2v/XdBgBU2B
WbqtyVnHSdJRNzFF0anroLavPXrkKTdoAiaKS8f5dojH4B4bFNPKDWFF32vkI75A
3GU8jxN47O4uQLuLjmge/wKWhN/XM/gE7fE5wY+aSBCMPwprL9kI4HxtskwVKN0c
Scs8cDz2bbwO7jypFp2Kgvz/UxAV2M0uveUaUPfU1LR5H1xmfxVDKeMNbWnLh8Si
/2SKyt/jLNH+gfF6w5VhHcKXq+z5HLrzQ0BQmqEGyUR3GhiAzMuxKdVijtlY6eJo
x5ATwemAjrgBNgMCeNzG1rSJ2x2cC4VU+ltfeLw1kxpbOLg7B2TAuu0R35f41DGk
HrgHh8zqbvEZqopRNH1Q3Bv5K4YE0GS/sLQ0I4zm2CKDV9s+pRz0jX8YKBmjIZwZ
ZbWasdeotKxZ2C78UG8oELmmZPP6i7iHng6ctR/vIVQO6VhfXewgyH0jROq5IAHK
ZHT5MbQGscneiCNgc7WU+vVzbdNhDkdS0wYnY2dkVcSVj/3rIGl6LeuwEN7+4g47
4EChcPuUOgKDevnPGbQ6jY8Q826GBTn49JFiE06Pu4Eie+OKeDvREStRu54Cq5FM
0F0wee6cD+4WoV/lFiKWbHOr5TTNJ+d+krEBSobTBsJ/jRe+0lXdwXalsTI8OIR1
6XVr32BnUV4IV/c4dIu7G9nGxoEKewGMS2Ge5Wql+e3/cxnwkk1zqKMBcldMrAgB
NJdUMGufifzcbTghaKlaCLskh+/qttJpl6s0A1bsQk/ERFxaBwr1dOtLTgug8AbX
RLDVs/rZBoGoz0rYdc4MmWUbVurlivfOOFY6wTMvin2KC7FfK0Q9QqcYOVX6TCCt
NsIjsNVAEB9wu+m8nX6MHNWZWLQgGteoOcqbOzekAmCy3cLevTZd+ocfLceGOXDd
lFFEmAN7O6hFVM8075ZzmnC8c7AmZH2ri9WVelRJ4kLlhdt/nMM7xVWQ9rW4a6Zu
an+M3lTJ+PaXesMuZN8A/v4F3XoAYI+NGnuZ/Jbr0F0I6Rw6F/kFMmaSzSvIcMzV
Ss3C8NAItqZrqx8i1hzyj3xKa+Qn6KgGjrirRCANUPaosyfeCtIp4zy7mc5Azd8P
xWkzTUcw3FT9I+5ny7kjrrz2A9I4lmCsJuaoFoyoQ1SRUJWizoweWI21DRqmO19S
8zocjhPl3BMJTbqVdF2XVsA3ifwsaswdEG06UbhDscBzA8jT+e5MCkBkKyqZ+I0C
XNUrR1w3WjwaDjHCwG6Jg6ESVIA/w4zZuJ9Ls2CwLPFbG+RoKHprjpxXi0YNMpeB
9mmU8mVC+4WzOU/ATzJKZWW/Qz4EshK8UquiO/Sjnvq/NydhPNQLBL5dfj8x/RqA
jkKXRrUj2ZKz42rFG0dLxCGDnBazvxLqvRrhUL7NDVFjb6qT/SKe+eDBrJKzvsRV
5o15E4a3IZCytb5fC2yn6xZCr1MN6kQqx5eAC3NgcSffZK1Sma5WzD6bEltT11/o
81ZfFKxcSzlbrf9onMnvPXpbblk7BTj9qpOn11hDYIdrugwoI+sov14lCd/nC76J
DEtjw7fHR225Xfl4iILBzibhRcaHKxd2l+Z/8IgsFD72tbgoD2wLVH8udMOeLI+D
S3wLaPi1oMSLS/aJiJrlUnA6Lw59bIi+7JgwixQ9H8gGsXslPCNBG7EGHemmXy4v
0X87GWzAoeYV1pYF3j2CGgd0H9AuqS8EZmesj8xfOsKf2MN4/oOU8I/W1LAJqNZ0
wJ9e6aih9ZdX7BUvVDnv9A2MLmJMSPgeXbCciSjcRdb5e5bWuy2KHA57i6DCG6+2
Idf/N23iuKGhpFbyzATRo1YVIcvX9r41TfxhiUbnsccxNnnNeokhcW8B33HyNXaB
Km24zZhOQR8ysxRl5sttezbc/z6DTM1xckQZMyezPsv+TxjkAXHYSobGrGXQ9H+v
5YbL1Ed0zh4zkJ0OXtlyFkGPau7XhqNlYo6KgWn5rIoOfpxG7y8lpQrIxQapxFsn
CsVslGaPvjjUx/IlRb1sRTveLPBGnShjesAuk8O7nByqzXu5qAhfO9IQfnfLYmM1
EuWw+a+hYe3HEzv9Ce0KrXYDYTRnwvyJexXzJ1rAIWloFaQnYJ4HxbXxg/6PojmX
r3U1h6kmsfOoj76u0jJikmpBdvU0n3ixsVF23KzLajdEOGVaqTaMT5qOBxZSqhSb
JF38nMlTaP4W0uJqmy0R2ERJ0rbE6K7pyLI79kOYcHTTr2qmXIR0J2omVSzOt6Vp
chMM086IZH1w2mGJA68f1liv1CExHVxetl9cBEHeMTVk3IysQ0zNBJuBC6qfQYBO
H4q9oQv/vevXYT6QgL2UJmY4s37SYx2NB6UKSu/SfiOzKFyy1wR07MiAMW4JAbmI
MW83aNDGAS9HtM7KDW8VD3SCUxoBoCd4dZ1BJmvSOlsU3UDola78BlcCknpTURgi
fFja4HcbMwm1l2Kn8ns4b/gr2TuGUBWiIpso2g1s/Z24/nTtOyQH2De/bfqOqtqn
wN9TNnQF5nMKAJAl/eDX3Bs6qQn9Eo+r1pLWu4M+G4iKeOyhvlY0uBSx7V6ASd6d
PIajVwDcwB7Tjsvtw3SpkyFNXyfrV29PA406JRXsHT2EZZUsKQyH6IufA9ztKLGg
1bFcd2eDqx04Vr6CRcC/1v69H/vdGSclDc5xEgenLERts9M1X0CAZrXAxC5c82EC
sSExqt6acmuWB6bK33p2h8s/KsGtyJG3q8LlvvP8GLHmA1+d3jNiW9DDrbOljpn+
Bjkwv1jaatkWi2GwAPtEDtpsho+OWnMB9dANwjWU+MR3Zj0dE9xQbkXS1bTR3neT
Tpn2luGSZ0A82xl41rEoD4apB8VTzpe+VZKcA356L4F+Amse/kAKiVY0bPSejb1C
t2dvTfBNAEyjNVa3GvUdQxZHONiMxOA+FPwo0EBuGE4e9LrsHGxG+SsnlL5F351o
tt6i7FeQgSmUPSymn6GXGj6rqhtAUdsEfBmCx9fxbQnCn38O0gx34B+76/EX7n2H
2YGcS/ewHvUckZTosfM0Oo+LnY7tk0tsWbOCEWHTkGB6sNX/eSRQqr2EXTGMxbWy
KYbJKCXgmUlpcJ4EKk1P7hKkBjM23rAHkgsr+4fvJSyCVpE1ShMwUa5y/idESxQc
ziBPAoHpBQbNMMqU/rjNGH9jvA2l4KLGPGrpfi3xxtPYYDcElATQz30Ge/lfpGbb
vjMP2mVKY9qgUdgi1Bsz0VRDSZhpB7HyUW84z2rjgCEED5VRnpaSxRJE6ttaYVQf
KsjHBZMKsPfrfl4FtLXHmhDAYw4zGcNPzc9EJmqu1dzINP+IKfIPRW4cflyV6zLa
nwRdz9SzQK54ijwD+dXYncjR5md0K7JeBf+MTBQU4WMedGGQuUDCFRxvR2Tjl+10
KZI/aYjiadYHMzGLlt1Xjavit60EiCuV494c+gdNrC9rz8fMgTMSZ8F0UZrtQ/z6
NU7GOY2Sb9zhOXcoauOx5w6+q+IxNqDTh15QLJlIZLvheWGzEcEgBcabg8712qio
3OBn89cXK8EfgYHoMkJd+KRRCaPfP5eIu1XnfRXKWonw3jOWnlu/m5bNbNwAKaA5
hGSbDY+2+tNxTEu0KhYfzFVsYSnoso1xEFSB8ZNTJYWuP/ZyNeIgoXRX4grRTIXD
5lMQrWj2XFqbrQ5ektZ/G77SYCfJO4jL9fjcdBYcMMpXm02N4axLF9dbDULK15FP
n2s4hHgtuYJ455SHXVRV9Rg0qVXQGdqpEAVf0UtKWuMKTDW0dH6XOPjZmmZYGcqp
vUfy5FN3OW02oF+ni2JESZ59baMOCwBXwVhP8BeUrxihYdAvF0ZWCFLD8bfD4WRE
ktfWMPy7X8/G9UJU1sBkIAqzimIg/uCoMMkVYqgPYGMy7kb3oQ5wJPKtUTcM3xHj
ajX7NmbP6c51jTiCJi+4vm1J/txQ0tdr9Nbp/ZEXdzcTqBwtH1NpgldHEWCVuDpO
LiedeD77TTlz61WWMAm0QxbIRSYE8Ts5hQupIocF06WVjuN/XdTFN/0xc/vEejhG
aMn9mqLlq/qnSPdA8LoRZGjjJoJfZVqGOB76iJm14vII82Zr5Xj1ttsgNV7EuxO6
vWK7AIMfQfhZAJWaXNgrwkl9uYhjgpWkaCweznk9YMfq7XNyz+EE7ulST2cPJ5Jd
4Wwdkx8ivRzKdhusKWhWDU6XggmqoA5soIiz482ElF15Q3IyIzQJr7AkNdaHBzzm
CyMhIxXIfDRSDycQfCqy8k/FMejC9+RJAfkronTPbOxpLN+w+K46GEFGXBBSrRwO
qQ+1H769tKh8zKTy4qnfryLVr0nqBI3ReZGtG2P5phxYKFkRaAD2g77ThhevF3Oi
FAk1lu5Lpafe1pwHjF30VpDmEk4hEpvdv0si12cNSsBg9FH8ZsizxSYfjL/tz9L+
1QELKEI6fdFq2sS+MVsQdirgVvBDT0BdTgOel52QP3sYN1YkQtcVLlj/d82cYUVa
izgYwiJz1m5SyiqMoU32x/0+gOglosC7rhJlRUDMzPEFzePywARYlEGzL96rLipC
kgte+I68NbeGSD2BBvV1aWgYOqBSOrFVuOvaHVb4Uw3NyuLRxKfOoYl3JUyMspx4
1rgmiTSRrYIhuGkgPeFFV8oXlpWJcuEHPJHorJlfp0hER06yqklZquHh7ug94Z3y
IIN8fzvLTMg3WY4DAkEB7rwyalSYrohqB41GouNd6uq+W803uTgE/1K1nwH1epMj
+qaDmDxIYl+P7QDUoJSRxjGNVBupofivSZ5AzK6m3IXWYMCxRNYqueJEKWB41TtP
xWb1x7zRidF7n88/s2RG3pWZSD1qhz5O9ZnmfJUj0G6jmtPIt1NKxFuEgEGKX7LF
AswvcfxmNvftCZR/A5IdmGWPhYh8321SvO/bOZ8x64SPZGTiVIPBom0hpmOvI0PH
2rM4stZWtJeQ0svX7jHdxowJNgJV8XERc8ixoQ85MGCgQfKdNQAG837bsF3qb2Sx
QM4Ye7bAg6EIev0kxbLOCmFBye7plhCEN7bWkGrctR31xGSo7BXQGk32+PFmbM8Q
vOe3x1iTfF2OkqP7PWiXJzDIlFSwEFeas/FelBrmEfnQyo3S0Q/axgw9XjwTQfBB
dDvGbhGOcS/vbCEOWGp63gZ6Rpfsw4qQu+SdB+NEKuPKu3SqZI3/lGlAHVfk1D1R
K6HRxCQydiI0kxQQLcC8p5wa64FH/SN0uD3zuIj4h1TsmbLwWdu9Cd4AxtefBHcC
Csh2hywmbirT6iIyGhol82059o0YTYLrk5+mDtbOHu2z9gXjJOX7zBOfg3qDssZt
Et71SdDGMCwRPe/1uIcT8YDdb+qgLD03gEiQK/Z++pq9R8Nfuzgve+21IZYyxini
wnr0qEGDemolGQ+zysmudEed1XXd2i6ouCo+cqLBxUsdllKz9l8pRgkeNJe33WVh
J3gJaVcRM26qXWbEWorBZiQBOHIcJsaoqJAAJEfeSKULBQlC6kofd8u2qHIXiWs/
az2ZxLqsOGrZKlg08qgzHkNwQS3Flxbv4VfR0Ygg5XIyiis3V9Pfk2VgqSgu8BAi
rP7lQPDzviHTUL5nggWafZHFmCUTdu+RWku7n4i+02xI4i0apAr+wpxGONZg1ZxT
x/cMfsJrMqVM8DTTFX3wn3Z+SPRIw8YWjwUoomZK6IdFMBjPjVUWls1QKjkVqxuk
vnKh3KIlwRIuedsQ3afY0LVvzknopitY9p1W2tICg3NEXUNG9zVo3EFgi8V5LjMG
INzbPOW33A0ZUGzHwjvVv9cBWSt07qhjlxoYsWZwnBkBUQwwIib+3nYtvnzo6ikB
HLeqIV3ImOnLPbYLswgFXzBTp8VDvpGRsT6uYtaIlLo2ExgxCYUuwpooXsh3QXZk
bz8yBkq5W4pEDSDxEhvgayVhm7hOeap3O+GmQJ37ph9LA+Xo7zCyywzb0dgewlLI
RpINEjsikxuqKnzZjYlXNRJRd1v4BkqLeyRgGlvxu9QoHJa/XpZlEyCnPPQAiqK5
bd8QzLvX7EsTjk7vNXp2mwuPt24chMt2dHV2go95RNU8MEUy150cHrTrA4kjJqWm
FNbRzHT7+t5g8BIXFNWanO/wzRQ7PZbskdLKQDXwUN8LjlMf4FgZ0ueeARwYqkOG
0qEGDdL/QiDD4mH9Tee8jTEy2NW6R7hYypt9ABQ7Jvi79MCr3HkTETalB5KnQo8u
l8FswYwKv6ymUad9mMicpX8e2j7ZgKG2JtriUcMm9q9q40zSflxVPk4moXjGvssC
yuBk/eJMqi2/WGK3zrPTpDrE70zz8Zl85/VXeSqjV9lnkv8LAqiHypPmTK5iwRMk
NMmiC/vzj2cjw6TxZZxuzzbP97E5UvsvXxXNVh7tXymqbnEZz/SF5wMv4s5DBMPP
nHez++VkxaPMfcaAGIzSxlit3cc2HZ3SVJee2FUqZMYpDPEhO+GBbSuR4Sg8uO36
lDEHG1Uz9DEYuiaONXTwU119F0yJg0gJD5ZGwNDhn0IOKaUigwjHJpOSBL8ipVk3
7OgO57xH0iTO26kqq6o7FwcHD16PfFd0sZkbEwyrpiduR/2MCQ58k3Xkk9gOv5fz
7r9sqtw8+ukAjpwrKADferRbkpIwRgRP5eAFoVJNJAECUYtPTQr/dXfhaYgtyd/k
cBIldt+WzNyhv/8TX2gAiHy9hQybRDDc0OI96fDKRmslWwv+OhyfiBWZPrk8fuud
5j11DsiohxEos5diEwP+0L4aNtR8iOt9w3QLelFydFoamfFOFgajBQXOH47fDAde
R+Rm6OLi0YpzFJvvsYLYzdC2qHVmP7wFeeISFOl8zr/A8pcWDthDp/gng+cpzCZt
oF/HAvTm/HJqUWvhy6IllO0n/faYHtVwSXj8NgvJPtk2NbpHe14rF+DF/tcgDwTX
nt3GDu5GYo5m3ODNjCmRJWI65FEM6TAECCJrrcRmNof4+C9WlvFFrEq+C6oIJSDt
70XqF1B2YZmnPZhm29LW723AU7Hq1N6qWDpSi6oY5GZ6h86peklnOKIiDKFQXkD3
O4w1Qcl095Uf1ngCATomuL15RO9LVeXxDFchnnScV3803V/nbAqd+5emRonhtluA
9m8gCd6/b9T41QOOZTej4JqomWAdjFZ/HHA6szkWWML2mdwxgsVnyiCwNyZqaGzk
UlUMCWYsufcWXy382A6RTJ5mrdwM+wtpxZ/Pjhq2QPAKSUhsGJRVLfTn9djQl/Rx
bgomFWhbP4ca4i9lHft7sy/bZy5f5ZH1Gg3kz/gh4qmOj8lWehM15/EDlR1Nkja2
kQSgkvSHd7X77xPOuPHHEUjSiSGWlrtV2M4RmfZIK3EG9ON5GccBL13f+NhZ4Te3
KREjeYtyyd1R9nO8przPP+MTQWgPXHqWoeOU+J1K3tgLG6iCrk7CRr8qcne/tLlD
gPH6ylzgj8pOTYMKsj59OQkjl20lrrU5DTwwDwqt3HGSsr95OdD9Nuc3i01I4tRf
KOYmKnDkuzlWcd9YNSN1Ztq9piTnVnA/GG83evTWD2zCMdEzRwZqw307xjMi/X88
HBCHVnEaJ6pPw7kBYsdiS897GUXQSWEsu4Aq411NJaUiCOe2I1BQvYStIHGU8dPa
85n5b7wg9hN6lt/xePYoFj9e9xr2bpk2SZ1OE7hl++BDPCTi31ZzdHNdO47ynweW
agcFoJBDLIv/LBtvDaHgZBA77YWpOa1+vw1P0nuAH4FQG7401xIzHBp1mwK09GNr
MezCEP1q99zi47XqpFgj80QxNe0B0wQewR3i7LSAJymjeqpV3c6QSZ6+k2edWUiB
cjhpXlXvvTKjy4/4QDRu5oqMyHnzaOiAhjhnKCX6RsTC96v4v973CXuxzbG/tkii
OvniqFHEmLGUilU0/a+r1eLdLZTeQWngdQxx0LGlVFv2m5JRiv4i9ZYDiLaxPkff
hvWO6hfRhsm5iI3PnpvV/xcru8Y6uBe6AtpeN9ujr8bK3bkArnYrh2eNVuAAM3OF
hXgmCXSCY+Uja+7CUfmhHjXAOj3jS//9/5fxUpKL3vMYRudi1K6/OVdHgUtFM/ab
1994M6aFYkgY/qotnRRqpRsnbm7FZojwwO7f+5FoVPQg4lJO9oNfxywrfkttZ+7f
356mIxk0LU8iJSWi6kgBEQJ9hGYXTTZzUSEA/CLeDbCSC+JqUAbmqYqFKtKU36E4
0KqzP4Km4cWrKHnP0uoYZF/cSrtHx5hs084HBcqKzEczTwPSxz5bEyzDU9Yy2+m/
Aaix5bBVoNNAo6iV9xT9a3PrUYomvyJDChD4qQUTvv8gsRCIr8HLNmIEtEnCatVq
YcoOe/yeZg91qT/dWpUh3DWpPsjUFAZkr51FO2BWOgWLDElPiEIZBTnkb8Hg5Gio
3Iw3LJltBVo6HWXGmW+u0A6aU7XAMnw1lIcpDwJjOgSVuEz5Nd7+x6bfoa4wTbDS
bbhv42ILPSrVfMNxDBOnpdXnJWGEzxcjNqRev6PRWwjn9mMQXQe4oyBKw7zx4KTU
SzApOQ6ERMna3k7boUn1AMQ3ZHyZ3hrMHNVtQkV7rDnx7dZkCQzapRun6pAReOnV
9gh1stVYjT6+QdQB3p7ccFpjAOA+miL7UdHazMkhPNiOniMUFb0B1wNx5+8MIinl
SyKztQH2abrVw6Mq2nkZlkwIzdnWCgnnqJvJkJ/xJP2/TbQ+ddW91yh/YeCL9jNR
NabD9+GYCbIwvob5a/HAUXIPCsQn1j+VQqsb8rE2puNBzlEaRLyfFsdcJe9NZkMP
zKrfjmDIqenrPhMbMJfYzqt8vBYCUHd8AycNg2BSYtp1uM4gnVV1WbdVSpBBkAl1
V2rJg5c+f4dUG/9aDWLJsistcC6Lt57jco1SRpKIQMufurgP0Lar2S91fqExle4V
AtU83C6ZavHUz4YAtpgntFW5cllQ31uGm4tgRbCZ3UpLuV3Z5O41EkwRUSpcGAEE
jIicvw8EGBLDmyTPabNPTZg/r9OwE4FEsA7Rv6l4z8K9zd/7lGeUltuqyErQVm0D
B6JEOJM/1Fz+TxLhJyQ3wr9bdWDNMN2UdBzXyqErolCurLuV5K0A7C7LKDI3MJGw
GzvDPM5S+9Wea71aoIyve/unjH9Fc/BTOQavZ5MJxQQReZwLEYxnhp9HFEnAsFv1
VXZ5cARbsjPIG+NkrPwmyLUoEgQ7+q+Z43O8EOIvKv2J7Uit+OL8U1/lRAW7JMd5
WYx0zDwmtEwR9Dfhk16o7Un3ZJ5y63Mpuk6Yd1hAUtxicKDfhOFKDpAAPhjr0zgK
3PMbdAqBDLvT1KXEKv7FMWNSityuegTowO/HGm+YYQNl3hRp9R4iyjMEjYd2TpOd
qwvZNwLboBcIDE65YoEHxN5bsfgEWR9YqQjKuTH8/lEOUEpEOU+penQgxB/2sYC+
vP5fzcXQ5iEI9MJhmx7DHRF/3FZliEoPZZkhdLO/PHEc+9B6fhNiWQhsxFydGIgL
BKA1wL7nNV7EGP6ctS99TihaHt21lx9jZUiJREWpdZnpbjdj9jZrVvP0ApLCKJB4
UQD357imugIKH9jpwmOvKkNq1KjJQ+TKBHV5LQW1ZP8yB1vypFKw633n210KJvbM
Zqvx8v00LMbYiA8guLirEV99HbF/iKZi/2qXxT4rqFrzopd6Mcp2lDk+EblprhJU
tIiH0BHBFBHckvbi74dn9vuJ7gVp/rPhxeyX+WffJnYLvOqB7broB0AXrET27ANi
jhTf06DeqnlBBVj0S9saP40hwAcqHc5K7LSqXdbzuMNot57/9AwG+zKvIpt0KKDY
0/oqF5VbPRZzyhN2v7fZr8eio/rolqSG4xvgkPY3OWGRUb1HlLN4sUbOjJisayml
3XeS+L/dpu4lIkM+Cc6BgUIv1NaLfUOR8foKPnZMWdOBnzEZ5s2K9pUbjywJi1A7
xy7+RSMfKIHdVNFI/8jDw1Rx02N2rZuN5OKL4F77AzEyOSmTD3qelsTVz1KlZQhv
YEf38uXEU4R+2+o5WeZVE5HR67JeqKgaXXBJGcjkpDKzEC5yXua8AmqqMHkk/IB5
2BLqt4AB35u7EHWZ3li3UNQyI7KFL8C3xYkQ3sif22Ga/ZFBpEi1DkOP+7zYjGlD
2XVvwDr7wGGmL0IjkyQ5i82PeVaNzm5vCQK2ueu3pRr/UWtnSSzTdHPEtCIdVpoe
zfvVoe/c8g7nJLYpmq6mw26hLTPQl3nirUH4EvP+Az6VaqgtOKMtnXDCIwBcUbt9
0J2VBTOKPCoa/Kr/Ei1fNZ1WHsBfjlqsYWez7aWwKAv8x7jePsizCjp3GVkMQdFg
NpuELFySEkqflp3DVjQBgdGV2raBiFAfF/J/U/modJhUxbUGjgP6asrcUGNm8D3I
zB3nKOo67epxGu/cP4/82AIxkJXQDd+9GgWgDengUv5XbhPWNNIKFn1MrCJ7G3OU
c61TiKz+/v1HhOSmlQDvqjrNjEWTOHvPtZQPU+WOQHwzmyeZZ9+HDPnx3onDLmEt
sRVVoVnLwjH8DqD0MjrCJ2JR6jtGp91pnNrt98se6+JmKK7No9D4u6+CbXuKhVls
K7eKyyAaEl9zQ14hQ9B909tF7Q8LkQI2Pp2jG3WBZs2pNvmOivNhrfFSnusqTUXA
yuDeChOJ1DdtTOgRCo4NH4l5A8Qw+f4CLNzfsoBhR5uawQDe6HlcVEgeTkX8aMY5
gTbgVQn6q095tzpAp1c2P7TAErXvVGejFMoroOeRcuM42NM9a9f2x1xPWzu8eQ+J
/ZsDXTuKHr2L2wA0Nj7p9ox3o+WoltCi7TSW6vtoCTcZCGQ7t+JdK7sIJCpIkpyt
gaO54iPjDdqwbES8K9BVnSsarXrMrTvkAy7Zq43i2DAeVLLRBPWqTB6KQWUaSATl
tCIhl7j/arSWkH66QYHfKaZaWaqOrFeFe9+a3IWh2R98wAUUKG4cPp7pJOjauC1L
5bxQ3XVNu6jdsYllb2AYoPxYGl/Pi25XZmYwoYaD/YeJ+6J4eppGH15JA6SSez6b
0aIwjzCx+2W3OeWiya8tg4w0UvVE6I6w5lPPHcJnSYAntkmFO66pW9dqRK3G5LJU
tnRr7Ei/PUCd0ikU1wa8VgKf64kBauEGclzzIa92ESAxvm0/WOadEPHPj99gV8ex
0a7rbQpKgZobWe6tT+kM9mAaQUSHcTmt0KR8+iD0zFOa8EZYKucIOINYXXWbjsHs
WOiJ6QDoV9KkeQlrRP3Hq4ylTf1Rbryw3vFSSHcz4fbVAaml6a0ilSYQ79F1YLug
RhLu7oWyIY6BBRZgLNaSHVCQyGuyYWmtGKUXP21rrxAuAfAxUhU85z4PNvHR6Bl6
kAVxL5yNSRQjcyJCAr3CyqFvAYHXYANhLTLcNRn834QnVtLD1tI8zfmbZiMtJ4sG
FU2/wjH80+WAZqoHORx5wFBSO3VcpCvnKcEJKmhvUb9viQ/IKF915KM/N477eYf0
AX/rXRtfVYMBqvpnw5Bmn2ZxKcAgGYHMHcocemQQ3RhfCW0oxAXiElyKwSYNe05+
hm0yGXmRonpC2Zb7Pvc4JhBXVcTiqX29x9Kih26HNuJn2Gxe/+IilPXpoCRHetnh
0xV38oVFSbauwF/9G3X0AqJk7T7f5wnflnS8Wmo1lmLl+ZpGZcL1OxWBZOfEL1gn
iBaYy3MTPEiUe12Nl+cGExNJLRkCm+3wkJ7qzir5LF7uaPcgXeXsTocqKd3aDAgT
BBjzrTa7zZPjuqfTk7ZBpwMOENsiGER72TMV4qAm/OPwvRfJClNdpumCSy4Nlbyl
3GpEjuOHKStTQNgz7cYqDti0GKmYJn98+5/mRQ9g7LglEN7TQ9Mx9E4wdH9EAOIu
I9sN54TMWJy/hPZ8aiGv5a/A5RmbiMnnslVhUKJrqYa8x0PnvQ9ilhlNjolQlTh2
t4YG3e1IJt4L7D/vWpy4/Ef/uyFSwMN3LJi/H2PoFg5EQPlj5Ke9GFq6Ov6ckyU3
LHwueV7ofFrTW1s4jjwHq68Prfk3MsC75VQK4uoPWBADsVl1Fdt2OTFrajpz5a03
L+2bgV93UiLug7ft/4DZeQfKxFD0X7vxeFPAcG5lmA6oZP29lcvxfP9rZn5TLgou
7zPCvvCAPXL/PADoTWjku3zv6zl1AMbliPI8slKXXIIggAzIuA2WsoKCT8amDcDV
UAE8ZqdrMXoLjAk0mR4K7VHO2vQvHRlVXbYQWK8PHp0FUUWYyAZNkFo5fV4qbjDD
QxAxmGxm3Cb4Cv+vwIi5x3OOXxVeY0zW309PlgTCCj1PfkiO1UUYDnQFcMZ0Do2F
jpLZDqZg5S4+JZioHuqkS8g2WRGAEJW/3HzC9qoaIEJlA/zsBHJZt3KQjb6PQQt4
kU0Nyqx4tnEJ/YHGqJB1yNyIQQkJE8hRwp+vkTCW4ONUUs2NplM93Wm+1yTRDvNY
X1qs5CDReK9LgYVXS8EcmXmbAZeHo+S+r+pLVobIM3oeXUMwpEakKngHOlU1UGFu
nSqIGSLPx3rs2IR7Nyk11Idjuzpkev0N0SYhfN4R3W65f63AuykZ5G9WoQEGnqoD
CYmJFuBhAh0P+Z7DkAaRUVkdz8Qhy1ZpcRRYIl00Xm1j4uZSCgAGF5Po9zHhikd5
468cFiI1kbzjVr9VkF18dgCRqY60P6t8Qok4Ll2aGSb5qDCgK1TNmnsAjlYLgw5j
mxjCvC9K/6n7reASsakwxiLluR+4pkLyhRCwDvLn2UrV/OLImJwkACCKwwmj+E++
YIkNRO0Mxhuip3FrFI3CjsGcvDOieCyIyzCmoRYPWLJEeV3ZwwobF35RFcIMzyOf
gc6Yu3+nH1xyxy5ktSrGO2sQLf4S2OJpbwWZ1tkYjyDjONTY6174sc0GMY2iRD7U
m7Y06MV6koolHX7Xj741wNGiDYk5bkuKlXbjSnYD+nmBCkwjgRrvShbQrw9BrqXD
oyuaOHNUUcIYt72NvJ4HLf32ip6nvjIN2LhOi0A2vDU9kKWJZHGX/2o2YRKdpv9n
lHhhmL0y4/e19nYRIXY54lq3TBwWNnoBdhtt5sjcfFDf5uo22FontFvmwHzAHuQg
l5gpq2PgmMXOJ9sjA6G4AN16jnXtOZpHls5BjM4umQ8pD45DY4TP4sK65jveCyEr
RxmxUZh4DRBSLIJqjMgztfkWj3bWiGJa0VjEi9b2LbaNaZ7+kcW3uGIHR2C/AnqZ
pm2mKg977pxgzMM+YakkKDhhKyobjuApGgFvije9n+hQuAOHHvX1UnaRUxiZYNC8
dKIOo4CviGnxvv9lRaRvCpemiUExkAkEKalRF4snfZj8C2LKQ4sh96/PH9eyVgqk
dFh/HvGrr6yH/Eak6xcow+u6uQZptopvcXkAzEV1B7YWTReFSjxcs1S+PdvJgezG
z4aBxL0PtwgqS0JFYQrexKPs6+Wb1pnH0YfY+1jb9MJK9J9vdLJ2seWFCcQdF3Zy
TlodoDVayhOqdag20+YUONgFUUTMySE76mITFgnxEwSQSlNBV3k4y5reJ8qher2I
trj2QLLSd3NCE2hCzdrz3xhINVq/L6ewauUa3uOpDyQc2c+3PQ6Pm6PCs1tX76KP
YrI0Zo6ozDwen0PL26Pb9qyNyEy7WMUmuMZ2gU2mDmaB8RGA3mmWtLme+sjpG2ec
/vwtJJi67sD+cpKN2skNJtl4v2/i6hO3S4ouGdaKkRPO2B6Nak1/Nlj1K92YLOJr
lTpebWYXIaWfRbbLdbYifoMDEA3os8J6qyZ3V/9w07o9Z3oMFDPm+yPDYnicOpCi
LCS6mfBoVQC1nw373stNRQie+M7XaBwsFSCWNJQU+m87N//1rX0fEixKgklueSLR
BFfulKZeHENQnyxjtJV9PPRpUnhznmqLKLY08uHVNQoO0flpLmpsoYyxvHUyLPzE
UhHiXdHrGAnne+5/0a/DYqq1vbIo6TDxYPnhMKDpH724juOs25sQuf7ISVE3R4Mo
/lxv1T/NQOyskOTsGkVBZoJDWFSbg6Z+xM/nkBxzMs82inFBTLIW5wfazPfSx7mj
KDpdbB2vJ49KGmV0a3fk1cf8e3RBczmeyv7mraKoFnvLTjialz/SVxpIr6+Dymor
WadYqP7MNPzJ2DxDj6a21QggXBKQkralQR5xlOT4J0bYTt2DidrpPMsvQwJWGMDn
XNqjH0lWOUxL79yXui7AftRZJr961BvwHl7vW9fr+m73K7C6umYSEwqy24KsPCKY
rP3qXCdchhLSMoLbTiHMx9ht5avNchHrUJLU0tT89khAuCfQlo9r0hloYGeztFm7
fAZO1AqMg4IjNDhyNOzqkK/YA9vwwUDBSYfD+bdFvgXBsGLBtDMEb+2f24LYGddN
gzRPCOKyfn6Rd53U1nJYyeyOSAQ5pIQXntkAycjoZIxIfo0s07S+NaprogbbNB4C
wbNpKvgL8bRHMLGxt71Q+6JT8Nl4T3lTowrvPv7qOVM6VPrGlLEwjnFKwcbCuohe
qR/alMdEdoRPzVBHrHTfP8wMczqvBJfcDS7dhO4OQPWH4hDbH+8dLxWDgk0QrmTm
EHuW8LbAG7BARs6j3207kfFWPuR0jZK/ZQomzSJgM1Pc0nHikNK5csxbb0txFndP
MOYN6u3WuagpAQNYwDYqDU2K43FD9qBenXsrUr6uVCJwLVdwxwghBRB0/SapGVf5
74C5mbf4dakJLrRRyS4PU+u+M+ZtD3tbgZ4XpxYpnAUxITXhymQjlcgSO6i1V0y8
0Vyfb6UOB99SDbiFNhDNonE13nH1TyffkAKQdeJG7i1LDsXTnJ5jl6wXnTSm6ZHl
oTnGGYlZeYZid7mJCwDnDJXfW6pa3qxVsdUm6ntC+jbUipUwhJOUuwth+ppSakpV
O6gX3rjHV3MUigQEM+Mn4oBUylQ+ij1eSdVLvAB9OZ509KpX+QDgXth2vYRlYAhn
d9X1iCvVPOfrKcjY+/skam7oEcA1qR/9KP1KQFYOtq44BsITjEfYGwZ/sOVkzJkC
C1n7TdpWJ1ILFevQla6Sf5B8P4zvfwVKe8FsoiHrj/dzoW3DGk2pY16v+n0Z06dD
eQ6mHwK+tIx2F9H3PAcCJVRrGRgC5qhxdZeO45ArynBCV4dIdCQnYW1CASYkW9ze
S+wuN7Gkgcs+IAo5j0ALg4EV3dbDSvlcToQ9CipbOszEWx3YPh5a1y4j9xzmrQhj
rkkVoK+6At6+DBg70iXOVXBhHP0Z1/e/NLVtxBzIsCoyEvmMU7+uVJteJA1PZpiH
i7L37y5VmUioMFmI3ULBAZmRwlQmjYJKRHuJNAUYo7rBIeDkXRqV5aElrofPI0Ov
5UW1I4E3W6js6Kh5U3Rem9gcKwJmyltMASeBE74xQ8IDuCGSgf/xCkw2lyKCJ+vW
6rBjJEcWGgaOWiyeM5yyOKuPHSQjhZHnL86mZ2XRUnG8r/W9rEO5bW8i/+3i+yPX
A9GpXq4BRwCzO79ay1ncl3+SJpLEoK33NJTbZgSyJxgKX+cuAxpMEn4QaZcbBNdN
bR6Vljr3hwSpPgtv0gDr2UGDiFWRQgX0PJRvIE/bWgaSHflIFmiVOvCj+95nRz70
gYS3lVWWyWtvu/Et7yrRrkL6g+LlQqdOQngqF08EJMIhw3c6sCBQoP2i61MeXLCD
ilXNiHYHAXPnGkRfRqMxgmKtMIaIqdBhoiRePASfXy4r68tJ9RtPzB6dBCjLocJA
lwLTDZWaiNcMT7Q86m6eYHriwOWdPbdCNu/Kj+EPrevWqzvHa7Ek9edZL7GTA3aB
Us40DYY34yh+VHqwbktrPUpRSXRRBo2ryKVf9tWWWMzd5J5SOYyVJR3eIzNKKY7n
9dSKU0Nc87h10/Wwf3ytRunF9rL9v+p04HyjkHvbSup2aOTsm9xQgOJFTEmwQUdh
b3gYg395ELmaRBSZ+tHWIgR1VtDxIBcsNeKTcg9itn5TRcMaSndzM1rS+v/d2Rf0
kd56FR0jZVkFz0xMiffjwsvWb0+1ckcBvAUjfoAZASv1dlmuxVDetpD9cHWVLqNO
8OYD0YvYyX/ikl8ADpnOn3kmiKgIIrXY+sC09zlGDRg+pzjbMwpXa+7TS5q5W6L3
o9R6IubavDX96n+84XBe2Put6sQJeOECYvy8m068HYdpSEIHQOc9E7vXpQK/6hER
56aQAg44+ClNGn+X1g9OYvwSdJJoiO4dALVxjwDVfuIgQwuLvpYr++5pHo3A0cAb
tRDvgpJQfWHk3xxU4hfAVOT3k1x0UbkUJxG75Vn0qZwMSMKxpojKBHwmAFYLJI4/
YeAe0Ct/OYshXarNVRpY6AqmivAlJfi06thknZ0XGRyA0kMFQQt3mMAtHFaR4I7j
RbdgRsaQfRB8bgb9RTkDswojxhsjMw7CX7zFai+l0SPI7Jih9xIgk7o0L3mEalYV
Iep+ZAsdGJzRSy28ASG1BMEesGe1XQocfKCdrQrHyuX0Agw7+IMH5XLjc4K2uhtE
O0jYMHMw6WdoBhS3qhuTIFI+rdzgjGxCA8UZiEAz22wRB19fHKuxJpju+JDUqYXe
XcZA4KvaZVCwne7diyP8r+IGHZXdZeeI1gZ26w1E4RBNTxSQZLuhAofpsczc2Yyx
vcZ5j/kfz4IP0vV51uQDT+3D/6TooOUdkDlyIodcFucFZhjACzcI2QI3/SQl4PbH
X2JnzWOS9tDEX67WY9g0C+wXw0xlb7L6f/4JC49Tb/QdFW9ZlBSfOg55rVTvWVId
+OTUINRnFj2WjoDozaD+7939R9zfKPKCvgQs9j1DGoXTFknXK6QPU0+E6yX/Ta1m
RxJ4Ray5QkAKxf4j7bBJeqbR5pHmOD03PjorWemThVFAWSudrIW6eM+5sbqiP/Es
JJ29frqL6ctpN/PdrIoR153qN8QC2Fnjzxnq6PFBAGn3rvnoNAftOCwi1xcLTXRa
3LTG7rTb3In9+QErH6EocrYk267yWW79k1KJbmP+pEky7Sd+CQ+TUos1zqKFsGEj
egA3l/E8BGWuLS4NnK4lOoYSH++QgEQ9MZribnYDXeWMN/yqH266r6tKjhumedsb
lXmPZnlZowakQh496oRF6WqQzVC3G9u7obmDnXoEtdYJUChVmgsmDXekGcBQw5wT
AuzVFQQRl1r06FNYC4/1eNdzz4B5rRwBuY/Uv8TBUBmXVlpkRsnYx/ewIfNKbFdH
/X7YhlVuZOrOcKHIU08gK4ma+bCmDclH0bKrmo0ljosw4tRsZwfNFqm8C46guH8b
02m7f5p4O//kOIXfuy/4fzM5e0Ef9gmqFlzd5q91/XCGCIPGz7rwFzajYmopewTh
ra/GRrKX7XRkVL8NBzzNPHb8p1/sLz9rrXBBa2BYiu5Nt/exF0CQRpbquyno45fi
Tro2ULsLccX88hqlKntk+xUIGM2jm66yZ3+zpYfB+AY3GPy7CEhdFfQF1lpF96WL
1ODKkEJP8zijH6n6/SJN400x/pB6N0rA9NoNA+Ogo97zd/tp8pDYqPRGa0Wlt3sz
qg3TRM8Z7WolwahI09nlgQnrg9Py3MaBUuzOLk2slucsf+kprrpghXUTBukWL/1P
1QWAJYhU5MMKFeKYDSFS0Ng5PSLZYqd7Mfn9XvawrOXMHDoJ4XAqwnmyV4dbuUiw
cILJXAOnGIrDmo3p03oHtxu+CXGs/QkUHeU764KFu6xMHxfybxU4LGvloRAfW9Hn
RYOzCvd0s3gAl8lUT/ZEOjrFdauB/Z0d7n3dBHkO6TkJZrIOSwfQE5EHc9OpQ6gp
4PSMAG4XxrrPI6CU7N2IxWuLOHT/3wQXc1ahaYw+xjb+CQEKzNSJnXe4QMehSQBZ
KfdPJT/ox52DbH9kIFs05PfReJ2UunW7Ajg+xgWmQ11J32XYqKXdiP3fjn6yUgt4
8wfK5kK1tuNKQOh46O8ShZNJm0Yd8tFFH7OHK5R77RxlNG04NU8ED+oR6iwupTkR
JmqRbTb9OGXKcLO2zWSJe9lrEMzlh7t1ZAK8QaFYzaukkG+wcS4u+hrdm1644gbX
gbUJ6/YkwFuuu1WiLpcsG7TAdStD3SE33nC+WxGeAtU5fSmm1grLQxudDqmND+s7
x8JrBqh5JUvv+EPOG+UPP0v0gXhKCFHGa42HYU5YxBSWoHmvIZA5FBG3tcOE8wdK
0J8kmZuGoEqWXx7+w7MaOD5GLfyTGi7ynejiL6ZW2FymtafbKJJb+0dbr5rnM7J6
xM7SE82+8ub/1zGxHIgeI2GluBp8QwuinctXpV5gmegLxeO/oM12Ife41DKe07Up
8TjHmuF+1JNRf5jrlUjyCr+ZQoeAh8K5mPkhFk5qAeEavBmNPIHF0sb7QelDcmTq
SfROwWeap3JGBWeMc1yt6Z9em3x//N+ZwbW0KNWnnzcl0yhwOKzswZ4DyiVxtZ1h
V8+T5xfPAg5LPsvsmPRyE7Xl0heHlOoqSyPGiUeCvi7Gmf3CIgQuXTI9kbIb+NeK
xnV3mRAlcoXO/zUguVzdxc0rhM+iHKriJ98U5/v6gzbDTlX4jfyZFJKU3pGL3ieq
Pt5xCA7WVx+HUnCS7ubx6kwwJIzYHQHmYcRRHciI80CztDRh/Cffr2UQShgjtXXs
ff7lUazxJzx1VvH4oXcWTRdMVvbSv9P/wY/Z2jZIXGAwDv14+KxGunyulA9UNqW0
V9i4Cq5z8dGaHb7NfrmlcGiDjt7v3yXnhKWR4LuSvKr6KnVIhLe2SPYjUOSu8ViZ
O/dfohlhwD9bZ/vO27FY9qxRHJN4vIz5vezw/7T/MDhlygVOyOf+aJEkDAB1HWE0
3HqQxZXW7Hy+bkEHQp1SdrD6za9Lc6D09BEjY5ahIr9IvhQG1wh2+9wt0Yj7Zh2D
A+nVeZ4UDDjoI43dglBvcyg7nRbfHQdPodJ+TseIZ9kugGxGa94riuVvu61MWKjN
2mSHNI+WgpRnHO7bP2oe7UoZdkkWIqqTcIuGYiVDK0ymCHnUT1cmGqtFo14AF14t
2To6htd23mwFAUHdsDS2IMUaXSHQx7WI/S7ucV/izOV3FF178cBKKTc0AcqpfJoF
MmnDCGxjnN9BUKUsa9sIMkQZHMo6+7YE9I5h2MmECUhx4VJcYJbWMECGN234fNBv
hhuk5NBLRYEm+d7dccXUmbgzi6lbb+QBR79lvRytlF034ZwR4TWIFUPliBz/UBZK
wR8RdzaDebrxEu69ctPkFACCc5BRpfU3GrQ2PnZF5IvH/mt+uqWL0ALAEV9V2WNh
0+bZAnTswLCIO48+7CAcCe5vCEBdtCMntsnF72TpuZaH9e7a7eyoZ10fV2QVMXwX
HJW2vGIKu2w81unPHOW6c6/PRs9lJTXG/yt2UlXhNBlM9K0SGGE8j7GalNv5s14+
g+u1Kt1INn3/gMng0u2KM33YQ1fFCBY6uy14sbAGDWTrmaXn7i/QVaMhPF0RiugJ
c1t0+dL9CnvNxHkKfnZsFecRUpzVjstqu/HjYZKZcYkbo1luLVmEbkbuXyYabJWK
lHt5yYv4ChpBWEcXn/aALGwZPv4hWWxdpm89YY4bu8kq+4BSPzxYhaDZoRSlhTCA
qYM0bj5AikuzZOp6GnN+eMakPtkxkWXMkybvrGdPXMDKGpIdXSxj5ewospMicj4X
9hp9GTSHk32BrFrctFrUs24MensoX6VjmWd1RvME1bvgyLbvJKzUuSD6g0JrpsjT
RCeCY9GqrAv9Z74BeSGhuCtX74f5OMBzT7WeKHbfp1KJHvZAG82kUaoVD8GvOrth
9ZQJbuHXLMKpgAAPtCspJlrM1f/AuxdYE/qHZkDkNSsPUFD9SKLx7a5HWR1QJu2q
cspp96psC5wEKSYlwQcUFxRHpNOCsXovHW1QOwD4E2zNCtfmmArduMkhMwzTpzsN
LMrLvmbuGC2KKECGDOzdFd/9eZERvZKYLUMzVQp7i69EcMwJhodJ8AzmCjjgKpaE
4c+B6fmwCRZRUbaFuyLpacgJZBadGsR13U7oNxqsMVLqonhqteogE69xJeV71NuD
sVm6Lzw2oYCamW6p6BjshjrWdMemqL5/5HKUOi0eBZNkevkgbE3onFz40hXaZtdB
08GNrWszoETLGCqq/lraxWHjxAhxnSnBahjdV3j61MurqIcbQK04rmJwmZOBYlim
1TrG3/Q9YHnytKguFOq9CusAqby/HPFmmlo5ZsEaPRDMQXDOIWYNYRevs4nu/ll6
GzCHxYpCjPj/x2FiqQ6tfAPvBWShvMuQvglKSUCanHD1XblAnX180o7myQWXVUVB
GfUxMZZYo2PxwopPD5o9lX/gJ3AJ8TrOnStOmIIDFsrVObxE5/jSPTwCfU+IDsWF
J+JLfpJUySVeahgbTJA90tZd/lhdBQQulFuv/D2M+tSan4ah/w7MEJ1kc4GgQ3k9
SeZ+B2nLqVcERwg0faiFdG0Kbyu6QGNzLpUKvjc3Wbole5hDRBQiOB2vCHepEnVH
Mg3+NRDhJpsMR7SWbeptrEFWQXoyvIreNcrqdCWKVFhAYVBFxQvr2fXC2WF0Duth
QA76phz1bUmpczSqfNhjTbZG6y3i6O7RlePDFL4ueTDLEhRPnwDEKsdXaRBJPYuL
TDgPlwADGn2kzsOIj6ZrO479rOjurVgDpHdfAR3o0nGGy6mIpQY6uZJkEsmGJ50e
Rqv9nuc8AfV8TQ+jJ2ThW63TsdiK/6iOQtONG6oquBpwlcETeb+nvhklk9vySlt1
KZxeXO/prm/d01OgLQp8Jn87uBGmMb+5VJTkDk5i//LuR5/AjMf0KkRYNnHsdqO0
S9q6lkazTbbQ/6fDZq1PDqvK/fZOhbn0fpg5tLp5uGJGvoS7dPOY7U469znMlZgz
YxZem9w0a3iCp4qAEWQhUcLodLs8cbsgwskB615CuBLatpBX1m5JYD2nXS93WQxb
yjt8SULxRfiaTH+/2YxMBdVIYWSacufGA/WMUKIpCJgL7DX9EGqjZFijPrBM+/jN
2qhg9gGTOALvYil4xKbUoTTaXOj0de93Nd9IRgd+/z+SegrLIMkEGhfrfecwiptA
eoUa8elvon34AJoQw0t1pfEww7TEhqS90MtgZLhPxK9HAYDGEh6Lyv+4X0JeNg/o
TqtQ0ma7YcnjPx7BrQL7M6+47SpH1YwfIVc3U309KN0kOCLHAVMDpCV2jabaATQ0
Stu9n4RPk7gJWrpR2J6VsL+mQAx6c7RqR6lfBwmW1U0rBZcA38lxTStwy3Kt2o/j
6boA2RtvZpMG5XIjdxYYXlMt8cvaiHjKFgJm5SExceQn8v0ocX7S79g5hP03+Tul
eK18JIKCRPOaFO+0WQHyAeYbiNreJuP69IpIN0S0fH+uHClQFjA+lkBfXT3/GWQs
ugYryFrk9PGdtgdtRSk+9jJzwr9U8b+pTSfjBrcYJ8OCVtFGsimW/TIhKVrtdlpZ
YX70zepmEfj4t27B4FdVeCxJNSZ4wwPWuwXrXvC1uTjqkDrZHe4yKQsFFmfKILik
OI2mV+xbZ5xpWVf1BpDAAx/jGwKozSqp9aJOLDUq7ZTcYmLL3HtQuRiO1e8OZAIG
Gvi3EY3LgEAhPuzB90M6iW0aMos6F+F4SSEI55qS6bDamLpof+2DhFoTaTeiC+ef
UHZZOI3cUT4KKFBIDoY6f4WDxVy2ikbSuu0183icSbq9CqRQYFdWmHtz0pJD5Aaq
wPimdicbPlXKG9uvLKwEhU+60mKRS1YkSeUrjqnYjd3pMXfRSyIRUn6Cj5ftEevn
vRfVITL4cD/NAzqaDEE6lvNlR4FCfxL/ctoy/GLjV+p+y6e9I8VNDY3lP8IniPKC
K3473XL+SLIH6r1KXAbTKVHDfnHjNUZcN5Xe6Dp6XZf19z5brb4TqPOnr4gDg1eV
p9dAGoGYjtOQaWiV26Fuxcf7vHi5IUMDcwwbNLNdcb2pdtB5GekHsaU5vzQUG9AD
Jzj6t+beuhPwjNacH6XoynETQEvNkwoNs0H/DCDkiFLWUU1bTlHx9shSkTEc48bs
ITFXv/cJIfPaWRJm00kKT1+/+Otwh8JIuscYZeigbAYJabaJPBuzPay8alGkYt3F
cFZxiV+XkPOnn8Tca2cxS0sJIaqDKsJYMvuU0BA3eUci4qZGKxmkwCkjOlVs8ihQ
a54QolgRff0lZMPHjCOYCsm0nDT3pzsO61SDYg8hmE45I414MTJaPoc6aLVg84J+
1OBYWNntaFm/9U6MYYTdj99zsXlBRzGXRs8X4ljbwr2iIjU512+A5+vA4icaGM0o
uWBnjao146j+8oDf6rvvmeknEmBMYdFN7GZCXyMdAcuymCga2z0WPpz3GoNhvt+y
BH1ep9KYX4f5dIMK+PFsINo60esnlUfFt7WVmpE42+HNA/DlCdOrkqvgetdxuxtt
6vPsl7egVd/QSyI4dBBDLhUHfM+/d0fYX+LMDvW5u0ixh2LzHOGbUKnccNSv+bKm
zncC6vjjt4In4Tze4PIGukVFMgS+b5fXJlETuPy4mVPvoJhPCOrR+3FyIfH19otp
s0KJfOo9Wlo7IBiS4ypUVGXkctdUe+3sG2kXxrVBBxruly0u+Kz8kfS44+TwvQyU
Ls+PT3Xe0ixtSzR1giZ841qFYCxRuXVFtGiTmalSxzTCnSwwMXFl5hFjfubbzltD
Th67ewFnEHJgi14nj1oKgmeif24nmpTOpYUendWbsXkigcdjK/41ZfG4Ibnx2UOY
gqVOS0uu5yGatuKwa8ToIiAXT3tP+/e71kh4xn1Yi+11wyQ9mVl9KmR1jYZkFQK6
rBTfCT5BLw3cFTys0DZeuJQj21EwS7nOpLSTtWxmB5c79ft/r1iUq6iDJD0HS/kI
5dTFOhVK9HpUkbVhFCnHJRB6DGkbMfxUKpGc6U/lo09pGtjCyCPhuKa0JH22t3L2
can6TWihGmHd1CVmfBfivbudi+aD0VNmMm8Qjp13Rx47y9PCFsDcuN2F8u4Sq9bO
zbkSccfk6u2acUQpZQTv2B/vLKxueHZXiWdJmf6GPoSX9QO76/GXjTh6fgzrUu/X
N2sYela4vXlwORQfjPQLDSxypkZ70st2D23o8I34D+A8K7JK/JxAocmvSe8B0Fn1
qgLSqHOKX0AWZv2PzqvSe4Bul4boqiDMgmvbHt8HNjj0EDKLfPB4hdiqBECOSVSm
bwh8XvKvxyXGtEt2MfMK0T3/RBJHO7DD68aHEZg+Ytx9Xj/RTYjLiIO12eygqRYz
kPjQDUoNxz2e/ki+2EgujK4O3m5HF6LG9A79dqVt7waLyPbGgC3FH0mJDI6fe/zz
vL4FtJv6/En/AdBgvY8MyymHPRaOeslVmptTiMV8PFb95amZ9iWDwZY1Zmt4lRNp
xrZEgKRSLzY5N1Q8/N1lE8OLt4m/AOWmbtUk8dK53EIFVUIk5xjqtQmbfjSEgiGo
wqB6YunPAZzYFfqYIHsDS0M/I1SEE0m+U6QQBPZzh5S41buUR5SMtponChXmQN2l
wrNHWnzhhSNM0XU/dERbnVq5kmY0xnjUwr68XmMPo6IxWH2F08iJ/62DJ1ayALag
9Tl1G0y5CwptZrqHApnG3s85rHl2HQn5/ky2o5OSjDETS9EOeH5PASglsVZg2XLk
rM5MTcJBwEJFWPRzYPHdR/k56f31P27u3+0ebyCfnXCtZMsBXnnbRTaTKgbLPBOW
K+grg12CbSMX8Zo/hVJgY5l7Dhd2h4ieRgjxQLK9v/9EEYZ56uNz1KefOAFh769g
vMVjqDuP6O93E3tBcpZOYrteWht5C/hBHzTYvVeplO9+FEWD18a72wTQarbeNFdN
8dmWa65OkOzHxSpJ5ZJRB6tDffFtt+56JvTUHJ8klyz6plnr2JziJiK5mAjJy/+J
Cc21qExK44iBeEsPrdi+p+cZD6F5eOdNv0sd/1Y6r7u7BDv5N5p3wNt1WHzrJ+OX
0FSCL5m5yw6NxmMaSQl/PZzeLCB22dx8bfU0Vnx9wj5+70lf1cyUISPbDQ7/cqiL
gWhDVkRF41Pb/AiK2MFv6qGJvyPYM6eY03NW01M4szJAx2thTshQbags0/EsBgCQ
laSHPpBMqNLjbH+suyXxtTgdEvMusOtu4wh+s2aM1UW+vtOoP5/8e0TnTWMmZnda
eMEJquc/qijDtX8Y0Jw1qDdSB4l4k7uMeT0SiAPyhvQbSTdkcLQKpgXlQxKv7KAM
z4VAHWXpMhz+rtm+EGIMRiAiCUWJwCnqORfzDN5H+/SeJmO/LqyPjTbF/DUKJaF2
p8/t9QsysacMPsEIBk1h1w20p4xTzSlrt2mwj4jd9AiAnK4o51Lab9iFUsijGW0B
YgA++ZPosBvv1BKeH5RrsPStrozS9ZSr3IOIrV5T0HwBXWeaF4MsHhG4uttoHENe
203J7xUfKSaMat096t8etlldG9Sy6+i3v7Mt2915g6FPOgRmqN7ziwjgGkppvude
h/Tmr0FbtPlsQwQaxt056yNhu4anOSZps6s5BiJQCGeZvHPTJioRAvmJphuoKlQG
N+gR7cbCHf28R/95eVeSFhRaAhM9BPE1p1I9mrdsHWVxPkIMNOSIDjOgrTkgirsK
dnHczLbNNKYtEctZ1ZqPFTmDHS7W1oGXmHmOvwmVnuw4IccZ+95J7KIHrJqohAyw
5FJRpOrRApu67yLltbWNqtB2xkHlPsAeGx2xnO+3l91nfZjdTAny/WLLLfreGp7A
wpo2aH2n29qdYv8C3Ckav+4NW0Jkn+tfm6neDTq3nrHKM63w3MMvuFD1vRWPyiUA
+9tKexjkI3F2m7ReiD2QHhnYy717xMDh05blD0n02Aip65o0hoZj4O+3Qfn6yFba
68RWaByzv1xWCoPmUjZTydEcTTSrCtbidtE2aphjl3ibztqCJrB/nsbRF7JvcQhO
ra1/KXOxowkGyMSn23Y+BnrWiO35BY9u0RoILq3x72CCo3TpaXaLglzx08O2Lbsx
Ccbg345kjMfJ9YuA5On4tvrY5ptoo/vdcdDIF28UzCSx/2fuludE5OoXvnzkt82Q
rovu34K3KHW3rutZR5zkgj0gmgnRlmSR2FbndzkQwiDGx/yh5OvHexbPIqsjOcZh
L8wSsXwSBhMwJsUuTyhimALlbHu3cSRqQ3MO5u0EOBRmJuGoTiS1CSncwiXgxO84
uX1p+TdFEoh5XQnNL4oRGMYXd/SwJS9EAsRfVp1/mvFGFUNGJVkoiXFCk75yAe4S
KKId1bN+/SA+hf8ItrY31q1SpStEcRAx8JpiHl7y9kf36eh8VH8atWVZYKvk3oUi
mJvTPC8m0F32zYiAsLdEnEAK7lyPoJHbjICmMMFlg9m/62mzLB4MMeYafFdOr1hs
tseZs7XRaqe5aiDdVayJQVEIisaMfxsWMTWkF3fsmxjbQCOyG7I2znlk9TWFDI4Q
pPdam/Mv6sZhIdaxrkyz0PP2Y9NO2MY6+6FKhBGqOeh/kc71/5Xd/2j7AHwN0zw/
EtRsUk2v1c/gYmzlAwaG5YaO5ZJ2/xPKAt2E2yBAVw4uGjmpNR0Xjd1qt17SHEW3
ttbVehvN/VgYei3A/yMmZvW2Y4F0rEEnVRa2JxVHDZEvkTECsITMaA1eryHFXG4/
J7F87eo9uN9JOPL+hRIbxQzMI0r/pGCZ6Qw+TO5CDHOE6ICyH8DNAU6WJDfVl2Kw
DiY+BlYcQ3tHV31csJOmkejXtRAFT88H3Eb4pTszG8Dw7VstocQ5EUdCwEf1i3wr
Ek7SZ6QPbxSRQ8MBggzvaHaVU64GaD2MpcVRaPLlnAWuI7DilhS9HU7I0JzuU0GA
Q14fNaPf7pqkfemwdfm/36V90oMty1VlIAHjiVjDo70zW8KrSsa7BpSCFqkCmElE
O/pCwOxdv2819GEVGXzw3Wf6oNQltcBEC5T+vLoN5k/ZSYThzirPDuF5onZCzYar
tmA6pBvehAfVoE75Pai+gRV9pV+DoTFXXG7vlDkBJlP1qmyy5OWKWXC46k0Iev5Z
fSIhSt65KD/WJnTkRXpig8eLWcdv8MaXC2GtWFg15b1/B8jKBfjOSh4sfDDeSK9X
D0v6nj+u4GOUzd+ckls8JJgjdt0KKkoWHZtD0dDxB3FRUuXPoTzfZGz3cnLNUYlV
HsX4nrOZX7rlpwDyRPCAIbufDngnRhhfAwInEtcvoDD3JWVnPYYdNtC5m2UQKXMr
jfAV5azlYjBibAXb1HYYyaxwHwrx4zMrYATVPM/+B3chWrowdELPxeDB4n8/iVFd
tKV44oLVo8zbXgRtrcYLJRC7MsegBvYgU6ERy6r69LWqJZxv4la7JR77V6f8c3/Z
wWCyzHME9HtCmj5qeHXoAKWRxo6KSqoLzFPNvPKn+DyI3oxSn/2qv7TGSwMSiCyX
2brrLPQExF866s7RwvnI9PRPhyQFIIliHiKlw7RojRamfJ2Z/PAJNJRSgqr1erer
FfvxY9/XtOe0rMhrqckk4rcMOyG3vFDn8P+6JLBr48eJ+0N1eKFq2oBmWBdI+lv5
VC/sfF0HEaFbPkwJOLcs/kO/ambDgXnqOvhcOUR1BD+PAF5C/c/JxcyJdX831l5z
kuefcpmpmCyZqIeapUuM1Ljsz7phnQXWn8mzJiARItwc1tsJFCJpAW9TbvEsdSrn
iNO2yxwEybALECAw9x9RD+xUWdrnOn37ZKqNiqyNioYwk7gKXrUcJ0E247YXe+1a
+DGKMp9NqEnh84UfiP3WGVusoPh9RLpWZGUin20IXvZl+UqQT3bhpQKW74ZHUrSp
odvFeNeUeQxp9qBaGrxWGxiuWodJArJoBVZbdXURSQOkWe/S09wffhdO5z3TbkQ9
rzxplJATksdKrvjHXGCR/Uq3IwiERGwoGp2K3boQGSvYk5rYPa2p0kvnI33r1fqt
zJ3FO0t6W7N8JVnorhQgEl2UZEdNmuCWW7J6tSkhSJob8Vi7FYW0wjGB8cl9dgfh
6/vl+Mn804T5X+cFUPKeJxFnnQziQibra198fa0Gd8muhfImBYICQfF1qJR5SwPW
0QAV8eDprAsYqH74B8IpO4XDHC/itC16Az5tW63yB1eEwiKve7EjH7+NyNZHHU71
7+5ROcuZEpLqk58/PGCPBuTmu7njg3d4TBXicxEBEWHOiwFGoBjRermtIlS18JsP
AO5CutxD9W7D2T0rErZciqqgnaMvmeOn/2fuz8vru0+9MEGw/VwBsg9g/30O9+/w
ORNmSkPWXSaH/KDqiAbNYW1GOmQ15h3aAliCmNv9GDTXOY3Fb6WE1HRHkZ0zmcYs
qw6u4IkpnRVf8DsvtFfI6grI4Jq0PBC7oHBf7YGQQo2ynLdqbtT+apgtzGZbNGq0
ueH48ErYyLKDvIijUTEVjBrGTNkcdRlkFgENKKwiJsHfXIXorVBf3HO18SSJC8I9
0JXJy4Ae5a2hc6UKTbhhNlo2OeaMhF1qsdOpvxsLAJzhhhffrWpmVTFuByDC5uH9
AyIeBBTbAw7owvY+7URNYE+TwiFU85IgTOdKQZmGR8zOIMUq/gQE5yPSbinOe7nU
oBAHj0GtoWONSud3En65xOdDHIWvBMlQjqqPaQj+fzZcps+myVTHKxLHVX6p09uW
z1ErsK/46CTO0tofm6ujs9f4gRjnDSxTiCtHiarjHb+hFg7h6qPfBJ2FLChuo+V6
nv2nWAicZx8/huf7ClRsqsKxFiuLEY+FpqQfIjWel+UpG4xW0JdRcxvX0Y5/vlfl
X9Yx+87MY3EkpNKXnVknlVfXolXp9AogWYGKtLbN5Z7S9P5xyHuAlU+rkIsR8Rz5
Lk/t9b/bntXmlFQhswA85RecWDn0W50+3iyk3JRS13XBrS64R90OwOwOoXXK0qOi
iQ4zyGJGVTlKChMzNPkt8Urtc/EyKwRiZCY5mXnyICPlzY8qjlmMzeyb5up6dyRb
tjA8k2iMgGzp78U0CQP/ENcLoTqY8/dOXA5X25vJ6Rfp/StYz9ujO4rsbDSx/6ks
EXP3M2jaOuy1bpss0dN56AIWNn8ZX23FSlrebCwPo3hulPmD/1LZGufesTE2LqQt
dEgq0MFOYQ3s4A+ERTSnpew8d8noXRbshz+KckrIlsgAp+z7iFx6XV9wdfyedCxs
iiQR9lOrBEtV2iZJoUP91zcwS1Nc2l8RbY8OoFfxeFDB2P9oKC360ZEbiJ8TK0QK
6JYKwD7QlZcNkFuNguMJZj/9mTxFkYbkpCAML3ussr/aEKDByf3cf0BLmhnrOTmJ
GcKkF+xck2BkyHqJvyZP6XwZaM8uK+g46YVVWeEj+tITMx2rC7OPP+BuJfLN4ZIC
Ym1ZHvadix4kp37ft+RYZJcmzd+Mvj3hAMoC7IBUcAZrJ0N1Ds0EXjLVLV3nhuNc
BqwPsTqsTo8xjEodHektT46h2aLHMMu49Ygn0O0ut7jO+zGMMl/K8IXlCffgrlaP
HpfAuPSK4FJn9AoLXDAEfzHKGrhZ0H7omgJlAVcJVzP7ev4qYBOZNxQuqoTbzPBo
HJKNuNBOcFurNdog5pLIS91cqQRrdu6yzy4m898D3D1pzr8annBijvG3tEs8OjVi
EXBILQsHbCYuPbxC8bGI6xHwAng42ohXSXvG3drUrKeXpt9sbVZFCCqH0iM7IkBX
w0imDpo/AAE2NAx+Fyrdy/wDTHOvyz4TuTAGgJK6DMKPgDqTDPn1emZ2zjHJ4jq1
TThLy4y1JdM9b5xZ6YnOIzgRe2LNFO2+UYulw/BeVNYj1M1B+d3ucBz3bAN6EiwC
SQBzlcXNTHOlmQN65I+PS2NL3QCRtv32mFLmnwwFNqxbkkPuB0cXWNBEOS380+/n
gjt+x7NDMTA6DO/Fd33GgAg0YhFgyEBuhXFYBF0Q2KjCj3xNEHx9AITPCAo1P/KB
PTvyBjotk4WPx5IWcqg1Q3IgoSPNZKt4gTBFXL64MKLwpIDRyD/BVuGPLWzUqJNO
kXewWTR0MxOzAk6g7ceuRhUjNvvEDWLU/SzBbc4NK30i7w2zvuw8Nu112Js3DUdB
eDHYxLClbMfFRFR1yu2nqr4MXEjklXwKVkG4ERz6820d3gdRSW6F5TKRNbsoZ9Fh
SFSy2bpXjamkvynDNCW7ysZCeYxD2/VdoQLnH4x28kSy2xjI9ao/6xU42LAmU4/g
9PzfU6+ZoIuzYqoSzRX2E+uABn+XhVbou82gsHhDvp+avLbJzytKRgug9iraxSLs
yjwUi8ROK/nNBex1BVY6cufcyU9Xl6+HwEq902CzBJEQqy/II4TvvTNC/BBcFqr0
TZcPyW/0t5hhDonL6KbFcVAe86RwVPmZFLyTrzP0T5eV7N2AsZI3P6iqMW54I4vm
v7vB9wluZmaAUoXLALwiWEslOrYAA0JMKQUmO2NIP3zkfyUNwBhrrQytx7eu3PjY
syd95M/B5VxlljIE8dD3Atbj4MawjT9rUjLG7N5YXCXlSkEdXsuCE3Oa0DhsZ/eg
5VQiTscy9mKviD7y82B2tq0ie+/EGa0wlhzitpXj1jHwyiQl5q3Ea5w5c4ycHWeP
n/0yezeecj6Lg0hpMm5+JCEMhVHAsEqn/CzddGYGLoleIGNZPWxk32YeIwRGWNXV
k3TVoTeRsO7u31ZllcEnQRJMGzRKdLT2gUWybbkqBmka6OpADTCjuc0gj+7KcFCL
sZGnNSKIfsHDEcWsKVdFj/0tlj7w6R45DMRMq2A2f9HnREDqi9kN0QzAGNeS4dxF
Pdj6eAT9UebIvClLJzarA1Sl8bNyYra+gMJVpxEL4SzGEPwJxmg1Wxz/s/ChgsDa
C9V/BiV24XWe/DFvcLU1cSMSoDQfTljg+jgqTPHwdCTvJsAuOZIEq9D/Thf2HEwE
QzbbtA/tEmNjAd2+10HTAPs7oI5aNcyYuwi3Ga1PAPgXVLWHB/VF+Xvv2rAMAe8r
WaIS+cAFEWjDKTGLsB8un2UmCvpDS1XSBquUIdqxeVJ1CyTYZ18iDAotQmTt+squ
eBijvpz1jXVYikwkL28DZMMIDOr1gsvKRVToxrTifFpXFJuAL8CL7F+Hz28/1K0R
be9i0nmwE9z7kuFeKK/Nyve6kHIWFEhn5sZ6nTT1RjV3jnVgQYXyJhk4h2RXDhRc
n67Tv6syz/GX5HFqWfx/cTHojeYcGiYUECPCKmaGHQ2kS9wJBAKuEZnoKmCE61MJ
M/xXuaCWDOKqa4UAtTmr/VwQmxzehxqfyqd72W+FkmCqpvprK7Q3bI9t0J6nSUXd
v4u+r/t9RmpPSmJDu5Wz7HYR/fgwoBiqcrRIF3LMGu0rDBoRmmXLdnk1xv0outaR
TE11Y1N80BXngMfStQpvLqdZMZp8VVFz/B6eQj3o+ZLmr8A67X1TvFGgglq7LmRd
2hBf329tGxgHKwsvx71WbM2iT0Qb+Z6T7CcmO01hAKqJRmnICrpDKrNSLWB2x8kk
WBx/R2hjlqyZYFoSjiQz5RTfBRuR7KE5Puyo9ykwpiCjQC3tfAUOpvKIdRSFvkUx
H4WAAkNPh2FXmDU79zNxzHDMBxfi8PaZMAfMbNxQqVp5Hhsx3oIO7Hl/xauE2acT
VoYdMOxaKQaUS2wKmG4NugcJa0jJx6qP/DPL9T6rzMmVYR1ikPgvaz9wPmQW1sdk
/Jr4cgwNQRLZC2xWAzIZw+oYJcxDs920kQgXJs+MRZ4/Q/T6R3zjF4rk82c9G1bs
gTkQqBkvx61p2Sm0o/WWwjmgj5CpzCcuKfOwBVdVJiqkKxDQ+WS1Th7dIgjp7KIk
enBSuWN3MitmZBHlqX2Bm6BH3zBZaja6SiHqepPUj9lIq8WxxZ6B1U4fwZUDfwul
MBlUuoHe3Bt301kQbo03bVHeVKnZr9dES52NSNRLB6y5Qjspj+GXR0BcMi9SrhY+
q+Puug/GBwan3/gfaTsVhNhIAxn4v8oSQgl+iX+ZV8O2vrKDMI3p/lOUISFydPcQ
0scF8+g6+STW8ou/mCRw4xDP9QDpcxPoU9aOLAcKmspSzrQ1oJmpZSKlQ35Plix4
hxCkzzarwsTc8rCZIY3heJrpykceK4+ZwNKhAcHbwTKZhxctItFoECKYqKK3n5fq
RqBxEN0lW5GzMk4xkpnM9OGmJhhbzGCg7994U48Wrlw8gGb6m2oaIjhdJ+GVHieB
pbnuk5u4hY7tVt0h5dtajByKav4qmQn+L9nFAk2aqCiwZXChYhMvSzQXayhs/fBE
b0dRW1g4VVtinb0ZYF59+Ikl00P2v7o7v9RHfAz0vSNas13VBlTKElzNsGP9L8tO
uqdZxjbYeuynQryGbwmjRaVpvloraa2pSTaufh1Auqp7AipNLZPP6QACpxIVV6qT
zywff0I1p3v7/zHAluOGIcMN20BkPk7sbaejruelV0du46v9zeZn2ngu3OzEy4Gp
ERId5PZktLSmCGBxWlWiMTv8a+NQUasKjQDqumKYiK9h5U5H1ch9drCAHfas4Xsh
hDxNmkctXIWrnoQ7VCnwo6Kp37gW+6EWeoeGIWFf47VwphmmdNr+cJvEnCuh8o73
CK1DasbTBDCLV4bTx70LJu8QAbPu+zDC4bfYgO30C2cxRl2lhRynH5dWBZ8vRlcs
qRXmPl3c9SD+HAI55VE4ftsqTZ0ct8OkrjuESp5OK6ft3cc4S8bzGOY8KHJ/FBa2
rKjGgjG/i93idAKnTcs6uVBNLKdr8yb2LoiUKcn11ih2H4nnsobS6l1ski6bpnko
7s1g7DScjzkQ8DRkDDLDK6ia+w30RnoLC8qC0njfLtICZJHM1KWGOHMRSBIabIy8
biCDDmD2SihVLnHNjYZRFcwdPy7Z3b9lB8PoB+OjY7CXUyjiUCJ8mlP4SS//dVhi
Rkroxg0l2SEsFNz0NZ8Bw64z2Zqaxmk/7H5+5ubGOpw9znEb2x0bWHR6hmZ9FK5Q
+F7wF7gItkvzu3Q73rt+JxSrQ4v/w+rnna5/by1w+bcKkO+q/kWEBGr1hL+Q9Zpc
VIjDfpQx145ZcrCCH+iRzdtyjBNviCkPy5zLxM1XyC37pV+RaI5X00HuQS+/E6tK
6sVR64gKV2sKpcOskiwf5LHCtiebcAjYZ/usZ/xJWFgOA3+vocMs+rAlI4x8hPtW
mBJUnwSzIf0+NZh8T414rMILeSKDZAv3FGSc3zdXQ0qFcE1AER34nfPrpoMIvnTg
1s7XJHuqDBKcDgRrXsPbGuKIubR/r3UKKHogB7aPrlkRCPAPbsG37F2/T8axmi+X
QdbdIqcTHp6JOxxUQcdsMpiev33oPDWQf3cN8+wISTjw/0YSlH90JPoRvABz/XSd
63hDMG9299HOUZ3uK3ZCwbRRBxnq69n6VUQL6MWBLXvsj2AULGtgy2TcKO3V697x
RGRl75MVbwRFFDhpXe3PJdoW3S+ezN2+AdkUHREUgSJ52C58tQ3DueEywYgXc+5C
LjbSqiRSyic/2zjDpvBtA2NvjGULGQiwKzgWQwsVOgd2IspNuVuclbQjI7Qwg3MT
PUDHwLudWXZUIE2hB8Jj5QtSZfe8+gXgtOFLH46ftdVNGTZUDzvOpghjEc0VtIzo
HKhTQ+IWPpinfae8MBAIaWmviWgqFs8vaDqo51sYJ+MX5yfP5XOPLjuJaFNF5qXj
U/Dr/oVpTcyTP28RhspcRBMCY/FMaxfBZsHT/jF5o2uOSRjY8A2sf9vvG9nClROV
NU19Zk2ZfF+QmmIYfFN6LMRM/P7iN4AibcrkTRIpFCqRYn4EmW6jUlWHuWdPsYJW
4IMXowCS4NbLn+ZNlW4FbNfNA0gKKc+3sznllTux8pVUiIJZ6zEGPBdaxuTZ1FIv
Mvh+FzsE/CTaPEwQaXhLEaZRwSnOc5jGIJWfXriM+9WDrrc3YhqbG1J9cwhXtgAt
RDMwQCgqPf9WuB0F5XHgMdBROB0QqqjCaUf+wtAg1t63SQxO17e73D2CzcFyx4Ie
IOJ9riY3xRth8He5E/PexDHqwzoCjfAgR08mkNgi3OiqIVcPggKYGWk+oSA+g49A
CkkK4qkOC5Mv9RZ61au3tgElWaGzsEiGfVexbmFT9vn+l2Fky2Fi6OxRqIoMg3YM
sdo9C5vqnrD0Z4pS2pAB4m/hzkFSrKuMZaMxWZyqBdplIvupmH4gRlEtPd+2SSRo
rFqWMbPaVin5A0iYyiomKyH6al59YMcuLZGmXJBmwTydcN3rveSsCM+mjrTGueZ3
PkCVk0x+AVJ6uuM3nlcL4lfnZxM6+EjDnNAB4xTfaVNK9k3nO8BSMW+FFsmyaEXu
r5i3Y9/7UggoZ4dfQLKoMOO/rR1NlBEOjL2SfbDabA2kW4Ml+c6wnvKUWLeh+lm7
Xt/vLaLsq1EKn9YGBLo4ZppFbOqh0pCPuAdgSKe+gJ/0v+0VyKtkZ2ByQwkseYgv
x28O7PJVIRvVp2wjR77ReclAJqljm7rorNMBMnLcHJVotuLyVrm7Koa9S0SnlwU5
1qQMw2hc8dI6tcf7V6Py6aDP60Pbxt8Pdv1zYsD4SvAirAWh9Z/o0b7XwJbmenYZ
zEWk8+vcVOVtMSDq5vtQsx7DVPvE7lvhiAtlM08LiDCrR3NROd+Ds+SHv0YZowDQ
c5Ji7sDGJCfRB55WaF8og2Asjy1DOyWNUrA1Ep0VnbOUFt7OhGJuWM2DAMKmpexh
Ch3B6oHg4xw/tO8QCKqxYg3gcTM/xow785ErD2XJnl7zZMkC4hEdzupJ3wXPByeM
zfp0J0iVeoqTwufdCGZCCkZkrhAQerq2oNlu+pStxZLX0zEPh4doILk7j39VxoYf
qj3T02zMfMDhPyvo0lb+zJEJSYVYrqRXVSXUVCo9iwvD2tc6eUorH0TBFNA6vXF0
zbLaVThdBDIm4xqecC52CoW80BkLGOjbKUdXc4IK7fAMClmI3GGfavC2IS8hzTCZ
xqd4NI/kQy480RcKl3MsSgXuXdT/47mVJBqZwsJrZ+IQquNcCfTjvSQZYodGQWYO
is1JkHumgWlpMLBkz7+l8OuGdB1oxHXv6miZL3kRohAKuVj5BvCAACmXtjcVGMEv
i5ecn5QhU77YQHZL1Fk+GbeGtVM9znq9Z6Uny6qyVmugus4KUR+BasMkm+TSPCpc
0SWd6LX7y8jOgqFueLv39Jkwz5kRnygbPxARvQdCOHnPG0Na9rNNgF4o6JtOvF8n
UvWQIyrgJEr+Db3FrcunnJZrO6mam/CzE1LnrZ1p1/QxHVz1vdwqoAcWlXRoiM36
0s4cKR0YBD+Ko6yZkwBZdMeaUoz5eIlIL1q3GjBaQNgVRvSskv9NGVp8ssZpDnHL
eYHE3nvs3EjA6S3QMVR9n5BnGVunIjalafuPvM30LMloMa1cBp5a8MOvcN0CCPgm
UIJ6y8fzIJeilrNz3eJyHNyUbnaHK5BsCZD23lfsRbWC7k3bHZHfF+dz1xm1RUxl
5ve5g02d1rCns7WGWRwc14dP9FWjKz2ytyVxtqJu52hkDZPc+IZxGRQg1nU9A/4y
1dE/E1XwslvTE1CP/de6Fujdk6isYVAsHwN9pSa5y95/NTnQNtk3cwtse9D4fhBe
KfqkTdc8vpRZIxF8ZhB9Rrxykszkc3I0ooTSiHimjFwFaLx7Z9j63L9XwwZBuGYm
4IhEjd2/a4hlTQMCM57V1VBUp9oHzoGkkTWNk1S3k6IghZyAgCIA5L5WxyBZaw/Q
dFwMBiSZ83fYEIT+W42MsmGxId9umAm2PxGmrok4TnZ131Zeryxf18jIcaMn4V4z
EEWyWD857yhpKeUjjjaPD+k4Nx+/iG9a+xy0zgU1yplwk2Y+4NxRxtVRVKia0VVb
77COeL+GWJd4w6ovz0SEi0ZfSytlFYGPPiFGl0OvZLCf3739QgDamsnvsS0pbiEJ
XpMSTZ1H8jAAynRV2ws9cuOSQ3LaefoDV/UK0BMlivxTgmpDkA7p1wjcvPbwJvHD
PlOcgGCNFo95KZoQZshVst7MPNWSeWJd9lcVyNR1TyYhsdSFeH7QV+0bhBTscgxB
/qbjlB0MC/zCNoFnzrE/fH3Dx7h1/6XirCiXmfA50fjgwR/ZsW4FwcJp9kusK+RH
AV0UZTJ3Wx6wNhCrC+M3ioL7OmxetqN0Ei96x5QKcdAQ1krdi1JwqUShSancGu7k
+u8Zo4nd6xgRJ8djGqJ1RXUqgx+yur1Teyz5YyFU91qEgV3HK8gj5T3xdKy/ZZfw
uxVwUntPvzInZYGh4A34FWx3ok0xBP0rcvtknHfJmuB2WkNQLSCKzD2LOZ7XiqPY
WWjiemprdf0icRCQD2PjmURHIMSAlYgIJ4woRCW3EPViaW2oe1yCbBgqAztFrrQ0
dTDjFAHPUvhWLMGhiOjUCP2UT2lfS+3XXksWSBseQM8o+S/mZSFPnF0uQYvROb/r
jQMP0fWcLxFpaRjGmDe+H2b2B3s7p9pfzfWu/ohVhaR13E+lvL69Rzq61ax+Ijk9
Qpg4ccf9o2WWAdO7jg8ktHZWiHXKPhzP33gy7FOwXJ0ifGu0ygf/5VF+I3DitKc0
z+eVBYcSMqoeF0IIc1JZ5zA/wPQErs8JzBbLmUswlR4ct3pn8WC0Phygde5iJt1G
r620iOgrFJ8DwIm7KkWb7lBlv50V2AmK88jesf/EOliEofysg11LZ6AkKKs3AcyI
QdgrLAoCdGLP0s0SHn00b5zcRiUIKR/Xh+UmjCIhlyz1bA3ZVJwcD4JDohWZvdNG
fYNM6wdJ7m74c8tLWOaXKgIf3+Xq8Wn7ywBhYMeldDJotiqJghW5nL67xjg167iQ
wf93CXfBq5o3TIFVF3XsTpTux1BJSR1BSrw0pfT0FgK8w32oMe91USUtqfKaQpSz
bBaoQ6SacOYzAfleWjEvurAspSFaXek6fERKc6p90gAAlk6yG7KPRt+m1rSR9fiP
KKDXJZDP9lHDyS7j9BCa2RcrySZ0i99Q5EXrT06XrkStpzxJ5yzTpEObdAjG6FW3
Ft6anhaqNNuiqfV9O5KUKDXgzzi4zQORBXo8r6K4RIh7qoRZTEhAwFXAafTPBgqE
w8w8Nn8I4gDUYStdY63/Tp+c7xiI1mGqVaeEGNzuQLV6savAlnzgg1sTNbUWtBvI
0EququlHkz4/tu1gAbvvwMoGZZ7kg2c9VJTDEEPYHET/CsUMIGA5i9kVo0CChXAA
m/i9Wl8AiIBT6cLRQt9STnoz8J8DshZV3FqcHxHJtdDiw7N2RrQ7ItGgvxH7ukGw
7MfTQSGpT7glgNpqGNhGFtBAxEzydK6QzMokZFkfkK+P3ecI0KEN/pyKrtsK/hZu
nyczvORjlLq3vQE1/8TIeVY2D63YsN1vfGkcWYt1tlwOcEhVu6KU9RaNUppSDgnq
5dBv/PRnQ5Sa/E4iNGNcUPWHSiXB6nE6xwrcVwqAfJrU6dEIv6Gmjh6080wTZ14z
s/JRiIjQJ2Ht+1PqRXHM+CaRUS5bV4F5YfTiFEcQVf9SVwzTulk+aErbdBmTbiQX
AnwRsiE7hg5xYocgrBP04FbRBVX8xEXMoQH1FQoIey8Sok488REqkeW6F1g014An
wYZe177M9+9nN3TgQmQjL/4tMzUZSNJTKzH6ThU8X9zsV7m9y2Z3mQIm+WQ3Mg+R
jaor1ysaBmTNlrdveeTy1jvXVEbRnsZ7XUKDYgoVZY6Xsoah4tqJQCHL4scPQIOS
Fra8CCARMUL8fdZj5LB1m+UUh3sJEZlmKEB9Ioi+7vYYt2ee+k/1Mm11o6EUkTNm
yjr5PUSokQo8c+DJ+0GQcL4UJDCu8c7AvMqs2Xa36P+uo+R2YphXfv1IzXmJsXbc
Qotr1A7SAbOfO185orhJKwXgSIY0hExa/QKZ82SD9uyfQdWdVRE2e9/1ryVF2qAy
VlBmYRBmv2l/tZeSYoANC9ON7oCFwIBlsoGSjwWyKPhyNBBvGRn5XzIgHQPAOK0T
tYyq2Vw429rWfrBUdZR9EprsQXd0V/tq0YjpttrG698lmHuQJQ7vpl7K29YAJKoW
HkC5gkOrf6PelK75X7z73PBO9sBnFNCVr3P2CFwAoAOVgH9FRQebKi5P8lN821XS
hmfcnwzxDenbHG2QzKZ6SWtnwetseLT1UpgE7qvzZFifl4ovPHPOIl/Qu/+Rm+MV
lDdBSTmxri+vl7xJbO6rI7yQofMxXsJ8LZT3yQm17vYWS9pmgIZnkv4Pjdm6emcO
ZXHibHPe+zeVNyJFdPDydx7lqP5DnSLT+oEPw2hBbP/C+31yzTU1HcnuXOKBzS9a
b5hRTP3wrUiLHG5Q12WGDWn3KQhUdhvE3sR+ZREpvcrKKtX14mgoKXfNyEG2FVyN
q61A+SZyjAg3yREe6WPWeAHbrp+iN4IIY7nAOXfZquH9+xYiocqc7kBhG0wV0QkN
rogClkcHNNmVZbvHE9jRpblfJotguYUr+tKtFXpW7wJze26w/kuxhgO6nJOioW8H
XKTXqpbPpMsXmz5QYX45Qh0LJwl4wgM51PeSmboJGHDfkuaydhrJCu39M4lpIqH1
6xa9SFXmV0FAiVGxkyW0lz+JWxET3uc/zT4tqJVK4ItHAJPUmOxzOei+oiULiubH
VqeZaJicq9V67HR9CUw1rqMRabKIw5ZZ/EdvSImihnvZo7BBb4ElwXmS1kW6ABTn
b+qeO3RyBWlSm61op/hyl4Pg926qlvhg7jtSGuFcm0+9iEnDY+cNWNvejvG0CI8d
stmAzjxkRM7soksn2MNN5LnPqeI5JKYap3NKPjsFzXWxne/fK5BKHfESRNGwPtmr
QV0pYhJFIHpT+8pdpFK6qD+dQepGsBQ+ay+WmQywtthpST9joMbPP+JdKQyWxRkm
9OqtFDY71FShfhE4LZSgY5CJdHXZuoMvpo1M2IlOAc59cUdJuOByMU+XPclUmKzz
rGXkeObuyE/9EW5Caa5S3XMFjOmd3kXLKxaNxxwxX4Sd+WkOEli8cExJKnpaIiNj
sEhw/IWTwHwk7JrBPEXhw90j0sefENltwmNKe/ufW2InskiGFmrWtCmb8ZXVYgvh
ogP/FrApJ4IheW2Uxkbcz9FHorPpjLwNbktAX82VMmWesJGpb/h17eNkxR5Gdwqm
Zvtbu3EfhK1/2vROpmNTVbeMd88k6fmZE/u64clGhUSky7aX97yT007AM5jSBwjm
XftgLhD/VHK2IAIf3CTVgfwwUk6VvQTABTrAYYo9p1N2wj1KdL9rjdwygey1Wf7K
UeFGgS2kQtLTvKeqES6/5k9iSDe1onSDPR/G9CuzzAnoLJ87Z7/1Rod1Cb13QKxP
uTA8jGy8xS3e/jEn9sC1yMhhw5sMFGL2lNiWL9PT3ThsUF8DBLW3hifv5d9c9uVC
MxTFSrVc2XI6J3Yt4Zez3xOljYuFonlA8UzTKTmhR0c1ammhxQ8DvMoXcL5eUXML
QONdRjMtl6vMLd5MZ6lpIOa2qz35TEKW5sVFcnidlywy+lBFPRd8oJifwKV9BBDe
TxHf+y3jklZ1k0MABQIJtRqP8NAElpyk9D4iadkljCMFUGzCoo0l49Lc+oPnoehX
PSR/CC60Zn4oyDr0N1mbowihtNJIf5BfWRhpK+j4n5r/XsL65+tV3CmvJCyl7DT4
uVPnUJwSxKFpkYcD4LauDbuo+pgMoVceR5wGgByIkjr1AHu08GfWsAqSn8GZo4G5
OQN7cCl+bKPrCIuh+iFcy/gLVRLoWaQLaZ0Snvy4GVRIsR4Nl+RFnnCbWZzKBo2V
0pUeuom1rUj1Kuv/nwg4mtM9cmt9NXL2xkB6/oSFC6c2MgzBnXO7JhKLLomtqoSr
+nMuh+xYwx25SdEUk85YTIgt9UyvsWCmjcQuisrYq+5DSYO4WsRQG2wC1XxuErVV
nj3CyXIgOeWK9fzvXKfair9gKxmbW/HmiGmZr4ojLAYVK0CA8clSbTV+Cfbj5z6d
VS5mUxFRH21KTI00xxwVMs4Jm6Cta8eB3Cu+3WK/lsm5RT6HHexrl3vJoFq4OfYa
0OXvRfqBJaId3FcOTo1G+6L9W/i8LhK2kOZ77k67B+uhMXf6NqHMMJQV9JvSfuLV
0c8YereFyqIhCBzg1lYXfRhSZuTyLEp/Ma/b89IGwm2qj4kWUKkJWv2xSO6KxigG
6bgI64/M/e5yeA5GimyV/iqZ3Et+zSQaLdXwaSTGTvcX9+CzNYdxiICXKlq2a4B6
6AHl9xGE88DL4dt99Bs/azaEnu0PKrHuF+yPHtVWO2s+1ZCAxaQkkIdrIoAEsozD
wyAGrinJj1ampO5dPwlKpXrOXB5TPrINHdOzWLPCIWXROd7vXS22uuFgNSqcd+oL
d6CiCVq+zdTAjOwDZ26Jke81UsijAKT1ikOO2g4KD4CYfg+TGbqtz3pRs5nTfCo4
GSaaxEAkfKZPgsWKJy4aIAdUWfjxXPOAjy5QwyG//+IxnokIIU6WlQoDNkxTAEE/
9BrTYy4ZSdlotvLUPJouq7/m0cIIhlD0a+ar+ksdx3SF4nmKoXRJNDOz4mHoGVEe
+gim3ivknjHSaNM9puzN2RV+6VNGZ0dw4j0lCguDQioHrUtNZep8v6AyRaIHD6C4
xF5jByrbcPabaVkH4uSfwnEQMGClxlCgox7E8AQCrGTekxiaC+JS+Wi/REg9JQ0x
uzlvaMzNYk8tPChOyR9dKVKWcXQ96DbmIUT3qsW0JYPIIOrjZ9Mk9i/L93ZfZWxJ
3DkeP6tirvCDUFZaZmX0g8jgu+4XdzD2RFQSCPqilj8nWOp2XS7LFVnXP/Bwrp0x
o8IrFqtyAaB6Kb3nOlYkT6H8vsd93EHcozZbbrtzX70ZO7Z3m3C53YT7EBM8If5y
7sFpVehHsoSuVw4YpQMw4SzjgfVdd70iQ3LZ/Z/YERUl1gTMbdf+uUs0BzsroGDc
eMotM8uVwZmKJyuw2cE/WbHZTsvl7QV52nsP3ao69GWj6sLUMV0EFAqFmiaozfN/
MstLHemRzBYd6lIgtUnLQaK3qtdoPb82qAbUZqPVoTelXAyyI5eaRimMdZA+JBk8
H52qlVVwYIJzSK7vRedZSE/r9SNRR/hmnLAIbUXX3UEY2Oi2JIrfWyxFRRwIm54n
AOF+Xy9Pb9uovrh6MFOP6z+6+F7lihssoDhSNLsB9ZJHQRmKb0hNya7dnnB6swX5
e6aQ4Lmqe0HaA5B44OZ7Sr/T/mY+H3sDqdv5oIgCvfSAYCKUTQtdq/4vVMBBAy4E
Ln0JGovUMQwezevQlKlFRd02RnhLCylnz82+tKZgGiC18Xug70HA1qGhLUZFtITO
1t+gIidBKuCEXacVqoOL4FzD+BTh3YMN/DgqRntkpP5Kgsfu/grE5bqQmY78Vfpg
x43vL8QVLjLW5T/0uusin6yuafK3TV3LtyWvVNG66caAhZFphDnCX57iJy8kzqd6
u3OtBfa4fhdm0wJ5WBRAYIbVWRVkmgqMmkxRxks5bHy09a+8299heWJok+Adj6zP
CFMUg9RaWasp3+86CsWeHgwZyYqsvCfs3xazv7Y8c2W+6E0cfm9M84ezkKM42eFP
ATtJW8BRHN3BDFrzYOd06KqD5nzDIN2LfDgGm76a4QpFovZg30Cz6EOKnZhiBl3x
0e6sbayI2N6iHWfjm95t8ivvhfIgIJ6I2vF4jwWtck8XwD8leTgGoUgUKD7KQHDD
BMAVoaf1KjecqsgrY+12XV6V+rC7MQynKt08QUL2O0aqTaDY0cvD+ZT/7no4joqv
8chrJfJIBwm4eaF9gKWssHMLwdh2znvcuHesPyFFxWVbIXbqEWlByAGvfRdXkn19
n8Oo4I9GpvO9NpKuRxJtjHEHgCku2dGwFl2xakcLy69zK4q+TChl1r0fk7oJguOi
KMV6bPInWSaRl20A7x+0Q2Nh/xsqzR8OHd3msP7rLOOpf5rlNzv0gBYItXG4zzPr
Vq46fCdpE6cBjONbFdZg/X6UqvUauVG/DK+S6ig5et21lNiiNnJgk0pUiaoNqMNs
CF2s+UnFfWZXSlgPmiQPh1MaEEmffb3ehqfIUF4P0GTD3/rd8G6C/H5L6hCbXLz/
TSC1gTNDvxSzO85sh6LEe21ThVcC4iOEIk2YeaAsYI3r0mnRHUYAH++UZ1qWB7Ma
y2wYOnNjVsr2znevfPQQOY48lODboRM4SNBC7BxmFLZLAHFxcP+lhrpZBeijGmws
6bndZ3D3Y7xyiStDQK1ZzaveUr4rS6gfJsrD2NPbddcCugqqM6zUO6RqqsutrKny
U49arREjyrBGHQfrtX0j+xhvjaLYr0AP9wWHvth+3ZlJns74HyuvEyTlEGarhbJE
8Zm3Ky8/+yVf/PqL3KhF+soWnbpcObgc70kcEdSgluylBuGj0pIwuOuohabNtYEp
QDJOXo4G9SmHvmTw+5At47ocFe6aKou+ySB+o19OtUAUCfoof71gEOaqreRVPhn9
cWczjVIwWDbhmD2AzGJT0Qs2Jlw8vgd78nXn0hu0sy9LmDXgIr/ZooKwdGTBLdLw
ZJskw7DQPW2Xj+tM+Sv50V4VIP6RKXjtcjITH4GSwaNa3iswHYcA0Wa8pNAd9EmR
oJKPHmvDLpDljlE/s+HJsLyf/L9F8aEC0JmDryMByb8K4tZJbDux59LNbXvwreQ8
1RjtPELty6nJ2T24paDNqOQFoQwVBX1uHggqre0itx/hEeEj9b9BEZptSRO13xYF
QOg38TP770VWJEX71uaWcV1tNkdlrKOT10F3fgaZyDmZsjSjVbuAwEspbvwT8LaM
mnG9lD4g7SAfdQiJMX3XhbnvMFXraTDZccRLZHKMISzle25xMZgIp5LHLLs0ZMhZ
XFGRcfRw+OnOrYBbM+GK7Qg6y+6YyU+zkoZdp1H9+MvNeEle3xcFX5oM43wo67Sp
R5otYvWB38CqCT5IngUC/X4bRhQNpZMChBgpmq/Ou2VWk+FubJQWOP3fDAgUQpSy
zMNYIa+UULiexiI3d+SNQIi3K7zr5Y9XATD3NVfRIZIu6A+XoquZz1zcZf4PNOwo
slqi7Uavd9zadWiGrqjU1PSajaRa443CJAKj1WUtJz9dOnTdocD8IBYeQXYrnMf0
FQkoFuQLGBwBFfISiEAN0+3ODxHT45Y3YgRysue3ivU3VQ5eLa8rsE157HewSIoX
HWPTRrQZEmYN4mnL7tPeMi4+edzKFhbbv5zHG/u3n3kIkItOy0suqb7etK8R2hck
MfDn9l5Yd7usey2y7747WCmI/n3eX5Dm2cc52tNgDCHCgEHd3zsk4DYRGc8mYOf4
F4eZqdDE/i3anU4Jsk58WMi791f/TPBWYXRyxmo/+v/Y2WNr1cpOG3xXKDi7k9MA
YOOl6t0mAFE8pUHbEw/zTgprHd3Ot4VOcOpRjVAFVdIrlZWlXhgtVLA5sKjZvnvh
VxE3pT2AYOuQILYYQEpqYg8P+bx1/NlLOcU+CXwL7Ax1Kjj8t0nFYRdhXnZaYkEx
X842zTK6jfTNeHLOaypNpK2kJ+wiIQ1F76ANixqOuT2Vy8hPlCOtsdJBOxWw7tOD
ve0r0hVBbPujhYRY6b9AQvVY2SW7Ucuvo9MrgTJyjolyzEe3VT/AVe6mm1+JCgdC
tD3Hd3GDwf7qLfhi6ip9TuzHtUg0dSbR4O19fphn4vgbKAK9M7wCzluF/2ub0Rf3
ZHnJJHUysNZsdyHLseNNmnVjzkA5r6HqEOcv9OuIw168HE7bF0f4JSmWwnLhm00c
fGfm4AgOB5ECF9AOmMlLsh0aBkfVHDHnmmTfREafw95wvt+xT/vGIrlw6sfsLCq8
jJxSIRfz3X7a0zxtRrQuefhDH6vVVyeSmSTrZ7alEGgkYg1khwJnWjzaNMFVacT5
qjfilEotk7jzdCCboz1jY6fLSUaPBvdGOZ4VtjvYKB1uX/3RzfJ/o8X/bFDEAb7l
hjUNoaEISyYqiUnm92GZ7QvZl05IEISPfvxTCsifEcco+atPAtbU4Rim+tSCJmOY
qvURbbqTGj6cfAJ4Snr58ks7ODHAU/AHM3Gpo4YNg+rbTr3OxeEoGFwCVkCIgqfT
L8K54M2wzrI5kexGJrFceLOwXt90XZY3Y/gUfrghiyX3jJAnV+SgOTK9D8f23VAC
BdsKAGGO4MUcpTNsdYLltRsQtnSMtoxlLIx7uJvGyOeV3tMW5yaUMFp/MiSDA7/t
Nl7kEAdeGe3CkmL5O7yjEfiEoqwuyURsIfcimxShqIYo2epG6TlhRckS2gtVK82O
fy9pkYYVV52m5wFoC9OD9YRBSSwum5vtnhhSq+7cHwvz+rgU7iRNnPlM7WH6Ecml
bEUMIBfSpTYELntg1hrwLT4G4vW61yS6jlyqs7K0a4GhDwqs+J9GUVERV6iOAed6
Z2XW+MaNoHDKTDzBHF8kRPbxPnce06BlbnJ9XGKLAn3joP5huhevKU3RsTi9U+Ab
2d0zvT9EVA+WK/fPR5TN4Xu1uTTShNHsOI2PYwxDTbNIb9se1PqXUMfQiGDbyJvk
JEG4lBqEn32isMqUrs9guFvByeZvR43o8u6VBTRYH5/tQxxI6x3m8huxiuckuSx8
u02Jv8tkkUEEmyKOLS06TiI4JRMxJeezK+DOlmoS69HUjRTR+AEyRRAQxAtQXLpp
rEknOnCHWEC6xXxXfkE5cgySZWAUu6EDHX9N6jCuZ7AlmVGMtrTu9inyBPhZeROT
s5ZDRXIKzUw0shTlfH9nonm/dNwxLn5jg0LdN07gqgHNhwZrB6GuqLX1dSLl61U3
AZQjMY3yJKtdBZBZfo6/b269TJ6qzVxQKu+UspSLMWXOw1zCRBfwkrSxVEyZmJ4p
JtZawGrAqXakAxJ6jQc7rDwwLcgq1mrKuf2fZA2oFpDLrVy4CiwQ/Sy2Z8c8dncC
RiqFkbbimqjx9vuHXGm3ibU7VdzlyHRT/tjrQuXXpBPbsti0PFvaszoHABBolkpW
KGu12ZxEY+xMmFoPSKKmCFkvcD0GHjhWiGc6Qyh6KJNqO/vJ/0P0g44Yvk6JEika
sQRQj/f2W7jOn1BGC+5aK4xTNO99NGUiY735R/u6Fv77FT07BYmMECdTVDUM+Ypu
zQLkEmAzhXrhVCZu/Bp9WAkFlsHGhA07YVUQAHXnOjFxTfmm+43TEUABiD3h51Yz
Wqft9LSuU1qySS51CHjKRPnsfEp6sh7U1ZBSYP4/JSzXy+2k+jDKJnvwisqg6yUW
VIe2+5DSVuyo/RfPN3J9mOV/LsZg2nGUTYMF+kqvy3IY7jGJByJwST5BYwCidSO1
it6R2ggCP2OCIh+m13LiaJvqIr7ncQT+LpfxA9saGPWvG7FcYJRHm1YHoqIvZQa4
HOQlB84330wuA6+lJtYDLkE6cIsIJXq5wgJXEutqiQaAoExj00KyQ9jw1yM3WwF1
IYwn7BQEdRczRmiMAZsTQkQYdVde2CKZohCVUO/aQaqw2LVGDBRx7pP6xwj5TSd/
kcGmnElUj67/mfx4taLqFA10w6YIW0Rg7CInDeOqcdHyRLsbRjRxyLjAFzKjBWoz
/gfF/ta92yjWBoAzxODpW4h7I1Z2z2bi4W9QbIkmIAIuyZNqbY2wvM/ibAF1UB1f
eqe/+sTYnGGqD2sK4PE7WLpNpR0/5GtxTEX2OJmzQEQYx6ztHC0ktcGVO8fSs09h
QpjpF+mdKLCboeSeoVWMBWNFsevFKRoaOPsn5Lg2H2WzrzhAJv+rMuWgKL0Yp/Db
ZEDCBn8ZAVcZsdeTsGoNUPzLicyjZ/Gpwcl5fvcWLjwi05QEhP+2pBupDmcR6CvJ
MinnaMSP17qq3QDKVCkkzxcyGQc3c5lrr9xZ/YlFMpgKggTX0tJ1qF3fZa/3CRuS
VEWq8qdlWRp8nEpdGdCa4uJ/Nu0vNmgRV0ut20sNN/kohv80HY6bpYE51+ZaCyg8
7zJp3No6iQnCLVHqqpn724l+fKZW4cCvblKy/OCEr8XfnFvMBK5miXL0crOgGXPc
p8PHyadWxDWDZuUZfDQmrdH7rsTW8sOE2HR8GPpAJszZ/zAPAmBSMMQgQq4MLcpI
TBlrl9U3HumRqa6jzIvV2ywtiF1TkYitoRb2ZOIpO/2uIn+Zsj4JzrrYdqRRD8ia
9FGUR2S9HPgBsTpj3gcjqPl+kbByuZzacxxMctfxzyihcxbMMtnbIvJsWC2Nnxcc
POuNyGUmhfJOzy73d5AjvbxIunz93MguiKMQHJPxiX2WfkylxrZpyn79ylEE/81V
hI+lV/IuXYJDi2g6no+mpQ0JRm0OWt/JReIOA2nqoOXTqDChZ9yY/fo23xHLsAtZ
H/lyQcATcKbZ6G8HBquoWky4LZRBVu2PJ/7n/jbz/v8BMm5yXN7m5pJHs2J7A+7m
+iVJgy0JSTsJ628EP/dRQClwg13D7GkTdpTQlslGKf66HtImYLlmnbq40DowqLKB
w3bPL6CapivA609uezDkQu8sj1eaWxyZe8veGRMy0tpmEMQ3rj0nBbdVmhdUlyuv
Tm0PticYeGTJdy5gUCabxelyWs9PlySd+Fk5173hR9SRLrYxSwtyr+Tmnw1ACXaf
mTUvsqB/ne5ZBFcMWJVdjN1L+equaFk0Vv3co1o7I8jvusBGqFH+XllzBo7hpYSp
NVOSJhydbMNYfoIWa4LdZWbw8mxKG1TY1orysFE2DcM/QpShz6yHStlT7PNIM3xR
nllVorUXg2vGyzK9Ix4HN+GTd1QdWZXw/rhvGzvuxnQlN2WQuQuZOCCpJFPuNdeA
c4yMheMTRRKsDLR4chUg4o53qrTlkZfpamLVvAUX1hqjRjQi8A328ItnCZtZIIkP
g19WAAqxG8XpH4eCk4LvD0UvpJ7c+bo3VGEP7ZIafUEhyzs/CLtvdzklyBY/nwPt
MEjURFImJox/SOlyLLDwRUAX3fY5oWxJjvaddoetVdsy72s3zELATbh2CxSEhQRs
TiS1oV0DDJlCw7kiKDDo74ujXAeg6EgiJfaDiW/84ftZ8JqbBcKDkFMN0xmpArz5
Xn6KSfFnVxlptt+g/vLxjYlg4ZjTV+Mh5s/LvWUTkoNHmfyAQnZs8Z0QHZVn0cWC
OBG1ekfOP269XWq/AcJ7COK+xahLmNQU2lVmFDL8Q+PmjDDhkdUMwqiJDPGmpOhN
8YfCMvUtdimClBuaaleFJrG1eYYGZxSMQzS4YFCcGl+U/75xuTVV9wL9mTo5axV9
bRmdqOXptHN0uQ1jct/IyV6vpULglqIwiUWfkf9lopS4EN+HqH0fM7n4fL5PKNEZ
gNcqxk5kgGl1bK8a1IlvdEFlJyw+pfeXfE+bEtxd/dOO8x3RB7escOTeyb/Bn+Er
9KeHU1r1Rivmf3M4x3t3WcxxljbMGlflVRZoMYV/PFok+TSV5/+8ofU1YyJJB+Ao
MorvWiegrcpokS8KcfeOg9VHIpL43EMHqAiDznSCy6Y/bSl3b4dWjX2SHFnPra3w
gjS4OTx8G2fFkwwObRCfYkZQN7SJCcAyZWnvl58m6J9BP3I9ch8TlaXKc46qYOxd
wcPF+WjTLsSXNtMOUA5wexNnNWwlrucxc+qQhEQrYxYNbd0eAMSICzXBL8AgSvKI
wqEZjeHsyiD9sDAOMxHzqCMYKQ/bOtLzPyDtew/EhRWTZb4kLYEKLFTCFKYxe2uU
IqMid+6rwNZhlWRY16YhDJbLY4lzpjO1/Zn7+h89lyQk36f8CHrRClMRCaZ6ju2j
mHRv42GQ9scGR3/fXDDWKQn+VCL0WGmWdKvsEbmHtCIJovxKoQdf3I0i6gLjHW6T
MRfpbWYJUml3Q5Jl8lCW5z4fl0j2wIrntZb1wM4w/vRf0VUb80xhgpVWlE25INbb
lIXJxN5nZ1z8ihXk3OwkTC4qD8i4cYMlsABKTnBFwRrP0UAPG02XiNYGluWapvTe
y1TEjX0N7ErKdhZOYxL58xjH5p1YR8flu2vsRSXarsz98qWahTXwShPyWlot/UZ7
29ccF3HOD32tciCPx+8IKOA6Y+ohJLz4kSxgtldRPtWX4ndo2v7WMpbazlD4W/VZ
0TC8Y7BQ66nvw15JwVYqEhSzc9v5PlOq/cgpwbtQWCtRLimHv/rcnJQs4iZPLz5B
oAqNdcf3LnvyuVv4G13O+ZOLPd3SbA3VN6BRwQMAfN88jJaKmhfnVBobwgTgqtPb
Yiae4lhcPNkYboPjxoBJYXtN05Q5PN+SjUiU2O1XWCBGoiSCLFFyyvQTkl9XKmq3
Uw3WxrvLld7w9W0A/DGXd7N/oMdETw+9sH/SqbDzaf49qyZ0lgjZfVxwuozyFrkX
PREWvj4gFPxdQ9cPdFUfeXSOC8l4AvP/roQfUaeU++exbMiDWHMott20d9wzO3Ch
ybVzX3TjPboUTA8FqOWjTiKZHhj4OsMMpM7npRv78ltsmjxK/nGXaiLXARv4VweD
RRe6TieyP1FgYFYiXyY+m3y2ZT/2mn8eNmt9ufQ49Fw90MUQTmyVRw4d19tZJI7x
whXQJOb2ygbXMB/rGrykOGjgusYEAhwl1uqv2SvKyd+0kMJCZaVVQ5/Pr1LoxLJQ
VeOu338r5LDjZ05HdZanV29jcUqw2yFZH+jPyBTZFFDul1gAHGgKz2VVEKE10FYS
qzOEjPAmMnXoUw9n9nkS1525qDaMNNk0in4LJTcY1LHKXekcuZP843um/UooACs5
iX67fq6v1XtYzJZIfPl9+aAAhK1696H+rpZ2mBw+UJ4Hxv5aXgsK1pETwQpeTolM
lxT2UgmMoQL0Wt66PrNo+l/5ZfQX+hJ/3GC4aDBAhTFb0vHgDoO6XBGDdgvO2xB+
QbzeRyKTX2tJNFJoe1FQMnJO0dJmoDRmWbknmMhzHcj/4kcLvmVgLIsc4UEa2hbZ
Jitn84sXRpn0vAoKhRUV5nRYRdtuw8kVrEKVfeqPPCU3qbMbMNCmR24eujXeXJXl
45a8uOP5SqbcBJ1/hMW4mxS4p+a6h5mcbqrPE4b+AHsxT3p0kPjmz5ktcOiy9AzL
Ud5ODw0Z69pXu3b+RxKRBWlCCKCbYCOdHTmwAHevNMH2mX7kuaSM59kEQ6gcAu1x
kSQGMcSTMCjhUWvOBpt85CLMy636SFkkYtwn4+YmDsLVcy8pte4dJPZuAvDtBZcI
sqD7bDaWJFTsI9NHjtlcL0Wm3Mf75McO/+jaRH26+0I6hSbn6naRKGD784DhWzHb
WFHa/wb69bJehKd14tJIP3Kb85Gm26ay2gdUWzoQiaqaEg1FYnKmdIrAcg2hXibf
wPOOSNnDlUbXM17QuXzMw2gHce9F0t0VRWSufzn+cSkErtWv6fGk68h2PqrA4iIi
/eHqxT9xSg+G8zMKvApOJSBdlVIqzKkT2RBrs9QpbZtjYXK9iX9DSdZE4U9lyv3l
2AdoLynjqs3mrKNCr/uv2we4J24SuyqFJjjrP5VCu1rjClxeTHMa6DXPMX3usxZJ
U/hEdnmNyIrKnZdxn4IhUeDwIdNML54hyaX80ZH+fyc9wjmcorqUfz2bbUapX+Ob
JCMl7INuMglGFS0pwr91DnGFwZq7pfXk2qCMfU62fS6uiUPH+rc5A0NI2/G4OOi6
FE+CWTqiE6rAlpGWnypCCnPWjcxcSh/nLFgpeP4fZQTPoONt7eY+48O7ffa+Lgwc
Cp8gO5SlEJ2xdmi0LaGlGwD/z+aEjw7pbuE9tWqeF1UZbCszuzTX0FiQES+gUHyW
IFS9GojHxXgnZFxMQyS21CBq1pYDRm2l9lbxgMqqyAqdD5h6UBNOYxaGEGSmHOMI
/LH2wDOlIN3wy20cWz65UYXOR1pxezqHxuM4S8MSik4DLVp7gva5JoBIHLhZbjBP
boR0/q34JWnPr/yD/BliRd4dxUMCHINJMebMzbwOed3TO8+nAvsdpXxTPsjW6BSD
l8GfRGg7BWnT3aWincpxGKVYX3PrmuAaJ2rlnAObnQB4JkmAUMsDgQffTop+Ymw6
u+U9ped/8e/Zy4231MrHlR17pzj2zwMZccwli2ITHy0js35dAY7TTp7m4n1YxJMT
RiMkrgBMn0KXxgRZxxGg4mMg8RosB1G4PaH+IePKV52MgvCMhMw8mYejHY22tVqw
3LN6sxanhoBtNAwBYMMxMzB4uJ9L/Jlr2+syBMArdc5THuOMxTeFFFvWkSkvm5WV
pFeMsy6GVpEzJ9up1PuYPT57pu6qnRaRdkrtmZRjIKZz6pofxpUq+fFy1WE0xaza
jAA1s1oVOtcgCoYqzk5Sse9xzAJiOOSqPJXOUZF+w54fL5qp352+BpMa/qE7QaWq
94MlU7UoyYWYVrsO+YWJ/rFyRKi1Ujk//4MZUZZyvz1v3eNI3JtrR8gqDJzkTrN6
YJIuT+xd6ymGjdoIZzLYSJB6ARa+uF+U1ZPTvn9rfIDDlTWrjxhqnSIyd6FjEnA4
ICISp2/QXylYrQ/GocG5fyzIt6AC4ic31oPtbX9IpTEhy0d0t82Vm1sVGuIu0Og6
nco47bsEzmJ99PmB5y47vqnzGdmZBCqcrKWGV48k0/6ywpWAdLLLtraDRMLFYovd
RrbWpvrAh3zbGPzXDPjVypUabO6lUJeJDfgw0o9qlyB0UzYZLoaAL0YOx229ZlyF
0p3tcR1vnw7Ye2nCE09unakFFMiC/dDH5tX4JJWgJpy1pf3rzuLoJ7HaOp1ebkmG
X7EB//lTiyuK1GGTvFkbNIc1pzPJG3FkQ/u5JXpIBPNH4CTdQlb1t8xSXpZWEM8A
xKT274nNwBzJ8Nq9YyFYL8pUVpL8dFjkvoCJphcUumsFOmlUPafk0lPn2Bm1h6gj
0hKk75/5sb9lLN3M1A8LbtYHiKDn1SUwe9oTERkEps6tovvoTKze8ueFd/1LJQ7u
AqxrWhLZY7PyW+OUSXmGjcYyS2bEko6ysnIzsZAt7r0TciaocYC2g4DyGXd6OUGo
vBHy9U2FaUPiv5XsssMNkafjv294lijocI2PvgnAPWe+Y3qWIFOzE1l8avvERGtW
5wqplJrJEZeNdCgCKVOkVM3lpcADlBEJVLwXXTsqsc5fbWsY6/VmxjxkVrFD9wlz
bsymBKZvmKRO/ibAaobK0mWhbRtoZ+Fd+yqj+EitEM1GA4KHkU44ivcKgA3oQSZS
/sSx/HVh8sVU4CWUD0N5VIrknF+9mPJzSN1IGNCVGlYHlBTM0iElF4L0JhD6fm4/
n7+SrPswiQY0Q53dT1uj8l+7FcQvWlleByngvLsRXnZ8fvT+J/IX6IYxASuizIXn
3FNBWBk05EHIpreOC2wbjsN0Sn0jUo3rAbvgqvGuFNBbwrYzawXMwKCCx0qKuD4U
NH60y1ric2Ivxd0fWoWJDw2lcSVqBA6lCn2YiT0Q0GRG2OUFb2yF8NcFZ4USy23S
z91Rfl7d/ipokYRU++pfCpN6cUcxWoGAck9F4wqx1TlmXLWO5yNVXqiu/ctTl7bI
mtlsKqWjBza4hAQDbAxDwcIEsL/CvJpTYNWrrrr+Tx5s4GhjKaOiPsujH2dMUanj
0dd2J1JqldEO9mPv9ONZcxNqMURW+W7SpmlUxgWPaVandtJhnj8dW1OaoNep6YvJ
0LPuErWNnlzgFvADWvAGfRc0EsGCV1rRbIihb6qDmRzUwuclI+tS+fJRzMMH5/9e
vBfxROReAgCEB4Y4hvOVpIWNPPCIWfClmrXeAf4sF6Cy97VY3PzJYaYXC1TGXDGA
COknBR/izVRJtxACT5MJ+XwKLiLTRmRZjJA4TzOQdCbQWX6LPJjuzOJIZBOQEpMX
W3Tqw61Xcd9Sg0NJsa3SzKHWuJDJWJUbgnJ9SLAkzRoY0LJlXNDJ89VLRH1y3/z8
xCDmF4GNyiOLSMc8oLDv1R/1CqLyNLCAsrzKXqDTkw+HLOrmE7yBsGk6flxdvl6T
Ka+5Q4DeG9u1Bd13J/yC0Dtk7YyFlsbbOrUWqd5sgS1jGPd/Egq7N1kAJBMdVoXh
+Gn9qiOnZQCiqiqJvZFcFt3SgcnCqAm1cIebnNx1vrxS/6Q/XA/waGLe2+ob6vGE
cMQ13ajQOoAwN5iSpz+GnL7G2SvhDoGZV8zFumb2puZiO8Zd9Vrb9VGpTYd/IeSR
ox5DffEIr6TdZx8+4yV/w10guYvsw2VO0kseFk0Mz9eAGUOx9qJ6+/W1uC1N9DOS
A5Dt1H3ge1+gEFvZ4GA6l/JJe1VA5nk31MTHDlRiiaVI5ZbIWTUZGaVmboqxzZIf
0C6W4fErMWO7pnQv8YJC5RiZSVJxLlsbmE36IYLV2GAMDOYBhhJQgHEBEw3U0ygE
Hha3ByMo7nXdlg8pW6sBLmu0vR8H6cF0I9Kelk9jaLp+smF6ZRQ1e87f81mRIc//
B6/joRL0CcmK+PvOOQXlUdtoaksss9NsuJBe1sMbKlOLvRyYtb8ok6GUMpec5dRl
JFWBoKuJMF8RvR0W9/uMO5HIHtdOPblNRrEVPc5l25XEMwcG1pFZGoGCYxu9vHmM
+gdVHn/992FA0T2WqdYBm1rkc5RBAn85d9nAea+lXbiH3m/9RVVYUnUinakxOF8w
UwMsjo0HUKuG1A/MD6c8EocqxLXxb4cBfdaSMt6RYNO0xJD5V82yCsIwNLANBshH
t0NVL/WGY7BmugRMk0NertEYIw2cHLf03ctodFxpYOxA14/Y4SJMmSLMeIw73hJ1
oEwmMnXYKl1XndUzzVONzqNUKgGwXvMdOeZfou8xrhVhSPk6Rmz47xBMbj7aPzAd
HHlV5WZoY8x86ahAhn98oq0JGYGN05lY0qD7N0RZ67Ru51Ri+5agQ3lDVUfB6k2x
TSQuJ2XnIs75Y2ZOq+VXtjHAZ7YV46DDWeu7ozYmhZr4iA9oJPsWVg5Q3fgxRZ5o
fCUVc6KmrN4r6cX+x1hHj5U0FxRRZG+QaJVuqaL1idRHQP2wYYs33IJRkmr2KHFV
glsV6IQSzn7u7dEcNSLGVo27zrh5tEK6rZCAP93rTfvnuGKvZLK+cIPk6BQXrVg9
4ch6nL/RpLvw+9uQAxyje9dVrr59iN6P6hf9dFXMwh9cxOoWjLh6e4qgjGdtDtIr
1W+uS48N+YvIcI4HQOtHSA3sBUogKrgVorsQwcAKw+HsPqMp1Dx6MPIg3vUw1QwD
gMrEnaQQvfR0ZSIBFzCZp1i+0rzMZLPJQklsLesS5wa8bx9it1jCYC1BUQfqNPQt
EMOIOHmCVLa+6bABcl49E/71BKxBuzGeZyhGgnQ7Y9qCrWnmawQJg9kCTAHqDSVi
/bCPP/l18IozPwaXJiyOE67cLfTkkndSYh/vlYmonmwbDqVW90Ak+MXv8+FpqKuv
3AGPTQRZt27G+wlcSM7tyK/ygba28+sCNMIy3n1EjN5hZJCgSyioX2TOx+S2sex3
OVcsVSEAK1trACaqDsQs/y/Ddv7wzXzc713GO9BuFyU5QUvDGPdwWGrl/i551r8i
VXLT9x1gMCpjpQqfRhDZtDSp5muwnts4ogEWYbCJdJBKHkMiI4+cz2OfcryXOXhc
YRhzPC2L2nHBsWMeY6foDC2ODGZPwcC5/au2FbeXFSZGeQEi/wwe+7wISqMWfBz4
8ojfOYZgpMdeYC1Sqb6Cfj+tEphFxkBZ1vgem2UP+XXy6EbofxcTTNyw452G9qOM
ZPVM6pC01ADfAz3c431miw+PFHStm4kHZxziYyURTaP2OpQUHOhWhDJmBpdkzp5j
lDHpEU0Kc3DkTaXAW+wy/zQ1JJBja/idsT5dH5UoFrPh8IqReqARYA7krRS/gJ3a
Hw81H564FrdoNyAHmD+E+l+riOKq6bUshdVY4QCXcUclg07HNtHE+6ZDCQ6brzRs
13KsG1V3xZXvSdufLTheC1NwE3b90Ufxg0xDSVswALDRlSW1m9dlaocFgaoojoAL
3M85v5x70DqxfUBYNc2EI11FPWC72nD2Aj+eVqTaduHSVFVs2mENtULGTwshyVER
2+rLkuFJVs8litFSrT6UQpNi8DRXlbTDhP6Ozx13K6r4yhQEvSWIIzGDEUguDRSm
qrQAgtuohM9+VNCkGdj+2l/DXoiq9Ty6JwGe9q2r0/jCPlHdBlNIqLDi3u5g9EQ2
+P7iqPhqPhylTL2CgFOEBb+T69parZ0Wgl8uVmRaadql9HzmbO3vQAJNIs8VZi3M
zKuqvaQOCW78URMrtntj+fDSfUTxEjjWBMdM26EAa/kqB7nltSuX4tsHb1xVJWAg
XOPjXRoWvtsWVpWXwnKEsl45u1QWIkiH3myPuPpSoUlRLTRYAa4l1FV0dwz2t5DF
HV2Lb4vuJeW0qS295NVwoB2C9Q/P7KLPhl91X42fc+8DhjwQWoDkjk6zDSgIwAbc
SQwhCw5iEdVZgaAMF82xVEZs3xNU9gh/HW7sivtYPsiqeCMd9LY4s2sjxMFRTFUj
Yl5ECHGBXrFJZHpU3X9SlxSe/Qkikbi4vsxvLKjFna6GzaRifvEfQLe+qYmr+nT8
snCQS8citkbif/UaVDbs+3wyTSw/zfk7icVYb/p8mJGrGMUPNmYHIJc0tXueu3yv
iRulA6s4WHDOMkgA1gmG3cX+zcDjfRA0etfjIcjq9yvCn4XtGvRvYnYhW6Ps3003
5APrUisRfk/A4BXwUMb+sVS/7AsTJHaTp4inB8uMvK8iYcaOnaYLUvVLMhksYK3i
7NKQv8ul0QmxjfcL2KpfQa5W+YkiGH+BpSMX2rHA1n2SYE1OjViSyky6TTrXHtEK
UDcXKYqCxgSFKPUNA4y3kVZsb5Pydar1Tl+tc3pv4Iz6xN4yHy52xSNXmawIwFtA
nYxM48iQ1JOmaDKIR1caay4EOf3jsDU1tSvLkEyo7A7ZQ9aQ8gAo1odJ6e0FajF+
7UHVyVIWhpKUcPbU4fWKCOJTdRwF8j1BFu9WM3vgtgme4FQxvvk1Oxey9B1OcD8u
YhlBxgL799XE2Bf2CjqScsj2DpeXomEcFr7Q01GZxSQsbgZ66pr4AQuogPeSlj8K
PoThcfASpbJ855UPgOWa/qinRyy3VDXntjU/0Lw0aENGXNiTR27O7dEI8RzIYnqu
T4b0NbQgoKo13sXyTAWCiBhLItr50CzimrSbb713RNbAyjyN7Smi51T6yDNzyWWL
STpJUrojG8ybk1JTlOEoq0F5D0abvfAa1K3AUxe7JR2D1Tpnp2skisL3xutqiLOs
05Imxe2wGt1si1Y4oFq2owQ8e4iq/le+rNU3fYfHJrU53gPV0RsxrT+QqKO0pJff
KnLsgzPr/clZcFqZeCWYbyWFILQMUUrLejE8dipUEHIqm2sY2wZD2ys6KIkI3tYF
reogMBwyq08eV7/20+zXw6YO8DUiLnt5l9PozwESKqpw+AD/GD4EZq8fknvRknLl
AWiYLSLAwe9xOOS09HWHPGRvz07kQEdrZPBH6eCxAOYIM2hKX3jRoWBuNFDCVRbk
8hs9LSz7+P59aWkapAwBdQ9Dfzfab3vkLGB7LLvpttv0OH8FFbPjCWFlPTYSrSg4
9pdVptM+GNOjadDApzoIJOHbhMbN9uGj90p/4Ye6Cs7CD4nQF6FA7OE+AX4zTbxF
/jnATUmm0EIaC1h+XGlFDticpR+4qQOHsmZffFNM+DBzznDXHW3spleTsr2jL4nJ
B95aTPn2rNnbnaSLVEkY1BUcdKWaoUUHU+J90d5p21PfgSx4cqnjVvTkW9cO78Qz
ReDIgkymR6c7GjjZIebTUap/3WpypfCgom/Ms6RZd6vQGpqnB8TC6s5vKeXs5hxW
EnBM62Y8JeOX80nGmshSkcsKzSetrHNqq5vlypOlV2oa4bcd79T4ZWv5NBNKruAI
Vb+WYIS6KU61ny2KwBo5dWXwuYgjWPk6aRa4idUBheAiUOpO+0isSc54sYE+fonB
vq1U+3mvwmiPu4xSu2A2lE2FGMiIjnuMZtj0Lvz90/Ih69IIfGn+9iXRT+/iaiYu
hnYAqMpOGtnvZyvwbgEyToxayz8/FgZ2PBfjqAm0Ua2b23ucpGQG1NSkuZDYaR31
a13dqTo1R2Ji8LQ8RaReHXo4e4ngyMqsYIBOGX4TWrIGm0yIu8erhlXs1lDSilsc
Qoj+SpKI2bBOEZo8pBJ5H5c3QRzO6mqaE+FNK7cMS9otiwDwPqttqlYesICBb0hL
J9RxDuzMX9c4Jig8cdroWA9w7L2zRQje9VGIvNlCLoNF6E65cEtNpr2UMdyJ8mGI
RCPnBQ6pd6JXeOeRAd0gyq51zje6fb1NZWcY1y+TU7SnnRVli+wRA5SIxRdEDzFn
EpDzJJMLJmSN3ciSWFj49ELEDlckrWNvpfc6O9zdc8sCDpe1YvnNwie5EsQNJMi5
ZWIQrygWfZi4Ckd8hR6lpR+ynkVg1YN32TVOE6u2a+QMPca1IWPtpcKPqixFs1dq
LRlD9xOhahbNC5k6gQKoTGom9BuacAJUw3DXvxFeilKjDyHky6MZasjIHo1MiQ+I
joRqQON6cscpJkJh1HG9o09hgXv51vAcvHvN3HWcz5pD4uagGfvVfAMWpNdq/i4c
x28fWtzM62/lHavd+3LRAq/KS0hP5wku7tHphQjnBGGm8Fxvrj3JU3/J0hG9Pwhn
lH5tCpR4wrX1VvpGsuc0jaC9eHDNWu23qApORekFjEDbigfpIHEmWYgc8Pi1hRNF
jOc68gtmAr/5MfpbmgCKueuGpCR34V3CVMYdDTww0ijNEehgWJtwoKKUCirLALW7
2Pz+AgOcxJ+Paq0NS28n7KWewoFK4qD9RyIVtJ/wKP99AAdufCICgau17DAiLYCX
HEUr865r4f+6xOtuaml6hT2VnO9k61tVRYrkU9LcG73+s0qDMGcOBZ4Or48Hhyo+
wZ/htXKtNjDoOgN10uuEjY2JlqBk01UXkmr4ffDNSeqgtOF0+DQl9dSa+vFh3z6Q
zrpdUOd9zhvOKpFEsLCe1US5up3P3TJVl7qlAWnHc8OGFFmrQhG1i0MpiyzATdwA
B5Lm3ifRRTJyhQIf/VLytVYFK4hOpPJRMyG3IqZaQD2ywGp1xq1zsh5qOjNeO4mY
EqYqzGy7uoI9nIzE4/JQkSniIZb8gBz27O+AWqkv0NSlD5SmflVdlFAJ5cH2Jmwe
kcKjYKZ5QCIUlZ43w97YzGE5+yypDlmcRvpBYTRLgWbJx5WGGTclZSNQN/SGZgTx
hCxxISfejd77ZlHnWuV1rq1t0ErsKPs89gro5TT4qT84bFpdBrYNIy9XfgigD8X3
CX5AKsc1KyHa+U2czM83Ge8UyMqz9XZznzT4xP8VYAjur9yAzcfWVpVW3H7qdE1/
pHNcx/qMRglCAcB3yTvxMspy/a8TbIfi9zXKdbweqX5AYPgVsLRUTmwUcKs91qhZ
vt3omtRny0CngNPzxm22rqyj/G6bVP1ktEi/6nIqvCJYriGRotNfguOptA3IghS9
qVAlGrhTWMOz2WWnaKBCiezYIxsotMx05qmLTFbdHtnVyYnK5/w3E2AfkUXyVao3
dzCP6IqflQx3bp+gXdgkkH6Me0eVTScbfCSvEcBGh9LYUfa7ubul+NQ4h9E34qMW
ZcCf7ioxHBTetmuKZvrVx1oYZAdcOml7PUEYZ53CQEo2FeNzzrulUx55b4RbJUaI
wjhu+NeezgS8w4RfdewGEL0oVKypojQahh9cV7pKKf3XO1T44nFrb5M7657X4zaN
rW3uQCsJKsujN2eZADicAfMo1K3InT3U1+PBnwrAquKMOODirIbhPH++PgJyUI60
TSQvV9L2ABXAnx6JWE/Sd/ag9YFE9Qp0asoi+/88OIM8Y1Tq7agvRP3GIb1MZp4d
2uQE0DBPzzr/Wpp9kV8EBgozICVycmFPMVBUH+lEvLI/Nn8wvPoNzouK2vpc3RgQ
WIX7Tt3yZuD42TdnKqg7UrB3DIfmln/lnd09YjYYzWBFWx74DDUpgoT7IG5J9ZRT
/CrkblPjUM3rwqO/HkEYJ3y1ETci0jqaBJFPrJ+SLWL9obniz8sYzcmd3pQu/DW9
2dwEmf/S6yRGbyFbJIGdJkw/qexyA07pC8H5gLxDH7nrDiBezjl0A34qVHILFyGx
skwOU535IQSLGlWg/1CqOjCtcL6ttaizp9mKf/fvoyBxHAqdjnG1VWB6G/TB+Hkr
FwflubZz7NhlPygEY5px6CxMvw0T92LpwU7xdU3Ry3tyuO4OQmAysOgd7UfD9h/u
UXXjepoXfT/JGM72/VTvYpsDJ+2N0GJGSHgbwPPdbA3JIK323wFq939sVtSUe2ux
wf50u49uUZhM7H0GMRhZjk6ruOh4bWGMbctVs+TGozO8qCfTp3UuNaghbSRWQ84E
/820lzzjJKE5tmNQMouRMmkSkJXStRwryNW/CAH66SrC12KO1WQPGZKmRs6RxE7w
6MqwK6PqDbaBxJYMTyQVDpeOW9398Ngju4VQh76r4XzvEVJSggWx4UpjE7eihTOB
s4RcbFkpdd+hCdeBIu753odOz5F3arxzlzOXl01JxKC3KduQltSWwgXozQqVHWa5
BIo8WS8tcVN04pHPX8UCHigmmWIjM4OwsGnlL4TukPQAeicZR9GGB9HtjXy5QQmG
0FWs6SIV0ifrRZfWXDLgOl6bFDjMUmEEOP18+dJ34p9kfi4KZo5a60zd6HLRjAuA
frnsG9MWxpf4krCv+KX+5Ow7TwjmeBjwt4sauUDTjueRp4WnbsSMHZ+K3c+JMojG
5KB1H/jNkZ2bliq2WVpEfhkpQdT/67+9LivNpo80qRGTH+Gk7MvFaCAKUgTeKdTq
LE0tV/N1NoC9NZWVHlWGqA1DkLldzHTcR52wmJV+BzlCjL2z1oC/n67TokiVe5CX
PCCDnbiewOEhM48WXfDZTutTsGsgKN1WOgKaY5TvCRZq9qLYKUUrETEPUvFyf4AL
7mdcPv0POQji5z2T4JbKDuQmkOUzJnKNR3lWNnn+nKRLT925s4LV64FwfrNQ6FMO
3NwuXfAmKQ+l6pO9/75zD1Qy7YcTxnXAJ/IV+POvSYyA7aKqTGHEfXCFs0bOWmLy
uesDTQ/OVuNJwaqCfXPRQBKHMxXE8GeQ6lE+oGjbWmF50JRTqthkSNqDUVhkXPiY
RYInhUMSWNAeKWEdSaOsMM4xUP7hX5IhfN4NCVukUjyx7/XHie+z6wmtbr16ubQU
hpW36JBxIvsOMPsafP2NW/Nr09VaJA+4M6XiEPEei4ZkKEwU4e+4+gqvt+gHgZyS
T0re5mdbpp3Ywtj395hSzqWuT9NakgVg2N74UsbmrDAcS/cvGMoJrn6nEQj0gJOj
TD0BlQVnGyxVgyIOayvhD7RIJQ/zugtXOi80EbhayYd1kRyAi2ofb5AaOobbt636
/La6gJzH3tWXaYpD8fYuuSpd3iYUZr2pak1j/Iqwbhhw6OkajFiuZBXc46kR34TY
6SeuQu1TAdMBZ5RT9BrtGvRvTavQouTol5t3ULfgts/BiLGwMqGSogQL3+kwN6JV
YLMqeqEt4RNDCk5oVH36AnrIfHWYxveqnV2IsZF0Qh+rXJonzeDk2JgJg0LDP/yp
Vfpuu7F1+hexccTHXlV7xCQyW15PkxLVdFO2kQ9UI+1pvOxKnnBcgKvXySMTr3KE
wWiYvb8z/1rWDpAUbs46s1Nd5Tz05XPt0nxUMOadCh7Dk6mzEm/CqAxTVUvRjuLY
iUqXS1JKodVWyDjwB5KVwwlfUXO+gQRP5edx0gcUimez4KIj6fYv+Uvz5aEsn4qI
QKSHtROS5zNXu9oXbXqEjWGh+ZMrDYGwITuoSO7oEvJFWYo7BVN9sMm8oqfskamR
stiGfp/7u9YzVKwkULKymCam8QffwhjOtPv60ad1L94hZxWnpeAMehkojuQe8oAs
4Eowfk7lUZpGnjqDP/vg2DJPkzPxSNLQg+/BSp0wWZqixqxdQwl9ibBOb9hCJPeU
m26UZCOKQfyWn0gJnTY/KP1+gG/Ml3RPSecpReH8T1RUhR801lJ3agk3T321/hrk
JRC3QsiMMsWBUcPUTdUd6ySH/00iSiWvURmLqxB0oSdgaendFO96cN/uv4J8ap8m
WP4p7w8aVM0O2YCpxHEDLplS2wFToWjDPGodUuZRXShvctZXzvk1EB4oFdeSdm+c
qFdgFqaE+gvWGVmg92Ac8kV6N4f4Y/UdnsY7JohhjFrGKxjABL7nDJKxQx8HVEuW
YQ7zakvJ6WZ5etooWtC3+Ma1mNCcL4n57uqzex+2YqlCtZXCtiSsXkf1LhUzhrK3
Vy6U22VpMJImXCwcUunRGJF7eDzpIiNQQfZzExYZcMueNUw9AYNRsMziirImSv7J
uQ7KWJxiljYLsrnwOgWXV002AIy+gP98lys+d2erx1yIMo7zxhD9n/KnWxQgC5gP
rjr/e7QXQ1aJLtTsbbORbXCpdY5/AFFWBfLlg+4TRbZZsQ0KPKrwa2/Y9pLB4zKI
gb+/U0GUb6YGUS3WVz2Tq34pjzAjUz0621WkSFEYJ1Mx8x1ZkADgiuyLkpakUj35
cPXeuAVv/ZlYw94Q5WtBmqFG7angh3ZQWjI5W2UxW4U7MHkQ+HgLGPMG/JWOKEK0
0FVHgoW0JH/EuuAVt0G1qKZAg9TuBRroRAIGl9D77H0qwAGdjPsk7JvS4EM6VIA5
9zX6t0+3uQGokHEdsEi+W2ZMLTmY55wEAquF0mdtrqIPGPGM3xt38EZIy7azIXsk
/DOimn2M67vEX40qddXjUU1FExUEaqE2hKxo4wr3NufNfkKZ+Cviv2sut0uu92Ax
n39Nkzhp47KD+kysBh0bEmtQB+/y4hzzmgaZeYxmGvDVsbhIJo4lTtjPOJw11pFZ
tdUM5UiWfmfnFJ06GaWDxei0MjaGnnzH7rkFiNF7Mw0d3gvoAZ+zEHjyBAlhNe7X
l2eMhvhXR+L7J+ToNobbkUntO40aQQ0aPtTDHi8OCk4vJAB3qNLyqwu1fFSo6P/9
f4wObK50fIGjMSQvkosNcbO1JB8z/YMRGUiwlS7D6kPby7rUqFJYM7cLh6lbnXWy
A5/iEAqPaLh7gYnCHvqApS+wihQFN/LLEXerzSTpFXLDKxL/UTIhXFfVj/e0crnS
awad/wFnXZJW27bvsNKKeL3c9ZgP8ffAzOUkMYYIoaZfa2lgUAddoj+cg6RclxPo
2qKheCR+TFCSiapb29fsEa4UsRDHmGOt9KjNQ9E7Zwgiosm8O6BIA5ND7ejHqbWa
W2h5jflaBfYSrRPuNTR8q2H6JAlo4KIGkCmnB26BBI+E1L84+b5lJeLDL0outXCG
kmVStldbN8es3Y+uj5KTU/0jvMZw4ZBe9Q+PwLMfJ0jRwgetRZ7P6tKmy8shvAHi
/klq+45uLF51EXIXfhogntNPdkQ2zmwQcgtjaRIXKWLtLay4vaiXbdfw7gAHuK6f
Qp4GsyyNAdMg3sCeLsjoodkNBuyOUTLsBh29WUw4swk6H8ae2cEJ1onpFRu7lmFd
5S1c3RZPnQBQfP2f1cO4KRx2omfU73mK18bOGA47s3tQq0auvzewyOmriUc7MFGb
xTSoy0NYlByXOO0UsTgp98GhxDn1XxaR6lNVBetbvCi83AaOtFH79AMDxlb5iYxN
DjsNVKCcH4T2hPGN/HGPcYz8/w+mXRkUtkQiw5jaCA1t118FbpSdG43z8WeqX4PX
u1+mKv3na0sg2bjCT+srxzR/WiD+Uc2P4xbTtpVW54d49jx6wz/Y75ZWehwW/B97
iBafYs0kPqP4U2c7KUMgLIlIyYXcMhzzgyvtYLql953w/0k4hD5u9D6Dvwo+P7U3
BSZP9/ys6RPZ/tv3QRPPMJgt8VU6fCf8V5IlXMxHjF4doGgVY4c64SyTDSOZPKHC
ORg78Dv7IyXLFCuHaPS4iEmi2+r2zRi86dUfLdrS06KYdvUyaj0dEcsjug83V7/L
AYIqxDdzilsaYUVxZCn46zTfs4Ta6uZMEoXl3vR9cN0dSxV0dfFyHMTewB8POjiX
uQljFvU8NCFzpNbggcAWBfXdZgVWYaDQnqpT3aMaycZhKxeZHfU6Y6GwrNuGtCOO
F1PBF2n7e76Ts9HByn6NoaDT0VCoC+01Ue69AWyopjpKiSSEEDn5oXzUTiDULlkR
u+8l1muEGJnHgetF0YZdZH8T1E0i8Vl6QOs9tR9yNG1+BTDsRkb6rghscg7VofZU
M/UH9Ye0wQDsRghoI6fTqaW2KNcetPSI7pFXsDqLrwWGRlPtwgZu7a7xY5hHmsb8
XIx5OTT/TOEBByKg+vecfCNEnNFdy7gw/1l7cTn278dg3+MKkR5u3HMZA9FR8EDP
B0BUkHZjlF70zZuUNCliKuxz1lEfZp/TsL0Jx5bsVDq3+wCp4u58ibRLbH7KQQUF
V6tyz+vcJNygSsijRerwbmNq0/wUdSKxZxmdyl86QVU3QbfLeZ9Wzg1yS13gLM4b
hVf7iQaDBD58ivGskHC3sWcyWh1lfBTM4kIGRe8vJyseT58uy0ow446cjy0Facgj
bBwkjwsaXD7khIyURzA72BWBQ0jWmK/BW1fHzKlXkfDKUlKIBwwsW8OrXw5dvt+Q
RPyNVO/krFp82f0ulFQh54JMgnJhMcJINcM2NVPEU9Hx75CV5n4+L2LhoUZheI+O
F5o1UEbvE8om5ghQm5L1V7YsiHBxyVJIta0hmaP+uEMjmSX119Sk5GpG4W2EGd2b
1aZs792voaedACVsLBUE8gmsC4IgvGiMM0q61YViU86LNTfwy2r1JCe3QZpp0UWT
vIpyIb9pTBZSoOhOBQX1WPHarwBrM+nmJQezKNCVVvLrViReD8kP7Bin+9buL5YM
Et7Xfzno+DqJ9IxuNWd4NXWYLhzODOnySgbWUPDtZ9isRtq4HxcVEeBw8d/ZwFlM
keTPTwsfcTpCE03syzYWhd3kVMnC4wzbeW5e1rPJcMpYqVr2sh/oqy5R1qQnZ+6N
ZVc7GBsP5Y9jb4KT8bKRO1TmU9ZfUSKbJFGgD5kZboWyQxsXtJ8KyrlH/RXUHune
Z9tRMS5wPb83twOWsFQ+09d5SGHmx0gOXA8A5+r0AtluUIHtfMbbZS4b5mSLhAEQ
pomWEc6EPD+G0LGPFjUhW5QkJre2p1h0JrnuWpCxf6Hl48741UI9LTdrTvJSVKZQ
bm5kwVQ80nsY6KAnFZWWZFyZAITqaqxYlgQn2d+Z6PwrChE972PW4iZTcbxkldfq
Qls3mxTrY1z4SNHNou2VH8N/cUTDMQiij7XsCvGGucg//g/xKiL8Lgtiu/ZUNgKV
PQQ4gLgpCV0l7mwst+IA/2fVFJlwP7CpKGNU15ucriCUrYfQgpla2aBJU7gQGiwF
TPBJXaVe9HDf4c7YziF1Saz9QJ0bg/ddhjgn4C1qYpeb55hX8SAHsazaS9bU5qyG
hz6gdC50ELMBVrIrF4nb8p+62zcXYgwVmKXOIt5If8gU1R6MZFcypQmV/0aS3Hc/
MhAkF003dGgLsQsJmBm9k7nUAutWg3KMzxk6UjtGUiD26U/i+nTZpaddm/L6fuW/
Lj175RwBiyni3Wyr7I9XUBQLU2oEmUAOGzdVjUkDvFRlQw3nTxP8sKDFx2pK8MdU
tZaYVd/pZjDcQpkGzwUYBK3fDgsfU4robpdlgMk13unrOz/fzMbKUUc6GCccnbr3
c7fhtg/DoC6ymyK6lhWVqW5T4EzC70vPwRXInAwKSLjYR0SFzfby+TxncSoabzsW
zyooxJ5uqANPOwgTKph0oXLNPt4fzl8i2WAjz3HqyGkFqLspoFBs1sy/pObawbIw
4x2HnVG3sjrmAnxlZZw0akWWEh+LOzODH0Ql/O3f5SYYmLE8H7MqW3KG8F1s6+Lc
3S/Tuiv+zhLlvsO0ifocnPcpvgf0g/l9U4SOEIKk7fXMcYsWHhYSJZuM6FCeDOYr
vop+GXO6L11kd7+QbEKN0+xAcKGc9LlUWqqrGwFssTLiWlQJR2y7JgNAzRE4X4/b
Q4Pqa0rSFsd9nMOFKo6uvNSwlwH86iKUH733IYfWoMwQO6a9imOP+vFi3/Eyev0d
5pj3bva51XyEvQe9IEHxFXYIPABRbe7oyQdOoaiF+Ysl+Ge1Tlo/iDqRTqDUKI73
dxdvWbw6x/eMBrgDrggWyRFEeqsbG7gXhfLpSzfrSkQOYq/wi85Fs8TyD6kcFU6b
gzlsNrVYTO4E53PbsLUO5jqw5djhIwWaJBvOeGArmvI9imYrTuzqNMyLAIyF+71W
An1pM0nxNUqfQP11s/wmsc+UWYKEZ0AQey7DRwLoARSrSvVIRU+YTARvFbJxKcE5
zjVyga9QAc8IMnpzqxtXaUrhcr5Fdu+7SADIcfTSzydqTpkUtJmgFCs+DAOu65O4
ZTTgW485mb4Ed1xw8+limAG1ugvUFPXwGmCac9rkrltcRgr4yBygKxxEJLvGiUjN
P6qxBBhpEbuEdbkMYKPC7ml2UUeTVwkTyD/abB0Dk0bHlHpDUBJAdtPbJ2OClvWP
B+ukq+HPyRhoCaMtAnO5dAPRcf7YCU+O1khTd6/DhdhdTIXY2VpezIR4zVG/1RgA
g+lKlCAw3e6id9n+MFq47V500WPYvrQ2KmbmU7DBtXAi2ymzfajjQrTawvKWUww4
1RZ4wrvI8gWUgEliPSqgRAbc3GcLIQgXVpopT+t3dXBt6e+qhFJJuJSRrX2Sh9hS
NCfNFMIgKDP1qWyexILoZ/E/f2BIqPBKeN2l5Mr/ROm+3C3BdUhhGjnfzsXxpyuG
Xw70ppNd7PKdn9gxQSKYJkRWaT2OEcJ0RlumXNcRbRE0zyvkVql1fNteXH3jsU6A
dLwvXi1Rj9x+F8ll0eH3Cepw9HQRMZovQOeR1vTTHGMvxCj1+neESaYrHGUA9puY
IBncP1YOZQlhj5pGVrDY3CpbPJrO9Wb1zAEjofnpG9jnH6hoYS/5KD1sM022N9fA
+XLQq+Hb6uIZkf8mmFp2xQHOBdMPsyMmjhYU46W2IJb+ccSim1DTas9VHCBHPcjS
v+K4Ti/gUxqKEUb5RKzPbPjBPt0pwmx5Nn/60t+iujw9nyrMw+J6CbBnFIg6t54F
3m79Kn0nV68HdJwFZNlNmabjic7swM1yxBh/ONn2zCW9/xdR4XIwJtNsmuT8NYAB
A5v1OS20jE8UZJxQjQ9hGiDiLcCU8cNuYmKJ4ZFKqc72Ry8oscv2V3Dg+qHehI2M
DZO2qTOMQXM/hPDuBlt5b2NEV7OqYbCmScWwtqvLAjkU25s01CNNDtpnFaM7AKYM
uD+thDGYQfsY0YPUv14GSLRUEsI3blSktqGLz4veZ8Oj4NsdConJikypK9lPxzpt
CV47mQIafkWix21pbQ/oAARXBovVvfl0QN0NQJ6vNC1NGccgdRXgi2+QbrFiJB64
EDCnWFv1qDZa3ZvWLvTR49Jk+EOcYVKbkR805AdLAAnD0CVZ19PCNt58aETpK7d6
Rdf87A9TE31PqCumb1BbAzLj5wYhMBXK03TIvUkhh4bfnskN2XhLDjekD90uYGY6
cqh+1U858kenFFbgx610FHSCzM2NukBtPkrtk0GYqxd2s9ZCH45WUkbvszTLJDEd
xGVeLCxW+XbtZRBf0ZlAEChugFdUjkQkskwYKXvIpGLzbUi53gm7bYv7b+XxuOTa
mBYybn2Hb6nc/syGUAI6VdrFFj18NfVsjwJSBGU8mIQHyga4gCZVniUsK4Ty5NAx
QAqnQx8LIPCwWn1jPulCKIvLVunICa0P46B4dmpof79jxCjxki/u37kqxzbtKEOu
ryxfHKZ/acbPPuMAm7YD1KIytFawVvchcbMGNwE83KfT2uOqjrUr8rxJBfI7tf00
teUVTBkOFay76dnAW6Bt8TwnTdB0fc3tnwyW/w+biiDl8gp7J/kk9jNI1iebkuv+
8AUGIxcZW6rm/aV9UwwqiM8pZdISbhUh9zGtiZhjhOucwHyz4yW7XbGSxpDLps4S
j0tROE/4K8kQlsxzTJ7bwrBORjyPLSSLSfVryyUDCi9dm/kmjYPlgdcmVoqmEFYc
YLLEShwbOSF+xtsnnZ3gkPFwYboo5KCHsPh/ll+0COrxSE1/jgHkafltJMlS/UJV
+4kUA1w2c752APrPJx/eHDUUPGbA8sx1imRfZGip8BP93iFGkLRyRMe0N+ocK1Yn
C6DJKU7j3wNelf6XD06+zpnqgYHOe/rlGxxzGM916vQxJKRGazNp+hv0J5ijZLit
yJ4rXwJ7/222vQzeT7gGlCVMIQozz0wCJW1eBIEQhktibDiSa3kxFgrQ8HO7O9DS
JnfAUpkBIdeH/xki6ldPPICWvMbJAq9RmkBv9XJCy1mODwfcXS/Lza3AKiXAEK1f
xmvXSzgSkyHFmZh4oAt3lnQch4QgXj+NN4q9x952w95RxuIFYXNY+KehDcTD/JCO
KG+3crlLDMb70fS++T2d7ipEw+7lBb8I3TTejPnT1iYlLV9LrvlrrAU2NTh4Z2WE
Giveq3A3QVoz8DOcVXaRFtWbQVnvinxQjS2p0ppFYgYB3wXk8hLbV4cBGZlWHuK1
rVtJJhLZkLaS9g2dKCCRLGSNMMPPcm1H2/HjgfjZHNcWEGBkU2gYsSl1qBbuCSQA
ycj04KoMiVtYhWG9IG82W9fP1H0FjJ0MCrCTiOwK7NrSrxE2bKdPt0L1ttSRPQhJ
WBLX7Sei4kmZKS3FaaubUOJBzLX71Fu8u40mtXoyZZT3ozr+Ms5Dmv4COs1l5zeJ
EqY4/UwRlAPsFAS0Zv5AoiBqMy12pzQDCKpozmjd/Rv5TosCwdupwgeVFwA6fL6b
CDt9Yo5Vln8/53mQWh03y194sqfc1aR5vxsxqXNZImxtdAv5RjBOdXvm3/+ofv9l
65HE2lWwkPlBmTaBbgi/XQbZmTi5JZAz2leu4jI2lW/TPC37bph9kLtYI4Ivtu6a
klhlrupdfi7QMU+yIknOjGGQWQxANO6CA5VuDZdDuaiqx6rMVXEi59xsnpCHUrfQ
deBRA84CTCDiG61rY3OxPeTAyeZzHvxggcpTbHStBkv3oPcVkxOXmZU06tchi2Wq
dCNPx1Z9p+jqpH7nbNHqbcTgspwFnJsmpegK3ltezCCvD1JePOamVYXrVbyoFIlM
qTNB94PVj+Nc8R59F/3+eNpqvO61wyCyePJ5RyD0Kuu88Iu3kfF3LgLIX/qiefPK
MIJDps9DWq83e4CyVp10ouNUIROfXTbq5IX9fSBKjcqAuRdyXxtKsWzCeK4lraEN
6HI4HMCzkaCKN+kL20pJTkyL47R1kWVPLPVg6V8/5MM5YYYhwq2ZW917Ydg+a7Gy
vBch6y1+F4p8UIJPWwWhNS03ur5oLHKS7V/OJCc5HeGVzGukQqA8/NDwRCYMnqdm
IchVLPfOUwrBdZ48RgS8gCKiFVn4lxkjQCDFX1EhjFFzpqgYSvvL4IILkkr32L8W
GduxxnvmuorIgsMhgxgN4WxVqDXvj0sMSqPtR++s/VMUzFukU8gD2RmJvcM7Thfa
P4VdB6rX3KJUXdINthn4KAi+BkIKBqHBaVR8dw6fdu3l3ucdx20gdJExWQ6cE9kn
wDPRJMADOKDlVNPZ2t5RIgTIM6HLWH4l0oi6XvJU0f+mih+Hua9JYK1/JTwSb/VX
5cq1kUnEoWO0/i0y/oeiQmCWgYLP6urGGT7SmddYZSrhhraQxaztpeHCc4EwsDKH
3Mn0CJyU5dkVlSPKHAvFPeZ82V75TMbKnuE4c8GbFhe4BOLS36xeQLHo6ULxD82G
G4+yNJ8dnCknWfzETpmQ3COVZCZbSiwKBykKva7rXxlQWkwTZ602HcIF7raFNzPu
qXjSn7TwiFW04EClq3jTDlfP5qoS9BQMDciDX/ImuhD2gdX/DypSHL/+yUjy2tSF
ZhU9jP9yLH90xzTeZQ4U2q/rgSG+xoKqKF/4UMffYTMMg6iQvpnOWSnmpLeBzk3E
AEiBWmhVc2zpVtznOB/8I4/25XS9eHToIxmtJNtat68OkLrY2AI2N4Mb6w5lVKyD
meuAQ3B7gglkJ1mLircdO0j1JkEI96RXKvxooUAGBdVm49eXHLZS2igm2YZChKtL
LP9w93Yn8wezLlR15GiNF+5InSGTiPD4kDCmQrYVWrR0g6Sx52ZWUfdUSzA0ae2X
IfYZ2QQie9RkxG/yU3+hPOgfjybq/cBJR3Y+tpMA4Y3u0uwmftbNKZdm9LcxbQxI
2KEvzvFUKW+BC6UG7tRrKf3rY8F6YriztNPDLdOYXPqpBz3fjFvkD0dBMsICuP3a
/F8CdiUYPMf3mt6jDuDz2KHtiOht2Y+M6++tNBr6L8E76j7yGcJIvkCNuVJwpfwt
HATXNCz2FqJBKj+2iqlRvXuMERFAF3U+vrUd+Veeb529iNBPef4mi+2OtL9jxaQD
llMrsDZJvuMkdybYqDC4dHMk8bhXx8IEumqm4Kxk471CaSgXG0gEd2/Twf4gU6Bn
lKkqSlZ41HD0pHf+lM2JY2OYSU7QFkSPPs+3W0SzXPCZK8gFVXp+8GhA83EFQHiO
L+sevaEX+zplpiTOkZoQg5kRsDUSQkO8hIUda4vQrJ+v5QIiqTKS2row+atOEC8N
gMG4tpoWRt30k5b5ZeQnk2uoJN1o3oSG9B2awJSzLnRlQtLWWimBKavu92sKmLYq
j+PhFPve+unB3bVFJaEOagVkVZY+39BMA1VptJSCq3GgWzy5unD5RkbXdfkXPnox
/x31f60/3+EV4Eof72Q5E4wQaJTbmoSNXz4/fxjtSxrKF0FWef9o3IOf/0bmhkDS
tlCZnOeA73e6/4yzbqH1hCzulv2W+Gno0DmZJey5fq/Rt1rJAymYuE8FZV4XL2Ot
zOwIzKdRQsNjDtRKDPlWSQdPGCO10t6DPLsgLKaRNPDSyNuxEYMlckmsQSAdratO
SSumUbnWrYX4PXG1FJPDyN7TnK8FOglqOD8UM3wsWIQfZK3j6Fvs6AxHeH/7t/3F
mcYLDv6IUxYVvH1NpyxI0JZDm/lesIcRUnBe/xdcWxudITi+Magph7MMxLorNdMr
lSwc+BP4LFvPVVWrw2ImYrHMSRw8zJ/PfbUGLDh90w12wh2ceESS8//y2L2PMD4K
xtzA3yjQrNh8Mk58K9C4lDTL+QlVE2HOC/jCub9MFssB+QQQG5agHQSwy//hImX6
xjz7QOky8B/sIhmqzEA7/xm7wXvpvB68s/O6iIYWZU4WIlWLmoeKNa30gKN6ERM4
H4vq0iVP5qH16gNNKshNfOmGtQr4AatQ5zRHC1uAQSk/wHz6P5xf8Umy9e3Um1x0
hKg/uIoyk+CNvcKUX4rONqNx3jCTXRCDY75QRA00k9cvSWCUqZj3kC1auOaU45mt
NNvVUDMaq8zSSU00cIqHiXmxvKSsmTInggazwG3cW+w2GQ2TnCGd/ECQFwyiGEaD
Zbi2w9aqnBVKwYGAjDhoRF9fOMFvMqbzc6P1cKpCpq/TCM7wP7MaCS/gBnXDi+IO
L5zDAi6tGPKnXWyLTze6JEUnR2gQUsmt7tZv8Qj+8R/E8yWLg7UXo7E63Q65Ej4Z
GuKeFVP/y9gd0pJdtsHaJjvNCubyBomGqU7U5y/xxOMT8A6Hhh6IzNjTRkqoQsOG
DOoVgeH0JHLOZQuZgwNu29oR9zrWSDs3qu+lNb7ASElHFRSiTxwA7ln0+jAU54xD
hujprJcY6YIrtP//sfgIocEJf4jBuf1rjdvO3P1E+ZLLkrxdxZE8optFqo+nBaUU
OlDpW/zhcwhVCxdOVaGAlLn0uQnoUPBDfUtKXq46wGTpMyTsLEu+UsIl0890qvcS
XMMfWKWTbiyBTLDZAi0OOnKkEAhNTXJYmY/avXfkySAjY4G17ntgWbTPsBhYqlNd
vCNI0oX4t+6BrGdQ/CWUuh6Rx5zvkN276+nCMwvO/tuzUpuUAnxmv49dIVz/mZ4z
VQnkgnPjaPSyGjs3j/0l8BcMpWonfLP4oIwqkVt1U6q0FTTuSxHYXAiYSy4gh6Le
Anv3a+6PIQKW43qDrMX7pwC4wNEbreEHDEz8jf4LzIasuObvQD1Tdcpnet//6KvS
flQyVIaBeNSUM7x3q2Dx3M3eJsxFy52nUHsdpow4Z8pcItEuXYvEDJAh2CKI258N
z9qVO6lTvVbmlbaAfTPObqamEqe5v007rEtToXbG3FEI9T3nwldkvBgz1VCQKYTK
St9jW/sDoYxSGvumypoRWyAPnnfvmhEML9AA0TvDoot7X7mqo8ybv6awex0Im20a
pazcFLeD0XYmjAPF+ZmQV6vKj6VYID+jaoH9et7iBW+XTpFwLIc7YIa06yokiaoJ
txCpwZ1YZ1kZE/WJMcukgoN+bpOjIY5dj7C23eerSjkqZG/HGPB9e0YoFLzUrUwH
NxAA2kiBRCJjjeY+E1qndlMXISeD5iGQsIALd1cOlYRK6nre3GaKHGUdXkuI4E2u
TeR8JQSH5rx20VXiijBy+6ef8ysxsFzZoXv3ctRAe1rS5dt27fcGk2k2jtPE/nDB
wskGsrkbWNpZKSjnxlApiDgtHShzsjfk5Ypo+JIXdWp7oitbmvOTf1i42DfRb7Ni
46JCc9eDrA2GEeGqw+PbCHdjJvZxiBPVNHE25tdO0XhrgrCzRrC13J3e/nzHiBYR
qqUYeByIpREg8WiZv09Mgo1S2lRWt8Bfr1NCJl6Mi3UuIdOakeHG0UbTbp0idp0n
Q4WxIXSRUXClkx6OCJh6f2gYkNOUK+fq0Liy0F2Jd18raVBhcP0kVOUqeJEJS5oo
fVyw52lUDbNA/dkzdyRjKozj6zNIGi7Lepbv0ecGqZDnDFwxUsPoprz+BZ4krXoy
Rz8HErgg5W5OqUi+rlojDBeWdVRC2/y9y6yH+btZ0xAOLvQCfPpau5C2SceqoidM
pUeHG3OMrEhb5r+WAub36Vn3MkPPQFQE/kHCyA/wc2EaQsE05fJArDZGp6EQ3VoI
a//LQ6g6kQC6d/pcpqSZl4CUoDtb2q+WMKjKo0CnzO/x5SeRSTVMmf+Vc7SvSPFU
xOsK/Mn72f0z3N0EIHfIEuHxZiKor9neC/TnhGft2qN1sI5FmdRGnPT5VYytVsPq
PNBYCLL+YLIR8m4sy6YUue7Mji3ZI89Qa2VnOSiEwKi0fR5EogwAXPXiz3IDiYM+
mORTc5OgKw24c/QQSJ0tUa6iP3m8i/o9xc4SPxBMm8b5iDVV4ODzvNhKlUpSgQij
A/t3yeTQxsmswmdE97WCCvRAoftWlopTevR+MleBQ8YkswMueDD8O+q9vNkGd6T+
1r8LnbcCMj2Rzpp1FRpbwgoszIoGsz6WOkFC1gn7u/s2P+QsvaFW/ZgEViBT0iyj
EL48P1futDWCs8iiLCzus/XfTPb2BkuL2FtAkwh+nAoqIa0rmHyy9y8lt/Y9sLLg
EjcRL2caBhaCWQYfTFHCx+mKrxJfqMR4nDiJsvoPLSemhh2p8goB+JX2mf6rbE0I
lbMMycrqlUNM4p5zGEgI7R4XIdjG6ofjLnM0/wcuC40CU73yFfMBMqharzBlP3C+
8ePsN8kMGVy16Ohd1JyttmsJeexWaYvjmUfWPrmJk09HCCZ7ONbMQP/ZsaoxmAVD
TSTAOuGkq1E2G51CrfKC/LdHmWs4aXTnUrheMTlStrJ6+dwjzCqNUO4KSFfJI936
terd/RDsUMMKZdGymNcyeabeYsvgDNA7QkLdKYsacIQF9/VleyrQt+RYUY+JTHVm
urEAHIwAYVpG9Xo0yiHdIqzmad43YijGh9uaoE1ww4AT07zFnxGeJARgPJrOys54
jKfGO7UQgSY3ZvLKo2QDmaqIuca4f7E7POM1eiE2VDgeb5630qmABNubYIYm2iRI
nk6v2kRPNUjHbNJM3k24w7PXcHp7VD/SfO6gvYaXVuMmH0JoT9a+wmV7aKJq7i0n
I5+dkky0c/vJfTcAi9ZWoJ2C5TyyHkzratu/DzDZepz3uflkmGLqY947VYJ9NLq8
GAS+J48zKa4bF5UwQkdg+TMamz+GFYnuTPFqReuzCMQZAQdDNy3Qv8lJOgA5+ZK7
0Eut3fCYStcgVyefDDrEnOikd2Kl1CT42W22s/BUp7DFGcoR2uZmzgBvH9SCP4Ld
TDT1xpGF1i2zBWhq21q1SuPccQEone7XJMx+PjScQHVvyeCtowsmStMbrK7vTNMo
/R2A/kXO94xtLF7/HPBbffP939xd342oA60HBExykg36D+N0om7fuOXcRg/2jA0d
qT0NtZkjXucJiwueTV8uwepX3ZAcIi1jasGNqnYQCECYNmBFaTrTIeGPgkASo+ZB
F8HcXmnBgJfOyaD9FBL9Z7r00CEsU8gyKu3HAIjBESMZdD+Lm+1sT9oJPiDHi+94
yMpZjmK/NiNwptEro9SWQjw4hf29GibiLITf9rxHSRAcfg7gchTi71Of7ozaOlB2
ab4WiG4SLzhpPezqffXOlEGz/KvVGT3PSXzkn1UtxuavQ23SC2QNeTf/klp8o6jb
ruKLDBotV+6dFgcg1ki8kB1LiI3gqtyGa8+2AMRYrC78pz5foW6dhKMJiXssHA0n
kRiFprsqZcQwV/WGs8yzFUtSrbZIKgVnotDz/iHeq4cx1kirTtOujb/1JS9Ob+vr
kNSdxD+9ZiDlbIOat+F6DQnx3bbCsKbBRVHOBYHRWTjIn7fol+NdGDBKNnT8s9j3
4XEcEFzgNewOQRWhhP+NBUUsIeuHK0YYmeWkEXia9qrSivmUZG12aArZFMfSBeOz
rSSAPL5rRmpx8EDirQUX7hAQxChDdiClNUNihL54hkv2YYI6F8APSkW0FXh1lo7U
9cvolLL+Mu86rr78jmp9MFbxyvbdPS3sA0h6rJ42hO8odChA2pcwmV64XQ7c1InT
RXjT2aTCiXgTjv0sej5A/68K+W3HHZfCVQTD89LcN+ptYhoSSRMF3kpOPvewh978
HtIGkQc/ueSWBjtXcOlc3iZcwHruf5RnhmNAmp8z4OkV7PDFBiksumqlzIwVf2ak
F6oSnSEB058f3tcIS2/LRvJGFBsaUJixA43mh26403QSkJtbhNqvp+DzhTvO3Wdc
c9R4tIe9Bez2HmmehlJiWmQIibJ5H8on9gwOpBsnXf+fWugrBxFpHEZbrONORdvt
V+tCynBypovuxjogvm2akjYoHmerIMeM+/xlzQc7UFG+chQ6cZ1iNTMONl56g1a4
cqveP2U+bo0kwAA3mrPKE7MO3/BRJUvbL2TfuIhpT4hpD/Lrn6vg0EL/29QKU0K+
UvjwENwE90WD6X4JUWZKs7QznczVHv0+ufRt3tB9bWofzLJVJxOPUnnms9kXdjzI
CZcAQCTCghR8JznlSCpBJPkQyeldeDLhykG8iSTEhDPmbhkDzdbGYWPL+nOHRSXE
70E6FR3DIuptWhT9WtIlwg1lgenc8JH4w2b662g1aT5xbg9qbfGwtYvD4KT2TsE0
AKgqhpBa5oHhgiQ1RHpML3H8iAywi76RjfANbi3isMaqlcMR+gA4NU6PmRa4kE7V
O8TXXfvwgqW81XkUPksNBO8dmwlMKipYs0O37v4i3JhZtd/9vR044Qbi1Y3ZLe4c
DUNzFdHSTyjrbYJIiSmm/W5TSTkamC5LPP2ezAP24zHIwA5xxAu4acWdxV60P2RP
bbqxRUOkfmz8WQWnC2kqC5ydOlFMiaS04EPvSsJ5RYxGiu4VKvmHx8zYdsgSW5g0
2vGLJBhAjCqoKkT7SO6LEQlaSYa+xQzViPTMdwCKHGHfKEAT79MbY147OO7MvCqd
dEQDUkgAnlFWURrc74KA/JB0tLVixLSGPLN+b6OoIDQVJTwhJ+D92ChtpvudWThU
waH/fFpLWNXRJBKDe4uopyNw4e8jIWMHNp0vCLCzrjl32IECS4NrnebU5fKjghxX
Ygh7eN2X/hd20vgV6KCFwiupMY5RnCyOCBzB4RTAG8PIDKkmzJXyNcTQnFhS/XuC
Tx+qEWxSx20PCJB69DLFHmPNbvagHmuoN8LglbJXk+YARyxuL6FxbLIzdu6mRpb2
8S6UGxmxy9v8nu+mqXuqvVUE0nEQeIB6IsO8/Cj6iUCeOdIFLPZ+NvfTjMrSFCRC
QCQFwypYnkVDFmvTmt6WrR5k64mQ4XOzHGTLsoPkTFb2XI2P7bxMuJOUdz+xBPMy
br8517aVn3yrFLR6RDqOg09c/2atHtHxQnKaiJdtS3/G9LV06zJOQhz7c2GCoUv0
RJdAAysks1Zr8ogRPwrlK/XkC8gci8gRrwHwTAEm+oS2COMNjZ/IHzLqmzMUT2Lr
V+1F1A4MsVPE8jQOBhQ4QtImyXoxODnesaUxmM4ahWM62TwHnQx39UduC0h/Xb/D
YBCkPwqxpHvQNqR88A3iFZ/Wph9wmU/rfwYdNezt/iz1ghOfA+qKSLuA/w4Q2xfz
8ra55mkPeNjIsZLW0ZbfpYymRsM1hj/sowh/m//5hH+LhNsFdHXJGyz05b5I6cA7
C09ijcvU1UXzEfr5wfK6EbzxYP05IZE72M/fp8RHEsEg6uKT8/tozk3Vg+osPR+D
6z5T/U1iWYon6ffnj/jmzxPLBt8nxCAwsrDNI9g8ZPKZntz3/hqTDJdIgpMTH134
/V4GW3MBTf7FJYGQ0P0IpG2oW/4fx7mxJ9V7WMy3c3SkDA0/iLvSzaL+FbPCo0fW
YJI+SI9ER2+AgwYBVBoqNj42vxn3TYaW7s88H/KmgpfVCZn8ZBWD0K4VPWnH0Tf6
s0a7snxcIcxPoUobEJMYhMmq+ovstq30b50064CQV6pUxcem5S2EHCBZwqfK/k/0
c6hM0mLHfIFDtSI1GjVCONGvfpKKiiEfOY2h1PyrTcNTDfIicGcT6Ck/ksY49YJk
WPIoHOMMvjBXFzEcS6zJKiJ/12zxGHzfFbWMVEYD8lIFDaVLXJgboyOTonbO6Fa8
T7RRoJk15QFHDhNUqsAaJ5AX4CndeYC11osLm8+k6Hj4GBPPKYsutoKGr+VIBdQm
1wl7OddpJbUXobMMnsJe/1TN8erZVQD0UkXUcSbcFgTicN9Ve3cYOpXbvNrZVdD9
/ACYRzLvXuvv435TmEZwdc2pcOspp9IiVyuig8X1EWIWQwoMyXLk9KS7Ykkk04Gu
5Bml3fJf99VIyP/bKMJLQTYhIbmddvfDti8cYrAStmahZh2gb0JAJHJVY2gEg0pq
KVec53Hmt0xMF5jlC5O0doro08KPtpAVjYE6EHL4J9FTa/Tyq2NNA+Ycpiiol6oM
m1ov2SdmauWMbeiK7o5Jb3Hd3mLq3srE9+gZGaHv4cbginAbkmYFFjgVjuuq9taS
LpoiTyktCDjc4hR9KX2mp91E5ipvcv9VXGJQf5Fx+qgP2o/qM96HMwXz2LI+OH1U
qL68UKSZ3lfjF33UXTT4rbM5pt2d8wqyd9djZ+Qw+smnhXenkh/BsBo27hj/NNkn
D3Qkx3KguCiK2LDJpMtdR86sag0JKKFw0MYBk2ZQmntkSC4XhbC3p65Xdye0Zr42
OrtAvjPuo7kKtbNYpT6W2SqyabDpgBgKbsc5Fi0PA/KBFthCgexe5DxsEOAFyWip
aRNtXHTvGRoJILUG4F3bpbafbYOrZZ4zCoVUDVspkLI3pFU4lsf3bZdDv4ldcWKB
qmpbh7DRRBHD14z8Ctt5JQ2slQQtj9NXxQ72k/iP5NrSGJhM1sKVIbRRzv6Oymik
UqQPw2sjGnXbIS3IL9J+roBgYEkhje+2ZRgA75VX43kdXhZL4Mzc+kVfwLQfHFMm
dIizPeEBcpBodLReVHx4FG1UcB9V1GaeECupgy/pY7HlvHGbM6oZ6zOe0laEabzi
om6b0ai+ii0I1ndI6E/q1DZ7YfHU2JyiKpw+ZWlE7ic9wF5R1SzR4QLecSPy/4t8
3K2Efe39ZdxbpQgu51rYgv9FZ7Dc9dv25tcqYOmA4ZiyW6e55uq7dF3+5Lrx5+Oj
XuYPOhagxPYiD7PyWDcAFr/BORUSeG6KzTYTPKCO90EUDInm9G6vneYJHaHY+bGB
lelYH78fVWxURAjqJbL3/uXVAwTuJ75JBW2ygAxcrWvz433GRE/crIjVcDXYFVbD
6eutmgeQYTqEFIUxJkqzPF/qw6nHWd7U1v/4VbfyO9PoG7vUjIOYQsETrq3e/g4X
Ac7sQPLHEwUCs5j8Jd59Xv1PbfhpkAF96BiWqVRwFjtPfoim9wV5dHX65MKMDyH3
WGLac8rXfSRSsnXTOLTMlrFK283EUbagYVIWO34uYfw1krupKo4tY/+g2I1BHhWQ
q5mJ/QwLyBOIP+iAirM0O1COjnCMip/mPWiL2zOSnHeLfAc+6gztF05F0AQiwiWS
rRkJhQ2ykbGHGJFO/Nxbc0nFBMmzK4gA3Kltm2TAsErv/GJt4mE+/3YXgv2t7kbO
DUE2IzK4LBX/nMnCOBEmh9jE1QDW5eWO4+Shf0rC96gqzpUQbrtKpaPsIgowwF3A
xvwx/EHTp2MIVMCehWYyhUveWIl2nWF/Db8WTOElaMnT+eamiNFmaUk7h2+XLQHq
HfnjtFqnalcaDWKGjFYsey24YE2Ir/OPZmAy/ZIvU1PBRNaF0P3zAAMO2+HGZ2tk
8HoxXBV6MrmcPNRTTKY/VL62N67szxuG+L9HNeyBH12fk4gHdX0cNEuolLZmFhrs
PHP3jzP0mz+StAoUDhbiNQYkbVkV/DMfybuis7sxk6snRg4x/fsFFSuyVrEESt3Q
7VdIU7RdFuHRj72ErYEQytZEUwUP/J+FwbKwJh+g/GBvFqwa4ul9lb5kuG0MQ0Mj
u0yvd5IWWJKx1V09xJB1nXXmlt+wFuEg9k8lf9SDYEJbXeaLUBn+M9L2bQycR0ZA
rQsCKl89KvaGjea1tEUKPw3PniwDI9W8cx7cxYRcXndvbt8RXV/lBIAkmTn6Bloq
ITTji2M5Ivh90lToT+3/ppRZOn2e6Ih3bSOiFaxzihqYUv1/vOu/EcFHkc2vE+Dc
vJkZSsiOr+Mg2/SWJpNbmx0WjkVnMyzvzSuHawEk9Vvjro+Z25hN0G/gnC2kMj3V
Et8jf6q9qqHU7C42cpj7qAdHAWrYPbDiAVqTBxcdmlqMWDkQRqV2gkhh6ibxvbMK
D5rKAoIqq/wxT+NipZI9FxAy9tH6oD5xpoZ7S20MEU2J07fKGqdIwasxqoW3pB/h
fFh2+dF/SF9QCmDBZh+5/J5vJkm7EbF6QmeIa2FDgEGgNXOwGjReV0eLdFNUd8V7
Eme0wKbrAeQlggZNWKOKxeN8h0ABGAYHjvJnPne55XIInj0JM/nCjerMtMNpG3nH
9LlryyBwIU64flWwcVneIErXG03NM5OGMKqGiwMA4MDbYRfeDMrYBSw3rzTgFTUg
nJO7HeQY7ybUV484iUhQzQlldoDNWdmRIf3DQS/lQwM+IJ9v80++0PkVEPBOb1Zp
o8SEZwK2/5X5Gvm0qnT6XB6KoAVKmPK5PAGQOJUi8jHpzipk8zQ0eb25ZV0mfSCx
OUqn9lhnbgoDH1hA7Nwm3KeCS0tJ0BDeb4KfOQiZtwRiZuio0c67YQ8eaJY0AgZ5
CcXV1nr0zdsEo501qG5vh42T322iob1+3/lq4OGcSrOadiNQPIjnr9Ctr3lsMObv
CesU7ww5KDDGtaoiDrDlVwcly3/XrOeHMAdVIZK9HK/uLgKGyAQRU30sTw2N/euY
W1aGEW5ws4Yw02udFZxFnUEnxrbm9gKX2SIlKrtRsX59SW+l3R9n2MEZ/hlmB/+r
UWgFb1gVcWe78qcF47O9zQXrts+E0o5bdrY20lKxs33doNqlKvD/i8gL1qAhjxkz
yYK4PtdCmxOyBfGTwMup44w3MdQQILKLK0hdv/a3G0VCCkGNDBmwaOnNyqfXGONa
LluPD7OVi6NYUPWgX3Fn6v4JxvzHThSo4fQFN+KU6ZvfhZ1MBhTFBpdKb+Zf9GrE
xUPcQndHSUeuIg332KPv+wSEC/9F+tyAut/VhYzSNOMIpwbjlgV88cpQunp+TDoI
l6EQpXTSomfmzZIzirKVhgqkxasZMMoFWTu/RW7RQGs1/2Ab01mEK42bt9uTia8C
OhXLs/uFqLdupsnb9gxQOuMbstSsc0d+363UX4vhQNB/S4xkEJHnYhdLMY2Ooci/
vIFBOLRJSBgXHQKsFYItHg4M95RwhD0hPTFmTKEo9C/mXduPxxfHVVfNdml8l7MW
8vMVvSFOx8Az1SHlc2c41au12f5CNxBBaIpTiQT6/1m6YTyQ17gFNkQzsiz6etjR
nJL1K/9+QhC5pux1hV+pxm4sPBT1EDmG1+ogRnXaFUg1GytXcMBZt/p+50/xICud
WDQ0orufCSctbEKHFpvQ2pIWGk7LwX9lzk1fT3dNjazB+XWWINPbIDMMiNGTWH+K
mccakAtLjvc78LuFPvnPUgW2YFRK+tyuS4dr/VZmtmfFO8Jhz1XhKsVEa42sXbU7
09zRTl08NdVWU9exRLMA6pjnzWG8GnOrhaBQNXZp9zGdq3jDPLYZSwDdCPD1lvV5
+FbSWR5BCiUoIcNRzSi+NMqN/TUFzF6wbFh0VwLc+2sDwEo6+LRlOc1MPaF/WayT
YMRPMzcvPUcMuOzCBv77BqxSuMMLtxkjmQ5SK5+Hc5aMH1sig4hD4O/JNq+ShDPW
/6Edrr0XDsmN5+d+LXm5oQugFsclE+d8EtM3q5R2xS5TWE9nhNJzJfvWAXw9Dqa3
l5uV8IIY65cQ2kUb2mF8OxBbnHH/Zhei0T8EyroZkPzmBFH2TjeLkzP/i0O5FP/C
ThYunmXFwtOapBM9iieXip4YcMKl3oLIzEHEReSbhwIPFbr2SGppfSaU+GWxOM8c
xj+SvqTIg4dXW8w5Unny84Qrqje7/IwGhu3pI5ZI2d5gVZqjknE+D1X+qMREdkAG
UbGlMIcAfqEqNSgjaCZmsbTEP/L8lEOaqqrK1KDeEO1LgWaDi4e+JUPV1YsB3R3v
Ge1DaC8bTk1rDL6uZqjXGY4Y03UJuSumcgg2YKKcpT2JdPBES+cHjvA25CFDB2Bt
SxPVJqN6xCLQBx35ztjZKNRaoODICGFx4bVfPGzNe+pMXmOJq9vLRVHCZzOuwKho
5+vInYDvCA7Sn3IxRT/ciGxXMXKeCxpRNeg5lPtGQE5CVFmJEZb/kauVztZdcxDf
eO6fIv57M74C6cNqWQxjrFJYZFQISzyRrKQXq4t9CLySa0peMccoh/XrYZdycNuF
X1Sxz7TM6466M5eRsz0Qvcp9769WUPuMuv4EYlIF1PrWpoRa4tZkIgh0AAH7V3Bm
cdP+4mqGf3W71+NlvBDhFUWZ3DSUljZadtWdb5kc/oe41c5/Bylrzd3QIeMF5JdZ
l0ZAV4vwgegyyK6eMTEGZjaBhqHfc63ub3tfMjZ3AMw8flqQbN91lw/AYPEFnhAr
wicYKN8Yvw1UBZb5nvopEt4LX8KxsR/F2lTLw8JxE5g/dLPqFMg9XT8pda4ZrU9P
0L29NqhbeZOIL6+cgATvjJ/JOu40MG+fiQ46iPScyRvREjl7DUov3JVDG7pw42g0
ykPk0IorPjzFUC9hh/cOxXmBqZdOfxLhoPuYdkQRbM8Dhbj45fapIHBSogVDhhhh
VEjWaFuNUUqRIOa2wFnudCxmY5MAYnCkjUzNpQS1n7XvZ1hF7RA+han47FUuXTUC
FTHDAvSyn6HwNvoLXJS0hBTwatHeWPmfFNWEfTr6bxJvm6OTzxjYHldlsBZ36ie6
0J++jgnArDsa4RJ1WDbcNHUWvI8kkha6ukLX0e6aJ/QimMMt+7Y9O2OQMUM8hUoC
ZFeO7Gze4TC/9IYTZ0r8J6zlgZ6zqehkvTk0W8L5CEi3kssFJBSW26Ks7JZlwns/
EJIlinO4wZHnNcaEb7tw0QUhO3lxixugN83v0hLMsbfPR4zmksv4rnLnUC1jfCJ+
nIypsmHBAka0TstwBHfPjAQSgj+7LIS8Qsq3fj3ZRR1P/iJxqg2C8dt9KgUqLIz3
K81SofbHIee4AqYIAr67v87K3mMJaYRpF4Tu6T8dhtl2INRSJzJF45XJy8vGUnsn
ht+ZARG3dc7OfseCWY/wohEy45UjQgujoSXWxYAt1zO0yIxgQwEY7l4V0c+wXdXJ
XE/ANctM79mg2ivs/9NjqP7sloohn2zjXWXXX1I266hTw6Ed85Sn7D5AD2dR5RF6
guyCHeeKvDygkkMp6rmdHRQAa+xfCWsu3qzeHmXaqxU2pTdqr3IRmxD2ypRWAB7Q
eI0hyokejL2upblr5GXtU5PJsSDzOTcTjb8wb3Xb+T60fqMCyMBGNwqQJnNuu1xg
myxMMpUPgjjFolRfllkqsQ1pvXONwhrqEUn6uJBy9+Pa/QHQ2Xs764UBvrfJvT6b
8b+dUnlwa23otrMl20X0S9UCc3psv1ObOoWIAj2pV8mAckcctkxPKgAEVe7oeXsM
Qj77K+Hve+AUK4AdqSsHt58XdYJNb1IJLHvrKD5vn53hiCnSmjrYUQD0Xa6pc6Nk
jiyisCzDtrBw6bhtD4jV1EVkNKFCVlsMRob3VPjdD5ckSymeUe3oKitktHbzJMmJ
hF1Jb3lNuAbjXsf7ybbckvxaZMH5NnUPIq+gjXNQCD2upvIDfMrTTAiwRQ8jigLC
VjuAqmDk9+93b6lWYMgrr7mwG5ECslMNFczfoSOFS/MPIaKhqELgEMSFdAHGFPS7
cEqH+ZNcb8V2cKnplXOdNDTG/PVxMaSS0e9Xuothpp5VfSrwi2JauRWorardWbNY
L7ZIulBPoO0DJ7qT19oAQ8doCyAGYMi6QG1okN2yEIFCQI5WXeXGtaLWaAar3CoX
moKabeANovnxejCob9SByr67RN95hgNebCMNmKAOiFcjdQ/8YCfMDz4mGlxeY9gR
eY8F9nH7gjfQ49MdV2CZLutmAwZLsgOkXOlQRhK9VbRcQyDWKhu+OmSzA83wyqxW
EAuLMALUNcaBrsk0GGCiMgfcUqMY0pnMdK62Rdva+UKYO5MhDgq3yJ/87x2sfNbR
i8YqEarzhr5+7qtvGQX0dpQWRRvinocyX0dL6rShSs6GR3W7tyKNONA1c5qMH46T
3JrcNLMJUsuYTl2S5LI3dsjOw8kHxIPLu17hkdldEM7VCKp4+THE0hCF97lXWPcl
J0oiMWzKxK27DBTrVHBIVkM8LL9/gP4ccmtSY0wp5gDJUw3G+79Xn20Bii1weZUX
GWEsze8tR1MFeHLG4Ydt75EEKA8pvC/zQZmrsqdyqbRph+lsI2w0dxS/5XqNf4lf
L+vwKoyUee+9F0ePGtEtlZARNw4fkUoWWfqNsPvi+bCaLGc2Me1XGvi3wOngMMrd
Q6UqUZ9ZP7FFSYHrmoWkvDhKVLdGggy10bUvHWJf3vzKQQhCfhnUvMya7bPJEmMz
Em3dOpwGpzoYY19621mXq6809sWIGzIB3QD//RauILrTAqJop5R5eBqzLgRPiSje
koimKXI/SPjgDV9JPIPlrsnrAT16uyNWbeOUPynFgj0Gwn8dnyWCmgImdkyq9OwP
kFfWX8aBh+MEqJOrf4x9bLxzp0//sZBXihrBumV3ts25hw8EU/idscN3p5QZXqlw
8p0QMI863yrwRFB+R5R2p2mLDIzeFY4/zba2aVU10gy5CdPCef031Gop3KWV9VZL
ZpChobHsDdm+o1PBNtUyy3Wee9I/KkvEyUMrAgRQ7AfDMbDbnEMmO/RJFqC9Y44x
aGWY/rThQYifPl5UEDXwRkRj/SYK5OImR18pE1pABwkwWbwTLwqnNtnEfD9JPsaA
ZhqbIVppsXYQBds9P6YteJNsoFZxU31qWYcoAY1olYPZ8mPfp4YqOIXwTBYAspIe
B5cl+haWOeNbrtPkGy7PTS7dpCmB/XWGQnCIUIlTfEBm4PyNWIb/V3LEBYV/Sxpv
eEjkLxPwX80STExiTtDYJAKw5QgayRIu1eK7hSVh3ZFlBgwziZSaDRKtbP/fTV95
9GXejQ8sl2NuscDZ0snAQKjLA0hkhI+WSbz/vb6scHxaVqJuVDnPwa257JUBA2kH
ZPARVT6joDWuaVCy+UDIGWimjCs0GSFUQEfLJOTMp9M2K8NBQ7ZGmUItwu/fijhK
Po5VZoulsqUldRMwDK7t7yzPqgrWRKAHAQSzGBKJzlYDAhOgG9Z9dKccMXrk9z0P
UmiHI67ZCzfMI8vlvesY3z+w9Gw4u/qIxB5i9Mrrs09j0A2SyXzLl2stIyTH62VN
ElFHw2BkPUwa+4Xw8JuAUTwh9v0xsCW10um0tvXl6HHDmPNAdheUIGJyAyYj6hIu
OjALbu+SGXRQfHQxjcmRDnuDFyr3Pt9Up8Ec2CB5XYNmC3jfOR4vJO3f71V3dSm7
aWYfJrhdoMPskwAOI7628hQ2kEkPeqxR06QPK8g2OCbcA8m5hVwIb9ZPMXXDjsAn
ZKxkqZ1ipADV5smoO1xTVhVK1+qUY9kBUjflRSzxA2UWKz9+8jbMPlBS3MmVTonm
xu8oyGeDqWjYpwOusnPZOxmqDgpWZF+FdjJ4XhTzITXof7k7h337PAMq79pHJqLL
onEVL+3z98297QkMnqQom+S8igsOyZz9SRs4Gs1yFRHxS/GYGWzax+XezkjjDit/
ECQSuZErw8ZL5luItT27JTv8N+i6uxQQupp/ltoGvOl07wjW2HNR6nVq8xyNjRcX
q+mvinuBzOi9P9JyR/jWSju3aEb7hHWzwdBJWgAhjzdKy9TRsDKzYRkhXVqY+iH3
SrYL3FnImiVcK9/bai0pUZDwp88g6sNB3GYoTtTQLTAO7C1VoALV4NApDKMS1vnL
ceW0AQ/nK5mr5JlcGcbPDN5nH0W/Fab3SR/dwNrlxoRY1yGGB76fN6ksINofU45T
k4ygFoNpgcUiQkviiPS0HdGOFrPWJYnQtFQQCULYK2082kg+BVH3tCcfxqsJ0yB+
G1JdRB3d1ygJV5IHMnMJuba1Ni353JKyTkoH0m11xxpYAR9LG3INzLss58q/dI1l
l3Kl+sp9mCi6+5AayS1MCssyuVB/HNCYWqByuNkrw3f3FN8/TvgMooli5yqf0WKk
u4DmeIlS210lCMaIztbB5A330OPW3n9fGvyNq9XCxC6bZ9nxuBtWTmj9u0KGtE7c
VvEalrqmQvRSCo7bv2NIxV0e9LwypYSIL0k1YcwouNZtR2ElGJPwq6DrZ/RK9qhl
cF77Kkh+JD2I+x+Rk+3VSamnQ5wC0Hlw2YeItMwwp+5ANB/WUi1VKiIfPUlbshBr
GB7UpTQqQBEDA9VoumFEYWoRWxRgMzlK3sS7+LJ3AzLQRf1FjWCLlHlAdY+O+fs6
Yu1t97/gcFNaP4IwWEJ7rqOD2B2FJ1gHQ2lI4HU1NhlU9GpcOrZYZjEmhllDcGCT
pbmsofWmBZeW+3gCxauyq4XYXxn/iNgm2hXJu3Mx1Q0WMHP3OUjThbhV3MMZDPrd
GhCtfycUmGBVmdDKwWtKJWTAaphbtuRARUKihhJHgC6/InHWkykYl7RdLkKFjMxr
voJcJbTLGLpaUchkkMRosPze5z/OCI8KHQ3omqrZP2NefnHPUOR3M7bN+/sgnbFl
zxzCIDzifietiO5Ww9ocdvdwkBguA+Rc0s6bd9sFWrULGNd017bQDYtyFeDLIZiI
vioLu9rFfOz1dXIjuO3tz5bJiAQonajMzNM6Mrn+Fe3KfZtTnmurlo6eqkrmoGHD
hzv69hsWlqR9K86tutlwis+VJkjCs0m4xHFyMGOUJ4TnTi5uneVroMGT3CSXe6kq
08RdMfrqKaziChj69ZK8XYbul7cnGeUQg3QH+1QUErtfv815FaIapD5ZUIAdX6n1
4tDD7ptlyQCwOo/MCqP7BKmxZerGDF63FwnKfwEwgrMFFEVJ6CQxNPJpxGSyBZ3E
wCiXMSJ6ewSfEJpFSu0lCq5QAZ++7dMhpXhpiNuhacwoC5F0EjZjDIL4+o17R64n
wVdbVH2B+S/bFdos2bJQoAHltXMcgNvTVTjOrbisvWp9N13tK16qR8Wa4hfeO7Cl
HjdF+yq1KBPtU3ICXJykxwERgQbPXL3syWVFe5WA1l567r9zfQ37Wv2NHXNp5Lor
8V+MAIq4bkdbi09U2rrs8PMgjYMKUGier09vIqUGHFyN34Q0VR/AYk5WuWTi5+Jx
k6RZ4QHNotxZ20YXHJgvWzuu0S5goCTkXfvG2eSyXwdSQwRRu69i5MKUz7GQxuwA
/gawlLMGLqGqyoOsur5F+cPnnVe1sTu7uLc+ansF2jkxQzMSUd/cxnDwdUQhAARC
yA/jXjKjlBpf8fe2YMS2BKy4FTVnzfo/5v1+a4N1L+Gb7OOB0tiwLrkEMqt4O65H
6uG6N84VD097+b4ecw9dPpwziFm/S/o6OMoA26baNnFNuvu93nZlqgelZqY8y1NV
1QdWsJRv955rd4LbR5p4L1iy2Iw7eRDWsmovEtRnddWnJ6sQMbGqe6hm2P34n3Rw
4CSrPG7tAR4UTm11N+sRHUh8tAZz+J0oDgsx5nS3u7ViXMQyZls5P/D/nYa3z7AF
FvFAgL4INrROiXSPLktUrMPZiWPMeR1v1iFy8kEFlVFhHKXjzckuPtA4SW+nBlPB
nG/fkynaromypiA+4E93GDhx+6FlPlHmWeW4fzHmEvBpJ2ar3IRrRNL63LLfgCQa
HUcdurdVpICKfQELnaZYw68u3hjYGuwk2D0dV3wz5ajKZ2cMeR2iYawBHmHQdRMV
9wGoK3aDUGoEcD0/t8/YZuThz4yuAS246X4+gcxwTyMS4TyHhtqueM3Ac8+7ZTgF
ipAzzySBu2B/o5oIgtEcL0fVIYZSuSrv1yaAPYl7XZ0pI5P0PrswCYGyh1Z1jAuY
hsexTGJdO0s8nssm099O/ENsjxyIZaFXBX7ts4Q4JYf1ZTLtu6IaWqc5ZlPlWcwH
5gbmLM5HsC9UyTtmoJc3Met2Buu/dhyzWITWnlLgsF1qCn8pk31ljCdotBQyx/Vg
vByNYLLVcHe5Ypy6+N5Zfbw038xyd3WZAaccZnqDy/5K2Yt3EW9NFi2zoZPmO4eu
/6vsBTlyG/3XeeBS4ofsJY71KH7yXLhsQLVQFPahht41tgVxa13CTJ7XxrUcLd5e
5IHjblPefpFmxiR9dRI/YXejFhkU8aQ3vyeHV6BkU+ay1VFlSbmoJn/BQPypUcxh
/zNiS+LEvt2RTrx9Fx5jOpVQ/Ch/BDDsZFqQStu2soO9X3ODTpO6/4J/gyh+QWUe
/ledbzqs26J/xpeg8gtOLt6+YFI7VshogzbmrInanCUaF5pnvXInQImHLKWA02Os
MiemZWMqCz36tS+XfgmlDRzWcHG0RA9eNcaM013qQ8omNivugSzW25Bsj1vRJjjx
1dZaijqWgNROQ5A2iF5Sf1yezYY54EZ+aGUv3XLoo8mk3zDgrZhLM9NUgI25yN8R
PbmI4I2v3oETXHYN9eHL2wd73JRDgsAfMDAbYVlz/m9PJgDLswgiVqpeAX8SnPQk
SgREdmtp3BUSn/xQPBDoLsRDk9Xnt/x7sVxBIOlJ7A6IAe/QG29aDoi1KJ0QroM9
1o6qjV08A8Rg/Lme1DNo4KkV/Cc1NBwGYZ1d80keSZBL8oguNZ5+cFae6IuuHEnR
O8xqi+4++xhKsePUaplJN5qG2/k5l2l+j6Jbkqsr2MPNwy7pr/mAOKn1x8wWd3wL
m9OzcMxD5v1rZfA3M+SDF27wScnPb9AhC2M2HkxTpI5N+GSqZevnqv3iRxpqPuBP
mo8cF6Dx42Ln3G1W7b4TOjTI/hTHY3CADyBOvOrzOObrM5twQnK2DjVqVJZFqgtF
+uHLK+ChUMAKY+UaLsWncutvqNXCIP7nJoAKKudY9LzIGDns5E5+fCKUP505iRK2
XKnW1OZ5E7soR/CKRePA4kkTSbhal1yyBWE0lbMgD9NHbBPs02diEeLb57qrr3z5
+92yE1eO1qiDCkmLKXKsw5r27DZwVexM5tJdSTJLEDHsLfNhtxIB3e3yEB+YdixJ
w3wrsUJWqoGJVabXEl39PzeYpT4XtB2akrWoCng0SAtfBlW2fnk28cWOrs3jlx8y
aqz366InobnkVbKDAJcqmN2TfZYFU8BjdXZZL3RbXwa90OSr0qp0L+7m5AQT1gvd
v2+h4PbNhY2Sxsm3gKQ/z3C3SymaoUHXFvXk5QGlJ7poK+45Y9YibWMycWoOfLDl
G4vkBfXp5TLP3BEsgT/My/tgw8ra9E2qK6PvLwiNlsBa97flAuMZw5DwdLNi4lsi
O78UY6yFYNTAQvBmxijPrDcrgjjDUAQY0gBvF42d8NjRU5qewRpSw630qlk9k5+d
FXMGBmDiyzh+GCX5BKYMf1I7Tlm5qvic1HFrWGvpoOvKSkZHgZ4SuJ7zVoPMm02H
r/gpTa4uwoUsb24Ek/1Ae4DijVbZfSw8/5I5ibaz8fgs5nZ2hyI3b3eIjw+0Nd3R
+XYH9ofmyZwlv0OhQf2lG7t7wq1dpON/6DmcUaTV2oBxmnkwbB00SzKrZhpMAbQ2
yg8D3dKY4gLjK9DfwSdL33UGFidrhG0CvNTCppIfzlvzfsXRGEty7R/CRx3b6/6v
TD8RbvhEzRUTxZdeoEopLKIF9DeQlLd3IFfD3ZYZwvuPvHgny6jpA9cEeoe+SlY9
PNxWXTDMQDGhb5AudMfDL0c3j1earASBhSj1ZXO8f6vbCRoWDfGQnkKRVkPg3ulD
214XXbuqOvD+61GPHM+MifoyLWwW8v15p68LFEm1iIcOYnwYbrpssh52uLXfnFA4
G4QfT9me3wA6hDeaxz5nFRGdhQXKOJijAtTcePFvESsiYRYduLzJTghPye3ppZpc
5FHnxGtNp727yyg7DUrcsphKRwl5SGT6XUeRYS9D+I6o/MNOrNNKzJ0kmAeXQYVm
NYkhwzAPCjdxj+rpQciFxjZYt8k9iaDfJOb41d4KPb4EMya9K/O45Ng9i4gDwX2h
Oj3prfOzmC67xEriMDumfN3ZPdF8zSS0mwUTpG5NPg5TkQtSbM+wh01SJy0kkR13
g5DEiHkynNGbKjIphZS8LQj58pXZL0JNwS9FoWL6qhf1AMVnq9yXN7/xW5Rm98Qo
TLpKi3BwPcbYEGch71CnMTZIOF8QUdwshPKFPGnBGSbFmYwaauRYBOVk6AIE2j6P
gwUwCcsyBQD97BQDXZ+QFyF+828TkmI08QC03Y0wqxVHyzzvvta6A9s3dVukEcCk
lzlKAPqUoZYTh1i7WRgBrKBcSRrVJ+fMv5eMpzcidp+0DoA57a596q5J08M6AmPK
Iqn9YtsXTiR6IrZnhaadpBnDFHbnhkghi9a6b5LtyYv8hQ3NTiVJl0X8WxrmD760
WM7nc9RP+KOthBxiblXL0F4ih2qoXesfyIEa+zN/oNtfX60oCvFFWVKqwzpmS0Ml
bOooXNu86gJS5lB2NntvGsq56n7cS74cOutK7lpJ7f607gmwZJMse0TQtklxm73D
LgAp3Zf0DC1qXOAE/7RRnKGYzL0+OzFl9qggqM+qNQDDUdcF1c6wTAEJr2AqnoFY
p1cNcJqlycUyHELKxucmCBAUKUyCnoPlGRMqaceml6ucu6yViugQ1/NziQQJgTux
20t/nSi9bYUSTcwdILyY8Aw/GrPm8q+bELRMtFoqYDnkcCIY1gZ72yM5wICf3kjV
AGQnOXMHj/ggIltCMhoWd+kBa8Az6h99++olnuaX+2XhFvuKqCkLj8vZWaKjdpb1
IPHglKRnIgtmjD/O7v49cJ5TacJKM7FHg3uZ792C1eFSHikS1wBup7YnCOPiYeaP
aiB14avrJ0D12z4RIifJ46KRfo1TZ93MsqAjmQ/VH7QJ56B1gqmeD2NhnsUiENZv
ULu86jXyb6JnCETS6GrUKaVWDI7rABr060+6V+oqwFLAlYjsFvqtkzTy2VFCVq6v
VdoH5V10LTWDLuh7y9ullZNZpPRDkUz1elhYfvj24WheAvFMQxRVpKAGZjIAi6C9
U9evBe3Sf0qN1sz4fNiYte84Cl18bx21N7r+oPLrxV9tp8OkDzR7TUA7PvlYuvZR
8w35Eh2qyEBMcmSuXU52reGDYNLbbvdxVtQx+C2Gz5vVi8oXM7os6egV8ajDJC5F
h0HM47WALAP/6g6WKjIshJ8StXNv+PAgz5/DljThbwSMjFAl1Mgu68dqKZKXrE73
feBZ1A4gRPl7MBXHGwEWL2ZxlHWARAYhU/brUOeNQydqj1hr9oZanf50IkgfTi75
tHohpHpB9aT57ZQqcotvVDu5inu0M8IgQUs+dVfbQx4qS+rbC9GlaVrWVyUrZxw5
ktKPQtUqhzRTEsAkc5wg896vqy70dneRTgQ3pQM+qhoMaIHsqREJe2KqFP25E6GB
RzDeVpguXBzalXTWIMV6EObKl//Cb8VunGCGixlDobWMzyveRQHTXOjpbMPgu/mq
FxDpUckhafpTRLkt0+u+tHuZHqFaQteuOr0vSdPyqLAAb6Nwq29CQUth0YJPcUdE
gSswhTHTJrsnEKaY5zN+A57/A6cDjLa2S1gLucIT3HBAXKb5h0OI7gpDSKTAXHhz
bFN8z6INlCulnOa0TjgUsQo0JbVVv+z3XrATHlRFT9/BtySv8aS0gf99p2OlKi86
wuxgHCc25bYN5nx1FbemA2LCox80Us7rejU7elbpT0ucT4X3a9E5ZCvvTKkYKigL
DaXHB7+ONNezX4HoUILRiJz+GwHQWJ8yuxZJbhhYUcim8cAK2/jWKfCJr8bFuQMW
MaIijJQwHB6oGSlQ7j6YYkdZKv2ahGKmd7YIxfCg+OlEgzPmUCeZ7kRjrEAVIivN
vt9olK0VqPfRBkhSIz8ZLK3MMsTMAx2KdyuAYXaw61GixFGvEAdPvVRvJ9lXWR7k
gDPvNKCfjUp0rqn0d8Xmfpp0thf2RgOTojhZTAa9zOxrhCXbTT/fzh4c4zktE3Ll
xc8K1+FWafP2sWgDtdDheR/dngUvnfsdClbSAhH9TaBU94zhJYhL7rR3b5HAzk5l
bS+IJ7hGel5UzG/4HlHbNa6Nz/6ZhZrXAeuKMA6vcRA8umIemucQ3UH91T8r5/Qv
vdW/uSpUhFdidYVyjJ9gk5281JzwvtyEfvXFwb5/9VzMbuBsp0aDxL7T2THDxQMe
2eULz/CfdLoBNBQZ42TX481Q48HZ/ZbufFgL3iDgbawRjiMwjy+B1cW6T7spEzAL
P9ix8LNz+9lWJwW4xu5Nmg+8Tou4vL9kGEPNMDHLJcqFjSdUxiGdJtnKnFQJh78/
6O73ATwx+fAll+QiohHujnNvbP+Iu3VHUaKjPXjqgPkRyM/T+tzK1VeCWl1zmMOh
meN0pxmLWHmHWcSzkGRQkZK85Fi2OwS45LuXPWMcGQAUEbGaQgiLjThMeF4OgRl9
evnFFgJOevkJwYThtP/uYqisXdE9oBqWAyus1CWgN+wkvSRLbSxKF4w4IF0Fm51Z
1o/ElaHpeVGCB5BwDFE5q/wHlwDK4nmzaL4lQKBy/2k7vCd8GXFtl0Ln8MpSdpUr
RiAIjeomLMn9L122c7tVWdGQ+bLs9t2pv4yYVlffasVjHJjHt3XiuBZo8vckIHD6
UnL1B2FIgJZmaMcHuXlVwoG5/XicvAPexYYl4iQ1TKZlnamXDd/5xUuXEmEN1EfT
b3PPXYYr1+zf307HRApFLn5xb7vwor9XS8U/GoXq2CqSpldLggudhuaLosnmP3q2
xMK6DD+9on+nDp1ROdYOQjQp9qoq7CigvihAcj95FtvveUCVuAVbusg/HiXGSGwD
n8sRQ2YdfLjNzz/ShzNcRiWFhDOSjd4N+NdcybusLHiKiDXy6pN+lHZhLMlZYb8V
YLMOo0oFGOv7TWRL3L8NhtGpRBhjXdbAHJXFIVFUPcPnGse31ZCYdiuRNxdGkGvf
kMeidjvXVWhGQyyuOJ4AaDcd9OeGLSrjyLJ3Gs1PVmG5Oi+WrZyqZCrIEtVPd1dd
Ynn1mOe8C6bADH/2TnVC5QesAw1V4xSq2lgymzrdMPLFNnaYb8dwovyHynumEfZi
gLldJVSZ9sXon57yjgKWXV/A0lGSEfdvjaBi8YQq6ls4/jrWPFlnhbGgu/vGlFo0
4QBjQ1aXkUjHGgQpDZpAZnRJzZ00o5CP1iCEohLl5OJIaYLrFgDaytNvIVfRPQyr
gANgvl7/JvC1HeqaKh21ipoVLCa+Ge1G676WN21aYJnn5Ix3V8RW2t5h4cOWyYhj
oUPYcP4OfPyf8fYgZvJlDx+elfN4DI+qE5I4EQxbi0kfi8dv3XHxYDEMEGzzrfK5
zC6TRuPWipSPdi7veMHUocVMJnDRHH8I8f8eaXHJTXfzNoxGetFCyJVI4lGuOBdu
P5RxO7OQhPpYCeLLS+U8tvv7Djylqc0giEGESQ5gAHy1bFY8Oif94c5nsNaHZfRZ
bsWcFZw9zgXHdhVGJKinvPrK1/NJEHJrfIXGOX3WDbOt5cD7ImXk1y+xjtD4dorK
WGk6wLw4oySaiz2zkxIQe1Xs2qAdV9EGBHOPRSUQ5mVfGJLcSMXEP8hbyolgEKCt
Ke6gYZ3mzW8+ZPgPGKfsxWGccV7+veUx0nNzT8gb2LrwJ1M9wYIx/y/ZuwkHfjcp
/VwokliE51FsJ3m/pygidTfqFQB1YMb6cTWTQH6MVLAaB/Y845elUnkYpQPPdIYF
oezwv4Nrw50vxW05j6zvGNXMcFa7IV4q0Su50ZvN70hGNO+kyF/i3HlGjhp7hzWC
Ge/+DjUc9CjuNJJSzurhsVIKJfBB1/D5vCgpqNEkPNnksdEtRlEYDwHKP3fW8nak
Tup0Y3C/b1XlIaIvf6S3IKDycMAKcKJXJofwLulVE+DeuXdb7tKfmz80km93elge
KfYVN3IJlPpPk2nyMtTntFFhYZPt30tPby/H0AFLUllWqOuTlBgUZp4wF8UghBMl
FZfx+WK71QIrKRSa/2ToLeefLCjhdUuZch8o/MM1zeP/rZlC3aZGYqc2E8PmEeOr
Z1RNpq2qIGTToHyEfkVkAuaFaFeIvFCmSdQraJir6ifVmAoeNKG5uUYDM/4aDDqE
ZB7UWLezYAwhTnshSacEvWW2lu/CqJ/qNFBH3g4fsxhRSecfTJRBLz39FjltL/8H
k+DZ4kkapQQ0xOLGhyQHx+RdK5VzfMA/SJlMiosKpwQauEo7Vcq62tXNs52/m5m4
TVNt3m1UwX25z3Fx9uCKIk23v1BPw4zOEkEUlXD6TmLWHLY/jKgRmVPo2caXnvAH
HyrhLbKNOweZwwnmDXUsI3Ig9bEJnc8gJAIm0/umJTVEB4S3XOpe/7a7JAWAf/ho
mnj3rQEn3oZSWiBaKRKz7GgS/WmjcP8YmcOcW/cWq59kyc77isDx/lfNOCTdyOEl
BbwC92e2o5SvweHQ0dolINBzD52ciK7X5ZjCZEVTRLSyW0Eesw4wb8Hu4o1dUmB+
PGc5NQ/K2tO4NfxiBsVez0n5QFsgUyL3KHKvEkWlFl4VSTPxgjrh1Lv3g3vMtM7o
LkS7riL+qDM3Rp1MaT2pcPzBmHCUJyswUHnnGjG9ZLkv9Qpz/YgcrYjpG9Hq89Yt
VAAgocmEYGVGiQha6Crv8y56pWhcTDU0OOabW6Qb/fKE55jnOAGOx8PIFJkL7SEf
ZNFsVXhPYA1cbBBso+uEK/aizi3G9I/haZ2c7W5LYcX5joF5/cWkGhkPkdKfilTT
56nJ0E5qOrKdIQzDnK9VSeiM7po0GNks+EBqMy8G1PbEt4xt90D1Pkh5/+Bhk6zW
0sZvF3vDObS9fQ/RiCt34ia8zIFl8ZkTq0TqUyU+auGojD2upGn+l1oAXUCwhYrh
97++soGAFI1OmHmbvY/CExjD6AjEsbuMgMH95ao0QjUxQ+S3nKJOIoHaS9/mu4BU
6huU78Jz+8DXFf5zo/7twwDacWDVdV3HE0xmeIef5zdjnqBzzku7ezPwikk4FWtY
+AZE/QXsqUKCe8LFGW9QCKb+zHhBf+0gtgyvZzp7Z46+0b6frOuPWHllvApJLSj+
2tWMbakTbLA8QeJuZ72Hy2zSopH2zZKtwl7ILVGh4z46YVXQph1UfTYnk016htdW
ovaxRkX7viaO9IhZqHxPToEl6xHimYxiix9tt8z4MTNJGJ+p8GmRiyW/0J/W7u1D
S6PwB1dFZj8oIPeE3MOnOghmjayTvWUk3z+Hqi2fqYW0RFtQK7TNCUB6j/joSswN
tmMu5IA/hh0tuA8xeWBU3ybMeXX666XNGHCbm2f93offa7piDXGV1OPxoFGkQmY6
BciKuKqjZM3Q+W/IA+sy2T3YeESCbRmSkDKTdpS6T1JvPUPeh2pso2FE5mfkMMiQ
CWMQ5eVZtIw4tWNlNHTPS4XIF3Qo8WwJ7Qul7pWxXbV/uQsIMcrK5elfV8tNs//n
2BLd8hI1HowpUHTgl2ZhE6kSI36FqCzJRYbuDEVqfDhyvt8pwND3s9fmE86Plrwk
A/AppPP/hyK8rUhq8/2bRgH9YfMCwR4cn9VLglopoEQZDGAuukDUauTpPNI7H7mM
li1LJePB9At4sL7EaMxaAhEtasYyAu5ANyT/Uk66vyGUdQXdzBWKnquPE8KqpdS2
aOA0Vq1h0T2eZS+PacwSUsQ5WL0ScSWNCaUHmdO85gkgp8YJgC/jmfYpJZ89JRUc
4ISzK/b7AMvQA76OVegN9e3KpbT7L+MYxhUtwVuUlN3diO1hjV3v2mON8yXq4rC8
pCb0M7ZUBoO9vVvsoiQMcy/r4WD0d+2xiQmdp11FXxdS54a+9voC2se/PwwSwLPF
RaWL9v0Lonx8GJHBuFvypOFO+Ma3kwH2GP+TMj6xxaVUO2OP6HBicqAVmVemmeKE
9CWYrX9h7+xNwYA4xbZUwAjE3Oo4dJW45mNmw0lIBqQ3nccnwyz/0YaDBhsPT7rO
e+9v8NxPM7ye/takSwqihWesErvK6mPgucs7T/7EKvn1MFZism4Acpdm6ExGnYHZ
1Z5/jFGWlAxAI0QdAgfpPpd3GrIvGoEP9nxWyrqGvVVhowulbNNcU9K3PbDbEIcw
bJZ2mfxtqFEBGmPcMrfVECuC+Ps2HMRRLcHw0tpPUzRzd/oDi7/1sNenMpZZlvKl
7TuooTzZwG5UZjc1AkwbRmb2BZmn9zzfymjnmxAacG5Obpn8qfHKGxkwbkh75htd
HE2K/htD5jJY8NUSHrMbuJjv55fcqEtjdbtTKqvilMBVAPd1XB3ZJ4dBSVvVwsMy
erQ7NQ3UoMzZDcxb1tsOtIu4bXrynF38ObURql5PHeLklitfUI9PyUP1tcPd3wuV
I6hliBR4wxpk0plvHAbn37wEtL69eAMQ8lF6eUQmkQW8COrTcLpnudwBHqtJx0+L
8vklU00GpSN5C0eWNUcgF9EGTXAhR0Kx5luGxPZsK4apYmDdu/dnobQHLAOXDLnB
JTyKXGYDENalQBMv/6LwPDuhp1drMkFc5CBDpeYkkNfuQIVO4V2zQCNNOF4Hrv+A
G4kAK0+6ooe+ktwLzKhRVwk1NG53sWQ896JvxzN+GOz2rr8NSS1X+X3Y8FLzHY04
WcOADo4gVy0MYgR8iqneuQSsZYWzCzpgQrIrstP36eiaLwJi2vCaKCfnb7rgkvXE
pVnWZb1iQ+t5apZ3A3Nzd8R4wi6FLcPsmehWA93Ky3Tbf2Z2xGoqBHUDpx9WSr+a
Jl0ck/74rEjA8NWDG128HZJxm55PDxKzQHgj3Ouv0R9VxAts+AE/xHgzfZIvgt7r
IJJbynyXExYhkfasTTmqMuzS7fn1tw8cbkGPEKeUxOzhU9NGZbXHuQFp3lMXNLyZ
V0iDNBLOjj5uXAwFeIwS8ojUMUpcZ/mSs3xdXveQPbPyFBTeT6TUyxH5FWd0KFr0
zNtr3+OgNG4Jj2t3sjy7fl7l+vk968Ua3zoST6INYW7Vb9bZaLwrRxP+GeFa7Pyt
rmCq36INGIO8guUduNWg8qwFjvY+fBzy0B7MgcM0T41d5ouFf7bMcH1C3lUbrzBI
bWWu3MYQtqZOBESIIWj0CtB+nR28FjOHPlCMaRqVvsyFj0komt0rFOPh91se1w8y
46cuSAg4RMIRphlYpONCDS9ta4PlroJw5WarBbbZv3qp6pCIP/+9r+gFuf2I5x3a
rYPL1UhMwmT39qgSlkyUkVkgtugLXqzzzuwVaoefxWGQXiaa7HfOfb0xWkivdlnI
H0ktfjUPAnd/i+ouUjlsaxvK6pwPwiVOY5tWvc5DZv7x190gv4zGV0DcSTtwzrqr
qPk2T2xIBkt7rT6v8ZcrwD8rMT/AK5tfj8+hFnazGM5bEMBZy5D/Hbj5EhGMeI83
ajgoS6BA8uHlMEIhApNXbhTkXmStt7wYCNV2k/qiy4BVrZk37cPyDMpEVzHqFinS
HN9PAiUXRlvMRBFJtZcQZs1oWAaVxpz+6sY1zhLVDgCSNgyQiswpzhQ2WYmL6Z6E
J/yi6beL5kORjeiNCty9VovlvS+zP3+2XlBiJiIklyqo8zHMWhbuWVZ3QMzZ5uYn
B+S5L6BuHnPmM6LdlYr+CZkUtm2jnYp7aIoMnZ4lht11hTFJyynwVQ7oCbs2rQ4a
oCvLNiV3iTQj4J54uy92VpmpLCdrEXjWdIqNC1/wMfjvBq7vqZwz49fnCPz1DHhS
rwOIFufUDi62Ulq6D985ZGwlNYEhAPN71CwIrQtLPzt/zgkBmhqUUsPX+8CYdmU3
PK02nVEsiwqocwJnoRJWyYW7lMSL/OgAaT5SG4O1E6TGflGOt09pcF+RsU2vnbLV
yMCH8zTQFrpfANWWYiJTEjlNtvs4WF9vjejcLLVGHRowb5LP8weJ8DO6EeohouI9
fahqfQ+uiGd/Sl2JAm6fVInxtTb0ksE+HrRArTLIad5JTfN5nLw13tpHjRqT6xB2
NAAKYrPWmrqVd91SUFO2+bkj90ahgR06pHHFv1KPLRgBRF+hj7sMRzPB925R05pK
RyHcbw/+vZnmQCihICRdizrq+NFWlTGn1QEFuYWFPP7urejlYOUpgPGu3WWVaRtY
5Y5UcoWUebxXC13xvYB8/LEuPRqZO7BLSxyVZTAjjNIpfESQ2DXyh8fX4UfBEzbO
b6lI6tMUeRj9OK1HxMBjgBqNzXzIiDWB6G+xq07fYKtEOjTja7kb5jJyeE5QT5MA
4saQledmMyTmEOQjB1JqRl3iEf2PGm0cIkW37T8LqkUuW4CxFSH3KYyCWN2IC1dU
muqDPkF9UUGzGkDtDuzjdlJ82iu377vNmL7zMKSS6lFbn5aK6NZs0YWvCq0IuiNa
+7jC49Wll7sieAia/qm2qXwqwNdMMEiYz/ApJRM0l59BguPxyQjsWhEuIT82jIWH
x33zvFZvJyoFfoBguh9H9bFoBFGibznZfwE/Mw0HR7R8EPUBuqIFZm6NQaAflRZz
dgMjFpJVu76dTgpagCbC10PFPQg0C3IdRHI8EP8JMlM2E3C7mcbVOA53I8wcVtxh
YJ1FDcc2GCw0rIrmgg3jt7JHkea7GJTPUmDi4BUJrm6SdWtEigMSjU+knR5CUjR3
NLa0V3AWOVxID6HDFMTTn5y8Q9J2ZXQ9mGPCP5bvm8/ioPBn0PP4rSQZq3tvkBPp
AzLmLCN5+sEL/B2Bkg4inAJI7FZtNGYMYGmCnVSd6+JsBLB/GBw4VcDJcyrqG1DJ
NEfp555veSXITHXDQeY5/tgBLtJTFy+UQQjpRO/ZkAlvNZabpkK9zAfsfaQvKAJ5
vlFccAAO23OzlRsnxR85u+1BERPIpUILCis7PPPRYdc6qKlIw5NYgadHsa16gefH
cDUvxrJHuu405NJMmZUTRId8HAfQ4DbspfcN9FP2ch/f/YMAoFPmTsPDzX1keuR0
dr8KnXSgaiLrHtP3HapeTzTKjNfGXJQB+VXf7P9OxvZ+t1sD8FYBEI0JUiirTNPS
9ZGuGiKkAf5pr0cx9bRwjGu1ujbKD5VeVE117/K6sEOyN+eT8p99dIin8aqzb2gF
dqMhleoFrzJBFN4ql+1phH/cRGjUdGEPbp9BFBxOa25O7syfGXpZyxRhdUtaB9D9
wsiC00VB9bcnnoOUEZ622kATIm1+xjVWwMzjmZSklLjgRm0derwD/YU00vSNuxRx
hpE5pX4yLtH4lSb3YLNSfJic9hwo1kVsu+AyH6J//1Nsu5sV9n42mqqjOnrCqW60
WsTu/aTSDbi/dxT9rpWbTYlUnoKtv0/pU3YPcD0q1HtjaGBo4P6yw4NOdzGA5KJh
8wPlS2kayCzs0DbAwDMU2DNOm8gN+faSifqnRPp3kKh5wNQ69qHwEbshlaFgKtrL
psvoCrGg0mpbKc+dFYEcZeiSjfXOpYf+Kl1MpkbPym6y2w4WOLllp8inqT/7QwBk
1u2gt1E5rBEK6QOB3+OnO4UYvcPNsVJk/pqo5kiBzS1Mr2fB0Ly+FyUP9sAwRZrR
FcGvRA1wLt50oc+3QhJknRYzZM03g6F9UEZJeUGRRZp9pqpEOU/l8Cgto1RGIuf3
ODeD9ooDebYXjpxKcqO8wXwbrDiMW8XXlc2XEg9b+3F6Nr+JlrD0lcw4j7/bsjSM
KlcqE/vLE8jbb1EZLRLnG+vD6t04R8eTE6xOAhf+8G4b0rJY+5ierniZPZfo+fGi
42npEwYh+0caegiBZo/pCPvGeCQNnY+fJfhfYq4U0myDvRA7E0kJx0cwJgp6DY1v
ib1t8BMkMTy8eOetISXjBt3eb45KNX7eDxJsYaJAlMT8YgRieAz9NVNLvE7xlPX7
XCF8T9T1/ee1b1MsYb6udGQXM1Iu57Li4wEYF0bmBo6Lajg6MYj/2Qlrd7+rsUu5
CcgXOj5jbIoOhRo+A2eGBHNpqlhsZHrnAModoxIJTc+GhmTW8f/oOfBzkx2wspsY
m1heh+4nTyhCXZd6IXw9QVz8tCnWWt5tYuv8vAnMzeFVmgmGBFs6WzRBZ4ZOldx2
JTW9U49WrpS5BzEL/evBmWKh2X2+LFRZjB5z92hTXf5NPrurvS6pYB1EOFfyR5Xu
eDTM5RaCge4Xsqk3duK87oE6YOeDRb2wunygHHvy2cFW84ApR7KSgR9oNBc9U796
G/HAqIDV04nXnbqF9N1UV5EUhhOg+xL1WpQvEu0B/flSoH2FMu2XwCTeW8ljAevV
EQgZvyYu4G83nSLN6XIhgEiRVg/rE+Bpyy1jeceNw10WUDp0xHII7XnKxo5Gau6u
4TV2U8YT0J7oHZX7CeS8nb9ZsKvYrkY0Ui5t5McEoP2kZROz/UR2jL1mqsY5wRm7
7Duyut/BzieuTE780WpCch0VSpOm0yz2TL2ReWslfWMIES9Dmf9pEPpDIQzabv6A
Orn8m6WTq+C4DCRBTFemLiaOuW6e9vRmvi8PYet1YNGqwe6T/TKN9GBKpo3bODrS
1gSzlAF5UREPJ8vaWIvS1XOj0nroHH4fuiad5M+14zE6LZzxFpW0sRIdJ8FwcupY
LTLpcMmgCLuS7qXs/FVN92tUA3oxXZeBDlVGg0Sl0ZAWKp44G4FD+GYSrw0qS/Jp
/cST5b8GwEZlWlx/7e1vcPsgHuugkWql+g6+Jh2K1yQifcq38QMRlpwQl7vjY1dW
UMrhyv/a49/Mye8SAtiA4b1Y16ZXVlTNzdYLqROrckKHPFUsBDqWgCqyNqaYilLe
6ezy/tXlMs58xIyOBFcSiLnwOMiuhfT0LaaktLsapikTRvgCVBuYHRhFoGQb3T1c
CX2NJjsW0l8fLd3Od0kGUuU+CpwJVdbdhus5ibAYZtMLaroxeZcOs91gSDsyxa4D
uZu884APpdqj8WQdeJtK67BYan8BpQzM4xBdnO5Z2vs3+HekZDOb5ryGBmlO1+Rw
xIPCtwguT2R8VPFTB27huOm0+HQZSbR833NiA44sc3i2I7qyg0jG4uluXwGaypYP
dJPMPDGwEV6heCCrxn2OaPd2eMBTWTVUL3weLgxyzR/jXaoObPubvKLDx0RFhx9W
4feUjZraBNb26KvLxWcKQrXmGmP/AAFdMW1PXf6Cp/ifwMNWTwjOXORJp+to4dzG
l55hWJR40G51WOEXehrflJt6GiEMl1xtgC/3/tqbxUrOGMrdRupzEvD7/LhVUgFs
Ku7ZmAu4B5Na95yyYtMcu0CztmGwXvXIsPSnudxZbQnzK8xzWf6qRvFziebLOkwe
EVFrpoOIqu3N+eEOGe7VnCXE6GA3idIFHO0Ri8LN01Kcd/UhohAmA2f4asb0x8o7
b0vG4wkgJiSL1BfNyWXvnR4gPdREucIXaf/a5PSqdRpKTFi8Scq7aYqSS6rfCwhv
Q4DL1sVJI95HHxahGdCDINfEjBbtFYlu63HH6zwwsBcDlUFhblL+jY19hBSpFWMR
2IVVJKtI8I9OJHn8/nPiyUTYC+Rh1fZyelBavbiBnw+44HKnlqna1Q5oV6QJa6fV
s6thbX3LPx0C50SGM8bcaTBYCB+hyceX1WZeyblyf/zVlWMUnPNBlxiToleHsByX
PovdqkzBbmzpQDz4eGylwCje5h1pP5X3QIkg1g9dWqc8ij5XR/l4S3ty8gwCd4PI
nqsuC/ZA8IB4luUEVTOqaDH0mh3bLgHw4YEN8PMvmsJrbzhl7m12F28dg2JmR/pT
vL532KXEnwLZHHZue5pH00munNbsElzfwrkohsgoN4BTq8/Cgnlmg2fvqh/WsJ+a
lQEjE94N7x/Rbib0fKy+VpcKp+nEHH3RBbltkpbI3xYpkcM1MuwUbzy6SZsiGYBI
3DTGc04GpADkKWpI79wxaacEcOHmRNFOkb9MTVBWmxfS9mWjJVlETkxNAIOIQUo3
69RyYWYyNU7c5jMWO/sPFR84ENgxajRymbJwshOn9ZbSL7/ubF39N/fouZWS2KqE
zmn/iQ757eK4+lp7Y4d93nnRUTi12Dv2NYyNq7As+4hn0qTujfBzOM/34OvS+fc9
SPkRS2Hahp5oYGkMnMc+3twblTSKbp+Xg6DIeq2cACt15WM6wqph9kAaY/VgQWBv
r4sFfezrlMgYPy01QFVVaWp/4mnE13CZ/b395W+ZhxSLw++kv/gCv7p5C00aFP2j
wqU+2buTTxB5DPh74XJFWCGdmObOB+yfLV2p6dsf5k053StxB7azkPG9DABg/Vie
WNYvfaofc6bv0nnWE4JdeijBk3lLH76czDIodMhJsD6ojAfTIKEh3Z3opGj64o29
t1olXqiSHmrr3EQMD1CWFRnhY9GSHrnO9YpUduaI8uJceqaG98NQDM9w0a8jUpM5
91OBRsNLDKBHTf0Kq8ZXyfxjVhO3LwWfYEqi4DQeZyKURyix23m09L7azNOLJbni
gpU1DfqR7pP/+EK1bWRk3KhlHLbZ3ytpI9AFKuITBIT4kyM+aas7oB8ud45sM5vn
ahVF+b/kIzorRTks2CKiJT2bEqWI7/hI4GYQNivGLFUz5cexpNNXGOneUVjzPt3I
5uV8nvlxJyHVRnvIn/MO40xv1lszHcNW7RKD+DHl5UjBSo7zMKJ426egpS0EYZqz
yDWmwqWghRBGRd3p2cUopM3+2mlV6G2IdfE2H1+MJ75tvqskLd/SsKi1GFShqPMN
yCxbjGpd5JWw7v1Qhi6TIWSC3NCkZhIIQxgyYUewQLbQHafnWzTveYWyBd5TSVfa
qjtTFJmz8/AXMJWBXjp5qGEGCE+klF0UlojlG5g4i1j1KlNt64Hskz+5wD+DmDsf
0nmYqSEmb6PktRdG75dnavkRG9GhuYNwitmbigmf4L3Fp/SpJcl2Wqz8XpH01Hsy
X6OHu8kHliLZzX0gkSUIPa/JWpr1eir+C7X2tVbKgeU/K8YzwWSANy1OzogmCtYw
pSSmfVyIqAa6E/e62yttj8SAVTFgu5JZ2gz5ZAFQ0G9MrSzKQHDNHbXdKfJlqnLq
k/E0puH5EswOMc2z7/GmNl6ZWDoS+s+FBURq8zdaHX8A9WIqeRu53qbSw1YOMMLy
ArM3t07hR0XMtolD+6k9XkK6J/llJ7309EUkykAS7Bs9DI+U5enjIIIDsPlGw86g
IURKavXo+lcr2aNRySS/1xAWx26nnquSo/S+qyEH8fIAmJSds/H2PAVd5gKJsdfB
vuD6GszVqRcH8k4IHYRVWQJezRK+Z1NeGsENvg30s3dUzK+wCCdn+hK3aw09NHG5
O2DMp66cefMiBqGbpMW4Ni2fPOo4bMVNTZ/px6BTEEUlEpGWTeQreO7lBkNRNjgz
jkjxzm5k4aimyoVN/s0LOXSyfIpYHSxcIFrLGD/LKYwgNF+s4DccKxeg/OeUuJJP
a9avwP/ZOfRAED4SOnMX54SCLxWhSRi27hepX8NKHeWhZhRZf0Z+f+LKOTg43pQ5
QoMSN4J6Lt8qO2EAHZOZ0JMTDSRhfRA5PC2uDjaeeM6YTlJoLOiNfyQeiB79aZ/5
Y8i3/+YaW3zlsQA5aDWPIRwmoPVcGyt6gU6488wvgJ+iKRzvHJiuM2GMKz6hj91o
70+owN1RuLmhGfEzVcS1idgtjSnCwlo4OiGqrfdoR8KfeUoJ5pP/+47OOAzaCY4j
kgOEUB/Z9mdMfIFzh+OJVCBIXETqoYa/00itJoUubmSlA+1HVq3Ke1KAP2pQk9WP
axIrDskcduKju0jxbZF03LnmjnIXc0VNnto2MeeyGjBU92SQ05YlcBDGsk05xh0Y
9zEpfar7dcPAJ6YL3ZqBPZVoHidBFGV3P5A3xrjbfX4LqqgmZ66jFFhJ2IqeTqbd
eC30BZ+L9wfjIBMYF5DD1EXTH7XD/YJywDJZsNfiMb7HMQBpQLBUafibl71vv5RP
MpZ3qWkLIab0mqpO5pQqCa48gIExPlyQS80jbhPBCwl8vfSNzDXgYDJWXo/T+7Aa
To4pwmoXyXMI2HV/RnHP5omP+b38D1n+Z65sy6E4kR1/KXOVT/ZaOyqMGLaaAmw7
gom0t9nbeokY9uvGNDm+y17bZDeeComySnhnTckC6hI3IpFMURIPz9rVm5RBlpVa
2UwQVC0G8zGk5A4FtS2RMe04RCkRXEr7FQZN5hsbGUXeLHevSBx/62sF1fqVu4yn
1f7fPL/UMNapS+TC9bFD911uu5LaE1CleBwTv/5Q9IT6P8Sw523AssL9WKUKFNln
bTvvPFikYJbGzywYBfZc3mkTz6NevN/at16Vyr//DCPD1b2RYnLK+DEd3ip/y8dI
3oNJeOI9a6DaKUMfEJDCa4hDJQym6VT4cewVSlA7iIpMqZgkQLpjhfObjOZM0khV
PHU/Fm0jy2mkD5GHTS5wwZq408P4/BxCBEZ2YNM9wtIU/caeQXwomxR+tO8rx0VD
IQuOJmjreN2tJYPBo+5SRTNgj77800loFOysEHG6gAWTW7KaKA6/3TKra9S+r8Xx
rs3tOpWEj19HR8W2AQ/1WYSBI52rRgvmrAYnL7zhKbzDCHmWWa+WQU1m8X3kHGja
kAqF9A5U2Eg2sFxloW1Is7koappS+z5+auABoEuEhSkzxA0PyBhfLzkl2am5QSmN
MQt8EenOftrAu+/bLAb6i17Nl9zME+zL+DKnL7Lpv6hFndT42HfOKzSIf+2nKzyS
uoHQh0zn8qOeaAI86ukIZxtr0ICnP02GlBpMfxRftTiJWciKuvZg7VubRdfATJvc
bC9DbfGL+xAl+5O0JLA6ScXJ0KSNBtIjAStqyzCqKh/P1xqjp1Ih3Hj4LzDkypBQ
oMuaaJ8XGhiq0vzLvUMN14a0yJ512BAkEVjUNbWxAwWL/p+VJJZ+h3RHaS8z8rqg
/7JLfZYOaJtNCNF3NuLtBPMguyV0MuKomS59kH09N9N5oG6gfItrnyBLH4+ulBQx
iL5pmDUdaSZ4pg95wQCvVX1A1+OXFP9+eNrRD9XcPhiyRXSKcWN5AP1kX2gd7W18
MMjJBizvsdOMWdjMfkm5JAghgFtH94oSB6tgolNqA6KGHNwkEU2yByFY5t2K2GYK
dPfsIHQmRxl4vnJ4TrGwC0z0s7AUBorAaM9HOb26qo/TOrJDPWyMlIb80hhJuvQe
3KJzw+D1PlG1nZtG0tTjo4FOjcsPYxrq79tN8gBPX9bgmNn1uNgV4LZWzPjqqul3
apzzdskcxhvlps3XfkRVU4pnU7fJMs+AbDY/4AweSv0VDcW0Kai0H/OiJz96dGJ5
I9BIY1SuDesQNWqsIU7Q9oVumBcMzg4DrSpOTDbh8RoKd+IR5DRFG32Uh7ETUCGA
RoMhmH2zTvQ+7hVvuX5rleWjatqOUwcPTeEc5uNl5YjfYpF5JAlmrl6ckrnPptWp
lgxFiqKtjLaK7cDCeKOBX0vZs+1CUATFOpgA1c7GEeEp5IdhQRzKN37NVxWYxB7r
KXTLXjJZDA5b24tOsRKzZJ4hfg0wYVPHN+K8cIxKnptZKNX8oaMo01ve04c4eh+n
Ej5iuq5Z6SgpUjkdeFpcJAQtanZLjeAiovXEfj06xVJK+PDouFi7rJS1N23T6phB
1IGEhwLhG9oVlPu+S9eyp6dlog5VkDZQNrZmkiPSsKFuvy2+yGEkU4olHHCaR3eF
x0PSUkbTbToftQe4a/XPCQ+jXCRkpaH9Xr+qNh3TvShmUR2JfuyG1ucHpL/6azm5
CFrAkUDlTV/XmO6APOBoTWUC2iw22sonzb2TOVRgjfnW/ASStaGSKkaFWyxjKfuq
HrR6bQB62iPp74T3V0HI5J/5Nl2QII/RDQWD1l9Wp6TVbdujd2MeTCHCDq5h7PJA
VujuhorUV9NfcHcLDucbzuw1OkkSRcX/0PVY49syPyzkxrkywRE5fZcx+UF9kNM1
iCL47xLuUh/V6r+jXixXmoAbB+BL80QoGdurgiluuB6ph+T+9U+TI0K2vFOcHOB9
f13R1DU1SE9UwqLDxC46YrPq6CqWxY2LME3SZZ2XdqN+BnWtiMkOSRQQHgCFhVWR
jMCg6RV8+TDAR+cKQL30sW82rwFoVr7FI0eyzNMXtdU3XIOP+kN332iFG2suh9hH
2UPMNVaeAxMxrP+meoP0bZ8NsE4zq4fQGpzRvM0EZr/nxHVbD/s7al6tuxiAlGA1
xSLvFIt857byYRoi2mANfLcEsvMa3/IRwgwOwuhM1jB2vDjYQ3Tkg0va2Ac5QZ5G
m8BRMJ3o5YRN1kN+lOZmzGDnIiGUjqd1f0Lnctm69Egy3/vhZjJjnk1QpiGGEOUC
zjIU/1udpC9xajQJ9rnpTkza2vKMVjX6D6cIN9TRd0Td8fwXykdp6QxBCWW3Jhqs
qvaOGp17jaaBcxQM64VchVK1w/zcU9wt+KCHd1eO2SK+ok8le+puZliaGQnySc1a
FioFtX9vGR6r0qztq8CMRFTMJkBfpVPgk52LqqvKi4iVSA7UCqv5Od2aT5prhFjz
j/GJ8clDP03B2ajqL6UDaHQD/9QxOp748ytsnqA6EoFITujOaQPFmyJfs6sbosXJ
dKRh/IkWIvpln8qHgsPAcE8UFJILPcOmBpbAAxq0Wp0EcipIVf7Fgn2cOXkNxu2d
eo8qBr6IG+9I1uNUILDWvMFM0mtzWu6/IzDpqx0zuUlb3e0sWMRygDYgSr5x7T2n
xT/6786awhaK59xJcGHir4cSkkiJ9Bj2yhdtC7XgQxg+QUxpFYD2n7db02zO66/1
lT3S39rcxRn9G9J4XqmAYyfF9sk3LlSCgNaWFqtUegH0DZ+I6JoZ+O1gMlgR3ikM
dD0fWflwFy8HOy3wOE8cz3bM9t9JFexAhxmRie57vbsKG0chdn9c55ym49rR9Qdc
7cal3z7KDU2JlDu2kv8wPmasEQtyw4zi6NThRMe6WhLeL7L6r5MtmqbasdxmJ5BR
4uMzD0QBeSs36+iWrhb2t7pGwLios5FPe86u9iMtVppU64iIAk0LkUCEEPoVLAk1
IOREuaFHtgJRbaIGkkW3Ev6GCvF7wI2jR6/oyaRm25K6Zt0bwOT0RO3s1DGkScYp
/ePsJnRORph+jApPVbss/P9idrrUZwge++1VNOf+Q0F2hU2ybaYglCVF6zs0KsSp
R2T7wdBT0+5l/gyog3P2KHv+/Z22kBbJoiXK49YexfqY0nwb/huJwn85rAoLYZhK
Aqm6Q/ReHIRV8bnfkHRSwU4B1nB8v+92543Ufllcj1LJmni8lUlOWcPKIgAEzD0v
UPVLKX8Rpa/1u4tpnqlb1FUpC7yMRaGJlWAsxSC3d09EX0Ix6z5KGP5uO/YgzstU
MDFCP6OO5h7ol3o1WG28h/SQa/SdtJEEnnfhXRhxvVLEzG26mtBxOhRa1CBYVSzn
JeNBX2Fod91lIJgufcXGzNP93ujnzs+LCao71weHwk2yw1GvJtELkjwKeYcJhRmc
94uZKBMA0Y5R5jzovT+YN9lxyo9itTYn6Tk0FvacCC2RqtkCP8o8wXVyKCe4Hi/6
zJ3hICEpymNwcKixJ52sPYPb9poHCpK24+QMhOK2Gdb2zN3WL12ZNvxf/dD687Ro
tBK57ssB3vJjFlgXgrDTftqrzdoQxr4vsTuIy3T/f4lKBEkJjGazdiwBgm0nBDK+
ObGacOLrlOv7/NfvbJNSzZAIg5z+5VlwWWUqj8ERt4qspF7hvm9glMp4ljs1w8Im
S+4MiYn/s1NSw8Z+8V27qxJg3zeERPVGs/0dDez4hSFhhmoMhk8QRi1dBt8sP2lM
+ntXa3WFB8a7K3hddfQm9Wg4MMCeaJn4yKlCj/1tggzOyMHshpGlAYSPqYsyUC42
Z/+Wup3MQkvDKHRqG/ML5zyGB3N9bCvHf1vycoAjzwO9YpcFGJM/ogFCh6TwZrUy
zef/ERatNTOl6GE0kUZoVXhBxNvMjAef/+YSnkpZ5eX2ZHTmRpPUaq+2fqW5nni8
++YSlFJvo7sbIyt0UshLGLKH5w/0T65NXHri+gIPiL9RE3LNqh0mC+ka11oI6lp8
r2N42zukKU5ndyOeqpvzuINFv9IfNH5dPdPr72wK62CfG2c2/C2UmlaHxZ3TYFPH
hRgLSfpJqQ7bGB0WTA+2pZVixGpG58b58c3IO/iLV4CC+15WUAFWp/tPqJeA+BDD
IwFLXkMwgEZq+mgbkF6SabH2wt3gMpLzzVfF9+igA6Y9rKXYMguSgh5NgdtU2ZP1
X6GPs0kfOAOyyAMabR63MKYGPBNqad1L1cGnDVNMBD0/eOLmPzjbJzdAsOjWOPp1
az6u5ZBSCe0XXwBM9gfXq/99EjVB52taReLfpMy0iWfotO1aMrsu0qX3TFnOh9zU
U36xGvLsRO/biz2jDj//jl2Ucz5EkAO21DV3PQgUrz0Mw7xclVIP/ONcKh/aUqKL
AqCcJSCCyn8EnbbZLub7qUgvRkHbmz0MfQrzFRhcGiKNoeoIXnqIOg4Fd9HTla9n
ieURlOPknXpm62SKns07MWB8hWuuijqSVLdRbEzizyjrcrt6fP3XTavhnLSxQzo0
NJJWgU19HcquYS7So3Fgf48wj6TWKQlsosZd0erqHCvhsOzJick1JKlUb7yrN6Gh
dapNyHuWLUMk9uD+KJTKO+pCq/moMJ2uoPylqvgRtYQHrjb7AnFc1dc5/eX2mRQ/
71rEn8ns0Vdmism9iRL00yuqHkoj7Sl+wTFUIa8VKLEAATTZkzDKuFHIxQ7v50qW
q7C/wjvQjb+KCLWKkd/m4sx9xEzQJSr7bA51x8TLctO1wPRVlWGDZr7bn1xH55Rp
6qM7YeEwx5ro48pK1E9tYQtGYMVEsdDpIq891u+WQfGAZ7gdZRERWOiDjvJc8oU3
iXbVbX9RXY6f7iJF6rmV+XJVxD2nRyfHMaZKu30dxjyHyGg4o9p32q/oLa9v9wK2
O9/OP8lMN4XiPgnnrTH7Cb5jsBeXQI3+WJ815EcdP4B2q8QV7Uif0uA2Jei1JxcK
D+PE5i/p+KiE3wVxnelxx5XOV8slHc4bxCF2NBvGu8DUumek0rqxdcyV1dmwwqku
a7A6Ru0EfmxWOUI6Hm6flnUJOszyfngdJCi+e6NergIVGeBYz3e3XUMk01TZ09Fn
JDkqNeximAIlzA1tDrChUSTWpokmD4oOBfAAksuqLgJ827UwivES6ACY7M/P85RL
YRLu13CVekXiuLG4PMeClzi8JBHRezht1jcbi/CzctAbMYbQnx1WvjTE+KjaFyX6
UmLOPaitAguFpWdkAWLnruRoo2DVzlBOJ3Kz3StD1M5GhjNM/SQoiHNg7DHsQAyx
sWeh+8k9y9HoMOlZFcqyihxDoc4iZ06qPFWX/3XfWlM0IBsF6xu921ltuqBwqud9
TmkD/ORVIUM/LpLt5fP8pzZIeUslp4fx3b9xTFqW704SlCFRp3C2gBIoqOxXhv6U
IC+q4RTPs9q2zPWl1fktvf+MIy8OhahgIUyg3ap1TV3ZcoaLsAXnXDH2W3OvhR1r
mJpPCJBV0CTGFdGhzX54XsJd6WxpSyIe5koKlfjoJNQbfrsj0SxOxFJq0afH2TWn
7mxIvsCVhZ4ejM9fS6Qkh09R/tulL5cidwbWwSTJYkSCC5tDO8ZceAdPPnySjLHG
/IS8CUpOSeZdg+P4XyW0H2h07NVx4SsuYNFUH5SlUXTDdUHZTqBHHnYpxxG5qS1Q
Bn/Ns5S9vzDg/Zylggqe70Ek3BOtbVaNIksKazPi3YlMYfkbUIp0+eX4nIISm+DK
qgX67ZuWcLzdFaQaqlgfA85UTmXdfY2aaFaJG+DpeIHjtW2zW9sY6Ga6YR1DnISl
dWbVSimrO0TfnKF6dLpbtyMFVN51wOdICuVR8kGYOztELMXtsjsaDySpB1zpAUgb
nStRtQBOfNYpOMPdxuA/7hlkLjPP/o8rpEk1hGdqN/vb5WgwgABtd+j+GQ3dLtCl
HamF2XoTjOopyBg+w5piSemU1naBP3LKB7rXlEhcujkrrz6rUtF3eKmO8RRTCKG5
T4aAEOA7L7Ujsvgk4oLxR4mVCpa04WgA616AvAq0cC/Gu+rWtfVRd9GXsybS8dB3
8sAP5zpvOooG1v8gI3nZKs8altjHTyleQVSfKOhvVlbtfT7kMO7h1HBM3Q1FYTT0
tct1o14y2nkJZXr9/AY2XdtRIGFj3pmJgmxAwxhz8hoe1MH2sqzwlInF3O6d8leR
ELUmnF7hPv0wEiADbrZe1yKnpwzT98lMABLNCzkGhttt9j3LGVbEXOBLxUxTXUYn
giEZjCLGgmhqhAGK5s2/qEQ6NOLv+d3eLkWNdhKhxud7icr0d+oKUZE5+FpeYEL6
sXZEObX6jrtr3fg8QWIjrGIAg6ysR6G+VgY6cQHbFG1a0l3w43h63jAXQgpsD/Jq
aPS/zSvM/6FNa3c9cvdnEd7VjnCMPales4mnWNoyzXdtk8QZleZP9huiNS2Fs9I2
Rl3fVt8PtIPZ7OH6dG9CQgW4eX8bADI+EDWhBOUT7XugK5WvBwd+7iX0A7IJ4x24
WTHu5wyc9J5llbGWDVvNZOsCHJs2lm750rYzfPkiBnRvZ5I2WCO3CebKTT8s/Hgb
zJ7jkMWPs7rCHeXXCIlCGXaVwKTqAUWs9N1gDpG2iYJpkkgcBz7vQemM8IHds4uE
wbzh+LzwnqTKKmZ7L6am40Tb6BpdWNRcvHuv1CU6LIRQ2DyDKKiZsj+e+MUHA57H
G1KqwbNmzbc8mAGEEvqfKgHgNQwUvplrggAlQik7ZONyd/devkrEuUSSMchrWZJF
5pAWVrzk7LZL7wJbtrNCtS3rrN2w3arHqEz2wN6kxeKs/0d8VtBf24O0fcNlAjo6
aBoa3ZNkx5XdcvEHb9lPijBdz2f8Ua1acqNtWCoyV1iAuCscxLOwrm0iPjTWOYGS
/518w218U6QH+9pIIiqfkBXFdHO7Dj+oI8ktOUlpA5JYCPe6/4fCnDkroQHiEv7N
KsmTHGq5FVJgRFa2ndf2IfakDYhJWM7eyVOquNOxg/FnHLP1s1cxsTuQ8XtMWKQ4
Dfv8mQgf4Kw+jKvbJcYncTE2p50Anop9Uvu3IVa5oi8QCpPpvDS7fqZDh7BKQV2W
1WWyAFsiK1xbuBbUMK2pqfCIJwzOJErGgK5WJvZFgTXJKQKUR9exdVscXgu2Jslk
imZ+HKb8MnzNDGKx9KhDSdLaP1RQMFHXlSnoJdyap9cdnFxODaJeEQT7JxxaBgyE
D2UxkKzRLVj8BuqIMeqJZj3Ks1hlMUESRa6a5dJnkegEjoC+UWPXZG5N8wCzg02f
0E5Te0zwknNWtCxLJ+t+SSZDucN27YUpoLBUIci9MsdAGhU6woNBZqFkNsDYPWI8
VSVABGEoxy46YFScT/h+UaNCkhT49QEm00hcqiqxMgYBWxjNy2FOBbG/IvlO/rUc
XQfwQBWKvmv1YjKZong9MZ62nMRbYphz7ZdW8ap8cMkFgGvSRzySbQZSmzDvzLRy
yeD4cnKAebSgtmcSUKqWRuhg1BoBB02r9Jplj4BuxFSS6zlfYI6eypcb9cwmFT5M
Hq8b+WjHtdemaiJ7sgm4z5g4GOvVPrG1UFe+ou1Xb38z0Lu+JmkGRQC8rH//W19q
Q6co2pORMVkw2flZjgK0woSFyDpfihmlftRF+ZY07N/gB5jba/hO7YHhcIencHLW
nlSU/FJAsIBIcCt8YUTcMAKz59nnp8ys3T8SJQqNb/jWJfutlhgOvpOLeeVAudMq
Cs+CpxTFtSuIOeOEj9knMmjiz5GuGq0dTRZOUaGWVhspdBb15tvBC0okfGTAM+pi
Cc5/2ep0RpaTF7lfhguednK9zFwnFDQBbQRst0+oSxzZ6uMOj0gXzQdViah9tttj
1hwOshccATwjc1oOYfyB+eLk8KR7MyWgN5I4x3BBKcVxC2+ZUAXiOj0PROBkjzhc
ORZG8fnPPWMP2eXUhccA4goHFcPaQKvKx3Y3QnJIo73O7na6tO/difZbXH8cgOe3
o6AGIHkUj6WDv8dB/j21hGCCVWx+XXJ9IP9VTUEGT9IULpW1zIfuVMaoMK4RdIJE
od7iei1AJgzjPOBLe0rPwzfoCI7VEeeaorCRilEYg35/XHpphjk+35qaEPSLi9DR
OO6yfVmu7ikk3MqbBbmO3XCe0vFksMf0yKN5T2Ga9r/rOrQ5e6Tg1+rGT4gvEl1Z
gjIpVO7UrIBGz9cMom9CDl549fzFquoPPj1g4AcvqeGm3Qh9aiSAfulThUYMtaWC
Vl/4Abh6vCYxvRxLjreCdDxRR3i7Pr7utzQ63n2tjxdTcIpBenOOV1zg9t4zVcOd
vIagBOrMjqHuOMPg6IdF6L5uk0NyH9XHkQVBWNJxgxG3r0tmD6Lxr7dYuK8fCBiq
2YhGudh29iGMoBeXvm9Z6I9acVIquvufPNZqgQPHbMvr7p0ytIvy1BwX7kWt5tje
ja4ePNwirVlhOHvQymB+FiQYUNvZXfdZZ+E/sUY82pRZcYjPS1jyNBcutD9re9gk
2Dhdb1qmTZYRF0tM19a18WmOfNvJhV5n+UDulUDHUwfdJ+fTf0Q3JMqi7vEObU1A
Z+lmgNhQX0BuUxZTPHsFSq/mho56HbxFfYTFYkBvUZfzV55ztNMK6g04psQnS7Sv
LaS2npqJPVfCnRPGjbCSDGnYXD3pvBFJrJhiwJc8AVy+Jfg2MWKo3Bty9yZno/dV
m9Gb5URkU7yVmolDWzL7X4Juh/MOscroxdEIy6NznY+N780+6u69X2Q4mZ1MfHD4
ST4E8/87Ptssl4fK9R8miw69Ozg4UWsIR4EKZFvHAvsCDyeYjSOJsVDcpDE3cgr9
ggts64aFXZKYMeMaJcq/ikUlxH0cSK2eC2k2rsv1cYKtNdP6P6aNG10SWwkeXIln
zQz+auJTR6X8Jai7ka+PdW4bMTvW9XOLvNAnRa6Fet6TQcvgEK8sO9WQZ+JSGI6o
yFG9NwnSnk4e1Zq+MR8PtYlixRQD1U3mXDvtsC7raSGRnMUpz2qrHpYx9luRdINe
pMpb2X1YQa7oygBtHmURrZKwUTViU/x1PHDYnD631JghT5X8ir5zWMkujCahS/fk
ql0D7MaQSxAHipFgTWHa2AVpw6Po1d/lpD3mLfI82BPrGeMPka7mRXRJ5fnk5b1v
ZgBPSc3elKZNS8AeaX8Jx54VenltRtgiV0rYQeiuHjyCDLKmhFXzOjRNV0Zv3yOe
/Hegvz0UX1R27PIadudQvHM3cb5kSafcaQlT7mIX+J4XMK7uPzko65aiNNRcDIH8
U/oNAS1/lA+LFd9lJDN0Tbkjpc/chlpkRiPT37yb+13+hZw9rbWMc0iNk9fPAzd1
NEmK4m5iQ6pZk3cV/DLQ59jQurFH2QWLiUXu83sL1jqYwyqwdjmsap2SnQD04atQ
hHHGNXJuT6nV9qw8yQzwHI8kj41gmEPTEZJ2wsLgrC2hJ5lF3eDmH7DXbnFk0uYr
qd+N3xKkJZZG4r5+rWfzelafJ+2Yttjv18/3j9foZ7g0bgGf1ULQuBS+X+c7B8bv
aGZXIGQCwNrOKXW7GodP+1nZNrFykVvAzYUeNUiszeLbtOoTqBxpfC5fXyAOIw6c
YqaTfXKtXMkocH2zSLlhY8LJj+xOP/yRtRL9rhsqDFMCS9TUGZZ7+C1Rq49EQ6c9
ZRpHUCm3nDv/XCr9lRNHgd50gDIJxOLyt8Ciiqyn90MyhjhR5Vfu62nnhcYwfJvU
bPWc6C0wEhyYijfjZ/ELHetH5wrESfr7y2BpDO44Lx/LYuOEBW05dTHLYN3oYGgm
49xsmOXL1PwZljJ0g0k91CFPxXVZ5Nu7sfw9oYlhh85R8pbbo1+C0xEXQnjpg3yc
hMWrlEkOJkRD9FZXh6SmjLgVrf8c+6XfY4WlDO/HBD6h8wInsRZLq1qr4/oaEl04
qSZWZ1P8fu9XOwapsPVJVxaXPTmc41aLkit+gSnRteKljXD6KiYeV7T/BIIAF6ur
oe0kI+rUGHP8guOXeogSdoMqXE2S2nst4anoo07jtIqfrLnj62Qp3wBK8+SJUhho
HuS+ON2lwNlXannog38lew1tBJZyaC4l99QifhmALqhiVoZgTUzlMHRI0jUTl2FY
m2txrDFX210CiWnETPkkCgixTB+w/2FH0vHCIIUn4bHdwmAib3VViZqndsDjUeUR
fQD+MYrOGl9YJzCY3qiJUEa1escbFiBKe2DA3B2hdwZ07+z/9QlcdIkynGhM8dqP
033ERfHtUysVJPtB1oeVeSHMmveS/CTa/PA6bXQcaBNSPL9uSLN0TLOXbHqXqnxr
R5bq7iUSRViEPeCJ18Q9BvhlskK5LOfASOSXO5EGV3FXIV4yQ1b4VjTK7tUvDKsf
JM0WPrgFCrlNsg8yp0qqb/rHUDgWdUNVBcodU2xXMxhaYRXDJFnPOA/M3UWEWB+n
msoVKXmDv+1Bi3mTSGOw/aGOFDlPMBtpTlsLqYdfN17wJSRqci6uXY9buwL51zu9
vqqa0Dcs/M0IvrPulxszYnIADZ+DY5sxfznQMA062TegoG6OVUK6tldP9qXl26p5
4LZ9fi8wmr3lqKmHu9H3VTI6Oy8hGr7E4yyeOKWggMA6A8f75uckQHiIPrDrSE30
FnC8z0m3ZxoSgvDfwNMa8RPXw971FB9aI1dTyZzIqUB0qQAiObA8LPrKxcG/sQHT
szjGIYSxEevM+4pxk19hbVofjnCJf5nH06mthpP5LyFyEOm8OovA3K42b0ocOCmu
DPz+VnhhJPVxIUSeRR1C7h6qGTgZpuyTmA46BzxAMNJ4h661lgYQwAnZC7U6WUyd
YIpNDSU4kBlQ5ai+2smwTFFS2QYmIYHGv7kQHw8uobtOeM/5XVvlv24YMRtQ9cG8
AZ6AzSMEe+ZhQJoQU5TFyj9cVicYyJJgD1/dIAN2oLB8mscR1ZEOIiZp3aBnJiRZ
TIwsTlz76e6cR2e2ZFgD9rjYk9NXOhMgJU4HB9opAbICSSlxuTLg1kY84hLtZp6J
iT9FbECtO2+75EK46KvHBgUOLZZHVNhnO5S62PzK4GmoPqohyutuw6/cUnZ/zcW4
N3iwstDI9tRlOeZNAjvROYIS5fm7WTQ0uuARsvaxKRxbvHAWZlRXYPvdL9DnTe6H
Uvd7cFZJK48zV2GDNNh6O6x+wRUCNw/5GZXXbtbIJNXv5xwQ3t8PuKYiqrHUr873
4sfqKPcwfZZJ8/OKnYzZI3voQgpDUXIAR1yrdTk7D41aOztN9av2ydicf9H0fN18
zTMKS15b+0hVdbWMVGXkiU6C8c8eRMwqkHxvaIXOrS386N59TxCXRks1G8EUy/sD
JBk9oHz3e/No53h9E7rbeVluFny9UIgb6IrZ+x54VvX0H6YLpIbIF78I3FX4puhG
YlorDK26mLmwF/4Upn0vmwQ6vyTAwe40AdnyQ0g8srR/gl4Zbsm/xQhivokZjmC9
wHtoArI8ZyBqon7IdfjsEdHUvDZVAtrTiBvybPHppUlH/31fcyzVH1qtOtq+vEap
VuLMlDDk0IszSQ7i1oiUIy5KBd8n9WeEYBKYlBUKey2YonppRJNSoEEBbZ2wfqqX
E4GbO1MXBTboOehGUDdJ4mFI7YFP94jqxv+oj1asyGtj0q6v3mjRafq0VOhwRtd1
mKIEUhhjh8l5601zr+wKGCMil7Q5PGtXfAwOuQF/6frJixV+9h2TmvH7TuiffPrV
vnBzUlL84NDWNLYzb420DSlucSo4uFBRiZnULENhhys9SVJFp6reVE0nzaa83Qx8
Jm2ohKy2Zq3CGfbSXGd7bF21lPmAh+bAZyJk5I7w3GWFUM8INXdGcYw6ieNvY8Ub
uYp8qGPR4eA6fXbAeVGLtHUNJiFfNW26HGozKWd+LvKzEaOfz9JT2cPCymU4h19P
I5LzRMeyI4t/GM+5V0OGBCrJe84ZzkUwSmbnHeZwHu2O8f+1Xn9Ad4O4E09fYXQL
ANT+RDK9oDPUv2uXxgdAHOc6BVsZ7mmtGPVpgfGgEP6pRpNcwiqb7gXpPnWN9QzT
r/ABqd47N0wZBASSlC0hHnDkRKCuut8ccDZyjkpotQSputJpC43Mb4+KRLxEW6xk
gnFqTSUzlujC6918wjlz+9dk1OLLi3vXacHO4cnGHfKd9lLP9f8kNr9L47hlyPkX
Gm8dYoweHF6hgFOnpLYJ5N8mKqUW9c/tS6gKoTn/ND5T3dBW7LohwCMM+r0xogMK
yw0LMkstq9sDtqlBHBIHJdBwPSZczk/ZO+UNoy7vcjMPRb373KGuL1le+gBAjFVt
iMW3XyEaqsppfK/5f+X7j1oassV61Hrdh7EQ+RTuOORodUiWz2QRlFSy7TFnDn2b
+6PbDCnD83SZZWb55q6tlf7YgIAMveEozy11Fz7Pf3c5AMylWhw3BOO4bY8QqUri
Tmj8HKpLxEEF3TV+X39qGZ/8xmEVD3HtM9W11YanX2Uvrw9z7PHbVpCBlOWsB26x
HIWr2GlpLyPmSnvgz5HaXyWoPArj81OTcGzpwrTY/DcETrS1gNbv88Lr6poY/lBh
acGKXoQ6mU7mWzXDv+Hc02WSK+pjRGeZx/E3CWRd4p2UPIGSL1wbw2vuqXUj8sro
LXZ3VgTSTmQdWUAj+/P9VYQ7+f5MRfhbIussntCbRoeuw+TQ8hQBGgPzj+SI2RzS
qrduVsUCeJt5Aj+iu/yDNoWwUUU8Xa8BfmDagw41KJU9BkAYFlPqKsLHwTTHuQR4
3ZW4ekorOQTXZ5rhZn0ag3zVGYqTUaMfKfpm7wnz+6vOt0/dBkNJ+/+tWQep3QOA
WEgayeNr1Cjf5hwAcR2cTHArtRF/YXnNbzfYaE1bXdan5yysN2gz5DjjXuDWtc4m
UoL1nBTW2YryjSJBwX1PKSsHQThEXC9IoZ81jMEGSPevrtfZMcM0S4Wi8KsuDSKR
hIUu4HgKz3t9C/8+Sc8XVNAG1QOyXQn1T45fgjS6zLyZHQDzHRPdHMJ+MBywd+Kl
P+d8k+IjP7nr+G9AA575T9vh2V4G2jORgV2s/ckIkCWbRmiysaFuZxLfWENWi56C
m70DHJvy4+leU0y+H3tlMKRschNV79I064im2H5Or7tgD4zc1PaWJhgZo4VKVm4l
W/zdgky+7lttOZPVlimgjuhs1aT/1fQMZZVxA1HqEyT2OKi2eQhR2eOrgXrb396l
yNxERvIYo63wV4FTn/JukB0aGuQtyWAHCCwyy8jr+Cx6xw0KEd2OKszaw/AePY3W
YXHXT9AbMJ5ekFhIrE0hhB0Wg98y5DrmDV4osJgRRfeodTc+W8KQQda/QM9PwJv5
1VFtsD4fERm26hSEVTYSL32slN2FRjIVRtWEmHzcao095YvwtXl3WWMIwmYR6Q4i
OP3jEcFfig/KZvL+4t6DYsEoK53DkWCuCwPs5+sHXN+u2zqcCt7vIclzM/Lq3mEN
g60Z9EEZ+L3c9CPmpSjr/gXC21ixwNyQNb9aJcD3pFqt6WOe72vgwLYIlQ+lD8XO
/D5nazOX4lWExQavvt5FxInhVCME4etbB/P/xZLCUfCO3Fp1ajgSqOeNuI2XIoeb
UJP8vIPVy3h9WSUhZ8o1X2eUvglWRWkqoqPmtesO3UjB6DWoR/hkSIS27qKJK/+A
479Ez/vtx/hS6h1qJkCo3lE8U5KdBKAINFj8AHzQFpKTUkWSLbZPFZ9yJmTtRML9
FLzZZzAbou/phvMU0WwfgGd5WacEw7LtJrSgIygvk8t+HvZMFLgz3WBEZZZMadbJ
hr6DhFIVNTAQ6gvLp0msg6EOkACc3hSKLEg8dlZHP/sF1H5XiXff0kDeGH+cToar
iGyc2vTvtj7TonQ3yoHyzuIXtHCyaTEN3/tOc7RCfoykilmKJGni5ANMtJPbdkw7
9VxZF/PMnN/ykJMp6EyYAKS6rGZnCxniyp3deYLpx/viM9HkOLd4GDQd8/p6yjNb
dnG5UAi3+cq0gtRolKxoFRM10SjR1o8SjTMsuzzkaxTZwKVauugTRLuZ2P75pSOV
Ln3x8EZM86HNtx/41MwyUDZ+iNAAvE8xOQiHVW2fyPt410WQq0Uoy47xXceDRsFq
6++/onnd6cJnLRbqC3q11sjsbKMDkDvzeqAQhWA97D0Yc8eY8KfIBgUvNoQDtuPi
uLEnrBB1Lthgpf7WojssB/IBimS2IwTHssKK4CxscyMqppXnSp439t4DMNzaqinQ
hhCy3DAFvudydos1jmtwI+ItDEzGbpcf/WaQIMo5G6TjsSrlGsyZc0wEZzg3Gp/C
q+Kxwr1Yc9bblKXxk93zExNKNuPo3ett/k1WsvP/c0RxPv0mb7GQPLlyMa/2xpBv
dMDa/JVOUdUD7ly6VoftUt6thSAzKSq1GpEFAxZ2E8rYwfyD9ie6sHprXtUdfbyA
JClvF6mfMohJVVPrnkUSJuLzOxe8R0x2Sqp/jtkTj8Nzci7xlngDYkQfIYwxpa2m
8lZYiRR3AesE1OPPBwPnMPL6WLUWI9megPY95YGQrVhCkbc0atYo2S/eVB6ZYOqr
+BaUjUbroT1xTU2f1lUdVyX8+Fsj8wgv1NFJycMhP/Bmq93kO51skaxNo6ocM+NW
Xe7QfqMYZoLNt4U5bcGrycrhWmwStXr0Bk8wgdAhdiKcbkUgRMFyb+jdsen8Rk8b
JsQe7oIBYFDg12lIJ4Dzo4lP97mt+sWb8OrMbEpjy2WgDngJobfRAKLF6bA7of1C
fWEVCNAPyfMMPNqRzt57ANYdU2IGFCod5IQurnVyj6NUlNAleBw7NgAd+N1LzZBS
CbNZ5QaRYHsfcZvX9nNBAdZ5r0DV6J0RUgGYsFl7phHlfGPOmtpfKvvmofFLqVdQ
Fx5n6KJU5bToOimoDIL7ZwEpsEjuvWFidi4785PLpOco1hP8RCHz5VU52H5I0HEl
SPv+R3lnOsG7eou/wnQQMqr3kmWx+i3+kdmE1+rxaq9xodtJjLoH4qN8sAZR7SMG
XVkUacI0reaZOcvox7+81jbxt7gQJRqMOjfF0dPomxG6YfblJaVSQz/D5EwxvxLl
aOexFqFWSkzALno0DbaXX4XNBpenR4vFIgvtSZdA5Yi7aHWqWhqXdWUVO38JHqHP
PEPNkzgcskVqBeivX/XDxJPEadSTsg4TCe3mJTmlNn0fRoAMmHRsgjctItrodlJ8
vP113bYu9JJV2zgfYMnOC1w7lefTD5nhNJV4b+TOUMeZIHpfIgxe1bRiUqY1pJGn
SZ2vYtM4ETpHoZdrJWUaeWocViWwWgVPHDEAJujyzjTS3uxotoGnl5NNcTFh74vv
cO7gEhyJ7uyFK/62EkowrpUsFzk6i0aK4JsphSstiCPs/bSnE0Rd1oqGUABvKTEl
olN+F+gZoQPUBe5a8qk21QJ0BH9efdyVLfJHwd/qlzm8PCiXeki2nJYvwL837cK6
FDMNEnIEuDUxTvnl/9q6YLjAuPJtsBCcRaQzCDXhVGv24cq9NA7vzU0vrHMDf1et
++rZXGcaYdu3w1mF5QLayZUeZDHdF3fDFIMV6If6O1v0KitEBXWgRZpe5KxrKe/B
eYengoYFUY0tpuKbr9HHBWPsqMz8AsCrnGYTd9rafAj6Mf3bBeAZhGhUm8Nvithc
XNgv3McpNv+DqlNx21H9jjomxvc8hOGOxcLyGZq9TD90kgnINh6Fe4xSEVXUJLy3
2lBBbMgSo8DpNiH7YziupbJrB4c1Y/A4eEAMcgtwh5ltmNdIfjj1ESAikffFWZ+8
G+GipnS9ZVX2iEKt/a3l0ShVtfgnKOLDpOiQm1tWHIk3g7lUdQZ42d7dXeRVwDJG
t0Dg1+LQcr3CkkZsv4ZDwOeWrH6kwlAkuwRoR15Wc+CYt0+9grHtv3cj1p6uiUqa
Y1LMk0X3wqnnusE88WmeYfPkisCESgw2/OlMnBPnPGCIaXu+UeeWiArFbu+u5nZ0
gm5X1uhdOCr9nOx5+6O8PaKjxF0lVGf0S7+IC0/E+F7F1jGW/4Hqj7PPzpsvDH9t
atf1r+4oVyffX4QR+gf2YUI4X1DH7cTEOCxVVX8HMhWVl+mh10yT1szrBeurSKOE
CGHx2PxDELfY+g9Hac1rSIfj+UoYGP/o7JD+kBQuCchWv9Vuym793ilfjSu49XaV
P/f02Ueiy5W8XFkuH4yCLbZOTBbOk3SE66qY5XFP0lhV1B6Eez8UYHehr9anh1Up
VXm9P656Txo+RXOgP2cR4m7Al7v72xcUiWI9SUbWFeBalPGXQNtLF6h7ps/LN/Hi
3EHSaWMzLkbAXr7+sNPdp07jto5M42cDtTZMjvTqdmq1KotXQoO1Rp0MhpueZbNc
Mvz/veiFvL/M9xz8QYXCbt7hTPqNsSsJiqGRLtLEuTVB6d6wPF8IyG84MVjK2CCr
D7OOWK+eA8nwfA/zrmpQ1SpBX2Y/bMZYT68WZAqaArJF7MVduV36qqWWvw9UVU8v
YdM/fPUz+5BXrxdYSTPLCD9Sg69EZS4/7+0s0a1gqfTWDFxvCwWFGZVAOmyvEmB5
bDGMmMal5T7HJeB5VscLW1Peu4uIwsK4V2yPVESgLiaKih1m3rCzjR5MIquIVEO4
bk9/KSY12uY42NEjK+mFSP8NU3tPebwrFM6qhlXsEEjKd9iolPyzpzYb0qn5X7fy
lKoQBFs1unwDy9askaTx6rrScSp2Y+zezXZvqbx+7iQtvxVafMZyB1ZgMaC9KT2p
GcamEWAq3UdUEZ/ymgfsa5eX0geHSul/COMil7BTDLoiirDjjLYdV/67FehSU1xV
ORhrV4vYsizFCaVTyUdLCEh8vh0BqVTqTiTQJ1nxXC0TwV7uVQM3Firns/XMCGNE
UqdWvcuys6toyB0+f0DxXs81KOjxr39MOFc1WZh1bU42I7Vo1t3pOSfq8ELNOilD
l19tt6VWxhsL8uebvAYiktcJCZQbsP44skasWW50yrFB1eLjquW+Sq/HvgnSz5oa
vs70QJPrw/2wLbXCx4vZU7ZjSF6YeOY0fTD8BGpI0y124a+IKFIdBd3/HgrTUINP
tRVg5v3W5wvaYpIJ7/eBblyJw+cthcH2smph+6cArzv6t5/j0YyoiUFnyvPhH035
+HOijokUpqXKGHGpY/OAhJZUc3BD2ZBWnpiQxWKSq08MNBkR3+MSUysiyWWmXL89
LNVZ++5m8ydwqVqEHrYjj/ykWVsrmBLupADhhr4OT3RDt4OuCjc1jVlbn5aQVWTB
E/gdsgLDViTRKkdDYG27AmJgPUCpAwtmLfcI3lKpTpqFnUriR8DfyAUtNc11emyV
j5Hgx53ycJUcWYvzP80Q3SkMGP1Hj/dEiS6dqRBrz0UBDJYm/g9x8YetXqGJiNVk
b2IsDi4QybqwpfSM5MP1lkz42wO79gVgqybQ5fbZMeKRhKq0AMYq9oEgZ4b5x/zq
hqUCLGYfMBIIYJIe9Y1gKyX7QBHjHdLP90h4OHpx5aBxYYpFIBAST6PJywDopX6S
zvJoxFZvJ/m5PYJZO22yUhAzichQ2g8BikPKZPwX7kVjF3smT8p0bIIEhuo0CJ2e
U2UblH2l9HFwgs0SM4AhN9U/cYaCY1G+c1MyJzOkG8KoDOri65V9GvPbBdjYcx7a
u6j84+RYZXP4xYq3ABK+ruBbjbR+/ioowtcV7Tf0baPiJ9wRqgoZhD9WsYbn6wAO
TjHNqQdmS00VUxEU6VgPkGcJGuWPiU/b/9w+LDYcQCaxcNSjIaVf0UQDvLxwdwlY
kEGLLBKlnHYimUIb+AsUNmDfbjdR4OHy4+5PVfxl8kMTNKKEIPD1ql7/XMAGQpyj
IJ+cKv0TH9oQAdiCbWLvrycr3y3rGCA+x9OK7axzALoSr5Cl/Lrf4GciTq+r7neg
ZNlHcMj1zgzsX9panjgOymCdaCim/Wx7P0yh7GweCY1+4DuhKKvXHewKMK/XY8Px
ufwiGQa/Ixawe/Be9Eirdds5EreF2pX5gHe0i4Z9Jkh6abKPn3YRCXqHjPjG94oQ
KgpRH0Kd0R8ND1eLNv4W9cu6r78W5sLkOxNWiwo5llaEmtq3agrpOU7Qy4mY2QlG
R0n10jxPvjziDgHusJiLINg7O8bCaW0HEnDUZmhFme4f7XK5q4751oTDGFJLba8l
oyor6YUhqXrCTJPOtcHXw9tBfNoubcsyl+YkH1mLM23FEc1jwx9QWlkXRORUx8IF
9RfoBGKJm/oGgFuPhkNspRUS+t8G7DyjwdSklu5Vu7JCkLh+ucWQWQZYX6L2GtB9
boJx8wEHgi39edh45WwXbvO2cr0tMjC4WaOqjVlPzerRf+lo4N5EZwHaLg23hyIN
qDxOJAJRKtTfup0Zw3rSnwdsAjHuU5jpZ0AqmXAJP3XnBymnSfqDRNb3839XXXjo
k40+AAcvxi75baClC9OcPsIHi9quDrJrX9Z8SaRCs6Gu+6GO6w8UQqwb8bJKouHo
S73FsP34aaBel6LLkX5CQs3wrKrmmUyvMb1pKp6FoNsn9u8J/zKblh+JiP/Zw3f9
dBVgiSTfbILg31aW7bPJnn8Fu3DSLZuyi99xGm/IP6Hq/HJba3sdYsMTzcNn8f/M
WtO6h8PRxGJ23gAsslSyvRs6FyFyHWevoASKY6ahTMZ8RgAevxwE1c9d0zwW4SCs
Nm00PT4ma6PB9bnuI8eAePSjjeASPSanHrucP63aWlBiXYSuMGbK9Fnrq2vSm+3Q
FvhoF2Y0ue0NQi8Zux4bU6bUel3J2XlvhNRRVwlCDmW+pI+Z8LLB8wWw63p9BeCe
Cx47HpB9v3l7TFOEF8ToVp8+qjQk63muF4vV8BXR1nwK+4rn48D4A2tvfvE8UNSn
/thC0ol0mH0lolm74qEf3TfQuzqbfHE7CI+AUjEd1WEDctJb+IysF9mWUNaD7UZ7
V6FRRPiJldwzqQzjQcdWMexWz7yO3+Ci4HBTIJnXXar4hyfpibfcj/w3bIWRlh0e
qRzBTVCWOd9kyXP9ecDD/yx7VXB6MynmTOlAGPWXTG0WGqNB2ieZWT1L/3bM9zku
VnrqIK2jLAnN/9SRNr+GYWIXa1o2yH2JjLU2nPr/EQRRhq7P0E/LM8mGk4u7quN1
rk1t55e7wnIoDUfayBCZBwMiWKKpLPLD8naLK2yT4lMfAeaYm78sVRlD+Rn/snkq
LsMD8UgkAJ0yWoJosj6U2c5UfiojKrh6xrNnNcSU3f1PyTzMGkcOOtwM5rMm3QPM
RmPiUZuULVVZBXJEa5HQAlJNDSHxwE4du8S2u34EJpCEolY8wBkUq+96B26nmGDg
1qKmoyeQng2nbd98NsRWEfaJ5Kc9mfbk+t7LYQy1EpP97Q5pCwSI8QrQsYoKy5I+
imyc21Z3fPSxYwzX2ek78PHrHojqlFYkmJ6WaxPHpU8+oY7PvR2mTlrl8/lQ0inc
nVw9qK1S956VV2o1gkFI7zJ259Ci8IzEbbsOlY3ZKWkLJ1s7dSrNCSfp5QjKBDVG
4chA4zWhYpzGB8jRBoLXZBPdpd3DXT8nXBQy4VmU3N6n+WH7OSaMGu81weOqlYPy
b5e5gWIXjBWs6ZprPFw9oyeR3gb2kaADeXLuvygSE8zHavX4/1JllyotIM/A/shC
7sUUhEwOK6mRSKrpFQY338u8xLEKsJGiisoitChkEeKRhMd1EIin0pFj+LmtQZiB
RGK6kxIBtE9ge+S53bkvBr6mAXaQEVwKMJvoI7XhxBM0akzoBiILDOUHsRKvXDXz
DGDLMaYTDgUinCZPBPc7hplNZ0BjBRPvRGVp/w1l86pMWLqoa7xkOVYuoW7X16Zx
JAXenKBkkVwslxwchsV+BPFFqi7oI6yom9kursffUTZ2qjfjZWxUfLJb43avGTc5
8F1/A06CVjx49cm+7YaDPTWJnfKhxCCU5/jky8uZOsHqmuVylj84qYwz2Cqffavg
ap8dpNu0ZegkQsjGhWur9NDA0dVHtMtShzUFKMy8cJxYZR+hd52phaYsCC4UMw8s
L/u5tEDs8idPTbXKSdTsAwrd9pQV5bq78PGjQxKvpPFJHNgmNqxw2LaQwxIFyaj1
qFWzm7uTwhun/23/4XpBOo67WhcbhK8ZjV0IrxiHUpsE933WxGBcWQ5IRIQqL/4D
BwVzO736V28tKt+Q0xM4MSOXnI8uZB8Tat1zgvpyyB/iRGvelotXyAnVm+he7N/7
ZCL5MQdDRXMaLYrerNM783vaf/PqUdvNkGeqVlCc/o8IafR5TAKEfsYbObcaINrg
u5QRC/pcWjCfZ0Zw9UAsq9LymcnuSMSyCfrebKzkWpg9e5CzPiH1uzDTqmylRd5p
yn/RLJK/6rlqd0r3RM6egOLaFKgmD/y8qrE1v4fKhmwHNME9cWP+i257/TtH2mmz
CziY3eFs8ONBkSytiV+zsmApZ1jJRXDGH7u7fEP5To9kgeGsd3bGSL1Xbb4C1JoI
YuNpEZHG1W3P0o+4Jwhn3jQNv1h7DKBNYvg6UuEbasHSrPORo4Gy7xYtd9WeSF5M
xOLKlUruNr9IreuXtiRiSsEN78aNf7LvLEiKdc9HHDWNWB+VykO9+eV6TP16JcFX
v7rWfvB9HJebgh0k73pLD4VAbVDueJ4h7j7S4LVqjkEZoDVa/v4D45q4DwEYBIi9
14+g1mbuO0y3i3PU0EWmVo79JePVJZxqiSMYJGe63qSrjkTCkr26bWGJKlZsYUpp
eufygQcypQxthpJUybNSVXBFn3YSl/n/stuQ1M7HLGjyb6HzNXMCYcL20IDX3oP4
eAC+pJfgQrOeYGyLTnJnU6UAo5i1/DSF7SMjlGgiFtsBTqYgQzd+5I+5Qfh6nibI
T7ex5kPiZD4+IPSasE+SZQR+auV45CfYn/VdYniO4YjHtkkkHP9MLHxZYqOzOP75
plnRA1iknDZZpIWyES7vT37UXj7PttmRgQ3WuTmmqnHNSNqiUPXpjSUug11ktu+y
tn6HxybL+ePDyPVbjQiX5sFR9x4iHSwxmv/kLmvlR71votW3+llga4uObKM/xSDp
3hrMVwHQyK0g/DuMKFhLWPbE11c0gWwN6gTO3EEc6Rbwde6QXCsWKvZf4E8EFRgY
LK7FXa4sj4QLu8aHB2JyzhJHdyi3/4kvZkteh1i563fvMUPxXoGzm8b/MBwzw75B
EFxZzU/4iPea8A4IAVBc+1774aYgIGF3IHusvL9lK0xrR/OSizanXlJJTEzEFqEb
ucf2LvH/8k9DSLe8sKAkNbQ73YE0C17MlJN6Qn2PT1oZz8PumORU62LBxqM1uYNX
cbf3b0VpyL/gqSpFZ61GibCy8BVpZlhXbIPax0UbKRAGZlzUgO6CFN0suuWvm/SF
hTHWnySVpEKzVekfV+t7p5t762LAxIIUImlVHr1iMOVvw9jMfEtDzIeT5baeBvWs
7ooYPlO5ZIOM5qVSPXutMgNqUwNNTvKxzlagjtopn8H/KMSx/+YIhEEZyDyNzlvd
tlWPgq7VooK1tPPnDIuDRBXKA2jKfP7/VRuf9mCC/qFUDR37ggUZicDbUbGjI0S6
8gOahx9C8jeNhDt04bqEGBfVMWuWibIYyXK6t8NPf0+pB3yOLT6NaNHvNEXkQL+n
WudA3szpLitFHpzy8kY659+ZJAclog4D+D5k0n3VE4hSIQ4bqed3aH2LapHNILSn
wClTGox79bHTmr3D9yQ/83wtwSDZHqxkpFAdRwnYzGwJAQ4qckXxFPnyDtV+w9s/
xaM9VTYOAPCiaIiZKLASvWFFAHBk4u1KJhvcDzyzPmlxiXpgllM205KvzhDN6rhe
RhiKVqfKo2C5pibblAupGXhYQYQX5E5+vmG8peHqzUxDPqrHZ20+BhWDkmMwbK9I
FDj0nAZp8o0zAhuMp02oIgWHRblmqYvRVaq0wQT0RsQZMazXX2U0RzV8zetOahOY
pGrX8Oras7rqZT3CXuKfpaC6+ixUvgwoI7lAz8cyBf1fmm4W//hZZyuEfl0egvwU
I0XMq32bvlk3x9084mA2rT6N/zjQpfyDrytyDS5f5uWcwChevOCus96Dvf6mERc9
0Id8KxOclmAyzEvIZzIsWy+SAC6oaZ/U5ghW2E2N3lSBznzOj2Em5NkmlWWwtjXL
1KrTjm+jvkYlVintnjJ/z8Ovx4XSqFzXs9JhUgzvi+Y5SL8JN5eiKH2hFNoGxwYM
79wn1BYrsZgaDncR7IX2StHTHQ6olUHHqkN/83DhSqVz08zs31XNdpnreeBpfQ9U
MF8Ytt3sSOw8Rj6D0bRT9A25dUVISbEdREf9gvjr4tnpkxdUtLDEuFFgAo91Z4Fe
MHdr0DdsgkSQQKC81Ry4UKYcJ25tsiKDbciqT6bqWAD7BNZMTcTeYufwDhRkj/NG
dY0TKzm0KwNDaNWWaVzX3InKzGsTb6/PflNn127HsHZ1ZvLAQoTjsvAq/Rl8rxit
oA6c9GBEpjMmTpi6NnHr//K0NoGkO8lidiWfoaVoXWXi243oPuFtofo24IYmlWJ2
umIZSmQVmxBUKCSFXYkCt7vtOgB4zJdctLnZyZgMd1NWJtAtscMjVoKa2d4jCkr4
SaBs03AnHKzvkpTifcWLcAZkfNg+Qgtk6TClVvfkBMlXakDLbdh0a+BTPkU9hTiP
/mTHWZgj9olpiW/6omRQPGbhqqXhaQ+eP79pbDgqSqXhsnPoJqDHbsJDLnZsAIxx
MZvy3mM2BkjszDZO37dYk3T3USfgmJYyeAhTWL5IPsTgDHszfD0VkdqJo4XE8pHn
Xhltorkr0b9qN3mbKNawgCC8bT6VyZRwhZPsZKNQaTaiXGl1l11z5oV7W3u0Fuev
iyhCrSuijDM7ovBS2yLy8JiG9DPhjQ2EBWA15jZDT75WBElROACkCgVAUdH+CCe9
QAWxy8ir4dvCMQaSAu8icT++JMdRCG4J6xdZ/4054WqHEol+RzwCGnKYNlanGJlD
nPRTlxdBx+wAZVqd+rogVXudN6rdhU+B41Fo4+98brqrGX7gkXGNdsvE3KRyasPg
b85nA3rC/Ea7nyN9VtVU9oOpjcgU49uFfqrBAfdXXkv4llo9W+vSPdi/59WGcUGE
DJDI4Z3fDNjSEhtwwVscohpyfvNU2gx9czNFT8zSLJ3AkTc8DyEOOXzC5ZIMJhvd
an6BKBHpmyaDWpD9L5tGrjoPc2F6bNQNWztwhCe1GKjk3XqADSawhgeDiLGZaYG9
DHgkRH/CNNs/PEKjwWCOL4DR3KWHJl/xcBss1MsVR4fHJq1XykiWOABtCLdXcsrr
aB9ocdS4pQDm7mjlIhEsM0rPFUN3Ps7hihBcaCUeeFaCZ+3rqHenZpXk3e7PPVax
wQP34IEJpzL2kNsq1VQFWTUt0ivBHN65qkeDoMIuBcsJ/5AC14lC+VGDt1l1RH79
/YIjH/vMNODLyw5XwGPifFf365zru2gFSjdLg9epNbzz6VgL38ijVwRlMSH5j/w3
61OU2OqfEAL+XadPfrh4P04wKMiaXzki/ZXXBjn0W2o5zWfOUfV7yaLd6DURd7Fs
OLLJFzg8hHvyQDanVOOeTY4JVoSG5RcrBgsjfsZf9c0vJkIwhIyGfv0Xc5mKiWXN
A7fgnczZw9Cil+Vrc3HyMXQZJVdxJfPOGLQSN2x7TwPwPxxiix5DngFDfOzuxhW5
svgvX6pkEeW8EfX3/mMI/UaZc7c3gw9cx4uO3vukfTYPU7a9VA6YzB02Y2k0eYho
27/d0BPMg3/OmK3GNlyqxX2v/D1Y8Ug9AIdS6we+2nf7CHS61QViNovBbk2FQ5c9
SVsz57QzD3EcPb9igaPDVXv6FLTeZ7Vikn2e8Y9JhnghqeqqqSZzIuNCyQCjDCpb
+sLruCH63NdMk4UJemMw3W6dosqJlHtg1aaghdeo5jQMOI7n3/kEAIdbIlGN7myh
h/JZw3L1ofwxBdJCn2/Bt7C8cAVh2Ioa1tveX4Uhb9HNj6AJqZrDlpA+bYxJ89u+
jCESmSD6YwDG83opy7q8itUUZsFAsGaXCJZ3Aa2S76TdJ/0zw0vpZkGMBTKfZ1HT
KqKXUK2BPfIpqxPJ566RFiup4NqYDpoUpUcqrL696y9U+eRH5+g4yIiXmOaGbN5E
ZRXMcy7RW/b1zq6yILSAxA7ZcRNxKzD+JwqM3s8EZWorzRzFsDyS06H0bPlknXLe
yXyOVtCPhEbxRWK4L0lYRLbQn1/kuVKtJAtps0MKKJUUjI24TGft0HL+Qio1/B4M
lPIsQmgFag3AH6egFMmHglRiyHiKdsPHkhQ0wFcPsqVw5M3pnqad919Dj2uzG65G
U/4fdcoQbc5ZfJRu0VZ602+jH8xY7ZguUru7b9uADkXL3XgoW8d3v40fP7YfvFTx
IcZ4Wsh1qwpP8WVZYyFf8qyyug34WV8Egg/1Gn9Civo0QOYnOsuK9+04BNsXOcWV
RZ7aIfgmBvsplC6bUAOknukvAsHlWhIiWXeybbWnI0a+Wj+FlP3l0z5mZcIUxVk8
+MCF6N1od8xUEVYaz8sRYGlgKeJUsVXx5VQusS6gs0gZBUIlA4UZJvtWPWiavlnq
9Moo6rnPBecrh8xQeUN7BjbH20vwG0hX+1Ba/Gq0WwYk67jJU0P5lEJ5ZmGeio+j
tLc2expD1yCFiHg+VVz0OFqX748KcGmr2MT2kT2lHmA027X0lZhsNMl5yYTBFxwO
XuFY3AmkTfpYzQ01pt+PZeXB7Qui/GTtvhy7LlhviHrAaR4wyDOCGBFRZnlPY7Q8
SL7gYzv4oGfCvOWWfiAMsLiBI3EGqlD5igXrx6rae2c5HTFcraxObnH+WO78u4aN
MeL1tvgtT5Koue64UO0XIsrxZRC09WAxn3y1bWjFS0kFQ9m2PMjQpF9vXLbPQ9TC
C3f5N2zfQhiUnPF9CfpsOAkLJ2ZASIHnLGF3CRHm6+MeafXPkzpsLUWxrh7r9CZw
lQhuh9IkjIp9yIvyU+xjjE3j/81do6YG5zDidMd1xXYy/ZNZv63z+emQrSapdhEV
6tqrnbZ784Rpx5nj7P5m9GgNwbzyN2tb5N4btSNhC/6MhLLIwRxXbO4VDsUiO64n
4+22n5JUaT1kYnc0+BqY/0J2ytoi7Xul8JrEkZ9q37H1fb5ezbenFOUnIjTTx+JC
xl1Sbc2Vjd9NEqQz9MOkJh9UDGBAS128jzPv4f6s3ORjGHLGnxtCF3/eDDrSog2y
9AaV6Skf56Vkapn/EIUiABeazc/eGG3mVZrmlXipW791Erna8X64/RQDbd5VrVsQ
PI3LCyb92p2fY/Xk7aKGtty+omDFZ9bVv+MKyIRhmEQQ+lLMaYEM90A76pXF0cIa
HhE3DpBaAJpjcc4qpBfDXfbK3/RSQWPVkrY5TGL+FhG4JY9zWLJL1QFmEduLL9pp
UMQCEklsV2GlwdZLAWQmHeyAAFjwIsrwmA/GwduTPy8oJHw1ZOREBPk3S8/yGFq3
X4sP8hFnaTyTpTb7UHidfps41ph7+On2Zy5z84UjCwt+16ADS+6XfPEZld/K9CQV
NsBrOXy0FgPi1ZPS+WjBb4iXBjv8aK0WDxfgQQNMoAOUh/skYzlIXgYsrJJYL8J3
xmqQeAjj333sNdYKeyTSyFRewk03v0RbUbXNKrMu626xQCNYC60YTOMgwtrnYl9K
fIn+pRVevbqY32cqY750VKjurTSXE6E5ImgeCKXg/wIdRl96Xb75UdRKjY/TwFTq
en1ty0ByQryShRfBPmojPW6H+d1fdoAsw8K4SHoEiv9Oug/TAHRL1gZ8D8DKuYtM
QrbWVVzgl2eu2/3tNGqwC23CLFa2RFAKnrb01HVxvjb8MUjn1MtlIC/nhc3qcoir
GuidJkmpvAb1DRZnmDvDa78Rkyvtm7U38XZak9gzMZBqmT3GXHZy4I4qWKRDJCjd
j9hF96nj2fHugpvtoOmLUbN3KM80mp0/4dHCGEzG0pPPsslFZMfPAcSdt+iB10a6
LA/VA3WVsVbrQ0LiRcAGqc12Z4AjsKu7IhsNLELFQZu2pLvPSUvl0z/RvejBxCpG
8qD//6s0vIQBXbStWg2z+YKJxO8OGasa9dN0V7IMvjI9Uy8nYZjIzHSE+StTaUx6
3EWNMHsKE/Z9SFZfn4MVE1kXL+z8KNmGjYbbgNLeCaWLz6m1JfupyHrF90GKNoaZ
v/rV1ZQGMI9+1a7kHCBit0MwCKy10wmBFFnwEcUOBPDQw0Yfvi7B8hSS47H1f1oh
VbHLeiTed/cF5qPKrVizmpFoPCZiJfB21U02lxr22cTlaBZ17zPTgj1Oux9cKYQi
fRyS9acMG5Ivrg5QgSD7djxuZi5ck1qbMIeziTlh0Kz3fczfe862e6INg0cbhq4k
WWBlPg9QXNxWb8nyaF0g9ppcAk5Xfp8ajLlW5LlULXsp57nqNHT6AGgeIiy9S1lh
F4m4+16eG9tZkiVZ46op8BSo4pqiCeIqoNbSv8PM0dirEeYSYESyAWpJUFx5xKyn
HFVzJK+rSCsA47rqZ4l9S1AJSBL7jazFegmPYYWabp/KS+PuYx3SwZiivpawxdOw
9diDZXQVqhepZbxZvoKOfR4xJAGhCuBUeSUu4IdnFuEKcVb+ilKpvYMm4nOC6v0V
Py7Dgp4E/fcbFudJY30RcnBALE0oHmbefXyZSuP8QDumq+/X4okUkbJUEsETYemC
pqk1chhkpv8Zu3iU6Yt149By/4Yfr0rLC0Iatpg5W1gFlNxKZPC5IMux4MbVTRas
i2KtYbWFt+NH9IsE23aNktgWMNp3fJMJrxjJ1MQg4PwbnwZ0a9MbvVSgzsdNhZ4A
Jkznj5wzTe3q8fcFZ2s9sr0fK3h0EZ0AIwjDcQk3iCReI/iJYkeDJ558r0CvS1wo
QRD5IPK+fW7J7vW/LikFbE69zNy7yJvRiSx3yR8qSQunKmh6cMcjJ5T9qShvwdpq
n3wqjghrWZspjA6nHLM3Am9ADwqcCdI8iCjajcVIJzK3IxbzRq42IbjHAGdDCdKq
uKrdI92DmhnY8QY96AAbL47z7UWVG4fM++1EaFtoAuAHBo8Erq/h1flojAYYEuIS
SFZKqKZqxrIw/a3VsPFpUyYn0XpETEDeth1PEX6CJLi8QHaH/wAKert016L5R1ya
Yyus85bsaC8OiZAuZSMMCVsDvx8twvJCx6CdXm58l7qV3yAZR1kyCWTYfa3Lk+IO
ImXlhYuT0wQvm4JBPBg/W32K4hpUzkXvZ7+xq9kWsbRA9MTOQTy78WOjV/02Rpyl
6oGbyZfU6bAqTF2th3r7UyNx1TAZReLXCwqqDjzQWz7jNOdDkSoFuqn6kfaqQFdS
i85B1aeBjEfgUNVMKQpWFUpGjsXyka3or7v8pinuw4ZjheocnorQY0xQeeE/CQ9D
DIHbMlerZ/aBuwLGVGOwzSWzGrnQ/BahlbEQ2ep8Ed6u15/f8ztCL6dqB1HMMiA1
UoNdeSoZmwVTrMvSIqisKYrC1HHYjUD4g1CmBh0NILTq6l7Bo5saQ0xV/0OwMei2
ajTqIToCeyZhHlYguQfNZfwcafay3tfNOJetmaKW13gR/CzrcDGLgtVPqLSk0obl
EnGZgkWAPK59HqTGQuLgcw9rHRg68xcKj/pPBXMKHVT7K8N49lbyJD3ZNapXUny1
EBjsfSuuQqoAzmhIZDxPsSysQdvU93OvEnoswwNF9QIDyON4UOTgRkjry+UM4pMN
Ht98VSLTKHshGDNAcsAP/7VToT/ItXdCtWe/jhLmHUSFIUV4EqrAFg1OOHSDT22D
QgJ5u5ZGJSb6kFULw8DEMVjxqLKfNL9Pir12Co9jO8mkRQOGGahXcyPKhR4wuhqu
F74LxpjFxjOrDlQ5dfYTqj/fbrEtK7NbK92MBD4m1OpoXqKf+1WEI7wewXYqxJ7i
RVqmFXrw2bMT6B+ySc5aOw7ayF/3LAuD0SPwa2Pc3NN7E5tmX+Zb8JJzIv3+adUl
jfupsnjzeXOv5DpsOq1MbUdrvhCZolPn4EB+kelo5IaO/XI7Zfixei8s8M9uMepS
AsHFfDpJgBIj49Zy2BRUT9G6jc0psr5IEI6KfyN9KinNMVTVZvXD36HpNafKsYSh
y0MSc8wk+aWAAHud6yHolC2/boRU0uyz7Q57OCgOylqY/nlPmz0KNRK699Gt/AUG
KS43DZl4dI/DH+LzXCXVzvnFZZaO63UdGw8WENWlmL9ww7AfX0Haj67gVwMp/awM
VnKdDjU226seNJeq2K9lzTPqD8hFt3iGAM8vqqwbGEHP720lfKq57htl6392AGCV
AJktzFBydaJvrjiJA63Qlbrir0aOMAZNyhAkEUpQ/oRfDRSnJYxAYyDVNPnZLIAE
8vIN5aB35VKaJMt4FHafQro/64Nf6SYCztzHegEGB4Ysl+KcwOlPZHYTr7aVzh9j
QOBs9PV3PO/RLSeIZGC6IAPF5RF2LqGa07CGNqc6Ye6PwCEJzMrsIaNIWNbuX7+j
4y+ZZ0CPOFf1CYJEF0yWYroLJ7HO84hudYXKaVNXTEJVOAc/0ZLRzm5dXC4ctA58
gMef24xCZ8uSmamom1tCXjT8nrf4f+biTXHNStLs7D62RVyi1L7mZHm+2jI3uBg9
NmOD7xrIhUo+z4L57BDJBnGHjnPqX5V/2+oYYGsK+RR6CeAwSBmIwf93B5OimY7A
mDWqxTjpbvCorM8bsDTLf+u7cYOuCt2BSFj94QUnYikxvvMpno9ihKfzBcbB0ZsB
1DWt2Q7MuZGLJGX2DmiBE73VmYkD0FG6uhQSrG+n6i7wZR8XZm+VHgWsexBsppnS
rGKFgnri2O1n3hovqEeYo4H4TiG49W14de+WgRs/5DTGxBgn4N5q4kljXs02ysbA
Aw9Zcyoeg+XLb/P9fWicCK45ijN0ojhrOIwMhl/5Cs0uRI1oNaFvUoRoLa6D286S
fSGSw7l+HjTzXeQe2cRily8tBhFdV/GIcyH67QTxJVY+T51IjLfFCE10SgYHqq4n
ek38C4CkEeDcasD+JJP2k/jlfRog0j96NLz1KdbYCObjUlajAh/HuS08PzmCkkWl
/paQX6B6V3PI40oXyjn9y5bwgnsxK7OelCC8tGz86OsewXSDuZSgODghqTz/nBj9
weRW8ktMQQYsHNWtqdsmZLJFo//rVQF646BcXACY3nmsz8pQzc11k7o92SmlPA8Y
W3BmjYhyY+2lEpYdIhEC8I/OgiRQw/isyD9eD0PmIXJfX8/yTLntQGZEyRwwn6no
XsK2gWxmZz7cshCPBuz8Am0S92Ms9yrdyEOphV44mGr/mqzLOZgVHV/8c7+/F7nW
/uS+9jvT7hZ94tor2toYDcU83txg9fl5Yck/4H9LAs/8wPGCQpNezEG/iu8wIxIc
g5uQG5MrZhLkhDtx1xYb8uR5Bj1h1YcbY9HPZuKlotUoHvNrAqJKKrl+vG4mcs49
lmrKsj9BVmlQB0mhJyQnBiz3HnGU0BG1FtD8CPrfcPOAMg7yB72r3X99R9ax4yJ4
4WcuhBaFwcUnr5DtWNh2tfI7J0ACuCw5/7AqdBoCU17x3THQdSe+0r8zkF/eGSPp
svoHLVJmDtENcfuZB4hqIKzaePudvKkMoSyjrpSTEQbeAwzRrRhiQ5VFL9v8d8us
74Wa085oagxKIJlcqVlqpbkJZy8dnOcjOdBU+MVSeQODho1E515tlN3SmDlcRYFq
GNm/WEhXaYmMOW+dWt6WAX62R1JxxpyDC7yKPn052D/Ald1uWlbB/lXaYOfAQM0l
vNA9/yZiCtfSa7hjWFtaiXAyIP175W5nASdCBRIU1ThMLrQ0T3gDYda4Xj32Q5x3
qToEKaRSxoHnwDjsqqNnEDkdm9KfM6n2u3yHZMyCrIaM9ra9dmijT0UovCreOMMU
OieB+5rNF5Co1ypzEDEJmKPE8FfMFARaJPywtd/ybuwmGqvLcRx3BkE/qhEpg+6h
Vnp9SK31N2kAxui3YrBBAlzFlJ/1xHV/wR3SdFgV4smigz8jOmm8FUwI2a7MDc62
Q5JJJ7+lFmeNO0j4pbuQiZt8GDBvXFmM2tHJVns7Mg0rgPABD1pYxhuXHIuz+Nru
qQJgd+oR+vC75EBWBBnaXKg0w5U3q2+GHk069o6ackn/vfoEBVNbealVTzepZvW/
8VIoSsqCk+tZr7blF6NM2V1+hdrn3dJ1eYsxd+H6uf2sjMkABYvdI0ubZPlepmFa
MaKNnyF5h4Rbstc+mJUGsu1JtnhaQQV3dDcGYF1ef95SA3qYYyztyzWrlLRaYSBk
Puh5byP5RYjIR4trX+hr6g5ptvHbUM0WNggFTxBP1BivGvF6bYuA2EVjyqTP+0h5
oFnFtGRoNicXj62vGixQgHzju9illc46UhzGHRUmAw4fnu1xcMfgjnbsWdnVXyCx
z5jb/Q8J7UThib8MipggRntAwr5hrlGdmO3sDXV10l2BCkIdf6sRA/JjqkRrl4NT
1BWSY/7xUzI5napOAnlFd4ygNBwweaSNt1Zt5Scyp+jqRoJcXf1doX0v28b94Tcm
RtWQcZoK1s2MjufVTTPlG88tK78orIzwMdMvcrnPDNnkq+xTeu1pT7RzZWsq123y
JKVQBeT8SgDl5KysYE+ullMWwct/Bxf02WLvB+y/7ZbRSTuwsjY2b43SMx0H0GQv
A1u2iaZTPf3W0GypGU+EFba/oldJsghO/swA4w2uw3xdsP3AAfEJJMWmgmh+AST7
1imNmwWhU1Bw/20fcAVicyjyjqkRFu98ZQIZ9w1vQntEpGUImCcvE+4luqxLaUo0
LyWC/v4AzBoxbdc8nNhLm/whibjzX0Ka2Z5kq7pTajoU5INWs3ZoEBu7VzPvF2S+
BWStRej8dV5vDM1ghxun5Z3Eq7Qh4GiR++SkTFFyNRuRlIHh50mlUuDfh/S2jby6
Egy6etatA5AJHLIhk31e5l8Vo/rRc5NbKFLvZBcX6oADiz693qbIC9onFcIMnwEr
CZS8QTeM7gtCv4t2wyph7GKUT4Fiw4/4pSEW4RjF6jH9Wl8pcboJIjZQ0My0y6Vj
isYY9bQHwFQIeU94CxOLwqgqR0JudGsdYOg+p2s3xkYDkmi5isDGQ4R/pW6ggpeb
pSGG3+taIuVFDzsamrtXz9WMu9heWMdgI3dElhcIPnSQ+8adMPsxOwUtQspjT/RS
ASn+e5IR4y5sDo43CMVZeba7qd9fV09LSxl04kWFPEabmxtP8f4PsHQ45o+Xwwy/
4eTfjjWKBbCgMuk+tJ0MGJUmKsQ0FvI7jJozOJMAychfS5oRdhr5RMJKIJJ4dQHe
Td0EGVR13Bu+Jj3/ZR2sUdWueCpVeTMbAtCLUOaOf6ZFG9vJVP2FcBcMOaChDY+G
BVH0TQJ4j66iksJ1wfOTcG1QBbFuJepwrsf6rmufLAv6BHW/+KhT4tR+9SPuVVLC
3rbApomFt6k6rDvyWOjaCT3f97yPCZDS4PO3eHz13mO2v8h+9i1B5qE9WT0DSArd
BvzYck55J8yv2vjMV8NuPd5RnEbM+iGI2W2twm/H11TPfvgq2ZHLlT8pdkf4idxN
J5AcvXgIcoMaVgeZnMOz8Qx/IGi8KwSUovR50FE2qLd3tQW9N+BkMzYfxppb8FZ1
Ror2lHBoQOkhE6XVTVuEr5Dn1EYAsLN3uzA1A3Zu9N1dLeYga6sb6nUfLeNBLV6R
AO8rA0W1E0m89qQZU9QxS+uMzA6WDFZczJMiA4yLlHuL61MkHiVOXDQJbBPcB4L8
ZUCWnoffDr8FLZyO3SSmcqh1EnD0BQbbp7qVRsOjzYLUcHBGlxK9TuduSRImYReF
/rp0Wzy2v+VAirnpLn5g8U8EeZIxZKzkCvLHA5PEKn6aF40+lWlrGVMVRliO8qTB
A2R6gSL4dz53NJzSdDRM6vD5jxuSFbTKijTffre6Qal60TNGx6+BOfVFOcLlxQWl
nmAxLDfAXZr/9kW34YHPXwxm6qtrbDU4QvOge3WxegH0/Lb9ICh/Kj9WiVmWpSUH
PHTbU785vfkB1LLT6x6PLn5OSb/j5AQ1J5SWfnzmpssPsyQAV5gqVsjr8TAMUaDZ
MgHDfimZB8XMGMofJo/j9j8eJMETE9raQKDCjYNohV8eOQTCkrmcbqWWhPykD/lN
GtubDHFIgpJdjtkUvdRC6v2k7FHgReqraw1sNYHerJy7LmlxOxnmVZMJ1S3DG3ly
Sb3LF7+IdaNrL+nj2W8/49aHQc9kpPuX6ORC0IhIUvFEiwvG7fWpAOVhWArc2bbJ
795sMTKHCUTU6mPED5RR+gQ9l7Gn8JMdnNzfzt9PlVm3zy3GNjC1SqXK1B2iM71M
qYCoo3scJg+R54CKOXqLSHK6pL/XCJlpGzhM9QAPz46twYezDzk1G5Scaoml0N/F
HFQDXFtpmiobFhM0/L8XBJa9yWzOc8drCFRGJbreJ2wpJz6bEpOXXUDl7Hv8C/I3
0y/XgQD+GIzUSuWx975zCz6SRR+VO67rWPP+O9pP80+V5T5Vgrevt9QLl2/2J1By
nH5B1dCOiyVrGN1v8ITosQdxL3DpUvXh/2IBAAOgca56Ppuu+wBtyktem2hh4pET
Y/p9klpSdiMsnPQ/d9uQClMjOvAzXdZMka5I3NHmLRaP2XdMQTcPPUSP+ZcV3nS8
8eV8u2ZVzam9kRzX8i1dKD5p7jpblAsrIDIyqO0mJkwOH1EJZFZt5wyvrJT/msag
YULwGRME7icg4vXK0xDKowyd74n5Tz9dWiR8moI7tRPNXEK/kn8BNKNOc35YrjvK
Fb1KFXU1gDk+keDIW5pltzA512nxFLkkbvclBQ4pExPpAku+9hF2wqBoWr11brDp
gxM5sT/8zjL9EwA8WHn9S72xAhoNbbpcq8/k2I9Z2H084g25pJZWhy3Xy8EXIvGx
9GdvvHe9dRntNYUP+Vb84hw6ubyoCbLVvzGU+ljBkIV3epkAp0I0zOf4MdybxZ+O
Gt9RKXTU2vH3GFOSBQCGdpTiJS0VLd3FX0Vnktmb2hFkE5NgewdDhlICv0K0jfPS
U979/NbU/Y3aLG1wiSJaxrE9o2ZrfxaQypv64OngTbqSXQeGDEfibr5WkpupN87s
jLBkKF1kl98gnH2MIkFjcuxX8wLL6rG76U5k97kVk/l7GWD37J170nvgzWD+K9eC
lgobKareTpQ0bYHapprktaqUvF7oE4j8NQz9QrpaaDLQHinF0E104nRhm2Tm2eUG
t+oai58TTY3nLk58uMV9HN4OSmNJHtqK0woTGaf8n+9zzzwOm6XH3CxBQuo4NyBy
9rZJtk/3Md+r2CWWUFb6cAzWq1krWnw/0MyBanzHZNf2q2G0WDYC82kMtzsKBkBZ
SwUu12n19LxS3kGF25kgfRMONX3R4qFJqeWBr6mQyKRlpefM9r5mDwCIKDrL7Ekr
hOWnRcjJ6reHPh8HHcXxCOlO2dW98GFV7pr3SoicUvwakIHGHYOCK7qtZTpnSwt3
DwUOmQzlVH7sXWj2blDnGUf46rTzLj8VMvnKef4bvsZXBz5ekmiu/eVRIb2Q8Bba
fslAIeUFqDaHDT5UCMDVu9FK73VyeXHUxDeIJLzwFDisXhHoxmYJ4zPsYN+gtlbX
7yZH0T8dwyFzYcwuHw11KymBH/NBkPuulzyiAAA/+pHiWscrh+86tVDcawq7OiZN
H/+iSgZeEGmTkeNonO/VaygQxtK/mK88BnabKnltkreEhHBuDb3D5oO4z1Efbo9S
8h2cMRjxY7o2bfDcR4/31zyEOQtExwdqz0O5ODDWRzP8USBL1IBUTPvGfI75od1M
Vt/zQUG9ELclYGGPRc08JkSX+NGxUJt3RP8IN60Ib7332qpjHsSMtVc3OCAE6N3g
GKHZWBKY14J8a0KJBpd9PIBMem7klObuoyDG4OddF0Rr5Z9onw1J3OaeHYEa6OX1
qjWXN25KI33C+yC9uny4ls7QzvW40jiHKzi2wzkmOdikMWOk9SzuTXnrYn8S3DNB
wemt+GrFtdmLI503AOR1sCQEXcKvwsPaG9a5yxHwW0Xuow1eh+gUHEVMgtmqKjLY
eyEmVeHnTfuhWGYfwoLjExwg895LsuPpihv71WxTEHTOhB+pWdHUTd8awkCkA4lK
xupiRy3YrOgIezwGOd2vSWrWG+ai+jlQD5LpZ1T/WBExwKbR+u3v2KCLQogHzgTh
PGFovkRXJSgAp5l065MbvDaEelKl36IIjXTyg719ahS4FjBhK0Hz3udUSenxQ5zO
/3n8OelErspD7bMM8N4nA6AOld+uDvJxUeDhkvaaFatoqMulYFkDA+wbJ3rc2q77
8R/knGtYVUMre6TWt5XiMRBAmJT/5siIWSWsgq4WLg90zGek/Q9ok+qfdOaWU5zM
m1xscp9W496Xcj7FmL7/eySynkCdnHdXTf3PE84LIzXb0kQxUmAChtGHAO/pddiM
J2Aj/x6RqePwBNb2OCNp/0d+4w4NNEkakonx9s/e0tfsnOtAsVvB3ORIRfAa3CcO
dth/n8BRrRPNh1m/ShZrXM788xB2UYu839geu3O/M6OF6o4k4Vcdz0IiRHI1sD0U
Cb5jqlIy5m3t9GNjBbbEPXhGnfJBuamnvdeFSpakTllZXz/M1Ba1k3qCVqearrbX
U17ZVieD2VbIBCQcnLDh9irDqwfeTIsjJ6VRDnqQDn4TbBXkj923Mtv68pl9vBt4
SpcZk56bWLgF2Y7mEOtPB9tmgpvLf0AFcsZ9wGE70dvt0BNfeSc7BJ2Tfrh9RNYj
KKKXoJz1KkkIkfyinRwJdvOKq/QkUWEAimhE5LubSOT6NAAdrM1jOBG1uwaB6EAu
xR5dojH7pzwsv3R87Zl6Tm2nxRReuGCyxbBghPDWn4rkFoNxTW80+HrDVXqbnFF4
aIsKnqVlhqd+vU8+O5N+STgX/9lfZuO2WJi3HWZgR0kSsITe8M0rg5Znyt79j/44
BkgXbz9rKDzZedgra+dJxzydeDsyCBdLrY/3VLJK2m1l2Zg8j1kxUhgF87pK66Ja
tLtuHRzCcMfOSWXRlcyuVGqir99fqW8PNcEiABcvVNQnXvEZbyj9FSMd2gM9bfAA
67G8lIl5AwLdyARlZ6hZ2nr53PtK34FgDoXTjKiGWcafddqdcaCz0KbJwtF8SaFs
zYcyf9Y1+TpIveU046bxPGN4LGHlWdud/VBdM7TdSuOLVUi/CUidMEhLxhI1k4ZA
JboaXZMaCmHDxZa79a6FsRfhQWDFT9hnPbz8pK8/gv8o/BZdPNoboPPchZnl0BoL
6X6y0xi4E9UQdUk6B3vSaDpG4DuzGVX/soEf0Y2TFg9vnywPKbVI5B6wZhJJyepQ
tx0wTEjn6dhcEDeBjy2yPv6TIU6NzaCGTbPtPByOUsN6+8t/ymSmJFgUQ+6p/qIc
1/w0gBjMrOqrx60iTX+Z0tWu/Yhq3LOJV5jrD5ZSA8S+4m05/ZqYNhieqEdslEQx
JU6zpYvJDPmw8NrL1JknrXSKEmCk6944Ou1/2PkGFXrQbEdZfLq1dBr48tIVqri/
SAUQmLUeyIwDrZ+0YwhhARozDuoRamjeL5EtGo1wpN5LofrKIFz198czBXvSfhXY
gJOceigdGvOla8M8vhNx/iCUPgG/B+751R9uj19EbBVC6mG52JT6VK6I59REr9Rm
boprWEcCJ+Njbyy2RtQqGgKCUWyHUer5dm/Fk72J/JWnukCdFDqr+GP3CI1wJUT+
5qyXvuNOdIb9tMOQG//e6qacPIH3HPNnj71sJJ9pLV+2WYahNTa3Ble3wa+Y/Tt/
04ALPHkwGpacOESLiVChYAFZnnbRcr5MpN6w3lFQ6m0Wa3h4fKI8PYSfFCtFpnVS
0gpToAF8wmRcB0guBQ9Qo91ibIXEFeu100WABBg7zVZZENjvs+W8oqXgjaF01RJ/
wZBaoR66N89eI3zQT8S+STb62Ly6B10XsEHazKphigip/qXd6fDDkwxBfpOz9Ftd
brwZld0QakIVGaeh6LbPvB7kR4jwq3RZ1t1666R+PQDleC8vPqE1QZ94CoFBHoDJ
aFW/SWw/pOERhKKuwWn3PC9cLzndZ1oH2p9z3nSwnBXfqc9MMT/Jes6ImeLyRhZa
ru8XsvHvdsHdNLSsQq+qBifRvqkB5U/Kbg/gEzA9vfMNU0uuuZC4mlNztKhcX56R
JMleSHxxx83sOdMsUo+0kRNq1JM16gTDKRf/CgDECx4rfHzhsFm2afPCEklnrTof
YGKyjhZaLFfuPWB15e/MigVrN6hCxZug8K2FgwXJBXmEFf6hyFnVPk6iSbFZOTqO
YUKtmAtJ/Dhq+wyGT53/n7vbnuzy1GGzyrtzJneY3orNxdK06dq0G2WLyH3rERM5
Qu40UIVQ0JlKon7172M8x1tuTidLbMgub1T2njgUWiWqfs2uzzs37t1DkGPywARM
tRZRj7lE6h3kT8s/5abtZkc0DP99aGIjI4BPLoepWxb6s7jz2045cX3xNsJQCPHI
TGKvlqxBXIx0jeWaXMe7ApgB2wY1hAli9yJPkODUrg1tpaRj41hr5hJlrfFxz50g
2sqGs/Kc6wEdYJpgdUn3htcrPlEieKGzQzOZGn4DO3LnFCrWMINnCLQyVMz8womi
SPUo0Toz76spJuttawz1ESrZamYhM2v5Nbk//r4HGf6A5890jeEEyTgTCnUDz5Re
deibtOx5ta9woAkr0M+Z0GNFxXowKQ0D523pxXP1T8YdftoN9ATQmrR13OGXMQ+i
1k9/AuPcI21/iHU0FVWmkKVvwLe0HlShouKgb5LvEmzYn2caKT3kRjnafLiZXUEr
wWQszAK/pchWN2D/wQPn5V7+VQtKtjFGx2Mm2/8hXkfoxIQEssmReuXyTwE3NNap
BIwO5WcCRoutR3CHrWX5G+Wqb/CCcZq/IS5lwp0XYZndkTZ+222XqqzeNY2kwgOf
Zn6jklOmcWirnjhu41QMdt0hkeqZp4MrSa1p286xM7wNori+A1HMAJpYbglzOn9S
86eye9WpI0E4b8GRIz3BLNkmzM6RhqqY3iyrjZqM2t1OusP/q4Iaiw1s7mZ3tc9+
dweOjXJX7ZghljB00TesuPNFus83eVJVyOFkYAninc7RfxBYYNlETk+YAivSWrOc
ETkARUaTqo2r1oEeqa4OcrDHDbBsTqs3OM3KgmTFqUW4Ws6pJJ/A4WFuJ8Cl1MRr
sjMSDcy9Ge9w4zfiWzN8LbNxs5ZBIjSZBvapfNQ6hf33sCzlLfQ7JUhwr16H0agq
OysOYN6o9+oUhBfcA3TywNDFG0N2vTbYbs3eQOwzElHbe5kPIOx6kARnrJ/zTOFy
VqrR0jcCO66MV7zIuqaUFutKYQ+/A3Gnymjbi6dcUs5uLpbYECYKkpceZZGcULU5
ChU7oc5XuUjUfXxql2vn+lTrbp7Pcvq17vDinoy0jGr4OmDGOYltph5K6HZLR/MX
8BGM6tWN2owwahoOkiJI2ms37ZKfVGfJIqwTW79Oswgxc8ErdXQzMME65z2EDRAV
4AMIB4x8aAwLXlTO/l9T7Q0pY64HICsJVSPZSNnosk1J+E/E7JIs2UOHK5FY1e5q
HVoXd80hIkPO3w839W0JyRM+UeYcktDkfAagA6g1Ronpp9255EY75UoSnRAVHdLk
AxaymVLVCrL83JV+HGTT4Yuuomgzplz1eTGFAhs6ED4H4DU//IhRHoUJT7/SWRPS
j/4zirlz4IirLyorRTSLoQCOTBK+67sElySeIBSOwMyDMJxtA0KaXBU/h3eKYAXg
b+Pf4zaPEt5ynpcO41zVjLpI/kXTh7qwvDAo8h3DLENFbE8+4mPgMaMJsNk1JdTh
qn7oZYP6D9N3NQYyD3ZJ3SFtTAVc/eRrNO/0uyXem9UGqvGsKLB9nRCFPgobBQuU
OqIPS9o24/0YYC84NdjNAWf8iq0Bfx6IsqDPLuL1j+aDbJE4OoXJpJ1lpnkhRK9B
P/B7CS9HEOn6l2zLRYntSHhXxVjV5Tv4R8OrrU7LEreA4m5XK5JgtKbcb8MpFF2a
jledpJKl0Yc2jL4VO7qEuKlwaq63cvQRXizbdLai2C58B+iqNIKMwe7/Sf5Z9Z12
NjnUJ/nUUSunm29j82JETsRu+afu8/Et+YomWpDPApPSBBfncROSWCGMcP5mR2Af
PP6Vr6Hk+84C+DSPXCdQHWs5+SJ6gqWvBPnETZPfsdAKkf9nY1T/wZxjl0O4Io3Z
VJx7Or1j7vj72dD7kg/yvnrJQVFbrAYSnXqOC6f12KZqwawg056VAug96G2LmzCb
YqUosyibtkOItcNPPjxMNMMpOnd0oev9j53NfrE5x7uWVUZZrHAGu9ih6tpQJXNL
P6j1Hu6J4VmiwDzn2qT36wqX6UQArPEVoe0ayuFErUADfzVtL4fX/87z9gT31+Tz
pksmyIusBQ/A4TtkmGC3QTSxHovwb9WtBUxYLTt5pNHczjjgejFoTXsd0KSvjFvK
qc+JR6iyAmxZBXifl7bcm7c3nolTdXewtHiYpTH7Gf63CjAVMxiUzH4iJjbNUb/G
USup4i7WrDHcrskv/D8oKsGTV9vUA3lc+jwU+o+LoAyoaaBeHhLj0AJb/7dzUnp5
jr5FdZZLNdIHYM5gKCGF4jdBt9X9vqizVKJPhA137FQNWuOMdFyD2gVHTr2EwfvS
rKS4hpoQu2vSJzsO8gQ4qBtis9YgfpwHe7vbHDpogT7iws3BYTJV0U828ikRuYf7
SvdgL8YAakDr199DmLryBqkJMWPOM4hbmvvsFZuQISNgxwaDjiuMLsu2BlYNdcNy
ml3/83d2U9B+Ilbj0+n+kIQQ3AehK75AHulZeBlVygaw9sGeCGtb8y0vTzRnkh7y
qjKZVBuQ//vP79odXSaUXQWinjVjUdck/KIpIIEM2MfAbeXvLVqxCYov8PPOgKaJ
g/50WBLEtcvCBplyvv1AqC8WUrK7n8e4nZVcGhN2QzgZPt1ZjA7ef/cAjAAM6DMX
JaAPmvpGvgrAJHWJ+Gga6xBxVsR818Mqs14mXaVeKNIKwiVWv4A8arFDZZd0iH0a
KxhHE8UVvPZmTckcbxm8IrqHnqeNDdikSnrGk8Yd+4HbHc3j6gSiKq2x7x5s5Lmj
WSXeF0EwsyCX1ggmWCB+m1Xj1x+2zbd3JBZWAT7HuZn/lWLqEsKJLP93IlAT7E3/
kMuks++vToo0J9P4LprgJ/zr1J6zD47TNNfC7VybRY1F9ibn+wS1oJu2c5xaynWa
M7YYiBly5eDZXzKeAMdu65EN/eAx2plrmMOZ/W6u1skfX84WAVDBZrbzoXtp7KJ3
rIRwZkGkd0zynPMEyVUJoaJoYlMBTHKU/ktw095PuUUWtrc9jTuq9NfMk0SKG8AE
1fgJIS0RekxaWpdIJzhld82kcaBFSPxV7YhyC121CEIaIFD+eU3sBT7NtKshqsbQ
GPC9aDUGVbpx9ejvLX+efFrUM9mIBqPVwVurVmwF8taCkEFCfqWDJJ9plJrDnHrp
TyDUeBdzKucRAgae5aGq2lSFT9lIAkf2yJHPkdIUzk2VQdcgs4bpyXEEvaSb3hiC
Rm6RUTo/rMsKwj0TVzurKAJ/qpoDTw2IEilSILOk5+07aSWTOxNdBDh0ytg971hb
//+wrJwgXDC7jpLj00jgXsWeZgS6BVuqlokFKoeDEmcOxm2XP/ZdJR2SKnG5pDtX
UV/3VNzc6LTEg+T19PrzsoKJscYvc7pdPNyljY73ryrBmgF4QzRAsjLtr8DLpiyv
GI8FNDCd3m7i4dHomsM/qI34nt7y8N4A1nvpTy3IOUArVhVQUJfsMGqhx53suwUD
rW+e4LPYDHNRsJ0mfS78K1Hv59dNjmfQxWcHCF0R/d8Z/ZRWNQp1IJ0lZtQO/7uC
NKuqLAyalsh/PuqQV3Dw3bki29t7L9C376eqx/hhzbrjTvtodql1A4CPcbz97c8e
dPMeGrh/47l/Qn9lqSFRtZvhs1peasP0QTLBb/QfJ0hwLGZ3/ghd7elEIyBZwXU6
zXwhaMJXpqWUozsNVlShRosl4c59QJYXIm6FlcXTuto01mSpGi4MoLFi46bJNnQg
H2eo3cB2A14toIeYgh24KyV+jgRGnuhwdIBIdVB64IlnGLPqgnyOclcBlF06XHvv
tCgzdBfDSuP5F3XBvB87OjaC4MZGExUWp2K9+1d6451Ob+qKdULxfIigA+VWRPHQ
5v+j/jrW6lsyHh3zJnooMM8xsKzerPiqJdHMvqrXQWqM8bsJYLCH39yNSbomQWwd
MHeWvrbRl/kzEMwFinRaw0Og+gpk6PEwpf6J+y90lJYGARwuPevaVs3j/4a2VORO
XzFbIgams9+Q2oWJ3D1zHECuD3YLX/uGh+12N3u3pqhWAFz9Ay1MFVc1UHBBGROF
rC4PKv2MHOv9CpwydQB3+cud2nfvE/nts5+w0s/IbEpFgPDWKY+T/11ap7de0Xuh
y03ZdXdzutbdGRMaWJgMcNXXJAlC1kEblkBB+6eL4VuSNT+dxwvZC62sZxQNV4di
Ufm0SPNkmljSmkPhfhQH+UK+Z0M5gkNt9J0S+dLpGylpnGPEAO9Ku66V7eyQvsAz
ZtUSKLWk0NpRnhO/Q5F1+UXA1s2aJCoTm1Yfu4ycdmktdocaW5UsTk8Eo+ywM9QN
2wtZIDjR2wB7lmIFP0h5A+iw7O34MlY82Xg7Pri9aCnbiNSTnkMIxr/9sBWICDXn
VjVbdpJfS1occ9dYt68AlkC7HUlAPc5zAOlzWW9I9IK2a24k65/qnIjA4a5CaaLC
5SG5RvRTVmyKNH+Vtsohmpy4u8CW5V1vTViMngUEcrgwA3xL4yLUtQIfbxb9sBbn
dEhPZRpUcPtnm05/Ct1jJ72WFDA0rFIZQgxjUaWOdN/Dn3+wg+H1dhSFtCJ+aMJz
Xrtq/BKfG6AgQOT2iHXtppj13i3cQVedG4jBMPo2VHEHGcebA6d+yYgHTwu/wZ/o
O2ObNF6lzf2EVdsHqV6gq0Kgnql+SCunglVT/ZRzLIJqTpwAJFiXT1FR5fK3oxHR
PVrYbSwktg1QIwzEzkftINcnrNV4YoIYKCvEIYXeTTj5sOgHaA6r4vPm7ikgqO8x
oVSskVZDFWITjrH18OFMHaixO0PjRuMrzEypK2E48FLEg0+i/KELQB37QaWDEC8m
GGyAXv2/WgBw7/vo2TccAGgRox8Q8QJ7OlMAfoBSOoOcKi6TqmJe1vj83uzKmyqp
tDANlRA695p950n30ZZ81yZEF2secM+OP8ek+y0UqZxIEKWQ83brtWwoiK3K8H8r
EmT5Q3PESEnt+tO7RilEp1mShkWgmmPV0vKyxMvRtZUMegennjl0uIqa9UnBGoIy
wkMXnTm3nLyEjQwMqeI+FGYp+Im3q8+RDRNYByTXk7Q9s4WNc/iWtbEk/h8n8jDS
hEdzXO+CLIS5DRq52GIOEuF8OYEdjaz8Pp0BeeFpkgKCcFLKSYTuTKK9eu9ERoFq
d/ynKJlEt0al7wHRwm8k1kx6MQLud0b26ZWAQ4tIYUBvMorHNd8TNYjz/NohL8SE
3eyQ5UdAE56To/54vYQrgvzlBo9miG4zYBaNm41m2rQv4GDKch/bwlDGCdgN7FS9
v8jxsqjhqsbxunUOgVZdegTY0cr3nlnQFGD9Nvv3K2K2Vq9DqZrHxszAsjoEFl7h
2I+SP+Vq5z0bwMa1uTpfWke+qdp/CtPZ2xkzD09TiusaHXqHQFrW7vMZsBWu0wQt
csY1uAVsqWHNjN7zQPhUcTCaxVoH+DyQI38LensRB3ixZGjHIhuE0N85KEThQox1
gA4/BaNTbVV02jfJYwdHI7F2UdYxzSd+FPHga+4eAGV/Q/kdijatpeQqNzT3GaNf
VurBRLP3ok/DzR2v71Ah+u9K4HqHBeuQvjKpCaEsH+qphvhRUd3s1xeZqEvJQiQC
90nRzm1+O5zY8ULA84b+Q60e85ebTxqpGurrqKTTVvF8r0H2eqNioeK+GZWzn4N2
5BZ9z+V9Q/TbsYv7o+Ldk4xMfB843nJeTnhZzIddPhxlre2vYOnotJuWaxjdezXl
7aFM7kHpg0BS6o+7uQzHFP8uBiBKenrkNc8P+jPzlW6v+FBRsiYkYtf9rK9IFKtQ
rS++GaYajgNSQcg3SSMFYaBlWzEtKMVApFBwWTMzGDb+IBFWfoZRl5B4hqI86Nui
jIkgIbvXipjgvFXMoHtzU09C3ZYGS/VbJnVWfJ3Qw/Dk7pjbKBBmdgSqFsvbVmLu
IhO7Rb8YbMTp9jT+t2VyFhCOr2i9iIXHM6ewXaFQk95GgQGKt042p0f12XiGNC5Z
6nrsxnXKJwD6ds8qkrWQzFg0qQJccxoMHzxVaBt4emyUAi37nPw7z4MshXBJY8r4
P7sVat6Jerht9YuFZh1rFyqr0CDNgrPBTy12PluvsPnLc0PJpFHZcj1PI8NnCewk
G3ZG2WxdatRMvZ7oBlQwC7wzoK1GGoqv1hwi5vJkHsAShs5eMCzWLTXqyz0OTNKd
hbHQibZRcwbw1QqlKo3ckkB5p3Sb8XVozAprrEkillhCwGc5NqqNlxA8ejiofCu6
qgjd4xC3G51deMZjTbr140hNnEr75LJjNIIPf/91h6uk52loYcs7A8oh6mwb1eTV
k+bSakdkQqn9eLR8UI4a0vb83cwTH1YZMq8C2J4RNGsIc8/G6pCnc/0bjHuu6ueY
0MQoIXcYz/eRJMEtnghcV7goM+HbC5n5bKuEPDYqnZbgzmLLgDboWW09OZjZ3/q9
6bLe4M18w0W0PLIFhMSM+dVYCG73+sTPsfcmC6JRTJbQs1aKuhpnneSDXT4vN8Y2
UeN+0P/P3sxM07XDAYwbPrBXfMtHcaSYkJfh+TKIP7HBOqn51cusa8bMKa28pLLC
faZiDJkxZSaoRcvJLXRCvNMdHabHd9KckJdzKPn6urttTGupD0DUZMzwPgh2ZcU3
uJU1Z222+nIpKKbMZpwTP/nEZyDmnT3S4btn/jua8TJOn3s94uSvajW1dHfuWvFq
0yuZOyb6LbGA0AfD56Rkf9VDiL3v6KPcDJIMqgw7gBhJR5v0aNJCj5du1Ce2z48Y
gQ9DUUnJhmqUeoFGjt8n22VsJSRavwJ9LUsaicSaZb95bpPozqsXGRleYOttHJxm
Ldw4iJtO1le03Dq5ZOX4XRAwkc+FLmUJn+qhrHhGmUYpq7fmRG3gUhVFqYaZ9UWw
SezA9HMEP1WgHzd7XA7LcKgelBvOZWMniDMXNo6vjtejzrRVfKbuoROvcT9X74gC
/sikIRydALwwGJGKNnDDNUwqM0rBXyVK36CfQjW9qoYg10sQsgzpb9S4SBYk1RZg
+k7fq3owZSEXwQFDVKKsMRKrFjovV4RdwUS4ukqfHRVkzEgNtZGySzz46W7meQis
n2X6hUPZ/OpzASBVjrhGYRTgHaAB/TsTTSRIY8b/i5HSdYYaazpn9LZIiK2KxMxF
oAMwG75BGpP9KjoMq6Er3j3yyFzjHTV5Zrw9SX58xbLPMuwqf00Iw18Q1f03cWqI
jT2zC/1k0NpIJkcaWPefIf1Jnna967cbiUpOnqGt/XzSO+3Ecy1ZfzMc+t37pp/c
pwGJzqnkPCo4v5uLlOca9nea/ylPjkTUbi40gaK2faf0+/Ct4YqW4E7GEMMGOgoO
2DZL6xogsjzmfQGwSlWOI0nHxggrCd2Tqqqt3ZIR1EGaidcFyfqPB5zOvG0AZDWH
Z3RYELcgOnTP76NLO37NPHAEJQmBwLg/OwbYmKMaZGBX/QXGg55stl5OaY94udfN
qjcXgrSv5B+BOr6A+JhEYvXdvrsZBkVH1MfvtO5X6wovAALvFVumfBjDjwjEqYG6
u8TIxW+HCbZCpXuYFGaOG//u351bw1HO3X9NXra/0bsXoMMHvz+rNsUtPdZjEXHC
z+eWblY4rv6sBF2MWgRiEyRSMsh/Pa1efb8oJZkjg+Ae+wbVBfz0vXDrKIzVbds1
eGFS1GITcSTHjrRJ/YX+miazmsyMnfYP2IqUr6Y9r64gc7weXIZaAL+S5Cp43e9g
+zRLD9PvhsmI/tnLN9EUhE7Sx+i7jf2yr0prcTzTnkqMWoS/FvXsXUfzBCmrfrBf
uJlnnq5q9IV2Suq5SOGlfpEtb9pXM/TfpqW3UResSPAHvRCShEmFsFor6z067VTQ
G4bEvQg24CjD7ggd22SfPKSRHVbvV2U/qcOXYg6H3mh1vJ9tU2ww34NNiQLK7/eS
NfptwYab99xhyLrU9Jh7yfXJMHYERVHGWjX+i/LftkZRHmKi6MB7qKTAez4AYPeN
HZLUi7lNnzpG78qg6QszIHMs+uPU2hj0vIq+3PrdWQBIWcr4vqhPYQG+vBCZ2MTL
rPulssyAQY5x1OfjtYNcfeKbs3iGzM1e6zADtvk4Rx3uwF+i2j6NQrMxkgPyoFyR
SCQ/9kWoWNUJjbaVgiuJmf72qBZ9f9/WZiF4l6chUNWZF+SpytC62UhSuYmxicRr
x+KT89Dvj0rBWnxEekI9s/hz41mt5pjbveqbYvxrJmnFg76LmZXA0/JhAgIqPYVo
kUgudZT13tbImFidkeYXHvxQYhuBpgbxTPbgbxHIcjfuuXG8UhgaLIVbT6U3sJBP
algX3QR3wVpAD8usxxoFOJS5GattQgbGs+C+ZPl613DQMEVzZCXo6iTpz5OJWbRX
eMa29i8IGvPzuAc2AwuhiBSq0g2Ovfp0yr0DpzQREXMSthVBA416qs7VnUpFRQ6c
6Xwjb1swtqgJEEXSC9cyPZ8lrE+yZlCc1Y7Ddbj/BSyeWkrDe8dIlXsdWSzfHrDu
iTNs/lo9GImXD7ESMYI4WeZLoXDYxWueFCFbMTpUI93aFTEz44Qurk2fPoFGTxVO
7WKjxyPu+Esouf6BqXUQyut+5xCg1X4qbD1A2566D+3CBC/hw6k6BHVFs4DWFmrf
SNixtmUd65c063InFdlDlecVDgytuPW6HuzANfDyLaw/akq/xABs2BabTviIIZBR
lRXpbPZE91HYpBFv/2baE6uauziEVBsPzaU1povJXSeMEFjT1aynmhS5ODchpL2m
9ZJx+D7BVbD3Hdnbk35aCzCRH9bKS5RTqp3ola4vAff0r3hagPJUaAj70/xEMxYo
ylpBZaTYy2VaFz/F5QQIxt+cDus6IgkSYoSiFs9P00jIqxNsCOBg/e+fQ+WOi8b3
qyrkXE5sMetrAt1ezYYUHbteUw0tpRiCy3we8k5QNnyPA7qKYITqHRxsbQHI1nfa
w3z+CWmMplAimB4z5Lilc98/z7k1xBi2CJRe1kD59ZvEoPcpPOR4akgAnx2l3wzv
HiallJ1ntxg0ZtZqyqKG5MNhClcSM4EqNQkYRQxBqzLgjCi0x1PRdtVV0LEyTo/n
lLwcK1vTFWJvehD+7nMrnrOY2TvxYqW1OhDh9nGf7hXDPajPRqUQ05yq2yfKek27
040AJ+KmUZqM9Gp/2bQLnn2/pq7N5iF/d7lSH12Ozlo6kC4wXwEOdz9rUebvGBJ4
FMz8Vqim/rog0JWQ8ifDqPApCMS0VnOUayf/m4tlrFp4Ryr1iGuc0AgS5She34db
AZfiVsKN2E0LBobH/H/3raxclybRtFlXoNde/yFEhgO8rOOAH7yTbQsOUIkCp9I0
9p+VGrJTs+a9ucvS9ioxKo7phVe3KjM+AIdPSjH4WAB64BwBE2inzaWNMPI8knYc
9FKH2Clr+Z1BmyRcuMwyrNp+Fna4PE3lpATJGFSkgFsjYcsBeS3+dOCTNQQarVG4
NXDcGKG04eGxBI/RUyq6AfQjxEuZxa0/25nc8XIrQWG9TZYCbtFygwNN/osQMyoN
qtKi5sU1H2ioORfz4CkjIxt+0TCpyh1WPuVIU9gMNqZG3FIQMC+8zfjVzOB9thkG
whepsRCCcK22t6mdjrrrPrgBg/BKF2MhbQ1ewhvHAgxgEo4ZxgWo8cRObcyhjLpp
4OIvMepYu3yHKiLqwPildHicS2k2++3vSFOoRFQ8vClWhK/yJjZsmbzItacQ36Ud
2WukVtaMLWCzMleAlUm/UOtaMZzllXbKgx3ba6Wut+JLy64iwO3N95ihBqH7nXUg
bBulBHVTJ5AACNTc/+dFZ+2E4GCBDGH1I5agRkt6G1gxMhUtY+FnuqhSDFyG/8M0
IRD7cRLABkEk0uTzSUKY3ZChLk6K3AbA461ITmyYeHJjCc8fcfYVtevL8Akeog9Q
psxiENf6Qr8cpf+sxPuoDiD3sZz8HCy43snv2gMUxziuYRk2Ch4023T9jHLmhSDR
hV1shMtrwqqVi/GncJ86EU8Mz/B8BIqU4Px0IXpm4zZyhOhk7+8igOTBhq30tqes
3AqplSA4zBLoLPGSkbt2vp1L2ijCOX0yLgEMt/5gLsvK92ZORlmeBTpU3ExR4HRY
BibRgYgxOrM2+qovtjvWD3kFXDzA9XA4dXVIkFNfoo77TJqE8Wd/ACEjtROtRHaW
gVX7csRmGWbyNo3ErzRGV7UsuHzQLB/lUr2tB0B4gYCtPF5zYTRwPbAJfjVZLajE
BAMEKGkLBlVAeiqq0m5SlAeayIRq1ABsozEmqKH8eOUwk0rTNuD6NoLQ1Zq4j4h1
H/O4REEafyErhZ0Poiqzj7+vDAkltg27frx4jqZhwfZktyMgKjz3K2JOVGRqL1Ev
8LelieTCu341HElaOJ+gNJM2UNyoomGAywg2K0Hpx9n0wigcP5KbcgJfy/6sWO97
GoHROAHCc0aVVvR9qfLd1li5wCYZt57ltuXl8lpGHjvaJW5dIPH/bDqJH/4EXc9P
WSzjndx4Cu9zQGR/JU1D6QmtdenaWHdPgiX4Tn0xgX1kun5ahom3fBGjxQT5cCxI
PVJd9oy+6BOeSuMdyk7//Z1OeFt9pI5+kZntdbmAi/OtZYizbJA2OzZTBe+GUQ7x
T+h0iusUM+bjw3BenpiMEbLr3ZcBwy/efsNNL1Xz8/VSSWXYmMcuFIu9HVPF+PxU
acWvVmF1+xJ1JhduVRpxrN2ZGKXtK7qFSPcKjUt7AWgIQCivxOLyY2bGUWHSva5/
lyLNKkWS0Zl4AaFC2Fquw77iGVxCEefaGyOfsBa72eVPYvXkavkXAdK4FNtVcKQG
WxctLKSx+9HYtV4f0aE6AaWmXmZRjjz7EObsrntXcbwfGI7s7UUMnBQrbEMzWj1k
vK41iX7QksRVTf27wMWGq/dnUJC3WC/r0+zyRR0v4J7Ajdj6W5EdAntJp6s49nip
THoYv3kmUrAnFi6iuSupslZVMaiybYj1jzMX+coxCOLF97pkZ4iQHIY+vVOwAiCN
w7y8BHVUjeP0dTHA1A7x7KlEMt28O18hSx38454Vko161dAyARGiEbNnTaqc2/mp
eVrXsG1myV0t0fjgOlXRk6u//Io2KzJhuh5O+gBwway9HN/xTGFC5JE/7dopgAgT
qUWgMImcGAM43+RhlkslQtAsvjPwx2A6zuakuCq4p3JhJo2BknpIbhgAKXB7FoOE
c6Oa1+16gJwQVfvGg5n01FBNM70GJApqY1qsKqO3aYMLJBBs8D6l5ZwmahEna6Ns
DxEG46CMJ4RQO4gzPIagHrXUMQYZAHuK0XVyyzyjYiDQ9MNVjI4p5VMuKBB8Dp3U
p3PjWUF73D8q9hb9BAGG8tqPfEAuYuTwUY0FD1abb/sAsbX3lAUE1SxzvsfhpIv7
rU8jiu8OK+cYBxHYvl8OyjoGpUJVDSn6f5f2DxaC8tabPmeEOs/ct1yHU7AHretf
d4yUSvex0lLO99kOs4MGrqVSshnfEwcQZheVk0JUVxmorcKA1MmiYy7g0dhEJ75a
3wulqP5KVs4fsLAl7xPGuXy2hA0XuzfUHMSJFI66Oi3xF1LVwk4DN7Wv4sPUf7m6
gDWdQrllUF0YPTA1LO0Wazu3UkWkgAFeYADhAAtF2KQxSkujj7YTxZlUl27dqANJ
gi+SKIrmDPC+Nhek6ZabEB3lAo4qfBZVxQdA9Kr8T+5pfDyJwkOzjBp/dy52nZoE
+L1UHq6wrLjmbmIqR1I8GUYYHM742pg+cW/sCVkDDmx/Ps5C1em4bTaOkUy0+w63
gXt2Wv3XhJQI69vEl4ACoh5c+qM3r0sXBzk4I3KVX3U6iuOg3jMO17maMDcz7ti0
7V5ypsC6GWOMfeYRY8xTqhonAs/9p6ZvJ7jqxvsktHql1fK0ZEcYrQbsqpNkT4zX
7vYQ4l87uJxmVb3qecqhini6uUn0e14um7iTk0UjIlIIuuN1f2P2YOdXKErSwfW1
MHHBWOX8RTpnE9wlxgEeApzFDQQ/upnL7YznlYGlM09uO5I1CZ+5Lmbj0IU3hBmj
ysjnmysN5T29Lw9YMiqa5WfgfQd9hgU+Us876dIJx8tV2nw/ypAugu9l3vxTo8gj
wOg/z6aIERdiPKT9jdJ761U2zGZ3siLFFH/Vosu5kHgSDTNUBwUm8xyrKf5zO/HV
Ze3A5gqhvr4p6eR0Oox5iDPKXAyhBF1ndhY+DKW9cj3ENPhcCuIJ3Mvgt0qE9DGL
cTDntoZvf5M+UkN81EFi/di1aPujS9utY6nbks7+yseyPk4dw7ew2kR5dJc4c5zr
vzi3tVCWYsfAAtOcV8aGsgo4mYutfYoct70SKpIlUOLzr6vTowQF7I/prJS2fd1G
7LdMq+wR0UGEEyNZmhsDaAE5P5ZQDefLmYWuEqr71/v9B6oe4Hi/WwPyrKpaYtNg
zN0iRtlJt2K3jjyXwt6OPjhyg2VNW51QjkKFPbWH6dl27QUQUnuWYgsHYhNXEM9x
9Q6pDttfBltEe3d9Q9MfgNT1qrlRqS0dh2BufdMXaT5hkNwdrLcKChcrxgShZ1am
Jny2BOWDrFeAY4z3xXNMldzY/57gekcr/BtM9xlV++vhRMZNNIslIyWWFIC2E7xw
VflBnBB1mjnTRDocd4CyiHkGyIyA4oeundmQHEML64JQW95gLX0ASJHAlUhUG7jx
Kmr8UvZP4197hNlQAamYRxIIDeH26rW/ZCE2bqvsqPK/bZurZFVxc00mFbJ9ropb
2gi5+mi8Yd1xV1v2W4xQGUc2ZQscAKZF9HPOns/b0AC0nJV1gslVB86HKcoMDhFC
Tx9mEGCGeEYAXDQXhttkFRTT1DHQZeAuE6BKygCIRIO68knwv6V+cJ5yAEBVhQsv
vOoOIAX718guYYmZym+GTBZ3eOKQ6LejeKYqgv3S/pG+V/VtW6R9WFlLxHqJNpXA
t1voSR+qRtucrLfij1tlTPf6p/7YtdSspN/Iq8AiAsDnx4qNRlU65uwiO0q9mTac
xCJrxA4NUf7+GQ/bgy+mp+gBKjYAppX41a4LgOKDsnbLmeN9gmio+1YK3wyjJI5M
MMX3NV2x70cQJ6YKtInGNzaSlJEisycUDjC99RyUCg79SVhj8unRIBiWjpjKRyNE
RoDhAkLvQoe8/KUyrsszk4Tc6OKp6+NVlTndpCeS8oa7f6p3sdYHjZISfEAGywCg
wg5yNMOp1AueyQ7I4h3Gq5arKoA1qP3IyOIhzDQipupck7IGpKaJJT3VpeXObCGH
ENHq6Qv2gQizIzlROFpNm+R2jCexxLvFSP/ABTMEZu2Q+UdUmAcYNFuutZ6ab0c/
xmruJHxkTqRIj+8HekcxYasgR+/A2WLXu2WG2zgutnRQ00yiMfJ786blDhm929Q1
AcHaj3LmNr0iV8aEpO1+bYXTyFsOXn6FGrWGb1QP+lqP0nKC0a3vH7dcYD5KS6xd
kzdfg9mIY0BXw/AAjdW6DsNJAAsHZN6aI8M7Edm7IlIEhhgfcWMSlQlhyU24tqbe
MaZtCeuq6ksKHRKhpyl2U2Wlpr6I/X4zeH/i70cy3PAQotz+N7bNZ4sCxqTrzTTt
ViVT/r8oDVdxCrXJbU3CniqFIDpbLGIigozh+mb6bdLj2+jFqxSDbNK21WDdQbIW
gZ9qhzjLf/Y09+ds/mtt+BDDHkZzBCmeLUMaNqMSFu0dzSiSJf2bpZ2ZZtcxcTBw
yNjv/p99zBFVb0YSxnfEM4/z9anlgtNtEqk6UqSlKH44XH55sRfQ4GdU1iv2MhOg
XvuNkWoN1OUzTRtZVqByXHgrTyv0fDGT6QiMe93Mk+bsHDMj/uVkf88HzJGtdxr3
k4/GRE/wvTc5u4Lt58AO+DnUJkWL6MuVwupFa0bS02YS3aelcqNIAmJVRtpsNw7v
iEU5KrlB37wtlzrpCShL0juItea3mRVvYVFbJ09ud5nBFcVbTzk6zxYTsNYSxgmQ
YF1NHfQ6/xnwy/EKyXte+eX9trqEGlKnIgyfejDJCd9jtcWpJwCRyv9C/F9pgO3Q
KzInMI3QQXhn2kTSEfFXwEzv8aTAx8f4ra6osvfho2Dmo6VE2mljR+bx27TbBLET
FOELnsB5rJ5bPBp9UtYf2AwooZm8JFVZD16SYpjexJU/4yDEzbtaBbl8eeSxxCUO
O1d0okG+8/s5tmLWfu1ecxFS5ZXR/JQvLW9fyVuky7zX1WD8oWrC9+1+N22vWTUq
UhSZNQv7bjXIiEduLQGyBXzCFU/nIPQNMsCMgmenOxmk+1eFagbmpQ/KK7LCxDaT
OPbCcC/tRciyCk0m1+NPHWxBKfo44EHOGQN/RVo+I6CCLqizfsX6rv1wA1/NKnmD
jS+FZz5sVCVi5TF6M0x/McTuvlEMNrKCBr1kzIZl5Hi/owhFJYc7BsDlkW9YamVC
0+8njNW5bdYQU6r3P0LwcO27GD8XA3ducoWCO0QlxZeC+BoyqQc8tGM2FNHz/NDE
U7qTn23ifVa2aZrMlqxw8dfNTTBNO//G84/R/ripraT5t13yRCkrl2PcBIehCIbB
czI7AKYoN+pq1U031sb9hMIbl/QxHEHLeDwXJTO+kl+bLbpXKL3xPRzyEhhedock
Tl7AxxJ3LFSu9vaTkhLjRRlvLyqrFttdffdphy5cOUE5iW6sGVLgKpKhlPJY7NGS
7uw4I+YoZXj8caMbLIAJkX/Dtbt0FjCasZSKDbJKsKO8n5fJwsRDML4w/Q23hbSR
kiOQ8WOIuSwHRI8EIQZHW3+7cXp7KosciFd74u6MjIijHbB5u5Cm8ojDpRnpXrOe
z/6aOSIoHTRL7nGR/YMDvBQziU5pu16JAXcjv3aJjA/WhlCEqsOzIrEjBxvtmgBz
SCf6TKlutpgElZvePO1miAMMOucKmqaMpk51rB3XJHuETNKEoivwrzk8Z3emJhV3
C4eHx41gXZCAf7USF5ikgjT+1pGVrLEHkoGgbLz0w1VAeGQSCJWTsmPmIklO90B6
jc58Qa2R/SaryZhRLWu9/bk9xbPQy+1ZXb7yFMmJ4dgXGchBCSQUnU/VOveW3RN2
a+O+wryUC5XLvJaysGS8r3f6yaIg5eaT7tlQu/dJSQ5XZ3DrXyvkgHirKYdZJO6Z
SkYjozQKpujb+AhBt/3R7d1lHVxndD6xIp26Pxv3SxbZT9aRA6UCINIoK/qq02Zr
+TaKQ7HIx2g32c2P2K60r6PEsotxpsrpNuJxUImxsMcKHEBS10XtAxBNp0gfV2EP
SnH6PTaceqMjq3XgHFqm/kmDDbjH5dQfXc1pf8L8SRagQCUgrSbCeG6hkMfeHMFu
qIOEvgUFFfjANlKGjUQu6wq6ATe8mafNBFL16j05GbX3TUTDeJmDlNpRRD0ZNKtj
rm/5PcA0Y/aTrI7aQ9Sf4v8MrTWsFI6fziWzXWxkfeX/Zrm/TTRAObzXJoyuuVfR
HYZc5UrKoB8/78YqDKwO4h9yYIEnkSD1VrQNthqCqwEzKNn6q1KYCYZXqIYDxg81
fk60e1Iz7/Wc4r0ZcqmGmkAXi1HGUe6iAxTUMUlZwzSQn96jnOYNpGBNkOFoIsnk
4FUJaKzAiAMLvgcPwKHiZon/pKIy+kIvrjRA5qiV/weysgKmWpnut8qWiNwlmYJe
zQlKZRY+31k5JK54+LjCRxlRsEyD/D6DJvSbNETWF9do8mxCuq3L4xweGKGAr3uB
rj87r8W3KQpopBe8Vc4nFSXC115Z2w5Reis+bFdnH8W87FtJ5msUdReV6b+6oqad
zvbINlTf4LgvzDPQE8M2Lw7bbpR45V/cNT31DEm0c1fNoFNyKhjnrqCsP9+7P4OT
Czdt7f8BXiRe/3el2GqbSSNfd8EGeOwfPldpdecMzu8k/Ke5UEVNVOw2ziodkBDf
2hrCo9i8N/aqQ3K3zpEBS8PKJz0qDZpsci9aq+yuJnHziXNZmY08EJv8w997w2Kl
RMVjrWITe99JNh/Y0GPAArWMmmToczPEr2t1IdiXBYsfOmQKZEdFUCqzOe1zuMIp
xuWuTSrlVeZv5QL2IXF+/rtx8ZOjP0bxaHNLkRoCNeR8ZzGiZNrvm36pyJjI1k2y
tymguvLi/FLo5F0uTe7hd9x0ip5872LDxPJuoPMy0AV6QzssbVtmM6bTHexd94X8
GBQUrQBbnO834Vm6F0JwKN8umfgxH/X700lYVTBNi0xPAV+xt0HOGb73a2omrb3/
9AOA0VKL0hkgK9/znckCEbVPADWzqOm8MvQmpvYjPXyr5RRKINNsCz3eoDs9IoYJ
Tbst1uHalXbDc6yBB8mtnR4/kMlmoCz4VJ0xSn339PGTdlBw4jlKZVHNjBn6wNx4
rqOWslY53+WNtX344UZpBZ59Ues3+6CfPm6FlTsEtczuAkRwLRmt0BKN91T2GzWS
xYMlSg1qstnYUKOT1jfdbfkVtAMB/aq9wruXY53bCmg5kLHxWtZfzhorL1FZ4rGx
cnu4kl66fSQjdINQ705Lw0RNHN511UEQND4MauD0Nbarx2JxclEFwdic8I3GDaKC
ApXu+9zvs4ET0eFaZ37o/KRtpNgzNKOrijG7JD7ss1+tcPaVlkAikBG5TiI7zwxR
v+t33BELCoSpq8onDsazMgFA3ntNg+lQ1M6hQnAAO1tKIC0WvJHM7rkHxdj6i8S6
F0Dqva+Orc8grfj61R6MtVy2vpIoibQPfZiQfFXj/U9awyMT0iHgBtFi53T8jK94
7RF791kUAXHxmZo3+dFvClvvaBuUEpxW9Jac1JPkZWKM5BNv8vwr+omLl8r/hMgn
18xLre+ATJSVvLrZnc9S9+UyDjM73j8/NkcuEj6linsTpYvjF2q0+wW2YZUZmeKH
7m7otnOKH1GejNzSYq8sgvdsb5ES6a0uf5o4t86UU9mc8UaFLNnT5Nvm2UcmOMLq
lFaljPJ8EW7qYzNEBA92AWfsH5C13Q2OMrzlO/9HUfEfkIl3bQkBFr9O4sL4ZSNq
mFkpdBzT8JgTyR84W6WqO+IrS36Iv8EaE9tvq4kHwXk02Jd8WTG6Hm0vwQpT6cfo
Lr6PjQM5MT7w/2fzAtjBdZsp+OZJQiSyv7q4gFH1bruF430t5YT+kB3TwxuYIglG
CxbM+9/TJBywNRkIMaqH5Sv7GT3vOuUVP7RSBiE+47I8JUZ+hT4pZMhrmR89oP+m
0g6R6VLlRdr4owK1AaEatBCxcbSM6hSiCiNum7kjv0K6ETRT9IEMHivz/6+pOX3a
88RKDrc/vIhAzXzdNGvQFbRGZKCfRtH8ULo/biBkmTq42/6HiLzvY+U/6VYyqZr8
nTQJjvfuqjDk/DSu2siO5u4yamuPb3fmShrPmAI4XM2VkIWRpkj7dVvTuktN5eOV
nO/YsmJDG+h3VMsM298p1oNS0SkcTtYeJN5s3BUQqhUCD88RKe8tOu5W6BpNGqM4
uM7KrdWhMooyf4skpXWhtxFTYFuBZ29zaX/odTm24KPcde60CTDjm31ipem1eQyT
aX4TsXk53Q3hrc9tMYlJQsjSu4QwZkg0V4DpOia5/fpu09VQ8w/M3uvBrhASssg4
VRYdJoExAgLftKsrd3yZpzh15yde2n/EF5La3tZPWk6BqkT+1HSYOyQGoFJwYkYD
cC8H3eUYC0KROOMVFwfy3BsabdkNWr5UjIL1oTsHzClNMIRQhFmYH4/hY9/JSFxx
G1lcGNFXj5nBsKoJ9J/F3gtDdlIEsTuXW+/BIShws1musxL5O94+Ye5BFpx+srDT
c+mq08iTAklHC01tzTebHVHnSI4E6YP2rB4QxtDZs0xb/DjwK3aNSrASqpdr/N0b
WSayAH9oqfQ7rS0B0YCfwCkaS9c2WZiMYXNJH2Os3Hd5eSjUxagC/c54bK8S7k+B
lCRN7Ojxw6i4o+1kCTVp6kdvT0fDe0FqTjqYm63rxpvhmkihk5tLXKeq/PfObHE6
SIv56BgXpydcR9ELeHoW1j+1ootL2JupysbeHpafnZpQya8X4WGjUEVVnNjN2fsg
aLxLNwsvy5o+nhpgjp0ix+QFoKIup0z24x74ZaZkhimyN7x3C4OtRtNrM54X+n4H
kxlF1yehZKOp72RDFTfzy8MLYxXAR6MEhL5V0N+Sfua+PKVE/bHNfbfWbYCtAdgC
4WSRerSvk/HJfayyLnSU7qAxsCz/qsXvuL7jjDoJa6PcQCYN6umKOgg0zCKZlWaY
LiVdk5Bl2nQt65alHljsXVV9EIJJDBkwqcUJbSIt7i1LK4QuOvNHdmvCQw7rdd3W
0fHef8YfvOWXjGk3V6/C/E8yogwzVRhf2j8VzDWvu5V1wjr9DmYAZxWMzf4c0t1V
qoxHPpWp9TfWD5uT5MdEAtwAqikON6hf0ZwYo2FZUQ8u+WtKAGJmCcUS6E6RLtII
eVJkssjE8ac5Ye4yycHz3dstJJfJjcacs/I2gX2FDALXWMGXz7DF9/oXaRFvU4oT
33FQXxXYdG05HWbLd0oBFbX3GyzX1z4xdeg6OMKAgD5iV8OR2UBV+m6WtawPLxI1
4TgcbuKL0D3H86U/m97Ro5aJl+8LkqG44uGvhLPVMR5fhiobL40woVgcw5Vrei7E
X05eeDBLN/dNqQ59GVEI7mvwC8oQ1TNZAqqVXgiSlymDNNazDpBuq+Cq+qBYqN8G
yioHbAZkF2tj1NeHdnukuVENX8en1Vic6OrnUnQPOGHyJhm1hj57eWANMVa3t8Qz
PN0VSsQzi25xXqyH0nRedEC66ecHUabQqwn1enjreVbpkatufmpCiVq8TsFLoSCL
+F/WJXXXXK1PwrJNgtITLcerDEPWdmWMpTvyYMH9Z9CuhJSbhbjVZFK1MqSdbop9
HQakhJw0YGgfbYmI+f9GX39aeAlNkKrYBYZBdfPJwzgwbYdkELdcNrvccxvK3Hg2
tNWwUvE5fezgk3rnmnjqNKd1mwQfWfBysZyT7FBlebL/vdyC1Wofo41+FPkHoFPK
mYHLS52OWNAcrzHuZidoo0R4aswsGfOhVYEU+rfkg0mEMpHRDCsW2KIxkQ7bcEOw
+eBtlB8cxnkEh9iOQto35bXllszfcHDI6RWuJOYdJKeGQ9c78sQqS4lKGFN47/pW
iPhwAJMQdijbWiQPYkwwRcJDH5ykPExWkOtlmWRm2S4dZJvdwC1m5SSybj2YYJJ9
ONwEScaHnRoL0Eb4taC2Xz4CpZ6NOsXBBYFw45ZzoIv0oPaj31UArJjSmN45ArqO
MdhQTisOP6uAZfl+zV0SGxRJ5SBVcOPaD9CvQqUq6mXnOl2rvTPAwuXxBRuPAUhR
botgLVV3wdtOqlnftRVZU0oSS5RbZZLG1vtDa2+bQLPFxjwbyGZg7txT7eKJcAj3
eFYFyuGDcgZPSNvI5Bx5JoKxSse0xkvgXijaGTpMr3Q8LLDeseljorSRFJNJ7gth
03SrNr1WHMFKaD4AedWLhHBHUOf0RoeutXowcGSZrNWAiUpQel7xkWEUzYjkn8nh
MGBFJricA+RRGwCmDq283x4/cySD7byJTyccWddwfJvJ0eTUHjBCpCpouKaqtibC
tf4ULRscBc1TmX8GkwGnogN4ahjVBCzGWBv1pGizkiDCimIBtUJdjgTe/QzRayqo
4lt2zAyRcwpaiKUXGVQMHRMw7R7MNHHkx+oBhEobzI3BZ74JKh457j1lZ7D41ym0
pAllCy7+zY+kiOY+TtWxpg6X9szJDax9U2iizMBZPoqkA7qbRIdTva3UFcVdjp3v
CMWk+LTGA6fcDCv/fOsM7xGJ7Qo9RPGxV5+bP6DMf2DavNbSTmnUnX68iWsHPvfh
nsjUacuSDC7DVv9vnRqXjDqCKqYwHIumW8yNur4uJToHdZbmxhvo5W8xHktyhM8Z
idyXbTlGoOT/eyREEcDpZkhJFAcQs+kCddVgvT743xCc1/QKqyhWLITp88yFseqX
AlM7Pl/wCeSlv3cB4pSkTOtUTyqgwSInLCH2ziInarfkTzew65+oUihXgnpJW5+D
5CnOTE5QsioQGDWKmE2BHrocnUh3pWviph5JH2eXCOyjzP74AHI8KaZyQmrgm6em
Fs83Cu8PWFOwnNdvCNJ2qfDueJ8oKzXIRSBw5YU+Bp/X/ht5lOwKtIcJeOvi6nLJ
PLjt65jfwDASlaXNONq58BhZ/giP26KgXF5PZHhwigmuBCZ6jJjN15geqVxx1lZ8
tggbl30lbhnqqZh4uk1+aYATXTVv6N/LXbbD0SYlFramoX4R6BnmJMT1H61+t4pC
fbxUAOdT+hFdUwCe1UJHNs7pDQQVkB8XrnjdicNB5pkRjuKHaXC9lHJfkXJOOye7
IJG+4bIdKq3+ANG4oWwmJt5A35Jljsy4nTW98Vc+T1Az5hDwO/HZjfazM4EPQht2
IAGFGzMQQ1BE6NrpUvsyx00d6QdV/yCKPYx1FG1hw+to7Qljia8VFLFNR+7Ik+Ws
Ik25x7O9aYSmdQ9ICxr/uL7JgcrmeQufmi9qPWN/gLieZA3vY2MCmzxgcJZFnVzT
ApUDhgIrx5ACd+N3IHKZ6PGeXwhNlZUvCZ6kXe67z3BUgyEvRf3b9Z69DqvEqmba
tk6MCsAP235iqWNtXFUWuhWE9kdCsouFMr0EMchIG8m5oEEgomGtlixXmYgSN/WB
Cyc8LgH6T68V2u7GhjZ6Caj2IxGpDmM76eHG3PwAsHQD7SfYfPFYs7Xzn0nfUM1c
ScYA54UzOTlMarmxsxXb6xPR4MddJUeUZ6NANi1UOhKooGYrDpuNqb+lH/pF9aqE
T5qEa03BztMBJD/cQZzSMtxMm06IY9RSnnrrpFUH67vu/VsRy+LM7JIA8nDziYMg
WJhzKTR7k4TWtwTyrEzHPSnrPv13V0FUG/+edYwdto0/ROdNioDbjAaEcS2u9/wm
BB19tVh8yEZSOTcq8u+5TJXqgwDpGVPVrLXV0QI6fii8SUi0ZbDkMCuDfJjjeDXS
nZ/tozHDADUQtUx7cLXteQFFgsESUi/Qa36lN5JTx6hawnQpFRvrE5U2x4fj7+db
v8LxTL02x+ZLk3+PlXUAsK+eo0wRYi6lOP0+oKpBjLH5g9goUf916unXDUF3oS9H
ZCKxNrC6XkQTN1lbTy8F28idoCB/Hk2kxmUkDyikAtioHwxrIOBPbhaDZYlLsCZU
zjAm8UTrmemrUAoFdcgWSh8QaYHISo/70F9NCfrgSbogroACGMDg2qSb2gfCH4p9
O/cXaXJd/jt+9E6rbvAPtkfCDigo7bxvOtxkCDA04+nvLAvBKyilfn6ci+0cnULm
PKdytdaeK9lqNa94o2VBiN77g+OKCBweN1jjA/gMtAdzUvrIco2pO92MfYViFQLo
9vyIuJp+TCEgvv/edgkA+2vIyxOPD5Kt36IE/pNfAD00Pq2ScPTsE8pY50UYki8o
n6DUvLe39+JlNxlhUVg+z4o9omGu3olKuLk7hLSzDVLvRYNXekkQmll615CAxVz0
QRczIhL2hnAa7bBwX3sTuUenPYmyPPboyQpzd9pUiEHPEKy5P5nWpCyvZgdL578H
eiVehZfkqz+ac3GWa/lD34va/QIB1XMW0Ejs2r+mH6cqpuEG9qhdmdy9A9RG0H9/
AOWsqem9oabyuQjQjbeIwEfAfUDVwMsK6HTgqU6K8Kmo+zzQdi26iBH87NZTEqIp
/3Dch64BdN5RXp+Q83vzfoKCDWR6DlVmDj057wxQeKegY1wDs+edd4xwyoVOhoRJ
0sz7EuSHq7MfZnHDLHIPlwEiA8A39Ik4NISrg8bPwk2uXL1z7hYclJaRTvF4ZHUq
FjWE+U8ATLLsIFwNlugP7TGd9K41hnyDqKEeVHOtHfcB+Ud3EIWOpL/4caDqay+7
BhJWwLyBOHmPYflKV6B6JIfsfnCzEu775jFApbtHfsLcY+7k+n52AIF2dbJXy00s
PRM73S8byrN1xKzukaDXm+17/o/cIiLMr+2CmNMUl0pe4snjBQWaCyu8YwsTS9Yr
8tgb4D8lWB4vDfOEAXIxO+Q0lhXEefg/KIznLuNR0SsjVko4RP1Lg5txa3a6VeIl
mDjHNC2rJrHhsJBUvo7b5P7gvWublO38ylFuev33o890/M5NevqMGVSoTSqhOUEo
jJhgTk36Tswp8bb0SJkCiRi02XNcg9z0K+Kl86G0d+9/HfBOx2uYrspO2NLYsrg/
HXrXOd3AnjsO91gFG1QrMIEYEJyJwybp2lM+HGZLVP/0fzxCIitTXLQntJGF3kQP
yEXnrg7/RkrhGb0jueqDT8cIU34vSaC4Ji9E+I9tQi9QtNtWSLNcdG7DsWsJCtf2
9JWJ+WRkHPmgVmEZTIN4gwaDP34pKUGy4KAaFgJPvhyqK8cf2b4c/HRhBcZH7bbD
Z27jEkvhkwb3exotFNL6Of/j9uHdtpAGTCENqW8y5KxtKPQrYIgzyWQaXBBSFE/K
opV741dfYLM44/QmPL9fncsWd8emfCN91Aj7H5xPZ2sEEaNdi8Npi8r0RQhhnX13
REPE07N6+qY0PeA7CFliPkZcSuRPjYPM1u9x9r9IuQwdehl3M2VW11j+FD01ud+q
XJLya+8UR4/Rk3b3aiviGeRzys73p65qN0eArSNGrXtUFP8lQnURrib1UwjNOYeO
LWSJVRCUDwIGXG5ZTgDTejBSWcTNIqVBIr/ic/Lq9Z8cNZhDHfpBVM1RbKPxi0nv
elTXVQTyE4GO1+jKAeR1cvrAP1S4lkMQ9p6ciPRSrVp64QHju63nij9d6DEhTY/F
KeLKVh9Y00yGIK2x7BhMPt78TmGWT5hH8vlbNoHBRJ3LNq2SiqoN/Qr9bnYYHetz
N5a0V4ITleJWJUd2NEYV6ify3tdVYSTG44txQ3iarvplw5MBDIXyOwXr8vh5BftP
YEh6lp462iEfCDuLGyEfq4WilVEP1hsIn1chz1ka+slONQrSYF707y6lmcZUcvj9
gLn6RpxkoWvbC82+WB3sKxq0BsUaCAIchMkO1n7eebEIoHWLH6Udvrql5EjhfTui
JOlgR89vAuGq4ms3CmdOyEoQjktc4Ri/x10fQnzW/OfClLQxb4riiWd4NTBKezjW
gv30PCSYnHAuGj3eP0lQmNeRYlZWkiwjZ0Cg2qAg7XgwjEMkc5IjQYQyBa6GcHA9
sK9MwRaSvrMeD+HrLfCXL15filUcck+M716zUeVBefmCg3KoUIqpX6ga/RHp8srr
eW4jaW2EigFAR3q+blo9nztxpgr4eP70FkIf2m7eoBYlQnaPIRlXcevRkQta4NEE
UfYUdXWVgRQhdkf63w0gU+fHMRBDTuJmOQFWmJ4okxMbHkDEHzPI+eQKT9pNHmXM
zq2Bdn9Jkt/9RBWCNn35wAbS3Bwk2TBiEEPqXgafKuluvOKRbxhSNz/CymXVCH41
Xl/NIIEj+VlR94e16mUA/LTp1AWTjobHWtzU23uvYX+bH4vM3+5Kos6xb9UJ6jKX
GvJ8GC1I7/PGA7uB515OGtjeq0EN+3mEDAO+cIUsUF2UtC+vafEFfzvq1/aqQpQm
Wf6Hc12TpLJD98gKIqFCZzzcGcAVyHdIE+e106q3musL/si/+sdC9fuEJiQ+8slB
lF7MlFxIODPnzNm+hqBnIs6p+PwNmFNiO0ycmrSgjCWOxprHeJt1pdwLHgs2Gnms
9uLm7oSptgd03GLiqBn1RwDnq+PTu8xkteqBjLybvpOu5rs1dZU8zaylgcKzNuvT
W4UFUO4xsxmidIGJJqJOEb1DXaAS2cTBmhxGE1QDt9zFrEB0x5wy94jSOexwG3V4
Od5BRvNe5H4uvx/GURItsCRa98a2cqh2YYNwcoAoeAVgNPWnMu5ymHC9uyO+9vQ5
cfG129C8XOaJ9s0j2+bkUYv4AY3MAAHqxDo8sBCjxpE1Yzm8sywMYe3ZOV+VqITL
HJiBR+gJFEXTRFmY+LDC9CBhWxMk/db3ruROWmFAvinaVadak3VuOrfFGv5enj6L
nXDKyl6JxAuIPPIwJtENlOGI50ACwWGwp9MYi0MSEUvzPPdnNVPq/acoBpIASyF9
BgWu7X0lrLxFU83hT/67noFJvcgQ8PXHV1UKQNBhiGYO54b87NDJpU6Db7oTnj3j
WKG+iUOO8UqktrMiehGapDs7SSY8Gab+DbiXg2bFh21W2sGCyLZQsByYV5hKmTBh
d6dQPOrdwQjff2lKdsI+OgSlc5lscrJMgnHN/91m8msJkaWuvIYRdHyFblguSwrY
QD91nzwKUd4ieFLzZLxNvGTxYC604NGX98ZfsdneIU/bcNpt1z8uDtjfBPYYXd5A
WgW3TFgSdP0lNhhLCtB52Gi1Nlq05zzdobZwuU8QuJyPZljCl4PUdxzK0yVNrSKd
tPlw+kEHKnf1YIhjIyawVPPj1+f6RSS8Nn20AuZEILpAE85h9ld+1a68hWM9jUsW
Oa+b6oVslTEfOJfS4R2NGoJBqXyIyRbFEQERzU1xmEfSdwKBgH1J0OXRwlpaS78Q
Tt6XUAS6C+j1O2sxfGvMmzxQItY/4PWmwcS4flPkW7Gy7KodCKL1ryH4deyKZ+Za
N+RilSw4YForIIy1fXAqe8LYl80se4l+qA6eMKsvY7sTffEp7M6Hp467dB0bBtX6
5XBBGFptxH0llRL5yu4zxrzz7FfbjdH1WCxEKNv5Ed59t9/tvLl3OhP6DkCMjENG
msl+V7Qb7HSV6unpzqSeNyyE1LBsrPX7MoAxdJJDT18f2giC/NmRSm6v4ajILfxi
83bgQF9UTxWmA6JtBxCEb39o7ZXy0UYO5ZzEnl+dHHgD9GRGW+s7B/gec59IMjAD
4gHdQ5pCHBS6trIPKu+XU7kXciDru0udW6ldQ/m2kAfX72fa4TICAS0bG4uTGjZU
U0XWQJmjJneCK5SPedCE/u/NLiaCQ59kp/4vptno/D43884BnO06udjwbKT/yWAF
7OzN5sS76UB14crv0mI/CVvJT58HyZNLNxuqa7b/yNMDJ5335PQXRVo/fdIF8FwH
ayaa20NN3XXSQUHO797ySbJY5+03DUV7DfqERba7n+KXWV4+dQu+dxRLhYFN7a6G
RFn+Egqvij9dRfqxqK7DI+Y7/xDJms3tEbnQetbxLH9++fXZWxeRxrRy2F/8/Wnf
p2utd8Cq04H9djZV5k9CDKj4TGLLWVVD1x6gFV5vZs4jXR23MLxyZRzCIT+6xJgY
pBFWIV843anDspcZK3B6tINT9oalHzPuJzTLfC+PIEf2Um52sage4Kt5yoqn7A5h
jHAqrT377EyCjpbrO6V+HJgdDn+oV4Hzxm30KKCb51t3oqIn40LxDkejPSPsD34O
VhGli/g58NV6hT24vNL4SGqvyDOqPQ129MGlYMeGMWa91EsDvTNsjepF7Dsyws9u
RH8IRxZJMebY/3DEqXKMgbKEtvY8pVrbdXULUPKqxhVE1vtlNWs0yPwy3EicQdN7
1chNexA79zW4K/LeG3QzzhmZDtHzxx6drXuQtolr6HQKzNqsMaU7JG1BMoJe2n8H
Q+HFnq77dw2JYGPP4S1AbLz48KJZFHOq9mgTPonsvxxjA4dz1PiAxsWf+YDhdr2P
PnIPs6DzL250z8z38Olv5KXzKhHerjoiiMyuSLbj4dpTKIiEvlmx+E3xKHbUAfF7
uAdijrotN4bh30q41oXbezM0tOi4z4BdtKL2EUrkxnluylczELpG+/6ItS0BcHis
V1/KS8cj1M6lt+KjyvT2fgqYetRSqKgERJXN6mJZIRNNBmu80dsjfXRi+CB8Mdgc
Ek6hJ2/2IHSyH+0JC/4yHE9e4no1g15j1eYNtfI2zPFUOjGaZS9nF5SHa5CbB3Ra
MZYbucrNmnK6QD9ss7g7OovkCogs+W31C0vKRcLjUTrqAdbku/IUsIUTSV00vCNh
nDLVTAy0g8qug6SrTEnOj9Cg82jAu9bZdppsC715XQ5+4pxyWS49LH8DRBEgZ6fe
NeYCWNHfidEe/mLkc7pQkY2L0zBMZtu7rIimOE8DWTZbIsrc33kR8lGTdyssW48b
EB2Ub5ghqXN2Tg7moQtW8DFr+vqSdlnh+v3dFT84jIvFWsob3Sz0EMU6nIvZCxCu
AGftpRJhLy6nnqvj2mE07/IdxadT6nOR6k3UreUIpjV+xJ/VYMV6UjBcAuWMuZIP
ybR33TOtIdnu23LzQz33nCeo2AYgoQyGTZzP0yLmzYXyIGI52g4NzLtFV9ck1MxY
4E7/XyDOYPpCbKflibt1IG2jDUPuBnKYtqG/oVsjXZXp2OT22uG5QRsKWYQiAIxz
qcbZM6KoowUtSKLLtcM6EM2+lAMCCur6AJHPkf3rytSLvHQ3rzsaH4MxJOkp0Rdp
YIj2+Z+gyS+RvpsPoD71/H2Zzcgc2E6EGz1i6vF5LOAqgzvLSpR7mmNUTbEMp4Ov
5oOMGC6bOEgOeTxTzKwbF6wbYxz/E+bAEyoW5AN4U2dFqM8ar4AvxEgwB3AnA75R
gFGqL7xLnunGnxngj3j8jWcDepWe+wKwIc3le7H5iiXRIXRGWSfHSaCdnORsZg/X
+hIPd26HLE48ZvIdeAUidSLZs1iNKoVAVAxI8VlHtqVjxjrB1VfXbdPtIlInPM6i
oLJhpF1GYjczeQxZ5iJoBZ2LdMnaw26c/LEP93f7VE+dSQD+7nZtlESYNnmdAZ4U
RqyrCK2bVWkwtDLbqLCUrLfaDemTnHbxdQda/VumsEfkB4kZEgp9M0NoOiqR/2Qq
xnblbbbQck/fi/0zZZGerRT6geyU4Me/fSewxH/fOuK3/1RBb7bReD9GCPPU+Wu1
X+nzOrpQDDZdfIwBT423yOw+CV+fZy70/zaTIU419MaQtTGwQF5oQ3JbfCuuc/F8
NEveKxcYObJeA6e6JZDcCuacAMGQHrM9uDzVtG+TDzEzCn0FWZ/ZX9gSXjtcEW02
18WXpgsV0Udj9BBt72eWmIJYPwZ/OOZ9erC8XAvX3hlRZ/RD9dfvlD3S1XyJk2Zc
GEFRQy3iYTNmXJpitHlI1hYAHHiwOTSWIouo8M5X1mMRuokTg38JYvtEuB5kf676
76zf8VXHKnqMuBVLq9Dh++fGSY10ejR7DsVcTFxk43udRRMlE4gZGypD49upAHIJ
Uj1iUFXMjNX3al4Vf+P9OTi6AIZ6WZrCjzFYmejFSceOWHhCvfUUmwswTogonY2u
1ev1c0aP/cQgZkc3c/IGpTLZui7qqQ8/y1voktJtdexZrKzTatrYLxBh+C08PRcE
URMzclmDNy2IPo9ra4x4lWlbnvI3NkPVD/fVS6RMQ6RFlaqF72YgE4e+xb4S2u3s
zG8eU6IM3EQCeO0mAS/OnzECTRO03I016Ni75Ax79DOLwqqFZV77tr5qtlBH4bo7
5MDWdkUGmwjOZRbE9+VqIHpLRdRnzoVe5mPulSOqrHiuFn2yl3VIhlbZISLL5e+m
zhD313J5XWJMpR1DaZF20LSmyqFHyXYXs86LiIB6pYeg2HOJtfEgedkey9o+IAgQ
4cNHvfKEUn4dbaeoCgX2XlTNuBXjT84chO4AHzw3/g0qcnTpI+IaFL32IaRZuFpQ
qU6cHSnYIKi13p81fH1mbNGywuRGmqU5nzT7sG5cpR4Ibq2xVFijKRGcRyN1Vv26
lH05AdWUgQLcSe0SOWJGqmwd1wqLQs4zONmBXfyudT9Ss2ifaxxx9zmHNOXdZxWt
U9t5UOJTPQmY71yQbSePJ2DOwWyZxpNbMyzdFX4Y8cyLyGG1Wea8+c9+7jmIwEUQ
6OmgqFMykUnEkUyuwQjCnjF2CstwFb4QZNYoLMo78jq/CLdcK90wp0KOtiq1NEl7
ezlErsnF185KgP6UTnm2gux6rGifPLrZIKPo7yyiye+rCz7ovSylPuR3LIr9/91v
IL2T+ps5FmEIRQy4Mk517jyQ5u0Hwy+BuWPgGbx0tEgnxWd044ALYktGls3pwPKo
1S7AhAuH5fZe4tiISU4EijE9St9GxMNIRJDFQtNlv1MDlF1/pcv3csM5FVOl/Xwt
r6nrxzoNS/65SZBZFjUNtUMcn1I1Uku/jKPl7OSbg59ixqFMdK9mmvBpmbCWSJ8y
m8g3lcSJIR2zTXfyxb36xuBZm3z1kPPoX2VHG/mDFXMT8YuxAq+PxV9nwzBWVr2r
Z7y9T+ajcS8NDQisLnZ0MArtTdV6Yu0/coJ01zYNBcGYy/srxaf5gaBjjSRJ582k
yY4BX46Nnm//MsCGt/e14hmLInSNZgHBQaiuFRCKV1LETt62VRstgW4YkctVg1B2
kSZ7TPl43Xh/1qFs+rc2/ZjIaBZXqIkFtVDaK/j4MZ3IyKIm5+4Ub6fb3KrzoEBM
xp8GQn25WpMdMdU7ef0GKIkY9106mKPL0+oad5l6Wo4RYxRvfNleO+l9t/rvBrji
/Tye7YJpG9Fzqn/H3lbvAp8JDjUaQvW+pVgxv0fl1doRpMUB8fCgN9jkkokLoD+i
KcTMzyJlhtkm2o5Y0LyIqlk35hTKs4suQdZ7dm4QTCXgkSDuJdUajAg/4AgAPOs4
Hzt2zl97fAfVC84DJQmd+1LEsctFwI44V01P35/Z5bToYQBdaeAD6z6uYubtEdrc
iodDU9i4q4sd54NjkJj7ZMip/hfydJRhUt1GGYtX1BDi+o3KNBqN79ZN21dGViGW
eq+tvTOPlbFLNmhxaVTz89DasUtJbCJP9WrvLCP71gLW6VHOpEWymm11/jApPhTG
ViB/BaY/iJhyGufNr6pOvpiU48W7jSvjVdg7H+ezbnf/jQUrStOxbpM6p+EingUj
wZ8mWzn96eef4TLua7fcWDvJlfEDyu1svwFdC1nzzBgev/0J3ejd5WXlXQerMcOr
H7zeNfefu7Qir23am2H/KIMKJ1yMvvDsYL+q3Hv9wQH+YJoZwc52olyPmIuh7VuC
6xDu2dtCQmxFb6nYE25HK9MQQR/Ysn2K6Y0I7C8NE2dFk0agnLL1GPDQSJ9aIsbV
HDc5R1GslV2OFNRkjm3BTtZFN5odUZZhuQ8aEX1ke0rgrT4sZmnv7E2/xceIUspn
847kDW0sQo6GKobU+CYw+R7EAAbbeTXfECXVADYemH5ZSoHYRGJGeF28AHce50qJ
D4FoMdKfOR+xpG3aDCXhZt9OVfJXeQZM6Opzcssk1jR2fNqoLGguSDrxRGdqFAgK
zSG6B+lYhNBeDKc/u6TVU1DEXVfI28vYVx8GWFDTLj/8FIWZA9TZFtDezDc9plBP
KdxNkqty00KnHMOZujIR4fJ4b++jKnoYxuVkWCSu/xlqj2QKFudhiKmm7BYVuwjc
pLquKlASXxzaQnEFKUe0yLJ/cQx3XxT20xnE5idxt7FZOTmoMCgen0zePKBd+Lsk
yw9lcNzaGYsdr5BFtc9HXL4ffQNSZYHoufM84Yd39pLimf6AJfDWKfkXFWvi0PKc
BmTV0qcaPmjtB0JaLutAnkqs0Ph1AbDI4pDMvFPRhysPwo+zSNyku6IoRxqXYjEW
WqsZrPzdmMLCMY/nyYMhxzmGj38uFgWtwZRbqsHdeLdtY1K0gZeYKVddkegvoq8I
HxlQM83xGnws7dXPsD/Byb1xtlyDDV3XGUOOm/GPnD5URB0vaMKuZNWWkLYT4Htc
SGwBZvp7jH0xVIV5Cx+cDUcFS8jwK9LjP6RRBN9UDUhfZrDP62nx6GH6CmsPCZ7N
yCuzRHu4X6sdB2uFSLz3/qu5gSl/XnXNsdSiaMEwXMW1SUQuO3U0PGjZ/LzwrcKJ
S+hXmBnA3sB5f3hzh/aIPhwkWxhSSxpgcKx+9q/6JiDpsoWgORNEqNd7A641l85o
A9HeuK5El82OyLBpHE3Jm56yVPpt3v7Yh2iM0eoKJs3dRWvuRp20SWPVGkbk8HC3
oBxVJL/hK/Wsqsi8sNDRftx25VnPA+LgaMqY8VEY+OACfHn8IwLyjfTz/8HdMaAU
TRivaw2y/ntBXdxVw5wY98cO0v1besQFvK1K0E8BSzJBmuPDW5ShM6PhaEK89LHC
lfuAwuCbh2cauKfRDgE/pkWwQcBEIj3Lk8zg+uVbZ8Jl7/9bSvDTD7oYR1WBtXO7
RDmGYLNgOxslDFwn5rRO1ezahfuLm3+t3vSDrRGm75Z+ZMM9NztE3BPvOfmQS8Eo
JyH7Juz+8d+esuuzjRXVrCrMP4WHLRhzVq2EEw3OyVEVunbWVmlmNk5rhU455RpJ
ufFN8akJbh2ouowcNf3VWKzXYdUf5LGe9+03HE3lTKRosCjJ16AUUaJd/NseAcvc
RHKvzdyyhUy+i4Y1Pz6D6xeSaQOcg9jTB38dJkPw6yO18LhmT5kyPV6danA5olgf
5rY/D3vDV86NOMBqtKKC5YpahrXLWNGD6uqnHoYFvNlvU+WcIN+wp0z2AbEsR4re
3/NzDTGkT50zLV36U4mHRkX9ghDRYepfaG3y3xyYRTbFtTjB4Gk8HAHiPv3Ph06T
L6h0yZVE1B3dmO1VLLCMAlD3aFWS6hVjaOLtbJ2lhfnu9DX0HmiNOQXPrW+aAEoU
VmUmZZyrqIjEbO8Up5cbb2P2+UjxK/bgHbIpYpQzYWfAhNvdOh761sRgrGxm/I6U
i+sT8I9I+iOYKv3xhz4K0oAZiNdnyAYQzI1+Z56L+Gb8kB3Z0ygtfB5AMdXbznLt
laM2phl6pxdyT8xBYjAFNUBKQAuO4rramS5BlJbRwLklq3bVg5WBLW5jjZH4ZETG
FDzNhfnQIL9ouMbwtysFupIkqH9FP+JGGryFHbBlerUBOcTMwJDWk0zVezZxRFNa
tycKPrQSNZiEz1LuOqhkZ3Ci4zeiBl6tIrFZSfzT2ZSMdjcd5H44VSVWYmQOF2oQ
11hqhj+5VEBMjJrmAyDPkC56gMyzUnyYDa7ShqPnBldWuDQry700HKopEhRE/3jC
D7gwl45sL2h7YqT4qKEEWy5QVNxJn0Ghx5So1rWffxWFS7iaJjAHpho7bcqoSbz5
uvpshkYIx3vC0MuYPufDVV0H0IeAM8JRtyWKv6OdYKTAZ9nu0AXb1aCgEotHUw8Y
ItcrIjZ1EHjIY+Ijbad+VR5pxkE3/E9bTWDKbkCo7XEpraR0s8rcRBEPDeMvv2cI
+RwznAjR7c3niAZ6K7f+U6y0OmarKVu8pNfQNlVnRSREqMxn9VdSgKbtCza0lYuA
4cgtUzR0kPF2ScvATV9rAJrT50XHkLJ3DA+l2yu3LiFtTVhItGEAT1X3v7/IG93Z
WnI2431dlRlOSr5BTusk70ZC7pjLqiMQMsN6sJyv8Xe2E3+o3afUh66wKtJsUuby
q0S9Ng20qmmd50cfxWr/5pSfKF7a1H8nhqGgJH/UvDtT6cNyLPzub3/W8G0w133r
veSOoAURlLnW2433U2tf8MpBkf//7CHpPS4iEW3cM4Y/XCwjTbTWEHY+PhJsOnUc
NBXQB1l43GQLtZtwfkbng9R+kdCWKU4pVqXHnGU0nZpODmfDkBdVigGxMQR4Dw2I
9KxB6D+JMDAm+ra9zkaPfPjq7eY/hCj6BWBRnwEGBkToPl350K7YkST450OUIkfA
pPtm2/EBIJs5JlnuRC1IMicYPWIXKwcltdXali6SBONwFIgYzKBFLZjMMq1Y0HNt
yi3tl1LK9rUCfK/VugsKlL50Ud5cInAwS0z4ELxuTClmqSO0zTErSkBXdHOeYjTI
GQtHmpkvFYjybbmafmLYj1QrU1tUFJfnGQccSpdrMS5pUoMqor3ZALMHmXC3S1dF
rfvoyv7jnMlrPzK6hzsV2rorFnbIZklyKsrsQ9OIbt/XG5Q29oCh1l0MBAtJo4rR
frESGJDRuOtqVGu5CD4koue/jLamBRvqryYxFbvP4rNUF2t85fzKfzG2c2nIzYBB
IFYJQVEUNUg6XZEVJCeVd1PeJJAdtCN70lg3wCwAOM9e3f+DC0vEgnkBTPaAaV37
0C3dvpK1NA9bwGiMfLBZdhqxea0BczOZXlNXN/b1ZJFcWslvLxKTzzOZhjEFr2v1
/0Z8Z+OiJDcX4tBr8150GpcALPTNcSz3o+Fp/5QfYVtV4Xoh5KR1HgTf+lfeNL4M
yVtp+sAONYUU0VSHlsBBzfkdk9tmOKisFBENxxHG2B3dxZm05uVAjBNXbQT1Ury4
3YYkaJYB5NXW75QG3pc7HGWn3RpFC59+QE4c5ouUrg2gbvY144+SjgVWwEx7DbEr
TRziNtr1g4Zo0qIurcScLakGv9peVyG3Ozph+PkdoxzQURADGRNVWD0NUVM+cT9n
gqw48Yd2nWsk/ZXtPUOlO9oT3MTi6c3j/1ayeW2rrXdPZrAjBSS9BB2D7U3k0ofO
GgdjJlIt9etZy7w3tA2ZaL6Vkl0G27DKqJ5N+2h8s7AImFh418WOj0SVxqXPH6Zr
95uVSaX/ghXjdTh484JuxXX1KsHI36tMICdxNCxB5hhgWMIz1OJpKSnYNVbc4cG/
pdEtvNEscQGOSvKpvQyX36yWBxgyMpGB25r7Vl8iWpEadEFOIanGeuj1ecerdIwj
rOp6zZMpOXKUPVY/OQVpgoO3rpT9hxadogvejxEQSHioaz4Zp0yX64EqZXHoZ9td
b9WvBM8mD8I3+29s4k8KW1jt+u5KAUl9b6G6r+zv2tqtqp35WPO1PDzojAXlcuCf
T6JXmZIz/DNmzh60QNOvgMgk8V6NFchQ8p4QQl82hupH7/KQra8tzsbHTtUlR+4D
/wJp5ljVtW41nITNUqqP7FEcFpB28vkagzIyedZwU4G0s/xNGKIiX5Cc/zt6F267
5nYrKFvb329A8ObhMWvedCNkWzlu9uy3yrYTT47BY206037O+/3eAlLEHFoP9WHQ
WO1vt3b2XpT7o9XvZL1Pwep59XIR3WHS6QgQEpTK7hrO4FJSRo1aIbsNGdUsSJLq
BjAtQBR/gPeH8JIwbToQCGujSWQIpbmSHB1XEu5xZc55Rg/2Qq87HiHJTfHe0CWR
unMll5nrX9JqwLy0FWwLYUNr7qFqQ64JHTmyy0bJiNiLC82q7TAr2HEQgPahgRzs
SSg9IvztJ9oHu6O2pjQeKSyKy6CDhtVwyz6c48PqWUSdID42gVebHqzauwrYVxIj
MExTM94g1u5do2cXBr4O9o826VD2oJB/Hi/6g5hdsvT0g1hEcBS3h64dxLyhiVN7
SA7cWVBfO8g+E0WR8n/LA72PelP+e2NMkFnZArb5JXcm/ihzklpEjInpSOPJSEO4
v4yyV6TsXTw2+mw/c+Sfb04Kq2ZFal+Mryd32ZNidKgJYD+AH4EIwsP+inR8E0Y2
9y9BZiyy2huMUVLddRIOJyoJ3fbYnDtZm32+Z0yITmLFithvEKcgCSDj0L/QywTO
8jWGBSYqxa8RGztmJAuAP4EtA7LBZ5k1t695f9Esde8b0v3+UFUqCK0YM/GBxiNY
430nVec6uXe4v+sCjeDxMCJ+zlf1+zmDGHrwOMpBNBCNBYdZGZMxNACRQbEgYEaF
spIdJxk1tPDmOAahgHmL4spozv8NSgXdcG0ryictc30xb7+ASl8KdggMAxJMyctd
Tnx+tDU7ppIafEFWB53HAj7dPcUB3XCwe9Ma8eXwvhGIKZoueTM5sfWHAYdZv91Y
X/BwyKK2NBMRlHb6ljTZehA8HTnaTHzxkqphwXWKfQAmJ9PMbZoNjCHG4JsMKD2B
xYl4LWfLzPPOzFH15sva88mywsGqPjJ0fwkGTwlHKfG07v0sCDBSZxKhbIuiJYXp
it1NqND87lWwCwGMT/6h7QXZSCvfJmTvseNy9If8AWfUPYSSw4iT9JXMDLSQcRWm
MT5YTnVRKGCV8IPBQuh4TuJILPGrTpO9pJgkWFO+zGjlgsSWcBZxYMw7UISPhFku
+dE4GUfrNd0x2MpC7EdclEpgTU4B7dv8Bri9lIGUcyZQEOGtFTTMKqLI2elO38UO
vkWRQXp2clIFGVEI/bjU3cP6XysDLkT90k9li5EewmMukN20BZRluaMxIBWWUYgB
taksvhGWcHrsfxCjIHz/nkq2S/JfhN/FOUJk4Ev7JO/TlS9tvYn7HSYWJNp/fv+q
QNMnaT8TZqDGXoWM+B0FsXR46BLK/19dusQ6gK/AAyEpBeg5stwJlO6fPKIlsCeZ
YEfRau2O51zlkQHlTMJMcKQJ184GWzMY/6dI9UbtFhBwe8gUERj+EjFadCK3mFR+
jo2B9Vvnl3qzniHXe/T9NIbYFjuK3otoTXINLghlEKNo8rlHVSzUyWtdMBVwUUN9
N2M4a9DKWdcmExVaSqdwkSnmEDQCoRkLaXWFNhDo1cZ4a30kS9S8EBM3IFEWrLvp
haKxexzDXcwG/HgwjU4QzedgQVXOc6UyzIfqLBPDwD4+PdR5rAbFD2F3aNxyIXDG
1E7e53UXQQjoRuJE2cKJHkvn4aGBB+iGARG73W56NViy+9jxCIy/1uOh3SPVB3ge
L/ERAomLwAY3LVlLyGZzdIwT3PjEWksjGJ27zdqvNG+YkcrznaeLc7430VZflV8m
R7ahwmFn7IRYLiEPeuGcwGBld9nnZQu1WhkGu3gDYjIWcPokCC7YA+zaqTcbzLDt
E0UwoK0QJkznl0f9fuVq2ANxnJz9c8J6DJ5SFvBjyaLD0tSYVMOs0EdDffEWJW7V
0vyjteykKGFh6SSO8/vVuKC+i2zeYHNG9KVYE1so9EbZKZeFTczd/6R3NBdhPWeS
JrFllnGLYAO9q57mgCJvXeSUjxL2RDp8y0UD7gBToPHX9fZGXsnuuZU1G84DtiJt
iTHqA4Zh0FNsLDrqbL6Kc0Imr6nMNyzMgLyKvXwvSnCACsCjNSyo3/aJuLFqMdTA
eVVMb9UKkHxry3Qguxy07lJPG1euf8cg8mcgrkFQzdWXmhjsXWrhOW8eSYN+1EMu
NUVNQzdF43Dz9piSHgXV+wU3R7CCMp0tV6eiX9Y8OrnL7qYkO8C3aD8ixbgrZ/ol
WL5Ojp5Z+Pz4eNHDaKDpS0wNSM3YVM/G06Z1VXrULSQ0u5MR+Ogh58VNGbOScy9Q
iMx2yimuMey3ILxIRMJ0dkQQgJeY4LKDEEqWoW8AnhSMt9yPlRA5m2VxIAn4LVQz
qxOJXtIp2O8Pbyz1wWoL8IDWyR8PiwQ69EXW3yjRQYhNLMAuSJmlP01+IXl9h7gk
5o6vqUF4xktv5RB3V05ChvmKp73FvKTw9VqJ0xA6QazpIzcxyr3DxXpsqv8MZr0F
FvVHqO7KktvssBlGd7SQnXvIYW4uM64bopFCVli6yX7/T7i7Y8cp5VqCYUEudwNw
MpFcSP9fBNjwEVKhtlP+GhMHueWq5FgpwzU0z3+9iOQIbEr0hAXcQhnD6jFlblw6
5LH8sNWgzt61RiEcqNKzveHXYmJxLd44OaVlL+Mwd4Q8nwdonY0xmsVGzTjxOw9V
7sXdBN7A2tICQA49N5QfEeNghWVzX6gqtD+gRJO2S5hi8IMF+wtoSqfMO8GF2otT
TpJ3ayOX6hHKr3QGIiR8McL3ZtdYq1WgCFzgo8avs4XX5SK7hVMhD6D0zYV/D/ah
SD2l0Of1phb/IwyMWE98izlGsk++oEREROMX6XK4LjGrEnnpS0IHaeMGKDXBOZdR
OwqwQlwZYfcmn/97/u2j13Snix8cDvI4A83zGH39RAjowdITDzAJ6W97KwAg7+5o
ZwcTEuBglf3n+gSD318G5M5C65/2vdujzv5szjvV6VU/Pd0/Tj2qq9s2kvaYtH1v
iBZudPLuqAx8ehuoyNysqbihH1NlmIrqYFJvQxLuuf4BBFx+L6JGllamMbiZ9FpB
WKHcokzSYTWKeyiokm+rLpxaYhtY60CL1whp5bTrszo9J8E4Kw2jjfcafQjTExxV
spnLP42WSP26b87gdKsuyDwke2lejOm2RBt946TW+b502S8pxXMMraGz6gsHkLv2
63XyRnLeeUF262WCnliYwrKO2FHtluXmrwye2dUKQhssw2ZQqpIee7uzZiiCD4Wh
hL/zc9WI1rVhlMCuiAfN8l7ymSJ0NIVBqt7krCiC40+LqYdpoUEp7HGXNovDMQrO
533UxB6BUwDrn9Y/10tpApHr6vqRBeluqual4UhlxuRGXFyBJ4ontK+4JYHi/cdJ
QRzN5RkJAo43L7dJrVV8F4/+OQN3j9vGLAsUorx3C2dZ9dpF5FD5Iqj3tIBiifKQ
eIrw0XZbG7y2BjJXA2zxcjIMifwnJWVbJ9H20hw/tyDV/2IL9VJQg2b7kOcZB+8U
oM9y24E868UJbbDlK5KYZQF0Wcpw3H1306iA1pDZd6c3DiV0fnqwMM1vghSzSOlm
s1PNT44GMCB+zLSB3wowJXivPDw4ruCgiBYXnKHN0YN7W3+zzeeEMiuqoKtpACxW
YjNArTXhE96HQVLEjcCvtau9VMnSIMy+DfWMXm9OBcBOKwMchg11xinYZlzjLN2H
sIE0WXDxDZfWNFuFoF0yBLN48sjva6PuXiuE/TCGXRo/Y7NW2/gfGI3NB6Q33S28
7PxAmS1Ox9Qy4TKzLIf0o3NbJkau99CZvTueTHi1jyzlmcS7JJbJWlsEVlpoz5Eq
l1TsPamty3Ldtzcv3ZvLW3/lo2oJ+YK32hHxt40TNm5bsGxbGEju/MSTFGpCHYx9
ta55UYpxtGKwBg/lFQazD8R8RARNR1XvY76+66yLryvyTCr/Y9J9/kbuYJmkzeHW
IVXfQJ5t5saGIdCLQ0PMR9a8NItWVPcWB5PP5hlB9faXnqbfy6TzLRBRRRWo8fXO
g330AKamPkdk24ETj83l2B/hgEQFLVkra8chmLgpZmfw2vk+utpLji/V7u/yO+qt
Hk+SHMqGkrvYnQOIvRoAcX0LHv3MxFa6Kmsufmj9BKaIsWtHpxaGF4HEhf5OwTJx
PHD8Y806DLwZXdl7kWFfQ7l9YeYe+mi7AC/a0/PK88MOors4TDeNn/uKo6xWtQNs
LZjWHVDSADMhU4nziPdLbKHGn/fQvZJi8DSaBHbEDCx5Z+iYzW/CM0fMTPJxNcUl
W8NkZYd1SSjGjIIdnZSqMTYPo/ibbuuhCSBdhuzv6HilT1HDSsr5huMaVmG3zu9p
E1Gk55roAu/jQMtbO59ndMmK3gHJEmI/iDWy+m/IJca9MmHo7d6+HrzBsgr/X6fc
ysb0U+Kx0s427LOVXhZif/uwkrw9Nv8zAq5/jp03ce3FxxuP/1DPEyrdWYi4pEzq
tjemfZKjeVAsjrXGZCbODWJtcxlRhBwkFH53kZfI1yXEJOds4rBiGYHjzoQb733r
WzkQOfaKJn6VD2UOE2dFG5wKLf+T+fnPko6U9nhd+R/vn+G/asuemQiDqNyGEeTw
J96+MQeqBQcYEFxvc0x0WAvkjH6D36Hcomojn6aYk1/8g8QtiKXUgOagsz8s0bCL
BnEO9PlGW096EqgYjn3NiogcjgEZRr7+1x7Vpn/zvkDYj6CnySu4wwLbSXUQqVj0
gPpbvJcy6SXFCspAvyAEQIM9QpgCXIJ+7uCtIgzbexpBnV9OSc1p0TLw67O6onu4
xC5Fji8wIUvuqzHCHB8g5xehgxOXTqrrSyH4KP3qWUvD/x+zp1NM7Cjik4+Mq268
v2E1rR9wlMBykHxnnN+OUDnVT6rR1rkGkDyEQq4BqyAaTczRTxnNUKPxtVawhZr2
rV5fnTcx14FUmNrE2zXJRdPUgfVqoNP1iNDDTcwxOhG/8ByClA7y50CoMmQLx4v+
4ePA17KHoH6+sVrufp8AxJoYoYso97uClu5Uo4jbTvxbtZ01ySAimH2VTnJcEpTE
tZEcnQPEV/pdIL92Tua4aMTlXXfMlFDofRjexQm7ec7NkwOMeiLgSYb2oDDq1fgo
X3+pN1Yip0zoNsBKI6J6dqNSpwB78WUIUZBRKONdPVm0tNdOMpBvKk3sVgTB/K8G
JEwo1je/mr8trm5hMOHwaYMLXEDxAyWHOMTmVmkt8Fj2TSO1/k4cm8HbgimWZZnX
39lhb429nZI+bTQuoQnAUdayX2sUe1c6+hDhkfyY90egn9WtSD9C/MmtYK/MgP9o
tSPnUbhVRS0XcOObAFaZPslKHundHqG3m0QxntB3BalDnMnRWetpgIR4gMeYxKuh
npaqH9smxODAgGT55Eoyzry9G4d8MSO+X6NR1P5dm0CJ8qKCZosUa/dOWnY0N9z4
tZopUVPEvEYMVH2zelbikEgvNeXtUyf7aQjjKf8V/j3D65qSRRkjMUzltVluSaMR
OxoWVMjSzqHA7AOcCje+PMWQdv+ifRm3VklC8tg1wBHc+dk/7nWAxwHtfChJi/Wm
MmnaL74n3wymSHm1gZ/J04GuCOSqooqxHL3lFJmcwP5+yF6/PRQyoygdQ3fX6b+6
BiV0tb8VizGmSRIylMcq5U5ZpIMr4juf15MZ9WdJB0qm7f+TSuY6lj4GZ6yK1dd/
5ZapLj6PxTSTovK+0W7KaRBA1qEWhYHo5bj+GhieAXYOgX4a1fBnOF81jVTfBabk
eRm+y0QA66HR/UUM5Z6dXPbyKV6ewDpYR6nuOG4MxTAGJXdMGd894Tv2XCaWC3IC
qQPqYgLlCyZrsUBWUMpEtt3Nc03kSc1ntDPia6PEiiZOLa5gc2/rtz367bkvGDAE
t4wqJpywYLhVmuY0+nUTCoXcSaCbXhuNZUgoAxYcBr3UIy33+bczUmHukOt7LASA
QV6t3NJm+gpDsS8tdhRnSXoLKJ9xrK/2lhXfCcL+NdYKQQslCZ5WtNholLi6ymOz
ZYahm3gP4SJoKQ/WnM3QiPWZ/unA5r8Ix3JKhtPWdbtqp571tP1pt5EWdUFdP+Hp
dQ7hbx6ORFAwgfpOSK3qqGyfRWz+KRckQNoG9Cujnmz8zMVrkuBD4sUKjlJnqoS/
R8RiJWBwPD+hs/E0DeOK7A9JxIkX+19KN/j9ggeP0Nqz9k9OJJkVhaX+LDBBlWxI
NfRLUtpMLt5ID6udTreoaxlavYT76sG67kWMEXleG5qrtRdadrKgd4qaVj97SDba
QbPDVsiFSn2IzH3rkiNTjs9QOkuRFh38Iyjz23Ms4PJd871HEB2fCO+nkzLnqpj8
/tkq3H1pZVKbShekA/KOLXGnNsS8YQERQyS49/ELhdMs3dMUtRjmmBYizkD0aICu
5X/l3/qXUDAVDWTNC5CLo6VHl7pEpEqujrzA1++CQeWCoywYQtpiOMhyr1p4FfYE
q2AEaYJQz8RqddX99+ihApqSos2aT9AMFP0GiKxO1hU4HL48Nm70xiZZvrkepIJi
YUECoVwP57KJdOi6jfIER6YTKEgp8Fs7rDRf5BX77x72S4Yp3zo+Xtr5b6DBKo2w
E8ERbRaZgu/tfajVMHS3vOy6W3lmiETMHWJ0Rk81eod8e+p0MY76VKgB+LpvwaTG
3ZUId7Mkhm43tBjHd8fuzx2o1ZQRmh8/jf7tmD3YmK0cr6lpf1FKvD8NHz3sLo82
pC/R4wksjAZAq6FpMyoDZsF5ilQWUG47yQVgqKjTeuSptrMuFcwKm40OH0XRbU2W
5ZEQXDiL1xqFNrLK93nTr/VcRvDK2Rnj3d+KtTWwXE8VKyMsXd7uEcQsZLWqn470
PEIGyheY7INv0vKRAipSTa6594l+w22kZs/zXHyprG5GtmrRBZI2LH9mcLdGdp3p
PPFAxyMkvlQc1F9BTxQNL2tBs1lhYgfzK9aC3QskkRRucL3s2fCbM0hxzV/UIiUI
/rt8w220DERUArg2xvg1YH26K3zPpf9cIcJLk90uLMNv37zx3V4a8a/3Jymu8xo/
E6SazxtlHSSHaMoLUzfUIst28Ml2eujnuXaY6s5/JzjCbwPk10DK9BbTnW/YC3CC
SPd70sducTPDTyrbVtQORLiT4PyVyOrmew8pyBdPB0H3Kx4GMVDXfW+e5zAG/1MN
88RvYERpD3NoU9gKU/m8RlOcz1Hfu7j8TWLLsVRxlUT8N1XoPk2TlsoaUFPuqbrK
GBWUgB2tSwipP592M55y35AqCVGOAOxIekGxymRtAIJsKZZx0U0OCaQanmXSNhRd
Wgput8aXp/9Dj6HpJLeiJxzL8IbLzZ9weLoFByLAK7PXd/f4SNke/rJo7bz79Z1k
9iYMmsTAFqsl+uUqIKuwb3HVaoMobFrw5x9P4LLrNInv/MM9CosyxaXnKyHsqoWW
/HAHhTttj24tY2ix6duZ49+UDLvalnudjXYihOl9CFTx9Owyy0OgLFehMcOMTgJZ
4xy+ASGtvd0D6Xj8ZRXzZg9hVR9uLm/2wJfDsWb/63WL/hd/kjYNYwtBbE44GDgE
ItSieL62zCu9SYNZJ2UkhDmDORvHuKpXAxLawu1kIVCf+RwwNtQdhW877urjupZX
xgtoc1I1uUTLJnyn8xTquAXYil/P/J6tYcw75hk0eTDOr4PVAIDT1UWhDY7iwVSO
stV4mJUtrGcBQkgrMKzWAI+wxtEZHDpAWCF+0pVmEf8izwnjPnOLzvWxKrWIrprF
hUd8/aMJPAN/B+/gofefcRshY2n2vbcgyLEpeogFUYdafJqaI1Rw7XBaYPtnzRWu
FevOAbcRgZu9mBhG3+Hvnj7N2DqgKcDXUNfj2hs7PiR9Ai9yduCKC2r4Fad6z5sj
uNmLMhjEcxQs70/iH25h3H/LZm5bjdIpSxJSS+gUQJET4Ap8yoW8Jb9nhEgVSsk0
Mp3JmIfUyY1b7zWCePrAMsA/m4pEnY8KCTuOeG1b6DfTqA9ThQscOHQacn7nQLYv
35dHtY5aZAxSWBfih7poMLNV0hEh4n26odRe9q7VlihRffyigvmnM58FMtA6pkGW
Emb01FLsmLmYuZNT50OH60iWvQCRzqkBiLm6aTYrZFqPYdbaR4mto1VZYC6ArKui
UssLMK7LYldarbxmR/M7ohEelbe7ph1XZABc3qbJjw0haKcNQCF31+BaS2Gis53U
30icJ7WfGlqcwi33riK/2HMwOX9UoR5+XRtaSPch/A4SbesJmUdn06Qq/zLqdmXg
QY+3SBg5hfbeMYDu4Hoiu7M21h5jWai+yy0dg+azcQISaf8dCaM6Q10JZzrZT4m6
x1GVzZDWe3pjW8QwyS13W2wEU2IMcJenPkM0hySvbWcPqOThaXvjroODinQbuR4U
K3xQDEBP5matD8CTDloiQG3dzih8UJVFGfKLNXa7xvEFQqncKOsGH92oR1SH0/IS
7/6ne+yitGWtppxA4ziihQKaTDEFhGE4Nfg9UPJehlz9ROIlAe6IAITRqpF4EJus
/Yd+2QuWbuul5AaoNHvrqo2qL1enC6im4zZODv7m3sqZMMCBckMGHftGpgjLqkJU
h8lnsCsYkVYCY/JwSFz1YBXH/C2lfjzIApP2LnpfbMHyb8rUo7DsBRpW11RGy3Wm
glBeYAqlvNoJVOKsnRPzzn6mCyw+R5RkFIxrsTocMCv2/PRn8iiaPG6V/X059S7N
BSaps5NQZPvIJObWMukrhRiv0p2bmNuMpzlIbfCEprERYlxpfvXW+uNe4JxUaX97
tEWj57f70jLTQETpTgZ2cnUaQJjem8WHMk/6m6BF6dl3HQS+qruYBOytt+7jxfn9
0gbd/WXQidrt6PjmMCYHSOvw5K0TNUU/riIjSCnJ2c7k/cVIRP4PyplLPGwJ1lfk
kbtjdENsH9SaKJi8n14MALq6n0w+IgsRa1mXeFJlVOMqHJy9pWszwENEaisPxTph
r6CHRu6BKG9nxqLoAwmVUPDh0aQfbBrhRKju2/Kgs9f/eXM+kB46/Dzp61mc/fMF
BqoS/XVm+XkhHVVmjFeRzkYGfm0l6BKoYMhX/8GKxRraBNAL0MFFS1q1O3R2ZMCT
mSZOkbZ5KvLFf/NeqbJwFPiShdwH4S5L9MpvBrPz5uw7H+VKiIUyLBg7RrWLxTFI
op4l+jvjH/x7diGYmnGBSn3rQ90bKwwspuhN8zJfT+baze/ooZCA+cf/v+nJGcLX
res0zqMZNylvrG2HLj9nNPPzdnqGb8O/urZMOjL8ZYhXxb/H63OyogMQPqOsONND
x6oPRonjms2JhHAJ8wYEAyKVSuj7CxPA6TZqaBhkRwRRzLQolOXqK8CQ+nNqrq5L
qptcuASpZ6+hOyVX/4VIQmBXrLXL511m1qdk2n4nv3S/PgssRt9trCwql9ktBYMH
KZiidDUOsFLG86WlUlhzvWUubZiQMM+llMjJo4SqWhAhPFMcoBxB7sUqdtotMCpo
EhGZhAfVFli1Mz+VFtxiGpv/NtwxvQOVzB/VMs9Px2gfwdf/Sae35k6acP54brC0
81ExBnJNHpc819tmUAmeFOviDWEv0yddXRGyxREtKayxlNEKc0xo+F7II0h1sH8f
0NxWFzY8AQpYGsUBSYfee09i9jw9RqXJeztrMDCh79aEYWj5NmNM+WwlbTraq5m5
sqJhZJCQhTM0EFdc8AzfjKXHtasqpDd9mhcPsdGjkWAb8nWiZYOLlJ6CE2NDR7at
RK/+hhFNa61SVJVg91U4kZPO4Mcq+Ztjd5ppZgd+X8URaLdgZQgiHFRldP6aHTuF
DsAvQVe9dvEDFKxYJcKwNSkg4DoozR/B8Jv7Ff5xxSXqSAJftP06a6mW7In9fQlQ
EIZfqKJyZoIvAqVSeWJ+dQEFojKYLglVKvBxjMpBkLvDmfHAXrAvxFZBgf0yQKfX
wjHVez9hiosxBAkfHKqBSn7JAUr1YsqWo5NKljdXxLHFBjWt4rigMCtTHJtnIR3n
qLlcW/Onas/cYHHqFlhDRBCknZV3Dx0uIONNedFpwSWPCTBKXlh2IugbUF6ho1IY
Vk8hYwVAsUjCaomwzRUp+sDjYk9ZuN4jtmPNC8Xu9UfB3b/YQBbooPzCS1IgcYEh
xkfdBoD92siBTUanQFClBjYKqH8iqdtaFtmnQWjWu/uaEEzcH1Ypckx3oA7uRGxi
DT2SBFc0Fc12468W6Ui+cj93ujGCkmEPHHyxKAka5QdRHDxroL962KiadyoUBNQL
3BBR9I43miQv+6cNBQXeIKXWaMGGANQ0fdm0bnQVcGHeFS5cQbdh7iyMlzaO7sz/
cR1B0seWy6Ekifod+XsTknol+l4nRu6wHFxT4OLzFNibwxZcpSoQonK1Oxzx+GX7
moQuT0OxuFxGIivFHvOCsOLu3tlUR0XKXCfrlSstuKmkxOkFiYA52WPAYJDdiurF
UMuIKSlqj/py1hRCPFGXRKXt7Ns/LTh63AjjKZu6pvEbmbEbJ2m+RF/VqarFeflr
tu89bJj7An5OJ15VDRCbX/urRYKxAtytcOg12TartDeKdjQ3baf6hSkFhKTdR/dM
Sez82fxZxWlgp/JPHA2rqkz0a7YW4097B88cFzslYDR/WuB9hNQ8bmb6+BEcKubR
53vB7dJb9Wp8uGIQA+OgJiG27W/UqoHudaB+FpnwBX1BlJP0mHtVFUgoZUCzM6Me
34xVAT4rK9x3miI9uE7f5WfP69RjPsw+iLwM8JeeU2ryEIjE7hirJ01Bc1zVb7bT
MgVl88UuURd/w0BvQ5sx3OjewsIKQ2sFCr9SNXK3+wqaI1Ie/W/ah0wF+T+/K9ye
L42S0a6eTNR7Zk3f3Fx4uUhwldVNdaSbgCQ2iNwLhzUP74hbnbl7ZrHDXOi1Me/G
spqahwgfxl75HXzoUMf0Bu9uIVdnPDhjSw0odpNgCAddIOtFQDlGGu/tnPeLx0oi
VdoPqcWuqnMroGnoPOVJDh8w2IAc+PgVbxyiG7jCUF42+ACNy1smXdxAfC1Dsr9H
d9TQXCVjE+fBJm4JE79bAvD4ZsipcTBCHeUxkrRqHfHPeVoO1skq0Svzrv3BqNiK
Tw7okwzdp7BZTivB4k9QHLlc7VOnU32SlM7LHd3PSRPPKEB4+CxdEwt8l581srBw
lD30cxm/VM1/dthxDjRh9TJWlLunlFZa/Vfl6Z9hS91XJL2Jb7F5wXyLJ6vqdK4B
W0N9+LiSRQNUxjJr2jpP/lTQDG515dtrK8xLcwf0/ChGYFK70poe+QFDL2+vf+2V
/WH7WbZdc222/XawiXsiF/9iGNSjtbtSTYJjNHaJQ/8IKPlxUflhCFT1GIicqkPH
aynUB1IrYfbjXi0ngwkt3pmeN+KXARbWG0utUO3GPL3RQ1JKoVlV0Rc8AwqHT1Sv
VDwhB4TYUbxCNm1RjEHFYr6zqxK3AhAnOCIgnyschrBxfnXW81yHTzsLnQXRXZ9u
jY0kba04FTBz0zXdk8DP7Ktd+qzvHB6vTV+ViUjCTgslA/LMWuh/ZorNydqjPCFP
8OqsyQB6P1mWRel/NhH1jYf3l258igBZVs6OJzz5rvl4ZlyaOQjAaYpyBmmPXYpG
sP7HWWC10WORlYE+UIIy/2SbjutabBmO3t+FvIGVM8Aq/C4KktRfP67U4tS/bcEN
Intal9raq6s2GTNwvl8JatuYtDFv9LZj4zGA/nCp3bCN9uC2QXLac8p/8BgObdqn
ojLqtw2O2BuD9Xiu95VHV/4CpL5qwblmViwjxOsdRHW/HZh4jI+lRPiGbeMJh+CV
fVSW+X5OTTugGu2T9jS97UDkRoLgX8rESZr8dSwcx+BYh95x4jww7SgV67L08YHR
uzDWkyhycgFQjkc+m7k+bkEJI2jYaMNW3ZEIDDexyQhJx8JTMlXNrZuxoUC3l3Di
tCjcTfRrBlXrdQLavDj6BlgIkDhwBa0fZEDj9CaoVvCSYj2G6jXA5NcTK95Uxbx7
31SEvdfDYUGMNdpFviFCO+G9bBi+w6w0bigNZbAp7nTD8FtD8lstnHO3J3AI0h09
+z6jEL+2LeaZvGkWOSlN797OmkIgkOvK71ct1WqarJAsrZMAKQi3FgxcxZSHDsMl
8aYz89MuvwljR1e4TG5DhkdKvVTweOPAQCL4SmhbNdnnzz4STSmkmGNFSmCTR6+t
NPYxo4oPJ79lDMY59xDY4xtQvLcTaIkmcAaCSQm6bg1SfvH7Ej2tCyzJNjSFT83R
pc4qoNQUmHihLX8mf3oCSGUgnUhl/BNwlGc14JJuJ2m+g+Gv6cHMTRU+NTQPeu9O
A7OVbIjFhRHGMWxvbnxVBAnmDDlKYyBNc++heeDmew4E7VfWgBePxrlRNAluYRom
lvho/4yiNwV6RK3uZ/YffSWISFS0Uw79qc7HW/tZXkLjF6ZjkK/KXL17BEhA+4DW
o2ee6wm73QZdC1uEFB8uizQzZvfoFEciRYOh/ybdFLiSWUENIMK15oKak1ExoEFu
7ylR7l4MY2tEVlQE2raVhacaEd4nLfLUfqm+cbuzOg8aT9tfm06ReaU9g5W+aUo/
P03WTgazJsiF0pThxfEBX/In/bKtO6kcjlhya0BCh4TzP50aVtW6VkeKXNth9R/o
8B2IQWf3RBKQIeSZH2spTXiNH1INmW5cf4ey+fOEOZyLnwqmZEDUS9n9I4ubnSF2
K0NSkT+hNIJk8FrgWjmaLPsUaaYrLRU5ltPvi6dpZWbg0Uz/9GFiI7bIUmyESxOy
lApyLm1uXejKYz18DXt6MLrsQumUDdlcUbH4KHVgwcnk6SnyPkZ7EWdjBeNR7Wm5
to6JKJ2M4hpJXt3PUn23SHXQ5CIvmTNrv6Q1ZeUvgq9kTSczXBQEPwtEokep+66w
mAjBMOeK3C7hijtZswVv+C0dtmRqd6uu+VuyzWNK6luvF/OpEnap8Z7jan9VdVa5
qHvGgwBJo5320zjMCgsRZu035LDDAz4mxBVYFBkUbh0O8B2kNq/0FlWzQfkloxQf
geCi9FgJH55JdNB4hSlquVIBUoz+yoEuTCMAeDZd2EzqH6G0dhOv7WgoF+LbbXO5
Oa+nJprgVHuyoAw2nN8GcllVRToUAgIn6lAvkSm3ugcEynw5butW1zyZgNIzPQzR
uV5bdwwI05FcDOU8HV1WUXTywNOJNnwTA9j6n6+Mb/KMefEw0FXtsa8jmudqybfN
E4/wbUCpD/hPLEerhbuUKEx07MPvC6AmWB7P/RMGQZr0Faacuk2ZwpxZDmyVJfjr
E4JWWCqgwhhRli98v9nqCnTwMu2MBjmhtisJbhZq8ALED8Xwwa/wd+LuNYYbvhNW
CYQdkPz75bnF6AyuA8lnq5Q+ekRNMWsMXD+ir4t2hmRPCDy135raIPpIpKYtkQYT
ez5xx1yM8rm/nPdIie2AxiH9rZTwt/idXTjfmlg4pAx9udkERW06RDXkaQD+EC+2
LHh/MG3MZzlQU1rxfMcD2uFexY8VhQ0gcggkOmWzYNwGgCVO/f+1r3fy+QgJU7X+
wgf5HSCvBppvtqRxgNTiiGw4FbnHX4w1qbMKbf+BWxPktMOv+YPizV9yEogAl20U
HvqKX/pw3gC5Ksw6YXeznEHabaw3MhObzfrjcE8VrfGBPmeZ+ic8zk3wKjF65wZu
9oleLdnQ/C1gVQq8VyMiXMorbE8XkBDWRWwixC4Ub/k023Do66JC+H/XJ+NYH5lk
cnSuj0QyYk88G0iAkLyBycnWqiMiVMKdRokiktby1npI/R+zZAnyzP1H90iBmEyS
I5zMpIYmp117RydYKaCSfhdsTfAcHkwwzetWII9BM3xk5zArpHfe9GLgfuREk3GE
kldlaVXnwnYV4ou7exLeouPEi36HjdhI9L31lqWo1M19DGKv2t5x0/8JcWdFdx+7
4iW4pnXuMEwJ0YIBavmUNYcL+vj3jHL76mETdvgpYnNw/r791AO8c0TO+uhIbg8e
agxL1Hn2gYtsGUcUPzhETVibQKkdrTJ4uSrULuKHSsBz6s4es/cFfWAE2fYNUAMv
VC86yn5nufiSjifaL7+k82PxKLZnz1EFCFYysaF8msp/y835IIZxoC3wO5MMEZLA
RLv9rGYh6qahmZFpdihoHP8R6YQEBpj/ioysWWVts5SAgrzuMiaiFKbhDjbQuNDx
i0wpHSC9q59T0QUsVLMAzIAtAt8nYm0Hexir+kcL16sMT6MWN+8KJ8TFknTSXbrV
WrCpKbrHi1kZDCA7zUCsUJ9pcn8BIKesNX6/XgmDX2G57t0bjv38S98Ogdft/KEv
wIJU3fakGc/j2x4fX3FF/Ai8zyL/dRkbVhXlMajOZbLTjsx5yRSmp8EQ4PnZJDv0
R01ElX4rNgh69T4qbuL2SazPkPo5U5bw2eKRT61t+1cb2iVQTqgfVlqH81z/MeY+
1yXG+Tk+xropeh9PEKrorV5It/+uCp9yge9m06orvPnwfNV97BqvP+dDoL88RYH3
kqbJIc+t6zIjNkP0gD/gP0XU7mtFHZyRutgyvlaa6IixjmXghKFJuA6bW08qioEx
849Hgmu/NjjkOmd3NhVMEZYM+svZYmNmWAn/crkh/FAg4MBYTq/dQUuK8aEF3tlT
sk0B4/cInxyQN/MU3C/+z/jFUpL419CpdI8flQifrvXsscQGxdJSMoipi10J//8h
CUrQBUgwk3Ytn2/2r2PzFVnp9pUANsDHVoUMY1FWqvXxb4jg4BXMgjUdoG3futkk
ry6DpIHZaATN+Xb0Qg2YZ7/7qtuMnS6NwC9K0b6s0yaBbZlW6+O6GByddcSbqb4p
7+rWejaeI9hDlOezIqqyxvQIcB5AonlHzFvqhG5skTjXe/9yqIVoMikvN3m4HwmK
xnLImRLxNSqCvb/nmjapDkfaCCS+D95lY8/2dlwHNB/YO+bME6rVnRvh4we+qTeg
pYkyEtbt2f3M8QHL7c79apHQgEoBAyiJ115Njo96AJY3zPyDW5/g7hxBcBv4KVD7
Ny77dK9s4mEaI53XrkxYyZPrGqwLltmI32no4C/3hGgvcC0AGIhsva1nhBya5hiy
YI3NW+rB9MRMHGpYLyc1sbwWMPSa/UshILS8nqKiC5wj1jYfn/km0EjxCaFP+31t
oDkJqCv0rkIZDNUSD1hvAt4QvBatR7LPdz1w36p59gkOACRdQqfbZXERTFnQJ8al
d4pS8ZX1t6dkDpjZV31Nb+zghWFYo8a4rbfngvvvsYxWpJ+LPE0zg8GmZqQrYOwT
wNQmhio9aYG8LSsEER3SvTNd8VBeEqsFthY08j91gLAkz/zQ7i3NNsyiVSOPJRIt
VA4m4f9+h/crZcelJewKP0WiCZLCTmhCpOcwXJla9dBWyKcE8/fg6rfXWmgD7wKj
bPYPPuglnJxufpknTI5PK7SpnSZZEupU9n/nIGWl32M1CWRnPJ0Wjw5MgAZZySDd
dZVJXWskXcbFd+OlfwR3CkqcBBqQqva2lXx4Kg5RZwJw/IIIALu4xG8WBXRFpQ4e
jsHIgiAd5z17Fsobb59ZoP+2Q7YSs+pizXw9tQZd5lARdgWra2iUiVxo8Qzzj+vP
sy2vvObS57cOjq0DFhZQI87QmnW1En/YIlNVwNAPPZZTLzebEf/4jRAkRMXwLoHT
GRy6D9ENbB87UKRUMwcjVPG987wNeEi8Gwju0R6TQmR69oIch5zAXdl9inhAD2Vq
ZMiTolStHWNxjCTkfftW52CsD/3PvHdXEAZPTwiL+a9nNBjSuVeJv9KbWAJo+Wqr
2i8dPRTr8U4mrsJpgkfdZ0hDJTU4tng5OevRopqChEOtndEsZHWFbaevsfOHJnnL
6yMSn59RtLzxWf6Iu9x1HwmyIEf54lAu2hHm8KZefRT+0/xmSU89cjjHmhRBQEwi
mI63zY46HD7gK8Aba4nZT5qUE8GNIls5VsVWmhFNQ3Lh73jihXqNk7QZrXMzsnvJ
hAeGnQWTodifuZ3zVZgg6mi8k8YlTmzjwfn6I8YiGxksfZqaUoxaQ8FLRHV0iH58
0cGzb/pzdeTDYHKrVD85c/iQmwl8k7PjXHqw23EpcBFPQiaFHuxcWOUNSKuw+PVa
KHnBwthDsDo15REh/j5Y+h2JqROaZVRZ7+zlZwdMuvyPlXqk27ajTbmC6n5yUj/f
cteRNEYe6oVrFpuqjhbX9Xlax0lEALCwVeBW5OAirsL9+JYfMnCQtfN78ZIf3tiu
/gb3pi7UBqu5LMZhheWXQBVNrjQWDqGioIfn7jnvR94Ue3Mg449qc9eEQ1VqwUzN
JpNmaYjF0mIjtkhDybjkJkzlvLldFxsba4RdL/HhMT6qC5GQBKk/2PYDepgt4XmZ
qGCnbO0Icu89Nt7k1qgW0b5lWxnmBCpzo0GSHx7y0pRWJkaGZZ3OrZ78Chk0frqb
UROiYXtCRgLjQhM4A74UeEe9c6nzz6ZG3BulXiA7O9wzzEPGmwmdykUamihgPJS4
uxqrnnMQwDgmaH2eRgApN74lBajkz2AFwrPt7pDlE6ZwhdQM23hzFEwJlb5zPayv
ag2vGdutTAChoreisoybvECIdWdLe3Iosq9MDU6bz+ai2NofaR5zmqrBA+Kkj3hP
ulC2JUDqBi3JWpRlNfkNenRfALmEZmuPljvzfrZZSGKIm+tfQ9H82bpQ81Jxb1Bx
VmmOadCBjqEMLrCQnCmsOeCofcfGzWJH7u6eImNxxtY7qZ2oGZEWFMGbV9iVRWBG
ZxDiv4uTFToXibvNqtMcKYfjmgC/LOarDHXPuLY7+pvN5xOO6y4FNLYE67OHqI/L
CoEzyW283iEv1QYItiG+bq5B+NO+YpzrkoCsdITOdHZo+Ctc0bAbcTQEb8cAjVKi
IlVqdipk1pkglDILrnuCUqq1UDhQnT/cstBtyUCHJ5A25AL9TBuycqaM/S/cIIt6
zS2C+4yaj59wypeCBPD08IFjdYFvG9+EoynkO8BkDrJPJ+qJs8YfR8aGD9rDq4hZ
BBb7PQpgkhEYBNBDVz8llmIUY6OSRupAeasIOvyPHmSrjfc0QzdJJWu1zhny7e2F
F54gxEsDnclrktvKsKmvY77SvH4+DFf2txekAy5JMqWSpRB1G/FajDOk08eKKFUZ
OkDOGRQGywtzmf0wPMXt8plYxa94ba6KtXsiD2er4fy+yX5UYHwEs5UXNopYAPBp
CHmGk+vyZf+Fh0Gmxa596cuIsHRz3Qs4UN43uu6QS5fF0xKLUmYTCpGQ2CZ0FW8v
sUjRPvjmm2M7AzDZG3/m7LgBXBPjjRZPG6xkAmzD9Lt1R9REs/Kd66/F96Bi8elF
008djM9iikcm5n9bHx8JhrG6BbIfJ8pz3x2d6i0cGSbDKA//QbplkwER/nFvucSy
yuiopMJlIfGYsrG8g+Bfj2KTpgF3nhIuk3sm3J55HZkK6C//9LKtgEBMaIjmxlr3
FI4X33ttMSGvMhqeiEIh2d6bAl2g0CLmUaHiZ1mFJobdYBHhikS9mHVPaHIlIQ0T
22IG55y3whEYN4jNx6MJjrgZh7U92Lm2m5qvisPMCpm+Tox3cd/ivY+VfHMXTasT
7sMZ/aXzAzBAMBlC48cnf3v/0mnExCrhgPKhB1f7KY4efrSPcNMGs3GitC/p2/aE
3uxXcA82W1aBeeLBFdaglQebQUbwTVlaAmFY0LLlrHYibCWZ8QzwG7wVtptjBaGi
RUhaINPDW6KsoNYbDeuqsBDydY5xaEmzR9wy+o0CiWz7oreXQPpdqZikPMpV8s4b
Stmmza0MClpFto/1ANsGfHTRNxj9IfM6iM15QOdIIi0SJoKLUo9K7vUQxK6JO86T
DerHRspgsp4VTG4DGN0Hjhn+wv5nb3dogP+F6Q9djM9w6FNGdnL3O9r8zlCX29+P
iFznOwfkCYXML0mwF81GAWdfu0Mi99WD/Sc4gDLboSVcK5I2SLDVhh6U44JpKfPP
htNwgeDysy3UmPTp/wSU+BlZiMPDtlI36OVN9atGMGGiIPMFxZv3wOUghbzyDZq2
beFXf3B8YwtdTvi4pTbkf6UMkc8kCz/6JVEbZkmjD/aInu4xGDa3274Pf1O/ALBd
c+VVAkWFhmM6AOFOtbaXmUWnzrgW7ViLUA9qXzUJ3EufsDCtPdcaGWQL1uMeW/9v
yO4od631NSUt3u6jTEkvjHnfYRoNF/I9X689DbbGr+WzSJi5cq/6Ja20x9I1goPg
7AjeOzV0KrwCWA7RKv2oyIW3wuP3Ns8DfbqZhXihxAYPfE4tVNYcnw6fJfn0tBeQ
ne28GdcEaUz4w/3dIp9ZsvJaKRKiPbZDp244H6jpaG4h/tV4SLVloKjDglH9xHBL
bHJLOnAXWRjP2BxDBdTx2Kfve1NpUipCYyVHUAd5gkEd5kEHzGEAC6oK3movZPv+
NY4fBDxy++7ZG1WAdiGQYqxSRnlt8IDGYEzwafsEkb/AMbCsQ5VIiM87QYS0VMTq
/6gG6EC+tG639NWDN3Zs2CIe1+RGRo+R549082RbhUynnpW6+YyQyuW4Rqc/9Viz
Z0IjQGT6+DoEbDywfH+o5Qu45VF+vsEJHtxWrNfrepjYSUAsllS69UvoJhruenVy
+IY8VJkczP0w7NI3IxbQp0jsnPmmCC7ujTGioCEowD1Re3JK4haDnnPbJVoPb2tK
pykGmBjWsILsi4TbpF17jDLnXgX52SEWBKEhbTsHwjz6H4yMmWIa1TT/rj+jrsR5
TrVthYbM7AKQLowO9Tl9mtPOHn+vZNRwHj0xEBkangFJ4hMVbaLcrfr2xsqgiFJg
AVO0wYvkq7OELwyQl/8Kr74ORvoAAW4DwX6G1mDXgl/meQTC22jdw7XcGsgcKFpy
7u4L9p/alVM0qGeYn6C9I9bcOJB3tEHSG6wpnhFG75W88wj6WH7YY0sOAWxiu3Fm
WtNPhm9o/41tUfNwq5Vt6+5CxIoODHuyJ9JjPJf0tajaREuUWKBwdz3FORuH++7R
RlRlp659nztazijHRl/vG87+/4sPIdO8WA0DPlq5BhB56VATjKYfhiE70tPX9ejD
bqtX9Vs6xE/Q/KOXfLqaFr+EIH7YXrXyh2ZsLmHbuY55f9w9+yrLRa7kQjIS8Dfq
UW6A1Saztv2OjLV5e3YAmVonaVd1Md49HU/2S868AQ2/Wsrt8Mvjf0n8ojQe4V2d
vko/hAw5C3O1VwtFAhRSuzyBYTRGHWRCt6LFGVFNqf0GkIj+pdMenjnlfdydMNZ6
s5M85oudEEJVrr7NBPD6ESZWuubdgZlXlXW/Rl7bCOf2pIrVosq6EUxjCEmdKzp1
sXhvCdqwMnVp35/cWOfWUCUsUvut7P8cbWKcoLxbXEPE6OD8HeUwkE+630TxhWCa
TbDo/m5d5TGj/TdurnSvlgz/Keb4NPSHFD/S6Z4JoUDI9PGvlMAMjfcfNkf224HT
1hQgoUXwHdGir2k/YvtGqqAmHST+x5hxDfcg2JJhkQNd+2A3BRHqRfFK1Pp/QY+7
5MEu4ychQxLyrqTs2P/9bsxHVBVRp0dJr1Ps54sl/K1XqkdzW1wFPYLaEmyOj51O
/xp3+X0ZPgIuSieXcw5X+SZmmnsKaB8gjvNtntJL/4Zo3gTOjc/viAm/NobhWnKg
q55PEktTOr7zTqPzMuT14XlvpEpnbGSaNqTntFyIJAl4inkRMI8dYWreKpVYr55B
PG/DDuIwvMlugscyczc5n5yE/28hs1O6PVIyAwcgUBxmWucJboQvphz/nRXAEPlR
hJi8n70kosLk0VnGg/22Na+aF9DIFt0CUM+/cBPVWvpvxtygeiW1K3W51FGsIBYK
p+ZQSPCoxp7a63vVu552NCvXyFNNN34wRgbJzsuSDrdWtFqm5c/XBfh2/eM/lD+l
KtpXasd8tV1uCgiyvtacuvOUCMZYETmaZD0gGLhsjVLvTtOKmm/Ilu+XMDUwbiUC
wKZjAIMP0hM7+czxFAVsGRm4sSGIzhvtEqcK1FKOZZoJj7mBRzUgM8q70+WQrmAa
suaSPrMLdcr76+0oBCfG6lCd9EKPMW6AKSaRbVUidw/GtrSxmSV4n+wBUKskw0Mf
UMdqEsDAkK/3AxQLWSh9jBFDWGHMlvA1pBFPko7ca3lowvMiSLk8VGVfNHcsNKyL
62UoL1jKNXn2sWMheEkjDOPkRXQP+TZQr5SWEGuYBnyBaK0ukiE9gis5+tM18VgO
m2Qfkk/+mcGhDWf8oGZrISddGHFFIzlF60+WFSroOd5XT94O2d81MlusOFqLK0U+
n1SGFchNwspc6HqDUV+heimaSzNlBAq4b7dtMRyk/0fgOze2UcwZriieWhHbIH+A
ehOdWutw00t/Ghp/pkKdqXgK4rvDn4KeHzpFrOoLVDVPvCTZY3DhbKp2Gi6sUMV6
fmpcbY+p9++hywU8Dya9Ts2ZL38/etCMCeyPdx0ySTT5ykiZsGXOb/7kDRyDqAPh
Wry1F/V8lKcwLn1jG7zLpyO3yxu/+xkIusIQeBrkBcEXnFdzZFn7x5WsgbSmN09Z
8w3abPrYoS1/ZD5OAhYKWAw1hlBwTU09jbHHqI+w205iGL0jgFZ6W/+gGm64ry83
vBDrlVNET6jbWXSzfNHUaZaWsCm4DTSAQczObMhu3WGug53hhsPO5xLvhZm+lHRm
Rn0pjhhZ7mSrICilRn1OQV8SqlH2+1MYdzlrhNibczoXWJ/mvugnaNMBTLfNhrwC
qjslSlNS2TRbeOo3hLyZ/CzdiFrw+amF9YWNek6aiKyF+Z6T+tJlQzyVbQ7hb8NO
laV+ebCt7V9d3GnC1IDofOERnlAMy2i2PXpp15AVqngkFffJO2q7niSuoepuqVO6
Rx+7adhj3qEBbdNt+ONXbBSSzd1DlgWF7NeAvwFx6vU0S/xtHdagAxQ+sxzgJtLX
9kbam+54a4fwaLBHWcxiWU1rdLhpLNZZJrI4A6dRJVTfe2NfR3pS65OMKimpmU4K
11fHWrFN0zuF6+p9w2DD5338rAcxm/F2tv9HipC4CEFPygzzxPonWQsIu42sJ0Vs
/MKFQoRd79+HbH142iI/Un0rbOiWAHzul+X6vl6VpN7WOtjFriklNY3Yyb02Ek64
y2KN0sreBwytdRQKPNp2fRW0tsie6kAzlTmL3kyQsilt1LlysYjXdAKs9Z5xDBo5
EYW08kVwvvVQjl70G7tqVmKv72qn25WaYeIjW1ozs7nSs+X7013k+YkDH8s3DpY9
ECbVqfnkqlxR4Wbyp4MAiDq/3WYWVVBHVt8PdQHO0oZP8KKm3FG714pd0qZj5Eac
ugfCFQvYSxgp91s+3T/z7R69+0RQdYEtd9z9IUDJQLzf8HKdYOxZvGhAnKa7sfB4
XlGmL8vQCdoJwNd2FPcZTi+5KrMtMdMejeNjB0aKYr/5MdDsJxWuGfrFyrcsaJjD
cwqzLdreFx+3WHOiC2GVtE+syuPBgtXJrHSVuRIsbgspCW3amMPrWG/VaFKalzqu
wpYeRmOgPKq9bHyFuwK+eh9GHn5lYwQ61hrQB40S7R0JKibSD+Ld04aI5S/Jd8bk
F+YLEMm/HN2mx3J1IpWQDltvNTSuYM0X8kmOSplaF04s6v/SE1/hGlnFu1HvWonM
GdwgY064CjfMWg+KdTvx8992EAl+pJkFcSjxMm+metTWfdNXFNHbRQhgqcH8buch
BWSj45W0k/eMJz8wH/GQR6ovuQ1kL/KvzRpf4GeNj7gRuGlBtX3WHtnmY/zkTmH+
0I99HVEuYUKGFvZHfg7hZCUXYPCHnoa3XRQOYOb6hFjhPS2A/xcRq8fD1z3iN9Sm
lHpqXvYXYoFfCg3ZCcTdMqFlhD9VVUAdr71mhqSEp4ofjY8mZ2Yj7PLp2eWM/prH
+T6Hh+fEvv2dtBpMM8suXgSxu307A7wgRVDF1gAw3IFfFlcx+cDAbeEAOD/u871D
wQ/hlZ29wn3NF/fD7hL64I4lWTjXxRDYGeNxoKWj67HWQQ8TV1aJssC+LpjkpSN9
YHHgXTCNQ9INw16gO6HoKHhQwfmlFqvmYmNJoleNo84QvfvgFIrsNrXQJ5xbvotr
SA23Oq+/6hAWHAo0B3kZ+AYed/MptkXnAvRrLi58sgQsRCgI3hj0v+mI5eXDieH0
MDybnzq7Bq5ApUM+xzQ6QftFVB9bq9xORKssorBXkXN2mZbPJ2uK4Fm0h1dLAf5/
3D+V7RQvFmLARkYJ0/wZP11EjfbKJFq/Qi2dfmZvApMCNPeUXOq8Ij2owP9Yx4RX
/fmpUJoYP+NIwUo7BPfUa6SK0u8bxf9atSCibyjL20SgpAxQ6lF5eoWNfUp9jR94
oqULOP+yb8PQLAO81M3OWXQMdGtCUNbAJ1L+89d2Nl7ClQpTI9GQV6zfPXlnIe8R
4lYcljWwmg3EHH7Ax/CBdU8nkyfqyvTiIms67tbp3ijn2oTtOqAwrVvQV0y3AEnf
nt7iUZHd+CGGwz97mxcaaPf3iSEWtPaZhDyvWps9FigQcsNtclxoMvWPLIWFEuZf
2NTWJRkQbIxIir5WRFrzETjycifWb/a06NfGg14qAh8InlnyPPgMJ6wABXgolaFE
LzDfsAHBok4/DmrfgYwYu/1jxhSc4hCbFfxtP+4+Uk6S3oyEcBzhOKj2eKyPSQ6O
Y4SjjNZVv3NOIPsYrtJUOeUriDUBQMklHfRKnkeG0WONsTlYBQG7luLcLAuD/cCx
QSBoqzp14i7nCPKTL+XOiufx1bkkw3efxcyRPGiLegCDe6bxZOr48f6EDuTnpL+d
X+kgggvG3tTvAMFC7J06KzOkQ/xSmvsDKPNBcKCmaxYwf3saImxxgKAVdsaSVOcZ
cT8oKHsPoRapsyZKJz1qiUAW/0y6XgteCMHxUzYH4K2vk5UH/m06qyTpHlTZJxa1
dLVmwlKceaHIvBq2SaaGoOVHPZU9/IXPZZ2vyCpaSSYh67t2Honl7nSHDI3cf64s
GxwJzCLYAcvJjomQskQEftW61VigO64v8/uWybOGeT4FA29HjiMZorFs/ZrkmjVC
6+ZuUBCtT2lnxFkPvxafuso0hNIg/qffbQXAf5FCEQHAPEgak/x9fQTKR6JS1WaP
ArBKMLpvApdC6iUYl1Qlz9VR0iiWlCiQ2CWDb80FeY2BA4hiuW/K++0ACOoew1pT
WS2E+yHlyo9EOdK8eB96ixezD0xppk9j6Xqpo/OSh7yJIgkM3ZWQIYHJp8diaxle
QlJa57tL+fCd3sJt38WjYYoIm3QnPB/yw0ws4h9aA5PJGojOpFzbgWQhEashZ1yQ
CALYf9wkip1QdKNiYSDuZqqqJnD4wzq5PSjOElkyzN2GOJQSWXkTBTv7l16PZFDX
l6WGF/co8IpXwqX5pU+CIZA05RJJniKiLVajuOPoA741YAOTX/CArFdBEjevmlBZ
4b7W9Po138EXxSjpV7LUdo+SHHaXADwxG/kSOKV9ELcnZwddcLdcdyrLJQ065RhZ
AyWA+Nkh7TOWa8PoI5Ju9aOKMOgkiLQTcMegcPaZjGV40RFTi8zfbKRZkXlu1gXo
KSTbspNB5XLdcg8vQ4ufA13NR70rncOS1UEw0EoHNpe7UyXpSGMSRsSS2yLfnH5d
VLYXKlMLjkja2aoOuUCZye7FGaanbthaMDUEFTvoRqVQ24m909YYFyGHND6yzbGG
jC7/R++E+kzRKtwO4dvSldOKoIWdZAwRCABq+SBOlwKB3giJ9L9deXYlGzyRdOYI
KWgfYXGpHpIKSZQdkTih528BH+zwdJC2wIqcCCbCr/iP33vZ1Ij66vf8h1/nqVAq
76bmYrPuQEO8sOooA0+WFOsMcK/hWZP7cxkfGRL++x8KtGm4XTVEGcafcA5jDnjD
Uo6wnbgcVx9LqI4CI6rJTGjR94Eg+CYN9Kv/TSiiN8as3IKSgZEKh+n/eK/HKeH8
20tibYuF2dPEbGzOKF7WSUdNOOkkkxIb5mDXjKeMyJiMPLa+wfWhaSnrdBqVNhkA
YK1mgx0NDdxRYCxmwKE2c6vvpBLa9emGYFNc99GLJwV3WjEPaEyAF7E0nWJwmDH3
qH7OQ2UzvqyZS5f8rQHadLi5TIzeDOsmOtGr5G7IpFY2Gcs52b8tNRRvgNQT5iqP
60U5mBKDU8wRo6xJ8/s/wUcSN7K7cElH8kPHbe+Bc+6nRDJ1IxIKKcOaoAjUPZ5a
hIio95SQCmSSfPf20WHPCwESeN1lUEty7KcO3Qd0fZ5nF2wtlDC2LjMsQ2b0Rdrw
m/vVY2R73sufGNtN7WY3ubMDbPAl82OoD3ggP8x6j1M/vFIkevAxhdgcDgKp49JR
q14YgdQfuomnqA74AFZKIoV4+wjI2m5QDJcgFaDn+pwsdBGD2tLdsT6hlQMwurN/
GywpbbEWb311nj8dcpfvBTxxSZbID9JEx1znkLyG1yTMroamxf9VFfcapub+Fpy/
78G65x1y+l0Kd6hssMBIzEb2znfTGFk3guoP8cMQlGAtmSWwA+dfdE4/Z7ztsT5P
3/kCcwfcHA22RN+SWUviX0UvV2/J7Fvvjux6k0XAbcRvtwrmucypGN60rs72Be6D
cK00TZI7dP8Z3lwg9juqc0OKUpajB/WJ50s2C8bNqUWmcxjC00q2T8FwEhJEDBD5
nJIe3q0rW8IgOyvsJQ1XwYHxwhNv+CMLVcHmv6az2Pij9vSxI64aSx4U0D74SXAW
Sy+A+v0VWSjhrtb7NpSDNrhTx0eeluckUB4QY0leAa0X6FH+U1VCihoeL5ppMHYg
9KDfb2skEYHG/p4DnRQii6gbSPiRIXOVZXBPhSFQ11UfyjiuZrlq3D1fNTkvYhH2
/SKC5fgGgwmgrgbu4Zf0Bau1QUwmX5khq12rnALGxw37uypf5sLgvjDA7U5WUh1g
e3LDjBEkmYTofXsbrpnbFEkGMiyY+9MOL9pIoFGMV7E78t76eJxNuw8F88sNlx93
K68DTe85DIZa8zzePYwUQ1gxtPngDVRGfjxVfaCZvh039VZkewpbN+OQ22qfzzLn
YTjC9b8l9RjSwP4Ghc158R5WYSvSMY9LdBKjT4R7HeB4O8aS9z36ILwp7G0S7Zn2
deifX5VSWHc6eLSxxiMuykYM12VQ8O8l1Kh9GIqRWrzIc2/HX52vuFMRdofo0t9Y
hjhRJlTmATwIBmxNLGwYmI+5+2DD/74paEvFGou5XMYVFjMGGECnTgbH9X6d2UQO
kpSNJyq2ILjDcEFpGKHXvRFspWFkity0d27kcssyrS63ZwXAeEQAZ67tuBYLTiFw
P12tAHYa/eIEJhPzxjG76r9NbwK7E/wfGAaVj354RviA9RCJ07AqXAIGyCzWTBrd
KnJW2STVmcafOWSOqssDbQu7qzDOeKXaR9Gp6VEZGbYtCz/bZxQRwBauHWeGMoOu
VEPv1jh5JGRO9d+ENzU8nuYpcjLE172GZrFUjhAXKshnKJNMAcV1jfqyLsTLQJ9N
VDc2TeXhOaFw20Jt7X7XFYPnAocA7arsHMymASzOuGlnkVvvk6FjvVIE+GowbDVq
OHf/W2cbgq9dJGgODIV7nbNk2dhCwrp3w1Ki4k5fA9ifHlSLqmpPLNKAr21HKxE7
245G5ER80N5ji45wh1Xv2TrpA3W+JCoLdnp6Z0uaLNe75M5GOhWdSt7E5avuJHo8
LxNwqDDheQk823mnvACAfUZ4S1NTxPnoLMfYVorLDSpUP4ABlt1aLlzfCFX8ntVA
l9ilshn90O55yIUc9ebxfu2LN0xWfMmqYyy2FatYGSL27JeEh+otdi/2Ei+gkoBQ
oMhQiSLYSfB2Xc/ApWvC+ZWYVs73IMzPn3m1cK6jh6hgqPUFcSChh5QSl87QIXRX
JpqykgSpiq4H51ftq9Lvaii3OgrKj1Bm3Grby01I/pEDyofLtm1oUUjXBH0lPb2G
85tMkhncOx1SgRYWyf8sn8ykkZTwqixjhO+RhfQ+VxHgUA3h0nqeVSkf4HdnteId
QkAyLk/yujWTJgTiH0AOpDqPC6LIrxtYVfTLg5LA4RymNhGFDgMRxablpyk2Vz5K
WFo5sf4gkNk+5iJmjznwJ2bwG0aX3Gnoy+xVRFJMwd7nE9kmnNsKl6ZYJPGTHAVt
hgOMgAqyz3QOdC80IYNgGEcffqTmzkZxudXGs1tZYa94w293dUaJ8aglcsVSByAH
e0z+EAIqxIjWN6RcyKa4rh1VRHePDBHvzYP1z9/SBqgSM6iDKEThG2S9aiu1L0g/
6zff+HMnaoPJH8p5+1pzSk70k7esocmTOnUqcjWcQFLjnbWLiU0gf5TpwyFGY03L
jMV5/VJzIlTsl/gUiVvyLr9HGIoSSAfiVIXpB27Su9GQRhk8rNpIBp6odsD3Q3Yc
wzlIdTz0c8sX0aDg3mn1Sa9fvz+r919FoiXrfNfgZu2kyhvZUjnmDNtSTpXe6iN7
Y4BRUnk14Be4FEYMRdk2JJcOtn1oHHKuVbEE58x1brcegui/r6SdCehIL8FhiPmZ
PGK/zp7RAgh27VZLEu5SL0qMabsckKLktIn/PI1DolYtbD8QdceUR6p8iZY3UjE+
8E6gpnuVqg4HYeUMNoxDIGtv71UJ9JebaGxwZLP6U6EA6K3pit8zpOneL3O1KVyB
2LLojKGL3ldkGAjY6FI2Qaq6tnSeHpfu1vJK2FKi9EsYx+yRQP85hVKFTRnXeZY9
35StBVTbP5yUjH6XgphUgJuFNhj4dzKd8t/FRa+ZMUI7nbA/+lfk9NupNFJjVDCF
DyMT5VGN+0/KGunoaAKmstiOJOgAdyaFYOV5kk0Bqhnh6DKlHPdoMHOz3nVcKG2B
Xu1s4qHoOl1EoReh0etQ+RTCBaF1GtIXltEtGdt7r5cwGD2Idj04rrIZgHdSRRoe
z5ZxAA+y54gLH2JCmrDJAtOFx5w24M/B0GCnRkdYHlvvXgdVUaQdkbJ8bxj55i6w
ntLuYFW47T0rSv6URZdfSFtFDSKCISmiCDNa8tBW6bJ0XUumxTWRdY9V32oE2HCo
IUKoYGrY9AsVx732MoQsJIHr0+KmftJWbKeoIgH+i4FkV0uR7URaVNXXqSR42Npz
045fPGSP1nexn6L+9Rc2+3quGnv8FgVaXKCl5D5M74EmB6SKP4JZuNRw0oz7wFwb
ZLqtG529/Tbc65/zoHyHnqjXZYk+BQJHySMItqU+uctcJyyV+qKl40Lwffsg8CJJ
MCrycr+4nBVRECsiVQ9DF48QXQui8QDuDZYVMvP5nhJ50PIeWPY9L1bozZntsZ9j
yVZ31Nr2iWZBkuiEvXfSZBqYLqGrtDuGtoFZXxDnL0v1njJE4EQAJrJXlOBaXu/y
lneA4O3uDY091wIiWAYPIfzOt/6BhDKC/45bpzRDTFDz191XRRGKsBlpNXismHwI
JtSLCaZwAsQX9XYmj1Q4tOK+Y/XPBUfz2SbaYJuaLe/kjEDaYDGUK2E/XxsZpYTY
nburbnvrduSJVci4QRgmEUFchl8PxE2eiQ/Y5ymL/kBx5A65M2UDsafAq6iNSM6r
ZHdMwzUuiygeCZ5IAu1KsyOnv23uiZW6UleyWLdbZSczZwrWOrPQum08dHCCr/MB
+YaW/xmWDRxi4BFvKJ2yPBQEYvLASWmDcN+KXKJa/TFr2JTI/oS6K9XBi4mlyo5A
okqV90SFDcakVXZdFyqbDQVs8g9k80MjtAkuBVEUpeeC3NRic4CT49a3VZUZTH/D
gWlv8LDzhAkOirlYYCc/MlL916zkdOoBt2f+MMtQnqWtIoN2s3IeQzprRgvySyEd
bq//VvpGILIMYCBUz5agdEUpWEA8AlYwoeDqNvmL8HsHr+De3ympCdrA7pNALYoj
wJ283HbWPH2Ed/30tB8RCL/EeSgoi6TUTbQmWb2n9teUU50kNEmRd/gAPhz6JAfb
OTr1S+ws8A/oJTMZA/ZNabLD6ckjV18TBeV0miGMRvKjt8xfXiF0zZDRJyRXU59G
QgGoIaKsNoBcmKAmkL46KtSwetsbPVhYdlQv+XZN/UailYifkyPjeQQLQNbgJ0Yk
goEj4+9IuXudGkZPnXKGMjtZThEh3Zb7V1hqttYCWBABkln2eaMTjp9ekFI7r7dd
zdTW4rTJfF8eP3HtJBHpfb9aXc3imDoRA0qz1N+m4rurKkmCFFxJ3GGfdazjp+fE
lz3gyKIwOOAFBX2kHQxrrtW5EsjNn1LxuN8K0Ipn7vQENvV4EC0s6t2KOakRuGqq
nPfZf+WAq7/Ik3i+MZ3yGmVZplhZMFha+H6fTDjtxKdYh5gf3vHvD5V+AUOXBbaJ
S/3e8q4sZkGwUreCNX1emG14WewvS/GpTJ1cgGbiz8PWlKesm+DQif6wjkaP3YFy
g/lgRnVCeM3rr28OlLsz9g0noYGU0q3IsM/PtTpoyECchc61emxr6UkPtDLgLQel
brRk1v/+TNkiXdTGi2ylmxR3ndQe8oJhr2Z2AMU9SaHuriS/pnwlaIGdnSFfXKDy
7nN5ZZvzr9t1nWr8EHLD94KPOn5EcoKK5KhtvO4SmyV7AF1YhE3CQ5bEnVfNdPhs
BLFLmXNjvWMPgJKw5XnOjmx8j7ammdoS7ygKcFMcpzDjcQpRn3RUWEN0QCJUVKnI
T3nq/jJFhaBb/UAVvXp1f+pgWDHK1ZtNJtOBK6H0FOcnEJnUs6WyapcwXpq1buEv
TYrc1KLxmEADQn8UODoqZwySes6lJYQWGsbkgcUtCdN5neoex7hKZerOM+Ps694v
m0osb1KQRAjZ+tmpKZEZ2cO/JhVrlvfOyLNp55jgn3f8SzdaFMnAd/WlX9CB5NW1
7T+I7OkB+Dw3FkLBQhsP+I2na3fRqZkJiqC572oIbYKSoivVZLJocqK+vDBnK8nh
9dO726oR1jVHqy3YpsoaNKlbcGwm7vm49FU8h+Ho2v2QQsyPPkQD7SvuV916KDtU
eb90TL+RXqpS0qcngGWuHsuCYcbPuL/uvGLQOQ1UFeiaDPAERaPBWaK4zNyZl+wj
ld9uLRruC0ajNWQOKO0NpUM8M8NCr/x5/5aFEnS9vENcRjrAIBy3BB+sw9VhZk6x
7S98QkFQ6gfGjmOVu7AXsBS+JOIVOPMmXSvPp16Zfc5Msfe8E3RFozBpQ/kr6L7N
h2YXTzRqvpDDdRtq08M82Kr6e/N6YXG5GdIOwy2QSxq7lKiybwqfGFRmMvHubD94
DANQ3jPsBCNV2n8mfcpbKQkxJJeKxetnbN1btkHYUWRJXzq/xUoxWknbUhroYwXP
hLXSur7K0iaEOkixI7ch2QwgXic7FD36igWV2zgQbiXFnkBWNVU7QPBcgCa/Be5O
7i0WPsy1K3RyQMe2uXEnmF99vejgrc9xuiwUFhjODoO2PGwf6GX/WAAAYJDcy7P1
lW9Ha2C4TeRc3YA+H/TAkid2j2bqGJNElDYRm3e9RK68X4NUELnUGYd4rALq35XR
b3rz3877LPiqL4ucAUFKzQsbQRGd/ivOZ0hHxlL2iCQ+pqQ6nd4vilgjeCsHhmBi
nm8LmwhmmtBSXbCqycQhTtORVe1+RH2spqXedA0ZAQmDK2pMeCh3xQMfEMF/1F4F
seUfJb/GW/CMdTSqT5zcz+1FblUFzs23f42LIXgtgdwzuMnrwS1CGU79GRHwMwSU
zkNRzoO5VJRES7xpm6C42nv4D0/texHoxcXBL5eGthd+c4o/TyKE20+m42B/+/kj
oGidS9pwP+XUh1ub9ZKtoAM1fGZmqo6QsdWaSuEvT+a9fojbZp4EPF0ZkUiNItxc
qIh8GarbZ5nab285Gdtv0Amk+R30H9ln7W0DPI76E4EHDWxCyM3YNmah42duX2pZ
TNsPUsswP2jGSc4Wavjt3hVaLXBm3y1ZfdsQfMy4qRFZdHiV9kqjEXYrvgOCQiOl
6yDKWZRDXlHZZg1e+1OnZPT6jvJCDjAVjxjcMTAkNU9Ub9b35TXiVFGxLhCHDt2U
qluh6ZQXvWGCmjsfb9z06hO6wPfY1jNA+I2aCIHK8PFoBtDvdC1EpWnyYfqei/Dz
F8Sg3/Gfy+OyDwaYKhtnq1xtC+kLPrvt69fQs7H6BWQr7ucf5Xc5FSfDMUBRKFGE
/FD2QAl8RXvpC4Mgqio1se2eA5mUb10b3zqdaZpjzSWj/8BD6+oPd/BavWIxhBRC
AMRqj22bIXYEb2BslI5GwgC1Q79V3sU6DiXA3a62+RkHh9BwqzQQO4Mctxft0ZEG
kQcG2MTMLopYG7gWzlUqxsi2VQDmEGLFTuwfBEjLKnoZi4kzlCmsAYdJ9k/nKemT
tP0+bnHgi0KOc8dEOwc0HiywQsmmpp0Q8urgTuOV4QCH+AQDnJaWZttgilk5dxzU
4tLvi2CvyqVNKAgvIS3EJsmivV3GXcZj2drmZ2GVTbCwIDr+WPUNQjGi5ziPk91Q
yLlmpziwlPgNwsoDBNXxpKxInAXkXYUoZXbu6TzYYBmTrgK7DOf/fCDPyU2TD/Kx
O1YCLlfKpZ8e1nuV27kXHADHAt5acAGOEcMiRZPIxmK57LUpgjA87F/vSgdBfWaJ
422wSqPcwFcWClwQ6z60iYY+XTEYKGMM0Unc6bvUUSIZQbXa4cByNH0YZx88OMkZ
aTI+BvMTGOinsRh5NxlcmHWMdGGjAaJV3PhNV/J2Ktc8ukulKaLs/FOhweeSQSTA
msAZnisgcksF5aMcpMdwDuOrQvwuUXbHae12xF9eTs0fyk7FSSJPcoTV9/Hi3tJD
hoIkJArsmOtmAV0Gq59y8w4A8q33aaCV9efR6DAiGW0Z7SGEuYNz8SpGu2TfirMh
56elNctipXt/dRaIZsmJrsTpBcWqHipvQLUM66AsBCMc/uMua+F7T+Iqo8MBwdgH
xTtsK96OD4EGSDmo5FcaYK7Ogt9lHJwxlaGIVIulBT3jQif/j49UH9mnigvUpLg1
5hrpbSqkppnRiiapkn/rsfrhE11XiWcqFTbZcNUjOL5cS3eQInf4xjL/YDSUh8EI
e5UVZCLzwhJAIVMZcviFrSbinOQuX9PwxvlpdmfAld1QVKnNER/EyQCW+swX1hfm
Qq8enCjYRRFbm8yvMNHu++A+JJCblVsWO0bjMPPnpKKcX6qse87+kvH3EbYmhz6K
pHcTF7ga/eJrx7TP6ylRXgw/uTHtsSe4TQZFFa+Q4JfFpg6RGhSL/QdstpXQSLiU
PR0qsCpK5zXlot+kUsAyI3aUGI5PKoLCziSWx1WGHT0ez5s9SaxfEi3QXpgO3PN/
3mX++x2nhfLcVYbs1ILZjG+J/JvZmBekWGYDvTGluA2cngHU1fFy1U19PsHdyrIh
YVMJLygROKBSrKlIPRCSib0a19Bv1ayjAPgqX2ttIaPLirr4HI66i/yJWisgWM/d
PwtHcoM13UKv3nhxEf3rdGvPQEpXQs68dn3PIdz11Qa/JTBo9sZDs0SOszo65Vp/
9iT1qxKK+3PJnOWwMBmndgllKsc8on72ya43bfnM65GalH8ntcKKq35tsbOE9ViD
RUquwmelpci2YUR/M6xU53ybAVUtvK43fykCu5Ujt9JU3o/imKMTWwCn5wcHGlL4
5BQgbU/qBeA94AlwcHlI5DjWOUuBQLz+2HjOT9H/yA4ZX72qodUWrUUn4MbMslAA
RV2T+kwBeezBHpaifuKKx4JpD14PslfFEBeapw2H8SzrFdvEPa7k57gHQG/iCiDn
s2pCPRDNZGx1r+pKlPzx8SUiXPDFSCQHpk4sxGziN5ydV5GFeHlCmvGsocMSKoVY
FFDbneNZL1VQZ1VR8F7dDeAEZ5b1osfCsLR2OusL+0eS/nK0xJLEqB+aFyGqXpr5
t6wqMIwhwMcPta5ZhPd9Yit44ipNgyTUvLvrlfRhGxDmam/fRRrDPIqueRWpRgS3
sXLUSPoF+Vi8zOKy+7glgSbZSzzTfKB0Dzj/IW8aqLrdlS9cAv6boE9/EWJJJn/D
bjfsB2QpAAKUSDzBb3Jvj7rhCOadEUp2Q5Zau/gUEBTYOJbSGfU57etLAvZdPeZL
mzSHPo8NhLD8uC2zTS+7IkSyX7YAgNuUro6vsBpnRhXLFGEwsBZsZGpoZJ+NlJdS
y1bLpQyEuhHQcQPDjxSfZpiuT5uc1oThQEkBhoEYbSCU814o6/euDlOmjKw24ogQ
FFdrXNOpcE/TKL2wRP9seMdnulPa44ZOEVU7eJC2c+kVWVhAzfY1ej+bi8PsPXwF
R2axSmFxTy+qLTbSxYVp5fILXjmZgRQQcbqvvaD64nLRydaMVYWhe0Fe1zpNW+RR
HG82YpFfsx9b/IqNBT0L0s5wc1ivuSCEahFavfDvRGCwiLAepAGp/GBG3of/ilOn
xrDQNh1bN7XNv0lozFZNh2MKUNpOmUw12W4tqYEcty6XNywBpze1qpsRLpG9UL+m
LMuHtARLtIcralT/cwLq9mvzJMBRAsBQcD4kyIfAZ4pg+e8kuDJV/NwHDfJOyUSR
3Nw2p0JYxig5U2X4CL+5XDdrY/hMdBMS7N3DXA/6mXp/9SSZ48jUwGTU6uSlBhAQ
IIAmN8GIyOWPrwObWsSdiSYrodHrebRVcga+QGPr9PRUzL9vjK++ZJLYUXxsopz0
MzqLiZX91uLLYAs8haI4HRMNsofwWZPvW01Ic7xEA8u6IXNQv+Y+LzJRodIvYfzm
i0vXk0tUGbn9Yqar0k1nmHan5fm/9XrPICKkbd18vmfh4lyNuOuNmA8rqhFx9t+q
dAfO4V2IOuzfDYlwaLmuu1ao7kdLGYw0dx8ymQhFpF+CCOlvOvKzISJAcYV3k4Ng
ziblGrsCIH7l5fkTOCbtwGOY/yBhAG/Ss6Jywv2bLQCy8ZEGliP0tYBKU3tZ4L8f
2DCPnSLg32YxiopbSKSWU6H0CdFvcXQcgZJYyRmKhYeX04R3uiqdRRO9BXT7jx6N
isoiEmEQNZ09EnVbn7LbUlBjrtoqVzqZ6zK9dfu3uO+SwsJytWJvyruzDdmOygyG
TOmr2sa3LGNvdmDLRcw5rLp9icJnPPiJHXvd6f+aQnTZefYYT4voSIRnI1jWPZrY
XYFkj2Au8bnidAA8HdKM0kIopZG2Fe4m2M2J+wc4BK8j9S145ML81vFFG3ddnKVz
2Wwn6oNcKbjftWhVS37apizvXgHfdqzpd39Aj5UBHiGBlu0MK6AKN0z8WJf39OAu
4mS7m9EgCVspBMlRBzJw3iBxKFLyNQN5It7iK/Ef6k8mDCYZKbs/Dnk4cYSZp0yw
qo3ONbGZqUyb1zvWZNaE0mLXGb13OGCPsR8uPAMzhlr/IPluS1yRc4WijW2yiw1o
MK8aIvZYvm6QXb/OR3oVe0fT1Fe8NLtFaOfsMVn7nPdqcrEj6pbm/uJMxajtTxcN
KlrwqBOvPdYNvj2XMF9BZYSmRHq50Zrn1w3votIdFsd6KqlKpecHEUPB1CSlAUSL
jjXfW8bxWI9RwBE3TmSMguKf43yFR4zmeKIYjU6tDfqoin/SCct5MHh+CsF11mqY
IcON6AjxE+II7X/lwdnKSXcYSZgQixdMmRR9R9DXsxhimfTNm3+ZCWPCqTCxsiqu
k5899+/h9EJmgFQVXFdaPaUPiUy30Aa9ZqQM0zzi67870g+2TpH0xgU6yf/TN1Dy
WlKbq6Rxxu+IjI/esnqbwox0iJsZfm8OjqG8OOa7zHc9p+HkBJxCGmKzLcWyCN4w
gNTzGp0P4+zuHBv6tWZtmfnXK9KT8SDEfFeFPfgNU0SWAU8r0gTPzRPDxL3PcEx/
ababCJKbG9jn4iCEQ9dZVeon61W4NNYuSldNTQR0SBIDjGRboEvnN7FmXYyXm17z
L+UZOvSQitv664R+5LaJGlJf6zLfDcYQojlZGW5+bB7fVIXxdVPSHfSyjHjy2ppp
lx4cdEsWQ0YPCLHPO4F3PdQGf8OU9DAQX2+FvTgu4GjcU0MPv9Z299e2aUURuDOF
NQcjw5Xdi3jF6IxduJPzF0V0p1/y4++NyYpsBtTdOBLknWBnB/0gtLRg9Lb1LZdR
lN5OedRoRtiBzWrE1CCaeu8vnxiQThOa5mYJ0Giyo1sl/QQ7+m/imVDg71YFfZTF
JYmZwiPEoF58cNF7t52VmHP36lw+p3RiRwi/vn0pzMZ1Arc/BnhWuU5iD+dlDGZ1
gjte8ZxecaD1k2jaLvHJ2y9QapD84JIEQ3P7Rw7bhPrqBl/x5krMnHBnMObcUuHf
O5N8dUoeE5dD6a5iCGfDCDfDfRKbTGgsIl/VQ0q+X5bYLEwr5gctTfZUqqDsV+NA
wFIFcwb6x397ttq26kCHsrUubrxFh3fP5I4KDXsa3XWFRMB9cMFQ0NRju15RlBhf
RkkRiFzcsJWxiGh4gayCuBJfofFIs3J2+jCnbMVLs6KzyulGAghqgtvRm/G1E/wC
rkO5kRNKVNBEQpJgXsa3kOjfkj+2F0Mp1kcWp0yn+XpSlTjA/W3frLW6AhEgSc1K
3kIwwxiWDB5eYeXZEomCbTXYvIbiNKB3kfielXNL7SE06s18oMFVm4XRZuXwqh4t
wSPIszHf8eTOFgvFQ3cueJ2TLgyygDZwculpyikRSPgjBK+XaTBPAje7mw9ILvLA
SoVoCXj31GKxRvsk2q8Mc3cIJiWq83NT0YKLv1Kv9M4nhuHzkqU3pcygUwsdz/xL
GIXgwTQamuiwYK5jq6rmB52fejPyV3IQzXoLon4WPcVKtcfe+N+BHZ6gQxJBx7lP
YKHK3WBUHCPZX9KXmrtZyalGcW0b3aMnUz1iWo4vEB+ExZ/YS+0Ysrff56C/WuG4
rCwIlzJnhD6GDNU/RcE/0jdMsdCQBVIzgvj/xPM3d/hi5m+o/UiUFUpWHG4mme+e
srpzt8QMW1wXcUTLZyx5zihHEfPk4+hCVqGMLp4JuUKCLR2536vkCKyWbKRpboiS
okK7lt1T+MnxaHSQx2+IIVcfNooF1xny/Cm3UQT6hYWFHwvIh7BO4WeikRFT8swx
+N2nMmbEW4nJ15y9dT0dvrVopUFPkoKTS2SRl2aqg53UbUJgzMp2CLP6XzqiM4Ck
wB0ba1fflt7kA1fK+OQP4VxW/PM4V5pRmlbMrci/A3ZDvYA274drkKe89OE57nrn
YT5JLIY+TtXGFrxiXeb2fuNfF/3ZUcL282vF3iJ+Q2o9tvR+m9nSoRIFHfFQJwXt
V6gvYHcy6ta/RVrv9KQLpeJ3SUKdzLYHQRDS91ZuTWEnhC/NrADGlf77c/deRYpt
PPqVPt+6dJWe+e/QtH8rqWv54dnRexvXTe/rluxpAYuQ2q/j2gr3aeFPTlw/KMEZ
Y9LHHXwO6R3JEK4/nBj4FC2G0ynz9OBJjA4YZ6bFAVVigdj+SKnMMINVAImLsPpt
oGXIsMznYCW6XW4Y1OXnnT1f1chy8IUhkGv37MGwBoY2fzNcHJy+vw2130NI7eZY
NiqpqDcVjHgRsRX3/AChnhh5MV/k6/nB6PXQZhrIh45WrBQQ/0rd7fDBqs88ozKX
mWB1diJR8TYAeUt8vf6qej6YFAwrQdtPjRzqI0No+I3fBAg3UQyN2Y0jFJX3VTVH
zW9fhrxXku93+SsAWOMVtN+i4FA99qJd0uNwio+M1O3in+lLSGPXyWRtHfFacqFF
XFPXFtW9cNdIORNlGfJKJGnk/2Npqirzo5/uHVrhtyP5WoJtDb56W9+TxSr/zNTB
zUAjbFSaTKPSepI8Z5mip0Nfk5uJ5AwPyuO0G4p2CvLsIy4S/6CRpXi3bVOqbe6H
Y5PvPVfmqq1dUhiIppEu7CDl0OA4hVbuQUU1LB/sBTGDnTyvghvEVFkuFFuEp+j7
0/vWqv0V3GprbEoaF2VzxVpSlljuoKNpl0/VUsXPKstfDtnNLPqACgMdCeOpbWF0
0u24PMkYBvdGO/2DCVJkcvf0JPBmuW6rF+EYv/4w0q8npyuUz/P7CZ51++BN4Ohn
1mTToP+qjWGGlA29R4DnP4ycXOzMlHI9IWmn+yFnSyrvH6ZaFHCcHmWIGHi8FkZA
58lFPfAuoBt3EV2U9MCfg3ULEqHpVurt05g+QXAKsQ48R4Bc65TLYuD1AOAgYxOb
luyAr2BZpXEu7CFt/2XpyRfnWtoMT366AyrtnP1e4KBwpHIIwpOH1DpanGFz7gea
LZSlCdeLTFzpfVZTlX/9fy6Y8doeMX1cDlDbZ3NWSBqLRLgv3Sl9qx3OlVkBYLgN
/i9gHefJIvQNA5UilCdfXeMb4jYd1BlQzXWM1ufHatr0cWglv+X7G7booWcgdp0U
wtTtqY1eJTqQoUCiVrlkm19w2WdfwYVYJHN1nQGdBCJ1Q59dKgFGuMU2zUj9TP/5
YjpayQDvmQWB5ezIJ0OFnZItddFdZ9tpAv6prWSc6oURMcOdMvKsTDBkLbVzWuas
tQPgF2OfRKynOZsGjzhOnsid7m7fA3+2cD7g5Xqv+vFxQ1j19eYbQErNr04Ezak5
2tGN8AgMmF7FaMd5h36+JJRh3TkDbcnIeH5AHYW/evswSdxGzWDqHQqVrFXphn9l
UVzxYZY6P43JEA/8GnopbtuuCV2p7so71x2/8u2lEq6abugUY8uA57jG4H7TVyXV
yKunCxOxjN+YxxASPmFcMdRLLbKpx1T+mQSi6sWsHaJevsKmdXaQXbN3brm1Xb1p
15M/1hNFCBTI46EQQG+hho0Gf0UoUURqw2Q1L2l14qIJiw0yvV2A4p5uxmS6I1g8
Vht59X7RXO+zq+pWykKntpdpBhW9QpHjyravcUQTbx/iGjLJZjD6pOatJv2fnvkO
zfSluT/kIXSAuMpHeh995kKFST2s8fmB8VTMEAununfosut9EFmdvwy96D6vnnqp
cGWDDYZBQ1V6N0jHAkqFecVlCU0dYc2eDVSiWNnIFCZTYSljBWLkdKG2JePmSTmH
M73V8Jp/0zFWvl1VcJ7wqjXwVVNrpdLwoSEfkAYRgBvuPsHgr1bx8m5hKxr/fUSV
Igx8WZkbQ4MUJ036uBRGBATScoMn7L4sGIJsW0ANMb7j9T9krMy1IkGTiUUSilO7
Ae+5HYpqxGvB2GFbs4aifpftf+AwjoqOBbE7K3v0Bkt6x2v2Nz9IAhnqvAWMy5FH
ZfQashdkUkGWeGzq1jRoWUmmBwmeYQX1KBVM4dZmsVtP+iyypXIjhs6ynNwQZL4/
bugL3cTRZnePp3shMIOBYpt4lo6PmvY7T+iRWVPl7Pg4kZOonh27v6W755Rpsap7
tdhX/UxSgxgDqh9uLVf0+qn3DbMGnZ4hxKyHeTP/ePn0ntwIcfYg9FL8fRufhPYf
IUAl6Monew+YlIYb8SRBMZuJxaYe/pFB/FHoHJY7YaL7k9qxEu+k+9vFuwh5Dk64
P43X67BdQHher45CXibWVjrbeqKvPWVpqggCthw9ZS9yyB1Mc8VY9ccNhL5o1DZU
U105LzbtqyqH9QpZ5K1SR780rhgIdF+H92cqTZgpHQ0fuYC2kAZZDcT8fOgQyKfY
QWLeCD7dY9vYk5koJuUhSH4yqZRwZEcDdq686p9FJayBdBw0qZaWGN75/yd+ky8i
/U9uUwJ3WiOTIHVof08zzemGIIHrLiGUV40orXr4cbxkCpMx0MkA/BwYA4E6Tv4r
OWeGEbqiJ98aJ4hW4Od9929bkydp1FWOa6QYZewhsslziRlRJCfB+kXzMh21yRQP
DA+Sx3EKJxuLm60FHHCLtuXIZbiEXAHfAqe1qG9jiCAWruGcdmIxv82zanL+JM6Q
z83aKrrJy9dfHzA0/2dJbwWgQHKCFZ9gJKyQ1r/lgQ0XpxULGs+rf276j+rfsZ6A
4dbAErLspC02wzxxaK/Q3jLiTnQgyxOCE7QDye6V5a3kkxYT6kDCwkYzATebfXME
miFHfSKin/EpmNe8O7ls+bY6ZGlNLA4LbIj3HvKWWJS9nisPjBqbEDwuvD9zgH5Z
48rdoUmm3f8wkEdgJxWwS3YJfYqrXY2pnsXqYIn5VaEd/8A/CUGlhP2Q1+TzQa0g
OshP1yWpWtqh7uCUOId4NNwzPY7qQycOMv5FoB9/159hNrgPvtgvv29QvTSVQ8N1
WJC1z9zKJ2KlhYDVaH5dPPKlqyus6xHKdVqAnslHHz9xosq0+X4B7B11jVr1+l6W
kH5tFSm1kh23B6Lh6XpJ4eiGRplzTST7oZJ4JKejqpE9g52ezwztRYixpRTMJjZ6
LE5wFg1Z9z+QFOCYw/8NCQGYiorZtmPZHEnC8xqs2fqcG+7JZY8tUnP3RzS/vIWo
nw27B5IZCaiYlqBfkUAjwJtm8UpqZjK674RGH9PkjY5jC1kXJzwYONiedTbFVeyA
CvvD5HA1NUbWO5Iga2GT7AhFwMU/KpNtlEqDnX4ujU3EDh1DSf6GGPvAr/zXb+rD
y/iWjk5+DTg0JDpSJkq25t+jz3A+FcZRLCtvHMIDjJwAiH0V/nCbh2qUEjmDS2AW
t1aiw5OKWSgvLwHavGvCFJn2MdhKSYuhL/MEWYNW+hfkni5i0Fn0qur3cHMvHKbJ
wjCIa3vM3CP06jaXn0CybYc5q+VrWJePbBvkQloaYAPt9iDY/fFh4UnLe+LICXmb
M3hCXaMPM3neAbj49gaLygIqqtjea1MMaBgDFZFzxeUVE59UsBWxGj13NoGbt2xp
pdSL6vCCHVlIHK2KGA+Tc5GapcxMNp1wabaIEqIyLLGh+e6aZ6pR/X5JGWSOaxwO
Swi694Y3aT1OjaHnAf0eeuAI5rljiqPCsY8apWbhMYIuJNBDqKjTNWRI9IjhUHQh
cPNHpOxzF5gv4JM+rrq8tx25W7zNGfVIQJb9jJyQ2VhvanMUjVd1Rj8xQSr7tdX0
xWqpXloBKCxraxQu8DayFN4J/o+OCGgyd445v2xfbcXVfVNXTeQT1rP1d5PCiS7Y
1Hby7lX6mCCBYCnorSyFawMBwnQST93h9EhxUlfc290YqnozN7GgEnRBU76K0gm7
fhk/pfEYEnXdihRY60wRQq9a7rKtNN/jS/+XP7XPJgWHxQfVBr02XoX+PC31Jd0I
LVfFGx0zR42brQfnaazTU2lVnsj/DPcgdvqNZ/+QqmD3foIJB41es0z4ud5Dc2IT
NoROALu04q23cxNhopWLs4JPsZlpQg7RBGwz6uB6i7OmS3ElDHz2+aBZD3znACTX
R6qPdc6mpu/n37VlxQIEBytdj2L+OeEbcrDd8wvosne1g3IvzJbH3GCSSeeONyyo
MysabrZUB969389lgf9YlTbBAosE6x1qkBAWafHrUFgGJk7SfBy9pYZXa/apJpy9
2JUTegPsPFEINs3Ea+5rXx8yThmFGkEJHDjQ9VYA9oK/NZdScbbR+WCbqg4jMREc
lPJFL/HKbEFA6qMgXrWIBGgl92vxo3T+n6vC/6yLm4NskqzYaKhG/Uqv9oaPqXxD
ZLt7ZA/NJ0J+Cjf/XuWWn0ypjcIKyhBAX4CuE8CXB0XLMATJgYvCFQmuZddIc7On
IFp3gCVygsugCcftZBN9MqtVzroK+1LXkWVKLvogxBOhXQHg+tUZtDveLRt7YMrJ
72sTjtPoNC8He6TJDe8ZE7/jzjzCIgmqXzL9tFqirDes3VkTS+SCzswlOy1xj/dO
7cBhg+fBLFnCKYvoDwym+Q3+nzloLTExCnWZBSXac6wGaLGOW6nk5U3SMz5Vr/MQ
CrvVRMZC14MhzW1TkSabJk5KoEfNZM4DDKz1PmikyVdAwvEzDF42QJiWNKdo4WAs
XQXEqdSS/bKH+hQBa/N1qIo5dbCpT7reN4Tt/j5uEa3hcyTk/2ab2/JuryFzUk6G
wX1FtzXwUybGl3GUWOUVIVqmgNr+o8t9RD2dL9B8S1rNtJCU6Y1NFvPH4KqXteOa
MnrvGNP59V2xxpp4rky3X444o7eFg8nPH+Jqvelz7oRcLysZckMsFB1tQ0Op8V5w
6U+Psy1N42dA9j3/0oFP6Q6n0Ia3hdQwAOQzmZk+N6EceiM93Vhylaqu23Skw5wz
tU1+g1CeNNmQALKiggbGpGAOqrUZLcptsMk0cyb3dh0lyadYE1KIGL8sF6l96dX7
ax1AnXjEa/Rca9F6+i5ASBH6mZVr7KXp6qjpYb8/wccegfeO1GXDHnVdcdktbx/u
Xrt1IMlUhbivwlFjJtkUpMoeq1q4s4OsuLxTiSVG2vrOczTxtZ+CFqrwFSKLXhuX
6aOCaFtXoOcXTrOQqMuw0VU36fdJ9bcndAnpVM7UDydT76bD499mdcnnlSPz8EnR
YPrqmhu0oQxaodTIxHo7Shk3U73Dhdvhu41Rl4SHRwUVDhQrzWvng8f15812vvvN
cqWNeJqVFl0PBycmgmS82r1WCp+QhWoEeWp1/C15uLpnYaylvijDUVOX7CWRoQkq
OAGZ/okY/rp0El+3mV4NlWYPpQ9f2lYffaTOAqAfr12BCNAqyQtI1nN1vsS0VJMX
nvNBkazl0WD8VVe/LmfuNWUvsYKoRIkrj1tICA1qnxiX9BFF7eJd3u4xqA0K83CC
7dV9Z9p65wBqpdddaswjWYbfHjc7aYFEF8FQTjKROXlRFC0vu/1csXGhqJcZwuAa
KP+IGwuYYNqlE2dDhyRt5Gwg3NnXmSlwRD/CrozYqFweW9IIlAFO5FaP9OUN5cmD
tn7JqEQZVbK5BFBagABEwdUjx8KO/TnTHNK8STNGYd5A2DK5k6eWX4jz56wkrq4J
WhCrT/FbyFlZXW3d5W7q6Pf2xjrWH7gbtidvoz2+zf/P8gNNh7C7akD2PZGdLQau
6WKuzrnsZTmDwiCrxNGbwiYhi6xQyOy43rfVMVoMkNk65gP/5sHIKiZYsH5kpa3r
M3zYhnr38z8jdC6hKT49oLXI1Zpp4ds+7+SzEiZShPwhqx4I4Q3fzDEaEfj5N7Rh
Na5vOFJ13MFBy2R4nzjUCb0ZtJ09nJzcu8eZ4OpAtPl4b6g/i7Gf6x7QCU2Ai3zY
RBWVckcLpNa6PvOkAguWYa8RqbU7TUuPR6fSEu+OWGBiT1KfRV/IxtO5cry90HNb
xLwOEwDaW4eMdSAQt9YotjCky3cPS2bKbBDjzpwckugjsihqv0qZ5dmzXbQe8/PU
0TYtJ9hbo6OF1MtdEcVhEu8a7wGYm9z9KJoFvaPEvmcZCTrJqjwmIFVy3ge7Qte/
Sgy6VZy8ABiBbZ0lxT10yOHZfozC6Ok4SzIvyHjOEQGmbCEt5aSwT00jg5Ly6enI
lYqcQWDKW8ZlUx7Ljq+xhCNuFvG7fuauv7azlKApEp72pkt/M/PmXxnxmeKqWb/4
uSzYSQ+DB6rZAIAJb3rkJVLwLxgKaWQYeeMsRGLpnh4Wj5cOH8VQH3AZBQwneH7l
0RxoAM4kRnXTw4zyedxAZ765S7TBqAVYrSFEKcOxyjMNt3X4KtQO9GFZJU03PMnO
a/BYa9PLw8OA9a8oTV785LyxbYi1K+yQAm4VfOCSSIQ41DAef6PKLohC/i4Kj3Yu
7Z2AAYfU8V0kIr/8Waurc9khnoRq3oGlSa63JCCfLmDgb1rwC3pMBYnSnzEc/A/y
ymrHyZr29C4VgtWIUy7wASRaX6cQqILFG08rA+uRzgh51PKMIN2xwM+Bb6QzttQS
qA71f1gCpbiFIxzmsBj9fo+KpEcXsiGeWvYJ0zvBD9MQtBuvT1jEAW/NZzLfB43B
xLTsmxyzcTP+78GOZKBEPOZp1McnZ/mdGrWdLSKCBz1R7q6hzW6GeWYczEfMQE/B
6iA0wzDOr7HEdWRkOJPOWCl8vOzZs5K0BXA40JlB4JdgcNUc2egq7IBoXTe0LxSF
klkpgtrfznfqyyhZ4SNZmcNeds6OvdeGRXDDWLlWHSnsXRsY9UuDvKrCvAjLM/i9
RG+7GnvlnP5gJjeid8eDEFVhGb+BG1OA6pZ1cGasvMKoyfWe305zzISzJK8T1R85
YlK6jd98u5RCaBT/aedumBcmgKWmYpDD/1fF02Wlx/6/uCGMHBFVK5KEcxLeSGQo
Cv6T8f9vutiE7NVCviWag4r6R7FJ1cKK0hXDv5UY0Aiyava0QhLn/7arA+zQCrpc
Tje7eYXXBVkXRFH9tFdhiytf58/rqxioIPpY9xK14vRafQNb2QSgWWCKcXhOZCOJ
y371eTab7jCOFCQ/Y+2S5na/rrJJeQix51UQTc4hXP1BXq0+d7RkX1LdRuH0kayy
R8Nw9gekaFbX/ZXz9A66Z5tfVVS+PLCw1vGyB2iK8Ot7wOjYGqunGZUaSOR/MEKs
jYQB2IncArSP/uSUQ3FuKFfd5mUu3GV8Scn8mNcxuA1qqoQmYeVUbnwqjwO18QQF
FjfsC920omYalX6UC14piYgU0TFRq75wQRklecR4kmeiAPoa1Z8UWtlqUcPCXMb6
RNV4NwG0AUIJ1iRaNvIJLmasDpfBmzbT6F2FNyqSAMdWoA0xs8fCAkE0EcWlq/jC
p0oj55zdJVbqCiBnBO724Hn88wGnvc558drD1fNXylZjoucoAFcJUfWEGcLX2/83
433OWDV6SeLRlm2KTL9DkNM4vsP0eCbC5zrZd8k8hcHpiu1ZpAYIGOCBYsOwXbdx
mIRsem94xTKJPstJmoRUGDDdMvwiobS/1l5WqoaHPyKzqpuIVgbADqvHS3IZNMVo
C27FdU2kFChtBEF3k6kqpnsCK3Z39nrsJ4MfNL3pEn0s03DMPyuRJHMvxlafg/Nh
UcWdys2amiX/KGT5W3x9EQL0TKbUski7CWin6ukoEQ1EaJ8hQKPjGNuxAD0S/eWA
CCVDbLx5QWi06+ZZWML8GCPwQUiTbi8+VNuAon3lKoRcoONC/6OwGKqDeUkj9XZj
sXlZP6kExFPmJOpdNmEIpvBL8jtMJpf7I4ia3iBgSpuAPGyKg6u43eCuVynCamTD
qo4PctEZNEzzJm0GV42MOUDeJpYI3N+oZ1qIexbDKbZjM1r8+I+aogDXAxQsm1RS
C0KBu1qveKjzOtIRDKwRVZOwCnwGpZt7u94MXP12yA6RobpzeOgxHkyWJIadwy2p
lfbDd6oKeH+q2RmH9WDlgmGcIi61U8fqbKP9VXUhebtZ/q2okAdYmFQsfnFqVUUr
xb3fl5zz6Bqyiw5TizhaL6cPRYwRJWtcgRYCFPzD2cQEZASnGz+Yk4y1fscwE6sX
SOxPn1yQjoR4W0uSkW6h9ItW4feT/IG0dxyAt/8lcjxkyid02rPWAPQDkPo5uyJd
g75iiE72l6vbCKQWOnUEtuX/qZi8prXWHm2U896HgDtYM9qPPTH1eXkVZbA18wqq
+oM2MyZVKYtnPFUbInGTc9XAFWxCK6NhOAXjt4xeOHN2NRaH44thtf2LKtidHYMM
DtQQcCHa5XmnxGbPTnNeSHaNnqvU/uHenI0CmvC0r7lzkP9uPc6NoUtDzJs/TMHO
3rAtztrGTuzqdDfPocvzQjimqeAW7OriN0fj9wwKpo1UeqEnk5I+jCSVsjtLmUL7
ZvKlmroXn4C/vTtD6ydGicB1Z0D4vXJ02OA9fHCvjnlPGrMdxAG8pDtN5+BdEL5R
TuBdL1MU16hFvz3fHcIVgj5ICcvQlkx8CvM3Gibs5H0bS9CIhgHcY1KsNfiPucrl
UIpjAHO3qjixUo+ybbCTZxgywKZ5JQHdZPNxZEXKF/TkzXc0XdMwdONzVYwwP9qV
ZgG5TJeoMApjFyMuy0uXFK31bc0FqYRMyhroMVJmYPb1wcEdXUadM8xIZpTSdFeF
vP4HkQPb47+rD9PUtWryUXltBvPdHLq3qKy6D+tETA9n7uxf3lTfMpfWFoDPQdvi
ysCZbJGRI7yrUqjtKPcnw47dySa9l0N8dQrRzjUCouDOz4UthIKKyGMAiaMTKZDe
0ebmEDgHJxhVs+8MPNAWAdO/viHs1xnsQwDLjnP8F3jpf6YmlAJ8FfKzSZAa1uqM
lmJVKVjqNRoNF26vS+sxlVd87KqInwuvu+4r7kjttKPf1uRnjsgrcUOaEdXjDA1s
m8YOKS2ZCmtMUVdz0fPtcVARipDiucx64oUJaW2C29gAiO8EwxXOCRx60u8Y0fCO
sCRdPmciPErB/zjymBh7dKrLXly/BC0YN7AdIIFrjd0NcNOsj1BCRLr6S1+Cx11q
+Az2banRW61u0rsqjJrnfdUdOF4y1TbYoYjf5tuZ4hcDk+WEtbD30pPLgmn5nPJo
ZiJO2AJeNKrJukc8SYt7Prms5VD6rLL9MYDon7Faf4WPkUXP5MdOlSrMhgqo94mQ
TVV32KMEXZ7U1EyizRxP2lSssSWT/7tRTmVOjpHB37mKV5IVZRdUv7MzigGgDG2r
oVRfjgPqV4hCTMvn1OL1Jm0drnPDQhrHNB3Z2Qpld2/A48uxuOyOHZjfh20WyrVK
ki6ZMG44PAyPBjJ0Esk4WyjHnSOtPc1c1f3Mm7T7eeENlNSVboreE/20C7SNuG2G
JlamhkJNBo7SzZ+6WDDop37206Z0ZnzmY+jI8szHoOhpKTCIf0p2ePt7dvID8dD7
qamm2rdAx4L7BvlFUZCyXjgaXuKPQp4sdBxOpxfxIeippxwe1t8+/jdYpY4YI508
SfAer7HMc4XgzE4gS05UnTpuxF9v3Jr/iKWYGI58+V4bqEtH1HI9o7M0ZpY2rKBG
URPZXE7xtJspYcvFM6Z7Ye033OwrFrlGdJljEam4ZlOGtNfG1k8j8Kjs0Yl8A0GL
+gNHwazPKYF45XPIOzgptPrh70af2KGVunpvHHfhYEqBVWu8sASYE/QGxDobYp2i
5b4kvPcKDfPuFclzOHeEjoTvd8dW+nWG/ImWr2xr5SgRPF4iR0XAb/rfxMH8TBt/
qTQqNpv50/yhbXuEWVJktOhIIBxnfDcj6GxxZTe3/MVeLdB1mMNMWcuSfed62l98
ezdFJVPEIcuQtn75IEaLFNbM2KwmAL/bvhqMMyWxQw6NwPZkWFla4uvVsrUrcDU/
DoiGs9oVdMr32vRIRH2Lk5J9Agbjh4OM896+LU0NcfyufBz7iDvJHfoat8CUYW3N
xOyfTp1pZ5oO4XShYgLM/MnsZWEkAN8IpLhfOvA2ERNwg72ydYjJBZ+eNoECoLLW
i9OkPX/1VYCCevPU9bjCfLmrSXB8YbfDMJc3E6J1D6m5tC6ZFDgKD3uRulOprbOc
upiwFAISaXYOLiabbQLmkMqk1pExGC5pJZTF4i8J6wsJ0RUscTkeD6sTMnC9nesS
wqu6jLxlFF+IVifKO8cLmftjg6PuPsXPVg9FxYcb90DdQzA/M26LBrFMgNHz3Imt
OlZhLr77lxLXlMI7jvGxOfcgzp69blt4ofKo6aqYhjeyC5Lt60/07MrDf79AzSmS
b8q/7p48NHF/eP0yqdQtckpgdVvKAdeikpbxVLQifV/wPSdcTQXF0unCgtNfsSfF
LMidklKT+ldkNphZckmwXP8wsMCGsIsbwES1AOQMtlLgfZlc8d9zdba/d/OfdHuR
rToNaHcOe1/iIIWKW6cCgUv4Xn+qmCNHjb35P1KRCQxyeMqHcfVDUTPMlVm8jLOY
QJV1T3Y/UYeBXEoVCd45QyC0lcsEpgerJLP2a/DX6/mMTDyqjrnQWKFmjKZlPgLv
foO0LQPuYapqze7jMFFeAgtt0xNgo20CRBMYEHl3zYCGl3gsaQ1Uirg+E56TTm/3
pBKHvbj7zRQWnGJ5JR353rTHh94XC+bzaof5DvU3MbIDJAiz/PfWLsRUlYWCv2dI
kFf89CaQt/nfgCatuYfppqm6EN7/tfR8Uwwj0mlR9QNzqpzlA+P9AqCcxZZwFx9c
qsJ6yUCrK9YOlHDdydl8wzq+59qJn9HkFSb7dx+tuxrVhfckPfoojuH/k89b3GqZ
kTdQOqiYLqHslsMWBd6nwk9L48QxFk/mlE57HAeriUvW/+QnDjIHeqylzFQShyTl
h4/xcZQRI+UxL/Cm4fOfxWPd5zff7ukvYlNOzxav5r6T2vkwBuoh4XSp+xyPlw+A
LyZGNL3TVXOo9XuYiZ8JCU7MFnhxh6QE8GVz3vn61uLEWuEUW2/35LTYSCeDvXps
V5HAXXpDPNsDT2VoI9L0Tx2VTuWi7hFHe6rfKMhYIaBgXg8d9ERaR9Vxoy/2t28W
tAmc4YnuU91VLNQFdrTMCwe3lluVuyZgdqnqFG5OsCM3XTCdIb/PAYt9kxsyaKVg
zH36rnxHgmyn3EEy/I9zDdQ/7Nohzc7P5+XdUbyop7Z51V67DxcuInTsmL0YfgXv
XN1O1SNqtAtuqL7au76QXsbccQhPbo8qhGLnYxLVx34PPEJ2qLaPsgvL0cPC7Hvg
iiBNA3nACSakJ58JfKOUm3p0ogvmwDbTudks0SQJnVx6GSZ8liOIaPkN7YxBsUEx
qzwpKFqXjBh/Pq5FMhBPBwPSFQTvfDRHImwFzDaEodxNhMpplULYTwW305Rd3aYZ
NkX75mdf1p1uYvW1/ZFB8dyWGLiG3Rw5dSm5/zJK6m2VgvISx+zWIa/SbxAMWUJD
qb0PWqWHDm7v/pge3vZ9IXQpJMr1FypkGaGnDDmTqIMXJViF65ANjSpcNgjbM2XI
kPbKpHBMsJsMtGJRxgT62Q82x4aCibB8dMus7lFmqB9AbJjuxEbhEKoeeGPyZQjt
JLGJNO820QTmPjdgiLlt1bnf+4zdXImS6tp1d5RpKCbR2xgxqNlykuKvTr6/pWTw
q2aRA6OD0Gn5zy1ZpcEc2S7ErWmft47RZJZHDzoFE+O1lxJ2Vpg9DbFJn/IgKFGJ
NARQxVZPh6TQO7chH25CjCBaVUNY/GGXs06pDEk9Bdpxg/fi6i6JxiEyAMKy3IHl
JXy8P0G00mc6BSJQ9OGCzYOD8v3/YRp6PXX4ktz2P4GA+LV2DXjz4bRQgS8ETFGq
vlIJbjY5997TGKMSwgIlkkV+Dgq0ZIt8C7J4C07XpuY6IBn4XWqq850m36F+dkjU
b4ydUG2K+VKUMZMz4VY3oRFaQyc9+6iYIhLDaNYVg+pgXRagkL4uZdDfvmtVg07L
qKYFywShwV1yLN/C7uterF2pjEJsxT29dm9n3LjSIwcKllo6PUq1YWOqPwWBG5Gi
nt2ShnfOhjZPdkb4+kVvgp3h5kvFwGbExcy+/RwP35yGdHrI75t37F8kIAh8LJkE
IOl3H0Fn4cf/TPIkrazBA70i4MSOsgKsSxyu1eRIeAXtLLUHpf3o9YW406mgHMsc
0EAf4Mmou3lpaortiDxHWgO4N4qy0QHN8PeUVNlh+QCIFhh4DTJz1NJNIqNy+z2o
7yXeLWHzwxMK3qm+jFqnIAPfXNYmRx2oGoSFis9FIC5LhvaMA0yoICQhPDY01c6X
XrHlN+33tZ7W1hE9t31z4bLQ4cFVFGk0/tDyPfMfUJy/gWxcXha6emcfVG+T0ML7
Wla4QUBoq4zIdUcZe3giJunRmpIXv7Vbo884HvVtCPlj4IDI3+7sjvTGrYVGByNv
9PKEE8u3fBdV5e7Xv9JcR7HoSGiQaM/lT3TWfytTOrENd9mLyh7fsQcW2rNBj3vu
hSEM1Ds7uueK58R30Z40SrqJHJHzv930rLfYCBApMvjCbmCWBfjKdrHjzFqxYaG4
Y0oH14Wo2Aut75tZLei9H/23wjTTeJUoEBm8yY2hOYkBjLim9AgT3VOrczOn1yio
8QcEqxl9clMJHAMcKH1fUXXt4JVMbVZd1qFXe61ArXLGmDG4RpQRrSPqdns04fZE
6I+Ri1k6N3KTi5YqxGpPykSIVia9putM6eFd4owXy7H4jpzyXuMJGY0QkCeUNUq9
ThysYb2mQyRg8d7zGtQGD9T+hNagrN8ZZgIw4LJ206/jYy/8umlAtos3xqlAk8xY
KD+dtl96epMzUzUN3ZbPkejuPBHL6NM/apMJ8MW+3KWc0swLXPuEVOSex6EH12fJ
5szQPTAzRJMcwdMUCXadojSV61dx0txP4ehuAo1cBq++QYWb5nm/eIFuO9O07JD/
82vuz7xy6O8E758YoqywygWWLjSskN5SwSNd43DRiZ38eGW9oUqUP9a1tS0vWiQN
CnL7e+G2eHKpQP2v1+vwLH44dMfBdPUsngLP9NMkNWQQf6vbGkIYmonbwB7BnKd7
8wQ3Bt9wyku6zXhgYy3dD888cB+ivcEFo4C9FeS5aE7dx3/+7VqjBC1dnsnokAex
0cHyRjQgR9QHaZEMtKLbTypCPQw2BKtQU+9n4eHfFI4TtoFR/y8TeMqxq4h5uDeu
ZfAThgUNkvxCQs6P8r8vYJXrbpOqS6ES6NqVGeitnItVzOEOBqcnqtB1yLEEk/cl
bHK5M42sLd4HLl8roUfLybSft48nqa94QbNj5jX9ScTH5RYZPyHUp2zdWIbzc30t
JNukbE5NI3UB4cuGEQqvcsMCkggfTK2h4B7UO17a4SbUZwUKE6S0hkGa7SabEco8
AiWCDL6JSRJfzgWlCq9KckvpJ9wZdEo2zhplqfaGbGamDRVkpPPG/v5tq35anCbM
rGzxrA0DUgf2J7ZseRCBEyX5gSBilr7sA+cAzRd6aHFbot1PH3FnNyrHiAbTS6xl
8tU7PooTZNOPxGe/5g7Ev7hctx8caS+0d6XhXu29/7QxtVMJLyoNhA194H1lZn3a
lo61AbW4059rNpmMLL81wjwVDccnRS+RaXzzi7wto8qNNgQLKWCh1XnvABLuAPJc
nCxthl9HkpAy4CtcDpidTVRxoRmFS1u5oAS3H8JjK8PIYuEA0N0zP+nnEvATqnKx
puQPFlRTHOLGwktkLjd1quqRmuybOENS6Xz/9MmIMrC9wiib6l7PkhKVYtR9VzOC
YzUotcz2pNgSJwoP2VT7Vx5hUyRIUZRFXCYI18Q7UMWdqPshLVOllAkX9GAWqLeq
AjfYMRSUZw7YEM+MMmPnsuAgDYYtS50U9NxSJIaP18kNG9MPy5uhQox3FQApphjG
9XCTXZTDONaI7g6kTUWyIdDESAeYGqZ3Ss/PlaBMSMF6kpMjUivJIicbvYnJBVHE
RJN9oleq55/ZskEGf2YEcP/fwqZcTrYmQ6WBinCzqw0hT+U9RgBiD3/S4Zh/2A/d
tUfrK/tv77Vl7ks6UorWHfEBogLmoSQtaZYWR2qobmmted3phoFn/hNI8BCDxi3O
+R4dxWZEeRfeoZ9VNlr5R9GoAjEDy/q73a3gsejyGK7CRQk3phtmhVbg110cRk0n
BfuU56tEEyE0Ows9Bp1LoM/c7yt5eEU9oijJ3+5RY/krI1mBnQn3C1rtmljdDA64
4diJeQa5uHH1D0gHi59p27UG575d7WetPn3E7ThZ3sjAE+JnE22PkMClCFBWFqyB
gY6CxsFqXjhq/woWzEiQnOwl3TZBun7gv/yznkka/y+04oQox7vqYxbjEDWzTdQC
tNwvYhUAfTgTxfq0up1+s2dn85y0qCjZ1PMengnCtUS7nGDtcdhzXb4bnKAtmIXf
WjmjnCx7lMpmnzzmN5Ti1BOiZD6RZUy/yFxa+yt5DnpQa+HPUP0Jpm02RgieHjBX
a6K7lZ8vBSml2grekbS5PTijokgIcluoOiYgLyarF3PoZg+Y1r0HOG1JQ7CAxTFI
ohpVFPE9WoUtkMU636zkmWqZrnQw5+2/DaAuF8O51A7O9/DsuiY7I/vaQJWfvdXF
thPyDMnibGCc8yYlt+miQaCfdUd4kaYeJ0f0Xi5SLMDnlH6aT7vFEptgqihlFkdi
KqMM0cXSMMlQnxyH8SjVFKWQjD9NE8DBLIRxWFhIsO6EPAy+7zXc4EEgsUwIv1RX
YXA0aVSM82/GsAdGPd0aEIqPJF4pzlfrsO5CUM6c3kQBdSs/YcEZkiyTw8pmJLVA
8K/wnkmKBjZnpUIGFzT1Z8kYL3Jb3+B7Mqb9a6cpgOj/2kI0B7rb/5cZ65bYshL9
FPo9QsU4h1dcH+ciMSsvqcbuOiYwiPdbkkTWHd+iJg3YK7pBRfC9O/EHhwG8DAwk
XbcEvhqDieU6IkdK7TIotjIjdA5JfFXNA4a/edyaHD9MV0/UaNaplMpcOKhbt4PL
Mg8lBUSCtoOhVXL4tEyPqha+wRMk1yGUlMZvqb1oRdORXkERvh4icTeTNri8iUXy
Y3oiINCNHFzSnvGuQpG4s9MeQppUfVc49V0bkJqoKV8B5Ffk1UYbRV7tLjTCif5g
8BDJF/C2CgC2fn7GG+7LrF/wywY3YvaSFhrwP+O0+2s8NbstKLGeegeZ94CqeDJU
DJKL557c3J2P7J2Aj3LGjm8Fg0XL5YS+35d9M7xLyzxCN7Y2MFf2nXm4FlbbHEfD
QbJVufvOLOw04nr76pZ/oVadpTvJrnrxw3YYeXO5j4nzZeg0dDdAYdeojqy1xMBw
Ys+CP2F2Ng/Gl4u95ti3ZXxM5OB90BQKLExo5iJ1nObB+wK1SqMOV0EFl/3lMk2e
IzSwiIWF+OaXiNiGsCORaJ4VGqnjQb/14M9lgQ1niI1RsC2ZMKEDBAavSntEb1gA
YRzQbBiL/wKK0U1ArM/XeV5XvKSQe1tOHEA1FsOwOsAbOEwL9MujdFB0mOcGcTuz
rr+5IYS9ZA7ZkYC06VFCgO+2+B2ATLukcVrZYv8YF5gbKhXGRJsqsARPsDceCl2Z
rmDGxhnpL9DPDOeL58NRFUsBCRnJF5lZ7X3O8eol53Uz6DOveGUw/C1A+iW4HhOO
JWCqPiZujAEnCWYeuzQHJOYvqd4W+V2NqdkQVoDKIVG3i8eTTfu0xopYQVlM3732
VWJj382esroOvY601NGY1wDQ/tTvMyjVqecfJE1I9eghs1e7onK6/htRgb/HOJCv
FIFHSlecdvswmgCcY8d8mA8d/9SfdmqngqQuZywJ2zFlUijsx8/d6HRpddC25yMg
gtApa1W+muOLJxlnoiFQrSoHROvR26eYL1g1sMepZVrTq3I5aCfa8gBof7PpscIx
VRSDP5YcqzJgvdVQMV8OOF39vI8TmKqmLp8UkUL2pS66ZO4IbCxgXWTvNP3/lktx
hNsZxgtRYYOzCkZlhAH6JEl7vb8ezyh5LclC99uRTd2cjfqDeSCZFqOXSm7qNeg3
YKe7cp7tsK0fK1xjZPkI/ERYppLhc9zjY72Dz+DTRkmtZ35Y7ap+vETiDJYcInVR
gQzXikftYZq76Co7IDGIe6W1ILozY7qw8+x/1ETsHHx0vdXlag35tzXgAL/2tGB8
MSntCTmyXxZ2VUkI3do2mGqM/pdOP6yRq8YG10UmIRe0byUiqJOAbetB/RxmKHrV
LdBpGSHBwzX8e/GXOXSEneXcp9A3/LwBB2svXlIivp2mFTBkQkkSqAHFBNs2Q6bc
vBIA8KbtWChhmP60cxVPKm7iMDGujN3tTPuM58UmRmGNr2vX4+u9kS3+bKdEAFdW
A7JaIHX+/4DK+GOMzeicbjA6lB456gl4HrE3wlqSRiYwlRsKqjnCLNvr8CtVZlux
vqPaIs46bkszTuK/0bLXaFAW/Ea6Qf2z03EVXctxzCHJyd9TeiS2EUvsBLBcO3ka
T4SwmiOppBOOjMCgCviC1949uwrFrxkkhPoar+Wm8tEq7CBOyWChK0lFoePVpk4g
stwzT5pAmZYO7AEzukl55jvdzk5idWYRABfNY009PlcSMs0dXYs5DaSss3ewEu/R
ec9o5jBATh7x7jrvdFWQmmIby9AyB1p9JIVa7cXD70FCPONtDPN8qC0UBKTvovTt
rT9v2r2Sxu+VyUq0dC3ZpDVWG1nbojfzdQq9ukL1hCJiz3qI9pHjZGdr0sqQFX47
OBTzltlyY0l1+WByV9HkRgRIHT96QPgm8rwYZcH4jAwr0fy3QSOCNovZlusT32ms
nh4u/qtM28tsF8K5UzrlDvnaOqONNJYiNMoloQhny+UabuufncjurbQw76bNbScA
oggyvwitg/XO9Vg5HzqsmKa1QxiubZB84V0QMYLzqRuaFPbMPkgrcvVEBXcoZ0ph
H8hCYcT+iAD2KJe87sggwA+7dLu0y5yvmt64N1OHn9nR+KjRqzSG6eRSRNxtRgDT
N3qXZtSLPDOaNSWgoDFkYYNRye5KvAk25eUwjgKf/1dhiONA3rrZPJMjc6x2VWR6
yE9HUine1jsUTwMz1FFPLQgSnhxeXAJ+NIRfjPCOrdJ1P6cLs4HxKE6Dawz6mKoC
5ur6AYENr6k8b/Xod2L+3dPtmywKXr6ybFO4Py3mYpxYMpB7K2VyGPYLMO4vQVM8
mOwoAHjfFnm1FP065DDen+7IF1KXQ6+RUkcIZyxwcll3bP7qRihi/SB8lEyuP1oH
zjcyamUugK+fXgE/XlnioCIPpmVm5CgjZQwnKXdMdZtXf5+gWW9Ir1+r+7TGBZAe
ma8aqcpONiq9DVsnfpprT7VETeNYgxzEEtIU8yjN1Blo6lkROTMJCbyj3eLF3DCP
3qUTCbdE9d+tzGTE+ytBZxPEH4NmCRYMemjP09SslWxViI/8gsxFECwYlrA1n6xm
hvSFZL6KuKBdVtkMduMWGCtkNhqKjOEzn+ZqeuvZ7Vd3DhM+FmTzeubYWnTifP0s
NxN8UmhX1/rwZB23IfQu86wD48kXIN5THIbqfDeyeilTIUw/gQ2kHgOH6F+I9gkZ
gZDnl1vbhkOSFFi65gYeH/vxSbeGFqWb/0meWSY71InBEkKwNdtvmkdK8u8P/rNI
U65VVuUSadpynlCkdNQVaidZTsPhB2mjTFfg4I+yf1CRNZWU63I7n4Qid5cYdiWz
DeJ+YBv9ZRvl8K61S05S9A2egFE7598ZHbikCWYah+RaJSlIEW04F0y6Lbw7nm4Z
D4Ss6Gw0CgknE0Cv+Y/DXVWpivOMsODuZC2yd9favIgbKN5h1EnnfxeN6qJKfpVk
/wdBqxG/rkysgnQmLaqdhTFxY+rvMhoktissKuPcxCDLOV4qXpe6XU//HTtcsIAX
YubrczLrkXfLNIseqnfbmVCay208Qtp5O7gIS4Eey8YbtRZ3te40S7z+yP01hPS9
5A90IQQLTDYCDSRWKjbpiB9yFl6K4FFiBfealTW7xQLOqJYg7rO3CrquEL3sUS6q
6cKN9ZCWZwwmnPipn/mLHGw/y+16+Ym/F+9HfIAM32La9+pzu1xiA+lwmJyRlWU+
+zVXFj40rqGjRLPGHaMDiFNad5kHk4SIk9x/35DzqNRV2MEoVYtgHtSjAeA+l1pd
5U8v1wzE0+n3UXIdsLK0JgCIIhfDeZNoVdRShf0VhhhugfoCeqenorrUrl/inLTi
G37HSl1vuBp4FjoN3CKcvhsMM0aTJv5HXsx8eWCGzzUzx2gK23QELYAlEDhFHhER
rGm1YDpW3tSfeDaKMaZMAGzkuPOnnit9PXrTWI63dt1F1TB3Gk6Zf7hEFyNEDYsb
QeR9TXG7vDXKLSVJWCrXNUHqHCiQmjj9y+fxZQ/WT7ffznLRix4qFvRR0ddV6P1H
/NYYTq2nb4t3/NdP36iwrvIDevQWmMJHV2t5HyOmIx98/KosfclseYofGEkxpflY
MMXqVYTMxFP4XmQJ+Ju12Kjb5HS2X+UCjg20yhy2SNlFJgCgsX9uqW6vhRaf9S1D
u2X1U7J6mWyS+gWmhdMUNUf0gYxhHbemAo+Ucshbiiy9+pS5GWMASxBB2RHYzMK1
wVfId2jdeetiekYjHzGqKr5XN8uUHJ2h9YirF/+Fq45FEMSSuxo4cm7XBymFqVV7
Jtchk8jrk/ysuZ7ezPZ4T4lu2XsT3gxIOMX7AKbfd+TwJ7okBjAYCyBNPpBC44NU
WZr/Da0ErUB8W6D49bkQ0b2NS5DhgFJRhIFAstnBm03QE7DFJ4Fe5Mwn2t66+HEV
Vw/cj2R7PFq2n3ctELll7wQwhk8WydU8CjM8Ds+oENUu2+KeyVerpwCMLb5L6u+O
Cij5j2EQKEnY5rc2vyKy/UJpi7nI9A+8IeW0wvf3ffC1AM8/Efz5wteubGSotVs1
TBNjd0cs+3YjTHk0Nl8rWoWEbM+CY6LWLiwhvIbsxg4JRpjkSvL4ZTyb6FmdgZ5M
d8yyNLwLsyslmjsS8SRRpDQL+zZJxby914Q3epJAR/nIha0+Y2K/vz86QpmCBVqC
31oc/GpxXW25ri0YsC5cUlTnREb8LNoWDxSTxvkY6Z7velckPifgfu+BjuSF5Yfm
bhhqAiAw8v8iPwFjEK3o/Xa1DUPkI8em79xq7AzMp4tug2HheqvScD0NAcvboK2/
2eCkM04cwU9YkgHkLCgFgATbmdTZjS4ML6OoFjIRDFRdX/7SCWCu9IvwkPUvtzI4
DwwYkXB6mGr8WBKYYHetB4c9fuzv0Q1IBUC8AFlaqBRdVmaTZnTmGEXCj+nJSieC
yYCG91l/NyZEquGmGWDG+rNdx2X116rRPjH206X2T8w/ya+w/IKQU38El+Kfp8lx
IiuZDTamx1A8/QRhES3WJFyv6cEw+iJ4KYu2phNClWtJIv+SQAMLrnaejrgNnY7U
CszX7iaSJnEup6FLSpb7o+pzbbVvsRbJvnV+rBJ7GVsF2ZWUOMwxEb0r/+ebGFtL
mCDRsxNFXbFJVr8cGEOzp1uWZEBoKhD4cpvJVHiBPmkO/Aw2T29EGbLqDlUz095l
bjw6w2jGgKvgHLafcYcXhohkhy18Ueq08QdFbj2brM60p5nTG7Ebsmzk11GldqEv
UPaeYMSAs0b6cSBg0hC7GtjwztwXQs2HXqOGJk/9nH6184XpwhqBRuitFM+OdPeK
pthQPKOSyqvTjLHK6C4s4Fwg4GjGgsKcyaWwcMwMGKLDmncnQ4ZjouQXL7hueAng
74pA/0iQrFxOJrBMlSbO1lOlh8TbnyGlNbavI5BzPiN9JhwOZyLLizOqS0dUomD8
V5kZb1LKLMU5+VJlr+KQHqR5vCVfrvb8YbPw+rWKYtBTtvoKJsSHRE5y6XYSlpux
KVyZT4LUjYWCHpSEqx479x3qBfi5rvcJIq1ccVl8rgpXv2UOsAXanVll97F3DE8F
g0lw4KpgoIUKkD0jJeMo1w3a6lb89CzD7xM870EU9T1m29KcNB3hcbNDc1sfl6Gq
17G6QviWen6gqbC4oXGPsNmGxcRvz7dYi9DeYeEIWkGxYOeCUCU9if+b5yD20trm
SQc3LPZCrE4bEwCIaQX5RXd12CiCwdyNHXQwpdcTO1SzzWbFVCERTkiwkoSDknjh
B2aTRplXQt1SOdnyse7qwL8ZugEn9EmSoIh6bUXm1iHUHOufBBKXpSbgJxyibYCN
/DLg3kBdueAowKmSWE8H4dTLtRwWcjpE3sduklrdwtL5u/Z2OgS0NYZ06t+2EfMj
zZvaqs2gIIDwe6lwBa3o0DPAEqsig7SmyD+AB4iwn9bAkI20atEb+KJUDcJwftii
6sHhiRJGIK2K7vxBAGMTDUKdCcNTD2uZdSlPTiLD1RjkVP9eKgi3168fqJ3R6Cu6
0BxTn2qxPJ0cS/Ji/MUdbF8xqGWWPt/ycYmIWtK2i+qwbKsYm7+Gwcqdlj6tCaUH
yM4wM+n5hPvFpJKxHjojNAtd9YgsO7c+snUpGQfZZHS3BG4q5wfhLH2ZWj6HwQWz
IbApbMSMdxEp/6HbnyBFeaq4AcFpBpzUBKN+4EAG+zPnzVhgmuThU94weSeZlfgf
Agnzv9eRGREgwqSnsjkX0c7t+4TUlWhnMWJn9GMmkia3QJ63vnxvGT+xOqOuN1/1
jvQUSIy1Q/KkyKfvVb/U4pFq04scREMWMNtS51FlObyqVFclauYAHF+IggJpVP+7
U3pkIyaJz/AVr7s9iT0es3AiWR9bwNaUCfo3lQdfkbMGxeiSw9dznmXHHpwZamD0
IMt91snggohFIuv7huaj04KQPVANfOLNacn2pbUvT2LSpwgzdpaO7cU5wpEIblQX
LJm/461VabRfGTMy3a8F/eUbEDupJ2iBeIR0892UDsIom1s4mvThnORp3u1Sc0je
J7VHShcBPPRKttFW9lh7H9ZnSiTO0BfbLUFlGkF7UOYpE5YwuMtFSQPlA5tLKw/9
ywPbEzP2vj+Alr/UrIa0knVzyhoRzMllTyQbNaO8kzloTwwELPHwRgLXf6h1NgJI
NnSAVV+DN8pp+62krD5cwNRxqC6JuCpxiEoBxi28+4+J5dEurlZKvIKNsGKIdSE2
fRKuwAYblLVJV1Z0WN+l/e7kGtCYdKVcNkT4KioVZ5tauzpM9DvcpBjcK2vymY4r
xFfYCHk2kZlKCHKaTmR8PRekUMKBqlHseh+D2oaK1f61KbXXxfDqeLlPspb94ktS
NMpxiiAGYgMk5mDqinj69iSzWWb/SX5pbzBCYs3KqBM4fZkDXbj5wJm2A5GNzvQd
nTF6UlmjxlN5/ZLUosD6LaORofidc09+RaGmXBr8Z53Ehhh7NyzJHtR/lK0cEqUC
n+JqUcHPOMZ9OHCEUAKP8UZ78VxykGpurU5UUyDBBoPb/CzmbtBuLMoedTjpvfnB
qDDMOdr/KeDQI2Noi3jYApPXYv9kfdqWcreIxzmwtRuCVAt5oM/5Jkk+uSkmx8g8
0+B/jZ2QssYyOBdfZ5LRp/Drmq1DymFHVO8wr6YOXSnZmiFov8H7Er1otwmcHJaT
BTvjOcV2GT1IgELbwY4Wrl4wYmQZ1nEaQ4yLRb5JFRKays381yzNXt/DnbffoFUz
DWVPR7zFxTi++Jpb3PYJq94Bh9s5egJ+E7weya0gGlapu4Ci49942hj0ggLz/v7q
OfbEQprGGCEDsOsJEvClCYqAQacxFQDvPxHeh44ZDdCUI7kBhgHPXgNEXwCSa+WD
8f/XX52ZHIzyFsKKrkeqywM0hzti38Um/O2RpDnacnQ8sI+9/NVTrtUztpBEMFqy
uDDOv6X/uGghb4UDIYb9YbAheeD8fHY2/u6OVb/g5ciPhsPQHxA/3gDLGZ7z4B/X
RvNilxHhfKZes5WFKA/pNupFyd0UTo3fYssNyNgWWCapqeydjE2YhmcCzD6mk9gk
vpYD3dFOqlMaG05qsZsq0pDqD0w9O9CH2nSm2Fz8P00HThGOItBjaQqcjkcGksFf
L0Fd1cT3hJHWX25Zxr2kL/lMnKk7EO2Opy/uiM5wMDDpQKY/QGq8Sucd/0721LND
8aa/F1rHTrsK8V4V980Il4EI528K/RL3QUUGorlQbFsBv+bG2wrf9F/6PacOM8U6
4W7Os4aqeeCZwdgZGbOP9gztuwMqfnl/LltKcJgR6hTq32rF8OTR5jbtdfKPo9vT
QGJkm6Fb8uuvS1k78UzJ4P8ZEXaexta/hZUSy+lOvTCMklIBnPhcNC6B+crBelyi
y4InmuI7SlkNS0eSiqVk5VGEY/CcPVgQCGsYMUvwGT7jna8CAGxD4fDM/Qht15AM
xERB13P3bEb2I3EWIXYQ7QAr5xgBzbCyzShPJcwYDYiIESd9MT0KvdDHlJuz42XV
usCv4Zl2b71utdjfoznb/+lugG3O0ymWv0xViazjSVOCQkz8wIcoml1JA49jwoe7
lLnbJysX3TLjl6q3OzzD1u9fztg0zk5jFQCqqiydxI8oaPH1W/dmpWBsL/B2JCXc
EC5aAEwOWU7KxiYr1L3oEJ8mUiE1soPNBX1Btri/BsSsesWdIN4WoIWNCcwzn7G1
iQAPlTNjNDLKcW4CavZThtDG1sx7MweOITlKHUEp23KZ2irf02YavlOP9wjRcYma
j7KCoD2iYZPbkcZIgVQMChkq0kejfSngj7TFNrnaRO6uUPP8ryOrciJFOgbZLDpA
IGobl+MviqJJ6vvsaDi41Frdb5pyJNmL7Fh0vG5xHBOL0EmTQQ9uG8jF23ifAzIv
0D5y7WQqs6QEHBhPhR4qF//KoNQvjY6MdptSnT87Y3ZzObyZK8a7pq88RWrXr6UU
rGMWZdiygcYX12TMkJYoxaf2xXZFujS/np3uej1rfHJBNVJ6/vQ0G+F8uUu9LL/k
NmZHE3reZw3IkSGxH3T3BEYzjIbtZN1ZvaUba5WvT3tqQ6d7kQKvffAGUm3Huhks
4lRl5KYO5c2EwFmbMOnhyYPZAJ0T/acd6bRk6rlG80MpXNaXweRf9QmeD1AY2IPV
MWUFHPlYj6Gn44Z/NmEwZhtzXUnReI+Fe+n7Z11gX4J4VA2jbdmKCW02WRXtK3Sx
POVdCZAg3um0ntraulZCePg2nTFpwylWI66lHRYOXKPPbTeYhUqyp3QOS5q42+nR
BahZSmFkUHxAn6UZkb05DPO87VKKGGHF7eTY4LDh8euq30eBwSLh0v4cjmY6CIbz
fKiY1krf/ADH1AzpwWXcvPz5rlKDnIdx9VDe+mBHRuC/VXCdT5CywhQipqUdKwJk
1I8YvmXAth7WAzJrhCoIKGl5no9+vKAlDZbrem0d3D6A/elnD0ghueaK3JYxYwbZ
ke9dECySqwFzOdx3rQgfXByC1s+AknqXHKP8l9vUXT12NKTnVv40nBfFhKv0mN+a
4+mi6SPS2UbDIGqIqWzMBEGy0IeG1712UPH1EEtXqivKM9d0hCstWUv31iZ73mlq
Hm2jRlSyJvbPcq96IogXxts8MjwCqDFEJLGFTEIBq2pFkx6hR9MIumaqoRCuffcM
PKyjnvZALwdkWcrp8PfyEMZ5dhXcjrbgQssan5GIFERzs6jUVY0jHw3lyDCBO1+V
hc8uOUXNDDv+il0a8l4B+8US5WfjTZEny3gY7gVzSutuWZCv+SLx8PUaTXUgce4m
2SvqOmV4Lm33ibC8HK/my1c80E5PW/bN93VHFuk1T2xSK5zGv8VqT+sPWGtKXbNX
EiIFaQI1xyFDBZWbWOLsovugHxfke2N5Csv5hvbN1PCX0yxPBLGTqI+2P0J8aXeR
PFATmNYoFL7Y/x9Q+2zz7LWcxEFHLbybrHXyV0iEKw414y1PUxU5y3gZgAAEur/b
FFXUNCFMJbTpncS3+4khffIWlyJDLJOOpipNBETUrdrxNNBACfUGGvY67ekD5Ykk
kf+As4KAqrjOyKBgtwd1r1yqZmVkT1elpkEzNmn+wSzQFtB7FCfTJ1thNSlSMtCI
Y+JHjdnp6V6429u/deNINH2dg5S9fhd47IH51ZO+1f4rqJUOP3GUQTyF9KZDPqa+
EgcFC3oFaLdXJRrA4c59EMPG+jNn+/fBJnH7aBKv2Re5KkC8YxNbeJs9lQQo1zL+
Ft1UGreNU86vcApCkxSQQ0d3n221wgg5OGlWOPscZVdtmJOUUUr9powRR8p9fZo9
UFZyciumkpzI8WS7CivIzOpnv9+o6ER2aIffnqk0IdoGSzrcrkaFc8MT/R8tWAYc
iCHvaY3H6jgX485fc4vrYGuyMlwXzMksfi+SW3OWLa4z0tgsoGSdxlP0QiPz2Vzr
RKVz+97MoqdSS1iVWeSaxeuFu7WQ3VycxrvrU2Xa522APN9QAgcy8WvNV2mG3k6r
DDmf6QHOwFShlre2pyZdPmwrxryDu6TD2V7XanM/vlBan5VBlTkFW0oBGEyUEExQ
OxVT6P4Gj1JpQoxKSINSn839vSaM8yNmVo6yYnBvkN9UZ3lPRYzDvGYDOx9tL7Rl
aIdEY6j9SpWwLtWFs1V4jLOktlzwLAAHrVleFV9M/52K9A8Uo7MVm3QNN8UyzldI
K/C39ujt03IFiDOYDm8mk2nt0SfR3j+Ck3Bvxv6evdzpgx8O5OMwzWlNrJPLT7LY
pmBP17J9c0GrP3H5IYkRYzaFfPCRYwhMlp9sMYKPipcUEB/3b6rt2+bEySVW4nJL
2tWBb3RCzr7XU3f4GLp+f7Jn38t3Y/eeorHgr3ctI07oa+rdiqmiVIY3eO4uslzC
EDkyf+wuQN49uwh4BERixrbXBkZRu3slLC/RSYkh03jzkSDB1ZD55UMI4GcTBT52
vV/dGLOcpD8997Y6+BUlx571awnSMXQ/9DAnnTZPohsTxEc4FxbCZ96yF5wAq4qr
CmOqkAJPqQO/0Gre+RLiLSQMfuI9/2Bc8KWDHrOImaPJcy++4I5OkOZL88qXac0o
2DqxYlNDQC/v+IoEJNa1rgOcC+fL3Fs73udLlQSI1K1DtvlMdEutwjTUCfqinyTv
fDHeZbqtTCF3xe+2Q+DdMQMW9j3LhP25BQLvqAIlAITNB5z3FznyOqj8Sparwexq
3J2iZy3sIQ4mK1W3vzI+rGlOq7LQsndzOkG7lSc6iImnjrITF85JoJHT78iJmyHa
MsnCBUGEmpo9JMLZCjPS7OAlJWnywdW71SaHriVexET016wil0l26UqrSB3Dtjsk
JyRffsCKNaeGv1CvdqhzN+Q6j1AUEiiZd3GZsut05mEfRY3E09Gy3DfOr/hT7UNK
/ri0hVATFXYtjcDpFEggiqfqKytQV8lgDx+PoPB58+BAnTrx0ctEH36LZ9GfhwFl
tElO3aXGaOMikA+6i9TJ/RJPLpXg5B4DsvErNEVDmfKmDYYFPlCiAqWEXtq3Z9NV
u7gBH4+LPAo/ee3gXHXxyvEMx3LxHp4xv+9U6UGhLGzi61uCU0TuxVHITFMBe869
zCepwqo/NjRUS0hPd69CUb1H7qDSgfKZoj9S9SbtvwKNSPtNNCdUogENaUN2nInV
cxdkBcAubF+JzranlhlyB051MBwiyQAhbQIJ3+kLM1uILh9hffOIklBFMDIHamoU
PJzn7+BlFA3WQfHljI2mm94t6gXNB+Mb87WTzI6ZcgWP5KTB27m+w3bp6+pKmI1b
zQ3oYZmqp4wxPphrC+BAOE44jyq5hZmZDMixFVBDiBSNHafjPzARRx4bNftFzUW+
cqmGnZhye5LcHKx6Ueb+ls9XQqTkppyBona81zaKcOSu+E3wUmeXdDmPJi+45CXC
w66mAsZMAaUeS0c91nNbFVtDoajvJSFfD3HXM8Z+Po+B9qDBv6FiqZu/7S5sIV2I
xA79WBeLi67Z1OG2pEZDp4KYT0OycC/XE+sgQ+b6cxkI1nu+lpZrrogXo9HHugfV
kNoGJmEUNeOnPcd3R8rc28lKn+JYg9qFbEwdG6Y0Y5bpyF/XoH5QZaKxLhPBStAJ
DqKxyzuiTpSxlrDdynx8SLMMXehHf+U0V9b7uEL53GRb5CX6RnakuXSzHEHtIZwF
+/MLmczUUkjN1a1yGJPw1bV1PvPDn7zcS7BtWq98LscFJ0PKhXcgejtsGXIzJtLM
hn6GVS0hVFeX1+Wx4zdNIpuvsdBp4qzw9t3OQmBAIazojT2xi72hnjhRLXxq4yzA
+PRRCIuZal6nDNK5VxZOHUDSq3opHriSvdjl7sOnqTPiZp+kJy22cvRrobv8QnlA
umTxsBXwRJPreJz/mlUJ1nY6DqNHG7aRJkmGrVppU0yWEmTaSwSQOhfoDhJazqsI
WlXuj1KWuq3OsAutRBJLqKhncRT+wEPx4k63Pvfs1aM4+K4PwzYgsGf+t47WMTHy
V8tcNRjH5dThOOM02itl6deFO/8s/5yxZ+odwZfnJngWYBz2yejkI2VCRCAscIpZ
19jC3k8UwnbM0Z089puw0XqOlqLzz75yHDJepB/CqoEw9XyFyVyZRXqFgVXRsiYc
nLGNkZwAPvJvldA55nvJmt7zjxT1uvsGTZ8lCJY1I+sZcjtJLGBD1tioYB0eweDZ
ZW/sOUiB0d5WNolpsvUTnkFfK70Fobb3v90R5YyhUiwuf9AL4OwSMMOlK72GHxEF
LR/JdpncWkdlTTgA9Dbvu9l8tTRa2ENPGlEKn8qkRSA8+DA9vxCo7R21o9g4cVGF
TWTUYKYna7LZiEO5x9O1Svi9vQteHKjjzWeFv3/6OtWvgG7wFRNkU/qXa/St3e3k
42vNNUnqeRed3/54b9/S4eaeWUui8cZ+BBmcXMVjdPQoFEFnNbhI4bf4ymPUQIBT
wSPBI3nV/mjbyyG8A6SBD/VvldvxXs655YpRwimIfWSwxug5UbveFXDX2ZngUcuf
ze1YVmedEgzaw7yGlGdV5f7S1+nCdHzxMEsgn7DmHyet/hF2alWEBl4JjM0sGGh3
S3xq6S7vUcDX4rPOM52s33XvIdQOq2aj41gTz3hClrxD/CLtsNpJoW/e4XuTK2yM
idPPFiNDb7ByMdl6LvdINzmqi5dknnCFGjvIAMruOkUBQJUEHryLW7/Oa895C8IO
8MifseGJi165siUhUYux2TorVH0LnkWI4Z7zlK5TKG+/7Jte50xN354o1er+D1rh
Erz+4ble/gV078s/pmhf62ARGwlBgJOyViObh7f+jGZIWPODKfm7iIsLOfqEOFoS
iZc21zh6jVw089Wua+vU9hQoA/CgafNXcnj93nC+daRN6WDzzMaloqqr/rUVnyir
B+6PTQbqOEzylLygwI0V7+ovIm/4tORA7KBxbQPuJPaw4MWq01S4ahqZVgnjdtsD
utaJzz0jVG3vGzDLsInX+9jeue/C0weAl7zWD43BaF5/8DzqXIzxxfkkZ+SZi46j
7va/x3e7CUkH+lye+yb341Xzn0VKlnJeh3a6z11wMnG7oSUfQhkQ/2gxSCqbXf8x
ChAv8X4TnEwFh1aBbAGvvB+NpWGNVwps55TSLbLLZPU768qRYDIsoAnQcCXh7xsD
6lnDS1RoadCdyd8AAxBlqnsCfuIJSITxdkV6CeBcT6P0fsg1R4d8fVAXoZ9Ha/od
b1aB9Hct2uhraz3F0C42mX7/rvfUE4MJt+vFYNQc0JKzFymNCQQRFDOnjCaOuEfr
DY3WyaMtcrfq/64iUUInWY3whMhnO5vz7H7OONSWyv8/Ah6WVe4Qmr2B4L3Ry0N1
d6rfpeFSQLKvbif6QJ+b8vcOzCqPbzbMFu44+2QWWNEUJSFFOpYz6dzlnFxjYTlr
0Bshj0jLmC+qyxvJbM+gEApxNGNTCtnOrmMLGWUIu0/ik1oSyJQp9v2kRnLxaMeq
p6kl1qgGiL+YEP1tomzVc15Ab9PGdG06E6YhxIxys8RLuyb1IK5dRb00Cil2Rn4l
XVsHapzcimxLSXn3DM0TLDKxcNKkFCdhdymrqRYB/TSSQe6GTWdP4twVQzGDRujX
cSl/g4STn97blyNdm8QWeC6JmaCmaZqr/RyQE/dSUYDRZPfDKBL+AnFFqZBp1PBS
NPBLRj+eZYbNgPWgfMAFcNfuaEH+lQYb2KE9Cl6Dqdc7gqvG4Z9PakgHdim4E1+d
nxrKhQG/3ohtxPyT4ODufburj8TLeEnJlh+QC9VRdWJB6KQdAMsbzM+0IGRqjFh7
lmd83EuvDG28jCSJQH2Z+0bGT753o1tKVwOHqkgSSzwqMjicnMcIvpxuKjsTh1/r
5yrWkmKUPCKTi1W0uooxePrly6fZRZ+6bXkN2WGpFsjWplgo/yxadlRCtGgjXNLI
WbORWEZqibL9a8CuTu3xTlz+8+b3y4rl/o5ObFwa6eqr315ziHEnv284JoDdW0fK
BYoObgBLtpP2q1qrFyabZ1daXSJ2ckZ849+LbA4+G+l01/XLLJTu4hCKDwyO5SjZ
B+xf8QeU99csVsIVVt/QwBGOWRPzzJN8b5701P0WQ4nM/Acvc77dZQNAQ0qGOG0K
iy2Pk54n7dVTYb+dsUR9fMuUOKwEV4q7HDZaaOUtDSN2a1PpxyRVIme7PFlZn7oU
nU5Ymo6N2M6Y47f5YOniW1HXXy5ByALerfTOtWL+BygCrw8Ne+lUmqmCVsXDX1w4
3AEgTQTzlNZD56oWTG0p0PgDj44xPQ/MJsYaxSoSv0M1+r5bpkvMgFFhQ1frgN5q
vgUEq+OFromONnC8dIaN4oleX4mx8KVVxIoCKdP5X7My4+sOAAClX0Q+PDqJz3K1
3TfzAyk5LCguYOr32yYrQjIgvq139alYLpR1azZKl6bgE2qYzx9rDWC8Dbo+RWG+
HERUexTHt1mlJ/zPmvvH4IYXMornT6unmL0jUgKQxqiL+t4HPGwrrq//vVwX61av
uoJlPnokL1GrQ+YqkkHLFi9l7kjMJxOiv5oefcnm0jgG7f3nFUHZVEuAP+OldWhi
qWZEycyazqnpWUJTOUfyexKrhTlYTZHw4rpNbT5k5LkA55XPTgeC3nzdIcNN+er1
lBuGKNpaCoa4UeT4qe8IzuS/AAL1JG4iuY0F296a00CsqCMA/QDtaQbcg6qUy57i
DIakrEqChdE6weRB3MCkziaOSek8O97Xh+I+0ItW43HkkD2ajMeuv7gP/EVuGuvn
ztXHJ6+W4Rtr3XAW4+Ldvx4+dgp74muIZYyLM5D2omKjRF88xHALF2aVehUKJTyB
vEkEQTOnd0x7MrzS8lTyp+SyikCKKE5wMfoD3nnNkzu0pYwFBgRuBfdddZHgS0xx
kP8zjutCu12BXY4n1FSauhX9Wo+TsJTbnRIYXiT5rXyg2+NjQYqDBkkPECMaVAHE
4wKQD/7FNq5sIPQR3RffuS3hj1uDWv/HfiUY9ysRVACZBb29WvE3HumF64mnjnZT
mnJp6bg7F1VD4DJaRuDXdjm6eHC/vLgOoTXdYNwq8c9FdL97MGA7OLObDkCx4WxD
Wx+BSXl8RupEuxb5jih70bEgsNW2nZmSG5aPaKQ2kdG9GC7aXHH9sEFtKqtSilUq
46kwlyF61721RS0pcOu8XjHqruHePMYXevlnfKRyC2hcXqXrigmerWVABRYa/W8P
pxX4aQbWV1CfC0QDs6zmdsj8Bs/MDixOtvXipRR3AJWz8Utdf8t8AKjDkir1rKp9
x4e0YPNoSbdUX6h6eruJ9/YaSiQeh/fzpWE8O2o8exsv6pKKIrxrRZ6/U5tp+Jp7
Jp0Qe0HMOwnP5OCwaR6hNVpcIwf0SlRe2nRGiJCialuqSZI1IXZh+gHERMeeDAcF
oLpLbVRz0RrVpR43sfIa8ciDTMpPi5S00s9OzYLU8SFIKPmGHALon//iAOO8AL/Q
SrDo6hV0b7+y3YPnVVuvB8X66yogRo6Xf0y+/qfepBxw6Y1Lasyg8mNoUP0Mmbm+
PgqRfV6aW4OvzF7WebCd4Li40aa8ZqUsOTu++vUErV7KUWnCIEIxbtji5E6xOFPG
91ExXGBVpMT9o3z2gx8HcXeUynBOseUm7D0hbYhujf2+S+D+ehRnqs6X5wPpB52Q
W1g6LR3M2xu4PsEK0kOONTejYLMBu/q4RIk75QgEErhcjBn+VCcydREFLhSU+EZl
qOYJfsq9AQ/aLmM+ZoI0ztQzmR+nLCGkyzJqjf8UZc9cm2suOitjjCbbqDTPSpkE
g+jNQXlOkJS7Jxi5OppNd4iOHzX2MWGAggSpOHYQ9YtC624e26DRVOyjizc00DpA
jEr/Vo4WCa8fKub6nWVmgVIoAUkygVsuug2FlK/NPTIlTRiu5Lq81F7m43m9MsHW
9h5YzEn4sJXzEbuf74WU+KIw4s8z4At69ODMBEiNGor5Xd7BxJNI5vhaoq+kJGxV
4QdNZQFnZqouZtgpjqFlDAtBM3ZuQ+eA9XVs4jYp12/kSAA4kuOmtUcK7Zcx1Tn2
cjjwqn/0oSCu2g0KNKiBB6zEMLyRPKjJGAt/MJ1Zykn1rAAGcLVX+yeM60EthUdb
OxqzXoNps9X+v2qWIfCwY5tHmS80vy8Kod6fv4OB2raybv+Y42AA+NEwXshzm/Rz
hyzxgddlTLTpuG5yXzGyMm56T040gUgBqomxXxDP/HvbqcHmq1iER6oRRUQ4EArh
9/yEqMLRBoPiilR/S7TYRC2gq1nlcX0jaC2eR96HxNBKtx/EBgo/WHxiEZKprXwe
8es5GfJ/1SroVKnO3gNETgGXUGwejKCp190NHP6kCCfpqHK6tj1cClGO92WbsrGx
/haNYVPa4VF5kbFMWWd1UkgtoQVWFwWEIN1pVputr4LwVhzUDYlAIayKdODHOlyw
POmajRAzmHMdlvDAzWyY1UuvCTk6uFg7WVytm3YlxPdEXYEcFTLrgFn38mnJROCD
Dg6LeU9W+U6UeHKkrGituQcanuHUP+DVf15Nrrxj0N0lnup9fnWQxV3qFvwpUUmH
76nvGqnx857xKb068+qPFieqsBgUoR9Kg7lm5WtZocYHxaASXHMJxsLQBKkWDlIq
gZsnP6g0VOmzOyi83elwd3Hdz4wgEuA/GCXxNzrQBvHauPULdxL/lmgfnWlzGV6C
eaeiUay/fLj33SlhzFLzMjjqkXk1VVe/bz5jjNpGgfoP5qAP/ksjEy6pqlR0XNdV
X6IxOwn3H/dj9xmbTLDXNUW/Pjc4wm/SoUXH2CJBtmmRhq7qiAtA/Sk2e5/I8Vhy
pPn7MvpSHeLHVi/b4B/koAzTZg7ORnBcbzUrLjv8aQrL7bUa6VJyVJdWEW/ZadK+
wJhAYwo1Umw30HGow13hIkAQ6AH6OhZD+PojSGx9PcY2ENats9rdp/E2UVj/E8Ls
FXdb/MsTp+yjwcYVBKWR7yBxaRtjn722Dmgf3IWsivX5mnx1spKjeuyPpBC6Yq+W
/vpun2mb1qmheAORrAg+W9C28RmTkoBBXcajRyA2Nw9XmCrIGBHUP1IqlFzGSv2W
WodXfKUNt49XHxcLhaFwSK4zzTqkSQofspKua1PrTTMWjkKxf0MQxWxvJggYbv2o
WDLpd2KfiXbYuEDioWGFfhjldAjxcAp1OpPKveB92OCh+26OfsDasplCWQI9QuOe
iMTvfo8asjiEkibOEgqqMSvc4cyeHoL9JnxnOJuM/ee7wuohLpagst+IKqhlNp/Q
WPdPyRjs/GyE4yfiApX59BrV5/tQlyIusQfvKl6cRJ5xbDZ6+IzjQHeR/6/NABZd
wdVLPRpIVreF/SVSKr1quIMnl03KQoCiTUsvgfLebJUDK0qiv7NRNBnZq9BEWbEJ
PjwheAIAh+YAMxvLUX1AToG7SY7Mv6S2Rqj2blA7Mn+YFvEFa4buXzyWVz/Kouce
b/dxnt0qOmViUNo0ndNMm99d9QVbpZrbcMyENT9D8wye+pyXT/zYwYNZvL334DkL
RTHiEmjTNgBmewM4aZod6hAZ2MHcYTlBqizS0DsjXSNb7k7HEnPH3WVy8l0jIZtX
gXNT7uZc3h8XDDtKogx9qQv/H1OESDFvJC9rl9s4wirbcJuo8/DDWsX/l/arqeag
YkBL3Oy7ibKCGqjX86wsSx0u57P+wnJsBud+HSuLnTCtDOPsAC9jzOdy44qq2D7L
ZHuG+PPBrlmHM0UZt302WPGfvs2AgQa6yYclpHiiHibL4W+LShvMeT8QszJKDrec
/uQYgs1mtzrYBnjV1QQEGjvdMnPQfvDwb23VfemGLWpFiggg6nGbQrsKSmDxijT7
uVQXUmtFUMwTEBG5lUBGb0+PrG5LrbPyQSR517eZ1/MS1UJOZJFrTDdq06h95IAE
8dAn9O6JHNx2vnfxZvSwTb0CUMO86zkUynzVOkwfJ3buGooC3YoEaNO3IR0Sz+ht
AnhFafkdnkLTdxzE4ArDzoc9bqSu+Ts4wFAewGtxS6Vt9DWOJkopndYPFsLoC5qf
QpDwnHlQmiirR/QX7C0fakHWlpEoPq/KGgI1K0BEbpGh5IMXgw6yJzPvV55qgd/U
3iJPdDqURHu61ECQSMXVCe7I2WJ7FIB6hNNLkbze8ul1a0CDgehFTfaLNbaPp666
Vf5dB1cm4Z1dzATBLPk5S9a2bD9oTMW5yPcFMZUiTb6h9TDMR3BWEXXbU3MpPqG9
WxAKC7Wved15wsFSdenL8WsWQxsNpusQq0hzE95kBS0nOA79D8LD5IyObd+AexkB
1CZFI3Lj8fjsk5pRtMd0q45UIb0lrdrbsjXJgzmpq/MRpyL2GSkUt1pXCGE1umqF
WITMK6SYdYqWGFA2jsHe1I2QgBkv0OQwEjzvNJv3iSjfVy4Hx+5KOZcnKG+tzXc5
bj5FgewMdQQ8gtVlGowEMerQK47/GHSMUfVOydxHFKqyDTY5l9JcysKn06e2sS4l
GUab202EPY3isYqHeXvbnZIs92edeWJU2kGpRrylH4BTUAMfi81sdMtlafLwtzL3
IoNaV4XCEHUXy3Pv373XWL5i1LGmgG1bz3aZ6rksQDmiz3yo7BKcpX0yb0XQM+I6
b6vFLI/V/sEpqBhNHj09MAH5tizPb86JK+d3cEEzlMrpjHJXDCFIXcjp/25BdBsA
+j+09ZLQMwfgaNqGtKPH1BMJuiJtJOS4F4SoUgfZhhnRvTpwCGnd7URwEqRqOcsK
7HOc6aC44GBA15iB2OfdvW/KMDwHudyrZD9cHj/tCDqD7wEJ6K4KYjnRBUHk28vh
+aIGC1w3EJNfbZIbAbK2fz65aqmFYUmNl+WzXE05jZvStOUga1Y8Msv+XLvB7Moc
0lTyzldToOl1RFSyLY5CRDHCwGiq8h+EfCJcCzn8dMkDw158LYrF7Qmm2qSZBhmd
mShkyDMwjjgIY2egbUuSXcYAQReJg2wSNE2rArRXrXrIqFoJ9nIc48XgZpszU6yF
UVyWPyah1dcOFKTfw+jp2GCprsMkzJ9lUkDJBpTGTHs2NFuy9ThKZhLM/z4uky7q
KkNp6huJAWWg0yRxN5m1QwaqeUM+R2YJ5V/jop4xC/4GvU7ljR5uznh5i0cMDkXU
8OdNl2JzwYzKeD63Ta4NWks4ZwSBp0ARGI/AK4MO/k7HFrGwKl+MOaIOeEv4rU8K
wa0W42JH4iEy6nkKGGZB4FaWTIHbx7bWanLYGwahuDH+UjQm1Ry3Rvsyl1p2fo92
fPefQjr7TbzVVkaCkV0rPnQ0sWclk1S5HzaVsSeDGn6iiw9ffyqDoSvdV9qeWD9Y
xobE0Ftwn10OFDD2jYRhIZqCfQJtxwyqDZ4CPlIWbU8jdRbrJTJWoSk5Ec5fOS7q
3GnRmXjQXL+FTUsM+WF1szlpq4IY71eP+XagAJpUKojqMwLbRglro+ALgK14dg+o
aOWNWT/B3NGq75p0uJpfOfnxbeEzn5/YDtixCo99sugPisFHRxaemHJ6anmsjBaR
ZfShxAw9PaO/P5RBXVbmZXdnam5LeoAonE4OxjPITshWZVqBBlTPLES+mytLllgl
vz3Vv0bn4ZNZbLiXNDAPAuRy4skoV9n7/9bedQ1RKtvMcx6o7jx9YSeE8wjiKOQw
9g52pdOPtyxwpoxJWKznz1TFpaT6tWqr5yOjyLzsq/zO8ny3pcGE2bsnRI5JszFE
96lkOcvAlOShUSBb5ZZgKgkvds0jhrsM21JNXFIJkNEgczl3FctDwP+AEE9tQnd3
1zLHjlIaHjDN4Lrj0a+O2IXdgMIUaH7QwRzWcidvCnhzDm6oZHwwfieaw7Gm6JHS
OT1nSRsN2haGZQjzd6CbQgyS0iVgxCIDPj8HPFGP7JuYy3LRkAl6zb+epB/yFjY+
RU0lF+sBPoSfxe/h/D2aE+PBGFQx9SAj561lc+eVDHNnd82fl0IcWZJ7ye77Aj8q
WBuX7mVGjxB6bdUBDQzFeub94smPK5/SJw/Bx2ZmulShJQMDOGYVXunY8ICoXg21
YFV654oxGZ84u6kd49TilNjFVBGvlA/njCro1vOm2PaGQij4ObZbLzBlVd6AVZeB
0NsrCmmZbfdinaJg54qZeOdzlcM9aOD4zagoFy2Wjzfg6WTldI/SORjBMzzKAuAE
Qb9VOscBtiNpj2TRWG0MCzl4eWDS2J9IHtz0WoYbLiENOew9wHyAY/ILShiwOMc8
oxryrIeZPEoL15laM2Tn3XzewYvcuOZV0VF14b20Nvp7pwqt/lC4w+mPNgdfBcbr
6lhFrIGLpaHosayqYeRt5RY+3FF++pM4wJsgZ+4ko4NWGzCBgvVLOuO8Oa+0qqFO
J7eZ8hLASn4XnlLIfVB68Kn0C6Pp3r6T5YHWpB9pX71ljPfQtQUTj6cYjDYNFZPz
3InWmla8RywzcisxrCUUXROcVASZjx8eGcjjQuH40LPVCPxr0+oMujrHfXe/QiZ4
0ZjdjLPq4SnT1srbYQoY/mfPGBfMz684RXx8pi9dSYovLNK+d1cujHooOBdcccpF
sODndEnQNfwWHq3XtIUlUhC9e8k5bQih7V572YHYUWuCx6tx7r5ZDX6nXQyJGWFe
m9/PcgzXgP0pe/GReJn5FCgtS4AVp6ceGdvxPOdwDwQbb5g+waW8jKl4jwz4deZQ
g5IhxYGqg6W3ygamYl4O3N7b+glM5Sf0uYDAFQERxLcgy0jqaCjvn5eaUMYYQrOM
7MlPMxDp7nMmIubH/0GhHkoiAv4gCeH/AX0Ce/rcfVwQAXQ/9OmYgaUJZ6DCOqy8
QpJ4cUpNlBYESNm7zCg0N7d+MPN0gTs453fOjBspavL/qdFnH6JViR2d8+X3LNW3
yg2rSZmdzv3tyUCxcBBgOuf+/fqO/3YtafYadS27sMeZpBzISjEyc7hvDsOeTAZH
kODGBrp7SEJibEc0iZmNZXzThvaClmoj4tmD7xykjTfGD/w45Fdq6YZRpPYKiHFv
LwdE57LemIz9wDiN6vFjUOgjraXfusFNuHjLuFW6VmHVOQhfBsQgvjH2DmX1H5ir
ZIG8BCfo5wEjPibJZRUT4d/QbqI32+fQxcTXeyJPvOTXFG0ppSUi+a780pbzMa//
ks4+8hS8LhmCaMdhsHsQoTJdaUTsqh65/3bWNn2dxDJWzzMTHZuKBwRWaxNajRnL
Cg+kHiJ8pbxoxCFbEq+oPljcNmQLeS0eNYF4M9ieKMg7Q6XalisqOw1dcWQTSMjU
3DCDeq50dYk8dJcY0PLPvw9RldbWNy+YHb2hla7wY3aL+Fpja03qtlq06BqX6x7O
eU+KyEsveJvHqjErevzULkUj9XAHyGfJiLiH3+TvpgoMciX3v7n1d2Dvk5dj/1OW
LuMeipugfYuUx04NB8KQjaYNyrpoLVkYRWDUk95HD1o7wTVGfktoBYnguVvKLpPR
+4lTfCcZqzWD+jgwhh7rz5Vh682TZrJDworDmgkW0iEIlYH+27GMxlzE6qkn2Cl4
iNHl6+Z8PUjWMkROW45qSsI9Z+sRA7IhlYqB/7iwUucrsxb8j++XOxylF4cfwa9k
WzDpM+Q0RgSCYlUwLFKW7uTN0YXINMezHjF203XRWH+ZoJPsCnKs0x584DAUJRA1
dlC6fuVoUEF29niypHXokzpOADypwdHAJpf35vYW+XYu52h1/RdYXnQR4c5GimL1
2POaUhR1rdakaUBCPe2yCEea7Wy99ANxt7KJH4wf1624xKXsapUDf+t2IhSXfRri
YSPgnALZwOUqfuPHpsZ5BbslBJNl//lunAa1SXgbyUFRubEFiPNzIm2D5jngBJNs
3j4GAMmNyw/Bt5SgwJtA5nBONl5Z6lOtxBNoesy5hq0xU0CL+ZSN02UBs3beILHh
4xUDCfqgPurxUP412pHjlKCbKovMXdmf7utsfqxWJL+a7nFLHG5qReX95+wuoP32
uO6aLhBvA4QjeKNVn65Im1sSbEz9ssbxxsw4nJJ0w0ysnkCZ/YYfOO6XhUQVYun1
ndW6qgkUBiW2vjA/tsJn4hOCcmtXVvUeyxfKvh0TibSS/rPAAnfTHHs52dDBIl1w
vW+CqFryL131QsEzz5W9LlO7TmeW3UJhBJzDJRQ6f9zDdyvtEEisEI9v6TfSbHRs
19T01iRCohIFcj2wkDLgIa/78TZnpS8FtL8WIFzC2KExAjTJqEpc8fFEn5U9SF8V
8++uwaRQAjrvOLR8Z+78vCjpFcQ/mh5k48a3aK8mk94TLhvluvIGfhpLuix+vqSC
qR9KbYaMt9/3u4I6DqrULbNzP7FYXWwR0yaToZctpwdQqnDybhML1iWLTf5Dbz2O
Mt2GO72ef8ql/NgrsivbeJYPmpb6xbfMshc1tF1d67xkIz0qhlP51qq1a6pWdvjo
whtl8ur8IBg8Ego66pOzV5IorWiwuNai01gGI/WYPvOcTGzFwzTkYZBSo6Pbs0XP
OKUpxtvdhE3Y3DOGjpz8akEzspcb++os+owsw7yISTcl5WuhvxIWUvVq+Ls1b/0z
kUko0KPe6dX8sZFeTccptxMU8yLx1qm73BmrucHiHKDq7urwFMLwFRZjEDDShlXl
IazBMjoKZm8jFiLUEKNpEBe8j5/GTRBPXPUhphi17QKYtIuJDErNgb2fKa8kDqV6
hxe5Rn/o7mQbYrP5FcPvZfDqSD1F/MrCuO4oK4sOmLsiEJC8zKwksSltLs6uS3Av
iZW0WwvD46Hq+3YzmEgSnw1/SYaRWpp/qRJ0oVKHOT8RVYROISSA9ksAV9SAABxr
BuWdJ1w5RFGopD/3czWYvsb4xXeMnAHXvPEF4jxzNK4AB/yhBEmysHCKeIxlpkRZ
KKZ5GJt4sWoGOEzcYHRhPYxvqQL1kT2UmIIhAwDQ0QUSqGu0ydKBi3bCnzVD2FUv
IyYBGu9AKkVwe+IYCwceMo4iGVRirBv6qMhqYP1htvaxu4wi8c5GWvODhc0wdqwZ
WdA69lYC9fS9CZ3FXWFNsFiMM/IxcZ9qMlxLkR607KLjWOa3JBK4CBGQlvgDv8oq
7T+T/rRuUlW2KPWkHG9kdgaNSX+iuJAXYKTgnXxSelnn1FpDioum87oJFqsx4bI9
W2e7Ua6U9YX/7+sGc09AZ2CsL6ix/zhXOWa4vVjbOatAdNQV0jpHhqR1cDUHmdBA
xeranneN0h7mAeDcuv6GgsvXlIgLsOpNiqZic/AuHICKjUeux2kJSWI0zyRAlCIE
7QHz8g5g2s0RJoB7k8hRaRPb3Urmi6TcQRnfM605D0FDh0pZxPWbhxjk80Nb8NDi
OXhhTP8BqXxiuizwiB+EDmklbHjY8BYMBMOazdB07BB3ANqIMnJ9nbBLno2gkjin
4zLXSouL7Aw8vUrZHnh2dpGCjoJD+Uovp6oEMmmW0ff4H/qhGzuVIO9Z7Udbf/jy
Q4d9WGTB7mU4zWNGYC/b4Zju/raRQmmgQostNpeC1e1gxxd1kRW1RIdZOfW81mLN
s8PwKAXwB4mf5/n/bFCdKbfVXa3D/0xsX2motlLBvA1leEiGcMso0FQXy4FJZxCx
vLYEQTYL+DkPje+agqsqkbxlDuLBfuTpobIuwt4AlJGh5fvxTRWn0cO5SadOe08Z
Kn0qjGxLWzzsfZOsW9W4XQOd7TsxehCx6e6e0zpYdxv1aSbL0U1KJC4Vc3dzNc/X
ADlNKGKdZuUrlss6YWvI1krZ/QaNMmRrvo35vT9wzsZLRKrN+sJI0NsZUBVIkg3W
KdymXkTn8JCGOgZ8xrPsUtUfUO6NbOuEEc2D9UNRerHtehS+mA6ao089QvdFXu7F
RLSGkiFxT5jviWnsRUCVfdXYFlIzC5C3y7VJX5KRDpTYIXGyEpZsdnC2IBGCmooJ
a7wAxn4H4qiPWkU69fqxQ+vxjLHPRejYpzUlq1Ej1W06A57/zCfTVp+ecDRvVZYJ
Lag1aqWygAhPw1785w9dUVL/nAnHll7vv8xtBaqPxHlKdS1jwnUApQjOEkUpeW47
vmhO5b09dCM6USTQsKtr8xSbEpIC9UxzvfmZrGBqCFNktHUj/e3Hi5kqUJk0NGQM
y1AEAjZgcNArRIcRHbWiY/+O9cvy1wT4aQvsXW28eWMjP3IAnjuCkmyZfARaXTGQ
Uqc00hlE8ewDctdgvCNdxitYw+RGJ9hLtu2BQibfBrL4/YkND7KuXpVAfFoDZE/l
mddW/3f/UUpnfwTuME767nZCrN3GwnEUzui5RKrWbQJhmQ7LGoAv+iBCPI/VY23X
S/pzKMz/A51lUNkuJ8yJfU/HXGi4dhHu2jlmeze9ImomXY6WLpA3Q1lhpYToK2XB
jHo7sW/EX3vpByC0aMFzHzxm4zzpovPLfnraQXwY7M5u63jv21VlRAR5oUrLcELM
dieYSnkjBRb30E74tmEy6XWKKdrOb1u4jnJddazw7nVSZrRImsjKPtxeYawMeATd
seC2iN5rDuvK5W666mtkd0WR8BudNuJcM65ythn9vVneJyRWStAv3WW2pCnEYllD
w6aZiQqSyNk2b+4wg3ChvsBmReW1Fwvc3cQZuSuOJ08rAtAPgZUkoGqea8J77F2y
vUT+IWF0lvUZZKYJcJqsGqLQWB3oRHagGdoiGFHm7c+KoWn40Lsu14QS1QqGokK8
itezA7Hai2DPlZVQG8WEpWJLs5I/OWL0NtpXVJFZpH2zctrQ0EKxq3BiaHxw8CT1
okjFhsYwvXS8I0dSG8mI9ZmjNthGcIWTNgHfB0RRvmur8SgG1T6JwFEWBGHA3icS
Wq6ViWW4p8j3HRNelZoiF/b37kMoY1QZIhX4NClOA9ZZnvUVlzBsF/kjm7E/cyaZ
D/M2wmj6yhqx8Xas443UI5LCFickdhz9QCEVYCg7ya2uGsbWOlH0PjUSzR1+O7/X
SGs+PA45bYZMoEwUMSvPUkbQL2MeD4EcFShIxL4h0WlTLcMwSvAOEsKvwriY3Etu
lWcyhA0cAkvc98DVruOgLr0zDxcvsleaOQ7qGuruTODYWhF6ejzUefF7kNJf5jg8
dWZUfyYMJm6/+MkM2WsyiTeZqRLeiUn387pNrmJ1oo9L/D2Vbs0N7xZH3vsiNvNi
s3TC4SqXsucxjKCBj9gLMv1A5aTVXJDw/qKWUTS+VG3pLQi3QL8yoqUMXDBpHFIC
0uet3D18s4ioYlkPxgX3KY5Fbs5mbu5TOAgGUjDD1t8FaHD+5XicOLTpknjvD91w
/c0Oe1XuEAW9NfmoarosCxWSBkRdQjqLWnUVHnPbwaC2u1SQaW/7CPA6U/Bm5eOG
nwKBqSje8p7T9Yrtk3TFzieAVtRzvKaZBOlFTauEgnyei9l+aRswCy61IHpKW/tI
519wz4fQ8NaXxrXihzMVy3B8tfApYlSOFmSnFpXhfvsFvU+v0gsk8dlJsZ+qnIYJ
Mq3qeVivE7d5xr+amQ7eEUKX+oKe9tNiPYgiLzztjXbmdRBIojGEsKL74aUwJFnu
ooeIO7JkhBAhl0dh0+MiwNvMRqaW7OwiuZiWgYUNjVJxVomQ8SC/8zBO3pmtlEZt
OR1InT7Aj/AOdXR+xNKWjuR7ZQ5xxfME/+zAyuIwjztbkca6sgAQ74KPi6iEnb/w
ygVX4THq+aPKYdwwHFOZmMavIejpck00lg1ou/FzAy36XnB8cQUiwa3kJbUf24b1
F6dVydliU6XEjl7zUsz0V737rOqT2rXSABp5j4x5RBvx6PDnmykskjwEeRQSh4ve
6GvwhEkyXcEixLhW+k9WFFQ/+ofA0cljLB8v7iEVDwoRJvSwG9RKhACO8sWrZR6I
xfogtiEOx2GqcZNIlCIqYhkxyfs/CFnwdIgmvRJOeUmnEiPhBk2sNPGbho3hBjxK
uXQb7SbnA6rYPtKAIjzQPwd6EhWTxN5xC7JwfxcefQRSxSQjQuhEOi+GEV7yAgnS
u81VTMh/XaWX80IWxVMf9VoXpIs5XPWEVIwnRmyP2AysudWEgEu3QcAkuDa/6FhX
9IbGJT8ZP3xCWmbcZRPGm9rYKLMzW2bIq3CW0EluzKt7zFMd+e8+DWnJBAj2kxW/
RUdDe1oYy0Y/MS22LA1nPX4aAlHaSPE7gxoCFP5nsVRXE4rOVKJ21C2qbUc1OM/V
aIXklObzzdJ6dcMgqMukPas/fDPmTSXkOXvPC6iPxr4yDnY8bPu8jSAuoQxef4Zu
cDIhbBz2Z1cfiLtLtHTWTVoDiHDdOiixuo1aZ+Fwcau3i9aihqT0KVsyK/LVVtvQ
3fF6NHoF5MqJAgpFb7Mn91DLhpjVZ+Wvho2UK1+9/Th2FbQbLhg58H3nPZjtyWKS
vOvkCfdkRUbUAAh4b94Lc64tfmcE2jVNhhRKdoi8OepkZotdbma6DW7+u7B1lybk
ONJqb/9KVCCof2kiH45+vO2vKCNllma3h4NnO6LlA3wfsgPax2xc5mYfXF44vRuo
d1k2bUF9FriFUOKf5IB3fx0eoFIU+TUaCsmOg0gE9AxDrUTlaCtJdi6rAXFZhDKb
OlDeNAvgL2YLNVTmL2pklDGsubprH6ZM9L+Owdpb7gEsIM37CAoH4U0x/wh5wGx2
D/mSOqTdWReEdegYd4En3k3/JaN4jsUAU9z1R7hxUZ5/FaPxKE3pXAAmNV6y/6pV
x08Ef7q9PlHlRjjVHj8z12FIuZiKrXXsi+hn7++uFhwT+xd0AEb0tUzqoVy63kN/
/NuUfa8St6msavi5OGGrWGCLl+dWx15Lv1q/YNRcKMYEcMgUQuIOYPI60VYoq3c7
+txpAWdDia3ehLeA/j99/Q0WeAimGMwdh1WiVFNbXhLYJuVc4l3x+kKxbvJyOFtY
CQXjz0T1BJrCEGODCjwD3jA0mZi/xtlo3ikG+bIMEj0QsC5pcCbprOFrokXy8QOJ
3cc27BdPvgQKKkYcBe/1m+0UYoWgztpQuMDfjoY/oTtBVZoJnGnJMdSok6X8ouIZ
xxLErWlMtE75MM+kezuFX25X35f24ZetRxIcKsTdHuiAOUw1IHJ1BhfDSo3vz/68
fRE+EnIlpeLiDTy1goNi89xxeXbJDU32cg2UQ89tktEWu8pN/WEzUK4/0rCpzEye
O9nKYZ6+ea7mOc3itEx/3T0AyznitRuTBMITK3W3zoUeXBovyxebu07wnGEOfHu8
sWxTMzeRjKkkfz411Wjrj8MDduwMU7Rx3G/5zWtXXMfbkkYgsaqpOGYlHETsuVoc
o2kx1FYpifWymE4oPPWzQjA1GRAYQblcH+O27XfkYw2jeVVVm8xVwjyiCKPCPbH4
DcPqMTZVeboWF7/J4UHSVnjVhNJU/smmV0bCkJTnnNmmdfDAcXpc1qKkUdC03Aoy
nHGE8ZQhh0DE+ycnXrTy0RgJZViXE5iEakbA8c+AdwxLzdmF/lVARBKJ1chTAcsj
UTSwBF3t2gWEwN6Ig6xyoFvad/0k0Uf+EQq+FlZmyPt97c1Ryrj2AeOMJWoyNhpD
2iFY7q9Oh+4jywMI0Vj+hl1szhFGY8n116rZp8gMtIkP7cL/rjr/hYpQtTDQYYL7
Vyjzm8aCsdGh2UBATRzfqojrx8IihVRH6RExnnIS6Zwkm8w/ROgruqrSizGE3keH
dP/B3BVeX9/MpWYUTm5x7//MLCKnmceWweNg/VoAWW+bV5UR0FvbE/PBWtPtXuwu
MxS7InJtJyjETvFXSGGXdRJOQQXaBgRUF+Dl/buWLI/L3XDs8lSmOwJONfqcSwP0
z+zQgtcsnNBSUWA7YHx7wIi6F8jXgLy3FbSJTizMjgXrI93NWmf7691H2F6r8dsp
RwO9HB4xUqgnqaA/1U0faceNfEKbMp7BAjlGn0LpXVOTMsT1BDYvFS5KRXT3Mwch
lrsD8jqXjd1BgurwdtR7oXSfw4Ci6HoflaOCe6euPvy70Z7zL396jY1aBLb2rFt6
6sWQseG6Kgwrw6yf0zIzufC/pj+l4H7NtzaQ4IkVZOyxFDoO5ZJbIT93AhsXZjtI
duClwSLbGaTkCxF+s0R4GP4zzTHFi3Ie7J0Jh+5GATud3UmHESQsUDgmZIv+XaH+
4YO3bFvrAlHvyXj+RHTgvHVUDeARjRTTODNAQdYTALxOpcrx/23PGaL2dlE2H9qs
2A6Y1o2xfMnRDFszSpX/FMlx/F3tZNCtZWUUcnkvD+4M6OcactGV3yaNbOOyyuxi
Aqg+ORmzKXiZc27fBB+gS7qg0JtCoZ6Aq4mOvLwY/HORnt7joc/VQCZ/a2hmigUZ
1LRJ+MC6f9Oe0wuI3JZ91NZXWe9Mmh99iAHmTpKUvsQZ5RRDu6qdvMiJ1Jhyg3XT
Fry89J4xcXzQEgLqIVO5GdBsX7jJne2mVDPD5imSHqjzFmyg6vuS4s6d8GW917Uz
LMfLOskFwKk5ErNZMXDcs/WjZ6P6MBPNyZRbwMOWcGcOm6OXyXpUpiRQIKwn/F9+
PbB6ChJPyYiNM6hsUiK7qLB75Wh/VFBpcBlWrVC746mGlL/phtluSbJEV+n0FbSY
XC+KoTyyY6fs65daUdt2Z4Qc2e7Aa9mtBYYRLJS+3amOOvBavE19phioQ507PC2b
Poy3v9WEqdQkt3uYEsQzM7XdfVqwp084qOpKE4emRJr3Org35RaMCuxBB5e9XzLn
2/ISzS6/Q3YCQy7CAcrHvjAPibJovB0gPD39ry3s1HMxzWoc8Kgya2KrDFHRbsdn
mymAHd5Pc6kBaUXd2yaL8LF/bM9NOEra63sJN6QLrxxLZ/8FFsIbOq0tjxMwijS6
FSF4qCwtD/I6Ct16TY28IfCnAuXt88/rtzcaidbt9Vyh+AZTiJGAQgKpfJnJquL3
XGLxfGX22p1b7hE8pXJ8x4yqt9UIvq7BHnxJWmTNU1aFF670GvhL5xLMRMB560hO
ZiXO/rCTfWNRBRS799ksAE8vdGM11sI1uxM+f8WeLUUaVFE9fl2hPMS0Yj6hlNDK
PaM06tNebd/HbRBzkaDClKGnXMrrgq8z65pbaCH3V3NBMyqjJuPA9mwwm0uqs6vH
hxNZ1RAgOwg35olsn/+j4IuyJ7FrdC9arFuGKVrXKsIAdF+Px99PNU9Gwkd99JNi
+crvOWOCBT4oiod4GI1nhqxlDoMmbEBY7n0GAp57ghp+BX/4URmStyya8RjlBpjd
++DpxtKZKt+BnDJQtGTKIvoW2OHSK+3rJjFhAC0DC1seF0RqkuElLyprgUo+kBGt
nWEuqg4FItGjlxSvBUEaOv5xaENZaJuLR1YeouST6aVu4wCXVGHjwesXqIi8prvy
T9hfOT31f0BWf27wiln0NvBgOGLqzpZ3cbmWUsiNAMCIod2vjcMMKmumqKfglOiI
41Rq2fue1S7wUkvyTYFSxejE42Tc2UUXJzM8g6gOJDd45vD3+VK8mqX4r4O1kgFD
Zyq7R4aMhNAebmj3zj1FAl/VQIwlcxmY85CwB+TeqyhvUvCo8IilnuS/UvWFjoX/
4F8+WZ4TAXov9bQYkqg0XcH1SM417/z/fvWpvivfEVPA5ZWJOD6NGiUNUOwlws25
7QtnZX2aQHzNrWRst06aFfPVXV91YYJJiiKF0FbRTHY/2jCIDG/51MhKNaXFCm8z
maoFLZX+W79wnI5KsfjZNWEM7UBhTxWjTlT8GB5ejqyhpU1Hd8Xt3afWtig2a3AJ
i4HcppesRimWWgM0E/mH9+TE4bHYRSqDZXLv/S7d0rETv6C0fvTJ5EBQ5LVLKMkB
4Oao4qbxuZf2GyxCgSwkQYycOcEXlGgJuQ6zUTFrQrs5oNnmGlh00sObpQ78A5re
h3+ABtX+3IhbFxAeb1GZ3rCFt1kWf/6L+QdhT2x60w9SqckIlEM0VChnv+W9eKdf
kS28edS01Rruvkd4xBKPibQlE8G3D6QkFDDMx52r+wMNHFTh5NXGDE1YriOTgYLL
ciDocmgMBLZ9UyZMH3KJYDqFKNQTp+zQsfO36oN9BRUiwpBBhoQGwpvyOGvGKTI9
S3chW6noNJ4p39Zu2Iy8/+RT9gjlTV8U26kbON9BbL8aHkSWcr/iQ97Mpnb+1+ds
nXYTsNO0gYzvShK+6SH+VSnJtqz4ebfuzSdm93rHb5wj4RndMKLwSkVhDMtdIkKT
86KUYd7mW9BGZQYlrgg0yfduZAyVUg2v7cMF9kAdB4zHmry7paT0GZU45RGLjE5E
1qN4lVZA6bHYbJxbPPOyzzOPe0o9C3GzRi69wf4Cbv4bPMEaOS0NY7I/nrIrYa83
9thjRuOj40jC3JmbTq4n00e24lPQfbhgx6ymayJdu4fcqCFfn3jnGVQoj7kDBWuP
bW01SkFjwSbh3Ag+uUSkD7PS12HXwq/VeOWOD6jDbadJPjOgR0lvKWzJiDitdbob
0jtxwl55oWC/0XRFZWIgUsO3z4kvpwxzIA7pR20NS3kL29ZIz5k38cRB3hZTO9AE
k3Qz9uPlloEEV/YyxW28BylNjrex1ycbk6G7qX5RqROiHrrl1yn9BYePEj89SwWD
hYprGrTIErrQ+Jw4ByR727+HKgo03eL8dM4ehecdWuyb2rrF9yOJTEwAtrkzn4EQ
xFOV9g3lriR751yM4hvjm7eUdatMaYe/+INSBEgB0zKB+WqILKmgrj6t+WFeaWEk
Urvwu62uICryrczqMP0g6mRpJzsH4Csm9nSJen5ZenyJK5RnI/9PrecUMlUU9B5E
bJ4IVnFznABkxn38XqqPPVqkq6ezvod3lqj10XQv3DGqjJqT5vMezefptl28MJlX
mFd8wp+cmOBNxFbejL/IhxVFv1dmBrxwcMy63uKU+FHag5iG4gRPaPUyEK4du0IM
WeQCAlhqrZqzB3vVNdhJjWgDQl0XrwYFHkCyTDC8XxSHb7IibFrIuMLuartQ69YI
IjOgUdLJjiBx3Pqj6BFi2+bShCoJ/B2thG0GOaAQem8gZUSrfhSc+EiQbQWGXkgL
qhGfZiZHXq8jJQupYZOudNTOL4L/ibL6lFz5pdUTUIadQnsakvWfCr5DTnPijh/M
ZsxAITCchl6bF1HVD2hFWG6G01kNXoSndUIsRsj1XAeAAxBKVUd3tR+9Cr82wtlc
UsU9cVsHQ1V0dCS/YLqlYc43Jm9hXXJ1Vk0i+mtxIOZrmZ4dact7oZUptJHbdflc
n6viuTokDdMiDcwaWJjosac0EXaVvjfqOJk1IPdqjfc7eRBvklhfv4CTbm1/boac
2h1mRF6UXOlXDgoZxsB1q4CYpdUSJ0hH6QXWtNy9kToHcDA47ZrHA1nZpzS6uXT9
upY9Q0/RhDtbEAWlCWlZaGReqeUoKu2tLvnD6L5IfViNMFf5icIO8ENFN0bYzuGS
H0GX2Ihzg5RQgKEdu3ogYFZqQvDQ5wEceNLCI3yVOkyJzgdvweBTkJ78NebIdxkq
BfnI3hNBfVjVcZihvZprykSWKg5fv4eZi1AqZ3fq483UM5JUpLYV6ZoKjct/bbx4
egC68y0NiYr3RNhaUmeudleL3X6yPv5a/raS3kDH/llf/1K05k3+zsmeEUjf/TvV
ATsY4P37AiIV5YLh1O9Tp8DfHlJPzzng+HJh6MFRMw2mmreVuP6svLY+S9BzURfh
Xp9e4u/Qj79x1LOys62DrUGhWe551saL+mK2jBFjU7ApwypPBEGzEuQFpKJHcOi4
zK1zZXZlpCb9hPTUYtQURRf0osLGdrpkTJY3QMeGfuMq6sKkNE9OuozR0l/BQT4u
WMSQnrBQwV5e03G41UjmGWgaUy4rU1he58qsaXG094Hqy3AH7o3a+AiRZFOMrdie
JzDqf5wLqby87qq0eS1+MOiNYJcKQjzCW2IUS8YBKMxb+kSax2QyOEYssTj8lr9s
BCRQd9CsqzG7wYYP8twhpI/uQh2YFE3LCo88u2O2OIrgz7NzNuRbPbjqU1YKsC2K
/4BGhlBlUT/LBFIR/tHdM/awfqEXeuUfDgWsDn9dttTN5wZ+nIThvtMYXNiEckFp
mbgOsFhk6hkj6NApV2+cLJj22NN4QrUv7NrXZCPt2SSQqxzicWK4Re4H5hkch/zj
ddv0h+h9xF5Y77yCvmTCfeiZFZhk7EHiDukuCmDCF2yCdTg6/IjmdKJf4IfLs/qz
H8oRiM7mfuvycVuVodJU6eubfRLdvsjdXxUyCCI3P5wmHJByW/hhK5HYkzlP/1PE
/3lAvxlIBmicxagsvt5mbOKBB9UWyWhLaHgrh1TECuY4ns2tXlYD/eh36whoKWJB
e+acyyGZhthwLSZ/CDLmT5hH1ErTqHNP0TW8so8do3pr3VFhfQBIVrB3SV1Psrgb
WNrs4JPzx8DQa65QtTd/8ILYRQBcLLUErafvoj7HEH8IR9L+6oWboXUbSu44PV/v
7xod83r/tME6ND0r1OcTeiS8CGo3X7fFaCrjO868R2YrF+pNQUzgMlTl/m70jq5K
BZUYwNCuIoQCD7pEA+gJ5hLWqTUqNxT2cKIJgyiqNZ69CzZXsxlTfWRNqszxPnv5
/nFX83rTlw21y7M1MLv2zBbePamPiYLz0YSIYaEUNH0v9rhthXvaY3ANEJa3PhRS
kPUaHQ3iDvOZ5CWtc18kT8ryP3LCM+OlXlwA6QNI8fB2S7K78GTSVnN5CkDeUXHm
cBTA+1Nr1N33tm/tITz+tD1hLi3MAjV+Vp97BqQXbIUsGWSmR9cXDVH8Fgbc0JVb
4SCdX3mBrumTas/6P0sFMC+wM5gD5FQAi5Ma1zW2OznV9Z0aKwOca5IrbIobs352
KKq8WxJK0kL4dFBYJI4rbAoLj0Ss+eJB1L62900r1mqJgpN0oyP6MjJBP7iDrnw8
1RQ+t6+K2720ebjKFm46GN2b1S1nc8wn0/EFqdYvkmn7Z3i3uaD5s6qt1sld7ltb
sqPZTPSVj9A2KaGZ0BU0MaFrOxTb+7gYI4dFv8xycV0o82SVenPmm3mCjVGsID5b
NbLk2uIgwBWV6pfj3cTPOkYRE7OPhP86GY2vzyT7tU78ozBMOXBng8H1EQzkcXum
Jek+hmA4y9dc5sPFnXMWBfM7TSVBxBDhlgQup3XzYlvguOpKZZ+0LY18FshanYAt
GTgpohsbdJ9XYQ99SxGGPxdf9AJrzcZvLUHl3vWucQBU4J3MKglN9tTMBuvxgYPA
e6tTVZ0VRXM+lrG7vNIYPLKADfQfQ9SpRb+enMajkqlrQ/A2IOHXKhE7m0nQ438R
/6YdRRJqqCeIow+SR11lhKyfHXOUFf8UUJJ3c3ezjCEoL0y/keWFmPx47zZG31+8
NcgvgE2adMh+8xGM+nRQScVGgDIePXj4FRXWO8IldbqQ53BKPswJXJWVeISvIN5P
KNAft+gXs3lmkMNuqMPoXA2BZSUJ4LgIt8XHIpUNF0PINQWsD/z6eDrjm323lK4Z
K1KKVYmKI84/ZmSE2x02kKPV5ET5uAGvKO3mEv4sevhUSQ67fkvqDziQLQC1Vqaj
QUS1RhGXgqKXFePEUErbTh3hiKVfENJ+wtaGfzsIPPw6jvAzvLAeP9ehlplyOBQI
lZRlAx2FNezD2YwbcC/LUSCmT8vUPPiEw+OO7FszWa9P5x4OEugH/2mB9iAqZ0Zx
mf/eM0ioyUuumWHbO6ufffK3+ZWiDeU8kmFtRJWB6AapYhuOum/fkkLvVgxjTs+h
ZED7pAp0rb8sdnmTh/2v4FTNBb4rvlsELTLngsrsa2Mhyn68WMAOb0A3O8jCXsv1
b8NkYWbIk+3WG++30LBvluHm7+RMQQCpYaSuMmRWFzl5Mssn6r8i0Z3xYgXC50AU
FgnTITBfd0X106+y2retzkoMG6TfWvld8YUVAin8K/Y/9Iz5Zs9XbfKb4Rj+QUjf
uTeWhE3+uokwEdZdduDDSrzJpxysIEJ/QwAlGoKyZZnfT5cp9aazUjapvhen4Lv7
ODRcBiiWAJOOYl9XOWrKjtjmXkuUbeWm8y7eL3YwHbsyBITLVg5LBc1n1thY9q0g
SHxA1Y0EXZMrunOoeQUdQ+YCsARB0So3+qIB24Tz+ZxsuQVALjGLoa1pwF6Bii6P
7pYEWU22D4U8CWV3m9QIX5XaD3I4mJZ3T1wbyvxtHBqIOLfsm+VMnHS5FFQnN2eq
ELq6tlzJl66jaXiQ01XMNZni21Mkkk5ekzmdRL2GwSgmWtHSq5hzZ1PObp+Ni5w2
dLmpjAF/odvsMTFyn4tuNfS93zpfydRXVE5B627AI3jreVMjXI3d3u7mjVyFdPEN
J56qpdFnMGDgaGVWBf5pr5N8UY0aoEqI9FVcngb32GPma5f5D1uTop6my46Dvpnu
/+BFO4dHVAvvSo1dsWzT3ntBe5X02sLsBNqjt9UPMuFZmXNlWT87si2o5bI1XutM
hNjAQ6KJsTztFYyRgRbjZxdT06HIL8hSeLcOEdPZQah0MV1mFC3HrbTWLC12gIKV
zJ0SCJ4ygw98nJ3DB/wiWO4aVy6Cgto9jntyGvqjWu94BWyJnnKKm/SBtq/sdmib
RZGuFB1EEBFJ+1SUH34+HoisDBicIsagEcV7wVX5bygKLxuMm0nWF5+mPqSuOcOd
od9MteQLPwst3IKBAHh4yYY3z1+s+4p7e82NPKT2AlgGrXwFIg3Ofw5nMuOyjoXu
mXqY7dVNGIOhCCIdQD1AnyrNWy4h8amDBhakwnPBunvpSggBPwKSNJY4POiUtJ/i
hXBirK/IpDgYhlVPyIKMQ26+hy+FQ1dDwJRq4fVsZcC3b+6k4L6ufF+4AiPSMLY9
oLYv7aBATNZnUr+tIGScwgl7eYT8M10/qNkYY186UXSutmgbwure9WzLX8MbErgF
wvSKrL8JEVL+WAoLAgWO/Tpp5jTNaDtOPiI60jv8QaPooedbtQI+tP7EzSNi543m
CpA16pPgVTQiZlYc1Zn6j4lwFgKpZ9V+YmSHvKhHjYzRba59sZCuqOHt+yY/mwjr
kmhgWhFCPBJd+UiHq3PZfUXnCd1I44OQTCvduNCyWteEwf5wX14z5Jh/dNoDe2qG
Ct6dEDPFJr6s/l2EK0M3Mrgri6noRrqHy3Kx0gog8ws7Z7+pJF5tJyD7Sqk0Z73a
X83AjTyc7BkBVAdOXcINPRmJh1vtIIK8D48CGMd2rcWCPXi5X/O+bnYNqRQP3xx3
94yw+3h2M6G2+ScjByJJ6TZB338LNxdbkYdvQAMa0SQ1JGL2GiV+qtUdTGFHTR05
1MeN2fdbsK09kYRk66PHv/gPjpkJf91EvJ57yhYnxv9qF8Espe6muonzNMa2NKDA
50BCLLZ925UEs4LR2nyEaRv9C0wYcNZXOdG+rkIGQYUrtShpAPD7dr63Uhd0eY4z
la7VPYOkaTsyG4QIBl5xKMdth7JPzWicAUAls5Hm8DIJ3uODOf1s41PorYCmEkhl
sd76HPC8SIf81X9pXqq8CnGNBZiwFlSzhTYrFkyuhzoyDuWEJdyR950+Uc4h3FuV
vcRHsIYIWT1Vpe/GPy6X0LwRcV0Ap4vQZBewuaUWJ4S7esI2XtwvstNXuDGrcn/C
Xn0ucH0MvMKCJbLAZRZCoZclsWykhdqHQC9o8vs7aM971s6hOniSN75OUHuA9OLi
cHxtSkOomq7t0o0DDazI889RODyQI0mjshTcl6fmxu9beJ6TOu0Z1y4dVlhlujQm
NUE3vdTX7O+IQ6I3KLRsnN8pxqghz1Rzx/fHXLj8bKgUw1b7WSfdcEcMV3iJKcTG
A2WP1yphxwTo2MTGCBAYDOK3MCZmgTSvqWn5V7/K1EUh4tyuP/iuRuvipU4tu90p
gFHjG7naSN8wmcsitEGHHg2A2K+3ZXVLnDQiRINdr63B+KXrDHY6f/gAgFZcYK2B
c/rG9AoVmFGac69/RYD4/EeeaP3qjVL0t3AEm9tFmdEu2MYTgv8zFipbVvA4XQNJ
U8LoEcDjZAbSziTHKgxnObzVDeIg1hfD7XrBjUSgekD7xW1V3U3J4XOfV2a3pZiL
OfEfpp1DhIpZ5xtSfgeaR9aaNYuZswXPfwVC4Y6M1DZnecM5ErQ0DZVp8jy99c6e
cAmcVX3rxXqPg33sfNjdm4XCy+qlro2VqwTsGy1iCnWVAHum8DJ1tebvolY5x6DM
toyV9t9/BFd6npG1kSGAOJBeJAzfv5nPIpD+Rl/Ea7qRO4NRv6ToAsxcmY13KBI2
Jsy/md+EOhxlPHKwqp0KibyR6pHLrq2BMROEdnnfBl3qeWiI3ApFC4wTdpE/kvty
GCPfvtTPoT2tn4ZY664+gctDTg6NeJz55M9OSjSl0xnnchdR2qFUuXTjTAjHoU09
n6PlGnMm/aNY6Yv9g3xGGKDMHOTsQjNO9jp5TyGJE4iJ2hf0m3Vm1dNfiv+ZX4M4
MiXrrzyxhVJVDYH+G5ARrxxOu1D+vJFkmBsUlRLWNJYO3YV94nus0aIXQScq3p+L
fw8r5nIErI0SKB7DMPSfymz/A77zm5+h5a0zpudmx0qn8h9EkuZ7t1xHbydSQnbH
Zwb1bXLtKAxp986+mFMLxV/s2hL01K+QKvAp6E5GT/p4r42H4L/1d/Td3Mz9NuWW
QeYQHNK9KsNG8hqPDvO7lg/dqL7rkmw4M8c6Nh/iWDRdtCKZXgfBZvUWF9SRhWeA
kdqHoiIK//3dHBlk6XNGVTiwNJejQi9Omugs9h+a356gVRYbYJCYoLUzt33XdEuh
81or9Rxm4pvyQxLctpY7wx47mPdLZarAwCsd/DdrXvmw1Y8VCOh8hM4VwbQjSpT1
+y0Zbah+HWpeLnfiHSa2E0ifxcrfUl2QbNbAVLMAAw2+axPmtljeVloFQGT8lPTT
VrNNa93i027fBe4vL9iVEnP/ILogHXOQyujVoNC16upqxPO7un5cU1bkf3klfA/M
m+x2ZXNP6KRzDyBu4W6jxgu/x2r03PKZp2UWbqQUQ4kkHvuB+/J7pXqKgqMci3J4
VSS+IuBxUnBiNLkmt+NM/DyUDtooHqnGqiKorcA1zQecm4BZ7RQzQ6k4uDw2Lfst
Kaq4qROWw62Sm8BrXh3qHvgnRVv/zR2+6JoR5i3jHHtwravfInjxQoEOWOAWjsCp
QLf5I+9IIncJmwjmJ3c44/M2q0iy4IqNH1JqXCvkX8uHAgq/f8XvaaXFciW4Iq/K
NA/+QM9NufAJriIfXuDoUmU2gLVJ279ztMv6z7cIvKxCLRDWGCjzBEDzRnPORfiQ
Uytvqu9lyS++h+8Ve7L+vq0s7OqD/TsKWZsqgktPFqvllot0+TY0PFLUXMQ7ftYw
xVK191NVH+l5qK7gsvJmA8MWIrR+DksJYIfvdFeyihkZ3/ZDjl8j/4gcPbj7s189
TV4zuXo6k7jMqHfoHyGiELsDcr29lNrfLN15w6AFJod7/dLT9cG1wxQppTL4VvJ0
DhjZUU7/dL9nJNTdOhGXKVhuvSHCVa5rP/Tjmb/6mKCVEIZuYu5VQ8oDpU/+EpRX
m4VUrzB0mAEpMO6fUYSO/V5cTJ1aedbrlNLQC1fKxKJ4NcKl4n5+miU6tlYEMvdO
goAFcnAkHa/DqIzX3FY7AUDPiERYIdXdqqYQjjOmdlLgSlQ+p4zmbLL1VWXIDX2c
71p2spHeR24heZ2fu4Jji2fPSN9wOCjK2e0orM0lkI15fs9d/+n7b2whkE9sDjU1
2hx37fOOgMqJ5NABPJ0iCRhiKpYuzrLIk3RLCuUtgb1RCxLY7W+JRgpqt3PGn2UO
2p5IhdKZ0zLaTfE/iA2LKmDapUUWLQGos6ZeEWvA2Z4cSiUtGo+R3INI2n2SlrqO
mV6TVlUdFF2AoYHKNAHj2mR81/TzZpTEYzPiixdeJTzIwE/TOjIi7d/OiyADiGxc
Lj1US2WtAHyeixchmD8MxsLjHWVNsd5fzZEMke+Lw8QZmpm7xXpVa4CqwpKyjVhG
D5nGeDUmpouLb16nXupkmynSu1sStSdvGAxPzLi3Jl9tc4Q0e7YrUInA60T+ZQYA
TKnBq454z88shRivOIVfzJUEMQH/Q9H7YKuRX0VILzCAlM0SqjSiJv/rYCziVhh7
C7U5WaZHv6nrDEG6p1DV6AiBMTm2IG7AooV51JVilVD4wF5Zm7Q4yToYVGsvami9
6aM/aJMbprini/t+f8vuQPVVh+p8nEKKu1vFfWzZY5ZyLqNXcwwoPIVLINRnI4Qw
mP2vPTIqPuVFnEHcZ/KY8RaEVRs0GPteCiRxVa47VrwPJW7nW6HqVb0xeL0KwE/5
OjKt9BX7WUDpbdYprzqkSJvPM6e70YYOQJK/TuuDTHrB03b4rFbwWVL7meHfQVYl
mBw/Uyzdey/7eBPEnrbLRCG3TSsd9T3h5KbC1BMlGKB2xWyuervd0EXB7m8wTtAP
1oyfRDuHyRptj84faGAOoNfKNkq0taQzo64CVL/U/564MOnmZTIN4evyG3p98i8E
V9YnTjUqkaCL5ixjiUQUfJg4Lo9KW26NDJeUwIQ3OZ0m9YpsSGoBIPNojxVEW3th
ZMVlwXBksYNcff8vD+9Hn02bEq2CLu2cHdWyWqXrdhkk8fT7HSr67SDSyvjJLuPr
d8LsFOnb4WCtMFs45piSeqdmG6rfF3rEl8qYL9iWUFnp+hhYn96mcx4WSy30DgJT
BvAZSZmsEq3phCC3yN6YsgVOkL9Df+VF5uAyQ9SOS/Q8Ul/Km/Xt+4a8z6Pa5KdK
1rWIKWpUKkufOJb7FvDWpr56WBhtN/OPsH7z7jJieQNhXB4OSgq0hshZbR2toGvV
1qABdcUQZvwWP5d2ChKDe+xH06Jzd1Xa7Ugjm/8rEySWxypRP9JPiG+JrrU2n2t6
qrTeMyMH5mmfbPTqMvNWPu/6QglN/1TZbhQMusByb+C/yslEGogpVcnsjSMVOhV5
fO52GkFqihSdfYhMS+X3zBXRMl51CaTxe6PvXS6fZdI9K/krYOfeelB70apG5osJ
srSqXlKT2YcevluAUukGQ2c1///sceEyjhurhrR52Tb/s53zQY5W3sHRljHajpnl
dQR7L4teNDUtHTvHeVZY1aln7/wI4FPl2aR6lwSLSXTt7hush1ApqmdUfmR8ickZ
fOIV6m0d0QEGkvF2B6E3xqd+J15y7GCp0/lRhJzrMLuoEMW0xKV9f9dDYgQ+Qv1N
mXvgokg0j3hjwGL63MiKEzOF5UJhbSaST/4SWoiVLVBErmJQ/KfjG3SfdBSJN7WN
VopWT2lopaCanAuJ+DUBnHe6gH8lPRxqWK6riP3OFhrVxNfy5wHxQ9OJd6PQpldF
Aa+jR+dbcyShGoVzNkeK2HHfPzqSMAhDMT9vkhBWKZ3YWb5Ml2BR5o5O0nbYhCAv
xv1zC6+W9PYOIy9pWdAI+ss56X0dxB/vPYkVJkhEAsJh1lL/c2x4/4A7kLHQ41nv
aZ+/s0fK+AltK/KarKvaUXnuf87hkU3vFN/QyJ6c1T9j9yJA1UjTXKfwhCswRWdf
NioCR2hDWsl4LehBp0gpucqQu7IuWyNKQeiCBIEoPNZJL2Cu7XwL8PBQop8LzdQV
nGDrZ+Io/Rd54Ddd3lw+bbywtpDDABOPY+0Zhn3vfGiND1PADi/GDUZuhmdKP1gB
LCDqk4Nk2aco8B0x8fLf8K97uuilsTFSKC6OLurvVnsWwWWKjMAYWxR97YiFWC+S
SLNoLse4W4CkQtMVTEuoStv9x1jUpyhz9STu0EJgOd7zikCUWdY9T1TlfTXSh/CI
fKz3w/n/US1y6phMi9xCpQBtkmaHgnMDzLKDAyQ//p2biIVy0qjZLG8cDz58Bqd0
9CKuji1BZOc+R/eyLWdsgWEAH4pCLhO2ZEWX3//w7x6B23unS0K/BE1k/7UCIynW
Zig6hypdzxl4nJ8qBy7LbUrwFXZXHxb3DYWSGvK2thXlHA1AwAC0SufOwRLaw9et
7QqfYTh4o4psovkmboS3LkADuxyiTG3Nm/rJFwHBeWd2UVYbTlzJYk+5QP+al06p
SCKGyTkXGvCm4TCYYYZmYhkpAQe7arTloixzBaRMvscIt1wTTAq5MBo1JdhOFH8O
KWJ3IcCGXcsrZujYJ0wlTU6FyCVA07KsOK3zHIiuShrLALQdOh066zN52exir090
1ku/e4myR0zt69Mu2tbwU/JSQrWCGN+sup8KtUTJOB8ZR8jAm0WDzEazA58xlPU/
p1aEITcNHInvfELuauqCmLjfX48vXYtsI+WAYowfeDCP4Rm/nggze0kB1ZSHyP/A
5e4UhTbuzeyCUXO/4CU+R1iBHAzwR3uLamR8oe9MCGBTtpOXV5sysja17mxmQZhM
RBpKszFzpFCIQka31fE5YD1Vv6UhVKPKWIRqnWadXhDvq9API9Zr5WeYXQ3iWzqj
21nidB3Wk58bjdYWisS2BSewP1Tl1EqM80JOZpupY++y3Epxus+dj/p7zEMmD63C
zI4/Qb2sRajrBDRnZx5Hs8GsSqq6C3rZepiun75/fEnh78rMPlSIAcFim4ONhU/J
27IGXLJdochOC4uYi5ptlh0PtJo5xyRQog9IBv0t1eqihfPsjvtgCsrz3YsSlJAk
ptBzx4ky1P5ejxRc3wUEGrB7auKv0BGrnTYQpca2kL0eEssdTeT+cPZLg9Lcng8o
/ahMXmq6YNU7xlKSdZYAB6hsRGty9AlQTK0eK01iCdq++s+0aeH62nMAGyNxAp5z
rA6h1WYF2evAM1dGzv7Edn1VQrjEWCSf2o5FJyU2LI0Lii6NKaYRPDCKw3ki79ZW
rhZfGiTG3wgkCWVyI4bVN5guZNaYpux7E3y97NREW/n+BbHmuvNlo0PXaIlB+AzB
RW9MK2fOto/stOjLZzr6cIS/E+PA/C85YJ1yprsw3ESww//h3lmwb62BFESsW5iK
YavK7HniOYRjCB8jYRtxUUANJ1VGDP0pKNMwP896ty4WLAOmq3/ZA16qDAaFpdoI
5EbHt3HKB+cMAiJlgnP/cBTTaUi2LztW2ngvDbgsYLvSnYY23m+Bc6zXnxoGK/gc
XuvtfiLoHUADl2kKlp2NfPGUHwqxPkuTF4Zjmpw0tOLlFbIflHcyzWiDXBHWqWri
cuOc7jX9C2lN/JC73ZDbCNhKMiAJYudaONdFrLinzUn/KTf8g6LTo4+xAfk3Geq6
C9iQQNN7uIDQHMwa2lKDT0VUWVr5NmocI3CuLflrzaHawmT43Uv2OuZ/32C3ITf5
ri9zewTa5oHXOV7YfISxgSHgjqhkjF8bQMXn+sRZ6sMiNrL+Zt3b7yTWe3CnUxwy
44hB2SpiLTR2sOaQqX+YGdlDXPSE/l1MC9K28KNLeM3qg6J89u/6wd1NpeoXcKuz
l2rG98BsULBqvxCDYaYaao96ibsI2t1Hb4UbCPRhknwRV8p8UbIIxAPPi2rGp3iv
jR+pOeWoGGkhaHYTR3j9AxF5x5I2lAwGArg4D/sjmL8Gk4kTle6AvGkG/PhH52cb
g+yhfHvqQPQIGIzqcj5i3w6Pp7sghrQmNhsXyGwiwCFq3XVJAzK1ja1GMlyGfZAF
xsvIPCcsKsWUxONeH1WcMl9PR9gn8hfZG9JbX61pwB/xyg7cX7JrzCZTIbHli4+X
ZMZ8eTkQ0ce2nclwtxXdGpq0H2+scI1GQZBiPNBUCcQ6BYYxsgxk68VW61HpBMcr
AC+6AHBcOxlBdg9zuI2ITeLgyciV4BAgfMECF18g72F3ItbcZVPT/mGG/ZMyVyv3
M+4KWDkblOaBRCdFrC9c+bswoMP7CiED4C0Kv/rfFhptkUa9JejHhYrb/wCyogu6
dZjaD3aGGSLezfBIGAPu/YL7Y5pdelE/nz5r8L4V81oU0Ask2CDixXdQgSiqHs/n
QlSC0k5CYNKxObgQFQjlpa/isdpH/oxP+g8Oipd3nLQRU0KRwYv5GQWkNR9/L5lO
7LYTlvPyxH2dlK7Jv1m5B4yza/+kmXeRZFWxXWAbUDngtJAtIKsVr7Vm8UIwrTXy
sAV93cXiUqqn7/TVpm2ZSuY+PkQZLzfuPrTpb2ghIvbsJokUwJ5MW7db9jspid8n
N3um/H/LW3UKZ/1o2u0gS2qS53kuGYwexMKvcwjlD1IOmh/gywPWV0ITGgvmaTO5
sBC1EzNzB55uQMr447Yfymbvds6pRc+wg8bv2uj9G5ZWMPT3pyx2MO+Vex99QfXn
veE93y6PIp2Cg85Ath010JK44tOmDzoBufIU9kXMbZvuBLOyp0/NI7Mxdd146uA7
ZfkuyTM0mq1DUGFVeGeu6FiAQGw9I89g9dAIsknvulA0Lx/kiKmlmSESeUGviLDk
2KobSnqRRxWZOArAyXajWp3XrO2GsxR1gjKq3RwBO3Rt4c95nb4RCDcApresug23
xY8XdncQnZcANE34dNEPumuXt2dfz+IWhKPkOONEb7Wf/IXFqInz7YrcV3jXexfW
bHaJP81yooqCUCpcRFfxcb16gqKd0ZUmVQk6dUsAHGA8efNf/ugfitiXwTbID2lC
639Lc66fJMi2794uYXHOE5Z1vjoWFLlVLUsvBIX+e8t2r87avKSVlbkotL9CdkSR
ke5ffhP9I2QL1n64pOBL+UV9z/pH+N7nnnCL7SIGsljzRpTT+NK1H+4IEbkxnpps
zimnlIddJv2IjiNPwrXSvNeWPgaSgEleTxJpYmXrsd+sa/Nev8hHui4LeBgOpwE+
eGv0Kq+nBvIfKYHUdo3ZU6n9tWLBI1ofvodEzzpete0gRZvkza95F8st6E89xJjU
uHvv5ifa80dlqSo345ofLCzvlc//lJjndMP4y0R0uMC79NZ3xQSJTYHrJBSE83aa
9GU6Mu5+hrFDxCHQ59oe0REfCCnUazwB0ZzazPenlwPPZmvPR+GVIepKtEUMLER3
JTyMW2gRJh1r8/j2tV8kf9XtYtdx4fYXCUBVqBTz6hcbppH863wVmoP4xTafRqz6
DRXspdBYBzAw56a42pyhbUtMEw1mWJGrd5tQ9NdDkJVQHkE3ZBcCrTD7ZydkFN9E
sDDNL+7sXFMA1yVje6oG6BQn38Jrm0uWeSk8Ec0z5oR17Fu8EuFJ1ykzpDqQWF7D
kZz3L3azXqr+qH6WFbL+A/0fYls0hxHciM4mApl6aok+5yeZv+8VOHDlmE/TUlZi
uI2Oqltzfl5dXS0FMtki1NJMOTQM+f9i+sZiQKnxGJVC4i6KuWHUrFjgBOg2/P8w
vNd6dQdffrTP2Hqhn2lzHvBgT9YTt+/SjqrGPT7WRs8K3UYvJhZ2kXAyQzNFEz6f
LRlJZyc67j34GYtkk8V76tevSre0hX+G+KdjbB2j9a4ByhFiHIJ/MduSFgYzFL+P
elUcWgZ6MmZWqg/8joDY/r3hDlPd3jCpsI/G0bntka9yX6KAGV2U3xZzh4EnFlOT
5YpalueNTZChugVNMYQNl7FsBHLmPjQksFXalcrsCU345c90yKbJ/nNaHx94tTcn
51nSz+HfiVHIWNpu2MB5x3QY3aKuc6jrr7FM7qxvfrzMWL5V3EMsbJzVwOpmOPxC
bwOhJ3WTEkBijvB/ISARJERw47MqRKn6geFvvm90VFJtUzbL4RBFDs2mv401IhGT
JOngjHxnoJ11TlpsGhhyfWLxtclqX97IJ4pEbYSAkT37Itx3qp5WR9E5Er5iwYIh
XoAV5/GeO2Aqyybi7rYzB6B6+Ml3RlvOXKYrAm1MRRuSIG8/yWzQJujgTcVEG9Vr
3YdFi9zan6AJTNhy/zIMXu94mZ5jL5fvU+memdqhJcdtz9nv7ox6Oa2rzqEzEf3U
TzscHs1SU26K4jU8isqjoq11rqMf01u+Za2pOGjBmvMrF/L3Fqy7zP43VRcA7iCF
jOSRCWSWHF0Yrk1urfNqVIm4Xhf1phrkxmNSCvjOZzaa7QOkd8/xWsnnSP0NGikQ
cG5kjsZ6kWo7QihFuc7EIdx65JOKjfUHtuvDYxXIaPzPReNJfN6VFepqkXl1MD1/
/K74M22o9VySXCfqwAmKpBbAoNNSs9Ss6FL3bqBhBHORgiRTRPnwYjlkmAF27jBn
K6DO9WxbeNW2R/csoNVI1OOGTahTwgCC2O2KN1utYA4SR5M+gshG0f2egrKQnmG4
1LFiMplqra+tGmiEk+nrpc9IuwjxRPy9zQQ5E117jehiCDWBisRG3qRWLe0qii0y
e0+WTRTuWBvDAWzGtQ+oBaR3405qEXmw+SF+uHT43VrHC7s1rUIEluy/I21AtXZr
+9dapJulkWU8f1s/XB1nw4vahfaN39t+VyrnGGfih6GQiGtXKBgmTkNpuu65wuh0
b5K+U7VxDZPONMoHSZiLJfVUx/4MwxI0+nbU3fWxlTcM04GQEVhx5NGXqccUkwXE
fqkwN+gbKFO525fTG6B6oWCZaG6I4ZUtKz+UGIppdD1hrJ0oIf/eyCoFv/bLWDQD
cN3UCtryq7YCWPNROkW8q5QVDXIsZ/OFwQiMvb/oeafZ1wMYFQzpiuh2W8h3YsIr
ZU6jKd3dPOs2O/akt/XHj4OSWGFlbYuFatbdsKoIRXA6ZxyO+wNP9cnv53yFO+PJ
g847okDal3L0HDaskl5G8Zj8Wn5OjYyrWkPmHginMumpL2u99VNriINiVSDZ2vHa
dUPKusLbS/Ih8IOz69X1nubcItyd6wjEHwt0ZcH954M9nB5cBPoSRqf4Z1mh3kBQ
FasDQsoXJ0JlDO6e/e8Yd1eHTR9wDPLCGjLA52y5qaJV6vUVy6XN+ODjVXhf+xwl
8vnuWKJ3UWG04kREP7KOkD8PT/xLAbTdOstrmlu6FZt7VNNnI2/aPq42IzMud8nc
0su88gc9gIr9p9Gs6ZdNxAs3K8wx5BHjad8xAaCtiuXYuxVtOVQlMCx6dhMnRltx
fLplrJ7Sv1HWiatiDP2H43J3MgS0ncRtA6rnDfo/jjZ5OUnK+qzV5KuTtKJZoA+/
0d37NMN34TIsmvYodbIhhVxVhFiASTdt5vXBck2z5ZN2NddwhyoDAr7F/7nx+y/r
4E7KUwlHD5+tAHQA5h3vwOt5Pi/xhbRqxdvxkET+NVKyIu26zC6c2AC2hItk1asD
4PSIJleUVzc0j1FbeO+ROYEyeFDvTiZi9du3NovJtJvGkEclKVCHuvN5WKgPFjfc
YYyXxGAMU8g4auluOjEzuvk9Y4sn+rXsYMFuvo022TsePAR/QFcC2nptNN1c4Ddn
cJxIOKI2/ZINJUm961PcwYVfGSN/okHcKKfR1zA+vWODRTavDiJPh/v6EydqClnJ
53bOUXtCZsV+jjgmJsPeQj875JqrdYTh587Ot4a8UbX0b2l1ce/+GztTS9dcaYiV
3B8zR+Hx+rWLq/4okgTqXuxEZv/aQdfhhfrEghd/fh6hp3EsMxlgvg1xM/68l/rf
1fHrY1dVudlXKzExVxouhJ/fUZExKfCOvJJnT+9dBrSeqDKWcpjhUcwWtpf0sLQ0
O8LihkLLck5dMjiAUSrzSHZOcfI+nv3shqgTbpJ4Ii3qsmaEHFkfNWQ7N+/0+Sdq
jG2Cwc0BEZr9z0Et85Mrcme7I8+77HIhqiFFzjUchwIiyIasqHSnuX1FvahRU4kt
ZrZxwzO1sjQzsHPs4Z3M1LYC3evKvLbZFJgKXLPsdQYyUyyUns89JlrjyjDE86JY
02Y1SdpkjnslNekJnxykBpJuq3tZUD99+Iz1QdhbCk5aAJMG7AP+d8OEYK6fOe4b
Ab+jgWI92Z3IH4p1tdcavpPgnu43Xu8SO8rUIoSnyONjSKAW3jARMwqpekHKU5Uf
HZJFI2gUIQWseG6r/Ild53NJQTxFUKxjnOPTaaj6ykYnKAalExkU0RK4Xp8Oo+JK
2PeYnKIAxmrpre3duGuJbUKxs5/4QBv5fYFM+p4lp0II6sorx+aBeIf4vc+oGmqd
SFFXM05HZREcA+ltaWG/Ma1OLjy25kSCeP8JYLJgk3HkQCakkDS9IqCLzUcyM8lx
LtIqnf6HS6jom/kOE8jSibW7U8ydr7VIkwxUdU1iwMJzK2nXa2RNLk/sHtzoUkSz
oFhIT6AkvwoT2STMawQiQn9Pp97fD5XvuuqZ3Kyyq5FClG5aWoWyEz4stOxP/4TF
HKPQKbW7usSjRt6mVRSCZsd9LZA5i9E5/MjMbU0X5hzHMY8ZWKSKH0fOmGkBAPxq
WBVUi0ON5EkZg6unuuEyFMIGSNAlCSN6hlRVb86KJK1tg6PUew/ExLjxn9Ry1nGz
ajdjTfjThAk3MNSKiwPyGtMNRItDgwp9nFsJvZkrLC+8NTBdl3zZ5DunTv3Qfs36
YeWKf3oEihfTZejG3bSpaVG88hQMdZ9wauNsS9/NmZ/TGFmHkaJ2IIW8p5V0avo9
eDJWXOZIohtHgrkmF+Mj0j7ZCxCqYDrbSx1akdDSv8HCa888ggPBI3ltupgzlEQZ
bGQpSRJs36e2+4Kq9/27plGEkloQxuH8EXwYCei651BypeTjGy2JcGubgD92VZ63
hFQc1tLDus+6EanzM3ZaznQk/fU8PbBFew8NcNucsZZiYJEoeYxxvGe1d4+x0LVA
9gfhQqsK8CDjU6Sy7pSWAHXBNOExbCYrTU5ZzMgPAf3xTY+XAgdwyMugdSFnjBnN
gFNF/VXeXE8iK+SWr9zJdkM9AHFbVoyRLfZ7zPkkidgG6AC32zn63h5t0lNNRa3H
TTP3rAE+blg6BWL/AbFoyXz8rBYNFydzk8RDoQZ9HPB9evZDjIdorZCIrPiE7hKi
L8ewwDjVYBg3s5taWLGekYkJvVL318e2s/3w8W5z2665jk4SNU2ql4BLOorvkbMn
rxtB2dWTjVD6qQSGkhbMIfL3ATO1sk98cQLYZggYR3cSmTbsBLozK9qzfZSg98+y
CrQei3IImh48SSy7Jag+wfc+QTEcSfi7OGGqJmK5FQaYLOdrks35vO8DFuAg/AYU
lNNH0RuD3Xs1isQxxXbWzAq5KUqZppHl6/9Y5PPLjrHHULc2/HxXefLDwRKtj4dL
xB8cqm3ZkRl9sDYnbRxrWqlw8L/ka48ufrsyhEl1axvWvC4iI5U6dYvRmAxdHLOQ
1bkQZ+Eb24Dz3jUyxqOJRliT/WT4F+triF2YU4pGwhyQnn0exGDbrOiHDEJPD3z0
hvDNkTqsnWOh4HjI4uM/0FqkLmwAfPXtHGtcfB+dMZ0PUnBpx1qKjPzpD2i2zErX
xIOEBFsdFjRiW/eXavN8fa5xYFyWgRb7vifm2jszk7xyo8Wj0km7hUMuMIceTmuM
HwKMQET/kzbtVVrzQraq9gx4iAwH1Irvq3CyfwSMHoDgK5073umsHQ3lmmVdRnno
D8Wj78lzd0TlCZcDbZ1dINDRf5wiHhuA0YaudbpJEKmh3Wy1iV9HEtNJv7bR4eQP
JA6P8M+KdiLJ3bxstwRNSMSqSwbyhrpooG3StQhuUOU664Yk7UYAX1D4LsgrZsnu
hYSUAZNWUpNNxTZY+6AYlI0WFZI3dVpN6+H7RNRoUPuc2GFqiMfYismQGcSRoio6
HQJz9vcIMxXABp7nYIuKf3kHpnR/g/1BwosGIt9rdeGkPp3y3ol7QKu2pBjiBnsJ
qiv3jCn7l86RkLo3koCUK6vqboW7PkQpA1XUGouSSxFT7Gyb49uKpLsmnDo+j1yU
3ltGSl/HmpE8rYfMRotB+bsc4dNDnEQUOFgtxuAOHvP9gGhX+7Ouh/arG9G4MGvl
Io0AVMZeFEt0kNaG2IxsM45XOhfJhHSUiRLYaqM23jMzVb06ovrYTtRfw8KUqcmv
06pD8wm420RjS3PqHWU6mmSLbYntz6JrNnCbSQknCPblMUaIEp2kLc7TiHwjMi3o
8DSUZGA5nZGFgs2K/nw3j+kMZ/XhdRUyjcwdkYiX9ZYyl9RZgXK18AzaAJYC4Wli
xMwPLeUQ1z4xcOBlNZ0H8hgUVyjczwe3hkZtBKvM4krLA40Mu6+m1nF6QpyniES3
Ko4Y026PB5TdPeCNoy12qK6DyIPmn4TX9vEXWG1a9IREpreJhKY3Nh+QHTMFMgzD
IxJBxiWFnKokvJREoMUDCq0+FWbSZG9Qr+bJscf4iBegcC+pHmoeT97UvrxyAPlD
EMFmGGAdoBbT4+PXxWRThCd5pBWBxNrn60VSL1AvDzaQgsIhP5nfGfzyEUp8iy6V
Wst/teFtWaS+xnZ5rDJqMtYbQfngMoauvudDkbTwvlHZqSm7M/NRh+p6lQ7sM3B7
wmQUxT7krIkgu29Kx4i5d9/nm5eqpeMsWyI03T3cfIYI4qXlhWCyemjYHeVNroQi
142c0+R7LRfAo3l6iixn3pb1cMkGcJtpZwvLYI83vhz6fVzjOOKn2CjcvYsyT9Nq
7CTyF4REEI8SW3M6JYsYjG9txO4Kr5sZxZxI7N9LdZs6Itz+TmqJ5K8yTJhAJaV6
8mOSaJzp5yGRDfOrjg/rypwM1Z8/fILoYyxW3WZE0HX0iMJnKGH2oDekjACv3duf
YCI4/TnCXqJ8pqsS8EOvdxYhmt5N/QugHYBHvtXGTM4e7FHXlasAJshWclXCiUGW
UuAIXSodf9JnFAeAWHJcDyVGUWaZTXNJU4V1OHskq189LTO+9ggoTd5ZQHB6ymO/
cD57Wh0o65P4tPy8X/OWGnDwWTgR3IBRO6gnXGDdUtWl7AT8zIJr1z1ddzm0/cHe
AwsUaG+t2neBx/IiBbsrEq4qTYiVHvnCg1Vi9EtoY0A44GK/vjhywrtTmDpJ6+ZL
GNq87eTOYXuuTKam232CzQwbW2E5qYXG2HqQ7guxZvRp5+k0S0b/mVQu3g4eQ5PC
8d6G9/YvuLChBgoYvM5Jqp5Ng5u6nEsrN2zZsvh/qSYfh+rTv1xJZbyYWjOlm96H
DBegvTjimy1NguDi5SLE7FwEnrBfR03KhPpBWoOJUNY9/chxsVtyxWAK7pBFI1CZ
HIfVpwBkU37f9e6ovLda1YERPeiVvFInu/yFDxQmandvHIB9gIb7huqHmns+F3qy
xuwYSNi7QIb22lsqY58vFcTSwH5j8SgXZtL1wq5e27LsQwM2va3jBYG6skE628KU
/oAF55FmNTKyQTrsuRUnZO6Bdp/acavRf2pKRr6BpHn3hs28jESbAtzk3TZb2NoS
LOd6RLmAtGmFSQAZXE9QTcSun79KNEIno9D096DY5OUc7cXK1c2VQ0vlv9+LmZYF
Rhz7ZyAwaHITMQnQuKLiDUkA+rmnZkc/KR9Qe7ppix1HgwXgTxymlM2Wvl3IY+D9
FQl2/d68DyhEUEbMgEuYuPgNp85urzuNDTYaS10dRe40RMjaH6m1Lh627RwPO63B
zgQxIWADJROf7tDwKP1PyxO9HBQHpOESUNlH2GhIVdl5XuBYkLa3rA/KfDYyVkrI
tXOv4ojlcwKqkRFuqwLgHe4WdSroOMsYhTntPXETisEDM0ZHvXaN0W6OEJwlQiCJ
jb4EwZl1K4a7ppHR+h2q0QSjkT+tfUn5bYU0T1njtb43OrxElZQwq6RwOIRBODLO
Y5K3USjlBgDuTbloIP/FuFGiQ3d718PaOUP+Q2DOCyakSnvR5SW19zKmuKOM2Ekh
TD/YdvafY2gYISmbNDXBBFZwxlNGzEE56AFZdUahRYCIJNQI9H+BlZl4s4cO3Tw8
o54pdCtzebNYB/xfdUza6sbt6SNBLlTYApBmgdId/ishIWehvGKNWyxHj3QsqISW
yytZJzNRhi16bIKbVLdwQvD1xwhRdH2HBCocfaQ0cZwZe2dtu1p1EM4NPLdufNUb
VS5SmmH1hiwnSaHfsSCkYKT3PmiOVvXorVWkWKRZe6kftHSRkoKJRoKo39A5TGgV
+zawZAlYRXi1OI+MdCnQnxCpEW9Zzm6+0NxsPato0D2FtSysIapfdQiT/ICRPctf
H9DEU/j6WT9HtpVFy1n4pXy8BU7C9qbC0uK/Y4oa4IfHeKTVqRjyDQymRFITm0G3
+yMiAv3PUlP0peNUw1Cafs1qkBWpAWTWjjbBoAethXz9KpPqNEnRHCk/Vo7egF7+
eQPdWFMuc1Z0gX0T5trDyFIo4bB9BWyMk9iPbjQDRtRpNCSnlXtj9qyYw96nOxSd
bJVK0BFvuZANavE5uuXh93R4STP8TgwnvR4RxpsqqcnU344tG9lPsZXt40K247WW
TLKBp0zhMhBbHBET4y7nEREG1rpZYBGUoOM7Nc5doawwjXQc2kKRhJuBdinyUJ8t
ZZojx0wwqudQVrKodtSYHQXzYTDJ0Rg/Be7VXtNZXVIDJfqPqTjd8rVgjvllSxS/
bCpmUxIYXQIO+ogkpK570Ew4iLyB/axrdhKj9qsFczIqf3gYbxrY5TwffzdZ6wtK
Dg+0FpI10JHHI9i/2T0IO0LeGsLe0fVXkLk6CGaWVj4ldY61FKdBRyuiXgsIy2D4
AnhunpDHAJ/HXjQpaqNRyi9xfMUUfu/VRA46hIvRIXmV+rEwE1cfQdppcZt3I/Mk
5Jro3+hxzge6WC7ye9eXXUZ4m64mML2KLm/4iOMXrpWQQsZDkmvD06VHBg0/G+x2
P0wlJoE1ZgAy3BS7myut4veJkRagTxaJKJ3lv+gbmK1F+3L0iiFOvQzveaeQdpxV
5yKY7CAe6LWvV5YnAj3ZskgmDH1lTcwDE2p1wy9Li6T4dyLmzkPRpkwW/zDJqugd
7D/gIn0TSIek4BSD+B6I28Hidva5Zx+UEUJnANQvXhG1sshrSdTj9sXM7PN0jFul
GXbfO0zV2VbfWFJ6K05AQRmshEm8UkiL056tE+WsdtqmJGIRzqkNQnC5k5uJGt1O
4CLAJ7Q9Z+0/c6rvUZ5TVh4PJQzn7DbVjnU/5V/OXtsBHHRK2zhzzN+8awOFXS6Z
IPN9dTrc6zFWp8gFzQ/9WFpc+IRarXvv9spW5Xl/JCDnpuqlOK6LzZ9iQRnhrups
givYd8DPzXQpuqdO5rKWgZ9aTUHM2Jse4ohbmABcp94T5THwBPlJWirdC00ib7mv
JhYYuFZD5YQoa1iLNtXZ2DlDH/HKplmnxnY+LuDJNJLlsUVnmQ4ZwBLfi7DAJSeA
KwlbyoZfxPMrScxrcfUsVWvcFHnVp2Uj3QuSlykTpemKWGIK1DL4aZxxQ9UQC19f
mCtMYhbkTXCVfmxS7WjykPikJcvk+pMuSBdpsG5U9MQLH/ZeHT8IP7mY9KAJPd5S
Z/cA6WzrkSxkxXAsQ3BLBV7xIC97sqcmDZqNitCzDVCbEYXf8+70YEumy/CxhXR7
owlKMLWRGcALHcdFonc7bTYeg55p5iupdLTLli5urwuRN3Bh7jaTpgCVAYu+duKI
sY2VBNcKu2AM70bJOYnBOdVtf7emDhHpJOfzI+V89QCyPKhhfBhU2Y6NlK7+ycNm
RHlU3haQnjldktxjrxcxqnFd1JQCEqjlUcBD35Ur7k23z+y6snc/mrea5ZC4MljF
NUra0J7aNcgsHXWCOEHW2GEq91yT0IHJtfw3mWrHA6v5/GcVUPLfkAZEAiSx2Cl9
q1hAR0XxFSVLvEiceLOdwb7p9tu4hJtHhSIwNWtb2YWApYkZkoDrJPZBMoRVYlwr
gS/Gkh8ZOUkqyFeyn8asJOXpyPn5GRwIibyl7q1m3zXlVKe5PRQRS57MwFshYz36
zfZGjBf1X0qmZimsrh3FkaX7bOYWQdjGf4EmOokW6sC5adjE9aRK3/BOA3AOYVOl
jDxuVeu9EMjRPw/yWNeIU1e1CriWT0N1rW6vlPPDDGF6eMXVy0LNes8Xyu0/Kwyx
tI9H6rz9rIVBiAxt5lKl9q/Wp8Vu303qRoGGTP/pmBLgPV4W1DNHQejRSAwH3hfd
UituO82dvTYksPWzXqXu0Q71ogK6eFBXvatlL4l3EEg3AnTr03TVqSxDLNUs//qk
qhLcrvzn92TzV5zUuElf+otf8AlBwP94sjiBLX25ze9NartLPLWVT53dXbCg+Yka
x8wLD0+rVPqsjZinmmiptg8IcnnNZ2iB0TVl6vO9zWEHmXMLPGnL/IBhGi7Kpuzr
h7F5Cu+cZZ2IgLYyg/5pmliPu7td3ICyrQ5+iXPq+4+9SoT4CspJuQ1WPlNqgYnC
R25KfGGyAzk+PljE2xXBt5aYUmjBvdhblsyLOss3FpOR90jl61OdtpcOMcLFwVjX
a2sVn/lnxNAIR8UkRBNgtLVXAdCSOGnQwHUaDdAR0Uqi+Pfq1ccFvKp7MOpiyzFe
W1AWECQKHFAB4dCDtnbH+0qfDawwL7nJLBVKSv7iQvEwbvqy+OwLI02H/8cQLURZ
C7kqIggKDXGaOhrHgZ4CK9JUK7fF82PlOF1WK+QlEWZYBXp10WnQNMIIO9n2kyF3
w+dfmyHkZ8P2ufnwyKhXgWKmQmhYe6IW0R9ZhVvKUVPmZ2oAXk68dHnVFmvjwT+W
DMa9cKG2/pkF1aL+s7rJT5OfgaikBiRE1I0HsdLIfwsLnE8MKZSRAXXd6f0H86eN
Uj+T1/WKRAjfPSJoGDl5vOtsxPfu63I/A0fW6Rew4+AuauGbN+hBs0VoT+E4STeI
o/RkU0jnd/8FgPR+bq1UW133MBNUwkZX2kMDFGXuoAPWyBpqEokkW5bMKJ3UTafp
eFVUKMb45cFMA7AQ40wYQwnugGhAVrl/IQqDZhfoZEFAA0jFumuURDf8ZI/O3zQh
cetRiPSNx2dW3bU/cld9sot7Ngurp8jbXsMEWLsHHGMc+6F0GZpUBlb6qdsOCzej
qBVVPO4hjqzicxyZ5xKvYpS8yHuuW1p5dFWT33Fbm/VD4tWqJNnPXXvPRv2aDmRx
WjujD3b8dsOiDdxQDSaq3vVjgYhNAX6/vBcTlcIWMlamxyOkD+siEf1Cv8ydGvCT
3OU99xxAQpcoSO0v7AM65ALhLSuxCwSJwAfz3OtVoAcA5qpZ2eAjxnLC7doPcKOn
6FUuxT1upIwsS2Lh9htQuMhOefNjY+9putng9Ab1iDTiuTixJU/EWoof6Gd/v1xM
RykYkjHQDaOqyE4tZ7eTqrJ/gYhvAk9pFNcT6RNNUe6wlaxv0uYQ3Qus3LxrU2we
uc6znXkgW0LcQmWLobvRI8N15jXo5/jJWijeMgUSQyxO7CCK/TiUlluD5sDy1Z1Y
Vr+Eu2m6uiCb3SX63uL9BoxKVipGTi9oo0EUF7aSa8+3aAS/9LIEJd5wc12Vh1cp
OXN1JHDLWjF5f4u4j1ALIa/eMEWUGetPIClV7l1AlaM2bEX8BQIXSIf8vOTQExrC
P1nUfGvyuYaev9ACI5sbOxO91gS3r8auYUI70yl9MQu6C0+qJ4oqVkMoFLd5/Jkw
+Ir7Xh0z7dAPNWWiUgc9vXazW7B2ggbZfX+fJMCvd60aT45Vya+alkdkFxFoPSqI
z9AH9hYxbUvSQbK3VOkeHW/6U5TmosxN9hNQJO19g7R1yCsh4TVjwZzGQKpvLj7e
ltNiHCmdbE6Ubdavs5zLRMcMH17asjH4PHMPhKTWus8p/szCDawYdDybyh9EJDMO
qFhrlUDx2JpMc4RGv1XCIRZJ/sLJe0Vb7FgKe+Vgf+m94SvTlG0HxBPldUaFhEcB
9aO+kSfWfWrp/Gjx9oj9a+qMC6TS4YBM7QGaMyw4EjVPK+yzhSI+Q9hSEOTbTmNe
EkSPpEjERO0RXvdtfZfmZim3fGdSFxB0Y49S4jUklqwAu7B7EwTha4OzvRORDgOb
Al1fMI40Vs4zrZmZsdtJgbJqxdVvOpfqLJDS9kxGmJ++8tYKBXfaoCt7pQsnnyXu
uTjqPm782cACNmDJQhmju+t5XAJaGpqzzYq6eQMMEz559MkGjpBmJcrErBtfmO46
Eb+XFUsX9gvX0735t8n63kwu03ag4VPnD+E7uqpSdAO0jaCFltZGbjsfP2B5AvJj
IU/oJumIjeUMuBlH3Zt8SLjSu8kKm6sfqp5hG5RyAcNN6VWnUNiUGzce7XO+miWD
u8TBIL61CO5H6yHWPZaStqy6u5ivUMIZuwHTVUx9c0yrllfATje7k93baMUmXAMN
Qvok+wAJuzsskvSRYFkSJhlDqLqam/07itaObloj5QKfUEK9FgXZrIP0uQnu9RTH
fOmCxSNuGxhRHbDj8hB9sSfGVcTI+BCRdtBOgx1tgvhhwUFITI0kXHrjTiGZ9gNj
xHM5eHL/ZGBubPprpjBpTubJ2UGPlI14tcO2Rmd6/HaHFom8NXF8zm6TU/y/+LPZ
xUl/M0QXWjRG7k6ZF1lGrrBNcm33/CSki8NiTxKZNR8ISew7o/SB55bPWdqLV+2A
0b6nZXF1GdoYVbV+SK+nJVEkzlcciLdVWRadtiKVDgUvHmjikczVpxmzOTryrnM9
9QUWlvcHN+y9eEaIiuphvTRKEQ0XtTKpsQOqrs+P/wuFHcGSSHsZxOSmW++q/wwq
bhHeX0Q56Rejd+FkEpsmbxySzYSg0Kmx23jiget/hVS8n5ExiU8zMINWgoTZKxae
YZ+B6Gi6+2LSWkvqBbrVwqKxc4Yzg22sUjAUV/A6dFC2vFzqQtP9a5MNi0YXUJqZ
grioPeKKm5wkMyDmjWOw9qjO4Bj7ri950toW6gWD9KMKaehcIKaRRAqqNleet8X0
VFQt6e96doRZLai4v4KBb+ji5jIsUWG8cEXIvFkjK0Mev9wt76IPTlamMaujwfAP
KexgV/bNPrtfV/5pJoSXD3MmdAsNCw86/siLpBReHCPT+U3g3MfEtE7Yr9dGwiTL
Y++bqU5ZQ0B6Tt9fl/+rXDDQWXbRNULNgqQja9CkD8i+BZue74OswWDC0mAsKmAI
6TfuN2p33rS7uozD/ABRat/luAIhayDmwHinUPWtg6Bl49qrDrl9KZ0JhRUI29l0
Qc+r2aHEqN42gBM2SCKwDTTTl383Pj4k61o7xchluxAW8w3P8VwcQsS4b3QyTxX2
cQHPNQwNcH/427HfMb1IytfBbM6GdXtnuRsscjy5QRX6lcjPCzDjHGof54c4NLDf
Hu6EgR4NRvujzjHF+HaBrScJlSujrMHUuEJCz1BNNUcHbuq3ys3vHZIUxSJd52R1
6dZSmh7EKod0zLy3VzMAMvjC27e9OJ7yWqVRT2PPOhfVmFxu30U9tLitfv6ZLHM8
7DSRIJoI9yDxMsP5OWp07uNl+wtNgsiTFEbjF8xJcU+gCdCoF1OWowzRVAjlN/Pd
HFOjKVx3fmdPl7Op5SW9NY/gRtzrGITVmXTjYp8yoZg8wLvNKlvKXcBK+LynRb+s
DXymSRlveG9fzW9zCI1RK67Z6k5agpVhprQ7KxP+6U2MfFW2WUz5me7mTSPQlf2H
lTkkL+aFm0FZTg5HKcPXQ1E41TJvw+UCHqbzZ8zipsM9we1+xpMtyOBE1WRdSSKQ
2NGqR/Yho0XsKJzT+amQjvPRtD4S3o2FxgRUMtGSvfUutT2b9sjS6Xekcguxu8IS
s6BRQWaABlOSway5HVDbfweehZoETUt3CKuMLT/GSNI+c0CtDswEPaRn/zO2oO2r
thTQpRhtpGf4Rhy+ywyjjfqsSYeWQxHht4IuTfr7XNnuBVMilLawpZnseoxdIaqP
TnsLeu5pf8hcLp+MlbccagnaiFoFdvhJBJe5gMgo4xDRJHqBL+tXJrXQzdLpOZoM
QoGvSEb6o2QXZzHy8x27RZO/UHHq3cW/wqztBCAxCCOFTBxrRrOk5sQOYCxTKi5G
uUdTMHl2W1I0jp7BZcYKolcJ6IzD+ceCJa+QgNmnv9chWQpz8zG/C4s/bfCXGoKK
i7qb18mi6S7/u20tz3atuH+sgKry6flKNtP+Byf+3bc9LqT4JcXNwDVMqrXXVIig
35pX/qzpV+viaY584EvxnBmQLBT5F72K82GepqvAMJpwUIZKIofsUC5MIPM603LD
5FPogODSdyEPXU+g68fsjAxcK2ykebXCZ6sjDtPzQ7PXlpGPPqrTZjkUKY+hPOrw
iQVtvboyVJD8YPSP691c/1oQM4NtuMbUBiZCCoxXx71ejpiR38HtXgYCdl/ghULr
tjcmfNjhNAlFBU6RWwD0kDFXgETY75zk4vC7R3wpq47Ugo/mnKf3K41Bcbes7XZA
UF1Iqkm8+YcJSW4+bevePSt3YELudks1+Lu1ARNxQV1481RHqFIJJGMkUcs1cNkR
5KYiw/QiIHKAAxqDJFIHtV5GBgN0rTZVkYyQcK+sBhe0vNFo6TYjED3NOBrtiXrp
PD9HxfmC4OoLyovp1eogPnguxnrwf8SImvCm/k4H6qYxIaS7B05ZCrb3fgc53bYo
LOUxKx20Ue0lRYQIsFJ/nrWawOPiBe5XSBxO4RuIzsFMSPqyK/UFoMQqH9Jiquwj
GrOIpYhBHHqY/RVB6wTlDkmSPnMHAM7DSNTWvxXELAKIM9jXFUuaHISg15s4BOqN
sdK2bQ4OivMPrxorhxAxIzrY9+S8qY0EP8JWqnOrs1T0pFiFdSRPS+cBLaZ3rRRg
xbkwMUIxPGOa2PwC+RM7BBrhdFoYTJ2c+KbLg2V0MZmbYOcHI5EiLPArg32X38bT
/+A6nRDdypcy1/rE3GRoxv73eRzzDn8cF4XSB5DwButtreCg2V446p7xR6n9rXbA
vxbI/bEkUabS3JMCu5dYuO0N/LW8PZcezpMSFsK68IJ7Soh64i6L5aHC5xswTdPP
UAd/uPlYmGzSyfjb29Y70HP4ZQL+ryRH8sE6hmMjp9H4sIL1tbIz00pRByqp6vzp
R4l1y3eEyDmIka4EXf+B+ZkVNpikIPOK5cTnEvaMUuITGxy7ObqL7SZNBk1tYqwW
t+qZX+5jAYasNBZqJMMHxMXmrrRR0u8ygvZgPmJ3yUTyf8lqZjtSsA+f1Iu8or4R
fcHjj6kHBBZUo6X1P7f+rdlLTrRsZs9Yc8ZOoq2pFhCbj+TcJZaMCTmp8iBPjE2r
jj2PMg8YNK1GW8wrz08jXP/C2hwD4c2ThUpTgMCvDN4/a2LIvv39lhJN6SUMTcfu
nTBPGAWVlwKmh6OmC0P2hCIL6ZoJSRObRATqXoK3iz7Q5Lxs+zAE6/s8kJd59QK6
bP+OoPQdDeCUi/El42/CdAUt3O96t/1hzKq2jk4TVeyLnvV9j5IoErp6NxxX2ndG
j1Nxs2xehrNLAZQVi0a2Z6Z2nt/OHzxXas8DRYqjT4FLQBinJJbx3M8B40zWOc9Q
TsXZMZmTfH3K4OuWXRcBVazXTOhQgAr6rGluAFo0VdiB7JsVGafpfgN5Hz2Wb9AI
/8qqb63jivvbDjTEwYY46AxQncbCh/SdIoyJR+eQjqSIKNK1vKyDPsM0aMe47t9z
0Xwqg/tp6thauWDWGIjTjuPsc5AhuoqMhpY+lJMc/60Ne7u55P5rf+CcN29k4yNa
4gB32xkIrTchnpyBj3C5Fqf/iF6JU1avXw0TP/ME4hePuRRgC7fIIkPRCOINOYV9
ZPpQIo1+7vY8SWfQlTwfTq9hnbYzGKQNxbsut2ox0S7hXIUL3kMr7MF+N4kFOkFG
QI1R/k27EnrAYQ5jzRaE16s/lV9A9Jz18CFt9DW4nnww5KnzXoJE8PyusymR3jml
m6DexXdo4UsVssSyHOdakV5Rg1PMPoaFr7A/K/LGMtCq6EvjOOjOOyTnplqQe4aM
BuqdxaMkboDu6DKvpDjWy2NnUczjjo2CUMm+oxyjCgv6Mmzp9ZWuROsEMUMzTV/D
sfScPQsRaZ44Z40gx88tK9zue2qh7L8wPb/F0E1VKMzSZeGOg95Y6C3W1R0f67Dv
KGoqp4mu2GThF6u701FPclB4fq9pZFLYg3z3BcghGFDR3kE+c8mUEem407tN2ivl
viz2A+iHKa1Zj10A/Zia1H84z1A2zPj/G1FQ20sMSFlVyJh+jdj25ZJPqwF6oOPw
dolLJQtzCxGibu+cyf6lyTDIB03RUwjmthgE7lFMYqGgTbY+I0GV4rrw+d57jSIi
ybiXOYpr5uuowShUMURx5M0uzhS3sq4RsGrrjcP62iOUhPeXkNiqOq21+ynXCqaC
VmY1ijOSncnpZvFin89JNxlBAfo/7elG02NQR9ez0Wf1u8d6aX4AjyE54/tusnV/
HufzZqNUxvauXoSQgZummgC9eDisWUpdzvuaOeYrjGwsALrvEUpBInCRdhwtY7Xk
ZW/H57rrk1Gdt523yX5jeri7OqKNi5VRcWMSPrxEWvLSvzL1Fn4bOyFr3hPXuUck
LLa0cO5Nye6Wfk0fvitWxMIl134b4rwyiWTV+rRhkSsXmkJHpvmXUrc9mWrqCPBY
PD0Hke+fiVDMicxxzCuqvhsE5j/EIhYe0WFMZGyaGzSh/R6rGDFGYlEmhjJX0Ro0
ayl+ch5TcegzBGxW2AfGrGr7lFQpSD7XHFpxTgTxL9XDsmYk0rWzD4X1aWXe+Lk0
ylVdAKsZLIZyHvTL8wyet/R5QlwoOB5cGvQbE/jI4I4Q4+BZa8r2HDOSIy7iW4G6
PATGRmaBu6+d0CtExEMQoa4cHWHTgYNCUitww4ruWt4ghqLrptxGI21eQwMzjVck
5jZ4HskWCnYZQvBYP8VXLGRq2/B/zH+SAp6z6HrSWBEuabnTfho3JaqqdjNpAlwq
ryjCyv4ZzsniWpfFhIWbN41KHAzEeoHhYCZxEfkxx85aCldDjllIzdbdEv6qi7Qz
JopAnuQnV7IWRWg4aD8Wu5k+CUihE4fsGMSg0HLWluFSFpOwdiMK8W93kSN9+3yH
TO0Q8ijE8VHS4ASI8jvQECrLL8QNv+ZzKq8u7xDyFAsiNvEALnHiOSNqrBaqZPOg
LgmttcMy7bvbglZJOQlvHAVD1EkdzfQHayFDHZHl4VR/0hnhatts8QvT8BGGfVId
XKPNAkaIWwc9dCMJDx/7myXm2i4EcL3WHzCZl9wSXMBe9ZymugcGaBr0jJHWY9Wk
9kFWMScHh89chYq8FrsMxEiJxRM8sRRvpmNA4CTHSKf/DkiecxbE7x6KYQIk/TIs
zFDvQ61Cu5s0Mf/C2GpIPlOJQNCpnomNY0rSDqCbM6cGl+rV8MvlZvwGHRFBkfUw
Bz40odB272r+/Qdh6IZ72mblg2ZIs+X4uDQOh1jGm2uVnJ/uc/4LQ0IJHKHpGObr
ei41l3GZbQOAWBoMU+CCAtl/3yUWmawnDol3xv+XPCcmetAjieNsipU7zCNuFD5e
QFd9/1scn/XrsKPsOWPm6zjuxir/ow4t3NtRBji02gQ3kudhpsCW4ivJYbeUnYYC
5xSaATTiH8cUv/f4W7L/XYSvUJ9rYeUtHH1xUKqk2LHgaqfuwDn4di0A98jjbtPF
5Y+gQf3qByPctEfmFMZtQZ9CgFj5HMbIYqMsnJDt2k9LdaWDTNzEDmKnGdRXZbqj
HrC4mDFQVNEq4RViIfqnYXkxSO4eWAR7yzMauHI9Qupn3YyBcfBqacbpHE2petnF
O/sXXThtFCxujwjEyIjY6uJr0hWtr+6J9mwRL2B1VWLsUrezRevXK58egN1lFN13
i1WAg6FHauQr+ULWlEdrxrfiSBx59FIhiY5e73OhRl8ErK21PXyaMYFmtljNJJKI
9CM9tPmJm1vO4lG6snVvxpPIhxxS8kKBoghcpdKSvpBexcEY9mLKM9Ah03Yy3qpC
9taby5kbVu0QpSt79W7YRDT1sxWKNcTIyHrIQ9ktilZzSV/LAqlPef9y5mpQxomA
i6DkRG5Yz//VsibPodFjXQbw9KSsOtHu6PGzqIYT/7FF3AbXr9t868aHhMwBJ4in
i1hSkZ3ndGFtziDzz007jKLt/r4jCfuWF7eI0WqkkRY8sQkC1JnMTZfjoKggdUnr
n3soxV+gMwyO4NqNP1hOS4UP3wbgAiu+rFCbjDPbuEwY/eTK6fndF0/eqllIg/TC
4gS+ZqXDEY1QDeJZ1ADdr9VQCiPcpWthg91It+iiKIMBucnJqQV0C3RVr1uRLe1T
/31S4Jka8kFMsQcZaNQzWrrYbqfip/OpqqJigHnn08Oia+R0Mi096JHudeYnQ7yT
QZRbTYv3jSi2QzmTevEQP7Ex+v92PGMKQBFvubsgeLpekYfLnz7zyfVmvLzft/HA
PNXIekBvGrnjy9jrcfF4f+Z2l01eLwy8E6XUrpGublmQuom2b73sgMs5eZuGdY0b
mRyDtKlKgWnpIopudnVDaOnpvxG/4J+MhRJygnRBIzM1TheAGvd+Ahaq3DnYP5n9
SkGOJ5NFL/fhy8MUYe9+NA4sutLLGVa2UoWa2ScNSrNkKzSfZ+N4G+sZYevmP71Z
gaPzLKDbSZBXD9Qnj7+3frpVIkcupFA/te8NCWFTz+15PZERcvdMHqMpuPq+QBM3
3EUHM0THyZL/9IsiQN+wkyXv3+16rrkX656TVS30ipxI2BDDIHYCpX0XTthCRBrb
qbsQDw+Jzwbjm1QX5OyHnkuMpWHfTGrex3uDLNCXK7VVCjph9XjHtbgZRHlvVs5H
MjSZlucvKZtnE1KqLnDGE1vX6Q7v+a+lWNMvejefy9tEzhC4AwBTL2er3SbN2pCD
PfGCDXaBL6m2hFzxAHfot80qNV7j7BLzU8vHuqH8hQc49OddVNlOgITn0RO0ZUXm
7pfXcc0etfe47FkflbGHAZvLquaWAmQ+EQVN1GBfU8s5fVu55VWkpa4OUDaNbBXm
zoOKkUfyB2JJ52ImPPFgZ5APtTiz+7FKBIFdWgOn4eULju+wSpRAdeOn4/MmpkTh
CE6FYdnX9BCUgVRiT7B4yzUjrQSuNKoAXJUZ0Qrt7a1e2S/2N3XVz6k6ebjnlv5e
hvOtgKvi84r14O3f62W0YBO5Aqd+HPZmJTN9PBJhhmK0DNhKjq8Qy4Hkk3yvHWLM
927OxmvOktezmdzFseyNwcMMS9GmuN7uKYZSWet0wiunW6GKo8Wgv/dZNVoXdt6v
4maoMhZ9TViaesMGLfT00lauV82T5cIHJXbcjQh33qn7/FNrapy1RSTwC4gROUS2
79+xN1437IssYNRNPKtXUd8gzTmrZ1c/RVbfUxCvuEy8zBgEH/Wy58+cgGrNoXHd
1twxWgmj04Tgu0ChOSWQYB2t3XToEOor6LoSUx9UepdeLLKcdseiSxNFBYwuN0Kz
Aqn1asijrgczH3QY3sBNAmuii3a18ZTZeMkg/YwkSwQZGNGzy3uu0qfkVaY+hYqc
2UKv6jSzExh56xPBuwXpuvV2FbQ4DBg4T7+LIwV5X2uw4pvGf/ngGfSTsfJLFD5Y
EZeHb2buA2aMPxojD1SunrSr7juPHyKPM1edPHCCIk7O8xtvmRwxd1XvfZWA/rla
vyNEqm4h5ClZGVXqdsRK6B9In1ApHWJOVA8bYchVUqp+LmJ8h7YEK5D02PxZQr3X
/G6CaY08vTqEj+i5NCvCQEjWUgj4Oi2PKDmTjhORabMdLFrTOvCCldj8ORu1zcAI
qto/QyCFJSoNHMTxercNCuddoYoh7htvNjfNwEo/rzEHDYuJ3hOJ33tjp8GadU2v
EAwuTVZyDonAbjB6VpygmxL/KhUIji4NArppfq/1U+RiR6w6PbtWFgrgHxgusJrk
0D1ZeALiHRvz4dmNjdPLp1wLeBI+0DOxwTNwWt/t/LzTNXo0nM3xmAj4846jOAK6
+p0Sth9sxsVdzynke3WeomvLnyvkHwDQPPqMX/2PYxOBrliVr3BJeftpwZrqZsIW
xErUC3zm2ph36ewQriQsJ7eAy1Nh5CSrWSu/mcLBCQcR1VSg7adGyVRNBrDBIXci
8tTtA6JXy1TINDaSbSeVpRUT89RWPbghs42XwziIyaMO5rw+Yy5ukJek6fJK+yqu
Amixk6syZvAxb2Rk6LSycDXd85Gr4q5ZEiWQ6TtwJ2JUw/SVnuK9YX232yxHnI3C
PAe3tIkulvvFurI3nVyyzU6CqwQvoxmq1emXCk2FGK12NrfY0ZBa9I0T2brgs/93
XPDS5UYkRa6WygGGLNe2DDvGg0px0qwCYWNfP3PWBcgIsLIeWecw2Xh6Vxx4gRlp
URGcOKFHeZTExt07NCq4PkDQvyTBMMwNhqGQx30xUom2l4z2oMuQZxm3UPGxt8ku
06NBmUO/2k/p8xBA4niT+Pci2gW7SFZMAIhT/eaNW7xO7RbDJ4Es8w9gYMEiixXn
Qmwj2dbHXXm7P+/FWa+PqCg6eE3caO1bat975kFmLExrbwYX4WdkGltwcwCAS2WS
QrUtmZJ10ZeKuucD7ky7Qmhwe9DX0UaRpELWKuij02sPpYD1HE5ODczUXbsLLVFN
zNDSj764PL2xb4E07h8R58vDkR33Ld1WVfL9uXw1c00pY/RMeEkknWl9qJ6XFYqK
d+KP0kwPFuJVv+ECKQuc1A73PlhwlOuuZ9F+kBFvP46QhFtgRcOUcoua7hl9NOiD
XbNNp8ZS79IpSLafRBpFL79igUXE1YLB3rYRVJ56us+s8jEppGvKbMm9JMuVyG29
z1LjVDi/Nao2jEoHaQwUJaUQolIkDsDPt8xNHmYX9kMPZMrlbicFzSLQ2GNBDTnn
MnUb9mZ9agEtaB9nC2ahFvdYgHTIWRwMZCPAbomKxjhe4rvyA1Z6KWJnhwj3ovdl
2ouKzPIM/gpptVZUgToIRTSZVn5uELmea1Sn8ehLD2rmbyASs980bjJWifUr2rZc
mRfEJ9eW72rIHjIJDHZTZkigrnlRhSXpZC83k32ssnu1nhjRKYFX3YNaCGGnjZTb
nkPFbobzie0DROdxzAfsvSPG/TLN6WqvDPOLFeH2GB1XAx9DJeZneGf/Gpdpz/qG
0sl3qAL9Mhc6cd4bAjRGPEzQ2kyAckdfdzXyinyDNgfiGTej83t6r9/tQLkMhN1y
ImCwyXmQ4kvyL6itTmed4sqv4ctFLYOMsAMo9fcFE0MwCNvkdcXjkvSmQwgWXK5r
b2lNHAywX70eJCcPNSyBmo7O8dlO7zURd5VGc0E7iK5gBM8Y/1ZdzYvAkczR85lw
PJ8TkGHEk5BhQpNmUpMN0mLXByvnSZuGOodv4/8jyOhUgei+99U7fBUxerQd8rkH
k91kWxBH+B1Vr8Buvjmddla59+iVE2NjiiydAM8mAWcvf/Q6hhQzDlSNV4et6MsB
/2pG4MWDbHcLnweawfcikzooMqUXM2X6CpzoMavrikr2OBJB7a+lBFp4QWNH2c0S
SSyXXNychsvVue8RFo9VlG3cPuy+DJ7vDAGOh2AbbCXq5z7u4vsR1FohhaZjVnVW
hqtn7h3luTeYc/S08a8LlKg5z/hy/czqRyIui3F50L9OBEuDhjFH+cgz3xLetq9I
kBJQl/xND6FAhu+Uh1GMfIW7G6bkCmcj0SOfDSKYyl+NKmLO8tOWo0O81iWeyzx1
eOth6nSLqsyQyU8Jlq81ihNI0cTRMJEfNrd3VfXvh4P68BygcZSsrhlGSuh0ZBUF
PNh25yseBnFsFbXozRZnyGTOInOJcKvo/D63KuHPFz0/7fP1Vd7Gp7aTt7KXas8A
7o1nkGPk2xkc6RYY6XeZGUtzW6a4FYzxp2MwP62xxyW7gAUfDc4IwXCgyoiNTeL6
6BIyh9U1efMS2hBrgkitO37tLRwbj0THXS9Bs2Kh/FB+VQ6SWR2i1BcLFVuf0/6Z
fU7vyChXxWEd4sKlqVtqdQ8h5A/eZ60hIz6xIHHJ9Ngpicf5foCFRWN8BR9JeFpN
c1RFBIXaRB4siar5HfzQM0EzdjjOXzi/xBLlYt1Zis7b3qnPkvCxns37O7Jw19aM
0C+VdTcc+c6PmGTqIfNNAjswpQdRTaF0/i0GfodMaIN8av72Ke4CiEaw1Z3acbRp
Rs80/KJV1n44Umj20FYMvirYKB+MQik8I+eImF341jbcNhFxBByAPng2WpYdsaVs
xsBuS7pCJyiCyNYxIYEWGikKIR8c8sEMDS1aP0eiEe66d0w5wPBEpzUXHnYhU3BH
VZyC4BAn6vLjJwdvJ6H3keov9vwnVT1gVY0CQBRNHsN5p3MiG78V/dg6T2u76BXi
HXLV/Tu31bsiA9rstyJNwhNMUHc4wh97h91dy/teIRKw8y+CQVIVfLaGcxrWWbyX
6v9uTNxZdXN/01JmRvIBn+ChNVJIjs1Zisq3UVQfJTTEAIcpQ+IDLeGaNxy/wFeZ
Yuv/vlB+ikU394C0btlhwYWXH023cB2BR5vetUjf02ddWF+Whpl+Plajknn2xlo+
Kq+uOzuGjDuvw/F1a/VSUjuJ+Hwdh+yX4tz4JOaTkEqwmxJx9V818jduGjzHCFov
F2bbtkJSoqjril+yfrW13S9AA02T8GE+qt9WVso8tiGn6FM9lLm1LjkygJqizh55
IT3xF3dQPwFucRh7w0y70zCC7CQ4bKktICqniaVJwdTQE6MF35XyIn/TOh/wTMi3
87uMsj+nji/p4/fdnRApnJsKKTFdYS5XZZt6ZfFnf2E8MKge1R5B4A7QO5Am3kKF
Es9tew5zrmXEd/uvWLnfuAAFaCe7RqseBUMlmy56GAQBXC1+kMwltbJhW1yWZN/k
2bKHIWkJZLZXWIkWaURBZeU+mMKjsutTQfjBRagtnSBh3P/dTcOczv9wjKPqo0nZ
kkEVk7phfjKbVJggehnSmAxxrsaNAAkp5exnirg9T3p1yqQ/zEJcgIHt5RkEzAbP
fzi1oLk6zZ6LUD4hAPoE/9XwKk5sWWy5u9vtOfmRl/2bo2VOlhKWDQkp3nrqVkau
CXz0oPpmUoEGk+Slg/RjVT11qPgjIa/wu3XNxijq5sEYOolUyBYz5bS+bmW0iPDT
hn2ZO6W6+WW7SxpZW7W7pQX96APNijN0ttEFN0ljM8gaPryqbww7kBC9XAa/DODw
cOk4/EAzrIEzwofoV1JDWpCoAmXeE+DRYNq6cypNtnbGWzWtlmnlV+URGGNh0TmJ
VHRhe/nbuKedwpT5Q7cTb4n7PbDmYkIP/Rj0lYCMVNI8rC0hV8JzlXzEaXYRUnAD
BOzYmY9eELRctaF7O38gnc289sZMtsWoL1OCJFW7ZNt9kA75JQOqpzi0wCFZzyQ+
ewhF9jfovkSHDS4cFw3NFgfaUxziSA4MAalDj3UrtSKjv3LaQbyFERdz47vsRpV0
UOQPMJ6z2UppWWerEn/XjgMUg+UeZPrefdNP5c0RHdNlb8igGSszdveVXmkarcoY
l9AEFYwn9MvxAWl51tas7H/UnBqNZs3+qHcuC0h+MMS7n7riXMDMX1ttsnG/s5Mt
ahXZHlvkwl5ooxOE1HhpmT+QB7l8j1apG/RqUYxJ3hRzidyPwpWSNCudqHSsCY83
rHv6GNTpAXelRJKc8iLFQm+KX5Ti6s5dl5mXQPxoMBrye0jeKHkSi2ksOd36JNJg
mcOQcjtls5uyGfMUk5pEBhXWnQowXI29zEkHfHr2db/KfgYpKt1quaerjQnsjZ0F
UYb9mppK0ZYZi7ZRbo7TGyq/gMud3cPOW3F0xnyfIKfxjP39uGBgot6ebA8Wgq3l
vpdW3SIC0FYUkclME9aQ/7H5w0npdvB6iNlfPLg6llQqBkq00GeSrlq18eHwg+k/
AH0WXElNkhFcIPZqHDC0eBxm66dX//4m4ixEKr5032CCGNcjWKcAc3o+u5lRuB9v
yedGkLKAU++uBuEu+9MSESR3dkF0zWXuPCO1i09FJ3hTuQwnSibvhqwBuPZ2sZ5C
DGhNwlJFDH/SFWnYF1EfizGzOYXEF2v81QnDHU2Ksnkh0NzSZKLQyXOsAwNeMEMx
Xx4yuXF9gKfJS9icYA+ShMu9DxBbiEA77vv2CWUX1lCV+2xevkfqxOS9M9b9kwDm
+2AQZNatBag75WhVjjWN819kepWCSvqSmr4twLKMU0VqJ6jW5MwtSP77vagp/RwV
JiqgV58slYhy6jY3qn57ZYfRWsmS8X6SOnOF7offj4G/TXZBI93mB6s96IApDrDP
CKy7XSwkul/cnWb2N68RO02yvdLQhHKGoQkTQiHf8PRepehg8ahk+XGLpzLk3+lL
moEsDT2+TSCaeO0ovJZ04iu1bzYwEjdUrk2NhSYvxrfYSpD2Eu06xkx3GdFo8hnM
eyh/bfy+Qh0R6jDP4xn4UJRkMFez1pHYOfQpDDG32hUtqsQdR4InfiKq9Ip4TwCl
4ch+RPTXwSHxczRvf1v0zVYwx8mf+KSFo+A3QchVHu0wBaplAL003KPrYCZShrbY
+jYR3+CE5m1FRcejbj2g4qbeH0PzeRWRS0f3UziObUOf4OfNOBIVvbRgALQepldb
FoSOduRJH+jgcj68xmrpubk6ssTtiLZRi++wmWJjKTSjg7FSLOfUYNPmE03mrwU0
sKMbP56RebKaNgoXWN6mRfET2MCZ6XvRdHc/6nJ5zuQDDEM3je0PFSMiIwo8o+Gs
MZrvE40SI5M3qUSQnLmsHT4GlTEovZGx7p53KnPXrYArM9a1+OaaWGptggcIC3l/
MjunB4cgCzwkhrmknMVC79CZk8d1vAeINChefLLJ5MuHH05gBYWPQE7b6ywuzlPK
rBkoY+wYTY3awcH1f7BVLUb3YLDCgw+XHCLmwMfCER70filtEXyT7rFN/+dOcILA
bLIgxKuFZhmtqGU4WHXQorhjRilOxT+RR06MgZL0MHKwYRDDwbsDYxcGSfOQjwSf
1bhVvtEEvL2hLKXenAHf1SAYL6Om+PH1nMVV//ki40gI0UD41k/JpzUetMtZyyF1
GpK05dpdzDs4WnWHV4t7+k+cLWNf9jtHi72gCgYd+165PkQR2ciiEFcG9OTKTknO
vfrps/p3IY5IvIWpeq9hcT27TNhJqgjRKis1Jw97GLC9gJhW6t/kXT3Wf01LhL3X
AoIE3HYhKOojRRTbPZM7G3c1hNTsd3cqzRaUey44jSWcgdgYoYP0C9D3nEw2SUCV
nZO4/0w07KrChd7GEnewIIQukAercxCqyLbg2DYkeKLSGsRzTEyUqQfzEFe4/X7x
9UFC7O3ZXWpFh2ZtuiWz64W87ScCWsC4bafSNFNATHxCZ2cBUVL5lKy/9KnjAVwU
fEHZB/dP2mTl3DoBurNgazwgH+LJDjAh3Q6jY/XW2D1GHvtjiM84e0NLVXkA0bf7
zk56xisq9a3VwR1sTaL2OQ5HsuGfF3xJJtwWnHs6GnSPPHt3AH+q3+r6CDrsUZED
ayHFgQc7u2cwwqljlIjlAcr+yQI0OGIgQ/sXuxMD2Lr1vtU6JNc1EqiZHQEvxw74
CmeQnKoFZNdSHmBrB5UPN9Eay6nNg8uV4bvfoImdkNrUGqjyId8HFKalEzRzOcFl
xiD5NrdRRo8A/bgZExTn/jc8EIN3KNYhSG2OUxIe8fA6Vn9vgX2rpVsF+LQbHqAE
ka/MIZADz2yNQEgC39Rabn9Qz5K1Z70PGDM7rRgQNyGHibw+YmeUEN1m3EAEnc+w
tuj1JLGnduO8zZJSUm3fEkCQN3PIkTa2x2LNWur3sgHlbskfcKerxh+QNimUm0Io
dnddRhOn0fDaLwyg39mdnRzVBgVBZ8+GfZWejvGki2P6h7ZT8FuOSEkm3JC2YpF1
FQb4buU/IAmNwPT4kJDdOtVVjLxjKqLdoc9e4YyStjLFzwSFiNQS3vuSZbTYzeMs
L7ep+gxLLW9SgdJVbXksYSb8zdhdMEWIMiXqQqXrMS/p5jiRO5/ea1BN1CRY3Ql0
Fzvl+1BATiMzNH7+o8lVYKGKFP8NVARsi+lpSJkJRnID0ouNp48OfV4mXdczL6cq
gK0ht2dSQFCLBKJiU5/OKKSPNBQeJXgeCSd4PooowPtWZZb5arj2Z/eyBnK9CTKw
aCual8ZDoRPoWaFn5tpFCwMokVABE0WFZ4QlJ/BZtZ5Aqo1ljSecxlsjVeaGuMiS
F/BgNE0mK4ZKk7oJaY8fv3GGU692fFhAk+nsEdGFxCCKGpWm8jaVYDCTMMgjz3J3
msd+dmWfAqG2AuX5+lZFy8nuhA/8rHnhyVb1GwfUQiGxIlcQEHiyXrb6ouff9nnI
quwHokh7vaBjH8cPRfzM7o8sRWEMiXiMmbEi1RuGy0BaPgU21XMFiJjLufXaOXRp
kLHrY5BAz5S0cIsWZTqI2bUC1EaK5w+f+SL3khgMVpM7xbUxAvT+14E3etNApdGG
gy4tgzz+kB8YY0N7ykjIn8jTlOjRjA1ak6aMLLuq1REucmyeNU6FDbblMeRSi47a
wtWF+RuLnncIL/+EDqtTYbhOrCEAtpLNDvW2GdgeS9H2Bde9uipUFOFxI+4lfhZE
B7ogLiqAe2sG5of3oQraEBNi/wzCIzltc3fFlde2AA9e1moaCf6jEkCPTO6Kvohe
QqxhH4tblRyMKRRt0QZzOrA5LAyI34epKDizH34SSRFq9wJjzK72L6BSil4W87mO
Ny7Vxpv0BJMrhAudvVaUuyLwXeuWhM0lLCcmoVUqkMKPVj0xoSebLCJpQJ5A5W0c
8uCxkNlVGqEai4A4RdgDmu1kvmd+CmwNcI13JdbsnYbkCUeINudEeWnq7NTOC9sv
xm77PVPJPrt7hKSFCeiXDypHkaaq8oOtoJfyB42ZmjElYUcV63J3EupC92Losc6M
I0WS4TFxVYUtYlqS7JsIo4G6UGScPpuKIN1pErU8QcZnjwvXfgGOYemdSJf7TNsq
WR4d51C9j4g4ytwsyLJI44xwBWo4zA7uw9QHrrNiAYC0p9N7hvKbvU6LMUfMFYQW
TZ4pMJwUaBCvNnbkN3vphQ8tDWSBjHWfu9A8JHk7ebZocNFRFPHXvNJjmYO8DsFt
WfflJi3fK/nzjnfavE/kADuegx8umvX7GcI1IqSG91pYIYsOYiiz6wl2KOyrCyMW
+W29Z4wxh0BVdEdXeBqA6W9B39gUiZj+DrvLsD/Ub2PL5aNeLhfE6gtlLLxl0UFq
1AvAER+NLd94iP22JEu+fsINaupoAGdXVLjAEmMg7eqXFwZ3NgaVHDNIZJWriKEK
PQ7nJ0b4Z8POq/rqNpYqd5ZSnxxkZdaFj2h2/4f+OGtXrC7iLnx1RP/4Tn0c1TY6
VoTIWTuqeKekHZBemMT4RpeqaOXSTEXl8svh+yMU8QcF65DhteNLtNLm/Axl4npg
cCPEG8S+xYBEeT+PPEdsNT3vazUDyKlwbw0A5FG4UgyjqV9csT4dWaGG5+N/F44+
svTBFZxU2fTWxbIQaI/Jm1+3/J+JwCGJ7PkQP5ESh183z8/zP/kKsj7Zp8j4BNPm
Cc3DQBJf7xE99uVoSXYEqXjc66+Zckhy9/3ApGLeBykY1VinjI+sdTu2ZCzfb25t
4MQX14gFHZzhAHHX0FTRGqDM7PRPfLSpGYDD+yjdKAex4V4MPSa+vwVMn/hQM4vv
OcGu1KSE59/Im0EXeqi5jveEAaK0QO8ASrMRWTBUy7LP5yhJiI7sFdFphee2st/t
+t4RXxErImnhY4CnejYvbHhrwyOvDldX0jiWGicaaVwEhDm9rXFWDSnD/1xRpR3Q
6+5w54HP0tXGrzKILBzqX/w/sfSP+mJzedWjxcXsDK0xfa3Zk1XBSGOQc3IvhvmG
b5VCChQk3OyFkKSF0Hs2NvUD4vuckOd9PIrMXt2XepENY/2iYpPrXtqMi/vT//mu
3j/mINChqExcxQz6si1PN+jjWyqoHcSj/xjtYIESDNsadOkJfNwy1c1QRxplGfB9
SU5qEv53naxrI7GTkcSnL5wJyA/pk3AJ/CulpvBYi8kZku75y9im4+RTkWikKRpg
ykyV/4MRqrl9xu1ID6rF42X7uvY389LFKzUvLEZdvQHnYxDpi7yEsqs14O4wj+yZ
YzdjjBPlN/Ut5TaAuc90ATS/xbXiq92bTlASP8/BS7d15Rs/iDZ693Tm2du7eqOg
CdM5TyTrF87EfZYI952A+8JZoWDQEpmMrgzEgkU6EDfWbOpBZR+kciI+jG49NLXt
6prpIhnSWujfot2nOhmBCfx/v/z8Xowt6m5qufL9Aulpaf+5I7j9kHmpYkuV8zGu
aSfadjkw+ionjea65JjYoSonoDV0WSg/PdA0unjv+EYFPAXaUh39bns2zKG7iW82
66D0lW1LnEiv2JU0r+fgyKOaMAyAiT1qzFioqKv319iNKD0fWHeNH12dFW/BU9kT
hSEJ6HyIDFBGB2D6OBtewx71lE1V0EcJjaLuhSuTbUnZ4643vVdPtZPFxDxj4xC1
+ec6hSyUIMGJXwGRNYCbdxXErcNZbul2f0X25flGrOCCKZspjw+M/3q1R+BxYJ8L
VMeqa2+TvPObmJCQeEYu5H0Hc+YojfphuMltUqKe2PTJm1BoHjx1jY4RaBJzsWdh
t6EGVYUo+xloFi8LRSFG9SONv8TXIgk9+RFfaxORvkryDr9fWzs8VSr77S81GKjW
AHUiWLKlHg0DYeC1pcltPhL7bxwjbIG7/gyQ55HzoJIqLVvor+9zFvTP95iGIKbw
YBQlC0dVEM0hMyuJmpzOAN3LN7rtjJECX9kxNzE/FNi/wwGADHF8hxwj+z7QMxF3
GkYhCIoCND4mwr6vhcwVNh7LyOwf7dtgq8366jr/zNkio1v3tnHxw5NUVzLNbgPT
5z8enCrdf5IwZRxY12SEvOh1UwNQvFqUTp6idhSPQhvcpFDVIBkZ4sMRwKAAMWit
ct7xTooIDGLOrgH34XF94FznhecpwqbVCdM5mc4oS+tYrviDOGoybOQHI8eDcdBb
NZNNukQiYW385WqE4yoewgtif0Nxa7zhn6xXmrTE1qZ3U1/roowWYMCVWe0G4SEo
DZ9w8uIM3uPmT2HdSR0qRTZKH/laK65rUbx0O2cI1VFFWqns7SQD27R8Ds3FiIDl
SealkvXGz1b53O7Zz4Z0wEcjsfvIB5P5No/LQHMFNjTKpMtqIef+0uvHvhdX4WaH
5IpLeqYiEXzYBfJ/QbX4B12LD1dATwvRUB+0mle5yWd/aTYbqh0bfFiJMtZulWiZ
+j/d0J1Q1nayqGGEkKDlJYSVUkqxkuBx2Ata2OUWGltx+cdF0nsAKzETP2ofE/Qx
JDatGahf0g81W+QS77271b3DMcVWN3VYKu36RVE7TduuFj3NMGV3qLC7QJC7Mi1I
bxcudL7UtxhpiBV1RkWCqVFZHg/U0/N/CPD5ER/gGZkG6GegPDdzHykKGAtUdVvG
w1QESA0YsjdpgGKprIKUgvG/215AwSr+Oe4//C2atsJLyYG/nDEDNs4rj6/KIJWV
YOdFoMeliTAOWoR1W2jcuSRDbzWElBO/S3cAlac0vRpVhcdyWdsoX5QLGxInMLQa
b37VvVh7XLxFAhbvMrXV30CNZ4DFsRn7Xv2heoPV3/HI5UntdDdagyEtLBo+Hwy6
2vX2dJEdETnl0GUSM3pgtlwv/IelnJ08DAY4uBDGnlB4An8kc03TFcjWv0CCf6mZ
bylt6T8YHHDjW9Lbib7PNWXBqz+yoibPuPdbwDxB/dxoAW5gsYGks0Je8jHwib9d
+C2hKhilh7J7jvqhC9XYfpzXneyGTH84N4a8g1KTqLttU24Kvw6uwjOsFmmigg4D
tUQpIMfKmLzLcpn+C41wCZ0xlw1WtaE171fADayASJMgnkST9O7Up7+6f5HIIjeD
DwZ/GKsEXCUxMceY4mQBa1+1GgX4ZVYPq/G/6QZ8dhFMMhCRKUCFEYVWAPyo1FiZ
XaNIfXlCqArrtIWprlXbfxGK4JndROaus8elp9QDyOR+jDYG16lZDRc/i0bj6oEO
8rPehxt9XXNSLWJkFF/y4Hb+ynA4qO7g5SAHzgkhCEQCFjT8bSra7uGzNCBq7f6P
F4xrefxhjqLG6N4i/HgA1FdruKsXSPqJJeNoCF2REgiZVSPkj3gC5c1hMBzK56+W
SpylyaSs0fEM0N+/AM9igdDqWtSEzlmb/YQuw9oKUmaw6kntCqy3ss3kSX2PPk0R
HCBwprWeymDcusDuyasoK2dgb6bJX/bJxH6SfdB6ZZS2qiYxud7adyqsQ0Pa2doj
i0e0A8sJt1f6oyxI/K5Viu+QLn6mPNytwIH5G12F0BEgMKnzvoi3nV0x9nanGlA2
Y8KlOxQeXdG6i6trS4j5kSdx8bv5IKWA0jCnXu55ekckYQ2gH672+TpghWFE4CgW
lT1KiDXFKL73tJatn+EWVdCj/joKMYH/DnTbHzuO98byc8KNiEewlEfc9ry0gABS
2GC+CsonIrIGV2dDFXyHeM+J2DVuD36kQYp7oq/PSsKDA3OoWIqVR7ZkLvmmpGSj
D4HWjp05GkLdrM47kV0zdEOi3SIQWNq8wurrATt3hW2A1vveyGdpbg1RJQeJ6kni
HSBgqTyPlJcSLsTgw0JMkQ8Qu0lOMpeXeWI4I8mXl49shdLubuxUkCE0j4oP6Feq
n2VH3VYMjcrXxokhEO3OMxa9gDZCnBlDnw6frb36uZnElOG762mfjMmOJLnmu8l7
8zjc1regp2ONiXUgnNYP+2jIah3fZQh0bIdb//5OP3kIFO5WOjy63PUkSz6zkh3Z
lJmSh0fQA9QHDlUQSkiFQSJ5jd5RoE3tLUFsSwRYuO8yWh735LF94RkkI3GE/N/H
lqNP/PHlnY/6TpDMRjSCPz3nIK/UW9CD28xoeW7WrivFdOIu2cwsfLogOwHsgySy
m5C2lPQ1PLFbikqRHm3Pn6auGX1QIdRZ1Zn9JAcGI4AOBkPg5HNZv//1Gb3K7IAY
hD2Rv8aMeZa9RDru/kMbJlXz3CrKvpeHll1c0RcHZA695gLepifcVrKRa80o8xc7
DQKqxdV+ZyK2cDO8QZc14bVphuUFxFzhDYm2oHxNq8+2Orp8Otiy+88/9/kXNRir
6lWwZBKDb5Hhjns0UQa5aEUvXF1apmkMQHXoFnKIlRRDzD1RxtD1SIGfZEcN/YsJ
Ci+kdt6/HUGh1OScSBORq2IGL7isNqrEdG1kYJmxQD5s4EjjNRyxTw9JFk/er4Gq
XVvN+6onymQBR9s1aLOYofz9nqFGB0ZlogQxvvbKc3yMICMbrQyD3OcvZvv23o7Y
XPRmyz0cnzUz+95HURgHTgDsSLl9aa4Mw+zSXIgC6egboBc3UJ4GloMxcPPe/SKZ
JkY6RmaxPitXwLgP8XL3cU2I4UNqJ8zFrzfZSwEmEqILb2+KVch7pfXTlw5Cr/MT
JWRiG8yVPQCLsACnvXNuVXujILzGMzAkYG/NhVfq7XALVoxWD9ytBa6aSLM3GXLr
tUkoz6XtiRB8i+Sip9aU9k/Q67UshXF5fjSLZqCqy7QtQ/Ys3/xPxTfqjQxoquBW
/ST+2EAiMvBGz9PRD1tL067L1pXcY2l2vw/Qx8Nf9LzgwYSbFzeoho4AxJZoGMyQ
g+fU2aHlsCp6AWCRKxW5GCX5R13hAE9uLgtIx+O2v2dFuNLo+LLr1fJqUxR5Q4Ef
e5VnFjakgayhDZMWyuNHEEFLT5k5k9huRSb2on+2SU/L82h1ahTeMUllVuMBwQtG
ae/juBHfi1ek7BMilVAk4lYQhgx3cL+4AuMpkTs+iLR1NaKvdhsxBALCu5YyF1aV
jAN2Wz4AEu5J3nQO3SPG12/Psp9pL8AcCY++J2+Zcq5t0kJUdIWfJyeuI+tYbeKz
mfnI03TGPg3ZIOLqHuUEEHPPHI0qZiMmmkArO41AYmoV2D7oUJNtLskfYdB/Nddg
PSdSaMkyBKnvWx2q5RbJlHIBBSNBff1jxcn16D+Q9NQoh8MxvrcIwcyF6/y5unwP
5hQNtvRJXMdBPqjc1E7SHezMB/l3kVa/bwi4z6BLSa7RcWymnqN8DUo5Nfeac2QT
z05RSBlJyruKeWBJpWJi7+Id5GyIlKsCm7qowEGk4pTmBEXuFvW6CerEKz0F+yDR
oKrdrjaWzzZI/CCRrOFfMly+PQdZi7KY2AMbLkItVZQw/9lGz9yyw/Go/V8BfCkY
vSDjJvHvkTSnT/Mis8vAyLDtOZk40M/T8njjRfkE4qPWhRWQ6dCf5ECAzWbG9qun
6vbrJI1b4y0w///A6bWquZzueGCN5ZnCCAVcPrvTGqBYV70zRWC2/paWx8MbaiIc
E45j08XnGDDC8o3DZVHeXW3fUaRQ9ITIevEwD2vsgwX1n7yWCjXxFnskt/1pcANn
fbTVI7SRplROp2Xlsqijz/ZpKclb1kx5/ebefBm6F+5osTQ7D0wlhbClq8FnSibN
C8+5qRuJLlUsyaeAYu3nZSz/kcBwvNrykVcCBuId68qHt0U2Pa03mDWy7koJR2Ba
HU3SQ7dJ4fefNd1p1YtKwgOw5j4sVUBInjh49nzONhXQMFJfj28ku5r9mjX2XaAN
ZvhoBWUCkhggIJUa/azL0MD+n/fSilSDiGXGpuOyyQYw6BiIsB8MyTPqJTbogWBz
+X77uCikqjemF3P8cQhQI5XEVPm5ySmg3m62ASP1GdRPZ6HZqFEZuK33Rwexwm3B
+sgDRxOd4fZ3HUmwwTWwy9VazGf/B1MReDGxilOBdzz/nEbmWvzxZeJ4jZW2nu/1
ObH3jrPdbNY5GIAWT7l70mQOaQKQWaDsecGPJIpVox7wr8nPuGjOW0Ue0PZYmxEy
1RRN7ntq9Gl2F6qBcnTQcbh2hKhEUwKbrCyjpmDFJGZSnR1AvhNYgTIlEvWpukaO
JQLvSSi1ffveHBGXB/hv9fGmutAKXj111HRld5KypVc8p6fCH/2Z4pPNWannzknI
mCl+2RrQUE5TwbeCQfBIKhgUfvP30SwOMhEM4wFnyBjL5VSZWsQVK01vGd68IOMA
Ab6ra1FMLGAmz4b/96EkV21VpFK3sCmMcFm+3hYV0zxXN4sqBP+4AeHprNB7spAI
fvf+vzdmE2BRf21dKmRBbQdXYpuAKFA3Vu1PMqJGB9/vxOOVLfYEvuM1Ux0roEHj
YhlKge4dFAxQTgUQ3FjnJC4/OdY2iaUSDpecH4S/iFzVjJGxpAw9vWxVmj/HfK4Y
J3eJ0d8291Fp7L1aQpiMEZE4Gl2cJ0MfEO+Z7b2XR4rRy3Vppj8sUjWPuF9wbgx8
PpY7+/sno2vkmVe34CViZe3qRuVTdBBgc9hfEqVQJsCSY8f9iBZp1Zl4r2FXjEvS
ibEjigGWUAX1qCXBiWVfRj7VJefKj/39FNFNhi6IgYSrQE3134+j/qa5PW+2i1Dd
wZ7eLrA3CWBtFH6LGOfxeWlpbtaYNX2PtoahHaXE4VSZWNAOwIyl6r1lmQbjkeyT
aKPLg+YyJNXWm1O/fO4E3h+EZ+L36QMvhMDAIQDhD2tJaOi1a5YD+B/noeBceCxK
Pm8/m7z35UxuIA+vDjtnGT80OY9nXlkBrbbcbRw/UO/YBYl2Z5MaEmEpf7r+fnGH
qwyRVgYn34GbfO27c7iwKtUjVOHgwCsBk59HX8y9jGAPbs787kSg5D40CFfWlfHT
bTBYg0vtxDQPGrmcfj4GV+UqpD447zzOuR409bqu7FUPmOGRJqXNd82NIch+HYkR
cwXIdvL8Cn90r5Y0pe4Y7FmOT57HF1i6x5xQucxYFPDU2PYnUKA9wVweAeqlbSp9
kWeZzkeZcXoCHs0Cv5sFliiZEv+vIt9WeUhM2QKbCtHFCH01TdQAlH0btnxQug6M
fMFDLKJiciLPij64Ti0g1BKTGCak6B9+SSs45S0NOn+ox4dessNvTzfzoAjpTESp
J78gniJzm4lZ1d5s8QJouDoYD+mZ8EYsIgxPb9Bl5vhTstiqygLV8dlDJ1YMIRYG
PwhXooBUNqejxUFSJ7meqaRLb5yPElZkjpuIq18Dr+IwAqETppDdSt3GfuHZ5DXF
4vJ6ugNHtF+aegmdDzdTwgFG/jU/dVfcXft4eTqwvMx/Lvx/jQPfySqHr/7hGj1E
nnICwJMAQDAMntJGwH3YZxF2GQRyhf3NKygYJ+od+Kst7BTdkZq/850VdjrqMn2Z
uJ4MsZhVulB97owNK2YTnh72UNKxysndYFr+6SqP7lk040dFTLPd2inYQhXRsbA0
I/h1wzR/lwWTOyVKD3ViRNNZ4hOGTwPKBtyn42wok66jFVVpSGEDolYg28priGeL
SFxl8jvt4tO8u2tGj2py37NWm+xPUXIq4Yxjl7LGzpoiSM+l2xP98j/4RxknrITa
O/5zmddRxSM/TTsXPl8U5P4btApqsDsVsqZj6WUxC8CiVuVHhy28RKF3gkhvbSG3
V/1P6Kt8LnSxnb81uPH/J1XQRw9VYMaVibotcx5hTGyAFhKCQt/AFCVmMiwUDdpQ
rA5v6uMT28eRI/SRQYgt+9NbC6uKCRoyaDzoO+k6Ixjjh30TSVm0xjjHxENh7X3v
HcYkGroh2iG9No+3AvbejqWtsFuDxPQZsExyVNoEEOxlUMGbo3t42LBt70dq9la5
dYTzRUfX263vxjHi26Vodzl/PSSy9I6pyll+ShuE7eSsyypJRCSS7gJU3jbgOvDF
VSbp447F0Acm1MOGvLvqtV9mvd+HXNKnieFhHkTXyIFXl8wp90sgvz8vDJV+y2uO
M8rDjhzfZeN4Fi7ZJBpwbvSGGXzI1nW+0S6tPwgJXunNyexAUPQGMm1gv9NsHFWW
41xIUUUfD//zpJePTXR/QVrA0fGklkvVuIpdSlwDeUaD5R3JqlDPL8N3JToBbqRu
+KACLazQ9GEU08A2m44P6cLmxm92y3IO4tTMbhCRzZSvt+ZMnOK7CwvrNVUEqs0H
YRc1O+H4We68WkN69y/Ob+sRGejXwJyDJJGncTI/lud7znVXkOrkhGhxz8di7QsX
RAYEn+Ast7zlS1yW3K/wrrJMMUX3B8RiJlvMydfg/9jKK/kVbJOve1uuFNHvZq0m
GLvMy60CzidhP+pJDcNT9lTXYAkgXnCl4iij7aN4W/ADhAQA0L0MyvmtmOGJC10h
AgN6KA22UWGManqwgR/MjzLBelt41oMt/YxuWGR+N6H2VzjDlIOqD5oKp6m/8THr
5d7XeK6+uCuq/Mk/ho4OKNiOKyJ6NLKc/xPvqguoly+QBnueLFPDEyGmuSZKcn6Y
xvDj/EpquBEJOv2b2yd2PgeRNFdmv0N923/O6mYIAE9WDAKQEQtrnduU3or2YhsT
9XHxg/u9FwNTrNpzYgr1KKgqJ36aERl1cCyDWPX2SIycul88jSDJhBZQGIT9JhRy
eno3lKFJWQ4AInRqOP5ftLnhh4EvyzZGtIbThRoCzjUcdViJP8x317QIR00sn8hN
HKXffEiicvHxZMIihWHZAo9ld1tdx9FwMDQYrumQx/3i4pEF3DKbWYzSdir176Sw
KuCsE1IE/dwuxH4iQ/Ee9CBS1D/XHOciA2cBOCkzpid/1OHAuZBPDSnO+gmmszXq
bJusPs7/xWfKi9LqoNdJmzEAoPCg9ok2zI4uPQ0vXiDthsIyrm+ozBXGO5keaezR
YkZJUW9Fg36vkziT+ACLmPcR77kQFg/XLweEBsQWfkNNVAMB0ylEFtCY155uiOm7
r9f1vYZy7B5vc7eK2rrJfeffIJB/nyj3nDZ//oU2kB0RfhXXizdCUDg7otJ/OqzD
hSk36c9zPUH+79xhEhA/dwx7yTdE3A2AWJJ1d7ri99QbSY9fHzdDDqKtL4C6UKqI
lfACeoqJuQ6cgCS3StFXrOon1a2pFy/6Rxg3nTm5ZVhpdgG6W+fB4VfvcIOvJlHY
+7BABLjLY0g10016SpugMp9g4JF8r0N+qVEAjX2sLPKDK4Z9LrcNGeKHaggAx2Su
0us46FbRV0it2tZOWvvH5nSEkMCs6gzbBRQiGzAR+W4IH39GDcFnM8chva2wuq3i
TYIMrKK+iWYEolJTvIKpJ++4prUCWs19SWvlfhTrmJWsiMj5t2k7xQOp3v1AWMeo
PkRyo7xO9GPFDkP6+Coqr8zNk9/XkfJZY2wNhk/y4UgqP1qrTQ/IMbvsmj9nHCQN
kxzS320Yyo3WZeMeo7zwGoe9TbTRhvMVi9wj6irImlCS3dwiIvS8eGG5zuldt0rd
SG8q1KWR33SyWuOOH1Lw150OKHpFg+4zge6NeUeDDnUgKj9vAR8Z4Gue6MzxX80F
s07laJ9oUnft3rjH/ZM8JbcVRZ+DRjExr22brg8jOjVWaMv7jAVVOi8J3KVtJx6X
8yZypKYAR4HDXpPDSOXeGfoZy3by+9O/FADaJ6MADIQxgXma4PPv5nz4DVPj+hwE
6SBlkcyMn6ZnXiro38kMf3RI8NcuBQpCZb9UHQ3z9Lpjre67yTmm1rUPiRzk6qC7
+KAm+Xcxve/ocUVwtshVDRSxjv8MzsgDtc/hWAHqkulZOJksuw8e3kFemi3Ray/i
APfCyV9s5HcQZZ332uHsCyde/7QGyU80nQiHXLjzEFOX9c0DlciQ+I33p8aFJAJF
pM+pJ1DYxpanl+z820IHAeAgMlCwJxWOaU9eV3ntneZu0WfO6sbbrQ4774L+preh
p8alQDM4CaWhZJjaDRfRjWGx1n7tEsBCaxUJmcZ+QBKZs1A+jdKAlpdoo9dLA+Fz
L+jU0r2p40cDrwCQR9J3xL7dCEGLhcdTKZgs9pyI7cvMa7GspXbyHTNDD2YuxFwJ
u42fY2kntV/H1uaON8geJiRzVAMWwM0EOSva+T9GYCZmi+n9YRz/ZumTF9MkK9XP
hETwkJ4g+uDHDf8AV2g0bhVKFxbfcJF/c7E8+U8lyHi21eHR5H9TFpU6fEHPbIID
+QzaU4zNL9rcqJu1aFY56r39KFffDntUGSRybtQTsc3Md72sCqTRPly4ChFRDI8L
tpjyf+0i5K10K1yrRGH0f3EUVTqnL1qKWsv4ywUKAToxp/jS3/eCbiRqAoAyV5qP
a68WhDxp0FHSkWRDkbye+cue2oDRky/lwMTBmLEEquMgF84YFMgUg8ngBV80tb9G
DyJtGqDhvmO5l6bVCq+g7t/XUVuOlaWpjzFGtKOpgrZTCMorbEqOKb1tu9p1u/FR
lhevq+gc4wO7i0rTdeEsB1cTWUjTnt0l0tog68MQBDSpkauj8ZtcmgjhCIGxfCfA
mvuIZ9sVMJ/W2eBr1tFCaQnL69xxzOFf1W7ifeJbTZer7naey+/w+So1qMzEask8
mAtyWZI8aczO+0JYFTTVi5Bm9CzMDXuuQQHwlKpArvH19udNV+nvvHm/mtj9i8iw
eBjMLR61egZ2+Lr+NYbMRX5Rz5QC1THo6DNzqim92zoOdFjpyE8vSnMd+a+wwejl
PjKkgfzmtLif1QNJPokXkDEHK2fyq81HXJp58JO5EpMPYpYi9Ez0GnTj7qadaxeQ
rIw5/MQNKIFad6JQkX5bVuJPk5sqgNnvmv7+ARsB376VgFkVvqsh/zzf/sfM2qeU
J9Y6Mb9KYwxEd0udI4NvrwO/wDkate5szsWxDSTbdf7QNUgnNca0qcXUGa4wNrDg
Mxg6pt6ZULzzLfCz/cc8o9PybA4yccos7UFt+ZbPmTtuBUhXGFDIX4jvqvMq+k6N
Wp8U7AkQsgqE3ab796xVXDYr5oNUPqkRu10+2plFmZ4YVAHqUV/Y1qtGBViWadeM
jc6cCsFl/mmLcjfHLfbJkvci7uZ6G1ENUd/E78dYkUh2PiDYHXR6r0RSPOm5v8Gr
YKC5tMBGbHRt/XaV9/fqQKbcc2x6RvbGuwIhs9fVEfYxrp8s7EHaQ6P7c4POvRk+
6NoG8t9haYz4ddIQwrlkhRnkwvDW/KGqF5jLm4qcKQBazjGMpAPmj/mIGcDvx4xH
oBS2inrAgMni6xpXaYtkxarmOzs5ec3udLs8l6ts4rgxVNcTrDCjfKI3Riox76AG
5RLi8bhR+d2I9g4CrUQsTfY7OmSDUU5e5lJeU4lnq5FnfFC8YKy2VmbK7Vo7qbAY
SWTpmeRRInCkfooy/txDGH2txqmnfm7y4b1X2cqGdXqmgYbhfuoK2jL64v7ahvzX
UG9me1dfSp/6MZ1YtghgYMfXumy/eRssfw/hp6raBbkVrzUsNTPFwtirV097SMkg
9roM0dBWtym2uV+IRRBx9dVyJcoxOLzr1j/xD2SuAbwKd3DSU3bdtoQljY4hn31S
16gZJA5FPCKLUbjaTWw4Q/bDB2Equ+ZrisoRmdJrsRR+C4CJb97xckRbUlJQp9wI
nVZ1iKp3pdbaGsdJtBf2LbVxHKfcwHxJzHd0Xe8lOyz1OJ9sbK4i7RZ2+4Kjo8j5
coNeR6PFs81DiFCtm7TCrXR0XnHn1pnIT2akRNe1RaM7YklYzEnVx7zSNEJ+zzzq
qEgJYBcrYQaA5zXqY6X0B3YTdoy8iA1FGUT2+dNiq+/t0pkhDfuNiVLoKbp+8iNs
2KooKCjcXL0ZjHFG+W6qmBB6WspvzYaBZ05Th/dKAgVi9lov1PwdqdKOxRwHm37E
hbdlLxYNMJuNfVTyJqWr6iDvgm4vRTc/dKbVcYL1h/+7/8IfYD/mnWOP06fYFs5a
yVwdA6MO0cmFD4tsmtQhmU6X0UuwlTs+D1FcEaoxJ5vK98i7CtGPfz5rjnu4DmcL
unVQvg9aEp+L9ymEecrfgZQbED8UnGryoJ+S4F2hwQoPR6TuKHoZy9V9NHEtB+Na
Dk3aMjCtPqYwFTeZGWwuZ5ChsK7HMUnb15/U/T/bCUVPLbJ+LiBrDBvd2KWuVmuH
UH9z78DKIsz394oSybBfRhNLr1DeGzAnxJcyXPvxNNH21nD5spYgCDgMwYBsf8NL
Xv63Vq47kRRTugSaCFkQnteAqPs7YX3bFaaAOFneHn4feB83F9yJ7mDcf01JLAe2
FR8s4pWrBXFcHS7Mdtcmuj11Cm5KOHXLhD/Lsha1jd7JrKFR23B3dHC/28LaKxy8
SCu/+9ZFzSVK9y+oLVYcW26h3KJ3AndtjGdoYN7vHLvWYfjSaG5JG/YQAAzU2fwC
UL3tc+tUGMetVTuFdN/Vfzd1hBC8E3YQ4gkqizGObZ+yZuI96FTN5lUfGsdwfOx2
T0TP/otnXXQ6iQ14jurZcCAw3Qcts8Ck0c6BWEONe38LHWJ7isxcnI+mnXAtU5DU
tO59k9kmMuANWvHXQsKzTKWQKKLD1XOZV+84k4QmIh1gDEhwK+WykyWexc5X4Mu3
V1ZC3jV3GUX30sfMst5KxXiOlEmibvZWkMj2K+h+bJuimuLSJZun7A/tPyLH3yGn
V97K+z+nR121LmNWLMTcz+arkzgSFblZMROdbFPXI3WM82UsBpXQXH77g9gV/5SX
7Qx8DjrGyjaHiJLk/Hof6J4LZ8C+FUziLinP8ndWgllhl0iBr6MCL2t09D26UFap
CenNG2v0KczsuJV0MFfzybmOPTeIQx9FE0VedCzLEW2iFd1VN923JY0pSj3RAJBh
BnNYgrwh93OFKhHdVNtf6faVcsJ56Y3gmp0uT9pY7RbxBG/jO5IIxuDPQuQguX/Z
Jzkq3NLKwIjK8BrqHdZMgAKRgTUH1RTK9NmX41MguVcEfnwj/FvcyZKiaUd9eVPZ
hX12v75iPHhXSj01jLA0I6E6dfFSVcJk8fh320bTJDiFClV63pQBAxYy/Zq07s0D
dQ2weF4fUaMd+/THMQwsDmraRF7w7s079TnU7YZNM1qKWzV/TZwWZRo8neGht1Ua
JeFpTq9vg8Lx/01Fm9Vtq0/uaAz/DEiu6NTgEj+Xf36xIgBzDeIt8ofUR9v8yY/B
E1zDcMaJcaRrjOAse7lpd3BKGCgpwqQtrODdE/M4gBe2ItvUuoa8TqoqeqVBPv2A
GxvecSn7M+yu/V86yyfifReJrvmv4a0IJ+Us4Ox5oOMlwGw50iYneAJwx0jJf7Mu
2wPIyKeEazEpHUXZeYFVMXJDJ6kWj40Qx+b6omUHum/crR1ajcVtJEQW0n1z6zGq
9Rb38S5vzu8e9E8OKjN4RqZFrPJKQqkOfi2Q6fPgo0j2c3CpJbQL4BGOn9fat+WF
DvUc659Cy+rc3orvFZFMzP9KrlIHfkikttZ9Nnh3pRTlXDpKTz9HIS0sLJ3ohOPF
g0V0LLTNlzMIhfrtkSVdbUz9XLQfEBx/l/oyeHTgPmX5dmUdscYU0M9KCI+3kBXO
fdWLIPkZJjJ+jPcZ56e1vprlJggsrig54iNrBKJnXro5cMtygqSOI24D2U6jckS0
Mv41lIQbe7MowJpqT2gnm+Kb6DE1wL9q+yszUyC7nIaA6GADOBphkJjXj5gzPQ3b
mmq15wBNJ1hjmaIlo2g0/pdgEOcLqO/ZyhQaYl8di6oYkR5Qz7YDD8+mK08pfkxL
WEIAaQeiKb/OUZ6dONWDn7Kd9fONebQYwoEGdbqIFsrtynIPDutM9oSjsuSHiUYV
Dh4JZhmpgcYSmH7Rk/CoVMSgs53HDPr6aE1+PzZB/I/x2YK2mgk7E1RWSRAghgqs
2WZyyxLwGQC1bb3TPQoQjFgJvb56hVOctdv5tLRegSeiZiMANt4bJqI+iLZusmLn
7Xv/8GN7+ob/LmuTRwoUMdsc+z6zWlVgySgHxcXZJwn+PGpWHg1BtUvswuoiAd8P
dJki0o0qFWvnryLkzKIr7V3azPX4U0zDR/Yw7M32mngnJ3uPGFgtq2LRMWTWiFsU
ebRK9Rf3Zl01gVYC0Ktr/73M4GMICoMejsKgipp4eLRVnFtfUC4aSEfwu04bzQJr
zrY9VPvzA90dnBr7M5Q53ClKQ3K3zg2c+oGTcE34ayX4sV+G8h38lUgJjOAUPiLm
/uVQpC9VPWyXLdUMXhT+SJdSE2lR6HeoV7FKw3X/YZgfjL2Iuis3l/VMNtqElld0
v2OkRY3qMwVX1/ZP3DvypCS2pacp/LuXkIjjcIi0RarOYN9iha6x+6v4Z7MC9FAp
Bn1p759QYjLCdGTGaEsCILOw+2rAr+724agIP656tmW74cAex4TpSFtjqtNRsEfE
tJECGQPLvOOaVMdR+QgijUJtckJT8XSPhp+EGDu5KxE9ZYfwtXrRqaKFUWsweWUJ
b+ZihFKSDd82H+elr+Jf1YMxdX0px4WSCu01r3BY7GQ/iumiawcK5vcEjzyvYPks
U4H2aXLRsSLvPXG+kivWDr6H2Ji0ZiwbcOZ0nslriFQVI8lo9UDLTBTvvwJgz8KA
mDE7Dh8l7qaiqVhfU8fJQk92r/8Uxh6ash7k9B1eWJ2oPVxWb0RfPV/B7w88U5o9
7FS33NnfoJIBCtzYda/Yk1KUBfkPZR5k3CSvKT/eIvgYdF1VoVhwpGaBoDfb3rN3
+F3dq3YMgRMH92YwqlGtFhRL4LtLfJbEkly7r128dkAfrpp39HhCXWMYj27L1Cnk
1KI78em89IDqOLXC9qBHmUScK+G/gDaYUf7yEUJtZTAkZ6Z1VEO3P/m1weKgdiB4
pACp/XSLjP4SiEHIKfsrQTJ3+8Hx/E5pwW47EUnYPm9c5g0gTBC8AHnDj464vVG1
mH4qBJj7yP2zgPBQYXGw6uIA61FTTXc/oizhH0YKnUkIdXVwH0qqeGsOGeWsYnPx
8xi3aXveEzATkSvSOJTLBU5aye3yWLQU8CDE2bMm/unumgyINgYYuq5e5KLAe/O+
SuiSv6ouVBpksDFsUj4I31drsYES985VwrP+rxvMpD5cHcpVCTgrTECIqd0N/E2f
Cy0cpibqahlvqi9tzPS5LghiCEYU4wgeKc/rOfr9rvOZHK73qqwFpr0EHN27YdL0
V8t+E1mSd/mcNjmjI0CI3DJluG7YDPQ5Z7SyLVCqmhN45u5GP4dv15XbzyIXWQ4j
+udDOHHAvc1bgu2bSGFx+y59llBxGkJ0AaUERa1VW10Jt268oAuN6xXXcaCW9sWO
3JxxJJa9a/YYnS9MkHOfGl1aIqehKsjunq14x1Ap08u6xW/YpCuxZo3w9W2+NCpn
9eNUN7b6XZmGIeWIiIIRZ97eDymLVWGHWm96KfjEou/RumJjK1aevzA6367QIKTE
KEjMgYLAQ30L1zVHLhhL9NkKK9UHJr2w7OrhaPTp1u43Q1P010VGW+51I91ZhmGm
GIPBAdGRTrfT33/A7v9KHUQLSY5MU0Whu4miVMk8tktLyiHO7LdrNKLRw3JBQUPf
ZKAbjAoWMe6Oqp1Wv4sE02Ko+7w+eI1NO/f0CUcsOQTrT3TEe5DYMShlu5Gwq370
rp2Icmyz6dzwEmVdZHNzU0iWnIL7dIHS9r1L2c3Ui65IRtloYu+e7FwO1RgdkOZz
wjKMKxLFHLLu9FbrRqUs9XGWZu2cea3PyJCsUHYnbkrQaRgC17Mal4g5e9B4Uuka
fSaFfgbd4ox6rSRNo8I2PDLT/bjUMZkQTEE07mmxky798SxUy5SKhqbtYo2GHBdb
m7ki50vuBgwUmVEuhVszZ9idZ9dJL1IbCCWTfKcyL8Ke856P+GaWH0tAEUCmTEEm
6zjUxXCiz+bBEnTmXUzCsKioHSRcz6RAQZb+lN+S48rFJHfTwwoKmXCpwzmm1zk+
wjKXl7eOpJgNgnwk1CWRxrYSZc5kzw7yW1ANhbUVeKAs5EH3Ko9tmrUuL8O0DnCQ
E4RHix5rjkBTgSFdOoNaOB5e7rudwO+u3lVkiPfOBbnJ2PjnI1rwaf1Y0UOlIIkl
nNa4YzDLDYjRl31J80fadhKFPInI1B5BIGCzI515KJxLpkP+D0pXON7PdvF/ANe8
OVaW0H590E8ZuvJTb7Q1Flw67kU4WJ/yQKvA9f6DooXLIHdCcRnGBGjzpITHig/j
qN90t0KYk8BbsVhEwg5k1U9+OM8VEXrtYYoL3z+FtQcu9P6mdisNkRZiKluMWjs9
kW/nTe4N0X+fDcgA6/ORLGbSndX6Zz4MqxLTPKNf1LASnByiQG7kic15BDQas9US
kha0mNR7A/6cpQrsiyDOl9i4UuFLxIICFQKaUFvcgOs6prtsfH3IovDT6KxQK/iX
2ufy2nICOhHeYjUw2/xqqFxpZODs+16C/z+SpZJ1y6ffcsl1DyJKMZ512abVuh0c
aAXaIyFF3nleE7H7gAn+6euzYqPfV2spcm6DnqQaQePirMZD3ut0dFoQlyEdAzir
N5JBPXa4a32K19kdDbDT6eeXBptClcwuNARSHWlcsDy5HHFmgGxq2rDx+TzvrnMa
+mf088x/kiEI1beTHpRMlznJU+18ml3TOV91+kpvhqKRLH3k3Vwe2FKGOOwdjn/W
U6enLB2B1q26VLcrIKPLdQ/hBmyWhAvOpF6/WABJuubDu7m8pV0K6xrRG6C1selB
+6wr2B2hmpEp0q/1qX4W1BDNWp/v61fQ2m8k56uGIXnzWsvmrdx4eYjilmvH/Fuj
EdFOcAQRw6OWJCf3gTd1+SKsn3L8iHD1MKbK3g0pIIHaZxtZbqGG7AXQPjBm2Bcd
SuZYo8bQvBkxvMtb2IEz+so73vWQZw+cNb8/Zxxvx6FWABr1e7J3DKqdiWGxgwCO
rdG1SGOwmNrbmvYFFUss8U88pu/GFfeDpLRGF4E/fo5iBpyVOqrlaFR58IfcTWTq
k0zCzV0Ciq93E6+2p6j81cngJzDEQfAdgZ1lPOaauBDzZ+4y59DUMw1wcOyLaeNe
AdMaMkPUdBFfiL4XYjvoqMx11wZYg0V10tH6/d+AuLg2RZcfZi9XY7nEw39VI1gd
QohbWFdDRiACm+fC7VZMkEPqVxbsJhfH5/G3n9H5ZpdXk7WXnC4uVn+ELZXmR3zY
hO4uodLltXIwJBMvPHJKHDrH2W8ussxZQUJZACfFf9HpS4shA4jkHCSEdNKCRpvK
oBXo+fu+SLGAfbF8afP7RSWQe0iB9VdwoXeE1p0/ptJvGqjTLMP0iZdJTxtCIgLl
JmDGIDGs6MK5SuNptD/iCAsmWF4ASHD5Upha/UZRkOswOwCVgbEyBDMMQaWGc66B
umKemEDyrrUxkJ2JeJ8PC1g4zNCHnjYUyz2uJkoCq6nHextpzRALhgFhpuHiMqxC
FkszBvLyooiGw9PpoGKj7x8bQzVAmpRUe12NKh7TpRJQJy6jF5l0mczooUFPqyL5
0sEuMpWaMB3AXrlIJ2F1Ry29icxPgPztv7xbhOWXjx+Pp9IEebVGUeLUF8XS+AtB
SJ4hsp6eEtfgJm6nauDHv/7mD5KD4tcv1z3XKwfyjQIuPTauPo0vz4WW+Xn39YsP
+c3K383fP25mt43ZCU5rGgKTNNDC33eI53mcBPifk4nYPCWyGV0+WhpeDv9rypJ5
ar/bL3K6B7W2KiXRKpnKNMiqVK7JnZX4gfkEuLOy0kVEzcKpOMs9geI7Id7talZ2
saZKD3O+qEbdEwcitw0YcX42WsoYByYgSUvVBAxIL3Uw66bZDmtrZHeTvbzOCYkj
JlzOFe/exdbExgZTzO0sXhRC9sgvMAgVsnwsuuX2yo4rECea02vaTNOacSygAiwr
FUlS7hhVNbYODflLAF5PsE7VhVSQ9Hc5ZBpFrsMaqzPYobjor9YOMPhfredmTTyP
mTeIiAxhrbLnYltPBHB6DtKBrkdQWpC0dzVSGygTuDlCBDcgp+8OmKEoybjj2fqg
U3XNd9+ugK2c+5YXo5pKBI+67iR3UFTMhx/JIKDHzFyBV/DiiBgjY4TXECUKua2W
amwWirkQUdyx1JLoF7KMaQd06Nauxs5mlroNdTdo2qlESgLbNYzY8ohbDTBozrZl
0XJRkdHcfbD8syJ6UAOrxoJeKbapwsk2lg+nPLGXQOlcnaPeWWLXqakTD8FAXojz
0z+q3/K7yOASGX0i/eLVtaSvr0hoOpcbceyVXVmdQkja3fFqUcaxzTQv+7kiPP8X
Ff0XfY5Q6D0ZzU0nXBKDXEE4wz+/iJsupgEhL0rin1oKtmA7NgVcMnDlzsumOCUf
AFTx1b0W2jX+/28P/The1mH0qsnKs8vOsYUbVlB8UtJDIyIHUuLJG9XVlQM/YCl3
T+Zt6Y6o7CVIIWKwXxL3apPdldxLMw3BG23/dZl+glhYeNJA5F/g/gLujVWF9tBl
Jejz9blnuggfXRb5uhRFIZkTx2YICLRFIW4GDGWKPq4GaqzS3cgWoaomcJvCsW+b
Gwal5o7K9nP5YzZXrqxFMv7/Drssvmu1nMNuPoShCGG1gST1Z0+aE6Ebt7p6LuXN
lvy8Rvfr0/ATSQmPsFIZN0tndJEPp3k0yFwkux7MCcLe2CmLcMXinXPO9o/fKG5f
TjaULWP9Kbyd2PfxnP41mbcZMMExqYtNON4vgBc/vj+7k7+0EloadUqL5otycqNg
I5H1eszK0j6xrpBnQ+T91wEVLnqg1QzsuU0Efxtb75I/EYPbSwia3pPUCsCcSvZ7
Arg1kmz2RXc2P1QUoY5bZ348ED+ePMfvYsfc7F0AEFU+sfup96O3NFJglsXXJsj2
RURST696SaTT+1PAzIQ1DC79aZQEJ1cOQ6MK1eJqqU8HVn+ZJnuRAI62qEb/bcy5
UG1LRUZ6oLxR5c5KATrwtwPlLcm7Y1aGg0GRuL1tndqpikCc2M/yI2+I4M6OZVHp
RJONLwfOxbjAEtPNIBIqURvFTwfg/QG3xPgXP+cFI0MNaGu44Ptz5G8ELBNJLx/R
l1axCNR01ZaIjT62QdKGZ7DEoO76rCYAW9GGJJhndZ4EI1Hr/lbQwUbCywvpudLZ
L1L2EgLCc79LhLZpgQGgdZUbUBua+wE/cTIYo7taN4TXxGN76+rRolXIxVF+yq4E
j8zyfRlixaprKjGhagu+QpGgjcUcJmjV/PN2Kz0SU26sE0Sa0N7wcRazUKaR1t8i
qWobbeKRSC8vKMSI6BQw7ImCc+MyCVyZEXfs7cD0SEasIeqA/2ufsFrOy+zhsCSI
MyGTKR9Bk8AovSY9CrIvSJN1x0TMD+G3JoWNjPw39cZdLOsxUwAGMWtyrpW6UAeQ
4y86x/wh/8C0lKVHVpenUg8c2ZgDQdQnHY11bp9l63h5LIbsjRsb0ECG7Beb6z9z
LY/+KzowyrAryOvrPWFoSfBswYU3l8mU1mO2/v6SeDXKpqlZ637QrrSj1X+OtJX7
EQEBN3dWPQ0YfyGV7uC1UW1crxnK7+Xl8SrsVYvCWzfWq01gH7ytJsb9AOd7wtft
u/vDfZRhl7vkuI3vPxf5ZVjPwecsHLO8sCWuU2fTIo8qRT0IndcEJfj0tmkc2nu+
woLKFM6snkm2G+vuPkiN4Ja8SqbTISoid22LHky3h1VIOpCoRNQhKRJL83zFMXQn
qreo5nZxw51FXCnvCdGCgfWsQL3JafkKIKQWL6p5FsE6SCMyf7i5GZX9VJIp1RBI
fGncIcazx541g8fPqeiOA7RYhC+LhXAK5b8JGqccOcAW6mHnja9oYUK2TFyCKk1K
4trVgI1sz9qGMM1No4cF1xLkkkwwXUn0Vl9ZtQCVS8GA37GmomwawILCBP3fKYFa
1JfzSOntQh2nr9dYxTVvhkZHScau1gtKzEG0e0gPWdHAJyZHJvAFtD4AFrhdoiF9
zml5MrNm0zFO664cWz76YShr1dGRVrRVjGMv4trppLql83wuLL4G9ET53AgUFA6F
DkJfzNU0Pnr9oQ4L9VpvjV0fCwmiTTIe+u2Gbmrilq9wk2OaIXSASH/WKSRbilww
h1xqKNICYMBHFr4DqTLt0Tec+pb0+QbDygCykN6BuF5eHwjabtvU1JgqEvTcbRnP
/JBZSWhfxJR8lSECA75AaF2hHzcjFMBkj8fz9vUAj8XHWggHMPugGFDB3JXPtiLY
mlBafhehR4QKR/XMhIczUr+38Boet0ToIhpp4Yf9vWeqnBm1mve5GFwVZTlYjlmN
T0Nh/j5QMW2s7/2ABoGedRAtW+A6URI+PvYkD9d9uBeu8BS2E/RpuAwW9dAnSBr2
ctvskdFfGp4wVlWxi5lAzIXYX1z5k72uwic0coM1ZHPx+eE5sE6ruT0Os15SNcGX
3iAyp91++z4vND/+ae/nExPMh9TcQeWsMV6xjjaPa6akUDC83hqeJijUBfF4RH04
NVGm18oC2fA2RPQUJolviLojAQafFlv7vtO3Ox5vb0X4o2z1sSscN3oIVQFJf6Km
vKkDk8EywRg1N9Ce0N0Tgue4yaJVKhqXx3PeiFz9owntXoHvlM2sAWUoimZVgzrl
YW2BxWL6JQZ/YwNxjqx7xtUWd3m9yDGh+jHaQ0BXZETd86/GTJzl/VU9QvrEdULT
Z1WM6QF3V9K0XqwebWlrOOYd/CGwy2XQ8Q6/MDHrnsT/MHJJxmqyNj5Jw4e+6ZJn
EU5iBX2z3fd/fqH1W3MOnUwrMEetl7ws9s7ibc4MZxXDeLpZVfaPFH4WjXLRZ2VP
wX7V2C9nOvFGaE2I79KuZ0Smv4qf89n0U7yJDIxU/MUk2UT5mYwMljUxBrb0wr6A
hnQpPIRWItV+xk/sirZ3Zj7jH0jgSb1r0f/1BUeIlGtJATqIPSEfKhJj2h28ywLj
9Ff1+g8sHq/92mYqPYqd16HcEb/ATZeEgpdhwQ1qXFukePAx7Epd4j6Y4RUTIvWK
UXn+D2TbJoRgNuThQDOr3/9T1Q6h9WV6EtUHx9vqlazl3w3O7lpMDOrTmXQpXUJl
utbb1wGV7CQ+u35tenhPih/BpvluVUVFK4v71EDaT1PS5s/sl+iIjj2+8tZUMPe3
QcnaSgBJwSG+8WtbtFOCMzd6QuK09y1EH+YyZD2teTVXUjYbSsYblIApH8/LiaYu
PRSBshrcJVOMzwVdpdux3WNaXjskGXdSxmVKOkcMiea2GKJck+1Xa2A2+SRaNWCL
h/pJfidoBEtaGu4P1cJeVnDWFrnEIQDxszfxGaS9apOqxIs0p0HaSUPSG0yXEHer
xZLby/HEsJ1sHDleVxmzQNoCn88PERgArdCwP9LQ3mdn+GbkMAuj/zRusPcaMUQf
1ussmUf3AguSWCgyIApIo4irfquLwd491pCJcLjkrtdlRHnPAHkvKvdK+ZFQlzX1
hz9h6KPh2Dd9K3jFhimSjRNGdRf8247uO+S7kfPCpC2x3kzhUkuWPiBkV9NPCAMr
Hs1xw4HxX077IZGpSwJxdbbuGItIZmfORaDKCX3zomtlXQV2yQoDo1ZlueqP2gzf
jfltFvi0c0FlkGho3qrBik20cDmQSYST7s74uMCB8Q+F6DhZNPmGQvP/8bhofO2V
FpR2EB77XKqGRllQBRqfhWYDf72IYzHIScJfbbRfDkzcfJLbeS49dPtUano9J3MW
QtX82gsNGE6CbBPZ+RNeaQR0s8bc1dgCKpYIVlZANR5tNKLdFACzq7VEYc7vdhWT
4wrMTVftDKb09poX6dQoSG48fwlsNgOTRd8qOKy4w6N3I1bdHaCwqWJrkYoxxuv2
2/kRiiyNz1jyBJ60s9oXQv3SyF0NHLwMCfRSnlTq8iMA54H7DYqLuYE0XNgV4Aea
jmFI+590ERGAJXzaVSrHAxsuif5IcLHH+FKB5SoNLXXyv2JQDtMSmMNEWSshY1Jp
tRtw7ImMgph8ZqLZqRg4Y3mjTERnQobOppoKg9MWY2sWdyFVsBrKydjVGxLaJXI2
t/CJ46cRXljB6m7aQF+dqLR7EihHu+DdLaZC0VP4tnCVOJ/WFURh24NGV4E/+w1g
T0+2uuTg7a3wSCDg8YL43MBK3iHaQAv4MKqolvXEo6hMQdmSnoyncCkzurmCm3ax
W3RhUfCSawNdkiMkxkui6a0+dsQXbepmGtM/dIl5OSaJtdQyKHqyDvCTeK46b+XS
pHMhGLD1r+M6OnFl4aNaHbUj+j8qACR6xRXa8c2jqZRsd0OiDaR1boBqlGjqaDso
eqgASztEGpyS+23NM15z2U0O7XL8QLe7xb163igxfbVzXSRNiDKe5KNoOiLYp2G+
O72qmnHRhpHE0SE43B0yFhaTJSrm7JxJ/pMxAjenQcjbA2cnsyjnArkR0gRgKD2P
dqLuggkGHDtIINsJTKspq6HT+IhvLLOFunUCv3ZzO4IQvb9e6mHZAgQgXMEgyHrr
HXRmeG7VX8ku/E/wltr71NXAqDRZBkWiuAIVhS4+Meb48AklAqTrupuVKgQmMKRG
TEpG0iJXxbCJuwG/ZK1BQcfk8uC8MizyRJHj8VZ42cGu9pU166wqOu8JdsUFIX5Q
R+hEP1/OwxQYQb8a0byZASP9W7A642nd1HeU0gUf2/k1C4ISe1UIai/IvPq1jYNv
XzBxFgWy2gOpyqOGBceW6d1zTatAud8jc/+SR0zmQa85Po2fM0s/k2ssJbzqQRsj
LCWagGxAtkh0A/t5moWDqYjii8BwS1AUN4uTpOZ1Rqe+2KEmi0jZABAIaFRtA+N6
t2VIT7siWDJF9QeB0JpMYnH1gVys36bO2OI6bHLf2I/qXBN+FqtC2gkVNU2yM5DE
iNba53+od6czv/ijgUI+HUoUm8GpHM7PKO3AUs8ajGagO7I4OsK2iB81H4G5l76D
5L0Z7wJnDWs0va2s3dSv8MRt5FufA03LjQeePubsHfHEaXpVOT+JW0rvcr0ekIOI
huSrZP5065ilw6tooX2UdAkNXGIw+aJzi7+tzjCbmh1v6tu1UFdKAZAs2nroGVVo
uR8n6STyyKq8JhRi+b5CiUJmaIAFPaEK9fXOX2aWWo/GnsxVbOXAnCy8hjv7tL9E
zxuc6JzUyEorcRw2xomSJNe1X/wCRnKs7tSu/pwvHC4wg22DgMDVJgTMjhQ4jv0g
hqt0AZGWVwkC9b0OW07LpSz8dwr+UmfYp9eGxbPPaoTsqq3fz7Pfrfw+HGp0GJib
VtGRpopAwjaJPhyrQtnEt+gfE9KkIeViUFqms7sTtC7WtL+f0N1LgmGn5hM0350X
l10kJ1+VqBvHgCFtNB12AB0+Bx0e1mSqg/o2tLunNzF9WhaH9tSFgDm1xwmVlV19
Fl1hKQr2J50vOtk2l9HY6eDtR39iOhiWPoEgnlzJuMz5/oEBcQA1Ia4BFWLSUXhV
moFj0r2R7WQySp++Rsnqogj3g1cVlZuqJPiVUyGSwvb1UcCj3q7IOWnQ+7A8wg2D
0sVEZAD0igQcEvy0SBQJroIvV8IZGgRCEdPEXRvaWCUjxeNpmXtrXN4H2xpzpoth
C6vYaikyQUNztdNLvVeMx/Uw/hkfNjcUy4JyU/v/deLKzv+grkz+I2BkysRi3pCT
aEpkoqMCDNRoDB4+83VopHoowsO8/uXu+OPkNqXdGpMliWZCleTSPhKS2vJD3f0d
JjrAHBtU91eww0zbbX+mLKzd1imBA9buo7CL3ZzjrHEJErHEqqF6XU1C6/hxntzv
YOiKyOdzBa1wPPapmvkjoX841RcmZKVtEipyzGD+RDmiN1C8B2SHIvk6wnPHdtib
+0FbS4RUJbfoxlv5PTzwd8NXP5iBgl+esTLCEAY5cjpHn8g81PzuFkT45uoS5T6l
oVvFzJckgfiCWSCojWbiDZ+mpnWV3vzdVT4Fs44sPBh30zGyPpPYLXq62NyxPq0W
8KIWNTxrHx4VPv9kCG3NFq+nDkH1jcp+RynlXo4vG2xQ6aAiZWyHDkJOEhNAmGPR
7SfuvXY4lsTFuAxuSlJDOezlI+nhgV5rpoSbwaBZOezmWYY823hjUjArEPRA5zKw
XbP7JA59pNCkryyqftlSJYxnHlm/RjKZW1ORit+6BuErBHOUaMKjURsSKmrU2Zwx
GqbLQ6nk31sTAfsWxLiWBn5Hlp/935+zyiFK62oE6Td6IkUNdNNHKEXZMxuQ5+GV
E3nI6z4Q6/0P/N4bvFQ9nL0cd2LVd2YdVs7WKf5jAMaJC4RuQCkK38RCZHlWqIxv
tCX6A1LlJMJ4Gx76s7kgzmzgRWwyMLlVP16m7ueOnd/069H+Y3Qs9cMDvwEK6Ohz
DpoEBY2T7x+H6IaRnGy5PA/XwaR90FReFS4crE4VKkzOwbr0TX0UUX0WuzC9kUxI
8+pWfsfeC6vMJgc45fYR6CrrcYmL//JE6be0lw3Q9E798evYr6OlJQ6YpBAYdXqW
OtmoCaYYK+HOuUfB7KWdOWuQY9kXN+QHOhEBFxl7QlfbFM0DbGa3PfJ7ytHkVi2b
V6nzDsDWdIbv6d9+9BS+FkfMO2NHRfNQlJRXb93YYflD7CEAOJ7DPZg7XRy3KJxe
aLBMyok7BT2YKijBW8PeN6elnGia1Os2h3WDH75BTfDfPxNKA+3a43mXXLxkusAB
k3CJnZxSsL02nLUMCNSflOFSeMAmckacTjDbRLIySEZN22O5szd0Tt+pYVe1Wi2b
BcpKR3uuR1QA1e5xmqC8UlESfiIZMZ2+qlzHfAWGAFB0jq9l93+Mfq7Zeyrv32J0
GLI92FIzKFRPlqqCLfD8JybvS2ipqPafmKmY4MWJ+hJ5H8jFHUympm35OHuoSwQ3
zYuXBUMbAeRtmWnB69OhCzHtI+Nc6/FjcPP4VsTetq+AJ4cSfsSmdYMA58svf4aE
72Cd8ES63lO8JiLyefkgnOmI+8zpgHCl3F3ZOlRRUtFvjy7yZmUD6QyaS8PZlSSz
mZH3iCPafWWHMCd3fe4EDhUMPnQREqPw6bjs2n2U7+Gh4U/N9iu0Lb8X31VY9W/c
fouDY48f5pQSwrVE8s02pX+dMYYy4+pvKW/Udmwaxuj4TITGAh+QHgatr+HIq/rm
MmjxhvSrAoaOJbkGQQ1J96gdYqVITKyMk3jap2GghzcOuCQQJ8lQ9Y9S3JGjuWIC
DDyGuE/oy0UlBn8tvBze1CkE8YTFDMtld5NiJTxVHu817vxjwGVbb8Y28U5ufrDw
X8EnF26m4rkF2V/p5q5IO7jQSLWdUjPpWUhGyHfLP6tJC4OoM6q30TG6IRMOgs4W
W1qEEncOxFrt7JFHppOVuG7uGAEWjIfYpl2p2ju29HCuNvKCJGSL3+hdrFuGKnk1
W90MVRSvKsfI44tGfxtn21x30+UDmPwhySpUZy/c2+U0Id0LFBuUMQzrp37luD/v
X8uuHNLDF6Ob4+6fURMGF0wFWekh4BV9xwKx91ObKR+U7fKi2i//3KFN/MInXkgA
hVaOxT3jTJJzKN955Q0MpDDVi346cvy23/rm644a9lzEREX06Nie/q+Chbug1txL
J3bztILyP7gQZerI3aAQ8U0aMD+S3v5YefV2lqqHzDMX4xI1Y1MMJYDAUvVR/9x5
zZbwsXMo41v9hzRVh9NstmaRMFK5yFlIvoP5ejBOTU1vlD/JfHC4AUoBORSVd/K5
sKo38yg+IufhCDmLU3NOPuh52stcpjaxDAmrzGa32ZPkv3Fq+P+MaxHqcscNuIxV
IOylwJpc8HpUltqMf2YVaF/Rm4I4gOatlq90VJDjC8s4dK6eos2s+FbSczuwmKlH
x+EZ+QZ0alaXx1i1M0dJP3m/wmSiHN8MeYiLIBh4mZdxteixcmsbH+hO9ZJTvaSg
7mvTadiKJOQ6HdsGQ0ZdJQfDnVQ6Bg7ai3HXR+mxhwdeUywJZDGUHuFrR+9j2U4m
1GYpzR3aS0hmf/li0TxN72Ue6QOhAYWRfmIyG9Prwg0SLr3jCN7643CEV5M820BA
/PvhU3N+Y1Xj2eZKyXjOk8CIqzgaljFdIUedwvk4jHXS0ze4Z3DFpgbXhIgn0WPb
Zby+2vEnjmktDlOW7wyRjpfxuGT9jb/XGmI06/aZR4cjjpj1iwWVIwOdIb2xU5Hv
lULQhJFrGYXpWUlB/W1hVK+lClv/0oM1xzJuKEliuuOa/QGDjfPlyIB6oLgwGW2A
RJVNwm4vSPlufOSVbQvQRhFr6P9kAKQkzR5RvROQHxt8ruS0pw2AYgI6cm+sKt46
b76E6rZjSlbZtbXRMTVjF2EjA+TbSBMeS7jKcyNfLMkl9cRoJAVETfEAd1scTpmc
LLBCLYQL37LqVjhb6vg2APXRTfSgbJErZbGnJejYRUr86y+M4OzJ7wQH/i4kSsMh
OehkMqBV5gJcp79DHGS3YXbWBTfI0TQTkKxoDw/FyfJlf/X1zJUrO9Yhqkry4d2o
ZkHx+W5kX4CMyKth+W96eF4DF4diJ29t1t2Q6pkszSRohPb7wn66NTVovZc9+foC
CWV8eo6hxVVGN3NPgksthjeB+U7htD7MB0AanFZKbChTKCbZc+kIkczsOv5uK40h
7hFsoLyozRySpLcICVKtarLJBrnxRFFUfMH/aGpKuYfunEhDNEU6k2RQWD3c9OjW
T5QF6WkHeG4KReHPwb8FGP5GTO4zRxwyGMqdQNISDWF5B/pkr+RqB01mvctK8DCz
DZ+eNJWpZxiQc1gl/VHVQ1JWKAlkWXqD16173dfUXhjW6PYuFiM6iMoV6ybOmdTk
EgxfZYzyLAyrARHxbX/DnZtY8cK1Oo31pHw/+dDNHIVj9xf/X5XjubPOWgh8C8fu
WRVuhpl+tUyXbKUlVWPWwKUu1LxYdjnfY+V+Tpob9aDaCUkavsKgWY5WRWETbYjC
GGBQmPzbVJt2fa5UnDX4IrmwOsOV9ecLz5amGitGE/FaRCdvgTJX9U9Gp56+otct
ZpJTHCsfwNfuzPKIFrsBz5sdVXeuDoNbNft5y05lPRq2CQtmikQPX2mvLYCGRDSg
00MD1nm3B6DFS9yBTTg03h/Gct+IJDA802v6MQTk7o0ee/FPzrSRUCfRf8Ld2pOV
YNdX4m8hPrWOuaDO0pSwv3MS5aD8NVMtye/UTzYNFVwL7HqNvgUtJgykyPTG42IC
+/Pz0wR/KCFXMxz4iSkmoI/Pzfa9uUmxOxMv+mDyGngsbdUvd2RpcNX2f19AfURL
exHaoW3S9Py7SFRDGA1x48blZV7MUY45EZfxj2+m6LtZaZERenqOR9iCA5XHpYDd
MDCQRv/nT+N/0+0OCrC8FtqfMCokoxOH8QnZn2AXd58auniON1fUn5uavfGfh0Bc
Kw1mhMgZXS8df9KJzr9Pc/vjJR1xe36GS94YihKYhAjjJLTOUBndnQOrWQLV1Uou
mtbC6Xn2UndoEAL7CGPFJgZH4e5ykaGjyB4/MsVvym/ryZn79Tz//YR1yR2qE+kg
Ld94Pj3S3shCHD+FbnyZ8sr3fspkuZxQy16A7e82J6fW7z/k7uNxBT/XxvE7m9Qa
TE1uqWyMAfVhmNlT7ixO6SReHvgB5Crg8NQjqPf7v/HLZ1M7qFlhT96Ql8tGMhii
7nEM7K6G5TUQSvOCCXFbH4deZyJ+zvIT5uFPwGh7gUU81u+wVeUJxtRaSHK8NNEi
aToTE/E/CA/6MUAUd0u2re/p9E4vFX7wmA4P74km1ARw6zRNdTnSbp1HLuZ8g66R
4TcSc+QVYqDOkXK4jmIxTrWziMR4w30fXRg3yTHT0+vm2Z/nTNHKb0DlfE7XqryU
XvS1xf9dldCtxtxiF+GAwbyFMGzloCg/YUFVLA9THe/YucourDX9GeYCbU2ESku1
i0z86udUz7+E45O0oWMGaGBlWnSknoU/h3Y5G2hBj7sggxpzLPXpf4sVi1dXKShP
dptQKtYp+w4D9rpV/mSAUs2nLsDB3saubEJl0VSQO6gR9WHOtpKYyeqCnAxerMom
O4okIQGqlQczOOOZiYEu9te0rPvTgaemdPm+KUpAyPWjl5FGgetfqnxRqnwddVxY
7EDy3yCsqcVJ/jI2veWlJ3+AkL6AKB8bzueGAz2nbKFBxYu9OaFdbqb6L9N+CbQh
Rb9Op1a0CCOuLV6PoV9aJvjHoY4GUdhWARzeBiGan8DiB/CLwU6HWnZQyk3KSN9v
pEiDrJPeL2WB+Knbzcs9F4oZosTkMJdX1/CVFlK+WiuXBriw30aMUprw1quqNM0Y
nU1tHi58wVoyTK2OzFA3Y+qnMcM5TWEsRZuE+z7NMjehyXUtmTOR9atcB0dvk+Xl
2yVQRiilz0bQCzuMAshMg4/eEjtmoclNlZ4BdYwelvovQ0LOpf0rZN2ruAkcAEjc
jrUCn0CVym3+p5+3IzRC2Qy3tn0uXdKtwgZUgwyuwMLdOFmupILYOzVOGzOZtVkM
a27rHZ32vaiKk4bvKMP6kMEiBXafMofigzrYIEWJ6sCp8hhhgsiLRr1sfV+B2zfV
jgcVqqRdTdPtxUaxl0IxyUvWw+lJ1YTXBcPFDLXCrg1zQskOigbaSA07HDtxOc2h
y2thuDH5HcZmra6mFMJNGkJxD4Bg8KMpPyOrYq7KC7S4of7uMOfB4U/gtMSrfiew
fMY5CWsLuCpuihuMfDHLxFfhYDA7uBdhjKAetthK5uEsefpSElVEShbc/ZCprlyW
17VEXnk888N2JdX/i2PfqkQWjiVVDXBs2IFJSLDvCGMZv/0pc6IXSubtqlOV2O5L
HJqQQYU2rWTAFPhRJyxaZxU3N2bSW9WYXGgr8MXvfHYIhMaddwLh7bM3wsGTN2gx
dheZI4VFe4GdGeiaB/EwbAff3hqgD4HBKDYbHD+H9lPKp62/fOKDOWSyXCjRBqeA
kV7U5WGGEx69qMc3FcFDpFJTR+mTM5El2vjRWSTmqozMt4rBNnuIuEprZqPPdsiD
57l5EWtRek5ACYrdaXhe7RgQC/s/xTw8kUpGHY01egUuBLdUI/7x2IsuRPYjgL2g
VPf0Dt7H3T3ajzFHd9bSeJrYH/cryjwoazhrLJB2kqAV0F01ihev0H2vmiLjm50N
bnfvCIbLrR89/RQu3tP58SVtiBZbMAyF6er4d5l2USBcYIAgZtsKlauDjIABnxoy
l+h9obPtKHn61HjVkTvWPP1+DAAl8Bc44r+hwzYTXToSROO0z9mEivdhH3d/cAeB
YgNp77nb6pGuZwuAMy1gLZnnSZ59BwFlwvWYW+EIQbiLU7Mo1j3BcpU+FGwkGYMl
AjWcyMH4+whusKwVSmD7Ffxx6e92fuskpyRehTuoDwtErVXkjZ6cMIhvG3mTL/A+
zoKfHFI1H6nGZ885+jdJpbMnpPbatq65Da0teq9z5KIE/AwrIaqwBYDAYxKGebKJ
2NQb9rWe1cYtUHNWCHViXbVQV3PnEZVe1vOkp+hCDQQOMQ389VIGgCe6mVowaEVx
c0/7sxmq4aa5acmSxJnJ37yGmmZfEcmD+TtBvNxeLffGgZsNEDHnfNo9bgP2YZxY
wmi/DUS1EXasAAnlqF62u7+aVX0F7rujWAkGe0sFH8K5v0IklawF92bp6GU50GgO
vjB1HhSeSkVT+QmIty5fql8cB19TQOwdF7K5OyIcyEo4i6e84ZecEfTl1h7tzfq7
r82iqjRXDUYWdXd+9xLR+BttdWL7cJoR4J8HW7CLsjSBqM8dm8waWqVwpzvZhxtT
+e4pX51IJ5M7gFWiYpS4+L1GajfcivBU7y0RaHiLR/eS75zhdY6perq0B76f6pi3
UHDAPLn5qVqL3AUFNhevECvjfC49j7i9Se3wVfgzLxa66FPkvlu+ZZhFwxgWWt+n
yQ/ealM7OnNyakGyDA3KiKC7KXubmoK9B8TyYUgXFuRSgRviyN27lm1fnH464ONR
7mH3+m2d03G9NmSzfVKCHOMH2Kvg0Imbves0BWis8SZRRmc2jUbcncPOOxMIXBSD
7PsDn1ERkJa7033mvO+xeS/mfmiHatwrnJfSShDLTCEGjX7e61Ev3Fl/YQjYIex0
FRka9tHvUT4sej9gJbzMi8+qedMvlpdGEy4+G9+X55yaofwufSRUsk/yrsydnJhc
336r0Trs5Y8C5LXIZFyuoTCIsbbt9vksq4VZD7uoX2VhKyB+BbE2dFlXx1J95XOX
4b7/AaEiyt1Ai2RwCWMcHQX6+8PBJHdlx+B5rrtj/bWK6NLLh0V7w4e/MSUhyLOt
k+DImBVn+eFSoyWT7x+ujnI84HDav3OSuvcdQTc/AX3RZ9VljaVptpz4geeQNC1O
QFSuSwlf13rO5wTe9e2DBThA2Cx6qHBV+qCqFZ6fyViQX1t/PD4D8LBH77Zx06MG
m/5AapRTgqzE/rMAW6cud64Ue0uBAXkxN7xVYkklicIDTgB+EIP2kCCmmDIwfJ5j
u0q7gX13lJNT3c0JHzjm/i9XkVENsxVFxkmNunWiLks236DW4zigUVlc+mtT61af
9gQjDB0F6UsZAlzPUeJj0MIJv7yYT2N6ULKoSlsW8I9Mv60CBr0WkEZUzFMxeUeM
tE18EGPxGPF2muto+6d+kRXasbMaTlsRjsY4RkM1LrWUGXiuHmHNcGo6YFrdWALr
k5eqYJS9xd2xbZ+BRapLUJ6VIHhNHf1X2eAlC53PIlUpiqmhhyh2BAFEIba5hWhC
7dx/zAXwBNUUWx5Ux1TLxlGeqXp7ZOQzkcjuK33BOqfEj0FivhQsnQ0h7Q3MOAoq
GheQsuEfY5nM6EE4o/m0pf1hIMJeTfXWLhViy4leh7o1L2fQxOgRTPWpbClu8Gsv
Ak9V7Ue6goHrq8spq7iyq6NwtOeRdo0Os1NCahgZ5ClrGJAOKeuppfyCISb1/rmc
uEa6p81ZjyPksUmcHOFt4ka4jEHYnjPh7cwf/TZmlSL6caDM7mfc08neaR5rYjpv
pX97c3cgc2rm9RvgV54rBXZlPa9rLM68paf8Ynh8FFzO+v7qsgXW2o941EzuAxFP
1rBprPSxgUsouggJe44ydQRtZFntGB8y7Old2TF3kD0OUrvxjXAyyrN1yJYv0JW2
zrmFo4AK64iHQMgKin0r2U5QGcT8xurKSETEvx24lzLWdUANdE3NMlQaV/Lx40q4
zwjEGgrB/+2VUXwoHPDps/vZSNaUsfibunXB/Id16f5OcWyLrG92a+NtVjk4KQnK
K0FSqWrhmbsmdHEeKtPPMAv3JCHqxeUAS7ni1eIbrBIe4hdgJI6Acd9YUEeuBn/c
QkUQlzhYtXwh3UzCernEweRHph1GmN4oMSxhXYuQikbbmfseEidCKVJ+pKU1YBIM
XzOzXfIdCxxjbaT2lByr9jIE+PQHinmGkxfhjE6Wze+jYAH0XrCJ124mUyPu5O+m
1N/9bLVXyT+FmSjQQqQ05CGglvZCkWNdZkZy/Ia5BvHo813Ydv2aa4+3K/yfkXeV
aIbBcAX7OiG25Ocaapw/Pgc8RLixgIWDVxO3dStQb83WAscP/MJRRYfx2MQhZo3D
qU1W4ht9ekFVhwWoVonV2Uy3fmLMMKTxKQUPL/NHrGLgkSggElkLbV9IBbUsaqlJ
Skjke6MUUQMTZj7XUALqEdZozPT1W49vgt5LaiSuZfkxTtTYlijfJEOs/RTW/lfl
ZKbT5bToisVTWHslxET/H90Uaf05pARrxfiJSngpJndw9zwzGuULZQFYsEcqydi6
p10ZFQYbdYlQfjyYtF0ApR//Nq0fm/7DWi0LuDHo7MZZSSYGOULez30j9WoJGmw8
+x+ndjmF2MrlCjH18/695N7jEymG4RKRvAHy5WV9uVGG9xRfJEFYc04hDdLvMvpq
zr2E7gD2YfosK0P+38/2hncjepouFaIhZn+56NwQ8ZoiTQwW2T5NFsf6Ouquq69O
DGcwcA2lnfaGbliWDMm7VZHaHYhfpz2IuI4+zC4v76ZjRLNdfvktiO9PWKb1ZRDi
ctPsI+MGtyuhPXAypyribTYK6z2+Py82V7BZI3aZNOKNZOfH8PJmhiEyK2pi2xwD
0yZi3ksPPuQT05eXXx5hFlmlEILTWuzAfDXYRrf4EQ3dygpgdRZ9L+BkgFKk2/M8
i0wzS6Lze8v9aUYwJIP7mdy/qQvj963J4ENQ3l29xZTtzlP6foFco+fCqkLepHgU
qS9N5rJi84ZAINl+bv89zMDRCSjhn3g7PRmFBFTmiifz+E1N+2Sfsv+yHIFf0p9Q
HxoXOS0a7guh7M+V4Lbk2AKjh+6ynNvavceZwlFtnPPg0HI40k9weRri7d/c+FeH
H71Vxrp0B+RwUCYU4kotQsvMoLfOlkpBVe3igyW76pYj5on4BzWx5ewaeXyEfwsT
6mL+t9t4U/Ad18Ei2z3qieq5AQS2Wcm2ik+QlBCKPbI0/W9z8DYpzhzL9+kF7M4v
KC0REfyhehwfdeA0+7IuipJlp7pXQ+Yo02ysKF7yaZcJryUBhZMeIWnc0UxwtiMi
odjgw29nt371fa3fD8PZkbu+9MEvgt4nLteZ0JL5bOhtdX+hx8UyQIKLbdPxguX+
73hppOsK9WzVSz+FVEXO6naNcwaNHKgtlZZsl+9JV49pYT+DgfvF50RDOCPFDoEC
lxfQUMt2RfqYzadzep3f/gDUj7BX/7e6NduckRQq/9SD+mFxRENWSAHwu4kr58Vp
zA0RtgUg4sR3+1CfffKalyA/GXIiG3mHa6UcouXOpz7OhUeUDfha49IINpG9YqaN
81dNmV/V6I9E9aKuDbQJzTWAHiUHwig/a7lgm+/UX2ftt/1mAKF6+MawRzPjx2Gj
J1Mah9paghrRRP3AneAK699FAzGVckeFC1cx9Aa4p6kDkhLfcxtCD5di3HODOdXB
auyey0NOJBBy6l6SjyVLm7tiCwzJMVwjp4oBr+WUFc9q9SIqmvMAev7DcDQtgqa0
cIkJGAsCUKSRiD0iSx+vaG7RTQJBP7XKJLV0uuEvGePZljdaxLKNJIXljKwVZgFy
OPNVEZ82Qft/3p7xLGA2hSc+XdPAyVLCsrN1gQgkMfZvCohUTvRHUx+eVGZRmwu/
veV6ZjbX86U65rIXVW3dFTQUs9axy1ll1IGvxR6pAimByjYyhTosG047wbxVezUd
IC2irJQDrl0mlSLkOWJZb56nahaxnbICjQmI5DdwoF7PtS5cCg5VdnnRTKcDBOcs
L50FFUp9NzOyrLCPtSwCBN0JC0ZXAQhb3bNemTd7mSeRjz642lorN1qZcBN/398T
PopiSp3av+SAeCbZk5GanNuvD/Wi//ClvQm4tBnJ+9ld6tyF4hDSBjsvGLPknOP7
Piv1p/FjEkv06Bb9wlv031pFgN8IjZx3mBW/N0u8PxQQIkeg7mmnqpAR8tVsd/sg
LFi0+Pkn5fUF43embXH8KwFPPLbgF4vU2eMBh9IMlpL643mYinMp6BerzT/BubMh
x8COqKyCWAoPCc679NGe+fjHOV7FYFQxESSHyJXGNQXEv4vP7nadYhJv5BUrlEav
yQhnmaH28gZleAq0PFQ/BfRJESctdxSbjElQSNpIKPAd0mBSnXfsOcnLSGfVbGup
ao2B/3nhq1fFlCqP+bOw/zO817VIHwP6DiORtaZVcuPnIPnDN19uaCmSQiQTPEUY
/YGobjMQALKyh+LqK4UqPgUsyptWupTaJIQg7GMiUk7sALIspzPAIXt+120dWx0H
w8Rn4T1dUnYWEW6J6n+dyRSM5U0QD7kL2BlDy9I0XF2KeJqX/sQLprlZLyaf+fw8
96NwCPQCvAX2eggsZdddnUtKpxvl2zyrrWmzwlBOlmXzBqer2JZWKAA+QgCmhNOc
wOjJVxxOC3bXsonBiRZM9ycqe0O1GU07k1hj8Fs/Wjglxad2t4w5PwuJgqgrvA1g
uXijSGd/FSXIbMxobMUn70EVnDAza922H3oLB8mvk6DRtp/fnokM2TMcjKhESKNd
AbqD+gfXKGwPJPdmfX23euV0+Qqit1O1LrGefeiM7v64ilLaalW/mQYEvbCJj/Ee
ngCLjBjiCSDAQ5KN5WRreiJwOLxstewngfL83XzeDELuSrxOWqtPDwyzt47nZnN8
DKGpBtDY/KPm5ywTZpPiP/Un8BJOyMuTrtrWUKb/X3lcVR9eRwCH/DcqwQyiLjHN
Gi/LXRMlR5HwRWIyO9t83sfqHJPU/ueO16S7MmXvYqvJsaf9+vPVnzIfjm/RbcIU
UXJhdVE7n1M4dpZX58ctyNcJOecDWXgDYiJ/tKMzPJTMKO7OjIDXAda4oxGSs//I
5eijZYXxBcyTp/UnlpAdQJoRdsNmFneA59QI5E0XjzCjYOjj99tHyy+RKqDQ+9vR
vOCZ9tdiFKx3D5ZvO62zZsRhZRmLUeu3bu5SG60bVKLgqy8TlIVKlgrP5QA6wNEb
wTopo2CbVW1Wr4bVvP4ppVuvPx0a5V+G94KgVwjlIzHnxbEcgYuBm/8wIost8Fpj
t3D0v/n9I7ZcYT9uhJ09NAc5H/r2uo2I4ZLSyTD603oM5rtsMGSIxvE74xUHOtHV
Hw8SwdWZrIMx+Y8AUCOjpigjOd0Dy+8v4n20IELGGaAnDPcueG3uxDs79uXZFOZb
n7sDHwRA1ceyyevLC/Y/79jFA0oW8F/vjcQ7VTMZLr7xWGm8OW5kdeELnFq+VxhS
yfetlCQt0OWDH6M6FHGdx08GA6k8Us/c+ToDMXp2BphWsoqLp2ACCEWV5PnzvmKY
g6OhnVHV2TT5BE5YbbNxoJezuv1ScjnCv3fs0GS4/YIChHcOyr7dtu/zRDklmVbL
dbQtu+Su7GU31z6JZPbEPPY/HILOTSrEd5W8gsukdEov1QnALbtwL54w2Yv9MSwC
2s9yyID3R+c7MqIu4yIKRHazc5sGNV/sYo6kJ4ZDmlCy6PisfYREqg9OCRqqtPap
dNLcEDNnLJVbDdSw6blVTarMPvg0iA5b/n8zo9bRZJWUJgMSI+S2w2LKvgLhiudR
8DZXo2X0D3ZWsOWUqQtsNFChhfIjTSllqluq9RljA2tJ3C9JcNDH/E86N5u7pVOY
vYoMEZEEKQhdVULz7DOXP1nihquYoyp8Yt1M9qW9rxa+H/rChaPjWy8jrjqgFBe4
0o6YEbehgLV62QqYRxwDnCODJ/214hYHm6CT8ZGxmeHuXocc6l/1/YvRVi9VKBSo
DfwOvEvRfnoSEqCvPfO1K3TlRhMJ0C7yD90/BRgFPdpNsG18HgSxN4XI4FepikNS
AY0b01S25H/hjd9TX0mEgC8c2Ceh7N/I+SaEhFMpN1oYn7dqsnr2iykN5VFmjMeI
4fAepRWrL5xROVZ4NRMBlPNq0rfc9V+GnMgxh8pBlqra8iQX51LsUL9VSLgfSPP2
lLYEpmSbSzodt9iOADOW8Z3LFvyM45mvMy9kKKtP1zCO04kCUS1s/ru42ZiPHhX2
eSpL9MQJIi/Xv28/mn0zH4Fub+GSYhJGiSHdgMCW0WnqpKDcPDT8RM568WXLRsCV
7SnE2UiUDzjyf3uih4SokxCr46R+Kx0p0UI6dQIGxPkupVR+aVffTJV6vRF6QcHA
NdgTHIdJMPJKuzwvXTHcP3aqzTctXOlCEnsuLR5xKTPgY9q1XKh4B2Q95sb6CvpH
dEs6cX5vP4eZ31smOrL1ZWQUUhm2awfhMD2BrgJLgy7ljCdjLsqMRdiStuJYuY22
TZSVIqr467OKyCiquyDiFl7dkim6+u7E/RYq56Vv6FMjF9PJFRBrbmvibKhiDVJT
X75qp0+1fZDiUXSVmx612Cf1I+7rTV8GX0dzWqEJN3strUCcycgaWiKhIt463Imm
Pef5xRyU8JPeYRUVvPJTTEzQcABfCHGCc1sQMNNUWZTMbAtlQUthKVKFG8v6HZg3
3wcfu2VuDlaNbHJibikrjmSrY//l03AsDV9iIEdD9ns7LRaQBF7xqx5UtAsTp8Yg
toDyzEBhuGM7mgPZM6egF3Z85BQbDncY0tSjPg2Glife+JvfL8KC2bQdUBP4xDtW
ow2x/o6pX7qhOyi7c29DXgPos8ECtX79EDAmsf8Y6O8u5DsFWRr/DCOeUR5uqlyR
f1ezarKrqpa0pKseVSFAkD0H0ohlwlYy1RcDxo/plIO7av1jzW0Y+rqctnlQXqoN
whLIJ1t2tSlrIZ/g7rv7i/4qfLUlQN3/bXX12dA7QHNE1Qq8QWsxFFcn55o3Mij5
h4UHslof/EaKte20kqPdWgm8Pmx0qRzf2D/sC9qMumjRbU3pDVgINmIKa3seAEli
hcRIoaUVu/WAZ1WcK2CVigHuZQq/oK8GEWToE4MUtETIygCe7Jq8eultEBImwE0V
J/Q/mIrksqiVm49RCHzleYVBsTspJ03hLRAvLy+7f4rtWFxHo0XmAb/rzVwKJx93
/eezyjdsMaGVVlCY64F+IE84Zp/QFLaXTuqclJbTSj6d3TltfU1HLDzVw1EOUXV3
FPg9q7E0oYO7D5rPkOgeXcNidGZiH6bFbiKly09k4tfNgU6fQQZRik/j6hr+GfcX
Ax1ctnV/FG7GNWIuwbNv+cKRP0klCx1/0sOuCZOAkxZEsZ5tLmZZw+CvxRLr9/MS
Rwz4m286Tw89LS5kJoqcYAlwIYxMBdWgy33xa8NaiJE1XNHidI9Gd26BzmQVPjQL
qWgcHdtJu/6UmpwmCi6tBMySR2oklY98FArYUY5q3qB6kmH7+8Ljt+hAs4urkJPC
5DD3gz8uhNs0PsGfopd8ctzOZP9/zXU1IyDIdXA9lxSFDVbt5tIIN/kzaoj1iV7f
0H701muqvByZrh4e55jo7inf3cX1nZL6J7XuNwqJ7ByRNw6QYSlkOObMIhrwQwYZ
vl4WRFj8IonWsEY76JA7kaaus+TL7V7udh1qWQvu74wf/sPQtWWgd/Eb2w9Q9Yat
UuQ6aKVRvE0qpvsxqykvLm4FYP5uiwUDm+HaZuFjFJ/Vlf0DJRWYuB8EoovXzXfs
6rdaqg4o6F9uW/9AYJY11mVNzr4q4kHyInzKH7PHERqKIGQnXpyaaVIVrNQJFVPH
P4ICOTVgnTrcWJEez/qRtoy+mLKpItAShin9XdRnmGYRuXJk6e3yd44f2oYP3guV
MsRiJkpKStmovGgeOZbkzaQd3LjPj8hiTU9WbBvf6plKWMNTb42OICxrZ+wpdhRv
98Ub5sqP1HEc9nUY6pLlPD0nv5bmJcVJll6T8fupi3YR+acUnhIahIo/wHDIcbgE
tdujQ6YsPKJJBNzZziRhRMX2opnsmNqQgpO+LnbUIIn6ZdLvefUnSbP3N+Je5UL9
uWNKXJ8dKc4+EijfjJyorBeq+1HpRbcWZFYwK8by5fFegunuLRHH03pTQUD7xkEW
xTJf98GlE08uhlxaVW+KNnFZM6HJ1Qi5Vts08W/hVIwgNKJOTupEuELxBX7PW0DZ
6kq1WQIcEz+z9HdFgCuI8ML8UriRzCZY/2gzFXKxQYVkWJn7tstD424HlEgOi5d9
6ftkdzyAClgf4LuYGq2IyAo0guN5BABWmLeimZ9DIaRMxEPM4zfRjmjLBFQlkElh
69TtGNt136/UqfvJSlfpJArgWnEYaIwTb2AYhCvia5ktPp2+H0+5ZlUjObYYhRPw
a0a2iDYuh/xFhsqDSbw1Gk8mbi1HCrI3KUOf6AmoKH9xm4LCmtMmOmV3EHVwkDXa
UhVulfX5iZoASRcSzo5Xz3fEH0/AkO8b3g6+otFlLkJKr/Hu9gW09Et9cl7Wf9JZ
wpXmnwcktCJgpl7jm7dkl4erV0r3GU0rft4fkJIrRBlJBjvGQVUJ/tFWT5cLJbpl
lNqPVqyUAHVGMkPwIy5gewa/XIN+e+2dTDz8SNzKbKk2HMjenUi/202/pZgSwkPe
P5WGt91tfyLqWubq6EgUdvoqdqB3xUdE6g46QRdchGIQJbHB2rr4YrqbxyAbZlpc
2j1HDBnTxfO2fNuR0LXmiVu2Yr1O7gYWqzDaQCebywz6hhWRmeceFDuJZgTQovcx
acxMwyrB5Hew45Ye1Qx8y3NMvmLvEp9RGtMY2LoRw4OKyNaRHBCCp9P5x07DpYQU
awVSzNjtRDVrWdal0mZH17YZ2enq0Sm3SCr2k7A3maGcRvd4yEEIyaQOUI+Plg2p
Snu3yoq/Y+tzhRTVz+XAIvrxRO/bn6vc9HJT2wTeEltQRTN/eyww7JqWccweBwAo
xIKKFI0+3VSTK3UHmi7P99dDICF5wk4jbUeTy9tUe4CLCmF/yND+mkn1yphfFyAs
ST8JbwPMPvfq25lsrlumFWFxemYs5XqUUonDqTslo2gGiiZS4gZRuk97btZzieOX
NyrVBVnHoCwpJZzKXtD54zztExxQza5hE90M1x4rB0wl8OiZluGHU6NxvVxXB0op
NDfDPJgYlwWGtvE31adYvyKiCgOHw5If2qC3oUWsRH4S3cJTC0HIfh6h8rVdTWPt
W3OYSl7Sx0YORgXHJ2Xvix/WpoNv0fqXzQKXckEvfHmkVORIR6M/N3fIRqtblJRR
PNlShD2YY1WPuS76+u6t2IxdFsRPWpCZlr5H5fNB778TDvn83ADk/g1uwSNb2iZX
pTrWlivFXYJv/Dt7md9ejMoGbFRlvLl9aWxMxTJZbM91tcQGIHNR7Ow1Xo9SrVPj
qCD3c2YggcDY0+e8/WVDgJiBtapYcOaYKAZGLdtdc4zqAyzTXCxurE1fQNq+0MNS
pK9cJTkbeXrSdSa5pMtHzCXGkiVZNvlPSoBOualGDMD/mX3IHfV3dbyUbCJK3dhq
RgjdXIXQ7yHlSMMeTZClWUkBNO1beMtwrp3T/qOBf5F9Fwlmz54blpJ9hGuIc9cZ
302BduKpdSGLcG7XGfqXeljdiQK8nFCF5VqrskhHI8aK/5aUBmeL2YZJPHt8DM03
XVDoU5TX6NLFOYVtMMZMIHW9oJBVfN4GDSHBZTMB4QZ7nphey8yW6qBWFx9xXFYD
MHKYMWMb6G39LAUq8vm5U9+tM4h4mRsUy0B/Z/UmNc5wZTzlI6OAE9dPMbImgCm1
hUNzRQLBC3cEUfwYcxKXZqCZTZVbhFMsy741g07P4jpFPBEDlVDjJ/uswmCgL1L+
eSKYjdq6CfdgdpH95op3PXynAzHiq58R+2fGeq5yAysTs+4RJlWe5yoSuYOh65Pk
+4bZM+nJ/fqbMKOJOh/SW4HXpRBMnzApUEDVr4uOGQfv7ikWGYplpnu9nD7EujGx
/ToZfRDkyq24PQHgK7BmJ/wmu5Zdp48BnFW2FmmKE+0oQdTmwrX0hhfik2n063//
Csgx9AApghP+c4yb+I/WWpHOgkNxBc1V4JOOy59ppd6sk+BVfJKmgjozPHnRvKw2
Veld9rWgrrg21Ti81rBPh8sVnLUgEJERz/lEokdfeRWhhyl+2bqGSFhXLcCJ3moc
GFpkxOAkO5sl4v59DXvW/Wrc/c+Tp9WB70Q18MoxjNsckTx5HO877Hu1lSl2TTI7
JVSN29nQP7GBYFDA4jdM+um0bc6HggJr5gKTA2SA8lOrGBqU7Q3/YFcZig7MkGnR
W3u+kL7bAaVR0o9IqJjHkf3BXclALljMPe8FTAg20065XO2tiQr8spSXvDm9OhS7
pw7w8ljyvVLKigx4aDLhvwkt1SNC4OOXZwyVcSSf2FWkutd/syI+OiM7Q0aRsDfF
laIAoxtdvUakQRFnMHj+etqHhSVfMUS4FHpeYFRs7MOMIS6qB5XSW0fXXkSZbdXP
wX07PtfdBZj0rHiPMyDbu1oUuoqd7VQLqLujrx3VzM6SUYQlZcnjJm9UXTdUKeiS
JYffxVU9CwY3UHFlvP1I6mqhCzlbSA0xwf8Zza1b1eI879Rms1jxWa3+fNm0eJSm
dEmMAbSZx3bmNwDVZ4127gqlQEIjPjEe5dpgB+ZgLKoP4rZ0dAXKKfFrvZtOTMJq
f+6kx8hKkMIYLhY0fkIjqMyt6pVL8S39fNmZMUrYab4Oepn+A1Rt8ZgH6lXqUZot
nl0yX31tXiqpvPQjiEfgXkVPrZRFAlIlexmtziaKeck1JtvbXXCbyw/Xfhwa80Cm
iaJVnFq76H0bbooAXrbpRcqykvCwH0IivAGg2WukPKDEFaZY5G8gAdkfwtZl68SH
8i+g1D2hycDK7fOOrui0P1KSj8yeAaT5AJtaNxoKHixTntZ375T4Pvy8KwylMa9Z
djbrST4F3+Tulf5GC2vC6F9FvRuI3rOyo6BNSqwTYSvtYY1aTyz7dBMccyxUrsmc
FYWL6FtZHFFDQYWXncX8TAQqt2CZVtozza6cM/MNUkD764YQ/BonZCamowykIZIN
u+DAptSA3Y7z+1zuTB9qEhqYHAxyFyQMtpi6d4MIxMq5EZ0jvTSBexv4YoYTRwsh
G+UJfXeXCWeiUqNciI0VbJwOrufYAuggixpoDIFnIsdE7hiJNAt0kl4PAB1JihD2
9HinPFo0ZbW703TONs8tQVfZEF8hNO/xfU6i581M0MPBVhMYFFK5s58CNjoisX47
kheXjRI/PnuV9lpigSha7elRk+co5MsPIULnx0kTxCVq+sb77rSRidolNgvuILes
HMumhoQ+9iH5kVRf8m/yJ4XSQvjtfMXMksgqmGcvgaN4Lo5eSsKjPbSzn7zmsVR2
yltA7mDXenWEVo2MGuF3nTbW6H2sto6g7+tzxkFQKEVahUJYXIfggzeqpZDpTgMh
xGi1cj68SHc2wDnjq83BqvhTL0C52rbTK7SLyZVCnTsqM/rfboGq00V2Z94PWQhZ
kfWtj46n8qKXthqjo/4HN//ZJFzBBEvWdwKNuDioPZWj4J5RM0MLlzlisL4yTPaB
r9tfGxDqwBK3RgSoPOdKwduDyOmO3mYe+42EY1QZeqUNsOikr1WdTTTHCoU7uQ26
GEtdXEnLR6Yr21x/KKCT1GANMkVPzcw/vHotHtK4sIKAaGgGGpwNPP978bor3Nsh
JWA7jqRdq6ykJ98MzkEyMkCx+sTzQW9A68aPr2DNkSeFJtX7mmaE6rR8S6G+j6yJ
KUW+ZqDrKmKsf5P3TxdpoDP2c0Ipdx8qZI+fpMo1+v9FjmJPDjauarT2KGYYNeic
OZbBEFwZieHEH3hhzPJBP9gRd5egGHs4TZW2ThWSP/5ssRRbOi+vlOukW/uwnwTN
yYgnISvlmaZcQjuUd/4ulN/bi4RLZ8owzOzvQce0ewnceULqyMTOboLK1zNbDLla
aSzoK1m1asOjYKGmw59IeZJVICm87AHKQGsaQx69TlfpgdyrwMZoQ1eflbcdHlK/
RfwMowofFUzDvdj96nsQJV3Db7wzO6C21sUBfD9evJkU7uEAzBgAfpOgxjmLBWU2
BFyG5jQdXjTnhxUYmguHMbHkgEwW+GmlwKutJTBOGEI5XaHXBQCNYcbLN9xjF1FV
4mb3cm4TRrsQ6xq2S3i3hmP/Z1cuth8dgSSNkaKSEZJvVXrA1pwYNUccLznhY117
YjaMAFBBwNfRHFMJL0rEA7PiWAOg5y9c4a7Zi64LUtUUuA44HdvTU+OiT2UvQBMY
xaLJ7KdUAOqHl5GguKKv87JoKLsdeXmzJspdEVy03s5UH2vNgLhFgjVJQOg4FAoP
c704okzn+Nxl4gYldlt3cABYGzAClU7EaCOiKnDL/0GFPwgR9c9kAwpnRvLBKwgn
bm1fK+TK12V6rtRENy+jB/yX7II5ukshsrQuZPt4K6s6eMBoiWzrCPFn1rOWrPzE
Z3+ewVLl7VIP7C5rVQaLf2dVGPgNka05rVCEvYkjhp5jOs3RkwPEX3kJsTMLyDXt
m1Z9G01aw32xMmZA5ntxV3dsDjOrhMdnJjdOGZRtFxFJ42wqb/HMHR022T80OdcH
LYrg/yV5MRywVpr92J1TyjBo85ql3jKgAG0wArcQO2CH13uy6KosjpYmnX59OVA9
WgwbOaidJvb2eh4dQbKF/YK+56JaicvIc1nSvH2O0my+ErsZPfrJfVNMFQ/zX/hG
Taecx9kvb0c5EtcsJhomFTeUjxGoxl980Xs+YprL9UpOxOtmm0WOnLfKlWvrr2/M
jihWcc1ieEQ7OLdnZI2bMQggH1ibuHZNwafD7ypF4oWUPuzrP/gOUO1g2tvF2z4i
upr4YgFOiodTNBS4yevv9cXOj9LUr5Va7tnT6AzW/UJS3mVoUMmBeq8SpInUbATV
Pi6bsBIfVrWScjm6AhXDCVepEjUJ4n3DcXd2tClsWK6GBAnmywd8egO1U3RT3iir
5q4PBCfZYc68txVkE1XkonfhUAkrA0NxP6BF5ObivDJQxvhf1CkmPXQQuDzmop/4
kbbFiUpG02VeHYVdGgNTNiXAg2K72fawc6CPm9xOHA08PzUOfnEY3KahtwnyqZ87
c0YESIW12cGrbJD1OvgRWHcxEtkuancwi4ssk3xHL0rTJDA0bC2tzm1fYJp8O21f
HUAwoCqTVFVTgZcamh4DsrgWTM0wiNaIoGUtdDoN59kRaHWbIIPd6tbEzuo6KBwv
0eakAEpjGF4I3SgSky+QuPnZJKo+sOlEKwpBEbMikrW4xAwX2XnBrlR27Wwv+pxw
vPEi794dlIaP1dh5f1CXS5uCtzC10BXxNMLPo1hnD5PyGMQu0WaBqfvDeob54VN2
WpgSfp9U0Ua51ZGHWHMsAdolPmT7iAkhvJPkbMbtXq2sJyCZq1lF3/lnNmni4wVX
So1+vYSyoPWm3C2l6pjBy+fX+2YyWX3N54Ve8I5EOa3L54282y55OX+uwE40472g
pI1QbfpUfawsNkPXsaKo1I0vchGk4HblxwSKKaHMd3R/NGpsuyQl3KtQHijjq3rp
mGhqjRKSqByfO3MVZBovcd/wu85LnSPISW4RXSuQf2Kfvrc3Yu2FVpfRMYGtwLsh
sFrWSpTh4n0kzRhPPPhH6C5cZB+Uh+BdNSP2xaD1upiUSGfqDPiXV2oqLo2rukgY
ZJVWgAVmVzyQJ+nBufMTdpvH/hSnmv1twQz0gKW2O+8bkc15i8FCzPu5sNbARvcm
iffMk4wGUqDkQvnzYVQR1rB6R7DP1RBP2e9Z6YFX62NbFXVha5WT8NUYdyMqrJkC
TRGIBfYBXMkfzteCYFeqy5ov+KbmnjgHUUtTljO1ThrznnvWnoGpq/ZkDapFMnz3
dMvBnEj5zniinrlPKQxckIkUslVIGRUKTUmQqVWWsJTcsgQg8Xh1ADW6pWxWoLhg
UKhsvbSNEslKWvxyK0CIsyfU0QqEMFrG+JSjp0/9dR6Qkgjw6Mg8HZ0fzAUsScXP
Ejdg7uXGjrMBpC+dM4kKa28C9IleG0y0ATi/UZqhTiVFcrNe4ZIcX2F0eMV3tA4i
ed9RnFOUtAx4Cxx0MaBQhNGLj4H3B7xvSpZDWD3Wcq0QrgPq3jW/cIq4YfJ6i5W/
EPotUyA0GiT0yT5J/CtORVahEgg4sPfOSel80b/gb7kyYqqY5VqlYGjd62Yb31Vy
gGdot0oWxyzTK5/q1I0cm4j6RmEUSSB5gE7uLEf7U4HJjfdnO2vRrCSxtFI74B1L
A3CsUCUcTodLcr70jvzv8RF4za5l9h2sk/i6PupIJpuXgnBHjpjKr8RRItl960d5
BlqGEEcswwYVir/Z5yhJKkpfyR9CrUjuqoZ45ZMt9hfJ2vuTJEbLao1sx+iMkO5m
zS+SXb/mgplSQONLtOjLykSDU0ypJYI7cIF0XKN20W9+olpmXrhbAOmFuyxrSEJo
1rwGEG2vzM4n6sAvlj2Jef3emPNEJ90vq3xuKTV+jHTYStXdce7Jmtqr6eDyptPB
SnxXTppBk7rnDFOKqYpArEVLKWE4hxtJdlzNfHfoccivOyExRbGvNeC16cTgHjtu
rkjAHB2ZX5QwIg/MHmvCRpt0nWRf+i2UYkejoroJV5ebCUAMDUkevJk9eTuJJW1f
bfV7j1DBGyBcjHPAwd1rUb5u++gvh/9VGckaruJqy0LitHwYg8xkLYkFzKQb9Bu9
Vpv1OhUhJBCGji33pil7FZvmWD3VLVPK0jtK9DGxckf/9afmEnLXBZ+PAhuKQEMU
N9MHz3ZKvvoXhhi6HCB8dZq+DTylT94mPMAFU2tbTmzmMnfdMKyyo9iE8JJXFqUk
tplYaIcsOlLR6wx8FVthcHaDjeU7bgd3gmDP6mmTDDHZGi/t/Zctq6mG9YiRnmq7
x/ed1vQXc01PRzeDKRsy6FcfiQh5npiS/aE81DL9cfIobsB3twJ1cWbkt6wRIFO7
jFBRiq2BZKynhWCFy0aaJHreTmGHACqyqaB+0nhhmwcDnPg7EWiCjswDBfzc8uW1
dOuiIPegcRV2vB2Mm0BwXEWpxDNV4r8EHhiCvkALfvuiIwooAgeUQ8vbmV8SYMOJ
4/pvEv9FATX8uOty0FlvAdmAPVP9cz73j16OIrYVnxgZQQlJx+BBZHkdLFqm71XI
nU98aobCWK166CSvoLBOLob6n32LmVPQoFqgaTWgbxKKrAtvLOpc1V0hqOqpKBbQ
+nGPpSpkS5ouua5mKPzlL4lX86WE+u5sm/zHUm8YBNuecbdCBoWq1Q4WyLkyAsj4
dtKf5uFrLJl3cRWM44cTEafvyLwpqit+8hbXDa3xqSNoF06cgFzyGIp++HeTuLlg
LBmbYeLsnuN9YUvZDexRYVrOgxVgxBUA+ShzKahf1bEJxoX2lsGecleParAZ/Ntp
KDZL9D40Vw0b51U9mjWx6cX4RbaJszQ1O4IfjOwFrhSo16cK5KXKB66fpIFUAUWX
HXoG6SHkG3Yp/xlMqe+bEOC14JPuDXcu2G2aNa+5NiGrRfn8BM+3wlkXLFChPgKd
nGA1bkZACNhulo1BMugdeQSVU+PZogYnR1BO9Zitepwa5XqHQTmhorwbK2k86NRW
YFpZB8V7bbLynXbPdOxEvvkq6kGMu4k/fP7f27uH3JVnQZvnK0AnZLdh8V9ewh2R
J3gcz6CocVQAhEGH8EeqcHhRk7ileajUUr3MXjWkwnC5eYZu5kaL2vlvCzd62PJd
qUMVA7If5UDW0+2ZR1Q1pR3fL+0o/Iik+MRn6CrJzM020TGsIVb6JaCiRfb1BBuY
TNnH1xtUYkg30FL83foM77wfF8ANrHKz3nAq104452nrJ4NyZl+Fvv9lqebbJee9
+lsZTkg9awO40IrH3p7nn9Ax+a/ch4Sv6/7kOb/ltOj2opL6Yic2sg7Dwd+TRvLX
bvCVVaEFbMBNR/xb6/rAYoCinB4aNIeJD7v9v8DZWU80LO1caLF4hP+BZR+/T2rv
cAMAgmBSIm+P01OZLTZh9wcQdD7wK1ypfS1vdVUf4DZ5Xt5nqrLBkjzSlB6GTCJq
V5fW8eep/psv1a+ATjaf6Khd0a7LiVn3kO751x3JxGE1GDA3E9DX69RLTdUEP/GB
A+0PQM+pLLpLz1znk8/lg1AxEZw4pdHIu6NOYvBJpg0WI3NLAnGNdSRVlqLzBqO2
4XL8ydUuwytWbK3rRexX9BGE/ILWNaLhcEYjLAlk77p0HwWO/rgLWDmlkE2U3oib
YBp6zEF3u/9FnzEuzSMx2FD3gRSW7G++UVEiJXzFjvyd31kMVLN4+8s2CNvK0Ych
HKBrE5wS8lpfO6lWrNwugvC/dIsNieG3wJta9lqm0MgL5g7r4KH+7r+2MT6vVcK6
0zY3fb11jC8UtqfeklvdRrXD8ydI8kmI+70c+Ip7hKtgUqAUWmg4EDMB3r/ex3DX
ZwFzTq1LtU3Df4/jVVxXeittD/RPazE1sZAkPF2n+NOyYIifFAB1qxSn9AjYmbLF
yTF2ft2mcXL2LQjiBbcwSN2mka54WR3aG7v+D6/+JlFd5+tVn995+Mygfs1QdJUK
EFtJ3N6Rq1lv4+0vqJMO2n5mS6ScAKX7vf5pLfz061mBnBYzqn36SGoJeMKa1Qz1
0EyhDon8FgLDAIuX3W5CohwlQjyp+y7Loxreh+o4+aybpO/NHo+fGwewZRpq9kNv
5zDdb/hnVx+G/NbRMdDd++NIkHOAhaHLn1zjN6Fnwuvb+JysXQuyFWtcXDAgJP1q
CNCuPgNqP/yTjfvGZOmWw4vytSCh9D4rq7yFGowxpHRNlmSvj5pHfFHSudcSZZak
vjdsRXyTOrC1Al4NJ9T46hRO9jtXTKVmrYqLy/LOrRYTYo79qNofrEmved/DYmjD
iEr9v9xmdiwFAomvounZp3z1jrhQyAqud3xdM8Ljb9RrPivwsOpYD5PqtrBiIpnH
HuhR3TiZweDildTnSogSwpzACIZhpDBo4fqRCFMo+fcYYxBSk6VPjfQGRcWjMqEW
XyD4SVsvErmdJCzAzkZDMiVAJlbDrz8pbHFK3lp53Jfm7xXxm8F1ns3BbJ2Agq6i
BanmXLipu3aTgg4j5ox889+1WiXAGNc2ZN/3kd9c/jOczHC5qfoTAEuNBRsQ2UK7
EENOWkdNPAVIyQOkQIl50NUqd0nOdXcdI64vOYnHsBNxz9QqG7m0XSvJjbICjoof
JXjnX++L/Tbww59rXzqxQieoUEsmr40Xt6BLRgwCSnDRgEhTN1lHUBJhhIjslWDE
+DPzCJvcg//hqr750Jh37LyOLv7aov9HYUY+71MOIyvvNhcuwjKKtjPLJYJkf3sb
fGaDhi9/pAlgAte9w8ymXeJHGDLqRG8MnajBiD+PwqnnFW9BAfLTSibDVDQvdjnN
zufmM4/XPpmxKVOdTGVaJONUE68TtLSZ8FjLkQo92WerYHIknuSnd2g2YC0qK2hq
hWP9s5TN26FGjr/7/dp05nmjVGgVveEyQI5w3NqrQBmtBOw7Z10wopbhKZ6n84a/
lsFX+g4dwoYhWOE8N0O8oGyk+dB149CHX4tVJiUqDn1JO1/hXmqs9SJGzEBMgZIR
WxJwAd5OgNzEnzja+u6KnPxYQnvLYh7VnCjQIBGRyBjWG7VEsvXkln9j6OEaVIzz
h+ssBosJgC+VedesJwRVGp8Hrc1Ckt3FJHoqZcwHP9sUovWY5+7vL/ghdkA7Emx4
Afl/6CfWOxV39z9ZSnHZOJw1yK+/GYMSJt0nPZEV5QdXSDmaeO3J9kS+CqUa7i0G
3bRBnzaatPRXd6hwBuZqXA2FdyOR2MbDnGb8UPGP16r4YO+TpYEBk+DQkDcLFYq4
zWX+YCbgTToTEK/A3qRxLKPjdzimDKVzyln93s1quJZlkwGGSHjolhDGk7Q0QrYV
MwRBqXwif5Zt8eTPJAOhQHLAuidsheg7Ik+F5tzfxm1jpZgIia/pdkG4jIiwFs16
UMZ7da72ZNRGoY8RJrZM3UDHN5rQMSlz1UKLGbwE8mbHm2h8MTiWQkDKe6dD1Tu6
m+wWp5xJ744+ghWsO6Uj3shEmWGM4SeQ/b4wuTnKv/P53RRiHklwHTYxMUNs9Kox
aTcDIb/qZKhjragiUyC3V9wjGU33IHpf++HjtXNoV3MyqRto1pDDF35jrt+v4wLa
eLDmPcKGndXtFudl5TcK6O6afc+w58assie/qllD1X11xdGOoOK5lK2G30ftnNTK
2A7BU+b/t0aiEOKTxcGSr1K/McjdfS6D31rsBI2vVFqkyGRpdpRgD1hayoapQmet
C8ZGLPQL8QrEhCSa3xdDWnTXcF7j9AjlTwq0mjDVW9F2LXtlSY8D/J2k1J91u9Td
v0kWgVWx0of0cELeIXB45xZp7HWLjTITC6iIoVY5toJXsfcbq1IRzUckNe+IBcDQ
OmwudUKlVQqkO5VZ9cMIVsBl9BxtdYwNq4uxhZeLY8odsS3Lg4IAhJK5Hi8QZzX/
z3DtZG4VFBamN+KY2oT+/wFiuOi4Fr1XckptzcmngzzEgFQnnNGybZLdI5TiLcva
SwbKRmB5il/wY9+2k6DJzgGjcd3hPpI6oIwAudn1SSbhh+X3S+NHGpc92hSZEPzj
RzKJRQ4WI+qzG6bGoavCZm3xSn+mVstH2PiAPUG/EDLTffO2AwF3R016V+vwLGBR
a60L8vCw0NTvJE5mLwv4Mm4xcBssG0rOHDGOd5jHeJx1Es4TQYI3rNEblyraU0ua
t74jOvmZcvGO2bRccF1zaNEiS4wxMsQc57LbyZA0+qXc9lsgE54xQ1++l0Q+qsIZ
w/GROL+TS1NDPFkcSlZY/bOSnQDs4/ZMPH5hakaSd9mjDUiOqbko0M5cwlSKBbim
SvlOwKp0L4F55yjOtUlRbZUTAO3AISYcHpLPJol49bagbD4W9birUZfx6ndQuWzN
IgXEqrAoDpPBt/T2L6Oe5leaDpW73lywFhj+RifM6tzN6uWfIRY3lIZ9Gy5Hb7CE
ecrdbEDJpos6/gthMJqVCh7nwca+JmHM6iczHYnHmrocn5lLNx91J3JS4WcuXOe9
ZeNnfq6KjlGVAWX+37xdk1wa7xmgbX28y+6wrs643s2IVFKqO4fDIyokiIS1jUpv
OFmdJ8FdbRjuPFwYBXkj8zvn8joD6GRxGl7Spls0bq3+aDHhqSZ4pwV/iA49apO1
y8as1e+XHz4hfc7mbTX1lepnXLnmslyfWQ6qRL0OUvHJrHVU13GvHRsOYFQzM5zZ
kSM44ktFzDZrZOq4o7yVqXGGwh64jT0u24CZju3hUAN/38XpTkEiYQcUcifDvE8h
hpIYJ/FOe+f+iU1oP6STqum0aSkXeBuo1nNIiZGFy7RngaaMDZYfyIvLWO+6tDCd
duiEryPN6fRz4FjTYc3L9c9WrT8I31fazc/ZR3XxOYHzbi96/rPLiA9tS04lsjMj
a78Tkt0v6jkWCdfNEVUVgI4UI72REruC091t/erR6wklSEEdRF3oWw5MgClWXaly
mCcPj9GrXnxG4lo/hpRRaWilSfwX5cjd1s75fzJrDj9AslkZAIxwudiIzvd5wwVO
o7D9jQsqNy+avUhvixj2rWyMJrFN8hz95W45pYgg595BCGtvfbflzpRIeuL+aT8n
F/B5MDJQ9Njv3/825OL6nYpAs8i6tk7k4/oaBEhMCIuy2fY7xNr7G6krgGTpofHI
9Dz9/t3TvQsSodJTe8CyT7IRQmoiMaR3GMQjvH8jRXhWFwGTd4ksBOZIPVUG/Nv0
Jx/TYovALg4BhRRRwH5d7jjD1vs0Fzm77rrhMcC27H+0PkS6NsZsBj98LlqJZR9W
sTms9PuTiU3cJf0QMPkf7si2dLfUGY0/hhMVyTxSv9gy0FKhU+r8Srgl60XNNXs5
JQ4Y395kzXldDQkTKM6IhpcXosc0mgLZm1IhErRuSapXn/Ft8Jk0Vk33sGY3mtqS
OCHNLbpd4VZ6mVhQG2C+H9gL+QLaVKrJmQ8Fu12ZiQODmzCVuYSEZZf2pxUa+J4J
zcg4dydHQd9XtHml72js0H8H1dzVnURh+M0iOVXlNv4LXEjgbZ+icnlQdE8b79Pe
ksNh0eL33yzzdT26/6AiDDm8FPAB1nThMWBppytQ38lzp5h47sY3lQM0K9t7wje6
Zs9hGLCiaL1JeaFDjH76pX+jd4zAPv48/p/Gbol+V6oOQzAvtg8Fltfx1ix4HmcH
0gQ9uquc0O7m/c7pvUqU2/vWepVcCitQC3/w8Sl+mVRXRG8TqVLC5ltqEAm241sj
7HuOHdR2TuMnRgVNewUPwLS7vr/PzSKogisjZz+LyK6FB2NnP4tCHsgqYwpSiLEC
hRJk2DsC7I4uOOaw+8Iwu9mXPLlOOkTxSc2JfgFw87NxbGoQAAxtdWHsBZIg9Zt/
iEmpBKSLWRNu37G3ydQXOOL7f9uHLxUQSSaU9sXUSo68GXHJRAEy/T9pWMmQBPLG
jBqZhYxE+Sl7gM+FneUNWKwf18rFc4ykLweKkKF+/tEMNoMpi9jhSMfpNi/vMO8Y
+me6JNmjkHgbSu0kM51hgSHhqCfbaTjpLs+HEAyzffBwY+VBxQ+b2y766/gr1wNj
kXVJqZs+xWt9fQX96fOKDmwHPAuz4j4aClJxj/syLkB1EPk5k684atkIt3llL8cH
QJegY2fF5Ae4KJkePMPpPHZFIZsnWq1Z/wlza3xICLpBVxEyRUXa5Qp+Dx6Fya3j
n2za9mCqyaOmlO5jyIUw3/t0lCNYYcUFLKKPZH6TD1wmFMSxWZjtQl1h+01RSE7i
GxzdFbAseksM+aiyDrK6kqNXSgVm2aB9Z0jwyTsepgblzMjG0z8+1yQn6ab2Uvk8
oofAWaRtfBkxlq13nY5qElM4ta8Yi6YjF0wWg6W/IVwurtvCywnkclQWAOxCrvHm
aZv7itGJNyPJ0vWrGFY8m9e+/qITet/+XxG2RA3KQ7C0TPdNzFMBdpK4Fa9kWGGg
tL2HLPzw77Y7cU4TCLAh7wGHqlSneVy3tvWmPpkMayY+dLCz5gH7x6J6l7y3kEbw
lXR5dHaECqZoSnG1gwhAIplh1Qh0WmmVcOHH3Qw/PWtPKk77OBhpTuDwtbmrbCmT
LEA6NU8uTfilZt0S+q/Nit1iUWeOdQezVUtUAeV8KLG7yA+MC32NJYaoR8vuAsU3
0WDL0v3QY2g3a4NvBMqZgVgWtqUuUQ+MCl3/Q00OuNSInKP6fIBrArk5tF+5Y27a
ipkOlilfUtr+QqOz7KSxT2vVcHSP2t8mtPdryDvIl+KWD39HY5nYLNR86TqHo1Rn
ESXZt3Zc0X9kUsFA8+C9dmEZ4ahRMdpcicQignoXXRwuPG8XCT+ynkIWWZJbHojQ
8QYne3zdGbANhZ6T48H3qU11f7J7BqUciKcPD2p6Ee0fkQFovYJYrSYfvvsdXEoj
6Rb1twiZS1HQ7bRtTy5Jg4+P3dQaRQATvqUTiErA2pNcrtBpOuqVHJAF9rf87NWC
FVTz5X4c1EOlaEC6f/tA1/+wHOJVbmZfH7k5R1Ql/ZBWbqU6s7Sjw0tgy6OMmSF1
bmwgNk1ZeEhw5DQT1b9/bmnEFRorMPJr5YbmA/x+kvpF5Q8msbyRUZpgVGt6b+SM
QYKWRtrSOxTpPdtMTp1NI6Z8geMdpPaC6JaHc7k+y71/gfhtoQiataW+91woJPz9
FZkW9if23YfSey/ABmzgM5ZyvU3z16libayVHvZPce6zS3vDdnALMBeRh8zwlHLt
231roDhGUPjTakxykC8Emilxr4SrrSutOOdnEuw9bsyoR0PGLYWWbkzYLR62q58R
1byvIvA2YFNhISceNuHzXUdosQi1hHHk3APY3ppSnfwNJR9kxtpQg91kPCfHOrNF
0/b0zgs4g/omUcpHL2UbpgCtDyANs0NakDl56UV51c6AMlwAdL4iwgFL1DUvxnN+
XYMD0hggv0VpvDTrPeW6F1F31fKVS27+JWXIWOAE4zzUkmqsYZluVNWj7ZDpEFAA
SW26kbSqxiwIAhVm3NZHdq68FOBxW5UutILYkG6Q2FUdrShjmgeZhxn4XFMUgIor
jc+ZXbo3ehZ/uMFzoGxLp4fyo+A2fOl5O6nYF6t08QYTpLmqWSZKOz4oSHcaYuKW
AVF9U2UoaGlnWglKYTGFCppijf24ibFr9bJ5B/kHC14/vT7ep4PSw3VKYmfayLhm
9YZDJLrXI3TWDTOy3n+LXqwp+URT2CTC5N79REAy9NTAu29sYCjJp8YfD/Z37GJW
Dt/v7Odb9aHPelPcS0TSOmKjORQem+PHt+k+fCGUBCwCJEwDEyPeo8h4sRmX7xh1
qAPR/TxRei8dlokzFs002Y+Fyzwypw7KW7yccxcSA0KVjMLpeSBJ6Pwzs1vsLlVU
Vugvu0dlmmNf/xDsE1c9AWZAbSenNFzfqTkKQeGJAHg7VHMQ7X8F0EP5yPxmLH19
rS+lnXHHICZXffFaFL+dCES3ojGT5sRHB7DW21WEVH3hLFzHrIHPHqON9nsibvf7
9RfUUZr+akYeH9nWO5KqMhzmuF7ECLaf0gPV2H9gj4kn8NVIK1toiF50wCy4gbMG
dSxNyoa+hk5RvaQbyVEwdGIhNsPTtk3xUYEZAfIbd04mlrgFfknjwLWW0qX9kFyS
DMgmcER4sVoQEV/FbDEap4lv7lSTxVHc66206rAumf1p0afCh2b2ER/3VcXN+1ca
vzbs8947uLTc/Le7srkA6hpxYkm8EfmV/4zAkjH/t0D8EudQb03S7yz7Zc750R7n
h+qxNkAp9sIFHNF/CUHhEMXNIe89Hf1MoILRfqfu4FZV+wOHNmDJkopMVHSxLm19
XKhAa/FENT4q8pfLl3TTvHFfs+zAMy0z8MF8CQnyEMtrJknABDuoiInD9Oj1d1zw
3w27URl95sHx7sS19mNBAEmY4Ts8Mo9uyYcwkQDPZiFHeKn8HOW7QGnvk0N4V2el
xB9Zmgav+kwsSPfiAtYsIF8TH9lr+Bc2Q2l0XYxrWm2k/dgAkKzNyN4EKsoOeVrQ
Zsw1PDIv8AMcUHGXQCNDHjAuteoSkMMVhfPcIg5a9WqAv1SsZCKjdi52AhuaUr6s
yp2XskQFQrSFhXQO/fLNeWfi08rboebGEk2rl7Y5nk4N8z7Ew03vH0sP3GC0SP+R
k1T6pQvwNR/n+2LrxcpXOJ5+z0OBd5rKhtwg7FVM8E4SZ9LZ6epncAov+jxra5OL
Dir+3yTk33casyPkwejvCW8ge/CsmyVyViNanIiEMtWup0sKETxLIg/9Rji6WNUY
EyX3dwlwUHaXY5MWSPkB4H9LP7z2ws8+8IRr2d0/zhdefikAa+g8y+3QH2s6u68g
N8AQe2EW74qr8JRSFnNBxrTNLAWxHbX+hi7l+hAykho3gVw+QvEW2uE58z3bN9iC
e9ivA2yV2nU6mOb0DpsdCuyPkPojbokAVthsKFqYui+OrVzKB1R48ElGnhS+zTt7
ttdBv91jQ3+r86oAl8+lzvmmi/MLWALEvOePcBZlXdLR85/npFvll4k0fo/xndWh
ubzGDXjGazp0K71zatrSdAZ0OLUXX+PA/nAVJr1lVGfbfvySyuPwZNUyDKK+55dg
MOxaO8qD3lXGz/B0yOr0ZHA5MfbPIr5m67jyJH3cjyttVrKNZLYCZg+sEy6NdCbu
NIBkf7G8/UB4RD7eWnnfbQR0Pm+JJo+Xit5a3hbh1RTR12Pk/1NOI8yKxb4AXwPx
IM17Dd321kweanU5NTP7rtvlAUJTK96iXELXf8jClsoVT4u6V6u7ZssVtTGp6Ehb
q+8zxyl85995fofG9TUj6W8c5jAcHG4fEQcsfDntraPRb3M4PuAfhtgADfN8dGeG
gtIA6qLgrTVC7IzNj+zLjpnb9+Ra9bhFKWgym9qGsnaNWHIg5x7HVyjctCP4C48r
fqcwM2+bTXEFYv25S3XC+pXsRWRLjaniWZUWFl2zyiAddjRihoxP312YnkZIlOhn
l6mcP6vY7D8kWC+wIAAmG3mKAFkF6HQdtNUXlsnQ2X9hZLeKX5k1TijhIXGcOBy0
MHd9ixQWlJdGOinCOZbBrhKi75RAsktUoJk8U3BZEXd37g/XXvlHg4RvbjlWKJQR
7LaUZ0sAAF+jHFOKtzS3XFcjMHbcntFoslHYCeVgAuZTcuka0Th05oT0vBy+brao
TjZLdt9ijhzSz4OQRSSEWGs7kTDYCRg4ogH8AZ2JhHShN+iy7/3785HmkBc6MLvQ
QB88nL33/ZM2ROcKWvkmW3XE14aFhbRUfbKXBjZ5Hw1Hzg29ZWgYK/QqRd7XR8F3
tAzeKDcU20y+LkrtQhoMzOzmSwVWuVzZu3VMsLzFZCYuQaAkoXyXqr6Y2aqxCZHf
bt4tE7bscC8HSOUjN0F3wMOsxLvEyp5BKh9OJALHTIYw9852fT70wk+vwab/sqMW
OUa6luOWKCUo3Ffq4T6RjeVQh2OcGSfJb9DCTDIATVwNO68rKZeAFkNoptaMIVDu
TmgiJdVPyN7AXm4Y3Tq4PdWeXlcrkeU/b3jgYRs93colUOllmwqXAalP6UryygWi
NchAWxDTZVg42CpDykYbiLhY6T76BjH7bUyonKDEu/mL+dSu0X8+BQXlUH/Vae+s
3akgH2yS7oeu1cxC/8iGxeo7k7dFAEvy8+Kq/ceIaP7PxiWu4F5qXwC9Q6fKF+KW
jZG51uA4gPGq7U3jGkJIgHAQWJIVMS750X94Wfn7vRubSvmRoWLV7pImB+kgcN6w
xIXaCIM/GdkWKvcF7tIogNFMCLoNKwLOn+aBsCOdfo3ELsWtJRo1HCnyPQzBsgwA
i9w4tSTIoLXSje3lBXS9Ms1fQwwbZcx5TDlYs0z5Ius7nr1GfCXaInW6cN7t791T
XzMQA4R4gwLVQzHst7He29QPAsXM3MGAcho40j4PhApvckWlDeHmuT54Eez5iimK
2KDp03dz//Gn5XtLh6OiL86D6Hkp+YlCK+bWUam8Ist2D7PZBjvyd4Q9QSp/FvWt
D6gOWEyUazyWtjrcS5TH2jcKYspGsYTJ+fY5TDD3gwstJdXNYCGXrcM5nyxKQc1R
flsyOMwZjC1H5P8gVcqBxffmNn5+GnB2quPss2laPV40/Ddf0Nx3kcqRy5IAn9Zc
T84xNRY9no3Bv6ZuST4REnEH8IWSbug0ghq1EZJxhUINyKRolcaA0gf7GoPcYEVy
58oHHKOqRMyrucqOEgkFPif8SMXqqMLd6EKWDD429MQ6Bo1kkUpKeKq0YeN/u6b0
qf6Jcf6MDaT9SR7NhWdUdWxjK7E/hqmw0lKGfQ6O2ivsYcdmtPhrFrAVAQ2TbqkE
QGHa170CVAf8hJEKqhDhmRq3ZUcs76hCFcJqv0zg4XK/uTaYqdwV1I2aACrSEIIa
tVQkc14MMGDB/sasV5owgJCfXTDAzhn/ndasabMSjJcDraCSCXIp8OMiYCe8d9MV
zqqIHb8hpeBuHA/vs2BYmzgYYceS32A9IpOv1K+t67w8Jg9rxoio5KOjRtwWRzZH
O8wHayao8Y93pXKSareGfwY+bEFrNyiI+fbzb6v3wBelFpldSbQ0XnHWSZwFgHWo
lKVzcCGrG1EJL0QXjr7dHwzDtudrMZVt8zl+Rs9eaxwIHDPd56obw5WPami7wdJt
3PpI00jIMH46JTMYO7lHzrBKHHqXGwIL/a5OA8E6ZgzDuaqvlLwHXvC//9xKPEsw
gKUkY7VKsO4IQtXQzx+mOTMqIzoATOOj2a4lgtjbypAwvbsb53lu/WFw9Y3JhLIr
ekpDeZMJw908C6nAbian+r+9JmLweOe5lcRqNWnHrTQdcMdOW1gHorRcfQjGNErx
lqU/vZxjKZ1t7JGhiDjCp4gcYSFg5NU2c6dugYLrB+mmd+X54mtAE+yqE6WpFEEW
icaUktbPVX9uGJBf4Ly3tNr04zEolV3iLBb6BdiibQDQxV+1swR6ROKIShIl35SR
RqUVObXL2dLq7nRCUoP86zFMrVj0QloiDw+isRshrRgQD1IqvnsGIX4Hxrw4U/TC
1gEOJtHwI6h0Nh6KusISx+pyrFJU6vTeJ5VmBzfkRVH9d2rk+OMQstyqxeasatoB
63cEzkiIiU/UdCNNwUx4qTanZKUNuWYwbwAllbAhcFWCj1YXQD7l+Hv5uoWh+1/d
gNDEjyUx1VCzuisHbvvEpTIGQhYuiZy7ZAHsaM4aB7dywBXBIiuG46b+MtW2XSL2
9BtBOTeCiKBS0YsQZsuRx4Rxpw/d0Ejr5l+52KHsI40EzPRc7YsPA1+KV1z2NeQH
/uaDrGqcrn+QATb9+Ht9Wi+Ud0cyTC0RH5Uz7X3T2pqgC0kiWtknMFT5ic9jC2k+
X0in9KSKcicG7JXP5YZ4BKTgPvsJbHPTPYGUgxsiGslGjdVjGomfLvr/dTf0gpLU
fktc7V3jFZF+uVrEeQamglYnbDo1noffSnF4cyRKkaRfr4hpHwzHW1bfz6xzE/I7
kcxx/Ku0f+3szkW9Pltl8gX5+MvLGKAzzR7C4zCZpbVzeyzOwBcKoar7zrrT5E1v
l3ucJLmJh50RkUIFofmQ8g5BYE4jD6ClQc5lxwdkitMdkZDpyN+XLbRqzZdjs4yr
3IqjhCcbWgiBgUxIt3V7vvq6BpDvG1wDfk54O4FK0Zel4DTetAGhfn1FGfibbVan
htRC6V+aM4rZNaQrrbcd+k6se1usGOYhh6iKyVdg9bJHeIq9gdZhsuCF82/fY0NV
4gu/t9/DQBbM3rW0y9gKq6lyLI9DDY4BcOUn0+Ly1WIc6Trv2SwLWc32649dQoGs
DKj/B7Mc7TAFtjlBPcV1e/YoMs3qDfCgbNmCpWYOdwICn012HjhbXPDm9XwwgkfT
ET+rBcB7EZnwKiGaKa+N16ZIig/J1lGf/y4ZjPhTd29DPDeL2ygoT6NTcZSwShAt
qdIXZJYqBYXtunrw7+Pcbx7OUF4569B62a/pOQRtc+eLtrKEKKlYGOQlVmZ/wj0Y
gN5rSpuf9RVlu4COc641fh2GqnTF4CcD0wyKUL3WIegDd0xGaERAFrxzEOYq19Bx
6oMRzlrRIu95S1zrTg46yfKzJsTjzaC34opBa9OaqSYuU06LZxLbEXsNbgxqzkv9
AFwSmmDhLYtS7U7D/DeyzpqdnpIHMBd6BotQraE7er8FfALVIVqx4TRW5kG4W/Qz
7m6Lw8LmgkUu2HeVUQA+STHTcmD9DzzqXu6HzPRpqRoV0yIXDlBQCSig33lAK59l
quMb0a+sHOBDjawA7cFT0yBCfm8/emy6T0cOtSLlKhihJd5DVz8WR6x10nuZjLvj
QdGD6Lee7u+HUMk0NvTAMx8O+OX04lZ9/q6wxKGlWnNE9rsDB7aLKZUSGmXrz3H3
kIG1tz6bygdpwHNW6YIQzmEQ6ej1kUfRVyN2a0CrC5EyWRUzKHv5LXWN8y4IrWHB
hBCHRxxcUXUFYk/RYuM1O8xp/R3CpQWy5gCRQENniqMVsiXQIo14Un+mux639W3T
y5kKA0P2TcJamvcOCBvKx1Q5adMZ7bsHhzQrTmK1zk7gT6ChL94p4FDQkeg5er2q
iQnZ9+PnPZyojpR/jZBsX4Um1kRwNpYZEEe275WQu0f8Tce+xyH7VYgAdNEIOuhi
xLMsPqTJSNCLru6zGWX4phtbyXBqgqhN/GVE0snqzuixJEFa7qPkwm1K0kV4nxZk
CDZVHtTvKtgX8eVeZyd9WwFhmiMrBDOGjr6wVFLCTUN/qChkEisVqo6incdF3Urb
bavSJeoOMmS+d4u7Fx3yU7zqhDJwRN//RtaMTFXvzA3rEBRSJA4f8x1JftgvGsst
qWsClIy/8802VIAfmjTEUYEnsuWWQ3/1axVUCCaFpTqSTybnmI2zKIh2v77OII8c
+By4DX1gnAAbqUVk5Eb5yhzaif4AqLv/RslnYsjv1VgTq3Dp93YUkctSEpAB/AQB
ar91/hgwH6wOdD+EfkJVWgpiiVaWzZlxi6i6ZJUFgH//tEohPay8xs8iNANd7OC7
+xukyo2d/Gp2MQi4G5T2t41zkFj3lmNMtncEj4XCSaaPa4AQg4gfd6rBk5dUSTWW
cKFvAko/jTBn3/8lih1RzxWXpdS5YGOWfTYxTrw2w/SkZz2hBhfr5O44agKDhjVu
IK70JIkGRSuVOsgQEXl3dAHJUgAkgh+9Wtqj5T9aihpIxxAsRmoQud8M5ViGW+nZ
rBM/E/p6f2nODKF2fSSxaH4r/I+Wf4aQbEOAL4PcRpvO82I3QcCVqblJlyPs1y6s
NNPb7uFHCnANB4HNolMHOOuAXCG19PDNabi1MTrzQlf0AwbTuRHdmCpUCPBpscVV
ShxIiz4lsZv75PU7qPitq8x76NktnIaLmIQGtDWqXaxzCJF9UCKuQ/Xrh13BceTh
hIIACOBn5UrCgp9g0JQtnv9dqXyzVWlE5z7xSobk0HynKTRMmRzY8qUiV+kqfuMd
2H+KnpTy5UYkbSJdqWyZsqy24LuHrdP1gdj8BTbPvZh4KgLOgOxgSjwy5H2fIkPU
wfZULofY5R13zePx3RogVV59l6gs7RMRLKXVWJzQWr2kcWk2j6Qg89Xx8v72Xtpx
R/ffUAFJSPSX4GcIt38PBw4IR6/o2fygFgjUI4vY9gteRtX09Pnhaen28vpCi/9C
C5M0QUCB45Swi3twzOLwKemL9i1YJeK+gI/VdrEzwEUeTVzVVZibgo0lfaMNvsMd
7GBVer7hPTy058iMDrWCJfoLEh6Qf5IgWV9HWGz0GmwB7bdHU+/OkUYQDG0KhRdP
5Mj0ot/75ROVzQyFyiN/lLZmvtkRurOnns5QbrUqyWSMsb8ADf58+6ccPUcc/gVL
QKVWDpVKvDqjuwthNBs9wBQd+ROc8a+ii/qMilJgonxkq7f5r/SQpj25iFLWHIpm
3yzQ+aRsBy3AbzAfMve2wMRb0tOxWXkoijeBflUpspUqAipqhVY51M8iXjboWT6Z
GJXrwQUxaZ+1De6dsE82eUo/r/dUkwRDn7m9gOKb1jho2HyN/psSwTQpyh5W+SdM
nqiFBg74rivGFIaLgMwG4MLp/lzBVZB/aXygfqFWSRnZvy1pwlCo/VD5aaNLNoXB
+NI/x5n2YLYSa6ZMsuVg6fT/9xX0YxklYzdHWljhgS000QceAmWFkF1iwuQ1tIHm
hRUCjPu0gV9Vw/3gLp8CFYxE7/QCjIIdr1IH1C7SbtZsupfl7Scv8AYZv2u3YR37
P4KLk7Ry5yLvTc3cBKYA4/fss+/qHELJLDakN31SrFfhVOnbnkd1Db6AIZBsQGx/
nRk+z4+RLcnidEcp5UROwX4kwGOYCKpDQmrEyhC/C73bTyJenq0bsZv5gaGSYves
Uqi7MqP8Cb4JGumIyywgxbvlaTR3pPnb2UX2w1tLZamYkR4aZy9LeZ8eUwSwWYMK
v5gnQo4Jio60l02ICCl13CXF2s6aT9rQrBSP8CdAUkPBbjFB/y6+0N+iDcv0EB3G
TflW/k+3yRUEgceeboSm8zKW5eJX9LYah9Ye15XX5N98qXGtbNQLqHbyFpy6n+Wx
KQL1n7qb8IVQyBeOqje1SRSJAn+LpIiQFsAVFmQ0dS0KHLvmX67QiUQb22Is/4Ey
4cXnidBeCNdhEBTXzRtpxKfYHLSJe3BV3L0ONfu/ZZbj3l9H0CmRXD8dPBdBbg8c
ICxctc1tktYXG/hU+H0K8oCEmOKRCuyBluq9o5AHv8dugLd3x/FMx2uRPTuawLUn
Y/WeYWR3f7t3EpDco+PY338vIVfFMVrvQ7iHkjFIVhFyGb92AN99qg8aNvtaXqZF
pALL4HcpuOSXhdQ/6SnkwVOQ9q+4i5+zMuR4OpLTLiyUXA+lpd9EgS0+VYQm242w
AJMGytkavzMN8p9OI/2BlR9cxfp4YHB2UHbraewxrX7pDJJ9lAR56JGDbdh6cfFF
rcYpA2eVzzNYHIAZByQIDFGG2kpm+XvwXMz0QASqg6AlUN9sC+CbGs7bSJ140DRI
ua9hYcDI5NBX46MPRKcSIrOBSJ32RaHySnyyckm3ZMKdlbqyRXvkP+x4mepQLMV3
J//13E7MpW57X/0tgUk519S7FXo3mZSx5zYaZGlcrK38gczCWuds8SlPdBJ8K2HC
msAJu5gdYNvl2aVhVhTKmL+8Se62/Wy+/eot5cf6ZcKEedEQswgQ+rktvNwgd+m4
S0pYJCo2AzVP4+8RbGzrICzx987WCSN5g26ROXKJ3+AVtvzU3J50Lq5bO9nqjQ2g
er92KRtLuaEWS+aHoDn7Lz3z0ZdIyKpxUHRHrl/quNK60oPE97tmGR+hGt0xaLVV
zCpWk8UDXd0Jt8mEpOi+o8aeg3I74ZzqD1kygUL9wOY00//6uBSk/xDudWVVZVde
8gK+1ipbVt/LfUTJlHcFSaqsxGMC0uywXVmxXlnVUF9TXeWqi9nByMw95VPFmpVE
upU3VU3iN822grQ24lY7jZwgu8u4OQFrlWcsbYfuGYkUq+5yN6tBCkwW02LsfgrG
bsJM92NClrShAIbW24DtR2mtIjPHYLSAzNoZhU+UlgDtymwwMOhQkseCmPuMAvVy
gUiVfRH9qMvS0FhufU12FnG494/yNHLHvs+kPWZa4nhkgOl/M5FQa6C1j9ua7hLk
JpQX1o/2ImplTWbYmFbjPH2LLor4g5yqnIwDUtkaHFZsS+Z1xBU8LYDc4TKkUMhn
DQc1umvfdB6KMwqzKAiyopy9Szv2d/deyh008ydnaHmkZJOsQqMVFLMQjFsBiv5+
KuECBJ1xRHvx8Y9hJoKL4vzMaQ5xMQ1e9TVgk95B2n18PezcHP+l5YauKj3J2xXj
YFN0SYbJ6QC8wsd6nCzcfSTHEPglAFP0JkyAAfY7iyRHrKS+ifiMWPVqHCEfRa3h
seh5JR7QESQp9WZ+cEp9LDg4bD2XwrLiGZ/OYE47+cZ68oErllFT5I7+a2dW53Ne
fIVVOe39dpVHqKp7w/BTZPDouQssaCky3LoP/TzfOrV0sIEmtEG3bLi/emm9kkJ/
mj+B6C9q7jLiECgTOxLV4cyMS+Oo7BITt96SJyeotHOfU51NkyeGPleNo7XJZWXa
seq94CI8Rx7bCQctKqM/rxNVTyCB8NkU5KuIMCOlayTcmNWtJ/lYkREspeMXOGKi
rKnpenDzhPOBoVwgdtLytQTF5C/rfc2YRnut7gD88L3or7ktUbyOEBdvuHXRZAsm
JF0ZKMYibzNL9SfopUT1Dqb4O1vglRZ927oKuIG7JwdvPQigiCHix3H6QU5F2BAN
kgScPSmIxxKgcYhNWmi5GO/ayGLZwo0iEtNH0jefwuaUz1MdXmMmth0KODqZSYeR
Y7nZWZXOFhMkv88YYsKVWc38Qi+rcgV1/xLqqNeIewtQ+MQ3eC7Mns+jeWLtH2zr
IyEqZjBn5ItAuupEjSliA1HFiM5FEsoVpK+9Wv54kEZpGl5jBG2jMlvefLtAAIBT
7f9kNnkK2bug41BqwdQgnN1LyN7fTFMgWa3ymxIBd4uhkZpmHqE0avoKaafTKjAx
g2iqZMGQXKOdxx2IzSuoI8Qo0yFh8HEW2od/p70pA8BzLaj11mAIrIEL68CmW4tE
4huarEFCb3Li2g15QfYYuPTYlBuDfL0e7s7pTQC6vRWBATK/XbX44AKaH6TQrnla
PW/xGGpL4CD94Yn3+o8Mnp48qULaITClNRbqGLb+xg0p0x6q18q9bPhv3pHDHYrA
m14GDyIIyiHhxir3gpH54VP07DqIJZu5a71GKUQbwC3y2HhDC5Fb5Ftzlpb8ulkp
fWnqdsVWeALVJ/4C4e7ofaAreyay+MgO/sF8+krvZ4Xqc9dkeZJA8BY2gyq4Lr4s
XJrBosOf5V6HDD/HlHP3EdI2dAS/EznVO4shHryll46SC6gPBJDH8TI0vPqiS3qI
3FyopF9O+iwA06nUr8OuULHTpnq3x6XsCR4onfmPKwaEBYn4YuInfxXBwyFBDgaf
ENIGs3+7fXlMdur9xYGIEKOOXkorjPSecT6UqL+vpLlx7QfldYXrT2Mt+cqxeoHB
CbGG4CE9jdxeQv4ZyN1NRFTlvVmFzHmeh4vucZcCToWPvA/GVq0ClFMUdDlujIq7
3PXWcpHDq2FzLERJLX57+6EF5xk5SbisTNfF+X9lvsf+go/seCPsLH3yO08fJqoT
DIkiJUleadDdAv8LAcQNGHUWjrB1sgdtY+6rKjTzhnAxOQ0EZ84ynY5MkQID0AAG
5/zPiKtvF2QwZEGUGQEGbgIXY+P6fIo6yANLlWnzsY3zO1pKjztf4alVKSuH0XJL
T45aM3lnRrVwQ9RvynXJCdFYDEQ/1leqj+hMkX4DwwmWMRRH38Rm4JxgoEjIQkm+
iM341r2A52g5iUmE06lzYuXfg9Ue0En9wlkiiAvG91BufBAS/EzaPY+HNY8Ol5Ql
ouWFRpsgih7UlEP/pSkkCW8t4Jo468DPQdvuGAjJpAKNPeTDq2t40Fy/VXdBxpcU
3HqelK4zu3yzvTODAZdfPx/M2bafCz2RRS8q5CiE/Cx/7BZzQuj4YRRZW08TU3fH
z7kKEUigbhXxSlx0ilQGZ3zZiqsfgwWKUBHaRbjt/B+D9A020BGNHqgvxd1yroeU
osiOnu0izmhkv5V2+Wqy4/rk+w5t0ZkOZgKKNXtQCRQcVcSRwB9jINiYo03QIUzH
poSJ0x06fhDZlZ3u3xntVdlIzwyi0Zp8mGkxAnrxtl5iPqvOVb/RR2fQaPdCDP3/
lcPHJDrklPPTtHFUAAbnWIYwV07H/EGYSDFt7VNWqE2MQFm9ASQL8GUVng/frKt5
jAryoRw6No2h/xXdC4q7Gv+PzGAAju//M1sii2Yci8tt1iOOt6x9cRw0EMBFQq2u
IxeW5f6Crqde/PS9ycuIe3pGbKLuym48sG85KUWRXybAuxCVh1Gm1fWHokLqqlAH
0kBA/YtA8i85S2TpNKx/ZW128Dp+3jJrba7tY0EbA/yjzVH1fso6oVTYVWXANNlX
4TySeC7YST6d6occmx96BNUY6KjxMpAaOTf15nu48dMYEpz/VYcWV100Tr9Bau1Q
mu1FbaWA3JkVAeCIOpiSlt0bYneMFJRzH1L+tfw4oiL3GUN0Sp14CwU2ujEJ1mpQ
ZBv2+b9HHxqaySnETu5685jkONzeJR1oadSbdvP5bTZ4a0MeOAUARaDGqms1dg7O
IncaQmqb+nXG1ykJvmZqnZSoUaDQXbZr61kDZrU+zW6fH4OjaLtLgmewgifsoKAo
c46nnO5q1uXs4VzcpLgDfCGn9/k7mEpq+eCR5SjxfjTEf/Lg7P7hOoS4ivTLmB9U
XjAapRIaC95V/gOa5F/I12AoDg3w3o75TZRxYAAAaiopmPgRGHleu+ySM01i27ro
zW3OjNtpoNnjjA7a9tm++JciikBO7knDpDMe0YsgWtTXXXoSOhHOKFWoA1gWQeWo
YzahhHDgSbEXaRf8vFjZ2SBqbqfmyokp5zGxClIgkLnA9rWjYuUhOZ2X1a3YIeqc
W2XdkRY/6y6Q/zVKSa6uukURwr/FSC4Vni9yC2tPb3Mvfwdi6IsHs49oLLG7C70Z
zAowlWeYsdR208SyxQnbYC8UWQYWveW9YtH+heZbNAbQW49Xb9HBpHlsfNIHEi7i
eXAGLeq6tWpMpniWp23s5S3YBEAShh1AePTQW7Q8ALeqzEYINcFRjawYdChKZp+3
Jy2d1yaV0r3lqgKcDTm9R/VbmaCirLhIQqopB4LHYvgSMMaKlsjov/PoHQnFX68f
O/81B2T3y1yQRL1IlY8vuznYFMOKyrv5NPT6Y0omzkvZWjAJHzUqw9E19CyICR99
aC6rU6QQEvKIF29vRq/CFiyF48tuzbiHNmZXciD7Uk1XPof8rNgRrUy4JUC8DbZ5
bZUTr2CUDTtNmHx9NaCAj4jB3POIf6UoFV1+ST0gHvoaSZZJYw3ot7gn26auEzBt
2Ux027L3pXJFSNtEp/Zg8iv+dCfKLfCJQBK7wv7qmec+E+Tk8460rvJd1wB84CXT
1BeS6Ok04PQUzTP+uX9nBWTcmiXOIRyxlhudTGAV2IPmxYj1zDAwPQtqWclzgd4H
VT401g8tgeZmT2AF+1fEbMAXmfF4bu+5pDlXqJEa4rqLE0SwtW5lkvvNtPyCtKuW
hK7z0Tj4RwLkwEtYIkcMiWX+k3YdK5MwQx7TmrUAqRUG432K4zzO3CVCT68+kJy6
VwB9LtE4xv7mh5gaD+Qe5y5CZ8OL10z6il9qbVC3JPr9zIp/SNAavEE/uGDE5+6U
jKV/dzb+BxTChsd0t0gdpSRoPffmPXiCMus8RseLCCiWw45wehfswbvQ03lDqr54
gY7DKekLGjFc8ONFkmchT+3nMxr4B6AGA4tXba7BjmplS+aUT4ONwhXXfa2MMGkk
sOqrivhvRc0ibJxBEUjXFAaG+lIv7HwEo1RujR477Ih5Dwey+tyu6h/CG0Om7xRV
ldBrnkyI21sqXRlU15AvhwQdLnDXS4J4sn/zL/p+UW1oCsyI9whetaJ6tCsNu/jl
P3LPliMWUeaj1T8fIRyT8O4XaCf3oXdxUAml3xQx4e4xjwqF70PXIH5Uhb3piXGa
ZmI5EojZnc9r0CcuPl2z+3he8QdTs2U6LIl/D/40ASoKVOOZhO2nH0Etx5hFQmAI
hSqB8SacbBIPM8o2d8JdBPmEQUlTv0h7qfIWfr4v3dphSv/YsdCBggD58KSN6XzZ
QPnL9vGkLh6YFttL1eyGfWQ8nxQHaiu6f2sc0mgGk8ehbfK/Y86hslPihdo7EDkc
XvcEJAv28T1e5wZH4OO07DhtX7p0ic/U4nvyrVa8K1GEdAzn0KV+m05VxpwEUDkG
LKm/yErbH/7Oc6vO3XJ5h+5pI+UOzq92u3IgOoGX2UXxMrgpu+KoKQWxjALNXkKS
grBGCqYMvuWKGBrZiC5gDHje+v8jhGADZSqi8NLcZQNcAUMAEYdXMXDSCNMMWiS7
qbucKL6z9mcB1QIk/rJjzH2ZjTNhBQvwkobCmlF6fps3SUAt5GO4VxY+ukB5NnAI
IxaydUFZhgOq2bLnxbV6GLzQ5jTxiS8xlptXntlZF1CGLqmQp/iPGkghTQfI06EN
3NASwjjswfLPAGTUW6hEzj3Fo5di66q2UGpVharYx6YDGYj1gdH+OEQRUZgEjEIs
QAS4D5emvUxm6Ztm1mfQyDCtpL0XaS5siBPiVUtCklQkArk7XQZeHnIk7hwIY/i4
9qP8UtdDikPJfFZ6JCk2i9GFTyZ0IVkAXkGUIXEODSXmn32tCaJ+3/DJOD+hRrMz
Fu/UBGmD0almN6orMfgQAPcMR2GIxz5ZJmMdoHjifelGl5St6tdSl1bCcaHe+qZD
sxoxBewg8B2v1nNeQ64bJrkOaGt7zkUKtXB4zwa9Ti9cUWWGESU1jL8Ddsq/4Zi9
z/0QM1DCYUGh4U0+a7D3vODl9QpqOIaq/yXsek1pUQzOKpzHKEp4o2xNxLl2GIu0
G9boIpTqFfQDyWnPxCXN8Gzx8+NP+n8SgDpHlljSVBl9JlmLsGs9x5ICW/EnocB6
1bqALN68AJDFerBDTe/FHn+zlgHDXDAQfFx8N2dEylD+EkSHH83iqIvamR3Xi4wK
Kh4xT4kwBytpwOAcX8b8+tz6DlfTIera3LdLc4CHigXzawRRmqta9C6UkpFrlYuF
y51N5IvyenrVpufRSU/gy5PSl6pa4Lpi5rZ7J03OGBr+g4arJQwdZ3UysAZVQEN7
pfzabhX94+0HsOYvlNmCBph3W/0X7fR+AYOvSl6NVeFhnXsk+25FIRvilBxTWfos
JaDL/OZ4vo/549b451ZW/Ks65Uk+/YJrsr4Buu8GmbslfGgG5IbMT3HO/rzMRh6Y
g0UCx6EuiK5LlegQ/pc/CHO/Ki0nCwYSK/YVwMuKOjHxsGE/mDgaQ/7lIJLmkATw
KQFbpKcTPYgaG8cOzgMhkwUhLSjISFmqGqjKur+KJxeDsLJDTo2WS7PBN65N10Ou
LWN3FHWP+Mr/K7kQCwnVGYKIh3huakTbTo/Btco7tp1nMNi8BzY/DhhDhx7RtdUi
PNrLnIIak+exg7irodGrZXwwGBV0IGmSGbWM5gpgObDxSgh1XhuD915LdI/oURzW
5SxWzpC9e+4uX/czcElZaL3qetMA/WSj2tfHzC545/XmuGMKSmdXV0F6kLVXkfgZ
EgXs77IQMilZr7ANrSiL+2qi59hgmhlUPzO0h5HgToF1b/qJ6qhjvJ1+A7rmbOtB
y6mE+ETvOYKRdC11AxG0ZkCiaBT1WPZcIwnim3TJFKMKgkEZueUKRbN7p4AlRgDK
5kTmoWB+7ItswS214cSjplh4DC8v24S0DbwuTABO+gFmSRukYaodVrzDlA+x1Ch4
TPasa8FkRNGnefQA2yBq5/FtYrFwFoictKJoJdOZGGknbBOB7y9+qEQpq+whZaiU
DqL3oKc+LOktLN/BTMHZ2r6Gn95vuaBAqRMQpUhC+ieAKi1yr5UQXGWw2hj605xS
vSSX0/L8/q/BGctNbhtqcUn5RQiuMDHDpF3PMsESAiRgLFnetgdjM4AojPo4dxdO
5f0OiXdX4YhanBBXSDzWdJ8bKG3pvK5GXHIX84edrfG888hSwlxt0tsn+CLslVX8
RCfaM7Xy3qHvJw0vZazIgkvQLw9aCVKa3Nl9SxCuXnWVLtDOUKQqPXyxdsRKIc7w
pxJB/ZG2U3jb1y61mQfEjLdHFG1/I1N1ikoL+voBLIhi6/p5rz5paM5V+tbR7rWD
zFxseZjH+Wo9UxlnAs8Jrrcy8ikIDbDw6zKxrkwgh5FRDsy0ZxO88p3WqSXwApj6
6A4wnqQfjQUDvoGPeoY3DuIyixGVFAEenE2erfCv/rx2hSBbz8OZ8wF6N+xuAC2s
+ClMbNT2wUwfX0ATgY7QGaLurxU6nRzpo0qG0r2bn+l0KqKRC76vW4frmU+eWl8Q
OJ8bXuIeha8iJ1vDI7xdhum2MdVK51uEyleIcUrr19wMkMpMG4lPjm9iQe41+Ds6
lTFFYhyEqhKPkz/qDkex5jQ0n9tYMjvWg2xYJeSnBDnh9YAi0BgrPDry7HmV59vQ
J0cQWsOwzHKTL05OOVynRNBBZMZdGHHGGkBtRVucCt4Nu/ibnltPeN4cXxzKs3iS
5b0R75uVpQ7MEaI6yKuBEBn61qgLDM2Ou6ca+KZhMN7dtj2fkFb8XlBhjWV6bfSA
m5HU4LUDLOOjKO73BVf7DrFbrHuGfSxoIXt9miwUaNWlxSRXmdtFRjOVnE+7Q/X8
Tinszt3MFBJ8sGbVoOZq++GqpIjrWgy9e1NTaZ2xW3qCOGoCxdGbK35j0My1hWPY
VvaNaqizgfYZOcta+SqcBHkHjv2VEeYbIH/3GyjNzQfzOKyBXOFNWSt/Q9e7ixqT
23orFvYdcGJbSOayVijkSUoz9Tc87MJbgogJ5gFzMEYmA3i9szVlHqPKYvW7GkGx
ZTs2NB/dmxVZuDPDQ1fpf6ocZPax+uL0DNKsmSmArBSuV5j/dkYVhr23+UfmAWuj
7aLdeHRe1oVCkMaouXFVsEalc5wpj1xZt+IxzlKn8R9sBlH5E4z+j5kW7QwBeIgq
edr+rRPp2qTy/MMlFw0SFg70DY1Zp02Rg0XIFtg+L3kUo2gJrWzhdauIuNIDuim+
XKcOaAXAxCD9sO74JrE/NQPl2o1q/LhoM8tBopYMZRhA+IYcXorM0fUhV7whgSxs
Ebbklx+E+LgOWV/namnJ1bFjJJVb6qdBJc8tm52FzxYlzdUasFJbQsBDWE9JA5FS
NEWwvU6TJ/0xdK/2hwMZfJLg4aEx67IbPyz3VYdlgv4ptuQp3a+98mfJ2oIS5m7p
bLsdyvfv5oxY58bJ2BAsCCxKUkWrXYyV9QuhQinBk6IYsMtMaPWZKGoT1yuzIVA6
Pax0l89R77Skvr2Lp23IVuGf4dfeO+cDQwsWK1cF4kv0FhuAMsU9ZlOe5SPIWqQL
V6HzW+8F67VEuY8rTCtzq6RhFHZsBWClHC19QAo6KmTURIj/eCWYu6xGQiHgAWpA
93nDIsPHfy9AtJEEPUqnNieYoVaE4tvq8lOTSWVE5k+Jm6gVy1ypKWDcJz/CJa2v
hui9LFy07vgCaD7FBlBWh0sDu6XZaxLMjsWFr+V2Fi8cjW7XG1bRnP413vPsxIcf
d0G0Y4ViEW81QrGLfSh17k45BOwyW+jkLe5QpC0Y/6PXuEQL7p1AxfORrsbHBBHu
Ta/NShOKqJAJ4GOMUAeY92y6sd6wbIshJMQKAml/FfedZ4lxFWAymnYbxq+Z2YNb
ffWlw/9sg3VC34YUdklehYWbgIciCy9bwugw8R2cHLn3uM0Y26nCe2wTzWd3Mq5E
W7JIrevhx0FMJHCpTFFi0qPu/PaDvM5DszVoNtK2MD8O+8J9Pz+3GeWf6DljrlfP
+rCqdBMxg+GqvChhkvG0qG3m4O0Z2ABrzb8mhx99vth9hZZbFtk9+E8Gsxnwebtu
yfnRDJoB0e3wFzb2NRcN+xxNsMrTxGp3t7XHm0M78/JJMC1ToZXuNE9bvugvLF1u
HaEnyIxs9em8++CXNka14Et8B7c4zUf8PmAt3AgHPhig/e/vs3FmSX0BkY9Ooiv8
QqSocImpbI0SPv5y0FbZHc7T9cz6C4Cm6leix/hLdgYtb5KxbIfsHa8KJKgO3GGV
lrsdCtd/5o+u+Z0VZ/TVisykoTOh+VRBuvgNASv5txL6uDJoKVJR4Ds016sl6C4S
wN687Y/Js6c0JoH0Zku2BeZb1gttMeaxaE2v4nHMBbLFSvVDtsbhxKo/q7VbCRc5
jB5WCnEDXtbApYE3OhDz16PP00budWOoa01E7LDAj2wa/oZ5ZE7hyC6cxtqBJ9+w
57fikETzo/8pzYWDTXAm7XU87xxWeqfE6LI2UVfj0Kdz41W2Ye4aJcADLa1CdclU
1RLaBA8hK/+LvmCIhYoPKoHFaXxyVB1ZLxSqW7iRV4ZeCFZgmBBM9w2aDB7lUkuz
AboPnRJ2phjbpqhaOyLs157KQtG/iNUlEag6Mhjhl90TWnsF2Bd2vF+tv/tc9+Ve
aSQoV8mzDqMT6n9V2pzcUDnEOyAlFUBw2K7fHwLQFAltoWDzlDPnzQECpE9yX0od
wQOfdNTw2Zzj83ubW/O3od4sW/wKNPmpGJn0EZJC/WEbCL3jBS7eAXjrZvsgqD+5
cKg3H+XbeokUD3+vw9CL7gwxKRt5KtTcsj08gkZw0I617mZZVa1+KVQd2Pz2tqzD
l4cUj7K9KwmQoDZA57Qudi+3S7F3a1KR/Xr2pHk9UQv8GuFsYv+zlV7GHi4LMupN
xLKi0Bd8a7yiND1lS7H/FQG4WfziCFeJgHhfPFr9868NCCJxTcn3S+YuD5LOWhl3
UXbxMoqUiKe5aGX6kPQ4W+IJFWLOK/jMwWKnMggOYZT0juBOveDYuxfPu8yFdyNJ
SOYomi3JDQw7hxam3KZP3PtH5xklUR3L/04xutjBrwkcjSxzMRT1urb3jIE+HEfG
s4cZ96RzldLoIQlXCpm8734+BDcT2eoyTzCrBI59gobFiyaHKvx9Qk7p+m0Ixinn
4Ow8v/WH0yM1xcjyESYGVDezrSLQ7Lgrfgpjq1f2uonGfomoL/j8Q9SBfhslhe/4
bgxsv5vft7quT3VAG8ylbGk/cE4aa76UHtBZzVRBiHjToAaQm8QbWHcrrmc1s/aY
YxwXT7OUkkyuFdk0kWSL9SNAUZVGIoNtk9LVj1/OieoYjyiq/s3QVWq/QNZ6iZOX
OyemT4YvZlID22vmHXZ7J571qpVXpOklY/9ceF1dF0p3Bjw4HtzzB8f0rtGNHOwF
mQeTB09gtpvgqta4A7JEtBAZhylkC/L93BNerBEKqCOaTdZBi8a9ptK+U4gYAIk5
q7TfIgAl0RepNS/HpOwssbmbgRh91ztOHM+Frss6LX3a88ZnLMZxsMpX4lUGq4Zv
pWOiUJ8JNlJbgKza/s1OGOmSuOyWpzfGSC0VddjVOr7s17wfgc/yl0/pEiuI26UT
3o4w9XL6h4Jasejhz+y6keThWFeno1auLpk+4oahvWjAqZuxc/PX1/KbQk/R+WYi
O0qNI1HOzOWoS/NZbs3aShBTwjV80YZdynrnqF2A7N5SOjrpdLbU1USLAPA4r7Os
F7QrnWpp7wtr2yo0LR0qixUWktMguBH1dnf2Hd0MupJiTyHITia/iMTfUrj7qlI1
XmgPRHssnfeZqBlI898zZl+XYMu8xqMz47yXI2BcIv2i5G8ona/DZ5pTiP5SxayT
zq4a1i+e/ILaKDHF568Yui4En0dtZj7v717szfW9bCCcEDOPPSbeJd1YbIFy36v6
KX4QFE1doNC0nAe1WAkND4j+SrS/RiAKcRA/1j9xU3qIpgSrshlJD45cpDilHFKZ
QKEW21pOOsjI6fdH4lrHGoTXceyQRz7SR5ztfzENzkjnfkxvD4tANNQU3Z/rcOPZ
WbMOtLJaikAxh1cnp5+iX88YCXaHTB4AjqsFV1B9+vJAY6sgRHz7e6DYzNoZQzHu
hOOSEJ+1MHn5m0YguryqzbQVh2UrOzic9KNPYrHwxPG1EXDDNk7p3RfvQhFku503
xoliQX0VEssi02lSB39q29/x/3sRWtMKXiiF9CMhilR1J45+k1d2gHIb9dgwinIG
4K7VHHr3aHh4TpnmEqPmANdSREObvHjAGX5BL2poKzLmlNypGHNin4Yd9Wn32Nse
FoCOCJWIfxURJpPyigBMw3XfRtjBvbXaRM5O6aOGhUVLZmYXcpMGN44oI+LJyu0o
+gP8BK4/R7mAekYL4D6MjRlf0UKLuOVWLbzeqwNktMalHm363jeas+GszsYxHGKQ
gfATYeEBab3u0bmyxa2F1PmYPS2WpUO/XSk5ZH0/10NKVpjw/egdrpwZwUfQ2DyG
j9aZF5Od4iUsvPq1sO6DdAv/53FrlXl8MEYcHI+mcHAI8XMOk45hBO+gOLW7EA9a
bn8HD3wsVaSIi0kgcKdQKo1vUcrXaxQt/5j1AyQMyUxk/ZAIWVtjBYUqJn+siUjD
BWrS4/h02SIKOMhGNKLdvVi63/uuxD1Vkmp0wX2X/jr/GF9DA6iyQSh6ZtB5XSWe
uCtTE/DWo5LUITerG9D+e8GzDEnOD8TOYfEoVQXu+xgOkObRhPl1J6ugNTo2xkCp
6IlvOqUuDFhyG2hmtwhvON7vBe65noWID5Ymk6y58EWJCDBFbUz96zZJPUYjVyGA
yd6bzzLEfrL1mfp0AycOr8z2g7SJi4YRHX0rrIQY8YdqBi+st5u2/waXvWeojLSb
zxzOOM6ZrMlaHFaDSLSZp553epCU+/ypMeZB6tM0pnv5XNM2sTFSesctqBjtb/Kl
HeJzEMOQ8T46LEBW13d7vdzsSj4EzlcUC1UZ0KutiX8S8V6lt0XJGSS2BAgxRw54
xadR9sZq9jRLA3XDYRU0R5s3CVWV5Y9W6ZoazGiJYg3SYZFi/0couHJr91CNPTIn
Za90502Ly9IaDJh9Kx+CWqE6BGyIl8rJyxXGIyiESUK2/Tq1SrNoa34wIJBBsPeS
QGuWPiFT3SmabO1+BDfGjzzeLkhBLCfNZOtvXZBIlH58LJ24/VvgIkdtNJOFGp12
NIF7CF8w7bTUubW2TDzwDqE0ofyW4EBJkTx2YeGXGhDmTvHqHUQUGvcYufTNEFvd
gHk6UlnBSj5tOLje44aTwgt62hB3C39Izzmn3KJdKOcfrzH1taqSKL0rw1sm9Vub
8MeE7TstAT6g1B/xcnOZbOi4EvLvOsZNYxjUky3+3FBaRjavnPt74D/JhMD1rfa0
iY3r9KDj3XLAYLxp1J2vThcRYoG83NnLwMbOyL9pAHJILhAzBrpBqzJK91zjK1rN
/aGgQ4dHfDGsQmufCUgFCObgBzBZGa7BJAv/mUHd7jwXw5K6J/1KrOGqL2wMOOE6
4eq2FrbKhDKJ9gQJSdg7XrFH47wypHahy6Go07FOON1TN8cb4x1eejBNyQjRs5kn
15CF9sjX0pO1iNbRpRXAEN+emxRcerHM3x4qKvLOk/SZ9U0zDxjhKiG5VJ9sVPRg
ghi24qtiVi9kc5hrK7tefjkA2vMVMO4VujNIlrVYYAyYdtXS+TbfKCWvNIsJshBK
nJO8gssyq2KdA0gXhMgKNtBnOIjzahueA2763JlhrJeTQzeiWdv4yMgD7yQDzeAC
diU3dvv9eBvZ8olXu+pr3CQtjfZ0dxRMnoNxTNgsZIzhpI+oBeUiSrrUF5B4imXj
YtWAvhFLOlXcxI13lZvPX5Vw/Par2sM1qDtMWb+f9g9M4AsFJtpJwP25uigKKQ8U
yEY6qwx4uhHx0zt+A0KrMdzDfnHGJV33MU5GeYknSwQ9aQ3nA4mGtZZ0aloQxSMH
QvKmYTLd15yQ+axxB7+UZouxGVgSenTae6XqEZArCny5ohNU2jjqvnX9gherFzuf
rdb2Ebl9AWL4ZWpS9X/O7Q2aIbsNrc9+9x6ICDjal7q11eeSRYFoBp56+1OZyGfl
6kDnM+fk7DrEyLaXoP7b+4Ct0fLxW+2oz3XLSmB9jB8Mcda84q5hI6s5T8XWNe0e
HqmNypsJOxdZ1iE37FtK3ehQyF7+EVDQxaEv+zO320CqEPHtVMW3CbuVsRHOmEmh
q7CliaS1mqMKH8p3Ye33/KX80N4l7/kbKZm4x0RxqgD56+A/qpEMvxlZMfQoIzlZ
mhJmXNyVCbO7suMyqNgsQwttpcy7kWzTc8pjmIz5sSVAtnSYe6RKFWNGwoLSTpwh
kXuTbTeo+hc/0pvHaU0brJn7f3LviIKYW/WGR8qd07ymyYeH7cHn+uUsNJcTGL0t
ek6AeFpCiZB8sKEdiBVXBkG2+W3ohSCyABrwONjEG+PZBdMmlhJIXFV1gKDzmcx6
8Oh+5+nStfR2GMslG9kFjDDVcAPbVFdHMlN5pfBuaiLky9se2PMkMHTWszVAhAFw
46xoJXGIY8T9b0Zj7a7ClkFlZtPnB2PDwpSPW6mYj5XW0QEU0gscPYE2vY4Z8sR1
On3/XlDat8A2ivS602e6Kkb5zLNKV3ylZiwSvgVAUpxzXlr2G87b+LfhMPdAc8st
NJi76wNi4Ln79fv1TVYD0Gkmd84fHYjLmvkEUP+4hQCtgTtGWZJvAhg4DeBOwLxl
ol0Yq/1X4O++zhflQCHRvivbDJI8+HQ+oaoEWwpJ/uo/YzLxrz+vxTmQyU2ix2Ok
Bq71CRDd4O3ONpO4JmLkZC28VDNvGHD2rbpF8eAP92TmCFy8ZB8p1LDiFu3gDDex
2FG4L5u/gdkZqiXs8EGmac3re5Zr/VX58+J+01ZNOLysBkUZTI2P0rlaUE/+gGUk
xxa8sYP3V+xrCpOr7t41cUacw7j10p43d9Q1uXUeUB6xg+Vkn3mN7xEz0uWwCoNp
wbUaxo4pF9xGUsmbUqGCBlNYRWXKVmh/tAA5kt4i43QvGcirXe01gbQucUjNlzoH
1sg6LBGN/B7uYkwgJ4MWJ5izI1JlOdFYJD+urUGPmMkTIf7vuhX6hVcia+ysPUL3
FpQN7oI37xEKyrgiaROKSNVpkYuCCBkNOdNuK6MHfgaFQsw3qiyx9n++wPiNy6uM
SzmRy4T7GhAq0OgJTayof7eKAOnl9iHJ+CX8NUbiitcuKMsN27cdkb/hiupJnYs/
dnGguIPpfnKnOP6RMb+fbXPLqf6sOEYN1dq1TXkllImhBPsTyB2dli4/eJ0ozRLm
Ua1LUsunuQhIygBUxMxGg1Dr79pkaA0SZu71YFLjnEnIw8ZfGibdZI/TpgTR2xaV
Bf5QrjFmuimuOoBZtwTM7GyqRwbhzXZ12MBKcax9zlKf7mylFCtNfZh+6l/hWlo9
cK+pG26PGhV83KDX2Gg7k1G2UAc/BBhWQJudiDfZmFwWhx1Nf7ifrmi4VwxH6Q1m
vBabrWwt1D2Oetu41jXC560LWusgu93LGlQ7tM8k2z3QS8VzQIvUannbhK84edlK
fLix4Erf9NmLXQiUcrykHPH+SnDScVMZuSW/zvNmYUvK5QOyv2O384mfBpBU0u+i
hp8EfyRsTftnabMfG79eP8Z6yP42VPHkAelNnAoeS6CL+bY7umlU9Bfu4v4yjxku
j9cknH33BqNqCsXRJQoeAUMgU2zCHoyLj6vjavb6J9hO8Nl1cBVVnNjmf+LPKfjJ
RbOgZV5NQ66/lAxV8DqMkXoTAgNv9bBjzY1OTxKlxiKtVsAfRtt+YNBjEncjJ2/e
v74KAq+ZBU6E01mf5zKNopn3lC1NSFn4muQtB++vKe1SIiqZ84FzQ7gssdp09kYn
gWYyrOUV7+W04ErO46ZOhxu3+VbLK/Og0Ah3sbflxdYffqa5F4EJfdTAHSaovBAH
C6+fmRLW79Ny45XDFvnUwOJjIWbhkh7ANbVITzJYTNg6PAP0rQkmkyVVaH3GyTvs
zmh9pmp8wqMxjkOgdLrLFjoupZJA3ppG+dIJw4dzWYFJa1ZvJnTQqVdi0dGIX64C
s2IbIzR/rZhJilBWyF3yRDKZyGlBlDZaHDYdvZ/bn/ip/EpVQ19x2Io+gGV46EQ/
cgkomUlkvznOW1cMNcSqcjDnzHsdKlkzyPIbK7+lR06jIMoUGkO1dIRuP3kL0sg1
XAVdFm/agbkt2VcMJOBw9RZLKY7FQ8RnNcERYbgkhj/sBZOUg/VOiPfpA+SkmrlT
jMSXen7njH7Kwcu4vLPdeKF26OERLHSd2UwZ+GsaYPw/iO71HfKOSg1woDgajQeu
N5KNy0XqCcfkVqBVt+sXZtInvNAzif6w1InlWSbLgrmaBmTc442G7Gkq7ALTOXFj
2lwRtGLKk8QRnkaB0WjuUbQko9Itlpq0fox97UOPbDtKZsBPeZWLeW9IGYhh3MJU
OV2o3UmrowcOv0TI8rHzPGiLfOYxGIF33EMJ5EiKE7BVCSuKiJvLRg+I5nHRv9Sk
tezXs08D3BrJWtlQl6YBxbdSTbE9FoeXLnJQSSd7ZLAXkCbnu6faNdWwhZntBUOJ
0rCefuNY7+SmzkPE7gt0NTQ7pf3ompxe6rCG27xokK9v8DLsThbvzztvfaVgRuns
PYvONGPsYiCub7Q1ibL0by7hl+lfwfwqIgoyEC9eYzZyRDeQiCPQrGjOMronsobu
ozECb+ERnTuAqiMJQu53I375LWob6RZn1c73XUSlfaZV6pGNKwrQarMuTf50MpvU
5EXdRGM2uZWjRPiIWieDWwBAQUOqqQt3YuNWL2XaDHpMlF43I8jPHvwkFkzmG+P3
3tk/bOS4bacfn/w9vtRKz1wc3c8brP4NCjfHqhWLap4ev6xoaAxkHV5XZ+KriFnU
Fll9DNA69kuPWXrVXcZQeakMsr5y+JKPZaKaPHCwxEjiZpt0yvxkddb5aofzMn2n
bAWWQvodMvigw89Mn78NROvBrAoYTPAgp8zleYOIsK9rELvNpaO4XgNKNeBlaMlN
faibJTVHt3Dg4bHfLqYEqfAHFlXgbhNqTflET0z4KxeHX2e9QBZ7on23rkeJzR8c
3geEoE3VXCNgwDdVF8XlyoAyljeFEUTOCQ9iHU2Tp8/Dglf5hiovSNVQWd7aeIc1
BSH5hAQhDMnkd37YbX7tJHYHeTfxCn5/BjJpwmLfEJ05p1Pp3NywLJ9nz4LSLxbK
IjusZJPyEXGInQmyrv+3qk2p0wMM9QYrbATxGNRcsrEGkdNIKw84km2KwwgDBTb/
Hr2KBzNOIRfw/79eatx57OY9Up6fIwrr3/eq78sVjhux1GpYjA5dIBoCXPiprEbS
4C7pPahxuRyKL9982T/vO5/P0alPWdHsC8uqlPsIOC2gSVsJ50VHEonv/ykLrrf0
HlSjinBVNtDAbZBz3/B6BNGt6gTUqXDA9Y5c4Rx5sAEsr4qRqRUEV7kQxLMkv+/d
+oavhn7adtPDTouglHNo6oQiKHhVOIJig87kYkZJEePqf2Ca0oP1MNj4BoVpaaaF
1/1VGYJkdohb5b5vHb5ZS+gEfdzy4hpv2DTw3+mEUJzMpgaNyH34bLzJ9GjleQEq
yUmSC2ferEPFkY3VDBgYL0lqX1eFMiU0fzx+HzzAmlBbwLcfv0K0GRotcY9+ftnP
gDm0HCZlbRYCYMxjSEqMftlKcdKgcJcYTEAKC7FWSPxwJR3wUkRrFz4apVi+A5F3
gYT85aMHAdJbemvqhWVt0TWvc7FIioQpC49mY6FizjnlDIeTfpxGylXA43JqutQo
c8XNgD4xgy/pmJVHgDHZyxAL2O4H2jgDan9XescrIumyOzbQ8d/7ogJe5aCNRdJr
zC32Lw1oP7cFQei7s/37/y39YRUJ5muBFbrQGa4TEbkVjuGLYGxRSweHA2q3IUuo
oe/PRDUZjjim8EmydNb2ASPfvmpey7AxqVHWjJqZ4dT6SxfNDpU9JIvG587dxFl/
3bG3S5jIrqkI3mUVlaMe2BmVAPnFcGRpqKyUBN9QFEZ8797jmPMINIwTv9EIkujh
5OTx5X5tvKesErJbPtWQjPhELmRaASXNZlx1v65ovW6eRAKGQLJOxdkp6jFRh595
3Qf5bRNPzY2rVvYoN+r6Fg0KN2ETLaYMrWqSgon5PCZI5wH1g8HPutc3heLm8TgF
cH7RYH/WZaZIGgBqlOG2WTOhvI0vXdZ6biHQO5rVxlWTgnlNHSxlt7VpcjRYAMC4
EYY4MhzbdfyeCs/FRkq4uawkO27EC44OwEqlGZL3ESpvQD8jJiDnleJpKHz3MBQc
J5QNoNNgSStastiV6Pk2ay3DVxIinLtqboLnw/bvtxq8lwx3ojA2jz6ZPJp+jcV8
Q2lmqxseBgEi1U3PjshhPvViop8Jr8akREc1vpLgT4giAqGVP7qpkSPGOa23IQ+z
bY2K/23hEOTYUyD2cHc2ixo2Z1izSoqdABnh7M5lmf9XI8pBxpuxktBBKU4lA7t+
CfrS4r4TQUeKj7yAkNFRD3jC7QLETBzoIQaH6mkmQuSMLGAh/ynFAoDRd6BoYDBu
95u9rweTI0SKOOtFD/4qjhb6k9ST9YLzrI3OylLRTGN99jSa1gINV6xw4VoLpQPe
dSaRfzU1HZ6HuSZLatmnnjXSiel44en3qjuRBYhVqJA3xZ77axvsmopuny2dHiA0
f1zWFhKHmHWvoYVc70KufqFwPuRauZhz8fW6m96p2abW90JTijG0r2p+pvHta9Dn
LYk/4l2WI1hojgoNQposcL75zSMazFbhS1hyld5PW3WD7iiyi034yEaNt1r274iN
xgXGUbwsU83aX4tBunDQsyxTM0siFe3yRqDOU/3m9reHETrEZ87472MuyooMKCZT
YV/GTe06Y65Tm516s1Y5jgrBtoMUSvacO0VsoGDercQBnVZ19DXqgezKZHSSspxO
mwASNpkeUzijGR4YSoWfjqV08WMReSdshu2g1QWOaxfK3nURXGXRHxOzCMPNcpBG
QK57xJjE567SiL+cGBwRsq/eOS9FJcEHGqBmEaN6DZTblIME8P8hSwTAlAUoNcq9
HdP+kY+4lgenFi+dGz1Vg0Yv/LjiNj8S5Hr6tMspb3f4dwDd/+C/4CymiCuL+K5V
SRkHEn0Bb72E40gfsq/4oOKf7HuLOTjNy5QtFMOQoGwmUYPp42PDzXMCJUrIYzcF
5ijkoK9P9WDpfibEZhuvPyP36WZJlfT1hci3xz9DhRCvwRziH43vctC7YpkocYSH
Fi/FgK/dp4k4vy70puWpVjhz2FRs2TBLGL/k2YATBfw/TRfKYmgjsmurIy72q0JV
Pn43SyUWOs37QlCcJplXmZqfpqohuHvUEQvhhk8Qqi30SCMjRuO/ayddOyPeBm4t
l1Y9azBHn/XNP6RMDfiTasQNgf+P3Sp55jMRM+O18mXRhkxyD6wA78cmkAVCzKJJ
JJE8sN6x0dqgQgOzluUrEXS2+XCYgFMrOWg6P80a/U0VPpAQ4fyIb/Kmw2t2Fl22
swhES7HeLM5YRM0/Zh/bbREoIS5cCnQkLAkoUNOTIH3zxczdrmIdHPQHRXMBh59v
CGZS2lG5hj1UY/ZgsRgOpCIgIcxTLz5NVKHOhxuM4iTPmkWxCT5Jx67NuOEkmlym
M9HK2GCMIvL+ZI4s/BBx7YP9lihb/6ryFX/kd69mXAXbqZKe5FsEGHTWm7DTSAzG
eA8TiYYQvIRD+QSUZMhNRKSg+nb9EgtkIxfezZGqK5cJ36ePayhwYUTB2KEn5H/P
DBBUEHgTf+goSRzbuHsdaLNXYukhLuwbMbwWU2yMZOodrnPuP9COy058+yjR746h
0iy4QVHVQBCiHDCRUFiedd+cK1OAzo5D3NYgUQupsPHvSL5mzpgE2wxQUfEEQs3j
Mc6pXSxjy+wiihkGFEcGmJfI3o4hlkTiDh/oT1cO6alowtQDsDOCUDHj2Uaopxj8
uI2xJFfizbcH/4vWv3fRrfmhZTVdpvv7DTS2FbS641Y72MtHm3dPeII+HkXVhWC4
GW+EOhOSxXG9icGlI7Vv4WakXEGgL2iq9W6KjSchJB4tEW7GXN5oS4P2aKJmXnpe
FIEv2XTHMxquhayXiwjqdEu+9mTGX3GeyNsx7FktDizPK0bwgG7gPIH3j4PHltzH
pF2FhwhtXzs6RF2YF0cPbGnFm1NIX5njWa+mo1swVFXdJ3QhtPezBsS/znNqJMYy
aC8wgAc8As4dggEsdXdgWdCS654NcjB87wdfiRTRkWUMK46VagFyA644aE7/eYVH
Ftf5PAED8CZzpE/kxQjvXUt+d+7/Dy/04gRAPsonK/HqZzxfprgOt2rUEG4xNa6o
ziSfNZDFHAryn3E27VweEixHh1PAFx/KQ2381I9AsxZtyaobGdSR9JZhulWz08OC
Yiyu8P+p7fYUgVe0MBz9BUJgVmAgZZ2D0y0Ylu7xBIkJeYD/kcizCGAXrmFbwnQv
jm+F3fmoXFkqN6OAjjbUMWJgrsgsd6eiw9c6O1WYpOE5Dxiuj2zdRqNYl5y5pb1a
mR5bdk19eQB7xFESN0s5h5p0YiHTdADqmC+rDUceNxHlNTG+/bTR92MvtdnspIWz
UF5qg7w3ZbHuSzYxNMcSRHvbuMtFr5YqdHM1CVKrK7g64W+EZMfnwmch5Mr27GOY
satXmOJNRdRXwDW8xcYIKf3/mge0k5iCISj03mpDAZTM13vaMG8xpue7O9QB5j5Q
cgykkiRCxen0H8WI/JP9e5dDcbHX9qf/tUlgbZNMF9lhFuAfv7UkOK9W+pzgnMzt
QXsSAV/BqsSWsd+i3TcnrmpU8NUqnz4wWAVtIpVFx67rV9ygBsqGbuX2CV14cOVy
vGUNtthpmJh1qrPAZvG0hnOHSAH06PrGUvDQY3Oa69ldcXuXXNX0MRlxMOE6VVon
a4Nin7XEUIuzjGa5AVly2YtZMTpCcCfHJGkcIcfN8511eTXfa9+H3+ItFNee2kDR
LbsTmboigUQnIImvC1C2IrMr75AYuQ+WjyqMchkITfVgICW9NMaGAiwybZMg3mWQ
ruqiwGGDhn2hOpVndihyBqkgfe8Brjo/my3jM55uQx8pGBFL9u7z7eSsWyi9JGM0
nKZAASMn4zPLa6lpRGtxZEhuVtQ4A+/qSPKM6WWg3AS8wpY6EhsFUl40HSIL9VXv
BVrmx9zfFq1VLYZFraCtHPLxV1Gu/LjFRrztBvJp9obNZvCsO3n2VSpUH3jlkxe6
B95WOr2kdk5V+wsEoC2Nn3kpx3OIiiH94k/d6Fl4d/MfVg7v/GTEzlbcyVvDr848
SMWbspP/iXgN21XPcVIpVKOc/jhT+AMHeEhDTESIjZvQLg/jV9C1fxmh4auVb3mc
2JoXX0jsNMRhxMrKj+clbosfdeMt/VQ+WEMWZgdt+HWFhyaCVETuh0yOpFNPytjC
gT2mve8TNMr0ikv2wNw8t6tnhTIujPseYksdvMxiSjjGcHp+KHF46RM7HcI1KEhq
vO4Mr5fe3tV3jvKQdpRHT4HUKS8l2oFtmKfW4aQfBOgWJDiI3RJEA4CnDT0s/v2K
BZkaEGWapHUAnSfaPu+JB10gXKzD+nKxCRldXfvj3cVTnGiNLFJP5zOJ8KBTS5QO
usSjuhgLII1mNEG17xhgUQpSV1EmP1zp5Cvkhb0nqqM30hGzhOjJYlnfATVe9IV5
0VZlh5WfZfey9SKWt3TntZBN+u6IaQaqvp2Ci9eKPrIDO4GkzYqan5uWoWXM/3H1
f6zdgh6f2mVZ/I2xN75rMg3pqB9h9c/k6caMBiL6sYKsY+UZfo/HtVGbtZDfjHMo
7J+bRASn1wIhgSVFxCzhdBe3J3ur5nlDKDMShWTs/6m9KVvHquUPPnGwLeuiy1CS
e/OHrRagdNeuv4JlAPzq8W1Qwc8pkKXVUTjUL0ehKb5AmEWMLDRbUNKCF2tcxIP+
zhev15VBhL8BnajUe/osKD98dq1r/dYjVGj/3NqLlwy1ER/04tmvY+6ZRImvkVWQ
2OXMoQAdwVzlzSLCi7uVYvZHbFTGTO7DEx3Tgsq7AuRSkIu50yRFiHGrjIijuhD1
ad0505CJsjEMImaqldMyKz/HWQfalusMN3tT8gP6JZi9eeXkcnHiuUNmOjRxc6u2
W3Um+uykReTNwchY1sOkf0kqoJN8lCTyk0HDaogvOl3wZWRMgpaJeqjSM1TMgozn
oflMMvoO77o+kK/FotubNHr2mvS+/yelpGYvam44btWFJL51rZdPCtO/hVhS6eIV
FC9+9uMHzOkbmRAiNu5jEmJhvVlH8QqyM+stOzpy0ruJ6/XoEqHksemnZwwNFw+3
NHnP/lAKdhKLqEgVzl/mLIQLPZPh10hGXwVGcRq0qoFG+XHWu+qpnTPBlNnAvZzN
+xylp9fImtFWjLABdkfKPfgzx/LXYmNgq0QyBkCXQqm7rGYl9lKDwXaW5PVuZXIr
duFxWX8iboMBRVhyRCzaE1cvfbOp0Q8eYlWWYf10FWBG5/GVNgE4R+kHOjyF8bt/
SWLt8Oj3uvOvHP8WfYcFLeyMuFPUuZSFiU+EcYD7tbCdAPhwcdhPrui/CppoDNRn
aStn+Y+Zn0dWC9Q4eNNnsNpBdy8Aj7dN56nDuBLi8tGT3iJ5VgEvFWa8b6QOhxrd
qYjnFnh3wU5VRjzaXkAET062srHmYmejyze412LWnHer/vTJnGCEgXBEGsWbvVrC
qlpeXm/5c6joKh3nLLTg6CgJ+hlint+8gJ3Q/Hjakrf4zCm7kXRaaW1zAZQFBbdr
+rHSZ1Ieh+ahOoGROxkT0KPmRH76BJgYFucjFeLcfsiBOWEI8/JuUfT58xObvz0J
R9cezSFM4wNR1fsgz+1guL4lNynaZjFb3E2S0BF3O2OKhYDIsj1Vxnng75X0JW1P
gXeDeBS9dZwocOo0QcSyHKEmqWkmetenc7ICGHavFElsSYXUukAAdgkyXjLi50ww
oT8U5jITZuo9dGOiGg7R+szSYSKsupgtmhx3Klb+fngOLEc4jd0QWO4Us5kBPUR3
KjL+uKR350aX7YW+V4pEFmUJh2rIJFe/aR0pCsodPak6GrCEhAzVJnH4UAJjUIyK
zB2mRT/9bl6qxGhkxH98rDjWZaKFpLwqV8tnMJpfmWVoKuq7m5Fww3bnkNhacsCC
DqWXQSzaCPjvN3Vzm9enw4NXkvTRnsWIQO1s/YcKo5WqjAI/fAWcer2s04kJBNOZ
WxMn624LryKCJll/rIQO2lsje+V5FHEnue99j9mgrSjUeHlh53g2pkP6fyIpQTPD
mr1rDKTlwEGxcVYGFEWQQiMNuCwArwXJhZpiWVDk2BhgBV2yW8V9pEAHph9K0m+m
axhPGWkNOPUKuuAbuxPmla61TiOVK/g+9IcTZEu1AQ4zm38BjauUf5MPYp6rt/g2
zZ39dFOlFyifU0uwyzMh99/PgSXx9NOsmmElClpevh9cpDZWB8kRSTZcnTLZtlB6
5UT07zHJc0hkbclfbkazWU7OApFgre9uH+n12KV6nVybkZqQlPe8mQ0/G3oxkNQX
gqp/i9moTA/H55htxKIYYXjkeGifaIMzgE8qz3oFtWHXMDSa3ix7Wx7oS6OSm4Nb
ObkuTBMik75jTznvKRNIM+1f0hkNO3v5t4Gn2fABP09cbsmxAueW1Y1WT0nMHRUM
COayS1eY+sSg9oyKJRDyXfe8mQ7SLyYcoS5C/VIFdkgXOscA+Q09Boo1aoYU+mKW
9oOX0RAsGdKAiLnJ5vl1EuWmsEEVeWl8npLdO/7t3cCibmyc0HnbxqMDEdxC6xxF
+n9DNgD3lxx3LCurPZUKgr0AgAkd1q4vehMifYaVHmF3yhm2v0xa3SuvdlIQDCGH
CYF96wZii4s/lpupUYuT6m39YtgA5hyJimcIY43k+nEaobxiGe+KwhdoatNoRx5e
torpaj2nEICRsY3l+ueN3Rps2tdKTorTjP/q2/3qMm77lhXcMfQrnIkpRk4AkIs/
5ZX9tpwEkTVHcKgn0DIZ1zRz3QjJJafTndUcEHPyNk0mwLXfyIA5neHEeJkvbrn4
qeEdnZiN+7H5z1JZ5kMFP92BRXg3PZsS9SEpNVzKW4ctKwp0J4NprdHdmONwSQqc
P0+isGfAAkaiKBIOdvM1meV+gQvIyIKt9q7d+Pd1GFxo74YKpx06kGfSHhAq+mn4
mv/1pX11mwHAf9NHLoi5uUQlESgP8JdEh4DWiJvPzLvc9eAtl18iDqE44ndiqpfn
2iIh1vCx5Fpmdu/ERULtYWk37nh85HkUULd0SdEnTHgqYr4xu+Gec/qzzk4ogsju
kQMIeUYUi7SEhOeHT/JM1QQSORkT8QKN0oV3OFhOHW+kcgkUr6l1C/iMDhj6Nd/c
vsUEmxVpCuTR0UkGEWOAXuO5oSDMaU87o5y2AbOToWfm916ezPE70jbZspMfC0L5
2quSg3ucE2+7esPLXwPL2aXWI9m5agYWEAqqTnh8OHJ+gLlpQzbzOPRR5Mn8s5eQ
5HmeEUvX/IfxdJTws8H04Sa1lmLfHIVTYLEG+IxM+yY1GrabMwWvdnndWFZGD2WN
CXJw5jW/qoiTBMhBXGPfxPSJce67jVvyMs2noqXOzBmVngYJydoiPV4D8qKm0TNO
Mvd4u2SnSLLpwYsr9l3wepxJsYsoiq+Fs07kw53GXFQeLt663lvKh6+xSBH4xXJM
pyhkpZ2tCywPs4OeZCoAefnBIlN62XsmE58nNdtiwm7mOR8k191l+V8a3L2ezqmt
ZCWp0kQ9qUXJ0WjBmrGuMWQbKtl2ttSKbr3iG4ASP5XY4EeNxHDK3hWSiaro3EWQ
WhugZDFwNId9EXtlX2smf4RMuW5DPXet202tcd9nC9O1+jncdvYXH/hcDGt/bQ7u
nIxzULgaCQbTYwaLWfStHyHGb+SDdqprH1fXe9NEi8dDnd9p0FJ+qpfQZt7yBr9w
bmcmaB7djePLgokG90YAzgeoA9Yp47Pbt6IWzA9mViFPMsvQ/8xkzigS0S6EwH33
QOggTlU3qsEJ7recvE+/sv8BsdjSPMItQfTWqrQPnymT9m1SB2rqNTpR6jtV/V8C
SKk1B619Gb+waC7/C9zPk1uyaw77Sg3bFtfj+OPYO9fLMYdPCsrd+bHVE0SAgUs3
83TNNmvAoQNw6OWFa32DPBR9Sf6ccv7IgFl9jOVSkBQDYMF9K/d2pL/+INte4zii
ZBfLcITmzb3huUu65BQEciUnOd9feMZdQsXu1Q3Rfsb4iOINMQFIC/YIAYSbgsaq
mPhmYQ3Bn/wXQOXcJAiq0S8+LEC1AaU5crFxgacRLFc512THbRQlR3Wp6DhQw6nW
c958xY2tSHgpFWF6aD3WofvxEmTuVFsbgQE6RuDU+vKYZryPIzgKh4tqmoFTCnWn
YpzhCBVc6iL+MVhfR6b7GfnreTOrDEQ5g9Khl6YaaJ+OCKZkYvUV4oCPPI0yLyqY
hUWWlJL0+fdgbxD0mPOwKQXVp2/clOnvRfTifSYqBa4sG7MSZ/jMjgZxIWdzpZ+Z
G1S63kni1FyOcCGHbseKDKp3GyF1mWKTgolQIVJrZdMDEus4fXoUpuH2SDLazrTg
xci9i5+mhWluCJpdLCymvVfZeaJv0HX5wT+tNVggaPyLy7fyfsFfrPk9oITc9dt9
siK3TNS3WEmEE4idkxGgEi4pb3BZWpwjEVxkZbe/HIKLPPidFPM64OeLTEi8G3il
nRL0XrqIJzYk/GAK6oBpLN0Bj5Bbl5YBiQRigKsjMtrtX4sQVAn7Ft499Go0KLbp
nOoHgMpT3kEfQtTMyjSYxApKhrJN26ZUF//zr2jenm0UxwxDQB3hPfXF5Il8H+5B
UNQN4J4r2cKZc71g7ZwWo3V8WAsVmx+xBuoI55UHivX9hHKqIq1re4by0tO42TIa
wYmxCbOK+TafZXrulurFeZjx0Z1lhm1j2l92BycsZCWFFICTKUeMtR/XHuVkGt0H
ReFlaqzBjDV5UmF6+9u5D2wuHO7+NSkkRMFLzhbkfZ1xUGnLWLVvBLXGG0kUjNUY
pikn7GFsWt8Bd0i2F5Poz3uSn1MGKz6lZjqbxvdZhsKDo0O0QG550X7D5ZX8hdbH
LHz1B2wzrBzk32OVGwU50pQG/tXig6C9ASJHmNQsCJNxifDF4lWNx4TLE4z5dKV7
SdkBBFarF89fZDuf5jXfVyBdPgUyZXN9SEN0G3/o+YEzvbaxMWX6GXeDjb/O1Y47
Cdaa+a4wPaYDF8UN85xD34nnqKYCEI9eerFYXC4zTdF62n3KZWNSWpxgIvci8tcw
2/AMI91Oe1Z6fsc10bTbcLTK1nmMnToMIzaeGEQQU7n3SjVX0n5RxDZ5QDbq/aIt
jHMjcO1FUsPbB2757/bwUofMzGEvkky1ymeGycWWn+47uAt30BZgzdrwaIERxgsY
8ibMVt6AbRAl0yOU9uNoc3lzoVY5U9yPnV/GtW0gncD1PZTcDZfVSbHC4WfY9sJl
eOQu0TY6rsh88+ZKW9Kzpg1JGboFCatZzVRDTX4HRf5GCNuDFRylSy1aMHMawZMu
WJ9P9x63q0tp/tZ4sYYxxKfBPKCpwfTCfluCAW4ewehpW4+s3Tao9FmSov2mdyyv
vxuSogbTREZuRApVygM2mj9SNml+edbrFuERVv0EKgRV76NhnaXEfi2O9GrUCHoD
rJ04B8nV2VCaLL6Cw5cvLZJwPeJkHOO+ZEn2SPJ8p2/dYPoFv2jCk8ytOOxQhVyg
wG+M50wLMF1DpUwSVUwCp9RHjqN/gAjnXrqoBx4VNMwxlo4jKctgTTfhU3NXX4Tl
pnMFq104UbEVvkIumW9abMulSI496YQEuCoeDifdpThUTmAT8mCH5mZezvUV20jn
POrT6zAX1YuOmNNzpto1aJGzGcxK3/DI8JnQSuqSbVzS1BV7VuX65zT3Rgf4K2u6
qmY9xLCHIFK6VKPe2/V91A+eb5OaUZceQ3ogrwZr8oiEA9Mi8/+t0w19O9FDB9NY
L0J88fiKO6c/kBgksIdoUK0cV7/2GgV7YSMpzCT6w/o2A6+fqm6Lwbylqd2JBRvB
9WIbFb65jkl48avPi2LfBwv2EndWGFPKBZm1nOeYfy5VCe6sp+16Ha1VADmXDiwc
NZNR0hqY7X7CpzcpI4E6ohiuRQ6654lYsMw9occFa76shsqlGvHONuloeY3WhqQK
B7zQhlaZcyMejSfjRYOmQajtOcbgUMOjM5TgOBsNGUZbWcP6B7L4xZLs6LPituV7
7x36Sx7Sj+EGkS+TV9x7/Z5/L/VomNMpw0OH5cTbUveA96aoeWJq6QfFnr+y5xgU
MdyCOHsU949H2/gIpsyyj8cb0NtMFOijQMjoN1QO3q1WVsxAoQb8VTkISCp8CKnF
QleOmw73MgeYiAmr9/G1sQShGIusO3iVteiav1bKH0Q9P57l4rODyZJI6ihs7hcB
SLqu+K9QtzTFLidcjPpg2HdYc8/rWJreGg6m+OOqdjyQxM3sasqM3nCn207JIc4P
2/xkviNbUuB/C3tToZdCneZS14S7JfdzZxEc1uUKt64sAJWoAAqn8g7BVSS0MMp5
nm0d0YjLNXatr7GDwdeerR8FaJSsLJ+dURScEWepOjPjIL/FdZdJFVfTJFFGpdnm
Nc53XkB6ass/ANnCLL954GPNfZdDe2D8TzbBAUPa7COlh5xApYQ7iS2bIEWKp/fQ
co57HM7I3yhfB8C+/6ELhLD9iXgTHBQ5tx2qYzYZ1bnGMspk5DLE0aSovBsAlleh
yeXRjoAllLEDGblEqTzRfiChI4ZXqMMSm7krO09AyjRUiYeQmFndyxFSQNz80Bw6
8PVSTK1yGIxXgQb/CjIXvcyJgyfhFwIa5i5oyRnO+ykHtwLJTIdKeUSEIDZy9xkr
cr4/ex8rxHtEa3wUroGepxf4CXBQD7x1vn3j3iNdAQmkUjm7qfvAJfPaOonzTvOT
+18/hgVDF9Sr4TtGQTodadfzKD0zAS2AuKb/gUVDOCPBXjvAOhc93D+D9rYAl+uP
RSRj5UbF7k2EH1vmTzAaGMQ0Fa5TgBcEggqrXuhV/mD/QVHG0VKUVc+fk4AMW4+X
ryGQQuIpINDUcilcPDj3DZUydeKezAqibZhHhPD7rxcLStaDSjEW3O+NjPn4uejf
KSxpfez5+kdPDag1js05KFuzs5rBJVD5gJOIpHB7JL6cub2cuVIcGsOoeEK4p7mB
R9/r8v6yQUnJcgz7n+Tn21/EICVm3sHgLVuWnfpK0DbSw7PLQm/jWChYiDtUH3p2
hlqo1sTjXMgAQ00/+SjatjO5aHkqEJYZFQ1HdvvbqD+3X1CcpVsiiIJKnINC7y27
sA3/TKdl0Frj9Mf4mg11MAH2JUWtdHcjflFyv3pKVTBA4yMPj+u2FZBnyQpKrNH3
obuK8cxYXxtdT05urksLfXTnM0m0OH/ID9hI2epjh0Ft0U5WFtohu7w5wnB6KdW2
bvRt4nw8JyVmAWBt8/2MMg/XAZ7cpYbBa6BM67Sfu38L+k+2UwBCdAqve2+g050l
FJfDbWvxYCKcweNiUijjXsCXLbaekVwQ/jbAmsM0kF/Ck4ddpLa8/kTt7L8H5Cqe
nfOEGJ3peqr3/wIs5CxGvVIqKDO5gGqKU6CTVsRO4N3Dp4TJFpm0Qq22m5MkUeMn
42y15d7NDLCrECgmMyin2S54PH7cuIxnRYPeQMAXEalzqWCZO5+E9vWEgtBtYf4E
QCBrz9UAlv1pGEweEb3z1bI6FJGmZcmL38DFshYPtrJUvhZ4ZqnewtoO0Yp4CVHw
VE5JOTfLkAkQSV5dVCXlTvrWpO3T8BM/Y80fn/pojzqPrEcq+rv+TJmB4tgaskKT
AcC/jZoD4eFin4Agec6XYQx8Vha4teBE+urOsQmackhXEuQuH6amejLjKIMor2VN
L71qoUYHkZEUCuGiOk/mCzcnomP88+Mho4AYkYPfCgr1pwXWuZYC/N88PU9Elg8U
m4R+FK2wArK7lq4gqW8aeScb8bJR8f+UyAJUXshvAa2Ti6jUJXEA7i92qd3A4+70
a+SlO3IKYcH62ivNBLaEG1J7zv30Pj8gPiiPSnueXCp4diB+CQxIQhMRM6jVndqE
a7bx0rkYXjow++k3bjfXjMiNWQKKlblkeM22UiLu9E/L7pu9TzZ0PszS3RCOpBKA
roaYqzG9eGkyoukR4B8H9jUPpPPqPqCW8rcFESYTEVRFqmUkqSeZDx20vq2eaCgu
hfHj60YjNBOhemSOXOwFjdc4EYgGQ9WvGN1Ub8aJlacQcPoN3slaPGxtd/sfvLD+
jkFAthNcJvonl6urAvw5BHNpl0KNeStMq3NdxHX6QVDKyDNXsXVMLSs9pCvjPONw
d1+P4umqDXsi8HlNJxLDiGLSvf1u55FsPEEfDBtwTmG8ZGGwP0sIsjIIIfyyZagH
xUe6eVR5/ktOmRgrnXEkiMb3M3dH3qTiP5MA0Ffy21iSqwvxXf+dX48xV4sULGku
8OL25sFR3i+9I1SCHCYA+p8DjI5HSTPmc/oTJCe6vHxDFyg2kwWvyyIH/qihMs9C
a+cAgWLPabfu3WP9mqmVNElOmFfvPrA95f+1MYpazkP+nE6sE6dcoh8AWBsw8pzT
bgqinf5iZ0h9jhZIt8EwkwJoA+TlvvZXOuLUuga095w4P3cQLDRw84bT+vwUMIko
Sw0Ztj9MON6WrSiatiOs0ZSwQdlhqcPo/BhFZYBAt+QgBDTrOnxQz8wej3gbPr/7
FiovDCFS5xN4no04jrjte5BVKrc68dtbFFxKbu8QQ+UVyJfwjbfAx9VxjOMCpYOi
uZ/M8iEcbfa/dOxTuMKv8ShgjuzK2V2O7MNo2qMpBXKJ0QHj6b51BQmSlRIOkN3+
vwtaKHZ+Ccbmg4JSESUilVXVbKquYmO/lEqILANm6dubpadfou2lpfYM/dza2oZG
ELYLN6Hq7aImAsrUYKtk4+xkCZIU+OoNlRG0DBnm89ZpLHiIf7ZZhU5nnPlugz8e
BlwsdT9MW0H4OxTFa8nLfMkm01WYROndawhrusGE8KA25THJvkQ91bDS0LzVHKG5
b1BbMTcAovZ7MPpYXFZk+c5emCkhUn2qEjszTMZut+DAKGdIZbL9kejWxApgW/aC
1O39l34JdExHMnnySBhGebTSrQ8lBNc7Cl9o8VHFL1hunBxehr2mhPGdFmFrsSKm
gja71eUso7iirISgs7Cra2MpEDB+KhB1VRDoxbGHTSOkyW0JScgSzQ05NtBYXmR2
X5544lNnpzJagzaPutg276E9CK3nI3dHKR1zg9ZTfd48MMVfnNF94rNAx4J6BYaO
3X5GkClxbl8bCtwgc7m9dC/ENPNPan62OBST3lT0hG5boysIscqwo+wIJx46YKdO
lbzvw2ASI6I/YOQ+ymoDFBxxojgZX6DsDHZcF6tOGtUW7thRVtyTzT0vEouOvZb3
zhpD1IhogRMsnZuq4oJQtx7f33wWHZq6fmc9TxDp2J/N8sbJZqOXVrTuRFtFgI50
ZBDrCQ4Ojl2sjoA2pz1859/9cCxo7NfFg6fKQ+zRv+4qAPJoalRPmAadFih5TQMP
VErd2MZNpFMPoX4JNx/zv4zYMTMrHfErTa8M6tvBQTaE1xIJCnlXEX9+ZP9k9sDG
Z0dQVVO5f+rrbAWjqxkqr6szCv8CDOtvIThr6JZXi+3y8Do6YW7xwrKduGDBXVsx
YBZbROgadA5J3/1GVyOddsRh8Z+5hP/GOF8M6bXgcHOqbjyKwRjjuyiPExT2YVhi
1E8lyUJ4oIQbENPo1KG4OGsKCHGYfXNBWrMP+1WzrUVtdzsjGSKGmE7K4kTKzey/
l8O1CRA2yULMzO1iIWR1R5MW56uCi8Nsg+OtyWgUMT23N2GmoxndJ59qS8wb/Bdz
LNTB837VV6G6pT5jV5PSm6Tr7jKAFpC6EpoLq45frQtm7V3E6ntImW3fPzp3g/WP
Nk8zR2fzYgWONHs6ghTdYr0QAZRPjUem3lHmykw9T+4+WYbTcC5IYMXr7njw/OAh
guRx/TeWwE1pvOuPxmgCfvkRlGVFIsbTXWW9OxTl0Lg5ed7ENXyTLVcxE/qehBOM
wUymT8hN8CiU03QqBVm4YisE6d5v9aFx6sgiucJ9W1EO5AXcp0sVHD7UV14JtGep
gx5aD/m8RglnFwxkQZ144nbT6SVk85UpuEEl/LF8WZOOHuZIHWq1mnX5lnTtuVwt
KhLhwRlz4aqORc9dtGaAYWgDl3aaPpSMye7wPiNM6KwaDd+Mg6fV0q9Yk/WiG00o
UY4ET5cqU3MN/ciKNjvN6QwV38m3kPLTJh85+3KbxVZDmkiYIk6G48BxNQ4bCLMM
dSR9A91ppsvqlLvlu5D4GcgDzo1oKlT9MvSajIttNno12FKltLttv6O9gYNG0di3
7zoX8/xwB6B6XXnzdeB3kb7vI7lxmvHQgxF+GDGWlqdNBaJ/utfRm5etg3XVRYJ8
XfYIIZzXTX3l1EVpXss/pAim5v30MKUWlTLzvhhZD9+fQuLvF3WpekSm9oOcNjwO
udCrdmSVxKJErc94iTG3r7VSLGcW2PLdlQh36fLC9FOzN0gaSttGUI/292PxBre6
yRwjwXMm8YEma1irna4Cuj9t20vvnCh/+4z8eW37DstmSUBBlik04v0IurckH8y5
o1CFv6RYqYxA/3xQsxvJ5KHoHKQGsXF/56jkc9BdHpc9d5pPb3Qg2rMWJsBUDhPw
TCgtwMgeROb5RdNO9qZAV4viiSvAb/0IfiHtmimc/H9usvrLXML4ixW+QQIMz4NL
il+kzndSbaddAOdjekA1nTWJCRBr+pMr61X6ryo3T5KU4ujL3a69OhICcIlo/C6J
0tx+6DzjKLYi2uUHBL5soUO587viiOC948zCZ4umyGueWVXb/8XC/78ReP92N8wu
HUC28UKwzHuoSKVlWy6qjKCiObvi4Nszc1l6RDCouXCgwew9FfZiYKLdjJ5tHsys
vKo18uh8uAc9NbuEJ2hn3/QWLhGwhLfkNhK8qSkZJQ+m7GE3Bgf2iOSyYeYUGqru
1xAOV5jj1F+r8rpBo1mdIMKT99yBec5PCxuAb9vbqvpCESQGh8sZxBBvUaLSCUqI
ztjygtcnUYqjC6K49wwq2D1rX528oSYjhMLj9GN4Gi0/kPhJf78TnzKRlYhAVa1c
AwXm3WMeQeoARuRnNupjzvXuey+iWzAPe7UF01Ag015n8R0J+9lJSHOVR7TcxSFd
HYZoQMeyELUXEOQ1iQYwpsM1Pg0+xuhQUXpgp7edM8U1f/0GJB1EQCjswDYKI/4Y
HtEmXoyXFnbQ63CKDVq/STJh+1DCb+mhMW9jVkaNzxhh+5Nl8yGFKPr7zcLjlXTR
vLRvBRlR7OWdkL72n+JDFcWQLfEsvDSvDNLLs0fGdQOT2QnpzD1sAUHVSVNXxjNA
TBE3U5ZLKojC/ROp2sTue86kBpPc1OhSMJmF4mYXheiOq3Yp+x34rZkYkc/PEtJ4
Trz5jlWqZmIbUZ1/J4pGuC0K+T7R6BO5WtSMvdwgToM6iYzCDaLfSw3BIXXUdRpJ
fRG4pGKohKkFW7/LCbGJ4IG0pTtMAS96RdtOMXXhyzFzxYobobE/Qlu/l7hMisDG
QHmpiF3x2Fp8l6Zfr6ygHDKEtSO8i5VwJH08/kxXUNbeBQPj+qrUTjGiYbGF9Rrz
5kSSDlCFti7vy5fCpVHq3OcX9GcWKkGP1xps0d2hKzn0jXqnjxZ1uHDlEBWu9RT5
ootmnhYYIPXfQhm2REdwkQ2MyrYd72TdQldt8Hd2yUuoVa9l6MHFkzGll95WGTtn
XxkhB+NN+WmUJjm/f9loFIzBphFNCLjvFLm4MY4fDeCaR8CcR069sWr/1MpV6HxV
EC5qQxiirmj5HgdG1vBC6vOZmqblf5Iio7ktcndKckt3w/X9YIPBdTGwgQ2Rdu9/
en5+JSYQoBzqx2T3aVmIBDjFq+8f0WIBtmD5c6P0igjUb+U1YdxzPiijmeD6F4Vm
7/MIS9XHQQCGPFfRKYH9GH5J7aq2Mv0bssK4DWRp0/wqeZDc2xK87PWtV8e7aUwV
zFG52QB/FptKD8ZE0IA71xWANiSNWDu8yOxL+pzCG+4Mmi5RReGj+n/wnA+qmFVE
EuME+lPOehOMdhPbK4EgiDgK6fl7dsXZsoZ/s0X2ft74Boz9apbB4SmxNnxl/aHV
OUE4Elawz9kATVxz56JzIMKDRC1RMx0iM4jr6vLhyE5iqEjlUfR62MGQ+auqQNRP
Nkt2J+VuVA8TI5cRKaCWS+Djd8oH55QbV9+rO90XAONzrfRAi2mPNug/zCudiOZG
IsxR+yE+Yf3MjeqCM4PcRMrzQUU+up7YDO2kJAeFbL41dWGWh4cL9mNFP9nE7UxD
kx4xJbi4GcvtLiGhB5i3Fz21JfhCnfo5mdg+551ozr6agNiLL7DaC09P6fbZiBD1
g+IqqnSUiQ4EiU/hcNimcea2ht/ErQJrKPCFgztJTxbAzOOSyWKIbBBvPp6NrTBj
sk1DOgwxbnw6B8kIiLmhdHdDxNtYjEyNa3zjFgv16UZI/vKC+cAyJSsncXym8T/O
mifurSbCTT61Ip12zCTYQKbBSonPwrEIH11LPF9bVeVTPUJtbshYeRbIQibfRFJc
wIdVjnDHta3nRqt0jbaVp/ABbjNYa/Jpuv3YfNgd73LMrZxvuwTY2CHiNBWD1QHE
3FR0gsrglHRbPl0xdSGN90vSt49FdASc8PqXlaF58N0aV+Jd74sKOb3KCOvY6YKC
F6+K3MU5aPI/az/0syeu4B0CPZ7nqKPnQG1gjHfhFOiyV85qG9vFBZSVsxBhLSVu
KCGWw+xUjkY6nqurIGV8sl1rJjqjbuPh69W0Kcr6DM+eP6SHdsKbyvs7Z6zH70aN
gZ7TVlPU+u1sADlTiKYeRKRPO6BPj2n/ldIohqbYJH6vLCOUVVnqF/8ySbTC3X3q
O97M6J1YZ1uCLzRLVNGEH28RdbYZ8FOLgnLsRwuz2rUq9qimvudlCtZlEWSRxaZC
RE4iREDJxMbNvGXEP1mEucOpXOUcId63lPDE6l3vSoVeD4vdlfeN0wSYhc8EMcY2
qjmoN2O4frrCBtSus3EUFJssHo+jr/IglN5IQlabk48K1X0FatA5wmTb0YU4YLqP
vOjZ2XS8cHzPDMzxhQnkzwH3WYgS4dlEu6KqZndtc+XUwB3MyN9jMvpjWDsOqfRy
aESA1QlfHwNa3cp+k1DLWJ+6snH2Va/GrN7OUIElmqBPXQFeWGCW6cOB9Aof7OEQ
miVqh9yMacxSUnHVyZmo+vUJvnPalzhZtAwNKhmxzfIHCUZDY0R1pyhYnabScvmK
Rmn6V9I14p70V1QOcTEdgYvjkn0l9eCSIR9q3DcLOkVSbRdEbcsmE1ZdkT3HZMAk
kzXpRP2KDH6/33wecxPZoObf04eqOlTObqq3r2Epc1L1U9IxZ7G8SqPTmXSbkB+8
gbjBT+0b9kwx52fY0PCKCYeFelg1hIdZEGmq1H+f7n8YMfMmgZ+J0v1y5FlBYbOO
ny3CoPKGN3PPHbsGjCQBJX3zDMylqHAGrMeuenYnOAvzRO7sl5udkPUZLNVyfDpt
7VsT2KT+LRtMiZ2sY8BhynDHq5UYc2J9BGeucVTRAa1Xb5prF+V6pU/Hne6I4hHu
rUausg0mCf76Zo+i1S8LywDdeOiYXpf59IpTn08fw3MMeKeUjBGiUqycdRjCBH9x
jB3McWUHp78aYJihdhOiIXCIPQPsxUPg2jlfw22uv8QPAzSBAwXVvjNSnsJGVYN5
IVc4cnOfz3N9kNOYNhCU1bPKjpxWM3rqzRK7T3fuFuVPcVvRlRrO6iUqf6R1Nydo
wbFk1kiPCIUE8q/xi40BhAY5g7JkZVeSii5cN0ZUmyH17pYXpv7yjQ4R2/ipHL5U
h6XYp8W6LyUa1W5J1XU/Fl9SLsYHQ1Lxctqe2oNJpMpL+WrPRJtjdKA5HAjr40Fs
uDpj6/o0SwkHZtm4tRTW3w5Eqb6yAl81lSAlvKT4STLOYOeYxLoFQ3Hnoko0Ufw/
AMFGdGlZccUxJJ7+mbfIwuWxG0wCELhoYvbRP0HZd0pE7eKXBlEui4GF9HftG0Nc
6eqRPz5u+wXzwt56aTnUd+5y072BUYKzC6OjOMk6f1LNB7p4KOeFJeTmE8Gs8WEy
O5YuShiMWug2KR1C5jQa+MafKcF/4nb6zwedET7E64VPSJ2qMhuX9yIZ3EEEATH4
8Ar3MJqTQzc+n7dhn6WmrbGlbISMCBeiV/yhThHH3phqw8QMOf0x2gMu4Zy3yWzm
MeLv2wmefjsyO3tXnnRdZlIoGlW07qsx04k47swCvlEAFKBetxHg613pvx1YdQHw
U3ELdej1k+X6h9nbAGS8/D9a97/QJfrkelUD/ooUozx0B871U5vLCD+kwQzM5dU9
EM3BsxTbDwBIkKLMft6rd2JCK5/g7QGnxfrq1xXNLIuZ4uX7y7NXF8Njy9R7q/8/
h7Aikd8vJaNPcL7HLtEFahO1pJ4Q3AHzCiANCaE6vwcCJkKm/5YW3CcEl8IJ2VR4
1/ZdZggruVciVyIAW7+KPk0vimsgV70KCDgP/TASjPrGf4v6FsK2PkLEIf8O5GXK
p55sSgvtzLAF/zTRgXScI+gTtkFov4F4DSNuiCerPQMuun+Y7b6rvght5tCgOq63
2Tw7wp98dhDgfZHOqiqRVmRLQEFDbU3D09h0oI/iADP4W6fo/HqmTNJxwGUzCjTy
XXiNW5sXBLChqLlsHkaIBIDCTlsbKBHg4CMyz3R74RBPESSNVJPfnY3rfQFoDe+R
8+4L6d8XYqzIEbrzf6HkuPEAATQD1S+GaH9D+yvOE2RGztpag5X6cIOf4ALgmn7C
DkydX1AcjnP414vA9kUrGr0fU9aCgUS+gXiYdtcqKvp/thuTGDsY11gK1UCKVooN
QlJD+dNQVPjccaXbociKJZVucN1lZERRRNn9bR2Qmu3nJU15l4woDv97EEQo1QmR
AA8OyaZZtmSz6i0ewLImJRfzJxkkBWA1XX3UzrkMh7+kIK2WVNpoTlAZ6nNN4x90
4/XFfAHNnDQbMWzDpZfdDNtOtL3WCmr9bT1SYn09Mdk4IreR1I6tIHIguBfMnSbV
cYh1Wr8YaG2pNbwzmUGixmnmums7xFUXCxgp3PubwJjduqM+E8Bn0EVPmlAEIYOA
YJP4N3vjA+uDeaE/DcZUwVhfT8YjbbchZlRW5+VvRnZwI6n/eewDlmFjj9tz0qqw
Nf/n3R6uvgISqdN6iVmlbrvxoXaQVv4kGUDdFAWQ35y5mUTL0c5fGiFDefsTK/Uc
KdEVQU6IScQ5+LF9h5wQrA52V8qa9HOKGZ5KvbRanQwNDLUH7Pei1IT1bOsLBJYB
D81hcyP7AWlFC0gkbdSqgofgK4t6NpIoyLdxGjqEwBrCIGhYvsc5m4jWB+DtKqR0
9FM8i7JV2XTr/Uy3ZLez5UjM55/bY32PVqyjaxjbI0yX6V0bAVi68i+Ccd4brZCf
DJeJn6s7Z0PzQ/8DZaux/QU9VWMOVvG7YmPbUsAAspXLvJXZo767NpdHbFdy3KVq
FQ0YJ4IvkFwdNeCgbNCqtCmWw5MTgHG9XnDPQ8XPH/Q7otUhpCGH2/F2VFreQcBe
Zn88KkofxDyJpgyk8e+sv95G1dtTZPZrCzCki4cLVaUCLVK3NIsOiqaCIQzIAMAI
uodFwWCC2e2x/2S16KZLImxFv34+9rB8OSjSD7JX6LdFxc+nP64DEqYMMOkCNUnV
DwhpixJ5xLmMwkC6QZG6d8ipua+Vz4bbnwtw3AJeqD3EyZJFaxbTBOKPFJU1kyf8
SIXm0vM+qrOvSpVKTwEEaNORoppxpfIf2J+1T/2a8QtR/UEPzOsR/uJP9TKIF2H3
lECVm5WVOhWufGMSXTaHcGlJWxYOoJ4UZGYDveVzr2eutISIVa1KXCzxwTUxk3F4
3dn+hvX7WcVXXJ0j74ALrK8hWJ9CV1poIB8aqCQVVLDyp4+qBCFE3kpwpu84Gi7n
gtjOrTNDHTbrVKDkFbNG/Fwsizd4xrUvGIYAKFQSK0977AYL7NPLR5l8uCAXQTKS
fTvo+dbGquhGfVmhhMhUgi9qQkjCBOCeMy+YbZ0dA/oP6Jy5ItJjZxsVlyYZhZ/n
498QAXdi4fJNQ1gABDkhG69rw9cn+trXlWaWh+tp7v5crCbO9x0eZuqoUXNPq6Zw
UAJvbisCMth52kP3xabS9XknSyAlf5xJWRRCrdyJ8Ns+NllbLbvC2WMpLDyJzPZ8
biGUuQ8LFTEleb+a+T7LuZylpLWD2YjYou6b6Wr4RrjIYrggMo4BHsGlLgLYn70J
7DtwqexmXED+IFtvkOhLZumamcqx3AriH73dVCpVPBBGP5JL1ExWZiVgKkM32YbJ
AKKPmFW1Nt0lcJh2jWO95awOvKE+upQRHaMfdX8wafgg0EU/a4+yNjHRABX/y6w4
LkngUy0FrCo0FjSFaZbIcPjn/ABkOIwhYEoAqPXVf6F919E4haVK1bpF2/m6Arr1
54jtxh1NDvBVm12w/7Fie9vlfZppF2k3dLwPEvOVIUwi4T4kWcOqeCJygERlzEnU
pc7HJK9UOj2Y4gmYdwgvsBgyFBBle+TbwP6bSEBhMznNsWKvYa8bC1CJ4Wp2JC+d
pw/PcL86PheQJTEFMoUugf+zMH2lOf+MpPUthmefDnPuLRspWgl7sZfJRgCzZb3b
VhQU89Y0l0DTWyCetXx09z/2FkFIOkiraxyFT4j0n7xa28qavnCWXl8ON2hM6a0v
/psMS06i2en8Rrh3c0RVH3fpNhxdejOON1Al5YQ+YpJv1eZPpN+P/gcYH2P/iaqn
co84BfxTeFidyIUS1FOUW2cvJjZeq4rwYelQFo0IzLh2UVOT6AKP11Q2BXGc+QjZ
4BzYoLcMUktbDust+pwHdiEg7zo1mLpSk37k1a5TgGRff+reV4jwj7/omP0NJxn7
V+naCGx8ajZxXYjAGwqDr0RoHQvS+bxCLyOqcvq7Z7Vw5k/uD3IJnOcNxWl+tQRl
rpuZnozu8FbDjAeDf+/FTGEe1xSfPtjIb8BRw2Sj+EG86URvzlXWhys9fu1S60Jh
zUOPcjwH4SlQkccONjlFwsjAUVctMGdgSZw/t5SCI27YY2MMzrtLP5K2VYGnwH6Y
iQXRtyvLbRkEB4xk0bU5B+CikRQY6PlFaUKYZFwMyQPC7rnIFNBblVR5AMtahV4D
isacZMfvcRYDhGCuX6luYk/y+JIVol3qUrvXrJl/Y26+rvHwuqo3LW6Da8SLevJ6
pnN/+tM6OmIXanvEa1YUisg37PIOOhUK603EZ4DHjnG8VKxMNWCH0xAIIJliOCjr
ZPK9jbFCsXuLW0uuv5JsWlI45NRdhwtQl54LRJTMTsW+mw2cfD8pY4t/kHhmKdSk
6NK6tA0Uq/Pj8dkMnqGbVEb2hueKun5cSWnAHILI59YJ43OBwxysBMPWkImRZNl4
n6xY4V/2fIYPPeLqZiHX3wQ5LVV8NWMDaeS7dM8mgpfZA0kBWuRMwyES7es1/C1d
KTYyp4NpDnqfiMTaM3t9R0YGKJ853PR2J1WlaIwuw2c2fmpcc/Q13AeO5f+hMDlN
AqnKGUr+SMpZ1tJArc/FylgKniDLescSwZwkZNk+qdyZRGxnnT+vQBFW12MIbSVC
lCGkvqfNy9fQNY/YD5dxBS/MQ176hNjxpAv7H103KwQESb0VZXhN/zs/KmPYR8Pm
FQhb1WwN1s6gSr9HnaEkSV+b8K16J5XA+GM+1AwbMR3W245lKXmKj4mxNYZWOHd1
HZA6mmTHLqvuVcVw+kniYA6vxb698x0NPOIoH3tFMtEwFBhP8j2TzmYZ7fBTsZsl
Hjw9jbdc0N6Hvn4M/tRaqsJJ11dqa7L/7Mc9AZYlcE2vqv8F6fNnRBi9tU528SRu
xglsgLhxmYvyP4FxPc9VpvcuunaowlfjYZvJDzyT9T/pkjtghFWjicSHn1O0VG0e
70KQa4K2x8dDD951ILrNBE8EtGttNezeew92co6Y3knK+khqdk9A2ohANZ3S1Xk/
7ZUMuNvUxwk8WITAaYsKInggOwEH3tTBXUB2UAafTJwYl1W6PNhZ4AZygNv6YylN
kyXAPIQ9d7nVQ4c3d/PmvHZ4I0dxOlDO1gvksbPX2BWU9ec51mNaTkKjli25+R7N
jA1wJx3Vi2I3Uwj8P1mhSfDb45764GmVTE/v4YKZUoV+J1iV4XNBkxV2PzSqhEvo
ZwhphKgXHBAkWU6IQCw+EHW6LFqugrW2oKRazuJFRfAgG79go2/MRawlJLW0f440
j+MxQZwowSmwYtP7DvaGbDa4TqZzasuNlxd4wh4gh5OAxCmw/6X5obVYc/2VoOtk
kvHquqdjcyUZkofszTvbq4NFv6bvczrraCnJ+75IKvtsSVSiNay7qUqzWkLP1FFc
YVDtmXsixgczt17WIpkcsN5APhJu+0Oy0ChlZGFoNoTJbWQTCIV1NsxjdpdXHu5o
xJggmTJ9Qx9p1TOnQ953ff5Ain/bWrCDQbhnlGaaGMHXtM5zgNJnrvQ5VZ0S1Wdz
USBnn1LMCu1uLLJQ98Rora2IbtIISoCOOn5+SsF8ED18IbCKSyzcxKTeiYq+irce
BZGUEwUE+k38MBK10FjAkJjhBR3ZW/ilCA7CUPrWK3i1lHu2vMt2afTyYHvVjaGH
GdqQmr0Mt2S4ZnetJtgfpyE+nMgCS9KcspkAzTb1q2QG4ft/Fp7G0mYaWC+rev+P
dlJxIlOW7yFShW6WOmjWtnT5ooX2AK3quJPP7poUueoC1oGYcc3POj4uuP5kE6BW
+nNwD/dGXqzd8MsrdMvrcykTVwmgP/L5hKbwIoocDsOw1fnCkGFlqIpviN94heuN
1iANCBepPR5KT1dXiq0QEvIaJzYWXjqgZEMaEs5+mq8/G2IwKhA0nlUP9bmVaYuh
5TmQfNBsW0kVM5MlE+J8t7Uo7hujT7x7u32DJ1JiJ8cFySfGi4E5Vx9z013JqyzI
SIKZvJiHwduPuUgmla1mVtIjqyWENMla5zCYog1IIh3eacnuE1ie/AO1S6ndR3u5
9vz7+eOi+pVKIPI6lXEFuTeeHn6CN6tgR8H/uy3hanPEq4zFr223ZZEtTokYGs/m
bbuA8h10HOAD522kgP+iZ6M/7yj37Mfj4YKFy4+mLh6MqT7So/Xrk7YM14xFMa78
2PBK/82+gf/W/Jp8eYFx7Z95D4iDOMGtfom7LehmrNyn/31MiLfBgjgEvNHjSdLq
5xOqwsvSbF8c92G5pg/v7YTyibtZZLIz2877qvFVWwsisUmqrzSy2r/eKdvo3x7b
MwgOYmUBc0a9d048dx784qO2i+0qB/55WCqqvi9g8Yfnn88opRm6tpNd+ECh8dBA
648ci/PRlqShpnJ6cIyEC0lEaWdO4mf9UFkXSxvXl4AFkZBo2g0R0kurdeEIKkiK
G/VVCjdMHVgNGDBEN1DmURfqgz0IcwXau6yfIpIE+giE9U+ddgGTjvq3EW/yNFk2
b29lpGkKqCjnUJjt7dlcX6Tu1vc9maADJ5Ep4DonQ9hrLU0Ir9wgzkO0JzYVJhFc
F7ysBc4Hh6a6tFw1HefJx9msQZH9GR6AfCyYjDN8a9ApXz46Z/m06J2YumFnBQFZ
gryUT5byYRVN2Nz44DuV8AGBZuJJtL6RdFSxqz39A0Eojqy/VleWffTV4z9EOWNG
KiukBkxadRi3LyvuNOY1N0INr4HXn3UFodhACRPnrQws3MkMWn35awW8CH93ccFl
SDol1VG2Ik5KOy6UljieyQtOVOIB2WEpjw/G8Fq/FxNxhXw7Qs+mTgZoAyGz0MTg
lQA6/NfIL4yZavLWj24uz/2dXobysnT+rRjWOpCp2RzTBcvgUSw00JDbFH+nGkye
bBH6TDHuBP2AGiy+F70ik5WUVvUJeOqDd2vOm+h2VMZfUyiWndYC7SwhuWcbIvZ9
PtppaJBW1313bBv8cEt4demPQFKzgmD5weS2z0RoMI3uaFYLWFsVpFCPAKrRWiny
TauSoGUmmbxOud9kVeIq3Q4vEoC6pt0dh0sgE2F/fvtUVnwyq4/p6sJBMaBv9rc9
GLd38631UnXBsEpgl/iyM9WkRZ4wt7EHyAyX1LD1jebODp/ygRqg5Uk6rb32F0ez
pHPLPjIwaoq/oqH7U77v1eqDh/G2oDAyRMXwmlY0i/w7SX0GDrvyRu323Madx5jc
6YIzWiIsXkDVldyPUZrGWNRJZrFL0rIEczlD+41b0MLPvgF8HKso4aS1x8kTTjD+
ZgkS2x2MZnZuPZ0hccmUO5go7Fjj8rPrJ9d25WdYCBrDHIhOHkzGNCwJRg7xIeNq
Sd3OLa3/dL2ojMTf5Ly8bKbQStCOKDvNj+9mJo+2mmx+8NAiZ1Qm1wvohnpoQBUw
F3jyuDK9GH8fuw4f5V7lL0wYCzO+/O9KDJRJLPs6Ho3fov4Kz/JN04BjvesGGr0d
SdoQLx/Stpcjp56aLZOIs60vZolgSmnMsrC4IQa5PlplqKDvfyR7HUfstR0rE8hd
8BioT+pNp1fw4DHsv/VqVYERdRLn6bv6mGSk/3MMDSMQE6ggZgQkM6oFa3k1bVon
Qw4m2HSqUxCd0LheZgcJLXnEQPecICYk250JNTsSRcmN4v1uCI9leKvRL9p+a8Ya
BpShNyaIJtN13jahhu+t9KEXUEX0W8f2BH8T0Njcixw+oMZv/Pma/qrmftubFO9i
0p9ZSSQgKb9bo9y3ycDYcaGNioEltiamhTukTyYmn0dqURxCARSaamk2RjI8/GJq
18dyzEzrgWZ4xzp5N6+v8ecLpvu5XLXTsCpJv/b2W+hSK3kz7Kjdre7en5lIBoso
Qqv5JcLLlkxQIOcPsBfv72n8+XtZyuG75LfckEIEFC/5cd6pUZO3fwd6WeGUsZSM
uTIsXYZZ39nAKeOPB3zsqGylIeg1opPpVvI2Aavj7hNsqsSc11wpZd+0W2eKP56G
L+aY4a0bCDwQ5wQw4mZDzw0hyY6rO+EBBXhKwzehGP33YTTPqXIrrTuJW672ukOb
X6DsJSuDKx/J8+ikTcj3qrY3IG2EdMsydv4eqRVCiRoDONVV8scmjufd2zxrnWyb
n6hSmR5m8aIjr8YyxYNC6EjrBl3zOnpb6/5nYq63zi3JN1QeCO8PY9kQm/t2J0MA
+ypAXQ2EqrqDVd4xHyGrV0Lar76jBQhpUSOXhVXEicie+qObAGx/ofANhpO6mD4z
GWL2jby6u5B2iDilhfyiqqQKCrhq/84Em9ox5ozH3LAY8WhGzSxBSySX/ZpIXfLW
74CF4JFnfKQmSfb1QpXM4RmMFr3qsWBxHcm2trcgvioIBV026rCkywBOUFs2fVLf
SF6oBaLwXCkF19yoy0itJhBcdTuRch9CeqIkOH2bh8mXKYkyNwqy6SjR17AddCI4
PlaB2G/ItA0Zy6P7LohLc+QZRGQ6XGgwK+E4w7s2PKqiG86+7xX7AIbHv04GF5Bo
vqMTYt3uzu+GeF509TA9vA52Klmq8G29j+zkBL0F+cSJ1kkf3SU1MAq/uQfXttYT
k13VeLBuPIj1WqR9Gf+luPXldJxDJhs2cAmRKY2cTipzql+ePiG9jV6ebIuZQ4BF
fQSrSLX3ycNmhf0mb/zX3/oQe5ksauRlx+050ERxUXgu+8FWCWvIRBDJ+OMBVI0Y
hpKElee++n9ZiMi24Cj8okVtTk7z5JM5MWmR+gL9OvbCzfuIxvysjZHkVWjdtgiQ
G5fAxRUKlLnbnjx6ibDpdYt/D4UwAjg7jbSmpLSu9ciH1+egG6jrWwuNlKzbJGlA
lXux6wb2HANeCZsDx/p2Kr6Inx2iLP014qa/RGkClPIUBC+bUNLhJlVvDc/GlJIx
K5kGphSAzEMcF9Ing+Rx77GGG9iTbE62ZC7gjDgX5pYeJvLVXKyyDZ0yDWaQIFPJ
fQrIjUc5RqnsS9BRccFXcY6S6DVhDDva6tuF19xmB2VCBaLa8hrdQADbzKTlvOdy
hjv6SLVZdeT0xBJB2EmrgKSwoxlaZI6ntY/1i7mOBeIeq7L5+W6qlzhrqg61jCnp
GUUi2PvC2/itSrr9D7iaTIO2gMLeDUkc5XePZj63AMMMwp/DzQdPtZp4gw841Qvh
yvXPAGS6CXQtYeWESUXEKv2c0i4B/7p3DoyXnRwS7VsoHdbFI3veKd4tKcDxdqFc
qIqOkMdRMlmIwX9l0x8LPReJLlKDJNWJr4BwzNpyymKC0IRzxwGhrY6NXyOno7Ki
AjJMaqqZRJ7NEpH/+juFJbTUzENxpNt0UPEHtZNYR8Zx3cU/lKBY1HcArHaMm2oT
ZuUHsamgAdjcVZftlRT9CwZ/p3jEIbBjk/g2IlPiW5W8ok/EnxkQ9Gtd2nLQJoB0
EnK0a463tSZ6qgkT8LYniwrVhFz4g/K1B2RxDNTabL0OWFKrI5WhR1LSQLK3j9kP
uYuqrxrqKlWaCCkYaod1Y7lXYWLdF4EmYQOQoPk01sa5SULse8rEI5Sbs6E9RX++
EZj9CppvLg/3ZPOGO035tNxRuR8RPNapXzlnp5E0zVW2g+xJga/qb17zlrGe9QtT
I4KPUypfSUffj/WEM1Qe7/J5RkA22BOzGPVCJwVObxteyvipkMJ2Gy8agtK5mz9g
ZrYC3fBsRMy7ju/FimPlFgA5QpMVer11CHJ9wRUckvUWMaV2uZZVmEegj6qa86hU
ho/fL3vDxH/2EeR0534xQREtpxUBZtB2dVwZZwQqjTOl0+NfVQcZEe4lfz7Mz3GB
wG65tEbj1RyUICbSJQr0vEcf1L0Qx4tPq6Z4Ei+qxEB3idy0Nsdj6Ku1b4J3O7/U
IaVgHX5xxFQvODfcEnChZeyMnkmLnDczaVRJDOpvbzZBmEkrQT7C476Aj8zYqABK
yhemFtBBbcNoBuh+rlu+5qDh9pO6jxUiemFacNA7tqbqdhut751CY5JSIvbDPtBI
rLZylnXjK/asaZxkDBwsasGT5+beHyTNwCbteaICWmIQ1rVuoMP/O5sJU2se09ab
ZD58kDOqpIJ4YeB4THK1GiPU+E4CM+IOzyGPUtHWoxYkcnijHLIhpvtmdnqR0mOV
E7Q28y8TTna2F/2QOVg88+DxRUyAOWDdI5KQXo+o/25SaZ3P4yOysxZCeJsK8/Uz
C4K0QtmcdmgNpffrjoWjsAbj/iB0eNXc7KacqPeyLIwDNFL3MFQRpR4ems5Q0HpK
rbVsFVqvTlFRoGFucprIEA4PMcmUS5LoGoQQZ4qKNNDzHNV5rnq0eyX2lxccU8U4
z+kmnfii30dCTaE8tHgGcIg4y7UD/kihbZukHVRht/YynfMMJHPn90YMckGhmuyd
Ftj+AHP4OSPsGCAVVnigTzkPErUVf7mbag9nr6RdmY+zV5oKAD0/9s66qFa/28//
TNYEZiH4WQhQQ8xyOtVsKdSf2jf6FapC1zhL7cadhpRddp7Jt63ummJ5NZOWwjpR
CqIYUt9xgDAwRDlfGueVUr7KderObefsK+pYBTL1ZFPHZb8P3X5Kqq7Qf6j5Syyi
Zl69TrauH9Rp8n6L+jbD07sheAxbcUTexOE50EwhTT1Z4CnHTOxvNdbZJzeMAEdZ
dpcRyDwqEja3OItjOjIkcmkUvcrqPWGVUpbCYHiYkLJTsu6KBGxbIQB/qEkWNgvp
jC27tinrLgqh0TKgN0dzkItwLpYi8Qo742wv8uRr0eCr+k4Cyy96u7ippGUy9ibC
a8ZxWSCETZKvxnVZmbpMACZAs/dYOwIRdwdm3O5PfIdnzILzhe9nA3YvnYeGA1p9
9k2Ur/MLKDdU3rB9FndSWSFKilEYoj6SYob+Dq6mlTbK8J9VyZxCYjbjYCX9W9qU
+HM4QDlEnVIWSl0/QpL9XhPSgHncCgM8amYbxjdnMcCk8k2REVvY2y9Jmih6U/fq
w/hC77T2+/NRCUr3uIKJvcFGjKKbSyNcNyO/6INp7MqoxQE/Hhm1Oq+7thZ968AC
fe7gGTXmAj/zaGh4hAdegY0yeo32Aukd2FIYtEF5q/HiGPSAvJmyTPHPhqQFmc3C
6sfs9+T7tzwljbpfken+bz+Q03wWcUoN2uKVhbOWBycLkQjwrR2GmkBhTbOMv+LL
gv5cHPSgD85uef1YTVXWxj6wI56fm/NYEKwjpMf1ehrTUXMzNNiBctFM5kZU2+sg
5bYReTni4QrCYvFY0vPm1942m9z8/Mghsfwo+mdhM8taC8IubgHOVAjBd2fk145J
dm5NcGnoozETbtlyRbW0sShn0/XPHs5fL6a2qouwATx82t2SX3R7XopWj5XpsO6/
aACoscMUbvzXhYSIVIAI7AN3vf7jApZCCXg6CGRnPW1zJ5ClN0TZFuiWy1ayyYhz
OLDzwJQNFbdfWa4G59hheDUs1hD7/JlyLGg8zTgOJrOrNVYUJ9mGvON82f27J7Xf
NtI9c5mleoLKN3wfvKVYmVWUvO5JyWIFosQOo7g2r2VDDBeaq0b+CGj35FYnCBq3
Os5/LKDay1l7nVtxjIMNJ98810sZy1vmfq5dcT9RZyh92junxMZCTyZT4uHfnshI
YT/2saazLpD8MObfUXliRYAu0yYh+s+e0b4OD1uhcdWII/tNhZ6o+SCr/W56tgZ5
oqIynurds9Ojab8qPDK6fnEBONAZlyAVJauB0AtyMauR4AcP2A+6F4Q1J5pSDLpo
ziESGq0v8cN2xmN84NpAWzwZFAg4gJ7spwc/Qrur5kOVQIMgAcZTDlKL/nA6aY03
AwTfcsbZBXdR7RyHHnVwLtFOvjMKey0O9jefL0l7wxiiz5C9ueKWa9Ru6p1hxpxA
AUiRXTvaeZ7qGRfFzhCQkcH4u8PnimQYQpcqTExUsi1ZY0rABVgUeiwxWLOylaTK
jQYjma+VR9ucCF8JHz+xZxagCGX7kxVK7HsJy/hm0rrpWIS+U7PoN8YPHdO83CPk
CvNqPKCNN1meq0wG7EZKfAf3usCpH1wReCFvJyG/BOkMemhw68WyNMCnM4bxbhF5
po/u2DcGevVH0wPR5yCRVtQHfuhRrNEBDVs0Ylkrq/d/D7b65KVx3/Dqsow7eRkD
D7Ud/Jj7jUBHISOjS3Gyf66VGToaLVgaNcF1d52qU1loqYLAhxZg5+lPnkmi6Ky2
H1V3kxw2wCxJeaMQLP/mmqr4ul7EGXjdQVqN/t7o5Kiw18uBBAeaYVKJLYPKTG2o
A4fipfV6/p4QfgmeIiD4VdC/oynOonJxZCG7EiVlNMUgAHZbl2NgTUxkKpjfjlU2
pS1LNeFcfIsRmHwiYzBw1UItAvM1SAlO0P6jjhqIN14Rep8INeaBPLwCf+4T2Opd
PXuPOJ3arNa0bZDK4wH2VAsSe3z26JtRZGFnLm5Swj2fvRtMj+0LIFiYblGZ+U36
MaOpOX5MBE2ETkoNOaf7lFM1/7FekwMo9lvyyEIwIu9Q/9R8DoBwe2Kvglj5A8AC
KExLU3oczwc9U6Ienqe0uk9oQ3yEf4cSJGAW0SgPBghe5Do4KTE1zBbxd+wxHR5w
gGaf2l1b9115VoQnx+qnlZEKQxRmMIqT1Tg2P5AV2F5DLXI0iEcCOKiw6Bunp8Ja
JSqApze1OQe5OOs6DafyxolVZKiUfh6IcK9q3wVhb/qy8GsGHoxI34sSYs3FEckH
pchfQXyltpAMzZnroQvAnKJLLIkqY/yn9OZKyfZXr6+oCsH/2SZvEjxBwmRWuHtK
6u6nIw4JC5565pPDROIbQ6rxI36FTtxL8K2B+XSoGelLDFw5GWcXw2+aPrmDDsKE
/83AizXn3pwl2Hp2H4U2VxK8T5K2myEP/0FtuYTA/tGljaVjGVl8ikWxhDdDcKk7
Tmv6irLmynABAkfOW8Rz7oURbxGsfOodSBR0WytgNRbIVEbtX8h50B6f/hEC4TVU
BHdj7Ym0ZO13P7R7bSvbI5Wi9Brp2HpweUJlcxqoUx/3xmH6ctdTHl/6jpsGKGxL
QrEEtTrXhX6CM3Do750HEmhuucKlNBjS8vUu5ZFjEHjmU+SNr4vnGR8cmtFQrVTI
GLNJ8uuOB0JlosL8pP3/w63aXti49eJUr9Zp81di9qJ8LFT3fjrB8zjQoCzbPVyK
fXdR8CoGk2UhPNOAbMkK09ZZfqiQddeVRKrIhF4da58n9mzTp1uFIk50DwmCxP1x
z/HSstjsjmSatjttAo6x2mEWXMvF05SFPOb9vBrEtWBj7RKFCN+LsZMMrkrzwhHR
DVCwPt8Nua2pBjWCKZbyVFfSWMzlF5D8pGWzmDuuLmfk6aEKmTZhF5OGDcTxfVI8
5OoptpD4TF0AoRRdxZqhbh7liCNn5ks67F9ix4l/wuZ741ZrPSsd7+N7vNgOtH84
hWhktaQtAaNJ+g+w9T3zrBsfdKkV4HcjBBk5l4IjObRHXHTx41N8CNPKgo1Fk9fi
zKDFGKjSSqX0mJMiTCARR4DOzDVHR8QvxbHhVGCSobYST3EW7j579u7TvLbJ6iSA
ytu9gMUBwBjGZ2kfsfi4IfoqoMSGQ/GpYJWufFeV26PkjCqtDbhEcJXmYHDBHuN9
WFU23SPAepmP62+jRBkx4vVCrTkEK1nfORVNLL3QiTm0cqV/PyEYngFPhWXlwN89
ZAI1Ok2aa1P8h141TgxE+kR/So87vAim3oKtiX89R9O491rhtW+zOcasmN36+xp1
iC7KttWQRzUY7LLDYXfZbu40gYP+RYWS5nj7Qy2ubSLNUh7GsNKOZFIpbfsRM6R+
ktyix/ALevvfGNMbVH4tV8/8q84enfcrSxSqs52P5JRvdyQjEPP5W9q6qKjzX4Qo
D1zxqu7H5tGtj/g/iSVSxW/J2ECCOirBfNCgOv+Kg7nzVjSLSpVZQABuVSwj0qxp
pyAtQ/r2Zgal4TLkVUG+WGvNObRC/rE8NrYtGaiyGstEXdlnHEGmEqML//S5skq/
7DdA3/zcygfAMoosAyUtD8ZbRnqwE6jlxJEU6tlciQAn/BDVs328Gr2cAxjVjMmn
Zl7uK/WquwuWudPGUeDRDSgYfi0x4CqWlQLczHFIR8DBeE8qQqP36bVxNGa8dFQE
a3sMYkt9OC2N8amWehWwUnpeyLzQeHN/oljyXEdROCWOXca4F09i7AkSRAePMQ25
+sRz5SFN/DpP8qZJsgzIdUrFcg+jFse0i7hmLaECRiot96gM6KN78CuiZSjSj4zb
5BJEeksJxPnaR3IFWIn4Yi77+tZ3JbxrClaZqK9GA66lwp0AI9++aQKKmrFNlTDR
C58DZZS+V7zyfRBpm00ytB70gNZRyVHY3Mfc8wUlH1aGnkk59jTCYB/UPRLDszAe
6aUjujChufpz+fze7U/xbohXf/lhfD/5Imw7QyDsnuIc7RJ4mHFsVlXmac2Rf0bi
CDBnUEPoSAXzCOtbGnm6ndhTy8A74I07ZiDjIDwm6G82RfoQw7WmMPU1gebCLB2C
2cbSCuc6MbqMOKxflvduuA4UwfhEUUrQge1Un4dswvs7qAHorlA40WToz23iQ7Yx
npLamlm1rqTHqD2U/vDRw1UXRPuL3jEaBCN06Hn8f2fZ1ogMm7XS8XkbBSjtwDhu
rC0Tcr47HH0g/B4HXwlYv4vjgJ1Z06WHKYZMeVSK4C2UgfAWNx/kU+8EKqG/fdMt
ORud+bH68HV+TeosBzdvTMBRgbHmmkEKRwrcjfnEAoRM61Gu8eplv32tIusTbl66
6ABzUIGqHHIXUuxh0p2cvlM+U+JjjFVp+RaCVBYLOgotS19z2HZJ2XfU8pjBLdup
eyijFR7eQeTnjkAFaTi4nv3c99S9XrZ4k7rOYjpsJ7F1qDji4qPL4Zz/qW0jlkGP
t3aC7EsFGPhk2t+LHKce38TLQDzYWoW3FiF8jw552LgC/Jaus4Ej/G0sWmuzNPtH
eh6u5Uo0FHAlQkFBreh7k/1KwTTe/oqB78GUarP8HBMgt2Mx+/PIKNFPJtpj/A+S
sZSvW6BgRoDhZTk/AKGx8+LTVVDN8GYOJ5MX/hvBeQL9zcFMRNZ6zpWOAz1S3RcL
i95Qqrh9NAORgQLYuAfO0csM+e4FEnFcN9xXkGA2VaXwvK5RuuDJm3FjxITGT1gC
QwCOhOK/+ZDG949JmxTob0bZTm6TZmY3eOlba5uJs/cnDmc+SIJqj3bv67RJKHxd
sWmSARdCCGrcUAOFryJ5JNkrUJWBzlmOFjfjhTyCWfGIQHMRYa8/iJJApgFtCk39
e6ACYN4pw+ovwK9SO6Oum21/2LmmEqSLzvEmkQJBai+rogsTt+yU7ilksCGHrHyT
YAm2fwcPIcDO1ZjRIsz14ghHvatt5GQmJVIEaWejZq+iRcg+cxIrEySTuM8unHSn
hmZI1/7cE8hs8tyLCaP5e9yICKo+ESFIjL7BbhH6F731l0tLbEzYe00+FIkaBXuF
IytGWhgSiQ7ULzm+PfAmhf3I/859Mq6n39a7Ny8qog8lytUswh+cvi5EiYPrvbrl
5jWGHFonFeojYQQMXcqy3/10DzID326ewnnhrN2ymtbcmvDi7FE03A4JIdsXGqi6
awsjPJD4IlLPEWL+34Usog0FElNCpt2qIlaWQ1XvcoXIrwwOk8UkdQkzfTvkg7Ts
6iw5LytpmpfApPnTUctgv95SEN+5EtRcaW84z13Uusp7ZfHfQCLsrgX9shssWE32
h+AufmY7Qs/Mx5rhcLv/qNeCJ4w6x6oietp2oljnXW2nsnqf3r6if6NeSbcfXbcO
Rsp3ndl5UPkvHSvieGkaqThcu9tnUmVxcFQ5W8xbD3wPpJRsq588o8/RReVwo7OB
yZkFXt5tOTfl/AXqDOKCCE0pq1UeklTOpKq7PKRLWYdDnK3OT6GNsslNPhww2ZWk
1+ZQwgF3VgfJlVnDSGJ3uiRrwMR9Tx90c50ujjxX6KYl7WF3ktC3/HdpyD5qfHKJ
91cRngIUdMkUd/1Zry/pwD1hxdccogXpL2Pu/5PzI81aeMvto9dj7UphjmN9X6LI
dk5VE+3/DaFN66lIwv94iHHTPbKkow2Srl7v2BAe7Rz4lBe8S/xASRjovrRp39mH
LWqWzk0DHs075gyCGRY7midWnCGiu3ceabwAMy3ufYARd5PyamfjZkIqA1dmejDR
DaBqTkEs2m8AGBozZTF4qXoTj9R1spRsdP8C7waXHv4UbdjXyJvLmjiTRAqjh/Lz
eiImSpQQfIbz1Nzu19dp+uhQ16CPw21yfLB4etY7bGTOFpK5dEBfiYa33HjGOwDi
1oEbI9tux8Cg7GO/aMWT4qgwUiq9eGXig/AE4nxb6poUHUc2HvCVhnncGbS2q2jy
VrZak/6Gp4UEq3U+hhxH+FXiJ4yUTBWaeUyVkU8GmAUy8lemmZwYfLDPuaLzgCeG
jucGhNZMHDXmd5jDeIXfndBn3BIe1C4IfBRb9bwu+oQU3/Z5Y0GlnCSQYt7zBf1i
Pm8N0wgSYZTQ5CZjeM9bdQ8TjSfkX9HTvs1kV0NsYhpiqyvOMgdAHQn1UUCXOS3X
tTCsxqYPtFzwUQU5zsugs7k5z2O1DryusPjhz2gKKhs/n/TM2tJhI85RdOnIUVy4
Dg1iSAo9RXCHwm5P0k5iQYid8sOpgmGiKQUAG6e0SwkG7GkCXn4vLYUkXCUZHgvf
IGYi0SJ+w/PT3Rd0ftlKFdGEqodQfLyncd40y9VlJJ9fmO5l0c28tZVHpaoUuZJT
rLUVB4y9bZ/RcelpuUTlvD3kkWeHs5QoyJCH3qfG07EuWqibNjMuUhUcys0d1vNr
yTxMV0cPsCctdZ6mGFDPKXj93NuYsMH570/lchmzjW1UboifTNpab/5giGjRgG+z
NFR2YgQlbJJxAFg5W+WoIzi8jWdaP63hBrN/oiuOztWGWfo5/h2BlJi2PJEIGMeW
Hbhjm23WPpekfIq018IF7dpheBV/w9g/8P/FhTf2n/uU3SnQunnYnOdrG4wBvtUO
iqIMF+gJy7x82828OLIUskTASYOrUtYdx5thMx+TzQBq3LDpNg8vVuX3Ty9Jx9JV
iFt7+NcvqtRJYFXoQnQmPI56vCZvOD9iCSvZILO78BJmg0AYPY+V0QrT/ne2RL7T
N+xjOz9ARTH8ENl0SgQweFNJTAeCWX97dxnvOy8S2BIkKgOBVGeJNFOQYX8TbRqx
jXqMO4hEHvGcChzMSGbL2nMURwha37skyvoggKS7hvLVS2Qh1SFzvxqiH7UEk9m/
+NPkFFbp6zTRdKvmZ8W+LISK1ghmYfAvlY1rVvHwqxCJUHYx1Ez7dExtKxg42UZd
EnvajbIVZncW9MKuH2uiqkGyspYFvgj6pNp/OCX0mX8MNilUoXOLJgcnZT1lbdMc
nxQZKyJ98KJlsDgk7Vip406CgRUkEd9NHe/6WQUpMQ7BH1BXWpsuMFuqihDe9Lmz
IaieH48pXtZZpf/10XTZuPQLXDQPC8CwOcCG9kM/1FFeD0MKKwy5o3ejHO5zNNb/
svkbV+kjSvwXrCFF0QpUbilRcjqmLF2hR2syeqI+Tg3JoG1inf+uwGyKZDRfn/Nz
Q1N+qUvMKc0swQ2vi3KrLa+EWOSx7K3GmgUz3oqXBwxKVTZ4j2R9gDHOXbCdfgc5
OtI5XrTlxeC6nQzH6BkVj/fOtKpsiB4rzvFg6gstC2KfHtid3WglmSCuHgZbIX1r
WTxawi1lBjpiKq97/Os9DVXED38EZ53yPeWXkXtWKT1mus5ODk2FV2R+d6EaJK53
1iqO2sA2yKK7p7U+GL4pvyPktey3cPBu/pz0cs4A+mYDU1DGGMbLwg6/w1e9IG6f
Sv8CTvrwD8iFelrDcORtqO9r7nw1ZLUKRiDObIXYgCAMiIUmbIRNzd8bwXxdWTa4
VMz0CFjlJ6v/Tgp7f5nKQeih0tPNuPhOxaS1fefKLFqs/1QFS+9N1uPx7pdmW/XP
f42vyzhqYM4bw9pw4Yhefr5zqzY37qLKva1la3+HaXBEkp4c7kmNLCSG2f8mwfx3
mOsDGoaQD0CGoBSE8DZfzD+SWh4bltHDlPEGwOa5XUPlgPiApLEpCAQ+U/IPznux
8kVX4VqmdtttNkExIfaz0fqabWun44zLeqZiO06pBhdcbUhxj2w9c7LIwvWAH+wq
IY5M5QEMmpdaGtn+Cckbh/yvNT+lrDGB3PrHFkAmkb7DhEM9UHddF2dp6b5WTnn0
vQJkifu1rsDNH0ypWdIYP/CPd8CL3vBKlYzXmDrdnqG4fUErFjACVus9BmRYJds2
dUwBxZoOdxPYlozImVGbF9l8isuXk6xNBdciLKhQmkDB0T25eGeDcJMHOU5HOf7x
qLgtwl7sHxaLFI9DRoGLMePQZqJXK48Z60uH17U/72r8s9LCI3H9Aa/GaMexdhJk
n5hd0cWTWRNiYjO/QySI25LN3WrZaJV3CW949kou5nXgu09GSyAtnDUr9bg+SntR
1KwBY7EWLw9PvuhRG5Loa8RbXycLXAmZ4/mPVmvOCBWLbxIaLhaTIMtxxnob3QB1
d/LRHYrXpQ5iqKWW/8ZxVbjO+ruiyVeFSqnRDLFfnxKMxl4Hbj+jQcWD4gZatXSx
q4hetRM0fFRIiWkHCyFhKac2ZndvSlWl/cZCnW6zRGFSbMFSX8SktY6DVTRYs2eI
we2EkV3Gc383Z416BYr+plKsnHkpe1h7jJN+grJybg0AQYd4DW3V3sZ26uw17fXY
qBejfvVclGyqP/Y4N5YU6bDlCFfay67JlutWPdJsL0f3HZzXrPSKGBJIWSDsk5CE
imERTe9EolCitrcr0vK8gSO5iB3YSOIeeEtcnyc25KdAFSAptL3M0YvQ9HloOWEF
IEiBsTgU313O8tu5oMeIB+1n8AMJ6UEssqAhoWQbdanjbns+PTrN1IcgnLsoRh86
FMsqgAfmUB15NZL59n7TnfbrXyds1JLuCUg3MM8jDUlYfVXSJeb/THd4u/Pnv38h
f3aMVXGp0zeAckiy+2z9lrcqoDINHix00uNHpyBEOzEu4YlGYs9ELloq1bNrAxKl
nOiZqZXny5FxfODUx+0TsZxAVjkxvS4dwkIiMfpQ97B+aWA8+zroi/7GVztSzQC4
MAQDINYohC6RJbjFJOKsjWQKz8q3p7y9alcTMTLXMP44qHCreK5JxEFfZKB6BUDZ
6qvgd+FoZN2WWieIApyFEOoGadTqKo2hLggaPSNcYZJj1GUvL4xb690APp0e9X/j
HH7ZBU5s20+77RBqPR5oP/urF2ZEaTcT7JD5cg+qoBunCrAMhxYRy8Vba+wB/mgK
18w0b1qAEb+cUy+QqCV21osd+6zTvx68kOojIunNspfBhdDy7vp395BcCh9LNU8r
5hVhM6qfJ0RjT1G0NqKcnbMd9g9mzE9guzbjlgJecDb2UteFB379QfD+p5WEEAir
MaskIMFzQDror5BPil7F9R9iB68HaT1rTkqV3KzAz9FLSOpOEpy9JHU00T3S2R6i
CmtxP8eNFm/ASF6npDCdwFG9KY5+8/y3rVSIfuayh18FqrX5gqQdh30DiYw+133S
UJbCUupCDoVWKXODdjC/qpeCcsa2sn7PUonIpjn/n1dzMTpPT6QJZXOHYoLm0nNp
EM67Y1CnXaxULIrnjzNe1w9FjqrLlkSIfOkywGFdm9TW8xe6pupFqZR5PS5AKGWT
LpwIMxDN0W10Ev+PytK/XnQAKy00piDx5HQ64pDSs4H4iM3JUeBK1AjCDOcV4CZg
4Vc1AS9/N1IZpXaiEVHm679DrZopHRPlAAuj8YQ0E8dtuc7Co1fE5OzR1r62PFeI
/c/eaFbuuW3AZGUyZBZmw7hKjM3meWBVMfwueoOSrBXuWwdo2BKpRtsvT3VBuBnD
v8LRt3tBpx0eZnKCkCsQaGYFocjhG/2s7xvXGyKCQ7qFLnCi+eCDm9Kicvwz5/J8
2yl1eVHWhym5iNQm+Yo94MxzE6pTetX9o7WuEf7jm2/e6/9dc74poneDYBgh3vHC
C6mGAP1mCpSYiXyWg38eNQw/TxaIJl9H+wpyzne6J5MqHqfZreSlLqLL8ezEJoCO
86b/cSM813Fl2og+H3BSlXSNlG7k0FgXlipMLXBg07sHcdQX4D0YDjdHNVBn2/pr
K7v1JYBvT8yQ2exl5jy3GDt8HwsY7xPmetiCQpbNXwQqoMUnMB9I3nyDO9kVhiWS
r78qBR8uADmsKdmMXH+Ks06wHvZuaSplT7waE8TX5us9cqoXsO+9SlrXVGeAq3my
zI7Z1k7zbHmv/02ROOPbiCZ2fCIS5on+k5YiUehjnH9tilA4EppZto45J4ueYfC3
PcYIKy5/jcBXHD16Qd1sxlD+1SWqb/bRO+VX7MJYC2SJvE6+yvyoVF8zmJlzA7m5
JHkC4Q97Cu5pHoXSQQa9AI+N5ejgXHXC0yT4yRQup28C735uJJIkipJvoALW/4An
P8a0ExCW/jJVp4TyxEnNzsdufYgwURhWQ/ILS9cFCRFplQzde6GtxwYWwdpapJGZ
xz7LAcZxPRictdYSGucq9ylhBk+4Y2cMyvIGuZeNWzCtLoA+52uvaiK2et46kWze
0/Lu0P1yTkTS04jSfnVy6rlpCsbpfPdW9wt0Vy4NFWBvCnqRLzcy6NTyJIsYGwOc
IXVcCg0yNk1JZQirnJocGzQ3r/NpQD9x5o0RJvx9YaTFvLRtu7nQQcmQ7VBfGFon
TDgEzYmCdp6MLb1JXFkW90W92sgtbV2xDOgewMF6fR3gkOepOmjx+t7htREedsVE
BmnbqirXA3XAFl5r5Kjn2v5t8vHQtIjod/UzA1YSiSr5AJRyY+XG3DOWZz0hwFfO
DfjvT7ZVCppJd527pECSrR2RveyaBoyLVa3aXIKFGolZ/Ow1sZoGYIvkUbU5F2Nl
M7l64FQapFMK2C+NT1/xqiwlmU+D3G4WcJem9v4rb9CUMFOh8ETpbb27uE3I7w86
eBl7ILSoCYxboj6ZfcY2aswSYgmmV8KwpJF6iTM+gaNSPsPjGjrze9gEXYBi1UTj
tsartb+x/zUqOPbhzWL3TdKAF3gp0j7SOthti5um0d19sMoZpAgjcAs4GL7NRWkh
yFWRXkCVeOLrV4IdjCraw7eAmrfujvf94ynidp7Qjy6SwwkphjOihHu0VnO/hW+X
WVuwaHRn34ahhlv804+wVPuGR8BIhPplD5MsTtfrQwQhA8VnReZlZ92Th3mW5R2D
UKw6Jb+6JDqt2m44onkRbOBLQPMcvwsYrD7qc6tD2cwmeyhMhurW6XJpNCYYNbLK
L1bDvDhrgxFVhadFn4m1D1P3gvCYdf2+yznoYPD3hEzsDtWI52rNLqS3YU+vGJuT
fqr7tnjM03E2xVjmsF+zcI7b6DsN9JTP8jAbPXmkedF+GKq3sVM3WjLtOyik6X9t
Xb5GvHLRjDdVXWIEpJdFev7Ediy2MzDxVpiX4MqaTCHxl599FNm0IUhLSwgmYXVK
THn1R+8fkGWYBEesgE7hfbGeQ83yAwYpMcHpfqsz2DvUFFTYMkvKMhtYPK6Q1RN1
SFqfBq10kJWU7/pBdzckOVD0AdfKkMYrqj+CAkKlygvujz5HpI5GhkfE0Pus4PZ7
y91UVAQnii8mqRgXVC4TGtyXNd45QWRzjdb+SFuDvNnD0maQXNjUYMgE0wrNzVYN
SeCjjVZGi4YMUD7c/e5rsVwtUFSPpP+lNiginWGahwnDMQn2ZLvQDTU90rhP1Urr
Sju2akOK003eEYq468/AkQE/V6WpYIfwfF5ieR3AObyQgtWgP4NFNGLHUTLfL7/e
xcBnEv6yVLu7r5z+NRcGpmQ4RAkEQCYN2Y8BkLy6VpXt6du4BOHyuYe5X/VggFeH
KaY+joslq1AKOeg0vg35ydmHUZlcVw+T/Xw/MyVGMAerEJz6cuvZqr//NvURmbCo
9YnEnEugSXTx/Gd1WvqPknnDj1YoDPfj9OSG3O3bqESrE1SKI2QZkegSb0cgwmVD
jUY1zRDQIt0QbSsXqNH0sn+EtauOEqklJ0XitoInvpPqPJpGeOpX8Tac2o9OAVnm
75aBD0JYMhMywsCzD53U1efeT77aok7VOnYRMmr/B2ZCaM/HOMHDu6NjBi9BHSxE
cEpbG6ygkMYkOlOeosZYIUWuWsRhXKAumgE9odhsDdmVTq7s8FlxEOkUTnqU3l+M
KfBLYXqLYyVRMG5Tr4SSfISykQ3CczEoEEj1D1FmaNq4A6uyaE1HUN4T6yLq1RZq
HSv2cgoriytxX5FAhhhzn30sDCbIKDs1qQsHwRqn4bW5exqYBFJSVT/CFIf2JvLz
wXvUc02QlW/dQ6+5reCBCatlZ8qXHKvWlIMmmxqcJgOzFvP8PU2iLNbItHNxnM+0
eeV2BpbgPRzQpcdP4s8f7Sn/PHYRXaqN55Q4hRN1e8OtmvKZZ5823tuZsGkMILgJ
J6Fy9SKkwSyOj/V0h9Ijd4rXFfckNJe8Sv9oWzQgXewKXFLEGt+8eOxdCoOc3RnU
t1XDreGse4q7TOkGFSnHe4JDVlYnVZX6g3yiJ/EKfMUlpUmYHxJbUchXpYW4lqp4
4rqGkicRa0yg6+ZRjHM3tQE437POr1VcIjnug7CPyMcIMFoyi/KngQBa1ftqDsw6
gsQ45kBGOy0ms5rH3CygvE7/OIjkZRgPaNDqHMH2f1Li6UJpDXitOQlbwqts7Bf3
2UW6MjXdaq0LGJjk4SoQM09r1smJGCWiRFtUv1R+Wx/iKVM1URKrXJW1VSXlDdCH
nwYmKYhH2o4Q91iaSpR3aJj08qd1eImt42ZzTgJizI81iNdtkNV5nY77om8IinWF
NTY4CYZJRMWBVsQZlejIP7tyI/vkBWLoGITE5kCfSm6/yFn6AKSFmHau9JWhUtkz
YVBrFLkDFAKNSbZQPtnGyXq/FhpHG4RZhKoU6jmkb4pLVeVaKC0zErtmZf8gXpL3
Ult89SPOxJfaG6DLSN3pjP7AZgkskDPXTGMfkJAj+nqM3vnaBH8uR7MyPLSpBLUV
8U74XLNOX4ZE+zOi+59Mk7beZQwesvqtdMLGA7u5fbPSP2Q+jRfSPxS1Rd1Rn2PQ
5HGPaQ+g2F5f87ibYf3jk0zZ1LOkw3tXNEgR19ySF12mBgyghHkfAZmePJR/JBiU
Td7WhCigIBuGCcB2MiSzlK8/hr53e/v7sleQRV5z16e+S5w6Zw68h5WrVFvc1OTD
EvX2tJPhLBvhDWdOHvZMz5jUnkupGWcrQABub6YigKNiCNcnUdAUgCAZW4ZP2Qho
yZPZM1QwVsxYfhPwYtRBRdByJEmgCt426IcDOL+JjNm7uJcupRZJCXivXDQzapqV
WqYR6NqcFBpjlgkr2xgjOlQp1MlaELz12bYyxe6U2DHJ+Nh/eymSAxblrsZr62xa
pSdtvdP2IFCzHRwNcPLDWyoT2Gp0BANml4K6Co7RNyWoIo9OxxAyjK9O0f9d13ff
8iL38Eb2/t/UAkTGxdpw2nSb+kwzplQZ5pA/OS1sVham35EimU4nhsSH2z41ruMf
lcHGWLfd9xjEdJVoDbQ7JQ26QGb43+tyWhMt2P/Ycvss6785o3ihJIAhayWY7d+Z
tR57M1l3PsuxL9mnCV2Y/oHQuobj2wXW7tuUqKnkVcnFEBw3SO+NMtamN028MEft
2OPJlRMIucKbMAcdO2NrNEOahb8Yy9XnYWh9GPVD/DPe+I+cJ5HtEwExtJTqRHcI
GlsWidFNELfniy3yAyHGKy5CHayMoIThSI4ieq0+bNDFIfrYT25kg2zpuBBVDChy
BOPVQ6Y7ABPOFXd2VqeD1tkm2GNXxPeWsy+9Ju4kRWfWC53/aDu2eYIpkUpZtuPf
CHqx9vKQZXykt1TrFHS5VTbv8jPRORotlIrlmE1r5Ch0gfTaQUWU/mHayRD5+Mr8
vQaGqWy/pDbA7VxwpFl4/7JbC97l9jeQ/XkxLlhLrfGlcB3MSCqZ45iramhXyqUp
nFpg3FBPmBxln8aFRinjytywzmi8v6/UypGxeGktpSMrP1sc7819dfhRZXVnpHit
1IdEnOwRBeWQRyJFuiywFFNXJxzNGHPDlOrZRV6Im2aLxnVLc5DuAUvRSjYt2VJz
OnRfu0aQ/gssLWsAaW2pQOwpj7DH+k02esEl4leNO6lxR9VnFVcGCBA+aPUvP98y
yn/IR6KD0cpjVu9jlYSAPyrhWGEJ1AiW/r5yJ7wuTB/Qww1YGDZA4gBMFpvPiTO0
tieLowxHB2c3uqWGSJfQwrPCCv8I81H/CLC+i+coUVW2m1F/PiQ4XfeINazIT16P
sNWAgjwPaY3Ywt/LTrYGgm+juT83CcF8YUwSu+Ljf1+baykvVFspJWwEko2Dumt7
6F8lvZHTRyDaALAeLTOBEGUeGkMDBsF9PJxommUqridjHAXoXaxTzUXGmTIsUqUQ
XipeVk797KZC6rGLkB3lgRUbo3a6ETS8zNAE/P5Pu76GehXOKObKdYjpyZmn5XgP
nuT1LgXoggdR/GY9sshEeY+6EXkwLdw8YJM+E/IZBnv2e0OTjX75mFpf58nltYHU
nGGrKEbrd+ibt4Z4qgZG1qJG8xvWvL5IBa3PXs74a13cgh5sSb+k5A7fT8FfnHz1
DSEiXYI53B+a35OfgessvoPhUfRHqvRqCoLVDdJOs/895Moof7dBoUWz8VxSko85
kVK3Hh5HQnQKB+BN4k8PR6j548FZv0u9xoSSnqiqvTqFIt63MOTGBDU0nWWAliHD
aNcrIzksYlaEBi2KVEhaWvoDQeX0/wscOH8Px3TbQQ2tHkLjglSjn04OthMC5cJi
fheoZihIo4ctDVVSeEeAqwnOwftnNEvGLwt0dj5mr2gqM1kcq3MAmagKEdmpnzpk
9qIl7HS5VZKgLHHXkEPIC9v2OO009U0390xVhVyymkVctl3Hub9GTkhw+I3GW1Hk
GemaZ8M0XLlcx8MRV9nTTJnXm08fn57xd/CIJjmsvCU5rsmdZmQEMNvh2PhWc5Gq
yydnLUeFd9WFzDjUQUM178CfiZXozveRQhhiNshdM5fLoYt2n6FI1YLPMK3nm78B
qc7p8Llg0JNX0dwgtqkH4atKlQnssgqWDtIp7U2A6jG51IQ73jEwZ1hnSGoJZ8lz
UqtsO7vHe4L45TxwLZ9V9r3Utmra7CBfkEdYzI1LNxacrW7aT1P/WSQdkdot4nYC
RmV+3Gqm6v9JdZqdgYOX8iWoG1LV1xDkLyDDZfkbgoDVQfINK/GSrgDxHwQ6Xo4k
MDCRdpOCKaozqg971A9yF9+8zKT20sQjI5KEkkffhI4f/F2CnGI5/iNtstQW42rD
CSNSRqof/k/2J52wIKc/YF0kIZlWbrB9wChf+ffMt0fdZ5gdTpjF2Gs3eSKOf1bX
qhxgrHlovzchyDHV+6/YQ680KjKX0FZqPF7pyU4F+pxKTbz6Ru44N2BF1+/dhFc/
eUlFcDRK9l8fXtMaJqx/DZZdkbHue/WzaYD/kAzOAgO2JYfgX5jdrJoLXq3q1NxX
f3rV/Jl9vN0SJAC3lakXQt8zBUlzjsOpN8j2AI20nJR0MXtpXOalOkVkVJBos2Ys
u49YdAFwN5RsLAL0j9lpbIiqPoSKlHaF8TWSfkAS4uQlizIiDL63EEE2ni4VDxaM
YypEBpRcpMi2XCpCQwH1Aah7iep+8sAlg57/2PcYylwMJ7bOl2hZK7UAnIquYD3F
3t1C3q8rPJviAAanAfqmOzI8WjS+nBDjXsOxWekMyHPYpAFKvNFLF9ovtnxabnEA
gOSURBXXulLbnz8mjd1/1joGxKtXe0rs6F3NJAkprlQ8Bki0bL04XNgeU9RvZp4E
hu4DCCzq06G2u27kfhZiy7BGRy27FPNqm9a6OnIXma/aSDpZyA7TE2FDA6NGeLMT
k+cqNmRxbkuIlAM/aGxyviCAQaoGBcKfdZsS49gmrMfDKHlwcB1idKS1Nlv+dqrS
+54gwc7q2AoKM2NfmmBFLfxrl1FB/saEoh/1RLdTpsszaURk7/sboP8/IpuZGnHP
IhQUdONyThL0FLCVt6YUyfz3D+Sl6fftOCpj50H3KzBtVHc25KbgLG7wL6R0UrKp
7CrzIWClZSX8srJq5zdXLMhX0Z0612u14xQlPitBdT+OPFQqTr1j64nZlG6Qg3GA
0TGHCFIVx/MoYQ1DR5IygJJTGePD/7yMv2YUijwCwnY3M0Ub7sup/MCesG9eYqHP
Neax7rX0+mtKqIJbtYaqIWH9tGgzdSCVdHowT/d+E7GZ5OE+WktaX7MTdXsHwCqx
Hoj4J6mUBKeHRxhnxuQxWWbq99CmgmtcHi4HI8OkwfDJIB2tk3yQSSGgp9Sadro5
WMsMSi6LDyNy3U1zMOWBPmZ6oX1A26DQHSiqtlL1lUmvkK/D7wOHPatyxFxvtLIt
m4pP9nRX7p9mbWj08KvYGLqOIZLMS6whbvpTtqkKzyEnpgBkme7qxvwS5r9ylki3
TLMeOwtTGcGo4k1kAaKP/92zQbLL8v/zVxPZPNxLNTLLqkoFQsXwG/kKJ9N4sg2N
5QHIsXq/hYz6VXNGxaIi0j7Yp4B6VctfYzAkjWnsFQxZGJ32dO2AHgccMwd+GOv/
3v/XIDwYIpa+613TR8aCCNaO4MiBYdP2anvK4JL340Meserxy87oCdn3tgb7anQK
DI/VO13oHoVGTXHR5e88t5iNAuD1w4eoL+FGHbrsPP+lnRaTjMsPdS+wAw9Amrbx
7A0P67zUhBNrpSSoUWIPUugwpCZH04jPJ3tHcdabmpet1ABoyZQaPhnt29E9HXnZ
VshCGvw9U3Rh8Bn5wxyp3OoiT4YHm17ZLL/zPTNzedb//cLu0y9lzjWToGhF9k8j
JL7UNy0k45NUAFvgEPGR8o9WhZV7T5rEcXWVyMVJJ+wNiEAjB70JlLJZw3R6HskG
Sdare3XSRTwfpHbq/KXnOBfiw7jjMpGmChSZolyLUKqB5hFZNNcqfRxdEZabaYtR
7/ahkJAWXohhpXGBpTupwIyXZzPx5CBXtLj83BJKWt355oxYKhNQlGY3yCcuWi4D
t5XdfioAESjEMAs1AXIDaJUz3kSPdEwvdp3Tzy7WqZpkeLwlreEyjkhfQjhL5cOo
0jj1xtPFhvf1dJaD3O4lMfdiz5K0uIlVqHitqKb7CJ5lN+NalsLkEEsg/HMyGOx6
Vjs7crW5+l8WSFK/aQmaxUhC3rbR+D0Z02WDXwzcBZpOUx9SsWUfVt55bNYNCVFG
6I0RbJREy2ycv/ABvtuBn5LYx6BDpDD34IJvLDkHxOhQvqNyazZx5HwGfzGKWvrg
PeSWBqwifXJzkMiIcxG6JMjVlpUwzdPcKn86YtKSYllOObCWVdlnigJCu3oiupGh
9DybcgeDuLo+H5ibHCY/vQhsc6RgDfrp4fY9QzxuZqkYPH2Z31Iu8b5lrYdaOIZ8
kIUvBc1jBk94yfEmU4Ni/yxa1ieYb+vd6swY0LSyQSSLuAcQWXifRuB374yU2mkW
er5qSuWF/kEC1zg5/O/9lByExrrhPAOVWeOSlSN0rw1ikzfst17ec8WC4yOTNXIX
qbmWjpxL4Ls43R2U6EZrC5raCvoObb42Mu8eWmdS/zo6J6M55HxB6ZCZ36CmB6DF
nuemS+MxGkwaKW1Y0UYa7ilJ/XBJGUXlVr2H2dBzCiLAolv+S4VkfNnjBR89mxdC
PuMFZPRk9cA30sWkMjeimd4IazHpNmDr02Erutc6NFAl5fh7gjDjsWVj11AfDI4E
axt5aBEEAqKRva6tfKcABV8NxcoWgxCKqM40rBlCMffTYOehMQ/KF6ZPdOHPV35d
INMnAU2+NRT412J1eKZ0K4N8kvwzpNeAnBnciWU84NAwbIZBUIqw2uBzymklwnNN
qkqcvO5ZAaJWa+8JL/ReUa0PWGOVBUlnA69MlVGd0MFcokPW1j/jaFTwvFmMgG8D
K7u8rVtmeTCceySxQgOErx8/qWZHIMdJKad1kBZMIowhmKF1yR3DhLq9I0SUrUfF
CF4anfqUCLCQ0m6eYb7mcuUdnr/gXA3DCXFVrE4pqGC+pLCt+FQ7DjxMD3d0TV5a
oZ6WM9jD6O0GfZbPVreEIGgfY3gqdEReAGbsujHCmgYvHD/fss2/3EOsF5GhCSx+
a4HJAT3o5E9OriFgnX78xVO5V6/KlrFliMejavaSn3O8dO8v9uL86+OjPTT6MQTN
cxoFxrALlHhgXN3mop2ox8eN74EPIjRNG66rZc6UfymTeHdtNRZ//L4jdS0O/KO9
XyCF6K1q8HHtA1TI6I/5CG6LPHDIY+dUT4LEoSsbQePd9BINXPwbGnhOzeWMwfSJ
KewxSHvj2w03TmUQDnlk+Yq+KTVjE53/TX7oUwpje/JEH0IH9TbCnYnC2KYPdjEf
Pf9lXopCJvNkSb92NG0CpbxdauUEf6LfUtatTULsnJlw8uYx7GZr8hHUpTEsFSR3
lIng4ysxrIvZoTfoyASclAXSibbBW4hiT8hJtmJj3RBbjfPizWNH8vU+qvadmlkM
X4iM6nvmbWCFcfbDig/vWyAiOEolBiqmqPV+dFA8R+WAbXeCYwtacGgOibHgOhGX
zsPRQIN65A4Xv2jodHpZRsHIAJIbrheW+tJFhkHGkxGwavXhqyYRenCKi31hlkEb
cbZ7jD25XSIt/Wl4gHnH/FgXDhgsBu5XEu97xDaR1ReVZngd54U6D6974mTex/I5
YhBLyi3FSecqsn8EGVfT+xX5vsPi9Ehtbqp/zCaX5iT0Eoq1ry/6rgdqIv7uiJYt
t/9rWxOnNOhxdgW+T5Xd8ZCQ57KosqVCW5Yfhb1RgDoHnxJDVAQisTnBn6+alCzJ
7zVpYJwYQk1W/Vl6PYqYtuuiCXtN7SJ21YS5iUIJbK2bUtIoOa/atsoKmLPZDpvD
o6wnrqmFPXwCn6hOWQTqj53K6kiIDJQRrj5JXygIDi81NPTyPw/ZRPhB7GVFkzlI
dsLB5Q9oNXfwLePPCTGk9KNhzWfTaG1rUa1PkdfXsen2hkSiuRt3uR3dNoBVVjcX
qYOa3o/yjfsp4cMsRXMocTLcHEcdj4+SPnj7th6NduC9Ia3t5LGt1oV2m7Bo7KZK
km8dHf4W+pUYgd6sMMG1ayDSGJc2LzzgntkHU5t6SEvyDsbvU9Js8lyMDO6VmE+Z
GfFvPK1flGmmJgLZvPKAoggpCIlC9qAq3FR66sPGXxgiybDCfwfmEVGpf8cFD7Q/
3ktIV6t7/Gg8n+AxYEo6alYN0TKrS0dp55EvgcJzFUPxBDSl77wfjdHvLHEqSexx
J1g/CaOG545twedgJaz6h8lNwOlFsp7p2wsJa18AL+FbXWaeo7/ldXmshm4QmHJr
6/lQIcAKzdXXn/l4EnvoPimhieV7CxSecLJRcs9ipJMQgDi7vNWlPFY20aoee5dk
Ozo3k3JYX5+X4jTPuHt8AxMmcRPYMwJvLXK0pClvfl+0rZdNyyLO5A6qjnUytOWJ
BXpYF+RB/edE7Hk+vdlIkaGc0kYtCqYYfJi+JIkl0PS/xxkd2rsiuWZ73/TFgzPt
qPHGput9nikZyygAksD0ov8IGdzJ3YI3Mg1mudr9mS9jkNqGovfPQaV2vBL1rW6b
+EFrd4k4G8XTpwbHoWd5l81BJgQs9GGYY7YOQhpBpj1atOGuhH7no03cTF//JeB4
/WFUIgWfjhXqa9e3fygCjyeB9s41BeyspldRyhxmBmsV/frMzvIUncBh0jxz3mM5
PjymPIWAD7baQudWTWw4k54d6IYokqlNpx7S3Aei6q1fyBoR0o7kSbm4gR0HuOLp
GE1osJcBuAHYG9Ritczja9d6D9+WqRKzH4/AgYhRSowLozlA6ceMyfoRFknO1UdK
y+2KoKIOpvgoT3CSGu7+1KZ98ec309VfVEmMoAcfpP8llBm/UoMT/jEDcginiUPQ
HWMC6ahv2/uK/WAZih0KcQlrn3QDlnm18hE1DRiFH2vB3GnvpPToz0LR8KrtVzb/
APgOwmKughaKn/JybDbVrLEeiD8OMaA4+a+uWZ+5vE9v1RKaa3Vt7TPesIJhEdFU
BmZFHnCCgI9xPJBrMVJVB1/PdMxgPxxJXIjhy2UEFg8X0AuJ5lebxhFlxrAWk34H
WKUmevcfddo0ClkmvU7g3Bq6N4uTmIJg5zMH/kQfu7be5Pa+XkxoOjRhKglPc461
YSjpWGCu/jQOMcLYT9UJsj7rw9BxBoibJZA9cg9Pp2D2RmrJPZqMkQRgmrEGCQv1
VeCoBuOJyWVxkDCkRJHmwS3ADYMIGnvFy7m3CRSAva9XgaeGGJnA6KrOi1nBHU+k
eHZdLHAqVfFoEAO+16M6fDAhycfbb6deUxyYX4njTMuS2Rrfr6YPFv7ug8KxTBMM
Ix1MVML0jTnQKq21IStrrgztGXLWQe1xX5UJWzXeHPqwSmzcrJOozmCKzKzGweLP
eTfIIVvfJBB2sF5ltW3CfyldfhbC8A/Ylqfl2YouPmv9vqKajoNv9NxZomuGitf2
4dGEVmiBp7RbLZL1pqX4GumdPn56NpOSuJH10M1MBBmqF+BHhJroLwpihamDmtsY
GcbGC83dNgipj4TKxT4TJuXPWpzjOLXYL7Xl5l6jSiMU7CGhtijtIgSY10o8iQMg
oS5KqKz/9UZxpul6mcOTGy58MOX8Bs7Lc78gHQQBC/BjB5rMPMkOo11ZBkA8j4S3
NnbJ+fqaI4v9KYEobDoBTqQR9tD8VM5y9WO6dJhg2Ww228N2H4sChTJMuwD0s7hl
I/9oMVQ8SAVa2x5Mmsg2pCwTs7HzCTXL6d9UN8zbEJnk1QDvtdww2nl3iz0iHoOz
T9RpjLwnYcfkgS9aOIa81ZEevwmJR0uCZCMZhPRul8cCkIBKMuvGXINIyjRKCbFs
da8Dk9/N5Ssggy5kMzY7S0B3MhPkCNgeHymKog4lUz2k06yUeQkUJLvJ9n0FxW+w
ITRyN9LwQkhV7vkEXK9mfB4/yWH9ypim3ZhjJ4dpFdu5CRk3h7a9fnC6thbheMD+
+mjMYo312g4Aq7e0HzZP+hN+10nTTkHvV8160wUVo8mmnj0Yi7ItBwD+qYf2lciZ
GCtR24BR5n0jPKTlvtQOALHwwWSFpOITl6B1EsFJR2dTNl2Rxe3tcOZXr9ti1tNA
/sFtI+VGZ5ibvI8sQramcuR6WF1YKYONIlfd0yTJhp2YT18EAkgqsgOLd7inkLFC
WGURFBz3uP/2H64+J2MVTkRPjBl+8VFziDJsugDoo8VH+LrPZGCwkJyS0yzGK+2/
SibpY/EJ1dytLFknAK/szmX8KpHHvyCHkpCzGwm2TfiaHGGY5oLdCKhWvg2NFZiH
J4khxzlkvic6Zu68GXpjUsgFfmc7BZaLxFxoJ0EqpS2U9mza5m3qRWpoLzhfNCT8
29xOwC+2oazu8aLGkz3d0os2H/Z8mahNPlSNoNfniGiIR1oHHXzapEig8dvVE6ug
ZlNJBHLhuNyOg/ewwGWdMUIYN6PInFWsWE2VeyJWolv+Z3GdfDPc04BWCfzGP9rg
r5lhd1QjxVUsVbDtoJB7ecDCt9tNmGX32X174xPvHc4ZMO+DWpiD5vpV58Ci224O
tDQ+TlR2tH4R1cqv2aO5ZJrKgTk9+ZJpFE7BdY7Sr2nEO+dS5bmzROBCeyarj0YL
Cy2nSuMlaywjGPZb/YVuIdfzrPplSLZoJixIhkhwxNhy7sSfxJeLJSfBrHk5aOES
HwJub/yxxYXUWaH9VDNesQg8uxHYElFUEVMaDefDXtyVqOz3cBIPShIWiCfeH/LT
i+EWrjJJczWqDRAvD/59Plfybm2JopA+LGCOBfIWXmfTy8OzUNd/d57oyu7hk3xi
OhCYuXtYSnF9kWXllCeEtyBrBQizTFrU8DCnj0EDQICnZRII4mKR6rF2kxNH7lDd
W36xGh0Kb4jzQUumisUZk7gmxVLDCC5vc5qdZYcWnZieL2aLKRTWMASUjVrFrWBd
ZruEU+Bqpsp9GtZRyff70LTWfunOrKJgeHyWSbHL7roXYSR24uSXmNY0LPOH4QUB
nvHUGn8FjYnkWfYzoXUZOmbmgwG9i610mjC772LNGwxupPcXVRQ6MQdJAEsY73GN
zerIT1jy8aTSDZsd5yd8i1xIUlD0yRntbnqA8BqQQ/C+XEwNmQtBbtjXaGaux3XK
STEi3ACpbE9jHVKvcEzSrXz7VWSbV92JBabYyxrLl8ab/Ne5olhnTDZyKrBWoO72
WyrHTAh4Q7fmA9ACB5HlVhv/nPvOjAaHTocKr97PqSH87BLXuEdDo4mS37qtOLJO
qx2LHDnCgff/IqtxDNDOo15LVhEV9bwrY6bYLmFsOq4h6G/cZxnlI7K34SbH5Ug+
w2SrGhebspZblkJshvPTrp7hMI0me7kXXmsEpbvexqQtkx8CdfnT2/fbi84hxMUa
rrnTLaDwWd1Wr6utF1nlwhzt6nSrHXilJZ6hIcCgJ7sapEdTo2mufekS30QU1ZhD
nwCTShKypQsIQESMQEKbPA1gZCWxFBgknGkwlsAicZ1FWhCGCnuGErznHushDfyO
dksWksRVy2Xz3DdOZb0Es238xydFYiV3CwDQNx09B3/Gg7jd2qMvUKB3m8OLqZz7
iTfZeRk/g+fNGU2Eo9pNq0eIahW+ba5QCEslY8LxK0djBeYyryabhSxqLC8fBLvk
xyCyyKH5JVZTFR7Z/Da4D3QwFGDIY4+gqORy1++8N/VbBM3SBZqHGqkaw4PjM2Fa
T6Uxzmy5pOLgI35nE7dnkduNKkZGbbotn2r3AchJsFpIWTWL0vx8xB8kevvo4c/g
NlS5ZcDpj+qKNGkQCeVQDUCO4JmajabeH6D2zIQ1HMKvHuDnlV/0LChqgG2JrlsJ
yOpDrRq3+RlSsQF4qS5uc4fpxzEOvAXXazmnXN6WnzTwC2k1qnGk8kCFnjepVMFz
zpxCtr8rdcmYpva9Fx4kkCBao/QtOugHLTAk2hnAg7l+aclj8ygNIn70v3DEkN+z
1/98PTwz1Y1WsYzxlMVpbTwd0GSAy2CXVZD0B3qSIi+Ffi0vGScofeShre0Ksqs1
DJAtuNC8sZtpb5jW/dbcQqTVECV8NCRjyCMMdB3DwM1u16nsKioppFBnRC1PNDIa
ECtKDWKEfGlSgdO5JYR2DTqiUtMsnN9uQsWTMydHGePry8OzrKCKckhNMDjiUK2K
boflFfTn4KlFtQC4fs/ZOD4XFijxAhKksjNXsFI5oJH+WS0b+5jMwwiV8Iysxnzl
5v1T5IlmUNCyCNVrIFPssZu8bRxqFhLbNzzwoLBIcOSkAc/xRfmtAO0FZQGDX5/x
3ZTPQc7LC2CQOK4nBYdatx/rWs+U++SDwnMLSqz9XK/8HYWHiZ10LdUvzfJKQCqh
q04WtJRilwtRNV/OrCTYqprQltZ8WVKg0iL5NAhO+AXLXXiNCFUgZmK478XsMbX3
zjazyUVWbhf9v9qH/qgcKJsfBtu8J01buaP2P46mMb+N3FFgxIkVbO3VrTgKiWLy
q+ldFU87uPrtfq/7AEqcJDJQlBaCui9YntC1qV4L7gD4B1g+vfej/8b/wUT1cJNM
/F3CzLrhH6sBmSFx8ghYbDo2HpnV4GYqRGTCtoURoTd+nIGh9nk+9YQ+suO3caBv
x5Zb8VTJ67blvm0FiEsWhrn1MuPE7Jt3Wq1GSvR0lkiksKDDXfkScEbVdgDFnLkq
yNhdRhrv6FabjRMeIVHO810PMsLNcDGZq4j8eBepCTuclV1gqCHws9bKh5iYR/bx
6JSppnmVJMzjKnqOeC045P9hWZow5Z37aep5xlWj+wbl/MFifParBfFzRaZpmVMT
E6a2aNzvKbq82+C7HwzGv+wH8B2DnlI/huyZYoTvxCirWbL6go7Ps3UsUTF3Zvyt
gzplhXElK/z+gyhiLYralVy2diilgkpecHerum/bKvyzQCLJTG8o9Zbtx0mj6P/z
c2m8b6K+SSYi4FHfo5j+nLDAK7KPPhjl+zC0+ucCxzCoEOozRWCdOjDMRuHTddm4
t56WVuifZeKlPjwDk+uvyTHXsgh9KUyfdvZpMmFSqQQeglJgyQxuvoAfL7iUv+Ch
tPVS0dM9Yd8DwmMwVAkv+k4Ai9gytl5FkzsQdb7IHe93Xm/EjhyWnZjpmZCXbeSj
EbZgK4wf141rrBlhpppvUsIqHKAnNTy6+2P5UCz5h27xM7DMI93e95zIyk9xDcGh
cygLy+cuq6Jzg58Ersm5zbKd2MmvdOhNKEVgz22vimCnvNGSOnVnDXb+h4AA6QVo
HWVMACeSy4Fo078rrWZDKEeZSRiQhC3dnjomFKerNQIgfUBrD8JCpoZ0Pq4EVPjl
MsKtD3QBxQJopXVcEe39uAstiSfPBmzJlvAONZch278iURZzoD7IZyoLLpcjdP36
zM4txUSz3oPS+Rzgxb9iDi+Kd1IZjXP6NcN4VBvat3IDPv8XudGyTuqKJ7lLupW9
YTs4wJEUUdgH5NuiJZvIaIWAz6M9/9iW4VjguUVO+yRuiYQ4087F2sEzhdvgZzZW
J6j+cLc6f2fy7ciKJk2UVwuEXn+Hn/UcpG5iQ47FZt3VGzgoXtAQVee4tGxLzvk4
uqmUBvRASmv2XOipJSsom8lDCaaCJ+42ytz8vAl8aV3TVrnVAC+vXbKIGMjzFOaE
uzZK2IvAE+ZNakiR5lN2iINAdIcgTcc5pWxxpfbJbQWwJnO06Vg5dJErsP5OU3Mu
MkbV0Sc7w5aIfqNvZsuEjVi+vd7eQ7EOZWSKZMXCH9G29gx6kyKOSlx9UsxWLyp9
503eWzvR7X1gFZsuVk1wYSMzzsgB1LsiHBE1ClmLq4r9Qs63lQQCm7cnx1bGIaMu
SKJcAy8uwIy8bEAbHjWnsOMQKAzizUbWtyTayDVo3nH/3Q0N/KdGno7DuXJMjheN
ZVVrURiVyTpsbf4c02dc0ZyLCsTbeQg5+FBOuvSJn1dGjXDg5mwCbfm/VxZuEEAe
KhviFvMXj/6dZbBxrn/F9PgiXZ2Fuf1IU6CVq6XfStKnCcF+CylL1EW/j3FhwngN
fhSpHgozgB5AbKyrmrwk56tbiGcQ839mv3Tkf/+wR0q43C0Gddlka4JIotQVnZxA
1FQM1JHAsGsI5wrpcYrCqJ9j1wTy8D3fNZX5qqg19AnwIKWcMmbI3HQc/dSlN3DE
XsDfYICbQjJspQhU7x8v2cBhm2XXnBqVCn/gm9/pkVBXGkkwtFXC8gr4GNXQBtML
GWwoKwTs8WF6xLxZCyTNWfhV21DeDgS3fSAuWQgCcBn4tYuwZgrU8ItyYCvHB8o2
JISqArL1PSw6/zr1beLD/eoiTw8k+jZxVQKIWtMw4h8cyRql8ltZscBzh9muBump
IkgHFWfFcNubmyAU6Jjukji81D3nXY/hVv7GBmo37SzoPLJVCpDvgIm35ABdzxji
46uhtqkVVRdPGipXO7UdGDalNQCxVxRA0RXhIEkQOwIDzcza/ym14IJHxLqUv5NS
prB9JYdQWJvBhqrY4jij3xOdv+RD03SF8bveXkRb7hNFEK1xZ2b5lCbIW/pV15pM
agCAJLF7pizLNNw+odzza1qT3AcziSAiPYq9mifBT3pimU6G/TtvL71vK/BC9tO1
vDX4hg7anh8L0z2ZcrzxsaoPGYbFZbndxv/hPN5KQQh+1hLadfjbZ/Qd0OlR24qU
bMJefYdOqE9Yo4/PoBot1GphmQwYXVhdiJG8rH+YkIWSbvlKV8rOrP1dRSHLpAIT
ZvjmTNoDmBWrjLTnQ8W5ZymB2h9/TKRLICbgQN4V4lNW6W9nKghYV438z57HfBEV
jJb2DfoCM1N+iy9+U1UhLDMpd9HxrwYGy/Vvn/+QTzSB7tLhkFWEHFWqWZ5QYF6o
s/DjAKmAsgC18qbLALH6pq6Cvn19f+nVn0SLStgwBO7h/jsace4UUMfqWOG4Pbjg
SR5F4cJxSfz8QSukKfgrpf5NX5t/2k91USj28qscM7C9sP9em8OMPOdj1rZZ1hmY
rZKsMoZU7LlfY+ti9mR51IQFNqXAVjpB/TVI4B2lgXF340PASpvr9E7HsWodS4xL
NwoSUD5ddj5SRvLtAjR2Q/xUIMN1f4LHfbjWgt34f/w7GbHPGCZtdHKrlWMnxkba
cTq9gALYAVhJ2Jcy3DZLuD3aJGuT13raClmwd75anqGRVjFWl5Tq/EBe63QIIjuv
mlDpflmhmIbpnm7n0J/f93/LubjRusAP5Bb92Fqypk76tI0phdzVpWgbyjQUPikG
Tw/r90bRHf6qX2AxNfxO8fRjnuCCO6dKZgRv2fEi1BxDhG94st/s6PVduKhWHgxs
SfJvn1LyClTk/CQfDetwvywqyqDdUTa6T5UCFLTu55ivfkPvvT9VuQPXuQ1uoDhq
w3cNz/sraQlES3fFRyzIaTEJd/eeHdn3nuEkz0XtV4yr16z7orb/fNi/YZxVTT+2
qZb7tsGjCNwm1g6zydZ6jNoePsSu0U0O+29TGV7qB21+ajEocsVCE1IYb+xRfgMv
hKrCoOFBrs4UEKsox1LrISQzamXI7Xp1WUiA8glCrK4xSnkgGQOFne7SWXEBHwcP
rF4aeOAjuq79ygR91W1b2RF+puPKIX0vQDAnJ2GcgxNeaDrxP0neJGQdThr70P9U
JhqwgobVIlFEi68aaCL2bPlvGz2bfwmDX/mHj+TrupSVqSPjupOZJt+pQ2e66h53
zoztcBbeeLb3dyahNREWvFvY287GQ3Y6M4TlVl4iXJrrXXlDdGPL0NBKsTExrC0g
wzvlvTROiyMrE6Q6K3vO0+HTMHcSFawYr/IHD46h3Yt3J5Am7QsNtdXATkack+JK
W0FwiinO8XxNa5TZsiElFYB3pw1b0jf7fmzIIC0E3NP5e2tie2MFj1USPIECfuYk
Q+hozjISELrkAtNAL0vo1+G4cI3OShIggDqH3CJaBbdJB4QJdQoa5o+T98lDdszz
qFVaI02yNfKAzFIA7p2cszgkjijv7bUtK6zFE+ym7K4lPFU7IClYsfe2+7JvptWH
m3s2a/7kZEp/TaWv3hMjoguRqaTji8f5uIVLVbQr6uUFlVQWTZCnjqCZWHzgHTxk
QHofW8iAoxXR09SkS89odv0QGeBsWX1CnTDuv/mi5XJ+PASEryJpA3JBeX4IBadB
EN+IC6JEL3lhLYx6PRsipttjcFU2/mxVSYpp7I/jJuFoqpBpoXyPw6MkykFVlR+1
byG6cqfh/tAtW+RlEtFmPzvkrNbP07C6qTW56LRlhKwa/oNJPM6ARXx9T1FPjxGF
dfZo+/vAGApuLT/qX/jmwlIuDgDUbjbYanuSa0pDYB8DKauy2tLqmtZAIf6RFEOP
rAfNA5KLJIZKtOqwan7XHALZZvWrC3NrjIRc2/RkF0M75kcKwhGs+BJvWd9KEgY8
VD28UZ9tsC9QmzOQDLgvEPfOLjB35IRBwkheuIyICbcR0KEEYQFbQRoyM217tKd7
AgMy4V9djkmSnTZ+C1mhPgCVQCD2dyEYIzFp5qzxdpmLLVIBMbUC5KKMw4Wmqwcv
/Y7rgNeFrsRroAnvaIPotMdVrlPb04BhoT96y15mHU9CSbBd1vEAntrOcYH7b5Hz
nsXUtiBVScawvXWn5HabAESc8IeSh9H/TBmKwB7+nzD00VmjY+pssnCueMH3mW8m
iioxMm8yluInlmV+SuMlQeZNMZ00qrgQdfxubLYxoEWeyLLTnnY5FstiFseCM9zY
H61kzeW0W+79eV9pTyS+ZHGSYlHBbyl+Ghx0IOTrBrvTil6eoaLCExLzlMDyWI6U
GaY+BPdm2W+BkIOdFaum24h5MWqCOhAHnzhGOVOkKFifGl7lisOjGXtcTHlJB1eY
as8KZPPJYbw8FOF1ORCzSTzXbNtg4kNsemJ+OPudIKgRtZ7SqQNVnwhdI6dznbcI
AF2uMxEPSu7Ft9KqJTBVRiGtpQhY+f8XuPa6xkWXYCpKvHazzBYd5ELqFzM4aban
wumliRbHUaOyTXczo+yW5V5rLQlJ1ryWI9nz68ooouut3mEQQYLRu7el1E6F5EAC
Tty9IwxxXQq6YH5Ehxhn7kpdp+Rc0VJ9jf/PK6WrE06ycrQpl2bcGWQDM15CKu8U
eIuD8vR+dZOqOcC3aGyfoXxhSS9ENkVVc63IrKrlv3jltPI8vFi7IoNLmZDqfwDn
RrFfv6ru2+lwBaNfaJFlMN6qf+Ez3lhO83KR7598x2MgNLG5/FzS++AiB/o2kWBI
T4gbDfSqfxoP3Wf/lydFPy40yrv3Mz3BSBqtRIJ96BbchKHvWpVRPC3v2LtrmkjX
fqUc+TujI3fO3M6FqoJyS/QmFCaDCH/AAqNAxCd9rkTlkFYjpIcu3A9fSGIsdlWU
zmYfJL4q7oZhh6UXOBTIfvkfSaMKCQxxH6GTEjemhKBu8dJs8LtS3nQhtnp95bJE
4UsuI6Z/NXKagDgDTX/HmpMX71WTmEptr4AbiBZQW5LfpIvTb6NgtZmc2uL4aP9p
9EVH6ci8CxhBx9SUSC4QF6dvBhfLIv7da1sX9/08gUDZ9c7nMdYlTUAKwfhDCMwn
e33fi/Wpy55S8K3yr9r5jos4HmuPTUHV11FB5kTFbSsAiEXCfArDDcqH5FHwnBa7
eOLKMzdx+Rhr3tJzkbC7yxn3gwhcfdMJP8oU2J7LbpWwFjk0ZA3ThXZ3jbqBHFlK
xMsqTgA4g2Ta3+ZaKWBgrUFSoKVoCO1Y+7ATEalEGWFL8M8g/jGR7KtQN7v2OOOR
D6rr6m4hN5WMmLKgrIqHj3QFjz+jQGYhZyKUahPs0sBR9FUvkr+wv8KuN5h6RpjB
aqgNu2wnAto6CZclG8V0dHDDH/7bYmdKYXg6rd1bAsvQ+9lUQp93PokJIOPJNhvF
eC2zMCAYRE9VraFTQnWtqKWQu4L0PODOrv4zKfkTmCHmc0m96hwZ22n6NOesbp5l
l8JHYC6Fyq+FdoJG+wRDctETevME3PgzCm35tZWZRe/V5EtA55vCEN2D+rTL+hfO
Yn9s7WPi+KiLP2Q2/udfNKuUxCjkXUcXO/i1GAtwBsAfpXkysvqWRZ8G/EzzhSIe
zcSYeE41KXBgzCRdnyOkyXPkA+NpyoZqaLPZbhNDO9AcOXn7ecp10PP+88V4GJqI
VhMaPrMJbitTeT6NsNjF2xHyIdDUcxf9H/ParIaZ6v5rNX1dP7Hz70oIwzv8fIYT
OCpH9lo7/CSeKItCUZKXL+Aw7nnEEhYQ+QkpHPWx0+qTPY6pX5Hw1W3aYsoob1mo
ufz1u8ICOYbR1/R7jDS3gK7JOYNvVcQwpBYaQSTtIHLe4E8MzQKzQVxIvLLMpvYz
Y7M7zV7xE4MMTGzAu6nXad2f2gtbd+Q+CIy4BhvWxuY7ZtHnu8HskQQ/SwYuNenw
IlXH0usfzHJaI9K3iHvglxKWuYFWNUDeLY3myvitri/CqvhPERjc+qecYUEWzMuq
FrK5Wng2o7PCSMr8Zw9IEr2J+WaYVU5buGMnace+NcFk96LQ2WxQCEqTemuHi/mv
9zOgUXOTLgZ8ViNYYjOUW2If5+RbWArlxvD52bO1n9EnGMBx3ul0lmJI9+a/Bp9V
y71tAabNzzZHyG4BleGxG2JafEu57yb9DiPteRZePuwp+W7Fvw6JGympGGG7S1VK
03GDDiof5ueQBcvX7juCP08Bt5ke8IY1c++3exYigkS0+LSacBDqsElHeiBCzoIB
oGiBnkQXp2EGaaJYRMzuE61JVmGA9irCr9yRWUyKnP2vRRrfAHCM1nuop3Y79Lwu
lCgwdIwEg5oWl1bCKeWxH8nUQo5ctkMruTnzLRd1OodhH87pilig8w/oHCfnIa+J
si6l8sR5TQbMGxLo22jLXOt9Alq1dVyuIlMCNpSQmNLja5+iPMlZKsJecvJNx4wK
JPAMKO3LhrQKT/mQwauK7QvoM6QhETIU4kxlGsZKHYfdy7hnalNuVoLpeqJ4Xucq
eI2xoKindU1XAhpyD1xfoTsM6bP67TKMmB6pawdO4PXWIcJ1vXkWBK9MWR1PDpyh
uy8h6bxe/fvxUdpwBbQ94qGHjpxmer8aZUAdStd8X3bwgYVsMbMPloZ3jvkhE/eG
e0aQnw3N6mN/QlM6/Jk532Ryg4nOSQRrFZHx4RwFsnTv/Qcgesd5yukr7ABYGkTd
clZOExGM9CcIejQULvGu+h4cB3qzhLuUucGyosmI8mTS+T7DkDzOkFKGjwKwe56w
WJV2ZnBK1m58FFGQ4liVd4ck6jH4h8wvyGgk54RLBo1do6FOdwwxtFsgZMYx4h1j
23wxAE5V9OLO+UWcdaO26qDeOyvPkXmkRhAXXN7z6X/u6BsRkY4qq25BEMTzSag8
o/OBY25qlX0fQCuRWXu9uAU8KM9HArRQWFUUEr6bll/ewNLcUuWxg015ITz1Fhmc
7JrZUK7RMm+9m9lCMW4dMylMYZO2NtQHqkujjg4FZAElY9XmRruhAxWX5uqGd5NO
b7MzkjBjirocPi/qTx8Q5R5cDtpfIBxdAaFaRCYHIXMKsYpLBr1g+0apH+AOpxFb
QujbZzV2cb8XL8vqgXVcDSRg4TijicI8unn2G12VXe7MdhSZFmIdlUJArm+GpiOB
2cdxrVLHsycpRTlGL3fMHvS1ctKSFLNbaXseFXkVRQb07RnpEGczXihWr3QslORN
AFH/4YmY40d7JgfFXynPIBogl3klLrilM4W7X0h++azHBkl1io3Bm+nBd4Cc1L80
9z12RKWsLjYmgSPzQBOnQwtiijOLMD/mNJnaz8OyE/NJXKr7sqwyPDOmJ6X5RCHT
9lUNaBTnreCQc/HtYFrvdHcT/d0VLv/uOhPtdqU1R0USVM3FzX3OJT3CplaW4N9X
+aW9Gl/g0/ZGUxE+EkCWddMDGZn3Kc8sWVboq2fvsN4Eeadlv3APfSxgmeUir+dU
KjVafyoKV2msQIrHqjOOy5mmhqF/E8uAemvOmFIbLLo3LDCe341Q/g7Ieo3yy+Kf
eQ115w+UoKv2Pmo/fpfN634s00cxRl8RUrrrRyZ/bdSLclefCbHurVgrtiTakoMU
F6F0UM/LJFOohHPzk+GCCl+r8uGr5kl3wSPxszV3JyBob7UJpjt80uaeBG6HXRre
LR88OiuF8kVMpDIc8JXaWK0OYGOm7UQ8P4wtAmRK2D28U9T0eTnIGjNdcWJTM6VJ
lSomQnGjT4kkkK6C5C8rU11Pru94dCfYYGU7ZOSkGsHO8u/JBhBVJWLkkK3501cg
auj6uudfxryvXSg7aoCUZkT/97ANe+q52YhiRU1hi5rEEm3K+GojXLIzo3NOk/Bm
rtdSADEThMhxV3vQ2yMbWP85psu/o+QFEteibIjhLg5XJgxUC4f9RDTqo1xejkNa
iyQWj4tH0MafgvOR/OsJzJ421SnFDHVxeNYTWg9P7FXmgcHQ4nng/L3TDHCWNXSY
qKzXQQw1tWH2189BNJUpI16QFR4C4T+9xJWWeUOiodDEzrJvliXVpOC2ln+1VvMv
yV0jjvuQmKOh76i24nI33V8ErD0YECJDg9JfQTAArVYvpbkZk633CiwKCpoHpyMJ
HBU7bg/PLx2KggYHgZeYsQab+5JwPmuaxaZsqUlIAx5+o2gWv8OgpmTsZ/7aUy9K
y0v5sQ9UJtU9rNKwY7ndjr31aZtnaVED9NJaGovUdQji7lE9dyceMw4rUCp7+uI7
PHhvX5qncW6OCjSw5t9JSMEU+CczD+bLFT3xCQ/6te1KCx4M9kbPePAGsCtyRw6h
6T8i9+CsmmjUuIFfi5yVmXj1aEnEWrJutUY+gxiWQb+BJepggmaSOHTQWQ7t21dD
Q499gLg1h8YCWZkrOtDG+Xh7JWhbQvO9poOoCK6itM7pV8Pyw8YU9n1gpK6j96oS
f1XDtidAP3Sq0vgH/5rPeWxI6/Mn11OQa5n0IcXCqXXllPxRRzXfkC7KKRlKo5FB
dwghTvIcUmZ895tUTdZPvsCju6pcTahQnUoTEh5Rv+adeyrGPMpmVVvh+K1zSFci
D6dooo1uPAhBkQrqH+608vMGu7HtjgaSYFe3EKyeJFnx3hgtp3mJJnoS2vBvMcys
D5vSHQIZZjLYKzq8s9sCiZOBzgVlTk7GPUOVC3Dg/HOPRgM0pNwK80H1Vn1ka50N
aAIzgoML99MGON1/OI6eeBCbJJ0RhrsogxuLjro6IC9akzTsGMbMa8lHwnsAkdV0
3D1Vzyc/HlURDHJPAkivU5+fniNQP1Ev3yGLE3t214lRDPSQDLy43yPzcsncX+RH
fROnNS8rGuoVLYyK2zm0gYfHUKPruhc9w3t4GWiVGkbpDgUTTdZAzehrh+2ji5IY
m9VNHJNFtr0QRZ/+fYCMYX6AGeF7ldNr5+ei9wgnZtiCh1FibPHgN33E7/1GBgik
Lz8LNDvlQTszVUd8TJvw8ZYO0IG/53FYaJnyK5bON3Ys7Qq+6ysRhnU0RT4ym30Q
9UIEmX8HKci5WY8ToQmHThK2R+5X9+Ki+8/OY8HSpgxRPS/MzzKhEs0YJsQe7aC9
14ABqQ99gISAZTLqPZZDF/tLYMkrngJoJE4h2eS9Q/PflOlUrr8Mft7ZolYNjat+
Bkt+PSQj4guSogYCjjZ4JZrR9t/XKlAZB/7UmAALMpW60XYrZSOWl4B0o3ojGf36
3G8rNqppSGg4w/xOQfHLfM0dK0J16qTBbIoOsRc2Rmrbolk39gj7KyBvoixVy/6X
YHAdoIjmmXoPqVM2hEmy/sIMoAGBkUp8oIvCU2C8VhjqcwJFWtFUfwbPlstvGFhj
M3S7utkqUdawBAZV+ewRgS9c5Qq1pRWUjrIXrsq21WPo2MgCo+oC7Q/tZ4QD4l9P
o6TRk2OS3Sw1WAcbzydkvFqIg6pRmHTc23H1NnEv7J95XSpn5ZL4oj2CYa5WpH+I
KxxN2ToZWoewUigSoQ0Y52Xi5PbxoJBAf8lk2UYdAQIaI6fW1Gopyl5hsR/o2z1r
XVgyRCDLYW9EhbECZf0LTG9R5LePPvccs9kgXC1VcpIzvGHcaq+aw8XPqpU0kQZp
2c4J1YXajowbHBjrlY4Tk91icYMFP+BNEIxexCNUFZYdjSGV4dKtw2idMXh2/q7r
9ccY4PhWtjU7ncC0zdGSemRqWgAI/BSWv3l1/rEfIlQiUJCTBeJR+lD+5qDvL+SL
PyDV1TnXtW9ykGDWzW1FoWEbMKOUK7UeVvAoeDmYkJg/ejs24cavqW8bsPRXSZBU
a/1iKOpfBfdTdF/hd0u6vzONbQdm5OUxffaHro8ER7WvXP7EhQvYUde1RseuE5Ur
t4m5tpXvs3OwX3wRPHFAVEDIzAn0ueACKWXUenGvj8QcRE8jfoF3z1bhHkz2POQD
7Va5gJ0s1DX/AUohxMnoGm78qq9jrLHBMPe/JTBVUNBJYSZfES/83FMjCxuj+CO/
xKoTk/PPYN3QQXNbmvZ+vEbkRzRBfetODJakYZ5aHIVyIPT5zHyGb+fkyAx23b97
XUSBtcWkEs+WCmkIDVe9nlwkqG9V6F2I7ZZAmk/0k3IcGM4yNXu5kakP4nq7aVu9
EaEQV0l80Czn23pVqIt+iy8WawVNesqj5NP/M6CIm2oH6QbPCoL+5v7Ip1+8WSUI
Rtl27Z3UN8e8NFugGNFyt/8KUnWL4GgBxRJsMIHXvM4kggNbjP4lNl4oNg/nAXyQ
3iUgRSGEwqcatVXyqdxpJOCapkXIUtgDpxO7FbqKRXargVVeyYcVTFo2+gJWS1XH
gquUT/z4BmC6UPoQfblPOkSYkPO8mcQ2gb3OsYKnIFtnV8BHlWDgl7ZtKk62DGWT
ovQZNcBFGw80vV95gHTiF071RQOC5EJFgPqNmuM9qP74BLpxRZZfaPl9S/JIK5Fj
JVnm+nvYXmWin//An1LQOhumWIFoA2Bz1RZXh2G8JqCiDIQ6TOyFGfa1h0I3Lfm4
1RsRr2Yq3OXWRitrvy2ekBubWYYrxY+NfKNTXuAgT2gm50+zLpfykt0BU3Y2Wqdt
VyVZCA0gxtq4nHrNSyAaAWBnepO3C2dT8S7o/SN/tGz0VUkX5D2s85Pv0hr/kErE
mLMN2kyoKiLsT+rSP9J/5+Ks29+56Z5kfBYI0PMhGBIFipNRtXMsAj68tq2Drpr3
B7HXwe43Qj6/PwR7W2lCS/AQCtAUOW7jF65EshDddZujfl5SenMB5LZ9+D81Gxa+
wIdvfQzcUJ4RLzPBDF5RfD1Tr1XVmJmfZUVy5j/u+IMKYLTSWARcGuKG0oV9m+gl
meCVRqMMAGRDd4uaFOiAFpvn8AHuaizEa91LH6THomwFIgXhBwd25h2OFBENdY8h
5Y6+j8HNNnxejCUsAFQ72Y9qdNxkfDkPTRyzjme5BqRm3ebHxBmFakDvxhRn7K9j
4pXpnvBHnGRgZYE4yIcMD8PhaO0IgyZHQkydMFGFd5P7XP5q6V5pvdj98+/nFp73
4NYq9YXKWVe0sox7w2PXkqTvScS5X/QKt37CRKi457RTz148WyzbsnNLXZMANug6
VMsXp4cvMC+3AdJRg2H16eGqEtQGra/eWNiw2qgDi01ocPXitk7SJTvz2z75Zw3/
6QuSDGcC2l78160Pg0yn1K81fHyuumOLll959Ssq+itm1bhbKt5811Psl2TzJQQ4
eCFaNPREuC/XpQkk5kFlvix8eVlGGezabfvWea6OI5+vTkXux/1ipX2HWKLDrNyE
m5H0w9viewnWRsynRduoaQoT83hmH1fsNmyysjKKc4FYl2uiqxzLXYuopNQd3Rfp
o52w9ONl5+0R86/sN8BQYUSIe5RullaMyJ+gcBu/VgQ6koJctv+TzQkI6gzVL0xI
iEMf+3u3/nkONS7NB9GyCersXaj7w8uazJUCWXcJeUK56HzGyDySYvuNCty5aIV8
r1aBR+JvP6Nr33UhT5YcAA9g0MY/5c/j/0K8+5WydlZSSaYdQsLnUheBC1K7868Q
WXq2cJMyhaYkSwb8ZftCfBrXaT8CgpunX98b8kTKd/ju7AAH2bAhR+pj1ET8LR5b
mgUHgLcafBFj31QgOlQrPoRS4WkKh/emuCJj4HtbqqZeE6O4wlDR9LRLkc3vB4xm
ErDm1d/PYCeIKRqhVSHt6Gd506oxziyY9SKSAcDqWvzoGtGPtZVAiTGFcQuHADoO
N31lkIawMY9At6zkUFYLIour7s/KB81qILVr6Q+2KvJjRbSK5Dbn3dhUOPDs3JQe
TMnDPN+neaffTR6W4hwKdoP/iH6pvQfRQ6j+c2xaukCceGssiCtIOsohJJzXqwvb
AM56lTLHCISWwPF05ZwQAESY8+T7o/UPOLsK0sQ8IAHSHng6f12e1teswypqitVD
XzIcQxAFVvceFDW5YzuFHRt6r4in5Lz5Gjlxk5Xf5wDQRyYRRpEqybDMnXIE9rzj
+8s/oHtPzYl4n1L4AQBce+aSHHf7ftFgxTmNVLtyu3TbBp6WLQGA0K+qvDUuDuzf
vpUEdcc14pNXheYjlj2QrzaQg7gjJ2I1lnyWUv0ZzMZKFKv1c/QD45yDi3QWdRfL
h52/GRA3aZlpLbXpm6KWioMlZvebReIPcSQXt7JxhuIUm6WbsolhS92EGrAeGWZ5
VA1JPsmhfvpKZCS6nE0ey6kajt6xrYb42HJRhiEnUcV1YwOOqYdEj7TKrFmG7ESh
hEpBFh/MeHPMf7c6GCn3dzKAO7Zq4WvqwzCRRE/5FD2wiWESNoiF4jkFMok9xVhp
V+LSxB/y1Nn5Em+YAIHP2xEQEh1e0IvgERRyNwXKpPJoulXFE8nOYujI0NKPAmVr
JBoGiFtT4mKl38sgJHFCPT7PuQ2eV9Z/rxwai2nVK/gHenfXYFxxDPnRkyYqlNAx
vJFQm/OE/PWSiZP4KPK0Gv3VZg3anifMfXxmKHeMdeSxj85RUmmqSyPuAwhyBDvg
HmLyRlToW2oPFFuAgB7Od7TL/g3UDU1fZrA+Av2IUzdDa4KrekwOq/lvZ6ml9t9v
Tj0VG562wGp4LPZnfzY9Z/5F6iXp4sGVtfiHQDiBauy/Kz+v2H8rONLSa6ZnGcwI
i/3GOu6dyP0pk5eIOmX07Tj9MeShCJ8jKuFVXbrxKXDMC37yRsJ9cQHcSaERA1eO
LTp3YVKmpufgUzPaFaWT/8VXJTpfItfTOzpcpG89mwdelASLfLDHMzBabqlhImKU
RX6wMTftLBIxaHdXHSr2uSbH0mFB8Q5hqZfZkFZSsE9xQSktO7LQ//uEYo7Th8Pl
0VyDzOynyCoaC5hCvSCBMRoK1h/geK1NYwDkx14+X31n6cNg+jap+BS90DTxhkjs
lfaOei607hHk1Drnd/KuvnEdQZ3Pmr14Brc83ip1oFsbmN/fN4WFftxKF046bTFI
Vbl9wC20NSPgyu0cGisCMzryoPE6dzlE5E05bTigQurYRy9SKMzh5Yc23ybXcoDp
JLb0RegWsnRkLMYgARs+KPtJee2y4ZoveAU+4d0izROxaCp4v8SRSF2GyQhAKzWL
1IJ7FRkOft3SoelQcZrGJS/0iqKXBk13IFJstENTLt+1QKU0UD/LyxHcXicLqCME
O06NL36WnGRyCpQZLN1aacomcxk1lYEOUQmtWhVy5OWGtOUNdhgCQFSka/dQqwQA
v93M7GASc1oyVqetDnVHGKe8xQrHgsnO9obnZr/+LgbpwJKkbu8rl5WBX0mkSQge
MO8qoKZBXxGFFHeoI/VNMc8X9f3HALykpt5+NJT4FP4lV692i7qiNupvA+TAXPNJ
18JMkMkembkaDj7VEFxqpJISiynG3TKArF9+3EgwlHj6q/XQ1nqCtPkHJtg3iKi5
97TN1d9KAIsnFFk+91QeNLVK7GNLbxnxfl6lmAuemFEVzoxk2S3UWHd+h5J0N0lI
CRMhibWNusv3hDpW8TEsPt4SZ3m3FvI5Vx7kCRb2r+8EUfcQ+Xcyp2KmvWWgH1ug
ju6Nvoj11+zWTsm+1+EnrkITtrA/ddsCneM9nT7/RyXV9qDVp5osgEfbUN3xSEYv
kvfGtwKseerciwhLwD9mgN08DLMia80BUUWl4abL3qMdgcD7IPpjqx/sjfXDpTXg
baR5mPPhQoHIiH7MXUH+y9ZMwMxok4c4ma0CWriDQzrIe4/as+/OcdqCXYiwa6OP
8k+mmC8a4HRR1XwkjlMAZLv1shmi1LwZXOnlte0v7O5jW6H+XC6WCFD1AOmJTg/P
RHFfVHm0BmegmnNgly/MRFvKoFi39ja67uCruHeYPMXWPj4uJbLYDvRr+E1q1UEM
Bce1+rbaGBnc0YuccnW7uiYJkw4lsQ353th0qPAgItK+f0OqUnjq+nhc2FrG7bd6
nIEgk4gi2D0Ss+wq4WTZRCbdNiUC0bm4ew1x5P3uBNOIDJW3ERpwBh6XXXon5vu2
AlVylq+yGKDe2e89S6wlhi9egfzoY4crtYAh+Ze5mrLgxATiMPakg5mYvMKH1NUO
pB3uX6o48nWIj0ICcAOdjZONGtJxZSTCSQdfOvhoGISPOliF/UpZf3MLWxIJlraC
vXujUZBXITBsuD/n9NJVimdxaMjUuX9HWlLIMaaCMSEc6rQogj40lXKlstASmzhe
x5Xk3DGrf1oigeZ9T0Dh/hSEhTv7EGj0ttaRgFMWCoYRNNtxEm/jrI7MVeCjCUxO
6OUcAX0y1HUdYg2Ir3btgMgVqV9lW6mJJI13H2Hm8+BChcexLtj+4yeclHpLXBi5
C+sNyfMtjWFWZJM0ea0RDQDlFUwyTYdTjiFNUNBusGZDDGnXv5xCAvIdKMtWOXCf
p7lMtlIhrfSnfWKdZD0485nZZnsiheYq03GhrOd3jfcyn359DXUlxaAjd4046KQ6
lUtxC29IMp626B2r5VB4wo5tR8hHUmFxNpDeY/GBtwsvgcERpytCcz6fkQQbwSwG
Yj0JWKJB3bHoM0H93hXxW4xBl6zmaS0x/RbCB8xDhGSE1HSJ9lvh16c7tkzxaYYz
REAl28ESgKStd74T0a9O7MRMKmLlF3EJfzB/rjADaUd4EZwknV8M2DDwKfPWDaJj
lev5f3di0sxlZ1Pb9zcVDzjIlQ4KnP0rjF8LHnQjowL+Y3lmBjgh4jbY8g55mRGf
vm9gqoEZX4uavNC3vlYIPKmp9fefsP3hd/SoAZ9F+/ZAZCvecuz/56eqnthinvss
DNNBMlHRM0SdFjWnbDhGM0dYWPXWnPtXPSayzGvonG813/JRa6kK34s70HsIqayr
SK4DW7Oi/Ev2WPOoJ9vUT+mMk8U8ih9FDTK1QvdqolP2+gF6E6nVPnBJzxj/4osF
+BexVTU9E6h1crsCoSqBuXZNIhk2HhDnUhA0l5Rqw9KB/7xr64ERSAzuYFeQNNgg
z3Wc0GfxxaHYsfyrvFBM3ydisUuxu7YKjRi0XKmaGjSQ/CAoWN32s+mH8bCmNjtk
jnEE8NAPveS5Yw9zJ35s5x9kr11B4uHOayO1VaJTPW+3T5Wdy62Htx10R+v43X/E
xHg0ca3eESpWlQxomqRg4wVEn/gs65vbkYf5ux/89o0Z5fpZXwpvDrvRKEJHdSJ/
+guWYkH5vitwhnwLBBlur3B2M9CRfpA50Sp6j1aYwiTGMcc8QpT+HxXawNb3n+Py
p7lwT/uQmIRODy59pxbAhJMLt9SbKrxKxrzSCvvGOmptP6PWvv67vaThzCFWjVWQ
xliWw95SLqsRs5OayGZ7JtvjQ5YSMlH0gGG2k3IqQgfOrr3x14NKP9SLwgHvIXIr
UJqVdTQjYcmpppmWge4Vh4+hZcjFNAYqeYNYQAcC605oFGtPgO3NJ+iycDJR2ZM2
vkH9oxFjAXF2JFTpmJoMVV5wlP2sX7FI5Xt0EtS91acfIUGdPjtSx+kqhVc0chlC
Md6xkL0a5I0zJaFs70xznvHy3FnW5nnsBg25dwFz022IvBMnFgU7jBhlepD0A+pd
42A1fxpAsAPszzX5oznQgf9g1ZIcsL8ejRrF3pDpqYaKja3fD2ddL7slRGJoZm9s
AVmKq467zCGlbQazSsod/M+Uei2QSmXKzKG779Vx6idDYzdbnd1sk/NcYEz1B51K
TQXrDnjFF4a71PNmWqX6Iqx2Ba8kxuIPSxBVrJ+QquFgGbbb7MbiVl87X7BBxacA
mj758pu1ZhJ7YOefggU+V4mDP/x+h/BE1zbhmQ5BF90kHficTf/w0GNkfeeRDo6U
oE/wceFcfX8sUVHRGKs6SgRRG2ABTIJM+8gE/cJphkCOPkiUOgQ6llpri3ki7uEE
72dTkR6FR3WdAWu0N1c3h7JHEp61qNTfJzSmTF7WpaXFiRRecGh4K8O+JVAzLVqg
Es3fCSo6K61OaZ6LRrnRR5HxiX4hfLvFr7REVhBVJHaaSAEWKYd0M1Zm0f+Spdlg
lcBF6c6ByQizgmiimCI4GYdUZzHvent+Kkm46JeAwa8Hv8COQl+QGLgO2lGm6i6U
4BSAEXnoiQ/6yh7qAwsn7nWRe2f5UFwW9jc6BKU4xZZ0TPStldNuaB2LdEnLhcEj
6Jplhpsg3jQnhEmIBahhzh7aAB+9Mhh4HS5dr94s3mLCybhOiwU3aCZeH4gBqw5B
uDBf5VVVLxkdyUynPIQDyeojppA9MtkKG0LOJ7h6LyRZ5PdelOTCCZ+FHnatfy9q
CyJ1IArhmtBst4Yx91KJBbDbBqM+BWi40rT8dcOK2Gk2iZxrq4S5dx9eruTOryLp
84GdGHURZkYLi4VQ8LUGVirLrc5W2YWgJ+TOtkbVX+FEclj4t7z/FngJc+hIlh/6
Ur2LtICWSK3UAn+E42AxgTu121Mh5ioWcMdgaTqPDIAo/cp8ZY1hs2QQkUggmX2R
mykko4nanva35kCrLlIrzx3mlzjOSacBBAF0B1z5F/SScKhUevx8k2M7JlH5YwoJ
OV95tmZlAWiVwnRoaG9ZA5S1SkEE2q1sYkiUUHuiXINrM/IvO7oWy7AZp+OXLKiy
jwGDsdr3sxu6l/UGGLKteHDuWZjqRAG5QNwp9wuJqYzSuvyjt+AhY5FxuqT/EycG
+LUChZLqrwiGcVSGegWruPyxcrXftPUpBGS1SHQvnAil8DyJCuA9z3q3gBQuU88a
DjlBgqqEr9AutBUGj5iOz9BajGGRuKuPWBOtfs3lM/eKQCThR/Tkrs5qyR2owyKj
LPMKvxMErDHRRcH6+ykUytijEfclBJHX1DxLBff7sLiHxfWCvGfoo0vGJWvZOsqF
DcMr0MQ9aXhYFNIa8cm//fphtYyDoNJb95t9kLewOTUK8Rk91P74JclkSBzAysNP
W8Z92LsOB+hDdQYIsAHxNoYKf+c1pLEsa9J9Z2sjRaiwwVupDeyq5V05wnvTRoso
O17AQd0TwAYAaoAMBJ6z2vXLPojQ3Bm4oTbcYKt5CYHzldoalbZGZFb3WIBK4mSw
bzd8Uzsy8n45i1lpiTB+AWxG/ugEfsUXlgeE8OOnIuXGc5WMrSC7zZ/arPaG2LXa
/Ha6oqTXCuHA8AJgO2kPSOeNg8BLlFVe7QjXb+MAuPdBNDO6XMwHc5plggfDJV8e
N+qJSFBFvnIlIaXAQwGSQBb2ZEBEetngpwsAngN7BXR30VHORyCwTZZfJbb77xa1
yEakU2HA5yEe2CgzT0Y8rdOEcbSmK5YzryUGg9AzRQLijPmMp+NEaN02/1zRXY32
wC8SBdv3Bsvl4YtVYIq6VXAUQDkWvMrpVoHf+lM0XpKuROOU4c5H8qhJySgtJlB/
ncqVyqkkEXDe8KlI7n8Ax/V9K0Z1bVAYAF52n/zBrf4trzeivPdoRR6O4ud5BOwn
0mAJKYFDBfTsIznlPYdKfsXxWF1Umvw7Le9D3KouH9rlyzOWFT7WjmRvuV6PcClv
2/jm47jNhhCvGqB71omx9+vkc3K5aVxUNT0YnnBc0scWXTr492fjrGPynzCm7fIU
j4UpetEDSyU4Qp2HlHUEI5Psk9IiDuuuM7EAxl5EAvp+CJFoF6uum1V4JrXoKCMZ
1T4f6Yy/xyzHRjkGxi4kPev9XYjNJK6NSa0sZ8A8xaFUPTFV8ZejqAXbxvwTTbr7
Dv3QPbB/6Jegdi68K8cnDuUXJiqQ+/R1NHsOlFiMfi0cq6rFIAa8ImbOr+yKOF3U
OdJGboii+f3kwgiMlMmlaiRSzdzzNpRGvnPF76a+XDhe/LVZtb2udUGSzOFormsO
0hThY9D5tLskrz9FqXCoC/xJ+Oy8oPlQYVzyOJMscfmWRBI/3+7goLanQ/XsQuAW
FgjMzhfGpCZqPCuG28prPJ1StwhxBdK6qxMcR4NVRE20DuFoV1XAhJFuRmNEyvsX
sfNkLFI4LtB2p0hztNu6Ugs1InZXeHI+EiuSLqqVlA/QqDVsUq9k46a9y/HE2ch8
E8sFH8BsjqOgQFwu//KpYcJl0F0rJXdeMqsGDxcfUs431tM5RNXEkd615SG2cxoq
CBi08hPu3qcgB5UjxLE3pJN/95hwwoFElkz67jFGeuTu+JzbJlWnwU1EqxA7gD19
s3WA2m0F1nwGfm35GtzTCb3qesuqdsBp4TiiTLXtXwhNfV34dQfIiIPpSNtkivTa
vwP9aLy/tChBdPi4Jfan3lj/uBvrjywEFTDgelVq9d/qi/m0e9jlwkyb3u90dWHv
DfqWD3m4B4TaC+CL+2kVx/RuYalzzUeNcVtrzw95bZSCd2CtnhOeOWC9OUrPXwQ0
6KqbnwiV8VdDsbPGp8xemnfCe5XGAzMgjxi8M2TVChT6QUnuziz1BYmqFt5aJSlR
z5+5S455+FWoyVnbMJh+U9nwh9IA/bP8gg99q4UIjwLiSp9I/tBiU9facP9a8z2L
5h6n4/LH2F2o2dJD0wX3h22xo/rZ5IgFX3DOWQOdH5I0ziUP3Rd5VgTZ/fcWNBM7
vdAPpB8J+QMpSw+YyG7xvO9zd7hGg7eLug69O2c9WBCqOnCSXWdTwAWdmL7OoUbX
enmrwLgDA2oHnkKUQoO/6XOKXZco7ftDcBRQXla3Z5qEWDJy0Ih35khpbIbInb7W
nnZ1sP7txUz7Wk5KD4yYm9MGyBGU6KaynedVq2O/P5nudONMh32VsNGoJT4LZyb7
xEuuSH5x5BWlO5G9DKJ51wT7Jbrx78v6vNYcm5YAaty83cq+2SvVH1r+cRkxEU4f
+kRs6isMYAxP0CBJD2mON6/ivXrXoUUy3k6hFJ9golkDha2hEv5FRYZ5zHgiVVIj
8HmDMmfeO5yRwqHuSK3F/bPt/WgtlQWkAf20YckNQPvWKnjSD58JjBHfsTIN+KDS
JeLX2Xf4H+7WTNt6IWfOTEpmoPkfqCpYvIPcwePmPWPhTXAOB1aHT41cmnywq5NS
FwvE+yy8cj6qiktRFSCccjfOulzg/NFS1ALTUWoCng0Cy+rB1r6vKzJaKfszA6Iw
N3mkD40BFt4zWt/ZuWkbX+Eyl4+FSAAwNTaycYHbGKoS98dN6NBvIJ4bzs0VYzYY
bcFbK92eEBVhnSvjm1f57re0Xdw+3PFgMi2fMoWtwSMXHNpKkjB6I2R/83tNkXTz
0bgLNKC0h6vQ6tpCj4WcgWQWwy4I3TbZqksU0E+Gjk7+zMK6DKLqzydq4k0fFsIL
RmGphn+F2TfaufHsC1vDI4niU+Xj5P751OHxyl9CfBSOhJya7NgqfRwrEFx1RSrm
Tz8F0zZ07P74QGoXC8+OZv1iWNsbjYsaD4cE6ePUU3Lbo2VqNR//bqCerpWrSDxD
Lts0LzyhO0e8kvQQp3JWQhmwt4UNVF5KMgPLSP9UuYXUz5vJ4ND7zVYB2YdUDpfW
tpUv5LH55FbDYzNqSWRKqrtRnDzi5tKJOTnAtdbeVl4OMn1C1kHOvGHgIaRLZO7K
kKpsLi2m0ArOIklC0lef26zIxroP2UinkcVa9o50u6skqLFMQxPvZXn8a1CtBm+7
F1QLNdaVDVgSYanadtwfTsfXRGI4WBl+9DvXjU47SHKo/lzVIGpJBDDPFCKdpJqv
h3KH3zAMmxkcCwnv3lv1dGPOjipP5lUKJEhH+b6Z+Glj4g86VvAQFPkkvoQRC1lK
lsS2ofM2wnFJ4eVFwtK91UZCCnTD1sm8Kb/0d2SuSy1KGhdd/YuZeWnpG2oAbhFW
WQ0uFzzYMtATD9hkQsGIpLM4m+sESnbF55WycO7y/mkdgsHtQfMk2A0abcsuz97v
nFO7oWzzNdNLriwIbPUPRhbveEo18x6lrHkhsg7laxKi4gy4qjpu8PeLCQS3PI+W
ULzoeWq6q8MhjiaM0IKKVT1bRBFGhKEFejBclqsqGQEkGTl3hPuw9Fol/60gkjCN
RzEqrhGBszw/BEVAEUot00/icVX5zgUCsnPQ9Rk+YZkUNB1VKIEfyscRe3dwFU+D
22Mto9S/yyQrsi1kgHAgHL61OIatlVrb0f3gJfHdFCmTNnMbcPuwxYZMC7gMXS4k
ElJSDKsXQkc8KrXVVAX0lxWUzz2G7RIDimJZz8GKi1+a9jsU+QQ63+R9+6aKNZZA
vtEh54mvfOM57yRdwT1aY3jAP7MJNw2E43nVOiC6Oa47Cjpb4iH5Jgash+8IwDyj
qLuzMBuHrtMQFji/Nu/lvQouGUZg1/HrJ5CyEX4HoicYeIoHePJ7q6z8JVkarCPu
x4YuHdRNAY0bdS52m2d6qjnGicb83R+m4OmT86rBJjXwDbnjB13oTdbLvdnRcqER
jHxYiDI++F6h28cVsxj3OBqmtjyTbf91N6eZLe3FSnPfqjsEgrkmaCDMP+vACAc6
JwnXcqYNyBkyJQ1byooB/P6AHjszSbvacWkKp6MQE5AsvGSNuxkGmrH8lwnL/5gT
35hhyD5LN7yWEi+KBI9fptpiu+ZuhDtdCMOkYc/oYYZelxsAV0q/8jKVYLM3XPHQ
WTjY3jtoLcvS3WgYDPbJ34Z83GYf/zfv1Rf2HECQZmnRF2jY2XbFPhBEGhgwM3UB
7k46RsuDi6DbQGetHlbCuPYcgnpdgKgLF3aWg5EUEduwZEinCGByroW+fkQ77+t3
afjXgELEqzijlOrFh8ENKqeWeNhgrEjUJJ7TVdIT8l0VhuWYnEpjWTk5UPVRei/F
woeabFgfkaX6xkebCwxTgE4A9tjgx0oiNTXS9k7g4nInYGPoDq+zo9Afcg7cTHPe
Va1+d5SOUXBKuTcqJ4PXaAoZ8DI7zJ5gQMxun9APEtC35sEeQe4P7QoLASE4gjYf
ygBWM5YipXlTV8O7ujBgNPY63isSULzsxhL5Mc8Skvomg9dSbRL3uEbrE6m7EGvs
mG/UZtCNhVcHhHgZ9wSc5NT8JRmGeQGUrhgVieL8oarpqhh58n/fzHTjwepaXQX5
y9shwtigckX97EABsEBGvfQOdLflJoAvlXN5cXYmvdF8mz7Q4Klx+fF7WtudnpZT
/tUJqLYX8VN4OswJ8XwvTmjSPaUYiH1pl3YcZzFzfgKvfe4SG9s2rX2Qw8PSVqF3
WmZogxh4mqDl+F+c73+0hJLzmoiDKObjlkaUn5QmJm32PkYiv74rvzd1fs8+dJhP
eTAiuDkt3x/i4i/f7Tk/z1Cz1JP7WFmYTsbdxL8xAulO7oYJ47ZJHwLBUP8UlAMv
eQPgeDiTv2FGDL66pN2okcH6An3TL5T4Xx/Puiwq0zglFpfK/31+ZdRSrEQs02IA
x6opDM1NLw9I9Yvzg/m88/VflERd5QlVp+qYc4GJfRyutaTcKVVgXI9+n3Z5DumO
f6d3575yIOtIpnZjBFsYTF5VwVfPZ6lyM7D1dJOgq9QlIfAJXgF7uFkyVZE5pCFJ
lZy4w0eHA8XuCX4i5Y+q3TfDXQQpRTXNnM5zb9Y1lH8bNCe4HBcfnziL9m+2uOp9
zm16kgoHqnN8SKNhjAHbTm8kkmOvNwmHUPaUzI9TgRv3gwSgnkA5jND0VxncMs/b
mWIFfJxC9H2TiZtCyaC2zkABM3ENNVmuRKztKZ5cWc5BXd643ksCRZVUBK4VOrwl
AySYzN8I2QWfBtQdnGKnk8jqEQd19MtLKIIhJq+MwJCF6HRb6kQkoUVF9DpaRC6X
bLfo8l37QGH7pSOm3XWNNvB6aXtzEC3Kb2MMboNUzTpzTMtvEvkKG6tuKnOczjZV
BVQ0Z363fukcIT/CUHeZGpModDumOzLcrz2787U4q8xrpKsWtBFWmUYQB2nGDqz/
0oRQXXL47YH84KW6jltaotdI840twc+qcOrrYxSfaCkn4B/eiWjXFs8cKlkSqgcA
6kbMZFFvB0K4Z171JIT2858J8Ff82K2IWz6uEp7jsUZDWO2Da+jpuLHG8DB4a0Fz
uiuODs/VxtsrpPK8bw1tcbsQImz5kvTAfN44XgXOcD0KIgQ1J3gvxOOj/Kp0PkHV
u4WH+uSshxRWwqMA8ZTH4TskNilT5b07wmXzZ65iGdALEk0Xn90RB1R2FNpXWO7J
UpS+sT3C7Pl8KV9v8OA4Z/oxkjalZsIoZliZ+kveCx2VFMeBM9EpVDWCbx6wcURJ
3RBhtW9ZhzGaHh3E9Bw6FR/gYZiiq/Z4dUjsQuTiKqFcnmYhR/MjoODY7X1oF3Ii
qQ417eXP5zLcWpVy0Xn6r4q1JCxW7TMAYwbY9xkSMaZ/vWPhGjUPoZAYAElXCo/P
EX6oZ5aK6DbyyYuFPJwrPq7SoDYtEROINwMBO+gBry3dh13ldd1ekGP/i6XrafA5
EfBo6OAdCCXfuaGItSnWShqFYfy+laKPkQX1bToudGbQXPUQmmMJr8/WGmpqyDuB
TytE4YdQ6NM6iCnA127PHQM27oan8O9ffayHOtvz0HiJKLvlqCY4paer8LfsmCQH
Dc9brwJ/lKbGmRUNKZpa2F8rj/WcCnyLqTYY/HGbVfHhWvj/oOAbkW+u1DRf/WIv
+k1WeFQ7QAt9soyVKOmkqqxgJZBEzx2VHw5HH9bve5IwDW6VU/02ZLoykHKtoIkz
jBOmukl5EEpIPZnyPRvRCvd0MfgDQ8TGxmczF38jgFqdgipbF0IqPLKrHH7W9kp0
UVEc/QETO/YuD5xGLMM33+i0WGuB3Q+da8/Azkv4xKgWvbeRKDdyK3jYURP62Rj2
/BwO54o8G8Z+8LJdra6xJaV1xEBI/+3MYsVVzbdpc52cX0hwfXf+PBpDDnu7Kmj9
gcC6gGVaPFfNyLYTgv9NVoRf8k5TC75anlga7aB1BsmWf7WRbc80whh/osYGOzv8
DLxwzTUNy/yaYZWpAkBed0kYofNMjyQrlp4j07DjueJe+CDYifDrY2/f8HbioeCh
/2w0Wpnfvn4vVYMbNnLfXLuQQZDKf6lWbSGksTfbXPp/1jkIugwWCP+IRVROTMro
rVT38QhUy4s3VjBr4AhRCu7sNZ2bOZnlHgaDSgWoQqFmfV4jlTP34/SoJlTnD8CJ
PUwPe2LYmmARVx0LGinGUFq3PDJ8Lyp/+haypo2g5PFIUAauGUMSvvbJOGVlseVV
6Q4skuGtgtQsoo+o01Kw+VLNdjokrLOxLeQDlBFrKZT+fjtgNWonxP5ZoFApwfVt
TOvEeZ0dvmrpKetalTHH0SGNdME8NEb/PLuJry1PE74Nv1hv62bcSCGkqzsFw3Fd
C8jWiEFspE5oNSzK2pFgltmBC3C22yufN1MIxGU/lRIexMCji7yxVvNS+FtP6jlO
/uPR4lRWOVn0hbBA1ysYfG8DEOfeB6wU9ji/Qz+S6gp6CTWExxqqkkAnKDmcFTfc
Th55nQq4qB5HGFMFPHkMEs/OkjpFDH8/bGsLs9vMoyK/zuedir3K6+a4rmvpC/Vh
6Yss1wEh4CCFF/T4hGjzPTUYHIHjb7WHF5QvuPIAOW5xEekbBrAKzPSo+LQRXOz7
7Os/LO6Z3WIgfD6xvMfFrk3HUDeuMxRiIzpiUAaPiI8YCHW3tLKmPuidFkxtQ6vM
40p1ve5ZkWufZSMoKRnQmutChgIHE2iIK/7wU4ldud//ofoN8oAxszDjbAym153C
EVYi8NZ9Zbn/2yn2PgAWNldHd2FpibcDSwtxCuXHCNyIitkZgU9aYhJnaf15czK+
ychtjNhPqP2bfKjxv8p8/z+nIlxS2GGdQDHbsCbnLFRQ4ws/gW9WXofxLSn3ubJh
AkStnSHR65Wutyd94ifMg6aNJSt8jn+/V9ff+LYwDegiKveQgvgiT892Zm1JF5WZ
73RBfR3zONFCL9PEBAY3otMh3tcZQT71CwYAlA+kyO8TZ/EmX65Tmg/matE8c6xZ
tmjjS6DWg8b1QwHp2wn9vqyMP3viWHLt17/XBmERstXjYmx6VE0BwwsecZ+QAoFA
3ZzB+0DaxNMAgQkMJq/irTfdxkMcW7R369tN8qeWiE8U9LZNWOWR7vRBNZPLAklx
gfP3K249A8w3Ta+qZ2M4niTCfNRRms/jiEkcJHqyGLfw+8UeEUY2b/KMt0khOB/s
MBK9018AE1ojx0mTxRH+ta56zyE42VQGsBp1oGTOpL67CDvWsCvSyZRoY/qBjC59
anZzO3z44IG/EoGo+evBk46S4ixibjRO93Fn5nUIoB7E5fKirb8tpTgA6Iy66J+J
9h8lr3LNuZh1+cCVUHzcz4JgB+0ZN4FDdzEBZ3PIqc79bmADFaI+aMnwTUUKpuNJ
ND6bVPXSE+4JBNWC36wfwErk6ui3ZbRMNEcHN4W3OMIP3jc/yQHOLAOHzyMbK2xu
SbT9/WKQptEDCuCcc/xYA6DAT19Bcb2KrVFjbxpjegwqyB93qMzlCLVx6o/EzOnZ
bhns6GUlylRAELcnSQrd7i0PD3tuFlAj30zMZW+O+0lL6Gi7V73o1TyKt3KqpTne
/oBr/ClMypX+SY1kfxvyDfwy1j2Ql+ck/Nzi3LQBzHzvKtkq1jZ6pTg0hJG19pDV
mr3iTXYXoI9ZXy7xRt0tTqL+H0GgdGMRkYueqVdKRSnNJYSuXeyf9vPD1z5+uTXR
AZGEupGt4hWuF+RxpgbBjsQhkM/PR/kM3j92txhP19LT/i8CJeG68B0JlLsRpZ1o
m0Qkh/DRq/YFsj46aFw4vua9ybTujUbU+2hwYp0qppQz3B/Yu/QIP803OCBvKa4B
GiumpceQ/APAnrP5nUIpypcJcNv61Lf1X8Ir9KGa5FQg40swhd8w33RcrDPVxrHm
0htZwWVvxB+OJdY/DxpzTKH+1JeREkBR4/fjurWu+NGIzWSrj8zvRqNLpp4SFf47
qtIJvHKhY3Ydp/E5G+mJePIT3lE55MoRFDr6QKJAk4lezG/xvENEOV1pQ6i6r133
QAA2pof/XO3nrqUKEd0pXwCTzQlopniuGpFdPJi7PV1EfcOpawUIt2CxtBwBo5aC
UVjkBPOy+XUT828GR5FkHfnbUwlVfO5QWtOt0Mi+HAGQuqdcxL8eDDnMdOWRv07D
YX5e3baAmqC89pGFVY4spdeHK0JArlz6WQa1a85y4ovZPOEtFOyCJPMW+VgK1WJZ
+Bv4Irg51tRZ3MUYU0SKcWdqCCyCdfz+KuQ8amm/72sfgbpIQ8hjGR1n2/t2ukMw
ZPGp2V/lhbBqEu47Lmflw8GwRQli20+e5bxsUskx/6WlnDn9UqCxOow5dykFhr/S
PeXIhlUpSvEd7/H0gy+7zO9I5Cqx+iuvno7zzAkuVEdllRBbzLY5h5HtjLN+R07j
obzW/gkzKEi9aSWCb3SgmQqk/FnIqEYIQjF35meNwGiZIBY+tWm+HbbX1U//cjdP
iWJ1B6a8rj0fbNN52AHfmXup06aRauen79trJ7Z6gGjmFsZkFIfl7DAZHebq7M8x
YglGeJwcH8AjPiEJ+V8Dn9ChcVrAprkpBLy79LDryHslG9Cr+mU9vhkvPlAGbRAz
qRp6iVNemh+nKW+HcVEgU0XMNfuNXx1Wj0evueDvVpt4le5KfOgocIbOIJ/PMWyR
3FJqEBbOSWxm/zrKNjTt4mWD/D/QjK+6exWmBYOgeikxv5v03Yis3Q5aSJVj+1i/
K8mFCwX4aMTs2DKQZ1uAt2dsMc75DD02TqCFRLxSGbeUUCxVpDs4ZrKAQuXY/sA6
qYbJXxr/H9FGZvhJ3FHOsqudYzmkkuer5pDgm0KISMzYW5C/uzfUpPXlfQCQWQHR
Mznv+5EauSYrDIxZPDSzd5n6xwAR8uT5572/YqLqGcqHUDvDPTAPN/lMJPr2c7z0
l3OyLbky0ZuHAuHT9ZVA3wjWUyzyv7y1AsExA20ILqy0kYG3saXcRx/b+NZeDFcq
8h9mMkyBR/+u9knXUIbqgjhReCPAjBloI1u1scCeLGBPMQpDWKun6u5mJ9LaT1Au
E7q2peLX7D9ZgxAN2It8MTdybT1Q+rfR14qsOgH6LvJrDULIO3Ol6y3Q+bTpb8ZE
Gy/dWOa8+GsELGR3SgevKb6RgCqI04zW2bTZ11tDmY0A0Hs6LZmktsPQGRHpA47c
I6UnwFgaySll/8ckbZUyvrWY4Q01NHAfKbNrqzMBQ8bAGZ01nSzcRNdlfuYtrTx0
nDgYxBIF6k97U1BldDdggB2qe0KxLjA2kBEKVlQSAYEMD9ebyRQQFfyc6smlwBmj
DaDV8SYHrxQAL5F9yFKyZhAj2A+KIIa8z2NAaLVQXXtBuOG1LcrwXfhoAyQNgSNG
z1SpzgIeP+yOpO1DpH1DE8e3kxIJwIuGNRr8LvrCH5SKJWxsQuhoCE6S/qM2ZpmI
St7/bTteQeZ1V4liftwIJYOEjVoyS0JOj+SmRlzU9VfKaV5SBETM3EtjtO4MZ08o
fpUg038o1WY5gFa+sG51EHWcpvl8ddA/VhDfh0Emr3PBiedXmLaS6Mv5G/uqM/BJ
uFLbQvPmZiRFIIjKKwRrCbTH/q7gOoFzkqCzrAzGzfitYdwnKqZTsCn6hLKZkQaT
hC1YRdheZ+DcmhvAS12giAnwxu4Hbx05XUaSgFLwyVfX5VUkUIjrVRqZmAcp6ft1
2hciZEK/QXYsG/XozrSmOCj1TMT5iAxloTNHV0C6qmwS2Zo2AIhRY+zfQN1kbTcF
7p3qId9SeZZ6Yz4nF0+LyF3A7GiEYEFg/bl+XmuyAyDBFaE+prRayPVBfaxeeYBB
9/8cx4Po/JSjB3an9efQZTQLMLPbW+pyfCJi+C7Y+1CRh/G3EevGYOb61JEfgsSd
NZqFdJWSBU4dAL1ljAuUDFDSo7MBQLHsihzvoZxdd22vhA2UKxHtv9z1HzFWkoK6
qN++2CCt8v3c0U4F4zguDRUZqSSBmOEILSsMubl6lcfkQopBRsIjjNUqBemBiN5W
3JhUPcHmd9SiDyqViEoHhejr9cz3hXouDoWr9MHESvnk1cChtcOoJm9mjP6GeSLp
Un4hZwYaA8rFOOE2gkiOLIx56PpL6/5S99eok0heAZQsNwd88aLcC4681O5pU/Qp
WFoVP6t7PPHfKguFJlslOIYicLnkIAu4RHcm/ZLGLNFO9CLFD9pzdmKinvoueqGm
gNW+qOd5fqp0JF4gmL5xxj8i8dhsj94f5nfwGiYlipJQtykt/pEDszGAN2iND0SB
Tao9aUU9FkFjNHOFFzGW/t4a4FFLn11hWpUQvyPfgkFSMLqnG35zgVaEtA1eS7Kc
kuL4YRTOja5HRP9NYn9qLMYWYJEfznSVjawISTDp4hdcOv7KdqCGErg+VwyUof03
69hBJn6YZmKApBNNs0tc2Bf6w6SgOpyXi2t7nIhrnKDk6ZBLd6jYmZOeaV61Isgg
PgAc7Da2jJouLIRRR6uOi96jI/f7WcBDdOG27iYFwlXtBjxz1ORWyoBH8fJNHgQp
aYuYqv//k6MPEPS0NLU7zDyYvZo7mv0z/Vv4cuam0lXAQfPxIpxJsrxphQ/N5hCL
UPOgPhSQz2NnJfEJblg0YRrgy8kCWkvA9o3Kq4XSsjZ6eAZVYzmrDObR9za80Kx4
j2fB+rCfSQFsxBWZfiO2hXYpVuHu5bJ+XM1pDJlfRAMz7MXA/s0FTDcu9h6Kd+Hg
RbritK1a+yD71SuTvrtpTMixIr55U8odJALlJjw6JfpepwOzzPDuyekJCsBtlMcN
UfRK7L4cYlFGBF75lC/k8QzBU34XQEIPvWuEpXh9/V+QwMIb1BhEq9Lg1caH/mUQ
jHTttB0plT0rrENwHLO4WAz7aXqEyK6J42eUv5tgqXgfCizGt2p6qJVx4QhQTHE/
ezKill93zCOthRkU7VNT8juHvJcPT8xmclnSUbdUf4cfyCOj0YToN1S0OTFnShVs
CkH9/BzrW1SAM2wekBTQITDcgq8iLQaN2y0aak6EmYR1eQ0brT2TKzQ6NxwiacLg
URip8xZCRSAhOSTo+052/xW+uYW5+NUvzMsJjLgWxXTihvuBMSkpbWGThGxjri/9
+GLvEKrcg0pgXJ1HbGO4DEq6Uw3ko2QezxmTDhs1veA/Q0cYKb1LnJsswd0beCL6
bBPA/Ao4KbymsgVv8pQi5zQS0T5nRJbIKmC1293P6AiKCrZNZT+CkEvm1/TaXXnM
5xk3d12AuXuAhPWP/Ti1PQtEAtXvXFI9MMYZWQ93sFVlhrmhwI92hmcaJS+o753W
7dJOMIFA6iZREMLWBFUwVW/sAiqiLP2ZNNUiBbWsumHIJweyuaiPWb+jnEm5DeLV
aJe1+DEZ6+Fb7DcPrdla7ZAe1aWHL+tG3wdUvVg3fXAgtBCL48XM0m+zA7L0zhTg
POyEiZqIRbCCiBT8I5O1r4w7zpmIvu+jFHY+NZ/OW87pgAKBFlh9EqBw/3UZ+QC1
ZrsDIhWtOynf+t7wGS3NhMYXndDoi0h71OiNHD6uQXY375qz//YkRLvpSS6vZ23p
2ubZHAuZuwGRYQfTwCPyhlJSTsyHtMJu1qh88vNngE/fkwDRxm2Sf2GTwmxEGGpt
2P9BY25wUZFcvnCJtYIhJxo4eeVnF8hxHcp9tsZ4D5EmUYzVCxgMMArk1tGmzbnw
ynbF/lEc0kqY/eWOS8MsZCTw5X6uRCu2rphlTHJzEjvvEM4eVksqLr/mtwvh3ibW
tUA6atuW+l4VI2onwWwr1iTXjJQ4pD12ybd5HNNxQLuBaExwu6fbAMmitWteK7f3
Omy6XtcDm2OWjkDfZYjQU9Ae97TX1IGROW6cIvMhGtHyB6wM0PawVdTXzI/+H+3y
CqPI4QhXv5pDMDlyYTS3HAY6DdKtY7AVFF0AdRfctlf5KNbPdjWcjNd9hBBC9In8
EJLojTTLCZPMMN8INMc182M8ud6fFDSr2gRPvTZNyEFA3ofNxw7ztatE8r6Qc5J1
JP3C16XfWHU6HGGItVKPJJ0i1VkDG56oRvWFKDZ8MmOKnSExhjGK/zrHFZFKWTVi
LCKNdjtYbaDIgcSvHDaqEqdGcsHom/rp3zMceeketoWWk0t2CocH7gl4k/CVsKTC
Mzw8KByzG/gS6g4/X+NKkWBSb90g2bWP3gRWslQ9tyspRuK7UT5FKe1dSVPspSgN
PpKpR+7ubHXgGyFXmWlxNbr6q8p60VxgurTClrewA/QoGakm9eGNK4fiibNq4QJj
5v+bthzqgUjTCYHjYkEcR7q08KcTz0cDLJSAYnkuoDmqIH/X8H7jMDKppZBnzJIU
4fpoGQzQy7SKE9ERSxuQN2AXS7adx0KjVXI+4goVXdG6rBndvynpvWTvyG9lAiMb
YzTCYPccmJGCVpyjGGLjhqlng7yDVjRCkG5aY1lWvlazRHii0T4FrOjiinvVXV7i
bzTwSbtNMRvfjDFEJ0JOTMNuSohJYJ3QS0v7HFYX6HxvWJ5K9djJkKKxbfb6Skbg
rAp0mv5utj2MngkzVfstfLLQG/yD1140ZF9C+20eBu41d6AnoRItTw1LGoZ0xor3
Hfn20DSoE3pjf8e1DQOrRTG77sZFFjqtZIy88DIZSPkkPFh5MsNaVHo9cBH7jdOT
ba9b80oKyKb+FtIdCPEmqbGKbAX/jU8ll5Zu6VcQHi2TSYUQBl42etr/r80m3BZu
s1r8gMg3v4fGMJ2HizZx/NNKaY/AkPMFm/drF6QSp3Oeg9ZKlOOTxZO6fBhxcV4H
NpKp+e/+1CHhZSbpbYYeS1LIv7niCebqsxTQ/DeNQziWUDPfHzdLl0gTOdmVu+gU
R4uHkl2H77nlfM5G8Os+Q6QS6cnlNRXLYb+vJp45ymUWOAmtdWwdY93MgXc6w0yF
/SGkijaikROV0TIrdtxAK9Hlybaqngu1TPZ4BAVRya6P7EYctUh04pDhny4LHB7P
tRJu11NsMvAFVlxIx3doJMA/Swpb0VLHvQThDqRQfmDyu8+RN43NJykQqIpZHQqC
EH9Eg55ri5JTbRy4wFc9YKie6q8MjMjxu6yMqQ5z1q4qx/lPEDsgVa1GJJcOQH1f
oluYqa7uEZJzHnZ7qI96s5IEHaCqpCddO0ECUqT9dpSakVURbi2Zp5PPh7RrRw/3
o66ecU3wHMdEHgL82SR2lBGdQ7XO0lP9AHcP0lLc+AAKFctHo5NkuIZNpzahsF/k
WUuIHiNLz2YreHBUVycvD1HACjM6A9SzKopWAoswKUyTPl67MG4/AXVGAORtSyd8
a5o6JNEo6Zrpu5dou1IV7awvYp4aIa8xUeC0toaZrIHcou2SFyyQtu0IRC2+Pets
p+r3LJbraxF8abGPe/nd3h0Dqwa9DCIBaIrDv38bS3zxX+ypOvDxQwS0xOsjubDm
YcXnlm0mJ+sYcM8bbJFBwg5So5PZbu6Bnwbv4NbP8IXXHqbh0nBCWHjmnikKibj/
t0L2k2FUrL8QTihMjPO1a+jcU3s7b3YjoqU4rNEGbqlzKPGTiq53fH4ITp2pn/HL
5rp8OFKLT8h7gT+nSjO8LhlUtFUI5tU8DnQ2xkvApUPKIAaJCsvykLJAQmRtYWSp
/RxVmYKZuwNhQKqPEtyKix/kVc7/svsJr4p8sB+jcjr3116f6m4Uqi+pYeO3brvZ
HN+fuJO6fqYYj6qlrTHeGnctfwmSV9oQzwuvpRKC6QMl3nOTToaWdOMWR5vqjUk7
u7kYk142lEPXm9X5hHdSHMNAttp8+rw1aX3y7xQmAfxvdDXYKr9BH1hChebvLpj5
RCg1CKj5XYSx+PpyMgNo8D+Axu8WLI2Fp827H51CsIeOYX1XGIGDoStGI9uHij4P
BsrNnPQz4os9JK3xc45xLGp0eQT8qpJ07zDMm0OXSYVjarCYPNH8qlPHAfV/4abe
ZmFAlE3x6onGJ14kqUQ40X8cQ2jXLmV/yUkbCGtYo9nLtbAx/efP5ilHU+cRawsk
/ql/jaqNeBkseyhGwK6X6ItZifyrIzSkE0yPN2240VisHvmGnglD8fBEk9Ua+sNH
MqlAZR5x8K4A5q8al5fhdzbWfewC5T5V20hXLqAVV+g9l6SRJx7UZ/+m+ZFi2k/c
Y3CN/x/B29y6qxsByHu7YR1tMYZ3/DiFL/GohpkUJITKj7ODz8Zh1xzUk6cE2VQ0
nKhaD/X4HY9yKpFlzcn9HXVacPUoORu/W36BS23V7xK161jEzZGeHQikmTzuji5e
Xh7Q4GcMitDbBcj7uqEseuZWUP3oOLhCq4tAvMBYeY+YmnCawRBPgVGBcJepG8GJ
VP89LnuVK6G4ghmmVWqBXXiHm1QmAaOfFcSLu8rPRhyj7erWpTeICq6nVwmHESla
uQ13HtbFdiB+g+oYVofsf88U7bapflyu48QE9Nq70hmnKup5Jhz6WGQIdPtDPqvY
BkOY3lGc5Ng+ttpWlj5MNe4kgmbImu2QaGqwz9NsB2OmlZqQzA9BI19cCLv5J9Z2
b0/BDsrI0V9JgtDhGjWBPnK4SsTmhGl2SfB1TPouuVewIQJKhdVxmSTF7ukFbkPC
3jMmGnoqr3Bh1VV33OCznN/v9Vvca/CSgjquz4fhiI2ByNEIPtC68rhQR56EXC+a
WTM/nCwBGoHS9y5Wv31Vu9VRjpBKmnLvX47be4CNeWtXO8r95ZbVa5P3noc60kBU
hxtH19WAoEVHWfAdt5OzJe+i1jMznpe6piUmQ9DqO3g8RUjp/s7I+nQbU83SSogA
6UwP2ysAlE5TkjQwZJN2Rfqf8fFXRcbJvDaPySlzJ0O/yulanS9fCHqUlnEJl5Uk
ATffJEtbJrdHGatxJkdtIvUx9fhIdaQ8Zpc6vD2rmBU+x5195gK7pajLzC4W+X7h
aU3ooGFZ9iFMYuguOvVgKAiyVqG4kYHba5m3vmeSnpUJL6CDFG0KMNqsW46SKDo/
ihYPjLgkkOlgD/aGUzZNbIbuyfbxzLE1zL0lWZkLeTt+e5vB3GqNDVRSEJIh//hE
mh8FdSX6C8p5DsAKuBsNXSINABlCEP50pKEsOO3XEf/SvsfhXZ4xtZS6OzvmG0gn
iYYM8HwvtZiVWhrXqPSRlU8drVHLPyyDsoZI06sawnrGucwHBqR5Fj6u0yQzwiSX
aPH76JMMK4xscWOkmVARYPfqcvUkU3EloqYFvB1SWsRhQe+o07WFqb/VjMxCkLkh
wCX7/g5Yn6F+UrZfdY3J7Al2B03ylrqR0iXpV5WQQi7rxxQYs4kocdbkBoCkgN4v
XGHUhsSs9xplBWixK2kbpakHAorz0j0I/EiIXnWUMtIMN9Xmmo0xe7Tlxz+dpm1K
joEiQfYFVVyszS/+f2vrNAB4Owef6fv3Kw5dx8g6ygSdrH67By2dDxDQMumg9J7b
R3NCkAy82jn8gnuyptsV6hsWD73mzQOjg4j7JDjgUxG1scNNNyR+4uExge7rle3t
4U1bS6uNZZwoWHRs4ABvNltzstGPQ6XUaOsO5FWwOIuCufE/RQ3N6t/wbjbRc9W/
Xu32Pm+Zil3E4vHhPizqYgCjA0WS9UrWd4ga1u3K7fC4BnaQFZoY3pFwIxI9+8F4
SIQq0qexy5N4a+opzrAAWQKqAee/NIpBuN1MxTk+wGyMk5KwQth9D1yNdDAta6Tw
r7CMNpzxLtDrChYZ4qzdb0RD4+LpY5JFJ6Ha6scBCU10YzHwPc1OEVESyIBK6EKt
tdAikgfu7H1yxh3TMqIbtCp+gy/+3sgoRq3rRfLeVOLO2n+yjkxii0PdIFu2yOUu
GlaUeFdY+oBnK9gKvKh0NqHv+GJPxj396tZY2v7ieV+QUu+HyhROoepTaO9nv3aK
kbQVJnPo1SzR2M0C8GM8yTIctjoykw5LXjJLNBB54uFglvT2XoFC/YjR8QCA8+RK
2G5jGTfa8nbZwQNCrtMam1QiHmdSO5M0Zmlqzyjnk+Gi9AVDicWFNZnNNou03cqW
D/siocV8mVDFLmQ4ZxaYmY3IbcC6dOkV2M+lUG5oTiNWAkzCP1fOBBQf14tuN0K8
ciPYPypPTDMi4q7xPzDv9sOapDK2394F7Fddo6ERmEzWFCUgubI0iJjockj4XVrG
WW8lzAdWjI5EcFfsXrjcKq3oGEjemDmjxlxT7zQnyy7NdpsMF3/vsRT0yv9TgMWM
vhTwd96t7s+Sy6MX22vckeA72KvAqI1RFp6b+MUdKmKIxqvFuRfKiWylbvHWfTzx
xFFxAnPbDa09O6Z79yUWi6CVQg81VzZ05cmluMENaZSXnSu7K5K8Lb+49YVRRJLS
mvIy5jbzencLgdeYwctGgRnkZl7yKTR1LjENmNynDrBVRiLJPqcTgLOAA9dlQ7fg
IWd5PxhSZ31Z5ayPyZhATgmhOkxR+0FfYL55iyBwEsCC8tAyPIZaMOUu61HQB93e
0p2dmKwnuCEg7DVVVDMg/U5ArySKJRMzvgRFsawIehhASCRJF+QkIipod6YpLPqh
KrSPREpAkYuBy0ODwctrl2mBvHeWOwcduB4lhs1bJz6Cm0dL1OEbE7B4Od1wDJ+W
MzwaGJKHY04ZEoUrG7dkgSFey6+qAmAJlzyc2AW0tCP67kqotqb8t0ShbUSFZ487
MLMUlONW1ZFJsPxOZOK89O5jwLsGjgvMNL2kQc+rY+j6CM5WkgfFMiHlo0CqLg0G
8K/WTbfUbHjOy/b2OeTHaiT6u96iuJbrRwsAMH1x49LPMf+Bw7J7qvnjj+1JM/uj
efCIg/vxCMhGW8Dq6dfbtFWDuQ9rTUNmf/oWmjYG7mrw/prblel9lWUNdyhhD/0K
+G6eUCG/AzUgLH9rIzhAMN2L5vyoq1slwPal6Z5HmUnVUjsgpZxl5wknjg1aYJzP
tCyItgOpNKwshpsQe+q6VnOETrghODmM7ll3PTknreGdoS5TL/aNOAtyQQBap/jQ
orsTtaxix6mhAEJiMOy340c7+/JNmIqiHgeSA0d8ezvxRmh8WzTJIFNrdzoCwJ7r
/8sadIhRCPwyfL6j+ZMdWl5jPnvUfJTkrTtpDIlWjPWISztGBUIB3/4uq0vP1RWz
8cV2S5D9nrYvnymbQYq0+McNLdQnO6WMKfz3fA9o3/8q6A2z8xrguCuH1Ei4jqgw
ydsPDYlgU0VZPhg6jgRlZFIMdc4QONmvRosecr6zjpO7YgD9TXYZOnV+hf7TgjWX
c5D7foCMrozj5IvvZ+IyqV5++u+MWeqVjSTUmARmhnhBa+5tmVEf2OZ2CpBaclcy
2qkN5PWf2lZ9IDP2aGPKA7ezQcE1yjYOp0NydwKAOhYI35iDSYMCSqhDoCbB7E8d
brioJfOR5h8JlZe1jTJuOZBhNrYpZ69WINPVbjNJKlpZU58C9XW1G7Yh3UwtzUAI
ieMhNnAqeO1Lmk0Zh5I8wH7gn5BQ3G9JNl0EATbS8HJ4WSnhm8fMZCUb6L75YX8F
Y0cRxxXsdqPrv+ta6ByYDu4wbRjsnt3a/rhpftjh8lv23KkU7Zay7mmi8knCn7h0
SzNHbc5F/5XBfHRwrH6BFqdATUqTt66Y7vX2s6kkGif0e2VCSG8H50JLfT8q9N76
LyGQG2LN/hJL1nSESYieXxDClfTKW4IrFL0taC2HiGBAduazMUXFrDzvuhJVE+0e
79hij6pM4Jl1RfxpcznvyfFa9f5gIxdt8HZVROb7BqqtT2losGlnhSuJvOHNlDil
OTikhbspYGCAsr7YksHTMyFr6wh2AsqCgf7ShbMWprCOKyN7SkS+AuFRVV9QvtAJ
a6VJ1eVZF2ms4F7JgoMpHlukdGnj7a4FAETkPkLIivl0scM+s7KhCUwGfrnNysbZ
rjHip3fpALSxt3tBvjeUNk5Bj2hW9f9Cdw+r9fVGgwt44X+6DFT0LtT3pYL+mCJY
cx9pikBLzq42cBXLtSJX/IpV4Klwo6dcH7PhZScC2BmqubN5NSADrC2B26pzFJnH
Gdd7qkwyqgxpRK1SrdBCVymTv14BuuSA+7KqyFn0xoMtDWR6H94eIBhU6bqBaZVL
GKyByLrq1+aJH2frXAZVSV3lD/I8RgFZ+oBYFy/YhyTbAGoGV+lXz4KTOedzutuf
6zzwV2JKhbZN7nywNQzScdoY9WCHcnLOWlEMMT40nqw2S1nzOntHf6ez5g+fPjey
gG8Mm3w0+11GFUL0eTJpGtHGs/xwyEfxk3kxz+p4po8OicwgzTAyeqMK/I9Cw6BT
lLTyaT4zLxm/Ll2xuk/Jsu2w3+BC6AOkn0UqUtaOXBAToKpH3345SJvR8p2z5iTi
GvW8A8eIAXgaGryKLiRQ9YAyEMJXRyCYK582PIWNh6yk1lfft5yzVhdwtw5EjhDB
PYFh5/zFrqiEp6pNJmf1EmU224KXcLQcXccqmxtS2vqxRXkdsInZUwaXXqmmp1ny
DgoM5UNybGfpbuaA/HWdANqgcHZ63huq8aBtXJETDGhc6ZsegewXe2gjgjwYV1oe
uBP8Besh4lrDfF7wkOpDyTWdhvNXfoiyqZcrjOfpcD7rRJgtExcPJpMGon/E/708
FSp3rQGXdvM3WbKW80K0ngwLXCeTK9h11L2z+oJEhgvCp8npPGoVVszthXU4aKlN
t3e2ve8lzspqTlDMLAsGvpTekhtK9xoKl47vL9ws9y6WrL6P4vIrxYM56pJnz7EB
X/buP9C6H+mD3zh4f9okCNSF0c2zvv7bvteBF3ZQTKv3Md6ioLGHTmY57XmLJfF8
5ucXIzh8IjMklQNkPmnzIlKyyfp3h/rLuJ6jiQ/oeEVJIHR8lvIqVVW9eyeu00Ec
jXC0fOyjY61teRIp1plFB2Twx3jFnAKiPKzVRPfM/YV98KnOaZ6X6jbAG5xSvDfw
vo5Xt2W4gBIyIT77FpCnNHwlzM3KrxPOrzXvUKpiOTgOOFC5DFu7NoyFWLU9rT+n
ICopvJ0a5SNHmbeNESyq1FcJ7WFi/rUJE4ZqW9hGHVYlRziy8JwN/DUpa0yKzlwI
gVp20eIRRMySpgY4IFiRT88HaXCWTgk6neyirTiuVj2PMCfhz63fjg4rJO/p23pd
mAWOqAhUfV5wkWQhjAWPmXFuQasZApDKHvIYukiLw6FLq7Aq9QijvE1HsRwOtR/x
SR3ddG1t5qq07CmCtr5QXr9/5pAUF7iQGlQuuk2eobuOGw6Nc//NJDzXEAsqLb6O
XEO9rkJsPsfZFpLvQxA4gaWCSwzDwfUTKG8RG7ALwK8qEfuZ+MdQnhWhmPkLo8RS
tRQxFubpimFiEmHBR5ul1Ua+1QvWGuTwv9+hoCyC8/lz8nVaK9mrykDZ9Gn4OKwB
HBK7bD+wgoZ09AmJOGPg10GW0d7Nn45BF4FXKKN+HMJN/qk2nS2Vn9gHPAKA/Knu
Nb6jSy3SnzLDfaFm7o6UJAtSmgFQQ002XrT9UhtSLXJT6oKkhtyTi01pwMQ7UcAN
Xcz33EiRZJItnb/tW7yQ9M6yrRQWxbIiLQ2QpjSnsoQfxMTuCOujWWJc+xYHMNI5
5NHl5Y1zKOrO5mG4tMlycyVY/6N4jY7YSPjw74VHvU1AmRHLTnKSEGu5w3SJ89T2
GUJVcFM88MwHu5Gs+nt8EDeJdEf1ZRRc0sEB8Smf6Za+MMlnjXSvhRpmLWwvDP7A
mhMPI+Cj1nFEE8Rkd09aJ1/W3nvAnj7faiPF20HZ2wRM8600wffl3ebkhuvaUxCG
LrNvK6FTxLm07U+McT+rAqmLD+AzGwueP0+hyn3kfAwlGOQvBexg6wSAli/drbrV
7dS5vxThssFYbnsPToKa0FaBp/oI0LTNqhqyNjzDMVi+FCt/AV5KKV7AHPY8AABA
YinG6aEBaVKr83HFPGkBRq4+txBq8weJApX1rFjm/C+XUTLIk2sn01t77q+GoADE
o0porjgZcETT1FuINSZO4QujPRohzbD5t9q6BPzDj6K0Ld6jn27WYcu1J4l1QjzV
yDn7pqxDKByOG+NQd3tg0LObhXZra8MVrNasjXQIhxdqBBwqSl0ddA2zb8cNwzrb
6GMfL6k48NE9bnHICKnx9VqkcXS5Q21SjJde5cISDOqhlmXiWE2FSmjhtubiwW32
wWc+J1kDPjaxyZVSCssBgoInTjxZsPLfiPxg4mPy/W27oIbveRSBpBTHzbgEONrk
kbYOPkrhWWplZ2xnhHT3Iu3syda3RUDcgazoUDxfNQ9cxXspFBZ4estM3QmB87aN
iWgp4qm8/AdlHFiUjXoxJ6lN4+r+YZejtv6FvgyxSX3ujtFzt8SLcX/3nPiTmPb5
2S2IZsf5nuJcwvjWT0ZWilwvtGEGCAFKkZ3QulWxIUaXXMfW+a+REQYsSmGP1vus
ewfQRVhTig0u0gWtC6Gt7ZeynNGfyqEFlyD7zx66tkmx0V9o2QOL4sXdTaNTJIG3
FMfL2FBMHFaHZWXW2KGKfMX9Xm26bQv/XiaczHGtY5kv7y6wc7a9rrCOeVmHqqEj
PP91/EPsulo99tOI1twpq7VABt8Ftd9aD0bWMKfjQNbHbtz+wUynsNuskqNsPUUC
1PKb8bCKRql3j6GhJ9faQXOIZbOWqttXtTVl3qJyZCFAKW4Ug+Xb2ajsKRzvv/15
5kPjs0Mt2uDf+y2f8vRh4haUsQw7Es048VoARukHTtbCMJL5LBjXf/65rOby9O/A
7XmdPKIkYhAEZEtnTbnj5q1AiGdGDWGtWNQiQTMdJDKm/f3Hx3TyDgeIUBsNFXDb
idehwuiEcSEpA2KuHnuH9Ze5Tf5JaWTvRJQjgDcIP8idDgGgzzNH4k04X6fW1j/5
WWQbl9T00XCsxCB1jAXkKUp+48SdsElLx+ycvhxfH3DRfyNkhg2l0vrJcmwCgf7G
Hbj6lOSpPUz8lk774fiiVtNEE21o+ruc6qoBJPVuFajbNurrYkJJoMo/jAiWzDGs
JuXQkOhJKr70vZbq9P3fkYB4k/DRIWxw7PoYlziGo4ZhIvIU6i5NTW1uuWDxHSs7
9qSBXe0MqGaujaMaLjn9q+RAySzcdVmKW9g6LDdQya1Mz29IiCqqzrgDxAaYJZXh
E68gUPvjwU4jpBzTGaE84MxBr6iRSLwK9OfQIYYEja0QHPYE2l91C7HG5xwMWr0Y
jEOBXFbkHZzATCImP81Ds99XbRcO5YT+GjTRhBvLN01oabMfejwvqgujoE4Nk+iH
s9ZLc3ulu7tiBtZt5eF330Qq0v+tsE6c6FM9JgLZfMWDGwt1Z3fkL52JRKyCDdtr
+kZzTINu+PbZiy7oG9aV9+zM0XldFUb8itEziYAKbr+sQ9Mx2/60/rv9P73QkE/1
ZZikphJ1ucVZiq2EBP9ONsgckVAwmuqykX2Ba+jvlSkq0tVvd5w3BQ4U7vUHTdZl
BmvuK+oON9/5lMf4j3C0lc46Qgg2spQXw286vcJkVD7aT8fv2CXPZGTaE7igxRyq
GqHBxwLw2XQByz4Zbnz3TrubB5v0KfCD3efWK+RtF9L5mTbn99HDh8Y2MP82pDPZ
CoDItpaomWCLGaqKg4yropaLaMt7aI3YEHiqzZZ+xJSiVdc1NhkUlnIVgxAf4osH
7M8hFWdniwwnAb28zz8srmyNrQutRfoWhNMvVXjTxBBDa7j9QawlnKe7t/X5V78U
xsBdpSlwmJSSgEO6BTwuWikjFpFck/9cJtXYBPitGuGpsulibC2gVqtfkuczJOcI
osT7qNh3q29OlJbUJhsBuTkdUCITilAfMu+C0zMQz/SAp/rlB/0HYUqkE6/Gn6Xn
8zeufrkjSzsdV8ksh5xJYwoOphC5T/3QQoT6U6nB86SeJrzPjjE8c4hi2PuoZ0z6
brQWynye8/hzw3w2ewg7TIXxvwOibZU0aX5V5sn2lt7ciH+RHcQDFCM0LpHofTjv
FTJWmLENVKz/IwM1wl9Q0v+4vSAkgqSbszLCUkLUT9nvjGr1wbKhdkuXrdAnvgxi
68XgrRu4bKo2aScW90vEeX4PImLbMqRnT/2+pVAF8t5kdzUDju9cdktjFnXmxJyr
Kx7lJqbVHhsj9DD2/v16JamJl+fCclR2MKrzu/s8nULf7Vcny61hh5Xr3OgZrRp3
Bp+HGhmnFe+BQQFmS3lK9JMSt6wG5Zx/De+Izei4uPGVQ3TZKfeZvMnmYk7ziHDw
XuZpT2xOGW3opvVLX88Cp/4qzdaKDSKsTkHy7YVXVsAXb94bF4WRA4xo873pG6G9
7YKlCtACI58TP881GATCgpEBTQmwEjmfIyYDfU0bdfSN+ueOnfbIHRRIBhyiUMuG
CuZeM2Xo5SXIZ51b0E77fBDuGVeRQAnQN3zc1jmWG33iOuLF4gnCoxcgmvrkJ6Om
aCsrRBGNzCE3E59HbTlCXmpXsmyt1M7UyE+BhI17VJiMc8xuwVqr07R/r6JRo5Gj
SM33fCPEmvXeX4WOOJBPinuvziM78IctjdKCvjaR86oYJmkzMKfsGYvpk61MKuhu
xsgB8VBc2R9B+qxllUkqS85HKeTfxiF0ovdqJHz0CiJr+W0naEaGoU10DaiS32mS
znKuTU3HFlZXzFgzcScQvcDnjTiSDIA2fxpdZH4GUj67WLWQcbKElEqQDBN4xPRU
lfdpP/4La1Ua34SnSJDJ6uMQ6y2nnXT/VipyrSpEf4Ys+zh9R1iQ7zktHBHJHi46
h8T/u7GKaTJPY/g0aT2jAAuo3q1oCguvL9V6KTfIOcn2/Pohi5eQw8hq2pLBpiRk
kO55ULdad31RnEJrfGExn8Hi40jkJRV54x1OkuvM7CBiAlSx1r9PSQ/ZL5oKbhTq
Y3uio8SqMcAth9xk8sdnMZBxu8LBOsJUrP3q9vX5t5qyBWU0ccdJ3YtV4H38W3Rc
YdsVJl2F+VbigC/PhTfUDBxzYQ7/gSkHIoFAZbwnubpHAaMrKxXLjJRQan9nW7gI
e/W5qC2K5Xf2bxMVLJdGQM9U2fIuBEqr+Tk1lEQn0zJL3R+k+cSgmUxMe3UdnsOo
0FPmzMADkDF0BQrMXTy3dC8LJFGjO2SeBeRuii+zQ67Tob8IFVGs1X4Cp5p7oZif
qHzg8g4P3myZlfH9B6DMuZTxUP3R24WPG91HetNNxo6FvravFyyTuxXF/grqADwr
Fbc9GLSfhkqbglfrve+s8C7YGVBSz27SCZtSsXewkqHdHQOh3jSZs1tmH0DiHpvY
hmuAYMk9cp3Ym5uhxmVjrmZagWP2wK2lbO4ybJZqAnndO5NQm1nC39/y5lewbkBc
pK0ozik5J3sLHjkxnSaI1atGZzXY0VyIoziNqPjbU50zJlB8g0TW4y/ZgPlJ4S6w
WwX7ZaGQTV81nkuXlts7GIx5Na24Hm4Gcq4QX4oYwssXaq6PWJamWGqN4LXxw1uT
I7Q8Fc5WrzNVIQe03mAV6KyF2UkDX64ZuiTChb7zcbf+vBUEbtdU4pb3BCyEwvRR
b+dtdV72hvlezidRf66SNdTg2Ce1g+hD/UhSyoT2ogkwPVYLiyC6bzhRQsAIT5p+
e0sPKs7vA2dE+h/bi2PkSOQd52ACja6Cc0lZxq3goDzOQEtuK8AT6Hx4NjCxaTjs
qtuEPwOggOR745SSKPTMApkQFxVSM1QVqjl8uLn/DAPf/xrGwDa4G6Vdlv7NVRnr
IpmCqAQh4uSZuxUus4mwItCL4EVCEzvpcJkk1j66m9alPjG+eQ1IvaHLBHfyahKv
eR2c/iqdg8zGTnpmys9EGNtWhsBkWpxySRwxH2LHgBVPQKdqos5d0e9l/P4/iYCE
DrHX+yKjXvMP/7gAmRNa6yi9tope09cvFRxr7wv3k88ld+A3L0K/FX29Ap6Ye/lo
7JBt9hlqS4JdeDEXCNke02Bkhca2SMi5QvakGRg6869NfLjREyVIeVhaJ5cbWT2H
oP+0n1ahNgWNe4DuEFRK7DtMloQKVqfKfzOhm20xEiySn0V0ILgK/AFbR0SJuzI1
jLNbUHLohkfQFm++pG2SjIo+YAcw7m+GWCu974wi3lw1oRO9tpBwG6ZheH9oXaQt
W8aGEU9g9/oFZhJfUArtjLnzZAP060IZk7XP4nvrxWyRDlvSd0Ez3Z/aKrTubuOL
ETp66Jh/DxIbAKeF3XZ/sE+Vr2POMaIApPJutJ0louZWxh4FmPh0GM7kfmPCScr9
XekWeWMc+lvNmCwPTNqvumD9xJVg6cr44hMCUXvDBZfFolxfWcphYQRSjm1QEkSI
ihf+BKTlAvO3mkcluOGYiCn3/pgQLfS2m+60MTOQKHDDjR4d4Xlrl6IkWovU5FT5
Xl18OKpcShPPKX3egWgHthFu892PVjV3Mxp/rGjt9sb18m0faDLmh81WVR/MSBoj
I6j1dcl8DUbINIkyM8BSNroNJZaO7zMU/Vka3g2CDrB4fKgEFO4pKJ/UUJqhopaf
kifajqnKyLUave3pRaYMdvHoB7lsTcaTB7PwmGQi/7bXjb3l+rMkOwctGsbWQQV3
cRvrvxLKXN0jmYAHCCEjvUCnipPTK200+77X0HRkoMmPYZahVMdNTuWs+jVQlTuh
Ern4lGJbdA8NBvta3Vq878EVB9YNU66J3j0faAzOJhNYIbRfmoayayB1DY+jy6ga
8PKvuHWij3i/BHsUDACGycFWODFNq8p2dVoO3EXkDl65Nj4WOkk3JqMSkPU5icPx
oqVO5txsuWiUXtpwvC0E1Z1asEtW78tHJKdkKcHLzb84ktzCW5pv7E5c3ZMoabEQ
QQB2qPfBZNVngsX0cx3b1+cYQwXz0L+O+147KCi0ldNWZ84fN3/bbHTwurD6onCn
S8VINOIdJz5rXAKiPSkeni/1iPIqnkXiFGMVDF2lEZGCB7bazoT8Y7GW/Dc4esTx
APZ3J7z5vj0QLJ3x8DJHnQk7YrN2YSBuj8AsPUDGrc4pq1u0nktJ8iwi2w1K+n38
j51zm6382Rn5LhU/3qT8cLIUJEGtgV+fR5Wn/Lv9mnWrFWQzlEDoWSGe2UlF2VR4
GoMxxG9XrpVqBKB+Mg8YdaLK6rl+djXtuhyhU0X+Z4YcHfqh3sffibGYAm+cc1bt
zF/rShhK/muogthOl+54UdXvZoNkCunplUrFp/wVyle6ws9q5TpRLquLr5J0I2/g
gDZejqu+IuVjYDpEbwcrpyyhAY1mPj7CABxgTY+76917NI+3CWLAkq2sKB+uNJLS
eq5ffBWl/LFY/yb8b5GErZULlTYGn/zDYDc2K9/5C7I/qBb44c5dALHbpHvR5GON
VffxgoGGtrF88PqPvDcBmPIVuVmu7m3RAKt3/Ep4kVuuzk1NEdFaP6MbeePW30fa
ojFTcg4UnRPMi9U0pw+jzxluRKp97YrB1ODA6/6jzTrrc5j38JCdFzDFek3nqRPr
sb0zKQ4GOLBaYc2hm9nPnRrMmMXHBWgwl+fW4pGblJp6AvHHsnN9MWEF4Gc9lMCQ
a2dD5oiA3VbOr6U9+fRGKsyDUir6CQTVG93vhzXOIiyXIRLk9TIC9Ct7YYMVQySB
5cCn3g/4GZ1lIdDBxEDrqP+PxoKXDkLKx3ltzlt5SEJB4xKTrJgNBhc/0UONt682
nwXsDbBH7Nzps6tEzbJLh3qVSqPnBGwQ5hKLuZzXIoU14Pm64ZEezZjhvaD0vXO7
ocnFKdS5oTBrTUzDK8u86KBdXliQaXZIxk7P3JTX07+tSqk3XNCuhQioO219NzS3
l5XNnAAE5QI2YwYlYNnYmSgsYvddS/KGhgDqNeKbsl37bF0XMrkMWnGTAhCJZN/l
oj/Xw0QV85cn8aM0y8jLP63lWtyoGa3jMHEmC3J9LLZWM/qbD0cGF2U22Ki0Ld4y
XU5PrpYdPJYOaU4bEiA3KsaM2cNN24sOf5+rf3nC0bQB6FgVGkDyPFAcbQCAmrpp
LejPuSybklVAgH+y/5cZTAXPtRMTH1W4tlBj1UokAX/OyoadqyRfoaA/ot03Dn55
F1jrrjVpO7MLxS1vL/XZK6wh0GVGxHZXicXoOFPahVo+NmpYx0wctX+cn400Fs+1
TgMSBPjd480lDxkc6xkZek5hJ6ls9BWQUwws76CRMUJdA4qoQi6turJ9O7OFs/X8
2gVI6Ls2nIJ/zMRFJwrlU6xIjBQx+gvx2LIqDGtQZO6N9pHL/u9mQvbx6jkWm8au
qf3dwSO35VX8pa29rqpp3wqjCTxZvg4nk8Y/LtdGEd2hSsVT8g7jwRgLPvuRupBM
BAGuTQ+xfK8YkYaN+9N8xF8C467H+AO5ljyIvrGLolYYAkbPtkD/OYs2Uo7q39ca
OJnFWuAukuX+t1jnD6BEOQM3Xc9oZliFaqkEAMWO+aWOWemGVd068P9pg8ksyngw
bjnrkul8oeTJUyC9WEeCV7YbY8B9sn3wDZU9BTR0j/UCdvbKJnfkJeCUi5+rTeag
UlOKkD6ps3fwL0dzTlHhwNSNPfHFgbTkG4P17X2rYa/vuCO/ZbntFQXysPIx4DMb
zuQZZ5YCquhp3nSeyeumJuCRb5YRUhhRqKAqQD4VWpXOZdPFFrjARiePHPXrpuan
Ydr6zqBYwQpe+1SjIY6AOaRrAcqEb87s3kdI/h3qxvovFieAn0/ajxAfp7dgFKDx
AmXsMqMD0OjP0vcgVe3zBTcXxprBcDNpG52/0Su/RZkrn5deZiv7OQdBUbz7zlpS
1StzFnq+GzVmz1ZPCN4pY4tbO+VsA1GS4+js+X0q1XXr5d9j2zqwdn8HyDV35wUz
9PXw/vsEireb/nYD6UOBj8TzS3dXsgML9J6fJBYCWaIfB6B333CMEUojlz+sOTvb
xS41IG83AbfaB8D/MxOogWWozszb5c0+8r+XgeYFcWWRFS+EiJZQTOb6Yhi2zQ9W
Cp6/G+sQLjwq39WfUss9mqgobLvIm3vTFbapNH1szMZSTOKf+chjKsZ+3o5SuZbH
nK54i0FeOJ5nelONKFyJxbg3HjmRTDwslUXmric2uZ9t3QO2XAIUfFRYu+4+vkUc
U+0WdrH3aPY8Zr1jfm1hVF6D1ucg9sPzL1kVYelnmS5RfpxN/OZnxkGXdmn8RF93
DaTs3M2fHO/3C4vh/CjP3RKou/HxRhdjFZPAvbaYCaW/UQurhzs9cDCDMdOp0Lj6
0oBc2TLqg3vFWtPqw0VsenfO/XZqzuiCEJ6szarB9uQE5+zgH634KJZQzHkCE9Ce
GQBX75AGXxaN4EyetX7O6hPOmSx13Kpyyfi9x2M+8NUx6OMTk38JD18l43XMVjCa
/zhD0Zdx1tyz+dndrjijUnbl4bw65wt+vkHEc9WrDCIGe8yvqTkqADDcMdI08K7r
RrjGeDrfWdTOgOHkFzvJSsehLZS0CfRJFH9B/3Rha+3eZTnBFfDC1bvHf9/UZup+
oyBAnzqEaBcx74LY8qVGLJcMwByVcy3lluZkDA3ghFJyUSyahz+gkFvGqsr4rIyZ
BmTol8Mayz+xzXVNE6iEL+GDQ1p3W9MfjU+H+4CZSrOGAPPmMB1dAAeasKsGmQ88
iU80v1+HGeN0mmfm3+BqISIYOSdUC688iPIRJomMYmhWn8+Y1dFxPghStB9EO4em
H/1SvoIY+qeRqRpwAPE6zrTZwQA+iv2IXZH2k0SENEiRpjwvo1YQ1zrv8SrxziGT
VuRFztH1nppPxpuT2/9J8uuYT5Xqic1WEbUyi8cVpkw79O/xmqD+yebLGizYqpZF
tVUT1ybVcTKgGXb77stRSUnQB8JMVtImAl7k4nhdtyegrq2MXXyqjmrMbDnrx0l4
EjFTsSFQXjICmrbBHGvzV9W8CKvnWBiZgiSSZyxbz0bQU9A5I/gpt7QRGDAfex6t
hVNhr74nP3he89hi50Cp4bt/uMPLv+Ry/0y5SczEdg4wpJcaOILV6KhF8XXAeHSG
2fYhGkzTdIeOQyTvrkRySou1OjNIw/PJG4fmsQcFaTymeestDtymtdTg9xU3oVOz
je0MXcPystwRCOkZgA4twTkfBeCgCsPMGVA0LU9bAbO3J89kPSRu0nBgeWUW9g4V
c35RtwCP976uSFuX8PdbXW5ntGu8tkBid6D2iSAOP0ddDaJUnagK3FyfTEpw4IC9
P+4t5PU6otbHI9MFev5QZjoZJrLJet9UmqLJ25wgBGH/rLk7VWcMukwr1xmlQ3wu
HZ+8hP4sxWuHUVnWPJ+tn12YTgW8mSwZTyTlcbTmI4LHvL6dcSDv8sG+BMXsJOiD
kMS4pS0jPnz0AjQaJAMU2tof0a0Pxo9rzdagdSpeKv5Bm9ekRvEhdo+D+yXV7e6z
rPyzEIuIHTBanSdyTbF7sAjO6je6SUYWB2VNL1POXyjhb7KZLEwNWWVF+TGN1HSB
meQcKzNok6la8+eabYsUqELHH6nZbV4SLP1QavX5Xbgpp7tM9aK6tulRXNKzRycu
lylm1rc5KM52qB6dDhReFzj7fXczCWYaVPr9s6uTPFiodqjFlHzEidsqFaFcEslH
aUxXgN0gmwoik14+Urmu86oLkx/I+MO2SYY/EBt/soGwhsBtVt649XoZWXkNeGuj
DT3lGSSXAmvbpyNI4QapBWb657XJRqlZzperKLIHOOIC1p1LxM3qkK4vXbZuthN3
jU9/oaI9zMPc4Mby+fVFtl9Y1J0XOkM6R63S4+n2bbGm631erPVZtETDAF1pLEtj
vsljmIKzR0NvNoRk0cUwV2nhfhKP1ggqK2fEJ0DY3Cuat49RvAHZonZJsyGE7Vtr
az2ETLZGMn/8Vj2irPLChaND2dhRZmqnAyUkiCDifzqsLsPWfS+JsPOSV0JzhYsU
eT84nDqGVWTW4O+/SK60DXEWKO3CYX8MuVFMRhtRfjtKUEbaLyFLu07MVWz0WZe/
nXFNAIBZycD6tilfGWUHxiVM9xXEZ0uCFPfEeJX7yi3uyqWKfR+uLwjHQd5Ej0LG
Zn0f8ig2TSUVjwdlfqn41fGiFMfWXyz5d2nrlXQXZqmUgiVGLKhD0mvBXRj7wJpe
zltcPXbllq0XtA7Z1koCju7HvPNUdsAIFPf/htquh42hFGJ8OV0UMOPgHyL1OZDF
w9mwGuCX/mJXBdq+LWF+aEakcsGfEySc0Z02908YHoetGEa8xZnH/RtJyRMrfMOF
6neiP028Bvt8Vq8q5U/JWPnX2jpmZToyslHTYVud/ECF16r77n0LksLyeOgrcEke
cSOOyBAqZZ5EGu1N3Ab+O5TxLRDNioHRb+CMW/Xpw8S9La8Gy+U/mGO5giZqsIqm
QsISQyqEvNVDVn2dXJx03cZYieI6L1K3XJxwmrSznLZycyW320kuRtF+SNrzoi9f
U25wvvDyETrkdtxmloJIjiVj3y52u/RMbwTajvtLHWiT/VM9iFZrOdrEU2wJGorA
skM0MTfY5qPGTP8n7q309mxQVO8dZWli09sY/Z5g8xBmZdc4qtsBVhZ7OhWLh99a
MjiTURTsC1UAkD8Aw1J7H3CYVfyRxVdoU8ens6jZvVSXL9T1N6Fdw5OhOMVngZvg
L6KSnO1B631PGFveRVacRDvFDiNzDJc44Y7pcPeW1T4URN0fJpZYMYjCnKL2N7l1
6oz3UbGj2jL2SuaLNom+uvqs7fs+EuJ/ZdAAwZkLVHOW499/rQq6f6Ypvtb7mt9R
0oDDIZ8o+/KK7bFhcbKnF4/ZXHA7tlCRAMXMYdHar/ssZjj+mQwBc70slInnRclW
53SagBHETtO5PlLm50aksdIMvKRhcv15x+QlRu27LoHqljV1dGg0F6TzmuusnAw1
z0BfEY7m+rNomSunrgb/bZhhNI9uhS7vHdYNNPpYoFxbg0fw5uSimFMUY7Hlla89
ecHNATWc2xoIksTnZq1tSVJvNvkZbYwpIHNkIhSKlyMURzytJUcjZToRXoZAu7rr
HLS5BO98CEAntjmtyu0ovCSeMMhP8PU5OEkhZQVVbz5peQyHHlPE6vZCp3bGiyIL
rz0Mo6byTlSaFFMHWllfLz300I8DxmIpR9lVAkde8aXpLFW8H7G1FEIWRsfCREgQ
eLfjsdmSgvuYscZe35LV7ZQuBlPbRV+8mqLh7aVTRE3zhxqxV2qgYYepsjvGyUwZ
xEqDw0brBA6zKbXh7pWjg0zq1BWmA1aay6kwruKG8rvoagine/xbHB7eYm896g2z
rmxlpv603PLCnJ7z7FZnh2vJW9TuKFhUdfpsL3KtZuW4uybja83p75Oets2SnJaE
JYGYStg91Ljh7y7O9eVDlJ4Uq6km2aA3O3QXPMO4w8kBQz9nuSmBCczmgWzi+R/f
ija1rypHsjyCpmvfVo3wCHuLq5BR7qEhiiz4N2jCqPqhnZ9QAxboyUzoLvOApzg8
fjdSNi6zTuCo3fvSmblJE1uPeOoo3kHa3Us2OU4Pt+e3Vjh+FFzu/FDp5X5YAENS
RJbRnMbq/P6CeVumA8z6t0j2iggYP8ugV/bYsLiuohqpwg5eOl+O4hd9DqexJQ2H
f7V7yt8be+uK4sXB+nRJMRHBD5IPx1s4+Uwz60P56YmelOqhGuFW8yqkjOogAIBY
69UtU0/84cxVCgoWaNFeCbf+irKZVmyha94f9hB3Ej+fbtV7P3L3Q5niVIkkL7cw
VoorV+nuuH3kse6vP/MB1yWpxYtOjazOIqh5LagaZQMI+lxL+adM5vfTyfMCsz3R
ikHsSnnJ6UaKwT/m+rarYFRbC4ucAPno4vAZ5XGKWd4HhJaZdqq+82wYcs9Tz6/b
TLsRlkP+WgX5Um2u8pGTM4kVjTWOQU5D51YGbyGbanN+RRT9kVFWRaMYZF0Y4qcQ
DEe2omqY62YTbMDNmMp3B8mChCwEPVrF32zyZ1/13o2lriL7X2SBx1mrneDOIKKS
0IXcNCv8k7CqTyOeLUizUXISiKVL1+VQ9i/uYUdS2QfwBTG2YhcRFCarT0i99Ksw
iv9yNx2leQj+onisPcasmYabzYZWy4G+OZFwKZirEqPG7M++Q7r43uLPIw3NuCeF
viqDVzBVCFjh6GfHjloNo9vPSAn+/h6FL2ltWYRoQxksiwlcmDSymDbCekJMpC+X
WbvIBHSna3Ie3KMm0HsK8w2JwC+bGxSMNe2JIwnZZmovb3JfhwjqREEDokEpFiHE
ulPuC0cOnDbI7Y3G8eJt/DLXf3iXLw6gaDTxmE/uJ+tR4VdbDAqOVxR40252pKFj
xL9JdttG8gMXcd2j9YPhLcdlDmMO7muVOYzan89wKIoQR3OEHrCHjFxJmHzxSCU8
225IyDPrjskMU3QgcweujDVIzv0HybFuOGq9cyyzfytnXbOdt79bv9qRn5TB9X2k
X9CDRi4O3oquelhc3xx5jER1xTkK0ZzlQyK6zXydXe7SFtpRp1BceV20fDm2vWdc
sCAc3O+Z7oDF+mu7ejdGPJZnNvSGMTjlY8T3Z0lJiuZbE3nlvjc0UOWWLkQtYfyU
DyLDmE+U9fmZhDQoLQu+VI9SmQLUrXDalQHM10KOf4swDmjMkZp03Ji1p3ZbNpBw
tbtqkoIALzbvs0VZRJA6p34RlJgG9Mfvb4+1piyx7gfUL0XJ8/lic9yB5Eemxg0g
DoDnQ37vHgKPBdw4Lrsi6xrqq2dnRYFr6lay3IjTeJANN9WkmT/Ulj3WuS9K7Z7A
URh0W0FFf55tx5TOMHx4FIb1eIRIf1aUWMjGRQVpjYx/7fZ74eOb8I0kg+V05qvO
yp38wnDdVV7MaqZXSxIunYH9v7vH2LKTJIT32ng6BIauUi1mKXKHzuZvfY1HKGGY
+TVetG4tD0pLYQbQPoD5hMSb0qrwpY7ARSFoQAi6s6AvubqqOkwTZ6Hdiq9IvppE
VAbZS/xkDFTp7RgMaMDk6zg+Snh3TWmoQCcfPXpBKQL/oNR3RymkDJ7gAT99vpnu
N8gIPLda+VaRJvngHjTPXIB+ArxMGmYCatqDV5HhXg2KmaECi/haEtZFa3JcW1C8
VR0X360YUc1m1PkcowU7CwT38jHQth1Dv5OhuJOuarOmBlTV3DU5+nDtbH3NcfAa
uspIyZh0q4plGP1KiFuerkXapblJE5Medb71wadyXIwE8to8brGHYsUlkE7NNsdI
JEkz14DBMdl8LPX9hHfFtolznN10rpIywVdIy+enHFxwEdlU1aTywPmSJ/AGe8g1
dVYYvFgZKp9Uc/NeWiKHFhKUA41+Hg5imd9Tu6kjdTXRPfo/b9mihENh/mtZOtYK
IsNzzNC8IkGCg1MaMIpC8TgM1MDVVxxJoww0AfyJ8cfD6k0NMRcHn5e+UEKqyNvk
ob+CzvULfwPFXHA7fvt10FqkqneORN+8GSf4LyrlhjtrYCnp9JmQYBxFtx4IHnQU
lF61Tp5g7n778HMRdndKJ5abnLs6vhBGVpYVap0U4pLFWVGMKcdBmmArbPVf1Ore
OkJ0m4a1o4aPg1oiTZbOG8Qy3RJLnjrkzOhCyhFg/YdQMhzlmFGHRqS81nwYSuR6
NP0yFDY/p7t2YIX4A0vZETkt/LE3SvaYbkzmNI29llzs2Rb04Zqj4zSG+GDzeu1h
J/Qd38QdDaRd+vAxeIK6v/lEP3sBNmdZWJ7hRGUwUOcg5mnGvNH/ThWe7klgMJLm
oH91RaurR64t6+lOVGDz8H7ijp1sGcYsomDeA1SjorPelyhG73fc7ZwiAL/3soNN
acoUTBtCLJAbQz8Y6j7equU0aOzQT82iBk6iFDZ6kML4oHFgHAE21j6fAvueK9HA
OM/oBFmSrqQPBV+69XFh7/kvlAz07C6Yoh8KJkI0J58xmCyP20LBEl0ggTrRxpHR
aEv9JD3e7cPwYz1dmUYYHr4sIfDHjja4nqJghW0B8l599I30JnQBSyT38cqx5YLd
GZgKQdUTSkMF7GDGbdB1Z90rfhOMdFim5KJyWTqz53QjA8bypROYer3tK9rFgH2x
/uR/ed0L3o8vEP/74RZx+XylQPt5+dNFgAnS/el2oxaCCYng7+nvDdQBS2nPyGAD
+6N0J4SsLooxTzU+zy+0xnU499OMtwR8fJ6OPSaspO1q57NC+kRbkJQwivqaYq0n
+KZ4LQCvqsg84aTBsXe5z4cx+DBjJELiiBAWH3csJPzN4KMTXNIx6Vggk/B1xyR8
xiDwMZGjYQHXWQgqHgLRVJZNvE6eAxvtlD9HQPQD8xrpwXZVX4sWannK338osDTV
Euqcw/I/LaCktmmxfQg3cjHQRQTYyGPbBZshBdH5uYGoQnvb6x9XSzuIRz9uf22B
tSLz7wNLCFPmYLZ9F5oZcbnvGICXrsy16lyMy7X2cdZlilURDT8wPZkoavZI8i7Q
LQCP9ujJPov1tLEgiP6m316WBqQhvKCAIgbKkKJeAQNC6kUViNs+jtSHYBctUSzT
jQZAnImN6+kOrkmZQ2ffA9JARwHGHEibaFRnmtE7nvCnoW3/Mf42bP6pa0jj9DQ7
UajdUmAHGGLZjuzDLHDLLCG2Y9TGo/ccyKQETWhHoca5EiMlvrlch3cDSdF+lyjy
ChY2xkV72Lrer6JHQKWtVHH7avekuVJP0GP08cFksyTTyDE7wVoAXuDIe2KeKlc2
RqcYktNwUe4jRp6ep6IG8qoIjH9XkkavEHCP8JldBoNGOMl0gDnQMNcx5EpNpazq
DA85DVIRZ6EpQ50Fted/eXkn7aqQoBPHBkO9HEggPLoxX5cJ22nspewwFKxdkTmH
a7pCbIFdEHKjLbUdwhLxS8N6oABjSzlVYh1hrZMcgn5wb1RXe3hvy1P8vqckRuUh
0tD9M6Q+66ynhvg7L21LUOmUXIZgxIFn4IqWagD7nTio6T173zxCAas3/1XfKl21
RxzFsgXNCD+TditkBTyMH8ZVszPw7ryAmwJFnPEL1u9SXyutz5VVE6d6OuVoJQ6F
Iwr13/8wTYgMj98QgsGTv7xux9bZ8MczTzp/iyQkmQXV4XfnRtAHHu5xE8NzAw+y
TNNNDxElguwRdw6fEXG0oqpJhwZL6DT8icUV7Qw0vraHj8v8DYcpG1rWoG09fTkV
+gl2ekIA/Dki8u50005f3AP0n+G7wOtfpOiN9qrEJzOt5XRs3ModaIwdI7az3xIe
bYvWI8XxTKwHC/w4aMsz26ePDjD8accGgUrM2BYAtVCUa0iasT8H/etAQ2hJVfs3
8ZCHbSTowakvgF9kdLkugzMq0D4ySmY9PcfoGZsWXv79sYM6UIl1DzT8hZ+M4knA
WLHiDxffV6Lyu6jUu55s6uxecdRwcYxJ+Ot2SvOtGyZX8voxt5+v+tU8ASlI7xSY
FVtLZWyEuXLjPNgjaokacsGAr6dMo1t6sg2HSsU9ar/X8uy5weTbnRZieR94cqfL
cgnlfQxoqp0G21RDKY1V/rukAe2bxSKpuSPs25UMek/zwdNTSFoeh7ia0IjjDwOO
ShB8sIjuZkbKViZf19SZJ64ddqCDOWZdBW3GnaU5yKrP1+XGuebsknh8GFpHKdhW
/qBF4T50jvLQ9fGcXYbrzy8ndHrapt9KZbcTvP4b8mx1c5JfuLIThj7yw/VDiOn8
piuwe7S2En3XAbepKBU8iHwmjWc1SQhjytOLr5lgp94pM+1iVb1id+47hZPKh+XY
dCTL0KWZUCQTHwQ1XxGO3m9YYBzxE4nBLf0AC3ZSxl9ThYq1vdij06rzFuHoSLDE
OVmb1O0V1fplDlWWB+z4yIg9ehVc5WZSdn3g/38XQMg6LNkOXPmwxFJSTRTjR5Ca
6XmRr4TkJ/8fBr59PL6WsbZvZRkrO3QzAXHXx7QrxD4+BTqHUIqrrcne1GmEKUFL
i3TRu0Q2P6Hvz/zfiNZkPXLTxgGmDLNAkasNPThTYmcdzvcrQ20w7pC0rGnnawXQ
ounHuzSQxAZKsY5gBDgMWasTnydF2OHbOdVKAnmK7d15Hv2sphLevc+ZG6LDLgq8
W75+M33Paj/dCa9ABbnck8nrw6R1hrTEQO+JX/ILH0poUIDoXdBeTfA5Q1iAXFEx
kKQZhRrIQX2CT5JKfcYEkzYq8A5zKhbnsF/7gQupVf00PNFRvl31sSMYNjEX0bwg
hNj9ZJVs60wUEvCtL2ER5Nc0GmyMLH1x7FBfKJU67suMZU8BdCiiozvvTqGUSZFr
vFIEr4pQdox4V51KrmR2ct4Ufj01SiY134gXtvAO2GilLgF+8sIlT0o3+n/hnnTa
wdsvbBnMX86515vivGAnnfTJ8w8BQmUlOtUfq04fly+QQMHEHyMYZ639lNhrFtTL
AdbraEJYJq/RtfSjeJhtlypGX2OeIM8B50cXH/K3n/1wN6QzOE0i9eUOAyGhTNUC
H6ivdRBHtNWLz/Ue5FeCgyGEZZWXbshnuPdvbd64RGLI5qT/eOAQTeEIpeLTmVT+
40iyeZOHlqq/7ZIGjFF1Xy0IFV9ksit5XauFhcEydqBi6ubiyk3jOD0Nfx+b6m4F
/6Df2Ap0ewsukEb51LK8mL0n3rGATxFYFZgEXAkbtum9HIMpu7HQpIK+b1P5DX4Q
xeS0/3MMA3twaE4qIQxkPdPL3q07QkzoSuz7M8VW7kDYnUyIPEClNGnWLPHGgWpf
3NRkx/TiNgzqxrOZWIjX1+4JQ8Ds5wP2BinAGEUKuwwb2djlPWJZBOEkNzQzUpLg
PDXSOpKnbxRwxVH4KRxEy0dNYR8BkjWZffjRqGW4s9LSADVrSRXcja4XBOGvdA3T
LcfJsEABjTr32eN60IeKzWKtAuoCQwJFpOSFVlgGK2//yVZ65A5rA1FbupmHeoC1
dIJWt6eriSagmknR2mTMu+uK/KvJy5avt9FKbkaNHkNKz2RGmfIROeBihrDkoHF3
4cbrY4kE5OgmbJgnPEVN8poPA8Sijux+NOXAQhoZKuSZz5ClnCrmEoSfxz3PKnnP
ingS7Ln2fEBo1zBUzj0bZ8U7u0TCZNjDVdiGr0ciNMkBpn/SZdNdtgrxHcCqum0l
jpUqjWiVdJjuE+kHv71nmYYnUjp8anb+WdALFGHzc172xzBjbFhhlPL3Fd6RU1Ty
LwRyrnoYTP1UvczUN4548U1zJZm1enbJo1aZwjLRCaGAUe9RGz3TYRYkZcNpQS9s
tG+fR6gzVdRrwXqgo23aimKFgjSq01guqpD5vlJM1Rj8Xs3sGdFcs5ygX1DaTLS/
xJKnhhBJ7CSIz5o1J49/5gzJfRJBm1pTsY874gpJxhXv4yMJ9/WvVtIbT51yc44A
D3z1xYrb0hQMAg/9WjTOIXrykcqlnC3GHBxnN/0Oqzf15M/6yBl3IAy7oeteQ+zK
1GjSR+KHonxUk12ReMzvateOsBrVGNU5x3U3i7MIAobp07rzlUn2EFyS3IOiH4hA
xbHzMAL8nrshBkr0vRkkHU+h0cRpuAT5RT0VezYw6j9XVxKGALy4omb/QH4Nmf10
ixmyN69PwGNvjbdzafU/qaYh3JULAdVxGD09/S2vLlisK2a7ZfvonQvcT+aY76uF
s+DR8x1zXBKlbesQWC/FzU12Phm7D0LNiQrBg3IkbKHCjubgbTlxSt6W/7Rn71ZF
v6EaH+dizvIfH1wxDwmDFVrAcQJET/l5gz2k0DhphcB/xT4U1dkG+I6f3LQIbpkn
8rvYP/J88oJs5+rY/dC/pQCAMYkxAKdQYkjrPAgFZjI+1ug2XnuMDu4LCwWGs7sr
1D0zAbz59TQXKJEmMhEtye7GHG68SoAYTMBeyCrbtA6IxIOz2cc5+nm3ODOjH2px
a3G/YJYwlv4wAd0uW4zDKwkyg9r8tdOK8zKSxwUjYeRIBwmOdi+OjDYL15X4QB7J
WLYJkrqonheaUKDKh84JZNgjC2V9VY6XkcntLTrJ4iAi7SlONqlrdqf9pQ14Wdch
esT35O2b651VU/sgz5TyNxZcV6EZPEF1SdR1mG7mc5cwFCCrFB8WCyWiCwIVI8HS
bvFe2EPo9aBHntxoTkPvwF8rW/UTCU1h8DSooHm223/CaqdQhdEywe9xxJHOFg8b
tWT0njRuzns2LsLHc2IhEd9VxFV8TFiF4GGtmrbBWB992fjEfnKNvsBPgYD+UbOM
Vu35iM1gRe8PB8l03yWj48aUXzlC2sZTGMJpYNp91jcBzjXxFpyXwLjVbz8ui7Dc
bp3hVvMLxjmxJQa9wjSpnQ+iwDL4kuLXB65R/tfwoJ5yoGqnF4NG8/KF76Ev3vGP
o00QdhU65AWmLJmQB2ICHAb+vMSftc9F1ptCNevLA3XAgggUdWd98COWmh9GTHau
BUb+34EVaTJcCm9MR+1iUuBZC4vXF6wqSlXOvX0jI7ZS/GzEcqYsIVgQ8KUkutLE
4YmE9PWOUXLFfB/qNmu2bPL4VDAsJ5w3Q6sWgTKUHwuKjoVlfirGV7svGzeGEwO6
i0D27eazCgLe582NXDf8P/TnjOI0RRAl3v1xIlA+G+FAhJ+irczI/H24mcQi/ikO
0YNpaJhndv1i8muvRKE5OksuLSyQ4+oRqRCUmjAZuj3iBgcceJbjCdYHlUR33H6a
SIGoHjflfxvrrVGLdedk+rFUwKInt7qoMkSk9AtFD0fTgKxMGAky3ZrjqXWu71dS
Ri926EO4vHB1sihk1Dmslyl4b13tym0EKEjWYpqw4DEd5QklpaXr7Ah/1yqXeAjF
N2OYVmUSkBfImLcIhqFwj4jcCohPtDDi3tAcM9JkCVDMGzsghgABos1orezctOGU
5eHPYJPASIkWQ01KYvqHGfO1iwjgaIV7AOq6hVvaBKK6KUEO/soO6HL9AxiZfVVM
tW1oD0p1svk0EgkJVajZQ8GPeeEYxGsOnjNmNSv2PCUXRWio8DMaZB/heRNYjLsc
j2nswktwFdbhJNfUP2mW/kNdLs6Ks0Ibb9dkVDdI/uRwI8yUQShrHifuzDGCCw+d
40tUIAxbgDCOqz2PhGvkGBCmbBMFIqkBpKlbIGyIjTy7JMsjrHLuvf5JcoLWhMn6
+U/gI42qKZKorMBF8q7cQUU6Og4KtFtIxLbjugPeXZUjwayHA5SfN4uWKoy/ZoEH
6if9Xnqekg54+kuw4gmZwLIapb4VfrlgljTL8PPi9c7v22j9vX8UL4+2PdpyWeGG
n6vP1UPv3QKWqxebBhHxj4XvLEXVAVuTuuQBw6kTbqbVLRvPphD88WvcCWWWIJCZ
CgVDYSji0W2UgftN3dQC6JkEOFAIt9oVYYcA8CF1Vw5BOhBS7IE0CeCPDO+7X3y1
x+WAAFW0UUmWyqkfOKeA/L0oqrLotZjqz/JQhzJEKTulpdx3r09fxXC5xChTRZg+
kuXCuW8pQmeqAAigVQkgML4fu24PXRWSjnySxXjIYbrvInqm0XYHKiJCdMb+ilu/
GeAuq4F75KfQBgu3CT7BBgEJl5SfB4527vqr+rFSMj30VFVNcjQLao+mh1eQkGiq
vG8iZX8SR81x033QO6BVAJ22kKKmeG2wilCodB6mdztnkWAwUJhNKY2BevZdueja
Okn/jdBNfLoYPhjS8BKf6Tklnrsmd2o9YripUMaLmCnrqoZcy4mX1LbMXHrzkQm9
CKEvcIbBSKrZKLVk8KZv7k3gAgYpkzUvhJ14EJUXRojymJFd8kAUQOjWIPlw443k
xXv27NqJX+oYbnFWPtHj0ol0Tjm+Dmx58C1hSule3KAOy2JbKZ6St5A8L9zgFPNv
5qQKNQ4Ngx914vzhPoPNE1CYjIIhqRgob2FT5RbUXl4R8ECe/InifygKgXK/gOp2
V0gNtyawrVmM1FF43k1IGCVDiOFfqj8okICL0E7eZDDn0BG+ZANP/Mots2njbws9
r+gj1g8/gK1fukL/0L0jSq2cGztzHRB4YtGHq7b+B4wx8cLGaTOoA3FIJQbC3sCg
k5fl1PKJkIUhcIHzo0WSzeXq8u897XMU2QGhC4wNWWJctcEtMdeQdXxQPzdiLVnj
YvcmYIAZ7dwdrgha1kpT+95aqfq4WmOz0B+aYjq9rX9ztAz4kYrOOCNT707RS2uM
JF3ooUP3RYNevklPWC4QwbYADc2pHX8QOOT+4pKY8ZTXi9Ud3kaIsumMvsMAFthu
mTt0gYjqnleILQ/VXsyVO6aSou4VFwyY+XObVj1RYTFlUHYPaNqyEi0P18JdDDYi
fHlM1oQ96qVd+zZo6Ajo53L8U/qSO/JSsU8HvzhH2oEkCuv1tcUX0mh5FLIKqtcV
yWCabL3hEU5JWFRMOxnwT09uce0F4DTy5pNfVG4EU8RvJLuZ6QuFaHGKNKnj4yoK
biBWGsk4twGHpYNPhmfux1aT7HV8AuusKMV+Hz4R2Hs3mlwqyn7HU2wH/BIxaH4O
8W5C646RZNMGg93UkXgT3bBk5Q5mghigkrwIDFIezk/ccLU+eazXxIm+rs3m79Pp
2aHVHFMRutVNlfFaqGX8QLTaSfl25nuPMl0ioeR3SJK1QwU2mCA1y4nojUQ5qQUp
0FYZK2joWItmxWVBJ84iE6MlOG2FN2b073047IU0j4atRjNEFCFeGKfoBetwzND4
8xSKcz+SU1wsIOePDMzWCHin4VPwwiptOL2bhYTBUeHUX6qGXiOqmHDddAWDlvYi
5F90poVJxV8/Lu9s30rx8R8aQOHRZNBnDrgPcJMQidQuzr8/2VKejS/VvYvkCTRt
ywN/usHkoU2F7KAJOtEZEp6fAwOqlJAjPAXJVhHiwyK7TXiPuTWo0XMVUyhrNmgU
Mjt4JKNgxUKy1ndrHjpSv9dIBKA0PDHE9z1Xg/RatsfsuF0/QodqIKhMe34ppc1H
bjxZGWns3UwggR7qxa04uSDVw1nPtrBSFw0Cntug7p4fCihjOlo5WYFcHXaWSPFE
xaoD2a+dujfdNGYzbWEjA21qf6VEzeza8jmZc1smG9QdI6wDluhHNKezplnAz5SN
tUn1l9jrgsH3TUfJqYFD5xehi9zlZX9iWPJyaatVod4Hde5bt4pYCpDcOWwtY1IV
Yp+gkhY8t527e8LukLQG84XKJrLRAJVlICxLmDx8GtsbAIYi+jz8dG9ELo6vjHZH
w8TAswoyFk3Vfb7NH7uH7PYfI7bWxzmD0xiz5i9tvgxzLSaT6IKxKWcXsscnQPSM
iXiyo+3uiv9+/S34ZG+HnruP0sf+NT2LBKA3KmtG2DkZHO2EM+LZ3dtBZDFL6jvl
BRYzo3F/L2yvk1HkpL1d7w3BI44zUvyYLZyk+Jup19M8y181ziz2lTAUS9SLki8D
EDeUFmprALZkQuKSXUvaGYfb0qfcsL60uPbMvArN3usfQhZrOU7GEPwyGOV3iFnZ
QIEC0tejtQ1MWokX87yEQKhzqVNl5xsbNi3MfuV3GZWrilqAlAy6JJ/GB31Lj9D6
hLSRI+FANb0uIpPKZpWRvcOKR9W3JbZZkZP2urbPzpzFSyWLVBkPQgu+I3FhNOEz
Lx5pfhpOTHM91+YWPsykwYxp5V7CgpLDL3n9JSanrbpHTYqEbCiUFCvTEGMBdECZ
85FnhABJxi+1zOyM/IKfipWF5QZ3/opbY0CUxtxpfyeD+nb3cr5EWrb5moqS92tR
r9wTfYsp0kugwjOiJ2dlJmzf4H4PFxD34zQVKS7YDwA9MjX28t/df3ojGq2cYMfR
K+lmE7Q3C50uHLpKHNbe+9DNdRqtK938QoY6tydmBQfxPh592f0y2E3yN6iIsQ/L
nw5MF2QNEw7PfcDYtVUD2yonERSDZ4kKGoKCB09f3b4vwgmRFBu8DsFjcvo+Xdiw
j/OwxRp7DudVl4Fyt+gZeHKuApzUihUg3YTQrkSsNsZZ6IFq2iCgGLKqndBkdrzw
Ii/oLFp/R5mz/GWDQgORf3icHW/EEYX7DXpHZZnk1YkR4sAC2ckPGuHmcTHw2pCM
JpPQ+VJ6IbaMQnDdXzjrExlKrRwJbAzqF70B4TP+6A5rQh3jQOFV4h/quCRayq16
40rCJmXkbHgtr2d02j9EKr+xvvUtvCXQr4aem08l+nb0wLWnkJ6nGSVL3JLX2WiU
OJhb/dlfoBILLRd3Utl8wsxaCQuuZ6ov4tZ7Yltd5L/6WGmjLOO+OB/JrBxTBt3f
WO1MjRtLM3hXwf8NZdrBBY7+dp3Sk9yane4YA1d5kzIduzadDjdlZHd7rdViM1KW
+tBgLhxdJLmuRAbxHQT+HXQ7L5xI3IYrGpG5xc0prBUifZHGDEnnOxHWSqvWZRAI
0JLgrJ4b1oTCKAtuNIOHPX5mn2HPaSJEsGQ7sIAYUDMi6otJcJZL1DCFZ3TwrMTL
33JqL/DpqxJvWP5oL141dp7bSgcYD6PsLJCCCbZdm0MdHiKolulWyt91B5XQh5lb
7FQqU72bF6LlNbPlUwWY1nJPF3/8sLwqP+e3yAnpz8bTJBCXIDP0mn/wWr/nqogI
BBxnUPoMZCz0Hpe3v/pMC+eS6e5lM2EWqWt54oaGymdPvHLmVdRaV59RCnAWtvQV
e8OGNZ7iPqS82tsyZjZvPeK1TqH+ysYQyH3/FcZ/+Tbf+RZmWqM48Bh+vf4n03D5
9u9SL17X5RJI6YtRPz/tmhj29miQCO9kTyafC/GP9fXbPejZTVKs+KzhSLHz0e10
xkEBZq39heMUWp4WK9POtpNYUo7euosiffjLv8uTNnPUSioE2DfGmif/v28Kv4ED
czO4QbqZhZ/XP2o5kUfWpdOEiRXzHnaD+5oSMdDADv55TK/uks/5TAgHurMqk9z6
yy25C1DW68IANtK26fV8YSvsJdCM4DDtlIq7HLPoveSmQpYO8zVcw18xEgzntyxZ
xzLuspY3HWdX+rqJ0cLaEUmiUtMm7tHdCnQLtU5Nw6jw+bqAV3OvdDqQfcRFZtKt
yiBal3N5uTmK3xGkwF/akGZ12exAzOOwvYcJw1NjyQ6IEQXY9n2AK1jmMe2TkTUL
D1lZDSjtm7Da/JoEtzL0vdDF5EwHLSijUn9gvgPO9RRhhFxQEttM9da0FLas/uYA
vHWeGMJGOKuvTPhT+lNs8k8FeqzdgYLS2JrxAtVyMGYQ6+6B6Vu05aRPJNCiDpEi
oZaT/flIw8MORdr+UU7c87akA66jBeQ6vlkodvf2WgoQXCxW0FSvkmv/rwAcYtdF
zu7o790Tql+drHVfKsazI7YWL5enMm+Tx78Pa5R+n9D44CIDclEvGjYzzh7kg5Nv
Wrl4KzleZKyctHaEqcGBQR++c52QQ/GdV17XoaNj6cxS0r8YdJU0aGA93UrMCYwh
nYVoNQ0PXv0le8eIvYLM3Ad70cdBI6xnvzMdBs7DGHsmFqZnpk6qfG2RPTIkBBzs
JZKQsdW13D9J9cN9du52orNCerD4nZUPwkNmtMVUa+Il4P11saeZZH8lA3C0jzCL
uOs62W4xJkxW/Vk5Z9GnMgMvsbZxzkk6wc2YdbFRK/C24vXZEOVgys3dT98Z0z1V
h2E2+LLz5GgYFODJEg7mm4bIW7M+y/u5odmLINgd1LM59D4afFY/3A7yyrL9NO9v
sN1ja9z9Czf/v71FqhtDIiVGKprjZeOuEHTA50SLzukqFBmifOZTF+WmZIw47qR9
zNe1ptyiRzZV00yNUACNFFVgGQH1zk1AKZmkCFUOeG8osqoxmeO0nu7tZCMXAAmH
oeP1DkrndAY8OGq7Orf8E/kCdSVyMKSU0kbopmhLhRdzwQepH4CAo8nqgufv2ctY
g1PU/gLd1unuveegwDb8SWNCIRkTmkHG8t1Xu0xTHLfgojIrSvYdaWTuH2eUOAF5
REkhgkrVie+wXcZotEyIGn7Cey6k5BO096Sm3sWpId1QNyvEgWUcOCgW35Ke9xbu
sr6LvBft0rEd+kCjKMldhi//DjtnyYzzjPfbWuNnhPszaC6Zv2L5ZScGwR1DqlCp
lEHthqseSSFHqVZdcnJ5JGJMF00CHt8G2jTXL8e+yJej1hShXdINvpxI9QdLZdj0
x5hr0SxoHD3ph+g+KNIAYBRLdZeU/jTgCqigshe4el5PvoUahQzWO3I7wLZfq1X9
T/wPvRfajUb0IvD2RSBRQGZjtqQJDm+kygY1GaNuMINS2Ik5q3lcracHSOQ1a5ek
e6SDmXmsm9iglESw9BjTECykmly+MOvnshHJL9NuC6Syn+a9uzph6Szy3j86gKIX
ltUqasn2z9gl74iHcBJZOCd/rjIrJuXXlF1ozAUjAbz1Lo50d+auJgIINsYnBelv
DnW0jkonZLIzpn2HUiMu3WmLfwQjbMgtzMhUwLz3gIKc6eFeyW/+3/hkAWC84m8N
enRGiR9xKkHYUXcqgVXF1jMrGODCJksx4VwOLyKrhcWrToksmD3P57JFOolRzeAe
/8CSRN800fGRReEe06aq3GkBQonJ7lZem05H3VQUmCXoFZjnEzgVjhGHSmozTQ2X
fkE1QGA9GRuTIaVnochA16Myc4/1uIkFMhvTHAi7Hwh6Dviujc8f5VTsOURV0sm/
llBi/jdlhAOt+1T0mTLTCu6KdN6uTs9cwx7Ruf4VOPSx4LsiHmTKPOsJydU7RWnz
oZ31GmmP+a8uZoJrxzcgLsBIGO1JIHmGRjSIcVd/7QpByFRXOXwB1ofNJYKeAZdO
WvhM9G6ET4VXma6Ao4FbtBVNu+l0050SuVB0sz4ksVnZOmaYm9HirFqx3cWSLG0m
RL6zS4gNXlSE8Jk3xZ+5wfem843bHV1IO+fBGmr011Vuzjd11UrQzwxjjo3PsI4N
i9CiXZ9D08dCvDo8g1eAE27TMLm68h6vFAzWeeJmB6diLo9M+A9/61FSWt3Fs6Dz
ey42R6GtkOI97dzqQNSqEGOy2yIKtDMuP0P6St49ioRpyuGXFMB50Teq2CjSzTA9
t/OVjrdsB+ks6EtZGm/8i9VuLUhYPIKtX5gm5q7TIP30y5t7mmn8YGbShBgLEXWV
78Sf2cPYk1JpcHJFsMZEe7f+YW7PQWHjT3WrPZzTiO1TmjdDVtCmRSI31LbVhykk
/bKgnDBg3P+yzY5rRBpN+adnE7N1u5QzybB84SDPF+4PTMowNhcdKYfvZMImxw3T
poSjQJXUejLP88gL2IguqWQKVbmQPTAEMPWRHZkrRQUYgaodZH8xTiK5NWa4fbmt
YVSD+3YtrCeVxt8LUFQMVEM4OrLEoWyI9fQXXvoMuh4r8wa5MbEU6a1WGid1K64J
WE/TJkD41uSfCSw3JCrTRYBxZoXNDQ3W24MTqrtnR249tFDPjfjA2KSa8YBoQdrV
6an1/tn4dO3VOC801bwj1S7rNNvBpmBbpj9Lpp87fxihiLvvdNw7GWX90TLjQ4Fw
H8/JVTrEVwxV30KQ9u3avWIrdo8kPP0P1Pj7/CoOwPVJX5boOBOiI2s50I/Tk0W9
6ZMk3KmlHBgpifZq6jzMa4beoVNPDFYaURpUchgS0QsxcBXABhghmOFMJTJzy4QA
Qqyhtl0QNewfzv89M5C6toXMg0LO2HgeDlDf2LmnA+Kougcxkj12JBbWmerRfEaq
Behy2Fd4mt6DU2PPKP/+yiFgbwgrAzEDu4xBCbLWOq98LANVwIkQ+b2ZuEGL0S8j
hUV408F0IkDcym/KaRTnNdaECT2O1guI0TmZmP9q/TJqk27kYh+HORJ929NndN31
R35xhl0Htekn+MBK8Mdmf8Tym4qZYnQTbqnVxmoc3xMl2+N2cb3FYt3GLgOo4lGI
d28XaPtGN6Ivf62ntzVBi05jg4ZGNIGOyLs63dWUy1QR9ktrzvsZZN4QwJfT8Xx9
/g0k/vfHH6MJSu9ZTomrbJY8wxRFE4M1ot5AxWxBVNUFV07B05wU1XmF/aHZVOY+
okddzmbvwnNNmUwPMb+lFP0ANMsfIsE1uJ1SPAc/OhSAi9D8/xsti7N913L79iLg
OffGtCWK6HgOInpxmM4sPM0XJg5j1U1jkk2M09kbTBVEUW1HYlUFw/CPOAVjeLti
nF6uAmDT+Wz6ADo+k3M3R6MjZG9hJNpoaNAztWTRDau+Dju1478t69AAutGYWFrx
QMywh8mFQ3JxSxytTk9fg3MTUYP25Iogrvk5sqfWKcrbgyvGTL4H3hh1pqAnmSB3
5yNh4HesfLOTGS+roiPFaU7s3Aep3waH8cnHRCQ0EkyHueZ8dj56hR3jFiv+UAa6
wYBnLHJ3y3VL2x7Jz5kyzHE6wRi/+XIF3ecQ3dFR/mlVJ438wfGhimiNU8b78M3v
mmimNG0wu4mwGlG3Yi+z8FaklT3y9Wj5x9+5THexTo3XD6gDhieIC8JKeED/W9/I
Pf0nRZUHH2nBtkt6TberVIr1fPXAqRPdNmAH5jKAkiUfyatZqnM3HzYELXfFUmd1
LHayeU/DuIXFZetGpHCl9JtLW9LvFcBt2nz9cgeCOTmMxti7d5cPaELgpetwcoOV
2qWd0MVrSUZS1yY+m8wrhiZH81Ov67IG6qOWUTAWyzIQNFGimpoV4q7P05HrZ1wn
QH6RHtekW8B81v89hctj5foex7oPXq4ZGp0s/SIpwm81N2fakFjrRoHA5zl1fxYQ
XJi3sGaX310Ust558FhMqACUL00u3eb+eo704uiqQLmbl0g73bN7jDl2zzAUrzVb
cnrXUFz34bpdTaHBerLsmxsvc7IjxinNao+7J79pNW+LUV6CF4VdAeExv9KMO70c
5dm/V21BhSR2vCVsSxjp6AOF3uvmGgyGvFnaaFa/Pz+h4zeaxlLcvUK0MzxcKxsi
UH7Dn3RQTCWd6p8Tj7xfwN+EBltIcQyqGd1KP8JzWxq8duXrAs/jHt3H99DbpK92
cwTY5QQfoOF9aBuVKP6TSfm9paL6vF94RHvI8Ht7A4+8zWJNBjh/cZgyQjDLVHPu
0qdWxYN2QzwxylqgQ34o0AwezzDQz8VbQAcQzwf/m2kX4XzEjH2Tv/JfvHPib57x
OxvbdUURzZUUV6PpfRojD9n2Mo9ibFd9QVPiAKJm/ItNhPL3egYT9+Kei9PkuuBD
2uASLbvKLuhHx5ArpvsIz+7+OU6M2wiq/GFJiMGSHBITExVBLEFQvVVCQFWpRmqO
cPEfZI17dJFYrITC09+QKIXIrFzhQKtmmoDF4aviveZyhf198TpEUBO/FLImMQX3
lHa3HkEF71PfTgt/v3KQsmN4G0X5EAdsnG5BkMI8dybOknQmx0JaT+dargMsEEPJ
asCp2UUXttB4N8gnW9SQseSRAIriujVxFuNPzX6FiIQyAL6GzSc4tJac5JK1M9jy
+Xx5GIg/aeRWVzYtqyNXfklrZ9mSdXt5qtrL9hSc7b0UY87Of8X//spS0Wmb5te2
l2EgCTcfp6/6kln0uCmQIalYbbAMysV2UgVAK1EgPjIy9WLpSB3h+WqRUM1Au8kp
ZxUQITLLY//IUUX3syKJP1I2NgLb3khP2wTu00MxwjkuDYp17PP0pCxqcVbNPTZ7
7wBeEnNBhoJSBQhF/mE0bWCav4DEkvHwCD9jhg0wGeAU38clqufGjnO/1i75KByf
WUabY9yr8OE5DDQdTx8Vtua6X29ASn+SZLvA3EMGs+/EnCilwsXK5dvZUaCtt3Ti
YBAC/6lFJWvE3YASOel2OBbAaYWrV5+ZibP9bP1+L2jBxHfKrrKpKo2/7noJxMVI
efJpDADwivzkWaLu4Dj6Y2xpEoRX06/t62kZgb3wMced5brYXrS7HNYqHhH31XVo
+GEYFQqCoWyMCVvpq6PPhjW2z+5ECWU1MFPpi1U234RR3qIlqhHS25ZtdojASsog
Vnn0/XX34LUlqeipEbArcTPH2D0hduK6L6KP9A2G5mvkZ6lgv3JlIoR8VovKoIH0
l5mabmga9mC9w1jIUG8kPJxldHFyurWvhDexzKxnabb3WwXCcBslUpg6u6K07RxO
aYXnRFfk1tKu19eBHghnXU+xbAuLSh/guPWth4+VfbKkzTFFRFDLVh9yYog5U9fU
zhy2BbReZugUy32LC/5yGQoL334ZKN3ib9HLT8hOP2eQN3EM8FEzUX+jgZW4KQMw
OLI+nku9wjqO+yaTbdLNonB/IIDw6JJgcnwPUptJRRGGzRs++nkEgGxI/kjadQRE
nSX+38XXdaiYSffv2P++TQmva7N4C2eutpbhtF6vgCLhzdnzYkBsnp7OOC1JchN4
OlUX0ZDNQ2Tjs6cA70fXXmApowen0ppa5xsIBUtkrIaQzFPSJpNcr+3eM7eeEm82
SyFj5WJksGa2JgF5UPbY876XLDwsC05h21ZpWYj7wy6677JbVOwkH2fA0f4telJv
E6cCdRPi+C8A16ps1J1TifDmUEzZuejOqkYWT8HjaB6HSfBsu1pWCRrRWtaQNKtZ
jrOIx5hzVDHJCz4YUSllcdH7yyYSrab0K51t/l1rP3TlKN84IVacI5vpZz+gKebB
74naQKGrH5Wiic3Ft4jDfLFQ/Qn+v/++3w/SZhyySRG/5BRttnnSGv3rBBSHz3nA
SeowbSWlGCwVT8YbNHTq9hfw8g25iIiAGdh0EEbu9FYMb4EaEve4Rl+R3G3rjOFn
LoJRGPJbqoUA/GIKUAtMhLw6Z3od+8zzwJQ2Jwnvfv2rz05xcLoZS55/i18ZeUMm
Dn26onbvHwHBsMQG7ygSZ16nIImVqhxO+3Gofx0/wIC8aykHIsHfDkyfCiOMNIRV
/QadpZJIcygtznEhL1aS1wgCXAN76PSfdJsYaGvJMLOGF0nHKib5A3viwwb0dtgW
ducwVhochRXCQWqR25CXI2FLVKWYXZfT6S8VATXWL3hCDNElE9Ve2nnf9IdCQzUs
GgitzkseXuWzjG6J8LtDkkBhrApx5F4ptoDY1i3+ZKmenQwrv1dUwik0vIRNIL8S
zjkV30FjLnS0zeh3quUJcs0B8VyrsJ9D9S9F6zxqrh0C/kcxW/1JE/rD6BPJVaGw
vXzvbGj0kEdMiJ6QGhYp6CWzNb7al0IBgX3bnGP+rNDeVlLsErSR7wgD/Oi8L0rk
vEKIW7MM4dwE6653jSh1FNlMXRcaltDpyRm/aTGuHOCNVzzzdxMVOMDFrTjo0faT
C/87RUA2AOOVg5aKHGjTxuThV1kQNDYhw+Qai1MhCVxY42r+VIXWYI8mxhmuBzHu
w48ova7BJzwdUv2D+u5MJ25P7UWYYHZbXPtrAYMke8CXcdJeZ5oM6g3bLRewYMTe
Nr9AWfusavWWrC3hrcFHBGGps/2LP8jBeC9hvsYgnGgdTu+67Vu5/HJh2+fOCKF/
X5o8dUqg6wbVmoLWQFHQJ/Q0+szMc93jLHqGWSw6XSh/gSakikmcYu1IR2agttHu
tT9neBlqaPt9K+naf5dAG6nBjgdW1FjM/WIxJW3lX0svCjWqPfwDCZb04ldbgPGQ
ZIUxKIPbhnNVfSEejWxbz4+LwyE4J0iMFSTMvcAoJdAmQUKB6/hNAa1H3hJIdAQs
SbLld1LMoBVHjDa1dOkgB2Th2l52YT797K1J+pVq1FFum5r9e1tTI2Am25XKEqRa
gNxwH8MLrzi/WeE52mFcFf2fX8qHnR8aULhQQE9lc+bdpWqMCjclSu4Jil/zoPNX
O1eIDmg0imAwxBZEJdrfws6bPi384ZuNi79GGdk0WJbVl6uJnwVtI9tsd7X2wYA3
UyCiz9AGRsGCfBAgUk45O183hYwWxgojUrThNJPy01eZQelmqqBMXA7EydiGpfXp
hsDaLkUY3MZuas6AcP5Xs5hy8tCvGxk78W2m6Ff0zgVgnaXnx5nTNcF6It4wXpBv
QGEisI+gzCW9mLqi2hiDeSZz+aya9wXAQZ1U/wd1qjlIw9tuQ7h7rHEjSKRzra92
4HcKPfXP6lrOvRvmTCrtnHMcM/l2EPl7qDJ9nVJU4kWy3Qd4BHkcBajul5P4Y3HB
TBPFNWgPjDylhWKAvDBkEdR2ZpXwOawO7yOB2uYUcvnEsNb3pYCNU3RAYUXXdbBX
K+VZIOzbtAhPBN0yoRkQmbNGvWbAO6Z2vakZghFIKWiuPzu/MVKWhCVFRgJhiHbB
Kq96p/+Xf+3FIy/a/bSF7hBqepcWiNdfooZRaDQGEg3ipgvevt0svaN8l0RJ5Y5y
nIIXP7UtaL9MO57n/pfQO/khzvAtuNahlG/rmNup59BOL1+5uJ7tI6RwyLKyiP4e
QyJT8fQ9EjDQPIawUZ3sQ8RXA4pPOxu8wS2hK0Qnh5x7GYbBdCMCgMR9GkC5uBhk
gr3VTFt5iNB50u6ubDDK6L8lKfbaOv+hMUR+Y1dBHpjJ8I43MjSSYRgciSOqU1ms
NCP7IkNDSwSQq9gCtMbsGSJRdSxyBzz+tyCiy1RTAIBu+XPbLcDCeKWGFdnAWkPC
gfwdsR9/W6ZIjt9jhlWkSbtVp9RA+RHw0K8ewF7abKu0+aHVwnH9Kqw2HdY24ror
MhW4AQRe8D0/Hz+P9NevWX1OOoLsLjy2GdTmGgsSV4tJsvYoBmMEkw577OF5Yao2
Fq7xz7/oofYJ9GgOHTghjscGndnEtQEDuEpGYINbmoLNBryfjr+FOtkHhPhHJWaz
jQZhg081eShIcDQS5pbLuQPLMlqhJcQckMsj/y+95zC3IVlAgONS2Wl7fFec9Af3
Rt/1/TwkgljYmk+5U0ezKHPr9ngQO4rzXdY0Lr5cHcN69e/xAAqs3X71P/NtYvSM
hYfai4UNSKfHZGJDZD0Xw4/9lk6LUS48N339oJ/F047yT8Sd+CBTty7sIHt13kbt
OVvS3E6hFA3PHWj+38yA/Zw728Cy47fg0rzO0pR9+oJaeQjE70RnlNnOW3nafASY
zn9b/aKXEqXtTsqU4j/+axI/AoNk5yO9ZOQ9oG6Y+dSulGIo7FW284ZHBkZJrSm4
PrZlRMov5XgJkYStS+J+erdyuLium7hFJBGHMLeliBE0MNP93WOjIrmjyQDZpo+S
vZFceQOlISxqTMncZ5YdmNjOahlqf32s9zJrIv76WIMAgyNAsYiFi8JDppjNfOXm
+6IiDQDO0iggOwXynjD6iGbA0TicXvG9wwHPnRzmNAeEv1hSg23atNTC7/1c78a3
/WtYhnC7VYHZB3sXSGeQfm3QO0LcJB2ISce8uVc0+qnPqXJNUJU81eEFPSdmnHCA
N3xHPuk5WheMH4g4U+Ac9j6a+uk4RGbrqB4yTmOFaLFJNANQoaSGxJj/rsvuO9oA
BroQ+H/RLlLTP9R31mQb6sCtLM89JkMTlyWPcjL1n+ePpcEV9w6yObcaX/bCMn0F
gxRdUx9/+ykVUoiFbG7Nzad6mLzdPtRSvcN/J65aDojAOADyXFn/UyabptC/mCOq
C9Pmgldp4Ej/j3SdivbL+9GHFTtLNc1o7Ia6F5cEqtdsT7E9n5lFktGedqyyMjS7
EKDI7dXhmJbbchJFaO2ANWogaJIeVLcrIEl5/FYbUrurVLNXDKVy4rSRarnDOCk4
6HvGmqX2qg9Nh+1eqx9BEkzNRXbEM6ZTIF8/3YxG6/UHLIiJ8JSaRUAABCZH3Kmc
djBwIGBWV7n5QIcJDoq2ie6EN1tInnSHW59yKyIN1eaelzhI9ZdtYP+dwJQbqLP6
uhMTqt1kSV9oy51B+itJcvgACsSe2Rr2P9JGv7Vqw5aORu49wBfxGlyodnIC9rWI
QF9fIS68hkUNyS8yEsFX92OR0+9XGY7d9BRmQA0mqptyrFwbBlg8Zzr/j3zAOrQU
1TgfSmYUsKxxAdNp8DDECBXRzO3qstDLcoaOZ/vKhKSuZDRJEqDnAKvhodckEYuI
+k4elxAZzS9o53VJ5/R52qeJuXvxjd4TvBvtJDrXdCYGNNQy5oLTCFtCsSMxZgaV
YqKzfWGvqhfYpRMu8fGgztZnM8TdqfnMA5kY2nHtVIG0ZRtWjXJXHq/FG4weKXJ+
9jdLrRz2eLY/o9Onu/9Sh7AQfEt4tfOcWHot2hcb8mKmX7EfyxIwdwBTwxhYEWH3
kPOtsHBh2YAmaVi8YBIfy6tEiUNE8vTC+XUFjZGEYKzHNqGqcT/0iKVXJ7RLngDG
YpSQcTpXO+4YdYODVaKtCnaoYAveypmkeGX69/Ho0tyhq1r3el3sDS8JRMb2nd6f
ZzDGJph/kha747kiQ5+uRjX4tezW53qiweIE1+d35K3CTzE27yPKVP8LCoqKam8r
vzBaws2D7UetUDfZwgYLt6iVVn71hDeivFmBFfrxSVKYC9olETthKzEpu4IYViHZ
KTUQCv5fjmjpp6VF+/6mBHZBg2YhVSIlVWcTWv2HZ1ZDktyPZ9yw91yeSDd7Nw/8
mxSPm4abweLIBwhPe8QVWHWyCyYV2rZ/T1xlacWlhlvkAA4v1qgqlW9NtS1xyQyA
mnnn/nm2vDeeTIIxVJpKU2Ilbouvw5gU28xbzCvL97jzQLAjHKjr7u7HFQ71s/4B
E+zf5ntCsNIWJ28EU58qY3H79qfaIbojEtgnS8Ff0w85Iw/QgJsxcTRZy5L25vv7
zYUvGeii+7ZAZbrxupMv4SVvI16zjUpS+gr5LpEuwm5vxrhn949PdE0V/qinqvS+
AQjoEsVNxSTrBUJe0g63LRewAlud1l3IgJuTEA7hIxbA0DQc0RMdOo5DRhVJTEJb
Ks7DC6+/cN8Hf39/gVgQhmywoXSm3yiNwY7JMBoyFv/fzB2HcsKUdPOcB7nHvYCo
RP9TK/VQ4vFrGtF0WPGuRmXHb4vEssk+d3EMd34NAM8qA9xCr2hOphVvl/ZMUduY
TCj+emuXbtpuWiuHmwtASr3Xy2CwkXBtXXrw6Bo/cJFNgk/aoPB6U/gHZQYfLKfK
gzhQwUub8L5z3kTVkm/L+gRiBvXpCof/Ufxp6Wkkr7iR74WRcmjWvWelJsYfTdnf
rVKSeCsaeeJ/w/lBviTRA+cXUOxCyU0e/HD0zHyuJQUn7OidJhwEr2RdKk/u9Uu4
BmxYKTBEF8dQEq1RB4YhQn8/Ds4D3rgiBWCvUSI1kyotDls0km378xsDBLVRjA7f
yAoDbDH0QFl4sqX3lTGv0npQ54OAOEv350Wbur/QQQitwieM7ej+ncs9S2Qc0TDf
W3TReVTOaMDSJ/jpRLxZEtw1jGBDtau52tZTw8HKzcDgQyju9VjYwuXn4BIhZn2q
l1DxZzhK9UfvK8rzD7nP8sMC5sJHua9bIpxll2NOI8GE4YeVY28H+xorVYtwYc5w
cgG8jJvBvnkomTjRPzuOtwrdgPjaT2kXvrB9pyeu3Bzuf2SmhJ1KZbiEvGXuriDL
Jac+N021wLVMJTFmw1PuDdmbHDH/B56BNF8zZTUiltsGXTZBP8kJRD4x9HnT998Y
PIXvw2cL+MiGQmgWSR90k7Zn01JmUZ+H2kn+yOW2btjju6UsY+jjVDvkYeLGpQAG
5PAvE+oKLEJaDIjf1Hf9ycK7Qsm9xNmlr7//fFKTM2QTlFZGjFKyEoe1Uquxu6mC
7hn4u6HbCVl6UghZcjddUpDpUxOdyAnOC/yHkY+a3BWtJ5y2FJtUeyK2fj1o4FQn
PWBv8rqB7OwBzfd1oS1RsFs0/XOGZmMeoXhlBpOTIXWZ2PMv52o73eGNwy9phTB5
qjGxY7JXmhhi2Q5U3izsS/3QJAQ6BvRDPPCXee5RPFnCTsdiGA7unmqD58eUR5vv
YCimEYad41CgExsFms1MSlE2iRt7+dAFneD2/+3Cw53etqDHCiaaeVU2cgUsdl8n
XpVMjyXOAUfxzeU8GtIomHia3HJdo1ZZwmiuB8U+4HUx2qHcnjmTdiVk4/Dcyqja
59S5Yv37eBj+oDxXoCv/ZjBMExXbPU91LMbVakEI89vRz2DTtJxFw1o2TGeCrBm2
Tvw921O0FnnUyeJagOYDyPh+Zj6lBAjEkkPNEIY90RsQaoQD8ohvhJ7PBD6v6cdj
jJUrRYfXCYIHUnBCGN9XwUReXGPNeO/C7zVEElxHGfALOgAWBoPABj3TVIXO9ux7
6ZKVjYmC+BUhd1qahjgOlIb+9NGopuI8HyqrhXhOJ9u+v787LRN7q3tDKtCgi5NN
xo7V3npbdtGEvSZ4U8mpnujlDsrSQA4z0zQQPDYKihz5gUDWwhp1cnWuif/0cgkk
4F/9T0FiEakeGyd/1piCJ9lIj4OvFhwTZv2+FXT97NpDzzAxb2w7OGiDTdNDwnGH
vQvFLXCEEgwFmZOmEqeG2rIATUAb0UdaPZZxywcSB98ROywZ8hRTnUUaGIyXLD1B
Mtu7GDIb07xTjW03gVXdy4dMjpqq5NWZFfT/0NOr9Nf+VfI+TlSKTjspsZGdLE5F
2qSRKA5q128BWzGYXn+6tZ4uZ0SHyN8SUij3YiEYZENquD+eQ5hZtsXztqY7TmLP
xNs2C89r+uYsNCJc4eSyTwhksrMIQyN3hlFRKgx4x8Hgxk6K5mbSWxXuasB34vAa
OkIYf1qW33IC1ATuWo8VZu5OIpV1nz4eS0BXzfG85v8krMSt2H6KXOzB/rimLvXA
xVfZqZDLhHisnYXxzn1XxOdEYjDL18B85BkNdWmu9oD8Oyxtrl5hwn1LBU1bl3uY
Acl9oIPdKJQ+tmun5JNcw7+71LOIj67P9pjoV+kczgAt4aDIuoxzXTwDG5M0AtnK
yn/ln3yX8RZPoxQDC4reLd2exHGArttg5WF478BAdRxYXZ9KWspxEzEJ28USKdCY
mexhI0nc8J+N2w5HpI+iwrLjniUlynAF30ipw5J1N1flMwvIQmZ+4OYTuj32pQsh
eMwS67MkI6wbfxhpxIiXSMQKWHwM2XLXczRUNVN8XeMLVBI0Gt1CcJuikxNLzx9G
zKSNfpPtJvYYbH75TxBBWzqVRK5CnmZbKreK+UxpJaZo2W9t1qb0xB/s2FbeWrBN
I5XPD0kPSZXlR0eqrh+V0otLThG7DEKDFswRLUSZOfh7Wv4myir5StbYklAqOxBi
vg3OK46hTkqh+PEiS9qAaImXs+R31+gy9S6svkvkKiLbTwrI2fBuG8Gi+CxoVihc
AbTVQmmQr/XgaB69/Rgy6vDl6LeO1d/wQAOFg4FxqD9/rATHjumEJS+5B+styU2a
grpenkbXzGQEOHX998/67w3p0maHOQICUJzgDwdEl6okLyovgggFnkl+LyMB7pIt
mdTiXSdr14mPl2no6HBQV878LgF9klr/dBEVfZuISp8eW0jjYBN68I+l7KHy+Yib
S4dGgyeSD0xBUOHaWvi04AVPOEKlsGcN77oSx9J5hDGZOVGBWxkQ/bobbD9/rpyH
svK9NHoetngSjWOXdd/3fs/HUnG48zzSCgD7lRp+/wNkdrf2Xqz8yan+xAS55UvH
a1EV8qq/BcoofRp+efImtERteS0ycyF30E4lXi/mUSrFF5OE8m4S4ntJh0V9fYye
bmGMj6NdUaeRMbYYRX9jp0gfpLhvQrT8eJcNjCpLrSnTMKtzTbT6W5S6I+ix7Qnp
JQMl4U48qOl4EYjwv57JY1eEGRx7lID2IFBCpu2nDOSjRj9DNapXc+E/C7vUgMcM
iVjXdY7KMwr3QC8WFY9kMw4r3txOsekKxWttoR9DzIXzNlXs1JC9sPvT+sTNupKx
gtIXiu1beIrsHvP+PVmlxZyFDB8WvsIIsU9eWzaEK39/0eN1uhwgSZp9+Ecxv0q9
i5qs/76Mj7CCj53bKQXG+3N+I2QmM1BQtXoKBWoc+0p3FoF3mFNkvQrM+4hWgbWc
IBo+9plnM6/TXm8VpPhlgKp5PE4vEj1jMDYsMJKsUQf0y5m19IDW04yOhJ69Buwy
kNyiYWEv5bT97DmoPWbrwCFSUPHqa5sxVOp/HSjPJm9brA7b+PkGFKlXaI4J5m8O
e1vbFBtlhQgzttEzWHCIMTJwnf3LTimLVqMoGYOb8PTgESZ0UaohoG5f3t3K1C1C
+C42mGId+jEUXCoJNZBStfIcZIWQALAHBh5eJwjwq09yyxYfWsmtsLEVU18rPGfA
R2ALC9+BVmaQcqEe/ZlzOE8WI8Vd0O8Dk9VuXaLYWlQUTePvWVjHBAXWvzqmUXbh
giOt3X77FmhqgUgBLjlaxg9Yl4Oy7zymcpe6iExWVXtPQyYkoG4wAc0pWIh6eUJU
kn17maW7VxwccDrLmTfKefc5HcwumpOXPxoyJau/Gy4FnDMK/vwlXbO/1QLcCqrY
YqDqULBgt+id86hoaso5LG2oXEIcBnLrzWXcBvwSrgnTA5twDZz287oODmPFtJWJ
uN8erBYQB6o8PAOH+Ov4AwgY2PhYuiw4PuZZvvGIsXHzukzzi0tjxo0eZ75/2PeG
PISYsYZMYMVuHW0LzIHjkRRkDOdFLWBgEEl2wPhmCP6oIugSYzWfstBteIPkeP24
QoL+G7BdThO1Lxr8nrXDiIUvorkn+BZEUZAbakbFRnFKgClZ8uxCI+EfDCl6RQ48
Dua1bidBMnL5DRKxorD5ItX0j+lvBdyYrPM91baYFm5oQpwH/7AriUv6ogw6orHk
IYK/vibt1snSg6bLW/B8W+0uH1MLYEuWzz4iW3fT08uDAgPe6+17uV5TtME+V9AU
SS00lubYNIIFO/s+o5u4OByA0vQoLbLw5/Sec5Gr/KkFArz7mQw+T7YVi5I8QxrM
Vag48ekPuXKBzXAt0r7+edIWHbScL2Q0JGDFXtLFPSJxJ7WvFilJYOg+18QtwJ+W
4qbU6LcaiVUhJYzZbv055ZbKC2/l3kJ9CurOYxUatWjn9fCxdfh6fHFBAXBzv3rM
WKVUGWF4Gsfl+rrmloeJDzgaZfufShcTJONrfCPcMxw1vCsiy6fxtYAo8c+J1e1V
JcnwjET3ym61kdaehbo/hN93TdVHVjP+o0/jCQLwKihpwtIAMyurwkaFDwkK29vf
gW6Qoz7360sFwzKsi+fBP0jUl769tSvlo2CFMLLqZxWc3TcTKGKdJmhqQ/dspoYr
Nj78AnLHHEENcWJaL30tFHZ3+6npLQLz+gl1BLwdMFUZ9bMtC6a8FyMbGxWBGYaK
bZ1qlMgfopq5ss54/AlRrcBt4zFSUS9Azgq95frPE2Yd3AqQzUBtsWBruUztig3t
wfSe0JZaE23xw2IG6TeKCR3PHb1X6d1ScV3NotFdU+u+WhkTyIBp2/Az0Z/HWWuP
AVBPizHlOYBXYfQmR/yV1Hzk5KjuoAQLKUT2/z8HAjuj/azGrsvJhqY9hgPLo+5k
LFwmzFHLq66iqbkkCBR3GLquoQmP+OYiDsfDck7ohGPfAjd0UkoGbCghGdayEXna
HDCPnCRXgVm8oIyX3zxMg5zbedZ9yy2JINV9xnhkcGEMG7s4MIuVfZGlQJYWWtgu
djRBKPakJLW6/njq25HRJQSmuwrua0DN8i/d4Kyhc+zcEOUCy1ccKCp7tnGmQQu3
IhDcLX5+RXczD0jAqS4leGX22sh18sIr4mNAnuVQMZ/0MXfemrNKWftW5jZYhLuH
n8rpcGR7VXBeJ8/F3Jk9uUnK3mJG3MprTLJcjxiAEQXMK1mdyz0qJk/OIsTbGFrh
EqJUJ0HcxzacxOA2nacMWaRu8FQBsBm2DI9jZ8IcKqBr+scwoNIgjj/z1Hua5Cvb
Ax0hUjLuzKvgqwqaiaPeOU2vugKVh8yQWUzU8Wj/vQcNkIyKWPjzNmc7HWqypRW1
XQeYYk6X1cK/cLyHtZ2MbgHji9DtLhS5s57JwIW6+1vGaBfefJh8l6yDRMNkrbnI
zgKXFv4LSCyHjGSUpuNlaBVY8eF/m25dFkS3UhqCvTh6fvVpHS2bnYOww/ve1G6T
KOlukH+9UfMJ1FVqUSwTe57KuheJ86svzYrpFzF3IIAQjMQ57cNgtuNPRhfJREnQ
JB0c1nsSSDA+UXOzsnYTgtxDjxaUq9t+5M7bR0tbEd9zOhwdunFmIengWm+LhLUH
ZIl2e5uzpf4L2HSVRu7+Ubo88rRN5XVtB5i39POFg6d0i29QVVQCyLwc8bhNglPB
NfxGCQlUdw/Yd1EhbWVxlRIIORuQyoPaSdmUGLXx7xdHaR59WjIOEF842x+GLGH1
EdHJdPuz0tsLqUaiyduVWGxDUA/LkQKTydO/9LNQ7S/rVMxvQ2U+uPWYlFQHen69
G5ZZ+OkY/rQToGxZPGxceiduBxPBwOvm7JamBVZjqY/T0qaLB6kcOhdASmkeTeu/
eMnVt1C/1EDz9SRSLEMcLKR/ZWoW1rYahS+2yOzldqGip9DG3JZiJw10qSLNzOAf
ppDdHdpdSXMaioY1W+uRs6cxEpkEO/IhU7IsoFryDsgiZ0UClDrkGP3b9Fi4i+yD
1Llw71j8C6ZFVTfuoKv20O5LT5clOFViS0gv4pqljzV6jUa1UA2A+F+7RZQasyPc
4NU5q2sOtIvK4acwhYE/6vFe9C6B/avcOLgsPk5IZOzuWGHqcVk3qC0v0dtC9cNB
NmRWEyCNvD+iHinRUau58fKecD0ZgAOlyFKu0ofjZ2xZK6MU3Dn9wwZcTuACRykO
/OqOWPA2VLYitBSPE0QeiX+PUPpvktiBd3c9mDEfDtlbKOhus3HOMbqPNS680RoQ
dIymeUv6nCuY77sPIKxIGPdnjvRTiUa8mkZKFmQr4tcEYzQEo0UbDiRZmF1Ljcgk
8n3w6L+eNdRIUX9sjdsjxYXccis6PAOLjzuAsKpQC2HG1Gigk5a7KwYbCtVOdCn5
TzzhUwhe0gnIolU7frVdSt/ipiui7yaO+lj87C4K2iLG4BdehQ+HdrchNm5hGDqj
3j9vAwuqybgxp1V1Uy4N+S/IKNKUYZ5NUlil3ljqfq/EdSiEePhcJ6aWPjCDEAEO
iMOssjnEpLS1rCKiEH+YG1DLX6PVTCafV5e2tSsqNAvJd5X3MW/x2CRtb+XIhO2F
z9qQJZrYK1i4+NjydFIc3uJ9PVO6WcGj2q1bhJ5XCEk88YMI2hmjNgY+smkwZWuo
kqsJmwWbIi0N/lj/b+V0Pw109nBwQNtxUmXP+/CE4owq9vyiqVDKYJmIWPUvgBcw
u1WT+fJPh5bt5/y2Vo4Ofn1KArFRIN5Gj5obAX2cjoffPD+eJHr7oIejSs/NFW62
JX24XpBTjSwtgyeDdYTyAEp96g0WsOlh1d/u9dtviOjKh942sln7rpW6ZfGFTHDo
NdFvV5T/s7yAIYt4muepIiKuu1W+YnyH3mnZXvR54hbqLpNzUtO2WYcfJSSzL8/s
2SRdKl2sr2123JkFUQgvc7L7moUu9SBqqkeoa5GmhdeYhXaYfxZRuEbAnvWKN+Gy
Dm7859qL4sFuMtBiQwi86BE/OZsstEZMaV7QB/q+vb+lVAUBu77MQ46B2PYLnhC2
N1hGwallZDK08UuC8tNqiBDMz+d9wYIYZnJaXqO8sgaGbyOtVGO8LEzioLJZ/JQ5
hd7/W9PsmXxJZFyZaM4cnHHQ7jI9S3Z8b3SN5M5JY1ksvJHoIneJQnDTjl8Me6xn
yc20oZ1lQFZqjGz3/MCuxyLUH86twlvdqbB01TRWPQ8tc0zXp6+H/0ySLXzY90n0
8QH2uoekzbSo7pnGJQ9YesHZIjLqfvYOsKAWS1GBbegXUPZFoFPLfAsf+44OPKrm
5w1jzuR+ifmQsYrnFR3CqtU4HoHckfJ6eF0+nH7W9UQUIKXP1WHedjfgG5H5xZSb
wE1y6QKZdlMWI0ehxZBD611A4Etiph3IF36H/nZ4zEfgKQVlOh6peiKFpbPTeYst
9D2Ckv/Cyalkv1eWbLV30b4QEqB1v2L88S64FqSkekdmg1ehdH1A6l8Cv5OHbqlm
GQJNUn7evyCT7NE5kyTbwclnjcrmIb1LGOaigNUvAq6v51fvp9bqZyeDPFW9QDQi
hhHRSBaFoNH5fITBjCHLzizEw3zk1SbKR4QfanONJhAoO5+r3QLJLJlI601EOm8s
rLhXRfQFtidgYYHx5Thq3KRzUnbGz/0/9UANg8MIWdrQ40kuaHBNKGy5SsSMQghw
6PuKwobVpL3jQeL4rz8hNgc1o4UXsOK+y+9KaWCwQdGTT02SdlminSuh9jECwJUS
wckCFMWMMUINGULGl/p2YNUiOYSJGfmndSIv4a5Ap+pqCLv2KHekYF4yJFbVDPLC
5jOPEhTGZP1B/GYcyBGljGo5BKBR6gd/WiX4ULfDyCE9itwPoa2BABRkuK/F6pzo
69oGxlh669D4CbQgQsw1v7R51soDYpQM1J+XOecQV2emZfL27vYUUWgosFlyk6Il
IsEOK1o3Bbw2SVg6QrBpvvwRfHPftaewrjNQ/RHKSvKAb0mvtofkwZ1d3xS6g8Wk
hs+UPgwv0ymzPR3taonScEkQNjhJG4TOu0hnnWXsaoh3l+f/5R2c1djYYbBgUXg8
/hgFIOJcT37YRn3ZsuwsSPKGsHtP9kA3olIQ4sckKRidPJrL5fNPgGdGLBh6GIfT
uB2ste33s06TSxtOUr1YfFaT4BwX/SvcKcTAYOitYFLsMI0lQ7oz/wz90VPZY5Z5
8Z/PV4XqTEKNXgpkBdIHL13jU3lz+clAGazQsxIzGxVjB13XW0BU9A1Pj8qX69hg
v6sOKtUAjmltCOLzMJGKCv76TuHtTn+DNlasNeuucBSIYl29/mpTaDga+Hov86q6
nFLgrngDeSNGQM2Se0setM8asp49BNLZa6hSBVungbHlMjqa4kjjpNCPQo4E+0Wl
tWo/W4M51/iDDDQfF5AcKv3xRzEYGah0aXB4z47txM5XC0+RmhyYWIphJ/w5Azeq
CJjME+BioWmgD5V0Kk1lwek7YiYJuNsb0f0ECp6VT3nsutwAixAr2EQs7uU6894a
PWXs6yXK1F1fsgSx1+MJP00hMGDEyn0pjAGvKqQdBeWn08vhN9KmtyBOJeBbTS89
PMUBC8EGgS7Xhwgl1vKk8j+SmV/AFi84B3nUaCMfVPunu13BMXGAyqR9wm5pBpOD
Z53pLe/H+oGU7s9AiD3gATQnWVYzW6zPFvI9y3XoHgxa07B9r4fm83/Z1l2VERnd
iWKvXaLTi7xCweHTxHG6N17vDxvHKO+kUXOFPVnmP0cKVJGcrhMKiuIX007+Jp36
mQrJ+IIIMsh+RDFXQGBspbtz+k/YOyxtFi/0xU5Xg4MninyshA4QOueGoUC82Jjx
C/Bbga11fhL8FhERckUSPnUZcTmgnspBaotAJW3jJC7Xw34OzsGfbqhs8Ka66JWy
Yw3E71Z6p5iLgUGo09CMN8abNGQFeKIrVyHjXcyQieW4r9a7np3cAOeVsIFWWVTm
1NiY0GRkDep0EDPkVIF1wUI5tn35jjG05vvGqYHjChO3KCqrbtbVWbp818IBkzQx
J8xA/YDTZgicVs/7dvbocNYuCN2CVNVY7D/eh0djl7OLKSRYUQAh39W2vZq2hdNl
PzV9AvgaT6ChKBQax6a7Wc+ndkMqq8YcrIKwBfT86btVB2QA/lOUYa+w2wXqjmQd
YxSPVLlvj+A6CI8tY9/FC333lGugztfe/U/iToEUIUmGTzjOY1/d4bVucHGcQRGx
fjXrwWDU8UTs15mbW9P5JEf5uPJ1G0lT9i9WTt1CtQVtcEDsRV8TqyzEI0BzjTOG
tuIA3FHnV0XL0AiyGQ18jYzFJi0JGgmpstgmOWona4bJzVluNE+fFefemjcR8TvQ
hVgr+ahD3zc3KtLK3yIiR0y+wn9TZ8Zq3dIEDtOTvwT2xbZQl45AjQE/Q9ysB4Aw
9UvBtUI/3561L0rpXh1jsCuBbY7VGn4bUT3GxTZHslB/uSfHh3u5uzwlduu3YWXW
eMJmNzrMwv8AiZeIaf3ZH9VYwFC03f0EmOr8ysbvmYgbv+ppHhj6hNrd/dKbYbae
Eoi/FoesFmAq7WrfYX9aDvYDJ2lHnoJ3SV0UseiB/N9YmM+xhjcyw9wZqnc4aqdU
lMvrlVTlAxhseCHA9ndnIcwifjiBKeXrkbto8STZTnHb1RkVVRtqTEkZcdPr2iV7
AU3Rv6x4duWQ9n82hKyzLq60YNFoGKKPgQboRVr6hQsBLyGqYKFTEiS430g7Bceu
hsYFmkKCR0vSIQHk+rKILpAsyLN359YBW5GyENh/CaiswtFPTkJVHKHmsFJidcp3
b23nYIflp2DZuKXt+rY/FSq11IqexJo25UXGOou/3M+QL9fjqoFnWCbTrQPKMgIB
7FF12k1gor3s6aPJA4A8QpKLoDGL2v2qcIvmztD6BDB6+1lV/hj/HQdR3Pov3vuo
73DsEsOUdz9dlkus7uNyw4itCVeITS+3dnUltYUrpreAmz/AFNAkXQzFsmYPeI2v
qUVG1tX+N0C0544WgEXvSwMVWC0pfdss4I2/4p5mnNdpwMRLAq5dQ159mxAvEUiE
lALfmrvThbjE1YH38dVJ0OAOQ5+2laT2CLjvlZuu4MOxUoQja5u7dzOvcymZLQFK
J1pv6n6MzVL4LdxDZ27xtJY0KJxiAcINNxBWqWqqmtJNd4Gdlt1Ac5A2iIJMCDC7
Z6P30HqThK69+XSeyefjZxUN0BBFQvMg0UxaREjKqkShyQmgVnoAUb7DkuG3ege7
70zqZ0Zqi1UVdJZv8mY7/Xf+RQY35Rw0Ed5L7A/s36qLSPDopMWE0lSnKK5X2CI5
Z6uhW5ZDMGldyArGoaK3RPdSWDYJgk24gm+aw9pynHZWgyjyUAEgMdZHj9NRE/an
R5EM8XTri7I4Ks/6Uj9a3ZuXmY3RA1R7jNocBCk7gI9NU1u+rIO/tDygQs0jRLHi
wOSIBVdWI9o0eTHOvAYkjPeSCALpQodMZzWjkpM893m8K/q9tZziiPWdtKndngXe
kgbbEnVsrWpINqXyIrM747p0oCD0E1f3ua4pP7q8WNEjnrnEdBca/pU3sEQIxRP3
klY0OIUYOy8UxKJC4M3t8Yr3f564BNs4wQI2DDco80XTZUElk/xKjJdBqOalUUDr
FQ8QrdgDnGkkWUC9EJMnMzHSzIv5/SThSB2neWJCrSwFGk6l29D4xgfREpbr9h46
JJlrzPhYZwfkT3+shBrf5SxXzpUSU0dSxriY1zF3HfM6FpLoNULh3iQBkWPpj9UL
5kb7k/+BLyM62sydwRgZ8PptJjldvjdE6+r7eICA2klpKi8pAkRk8k1lo++RKnlN
F2kGS/2DPi0NREQDegTmOVrm3zANWnmnAInjJsVE1orguLOC2hAEEhaaJ8fi9Bp5
57dUfZuJPF6agI65Hao3c9HqBheqCq2xWG+D3n1D3Uk4jYI3ZrDUnixYi/AD8yE6
h+Lsp2f0o+wpEsRGFs74p8IaW2fC1rAtZpVSVbkY/t6AIby0MIEwYHZriuE5rIsX
Damogqh7Njdo9wPlJnO4N0F1fsl2lXMYEALMB92hFefZ7vbi7Vv+ysXIhdCW6PiD
7ZYXZs6+QM75+G7HBxKA6vGICfTdkqvo5cUBai9PU+3G+wnnc72Hc0D2Ruxx0/oQ
2I2B73Mycc76xjtJx2WIH4rN+P8Tk6zYC6Iyj4C5Y5R3ak+w00ursep+mwVKkZtH
5Yf5RUgPk3VK79+RjtpQFQ5rWTvHy/DADMxZo15kQ3FMXP8YWUT5VZJJfwhsJ0sl
3rgWedaaa49IwP0JhiXnMIioOqOvJFUkRCy73tiRdSl9j22oltYrxwsXMoAuCAyT
D23R5Kz5NzCY7Oi5KhquXcPBFGyruaQv9bI2Z6cBy/P9jJ/jK0fxkKwzbyzhgAe0
zL8NbuAQ43k0xUuTklxWDacA1ZOH957qQq18fBw3952GtpyO8z6lbhtKza21JI10
CC5AQVF2m9T2Hv5nsr2l29cZMNPAi8qxW4imTWTEYqtuBpe+hqNM8B0Ez2zKNRai
rZYj590mEk8s2u67swhZ5IkQ6b8AsAPLI3OiLNwD4C2OMwHlBB/9t4FP3ynMAinW
/WUD0JaHhZ4/0Upmhj6gtX3vi1K5krwkCjQqYeCyNZMDpRY3DUBqvq9BwF/uwT2M
geeLGvczcgrZO9We0maBYXozfL6OrmmlIBT+0a32ohTGvY5sKRRlNqslxRZmBp5r
fTWnUm7uNb0i8u6GtAKNcHAWqENnzSSzAEpw0dOnea1gK77FQRhsR9XibWEjR4fc
OTjlWkWpJ3H+9AHQeIbFdM5kYcO4sfzNK9YUSijW/2IUTCGl5GOjvTUTcTQvu6Gi
F7bBud1n7YMQRWgWVY/BBKo+x2bKLa2NTN+/u0wNcJgr4TRSfnjwrLZi1z6zcqQ0
iDH5+83l64plf3XczMyi8mWYE/ODSQAIILxgLg/NTkmTI9/aiXREzAFAApUfNftg
vtZdzu8/jr5ZooQkQDoXDGrDpmRtydYT2MGzZw/C3X77ZP29f9++7pKhF/17wSvq
YY7LVI/Q27DFPWpHclKf91QdBqy+b0AJeKv4TgZpnuuvFfITnGxckurqQ8isD9bd
VPUZ2GvvV9U6LT0hE/nZHYIH5jb/oHnJFoRNWiCw0ZkRBgMVlOZZ9LMoNjBXucJa
Zf9oeYmdvMzel96nLTKIDydaEeKJ8W02a8/U7sAr8NBIGc2hgo9AaSj+CJbEtzOP
EjRoVwax6gkMGqx+OMCT6cPx4ghSh/0k8Dl6/dxgVCU65EftNuHCyEffn9/6ggri
ovcmJOkR1Dfh1gyrOygEemWR0oOZ08zuZ4Ynvtway4mpchxHIdPjPQASYmir0hbi
0TjurQ4KdNxMWJaCE7lj/j9QgctmgVQ7uxagMCVKXaC/iT42ZJ+49jIh4HjytmjS
RWKRDmgzpJtCi9v2H3BezAvVuMKeGiilVR3ihqqb6gVvlqc8hvNHmanRG/1nFNKt
i/ZPPLeathj5NxNLCpKiDaL+k2YQey2+XmcsHQeHS5av/qq6doXChzgwcFhxoRRv
0y7n0vqkcix1Gcy/80qwaXn2TZJlHwCouYaax6NUCuZ7UJ87m8ECesVKqhe4j6+T
jTazcqdaattPc6vE8uZx7i5JhOmM40obGVPPjxDbVLN5ZeUUU/U0fL5+6PX5ypLU
mY2OaUNKue0n+jPZtUqA11U12TwRnyEDTWArE9I6Xkhw8qiE65vfd+cX5UcDKzek
KL6ZaSt5+wtmLP0xBezuQ6ZXLHLVqaTNkfxFPKaNt/G7nIRaM/hw9LfO8/nFOqpo
27RXmV8U6BdLvz3xcawpaf4TfYO4YEkluhoPNUrxOl0rusF/IkOA6m0tavznhJvL
w5wfuVHmu0U1RoK+tfmTTcztJrEmRt7TntnsZ6I0Rqay+SKJKE4Y6bJuF+A7owcL
rb7byrqB1xcy9F1SwDIT1juV2I1unUiMzdZWoPMg+TCz4+4wDNXaQCRzcKPH/HZd
ODkFfBbcMphcI2Vp4KxLihzBwTU1WWjMLFt1A/qzXv1OGXdeXlGLxUCMMdw9kQC4
yWLKbkUpGTHENSp++mA1LumzP3CuI/ktNnGTAMliyX6uYJY0kTgkyn+UrmqIhpEg
+12imD8Bj55QJMoTH8ZpvpmjzTCX1orHMXd/Ry/PupbXmwtPdV+1FTjXSfUb/NZT
kO72epeWheTcEAN7eZ+AnSF1mBE7rTcHEFYTJN+dLLML1Oe2d1F+egc0QhZtH22W
z+jg9FQQeBJaTmh2gzabBd9+ch2p6V95TWlCTL5Xw2AI+GCE+dL83Mk9yi9rW/Lj
LgkdKce7+mh9va7yS5jevDsbdnbPdsTW3EVaUPuTOtvKzUhr6WssJSISGFOX1W7x
D+j0v7ppAF2jBMyYHFtK+gpIy63c0H5iivi0DVzocztkb/gFvdqpA0bemwHHhZGB
Q7Q7RttwS3roAoLSsFE59yTYYP1vok6SLHEtUk4ctMe8y9v2JcZXKjuITTVmxEyC
CV95M7FRbu0CP4jgMhJR9AxrmiXD2B/K5Eu3tkrtAAE0L1sxIyyAFETgpyXFDIrv
Vno4X8WR7ecyEWtfvYDl/slSkM+hAkkppTwm2GTy+I6Q+iX2HA/uqPoZ8oY7ptEB
Gbb+oPWKvAq+Etm3KT7V/BWn6RVlPKy/7WPEQG/FS+24aksi+9kN2Ebg8XNyNJDU
Puof4hvTjR+5aOasI0UGf7CvQmfM4ns3Sf2PovjxiySuE7YrlpQGkSpEwuvCo3aR
Cw+RjcDlALmlgLjV+ml8MNvv1m2KL7Om7KOnaO2p6ONE7K4X6QXaRC2KkUkToUeC
19rJRnqOcMhmXmLXWawSwrVb/Ex+1AEdZdsek0aBlmt8JbCXDwQlwe819KbW4Qrc
Z9NklQGzNwYvqA6A9bPpiqgNxRFuhrh+gJyGsRdh5pKIwl3ybGxatTxfN7daVYsa
0iNVYJytpD2d43di+DvrUNnAELFnTc/3Bo86h1jQZx3cDF3uwIqZnrxeKso5PZRC
Mw7rXwXmbv8wK1r9qRjmmuTCxq06isju8awV3G5u4gn7cJfQQhvtPkaNhfPnNZaY
Es/ngGpgPsbXBieQEo3rWM0qqhk0VQTVU5OjlWGvtEcJ16W/riR6gxvAVhBdaK1J
Vi2Y/qz/IecWdy94SvRzrl6zVSxj+Hv5oDDbXeXr1pEcUAosIkrI/2MwddJ3P2zw
SnF2qh+l9jyS18cyZNr3tmJzJEK/czLe19iUf61l/b7rCnf3xg/FhPvZhYmdegJO
8+0RF0SpVMhZj+NpBFsBTMbhxYvMnGN/c1I6mWDrtxlbXf+vHxeUbQb1G3TUG4AE
J/LYNEP7WWcc5LwKSwRcP0h2Nef0yrlvZPj75NhFdkXRQiBIiuGZIyc/WuZLSo0/
tX6pL+FSkM1NlYTdCXAnXHygZFh5fnthskAYrndQCoQfOwe1KZ8Ipa+oTSLZzwUE
6Tm0QCzDto28MKbGw+WfnU9kH/repsZL9pEdS3k4J/vHlEB7b7wFA3x0cLEAxuAE
yTNRoplylltlWrJ/2zdbXoQV0zaBN5GlhK8FDRlnQXP227NDm9+4KHV4W1CYwqfj
nu+zo1nM8/yRo/BBxMB9l2RRa6msPfpbHPQpT5KhD7Ux/bsptpa5+0yBfcMhmVTB
K9tR4C0Q8ARmeeMgi+1sLw19PjKc47tuaUeEnUfITdK4x0WjbaS+sqGy++UkPoWo
3DnL3ZwxnLbJgCNbhJUbxa+lxh/s5sr7+LflFkfUJOo1dAcQtLlUkf9eQ9nhXcQz
77Tox9wQjFPFhkh3QKWmYHJrnjK8k2hjZwJXBJlvP6Sw55jScW58sL+YxGnW9kRl
/JzrK5/N0vrwc7PBQa+00ZIIDQkD4s9tx9KyKcgfng3FgW/MVnrZOek8c795J8TI
Ire6F0BAHXfftKQ6Xl7/9NQjDBXD98pEZr398TbJMaVwFIZN/Ms5mbeUPfr7QxGU
xOvrTiIeThxJfF3FLXz8O78hqRFnkTrDeNE+L9TaEw+9dKz0F/8rXwwExOwYkxZn
teOAHU/0n6KTmavN40NKz7Q9yQLXqpdvvErTNmEfZVMuyFuWr9ls9UK5Z1CgFswt
EBLwW3HEtG5ujgQz6Z+UbIcVhkAHo8+ZiIhjL31bqT4Vyev3meQcfKN2LabcCLmo
we2oDDzzLswEEjdKfxB1gml/sEBnTge8hLcU1Wke//nTic1DuuB6n1w27oitMfCB
CQorebkPICDE5FDwwihS0HQe62v1z6mUzMYGxI8KdopD4VXn4+zUnGbd/vbhi2y3
ZIc7pluXgQdBNV6KMMALaz7PfvJSE258oSVCtrk4GMLxp74HSj3PIqhwLnSZey+j
Qp+qxlq3XF1IgJVoKYNg/tJDJQdShycPTeQ3YJJ9Xkls0mIXKNHInw6hB6hVZe8a
mB8v0XcnIchNplKZNqxsxuNl+3K5TiY8sIMEZHWNePNmVNuKkph/QcRaD1kabgjP
VnNxUS94zyXAKpn9UIQBo00A/kY6v0IY1okWlM74zggXdmEYt1/9lMTv8EYxxA+6
gOORCrfGPsITJ65dYSWRz6S1rLzBJrSHgchWcU/3DjAChMCRXcS0wpAUy0uCBqTC
sfsr1NwPj1eMxQiSOHystuL4En/3ZgUramuDiZSZHJ5lSBsXcGdle0ncsWztMPAs
R+11WGDrU421nwulVW5IqA0jtUZoFmeA1K5TFaNb+eZsQpW5i2qRP/CZEx2zIf48
0/OfI70Oyv5M1XwcuVIRZe48GttIoFkiMJJ38jJrKTQ0y5bwYniWIWWhXLpOHKA7
X08kvsfLq2kElMXP6xzqjxo3JahsyvLeQBhjIVmcf9KRm/pJb3x2UzsipzSWQxOs
gVQnVAeIAfhwiXUBq8e/a3bJpKJGcUEl7g2Ohb6P4ypW+sSJ6YkmfEZW3S82AV2Y
esal/lOZHMMWu551IuQGq/jLKlrAJW+javYgIiuSPr6J7jUuDNOTtEpDmYwKpkXJ
rkzMhD6C7CA6BqPyqOOgOMteSzNnUPPhPcNIqcBI8XdTp12pEU2PUYWreMD3wv7F
LcBj2r43hx1s0hz9UKyqN1NJ8qJBn3TehTNDAQwjWcERUzL1ZFujzm7E8aFPj0AJ
tWMTb8oukJZ1CtAEGUcx7a89/1qY5yY4ADzdu+dk640PS11/U3+PR4QiTqHBunnW
0VHsOcNQQV7o+q3zvDACHKzPZ05LkLHjkYPfqoY6ip+1clsHgGzBa79a0vWYftXf
e97e2LqmL4IoxU6wFy6bEUygbXBDch8Dzx9lFyK3P7icx+vqaMKaky8x0suDGRTR
iOpUcgBrYEmewFkewuRNAfrHJohZ0BoWPTvZxGUSX3WndsrHKZ6lKRuWkbBuG0ko
QteXkEREFLb1N3xW8CZh3yCeu8CftjGYXJ524Yg0rOoqzMotR9PRYRaTRcrVWILu
XBzJAc1QImNk5cAme4DnBJA3r4+AUi4ccM8g2c+rZvJ8dgicaTPiIX693vK6cgQw
dD/d225jb0rx8Mhp9NI03BARXoecpWA2BTWlphxg46dRY37/Km8O32JYXUOM6YP0
71B5jyErTbYLG0FQQ+sa6EjEWy8wwa6Z4fto96ymfRmi2UT4bmSRHZifSndQ3Mog
3WbgXoiCUA4HF7mHf3D+WEXpM/fvTaozL8TuwWScRBvCt2HniCJaoF8p6OcMRW4I
8vxKV+g36PzenDuePbLNgdxrGlePvCuCA+ho1x8ol0mjLA61DZcRwczVJacDsAhU
ivTnGydJpWTCvy5lZJeV6FC3aEDtq9mpxeIq4VCxLObxZLA5iIqA6z0YPesFVMcP
/b43oU3bHrGXk/0AjJIQeEay+3hyVjJErVupHc4ccGK5bz5L1+P38a+g98GEJe9x
EqCFVbPk5Gwl7zZi+3ol+Rvz+S1SDXtTXtqWsh67hkDoUiWLYREfOvE15RjRZadr
QXfhAyfT0Sd3V7uBUICJ0s0f6pioxjvAW8PpI/xdbF9MAcoSv2A2nEEZXxViOSA8
9LgwIlIvy0YPzCc5WR8S8Fns/wK/pC3t36pBwrL8GjgLUiJmQYmzLVDO4aeJbrZX
a6gFDs1FmryoGx7lb4tCEYsCCVub2ilLK+ymfBGjpNGGKxjbaiO73Iy1oRb2IcWg
BLSHdwR89NfAC5tqtFYd9t8Ey891+y2u5RKSof11SwSgCZQ2oAfj5BAyldm4JmxF
Mi97Gf+VdcbVkxAFEqJLA4SYjbfObMFuiVNLDFRRXacf1F2s6BkqROD5GRpdm49p
Otg4BgdVDDYFy8N9TH2OaQICy2MIAih3oU8mMCVcD/yZkt2An47R5aqcQh3kLkiK
BpZbnuQR4jwkayeAyYJETiuMWbV/ymeEM8sPQpo953kKy+qSdrFz38utcOKVq/v2
TJB+/hzC8b8vnq6OTkOd+eWNzwL985Q4tmrDgaQBJ6kMwzZMFwu2t9ixGcC3ApqD
V11zoq66K1j+bnYJ4rLwZW+zIhY0wggh9r3Z+uo4zwDURYfB4IntUpjHykQeLAqO
70ABOUUcnZEBK6jzNeYTum3RznNUBCqYwhelTaEwaeTXYMyj/Aog3Pj0DaQYY/XQ
ikPCptni4SLbufzZgyPjfJSJZlU1jQuMFljrzb9Gj+0PljjZaty1OaHrnrla4ood
A2MeXSReeZ9qFjompOi6NarU7y5TZ5U7QvHKs0nmOsozAqXT+owojXzfYoxPYFLH
E0z5YqtgAaal5nDkm0WdoSzzojEzm1jcTlCHe9+ekILFwveX0P7n4X+JaFMkSiM5
YKPF+/lqDGPkM9j1cFSbp9pYA85SHd/6gNswhJjr+Z25KUyFj43KK+raZfP+hbSp
D9jZK+VNZwJlrvIzSXSjlR40unIBYye637f+cq8LLPd1d2xSa2axbqwTp8c1kI9U
HZmTNTpfoNItD+hALx8Aua4gzbe7fKISQoPp1wFsu+U431lT2joV1JdZsnHh++KN
jmuzvOsdMNyw9N2QCfjP+/IZkAWAEiw5KOM35HtVHVsLSAN0a394RC9UxDX0izNr
qpE3o/tkx7HDADv/CuE0QEBCvOJleenPpgpbdt9FRwqAo6LxmcqQUTdpude1RXZh
5DHB+QcZ+7w2O4R/u5MXFF2jSJtYCKugxNLiUTn2/+hBIuFNZjqdz7zsmdYa2ypy
BGBgIdBz5vhdCa94RB8a7RmOUr+Ud56hTI/2YK2SzPJqWLJjX0j/jeoh/Rok541J
TCIStvZ+zpJH5PDG3zy0QulZ2C+C7FatkxTeN9TMOiKb7R29bpQAsjdB2S6OhUJP
mkRoAj/al/dD7AhK99jTd9AdEATQ+BlPiGIspJ9ECKhYsYUGmTqRAeDueajWE2km
B8EsawVL8lptgf2WV1qJwjt5ySfp52SWRa67I5JUFyP4MXB6kfxqchsAbgvtHK9f
eFxkFaAk6iT095F5vZuRPGmmNbxpdXe0B9uu0LabRM0bBCw+uppAMpKBiGSpF+dy
DDM6QbO1WSw5h8zFKwHBb7j5FSi9Y3nRyPH2E3MaN6sRvy5Db7nshVqIJlUaJZ50
lLkGmbwfA3/5IBghiR3Dlf9DrPqk9gkiKNwJJZOQSoqB2o8ymUAnQWvKTSe5H8P3
wMMblDFOdMT5SUXWTHF1h+uThyUMv1VFjI36fk1JRLErdp+9oGxQQlfekNvNwhT3
7J4uMLspyCHtG9YGK2apJ6/FGVcMLUI5L8KGTcPsVPHuvbSOhxGa9zW0sEs80Bdo
dAHp8Cj4Ud68XQayWF9RUXkrjaLDe39ZdNMDp6qsUDCYsoE3xQ77YaJrEJe3WKD1
7thQZD1GkSUgrJ3HabJ50ERh0+90qA4GJydXNKnyM2VW3kcNYyJplbhLG5cSvu5s
9ZnkXtNI6IOhbMVXrR1DAp53eRmfbiF0kDXeqRwxAlE4pXKd+E3jRg0DKl62Trcn
EhZdD9x7UbOu+hmyXcTn3H67C2dkGjLVqpO7iQI+9xMl80re0vlULdzK4WOZANoi
99knebIc902EqtHRo47GuNsMEGYh1PW5/sPWjVRw91pvhLIHSEC+HBdb2JvMwNPi
tHe/GrD+p1zzOxrC34HdJeGkdkRIY1H4ATHeTCC1CCLEuTaPDMfLZpUm8sh0XWpV
pdULqJNlrJx9F0C1Vwy+rPOljGTXMKn1nX+10RJEa3WdP6EEfA5eT8ywI7Xq+4M2
yKGoeEPz17vOQFGuoW/tLGxrwDMPbbg/vxwsTBPsJnMvrWa1YDsE4EN0M0s/avsH
K9CApMJIAETZARrDchEAsjNMNovqYyWX2pjceUzCZDV1dISucP5yCddG2p1aFjxu
s1uZ9jV2S8KKuubHgWeFVIsv3k3mV3R5HsoXLXlFmM4zj28EL6HaMKxh6vIuFTx3
0nY6dh7VeU5DGMyBVtjL9uqcdL3Hkykw5VPV7WuotAZEjkeGUeQwIo+n1xsUti+C
//NWBi2jyxMydBfsc1CZW4HNDB1vkXkGZ4C2eeeR1YVgyjhvQrQad21Wl4C/M13E
BuEXm45w76cZcW+9CqFziV4QyRk8bwHy8X42BpG4Kd4xfX5zIFfCIbuz4SIZwjwD
HBx5vl7EXMegwJlRkcBgJ6KQhbGP2p+FCT8FFGLkTAZUyd4A0+fZOrzhrsm6FG81
fUrfRr0AoysEoGFqaxYm7bnJgbbEwJ8uD6z9VgH1HHvwhqfcFeYbFdeLFY/kH5As
paTyC479HNgOoH+J9Ix8SxANAyPsqbB8o5tNmUZ/y5fuoeLSmvdfKlY7aDx61+w6
Lhi9HhXPRJuGMb6Rp0rxZV/C4cXZboZ8slR5HVPK6EiMb6CZtcb+VG17hKgvp8yx
D6puzCSKEI1r3gbOJkonB6S+3wmjNaUTh1d1Vdvieq3K1vBYgtNEtaFWcrtUWEJe
JbXxaCWjj0V4ZbrOyEvalA+JDli6wvWMhNlrHMpFfucfbUE3ycl1K24135V0xxSD
gtiZnc1Bg+4L92MYFx7TdTiNvuw1y8IH6Z6e4SpQ+MOc2BKS/lMCUQVeXhjsUJmy
CFFcxQ4eUIydY1CmEUNco9N+W/0UudCz1X4NXX8zCc+MQDWj+VKJ/p4LwcIFQ7op
AocWHZFMCW4KHTxFBrw9TXI3NLCHwhIbYvYufdDY7MRhWKbl31Hko0Yxr65Bm312
ShP6waIp0D4EdhERw83jlMRYBEm4Nh1MgtTuAo0wm4Gib61K0mzfYQjsk+BoXrOn
JjL961DA1aD9iwpq/NvDLulssQgdB00u8p+HRaL5uEaibsNYLfonoFZHXqJL3w0D
GJBr/OH8IRzpvGKOYprdb8w3ffy3nyWLtb7ecNliUwOgzSRC2PkRTnxSG4jhQa+/
V6yCclKlPyz4OQPPKNCCgppP7n/eSCZFPjOztZdwhX8NgoI/SfYsuw+P87uqJzyb
XFC7erEm22D3W4nFjKR1YxreK55vAtief7Ll/ehwp4JhShld5yIICzVBNRpeCzpt
c37eYx1Jn0k1OlpuQn1aUhOLzNdbeoMswvVXanqdXklNzhk0dcOBeElJc7XUbHc6
nPf5Fl2A5GKYab9PolLG0xLDGQyl2Krs7AwoJ1XL12l9MMiyDlbV03rYHTwpa/Ly
4AOk7UWMFMhRIn4e+VZF9UrNf3FuYACnEQdrNX5hOTPoEO283rttI8oiU2YOKfBp
VomBhAO+4OzYlmuaOTF1vVTJcfy8r7SELnm4Ppi0FtqLiiPPUs13/8My46U0Jye8
8IKgWEpofo+LmGesvmA6+mcfT0xqcAUOmSgOyIeYI6NX+VNtsi7QSMMUiD9jFoA/
/rl9bUQxFl/qa6eUxTe3qlc7eGYzFGv5670imcvG/WIOeeeuNZVLigdVGsgtkp/v
14+FXgNvtxr5PXQsuMEPrG/lbtbZRJZeKYs7hhZqniMpvH/mYLl6eK4JZzX/vLOq
UE0nK27F31PkgRQzv6OhZI1tY2rC8xGnJnb+W7esteVkqukXeEVK/lT/XlgCK0K8
lj7mEPMB2r7cmXl42Qkmb0Zx5shkB7wIjbmREVEMO+8oIHhwdSyJGN2bxzEHva3E
IHOSHnFVZPzTXvUdrL8DkbRd/Qb257GpaewWXo/aZkufdrj79/LOgo9svX721kEh
7g0uLXkZSmD/ME6wrlCQ9GHVGLvaGE25u4jQIS71u+MGW2nykzQpai+OWVMIpIzf
LgvvH/2bxPCNke3+tYMhW+YaYfnYDG4kw+XFYCkEMRobEQWaWp3KQN6NvbnuvDEM
cOYwM5rWl3CElzgcbGTgUSc9uyNuFlSPYs7F0FMQrHYcz0zwuLWxN6q7l85dzhXq
3FbfRhE1ZXOpDlaZJMKle+5GudZB7F+EdHygS8CTZOD1KxVWD5OQorNVsTIONWTm
SiFSIP5AW2ZNe3MJ6njklZ4JkikjOONsemIHFQ1CtBXc6tBJsaVO4dnritrhu0ix
sGSo6Kf0kQAM8IRxTFrIxIngrUfIORhcTGWOsNB+rx8F37wA97B9N+Top4VlscuR
ClPzAFpLqR7sHZKRZRrOU0+eVwZTIuRbMhyDQNnPPL0Fp90ORO+LgOuOa/amCaGq
FGBlQBkAJftYjMgTL38KUZnVR6fdRF9mBqTlyi/4l2HB93n6epCfIFAYLVqm2JDM
lTWDDuw0RgEaO7TsrjZp5/ls0rTAiqiaqIzFgh/+AZaLPPNaGQUvbVNdFnI29gQQ
f5XZ1xG83/HdFNH+6NArWUmL0Eyp6nL/bjGY3eGJOyinjO5ZWtn80a37pWDYCfuG
u+qbJHOwIY77ags4CsYctsjF5qTTjZnosJ+orO2Nbjhl0fDguRGkuOVoPXy02YLr
njaT78PyVtimJAc0Cc5yxQF1Xd5wEBQf4XFcDSX+EBmIfRnx7YBtCwraZnABKb5l
su7keKWRkZ1I2kdPW6pL7Zuv0QZ29fUosaHVK0JmmNHzZ8iCAa0JBDR4iFpZivtP
Hxhx4mZ0gdNgrp5T7Y7o0CYGjlLIs/mcy/NIf48+6asUjepMid551rFEt5/6gMhI
ajKq0EC5VZNQbl2OPztcuLRjbetvdrRNI5DM030axJZF8/fCM0PcBiBCiH+t0D0B
sfQyBrxHqsxCRGuJjmIBsGzOYoQLcWbH/soMKIKr8gVdz1Nhqi5uwPdhWFKNESNj
u4YPUwQNn+4U1usQiZbOrJXZFUgK45khZNF4vCzcCwlB91zvDiBEO/zquZbcYCTz
h4ItqKb4V07oJFRLZLdraxGi+KXbglgpIPWTdkfusq5FAsN8Qwp/f9nr2ACX9KaB
zR02qLYFfbpeCk50Gy3vQcho8OohE0mw8cswKhKUS3llRo3NLyE3WMEkksODKwz0
a5N6qSinzJhnyy/ZLmXN/aFuaDVwe/9iilxYuRU0gD2ofjQvwXvIufuMi4/+j8s/
2LBV8Tvr7KcCBWtzMSVUK5uPv1lmnfrYK1/K+ND/cyFC2MlYZqwp+vKA+y9IVput
gUT6pB4WIpARLyasBTfiqRRCJXmGhgJOuYxC6BYm5PHqxC91X6CJDnUdyofiShI5
LPUe6adEj8LVlmYrRrkEiRluTDAqiNmZG2xeuzpWkkzCXWQbiFyMsZqtESXyXDAn
KTs98YSUmlfZ6JSNueP3wvBSWnaqxR6mmHZGFdkoDfQqsbA4UMbH1AUglPc8OeQS
Y0h91jvInxJoBTftXSKXRYJWUnYZERK4GcV3wGH7gBOuUbJ/GGeRHMYYwOzd7DX8
0WBfZnS9RAXWLYAn61cxRKOrnI9laXAKQCIJ/UX+6He7cFnle1RL8AylJM0Mu6Y5
QkcPr+pDr+EJDWnjorR1OuT9X8VX4tV8/bGT+xHyS/Hl3htyNQOOhIo4xzRTgK2m
Ihfd5dBs+NnQ1GXhBbhxLvZy639OR15z9gaH8cY+JIr9js/mymszwHAnVq4NFplP
EQoY0JfqPsmYJjaeJDbSJjekDAcmJfTZ452h74DBU8dIcWF+Z385KvPuQjYTIE8l
n7ajHe4vSvENPm8MqzuyF3xs43lw7JLnMIrorIPMKK1fFvK3+fYCZ8D7MpBXeQgL
WALsP3xWPtnSai4drpWGFIcxAg5IAqqage602luwN/L3xp7E6OGp/dLvy5LjK7rH
1wRRj9cAKp4jj2zbKhnmRz3jkmmekF6YjoufX3CVBxC2kuACQwIRYXcVexTnqjzS
bwRWOb6m0u+qpDrjK4zOeiX5zjHl8H5HjTWD6/+hD3W/ih/+HGm47BLX9h3P7yP8
8sdB8tqhuiGMYSAztNS0w+Zup1leOgV5o7Sb+fcQByQZdQNyaaXvAM9jcNtHTueM
iJt/B5/ulyuNCkUaGWJb6r57Qa2rceuezVuZYzMJb3mKSZiVaBc7jsMmUXagvrWG
Ogcii66dKRN04f65QW+tek7GGp56S8N6Dy53vqPNkewfxiyP1PRW/kMgIC/EsFE4
2UzF33qec9YvCfeGArzl9LAPZRIVi3YIS1pIZDU9u9Kk/002JAXEmAM5apdkbj0L
+d/znM995HuUH3qobCsWKbQuO5mxx8w7sIOK+FKW79BYqDUeYXiYifA2tMy/hI+l
zM/iHV0Oet6dgd8aiZGaG6PSnWvtyBKc6t6Yl+nIwlQUYe50uRF4lSl46OP0Y6Mv
6ijE+FHwx2DOuwXda+eLtK2jQjW0G5MCppY9tW588UNPuA3EEQE0vSRQ34o94eme
3jg1O4V74tMT+Stw70m/k2puHAguSS6LDgdYa9Fsse1FL62huq4pq523XQ9Fe/cD
Q8MVqjiiiE2XQ6wgWhzarNlpZKAi4VJl3QEsk8dkAQ0eH3G4WF7Xq25lNBkB+pjy
6mZxzX8k463Y0t4PFYNME0qNuZXJ/EZ8a2EgKtFKpoXrvOSJMW867P65+WY2R+uo
KgqvBBJrrQX68f4pzKpG0HZtbwZUlKW2UwnImBVkxxEA3e0MBRgRMojurpOWqji5
fyWpqyrb4G0dgeg2I/sHciDBUR4NV2I859iC3P0H2/rDdD99K0XE/s/syOaNqngC
PbsP7tn1CxjbCESSvrQ/2crhY1ecZKkQmlRFjyqnPhdpF/flhW9Wz3NT7TcxW7JO
jPwzhaHSP/w7Y0oNlAUCbyJjptHJkKdNt0hn1aL26tqR2ocE8V7DVQNpx5ropx4J
3osXSfv8ENgbA3GSzYhMU7uTF4FmSuvirxeZKHdosdWxnMZZghuTTKhEndX3unTQ
+4kFxsV2PveBvlkFhDXWVDG9le8brOJmWYy8CUTgJVQC6qSwDsRAJAziB2SBLHvt
bSvt27FRegti2W6tFzoSfAC4bfM1NhW3yo+RQWeNgQfbeOYcN8gCYAhwifr/q+LE
Y/rtwFRHXUAkBL4qmuzeIovUKWgYL7esPvzpWmG9obEZd2VcGdnge/b/4mOktxlR
dAtuRzO8ybfIAwym/rcDXvkF2OOfKSjZahg5LMZ2t/z0okHcVeetqn4ovNe/8TFC
vYdQvG7cOlBGq4QdvQOPlWCaXpwOJo9EfxyGyzxfcwUT6wZHdPLJy6ddXoATZIh7
WuvrVH391RjlAXxNGPOQihiOm6x0kyS9G16nnxec3OiyxEmbVaL/1ussHv+imU6A
kdrJe9942BzZKxlZgiu/fPXo1RtN+nm4bI5nkPbLijOJvunVn71rq8jrvLVYp6/j
m0EKwrHh9px4UTwTuCEwVFSwERPsX/kRSV3jyJ+q3aqPxtQ8+KSL6PeCE15OQkJh
VgaX3YIYoj51uNU9Xe0Yon9yYsaf6Xd+4hdUK6f06fxDTI9VrShJaVC3paVnaWmc
xBJjrIsZVlCMWXwRNT1PRMPuBGoryz6CDy6VpbkmTso/1Xozqu6cyFyMOQbMwgBp
Hq4QKQESitULgMQInEsDxPkbQ3fpjwy/hh/h1amGmFcU/6RPzlR0RyF4gX2J2gWK
DxGoXg4CmFLhmHq/emiOKa55T0UYeSdrlpREtbLdbE9dwHM8n89B0DXzUbgMn4eu
N8qEIk0+rJkAaSTQAmb1e9lEJ96mqmVzY80hjJRcUfMUsBHvkjXjvbaUCejoYh+H
VDqbkox+fztFLfXZ0wkYtkMrQ2Xue7Gr3UqADQEsXC/HGR9F3d36+fD8OHcGb53H
nT88sePUWGoCefmatHiDQKiarPUrymymrd0arjEeiNvJ9auUBLtKFv3UsU71StOz
1pVqhtusPhDVebZwKaO6/lVRcEqj5xF8wD3dNWYbelmNy6/+X3zXI4ShKw8yKH/V
xIe4j/YY4UDAl+aYTYzA0L02U+wCBi6O+XVCBLaWuQUcaDGvFAuGyGBE3NHK3NkU
AFImUxZ/tp+jkeBi6f4iWnvt5VTi4lLLSWvaw6vS+a4QhSiE0y98tbnoSPIP4RjR
jUC+bs4G1kD+NFTskqOK/5/c7aNFZ40wbGVNvdENoz+d9ClvH8yYo7mdG6frnNSx
6xnuhZ4L3MhqQhsYAayyxcIiEivSmnv21yIUmBvsADPHDc8XMCHw6VDke0WUjhpO
J5M5tE4bwcaP1xZo5oinSsWrHrfbNm0jCVA6vzi4BuVoB+tNOCVzWdhBFcyAUU4v
jlfdx8zS5jEMDi4vobON/yEUpoTW2x+RUs8c7V1yV1bpLar9aBs4OqyLeVSjbF7l
GtSD9SgGm9/pD0vvb5ncNkNgnfamvJDsQ/MlrmjOFcur0pb/YJ2Ux1o/A8p7d7rE
Ct7fNY38axlBU/Fg7gW0ifs3p8qgd6V9FqBH5/fXCDyb50OwpDZwUHxghnU3UCq8
SoR9JKqvyV03DhU1rprOuJsKHl/BxFDrV7X3KPa70+IJpC7GLsdBYi+NG2RTja2T
pUQd8cRRcErYYrMVKfpN0xdXNSFaLcBTUdstjMybwvXoUv+G6zTVmmzXWqGxadnH
/l3Wlu43Xq0/m8Gt77pY8Syur6sz/Qbr9zYkoNtU4KpGwqjqR1iM/68+OwObE4pr
rmgPtFwzYlBiFQT6N7/jB8R7iFrxVZdtPG+7CPSSZp321KnBz+EfTc+DEl0OYr6o
Vyp9ZuQuSyiieYSmN4884tzmJZMCOjNBH/l8E6Z92uBPc2gfoMSctJLApIpMWwqn
mzNDeev2BWVb1h/jVP0E+pLeDQipMw1ZhNzct9HgoL/dvs/Pmdo6pVHmHtNf8nqg
iROOK0i0Ngs+MQ2u5ly+wIS/hpYV2uPahiDGhWQLjshU+S3dnTGQdT+C8w6dr34Z
sJqwekcmlihmkl3IoyqD8jOxnPRW13lfpyJU80KWKeP5TdgmYt9S2MH+Sjv1JWKD
rt0YXF+ZNTtB6UTsrtC9caBBaT+gYEfUHUxpfBzFuLjs26m4CuDPGQp9vU3xEciz
eq7m4nwF5J7C5HPHsOY2T+8dK6PYT9tSjaXpOWvx26LFOGrvIC+G4E3XG61ftSqu
ShK+Dv14hsggVyEcSL7NJ6hkBqPohP9481ByuORTf4KWrPh4uIEVGExUM+xOBaU1
fFzd4VGV+n2yakGnCIRi2QUZgwmpvgYixl82+Z0i8MgrpfxtOlTpKFdfb0JjOGZB
62YWAqu7bpp/Hkifwu0pV60mF7FBsUeaNMJcz5tpQmCycnZlFQ5AWipuwaXERQtu
WlKaPxUFfaPU28GiEv/hczabKHxG4Q8yX7ByTxIQekCGEFU6oLRLzgQxVFdfS714
9gkHkpI8rv+CfUszssnge8Z8DZ6skMUCQjSlXIKuSdsyHRbk4mYzmU7YkV8mDJyQ
akqeCHop1qyCK9NJdzhXktVVGE6fQAmiRVRjSjicHic/Kbp7VgviHozXRNhdCPM9
LxYixZ7UgOTeey9po9OyjvBMo5D0WBoP3EopURwOWTa/oJ4SMLV1b+4pUxtKtYz6
IADBFH66vxwZ/Vcz2TEvwPmJODvP6i7wrD/UpO7LJX6LaXR+1tc+yDJe3k1ZL0xu
jsijgU0xaKgUwmrRcaYroLjKMIK/TWIFKC/8pDIG84uzIfjFzygvBriU536aimut
F66ScV4T6yOkQ71hax/lHzL7s/drUiRKCq8JYCVS+zYaSO928xiJLMJJSi/HR5Wi
axhtkY+jkjYhLygDtEtYWECC/ZgaLD4WUXGtiv74hn2Plo9tau2Ewd3LLYZOQwyi
KF4d88XYZCirgBJPs5HtZMf8XAZ7IpIpfjVod/bKQ9hSGGEa9SJNoVQtRTdadGxL
qSWouMKt4/eEkcscoKbEQ1gnAfCetQRDgC+pKGKxfbDGSDlfXxd5TQRt5vrpNOai
3rnhU3tJkR83JHMYhv/Oqi0qW+aMOBTTAoic15d3Pfwz/50pHhiu0QEX85YREnO+
V3jq6UJoiSodH9M6yLiXKEoVkYyiAXwcFmVYisv3XdBwYsBN+aVoGQYROBj0Q4hY
KlY+SKLUFgpPuQk7+2nAsKnLTqYZBEhQOKV0oJByZkxPdYb8BBHQTVf9glLS2vF0
nuVO4X1aFWYhsy8qv4gxCy8BgCyZbuHWXe27UpQvUXU2W9M2qKLvRLaw6Y4HaLfk
kxF7Ue2HX0ze9skDGaBNx4u9fljpo8MtvTMl2OJgIt8IRO46Ofb9d0cCxNNAIqKB
1b2CRKfW7cH9kV3k12SSq7Wy/z72uyI7Y4yRjtYAz8kE7PWscOFV61TP7kL3lVlr
Gb1jRYTKNYBmMtAWfR3UAhoNICEwoUYPAyOY6qj8QVii8o+ODWHDbAz95662OUXa
5RQhM9bdpXzIYSMiPlV/P/iLhdICCmQlQFIJce7/G6+yuCnyE9A1gUJEZhUKPnIO
zHYKtRhGMNPvU5IHmIFHNTuepAjGk5F7gqCm/yRjtJE4i/rKiFRXl6STcuGu6WUd
1tJk9jIwcaSQnMWyHCSQe6+Dunt334UOcyAQdeAxNm7nNWGLvx8DnBjiVkMBAEca
Zl14XoT8ah5kn72KUcC5xTO+Vw0ImkUOjMvZ0fDAviuqeBDxPEForZSHIEhpHXES
P1seNg3Kq7TJhODcP1Ov55cShynrf7A+94x5nRsJsVMopZXMTFuJaluLZygkK1uc
40JaOtMbzkdm9C5h8i2fO2orOMQ4TgL5Jpfwucn2AxtK9yrNFXeCPkluibsQVm0L
pX+f3ySQwDdWasUpwSx8Tzk+6Xcjh+Kgjal2HthVm+FLNNiIcjIEMdVpgO/+kkFD
hGwikR4+zHnPkxKWzCGfSP3G3vTvzf90EHyuy3FnDM8UeVaqCAYX941Y72HLiVPz
3CIAGNk6J/tXjSkN1VoNBQsLjbtTd/lAexmTbjTsfuk6ElEDZVFGerkk50ri8CSG
gVYFJCO2cemToVt9FVKionYwvUznCFvq5aUuK9H3QOQIEgBBDNJsXn0WeC4AV75V
LiOTAksby6NiTZ5N3skNv6m8BQgfaqNLtyp3HxnX+4RZPo18lb7Y80J4egqG/xt6
Lgbk9GS2398NDEkx4YkdA8VAaDOFzURBcCHlrKgjAXFCoXRTU4omm+SCqYZgc0fG
TPPD8ahWL9rm2zII4LCsGMNPD7hzU9fJpxs9LOCN8zgGwr0X32/AhM7lStwnpuTy
iJAfaHCvgy7ugGJCpOMto9TBFa8N8/6PrlCJKSRJM+eI8KJ/B/f/Gem8WzOS6ixj
C03MfBQdDBpIWQUcMajJme+HmHuqFHxn7ybmTonPsYqPkOsFDbLvDfNK37NGtGbL
7MvCItRUqzME+PDPQ2fOVW1RYiFkXyuNJWfOF+hik5UyLTVaifFjyTu2dEMkr15K
Xt/p6Ungxx+ruO020wsuwvWDHNgoq3UJRvuR17Y0y2wwur4upFR4x1Ixe8lnW9tP
dBxUW3ZyCxkXxXJqOjopELj8AEHiKvBnv6AQT3U35bc4XNmw27TMxnxWzbNhu6gt
kQOpRzxwg3auNbZ1KTH5l1EtAVgW+XPsPVLzVTocOLbcew1aPrMmrASl5+C+/N9t
MRrlCKHcu1dlxT///s/81Wicl8CdGr9NvH8+vcIIsiNll8jqzOnr9n37zByG3eth
HERBkKyLO7H/7barQ496VMIDy1Gxl2B8idPnkLJ19GukibwJFYE9h7NxV/XGiIOe
Rp6svXsiXyiSJWdqtQEt+eN3rcJlfVXxaVJ024EHC+rJgpHN4Y5m1UhwcXr3hMHx
KtAbGdhutrnL4MR1LoQNgfAKVIeY3XgDercEFMk0sSRjTqZWw4ic/CKFagx7dUkv
bgnG9iP+FHtS5O9DmorVjoO3kqOewNAVx1Pn3L5xIk4Ra2e98mMDmW9Y6KpCYa4f
zwsYJuKLQABcG+SDmnH2Qb0SFq06Hayft77Kgtg013FbxkCtuEDDZCjMHI4O3Lhs
oPwtkemW9y08uoaeoHbGVL4dQ/qz/ut9I7qGEG3UTTAgCCp6q1eHpph7I5GW0iZQ
WnRe9QJz9B7ke28HUkeeOMwEtX7tfX7XdjCMAq339xp3jFQ6S5OFDeeES6nh9M7H
AZTEt1uZlJWj4GySqGRW1Bi111PGbo6DA0rHEsbDg0FpHzwO7skcvfJEdwbXauUm
5frhMo81jtC2d4W0nY7AIVHz/im6eE2lZUk0+JQH+bQS1qs4vIl4u1o3kgkts/2H
k9cy+L5FFz+/oafeQ69Mcshl6e2m7e6fpw6mhDWrAwXFOkPlTjISfsqGEVaDf5zM
84EPc4B6S0vpwKlnhwv+caXuxZHIBK0RjVFXjU/rXRe/deMODDzdr93FJGX+BwEw
8yes69M6T3RaefuKVirpz5siFldTar4zZKvn6Ag94zirv/EHf6hiJQY6cOYdTOc1
Z7yFWNLCld6l3DKsEDpHXx9CcZOnYz1/IPZO+UnIsbCaY+PrPTvoIG493F2tdIu6
tDZnJW8oFoCYJZO1MmKg/dnsHFVzjhkj8hd820AhsSz7H5mItoLWQOE59xJDR04G
1/q6+rXoof9QAFgeAke/LYdURsf6c/GE9duMZLbKsz3Ber7IqsYVxf+lhL9nuEAg
ZF4QkniZCkT1ugzrLhSXIvtafID2tY/d4bIBRI0TpZCQl3XEAny+aVTCRi3GQ9Rt
BHR4hZovKutzaP3ou7rkA0/1/kA5cm0ONwD+ZCZvXO2EWaA5PwuDKxPt0Pv/pqGs
/U4XClGYxrrCe9sFcvFUXOQgcWNF1AuBlKWULhHKQTdlwXku448OV0NkquQzbCR/
m4BsXVNcIIemg/FPiE+wMc/yzCRZ6oxf4M9L4jStb8cKu1sTccShBMnwfAAe/2z0
j1UjLi8+KdA7dQUQ0qU3+AsQzwIV9bvnrX1JicyEj9koFWKxDkyO00x/ChSPvWqb
FUtRfvcEsr4HB8BzTdbExgV+cut/qC9QTStMWD1HcQ9KyJPh5FbfM9Jr5eZ0qea+
dx0eYPevBsxh6VJFt5S8KX/hZfrX1avRAVIlVJDEtZzhJMox8Ubfrs9xyMxcEUg5
jfOzGrm7EwYkK4i85dYKinN/CoqSLsF3uajtUHhij/ZMq9wMF7/W8uX8ZvUjdjlb
Y4pAy1QO5lFuVsTPdQ60CEPd8hTrnY/UkxwqhXvczkgDU4z+zOUCeIzoTdatDpN7
6JtRs11192Nd76lLxwLfTfJcewg6u/aCw3bLtWGyEWCEN+nNuKl8bWdiqSx4NniT
rhGsHomdnB3BsG2EmoQhrrC65G/H0siF65gUtuEDPzxsYFXtxS3e7pyPyKW5HRW0
lTmTqxgKceUThlabgPgbcY/2batuHj3f5C9zGw5yu34a2rxuSBr391HTQHc9RYkv
rbxz740cBDhvPwPz5Iy16+7z9arZzBt8rxw7YFL5DOAeg82wAUvzzA+mwVrNUl94
c7n4OAX/fPKsY/C6nkNwbsQeMU12p8/30AELaN713n2YnkiKiMI4jbfPccvUf7MG
wy3sFMHX9RFPUcA75haVDKbtSS4rjRLdG8H6lEH4+KAIXz8HS/s8+BxMXLFoEuk6
Wz/JXHayDIxHhLeCuBABjmq6jyyZQx+UL4l3TV3uCpM3d0h+COE+TsOif6cHt5Pr
xaFPpA4hepZJkSboGZpQKO52h3nmKFavpOTrPRmtDpyYnIRGW0R0mGPK/kciZH4Q
zUBMQDJUoizncNx5/tmrfpP2XwbMud+jxnc7nSubSauyTx8J4Kq7Bp4AvWHWLWrA
IFO1gj0dKAdhM0QejocI3dUww3yqhtvETyznOfk9DPGfbhM+ZvZ9gDKYWSgqJJ3X
0IC7rdHaI35YUtnU+japIgPozmN6+n9KHaYi8JyFOmRKYne3ZAJamRY4PCu2DoMz
bYERiEpl9UXRlUg/rTKQmp3R+k+KHi+YbQ+0Cpn3TR6BLcuR/nw17TseQKEDclKy
se/OH8gtKRjt+4Rjb0wI7Ktdn0JAhUaWgRK/JEH7f2G/r8qt43QzL7EDO/j+sJXb
o4eEada99TGEketCFouqgDNMuZoSEc0SOoNvDykjGzm5BwjgKwFRhP3EggIcDo37
bpcoKUczXWnvm+d2YDTON+dVaZs3+woRZZSEucewxrNNkGt3o3mvs9YZ5t+UDu30
Tf3nhSTeyLtLIkstRzoYE5fsT2E00yMLrlFrslk6axHlfPFkXNb01ZDxzGytcPfy
PR6lP9PhpV6rfSYIlNzKO3196W1nTuaaKHeWenQQOcL5FFa+xKm/daA3mxBypzIh
FHOkbq1Ecfqq6rQbL9OCUOfzBirh6k9r0/QHKoMNFt23cy0OtC2kwIHbuF776q5S
RfXma2Jt3Q8w+ayDsajKTgpzh7fwOGI2ZblHo9m2atEU8OX9D4ZXc7IjH69fwVRC
kACN4MO6sFvOA8W3nKAV8MHJ9WHQRwPqCugaEkRvxV/V3NT8kJOignC/YCfXgxBt
/sb4BPYsyrTzC/HygkFnNIDh3kno7W4aMTud8mXqoiLC8FXW1LAtGKkI36xpEf6x
XbmxxbXl6HkxewBFHbaDZPiKm+hKSwU21qJCTa1uKjGcETM8xZlBUdJJfmUFp9l/
3gVJSRgYMebohnUxn15qDWB0xn3H5dRfspXT8aitoIt3i6n6hWeZNNxc/KhoEcH3
HF2m6OqFL6C8nVNtmIpmDWMmJaL8WMioqpGWuN8+e++6mRWNhEfCqgb/CgsM0Rd6
k2DvQbDdtg3vL5GxEbD+/YHodng0v07rBLztkqNtLg0k7a8omJBfwyMyc/19W9uV
Ym1zcsmhpspjYUg8jw6g5HEmJ+yzCtchHpWNiLoxGENWd53RrA0ly+xqtqz5xwRb
A6jES+Gmd0XR3hBJW3baNFRlJv9CcKZOjPBbXHcPAFn1edD2fqZgY2zrUxCCETUi
WmDHxS8Fe7Jb3zcThSePDTy1W1f9zDnBQDC/c2sgtWZD8HakRPNUsp63G4vcxuKP
iAoRgcDA70ug4Sp02cmjVAhDP9u2H7Dp6zIOnKZwG4LBYDkQWPc4ZziBv3VRYGIt
aqEhWJYfEhN/qgouqrgNDIouZFS2a9HMbJEfrmVSy1FMKCpkj1RCc5m8HMI5PVU9
iJHMtwtpsWH/pc7PaD2JlJ65Nc8OoOzpTpmm0mou9lW5tXNlok9s1prqNCetIt9p
b0/2g0aSQfzouXlG+3ms6qVe4e31xTQdUiY5G8h2VzNviyqdyTfYQVmetXe/qr8j
lL6uXAdunQ6nnwS4I/34Fh1ip0+BLDOUKpTWxZoqZm/D6NM8nvAUTZe71N3st1RC
aZFZfedGHAGBzKoiQC0Qn8cbA86XBHLFFjtSSGaK+OSkYaEaI0c5ZFXJ+HZh1pkG
9Bn6uIzD2+y7NOYsSHvC7XZHSTlIf9nUPFUc8iK3oEut8OXY9FosL5wKZ2NsVIDL
BXscEYAeXNNxzFAjzHtGH9WsyRnkZxMU/PiRPfYv1KM7+W3MZiRBPPSHBCrNlBKD
r4An2vcNHReQBg93mpDfkRiI5nlOQa1dpbDdbckUn5OU5aAylrpcXDdC2to7/toe
TOMgEN2f2iT5XhBajaSw7s1fVIe5QZyZ1qoEJs5JuLoqHbCw4tjPNjvnOOOCYY/E
oq3EpT/Cht//tAWq8C0nwvvWdBgML+pQPvhdepK+x/ve6EfXTmxoUv2aRXjimWVl
Q8mBszdHa1IK6K59uhzAvycdVpQ7hvn2vUyIgbRieJzwwj83XATiaYOiupsNwY53
J3CdfzjYmOS8ARw0nJPLeStBx4wfKRdTm/JzvbQXh+lPXIvEdg7BvwGDZTM3q601
LzCDl3iJ2gEx61EmoezVQ/9stJFXH05DoKV9REy0rxUdRTuIed2NX4PX7Ovl+8+g
p+oAjR80YzgWZuE936d46lfsdDXrovWcNRZNdqO+N+oX6RSd5MNFHLGCkxuTFPNM
Y0WOoI3910xYfKD+3K7Q5uWYlRNQ66CM0Rc5ym6BA3Pekwyq5iSmqY+odYlvcGFg
2u9AeJDtqYlqX+DWrwp2yF0qxaMqvp8SN5MIUYZ+oC/traOSMhNq1rfLVo1wn8KO
EPHNGB7cmt2boV1BKSWmdewrTf55bMSFBSDHR7cbxnpdD4lNN1QFdcpQMderJFqZ
qMOVe7vBEqf3jnfNycRZFEceTJR4Bx2tQzR7mQLsFf7uCb9wnQlV/wTYKc1KUArV
rZld2gli9CwAVAT/RdMtAyYLICDqtdZ1Va/Vapw/tpLPkQH8jwpW6pRy578AnL8l
PzmaT6AmYHpGSSAu9FpHuvfiSSnC4fLz1xkr+Cc4t3OuYBGeX9s2LR77+4wn7SWr
tmah42ZzT6fTRQdo5XSFi1zREHbwQFtuqoHmuffo0aTUQoPb1hdKUC5D1bANd1P9
tzSxO/TD1eWsucAKVVHj4dsAXCpyE05hWhkl7lNB1G57VHLhM7Kcd3KS+qjbrnfx
iE0R9bvlJCS+ZYSEL7yB9HnKdFL+F/XsUkrXpowDJQf3YizNlFug3/eUxI4GKfZO
vdAE55lrYFwcAQeoVpsJqnLAYNKO/RYNz9WaWfd+2cL73ZSxlDJy1O4QzFlzXKD3
2qv7VExEgO1ca9e3RTdVQlgzuJBMAW6YX9Dr/uxRiDoHF0Xn2oI7NvreFpIWuCZ3
b++HRFrhlIs4B1LVIkaa8qUMxqrGqmHrtNxaq8tK5pJbiZliaVr9nHbQX4jUZZt5
moSG3ngJd3jOoBgI8JoBFFX22/JQYCnKrnUZYSRF8VNuuTxQgomKorGgfpUNbPP3
S80W5aVTQYl3deYIiQuBqgY+IBAxpkk3NWy+hsBC4cxo/oGgBmaCm3XiOj5574RX
wFU8icGfPNqkYiLqF5kd4QHO6fpG1hWIbxkveGppi/UDNmW2gW3OYkj9zJt94KQ6
nKbkwhCkoPCkgl6t+vVUer/Vu0NEXHeM4zdgqCJEe4QodklueG0uTwgT5wbr8uLF
K2G9fGXrTbLGIM3yrx+ZuP7dqjrhAoywEabaS+GGYrRcdKXWqzQCSor61yZc+uTi
7zmuh+sPx+bKYshE3nhgl++7/wyZKW3b7YzejBsi/CulDP9RpM3Wxqe1HENo6tdW
gP/gnW9tKeBuEwDW88ivExfftmBEfMAzjP9bckYX1sBMgg3k9mV2jCXLZeAtEDU1
4WvHCa1oCPYZMqnpwLTEsK/c8oA7o/tRhKv/Zs5Q08VpZN3X5XOmZA9G1R7XTdZ9
Bq+IgpRqbBHgP7uwH0MLWFqCLDDaipDG9VRKa6UAQk2XkvTxsETU3Kv/cqPHiz9F
z1W1zCyQl9bgPe6fcUJbL7GKsEyNo5wSlE2GmpdbfCPjVbpHkwEzhT39zwxVEbWm
sAE5VxAAra+y1ytBfcNkWgU2YJHCOsKm7Pq0rtqNjr2j6FYVfVlO/g0gzs5gOGvC
x+bGdaCFZY81JH0ISOqA7Nx+qP8Jd+N3cnvgzsT609Gw0PvNgXUCvQ8GrOGklsCb
9Mj4Lx11a/vH1axlHWY7zx6snk2R1LP0qTdJvCr61+LoSBJJuStifj3s0vAgPpl0
PDT6+SQypEvqrtFf0WQrfxCm680Ev0gVdpyIOVgds4FvUg/krhdjdR2NajIDKDb9
5Ld+GdIMgrE3RdkAZ46lDSsvoq30MnOuwHA0e8mxsIwo0BaqdpgAebOEcqnUjpX8
3uFPmxPYhjC7tdp4evdwkiR8/1Zlyz7IHsqGZQgXh3pO0XbbE7ZqxL+6okmHwoO5
RKG8MNIQSg2rCxTx/uLDuFaffPuBf143QQtTgi3lZj87jxV0X4c6PNH7P9b7qLMn
XhbFagorvW+l6bbGLMc/nYzo0NXCM45GK49kvkODczkNebhlitwrypk9/qQxqsV7
zAAsWiBh5OGApSILukCkzY6pCk10DevWmghybZ4ao8WLwCHW0lf5cADClYKzofpE
3oNvyHMyoQHCNC+Bxvcn2QzPgmr1iuGusXPJCl1UZGivxuReJ26TBB399xCOGLFO
31VW7RtB3xLjqrRa1Olgmiop68MOTf+xMSIdTngu02fY0GIeuij7btqcO2e1fEeu
811I9gRkvHy7uAY7cl1a8S68YZsaaF0+0bcgYkZWMT3bSN24MoIQJPM4tdQPgJxk
F/pPb8+LzVWFUL1YaTWNU2h2F/77kVDG5y1m1FWC4uI5nXS+e4Uos3E3qIbzVX0H
nUTjx7SDxws0n4MendVd8J/nh5Uf2ruhG9dXwj1Q55ugBYNzcBibKZ9q1HdboynN
fA/DJKcBeCe7P6cfGk1minWdADTwcczvQRLLaXus5Q2KCY083+7d75D9V/4PeGwi
B3d3dM1W7L6tjM0zrxBqQfKxKrtFnHtng4IL660yZFpvCwJwNyjHfL2nGrhWvrKA
ToYC5PEDTI3wNBESIIQEp1rrH3415dnvKjQGeTtVl1UmbgYNyvy0wP2qNyTlgk98
r81ghKeBq9l4pP+JCLrPhAhB0WtsGF4tBNmqS67WAC6nkUUJHCzs8/64UBTAZ2oV
HaLXEEkDS/KLTSoeWXnvGZEI6ktTj7ZEI7uA5+ff1kUdo5LEzqM6WbDvmC1Tf9xa
P++JAKgCEJmXNhxwsWSEsTRsHbr8ML0nFRCiY4BWbbxfRSUoHDOpG0grKXu3ebk3
HHG1xmrvFufeXD8VmvJU/T5aDJBe4lCYqX+97hyauD5OZuG0U8lBlg0QLy7i3msx
nSmoK/jlhndt5gjih5aE0yM+G+GIu1u7eSIsBRk5vPB7d/YFNJKClJscXfXUpE/B
bnnqo8UveVbK6ago4FUE39O+8/55WKattwQYSBAnOoszb1hKYCAPvjBM6ppnwiDU
vOvaW42m+exs34inq63wvKMUgq85gradwFQcwNI+wob/d5x5bZwuXau9hNayTmvH
r1i1Ew8PtgcS3A5UazZusoL5FanWJipsSP+LsN8w7y5fRRUkekZiLsQoMN5pEj9N
Ua8QrwsKv/0afDYkukQx6ts3BVQpd3B/dGMmUggwWqO8LTItDHVJDRBoqog8fuTQ
oNq+zAjX60qry4xCtLL4Al5qFpoG0a9IXPGcLnSouLt3Frer2D0loahYUZG0aV9g
pvYfFhUDFziOX+uiFNdAgPfCdvHG9aaYqv+vpeg3GGY32FeKGRzqtNuJNRKNfYmT
/ZaoVUF4qKKFG031se4ESTMC3OWw3lmyFJ4G1y7OJseADIo/H7KzO1LfCBwSSj2L
NikCtRs/lhmaDMANxhf38Y11C2kHh3VLMcuMOzcUqRr84P1SLyw1eS2yGLBEOZPz
zMb+t5vyDxGJNQ9de4tuP2by+f0MdRrvL6v6EcoK9BMphmh8xcwngPpHOL0eA7uB
7G+5gkhuUT2NMJW/wDDosod3Ivv3jk4DhV/fWCoUmu4I3a+o8IAnJ0d5uciuzFzx
F/SSHgcn32RaZPRfozaPxIdZkhon4j2/YCEHk8F5X3X/YVdVTZyRDNcTD0M8L7K1
XNdNT0qx196q7/XvhpJJ6EB07BZKD7tCA8EEchmM52zryAsQ76FRiGbJlFs2fTn/
CDxV7IK3YexMUkD0wnQyzpdCg+oXyNS7ak5K4x6h6xIfONy6agYrwvWEEyJbxBvb
jex3xzN9R/hIAkBkONaE7hx/JCPGCWR+Y6BK7mQbHt+4ktZOi0rs4KvDmVFFsTde
GDjOe0M9Vh5Z7OHMrSmdqXY+FXevoskcxEVm2FF9Bokr/SPU25xJvGEUhF1cUIEy
5gqes61flLlin0MMbtkiiQE/GnbbRBeKKO3gXmTG0MhK1utcB/rVet92KG94972c
X6m0xBBgZFuIXC44WRKxhhf64V/Dnah0G2Tctvlp6gFUWqp70EiM91Z+H4BribN1
54szlc9+I/NVUW8Hxh5sSpG9quBIBCQbOm1veQbhw1BDKLlw181Z8L6NwLNmX8qJ
VB2ILEE1HA+RXZ6eoe2C+lCSj3UWEd1CY8SgNdPFKHD0sOu1rLq7/ZtMHIle8sbV
mmJJDn2plnd+xNwSjk7o7A38tDZFtQT64GGWY1km06cwzhZ1Bd2C5jocy0yLhNFm
2UhtSnW+glajjzPHE2SXovt38V+Hzui3qg1WbLsrTvd3h/gYer9Xnu389Ki1fY76
qJO+vv9UZADOxc7itnoYewwdunyPT5sUuWMA4pnEcbnrKClZo9IIPT9NMzgiVhYF
StXQwROsTVxbMYJDGC0SaRE62x219/XTeA9YdBBJch23kwBwyNTQM9eZpu0ue56L
lThu/0vATftt6XXrgep7lu765qX67ccQ8DQnBmGWFEgzveFxD9vLqpFaUkqqwoBv
FjTrEdROr8FMzn9okUzEeh548OkDWp7ymqRC7bqurbRlGEiNkDtZ5V5gCm9NaEDQ
A3nL3ewFoLQe5fhEYRuI+d6M/eb3GsfzKRpq2avq+vdtf3mR8/9kL0+B304sr9wD
eTn891mQZcJPM7j/niFhARCTK5+EHG9EOLlE+bhxOorSR0A669geP0AntU98bXtL
9DkT8Hplj3RiIOideCvPgJQ06dAl5fd4lnKBRWYIYhpDDDAJ+XYs7eyk53EfSwcX
oxya9e3LBpb1ijfxVGUW5M1bcoX1NBSMPUy0kqriHAkWtvX2AIQ1K0ygTgZlmmjm
CrMSjgYLGd24MTjUGuXMSrqZMzxF3YkN9rc+F7nVtceiPyJumdPBW4uNWhV56Fh/
YQlAcBpSRzgPkQLWhXWhRiPr8GsAaMrSCdujhdWVWHvdywwbHKNae/5D7GfzjvxV
ufg8e5AeZ37cXocjhtsrddxnoNIseAxk5vjUm41ob+9tSpAL0aV92uC1UGW28rqj
NdwrBiR8O2z7qEOtklFYiZSL1oPxud3DwIvTacqxmb8mxHDlmpLjWovaxXfoTLZL
xyWGbhdros5Q9RMQIkjT4jFGkLUEm7gZ8nJBoPU0XJgqLQnIAjtO1m9LCEw67ML4
FXiwUZobiX4A9TeHEVLM/6B7A35LcNXd/AJXvq2ZprUv/fWEf5cWnPZUFgz1+0Sx
Lz5pKeYSDwrdSjEr0/iddxuaFc/5XnsmsYcEWIkK+tKCZ5JqLxnUB0KEVCPSjqKQ
4r0BRePzwAiRaUz+vJRvRAzSM56JadEHJfCW+W6nfF2cGKKGP9BErX1YXf4roRzG
uMHt16McAPmlJT4hPvrmxUZW214A+6yxh5IdFVU7zjuLzkmz3MT/LMT7TPagr4xj
IEyU7r6s8D7Msl4/Kufy31Wvu4qFDn55tRM1uSsVkQSc++7Xf2fc2CFQkj0I/3V6
Jf6I/vrkc/Iz7QU8V+Xnw+NII5U47QirY6r4hKhyMcFAWskn2KCzCE/NZUwJywRM
yeq5ROKJbuQ/H/Ywru3PgXM/wRELdNA3pL31wsO/c2nR8wAOFEmuK7vgYXBWkACa
qDms4EmRF43zLa/uaigmRWx/czCOB4V8d46F6Ok3ybYBlXm1AJ3SRi1exOd5iLAX
1J6nce30piaOPgf7OTl8oBEzhXre4o5VaP1lSvFhovvrU+r7cSxj/11PLTja8rLo
QV71bA+wUZY6JEQhzpLFFZ0kkGrH+I45H/0y6+TpDKL9ep2GAXetoCUARrJv1XDs
NId+6hkTKMIXH4leDnMnKNhpZcsVPPotvGLwET9Q/DF4FlUOBD9rSBypBwNjk4ME
uNezj4Qa98iuSZjDcSKpBJiNg4UZvZVUnJzZOZoAC70r1O5vPVrfrSOaLFIbwO65
lZnwpErG57Wfv58YyziRKSIZhYhfMrCBRVJo13gw2FxcRLb60JTLFsMaXhImEBEk
lE06JfI12LK8JM1wi3KnjaN9IIAjDNUPjSCyQAvwZWHin0MRNHbYAiGxpSGdTv0r
wwp+O3CH4rF5970mXnj8aA3BPqWjmTaa2C3t+3+DEFeRGgsnuZKPXT9drU72Dm/O
2xUu/FrTqhgwT88ofrfNFbixh43BeDvxoHWPTW+0cF1QvBMJ5N1SlpAyRNHmMS2O
/KAN7/nFMm9VpJ20UlOgpVPdq7ei4HF92ubjTaYIpFIk/e02xypypEKE3xb0jLf9
E2FGaBaFhqgdsjdRHVWydNkQyK+JmkK/Ot6cQuuFsvYvDxoEICfieBV+fd2L2C5i
gWf12fvRSJEnIU0CyBclpzDydwqvY/jxI6BiFOTcBmSToiIqJzeu1I6ag/VVC64U
Rv+u2jQCm5X54CBWaW/kuszLubLbvHhTFLN7Ytpy+UOF1CwC5ALjyV0FrmcmOvHv
5xX3R2vkTGaAttIEQp3g6boPo1dQ3Tb9uYhfWYwpxhAm+Rlb1sk54fXsh5bWFS5r
UspZPPYaJRXiCGlUeTYGV/Qok/dXhrrRpw3q5pyKekl7nmchY767J+jvIMlbcT6S
LpKFVI/kz7KBhLeOymjlgC9fyHe6Z8fOICndPHraZ9MMv3aTpcZJk75/z/k//06/
rgKv/fZBm/UERc5PeguZgbOvPyIzDIWwFKOTlnFDIHV3Jsa3ANFZFS4AeMT0yTV+
Vp6jcuJ+ZBIYUzPiYEEOfPtMu6IVqFHK81Sd61aYFWsJb8vpWYKUbuFiwv8vTrQq
jbBgJDQY5W1PH05LPuPtmKntTN6Dd0sy+8LFeyLQE9BzYZsLhRe9/9FLowlz2ryE
EdQEaO7FH8uIbB/CY+8aA7FaF2k4RrvznJRwHdHToyKPOaKYdsm05DE3tSWW2P9S
6xwasZv3wqFhOwjculNr9PzALBbRWzBwzhpluKpS/tBLWE+lq9rFpJZWyLSB1sN/
5PjlCv9m3PiWDHbqAl1JuOdLx8J7P+VCGl4UsPgV2bDvrEZAlv+85rK/Zysr+kd9
7N6cwBKeeIo4YsY49KQdaeotU2w3FwUiDtJloRNzLyBIa97wrm/elyN851TycAh9
JGHMq9RMhDoWTPlTm0ajU+jsxCwTHg1LvgD3858CyhqfQxXfJBlkOE39o+ojkrXH
T/waoBqBegZy5+2BdkTU+fhQ8IuDSvyqMWCHtKGCOQpIj/K9JUK3h475XBI+w/0h
5pS3bCTDS8GBW3Sm9DieqwboZAbX8GH4/+R2gNQDUoJTvvpVMhXPVrDj7Lx6Ik/U
UUEKEKjKWJrHYbDv2wDku066HoAL5O7wRuLP9cve0sT3spb4XJt0g7qPfxJEAqTG
MFxTfqM+46nU6Pzo5QW9YVoXBGSd2I+szfdFeSSNz9FgkLSLPXFAeWp/QWXh6CfO
2hvCAoJklvt77aRpNp5OmsRvLpJ6rjZbTYW5QoS5YkabPqOBIA50k9xFeWMTaq9v
35kOkmVT7cKpIQzXD/RdaBM0cg1GulQTyLXAQsixAwb7DxySnX0TNAJ9Pp/fWAUF
v6M/ZegLewtbsU0odJs9sE2KTHJKzqxkowBc3TBsXSVU8ZhAJbulDzfE5s56kNvw
yJqHaciN+CZABqeSDrGUBq80ifNgNkvbCJZ5bIVHE4n6IbiZrN/1UpdwqB6pWxtF
03ibtWy/bSqS8E7/oMqbbow5GH+pzW00FJFI/gUhouGFp0OplUi2A+8DecAddeuc
x6S7p7X75K/SK3w0JzQMq4eo1FA7JJAZlpxQ4WM1uhKD8v3sBFhu/TcIBwFyGB7R
G1i0maX9AN/4Lbejo9RttHcNXjQdsM0mFyTBUd9Fr+S9OlX8nK77pOW0xNSkQomS
aX65oWLPhuTzOjnvxqhfHmw6SldLpwvylBwuXxJF7a5VwDL5CUp/bu9L5gSHdxdE
Yd6tTfMc+oXumIRO3PmcDL6AOLrQk2ivThlZaEw4AnqTE+a7EbWWJJ+SRL9j+z6N
akh/27TdcnAu7Xc0cOtv3xfEq61IaFENu+hwTBrZye/qwcOqwXF+8/uw9QgjKvd8
to99/uwfgBVACT0eCG86VM0pRnUS6bI8fitqjb52A/xB58LgdmJrgmGGjUUP4hQF
0P8/pmb/yP0aw7lt92Hu59HVIalKmtuDzuUr7H0w1yabRkSqbzNYhPSXvJTPTjnt
/jM/Cx0cncynUHjIG3923ScXkuUWM+jPAdhxvGkTJDp06n7dBOPdiaAeH9lpWLTU
o0KWSmUkq2dTbYEpXLGPlmuEuRECYEX12hNd8Ep/TrB2cZED1j/6NqsClHrz1Pcd
qJqaypT+kHCqo7Pkw+0dh+w7hqX9m1qkxHcZMLBMv+9HsXZwKBmaaD9pp1gDfst5
aLa/VT6dNT3uFXgD9L9HtTB7vTWqMfVr3ObfvCa+BK5AZD8TrsHY5WEgYN2d4yhK
spZMizek2wbmdCybiJ/AHJTr4NV7B8EAobMv78i2eXudXVpKRnx1Npmnk1qQZ+Ck
AwxsKMjc8iSAYsvaIj8d4xVA27W3mQDonZM4zD8EHFYkD93UguOmePOTAf7lBGIt
tEIL02haPNNPZglpKgb6JxMwFLKyspwvtIPbjAXIj+Fkm6QYT1tMhSo2mI8dhRKN
RsLf0E1Fedg1pTzGpqC7es+3XTAC/Ypc9kGe92XfPTZG0KmxqCoR7wV+u8yuM8ti
3ewyIjeMsSY6MkiN8ABU+mQOFgIYjGWUGDelohY4FdR0mfytBcbN0KPTIgakV+UA
+A6y3q4kIVaqLcHFHAl9eadaIt/qvht0Cy0Fs1HYxd8JXQrSXBp2weOEBY5Bm3R/
knRnfTQwe8EM0l8JE3mCajhbeW0kMTQlZ7Q3TjQRkw3pU8vXyIhYgZNxGGzlUkTQ
m5rHg9jsfnY1l3Pt1eTdJHJ3Aew4EiktKRd6w3DL/m3R4Qxo/WNu0ZJGoQDRIjvG
ebcCJdp5mHcXEdbrJzOPXKDSKFufeBB5VM7cPgYqlCdw7hdc176BlGuxMLnzYd9E
/5Spl6q9mXNEn+1u0Pk0vPzj9qjvXzFbTEp8Ne5XCSPD9npCFjEBIkd+ZTF8aBWE
/vJG7c00c3Ok8T4P+waftno6dzrSpWkb6WqDyzPPYSN6wJSnBZyBxDjqCMKWhnHU
3Lhn0VYG+/3P624O4Qft9zx3WaE7ngvHAk3YQRvNk8tlCgCFIj+aZesNOMUstzRo
f083uA7dZ6hapegs34fU9m/2MYZDRzNXzRKS3QGb7Dr88nMCwbDHC2IhLYDa84Ug
BYqA9szyYQRNmy0j89rvzM72E4n/wZzLZ4Db9gW7KG8KHtK0BjlDS3Vj8GWe3M1t
jjm0Nsj7U8/qM99Ol8ed+8HPtIF/NwfoABBVApWTbGYU6XrYE5TWCIoD2Z/fwVaU
yM0ehVwG0YjjEKQGe9uPB/AwukXJRyQKliKh+s61NPAL46smrcBVIQQMQG2sPENT
S+M4dAR+348xiocd0QK6VarL9RtbEj80Fprln7Mt3MZDa5y5LY8otfAax13e1mr/
ehL4B6SjKCf+oVE1BC80jhBQPeK4IRIbTTX5ldsc+DY8x5Me9ZurMK0o8xsmtC/G
giDmuUS1AJEqDclomzy9yXJuxjmLU7rcc8Bw/5QTVKZzMrU/yUAcMm600/PHEFFH
Tv5x1/N0GmrJvznO4MEHcTgz8WK4/7OZqmPMMbUv9WuYyvNBT+9/3ca5G9T3HS6B
1nirIwPF2y8m72QLeX6fT3zEYhSriEs9RrgwXVQghDTUXlAZZyBd70Wqx1wxvJZP
B5Q9gdpIt1luCD8FnXV2hd0nddUw/dOtdwnP3p7giUYDOWIb0uxGNQGVvZpHSG90
ke+TXc+G7N2dBz5g7m9o05YaA/MX6qTgK91Eef7eZnqRzM/gNSmhDvyWQMMhD3NA
ahhR6pkrxJbErKUy46alSDK7l+vZXULLmnKiiSA4++iayZ4ON1Yy5F0UvvCFwofO
S//1Yiv7dVB+bqbldj/VhzKHeqte4wO4KMjWShcgzO62Vg3vLND8K2NRECBh8JWE
csFTD4W7/6batzOAij+6ktFVSh4dl1lBLko67l3F1f+3HoQSyfyoKZCK6B3D06UM
9AJZMhl+/mtRDnlQpWtlhi+tbDdc26fC8QMX8bzvpvrXrQrNQ8GPno3bF5hK8d43
C37cy7bFznyoEvSAQggr3Kt8YuBdPv01ZvoOxdZ0ItgqlGPi+jGtiRrallLBlAaa
Kpt78Y703huAR6DfLUDBNuBG08ZAYPBFEsXeX4DPr+3asHhQDqw2V7Gmp1Xus9sb
HU7N/Q37oFMMzvWQEjHjpbi67TRJzKoO8PQ6oifw77+IaBG5TgNSUA184PkosxIn
29zEWy2Bu+f7bXcnftI73M1M5SHswlbHcXgYfxN0/tdwJ54vxY+0pyCVQDx3Kurc
XgoL4u3LFtwHm0iwITnUqH+NrnWPNVBTv5sg2tKmJuz4HHsYv29wRpX/OlOLa/+E
eIabaBifiLvd6yotZrdBk+0RxpVyeHU+v/QYjJeXhGpF3sx66BeljReoFb3EOf4w
s8K0ruoaV6tg++ZQVzYHXnrkx9tOQ8ZaB0v2dE1z1bvOVMAVneFyrI9wgojQSW5h
lzPv4Sb+vm6vDfTzbE19EGYIxo8/GiAs4gjIolVbpUj8i3CEyqbCcpG3m/by7Au0
s/rjZ7PWu9HB5orKXIZsbLpGRWdzfFoDzAmwRGSDcj3vymOdo1SDCP/Jszk9tAIP
J58NJt/5LNy/JzB6yraWvZ2NCqVSEqeBY6jSsDCUhV7FXQEDhlvhalS9qmQQsixT
XcRM+NdfCpNExSOc3FBI2PvnOZ3VdhUMXbExBpmSsWjtDmxPMTdOOYL2KKVrJNtB
ifz/b8judEKoAb50OGy3+7NzDZrkiiKFXMn4l1kfhp1WxMEJkQKUcAK6rsfqNX8w
RId5dm5IgjhI+Afh0KPNvseGFhbB+Ilz3Ep/zb7SgSWMmYPU51JAR0yJw8mN+Ha8
v5+8Tp7q1MCC65967QcabX+b21h1/lTMeVcFKWWt5NI4wZQFE8U/7RUcQ6Huli+F
abxv1Z86lErvDhl1gYJctuwtYHJF36ZY4s7YBWDQPjLc5XqdzSP5srABH4aR5CPM
anK0ijaXPh1GM1QhA3Pdmua2hceAfs8B7uAn8ylh2lIT2yDjQ9rqxIAR11zlf/S9
By4fWG7KvqUGr/WdareBExS0Sm1ouTYZ91PffSaRCmj3JPMvc/f28FYfuAeW0Tpy
T8PIRWAugRTwHR0USWqN9f+sHmg9R302gaykcsXcXsJsnTdBsvtmKoMv1IXupAdG
GriDPnS95hoGg5b/XGHTlNb/AYyctUicGjR6VHLBICsPgcERui/y1/358X9fPxFg
ySfSJJaZOYCWl944d8m2yYntfUqFWzKqNNDrmC889WVHUE3QmKsWM+aABrpLVbfS
Z4hN1Gh4XeTmfULECBa+1UKw2QTU+kT28WhMI9utCKlVuuJUMeGVSX0PTCgmlto0
Onq2ViosSCl6v5T2w3nACK4LpqXeHBH4NDaivz6GE30BCC6CbZrdAbHzjsI340Qr
IH55ll9tB/k8TvNBwE5EF1OV63hrjS1IYo8H8vxns9uALQ/87UKe45K3putetW7L
hAZnZ1hEICcXb/gTrkpOGjqqIEVjxBhmlQ42uMaAWhkIvqnYBQFH3miUpQnpd/s2
fG6as953TvYnh9eH+GxpujoBz5ZNlfWFuEPA7eCU/kneF9fD9Moz0OYmJgID86q6
P1FBLR6DtDMLw/S9/KWxEE9mjYBY67/jr3mzoDd9DMmWHZMjO3xWn6OpMLZqZSs+
AMyWtybWhtEwRnJlIBS/sv7ryEFsA6vHDKMDpUOG+swixCP9cmc7E7wX6fqz9VEw
2ILolVVf78H6UbpsvEO7D9zn7wKiONYawrHwkejDb34+sc4dKQF/mjgvoWs9qNyH
MGQg/pw7cHH+4fU/ZOiT/CbnbJcPDD4tdXjyMf7aJa7pdw9AMXvQCaa0WeTsXtmq
glYpBYddOopFwmTcvq/8GeYXR/UjeP+mFljtq0shoLyc7QYg5uyLLLPOATK74HiV
TrYfcO50mahyQTQ+92+rwgvp1YUpNdWvozn3zo1GNTxbAIwA8q3Ktx9S6iPGm/1W
6WgznUuZZl+LJzB+9XUDJz+GxlMKMrdggzwoJecc4pb6LqJ1ISZVuYmQeoNZwERe
kdijOrKK923vlxVRRN18gXQY1Z9qbyG2HhD/FuMJj3ls4pzLz6qF8Y6tDJm8laBE
lTZmxIngq/wTaoHuVGQg+zkpOQLVjSYz+nSGUQ8HyxmnY6DzQbc6eWAVIlgt+avY
WQwShRKiusWPVmjCa7AI+rj8+WiV0943DJxG1IlZxRaxYwYLLFs1sUIQLrDmSBJ8
Mp03M16P6a0HRR7JWqCdX5Nkoj0ync47HniByjE74mZez9r1hqeUuARQ9jygQ+yC
DgArJTOPQGcGDk+ArIu00D/j23pAz1r/ALe0W7jImoakFPLUjkveZz9RHvX6IdQB
5MR82swWO6hI758p3FmBnuJj1xDTdf6SFlqoDWtgw8EMU+8RQIJOUJ4k09fCMJDA
syZAPIJfNZJFeUClUZsjEoF/fbNQ7ewhgvldPoTJ7NopdDFDpAGRBK3kt2N/wynm
JliJFBildTptJxhVXXLJ5KUrpxbElSaNAE99WbsKwyvedyYS9/VvzuimkSY5vZZp
J7KZoyxz5vehD4i71ryJx5/k4xwqSD7ap9+ikd1KUYtRdglwpVSIij911234HTmS
3LCMirbmMGNi/XmO1F3l4U2NMdu6lF+EQVe0uFG4yRgOdMlke+EWtPOmoLOcM46p
T1KDDnWdVlV/XxCqrt7w3oyBLQFuFVcbL/N1vqtZFbzYcLXCjj2oc8+1Remi+1Qf
XncfLncmDBBckNRITQjfSboYj5lEQlVgDupoGbYfJL10wMwn2bILAPoEj1kSBwiv
JKWx7UkBaw7XqVCFABFZMyaFL7C6YW9Akw+Sp/iBVxgnhmvIdtmBQjLOb41UBK8A
UoSY4DUHL6+eniMQsakTMTQVkqwfi8HYgfxflFg9ExASvdOzG4L1TFmWK4vo3D9/
jBhqlJ+M5zrew/3N+6Xs84ZT/23QE9itb+r3b6f0t87aCjmCWE+CWdKXOedjFkzW
Xl8NxvwXKV+dgWyin7UlRL5HLb8AyLyilUMV5dQ5q0YJhvWkufj7fUIyvgSXgPRT
dDiuxiZNzOdZOXxAuy73nGI21bN7blxZR2za8BRHkgracSwvwQR23qZBU7t6fps2
pD2wj7A87sZ+pdEHrgOOfb1eTq3hj3xWxri0kHprtNG2eNXGkztneFqkAlQhwLnf
KTabUYhd+S4cC3XNX9HKpbBvqI6/NVG3SZm2Fhc7SNg9WxHpL3K85BjEJbS7pZ0f
sKEjodPLMb8xRPpgNkkKFO2SXMIEqHX+Qbg5WpWm+doU2lTnAgF4hJ0WctZjz8N2
Sq3obqh2FIbmoYKLo1hOTVmrvZvTnFsTiN+tCQGi5GeW1eR/a/mb9IzPglaYdMsV
skSWQiRgArOGUEV/skggJpSUpRWZMsIX9ffgs+8RMjPv0YKoVEJUvU3cjQfVB9gI
Pfz7HgSAYP1Fooemu8A/TbTm4EhNohydKmTWZ0l7pF57UnNuqvPyaQPlU+ZoAV9p
vVyfczEdN7K7GpcDk/2tsNXX+vOigi0Udtz8HJ8KIE+imC5sxi9PMlVuv7aYwSTn
5EVMClVIZ73E2HJ13jE624M6mrOvxX90qjV2Y07Ffq1VG5Mhm/TrHwEduFiYLfdE
QDC2/WmPH/WMc56w2/E+OzYzuumpixakeDED8UldhTYQ2cPNJ7D9jLMTlYfsdzN5
BTvV73KtGmWd0ROEoKcT6mzws37V+ZjEbjKfBYCJNSBxRceWsCA8/nchJOcn7ZUf
x5crqBelJuViiakPVZNR5inN3mIGUlvRXpJUjUCG5INF+Y1WXNzGLyLM1nYnG5yx
0nsaoGLq7B+KkEPbQAr8jEmj+FKWQtkh5wa+esHboqfNnYF8qOE6wfr6YRpMDMhZ
s6pU0nYe4xRNRXbtRi6S7zjcPSiC6ZGm4sZqkplZJTGOnSlAYh8uSB49ojN/YYfq
Q2tyevgzvv/qW4m1H4phI/sjIBCgRScBsmmAyk2WZ6mipdqLWni6g7G276VnSqy9
tfkNFjWuR8KJ1Ha8s2q1Bd1n6jMHSHrgErKJHooiUKrzFIpenqtnxdRO//gZSRMI
9I/5NQKPb3YrJHw5gBU6Fm3uK0pPH052R1aVWXcFH016DC5Q1PNWtOxtjKg6u3L6
2aW3JscA1cSOHiLhw6AryByMPeZ5w/RI+K/sw3ufkYCSYxeL4G8pDOKZdV42KlpP
cL2z62GIpubRk04qVYg3b8xmD/pxP3fnY/hLBIos2u63Xbrj9jDJIAxALPvnnEr8
X1ul4G4sgq9RbC81+aUE5m5bwK3x5gqFLqnJgJwRyGj4mjfNV1B1G/uVgJpQAtMM
fdHyKL1X1KcudUKOZoSuGQFcSZheNQIkq2z/V7gZeB/zzhzca5MxZP+6lh7ljqQ6
1sFfpZlrcMkGP1gTFbOh2FtU9pCpisIX9VMdhdOjtyoxBlV/1MsXJxfCZxCRbe/J
ZxG/g3zxN/2WeaJNURXcDRhgvPv4Mk4IutQ2/mDVQsTz7TOpXhpq5Lyv0TXLHNev
vaehUc+PwPmLhyCwCNVw9X0DNPQIGwwEpkWtNug+rE3boi/m8E1RV7WzpXGT12k8
vM1I8ctSMkwKjRp993sjeiNQGJJ83pwGYjZEnCajBGSW+l/ZLlatIAfrojWDbP7J
U0dxLg5uJH9O9ZPL1v0svfdnQXMyJcYf54bgOaKLTTwaAjVUJVATqerSb1l0J6NO
u4kVfqWVMJyKyL+KmcvAFbY2nHGU31IdzKT2WkAr8A7NdwNkp/nbIFCIymsIBQth
4fNxpRyF1gQP6bo8G09nJ4qF4d0aHULfqQDQGLtFFiPIyP4skKOIsO6Q1LvBshUs
C3MPNsE7pnRsQ1FO1eFhFu0y9nMWy/dJVxvmK36cuq6+2/Qa9fTwZ/C5uaMkLLrb
yhlLh5qNOvtvfdJa31y+Q8ygRxQb2IddW+xnVYFvIKCfkHvR/Qlwxu2gMNEF2Z6+
jHkkQnhs+wKpDD0MgEf5som+BhJ2NGMWJwafbPJwmrkNeuRRTmG+H08ai2C4EAmO
+idRPpE8DG2jwjgg8W2AyPX+CTaoyFZfLITl4IyPy4Q8A0/eZ4C6Smv3WDYTde09
x50YYIGdIY991JL2M/MHap8QZHH1Rys6WpOP1uB6jsW01f53AgB3GKDzawspx/7o
7mNENpW3GxGOesex3TuTGxhNTjxH9oU7ZE52d4caoylKNfKIEqM5L9GmvNK2+naU
X4pA4o9Z+Yajo1gs9EDCHj/sxuPx60zld6bsVkOZTeLdAlf5kgQeMi6U3qYDqUpe
IyWombTEZ/b2tCj6SgAglm/gUhTjg0+jkPjRQAIjcVdlJVH+Goi3q5HxgLRFPUKi
k9FY9XphFUrjjIbh+JqdpG26zkcnlHe7ZsoaBJLiBX+xi9U/JyEsWpJ1A7E0YdJ+
XSwM5FY1dVAqtnlB2ReT2P6xvhbeFzbmA0aQ+9PPATjLV3QrQmM/zJjUrZVeHMQk
k5SDdK9AzOgW0H4bENkvaWse3f9yN+rC4x6v37cGkJPJ1zsALZhEMeHeSi1R/zIj
J7XEw3fheH8byLe1/BqAP+m5LIucTOFJu4jT2V5yTq2f66mMVRFoJP03+K27Qcbt
prPDyRyMJX/DLFfumR4JMFNtTfuRl5Ipq5XGAgJzb+7d4oEf4kHgy1tJJwMB8D1d
YMd8wfz8YjZyBswoxk1rK9BO11szGWWilFM7U8vmJn09FlZsXdqUtIWI8IdLc5+D
pCPijVjoAqgvqxumay1mOjOPKWSity8U/39TvtQ3VXwlzMmoGGaU8nFTxQQof43f
omUxJzuBxB69AMAOLywd0NDvJjSJAyyEQUdNsh66iYy6CaQEzyOj4AdTcvdPfWHd
8yX+nJdhTLvXGybjG3ZwDsmnANX+ENPBKwwSo5Kj+HPFc29hvjCbwOR1ldPDMHLx
QByrJW9Cn3XOBsBCGwHenETzCoIeDgYK0JLBYpcrxhGFxbtxKKeU/gDAa74/ALuk
tksaV0tR8eRiJs9J74jov0UEeSe6S4jFbbhoiy+xoozhjoOXtzte8AlyVzEqWZRA
N0EZLSI6Yu1asFsucM60w+5WQ5PpKqkw0+syltQOBibDrBcWvAXCAbq1c5m5Ejiz
U7DgnWZwqiZvwN7wQXruGdCDyaRFYZXxZEInaOsPELcT/rYysLVb5kSl3uIQ0SMn
GmgUXquykcUrXS6wm/upI3ZTSTSWfml2wVU7wUCERZmumpU9B6WHeV70yaHl39w2
pT4a33aSVHFYb6arqtEIdBxPLNPyiAYCamFKHgU4q6xJZCOWsB95O+e4rtGiGgVQ
Kwv1zjeN++xetUqNqBKpQSilwmEXvmNnHmACodDrJ8X62q+yveEMkbRToXKwTHnp
/lsuGVzZ4XUdVI1hmbVFqETQ1ly3pgQWOzWx939+Am7Y9jMCZ8Tm0PsC19V9qOYv
+88KIL1XaUqMbHAAJaAIru7qTfjPYO6mPoKu/7Mo5O1/+XJj7IXuG90JrJbd9KqX
RKlCvFgFEsV5ioVag0FQBfYF+JflzabUauxvQGb+OojCameV31QZ39roPIF/XxGM
+hL+6Nb0HhS7Wj/kRwHx30s/iJ9nWPkSMvuWTBvhUV3z1EVxBE4yGGj+skJPNUJ0
zeO4vksYdsAFvw+VCULhQd4urh0MvqsIqCHJZdVG6pn0BYWVL7XEyftSizbFxdX1
3tg7+TDuBLY/KsyPdU8j0H6HmNRI6i5smW7G+sPHHab003y1CHH/956SvViNF8rK
yRhsnbmzqJdQX7e+PkMApxk7yB+VpQVU5zmMn9ZRtcbSpH6Po3qbatt1QZfDPTii
Pa4xt2VRSVPOHe0hgEZuz3g0W8ZMeP2Hk07q2s0OrmMp9J/X3f6fg2oHqxlLySf+
eoq4Q7eejhu8NWTEkeGtP5Su+PrSa5PX458tnzXyYwIo3dZ0geGx2vDgFv4ZmZOv
LSISDDM9jJOMW+muiu2SIuIWClaKd2eNkSPgGjrf3Rl1gAK2sXsWtjigbQ9FaMp+
LQFaTDUPD4ufiXZeIZV/BQBmqdgB/y3XngGqCcvmkCu9YKblz6H2Hz7RxFkLWP/V
tz77MQ1zVdkja65jWVCQOaPHUnH9iWMjSfL+2Wq+SU3WwqZxtKczk9VMYf8LmS1S
sPuuY011k59ymrFxFrmpCnRDnRGkAVqppAXy8EkHrPc5qv8nB7jQnl1aKBnLRGjx
57uZM4YI83rlHgrXDarM4HoOqMbZeowdoTKibGbTYEWFoXe+drpXmJ1GM7LPozY4
MXEt+ofDfYbcE4sImfTx2x9fHKbclob4Kmyxs8K9P5dFB1V04TY99L+m5Od4ncxW
Ufysrij7Gsd1rlL2C8y3RZqKFC83GJeKrYucGTRj4vf2eG5kCozb48fVshKpy/CA
f2wW0i5CM2NNdnnwa+1sDvCVntlcKCEGXpUayBTYnfJE3mVqaimPCskrTja05Yas
Zc34R+kqQViRiLN/sOljFzZ/hEPj3NTpStxIidV2xEZRBvsT1Csx+M6T30/AZKcK
Ug9CLYu3IU8A67CCBbcrQjWEoHWP2jlisWgPV+k1krmKujF1cVifhb6cE0nQeXm+
Pgjh7QHPWH4EbS6I0+EuCA5OUfrXi6oDOvcYYak64eSOWssK4ETL1H+AR+bEYUaa
4YpV+xRiAQvU/EAgICg3b7dzfenQF9VZT6pq+iAWGlDm+wRkUwYzeptW8f5qTMTC
WX0WBWf2UYI4rSqQkNrElnP6dAPlQf/dWoZamBu9kOIOg5g9K52beFtVSVYWaNAx
7HEUiglmEuOerpT4w7wqKmF+kqU3YqZXkHQC3KTJB1AbuOKJzgVKh1A3/Tpx83xD
dH8v0OM8/sSKjdSPexuwpZpXCt6X7cjpi/A26DYSG/OazIe76aCSqBe9JsOrX6q6
AxBn7KOEIfU09gXqqO/VboI1bKWNlVHETQqzK6Yojvgzzpp3KS6vfEXyYlNaCb87
F/yaF4/tOpfNRptjTnmCX6iLDfloUSvdKHpMclpgG451PAv/8cuZwQzPQp/ejmmB
vizOvewd3B3wPJfn/qH0fgWpjW41SgsK7Mb+EZzscAB3uEZwFju/pe7ilvB96+vG
NXhp6K4F35rOQqKFEWiG5xL+9UxNe5iZ76WutYZqikyvzHk2Daw2qy2B/2WOI1ur
CIWaXzvdzxG4pMsIdb0UsW90KqW6AE/Cy3jVXmUFVv5jcvz2Lyq//+A4ww77qNEY
UA8i+jn1UJTeH0L2mz6Fv6iNQP5TDjnb4LqEfCKWS8x+gcEDshg4xyd80FuC0tf9
8Yb/twD1cMQXcWXQlVR1ipZhAdZ298Avvl7G8bBj21vHm20SUdnO/ntbCPOiYRJR
f+PmRYJcE3wmArR9+qikdnoyTyJ7FIGR2gFtVBtLwCFROpcJoBQ546PtqhPpIJF0
hGrTfFaDp9mAvTm7ddSQ6eatt4D9KVP+vGOqYkQvH+XTsepGZwyLnVbsIo3SBoK1
II79nf5tUxEJew8N9L6hW13NoBE6KrHZMVYgnA+bkEArOyFTH/uHeVypu1FaOBG7
Lf9H+YZyg2GVLDEH5vnLaTJc+eWfEL9r0P/97F1At3nN69lRq4zI/Faokj4NFJcb
IcNCQPqn+bNAQC9TpR+xed871zG81dveZR+NTM3CNoeEFjhHYR6jLXD+wF2uto7z
zhRvFCMzE8apgg8G5xLRl/ZOINy2iNkVnzNnWcvDQWZ8AkHlzfO7Rr9MWMZk6t3v
MAgYbHfaP4quj1Q2JN+lKCuzkp8vitfh4taGTD3s5Fv7C0z4r3JKmqvNKkAOVd+C
JHYii+SKM3+xSJya5quw+FlFh3NmREJUOsDy2DuGhSdPsqEPCS2iYwanp57hQ3kJ
aSwFjZOOfof3rSgYHnu+LXKW7C+TLU2QXB2tGTSyIp31IuiamV6wHioFItBU7mLx
7Kmci6zgeRcmVCw6hGqQdPUCK4GNQmSIe+6KXXLkUmwL4IpprTGQ2tYqSbJ2EUvK
OsOY3/N4o27zP//oYH/uwJrgZTWQKocgs6OXQ9KaQfa97KZMfkLf48irDbiMiWVJ
E0Rs9FfjpXAGPb5byDsaPcJ/8FXzsV/dxvlibkggAAJEbQzBj9RqzvF4bSe2YBb6
nWYFa8e7StqBKz7Mn9GUsQlkXQHtVq7nf4kYMMK/QRbjPOXnj3zj2idg6f03M9oQ
mWfsF6yigQ5FFMBEDk+aCfB17sR+qlxu0r8ckbq1CCPkVzY5SXjzG5DgjnWY7OsA
6wrpHHKPAGh4V0PLDiZnXsO5mQgUgVrBvO4EtyBxCHsRh2nnkybRsC1AmC4F+S/Y
Qa7H86mfy3vVkzCf51oNnWY3jdbycs8lQBVwtlqm1wT54vmDrXpNVxVMT5sHL5L1
kYwSpVe2hhijEE8tMccn96qn+bwuOScdg4hkRM/QZLcCiU65wbxFm9VCl99oe6e+
sHsj8Wtxhv4ylI+e2XLjjItmuS8zD9QTY3nJqb+JEg/wFeAXw4NCCJvOWtdrMwgL
13OHowiJ5MSsSlGk2rCL2UTwCbuwywcgMNVjPWszklBJbHhaM2yfFPAOjL3LhEUA
g7XiRuZKEohUoq60u/kp5T1oAHd8wmqIcmu3+XwsKErrovZ7M97SXesQ5hf9xy/d
CxSnjnExwkpucsvHnhVDRGjnndXWMEQ1q92yobr8jgx+pSq9suz/1q/CwfdxfWEn
yQI7rBP1hk500wq/x6C03pfmUjAyjfR9TcSEGRaelF2qEcCLNXba9J92RqoNQoZi
a3ttWwzPg5liPCT8Y+C0HRvgFbPx1eBgAMSlHacmhXAxbk/ylanj7VQGualyrN7e
+9OLWkGJbjGZ+reOQztMMJkq6OkYy/cOuXDVtS82YyipoHcGbrFAgc2NcMAe4+7O
oQFuiE26z/h9HrBd9QKy/jnKuWaE8ssBkXqxTR79ffgyPgjz9DwsEyVePujMlUBe
s9m4R9IwIlcn56ujhYphuL9bxiqivbOtMYOyapO8kBRM9Y1RNLFV9gVvXRwE8qD5
AwImyLZ7SanHp12FSyrnSVRhJiarLmwlfV+k6Qae8gavRMmVs14UyQql62/P1Q33
QZzmyOvQhcSAmaM3fgWjgoJHljPMnYMBqF0jylFUAjJSWCHk30yeKwrfbLOQ2Ejp
8yx83ITWCzPFK2qbqjpWICWAwSBkdetj2n6DsH79gNyj/J12akuKwX621UcaOEhz
YjD9ZEOKfPsjQNbAc+yqCQaelRz0L8bZzPk9Uxzt+oInuUzrr/GFFWHYnIa2edi5
LTOcdbcNE13wBRFGi30U33gPnn+v2rYe376BAqMavscuFOoaoo/YsOysALuHWdMH
62vgIjKRGwUUt1CbFJ/luY6crKy38T0qVApgXbyvUXdBBSp1KIOBLiMfG9IYa3MB
QtQquCqB9W0xEjLs693o2Tu6DhTxlziakGKx/2lbpXIuTIl0zBMek+afUyb8cyQ6
klu4KdS2urr8vrafb73e25AIoRcDNPY6okc9OGgvzNnyUF5wboENx0IPnFtsCbgd
NNiCcwvMzmPuT/WHIslqc5jtVcwVO6wZF1kP0bJFiM1iuLyj6s5Imx8Q2TELxVo0
TkP+GaYy+12nFmYzardENSPaeiQA+sj+7m/zKPfWAQnsjfJrz2wmibH+qHhHDuda
ljcTaFX7E2gZmc3Vmp19I0YF1I6ISyixbMqgynekbU+a4Ma7cFsZq9AUVHip2wuw
4xkHmMWlrY6I6DTVBgZ0VRBbz5g61dW5KDZo1FZt2iHNvK/pwSkv2uKrlVZ7vUkJ
CugPoShyriRQIlie/VmTqYAzqO6QRZN6KUDU7V5Pd+ZsbCtazGYTQzSnIBwV8eUU
oh62vgvUhNned4DR9PEj/fpzxOL/Fn1q1XOHzkxE0jNb/8Bp5qY139orI9HcnXzp
hBUhL1Bx7HPLyJJMUu8IkIll2akpzPkkSftgcLTFXgF6hAhYmR/NPj/J2wC+YxTK
y9lOvr5H7ddIShxMmF3vs++rVTUmMPPvDZI4WVqTpeLj8rZBlpoT2Koxut5eGzMJ
x4oXLLw0pWBD73SxSsS9S5NfS6T3hGiP5wl7Ru/ugHVvMo7BUVEq5ecSfXXRx2Ek
/a7oEnGkPjwSmyoARElK/QhP9tjrg8eD4mGsZCZ7prf+aUTIyjEQNJd/T2cDY4Wr
k4wbAybaCROC3VTh+yeSpnKUJ8DBTCWdHPsn9DVt+XrPwVC2ktFC+1AD3xPULQdF
Sg//l54PVJzqs1dic5Ofr9vL4EB9+yUtkohvMa1rzwUyutC5vo7st9uiFyyoaXYx
cAW05pzR75yeswM7j70GGZsSSGeoF9SRGwaT4HeAAbiCpaydKmkv3VkxX3UuC2iL
ZCMtVu/zV5W0XJ7ALV0OYcTqFC03eSTbIAmFhGl97ZP3C9tmUT3aiatRm+s/vrYQ
6MMJ+5nmW4O4mw3pn0xameRKGn2hjXJrBaiZCI6cBOFa8Y43kAzvIaERu7pqPhVa
QsEImjgi3cM5m15aRScOfWMXKh6wMVWOQFn4DgZXhYJUh1kmoA+oQ0S7/k1ig3z0
Tocv2mystxEDM91nOEonhObxeNQbIiAn8Oo0hJN2MAg1HA8qpDHYbuSOfF5fiKk5
84lh3U/S8rArwmgEJOEq5FAiO7+y66oJnuSu4+W/+KPfmBJpzQjM2orvnElK9N1/
M7vFkb9jZf9Jb9jYf4V9voTP1wh3ljXyUKLAVZf4ZDZLsP1GYYWbeEwX+yh1QYc5
i3cgpN+HLKeJvnHCD/X4Zrrmkh+kvtBZq5nilM8FLnIeO7YjKvJUu0t3th7kM097
5gFfEWLhC5hL/fHDRHCA+vQkU//m3rNsM6+9o63hHXDhR0XVuzN2wtmjP44bLpA4
M5mxrp8e49yuGKK5MImMFOngMpL0CC1tRJriadeF8ODDR4QIbDLS1R4qJ0zBZBjC
g5z9ONToqJTfLK0nOfEmw7gUbe1aQwqvKlGnMgLQYbA7Y4oNeuY9GScSW2fO4Odr
LhiH7mlyMb3m8I0g4P/1mJYctx/l5EijGcBClYskhRtgO7eCyj1uEOhEJyetMIgh
LBwUhblwSdThjja1sb5mWU0FPt6I06k1sBJ4HcenE9zvFzg/+1cNd8Anp71AJL8C
rjm51waPjsNZsuuXq31hhEXt5Zhvx06nn0Iih/AnyAplI7cwe/o2aI4HdOODc3N6
EkYgIsOubsv29jyoN21MH7z7k+UydiWK7FDsJ19RQ692tX2nZZi4Gmy3kGQheQ+2
a9uA+IZV6LAbaziDpfQ0aWWk4JPv35Q6wooAQxUuNOfJoFVYkCFtmcukMXJMEste
6GV0RyBSw/h0/Ed1Ag9VhgKlwnIzI9QjpintoR1JOE7lVRTa+Zkz6RoFg9uvnQ8+
Mq4dZPcZERg50zBN0s8lULXH19LvsCaRpnFxbXEcYFNIQPrBvbbOlmSmQd0fIBIY
yNNZ7HY1QKEcJGP72abMPN08/XNA0u80kfp/kj0ZBrWQRs2rN4NloNU9sr3z0YS6
FihWmIBRJLjkTFQw43ytlJnlQoL8Z2rRJrlf9i6mf4/Prp88KRoaqxp8mHkhQhh3
GcA/J01cBwTMz8FQZfwdUpaghZJ6+l2Z07k+kO8mS1OhsQmaftok0TOQB51Qi1cd
zIMYb2VKFyp2LWoJ/n551q+QLQCSpvHneNtB4g35woSLghPBTM0tlygP5JXkS5Sn
x2KbiJwr6YpvADIdGABuTZtU6h8z3hoLXyNIA526BBnqV+Fu/8UvqzZm6WlLvWWk
jRdETUeKy2JylJQTLWpwQf+pp5UD5wIvGW21ClxmvvGyCzP1ApnVeBJZCYmviKjM
efH9j3GE78T/ppbuTi4OtVc2xM3n4Q9xbN40g8yJF1vvT2k3WTjGa8PL3p8GZI1l
EsR3ukFw3r0Ey4za4fjWivDHPO6D0bvzVnn/tuvkFbZjLnI2eP3K5vZwC1fWcQHu
2huA39C7Jf3uDyCb8zNGdApsmJpUHzGtfv/5hqeZqnchaVoQZTAmijF6FjMVhOQA
lBD5+kZp7Ex6ybYwWe9sp5duNHiZG93Ujhdmv9H0M732zkojMdHgpQD7PBNFDwjK
06gB8Fk1uHySVouqhOs+CgMkzVtYLrOeiaVN2SYZKmY8+zZrrIKu6RzJTWNeCHxZ
erk6iSKIUbleqRVMym+zEjF1NpaP1PQj37314tEij2Wj9pHfXV30wfv6nxufNPWl
SsJAwcWw3KY1S+N8OEUABnH8XSNJXUNhu2LD4Lyd/IF/IxBxtARfjBHWFNDnhCl7
JzHWRrHOTD4mmyW38QQMxdISIORoo0HKS8CTmKqqbUfgFhALgXCA9GHOmoYnwVCe
ciuCnaIDDbH7fynxgutWmTCO5aSvtu8cbkgbjm4Gn3vrJrvmy9NM56PQO6VXB9yj
vn2rv3I565ekrK+/TvoiVpg1uJeGpk8kEOPP6xxNaR+iCZuAxBOXS+wu79ZI2EJS
3ByBfe+KiPRG4rttmcjZ5827iUNDe3+GfIwu9AMlP0BEhlFyIK8ONrccxpefEeRq
K0okYInRnYRt+FWli9jWqh7LKfi+iT7EnZQCWmoKwAETDDjoxpetp568kXdy/Qmb
Em/T6TY2OyZItX8CwF63BYS5WyR3KYj+8ZTcNUsrU6Jc2dekXPKrejtjAp0NyWu7
y94hzBjuiy+0mYubesipwVFAMtiIvvQW9Xy7CsBnMnrN/2PW7JbDd78FaiW3wjPJ
tAI0zBbncGhWHFxKNXB1rQTtY++SKDaYE3H9lSPADagK81EhI6nEM+LvweMQUzgj
0eSLMQffuU1ntdcnmqbltD760oFSFgHzPPOlCoRuFuM7QuC2uvMs09tfM0AaJRGT
xPWe5clNBVB6xg5vyOBsXu6Js2MWQlNyKs1Njhfq98Z7NPEdFpwaEpKIhBpjWtmH
7/wbSQ+ETIE5+NiNJBMCVDRh4sh4xoHFVC5Ddwk/tWZZ62rLIfjj1L9j5ae7qcDj
D71AuWaSQ5OrV67ccfo94zR8hAvhsoGjpLKkcLgU37+iss2cmhHIZpIXxBMYv4dr
VsjRbDvEITGy3SMhhihTl/NDnOuHr/Ci/zTnCMTiqkRBAvtBXrmCmFDT93uL8iK3
Oo/jLqFQEhTe8zsoZ+e4bYG2tKwuXyQiMQjXdDSEtQ3b2RxL7sC7G/45mnuzN5W7
17tIdLaYVQBcYhtpLykvOo+nsOlwr/UtjIx9WzQndjGBQtr7/E8xeGR40M5CLPpw
EOKKSHsVXld5+4nXCdinEQibc1hzMXNtVx6cw0ay1VJ7D5WaBd/+tV9esGi89y3z
tr07D6ZaEAfRNItwgAAv7iE0Kp+uPee/1672IdPxoa0RQ10lS5m0ORSTlmQ9wfIU
+uyfp3D4vtaFbrwnXz6UaI6xgck3kybM4i/3fJay2HHGB+VEZ04iIzs0qrgSeP7z
VXRB1JSP7aiNDzfSLD3xKZ+V+2JAU3oyP12/2iRTRMwBNPdAmLi70FvSMsfMv/WF
hHehSVU/Gc6UcOAT5SoZAzhpcXjiksxm6YBoHzaM/vyuqk68FbF74tU2IE3yzeVB
MideefH8PHRT9MtkuAlxtAmAet8JraYbkM90CgG7NaBAKKMYmubv43PnadWuzXMe
lB+XFBkdKzWfSUQriMUT1660BXdvmIBy63FYSkX/jvsPdhqnjyqXMKkjpq99arN1
vDGBe1ufIsDj9+edARjUVuC1PZBD8Uvt/fBKfGyvpvUeKugncga9zAbm1g2Oa658
v5xKv+7XkfENbMjvu5UIVJAwM+LrZZO1G+lStn22uTcfdNlndfz1b22qmQAfqny6
seM4mSimGdjuLhLmS98ozINdzAyD9bUOn+MEs2L9lUxRNe1Caa/PqASbKRGs1Kjj
s36okYcK29zlcsFpWDEMlYW/wcZyQigs7x2UVh41Z1glyAmpSZ+x7RGj3OF/Ohku
2nPSKMVuc1Wg1bwPGEKRsFrB/rRmujcLsKva1tr4shbmcxMzhNDAKZb61UpcWkRe
sp7+W1p/keosEa/7yauUqG+44V3SXgN264yA6Mt67N+h5+72LlDG4MxjGIQO8qQm
J3hUZB/iq2R3x5z2GI4FS52kVGb0Yupop2MbYszCUaz2TM4qyOniX2yEEB/fPZu+
9d4pDnhqf3hx/S7ooJz64X6BDIZ68Xg+3lwEBr4KJUHG7V4bQMraiLU6WCzhZ7rD
1upsdX4IvSYjZr6izX84g2vNHjEc+eQo09Z10c8gfDFmvbgIT1QAg/HOnoGM/gUn
MP/CVkYj0ltOrVdbtNv2LqddhPG+NdxIyzR0HVUK1u/QqY693ZebmJfMwLhaSorQ
8+MQvDi3v5kS1YiYrWDjIBD0ofpuJ5lJAlKW/RWygNjqblYEtMXj+cIkSGaYUWz5
jr7M9A0/6q4LjVo8Vg5cCq1xJi4MdhFtSlgaGULtUFhIGRTwWTlvciD+9yg/7QQE
IEiLWbdl/6MD40FlL9WXHk4TFtQD1ZVW5eA0xdK/v3GLlVrkrbLCvsCVa+54ulW1
Y21Hl+Dyntt1RQkkoRQg+cyBHkt2ufBXQkv9neqbfJuYluD7mWcd7vSnexuv9z3T
SsmY0lu838gQYTKcqZJe3zWGCxc8M1p/Eqpx8Gr7KKrhZegAAoKlemoFjQQqIJPU
lJNuf4R+829Vabt8Hhdto6Tw4BVzsFd8QXZjxez0ZzYDtcJnpvxm7Pp88nf5rRW2
gzjOzvso7ir1BdI9p75q5vGri7SETe0V8ZGzz9mq9H0jqMjQUS/ZchbZvb+Patbp
pL8DxwepgdvUQmU7IWmdTZomenIcp9PaPDNqhUYc1egFdGPEvTk7fr/hNcxnSKKf
CI13OrSmVC7aUI1cGpk4c+1DklGHXKiD6+3XBgHtE5GVCRIg9uPihOUObjI9FvnT
2gL4ZrY0nhFFxrMtqB8eZ6dUo2wXLq2/yDs353+mY9xTCpaXaNIzx6t10f85ptIW
7if6gTYEuKiGGn2SHvTZIpjrq4bV3VNdFfRLk0LccNI7kCcMr7IqNnM6XyfW4erX
F/JR6psH51PUmdx9swNuuTeIXzqyGcK/gUCPxhOWflYAcy1RzLYEe3Mzv165P5td
Vts8uePkFVy13XQwp56p7k9jwuFYCNnt2S/ylyta/jd9lEW8mwZ1Rbvx5mFTvjlw
byg2qUwdcsSB1trTVhIaBoRYYG43gXwGsZs1Kul0XrZaFq9C9Bt2YHmpe4OLwAGx
Pk5+zYdgoM+6dmtivMLAlKjMQIMFMuGsyyaDrsisXHyC+xeNuejp/dN3tij0mkvy
eHcsyXghSt1Yz0KCQNjUhK7jn/3tplXuu/m+c2KKvfPdZpAzjfjeaJ5jmdbcqtsa
Hb/QRdyy9vICPbUZNgIXYR4w7KuwTpl4cw1j0PPUHacbDy4qEZXC5ZO6o+WJVvi8
QNcJjPWMWYEOQndZFExpQlrVGwhMiMp070T5+tQGsOxCZ5RMaOLhwhWUPry6iDSo
JN7PMjaFpCZX/VSDl7sYc2C+bmkapEfHuYKubisCN6gsZqfbZAz8pJ7lCuFALpVk
JnKyHKgUVCncHOF9B8X/kjgfyeATWbdJDmPqjleLWs9VkJjn78BhpWB+TlLNQYZB
VG8yZvWkl6xYr1f6GpeDv28PIVxUNxKVLSFR7vP9sLGs2n4kamNTcK4xgHprrLVQ
L4waQlkESu0Yx/euHWRJ07Xv8bAUG9hpvGw8CuWPRGhOSy45jV3dWqDs3u1K/rWN
Luuq19vrD2yv8l69UPJxE7yVcQc0o86IsAQxInayEt4OKapr7LpykboZ3Yu+igl2
tNViJV+PiKULoRXsntz9iDnv77O5i8aAoW4dZG4W+0W1FJsSHxQqN2wNsrmsFBLj
8AsEpeTx8tT/eHLE5OhfSLuDgDhgQmPzFLo2EUP8+7+8mvruUYtM4DSN2XGhc4yv
4tjF7jw59ANgMtVPzYeFqZTjfvSSW9P2g3pVxIwIRDxJm7NX92gMBfo0qoV8C1wV
+JzDqKo/Vz9B/hFzfiiZ9BMRJq7rtZPhmZ1KUCsk7/BHvDxbxTTKIdDiL8Rggo4v
6amgg+G3SclXgzm/cJAXaXwkYuhaWsIaUWF+DMlvaZz4MXkQpS+I42qy8T9d4ynC
YRIqt5zy9cJPufIYga7KBv0fauKnxqHoE8kEuYtkOiPVOkAJG90j8ZtT36EM9MWo
LWJ909uXW0/ubFrhw2sTP4TsL5awEklUJGL3C8Oiq1iGZJ7mnS5DSp7tENYv2x9B
ASDXB/3N1swlTR5ha8Px80tMCYDvtWPJwHtV3ewmiiHlTznT2kJp876l3ANkmPpN
cUGg7hshcE8Skq0Eu+9yBaIBNL/XINLFC6xA6cuI8zBgpBJqOkYoZuWHb+I78WxT
ePvF5JKH7JPWFq7ES7+B7xJA8r/nkiRgfSxMywQH4vSyHbOyFcC3XzFe3tE+GRFa
oAOKgp279kfTZSczEej+WVuCwERzaEo4NqcPEN6Lus6c7qk3kbN0pEot/kTjq2d8
IiQvrlz0gEPEr8/n/1Lh0B8FGTGhZXS6H+Dv68TW1X+zbXtUQc2ldZjZa1VSrJNG
cl1PlNMxEcm3lKCOs8R7ldwWgT009635uLMQplYzDbeBy9jOTgJaCL21k5CoW7FZ
8LbenmeQnjo9E2n76XriUDGL0JUOWbRXgsfngNhDHI5NUi7NjlUE3meJxG8iIIDL
/S1EpDaSklN9hLxM6CG3mOAwspDAuActDkw+X/5FZTrw6KhI8yhsO3s+pp+oOOGC
lQVSEkNxgoBozZC6pZHW4tZak2GIT9roJmKhyE1Hv+3nORZZmGX84dl/LSzsqtRo
zYaGI22ATql8SlX6Jm+igc01V7W5DIICE4tO0qqvzrAu+zLxPi4hA8+8xLWlxL07
1k2z/ZJo+Pqn+9svJdDmKrWLnTCpJe1bjjf+JQ94rQb5iUAdVByYzZ7iInty78Pz
P2p0I9fs3h2Jx771hNxCWOCx4fyZThrwxjXNtcJiGBW8lFROJbnDZiGyjqLMpK46
Bv8Xgvww18qoU13QikETGvPCEuP4VJ4GosczI6vN4aNM23mcyVBIa8/qNgRyEufX
s8Zr2o33YD1HYvO1tlFKjCdLHg9KmqewZdUySlOPbDla1A0Z+SwzURl7Vw4gx9kG
bVOMlacN4hxCiqKIJiwrNmpILEZVc2cD5bgIn5s5gxoZigAQ/c7MkWTk++EjfrjF
kspdT7MDryaXJO8PRw6z2Q1fCBVwXodbygzW6kHUmZBp6KTJX/2TTeLSFkV/Dehd
EaPTZf7N74OTyRHRz8viVhs6HFjHDmxOCNppd+19VFnRxV0dwQlGv0OwD0P+zbJe
TGpur7ad2P85Mcrx90Lpnt/eT0ZVGxrSBuQB4VY0B6q0+6KbpFuUyHmmSaHU/FsI
iSeBj6IgLo9TblhlLLYl1HNY9ilgaFSHbJPeoxIiNR/48QkMP1hwnMzdgXcCiwUs
V65DdsJ0Duc8TZ2UmvTLWnmJS4Okmw8amWY5Fm3OepqEWRVhOexKIYuYCqsE1+k8
0gICaPU5/J74hdalXHa2ggZXZhC6kh5WfU4go5O7x/Vm6/HNgItYa1jtnjhgkn8B
FfAmDTaoJzzt4Xc+LNUgu0uNhT1fHp9tfsmkIJCqb2clkKoae38/t20H4F1YyMdl
OSnwQ2rCtSITnqJEGYvhVonKPLpSjb/+T6qV41K4W2S+IrclSqpCeb7DnLLWJ3/T
KE9qw+XC95CcRs/CrpycE19OwzcH2R8k/T3UbwHQlRF0VsrKMJ2NLYz/JBeda85y
9BxA2lVB63bl06cjm/F0YQbirWcEI2qf90FZAyu+ZZt/LXuM5v24apO6pTR+hGr0
Z6jR+jw2HzgQD+Mk6G2JEYCleAsFvAf61PxR1ayczceksm9bs6wYJzUGAW+0u1O0
pSfYzvABhSQ2X5x8lHF6V+JRqEkGC2CNRnYmorQYKTOPD8tUhrbRl3k1lEHi0JR6
Ba7DniY6J0jcxCG8OPkZsJdZSXBn63SuIrEf4SpoFdCp9Zvr0XVdikWcNeE79r1p
AYX+xz57HvQZXHaS+rqZ4igIqUjJFVek7Q2DS+0VLaIq3hIHndxTg5IZMlMqpbBX
qDpzJ3IAUp/q8YEWBzVdBK88L5jgetLzUNDGGplFNaGKXad+IdGzBnZEtXp3NXiA
xuDS4CZfypBHTzNN+nSdJm/wA6kBfvMvTDTD5CmDr14fX5TsHAdmtJRZFQOcIdHP
0SyFXbYKzmonBSG6jbOcJ8yTA7ptGT9NjLRY4YgxlJu7dnO5kE5V4YGBZ6R5QAIq
g3DbYr9TrvIpnQweYc23oVZ7PKUBt6Uq9THGTcUZInr3i/Bv7AoE1KsQAeNiDR6t
7WxiDrpG5J3Kon718444Ca6CKUNtDWPh4r9czTaMJCltkAJ52YAtCFnuyTt3D636
4W7SWewbD8SCHyOKQVg3XvTi6uXSnp1j/kHKVVd+HZXl0NhfLODKOVWzjkuqd2MG
E7m3rjN6i4SN4DX/pSYeiJWHxQcUHed2gbHu467r2RgaAAupFMlBAnAAaX6cN3Mm
0XJNgRB2+ac4OlxU4REaZ8pZJKahF/dcqRmtSdoYxhtF006FwqnybJhN11k0b3IX
V54Sf5lUjDnr3DfLBHixc5wFSi9mLoIuRXcfj1UUFV7y2wWdKDpYcw4RM5XqEIX4
jIWRBNwfV1Ti1GhHDN9TMZOJbPSAubjPxseJXuuEcQrf/FB9boF5rN4u4NpNhPJB
EDmYiBZyt2XIxgDm8sBScFDmG07AC9kZ6FAjH1nJ21Ybk+TCpxRegYE0xk8ywG6X
ocnbjvEkfC/uGMu39Ii7wsmZi/4tg4jTdTxY2lCyKt7W/4HXN8TOk+D+JLpnsAaR
if5V1bflAQf6t3Y52qf1uJU1O2M5AQ/1XO/5Ist22fHrpu9F1PJDYB5+nJLUfvPR
gOoMODHsTNTN4aKkAPAr/sv8tKh8t8irL8ZVA8szK2Ou/oH4nBsaZaqPMvLfDXc3
5AC0wN+QpXC2Nkk9zZpOkIu9AYhKk8bYAIznwR6UVB/pidFKUUFhJ/jO8AfjN+qx
GytzvilVIgsVoiMMsQKW+CicGT5vjGeSxs1daVT/2BfcEe7LSgsoExvViqB8QI3h
Mthu5AAgZyfZ60/lbs2oXjkwkU/FtW2IhYR+9q5B0NpceUIkeOI5yXOmskqu2s/R
t+/WGr8c9HB5KsExYczz3h0Kt7EDAWz8G+frMDV8s2tdJ3EimlSjd2T8IO4mWK5e
nQ35nsJdOGWcq/RwbNECNyLARO3Tm/QSHu0a6RbANMrvpNZWVyNxyeIZvIYqmnhU
J5Vya4fP4brJz6qcn4s8uN3oZT6fPMx3vr5gNry1lows9fQMky4It3LMlX8F7tn8
9x060MnQZKqcvzGNI6GqJBtCoAsjz+bQCWbOKnD+OHMS+CEfcWyK4Kt6FsGtRXGA
+Bo1l1imuOZtixe/nlohK1WqHOQ5SsJqIYztELHnZaFBDdkgQujLBCDeFDsGlQ77
W5s+NXRW9QF3cOsVdJmsNd2GwzWAWWrSB/EpmfUs9akyKLJ5htk1LGORxtlttDG0
qZaUxwibqiLKdzhioD+5GD2pX6+jhMgUPavSEUef5L4oCTrgEVFO9rlbYOxkW458
k0WwtQ9ZTpRgK3btk5F9IIPQNkRQrtDJGDh7T/jIWAlF5L0Ul1ic3METrobBx0MP
/MZTrq05hR+SLyL0QyMtQ1x2baWZtiFiBuH5Ehat8pgMbSZQUfzJ9ZXHaeJawZJc
HM4a8MXYE210nZy38b50ZvcssudBoQADM9AzCz+F1xMKM7/J9zkfeK8bUpRF9bLp
DE2ghh3sni8s5X6zZDudDgkrHhOrPNWpwP49LjA26wvLYWklt6BLzXWoNmxl2aT+
aZOH9+2hXZ5XLMuFNxN/7uwpf4IiwelERu8Eqo3Rywa6X1ojcbbSI9MvwjHRWFS8
H5MdhSIbi/m90b5ZJWMFVVyJEfvo4gSy5Av8Y7YG9UTEfTON83rXdt9fiAwRUqUv
WWV8D5wp1jKNURHbD145pR7owcoAWLg/8D9gG5vAM56w8MTOt2/hotUevBb0oYF7
rbdDlKhBB0xVFNley8sQUfefLp3Ko2ZM3QIZsr31KMthxkVdVZ9O0vykbBwE6HeI
/cGvkeU7Mt0P4ilU5DZ64HqBXzo0SYtB7eBt1mn8fpbeV1I6cA30tp38BtqDEFed
XK2VzDvg8EAZnaOSG+EyZxMzXiLoyk3ahQTZT1qFouRoSA9ODN4dhkdAFEbg2Jnr
0tfgkDOIFZjt7NfapVWMufWpEbLL5PtL71JmTUwVxPMY0W+C5PoPkimTlEhqLCQx
POgMViRij3jwkfST2Dn+jDXvMLFurvcd21pKL6qmGY6DKeswr76dkTEdUlLj1Lj/
IN/Pizqt04qCk3Gggm2s9sKODw5Zy0nlJDY7J3CRX1wIvrlx19vlhJDtR4wIGebG
/PvN3RPZ7Fxy/EVtqV5U1pCWHkTBBfFo+psF9e/Y7ciIxT0Ps8jX3RlkVahEHbZp
eCV4n8vs1hpKFkL3Ma222vCAXUc1n/utbIwDcmIkMrOv1ZawGZh7YMKxWBouSJDR
zYbavqM+b5eozR1+juerducKBBXaaPIZogX/+WaHlYYtYUO1WPOJhpjsL7IjYn0a
Yno9kZEWZxKybiU+8W2mUffIh88mT6jG3TkEYoeRQdchuIb+5mqOjjijetwlGAhj
ejt3V0c3DjuA6XIHsSCnjZPxlYTlPqUMaw3ENL8ujIOT9tcj2qbfTLtNHO/QVRDl
VGeMh9DKJO9vyBxcRjnGWNn5NITW6nEbQSUlWLIN8L4XV4Xv3DsZBnRT+6jK5EXg
W5cQRkIlHkVlkCrl+UcUD/pKQw2JVqIlxR3jNDEP6E8l2BXOdpZudnU50mueolOt
M9CvQqu++S3m4lTjDNNIL5nElb3DdFXvJ2mKr47sXKB39YlFl8BCVrtG/1PUe//8
+p8YcRghfMIyb/cf1O4xum2kfFTNbI84mrbgK4W7+HZzyrV6idQK8m4jdVu8Gw4+
1hM3DHDLVrtMRY4lGAr49RNO+XV3OWCMLfkuDKH9QlsqA6Elwt4yDaJ4Y6NXABMm
ScDtk+w4rm4G1smu9TpxZyQyO7xmc6TYUR9CizUjjf67autoLbhuACVftlGnv6yy
e6JPyYWaJHIybsPnrrUOu2+e8eGtSWISLIO8dPRs+Sl9RssVH2mXX62HEyGWuV+M
R8vSONQaimAaFxgDvIN8CZ2Zounfiz1waIGhVxhsbxeQ4pLXC38I2BJEHfMyYTF9
47fzHNagZOBnT8BtMFOBLsDlptoxAge1NEEBC9K1/lDTJxgT8cUd6JPeDjbPqMDU
GLDU6i6I8nwdQ6Gl7dbbyqyqHEazMqfxzrgvapF+j2bw6iuHwNLOYJ+XijKmfTBJ
0YVJh1dIYJB++c/vas0q/BLbxmV0a1HgUyDL0osKxJLALrTjAMbx2pFNV498f6Jo
tAFvyoOEZbcimTFio/pbJiNn5hFqnw1j9IrDIFtN1v6QAZT6N+3uqQR2xktB6No+
ssL24gP/5EkR+rBrDuMhYA+IPMo0g+r5tG2GcDaDqeWj3/iboU5PJWX97HUVz5ra
DACOR5P3BG2K8dJBzUH549jxl10eOG0XCUvu9YRAKhU4PfARBru7+I1JcOhghOUP
GYCs6xwbMoMb4j3RVvwpVYT66hUN9M/h/e8MbFnFQx+OleBSRwsYsdZd9yfD1zbp
h0qlsrAdDeAxwBVBom4RzTz4lurEWJoW4ao8Aq1RSPDVjyLGQ4qVtDgTGfUCDffJ
Euhln4Ex5xD8H9LWqqKYsfvG02cxlLQx9Gp3t9fr2ALOSFxRKfInJ2f2wMxls7C9
G+9INO7PKOi1bFk4Of6Kg52QZpYx4nHQxFpYkD+u4YpgBhbvXIihcNwGlepBulVc
bwQfjxTWrV/yE67zG5yWLs8rtjCz+BYUukNyBQsrrnsTy9zoBiMwbwfBzY9tAizV
+DI02SbJVy4qEbstydleIDk0CVY+l2DmcfyxTUNxG1oEItu2YSmqXVKQqWLJmjFu
rk5ZG5oOycWaz4q0lWefGMkybnRLUEihQxJST415g3gBlEh/RqIeZcgM/Kp4WiYC
WC7QsfpD8tEr/M4su7OIz3XeivwkL2h98qxdqTobIZhhuRh9pT/ZVeRCC9eNMEG7
QrVv0MObG6MBKdXXALfG7T3zZhIa/rYD4HzgqcRExBdoIz2NeS5tOwH121LCuPmM
ePWdMXiEr4RArgBNayXX5zshQLC6ImQ/xG+MIiADPKqD2zt1+gshYTIBVaqvYdez
cHbHc5Sh9YWSfZfA35hz0eiJsnvlp4pXQY+PDvj8VjG68y2hM6Ym8xXzf6+aPmqh
qzhInszJpYvfJY2n2SXFdDOUeoK9UNRVOhdpNAaQlKa8b7EtAE+L4kap48P0w71j
vmsqunK/A1I/mswVoLi1odZBcH4ybh7HmL17o7brBDWqyUZVwb3d7NwcrwLaALNL
wuGtBVt+AArqNE5+472GEu13WxTB6Y43D59erX+1Eprc+b5QLGKuc6eDOh7bVHgu
yq1AWwWp0/EWVgXPZTONvCT+XAml2XwJmroCo7iv7YKENPEBCbJukAwRTTsKQiHN
4ZsBCJBbxxbb7QdC3ZCR3F8vs1Fas0JCCWYMGCzNbho1GGhnR2ffPh++3JKpB5lR
2F/exOgRf0FINDKiNsVXpeWVN4GLJ2JJObRkthFNlmxyqAeVOIiU4BTl0GJduov4
IALJRIsfBhX+goEnyqS9izQO63thHaTEQNeD7IzSwjbHl2vn1zobgHGJ+UbF53Bx
HvuUBOQall+LM+hzOY5ZwuX/p/hR/s22M2mSl0GuAmPjO9t8wY7dkF0yhj2s2bfW
ZbA2uhQL2GIq3MAo5zLxC1dcxJtZ/n+MQ/N/rW68GJ5vJGwmA/BVzLEmjVU42t/z
V6omxyt8AVSpq7nY5NfNQbcaeY0bDRPdw7hWSy+qEzNZpuTmrvUyzMyan+z3oEsW
1Mf4UpZRfX05VhS1uPLGFJVjEqgM+aVT10gZ9gsCJApq6fOyroC41BxFM8v/UKOJ
w3xuBRE/MEP6PKMtjyTB0cDNJJipnJDdqa2wyY9WtXMXkNvx562UUgj5rdchpQTw
ot5fy/wFlse7jI3RZb/VkI6U64CyUYIeerCJgEObHuFAwUGxMy5d2zbjxy4x2wvE
w/yTJ+sALmELeoHNQPRZSZP4P8RVWbs5WCoP0w9tktwfpxNHsxuNjjB/P03InpvU
XXsGHbxH3JPqwVX29dR2HLdNBDKQldpL1AMx1Fo3nkqLcutaEjlVCTSkPZ3vMSVu
Xcv4aUfEgQbqiXn75scSBNVqUvDSECPO2vdXoFp9GkTybUXRW5h+rezL7odWh8hw
by3LberAM9zJJm/R/enKPpZJ/97AD8PL8gZIJbEAEvOCLbZVWgBGSYC7PrOghbvd
tZyTmEsxSlTe3B5onfAV+vVQ0LnKGB/kLFcEWVFf9bpOkKn8b0faAhjGNZR8S0SC
kSa3MRLGuk8Ixi/IWUly+CdNmtglILgrwHjQPWatTazhCf9GC+50+GjpDaOjkPNH
hz2RyfS/hIL9m2RZapt2fCPV0zVF4xFgg1vMOujn+8kS4eerChQLqbv8WrNUl1DM
SqjpdB3XkHgdO13b2Kylp/7FFAGA165wWHrLzUICikm1H172lPOsXtc/+Ln823sR
W5CTofqlHOxGisZkEBonADbgPpBOL5jF//vmNDcbZkHWN6WZpzlXjf3rzhMxGyGw
BGhj+3RO7f+Y+y9UCgNcO+J2gP4x7XaZjVxzt0z52W1DhNPHfBx6Gfmp8bEC7eHh
qwm8g0IYRoJlI1jbVepeiLer3oISMO9tLZfnYEoch+D5PNmOHhbA29AUk7ZCcAQU
cQqdCw9JaBo08hN/JbT8EecfcjOQiGP9LkpKoHdcaMh9bKkR+L8+yLgJ4qMIRXsx
oGV+DqkYzQ3my8/lsTuFi6w2EXCbO+wEBVDJgEUhw1iGonyV+KpI35qKQT3LTLKn
EYFOCR3+DJj7wcMLkH4lUPQK9hkYhDLStPfFcepBqHcfo8RNwSosmHCFJd2MxP+B
LqxwzXZVEZGGb+AJxDRgDp1sAx44hYXxOgGIc1QnWGSOXIRJY79E53xZGVYnC/ZU
RB7uvBzKBrBMCcEcMiWuD14N6+aPrf4jF2r6r01d1fB/OATFqA17JxEHMhzNfzHz
9oqlVCbeNgouXj3hoS85zacoRMQH0629OJK0TRq/yHObG9/X/d0FzMKpsON7i16o
3xWfWnsEVmnpk6nFqcHOxWSLWuEfSAj80Z9W/gCkDqPJ4nE8ObVWzcQ08r96TQLP
vXme9TZhfvRlgZl3mFoA2IiIU8N/Cm4mEDLruxBD10msa4iH6AWxeF2Z416YtDFu
9KC8IV31/QA48y1NUiln8w6iC8lKCGdfQitP0NA2WgYETTIv32X458vfGvxubml+
7HQ1/IXpwS7Wl49ZusvDOX23GEK7Rx6ck8q83NUcH0zsMmgGy7vZFE+Y6t34PXlv
l/aJuiStqYUve80B0lGqxlzmBJe9z/Ktvd6mMj/CJg9dS6JzEyp5/ZjJiuZcLM2t
/VSbj/e43XllfktDmBshPAJvI/0Hi+VL0GYKBd0stI48mxl6Q1jP4G1VBLs8cCgN
ZqgWztC0dCHuLYUgkTgAMyaG5RbjzMB2rt/5Op+LC+Qo2AZt670x1s2RAD8cc2AD
6q4Det7zNrGLECglju9EJUi552PgEj2ehUXyYLr8RaF3XAquSpmnmGmyQPpjfVcu
aiqzUTitXOYcd0Ss5m8Juksi324HA1LY8wZaLfXyKrHkmK8vxV7qOOts783oMWNx
87kYRA/KK5oFCusolBI+C0/lWxT48gCM4D9nIc2MqSInG59ZlzXDKZeuaUB8dsQT
fkcs1F6luaqBsJA4Z76vnox13/HgPSPlY4FJ7c4+6Jh5HnFdCskCzJISbNVwsTOZ
J3BZuHFnA4rsW1AB5NEia+T9RGk49WYHB4fTmHoESKckMsNMeJ/lO/hykfH24qxb
kqh2ay1R22vd6n+eVp0sU9okcNsYOKiVnm8WSoiXt06+BMQfhhfrQvhFqwnLD/68
p9ORcAFdUUqUwAtvE2a0cUn8SLvqzMOKRh0bh1czwXxhRSem3ny+IYdbBAxUu18Z
zuam9EzX3DsGUlfmFBls3J8pDvCAqWjH8CgqPipnKSR9xslaN3THbtpwbbL+Of7I
vHfYUMjuwdOOtZmgtlgizpdMGXlTRV366pCtXDWv8+h6s7tq6fzv35EsT1AUKctR
Dtn9YMco5LqAnGikgxYGDJTx9Stv9WGq5tOYo3jkCmLssKX7tcltawOLWJxm05Oq
WA8YzoYcRYN5TnSVEmvidEFkHPYF+nBChW439cb1fkiFmTMcRd7fqNsYGBjbuQTz
Cl4W4NoI6BSY/eaRMw1jcIj2h38BhSiFdFlEzfIrRzdDNjJs8JpzaSWlkkaoDnXT
at2sVCp8TiY3ImAWFvX/7jMKVNmfueH0G4s3WxulY09PVLgN6ikceh09ZNuHCwXH
BzRjbldPlCce1jbNtV6D0XLXrMG2YSdPkcBSQg+Vux1+yyLjwxIXhHoUxj4AgtRo
LMlcBf3uHqfM8tCO8qw64n+MR6OAnggqBd9SnNfIivMEtvUXdwxpA7hZsmoR+Iva
Hne3YOh5Lpiph9muv4s2vnhAUsc4MgMPmxO7oaIf81Y5QWwd4abtIK1IS8xVcHx5
RRFGVcjs+exagzXo8xzdonMQncnWf7sQbX6J9PmygTghb2jkT8Ed3tMH6nGCIzR2
SkXdNo/t8ZRHPzasBBZrx5GvMsmk3fB+pWuiaYchtlJgbOm4ZiWhDM1wh4+dDkJi
1a2rta1IzS8Ab51YwXgD/jc0fQGn4ByvhJAwBo1gXIPZ5TEhAUwg8odG1h3aTDdS
P0C5y8pl6+leXxhYQoNzEAlijcdbCshYfowFPgjeiUwsIJQq8ZvtbE1sJt1vg/aS
XHi9LBdiZiRNaO56hB97bfJVrUqeWFJYFtCZeV2K6Pi4XNOjrpaakxY4Ory00XlQ
J8zUFVhdBzw9K6bWOpklbSAkF4S+Kof4AiOQBfO8iHfs4QsQFqOYdZowgGLUTlmW
ScILdCylDSqehp4ninuzBAO/ZVYiiQClmmRrez4kx49J9WlRpo2EaSsI+nYpyOE9
jDIu9r1ll+q9Ld3TE10AybSYb9y797bElsZoT1cserNttts7g/jwvs5XmLvVsWZ/
GLfEhVdXxybeRdVNXR1eDVvPIiuq7dsK5SgY/p5BTsIJiiyUbYSM6OUtz68mW2IE
2/PAbE9hhJPWhI/LT+FBgYAE5uxDT7RhgRCaPXfe1mnNdMtG22FNtZtAJuHGu8/a
LmgwG2zp4A6w1RNYM/zqTsyzIOXXnowtjLRU667eR4wi6NOLU2VaiYDG73GIacaX
6iBYs/GSZ2gVY8Ulh/fre3w426gyPOejw5vRBtJdgSEA1XMydeDBJGovCzEp2U/S
uDtJuNS+l5dYys4zrQEZBHUG2jNU6ltbsc9jk8gv00w0r5FgsoAybrAuiO70XfRT
dpGpMiQqQDxIio96zKsSP9wWQGOCZDYdtd/lSJcee2SmIbVCdmkCZv1PhjNNEf2y
3Bz4lks/ffQeDyeJBQBuXf0QXVktbrtLcszB+RfffzybHbHcF17y8id2Uq7lLzX6
4d+C5/4m+T14NCpMvzZM35SPp2EkiMTrEPbSPuDT9bY36PJ5ET6noiPj/DFj3sU3
1GHuPiq9jl/g1Hrf/3hclELLyi2OpLx2fTezdYxgIagPTBqp6SKBmfhf+KxDnRWV
2nWLWZTihn/RktytV4rR7b9b1vZTDLvBuu6bzaOoF10GLEd0MtAJ0Gu5VSDrQ4s1
evurHP3NFy3lx2qLxP/Mwvt/xlRxuEzTQ797IfWqo/O7WD8C4qklpIJagoVGzRFQ
cINzuZPMG8gNkVZy0cIB0FkmwTUBWfmLlJrG7zmw571CHu/squHLN73ueMlP2zfb
+eNlsRPLj+p9Xr1/7es3sHpveUeT1e0C05jPKSEsXJ4KRZzyjtF86EufgXagE/Ql
gNGgavxFhftjrCKQbNBE+EnFeAsWfSC2JgsjHelbIBMCN91zjEkyL8LeK/koQmCV
dWNYKuB0UN9uJ/+vj+uyJDUN44G4mIv1xZ8y6/u8nH/uuPghBzTSr0A9mlm5fhPC
EXC1FlLM43ED4hzz0rFVwlUyUmTBE1ZWM/+7TgvtIq+IQ2oC3T2S6/kkYYfavh23
Pxvy9+Nn4CUQjJuWe+HWYrlDgmfc/Zeym5r8/szZlQt8oRft1iGCjj6TdZ5qW3De
QOY6Oq00s/wIp3Gp9ClHGCu+b1mKJ2NuNudphxt0URYKonaTvUJEuPLjOFisjrHb
XEfdwo0pusvH+ihMDCUOzZPzbAVQWT+59YtahKWUxkHqw+U/DvhToiJccVF003f6
sODue/reFWbNrvT5oR3MNpkvf2YDVnhQMf3zIsgm2y+qiDgGkJAdFtmNCSlWpn0q
8EJliknwct+6K53kL29GoMi9chYo30CqihSeftdRrumZuFsiSrY7jHaVe84iGde3
xUusvN3B+aenLlqB9XPmJdGSXj6UNnQnNH3p4Co1S7gGsNZmyFkgwTxhXQRDv0VG
tLaJe0j6F6K7bw17IJhegbdJHa27Hqz9ox37Z25bMz5yU3wk1siLOfly/R1mAOwO
I6t+cyAVIgMDb98tkiZwiXy4v6nqWVk89frg7xJsKPfdAI1bvcoTTRoaJVgXdMdu
DePbvUmmY5io7Q50FfoN7kg37qimr2o0EijKcFxnldudX5KoC6BCAboKBNm051N8
V7wws0o93GKPeJUZ6xxda7WjmQtnzAt1f9y4zx89DASAALBB2iFBj4evLMP02C5s
THhXWSG/tR7qxtvP1luLhgc/8CZu4WhdNPokgp93oon3cl6lcYt5I4TIAZHGg6bx
SNCwdyKidUzkUVermBcQfCdXDSmOCalngFMjBe6QBK/b67OXMzHHSHCwjpUCBQK1
KBGURXCAxOHIYOoyjTeLGfnSbouciTm5/TRrTRQ/PMOnH39DD3WlVPPanLtO//a0
hfBCa+OwoS0w94wxJHKWikn3+geJY6M3dBFUrpZl+DERt0nt+pnFNbSLbQNBOGxi
sM69IRUPpPzEhN4kzQ3ND7hQTeKf6GHstOZfSXkmIT15I9qff+x3SXVSdkyGXiPs
ojcFgoa/sEUiNYNHsRvaPU8MvXliDUY9zKLDInupENosmYlR3mEIpQZCBCfQYj1u
YnvGUeBqNGoVAKhajSZpIBmIwQ0z7XRA+UqKI+csCbfvVAzsllcSDkhePJBe6uHt
Gfe6d+vgCeGo0JuzBHgiF7LZ4dVAYKk2iftIiIGUl9fjO70XybVJUcL9ZbcRtmya
Pg6h2H02RmreuD50B7fxq85sBvQv32gUZ+s5m3VWesiImOAHAdz7HeROHZ0IbtfU
7guICNaS4vhf0BnpQzRUH5PF+eP33s1VSFxQDyqWDmSRPyDJsRLJZUYb/43cMP8Q
v95DBakhEXVu6TRf67u7l9hU6sqKtulWneb47pElcAV3ffry+/4kvAksDSY6Y+X3
Uwzhcu7SeyADqGsCWVMA6lLdGV/SPSxGhHqtzhivRUKC2bpaVvhJLQx/W8jO6z0y
di4FU3NaWVgFqZoxn+PZMs8mJW0M88DgPj1OHRgUz2dcjhtpje2ZJfi4esrYXAek
RjB0vATGYBMO6nswtkT98olw1AnXup7RbjeFU5LOMeois/2USvB0CukgOfbeRBCs
VbvGixFPr6ec0PTfwqwhzm3t9955SK6EHZeUwbNhX1DiMeYFuUBjhZIcdUgN519f
utLnMEbiBUyBSPn/nqfLLzrpoAitSzdp80h1O4trKjzdwa3ae2JHrCNCPMA2ryoV
vETa+tlGqHlz0ny11pxLZEHYZHkDAVHmoJueZNoNKyQ5S0dzBUEoX1PCXk7VNOP2
YtMCLDoD2x0NBlUx+DHXHn6PziJuzu8nZ2IA+SYGd7/wMtPbqQZkkMTUhO64VP9H
cQwiZRUlba3/YOe3vLZCpa8AQ8y85n4JPXs0ckvqZ6vbhrr5qG8YVDhz/vD13puQ
JGCtWlfaCURlu+GcYPPgKoSA8c1oIyF74iCwb10U/7WUPRmZpLbPi/o20wR/0FVD
YZL43Jp/QmC97ff3rlOpd0L9t211vK2yn1i7rvKG0ywlrbFcM3POeURrd2kYpw1I
H/pb2TAnRVKLAHrv1TPtMOa/O4/+9ps3XRYyaeCMgXe6NgSiRw/GfSJbfmMK91rs
SptfxjGWlXBEd3GN/KyEKY4+/P6LDN20yk1K9qhjMdkCycL3IXP8pySeOme5c9Yw
XaXGVGqQlpIQITH/fLH/jGpKNHuLtfZoykj/oEY2AgkTXe4uEQXeFVvYTMFl0d8q
T8byBD6QNAYhTI1/TioPRXqbXfjgRC64c7UPsJ0WoO9L4IkL1Ti014dQsHNy+8Mh
2xAyQkG2ittSMjdQ+fYTG57A5A2xHo6w0TI4I89ZxG54k327SoVvRv+hPiKEgcz2
kkNjVs8hiJbN2GRSc0Crg5ZCQ8t1sZMgNRhRWfEd1tuhkuUr6yM0NVerOOwexKjX
BeR3lgMy+cxdx0I9HkSiWyWoterq8wjZsviZLoX+vZ1qL412i/eZRK9yVoylMrmp
SW9En1hNBlcFS6ZA6R+IhD2sWCj/Mbd+uH8ow5uXRVDQw/21dqWKXo0fy/GBEyzi
L49xpiLBSHXax0wzbMquEjBhf8yIscIEny6d05ojY6VjNfh6xDjJADfFHH3WrMqj
tXhkaBsnXAJb+uxaP4go8PoPeBgQ7+szg1gAUOiX2waTxZ0VIuOhOqGYd5Gs8gXX
mABOy0TJ+KSRAaD7DWc4amWRukKjD08HPXDlPwTxvpqmatdhGhpxvujPLYb145uF
h/EuciRQFTzNz0+xOtdWz5AmpF7gixdeECDa6PpNJ0T9bzkOO0mgME6Lr3lJ5X0Q
WsutFRYi72ULVFI90d8qPYcKRCDeqBWzpzC3jLyPGsifY97WIcd6xXez9Q7RVZ6V
xJdFZGQ85d07XUxbF9u6ELSdoSqjGRU3uy5cJrfpfDYEskUkce2oGZgkaFht7oMi
rHshqYisEeJGNsVvnxD9c6QFPhFJ+OH3l5cts0bLmlYS9lwMhoaap/SNoNYDTX4N
kdKAmWHx+PZqzWRZeVMZA8b4SAcFpmOXNTSTXOnbKpLRrRnvVwuqlJ2h1Aci6xtK
lOHEv4015x21wEkcJr4b6KSTu8r8LeHMY9rEG+UFeUST+YwCdj5K/nLBDdYe5Xba
cfN14DKtZD9R5dbfBbmCnQYzwGe2+4AaFKMteuFcJ1GGYoGpSJzT6TDrh+BeTT3U
xEzhhGmq+FYQ0M/0DRHJQtBytR0ReloXuy7f05fg7GTVNEj2FretBxxIPxxHddwN
q5SihbfOP0mdabJUr+vJW3cmeFpfyeLBokETnTlabePAG4lNuNsm3DgY8R6TYixC
HOQfKPcpmdBar70gF1nZ0B4z4ykCGF7qpy5pdqb/aKFTh1JrHXjOMJeX05Yb61Dg
KGx8pBvDlf2bHm838lEjujU9ujxG4OL8W9ojL/3KnwKxvJwwF7rdFXlzpQ7RSwTc
1tA3UjfCbsZJ5WmSxBGsaxBoCsHZAVQiq6Y89GGzeu8V+uJ/BwjeQhdAAvTzcoj4
UhmxpMGKA3cUtx7zT23j7kar6dMcT5+ZnAyEHyFY/hITIb98aI626QbfcI0YKsAd
s+3phQ3tBi8EO0zz1MOJe3/pBcQ8sU4oIRiPWW72Eu+Fi4QFvWVWHUb5GEDnQ+Lg
vr+Jkybjx2CY6PL2Q7mcfe9QBCcFnYDw4uh5wf6v6HOJo44k/WmIoZUClLLmKrcd
AjGRVWTpPPlA5vEj95lWJ3dh78U65pyQmhIjkNh5erjo/KjMyWQ/SYl3NoddJjYs
XUw7F9p5x3ubdyydYJ372Ny1zMsHZMr9KtDtOlIKPqz0fAjdisFCrQxYlrS1F1vF
u9RMcYirJT6i4Zz13Mm4iHYluACQU0TAsRxz23XE8Te+gbWXMYJsFEmw6NQpRFFh
1bAy7g19DLc/DkykoSFlq+TG5mZvEVc8gv9A8Et0Po66ntUbIhtHb0svZBUOGUqC
UKIkASBMt45QDrLo3TJCHs/hT6UK2X83bVValz1/bb1EuFHfI8zxHEtEma+wL47Z
5Acbeo6gpMO0h2d4E3KsH8vgc2rf7etjsBUG73ht1/kPT31FgjzQK+GkW7EG8yxS
mn4a9dnWAX1HRQdbTRqTaPrs+4rhBl2mnWnb7fJ/iO6tfYdidpI60UkpPuaeAO7O
n1T0OW950ebB/sBg3uiMWgnaQALiXfy9chF1mYIGzbZ5nXq+tIBv4d8FIcqCHPWo
HnHanpsg1AzUQ5SrX6MLwoX8nxoHCyiTxuppudjHAmtbCD+vayVwtKQRBOrufBfs
AYzZxUMCul4/Guxdis1+I+g0t/j8y7gWfTRQ3tWxsIo1m0ClsqWRMX5J0ceJwRTx
V4pDa11vge1bzIunK1pPsRmICOoqjn1DDyjHK5oZFWoX+sFZ8gBBmllaxt45T7kk
jYmcYfT3ar5o/fXeolRYy06anZxaziKxGv/3EyuIIjqZnEj52yuS13fqe2u3Yp9l
ovIIF7yAegUNqxCDalblQGahp87Tpcg6X/bxUUQXxEj+HNJ59Apr/Ca/XrUu1D1I
fmRjr7kg4jp7xQFxzMqoOcu63D7q9mtZysa+G5xIZYLw9X2JYSAuxKIHPte92TsL
Z3WRhiTdwED1jt8ggiyD/zejRqpgAbIGHxui73l4/hhSV1eZXhUrHZRXoyAWW99n
PDRkAW/cxwRpKkodHdTZVMRVpCh3fZh8KxvTg5KsQNlnX4rvGe5yQwlrFR59A11q
/C4AFbTm3LlRLTL/1nFW1gaPd9ZGtyDaksD4/1EkoCAdmoTL8LEb96GHU+lksSgA
pyb2SoB03TX2XXTWo3ZIuQWB9Ket5o9bpi1ORoqFrYjXy563GxTZ8mlH1lQ1bv5m
/hcccJhBIhpyZtTjIYN9fX+zfNuMdUd0RJ8sCjoRIZFznK4vedEIxHI2qUOOfYN4
q48ULuYPYJFXEbgIyodIKLLbAVjLytT7qny8U1KhcsGKCfp7aU1Hr8vkKIrQwhBg
da2NEJKuwoY54sB4JQZlIJr0ljMyosPcu1z9FXIKlsfpSmfYFF31me0p2Prsg1Tu
a7Xqa+FnOgxgW9zlh/ml3u8Yh4V4nVwpFTaMeqO07ZaE08x4V6vw1O+py7E4GEwo
2Iu374vGgq8PV5ZQbQuAfCgXw4xNYhQDeXpneZINtIGb88Pu7e+we0UsWD4AGKzQ
puFNG2Xug/VN2cAQ6IsDLCOc2lWPA/dQczZz+T0xOVdsKJa1103L2sLOznqNAvIr
r0RHuhR6YNponrz3uWZNQ+2qqk40RhWRmSU7QYmbEuGCkmft/lB9zpVbcNNSHwtb
jll8E5pwNrNuSnhGps2sJQWmILh90tyIR8G4XYTc/k3MnHRkdnX/jA+eikiWlnmS
mQuUKixsntK32xvMbIOurG3KnSIpeL1DxfHqFL96O9Td8Qn+p6keO377aWfsmv9K
b7I3wXTwomQxzSPFMLbm4wVc7b/ocrF+otGonMB4QOdAsg3ZOW6D9nN5rbiuV6NM
iVWNakpLYM8ushEJPZUNIzFiG9sZ5YylNwlETRoLzkbBjqK3yMrQIumw3lUq8Slt
ypbFuPFgiZi15yT/po4VOxpoShoV5koH+gxOqKGeUOjGkHOu6NH0+FRLE2pO9D9p
QqhtLqm8PYiuq4PZcZj1ByIuBr3cVYehe8bYiFlhlltJGjpsGnjD75T8KlqBDv8a
f6/iXG6QGNJAfY2GDq290rc9rdSXEyditH7f6/uTQA3Dz+B+jIGclVtAyuylQs8t
Jri1RcoLN7f0RRKIsjaKOy3EtQhxGOvnNid9+lkE1O9YHptMRZW6r9gJH+XYi+Vb
p/ffiEBAh719K1a7TZPPxDImnD2P2aazVxVMmowm/RlggjjUeL1juz1UwNitKIhh
AWG2kCMKC5I8BGs/cy86pOl5n8pimXQe9fdpuEy0ppvDxG65ZU/bXbLpi3YZ6j0n
npu/0jNAESCqSQlvZVHrqMNClOd3guRNPg8zOyrI2CYmDhOlqDQarwlNtozc6m9P
JCz0KHj41G/fCro6OLg/sf5xJBFm/FQ0YS229HUk0r48y1MCqu3ftknXcSazKcvj
BttNCHSsfa8rPqFyxJRDQEdhDg2+q3gheffhE7PPWvAOz9IUn31Ix4eX0QGqHK+6
gODJQHLhJhSRQRpe/mQtAKGFNDynJ5I6GTe3nERxaFR/6at6L9APoTyUIdvnql3D
U/UXXKjtPtz0SUYA0igC1X8h7dBp0iJnaCNgDv/sfTe6wspcNPe5xG8bjvxsLUfE
siqbnGMjm173IocsF5Qm2e/ZB7MVtH37/wL4XhSJzDzLXTNSBcEo5y5sPWwIixHD
MUVD7SE2Lwf3XHzQ299/BZdmloYeOkwe6xTO+q2h7gSfcELLeOaMqcHaQCZaJdUB
x5tXfy8Rq6+J2kD03GWHi9GsGJVjrQm1lLNBzIKwg1S2whOTiM1rgEQlPvM4d2ax
4KHSk8o3DW3Rj+uSCgCrAkRlxxVLxxZr9kTT+rb7GFdkQz7YSR5+GqUCvedN7xY6
PcgM+B60tL0OxvOcRRaTZrVTrT1DTciNNmwmMylLYe24CiDWdtVSYWnjmTMYG+Lv
2a71uG5w/BLgBddsVXn62o5RA04cN/rZalYo6gMtaJRgIxD79uQtruERsKIFJyoa
q6CikvjM3Agt+bwcCGaQ4qjvUe4jWxN7cwEwgn9M0+nmMEY9zg/5q2VBORuOtjfH
HfCTHRHVyjz+wiEFldWGfZJ5KbjCBgWEVdDJR2/fSS6JzGyDQOYV6weYbOSESSH9
6rhRvXjYncsbTe4Fy9PFblrYm0lkxK7Caa2QevlZ55dwcrF2budZdxyXca5fAQkD
ityZ1tzHhTZhMBcezVUVYXh8ewwL13wxrLXge+xM4WSRo53UabXCzQVdYbgj4u3D
WJn9CzFheTYjNxoV/VfMOfY4dboiZBy891YjOuIg9KR67wo9Vx5wizW+JFliO24S
n9fykOTSCT8wqmPpgt/9WdUUs5kZAQTEi3XrnBlxhojF5UzAHesFsD7xeLiC0sfj
rzLsNhZjCgb5P9bza1z8Ht8YPXLM7w0nr76h7MWd5j3oOYZfFTg+6UR2PqbUxGfq
3ZhdqwrsqBvV3qhCo0mddY1zHfMm4jc2tiFCRe5guuYo/1mNQo7mEElRTzjXtcSI
rwY1Qs9kNrl8V0VyGjl73K8tjq7l29jXwgZbE813rEfEVQTToxccoDuXfuralh9a
aM3wVmWRCRjPbNSZQAoc9II85VtCpKPzUjdvCFMl+ho8M7sAWpsySJ9xj3Mozs9Q
2KJnnvWkwriG2olwvW9GQIIVkhqQHNa/mH6sUfDB+E2cenbfTYK1IVEAwMNAGnom
a6fR8MDumSmcgx5kOOVey4XnNW7+xKGxb4/zk5tGfB4EYWHgmEva+npEz+q3Hzq1
smBaxh/paj24Y+BjYowPIuShf6W6TtahgA1z4hEMRGFsv+B0PJt14CgzftCVnXwd
Ct+ozdPxyiSe/D1VQsouXZJcOUrzHmDGLZU8M8dfiOWKX4XIz7gTvVc4IGFFxJ+r
aKRNEgOC/12kiCjiysnRSa5OVeHlbbbL8GliDftRbx6flb9A0Q0h6/9G6p2STagO
k4GUCqtN7u9oOFKOg0xAJQWjBAbA0mPMv1SgSEBpwtCmega90Cm7YdSW1y66YIzd
xZFA6Y9FLYAX6IsDKMMaKZziJEyO/28oSOsoxq+yqndJS/6zEat6mNn0h9WPCoHL
IT1ER0fXtKZYFDFpVe54oAdaY3jQ6p8EKUGU7DlEJupkwl9lyPXRTsLoX2VuuJCo
wmOfzmFIlUx/GTs4BK0pebN2VEy42XmZ0fnN99gji02hY33ClBA3xzzupJU7AGqM
zeiLn9ecdzaYo4FIcm9YaztHo0RkhFwbxAFb5YmEjItrwUum4C6v2HAarGFeR7ag
IxLI+xyIwOUfFBmx0HJVC57D2RmAjERwv6BcHlHALJfRGrk1N17qcTS8hNI/nkQY
xKFytND2dFE+sEJ07tBwY2UoW7W7Rmo/0Au3MmEZl6vQ8HHGmaNB4cH9SUEUXAAb
gx6kI6vFgZ16qFN2PtBIbxvZkq4UXlcdvefdJb4kQls1ULYHTAlRpR1ui1A+OaQS
ww/zAUEaevZTV1jaCuq+7f3UxPXvVd99sH02G5xGPxHq3aLzIvVjLmlYytzQeUqF
IIbaZBba7F7mADwfcPawP2LaMZO53Lwx9DraG4S0mFT/Ij4frCOs22yavV/zXJTW
vX1kfgR4K8Oug8RIxPyTMpUCib2K6TU69janhxfFHZVOAfDuFyjYsJxb46OWftgU
XggXOZOOeZQdx88TUX6wdjwciSbk2NyaFM+Bs+okcQTe0XmXNC3dVaC6vkiaMJ3r
SCV5ZHDpHpFObHBIQK1ji0c771AAFISkwSmaAWhOlrDi9erL48vgh/iGuUtvhawb
2if83sMTq0tVDAzpRRq4wmKgcZl0uJ+p2CChGCBKmMBbwsy+Zc0XmGKXfjWBf846
tAYQ86koGvLz11ODY+WSmVK64nKyK53Q+u8JR53DC+y88cVJQU+NXHN8SfI5w0H9
8vdPrC01JKBzSl+6Aj3PqIUs/rCReE4H+NL/gQtKaz3U7pbvcU8Vo6szr3UMqfeT
+ZtmlVHRCwRdMzCl10EWKAhwHInMFfTr8H2RTqyBhVLH5tRvWFsR3eT7FrJR3l0/
F1CX/qPswMVbBTzm8iprMmhSjWOXghLkci6iIOKZUIh59ySy7QPqOo+ghQ+WqlzT
4EYXDjYXDzpEfuIAE5Lujbln2uk4CTCo+eaAwe5qMLtQzSo6bY2QMEmNoMhldGs5
j/p3shbCDmDVCtHaYCXBjp6nnU90+O1xwEHdszPT7PoIsA6A0rJ/kGpC7M+KfcuR
setuFfjL3gbbf81/RPFeMpYS5JPpy8kk86egGnJnkCDOLV3dOgNP3GVqlOfNdKff
cK/IAUg15eU7JJ7aYUOEXD1QQonMg4254JDOvov1np9snqoCdS0mKT2CkVOejPhi
+gsqV70qTFnzYrY0UzBUOnL/gQlyM7sidguNk7F1VYdPsrIpz5++w9EClT7FPyqR
D00yMeyLgcLFLv8HdoriW1RRmKLrbYw3L+1g0QcEqjPQIqMiq5XYLpal/F/ke3XG
ylHwBCAj6sarzwVvsDDQR/RHkggBREhn4BT1S9eY+9Kvl9iyf2JNhgoCfP6BZJST
c4QUT+8V1gQ+jivDySBo+tBSqwFV+87A+GcWJEMRnNnMomQwwaukJhO9OSfjGL/p
fb5TKxaCITTOTTA++aLsu0CJsAWAiNXVPpRlLRJiMDcODYFeGbeQF96pv1eWQkJn
7NqCYB7WMgW8nxUsomSfUxFwgGcr5LTQUli+5vmWAFYcoUiMEXsU3W5+VUuL5hFv
CKpArwDbo02GdoODKlFkfeg8jzbx2UN2QnQDK7S+Vpm7ohwB/0hS+g5n5BXpsO1l
GZJ6H7/W2OYb+SktIVmZKz8r1Zq1pU8B6OX6XjsQ6fT8mDVGljDR/3B+JILCNnve
PXxxBRlMfWeftf+jLRpmLe9jdAY0YDCV7LEgo30S0v676HRwAYe8SruQJEYe53D4
VYdEt1TMTME2Ge3u2csCGwDhpdq89tdPcrTLLB8iHDTkDo8tBV+HUY/0t2u2mluQ
i0GL+I1pUFHzPjPiwl7kaLdbGMwbazOLWj1wR8AnJi7ZSiaajW5h2GilYUTVJDxB
Yj+7xjZfQEiywh923v+/F2y0bkHoGzHjBksT9fkj0tXk0XSn3E9TNnc7PS9cu4hF
U0/1xhtQAjaIl7db9kG+WFVKYoeAlVUEmq2DibEOrpnG2Z18k0On5ZLoAQ4Fb+hp
hnxMVu1luNK/mEXb1AJXJF4AXwGcNbTKHt6S1aW9AfMObN4N7J6K94T+rDPimHRM
L4z0bx7z+eymexqFdCa7nob6f5nr/cQ3RESA30UWL3/UQxZ87vxAWIkAU0PS4tLp
6JtCUfljCe7gMzy6Cc9NPF49u7y/BCigSB2908vywGYcpvVmsroEpqnFPwjNqM3t
JMckuQd6DjiVrwPdmh5OpB01q8VWxTePYmOXCVr6TRkXLNHcd1Zo2Mqw76U5huCk
wurgGDxbgpkDbfXBSo9V8DhOACPYt4z0PjC5Xj1Jx6iaW68BLKxAUJrUEX5VUkGF
McZuyAN7Z0enh5dpsf0kFS6E2Cm/OYvLCRU3N0LYE2TlFhkdavhWiRuFpTCYdva0
Eh/MLHVnxOqpnt1pCEb+QkWojFq/mVt8PTFZwV5PyFdc4s1UNlR5w4JPVCUJjH8F
9N1QDn0bge9MjyLBdHDSQ/o3KEOo/85cKhZq1KKxxOdJ3Xpsx+sASDnKCU3tH/Lz
HKVkmVfCkae+j5OvZjiy0gszWRoOHU8kodY8Njhbx73l4r1Q5gaZl/WGkQyqUmFL
1xUDldRS1Tg6XPBh5s/pv75L5W6yo02kmSv1xXC9WE0crqFrJDKLnNwY1wDekM0g
YE5ZVnCQsgA2S1wEPqkV3N5OyAdo93ZScp5EtL3g8uiTBu1MlZp6qFuxGZ6l3f15
ZvzxPM/boDUh/97YEuFDhnD7ztb85PfYnpv1bU9nY7cRwrpIBWiFy8nQp06BBfUV
FhF4B1NrP2ca7/VupacDxS/RkAHvSeWn76CNI1X13m0ScKUtG0Xs7IwCClbzCTdY
4FwgKQfg7P6VCGPwyw/4sK3Ke1gh5k5hRAweOqVqwgHlr/eUDXNuMZfgLjJwoq/M
RLnnX7znXIDCq/Z1SumqX+d9HJoW5W4iBwAyq/Lq0VnIwpISR1jygyV4K+EKrj8f
6BU2KhaviMv6HLf2idLFW7qFdkHzHukWzhRi62bdYEK8SEd2Siuehexn3+PgSl9u
KUHcxyEle8r8ig3h22Pe/kY2rochnEfZhA4K0fbmT7lirGJzBJRq741GIzoZo9Oy
TSOkTNyAlkxWldhX6VsdcsLmW2gAGXndF2+iSIWULkDWAIZXJz7EowRxfPAyx3/W
rqw2MIjwk4aPlcpyeutgn34qt84rJdZDWPB4My0KB3OSJ41aQGYFNs8s4/Os2pKN
NNHIQWWjZMDCazZfCZ/IBZbey7SZXX/LBIZyPtlO9iMOTMMPOhOGY7/UHQHFnIad
xxNkzCG6Hk7x+XOaMT1tgZBQ3J0ZdHQgaeRELlHp+WjgGmhmKaV3nPZLYJEfG+5t
+F43ZqkhJQkQEF8FUAlIY8UXSvg+WGPbbBWhxmPcE1d1h84iOXSqLVytfqv0SVOF
uGF4xeIGJWNvo1QsG05uDh9AIz99qj6SRv7NFbBYvfSwQhx4aVb515bLYzs6B+Zf
67ZBDTjyLYE14CbZvFkWcebelYkv/IYSqdZ6HQsjmwF9WlAhiUNok5ibWehIv66G
jXz9KpCiPquUfIjeYXaWbted+3t5jVKRE/GdIp9Dn+1WW2jIPDxTXEtCXGAYcul5
Sd1e6y7CNYlGihei1mYPUEl/Xj5KVznXtF8NMAbmO8DN527uZAM/c1jlfTinWx2a
AfB8dw1j7RnqLjzFiq6v4BDjsYlERXkXu9BTwfbgDdhR9KCbnJnupXcDabxRwGk3
je3rrUv2Ef0mKzSi5tL7Wp4WxhRxk4ULSkf2B+lnQ/0CgPu3w1vQgofR8wGlHsFn
yrF/pMxJf7so1iHXpjfhNIvf3Vswqab7TSADWVGwRWji9KqdpqWD8cPxhsRRL+1k
emgYDqTddtAXfCjLcIREOcdXMFABkHKViRvBMPZR6xbhq3EbM1FHDPSAGewYTXqp
84AbcCk4aChmvoV9UX07X/TG4YA/r0GsAsf8k5TpfaHyplJTCHiEr1QHd7VP4XWg
MLFvJwDtVRhlyYTVfs4qebu2JGEO8dsTsL/U3jasIU3lwEbvp0TtosnRl+G87gKk
T/opY3vyhLwbrEyDwAf2qmJzQMsUI91nei1jc75txZfsqV65Q2mTbbaLeCF074f7
U7UDGXUJn/pc/8Dsr4g7UoE5un1hOcHmNhCHOiFWyYrJ4uPbhEK0Mpx/qlFjZIzs
N7NlKjMRoA9j6+lK3oCKn9qR85U/iC88PnWdY15FZ1ckWRGv/GcLGvJ231dTwZ8+
TpfUNZQ0hqMNXTEBwWIq5DcUJvl6s6Zy3SrwfdxY9LpoB1NCViUDphcz8WbwiOwq
Ag1fL6HAUGyNvtsVOR071zde+R7lzH1qiaf6K9OU5n1pV8YsGvYhlZYTTSOPIZ7w
/15/qZn1Ze3gj/Au7cP8aRYl5jx5I7/xa1pH9Sy3ALJcExXwyBONUlcLkOdSX8hS
GHatnHEjuc+K2dA9XuOrvRjBlrylWrqLLCi3zZ6WB2TW5bjPBbLYGG6nIlm2+P69
uXlYtIuyZRcPrVagFBaLCKhz69WWzjGR6n4qXG4Uss/POU8/j0amIn0gZOTPeO1z
QgAbjgOZuOwMj3yiXTK42x/9mMhO2vm0NJ9qybE2QkonOzN8OWFRIqDMApRn2Djx
msewD3AE+LclXXNff2aRrkv+l2pixXX9zX+5tXZwMWjc2hMiOilfmpGs5lXeg7ID
Mg6fmop+bfdmRl44Q2JYafSESOX6RnEoNybXTG6myK8p3hMTCCR3mXKx1U1eEGK7
iDteeR/BTKu6lyLcbzNxfMCBPI5K5pfgaLfY7PgQmM0RP3TQW+gUBvzprngV8q4q
xWIbMw/S5RQsNS3CFIXAv2xDIQisaOPEGcBdtmEMy1f9gnzrNf6sepzBAK9HBXIy
YSHAPsmFy7SqrZ4EcDl7shcQsHCuRF6VUePXBaa5P1s7d1Qvjf96l3sNxml8efYu
oERKlPU081ttGAzuPuLL4zow2hoozvTIdcDcapCPd4n2RPqJRpBn9hSaHE+EZKsu
NC/kqIV8aIycp+/VkXc/8VSzX3uSmgdWu9mcJ3LhKXAsEIe5llLPrj03Rz4inkGD
5+4ua5EuH9yFBrfcDcZkF6FErPCo8J3s6YuLhqNnsEIbVsawIlNIQ6uEeYidPcyI
Z/b1je2A2q2U4FztRw2M+JVQrmk5w2tVhErs/X3K0en2+xUWvKkUeWJMCxrJbYMc
EewlvHkZAZkc2owzjvsIbzAC5DfRNXmybPeluIWwB6h34el7CajhuNd85dETIVcu
go6ftfy65FqmiKcZV0w3EyyD8JLuOSTcOsKBMJddhrzoSRVixOtwpp1jN+DhUvvO
cDOPYxlSF3pn1V3gtOF/Lkl+G9YaFGj/wfAwhm+zKD51EkXfVl57TimeZiBzFBTz
fi+kpySYc97OUrggTCX4JSCgxefW91F20+Lk6WJTMgLhxwwXjLhE6e8Hs1nH+rN4
XI91xSOlGwJC21dLzszdtsCurCS9uxlJgnxvK7ackwpjJ6bPXmPnyG97veKnJjY9
zCV3oNhPBX16oMA5+sNMY+u/Mxeq9PZmn+8otSNV9uY+CXnFmrEf4tzbm1um5h5d
cPWOgcTr4SVIMQpuxswMQ0M/6xavAmQFBWJ772ddPhvxcXQHLkfDT/RgdEhDYB/g
//y86z3vnPlS/J639xoVjLLPA7a8upLRo/uwsThtP5M7KTDR8ck/7UafjLGCuy4w
bV6Fq7eStAWvMcKZE29svEJemzlLWknCHIKGpfXGS11g9tSlbYzYzhrbM7CSZYc6
J83dAH5ti6mb45MWzb4ErXBp6SMQ3ffLlDrhNb0pZBvIwAZQ+Sfe0GJgshG7tj7l
3Cyoy2QmPNzGoypXF9fkczpk8ha2Z8R15Qb9f7KSdK0SlVDe2VyLiCriX3YAav/5
KCTNoboETjoZGWBLRavcrw55baVszJ0u/f6AIYO+h+6u1PBz6I1Hardd6LeDZfuW
k1X05kxXgT1kt9eexW9cuftJrt0HsiqLrowOcPd8kTj/I/AoANP2gVJNwMzSsJDV
zhlv6PWqkYXtfa4+hs7Jl0TNRPsfZmVmRsyL3XjjPuvVIvl9lzq8zWn8JTG9Bxn9
Z2Gt5KlmYMxmA+A7NH9zTy6qtxmxgPZo8v2wsQw5sGCo+J1LU+O+zCTD2AIcQu2w
7SMOo4xvfvt1QtnXJqArl04OKO8/CNNXY6EgCUOeJ90NaLvsPP2jZ0QEho+HChY0
zUXsEjp1n+5ZApiEnKUEjqeoD13on6ADWs+vKGPkYKxcVvl2avtQZ5DI7QRMSC8l
erlwmL6Gu3XRTyL+OlLIw5EgSJXlMunjSekdXUiLVZxEqkPwt0MZ4GwzMDV7iEHa
uHTj0Dre5VE9Ju44v31MurOS79zYErUpZ5wSNnYwiI/3rwC98zHZiuGfWDOoMQkB
5HYNRSMhHEy08gJ9fWekOG8qUCapIoaQEfv2GNvEp70yYrd69kmqMwVK60hBry1g
IHxByrCNgRFhEvt4BiEf/oU7WXhnmPJHDSrJbc+OdaPK3qShdW0N9+gyqsFywQE4
bp0bUvfMmOdcmqr7cK0qa0rRO24LF8Ner5n1xDGDUBFMCE0uc8qIxA9zzkrOMi4S
zowHNlCoSnj1twe2GoZuZ+34FySbKQhomTIK5mQoUx7LDfkELkDZ6kGfIj2VDrC0
y3WrB2+dwsMFKf47QtSv2w8ZbnB8DpNaODnnHVeGpwGPgEt8OxcLL1vX9ytgEqgx
OtRk3nAKIyZjOen64rGuokPI3XPHWILnTbJYC9vOkbso4UdR79UXX7yOZ1Kvy9M1
wUz9t7wzrRpVgAHeitm6bCURcoTQ448w8lsz7iZsWsauoU2oMR48gMCFI3L8b0Gu
DTBhE3YEeg7wAHPFT8DfMrCNabhLdKYnlQh0x+8RaHNNa7BONFuSH/YDfd65ufQ7
gnzFjMrFXCU4GOzRxRuUNDhmNkPYV53bBWonQMc8HI/CkRd0kInjpihOn3uzdrhC
lPbVuD3LDiY6yihpKp6W7rIjs+7xrxWNuwT6Q5OEByKiJXC14qNQzNS09pR+Ujld
28X7RVGN9i2TJItnyXo177wbr68Aqynv5KYlaT6yB4UN/oGkvgWbw/1mMHXvDHg6
K9DP3PJgkLOHAw+xc/d2tNqIDMj6YzfWJztlR/qAQmy3s+SugaEP70udSB5hVw1T
y/6qjI+BCI7L+XiJJZTY4uAf+ksqjafVSDNja9UJg4kSRdboqL8Duu0lXzh6RiMz
1MjBOs367rE7j1iGobUxZzJIwe7O5dbGUez+viepahq0Z1htH8Qel9TR+lIyWZJe
vSEXh+HxORkr6UrYsqmtO07W/rmp7VffeC7fIhsSg/OjVsSP1In1Vt+isSiTv0NI
rdm5fomIcthiQzhrYV9rJ1mmkDBH6lbPBMo5gi8bGTiWG1MrehoHddSqelThMnpn
rcJO88Q6NyQt/bzARfchNesc+xHrH5RVElhlCUWzRKiLAL+nggUsx/I9AKiLMC+7
MZnEKmK1p1fl2QfmtQ/2m6ipX6+JC3esUC8MoW8ipaEO2BgrD+FPIdi/24lfGslX
dutToVyiN9/12GtUFzsSRkRlacrIsOoL7TARJJ0K0aZW3s6snMesxaZy8VLMFmFZ
UsgcddsHTxE54KWvnSr8Rcy3wZ6zzdSH2ZkV/JSIa8OdWnXLvCy7YLpwniDkHxYt
VGWrGgNU16BGtXp/BvKrRKtj1/hauZWlvmZxKz5KWNbXxejy2ANnDqIwdCUSyy6Y
gXfhLy8vs60jl0LjJ0SKP0NTh9fGcL5jsyNVC1YDr1KgY45+emc5i+IwUnBcUg2b
jVwjOKlgUG8Vi8zF5rmkUKdgXugkg6N96jq+pz49HOEdc4YBgcf75ofDVOWA73TN
ZXcFbPWLMvE+YnPv4AduwnFggoBJWzE9aaurDEoLK9nnUU/TdQVjpCwJCfk4ohFe
4iN81T8VI7aj3ZA5164NDybF/L5sjfio6cVMIkMr0/RFDxecdlsX4TsD1Yy6k9zh
ud6mDKmNMFmum3LdjmbULN5lVzSnuAz/1Wkkym0f3Mh4wBLc4fZNVTe3+a+U31OT
iCGOOA6cz7FceGtbBJxFuDLDVeK4dKYd7wmF//9pDjA4Z8xIoqGz1wpcQpu4tE+7
8ed6TOSahbFYAp3msVa9rfhnz4qSTRbeKd+XE5uJeb1uAd3lFnY6Bwnqn38ACBSz
fKP/1JfYLd7pzlT+dGyZyZ7LP6q207DlLYtduAbySB2puvE+rYnKXsZX85noQqyi
HDEBBHfc9nd2H5m1O/GitlJvbjoLEn3n49NeKy6EpSWKpa8+b4V++9biaDFrXHgi
2nQRXdRuT97qIDgvW1B5xyHj5fyCBXZ0Bz7YnrvcXCyqDXhd7AyUDVE8OIo2fzUy
O0dA7TieZVg6v9gBx4PuY3+jnHn6jsAwdz0t3ty+sZiGPvo6nBToWyjiOVlgU86B
C6YOC+YxuvdCBKhD3XbLa+IbGgtpCEXCHE/AZO/1B3NVUQHZjeHLCJYWCBmUJY7/
OndE32RVhcge3prcIdQZ8rVbu0HY7b+2H6d9WT4pDtaD3gW+ezUCw+DK3M//dsaG
gynl2DJvhzoiAIi+IJnSsWuDAQwP5yXWv06+i58Y9llR/ZOgT2K3w0+Blwkt9Cbz
u72nXNvLUiza7aBBACJ7CqlYB3oZHC2qgKymrsyVJt8tJDgvDvkGqYa71vskpLGg
7Ti9u/xz22MqbP2BIaPgtrd8DEC5BshXlWFqB7h1Vloel19ARJFTlauGjVHQsRrc
ljEhJTaahy+awajRc6NwIrxbmrAUTtE9jgFqY67GzWUpw832Yd5vUAPfMMHzOYYp
lYlerVK6b8akhJSWFioC3iCWJLuhXE9vGdY7sO51wvKm9Toc6WG9IZeB3y/XI4ZE
/zVz+mdLg206PVYI5OAxW6J7nT6Ol9lfdXhE5L8meO91GrCuAqeMOz+QX6cVKMSe
CDZ+tTO7d0Oyq2R+naXHyiEHe4XX/SfjJBxg0g+p58Vhjae6mBzXEOp7P0kNYoll
AKJxkkDoaAmapKdm+j2GoQAZP8lPGbBh4rixaMb7rWREpaWkohD9xJmQ3QArJL5A
49SDojfWjWjUZxxSOWffYLYwAngbM1d6Z9yV2g4SCqJFApE5TppqvZoPp6wfmloL
FoJqRc5izTogc8ZYqhzW2yfiMeE3jIO4g/iY0MvydSAi74X1vIsR9KkXChC+Aofb
wAkV/aheK+MaMTb1sC+5WrzcLaojKyxxJgKJP+T2YO3XKK+nQxBfJ15IO+XtZXW/
GmKrvpPS87W6wL/hgYk6aBH8ZeqXLitfPthqoLaRTwSmkRjcIYYNAlDKJTdSq3PC
bTztLpLs8+uOFQwpQt5xm2kesqjs2ZmZXQtdWyF+keoOt6yX5fmSTKrF13FDOmYh
bFpMlwBnoPDeMJMycTe/5DPUNcoccUdgatTb0HxcCPzwtSCFXM+8U6jSjaPJ/Yep
6b5B8IMyeT2xhT+WhyTdIfztnX1OHv/UguBKT1WwHLySaH1+9fKvyNvyHkptWzby
noxRNE69ADEOnYKo/xCEwGPTvWAA4S2nzW1hR16YeJeTeCkmzlLNDo7tqyjnVut+
i9RZeHnyXgaXIRcWtWuDcg2VWFmh8up7g3Whhf7iJXSEaGEr/aWFSvc8tNI2KGXO
84i1EaIMjFlf6vEr8gaO/ScAtoTPpZD3/8KE1K4cnUZ91bwzlHGzBjUOEl18EidF
U/MmA65F24SZd82dv8QtPeAw6xJkH+6ojWGkjD6nvk8eeEg9sdYG7V8Zgty7MjAU
d3TJxWffvi04/FUOgANdh2R5ienOcU8PJMwdWZbeJNXCuqnNMLBxI7DdVY7Tz9wj
HsrrWkEOwFGoOACrHHhyewGKKX9/fEdawbQR8zcpEWUFvrII9AFDNZO3ZbYWmAbE
kpMfqrKIh+3CdNYCDhRH4552qIeQ7KEHd2cyP+zJJJ5M3CWK8u7rHGCfZNn4bR5U
qpE5/5J5+r5sQrakCs7fwEXr2dYMiTZLS3lfHrN9VnMsM8aeRJprilKvBa6KiLmD
C0ZrVb1kR69QEGLlfrQLSox0osHAtwfYneaZFm/CddmXFwUpsvIQ8VeR4iC+FIwp
ONe8nbzSI4CxhPKZILhAgqySt7m5XVpDXkmKVT1DB+fFx6n6IErRNKGY9x8BUYKk
6klhkmqRsk8MLMFYagWAh8v7SSv677Ckv0n3qMg2ijZX3svrGcyi2G27QsGEPpl6
vnT2XT02p7+vlP42Us36t/5GjKpxKhv2f653Q9GKC/Jiz97i51RRJtreCFVMv49C
1c/kF5WXCg5PT++ELsWZ8kiZi6st22ZDpv8tEDAkXx0WgmhsDguiOeJFJHR+8ZaB
uDcE36UfaX7rikzvLeZhHjeCipLeochoExtg7aAxkdJVHRQhN3KaGySDp8CWEM8c
i6dTWr4qAyz5M+r5+/Q3Rnnj+5HnjOfWnicI8fED6gJHgeUi1755UG+U/FopF2ip
EqRbSlTN5mI9Rsng90R55ODe0OyPET3IraVcb4WzjsqUOWEEaA/uL24X0cirOERs
vrNpZAA3DDWYJCJAWdgbvlwGdpwydw+WD+427G6n0cRbymhBRry6EZmVTB+tKJa+
8mWVH6XcZoKXkH2ZbSNDAux3KJS8LmAEHXwt2H6K684Ow9uUXWJCZBqY53i6IPhs
goTTGkk0KmEdLjmfRP0W8yjzUBZSaJH0x2sZSnwuPjJ+H2eZvjsjfMW9UTCVYgFK
/W6wwFFDn4fW6KhiGqc2x+Xmd1a0Rno+JjM4VudNa6AD0W9M8kEgdCb/WBxn3t/s
5xUiOsuQG7uekXwOlz4YZUnA7hrLfBKfw3BPsla1K8IoOSbp2HH7EZV7WTzI0I5G
cX5Sy3zkqkuFoWX+SoYh3JL+OmBP3H4h5LKrBi9qPy/yhqBFeHyjk1c3PKeHkzfR
2JwHYJqHN32QdeghSQVK6rnI/8UbpOjG73fB3w/4EvIYjk7ijybEUB5Suq9ow6yl
QJvR59rHXt9mrplqXcUE7mwCRzvqAWU25C09muLH5b+dr541flleCcMvwUEzImGd
XjgWdSxV71RMqyInRKHfu7SBtNaqBi2SItQrrx5yFv6+YXT0vB00+aONR23D19+A
UpIVxp4Gs82lgAPst2hXCrLz4st1vBb9RXrlLagfUEzfBLL/qAYgIYiqQcfFFz7E
E+nQVIC487sV9fjgLW3ADx7cO5/8uIvfAjTcKkkuphfBtybuoOhbxm6vOLww41hy
MwMDRXM240cnVdfdFRCLPq4PILXSksrHwzpedFSrC5TZISte4Ss7jncw3l+QJTS6
WwG/Mac8cri/0KkaNkrVTln0pI4yKwF2CyBsMXcB0Pqkgq1ibpUW9IGziuQXieOB
0R3RylJXXbUgv/y7F/0jJU5IuBGJgdQNS8Zg18uLPInAZlfgE+eTPb0v6pE0PPP8
ttQDHL3hsXYtIsImZuLRb4hrJh02LMZi++KRJ7fdv0lS6c2XQUKypil7xweGKnGq
SsLrhNCyvUKjNaAJCD+/micGdsktqSdzQqXdBkKdK4wjmLQ8Xm7gznleCpdtvJJ1
YNpmd91Bl96adg5h77q834cuBHgYNHxJtrig79Q5bwcESpCkDghPewlCJOSsHrBW
pmpDD8VNghnoiUrPO3AB1DBmF/U9s0sHdKrX2zTM3lANstf67ED7vVS09MFdyADP
2UebMWKSPYsfuNdn3NWMDsOgFOrrfVVlADm8JUh1NtahOfbLMAN9TLxalI6WWpHj
TnUrlEH7Bz56tLHTEgwrBfpXTzE4vgAN26D34nLNJdGc69bSNcb1UVZFOgkDmYlM
dHlFTMqNM93/f0DRu9pYf2l7TQnWyakIRZKOdEbhuDBSdmJ7TTHp9aRzW1TMcmWL
qzzdgnLU7koAC+9dNl9j/fMAe1tHpjJdBxixY2XWXZ5JOGgmcfYWso5ibgcm3/pJ
2OqcJ42FP5XFuGM5WaTQoGIa9uXY8ulEz80MIIKSZAW9LyrxBkhKt8hp2ZPdSLqj
GQUN3zAWl+lShNs2dTilZQVcWd/d8nuAx86mgqnvLixsXxOwWxuh/I9ZjniMqap7
vwGxHxeq7tX13yxYmj1X3T7yh/FT9o+kw4cHfy76Lm/vTl7QH4UoRAymJQlVigls
IfV8JYlwWlqzVjMPNdPOcoY/7tCmzyEwcMrNp1F+xaB/rM9zBZd0X+i0RMKUAPsX
a0YS4H1bQ3aSxDYB3dIa295G9aozi+c+QrFi69AVtADgBYsPlcKtamJedl1Ms2/4
hgMMDmbtRrzDf/2m45V5jUpUrCWbO8RUqVCIMoV7Xisxx1mlQ1PfjNy6TNuAbtlp
8OyB1YSKnRi/TautISu6l9qxjYAMOWUsJPGThzwNzG3XWJKkAw7eAFbIAVRGUxv7
Zqs1QsRDJMUPth23x/qZ6Ege3xnZNCz6uZDDJi8oU8nBbApC0DSsS2dLtG4F2GXV
PgAXbdI70lHQIGILE092D0zvfGMxr/prUcP0LPhomfZvXTHor50aL5vZg3seWP05
HauzZXxlUY+25KjDa91xQMfoo8JKHjowOLVkqQ7ZTbdqJipBcjQpKO6xivIrOM10
SxxsLtz0m654bYfo34OVQ2eeFRUbY0jwFfmNWDkDDTNrV7iH7CyGYMEp57eNOBTa
FyTmS5cSiL5e1g3R03dLOckOihLGh+z4osbDqhXlvf7ctNzSOQSj+aCjwIqBg/4z
u2ajNjb8uvIkHkhRdfJUGYFMpX0zmEMyV48ARlF6qv6IC6OpgzNlmLtSAqAml1hc
kzs57+P915/FLe8msnxDlGHHj1w4JEc164secQJgp2mOxHH7A32kjhW33NiltuxW
h9PtwhItU7+7z10IrKxxUTeamAar0tvZZlDpaZ2v8GZoTYvv5NGki5apxMV0rA4X
ub0i88Z9yvtxb7JqEkMAr6JjwWumnkveOHjzRcMhATY7nOJ2rGs8+UKRkj0dnP9E
GOL8O0cpzDtCWHWZVrE1/vWRo4xki63UmhenyodH3Of/3E3BVxZ5ors2FoEVLRbr
aSkSdomfP49YpDIsladCgtWtKdFypXL+37Gzu3eECPlZHTiTiFpyXfmXbK3RcLy1
mWanDqdfXX7qoSrLuFISRG8IPKANRa2TmDo/RzxEiJaWMb6//31GSwve+jl+Iw9x
tqe5/dqNU48ntnZr/yreNpjr1s3WLYUsRCYHT5rB1VEarWUfl7Czyl/VEpwIIJ4D
cztK2Cr+ARf2tEjdgEdix2//mtta3d/YE3Yk428IdATV5f6ljJbiGsgge/lfyJEs
dgmp69/4XeNkhKZkUnnFJOB6mdqQpmUq7RBS+JNsdYRSG/wYAKqttEWPbavCVNPZ
fPdX+QlNa1bR5kEtsbuvt73jCe+RfHtZEZ1BEO7N6ev45YlSAU8sRH1yJseLQ7M3
AkeQv2j3JeMrVzAp35lpcCOnk5b52rzbJvVIGFqtcYfIIqBeQqVEFQqduDNScHpB
Sd1+GG7vypSfZqofnomCA4l3rMxQij9IesgDLYplyS0lQSrUc64F/yrtFwD82Zrd
ixMNBTGO3SqlOGca6Bgbh48bWQWsvKitk4BjrkZHCkBYAyjtx58Ce3bRQolUGr+0
fDvO/zqVosXBv0RK/tj2gifDy3Eq7TX6S3JXYNs8Z2Jje+9J8Zjg657qrlPdPf1g
dwI/wu2rBDL/zziHOPjxVVpKek/6T+AJTlwcIcf++F/JQGVGTry4EbkBtOXv3WTu
6i7Q2llnQ6rGe98v2fJ5sljCAwZWEkMg0IdWMkJjCxrs5c822SP3gFNb7R9cMHoA
nyS11QAQgdXyMMdBlSIL1DJ9qn5EqxjsaOb3y7YTi1X140y1HclhtWdyfRjRdkD/
dilzGb5M0ZTTdAyrg7wm0i40fzZBo7Mpkv824tQfk4p0c/yoc26mO/7nojMWgzEJ
V0jxOqu3d21532mK0/Qbo52iJQjJptu7/upwPHqG1Fy+ALQz0mZvxuNh+ZCvyiLc
VTtPQoeHaezH7CRHec9QR4pKOsxo4u4ndhYEqP5ROXaPmuC/JW+gSRx11sRxJHQd
MQnbKVS7ddpVZgtPMSEh6XJKrFcT0HE2QtTubguT0DU+Vi71Wjbjr8FWnMD9jwX7
wbDIGqwQPWVEjXokD1a99z6cA1FFBINqaJ9QnS5+PBeoJX11wCncUVTn0RytNREy
7XOEqw7moHvJvtofD1RnLJYP/TMtHdWblD+zZQGIZEhafxTenPuMWQUZCC/ecqRh
DUJreJ41/YCrm0Z9CECnI7YMnufp3cWmFy7yV+srNQ7CChBV0pAB0Qi3+8ZlfaWG
vudx8R3O96PnMMeIqLedMWsxrC7sqR5vi6eXOv4s3YWHCB2RlEc8o1c6CbrptaWO
SNVmUM0UFxTyhXMlKQkB1hx0OT1HZbNZGbHPHSQXh4o9gvk2xwf3yLTXVzqp6k8e
GuZmRMXMiZVXnekfaxrmyJa+X551ASK1+MCoF00pPLTLtzHA+ImM9hSmaYE8JoYo
5JHVph9/NJmcvk+xZgxxQCgihdf/AbtC//kX8TiZG8KeBotoFcLASLGBlKlwdeZb
6pPT18/JDFM1gI+y3lakbuCjVnlSqOh4rabtQmoWuYYKAmGj2E2GGJo6bgH7ahzC
3Da//72mfaJ8kXaMrhPZkUUs3xQm39/a3KC94vsD4JMSfhXXsIjkyCFAWjlLy3Go
EH3N+k3BH+c+yMtXjFMPYNvNlYsZYhNUULBrVnWjeLo5AIO9knATFkBo2RugdBEp
b7n6YKd3NUU3wzC/JgsxBXA18sM7V3XgRN8WAPOi1ABnCOyc6d7J32I492n5zNkK
q6r5aiXzqpc7u7KZf0cQC6OKazCeU+r61LQdHnjdSKymnCehS3jMjmvptQDvc0le
4dWGjLTlRdgWP3ArJatJDSbW76OQFfnE3PvHLfwbkuhkUCpjGLeqEJtsfocZE5UG
TlyJvH9gQbWJct2FCo4YXYSp25n4WY9Bw1kDZCRP2Y62Ym4FUqaKWLIcNnY9D7La
Tlu3xwxt8NFq/BeQoFhCQJ+7jFgybm0cSYsAktmeWri5LLqeneTCF+8z2g/F08Nq
B4j5q7MEIui/oeJHE58lPcdvd+6PA4J14HzdzUvhsTL8QPOCyTRc+qMrNzbJgeiE
9OHft5OpZVlolFEM/Y1BXc3UDkXOE+0UHnNn3+zFiU7yyQrIhNEFWdqz+dZhgqj9
oHcvDd3f0OAjMUOSiQThCsTdzpC0JV5HUcSrRbaXSlD3uq8TWs40wUYXxz3yjHoz
AxrS040485F0j6RYFssaU1ilfAwn9M43y1kjyXLDzO5ljfhsawbP/Sx2385dGbIl
7IxsLNeHNh6JRPqoasKIlJNcjssjjuGwcPbokVw0I/I/Mff3ui/FIPNFvEeLfhCJ
IOTd+4BkszBrd3rIUUxuLvDY8B7Nnnb1JhZZ13aKiTqzT2ZBxP8Hik5K/cT9Ixtb
KZXIERL4i/0wNGx8mDC7qu0F3Jkl/cZD3GQ5BF/aHfUb9qYvdP8syc/KjYMgtUWL
nRumHUXMwT/M4WxtGBkJumGTePrFkZBSPYM8HYJASZEAI3ZYjTjy/aXP1YtIw8Yv
qECPsZvnhk1L/bEgBc/ezPWUdrJrUgBHghA2lmw2vgM48z43Ol7fD/EbYdTatT7e
dXyYtSj259ZWdCHM81qafGlYmVh+vm7s+odN4zTAqfNKVklqosncUu3B1y2z3HQo
/UFwRw3+zNyzLK0pcvqsSJQq6ICtcqGfL9jSu94iKM2bHB51XI6y9jc98y2VdzZC
UvOfNQrIfQg6mWu7W9W7uIIGKctz2n8MKzpz6Gr1NnIu7MTU39g2Jcbj1uukuYly
reGqRRewiwHHeTroZMaRjqE0JgcKSANbwJHET2WxBnsbrwONAkRsXLNC9Pi55i1x
6Hdg4iUoxT5KMUuF38L1cQe6dolKPRMQ99yeeYnM/b/KI1kuae77UIucR+wA83+0
i6z589haHwMBFIpPWzBbTYjLn1zxDd8mjXBbhePEYa9bMHYbbzucKfa8uuIhVBRx
uFdnCYeDtqueYnNRQCV7I1hVK1FjUYskaauH5wszqLdNuDJxF9B4bsDHUnm+2sMa
r8Oq3pR2aB90NeIYwVxuCshxnYIMGcJhlSeAE/qm+W2yHh8fZfpTj4YFF9R2CUZW
Omwmfq7ib/y+5KC6+zXlyqIZTda5Ksw9nLsIA5RBwX7NSV2Mrx40D1CkWe+NwDPT
iUGlLLnyjOvAxxHYFJr8NNAWIY3K/OspBt4vnRsanZj1WEGG7fsz1riL56dwcuam
IcY0cb+3mZWwJFcwdFwA3c9NtcN1mNgMnk8Yw4o3b6z1Jm2TPdziWAmZ+ecK7q0V
+LsRev7KpTDdeH7LQEaxlWJdy7KHNXrCahWyijKHj0vfWXisuxkrC8jCmLSFVgaY
nUPTLnsGxilHo+DRHGgOhk92aZSLZbIxamSsy3VChh/NjmIqePZHCrA5DJmJkvTJ
WJthU6EafP6wCWibEFtbLKWGsHeAUYkTREcc5kJ88lHBwOWAboJRi+woIRuXhgtu
RzgNMsSK0y7+ebcbNOKhynYXt4mRoJpdTrI5JNTusOVtFyop/tn1Gs5s/qgzg8Rn
5c7aM5ULxG5zVz6HGEV3Yr/iCayduuP7g8rcn/cOUgysZBDXo/9wSm69UGdn/ANz
tgkxH0F2huRCcKGhvaOntY+9hhwLp5FEWj+CD+yyNpShKBfnOvScJuqJNLmjzn1u
FV0nK6ghT2ra93CK8jzrYy2NrynPYY3xJGvlPSOcB6chhOrbYh3IOoBdmoS6EX4F
gzepG81MyJpMfMZsHhdyDpbq2yVxONrE+tkY5Ziv5U2QBUKlCkQ+G/tDn7NNXZd6
t/zP4jW833cxGc891N2D+8Lfdz04sp1i99029XOAPpZgDFtXsi/jOljbS/Q3KW3x
Lg+1NtPibgMcW1yt/9YjEJAR72z9uIsYyKF9Tbuq4xRFPULMxp4Wn2lwYOblSNM8
B4XUYpnMYTmRD8eST98d/tXMqWePBFTM8wmSwxwk6KwhLuZvJRJC8GivW1YULJaB
3I6BE7MryP6EWMViEBzv2XmiCXSofXGRQ2VDBfClj5CraOVyGdAvacRVRE5VfwrD
MXqIbsplpjlpkBjmyIH/JRi5asiD1T5BwwbND2+Lal+418WhMhovBZrLVxhSy/bS
OGJGW0gHautI6FZzvcB+6MD+0lAnSNZN6sa+UYTVl63wLQlvr2mnmQOb0XkXmmuy
SX5fQw68+veXZfrHf/6G5U7iPJbC+FFfYnpLe3ssTHbtodVgSGI7Jasws9xLbvX1
VgOoZvi68gJvIsD7KuMJH8TKEvzD/Q+XwoSKue16Fy9OJCMJBhNHhsRNqCN8PKxX
NrMF4R7C7tRY+I4y+c6l1R+VlOFl896yQPx/T+Q3sgT5ZjPOxSydBXVrd0Q8y6+W
jphYsPlLBihXZRTQNVtfLp8muwWheqL1Z3lkWI+SNjfzL5+0+fj136S4q4ZLXxlG
vK15o2idscksGkcSAdMlcbSvLngriruMo753hEQ3XzUm/dzlqwS+rMt7TK9Cnwe9
bRLPlEKoeL2N2ejcma1S5y/mRnTZ//JSyHknBPqSJUp/QWWItCgLn/aAf5GmC+M2
I3vCgGiIrbBqJsKumQaPK8PH60woLf0B+XYN1KwdLfUqmxKefbmVqSOp2Xm5+584
WrCLxfa0ig6TQEB697PJCYFmbP6rWKuce/YK7Xs1TzAMZAzRaYRsuSFXufY3I6Qg
lH1YpMmgwKNt4pJE2eX73ickZpOcCM5LTfi90WfWNjrypmNwzuvu4p69WMI+pNgk
RlPlI0b2cnYC0xtIZJd6okueuhivri8qMUjNvognLUTgWw9n8LWx1wsUjbnkYXm8
NixVMFtu4X5ioVULBSzgU+nze2qaRJUVpZHha3R2LZI6hAqRYzlnnfzexKV3fB0D
3SRUXKRdy1sUnhJWu+P+Jn9mIz9vIGk6b6tsLmgWpIDNIFBBSid9cOmf03tJdioF
+2XCzXuD77OAsShjwOjEmIkuBMwS+vsDIok2lJ6yOgc1xVNbyNVBnqJiEmNY4fMk
GhG3+jSsw+8qmbcvuy3hYGWEYSxzs5SMq9XYCMbHIPK/d14qb9deeOfoEp6RrRTk
ZTgZYXQ5GH2dhzKb1KCd/3hAleV+Wu0ozY5sF/pa2eTVE2iyS9ekOMThSuBXIdfH
ySzoS9EjdsAxS179Gbn9zGuKVnS3/Hg0244CzxuHjOF0mlYEIBWa7wplBYY3G8uU
01pGSyCiwIE5cAC/icciZTCJBSzcmaC2bzTEGjbiF5tHBXCtBUIIUs6oR/cy/fW+
pBPorEmubKdNDT/n+IPOO7apGoZVxwPOW0DCMc/q6KnK4OEb5WUSJsXPyIGqTJbf
Yg0zKMZuwe0Va9IO6WccbbMdCsOsJ6V0FeYm3iiRDzhKMNfOlHOaovgI5RsJxnq8
prcvm39d72EJh0J+7oicmZtSp112a+ZWtNXch5LVTtBlZoOCa3rLGxPFwyCqfiiX
YRKFomuBZv5QPHiqCvCHH2wR2VH217aM/tmZ+wDpUlaUmEeCkCABBhG71qiDIE5D
OSPsChTxnHB4++bv/9gM1Tdy+yHbwxI209Mz99BZoGSahJlPrbmD+BInZ/Z1hlsl
llGIVAp9WN0qD2Px6vS7eg1cF60eKsrjmXfb+p3XWRBa3gbS8vhY6kurrRwpRiac
L7uT/S4S+4P6cTZlyyzni9QX/pzWCIOHu70AdMuZ3NCN3CO3bftbEQhcAdCzMrLO
+lksZfL1YQUKEy+sVGkKOuSzTVOUlvnIrKJnVIXKCpUo5f4Lar7FedWthSDlQDAC
E//gBXJRLE96+yFbDrei8KyHCAdq/VIg5gifnpNhwaQWT5ojGEXDecNiAkHKizFh
P7gYgd051/r3zp6NBQUUf9qm13jTCy58XN/aXnDjhxNrvy2ONiExVOdgTJyyfT9C
RNGzAhH5JfAP4ABglggMtlQiQSOcpguZRWvWIBHxAOCl84Q/gbt62pnbdvRYLSNQ
E9j5pmHuUnJLmEiqDsTF7vTsBZuo8aqsRQgZeL7vzk645tEpUMnlZleclVeurmqc
DtzFBO5VQRSGkZ90exPmTd6evT6tYTBPp2UKQ/TzfueoxH5jC4WLefprksz4iZWG
s2lUj7OhJDXQidjoBGX0V1Wt+VWPMQyGel3BoquQO5jfKURmFppe+5vZ1x3J8zfs
XKTwQEMHuhMUrXMOjEfgrFshJLgYw91wCgk80mcWeiWe1xEQ4bn0R/2GAeoJRMul
IpZt4k7UGSnIQqgD5F/YK6xRptGlAIgrg9/SKDLeJubCBzHXMT9ATUF1OE65nrm+
iPNXh5/AyR07atNnx6o6qbK9xqYfmVQmoWx6LC0xd+l0DBol9hHOoivmG38+F5cV
7RJMsBI1OfpWQgjVE9cqLA9WYbPwhoJVxMHDfbFG/s3jcqaOGTxbkeASlRw9A6bY
6X6FU6HTDJaQtqLUPSYv78GxgxPzosL2v2kt4X9NakYYPG+5lOMHPw7G3AY9knIA
qwaVjGQGpe+1bZVwbotuV3cLNZJOGrtwsWY8oYpM52GMFAV9yf10ZB04h+qWbKv3
RULKK7ZuaPvA15Q+6IWj6Sr6w0mf5iEPq2//xSCc/ufXY+W/ziedtMg0OJD9MoNH
0TEp5icz1fCmearUdLKqzyXRabTZisjN8CPKuW4CFu2XnkgNJQe4r9Meky6qiYag
VrRAIJrAo2NkI9FfBGKCUV2FIV5FXew83eGve22CtAplnIQmlzAKb2i4mk/CWcK2
JE0Rvq/DrErZ5WaPANGoaN2uWBXa6mFq+nuYQsOXgmDyHZXrUeMvXi22WUF0O1FN
gaJLsLq/Gew7GOLlmb/6H4kl+kiA5i5tHQri07ZriGmEOKY8WePa7fh+9eTj3TrW
boCJ8UEbg8OLfpklWhWvsrqdpGBmPOICR6YdJARX5XR+i/ul+c5nAXP/PP8EiaX5
T7HuHwTbuzmRD+Ztdyh9mqfAwGcDdgw+Zqc6uiZSiiTQtCM/97XFDXSN8HKez4mu
r30TEpPLRND+Aua8DVsVdMizx8NCVzMvkCFpKVyfwrbI/PNUcfv5KH0GRtjszoxT
rL6dmH/QHgfGk/1s6l9QH4UJA9RkufRqHQaTyxLk2AuljrwPg6XknVl9Oh/M81Ly
fCGQcfrBfI+TxgSoYrDyGIAXsTlRS6od3XTqsSRu7pAhzj2Pf2h+XccDIlRfb8zP
tFeWS/pjr2FOw8uIEyvjynLRFsk6Y+/4LUqkJUxkGgYz4Y1vwsGFrBH5KcsYQ/W8
Gvh0/nhYJOkRwDtIjQEGqyRQmnnSyuByheNJbG7b/zLXwO63cu+OVb3FvuhtArHW
JmYgc7UPdmD+WDeu1CIeadUulpaXJOLq5yY1GDVDVJV7OgjrmYFrwQMuxBZtYwY1
JwYK4/DU0DS+Ba8S0ODKW5j8QvxGyR224f66tqfXCX9Kj+0Hw/cHQcORIPGxLt1p
a75VHfMPFE/sLrJtj3V2RvlRTCKBaVJJCTUgPkZ7GnT/KUHAuoz14n3LrvwvYbC0
gn+S3v4cw9Xq25up4jolG5JOXnFuY7F3h7JB2lB4TUwLwmR05HhRaNuhaRa9SUE6
Xz0Lsl3A0GmQB/eqRyG/sz5tzX2ypSzBeCNlvnhv+pdX17wX6TEltSj+Cu8vGmU0
JIO7mYxNJq0GqNmjZtyyn4A65Y82nSTW4wSnlz2PqBHcMcug2LWGm7i3Mhmja/Qo
UXnpzQtjDvlSKB5Vv/jLIkyuDAg2QcYr0KOkFD2l+Wn59xucVYC/v/FBPLi8CfOl
ORPkX1ysueikkUDh7W052djVXvDwVoqBt9bX4+CyQtiB+egH0KMEA8+15EMgUOuf
yO5GU/9ksE8mrG9U15haMvl+KsponjpAiKI4MD8HrSZB8Uwc0aIyg2w4padxJpp0
NH7R7Ko8GTV7bdLvafukLyrCtYHoi3NTc/ZCtmOIYSYUEicEZ0E53qRkxroUQ+cT
UtxZAbSCj+yPXCuC3P6vUzalgps1/Z3WXCKo0Q3qjLavBvgBX3eE2ymymrjTisA7
mYq6VbqGoyLgiQZqAjhQpvD/8NngIqSYNJxhfygdevCcWtzY9BhDGWbNedzMc863
dh4ucqORbeNSoSJfoJy7EtRA4Xn1r6hT2jM9RbwiPsI7iVW3N6pdkFcszTc4rM+Q
3CwLwafq3xeI1e6DXbGxGWbz45NXgafhHnIK5OldSMFS685byHO/lB8aU5iu5T7f
AOm03c+oOEyW/nF+QRR+uH9iIKQi8ohoTiObbKTMJeejRqYd0udJKZ7IeSUO6q2J
vkhGvU0+98kNdOWzoBXg0jcq1M7DdJV/y/pis7BaINHDnm4EGYqvOJiZ6Xzhpvbc
81z2nhP7c+NOI/RL2ntdMvEC1JnW191ch3efw2ZseWaHbD88s14vmzkZuBAC/itF
OshjREaPjeO9fGS9zL3NhpceEiFyqbesb84WV4We8DCzVzU5mXd8zuXvywwOWlVL
5Wz6m2psJ5BmobNBQU7On0bdsAGovCaiCWBGs3VY90mqh8ohFiUIVUZ6akKeeVE5
cEof8/RP39PpfPbF5dLGPOfCTKVMTnL+v55PlH9IZp17rHPzLyWDcJWz2tT3EYXm
X0mUULBYBhN/gkr6mxP9TKZcFqMBM51AEJLT1/+FVQSt6Qsa1b98QotQx3zZwPt2
EMeMCurjYK9Q96eMZPmNsWcrGJS1us+5DGaNtWExIa/Kaeafd5kTkWAe1qZX62Ap
oAkkNK6ue2cXUXd7IJnNLk6qtN0toFkvC3WjD7sMCg/uJVUBF0AsB55ES9Qx06oN
wUI6NH/to0nFUMGQ8XVXBXMhA1DUM9SUYqvE258X9AXrvvueW8PgCMrac2E1795s
xp9DXrjsKoS4/6WjgCotIUSAzvzvaR9PsIib44px/I1UfBrquIOnBZ6JOm+xX9z4
+WZ8W9Z2M+jbTwwf5QmhyK2BtQtcGVY3eaOe6MvtNZmXCX4s64iVdttF7uIIRh8h
zBcUpV8QsaKzkqFKiKH76YzEBjUruIvPKqiBTHOSjdz8vL9GA+EvWrNRF+/OlJsi
77XqyMnEMZON8MZHvOx6QAXtV/ymDP+LjW97XDpRCE5xSb+zYMDEqww52jBj+A4q
W1qYmAtzsnPqbcm0egAqHKr/GXOIHPCTqscftyZmxnR0B+cTJS6+Xf0xKNT8qXob
CAUSIL/+AbvBIw+rz6flEPyEEMpG50lSUQJXculkgNKqVhFtNl5MWiP4NeqBzTqS
hJ3mMoBnxxOwqBujrH2Mooi6fE5CTvRWvBcVlQq7TUTcWq6tJDPoAt+K3yXRETur
RztI04MYD73EtTZy0Q+3sLY1W2kR8IjaTnXOZiJ6DuBCMWBLpYeZRlUfl7pwZWRo
vf/E1QGNebpH/HVf4mOL7kDqMNuRkf/wYlrZLdAm9lFruePPvxaod8aB0jllylxh
csBuwkLffh6BJ86k0qADqP1KStrIXqLiGyuRLn42baHyD4E+SflTtcVC6YfGzSpT
SgcIW2pLgDXgwHdmvVBK3mEqMfJURo1aE0wgI2xQnE6W++mmkV3IzxygUHUEyV3S
fnzclG3/CCF7Is2A3/DW83tXUJaSZuVPLmQSo3r7JOzpfRl+3He7OUZPNvkIMWqn
84fD/0DzFrXjMRw1As3AtQ18zQ5D/GE0PqnvT5DVMwhFKPsuMw+h8oy+L82+8YmB
YIbGFwKPQI9z03y3bpxwj/IWWEf1h1ERMmfk99/jgQOr0mZWRojYwK87V4HSwBnh
eW9kcmClIT/i1suvskS8Ja53hR3TJRv1emn186xTWXc6w82Vq2knhDXv9V9m2P6O
THsabfsK7OCIavQeJg/T+ywih4xTK/MMaNT9cuILPmiNtKtFdz0OtiomZLdyj23q
c+9zUvsXQVx4fmAZYCpHv3XdjQhBC/ahFW4+szlilp+k2KhIz4UvSihuTdAw7NhD
HDT1D0sP2NKrdgS/9RR690zXaimczCVtEVz+PziwkoEb3PGaSF/6Uok3FD09J7bk
AQz3+Q3Zy8IXqfWoXm07W2qc4/t79rYnM6lk/g2hXl1nuofxJboe53LftcYQ8Hw6
/zRcpS/+IIRt/htukJRdJDL2Kpg4tg2bYx/XFUHd9uTEMFGCKuhixKhuipvA32OX
ULjJIQHoXjkE0cu4NR44TMr3HWm4a3EJlutG0+4UJxvnz+7nte1mZ5c7INBkyl33
76J2ysPyHbEvi6EnJzcwH+AMQZmCX0jfaDVMOyZXqPWh0Yu3BbUSXL8Lv/YyNJSE
Ki8NXhTkk9thI+sqFP9VJVn8TaHWBwGZyFY3esGXir8hjD62UL38XR/9tEUNvZJB
7t1yGFVlfW1IB+yXKlxdP2iBb8ItUoRNtRJo6njymztf9vvE8kYdRpjSEWYdn7UF
4j7e+JR1plneI+KWDid9IFvzJ48zth95JVREmQnturZpPQOkUDzOBE2RnF+5OXys
CHXwuxQ8A2CKjbHK0+uVsUarNpc0FQzgHurhVWBcppCyeCPHrFm0V46awbEYZFpI
anXuJ5Jt/6QFtFN/5f40GovLw9YcoaoEjzInprpRJJh+py99PL53ONXaqnBYVPZ8
dqd0G/p/7Ujfb9228BpWhVpLCqmSo7vjd9qmBqtrRLGgzWX/4kRQRSveuBjD+Erb
Gk6gbDUH0EgV0DTGIFEYaRMfffmGmh9j/3fhdoFO9i/ti3F3xhoTP2YvFPy9Mebd
/3wI4Vu9/7bePM6AavdEr8aimk/DpdNjucXgow78R5qTA3GH/pRq9mdQCeBxOFTB
4crdc9sxd5SPaZwYdJnDAHp8YarBiEWA748jPuLZ765DqDRlSS02x1PhbJV+rF1E
tTQuVU3fiwHu8s8q6QGG5S4NRd8newDvjg0Knuruh75oEYnLLF5BfSWeyC7AuTvo
Mey+23sO3gd81X3jxhINaLhC0U5PQFgG0CWKa5sUYdQwBenNjxtFSB3jaRZDtEbU
mwxCMmHAmf70rmlw4/xehG42xPDpJwAf0aWdR8fefrhu7YRJ8fcap0gRIvbzt2oM
Lpmt67n5UIx3M1qZ+AGlfEzJ7oJxIiEueW9UIz0cqEdpo2GbaiwndV7Fn0gsICOH
H0TMlaC0K3NP8g9gwiGrZu6AyXJbHLK5/CMMDT0huumw16gb7/Xae3mjl8E19DgI
11GhQc9uV/Z0Gv6wBJaSWJwVtJ34LaWsEkhVVLRlAYuNtm2GLBSK8Zm8KnxEVvRg
IUHi477xH33qqUcsxTFi7HwmMOcpgoT145wNBlyfd+vYspOuNs48tty5auc80KAN
AHacPqPs7Rhx6t6+O5BMsN0jtPGe9xyt3r1hDJ9+DfdtDrrAQqGBtpMigAV0Ji7i
BB5dsAi+H112h2HIoFeymnGG5S59n37iRG9TaI5QZJwPc/1Eezuc9GYIv6r1Au+V
Ro+GFDLyR1Oh9Z8Y8mfv4CyX17U8urA1r5z+VT8TojyZHOZFM40q2hRAAjl4bIBR
u0jtec51ryIHtmbYG7YqIYsV7+uA+SeI1m5Rshril+cpeM+yx+kSDLvV4ILydefu
9Q3+J3ZDoUKnAP1A6XNxslaIG7DtWMRPAC3FBdAZ1j/WTOdKuz0pR8dKj/HKKXff
DaWrakzFBY2WqeEOzMWSNKxMIz/z47YlnH1tzDeJHYO8CvIyAPnumhA1hQOjn5So
2xlyN4T9AaeXpGlJhAM0+rkbxJ7HyvXMCpc4ZmQ+41n5Ev+J+wZ2OG8a+A8G/vFE
+WQtuaCPG3sBpuOExiO2MZEtinSh9/kcTdnddtqQjWfaraAOW1u3qOcSbgQ/0Tgz
sCMdqlaUTj9GAJQiqs+oA0Fr7UagqU513wLz2a4vvWgxWSPRFmmJgNbBd4BokSCf
JfxvwS/ErWD3UppwmOZwFV1lusaliBg5LyoYCEnkpZzFJvnCqvm2KsreAFflG7pj
SiPDucW2F4xNKRXbuT7CDp0Qe1S5ah62PNSQgNVp2BZ5B20s2TP9d0j1WSs1taUw
78Om0ka9JRKtHNvb03q1wtFHItjOT1p1coQG/1+1nIeBIx4JedRJtN5B2NQ08Y5g
OCtvcs3uIMdpy8q1m8DHPOzl2ED1ZV19wrdUov8luN5ChW/GaW47M1A1aHN3fC3X
oqC9qgdSroC0gUORZOvZd0UI2aU4tvYwgwHkqzpOSba+XGi+AiRGPwQWu+tGvlXr
dP1ejP3z2gGTIU6L1EPHBzC/avU4Jom17kt3EcFcymL/JQolSpzpzgzIiQFDmwz0
uIJehiL7RzFXgEhF/CFoJL0X4HbJemrvt2gfMTVHh6K9+6hiSpzcwutzgn0TTEu3
44VA6j/6CxjKP9NkFKFUZF9zdO6Khv7U7iM3PapXUJZL4x+UkZJbC+rkcu+yBi0m
hc9s05qmSWufZOc4LOI4HD2MTYaBzWsJSU6SEj0gvDNlmLSgQYUgAMUKejoOFKm6
G1E2X523Sp5U/6Tb4VTflmG6Xxhs704ONP/tAKOavWxHZLOOFMr8VyVqE+09mPAo
YvZU7shu5nKaosLtO2K48+PimlritWYR3nvK9qbXPEhxjYXcr3dbxv5LtyfOryXR
AknwciF28/qKLRx56wP8kQemy4uHlrte8JfWAKiFNpMr3ea9STr0btKVFmHGXK7b
dMgtb/JuCQGDwBYYxejDP6WvgEJa9Ed6I5ljDumm4GC1zDZvggzj0Ka0yjhW4l29
9Ninvz/uIRhSe9bG8/q0x+9led6mZkwUwZpfeSbigTLrFkp6c+hNBtFbImAI11vA
9XaQ9RBBpZjaVwXjlf893XeQT0BHopcP5807pkJCt8WEI+BZLZ6GWoQ+FcscVbuV
ADw93/0m2AuZ4alj4g6j7NOU9IOtkNmHNXDD24rDC73Y/wJT9zIsaX1lMO+RqZ6E
CtpNOMw1ZCxtrjDmLBSY8llHfu3in+RhxryCLuw3Vi/uVCq5xdRafx1n/cmeBdai
zearbJkE6C0iDWK9q08yVDu4gtgy3Iq+C04sCp3StkbooGwLnxNkrjXLv3I3/b02
NJPML/WG8v6vEOwPzrNRPKrH7maBfv5dMG+MVa939NqNpc81iqUF7rhrCBzIGI5W
mGoDeG306zfRbDH6vctg8nk9JHNUN8iNoESTn5mt2kuJRwoslQCP32Xko+ZUeB/C
mTpLl1uaQXSP1TAA3RZlDzVoxFFCVy1FVvMtL7ldkMk/GgB5STasomYh+06lKSOG
jNQO5lq3lvUBtFNSzA5d4yEMEBUSOF5tylmXQU0ag5Z+F2bkyrn/zqw7YgGp+1Uj
eEsiPuBELOpeszapmpogYp0uhs0UQ52Urt/3YJEBePF5gocHwMcCP4kFJWaQp5eK
rlysYvqxBxuPIF1XC65ahu5jyzCgkxiQcFeH8/1WCbGZ5i/2RhqYvFyMHPCOjWDr
r3PbEEFZpIXhFYrLIL7/qWYXqbLl72Mm2HgezYMFANHdU7d2ogpa5WwytxfbQwCU
VtHk4ahnWmRRy86TAKRXlHewf6nvY450dlxNM7OFzu8bbbqJl/0jjBxtKkYj5/2T
2h/Q4w50qPe/EKPlOxOhQIUF/R1B8eogA0HyLU5gImq72IglWA6DfsjMAiPn48nV
sX7XipvnoYkVzFSMRvamflBLCugpX6uuW5e1725BWlA/A5olvoIEuOJZPh0YXup1
a29enjSj0ZUMdDOQRUCS7XrgYFQ70x4/7YWJ9iWyIgXuM+tvW1hlrBySV3rgcVH7
aP8JUG1xaPf1mziWId4Qrh620bo3N3E9XOVBvlk1iIsqjJAP3/0uGPg2Jzee2b+Q
JemvvEGwOYnAZ6NxOfe493xMpaFAumI0uE657ed7JPCc36WfV7kYlTFyuSmvzw7l
CABCgtFOgbfBC6vJwyifQJBBSLgQOKsmgtsRu2IsebChvokz4SaH/MREmMwuhMdD
mAL7uDsW136wIuc4omt2oNMC35HTNPF9Aeql29d7qIblkFr9jD2OwnrYL7j37e8j
8gRNeHReSHEsT+tlNOZ+4LVQUJB7+nixsOPKEU3upHopPQqnGKRPwDlCFsfkzrF3
145wFPM7mPfBszXPR007b9cIfP8tMNRF4vq8hKmG5nLIUFkIVo+t9pZA0mfCy4Or
8LzyK8aynJQ9b/qVfiyUdpoFmv2nf7M+3fsljfRXvhtJDh1uLAeoqYokmnmFRyTt
yiBAhN02k+KaMQlOUYXxeH+hIg5xWjt7e5Xti27t8aHmII9vEAXa6X1Sd/EHLqPb
rZ2WPAcdzuggsBEUvTSjhqMhk23PAOpBa6sDE4kYSJjk2nfCGc8xkvOXz1cYtT5H
BxNU8EE1YknoU67WK3wzD3kJfmuftUznCFjAkFDjpvMwSOcPTIGhQVR58/D4wQ7o
Fr9EfVL0zLgvYJlUOvyGJezTRMITx7intX7W0ysMgfHjZ2pQtAbpNtrk2A7rTJIJ
WRfW7gwMkPKWHomzUQJIaprFkUAuK0FBwaiV0L8gka2VDmcFrH2gbqAhBQGTzr0X
MInWl/Fgzjh/OzAx0u0OZzr2yE5jvMlWfiVrE/LZvIwv+F8HNL8tfVy48xVR3NuX
/ql7VwR7yZFgxjtpBowrCvWTsio9r8pNLJRisfause+PqsA3k1h4xnaBt8tikwKh
BNKS0iJdxe8FvHlTts39bggxrMe5tiyH4ADS5S5WRaxfvtH9EtsGlgG6ScRzy7TS
7yLU5zZ36bc2bgFRXk/pe5r8c+rhBojvAJ4cfe7mVNYNajbhQuY8jSzLlhIAYeAa
n51we8I8V0+DFF/PedL3NeGcLMFgsLv2xC5FjeIA0l+BJNdskTy/Xen6rkCqiQoH
rXU8IWyXnOLuLGAUvKLLlpX8QjvroVYfUhrrjhrzBi6m9A4hIyRQbb38ebj4Coji
MaMTqalen0rEerDXoQzNWRMYRRtCDFvEwrZSTMgTmVjPRJyF1Vii9K+Z4D+DExbP
LdW6wgf5KoterL1zHdNduxQZ2h9rcuEUmJaRfrxAqpvYJIvMQt2zfr8sha5W2S8q
GL4gCI/HAauGhQ9nwUI6r+Veg1fktnvpBa7cWKZEQqc2rVZNq1KrYWnX246nUidW
QH/4xBw6xhSaGlwDrevCzmjPR2Ba1ZDzAmxRIVNOTzeXsi6jxG6ZmSTE9xOOsmxR
w98tMXQ+6kEKhRntsDsOZoIycvmaermpX125YwdTjTcnaPbupOT9389U9Vi9D6bf
zgJu5QOc12P5Q1d6BmGp+8Mu8qGEG9F5600ZuFgjUq8MqBI/S/gNxi+S+NFQ6qy7
QwAyYqt7G883PnO7wMNf5fAo83EVKcDL91DpK3MUM1R2HRdQOQD3F66atLRv5nvG
37Xo5VWQy7mTSz5TXKLB6OH2bgPnLwUW4Bnm1NezzDlHYuTU0Z6IaI68yOcDAN+m
UmuAX2oMafSOfw3tVdzLzn9GA3cvHLk5npiUbd+BZCdk9F8EBlbBde8Sre4LVYGA
LDa3vUhAx6mxP582fthkbFdXsD6h5nzvH6UC7p0PT+3vVPPX3Xkh68g7VR8y+wk0
Bc51AGdpuVpJS8Psyg1pR/3jedXS8YIJ5OkoC628WWH6faV5yimQrNBZPZdszcgA
Xs7WOqhsHM/kynhk5Xl680H4SNKS8mcmjoNdZ9lBSGp/2u2QOT67+NdrNODC/KBZ
alv8SPRUUflebyaHLcRnzs+Kai0U7u4oAQNy71HDnKpHLqcAyAEMvrfStIiv4//I
zZBIoI+iiLlcY+96PxC4YniBhvLV2R5gGjWga5nZj/kiLWlskiQ3MYO+nVaizdX5
2h5+2F4OJ1cPQfFykgC/kjKOfOBfFgmZRXMS/snImdFR2we2nup4gHbEDaViTlhe
JBdbptN7zOcCNNCZIGBsJbhOXOx8yWJ0GIapGqJ0q95a+2AsAQjXzIjJiOVxDgW0
xYR58w2rL9AjmX0Jj4qLYLHwfk/HpMGEEjIMjqRsZJnFFyOsLXXw3XFNzXbYV3GF
JcyHUlwr/5fxpM/7qd1EPGmDIQHiZjCvMkg83TzSYigQNJYw7jJiMuu7Gn/oDMp7
aVmwjkW/QTNu2fiCcw7YrFLKEYbv339rebpPgVtLhmsh1hezMJVC3HG8BU4YkrTu
3TqcCXqvcjLAtXKkFlV7qv0IzKx4gAxErsgPLJoHBvp0/sLDKhMzdS8eJn4mPmpm
aZ5zQVnUSXz4lWHlX+jYx+nx3It2LB+8vYP/KowWSrtcLYgaXYu4zAm+lqitQHCw
NTJ7964DOBdNjD0sTqeLxZ3bTiUe5/zsSUWbPw9kniGh+bJoJ4+AcPuoaMKorvss
UCFsuaDatAKUAcxuph6xuz9ybhVAXo3laQugcIaywv/ki/tabpJeZA4Jkz6lCqSy
dVCkPQhVM6EolMH/C2AsWR18xNnt4a1BBzKbw+KeUflPaweX37AbOw1OzymFb1Uz
z3wVULdHxGVwFHsxstCmJGHgt41cM/o1VjkSg0NzWdyWh5ojA1hBmt6hMD+wYewc
LB5EO2//bjNr7PKrZxF2FuOd429mfkfUqzfCt0PstOa/ttwAFtmiWdOWfHarrlUC
6B6v5uJmpmYuxOJoJHSlmbrX9XwPhJGrMjUFOzRjtPqTXupLV5csmg8NjGw1brBd
x4w2f+k41W2DiNrz+f/3jqkOndqcCjWv+/f1kvvHgij4FpxQZlR2NYKItEimZLrD
oVXPHhUFIvbD/G/5S6zJyk9qJjJ7t9z8R7c3qIzHFqAsvL9HIB+cgDGwVDhEzUPc
WiEzN5Ugnso+cP45Giw1hApHK7PfAL8gT51Xwh0fDbRWzcIvzWfoWwjIi6/96CrT
GYG2HU98UKYBry53ZTxmVVaOvfUFbWp/cz3msfc0aMMnmQ18eHzcpwEVIPnXeDd5
jD/ar1nzrZs1VYUrglwyHAgdaQLTYPmre1KLQoKPTy7yiIjicm7pz0tHswoe1rGT
eQbKk+39zVtytYCVOz3hKvJPKUZbpPUyokvxDA1oUk3mtP+F0RANwUWBeo11VHsp
+kbNW0DGGTTs9RSz1W+RNygBNKLG7UYg72L3IyBNOZJJse1nutH0W0EJTV0uVz4r
OHwR4VPPezUNoFmbC9x24DjImVO/EMTalv1GVgodd21C83VOXg6NhbIdPwVfrscg
j3pVl+xbLiHv1V/lbn81NO5FmZZOJGWRz6RCiQpaENfUhGgvVq9Um6vIG1Uib7zp
r7ygUPP4wCc2pB8M3pbOlgYiwmu9DGjaiNZCKdAbx939T9oYA2JrNM/JAPVnl74G
mumJsv8pjAg2RcCUnWSAp8SVnH2NJPtctPg1i+Df/nYKvvCG7RUtwFLhbG22EQRH
kRCb+wnDQtznEACsmKClhNT3XtyI9q2v/+k2vwqyfgs7UukDaBzcsyOeEjdaGRnN
yz7YLqkY9Pnl6ch150xwmIFdIQOKRnEd8HxiRu1CO5v0iSx2MV6XBhTBGNvwoyIa
kc74lJbwjOywY3DP/rbaNewJ2YEzKTCnAfMdRTu3pE1b3RcjSOOUG+zrpD8JzAX1
VguGIGblVU/u3dmGr63sQUnb7UlYe6oRXeE/VQwfpygbJpe4BuRmk/tUUYkf40TV
SmE1IYxcnIpRBwk4GJDNHbZXLtrxA3+p96F69E6YX3kmIaxlO/IK3MA2AQ04NTzj
l0SCUyYyDjzNhGcdobHO3Z51yidsv6tv5yohWaKqqKfjAMk/SlnLvYNPdYnzZcBd
8EfZFpU0Oyt782zOvgIZrUZBr6F2iswke0mpuXSPOun/TevB8CD8K/Hzs9wZFasv
HBBvyznu0o71DUjxl0mQl6Ev5y5KD8mg2p6CMYx4J43fX8XYOmHdhcR3vWLw3D/J
QGr/fDZeB0nEHv4gdNEBZD1O6UkVe0XwD0GfPfzau8rUT540KzHibmFEWpQuNwBK
42qDaAP58v6MRJww2YEiMnR08GzcmCaiX9WkrL4/6oQeM1TZl6TwXWuRCB19RMFT
r4tUj5DARSQtAwHA3HzydhjZWMEAcUD0a38ZSAk5PNxlESSMwjDvMTigafZHontR
nsFev7d+6kjMfRaHH709mJzkaxrRJzUMWzD83QEurqov4sNklsWumkcUWxhDsu/P
eMmnvJYc0m4drPC/U/IfHMpWzekuh0OAjYO00rH2bBRR3ItQDJsTUG3kZOOrPnJp
0YrxxOkwfEthtIbuUI+ZJS3fvc0XyIsV2riqCWREWeLXRLorfUkIMZtR+YJ9Jch7
cclDYGVg3YYXQ3gcBmuiygRc9sdZy/0vSXQjfTlpfynylbnwBkwu3Q7jJgqHpDpP
HJbvBAX2qTg8D2aU1fEp2nl2xUkTDjEaMU9POK6XLHvWA/DkGFTCgiixJ5bC4EOF
tLuObzgx2KhbG3um8u8FRToRBu1xWe8s9hnP0awM4MM/r+TDW4SseDQEWQaI3t5n
qkEf+Sj/QiTfn48f5oIOrzaSIkwoTCDCvE7IWgwpwhKxgzXieGGMTHwEiCYyC1Wb
wNI+8bGgQznrO3LbI7YWjlxAsnmIUjagwmL32+E908CKwWkpjMV0uNJTAgCKZ5Q2
ICGkTIhq2dLg/OFpUhNdWHw4Cv7gKQMw2NSiVBOhvonfF7V4qBeA1zmThSlC99XJ
a0SevIQjQgaqw8ULrTKbmATwfjkzlUyE8WFlz0WpayOGUlmHxyQSBkjx9iVKQtk5
gU7EQlieIHfmxmUQCPJ1GIf73CvfKuqis9UFgiKOflfVfmtgCdFNFJ3nBL3AVrq5
nmPBW12b+drtRtkWIdomR5lWhHdON1p+DkcTutuyDc9KXeu6wJnaI/bjoIbQMGOI
bnxeL6a9jfl28Fsd6Ckzq2/YpoVY8gIXigdmxCug0422gb0igXxfwpVnvW52+ljw
gKpcVhBFcr2r+uJ4ukcB2u9/3ejysxDl7GpvgQnOP69Nr3l0wLB1wMhE+NCpEcxb
ealslugecM/aEyjRfGH14X8qZz83+1+KCpoupSS2bjDcy2MfzFjcqMrsHC2gM8Pz
snnhk7QHzcrm4hQsZXqIJ+9Q8Of7dTAUz2y2Z5KTyn4+H6c4okfJcICYTuKq1bKr
TNwVQazmMb0WgGVGpGy1TFaTUIB2RZ40DYx+sgwccfwUFyBTlhfYu33WgPgRrdIQ
8bE4cd0NWi0MIxU8EgG4fLimCY5HqiMY9WeJeuveIL/eoFpw6l0M/2I9z5pzsNlZ
NXYcjkME2ZLNTOdt/HOeHiPbpPZ5NOwj5Cray8uc9Is03xS88kjvfBK0iaO6LjT4
2nI6QBQGv5fVqT3VokgaFA8btRXKSQP+PhMoSfBHVQjPCrbOnSBlx0i/AKTol0Xc
tO3YKZc9agudMS9TXnpsPCse7g2aM0dqX+gWyoUAeJ1Ec8jFUsPrp1cQM9AQxY6X
W6/TdIAUmjV940d3vElqjVmPnSsMF9RE940WFJFY/OfdgfIwle9nkAVIXziQc37V
v8MbKbbHsvGrE5xhlu0CiwdmMSdJGNiNB17G7xM1nX1wcW78GKCtF/Ycn1pVLiVN
s90J7rtg96SJd7gg9kedd79zAPeAY/mtL02PkqyabF0u8iNhP2y7dcsm+Ytlf4uY
CcQ1t4Yieg2RKG2KF0XQogsjbZvYy6g+Uv3kUrrIQfWD/UxaMagWZ72K0QtnVBD2
rQaU/0VbVhqfAE4eFasGhhl0pYlEj1ADuyhT8uK00f8mNsQyiqPeB62tSL7mZmLL
+o2rczzBIUnEZ0TyRTN9LuzuYI/EfvNJupvXTWb9IUnDFk+VVqLBd1SHTg9wg4jv
qqysGHfxUGlaRSr+li9/q7YtjJxwTIeT9L3l8giN/KDSyHGzmc5gI/ou3YMkV9pa
jTmlo0DAMsIdpQuFhJm9CMRhsGfLykpZODzAdEHdGlArjJ21iAf36aQzscJeVmxQ
dvSwuxNruIMcLPKuehBRYO4tuZGhWRachU8PemA2We1Tfgkb/x8XjKdr9ZNIS8W5
9n0dDH0hI1x4zQINbBUJyQuajx3yWEn1SFZOwA3bKMSrZqJcWrjbzBo1L4P/qCzB
W+LY/qYP+AzszLntb1JpOYo/2q8qnRwCekiw8h9Wb+2TpbWJi1fXaucGjAOGPxdB
/rN0thRp/6Foh5513DADfQ2UXnPjZU1trPNce+l/sRX89/eV8oBtlb54i5MQpyR5
I2dW9XYmB+fBlDySp9TWzs4ZxJRWTMKRNSZn3mtI1lTL2SOIOLESzCGzbYUw6YTX
/k4446z49zWavgKArVSYpfsN+TFmBqUh0J1wykh32hGYKIGR9yojHfXaa6EPYEQk
X69voGsApu7TI4ez5w5l6+LdD3aDuDX0+MImRXa0/Rg7slQNAQOCDE1UdqZX5+vN
bm/ueaVvWNzDAdE5eFsTarq2rhMsUwe1GsFJHqPn0ZkQxgmScv4eJwG3iS+bdZb4
x0K1OPVpDMAt7tXgYq9NHXCLk9zo6SDxfm5uqHc7Jro/Gfepe7e4NokX0S4VTo7+
QOMSgY4uBX5xSxvhrNAxNTcz4gAaiNJOY/xHMckiBKY3xMPF/GaDpVeZIkhfO8OS
CLIADBGo4w5QcbQOVMqXvn8TWqqlaB2Z4+rmqvdp5lHhIrqzBR6UjMg6ePtCS1j2
/EDzQq5P1yVoJkSlO/mBhBI3E7Mx4inGNSIL68YbjWQ0QA3UYKOO/wFTyQQxEVd8
caH6iD44mrgXxGL74v+hrj4RTiKJByu2k0mTILArh6b9PzBc25Po8wZG/8Btr3+X
AaSUaVTQOGP5op4olUKXm4x/FvAQJXq+9vvwkjoHB45y5RuDWA3fjWU48gaoHRwv
x36eRKYyG0H+AZgZEb2EHu6tlp63mAGOQGz1ClZoz5R+GIrrcF36jyb7bMcEv1kd
4a1mTg56jPBrprUc3ItL+Kkdhu6EEKugwis5ojtHzrlLIJVaRz7XBOj++g+HP6WZ
pnI03bcVbZJutk6IeNVoqsVWvLA5aD/5Ft4NPf9tqFO4nU50IZRap/KnU4XRwWvn
1kVOUdHziN7wmmkV7eKY0s6cUbABsmzs2hBR36vzjs9g0ll4fhCCVCyoQdiMUmAG
rBPnk9d2DfAA40k1P0CWG7duE9oQv3ivfPiXGgC25wrPLvMigpNh+70YuaNh6t9X
8N7HelaAlh+q+Ygyp303aScudMpVM9eb9xk7eppSqsJ2VXBW40JsxeHDbVtR8PEJ
TZBw5PeGzAiQ4z19hOYc8r5hDTQoGT1YM22nkPoD8MlVxap8we/A1JkxaA8sIXmo
T8K5P4orm5Ik2SEEmjOEvwQY6rnqli41IQ3nosfmjIPVvZuUpazaim+hR5++s6Sw
3PP845hnJSycAtKGldDKI7oYDaILvHcWTNIp3rKfe0xWxcLgq4d+YIe431sz+u+U
wOJtQhRepxYeZ2O2eiTnfGIUL4ernl3vq4kV2+Gca2lid3Qg/LZJsrh5u0r5q1AK
WIfOY6OYnoAVbbPDe7+wAfM5XNCVg6D+Sht2Z2iFr1NcLT+oaaQ7A98eBYgWPRo4
dxUKkLx4TO/hvQZi/shu6o3wrJ+rMC+i0hOqdpcGMey4+ljKsYXJYFaJQcxGbXvf
haWyk9fYEw6r1hEEPUq4eh8KuG/dInIJN09kWm8EC/4ivkqz5d9Gflc58N6PlWFD
YLxIzZQl4lDcsbHBuLeaq0/ep1kq9skIkcyTfWcN/R0ARfbCkx9CMCbCQttbhU/U
akdifq4kSHJY99ijHmjo9/lVEMgoqIoZJXDMKOKIVv0FCM9g0qoUyymipYpltH1V
AKUXestvJO3HebBwLXLm2UIPxC2ye6kcu+y5pqwKX1mt9i3GKdS2CwPhJLLvRFsh
s2HSr2Vl12slo+0NoGXzFCvJUDhmWqoND8eRGwRi56Ucapnn7uI0NquWh8DPC9pe
rTA3ZOJQ4DVsVcKFIOQIei4nqdaYoMgVv8OkaWf3uiaz2ucykwAv2CnXiQJp0Rj1
CkQYqymSXMybqXzJzeOuO1H2cAIhuL9TpIq5aAk/4+jQ/MtWywuYrHBQSrwYKas0
BrkY22xABqoKhigibZ48PBs50uqnfMeEPPYGgX+TWTalXPs5fxRkhwEhoKQDjbLT
q9juaWa1CXYJxpQc3623vC9NTBqFT+FQz4IQdtrmoBRyzMYbuGWrUFkYED+yHUfx
bRZRacr6+pDDVP5bSvf90pSSoAHab8zueT/M48pygM6nIVfv+ibzKSN8RkFl20aW
c0QAE7Kjhy5HYDSqmXafH481wuNIXNxrYcnWgBhkoGluYFKWOeDyhAlOf1cxYJKS
V3juD54yOxig49zgkCtE+HAdQxVhGGYpsjPYw7zsH1kHn0Sdiv5BFwAe1Ehkinha
t2XIDDJ6C0zwL2bPD+zGyqlB9Ebelzmyjdtty0L0MEP/YvyauaQEwqElhEEJUSPg
4JH/5Jozvl0HubDxxXZALOm5DpSUrEgkLQf7l76OaIbm1hZYBLVM8xJIFJzy1s50
LS76EJhtk5UXdv3APreJJHCaRqTMk61hAtmOhYvJ0LlYyALIU3r1cGgiA5XjxPHd
f56RCUjKRdGZq+Ll0dYEf4rADR/6tVvFB9rzXSjVryBfk5a3wbvre57oM/XCE1Tc
k6jzYq4o28h2dpzSg86KQ1qY6voE1UCvEBgmDjEZFO2dYYlpVNKKPDh/Pf7o+KNJ
gcQvEfgcKyAbi0XnCIW3/t5aJHHNpMmBSYXA+WPn3tdGMAjbzC6TJ4cn5to3mPM4
JhjjX05HSVvIsdhqRFhQ9+YRHKbj9SJDSJuEYu27HqqiZmObrVuHGoCW/fgKWPCa
NI/PgppQCcaMDIOMVyTiz9wkgDQm5AQ5ytx8eepAKxejmZzF3uQuUQXJ77yqlZ+C
FTfNKDlQAJ41rE3smCMKwdr4ihe+Vvrx9B4mqTIOCYovUdJfD0Cea6Hg0W6cvt6H
lQJXEkHMBZMpXTrc+/+9r4LP77ILRTTAwg735dd4g7c/kkhQLeqd4vQ6eWPUruoL
vqf6t+3T4Adev+b+gGKBYZhqPhOfCylgaohIj/jxn6M0f2ybrDQsjAZPIlou6v/U
5I06MWDXNwLpw2S60LwaFBURwqVStK46cA0A6/+ARs7jbvxIQFJTiBBiv0M7RkcS
Qcu1sTQFq7LU9mbEi1z1qHlm2t7ADW2vfV9f5KSqftwELBKb1qO1nykMj2a/7DPF
LLv0iasRIg7wJNxrFWi9vzNCKtZUrGQgVtUffwR4hWl7ffBJVEJ6uh/ahEMagJr9
6ui2mlYHcw0HYTA25GFr/nTv5/z/BL+zmNQ7qGMXgRu/E91eEQpXqsI2GeZg/uvT
dDLxlfJH8p+MtLFHMLcmARUtR2AChlmLxcIXvIMyikINLBZpAXG6TqBKwBGJ6zS+
UVwUzhH9IETgdD0nJosxZM8PYnWnaVgFucmlGSV2gMtA5h4F+6dH0DmWkpEzkAcO
iFAekgwJuuQMntJ0KcMNXardenZ4M3ezbbEv6u+saFTgP0y9BOvjoeCOvQMnqtD9
Bi8XygcMPhN4ny+QTSYlqP/xdrVONioowmqb1t/lrvHNphBoOoZFEY1dQDkP5JYP
l1HTD1VA3V1HlLZ5E6RwMT62lVAV8A9/9jfLuXyhyFOm4qSipwgulexMeArKRVug
eUIwl/5vYpq9X3lm5kzgCC2y8f4Dh3dctCjDOzCZIJcUXpZKDF91dPDBrqvTMZYn
PyLBjqN8P2ZJMAnfbg1+gfCJgPDalVGXy48ipSf718qEVS8mcDMl7UidRhfgtGTy
J9L18rK22yR6EbCkq/JrhimI2Ca+qL+onSC45I9qiC7rejE4oUvNDR5IkVRX4oyx
nwHvCf+HheUeaNHNGV+sTZ02tirsanxudj+AvEDUgsBj7A5cyB5hhxsdrvQk/UPf
rpn98C9hSP60a2kscs9LgRE5F9Q++7djTBMiKgfqKvHd2eT9hgH68BAJccb/fzXv
a8T684Bfkg5bzquxOW+Mvigsroks1TAd/wkEnoA+i8IW5/MwUpD3PXU/rooeTT7S
hfLptNIvxxvP6iGVBFsR1j+CJ7X3JZSYTAT1RWjfk9bZgFmYx6MjTcGLCNuq45Ol
FV3E+5p+iD/n3ZCFj9Cm96G9vXfDVe7uEvDeunpm08xmZTrPPFfu8wZhUcN3lFHb
fi+5ohg4Sr1ZiCycLnNBeuCBYiYUoZKTEWXtYOKWQ38eDgKt9tWShhx16Cb65W5p
GOiPYwRaIhG8r6r4Xpd04aAH7+9RRJMcB/VlR2lOqWFBUGOyCJQ7QDo+vz/uSdkf
UzvFj2OlXWW/YKjgoHGn7Is9v6YASHTzUH7CI6eCbhedIIecvxVv1Yh7OvPRO2Cb
8cn6aNizdskAii9Nm4Aho+ALx7mqH4it5N7N1ZA1Jl3rSFKY0fRcpCBQrvzDmK/R
p02qaBiFeMIcWpBOESchi9xGpytZQ3DedLLCyopYP3PM6Fe8MzieS7+sDNb9LSex
5aEqluRtKcxHhoU2ZfBJ6wiLFICCdaEynrhHesm/GaUPDP5yVe6OxHgG13tDl08y
x2BkljcfiqVT/b+UWhOKP2H6H3g4c8Jo0JtIizC8nr/3H0Szrk1dsbPuayeSz/PL
Nmw9Lje8OyKvxvL2Qfk6mfIv+gnE0qJfgrJ30h0hf1YdDSRytoD+AUuLzsyJdouk
7f4DJrckgApOrjqYAmquxXYTLWFv4IiOwygxwBNfsIXp7cmmFTWv/awk37l6zV2M
9j2pLJiOifYgl7cMgYhkieuCb6T0q4/+g7Y1JYPQZROfUR3SMLy2jcHqkLjT/FVb
Wf3mACR9tZmBN8V8/FrAdiI5KKbM6mi52PDkpR4tSamYlW7ss4JMrtdEwTJXoF32
z0kmmX8VTg0jpVCN0X72Z6WYSpKX8oTCGQb9blMZfkCjgMayokyjsat47XAN6ZNu
jsO9uKrlkIHFcWf0nX2ERnmbuGCjL8NvYboEMZ5P3l7hLjCagIKLBCoA9f2hd9SW
XqPZO59T6D4D6EpGF5tQAhweNoptYk6n5EyNnujZxnvB4IiN3EeQsYUXAc1af/38
UqnSXg2/5sLub+NTHd9znRPz7qqBEiBmfi79Ti3BMACF0sCgg9gW8YsgYuL/JuGS
BdSKKYMh8ObnUkzz/Z+EH9WDXPma2eHoXU8NYuE5qtfNZtJxeJ5dLevXWEQ2UDd5
q82wX74+MT98HAm642SwllYMkmq7tv1UpfzNVb7eSIvIgBABIgDAst+n/2i2vykg
TvPCQ1FMm2mwaqQjAQcXhBhASCgyNKVfq9KHpzB/BHNLR8hBWfRoMZ6DnJpvfE9j
ss5vz2O4069t7ml/v2sVYIRWdAtysgleNL540xntCu+BfSp45lJyHr6rqeuXwQCe
Fdvh05GgQ1FFT58E7VYjM9YDofZmpHUHfAVz7pgnRAdmp6MJpjZ8+L0jovMBoYxq
n3yotUclnuBzz82Mu/YOMo86x78ymaGfJ87DG+kowR+K35M4zvDHC0tGeJ4mBSn3
UyAb2Omv63vZWNESIsLNrjkQ3ABVGJS9ZMbFY6VuL4veEgHYvcmq+0jdZBElzqWY
pVosr99tpxvW7hYA+R31dxPQLM8afUfjqk5u+vPlHgjVxRNsYCEL1KWwUIMzacNF
ftDcL3D8iWwwj/RaXdzhlYW5BzAsYmNT+ni2/87A+msX/I/+styQGXZ2dpvMwwn1
WfXbIw1HC1Tv1hoL8LgofkdJcXKVnrDiHNwvmUlT/XYPRORwpHXaTuewxkJFjmAg
jC6wyXNjD4Y4JJ6NseANXEeNCmitxCh55tyuUtCTZ3KqaoWeg0aL6eGx25DJTNhr
a5ouir+gFUuMJKaEu0qL2vIRE+TLixwIvBA76WHQ7ZD/IFWVflb5yGk9PohRFJeV
E+PuQL22UqmLwD0FaC8781uVWGJdHAAmfx+VjR9d82yipz5yIrD3aeg7L/9EhS6r
ne+vTb0HLX86/Z8CNNcI8fhFzjq6TUauc5qqWGpDwWNnZXS2OF3YA4ZvOdBU/6bp
Bi+OjC3KeNmHaYzbcX3XWsaz+wWqwEzl3iYNT+Omuyfj/XHHInnybRMSRN5nZXAi
r1eG/D1PMzFaKmNkwcx+A0tqG9ndqLqJNYOj45HfNdPnnQJ9Je4+icoGIg2c1VcO
FofpAac1TlfE7lNgzhpGZp1Rk0Ma1SsSHo6hlbToFqm/lGA/tvIU3xsj+VILH+14
TZib90GWvs1mZuv9k9IlxUmsfnkt4mhBts0fow7Ut3qoertaeuhXUK0TuQ2q2Ttd
KQqvF3wUIjfFhidCkCzx+NJvIf4eNvoQaeqMVo5mwsFnEc2z5+/lYapnv4js7cKr
J8bm4LUjZMUi+CibB7uO/jt4+z5K4QW3oFizsv6iRD1M39Nhq8u/QFnzyoNuD+5U
6xALGK+llX1FdZEUl6XMN/XEQk7EEAhagm18xWJ/vIPXlrnVTAB5mcuwScwYXHeC
jzLRNeqBZSo+FmoYI0dSnKurTzQtKnI9fbU6WbGDBniKMeXKOzUFd5PHU1orlp6o
6A1c+L20PgqxjzYla05JzhGIIPiY7FF8++imwWvbQf/QMCVTzJ5QgT/dD9QccBZX
8hxBzXAVoA7BmQ6Qv/lx+ebNgoBYwm+BsHNaUmdMSAb/yOlczJXjBOwDUZDAlwC3
6NqRXnY8o/c/IRE2sSgOxo78hnbCD0h/k4OzwFNlApVcpmmsY3NxBX0jQ0we7tLO
VkkJUkqrbjU2V2nuycW6/Ga6jtIXJuB1BGMAeGG6ARVuTTzZIFhjEyaKxO4t7MNJ
7WM14HUWg1sNMZiIgsfKoTvIubipiSvtfM4eI9v0+OjS/Q9RG/YargW+z8qaa2A3
Yxzlbp8RK2YxaBu5Za9+846s0coXUqTT/+6sCloV8tptKsqJGata8kWhXUox39DM
E3dcWjmY4EM7sxRrqVJVo7OBQMjtUVYnx2LJeA6jZDrzF/HW5wCav1eN7gs4Bjf7
gy8SCrSvvd+2Z9yU2Lvz/+BlYdcUdKF0mdR8+vMV2nVK+6DO7knl5Qem20xWf6OU
z977WO4Ex+YbqAu/HA0FmqDnyqikfb6hzvOAubz54eSojHt0/eL3ol1m6gA9Zk12
aMRPIRxv8ofOY/z28oVtlWJ/ZDatF4ogICqrXIPjsVOXzBvxfJY3uVg1Bg57+Fa2
LjcMytPyXRo45+aUHJF4+Zib6qlFjBJ++pSDh7aryb2MaP7wvmFvmXf5NqozxbSK
+Edpn4sHg80ZalGOJ/sZDVP0yjp100pAK4ZPKv1cXasQGEz6vrSjQ3ofjTkAhTOP
TGsRvnUqRR2cZpnZfDuLVfxp88C1Y6R0hACuwsmpNVHH+D+dbVVFigclUD5VDDkz
gwDge1TNZGOw+ews0SF1AzqsVkze6IcoGp8K+cKz9dl6VbjY+9T3LmFfWmxbnakb
qwzPq2nc44PlhjfIr1j7byGyyQiKUqKnOjw6bCJorPXFYmxR8pb/ra7NUxU5y+9L
KnfGORLn+yN2IbpGq7T4ZWtjPRF6ILi43/rxa7YTdxSQzlZvlEM8eJYUoQV7CDwF
ugcKyu3pODIFjAvQTr4zvxEZTpoASyKWQHv1wNdFamBajfeVx54c7HXZ5Jyb1wde
qNM0Evl5ZmaQhFMzIMm8xnEssGxGqmywauTgzxfzT8jKHXRL/HfkYei58yrVN71y
QPTBQsRaHXCNdSe+nPXSYcfODF0w7PSKzCpG7hOzQd43P+3rkvhuGHnGFkU8zi67
U/r4rRyRRGdGlXbZ791kCH/XG+j3Zd5V2ARwovMnwG/Io5AheikLPNswiYSYzALP
pTox8IGA6ab9Q++hSbJkRbBgZUlRYUKmACcFElMvhhCEXxHVkQzXo04X6SVc1Hn1
VcNsTnXe4FGG9ZqVMzeOPE6Gigh5SyUdW7EUTby0J0xbL6SnJIw/gj6f6mIL1Djb
BPl9TUeISTkY4fQU9JzGlNnlztj5SrxpmMmbuxev3Q9A7dH9g9KBPCxF1MQzDX5Z
MEtiK30hUEdcd65lCUXjXso4NitOxyxXFI3kaaxpeKfonhbCTspUiJOz5DEItyW1
I7mduSqTd1kFojWdqYmrqS80bkfo7Gop6i2CAjpIzAvK/9v+5FxqwuC/BWEmjBCz
ZljFuRTAZIKhVMxgb69be+Ri+RwIcNC+D3wym+JVI+UGGgyd/glpTFfmxEEqKCA4
0bedOrzmKX06t8JqTiTkl9FsVl1MWTsjBEDw+J53oVvLfqYk7/dc7DoKRrvXNoSK
xg8pcBbtS9OxkUb+3/3AN8vgIR4kv0Kju0dgYPipif15hDk7rPiseBEe9salOlod
Wr2i0jWfkjzzFgdHzTxnzWZcMdGsqao0iDpkIsq2InQH6GdQ4ErepUwFNBkLLBAG
JlFg4Sntb9SNv+0X2PeUFfErxV8Wom+bk1LirLTzETz0Xk9Q011/pbwk4ACYg2b7
R7m9RJP2lvcaeQvEmpX46RobG7dTOFL4Rb95NSVPz71meyjISMCDuIkc1lsHENKo
awHG1yFEvSgCgwfoKwXI1dzOXPgwK37/frXkxolVTFqhimypLrKwnOL9QQdTsQvp
mW+oSvKc5QXpE8TePkLYbVtE2mHd4KGfJUM1/lvABJ1mJDqxoavEi9QmgJAsV6so
4W9CuJky2FAHdPvg2eJCQLjv1YVpvQCmGiyMmNxmST9Dv+buG/Igoctwm8a4puO3
IehHr6smwDCtDFDTfwxuO+/u/cMOioeEKIW2LY4zdUBU5sk53mEybgGP8n9dlqcV
nf+lu3JHxarkwWa23FPL0RlD/JQ72MQmXiOswm5rW5ypdybWd1cPx348HwrvFKCC
lwluAGX/BvzuR1sTODwFQnI8Q5ctplfFFB3Dzcj7AkvOfa744/qIn1+YWjEZf20J
YHrgPrtJwhYKPWTRKUBK+0BsIJtk7rnXMfhN+tPXadjQ3jMISl60r3H7dIo+QWig
ZdZx4cam2oLWWZ9WCTxatPacXiplokHklahotyFdE7oe6kEOQW/nBYTai7zkUHzK
DZ6IpbQPyQ/hnGdk5u0TXzaGJz7kujPxUlKbmG82c9tS84GQRyfI64uVARWqeqYJ
wYOZWesspeBnZqnMtmmNTheRCA7SGcQ2gMjT5w500CSV7/VM9h0AVKvW3qselCFI
EHYxqHMeM5pnD/l8JdWeueIQ3PYzw5QkBWAsEzi33wwyOPiDoK99KhQ4I4ncauBf
UBBQBtGhtXpTcdPXMsRYXjP/o/QLRCCKZk8ZLQg7prpX5Ypd5MXkdJ/9DFnEWwhy
lRrYNZgCKAlP/dCEyQ0PCAawodXAfcD09RSh0Cvmr4kpL5Q9aMOARY/YNmjIWy0c
eRMXG86Ynqx8XDk4jUH9MYDANU7UGFkyaKxpzyeIPi1uYwGellFXcf+A3SrvaREY
jVSJ3EtviX7/UhbwPbF9NsvQa/9TOWq70/SgxyaEpEE90a5T4fZU2ETIOug8QhjB
3YjrGX58e5HI+gHFIFmelHrFk0MDqL5T+p9jS7zVsOEwBKhBF1/nNmWSPPa2QBvx
628wIp+Q79YRXYbxz6qVhCLtu/SRHL+u2N7WRkMBCo2unBI32pto/22FQd80N8bQ
MbX5gQ/8q+WPUKyFCXIXdGnRMcdV73/4lPf4Of6ZXV5WhjojvyZ+cFD2KqJ072vG
x90hd9eS1QkVMBh9VO0XIiToVNYx6h5IjUusIm4qUK+DtTwj+aKBkkSkDr/kan7E
0vqAAkTLqm8mmJjPMt+6PqtqaPOJDWnUhZff+4cWnDXrh0Mpp3uY7/he4BtG0Ocu
X6zQff2TT9HTvcijZwFBv+lQfOonrch4GPsxPk7Swfgeugf0OVo5nG6BnT5nIZ6h
1bI1WjKFhoDytJLAWnUjC5jBN/a56uDG18H7NNMGJ6UBNP6Trx4WVwglhYeWSXxP
PecHBOk+JJiMkkAihujQC9FGtR7xzzthKuR078DvdT4sgJeZpYiJM60bWWOfMdqc
aj0VFZxJh8za2wxo4KG3UzD/5at9n+6c02lzg58R5bIVVbe0Box/2e7Tf1VT1WTk
GcrKyCzjmbKnvMsx7/OIDkKbZjxRkx6L5HGkhEZlWbDPtfDwWSvLyuRr+9Wrz+1y
5BhAyRyuCAx+w9mzjNomCYEUMvfqD+pnKnZ/ss9oYJVUxy6RoLZehyVTOPNnZ3lC
+W1Wugg5RIleMIWX4FrcupDM9lfXb5YbicDY6q1r+jeL/rMImd21Guw5QvgRsonJ
sBSN56R6qvixaQ/kuhShPXsCA8XW6MVT+z42erRqwYpUtvWuCmPiKN3w67yZzNXl
r2T5YKSevzuYXlkV3rhzho4jIV+aVrMnrEf8+dQ30YYg4Ik41h9DkyvLzO+hkrD7
hwxkjlALZNJr7cLmPu3LAlxesd+897moM24EMEkjt47iWwVP8nEgiqwhlfIIxEdQ
l0wQnp2e5p3iQMDuu3n/8VOTLyP+G13stcaFmrnSPyboonShzm6lI6rVs+2HIM6/
4k9sN4OJxgKeAzRodhMoV9TcjGR89WMl1noBfVTOjTzs/dhOeq7Ts0/1KdoHS9DO
SON+ONLCDuOxYsdcr8mBV59cdwgx0dGNs8d/2zM/aD5SHsvLkopxiy7Kf6+lll+P
Eu9naVMAHkILpF8lN83qA7ckEMtJxffb3cbKvL9Nn2XQ3RTvIbNmntNwWKF/qjUM
wuLyu94mLMzolM12jL1YTT3a9CXMqd5lSuaI3KSlMInubMljK+2ga4qpKYlHatmn
1hK4UupT6CflWf3CwpcjRkq/mAABYEyH9DNCGB5YJpjeOblYFUSgbCBZyILuAL9C
pQvfitz7HpdwHtC1oJZmmS2nAJOCVaz07Gtiv+jArA2Cza2SS3v0bqNwyJjENK+V
mTUpJgENHFyo/ocaO+Tbsts0XZYW30IrAXSYDVwVbQ+k5zXwxRBc2r/ZUEQCVy25
rsghQ/yEToeFpp/qfho+GF6fuSYdAXmfwklM+3NCuOCvyJ8Go3Q+OhFF0P9PtbJH
hmndIllWi0IySWnIS8Q3WSK206fnq9I7NlOOBsmOZzmqMRKfvz1jCyHptU9Na8dW
XNqRctvvOj5ZrWZA+PJARZpqLl6LGl5ZGcTgmMGJyFw7aLqU3mRnM1Mmu9DuXFkZ
gqSllonEX8JQNlri4s/k0tgbynRdGGKny73rloTeEtvsmZG6dnkM+XHmEn6qUtAs
PBF4BpNSYVouoyvjWyA4bLdrQcNbJZHYvQpna80dbhCrXtL/dEese8Qy3md/au5n
XHkh1OX/9fyY1yE2LfysuqsqmuTju6PZrp59dw1kp+RSyIMFCCuor8r2cHV4V2WY
nm11RiquD1cAnwjBOH2m66eP96Mq8bckMjbD+KWo+UDLq2twJR+PYqQw/Rf1iGDS
5zUJoVl03QyAl+ngboAsM2f9pMhd3X9NWjspLD2m0PTQ5W6jQ01z+RfFww2dtW/p
AyucxCNSURYpdYeBJQcTNCs/AJA1AGHcWwyXQhMqO8/3DQR2dm/DUsKg/P+P6cir
XUMfpkHKSxFILYQElBiTslYGYEN17G7uYbej4xgpl2cg19oXnws0X0O14QH+gjIB
/Eu686r5NFzxiGaL8rK4yRSnNBgdgnopS5Kxtp6fb2GIXMKz46suqqaaCfiORgOR
/vfP85c/faD7afzLFTXQvtOdHPy6x6lV817yCsM7EVCTFXv3KS2k9PO8Xgcxly1R
I0aBAXu9EydTmQDWHLDXb1HKCs8ZHsNLRppn2+EIrNy9WF5PBhvHStr1wydfuPFJ
+gCr5Z0cV6bQ4m+UapC/66XVdZjJWi8HYOVm+PUX1X+k7oXhaTic+aDi/uk5xb6n
LXnMixwdf+s5lrgL7wYb6EywtsZNEB08LfZPbhtc7cE+wKH7AT57tdT+CofUYgTy
+8S68isjbAbiSOB4//EC4IbeVFZKtqzlZS/qHx6cLrn+aH4beNHb2sA8oYdyl4zq
pHiQFKvjbFXTTKU/nPOHO+fMR+QdU+Ig6MQrdSm9VjILS8qANZ0AqZU8fo8w++kJ
twRBhkcMdTYfQI44yaTu+iO4pEAz85MNKzV4kJKxpdgpc/9o+x4w62NU+sDl/5De
vr+jO8FBu3NbKmGANaOAiQ1SJYzExFp2M/QSTBppJvl2Ub/aXMM5ONe3d1GsLboj
zoBPd1MyNjQt+vhS8o/kePVgxcV+wcUjhNMQruz2xdTWLhYMajRBUPXyUv9+4WYZ
CEjpFEDrlLUA9JIpahEknSAiY2EZqU3/iunhH2GrkUpY0jnrm+NNNtOEYygQbaOJ
JXRKTYhnnTQnM3n6EYCrIlxv395XfcU9sG7AnomeilBhAyTpV+K4KZUUfAmLQ5Zx
9pPbpm+WNUdmiiszKdOjg91IXGkQ0kMP+6Wexjre8lfl0vp/ONKvsnr9rGXW02uV
HB+2jAPFFwQ2SGV9YL1bSenatXd0WXlO86/iX17Q90bCknSuC1aDhZMo4dpxj42q
XsocPdoCcAnWVoemhObXQQT6r+YJ5ppqZWAQM5GFA5ZC+ZtPylhyiMQEAqC9VL0N
iDbLKYsxsq5/XJI6LYvkzzO1Fjz7NeqCIOE2spzNkisawkKRBtKNL0y71C9328F3
qbucV1aOZ+d/5ljYl7pRoNDRVaoAb6dAQJVQTU1cS36xVz1JDOc4YGJ4CH6fO+Op
9vML/hMSWLYy1lghrrDo9OoUoeF/6jYiDuFtH6L/bO4RrqZEd5mdgdRJ8cYkIrux
zUFShG+NuvIx5hgqlPBSYcb3Ma5PZe78Duqxcq2pMjrg323WSpstXswNoYmKAooP
Jw6zeGlT6Q+z1riijYgoM+LfolOZYc4M+nHuEeb2Frcro1akoQkN2WLMWkwDrULa
1BUqFR4C4wQksnpclMpbKJQXrj4H2+Pz+N68LFV48Gc1oraS0YssmTpTdHBD3P9S
pOR+lTTHaUNOba3MHHVFa2glns38BzFAHC1CpXMr58M3gzFm9rtERYyVWlrHm9pK
MVAST48J4YMh3fkJRlzXF7AAsFyQ0FqEdRzYDOjq8Dj/CPTPv9ecwfAExEUgjjOB
QEr6Piwpf5qfv+0cwZyzQDbi7UNnMngbmNZbYBJ95MmA/rbhY3bMO0DNWfjnLnj5
uqgbQL4THNdhOPB+gOCH9BqcSqTCnDg4kbqKOoWcxT5DiaORGALi2AMPmq9J/Fw1
iJewRbPPga+3hESBmnkpGK11hPadPs+oZALboWXot3Qd2FBNdi8PVxBGOJVWxWOx
DqP/TtzM5ywSb6XmBXV8n4eTytpqgTB9A1l3W569WsYFMQ3szLSEIz17FMvpAqle
juf12mqIaI2Sop0dJg0SuDS9+pCoMJuceM1H+ri/PCO6O24DPs/51L3LyS629Srs
iZj2ScKlD+lHYI1B3WiCb9PLIUva5cf5iriU5dR0LCQzpA1PiwVra2B63juOvy3d
LHwaZFbclucF0YKcFnMNL8Vp6vBHHs7FAA1qOPw9UcN0d4yinKeeDJfL6qeidyuL
Cjr4kwoBp7unYmkvlMvZorgQxCQbXU1+zfn0xgEK39+C4rUMYsPvBDBe/VeYvxhJ
rE0gcVlDY2DsWPyNXyzQWZie5yTdGj869Dq8Nk3wF8eBM/GV8eiRbcEg9KzxWECc
Q6Sne19iHUDAPbWAU9PUCdDZCfB5M4NTLloKTos60yAozdA1S6pUoZw7b4d+3BIF
LKoI5dkDQV7wPAUZ94b3gIF0fTKJNRNLtbsijUvip6aSXm/I41MHr3MNqFCI9MdC
3x8lk4KO+wHdGlY1LGISADMMYoOYWQXfxofq8y3yFfT805rCVDYygnNog41BygKd
tF+DXtZ3Uy/ewJQaZUtlXDI4Nu5J143EGK9TcWmf8tnUfoGMmMq4pnA9ydPGBZzn
g8HHpy00WlWYTjnVmtnnDN59kEjpfe0p1Ru4SWhAtulzWfgQIOfsdqfSYP7WIEun
W85jpa8lr5KgFnA8hkJbEwFz16IL47/d0TOCIqlCa/gxQ2+JpfGwpM3M4bdFILE1
fJebgMERzM+1z5lxZAvtIOA0JULH6B56qQ7lqn4+NacWoiDXlGqniSFdWkhEufES
EPPxRUWkePX/vKTHJRqpVL/htJahRYJ3TMxVM6aKYxY9v2T4erNOkE0E8J99zH32
tnxtRgekGgtJ2IyaZb7Ir8WzQbXN6NydmOwHRnasFRB/KWDLIWGzc34Si6VpqmKz
gVgbprvJYyOpAbgnUJqDH8i9ngMaX/k0+JeUvR2O7HQJ0zVUdVCIu7TW+49S7y1i
62WMqyyTMsKYt3vQQnGuL+aXoJnsPwYXIBdSvuHMqJjK9/JPOy90ewlC3XtZ41i8
cwCKvRz1Utk19AHx3bG258Q0ujJe/mIBlrtragsm6h2w5r92WMGN9iTdVlQMTFcl
i++eGe8vUt6V1NmJJtV6lE0QdF4LK4NXGkbFuy86Y9QcmLNexFlMEkcFllV81TZN
OdTUu2mLQ8IelCiC6ow8X/NTT80Jq7a2HRCRypbOLpjhQ1s7thUo4VMA0o2t+AYx
9m+0gA7V42EdF65YE5gpJt41/euCi68X56ggfH5GQ+t/XhbtkBx5lwgbV9+ks1KD
fboQZpQB878vNlqB1TnH6rnHLQBwoAPWA0X+o7F+C51LkByay+OCC8UyDHzFvief
vaYRrpcPBVf+0rrDXyMmU8wQFHtaiZP+1E7aO0+p2PGNKrr9rW0LLuKNF2M2ZmJg
pTloMx56Ui68RkmTLA9CtlNodZ1kMhnDrtyNX1Rihj7j1XyJztlqri2dAOdv8R4o
i9LsBVdpRbW8BwSRf2n43DololSK5t/GKGC3qi7V72bb3lroTYEQN7F5AaiWF3tZ
X/XicPk5bLdEK3x8JoC1RJXIqF/MxgzC0gvhleQPg1N33JV6tZjrKJcrwTP9rFz9
APQ8ct6BSaM899flAxUt54QUt+0H6E482mOvjg+2dCtS9O9Ts2Eb56pcQoZbgH0P
TPiyA5jz+KBguppI10YWgnghR4MvA36JSv15nHd8PN5X5Q7duy8r+Tx6X86YGMXi
76EyfUq9OF8VabVDtDVmHcsisBLe1AQ0ypuoZ1P37xC1X1nLf0m3kdOK/gqW0IcE
6S3+Gysdi0Akf6X57ioMD8tf2e9CzOHGTTlzrpooOSS6vFL7R8iDGuQSpY+2xcaK
RkUqscXMDKoX4VdlJV6noYpZgyt1xfy90rmdFBf2RyeqXOmB8+OZjF3T6XTUajL5
BPV6KZw4forUHQjQ5jpcOvykvqoVkgNEQiyHAGfsdhHFb/NWId0tRfNPgAQNfWWD
20DtSOfteWzO93hJvEqAZDlQNq2MaMSYt3tsYB1OD6AF8LWqkPZZelGHxY8bBK8Z
WdbS66Wqcb9i+MoY9eB0gSTyNX8DoAEOE+c6jLQc/AvUpdSoNSKdeIa+vBXSjBPv
MNH2VMDGaPxjkN+G9QuPhF5pqB+Bk9iFJBx+e8RdP7Xr9DizGQYt96HL27jVWGSL
bQGPnLWR8mvrmqNcn1DzKNoZI8zzg8eaVddyDovnj0UNjipi5sxebpx7sutMzg58
G0Ifl2MrPx/nZpg9liWubUBbcNPCh2LTB2NDZfZ044/m2HXx9wupU1RUj8l3fNe3
x4IEmQC9/dFs7NJsMMhmJJNzByq8m8R4DQw1GaoMTxKnkidRv+qK0bI78UMCl6T6
us1rKZTIbpxvCLAGflXzEJv3PljNemoveBfG82EUfYkUFRoBb4b+9lRB2yuKut4o
6EkLucq7t3S2EIEUjJvn4Q693weVI5qMUXvJNJdu8aGluIAx9DtUGYZJmYHCGdax
Z8Tn2wM7K58ZljSzPn3e7dWh6M/qzBt3NQaonqEq86rK1MO8WgPCV8oAAxXXYpLj
2SEDRcvDg38EobJUF/Ngp4fANQM1dRfO5X4kAe4XqQ3W2IwaPilCq785uJMBJIQv
4zKVoyRfPbiz8MNIE3lrm/dLUfYlJ74H5erdbtPQDqiCxc6Y0FteSaMx2ahfabX6
YlyzHJDjgeJ7zyytDpyWEhlA68uT+HHVtTC+evgZ/x4l1S3zXiS12hCIz/RU/Smg
Ai6kUBk9EQGWj9gwLWqA4P/f8RgOEdnHwcSxN4jA6gGXzaQMN5s6f208bOrCu65W
LBygqWvq6uJN5LfVCEo3L6c8K8BezA3t0NmZv9yj8I7VxOXHA0NrslnLefGd8zzg
f8jH9AVeZ9ZWV5MdY8FCzw1b5iictEm7yF3sIWIvirN2ZINOz/++W3wnbGkBwhjU
bBPolKA0BH33txxkkJ73qvKEZXV0LpK3QasUARiaAd6/Ri7EC/EwFBMRi8PAMS2W
ct6HsBIMlHwJorvtU7STxC1jutuik+F8e+pKmmWI9Cho0mKi7CyXYK2nUGnXIUep
qWSMPvgozDujnHGzrdv1cgz41hwqYb/c2ZJk7GJcdLjmgbxcWViV8RZn1VVjlDVm
5OovQITUuN8TfkEqZhJPUg/YhaxKhA+swDjpKN+dJ5X/0i/B0tiXPWX0edAE9iCn
TOgEyVlwMZdPd19s2qrkHjyf1JSnCzzH3Ptw1THB4Y8kTiTqK4dNR/ax/y3EycCE
UZdqA70Db6pTAjhO4hThjRKsCro3W0YZKybIeSJUUi/il9IM8fMK3K6HtE5DH2jG
bA1OIYhFe289808Hnb5k2PEZmgvwAiz1umJ9sfZXYJSv7O3ujeLGiZloIa1TrK8U
usKTAAqIrJ7tu6D55z4DroR2UD1Y6dZBCjPcIhV01IAd1JuXzVjLi15r+bdUyPFM
kc8OtDi6JS7EXRN7e8EQHo2Zh++KIMsL/aK7HMVybydv7cZCFPfYbpJQ8RZEIR85
g+s755zl2xX9La1TqeO+LudywnF3+lHBwGmyolerXmzRMypjP6V3w8djNLF9Ivev
quGapuZXDy/MF4corXx4pji8ITloMz5iLhuPFtfmJp9b9sfKUuKcpOtpkgCq1sp5
AUifdjKwFeXLlh/N79f5viFfraoGOC6NaBl24cu+hOG1jLDBxdQ5IfRNr7qmZK41
X10rqdvf0yzxOV7WvAcCtb9McX2u9JaD6B/VZpxXfamxFxfOmoax3SGiTxT7wPkq
Rvom+SEadNOtn6hut30mcEjjV+S55l3S+qGGqGjttR1bTVHCI9JEQhp7qILAVObJ
TofqLeg9txjBwWgvjbZczthc5DVvdAns4OvvCtwt7W8MW/PKUUpWuG9hSFX4CBUq
nmApvsouUI9hiY6YQO+rKsOX+9ZKl0txJHlEgoWMJTGOhd966vRuM3XWIwjAJ9JC
A3OH9puYvtCxUCwpMES7qyP9QQ4utsW5lK/jmzFfdqEokAybfj3No9S02VZ5HQdI
jJ0GzkP0r4XH2C3uZBsMAga3PSheajwypXgNLORvg4ivIUsUG0opGg07K6baIY6I
AzJpbe9990Uqr8SJFiksYH9WQhyldSp4Fz1bPF6GC9CTFCTGETEY+SaNtGa+8R9q
BplH6VNvsoBSUWH2sJ+DE11hX84lh1hb3e/zE6z6EJ8K+DBZakbG+TWnv1gguQMQ
6jh3vh+RmVUtQZmFrVZ/C2aMYOO/U17hD9cJRVxl8q8fxUgqL7Gwe3cTXrXI+WGT
2InFfIdCD5UDMWc6m6mZqR3nZIcgUeNSCcO7BE9n+FUOs2/IHf4vGiDF26hs/Z9g
Y1RH44c2SGjdUnvDS1se7tuy9Kln6j+yardcjDqQcGRBcIUZit0AIi4PsNr25wUW
3Kb6O7nh/A6z4OJrh+IaUsM6LcZxXJT8LCU9INZQki4mTbH24ljlbzQQbmVVNGjk
eUFJcZEVIPQ0/3e/UMjhoE7p6MtkN2WvDVDpnJspUOBM4veYWHODUGZpxwDayKMQ
EC9Pv4btnSgrgMKDdVetShwygAeAmZu6qGE33ZuRPpzdJk2JcsmwfftvXOfFoCQA
N9EYqz4WgskT+2lUTjELMJ0Gu8M/aOLl1m2PGU3jFNlMm/ufuLtFxsH/6hAJzh6s
nSOV30rtqHKP3UMkgozpTm95qpcXdDRLYEQ8FskRwPDRorzNtcms/1nIkg9Knb85
jcNv+0IvqMs1WGwYaEw2ny9CEo+FpUwsCTNFCaApieZsnzKTN73i9i0EglJIpJ54
EcAyM2KaqPR78PWpyGyXnvIV/EMCfbXjkO0lFpvwjAyG8Xz1wMkz9xNfiGTGoDKa
GQOm8xMCss4NKFikuALl0BuwXBTE8ImqTwioGWHj4PwwxubheUL8hxNdtSpfYc2p
GvTlS3ckQUXes99HNuV8lsiBVFft9nLoJWZKQVYhvPLiEtRBrBTK0HJhfr/Jd8y/
lqCydtnCNu8DuBcNI4NBG96noh3kzYPUR2Y1JsPdcIrjK7l+6YcIxbJb9nFZD88O
mNEIy+GJFzvlm/N5xermCPqlIvUMOEdg2z4GqnBZ6hGNMnHwUNSGzP14/NSonpTo
PrCWsp6GkRkKThYUYXrBEu8HZs6QgMbf6o2MvrNOjCXy5UD9CBr8lTlsWtoF1Lmh
uODgf5JbP7ehk5cMKb7rOi9bieztt/aC+T2LU5RLSnQEvfkJ5DM5txRvoMQ/ONxX
xfDMR0G75E3ni2HRzZihu/1tMNeboGTYyFeX7tLr6wHQHpoYtGAnbFsn5DM9d1rh
OpHiN7MMMOwYZfqWFrZ/fP+pAcru5I+tkFtOHNtl0323R441mu5YGBPvZt+K9ekv
lA7jrzGohR9aszNVHxzemxHlSXVHydlEQ2+3Mcm3ofVsLXhlbUe0vMoiL4j6urff
zjRCN/c07xiQvRBsSibARHpJFg2yTbuxUBbddcrLGAcCV/d8N8xbk9t1HK1MaXtz
1M5vLG7aggm5aLR9zknedtzlhmlxlmEXVYLUxdfwk8ccUS1GXKGKs/7xangsd9tf
wq699jgUPmEZlECh6fKT3JNiGH1phErLKkPJ9R3tiMZqjxcOIcIdQL5slVXMzbVd
4wxfhq8vlo+/M9pPu3QmXGZMH1wY8Uw6HZ0xWdqdQaUFEWz/+DHslIK6UmkGzaD2
vp4cO6reOqfkLw7LuIQMVseO650uFjqjQ7uzNtGbodViivDlMmRmJnyIkaNFbypS
/NH5G+2lH/0b+XlYWvt/uOuGI7OAjBLDOxjo+Dknc4byA5XaRM4n5BPIon6uZfBv
NevW924b8PWz7uCYnZFlX/NVgSTsZj3xOtwXfMklQXcAm+7lK9ZqqMJLIR9M72/c
iFUfgBJdLzxkk46zHfWi8pCdwgkOOSQuSbOLdQsjhqVdwoi9WR3xfBSTQNTq0iOa
h+5J5qFuOe8D87eK/Fvnds8TYEHKcde9ChfHzmZGjib+3e6vKHe0yBGF4CDUgQu+
j95Y/5rnItLaaMe2WWUi8Ea+0VPfS3eGUtZHhI50dDhbY7LvltnZOu1/RiwQT6lE
9FNUaiPVsOE//d8Ejn+ZrJAYRDV3CScpcFIUqfKYWAUnBS28NjREDaaapH+BgYrp
Kc83t0ecr6DInEfbmK72Wb0w3w6NONqmUVC7Fsp2UABbdrQ7k9J5Vkbmy1AYROIg
yz5JT8i4V+3ySYxPmS6q7t6I5P8O8AQ4Qza65aq3M6ZQvrFAafYK2a0WXjDYkuF1
AVLWjM4eee00/MZWZypH6ZFdFhui8Io9s2X/zFZq/QM94vHSr/FiO/i7nM7+/odA
arJI3FoVYtoffVtAzTLLp+1vcoTr1ootQNp1lG0ZmeQ5CFGBORBHMnG/YoaprSpE
aWhy0eomPD7+r9/fBHtOPnMTEVNkU+0cNcIY8yIyV9wniwINzm1rm7U3eK9TfNFC
uUEsNWmXWB6AJkuCUpyypw+thVrhyJwupatwf0SJfAHoAbn8eQ0JcxY3B9b6EbrM
A+RMexLcXHwYM612lTyCJjR57LXjsciZDpA1v8r/t2xcUebYzuvU5yY2fGroSRHo
UBVY1I13DzOXPZNIVra/PcGiYLFMfX51ZDch/ET51tMMlgmtCftnEqecH+jzNfUB
5wFmfh/rOs/TeMWbYONLAcpBOF1Lr1zx0ZmSMTaH003B2srkMljHD0XK4j/kEHEL
Lc+ZjybDCG3Bn16Vyhn6yUP0xWbLM3G3h9On+mLfHAhhTydrbCjGIgx537XPL2l4
XG+Ps/QEbLhIHZaqA1i6CxbZjH2ZLmTdbCGM3EnYzkXf6bOqqZVMVAaRF60ZFYsI
4xVCNlRIeS9RJrj6rB2pil8BkGf4IAtpVRvCXXDKMN6McmU9OGPl4rwZ7qh9U2F2
RxNqochT/zAwqNOaTCnnT9xggjUenXMd/ZF4LtXhL8kdm3/NIKmEO369Yjuu94CE
BgRMav5tP5QvUfCaPbVoE2thVEXacotQATU7kGptCh/CHCaWFvDKMU7XGK+9w2O6
D+8KxQYaVj/ag2FxQ5Zosb5b30zfvMWRXDDS9B2x/JFJd7pPif2FI+Hhtz+QR/jR
Q41+QwG+jAegkVL0za7nf8WkR3XbXeSlq9QbdTZCeiuk2yOVRSTw06dvywmcjV9h
J7tS3miU8RHkYSjC/cYpX0Wfkv7eshJtdQIOo0iBj3qgH/Jip0JSXaGqXy/yYgdE
uY4zYQJsWZi5526H5QbGlxlq5ERlYvER7IcRuUlWEksND+ADwVXKoexYo+P7gbwz
ViDjk+4sPw5dOLz07bZxgINqatSl8KDu7oXJSXqisl0Z+z2cZjUyYqNJXbzTTlP+
o0kkX0oJ3DcLE6szCaPJ3FXTVUg/GbjRmxAzOaZmw4dZ3FsUIbZTcalCIl8J1qM+
gPWL7UPRq0csQCJ4FSrWQrHAs0Tz/Sv2lAalImuAh9JvoSFb3CpI2h7jjVVhjl4j
Ld65mPzziW3rMyoWwC94/BkahXbl/1oVEw3ZOKfNZOhZHJCviVMI5M/oaadMyf0c
XpfMhECvlNlQC65oSUruWDLZgVkmw081tmjpMkgQFBYnbTcmnahoanDkB2kiw0vc
47tmCdMvWkWh+L7lACrDUDOzcrRq0FXs2yTI14dIJxrjHu/OURA+Qa7vKu9lmFOl
QOxbCzg6gTJ0OS7L9dPFVaPJ/SygOlDdh6UBKhottcT2OvBOxQw7qM4dOVTbo9/v
KamOKgwIuAD1aOVLB6sYNRZXbKIiNLDy7TpBgJnS/gr3Z0DPRFXDavLdH3FxiEgY
Zb4oxLgcbaDsaNREIhJr6DOCxc3mqaj5N5cfFpBdt8d9Mkh8SuVtb/iDyhcdYOAw
dhkT0p0+Ycl/eYZ9EHGVQEkSCaOTFP7usyxModsbOOa8WsQn4tbsbZ06hcZLSg7P
/8GgoiOTr56wybPMWzWsxeYY88KTu1KbAXl1nut0e2vDi5+RCk5nEnWDOZPt5zK6
hk4tj6zSU0gZ8/2sLP1YgLeFmhENbxJWTDGP3xgAZ+dD9ovNAHO8WEqX2V3O/lCN
XrlmzCNPKUVrpjKvkiW2wZcrWw4maLdEZI2kRB+gKIG+/QeedoRv4gdoFSsDRzp+
45J9yq8pUvCXik7aL5QYZpd7wMzJgbCst4fI1AheB7T6G42XfxGAyIkc95fGsQV1
Ts/yXTmA5vyiVOWALi4LwqEafDXMPfUqKdFeaDARuTiXWoz30+z47okrejLRQ8Bo
Rz0CUglmHHt0Z0rKZEwZr/yxu9azZupAIqk3gcHy90T2ohUhoBVZM+NhkIUFafPS
66y50rz/709fmXdeEXvMT1zr2LjuSJ60H/c8tWnC6bMEDrp6sG4ZGm6qe6GP1jaM
KFTZasG55uRjLKaaSyH0J04XReftb3ITzojzdWg4DED7CMyQi8jkFW7HrpkkgMn9
NxebQc95ImhO1Ljbdsm1h29kQdYP/jKn8JONck8AXvYsnWvRy2MKv8pES+l0J2Ue
RuVZQB0uiZQ0lde8KNxQv1Fdbt0aPvYB1zkuzgzzRbdp/ExsUxoZNSE2e03t/Ehp
2W0O86uTwHGPHQx0axaUcemCgkqP8uMOnJx7Fpe5HdNAp4/Z83y6JEkmZCNkMc92
YpkuzgjLs05rQm6eOqBjkjg3sVyr29FHqz/AnbDESVQi8CJrp2mRVqMe0M6eGPzM
KUTNwT2qXL9Dsp0h0IF8gwa7r5xRNOqNi2GrsuDkstr9DCl3fVeKLkq9KIsKVfFF
prrZiboZeAguNSGWQMYhrzP3dMbKlg/QSJ+t0mfzI91dGFol3mrfLehNeKZTaKOQ
2/xjnHrjpKO6Foquot6J7TwzJKdcV1KbHsNaxyXa0aivlAMYu7264amMWVxvmZqS
XlsIyE1i61qxKVn4VMujh3eUUhXUsYa0/7BA+zYppX4Y1qsAU75FApotr/MgCOlB
+ANZFiNsS03pdM3a/p+2SDq/B+bP9th4bUsxEj5eAVO9+EG5VHj3O1dH7rzciE3G
SZmMSdVt3BmEFqgw16oAcp2eDLBTJ4JDVh8RRx3Qbt2OpwCEPZmIaQbPLghfZRnX
TMKvhmP7EOXiIlYpjQZg1qKQ35hWuZ3/NtNAeeVrf1r5olCT0hOX3/kH/BdQA1WJ
GFlJ0ZHy67s1CVRtgdY8pWY+XTAi4Z2EAtQnspiWMgIZVGJtfWxRqrcH/CCOyt2G
Ropfemmmp9WvsJmIw3Vse+ZfH4Op1O8Xj2sfl20ZIiwinpadeCuSaYKmCRCPhvtw
PcY2OtCyTIRmk3kR27qbVaXNZIgl9gFXU7dnimpT4z732DtprkNCYtPnpVirDlNt
P2MUT4U/u+K3c0olBvU3mCXE1+F40bEg2kSD1/fYDW4S05eSPH/72XAHBSSicPY0
vUnDbuv/IU2RTKlK61hwcEWt8QctdYfTcl4drxCdO8kThpkMwOFRMIn6hIz0D/wV
0uUfs4nXtMVWFN5p0LK5g3uHHcrtiz9sZ/frpSKRqjYqoSC3/XwCgPKkpQnLt1MR
1xjSeQP78gzuOFwXkwH4NMRTWMT+9C8/ZCaoQz6S19IWVLRP/lZGD66JIDdgCyMo
KP6+0XWu8NrVOOM3oVowfp2mST+nBuocetKN1cOcscE7lYwOvF7o2spoKiJhMZzr
hOk7CgzY5Jjbg5/PQpOhzNX1V8QuZxEMYEzAMXmbM0bpS/KYTHHlFQrL3wdQIzcA
eiQ3ZG47cW2n6eUqIbDAvA2KSGwbQwAhmSNTdUGqul7jCyHApGduf44bA8+NhAvi
IgKOfCBLsZyfhAqlKNjxYeH/wMdlGZU9OEECZto4Q1K65vC0zJjkBKwXJO1mO8Oa
OXDl8EjmbSm9a0VMPsPkvknw1zKIj8W3eH+wm//KBNhlSi5DT848sB+7RAeMOX+w
ksy0BPPYtgef9vmZCBZdZu+Ri+jayEFbDWDLsolI7D155gxvjeqiGc+RJtSuUkDr
v+Oug9ub1iGzrdvLRzHWW4GioempOZOQ20v6Mt3UquvytHrEvqTxi+SzP8ewIAJE
Xp0U3DupUR+I1IE7WizRi2tYsywFi/61F4bfol4JHwTCoAcIDvyagAv1b6rLE+7i
lx2ZxpOjxwNNBatXry082YTwLOTYlJJXAv33oUv8WUvQxRl/b3KBq6tFv5f+5858
87a0uj3nbivfYVvSrINxdBEeGfYdwSZm5Xj9KA3oDYGpH9Bdnb5zSiCdYXSwP6TI
ITv/EAuggOq40bTrGoUyO9pzHMxCK+9KMkAJ6t/k8KZWLJqVJK72q1ZTWz/jda6U
NEanXRNcERCsvT4PsERf//TOHmezV6iLqGnF5IweZyC9BqwzaNHvA023siYMriEv
i4O94PJVxcl5ES4H64kF5MmQ9PVCfUv5Tt4m9NfqfUe2KhjJflRlY+plgBwMdsjW
/TgsuY34nYi5RiKiDcrxhjxseFNI6w8Us480mH2KXfXl0uXGbzv1frWE5lk9hXQG
ubm3320xtCM/QkPGKOHdXk+DsxdguOW++GXbdV2Sq6Ne7aA/ixeh3+RIkgGeZSoq
FvzxM3uebr3r4vblGxfA5GadmNASxWagjQJXX8EByrgwakHcKJPkv4+IjQHe/9JH
JdBezOcpWvel97TS5qWU3hhK1ZBetZ009997Ye/RkGE811GV59IfZYx86LgufPxl
Gck97wes/NT2jE+Xke5GgAfDpcHV9m3m4SAV+s/LECkJt6cCCFAYnv0ZxEThtiu5
Lfnm+ApPMuK6v38PunS3hZm0Ut8hLp7/DJ//eCx52VFzo1eCyfNoglWrT3IUvfwx
0MKKmrgDDCODNRR6Zf4XcfvNANKHLmX3E3tbL51cN9N7gE70bBc3GG8d/jvzWF7C
eV5FgR5Usfu5st+z1T/2sWAk2D1kydX2vmCTU4uAEZXAKUETkrRlmn/qgaFo+2XU
VX6+6CUjJud+li2RQlz+dx5GHslf9BwoZVNkrYq/iCOysGrXQRWLTT5UjreY1WKB
IoBRLm0q8pS51LywKzJ/76qErd3SH3JytRy3iy+q3/Jr/Q9HDg7MaZtYeD7obK53
NUPTmvu2Tj+5bXbI6Il6A+6GdHnQP7rL8hRJj1TyqEVV05yYQWdYsmTFbl6lpA4i
cBX84c8q95n9a41TiIwG+JsZJ7gBS5irDdtkyl2P9dx1YwgAAQlBqi2jWJuMDYmz
eOeR2S/w6TG+UZI0ESpRBki0EV+Elfirk01n/iOd78q5TIPAzNL+NCLbff1haLCq
vKUalmqDE0YgszbPGBu5UXEVxkJ/XwruhaKctem6l/hCKgZHwb1fOp2XJtq4dxRv
ft/tuzF0SgDJc80MZA/iNuEwvKL8cdNSIJoSz5Ub3zDv0Mtn398tL2QPfBo+bmLB
4qD1eWjpdq7MPLbALzYk+AKVIdzM364YIFrPLVsia4PYM+rnrBbYdrP+pYPYKPax
UHEGxTk/2UvlapxFPoHqD2oSZ4UBwrTPDwBWIg1BRqltXo1UkDUEY8wkk3zAIqBo
SBY4U04OAJ19YqetXYhFbJMkHJuNDw5vw1kXfSFgCFQli/zLtEsTGCh0dfpYGHiR
/VKgop1gJipCJNZVlLK7uuJ9F4CgcJSACLlDwcwmgZwby2iujeOToDuPDS96dLxr
ttMuTn01vEHvvERU8H6vGlIPBu00oNz5/DvOMHvOapVvEPlnFebNcl8GQpA3xP+a
S6jcdrPaXdn/Xq6ydXUFdfGKN8zUyo/uE0v/Zi7VYzHzTWs13K5oV8LGova2/FdE
YbXx+lAMHFNXBhvInTxhpmCKSyU3u2zRPpbDNXpiubIWZEM9CKraY2zgFEatSkza
LGYIyLIuGnLOcDWN966YTL7aUhky1gDNzc8XWnUs62giGTks9FBedDEEToi6Co5B
EWsVxbsH3ZapfR3tm3QAPUudxK4iacVLHYecWaLcdxz28yGxw/MDYsyq7Nd+pKzM
4ZK/RmVRczTH4cmpfGV4qet3HKwHj1Lnw5rRzauNZXAe8B49F7WTow/d5+pzH4lD
nzupW8pRnisuLKpoXZWZWcm30ty/aH+jZq+XtV9NSGMPwHyqhLJI2zT9AZiscF5N
mgcszoJ+pipaO1vat1HHVoUfkzqEojqTtanwnVHp1GlAbFj+lfAkWF15qj/XmXBb
SUT4nSWSlmR1QLUkdJyqNLeDripwHkuh5TZ8rEaq3S7pFqC7dsAMqBOqegP16GUS
L5NFv51W4ytiLollyz3mBxW8cvH2wpB4rjdo/RxHY5swKRJ8YI7OqxTWLVqCarHT
dfDDoG2vtGw1gXm8nqiRjKVfDT056b5FVl6zZH4HGJ5GjwwN/s2YuxbvT0GJayhS
6fukLf3g61Gj3TvKXEMKUmuoQeshGAS4DtDfmxislBu1nIyQgbJVGVQ1n5ILdNT2
BGg2hB1Ocj4auTQ9u+F3fLeJ0/Oe0MUXj5uX+RdwEDhTZBgMHaXeK1BjVV46CgMh
HeVMjvXCyLzguaIklQ023wjZpmZRTx4aXAXbs1+ETr5jskVcoMEZwYsQ5XusHsMW
XQVvkmFtZYJ2wT7mZMnMqEHiUjqyg5oZWP0mjK8QbleiYK0md9cEvNK1zWtMn5kL
rfIMkqQR6uvX+136+F4Iysatf4nMPfZAy1UU9QUJD8sXYGGeSPnQV/35mM1Yfuzd
ySD8VxmWyNN83SCKxdDstLMtYo7lD8JLIQHqeT4AbPF4/Ny9ilCY4Q/T/Z3PxsIe
K72jhgAPm53fvJ9VHlSqP1G8xOLbWBUTgbfOXrjj4jjH69yZKWn8QErmkcH4BTMZ
6rY5uEWCDOT6CyMKFNx1lR0PyVu4rdfdFs2xcW2APSYxoqeuAtS6dgkXgtGcEWVa
IFt0adLkqlKUQHwyP6q2ViBIWBU5Bx0pm5Khfu64srYRVqGRghWO2CH+e+feerl5
RfeUCJI3VkJv634KLXzWFnYP2QH556xgc07foBfPPNoeXcH6yhPbCBZia1BCrqTd
WcFaeKB76moUokRCSnqOkmWZb3GFie3e/MOAIh57YuBw8rE4HbEYnWN6n7P511R0
vAgtCe6RytsKRvPuVr/2yYya6T2HTENR69VIpbw76rN6rK+LrDpuc25RU3MLVFvp
Be5wiYuRgZDCf0qvZSBvLXx+NssiFdOtg7nOID8F0ZzSKG6XH4kss/1aYggFpVAr
urVahUlvDlKZPIKOEgSi2d+ifSBRMLFsuCwFSci4wDeFR/uM1TocEOmVfHBexaXN
+Zwo4ojWbUwbp4M06+MIzUJC0m3D8CIFeUdwAfnqb3MeaA07iD5eTdNz//M/qvd+
G9X8Lf9pBbZJrCXA2lysBCW6gDofcpL0YXMLROUy5+u4NQANVyp96OMS9gSF8shj
LpzAIV8/+UCmEuAhqoOogBcqRaIDCeFEe404fg9j2ENzrQOJvsHgejLzYxZYFJ+4
svu8h0ChslkRVgWX1w1Qfe2IrQsiIq3JyGP3aTheMa9lmUahFkNA6RfpdSmCg6F5
/XLu2k13slvh49gpa46zCfceUcysLUChy1/8bWiYbl0KSX3x1Gqhs3upt6Ut6O9w
R8HN8j2Fv7BS0vjR4aj6ytsMdsb8btbIJRLZMfczKHkdOW9T2b5K9VOUU2DaWUvK
TR8Oh4OGX03Ybqo0qQL3XI+GAUjrTtG/llNuLYhdkOdfMBuC5/gmmawrmLC89bQK
zHeRkedTi8nMiV3ivFKx2cwD6ilj4x6GfDrVH5CJdjrue0DtnhYFiAZ2GxCX78Cg
1mJKQANdDYbPCVEg/LrVLGrOy8Cz/A6J9/SMyMW2Inf+enlpKkGFxH/Q2gbnV7Jy
2G6zZuvMeqEZLdjaFSY8MiGFONtIQ3hEgUnwG070kDqZN7JQwtBYvDU8vP73pJV+
LeyupmVnOTi+nLuswZyHCmyeiiyh9Ok8tFGg9uWgS9FPstWoLGFJG+rnk8BnZ+k6
MFHfgvW6TZPSp3fUbg5Loh1fKdKyjYHmiNM//syU3XySS++KdU+0psHvn+D9e1MD
wSgdg+Ymw/0eUxbfnHEOl7x9QJpTebrWrj0TNC3DgJNBW738rpbvPfABdncC/lrX
KXEIz1T3MfCwA2lttOqGiS15e/xgKtWZD2S3XUhNF9fgbtcdMWmaYs4r6E27y9iL
nDw+K910FQ/EVtCuJSl2s+Pg5xIPGu/ivH6GQvGhPcKfR/lyiBUfeItwaee9n35r
C0yxL92YQeM2UtI3sRjY24g30MrLy+GjfxHwIfyGIEe4a3/mVJtl4qMmTNG8CBA0
b74JpEQMb6z4ZCXv2A9sHdVQCrb/S34FSxqHShG8Nk3kVTnlJgS42n1L0BTWOVtV
puAei7/gFhhvEww6RVMFUOkQacv5AMWuSfNnS71E5GetIqQd+N35vOGUTeOvoCIZ
FNM7uxnvikRI3yaIFgf1iCrzip0OA3Nya6h3N/kVCufP9qV4PzGOmG9V5QQVQFyS
S+ldjZAGd69+1cKPArDJrb2oCJCHHlqOljczCiJlijo4iJlgkoulPcfGiVRc8W8/
q6N8oZ9stg0cvTKBvda1kPsPgjcCbGhvvHs1CmHG1Gtmoqd4DBrCLzWeP4oPmzkB
CS37QYw8efKy42sAZknzEgFRflPbBzZOQW9iWE9RUngazUf7sb1ye85seEZwYYLP
A8v28wfc0dpiDMuDc9kDKu6sp45US6ZmO0xRwVHkL2NJNe2EaTb0kAjoXhdvnvmH
/BvJHEQN0GrWjugEhCCbzIJhbDrgv8X4wDb7yg9CgL7zP3FbCW95GSv+3BLF7fBL
MuLlPPX73ZHfO+ILSYHgTceQXU3ovklECmXlIyF+Hs6GHP0eF+i5KFFCbZCQ6RjX
m1N00tN+L3UnUSc+ymmFRORR3IVEqN/JsnT1LrvpJyEHEyYNYkJ/ZVuRdNhJYlJN
yVd4bQwH74S/9x2Ch+n++nw51+DfirT+unnwk8S3+vgKodaFzdiRoQ/lohCBzMj4
Ag8/dH8pGPGO2BKzOdyyEgJvLBSVeQsM4fshmfeqOJPQEdwNm3p8IgIF/3fPckL7
ptvBUs9hicvWXqhTkDYZ1UubmLqzZ7PHbyBct8KBVQdhrAchA1J1wxHQMEdBKihc
OuzxQTj+pkBN0YdbDII/z8PyVq7B4Wp7kSxPEcKHFTpPoeu9T+9gnOkU2n6qQbjn
7TvAD8LOTsw9FvxLq0WzwO1IrNFYN5Sj9aBLWJ4QNFx87A22A4xC89d/fWcLoavn
djmFzmMATueNdCXrQgH4Y80QRE2CZ/PSJ1rPDYxl7w++kbJqMPFGS04+c6HKHOHY
qZP8N4+/Pu/Wp9+6BA08AaMsoYQTPw4wlfNs27IOJ+Ekvn2vL4/wQdhS7vVRnJUm
QSQ0bV2vSIKWgnoeMdqyFORdTjwBbcf+uWqVmiC70TX0v0lXXYFumDkqEaOn1AEj
W2fgoapI2ufnDlfQuroVcz5V+at0tx8d8sfjYyeCOZGxAHUqERglcHRBQE7uJiy5
fU8IMUGUyoMCkMGASX2FwEumUNSSd29/rcEXyn15TMPfxBqhAwESbUdb9KyyvxE7
eCyU35yMix8sOFcqdpy9Cyc0RGAhN68SOs2CSjzr6kBNq78Eax81Cr7UskguvmJS
4c3rfPmsOftzJ7GOywsxOlx7MLOR0GLtKt94HrwbMdkv74CTtDwaMlOf4KXsSHtd
IfB83gb03l/vyZKq8OAfDEPDQKnPMcAYfEuXHxDJCoIUEhOXfE+/GriLoCQCfGdt
Fau4ZBKPlnxbJWyu3sgrr+MXwn7XkiM/xNyRi2bgsVjUBNnUU5Y8U+LWmIx9gr9F
yQwq3L2+/g7WLGAYPNfYWkzB+I7xk3uDGuJikVMzRji3EHlyKYGNX7afZK8uHaiQ
iMWMGhxjseyy5iK99N6xLc6zU0c9RNSDqlKESn3c1jplgHD1dFxZlSI99lXEb5DT
9f/n8/FrrXT7MT13cxM0Q+nw2i10VcrJphNAPxLhCJ0dT6p05z3XPwuad85SMPm5
aZwZsj7cVD3JXfeWgN3w0rr/4+0a50sApf4mSs8rGdbnfoTa2PKbXmB9ULkzcrNF
/JHxPY5zy2u9dB8tthv3raJuA+xVUHUz08hIDQRdzYESyjk9b9qfCRJXVZsMNQG3
gaA31sGYCjfao8C8UnPoK3zfnOUUqX/usPPH/8JP22g0qf/KEDYSI4Ilu9SN5liV
BItNzLNC1vtkpHtgeF4WbuUwEXfQrOg+rShXZwRKk3RYOrxM7dmuF1WFw9z8FXn3
TxZVvru2gm3wcK36mBS+J3V6uy0rgmfYTzVGhRQwecpK/28SVLS51pYKZNQ69mjT
PBWcfwSjdCbEAjgrpXcq/rOor1GXyNjymdMk/IuJJgX8uGcY32/iPQqmlSRbs743
wfisJzkw+q1IujrEjTFVaFuWf6fdRhCGg6kkKybS4YIddFU0efItMjoDSpVE6pA0
LrrD+KnINZAbyAQ04UIeBy6VBxcKPo3aICswHlttPVzx+YhaSnHdsI/mI4h77p96
K/yBJCtR6Uw7lOCl1wZSMPng2Bab81pH5HlRUwcGpILQQyjeRzBy3nRb7P8rEAQc
jKv1jbp7pQDheRSjrLkHLVJRNl61niqog1cvucyaXRadq9zJKYrJNdV0u5IZcrXx
QdAEzVItKQRnW7XgONSOmc7HwM1BssqTh/YEeK6w7t8TQVAFy0L/Frv0D1t+3X7o
/4CGTW1PPKV/vlfgy6mPCKCxlVgumb3pQuU/Gg4k3ZuTPBng5PFZgAvYwXcRTG5j
7WVbYc+q3xC1WSZxzFJ+Nmjjz/J3uSOtxNo0NPiGEEjPX7bJ6jmCX3iYPrtL1UtM
cF1Rnz0hSt/RLRxFMQdMdxSZyoZ+6PHQCeoBliptgYW07JIFj6kWEqSF47PCQUs9
pFKZhYlUkY228M3v3F22hbWGuaS9kpR0SJ2wej9qQwtF3nKfiJP7HDlD4Hx/bD/P
HgiqEoK8giDRT3l+wyF91g96GZ3F7PXIHwL1CmqHzzwumqBlWfU5L3XxoaW9418e
P7of+P87pj2fTDHZSsA/SvxxEbE9eoToUGEn3q3H38o2jKUuatM2M7+Lc5HxfMTb
bMhp8ffYSRgfSi5nEPGDsQa5N5x+EwiZIhr7J7kjZAgS0wFjTqnTXNWWDJAay2qh
HwevXxI/FFymjBki3hj95SqEeOCkHgQTx7Z+Dpgy051k6KjsDcoWdlWooxV6aogY
AGld2wbs2WRTfyWYNfhFrUKm1DmJgdoSjziaVI7JwA2gqaRO0nH7vxvuyD/Pm/oT
p1RyZrlGtm+nCk0NEot3dSs5QULVHM6cET/HmWinKyie+AGi5xnj5/ndvnyRenKq
cBdI4lqjQ6QNkp31dU11hUqDdlo9IAyNf7v6VwkIIO6xXroL3P05xNm9QqP8A8MU
37DqXbEs1utX8MqiyQs9os4JaUYUCTavruOfU/gom5NVamuJgtjiQwN/lyeP3szq
+Uh2iZeu/I93jhPrYtNqZcfi6jlfdDcGXGp/sSKsPEWp5ej+X6r/9Y24FySN8Yg3
2icJA6N27YuMCqZXEo5TugsxU+NmGdqf+gfUtxSHT8rUgZtyX7e0NNSRBn9aLna4
6OJXR8CY0mlDGefAX4EATZe8BRfl++npQN82iramEtfHWmnauz+xu0a8oFv2m4Sg
1SMVuFF6jWJcEN1kWblXEoBC6PhbR4TrFKksDbHFXBGKnVdqMnh828C3i1ew+rhu
Hfok5PxlTIeGUFTzLnrL+44koXA60CZz1oc838ugIWUkExDfq/q9piFKJTBNorPu
GHugia+ILiRgKCFqx/VI4jiVeBe6VnAWZPnLLOfcTV82eolmItISI/C7NcEd/NS7
a8WvzxZgPQY64QJRblAcoRi8W1MaRp4uaftnndmo2xReHOEWMmL361k02CdNsg0i
uvLPaH98SDC2qW598sZcZPMeCaWYpbfLQjxESlJLHUnpJnfxQ9CAag5yJGuGDuRl
flVdnLWNjGOuUdlAcrFTqa17bLyAZxeW+DHh9/p0GA9HlLIwp/AMRWgQZ+dKe3d6
AQOpHB8gbZr6Wq0pf7uFqKHadTncizkYAOcwK89GvN0S2vwug18/Ga74RSKriEYX
/zWWB35yjXXnsmAc3KQUcmr8OZmU1Ldm91amynVk5xauME8tddO3AaP9edlHd884
AGzlWZvUerKj4LMdpIStNpD5tJf2aAeiYcFCCkil6+GMpn4pT/USWyDzuh+jNuB1
6fVd7wJ0TDwIJqUwNELMDDmTqybwTKjB6wqNM06pftdPLIRfZWPA3HfD5F7dpHZ6
g8sGqRvu8aRVNC2FZQuI8UH0az4FabOmoV0znK3McUIkGlcS33O20h3Wv80aT1hI
Zu0H7vp7+bfXWdWAMRnZJgIuCFUqHwfvpb3rtlbru5JuspmwCDr55XqwQpfRvO/8
rOkYTBI+2zzsjlNjBm6RlTUx3HOdaAwi6b9OJMfUBwCgljx/j+dXb2xqxrGU+Jum
XSkuGct0jlLpVbebtJj/GOhpTKveuPt13FEhmkXIPiUMlqSPqCafYU+7Mbhe+1Vn
fbEImrwChoIHw90bX2gNvBWO0PVJ/Dt+TWtS8gvYYIjMPtqGET9KPeu2BXrkBj1q
0XDkhSLUsVLoI9ETGUX06vyxjyiVcL+T7ZiJUQbs9gEWLLuQA+no+8+N5wu0W+uU
bD97SZ8asLFzwNO7raa8qIRoCzHX0iHJcboc9DzTi0NC8SawfQ/4ZbKHwG30CWIk
u5aZGSQUZHhYrF2l8IytvB7NMzA+V0AStPjMKEIzzcHqS1U5lM4Icc3zZoxSTkse
h9Y8KDkxHUjoaDzq47Dbl7Xzr1sU7LKVqx97YFNrExPv8e3Tpp/U8OHIK8o9FP3b
fUPfKfu+kBOPcKfNgl6HgV3owFZklamyd1bLcUL2X+u2U1E8lusD1NZzlNLGN7OD
/3KKRnju9JjMufIUSO3ZhV0ULOaUHQHeINH7lJFD0er7oDR0B7Z2GL8ifRW8pATY
VaXG/ttYVitOYpp/gZCr0lAjkd2AGHZsNSBWIKdwz13ih5UxXEVK4BFyAWoAIg1I
fEmiuzW94iLrLWPWaBVnEdSnyMCEWEQg76wKt5pVWxdwkAufKEYqRaQZWq6zwZrQ
UimHfz0W93Ifq/j2YJXqfO3gsDvBbDnbjNzY/aRSSgYHyX4clBuzecyhd/nyqpXM
Jgg3Lmqbq/LZa68ODSzkckOUG/S46g6xrda81SotD4l6STm/K0cAdoYTXMcbauRI
nkNDHgMZwo8jrUAo+m0BcaSiZUGs4qSydOrSlSpAUnb5KvJmSytNK08G4p888Xi0
HWeE+e3xoefSPJH+MGdTE/qJE+D93b+85s2ZluoCsBa2rLK+SHRK1ekO8GOjQR9P
i0HQ2UEXj43t7hvIk1bGqFEH+hLxy06aJ2n5Ko7nFdK+4dGTF0W5jJwBJAJPWpZn
VUFkjUn6JobET/YDCWKy4+iybhB5rnDdSwIY8QhIm+s3xL5pjxmg7LAllUWU1+By
YtbdTubvGe4JgGTbBsSWRpyYmYG9acAKJv5Zpk0DfwvMzVTWgHF9xGZ89vZhoqpV
OIzr3tGKqCdZB7u2rWjoX2uA2mW4avGjnUPjXj9SvY+Py8iBZS53Dzf5GlvaaLIW
zpMuwidVH0kdBHySoe3LvaJ7iwgx+KQjo7yQHBift3cm5B7MefyJ5aqe8TKtjwQU
lzojeK7rbi8xSJBlnJhTAH4kmNaQxBJnZtAQu2cYFwOgPtH9TWkWz2zK3g3SbWhN
pWGy0Zhg88Cgux88mRH1ZY1XduJ9cEz/XOZiHWOBJw5y0buIwrKvZJURa3yHSYYl
I2ktd7vnUVM538GwyybzzpZvQKdceu9mnwfZsibNUbMi0dEoxrsyrFgw/oUyZEP9
o6cHFPvSFZ2lcDEm91xad28Klrg3EP2ShWmYoSiua8zvXG7P2peA4vTy6uIVq0Fr
0UkxK85wida1g0rS/jLl/r1LnfnPu231zqjJC1F5kw/goAfB6pI0oARoWXO+J8tr
AIGsMt1ioFsZdUcl/OI71lGZqZWiBYt6kbQdOLFPHO1DJ5ZnCeXZLTS+cOxhcHQd
0dMdi2DlNleEuKYCYXGumdJuL1SU7jQ4mw07xSyFr2RkoN1j6lZk3vXEmiV2dfbm
i0exP3IEeullKS6RbWzf5s/N6O6xfeXIrslfNCUmQWLJ1Z7g6iw6Jgqwn2Tt/BQn
HCko+8Fvc5ZNUG2N6KkkVwMmmvzbOYLicqv4CXJfl7LqmI21CqFPMZEB4w/plPQZ
5b9vDrHx5pbZSGxgM1t941pIR3bQSRRECQ8ethg13F/99kMLWLmfIC59Ukg4ZBTT
YbqR7hb60CTtOJFiyqEZyF+JqmLTvZ63AusCkcxaY9wxnBD8zBNunF8Zaisc1Qms
eFh32ZVFhPMUF8VMYmGQMoLCTjrmwCMQ6FUAB6t9Tg5s+DmTL/L3hDxzHe0OsFyQ
uQlDOuLx/HgITUK6faj5YEKfz+GHn9ACvvbiRDhNmf21slTwTn/7gs1YQZHuO61H
Y7yF6lc7xbNrwYCJ9J8mr/JmQRL3lvdme3ch08sweImrYDYghQCzT9learPb3e3l
ETCOSJ2p4bYNZnB/PjCI1oLBZ4k8ZOMRsvvnvtwCoRlzT0ymeLb4QTWX6Wgdf1As
HsPVlJMFiJ6vstfGcmCkfQTTDenC4y2AVKswVWlyo7jT2DdOwIR1jVQ3BYgVMnuP
l7MPUjtObylLcVtG1wFJir1sLw1WOjiPpfEaNxD9e4lOcLNuiOOV1E8/UODw/ebe
OZePqddITYDAZK6fJIALQTC+HyEHXk4hCipG+j1F6rn1Psgfrsg/Px4QhXEsOISu
JD+FvVTPFKJMUtpa50i6Fcz1N51XeAAhDBt9bqJSlwTi9YgAAit2qTOOTG6FLSrV
/bC8nQgqDJ1CP+zGEoARMt5Yb9t1gs4oA6bBEMtd7+UVL9gjHyHdVqh/HoLDzzzk
DeDUtsM255exZcKm/sPlU7CDoT+LycJt1X3NrJP43rIAJjShOxiA028nyyw0hk2R
ik4c3UfJ/W7SRbhQjtKo50HXSd4YXmwL1bS/icIZHhW6CBuSlzN9UEjwNkDQH9YY
5cHGtI0fX7f5bTOdG6ze6ENeiaKXMyR/11FVaCw67oAvKdzVoMQQ//FYHEAnRKMG
rrHcMo4REX4DlqkkeS9epRMrlmHAkZc2H3S7IDPITEyV+xhGaNO4sJsjDNdYnveA
kiyf1nxRNsaHWZBby04tmVF3wclxKXKDhmKfjPSJZaTR/ESTOanPm/aNHfSeLrmL
XjUpoae7ZSgU0YCeYmqS8qQ2YCa/K1MfpdIUR8Ya5IldQJotCy9Rge/pGvWFnZCW
yfGb41P9m0P2idqMBt8qAN43jRzWf4EQmZhbT/lO6pp3DsWqaaPqvf9A95HKHUvb
QbLIMrk3OnkKu0EeF/iS/Gw0GGutYTWoQrKvIdrqipsNPKVOievD09IyJIUhJ4YG
76l1T7sMQDECWkNLiwkYN3dUh5MZLA6mz+moYlKTxcVN874j2sYltTR9G1HJL3FN
bT9h9mHH8TCykCPnK1YDvPUM1UD5g23+pnFSJLpDBXI1kUJS3xzqTvhvKja5rBig
GwzbCX6qR166C8031Yz13/HM1DAbBSJvcs51jupNBLnqxVf0qwsFMZ8FNGxOkx6y
bd3Zgr3+s9gUYK171uf128Vv2MFtHJnqs0mRJLyHcQBa7MG+3WnGHxk3nPWVxGMX
IyVi4/IELX2Vtayzd5A1FvE8EKmaFYkLUCpBouHr0TPl+wpl9FGKUA/OYs0poPtL
iTmMHncyu3R8NvQuAhuuzmHTfi5zcGoBw+fICqgQgDCgsKWE/oLdep3S4+JJCTJq
Ra/FOK12l4SwxGXx2tXHMRq2ldIVlb5cIntxhSMuZ2Fc+BVkn6oUW739/atEIuSD
OmvD3fel8mRLipGZkKP6xRBiynW14ovsOlHMCCztXFW6Gzf/+zdO/IVZMlGNIRQ4
TBXtYGUPfUQHSHmfXBdbNBajHvM/CWMj747J6WXmZh1+ifQOhY4Ftckcl2dh3+zw
S7V5RkqsUW8HyUkw/OWYebyXENE7ESM1M+4GqjWbg1RR8Qsj+JUjG1ffrkpcbOLn
ECZQck1atLITo1xnLZe3Tcg3D21pJIxrOBpaC0/7gYWzuPMVxjYupgv1a5eWPuhd
u7lB/m7DL/qbMZPCpE/k1mAlTovSLrIv2tS5dPg01UWj1wN7J51VFOKBDI+UGQ/O
9g2hlEIbaqLZNyN/FDh0yBCqZaWwDE5td7KjXk1tbWrDLCM0ndiK45Ep6gZbmpg0
do/BzIiKX7ILgQ3NiFbyR1odugrytmfzvlUGGDahZrMdnp9BOgelqgYIO7jDztLo
kRM4wMPKObMP/O3OE111gASU8ypznFPmBHQuO+wyvCSSYUFToxHvZyVnaQgqebwN
kfCW1e7bXHCy+BhACk+RO+ohUe33fgG40EBxdgWxMOSgzcBh7v0X+6WRKmveq/d/
ps3UXjbxB/zvHqeiXTt4fDzOMR2tQipUrR1abw9ZZMiGh+su099sjbYoQR8xSiAV
yoBcDXmMNVSAejzcguwAmWfXjb2PEmzJPGN+z44mmGchv8g1sqh0bDLhT6b4DJZu
YZ3uNmlDj64zJBGR1R48KAhYhROw0D4FpFhEq1qceME1TmY1ow6arNSZm/y/G54K
R5gJsUyCOas8Jh2wX3Dgn2hXZApvQDsqoIgKv4xgfXjDVMpmydy5HzAzYrcJODFA
uCQKu13VSSAOugicgJkUwzrh2TjM715IG5M2NuoRTO+rBl/BMFYJj1lX6IdcYLwT
Ij7LKpEKG7xkRmLpL7KTsPfc0MmTp2B20DcJabTXAHEVozqCcT2HUN1GS5Z2sxYH
tH0DBkqIDF0S/j2G3MY9EvamBV4qPC8XeJL9JM0ZZx/C29prHIaDc+0fWXKDTy65
/wEQs58QDPMnv9v4XERsWPTBzeL1a586SqaGj8Au//hfh2Be/uWxlS0Emy3+Rd0u
k9mFnMQ9DII2OCPdG1v0RieLNSAVSFizfRyFaSsf/s8bef/OYJVGNv4/7hs6SHr1
qLs9ixFDNnAC6IKL7ECeZ7rlAbtBESQsRRromDLqRTda4ftFNy6/8tFgabyvtQvd
KosF12ZKSHLZVUjxQc/W0yNGTO6POTJJR0jcKMcVMv43A5umCU7KkVq5Zky+k8FW
ZqI7o3iwkE3QJKwcSUwBiTKFFrOFGshpq2vOrRn3J6iuPYN4vUFlXgYVjPVIT0Z2
nK+9YbgjupMA5srM8HcK6sm6ZpvbR9Wf3nMRFoZGAehjk6KY1iGgdyuaZkWwkCbk
nADmqEcBPzSmonRGZ9lx1Px7Ej/Jyq7WevD87+CLv8Aei8TqxQzHppE4ZI/9e/v3
Z/R8Oloz78YMiyjJIYPgS1Yk1zqb9u0VSaCX5maqqrgIHoK5vVZ/RnoV7/f7Fdlg
9xha19OVTsyrf/IRraGeiy0xqszqJJMm/P1OVd/r6ni6q8f7lbwM6D3QD9ONg4qS
TVcteuAYU0W2kIXE7qph16v+wDTEWM2R4n9TWHYdr3d6i8YJx0xaYEWQYhILs/8p
dHHW9JIFgjd5oMhMSKoDDmxg6oXP3CBohrardyFzGbbbK2CZuLyrFHDJg0cjrLQd
/sB87R/KEj1MCdKVkrBbNHIw0umyshe7NlWC8+rgNqONoDBiu9bN2Z2EHx1xY5xR
pWMkm1yPBDKiN+AeFsTyk8ycRczaw/lsiGY+Sp+q0hd22DBXZYhHdBEIFH/KGcjp
3z7tqVlxnNX+2JDdUbo+XnW2r/IHl2UKwBLI8JJxx20S/TBRbPZf03DOKgf4+C2W
aDgqQxnbeClNQixn92xwzoURmaFHYlNj80xar3gLf3dzMZXWG1C1tzrCjplEjZ5u
lVlLSQb3+Z07BoAlR805yYDBjTXgGl1X2mmdFPyJUnz9kpnnu6w7qaR4wf5WxE+N
S+IinrETo12ptJQoOYqebGF5D7A3NIv2+3UunFhEKgxM1s7/1Uk2WVp/fguKItlp
/aOj3UIzDI9Xsu4Cs1SDToty0XQY+D7TS+ijW4bNAwAi6XWIMeGHlFt9kDu/xSnC
zzU+XfGYBC6c0Zm3ZY/3LKZtjrLEBiHDCM5LS2n0g35+uzZekw1s5zWyYHPqAQHA
qoI+ZaAJqpp8yFgNgUZsLNc9aG7toS2sCF9RLyQA1HThXCygHJz2TfQJzd6glH4I
UDqdqVtjyVnLQ/yBmtgeND/BGs/rclGWrDcR41PTJ4yI1xcvXPNlal0GJTl7p4j2
+BxvuCz7aHiSl4OXANW6F66n3tdULTsvs5ROq9FzCEMpByu55DSItlJ4JyneyII0
tAMrVQan93h95ijV0R1hbDaSFGiI+FETNo4+rWpqVDU3rogTfsGkglsRT92kY3Jn
lc+7G+6vyB/NSKwMupfJTkR25JzAMujZVBsUk+RMV+/IVLqdCG1SabfrVeWCPCvz
AFaiTu7hWA60EB5CE1mnBEmRS81wd2EqmQxojy/elHQiaDn89yZzbzkB38BWYBmF
76JZ4IcANir72rso7lHQuwwC6RtLSUYmuDjX0acj5Eipk4VAtz2OxS1OQqLnkg4o
qPlM5o+E0d7B4w7haogsRV3DuIE6RsKoM27023F6b/yzrml5/I1pzyzpIS2vMgDA
qQpqHcLNQ4s5kuW94vQeKfRARMCjPqw5YNg6QuWK3s29GeSu+/jI7V9f06pWpQ+B
UTPKJFTx1hq/SKSn+ajTx934ZbFgDk/B9oDbk+dojHHOtQZFG1rMmu6ytp+yceZn
JJc5/Ec4YpxiXNUpr7M6TypsjtgfaK99Q4NCzZ03Arcnh/Js4d8xtYPcAMEbzWpX
ZMYvTw9oeCD43eDfzMiyxkkUVdrFoNar44/Uq7Bav56rD0qQQqfcu3E3n/acCL6p
PU3gSFag28M/FTqKmUh+ZxXOSATXOr3IQFBM08NFTKamZyMonO6Nlf8xpEqXPcMb
3YvVx4pxicL/8PTX5QGs0cjnHHhy7Ad6vVed/ueUQ4ox+EV81LNXNzK5gruvdf6K
eC9Eu51deponnCoaACkUyzSjIkLHFuIdjqZidIMT+a/MFvuH6S3JiZUBJWwi1vUP
zw4lcZS0XzpyLOTlnpk5f5s4H/v1fkre+tLxOWADpmPvFTejg21rMhkbQ9Z9qU2+
qSYuj4UvbCwm+W4vjDDgEM9m6frCh1nw+G/wKITUeQBInemDfLNG6fN8Z1JNduTV
lMec4uHB79WmjElC2mO6GJqcR4iqpDlomIlw6nfS18WYTTr9Rn9F4g83fM/fm71t
B/YQbXqE0OOZykfexsRyhkBupVT5j90kltqIsEYKqRIJL/AgkWK5eMi9SqASqBFV
ylF/XuaHoG+THY77AYUZWQwrfqIrCLd/zGhvq37JTJQTU7I5kco3ssNqgG7V/J3J
Jz4+ydtcKiKjBaOIrjDUAC7mZHeJF2NG7AC9Z4oBSLINtVjvujAwglgYnaMWdqso
rcoqrbVnKSQbhzDCgfC6gBwzBFuQK0TAssEUYpxdGKNwVd6FULBCYCHWnkhsJBQv
skx+FZFl0G18USFmuhIR5h2y8T7tbep6FI0bdcmbEkh2rtMH3tue73E5rmdlmWdt
wEVEj/HjvISY0HE0M9YooYdfFEJVUAxrEYXpKenk+eeSww3ZGMB9a11Cx8xO0b1U
UUP0eK74n2g5RA7soDs/s+QMV4JtopitoZTh+O0LlttX53FnKe2gm6L5wWfFTlRR
LukjeFb5zncq9ZRxXlAShFC0uCCc1dg8WS2blOjKToomtDPyHA4284Mv2T+JsnLn
xxLSA8q5lgy2QwtkgoLBN0cn3tKgmRsF+py65m0j1Z9o13S5XYgIu11HNuOhS5rF
tvO1NDKpAJLO3cJwtTVcyoWRGTbB8zWzZdGb4eCofM+SGGMDy53BEbcL15zbLxmk
MpIVgh0K8FC9G23kQTIky+RRnhjjJGvqhLEYe+6X9uhHqCA3H/0APrpGf6BIMjiQ
dYaWYpGhp4BxYVJ9oWYTu/lc9E6WltNMYqXg0UcyvpqNY8XmY8G+jppLCCwNFYU4
lNZjDxbpId6yL/bWYjvaa1RkCA8z2nHtQZ6r8iJzy7R4fAPdvdW7hJHyZDfwH01F
EwDZDL9ho0+AD5JuSq3YjFYH/7VOFXjdZPVbmvRno36kO4Uwl4xsXHI9astz9cLH
wiPQMTHAAkH5hLmLS9J/ccBC7/UW8pUScndEG7y5E9tNj851MEm2Y81l0CHlL/xp
754AmlUwd+I05ozhtTnUK2Jm6FKpRvKUEIfE/uZPoAJIjT5Rq8dyHvEYiw0CV8Cl
R0OWpbgNZyWpeLDsJgrKB9V35qeF9+6SVgPbsHNkv8pMewr+vm2BEnBH1sIf87Gj
X+mYkMXZoB3PMqyWklc7XPmePtVBvcTgsObTadIE5BfbZFXGRy2KPpO1cpLMSMXN
/mg+pjXkj6mYc5mqb2zxQf7dyvWJiKxQE01iz/VB6HNIQD3i9Y39jbnNKLiDcA7T
vFbLW+Hfdz4kLxzJg9LTNyDX3zj2tjQEKO9j7xffiNXmZ8Q9wtxLDixynNH75+nD
heziex0sWEOdDsWqIww5n52dZEl/8VJqmnshQfMj6NUcemavanquO2epRp/dcDJO
bl+50ayj/OhDtNRZdjTyjSAoc8R5PbTULXrMHs4Iv403x+X6HveLhe5ggyiQFNiG
GwjsswUXnZG5fcbdG3uui7ihefnLgfYn52ii0Hs1DdJJWNp5Sjj9+zGydT3PVSt4
YnTqrXn+9X4OM1+Q/DiAh/C+gN5d6HM5SEjdxo4znFNvKCEYqP77mMYUCyWLL3VV
uxk7c50i2HeVuU8+asBMhZ6vm1OZxoDrP8oDkOHRU+oA9IRNuRnMYqp9QXFIgafY
R0RNiw9icI3+PW99ArstWqjBlk8ScPqCFT40PYjW+Yv6pS3f/LU8TTZIZrEDz4z4
MnsRq+8fVGULyQp5Mqzk7yQIlwozraCF+SZa6cikciE+4ZfzmqxqQ050UF4ul5KE
8IERfG8bP98THDzVdErfVNKEHIU8smL/sfMnUE96jx9wcf+0jPXyQ70ATQT/L9d9
DCv0G2I78AReDtGOG0E40+VRQrnThSJyX/FB2O7K1qZWctcs/d/fnWB4aEDOdfwM
f8HZo3GYdqPuW+dZMPYOS4rHKj4R1BKxadYOKR1TanwyTfbc1w6IZPAi6yrEqxNr
6WwR5a7RUsqu6L+is3iYQM2of+tA2oESisebnmX3I3lgmWFEwDORPZu9sDnQKSK/
Rh3L1S+X4Quqyoq1k7xAjokZwBsqcuVw5xtSgo4qRY8Jwb+GYEJeFt6CQt68UoZE
aDm0xmRLdzv09Obv0g9VZUTdu7SLmQnbtTXiX7gbsTH324LxlYnA+VH0d2lJcmQL
RCmVycEfVPzT+70VguStb5+TaE8/MRU78rZW/gFSc2t1OyJZTWtlN7nHmoIapxvR
ecTwWfq/aJml7MO/zbVKGnZrlCCGVWziRqy/d2B51hgZcusFkM420JHR+iOl0Fz4
rI81JsOqta4wEzBa7NMuRrFyOd5kBb9Pzn/lTqB1DTBEFCmSWeexS/bT6u6JlDg1
VGcTr7Vr+umKuA3aKvfS17JPWCOB4aUWoYzfUl3CuLqkDgxizVjQA17I0RSuJaJR
73kB7+ytIkR3KpjglC+EkwLfFzhtZImFS5SIvVqSSraoyX8VOTE/5tKCCJO+cTl0
l9O7WL7+JIQbWp6MsVB9q6L4X3//p5JkcUZk0Z+tajkqr+wgUlP8urbEtehXlPZs
wveru+zN+SQe6FV5fHVlnBcAO+PvUe4b+fCnS8Tu6t+HKTi2pXJwD3hSkrd6d4Qv
MjlsMj49UFNqjRKcOAJZGHrA26Ji5cysgHIrKGdu9bhhuSXp+y7URTKKrdOnHJjX
5qv/PQPEFv6OD39dpCKBOKlbcYeiN0wAMsBPhGUDIOmGltQKPsJKFOV8qH2JEAhE
c2ydjrNrjIpl8lvVGX5328E0j1FShmJ5zCDVu7iLK3b5FyyfgH38CHJFwoiJyQ3C
Nuvj+yKecBl4BunajPu3519FFUSzzfMs5uEKwrPUiH2+fM5FQUw3iJLrc3vD7s3e
M6oLpUqbwb5QrYzVFLljZYti4l6N9NV12btLEt34C9rXh4nyh2UugAw9n830RDaW
975Rc/dzCK01PPHFfDYemiDyP59CfM6b4bif8nvijIPhTbebmGRezp/R3CynadZE
fc7hYk3I8WGRSDvhGLlhRujX0T8+4QpSf42XllNqSvPNhHXLHyoJmR3zxbePLsId
zU7f8XKUJxwqZIofzmP2zoDLLgXgb/OuJcaj5D7MDnldB8kdo7QatRC28bMdIUVZ
P0qjUc0HIIVlQ+X3GzTfKurZQCMYFcofIEO4+ZvQiS1O7l7l75kDlNmS6zqZG64o
4ODFs36LlPe7XBelXKQQB0oohdKi0hQveP/3cYQDTOMTCFIPvadPymF3Cdy0Hzv/
JHKL1vjvkKymHJb41gosfIA1oQAmFWTStyk8Vq2Etxn0H5kKl8M5vptTYZCJCtXm
nddjdH+4YCeUgMk82mF+v8VSTg6afvwvUG+9iZVlxkFe2d3EtSXKhj6UPdP1tGAi
elE2lBYQLLu6m7JGlPhHOPL/2aYIW39uduFjReHU9GpIch9fxcTLyckfv9m7wS0f
2xXoP6PZu9+Q6uorzMfx148fjABm7DX0TopkN/bO0oM/autbXp75HvOkFX2XC911
ogH61Ppy+ExByu7uVj/moO1ZuCBLAIm2vFxMgPN0PdjJS0UlQXc7xG3ffDuqSpqu
iOufW4izmq3j1aboftb+Xbc+rpwIsPMvF0M1fNYPJLIdjfv/MK5vGiQXsAkUZHIf
RSzFkQx9KY9Ooi0irGfa8FC9u7TCokxAmkfET64cq18/3RUEk4CS67tXY7Xnet7z
qJuaOojSg5WSQNKEFXP/snesuqZEhELcwONYQv2Jlkmy4Qx5z4Cf9wJu7iL6VWmg
I4ppYN+ekRTYGrwxTniEb2SQ0A+5V/E2DRd2Fgff3wMcJ/tv71IkbgE52/MBiBxj
1XioXUYeSzvbcN399xrH9PTpsduOO+n2uwDsrSe9S6L73UUqsF5Hz4IkE5lFL6+R
r8cf9UnTYk8bJYnPz2H757L/6Bi87JckbXLB06kVtR6+vHorw/nkRqXMg9IqRnY3
cfUWxGNkFKK+oHv8w5EPOGhR6F+hiauUJflTEWhSa2ziKhpxUNv+OIPCDw0UqprA
lN4kn7D/vpJrf738pOKcjoFKwz7ZCSC6nc03a29UGzTao1RcAgYySvvQZG7dQXgQ
QI3ZoIjW2UNTKuU3kNrMZK4zQtYwGt1b4VHrSZIN7cwvyBf4U9emuGMqkfplRP5H
HHDx39BGYuCf3gRxGWaxUJO3HCvjPWfwMg8CnKK311ikJdttUDKVEcSX4JpHuiL0
8GhKKLYz+YBg5OZZMUk2L7TwjAM71EisTL8sWibS9rygNEbMfuZiRo0Rq8XOFAsn
gYSSXrqoiNw44tsxBKW2X5m/S6wd2OJ5qu/MqC+w2fm+O1Tntstkd4FnfPzrf4hh
e4ZWkUsgwgPCVfnfcoDl9E1TcS3x6vslenWwkRWNGetAgcTG9BXjMyK4YaiycITp
xna8dbLEfd0WRPpWCqAamzFxnlj/fhu+LYhs9ImQcHZKUF2Xp5qg4L5wyR93nevf
akbRi+BmKCAzBy+tokPbZvnL01dy7BQ8nSqILtUDm5AA9blVTaQ9DMOoVvt7pirb
7hmeXl1OfoXVIjlJpBNKyPQyuK92Q1xpcniss6QnPBwEJC2TWICAaNK1jN0XlTdH
UV8dhqYOJFOBVvc+NQlv6eG1fCRnhid7or6p0qmfvrZPi/XVDzG3YDhVsnF3CcLQ
ibvJrTafcibP/8jLcvax+PAFlX1ng3FN3A/A8Q4/OVjo5J/kP6Hm7zpj+O5yMGFj
0dSXLhJ/p/LdC3aztAwql3nwVWc4wfDos8CrDBH8b1ZozxCZ+UeyX26EJRurUYAQ
dY5/V6VBY/7esZz21s/17J0jHWLGCRQgnN/UqrTPrul1Mzc6CbaAVe+8R0BIi0qi
bJPNyGbuSPoBZijFOIEDSWtHQO7EFe4Z+GNvFb1JoXW4Bd8KqJYxCEQw6dFHNH+o
trmngDckwzGiTVJCJDKko6lKJxBosw4LT39SNwsnHhDElSwDUxTgpmyTZOc5D2uf
N3LT+jlH6+fj5l861NnxxqvtbuEWVU67tsTP804dyjNgOe1Hqdhmk+xlf6dCqL3w
3AgKGvi66Mael32FPfEhRgxk8Nz1qx7pji8LPffaoo1xgzjp2e24rhwXM0BOd8BX
bT+CuZ3JWlfZmtZMsAlbUpOwy4SDNxf7tsYalVxhQVdghtwtc/neQv2CRbUwnPlD
j41TJNs6BPIJRK/OBKXzW+MZxuRoWKigKcb6Wnsrn26EY9mQ0+RiXWGJbUXRWr5I
TDzv6uI4M5LjJv1UgO5rK4IxAXrB97rRqs5FONrz/idgGn7hUWkmJ7BKemd/7LQF
tiJN6XpayyieqEOVWBAzyH0IxzDEjyYmq3UdKFzd66l5Qsiy2hnYDfzA2/Tsl8xb
PxxgCGx98iN53BrRelOgzPQ9xJSaU2R0HQZl0GC9nFcSuoE2Ps/QQ662Ml5FWpLh
ggOd+Jf6HE503l/hV9accGWwbyVeuZguelyEnq2fwPqa2ZrJAdkcNS1P+0f5LrjP
ZsZhh80ylMfsqOmzyvhL1JXeuXUJl1PHXavQt3lO10qPLGN9Vh+cfJlTxZwO1xSG
W06z3tBuJUCRmW7CAnjho6EAEZzmozfiiXq2NM+CaxYlA7B7AAyPPaIuucP38wkI
OkM4E+DCJSQ94Oaob7VRG9ixuO91GbzUuMK33fj4IxMQregr8+u+lRCAByqogGZi
OMpsvpsE+xr5yoH99AcYmumPTb9vvMm1jUuL1VFktDrmhDi2uWW5MULyoINMcSLM
fKVTMFKtFKE8Uj0J7I2pXEMqDAvJZGc6GA0N+Kq1ZhfrI/AA3gl0IguOXSQOuFLr
0AGHje+3zOFtpNE4gvpl+Kanm3cUUjp/9p1CbH7gLr2UjuQukh/qW4cFVqzxdJHA
XmAsBLm8Gw3tdMmHwVlux8ql06Zv+EkbrePf09D9je/05OI4dlwn+ZH4cBSPamja
2WMJzMRr2UYGKUm/m+xbD/sg36YSezRRqKxZBjOj4BUFhoJjJYc9ACf6BIhC2bT+
zLJTq+A1WWp9zPOmB7elGvj7x5xqTdG1zRW64V7UgdH9OXXuqiSw5CKX4Jmk7SAP
1078R0F2BYPIbbVS/6/dm7xJta4va9ZqMqKEO2d9xGS2n44UCsJQ4Gf7ed0E2BuJ
AwZyYRdqngEP5A0wir+eDNTXI8eC0MJ05Ed+FCYQmITowV/nxkFuKYm4qM+9NY0k
09Py3r50nPaNuXvUYOWJKZA0Bpfv/vqMqi/q5Nfb2c5e3vt88PJxI/yMZW+bv1yp
FwNtOUnlHYlkACbxZeNs/4K7IbYlrLJW/zQiem5E1BRUci6EHAgPz0rcl//YBZ/A
bm8RkWz48aGB2qZyoSd98Xf05ynzqqzTLqzMCd6NO5qLfoVChZdolkiWqjHHzd+A
M5SRbj5cSpFB6Ot+f5wX83lkBvylmPFmUVB2tz0n8UjQwZzveIGf+nak/XkX1crU
cqdGaf8woRmWLFkF+0lbWJMSTdcGJrEu1/o3aUDPh2AYJ7qMGbSa3caiiSQM8P7v
nl4oBj2KSNVVVc02CWz+H37+WnU4kuodMFL8w5VkzRpglItBj2a9HNCEJRfiRRDZ
1dlH7CUWtTiRM8TH+YLNSqSiTk16vPiagANYgSawwZ+WcA/nHsDOfSy1WhYa5SRr
JQl7Soocq0I6vrD1lS4kEYsopB1o/HDXx/M6VR3Ox12Aynv8Q8fMHj671eNxgbKL
ilBBY/fMmGnAAIPokGFRtWo9pxrEARIkQxTSK5wnWS1G4ilVx2da8+MshH6Rye1l
rze8IZjo2rU4kePMvV92hwhHPfiYLbwisF5qqhngeV3vfjECy96KOeIf/tseZK1F
9LsERHLXIuyqnQChbxHh4/3SFXB5O/SHEIiXxr+u2UpXR15CHCX6dlLjAvdtcP3N
M+ML+thbdC1uTR/DIJP/C4G8YrmaD09hORWjEC8eJYDjUchQL0N0fYx75HX+B3ys
qK5+g/qq397/pqhNVXqDE7yWBRZtDtzbusxGaTDmlCLHMiJohfI+IEe+/vVeBEZ8
yMTj/DnZ+gIxRJRwhhE+8u43JHyVSnEJql3UEsWI/DFJhGhgqozKsW7i4IW3Jb2Z
LYscC/yXBIdROtkLar/CfJAhL8OGejihnpH//JGjlLX6T59xSNhdw/hFS6aBteNl
aRIaiDb1aMEvVv2w/eOvB6TopOgfKcjIEVvGnFvBgqM/PBHVTEjBmZNmOp1J7XMt
qvqlwjbqYb5elHyaNA81fqOP3fqlFBEhGyuKFxhPXpJRN4hdFuN6eJwLQDm3oDVj
d5wC1VVOMmzH3oiE/sVZDGZW5BIJKi67GSYkiNmgHt3uCASms1Z79z+OUc3b1W9F
aq0xtUnZyYCM80DVTjStKFMWob8mzEa5+U83jydEAUT9/D11DaF9mVpIT0dUBa1m
I1ErnWX8rABsURjIRZip5IYlS2v3To0SOofsiQMVCn/QGYlIhDEzkW7SVLTKY+Sl
mOnEZn5U1J7cYIDRpP3gTV0XVdOLx2annXoq7O1Ceo5w7pZNKWsKkE+rPuOYNrae
Pf0Q0z/53w0wYuAyEGAaM2uBBpKDm+JnLEyNSQK3lq9LdNUBmEcG7oI5JC5UYnId
VfBmyxbJTeNNJGXX7MQoaunudjz6Ci5XrVmNkx/2U4+G8hUSjnBhw9itEPP8WefQ
LXdXKgksCZxKOePJLYByrJORZEYHMdd8IsyrnBkW/W0tdPXlicVgMiVN+EIl/iXB
ROn8ysMH2n6j9sCsQbdBs8vX1Uab/DvirySRqM5u47wkpc6keIGgyQm51ffv9WvE
L66dx9//u9MrBMBSoZG+BJfZj9cVV3Gw40oTn7zZTfit4pon+1vqRdnKXIIgI+1P
mVGdxKFBEj2gTQrIxMLhtCPdmoRVg4fiiMVUChrcEunp7Zbpr3UI/xHaiJcnYZ63
/a2E6DZjwEzQ+zuIQ2Ann2JzBDJxinPb6ZgC2y7MXgJ9q88zk/39eyBExe4OiQCU
I7akqAjP+Dx71mANHfHXDXKtht0tchZT/tbojRyrVMcZwLe2al0SoRdrPNi/Ik+s
RAROnNak5cZ/FkboA3uceFlVZnOckPb79VWpEQKwAZ+FgUpGnKW4ZaUb4IEjdB1z
beWRgr2Pqc1cI+Se0l71U5s6A8YgzMJLE9qdGvaYS2XcY/SmT9Q801M6uC6U4vOB
QVPPU/rKazq3JTE/MGnArhCYhe4BJ2fQB4zmV70zo33A5UB+nhFkzc/ImdiPImc0
M2Z+vWzyuKQomFb9JnS8IgJCQ7/Lq4AxiK1jYZt1PvjWsXV6uzv6RRVTKx3xhNBj
tFXaIHixEruAq1ri8z+Q3wicIThkeWvv2XVB9VQpT7D0I0C/yI6P5Fo8y+ytR0kS
COtaJUY++didUTOa8hUTyS+EWgwky5mVh/HjVWGu/5ZXVWatuabSyC+10Gni53mi
MvYnUSmpehdtgApBlicUUVKEEzq5iHvkSJw+zwV0Vo/DCrpax80ybd/x9i8uDq66
kkuFZ9jCOJ0T4ldVsYRbUsqr6i42V06xEKm5mXywWZy6dGpRlqC7FxREs1CgnTxY
52y0bWWyoOLLolsEeiyWF0NFRVQJ6qa0Vv07+2ChPV6YqiPQQwH8WoobNSeOOXwA
22NtT4Wj8813lMf1hoPVmKAWdqwEwCn9F/8bwU17ZiWGRMOLWMCzZeI7zgdQsWRq
yF0+2eTaVo74ssyTMfPv3N4881g1Ap1snyy2/wBPKS7IJ33c7GAE8wM+eD8MKUy+
NglXYQ17ZcrEC0HzXkPinxxMRE15NBlwnq6d9JPe+2wnogwTlFyHC87oF+GPMMdh
CV/KP+IO++EY+C9Sw6CczDGzR/wqk/Jst+xsaxZpvxcm+xeajP8cqYzceK6w3iPu
8oDF+cshrh4i9pAKy3zmZB7yJwPUeryCkOTuo/k+TNG0+0e/rE8UjVXT7SBzof5+
CgWlZWWR+cyMC9A8LYXq9G9TXnZr9JyeH4mqft82wG8jimlMD4GY4xIQQZKHTdh5
EvsHog+Qkyn3R8q3yekBPiGsMaS+aXpukxmqp/8gnIL9h1ZQ2cmBACNPGLZ0gCqH
t6LEnlhODtrxUJUrF/5OZF85Gix4YRy3tU7i7ZDjL4Ts/WcrSYoQ6Mk3N/EW7wjm
BRG+eRQ046hVSvtZWW9G+pUFD0I5SV7aS2JZx98MQy+NaQlG8GxZmjQQc4WEAv1X
ng85phyrvKm6rprq18O/Q0A7+pYiwitNlp0nI458LUS1RYhROWWicVJ0HT2qa7Ii
0m/gvqCKK/Je2TsFWxs0k2KBxF5F7v1CkhIglh+EVqYaRm1hARNsL029zWNBAfVz
bqnRiWUX8blWl+UCtJHrLqig/axsUlxIG7ZijCaNTsEuScS1m+IjMnpkqhEi+jK9
Z42tXieoJZwGtOLl9KEC1jxeM3rmCYaprOgI4DUoe9qYzCTDr6v/TQDdX0yDR7E0
ATPOQ50Gw9ymAZ7meCYVtxxITsGJCyc5if5hNEQ3tVm1gKhfIadMwehG93gMBPod
pzm3HongFRJL4WBtngj7LLhOFSpEArlvGTlDh5j0yG5KY5Eb1Do9k/Ly4VNpyPmK
/cgGvVLYsYRsKmTLV8KkGs2B5sl1sWuosYDxYY+mt6HzVu+KTyo19RzuaQk6NziV
dXguw+ejS4LL2HEqSsTn2T5ZffbL7rjT9EErVHEcnOyP6h0uFICgVJa5ooSZmCnC
+JDDmxQM1UXEJ/wbIHGRUgQrWeDBUDzOSdaGeBgWIoqEQwJGLEcL4VjZpuO4ro0C
BfT0PILGYME5Ontc+Z/Y+h2PoUqPzWDbJMUKlWpMWbDvbH7TxKdjmD9EJhDsyGA7
o3jFB4y5fKaLcvV81cv1DkXfuVB4eS9kXEyPvfwrQmcW3bGIoiUrg/UpCFZAcITV
5NQUkJfB0B5BznrGzO1Kj48HUZnGAGf2P9oT1X8sAbZk2scliV7c6swr0UvNJyMI
XW8m28DgGYfR/JoDcHgjwukXQRFesTaOjEx1lGZuC0+VnRFcV9F/sfyVAYz/EAsw
POQrViJYoSt1qSvqQZ0eZlrq6jg6NFje0UyEB2wNf2MqMJYBRHH3iCy2Z+wyNnXQ
NuObtUNssw5YIVDyvVgAdOdabua1YN1JrXkC/8/Qk3H4r7oc38yqyJzOVj+t9KE7
XaI41D3bYTPvxqBqd/JklogeersYv2oiA8UHI1MNif3sWAplb8w2BKYDCVFUABFl
q6sEgb0tYzck2nn2Temm2vAku41ZFMEjV9jUcDtinZc019npkhd9zWgfnXc9m6k2
xQzNA9m7rKG5hX9lUSLTnrnOSY0M4iyW7WjOiYzVX0Z2wPmEVXodj+p6cidRkcqa
EQSxBSZV7mVmIsxxZRxjKaawwV/+BLBIJQ4bFmHLzLNkY7z2VupJfCjoxdQcixv/
lMVdpdOunvBZgZKTP5jfcfiBdaHPjeq2oiIY0UYzBKCOeM1y5s52mVBBAYu4Evzt
5DsNN0n1FqxPFSpU/H3wDEOM+7fFjmKQD5bvaFbeD3wZ9MsGWPN6AIXSXE/I8R3m
+K97RPUEYY43UAvR4/rt5mqcMVr/77USGfpW5p8ThvCM5ucrVyxbgIoCCFypp/vf
YajEKkiWuRjnPGSTVIJzBPDDZQlwh1BHoStdpRKHc6KQq1uemXO1mx9JGQIl2xiH
XdIDllv8RkY1w1yAEBvwH6kW2FAkH7Vx/NqYllJJbFCw/wdk5dFfLB1mCsnFoCQ5
C1whbik4/dz8Y/LewqgYs9Mi2L2VxOGWVIpAiX7HJBi5fTyXnwOsdWNY08yzW3mt
1tDC+q9qp6KEbsdbrAiLf3XcWxsrkxHXpLVkVL+QsFrwSKvywoFLrW1nWHePBeZD
b/YeCruMbIBdFnBK97O+R2bp7L2EHuvNcWIQGfANq6CnlmH1Y/neEM7tHmpuG5df
oZUe0jkLQwP73ALCK5qjix9sw5pQOVW/zK0e40ir67xQVZY/mUHpn8Zqiv+h2EwA
aji1EDvMfOriurlBmoiNemwQcYwWg7e0rfVvW1Sq6RTh/kgSyKXx9IOD3q94OzWL
NUAhZpbeBOvNwaOg8xFL4TJndKEfrrxHosB+S5l2z7Eg2Rmhy6MXOpi2czut94ui
z+g8lY8UG3hW6n+r7QbcBwH1bpn9SQsOoZn5py7inJgzxzENNfmLWfCN25ImNptB
Y+gbvDIZ7yRjEl6lZ62BXDyhyU2Hk7I3EBVA03L8jdUrmo0j5WC9Tm/ParPNvB93
LmxxZGjJBTaOhd04PP3/JtehylLhaW/AInFCgekMf+LJST3UKl1fCggUkIJGlJHD
Ywth7jqUIxV0JMGvyguLT5HCZc8mSjx0ESqKpmivqR4JjjOeg0TO2pJcyxxSMvfU
jY/4b3arw6owzcedHR76Xos44ZNoFUEkSKm/rKFP/dcm2+0bEAFrjgoXOqE2Mf3L
rN8CRSPAezcX5LLfYJNGJfq+nTmD/v8MuI+ncr7hK4DQLEs8F0cXrWW727KAopC/
6z518SRwrPuy11P9e226eNOaP2DXU5jkIRoMzuEgBCPS42PZ13QaILMWXEQsf5+b
Clf/h6azcArqEk12NU609S42+iU+6DoydFo3O719kS0kuWr//k9bmlKr4ZMOHxbs
j0qCF+fLzeFgwcqopaBmJxQMonw8UvDQHYJOWh8koXqOohLIwmlfaeeTrHgUMcHd
ab5qju8s60IiIx8Q8XELhfqvNV6qiPwNFQejKGATfOrWGsMQvmqwdy8H46/jpyga
iSUt+yPBHNc1D4P9UsrZe4RSrAg3eDmK5VnTgr0urt6KEoSznzkz8J+x53gbcc6Q
Pl4QDJb0osDsov3JO91P2Yk9hir76tkyDx6SOjVCKfSA5HiLp2/TJ3z3SFvOVxnz
iQ4QjSto9Jz0UikB/balFfTU4YAGzghjui8G+asthEJjNd5LlowruWD1+oKlBb3g
M3Jejh6zIpbEJosHQ3dCRagovL+oiWTJQHsUEuXDvQLellyUr4qY89Qt/Nsn4rdo
3nIukCEtn7rHX/wQt+LZ1s0+5/V9wfg734xjmg2fq5ojpkMu6yUUmAiAtM92R0w5
ZLmo4QjEoH8VMekKvQ91ZSyXO/kKjTI58jczJNSBoLLMFAio0Zu8dAAoRFGM+A8i
5Hv50+V+TtE0VV4P4OocaCiSYsLtUWyexvKgMfSCLI7DykJitbhES68sqgbTGXNO
wqH0pZfDnIPcWjXKCjGvAsFgeaDO/YwdqkiBLMyhLjRFx7jgJsyyIRN4qwBgJKMV
D975YW4geXe+rpmjSVKKGyNEb4TIr0RuQfbMU6eZvPk08eSE1OacZqhY6FOI93AP
KDxoUuL505sXK09fiyvaP1Zm1yD/c1yLdIaDdkUdUWMDlM5OSkyWUZAJXXYsLgSF
3CXDfkV5X1luLg72WzONzbEFd0jhLcjtsG+opffpycPQRZb+I/ISEzGgiOMi3GH4
Pp8sMKN6TQubQE+gvZnhtYddNBIPmFcz+8QCuDavEKPBjqGbwV1kyAm3px206B+C
ge68DYSU5f/AyCeL9LVewlYNCchupO3q6sq6l0EzzcJJQKBoDjaWx2HoFDmB5oeL
7YyoOaRPJ35uEjky5/0Gd59oajXBZYaBFJZ2+hjqkoklG+BE9QxtQYklhpzDk7yA
OCBT7wx/28vCkHrqxtvE+4WmwRKto/ik8V1FvkxKTtD2Udq87RE5KbSMnRYdnX/t
XFzdvUsx+O7LeDgg8k+b23yQ8LKnpQTB8P4Ke5s/sa35G5N6DiPyWYTQVWUiZPN2
bwxXH0nAoP01DbC4ENg6pscW5g/bvWPsBVi0xsLcK+wDoW12/WYFJy23MAQjzmFS
y0MzkSsrGFZhMLtgmUE94cMNoJ9WRKfOHtkY3Z0Brv/HkyU1m02dQPMA/NBXkb5F
rwyZVgn+NCxywrvVhyQVH/zROUqchTa15hdnCDCOO4HxuVMTcKvsGeNrDxyLLwUy
dhUj5YYLRTbs5iufvNscCr3nr6BEFjWTqZ6Mh7uPkxFpQ9DLis6+K/C0Ts5PrrFF
Wq3Iq2Ah5Ensb5nhFThvF7bkEdkSAfKmuIXrLytFLorIAx+Qy/nXHP0ovPfNuI8P
vVFnBdtwhVgpufUgVqUMa/thZ30rGdEVYKUXU0u1BDvDsMf3cW32Axc6sKTZqfio
YoNiNjjRMs9ZCFyFGwcNgVBdqu2AI5cXL2DglI1yi0YNKK1n3dbNU8UbJ1xHZRyn
duTPAs1wPAXly4XWu4LvMLNFORWvPDAd4o4dPAALm9Z7tMsHz5urofD2psss5nBV
naFU6IOghlaRRrjT3B0sTLccGjQ2BrMdDIbj8D29AD4w3U8FhCoXmq/yx02H0J2m
MfX71UQ+VjnnuI2logQGGp6fvugKBAgopz2grJ99rG2jKcsDeaNADEie3+IgJ4Jz
WaHtDg7S9GOmtbd5OjeKCwu8taGxK5eFhzg6xltZrYOfc8AAGCJ6gUe4mN5TXGkc
Kcx0tqYD9OEL/gTUCadLFHjKhlUENNVQtTa5GkFMdi3AhAPE8rL7ErtJtxkbQMxW
oC7JNqyytYDyH3xTgu1WB/gCwul0zUBML8ey8q2jXaafDUzRcTUeaobtxFUGKER7
9KKP+guUSd35/K+hDFKao3KxO0WhYDY6F73Jct9cvoxl/fjw7nkzAi2jElQYbHaM
2njy54UWLSpWHwPzDi7o/iAM07I74kvh9Ud2fquYy3gUBHORKxzSzy0Io3mw3Q1L
/qf409tGFh/yvX8sloifW9b1OgLKMHQR1FsewWUtFGGqxDYVftw/OZKoQdRubyRn
gGZH6HqabU0SednIXCiYl+P58ev5LWtIDC52X2XyO94ZV10rOKnEOT/+AWEJ9f6y
HwSxOw+lhOiwGOiaEDi2Yvg7DbAODfnmYCp+U4eEnNI7FPSQCy3fEWDyB4IDuI3r
YMSLXgZbTFRUvY3PbR6APYF0z31jQ9R7HJl8lyE8+/+gHbox9WRqknc/cVhHtkRy
RWTqNyxORzEw46Kjxssq9Wb3DnCGlCfnwRO/bpcSD8t2rubq3Z8f6xU/NlOnMmW9
zl6ezSuDjmIxYzDdhWP+HfrUBtMpyOdjLPXHk4pGesybGfz3cXNRBG2rcuKnMs7B
85mVP8axVffso5L3fTdA3U5r3itvMJMqOgBQOH+q06U4Ertj2+oUDHD8Cn/IRPyK
/NKS+oZ6jIlkxZBMy0FABdLzqgIvLzOtNNv9sJCGWncoRGGEaqE6Gdogzk1uXHJQ
aCw/IvhKphERPKeGuKboP+t48sV4y5nr5RGqsiNw0CtfO7JaDXDXkq7rS/gp4ofD
Ba0h9MOL3LT5NdnJKecf/d6JZVp1adVsc+v3LN9oCFoiFTP+gZSi074dqEng/oLD
6gQ3cZjoJSQZpHrR5n2yygnwcrE2xhydAzy6EtGPxMgo9e9YHS8soxQ5o/m4IclI
XDyvbgAbqQm/nln8Eop0UW36smWvho+03mGQZYukYccQexx8a0kaVbMvzHQ1XcNX
IXHKgeyzyG7jL9n/3Ag75e+7MKU9O0ACbdk49DE7H1UVhqSXYkNlczqVZdyHYjV9
lhS7CxhUC7ZgL81wI5KMGBV53/Z89sLtxqI1iRgBorxqPBKQvUXbjHPfZvVQc5e0
AAg22zXWZ2akV1hI+wAEHP+Ud6Pb1RpR6Z/XdcvL27iaSh8ThJDBd0KlXq75B/j9
5Ba6U7qhTXBr8/tEoiL77eYMBJxofv4p2jbLmi5ljTQvxgUXF/GrU2XnHxQlB2tO
hQC2qKi+57OXZKgDPYdy1TQa9JZ2d5xRANCNt9ReJc0RRWCP0/l1xlojW2bony7H
qAb+GXRBwO2/8y77GTtiZd0Sn6yTsuSaOQJleYZHrEsdxavqJKvJ+c4cbx/47RHg
zzZD0K4Mk6OUZkScuyNJQGj9ikQ6U2ZT5MJCxYPV3u0fq+7wr9X+d+uYuSDMnRsk
rcmFwl2fx6QGDsqBuptYZFVevwUlwcYS06nH0KlHEtGvuQyXZnYmZ8jwh42EX1Px
ZRi3fSyErYpxsw5gJjgAiiucxD4nsAPnWxTbtfh59mQiQmgzILqiq/berfsJMNS9
t4JmYcdeiCFMoIGYHDF2SevRPmp4NDSx1x/5ZP4Ly3NaisQbpI/sk1mzwrPHatX9
fa6Fps/HAaR9V7tu2kDI/2xuFjaEXIB17/a8iJjwhGxgMrCeJg332aA23nwptjq7
jPMPQHKfFDwwXo0OWhE56BUJDggwcTtf3wM0lqpLUH22gSft1SsRhJbUCIWHGMuq
BWMQqyVhTSa7sQ9UkAg8GdfaAwD3AL2HBqK2xQ8c0pveZt2BhbZH3JhGKvz3QG3l
1pYo4OfZkSgKfzX7FdMzWajWhom0gTD5j78+Fp5P/ZOnPny3CGOjzXNVQydUCTvE
15MMp+RQVjjSybFVp90xQgBc0JRnpoIJdyQhur+AKQIAPojMj3omyIGhPEnj0QqD
9BkLaqT3dKptc4ATsgPeaJJoFpLhrS8buEXu25tWTo5VHRsImnfaeniJPsG1YwJM
wKr3BtWfkGEe33bpoZXMrC4OvIe0ewkH/TN05/uvezWDTo1sEgikfMQa98G61aOc
vfHbT9lHD1dIoPcfLewUhN0JejE9YCMhPkEE+3AHO+i4km4upDJd2lrLo39+dU31
eNBzWIk0Kul6/7N0AbB9Jr9sWChT8NDYyvFU/Tx79svxvRShlA14tQ5ptKJ18EIX
fApb12hZFw8ibCnzx1dFRJXrQ07U2EPdAPIo3dlNHsaLUsmtHh+YZiO1sowcmvNG
+lvxufQ+J1OSEQhFvZ/MHzt19Wf66ZoWL9XxQpHjtHTizvuJUwxMPWY26VhwKxng
OEmDuUomntbUYTP9HTB4mAMhPbeRn9burEB4dhGIeppgPxQexgFhlMr0KZ/GPAGX
CtlbAWJjuxmCpCuuapzcP665gvY923O7S4iHyTYKX7w/Yhf97FinBXKiUnqpSv1S
mpghTs6jxaKuWR0qDpCkqybEJyhyukT1qTqB5roRQh3z46KUxZPTl6dAso4jAFya
FKC2ccnk3Vg+vrr1KefyM6aYF+TekAZbt1VGZlpYjtJVDCMXTxZ+0Zi3XPOk1xlA
S7u5m72+9fqzH03YPHx/rLvyPrsaVhPFAy04+Y28VItILK5rsy5QxOkF/0bJs937
1wbK5V2e/GWUhQ901fowOvCnfOMjzBPZk13vidOfCidgmBcuzGHS3ID4OrnnjoSn
XKVSauB/uykSMx1lMzdEZOCcJHtu/4io2Xjjbd0Yg43BK8+5tKJzoJDrUoyA7EsS
GRoBUS6igSbmHJcsx+FEC3CRuyUTUPS2prjinVdhjiHKWIhBL/JXKEgK7Ejho7pO
W5oPpXIJ/A0B7jnUneDGX4fnnBZvD4nkg2e9MNMcly97la9+DvjrktifR1Nl33pJ
b6ohp4avuOOXk8DBYKAu63nXC5k54ZzqPZJjPHd+EfVay7TSMkpjKirHvvXvYvLr
R0WjdO+RMvF8jhZVs21GY+RbOri5RppaSz6+vzwEwL0FDaN3LIqQOloI0pfhpspz
GD5b0B23ZNSiWpkPgAyM14AnQHLdHTxrC2otI3ke8Y4QCQV3ONADHs+dyeYF8dqL
Xk6+7Iw9NnX9gaQx2+1AO97Amz59YKdxgQudwbKRSitA4lf1vGqwlfNk5nAIXg+v
SVU9gyLXrDUi/E/nrxtQiUUFOiLukth72b0VGMPbfh6yzHt7EjmLT/jN0OZaPl/g
bROb6XYDyxi57TMKuN5Ct4FMH/RUg7Q4wxvobATRI8MZ6Yc35i29Y6LJFTxr7PfK
rTCgUmV2QLVYVvXk+dlJZMF8SeIcQb+38Qa26EjBWnqyak7cnFeOfSmI0rD0qQ3z
ET0r5esj5ti09AoPgknO0NMeK+WWYTwW96XNDF/GJek4heTKbi+lFF0mU67DyOzy
dM2b4HXkUvddJY+331Na//fWr2BqxeO96psmqvgCtpPJnTN7iXs2y5W4SRSCCC6Z
RG5cuwZH+HkA9P2TqYOB7+0tlmOGSKeqqz65ry0yIjPAyYvkD960lsw62wA95Tah
VDhiy9cKohNHk3QTPK5J7nAPWdU4DsEk/+3UQe6MarUH5fKEdc4JQUA7yOLfHOW2
mt1NzVaPz2TBeGL4quIKFbYk5h84a8WDsatP6BSDTT1+noE5qcrHoR+OaEm99Yg9
USVnWhDZJjnruh03OJPDzCbszPnbpEbK01PLIL0kXFe6xUUKIrVtENk6f52Ob1Hj
WtE0N/PJg/XSj5DOvbGcjFb9Ow/42zq7nXgJsAHqx3fOKeOVU4oM4cw6uferPuvX
hHGrdZWXTrrlNTFlfE19j9WQrRJF/TReb63JNZGtycGGTyQtFgI426qyuaAW/jXR
w5xjvmGjzkhoSHfcgT78eo7ZUeABbUBkqnrjn9jAk91cS1dgD+1CcWnOKU0M6lCp
cpMQiNwmDEBJktbnRVURT62fdy3MLVgtxzBYE3KKuy0MZl63nhznTrGeZO+1Mmox
p/+LTheHyYMpz/Jsx4re65jQXkrMA/0xXqYYeDxOFiMShiqb5BDE/9i5jAW8sFCz
+EjQVW+VYCuUPGMIFw2dHzvzHjMNZPXpSFYrvKJuy4mpfZiN0Z8bTsMqpMm2zoCc
IgFAkCWmc8sGNTovxRtcKm15FSmWopjztRCVl575fmtQ5fdOZFaI9nN6HkKlRxYc
pyk6BUlvbIfd7qqTM5EQrWetHflmaSXSnScN47SwVshAYm7TQsw0S0nJG2ljfM1A
OtoYPzCz/gv5Ar+xrWJTKtkVEfSQ3sIO6rPQ/t8ZsD1G5s2V71Ngs2Ep6By8gBPg
s/+H8jpzNKl4lbl/fbZrV0K70ypvoYJ0xeeU15WyHyizgI3e5HN911KURT9U73XP
1/SwPpQUejmcv9lzfwU8On2xbq9CyGTYJzlNYH8ytTXVTV7l0dsCscsWcwDWL/ls
x1YTuZa2v0dOHz4eD9+otF8Qfn1OaUOKU2Smot/wXa5alVBUqFsmu5GbmGEua8ZZ
DVxrbjgYlUItsTO86ufD63UYInIopirYuAX53kLaZ5uHILYsoHzByE21lkhh7XTC
Z4j5qTmodCm6fSmyPcvL1l7XS6/N6BxzrRZi66CRdbS4DZZPrFaJQD3PPj7cdwMf
/Lg4VMaNUnRq/dexNj/QhYheSL6yEOGkMmaUfVjHb9O9U0Ur18CpabRO2fA/tp2S
doqC8YDKzouIzOP4ZuakUX54vViA4XSLTe2EA/TmLxPFKfRUi22cl8cwL2OR00mU
wUd8pxS0AeRqzw1x6+403Hq1cCgQx5TgFZcsceollsVVy6qYDzAVXq3vACNtpp1w
h6VtIzCQAeiqWHNHa6hTj44AtygwZwCRYABt/UX/CNL/HsEE0feeN5GwabQxdg/G
YvKZfVt63ZV+c4MHR9i6PFglFDoUNOhces27wRr9//cRWV6t2x9RzbnXFBLUr4V/
l3jXm1KgkCbjegOKovUhboo425boBp+Y+OPknRpzlTNSCzB0onek6EmSr6KRVoSC
jzXAsHES1Y5paeRpuyEUsPDumn9/K9uHY88+9t4OvHkklg2CmSb6LKhsffa1Yr6e
Co61lEcdLPU2ehLuQIRhpdPIaUEHukCr+s6HBjOy8iPWQpJ4IbmWHRKqc5eN5VUE
OEoLgXxze5fNv8g52SGFFHHzHBkg+2I3E8CpGa9Wg0FsPPWXuwbA+1hnu/Blag7G
eHXLQXW05upnhD9m31XMlxC9U2La49n+KaFRO6VAtXZJX5kTdk1IS2trwrhreyFN
l7HjLvX0XwXyTjL7WG9hdv6RNIa5bfj4C/equV6grPZ88e9EhH9qIbNHhKPh+IXk
gtw80/DvzeZd5+95IRZhlEf1D3j03N8BcBhooy2OtaWBIYK2CMRSBAs6yS1shJwL
4P+qkxeJ+oJ+EKbIw7lA8q9MYdJpci69bM2HvCCud3qkMzRIM+NH3hQC+om4rgcO
D4FyHfvQ9VIF3UoOkt08jJpi7nXfK/rV6xrWLbGejBUOYRX5QTpXt0rBPycgBE58
gakBSS6x/05lmjU2mkIfJKtshd5kc3MquN3R8a9lT3q2XHw89P3V17eeNi9H58nc
8Zzs5NOATEBQPzdfH9zhjU+oo9KMOb1b4PyhcG9xhkpi4WJqe+YICyV/KzWagt1p
hxEKupVTpjVh0gURhlc/Bn4KAF0WDgOwpL6SNQ07BaZiE3jhoVRskpP32t1g6H93
DKWmb7A90Kky9WOJSf6VZgES1lkrNnQ0IQhX2tVkYbZEIpK/IfCaHKOfbbG9vLGN
REySggrjz9pNYXHbMnR5ULt3sF3Csuax3EQUlHEZ4MoOgSzKAc9IogA3o49O6haR
oxo7WGGxEMXOvAHKIA2jqa6oMj5SQ4C0uZjY6/moinXuvM1aEhp34c/US4oczD8d
megTZuFBP6tP+ZE31aQPFrwxyjnKJYFxLyavAH6BpA/oXiztsedITBDpK8wHvVce
qI4Pgr0kVCbwHZ3H3eLqWlJyctj9MteFejwxwH9ZuJmuUlS3iC8YKn7in147Docg
Oxmpc6/dX5wIl3PfyIawxGhRYxAjYWQntbjXZX1TiSWfr/5fQe5LKPMRm0mg7lI8
CnOnaCxTnii6rR31kxppW2/052EjR4mzbXdRf/y6ZOd/O2U7U7zTSNhWMo/6F+Eh
aRZVvnvvyZYD62bDqOJjrJ/97U///tjzRAHb4VWYdWyMf8cNRBvR63l2NWSU6UuY
jybgTgM2v4fC+f//KX9y2Yj7fJOnMWDwb8LdWbBQc1ivBhDzw8ne5fBJsI1g+D8E
UVkwx8bxmKbaWzvXF1zR8d12IHYe1rSjwLOke3K/dpDRp3UmXWHdtMasChaycGUz
v2cRmZJjLVObJqG29blgq0/lcBjOjeCxrG21fMqKBC8fhx53JCyPjkhXNdg0FBcI
oUGT65fUbBuX5wXv3gA8cH715sNjW1YOKlLxT4KFQtyNLH6fgQgMzi5jsFFJu/Vd
bati3Uv89jnxYKtZF/taV9DZUCQ+l5yWcyzYwLrb45JcmSxU+NsBHl1IZUJH6mNI
B/R8tGa7yBhY2lyPA88jjXWmBjczUKEXFVKqjRtJ1+X6+j+QvAX+O6hvZ5I1xb+U
ts7Nw1oZOEkkRk2FqDswK93NhG5k7dOTJ8P29fWGZ9MiLItGgoTJXaKYmfGvCKGM
QvAj5EsVqhXFIJ9Cvhv50yBiuX2WVAdnyPzmA9slp+Xy52/dhYyikHCU86bkUfYf
V1mLQrfu4TYSMuv9or2oL8rDpBHamJjaS6CFqRmT90DPbmtAOT8r39EmnjeLl1Z3
TmXad3jYBj5Q4gbJcCgpuraq+GTQirx2fb1QSrWguUPVkfMx/FoUbj3XxVs0T/aA
Fq/ERhAhvbpILHjZg5ciFqjne4dnowTUHfATH39azeC5QW2PzhmNKDZEEHPyysQV
fiHf7YVcu11MK+KcLly8qPE3PEvutL2ce3dtJcPyeIHnbd1aUiyY2Bs/ARNcd+GE
ddWOaNpBPrC7dKOm+0C3NpL09NRDBEDqWPbWrA/H/npC5p+NPG4VrY3XVOtcFR0v
fLo5KVcnBM4bZkWTz9r+6m1wAnCceZOR/ahO84QbjlOD+XdHg2jAMFln11II726F
3Qk3/1Igj/jxzA4u0DSPaQqE42IPXl8D5kqv4IK4+0xM3egavs9omZP8jx5j6DCh
WW40fKD1nwMPQowJTBSUn1SAyXXT5etd/MtieR8DaBaBqU7l4JZtwLcKxhi0b7PY
/QU2cZk5vtz/FoZLqeOjtqr8PpoemESS/GbNYaz0Yc8mXc99FHRzvGrExC2+W19J
Tx1zr12/KwEbEFnLrQAiFIk4kk1wCc2LObwSK35DQ+TFldRZDNQMJ3Wj21k++nmw
k5W3pb7vlSMB1TjctE8YqTMQ4RRD6VOOXD5RLp4ELk8OCP9iN3fK6hA+94takSAc
WrExVTUOGxUAj4ZarbCllg0o3bci+5/0fXqYcJ7d7UTfJV7xg/QOHCbdzLUBs89h
ehGXxGo1hj4gLmgdc/6kbuCVc8fNa05yYuJF84RWhv0N5S7tSr8UGt+3cbe2i+A6
XLCaSpJ82gh50w25WwxwaMIoFo1v9FPgiZZPuV2ZQhZHXTRO2tVHYuf1fCeYjC/X
v5BaEI04FpMhEug4iMd4uYkO1WzazXr3sc2x32Ma6omIJB44hDDcZFJg85tMnWbV
MQ6yUjRkFXlrTj8piMgsK3bdEBAKlVHOnekSaLU5Vk5eMSQSCUuAbqrZqnt9lGqN
0HPapRJmLtbVKvsEoMlEMhQyQlE7OmDA+8IEfUQQ7EbthUXTFW1JHVz6fFmQmeiD
LqkMXeB6Fu9q2sgv3s8LMiRKLS4DQ1lBWwk4jh/tpbabcl5BEMofc616lDDg95md
uZqP7bbKxa+FtvcsiocRMHPM5kzFYuN2CFYdjCdg1zmw6JzU+1lVooxFuu/aioFx
ZRRdFF3JUMtZhNcpXBs9ue8AMpn+/dj9PAfxkKZXb9LAhfHBtoqhtie6zok+tQhP
mchuGkTbHVMv112+vE+2KRSSKmTtIkKb5ZukUkMeYq7uJldoI1oTs7EpDF5o8duA
b2l544whK8u5seBAtb2vJi3baIAzu6aqbStgK5j4w3m8XuVIBw7FOqUG4ATvew05
1WVoQ3Mjr1f1zGKbEha00iwldl9IDmBskkK4e+MVjR2BMPV9t2guuWR8jVmPz3L1
sv1NX6xuXpxuMxf0ejDhwuTkghkyCFSFbpiXzfHcI6koEYRW+Wl06Ve5tCIOV5SL
JhTKuqoTYjaEitg47vsDocRqmRXEhWE/XyMa/Ia8hVgxEI2nx9+GnSpgL3ou/KC4
fYqovH0bz18pbf6HluiqowZyBPl+foGKZ8En4OExoCQtvoYmjPFrPN/YpN9O4dN9
4IoOQo78R5zdNiTHvTH5oyNkshuS+pBla3meD1S9h9S/UqjRlEE60aWZB0AEZ9/V
fULpd78QTtlT8ZhOGX9bJAXm/4HYoN3IstW9HyArdRLErl9/O3OQlu4QOKN2ECe3
upYXYJ/W5mBAhpoisL5wsHxWzHgZNQ3LhAXSlYsB0C/TMsvHzqKMhA3FQFxsvZ9l
AoIcVKeOqFxgM2Qjk+d9Roms4645Iy9Kqt7HzXhpVYKIUNclMwuQqt1RmGcNS4Fn
4caA4xm2hQ0oQf76kHZDsrLkQgI4PS0i7AzOxhPLNhTF/FmoOMZXnfqWeyTmW1/+
xqygmzmT5mO9O/zuWA7b1PpdVqoyZ5URNhLCPqtktr0fZcg8Mob0gICCEFZxsdmK
iLFcJ7B6ZpMgPo0kerv0ti2X+hwCN0WA1MsglEEbUgbJCqqC4aL/JIwa8aRdtWft
ms5ovuhVNAPh2KvxYNfmVrW0W4Ng+A6Zti+O8mRTtXYmjIFN0LhMHGAt5yioLE5P
+PjSN7Uo/vaJ5+yOUs1Loo2hry6X25ehu8rqTk/KBBmCXxbCR1Xos/2XXWANAi3x
Ks724xUrZZr12gQmFl128qMPKJtcaFbJepSKrFgbJU4hN1/nmKw+q6aQHsnQBzPh
LSqfoK08iO42did9JamcVczIdWkreB0FocctWNIunKc7nsLX55eRYWDP7sXUHv6T
8pozoVN6nealKgfzxu21Nw2oliLJFnkKkuls5ocCqhVTQuP3n018JnaTMj5z0ykA
FjYydcUA3Z0B+GKIP+5sVaLbR04Y8V7bB2IYEAMputsFno3R4orJhaWm2Lwy6XMF
6hw8mD2DiGS3PmZj7pdOBDlXO69lbFV1QhViubWbY/C8gX/vhDJFRwirwJQoCxoA
ks/BCSGdLaHLuat70KeNBvGrhMSqXXB11bgfZtqhie6ReMMKgzdDng2YqjqgEjcw
rwqy8lwVNrx1gJlT2EkQmXtkCLSAmLQ67hPyZ3cqCzMdqS/R/ewbPfOqX1GqDL4p
hbduy1KY1HJkJi7qMmwY1Tegwy/72vrf8nEN3sEMlsYFZzsPVPw4CrKzZ7rZqu+W
q5/RXnr6kBXqHOMFMNsw/9T370+FwRuQTm5MHAuu2stMGcoEB+Yc96MurcWbrDZS
VExr/jqIXm9ReMwjX190jgTFBtMGehWIHm1MJsYOq0JaDOa9zms8zSntr9J5i7qC
CXVQELPB04KbV4e30AXDdR7IHokIlNox9DRhBY9MhbghOpiMnmC1fHokiFeXGJm3
ryyMRoj0QHKUzWIYfGVVwF6GoX7RFGa4Anr3Et+ybzCN/E269XRP1HdusjyGah/A
joXf7doB0WDrB6jEKgGK6flzSoJlqjZ5FMQ1pZg1IkmZC7jxvoaYZ1Ajiko6FU+w
waGYUH6VPBUb3R83iqkB50Mu3Wr58X+y1of8N9Vp6wfBA4DLzelAhhBHehjKBOwK
LyW+1fCTWtllk0bpFzSGGcZ199nlvBlwCIw4JbKQaVySb3xdtN/4JKz2aPGLL2SG
w1JhKHK4i/x5hcXlXKkwG0/a3SGKa0aHJw6QLtRgqzISRB2UfZTfRz8inn89ZPF7
x4S+j1ajoSFFy6Hz50G60mPt/YYkNfcell0h/XaTA56Ip4Xbgq5laOKggK5oWY2k
dF72Fhv7k4o1kw0S8V3Xu+2/RPC7jnbeajVad+nPp6Ma0c6k8hnOz4xJXCZez2tT
iIaPHPxKZFPaX5LghmoQEugk8PL3q3CF90Hsy+rlceSOxQ08Llxh8kdU1KaJy2b/
b9cHfmPtTsxaJr1FL1tBAiY2w+6CsNwwCCtzHfLoMs/XDVUvIxAifgb0g5Mr5/se
rVrgTc/5dKlCd95q7aZvMBNBLzZBXRfNWfU/E+C3U0/SwWODPJpkW3P3/JNNnps7
rYof4cfGV2JyVazBDoVZ2Fzoc+j4k27219VkL/2yAN78EQaPguyp6NG6Z6EKN0zQ
r/Y5SPf2OAyTvAYrlu+Rmzdu1CZ28J+QhRKonpXMcc4VffMZAE/KvrAPKZTjJ39T
NSJm4vVNorH4EQqxVWU/QNoJ33Xsbhf+4yFnXIkBq9y+G/VQMwVwEsF11xNc7P+r
ibS8+P43ujej7vVyjiy5puHXMLeDHcic5MoGxOxKZBqMTrp5EID1U+jst6bBB5Xf
ieb0xMVqynfKzqfB+Nv/EgA5W830DrZzDbXywyHlRsktza76cCsxThhjGigH/2Bk
2nuWlnAyH3L9iyVPalW+2juj2QBBKmpuhRyC6dooOczizXDib3f+9Jxodze53wz7
JVJJCuSA9dAMtZwpjuHDfXuGpUMSjA7ama9/7HDhwsQEgReAGL4Jd8nB0uUEhe8Z
E22j2UNoKzl5zmmneuliBeauI4NP8CAzg314cAYR35H8JZRNKKjk87sxoBJRsLJg
9GqOSfGX8AicloRwLmt/Wi7U/RYFrx74N4aW8VBfrJE33lMog7sWAaBoljKQU1vG
fcpoxYcG85Zkh4iOxzksxh4SnVZ8eCLTntPN5PHx+NCcvokKpehzswJMuFxCzOzK
26nIUlFlgSJNGSgtt65hMpjLgNf+7xtue0CmR+sy0eC5vr2+fK2DR521UKZfHMZU
1a727b3Q8m9WibROhy/VABiVnZd2GDBviN68JCjnrg7Th4+fN7MUQRQsAh+Htskw
/TER6DKdLldlGu0exSvnhc91lhFIFl++XUME0GbmBSBA6LyrYi94hfj/8gE7pIEW
3pCA0sSYgnS6OjlJVD5p7J7OvdnTh+xMQsOUecuiTXQUfMZqDT/NJojP+IvKDpkS
DJVA4O2KG90+k1koxaPt+RuL1iTRxNfeq73Aldj7JhgXiHtbhD1u80Uzvp10xQK8
6xiLTCfm3zEZCAxHG8F4V1N3Waeo/us/nRJFNl12VcrvUZFbeqDgl3NGiaZ+F3L2
arb+twTQ01OFWfcZyl2yYctwtr5oBt4kyXSLSQpa5RNV7gKXaPceS1IPYDy2AomP
3jbQyHBtnTfGRQIS7STiYyY35E2kCwzQdE8EfxXEbM1P+NOJUQ0hWMYkrSEy3wBy
Wz4nWux15tST1aIVXyRDhJ5pYnBbfPjOMUBlFDeFvBmIiwevG6/XOo6p0nLaSTKj
mETU2ei25x+TriTEeV4uoi5F/ok3rYz7ZxPIJrAKwEl9uCNNbiWJue4jV3S8CHRn
pRwYiZiQvY3BfFXU9ralu6yBaWNZVDRUrF6WXRrbcO/624mxhUPF4Sp5KXqKuVoN
q9I49tmjTixqtFQ1HqgTV7jxp3h+j+eE2pyt6Ev/fS1dNOJoiYoMB3e9//OubEvy
EMh8TMVpkdqkKSqCkkdynMeEfYEKV8kUOw9vj0sEnugVNATOIJxZv7ElQjD9UBTX
CA8vMx0TUe2b3dEHuZbRH9wlvFxHl6UlCs9X6bsYJb4G7iq/8+SV/3agbeFv1W01
Gjieq7umwJbeMJZS71vrkPxb9RVZJq5cqVHOPeMPLIIhKBmG0+/6Jbjjvk9dhl+v
XAid8kbwwY/UYYv5jb2SPipvIKNIRpzMDu1akZ7paHLT+9BsutQBqVKlkZt72H1n
wsjayDHYHwuW4tv2c+lX9n/VJ+/ShWO/EfXnOx0LRc22za46nflyzpmCcFe9AZHO
Qo+7iJPDWBegAAcywqbaLrfGxKoVqBS//PEqru2msBSR6Sd498uhrV2zfoE3G1Sk
bhAiENoB5xWfiggTf6n9X9MqZ3MbtwoOnbwXqvHoYqmOgcuXb+6t03SPzUDLDpUF
gQ8UiZaoTr9CP4+PCha3CkRobTXhIeIZQAEIvHhru9fHXLNSaWs0/9MnSDtu5UVT
2eVB04drk+tq650twM4TtSOOxbbMEw/MGBRmBU/+qPWmWEqNU7BLLIbHEgQEQ85Z
6Ca8rTvHJ0dvbn8XtksyJr4S5ctwj6YfjUrHtrb1lqInGy5kjUUbx5hHtFVWsDJa
QtSKRvy0WWahDKtgKNK8e9eHuWjD93wQMVUJx3REgDTw5XpkVAKkoS/yjsKnqVRB
fxoOyA8hRdLjmUysiDYyYTHHBNZoGM8UmxRValWnoGubgNmA+3I1y//z6CwQS0Z8
h1Omp8GDTfSb9qQNE8AkoDqbF3hVKlkABhyYoCpPPRt/MG7m1g6V+aYCLYF7G5Rr
7dswRVU61kBwXS6iPn4aUK20BGaOl8cKkCJ2Yj3XyorXzBPk9OSuT+qM1HW7OFgy
7bHhKqulTigxA8gcIV2O+da0wvuW4WV7stT8TYQB4LtYjWXqT0YSqXjpnnlHg8iy
pLZjU9huSDlTYgnIWzWuB3eI4xTKvY9aoc+bE4/MXdA38X2Ywd0Xc5n5P9UD1RgJ
SD6w9S4pjVNt+TxRQaodTGf4OWyYYpiZ/G8MbDo5IaWYLWPOz2g6MA1P9OO4/PhH
jwL1rHt2KOXG7gqV6f0fL3rwOdqPin5P2u02hwR7lMbcS8Kz/sdRe6tgWjeI+IBu
XeBh24JpmMm4Q6p8sMJMlNFbPpI21+vGn7RZ3RW6kmNjgvWv0amw06xX3W3eLhW8
WggLKG+RVCrghVmlmCiUW0tY8f6B0vLvOT6i67X5WDchGc0VpV+qElvS3cl8Hk08
eXxfSB+2IFc/WKY4BiA6/4/GvPOUDY7AUZL98YXdV/8QfyzLZ3MS9VcUlQic4UUh
HJKrfUdph7DWSQSLeNUvUXi16YxVh0ALmTseo4W5UK8G8ppD8/uARGzKihzWwfZ+
1JmKZJ/J46m54+UqhEI/E9lnjFThhf+LaKsNidRCB0qPKTkRViSFTFFyOsupz7oR
FIA8pPbwoCxxtyBqb2pxRevv9RoNDdASUchgD0pJJUiTDhghQoWJ4zempcnzUnuD
nCbQQ/aQxgqAkBoLVoRYbo62xqws8sXiZazevQkVTF5PHtLmrZqqiyy2AiGQcJav
pTpx7WjPCFDTTCtSn5xuM4hNG9D8YNp6vbsWxQDHJSACaTVxyQjNFu9bHsEb9mcv
061YfWXGadVv5c5Qe+WIHJzTLn9EIWXIGlyLO2XVxGDWRMDpUFv4aHuiKbZzVCWS
jcomoyd3K4d4vVcfHeEEfk2g68LFdnHyjtcaLcylIV9eC3Azily1JcsbPv4tnAU6
9I/J7uND8bLQBtyBlQiubbV71JpbniH4fnZeO4NVixBDQ4pLc0r7s2hrO+Jp2cP2
JEwNv7+ANJv/ABLVNUywRtfJXrMfEAtwkZ4AJETxdQ6IBOZiDp+tkDCGAucWKnBS
nhIXxnNDD7nsgpkJtAYVl9kxFYUXQ/jmGNpeOHf3TX8e/bnqzFBF6d0gycRMsCTf
i7YWoWlXDdkbQ/VernCRRxNRQfwmBXndjA78Ci4bshPbbFKFhWcKt8TS9jia5Ts+
O9P3NRtRKryrLeVnSi/0RyH3tQey1kqw4aQ/PQsKDFK9jh2/XtfSQ+0uULzCoBqx
YgmZUQs5gFW0BJb2U/xgcKWLsGrZsnlrp/IgyLmdNcRyPDpYTmjgjaxef5rkpnAe
TvVp5em8/tWaS2bpjb7f5HUjwaFwAR+A+s1lZDZtnnL4avuosyRk46pb+yE/gKSG
Tc+nKomKv/yPNHPQscKffuVslYtYx6aGku0I1JtydjvioZFBqSy4FoaRxEoWkuMG
pRiLVdslsZMR8T0iHXxiQjv2VWMx7A5DOoHwQmqdzH3PZboS78c/l09x05tRncLd
FSRk6zubWO8RuC4u3vqOkrx3hcshpEkRivuCYEBS4dzQLe/4ORd+0mIE+bv23ZP+
zvviujHAzp1td75BVwTBEis1O3Vh+1bfmKQRBapnmtUrbXk0cjWe/FQZo8u1pUgA
ruUDFBUSfPxRDBWm8dLF+1coe1bpg+58Wfw5UqYZpc47tmXq94sByDeJPkIUYlTK
Dva40FFZcjouS+GoKvZRqyJPYzuRbhkbReITc1xlbYdwdhe06OSqanBLr91jBeIb
Rm3qp284bDrbujQMxcO3LQio6o3febo18FOddpbOfSQQobaj9sw/uf1lMm/umLSt
G85eoFBiOVkBL+XTtlnXgdTdWHB8m4pDzeOnSdk6NMl7si1pP6PIWrAoxMWiz5U8
+r0fhyPcHkP4Y6fnqERfaM21iXKcaNxBi8r7f2LEY/lPRVBM3CrsZJHxISEdgo2Z
sE6FLV6IpV4RZJRFlotHqgOA6p6qYory6bSWo85SGfe3uhG4Oh+kQpwPb59TuaQT
a7q9r64K+nZjOuZFg5N2lLRn6vdRFixWlD49cYKD6xW+etEZOZJdWW6+keeRp5xg
hgkQZ86HLaM5/45YAEDew1ti3gjGLhH42FMDcm08fhKOzMxwN2an8N1o7DfyKHCl
Oprq5nwnRfX7HavCAREc2MRUC0KVu7uBEEjaq6dwmG0G8OTQjuHhQ+Onr7CNyMnQ
SMEa082cpgUCw+rEr8ksma4GcG/ExBZBVfoVCgvjU0pQaUtjybUsVZp3lGqCZzls
q/O4OTyaI047h85mKfcHcP6OoMDXeq0eb7yL2/1meHcl3F+QqVAVRd2Me9mbhFZy
r78VJv5AQ6ZVcm23S55QY7VuxCMyYEc8vH+fHup8t0fBkzO6auTuIXjHT0azJ2Uj
7+odQa0pBndLGNXvt3fqQXWsHDGEFu6wztU2592tSE2zfmZec+vHpJqxkyI4jsld
OT2DPcoZlE74/nMMD3kCJl/TEnCDIoAnYoPVhrTXoXGKoHfLzg5efPXy/7CWTH5M
1+w3cpr3nXiOCx/E7NcIFkT26TYVeJjXxpPD51rLDaBJe7RimK0nBcXqRePvEHmU
Y1tzQ0C7Q41yU+co0ylRdAA2RFEtUdBGN0/s5mkg+GVrsnbrjhzrmEHS1keswdTC
+a/2iTZImWe7XwGg6g51KaC8fWocsE+D1xwF5lpQcbgWEOr8e9IZeXGLy6eMQ3oX
45TfdgS5EbnqhqZb6/73fwuPz/M1Zthj/6WX8fNcV6pbszMO+QfD0fdtoEWiRTTF
4x/XDo8btNI9hVDOaz9AtG4l/ks0i5UlxfYAEgb0RZA0MySj9a1cK57w0PgtKr5s
Zrfg2rpQzgZRGeYH4Z7DASQB/S1MNJyUujJeRtULSz/1QDnxpea+gAOfpH6CyZ2x
1FI9nRPnU7Pdmb/x0CCPUxw1nyvbEQmo07fIaEQJ3b1BNiI6sp6XExyeZaxqnCWV
ZNvvp4YgVGct+oikh7BoFF9QREMqHem0JdN9mdcWZNnbmdyNjkr8gRFM3OpqclaX
StVhFVBUguwo47+tpCnlWFsT02EkLC1LM3fzQGoQUcl+bLmiNJXH8QEMo6xLNw2j
ue6HM0wH705JE8Zq3L88x1s3b8iVtR2wr1ktjPaPCqjRo02plvhIYRc5n6BGbkDQ
Zy6gJcd0GNqOl9oGJfHKSfFbloEppMnZsY7mbcLjykgAqHjr9b0Mwwagrvz20MZO
7QYO7IBuoHdLKzpNk4Mv5F2SJ8EnsgY7YJbLELwi0fhuHOozadDzSPlNsa6FPzcz
/JuRYr7Wxpdvvmwje2Y6QgxILPg5E/ao6AFPsAHucSyNagtRXdLpp/KcwmVzgbXG
xU9bidMPHdLzZlAseWW43VrEkQXbRT+BkyMz5Utp5K/yOkd4YgluufiQqai3xiB2
xW5nMNk8IC5x44MZnQ4knbmawP7pMtjwm5rN0HMXr/qK6mFS4sZhxSM+T5MxW1UI
f5jSlt4cEcXlwNplGcBhQEHzPj/p4E/yNMU6aOYe66tzGcN7a45xXaPSuHE9UWmX
nZ7IdbygsH/oq021e3ZYKli6Om3qOq1I6vHHEkS5WqrC/jF4c9S2/3+VKXaFY7AY
lSTBfLXJDyqNW9OU5ZLpEcSeF/SM3/t1iWUqM0MCK8FgGHAntppLDLoiBq0srvyF
zCFYLcoIQcWGi8qhKdp08If34im4INqgWguluWxH0NYTpCbsAbf5WImp3ZDCbr+o
POcRUxSH9GKAOsDxKvOTxHTdZQglKnpBEgB5/s57xjOjAdCqRH4/RiUyaF/v/2pd
bBSVhwudIyWi7V6uLmhQ4EvPoegz5FH/9rP0eCOM/LASPWptxBMvUNJBlmLuGVzO
+sO7Zu/RS3ms7wg3yw9CrfAWVVNrQ9JnWCZ0yyf+45luoee9kqHx4TpdlitkURAi
Wibw1vvdVIThQgAAyITshEyaJdWyef9yNf7BeuUswL+MiqvJxPvkdUsy5AvKfaqy
FA4XoPCxExMDXcVpiiRnSyIGwfofAEeh80tZGDTYVstdxjdiQMmkyL3HxDybpBkT
9YUBRM9/l1gwiNd50eRX/ws/M/ryoojp0g1to7tfVDxtvWmWINJHkZaA1x+r1nCT
8cDuxzBmovHHihLgTJmd23XIZdKAAd7IeY7XJWb3fSOPCBhS1QOtkXW6o7gnOYSN
eW7bqrkfbrEccJtyM7cpzr6DLrUW/RwYcXw6tidEzd5qyyRIF/yhIvn/HK7rtz5J
a6RYW8jaFLwFyMKS9zSOMKq3tGFYvFRlkcLJsEuIXs/Ll46yLsbKRPIu1gBmePMX
1sFWxEOa2tWsavr+PiMSWNhFQXhU1vgLmDMyXVUug9GXE80rRUVwgqjfowmOZXiu
70NSmNXy1y8xSaj4zsAafVKaec8kMDp/fPvLYsoD9sKpn3LlNCA62C6197Vw/OFu
QEGbwjvp2RmFeLI4XAiNIlINgC43/xXZP7dlqjdtedAhCpdpMK2k9RoPSKmJYqPg
Qt/Mt6OIG9v5/LxDdNgh7ZMOeqtOS9ihc2UmqkOZjCIo5xuLsbED+qxYQB9FPeX8
en3v0w7IccmKD2uaHUB4k7AnXTnXzhr3HkDCt0Phggemey47KgQ46nl6Y43Mdvd8
p9Cb+8Rx7iVX3R0AwtlKvG1vIMMkSHqdQ74HrQY8M1pdjsvzi5JJ6QN/7L0O8C4V
G0s+CnDJ7dnGnSL2yJxAnQv5vDkwRgM/fC2o7xtPA1A8W7P907orbt92psKv4TCL
sdxoYru3L+ffS4wGbtVmoB44IN4WA/Bh3PwGTE6qPwwg8APEoDe9kJtICM8dHdgw
krA/5Rh2nWdw1a/nvR1cdmTQKalnFq+1H9exPR9CG3qtGMkrsEOKKZARUHSfANCp
nAmGeXYSThSdRI0LiWICNPAwLsi9zusiyTjYrVqn0IffqAeWzxSfFtdI6M/UBziU
6sYG3tATASgjJ9QO0AbdfTT1esOwyluYCwwrWF5Ux3twwENZ2l9OOqIMCiVkBpA7
hiKlsoYtRQbuvwgo1IiwsXMeV8UmwHGB4lShjUdEKVbZspxbBls7CayVX+vG5IRp
PHN0T8bO1EQDoa5D/tYNbGxxWf1GWq8ygGZxqOmWesrV7R1QvfTXZ2yt0Jj/ndIy
JRB1OIbTkaSAeihGwkGIzdImi11DXEvS3URqzGXHVkMzfnH6pW0OPKija4UlR0bW
pPawVGiHzyjNEQ1Dihdei5TmXuHM/7QnBIr5qgnuZlbIOvXjl7jVGXtE/Y82dEtA
JsQ3BtQ3a0b11esMOSptjJ0yw6DgJcv/ssks+fz+mGRhVfLUgHy7uUzpO61apVPM
TRmi5BuIluoNHrFRf6BKpo+muDy6JZ1miYb4EJXC7b0xmfHVOqeqVLyo6ps8MHYe
PObpQOTFhqC07SYyM8qLwSNFBGCTbpHEM7duUSjMIIz6GxDfmiFD/3W9gHpWX/ol
0TKXRkhdnWQXvC+TsxSjLAZe/Zm0UtIJg3wLalTdaDi+glzrWvmbk2xiNhaV7EPe
VWNBOedFNlpx3D2O7YVaGsYECFde7N/qloASCI3g/D/Eu3cdnRAM/rRqBGIBKllK
AINiD3h5l41O0oIaiAfgHNfePUPt9HEtzoBfWnPXiF/qzNkL8J82CpAoxMHzAD3i
Omlp8qnJhkajJ7TGiGRNMBnVuitFyiQaTonmCCX2wbBJurLirgCmOLMi3OuXZvoS
30Vqw9o9v2uatmT9ICGH3jWJMpsaBrajS2jnuQBqftBPfxhIttPS1Es7PG9mvlAB
aNbhIuh3a0YNcwn/eg3iKbn1qDi7XU9MYwYxn9rQgnY77aS1BY+rPGfH5OBODW2F
ec14lqct2pXzGRWkSjz/c2RIhOPu5phjL7F41QJkE6D/73pfqWsh7UvqDlZLQOZ0
dvPxd0e+MbToH8RrQTQtDFLjq5w3OYrD/KbAynMyX+ZL/wqm9yxkUoYWnrlAIsj/
ydOr6JMwGYuwY3kqpJWzrTzLPmhkaQlNGCWvBfBUe2YWQEOYeDN4yUBTeI88ylij
tXD+trlhSF2v7KRzUSnc7Lv9y/bOMt+P1hmCYTIKcnmgHXgaZhlhYQ09hLD6bWZk
TouEeYujmI6Q9zQ0P7vZW45DeIF/MltdBTL8xP26gICGKo3UEijPN7hQSR2CAukH
xGY+fqDHB09sWk4z+81GjofWJRzWE3IpZgwH4eqY3bD63z6qF5qKigT/MXD08CiF
jumsj5yh2+BuhMF7Abz0e9iMQgNp1dOqfZ117JF5Q5YKv9bDCLUhniMSHlOu0Cr3
GyL18PGgcrw9yOjDkPZG7aNRNT1+ynNmBvMEwguJ6VNLr93dAykn+4Pq/G+pqeG2
P3SRs7PNLYV5UK/kkYf7m2zew1pFCopEHIHrX6G0TpGxdN4jdMhpMUIOCFkdAL/y
ZbH9R6OFioyrQ93jjixXJS4+MJ+tSD6+yzRJxOHZXgbMREI3VKc+LgG/ZqcSTjGP
BJ5YRcJrN3BVEY+hPwK62mgPi0KGW/B8x0vixogoqhDW+8GZQ+ptIw9y4nkSPQUJ
ENAIdpJOuyjwx2WX/xV3OJthGnBU8JtiKlR4uFoIbnHPVDb2wFjqQlEHPq5wrTWi
q5PVdXST87CDybUHtKo5o0gWtdvDmazhgivB/J+mB+0hN57+zOQYMFPfQhOM7h2z
Q/CW3ZVu75XegkMcwJwGh6GhS8sENRm+DcRjB29DGfLSNxLe506o9UZE0gfwB3V+
5A+5MpFrMvvA222XNyko3IG5E4YUxp32ecrH1DVT6wYYUAjG+juU9cZd4SPvqO5N
i1xo6TlNDx1WId+LCP/tmfHJSs+3YxfD+x/CSxhU2BM8y1mofUfwDOSc1LbLF7KB
OGmHm5b7lghewjeMZQxR+m4rio9lAMNWXA94ECrdmjSR4rZ3lgfFsZ08WdgX8yD6
G19EeeiL9krLp/Hxm5ylDvTdS2hAMbbGawgK+KE+cpT6wMl31Lp/3ijO0rxgKzXh
Lgg9UFDu0gobbGEfh5EWLJs4+r6wjhPVKVQw54rvicfEWD/8tK8ABEZ1yjuCKGQh
2OLSVVPxANLmPbc//rrVewXWvM3lUtzcZo97bS9Rx3AloMyY5KLVe7YTQ+CUXYnL
VQbV3rQfWkJiT4Ph+/6hQSDmZkoH6gX1P8pznzhL4fUvKxT5hLq9/DEKGR3roSn3
BCaqLGamY8NSEGV4t084gIYt/gJ/j47HWXCum523kB8BofOkeGSeBK/pWhkwsoeH
cjdp6IP6PZVT4Qql6a15OPckuELN9idb795BZCu+igV8VWroblw0P55qBNJJGq4L
FyRRwSc/jf7iGIk5BIRc4J0yWMqxzPEGpcUhkYE6ICqkm8vPcjDu3vH+z49+pvSo
Z3I9c3T/ECcLK3kHQAYVbmeyrvJh5Es1PEEpZXGBQAshz6WRqvH9t8P+/vFXanTB
gST6qYByy9Hkkr+1wjdCb9UkjCfoJzbTLWRgoyMa3f4FBPk2NWOMB+UkH8dELIsk
aHZloysIjNxqaEWnAUJEZ4fOYJPzyUZqVmUPzjHiJ/6xgcL0NmwQQaZKXlyschhN
888cnSYGniSsac1gmSCpzFVV6Taz/FAyL3op55cSoSf3FaKQH4mAYvgEHp4N7qaz
GQbGe8J6sxdYgqBrpUBzOba5EG6VjAkbrlbFjD3ezFMMAnG/m1AcnEp1cNwo1DXI
eREqToPjWZ/7opgwyPDQI2Ii8TZTHctnBtm8/gRkzSC1lk6JaIa8yrRFhaupYn2l
Thj+TP14LmLK615K6E02cIq3ixiHo1XAT7kweFeI+nwDCj7rm7auB6fxk3TFcupK
Tpr9a+rIJL8ccvdjFBpqSSqWmrK/VuxiT2MxZNr9Up3dtL/HvyuwqyvBIYshZLtt
xx3QfqIO7zfo4DtUHybfC17tDtnGXY/HdO5hbUMwfCJx9iobfze9ZjBv4jSDsWMu
EX3e6y4fGLQLIldOYsD89zAU6G1ctKC5VZEI74RRYvk4TfoRd6YTbwp7NT9nDs54
n/SMe/RS4upOEUOGYpddaTQw7G9HWwNt9kIxost3WnmtTrgmjSCEWsRXfhGBZh2T
FqDdUKlLRi3hTEMM3x9nVPmFXMKhDYlVxd2CT8TC8o00MXtLr+f+/TWslG1Bfwko
8AbWE0pjMO64fONS2h5VyvK6Vp53PIaPI6Z4+Rs/X/ltUXrButavTyjb/mAtn0jS
1Buozm0jMSlTF7OAPPbizBbc3MRY31UQe9TNiYDmAEF+IHmSLxkBlhz3hnMdOJNj
5yShgA7bxc0fwfPgVGrjqkzNiCtDPQWcycQfKDvHDldwMYi2VLuN8/QxCVxIQTq8
0QuFMlDcEf/FlVfR/YocMR25WXoI5Bi/9WqMkFGsKPzyn3twxyA3I+FySFXuA6/6
DgTBennt+ehUeTfC1h0rIiNLgamJBPN7bvqMEdNulCR2rD7NvGSJots5MEW9KhSC
R6HpJiWdbUpqE/ZqL/vY6cya9qCGKXvUfnwwnTJTjl1ViB1Mxa7bW27AEZeQKx4q
GjeMypgtFnB6zqODp6D+CEP/0JdRkBkkQCJXl4oxDWCZLNA+IdkRUwhGrqheOaH0
rfdIdcYH4B9v1W4krnB0de6DiMk/gPODoLI+YXabejZmy5vKN0jUParxi9iz4C58
LabDEaqAUoW/u5iw9SspIRdxB5NvMMm3PMF0z9M077iadpXK2e+BDNUE1RdOQMbY
wv6it5MangJdMproNyddGez56RLFGQT3nj/Ahxny7nwfHY9T5rUZp0LgOmVnGV05
9K2k7ouJvLiQT2ZFdJ2VGwIBUoVMOhbF7fGfQMZalpJa7UO+LzqikNLRu0z7alTn
NMckVWHcexPo4Ad39bIS68ofIn+SlmLU1lZaye007ryZx5kgbj4xX8pjDqMHoXqE
oRSYNpcgwZhxEV0J7Wrp8LfyJP9Ch2zMnFCeDBx9RpL0qMCAQEcE1BKx/D3BZ36b
AI6GT9/p11lwbwvtCX+5uaEJ7iZMjMlwlYPEsSbL6KMF791eg8rHXlLkQ8xBS1gD
dw9TLDm9JxiIWQe5tvXrepIAvrgu9J9WjTSRw2DSnwXARGSouw8xg2w40/4b077X
cLGWjV7Rf0p7VXZTKGfUp9xyZky5po+zG6JOTRdov1l5P540UOOD4shtYXNgO8WQ
rHXuiVSZfXp02CqWbVlhpYYiXIdGBuYHaz+Kvnf07a+sM3rJufmBs/9FkdoKPXZn
xBbrbiEIb6/J5mJ0uqQZ4HV/7WHkdPW/LDRtHf5NjLJzG/rs2w+qB5oJA3jOgMx8
oj6hh1lJP8i8vAN8P12yJAolE1LGmHwENiq/xRji4CX2C6iqPUYzG5NtKyuMO2Ti
kIw0Cd8+vYt2lL9iyQJFI7of4P3nUSkeXOrwZMmu8ZaXqHOz0tYbHtFsVRlXOEF9
nI5bAdb/R7YAlKbQz5StBbNpF4tZW5UbsOsLi9Khd2P8fXcI/OA4z8HE8XrjCZ1q
Lw6cW+M/8PM82UKMczI14EvbFQHWPeF0DURUT0diBDy3GhucY5vW9ss7Ca9dsuco
iHZspXwAZxzLUQg154tpDdAY1UBnKPq0pk7utdBSdTHQZPua/QNqQ7Im+ZVMS/GX
73sW9lLAFwH+MY6TszCJ6kU1VpuO+RCinkWLtFSzRiCDxnFzLKxVbgFLsMEwZbQb
mx2Kr8MvWLA5htLGnBYxA8h61ZG8209n4iF2RSEa42IkEOVA9abvApIIFOW5FMVU
SBNsbhpJST1A9OE14rS6/6XzIdMkSJv1ADn/JNzR8IKb/BfaucbOD4lLg1aF53WR
sS7CMAjYEGfPc8gPBV8Il4Hh0DMK5BySY1lCZnZbFHoAqJr9Jfh1LISY0R6AkbUG
X6lM7m5mSun03WRfob5drY2k1Gtj8psy4pED5I0prA35qaKT0q7mYBVFY6yV28IJ
HqQplyMu1nBINJrzKghneMGfp6GXKiPVIWKkzHy36hcvM56pXUIep7+5iWL/rB/Z
3eMKK6Rr8Km6ECeiZQdEesmTBuhKtT77tPQaBRyPtILtMrFctDE2ktXdOOq2py+d
BdPApkAWRDdsUzhmHq2d81G3OW2PZ9dnn8Sql9+M/gMt2UI1Nl95sjesNhBar0UC
8E51h2qEdRVRoabSpkhTCaeo6+0AjqiytLTPjaMyn556gUm2SPVY9I2KQy3eQYgW
flqMgmJVctn0kZ/035zcJ98ItB74V4NbRJfr2sXOj7So50eE43M4IoUmqDduu0RF
tNxpOH/ZlrxHeAXihkacA4C9pOMP0S1wQwYNJwc/VgiE8d+drtQth2g7BfRbcu53
AukghhWM1j5ab+Z+1S4BLJhia+fC1rJnlau8h3b8LeRL4IGcQE/ty58nncVO9xuE
ss5Gcm84jY6viGvv2//THcVYWpET9ZcpMJaDNZr7RQc1efC+/yOHEgTM0f3AMuI4
VLA+Tm0wdsYIQwBBg0llYUEUFE/sL3+bDY/NrcO85sCg9N1raG8DTJU5RIPi0uSU
ka4cH5uFhxvm7rabWE4bFHHU50H8Gf35iK4QQbb2jZCk+lE6csfjgwBeejOPiHh6
e5PeInTsVb8GQ9wJT+f3LTMDGGG1JLbulSkC0JA5c+tdAkJQu7nug2fJ9Sw7Vwzz
hVWZy3qQWSzU8U0W1o6KVtcpD57Dt2ElYkjA13SNtB4E0rkO4vQsMSVYg0xITygw
+hsr8wWgLyrYy0qOc4Ds5UQlvtkhJk7FxaTJHeOHo/JYdNW7nKv+gjPfsQO6JQDc
HDt185yZHEE2SF9vsNDltPhwNe6ni3Fc9vwIWs0WB381viP/sy7zl0udEby+TSia
wwhSMbn2wqB+E3qMyyshwnMJIurANw5WWzpNgmo6qzBvshhKZQ/0kGBkgUtJsIs5
oOYw5sqqLjd/VkmV2XVjW8C1fR+fvRNAiDknoxEIX01qChSFpvtf+setY+p9+swd
KR2nO27ZNiOD6LSFQnmQAyABP6XS/VocHd7d+RP1ZYKOuhbocsetRB9Qtt8VaP7U
3hQwmaN94Pikz0lMc5SLKn0Jc5BFHzQbYlVQMVA/Xj8dxaHT+UK9u1iDHrdQUG7g
3aWLURpnlvn25+/0B6DUkbZS2e+GeGbJlo0UTTLI0R09OeXYvqFQJzfUrrVFrNFy
MCdOPDZBJXGcdCDngbpxJf5vWMLanO8bHdRqgeRuzdeoSz1RoYQTIP3qqfbVh1Z4
xL7INisoeZJRYz4dOgpifEKYyKUP0m41O6UQUjaFMCOC9FtlUmzuLaiMcTyVWx3I
zFOrgJdi+MT68dnlUJ4ayNaxAnqBpsmVzTlk1sTyoWRHnTTu48rElGPuyfjx5JeY
P4FG/eiz36qGt6Nar78mwChHWgMOjHGGJjykX5+mL42YwTeIcRYhEGk2SEYw+TDv
Fp+JF3ZYgQpNLU+TK3VYXcNbGStYkeda09IBK/hU0vPSO9Qa0WqL5bTcIX+88Yq6
XPxYjqDQ2v0Vo856L4uuvrqeBPfogHQkUSJIH6ElVpaKSZSUvqkhbOufgnZiZJ9g
D78fQyzVeKEuVZn3/CDDYF93GveSz7ZSSyJWOWCYimNuj/Y/9BWhXEH4BovT0onD
qabOXDBjiwWU4ZeqRp/3woHZZK9r/onXO1Agz9Qx2xLt5HYtUXieqSMDoITNuYFP
orCp/ycmhZDLfhU0dKlJff5ppTyNU2dGGTgWMmEEPsGVZyTMV6vOwEMlqflq9FBg
72UlOGU5Ist1xGLLqqy6RUjuXnUWe/6M/w+//f+e5dTItMbwGAd62sv5PdbCCsW3
Bu/yW9BiS/g9Jy2PklDaVF4B/xtD0/D0HqS+eHS1INN6STUs4aF2QkW9BIeUCcsx
3G4+rhn8vafiyRIsReaSTdcWIE6K3ToxwN7XCOtcxMc7Tf+FlCce2oUwSUF4WkBA
gXwZcDD0QfIVJJ9XczREhWEYua0P0kWhEZoTScUoJdC8/XczbE7m8OFCuil+J0ta
EQNNaiF+vz6Fvq9bndBr4jbykDxm2EIQWi+KBwaD1Hfelq8PhXXy7PkMxN/4Voki
926vxszEx1LmFtazMU7eiOnoTBY9UcDDi2nHcPeZ2MMT6vcly+ywSbMMxulH8xgY
vtWmKPiv6KyeeXjaSp75EDD/dsPzKjq3MFR1SXZ/3RCvWnQ6mi56d+OdgBXBFwUZ
/gfTzWi8jOdpf19cxK/e2dOuNEgDNYZLVelN+fF0Vd2s9Fc1ef8bb5EGyjQpL6oz
8X+2zrqAXTfbL/Vnv8OuffMWei8Ws5BG9xz2hkcmqgxrWa7nL3jNNeQ8NaAGFdqp
rBAvDH8tkkEWUYJK/k1C8cPxr3ypSJ0Y720kn2NxuTu7eJellGhcyGv91VCHLLPW
PycEnRznxe0noeufXbZUFSI5t1YUE204YvmoyBwVkX1y5KpHdVtJVgkvYzUHEGJB
/zKPK+gAMwsJ8YXTDxhYVWsE2gHQp5Vqp6CsPH7RdIq1SzJ0LeNuhN7VGAWx545f
/UN/RVD8kMBIT0kUn/AcqeFOHRIAvT1Ddk/i2pAhSnarQgwZ1o0d9FriJFGGIkZj
Z9lYLLnxYmGw0aHZ0+fOWBnaKPvG02xHH22pOFSggAykNnF0ZTocUzVFYH2ChTh8
1LOove1ORTRaZNPzzruD44MTmdN0I0UBCB9quhoRmo5UBlGB/zXoOSVebzr5PnBW
vPKCzSz1QcdAwJw2nwlJwwQ63lP/z0r99BNP7FejWfYf5Rvjf/lFnuhlK+VZr27Q
juu1cAdFGq2b6iSRXVa+pmcKhSar5z8Z5rLafokEv209qI/Gg9r1C9jqlaQb5Jbp
68pLGCrU5PZ9osDRe8CyLAVXzSuIazN5PRO5ryH9ELFqKUK///CtPk9rxqoREUr0
r8YAUVByTzNIqxpVdUh1lz758BmTmw4qyDEQKJu0BN5cL8+YnqsCAXNqRlpwS016
/VG+QxsoGXxo1sF7AmT0gfrp1Q+dMHpK90FmWggDrit+DSwdP0XclK7wp022JVo4
06b3HW6nkeNMHU2r7Mb1gSLWsC15hEPmKeQaJ5BZCsphrCcnBGc1IjG8qSAUugnk
a2FD4B6uV41t7u1Bi/s9RWqc6m6WPB1ZCZhaaUzra1+tcQErueH+1TZIzXjqZARK
feRa5Iqbb4RqeKT0qCdBSxUTcQd8m/qEcQl60J8pg1JtFVtDGtxBI+Iio1Nia1lZ
4OkLQIv0EZEUqdq56w3OrAWO04XechgwTbtjH/H3+6y9lxp89T+nF1LBB7RtNK8U
2G59nAyERm2F7XR0LOPMod1yWgWbyo4bLoB92Z4ZrkSPcQFTJyG9rm3laBbAXpMT
ZbVm8y6Z7XoV/hUTjvOlOfablNlXDdNQSG+4M85HwF3XfJxSVHBh78J7bieLX8Nk
WaPABqWVCF5b9ap4kBBD0vMYop8uSslGvCD5IEy7DdOhY621CNGgqcKrjyN/XLN+
OwsKLHvEtVv3524SqIEo0X6v+MrZ+jIveX/pO9a0E/MCTK477fpd3xk73XY3Fahi
iIfYm3M14QFoKcpTZ9ji9ztNXolVSStpgc53Q2G9hcJ1z0AOcOCjL3AXsiKgD2Qa
jO80rzFaT5m4RHpaTvRA1ppUJgBqLbUeAoM3yhb+WxyX84zo6ntu2mYHqMxleFOx
Rwt/opCpjooQ/KXg0x7P+a10aNt8Xt7RLa4OhFragjY06TV/IPVQhyuo4PtMjQ0i
Ti0Z9QrAxw+g1nBUha+K0Mu+HPAS9IRZmNoL4qmW3D48hJSHSM22VjEwbSbZ9GVG
9yMugdwN1Zn0YaUO3M6EGlc2Hk9oaNZsoXWZLrJni+IBBwM9Z9g+phtS4t/Sq9bY
WcDhYjEvs6fNQAJynYR9ZloZuW/rNWZVQJOoi4QIxOnkf5KHnInuv2rBqsd9DXeD
VnAw8AgicjCXK+GXtW1KQdWrXJD40CZESETdNjXlan+Ck/HeFv77to4TZ5Vm8a/S
2xQ1c3Jp/Go+6+ZMlsqmZMGJxSZ6EFEs/77EY0XgKwIZI/YWXZLLMULrXV1oAwv0
8C0Dq/LrmP4LNPdxbyB6p/aQyzk5hgUDIlsWvDp2TLzsXv+Nc/ep+fBKd4JY/HhX
UzYJ9li7S0kRq5bK93shNKjcYBmPBVBhf4af5WxxwUm7zptjUtFrnEput6bAwH/h
4YkO/0Qnak+rrE1lKCjhI0wio9MGuCXceckJmG1sSjOyhWkt4vAUkW19s+nUa/A3
pniLJINE6y3VlLrwL/9zXkRyAGqIail96zW7I03u8Og3VpYJBIcG5F1r9lmJMDZE
GyW2HglbB672S8XuS/oZG305jpNC/0IXSW7mW3OAsboMetPOdLTQRetf3rHXzyBE
dF5wemRcJJZBu8mIky95Pj5RpmY3xRIw5md5AH61Qt8mbCDwoaOpWYcNiXMhfDPR
mo1AKmylo2ZtHt33gkXBxkZuTxDpSx5P7a0lddBpSUXnwiwpZ5b2DFJaewdfRUma
5rsKNaDa/x4yDWSBAG87ptgTtfmtUwTMdz73CEo7hzmSIFf9c1mWPhI6RU+aNXcE
5X21XufM1znBQYPQzqu5SZlvRvgPPe0kXYCUnancqvA8TnhBAQmRtTRz8mKFABRh
wOI2GthWUAkKNfy5zuxgtHy0Zs+1tNZY8EWlwYSwZss1KGmOK38cwqlkgU1HuYFc
bvLJyy4nPwv9WL9TR+fgES6wFZu+R1Zg5pdciOct1fAxXu8aP9GTQb179k9H/f3s
h0NGC+yoe9Mx9T7OYD/uzbihsyh9J2Ju9l8VuCtVzaDurmRqNlJTuTdAXp06zb8P
aomB63Dy9FUAhvxRvoNY2F18SCk78JMqpVX/Q9/fW/2+q5l2uoXWktsxj4tY/xt7
SY52eVQEpFTIre++AsnVB9fvTA+l6ZecJKeceY0GrZsFV1X7itPUFAP3j/2TjeJU
nvktqDRkK1M/RgjYsfMrkmXW+4yLN1Vay8feQJX+XYN3Jesuc3IecQ5hGMf29Bn8
56pbyiwd90Fp2zYFTGn+8z7tC+7mk1yTRdqi306Etwrl1embm1aj/64J2tu3Aeww
VKSyK2xBcouxFW06LVeXJt6IxF5AmMG4mVFMTtayiGKNW3Qfd/JlQ+nGhWTy+GI6
mZKwx0KZA8ihpr7hs+mcznzmHodrPLmTmtX1VV1HDZ5LqZZkNSH3TJlG4S8ZEBpy
B5PyGilaFkQaJq7473/hE1WQ7eoFiZzA1LUD2MHeC0Z7OeapbTBow4uYAY/1d+b0
uC/1v2RC9/qZOG2P6GwrY5LnG/UomBS0hnjyu7y5Cz/OTa6w/bvL4P5MvHJSx0FN
xkbcZNdnwTtSvf5pB+l1CMb5ZS7gmKrV3eOEIEGYs7POSyMDbgpSedQNZm2dX8Hz
fAu4dgYwHXWEFASRvaFYjC0baUgEQyH0AYVsGbcnUnQXhzMyE5q8D/ad40wB2O8n
Un9tTbd/4cRMdkJsxtRc/Y/p/BQqHrrz7qcR4dGULO10lkyZGn+YXe+ZEEUEcQr6
iTPmTKjORt8NbTB1Jm28cE+Ana2iIkWPAEfEqqAw21s6e9QM5xHkmOJsfvbztBIu
d7hAB2xnb9UEPGIOt+rT+F+Df5xpYuhcmCPURrvW8RpVKCRrGS+2nHRU8cqtCRzG
oSHYLq45vB7SVRYehIYjDn0IBnHv5ju0c/hLoYLXBAsd/u/eKSi0Qev8hFbTGMEs
+ya6sMT/nnJ3TsLBvlWhmsxjkxdNqXapUsU7YNfczCQUWtPSI8oGCbT9MVmcSEby
+J548gQywJAHLrabYQVEHdQABVEGGv7W4L1yWN28Gmc9k+kSZLsX46GWNMsH2Ijx
QAuNxt4L5DNTHDcT70LnYcKgiQVmPor0iat2OLddeQimhT2L7ycTRMSg0wLEPFhE
Ilk5PHmo5xRWuXe1z42M5s/3LnigRK4Yi3eXimD93p/3uwqo1zlCzAlPVCgcIiK+
BooVz1m+2kyaV9cSvmOZTWNTiDIxenx/tPN1Be6TYeb3fn6JGazVXLgtsUKb1/p4
y+Z81ISzjWS+iYFgwlurTpm7jHRYxzfNK0hGjzg5/QeUfjy0NQNM+nha/cDOimNI
urm/6YS27hXYXHOiMFHy4k3SpGQDaACOa/QyYD9T5wFurIMFPVP29YKNc6cNIJkb
86XD+NaUlvHji5E/dNfcZInHspNIAAaX4iAClLTVxv1P4Riyu/fD5A3YviZX8JGf
6y9AYG/zLcxoX+ZdysymvBMhcyklhixwhHcpX9VykWiHqL6mfO9iUfDmk3a0cVF6
5DTiY2Oy0m6QrcN2j+33g5N4CTmKEBdQa9BUshm/d7SsBfXU4WsXJTFXx8u0ePAa
3PkFi8NkUWS9hIJhrY9X8GY8+pDS4BqWBaSXyJ68HnQ2TnenQnt67aLBnoodKZYZ
m5irPGWi0gP4c5AF19SMWkv8POTvW2an1/OSWsknLIU0ieeIje7zEw1Ks20v71V/
6Wu4aV6/5zduC0rhkHE4UtGqS9uabvgqymVoFSop/3DUdHyYS2rcr6BLuJt/Bd3e
XZLKItQX3+c26Sr3giRlzh6K1RBtkddGReag4/YAkG/NydTnduwRxbKWMmKXUumf
8zlNHSu/BISBpqNIWH7Qr6w2SKtgTFNOE4ThZA4plVwpXL7DYmUomCIXfTvTeHIs
43zwWsttJYR69Yctaem+j48vAM1tmkew+QCXuCirPaqA8JUKRcvCQgYPyG6ZOuTn
DGDGqNGbEa09Nam3hH8LBVnh/CZ75H3tc/2JLIwLVAWX5qWTK7lQzbvCamcq8m3r
Y1JWXsV5cTuc6lFXX/lDy/CW/ExjHlZ1GajMsl5a1SBNs4cNBsdcb4kM2dSCtkXL
/eAH0anpqc332QOkqwg5pjhcS8mH+SVNYHyOuLJXsxdfkx98v288bNcLjBq8aZEl
pXdH7uL8qZ1xqzIlKhAWWvyFxKh8S3Rs9DK0H2+doFgi1d7E6H/oMLMetBq6Rv93
nICsxGwhm8onKEcveutjvnaZYkB9Br8ZzrW6f49ls75IDEs4utz1Jzw1nkcl0Pon
e7UHMjlJlxS1B39uxXmdZNAAgYQajH1YIpNYOxOKWqLTV0f4yQHp3xmfGZmRZBgp
wjXEGGlG8hVUyneCl5FrVmjw8w7D7lXrgDqpr5W+VxOqIsmP7NJrKctLfT5YpO29
mENRgB6qCV7TafYy68olAD9SSRXMlAJ1wwL6rdyJ1c1rITwB4Ox+GYSLyX9F6pXK
wZqPmzr5gXgJ3IDEq29oF7WyGK6frYmWemZOfDU30ByqlQuyl2wvzOstPN/CBJWL
Cu+lhG3/6bhWT6uU9HPHytot/LpGC+D0pkWfZNsB5HFAf7kb6viRJHNlmAuSgC3X
gHztyjPU+5BRx6mG8xRM2f7MWUub00pgLCOAv87Sp8V0BmZMunP12NPLpksT5jRH
tujthkp3h38DOp1U8gwbnz8+AohSieDwPQvxiQU8WX0SXO0OyfZOWyWLkbPraDb6
YJlK0DKMAYzTPQIyDbSO9FQanL2ihDzBqSpNq/aYrRwN2XRsMAedkyjYuWpWdV9L
PFjk4Z7xWyD+yqKFvRngOO6d1fUZpsnsUdD8JbK8Cid64cMEoXCH1KU0hyHSsRBT
U3ZMbNjT8G4ocehEUCQRYwySMVF6hMUYdwNUbAhPqYykmRI2y4410uJCg8Pi2Z0t
JNlN7+YrHIcIrsfqiP6fhS9XL+c0jYp8ag5cyAoOET9cSBbLn4WKYgR7Ojym21kH
haQKY97h6K40tztjMT7WEAZ6TxMzP/f1nNiMJNM9oVV8S2W8oJ0wMhAE3uNkXban
KNIxGCVrzO1oxM9p+z4QcrRWGWsV3D6ub891lhSOGfNUeXKpvVcMDIZaaZqoJRGV
IOxqZn76GWRN+HZ7Hrw1Wd83saoDUquH2YkuoiQ0of9TC6lGKgNUb0no6N+yCMxU
mWG1tYEiJp7cFsoL8Bgn0O6ppMYObD4P0ngCJdHzpa3Znuyh+IrmeCEbHivorCpj
ZnJkds0dwZFZTTyllPE4CuuME39HU4ao+jxjUegale541F70BkE3KLKGjOZFyN+k
bVCp0nw4Heq+TRP2nSMfmL5uzRlAvkEhzQv/DM6E4du4ge91av4mQBaytaK/msfY
//WHsFl/QzAhFKEVX0Z+D/YSTx/YXDHbLy+pEYVRY8J13JY4ldnW5dt5DavyYrVW
fF6mOYO4jmuqyi05mgNsxl0mwQQiuwDhrODs5EH/hJ1TdFLfEDvJXznfmITE/wKX
/pU2c5PEDoEyVWGez3jcBCiXmclYziqfHU8unHCzeqw2XH9xpP639zXrk23TcLaK
XGoKtHsmIP5WNJ8jp9VRIJclKtvcQNOBqwLEtT9fw8mCARrTzECZVAx0qJ1KO9it
ZdBWgAQLNNhCkVloa5d0VSLkQyEzaAHEGZ4zxBJdXpyLumdCPAwgVFcmAEUjWhA0
DfcmWw6w+OTqc+nQDZw8Yo37AkspdSLFcaXIpvw4X4L6Kw1DpCO9RiAgxP5lj9B2
r6QoeF4Pc4YsSdyDYYSksv1AIATC03PnyK2EsuoZcpkQP7nfqdS/nQcqd+behLaL
Ga2gEHoDFzxxvNBb0kJG7zogUW9keQ8QNkiRWiiblhBpb6v+HGAHu0keiHiPHk++
Ck8EdJFAkkF//jyEP6kN/YYOzBNfYBc4e2iNlYU3SFd6WvLM3Pjy7aznTNw5yCaB
3eOc3y+qCa8MV/RCFK24Sua7x0iP1riOQTKCguplkC5jej24zRYC/Rz0nAwvc20v
Owp2oTdAtxb6dkk49x/GLaQMiFO1dXFxuKRgLilVSkDpyyVdExvOM03FuiqgnOEx
8qgznA1T9Z6BRyw0S+A6so7YaQi5ctwRNym3EixJiPg8daQVwBGbi65hvyw/w8j9
6telsJFY+7VbN0eZe7BBsXsozcHsDrOmB45c54DLFi5wQnzJ1ETsrPM23I/cUW+4
tXuMRRc/vQdY1bngMmjpqI6zQ9U8TolOGq3zmPHAALJO52Y2q+WrNTMSextc2R2Q
DWc2wln24h9HekoifqCGAYIFic+MP3uWsU5qN+GRJ7Ls6Eq+rQ+eJlbod9GfBD/Z
wOBFEjPlgi2pLjp7vzsAs5jc/ditcmvKBZ+ctn/OTacGP4iOWanyAKLl0f2Mquta
YnwlO3s432ZWGKz6Lg7a0TZWl8NefGj/crrzL76sFFiDxj2J0Q+ooOPqFL+Ogl+W
v4vWLcFjMAkMtLrp/rd1jvrHP1DSpa+YTL4n4jYYfu1uckTS3Y80OhyR5a0hxFn7
Vpwf+GQOYJAzkh22Z4E0M6QwpbTBWs3KuvDgbBva3HrlwDrYMcCnI5i3MFRNshr+
s+IytHvwIKNNR1eS//gAhgEL+ig0qxVEAYoCzuXSYiW6Z2EJ7OURSmhCFH3nk2Mb
JLnkth0C1imkL2OzczTf8KwkuKotLDYjclcqeiDHxb+quSMVMzEkfTC38suM4h92
Y81Il36JATcz+jh/AHV/ifFGCy2DgkTeB8PLXr86UOY8aZlQwf27FNij1sQixZ0Z
Y/HEK0bkqMlJ5Md93Ua0rCFLHjPbn/ntMk2ngI+HYH9H/kuOLKwV+aj1SNDf3OQi
lDQDE4L7wN6u7knmccZ0atcBNMQRpx7slJIAAgWalLoUNLbovVzQgUdcb5+z2tSt
ZmhoSeqG1IzAkFJDq3fjW++YWQan1WLN7Sdyr5pkb/zfEb4oWxKJXEN5BNz8yWlF
bg6fvhTYd45hJGTkS/Pd2oPaYt0+mhi9S/Ru7olDkDsVNbL8Pblv031d8VJSrAqP
TLYUY7y5vFYISDt3PlWJi08iQ3dco0oTfx4ubvvCg822JHsuGPLWiZTyqdQGPeQO
xSek0+8hsBkDp4mP8LjM5Iw6iqTa7Xzp9ox/g7kS8D1xjAKr+wl4cryLDTkMVP1a
vtZYwbCE2thQKU0sp1D2Gfh++vQ3BmUyHEWrhRQhzj7btccF1/Dljzl26EqvrcWB
lpEqZT07Y57b3eR7x5pnoXKzP4ODY84Un/2pVusGioANeXVS6U6gPrdKmjZkilph
Ddd1gsm3KTJ/TGT6nei53ilJ32UQiDdt6MsglMV4N9+FHctMvfSy99Kf+TQtQ1cq
wd+eZi/yRvYd/X+E71SzcDRyUUcoC55IyCawmwT3LCcJHfiHEfjPoybt7HLzZVpQ
cZtY+J6rjxI8409P22JnWapFs4tyIOQMGsPBsL9Wby13vDdOqQtM8Ya6M9npCxnA
HAutofuchXwWCW4I2GbmDzfyzxA6J/5/t5KqoEpBSqWgbcpf05DEjva4iXB5trcm
JzGtkIqpmFasombhJ1og4q524bGj/HlwgLSdeXAJ6kjqNMyYUamRzekm72d3T0sf
GnHlBV0cRRLmLaHOzoiLzA+bld540C63S3Cw+C0HJq3VgOMzyUBE8TEP8U4Ifdbd
0S32zg6DxHDvlo2lve/2pUx5nPbCQ8Oac6bkHPTOZeDQvlmT4SQ46wFoY5Io31Cb
IJgTe9qZW8AXp6CIkAxpU0TlCDPLnXl5poy/us2dJ5I3J3Aqu/HD74jkn/RLX82U
4xOgT0ncq8uxegQW9m9bNNmkVPvr2gzsYqMxim/VPJhYCP5J24RoEirDQ7ngGNmr
rPgmKx3Jncvzwb/UunOxV0+RKvlVU4JUJAbU0YG90oj/aYCZDfzEHPQK3OkotQma
3jIwLPn+DStqWUFFH6KddIUsokdTC7nk65E01mDi7ZoddDTBwKpJA4jNAA8kGEnZ
CT9vCtH7wczlybfCwQWzmpWV6Jlky5doNrmJo3SncJXnIDpBF7hozNT+cH50kbM+
o8JsLf8jvBsHlmjVl8mvDcU59L56qoRw+YK1K7w3DTk6+TceQ6kdfq9AhgjTPGEr
B/qupICC0N6iyo3X0Ruamkmf9kX8nl7fXFiHhoniRfxZnzzqj6kjiHxEGPBGpDWd
LoDh+Tr8GVCd8cb6bVdeMGXGUsYKaKezd4pW9MQisi50wNALT0JksZ9LqJGI9is5
WnbCxnRi/QAFypibZDJJczB9KSU/Yx0wZMQLoliDFkjM8MhV/42iqx/OIDnAAAJM
PRF74ijaLdcB//4M5+W3QqnLUD+ZrcwfaXSMbuywzD1vkVukjtMac9VNVRV4OSk/
LewL+8302Hb6clAkYvdAD445pGwwL97+xCpHs+jB6vDlSKb3+RU/1J8RORz+bDAq
OCJv/aklD/aJ/FZY9nBcoUI4lBsjldnlRNTVecpQoWxHg9UjB8Im0rZjlXJdtAb0
qnPZbF75NPWH5Z5AoYM6K4inuPvup/1RBPvPoxoAaNvKn4Nem5oWxxMJUVz6n/vj
FeMXbyfa85tTa/hfGRIodt7NkOJ64en3XU6XE25rMp/d3gATeCvf0LBwR5IakC4B
qi4b6tAx3BDuo5KcsWr/QIbaIPlS5h/DJtLlck0zBAIjMSRtwoNz8PzVM9oGDNln
GKmj5ed/A3vXY2KiMsJQW3kY+AKF8Uv3VXxfYdbbnHqtV+m3+qzclgJjERZUKK3H
NwdRsN27FFMZDBx1aUW+Qr+8eBWNwnT27mH2EDA0XShAMYHr0EtcqQKTQ841I/Sh
hwki5pZ6+uYdDVCPCbIXhCnRzy6DcebCayln6x8iRKmVm3OiJ4UVuYdkc0eGNYzo
Ti5dt4aVURCDnfZTzb0aC9+xN+Cel3doNZ1DZLtvVOv5j1tZv4+WrX/qo4/Q2M2c
6bkZCbqXqBCCXC70CZbk0uwCSCEGdhVihd43C8jY5TzgTOVMfOvjlWDlL5jeKb6r
R9L/TxD49TU0a+/JVQbC/2NPa+Id5MoIp7IBpFzIhNrL9RLYxepYa0NYmlS6ekD3
wTMPQe7R+7APx/NZ14uL0hRq9bgBKN0tRp+R1eGgOBLfylOak+CsCq9qrp8F3sRO
FuvJm11JceKGe2rNuVdhjEEUZeXztt/OoRdftzaDunFkN+ZeYlI6dS9FTVPHQhoV
gZN56uLG0VPEmd/xOWJzE9jfc6gOIM4ccHxv0pta8c8oLSIim8ZMbTzr0WyotkDx
ixHJfpVHZ+C6LGO7hWOweMvxluCpbbvKrkHeKDVQByO7hMy4uSNR1HVMXLQ1CYI0
p9hn0BtowlHgpon/S2mEaamfBoomkvy/FBmn4cGaPryhGy1dWpw6YCgwp0IoCz6u
Xvz5+7qjtIuKkwd1kksUlRuOB/b/nA6/I8c3B1I2GzY9ex4d/wTHfvUCaPBjK22p
cK3R/lmEe6xdjHf/LY5ZOYDGjbeu0s04GfnH5qeqD+AgkyhRHvuI7wuYKi5jZM7U
0f4Az9VoYhBrxi4sZAYihlud7XMn3Hjf882bR74ZPe9aeiH2e+GZJcClAizALhe8
KZ94lMpFuLtMs2J6NlCq+v7EOrG14unEQWkZPGJeuUbchZ3+T9BvpWMv711LkoYs
WnzM3b9fI0Vh4PTSRDLFuKg5b8YAuGxbD7vmHG/aJn4oD9pkZF9mm8sxE0F6Arf4
byuaTHI0to+9jYQh1rIV8zwvLMMqfpVouW9Jk26oxfLrHP1sXkbdAqqGfAmZOLUq
cBSxHXbVokKwcsw9Jf8Rd2E4LvBnaXEl4gMiaeSwNKlfswD3KSefeBoaKiXu9T+H
HIb+qdTv99wKpfHDnC7y+H+jNt3yHcVRA6+Mo/fkofEXH1Li6h3eiKA3WM3kOrig
NJf5FS0u5TZ/QZ4RV6ODMTa/VaiAGLe51414H6YCnFVrGc7EjJKRApXEPJ61zvlg
/mIJ2OkfbpU0/uEAKOPUWyPc8LdzqEbZW6BbUC+qiKRHfnSvyQkodRhvxUCLg0Yz
ipCKx2P+wZl2J+Bre5rbRe3tBV7LS+Vh/aoOwkJJjjIMyufeVNaUN9vIzIEOQEtz
7GcFerFw4ykyXUwLbYRDnKzddtycY94Ozo4DG2F9AtJgiFuoBd9oFuvSb05M+/Om
qHpBOwIG8TEPXt497S+nMroFaIvklRdjpN7gTCk+jJ9p9m7KvfJjk6oRM6/k7daT
E1/NHJ1ykFVGXucX1WIaPa8NiLWuN3NCO8FXX2JaaNh3pFQuZXdPHjAhRa+lT3Cc
g5vJbXrtSFs22bEnSY79yN+f0DFmTy1JFfB3T8fB57nJihs8iy5Z2n5HwoOq42I3
snU57f8zzHrvlzZDbQe2fmPTAaQUdeXOLufwxMQiNm/uLlo2DaaprGFtcUd3NtYc
9vHBkPRzNitR+4uRVD3NUaxn3NQPxXohMYZNUMJYRxLeJPcFiHaudeDk2KJGmH6Z
NW85aZLCB4jQ3O3JByvkZeyLGopuDQqabmI6b3fy8XSf2rSp7BcwqI1TQOftuXKM
iLRuhSJWfM0WWljsrL/khG88cMLBEZnjpK8yDsZW0PG6m7/XisQkwdgADYZKuLsg
c/VuXpUgtrpWn3z1XDfdpSoceWW6EX9pPL7qYxFo35QWstvyBjen7u5shgbuUubq
JCs2stev20WHolz1Xx7yb6GKqMuvgDT4MusD3VesFJVAH9WG4LmeLb7sQvle7KXW
zkydmoDUCfQ6u2rgGmBA+7jP2FtjTXp7MDnG/5uaZhIDZjP7DGri/Bk+vBQlh/y7
7nFgTLaqFfIu/b20uLewnLZ+oWqCvLcA7LAb+E0tvVJEj/4WPbcF3qbsoOpXGbch
KhC2IgRPtKwSSlLfp9cTY3KMCnmT3hsahe27Qk2JfR/yky7CMPthMgftzk0+uH8G
z+E8VfuJc26tpD3PUuQQahPNe/+v8zTavavdk10JiaBmHqk41CbhO6INLsjOoMeh
0gAp9f3KAqIWRkEyFwYC0CdskGk2RdoubdYTymcg05jUa7QGyDfIsA088n1tmLkN
8ul+BpCcNaaEyCpxHIVOPwizGAsAMvkTxyHZuXopRxiLbxapYeG9+nAmBa64LkSQ
hWIK9ORzBiQdQI6H4z3Nj0nc26yDIG7K2qt9AnnE6L0sKZFwxhQYWg335CnSqhyZ
6PE70XaEAEMV/zDZ+mMndpAqUcF2HRVKB+7XYZIRSrVP3V8gitItvCq5zxid/m0q
9J27rZrmNgujNLA+zGulBtgVyPh94KVkuIjwBnZrCJqyF02MG8tWFtlZ1NshRFh4
O15Vc3L8gQmQno+pqvgz4JKk5OGmc97I72PYeceEMKkj240EP/sdmgsgZFP77aCG
vDv9006fSzoMS9wiYTJqnpjhO/SkPnI3YMudKg72TvvhzXAIAJagCCSAAxfMUYQK
sz98kQ0cIwanZ8iJUnGO1LnYgbgKQZvbce3+C7PkANP+znWtJfyZM1MMk7RaSlw3
xaTDDvLcFxoRtXnl77GAN9IcXKHZsyx35A3f97M6GH2cktWRkhvQNMzv2ztbRzzj
CSO3nNacXcg7ni1Es8J2nqrU0Qm0ODdSoVfowVOJsSsss00ewijoZB2Cla7CpVyO
nTiWU7YvAMi/VgWk7j/aEO5AKvkDqsDxm4URqU3skFe3aTfAhzA4XVIAoQnAl91r
+o7XoTmwiIhs8i7KTH1/K4bOnjN369197AQyM/bFjEqUUUoWoPJa8OSo3tWvjil6
r1lLqdETzIfvjSO+FhjbRUf+2MWf3d/34Nys2/mXqEtcCip9geOPP52qtSClObcL
lAJCyshBkvE6zc6t3ssjz6y1hieLCeglFhrrkEXRT62J/T9+0Purwav8V/owTfRS
mLfpQnIwzMIS/xLYQ98oD/RKvgIzkPnt1249zGclSLGbtk3PyLDnYWaVLT8MQpzm
52XyBreqaaNq1E3ypHcD8mcESHiN3l55hvBe6hb7b6EJapLQBlxsciGTYCMEdrn0
lc9FDcYUOQ6ogfvX5Zdu85rRE2FthCInjPk9hhx1Y+fGZa8orDXRzRMzyCxOl/RH
Yo3lbRxB/iFoRmuMZpwWTKEDxt8TB7nu3MnRHLXQ3X+rS1JMsiyD+8UnZzX+ceoR
4/iFjnnjkXRhQy28KOgeltYlMw+J7d8yiTXqw8ppkhel5JCs9T5mc9mPjKvcwX1G
3IwpxhLpIh0h5RYhE2DevlAZTzxdxZCMejBMq6rwuWaAxPXvZfRdZelkYb60aBsi
LApY894IJRd1A/ChUintBJJJUqeDqebJwYVSbA121N65VfRBlojCYu5r5ebJ6Nw7
CC911l6CNrCQUz0jSEywfz4w8LVyHP8TLw/yA837zC4KsEOtPcJ/vukkQ+MLgRK/
22kYhrdmQosN3+AeAUT5h3NaFkeIObuVQbRfVXUgPh80sBGonBrFHYCy3XXIx16h
oH0tiu1JE0dNLQ7JtDnOEoC07Ywfdef7hfF1137F2EJcpQVnviC4+rZyLCHVLRGd
CYzAv5oYEzeszvS/te+1etGeSU6WF6/B7kwm+bVXBhxetR+MEcWDQbUdEHGHo3o5
V4Vl+1nSFLS4St+EsZS9Tjtkp+w/SpKSgJ5GjwPG3X8s/Z679LSsXw4vILbfAz5R
4LY9swAol1zrYSrbpqH69VWvP3P3A5+6Kx16amFoUlBVjNtSHVXJRopl28aunGgu
zxomArDuSafPmvAiD9Nvn7f9NiDxp/Bf3R+h8vJ2mjKBvzdrRybl2BkjSud4GluV
85S5KYt8lO6O/gAaemO2l4FFoGPl0LhbfVM4PQaBNnAYb1k9E5l0uXsoqIvQvHkg
ecKGsiBe6iK+1LDdJCseciICkxHm7oDMeN+Jjyw1NCi8q/Io/rleKc2eBw+qJySx
xWtFhamtU0HcgPkH52WQERaA5XKP0Yo91gcqPvPUSDOqYCQ/Pn8ywaC6OAchGJVw
hlj/A59QwkmSEGa4oYQjSOiIpUAwcHA1tmSUt1IBQV5VmvGp30SwnHXygFHVnJbH
j7BXH68qCc3VsDhw5+RWd2gGnBcrpQHBmBDOJoM//OAnGBYCQ0E7RCrS3vaephiA
n3WG5iDdKWn5y7RmKbP1PVNkG/PbRei2phsL8A++uQdatu1iOaEc6q7g3TBEFc3Q
AN0uEnIsJ/4nk84IDpazhy+CvKQl5Htwk/yJqzUae7WF5bYLOyBvNuNgOIyIS/vv
/xobyccgIKpL1StG+RjZLndD9R9a7JP3AwzwDiJb7EtShT7xdP0i/w/L2PTCyqRs
YUoBy75kQ1D4Tze+KIy+SCNhsC2txqoOVxk/LhJtP+9lB16HjMVueBh6qHbe/PNV
yiUQPpXe7l6GhweA1eM6EWbCHJZMR/IbaYj7nQu8siF4p4NCZ1iogz+Khh38l18L
S4d41b0f2VaIsinl5SCN4Ljilja5GVEHtZ3iuGucfMqMRO03G+AsaX6Mz8ZimfwD
ee02ws+/YrMdyWgIiHG5RBtuU9ZxSlYrXW++HavJGXOTTVxT5ltJcv5QH7O5bT7g
9E0k2l4LFPsMFQqNfzU0wVXsa14po/eC48id05YjRC1BoivG/4RnE7s1C3gbhfjY
Yr/l/2xn1keHxiljQKL73qMxlRsL2AuIWQCD1TaqFXOStZjQnLNatxjhL4vtmpOH
h4wg+5rkDBVS8EWA5eg4+9vVPgg97ac58tkS2G+nW0kLokKH3yxbl2Y8T6ae6vEn
9vS3vjLulOfkeVHky3GGHfppZdms+YC5IFwn8TbX/MzOprIBil5bZj/BOOHEgDWD
EyC5w0jGu0wsay0O+v1uiqCbBeBusa8A4/MhMwvBosUR/nTYXq7Ait4O0dGbJu2T
JLzOhoe0GbjBAPfmPx8jQsaSzlPfEu2KDPEmjPI9CI2afeb/LlKaJKmvqB+llCWs
Kvsa8V/DRMM7ZoQ8RbiDyZeqwIYad01CqKr3Fyb4YHLg44PBk/hliid7ojn4+NN0
BBCudlWY7Bgfr2q/k8Y2nOCqlVxN7Jf8/3a5rnxEUNvyi+uXbSrFSfD2esgsCLv/
ApgowfG9EAnJO5CasIO4twaa0gGtCL3RM9U+feZkobWaX6STC1co53iAS+1qNJBc
qz8q9hO6r+nrFG6UaKEHJeN115nJvMSMZ5mclhRV1Jhb1MuGYFXMuy3nzJbMhIrm
FATa5A+Y012MgGXeouDHPRPNSxWwC/FfLjeEgUjBr3iQhEif6J+nnV3BVO5zClK2
Mey0XnL6SvPW+oz8vetYgQDgDvDf7hNSUQty7njWc4F6Sx5MMQLY6tjNApEgR2lS
+kmLmE0u4E5wOWkbPzp47hsUfBZJTcMGMkNhARSy0pIn0xWApc+cAICo6Lp8FvB/
tHEZUZoDUiiyK320UPxQbBFsEZj3FsMx/XJtP2aOVcz/fFbwR5zDVtwHDccfXVEv
mw2qE/LoxoIvSndCN9iBCrxRkcDM6tdFY6yyD1/DZZTaDaSRdCsjPOoIUp7EXHlh
h2jjghUqdc2aycAL+PI4UPiFuNYzgFZ9BfHrfEltFGXOy4hgOxqWC5E4MurSlsCC
Eo3k8F4RtIqdUDJoCWIPUtlGq/yHqnVmQ/P32wiFWN5Jt/FTVwQe4H4+vWD2ItSq
HRpRT1aKRDPw0Y5VHTdhRBrc6Ap320AN5qNUaIusn14+jScxGGUBF53wVe6Ugavo
CVUJ+whpOcCFZIepSFx/InEFYYzwLRH3A7rZg3Lmd7ppVkODV2j4f4y2vVbm+wLz
UV29skUS/4yxorBwYcrm5mzE5BNMkdIfOUxU20kJlToQIzpE3o9IA7YwIlEFQ5Hb
WYXqN7O2OfMWmzly9CHO++EhNLJbbieyy7/aeCybIMK1p6n0rYDqmv6g1hvuVBSz
Dkdw7akqOggWpLqOswuBsBzf6uwyAvWaNIveUzBz1ezxp2kzLp94vdaMLTXU76dM
ml8HErbZJN4xdqhbHvrWecKychh1ZhcvKEB9C4dUKetw74cW9daImvOdPcu9PIRa
iKX4IUZrzlxQ8PXtQRzKRBmcjVYn8zKOhmdwuovlO23zSFdkdk4uBZ9oGQZ5yrvN
ZE2p6VMWDV01SEwJTAsvOrh4VSStrd/wMOwt93j5iTu8KvDDz8draJMPzpYvQQ98
/4ZYS3IpxsQmeAHg1pNSa5E00/t5YKefNlyHCQj7ewi/gSIx+b3QbBAGUUJ+Vs0z
qEqNjk9G+pw4YEBUU4FW4vzxIhsl1ERkePN7XTlPQQhehAhVouEOHMs5kfhJvvzY
CkAKAMPNowhI/V9SgHsdL/vrwDd8vPZrwAi2gIgPwJ3QPV637LE674OmRii75p0E
sgSmzkaOnehqrZsp9V8nyGYYNboWxeyViKJNM8F4MDb8ikkydfW1qtL1pBe5wQLh
mzzf4KNaM1I0+90yItKHnOlhmNH0V8/621+KZ2RKTckzRb7I5R2hg3FRnceF/xws
de3Z/q0gsqLCt52mexiJr0222oA7HKFcCAUoqGlFPZo3vZyBc2AI0ACRw3QgKbF/
czoOQ9XvYzDYhpsv8IKU4F7it7W1381mSPzToRIPAH0s9U1Wb3Q1JgnAaXkRZgim
8yADBsk2vuXV9V/z81ZDWgPxmLHMqZtt+W7PxbFEPg+F+Ny9JH4xVYO9Ptr/i2GE
XpLf7crUe3GAEs1b8OjnCBaEzvpZG2QboadOHZnAj0+BklqN08/S+Q6ePgzfyZBc
PPKCPcH7A3KpF4lKGsud4Iq4P2km2GkKqkdkkVaXk1yYJKyf+NZsouRaaEfBCzke
XrGyCDHCYwq82N98dchOzwHDAV7BMEk9QDwfc9tI677oNAyByI200iSfBp5nE6bM
Ii40izqdmK1vU//nmwekp+v/a2R3Jr6nsISJhbXS9eVAPzqmsagM75qokD8iEiiB
wn0YIrEbnUI2D3grAhsFFCy4KpnB4/crE+Fl/2IFaXSu272WwA/8JEIG2vN9SH2n
ZlunbnkzWGBKlidPOpIWLa/tlfLIuq2PhYkqH7ZnmZ9sdtuqF9kf9f5fozV5DCLF
2H1unMzWCwEbwMEMlhj79nHh+oJJP0PQLKBueiXWf0b2dF1e4QAroX1aj/VaCFAq
NLsm6ggySFXV/Ckmc01xa55mBxI4sR/0SuwpWQ1zyPmFUQGQBP0B3Q4LRINxbBlw
NGqA5BPNeZ9XqyuMPxisN+RVDgrTAa+luZsaebArrVG6TYjQjjHVLUep+sa385wH
EaVlHV92HqurGD8ewlu0bdgnbZnEZkEhGJF2qHsKpFolURvq4Xr5PQAS/1pv0i8N
rhqsQxr8eWxOKoTNWjBJpDP/gqy6H34m54pQktyK26UylE6oUhlHQWIxmqtskJu9
sDjBP5gxdAA+7SY6j8S/nGECG+f5TdgE824yZcE6UTa37jqSRymk+fZ+xw/p8Pv9
D6S6UitzS9O70KYIe/2DBIZ8UV036yUpDfsAaIbOoC0oYCJb1UTDAcXefTZXZ6fN
z2uDoVTEI0+SKI14atd6UQ73jtQZaaE8E+wgXM5uMF7aqh/gohxIctbugbKm6M7v
wKvsq2Km5332rMDelbLnIhaT56DIbhaJoi1/b52DI5zDTfC4lRniJkW+JH+77HkP
T5R2TSv+blZSr8AX6GaZthOAeDAwYyp8ocDQ1MpVMKFzCr2jckp6HDPo0EkgenGt
nzhFgSQJ7j+7ZzBopSBW9xqP7NP6gjHlQcXDdXdQexi6LxQ9R+ltZo2uZmLB+sh4
k8cZkV4aLPECImlo90liQiXRbcymYqYwnX2SwxR/xzAp0EtoAVWYLBGJD0lFHZ1y
VrOx7VAyHkSPUe6/Myk2h0c2JUYV6e8eGtLsIJmGleeZcaByTawq0XUNAO63DLv0
On3IZ/o1qcN2Gdc0VR7mSGzKFrJXl9aCJHLLmWoZ+gi68K6N1zCR7qm1eOdr7jFg
rQ1l4CBn4CT5/zhoHEMa35aFP40+11BFtRZYa/8UjQdtdfCZdLKtIe1/B5j5V/lP
FvBW3G5IQ6ZhpKmaEzlcLYm7UiWXgSHbYVPQsqKtGgE9V5fNZ+s7mODKAYbMW58O
ce14qCsJ569/mpBO5tZG9fj+ZI7P1+wu3DEtuLwjXvkg8CBANhPFIF8bxVDcnhaK
0NEyOb2luHmJMYnGyCRe6DHSvNN15jcUY1+mG6euabTKSNcHGEZ04nkvopOE8aJZ
/39kUoYxBoJxPqX9+6BzEhSRzFIt5+wTqpilJKYD6UluhAX0v1P3Ibr+8nbL3yS/
UGQae/6O862XfnOSPIQHryiduNkFxDaVusWXGvdA9QlYUlA6a5f65tavP14QJ6Ce
CSTm+CYbKp1JoBQ3H17/814c8oJmw5hYoGZ+HIK2C2eG/3TN3GGEbrsut/J8PoSS
o2XUHKpDxSCyf3J/uZ5JMTnc/IBCoCXs3JiUNemREr5KF0vZx4dMkiOSuaqzRS+T
pmkpalqontewS2mqiJVW/CIu+39WgZV4FrpEekuxjTHRHitgIoK0pQNIH+GirvrW
NDEgJ4nmFq8SdFGiAmbl5xrqCT/3MY923qY2o4RZAZdUMYs/QCaeIWaJEgJYy5b1
vUxcDVmD7OFEkV9t8ataULzlbwlbBjCNHGS6E48HhypqT3qasctrW9z1QvsnVoMR
gOhb62uX9Xol+LjFnvW0Mg1jG9RYjrZ7q7Nw+KLTM/dxSyTDPCRP4Q8Ei5LvnBm5
c7mw7OSCPMAPLnmJVoeHuIU359VIp58F9PBT6knaSDP0rfhPMS9yCyXclKNI7tpE
MUOSUX6u69lr8/P5oAUpzCWJs9JI4sdhx5rA37H/Mz33hiI2fw7HhA3ZBTNuuKbP
JrTKF8c2TuMZlMXvdnw9LVE+bm9yzAUrMXRmLWgA0xfvuiw6gbbcckIrKNTp3r0d
5HlI3RXVfpdfbC7GqhuJ6dJUfX1obmtthqhfcTe+C6cQqPjVMPvtFTt6munK/KR7
qgk0nBDyrkcl87SynJgYNa9cgm8DrRXa78DGg28HfYAlU1QkmJC5TKp7wlUdBUEF
rsQxM9jKlf6R88Rnq9CfAX1Vhf7HXDhz77adNBGtoE19q6q//DdKzSS5wPGgDTtT
+196zjpUyNxCEJ2HXKidILgmPMkxCdESzb89eMHNpkZEoySRrnQKMlF+UfvCGXCn
luBqlCpkYvKztK2TbK0q/JJ10jTnDdhSIofx1yW6xsaWyvg8wl+f3RjB5NGaK/dQ
X7azYtMO74mIaFRmcXg11dEZPlJc1fDBxi4xCA56P3+EQfGLaDlQThKcachpHBoA
Bq32zwQlhhzA1c9DZoF5Hb/31vJHGGtaKv49U8tWXpxDViFIIEeiZl6cPI0VRrsI
+QcgntYmW47SG6cA7FYKaO+EATpXclngGLAVrEK8gOZLIrqcq3LA6yZ/SkpM73KS
U9txynhyVo7nMKkbQ6L6exJ2+mFbNi2qRodV3W2krwU0WfeTxiLMO3hlvLCcWOL6
QeStNBU/Ly63XJfHJzIc8hTsujCO3LsNTjfs0vEgYCR7M+sx4mgmUCt/jORtgON3
kAbLUfpkn3vYJQfceEfOOMuEsOzkmllpTbwalN0EDzSUHOnHko4MsfeaeplhruzN
NbrF6cVM347qmNAkZU+B6RH5IaVZny3JCuv8ylGuYREFa60inZOBbbYeYHom7CdE
vKbDfNd0jaPlhQ4MuJfUWC2L12YxBSZrXosDiRffKL1fIiMJlTZ+ZTOlz/pYXQ0o
LOMtFWD3q7oZzGBOJxqt8LZRTiKOfPgfAuujRIZ4LtV6lm3GnAVmK06K61ZXh0KS
fJrh//CuD2zA78Qg3hJBoqXDPakpxml7Ca4XTBLIHL56xKM4G+cADD7JZY/mz3LU
6lX24bvYYvVUyi/KQgGxyKMzAifHxH2TixjYpVHEL07rIijaoydS/2SNwIqr7ot5
fqtxQrAdfz5VtUyCggbkWu0IB+3L3mLULty1rmQoIpSEuhiUo62JOXu+sMlTtCxA
m3R9sc88M6U0D2cjrZgvOgkxsUag8GiL2+o0ZWrv1eJLD2ChhO4AOxXnODtP2D6C
chvK64dhIxL5xROopM3Ml1GyL8C/NfRH4D9OD2zTb4Y3ZKHAmv6opicJ7yTzGlTk
FES6RQUMQFaNYfwQAnBJAhuW3sDkQyJF3fy6BzQJurHyVhLfTuRZE19R3wAl4wY3
ig9ZxAecTWKoo6c+EGFwnd/PcGN4xhH2P0Tb8nzRsGZSv+BMxXiBfYd8QAmX/yjx
jpLLALzVQHTzRZ6dQYOPaA9AVDlMiKs5JZOzknibjPx7aSY2xGGmd1fTETpnQeHS
3Bb2UrtGfSNmcFlYmDRQNRYTCawwCA0m336sQyZdysaX1df4ZP8TTbLM60U2Zc9F
fZJ/Fm6FGbt5x0W+zxJnXCMtoc46JeujF7LqIEOvBlrMcJDY+IcGvO5LUIx9+bq+
9rMXNasBpyRcK06RYVzE8CooN5kMjkIExfaML3PHrFoQhd/A7XasIeBaKJri9EoT
6VrYTzH4HNbOop0lBdo66vgi5HMf1/EmUD1LUJIjubWDetujSJXmtC6X7mkF8zJ4
FZnygI17f9qrPzzy5C9JRs/fQnWrciS01o2TC8McO1YF1yee05hxDm7m8FqGoU2M
ocESFOedrsmH3D58hr8r4L30lXcei0VDlg/gFp96ml56FK3sYsvJNvNaKtkQKWRF
5lAbo4812iow+4MJaCToIU4mig15hl4lM2G//CPVz5b26Di0sjIVWM4rp2Sj8fnj
5d8mIQfB8+psiWl9ll48Yd3oqQNwTNKf+yZKXUa8F8bh92PzbC2LY7bwFkPf8Oro
xX50sagMGDLF0iBUVF0rIEc+onO6C+K0C9j8gYT1fuZCYb5a71OadQcxhuok/I56
Yd3AA/cEHCHf1eJ15IbDS/7ZWeHILKx9MGfxjrWpgBc8qkzF4I6BDDf03GDcU+YW
wvi+yYVEnGR8OlaMQpGjAgxAo/UsPcYYJrJCo63/v+a8igejRDxodiU/DcGDgHzb
uRlLHTqbba+2a7pjnu/IpizlCZ5ysAqd1cp3SES+2NfhemIb0yllGipXWO+onR2m
SACiK82WdWVM/w3E/2vXpIAgTl3gu4JjWHTcWFKwP6O7y+YQrGh0GNwpk4aL2+zw
xU7d1aWIcDwRVGveaofSZolrGvB27nQG4Ul7y6xFxPViZ0S2slapBkFxI3c5t2CS
i5ji39OinsVxGOu272oCnXiY5tw7h7pi6AlSDnJ4Zm24rDdCxFnjT5JqDOsBu2pN
NvicJ2J3TOVMtvY7FP2zQKHS2bpptJ8dYPfRGAiY9M6DBOKVh1WHyI1lR4l3RlR+
IEaleaREezgnfsPK1MSjJASQDMRie8OA+GVnw7wb3qzYrxQwXQiy/Lh6qcq6cVgY
GmAN4dSUuX6G9GOuH+8Eaqsv4+nbqwcB/HliMBn63sfxiSIn0nNic5HjeJBZ+McP
3hXzZRT+znExZxJybUhg7xG9t5kS/56gcpquhzj7G/1DvPv3wexHMgdUdJPBNBM8
Z6HKRPYe0Yt3+jUSpt5SjPR8/Zqk3wGCr61sx/9qf3OR+e6yF8gjALRWGPdhNy/3
Ncpr4jkl5yKl5WCgCp31gqehOoyE2y8Zd8Dq5o3ozrPOqxbkGG0RPfhvmGBK3krQ
Lukrjcnk1lYGRgOQ5ClHpHXZVfiJd7kQb4yh30jNhEhhnS+v2WyDRUXXHu+n5gvX
KxyGb9OFAwLyThQgelSxawJmD9FUilkllAlO2I//bkhGEpGBAkVrtaOSvu/eiSES
slsZpap826bEAUwV/8VYxme5XZEkM4AabtBHVo/WUBxvq7XvHkFtl4GzgGbLwHRc
ZpDXEG4hH4mNIWjZR25CuwZr0asclMnpSwIf62xPp4CboT6WNxsr1NTV3J6KrtEY
IKk1jfNtqE7l2Pp6sjDqI1KinWpKAUV6yAbsJ+JF0C3U/YMlKqDh/du7gP3KAKf+
XsQ22l6Rfwu11nz2lUp9XBbyOxHN6ZQ0PTpwbbUoMfvKAEoK6Dmx+eyH72qf3kLQ
e5WP7EHm2/B8FnhyZTPoXbaEf50P8fE5UaQWLRzZ03SoJO4lxLZSaoqRhpiKs6d/
Q1cSPWmtJSsfh7cMgZDZ5sSnm/AqdXkZFylePwVcx81Ujkdm9sNG5JegSYv7tI/w
gZT9ev0YxlLBo+Vg/tTwA3C1PEwmmO67t1CWpXnmRrng+ugCBKV1XnAsG2xPklvj
7YxnuUW9akcgSSz3jdrcDo9SZWXrBzQnoA0ATfHs4R7zIWWih3zTbw/v3PeRh5G9
D6LJ5mk2NZ3LdskBbNEafRwAXv5HCcUgrFZn1gdnHF74vtsZnJy2SYx/zFVFyPcA
D3mHIswdFYv8EZAa9gwRpcpNM9gVg8HK0ggCeJScT6uZOH59z1R0H9Vo8MVgv8YB
VSPnpuTvAZzIk0IBAPL7qXczPqwLeDoQ5aeFDMdkoRcsLm2IJDBSaHku4S/N801i
98fUElmKNzvnZKCi9ynV6ZC4L5y1veqwMNaCQsjuDExNTb+tWsRjbWvifu7FYqIz
o5OOVl4mswmckgcEQlxG/OguugTbU2JWewOKnSa9DKcfSij0cikDqv4mBJ5bmJMs
gvqOCUKKzAyianzgW389PEeHbnxl+/ZaLz5EbOqgNn1zAWWB52qgbdGHsFrUr3Ty
DOz+2RsHZqOj53Z0vn60rJQRjbe33rjlrY6hNWD8WhqYBLWQ8vWxc9mRRxWoB5Vh
SWSjv1RE/7zCDn+Gd+G6dAs52nN0h5G4Ict/chA3FmIhFuDOYjqFAnDkEuMMM2TN
CdvBeCIONRAPd3UvG8h2EOcQ9ZVKFcd2i6b74brWO1Yu452UNLs6o8pTN9kPq0nd
b/O+dgD5t6AMb8z99uO5s7+0PVCbwOwhFOQAtRk8HDx2Ph6e6ubPTNT/npIgO/u4
uHLeCjy5JeBlbJ6xYLnPDxJvyAJkXnpOmKXN6tlkKNo8LRTKN4wbyZA2ryPS7DUQ
r2VvegWjZRj6YHMB1lageiTDuqQ6M2jZ8WqkOzShrYLj+1zFEm280SeOdNaVcRAE
bFIXkc7n0Tu0QrLDPMtLW32ApTSb7w2bql4UTz39qJ13lQ3S8GesHJZHF3HjjMPT
VdqNmlOOJFH04KCrWCYHajWbLmQ0m5hSzVNpho6mY/4Ps4ZT0Ku0rMKReXKDhBv7
7BRleYLNo06knbK+G7UqVqjPc9SvdoKN/wpCR2+2OIOi/jLreqIHVEq0KKB8ixM0
kV6vbKvIsJBoE84vYnqPO3drpXR5s62NcQPyza5Ay1YP/kucsrfL2vAF/i7Lxi/H
JnAJRl/PXLz3ZvIOxBcu+akaM8oQ65Ji8rkQtbh2sMWThEX3NPYkNwteiWCS3hz4
8bi8HtCA3VyLzorWmhkB7NqlADI5yFB5B8hSJIoEdiAPVX9BgoixbUR+mH3vCnOp
C0QlsWa2tXxjH/BU+rJ/gt0+ngaCpnhaQO0sM1drMNmWODQ+JEB1w+vZBVwH9UwZ
EST4dfKutZhN0jbs2p4kFYSKPHNknO0D4fyfTBx+UapRczjDn26/L5boO7iIU56J
AAE5O1IiCLOYuXHjTFUqOVwh6VuGFVgZjcdoutQ6r7FpSqv+9QvBq4b/NHXCETTe
kOIVnxYZTRRpzbAzoA0qLr3rfHbKuioFaGbadXqoR/F4JHHFCf+QABRky4BrTmNd
VNmXBv237XzMt87rZK+FBjCKMDdlZZrYWZaK8rMPUHzTpf2Bu+drHQFEjyYn49Yn
nscxZKcv+InGaWvRQXiazNLeBIrM3x7IkWrB7lXrv4NOrcR39gXoRMA39eFdktsI
G7N8b+MXgl6AEXzQsf532MKJwQSNrapuZO6oY0jJWRYq/cdQwwTEJCzgf7EbSXaD
PLSF94ia0cBljzz26+FQcl+hv2U4eWxj4j9EUeAX53UhSydeprvJGNWplMYzdgvG
vHWxGVWLxtJYOPK07wjs7GDymazzj09/Htbt/y9N9fWTYsK49pCJkUJrFp/4hLTX
97Rl+qAe5dx2rtHugyLz4JRq5BsnZ07jT34EdPVN+HIH1TmigRg0MTOn+fDQUpUo
xZkr9K0etzo2eLdtklIxm2FnuIlQAbW1jzbsF8f5huZkcLz0/AsoobMucas3SOsC
EBzQuqnLt5JuO/qhsDQBVJFLXjaJ9a/IwPM8PlO1ng6hQ5FW3gTkWoK4hJvU2dR7
k2J76RST4zPd/mQBNErkM+sLdXw46RNIKol/CbACqgTJeb4pXABMxtyuRGYOy9T7
CKOXC+bgmB0kQuj7fYpVYcUg4uFqRs4g2+dMwfKzixPO84NpUw3M8PsSynYfoMDC
whC1xFkktHNbIPk20c+/itKsFvnOhhIwlsEdQxRtRDIrgFtNe3G7nMbslpyPyQcQ
I5KpMi1xVUI/BiXuLm4TRqq9V60g78NDsQv1eS4H+pXcp1NLNpBFITTphFH/XHH+
SCh8tYVkIGVsMFLYrR9a/RFYRqE2vb3og/DWlizVzGkU1YhS2dC+B8Ny2rBI2POC
8XVLpFB6HpM5Z/0ngVBl/Dmjh2ZGCeLDEo6RddRN/22w70FJ5B6GkII92CYocUd7
9Brey9bEzakJmCpOKNqOylR/eAanmGSOetPzYi7j4cf3RIyPSYdwOM78avhPr4I7
12qRuhBrtITlL2vv1DqPfEIOgUSJU+cfIpg/fJRDMCDFkwPzL59DC6yhWZYgf3S/
cJlrXeNEkb0X4vkJLv9OykzhBRA6lq3XE9n/QPD1LG2ubThhDEAXmS7sp2M49EmY
accJ8CF/3SIdWcTuRyCtZ8M+uwpwvYz2KQcGpR01mrDhn6JapatgjqGd/hJ00BAq
2pXbNpGoAmSrB98IL/93lmLtsGVL9vqmwizwHGtvYF4sC5/X5syfj75amoQFATcq
e0JuLL6bKf0EFHnBK9mUyMi9KiLQzLbpHwFg7GPBd5c07ZB1/tL/uJYHlQlIoi0/
5nGniNMGpFRqt73K7Dvg/L5mwNSxpzRofhs3pBk7GnlSo/gdfBXvo3zjCvxpBpy/
uuJ7PM/8uDITDDKt/iFzVwaVSil9ZdSFZtDY4d3LHGc6RuK8vBXTdCEDAf+V3dGt
9sc9A8FYRuRWOw8CCdIIxhwEZ0pxkxmOsY0UjlI8nwEXolGz6oCfuyjZtv5MfmLU
7kDpbGTJVpNxIO/bkYC0h2vsOcgU5lpTfeqxc3gYFeSzQs09FnRL3Y3r3+k7tZSu
zTM8J1fc6J7SnjGcKlsH6daH4Y6vaCYC5qCbGe8Ee+tklTrFcYgTIIi0HQ+QqcLx
Fwmyg07EJ+EYeBobD/xL3DQzUt1rtBkMzgNOr4kzKAGeNaEDu/iDRnhEMH83HbWg
jir1g68zXnUKKJgngfAEKStTX65WfTaFyO37NDatrEBUeXitQScYaRbICGVNpWim
qx4jLIGL78NFkSMiwf+x0paxkWbEdJXiPlVO76H3dtZAb1I/Lg5OLN1RNVWgS8mb
0rpkO6xqsCfCnzaawsulOIwTNqNTGxKktPtPWqgDc6DS/3SfmcgszjBr5x9P1LS2
1s57RkKqVNmOQm+9BN979S0gUDaKx8awWCzIlGD2k5JdQ5A10EwHeUQEEfN4tqGY
osEhIa8hEvqzBd3xp+YtvhAYFmwJkJFp45UUpR+So27ly8XzBgRzLDc1QzCdEYLN
m8a0bmFrhv94qhiMjW3O+3mCn6b9Mvmrtjpc2bobubHr/4fY/2mDtAGusYOqv52/
yZQNaozWzlHBzsoyAH8YzOwu8YgrIaupS1wfNJ+0kSIMQAgsCfc4hgots2AH0a90
twX3ULLxAf31iVTvpWZP45vRFE7CxPc0y1OuBdLauEo9WKssf1jtEdiH/kT7V4lK
bFWrLpc/uoXrK4/XjWw4YO9tRIMebDuWRgbwgMLZkg0QEfkuMa54hYXuTNB3Vwuc
zN5oSAZdHsyPQA3bwkQhGCEAFNSzZen18tEYQjPiG6VCTqBQjlU37kghfvzxzVYP
rS+0dcnjT3rBhrlKQrQmBMt+2ACghJjd3PJ3ddAH8mq2SGH17K3TI1G3mWgHUa5a
RgUwyYl2ECmG6H0mkEgb/T92zm2HcNy5BjcL67uNO2J63uYyBScwyC6hUvcyDc4q
2jDo7qxhCz60V4qgUaPKC4AnVJIqndXThrHPrkbNGGSZao++iiM4jCeStjdJKqqm
ZT4Dkwhqr1v3kAW64mai5gp4uyeIJvkvpHC0Ar4KViTwiDKOD/eII4lx7p/wDtGy
KiefaiTY5QZYoUrIHe1NecAfBmyAaKgf499wJRnfdE8gCnmElCssgr4Q9KsaP+Hb
6C9s+kX0wBVC0omtL6ZM2ULABqggVm1h2fbwTYumrMMHiCUGdyVyp6IkdocPWx9H
JeiKdG0iri5H0WKrG+LNrcCZ2D4xjfE1cAQLkb2odNwG/ypBtGzoktanUceuQMQi
v+iVhPu+v6unzhfhEEJjWwGDllU/9KaJ8JyD1O/21kJbEWKqaqcxNN4pk6oOXbO0
AhiLbV70doppcMzW1ZfK3YvsBIgr+AyT6g28bEkUzbXzWhSqc9t3T9fw8/WP4g/Q
EhZqT5ZQiyPk5v4S33UNwoYNim/+7z9EIfepoPjlNB7kL8mPQmqX5WfuwqEpgEBj
FZfKxMDbZ2CyS/YZ+3FADN/j0tre9AIt8EBIQrTVJJ4bvjwBWKLqnctH4VYgtL+T
+WqLnbQ4Zq8anv1CooxoJ3O3QmkQ9S+C5Ni1j5GtTwWG+joEjiRbbersvOkL7gyb
STy4OPIWNqbQ3F6wpH9SeTyExmh91Cyf9O8J38gk6EQ2NiS8HpHpbzwDQ0VvNYPy
e9YF34/SNNKPY3FShOCNdZXg2BxC8ROzMUNm/J74a5UuBJ03VyDSEGSqA8Z45cTv
z9mahee+9S3N7p7Dk7k22xjME0ocs693MjIJcpSauh+SEZ8pQwp2xvEbkDBOp3fr
tLyw6Q2YukTkLfVBrV1enZcsyql74fddhgoxORZ0WbfFSb8h0FivcvtJYAqaJFZ6
dOyR+OPg+Fn5VhTRLmNvYsauCTG+jljfvUfCooumwSOwobPwVrX+DrLGoIe1PS4e
tGL5g6JyuBeqY1q9NtTmUKgzH9OOZ1Zd6KfF1qYudiEmXeHVpGxUfVckvND2Uiix
YJS/CgOHV2GF9PdGgvXZyhZosc7hvel7uU3SugKGvFnJFEFbmjpgq2ErQQTZSdTa
WeG2skcNLp4VZ2SlClsZBo7FRGhTKBDxCl6R6cuMMYj9sE1LBP+0vpw2MY3xZ9Nu
jQjG9d/BPCIvgT27Nws4ccP73K/sUa3qfptRcE/EsN16CVmsu9huFlCwONsyqIQ4
4E/hRI3lLXFGVNul+SGpbWs0XQFATb0tgxG+QLFAtL4bnCQK9IzO+phfHUMhpbPD
tF67mQgsDh/YeMkR/R/08sVRFAhq5aWgyta5zDQCiMFHhldsnO4SzoL/DLt8Rdgg
YtTEOebxNya2zUJlOr5Ty0es4nIfP+v9fz2gNQnt5uesZJBtnp2nw0M0FbWPx7lo
RU08i1BmdYQdBWlEVreDfDy1T2ICY7uVXD5a4lsGV5tVL5kkgeu/oSLQpyCNWuXR
40vPJdrhH4+WcALwNuyk0SDZ3XG32qqSaSAqsDq2rlYgnQl/0Lei8pX6pySJ4NTe
t2KTX5+jRTsoSvzG+iNCzKKT3OQcCd4TlCtxeYZMCXwT0rVuCDeKwjqiVJVyQUau
YX17acj+KoSEYR+H/RG9vYVZfj9OmAMGqG7a+8HJKKI7CgoZe2C1QImARDexkJPa
jaeCIxxLqZQ3Ho2ui8chFZcXy7Zlayw6x0sir+YiIwiGRnqFJRiTrfo5Lt8uDTBU
blkXEZ1IrY0QD/lSeyZh6ZN60c//54updtCWNn5xQy8Pl9uNNwy39TYnndrNpwTX
VOx4K0/oL/GkC+5hqXc1+/W9zmI+jJtZygJ7a/avQ6q6An7g03cuKUc4sQXV5aiE
YeK4zSvfWSAoCU0JbEmXhipqWfTRR+5Xlfjqqp9tilTkPaIvYE7l9c2mFk1a6WJ0
Qsimc34Ojd69uK3qOnrb4GoF2CPtGq1aubR1igZlOFoJ8jG3aOrhxK7Ezr6kBNg4
We94TEgEMEQq86JhZ+pZpaEst8hAIuBH4UwYqEF+P3Fx2+x6Spw8sBDQcrrGFlJ2
2VlIs79BVGWMnGr+Kl4gt+mW8Q4ql2uIUYwAEj5whViu3qASBNwmLTGeB2zqHcqw
IND2xeDS+K5xpok127029GlmpB+Ne/Ux6LoxMK7rZsZaz66N09iKlci7ImuWS3FK
YZeAuyB1cBGqV/U5MMWVbZPeCZZ+htWlzgEBvhg6LtQ+zkvXMlx4280NeCa1N/Q7
/7I5v2rZgy48X83OGrvfql03n8mv66KxZseU1Gxni4YqxbLV0LArgAiAaGsRXbSQ
rkBNYWDEazl3oU2GYiKGlHB36ftz856j10qfFxUu/TyMi67Blk+KoWLnls6y98i0
ubxTrv3Aw8Nv+fqJGi5RO0uYTj9NgOSIdDkfs/utVYBn2QO1ISR8KbKst1IVWbyO
QWDXuuwh9/h+d9zpdRWLYap2K0Yirh4IOspCwAqN7HU7GhQackra+IcPAROphLp0
20cRBdaHJVbNNcb2E8jFyAXB0Blqkrr7HxTZgsf0THMQ6JENGzWk8bLXsPHXgwzv
VtOoLn4zk23t/BJxijhPKVNALw4wuBxAsxeWzLNGCc1+npvsVrdSDICO4etCxvUX
lWTCzoIDYuQGhNhDRbj5pJv6h5/J6KQINj1z0VQ1uErAKJjZ4sydni6IFYnAwBiZ
tA1hyhwYiLP8xbvtd5jLgozbMI5lDiU8sTEa+rl64zJe7IjbcQycTbqHWdLIVoZS
otRvUWH1ACQKdoAVV99G+LBMT5Bl0Zt9ygAzmUv9hV6Vr28WtdFHsycwm5Ww67yJ
DsoN8usFzzpkqMdkiExk0Pn2E3Fxg6rcFchLsIvjpKpWkoSFM5Y77mt64olQtSXu
4RdfI4EqgUkPW33s3IEqX0CT4Jw9dt7pBoEIzTnBQm8SF121zDizASnIXNM3jmBG
VxS8nwM0IyBtUzsVXm6mMDnI0Q1EYT81qRXOJtuPndNoNQRsFdMZ4ICL7VgOWlWK
R8ElaHiQjzCqMN0PgF7KGkjU6pwFU/Zn0hkJtrBM9d/cmMFavBBH0hIOn+isQ0qP
Y1yHVz8uk7kyylkSmyWnsvnJURMCqJygVd3ibDzI3+Awm/sWogKVzms07VdIpyvp
PHx7tyhcc77RqOB7yEquWhiOk2fynJX3J9FJxtoDRHE6T3IEbyQ6eIz7nQU/aNnj
SfZPez2hLl90jCsNARZHTbOcPB+X31DtKeCmm69wQvjZb35h1TmQ4Kvk/DGZYRpy
0zPDXb62S4Cts6vL1XxeV58R+GdU07jGu/aFmjHvlM2LioqIiMjs4x/JpkJ+oREf
4iSyLBpLiC+watjnkNRwQT0+IANXPV7YHOK7G041DZyCKB+Q+etTeF28iSutF+60
jaUqsmgxyYUJef+UnF2oYPOSzO+gIg3SSTzXcfzWDmY0RvwpGF7ObeLvSzd9HHIM
EbxvhE9MwEyna8/RZYd/d8nbmVSedoU3BSvFU9NwyIRvc9BsL01YwCV32EW4MTcL
MdQsIJeTtnLQdYeb7O6Jbb9wW7u0Kseb+3UpCtdc+67GrSlCVGySNiQD+9QUPPtb
7Egarw3VMF5oy5BEVCHBWilrII4JWTuaw8PMdylbuoEQUCWPEwEgHACcuw8AOcT6
94BVRZpORvXxBX6aNvFjNSdYvYZuqx35n3s2V8ws5X9/UfKH+vTOszP35vhW5MFe
dFirHumPhNwQ3hDrRXLKypwIZMqlvkONdcilia9qnKplCxdjuCCL5eGiE9eahseQ
Kaj6UTiFc4RyhaMDu0/NRp1mChsBms7k9jW5pZS8SJn9P7yIp64t99TJrNoSwFbg
BrvTyHi/X5qbyYXu2sTfov7nSZig26sN9cuL0d2LwR8txU3EtOvtFqpEy/oVy++f
RvUXH0LlRuCei0mH+6obAppt/qP7VdH5Bf3TdTmjEYpeHIy+xTEdD5xOdhdkH+9n
PJVbteBNIyyujrKgW/8SN7FWrl1UurMNgS7RQt0t7zFJeU4xiR1D43HdmTi0SDaw
yo5S/lDZw3y5Sy6+QFoEeN8+zRPy2O7ID/WfTxb3IphQViPSd0pI59tKs+5FjhBB
C7hsDRwVE6cVCZZcOCAZ/ZGzvegEm8ITQwkMaTV72Mmzft/2Kuwez6/3tH/Ho4cC
C5Pj6LJuB6eHHnSsCHZIvt/uQAe6+dyku6SX+CO1Yia4ILWWESHo2thZC2kPq6Tt
CUCwPeHXrho3fH5+1a3iogf5ATuUBgDZ/DHwGdsFES2w9xeH2r5I+hkHQ8JsYCph
LS88yBEqErhN3mdlYLVI73GcwsXK7ZjkuTFnt1ay29x/ZORE8QAtx8uTghO09+iV
YK/Hbn13Zis6INkiCGrNv5jkRQuPz8ZIt9e7V93ybp6iRtqJ+5mlSBSZZ0vEsZBL
AXJBRkpLmKXSo2lxyBDijAVPwHS6Waf/aUhsIkP2q1ogMMpyVO/OzN+xSYHQNnk4
BI0vZnBXvO9+XWjkx3R4SQTg9z1m1EnbZEq2db0RgkuDfdShunuzvmvq657iTC9f
rIcoKXPOZO6QF0Q1H2VXZayUOry9yBVM6rEL6Y+DqiSX/Ed3GJKoxhLs5/19Z2gg
PXLKStj+jb2zmNfLC7wQ3d4TCbh15oL20UvVzkeecIIk16jwc1+unyWBFX3szswm
0nceyGHs5iHlk9RROIsEkMR0Fvo7Nn/l7dfmmuLBM8gDiJ79pjPVGgrQM86+niyd
/6q92eJ7dtI9HC+IjF891Q0okBcTgCBPVGdPuqQnjNX0C6rkKQ9AfFEvMrwsFVfa
GfRK/fXbzFfpcL87C5rFuDoq6aXF+ckbu93vw03BCD6TqQa5/O2cFPa7uaKidroW
ruWATarkFEaTgOqh/fsJDnRV5NPgIAQ/3/HaJjhQO/qpFyZrutdVUUMnU4Z/zqWI
Rwu9YIJvOcRb9aDVpE0XrirMS9uw1qbTOOisVWR9OwYBwzmsZPlQuXc5glQ68e7c
Ex8jbvCW8ZIgGKbLMtKSNpB4HineQjF242GrBYIfP25wVzWTA0dhQH1LCO60dHIu
Z8V4IEPFZ0UbrfJ9HT5sxzw1VHfe8vwF0vDpwzF7H6c+Fnrrc+MyBebMz8U0Ag52
00CSTDaGrHtVFDEoxB5LoKw6FwViG4X3lEI0RJVLVX1w0k7dAFpH+tsffJduw2c5
qlOP2t54JkzZ1XRKZC+0a4cMruVG/KKcZwGY7/jcCwK7ZwQrtvscE83SO1qwOu+n
oOKAU0kzqGJltsXqexJATtgTnEZr/6yyhXY1EBf6zoVG2ildlazpCONsIrhuwpBc
uBDv4/oQ2Y4XnFiMZkb3BYMkkFrvYpgpuUkGWcMGqgTKxmjwcmvpdv2XqVN3OHjJ
0tHyynOHtQ2N+Wz/R58QnJ/xw3ad+JxFENoodxptnveNasmx1Gl+I3OWuzcdPHdZ
PxsWa5O3DHqHnMZxP7Qsrgj5Fg12O3Cz5Vrh1D4tNQWAOf10pVqt5rKr2If4VOGS
E09+6/7pcmSlIaxoYaJdO1gW9oOmekIvkwgnu7vY0yCoZ/6WbXVaQr+Cx6TVFQdq
vGOQaogEFZuGxmxCCUoZ1hU8a4MrqS6kZErEDnnxZRYw1DV/LlfuzPdfOEX+xyM+
15tBYNHACXsJwgV6BjE7pe+v2nWMqFQWJATxNhDW8Z9wf797J9PiDQESNUVba0xo
bxcPsLEWm2KZ1x2W+8YkkMM8ii+GhS7C264tnqu76cFBsj6kohbUpq7uvQXZZUKA
+njjdjlKQRst8zIGfZn70sgeq7xcPpC/2mH86Im4mSQSwtdGPIAnqZNtPvRfdRqi
s27u5wKMEqV6a81PvtjXv978WoYKmkPON0ouYFu3Y5LVj6xjAiHg0JZgndg3PNRP
Vo7NqacfK/eJadV3Fh94ouZyN0+kNsx47lh14WnQmoYY0WC+A62g6O85RW16KVAu
uIR5kPGSBtuqCfC1sYDckpALO9dc15BN8CDlq0hzBtVqgRLkIZ74KXD9Z/JOHDL+
LQ1PI7Hhv9w2r9GTzaS/bfVIOr+5IGWvY89aeW2xDmRaezOHCfIjklfBx3sRBvqT
2JMQOzilp3ZGG0bHsGh86CM+AL/wH6K6TU3ZoUyBcPBmsQjxo3zkG+bMhcRYFPsJ
tEYFpksZPASfgnq0k6E3RyP9ZH8zeGe4iI8bzq5Fk8MuCdEg4HTr0iMlrm2SEaDL
T2We95tCfSHs0AFc3F1TYMlioy5Hji5zf4fYlbMs7kAoFAkYrQWDfYEHknH8eIpU
TYFVCRN0YH0/zdDdTxlTAf3czhRFJ9j0j9P9rAyU4ZnEBe2NhguRT1dnPiWpsFZ2
d5CYfZ/om2kToRp5bbK18O3m8IR6VLEsQkDTJcHhxE1qhW2zCKWLr0kK5ni6PsBm
fSC/PCPcjEQBnpEs5DQVumIc6wlKsUiQWJWm4wnmhdwHudkKMF7wvSVgLiDsOzJo
zsByLnyKRG79lkC7Xhplan0G6d3UzjRuyMAUXI5+Xe3JK16YyR/1RlUO9NaoDpfQ
bJ1El5y5kWh9hcGKe82qTMgbdHnCNz+AhOo3LPJVQ/U+y6+c8F4MvgCFd0pbzgj0
c/5BphCmIFPkgPCkVyA0A6h5k2jPP951+VtXDkmi7lkmy9yPE2eySEao0K8n4i/P
7D5SbA+3w8fkWmui2U+y7s5U/YGhpMcoeKVcOe0dJZGm+30floCOj2YPImU1ssKo
42+azx5OxI5hfNDvFAw+shVLRj7jRbO5FR4Kw085GE0EBxJAz8WJucCEd4p4lOPJ
HM/mVHSi3ImzOupKB1C3McWDpVz8pW94pQLpLPpsERzEooQGbkXvd/51CploDtkE
OS+sKI5aTTS6+uAPSRZsOfZVknbUM2kWkZ7ixNbsCbx+efvsI0D2+1d6LFf6/fg1
Cduo5vTp8d/KayyMv48fsB21GccXtHYErK6YbqwG+DxZMRhgJubjnfDYw+VUrlwn
AGruYW56Ox7CD18oJOzrPsVJHHLXbCPZ9bH9G74wn40nYlErOItsmav3gyhIR9ek
UmQVRXrSppsJuUOr15vS2uJYoNDDlHU+Y+NDJhxxv3xDxVDcdzu6CucyusmVRGG1
US9ukENCVs8EFuRpFVry31iD3SQx5pHCLNQO62brAPDmrV1x7BRbb1wa7Z8tBDus
h6VAX0Ymu8dGYc1agtd3ihtIvNe7AcbRhEnzilfQrqxStiZp+dBvtp6RP/+guKp+
4BifW5+Q6E896rosTMSlzn9KNGFDqYuWRGaJE0x+Hh6h0T9cRcjF31oM1fUIVT16
IXS1rucoY9AFc8SxIZOEjQtHshLoZxSTBuinpUFsgF5zg7J+Fd+yQMyKvU5m7jCy
g/1wOydeyo3UDyZrfFKCqGH3j+9LwdtyXG+pmEWAa4U7IN4vWWIjv68XXx9f12Ku
4qIEo5v8XBoViyFAULbM8NxBAofZLzGghRGOizdvU+cwiThNhhTVE09xpxeOHcvn
139PEnQCX9AI63zxCMSVQxu4GHvFzjaQGA1gZ7thSlMC1JJ8R3tW5eijPeBL41J4
AZnp6qek3BltCcwda49jL+twuZVsiRSZ1AHsQj8cn+JKZJB9HQl2qoz/gqrg6/EP
9sxt/yrIvtvM0YrV6niDsUglAw4vj1pkhUU0MA3mo/LCFVZTDhrYj7H5nvr9eQV9
t9Mz3TYv5zaTuv2BM1A2H41AL6DSyxc6/vYTrFcn+I8CjR69BcwqLhj8FYhH2U9V
XJ1vHRSosrC4vHTCvJWTEfCvKEKhph7nJAkCnccPbY+llIbR0oS55KYGB8MPdlku
IsWRcvlKC1TqLp+EkF0d4pYK+yjo4JOajA4UMB467zHiUss8/zC32LL4HYuonn3m
5BHAnCSwSDZZhmOJ2onMQ91sYhVClWR/S76G3OxRkdhDUxGSml6MP5kO13Enhgul
gAAmYmuplhKrUi8htHNSLEIAeb7harVneUIf9vgs3Mz+V/Jj9biRsuQ68lZAYmd+
t5DhJ3DysO6V6jU7Fu9mlAQ585Ib4wXvfcu3FroCWC/VwhXkcZoFoKn8xcz5yUO/
dhFhFx+iuxFRhy3TzLFXWD3IS1pKyldSvMiK9AAIT6ZGImoOQj9LDuRqvlfM8nEB
O+WPvHUnreOSrzwmt0wnGxAGrBMn7PMWSY98KGmegxsdzYexnB5U96WKYo9v+/EH
wgUbNBjSlS1Sb3tIWg9/lc1hlS7Fh5aohIMdvrmPO2kKxM0uLNgxrqMKtoze59rZ
HwQCPYLfy5qU0gFpqrqaKpVyJMIGQiQG5oyQ0amXos26yrrgGu62xsgNtCUgddoo
iLKopG0812hXSNgmEiVeXFmCnMifbBmh4ljt8iU5tzIWLYdqHK0/TOhTGCHYchUS
Vfb+Ni5xI9XxBgAJwYsWRsfMmz3t03w4Ce3EIEUfSYRSb3XuqqML9zqcAHsItwfs
TttGUC3kKgug8ggwE9EXgTwkfGpWKp5hGAhTJe8jQkr+Y1JLPXj+r9RhJrLZclzI
zDneJ8TvfLDYy4dYljqt/EqUAKUEQwhOYUCL+7AcMhhYxzjNgBVUwWQcmz93r3Ne
j+19la2ZE40nK0PicnObvcNpmPnMbxanneDkttE+oLmT4lsuxJKZhA5z7qsFEmWZ
jSdHWHSjpn3ehZQK5zOVRQ39+W9ce32Du06c6SKRPLHf9YhTu1EA9AOHAw7vFo/h
ncH+N7b3kAyaIGyEHmkvR1mjgb+2hy2szwoLng7valkJw46x4zJGnpHH/T+KBmhb
CJDaoNXSt0itduuTTn6x8HA69zm/6zl2uK2Vbff70kvy9xSug5u0tXueqX12Qn/F
HOkzxtc3gDqcy9RXxkTkDmlA2JOTPyxSrjZtjkI6jHq0vzexFLmYHANtoySLBR0p
MWU/6P8/xvbSCuRc7SpxsdCXafnLy1uMyxYGTDJdqAWkmrvE/bD3TOqjM/e4W9Bk
Njy1w/kAS7YaVnGuaTQk/9sJnHsZ9G/jEniHS9n2OCHlMJAU2ucnuCzh50TPQjke
dNfTwXHcUpm/yO5UEh+0k3cWn2R2AwTQNOegAZdBhq0GtrwTHnV5Hc5XWs5yl1gY
nD5U2TGIiSOMadX1k5PWfbpo0yE/Axne/U+QVF4wfkbUBI4GuRBd8UM+4rB3cOoM
uvs5gsGJcmiGnq+8weP1cx8f+5J7TOn7qZHctHHYvhMslNebiiW/VZlDTgwSWRYk
iY3IDNhWfuaG2v/voClEixHiwjB6d1JXZPirmzx7G10Bl/ovxnRF0NkPE9wBkVKE
4Ta1Y4jRqXfO9KyHTg7zjm1nYJLvzCGdAcHEt3BfEHsuYw+pKtQ28KB9XeXyoPAw
L2xqRvNV9AU4d4QhPonz1yHoR1kFNkWuIQCcdxboGtVFaXzfeWRJD5vIldSDNq2v
HPBE0h1f7Jt6vEPj/L5y3+qFo1ji7epUCqJscrsO0siXP/2aX4BzGTc/U0dZJZ2A
8UCxAoqEfkmLYlLeI6OHyMu6kRCzqjFuwZStLyHVG7nhhknNE4z05fBH0xqBAotw
oW9JGEVdciH5DB+LI28IF5s2m5/M1CRMRV7ZgOAy6Qqixj1ATPbeuVfOQIW4HWnI
yaVUAscvvQzXEF0yBIWgn5G3cIj9xRsRXMZYtrJIfjmSaXQuvnYNZi9xAaWEJccs
AnQxjBTRGYp1bhcP5LnAxk6NNSw/IX8Rq9sq+K0q1QvvrOjpbFzNOjO3FFvgTuNn
pfrtKJs/zxwXGxKzDkg3qSEJk9XGP2p43fwSlHNG3P9RY9ejtix0KTPBEQk05o0q
mg+yaCXxliILAcm4TLIRAXKNFq0gIqKKthcg7BOAlmGcvQBP9K4cFTajL6Wp6fRO
pH0bQGp9SQMsElAWFDUKz1RkzxKivw8vsy62ZK2XzBprawLIH+Tx4zYeYd2Tt4Ve
yuSJbeHjMXUfhw70jrrBznjEXvrEoG5q0eJV+vnSHYXVDnDoYyWlVtDXmSUTdXlV
v18iEjO7Ix3AZAVnejalPlvcfJf6u7rFZkbANNgDkuQL7D3lj8ltc4g1qh0t+HOA
4zmibilMbsN79wdaFFEQA5c/qTnolY28aJwjLeGIZwhH31BPmSdMxbjWuluy4+2G
Fn/bokRSXhRdlZ7ZlHXVArydcLZc7BgZgYjRUuwhIPqoaOXM3OrUySDluQuuUNd2
pCqS2il9XB11ZI9iqrqsdLSil8Q/CTMdpULgIZ5JlqZOaiJwCN5bmNDFzQCefeSu
tjLon2/LC/kLkzGBRwhnWxQfHnT6G1jYGq8l3jw/CykQNnlVjKMuHIbBV3i1XYTi
uurVhh3v0JijaMuGIErecWw8nM8BIJ2+ACpyMrvUNetBojf4If5pVx432yT64NPL
+1mHI0WLiUcQRHkbDiFVmz3KfjDLsS8Og+tjG90VMaDqNlfCOJwNwI12uWeI+Brs
5cabrIzL0tZdUmfcQcmIScI8l4unI954umh3+CdtaVhXWaZYBDN+bQxJ1DPnwJl+
yG/AU8DXJmsBRWmKxEEa5S4RElYbEMDh3h5nk3hcCDggai5QD+lMZ6G7tHY9VX5m
N3skaNdSWePak/IoJSUq+xAob9GOmwX2SrfRphxfGM7fi5c7rZ396zE5/fj/JFh5
+qyg0EWDgdHdy1aPlvkP1KBaW71AO2qqqHOt5HAGstppth1FbAGgdOfXfSVzcDgu
It8xqkNmmEiQQVfM2NZ9LHIqaJ69xTbjp26E1DkYaQbh8dekCULEC6zMbHmA+8vx
xqnouwrkSJ1pCGy3TClgRvAGCAhJ9RWVYSc7dmnAiWtcR3Ho2rOm8doR45pNEtJ2
aAUvGy5xRpd5X49+/smLLFGIK89SOUVJ98yXDaQMfx8YKmjTSmEU+wFxGpwfIuUl
gH2oaAPW+y6Rj6CqCILYCcJvrY4+K3mbkEIxs60/rCJDbNRG4A5aIx7t2QSztAyT
pxdlniMuol7ACmJR604BdpiGCrfYlm1bMC7lsoJUI47oyjqP0QzWg/VPp+m89nuI
qK2VUk5mmjJbrnJMp3eIF6kDJgfCN/N9eFTD7g4LCuY1wq55Zvc1yhRswyYSh8/N
gIwjIt1M5wvwvrN8mHs1A5Kos16h/DRYjLMPXqMcr6v1BU2ezc/2DQv0+AbHLrAF
hq7UotcGTE7Bs74geDNvzt/7a+cFdSMd4Z/l9jKRius+w+PYHL53VTQfts6Vp6Zd
Rd6DS0iHiMmXAptH0wArK6zANZAtauZAnSpDUeTqkUVSOeXNL9ner6THPoc/RHGy
6+dzGcAPoUQ7tzi3Kj9USzuf+wP/Vm2cRjddxLOVjZGdYkQPamDM3NDp+LA7L+3P
sFwBeRZurQsncnH2qY9XDItvMRzG4ZETxqFaKB1/spitI2O025NcHynakpqL8n3b
q3XPEKR8j5XuqT4kLyuIk32UCdYESLUw4hy9jJ4K0hA17NhFF55im3Sf1bLpfNtn
nJxZy/juXEk7EZddzs0/3WcuwsjbfwnGFo+WJpFQIIR/dK4jjTCtKz74LIGlkpVM
kW7uP2v5q1Dz0NiqxZJtR4DsS6PMdaFT9bR5sDtuA/enGANbfStahGSxmLSW/ZQt
jekqs+qnlkXJ+zwlonJAr/iz9OBbjUwjukfT2knxHNPLFv5/ziWmzcHmroq4rWMz
/eJUsev8k7YHieXAywYf34fmXoNkRkL4O3MDMTc+A4wmbP2DYJXRQUArHrg/6d9r
r+6WG2uR7NArFVPSTrWVIbMpTNu6qyl+zmbvo4AgGPwRMh60i7hSNtM2+tG4no9N
E1e3qSdi5x4XQ8hCnbKFvm2HPD8U0A54wOe4CKXlyNy9ygfPWM7uxbQszD4qy8py
sC87aHncwrbpXC2cbBievPMzTs6eiODhTlIOSx0rszhwMq+/ZU4cAlIv6e/P/1P7
L3vkRbSOAmubXUV/rTlFM99owdZQ+HhELLp2LDAXBoYxVjkJf0dQcWsZ6aVXrEbR
RnX2UpCazvsOeFZSjw51GgeVyzva9jO8h0C4/AiiTSonhbIiGekdB0eBSIyRQupr
zQU8t+SK/JMLyAYxevRJIzp/m4a0Idr62bmlmmuHTOSDUPRxry19TpQ8+/7nFfdb
Ftp3ms79wBTFzUMhwY8KdPaV8JmAh1BFWcvRhnFgBvcDBIOQf0vzPiBKfAcr+nMC
if1w39MbK0EfBZz+je3fjCiMKQvVzFIhk/Ap3Okc8N10+Jvbwr80/ynwro5gaT9a
2VU1oX+Go4PsDPCv+aoymP7nrt4QvlMKtb/D2ozfVDzcP2/PQGKaSjlWYkoNjWm/
1iXcjILajwub5SOpIcCGgeqR/gNReycaMl6fitaSIC2biveE0lbTUYMMNbUMzMnp
iApzDTE0e82iTackm0jMZQIbztqo1t0+JcoxrmHQ7mCIKXfLl++wtcu/Kn05naJe
MOPAfhOm/PlFX1oFOWlzJD8+U9371Kbyyam+tQ0rQEU2L8O1QovIohSxb+8pbZAv
pfktODf0BWurqqNnv0vbYZGxS4n/CWRjD4LRlmK1cZnIt7RW1sFK74DUpbWy1OAx
0Uc20bvGDtO/+c6DuMGz1pPBJi/gVdWabCFg1IYrUXBMZMw1Tz8K4PdbvMhjgawZ
sED7rlrJZxC0pJB8wvFlUoOD9oE4ZtFkgqRjR0CsrJ4AaMMi7vWLommn4pJ67ark
nE/+/rHbBnY76DmUSd7ZEB1gkHDyn0ku2WxMuZmUxwj6zNaZg8vBDphEWlH7MzX1
Lw4r0AM3VwisjQIxqvauC7oX5bG2KgOG//Jd709W3hNQUm4f2ClyI38sbdsEIX7S
drAtzTCWdHite0dgyHYneq7EZsRF/TnYfC6913SnzDiOyGotN5GIff4at8eviwyr
Tvpc8J5Yhh8dSKDv6pJ3hKRIDF3FWkeF6CKri/ZT1Uo80Qn4RsPLj6r6NY5GfjgE
kd13SmM3yy5TO50UWkg7F8IfhdtplQsW8hJIImz6sSojnMFoPFG2wyi3O6/q+zGJ
lPKV9YaPP/xku1CrEJNWs8PVA0xpPK4OYQ2gEv7GBkUQ9Y/vuiMn2zIVHxqpilRN
CTw/ybhrqmn7TDvtLjoa4rGIYBz1zacqaSXHScOZHVgKXNjlK1YiYxtqErUSza3m
Bi7oJ7mtfDLWKk+TO0Z5KT6t2Ctl3x38thQ/gGfR/y19COdsq/4T9sgeXeOwxZJJ
KRScFibJnPycI49GIvoDVBZIx8y8zn89JkejmpUNukKKji+QI6MDLQ5lsssshEi6
1RD7C1h/heU/gPedOUheXIUAoX6lgYSx9vlE6s8Q4E3NcQ14tC/lCnY/TkW41yjF
wV4YcoZ1W3i9ptBwBECBsFjTcUTGtILj0TXx8vvT7RCX9SOGmKFVuzpepeCC3Qs0
dQCWqWxidIYnmvpcjlGK9vezxH/u339ygeBpmiaekmkVNt2Mvok8Nne2ID56MhG6
nJGIWZ60F//gzi7ZmXHG2CZmNy2O8QxABpxDsZq7na81xWJ3DCjWefavE9CAPeZQ
tIVHrH2AsC0erjveDHEQhAawsBD1r6t67NqB3FU0xMIAvdDmFm7C5AejNZbklAGX
l/91V4ZCaGIfNgBzfm8EW9I29ElrRVN03EC3N02tLFGkyJT2R7ttEoesRervRAG1
2gQ+xkYkK+rYL1FNDv8AP+dOTgiBBZfbUKRUB88pW2GiZzal9QC7awyKSWe5gWTu
4xM1aafc4fPUsl8ijl1BVa8RoFvyigey0WyGfdvkwsRfXU1vE4AvG9Rdl3Fgn2BB
g37GK8c0ONvNDTVPCBBxBerrmKI99mTjLgd4ZqFozWPhFLJi0WYylXQ+5XVbbC3O
Mr0lNIXYS9pp4YP9wyMBJ5outdXiwyxkNlARL0tUHsiwa6+7kyK2y7+zSPrHqtKI
ZgoVFr1yotw+cgJfdkHTVDrpbw0zpP9dkGLQGX4yW/dXLPKhqbOpNfiF0krK0sxZ
j7eMtYwxdkud/Ifqcs8eoKpPKGg/qmYn9fPVafj8xCw8zkO/xQC7gZ4dIIJp+gab
prsPId2VHyPfmxjUKXTkE1KnR9IOOBllRi94nw7u7oBFUsT3HxgqwWj84x999lM0
MGhKpOp8UrM44O5Q1ToG0AFmjQix8wMXe9ZRv4oAcrGfXSWU806il3fQhr9XgrYY
a7jSSwGtGpvxD2x5CLlgve0yP52N+F0YGL09cTm6hKyjqNc0gdpdXGlRfqPvfEOh
2mTtJixgLTuj1QoCOmlzpfp8VQbjZ6/JQbCUknnklLD0g547NDz9zzZcC5OBn2C5
USbYLDDnlEMyzDEI74EQtdn66uFUqhvkXXI4L5eVqLVc8/+kl9OGvdOrJ4HqZPii
p8aMMmmEajTs+fT4576BgVD4FmL4ze7AI83gSA0hfwfEDuk2r8EN2ymrd4oq+VXt
ipGY9iUcTYcbVXtUaYJVD2jN1Ya7SlRFGnukYeLJHhxiLNdu79LK6gGEalXou6Dp
n6Gy5k48274RF56d9XsMp+CBUqRxdckuvjwpfAuwhxJGFncCRXdzsyUEo4/1waGx
ft5LxoJUVzEzs9VpFpShEQalpJAeDX71prVGO5g9Uq+1se88BP3uVpTcYnOUBGi5
bgaKYbOegF1uHUPpFnyoC+hVgVAc6XOQG5bbQSbKs1xqMrwuSWCLdIsidnvXgM9J
hmmOJciJ+ClTHJp1MqwnbLUICAkFqrcp55hvOR8/A4K76JvVGJ457ipZ+2LYYB5S
Bl/8AjvHUavxJBF97z5+DHkjVZmyKa39+tOo3i9vzhVJgYa21rbqqwCtn4/wLwbB
857knalN936knrLeR6UdsE8W1BGWJmClKPQioBLPUhG444Ca+oRAF/DTfyJIGJkv
o+uhsd2WKBQ3XrnC5xeUlltDtJbscMWX8DJ6ocJuaB8L+j3zC6lPQvhZWqhAxaxF
2ypumx+rF7qYjVZQJL/yBg8YjYnUE/TkRY57WIwBNejC8zEEREs6h8oXqabUFVl4
rLRJ4h6TjTH1lfqBJicPjtPXKVX2Da52axMrm6duIaGzQZGqniaIzWJ+4dPuBpby
zq9xPuSMMAkFxN8wdNNF4CyCy+UHit8T8Z6nVHgzuwD6QbcHynBtxclSzZH6UuxH
/7tu9mD+jf68nIKgQKL7ecFMPGVfB3jUJKh4QuHCKqdYCQ7PkYwRAqhKSqK2R0Kd
+ipX2BINJ3TAhPmOJu1AcNOG3/bayfeJ7CmpwBpkWXAUw7c9hNC4ftH8SlvSUoCk
BjSxZSlDf6/mbBDYIBHp3cwmAJ5au/ACFqI+SSTWBWlFpWPnVUky0xXFhQCkM4Td
xmhHNcqaT03UuCgx9s/uKNsE2F5CkmX1BA65Ao+2jdgYsiiu9Y5fXVyJ0wBNyecN
P0fQJdPbIe5mf5IZmtuexwpX+/yHFyrXWFNMVtgd2xcl2rDm+66gKgTMOo8vOGr8
nX/YqJcJNWgRX9GtpucgycOAwY+VZXYQkVkUW0Bqb5DW47iL4rHC38vPteMWuW80
urne4jbOOAiIcnuF5+yVGDX2bHbS3RnCGxXqVOJHe/w7HVw80OoVTHr+kCjDjBgB
uWTLSXz1R11qeZmBamTSMhg2fqA7nUP8Z3F3wpMirmay6fdjtH3qN4kYheL2kEDU
F9bE1m9S0A25FFXqX/xKfP0JlvsH3vYLU8aUZFygUhroY68h/BgapJuROnRr8f9e
mzfXghTi3w42/mn7qRYxDtflov8UMb1JIpgb3oRi98j2W5IeJcIu/Ka4TJn/W0l4
2jU0HS3nneIwn2YXfU7Db1jP/cSW8qxFwbMW5XMrRnA2FUf4udqeI46KvzyicsMu
s5S8uTHa44m7XRJY3eRDBvNL5BuKKkHrQ8n6z9OQrAiIillAYtUfOM7s7qb/RYJX
wm5IkSsi8JWLwXfjTQ3psaQXtppwET/mCKIK5HFuPOXMjtcxajX6TMyJp7EDtdP7
ORhJNE3oIDU6PJGMqw7H3NW2WZG9Z44mmozXLpC2OEwoaotGkJ7OXWE+jgWuubxg
i3fPJj3vFFjSnQJAtdv0n1B1CVgq/A89tjNjfYHhxg27jF/qUJTNaJSRsuIvgaY0
gpqaRVxTX+cesJyrE7Pzxxx+YL8fUUYL9OCLsOPOUhvVpR3ZQRQz2n7j7VRyGzNJ
G0ko+hOGuoRs8Sa48SnL1MqOJ6oioL3gJBCvOtrsGPaJ5cOQ0g2fSZ/MjLdatFUB
/a35ZCSXlFJFlEI4qgJLqt91K8t5BXyOGX/xBLqVnAojcTOOr/oVLvvVPX53kayN
GdWbiLT5ncuY9Xcs3AO7JpeAR8PIZA+Sl7tTbTNaOx/KsqV4AXrbY9Y/veJlTdY1
rxDX+vkMfxiYyVbzgJ107yLK9rMgOpIjGhTZ8I6By6GG5kEdYUW6XDrPC4cRCKzt
B3Q1C/VIV90wLw6Wl3JNWm4c0gi1YMw7IEkD9wXQVxATbAixKJRN15PUeNtfG2oh
g0EZYv0MnRaz4Wmmf+awAhgP9IgXlQkkxKg4pY9/nNyQ7BoU7QQycZm8+dJwKRLU
BxLtKeLQcjrT3Dug3hnscRCNrnmIj451+Qlm1kR8VtN+P/qPF+xueyS0Fql/DoO9
ZJ59QwdhuRnB4pXiqsuWDU9yAoyiZBI5xzu0yk2WfqtoS6xr3QdED6FLMghzH3qr
Iq0yP9uVXW+nUWqFl8Vk9fVDOe2/Ra3l2rWrHbXYBUuZSkXPaDufWP3E4zd4eBCZ
m4xo26+7ifr2KiAGgsGpZmRaZ9iWb7mBryawRAkO1MM7mbMzMjog0dS8LR7XlOhn
EGX4oI06dvVwVMOtzkGmRQg3JyGpZKIRxHHrfabwzynkbRTh2DWRv6Weo/3EF+Ro
c4VDjhH/o35oy8kynFP5Te8FmZhBbtGy9cD3qjQpWVCE0R/r/yxIeeQUEH2rL2Hi
4uVy2WlcCdLT02JKCm/yhsw4pf3rcq8KAAexv16sXolALScx+YkerXhSUZQZB6/S
xkUcpbZYJ35DIs91bzV/b1Zp3OUEUgNDJDE3lkxjFEAZN/9gBBM12Q6PTdLP/F5S
R+Lexp1ouxbmAh1403RBApTyqNVxqw/9KUOB6ZZhdMLlSmLHx9c3Th5+CJiqoMaq
PVM2vLT2DupckPJuBDlHvlg/BSTCvGAxuuRGAC5h3pE4jC4STPKyAQAxetIjUkvx
O3QNwtjqUL/aUyElSYcb3Jabt4mMu2SCENoqi+Zxw01wKGtl5rEvI+yKbZkiZq4M
aBIJFhtq7q/zpnJjSURO0hjPEKmRzCnUKZul6g8Y03RnPRkk5/dQTc/re24APcZl
cp6iJpqBaOar81tNagZlo3Z6mupeJQoG6fP8+3Oqefc+3XxGDeWLyZGw6g5gZCro
GYkvo76C+HGp9lQ3HoPtSoRPZmTRLbPSddoeBSMD/4Y47fQZb3IYvlcU9VGp2U//
mxo0BPj4jihUoQlMa04/0RhEK39K5TE0/rtEPS4V3/1Hd2zGgJ679VkgzfXtgki4
aovOlFSYVlpNlMfdVPvwNjU7p3iC2hTkFdhPFJip+9fp1tE1/56xYPp4vq36NcGR
MsC2IhEvCHGEK28HAkpgPBKodhw578bqkCTAZepqM0AD7rnCg99vJ/Z0M8nVmhRE
aMY9h2survLoBBoyTWWlSeSciJXmc7et7yv+ffHWKzX6B9ONGrozVNy1xYqZ+4pB
Za1YEIvHDAoxEQy/xkx95eGcuRDsDJ9xJDO7fBjEjgtdL4rlH3PTSfPXGq3v8hb9
6f6YRTzU6mZNgQ4oP+KuJjsMsdrxNTuKQXJaQAJ1w47LkfNxbkd0speWGL69Card
+GBziEAYlDu56HJ7QhmoFBWSldO4okmWfcDFSD9RaE9A0H2Tgwi4Q5czN134XGSI
OZTuRqIeVSIXAIaKr2KFstg1Ga4ZLuueju0EABP3/4N5RlSQQ949eRCqvcivWZH6
SSaOw+mbYfsiKsyHoNk9m0mmndkqL7gVy5+O9Sz9dX40HB5tKjm+MYM8aZCdoNUF
Yx0zrg3fDwg4pdsiF2/IpniwTRYYbZ3whQ/pkSz9pSKU4byRJNZwqE1+tpaAss2/
oTHMXgSfhyutZQIogMC1+UjFTegAOopXFsN4NYJejrwYTumPzYOIBrzzCsGG6KBU
84tRK0yPg4iFzObryvFzKu4dmmlbW3P5E7VeIyW35bJInWeSJkqHh/ONEyht1Yun
bxGu4IVl6/S/tx+TmXTa/ideDjC7Gz488qrHXFOp+l338pkhaL0ji3X7ZY+CgFyH
aHgVWQfJMizNF81obiqyJl3Ol+a7hzYMeBTdMlCKTlEiOgbLy5yI0Oi1q1/tR4eM
6UuaBucBej9dMH021eHD6mUZM915cZh7ZIXd95Gc1r+S+U+Rf4tEDcaEp5RvYyl9
oqURg0UPbes8tcklFoN4fMlXFbbfDLxU9rHi+MY0AX4+H0+HhT6TNzIITr8+e8jp
yZMuCodcud2gcg3syqW+/KYnY4N6zMujFmejqIBrepBN2PL8rbMQpuucN+u6yGta
9MwKx8QzH+CzlabRVq/p+1CyHEqUFcOGTzFfRKOf39J0C+BydkywpL9RM/uAG07z
9kMOI3OlumpWrLvtuZ5F1U+5Wbr4K34t+YAMFiwX7bP5inMjUA8u3fyHGHgymSLc
QSnULdXlp05CL94Sxkcb4xI6W4sgdgz8DHkbTeFElBi4QTbiD0mwXc6C4G3PBKaC
8k8iPHFXkh0mvMBGToaqybxFIvhLQdkbNVDdZGCxFZRd9nVWnD+/l+DSRNNkPSJj
Aq/p3E+Ui97jfXcQUbkqbNemJJlaiN1qQ8ISVEYnIpcGr4c+DRdVK5VpsSVT8DzM
/vP/p4je/66JTorcX1WKT+OQEzGmZuY8QgPyZ9YlIQX6evRSFmoXhzzaSG8c8dOe
czilwaMXkJkFQaMWKTe04rWKRwe9qXPKOzAW0b9GD+pzbpMJkFKKYQ+UbGfN2GUC
1ZTxkEGUqJFprCNFV4ZtKueyZtWvLshaZtZot/wtlC8Xz6Kyjl2VBaLl5dz8JjxY
NEo9BFtrb3HAsJ1m8wxWxvxHG6QIHI9eW9wy2wbzNwuTEVqDgviDCJV/POZViT/v
dztBxBpe5bPhlr7WrEm51F3Cpcbjuv679OS+A7o5XSeW8GDV/GDgjz6q8/77fvWP
y5sM6hncAtKeor8mSpIUgIedzAKFbH+R7BfKrWWwQ+hR/1pSUlbMub618xuQOYG4
vH7XLYTnCBdvQwnd+E3jltDMaOe6cFyCuwE0NTjOcscSFDjrmmNsa21ZKBemQrMr
mhZ/iLoK6omry89kyClNxa/4x3VzySbA7FOZ8IAzqORdHDbflN6Jyw6oKJ+XhDYU
+oz9UA18+IA7IXayfRSPzIlE53kuLlnDdqffzCxcJK9sVhkM1kLU7xh9/4Yau7Tl
003HP930Y2lgmaJFlxyDFUdxQgZzHLFtOemtBEtPgTWSG8zrDv/xXmdrn4GTtZDO
5ndV10RzmbyStXK1Q92MRlPQzNxyciCtPYYKKkh7RKuvX48BRezFKxSstHfHrn4P
WcmcH7dTX4D8sPqrYZAvu5TIkril5OED6XHeaAmhbVxgdHvNrL2pbYLUwgu1kQm+
qvlMWPwrQd3/tTjnLtpsK7Jx9F977LyuFziwIQ8/qiuMrf21eugjJxo5AIlXUMKj
BqLVE3wiY02w+7EACSxZ4BLSmjb91LTD6tCEPanj8/DmqMTn/1VygsYpXuFTXIn/
OyWn+U1T00iH9+YJpA9BIWctBrodyF9uT1fzGzhIJkZQm20AcoUo746eKawOctyp
5kEaD6P6mbGa/NPh95ZIOdrZa17yQH5ZnPQ1INSd8Zbwm9V/3zeNhHvVMpnJ9iUb
pth/NYeFHUgv5OWDsxrQ5QijyhsUDw+Dv57rCHNVRj6OahAN6qTgnMP7QkHQHRld
cRI3IHWcGSUUXnfjxBQ3UYnTeU2GmPDG3vgKqI5nFmxUaD0L7tLTy3Ex3lWGbxtv
ViozABwZu+kES3K3rRr4YquAXJrwlUAcUS8M1RrcFHMGJaytTOr+PNVqSUmEVA/3
BbJ7sl9lbgUk/jZplMvwLZyX1RMiLTVPCVlu+BT1I7rBGdgZB7SkYX/nw37okQgn
PqKXEk25t0rXQsSP4R507A24Xdzfgy7bMfwvgfQOVfhs6kcGshrR1GlNZijMPZtL
/jBsgtTPLwEd7erYE02EdLLzO4oCa5qEdaMIZUcKcvGfKqZRSGfor0MXuRc95hGQ
1ontuto11AzfNwkCBCQhsDnbCniWEIQaMdmyyXMvegzP8PQ/lDz4GuD87y3NNBU7
pYWE/CedoA5R9xLHPSueqDMaquWiOkLKfk1bubPjR/+ipwHg/WliBdtfwh5H3oGJ
b6oVhFSYBsY9khaEKAQKqVo09ftctLsNyT8NIIuOV54gi/34bgNXoWWwAIrnrZli
tfIQzYZamqK3leM2LDOI16GudCZwDYzddLVdVWC+abTULkpE0OOjbAB63lLzAb7z
qCMhvjskvPDruehHnRxAgjh26QsLWX/O/PDZqVbK89WGJcTFng9b52YHIU9noOrP
wELbKN2JA5AJgrKWyShZDNzqlEv+J/jO6fOCHJS3PcpqTwa5J9VV+eq86cHPFMSz
drhIwys0zJhAKazDU7ja501NobJDqAnNGqwVh6lYHyOEcaHmeORyt3u7QIENfL3D
apV4GW4R8n9Nv8Ge5sQbWFRWF8QSMiMtiXYJXHXW2IMQtHhlOZjCvi0JoHgV6hsr
xuBUiUgODd4x6viQn1wOP1mUVtjNLF8xR9wldIIOikcKi0NizqxPftUfnGAeh4B5
LMNupRW0r+Eg05SN49XArTSOdSGilLnlFffBMxb8ZtLhIJY/ZrMxt9cUxnkZ2LnZ
d4UJMNEXDrGwhH4qYqVa83czxfdACOazWpVwclPAkN+i8b7kYNnhVrfjjX9UotxX
pRPXx3XuajN6diXNf5Ds3qnDpOx9Xbfx6DuvGl3/Y7L1aZb6UpIGgGzgcxcoezW4
mSu6+aE7JyRiDJ2R2kR+VHqALVtLrfdPnECyylrm7UE0gaYEh673kpz5rUnblvrS
6ZZywX/3iMkD6WZktGlwgUFTE8pQTPfC29YzcPSgc6i8Yhph2oR9o/M5+fCAnter
pGeD12gZHvYQzm1uVWA4DdJoYGnJZGegWB01YBfwCw3KSDdQizRXmFYQr5ZKIVYB
MiZ8YxLo85GgN8Uywq1jpoQAvAn3YZbcrTECip4DlM68riV9kLF3mjxCBFtyxevB
ZUY3lyhp09ez/mgQDMGfUhMU6xe72/6YwSvLPH9HuLWewc/x4/SCqUukT0ZnIlGd
5DLLPloo3ub/RUT5kKxpHSZwJMcPZu9hza4RhRRMrfRY21VnL5c7fWqb2P8RbO5C
SR3P7clJNlYl0iw/I0eBU7KFhmRH+o8QD7qeFIxHtbQ39t76cMTsu4jcLKecDnxc
Au9Zc/5CX8eboR6fb9BTIhKqMzS6DG6MP6ocE20L1opxQVN9zNldH/52lAOz3Xlk
S0UO75gjDU9zkGUY9bvpZBSkCYPsS0Cb55EHXvFJoQEHTaArDNUAjN+iCbqIF6+i
vOG+QTGDbv5wJpGu5wk7VIfOd6qQujzbwKLQwzGi5eoPB6ivQpQmWhrHdyvaH6Vo
nNAEVGoV6EKZcVf5eeoWxVnjYsfuefDM6FZnn9W4Qn4kuDl4EUsLD0Nz+dcUiqmX
LlB8OWj952vIXvUqkaDxqibbXErCAHVDVUv+jyWqRUTX1qW+zGreWLTBUUx0LZAy
bx0VrOgifOTp1sWWPx2d79EoNu/841+CSGhuc6I5ulNhDT3NXCTs3SVQ36VtuXeS
uqdk7fAKzTKfWQHdz/Tm44T8W12ugpV8cghttcOInKbljpBCm1RffN5WXlvQGIio
KGgQybT+g+mTU3HP8EjZHGA0Jz+AakfcL4O+VW2ngFOT8Pu9qlZgeFkqnEuCXkFI
G0irTCk2B/KNudUS91LlJorpkonuOuE7+FVlb6eb3K5cOqCtY7WqZK/tszbcCaKl
ntndkkFK/A1lEckhvLNg3fXje4BdQqj4cffQ7f1+3fmu4mm7n6LvmWhVgR88tNNz
CMCWgimoC+3aXTcpEwRHh7nLEUVRJLplzAYdfgwwnxdg5HEHt0sPFSuXWpOZmDG+
BjEIDx2qzIKa1ryDnF232fXoYlfW4xilZJzJwDIcBerzyfc9dzJUtVzYslkX1+MD
KJtw9y6c2Bnw4GsRFwsPGTcd3GreYeJ+QwVo3RbwHkZV/jFUIfxVvgEmSS4fXUn8
vGSftJhbmyf6/rohHjg+VXrjc1rTffrLHKVoUQASxmjOIKRt4MsmkbBGftodg1FL
iZSPXOzJM8RveyHkCV/72mkI9e7W0/PUya2aTLpO9AG0vLPsvVkQu3xsvCjoQ5of
llFwDC4TOwwoE0/qF4znVrG9Jq+OhVwopfA/MYYIwbuBz4RGOFm6b+qSZrxRcCV6
Q7OKpDGCZG4jfn6RRtThwwUq43CQTe763TtS2tqxAlvJMvs93k3T6y3YWpAj/Lwy
jttSKScia9Rtu8rAULZuhUi0+HYIetDh02FHBKD+rhPuKevJC5ew6Vrl1rie4Us7
MBdeoMiLIMNLECZqoIS+nQB3tba8qnDC49g6W/97OpfpwxmINXkB5BCtw/LakY1m
D/bG8THB46kL54gxtNlhrrhC36yqIuqWrWLDXrQGAB8k+N6eXghp/PQl7QPlY8Qh
vYTkPY/fHtvL+/8gp/CIc+DLNqYhi3Ize18Z3ud6jM2oyWNCom1tECCs1b4XnXzT
+s5FQ+XUIBz73LSjlYDyWYNRYXg/L2Batzc637nurc/HiJsZqfQWw8kmTTcM2mjP
K9ynF7P1E1+Njn2yapOnTUXVIf89MPdIKoxX392PcE6Pzom829J7EBLthJHrkp7x
vWOjKcKWukDmAIP1KydABJF7mY1KDLQZ322VpPzpkfNalV7IuK0nfzgEu1DdA64p
BONzHHs9wj/Nl3sobV7jZztnvMc2LWykcYFu+9sULQh84jHL34e/vFc1YEzLMooY
mgeGp+FxejcYQJkndHWUxPINpuTph+mx3rI1UXE3rLkUY2TRysUWx2a1NPMdi6Ku
Hu1W8HVvwjBNaAuMeEzGKfEQcvInTtowoba506Gn+6xNNRNdA6zlpKh/lNQH91iB
GuzlusR3GuqsLgIehzLNUIfUc001jQguu+gzQkZTxe/rKraMhTG/HeLR+qHifbsj
VDAeHZmO+824NMI+2atSsNGXiHgpMX3mGXBx84NvA66mxW+7ocdxLqCb+4eN3K55
KcbAzNU7MEkR7jlCAwTqjiP2cdLCrN+mNL2tEiCS+E684XaSrMfHcLVmYgY/g7Hj
QDFLSXPx45Ka6Qv/NrKjBa0oTzrguLnLcZ/ghV3FRKkQoBLFDYkGFxHzTY/bzC3s
2sX82UVsTOFZAtA/5/JQJHKiquqNsfljLw4ahLWacEv8fw2o+uprhgxQKgAcQ5xe
Hnz1YZRd0unncfvApW6NAabDz47mMbxTn08LqLltx7S5NYZogLBoQ8DavVD5PPMp
3S/mnm4lsfih4C7rCcqNc0OLxjKEscsJJSa+BYoLGhjOVAdKtetwMoxSpN3jdaON
nRcvrnbwRTqyJr/+pXtQMExQrhgu68CLmD5UZ8HoUpU33JNw2dyxzYGhjjlX9wyt
hiMRPVumiVIyKPqLaWwtAuHBvDhD6dUXDcGt4u3bJElMAJ5XsJ/a3MrDpGCRBwq7
VUU3ONZI/tlR0Nyd7gxnorK/e8UrjDdKnQxR7fmLCmntUOeYYT4YNEte30MpwCpO
udpuD92G0/Z4lG0j/nnpz3qgUO2qCIwejOt+HaYWkB84i4WNl3lF+aSt6fpP9bzT
WMcBOydul0GqKScbbejkizV9b06FzvgXvfAE1pilbj353rS1IbccYkl1BW25lttE
g2BrZ20U0tk/8uOhrRj8d3f5my7gL+vq6hgUmnWJZtbB7gJvm2zldEW8JgDWdrrs
qzCyQ0goasuCPP/TVeJs2xQ3Ym3f20mbldM9HB4jP9z9lzoPjtyEqijx/lwU5wmZ
MUuVHmJvjAIxx4M0pcoonvXQhRajtk684qQS9f6hskqeZcgzbx+aKyAkMN03lBFm
lFQmmfj+ruwbHjHVb/e1ub5p5UBvyPmcV7DjrVt8jOh2EKK+iP/GUKXl+V1PT3aW
5mof71T1F/uMbAi57wxoRWYgoTY7ZnRIlKeEDkTezs9FygaXkgESl6B8AElzM7o3
+O4EU05tW8cO7b9IXkYcyG38kQLbe09D5IVSZbt/FTXfM+JwqhaAk91dW98blGb9
CnMbvJZoRK3pntddFehTYVw1xgAybnfKKO5PKDDvOgp7+/jB1EJCwbtr+VmnfKHL
EwwSDw1IoySypb2JSsLOjiiNol/q52qMzFY0YniTvcEo6ZHTPWkXetNhcxcBVuME
uYRMY9U346z0MOHe6aa70+RGyyhC0QB6fLBV/MPjVwCZ0xHsew8xKMrYkZQAY1j9
2NU/WXqFaUPxeLXD7qVrM+1sC0ov2i4xQ9ErEdE3nhD7LeTs9VboCTzMlkNuQL0k
l6kRj3ZbRD1WNHSuTb63Bt75wuZJW8enSVparsPKr6IoQlz9TE9wAYtd0vsuRJ/L
iUqBdUb7w9VW0CVAaVC4Bb3KiNQJh7VPpFTzNA1aEz9usCPLDyegn45Op1yU+h3q
KGFrfXH3OUhHG0A8H+bUeEV/fzvILcRmYnW5vm5GIcG0vhvgdmgOnChRPvhxt2k/
dyF1wITZf5W3/zypE7w2UUbLg52i6cpcLq0/T+rjjDUKhLrCX2W2mtto68CdgbHH
ke7eBBqe8xlHJyPCW5ochX5a7SC6YSr/PZbdZqhJh2zmz8hzuT+6xevZbb1WYCBi
0RjWijaVRNm1XhVeZ61kzvFBZ7jKAt1ZoHzMA0jdYjpb8Ahg2Z9FpNV1kDG4BOhx
BD98ZZ1pxRjIWJ62LjrT+Xq8y0CVOzGB8I9lOVTE9t0cvZWWs/FT1+h0KUzERuzp
fWLko82R7lV+yC5T+juJYyiAnQQNHcUOl4VpeejIpxdN6OFzGvIOSGu6KSoikrtS
ALDlRZnvy5DcQZA7XL7phVrfC6FNO/y63CSyatMrKwddiGZC+MggmHTOiYEwK/A2
EM12Di6opBFninQU50IuI4SI14b1Qly5OeMMn0c1VCIrytn3e1KQJsCXSa86z6HJ
TDXZpIhkSdkA3SdpLCT4UAVrgIN50hWT4/CD/ZRPlN7XwrQZ405q2isxtYcgHAXB
UIgr7FPEX1x0HbO3isBslvfni0xg6cU4aErME685XBoez0SeyT1j2pUscJlMIdVH
jtPamoTBgX+inwtKtMCINIwkfWxXlwSELnCndGMdhUJUHDlEzzoaa9OZW/dq673N
UrHA8ldiPO2J9xU3t98CwkGPexUOCz5Blu+ZVB+L7cBpd0LalIThkee/1qw2zzvZ
rUnMRVkkjaDU2ZkgzPaL8/zwConb1emB10udPeLT31K5Gb01ghvEolC4cT44Aw/q
RalLm2+tYAFbTcNy0JLomuwMRUiDPTP7/keuY2fprEcbaMeIG75SLfhx3maNjzMM
4re6WFBKVAgnONJ9q/is/DdTWF4xWEf0H3QVYzzuEdB5EWkvTS20nTWawZu3g+iS
7MmAJ00JCKLoZpmEzZk0TmLnSQ6FzNw61KbbW6IKp+nHiN3Ku/AQY4/GKNFewGX5
Jy4U4QI5N8yYs/eef4yDv7mkVKrK7zXWhLp+RMLvjAXXuJagCTNCdJ5ktksTsVf8
WkdZy/KqemXKwumzSRr9jXzDkgLCu8M4Z9/u71ZBytVe/1t/wBnzNPlCh6KH/lrn
MLKWA+/rApKujJHfjr4GvO4uP2/NpeGe9bD+hIf/KRumAlfG37l7o2mG0OlBjdqr
uKUIOmuYhaC4eWxpI0C971rZv9YoYR8B4HfCRUvtVJ276cyu3P9BPPUY7G0BI9+E
O6mNkcMB0+rnwaFUCiBqeuUty2pm/0OFAyS+WuqkRYDxFmdgsTkkGP+CQ6bV5bG8
cCZJTcHSGjDLSXPZ7/+hw7Br6S4SdLgddcltfddfBDaXQnY+DtA7w6QFyPK7AuBk
Qwqfhf+DlNsDw1qvWLjDUq3ircuQU0NvbLqHqSWuXX2OLnKCNXiqNb06cckzLlT8
o3TKEuHEyf8FIzg7n7cbS701QlRo7IRJ/8WzCa6jpyChI9+qNBG5/czCFwLT1kKX
1pnKZ4lmCQlqlekfY+0oHvm/NlMaLS8a34FY9rtMS23cuZIdcVxj1smdgKdimSco
i2rbhjiUGGQfEQvn54rCrg+7UjkKUMjEo2kaERSHcNJRgmAmwM7+z4Y0OsDVQt5+
8zSYzTeFOXE3aMhTq3uOtE6vyC3Qp5g7MlBMtBvYd+CoH9/k0XCAGl3wOK7LmfSS
e04u0P9D91Eqx3LzWkpP0nsjN6HR6pi45YPiqXLOp8oMngNGSjRKJWArqnjXrnFD
Y4QrpnOlw7vle8zQBmu9B3IIEtDCryTNWGwUJ7TAXxcN1aN9dmgAAXm98mIQqgJM
j2ryMFIhoFDZj1QqqjKLstQkeLy94VvX6wVy/AnleacFlt6IAW2pzvf8YySQW+Yr
+uy1J+h95FXjtJ1nEYphhlSVq2MD5yHv2tyixi4gn2BWywt8Ky7yMz8bfvuNokZW
xTYj42C0hHpT5cueSP+dMpYtQkL4Eme7IPgJOR2EFKW1V5kiglyLOdaZ+dLnLSEH
lWEEMadxcuof9UAOHqKIhnIjnr5JHX7z25z8qGqJqBW2sVq8OW9TjR/Kpv4nbBmf
5n3vlGXmxTLjfSY7kILAgssHjh8bC6zwqeZgiDp4eLGN6V5JGlDFR+3sJavXWgZf
ZxmSUGCrgY825aCIjP7KKLAn/0NNJGWKzA9aixpilft42ZLMJNdpCK6zU33gTYez
0sUvEpqKktvr1QfAcmAnedPoUYmC7F1obT0haqjtTAwDMifGKDrGpwzAU/mg4pSh
mzVxewPc3TGW//SBaKXOYTyKP9ahNzJuQ208QWXjX+lzfT8gZbIJ5ooP3Cc94KPo
O09zbj9gvs3uCuIzLzRkm+Gu+FQgNSI1uK7UIpTQfCs4zKyz47tFGbLtZf+/gu1P
QwYjceejS8geu/b+zx4pUZhqO+fxXtUnpham8Yf5jketXGYf+FVVg42YsUgmvtMU
SCt2w1HswdU6WZGpU3cOCGp0u6yOINqeev0bTwVvUcP8f1A3yZacmXvWxjeWIzcx
G0297S2HPT6hRan5qTeyPNiaMhHucc1gVtl5wm5iOND4WdxjGGrycX/l/4Y9xoVl
WhgHi2R/ZGcEZrhzjCa4UeIRLScW5gv7skSn+ttJDLGA4ciMr0gULOJB4N3DixZb
SFyST305CQJJRaIN/1AWcsFs+LS8KzbxyXMs1KkQBI8DeBXW9x1JceaWr/dB5PMP
v/bCJdB5y/yYmIXW4NWqy08qhzp+ULrxJWRfg/1TYC2qQrFrJViUF70btnOiWEpq
eZ3JD8Gpg8ktyhbaG6UDdoN4nS4E9SMqpieXND/V7IGAi35Hm28I1oudHJtm97g9
II6CFz/9ntvyDzpzoM/pchtPq7mvflb7ME00dmOG1LbEY95qXePVPWaOn0MphRSh
C6C7cmoQh0z97f+FOKb1Hn6s2LRP0gDlAcH2q2KzsAe6lbW49KzVdpt84bdYgrf1
SzJHNu5p+jz2bSVfoH75Dh5yWiMuumpIpfMKb3cjMXRcqLsHzbU7EGUYyyjHBj8g
qzyOSwlUKHh+e0Z37xZGaQjPlTemg6hYWYWE8UbXQLLbIfWytkJegaTod74RsrhU
4YyWpN5R82itVOmBZOju0JYmdHZvJ4lAfqzBmJa4pbiwr56T+/GINgHg4NUkjNx7
hhBnRVko2aVP1n5i6bLJRyvCiixCukjbzZ6UZQMrIFfBVRBj7g2DOzxrCyEmumyx
BRC2MCjKonYEogvb3OQ0ZubqCpzcsMeo+WAimYTXgWdpXgWMfYSb4QAUGgjDGjGj
kgsfY+ADSYU1/HCHPSbam/JkrVBMWjr/+Njj3FCbA0jFflRxt24923SAXyGSR65c
eRZnysnZeD7gKeBhkkEqHL6nMbcKPSVNh0wMix5O/86cJ1g+fl1io7WGY2l7BYMH
OTGSNCnSVb7y7QSD5Et1eWuQ7CXl9wHO8x8qDoR/kVuCbYEYZGzn207eN/4jT0N3
z9p3l1RnyEXzRjNYMhpZR6LPpEYV7P3vph2AmKbiZ/povS5oAPweFlsvCnQCTbpt
yXhOkqdtKIyJNiAShc4y2IKIMYyQLUjs7wKttfChYxOxnbZjoLSzOIGZT4cgMLRP
70JYGpqKt/GIf6kc/sc+9/nd+zR9fOBpR7XI1hOG5mbBZctaRPFZru3+y799mzbK
N/OVBcuZD0ylokh2OJY2Zah4S21ZBL9QSFiKB1rbuBK+sdzyB4u8n2huI0hD7Nl7
mEA5ZorW0boRSkbsnEZefznsiqwW8kEcNPVaEX3YXTUuFtXAAijPGbIwouKK5qxj
cIhvc6mw0/QkLAr/CiLqjBlTb0u/6+9lo9DkdQXGKvXi4QEn4F2WVoI69E//nAXF
T2DF8hfZdp4j7/M1thMLfelYl4Vank6cKmZleJM7Cbmpr5zMZ9u0kfflr+K2musf
gZ0p4CPPhtlR/1lu/Ih3cIHYT72Vj1eLPvQXw27M9USm2O/OWh6V+D9Wd9mBj39C
IxOcdKn649fA7CbzaAdtPkcp5q8kARygnwCMaHSRrXl3ls4EupmIPwgqhy+U0fkx
45KG7sl/Ac58PDXVDW2bg4HzJhfhOiN3SBspYN0Ta86UO9aBmJ4iISkXgLY28FHj
YsYDID+5d/0XNJZyWwW3lu+EME0qaBHqGcwbHFw2itTc5zEn4dtSUDTQEkKKZJtr
slkszaVgSe7C5vzRvESRmoqQAtXwS1ooJ43NlPp9Kxp1gUra0LVH8o3HXDCv/ii8
sh6njgdCTT0rAx8A/jzarvhsCtemhjTpVcKjZ3MZlk6Oi6y40f+WHf7vBzED0ZpS
yUlmVfcnjaI75GtxrvBdaeCDCYNyJFvOFoQ6GeOZiEzd8q3QN1LmBHKsHa6Y2mgG
uUJvPqeppOqWNKP4m/Ah7DXiErky+gOUqqDkWascEGVed2ZCsz4zq3nMpcCeU5FS
2jyecfRQh74GCmaK5hoGdwaB1FU+/QEcnCD8lHJUS/lhiLcru61uxRpu7UBhsCvq
WF83vtwrW5OIECWZw4z+UQ4oGHpSyX3ziruDNZlH0Ygvf6KaAEcqPwlcB33AtEBD
eT152FObvjm3AGe4BO7RgXQ7YEts3hQonOv4eGp0Fk3YsRvVIi/uZPqNln2CLD2w
5DKqtDfLg3CZzW1LHpn4flFXGEOwtbGbmEtHwLxWJZLOxP+ouLVSEFiF+YzIt+y0
yztfUv7730/njobAi4mSa74dApZmhmToz/D5vwgEwB0skFFETsXwQEnBl8G+VLuC
ZXfufy2BMc91tHj0nqti70R3GPpi42ejpnT8nsiEACCN9euC1rA85ZYlCgQ5Nr5J
nY2ms0ISbhaLCr3DeNP68f89tMu20Vj1Pyb/Nv6DTJolUmB43C8UKlUpro39hCzv
QYrNANZZ63h7+pLCKDIc5kIrRDxAwC3V/iOvkcKyfBERwCzAeg2yxTxS/9SKbFTn
4JkRtbwtwivCzEYUkIGkmp/YTJIRRx/eT4Gq/05p+B2Klgl2UKaL4CJUMSFbTKyg
7nK22GnEgR/Xm3QSjJA5YGdUKJ+ThSa3jZu/6MEdm+n4K3TCtGRLCtWKGcEZROR2
D4T/LaJ2e/aUb5fPfV3wxFeJY/pQxNVL2avgIQro2gz3t5CqTPBhOu3V6xw59Y+n
5aqIUvtDDKfPN52RT9ZPqw9RCxqS94NZc3/c2b9/YyjMYVYEeh/nAQTq4lc3b67J
fViVq69NVfxB8THNweT2Wt3usTPo+znlq/Aqj/TJZJiT0b1Ty40voEPNpfWkjUcE
iooyO1hDHBJu71XKVOJs8g6nz8qnH3C1vxhPzDyvltENpaVrypgQ/qFyC6dBE+Z0
4ZFewLJd5v6njjE46dxaPINRPNXI4PTnyGjBoG1slRtMZxm0xkZy3hne2avN6pQk
fuG8XT4kajpvHdQLPoXD3U9VuW/7YPztqgCf6PTse4xVfty1i1N/1r8vZFXH1xrO
AkzqYl5xqm7lH4VZ6cT1UfweNht8dxzIioj8d/x+3P1XSD2yt0a9HKqHEPFntAgt
mCX1uoET0xqV5rj9u6RZmOLpjkr9N7OPnYvPcH4mXkvO8wwQcJQgw9no4Mh5n8yg
aScXB7XzvcV/d8iXz92WlSjn3y/4gWk9Z7uL6TmZ/nKqc8Pm9M9f/PQcgGOElda/
4YBe/lZ/wELCSOBFYpWsdJXdvWbedY7yy3NSGOoLehdxZPx/lATXRE7wZuXrHnRG
fMbdwQlinUd7P8WWkSXf7ZCe1Rkn+D1kgttoFP53uXABBiDStenqjwvl3N87hLIB
aiNaq1EbCN3fF5J02Mm16WczYjZ37an/p7e+EZ+ubwgfF7SD72wW/RJ2+aFa1NaJ
jeNditbLh+IjaJa4qdIK6osMG87sh16p9Z/hNC30pOFwnoc/lEognp6DoMy9HxcX
kj+yCThfVGL+YXvkQY2PxAtNbjBZorb8dWBcyPKi6G8qCJ379H2EeLxBnJ5AGDD1
jI2nwTJVqQYP0/zaqI3NTP0swnEgH/pi7FZ09gifTtzb2bXpkWh2GT+mjYkF27/+
0+aZA1ZoYieInLX2kzsVkk7MnOeCimVn88pOL0b1gAleV5eYf/co7ubphMeQ9mA3
TJaiLHr7IinF4WMG4D9cgVmRuC5P2jN/zSgoHZHhwg4aHrlZ4D1gMdB7imK2eQJg
ZwETIBCwmIIh8Mqhii4rcvnxD06OdIHH6ql0P/CmyV7AdJli5djYGMFs+bIwCNfz
EqXpp+wq3E3+wli0gTpJIIiYFH3V48zsapfpm5ESh4ZNc2cWJ4UgTmTZjpWQi4o1
p7HyTN88DgvBrWpyyz9PlV4O24/1731Vuv9CTH++hdFUmfyhrFpSbCxfAiH5Wjc7
qAgFiIyh/10EsFOX7LTw/v88J7BOe0AndUcVlu4z7vWH6q07i4aIsjEpm1l48Buh
aq19JDDD2F7UdmY8f1jZCqmSly0sp161CPcVQDZOM+sjUJRgIQLufYd7C8DJn8Hi
BE3VYPv2VfQ4XXx1SLxOwV00I1OSAvr8QRU8F4J29UHIz3QlFBHy74fA85MNBACs
g3ZHMS6G3vOKtx5CtUvV8K3OX8/lR0OyvlXHc9eMh3Wg/0xDPCLKzZDnNlmbEt+p
uKkZU6rR78jhfaf/sWqHIHYyA0C0y4E0ngFeIH1FV6kn287YXf0o8UrYXAIayWOz
EJk+Z0gRfK5VRRe9A1dmR0QMeKiI4P92s8BjIyYYBre6V8FMCYlZNfx2ErG1OwQR
gYjHCZ7ilWUZClsEqnnUmsyCGuGs2YHLj3xTRFNT/4JE8k1TFEFFuIESFBrSzzeM
fdCeJgCotSoQHdI/I5dbFl64IjLPRDAqYvv0OzFNR02NLp30XdQsQtXMxMmw3pdq
/e/WEDVZ2XLnIcq1qB5VlE+apIdfV6pJ4N01tmya3Irz7ZZrUNtb3W4o0cEU1bGY
ysInOXdA+9Q3lsdTJghtAm2BnP25Bb56j9gmXJG6tSudtgQhiQWdlKjyyXJZkavG
NQ4by4B5qy2qErb7/i/ssqrOMaqjTFS0nHUe4BNy7BxvbhgAhdKtwfgE9t81NEqr
7Yr60ztqRlzzjxHesdFl4Ut5jq5TVkImA4zFSf2DsdGC3wYja++QzGTBEaSLHcoI
N/FZ6/O703v2tXcHw60D7pb1/2gTE74FIaf3V4c5srA9UX8GoVtI2NUn8Qk4Hq8a
NC79VNPvSUu/BjHgtC9Gy6nkfMlbTA01/Yk6uYKgPrLsT1W8GsQhRkRYTTHwt4DM
LqjlV1RDPDlF5iOjtSeKDYG/FIQJ3I5sGkfFUgrt9zNwavN++U2L/QTwAS+emVVN
T8cO/BFxKBnGJOa/7ZTjCkxmfVXJqJoYpGnA8NyjayEhCz4xJarQ7DZtBTLjSScX
L/djAOweZxtZ9b8uAW+GlCOv95GUsWCpMiZhYO6o5sWcTlx11k+IOKhjSV/WZaeX
W7/DUUGR3Ti840BsQQagIcg32N8Gb3kYh7IimuT6getT1whU2WBNjYd5CspnMCBv
deUlF5wIOqA7HU+55T9BvjYAMZOWJjv7SEJ/FFD2nHU6bGsGUPngAnpc28xUL3mY
VeSgPkl6tkNyzUtjy/bqlIlJQLV7b28y0I4aKh3uY9tTmsyWZMos8kygWFtBdpvD
YsdxgFYeKLT+3ZEMkWeRM9p1qlI/rG7MX6sc3NIL0aGNFdUyERSbWXiWq8omB5Cz
fPlk7aIbaaSL8FnBJI+ghdZKWn+fJWUc0XU0I9YbzpD/qLRDUesfvCu7mpJIwdrQ
DSMweUFKK2mZc/lgZsK0gzRbdEoGO9bczFLtct2rzqOr1OA7B2xebh8mynmS+FLf
gzzyxWKXONPMet/OExgm83KcBDZE1NaVO7g+IorDwj8Yx70qE7kbSeYL+1D1ci3L
1I56VYCaNKlk3riDKP/zWP2rSvTJ7Br+uYz2AHqrkxVtF8k6NwSFLWLsf4eRxo0t
B6j4dkXRR5qXl/3mvnijFo4noMnoNHV+4BDxj8p+mOl+aKyIMKj2j+oZfXNgNJyq
Qmr++sSimFxIqb2w6sLj4O5Rxt3lBIJ0potvh6aoBaorMWbC5/jY1cYnNcoaETTq
2RSBzkfAWKEUBClF99cvRyjcb4NzcOoZKUqonsntoVP5coBQ/OYPZHSx7PyRf6qb
0tc0wbGRPv1lljEd0RRZGGLY+Pzo9SStnIXor9V56SjTwRLzFU4rmzIIfz+vfcQs
rrFiPJWQdZmIIbmPmrTkPi4WI5kmw6AMtUOB3pwC2ofKYC4fle+A/AKILJ8BTP/w
PSa42sMFtpRBwU9oNC6/6nyvCPOmzDbnjaivDAIsK47R0/gGaNJgkTgvYoH+wdmX
65tJLV463J3mnfqrGlpdSLfnwKNEXkX3ccsWqHvHn6e9kVaf8I8qFe/lQNA67IKz
qU8OkfWX67lAsiBvqwcvM5QSSg0VLc1KpOgBmz/OA7RTsuwdr7n73pGUabcnLPRA
EHWWU8ZV7Uk182MyKaN9q1ek/QEmtT1a/W7yTRUM6qcQkft5ZQbWOnn3yDH5ehCW
XdYD9unVRRYPipLQZ9TeIW54S6Bk4WD70WONxUyDysrRspqXwrvOX1x/t+caNbxu
IstJ5ArbHasIp7X0xkNntwAUDBrFMqyGZpXPrJMsD4PnjvlGrWaQe0dfJMvom2so
ZfMvZR2OpSYzJ9Ltjhd5Q4JmGdfdy6i1Q0g6Gq/GdQVgSqxjo7JTXoK0NBkOmL0o
EdXp0zId+A6psc1aaKuHJYO0W7mrnscG0SPmMbznS5t1IS8Qz7F60i5MgEsVIYwk
X29SlbsYa8/fGMi5+hjcHIE9Wz4FjP5/zWtkIqEIojs0q9Wi7nV33I1+D5jz4CBC
reo7sytrFzcoWpHUeGeS6R/r6yb7idTst0ypOf4aK/1vDBSyW45gKqTuWTQ1apI8
Cx0T4uGMl6RYWrQgSHb9nRNj0mP3MWZ7sYljLLdk2jM+z8Td246flfbCTiewF8DK
7AF/husGTq66GOFDXNuCPk2Yh5m5ht4H7sWwN7i7s1F+Z+Yd2017JLO0NjLR393H
MBLgJpjDaZFftsbUdZfiPJm12l/3ZXQ4c33+FJuu0NPz1z6R8X865jaG28iyE7Lw
qW2ST3HXMWvx3Rzvtjm6zwFUyA4F6WDs5BrHhogEKJp0XGGp3ciD9GFVRPwd8G8M
qCA12LlD6kYMyA/Ixyn0V5mudgm3H1vQ1mz7E87YfRfDNmpn/kAwZA1D7OKNdF+W
s0EsxMVQMN/CICArsVpbiCkusqMaQIsieQ2e2fLj6xmZY2h/cvfucnTiLAZRzjZL
4Wl0f+3WIbehbSbmZ6xjXt5odUJwwFflXuLmVXhFcHTHamdPr7vdUDVbTGhf34Hf
CQRJAg5zrCLKmTsTRy/DORO17i+AWRmxedvTqs3xXIMC7EuhgSi1J5Aa8vdPBP1G
gXI2CmyNwAhDjtscEdNegE8LeeWP5sT2ZRFRfsZN1/eE8bYPeMQezoyrtMv1Q+Dj
Y3UBnR8f4IfGwjONpyPjxwU4t1j/GZ0Ep/PAi+d6SOuuPiwALqTANXdUvD0q3ayQ
Tjals4jU4kufp94glXhWEpihfBdeLodYRxs0WUaICuNS5otwHqCCEqwXCRxXaFrP
H0LXmzvLLJSJ82/n4UHI7o4TPnZDjFiMSRsPncaWjOdCVx7YYA+aPWpuuIozIBKi
46AnAK3Snxrap079SsHfUCO0uqQUYZVJd9IwefX33y/rrWMZAzAnJL0Mv8glCHJh
Axdbr3EFWL8Fplk9SNUzpo5XLgbKfZkMNKyAyGE9oAXmssNJzPvGKwCjvI0uH8i9
i8z0dtEAeTnB0WPO8/NwDyxELK3oBXWqrF9yMjR2cxFHjUpTNy7SfN6zJyy3BFWF
ncXgXvPTxMswXNhz9OwbL1iYbM5w17ftvLC0vwEixennY0dEW6hK1E4Jyfyg7Pin
7+tWvnN4rca9onMeRfh/hOEV7rfIFqNoysWw3Dv56So0ZzBCNVCieTzKM6+83C1A
NBggNeXzb2WkRoYJQXZGch3I6kTEBLjR0WRLsrVruKkdHR8g1sKVkUyhTIyO88fP
+fJ7oh9in1cFIrPSFkBzJbmKmJrxPBFcA3ShqFeZ0SJLWMo7JnOqItj+Y1tLOwWr
stz4RjyGCJqqlA1j1r45d0CH3QKxdOalWgQGpSGHUlAJYl1UuxlC9qeV5Dft3U4j
BODJra+/mAQ27oNMEVu0EmBErRdQedckyqByzmwQI/vmgORZKfFO7bux8rFzofSd
1DX01qz9cbP9F8geB76nHLZ7/oAmHbo2FiYXe/IOGsxUdMRqrq4hRz3bxRGDXCOr
V+0i9/LBrIrYLd2U8uc8o/3egRguPNbArWrn8VtuTQqlbq3nYK/la8ZTl+5SwYPk
lOFjXA49kR2t3sKwT6x1V/jK/zqm5wl3QMgar8SlgHL/6u1Yhcg00MT2oIx5ESCY
o8gPxBjOocWp1dOVYtBSo+bQyN2Dcqw0F1MEbLUgB14mUG1BC61rpqypAl/EWTmU
u3tvgmDSBLCxuwtMekzoTCnClUNY4u0pxa10gk44KnuNOqBIMxKuTH9HRRxQfrZM
PW+ITVcdfhkqQhT7bGfndvEMADcOVXlN4w9LJ7nrtAbjX+yAxRHjBxNsy0CrpvPs
XlmiFMFp34aDhrUN0a4zS+C7wFcwCsCrupi9LJFcQPMMPwMrZxBVeHBBAl+IUUNY
HYEREqRfBfTcnwXpMT2jVaZBcsh2eHhj8enEbqlZ5iDvvh37lM6YsejgRAGvVA5P
468HFh8GTjW9PZqzlVUd4WvYMl+jMbJi052LEK9iCVeFPTSqiY2xVXN8tn7qIIk8
me7N16gCmatuemFkDeTCDtp4dOV/pAil05fC4oW5fg3p8/4EQw91x6Jj7w6Rgp5S
gkFVg8SWxGhBkL6Y65Q3K62i50QQc1DIxrlVMOsVHt8tgPXgJSwFqNJd83hg8J/J
S+MntcBw69N28BFqn3BbXUiu4/YKr985NNZW+LKy1Z62saFuVS5BZzg/NYJrvqdN
gBrx3kI5sDtAPOiXay7muR+THPwBYnjppvjoBS5VVCyMwzaHob4EHY3Me3vjBGFR
r4VDdkGmCdSrG7veY5JS5mvX1QHGIjwUF91oLSKmmJOZzSwBivzwTJRmp466LOiT
Zz1YV/NO5wjOGfH3uVJTxf3oab0bPm6Tp6W4JlVM35xG79PqoYAM9WAvQRE/Jz9C
V3Q/AH92+3j5p6u6nUlIKvVyQzKBNYeMBT7+IiUZXEMje/94V/pc0vDT89YWmsSt
99/Sd8D1LmdOFgnqP2R2hnGjdyS+ICvbKVwanzujKcY6gJ+5vZiPEDN0ga3rL5hf
Jt/OM+1m4vhTWByqqG/11TfXeCdtwhjpmVW9xg5wXJr0ALyLBQkQk7SziHu9IHix
wEeCbgdm89Kv7gNbHU7aAtf/ZVN6GLjlfwG3rmZfPx812lYoiYF95nvyeiQKKvlF
Scj6CscOwo9tpYALkCNUwSN/1m+yfJQB/oYQQTvN/XDEvpnOtSbnLHF/UOeqorO8
qb4rFxB9Vb3MBJNuX2pDPAYl1CUfAQB2DgS42uefjYosVQslBd/+ckmX0E7u0eiy
9TfvactJgrLfhqxYenaXO+BVT60HATyCkZK6RUAPwhH3KabN6WT6O/2OFjfkVlif
9/kzJRi0JPks+MWN28gQ6YK6TtA2VrT+XA7XwLPvDAEBTTBhIK9iG/btN35hNVNf
lhsHKAxwVvGGsu+gCV51PvXubuuzlAld66YFnm6vp3phVp8w6DX0GZ81/t3tkRce
ghNkAxG7CfvQQHbdIg+j4aNsQdzHCVSBfXntGscyl747VclO95JrADvyGxAX+AnT
Jo/290wzOsHPL4r+pNogzb9XJxmuK2WOe70wE0occT7+4FAsd3tFIW0II+tD2eBF
HhH7kX4hDZuZ4hIyMvxYF3exKwn5LV4nEZQMTU81b9x+c9Mxf3a+S23O1s1c7nxF
k659DiANi1zfGBrO98EjLPjno84bAScS79GE7ZX0Rbu9/ZEL/k1JT3nCtGeouyIi
az/fzageQ54o0gqxXRxmXbI+dLmzA9y0Cs4N7dvR2l0PlIEyG0XJjIy494BT56t8
rKc3s+I0gzytrdoJ8M4ZXg4g478RVOry9svEs7cOuTQUT/2qCBLwCs2bSm2tp/az
X5ntqWzOlFlczBA3KdGnsmINu5QukyTI1qCJoSg8T3Z0jtiFdcLmNHz1iqW2flsk
L0ca5emVIdH5fYSWy40g6A+Ba38GiM6a+TiqXizjYlHWZDdqydd1SwI8ln9EFKuR
P9erHvjhmXgIFwQU28KlJzZU1dC9BfOb5koOH46YmiWUAOGunK3bgKNz3p1jpckO
ofHtAnx9vuORvD8WuxOkmpGhZb0RUva6ih1CPwCfE2V0jW+BSbiPklcPGo4noze8
wHbp13YCj1VG+NDsE5lCDUE+U+eu3o+1B294+49TzOtAyQzh0tN3QZ21zxglbIMc
GpBuNmIc2SlCSoSjXcOYyHSATYw6z+WKAR48I5zAMUVYAUrb1nlv2cptu55ZNgrw
IALL/cFm0YHroo6D7NhUzgyZltSRMOFnGpVh+qdO+/x4E9/xwvuKzpyVWbx40Xma
JZOR1lYYV3H2rRg55Y/jyXgJ+QfphHUVxTJ/OzdDqf/An51FK+fq8+RwpYCdJ6Wh
kvcKGsZY19wOA8v0mHYSTW9o8y+z9ssU5NxE5Zxx3ne9Lx/LVfvHwEk9RtXpvtix
cPi2MQPv/YhpkiM48qEC2R5oSqJ7kc7yn604YtemLwmEISdhUKeO70Jj7tb2p9zt
jg9z/jRiK2WxAXENX/3NLtyfKPy/DVPr/oGzxkOqir3nmk7LgVW9C8vJPP02rI3h
QvNXW8KUq+jMlTqSXH9BGs7B4z7yHDO2zha/KZ2l4RC/APsyyV5C7zgc795ayP5L
7lKyf8myrNUfMQihRGtg8yuP6VUtCnfcIjhDPZh0oBK8tcLWYh0ItUZVJJmqSZ3/
av7CyjPt+yngYF4omPwA0c6xPQciwhqYI0CwC3TW+l7H21TJ/ZOFvuGnNBqMgQLm
LLtYqA1a7fI44uow6tQosD6yEicSgwaZbKdVT3FRfg8jjkKw44BxncqhV1ztlY7b
sgrN1TSGRRw7Svpkdypx0XEAM7cOy1k6mByMijIWerKcFblsMdI+xN8MykixUhHq
+WhewdFNmMPR6xacI7Jov6PitfZGtr/QWaNS2EjW2pcbReLT4dW02GN6cD92FSl3
H5uj1zGumEJBY5YR/movLVUUFc4Fm0MWmUrcJftGZk/A1/BZEVr5Smxrp5e4FvmC
QCypgmslHhomH8pjdV4z6SxvvbtS7i7eLUhZ5GslwP0ttCnZMF1izTyMGY9JHTVH
F/jpUurWLGfGLb0mrusrIV75SaSKblX4FCQ2gJL43wh+vD3QZoAK5VLFwOQm+wKV
DQ0OIo5ZBuk0jRJ/Io1OfM1pJgVbML4BeFv2Z2OlE+JuW7rFVwFgBgZi9NTpZ0eo
2mWY0QZMACBMWx+Jaj9rBJ6T5nrjQGcoL8bJs4AonqqTFLB9luUei8pk6NU/Zein
FWlCXOlq4+kUjijCbTKwykRdpa8QnSaxhiIuW8+CuBKUCZE7MiOEZycmnK5g1Pln
Y4FCMBM2weQThQDWw8bRZjzpkFT4XBlzIlUzfmADQ6NYOnXOQCE2MqkqhAxoZm5j
YcA/GBdhbAL2SNxQP42c4SgIlY8K5DHJ8c116NX4aRDqEi37Q3G6Lnb3npUjKZcT
gHAsElRLHkVyukr2qsHJIKr6GLEgjcZwZHHudI4AQvj/d/zN+pdwjDnMf4vvKELx
zMO2M5DidNXg2EVJfX29WjXC2Lf8I1g8IjxbpE3O/GFNCTcDs5nw1Sv7wJqf7gE6
HCyqJWQIsbeXn1SxCruj4C6z4QwMWZjWbZSDWg4VTmvtc11yAU0aCnCXp3Uod/zP
225l8qTWrWbcr6KaVG4F0xon9FO/TieqSHz77NJqqLpu4SNw46wmjUCru+hBOBiY
fFcMvU+Ykr32fHeBr5oUnjezmh9ugMXL7d6CA4xjpuytnrwLtmoC3ZoRkQBIDn+H
hi8Y2kiDgUOTrxxIGmzlLg/vRz0FHE1UsoJBOd73+h9OR/LpCpL6S59ButfJrLc8
1d7TDWU3jFCplcklA8kVCXFUqQAYVJofaMMJto7feIyAQTjUBC99b4CnFHOGu2Ev
LZ5Oqz4eOVQVqTkb4yY2FH8NgZnDAnr3OoohZWkzhNbIrPFqfpNe/3K+edOLhp9Z
u39uG1LnFKqYzFzSm8XRcfGJOKkZiV81y6XzXVnuKt7SBvRy3kprkVU/onG1ml/W
wFGOebcAuPEfaJ/3hVcrE3Fih1PcwVbbWDi+JpBQe81xAY5WJ+BDnbSDbnG39GLH
BdVR0NijXJvyroYIyN7jLvlV2TwRPDiKM96UghCq5nrAI+VbuunoKJAMEOmJ4Qzc
XomzUed8vWwSe+E6C43igFADdLJjhH455NztwAN3Lcansc4AzvLZk8+1e/LlZHYQ
RUgrYaNzXl5w3Tqctxha0lC/pkB6TCOcYLxFP6He3nBa/bgb9KUXrsky6yG/N3ae
+6qoBak+d+ihaVBgZtY2MTCC5BXMbWqUTCjQCYp8anX3Yik8xLC/Vi2wunc8gnX/
4PQI9gM6D12iT56JqrYj5Nm96Z36Hl1GJYaMq4Zgk38Skz2m1Z3r0fNYJoSHCVkD
R2gSMcE0CHFA3aW/Vjt/ntQPUkGLc+OhxWR4TAIf4p4x0B8DVQDy6hRmd7HCdWdf
2e8Iz/jOWrRc/okOiTN0MuNND3PHVsUAfR7nFJiDu2zyObc7MfqX3fG/Xvjy4zXv
c2MDazIBMKfaCVujzZSSBEzTku/FAtnGDEKhgXF23Ml4sRo33+ahLOMNCHX+H82R
4FCEqAEDP63LSjAr0dr5rAQehlsmTuHVuGLSKTDBOoJ3544PNMR0EwyOMvVQHMtr
ozrJRJ4RTTmn6oilvvgnYEY7M0zM1xFh69LZ/DzHB9kziXHmoOZEq0AY/X2UVfgW
yYlL7A2Ti4GDQw/MFqjlORZ+lO/UQNES4Sk1lSTn5cX88feSX0v2iRNmjx5Z6r+W
D/BGhiqn/UJoyUB4O7KD9rz/QVHhYJVaqc17SXmUeh7sQ2JKktRmwHr1T7UHJ3nZ
CwQ4erIq4R3MjlwhMP1ZzMj9bUpUjRC3azdy5OYlqG7M+TEEllICrc1lDvw47k0H
uJRxvIjPecheC21FFPru/Php9aZrWQNGb0k5caw/Ou0EdGT5JBByXsV+jjkn/Yr5
itZ6C4w8pv5YEhpqukqroPdtPwGLl7eOmfTiBXyxnpcUZZtlmUybmcYmTtPGjTQs
LHCfJcRWZKg+zcRI7sYI4bfYa/fCoW2dWU3S1jSS75FrCI4AAF8PMSbRA8fHWGBR
3a6VIQeJV3xja3y2EDWWSxxoH0P/tYi4j6F1EBJWRuUBgJhV/fH2qFVJSMlD4MC3
wiQfHZ11bafSUVSNOyTQEhbDEAuLoxMBbS1rRwJWrn98rxQGpkhqO/L51Uz9Ylgy
9YyE1QkdUNj/4FUYPSaeVF5AKTtpSNdfNbbW4eUWEHU0vUDd9SiUy50ND7fmRJLv
WCo5KnFTi5l5eA6iaRTmCYh9cQE1Qj9jHwYepVFoxvLAruhton8trGsujtlKVtny
bhx86WOq42Tc/x7M0BNcrDJEuhtJGPW42mET7zDXXOi4C/KLjXI7KrTB1oFjUdjM
X5fmV8MPbF7Gb5Y/gY/Pfhc/ULToYN+dMwZcpnXY9mfMcuKv8x33NaP9eB5HT3s6
rIfl/6jUYBg8j35bOkq4XAJAOkwKX1vobVt5tbOgip1ITHDfCtaBHLaL+XooD/DB
NWnhy0YSspvYThRvKlsBbCp7E4JT8UbgGPs4RfrG+Aq8Xr3cBKjtHCdyN8qDxIM9
k3x6GiBD5RFnqwye9/EFXUP+Cu5ZDQ1IyOqHR9obQ0iJE+FW1nUYCx7XTSk+LSR8
Kv2YxkkSUYSxk0EEjOSE+l3B+mvw0M1SM1EEkWDpyRM5NabuerqNsvWaVzOtTfIX
EuH4udBy39skYvZzuy1wg3jJZDQ7fwuiH3F8IJcEfqzHBNFrLffQFPRcckCsqf6Q
KwCXsK6gvQf3zAIiKKETC43xC65oDDo+/kfEKWCB/LAYb8ckkzJR7fij2oC9yPur
LdAHvjFqBb+KeDU4dYqtwtP9jhpXKLvB5yHIMVwdK2C6c01vEEvkjG4ic2zNjmfa
UAQVlTWmZnHcO9gC7xBTQ+lW0LXomTCRPSc7i+w+OIqfKj089Y/esneo5tejHvRZ
L5OzwF8L4tSyzMt4+T7tL1DJYQa+3VzG8zeeQxwrPIm0+gkdZnbhtuhovU8zGCPb
nRvcqj5XFGhZ1B2vdPeak4/LSVR8/g69alploBXjxcyiX0p0VJYIkDeugkzJ389T
4wPY/mc6/6Wt84WA9EVHpEepqh5DNQTm3vqrDKt4TNcQbBs4LLMIyCZqqnGmHqsS
OImGnxEeJZ1vf3ucEZJDvPFbDQkIuVNMSBG14LaMC6n07/Pd26wmhB027q/VSZtq
vUUxTJZlh1JO8/r+7SadPdmnIw7/m+MYcPwgF4jq8WbSjF4NYwVNn6rMQCzKTYV9
J0z5U2//e+sny8JVr6u3DgIq9ChPL5XaBLEWmX0/qqHtTA2BacryWyLiIxArCfmv
M2clQFCbqX3BozAEtx/BTzC+hMTBFeY5LFcoxuozrqMjwtaV3EzGZL/aa5hxyASE
wdOMw+XHMvj9gvUYEbHDctQmc1jpe2CZTUPw7M5XfAhB06LK6l7z3zQ0LdhNQeXv
ZvOd+6PcxjABNWRkOp7RG3ctv+/slDqGwQBpuewzASA8Vm1PEftI44GUbIlPRQdW
UWxbqta903Stew1pAt9zdMh9pRDxfZBe8mwyhI1URMBCAJguMN8+rFUCBoWgwgtc
WouclBPyU+aZ716fwYIkcs6nicMKOiwgawGmLjGFdAEtB9xuXcngLtHshR1YhwLw
jQ5IO73X43aiMRj4dvuZXCQxI3YfaPH5CEZUNFWJTX3CpJZTS8rFJxszwjq2uuUa
zMIekOr9Wi4qpV8YmpJzHStWsTZvCzfBDTgrSvFiRFIH2KY8j86uz7bf7BvlBcrO
SQhnLaosXGFZtEKU0TxspS66P63gp/DVOEosTppA5MSr3ZBSzFHv3QyPCJxt/PPK
7xves9rY1OZPsp1mSMU+VUxji6ldM5qNvbiY1EtDoDdfjgKlbxg2Tu2c80Sfwd9+
OZMn/sPGpPxmbihIYJFWAlH4b4rl23oJf35VjYdIQFI5zO7a5wJ7ig+hvFWp+sLd
OY1/jP/DhNreQCbtQhC67Qiy6LPiLbyVnJIglkFmzHla3nKmTXeDR+bM9KXHUHyt
zyFJAQ4ThgatIgzhvFSC//Ar7FR0iVx8+iGabiieTqpivp8S3hkKIl1UBnMW3BJm
REmHg9uvvVCGkGSOkRgti2fJWt8aIcfwU6f5g1bfV58mAprkB+SHwHm6wdcOXhuQ
jCJw06ScTlfdoHfFdB1nCTtGEpYBclY9T+YlXdijMZAkrnLRXCCCAc63a9wegKQs
bDcI8iJOtHv8toVC4IEQH7jrJyfskOLu1JhCRwVOXT36fiJZg6PBfsSEio69BM/q
vOEbUHeptxYGFklMKPmlZ1G3flvSU4KsZAFNziSNYpzPrNgbWVWlUj/oZGV1SrjR
1hl7uz635GseBedoFbQr6DCtc7e9WgLQp26L0xZlW0d5M7FnQtIiM/CqXhsFl0Xs
XVniNNkDh8KJaem8/DK3li+Dfc0iyzyc2Qw0PZGqxVdwkrAKyaik5ae4MS4w9jI3
RoWJnO81sYcxScBPXIeCc9VDBSMJfUxeo4YC16SM7KLYSWkvl7P/VtadIpnTdhxA
y1j1ZhI8s5Onw9n5IZdTRJRjGpu75zLPlRtKtnT3Jr4yvA3ZyOuBsdm39iltA9yw
DmND/31hNXOfsTLDCUjZgq7Jj13K6efu//RtL0wotqU74V25YndJAV0VyAEM77mQ
KfnO8PX8J/WOzO3lj5z6Z6p7sYuD7KPKAPIQXvnNN8fjlF8k0s/N1rKloNFF8gKS
XbRuce1/fQv9pitXyPzsaG1+1FDLjUjFclwZ6QyuhTQ0ZL9Gj9ArxohtmV+ehrND
Khu7TShGa+1/YhPxAzHnAats2MYT7eY5GfBViL0ogafgnMiGOBjMqg8j2SolMKs1
SKMAifPnxL26WN0WuKJYc95W8V4/aEutQfoIR4dT1O0syOQSkKBxMQGG1God9RBB
LP8t47qnxC5o4z/YPjc1JXFtPXkkw9CfC8yY3eAwTqNR+uSeXNIHe2BU4V93dif1
pbh9AY3lapRSy5Dpg0vCn6GRW9rVVePC0cp9nPGbiKj/KwYYWy0PvQoc+foJMsfW
Hw9x32xF8RAZWv1tmmh6C7SpO5xpcuL7LnJCFxhonKXlTzTwErOMczUi10Ut+mg0
KwV7XOuSerq0pd4QRw+uSORkA7qO8yF68b6vTaGE6DrBcRM4p7StaBOF+wCqzPbU
jQfqk99tZ4xVXBgfHZ0ad7dwdd4VP2fxMkzswKglEDIHlV0KZuI81D/vLz6TJauq
IbUo/ZnOdi7KZBHikekt2K293lJyluXpNcTVPoPA1l8BvG1Lv7HYv9Hzul7RYP3Q
2e/tgQXb5IB6Hja8kN9iHRxrX3AQSr7VxEh+yZ8hJWuvdSv4WgL0ksd2PYobpkhO
ZE+AX3C5oxIoalxuYILvKtpxPNZGRoBrAzrKBlAU0ruj/2HxVQzoZ/BtPry9waL1
DhT1TDkI4Bie+c0FcN0ZmTHg87rJViTeWr71xbI2qEAQhUmiCJUelrzuMoEr9Cq8
G/RVzLbVKz/o8g0c3IUcSVcS5E20Gu3G2ZS5VBhAHdA4fj4xXIJQCmH9gj2RmaIE
BBJXX53OwRjcThzsYLUenDOT9cxpU1cheA1UABeXI++PPcRb2vR66iHpkrUdP9Ul
Y/qwTktug6spetGv/NVpS+yQMtuVYaUI6DFrG567uwYUfPf5WpTfiVIGGmFSYQsm
sYkbOjbUfFDmORWxg0MCdroP3/SPyEDQmpEJtcRGudd3nWfnVNjruRROwPARvE2L
syzxvOL2G55XWS5w8XUdgklb+lmGVz6sxxJYmT4was+fizRd9FGRM4ZE+aumSdFz
EzjbBWTeU3pH8qXx2IBgqffpU+S9kXFynRCJKCQSLtI9s3Vd2pL4g2WTvy1iUKPF
qvaUkv+ouV8L2LsJGD+ipAtgDHPQvPmkOof8UL/2EynSEv/TdSEHN8yeOBYad4S/
JXwoy0NvdCWPVqRGhd9QeZSL/2EGD21iSKoidkgBJLmJgudfv7wJDrlq29YPZQBo
3QsDhTrwnXnlGrsxVPPvIWaZvml4gFbf7V8EDXz+10akkecyR6Ak0Dj7SoSjfDiy
dBYJDHzTpUSxH0+RvKm3NgUj6WXvrhBWw8O6NlVzXJyTHGCIJfeEBsv77vs/W8A1
xmBAR6FRH9COGxM6r8y3p2B9p/vF0Q0J6Q6KY3N8krzkxDcMRHtYtVypwF/drOPX
XekbMbiot7Y5wDMw5+aw1Ytg5o43NWFvSKhQWndFiAkxPUnMrFVkG4HDt2YnbvT7
69tuI8TaZgDhwqO/Az/JvrWRj/9dtN6fL+v5TalYTCilcj0n4iRivNIG/lHpaIWg
oCBgnwkgxbaEw3cndITU3PGHnC/RgvyfpZJsW8chByY/tQkHtcgx7zbyoOPrOSzX
lS2P4LWcYG52rkSqPSucPvKEEPf68iZvpSmPDeLuZAA9ylJJzsn2rK9xsvQO/GYn
+4ss7rBLqJmA/qJkWoJpYQqs6950wh/VQTQGcMSQTTyhvRqWM14zfl93wfdTXBYg
r2w2jS/LLe+rWTShuueZQWrCQuA5GCAVjyHlVnJz4PomkQdbAs/BeClEiFs3nk2r
XYcuh1oIh5m+7PmBVxAp76W9dEs+/3ODfC2NamaLnvhEGFQ+YW9eYVbbIaJhDiY5
gKJCTFvmUzuPnJFA+WMWe1vK31T4Io6Nma1UxpsyuRqlSUbovOaOVAbAe+mN8pP3
hLM0tOPwv6pFTdNxdZL1HhUo3QSvvngvZEl5jYgRboLXUmbSRMf+QJZTcevGElI9
bvdMUp8tA9FNkEG9Z9Tl26qAUB6/iKuGskhQzL/juNirxjtrzoTFmnnIZYdIswrU
RnTm2T4/N1PCWZo+BRAtyLboJaJfrRYZaNtBULraIbSe8uXe2NSmk45B1daUVDPJ
ox0QIpyGcy2in2B/q543o/7dH3BlFiA2XcWKS1oPsjTjEWaexV6Ij7dVYzFVUzUp
gdiWBdVX5BiSKCpY0DvvmIg96qIVkiCvoppMJoRPJoksNQmROiQGOjvEQbW/jtSZ
FvSd00f4Pv8LWSD6bGTbSbQIIAYnGuTzN//sNrSWmkOIi7EOauohVkBXxMcGyPT5
hWe1i1kY+l0epGYCXNi28lukZ6jHdRUoccOU95DjXPMA8ANsIgq9a/HZsUqaYKKD
kSoKDPenKuqz77TBw5IQLCotJsn7lc77vJqwyQC2XdT9f8SiZ+DFtfFiB36YZ62d
2XSm3bQmM4/QZD9KEKX2zOvsA2O1PEi9i+9tyqMhpJD/0+95ubDjYeh5xKAOkTTc
1DhU2IeUFKhChhT0TU5R3+1C6L0ud7X9zPN+XkNJlX6is6XZC2kpHC9pem2JUPkT
l0VUEwQ1+NvkaY3hYuEZqRS8Fc0w/YUhHu/YNLXNLPBKwkGGf5L9tnWB4HFUybFn
oFfsATWNL9nCTHTOe6Yo5kSlhG39oGCInR3tWmO7aGX/RjUe3vSN0V+NpgxSKLqL
6K0cKgVLv8T94W93BBFP45WIAMW9zvIGSe1bHIIjqdrlIejFgMjtsFp4vO4zcDQy
gVndqVoMszBlbL40e4ETc9GaySZS1kLc0nwn92RM6XnQVveMBlYxDUStAPvhPS4T
LP7yD6TYhLNyzju436XPHQq0iskk0uCT6h48H1urI44cgu6XUWBoSwSMnP5NHmUm
VfOX/TmTedUifBOPR+Ow2Bsc1/1673bAgBSe7MrE7t5tMh1oHqJKRylSBEslDPci
AF1UqiUs8QvRS+gjbZqQ+Wgq7v3TsDnjbSHfKWDqdfoduLa5e5Ogs3w3RkubCe7R
CjldE3/ZS36I9UTwZug+RHsQ0lRzzjhG9+4MwNsbffy4TYxeEidUtRdl0qvUZ7EM
uVbbY5AWKeZLaUu3LZ22bkhyBzdmIoXej76YNGQHIrqR75bvG1FNovOxlP3PiOUP
PF1svFaF711ZsyqcKbEOnxPDZXNFprQgThhsYzo9UzjrFFmrvdi2xqd+WEONNMOH
rrNpbwMedcEdNrxULo3Zs0iJocWSjGXPWbVp7fCLrQgcZw51kegu9n6EYC6Oj6tp
DvCrGDuKZFJAdNNgPdxhJJKBL/1bRCFwuU+6yZe0zRgC7f6MONYeWzI0zrw/g9RB
lI0xzVw3eLOdjEcKUaw55Mk8H1tDEby3vhaVQ3ea6EUe5zxo738q4pXFStk/j6Mf
zLg5RP83DuPtlo6GpOZTZgXO47KwDHWWYp7kGYYmfZV1pLdFgKXTwY3KCSzDrKkO
0HTsrVkGXTq1gEN8gM1LwJ1uPao1dSRx2AXKbG+C1wxLBTHwOG1UM+8NUHPMnhSe
wSqok/12lOIs1Zdc2jjILCOAN3+OZeoepQkrXnPF2DxqB59Bkwf23yvNEAJcPh//
9CaP9gocXiOfSdSK8vImCZ9alqjdN1sYuUqwCnPmSwxZ99EoWUkdnUxKixjX3BqQ
8HMmiBdVBIdnz33kGoHLS49vsUZpCLoSb9liKDkr8/EOXeLFF4pUr3mbnoG8j1XJ
wtrqxdc+CNrDyJHQS9QRyKMMOabkKMKE04WcsX6lo7HFhTf8mCaVOJYBvYWst7vd
e0MABrCz5PFznV3UCzFWXzh6r7jrSdyom2P9q4k4cxmdcQaMU6TIu7+Y789YkUIV
vq90vD8M2nw0A1YUokStOdLqnvxACB/xRXi2yTNHGm6Ucp2nQROiSQA5ryCFEXYc
f6ekQZ6uFc0sX4SmE2hXCIMYCcJTbpk+/wIw6hM6VTtqX45+zG3TxsxePMOOTTRm
aRyOxLP6BifreTGic1gMN4qzzAnzsd4NCsg5NNhmxf5AAZIlLm6NC2m4UWW39AUk
h8ReJpRaAtAPPDHb8+ZIPH+vuT5+Nh9pbVt56M3r3k6yOvY3fkXQj9JFvSTCK+pw
wBrUQG+8uYKkMbDyGYEe8WaHNoSphfH0x8L7eLtDKpFQr4e+8/gZgqBVxPKnuT9n
REWZqYGLmugXgIe6c8XqagLsxo2TOq61owdbnFLwxqxDpYYl5Lol4+p9JF3I4Pap
FhcmdI+WXyZ2aseOm1ivDbvzVkjNY2BZU9T3CKhhjfu33Jn9WjnCXxfYIZJgnzzk
Vt1o3jspnozyL6OyHrMZKL0aBK48Ek71Z879m0e/sNeqYJtYaJvrhAK9kr478HnN
29r/7FbSj13LnhPbxuMTD1wYkyeiZdGTmr4zyqIT5FFahiX9jXScwPbVqItnL479
ViWvN89Fshy4WqHSYKEa7VysZDoWPGTKVw0YQooXV2g12D39NA/1SE8dnyHqsPpt
mnz3vnX8k+jtmnEEF/Jdv3lX+D17GJjQGCgsKK7ayIilgYOCI4+HK5/ilEFaQWB9
36Dj1ESoPS9xOFec9Z75nFSEkXZYOCwZLoDYabA3dZJm87U5nD91EfsGw7CneLSF
7gAcrLcH3TG6PV80NVRK01w9wrmM5/bcNw97oeYhDoKK4ucsF2IBBc5xgxq8C+8Z
LU27Wr04FzlTd/RNOLMDtIsvV3igBp4i178pI4JXiTTrKAzCi+omlOse+s86WpH0
sOnWoNFlyhvg4UG/J6akrl4hy5sVrPO+Ei8qqbtOE0CKyEwtrvIvjP9vGGPWEzP+
87LAjAiWufFyJn09uff+Lp9D+ZrUCW+zh65kFeZCUFDVITjukacqxGA6Rd8lSTI+
jwYsj4ETpcUqZxQ28k9CYnaQCW4de5+RhS0sFOdDZBRmdyEClXkntlSYEGfHKfo1
cPmr8cyvwc2r+EAiN5oGB7LuzMh9M+ppnuwdDlwrJq+MDVSNoXkGqSLIwWRkImhO
rz/QfJaJJnp3IuyDCoY+keqG/mjTzkzdmGqGXwU00o/oL4bSIRzqgu2Jw66Ix3/V
XvJH14U1AeJ4pA/nLjO/+wCB1M6I08vbrCzoOTrYDk0+jCaQsoC7Bv/olIotlk7s
Og5q6iNqzjBJdv8NfPpSeTwTBfEuET6crq9Xhlpmu6W0iE2Bcg1+B+4/nHkYdwaB
BTj0ISNaEONlc1Hf2uf7qMZOfsPEtmqn7qatxk1HQegoIrNu22eZMDiNL6vUgixr
E25ylpBMHld2nzPMtmHH83PeGeVdH0aSAnmFX8KvgESinBHDMN73emZ41yUDjzPN
gJp//FtPjZ2ShA5Eec/yYwT0VoP14BjJOHIrUzmIF9/cctuVE2EgvoYrj4gBrWjj
A5kym3oi74V2paZ4M/XCI6h03r4QrPGWg8BYlBGqlT+1rpSgOT3zyKP4gv4nkX5O
Vso7lVlEgAEL/aztsSgoe7wlBRRn1FZJ4ve/uP2aV4X71Ash5ov9LPgxmGQm4sgu
BYr+VXYKmgbGA0JRkt/n4467lVH+Ot/PwiZJhxx00FxJWNcEKNYFcsenliuoz+U6
ugzgx3fxDPaselJeVJJdGZns4H1uxM5QGNDlTkPX1cgaxbMmn0FaNBMgnKwVqjXd
MCfwhQsut6IvidCW64LASBLpJ+iOlFoWeudwSUI6Tm0xdHGw/Wa0sfF6odFUGCu2
T4thCgH5UwhpXEfKca2IDKhKWPkP+2MhZQuC6nbeK3s9Zqy7AGpiIpZ3/HLKoQfa
8ZP7KkgJQecPKWG8aUinVrqxnoTMsihrBfXiT/BpF1a/Eju8q3QGsJPX2s9nd0FJ
lXLP41MMDRDcKGz7Tb38pggvgezbtoXA2yLcqyQ+ENbVQ1thqXoPwcGckyRLpY3r
+KYKg8hhdfKjGgnlO29NzwOpSqH/mxFuwWN8nj9Onab1fW0PmaCW6T+dLALKp4IK
gRNgMcOIolgRpadW4e2U9eQmithYroAtEdQTuxOeghNB7pU28ZoO3kvlHr2JBMF5
icYHhLMj8EWmIai1RV/u0m2sQkLRs2MyMSp9eoq9LnikoKDUIUYPg27rbfDO3D4K
gLlfiwR69t6Ng03V4Ifg60n7N63MEjnIE9vctq6B0CoZlHw5WpnAp0ITmNNGRN1L
5upNmmOHLK2IS7lr5XO3RBLMI9elo1RHj3rViIw1qZNLhg0167d7g+UvUznX8Pxd
HjgknlLB1PAAaINS/OlSYdD3lgzfhPCKvPZXNdT+GPx+5+JLwEKA3i9zLcbtK/FC
WgwbrFK8bEW4N5TQ6NBiyZ9VIVPmfBlHUjmG8qP7CxPGrJ5oeikXwA3zlYYQP0I1
OfzCGAB/RclsqEfNWepgcEf3Rz+Y0iO1j7qboTfl2214A0J76jmU5yuVSl7u2FVX
m92fviki5CKv/6wvpDeOXWfabYYoIWrOiuOlpwxR9Qs8EbNP2u71HAC40f2a+ZEL
79bFRuA78a0aqrhPaEmve6PLvUQGHSKn9gXc4MX9v0bTnNnKkC8ywyZm7LPeE100
eP5Q2wzlXGst0eD6BrqJsfidyISC4c67EmqddZ6Qz0vdMgjgD6ziJVQ6P/N9Z0eC
Gum+OLOHyIP/KoV8LA+iCRQqOS2SJALkgyvzI8jzCN9jPTyNdTMJ2sAoBW3ak9jU
UJkowzs8zuHtCk7wEN7V5DqW1dwZQ0Qln+BQi/j6h2TIN1eE4ULSElDz9OJF+2qd
hOC9yvlgGoaEzkvvE2oRqJtrdghWS0f4tHzahtLJYFxyT22mnKXCUFTHLEPIYy1N
WgUIqcNkLDKhtRu9lcqPYuNUJTq8MenZJtMI546/dvttHo6oB+h2x3Knh2J+24gg
WKInZqU0QmlSUEjDwjX9RceUEv3/NAEns6BE3gbKMH5knZGg9ovKfthoDQ/+D/XA
uEFQ/gs8X5cYyUwvCz6oIRz6TMr5Lh3+yx483MtanZcl9ymZBJ5y3s54LGk4fa9L
hmxn79/QllKbozq9bQsdBD/4kDeRNBHYRBg9pnx2EVDYlGH7+sJ0/j1j+6VczkPc
EU6QhmuQZpeHNrlxfWjft+deJwOemjfvB58NsSOHBdXzulvLhP+3P+RnIc9/5V+i
k/sjXoZ86fpdnxjvkTrcD8dxpxFp1lkE55/omexOTxXGjt/CG+RWOxSsEbs5CZ4N
TLwdmeGrh8rKiBAWwiuymMySBw8lP5zD2kY5E086VM/ZbyccbfYwDPZJx8B8B1t/
yk4qFQtB3bX+vxL1DyfUtWBXUA87ldO+JMkWldFW1jrl8LInPJt2gzX+5yDppk1t
3z9rzD5Bqv6Pb/US4cQgqKTpwYU5XXVXoacHowEeybRMQz/yG6z78z69aamm4U73
w0bbZcr1yzCPh6MttN83+Wlof7u2ar4eVpXTjE/H0O0qMasYFe036k1zTxwg412j
ZIqysVn+9H42dZzpBpe1zypqyW5luUQASc6o5ZL+ce8SC76QWKJAljSgkXSSFdN8
0bHNp5tfVjXO5YIh9MzJraJsZJLowQXKclX99IR7i4c7TvZMM501bpYB67cY/g3S
vJyVFltTeeEdjWeaJawBTHfudgdDdke0Ihyls4eLXEpId5+TFShYomEx5TZrvYRW
lgql825/fNZ/NA4aEQKU2WHTBsxqRqCCnAuG8hBJelb9Ynsux+ExPeY45lHPkAjH
kCrcyNp78HOVVZihLIf0OfSmvG6W/P9fw6Vay4/E/3A7YGhQFyMjigZ7Am7YZKQu
NFWm+ZMemeKpmrSstHtYxfCYiMuv/Ge7MkrQwDsRacnCNN/iP802DqQ82sxDOWsH
CwTnV2fi9NJyFU++Bl9CJ0gMaIkmuGbYUewPf3rYhi5OxKoJFlbAJo4xT61Cw6Mp
EvZwRGTzWj4w8Fx1D9aqPAa7sdV6bAtCo878yVHjNhnGtxT98vpskRJwMAnlQ7LL
c0cfCSGpXwjV/79672WhRkZtQJy6WeV7iM9wKKIydAZUYUQVKrQmptTsL+tjxUWC
DJyNPBkkoB3Vx7ugukrW0LC/zj5Ift8iSt2ggUR3lIyEe4SuXysDoWdeCvZEmuPU
+baPrztO0ZLY7vh4sCRxbNqw5peLGIgsEF5DRHUfOWQVB/ZcfK8OaXoZAjc3MEHa
w1hZ0we3A+7UHViNbUx0Gt3j8MdHogBVTPhflny+LFF7ZGw5fFMGldLR4ZByntYl
RqMVBtAOm3AYu84YuR9AKgssaZ0pplgDZqHesnWEts7yyRfz2RVhbHl31Fmd+yFL
I8c0yXBukBP/vhjKOdHHbxKOCGcQ4/QQmAclkYjXmEQbcRfwDsiWuxGXr/Tb2sJ4
uHz/m5am16e597gYU5WGYA/wpvFt5UmLwfgCPgOpxuAUDbMF1TnOQG75PDIJ261H
3UVMhicmN7er4u8yjjp96mxzcGSnx3xVhiCfBccqnH1C7Jk9PiZc+gGF1SCI2ghc
rRNPZL9OL1o+tuJNaEnKr3cQ7gBIAZWMqv0CrkA0s9Lm/pZKAiggdiAl+srLnsUb
7UKDJxc5za64cj5tgoJXdaJ0ASJf1cIC2gbhRIoNeuz/MnID9mXhIBGyFbvFTvu3
/uwnXfUlvQgF3THJllwiDFXvgTcUGiMmTAAvckgbhW14yfdTmKy99mu7d2uyVNME
DA/3lanX5stNtr3Pw8yIHHoNLP+BPBsuBRZt6n7oX2bsq89Xt8vXl1Z9DsBeaQFo
i6Nb6OtBRrGavNvlfGJrNdvbpKDHE4lACDGBXrZC3+fuFWsiet0oATpWMZVEUuYL
EsQ3I3WpTBB+jGIbhnZ6xhGHHYCxFo4EGvbWNO/KPfkpme2t2DRTH3pEBaKUIVV/
gDm0ThWvarQCJ0D46jL6m2v+D6/P/bBZPapUoOD8LjYD2tsRYvONmFM8XdwZZS6g
mmSSpikozvmRwPXJqonj9NjIeTRwggE5ZF7T+9qSqDQqGyOEJM/9ILs6Lzp6Bc4n
tmW7T/Dkft44mWg5bRuRC7FsoBQtviA2dOo/pM4YShAP+wYO0aoQY4+0V4UFvmh5
+7KERJCose+1bWZp2zq5gjUbjalQi7HfpXHaVwZJNENt20VEZyPPp3z40004gPjQ
jYkl4MUIZn77e+wOHM78LSbxA5MkqTBjHBf/JiU93MNp6+6ddDgeJp7WGsik3nQ+
M5IH4DVf3sS2omvGg3o0nZv5PxhPnK2PyHj18ViU329x+ttV16WRzBWYBOhQjm8i
gOHHyCCm+KeEQci+0IfpUJCiny7/G0W0n1FCzCWym9vpVJ94MK0Rjutjmyqgagra
PpnSZH4NRTl7c6/pzeGMH+xYMsfhO8PmOF0uBN279DLzjprfQ5qCDPwzlcGoBAYg
yum2MY0nNoKjbE+rchjqgj7BwjmQVMocsrg51JEmQoV4v7QO58d3u6To1fPWCvHV
cImbgW77JBwISvKiqN3uAbkC0HVsB35oyf/OJMicq1OstJvAddRfX8OXNEKXMS/j
k0CAutNObFJYkD+qcKZr200ngd1zafpQ4EzsWmROb/p3fdWVhHdPqVJRnXGVMh7E
EE5cbs2i7KXaof/dX4B0C1vHM6punUjBFrtN5vin9zdwN+bDJEHhD584uEkbVNUF
PhfxeZBjNDL/qv/R9zVSVBMJx7K0nS4vh7+CzG/eMlY0Kvam6hzOyfWbqBMBgG27
jWDTnm3jwzUqG7HIoXaBzgi2zlAyZIIYGZF2X4gLAGBC3mPk3Dv7GXle9twju21l
L4+o6TNoGellGL8Jpuxq9gQIlctXo4wmjHC65iIGs5Hhijw0zOtELU61TbIrOq2o
xOWnwxpNudynXp2JwIJzWMPToP/34aUWn+7IisyoDE2h39r6PtJVwg3F3u0S93HG
8mz6tRKrlh2qkZcPXBXwYV2hf9FNMFsQo2EEH/s1A3ZymiP7hQMFG7tdxy1X6HAO
2LKzbm+SIiKo44Xt5mBd/ty6AXw6wvw4FqsTAwZjKXUpfuzIGTmiYmUKV9ZH62Vd
qMqCgGz9tyACK6IveNrK7GXv4GsMzH+MxqO2guOPRuznM71jEfh1jkTwOGC1yhFc
Ah5eZbWWFp2WEjLBLA4/wRVrw1nv3X3iMnDjiJuGWyNKygj00vKNY/MIQdDcF+8R
pLV/EK6fLL01DSrX7lB0OQCRX9oD6axECkCSfIoSgynPyogVuCv5VtNfrtwZyYV6
Qn9a/55EmChMlFWfZmm04ESilHr5tJTvL8pNu2KDIT9jk1ZLfWa/ZpzNxgSaPr7S
Ew1qaximrlOzPFoCUAvUnVSyAzx1bh8aNlnwPbi8IJY/Lsix01Hb9jsZGApEGsmG
WuxAoVbOWKejPGflZ7RvM2KKFki38OrPSXtV42wBnBgqg0EVXzRsBbi0ywhhlt5e
VJAhqkFpB03HyKqutP7Y5sMW30YZRCQYwz8oED+ooZoLJIoyTgjv9hrS3IaUvMcd
tOH8AF3BKkYDNBUWvhKcqLDt3Bom+6Fga068ROAp2qzGTS8z0+0nNZSuKtwtarWs
TWQoDY/BKpw2kS8MGZuvVxGdjCUFvHjJszEanow6W+Axte+NTyqJklPx7m3W8U/+
NAuoB9hkv5tIGvcDC/OXGODWRVcvYvLUu6hd/DIApmZ+PDjGQwOjpnLxKKguYoXx
baH909vhlEiy/wxdf9+2cvrAIPhnoE1ZhiznS96kJGVWVC3A287SxAAME2gyN8xh
ZjhpUednHE2Mx5M1HgHP+lJuJPqZu6GLLTRrp8mtTb3EEKnZxMZAlrhq4473wn7J
6RyH5EBDuABBb5QUJEeWltFiAhNN7eV5nMwipvO5EpBJlh9prtZr67IHit8c7HLF
rYK71w4uFhcD4MRCHkS2sgz2xWnVaYdczFwuzOY4uq2xSrpmufZTEK9Vta+zxC/I
kZx81MNMJFwLqJwVbKwwpzeU/4ddJfcf+F5pTgxkJwZel5Khr4gUcASMAdNLClXR
uq1NnwjIDoxILVCdJXisKzA1gv8fq86lKvwrf78t3gnoK2kr5Ctb2+qW6iEOzEx8
4q4Q+GNLISYG5lWWIXtD3KgIb5x2HE53c0T1faTSaLIO9KcWOqUkz9CDV9k7rdcu
ZkxZyHj5URan9NXP5RxvNCbk7EaiItBY7Cy7B1VmiLfrcC7mkjIyZVorgcZrTs0+
YCc1GmEFf7c1caVfMwXzr+D1tbL+J8eVQOQ+VBcYXhcw+zlL2NgK4LfwgmjscK+n
s7bXFjrk5A9/5tDXyQOjNNyYE9Siarfh7lYelvtFj9ZyAVR2kWGAOUSW6sGIPg6W
eYq3/V1PYFAvVM/Td5kBazDsC7nGWvUw1RioVngM1Jb/CHEDg3fRSVqRIo774ZcP
/5sYe7xoXr7Lcwdu/ue2IQIoBrJdpGz8FA9kg+ZjJ1cxXzwDgAUQFkb2RVMgIuXi
DbXDccbv1Xc9gPiEw8fl6sAAP3sOra8LO7TnygT5v1IHNLtS1RqlbI+fJ1nfhihU
szDA/XOzjleWXJkpvJSVO85OiqQKzVySGwGD85eNcubtykc96LvcFnYN0p0mM8YC
oMHtqm6ShV7AyUbSwQiakD54Y4PzRuRqlj2F6ZAPEmbDyJJjzJeYLmGJ1LogkeAP
vhHd6ZDjGJtU0VTEfJ8jtcqQt07eZENFLMNZ90V2xDPqX2lirVF4ZGg5S9isdxT6
kqfp76HDPopVBLf2wVGIp3vBPjM/M0KQRjszXOqY+ERzCEzRKZo/Y146wpjLiyfH
22M8IwJdcJc/XfV1SvxSBxryK9sE9NtycpIQueQ1Ak1jDFFj+OFajAf4nHNGbqtP
H3Rckym3MvOlZUozSH8Gqe5AVVgSW/lhp5QYmwMX17L8IhvCtelggy1rSCBjEkWI
532j6kAtYzMaZkV+w7bB0Rthd7psjx6JvjZUmDCa/WAyAK+WoxcaN+XzLq/Ji4jQ
wToos1ylTtOsy3hn+4bh/QsWDXpo4azLgWgn7M8vx5mcXU0HWQaZxHN9P5oBZDX7
hE6+AOPt1ZhsS0uHK2AtXf/KnxP/MlhsBDn4N8oKU1e374qWKuGMFfDilB3jmGR1
rAPERtxqemOQf7WjCyKUEXvF61ZSzK7dclVnWkiqWaRONqqHsHFEcL4Whoan7IT5
ys8Hyu1ZLJS2NzFLM9Qp5bIZob/bV+m8C6pPdbYc09ZJL4bPYkEZTUGhSH5Ba+hT
XlegaZsbu68m4eD7OjkQjRhJx+IhTj9bfl2Q4Xx6I1Wyju3ly3uuzOnCchYvCanP
c+aTPhfgA6Q5O/Onlgkz3f9cGjB11dND8Is24Q7eHp5l15CLIz/w7xWN6L/AY3ut
6lS2hrouzebyVEbvR20HcliuAj6A+CNS5gXdGPw0jGkois2WDnoARAw7T7+UBH7I
/cDyoi6kd2N1qI9MiS//Pw7ImPN5iSKWaXNz4XeVsPQNoLUxgAkNNe0iuTcIvWSE
DL8Z4EPPKdgd453ToXvRq2KoTVF2+cDuKBXBt/tMwqXlDfOrTD79gvHjP0ZuaRG2
QFH/KYyJ7ImSdKF7Sd8/qpKSBiqZfiB8fqGZ0vb3rY5Zjgrbt15Nv6Bph7wN/5gl
ehy+Zrs3vS0yd+m07OYZ41+FMnLjBnGCpXHXbe9eIKox21/D9qKyI2BIkcBstv+3
Ya6acNvHdacRme7S7vyJ1sPfMidf97eVjOQwB3gP2ppB/18qfCTNi4TY44D5xsVD
OFezM2Uek1EENi6mxufF1LFAGzgGCVsqU4ozWEiKlEanUIxZIMkzSCHRoXjYc+SG
pO4T6LpLEuBBj4TDCB9XPdcUlNO7Lt9JDASAKq6RtAlklZzBPEaW9po3fY6IRPZT
eTPcs1EQxfnh788/zdAkWDM8MtFsPINTQlxQQbnlkSmS0P8jqJg5QRqNlPev4oQF
hwZoUL8iqooNW4dAFfR27mMyWPP2D2kgdfB3Lf1KGg8nnLp3lQPjDaZTHi4MWhgQ
Q0pR/zE48wr0jXiMQTJUonUT0hvmjaO8UY3xerr8oOIQ6VQmwdbADlIKbsstR2oc
Uu0JgsD3ox8HmYPLgnz1IWRWfw7LzTb06/+yS4z3xB2OCtGgjKJHXROJhDslmB0o
h1BKJqf6RVfT7yZt7V5w5081KtKWPfpp8mGZGJN9P46KciuTVDCYC3HBa8YH87yJ
7EZ14mBcH1C+TGEF4hpi7dcolzMO5HuxAT4DQygKz9XrIlpXTUDO7Gej7bCS54lV
RVtG5+v4yaPLml6702AurCCEq7GERmtQBJSdn5AvXZ7xYou1TRAznyQvaKCr+6hl
GQvhK/v2V+qj0lmfDHf528WHDA17/njGFCNiS2CgMFZln1/FxLgqKd4gZxjh7449
R/BtNrxmYfZmwM9Zg7Qc6rddUIKMN1gPyxoJOijYxsvCXFZwzC+7lj0iU2Kizxok
RjUMSJJ2IIRGiued7mgxcLmeFOJ0Ac2aoeJB8aXEQpAPnoHJDkGoYr9J9GA4rs1U
6XzMTRZykVNmuBG0Nhs3vpFv6KycFJ0Iy/LTbN60SFBNUDcyM8yBhY7lJjU8JVq2
nywqShN2qp5u4DepTiIj5TLyQks6jnClUrEkm7RnvduSzF6KBtxa8QWdMke1LaWB
ctjLpCgz/pzUWR4DLtrSLKqrGN+dT/vbyePqbHQS7ung3nr1hl+hUM9J3wuB+r8w
3vI54lI3+noEcjtTb1f+fuX+5lamaN0719Wz4pgpaRVxUr8g8eKrczOVe2hO6BFr
Ic7rhbSAC9B4UKiDPDEiN2uAWpLQpb6pLqUWWoIf+l7ofRHejwD1LfRprZgAqqZk
85XTFzvtNO9H4j6tbDdqE21tmYeSdE49jq1+2RFnl/BYTZWhBqQxH/wEu1vL+P8+
/iDEXEFZj0ZTa8V5TnvWoRxmsnK2wDWQuiUvhAjs9QZBBtPv8PyeMfMNMgsmAnqA
C674XEYTyhprBo76GYZycFMpfKZCcfzyJC163o0icCafvhmwJZOOIFXBaRc6QL69
rkmtD5gBSNbCPAkzKA10ZLnxa3m5wa7GFIlCDIAmL92y9XgwjlHtoLix09ORNZUU
I8kIcbanqzz9OPO7a+KGeDuZfaVqg5T6UNRVkVEaH6Xcr42DXXTgLwXN7PsluE/m
iK8y8GpH1sH8pPbNaxSlx8Ud3TfcxWYWDkOB+jUSo96ljtlsIl8pXrZ1ikQ7mAfM
z4ORqbRgi28cXJMN/K9F3LME/ALzXQvuRQd5OX5fd4YvVDbNGXNiijGVihiEgjnR
fzbDXJVS4oWfwB2omEtwKi/QrheBRQhqAkzE7tOvLZvt5upNAjRkJlU88X6tlbY1
emb+VCNssQB2pEdCJ+BrTxBB2754PdHbgclA1R8pn8b4crXSn6smk/PWy7GZu0sz
G5snBnVlJu9tNk+NjiZrf9uy7ZVoQTINjrz9RfnTi/a5XdQoJcBKtNpggXARDD48
TQU0UEETE7D39f6kWb0vlaYxh/54N+5VBFl7SUZspQ6xHd3qlBieRVXGPj4E8siB
V4zCorPNwSGAtlkJeP7S9rtlYX/RGRja8XFsT7TZzzFUZQmRUwcFSQecX6lQ3jk5
i0BSd13fZBTH+c8Y78/MfzRXNFJXAlALFLAc4jfxhnBnQx6i1f1x3qV+eBjjqya0
4QYnnU3xY0OIFWpQgmqCiwfF/v8+20cIyrypZC17pvUadW0LSrw3gszbEjvlIvhH
mojpUPCDM24Qs0mXJik7/Xh+sEAmJkvQP6mx6G8pBbKvxVq3hV6hlMesJ0jg/6Lm
dJkQ2OLEqQhyuB9Zm6PD0Xoyqk+qNwr/vRvig+4uHvCBPwrVbwaXoJFYrxZVQY5j
T3ZtBqHmoFhBPcZb+B0RrHxnWyK9PQFzjH6jjaG/oE0Hr/Dn5EtUpwO7o2teOmIs
VKRkmXXAtNtYCiG4dx3ePswrLWHgHy9xOP8/3ly+oGop9vM/4dCmYCNLVnqUw1J5
q1HFc6ppvfvXRJD5OQ3+4CuvErXvsFbMrt0+IblXBYqY8lU1B9ihb6DLORHLVoSO
SKGkVT6/20R1sZDzEubi8VkiAD+CRs+SfGa6evc0weWzkQm5/ldbmGObhJZxKinm
43JqpjW9BaUa7v/qbzrQyaRHs8lCVoRFeOrY6BnsVvtY0AC2LAYnqIiIM7+JZRTL
xsly7xUXj85eyll8REUGSX0+DDAJrsTBpDQiE4Caakxoq3reoEyUAA1NvX6s4cg2
hOvPQn7vsxZWsjp5NcG35dSUwcyX5tGspd9RXbx1zOGsiGAm18hid6FJoz3UYGf+
VPruTYZ14ju4pcms2Ru+LWoJcpG/InxEWMN8XC6jNeMLzlgkQ8noWjtLeBQxSFhw
wMkPZmJfrV5BfOL5LJsn1k22WcJFdwlLEKIBldWjNQ4eeoHtEyGjbGmgvqYiUPa9
bPx+PQ5qkO12mYb/JJhaU/QFk1duhKKfL1cFWOuGOc0d8IioxnRuCp9XnFFcKZuh
+Ng4l3WRujyrIKiVZSutleMB0oUCkIWhMxB3Ro7PjRCua5ZSET8dm+6lCWnXgzwe
tSMlfdvw8BoqpTlzi9xIOEgXQuItTH++yRVIoo5juz8PlTQXbLjB1etu24FXVgBo
x8oN67taUPJGxhJhUK+e/GJzWPYSQR7aXhz71yn21Wf1N4IFto6DCxyDtWsggLYM
9V41MG4kn7fI3FAalkrfBBsIq1uhxhq585Wiqz/QzqXwzVHbfE82plq8pYxM0H12
kZ/triFOj6L5str1WvtBF2poHkbmb13dRiv4/vslbZYIK/NlrXNM9Tk8UYckGutQ
NNa3O6YZivRyEcD+zPCxN7elKveC5wdsmEX3wXnbLdLlowvtiszwGx2qefOroztm
/xI8Klh0xcdxgC9X3PhOu2ZYeNuf38IYex2MBYyhckEaIxCBnHzyBVN8HvDx26s+
sUyBWRdsCm/56HiSEf9+MAE2j5N2ynGh4M8n7IRICAPQSD8QsCwZbu+yfjZTNX6w
Ek7GPe7lI8+NTbaH4wy0/ApX/5nUsDLe6EB5kzNCbXI1cUGzhp+E1wVcET6zghYo
zFBvUdd93kH/2NMNI47O30v78BSdt8MsKNWf4Jf4yHK07Pl+n2eg9p58V2f3LAnX
7QIVrdR+U01MfY+gEbNydgXP+3AF2UpZprkfA1fFOykdjBTjY0JqEbrXH+9vVq54
8zcZ7glfwbcdL6QKC3HTogRleA3Yf5G9nbtzh4Qp/DN8MUveoJgqvPoW3IHev/la
OohW+CX60llFuKL7axEUvlrIQQKl2BGu/XFE9Oyfo2QHSFvksvwybi6V3langxlr
1nbiE7mThEpovJNiT3FJmS6LJ3u/CDXPfYXePaYPHkTwvXIL/BjoAhpH6Be2U6hP
cC5ZQD0Abs+l8QKbRjegaMs+mhZDHwu3Kbb3JS4xJ6j0F6GCwvchtcPZZYU3v3l5
zIPMfZFmDUS2/7h0IR/d3aS/W6SYyB6IlcE810LIHmCBiVM28cW+csC200b7bXKk
sbWVRdD2dJ/tsXFtkwcJaDLn22y/agnuraI3IaeU5QDoaH7Ieuqh3uWxPd0QircW
OKzFFor9Ia0+TZi2t2//NYaunCMLJy+sp+a8yvGQ8VmCUqVdaft2AxGKI+45EwMC
AsCH8u+zxFop5TX1KjKEYF8cxV3ucKUAvu8fV5uSwi6TKJaK6IbRM49vA1oBcSrc
J7HDSEYDPHFA4Qox+NF5VEQNWhJFtxEzxp9fZsoKB8wI4os6Z1BQe8VKdTvcJS6X
wrfXeyZNxAj5WWVgyhMg5UTGc0TE+vd7DJxSttITyKDwEgZrjogNfxfVPite481Z
l6FJzacBCt8WWGZ8+c0ZL3yIlxB1Xgha0B1CsxriJmQESNgkFu53vmoY/KKI3SRu
aYNFJTkPl+y4S545ZOR5zuRn0DnlsVDeixHidJT46ESMNUa6BRovXOt5KK5BZOle
pl3bzWu3m7RedboY+E7SPvsUb83VazODLa7KvJiWW7XlLQ1sC7X/oqO9Zbwdk4N3
ILS585uRN70hshuqCvBLKCr0aUOxIeGTLvIg9Tdcd1o/ZQlyHyl9aUwNdOzQelGi
jv3LefiEjkx7/Xh7gSSVlN9WSqf8jNCpCaPd6McyIPvKsU4SvqNcUta1MLXXtTDu
VoW3vC+1yhUhclRTLF56mA3NnCd8A4/xFFhRThsu8PUrFB1oKnICNEcmk2tYo4Ti
S9JrDte/feMEpiUC+0XCsw3UDGbaB+LFL6QCtodAjy8zfnz3tfThyi5hzPJMfml4
vhCqU90NaRq6V6gr/Saegs4azNnKIIz7k6McC6d548OjAEOG/4eXSgYsGgwfvGHZ
fappwuGarZpAhkEq/kDYyniGeeipkNYAREgHdfA97TiL9Sg8Gh9l7q0QSqRVfFTj
06JOyJLZNFG8y5xNNyHrzRt2MOu8xUblBW3W0ucmZEcbM5eX4XVHx9YkGuhfsVBy
cwSIERLP6w9k8Oi02+et2mxkFPzGjcU3q7G+Cru0eqi9uYzE/JX1IRGBut2Qn5Fa
C56qUne05HKZ/bM1uKrMbzFX7/MqNyJK4ET2pqg/oLtD9GcfFY45/AjgukVv+hM5
weDqKd3fl6Tt3nxoND75uz32fNAK49k4xQIOs2OAxQcBAmB5AuaXfd4bPU87fxIN
ns4wS8gT6z4SxFnjk5FKwK21Bb4+6CQDUclWMzrKMxwnCz5pOMw80XaRfsbS4ble
s/c1pt19pBZyyY1OGWu4gCi0AMo+WLE5IloGdE5WLhLK3ZE8tt0vYnB3+1E06Qcw
8UuEDT+oPyHlWOhrnqPxg845rDR6iGgV+Mm4kf5hXKk1oBN2PUNbRuazl9di1wh7
8eVvGhhdRV3WdXo9ovnHdK7oWxwVbMtpGV5V4CmPjXc4fjadXTBVznaHf/0/notT
0Yqoka9kiGHCO+qISiSn4LKvvycTqNG4KSs1xABeNOZu4+vkd7iYjiYb/pwj0xo8
VFJPPlW1mIH4Va1ETgHV+lsTwAhxyML2F4xTI7RmfIi02gWILeJohITvuCmBewZQ
8tx9tePlsAUv9o8USnQ43Dn9IIQAXghYnGIfRKSsgL7Eg4tSgSlk75S7qTezok3S
g6OaBPsybqwzTJUVEZA+B8McbPI7+qJWcKIFs8ai72Uq2iZPV7+Wc/fte058i15r
sckeyqR+S6Lv0dDMTO+mqGmyTrONI4j5RdkrkJSZr8PV/MHDWQ8g6qlt/3V6y1qq
Q8B50ZgoyK3qOOiwnOVA0H4aYyKwfpJKuMHlu2IiCyLnAwfByLW3eihpVpPlrDIg
mUhyhcbu36i1wdWr4rszM3jRnUdJgobzP5ddcC1Wy2aJsLdAf209McZYMGjXhFng
tO3DnEMEQNsCgIdNfisLwNjxq9VlVyjJDG6KqXq4h0b9huCMV38i6f2GegboQmru
Yu3fiZB+H65ENk+wZLB//FG9BICC2GNY2cvgfKd29pt/yotgLzGB/OGHlQZ+sqbK
Olrg/PdK1e0nl0v6Z6ezwUgP9Zib6RJqYr+Q/YlvmsV02/8U3qlngLn6cNleVEK6
l9SGOPBOGp7VV2BHZIDXD/4PZrqAoGpaMPfebH+YxqxmI33GYWP42J22ZxtFOfvO
+Cx7D5QZmCIT4iZxRxERVosXtO2w1R8MINy5LsmcciTMomSk0OS4F7fXwo5oLgV7
2N3ajgSAlbCpb2nVtBbxWOMFtHab3SErFTB8QofbPSLu7DodtYPa4GmF2ncZYW1z
ahJgwQo3QEx94TEMwB9rB1zV94IfUY2nSwObc2LwIsjwEsWtg0rKzFWToDOd9zJW
aMuE/GR66f8FyBS5xC+wtJom6ltAam2qAJWlOR0v0VjtAPhlRiQ2bK57Lykd7xK2
Df3jJ9/lPOXsje6Xo3AXWzJCR5mV8vqfTLKVLtlHETriE3xjfAdXXCXa4DxO/qG6
SE9Oii/tqWsmblX4+ap6ZOLnUxHkXsLapB2PaPudwko5u5PDVoexhQ44UFGH/jOy
H+9UpFvu6tT0+XnLas4z0cXZZZhGqX/pKQZGPdz++SM2ZZNelqZQnJx2AcjBXm8n
6d4oXkvwik7yp9Dl3LKYUL126WWjN1TXe2AXPag4VcKelQJCWz34ShKXj8Gfl404
VK8B7wvURDiOUz5PWzRDclrGSxsmNwDITRNESwJkHB+a4uozxcyaowwvTpiI2rxF
4/bLMx714gQR37d8h2cWzP3c5awanlRD0xR/1Mj4rD46xiC82mcagjDqH6BUlpRF
kuTLhw+bVaEI+aTGqFIo/JCJ9O4OsJcySy1tXKz6IvJCXk6j47Wb+1o4nK2pwvYN
HXJhXpyk/6LgRD+JjjTyuo9UsUo2N8d7S6ZKVH6uz8t6L4O+3qYNFFf8kKSFWeQf
EN4KU509hWFW5wnC4jDnQTnM+rxHRYDXfYsxMgww81oZBv0kLNrXr6pW7xbtZI2X
DfA/jPX0m2/DPikJR1q2zw1xImFTT/7Aq/QgnRn9cUr2qDpnEc6lzv6YDxfoXx17
cgu42AfgiG9Rp6Weq1srjM1DCW8rEsgRS7cYXHqDGc/hNII3ZRuHzXi3WKhstkzV
BAqP27PBF5VqB6FMk9ITekl2wkREJG5c4/ZaYVWgleZXqJDsp+YXtDZFUhrLTF7l
fPowkg0UWpE5OHijTyod6l2hVbHozvrj/R39ohoj5ejbv3HXYZ3eafOFoKk4F1GC
SF90JPxOWj5qONL458aaJ/Vs2quwsQcRng6TdKR+7EBTbQVRV3/GK1EYY562qRSv
QMMgAEag8nkeH8WF1fdF+k2rwdPaXTunAVo0nuHhB33oAW4CZJW1ancg4c/IF9Pc
X22Vb8H2LTGKCzn4DopX0MIvYiSgepPyCdGC/SwdrZQJb5VYaINlt4UFewlu/0Sz
y5igWXIXaPJ2OF9rd33uREHLt+++dt86Ngk+om0W8OZ/yNogyXpOzi90RDul3r/Y
r57SzLDgSjbVldJUL4TSsk0dl92exwodyXuaLoUOSZHHqTAjgPYnJun7pcO9VMeN
XxTqB2VXyBoE01A5GQBS61djcmArSRHnnd+ONf1O+TNMQK505615f3M5+d7ADK3T
90ECj/dGu0MM1TKDtjoqeET1BYmdnZHOdIt5NmHcdxy+9NCDbe6J9HNxqYJdqwDs
RBX3nS+RwyMuFTBQ0lgaK65MMdbZPkJ59Oxecz73g5o1dO5SDCDNctjKoSwaS7Rw
xtDfZZ0mgp2Q73IFFUupgLPVU3KcKqtjzj2a2D1f6vLS8yFJ8XEVi6ePSZIHIlkr
5YwWprpWqMnX0WZjWU4AvSOrWN65Tv0EKL/1ui6DyaVqEqJ/AAuKWbuVDhpMZnN2
YJMijvPkbDy1gk1hafticFd2NTbCEszxqgH45V0Iplj3X/c+XImnTtHV5MZ/s7Gp
wjCTJ4C0LRmVMdzSY+tN+JUNZMBjY92NCJbdtl30ffFqGKDG50UT9/nJtWrru4b2
Lk2q6KpSRTI9ey7gRvnjgoWEl/c0JWHZ1Lgab1I7xtMB4Nc3mLGoOUjhwAxtQIUp
EzZ8NVHz9ZAWgNDb4y2H1eAqq3tALA9uyexpWFRx3ixb5y/xCkqUdXKfNH5xekTQ
4iKr/lHnnE729E4CT5fChjsuZpQuh34Z1SQxvIVwI6ZlBGfczxUfrAY8ALag0PJD
g1YrChI6dZ56Wo4fQxxhSTeIVQIf5NUcUVWsNlHt6dW1KrLlNC07UphjtVV27XFP
yGQrXOsMkL7RVk8ZAWmzuWmpGDEho1iNdPBN/NKVbbC6Q18/HFREv9rfOvyoj7H5
GwxS2YJrnHZKGh9ZcU1/f3MdCXpaSv7xZ+Ws6YiVsASXew6Fh4Zl7Bw8WYroLT6C
Mlf12j+Y9V2dkwA81lS8T1Yh5QB05UsEIkWEZzPkpVyw1pGJb5QFAy84kpiyAQ3G
HJ9djv4pPz+oQR7vUIvCrlaFih8fQ1HkS9g+1p3e1BMjGvAP/IH7Kdc1HCCEjTRx
2TGqr8U3k1llwlgD+h832/UUH20K7NXijDwG8IvwI2pQp1AH9KULsJg76BXas/Mb
8XMbs9XTyR0IiSaAE6Pe8rZrO+LY6uoIB+i8y7xhYuQcnTuImCfiXsyHgmrgLsoi
fN2dhvi4SQW1IEohqkuGPB3YOE/1Fzyg5JT42ufVagqA76Fk7CG9k7takEA+VIyP
tbubCYZ3jYkXY59T2RUedn5551Q9GTxR+PzNyFdZ62a43yUWB9uyVby+pD33Udsj
sjbdDohnlzed23ppWqsJAP0v6jQunelFjqG0uY8fevs2By91GM02IJiR7iNlTiKt
Letq08ToFcjxeyNBPoBl7/IvGlM8gN2JgcqK/6wnu0gYjJZQYBhNo/yGQspustSu
w6+mL/3WJflbZQYYFYxi8vYkXG3RwY3a3DkK427DIn57df2VtAVhfc5AQAcdFS7T
wimEl/6HFRVkV2hNbDMf3qOfx5VMmEW6f2pBMzNVbCJFmLfgpEuZMgfguAJgVseN
2q/4SvsRUbE3400QbcV65juprE+Ns3DRPL+As4quRKo9+lNqpEzdsSxwuEMcgMUY
iprmttroKwrtjxWfMJHIXVAjBJG4cJ2N1bqMyl8Cfkg3mxjxDOKbFy49H39yyvya
6hmxPR2eS1QJYVsS4uvn5S9onT0zelBzsfhH084t1tY6IkDh+FO1rzTYMdTDjE9N
MOQPBdQlpgE6jyphc7gM6QdsxOg/FDDVQbvBiBFdqjwG0g5EWtBZzgJwNumBdgrf
C/MTpcUz//DnNFh3VgZZ1OvVKcvkhZoQQEF2OQdLbCK636lFprmxuJOnLdmTlu6r
ZWoHIXCXOEL4cfwChD9jY50nUUVpKZ1rjV4n45JGXfWYhNqxslejpXA8ajx+mZi/
6j6gUnmLfRUk8F5oHKferen5erT80whlvIqfjN+WkfoO3J+Ur19Gr5+6H3j7aOtx
21R4Xmm/2NZS63jw9iH/W4aoFVXOxwBAWiQJFZA6G0Dfp+Ai4VK5Ew2/kKENSNgw
y8eaKfhMy/CTC9RKlS4gCYvp3rSC4+2jv70cUoWJh6rC7LBWrkqQYJ5ZpReHrtzd
AnLZAnKYGTicuHJ2nFOu2p4lqZhwSs2m5ps2mvzW0D1WKCakWPB/xi0SN1h7KISp
Cb7RROPRxUouQtdg58ZPsu44jVvd7NwRjbfPKZLl+Ji0QoeFn6UHDjX+VOeJAW8o
Qp7MgLxp4kvPO0TZ3tJj/H7Mp14AggfMGAyo43iDDwbGUOWUyEjp8MhR5qT7WtXq
eBC3Q7wjnJUcfNmew0fxBdGFo/o6/7STJLL26AbaP4/s4N4JbKtv6NTWWc3k1+ia
vdJbr2IpnRYlnFAr1RtUdw0ZbhEfJ8qG4jcawhJyqHQiYMA1ZN9+4lmQv8Dzr19V
19B398sKkJxajhWERspLTPR61oSu0m1Ot6xDcxpcVUg+l3yHBgq2v0XqSoBIwP9g
1Gb8zIVf0vVq5HAyV7L1vtyadR6/CnPAVxd1EL4DcGXiGi4wsf4grybTTImq/8Lq
V5Gnltbi3geJ9hiGqnRpY6rNuKpp+ys5LSyeQdqOlODGSN4XbOFfi4mKRD8E2n5A
5zRpiFSNNkrmraAdB66z9VAIV4loHjjc/ujN7HFwakcMzo1CAY2BfeyLKsOmI84K
ZGaiTGGXVOjHH1wipgcTYAs7E8GmRc1sXASJHwRm25eJ6PMt3dKJF8jFwmkYlX/w
OI8auk5T7bk8UbNaflNqO5Y9QNQUagx7mfHmkJP0gop4WVUXjwZn8hkEs7MvJXUt
iKSccebXEePQfeH68cFHSoNCVFItN59KhUbiqdqllnT/OrACO4WvY1hs72MUgPEk
JCfiMH0tS049/pCin9WQ3YvLkCme2LDTi4gFrd+L5dcvFkfeMf1R2hgJoUoaameT
TFMnnYflnsj2mrnqsK35aEKHh52MT78m4qpJMvSDgzAF/L/d+B3V/STKMRP8nmBZ
/GyE5w4rgBfBpMYGoQMhhyL0VTqhZ7s6Ml8FKX/HVhH52gzi4KKgn5M+fTDPTraX
mFeGUVpGiLBukcVd3jQvKyE0Pnv/B8lCKJsTSS+LHDF3YP2PFAe3713pUd6cs9Cn
gsI76U55y8X8xtFAf8JSz33CWz4Ktnq+qdaJeZ9QgooLzK7K+PxaC/UNIK14XVEo
W7Tpwy4NWjl1m4Vqd+thnvfoXcH+a+Grep1u3CtinIE0mZnD5zfZbADVg3dFB65L
JeeDmFSCNpo33Te0b62d7322ptzM93WAWpm2+5RXWHGDrICcjiFrI5IDmM4OGwWX
l4+lYzGE2wZSu8Ug0oZ0M7kcSPVatNbLCxXpiW2lVhfj5zpCdue0xTfUVuW/UzTr
9MGPRXCN5zirjE0qgJ8rguvuhnVkXIilHH/8RhFXs8ExxsBWrV16lBvGnE6jRgf/
pjEUMIR3Dgs4W+NRmY4IFd/gbtMSy/glAYHeRkoz1A75yvkIVM3X1uCaKFIR6NN+
yAfso6qsLAy41OZrl+7C/FQvTYNg6AXJJSkAP+GPgcA/yNeraWhKqmVAU+SjjN0c
COGzJ7X1uRGinVQj3DwQ863L6AgdN6OHXxAarbhxxtT7oIHD/mfUYJY2E0jE314S
V2FRN3d0R6uVLxNwXZJbEFGr6wtPWMbHp9QpNFCEz11wPHU1DkBeMNeMV89cH2JU
riUMeSjczVtufw8XcJHW5id6tURSglZ5p62KkcgfOVGlXGc6/MnrTPWXACZp3yNg
sLXNw5nM14wRu7kWPnuGI2shUi2azxHM+FaLST4b8BKpvQwzwhh5zsxdxTiravt3
LdtsNv5dsUgC/GbpBmO2zSyQa+oEHXINUMZWru48LpNAvidWzwNPCXyy2SICfI2T
EZLKW6GY4hQMIcCz0VGwfQv0LY2Dpyy616zo0O4T43yDoYYbMgac3VYKRciSPREY
TxumMlerrvfvA6TXkxGlC9WLysUfpwAlSfgF6xT0JyfV+/VXlPo6V1spgNqkwnVL
TOpAaMlTFlpF0lLrTqZDlVHYtVDrtmI8wHStooU9Q5R+Wsvtn6RGO0f1NjneE5y3
pMLXJh1BjMIlx5BXpIBFufH+ZupIvyz+cozO1V9VH/Ls3UuYqUyLvrVd/vvxQymS
eZopLqW/6dT3wINJCiSbbEEPD0xw4Su1QE8dbsxOlnr+pMHxGg+PKT0bLTTIqQ2B
7fB/9YOEbzQav1FqXmsj0G8jHJd3/6o7wMlo+sn9KDtimh5XGh+qOxuTDEVBZO55
xdsBAkYOKo1Lor6Q5JibtonjsySC7mhvGs/8UJdF3VhuqSIleZq9Z63J6wtT+Hlh
dsf5S5xyj+WIC15JIeWYDOddHI/O0wFxzT5jgAwka1yhhbbYyATP6/8Fm9J9PxIV
8nhvHDiO6qwCh4J2wqJrBWJELR8eYFpsgDamX5uwrNpmvIo6nO6SCZ/2g0DLEQvY
wLa00YM9wJG8HOdP4LQUWh11A6ctjTbbWASa0LzYC7zJignHbaPOqcWnNbi1/VZD
odbK4KbulCyiMgbp+8DbXLaTyPNy+oG3ig/3Mlm7Un0YJxkCjh4gq0ELpOdhiXzH
orvA4Gxo6x6xRYV5oWHOABziIu1UXKHUFxLS06Ee5cDXLLPcBR4fTyBXu9qt3kuP
UnUxUfCsi62SagG0MjxiOQv+aU4lf2NWGp6NmFJfGeYCe1u2xBOjxJP70n90VNqX
OpH/ko67YKAnGXF6Xq3QtR6QXLd/Q/lUzNQ2tB8LZHhYw63bplfznv2AqrvKWX/o
Li3DplY4LOkujODpyZWIgEpKaQ04CwDtHImiDZ3SC5u+zOBP4um17F9VY370UFlD
e97KsxGXFpF/CF/LehaLit5Xm6Dh0jMvENyVhi9sjur2EauR4c6JHZwDw39MvvC1
xDBNxoA0AKMgun8tF0FKA0io3vHFDxQOZS28dFrvXu6WbgxZNTSC9/vueOvKz9Lf
Kxid9/9cGQYHFHbAEmcfymzyogCc++RwsL+8MIBWa6L/WpkVYG7oyoENuwWaorwg
fhbGAlZlLeqiFXWBFaaEsCWm1JVKW+A7bf3SOHstXtb0GPc6dGQxxCKzIqdpSEKO
0HQRk+d1bg0Mgopu+z7J+wHXe9JhJug6z8REAIH2eorntH8XX32+g/OqPUeIaHwx
UcJRUVhTde7xxcBFDmj8AlRveZIHxNeSnXH481G09HO8HMdJ5Zx5XLwgP7dIRFnB
F471zDX5MxbIlqE0OkBUbsrNs/mCfIIQPt/APCx3XMYp/lxilqBlLnTmjtStLyWo
X/voDa4H+im2xFL74oY6Mcxc0Dc4b8yLrbZhvcKzZ6gU8jnZ6yXLeW/biuPHDgYi
RdcB2PYq7dsskShbpwWqMfNLEkD3XuI293iDEdwNUc+Nq9gPne31Zr3rvgeGVCo8
VBkHD2xeIjTcEPExCQL5uYg4DNbMfqnKKIsjiHcNjeTNABxfIi2j2cfFzBLZec08
hhvQidu5ohRzBuE4DwvPu4g49tepxi8R0iaGPi4VUMUhp3Walz5HjpvwEtQ6CwQp
6J9DfuK/fdYUiGFb7703BQwe9rYhEuAnziH2TYWk22KwDwMqoblhXmQVO0H/9Kkg
UzHKK5i3HxXoKaLGQo3YE510DUIY7EszUz0m2vI5vOXPg6S83niOy4A5s4Vw3Oxk
nkOdmOUwiX0WUGYD2cQQ5uoCMbyWHwKAOWzTPrxFlJsJ6Y61d/rf5FdF+juZV7IG
wU9OQi0fuLq314ISYbyKajHxTxACcCZrCdKgh+xuPFLa7Ukg+YQBOWKj8oUnn+ba
7dpfsAvap3fLxCcPRj6+htrf04zRfuDQVAHDQbU2eWB73MemwvY/qjM9/6KIDLjW
0q6hyUIxB7JVFUGfIwCyTeZkzCYyIyAem8Jxh2EsGZVlowWmnN9JDJ8k6/WviDsN
RPsd2TFHMoFyO4a2EqnyXk1hODYJdsZiVrVrFfemQm5RWUTygZ2k2Znsa5vnoMJ/
4XGnYPSwXzuslJnwv8IN2QmyxfTLZZEQvi5keA+rdvWPUMtqj4BsYwqS4awIgKI8
mXG7WTlXa4FOEv3RPC93etNeN8xvGRxKXENcg4vXqlRHltqNAha6TK8JfgXKDKDn
ptMWsLzspVnoAbfGk/TbFok7bNlwVJRvTTnB5D60ArVSyeCGpt9CKQO6IYgGBJYS
vwd6tu6t87OK10TROaQAXQae7mZC32shOOD2yMycFyVtth1sXW347Y2Ly8ISEd8E
TwGZBv63zHsP7XJ35QDYxCtBJqheH+0PcTNA1aJkkgm8gzhf1epWRBkDiL/6pwoB
Saaav1r1rPexUTX9qDlaB8hF8aZcTvhrlpWCXjpdMxPi3vRc9nvt6a6xzIAu/p7J
+FdQW+m4SMTGWgtbIxlinwgHMNnDSnmFEntL7y7Qd/t5rknd20YS6XHFeHXCEj3c
JZ0bxqkj0nhEb41k975n6gawO8GK7ZB2goYf7vw2rUgqFgFw5c2Wyfw7Agvlva7z
or+Gc0mHhbf5bd3Q2mbzG/NDRY3vg1UIXseR2FrVQp997X4cUevOOxgGGtjZPT8u
TO6mb4RMUPAjY1h1/RH15ONMJpUShmivFKIyqW+yN3d/my6KuyECDLfpOkRX7jOB
bvvzmpUjtfTOcL5JzZHrCe0XATWYlDai++z9SoK72bDCpekQr5y5d+bBeQtjBZpV
bGmIjnMYyP+wcTWNol9lBDVheUANRKgyjOr2dxHZwavfHMbeDpgG+NZjQkP8C0/b
Rx5E2uIKW+HguEesk0hhz9gHwompJfw2T3Eu+lj0ybnRrYNyBT/WmJ2icMn7kkoN
lHvUjSj7CAR4jQFspa199GsBYViKlKXifQ/C6mY25bCjLh2iKNdl2LWvC4oVKqHu
cVCbGzd6hLybshyURSo1POIMtwYcbuwNPLBzZv68mrjAHlqSRxouwWWqeKGAJBPj
UBRbjDwK3PDTHz3vFIBMc2kzfzaFP5xJtjnBfs/tmq3kdbyrGZosHwIvr7Oec1Mh
lGxG5E2+I9ot1yzuPKomj6xL6O6jHKsVFbtsimwHWIXb5s19BLDH6HYroZG2iyoU
wJFvRBEmBCyWD1Arv4zDVsN//ky3NjSL3rHnnt5RRtJagtvtxyEDWZQJyAfWa1as
zxxKUIjTTNTB8tODHSSP5S6sC2FKidu15TbBkezOV2BKUh1l96jggzVRNjyhfhPd
g7rOfNJ56O04AB9OtJDAtt4l1sNyPKxnAI69adT0DNGmhZkjiCQhFDa4ZwnA02xA
DJ3NeunQLZFQSe4zFmxvzePxaZLn+n8tSrYrf+f7VHSFb/1JKygnuWL0SdiC4k1i
A4aOhHl4EtxrwuUrZiJVmevncMzo7bi+BZkwvr533+ClCuOhYzgmMM2gtVQypOdJ
2oYdwmrhwR5YZ+CsK4DwHK87nbL0Ebhn9io3K7R+2GJRTjkTBzF0gbitBvi/gMsp
ZJm6vBfn81fKwo6+Ctj64Ensls5M153+XyGrFFGZB2ViQmWX757gsuMba2Aj6uwq
dD+tKKjIBn8iFChY4+ZwZ2ZHg8e+hsryXuTyuAX7Dz+rgB1QugckyTMQhN5qSE/C
Nt/kMbJAZRh9auW4abIKh055P5fWSlKfUEuiH1JSppwesR37AfuqVvAkMWf1cXzD
nxZeUUx1UGTykBVqsfEZDIlCS5Bw/BZt2rOnvRKdo/HSFXYK8OGFNiyKOXmLk1Wm
+GnDBqnfOcJtxYsVMSjTaauz8hSbSE34v+ol7aPfXMMUjSiSmgmUQ7XJzOfN4T3T
55eVazmTv2uATnmoy2SeASN0PlBzONAUkT6jihq7SYzw9WVY4dazc2+o4FAImAdY
dPQYUGa0HzIkpbhJb409XdR/trQyHkrarMA1rkYaqwv6CC8vf/plGosHh62TOC5m
lmxen/83LmYBFAet/waIar8EnvWiV85O/qfJQpg2ehw2DWWH5AutpiV84RcPzmrp
vRIZrJZSfMvlmmWN/gfVJyI5H1fj876C7OH8YR9DT0gjxX6g/nM9FCaV9SLomp8L
IcS7PU+IRX/oRuDAv1ztEcWplVHI+2MZGJofVQ+F0Sv77T7H3jYXjY8NXsW+QRIu
sTUqcHAMFp76d6EKoSl0AmYdvMlWZcXlO9sTRDXTSq+Fx8cL4zk2HQvg+6e4x+nd
xGdGj4swBJLfjsA2Kh5LnMoG0IEH8FYX0AddKr28NXYcYCwbNDm8CjjE+UqVpAI7
T8rM27XfBQS5RyBq/9SxAZ1os1oFxdosJhPHujM6Lh4UU2xJZWOsp1sAqh46R0Ol
LRtrRgF9Pj6qC8QKYowgyFTMCMAhEzC1SoLdoA8/ThUdYk+tM3F+0K/8i5gLGHdz
VkAwPMoszU0Kod3dn+Bq3m6r8gNgTPg7eCBZbvppNStqqbZqno5nqZrr/MiMqOk7
YZYUNdlTwM5tVdisrHIFaXLqbfLWzOqqq4Odq23IHWmlI1mFqsD2lez7rHBol3FH
3Yz6kkTi5TEv4lp95j5NR6njL0yqoebusQzi1gcV+ggFnDIZma1nqQZ57dKzzOyg
P/1c7lzqWUIF+BTfj26egtY8xVZm9ij5fzbHNxypSxceJHrxDKXyN7CJEUq9Dt+Q
gnot2h+Xsj0szaXNMmQV0nr+i3BtjIZlxU8XJ4LTTG5T9cowgYWufoAWBvGUrJ/h
siUeKpa9w5d/jJ1JjVQ/cOVARTIjk1R6oZlr0I3SZ/a3OeTz2QK7M06bkRxIzNpO
XcsZ8LQ8BCla0XNNWNQMAHv3g706gXYP0G/3Yy4qsNzdzreR/RoCYoSb7U8yvllo
qQN1lM8pL/TpvxkJraG2UKU9CffLWshXAoWhGCkPHwukZJdLxeids3RlGfVMwW5Y
jU+bBQ79eyNv6B8lb4Rw0GzmDqa+jfc4D+MTJz8a832zFwWHoT1ygXi9SB1veOWU
yaIPiJzYxc1KUYClLYYxpLy3IobAZek9k5sJQpqHX/ASAyfpFIlvvVjXiLoMZ3tZ
j1k0bV/ZMJ6P5R8XczzaRf9e23IenNECc8cnJX3HkOOa4hd3VyHqpS+UhHnJtKAE
/VwpS9dIzalA11QTQ/iMDP73aOIKnaagmJTR875qRTXRk3Cz9KcbGjw/wHYOOuhi
Pxb8ypKYCcxka6SH1gXn+wrLPH4YUoqMz/0Y/BsqpnPoikXTeMbaBtLXP03UnXKp
Zl2LqdAM/7xsf8MJaPiAE3S8jPnjEEjURbrvb4sXVGpXJEsvkxzvbt/0BIO2lKHj
4udgO9mfl1mK0KlF+BqjW3lllMxT7Kd0jxfwzFCb1s/Tnm8DiGEN3GXaFLfP16BB
4nj9/sUrW00643DZowWUfPVpYa2zj3ZmlhWLsLInBRVGY4UHOYAuPxwRve+rYTRG
xaKpFD4qkk3CVpU8IgE8kcCaTjm+1R67mTxaNp9vB1E5QuoJ+WWd78dwDw5oqg1k
JAF0F+IL27x1mBx/IZB3teR0Ibkg4gbrhN2Iy7apXwcxjs83L8XIxHAQl979ARRq
3TDtnGt+EFNYOxJWx5JyZ5GHUToz6OU2wG/xyolIzt9iWcCiBkXyXV41khW39DRp
Da9m1wizG5H5hwwIQwnMrVKyhnVBmjRMexC5IeK0PdC4VEEA/WLm+Y21FaMpP0Hm
+UBPiUeY0ioTqC6SX8K+kXQ7tEePvzOhMnRwGMty/GWp5ZXU11ZanyM41a1kCN3p
CmxR/1vG9sdT8RGLBYk2PkwTFUlRBflhwEKezEVOzXJEAwktQCVGjSQDmGio+9g8
31qpQEgb37isxW2Lul1Y4apDuPzQjh++Oh2yvm1ursxxC9m0WDtM/iEOGsdsLpNn
Z93CSH33Cyb69QLx9JwtzwIzqS5nL+6FPVI3A6s4kKSffTwiTxoQknH9BUeMJ41O
4bBM4os1ySVfju1W/mThIYgRYXFoIpaNcX9ZGCVpFIiDs6tdWfb/tZkHjvnUlpcK
SL45sYBbkjqQLjUVk2M3DMppYRBGshXdDpe7LrhAhURafNNhEyJ9PzN+McvdT+iq
3Dvi2IOXy/6gXBhhF7h7v7jMlY0RGGD3f3mstlGpk6Y7uZTTtEizOqx0mQbJBr00
Byqeoo5S2iM7H8KYpaWYSuSon8z5feev2lO3Ddf5e5mQXztll23OrKwkPa5v2bT2
VbtwwPu9twtTsNt5lhgcnlJzLhjroPkU1mcXk8+Kdvj+dqUaqzjZ3yh6TgeQR9Rf
vq0n0O/R1rm3LNf6z3CQII281UF1xeg37/QHmsd0eTHTpAhVisa6uLzP1qqjDJXO
HUC23euuqayqc2KRKkX38tcg4NeZD2PqKY4zDy+GQ1HRBMUeBHtCliuptt6CEebR
HARybLUJ0shT9dRPT31ayFXwkYNsHwnqVXjGR7OmB1bENZsUU7mDCQop7WJVVwRJ
Z8YJ0Jp4RvU9ZOeuxt4dl8nlEMmPCGjh3OGbCsjk5Ey2yJYr1GluCJcYIJGSJGe6
AFVj2UZd8d/fOjAdExRCHRRVQw/COIHF5fMEILrZDzdTDJqzQ1T2iwR+04ZXT7VG
H7rXLcUVQnojthI9OTwtIGeauUe6OO4Kqlgk4W3BvUPutj9XklR9tVCyowAE8AMP
LQjkbbGWB+NRbDu1U15Sn6K868bUCRY8/X9+yIomisqQTvvNJAZlDMgyGkqzn0Re
KLs6x5PAwKbyagm0o/CCpgb8xfPrvSk44tmPXBzPbk6xJOr8mD5kOvEUrHc3bAdn
sCmQNNIPbp3LPtMrzjSsuMWSgFT2IPB67XKsSVb/csOOI7qzMx3kMqtnzJVaeBMx
LLRrS8h4J5RBPgzf0G9zh9qSmy3qaBOt8HVtSdK5q1R2jdTZN4LeJ8Y5opwdAHgO
HU5SNtTKb+pin7umpGZLh+qN3wtr/NmKIOCu8QIRuQ02MtrF1dRda0vsdUfLWiqH
9z3oy3uzG0nTOVYxrHjzR/7TDe7RH/g36+CmNrTo81kvNmLQmQrbWyVxVIxWylVq
DDhbkAYzfoc75Snb3ATQyzh7ewh/RF4k+dB+eupCiMoSBtWXdw5i8bkv7kANVXBA
QYadtd0ik6Gd/AyLHxAkxr/AnfvOWx+c/rc6jT8rv2B3QUq+/oWWygKpn+Bq+Iex
tBh3X6upkQbrr9bXXaGGWKGp3tAwSxB3m5baiQbFNOe5xNWCbi1MCgVxNj/5iPnH
ynTFkywzXFaLcrBlHtOp5WrliaakzlTYk0mkTI+kRIcoXm9FqMqw1iHArOJbGtdv
AdYiOz23W0kkhCQOwFMSEHOP7gJ5rEapbJc1qmECebLDmBr0DkCH1WlSRT6585RY
gkl2c6XC3FbYsiSQb0TlBSIkbUT0A8nK0RCdwsVihJMvdeaLAranYWY5tE2U10e0
gA3WD7mubZRi7SSb4N5SERlxfAg4xEjdoZeu/9UBphpTGCgm2Rk6yoFm4bJ2PMx9
3qE+3m8Uus15mybBvDC2Stj4RmPrGEVPPAmnDk1/B9Ek80SFtGTeq/mKJLNNW9/N
1rC4dGAY0aCQmtDDbpbG7hRilpBF6Vwe9qiChYFWdy4mVeIwPoMTO1p23PRpLa7p
WvARE6QCfu0qgEQzZTpNnQEDp2lQ0cRu3nCZIoAifONKMCqc9b0cLEOH52eMtcq/
ARN99t8gsCWt1+qGHQ0afGwXh/8GMmJ7RRIsbtRJdVXYO6l7cX3aeFuPp0H0gmpg
jFo/MP1nSJkTTZLyhFa97EGvW6+aVFWsLPz9mESbSKfXQAWU/Urn9cDQQzm0CjBM
/Sb4IMc3HBq7R2oWJMY1efsIRHhgyTNtSpAiHf9TXre9bjf7fJVxyOK3GxfSyLAx
FwJ2wOcbbuaW8qEpl9iZnrHjeAmjsMaznNgpRAtU6QlPA32HyeRMg/W7Bnbs7aFT
sRxSph/7hucoDIZ5pm2rN/V9LQLSc7Lywu1YSudXOMbtiA+CKUFSFn/0NtWN7buw
xJgDXpfBlimEa+7tLdGC4JE4cyPb1sf9XPICgr023kgfFtmm5vMuTCi9HubqEgZi
1hZxADYZrsjaoDMuvWkjPSolubeYwd0JtMMhhSn8AL8zi9Ohd102BPPhvlvtR09D
VdhpLsqmL3ow9iDu0Lny5T13bjeY6IGLQOiNP6A4q8JwqGJ2SzkXRSrO4BT5t184
6zXfRny4KwtkQWeM47ipyIRANdcT9dnOYpCuQ0FPKHyvZ1Fk0KDyt8/iW5RnRMkS
+Q394EkSJzgOddfsgyaIFdM9iTsvVmqDu7YzatAozCGHdGeHolKMlOQ/DKkNwDVI
nKuYw7tN4aobDJfX8GiUW8++gGAgaKDe+389Mk7g/PRNOGpPtzZaHmGwkiFzYm33
UzzZYt/dj2ob+gFnGDb6uFYf+q6E/hPW++3hWrAWgAi4o6iKRSYF04zYU4zeTFiB
aKMvx0LlDx2PdaKsCWciAqUVrxk+sVmuht+sBT903RCVwA6EH6hGgUYLPzapP/tv
vkLVpwR/tOWVONP75TxauG2Ri6c4zw/WHFikiqLwJLdkWRoUudsK7VIq+k0D/JKF
c0ZCNDgZ3pZdi7Mh7V0bLS7V5At28OKDZTsvbgyhc3+50Y478VbqIjVMjNbRhswM
oBKWCp/1QDRWz1E3j6T2QWFEutUK3T0Ev66EOyA59E3sGy+yr8pAQbOdrpRlWFjv
hUniZKedzZB1ZBNNPsf/rxWOXFbSrpn5uQ23+xGSYZH9EniEjZyPsjwA0ZZKI6Bi
BasMzecmje7yuzk47TLPkviRdiarLqvBqH13FpDaASntivWBnXkylIvcdZIOkOGm
oyUTAxpy34ywb+aVbgZnQNUPf+oA2qEiOT+7opIhvEvGRS4EU1RQCbW/bMNocfZ4
aKDio/IYTKEwr7Pb4IqsVi1LPsOYL0XDiJK8hgqGrwfMorQSRzSEC2V0+2+72Yio
fUq+ChQ0S/AjR+6Pr5CcdRUgm5s8K6X5Mc/G3hXqZKZr8tZEXeSOkHUMTHZhPse7
Uc9BCKNcPsMImXboWrrSkrnsTXjdGFVktLeglOMQGbAu/wU0y6MhJM7KVfJhCAHa
I4nnYt3zIOoAxY8icR1Bl/VkevPOtOSQOyR9Zxes55hh5FIzsIUFaTe7b/YQs2Rh
D50PCR6XlFkGFIoK643J1EkwUurF88Dc+2maUg3idsva6/upO6+uVmHeaqLuR1qz
+BDLwdefLOgX+SH1rrEBjvAGiPo+7DtVfcq5VcXrAqfOc9pv9/GnLeJpcaCBPKUi
fSnGnXGH/v5m51g+dTjHLXfvawANGJEp7WtizfRTVx/YX8I80E1+ngOIKDycntCM
8KcfoY7ExtGAW8fQMkGYwqhQcYcrUJioXh3/cYmNdi2giNiR3H9ZemJso9rMHZa/
AuuDFwa50I35IYe+72AL+wTMiqEVsHEPeJ4YhxBaCRKMnit+z1pvbsMHD5HbjTI9
8gkH1/0OhP3cOXIQ+KaMF9Ppkm3eY+YKzks0GNCaz52blAWhXNKiEqTcdrytmk+/
Jkybx9mKDqKEH5W1Dm3TKASkE/CC69LJj+LCLLxtb9nEuodtajLLEhC3vwUWdt+U
w8jwc9vsHlewOMcl7U9I2zGcN7etd0eGq7p2JBp8G6WqmuEO+1NL8bbkoPtBdWOL
c8xOGMR89hBnmVvf4MHePX7/a2UeiY/jqvvhOXKwuH/Bn/9xJUGJlIEM5fMcJDHo
yOimZHqJVBlUukXwU35GqGgeNZgne6GiAeEjR0wEG0zjzgzE2tnk8nToGtgAnjGk
sdwvLcSFCFzlExiIxYIQCEKrCBuICgpKzZKtUSo/yReWgcnFJflES5tgEJkl/p+8
PyBjYdCAbheie2uS4gg7Ke71XN8Ixy25RmCk1VUiBMVPdAUvm+y5c6EqGNGzL+lC
l9ropJNpP6QLSOVtfHC0PuHQwqQeqjKbHpWXL4Lfb1Rkbbtjo5oDzQAxbWsAMxQt
bRauPvbdD29aTvdTRxNQ77FDN46tMlRXRcsW+MNxhqBvO6Kpy67Kcd/1W12KOAEq
I7eWkPw30WVJwyrGBPr9WzcDIs0GZBCdMj0Nh73Bqu2nYqTzwmsYxcJtv4fZ9Ja9
kovL9K6JW2C/vpP1I4A0E3uPog8qX8My1ocTm6T5hIev0OP8MCHTeGcEyew6NV9M
P9n+aI0lpNJxH2FIqFrGhEb9cyIYY4Y2lm6aMwiREqYwASmW9aODSv+U65/Gkwx0
8blelHftB8liYfQ13Mzq0OPpd5N8kRUhoxfgiAjghLo9W5Isjf8ZuMuneS5UOkJu
kHHru4RwXjTcqsALRHBPZ2tRqFVyWG2A0zQoyXyee1FjjXlv7YbXEV9hKlunEu8o
DyO2Dcias0KpHdILNZAbI0U+kqPbGQBbiy+ZvcsUwCGPceQ145XCH3WYcW4kjh4F
2pyJOCZXsS4UaSxjBTiAQjU5pvrQ4GDXOV54Mwge75bX6KPaHGUfJU6Ujv+79yhf
1Rrhc4OZ466P0cUyyS0nZUsBSrGuXm8keNVXHpGRoqfmfIUPi71lMGPUKx+OGM5Y
XSqASZbsDvnwoNAcex3CIiEGYfAMjy0CYhJSEE9f1cI7TqfZeMYOqRBeqjhuMqZq
JXcbYbyOsm0ZJQJW3epg1hGSCca4lHEK8qDcnS+Rar4SsJHNvumvi4wP+AZos6qX
++fbAUtV4KhBLXWasfS4ARoRlH04dFqS/aVdeJGaicMq28bC0LWwkAwO1kslIKVT
0xMLRiqx7QV4v8jDuiR4XMvJ2GdSetpOGyERMzxnnbLhVopwQAWR6ufZnS6QBsxF
mQ9JUrzjFwAm59m4MrJjiNzDbaVWlFuT/viBJsma32cYZpqUopwXKbMrFqo3e4ZG
PNs6KRN9QfKFtLdPlej7E/2bnp61j+j4D9QnMSWXZ+PRmAdiufJ9VcGGRTKWj4jO
l4i/2YimyeQAxIVCthYcQwcQLtnCBohbD2x/S1JqMh5Veb3rwLWVCVcV4YnYr1ZE
W0TgTPH87Z01j856qQiJYxLilWsV5NfRVFZUi7w1FwZ1IiPp7lqV1BhCiqP/eEFU
SUwXLlXvC3lufB4WswcSjG1i9jNhx8mtjKzg3lsGEsIIKLmxLuEqhL1zCu+CFgJ3
onx5dfI/+SyTUx4D3ItylYQRx0Sxa5mPfjLcnMf7/9knp84zi8T48S3c/d0SEZ5X
VUHRNIfUho21kk30bmuLHuWEaUO/QNuXe6Et3zDQBiHwXgpL93z66cNRdycE16Km
WbNyYtzc0Op8kTrbn5VG3uO8Vyn+EBKGw7halWciLqfdsTKfD+3im6PRwhKLtO1x
VVa6jhsRQTSv2wN3NgcDJ4LT1JBRRfe3OX48dCJo6I8XOgD28q/Vt5h7T9O+02QN
yWh12IDoRYBcLgZJu/y7WI6zleprVzjurtsfGa3w46NNY6qjM2yae/N8DDR+fXy4
5Zpyk2DCuHS8eO+WPBLms7EYKx4OT2jVD2EvRAkQWy0UK5kSEa2j+4LX6/QJBGHg
VAwsR4TG7T0koEByHIEnOtkiPu7fnSA1yYppJ1VcBtccOoick2cIWF+VPQeh/y1a
u6mRJi54PH7XLhR5w21Mnzrvtv05gJ1xLJ4zW5RJXHrkzbnx7rIy0x96985Xs8vQ
IW0e0AR0dTIoaP1ijEaA/8BOlxPaZvozKU61Gl7L0ZXggeXHmnOWuELXHpcDgmgH
KvNhstGTAQmXVI8si+GHZ3BLfk6uOnTP5MwlpmrU7jWFCB8zWYE6XP9mtY+HXu2d
sJVcR6cA8g0UeUaAatOKndtqEkwV3kp4CA3420c0r+kl60dXxMGytFkaixGRrfZ2
5DvDQgI30JOX0/qrpPrIfAywX/Ly7GIdypDT1JXc3HDW/cGbtZX13xIC/G8ltijB
EOWWXle/DtatwWJUYzt1LxXethzZSMPPw35MIoy663UF4JhU3+XYfYuWQ91mkBqU
7cNsjJNN5XyQOlqDT65tgoNy7BFvTwBImnQpC1AIfpVr5U+rgGdO27v2qKxSVdwu
spOLUsf1RFgWQkYgICN/hLkiurWV2M1IsqO7yTzSJ0ioQFKuSDC5R8HugZnnfcjn
uSh0Bw88k81aWGVd8gMRSgKDO3lq49kyN/8qcNIvVUDyYWlUqo1sFCEcvNidlRHN
ZXz4uve8ZkKwBQBxmNoLoU50GYTUbiJnPNn0oVE675y5kU2V9WoMK7C4jnWzSxum
3qvU+kH6BJxtsFGqv8P1kzbYABZUO86UNEh5Vs2DbfIf4DTar6HFfYOSaS2OXQND
l256cXYi8eakzLX/XvLtUzHyXrtBr/AHwuvearAloT172kI+H0IDGCTd2Lg00dtm
GCJS6CY+0MGqNcx7/UG9SEOmHos8/zW2tgww82W+BNd5RTrP7WBWyv61IO/BFvV4
ocC67p60e5+rOgluCEXcNSvotjUD5z/i9l2DZF36O29XaYJ7NDdnuC4yvieLsA8H
5N1eSlgKgOWtWw8TscEnd8mGftC0wp1n1V7W0om0n8DOGmrb453g7wV9MEmks4ov
zXAOtNS8PFu05glUYwkZQ96hIixX02r7W2sjk1vyX7sMPEAMl3wrypouG+KkRB3m
2VI27kIQTswEqle87U9P7/C6r3PyVU4b2Ejjo0RDCv55bCgaNVu7fz/CE2Z3ETQv
/LOg4qvA20wHTwpTVMNUSlFH+g6bsigmAiUUr1Pig4YWK7bbZDBgSZZ3un8SvDrb
E6Vnz5erWm/E4YwZZwFsmrZABNDMHJs6KB4trvN7pR0/H1OavQfmhDcpJv0JutDl
qvL2O6ogLzT3PUpwnjhYKo+4CO/2U8yIj3JeAH9+aIOXi9nZl4cip2jUz+vvsjoy
JS/IqO98/lnqrWlqzQI5tnAbLRS7vl/RDrTgYY4M2Fd50Y2t77xe4nYzMHtuUvBB
f761qUunc7NeME8dN5ylmRg5IuoKM/TcWKYJkHZC499+tAhDPMwisG5hizQgQwH+
9U8IL/eDU83OrjsfHjOTdUleAeMREaQkjgl840258Z+CXrIPwQK2EZOct1zJi+eB
B7I4XW/Ap4fVYsVC5lKTinXlIZ8efPElSe8+03Zp8JJ9TOUu07l6dKi5OgUw99O/
YhsZb7dPJAC4oOHh7MRbm3Jnwd+tgmOoZ9tSZf1yfnQz9640E5T7R2e5WAGKfW9P
aJsT5L5YZkTMGVhjtfaSdpdzHpHIV16nw3WJ9FpJLzNx11FngisIKcWqVf5wPsq6
k49Fs4kgYFev1upVO2aTXSl8cCxG5s4wip8mch6D+OlaIZ8LL/s6KxlPclfVqtrH
htxsf/PPTrPOzwbnvZ2ez8TnaywoVpR3d6N5HqpXOM0jfAYJTQRr/RxchnM80zmf
aZRxRaYciiR6O9yITE42AqZ82l/CqECYGPZ0YmwV+C1yp5SIKOxJAD0qSejvqyZ2
dgLDtLoU344126BTgqYNjTb102xSkkrbOP2ZZ7xdNLn76a36ZsSMLzJSulwrYh1s
LFB1UiupMp5dvvN57ir7rEZDUllEvuAIwHrTLtawMy3jBg7ALAZjX1eLJg7Rys1J
3Z7xBgTarifymOLWxus2jy5HohEJIDYCK95GH7+i+K72C4s8+QSWvHOqMSPI4u7a
77k9q5qHmO0dzkOsTgsrOLsX7Bi2U4CcyDNBsGg8oFNkMpePCuakpnkBod71uYMw
yrXag3CtXYddghXYgh2NPQ3XtI6D9CQAurT0LcP15ohjfiVL5UFjG5ItlYmlpENc
pv93C4PZFTxQeQVpJu1lPdP31RJsDzlXWlYYIi+CwUeODexcrIKiicmt8tHfF5nU
CREFtI3QGsLZXCNsuQbG7eqLumJNntcNVcBedBgPUP96jhi5XHshtHzRp8XgjZq6
6C7wAZkps7a13xP8eXiydjLngtsNRwD4mwOhXUPIfzzcjKhncrWOE1NbsNHRzZG9
BTwPfujK8PprpBZAGo/3asJD6QxU8k9g8jEis3gOKLBaWAtMBYaGTHUvBbXadkQW
Q9+A/wYd4nme+NgYGDtA0CmhqFF0VPP9zGK0tl8JyAM07ymFO31evo//TCuaQJsj
g1KxfWaMDiqNBh1qQPJyXKF2gUgLcfRambfCI+gw9UhnhSa252KSjo50VM/20xHa
D1sJhdsPONnJ7HZu2aI5/8PUkT583bb+zi09jhO9KFDwUk9L2fUxxHVVPU12sCtj
6XVEH8Txfl8tMxWLeIkwWUlD730epnWdv0z+nS3tbq6JMYdYVYQWx1N0mMF6XuYE
DHoozFJzuQjuXIycnqQDZKyEBiNvSyZNbknDGAw83/cP9FpS4+04pFnsxUuL6gEO
pHZQJ3t+ws688MxCOI6tAb/SvkpZTSYlw3hoR4rARFvOmrYYdTqr/BnO4Ik0MW/v
FvDtibIxQG6QYsv34rF0acLxUY3c/x+l+Evn1iODQB++Qq671MIXmI/O2v2HTX0x
ngHkgVaaN5JfqYUqigxjaBkWD1Z8Tb23d/1nBxfrL3dI3E9kF2IHQg+lZZ6u05na
HixwvllTtOeUAFmyomXnA43CDn/vSIfWY8ekcxKU/bUxBaOVvceH71vzfAJGdxma
HfsTvSso2pL4sHp4QMGGpitW/O02nHijM3SlZvvWWlvCCBHLCPynVIF7v1n9Q4bf
fodAo/+B4A2IR6fi7T0scV4RN+8uTa7AyJ4v9pv+yZ/ubiUF6NuCOZTb/q/OdskN
7NpD+MjR8fT1r3uIn+BpD13ooeIoTffOmiDH38zuLabR2/w3LfjVqDyQj/uMkFVR
jFmUmVvRdRI2k71u7lYL6d/mJSqxMEp1LWhf5heNJRP6bY4odDa0oDmG0H1eJr6B
LFwIiHP3LIRefBpNr2Z2Lf9HKMFS7TQceSFhb6dfZecRDTkJUvzCoqM6B4CriZLY
AYgixxK4HMBHc+zGUeWGsWiCAh135Oc+zPKZtz5EM8+B6tZEjarnFmtfXg+wFQIX
srCR8io/FC6yu4RzK6nDnt5PtbbqIm1B8DNkqfwZOxXt7SKgALYAlO2M7NmCuBTc
+hHLGNuhP1TYVDTEc/MyPngQQmB+UhdvCfhQL/hO2R75yZmKMuUFs9KTsiKg5G/K
HFcnPelAPcLwgqt87WrAetoy7tE2VaCRcqAs8X+laawfPrCYRYxAzxhEIgSTg/lK
o2/MjjGNwlrfJewmalWyEf9ki6WJAR/SjpYH7r8Pj6MtmN3e2d+mUI1jvugP/Ozf
ctAq+RQFDEryg0VzYZphRdDYRCpBoNhkDjCMCZ6uSoJVc6jvVZ/ldRhF7lU2U2xc
Kjfs+6zKzWYQnS3ccwaHAKuWPvmfd15h0UL4ppSPlXN5j6TD6D+ycSfsjwzXGPyN
1XNYDMPr0lHUmfRbTsNFt9i5Lni7thhhuIG0hA9HsLEn89yZ0AnshYhMnU+tCSax
mi+jVTJMR4Exs+77vNCD8oCylALo/MoyPBpZ9HGXBrxGJIOZwSKcCTyYzL/NmHBz
u6ETTWtKSg1F4UPNjab/fJf/oOSj5Q6a3LeyEV34F/NB/mknDx0IncEIhCRCrxSn
q61X06fVpjG1tpy24l2bNgD7Skrt+8XWsLOPRRk1NUMddNWCoIbi0qva2Hw98MCV
BnM6CRXAWi433rI2Un+LsOsy6vKMHS8moT6/h71WKb3YeKegRbC0vEE0QK6DMMS7
bCFgB2yypZe7af2YqGgLgWIgrxt7kvJt9VCNreZTadssuXrsyMzBF+wMrs4WBSf6
tCvwUGMGIdMe4X2dyAES38UAPEIZRA1fRYa8TdIhtF73Pg4G6Nxt71yve7MOMmdw
7Y9/UWuiC4yDD4m9EJEuNsxZPXGQFoxjDd4Un/AyXfR4glHpdf6XtCbRElYNvLlW
dmwPQ7gsq4TGzNiPQrs7Q0lNef/00mN8Ao0vKPo43cg1H/8cB/SjdkC9sx1cd5W9
iCt3d5v8UjIx6nwE47yi7vzNJGQpGJ/iyZyVqesc6SSj3z/0v2czZRTnj68hdiOr
sV3rLFE4zzowPe19FaYwc4hT1C9zo2NuXEajLWNUHBQkAi7I+nU+YdxRU9NQ2V8k
1m32nyg74noECbDqxxMZFs9JVxEjnzbzsJRAmvH39C0gfTh/I426fkERsslnmCbZ
U2j3+KFXRkkuEOjKLjRFFX5g0nB4Iz/lkBt6SLC0k0lKQRGH5z/0iWkd3OvRl0vG
XorFAYyhF+oXokOtnk92t/S9IqotNDoy3kdQAptf61D0asJ89g8tEEDZdcNLfcJ/
Udsd78Jg6joZUCwrBUhF0QG6ffhEpNX8c0xgCVE6AUQoVtT/1puIHyaYXpd/9Fjs
0pI83OwEsk3Hec/eLjFF7cbwEKgUKCDAT3LY88daAIpYonbpi+FaCr8bFVYyPxm8
kQBPFjyN16kZC5DzRzsNF9kC/w6Ru/B5v+Vs9Zb4r9SLKdUhQYbiTGH4Ja/Wvj24
6OPGj3DGRrZVxsWYjcu1mlTsZr2gtO9RLZorivv6YAbIP7JtJM8HIHY9/9Y87ptO
256m5bX4rZqWuntRMDnCst1h57QuyQRGue48v3k+Gzl0OVgsuSQXyj5VMdzkaU44
WbXms6u/uzClyjh7qV6ClZ3nwiHQ/cPNo8+KgXzBbGdsTddW1kEOyHjsqHRWPCtk
gSZ3U3ymbjR6U+tfHYdppwnvgFGWemOwhnarHMDOH3awow9SjE+T7kDgX3nbio1G
YwyzSByRC1f9awrTwIdTyKIjZkCnxCxxXp382ZjGrWCDY0LmhxB1Mp1M4UVipp10
LWtjykRrhis2cJFsVzV7RmeU0l0zhAoiaGDZUX2MmUGzOeO6/Y1e1z5O+j9vEUnF
9I6pXCRU2qHi4phtrzU87GT2ZjsiXlMDkXuIO0FO1Xee2C/NhSEm6T/Br9ZLroTX
zurbhD4120zYqUnT72j/KKMANAAvMDEPQ2SRU4egGQL5BT9cGc7V1j+KIawUBGhT
xX64bYh12bl4RPJhFLcnxbkmSaXx3u4DgTAijkd2lYOJ3Y7U0W+YVzV5SawpjsJn
PfSZ/rz7jS2le1KPUgm+CGquf1BZW71qebtRTIzZvwaM/tDLAem68IBaLDCk6k7H
45CtBcmzN8IB2NgQTCRkCc6HZk2+QkZsRbya8NXHbVuZa9K1293Cq3VbfOy5EDJF
ktY1dKUzqMytRozVrnNdDxx/+mLX01ebUgUWdsFAKDCTLGVF87rCLo/qTBcAosnP
rNdyR13AfK2ZpK/dSAqBJs1SXkWUfJAS4luKsP1ChamUYgbuHQiiQzZxRUavzOB/
rOc43/5PqQEG0q+uDudzxGFdKtGief4e3DV6+RqiJ8s1JJhZXClp/jzZr1kCc62B
lGtkejI3jHnyg99oSAEuZgdn4HpfESl1vfWdliYcUq4XoqZ5lDIjMYmA1C+Obo7h
4MloJYIoz/B4qidmJaZeCoWm6J7Rh+Ilr8o31GO6vFIUvPe4uwG6dHLu01ytw/W4
6PbZ55vBWE0FNJelHbADQm9N8RK/yCq7BIRdHDjb7q5L24xje261WcNaSVFtfGps
ap8OGWN3oLel2CvyNp5vGDXb8VTPAhceSwNKAdZYL0VmDjDlBSAIC3r6bYN1Kl61
N5NKgUA90O+LNBgHl0WCCXy9jKKgYSImEO/5+EDfya2qzIFGud6bG2QkC3qWzL04
K7lIksJ2nUPl4CAJZzopvp/ZYczY9LcYrYBqVko2JM6pGY5cK9GCn6FAqchqJoyY
vISPV+rbxEOgSShY1H3me5fQ8N85fTjVcTeYVKyxBMK6/mRUXRtpUBiI+FL8A0dr
/7kGA96gPlznN/qPu1u6WS86gYzsjByVq/nt9l/34N3fEjJ58zJ4ajG1KEXzok0U
3x5F5q3rrfxkoxffu4zJhRgjprrLOQL4Y/oW1UHzuTwY6/HUoZMWMZqUyGxS51ah
o+sizjJJO4us/d7En+RYI5XjW/2ygssKx7CwoDQH1sW3UBVzobQz0ed1Cy6ueZoM
r2pCUc7sGhRpUGP/RFzRat4EEC4bGp/gt3fKZBdFPOYWqRExhsmGi8Dd/J4nnL5D
JQos4wx2+KfZ2VFrnueOs+zZLWcnluePPOTIqAkuHxtqp4a82iMJ5iXge7ransRH
APb4zaaFxKeyKGHZxQZ5bS9m5mTzhXzOrPPspRMlkvRGwW09dfLucjG3m9754KHl
s38k38cqodgIFL9AOtc9ax1Ro+djk5rN3IY+3u+kREKq6UflI1ArhNjjAzTpPkEx
Pe9ryNEkYccF5XsChk2LOcL2im4Sdktt5YCjp2w9GMs2p/DKGIYcuB9ux/p+ntWK
c/flsH/oA9kvOUuTLN/EL4YBRrvsI/3Rfm90pebQS7JpHQRRVhPj1M3/3HHhD0Ls
GBXH8XgyNz4BPqlg+am8NLZr97OQU2SXgc+DDRVtxw3E7VTHj5CNboeX4XpwTot9
rSEwZHkJc8bwRr+gF4UmJEe0IuPOEXdQQIJRQjC6EQfYS92L9Mj49FvkVVTu2E9H
nIS/1/5qWixS243c+uoDgaK8mCvydjNxbcMZhFyT/hrQoVcE0E9NStSgkrDj+JWp
fdT4l7cNp1mmcqoG5n383KLVhTDBdbR/qemr4qxmXVMKd7SOtJgkNod6iRNDgwWP
4Ry0wGFpjex89dBJrxWmBCs7tMkXlOp58LtaL62W6Lbn/HaK7IvMeMaBFik5G/rQ
dCTkJRpcLZFqu28vSjs6YX0xVnQut5QdMZBi1YLBn0APNgD/BaqaQc+fR2mNAAzQ
L8iy2fWbDylfcOUYp9Yo+n271NQb+LjGdS1Grgi4K0kGzsslZvZYUzxiN3SA2IvH
7njBcs+ow7+tWWoQL5g0ovh7Zo/7q6etK0yydIzWGUG3bXjNVgi/DRMxmvl8Rdoh
hB0aU75vlufWWsqTNsFSqdrPi17Mg3+qoHWUxYmLfsBJtlQV+39MTOZuXkw1vOYs
9n2CQR55WAWTOJlWJ1v+DamGsIfBofjBFYiWgRDYrPX41aCHcO+DuGCcQf0xa0pu
RNyeuy2kA5Vx9VgELmu2l1q4NqKSAkteWfUE207+AQUsjbvoQyguJbiOE8PxPOEI
ZMui6TA9kHm2DPRSITB4rKv3L6afXoxV8UWmVP7K+blKcLRct7ydV+p+nLESgEyx
1t5uWtpGIDiTy7B2JLIRhIiR7s3XEN1c/9CNDYYZs//xqR1aVVDVqYQhAVIkvE0C
TXbONQxGzBkAwtwvHuZ75Ja4ZMg8+J/q4/kfJFewaljCVHqEwWTvlxDXegfuA2Gu
ZUiM8KcyvzZf4oZqp7kid+cCU0WwJlO0X+N1xdpFstLCICImPNj8RcJm5dY4QEVQ
WQ/YLIX4Y7SZ4FcwFIxP8pznQE3/bATRb5GsFfkCafK2X++ws9Hn/U2wF3Lj1/ue
/3LgNv+R3k0ydl5Nt0XzOyOHy67YtyYlVQT+wXiAik16JZh0hSAT9rtIXKEe30RM
CeKjEIk3WX+EDiQxZE+Icwdn8yYp36Jqc8Cy4cKlkp34dXXp8lIZ9C9+He6SJHyW
IpIXw/8ZhAcps5ZfJAgBEFojfjOeKGrWsDef4uDREeuilSA/Px5MjqfqqzUKh+uL
TrJDtfUdFbnu9x5nMGTYw1fLtrXbG0qyFf1otULrdY4BcowPKoaC1h9LbJybY+CS
RlyIpovt5LFcBeTkRAue03osagDH/4Y2hK3QpHiGTFGt1QeDvyJh6m6WjN/c9G4m
vfNKIAojR0fMcf8IT9rTpu/0KKQWFblNNAsPw/XiEJaw83jtPfnWrbvUywuHDnoz
02Ur6jLOAQZiotVG79UsUxZLJ4nsZUZL2TFdAnlC2kmW8+z4CgLss+cvtLQj9ies
eb6oyRZqojDWVBHEcAsl46yNvG1ho4zP+hQC3nZ7/zk445N8y9ArgCw/6xavXVNu
s29orp6nbzZDrg0199XOYRoA6LGr+w+7UJBVFGQRzWE6ckq8LMQUGR/9B4giKtjy
xVjBcWd2ECxwWtL6pSRgtepDJdx4TY5/KkLR9JYMc9/Tt4X4ZxtOHMuvoz+XIDmx
k9HHVqtox7W47GSySve6JCHz+mMvfntwu5X+luwYNMNR9QJUfAuU60f3MAV4VI0l
ICK/EjPkHOCPhfnJuciLtJaFk7mEZc0B2BLBaD2rMqxRTXh8lUxF3jecytmmWZlh
AUPBsx2O2kThYBn4SrT2Xebsn9vjoICwqnULz91gN4QG71+S/45pq0HqmLbfCdMv
Dnf+J+5cr7gML/zetZr/XPYpfHu+JvwFfbTMh2iK23gnOPb7SKhHVA9jZ+2gHVK5
ueyqTKnmFILOjQToZwwsjKhPuzSf0EL61h/29DCUs2nBDVAHB1fZLjJdnTvMXWTy
JMs0npkpnr2NbytZz1PR77MPn0R0O9TGPk+vLO5TglYqPcaGcUdGF0Lsfc2NUpK+
c2ZlZrjFE+Y3gmDX83PHcG1FypC/fWqhJiLd8pncUbuUYpoFjRFl34JEzWu5yuKa
XN8fZYeqH1IBw43PgVImukyubzVzN48n/617RytofaC0KTqS7dyyeZ1XbH9gMxXu
918IhV+sGTjN4pLohxu9NDboZ7+q75ruXhikP20UEM0iY8g+R7Sg0U0pvW+Ie8Zh
opWhgx7GABdQ2WTLGvuDR/OORzlTyv4CpjU6YmUkou8uJHPn/fOt8RuY9B2j7TZc
5wRO2LThKJQ6qPGzckYPM24+lru2WAVGwNgWGiXL1txZH/RhlZTgE8uJAt0FIvO/
gnCPnxDGGM0T1FmrV1kXMuDbOzCdXf1mEljN1g1fP3YCeN8ZbYWOwkMGLl+H55Xd
E69SfKvvn1O8grS3/jVRco6UINx8kMFycXxeiqjF2DQiLF8TNJ2B1rCkGxHqrTOM
Cv1ZMGEE28FZYwGQA4PWuZ8qnzYwajTJN+ikPCx17q+LOw/bXvArhCZp76AbRiIY
Ulhb6AbHswaf/pBnswKdBq6DGe80FKsPv/84OTyN77UUnaSL5SMK4/LduBeZed+p
Nxv5k0Ka62ec1xCZBAOx9vpH/pxdmSQpHQKKYj7F3qRvbYQVo2J/TAKG/sLWEGI8
auzATz5F764fdYIZzCMkixG2ywZ1okDENdTV9tbYDS9sPaudpoKIy/dd3uYHu2QD
NvrQSJTcylEuEFLFxHgIEagI06g03LwE8Ia05KR3RjhHdzz9HWmwm8b88snYgY6B
VSQo30NiSy2C1Ycmw3h6wSxtn/fpwVBZO3BsOKH/KDHI16JUOZTY96V/XdpH70AG
Lk8+guVXCMqj9oGqx4QklXL7n/ipfaCHP9u7NmpbI4na52ZprtbElMcKE6Zh002a
AaXYilK8UflfEPS29JhVOqrtcYZOyEPe4e3R8ggLC+y31rk0KO629CRG8b8hH4ab
mjBO8F1oQirU60zjcgn3lERhUrhD8OFwKjuxh0mJbQNya0kUrclWTuVpQMcHEy3e
vTJ1A4c8ZGs0cM9V5k8jkqfdF2rA7hzhqPDfbD1/Mwn0JDIwV0xRC8SCAUHrzI8M
/yHJxQFUXPMzZ9JENHsnq+dF5XRWcBtIg6RzGMKya2M1Fgss4yK6GQFVQdquc+M/
okdqK5CWsUxqh/2oK4oEZgJCn2nVPZLxKT9I8Gku8JANKxO0Dl19OU63xWaDU7nz
FcrVCcEkkg6R2+CE3xKSUiQYnU73/Ob1iWrjV88RpgKfoJ/4lIyZgIaRxVyRlbbD
hI6apPXe2zEqrEzfasEkh29V/JDBgspDoA+FTKY6XEht5rekpFLV/T0N0gZ+gREP
Zm9ZK2XufJrH3hHCQP8LQO1PQtrGuOTXV8GFoerN72g40QPRaKc901YLIq1Dr++B
ogx5JviJxe8RnJv2H9GoygV4Vfg7mibc2laW5RBsEXHKvI1AYyEbWBoRpUBQgdi3
cpIMn3CPOzkZqlZHKqGQd6nN6ebP9zpQjb3y8b1wxzeMbR4iGCbopx05z/pKlHqQ
MxVzn5Au/zmr+HphfpJHkZxi6MSpkkcpZ2J32OPw1qqIO27dwffXT7V7624uCmyI
sUQjupXjBRmTBzNlBksjZGgw9eEN2Oj7wNzlWxVOAFdQlTmxKBUzcn/bfIJhEZdO
YTvgpJir75TpNOmf/125cfPV53DRHJNjCY5Hojj1ttO2F463YZfEA0WgRYprzDWt
PjgaGv+wryoOQ3wZCJj9nPbqVSM+VXAOmomHo5qV3nQd5tOeQAZ5JrZtRQ2Nayy2
OP/z7CDvg8MVMCDtYotvnS996EnyNYcyLSg6LlDMvXQW1c+b0bVA1RGBNoPojgj1
VRg0l9QtnlexyiPGi4l6XRRJ2jFQP7MExO/LQquA7iI5LWXrCOYyGNhuIBXBHc3f
LdLfrxavtgbK0D8WnQ9J2bPtf5oajIQHwyPANoPKdjd40ZZZ6ulo1UQ0fH+C7yrC
p5HKv6Up27vhcR20T7PNFtY361T2fTRzgaxBoixMcKKGXTNb2rFjv+Q6NVBhWXr6
GncIPUmI1KoPINMNAaQEs/CBWky4krDflNFwQseqoTNnpW6SbwIUeUxTde5OT+H4
zeGwgg7EVcgy7tFMu0j7wFZmdEIzT7XNSdzMv+fk4CUUpQFnQhmr2y3sJvDgrPRy
9G5tpsgZW0PRzsTLZfUDUtTrxH/ZJR3dF666iEwNcIEjHrgDddNvl+EQ2gB8MP3e
Lw1vh8HdamBhLJDuTBZC5nKE+osB51CsncfDmjue3ot4dGZ6lzhOC5/HPlLR/lp5
6ZiU7PuF6aH4Ni7nV6t+VrgYxHHHKrponYnbEEtz21wJXGBpi/TE/BRvor32uPUH
yoRYTQae6X+JePQejytjdEvqCkFvq5F+WItZWVCpMlO483wuwQfwtA1vvRT0Wl7/
3z/kJBFQxoG8ceDGAfm71scb07qKZLm27HEm6agra+yelvEixtwlAroRefAzBcfy
GTyZQ6SbHyffsn9QO/7BLkhhtz9kwitlr5QG0Fd3/q0JM3dKhOts89Xky5ZXfrdB
O9aBXwQxPy2F+yrW68l8N4ZrngZLY4TuTeD3j7iyZ8qvHWgWdc3Yn1knJ6l8EcX3
xcMjZ4QNo97sdpIgLy+sDhfwKL7ox1W0VytEbLAgz+daLQvv6bK9cmrVN2x/5PDR
B5a4DGvj6e64czdJvqd0ZMM6t5+9M9e7IpHzuavLU0b6tfWMZ0E44gaCvsyJ+q5p
krtH1YrNcL5fBLt6msJHGx4ePjYy08HcPrY+feo4YIG1f5dj5LZlbgzuUDLRq5Pk
zFf4hUW+qERjCYN8mpO9yFaGPsY7wy/W9+fiiJvCOVLTcHX+xZUAOHRlzefH4BI2
CnRQGF1jOsRbzngyVCByZQxfOeLUqR0reeGh3482f4UHOdHMgYqfu3yl7Caux4z+
5akf/roN5bNPaUYv996OwXBAWZq4CeTPGZDM7TdyQy/NFI3+8GtFQi1VSDv+l7Al
K+Gv497Qwm/USBOgVWxybgfz0MvLAiF3aEeTG+xjfmOO+YIzaZsFCeboidTUCnjB
RoTRJZ2/BPtgoYDZAda/fr3OpWE8ngARzxvHhNfyFymyKLQwysYD00dHqZqJRZny
vh6ODts7mOkstdYPYNVQBjWwx2MjYq1aXNKL5iIZAntuzuNqN5GjYrPbXhZAg7D0
3CzQLa/y0aqCOQjC1s/+Hcx9M5VK7lN3wR1FZygBoWP66VGlkdyC8Ms+E476grEX
8TCWBp/TDM9PlUZugSJi0ka/yBUTk5AgRwuwnr8lRoJjKR1svwVhs62lXiBcTWN0
fWWqEM93ePEc8XDINHh5sinXgGsafe/riACPn5cxMXIHmw/j7H3yQDbYAMCFiDxs
CQ5CejyyuEQb9scO/U7rXSRVepIwWF9hYrtnBn1/M4F4z1MvbO/Qc5/+AOQLCd/h
sKo0CH/zNIfXxNVMpwo2jVXzxSQcyXX9XtHV7RrqQZ/T4pIabAXc95EEKn56cYKQ
nCEl4DAilBsBNqqgEgWRQ60BWM6mAjhpmUGAB61SXegVDNKZr9C0C+hFVzNU2b7j
ihe5CpvB3ZlfHE1kiIc9dd+/yE6CB3iSjC1iD8+J7/BRX0UJs2nDc27/KtkJTl0P
svDjmRl/R625J4kx5C+wqxqu3ZRTDH8ZUgGJWj9N6LIo1G7lMjxm9KKgSKXHcJHC
OaACA19xrG2l5UPgdbe38xIcJQkAGcPBPfqj0vgIliBxAZuz0xctH1jzBN6n/zkL
MwzuvZiXvPcJqTYTQW9N+rJrFD6Xb/+PBV8dokS/FEGZ7ie2S+aqoUy/ddk6yeY/
8+xn5COA9w0KvTvr+XOoUemYk9lMZj8HWCqqNeP/Fp/hSlGiquS1W4ziK7Bf0eO+
YEjf6deO7kPPVZ4NnPtala1lmSLBkd9UryWJWLlslihnSPxbfmYouqIylPPCeVyB
2tdyZKnCYxBSkYy10bK27Y+08GlSqtEqGpZtVXTeyZx4gz0OJj5wB07vFLLi113D
9Lk1iON8adAwLRp+7Ib9f1JIJc5HlX05md4OBQznWX5gIKxiYZTrfdwUgQ8f0s8g
BpyfXMfSy9xi3Ie2msaEZvUI5EKNZiwUxnArE2Wloo6cOHWKqb4Lbo5LDylNYr1J
nu9AooEPAIZwq0idw94q9L+1diBEaCBmu5lpyIFH0ptiQUlTDMdv8YAUogY4MuRK
ycq9PAZ1q4KQaZn9VGLJHEIAqYux9W1sxhUb5a5+NDMla2o8Djky74Z2ULpQtLg/
yp/zMyRIXBk2VcnNgSGTtdNRMuE6uRsf/G8yF+gf+wnkp/ytKnm0+RVRbA4ql0a7
UdSta32WaxTSpvRQxZrOWuOwxO2ZBgEcTzxCxv/BPkKvzFdX018q8dwwteZNB3Od
WkmOjFYCDagwAq5r5NqcqPIO9FYWMchXJ/krotDoGOSyYuSIefCNFJgZQGUgxPXL
thGpEsldAqKpBHCMHOMGNIROFeUH44amNalWpoxHXfk5qBN+6WwTdyCbIyLRKNdO
3osUN89eCQ9ntlqGJdxyZQH8BIdbpCqyO/NeOMVKEAqp33IAZBvtazr+rOYbuYec
ibVZOKSktCGxO4CvduwcSEL7Hj63MEDIfO6dNDQoBVukiw8PEIaDQe1xXHaG5O/C
45Ml4BqH0m3qSzGQqRj1yTzVm9Sy5n3NwQoD0Nvj1s+AjiRWObqznXRnVHzkSYS0
SgV8ZCklxs1VgSzLVGqD8+Q9ciZaEzTXseo7XORbvKjm4k2gn2XzQtXu5UaKRM4d
vXOG8diE7gpmXeAG1HUrk5S6NsF/lKcDLhhrcJ6EGAARQfUhntMZKsnU8IH2Sv4p
q7wgfqg+q1LN47gX1iEzHs/NED9OEmna/dmV6XWYbNq4bpXBweanylfoGsQ48yvt
BXKtoQEw88wnyoaWh6hEnKxlNPQxfOJ8nSVOROU3N4dWBrRH8ifcQuSWVggN3RGG
hn09VHALWbNP5U3WKkhDaLO+6j7UwzB7r+Ft6uyQCzhMIK3+Qu3YIDS/iWmOiagz
/Qg5nrvKLoQaYQBVKQO3ZjQT3S7K7mNxHbQ5v4dok062EnH1DL8+LSIK5PdK6sYz
BAQ5ZcGaGlhj6q/E43dyfLMogAWPA1MBR4YO73+ytuRABMc4L+P5H/uTpdpu/BEm
oQ1wnNcVfWaLkVth0D7kAsK6BCYO6dVK46ZtP1zZusMa/LpDoz7fwOBObSmGenBN
WegfHFGJHyz6Zc4ZtOnCHv1btw3IGD6B8a/q6U8hBSRWM7jOcuhXdOJReWV5SfTX
/mc6aNvxFf2Be+xXjGNdL2IH0iHxPPb/bNHaeA4vo7+ytaRkcYWQOtck/3JLJf1G
RnB/3gcH86Zfb3ByftKtbEW5htEtkk8zzU1mnaQzY0gqzfQK2c3wivIMmHLI+yML
QOzTS+GmvBCY30vyWYr+NXSluICnttDjv4FdfV9X+K50ZK0Fio7ojYEBfGzGqrLs
yDeTB8c28s0rv95j/9Ab+fwRQnJeYeozJcsaophEiBfVDZSkKcqQG6+MhaFwaBrT
hGMZDihSO7t9WR7T4iYrkOQS4zXlLPoNMRqPGKfrkXqoVS7XGfdqh5ACNpwfVUs1
MIJSgqYaYhKVw7C+9O4SZqos8hgylsapkZe3Hvl921FPoXYpLsKcdlvK4dwHE+fj
kedz+n22anp4r8gVaYHZpj8C9KpcsksHAFv4mqNssiEEvDQCbXitNjr8Gc1qxyS4
9XP5Fa5Ir/9kxtvU2dmFwoeK8QuASSdDoNTM7ObnjIqTxDm/chYilvhSKuSsMLF8
s0o7qVZPwEE+07WnSLxkq4oIZXjsM/ZGjGTCI23LsPKah6DX+zhYP6MnTQaQB5Uc
IO2VappCMTucJkc7VbcYS/V+lJg14o2WW2ontW+Nm2NT/1V5ehRucswtwKOgMrrr
AikkNNChp2psKo9/zwU3ALb5uH03z4FexHpTALkbzku5KyXBQOe8t0hWsh+KAsKA
KMzSw0+PqVECsxMOrJTawtC80C7YoHrYpevbdbGKBgOLkgoro03h51PL0R8GAqSl
5pRgDXbrudkDPmKDzdLbVoQThQLmRgIXs7Il/55A5UUSvWKSzy8RM2j9uFTE694c
Ji0ZV5RduPdokepFTlQ52ZkPiRW4MZLms0D6JNatSXGTHqMp5w7bbuKZnOMeTRdq
o072Y70P7WJK1MGDv5SsJ15FHwBF1q5aCOEoSvRfoGrQzcD2V44F4um+fJieRUnM
toU/pYIL3mPOiWpEtNqb/8c7jVlu2Xe7cG6qEEUPAblXRNrwGYnzy35BTg6L/8BQ
XhB+ptlIvxagoAFuBBPm7ta3T8XFkmVcIOKAoau2ILgFz89xHhAfRuf7GvcJTNFz
9CUK3yP6e39h34kmjO116WpJ4p4cGoZkEbxhe2e2oDUdvzMYXxFJErH47mBQDZpc
ooDoCLXQGZrN7X4w9U/4nZM5lTmSvMw53ik6HR7QiAf1dwiopHRTCoAjEP3yCQpn
52/pHpRL0YpZxaNbJH/DmeJFTBvQCTAc0lliFD8yU+pvy7ONaM8jz3P8pV95Jw50
tzMzsFOsvtqKkx+kf+/adGfi2or/WyXGBUfGk89UEiLV2MpIe+FWrAeb//YggGvI
T08IDMmRvz8lfwszfSmMAca4gX+zQfkukEHI2HBA7zNl3A8oKwrzoVSCOtsuzMqB
2Yjkcp7jDDLI0DiwRxIKjJu3N+M8R9YdF8li6ctjPDoeJN8h0XfjH+lW6ddQT3NJ
qZk4VO9PcToV5FygPj1BMtskSW5JxAxAXaV6iJUrkmDYiOlq0A+Pn2CDOYPbJOgG
Q+pNcfUPmmJ2Ze8xtnyLHgh/T6KEvlkIIoMNl+oXg/dyfBLn3NJt5pToKu4c3Jqd
KsidvJEjrn12DqAKb60e6lZkk+uh7yhQH5Bw1XlSYsDrLM1TX3nE2KqFczYvyy5p
OWY26v5KFBOhRFcp2jQS5AdhJmKzIuDMJMHzuhgVpQsUQfxbat7LFyT7tYfYstmg
7Y+VLWrXfnTvHCM6z6Q2Td8p/OldxPM9bTJntQNRm/0JkZdIj2DqwP4Uu1utzTlG
t161Lb77Fm5ayaBsGxjjDw12aaL8kjwVLxiqgxeL21i3zXTHPRWlsAhaTDSbxJ0Y
JFjlnUhknnPOw0DI86EygIIkOzFwfnVZmAc25H+QbB19J0HuCDHgrg5arGGPt4vC
FyXKgIlNwOFOkGBx+Ly0P4YSToqvKTVZxFdD9rx13cOTrMBkbIzLnh7ohDnxxfJc
RmiXEKOZDh+xyM/cNPG4ZFu4/ciz3bG8kGcXI7qU9J4WX8eP67FlnKVQbnljpNWM
45Xrmr3geQoCFpJG/iaKmAxK9srGkOFO2VnwAJqQYG4+jFnkAv1ShGid3uXEp6sk
aFYp789NI3Xyn9rYikXAckqNGfC3uaRHieLKup8uyatBI4ZTWPFX4+e13Kqacx3e
1jP9eMwS3qAtoDs7Cee17j86swjfrsE/yA6qgfii4qVcf95ikyUoirRa7zEn/IAP
ZqH1su+wLZ9lvIPAuApWPAIfdiJejAqQ9xhoGjauZi8F/KGB6//59BhircITydYr
t6oLHw/jZca57xEW3xOzU9VTGSc43PjOcKgKo4lBwW/+Yb9He3rR6zwNnG8llTDf
CsqMI55JuEznbTZmytaVJL+rbdndm5eJMGtAzjzpCv29yuDyYwQ6UtvWbQ2OMQ9D
JUIDJIN/GH+qZXTn1qIF5PsRSdhpXBjGrph/s02aH56P094U4q/H8P2yFFq39tzh
OiAgzSe7OKlSQo64xh49iN+iiYLUfhj213OyPZC9meJh63tMoYOYWfbq9lsB15kG
RsrYkBYL/eInjdUIRqE9oGaZvTOY65tOGLiz7AEmoIOn8qwP0DS06Gd20gtOFEuU
9UV0VT/WhYxJCchSrifWwDXelKjaga2bNJpMUGMVx56yc6CnjkjAF2m/NwY9Faq/
L0vt734qWzGSAZLGmCOMc3HWgQeCEmY7MPRkeOZ6MNVW9y5terkWNSB/IinEMNLK
jA+Ktd3K5Aghn1vNOrh5ddmbJnDVekmqyayfLm6n/azkv1f8EV7oNVlEPVQ4nqbI
5Bp3cEKgUDgfyEE5jk6bjIzxzIXpqFWFCfWQTTnZcS1MTwls2/vlFpVN6/Ll3W0F
ipH8fGpsSTK9uWcz+JFXtvWiwzQNcr/UCOSqCyH06yeJHDm+EM3Gi3HW5Li1JSC6
jCVb3J1n0BYn35Eq9laYqcFkrhce2NmkyN1MUwtYmnW6qIwS36W/Pnahl6bQ5EgN
cGPjYXZt2p8fqCUX7LpOMH4wUhLgMr6iFomqZdT30T3SOK3T9ddNTyI94OjvGATr
YrrXb6PY3PH93YS3qc3/e+jMiTLye668hKjXq1uPGu4QMkXsUNCN6bd8ssoErgh/
gNkYhGuzMUcqs0KSVypRpLBZqb2Xt5+YMJ76Uo78I+4ufM/X5A014IhNCDrXUL+y
ziDCrRvSC6exjMw6VONpoOGJVVBwN4eRTvAZT2bYqBR4HOmrNMj8Pn4QyWWwjs0B
fljO88j6K7mvy7OTAZePlI2UAgNNql2UArugZ5ogiPvfHmWdBlc1vnpk+OKn1mjL
F+gxLmgU7HFbpN1m3SFsTwm+vvjX7+ppeyrd/hX+y2O1dZcrVq5Qtv+1X+Z2qtxW
fF533Q/1NtjL0RG5ultonU87npQTJolQ934uyyEw3fI2LPK2IK6vO1ibmV2CeZqj
fx8Ra+XknRBBO+rKyAEIzdvIxAaP3u+97GrKfgo+bqn4ybV7MOq8Es3mQ+9GZ28k
r/6AMYEsOTa591QvDgwTt318LlJrMCrxH50dvmD4VnocaTW1vGG/hu0bZkJm3NcF
+1dVRzArua2ttn8EMBTLACJRjud2T451ZjNDnBsD3U2ZolU/K/AUE+P0zhHLWLJM
sXqFJqrDp4kaIp2ykVu6SrjQ0I9lyBtrSy8l5Q/5SrmoKoCV721R3h5TNnx0iZUR
vbTW/UZYMUXBDDnRlJxK9M1DlfmviS1c9UsvrAvwIS9OankYfDv6Z8PsZxGRt6q1
tpkBorOs6q7qYHn/ql8c5xVFFJRMapRT2i2TRyPpD6zUGlc6vHyDlHZigOEMJGB6
IBoWMMAs6cSMtOdMnAlYyRQ5/tfPpKVQqbFV1jj9bRQ++8wBKr03ufgRHpPEAejW
NxHrMizOEQzsQQ+eRSrSyRwY6NeGE7ZEFpRoBMZx2seQFMiemNhIztJX6DEZ1DY+
yXbXaVt5gztzxRDe7eOhVgMA2zyYH/MsS4yIJlndhqVC7/VAdYeq8coGMiP6ebfA
1fch6lGIBDTNvSIrPfzIRhZ4uXdNqp55n5IJu+Jf5q6DdRyYGgVK9r8svgkPQM/s
/oYaGllJZjTz9dp5YMOO8kQaZXEAK+y/rtj6nXl9n7gJNepXsbAI1Mbila9qMAxs
B9eeW61n1Zywoh9+P2TS+ndQWl+YwYjbTC8GXiE0F+FyXFcjF6s8s++LQFF07PT/
FPgJ/3YyEuvxINxX7pJKBnLA3jYw2n+rBsv1BESM91v7WdZUZ3oJ6qmpFFNAXuAM
KAwNaI/MCKdRTPvA8joD28EPlThR9Nk9tZTMD37i3QT615OeThwmjgH1Q1gb54XN
XlaICH90lIR2qp5ljoH+mWNTqpc/6d39ymAiqW0c5NNydn9FEu98J7AvuDHQpGwO
rP6VysyhoiovsubfBF+kmiyzOEGOvJSyoUo1ETL/FuInnxS8OqFSlPyEqN2r1H/p
gxtbCxshHAOD573rNQ40BBUETFN9yOiv4kldSP+Bu8mMROK7IqseP3BGxjG9dzLW
tNqLdG3F2Wzu6wAFZ/uPVVxAdH+HOq92PNP5JulcivGjuhbUeEkq9tPKcLmjDIwL
cIRaKRU14LQAmAK5Cmy7b/VOi98TqvpreIuM3eoabw+43TAO4lL78mduncGFZM5B
4LgR7XICt/oFom+NINEmn53lBj4vvHfZnqNpHn6xtmQ0oK42OeJXisGt2sUDALqL
1uX02UblXR6scGhTFd6WPeU8AgqCdnbMl+QaJKUG9z+5kw9OGJiSvfLgP9mh5ba7
R8HG+A/iB2RCTHoxxr/8GtSkKLY0ClRChuMH8HGG70WEbvQnOwfImEsZJ4Mf6Igg
+9fc662mqFdoi1ar2R35oVm+90LAPpPm6KPU1tuGDdCDIhoAskCnyVv8rvY6WLYt
cLh/+vB4CbXC+F9IaZTsmcIvA59gl36eX/s77+zbhVUC66gI8Z79NGy/xIGoJYD0
xS98K9PT8UpfKlttIL6lBEWaOVXpxVvG3EFpKnfw0b2ZBkOyeCa39JXSHI8uykVv
Uyo/2eqUGm4RjzHZKtQsQhjA65lO1zEAMX/Wirlf8y4EfXTiMbbWKaamIB4i+/W4
Kj8fpnDnKjoKy2aH2VvuHih0/9UI8vV+olWOOtv+dy9fPq50mlsdzjL4FYIvN6EK
+b8XagZorSJH9h4MvPqwHOyTC+9MU0N9wfqPv0nz8ewsyrKfysnTGeKIYhXFgMZo
isneZBxROO5/qIYQm/S7Kvb1cIQLbEwMmDIw71P1dJw8eP02tr8UMjOapCGN4cL/
7Ao9EX/Xw93qigH2Y4QXQq5rNRd9ST46yKHEJiQajFMMp9vELWHPio5E7Yiv3kDP
RjcSkxERwQqFXC1NFA1wx/bwiYBJEG1dbS6PaMjy/ldGQZ7DATuhMbK2EZBmPrJ7
s6V16OripbcDs/QWlOf8z8B2P3PhNkuXGL3tGKxPKPbTZBl2axOTmu3Nk9fuN3+K
gTfV4eiXtOofh7IGdL4eYR4YMqGNSwsDDO0hO3GMnsdk20PRSrXG62rXgczUxs2Q
UPNWwkPJAp+yw/gx+fXDuCxBAHFzwaLSwjbjCBN8fAdUBgOofuONeanSvy9UJibh
h3PvJ5lFfYAwxO6qrwp15WAjEeG6wwKcIH0W4QNFVYFAwpBF4PgPnULyTiBm5kwm
lCOgF0AZK6Z1BgQa340ltD07waeHApqMWN6S0n0kMEQwLuAo0hbueBkFQ6i5W/5m
SajzswUC8/8m7L3nqM9aTY7QythpjJs5Td+ofvEnO+rEyqQ4WiNOgZuqgKHw4vRJ
WW4o4AEEWGn/iXpMHc30cyRIGljGoNI6j3Rs2ptlJ9qGi4GAtj+saTynCEWTRRYA
4cmwr3a1ymw1hlI4IKwlwCkIi4+Lyrij2xT4sBt+cTKA9Y49Rs36j5DaGS3mLd5V
R3oscUTOr0EXOfT1cJdybpCBdCgzmmSkcVgJAEhX4KHQlTyUjT5QsUaujfBKljUU
y0e8HHnV3bOyEp0H56x7ajtqI4aMv+ixBkXPKGuFCcv9YHVLD1wAREU8ZtpNMS3S
PLA33Y7qgnSqwAVKO26cRVuq+y0IlvzePBtZBC3EkY2jQ1gL+zD/qr6N0XxsqGMb
pBmVsiz8P3KlmGuKCZTbK7QbNf5hosLvTNjJGzijulIslKCs3PKLXwZXgkUvtyiw
++6QVkM5v3X38qGmcIU7vUPfbyxnx11//VLJXqxn4oMnyLJ2i4Y1G4lretJGNMS+
b3cTFQBQjTbxZuRL/sX8zJGKgTzYAkgq7xHai6pstt66DtYkPHDM8LMLjtXGPoK0
FsrVbBbXCdR8l0rdY2zxa74PFR1Ux2p/kVyfVPrlr80sGWd5DM8d0OwjUwbKozk/
XueD+h36i8ier5/xEvE4i9VDPTCZpJW3ZcG5SIyE3j85SuZyQ9utQ5yGw7AXTqu7
tcqCc/OufHyH7UlzRDVBFrKF1L7zA6VGvsUKmQ5d6jPK59ulVgvuruDLH+eqkZ+v
N+HmAlDvzd8yjWFCEOoPUzsolantWaRS2BAZdrGatfmVW4Ox1DxOpArBYwEaLE1f
Sw/+EYGwgIYDAxqNnxKDFFyBhtfy0PAMMeIuu0DivXfj1z2Gc/MsHD6b0LrJDJuR
amTdH2iVAF3EFOgEfkPcYnsqheMlgUuAIFhrtB68eDm2A24v0xVompxtzKr+VV8D
HATbE/t37Tf6UOeAx8e1Nj6Blp6gxoB9W2yT8B7lhPfvqqe74y+5CfVA8nztZhUX
s5HKSSor2JUaYwtzUz0rHAmo3gzF8qaLdXUpQsyjAaSSLcfEa5UAhH4s/O9wv6xO
MpYttkdSh0/+UJOYgY5aJufM5dXqcUePLcetL5XF75jDoucMDzjsRBLXQ60J1Dzo
kolBeL6LGGLWXc1MesDFyFgmAujJ6bDeHEszZICgRsc8kCzFdjLnVKnXFFytNWIL
8bP0j/QsWqkiohkRvCSsBHAeGiN7Kk+LezU7phjAw3ywnMJ+Wo8j81bgRHq2r7PW
4XfyPXGN9RFFzBS+xDaR6gZIRfVwd9qY1AQRB5bPC0ggaM3fVdg9qhErAEH4JF8D
eO/6PgjTMA9t0JlChsDDWLVhOivQE+jd6801NxWqFFSD9dQObTpQSrsawHKScm1y
d/BchuIpyjt4NII0L3vu1Z02Lfk9LUWv8gK5ZuihG0lvMZBkA5NTJO4snQkJ9MC4
h0N8oTL45l2h3v/znnLYvPqjK5rNNVFyK9v15RXzFRqTZRowa9QmmRaiiVnUkQst
6AHkX0p1/cy6b6sGajeYoASM4loA6xCziwwQKW3sjgYujcsA3wLvRmczWcgbRVur
fEpS0doo7LkBQQeeBpcyqUErREKBl4Fs+dPWpnjpNvGAQLZgne/ElOMRLfx07Kzg
NApdoEGSUswkOZKWf0iAPstaPgCp9OXMP9MouBpjLJNIsZonIVZAGWGB5Mo++Hhr
POm1a2tBpFCRfqPdTbhs2UNs2RHIZzEJ/iEYiucuze2FShRbiKfBdRTaVdcQflti
CRxtzpyWuch+XCMbM6KXZLQiiV6bVkRY0AIqp11XfztS1SOsOI/4g43FeFHe+R3Q
fFojURIKHJi+6Vpew/g8UoEocVi9Om0CdBMwwjHr09yhPjsqWqS9jG8MHmmGazgz
9oUuqc6ifvnXLIdBkCm3yiK/VcNCdcLWVl6EW50gIxtJXABIpl0LNP9xLij2v4pd
yy9RIzB5Jg1vzC5DfHoKSnOyX2/s/Zp2H/CyqVNpzbYVeRXbZOvLGDsU5BdQbDmY
H/duIKtQNF2ybeBdKd5u0wp+Ref31YPQ5kazTyv8oFd3mA72g5S0ckBPcXc0AQ+3
zWou95DasKv/5G0FpayrcfT+tb+VUJJ+YicLNjf2jIOZOoyNa0F/1D27e3OGiiLz
XRgn3bb1S8EPAhmugrrV3g4B5kPmvlkJ9UvM5Du6YBWg8wJUs8Gie3sagT25jiMM
Ffz+1j7xs4BCCNjOxvG3Joa/Jc9K4hJG7bygKqLnybQD5b8GDHUfz4VRtGVnNnqH
XPJFrVJLu/Tq+GnTkrEo3KvtkaUNyR6aPj/IZvOXRSseQox1iiffJiyGWOtQ7TzY
RAHOU4n+Zly1ee5/vBGGKvGAZoEm0fKdXFptHdDpszVJk2izoxI2VDuG0ciQy2Uo
gTUceoN/x4ZTQRtMSh4O5AV/Ew6MwMdjxtZNKAy6qE9lq7mQq5pLlO3KMzSfjFeg
ih3136EKFQyOAoOCR4KSyV9d9tLlcasA+HNOLN7zJtUe5GTe+1Mk1E2nL19vyHVh
gkWQ2wgC11XCyiFZ4Vb9Uq9EGxg7hYpVHOb7NdtCWfKJliNMgRojsjvG1gu9lXuC
qJDMyuNw4Hb6jQVWSCar/0DoKTTzyG2iFoROV3dFXcY4NuoRGw8zzyndKqIC6lqZ
ZVdLwZLtNe1ebOJOGXwiWHwmpWHTbCuNXSd10bJlaf1CSPBJo+gK3WHNcdwM2JkH
xNCERgZa8DlGoRcwD0O5Y6IQLDG1OkmN+qigGNnLPH34XYDxz/rs+m52DbL/5HiD
5abvBSyMBiCiRK1Coyo+mlQf+7ZYFfn5Xp7NMnTF2XqW5EaYrhKvwyYfb2JhilFG
hUYtgNN/GfFLfoDdxJLyW3df1TtYKv3toJr+eVgRIkWlXNW4LzHg+nzTivSENpaA
7T4yvcmg87NPR5vkZiCjlsIP43JDLkRou8mmVB4uF2s9PTPD/aVXUBaS25qTkFYW
IUZYB4FIGLLRjwapCNkikLrKuKzbXMtV0h/zBrYvS17quFMzcagV4IFK+tBy3d19
4M+ciGvPMgGuGGJW/YGu+dBSy6rbyVn1UnSrGflquIEruFh2NIQTcaugCpaxmpkL
Ymbk8FRsAnjISBncKEVIQXkFuxCbB6yS3l9C1SpcPQaMUPLC5dwjLIFMyg90qCQF
063KiXQHrMXLnhXKY5Qn5RVfiP6Ej8il1nCP9JpmHle6REx/Mzlikzdk4D01DoGb
00dem2GLS52fGhU81FBDK15B6v2GGVldzIDEOoBE0Cw3nU9rY65JJS5+HKc1frc8
pLrMLmeo1slqtvhtjrgk0TF5hVQwzwe2zt/Izf+r8Oj6SYFESnzw110N+5uFKRbv
6tvTnY7nbJE1P1jUyjAY9nB9/B1Jwa1AMa3gOIXkEnHaXuQSxSYqrZanQqJbptm/
vY6HvOuims2pBJN7P3Gw0JRg4yXqrFqgg50sj8jRwu+1fdWAFY0Mkqr509RjfBHg
YEaQWWOqNNBCTnqaUJm86f8Pq4zoOkMToSHACqNyfJJ9gnERmx/IYCTFdpJOTZzl
5ykpmC5Hg7WIf4NMLUriXxEK8T/oJaoPJm8RkDn0Ei0cE7ViHgc+D5PYPxDb2fmO
5nQPNuTv81JcrfOI28QjMiBLnyNSoCwcjwvZckbX0mCkqWGjkVJDBLaUVJT5NYUE
UzPBaafTxxvpndhvz3+/9Iyh6euChGz5ekHXA1IHu5TZsdpuxLr4coOqtyiQrOhU
VJxl/nM5bcTqvD7rOovsMiX/0FNYQJXbxYPPHEVCtm6vsUlMdfsSbeJTXWO+sY6D
80RbP14/qTMlt6RaUYUQbePUu+jx5YbhxvlM/zTm4X7pR3qYehDpMNdDoxr8PiCs
vF649796vAGVIXU2v0U2XHYsOiqbucGoxE3AM2BxB44eWPNS93Nor5sIMvSPCfAR
EEwln1EimBFQuhaTb38P9wx25QU1/UVG5W3rabVyledh0x50XkYuBckBJVUuPkVJ
lTwWVLxClnyx0gWw5ZNH7a66GO0PZYMe+CgokPVKiqonC4KvLpjtPj5NS4WvKVRe
QMMVzBBmfp0Vmoz8wv6gO8Ndq9eo4Xs38R8+6DtcM+wr3U5jA0MmBCjZ0FkW/70Q
5PdkhtQa+pcwY0cb8miJDRc/HXjVJ8brGy/MHXjjLJ21YVY+c4otONgmiLmWfCFk
70IMSdmWd93Qjf5eq2ta6o3UtfrmT+k7BR3oAmbkfvDQ3/stz+VJhU+NcvZmRelt
mKb/wad/wopjCf3Mq3+sjwH35Etd9ENqENm3q+n0xg9wWIrZ3zIA33pY3p7Y9EYU
s0oqPtOLPKVYMxA9sPtJksxytnkrDVjUVQj3on8Z6JD2vPNO1t+Lx3A8zAj1f0JH
pzXFZ6786k6rNAfkc4PAo4+JRv+51NwpEEz7hSrnIP6ZgKbbXjlk0LmdFjd96vT4
kfvyeQK/che4GhCLu/eicZZaliCyD9+g6LiatzEMdn547SmB9A4gYGXEV9GYf8+s
GbKks/cKHZj0cmspSjOfteQoHjPr2/Adn4vu/RzasAwK/SEXcEml8ZGbs0lNmRTk
nF3/YYCaTkqpVLNBZ4TUhrVY+OHMwYlMzrKj7zGjt0izVmBvVKVqnm6VeCZEmQC+
bdyC/NOdRYQhuhLr7X+PylUNS0C7oA7j+FzxrHNnEDD+/QD5Qsrn9bNaT7YYPkqM
4o2QuTxocX8sgTR+JWXOi82cySo0RT0CCDRGLmGPzEJC9FOKHRnaqzvHzQr7/Bdn
QOcv0lW/6yaW3k5rRD4r1BOMteH96kTA1TDifc3DsozjcrHQCSZgT9BD5tY73ESY
qV/h/LuYXsfZ4FnTdslDAAKIonZyo+PXzFgL8a2o+BAzCPbKd5HS5yBQUSayMtnV
oQJ65viUTmTloH/vzo+bWqdnSJd0fBzmArcLwpS7sAFzApQel4SZ9GTAIFCKkkP9
jxccDG6nd3FHHFhf+ZKba/APoz5P6LRwxa41XdyV2XlNK2bgfKLgfKVExhdgWP8/
HCht1/ip4AEuMNmqlT6MdtF+jUO/0Tv7C20hh9JVElMifwtJswbyOgnsNTT77nJd
r090rlCPE+m6X7n9A5A+j6c3JHoxa59SLGOERJL1j0UlSZmRqgIVQNnKBJf/+SWg
ruWM7XGq8dP0L/7whftqbmj5q29VN1/8ORJ5WrKbzv48zb1AoSH8gynfUlxMikq2
IOtzlxxuoq9uO13KsNoTBfDvDuGyhuaz1i9fXk1wRrz3SLotqY4Ubh6NxCMoYhjM
XvUKWmLAEOhRutm9ETzF6IkZCWxM6aQ9aRxfvQ10Um5ufbVEw3FkBiB2OP7z1Hv8
TZNmDdztX1USeVoHJPkcse/Nfo4aAkBpXsOx/Dw6VfTscYtzG/97MKYgh9609iVT
caP9b/CoRdoixOnbrjNdocnzc6mN6sbXY5tH2B6Tpa9q9zq27QjHNiKlaTp+xB5L
9Nwny2GRy9j6wcWePuxeknMBT3e/iDToNfi/gRL7I+N2nZj9xUzh3Y57URdM+3Zc
oWtYiK/bwUYYfVlR45JyrdCE7atA5x3R7xs1m6AiEgoZVvziK8X6reriyPnSA72U
9zP3n8ZON6X0RYLEBOl4oibxA/WI+WE7q4HWkRAi2B4xYACzsu1M/mbf5e61dpdT
N2MKVUdIEj1jMsRarypHrjBOPhYAEkkgdT2XiixcwdC+Bw6GxTAjS7MTfjme7BRh
wN0SgoGt1T9y+nrUj1GN2Egb2bSGm8E6OXUgwRWyXFovs+Py4rnmdpdTrzFrDtcr
/JQ9WZh19Ri7kyrPggMENDMd7G2B0pT46J3fHMOprRCZqOaAnOLSrfCMUMBtOK73
EsfbG9Tw1YARm2pE93zuRK89F14+MLFeJNO58AAx8Zoe9IDwGC0OqUZTnMrsvZVs
WSI6zeHkHBSmTBpTQ9oX5U3f234xfsGHKmM3O6dG7Jcxl6yhDFJQG2/6jxXla2RI
Fj52fv+JGY+E2+zQu9vhpjHQ/x7Exo7wB11wft+AK5trUMnkOHYfwybPt5kMTPXV
l5DokvFC3TlLsETKCvdQnesD4aF2tj4m3H47rrMl5mQfYIIbUxGr/wCwmS29mxtL
XDLOruwuJyVmUWSLGSnt9CZrzoPNyv+iKgDSQuFVcDYVrV7iB7T3WXBgMpS6J/6Y
04DcMbHVbeitEL5cv9Pcpe9jI8PEQ8JYXwnTFro1aZECvhFLavS9T7krjElvsEef
fit8dz081Y+khYgE7ebVo/lLy7kqETvVkvmEKYa3zvTAcVogB29iIjnenw4DF+VH
Cz7MoCk66N+wrxhIV4Kn4rDj5KLUC5uYELDAPzikQ3RSppLiuYCwgO+v990GUPCE
7ecX47PfuxTpB3ZyLfOIz3TCdCXN1fVTK8XgopCzL3TXxhGzxYY82f5B739bSmZ2
qmHItAMkRSiQYJ6VIuHtrpuXu1apT69Ag3HDp38KvgT2dVeSTD+SC6OhNl/35C0N
kP+ahJzwFUJ8PAfdh8tLJ/9dv9tv19Dyczy+XI+ffertdBC8GWyVDVaeoTUUCihq
NRXAHXIF4pKtJbSNEILxtvjVXPp8mz1fzkQ4cWkvLAIYtdQheIK56aZw9So+frer
Z7GiXN5asg6CjviRUdX5CCZNQuxt2CCORs8pfWOJhPUnxyAHn25lbqB78djb8FNe
FoKr/Fn/4bdteU7mZrDSzVWmuywbeYzxaXB9UYT8Gi/N6W9nZy1masVbSMGxmB4U
LIHK6rQOkzLERfr3MCKIS28Twgf67l7DY5EoJYpTTvaxNAwrr3fDHM0/qdzyZrqw
6LaKNH4EY0qSjQyOBoGUFbqF122Fg4DucLGYtQu27zLzO3EYqGrVLbWvPjBh7RA1
G569JhwyTZqd4dyhKtkFI1bGFZUExn1dt4OqkBmcc4/cLCItjdbGwbge6havdkbL
zU5zUPrD/W5Rdwwx1oxIOcdIREjdo8m/r9FMXinrPxHJz4rOD4dN0ycCL0Pfwocd
eKPWZ9jVdXZ+jAuD6fJO6J21YKh7sk70QLLfRbb4yx/xf1pSeiGD1kMo3E4qhYSq
5tE1LkwUkHq6/wBlnLayA3dyak+XZ7YhjENDerrhK18nmzIXeOutgs09UQhgpGg1
dDC2YKqq/8K6Z2gTl/PfINLr+ZeHxFGhkh95JybCaIV/tnN1n5Eux1Qf9s0hJUzk
ExFRBVyV7C+Vsh4yUTQNjn7P4VlrYgjiBwTv/nHV9VXdKJU4sncL+RMsUigOpQyw
DKJyrYOHOP+BRI2eD/oWwhptb7T0gX1BYBMeZOpmdXoz1creyIqRNLeczAlAWCSY
lAefBbtLN+v6GLfFwLRtxAkEzF7drxthXUpwnI1/kYafJuzkUk7FgUfmMJF0a2KJ
Px8cyeomZLND8YH1ucVsey/MH5y73CpjBYTR/ahXyQd5Ioa0tz3u/eMkNOiKCqan
hxOqUydscc36eY0NSgUN9VlJpXRRXpb6AATW2Hys6KNyA6uvrm0gx4u6joRm3IoP
72Oa44aRsK9NDNnAgEaLz5Eo6y12DjACwOVWjdkJJitNd2hk4/qInm1xFUxHXS+g
QelcOxUmgI1+hu2fLkktfTDovsE9DOZWg1u5DRe41mXPescnXZHneRoxxODjThd6
CsIQK45jaMhYbvLqRexs0khbU8IwnaZxgXgRTkfaeQKyZqxcVcZjjtQJIj/1yhlT
Oi2PVrWxBkz15Wc/XNsyGS8yufRsVVL0vtOmlYcsqwM38wvgQ6SR7rFNG7uAV7Gz
Ywyp0bu96OIIqjHoNlaKF8XH4VEAd0dScoXj0uL69IHaRooAD0rWnJ+A1G6ouSF0
Jcvph8tvBscpTJKLoeZCZlxTzTVNtUz/fNMLm6fEI2fOgkvpNE0A0puQ7ImlNp4L
eZICq7JhieEBUwztY3XS4lho0wuxQl8PEWrDQ2MS/To4uP6eCpblpSpymetbuomn
Vp0P604M9OqBK486iWNnk32QWC7xlFmXCnEcBppZXtIMkIsV0l8HxbbaxNdpAHDb
TN2TAySZZCF9MV+HRRpNlItd/PhowtOpBrs8a/Iwtq5Pum8ifLrffUTnfmWebXzI
J3HmCoRJdjlIIwFqbLWeijxOskxI6dYGJ1wjdE0HC8Nc1HhYWVfA06zQ+7ssup0G
s+1TNRORna6/rJ9mKO4o3KVEfUTX8JNj6pNllYWz19LxuOyjMrj+W1X6nlGNVNgG
15x1PzPzOKrrvwSR/Bh/RHaWVnFZnsdoUbHs9bxGOmbkDYBJlv5K1+RvKTeXrFVS
srRCN3q4Y4yLvUHJHwKYlk2O+wgOvU1F+xZ+Z2LjlnzxGouU7AaLu9PZv5OeVkLT
+Y0DtHLyMu5m0HLq5tKJHaLOIPBNRwJLIfDeszifHmAan2PcfsAelsDYsWwpe4PI
y+kmALMCAXS4YVNx55XBw8zcn6s+MpmTsqhr6px24E8vkOyJdIn9NX1oix6ROaXK
9um+7q/oU+u9nh6I62sDCl4KcHhFbxxKSmBOuLUk55CQ+lYYQuiIFfv3Dw0d7UnK
CvrFjmDBYhM1qwkbnnxLqytu+pQIHX1BS1R4M4fBTQrmumdLcYUY039rL+Z6cvCJ
ZHN7SdYrceQjoYKYdmvzpZIUbEnFXZ/4683RWQ17cAfLrm4GbnWdc2ZryMbxaZo1
7U8wLIprpiFEb0/W5HlTnFHazbUfXAXjkufWYzKi7879eZSTIpG8S9fnNxEDRnFf
1MykWVa+q9ne1dw7qt1h+qyeg2/xUGETsywoZQsJwEbfbmLIxTAYhGdJEKRi0AGb
YjXXrcqo0rHjaFxauB7hH8pooDTDAVEU7ZYZAPD8E2Rfm9CCZey6QxVFzw5cDh9j
ID39LmevlskQy1PJKQg7D0w2I8LxRSHqbHMrRMwt0FdtjsVIRw2ZExehR23/+d6D
R+g+Qc6UHTBGxpEHD61ALRgubdoSvUVNu1bi2XDZTwIiL1SIFiuBRwFQiVk/31Vh
nR386l+NkAkkbr2dkk16D1CQdJG7MinFJoqV6bOGDhyvHD8q09gWaLPXmCvcBCsk
q95aBHPqjH1cO0zPR19EcZ0DyjZ1TXBsjGHdvDRshBT5wjXslTzrOyZWpu1QQTCi
PtOtFizz5X/0RBOm8gWgYxx2Ra8v1U0GnPp1tMcCh+8gPOBYxJd/H3Ou7pak9zEv
bI3+JEWJkwp+JXFKEyqdNewpFbCTuK5hGCo9eD71Gs17pX3BZYPclMVEoJ9Hlf1W
lZfwyo16fLymuz874dAp9lU+YrFnBRQapasxHOCo4ksd78dK/uppIPh9v2Ojh5gB
7t8HE1K0Gh3Yzlrbj9/ibRy+qN4sEB5JDdbAoALpWIcYw2HMvc/w67ssj8mV9qXh
xsyShBRxXuJvhGBJndGi9o7TUJrY9eYgV20/ANPXI/7U/v/7+0H+qZCavJ4umzkR
8au4qDhTaZjxyi4JX+OPSFnZTq2/sOyMIwdgdYyTxmgjH1EoDwhwTWe1e6cmpwGx
kCbgq4rZs1dY7uykbEKeGIHRHjwiUG96qw57T0drnpkAjkHexjQpsH/InYsKTtJd
z3SftKlNE8067qTwGUu9eDB0wOVjc7XR7iJFRTohVM8zoOkRKx+WQFu8FbrVz8Sp
lQfrfQoqOpBBpyIdGHPKH2TYf/gLcb5XT6LASBtpdDjpN3TOqIxBCbjB9lF8fUsw
RXDG84stD2eSQKQq1NtOuC8criBr/rKfBDpOs2dLLFHwoSmZ0mvUXdPpJz9cKqxI
0ik81AN1uvrTWrkzlY0j6MSxvKI4KOI1D2qSZrcpCsBbcPa1Ed+hFZ8V7BXfXfP1
F7lIcuUbVCku4OlL14ZNKqgOVCdkHnk2guzJpL2jXGL0ELeQtswvjcLxshnC0R4B
R2O6gQ1oDDC1O2mAnFRukfHyzL6koeB2X2vZkRXdUI858VevjbaLmlVhtypB/n7N
+iegZ0KmgItKJGyIaKYH8vK9FfkO1Pc+2BKpYZWKPOJkdeDWIvRuViZFHMiLkeJM
h00Bt+WICWepTn9u17yZOfcSVK2nWcCl5Qf9BIqLvAxy+7TUXUubrq5j/yTv9OdK
97OGfurZMyJzJfIScv2WIkMV/kEz5cblRRTdl5pdJB6to2h2E3ZtjCmA9DNEn2wx
v7TZMjkgav3OGem5lRkpLsrmfcl7A/55wmrYHzeTt6ZNaAsyB7sQioh6Yf/x/E8d
DGJ9hwFSVSK/hOg4VxZlR3GzK0tnJo3VwpDubHFZUfDu9kyBSeB+bU7Sh48xzv88
+Ntj2IeMgHG5dbUHg4OakiOSzEYsN7cEqh9PnnuYPovrOlu9deb/STE8fu6/f4Pp
myZc0DJGdze/sQ6sDN4ps3JZbtRC9m7HG2JjwYbkwt+ZQ5e4G+0QzeIEJTczOJa6
qCeT9DnbQOSRiWSmrcclTkWPH9ruiM90XlRoBXA3wWzqk7se6QS/iTWKgHtfasx9
blyNwKQ4OqbrKhSNj67WEwOLzQ5sZ4vZhBEEhdEpIKvOf9MR9hJ8UD0kwxrHMamC
1iPwnT/ec8OSZmWx2wYZgfpX0FUnf6M2YeNkSOLcK89f74JCN9TumAybAjaAA8+O
3miL5a03zfzIy6OAq5lLVnPWaVFRfYGYRN3zapYjsrcKdcOAuTWP07OFyJWOwlBT
pMeB+3z/8NPgSGqHe4j41sn+sDLpDziGpRTcOwLpjACgs9gvFft2YzPge4Ec7Uen
a6uLwDIHKMVKt5SDT2O/KHK4qKMF+Esxkj/PXufpeJH94nvLEpGReTFVeJSVAYmY
dNnJF71QyN827TzrgxoWg9DhmVYPWef3AmCP8lf+S+UN/iCT1V+Lfw9WGus62Q3A
42c/YZKQmZIPDtvzKSnsxfyRzVrSbPgFIKqqITc6PBU9xFlo/kUXGn8J94SFuuTO
htApay0N2qQStnW9+vNEYsgeNrvQdZuWq7nbW8tYupl/7xGEi5zLAVJlSytQ9EBH
PxkYiDBCbB52MitWhADp47OvmV1bi9U2Myr2DPgMJB9JbgLAtObPijyCCWV+FpwO
cy97QtRZqPPCKh9h0K09l/ROnAutJSqnQsH9/NT3eSW1lfekJeVeYukPwecqry78
NZHJTilomvPty0QSx79AFwUXjkF9yJ5NmUSqtPLbzzL2DjqTc98xLvverShRA+U8
L3vLTcnG4fEtrrnVpsPmKeh04gmZIzOgujmQ+22CjEwfSTVI9cEz66luHuJkh3NV
DeXYJsxylG8iT6kTza+U9uoogiJbZPV1KyIGGghOO/Zo29GeCUS/UuoWiFCi2HQ5
AEgkw9UpKzCMAKx4HcNaLyAPJppgbvyQl8H52ygG9P95K1S46DwmCLa8ohrK2T7M
yCzuAD1tk0s7hYFm1/EYTTHGuXfIVPfTvkdxy/nsp+vCkhcWSGE6p95CvPN0ks4o
nrGRvloS7x2T8lzw3pQw3XBR7cPnmnRxM1eOhRK/BpVQaWMh8Byj8V0DkUJO85bB
Pu89yv8/daQUZov34ae+wkqMsujwLRvnI2FI6NaTc/0yVbMN4R669gDQRGNf1P7S
9hhIXZcBe6O15iHo8vH/+APhgaTf9iA5Ohvz41b2mNu+LQjquA5f6P0uvv87IXYW
M9ZgTfICDDLKNdoVwsr9Z1kROC+HdvzN6C8NocJdsE8TMdzIjOoZNX4bfXjFKOV3
aa7HjP4qWP9HsoEsMTZb37U1Tg/wI5NNHslA1MTt4UUrYkM0tSzcFxnDF9OYSjM1
7pIeSKr5vayIK5/qAzEmc4EAkRMUyG/BBxkR8v+r++ymCxAu9VLffPOrstmVcjWa
SV/UzsXKoLRTouoF20m7OqbrOXx+I7+411VRQZLamdSaQ38HNlgiQ1Sgz+GkUUVG
CKW53wjK0LU7RtxYp9YyE5X2D2OHMyPpCBr9MBrvu3Yq4w5QWsonhrmvdolSvKpZ
QEY70DvgFcHmvFJdo3xZm48pcaCOX+OrGtri1ErDlHBu7iQXUjw0GlWg/WISqQof
mlNpjzy0kjgShYWeRxu7KJ52riLd9LkN3y9b2pTaPYKbcLnAOi9yI9bS5f8VaZcv
sKa0W9wW0u4xiLRdQwbRnpKmijVd3M01s+cpCjM14F6vHYh/gm08DHyI86214T1V
zduiqGe5Wl5lN5mvwA2NXZ0fm813QL8u9VF8VlV4UzvhA1LkBaQv6b6ximrxyymQ
izHZT8hp/H5UNi/Mq4mBPguU6lpPXizeCyLYnGqX1gQfDyGY/LylsXM1AauP30ln
q7904yAzyN8RoVWhOyMrKt9JywJB2br1CM2NxRlUhxSjgdxC+f86FxUwUx5BJmfD
m4rtUxKLcgQzCRNQX96tlACKUlEPmXnNsktGoi4UEiKOGSoVizhb5g7/23Bdhn6v
wopKM0vwMHem/NTtSl1aHSikLNtj1grQwc2AEqyRu7kgzeia67YdFirawoJR1V3A
uJVBHRJfhGxWIaHUxP5Dn5crTUc4Vl4GFfjDbds7mNMS27+Sl00MR6TmeSmcb2ux
VL7bKPuwzQXp9vovhsmxot19in19AO44l2GEXh03X9j/84OMefppTRpdnGLfcmCO
Cz4W7pVazvCTFrOBlf+FUxFbvg83K+W4JAYIUdJx773bJYwoCZKNmg+NQXPF2csB
kj0n3/BAVhj3WL63ETzVatUGCzybpbYTWjfAgsxoelj7XfLH7N7JovQac5NQIGEx
CmO3LIiBnxgyR/gZdyHbNmD5iyylCxbzRFagqfGNK2aOBny0ylQurk1lq+ZSNPol
XkJAVpntWt4VcugXJ3V50mN8KmqHkogsCsMwHKgwkQBcWW2mV9OBRu3widaA6p28
ZkA6ASeviSx7Z60EsO16b5cp6d5zi30HMVZUqS2tXtqXEa8MBoV8uJWJelT4QOo1
PWTuYh6yMmc3O36aVVM+NP3IITVEFZGP4ddTTqQDLiNPYaMrECHp9Ui13oGhTO+y
OaEgRoj6v4zbcSjRw3WoMAAOsZXn1Ra8Y3NBDcm3VgmpBWE5GTCQ6WrJqCTHmh4Q
8Y9yFn3E2B7iQ28i3Ehm8Mqr+w6BG9G3ol5ilIgDjOd+PPimbG3YGzDK+hoE8lWt
zYLkXjoWhNoZWIzr0thZj3F+7EsqoUnuwnalqKqWQW7M/yk0MdwD3a3XmnbTNK61
jcZQqWYAMrA0vYbUc7pp+36yzvcXqjUeQF4fYq/h/7QjxAKKooqp2cZrSWSQxbkX
wXOSlLt4trZjk3Oi8Zc90VuYxYlh24u2Dtju/fST0pQaNsbh7gT/9AnKdEZxCslD
96dVlBTSvXXBBVUy1+nSf4gXLjsB9zboPMrW2RGy/ZR068I/mpJuvZvtBnA+Go/y
dbaMhQGf+bTg7Q2H619CYcpFF437hQpz32ZUJUcGBd1VNYOu9HWeonKeeTEGzMSJ
N04kgtAjy+PK/42AyvOU/dew517Vf0yMoKxneluPfWQ+0BTHok/2GjvcpuHGBP3I
mEK32SiwVRsSE4FlFjQsWB6jHnSv4PPdF1Ew/AOaaKjbm8JKoyUbfvHVBemPq3i3
1KFO1YVPJ/gzB/uWBE+n05UqUNcgWjF8m0W2JMMYwj5lVtmPk5oDOVnLMFax1onX
o4YzI+piAh6kgKdTK8Tk0LfwJVUE2OZCJZ5Phuu5kE4Q+9TXuxboyklDc7OuAuLi
4xqEJhNE4Qo4BgpDF7Ogu1LJi4JrYmY/JUIGx2rn2O/ifAj9yU88wz4IzKwyFOvE
e4UGZYo41T4GiZkAWShz2hQLkimxkZr0rkGP7VY4ALRfl7IpxVGO8oJLHVpX2NA3
xmREqYOVdX3+k8fWlZlHLEv/IyMfGImS16rDEIEAMWzyGCHawGUv55/szo+rlq6a
M0259i0qXWXtg6VvzFDaqVZ6iNCGxdDMMSbjIC4jFJPtzKaKFm5ZNnnA7yshzJSf
zsOI9Y7z/jyau2A+LszTfh0lUdJyI2TxmZi0NBKuLslCPPeD+Q2Du1CCcLKn8eeK
LFwfL5WVmMkusPej9098EmEhD3l0oZwj8MX+34qCYwFx1gDR+mHh+UVW+rFUtrjU
9TpPAu68pg+2CwCYsPXkOQkfg9F86gNIGe303gGqyewcgjxy09O9iE1thvtT0+Gz
J6Tf37BKuK9k/XBz+j1ZeN768CygXzhtH11j7sMGmdSjBPG3rEPm6iMPHYhTVEdR
PvQruKD3y/f7fBuAlYwM1wnvORPqYf8A8GEITUw+sOB91/THh8Gl4kYDdcyLmsef
1tsdsQib2L5YhpNDSmE8zHg+oBv2KMVcrnp012Y615KKu2reoNzLEBQDSzqDxmOn
x4e0X9Y8qDQiCqMqjsQr/m0rD0Wtu1itKg2swzvJc2Vag1/qLMiiqtUHWh5hz1Ps
VFvoD8T0I0rlzqQLmSlf8UAHigzUt11lLWHcG93Y7w8ddYtzcDwvghu01gC+d6O0
ZJgH1qDNRdJ/NU8g3iscXyFieDAAj+PgXIxjCIz0hPMJEpK7EfwAKDDk2VRHLXU3
Iylfi+QcoNG8v/tuQktHa6ZxUlTYB813iESTioFvwu6blegeIem9LbKigNmA7pRz
R/y7EJwAHndm/ZdtLjOjJNpYnSlTtwmurwIm0YYmUy3hUQcE8rUOJ+c/5PO4vKXe
VZEquyoKt671AuWzOo3T3yU+rzyPxRZ25br7NrEbhVQEEiIO+0S2WrIUxUP3pU7Z
VTsp/ixI6F/qIKId5lS4v6N67HRl2Tc+sNsaUG+gF3OarQCU7lIGkTWuF9xmHvFD
3Zho+r08UzOhxvAB7FacGOMIPAxXehM7qHvkqdqdL6DwxboywVP0t/uJWQ1eF9pZ
4x1mVTaRCl84A7Tbc9omzkB/1M/4u6Otg4K6/MHsB1OJA5rgJUxTBan6sW8N1yij
t1CGCTfZnUH9dFNLSv76Kxa8AwG2G+rEEcpX5wjHWnlOAI0c6S+TL7Ba3as6+tWX
MENF9hR+Vnr/b7kgsbfuOIKkz6mj2f9pq+sg/b3bUkiK+s09IPc6Wfqd7T8/Wqd3
qwc3WnF88w6HW7FNaQvW7AjvUrtXo9KVE2hZAevm9DGdSwDTzuLKMiEYO3ZYYCm+
ku/VKicqRyZRvfqyCb7B2tdT/+5bOJDwFh/IW3RA3v/vCKEbTpm1hPby7/Xdny/S
vgHp67g4MQGnf0Ct2WKIH4VSTCp4r/8wcMBZ4rrYyn5JX2kMV1z2u6jCTdEJIo5O
vIlDq2BCrM7sATSgi3Q7JfnksqMu5uoqOVXv42JXhXEgVY9vNmxjyKt4ySQR2mWC
ShP5gRghWbABbq0y9nL+Jhqvx8B8FYzXsHFoengrDakjZ1iLTmsVdZEkWsMhsu1Z
Osem2xpMcVMUdmMpofHO58Zwln6YkbMDp6I4fByvPQndKEbayYq8XdRgc+VxPe79
yHlYayfCeXOzCz34U5ooDTaGTnPLIxKv8A9IRHMRbGXgwT56jSJyhTtj9HTQC8B/
OW5d+7urqyemHnNPClWZfA3SAGThNUsigu9tKRE42JYOi1n4voiX8GmRmUudfv17
KjJvxM6YuMpPVqBDAIfJhHOkVYA41BPtFFUX/QYRffPzNvGOV/Td/IDCxwyqbznO
n9hh98yKazu4xQqPVnBb/FJyb8qRHLpFOz9y8mi8Ey7tJd4YGYWmQrQ44yhCqdZz
6aIcvNu5AcL+M0bpSNYfzwayv+Og2LaMESxa0px+sQTIIthdOx99fK9YG2Sy4z1a
YMOyMg7RZxK2mT6ekhWhUfrCSs0X7rAiqmAqO/Lzp3EUKCvBkh/RXZdMVkGDTeBG
rDTqptiXA9o8t1bYWFjqn/7NCK7k2uhlm9SEn10k8hAr6xha7leZurAbx+D7nDqR
I7cwyZjcUoSGp3FgJoAXWyCibwQCPdY1ponmNktA/8ABQ4p5AL3+DUqoaClJWXev
Z1fxlg8wTIMiEGdjpqaJXeLtweP0JFPHHajoZbR/gwGuYsca8S7NqtBqMnGvIgbD
kcDLgdxTWS+bnQQgKopiskX43qCHT94ZkxzZtdAfZn7qdTga/mlZ2fLY7XpsxR/H
vgRiLGVZpb0jr3UJYWeKhZls+VRHrNpNUoCtoqti8QYC53wtBJEL+b5vWVG2lt9M
T+rGhPjppoS+PrFFmL30O1NO8yNaX4EpY0d557U8+mhMRMM9p7h6Kgh1HyJYo9GN
+HXU/8dhj9iqjitmMxW4e0A43fOlqx5M4pYEj1WC73VAVHy026BrBknlSYagjMbx
5MNKKlny411OvSGOdn8AEfj0Ku16edFtNvHM1KRq/GyGt3PEWnMWWrvp3XL/2gZh
uH9v0QfK29D8+glqmcbqzQPyH/27JRC+CNS2NIXozoBuhSwIdovjuTm0B3I+ofvf
A1Tw6ZMfdJL24m4w89MMxnZeNh/qozrAGDbCQoHIWUNXs1aOKp1WpODgcdN8MuJI
tHpYRTuKSiqSU09VRCciUqfGNjmMEoNIOzRAcJs7/hjVHH00tt7+xMVHCc3qzcEt
IAhSzCxxqfDd/zvPCtZJRmC2yz85YRBB/YiRoYJkwQbe//oTQ1o/5X74ErCtee3Y
/oSlXPoNkZ9eZGT6pa9xl/yF/jmBk5U0xBFOWGIhG4xmkGtHktaVqd/yuoS6PfYU
DGXLXfLiHPcFXJMxg4akea8sA9rxNC+3pnA2stjxARW4mGBug6Eoh1c8Z+1WMeyA
alA5tj2yLVMTTHsaDNpfjSMGaLG6buA8Bsg0uUbkEBIClEXkJRdKt/0Uh74Immn2
3TxotYopBjWJ9Jr7Tyq1PQ5tJJQ1BFmEvmWIrXjIv+l8Eb8KHP+CjGBEbS7Bhd08
BXHIO1HS8RRsLUPO7xFgVTe83o7IjpnBFsq4mxj6fJv8+L/xw9QnHm0Qlm8paPMl
hYHmed0Biu9p2MuYxhNA0OiNAaajcvV8EH7wMBXjzsoWoRs3KRrZ5LgZAhaZaEJx
h9hAODtqDJ6D8eXfbrzqUk/oFOQ6fzXanc7x663AVSMzRqr059iv33bzLKr1Zu1q
bBKmz6ICkU5wSs6vvRHx6rMhvTeE26biXkzYILfsUXO8ZETtEfrNmnkbb/Axsb9I
gnjy7Rne022gV8z0YYJurt5To4rwD2i6hLtigFC60jt/48oZSRJZrDvI8OjVV8gM
iLx0b+rTk6glLRQ2YDAzQidV5xhLdd11wQ4f3WjdKGKH+9EO7wrW56wDH0l0LVRX
uWgTdQUUl6sgfwH0KrAn+HYFD0AwzogSUZdwmnvGkWjrM96+yRI46yPVzeS8cqaV
zA4BgO5upnU5/SkYX8r3MyG08IbF56pqM+ER7kc1wLdBqtpM+R8uDlqlvBV9ouoV
NchmftUXvjay85QVEu/NbgIKxyC5pkXWbDfFBm/Lt5XiNFTSGglQ4OUSHVSshlf6
tvTpQVeZRFo0dusivxuuz//H3N4FxDF9Fu3TOkNTMss8Pnx8ILTecpV1xA0S/J4p
0y9tV1jch5iA/mkC6RO9TkLDbh1kTbzEMI7nT2HsZcmjq/9Y3U8TKyRp7rcydPxO
ZycKsLdEk2IE0Q/Ug2AkXhYxoN6jBm3M2BHz1u33blBPBcWsQ4L8u1jDYZo6WxzI
8NMxRS0KlkQQPHHy0aJBM+Kk2+w9ka8Hy2X4pn/IKu88RLsY4nX6Y9WecVolzqcr
WkGBMHdV4gEtO939omY+YA3+i+4diJHTBng/sKFOx455MfFCJ4MIfHiKNPTSifWc
mBApYO0TepyV0tXEjkOdIUm09lBHXGaWCMjwEIlcbOoanfcMxostkEYMNDA0JpLp
JZ4oM2GycP2425VHXA8GTqur0lO597CkXRwlJUQwn9FVQMOU/R72nnivJnVVDh1+
w1Yl7RllEFTq1cNNMY+bXNqAAt0yrZByTFWWVZxUUn2a04pwCc3j13KBmAm25ATC
4Ko4vzdYZGTrcvXNP6Yin+uUm0+Hkg1Ei/jq5C/OCPPjU9D/c6sfSTM36ryYOkKJ
HX7tydgrP5pZVPZn7RmamDuxQP36rztYsS4yQEsKaMIuYGKl7/Edcn9WgWnMn60Z
8EDFRC9KrBgPh0nG8tnh/YXOJQ006CzbVgpVd+osvizTCFimfLwSOTi/+8A2zCQf
fdkWUElOPChiSjsEWfPr3iwrqRci/Iu/vaEQF88o0z7eaJJvhWSoUbrNdCK+RdRI
H0IlCXhhbIa5B7ckRBGWcCravZyjvhRt6vBacFjXb0n3DlX8kKr0N4Y+VKkZ9Wwx
b39dBpeXFzorMO3KgcJfeWBfBiG75FlyjJiI6Ts3lxfIhFIqXjeLDhGfCO2iDGZb
1zTRZPYUTnoqN4/ygJl+pRZCf4FBmwsseQmFtEoYkNyXgijTBSTD69405SkqEHwz
XtZmuSeVbCNg1UcmMJSDoqH46MVdO5BQS1VO1gqA32JJw/Yv67d3DHVtP4mzAfn2
2YZg4tGXyLLus5FKK8rXH745Baok2xT4nTvMI2qBfTbINhb4lvhQpK4HHsSTPAcE
BZY6C3eKZhDjs7ju+6rifzLBuLQzD1XXjg7F+WQHHETZ/bSd39TnJKBl9b8x76c8
KVV4zQqGZMPU5hYYYOvf3LHn1KCpFEfpdDcHibGymNk5fgn7mApo+Ta3+kN+MIET
REOWS2WSjITUea2T5cNKVwic9PStDKo5j3TcDfaPKXsuv1d8dJgMrrXra530mrTj
TAq/2DK/uzCiCP0kxB/GcSlmSbO1zkvzYHd1DMhSgIYxErlcA7vSRIjfANEKbZtl
ncJ4RSMEamv4vMQNePpT73cCykK8GW80bei+FjjY9fEVW+DZxTDf9LjSetSh0Jm8
NjxMj1RrCFjhiSVTKEtLrCdBK3Ct20yggTpNQftdNDkh3Lf2FD3a6SFN1lbz6NP4
vTmxGMMhW5sDgfZvCXjk+vjKY99y3A1t4UGGMOD8dN8hDg1fcreiSxudGY/odIK6
Hlq562u45y/gIpI/AzcRnlLLyABYWweAQ+aDi4kXXF5U+cp4HZ8OnunTWhrloYrG
U4EkbiGuXN+tcR1GMRYSvK0qJ4BTzzwSwJu8ncOYBcw2FtI1y83ZCK/p/VA1VUDV
taG7Sbr+M9L6vpBmvlxDxxBbViWDN1U/jhmLYAYOdT+zu/0XNpOPa7ogtcvT98H3
Zv6SxuG2SLibjModD2lFI/rbLmhhoVEhajmK1dMEVXEuJRXZlwYT5Z/OR47S388e
GUP7M1TjZ6I/qjFpUAcTYyiT8yx62kZcXB3zFap1V/mdtMrte7HGEr40qW3iDR1g
y5KYyqKiHMFAwpzbT3UCgXBGwVMr8A76Yizl5F4cqpCu/RiSBpaAh6kj1kmch0nP
hsuNuBoDRgg2PYl62x+kjBK/o1p08o9KOrydceLZgO05ffSvWb9F4yVmmiXHcCx4
ClLfk+xxdesNtleL9KXTZxkrFRb8QckcB3bUt6PIIBirNkuBJFGE8nZNHkms9/fw
L2MzyjdldMTwj0tGxQbGiG9UN7kHwEvWe6sdDsDLETCSrOS8shMBDMJGyiZH5sYg
GkuT2Tp2ulEcXB/1zjvDk4zmUd3G/jGgv8j4X4NvPXclW0XNRLFuWKTQLejS55D+
Mue694GhO5n1A4WkRU7fidmjkSxbrafBK+4VWHbO7a3DFVSaCCn3HiVRniYiA9+0
EgD6xxSTJJYJ4Dw7sjlTsnr1iVBAVLeVbxevs07vj/3rQQa+44VfuF6/RiL2qTTX
2JpvtLp4AhycvUMaxuUAAY7WSJ4ZqNF59xGWyO16Zq64QxKlxWC5JRW3LA3ixX3j
HEWMScX57GKJFFYcrlfdR/B+gGG8wz55lpM0CsaO7J2PJW9e8x67fmY0WAY2x94c
asoiOZRyiTtgd6kKXLFZbvmDs9rm5P/TS4fkG9ybVioveLSNtRgNEI8Ab+dnRaci
+OJyqAApJgaRSCZeddBYoXsVukk5qmO9ISX8aswT2JThzAO6Y8no2sk11eii2f95
KSun6U79QzeJ7RwlfNJCAVG0YpxYnqQsdJ04fVsiMRe5liVAYjd/kANvYPZTa6p/
XHey5LP3TcJD1fsjIQ/JtH4wVDaPtkW8cq4d48V7QsNGoBHuboSdeGhg/Pz97XTV
AazX0sgo57B3iijJbUxtuSlucFiX6jB0iwKPXb+Lvd0JVuFAyCwKzNII9Vpwwi/o
xbxZHRUNskcE9yBn+tJjGCw8k4k6cFpPMSJP+IDOHuibS0Z38/Ftb/Cz2Pa7DQI2
/f82S4q3OpMXm+qJzYeuiQ7NeS/QUD90YSCgjpfxjWZj60V4FVs3zRIA0+TAsaC5
x9fgD6p3jJC7+sFly4JfHw56JfLALNHm85cp4mikDLTx3ZSZL/5VNc+L9s1cEgXe
wjb8Lcpx8dr4jaQTpntJVh6Olk/lky+eeXqdBWMdURnYXb+HwNMlKalT1u7OzV4M
sjrBiI27mO+Qd/MbvwNa22S8YSozuPFs7395mC8x1XtHrmGH2dwhiyDoYbXXM6zk
u/33WXjQttFUwdskacsxvFFfVKKj+iW2FXvsatVDxzQjHAX1iDU4qHKUsQ6627UG
Jexw02O2cZLOr/uE8QoYOv1/MZD3F3oWWUZp2zpjwOrac/7oVt1ayA/aAvU9jR9c
f0rXvBsP577yAIl82Lzvwk1fKtnNhHvX3JZoYFqLlD8MteW7HkJIxvrW1HcL3A70
ZuSj8gPCDTSoF3NtdWHf6eaTdDFhsYo0VCH+I1oFfQOu7cVnlp6FpbT5ms7pozZD
f6RjMeKW90jcSCYutV29tov7HgTViXGpSY5vcMYCccKYX/Vl/KJfVJOn2ITcEpZt
n4jZ8gccwAYYbBwxCvWy+UV9Nrw+kvhvyXekS3WPUAQfFF7nbI/1k1stEN7pNxz2
wwA4MYm0TS2m6GOYVnFsMJZnM8H1NsuYtuaaYNmgeVq0asRRvMjSRtcg+BEBGTBP
Uea4uBRHbY15l9Nt/c4P6tdl0dOoBADt+aRdVfhz0aGON5C3uPkYDWgZn+YK8VYa
Q2svSVRYLGKpU6nkNwUoSrD60jizgYUM64eaE4pWlJOqyf3v2J6s3q0TDOe8Z9Hj
gCz4xLTdGMoIGwCtgHUyFFuK1sDdytBv7qyp5xRfL5VxukQtBictdhQTGZHMNQJ/
8Vf+s3uEkmN8Kan5U80bMbV+ehIVn2yXQ65YS6yOSLh2hndzmh0PNlUKCSYnyK6a
FHB6tIYxgx+bjGRZxaPKcVS8lsEYzjjHiABPpTtHLPEvaViU7vap8SvITGhSsA9G
fyTjpg6IN04di+fMvCKw36ndjOxQWHaKfEl70JMvdbOl+L7fDGSAJhOdhKaLXFXH
KpgaASVQNV6JhOFkA/3+TkHLFSBqGZqMXywz1IhRyjIYsZA5KcRxW7bO/vprFhow
WSQ0aAj61o8Dw8PweqD/pemGosp8QsRZCEof4kPierJaBy7vHlilSLDtdNWg0WXj
cDyT6Wghl1Tg0laQEOU0ierDFGLKWW6pTnxl1FjgxX9WeBiSMv5rjYVTWh2VTV/v
U4pftwa9OY1/vecaCGPkLd4IFiqouy6GBdI4ssefx7E1AeuB8lymzNzx2tFSJ21j
2UR9TskY7Xc+PL5pzex7+1GKgmnFxhxGNufJkS4WnGiBr6IKgdKxCk8z2ZFyUw4Y
fZtAnrZjPP34mBuQw1cSc2eMWndsQDo0PhxS31Pz3kMd3u+bXVNdcrrRkM6uHhun
jbXWjO65LzXCzqWO2MM7w3Dsl25XE8AuGNDrWctwOBYIzikoK5ocLoepNkDfpWSq
U3EDGr+pkKhPjZtN5FdHEVRWZnXG2U72jcElDGq40Su6DwkqcZauq2cQyqlRoAmP
9JnMYpsKKTjEnuyfHUmA7Gz6tgXngyWCwoU/aibFLgjlyZP9oKUpWcPEGJRmhRCh
dRNF2DUd/sdugKThqffLDbCQy66XAzHncDUAgXyjkf0ZKs3eTAHeTdMknFZHL7TB
ejMxfeKT5pEDKUtgxuvb5dgh0Q3JyOSt6FmEDjTX2mf9FfLuZAfvC/EEjRrY7xnj
aqDbQXXv87KNXqSj7TBroRRYROa137AzQyHR04Lz3i9sIR78OEbkGdoq3tpk3oXb
ZFeuTtXxn3m4ykBc9a4YHjJcTgr8S5tsg7AyxBPuylmovGWl3c3p+mZY/iTrLZLg
WMB3GE6o4EQwMeEM96kXWtJ0/g91IHtWh0E7TT3eq6Zh8RDT6SYnUCVpT7hdLGtB
SskaHSQWhTpv1YW0i5Y8y+7kcNWvvU0sWUyxeU1CycelINqtGbEReGiBjpp9ZEzL
Nqd5ACaRkt2v72GVKrjZJ0W2ZCZuzduTDUA+cnAuMhVGRmnqdhvD5qJ2BGfY0UJI
skr5qtNDf4JuDeJ83eyxsuN2XZf0qA6Bdj4Cs/5tuDQ6iYjgDS64T/TGtz92MJcq
MAtPu2WtAjj+RIvMG5cQUFxo050pBmIZTPQnlrEVX4jpltxGlL10E77NbZH+njed
lCNKQP1ONn3xwqGff3Ma7RzpPD6Si+40wCd/MsGuU7cahw8yqnDcAVFVQtSaC/ju
d8zCA3YRA8ex3viyHivMuAqghkwtqQeygVXzzXCJ+lSrtHBuV1g2M7oejFXRGWvO
VELmeQlL1k1fRY09omVYOPHXXmTwRGDf/ivAFy8Lb5arXOjTx+1v6hP8DEKtZ1KE
nOI8SoHpxI9q6hj7AoaXDRIoQ/MaLORPPq5toGPnJSA6AKwmDC1d5cFMx2FkAzkE
JAKI94bJmyRXs/eIaT/yA0JUprTEkZgP1SyiCijqaTFG06T0BipxUuWHzRoOXaD2
mBvZMrE/wXa07aFwjNltelPP3hUfe6GRpbmBskFTxXDMq6E8HyCtnqVEBDk+PRrZ
UxK7SW/i/0rZndoQnpcQtf16XVDEh5Bhbo7yCOQan52GFGePCT5w8P9qNvaQX88L
/k1DXtQ6gQDqpiebE/Y4jpL0aml9mqISWSfeBvuVGco0R0i2xY4gTJ4ANI3wpDbD
VK2LYnRR3cwJBQoEnPrYHqs3TheDV+ag0alY8Rm+/se5p0SK1cNcU/3fOezZvcPu
Li0URo+ntMlqzKEBbJd1NNh/911dtlQh7kvxDhOq6WBklCfcL5yc+euFCtKAwo1B
RcsLjLyhHQq3KGDO12l1tJ5UM/p2TFCCyCTQQS0AVYZ1Vm6vuI8aOCNSkNAz40D9
QEelwLu8Boz8HbNTKAJYmZ5AWQ+S3D4v+tYfN+dsDsIP4yCDhIdjNpBut6Ub7QI6
N2SLq3SukvZBdT2ZnErrB67PO9ie2WftFAmx14cWTzEARON5ts8YjqNlIAgyVyfm
9JCsv3TvPrfqpdn5QC4c4dl0h45hc7pJlKpdR9ISXKXvmu1D7VLn+IlIrdBs/LTH
j1kvOkfxL6Nr9QaXUNYWUxCqztXK0PjFyzeA6kon44tSJ3tLP1yIXH417jy6BASc
wbgSwVvDiTZgfdomA9LEiD9EQxaaLI4r6rGDiywwoTBZovodNgPwL/Jqus8mtQOp
Cwf0wAqEHNkOQCN0s/GMVILTIxqc9W8TNxUUKy5YgHye7HQZpFjHxozi4e3C9Gw4
0mZ816PdL70oHBmmj3mA/CPck4/M46wHt5NjhbdX4XPxtsLIda10dlHY1HbW1l0Q
0jSQEyf0Evv1RjoZK6T+JeXiCAGHeWNFzRG7mnGTe3aZw5qvp6Omfj0LTNNPqrSg
6jW2AmonmA0Racz4ghd2PnkSLwJkbbkW+Zn2ItvWnzIy/iBBW3Vohf2EgaGUAX8H
c4yt+VRMqT1NJhQqP3UDbOdRX0BTEAoiKZbhQ+zxlWEYHZVcteibuE2KBGQ2/sGF
9fLQf6MT9VGCt3EhzgHNjCjqQoV35IPWTHiA90UHFoQJWS/c3B3VVQzuxJgd0kvb
S1+WB2FAJsDEDgkqO2yjcIt6kPk3DwjufHsX6fIQzZkreA573AIg1GXUmXOt64bi
y7ojpMNQvzTvPZX5nagzdSBqmoMjKQz1k8c3NB3EKzzrKAWbFZj8qAMH3O7UYlZ8
dnoZbDt5CHX2c07h8ZZYNx4dM22tzLqQMQy2bsyeNQCPiMvHdOPM5FyLCTJFJb2J
8scGTE3AdLJYc+eoWwDYipJd1IMgEhZtdQj43F+XXBnDGu/AtvxWIiRndY6lxhFk
CuAp6blVrYK7FKoABGbP0QjqAjaomc7I4A65wPSxQW0Q20ogjxsnYJ/ud4OMdx0p
2UFVeTa/bQsLidKYwg7ngmG6zVIZWKOg9vM+Xkda8wvso+oocubCXq5TFwuqaNhg
mXCramnwj8VZwxvNTLrc0y25V63vOy3zoxWdNoB+14Wp6SqnA6CxJ5f2jaHvVJvv
dbzy6YhPi3HAvoNjxMwVQR0vxRul3aeroYUmeqGrjWT5F7u3IcEtH3/xrurpFdRc
b2r+j9G0Sw6tz5NeNRvH60pJ5i5SzWrpZIbFLWpAYi4YZTc2iqT5BKYTWVcn19PJ
NnJXGD5gaJETx5jucETOLeirbwEnJ9PEXdMq0Qifs1AfqDNmUb+HfXKkZ09SsFCW
ePl6DGiNrDLsqfacwyyn6H+cCsPGtzi2FPo7mBiBSRsLke22+cabAIvejmDJi8ae
X+pj4yJOadM7SU76IXpGrhBFw2jSMdml4uQuyJq08e+4eCoto8+q7uAhuE5AM4cn
yxG9Q+vR4m4vCP/KWIK94wf4sja9yyTfNkPNXm+DZZXR7OkpxRuDi1+VCYvpC94X
Ge8Vgc2XvlMfzY2o+Eu9QBl9Q0D7mSL+ERJTm9fleV3z8mMu7ihbaiE32qCrX72f
4iKnVFRrroMwpfuVwbCHSUhpOvfZFPmqO5iLm37N6amKPF2rwc1IG/FPguGDTz+a
e2D1b/j+/4UOKxZp/MAsVEj570a43PLByeCws5q8DbuDAWxnYUGOCW20yef4Pb4v
4laqagWKIVFznP2zlgl3Fnph5HftdO1liNh7Mnq6WdiRhEL/PmxueP1t4nDFbiH8
2Lh3r2uuJQQ3N9LHJA/T1DtUbDPdkVAI4lfpmqjyQ1ux+aCMA/ab48z0KN4HC3p1
lMbXSe4wuVKdxlBmMRIvEpKpKAC2gvycXknJ44dVCpWXt9PAcG+2nr9ZgzOX4zMl
jeOP8FWuFQ8VAlqHTerCz1+lFch9UiXPuHIuj2KitmGWWEuQYG7BFgDgwMWrdCQs
+o7jvrRwDpqbdM63A/Ehwqi+gi18omEt7opefyAz0NSuP7S+j6rIpSO33XVyBapo
yIVEsts4p0GqSQseKe2hDxMKZMc/BCsfw6hBcT+p/c5eOo+h/jOF3OFWopMlUJGs
7Dd9v57JdpJ9X0DGkJyq5Xx/1kgJGueygL2Dx8X7XCm6L+ONCWmGupYU0gPcWy1j
vlhj430b/1LOE+MvhQEpByE/6k8mY3eQXTNZJvRgngOqnpoCzl5HyjdYRWEmX1t2
pTopxW8ggVuOJ/WjX+c9O6XqXR39BrknsUS/5XwmvgWi+V0JGFKgMo8WRksF+WOj
g5UDgkLXIGQELwhnITpMUIBWXTOPVV9qLJulb08mAyiHL3Kgm3Xs6S4BGQ3KEOJq
0gz2gus0+Nqz8oTN+MvEHui59X6gsVsfUQikTPxSrYgjTEo4GtDy1MUSAVa7zt+M
IhFBd2+yIuxbz3q4FZEdZ5+RwSEcQ1atQeAzVOI31wURYGA7t6fUOHDoUHpXBenV
r51UY7vE1PgOHtH+plZ5InrwAIQ/L3zcT1j3Gi6g/27dWXa3vlcSctKB6j1ct059
Gkbr+poUiINgGcsuQyYnHmzq8VWstthA8PDq+T2BF/+DuD2OWaT26vAD/A6aJ0/l
oV+mnGu3iOTnvXXJqataa4eaNc1sA0OjI2PRknssIJT3WG/A3c9+nKyXgmVLhd+2
U/qkVXlQuhnhSTgEM6s+Un9/QumQYZiqxQmob66j9xTB0N5r4YCfTA02hqlESlUB
K1qe2+betDF75yqUHyq6hY2zEgyKX8BcdfTpfqgTU9RtHcOlmqDJQvyed4Mf9DYK
P7oGiQiOiT32zK0dKdYhjVNkyT9ojlC2Mfih4JRDWL1ETS9bk4MWteUmZnlZQwm9
SWVFAGEkBRHrJk14mhYKaTzOe9+cmzXXxa57ii+OAyVlJT8dkzPQsNctW/FU0BJI
m/N6b+KqGQdGQ+W8KaRh6isT2faqgfZQUkJit/hGLdQiUAkx2L0sgbhOgW5lwpv1
BByVIIXjNMNJkB2/ywQDbMSRztJo9xM9n0/f1Y/MhMTLGtNR34N2KabKsFcP6mUd
My2DCYQXVYRpDFJtyMyU0Ggj8eXHlEIo4T1/jWPS+u6lMyrQ5A789BIHHptbLhLh
WWHjT52UQWMMEsnyY4KabIipn3NNXNbnCkzMM74HkXWuHf9pwljiG92gPdgTooIU
UbWGyFFuzmMrgcTyx45e3vjG2rUhR6XHCC3FAwo0EbgPvEY1/G10gDS1xCnUeVnf
2pyPQYjaXxNlphy9VVhLGDgQlDKZ9Eut3y7sE+f9IlV6KXmOePL8XVrAwMjwXWxO
suYNxdJs4dMAtNNwTPfqmbgGuBuebpdM2dk201Fii3k2unNpCoEK4Gd4snZnYnOQ
uD7D9QrrCSXXmWUI7ZYDO8comATvAI/jtHmDZJKHJgV7wUfqiyBWEPxnOxnWovx6
DGV9i7EBXL+agUKSObGeG4b8ajtO5yWsIaDd2HStBbjwvPh+1j+hll6X9+X3tkMR
mIACc6oP8zAbSfWpQbCnbVQw1Z0vysa839yZXRzaYqfUyzRr7gaRrolcLLPNUY5R
fV4XOASbwp8wEA3cRtFkNnFkGfdfrQASh57ATQpluXqN5u3eCH1eAYXTwgfNqeCh
i280xh4Vdy1kMODgAcrjUqM6Jcw1zND4iX+oZ8ATcqgzwnQGrjjMwgGAXQyBgHIZ
00s4p1zo87NNZa3LlmAyNa4i723/3CGrfVB2xDHjt5ig6HTTpScSgO2jc/D60bdE
Pi4Uxm5hYneqEEmrIwGfseG9/NlPoMLnIIVdXWN/LvDtqtELlGKJVANU/sSrZNAc
MMEpZRnKi0Nz/E0/BQIJcfgIOJ/mbKiV3C3FcsSr6Wxh4HKTj71jWdCEouaUbpxu
offLJSLJi9Tl7YDW8RrbBKKE3Hz8GamnPIoT1unlUS9CIUgfqLQG2j3PscvpeglI
ecXIkOaljwjbVAeKdtUAPPPhF2kB4LIsq8MIL5+VnxhV2l/ZaPMgNBt5iH1WCy6e
XO6o5rPUM2E19yeyY2Wd+PKLy0pf/qtDnyrlccj1GKm0o9oKdI9IeJai8OqB0Uvy
aHII/NOt0BecuT1FhqPnTu6y9nSAEUOwPqHQR7GR1Ad0zampZOD9o0zevAdj9B9G
hjEdYTluxIH9Mx+nJZT/B9j0isEEkmC0IaU7Etp/CjOb96s5P1iVEyXYuCbMnWW4
Rz/ef13xgt+xIU0SaaiP/huNBD308NjR4M/r7X2yre1xF3//WyePI+5UIlg4vDIk
bH399RGryi+HsUzsejJz4FKbmIjgge2lisn0AI8HjKDMkiVgc4ut+WHSD8l0J0J0
elorTjIQj6xu9m31Ppbu2BfyfNBiLIWO3LOO4gGKtZh5Z/Jft6PHdQ6POjLHOOnv
r7IJ8+52TitGxmrBwoF8YTUwOaW+i05R4/MZI1eTJHjhVNx9cTUIoLx//kpF1LUq
4V3zDQIlSkG17hfyxhzRsnYJyYKC5bPkJO9g4ARYXpZQlQzZJOAh8GoKHTxBuhg4
vvezvcxSEfxEpFt9JtQijVt0zZ+4sFnj/Ye60L7I/OOupAIrotJt2EFAUG+SV7tg
qZ2B/pNewOVggMK6ryME1mbhRHLYzqd6MHNjmENYVgbEaqzzAAmr40xzE0CscQMf
eCx9wU0tSDOJzIYpTUa+vDNlLcoYZdIGd/VX6ScKqc2Q35SXspzU3taXgLunJJ9T
fp62O768InqfCFbkgUvXCR4xuIzYFpMQKRmXnM1FWAsfbHPqkaPHQqodVLDTTxE/
iVpo6fxR1a7ntdcu1HyFYsYXtJo2Cm7w3DnnLerybZJGXrTz9aFo+nW0+Z5EX07u
yXSZFerUTZ4cc5TRL/zsNTHWnrFjriO2WSb7iLOlOk/XP7G4UOc6y1x7HaR8I3ko
a8hwIUf70X4wgScaSsO3ZRNMyskvP9aXBhjWWEXJnv5SF0R02i8x01L9ZGisOuea
Uz0aEGowTHHUEcS2euOyuHSrYJofX87taFzgxmKGViKQW5VgecZHC5V5JsVpfYG4
Nl0V5XcmtMZCZ8e66KIZA8M9jtUX52A4lvqbI+iy+ciQauvx6C8rtAgPRZBXyFPa
+MLFI4v4eYavgyEnPruW18LuXB4RBOR5u/gh+vzsvZrqfiOoCMoDsJSWWNFM+JhS
JDM+D1hsYs0pHbGv1vgGHcVAu17UATQkzVIFCZH29a01GNx8Q3xosNQmRSVv+BhJ
IIucSWN/ds0xDNS1KQ6A1LACPxnHG/Y7c9m2bXcG/iSWDfNDCjvsJC6v6UzT2j5T
BM/ddW2WPBhv6k7YiO6v0tgsIoYIJR4BeGqiQ4auMcVfjCldq+1Ejg3y3lo+LAqI
FHyGjLBGamdIQwe0k5S7/Qs6BH+L9NkVCOA2GTWkq+NpO0z3Ile9YiOPkn8wA+Wz
hWVguQK3AFhQjg+v+uOs7Fg90kKFIy9GqcAtIhap3VEyhoyWOeGpVU+k1dZ1jZaL
qmcbfrqHVvf/cw8F8AbMWIR97heGT010Ryzshsy8j6Y+PiFMYFnRvTfgDk8u14KN
31HUlnFJ9VBqX9l73hpS83zwa4Xo2ZxnUbMNjVaKeJGEWGZoEGD8RGMkzqP/2WoU
9T6CceEUVGCkMM/e8+BGHmSI+rA8FX26UxYfiIkDUgq18rbVJGOLxgwy2tcD96xt
HvOBxnoGbaSaagiLpjPQoIR8Z44/3Cd0ml/kMvJf8n7L25KG4XyVKoAq8Kdg/NHa
tN24FhiZQK+Rue0S82w3Oac0Fp45/ko/DKfuDAiKDqfAIuXnVKmHYBbGIO0dG5Z4
nhQ7oF/PT4At66/RQCEyBGNhilD8ZHxP6E67FfrkLor6tU1Dsr9Tiqw6TOJ5WHs8
/2jSYG3RWEi5qPe3jmHj6ai/C6zJsA6f0hp6rPy/0aHSgwQUEERy3pboMRJ4X0sw
ZmfWXrsv5RRSaAr5lg8qhzvUaDjc4crwE5AM9RJ9LHMtRhWSNygQKmkBODzMkZl2
phpest3YnoIWdtC/+793AtalLieP9DqGaNEICeRTTSPbvCiGmaLpJrsD8FxIYmJe
KQQdBo2BhUDSxjj5FoIGwL28ZGINRwfJ5QJTJ+HtciFy9Gzx+/j5EaM+gg4KO8OE
GsFYmkR26YCCSIY9SNoSRR1pSVbNBcEZ0I7FJaW0e4kTuc+K9CYfgGL20nFckm2t
RFxkIcrffuTrrxiIBArtGd0OIYZzaahn0HFDaLd6YpGaWW50nLtf+Yi8uSCpDFJw
KECBvh5RCHnE4Hx/0eNMe/niCDWAVcIWsSEwMBkW6RoVy/tfy+V0e7xYQ+28cArL
VxcXOlITqMCLv5si1RhNQ4ikEE4x5NlGXTlnjfWa9YfdyxZX1kDgKoT8j2o+MsK/
A4ivlctLsOmp/Wa4jVe2BcHU7Nw4FBf84Kb0lAkvT4vii6wEVTq5tjT1xEFp5CCJ
s1g8fUMy/dhn/pMhIxMHJXsNX8QO6eoR/Dn7++wO9ms7tkRKBAgM1MX/49trG0Ee
kJYC6y+D1gGp5bMljDT5Z4HRm3tU/Hf2W7iMBh3SF9VyOHry2ST0qp8hCuamMjxJ
3LRuQ2G2QqbysavQ57KV4Pt7b/uA5YLNMkXKN4zbT+yFDanhQTfmMpOdgrL4aqcO
0Se3RW/2+SvNM8Nkq/RgMNOPr/GzeQMxfVFM4PlnSX8rc6eyRf2Qbhs9wV6G9zFH
kvianpW7F5CbaETxE8ux4EgkL4o1W2JZZ6Hiz6WsAu3BeTKGbKVh1hfd8lc3nWY9
dRMgFGJf6/EOTLCO40bIltXMnK36MqrB1PFaFPo1rZlrdt4gFl4sz4OV7CP1c0/G
mT1Oskqh0f9xlsyArsd4CMAkdKNJIGa2AlAUrL1ABybvJFxc/0RpRCcLvDbQivz9
NfCoF1GrkS7b+wWFcxubWGVe6aEZJtfoPu7bXBre9wGyi4HWMwoQucurBeofdG2m
2qBpVL3IIgMAis6V+4dNpLeOpLg/qo/31nf9uLmKQCPpL0RDitK/AAeelNcrnmBK
5IEeiStkuemMZKqu1DXtKdVpT1o3G1irEbNDuPs0kfxBBAxVjGYE0YHUnwPetRtW
suqrLipgy5SJrwORaqxYsSB2M3tcXLbJAIhsu1TkfAxM33NhcHD3tta1FiuujZ75
/+LGXV965HLJfI0d47EKPPyc+tm3svtjayjV/lw6FWSqNdjOeLtdw9dwjUyz9bhL
c4AuN6es6kQAie7F2iHHtAtQTSZTAipAnru/4IsHjDpns3IMaWaCnmEOE7ThC1LB
dQnjBjAekckBo5TWjPMR3HvoUJH2kEp4D+VLM7CGSNf8T2W1a+gLaSQKj8kdSh8o
GrWP8kn5et8f5os50aFe3E5Qz7H9jPyE4ICw01IGLJs4al3fWiWRaCx5LeQ8Xg1s
CyVOf1XDyPFavfsPzkIIuELSg7rgc+ISzs2I41bbWwumtkx54URTs1ipsiHFSD4F
cAteZKL2VInTtmlIl55aN3v2WrW2tUgHBR62x6WBX01Iu9M6LIzXc+hJK+6wj7UB
2NkSvw8R4cO3s4ixo0MKW+qA3pxtDIAg2wDoys1/9u98TrRI+tH24Mas1k5LvKvB
jeT4VKM/6LG2XLiM1ppIfar9ml4BySZvgv5E327Ztw0eAGBD+XNOMcQTcyjGIyJI
gyk9upsHxtKyDk0TL+RFzgnSXAfoTrQ+ZJr0ak4O4FP3wWp8IpMXcclVpW2nXVpl
r+eDqIDZjABEpnxucGW2ASECHZBWagimmo5dqW/OvB0tClwjt0XZ9Z4s7+ZOtWj2
3mTSlPLOOgOA6nfPO0w8DIIuRB+2YIipQitZKXfIDtSaIHbCS8UZx2HEF8iOIh4Y
g9k0cd6f0R5tmnMGLJav4lgPIhKqxPMtmZx5FiMjW5JYYhJ/+lmdy6SmGqcD1Ar+
ZifOQuOfolQv4P1XnDy8C69BRFYja+dVhTurPySjw3yefGNCrS6A7Fr6F/8N8wA9
/4tKKDV30DJBCeeuUjumyCBmTG2cOJTo7xLBSbUTBIwDBC9ojBNWr7B7DJwWUZ3j
/KWI4QLo1XTMgS9Sv8r5kSLANQl6WLx0MiGNPi/u+em05535PCGkt4VMqQxdmyLg
GYMxZI8X7n9wHaonhgSd/95Z3sKwGnWW1nAqiUIJCZ3sy29m7pxUsj7znpDZdtU/
D77hgPMvMD80OL010y61sdri7BGeQfJCUw/dcawc7hubKNSr0JFCJ7rjrmg1CZHp
RIw+H1d7MJiQyWqij+zWzcsdSANwd0rw3G43izpT4pZ32oHmnzUAcd74fELqxGJG
wql0yjcvUYf3I7ehVofAPbDa7a/QRF0K+3ynzjF3uCG0ed2xyEYPLUehmJiqGnC+
Xu0cTuc7KD/43SQwd6ljMlly+ujHn080aOxBZGQPqeDkZiQ5N8cj16CtooGjevGG
na/6JLibRaDEvjmalNWPv8s4HIWS/zY8u70CJJBLbXvahfnKls2MjJn5WiUzWf9r
l1YXz+6rASzlhAPl30Iyk3ys1664kGllR4nNlmoQhm08pd8xLdlBIFZ5qYJf5o5f
dT+0zynd/f/MCHq32Ora7AgI4/iPtCzmOw0umPg9y0axrbhKtUToVcu+pH2vnrmU
PsBJjDuzsDVPG7AcbnQ54ZO+WQPJNpfWlt+WxK/gjan/F1urL6TpoaxH+fdKC18A
apfgDjq0w/CcizuLtyK6LIoCoumBVW8LFEVKoXscLuGS8r1IIwWSZjza4omdosod
uleWFD/1luGXoX/FrGkL0tf2Pwzd/gISeh/ta9sl5Qb23O3gVdDYqRuEYia0qsKh
ClCjId+xI3Tl9Cy0Hmk87QHzI0F0Sb3gtaReo0KIbAcaDtITfXu3OHAuJDobNrZt
lYF19CAiVUtHBmodMw2sELj5c3yrskXJ6E/0fOpkHUCm0IUzEtsmtYXr+cp0sSIV
ihkJFUOgITBPtFAhDddqJbzHAu5VrRmZ+YH22ShukDH3zt5lTZxxcCaykrArW9Jw
BQfbcR5xcDPyi4sPs3MOluULfS0kyB+xqN+MX6nxfuRVIvaEpLndSCoc++LYnsD3
Td393WtSnbV9bqmlvwCvQQjytGy2E5F4coN+JwkbZYCTXHw6HNVotFN7z8mUgUHc
ZRAgOlZbFu62hCz87S7ai9KTgXzcaljTbGKKopCJ+Uh6vHJJq5GL20iNFcigQubp
oBSqlFTrMbxeXOcrNXkwIAeU/yLeAw5Jm0mhosrI+30m/sOPzJ2DKM1pRi00hyB1
4Qri6TozfmyriuR44qmJABipDXMdAbnv3/Ss/7xSX6rf8tYSiTrvzftz8a3Qg9Ic
BspXBDA08Y+VAZCO6j0OKFnOY2jpD4bzhDw1Smt8yEdgpdonlnJzNOd20Df17jnz
mFMo3885oMHHSppNJkA9acOjCCy8eZrCiOMuFTxpn20Buj1Kmkzt6PTiZ8z3jekt
MoEnU8penIjNnadXO30alngTgVkiL4oXN4pwE9ZUCiEJy0SUWKCP+jFly9PbOs+v
CHn8vB+EYF23LBk1IfNr3O181pPSMIxl3Hn/VjX9MIYM3AJvB3uVMzUV0phrClhS
z1ihW5oYlDOIzqV1Sc3D6w33taSqiwFO/JEb4IenHJ0YumzSBMgiQISjVz5ZN1T9
BUzSOmlRSPDZgprhWX1sAtOsrtGDrsCX/Rm+x1hb46cLPB8RlaKH0vdn8eOngy/C
R9niVZPCc22FuCewhCIH2/cfUYruR6axcVdYHZd9AqS9pq3B3ZmUcwSNcpviP6Me
9WimPq9e+z391ItzWrgEXQob8eZo4/ORSfO4abZHQXwD3nJ6SgnbtR23FGUk9KmA
+nlgLOb6mfiaN3MqzFyWAQbX0XTONewbBtFaB0FsX2LXxnEMi2h6Ta3icNmP5vqu
hRc6A0UhWJanNhV+dLxKO+BVVMXt40AgmkFcWaO1T/vOOWRyx7zbsbVAnoOWkrDW
YxZSYv2ts/+lxMWaACWiaywq9SSROttyB9uN+Yfu4pshKsgYipJCkNJNVbQbHmcT
KKEGqbhjaUAtoV6JiAe7OJO6NI7lwOxLgcJ1Lau1mKcSIgqSzfTD+MjAeqqWhK/n
bHbskfq97M6xihzWya1YEWHLGSburEnbOfXt4Kxq4A40e1pjuRKNFnB+jpBd/pD4
IpZt2Ux0vKr/HKoVoSoDYNs5Lqo/IYEPwp9Rz4Qp2GzaEOqeFsCkeEnppyyBBPS6
BcarP/msT6pharHC7Ce2RCyyT/d4I0g1RQRZxtolCJvqRuHRkISEl/eztacEJP7o
Br//jzUc4Ts8e1R7budz2HozC8opcaaRqIYAcSMIaVGXEGAtS0isvJqeAEmMjGuH
SA0o0irOko0PWsef3rifu7cWntoK1DGVH4/4f8fdKVVxIwD1r4LyqvV7xAqqrJQl
xXEe2FniBzCMUAKsXlDj6bg1+7asqcajgPjnFBpvlgk8g7CRtOGVwK7/PJsLBLe8
ATkRVrzZLHSt8ncTSGP0mV+mORGERWrOIkUhkZrDJhmC2oZROwySaQ87JVybHpSM
05ce5aHrw+LI7r9DsRk17xgoBmouCR4RXhTQDSyeH5zdQJyPfgyzsZPQTrrWyVaE
o0QwNXVTXE4AO7ldLqzQseFNedvwgNm9Ih7KdhQonjCeiZ0zhcBLzI+C5dRdqtr8
YQzoUw8IwKIIUjZixY6vm7T81TZW83F6X8x+2Mx9jfToMj8u5Puuwzot/mCNC4bU
Cu2v+TBRGHpBp81j1lwxVKCo2EbGnt9Rv/P8Tzr3qsU8do3oWJrIpQNSFUQ8vumU
cFdkcO0DthzSZMXUNwpx+2JSXhXQl8++VYhqP3uMJLTEdHs5Xexr4VmrwRoh+1fD
0VRlasJn08TT/lY5I5TEojrmvl2TmzNFd/7HCQVO/GyVYSPEwA7nYkk44j4pubJ1
i1e/2HJbWpvhxmPcL70fu5alSEdgp2VCe5is8Me5aXEBBDXbu7+olTF7Wiu+aZCg
xSsUYUa6FVyGps3MUpm2UpjRJYSEaBclqi8IsArZ41lmNpqeuQP3YAoO2V8zBCjN
rqmaNyRDtYLsGpBNYEeZtfXo0fNMICtVRdp17Eld8YCucZs31txYr7p1gZRwDbF3
TqMUldVjwkyY+BGRxuCo00SECGTudr3n/GpqXH3Etfpasu9svHF1CuHVbH86zuNH
+PbR8d/j1Mhd+XDm6MtEGENtlTOb4jR9RlsqwpBh+jzKmLJP71D0GPMPNP0B2e7a
PpR1pAA6f11egaP0GLAJJMkFhIJh6+GKhH5BsLdNFwaupxinB/DtSwRk+XnKL/vf
cUeZa4iFiQtFu7ibVck7gaarAu+dC0UHFVcitEf8oozjfLZrIHi76nCuqc7NowXt
ryY6t7M1Xcn1z3EuDe8j83ftdD5xFiP5Z9ZFVC4fmZ/IBnmy7JaWWKp4aztDXVTb
hqXNgn0XlULBZyoPFA1QegYuatpoKxwnPQ00HNn2tE4gLohGYViG8KWdNHxD5Jiw
kWRaooey7Npc32Lh10TX0u4mvnHW2hWlmLQTzLABGS76G3K6KzFJYwTEZQvL3Gm/
TIBQQdrEbknDXomDWvyxOE/Zj8tF8Fxi+OPRBgsqX8Pvi+VTrMiUU1Yb/yaPqS88
h/Sp6X7ysvkBod+yKCJh+DB0DL1QX7CxEptDlgKk7OAcuiAzX64I1Z/JMScSTYR9
OGa+xbexwLCsL5r2JTBiFefeIw0V0ZGBP+EcWFToM0uviv9CoPDf2MgBVT6y+50S
H9V5hqVhDgWibqw1o8FeQ1WTyhsZxCAIN+d79jBx9bTCAmUt9WmXP2jPdaPITUrk
xw0xxcHqttaSDtFph4NbSoN0JKhIKJLZ/8xl7vYoRYCbsWTQ1L7/3mY5ex8etcuR
NPC+AXDTAIHLb6HlErD6akKsMow/aru/6GP5cTj9WMf20CYk8iJkr7YuQpoHOrqc
lus3mtaac0ZwRdPCg/muzlnQuabQDEZbFlnlf9iUGw2Tw/s6f+EZhAVl54UDXgO6
8XRV3Ny0aX2RdvweOnugi3UCSC+rScPZJpByAI9uUcpVROu+Zjvb1v23PCTpIOp7
7hfccd6gWk01uNn0o5yCPSNclFNZ+LzS3xgHDVWtV54/8R3/8XOtglmxFWRDXeCR
TkIghr+zZkDJaj0Cpr5HsYvCmnNnQR6+Sk78F9ro+ftVDsBIUl9J4L/vE1FpniWq
/Nl5Pyo2d1hY0JydrhsAtVjixAt+mknb/aJoo1BybZUrtqAcaagnVEXZSTzAs0qf
8unIDekxlAjvdNheP9O22nMXi2frP7XH0ugjjjDEmRoCDdzMQqVk4FdtHavRBOSZ
y/g1w31Kgdvfeb1WgW3r3XMMDfxTABszcerIX2FM7viQnp4V1ePRg4H+z157F/07
1wSTFnzTtFy2xtVnfDkgKn2v9QKCW1BL+Ef9OUkLZE+/N1AXlIiQ6f5J1wBifoT3
dLDFCOnHKaPMSiEXnW89RVeSZDs+c0nqFXWC8+YPHqoqrIHazLnpA4hufZvhDOX6
xSJubkheQRZIlSzEiSd3bWiaAQkH57MPj2iCTBsige7MRE2kJd3qZ3lX2tNQxf9J
0wb4zyROmkwj24K0CEXabjlL82SNH1CPXYJHQJXU3WxD+WucGjCkek54QatYatKt
mmzgywIhw04/VfFZ1TidmmyUSFLoJ5Miqd0ABzq/M5gjvVgI0WfncVcQ2bZSOlJN
RbBkhLadF0otX3/2cBvK6ltiHKsYjnO1zLkNfxb7RYhUowTDnV86cCYysOpggXj0
7wWTuKQS6cUcp7nY4woLoWjEkD+aOTaY7I3LIwwDUOPV6HXqAbIeZKucxwqvSXJE
sF1MSGX775tQWLwEok2nbRN6ma7RzwFuqMpDXG2iZbtpm6YAXo2Te8PfTBJaDMNV
pVUADlQRJ7X/wBgUMU7wqTaK0p/w2piDI7vDTgnq5YL4IEfYBC+FcaPSVeRXIW4d
DutGgvXwzxGJ3F4gYKUK3/O5Sd9eIROVHH0nR7EzJGtTTkdi/xa42pDiyu4M1J5l
ovNwRZidSmM4oHtJKk+hg2TZNWVMYFbxEOIUPUJxZi9B65eCxDY7pQO2UtYwoWyZ
IE1uz+PEaTKudY7U4ycroGu9x5UCSHmD2diWpRY7cU48ZILHOzK7NrFZKsVj+ySZ
ZrvEN2RUtO8tbfvYWQYrQksD1UiM3kLH9hlODRQBpskGrmHiQNoxDv53vmYFJ9K4
JQZkT1dtwzgkajWATJi+NhXX9RKay2HGQofX87M8Etb9U8dh9jo1MbOFPfUmBEKJ
yWRbuNegSyjmKTH5IEAMAWe3WNOslAb4mWGbemvLhwXp4GnCJR+w84FlM52YkxF4
YC260USYakwis2PoOjg2Cogo7sNkEmYGq9Jqt3PIgiYs1nTUokyrtgTUdet1P9P2
PRyflmft8RU/0O0nIh95IGboj9pwaBXfOFNUu9vIiiqjB/UTfwWeIHI55u4UGfOl
tg+h/O8E0vE2XiCsr06+jWQHjXZkKZvBRWgryYEx1DBCoSc3xQfb+qOscaisK5ER
v+I6MxE+tRShIRfD+IxRbXUjvmtpeiQ7g4Q7eiBOpQyqTG1TX46Ekvu8thR556KN
iEpZMH8POzYmK5rXjA9zvCHKZRv67ROMNxND0LoahftH1sFnCi3hcBEJ/8WTm5Hs
PV7s30P9QFLUh+m9m/SFZIJk3Op+oZeCIzjABra0VHSl2Qku03bNYSzhX9JWb+Lp
2qdUmnXqH3QqrUZglM1uSukJfdcXScFtrm0YPTx8ZogrqorJBmTdbuPrnEmiK2KP
sStiEywmcNoZy4Wccu1XKhxzlqbLq7RrEuTDopSd4nAFcafxxiKaqCFKHPc4259R
3WsuGfNNEG6/BltNzpr+MQ4XpDoEjjX/3dBwdx+JE4gm9huxRaLJEUqJocvQHu9g
qrIgG6KzhffgKGdLc/BCmmgCSOhO1BN+jDw5CYcb+ul9rhrgn9ZvoNOSWczpEkiG
h68YyKvuLti4+doKECAX6CtOhZ421BIUhTgm6GldAspz6Hfq6pNb/akQnIpVro8w
nz6DJkSV8MYoRS9h3d5q/tHZxBqYNtksnh8uKz3YVosgZapkfuBlgY+zdZXsZXQm
6KN4BfSAJ2Rve0VPcO/59qr6PcLFw7NhGVHq5+2BhCTUYY9NkkgJVaSP/wqfyn4w
AL1c67fvXZwhqRpB3oLBYcp4OWoUBay3VLrE8IdXV9+r3pq5CTUsOTIsIiAKoYio
1n7K0v3GJN2W54BeY9O4sZdVHL/fURnSDWrr5vnQUTqaKpP5MghCWvpXe0ecy4hs
/szOOt7MT0mWHmwCm7rkjkun+QhLU3R3gQlqZCRcnj7o5MzbJH1OQotFcH49ahbw
VmclO+uBV7VFgJqwO1QnVvOWtwG0uQwLn73xqp3g2TwbjVo3nqx1KfdmZibaSmjh
jlevVXSmVIlqTBUZRPshusFKxLxbspbXXbbfOaxknCvcxu7x073UteiPTotY5ayL
2Ba6Dt2KmkYqqqhFjXGCbmM/gj8XwRWznSo+dtyI5MaIl0qu4JWseA9V1K9Y4i9X
kV3A/7zV3qxdRMOCUyJSAt35gOE/bN4OgOdMDFJRJm6qEzuKDCYathiIJoJ6t12s
khMsJbQAdLmkXcrB5jGCxY8f3A8x0UjhwX4etmz7F4xchjj40r+0xmFE9u1MQGFn
5Z/ieovowBh+89G3aKDfvZDKJu7At7mRPOeWlBCVZBRqAey6S5pX745YEVSfVMOe
GZLlL9bOuEuc6roib1aNkljcRfOrDVQFErjzNnHR/5Qb1QFpF3vRsQNTs5gqt/9j
sKmlqDFbgthWjLdMlbehnZmBFawpfbB18V571OpTYSUY/DFWjcnpRs2x3pHwXpns
sh2IDz5tMHWcPOJuUS+xzXCOc5Ubdhd4TLlHvSC6/sUeTv+XhEjhf0UGj38w7pKA
eDw3Zdz7eBvBsEyF4ANSE18cRj//CAHoWz3oE0KPAbAWbnzGMyFfB4/wdtyjEHKx
oOvukEkCm942XDRGc25vLj8V1xJwI1aEl5dz2F8UWyT9URFt/FT/HpadsIEgHoQ/
ox6in8vEtkIQwTQ/z4U1tYXpCl6wLx6bAcydSpcj7vbftHYtVtRij9EIiaIct3b3
0YFeP6Nl65jB5wiQ/vEVtRisCOdGVVtGEmJKwN5h9AGxnAV5Nktn7nfXkN3t+PYN
hgHYh9BeR4B4ErL3a95VAC+fiki1iPRrEEozACMYyJ3pIxMH4NnkdDDURbuHCnlb
y7Dqb7jTJb1H0l0AhlppNlEULTrS7P0q2tykY4wpcDPZEmq/bzMTlVKYz++Kqpg8
By/4hvJlLk6UvGyllJdByqa4FY8PopZlEAFTW/P70pre73KgYlnPukuq5wJaiMMW
Ou1sSSFEov+eCiwXAlX4/s41ab8HgAlbkShqB+Rzl6xQ4PAWPBhBWYCSvoHjgua1
WXWggxf5XsRq9MShion2RM66HYDoSNqq1LV3I9EKsDqBCA2SwOSAFQwMjFjTj4/3
eMRaU2796i6qbDOR2hs0fGU1+ZNZ/0iXk7fZtv8k4ezyx5FdsPuqml6DnLWsFs6Q
9S5MjPLFQmOBs9M2QwbTcVd+XRpXJO5lM3a5DnnpqkIQnrmkpXeHIG7lPMuVc6xJ
/qpTuhWcvT15zVq7EuqrgfyVvpdZFixlPBJ+PkG+dvoGoYHyYNvp2WywYAATyvOG
euLdxh4K2Q0npyFJ3lGxCfT/C17d2xdEw6mwXhzyiqy7Q6/Uo4hOhcZbbExZFSyA
iIphaxh+Bs0M/z08Dl4nj3dkRzNILsUsZalG3trIBXc7gFxSI6f4QneLsD7iAblK
f14ENwvJywCJnExUBsfIvVElhAuSbGtYN8BhaKGHz7GeI3M6cHKME0zCx44q85T7
DrnjkBuhYFsLEDsCcdSp+44P/kCCG8O4D+P/6buzsXuuXyJqx3jQtq4p5TiVD4HS
ZYN0yNo1SNbrrNB161fnYRiX4WJGUxyt5Ni6/KvXtcCwULbaD1aAPwAbISfQUclq
1npyD/E1wWYpWtAeWnP9cfZL0Cf6EOmQfI+p0W/ZyT21qNT+UXcVK6kd6fZpC0Az
AIf6SllYxpFj7cKyhBBuRliFYsXnKA3JvlMNnYKRWfJox86gx0yk9rZCm/p4bMnz
ukJXch2ZU/2wTq2uw2Bf3ONN2n0BB2tFA5hlT8pDdK7txNzR2c/+lEkHrIqQ74jy
b31fKUtvDoJUk1gL+AcZVOTk8qXlLMqWnBoxrESUlAlCrt4+Mal7xLOfGktx0xL/
TuBcZu/l6UZsjY0hdLQAk360iPZPBtg0s+OQMN1+knnm6FrzVMC7ThU1UsWqBU2S
vyAqO3IN8sQdjzuyVIXj30oOXteuLfuBndxjFmO8HbfuGpAgJRW8o+FZ6pHkW7di
QRAEM5K9oOKVBDAtB5F4pK2r1LrQQhTioWJgwHSU+xphf2pp+6xhERNMTh4pRTrU
ZA+ibX2e9arFWjiI7y1IH9BGKVMj47Ov/hwu00RE4ftzs1/UzlbxR9sJpCh8GeUX
lL6u+wEt8ZWUwuMCGriQ1xkMhvFmP/VhWpT62AFF0JAU90hH1SjyU8QzpU0DN0Xj
BLldiqDh8j5tVswVE7k+MzmleNp6nbGgNRbXmP5kRFU9I/pMoDIdia8BBLkH3wc7
66SdxH+zVg4QuOeBm5PNCLFmgC06owN3Vm3H/sG9dQ/bPGq78qPXm/op1CDaAkZi
orCCOAvDqG6cbsWT8prcJnkreyLwpUFPx0qGZ1Ai7P61kOc+id57jgPAgqy/nTbb
GD2T6f4+zfZIgLhT81dd/GmA0wPy6OmUZrnWOKaRXG5vWy2xs233rVIHXYf5Yl3M
AQQQTzlDd+GxHCAw6Eh1XP9zwN9g39/4Wz84yzQpgeyptkgrfzfnLgcxMNid42xy
XvZeHMrDi6MI1CncxYcUBnI3bLrn19eOIvQqzjamjW3N8R1M7blfvyg6X6TlDvzo
ozQZmrVHpW0WaBM+MY3BfIhX0MhTIHCj3Uhm9w4h46f5lc52ptYEB5anIb0WpdFM
RU5LusS39TyelOPtF7RxuxKnrV02ic4je3R9CuYeJTKRac4YKUHiY6OGDVbNsG6e
NQ734jCRfx0mhOIM1nKK6xAPCDHfmoHrbGzABB9Uf6c1PsSLarDtwxSvqzxDSdbZ
vugOJBSKDT0+LyRLH2KN/LCDih4LypVHaWpaCLx48JXpxrdXzSUY9g56kPzUVwwd
7F6kjoTMipjifoKYV+q67BWRAvjN3JeSzpFckw09wNeiSWEunJfCC/HqetolhOqw
jpHRhq0SufX1sAMv0JHy79/+5tvPS6n9M5eu8ifuzZhDxYcU17GIkCR1npUDY1/k
8IqaVHVmxYXRmIedizwp8dJ5alYqJrYUdlqMSzQTPJKWmnb6bRxTOx8faHO+w1pF
pSr//9Ykfw0jiSveNGU2Qxm5v7LBf77wwlhgZ4cKs6Ga+IJWlzjMCNr1sy/oA2hD
NoPMRZiuuQ2w7J2kr838Nh4Jgm25vZ4AuKH+rEEHcwi1EKBT4k4PqeNKbaNiU+5S
XCGCGvQNyWk4cXGBedfwCcoGm7cb12Ss2WhEDsHARGhScD67o0svKir+YHz6fJ4J
xM2mYJoqagtshhmPsas7wtXkWgQUSY3BWKQ52wu2AhkuSv1taptsSAexSoZSyVt2
BfVqyg+t8Fkk/QoWHBquBBVQWTLUQOtefWXtx8NUqlgIMgD++HVfTlaD170REUqe
jX1g5PUj+SrwSZhrn/VWj7WSM2KChQNT5UlBVX01mc7Tv6sMinefmo+dbqlx7IGQ
fPdCvEr1gpGBprAjIcVzR1+x/SsEv4QfsFWHdtvy5zUxnvllOszsp4Pr/A761TeL
aYLX325d32oO5E1cCKoB45uaq9I6pHoK3CEo6/gJ9kdT9jjMLPxcIDa1Z+ym/F7H
cEXOA0uemsXg4hljMeT/0o0llcg4NvVo97S+6XYFey+yGKDPktv0GV/0LjBdlWFH
Xv3voRYPaRhzvpws9pSOxT5M3Vu67855Fd8jlRZsUYG1BhWRsCToTHn5uhjrFxHK
0k3VcpwqWlkdF4B49HrhBvsg+eI6Vdg1UrZlcVoW9q0oA0XwzdQisIzNm+WVG7U+
GuOg2pBDgLIaZwEZwObABZmuEgX62JL6BsMqd/EI7Dh+eW5pK/5dhwylFRnFYRSl
ANxpQA9vWs3fAqfBAjWMckl5CV9fAIfIGMSuz4sHCnRp0CTVHXbMG5OF7sU0vRWr
+Bi86mbmXoBr0uSl3wEBv1CfROQWpl5GG/auXWmfgY2xEPG5I21eBRnQIzQ6ybrC
i/kzZv8LYpr+aQJYc2+v8KvPf3CdoKp7zL7Y8n/vX754h9rn2QARJMYYVrvkA8fk
juvPAy1xrsiuYahS39NiDRfITDFqzOTxydzERhYrtbCF7Cl2LrMQzcujp9y3GpEo
0Vmxxi4/HoUEQ98ZabEaucqkoAPPowjzSHM2b1B4NEBKCuR+YfuyjnR3s6opqmMG
SOCQsQRaBOa+X61yo33OPrjmI5mBLhyjllt7o7xDTP/iPoV0EzMz99eNCbpDVKtj
5saDC3Ti2LFe3jctO6h2QsjNwBG/cJqOo0BhmzUOAFCp07bkFTKjlz+gQSo6T2Xb
UAe+wbqyGBzgBL3vK7qfPnKlkCsJojd6tFPRGmUrZ9T6FYnvlzhEc2XDux/aqbJU
woPOqjxZ/SiTEBBazi5J+JpvCeYx/LC+Ri/3ognWtxbo7/VwsXQExiW+umx1UXQS
E5xhCRFgHXdIzQWhN9I6mG1YUfwe9HbXKXwaAAdrVYD0EHy//YC7SXGeQSLbjl94
zK+XcPtMQymjE8caCavbnhZaCMhxqmDtLKKXANmhhOFoRE18AwgNvtYHO/jqonok
/DB0XxWnF0p60+5jdYfbM5QabsDAVAO09vahh8sN3XDf3comyRH7IrlpNA/lKRT8
cgE2ga9yMSXN9OLoirCZeomBHQWLsB+WCl0bX83dqWwADqyRrL4EEZjwGjQvuT41
WsS+lV3aMISueL/UPC6s3zHOMJoSdMp1kXkxkrIYYIlRgQJRk2iXX2llQUNPNKkd
QYhHwKb3rJgDIf3wBBR82vHmzX8rnw/pa1qgTR5MqkNRDCVulntt3/oijBoXne73
eazm02rwZhHO7+69IYBUUom2+udQMJcnpOgcQNJjS44DUNbrzz/6dFj1dWWZBpgG
QZFmqFF/PTgzB6IBHV+wBazpyTy0y3uKV/0o8mUuGx5VrL6GpO7oBJYYKq8hAnPM
BFqyE1ZX5K6DOopoEeHkUjJ/0Y4H/DHIJ2t4F6K3xtQprJyIyCpPhZbg2PPEwFa1
I1nLe56xn4GQj2P52IQipCzz2RwbXgrlpxisGuHZWj1E7utE/eYpMRqksOBh8URr
6IgSoiXm7yzgaYfvVYmr9vIDQ+brs7G+OBFsq7MWY0xe6YOuo9/l0RUcT0LgPtP/
JQLGJmA95ZgA4mFUmFgIRnCyqvH/k/WuEnVU+yW6GFTPCjsAE7A9g68dIjUZFIjH
CHP+fybuh1GNscC3SlK2HU3sTZJMlj8JqHPQcBLABRADU1Bptjwako+fJ8uUsFXh
oSN8XoFCbQ6eF+vfvln2oVOKa6IVU3RzthHd/XFehAb2ldMShPFzsoDxX4crAspV
oUXXexxlLDlBflsAKQitVRNZkMTJ44h3/9jenA6sjFCTn+F7iBnfwZ+asCyoPrCz
BKRp/rPXf8q309+q9qA8t3S+mpwY25UBCDverv1qwn22UgKJeqjJ2/wKe3j6QJAo
Ck2OAhkgXA3lwLIBqRle76Z6ARdyDhOtf75ni5oSO9STDKUyaeBbvfkogDTtavZF
PnvmVR/4Nkrj0fn4BElCYMY6u3uj6Q9dFKflcnWroDWLwkYH2g2JKAAQei35GYtX
5eDCBTCOmzvLs5hdQ77ODlVeZrYG91XcHYxPQnbFZxWg/7Q8P7itXysp+dBSapgE
MQWdzB4UUUgQdJ2SC3a5pBXpXHY9YaLa5M4GMn5M/3vl8kCl5SLgEgIMZ9Cz1iOW
KMx5eivstHvOkGmt350cBhqTWPxLZ6uJ1UJeOM/YpX75L8SZjXoyebsvBmKC1O8v
iJG7vuUMF+dupQEn1Da4vL0R6QKUbprUlegWJdAkLsua0n2L0Fuk2Kd2estj/mEZ
Q0kzIOU09OASzIARmcMR/DW/t7EboGskYTHH20aTv9Mdf/lYuWFVprg6ebR9Vz5b
Zwg8INCU63Ak14whu1KXmDl3QNu8qYZjvNs6jGDJkGqhN/8t5Nn2h0N3PfqTgpRV
h6DgTI/IGUVs9upaSATYMTwHy7I0qbC+iSzBYaFQ6ocad51wX4TA6NE5L19sDmyE
QHCJ0AQT3vVsG3fVWBaWTleviajB1W4qxn8YBA1JKaw/jTApgqqUBtFWCgyx9CQq
ju/JAf4cXbrg5ZbbiHLPUAQdxq0wy1N8yKbrvuFyOvR7nyFe8GRqsrSQydrVbEVm
YqLwIfKPXknB2vUP8/l6DHA61SRk13z7T3eU5J2qvY3vzs9ajG/aVkmYndxOsXF0
7uHnSgPA72JzLw2SrlqAlgKs5LDG2B96xKzGPZmKJtbzqQPKP37UEeF8Ir1uVaUA
Q2jnKTkrRtgoTg9h5J9v4uguGBO1zSgeGsZaeenhTi8QUHfr7vr1L0q1Ik4cQFRP
yPqA9ztQOOWbarOrz8DwDE2M/EqTAD9sIzT8LGaF5tAbDVSGo/vhZ2flQ1G+C3oN
2JL/96XM17yQq1oCNpuHaglS4c0VNuaHneLqqD4SqfkPqtR+wliibycJg4zLwXfu
91X/N/YQ+6nSEk1QrDmb0rJNuTg5HjH8k+r33UpTRtiENcmqNOFFhx5V/FCuIJ2n
KnPqx2YyCsTmUXrGKfXFXcT2ueSuvPEyF7HCakFmdBQYYxPuEDtATiTjytyd0wbc
P+hC911Yvs40p+fEi6Y6htlqHkJqEJ11q1It+5n3Hg96CGNFDQJUgmpXqifi6ST4
4gyjWw8+OVfljPZbQhLwqChkb6LUn05yd73ho13AQ5Br96BbZ3U9vqhTx/QsXbF8
S7IzowEafzXGReLmpB1uZWn1ggBa/Cd0lr3vVh8xftoHrcZkveAUDIeNHUJ6Z+Be
OBdhSzr1MYDC3Gpg+3dxLr0XmAWo8xptip+/XR299rXkcaYTBbKrAci/7tfVCWu0
Ri+IK4MpiQR+y27EA5CD0rUQlsOA1GPHy2i+owWcNzvjsa0mnzVlmw9+8FW3LzYa
uFk05ftgwZnv1DtoDxL3axRgwbh7oNqjEKAyYhzVSiYYmchPJMZGOVQbCGx/Tq5r
el4h+eqiTaRF5x/DYoS/wClHGZU54ae5nFDHoXfwg5zqweohfzBzhbkWK5S3KplV
ik5fjGL1HT1HZ2K0hOotQ/Eg0PjFwk2EwchiXVE3w5PQ2935V9XicX2EH6k6Idus
pKMdlvyMC9hSR5BQKlbs5XX5kH9ytox7BmgpcaFZGWPdl6zySOdnJLwUoZVcIKG4
Zq55R2nWfHUqgndzJtIX1oOH8l1H4EZWoG/3XRsnKzpM0FpFd9YgYyl5gn+uJPbh
oAr5lJCxfbLrorQJTJ/oC9n0FvGcX+ADXVJWv2CwEFNtE4pNVSg7H+2bBOc0e5BV
8qkHgBbvWuAl/JhCoXWYChzp9lExfaw891nCPUQPTXQJEMLHTlYoj61U+vvbI0kn
0ZkNsdelL+hxIk0rR4Mn86ih3ecPAQE4479fuRVPbySDioPk0pHBRIUxHisyyeiQ
ncMf5H3J0upnSezcikT4B6OrMN1Qkf/yZaCWUsZxdQC6xk3Ha7lHys6O7L7TgPzY
bg1FQ/Lgc8mR2uegnquIaE8WauTvaJXfAi8ERtXAj2Va/E3TMDUSFtZUaXk4PKso
53mLBeH/e08jhKoExX0tYZPu1HIgaFFBmaGUN4uH25/CcbrqQa3PN1Htywt+7+u9
N0LN+uHK/Q807y+cFR9ZoY/kjxIBeoWWKnx1h1QVikhF0WQjOdzJCh1JDW2F+Blo
tZWVJdOwtIVH303F8ENX1lKFQGREoFyRltfBp2eSx9Z44jpkEjonDFW0Rn//R8B5
AQsOi3jaFn/OokwNoDdNBl/vY8cnsG93tCjkpVKfGuaeZpkeHT36XiUFViKJQvDc
0JBe2ruyvxYlrzb49L390ue7WIJAhICK0DANgC79APhYv6KEzZgNa85WpBYTZzCB
IoQ6nPPn1yWCI+Apaj2WnGnWHAWh2ojyegv3oaUYwMIuOvZ61ScASjD6qkn/zSc4
iBXzSDxmOMRFUvuevgLiqwAK4B2aNX+7qR3JYxlB3q1vW4laKscFvBA/lf9amr1F
Ak5qB3ICj+OYsEIsL4fYFClB9C5dOcKjMwwWtx1l431/8qT3KTZFGhqcz7HQXhYV
zT8TFS/7o4QI8SwcamYLC2cGgS1bpB42kTwJ1kxY65K9PUyavyd0N1r7gqbJF4jX
3Lcz2NHNTHRk66doo2xV8oANjaW+q/kipS0XRQlhB9ag7f0TMxNkP46/9r2FFSWZ
psEXRj0hfKKkKsgUADGbiduy4VnTqJUzhP5GCbzPuAqKugAYZUt18opbg3fsN8GN
Y8wKskVBXjWwbbWuKWsyDMWSYtvihWbBitJAHqefWUSNwSZdJiMsAMCc9cEhb9Et
n18Ct6JP4IL+sSaaHTkIOFFqPSqqVJGj79yX68uDbYLyM9RRslKzZ3qD56ZEyLTV
ddyf9hnmZEv2zOEgiwojbzfjB0l2w1AKNrv0q1E0g3NYTgBkQW8gsDXTzpAnyzZc
/KatdoiDTUMfNuxceuQL+lKAhll4FHJ3AL5g23k/JWzD8BU7SEUGtVkOxr4UgTJV
a9xZub5xpM5rXXV6Clopm+P4/mXzmXWhTI3433inPNJ5uB44XHtb5o1ELhc2H54T
p9B+snwbT4KD/h2v/RKLEL92oCJpA7HtzfBdETYOd90nQe+WuBkvirx+3IBHWG3G
s/Dh7B5Cw7J+hCJdShglemJ1Q88PC7V8w8xUkFuvyJ1+qZItT81mCpsjHBQNXO8e
RhQyjlvJgaeIBORDeQ/Fyv2TrG2ev1xfkTx8Gc/+9uGwSfg1bYWmWe3mAGnil6vK
7LpVrGMQJGi5yMj6PJfkKqlfcPhn9bMii1lLC0Tdf8jMKtJjcy0kRvVRTy+u4DTg
5Wvd0kxgYQRe/pVBVrXwKVMRXCk2Gkb8bCbKL0W8Mkq0KUNLHwOPrBccJVVLu3jF
WfXY1C3YqX3kSc77ZxFy5y8ybXTDAQSDQgL2qczhu5EGOFd86bts8DQfx9VQc365
c6YEhqvG0W6Q8tneObRBs/KxUXVAhhJP6zlyIyV9mQxa8JyxfamPQioL/GxvvQKl
ghMd9Ewrx/F/7CR+LJhNjNISIDlbrNE4nAafcwXui5F6NFKaYe7/hCEoH0aX+1jH
0mhtP8LiuPG7AiOtGHvyD4HI5D1jrboJThwfKLDm0jJru3RHBwix4+m68D31eoLS
pKirSxlncRBo0B7PUFqBKpqOYKlX8BJSPBLyjIi6GFo8Bp3r77OFbFJ4UoaaPgtf
XmUfgbCctrJboheoFOVkdG0d2K/43wGiOGZrDZNuIb4WAmw7m9TwysjCtygPAbUo
57t80X6X5LrvbL4wRpPBCJWN/X0mFm+ZuquvfYs3+GnBpYnih36hNeVdfMq6TKQH
AnGLVvgPLZnhRntEfu4mJJqdt2hys666mmpuCTjXXQBxvEOTcTEqQlIvtONLwc+e
dSAanB2oFBQzmXixz3hBxfHuMiqzSr6sdnXK4iA1B7cBfx1lobGjFsmp/gC7zlUX
YADzv+yH1E07Iin35jYaUxQK6PmwtZwEmNd7BmHzh+GFYThGRyO0GuibPkkMI+C2
1WpJO7PH3GQRCtEpNgeGsN0sGoJPRYp/5cuY1mFguIA5HFKKgDoWXvFazPw9J4oQ
Bv54xOVhQ0ZKgo5aOIxq+bWHA1BUu2vJs3EB8zU/ZyI+nnYyhW9KBW2AIzEZyefL
d1gZ0EWWt2P26nkC+btcaL+bZm2y87TcgBw9l1eXCiI8PkJ7tZl0S5cme7F/y275
LTwf0OOYDyngIQkYWHh3edjfriqvabxSsBDnQ6gbE1okPmZcl8y+/BwRo0nVTt+l
KzZ/iWX6bII+VZ991hNE0XyXFlwKTc7bYuscpsiCSF02ImYkDEJEfeXpkyKIyi1A
HLDLKfzKRxQYF6zsonrgO8LxFIImsTQ5c7iv3LpDiTfwxlGnTVSshpP/OwWStwJG
pADRA7wpJMNUb1yvnGkl83+arKpvSoXq07NseITlp4aQDFaYP5fp3G8sKRSBSXFN
B1TQZwvGtA9mxziYdhCajBiSmBKnuTXXtZb3B4b9ogRsOXqr/2fD1z5zTqCU6lFu
DINOhJxp5Qh+cXD5xudQmxg0lLRdnhP8fUIPcIKJYuWoC0xCXqmfASUOrTvFGrl4
z/ZVKq0Cj47/TgLo5PdtM21evBxnk4MrfC6T/IUWPw4IIpb+ahbdU9NGxK2YounY
y7NSZOPMAGJrVJvQnKzokYksE+qKmb2xm08mp8MjEwojiCl3v+ow3+a27D+MSS9T
4sz0YyaIju5k8ak3LrRJdc6eC7JtY2VJ0UiMkTyfkEf7lEUlh3lQVdLK/DV6/w1P
f1nwrMES5KQR3FwTvKxC+mMyIRfkzjcnynSzllCp5WZ8nFmJv3H+ZNYrF8/5Cm1y
n+ZFOXL9HH9NjPep4KcXt/MdmTSdlB8QZZ81tRJD/oBFD46W/d8E9svNVsQSr92m
z5VIRdCxhwxu5Jak9oXxnAPonZwXegsXYc5/54s8IGWUhDjM7afTNGg5r7T1Amuv
ThbQ7gQ1RFY3iHF1oPNkJrMGWmwjrEN60+MfsnwdlsWOS1J3ksPGFh6xQq6N9NTc
npTDFVWr0mZahvXIfuGp3NyPPPHN02vBK3DIc12hgIogWiOkRf40+W+MZOOjcc3N
zYVj+eoP3nqU9s+EauTY9bz5XI71y/QA+JjdO+1/VVplg0pgTHESrqcbDK9q2PX6
UnaDx+kHhOuKZc/JrkwwhBJ9PQQD86ztCyj4yOvPbdYmHTINL6Noa07jipshT+Ht
TaZrMj44Ar5bID4EzYp0wNjWIsYymRR5X4oz4qjP7xKbNv1pxOPxP0UrYqYXRB01
vKHeIb+uXxrjSt6BCAphcWEPj+A5olLyYRHcoQTZNJrnRuSUy8j2zvbAvFfLiNJZ
r7l+UwPKWluR4PKx/rMH4lkLtKThavRRojDUYmooDaEkMFg73xfCHh5UeF06t+Sf
g+VfMZIA5bNjAlyFD8EAHVp4ncGQyJO4V69Mlv7IjIQ2CD7kOqozxZhCmK8wUP2G
Lvr8GUUqT8s/A364Rhtj6gK4TMYeUvtVlzN7/oe/cXeFDxQthCELrtZGCR2Eotre
fvGZyqLSIhJJAdjraLDu/eMEgwp5aZw4e/8YdaqU24HLtEmU+cvLzPq7PL1FAi5d
iJSwzr+S7xjPH/wRT7LPABGPg08CBrD30w9CvmDV3t5dHKSmBZBxM+8bZnK7AunJ
b3fRUiZJF7K3B5Yxo9eXxpJhMCYP1MVp1wE5BxUDzZIT6V4mhQjKaMwUD36F3u7n
YlVVgGUnxjGPvDzNzzl8h/fw0yNv8U74w7PY3bIuYeV/4Y5QhZLdd/Qxcgj5/GcH
Je3mJtddTmtOcVObHJkx5kUko4rP8VWCOx44RKxtWuSNmbXcOH2lsxqvFzgHik/h
pydKdfyy7Q3K14h57bOxnnzE7OF1YAL3FrGGbiyACqsiuNTTz6wkIzjTAFYYBWvi
HVIw5+gm69Kio6oA5WGSMd6T8DsCioaQmQ1m4TIWHrA6j0/4G6+Ytnw9XDQMfvB/
q43PnOgxRiFK/MSANI/p7PaESOiuhbBZBEtYWej/KD4EFliMEkFNEm7K994v/U+X
BCBaWpRlTPpL4IpDGKpgWrYtWJshCK651bFIwjj1za23+oCwk2cAV+HuE5CzGymv
Ae7jnxx6UbCYpyU0JHLPxeb1X/knDTSbKphXiZi02OBolRmahMKfg9vMwarauG7w
iQIWgxg6GgX09HmSTJL0wllEGNLRQbJ2vKsKR7ApfYwiDe8ZSaaJfCOeAS3lbEbM
jx29IAIsAKtvDepFSbt2YoVU3mwBFhV83NsZyICWAsDnjKbmuSw3KUQIAAVg4tf8
hxYBx/dkS8yoXmTofwcDta0bMe/38lJOnCmfSedChseT4Qt2WUMKeGqHXpzg3cIp
UPncKWaEmWi/HvDNHu1vHVuJAvBMJii/1nwNiQN3L6sMjvsIE4XKQQ4QVo/b9kU7
2X2TWwV9IUzjabcqZgYqKFZ7ILjZATNFrwUTpptv3bSR1tBxxQXuhL+cqVVNh3ne
ycBoUrjkTkM4OoFxTS5VJcr5ValfnonQOTE+RgfFZtmVWyx/mIIYESKG8gD4Ub+t
kM7Ssa+OTYnti+5kzJeR/9V8KCQQgfZJJ4nBsTNCZRZVBPoGJAuMJhZuoLN11xpu
Yt7Bd8kZfqGXu8b1oOGlGHMJGDI2gDbVPIMRpEk5ssjrdwzE/gGkM9A1pOqbAbdg
a/HbtPQu7MCz0yK7If9yOGiN2yhkZZWMCVVCAMulwvbja5kQBvfmS23s/oO/rUpD
Qf1tsraskQ9uCW5wqwgFkbcUIkozNlkbqnn4WQ3+/vSqdFq1HmXEeibkW9ecudFu
8Sbjs76AqBQAzSkt8FcUY9eFbuR9WV16ofMm395nE1ehwRuNCDiHNApMOUuLPlRf
YFoq7vFBlzg46VAEtGOgeZwQrFpH46Lbi9RzaZdq2CwoS8Je1RUGiomwK8N0lZHy
vVIsIG/ARrHVjP3lHmYkbBCWeq2wV3Z7mZogfy1uPAzCXbh7i8EGossBtaDrMOLY
COjcOmNv12iQ+WJq8neKn7UHGg7Vn2KIb2huL7mnPbkCT7CWQe1qkVNUkVK+ZNau
Qnaq24eFCGruRCxMdZNKnYyeWceWI5T4DARkQGmRPoNC6v3yzZ7bG9U3QFJLhIgT
QQjkA/aRZ9VPVHj1VXuZASEaXCU/yKavRwb3goxo70JkSmucS5e9Q+37ivAMpB6j
8m+laFqz27zEryZqyse41cwgp9sykKKKraUOX6Vhi/mUbP8WjFpDCeSeDf7U/VbP
wXb0EnV8St46BJVUsDfyvruR+vWeVlWMVLZmTuFOrE7WUNE32oSjrLHxp+9nRx42
i8p+JBzDpFoNLv4XNEwhNJriBoAxPW01yxaqMrt+9xhOebfvEUq2cHxubRHDkzbH
Qcy39SNowIuLauWycZwm05561V3XR4o3cTZjmUbPRACSDM3m/e8To8+43DgH+KNo
2yEoa7dJ8Do6AMZV/DrtEMQJ2nw86jn6qpkLG3S6pruqFzbqCR09qQ1JihVdt2Ot
qphc4CbW4Gt0Zclc5gSTMcrWy7YaioqrbS0B+pUOAgbFc/f6PM0WMOa/HYrnMA42
Kbsnud6fZI6OWbB5bkmIOHCEv8V+yaaqdCaLpk8qvobv9qDeUG2eYmMfIlXvlRtO
H7IxT//tF0rWC08QrEIHW8e6CBa0XmXalTE5vAiaKMfkxOEFF8EpH0KR47CGj85m
3CDENDY56qPQyAT1jzyB3Pko/7VhoF/yNCcqKdNWJth1eqK9XgRM3FGvskB7Z5+2
5GkUQh+wydbLiq/W38MlMzDQtiW9Qi++MzjdnCHaKiqdUiR7DrqWDioIoWq97/HX
THfFOErY8mzYMkcqrcDo4ZWDmewa8NYsTiZCrM3I7rqDZ2PfgAu7ikfraZRani/I
wuLjzFCDb9bvfxf+8edBHeln2HaC0v4i5oTJGIuUMAY0285uzVONUh7UfYv8rRYK
8y/9OZHFWcd+hbmnJ8pbpMGe7T2dwq8nx/EE2HpR0PjA2LZIvED2DenZmO3QLC7y
tV66shhHrguyvX6sYRhg6LdsH+eOQIBGvO/9Uc9ADY7LsU0SUOZwqkE/6h/sAL41
3Kb82n+Ul8xBrpCxlELYVobSP2HAAA5VVgkKFMfqZqiYjiPl7j0vf+GHS3NsnWXM
/MXBZORu6HZLQdNXZQx0xngMcsQbeEM27ngoYHFfp8iB4kWUSKHUwLQ1OvabWQA/
RT7MQsIPmP3Nyc8uqrPLHtFBdzL80XME1zm9qfIFnrFItU7fPWeUWVweT0l/dfyo
r+ky2j1sr0ND1LExBLmyT1uHcgRrDYEgv+VwaxhVv+JfCiVHv8LosQDItjyS49os
kiqcpF+AUtO26NXcj0rBjUXeVsKIdnUpj+Cae5tl9IFvQ/uuFkv10xb3HE0HO9lI
a/UssEhG8s2xkhlyEejcKdBPdru7oWdSDvrmyBwmA2dvVtEWNmFxL1OnTT4Tv9tB
ffqjAflE5h89JdfNUYsfLEnhjQs31/QF0s/mKVhDwReqyCMXyN1NYGmAQcf59fcW
tHerTF86vSkv6HEcPGokoJQtC0JBlpBJcGmZYzVZqgmu8AJ2T37bcqBSXwGGudg5
h1oagz0dZP2gymxL0cGzItrR20ZKc4udlLHFPWQC+QsHtH6EtiCu1acfd8Peylsr
5Rkmn59NmMoxEzc+UrvThH3H0fd618r3g5phH8VAULw8S35hRNIAFy4rI1Kmj5MD
9WRQgQxfts+I7UeymsK6HQ5NOCuXEy03/OONP9b7Y0rYgmSTsPSL4NKAbMaCq9ll
wlzK0Q83Q73emUE1jfBO98nb1Rr5/LNMdeUFIE3pvcdE0+PACAHN3nxuuZZ6lV6C
sNKwvXD/OwHD4P/Rl8tw4opiqzvCS/Q6CWQQMBB17afIZj6vguWX4Ko4qbg4+c6L
gY068YCXuS+9VRYhTSkvdc/RRAb6nQkAO5ZI4WDkkhWFFAlXA8A407Ik/8fU/pvV
EBg3ju0raOmgtKrZ7P77a48RufQvpQ6/ADBAJboIHJEXCNkuRYkEF/XCXhYkEiUY
V1tC74a3JCuDMVa27gnm9hKWqGmGLBnyrSwsddlt79qRH8d9DL59htMSFvMFNd8N
FdYYPDE5MQQbI5u1iy0qDQX2cAzC0LT+bSYoakKux0Bmr5IGbmn4gi4VdxYiAzh7
g525dkNAGHDAsFD9UN54XeEGIRULtVhrldV1hN0MR/UuyZmZbg4DeLOmKHe+Wl7J
FNr3KDx0MbUL3fs9u0uKA3J853dPXGnh8eBWH4OQuK0eB4qac6LIx7ZROiBESQPr
1W8ltJnw/YlMd+TBcrdEYeoayP+GZtJfXr/04cRKdrEtim74ONDdw7JSXHCObkCd
7tgnfeeR+tEYLNUFFr/wb+QMVHzO6meU8fIshHacXkJo/bVZPuatEwh/ZlfClxSs
tAz2tDSgf2AMlmoo4a2TliIxOQxN5pZJ0tSCS3odvv8oN2SZOVf2tTKE96Jano7N
Q1uDcf1p3TQtICadbKc+zRIKxavMaCKsYqTuz3Dg5HMQaXJJZtCyEf0Pw8YtqUAo
c4RJj1jR90H9gAINCBE4ipPr781FD+ga8HAPe0/wLkwhJ6Lvo3iDa7RhG2oH55So
xf69+Sst6xQm3HHWrJJTcQoVQZZDomPiorvAuUSK8ZejXGj42RS64zsWmftb/5ui
QROCCIvB0MHiOqW9huMDP2uewPrn1/2i5duHraAnHiXYsL8SiNiE/df5fB3ea8va
cBWpdZF/sLnuBA9XcAFrmXnsyIoTNa29xZsWcn0OWyozSFr4E4l5vkr42erblFYM
yJuQd1w6l7sVCbbqfTfPDaUdvFu+nRo6ZgVYWhbwVb9W9+1ZCfH6nWE7VsE7knAX
EUSiMkvbOVcAgfHNTu7FauMVYLrIZjMX+uVHWsu4vOXjde/2ZwLZVKUh9eKbT86Y
RXMXNQ8YD2z4ElciSyN1zmnVecvT862wRX2n/9PsF+sfN0abNjNrPWqqnSBUyN5A
F0KO8TigfwZQTr9lJwBlkPfmLLq8W2g6jep4s6Rx9skY7w+FR3cL82nVFUPEdRoj
t82GaeAYDkozYV/pusVWigCpDtoNjfhgCcV8imr5Q5OLNuUNaNzUZKhoQB+rGSmN
nsk/I5tfVWi/hs59HFap/GJmykmSy8epNH7PVx4kiaWPH0u8VjIZNDaP/m3U0dz8
ghlyEe9mA0matIWE4ytivnZnXN0Z64j1ZZm5zXlwwiM9KcF2FXWmOwBo1ARA2QAb
YnAYPIzV23jbisHS6RyDAIQXGYi+5ZQ5FSi1ax6YoQ8elkYJPXriQ0QN0nDAu1Uj
RybglppdHIoCacZXppKezNzk52QIZHPNG2+0x2nq8PQVmxUgtkmnKnY3jvw8+a++
hYwsrrczhUHZHwrz6DmnYkRlDzVfDFr/M+WfC6AKYdOUzOxbVNkNNqi2JkPpmwBv
kKJPqXlRhRqNugUmubg+Jbw3sEef1ThpbG8MU7+TfFwuC6/sjdccqOUofmghpOHY
NrqPUFkiA+863JBc5Q6tIuXNI02GslvTTIk2QeyFbL8JPzN4ROYiX55NREkaQWyn
yflierEx6ieTTD0RdDQxvM0AoURIB8OI1/Wrb3L6TvUHU/Jnr/l/ByWSp63nQ8rl
grh+wSEhf4NaLpZMYDackWAOANleGO2MF6lTqMygceszlhNrBv/JFFrxsLZ7FyiS
DBs16Gutvf+0T030n26kylyUtw3OVZ+9qsZ+aJyCriVo3aBVq5Gvwbf3zF3Edi7d
vRqRBrlNC9D8SyUnPtaPIYvWip+4rMQEuvejaCBnfKRsvvQp9UNMhHlDmYoi15zJ
lqhaualofw/RjFntB53LVeM1J6VicDgJvTnMJp+0fcZnE/UO0EckX8+VY+ZLWTFi
KR/bvzQl0jgkC4HJpTEn9859gaI8eh2kUCL01bI7BXziw4foArjMXA9BTRdrdfLA
HIp1rGBV2ORJBCaMIMcZ8VBhualIcTLejW2bJESXK7R275dBW6H/vqOhxZXEqFx6
li4CLDPZDNh7YribHdS0Xw0qaogGJKg+1lWW6TLkzwmqsfkJXtx33QWHB95OLebG
YhAvZJ4+4a66DbUoVDMy/P2Io8MuDZT+H6wP8m2Pp4rrA60M6EUFR/82D5FMbetK
hdt8zvLcp0bwiD2b9W24I+7JUXIUuuKXbpXOfY3s3q6DTdwP8VamuAuG5imFzAGA
YRXb5NjR63NqdZwrLD4npSBJQn3p8Oe5dY8+dsk5hQTYsjhc7v4bqNsibPuWGf7W
5NADMvxK35TW2wCw5s+jsrpfc3LCTyZN5R3Jez46YDATLDgme8U1f34ZPeAlNXDL
DjZJlBXUtNeyn/42ortrXdIB3Ca4RfMyTdhBdcChU9a4vloZhqMvqZXQl/4n+UQy
TZ5h7ry0k9z7ZAMU1pPV7s4HQSvVCd5Jg9fnFV5ARTGnJ7nOt4q0oWF3UOJxV+/c
CTMFKE9tLWfxbTV9RGc3Mg4yxfyfNv3Soc2moCGoKEn+2SXiApee1uvZycBW3p2Z
jkLV8dAbRh0y38ycjYu36G8f08WHsJjzTguA2uBrs59D0kafqLG2r1rLpEfXmYkf
PmbwNW7Blbm949KPw51dvXbWiaynucshRYZqWKozadn8h1exZfUtxWXojUdEOnaM
5AKQcGDbFVztjbGqmuNt3DG3hSe7HoT/1PtSinWCyzVzsUfvdlub1PvAlS3fDwk8
UEC17f51P4gIC9XtuRHIXE9nqzQpx0j/VIWMqrggkifWJ+inLY2uIbVPLYisRvPJ
qtgENz9+5tDDfqA8Tz37aw9UvB4xiTworCfx7WjmmtBMQZj6qpKjnNhTMZTzE+dE
JtQUqg4bIf3j8ebJBS9frum8jk/yPENt6H37rAAq67iUr11wa/LbJURW3dh5puyg
3bR4W83ut5CbsdcIGYoGDyeuVwgtRSBcxqbRPG49riYGhUf2cOJUiPwyEDblMyYn
xaILnlETbBRODnRwgNNf1j6LUTohs7gkkdHppZwvVQN+S1qrgCkLx828EHafIjLR
6UJ1XeCX9HI8c4f/EtwwO1Kox3uxVES6bgyhhnBHOlMSv2EBgfzU8u/DGbAXrLkH
/y7+6Cm/V5FZUglF2axHd7vHsPoMMOkRiR9HiOQflZL3GNEZmySLjv4qqIeWwVXW
/7ClDYppCJD9/4yoGqEKsPE+RWoWqi4cDyE2HNrLWqZScePyWfTNZcrZ6hWGLU4c
sdGLVrkmuZ4m6zX5ukc/JRu7ZcctiZ82bEyILzwPMkGJhnmJmhoH5v8zIJHV6Ywl
PSeI22g8Y4iTfvgGINCYG8NitmhcwIgx80plW27uiLWMqDO/3zZTDSIV/ny83urV
2jiBV8+L8LELAuyGXeIE4Nc1f3pLdPGFx8zrflF2M2BPNGyBV4a1y7nC/FxDwpj/
7Ae+GrJ8tugsFl7lwjqQWhd/Ob6n7AF1MywfVNLLRy6mtph9NLdKOnuqytYZTDoT
sRlAdYn/EEUaixVSn7uqiePTbfYOIlQDSdM/XOw/r9q8oCMvNl/kosdtcVWHEJh7
0nKcm9cF69lA3XEjHXOrD1tpUqItH+yCxZO4ZIooOr+ctsIdtGFFLB06aIDeUL8b
gcL08a5Ijawp+0RxN9vHsolZNun+nbfqU6y5cFVGhemDC1vWLFm7qYm6CI5kNT7j
pcvsP3fqxhrMvdB8F7MqYEEF1XAof7aIVyFF+xFN4aU+lg7nbKk0zDxjzfrmxRYo
pFvlQsVmQEtFBx1GdDPqRJ8Qf17U/K2vNSRZfAnAXHAdx7nt6cqQgj/6IYyP/x3x
s5zlxjSJoP+ZpmAkm28ifYOKw/TIj6v8QDPchz3ALxCaSfh2iHF155CR5SB4p9vq
JLGeQSlHiGT5AkBrVlNB6tldEUHYoKXrUV+QoqE6jHLD8AVTUkByMBIBbU9CgGGQ
gw1IM8py/vL56ExvcLfXPq0hS/mKGFdQMlbEJ3oC9o6DqKIg0bcirIfro1+mg/nh
M55ul+juetH58uE0WJPsAsV0PDkXib/mdoz3toDl+gGcHOTbk++921dOvG8R3lCv
xkWnaDt3k66K126l0wQqRr1YQSb/PivXK+xVnqUSAwhrs9aMxqU7+OkSK7D8afyB
5/rN0XNDUh1o9RUgVBTP+5B8R9eDTm6B1vj5PT6JNrYXfk42Gav4fagSkieOOz6z
cmBFskpJhA23haETls6fj0f/zVmpfVOBwBMXhugg7g68btwOmFiLufcn+ta5I8GY
c3sdbJ+y5osjMTxhiX6j3cb1h2hGVQ6/DXDbS8OWpGsQOkmy4SU+N2XUgyMf9yrE
bAGi0F+ZndSvOvn1KiRoZ3y3joEwqhqH2O0Xs5XYb3MRSoW7btaTr8VSjtnB+Mue
KdhmM3eUZC34KrGZXoBiPeEH1Dp31RJK0Rv/1rqBKuH+yaw0GsaeZmy36DMtB4Zy
2FenJjFLnLb3HTo6cd2xcsXxbcqJw7m5NHSar9e3Q/wS5BbyKR5oqCR5SS245q1i
UC1CqNggHOJIkKFa7m9mDdBeKIPY0FEQi9kf59SaD2XJp/6MfBBl3reLLxgekUJn
OcIfGhFCoY10e6Ly04x+EDMOvYhXcMiN7NO5nWPDVkPfmYPJUThj6M2b00m+9ZN/
GUYzyFDmJzCpEQW/bFFW6+7sAY9PM6lJCFI7/irfazUjwvibmtonjRLjFuOSMxMR
xzOUslTqKShgg5VnrVmfRdMCnCbcnFBSffm6Jnbixu+NQtuLVFhL0Bzegm1NZdan
HjTDIWYzsn9dym58vV4nGul/9TwzgDOmOh9IjbDWV9Uxh6W5/sR0ue/hL39tpsP6
bbNzHpiTBg+CRbbPaQzlJHsbL+sLF9eAvY7zVJXo1PnbdQ5xlS+vMUudsnEA18Q/
EXMmLz8kBovB0gMOwSbkdN9s6FN4KQHBQB8TEQDSIw6f0dA6dBCtYI/b6d6fct7P
efgI3WjCsHTF0fL4ULwxyJgNOY0YEWhGm9L7PvpfySutVaagqyACMEEV9jbL08sU
vyZW3dZLVVVRtMHeQrsg98rWDZRP4DNxdId8sfKv3IyAkmVD+L+Yw0rwC2R0an7j
E5zZ70T2OJRloNST7XHvyA3lPSzip7/Lovasob+27qFhEt+IENKS3spWGXfqAHeD
FvE9H/1b8Vsi5NgMXbIVjMxMPXJ4NeZq/dnu66/V8pVdEW1lUxcobcKA7nA2rsrh
pRWK9WQWuFwf/lseIvGrYmHg28MxXV7neOXfMi6VKmK0Gk7CLHRzhHYTcW2zXFCw
fhMbU0OTj/oCoO0dPj4a/zMWb8V8P0aeB9SWDU/8y9R2apO2uTDGQD7UxPmSX4ZR
h+Za71Hb49971h/sFYNeaIPUloBT8kHo4cPOTFyD+It07lIfA/lzjfZ6jeAKs6G3
Xi1/E2c/A3D54EIzim/7Oa/DtGTqE2cPZHiUbY7GsA5yiSKRKe/B949jC9uSQhu6
jNyK3dN8GHzPjYoZndsdMLXYu9I+VTOhRupPTg0ihbNdliL+aPceg4CKvBZpiqE4
TT0QXBBVZFK25nu37NXMcmFnh99QlVIKedX9ERTX0kkAQ8KCPnqPyoARroFZaeKu
K49e9ufHKqsRwlf37WFZLb0gWAohtjqJJISJdeF7+1FbCGFUAX218fpPejNn33fx
MMqCX4XaIXt4W1Yxr2+hKZGGMUtSi6geufTvO+Fs8PFCc8l4+dPW1AqAyvIBfIW+
rY7VkEFJLBfKHXDBU5OCM7KacS/HQT6h2PtbT4cEmbHQdJelEnp+5BR84JvXh2h3
t6n2ARdQjhcK8jG9h4uRMGIAPujZVcQICUL1mT3+4S+mFKMoamGsy/veUCr1NV4k
Y+c64R9UyLEkZXcSDES+Hn93MGjAV1jYXDrjwZ+dZ0tW0steUpVSzNBakzdI0ZZq
/wNviFlPMZyFxCoUEpyJoTBZZJIWrOaYeP5QzWgZaNt1ps4wRDb2pnKxgZX8y9o2
O77qiVaXiL66WKjy4X4cDfaDdVRmnY0VgRh/8T5DcyDPFNMBRk873qkj9/FegLhZ
0pyMoGOP26gsMLTTUAtHPd/hr1lPa8IvbX7LJWNgAGCs5ujgafDmNxOv0P26iiW8
9LIxOQ3zpBbxan1NP6tlDR9genXGHhPy/Z3DGVTakxAYrB2iCTJ0LErY3F4CJg3x
PUjiL0HJa/wZBx9gQeE50RkzF+scsYW/XUR0LkshL9XuTDkIimf2c0tlFITlBYZi
NXivJ4brU9/kvSVG8V+8uPqnppAzOg8FSeVgjb4O5bLvP49uZDsC6Rwhpb07r4Y2
OpZhklVJR+8gTV85noaCp3qq4SeFHFew5YZbRFRPlwrFcHAKoLk+D0WCmpskmwBE
7XyEJ7xKSNw7AlzeONp/hiLlQQD+KD/42XQlN+QZgNi4G3HiA9z6U1QTqdLJhNNi
S/pW9NGXccLn5KZPPMTtl/xCLu6kDo+OgG2Frh03mW7Nr3W5uVM8tlPoGaS8OL3c
2TXd2eWuAfSqydv+A2jxax4twFbDwvap3JMCBB/SKLyQQHeW6/NyM5SKo8De5bI8
SueUskx23Pr6gMwsLZeGqKXOwxbpP6b3OFHv6pf4ZBLojWldfYcZgA8wNlzxOMIR
GVutRjT+wXaVyC4z2CNVJ5EkMojHqZRqjBDcB8ZqUpM+QcOBd8HB8xlymUcYfHcl
sstQQNFQ1GntQq/d/XOgvCwdNnBxKsnGEKiOdvnqRaKH/m/QFnbU4G2BGhjORn/8
j4sVE0P4XHXSD2hTZpsyu1edyZZ/n0hlTG3uDi0JK8sGcR3GNH4t3hG1VoYVBJ5/
RBol05U6nLgfHcAeBcnE0xDtjYAiKVB/lFhQCPcrzTtpVF+RBbW8YFw9iRgLMl18
mw0BBL0H4fKQ7NYlx6YjbX3A52hhWf0KlwImeXDa8wW7Q7bR+snD5e0+Of2aXkyd
c3iNGnio2pEnl884ZRLtuL442m7LFEQ9p1t3cRCUJZGEAXsI1S/7Iqv74lumyFQd
jA2ooYLQDDSYltBGWGVO3NH7vJ1b6b0LKyzt0G9Supy7ln/+SAUEXUWQIG9xsCCX
vhRaO5OLqI+a6a0X/MTtI37XiSWrKX04EtNL+pFLiQDs1y1eYT6TNeXJeNNRrxs3
2Ypuw9dCFpvY8V/zTjaG3/HsluVMtmvGGX+fkdbVBaaYizLWXYx0wjKQgzoTM+mQ
J/+PQf6xE/YkGoZN4GDGRWZchjbA81EuoUH0WcYtJTOn6mZJ+Bk9XIFDyz5vQJiv
Ud89MFQaRwFQ/xznfkffGjaExatanuZ0R8VqWNjrF94haiIQF+QjWZAlPQ9ceCRr
XzjZ3DzbsZubh+virOZJdFJBjxAdM63oC5Mw7Bz2gNDwOr0/qM7W7HJRnK3wckh3
jRDRcjy+5n2lXVlUDOXtWlxRKflZ598ym3Se9DvBE/M3SP+nUHXrWCX4LXcexAhq
uUoQukRrr2N7RqA0rTo9XUJdWcjZJvXiVz4uPAWn/ieZfH2+Rd9gztq8U77pge58
ZWIvzur/wLUCN6jl20x53sWH5ipFIwOgapqu1uGrWwfdPTMiJ+B9LYq1lIWPRqyI
R+GreaP7rs4SnseJ1ULfSznNkS8NJQoSArLqEtOF4wLR3J5zeixPcltc1ezQHdB8
2VysfMnLTy5YcuJQI3FDmMk/iA/nm2M3FB4GSNOWm54JKJ8qTj1BiTCclBCfMSMR
kIjMsoFwJgF62Hta2AZ054n1Ug2xnhKhJ57Y253I+u2kYsZko7P6Mv9W/Li5xEwi
2fFWV/MVV/uxiIVcDRoF2foKFQ4BL53G5y49jjszqht6a0SLK1mkUQ7N3835Xt4p
IG9/aYAGfLnTIYSszVqQodpoEBnSsNWuQxrOD7yjM789tCFYgUww6WYRe2HWaPO5
ITcYm/u+rb7CWW/rC3StHrwi3z358ljP+fYvBHVyvJCO2SZ7yyfnt88L69VpDTNL
RaL7uq9tjPXufY3zHdvV7I06aWdXOmFrNhYgttuXsKLyx+cK4ChHjNr8w6evdy48
oGyaBboKpZi5uAMRa4gl32OFh/9d40eV7vRrUDGIEK9jn11o7tIJ4+jhj0TLFRjp
BZlkRjM/57/bHeFX897mWEZrPQSqLLWmUVWYri8GPtX0u6sc4V1GceA7PEJQrR5m
d5Yx5NSP848z/e9xiaBT3q9GIuTHeBPfmzn6axsiVqZApE5XVKBa5uksTV8+qN5c
OXyxC1fY08I0Sj0UGD9Vt6iPCI2292AR45GOBeriHqTXI9uHoMHfKnDRaN+Jdz9P
Vbcwy/ueGQV83xK43HUaNQSG8afwB7MCoRQbM/HBW0SP9HXI+c9eXMPDaK305rxj
9wfEqathF8ooNGIKFxCfBuU5Khavr0uJe/NRWYegcYAkQjBT6rajJtoKiVj35TPv
D6wni2We0JUeEp6aqNsynwwhJ04Wr62n7nfuz6sU7ahh2FDaik/C7fqTq/Vw2IEX
dCxp+oByKas9fk8nBc7MdFsOWhnmpPyyIZbcSg6is01QYbHjWjGj+a/uFG8NQyIe
TYweuE32weW2zOJ7IEPwg7Rfd4cDFFOooYB5c5X19O4lw+AIGcy9VSCXPdJleoDk
PY6wlX2G4qefh3aajCCI/dejdaQKjy3pp/3BGrQGTbLjNZLfA9kofnhq5W9SLXhN
fv/8Sen4wWdMybFosIWKWiDFmF2rziwKItwa7nYN4STfV/i2Vhgh49F3ygCISep1
30Cy5UhWC9WRcoZ9H95BaQkbOI/DpZ6X9GiwLcsvDeyKp45pWI+VM5/9ukZRiw52
8KzCHlcgHaNGu6WGMx9R50CWPLN8fsblX5ebFJy9OlIRE670g61b6LnyRXEr5ylr
jReiXs4AtAt2PYPm5ShsfFvl+PaZ4LztK1OaIfIJFQMCd+RKhM6FzlleuJPFTXnV
IKnme610igE0iDKL2FvNeiqebMCoWKRD3OQ326bm1kfyLG26/sAp6gXdHpChXjgR
0szSMRKnk0+SYDlrFyOi/ko9VJyvQydd600aq5UNmQYbhMvgPty2PMHy7x9wMRyV
xZIeJ+BUKpINt7PMfCDCzJTgi06xXzer/FdPePle/ZFA+IGTwkxrmbaY1BsgzYFi
zSy1dZY32tyrzdKuS2hm7OvMmyNOL4YC29DOFb/w4XLdsYAjtBFHbFE9oRlZo8u9
BPQc1w31tn8hhRA4ybr1lI1YTHAymlU91v6wH588/m1mdPXSp6faHTKI9ip5JycI
Zw5CU+vLH1rKo3AEN8QNRHKpCUOprk8Te8upNVmxfdVLsTo0Y3GNtv3+Ilq9pb25
5lzFkv45Ns3UVaSifFFRxXiiBRr+L1vtH+QhrnMQSaTM1iqTAWcstJD02XoQDZUO
fe6mVR0liqRRuacSk4fz2zmu/TyiUe+mIUR2lnTvg4+AqbZ/Iw8Mzq8oHN9vGwqC
p9PuUyhgL+oXrsLd1wt2H5aYSa7rvP8iQPYXNdxo1jnzcx7XU7f7W0a2MB6EwhcV
+FoJOW3A6xP9EkKr0i8MGNJDzz35oD3yKNAZXEXIG9YA4eSwQkpBn5Qvs0D1TQ7i
IAG/d4g+gVcJpi2PREWyXauw3GVSGWtZ8MTh4oC6tQ1pgIvyQ7vqmB5Zm8nF5Irm
+ueurvshKTbAum0WIKIcS7ArraOhe/uTshDgeYD0NCrJgOU5xt0VQo7eRpDeZ1Rp
iBVopS1puiIVkcqU/mS9OTQWludKAX+VZth6QcBl5ebU1INJRUN05XkfwjZdE2Y7
YdWMIcHbKYirsGfEk4DEZEF3lELcAybzPGsosMEH4bavJt4NQEINXQCOJFye9hBT
RY2Z14RVbko0Sr4y7qur4i7MH8a+iSja2hkgWYlg4Wky3r82KNv4eOrVQYYCCBBu
7P010prLIpO8EUB9Zho265G5ZV9ITnueR3fSMw+RZ0lQli/iXVYp0dclZHxbimjz
OyE4fMvPWd2OcOC22drWnYpxxONTItiZFEFwJSbdcOA07LIPch5PZtIfEizMN8iK
hBL1myxB0DVkrTRFRIH1X3JfIEFoHAEJgVS3dvtRTpaY7kngA4BPLkr++sPvIY6B
oq6Ik2RoTjtzZRtUerUMjGHYygwkdCjf5NODwO3SZYH1BDXg5MUOpzOvPE+Q/efi
xDksHjwhNwQSHLhKeXoexCPLSNS3ZW6yj7dZX/14nGIt3qExUiaSSFLpZva85XcS
dtPcNBav97y7en1JqZ3q/NxkOmT3qUwyTQTyq/oiLh6PJ3jMdkgpqDi98gPu5mrU
TUsoeNfFj/jS4sk6ACYpOLK9OzFeImkgys439zJnqUDnow8O6EkNYwOfqjitr2d0
UCj+lnX33aqTW8CHp+cr0bX4zK5BnwCZ1BQ7abjJWqRyhF/HigjTSakzblmMVLML
csZPpgfn6s2HbAg3K9w4Osq3AVm8CiCB98e6Sijm+/SJjvK6iWduvkNrkcObXwuT
3WWkkgoHPTGxT21OxzGlaB6BsxDduaUqrBn2DOGz4bpl6sNckwIqED6ig4OrvYFE
BoZKPLRNlQNZATZqoTTZuV6zdkIFfGmWLfLkspFASpci225oGc9v9ThusjHFZYEQ
lcXROEYnQTllzllJJVgh/CQAoDi2KVQS2OUS0sndBwPtwB6xpn6jLSof+QpF5/Gu
HbELzUlx3KxFmJTIZOt8KG649GQrdJYkmFN7SJsjEk1gh1+vc3xb2ppuBhpOYLWu
x8QuCkRfFVyImIFy0SydXkG4jCf76YbPqtCFyyqfbYWw99MJFEvDfWx8Hl212YDI
roys0rCeRCmKIgb7Ri/nlsLphn522mEgx77xsrY9LN2cSmS1mjZ4XhgzfJwFbBlJ
zDE5us4kLFioeCgPSx1qJ27kxxvTpGTGxOawLRC45bR/2hde8hWm9HKDsBwIDlX3
i8mXShKDFNw1jofzTDxsUbrmYpSsOtz4xkvmPKD/9qcbQR5Fy03hDT8KOiD4QQdm
KkAKrPOniTqeFYI1pMw2lFrhdfiFxh3YY/fRLI4K18g4uxd39NcWU37dhnAfco01
4ncK5+3KApec6a3Ae8No/H07R/6D/c30S29y5MD2c+aqdjDy1Vln7vLLIZVGRyCh
9TgC3aeawTxj6HnPKfkzmurSzDZF+rElN/Ry85W2xn4oCAeb79Vbns+DAvH4vhrZ
dm8e7ilMsMHstR/uGaqj/SloMLMwPkvpu3vGPO5k4sweCxfe6TM4r5YlKd4LSUGM
3Jk+dQVk5bbo/3bw3iKMiLW2aeFUO1Vha/KQbW9FeUL5jakGfZy+KFOe7MgD4B6S
gjnj+iM8BaH4BNM6/RaOWDM5Os1/+NdvhvScfacN37vfNi1a+q5f1grIVImjK129
ywEbFtSetoBOQ+I0z2irwCg6YJqPG8mriN/ABsB9FIFvddpM8FNByV7SQXbCowFA
W8huAVqd0D1A0sz9Gon6drK9YgEb4rAh8xab3KGNqr18uxlnEHGcNxGfL0HleSY2
6K6Gb5WPvrWAxiKdsgvjdo79nzf2MvL/E+o/m3PvhgT/hewArEV7CRxVSNecFUvv
VXasEkPq6Mls7NWTl8R059OS2O/6qPEgYBPlBxDAiD7b0t/AlW0Borc3Bftoe4gA
6yfk4MDwLF4iD3pOOX2G/nfXs7kdcdZJji1aVQ4NySKrbv2xURXlGC2zSUynbl/x
8+zakUYjae/S9z6cz/oT6Bx/ileSJKLU9NxT49/Wqgvj+HPuB+I838/4IwzMEDsD
SRVhLvq4OS2XWPE2XTlBLqDMzbhxBE6Vix7bLcW5fgEhfKcCSFYhioP5H5ZGhKCn
jO3aoRWRGAnz3n/5F58AmxIKDfzWav1v0LPunA+EGgleoRby5PQ7iTraF+RgRuTJ
7aGzK4+c/OIhII12QqzpAAjJdr2ws20BJwO2uk4o2azBnb5rv5jbVjOLetXHYqom
8Gh5npNzkumTu5MDQKlILGpJ/S2A+9XpioML1yOJygu9pyCTTTJPjm8s7QRZdxH2
/tTbJURhL0jUI2STci/99+OylC3zWz3j+4Qg+YRdr9FFT31keYKhwLjdKjCxKRVr
QPeINDle1vSrM+S6rtR24iaHjX6ZDQz419kEBaZ19JS16/NbeUjmne6QBfLIL4cc
8oktUj9NSIJ5N7mWmeUEl03ARK5nPkrEHBo9a326kFc9AkEcPze0cpYtAn+hrNaa
U3LZxPanJz9lnxQVOh9YKWQ2+vaWyxIfpveOwOBL6mk5BQMB475ExyvXZG61yS6W
PcBo2WTmo/pLELueaPCwx76daDw7wnf2ELc0OMgJOGrT5JIjGsn8Fc495byu3Nls
ENXhIGnyxAxmfvpLE7sxLfv0vUdHtxs17OS+Ys+3K8VFvR/p7yOXkqaNtPLLkbLU
D7jW7REZ79gqbD6R7WCZTbbPHZkauZeGNHwlBd8Uqofw0UkI3LPfoeJeVei87H4A
xA7axWCNOgLL2CVDunXGs3baplMQXrOdzmEtbj2Ps26nPjN7SbQsOgUsbf9P01Xb
QiyRQDvCtIhWvbxyJaVU7qPJN2LXwz3spISlNLYk9GjOyVb4srN1g9ZT4JWj3dx2
0B8YDjS+X8WuedShd37uTvb+vlTSbF5JfBmF3VUKVfvByUBCDxD0RC3td/+by4N2
zFfv8HPDErutYbJ8ik5SGVBBm6Ynmvg+dyO2VxjlV5oJ/gv+/NT4lopXhmoe6OoP
dtAD3wau0ltRi2liwT/2Q3yXZ4hwj56fPQjjNX2ah+/rajQmRtXdD2FGB0VS2zVB
gzi/RMk/pqVa+pIm4WpyOZRMqsVXPwT6ntu31BI1s+/pyczXYomJt3B4CzNRbKpM
ZzpWJM6m1KRVE4W8srCPSmOsNflmE+zDo5uCuuAlVovql56UDy8MYreKd603Bgjl
VkqtynC99MscF+ZvCApzjnV6GdkXp85WxY5OVhDlwYHjlJGiZAl/YdIAPHGo7sKg
Xbr/NUrJi6HcGIYk+X8YDFKg7wCGe2fxFx4KNQUhn04ru6R3ekG/3dzcLNjnfp/O
LPLCxOco44ZtfLGmhIhF4mYSX85wQUOPTaj8OhYE2BohNxEKWfCA87PI8UIjdU1t
kC7Z82nMEm809WpSMwoy9sKxGkQjGpeFtsWp++Y3c7h0JjIJBT73TGlPlACAQRF6
NTWFS4wQq3TAJAynka6wZHkjt5l7B6eDaezE7Xt3tG/xpwD8qC6yRGYeB9bsSGnB
Jtj+9z99j1WU4WZfjMugzTgIFcObg+hDWDixE3diKTCLTqiZPjjZMX2nQi8ueJ+e
2o81rFnXVBFteX4yrfz9IwVTDPtTe+h6K5RmtlsKSYyw4wsgSTi5Hlv8xucE4k/h
5zT/bb4yoD+4mHcb46nDFiBu6xZmPBev+xjAJogHpdc8/eqQHSIqOBRYhyigLJDD
Fqw/671e52m7+D5dkfHOBSWXk9wBVf3DjK91dAKZPwwfc2TA8h04z0YjfhM0b2RF
7KIA+nnpkhG3ICFDDx0SZDjJbr0P4JBwy0vafgGmj55kU/emOlG3VidofG87QyHq
7arbx5+liBoicqK+VgAggt6hKB4p40ZKmiMf+6kPwJo9tZVDF+yGr0NA7HdnoBN7
StdcjoeZNPNNWn+z7q/w6Ak1zUkGLvjhbpap1VphHljyZFQS0hukTMkhXNQDQavZ
zCt+IMG+4Lpc5uAq/HnQ+wYq/Cr/j44ksnz2alf1zRG7eBqrDGLOpBaBexds/a+t
vsrkVy/E/g7o05hf4Yxrq2dcxOaOF1ZUExCy71G8C6ikC1whKyeTObjGrycMuSqr
hjqCzRym/I8dzQzG2tTMtqMwyyGWT7dIBA1ghvaCbjFWGBjWRhwnifhW0fntF8Mm
ARUxzR6R0kMidCjCNujRaO6h42d1INItmP+SLz0NVSdh9VNCFYbiAYHb+ldf9JfB
/4kC7moYTKbiYGctn3YkpW7+chTGateBq8TGR5JMgJwmryFLITUPRGYF5oqY0cR7
sOSpbI7yyfPxxNNZBx4enrj/QGNezDFAxR19F2DTIcVJjNv6sfSvfFCc6myINgdU
zK8vwcbHSVXfWm5RYYBFEiG6B+nul3jQeMu7Xn/n1wdDN9m7rkofAD1DgWyXXOB4
IQxer12uKfUWzd8ltcmKh1UHCXFPJvKRiT8esAgRbgfzqj4LMLS98+U6mag/Sdn8
gS1c3epV6b0VxcC8wYhBtSL3q0oLowRIdwrGnmSU12e0vPOSBSJECm5n36SU9qR7
pFo9OnySCRfrOz0mSwc1ftXrink2UFRJn4pHm3BwZkbDCTld5yNN0jiQAaLHPqZ2
edB6D6rt2FSajxn4GjtwjZRcNVBxLYFHTgpYjlB3ZhYYTfiaygFyM2ot45miRDbC
qPzuuVAdWtSnW3DivG91M/NNYQ037wcj3TnVslfMmfxjkLQn8K/l58ZfKHX37qDm
TZey/TwJnykRDP0S01GdKnBfYNqLEmv4UXoWaWG3Ta6/6m5SyYoSGZL3MLwgjTec
y+Gi944D0XvOj/UvO+b+8rFpWhVQdIlRXJlMk++qPWX+ihxyXeg+Xq2v5sp154G5
S+gaK1XOV23VMeghwS3FDTU3phPMf/AdFLJjwhYB4YfjhczDjclWBGgAH6h6CEDg
FkXZtyDsxlZjwL8DimEDdLnzkoVo+YmJZpFo+MWtD1zWjt5yskpFQAQKcCiSyJi8
/N8czrLCiBn6q6AnuxkApytVBMahBFMFYP4VXo781M1Wag1v5Qg23Oe7c9NIo156
zZjA2/edfM9ggz4xO0lxDQQnXDmOJkTtkYLrE2MeVq6gHWRsvmYkmIwW6ocfSPvL
/phgrvqqmi4ylovCBxK9c6PilYN4bnMpvGInghPuQgO1P71Enq9z2dzl1fPaqbVq
zX5sh2hk90nncZi26TYBqK4r1OgCSxS7VhZOAeaqGJ9xrN2UNm1D+/ccBM8AKdiO
ntGPjdWanBv3vqCpwJt063h+ue0eaFMskPDIcfe7C+xQoxP6Fwan89erzRkHbTzd
n925p35rCmRjGX4k2bvnm89mSc6ErJ+vbjhUwfwQFpor8dv77zxjmMrAyUaX55Tw
TNEn5pGqr8w4xZnU6jvjwSxZseJyOO+jjJ95SA2jDyvtydi69kZAmb1Xh+jPocKH
Wp5YWSOQFsB2rKjCr7VbmnK53Z6989ezb4OxP+RoxRlG9Wx7+HrvP6Vmu54FTAvd
pepdRX7O4qEP9PNXeUqdKcsg5ovkpme8lbBMrGbcLrNEUDjkAVDPGcFbDC7mFXk/
WNnQ9cAdQx5FqJHJhFxNDhQLext7kAACeQh8qgbLEw9NnQJZvULpbi101WRx4bQp
AvQtEj8Uz/2/WUlMKUzdmsdnlmy4fLHzc9LE5lQoH/cFUqW9F9Hd0vlLlQB3zzTJ
cfc6woBhB2jPqgb7w9YkBRtojEAZ/0APqqeeiays5qNnQlqO+KLgkymJ7qfyR6JK
aKvVV0vi09Fm7FmwAVUc4AoFuWRmqVW25sLpW8j9190+pReHIWP1L+QAW5PCk1eZ
CtL3xGsNJkhgZXF495HDK7QP1eEQleZZySe0/rqeavo+7g0mnhzN1b8K+mc1ynsQ
PXSmb3k8BogwjuOM32Jrj06n8Bwp+yBZQRkDTBl5TRZ0VH6SLL26gxMRi5/v8cs+
oyhBo/F4h7YUHIf9CZ4PXP6qezJTHsSyWS4RULP6Ze/BkzMAWNpYHdJ2MHE/pfuc
med5FT2sfFeFLWbVkWPp5jTYc97E8zHdr3I92W24BXm3hKeAwm+SRbK90+pKIDb3
J82rLCpfHigcqAt0cIlKWQPpFZH19TrC+A53t8Y5G6ikejFnoVFCXsgfRUpdzCh6
u9rtbWy+OgA121/VD4cDz7xPdrrUpHsd+tvIaf7ZWasWkrmRV0C75WBEVmnA4crt
ChdJBms/NjSziuyCpTQQweUBR4gS+QCB9rqCrVYqHtcaSznoVLIiqGJerTqjlE42
AGQt2OrPsqeIQI4bDR7lshVAGsPvXGEo4kGvstl+8VXsgEQTMEHlKmaQl9LaSYs2
k+qD9dsTencXUjc4qiExXsCC2x0mwA+WtGV4vn+UzOrxlau3Jw4JZbyUSpyIMArA
fnhULAIgEmcXPXftg0ppyg4/yVDutmytE47USinmvAZX4MGgmlSbcDGTDDhX1VfM
5ZxP+34xUIgq2r7rte2tuvZVVADLRhZInYxM757pWXPn2Qo5XM/OeZF+BSXQE673
cth6f8TPvOM0TtcapKezqfHA/Bha4988vf7elk252vK29A9/P0GKNfgqnZaZC/bJ
aRkX8cotDqfa1LAok0ou77hJbLPMjEERPC5l56Pvqwrr0xvTIglJDM/CcmpASPOl
tJH6HK3gYND9EnGPn5flgZP+kRyWVaH3Tv38oPTz2hcOfWM6UGn5NeYeZlPUj54D
Ah2NQWf2f32cF8phUr9nmQue9d3ZOtKsRlpMhXwhZh1JUTw/IduxrAyMj2B64CzT
jdIiJowHUF2SS6NNKuDA1mYpmbbH+1wdpzSB+0OLae/NZvx3g2AEk2Ap1Liz491e
j5jmqJmlvlaymIE10E+kDDgOdW91RGMDADaouDyj5prcWRUiXZCzZkvFODs6fU8m
HAOgcVjaAfSHhQQkw5uy8x+VlhqdintRt8ewHKwVMHw4Pdi64hrbC+oMFMnNSNTE
3rEffmbzmFdqaMp4bPbfYzYEFiBrhaAs+HKMeg1APnhSh2uRh6BfGMNAkKfI1c54
wOBvC/II312PKDGl8+IeEyZvh+X6zwJduGOxTsId8wQeDpFjdOSHbO9LWPHphDM2
cZf9WQ18biZlrlOZalfktrcV8VfoWxnmtqqgQZbqiR4KNflVGEeT45mjff0CXhQ8
jc0Fy2SJyUfWMPlGBX1p4BMuvcSYW1XkqoNbRiA5r5c6L/eYsyisg2baHSiKLrRX
3xbFDMrTQSbhIM9ho90P3Ogh/nW2mvwohS2xJK1q5GR1+obbomz/+dq0myR8ivAk
VPxbE2L0bdQILPpWYPCkWYftjJILqqV8zOqUPfpEUlyasS103eRGSQL+V7BnDbdo
zxOA6Lzs/RbTA/952cUuV+c/7vpQplrKFFfgMJkqiVJehduSvh8QWNSSkdlLWPOV
zBOswVbCUo8U8vIpWyJpv+MKGk2DymRDVdATrSQxW7J98HzqolM6PUewy8NvuHZV
pcC1zZk0A3BPPQG492Zo0c2ubxPK8sCInILN+vIAaTX0xD//52kmlsnS/9ZLwent
HfdATYKyY7gEWUsSc0bTzeMexKO+8eOCFEfxkk1qj2+oOgkCdV22K1979v3YOAoL
gm81Jthy9vinhsgNKueCJU0EsLE+Y4H3rl/O7AerSRIVhxSuIjVUbpd7QY+Zuqef
G2OlnDCUOlMgHsIKyzuLc5gIPhZ4t7JjQefCVm0PDr/nB1WPwdn8x/XpiMB0Jaax
+2h9vAlI29PrKeLeBLLBsd5iXmINUM7POpQVNQxuKlRWVrn2O1GgHD+tgaifQVzz
RQ5dPhTqi/FihyMxt+6wN7CDC2xOj3RrIQjfMCfjzW3Ell3xPzKa6LG9ZEUUJ4+h
iIE26qtBd88iV1C6DNhKxOWF3TPe37OSBcf8YL2y0gmuJOby9rVbJ47fK76w1Tlj
fqcF2RYc4NWpw7skDmGtGRosFvYI8379Iqfz/uRuRsq7ge0uMYgG3LQ2vSbRQOzT
cg33hujN/pJGJzhqRnxl+zlMjCssSzEyCwIBTYGBzmVJWDNUKHlRsUTo45p8Njtd
KAHLnGllkgT+S5sR2opYatG0MdgMrikxlvo17PiPYuAqYc9TcxRc7Lf7KH+lDvBb
qsnPO5iimmYhYHh7uK3sspP86Shf66JsQizTXW6d2iH2dQgizo+Wl0f3eHiTM3ir
oAuYUW8XpUYXeAQfq8N14y1arUFszI0OAvLCAH926pLETL/EwXzeoXdW9XAbUvuC
aAF06XUuS6Elcip0/w2erMbsiDXL55ZoEBMvXNekkTER51LeRkpjp5eeYDcTTj8y
y3pwpFE7pWQwlNB/Evoz8WA5IPqxET4DyExGR46+9sRBkJWZhiOz+vBwAN1ehFJD
ciPkfH+ywHRloljxMgA8+ajxJFbl9HYOKr2o6IqMHXQIBDTK3Zxbmn6rG/Uj9b48
VOtgFxvXVA72ptMdz2cuG6fAd3nAfNbySpVBGMLm3zopfHnNjuKPKPvktKSSDjCJ
w4K0J7YuA3XfASPCOS9QmcsD36nGJz773hjeU0c8xg7c48hGyjjyPjnhezTNVWT4
9OCKcKGv67o4gDoxFFZBwq3jEJP8Yr5u7Ml5cuAIK1BL0m4YW5BolHXVhjRh1RDT
OKEGGwlMyS0aWO8nKzQHnzHUWeYhjv+LW7A+lw+gLV+hTkc3cMn7Em3fsN5tWRET
RsXoT0DBsulZqXDCC86MNZPCfMvobQqTHzN3z8LmhOEuLOGcv+QjGxsrH2IldIhr
UuIeqpC5169X6VfpiYa89JuCygjlZg4w/F8tVtolUw4w5zYOo8H5QyOmfl1RU8vZ
qHjlYz5g505DeFJZAnCi9Lmnpu6gtxj5AMyQ0btm5evjmmkL992h5Th1JxGmIaW2
S1B1sFnR+pWRrEZ/y9B1MHhuK/iSfryJTgljXUVPcKZ1yJIzHPVMYl38mBzAa25H
dA9ZwXVPAxs2utb1g5QGbpLd02JBFw1ACz0XxeqcCKmTOvljYtGxhTcR4ZtxbY9m
hZlqlGUb0ksE2Vfxb8DftyiedZieWTBp6ATThxDQTnArcMoz/kVSTNmp/S81wRdj
Hjg2xROIs4AJIi5+ZItMy5N000PI4NVHewH75LI/uKBLW3j2Dnf3BjAdpP9n0a07
0qqIaYFnsRY4CZLDwzNlMo5KBJi4gRQLtHdDNGnahFVrc+/9bovHDDqUpb6RfmBN
8SuaerbH9ZGDRzxzX8vHegr/EBlOqkgLUiZJkOetgx5SXh27osWAkDTUGsY1gFdc
xewtgKd3A11XRcoNQR4GdkzmM57nAtPqHTc1xiVXsOebyG82h9/DNGGe8g3t7Eha
tltjfHShakQpkoBAo7sIc1ZBEDLbDpGhmcv8tUO0O1+GqwBAiPINGlcBVrWfairI
QFGOQyFMIztYk5YtBqZ86Rt+pS2pq8GwBfMtuGBsznUY2z0K8VZWRfaWk5NWIbnn
N8vgSm+KjDJf5c3WOFNGjcuMJ7wcGN+T6YYCeJZCs0JykNw3IvkFD5Ue/ZceAnUt
XAe+OTYWofP3Mn0IW5vq8WM1JfBdMmjyDTEaNj+O+6Ob1hZROHtN63dtKa2i9KkM
TkS5lL8iiwjUkXsF6UudwxSHe7hxlxWHsu3VSz4kGy57VM/UvSZ+O8Z6c7syue8/
IJtQg1jiqWKYy4FBclhNEVBFDb6IaOWt3Ae0yYTgy5WWy/qq2UQbmstywcMI7cKm
J3miHL7JkKKfkrY1deDvrM/NLyW/V7w9/LBVZH+lUzHZfR2wuWCuSopNl+h2oexr
oLkaBVVhGckhCrYsOMRzMfuLi1QP3Kx852noYmhkgr2ZGvJCSwRKqBTkIdlf4Ajh
bqdtx0PIxVyyHdPK52toEdUx5AjfYe0TIfF3QZseS1gaAwRCn/60ubYBtzMhF6oQ
NBw+dk8a6GBx8sxNWMcul263GP3/ORcZBMQrQKggHvD6xMCNsOVE8jT7ai628N/l
NNrFyAL6Ao1FtX/WBMcihOS34HrA/0OHuPNC3MjbkSefUJuUwE9xamEPVOqiWvKv
TpouCHmUrFzm0JNcRMZa2+6x6wgr+F9Y0fkcvojpoH0L6Pz+HcT1v3vYXeqn2Lay
CL0szgI9kJUh7jn37IP4pdtolavVlYhN+Kd7Z3zvWXKUn2fzcuMPsrKtRPOs6/db
nHdiSHWvooIbRlmigRxjGtDtAX/lnkmFbDMUpZp2VZ1UnLdCsuaIB7uABcrZdszq
GmY69LKrddYpIO8B+fCGoujhZBNlUNdP6gqemCAzZ2rrA4V1wsz5kwr00fU4SneO
/EcXAgRT/gDfrCN8emE9dPGPSawHQNRZaFd6iuVZ8XcqU9bXPue4kixJS/bLl6zM
VH0Fs5IHvrqysWuovgzrATS2Bmz+MxFGw3f2eMEY8UC45bIc3Xp0E+UK9Fv56iJi
4Hy1u8DXhIh+4GqO4JiTqeX55CmzwwamwFSp8YVthVqwpg1Zc3C8lSbsBNTd/gKc
eAH84Yqhs4+ftAaW3b76d/ZDcAEQ4FUlStrXxC5q+X1Uxn87/ZDQ3kkKiRx8m1mi
dG8LjhQS9aSzdSpKCd78qKDGezPco2odWTg4dJFRuyQ+SKSvgglmjZckGoRJF2yg
95aJOB1uDES5fqhnCROxRUx/bUrRXYncDahN8VuQQkU4CT3zx293RTgJiuPGMd6B
oVrNPTh+GMS95b1hw2lUAxgCZdIaLoLC6fko/DmmIePDqH4LJne2QO494fllMjE1
lwSemxDpxrcn0PSrbxd8zJEfdD+xyjN9e31jPW9HSuVIw8VqTKt5S03QTgLeV3Zi
h5mjpweMYpUOWWvRs0ZWkjuEC7DO+7o4uTvRK9mjficLXeoA+GI6ZyIYFitgHoqZ
JKFVfb7yILT4eHybhaZIeJbt28S7X9a20ramX0le9VqSSozFUFoGRYusdbnfsze+
bGFzp5GxHVfxpIwmLRNTcWVDg9GOd+2tEcyJxoQ50I6zDWCSy8fILl8vHKZaqoqD
yjprx+kkuH2vJ9zCVSeuRK1Pq5KgdjAtBf7Z/LjwEfUEcNrLG6hqusb63X/HxNys
5OYpN7qfcFnL8ZMB50E4ZFGGRh5QNbQ6xuAxT2mne/NVXs8/LiV2rYmGCUrm6l7w
m49o5VEIMSNCOa8To1/DeKgn3j0s41FFaMivSxOiEEKriMlEtibBVlHZdG3eOrhb
efQSL6+c2VmFX0hR9djUH2APWhRRJgnkUTzxg+JNyKU17c7xKqtq8wQlFX7vIyF/
lIfU5E5ok5H4VM+f0hngAdoy6t91zlegapd7NTH+9w8OYFUk8BudphRE4KieC+O0
p1bQpDj3hi1xJJwQFbjkj4fNs2RiKFmUvvc+xS1Msr7vsRjqwV4e22EhEKxIokZ0
Vnb5EDp3AXUDV3/N+esmy1X0s7VmAE1k6ZPKqL+HIFXBQUdu/mcffKxCQ+77VS5j
UDyC4gqASOz2NRjwrbDLOUvBIagQXOHQAPbThWxExl7yli6g1u4bDQPAlpXScdnU
qiGigkcIy9jAiy84VfLNhBubNEJpPXZIf3UxzoAP7sZ+ojr3Q+XPkiOIsUp/nk0O
X8gzioJPslXrHHwtO+vNYEk6r8QFH6Mf1XYUS2P+SW9R8NRgY3wEbIzgXO+WuB92
EpuGE4eqVg6xsZUyZNSHyyY6KYqlsg0+9TIM7zwdyabZJq9pOslFumbgGRBz1Srz
gF84VvJhrjSPKnrwDOEwZzy70lAXZxbvgUHIuJK0rIObDhy1Ba+IrM/Wv/cs/0R2
LB6lQ4cLHF/XXDYTJcWOoeVu1XV1NcY9aiYpu+14x/iCklVdc/RzipY5sTprVFLR
h1ta3O0gJQZchLUZtrQDtxs0SukQ9dPh5ygCxZwDInuI6czOJLxWqyVsJCL6Ln1R
pdH/k/S9lQpOO2D7daz/JF3SvirqIl8/dx8+DDaVT8/yd30YKlyMde435bxXBghU
QxHVoeb5Lm3v99q1Of7y9u9Q2jGT1OKD0XNr4Dj7EPvfRS72FWTziHxC8q7a0K4A
KQCfOlDF0ih15psEP2QGjT6ZpuJcgT7b/w8+78Q5306Je2HLvCEzMqaP395FWUAq
lWP0oJ6ROu7KaOU47G1pFTuQCQ4V2q6CtYHbaqp/YOvKNXNJeA0xfEwSqS5N6LdA
W1+vN1VoWP/jAYWPg+gLv+OmY2Rdz53+YYGqUuNqm9VWutPEWUqpiq+if8UZ5eoX
YGPCWcw76a0VwWrwcWb7QNfY6L3EwuXKgz9zk7Lz7RyiH+jya/t1xFjYbiKRVYLo
6B0iIs6DighrV0sesd1X70U33jIFXMF8U6KiD2QTE4s5nQhmTrfwpHx2TgfdnhFi
e28gK9F/NJio/8fAplhXvOMBYlyhOPUgsIzo3IEQOgPNZxTgz4g5v2InHOM+kFYN
t/fXcZQ1pvsai6hdEdjD9/shPu5ch+8RPJXv8GR53e8IWLW8XZeN1VYdQFsW1T7a
+1ASboRbhyglPHSFn8cOdWXhjxhMCQetZZcsjIZjgzEzOf5zqge02QDzH4OA0+OZ
U8wxFYPUNaZce9QqTMRSBw+rS3J7LauHhvTz3t72ateekAh3dCJTEDDJB+CM7mUu
GpzIPMXaCVrGnnfJe5/qUtgs+G6SK6PKCWUknIBpPBTPlbCSB2XZ5HtLlqhyDGpi
hm5J1cIowYu6N8eSXu0cYdX2OqluwMkXpoHdjRvJmFOddsJWCPwd0Sw+NgR7f5gS
k/Tuich1SOQc9Z2L1ZMGnSGfukatw10UuNOFlpe1Bcurq4yq6cTxwV1Hxo5hwm98
Me2Ltf7Bc6GoZ429xuHKKq8WW0V6vFKM8BlChDh+MUxrFXxaesvTONV79Xb9/vYp
uHHaAFxEuFN+chDB0jWdYjDcIWogIGMm3wzGG6U1VfywW7fsH09eOwurIVSD+GRo
EfYVfQ0NqeBPuFXSi6D0YGA700D4+1VHcxMvXzJpgpzOTaAoBq+z5t6TlKzRCSrX
7JYzhRE9sYoUsvcJyGcupMl99JfKb4rg5CmT+xa1SS+Prm//Vs2P42lKKyL+S8RN
ny/HNeBtb59TFxvVZvWpu3r+99zYefDCJcHOwFMBnxFus+hD+tkD3cpuYNq70fZv
NRbyd7YtylKV05HFaiKCDf9n25730G5e3vxFSHX0vnvOVNhYefpaACI5n5jjtW60
uLieabT6QPunCBtnZRmNrw8pOj+ci/db308G9iM4XOCTQSmoJR5yFX7UjLjM1lT3
f4r7p0o+gZOK/Di3Rk+0z1svRZsSxRI4AQNk/+Khq4RkS4TyDKX5bRPWLr1Q4wm/
mOLeWv/U+OcpGb0S9JAbeiZ0pR8a1iRAP/vxWINwvxwwuPtYj0256Y2gN/mtdVVc
vewi2sNZ+earkkxyr5NPt16FXWdNFWs9NjHhKIM8DC35/xPYch+GZ8LIK/QgFL/N
Wx/I1vhAP8ELbHyMrIi8ZXFSJ3b8/fYOwB7EsJ5OjBg/5lk1+6/Y6HfRD+GRhfKS
Uh3d5+9rW/D+tWvYC+p7tY/VSL6EMUdqsHjFzQ4oOk3nqVbmgSLYgYKeZ1is54LB
sdEzISqWILbNb25460GIPVRMEWaHwmMFFCycCJ7xf8QF/qltwHT2+HpQ7Fy08Euo
KSqS5voLW67AORwTuA3BVI5fw9FaN10v2Ep2ODo5soqgTTdylEwZJ1hi8aGCnXgZ
3PAKgoHJziPrCs16x/gDEumOy3SrNNVUu5Z/6Kp9Qi6Gz9yvWnVWAUWAIRMgf4AP
G45VPf4MbIAdogwD8+5rnLs1XaRQnBASXiQMfkJa6fIUmS0+2DDra5EhMUANM7kv
EqLee2SMIlyCfbuAmizbHlMp9qTBo1CSkmJ1gehPvtY6J5+FSDQ++8Y5G/dj2SZv
VRT03O5Y2R9OwzLvT8OyM2PPGhxqfqebwNex/HOoFgFP/qdw4F89/G9SN7FRBheV
vVDWfF+hZvi7rFxERQ9qe8rZ5o6gyHoBeMyL/Y4/u5kNLCnbVU8buX3hM8Fr+Euf
Lysk1l7tYnUBGyUqfLNAh07Tx1K8H7zrKpj2IfbsTDR1wJq6ExIVtffBV/NrDEfN
e420HIlEJtdnUlbrhcSqRBAhWH9/8fyXX6SsyD+3CAV6Vgc26jcY5q5oZvXIesTO
Z7KD2Dg9IbBb4n0EfHZDNe7TNgFhqNXYvqq5222wjYCrDgMf9pG0YwULDYU4Qod0
2JDJXyYNi58+10zzLLAE0FTmEO19q7tmGw0EJjRmL4cM5nQioD3ZA8RXuj1W0aAG
XnycpZPtc/3QabUl70we55xxCBef8rsivsdw5orY8x6YNPWFmQfW+i+UFqKewoLB
fIsnWy1rjnvi7X8JQwi8tfOxXPu2pqw7ROZrmPnJ9pEcMPpOpoefdu7E5oBZyjQ0
jl2NPwdvysPOHaAN8ZtCpEzevnTv3wV0JETah1sJlDy476c0aUuAvXxNCgpJa3+h
Gb1xHZeoCVGDl0pDvfdRp5M+zcjdN5q8ACQcG9aAbjgu6J9VLqhcIE4cdYYxcuck
3vX2q2I0uu8+/2sAB8qSlmxZur5yhxAGhzNVFfOUu4/UTuFWMglyoM4K0ayN/VuS
87buUxfBknXCtltE2flMNjs1yaus67+CUfdgboOUfr3DoV0pU/ZPjPWP4wUzHzNq
9ns5wC5Z4dFleHCsyE/vIYvJ6NWY4PNR+diDKp53dcMblYCkU0zchuxqzF7Z1ZCz
TF0eQT6zWcO9WB2Wn5jetLoMvJPMcoysXNGUIaxn4QIHg3MJYC6T5Z4pyxf3Jn27
sq2Eb5j0AF8m9Rx2esAO75/Lp13ybBd1ffjaVJmnJ/gTp0iIg2iQ+tsErU3BuCZO
erU52jKEcPxr1Ha7UdQxwZLla1rSnGqpkZWdaScM6yjjDlvc98XTdU07xazDf2CC
L1+6MkSBFm5djb111egjWydYjDlk0chFll6MqtfPkzEMzgMCYrXehWyXrHv97XGG
Md2aVtAEuv8Ug9QNDOf4tfZPqdYZTaxk9o239HN8g5cRtn642zfHmW3qEjgvzIrF
QHGRmo5wK7/LwfZHa2kDQQn9pN3lPW5r+kXcctOMT+VoTwwKld0NA46fx+j+Gu6T
mrFGTctRBrg6GbXH96aM9iCQz9kqtBAbuKbkR6fmxMigAvaPnx0TWEP9kl23mY1O
G/VVd/Yoq6mY7+/kS8gYjPHnYPZQmC8UxkOPAvRUGTQzokRVrMdFHYYUozjmqye1
ur3DQls1UpTm32qsAqkVa1lUmgppYobGUohJlnCNdYGBgFo1mUO1Op1aZIESz1II
9qgPZ9H6Fv4bexgzabRUzKG3M1Epa9QDZsv+vflJ34wI8T6AcvCCItILG8LigvaL
x3xBfnxxVW7CLAg7elxWN5Dbbhpz3YlTFme53hzUsVF0QY5ItLEIb74M+DBdp7/c
AIp4h4i+id+Ou2V6Gb0vo1oks+r+68B7rQhPCjc0oyIV+ozw+chE1kKzkUIaFla3
CYvls4/Yv2gK8jR3cF53S9CiUn9KB7C68cMinqjAIoVwHh0cf5EY7hLS6DiY3off
WdYmjg4G8A8kbr+CsDSDoIx61FtgjPEgRVHqM0Yfkn0D2h772olE29pfgVSvTDSR
oJavCEUfa8638X6/u43/y7D7JZPKGl+Xff2Q1eW/3pN1EusE5Nkan9XQ3OUuXLqr
Zrdm2/cpxBgtR7cr6HtDATq2zjkm8VfMxr0/QARRXqdDd1Jk6K29ugj+e+11Ez55
bw6Ham/8bN2PDnWYZCREL1NOKuY/vuQqlqu63thK41rSCNdfmlO69I+KUm64Pe7D
HssVLpiqQnaPriOC+L2fSlCrOBt4IGntL4V/o+WLChPT8wreCVTq2gXmJoBu3k+D
4J4+0EhM18FezbzSu9M1qu2sVqkMe8AFBQFe3i0NA23+fs7i1M54lhy2JlfKoWJ8
nHEr8baPN4XnNveVpb69j7hj6edVXRDzXGGpIhmRTYccQHfU9yY330wQRCu8IneK
AE5l4ZPGjWJyScYqibTrhsU8rRlnc8FX+TYrHheE0qlv/iRxq4bdZgzyp9l55lct
+NN3paVHygLQSssM407HsPBmVb+vpLYbXIAhPMp+q14WgchiqOFdv+dlbE1SK27N
4yPJXhq6gnDKs2l+E+qe/hDENZRaMieDaZRSKy5XQ+2P8gSxRaBkAh04r7LbrcR1
qOTinfbB8/uMLI+9x+McJfwY6QAty9AIvjjNNKpvSP46yabPNl9boA1SLrU7PiXB
rBETHjAWkis4+fldKaj5InX5ruB60nRBpQ5cgVOkPqx+Z0eyVz5e2BUKyMflc2vx
bXIfxaMeqS+aMTLsZLM+WCC8J31/K9cHYHvo63dSj4GOdKpvWfqolW/xpPKQ7vbW
pUVnAucPcFO8k2YtYbFw2GzBdcqdMbhJzMrfHNkUigD8h61N3YNnAxyC1NSYEo3f
xB+5TIq/sJ+o3jFjpf/P2cDk4WCYpJgO3TiYfE0PMn1+ohkUcfK6k9YyiNhxWkRu
jUef2Y4P62+N1v+TqVF5preyjh4VMsQ7RnxVzHC5ML9FiqLq0vQj6yr38AyIGuAU
nwQmSgkdSyBYfJhrYKhUE9Lqi8uQt+rYDkCyKuGhtHcx1mxU9gwZCy/amdQlhSKX
0qWdkac2HaB8MWy1KfUXryGAHZTp5C1RAAHoxnevO/TnKc1PcsLPkKqMZPzeNaHn
L3AjFRM42U8B86uMaiHSfm/ck2hmaPMkWTR1vF/Swk5uaNrDnL6Hg070lLWazzR7
JQaEZ9TddMpBF1Y9TdEMJ3up9PruPEDjoSEm3NrwG8Nvstvkpsm7cabGlBezwq2c
XXAKTfLoojXiNjLcVdnveq2LZnA6f1IdoS0o6BrXOwS5DLqnZVYw9kYiUGQjkOzo
W1dMuaD5eBDPaP9v/jOq+MAlGuX/DmZxvYF0aHUFZrMBx94GfGp9aJsNyz+FVWR+
HZ1r4LRxj+xkaqObqFKtvkVj+qi/6m1toPweZptGYMBpRo7jnYN82opBKuT71rMH
M8FwSy1uszevvXmN16iZCRfcIPmy4TBGEJNA1RHkjRrTRyXJdFmxJz9k9acJuj2T
QNn0MB6KqfePgqCkQg1LgpMb8Rz0BO21MhJTziuaVjtZV+EEAqOMB5sR2G7qMgkD
HIdu7QK2fwRxS+yKBeLKOMbRvGllcas75m9NDMI91/LcHnQd1bVfWq9U7/6aj4kI
E6NatgrmFqAQLK/2fJhTObH0wqjHr9yI7Y+WJqDg4HqVaeOfYLL7ialLilDH64to
cNK4IRYK12ekTQWXN2ipdFvN5GF9FchABYr3kJpKMZXlof4Eo1dKWsg8YJhOjlNj
6BAn4bqVGcMec8+gPp/9hFhNRd/ZwX8iR7hjgZcQ3V5FtBhqAMOucOZLZ+JATwuM
744cx9CGW6TsaDjeb/56Kj0JZoRt3ZfQQLUmvR50DF5hkkzukaLOzIKxzsoK3QM4
f4GE7EmdTl36jAYsw6IlJb0xYwFY2r3p2wrzKHhbJ9P93QHZuUyRTpUaCKssjEQV
HERfgijnuI+ge4lB+2Ph2AP06o1qbi4Cl/DMyQMQHpAu9JCnDWUlyf8foJiAjo5F
/97a9sZ4lMmMjnSa5NbncD1vZo9XZWZMie0+vgir91ULXGf81Ud/B6acJ32xIfYj
jZg4i/00cnDyDrtuwwucumrmXo8RYLt6GelLzlkoIxQf8C7qtarNcqvIIaW8f3MS
PtUZUnG0omR4nl3+SM6PtpSpr2UF1H+r8VyweoTCKd67A/cEXXCuy405Cmog6vpz
bK3P2yaNCc7AN4zgLyDEFEatohFpraQ2RsG0G1+i2rbZPPcNeJuZsXEx9iwz7vnq
Mrrf1yfkK9rlHlK1XJNjL2KpJoH2UOg436J2IsZ0bIPnwFUzVGW3LH6xuJsEWLj1
0GC1WNNAsck0lQUdmNQQLy4qTF7w2VH7OCvkXmA+7f8BHIcC/UEXIzD84Q1HsFX/
nBdqlHRkIG5UrBZvUP8NV321tlvCb70le0DL+PmIrJFXDctzAI4764EH0Z53bmrx
qJusPUaI5J5clbA6GrE+dC9T9VmyMlK0/wPz/8q4nTCMEmFUA5PsjbDDodFyeiE7
f2W8yqxJYuHR1O2Sw2vMHM8sgiNjLHAF3fK/+B+MGDdnItlwRSYwPGqGNWOMwfnR
HGW+79pf33yt1nLrsKmY3aHZLEtNO4oI6Vvpy0eBxa0QKnEsInf29uOdl4q7H9Jz
VvrAMaDO7Ob6mTVq8Q727V7isOrECU5azF8t0IYkrReYMc2TiK8W+giVBY0Fyrb3
8MV1m94Ykfnwc4wE/hX1BccsWrzQiNpj8PsVir75k3IwaUL/pETKKQLMG6EpFvKg
SA5Ro0ZqAdbfTPvpQep9/+LVwvvztTy51QGWjvkLE1j9bq4bbnVHKubMx5LrLwU1
KhA1ChQNomDOMYxG/okaTrGgItMQGYNbRPTqEX7qRwdoP2ADA4we7uhLMbOEUSoT
h3cDPca2CqoTvq9UQbsaFJE6wmUAjBtWO4OwJ7LyQqZAXM2ai++paZiskD2IlpkU
pZ+qObAVG8gn3TfScR0Xeq9eC0XfHnZ1bbEA5E7+L8FkzNG/Iu/FuorihbU5HEYp
8mhmWNHgtJ+lJqlqGmdQABzE8lOk+fWLLNQqo/Y3vVNafCbJwn/liEgXYzqQHpAA
n639575pp1DT+nBr4Xrxnfyg5fIh0mKYxRBiHCXy+wpYVG9mrIPq7IqQSXpy7P+0
3OPVu7+K6wQXjqJUgV5ez/rWxHk/Q4XAFSLJwB9sSv7mukpBcZpxRbc5GHqNvrBW
RxspLtral1PYyZ9sLXZNJZN4sqXNj0qk+0+yOfvGidREYv6SnPNmW8areMZ+/mJf
Ru1i+lUcPit8bHt20yvspJC1AD41258UdMMuYOQLfFQN31gv9r+nq4tRyui6Il/c
1KsfX8cmHvq0DFN1XwjdDH3fqJ337/dsy1QPwDVcbVVripPaE1FbXGnTxhX805qs
G+EmnnH+mwxKBxDUQsDtutqqI52RDxJtT6QWQbWLXvnxwf5uGFIWsfyAWUH+i4E3
0fi1I6FxY0elDvtVG5vFdJDkSdPQSypPYOI1civgmrPLYzGr8k0iyd7qKhBqVL9B
p3wyOpWsNcTBAHTZWBREjLluRzZHs7YW5HW7M9h1fJZARQz36ta/if27X5XEu1df
m5ub6c2WRXveDp0n7/PSUglIvkPvkH4/ZX2Sc1dITuZPqx5yNf1dNEeyUkwjkzzu
SarMaFNyZ6+bz29ShRHXGs2BNAKfGsX0EqMf+dR9e/ci3BqObDTkNcd0NMF0XhQ2
hg5TQGEKd8pU1c5hiZIN3mhp1QHpCQFQdnyBbPUyQfy8oVLOktB8lJhCXWzF/w/D
gLE4oCocu/Jb7QISSzaNTQjgvp5tbaejBZdgsgRVD4ImNBGUDSz6LMAXrWv/UZRP
Z1PmDidgZ8IQf4QsibZp4cIXBCa+Hf+Syz1Pfjl8jC2q11pAjYpdzIm6F0MY7uEl
OyqhnDkHxGwlHmdsxc3NC3EsFljUS/KPiEQfGjbqjt3bVnnOGhK/9KONVa0952BO
0Q/Cdt8HQlUo580LkWYNZYuDU9YMmrw3mzQeMuI1w1W8iA8pG7C7d8jrFhW6f/60
V3MsXWerF7P8VeaHcCsfMeTFynP4iyWDiEEsvXItLpz7mioPGO8pEFlwsW93oVq/
rDgaNeIPHwSpWjDCk3pp3yPC3HatPFfC/K2k7nrNjPwY84IQTerCHBxYl0OPh85b
urShND8dsISCTtaXoE4Xi/E/h38WBhnkYVyW+evuhL0zvhw2niZIlJ5ucNLX3CNX
qpiP3fljfst46u0nZseieO5CD78TdzxRz6jjNuBSIhtykynIWlRu98VmEeCpL8Ri
YPVTXgO2uIUEZSDMmY+tT/yXgyYcZcjm7vnrB3F2WDid9VDsV7ygakt/8wMxpvBd
qpfR8ow4LqBboYWJ5cSMcZYyY2B7avSflR4xjTuMswQl3n8nPrh57LjLdfJixlvx
u/Ut01asY5STR2o1G0VSsFChSvtCriFNIbPvWQDHgWEyINF8Jt/LkJah2m2MTBvB
c+5NFs3RjfPS96kwiKla+5VoBoVIAdCO1Oh5HINsaL7NkUy8SEPE1TnvTOCtzd/i
JStX16aK+kbVUIX6DCEntvPiqZ3Ebb76tjz7eb9uowwQhCjCWXHCYWWN0u+ms9M6
3VUJ1hNVkOEXNX5E56cI8pqkNZGDN0tH9agM15qopR53QEALZpumNJUn/72a1eSX
m/g6UU4thg6pEKP+/ZX8MDmKKKlzTYfqVbnvgvqabODpN8gl1MVO/ZjYPg46+wba
K2aGwO469fS90WGw4wfUXAE0kyuKxslPAbYanSRlMzTjrk3t1QnUv/eIBvpTn6YQ
VyTCUNQ7lZ4l3ELb/Xq0opWVO1XnENdiVGbpUeKvuUvy+0eTQxnLPOZoS1p+baSN
5WXpmiESk2ue0A7emVFyfPAoJBVR/GcTzxJBDFd/DlxzXUJm+RX/wxFgEcrN8OIr
OKj+0pP1mcOtzEezkiU3mLZJW1EFpjVkvRjc34/nN5AGMbuUFF+0cb80dD0sDPN4
adVHnS8tGDFlvpb95DrMQiTsasw83L9UqwseJgHFCtjSon/jZYGmtIY3TdekYXK1
vkml63G1G8pGk4PnzGQUmh55KkoS6H00ukz6v5s6NEVvizlsZFtmMk4thYd0l0xs
qh8tySiqpsVLtSbfvSlRo2Jz6L4EJC0aWUNGNgey8nJGZEkJ71GdTw62qCNIzSWg
lTwKO0KO+2qFgCXpbtVr+g4cqC+rvvU1aZFnM7FY9LRboohxFsxRMm53mhCL/Vk0
r+6o3pCCLPUah2BrJTDfgTNZOP/xlaimrZRvbhqulQx7jRtGJyN36UKSnd1hu6hp
eVwO38jz59toMFbJANhBKwKRj5ijlSCAqYl8ffdV4m7N/bwhNCf7wLI/VfD/CgYx
x0wv72Oc4JhBrjJObTjl1nYpD8BOpq3EYMeQSXH12/Mrz7KWg2WSDhrt3OZtYCS9
L8YgjR8neleCewcj3Qm9jRI6xGo65prUcbkSddbUxPWJQSDgu49ej1KJ9lI0SmN/
PDc01FfXNtrJG4TP94nwbLhUfdtcXyT5zL1AxbRZWfdBRv/AJ4dBihELDQQH0tqB
o8+KuHUofhhD+MaDLV5b2RXlBizLJU9gqh01X/iuSrChEpreF8915+7xfen/jPUP
Xl/vwgeoU2NdTuA4dxL1tn1fNNyVbQaMR6inQVXrEwUIJlxfBwuIepx5m5thNSZt
R7jS3tcgtcYuuzu9jwsOZde+BMutKN7G7d7qY6bFu6uAjgleJiZjZW7ud7lNpvtA
UGxjGMYC2PdQTbQi4OJm4zQ0nIPjK0ZN3mn2I1EWFpQwjOiT86MqENpjgjm9rvij
TE86spSxknu6thBOAFXzGF9Pl97uDjUuh7YmMA2i5KMSwBMnRM48U/j20ubVofqf
U7/lAIbfDpo5u0komn4GHyQk51mkISXRQC8Gfik8yNgy1etX2+Qc3tLZp39ORKvj
a0+wsF0aAlvh0uboFPlqprAAjw7dDwbA9GCo1RujjV41/h1XFoO4POM42cFjzZJa
AVJczxIV4PltOUH+H2nn/QhKqsjY2yXYWccxH2waRv1wNW7w6SuJiJJIuhBUnzH8
jjlpNsvbgznDxWJCD5YPr8jnguM79QwrzjGrBNiGuUWyzd61MAu7KNPM003AjfOx
tnLJSLVSNGfVsNg5f5WiBmOltFBT7XZ2kVmsIuS/Nh6ByhaHJR3to68V7spaspu7
9cFIaJhBcduhdi2h4oeq+KibpYujmErqpS75tqObg2cQ51W+L6pQL4Fyy0J9CxDG
xu3KZt1P+RQYEG9Bju5g1EueHPuTSMTGRdmd0lxtrNdk+cIHA+2ROXqwq/Ub1p20
lvAUiSfiCx6+O+5xBLcXGAzts9hpuGkwO0SSfhdnrL0hAvdLFL8Q2wdwiMJ4lxWC
ASxXoF+KRqoA9ScXvQaa3FJxB0leT4RB3D34t1goXTGCoFRNfAzGUrLnrRT/JxC8
fsMLshOpV3PN1ZEfWpfqSrAgAS44AkQy4x+74wu0sGLwg3mBVNiCe32MGXBR+zJn
CrPw5I2x7GBNBkKWBHx7xgBWc5MiHmkavAQjKrKLWeLvVoBZ3kjLQ1sj+eDmWmbD
mghMR57VkgBUmmINgu9WtVTnDiSdcl3o6NpXwyZjVKFXmn7zhV3Tz0GkNtnMu/5z
Rx3ojeXWoKxrTgkXMUI10CMqOsS8SKNO3H+e/0IPdmHlK9Q0ArtkIvS8zxoJxKTm
6QgxLq5UF6U+6sZ4g5hAO27ibiHlD565vucxOX12jJ7DK6pa15jfh2xxpATqnEh2
iBYyf9m4M3BlLuzb3XaRfJ8AICsK+ZXuFxvgsSTNxSnF+oXBHtd46vu0O/ytOSaf
kPTpXfwG0glZIUyzylHLtEIQd/oLo7uGNee5AuKRSWqQt1GlBmrS0hwzPtnhuyQi
1trZmxHZG/Z/XhvjPbFJMdtzCGgJZsT69sKqnRf9SuTQwwhXgNt5ah5/11ezpqan
WhN3drQfDDmmd57QYo3XP2t7mKpcD5ArPRJ1ggMrwMaoOpdUDEgMsdq6kBtKecHi
4hkZ5HR6WXrw5DE9d2LAyYm6iprIdDYItplpzJ9cPVs5oxOZU56vF/pl78fKcAv2
GTXUqhnrX2OMyZb4c8dBEcHChwfLGnpTCfYE1tuwB9/Npvpl3z82POZwDsHIRjv7
zx3D8dw1Gp4GULR1ZYLibikT0/RYoV8Vkl/mmEFZkDfjtEiNGXygryvmKVA+b9EP
2wI569/fDbH78gGc7zOBcsMdBLHdVaGGLHrv1LWtQkGnFjrPVXLm6h8vMvLKpFKV
OP2MfBFpWCZh4oKunW7uzCc5WCglbZL01bvvDwVLn83dfaVoy2UZkMH37Ds3LoZG
iTZpzFHQUAM80g3+FiHojMIjbN+AjmCo5510Myf/eNaA6DsQcOhX6fizEN6kKNkT
+TcuDG6eYhk2cdgVDL9H7OA6vXaVceiXS8cJQSTxGP59dakaFE7GZmtWzQrWWY/+
2rlL7wKouLQeUtq4cSp0l3owZZOhbj5Xkv+scS9jSAUeFwED+9GPvIE8KFSKT13+
NjPu5DwIwPZg041yAmX7sZwfG9EQc37gOfVcLmfUZ7VxG5oQM2xLV37vRmKOlUN6
5fqdCk1KVxl9Ri857yCuiQN78afkXlx3ZjK6iiiYpRgZqhD4WVtpf2cn3eGnwL/F
dduX+IHme9uSQN3p1leg0z3aoR3VHvG1+kNLYQNmKMlRUTZv6K5Fjnoqt7AaxzUD
UmhY9guVSoBhFnu/xXQr8bZq2W7rheVLgG1iVzSONmymJfX8nZ3hB6qQRCN7r2BK
C/IRAO4S3Kiahjq42zK4Y0G8/Pno0n2rg05aD9WDEtytEqJiMoZrZ5mCwpA82k3t
j8lRakTx85YnKzUvI0mnu2KSGWE+6z0cDoRsKRWalp8sY+kDFBdyo7CF4vzIlSua
VThT5p2mUl8utRdh5NX41cOT5hVGnaA3uuRMoib19tQ7x7wY076oyt4GvkiaFe/f
lGeD9OtT21V3Iif+UuCYQt9/vc5jaN07G/Ivjm/L0bOv/jh1TWxOXDBoVHota0LW
Bxbs/KioGwIFAhY55RZYhru4KPbqKnIpuRLjfCJRGB/xrRTPtFLTRupun+FAzQ0v
SUPKW2VXd60D17voCLBT9VH+nc1mKuc4ts4SP5D658kw08BY7dALQYpLWTpPSEtv
6ai8SXglo6VBXbS5SoCfBzqDngCOTv4yhw3J4zN0HRPkf4TDEK38B/9Mc9foaOKG
mtVDx2OxEF3ScQALqqSHdmw6Q1oHG1T6xkhYLONCVLEu6kbL5cFDe/I7tCBSHxm2
zopYx9O/5DLkTm2x56mFpAsAOa7IPX9fol/OdhiDKn8m+ZS/LU05ThEEfPdCxPIV
mH4ivQcyK6Hu3Q+H2SKmECbmyI+ycaFoqQfUvalid81lcguFgCdTtxLpqGrOZTKS
wzBKN8R9aJ9S6yq+k50CEfA4/4brsHTDJQ2DsVXz6h2uD2UUWGPlquiVpWxjnd70
GgPL+HYD6+CkAqMxjm4MZ5SRzcVOGZzq9X0IHhHB1/MlS2/3+WzBpaknT7AyyVtG
KUXl4RdBgwxPZKweOfrWUiPbi+Mi9frMB+pdHOTabNljUDaabWcjUkSM/GX2UI/r
Ou137IvgYYruPe42J9Rl/6+t6YSK70JvoD58OvQkoO5me9nTcRRQWkNp8WFIJdbh
wAuxxwFPTQwUQsG+t9tkaM58oqyKZcVuXWWief2E9jIMzSDG25RRP8pJo+r0UR2Y
DIBIRo1AyqfcRGTFcPsamA5MsSjw2VbU+zseAZp1XNAIZlgVmQ8h7LUnOsglp4QW
ts9lMwBHDvt9lQJkP0wXSTQjEFohCScKl1WfF7ndrE35PAna5h5BxZfBticBO5ut
wjyJJTNy3iVk3K7Sb6oDe75EsVooqpZqX/P+NDyXbZBsPlB3LgNm+gubLruz/YaX
3Ek/vU/2CjAJ8sqk6gGSlDcOAUpHtB6z8g9G0mRbDc5kO8fHGFDxyIyqyvDcFCbG
L/nsZz4FctwKg3CROSP8f9WQSMXK2/FaNVuPoszoUp2dLLCcehfNRZehYuxAVdME
0jFz0YZKjhBrqcuegOZ/mWbizSkumdOqWdeSOuDkGdFGkZuwNwwcFQ7JrtaZvWIe
k8HOrLughKziazGA6ounisRGGeHRUgMs9FfbvAfT4s8rVsZ9j906KLFBuZw4/G3C
0q87huoliF3WAvH69rS7WZiCpRBDFKrIny5m6mfN1Xd9l/EgzCRFUCA7mjRmqPtH
UAN1hA75QxpgVBnCsqHEohTMsTuHnHa30Z+dSSpOKpbmNDZxvgJdEzoMfNwKZgSS
deFv7fOzUJaI5rZv3/5cSaec30S3m6GN/BKHrWwWPHlEHXD1+I4McaysXGgcEN++
2uatN+PEOeblgGnnzxnT7wSMBdWSoO0H+o/+ACkOLzh3R9pTHI26Yoghe0imaYbG
/HN4NzUWE/vBa6SFgpuTU27fI9EMBg9+tbbW9JtKv6EsgNNWkwCrjgyT+JgbgiGr
usC0isptHD+OKdMht2K2btdO+a40FehFC10Rq4BkV8D9u0heRROdjXOFX9xNaWeW
8YcPn5KuFluahKtJgXDKRl9qXv5OLRO3qfWPhkiq60jTy4AxrNs7alYH2TL5gZMi
Rs45U0MrcBO2oKmy8r7GaUvU7L3f62bGBvuT9opVAcFsnZIJHj8n0djc3o7sZH1d
2j1VEuDiHgbMGeMvys5wQaALsbQlFFU4XrfILkhtYcVd5nxatevCytN1I0MSzwfE
+leDvUi5AsiKge3Mbvs1jb/w+l7/yhw2NqFiVOCDWJP9f0/Thn5jW2sFkRMrZYrT
MnJ4Kw5OLJ8MV/IrJtFZME3NPUImALKCRogUq+/Q3O40E39QNBgH1ahvH43LFbFR
fOKO7Fl/415oi80gJiSUR1Nn2N//IWOEdosFRJFPTPHasj18jujDhNaI0ag5ZfQL
+UFKZ7ATvE/yHuETEyJgrLIW9TFAAE7kao5IQyf4l1Z56Zwk61qqmHIiS2kI0KiR
Qk0xMZ/YhL9GJYe/ZMnYVX0MN3YrwNljHnKceDnHrgzFPr+YusxWy8XmSMS9ky2l
vtFHH3lZT/Y7eWltaikA2/4z6cW6RGe/F1STxUsBN7NoRC7znHSvYK3C1P3ZTZNk
9Y7uIdpWhP6W1PLUhBbXkCpUDZxxm5zdA6HJAr0GUEAH4WWFPEUrmDDLrD24RFYx
NuThpqKUjmXt5zqH/ZDqZrinVCElKqkKNPzkpMmsOK0WyaU7dNaGOTK9N/2xxy9N
Uh8Kt/mkChRppmRX488Fu/PNFti/SUk2Z2XTOZppmpyd+eMzAcmPRV2stPNYDYnO
ccy2ZFEisCc8hBpq1tHWJNdg01IhLo0jhD9yYD4DOzrflVk2OAr5aG6tPCWme5Z5
LSWQw6bLb++nF7vo7vNzbvxEKqePZq5znQW2J6WkDzmsrgOZt0rOCX586Rr0Ls9r
y8jUhgsAdlJX77jaYnqyGbLqNGC0lTDdETnJqtAP1rT1TnkFUml7BH3gkp4w2YBG
wnrN47r6UFJTJaOfnj1TwqJ8Ko9njT5Xik1VwiK55NswBI4x6HAcPIxpgm1X4aWD
QZLeNnQK/9uCWt4dLH2OZU60kFFSPk9NvI6Npw2nTzKmGFfpF8Kx2WJcg+xIgq6A
uDbXpumaRPBQdGBLuNJErATsuA8mRK+VUsETaW4AtMoJs6e7J8x2Eaz3zgsvo92o
eD/MSJ/Gvg8LPuuPOC2pYtGh0nfPqNs7LA6z/ojgdDxSX4u2SO5fftCMh6CEDOCd
xXBBmoJLAcksCp/GmCzhRH4H9W4lhsr1BHW6A4g8aqKV0JdUscVAYrHP36W0+ilO
YtFpV7IMRnX577Hh3J8mXtgGfjo4PnJcL3kq6d3geiKWMjeuxrY7bvtD7igcfiQS
85rLCZSUdmgamtlbRQ0zBqD4ekUrHO5clu8mlyH39ZcjrUr+OaLEua63mWf+O3GD
KXJvUQB6q7MbLPlAwqIyqdky/IFLigFI/vBVDC/2HN6MCA+ehwVWg+60xhIXJmxY
+a7x/1+RkPXhiWafT5UslmAEmKm86m5w6V8rCCCy5fukwIYA31JaIpJAXxwh7W5G
R5fmBMnA+OEYXGjSdvlVQnrPoCPFhsJAYJJCj4kEzhdGcA75uPUDxuaXZiBZ4vj5
/g6Rm8mvf7Wby8W/ljQYG0uYNJJI8coErzrGEAk4CZQAs7J96rDJ4Zy6ot64CAA7
eQbuXxHNWy0Ufh2MULG9kFu0AiFSy7cntqSNETVTaVjwW1Nt2q57AydoD/w+g5vH
FxZEbfsT0q+hx2/eERXZoAgWTsAQDEFosszTHBWC0rX4sPO7+Z6v+2V9sTu5XDLx
MP1fG3tTCAhBw83zp73R2iP4exxkQWb6HlAYdFIiglN895P+Y6HNOmJaaHoR9eW6
9kjPF0HF2zJo1QR3roiiDzbWyvnpP4OPazU7wgXO5nMf8G7GjgrAdBpzSlN3/U/f
ngrUyZwsByQpiYkQuHOIqylRK8+qeiG6xlB1D/Sj3epkYTbt/6vG3KXOcMWrJAsA
mNMolzdC/gpUVMA9ib1mARDjoD631gwsQwLfE2sWU8gbLeWiQCKfk0gHIew4p6AT
q2Tqaf2X9GnsrMGJNYZSbzARjpcFP99FwKObwkTu71JX3JCx1EfrEU8QCxsIQEC2
apNlFrzI5CYRVCja/Z+Xw3+AY/xf6DcOvmIwhHQowSRG+YY3pOiIYH+ratXt77uE
ukkwf/nBvhUnK5sG6G2WyLfeOWraQH4NYUN5eQhEfHZWze1xqHPJeVCyPAiV4t8D
UlWKFOp8eynlUrBfun+2slgZFQPQsBkWdHOPp15P2on3mDiuSdUYHpFqivvhFPzh
cUgIFBHzG8an4vpp0bqt4JED5V2JW8VdrE1g/kvVbPcmikcJXGZUouu9o1G5fSNG
4lRWDJ+Np0WkRXaeNHyS2aLknE6KMlsJGoM/Z5eWsGEYr7Uzf/yMC9LNZcXWRaUS
5jnUzVveD+P9wqcjO8ZUH14h6daextWUgkWSjXbr8b4Mdg5aif7ijODL6Iz558f3
ypSvSlazvlHfK6o3ikl8yl1pwBLWPPeKe/sq402iHPlUq+90T9ey/Lxpl8qbbHha
ml5K5uJ+/+nzzFgDzRWZrvqYinYGi1xYWhABxsBDeVw/nFww0XMj1Uh9RaYHj0kZ
yyJPkTCB8uyYrXpiKiAHgJER5JCpk8oiJuF89vWgRxiHlP9qyS+O4oJIVyBs+KFT
X46Xsw5YRSJkRcNXmiwclVobslRmvWBuoY7ozwFrWQoQd2blVoohG8UvjzJZyfut
PGG3ActocQ0D5Mami1r1mxBq2NS5JExiL9YN1BcI315hktj5cev7+PNrNNyGbbej
mo5C9njWypYt9mox3XNshKD3RLgL8m6jl0vu4YaCzRprCSycMPthKTZn3FRkuPGE
j29HflK4KKA02Ne1rwwxCimE3Am8X7B/xK4YvFCADFY5DSq+0RcFyQFNksdhr3BS
6xpbWQuru3YuHXZSn4ppGm/vWJ7N1OSawAXZjFReRNm9UHy3gxzzqDX4lM+7fLtN
8/vi/imWba53BkYg+sLfDChYKS41ipMX27nuTeByhsyct4t9QYM0lY11UiaYAtmf
4rIP3m26e6E+7koljxlHnKZyp2+EIdYnH7hgfGODRwAkzQOVfSBuB2221t6jttCQ
5P1C/AO6gWTeYuPJFDO+Q31Xq7eNhjkRm08Bu9n8qT754rSiE/iGNzMCaEh/67Wq
LseBjw/3RPDmz2Q5OeP4MHF84DDhAixcEtZCQGL0XjGQx9zgTqw+0qGw59NxeZaZ
dLDAaagGtDnB30AnEJcA+c978bXTQT8WB86sAjZG1Mu4VS4qzdB2EuRjuhyMuITC
cEPaA+Nik1vLJ8hwho9yjbdM/qtFg0QMD+lxVPWMrJkuQRVmIJ653IzQEm0ybkGz
zickECqcb6aGW8j8sDlwPqC9dd7BRRnRfaQn95GAOvwsO+MqxFQhroFWjv+2pXbN
yhzw6HUH64Ak77VigQbapT0GYXCXf0yV2CFK9kZRCUH1I398MN5QgdUwtimy3+hZ
vV1zS9ZZ33NJhKhxy1iQUvDROCw73gntbhA293e6TLu0T3msgSpzzY46s9rtHfIw
gu+FJRmc2Kc0WDy4DSsuPc/7hkeqs1BOt2sfFZTavXiAXE80GTgeSW22PdtrHsW+
FFRByaN7/f+Nef55t6//mDqay0xttkYBOdo9/WTsk+AJtsChcZnZp6SetELDanGe
U2XvK14EILiHuAdFOc6Iatuc7L4mKQWfUOSr81Fn51J+f5N8zgf8SoxRa7vOCrnz
vNy5p5Oua5pQeuPsUzbkWzKw3dOond5XkjQYMyf0lUUMbphqNQcFhCNg/BBzlNCH
AIzRoOKnBHZuVwsmWH6fImMr0+20O62jmSaEyKW3tvczYocNXpUhR774Raxb1g/P
9wQQvQjQw+110OPrOuFaLJThtNo7d+famunq78F0ludw3rG+UE1cF7TZaAMOL4P6
2T3CHJiYTWRBVhEukqQNsNACM9id2iJvpFlWbE1S+P08dKmo43uWLCUu7nCul/Ry
uSvH7CHrVdfAxHsyIyLHXg2SDdBkdgqPumYdSZCD1mTOFmI9gbDjfIdYrzV+RF/Z
JqArm7IS06JUJMJvH+moeI5M104uju2dYHvKNRDq4vKNx/6NG2R8y2TOEDydfXWy
IqI14P5WRxaKLtX8V20mXLG57Qrjr8Q3/ThCblYh1eWghAz4Fv3D4Lj4QP3LwQYY
zRTXY0A4AcgQyVPalQgTt7y/cirfn85K0mVoZhVV5NjvXmdOpbZp3cbL5b1aGn/q
MP2btgFX10iYAykLyr1OFtHko2ZPavVmXuqr6Yne3++q40Tng8EjLi22v1l26INm
+bXyvuUv7AU257NrjFR51xZjlKso6mCyi+ZiV6ohYRzJ+RQiJ3RrXMBostRVjmq0
4DgQ91Xrie192pPMzfHXs0SpvvsrqhbHjcIX7VOZPxuSLRS9WFiir2easfY7I0VR
41V9LQmhQdYYpe8H0o1sNAf6Jxt5IxPgileEapqyjfyPgt0HeyXguPDR6ZEPhE6C
nTN01Br2oNQs186UUnzie2jOuUasYjcu8FLZ9FceYpLAThMiS5g9ZnYb8FzMKJJA
9O34eeUHDap+QXH4QdyDg3xVtJvLj4d2+AhzSoQGtHI3uYS175XdO8tsjz6lRMKs
9xWWRTCTcpZjOmnPbxOSbwOF5m6VpHNoV8kyEzJ5ppxa4Qqn/S8So22hUkqQNzDG
JITKqgh1WUk7XjZqMRcLhjGvnXlM+d6eUVzTZdfT0byVEHHhJdA6+kZY5NL/u4UV
zwSylvHunjmHMhjXHYajnkTeSXzs5Wj6C+o+eONe4KOSSlClp8PbWSQPXOQWrYlw
nYH6hw0Wg+L/RH4JG/WW8gSdzGG3AuMBeW0/xOU2P5Wsn7siX5ZZm/Le6yY5ZNtg
6kbgtEp8/eYmBZmgX6NdFVyA7G+cRe8AKLid7qgkwiXfVYx3ZWAI6Cbxhji9UNZK
vsH8m8eDQaEHhwQfsPG32Qj6Zkt9kFY/eZ1knGAw2zwH+sF6aRZ+nqtaCvhrTDF4
eG2OjydlWPDU7SGsj8f5TWE4B5nHHYnabU/sHvvhAjEjAxBeEpEarRF6jbiPDzBc
z/QvEkNF95Mtc+zIGhyidRUT6e4C9sYSjwfkFqUTH8ZlWv4cgFMkC4Fylt7P3sOa
0WznfvL1Ruszdct/wH3j5oguugKVks3LGpoSrqm/2mnvhA4DnxEIemUcSaBNTzdu
oFybTK62bc/FDShG7XuCcg20/PtSAioIQb84uLaDSeTrTgt2D+FyVhLWyheFVrFE
aaXOJWfd+HF+iLaZbC/rycLJa16DSFM9kce/6SCjZ4CgOETVIyx+MHIWfabTkxs4
7EiZZNA+rXTsN1uz4W1DsHYSnADjebxRtrGdFzcnGmtSUs0PPcq75JYwK2gi8k4s
F7ed1eaS1ZsPLPFWEoWSbzMP4rHp1z/LAJfC+dF6gmX/4HAbsPyaIScHlbv+Scs+
K2YOTnT//A095yuBZjQVh1TN3b4OBPHclBNzfIwImVXzpVU3JG+Ysr6U16P1OrwO
mkY+oI5uR9azczFRMBLtSAIXZXEDAdpYUngKQQeD5La7bMb2lqqM6oF5aN35CyFI
8SwudPN6mTA82wOrAncmeKIlM8A7NDWND7nC97Vw8Cpqgxn5ixeOrsfAE1wF5yVF
RH6WvmOkkNxrq1MKKEnO+wtpmK8+MGhgtozmO5XQD25zkV1XrToTbB+avqnjQXYH
MXprLMUY0Dx3S/xl07X3gso64706PikaUWN0MBS7mLRSDLRW1P6oTpMwOBGH5oYF
Wz1KrClRQ/G7DyTAlCxABK6kWUuyD7NqIeJcefbD4qF1FCSqfaF71iqKD+8mA0VO
TFF2OCToWvX2b8vpMd4dsy8McHY37qV+ty4ZkriBCXCDtc+ck3TqewMpdxn5YA8N
yHf0nhJYow1vfkJXUbHKUogVBBqlFUVG7XQJuRFzx2Hbi+L3wn6Cdmp4CGBy4gPt
6iE1HG2xD14JNDfw5Wq2ud7TeUxCGeXDhWZ8H5jGFYs97aMU16SdXWTGBsQHK//8
UqVWEqOhLOZ6EjLiRJyNq9K8pzF6wJlApEoUbe6zczBHySCvIONz2nRIVP8Ikz7O
YX/FST84qhK+hzrMZtgPXB/u4YUI6TLlGZXeH8iugohhnT8gPBy3ApHWGtBIM4E4
CLPMJIPgkp00z3vLEzHEATbPzWGjig6x6oTA/RxGfodbu6BU4Jfqam3l5vdML33e
bOaj6LVeoI4WGbzu/vhYtfuJq6G7Px1VhF83qmuWQFgRU7cc84Keh7PYeFOZfXVD
w6cnN0sl3FT4k3i+L772AFv6CAJDjo7hLNUcpyVzOy7XpXaLFWr2I/cRBjh+m8qY
c7iw6ilqWshlcZybvuH7gJeFfzfskR5w0SAlkpFAFkVTLYXN65AnLtH8qlp00wdV
H+CIbFIn61fHES15uu2xlDKRv6jujQdVzUgUKMjdOYMy1DgcNIaWI7CdH9WHljim
QUBVKqya2TuXJhz03S94ADPV++YDkjwlOAGGaCTomCu6/lZozo2y3pgTjsAxb+tO
da9fVARuAGN+OoKVxdeobAls+0m8JGTzWa1gqHUNJIKCgh07h5WI7gd1NdKJ5vRu
Jv57OqoEelLatugPrigZX546D8bjhvx5nC2GR9r314XtomHWaYZrhU3qbrdiLQNG
1qOTD6rpvSeYVZR/IPSA4ZVCsEXJAy8PAhbeHjqlAkqxXcq6TQVH10huVVuXlvBD
fuImJV2C56FdCp6J/sVjJJAQHghPSdH051GYra+c5Blqmj+TXPU4mx2McxD9FJT+
UIZDCShbcc/rZUeqn7I/tlA0qGBZPeADzTZh+P9jas+2SwQyAg/6jBt28qaj56xG
jifHrh74rxQeG7OCx6Xb0PDqfdf+XQG2TJWJ2MQL1tzkzit+FA0fwEm110tLz7kA
7AUxLORoxLMsuOUPkaonx7EtAn7NP3sFtE3/eVkvlJene/8OTQzfmIR5DYURdLom
oAgvL2fFav8RXkB3nhm987O2zTjGATxm0aYllAT8ptm2YPSAHMybIY3s8tC36m6A
uzQsAbU7aJ7oXUaseLewSkrSgfFlK6DxYUG8Uw8qPDYUCOVNs4DeGUgy6qaZdHTx
182dd7epcVCLYjkQipfKbxZPskSFeDgBkm+8JmMz0oKQ0AWlnRfMAlg/S6tp7Crb
n3QGAzgq6I4M6Hw3mzI8fyhlIs1GVLMgkOR+n0sLjdZ/tSl+9VjNAZtUFGcNNjRn
svV8xZHdhCud4hxiESoemP/Dc6PuSD4qUq7ZNIG7MMV5IaVLiWJUwJGCr13tVNKo
KXi5mi0Lo2ufayxKiYdKoY7ezYauLqEAUv6tbXUnwQolg2GDPQ+o704wOpHYfDCL
eLDGdRlWDVnEdWcJW3YjINibNskMLVoJ4lNxlAEgy7VBcZlBKCYr1DXhgsI9NOkz
kE6Ha+ffL0Dbf6evhYv48yN73b9XaRQ0GvYldnxDUMgtf6hh3VKLgqqTwR784Lx/
VwHaXlqkpai/gna4qfcXbzA/J+rrOcLzF5oGPhG53DyjOodU2mrdIqUU6cAksg/z
aWQX9sHOoTeYQ1Bkc7O+48e6Pymef4HZd18qegh49EeFpDv5/v+W+PaOQcbFsJIZ
9QErsX1HjTF2mNRwEnS9BtcKRAxHTLHkMNHWsPfRP6tl8jvzRoh8c2hSPFESb850
pcV5LZT9uk1bGZV0r8AhQyvj5e4SyY2n9mj0aUdNHwumKDwUQ/eMvcPfCC6Hh1fP
kDAZdY8S27s3Lsf7MYrIfsHVrAvHMXLy8TcgvUS5HtFBlNfvj1ZwhJ1lHDWxQ9gn
ztldrCcDjZV8ty29BNijepY374bLp3P80qLkCc/aZH7LN1mipCEp3eSCvYps8CVw
m/AMXIjuWkJoCJ7EUzQxoNvQf5HGbFqSbVPkXqGoqrgLCVein5sKxPtS18Yhv+CT
Haae7K4swJKM8JyF0yhCg0lbWSMMZH585U2pRL8mb1PUWr2FjmNN/2OlAjcKFUBY
UyAkuu4FjxpsX8ptRv+emhi54UGKj064j7CaqkVZl/9oAJheRFPGkbIHQHmNZymO
k00eyDVo0d2dX63MlLVnurvW4hv3PXQ7xJQFPBPrTkf8LBLpT2vBJgcypkt6mzAr
aJXH4Jx6AoIv9RvK0B1IaPdlB5+vuDXQJP//wM+9NLIMIjBFWKDR1jVYoclng5C8
x0CFI/NY7Db7yNrwjjjeefr2tCGHL/fPS8q4OHHUw00MVhf+rkUBsIY0CTQSqIjj
52Mx8Z+JaX3vuCNKTRzzfmsHn5L1krsdOyeVRzpJxnXF8gWealfSSz64iwxpOK6S
y3U/D1FiRLSr8I69m0DoWw4lCGBbU5QvS7HBrfD2GUIJKLs5tHVerELEJ0AZj0+x
y/ESJ/YYUl3TxL4v78YA7AbIYCX8RZKd1CONOJ1jq+NR0V86Dqql3tPGiZbnp7lR
udILHFHNVUjUk3RMjgSFFeZM/bzYIyDN64cLwxhXmePLvqXdwz+pWzPZr0jCx9Oa
2MyjPhc8snMBh6QdOfiYA3rbU5cLJLB4FpOp/nhfGTx87kp+dOnOGtqVIfiodX8c
/DBt7v81sR7Si/HgSMyd18tYzRmAWeGET9tLEeMdJA5iHw2NWPtyKsvDB++NWjNB
3lXZPZgVDPyoxWEMjlulKjKPzpu4+4nVT+hC0PJ6zf47z68qLIsNwTNjzZ4H6Yc+
cJYQlacaaZYeFF8DpdhvEK9aPxEmatytAfhyLuK93OG3g+WSfqch1mHdfJ8/WC9h
FXgE22+h5wygW4oFDlizLmBoottlBd1PY3rLhuW71AeWQn47jP7OjXw1SLk/Ms1z
4YS3FkvP0QLdpOmpByES/ZiTlSYn2FTDLXIzHtl/Y0guLRkJgZF88jvJkjc5HhIk
wwhxc9JwBAONaSfyt5UWzhSA4rseuQXyyu7qI5Cy/YKsuThn3Snyr7cSCss82EL2
3+FE26vd5xnoJCRm2fr08NBQHgaygiPrY9WAtRTdpAIBi7RD3Mk5xDG/J29cGaPV
Zu2ieblxKnzanHc6WAzQTVh05uKxwAQqb6eGxP+UPEt1xTAmXU8KwwpTrqDhUZKc
pjX1mj6u1PJpo77AR+nXfDRlX8OD5AB4dsyUwmG8X0nSo/L+hVfBhR6ndleSBUUG
yItoPgwojrguRnFZQ9XKXDnhx9BxzxP0ucKDHad9g3eUmZuqMiOgxid4EHH4XR0K
kiJsduJR+Sdqm2g+3IbWmWRaQnNBBk3KqCQGSQmrWnoIrUCAfGUtPNNDIwAlf+1V
k3llpJD5IdjNLIfOwdA5qH9SIidRQM0lETMsJhxtQAKMp1WCHVIQd+JZvjhBZ+RH
vlj/hC0rP7ozOQQDQzdWMpF39rnr1UTIyXvgnYftK2X4aegxp19/Hr94XFGAxw3Y
4r8pb/bktN57JFlxsD+exyAogGL2oh2pCMhbL4f+AjGoO2Aoije/Oy9ZP5Pgbwlw
p0QndRa2pzudZm78GnlmkuRCUFvYAzEpKcXpeqFhAs+FW6mGtx+r6rP+T21MNSFc
aeHamMbJ3ZFe7aXWBqZxeAhQ8zQuNfj02PONp6/tJyagmTmcSJx9RdXs8GwBBSef
vyxoMvAaeqPWuOYTHgezShuhkWSGjl+52/7I54eNO2ntNJABSUth9Jy98TW3BRUe
DyzoHk81mfAB6Hh/h4Rkw259ljVKZrRiuEvGf0GXF4SZ1i/FNKOi9vQ6Yblc9vfU
A8KIiIXKjmEgN6rY7EhpWDLfa+8fxwx4t7qfGv2LJxzPlKp4imeXJkYxKsfb5sfI
Qm28m6KYfxfmhwUTYSSYSHWVUqc/Bq3OkoIWMxc/Hg5bp7mRw5Fbdn3JfQSB59vV
x8VkzNgJvTc0P/7aGfH2tqx4ctNxca0YWUhWOHoZDUVca+66KCTOc3PkzVj16EdN
0OlEPTH+hTVpNGeR0nxse8ShBHn2IlwRWEytUXEJwTbNxap5+N9yafQQ+K0XsEFo
Dnek/Hxzlm6JIJIlyrQUpiPU8HwjpXA74NUVlGti7No3+sSVKBG/HSkfQcnDwqWF
Y72/buHqXCXOOcrwheirowO03RIedqAQFi4VatL9kIkuqgg8hE6CpFgkNPoKnLc4
Nw3IPhrziXGkVMpchQPfHhvcuB+WMp6O+tkvCpEzQv1miV7/WlEllOVERx+AM62L
fggy5CWkBKoPie/hPGpAHnssp/uTnDkg6OiR0Y6xD/kyBuU/1dkvzVjsYU83I7h2
fp70S6clxTmUjnAiuF4GJ7Q7WLcD76uQg9xAJlPjKGkfpwe4efKMo9g9jKic54qr
St+au75LSYlokVYBFwl15z4EedoYGnq1B4m7OqwyxzTuxv/jEFsFLcG5tyT89ewu
C3x1L/nkFwE3SJjh7+mhiyzdVsGOx6M3ixT5ZN8k6+50DQbrbnFCrwqojOqA8OA8
7GJ0r2uL+xZSoBznvGhiBUg7z1YPr6O2/9hBtSrinm5Rs+DEUcjow6WbVdo2/qkR
Fb/Wu5MI0Bn35CVfLbvqtvAXLsavWBN26V+ZbasSXLrLFopBC2NU9SPIg3ejboiA
XP93g4FxzenwUMT0yrFgwmc/hciyYflVzRS+MzOgrV7odWHWqBwKwNnRVdRQIxQW
IBJLnK0kq/Nqj0wGAF/QYO1lB70fwE2pbasNn0DbDFgVCu59HbUHRYydy4ZNuNvs
ArXgnHLKZHs7nly+R/o0AUHAuDTR51NG4o3As2QRAcRO23nmRHZ3NB9AbQMSVX4y
nVQAYbHU7EVCkK/Ziic62M93GxMRq7cDFR7utJk1nWCc6Ka9OVu3ldoZWrx3B5tD
XP9xQUe9qXFwZBApTWySLjsafDFM/4GNpzhLQ/2wM1GB5aQAcrGUzDb3NOpOO+ZJ
3pXJLnoy57a+DNUOmYJNM3R2Wxjife7DFQjuS+ZGP71tvvSz48eQHq1bwk+7rjrK
afBaXNolGvQ+LQ6+T6Ii4oWhsMUKtiBhHDz2Qj+WK+6M47vyWanDdifJfvomGeYa
RAiyrIYDtmgYcmg1qp+TJ4kDHNceiU52bzbxvWrGpHL6R/Va2uJULAT2jC+caqYW
MpvArII7ekH/y2y02KRtLqBy6d+DYibZswce/xxaXCiYYW1QKS3QfEpqa+RzdMUN
ld4FQtf9IVDP93tPhX4E/Tm+Tk9V8moX+SJFg6xnWbZq9Z3etPo0bBx8lOGAyrc/
F+7KqrA3xa8vy7FZxKGVb8CzNEvm9VqizfABIfeB1XJF15KihFmBZ7ttiZkniUdC
rc8UN6zU30bo/BS4RNxNuvbF10uvlWJR9pzGD77jDFPE/QiuH6V7yrBBIB1DY3h4
pMj4DUoqtgYTjxZKfmFxvhVVPXOm1uPS97ZmcF1fTwZD2X6HC94zJe7EuhXwQuDj
XpDuYBCKHt+HWTs4eulDvg+yd18o5hLBm5aGkmzolKHBFBk9ecC6sQSYxOQzIKy+
I7nJBHReJULrZvX16u77dmJ9LsThZGL6dUspMd5ZRdSU0yPjOevkoUI2YrfN+rho
szhbPBj3lH2H0oAe52KKB3HSHbZMFCswWcB5SlMqaCbP6LHLTfL886sKNbLDWhNl
iiSGD2b9XEH7WQSG2QooxwRIBPhnlgJEBEL50cRfFodrQl01eCYWaFOFeLqMyYmg
gR5kma+xS/+95doLmDLOG2qh1ruTjQHrvzEPO8t0mClWs9VYhfUul4bNH1xUQ7Iw
Am6i835oe7UWivAVQYatWVACrQqACwx+1aNMkXEE53OqkVcySGUZ2+S7f0htqucw
fdO6Ybeeq+oztgCBHiTNzm1pH+BxURjFoJkICfyeLxfw22CdXPW1zfywYzbN2SZ3
CJIfNgCfhqL7/sYoJdbgqjyxPBbT+VhXqCKVazJ8kVh/Y0h2uvwdLgW+dokXQUgn
e3Gz/YAmZtH/ZP8LUF8pKtTYCiiLkmjqUK91rH/YuUT8aoYY5oCI/41MJCH/rDrx
dTWosJiBkJNvg9c2h8SYzf89LhHngdcKGsFhlqKVg3VT8RYYPLw1CXsrhCj+1B4l
4YE5/h01epq25BJyuBjlz5xPhdrG9lDxLhyzm1Tf/LqDi9Kvc5zu40O6Dkc9uJBM
AFxiUbGpJPsc6I53BxnlhwC/pJ4iGjndh0OZAdqK4Fgi4fdle26h75YMu9niYo28
0drZduQN6K04s7OhO10vxr2IioWPK19Yk2W2dPDqgpK8qqg3MqwcZEtAEMY9VPSO
O6Sk1YsADmXwFNzzyFXWcPoBK80pxX0i3W7KDPIYGcNnprRSkNupLFL+ixcXciq7
HSJ/+pXBLkMmvSfyrpN4ZeUgl+pYDDNcG2OHaYfcFtA688hDjeELFWcZAD1DzDFT
y1wbJCif7G5PAoGp4LtNyww7JjHim+JmTGTXaUj4BLy+SuR/fJBIKa78Y1bJs+xO
53Ncv/qEaD4kTK++e4aB0c0IXOo3LpIwOlSvInlhx9nxZS3sUDTFWg479FQBvgjd
y3ekh/iDHNHCApGJc6JsITncpKmeqr0VrQTg72GGwPQwSk68DIJPvVdVoRYHZBUm
X6b8FJwdK+ieJUwxYHskSL0UIYBPkjq31T0YF6aj0C1lQdjBgt0oiy4/jqEW92qv
rVSA0D0rIytWKzjd04Ru6I3eyWxGx31GZhx8Jn0JXKZKyljeTOXo1uzuOIXBUHlz
suMHCEwYoOqU2qA1NBpEcwf7YUhjVHfI6k7idfzlRpRIckIWNye7iQEW83xVRhrf
UtAfqVBKxZdwH1q3KndC2WXPsQ4GdfivWa4ZEb2CyjgTeJgnUydK66MqfJDwvwDP
k+t/ZAhOOPVyjM+tWYGppQndN+UUViUuFfvh3mizxstritTXvRgU1TJANI6vk76l
F4PWvwdleiYXkOAY6AIXohWCvJspECa2CLPQoDPndm12Mt5eqbwyS76GYnKOo6LH
pqG2O43von4cawzIjN7+UjnCw6bijnFT0uwFfEgiXG+dlE4nt95EaFsmMDBtHBGT
6hBr13r7tse20b3Tey0KX9cQ2J8reHgxgJs4+L52EpKWnIwiSc9OJiZ+c5pzuILZ
sWYa6lmZzX/7XlKnkX99huqJcSlojvGEF+RtVYp6HZATuexhBMmIV36sKp4CmaFi
7KO3ZZxAqH8Lqet3jgD0RifDuhzpX28Zk8EBvc0mZs5Wl5OY+NcN/9msf6Hn09MN
GwNG1bXHRJgW3kKw7n9TmmoySU/OvL/q6vV+l5hXHh6uIrhQ2B5Fb1AXAR3iuYuU
VzvYallFX7MmN5NsrhfHPtqLngO2FqcD64YrWBiWwF+fg5A2JKRLSf9wY8qpv0Av
3qj13yP/v2KsXngIplBR/6yeohGEc2+4ymz/Va81eP/Y/2kSqzgoOptQDn2lt0nU
WZSkJTOq6HZWfhM8a+o/iT+eYxQBdpY1lQ4nwqPfQ9ihZKTi/4JSW5SDyfHoSjr7
GHCUteTLq5tajdkW2EBC+/DaR02OT5j2Q3Xi4DtPEirvRnJd2r+8nh7JPstOLb7E
RrXqXuArI/VLWfI0/QrOUpYqqq1tj/65BarPEbH7gtCjuzpOFuHQ95bTQoF3kiBe
wlGVaDxf284ad6S4lvVtCuFoyOtFUY2g49ojj4wn6QNEiYPbS6xc+6eKhmULw0WY
XdoWOoxY/Jp81PmVtZ4nvSWmj+5yquSS/OTnJw0kbTofpg/KiEX/B/5EP2Wr9bCM
tOjOlPrV6Sda80uugmLG72BXv6Ecr7nNlhFNOaGFQYaX2q6Vis8FpwcMuLXHoovm
sdeTvhL8rY76IGBrqq3ihCqcl4vSK20u/GQ9AJveFC8OJnN6pD/T9xxl66PthNey
0vOngSObNBFW+iENqElST5GHqp3KY6BcDk32Nu/5MzLQXRanjtUcbczjhwEqElid
7oIOtKMsjtmFUXjSf3/TuHAwhrVHs+sfQsPQjW4OfcEReM4kolhoCivYK1zBDEB2
v+//RF+pevQi/Q1WFW4xQt8cMmQjmqwI/9Z+945MowZHjoEIDEI/NmYjmZWReRg0
JeBTaOLThXOS1B8Ru457RYgpDDlk1E6p2YsVPDHbp5URHDPaQCY86EGEg4yVjnPl
Zm4GyV4XQHz5tj5k68TyGaE7WNGoqGWyis9DhjiT+z4QjfricHud3hnjschsz/Tb
Y/tv7NRJ2yb4AB6s4l9Jx7Pwm7qYHkBT2HI5NcixoH2AK8JBKbPzx29CcfsVJYLO
i7ypRFy3TzZzQboSjBsc+L5uGnRcTmPyOCet1etyAQjpQOVr89s7OT2JuvrkqwUR
J2xW+xKv0jcGsnQnUxbKW7EG+JdZCtzbyS1sA69zXwj6jzt0j9EvRl7nwpGp49/4
Y32TH/OIkhE1HhNFenFXmnYbeeQ6+Z/mXnhXTPjHT5Lctdpy14Kl52n1oUfuRV2a
1xHppO+cXL2lRJ2BIKTI5Dt5fikY39N8HCP8fihkjAAiV3o4AG9jA4hvJRejZuak
Rd0NIFC6g+l5rT/KnUFIDS1jHkhiHZKrr+bMwlJOWxEuUl8XjgtK/U4UCB67YCNL
Bf1z+e8kMUuANtrwMBuihlrkPnTfJK9CMm0Pr7g7NS8YfB2GrsASxbCWFkeseUBV
WT3Gsdgyqq6ybcm49DsduW3g8gpo8MZ/XTt+ezCyTq22+8bGtU08oC+DVh+SYSAc
bTGQ/h6yEwsjGypDR22pSxftllhzIEOnZfFYLjffFzm7s0FB3YtCu3mjqAuFIqSJ
k98hjPVrDZa4qfJX2Ne6KwQxK7w9bW4QOF57fS7p5c21MMPwV6r7btRJpwoFri3K
jNYmbKPqXhWNYQvw9uKJte64E5o5Xnbc1o9eDKVC0ljBxdogkuCUI6AX5jYfbnZB
CqG2Vccyk6Or/ssvCK1BVHMHhTr7y4IqYqqBKClvLBSWH6Px7tji66b7GAwLo7yF
098TubVn+WzEpp9e4LNbww0s8Fm9VCYsOHzVbiBgSQCwrv6ljEskYSRhmObqnwYD
TKOmbB4DH4Y9h2eTUKbqBt+NNki9K2i4KU0scK7ReXPhbzndfXIMNZe+nerQpS3b
rNl3qFG4pIy+JYyXRbZDPvbAZKlPfXYcCM8OtOGTa9uC/T6YLlnHQ7IpKAUL6hC+
Nf86kFlfWgUiI4Ge7Wx/uIDKx5zQhsWH/0r+MyPe9+Y8DzNsfVbsFj2IvkvkGcGV
Ell5SmGaakNAu4uRLfom1vsgNZQtpBSVUOvcAdxRmwNyfcw3A+auh8Scm2FYMMGD
O8fqstpii6gd+UwwWpxTJTxwJsPhuUW6hyYOk8R0PQxEEvevdYIVJzAH7vhPGuAU
dUpyXH84/WpqQ0Xwl+8Q+Nm5c0G4jJ73veGkyFikaYPw1Gvi7X2u7pikJ+bhcyOL
EnIXBAaIuE2/oUBHQlPX064cvfSRI6GoLjfQ2c+69IbqH33yAVHViHK5FHV/vsYg
AdkEl6sqLbnyHIViiY4KVNmkHRGFIWPBi816hJfLYP+EdjMCIlvoVqY+4egIXgWK
eVU2qeKaZulOqHtJ9W385iAoQB842wCXwrQAM2UjKcTt6MqooRywAktZD0VjQIG0
kCbxM4YuuxGPYrGZJEe3lEpaw5qH93oMLCiUkYww8I4WQ916MzW9XdvM3Qayzx4/
mUX1WiOVQSJXKX+TMdYiCtFrzA+b5UAtRugah40YeWHv2Dgi/3zK2yLrvZTzio4U
HazuXi9vIKoHx29tqqcQwKPBoBUrUKV7ecPeW3xFX7/K2P1m+tFYgESpT7/pfkE/
CnKTWgsM4T9aPDziDVaU5xQLKTqeMzZig0qiqzeu680TxbuU85l/yaGKZ9niEEoW
iBc1xLCP3SoF98DvDujJcjAawmaMce/bW5U21f5kmfd3d3g/l7lUOdtP9mk3LU9t
sB6J6iJWYuyLgJ9T0t+DOeAkJjt0of3lzZ94KUYFVW9vyc/5mAEqO0lnJ5nQAhr4
i8APRKbNJzR/8Ag/HJwqPwgQ2bEP13O/jYJc0RABYcLx7O2kn1jrTEXYBLrySLsj
bBVu506UnhAatYa7w62qCsMMrPmGTrv4mFSlMkuWiJaKvbGRMHV6GRkOodvkDQ2u
mUiwiRpcLd0Z+2vbwxz/0lz+dBiRsvh3UK20QIM4sKP/dZNpGDk7d24A4Wld3ksL
DfecrkssUMVXQ20msUSAc1RqqzpLnWyKHkRVSixL0H2xt7HUKxQzL7d30q+DE/0U
mUhDB3JhvR7FHcYblPvWssGawN/ND5tFaY/QmzpANgzCil4vanTyNfi5v3JDx1RY
ZwGqVTBeewq+WZAP1gQSwHp+0JpcUuS/6tbLIEUjfPKjDwYUQNWhY23zK8e/sjny
dFpZVNcwjeJelq0fNCSCh0lWpgErnL1Fem0eWaRXWsZcLRn/MAs/94q6B5EIanxa
uXWk3nTI22zS7Dlp8Uqkx606wrwWNN7oCpIEpAexMYDvckPqiTzkDOEwot1Pvn3e
Yco0Ql55YN7fRrWaTl1dmr673ytfVx2MARbXpBlj+3j0jfl3xVl7hKpXZk88ZOAM
/Hhp6LXPuQ3fU57JE95ooXI/3JeNZ35wsWx4jjnXgnDLIeDNdhQkqW2TfWGfIUuG
b1gKpocEEOgn+rrFlZNzPx6mVjF/fNwuZnm6QRQQ0ND3kKsNjTvYNZ52ejSCmpKA
nQKZph5NN6DOmQwGOZeYtnlP2RgcCWrQrknOmtjc7h0PtchFQ0v0LMDhHX/Di2q1
pxfAvxNeeQjFxot6NUGS+JbyLUIg0teMqWFq9EPtA82yEjEgwVskjeNk+e/twIId
ZaGQMvUhnskWmPKpO0itwXq9yrYJHbbrALCKv262p3Kj7Z4EkHBY0Ye8xaJP3/iX
W0yn6uK2pL7kSnNdEGvzN+6YfyzcHKLq9+jh3rySUzG/29AIn6w9hyuTeR1IaxEm
KjrDqj40B5l5F7GuUyynwIfKwRnGXQ/YbjNoqO9ZQKpeGYf0Ffddg8gzDUC/gaHU
k3sZwaAEXC5O8CeOKqPW3SXT/Ol2dU2MaIeCwgPIYU+069gxOeOl+U9ufhOXpNO0
hDec1U6wmAb17gaXQLr4tlDFp5vdmJZ1fqaN9gHBY3EuN9ovay+DcTS3eROsuTJu
qOKbGA3SkiaFsxTYQNPP5ktKsouApK+kti2jvOGTGNUYmWKr/4SC0lIcub8zqAq0
g9gyHA5jiLxJA22lzyu4UFlCds3i9bZwuoeSy02F4FjJGJaLLnkCHYrYOf+I2Tm/
lBRClRQv4Z28G0GdgPHONkGZJ2C9pgM1m3PpkR4fm9eA+8kvl2zP606on3kAwqzK
mKfaBrjRLXUWr2agF7gV73kGl7aDrd6Ga56ukrEwVgtPMmMVoOZFnWCGrdpMn5hH
gDWzJJLRYJcsghy0d/pnfYzStxi8fRwcP6wOWa6D45EG06hNyMAE809f3oaTXy1R
1EFRNbrNHian52fr5R7Z+FFB1h4o72atgLWBc46Au73Us7uVDnTWj9JOuLxjLKoQ
oEcF9hQQjvgd3GVK7y+yOoQf+8ZNqG3LnRPcKd+swc81fe86zdhTNcmasbBPdgFL
poZGYB7qaYtoUqnnrXQmG4+y83tFA8az2ptyXGgDhlB4Gfefphe7vtl3wAwDdZrV
Nzw2gmO7UG0/4hH7TdFO2xEXQahb4FsDtjdN8Wz+Y1BEEkDPH13CnjmZZRxclG99
GuWavbyhv/j0lEo/W/mpvPKOAS9+1szCdOj5HIahWp7J2PbQs3MnRTxXgWxgGDUg
NxCyRyHelxPAy6vVN+h4MuqdOLxhsKsy+8+vWFiG08KUllB4h2pNwOo0/x/N6oKr
NR0sVxwa/iwyQJt5bSxSzOuYvgdcwSO0hikQrin59oGyoawaMxyeKXrbadD+Sa3M
L5gqZAcN79YYFNhQ76XMeK2EdcVDes3zKZ1maNngFIgYTTwhBvvRNuHAcX9kEecS
obM4xVrfb4X9aAeQQXNBqnau3/QmNVaBof0+qnoFL5JYqifqN6XL82q+2YeddqFZ
JyuGbyS5IH4IfUt9Tczo9OAZ4gW+80P6yanO0I2qG0hFQQC70yGHZRcSQInGuJsO
KyBWEpLm2b8INpyG+bEIxL/rhHDur6L1Yt/0l7QJy9mVc2huv/1qRILmETKFzUxp
lUa6Qnr2LL0lE2cOhil2kBg3weWwVjDr1bm4TuqPTEDBcw05bo/O1v0/JLrxO5e/
vKfiFP86RbocUpI6bFNp0hNaWDLjCyasLIxYugL6KViLbgRKmzIjaTZDSQnC/WDR
j1ZrPN6AoWCezFKhDuJ643E8/rGfbIB2OK5nVarCuhHErCV2grgPijkgimIkQ+uo
qNDD+K86oyBMZSUCH0obDqlbL5WP5DaFIpf8yizvFPRFPXQKQrhH9ybzx2wjjTfF
Sy1CfdXBkIRwTOcPYch3ynwaz2fA1RvExaU8VTc3wNJflqdMpl+yY2SDrJQApYaE
V7ktdsXQ9gXGj1DUadzNX+tiJT6sGVrKqhtu4we5Svm+rNS5xLo9pDroa7gGuHIO
/9PTj5ZRFPwCm41ww7f/RF8DeSZnGgYTG3QStS8CLZ6DTHfQZi0LaGX/7lUHbD/r
+QtEFGQqf1sIhfqxUas4Z9ZRwG0d1SnUbAo8Eha4RFasxtyEHNPLSRz2092g8UTX
KIwDfCj4Aq9mkze3USE5CH+z9k/11vK/m9YWl90jCFrP820EuC/96NaV9kA9qtIM
P4QmP4FXHmne81MvzbskazUHMSpiDruQosMFowUu6WoYO9peem5/ea0r+sULLs1B
5Qxb2nyDVyFk9/TPi13t82IuQ0lWf7JeLPWF4+cecEJBcPNWPS+5NBCKVtBMGEyK
ZUVmNnhIEYgqeOE6KiqjlfZGGpnLmXXUJwgLv/GtsQaTgQztf6rGs8okQ6ZW0Yjt
UNvcz/5NH72AuHAbgxLrrMjSd/hwGwJ6M5xj/9QfuX53x+hIUx5C5C4cwi8x62L5
Lw7AK1fa42Uojy8KR7B2AXq9w32WAWJpTC869vAA1Ip1hvkt9W36q57SodSQmOhs
kLSdtXHG4LmIuhBcaCxi7nxql2wSas3mZH+J0GXGHHQ/rnH0XFrWKlDwzEMxxL/e
Tl7/wYr7khRn8sdOztXQ432SuAU5RvGzPmi/mAFPS4wp2A8cmvlfxwnwNyqgtIvK
WQK2cs4i18IUEx8/a6kQKDBhIzE066NFcsifgJ7bas9+jCDGFTaCa+raD4y2Reip
bTGBX83DB1ZpbSZcAfYeVjR83eweJnzWFN05B8eIecCREiK4ZS2b1kORrWQNZSx5
PKO8UYZlRul+R/9ACOcPBUUzPHE+4TAqXjJXyq0rnRKJ0QTeD7vzeASk86MDqK+2
TSrL2D8LkLpR/oeWJU9zlYFNorHrh1fOUd96sxQl3opvGPl29kxMMiIrNakRRYrE
iN6Ksyzl/VK6/L9+zsR2FgNTFjvNogo1dykV8nx4hO5lH6O2usfHlBmOmt1bcS9u
qoK6nY1QPewYfaCQT5Sh5jqcwtkG76Z3EiWKf1JjyQAcIcbemM0675BQKfwTMQo2
Iqq5p8/ldRBvBEzNxMejpKO5SdEpLA1GPt/zPHqqUR/zeT4CAeZ0WsbAQQ0njiXm
dcrqL/K800HzwCqQPBM44OjXUjJQtarhby7NMRh5aFufW/J0DocEpjMmKnUS4LNd
yEwr3pVdKOxu5QK2DmfBZCpKwDUZPM3Vo2apiOxwOOnpgYwjJ0etc4UNT3fcv+eI
rvKd5UBnLJDxC+jWvRfdnGs1dsR1AEeJ0y+OI3X17pze0frM1Jmo3kBNOCdGJWmg
kcU+bvOX5faNpMnXuDqrATA5y08kwd6Y/5jFwqZEWSuPlKTBZnek7EtQCwEvApwG
AUtD8wD9ktiIV7CWuQbwHtwQnCrktGuSrQ4SdkY9Ef0aM2gYnMmw+eDfIVNyXlf/
qNv4rNxrvKKol/Iz57mGRMdRrNqkObmOvffyGoDOjindMSqscqDOhsydGm7obUUF
TPnLSMtGc9a4f5DzwgZaGKqey7LywnAsxb+ySf3Ej15E51RiovZCqjdmkZES97Pn
TXYXKHT0930RN/mm0NCSks05B2xWfPvdyZ4R7pC79wzkG7HZpzyYQWWue8H9rJ+0
EdDbVzQUYC4mbXWIOGbk9JXkVz0hoXFPSlCNPsLFgvstUJ7D89u7uNcVsE/7FCr8
iH7oA8qIivzx/M24RkiQAM4u1HA8nLDyub0d9sv9icNl0dXgk2IAZE/Upkqtwz7A
e/XBg/JODgHsqgiSXvnJQusLw4aX9mhM8Zsi9zuwtTFG9rc5To83iSCbKjbGHGDz
0r7ManDMmcUjRDZhlNrx5/iIxlcunPemcrsxM2Qln15WIkyEMl8rXnr9xzIUW4Jp
D/uHs55K0vlzogQHcmAwcWN/HHSaY1to0ngah0pESjrbQX6qa+oyOGtLacWIMAFU
SMUYYzng2chnaVXJn8V1VS4MkP0BN3QwYw1rSX4MtMWzd8psV6kiuAGAX+v+waNQ
ncXqFW0ki7tYNUZerAFZGQMRD+wZSQuX/fuXzsdAZ+ZffSUpq0kD0ZDuBqeiTLsA
ptWXnaVuohwoZ+ZSa7V3TGGUv7ODuYcSNc4NU8KOSz3r6dJ5TcQ9JuflmOlJtNYP
6oc8JdtVsIuq7PgRcoA17tVpiFELQPjMc+rj2iwyyIkUwDcyBEjBt7UUMEl7dqDq
uvievxA7y4SZNeAgRvRC6EilfCCeXEIKvJ0R5ZyJkKajQlji3+XjWqPukai953CB
2mLYqZCln5w9jZ3G6d6QCMllNjAPtlcG2s+IJPS6DkTP7Q1pvoyxiBHMcy6ClUzZ
kxrrzGjny1WgumAmea5WvsSnnz70sIEYlV7YymwSixJUadLnLL4Cde3iMr3SaYZt
FVE5VrcHvJ57DDzONe8mEc6zxJlCp23mOsv6kqtRi4liVh2gSHPueUaeC2QwfavR
tanFZRJbcsHzX+MJs1Qx0MCRBF7td6swKqwCrQU971hXT2CMiL5G/SNzEPwBCois
3RguFp8I6Nsl/uY/WRggeOLZlPjwWRBZ6gNH8IhmpkNWplQvdEVG+f1nitevEzZf
vlWkgCV1HPVlVkr5nZHYTqGPagYdvK1uOb1W7Trstg2glHIYSrt6qem/OFAEnRh9
GA2j2bGBYwv87p509SaviGePDFQFchaSYdMjhsQsS29fzZ3kt6X8bHfUhchu0qGh
Fk2JCBm8TCONB/cyYi8/6vhjtUCTACX6cTypxSiLe5LtBtY67tDnD04z048qtvlx
zRiPey3mxaaD7QKpzZGJo5WHQPunQovEF/FpWZnUNxYSacG8S1M8BWEykX8h+5ZL
i7IghAYSQVxbNvKJajj01MULqLimLbHO96rshm+UwOxFc4XcAspqDIskHaLmWeju
L3zRHrkPh57Zpu0xBxFIciJfQUqaGfr+hEU5AHvLOW4SKMdNtmxk/TiUn/99giBr
TYIIFJUf0e9bVgs1Xwu2eguFsAm/w9WmoiGsF8JB/Lmxfh/kFnq65Ixf2TaropGF
RLXX16saOZlkiW6T7Yo4mu7oak1FuPeOU5Ka3jHSBWy1IBGzbBZpIxVoUM8N841H
t/yjRN50Pzir7zaM3jLAUKETLPeBoCvdAbtV4U6oPvGwUlKMpVcLBhm+9rqhwWUb
+hfnnNGaVgYJ2VsVr94XJZsi98dbXg1iZUPcHFXLXitImdMQVEnyTm3mMiEfcn8w
EwJabPVvsUOFNnn9/ul6r1z4iDkdCidZJvNYkHrd+e5O6GbBewkGEuOKOVjepgBu
I+2Raqy7Ywbtf1wqV89OrbbDiLrYg00oo1AQbN8h7gcgln3EX6w4yBTOWrlVtWAa
+FSsumiJ0OAaoN7y/b3gDHh7dFYSK0XXyWlf5b4/RvP+TJFS9JGV8bTSV0Urlt79
uuiK2SdzuV0pNLfu2MEju5K8g8k0p/hwSU7XuA/vlBbBSOsuBFw85EozluQ4L7EG
+amwDo4Iul6FHOxjVtrHKQ1F/jkYbtji15+LathR69RDFh50oBoRDP8aVG2+9Pd7
AWmvtMKVRO8l06uxGQNyH8OWOcXUjrb4D6emY8CxtCJlYS9usp+CsJWlpKqF6NDL
EqbQU9zJNnvkNE/CwKHGGynKnKSddNz0Sj2IBpUR6p7pMSc7okuUYQBZEEkou6iw
S8XKubIVIYKZafuEEy16NzxrYIhynwUKTKqBZsyIOAHbBA0jTwnEyb64b4KkOcfA
HT1x6a1OMjo4WNh6MmqyyXHtAULdp4HnhvSGYNsMQ7hJjyriFIge2wbOqr9o05YG
NIOZz6xbSEhNtQ6mq59xrH5VDmImMnL+BDps3zFNSrdCRcKip6CtGiK2zY/OipM3
ApbOZA04rSbKJ2v9joWAc9EHHUDZQNGAdeAhLc9wLdJSy3cIguXZ7zGPee3ToS6Z
EowRWsvbJ3XHdQKVFG8jekQDhFNaRnNQba7t9nFcQrrPcdc2UzjSkwu+qAFU1WDN
IqdAxG4dlt48zxg+hvPiJhrrP0ZPx1utj1+8g3cLTKjmilh0ypVTc7yN9rS4qTU3
Cmd2LJ56giP8lv7ft2ayvtXMdouXcF8QcaC0YoKeCiqU83v9qgsg+t334SYnv6er
elX1m6Y2j0LBKq4fMAIBCw/KA9qScKyFawDgtubJVVvGwd0qRV515rZqI3IninhM
g06tOAjtEBA0X3KW/3G+zch6gDjoItNWeb6vmPyiz1lzWmFD3wyfC7WtJR7E9uuC
mW05j6AGU3ihPCi9z2enfk+OzBzsX7EPj9UZZtZ9XMHdkF6yv7FNs4nUNL57G7Zh
i/3zyIFwCaKgSWJXDpyuZPgXa6pdQNRjpl/MmE4gqvy8rKJFeFS3EkG3Gf7yWF3E
x4HpNHeDlQtoBXy3CzCueCDX2SUF6gYZvs8DQn4qPEiLoP0lH+xHTMe3XY48Makz
nWPc4eHnpXxH3szNfx6gmSu1gcGjdCyenCdteSaTLfcy0pydGxdbzFmeFnDIf8X1
+tARjznnIT/2/Svv2/nonVYsQ+yXLpAsBtR2IQib5/pMoGizAarZpRVxLtYRhhqd
nqiVHAdTSOVsPxz3mf+MJMgbsFiRGpXSnuiFybGLzvrEy7JynvxQYQP1wm5HU487
haJ8OigPkceU/62GU8wyWE0A0tYSPPe+ShSBrrJ6DGYfal16y+5hTz0GU9zxWyPX
L7jZAi22herBHSbdip5HWHWesWfErq+qBBWxuhSR/pZ9iCKaGiD7sZ4y/RKpa6td
2kbc7R58tLpcfGy4bGboK29yZXkf556Z3tP7uW1hG/+HtiUDa9JFGGOKD9qwcm/W
o/jCrS94CUIL13Ilbs/GMDjXdOGxa2a9VrvnvxrZe/YXH/dBk7GF4/OqvY1SUByc
uJSrENI2FvdS5YXZUdutAR/NtJU1u6IPftEeYh1wNLICIT2htyaKoDI0bGmX064I
VSB+5sEqgoAVkUV75FAufjTWBKqlhDN326yOGnb2ISuiln7lvFGR/KvJSW1doR4S
8kRSFyOjUNEl5HcUNGARFOx+gUN5yKnegxMOHLUdOm5V6CdYTeVrrHw9uYawxkDL
RLrtc8mprvFYHk9wkaRe7ZSk/ckW6GqUNN/8dYyO9EnquDlTms1ZOefLu0LlXcU+
1/9kASoYEzff6QnOxZgxm4/60NNZt4wNl4qXNLZTuzZDmxzcSNiij4cimFvYarey
jgkRtv7CyNBnrIaZGaqPXmexlzOmIlM1eHiTI/S1MeuNThjczuyxO0x+0T3jqoXp
lXOtErc8SYzuBTvgqefrKXswRCeD3AlZad3x7m7QUbcJn1RAY+035vhpqVMHs1gD
+g+XparxiNKizV268RsroFd54po79a3AhNvMarGRx3jwkZyJe5EcM5Bs2YkgkT5l
0Z31F021rsumZNrrnfaDJIavOzFTrRsc+nGmNo69M+teWIpIw/QcLV+qUlBBBcw7
KhHhNTH2/jtfcqBt9ouaPUFBGYjU7feCC3E9DUSINSH48dj8ythPaQVw6mjsU3xd
FdhtgOUgEpQdYu6/KE5ACp9w9pLmRu3PWZJ/I8MP+m5HqeBWbPjnaHC/GnFBxOCj
x2Kvx6RXfHsgzkyB60aF20h+FxqjCITH2Pol3r4VcTU9V5u9XWubivTW/bth5yLj
1cz7yuQ2bWhvykU2EYKDzbJGzSmxliSffWqtubsern1W6Z9bCpiBOiF7DDmbklU8
e1jk4cAqs6E9/WsbsVDm0G8Z4RkECPFjw50I3Y0yMVskTDB9CPUvSM29KzuPxdLd
V+36tc37qnc0snyyv1YPjzrGT1tP1SwtTWfFCjvZbfzqlKSRBSme8bfH9ol0ErUl
SLOZGGbwJs2WZz/YYde5HDdPY5Pcyp2CSxW7fWausA4UWNxMRc83RRwpiRXUioeq
r4bztUKB92hEZ8P5hwtrra5gKaHhX3FrjpvIVZ6jMJ98yK5PlMlio0XRFLyfvTry
AgAWJRUXyo2DCV7ibTno65XTPz3JnZIGipWmXY7hYH/MaLZod9uBrtAbS7L2RV0L
cflAJnCN3odZz49w5KSM2j7JQD7/WBBvAQXMMbXF3tRgHhd8vtmPR/gmwH/97KlS
8fIqeHm3Xy2RCjVIc5Ya6fYCTulnrbBjxYH5TT8z94SsDIVCTmHujMi5NlhA426N
1tjBKNqzSF2pS8CltdD9nzj54Z9r0mr9MkLfhSNng3uNhvu+eyfnsJDMLbayT6mn
zHK/BOvhpWXO0yhLIP/DbISl/3Uf/py3RxddjTeFqjEdkr1HiFpS/pHF8tubtBaq
Jh1KQst2cHZk6OBPxzfGY8suiYJFqytneI1mIeqmKvqWgaChLvCuajjO6O7LVKmJ
OragaWW6IeQzhYpyuQ1RMLi8EUh5LBe9XZrDJRWjs3rmVLOvVui+SNVdMvLp+dw1
Q/WReerNeAmyGpGzupGRwkJme6yh8sTG5ltkLmHmGA1Ic88Zhs2TMdnPuAT6sqP1
w9DbpyUiiwmVWxrPEDjtDG5985G9DAYaFt0F/Ncp3bOuo0pODlcQ1btJ2XC6Moar
gI+57wxmTgcsSMeHj02jdgNlcXL1CRBnP70LEfUE91PHVqkzfuxkV6NtiKAoHcD/
N4UT/ijmxYTOWHD+4nBQyJkNQLS/OuHJPdG3uo0KLZC1gHYU1+5VQK7kh+I51Fzr
aJaDmNOvfl7yOmMAnbdlHVrgVMQ/14h8I9nvtgbBPRvs2QwUuhyvGVNS0lxppgM8
4C+EJIbMO4MgmZeLDWf6PlR0OZB25IivgQXNOIBrkAvakBQ6bTMTy+FyKwMgGpaC
BglYHh7gF27WSHGl4f4xy8R8pFKI2qZWc28AYTBx9UvenIjtU8xQV26L7O6OnTVQ
oh5A4X+g+BM1SSlyA4As1ZJ/4NpZafIOOvqwLBNz3nlkxcbSXfrjyhzytmnKTRUS
t4Z3DD7zjwxlWl+Tq6AdWTBDIaGBAGCWkGQ6sEpSCbG4th//IOw6bf7CdqfhBwSi
MpHVtYc76BhMUPcKIV+z8c/p8o40G0W20TwN+FcWftF+VWmVxIvI6beemSWbbrji
8vx+eQ/RI1hgv9luIdGBEVFxkQlJEK9h+76ilCEvKHBW5x3X6sv0l1y3WC7Ed06i
sTgk3MMPiEMoAGkRfMp0SZraDrefckNuyFrr0TTzlYu3rBMjO691hrJUrB0r6SvN
ayL+KP7IlyxSob6w/fRX1pJzivgtsLGnST+a8Sp3JwLukqrgqA/KfuNuDQaSno2b
dBgh74km0bAaXO0cFJxx8snIN98jJq2lSExgZB2Jt0zupRhZjhYCWX0zD0YX/1U0
CMKVsmrg8oi35a9JoNuCzSQBHyzU5U18Z9HjnsLIYu4ZHE1B2AGg+uPKkMPL5bQH
8icTYZkMvqHqZ9tLeC8bbfyxxm8t19TaJNTXckIo+WgxDpLOu32Up+mtFuyLmnfs
c5OYrcvcd/NkFJCnVTSHjwb1z1lQClVczmKy3S9qe3M1/DVG3VrlvFrdINAryN3Z
rLxfQUtOePEzIt0TqMQvfgpO3piWYMLr/Tp2UyiGUUdGVsUQZhU0fU8vXVSaPUGH
ZuzkwX7Wfcg3vgJUAzgRrh+6i+MXSjZJZMIvu5xHmNu8ntxchp4CodOCCZSDjGNX
RxKwh5A+aPX566ujP/o4nM+yvU05pSJjV/f/6JIjuLW3BhqcjH20W7bADdEAKGQm
z+E2/njk7I39c8bKOlMUOzpTTrOsAfQ3vvVjGdk0mohV4OJZt9r+A1nmZHVZea+t
fUxLtnuqLo7CBNxmwL0iC2DPB3AkX18fVrOySE18vhRfMmYQbWLCSaBIESSniwn9
Q5unK5e9WpKXBlSQVl5NPTcffbPHmVriKL8oGQt7+7Mgq8Kxy268BItKjbsJOoMO
mW38eZJ1us0aiGakAb6teBGVyI7zI6DTsXQrPTfcKwxUoBBQ3CxVkroGeH5280Ny
klB8McSgbzyUjTz/gox6Ldw7aGNkDu8gYEJGSX03Mq8GTCXVWCgd6OOmUpyMIhch
Axx+la1Iz1D8Qv2IZZ2JLl0S4/sPqfzpfKQFhgDBIrHPbIm14/+QfmPX+KRDpKa5
L/EW5fWvaFzYzM2Kb/HqE2zw6zNwzxlKakcEGNR7Jd4uwuaXzqtQE0ksnNKQubNR
k7d1S5Pe/YPoNBWRWynB7gjSwjcUVoTzX1yfXEbgUSEFYBN+aumU4FtQjvL7QMpz
DTDvG5iNKYvgltcfG7p9Z5jugCTuOof9Byb4WjVwyyIqSKaEHXLxg6k/PqMUTXPR
EMYl+Ti3u/IngtMTr2yppPAVnyQB3oTMABIKvaYhhlXPGJ1Ase1YPGVO/xGCUr29
e5YWo4yL0YYAlb7F4TmvCr7dB5pDM+krH2B/De3NHOxrxqMWAikj2D4zyePha/Aj
cs6I/0rBlErVebZFR/PB7UxJ+J0bJ5ipAR/jKGEv6w2BJWnRiSogV5ioIWm7BF1K
AHA9+WlyApV/OxRxg0yZgUsbyYOpm0ajmqTpyoVEfy4HqPjkKHxDTKFIDs1ejTrg
pl1me0lRG/l9c6vo4xgjyFd8abQt9KvRtJ2qiJxWF2m0+zIrVedfr98Jz2icTHnx
y04hdj5qy+VvXw33hkPKcWeWsYOlg4wJL6dhL8YNvShywvnXp4g1zHXAreFk3M5f
lWpBX1b3muitymkjnTQA6Z+vnUrxaDSQ/4op90L+QXDhdG/VLwKJmpnGaJlnWmmK
uRKhXBlFqzTKTVat4kJCcLakzTutMXCQ/j20DjEJ1FocKHw1SYEjURK6aOFtDMlY
PWL/Gq4YL4UqR1dVSffwFGa1rnlQGY98jrvVQ48ztIkmbnX/3XVjfJ0TRSfN602l
kkhNsC5fc0x99kPEAgouS/CBSLkLJmZxFIFqT5QqhFdelBIn5dKYWwffgB3W6m7i
L4XL3V62MeQAnn+kLWV7WcU5s/++rdc6ApUQlE/erar9HC1NzdL9Slyj3enJwiGD
odc3LvwEUo4pKeiuDTVxy/BiXvma6hSVOiFGboMBBCxvtjcDTghqpFH0Xcn5fa/K
DWig5tOHUaZNE43vK3rQrjFppwBwgQvkQivde15tZu71YWznZFGPQC1Etp4Fr6j0
JzPW2cm7YlGPGuJXRpMDasuIGYRVhNZMqTqWHwANjvVCDpResS/GQQ5NDUYR2fQX
3KtZRfDyGvGfNhlfOlVUHYDaSKLhnslUfImoXx+1Mg5wISK1vFmlwaDU2KbpK+QZ
uiXW+rKGyIyx+PMP+ZfA6WOqMlcEQJAKwUZtw89cQC9O3sVyUC7wFl4biFZ3whJz
qdwLSKEkVVWucDZea5MmxKnZ5yWu7MVCOylxLFjttj89wUVn/uSIKHNPDMMn5c4E
z0SeV2JShvuXvz1uZH33wiuzBClLt6bzK5WOOunINohQl4xNcgOZXzOrDSDkSliJ
4qFDYo8c1ciAmK+KP9+bts1nwVIFoVP+zyyNwg0PxB8ptTD2qLstkQKToHVgvdKV
OXYINC9T0dUnmIxwsRVxWSKAJAH1tobUN1SHEShnwS/4Dey/BMk+k1Y5P3CMfiqv
vZbVNwHXOYAlCfgPgh93LkeKm0HWKFMdWjpAoBze4BXitXP43o9ZwJ7wFy4WX3xb
eYsPobHidtae9Pd8ipYzA+41sHi6k6oi9yWnXwME6k7Zf5pMX8ntA4gl9BFtpe5Y
rt9tf51nr9H3bmyrlXhbINh0dWWkDSLx9Hhvh96LCjYqAx1IO0iRZOVAVTrCQEqO
/kO7k5SHc46++u1OLjZgyfbZWUQz0bl1nB0rO339v23NwSjire5gIiDLGTy3BT3y
zSad/1a8A6WxtsLguT+MHCnvbJvJZU7oFuul263WXUScicSE61XgBKcmKoB8FJLm
rY8wvYn4+FUd7hOxeEkOvPvzpF4qR8RmVn0rnseQ9HZ0MFugCre+aXgqf21g6OwV
XKqSLkOTLXEMr9sIZRTnwoUoUGvpZffHQRe7N7ZvqCoZKYF2M+wWPZGdnPjCbds9
t7lkjo0FegPN+nSYqrLyAWQZwgCYbvpIjP9bMwL1y+RcHf8XPP54Qiudolp2cdaG
KtlZvFSkEYdxp5prwZ0V8FEV3L+FHNhflqvfTwF52GNJvQ1rF/uydG2WHvMskqdq
zZQ9EI8NlRW4YkymPWpHYFMFV68cru5ejWLEzAp0qFrQ/MrIK3TvHiWDZddOis7t
ZUbRdUjpVeyMolj6cqq4I519YvVhPG1N1FIgA3hviBNZQ2avbyXA8pgfVQrnCq2L
q+ULaYWhmgbm0fEBZqFrMOO0Dql1Jzy4Sa0BqvWC5Lu5bM+1emmxzJj1xUp98O2d
zre04yL/UY/yEwhuuGFRKFMLrB2iXnFcj3cxdYNd8oZH4y7BtbC/8tFHWxZzGB32
BU+emnon/AGJAVG3NyD03HzkR48xDA1aFR46HRURyJmGfXJ24XIesFIJAHs1Tq4V
FOOJhD2lqaiPD2GOOPjLIIkvvlRVzFaJe91GpchoqxcGn+btBHBPKs+1GPs2wKn7
GdUlYKn2LBfto7wYUq8NNrKh85dLKn0KgbV9zuHBbC1XcmGQ2f91fqOOlRIwIQO+
RvMU4VpTrT8BE2455cwmUqWcf0wTS5wetZl82Mfkg8UghFfwSaQI9pXdVafj1L23
U9aLkiqRPu+O/GFzXQQug2ddKS1789tecEsaAL4EFDs6Hte0Vt1Aae57AWtVp1+8
R22cTJuZAXT3t04H3LY44VFpY2KYFbSRMbqcOcvnObxOPZ7U3Z4oGUdFxGZBHqy1
LR3VnvWwYUUQ67G5WoR30BrQQ6cjrO/joYXOG4omlFD+1GcmUQrR9wWE/HO2GZsC
RGNd8zOB+AGeIZ7KRua1RIed/Rl1eHzlNEtj0sVKWNKS0aSlUf9ON29JreF8iO/Y
FyYfkVMmpzDI1V38zheJVdAM3j6PWb+TPQf8TrP/y73/Apw//1L6XoEERdtGu0FN
lFpcoYYmmBeZbb6JzF0fIPb+2XqFHvBx1fUIe7vG/uUmHPHUw13zAKoKGM3Mhz31
BdTZ0d5k3ZT4xtjxdwe34dcNec4j5ktS1UBNaepJWmTv+C6tqEWgjoogYdCgcORQ
Fagxt1qSWwrb7DtUzQHNOpBgXW/x3b99l6xQzr1hkehhiPMBMhAmXPhUqsb8ZfeB
h7zSNUrP/M7YyjE6kpiMBwKjyhjvDa0K0+DPKT3Tr5ztdCmI7ce4j5ibe0V0ho8k
9ug13pBi09iKpo6eNjp2WuupI/24A/g9dGCkRigwOLyxHGIpcxbApdaCm2VRL+vP
V8l5G0FFom/NkpG9Yxb2FF/zJdaIv4b0vxEaFPJJtj5f4+U4sq21s3D0s+mp+VLw
Hokfu2OFB7jDIeKoLcrHClI/iBI8cZjSn2GSTpX9M/E2DtPI4uUYDREnbZFuX4ly
dyWc9mvZBDVxP+l8aXzgChLNY/tanOzUqcSIgtXm+jbzSkNoqHv6cic8R54Pq3cX
FxRNOftQqvcCSZlkCLHOde5Ci57jXOyF+pnQrWNVV6gDFdDmer1GtKEQDTztEzpN
fG4fvCFQD3tyNvOPZ1cr4EKvNNIzuqO14426IgjceRYcCP2mOQD/xXWXAuDqN+LZ
EafqkPfYm2XcFCrIDB73r5epf9+EyytxsLT1NGW6uFE7F+wO8IHTv7MlSiq2G1wr
WYvUbgojHCRqKS0GKhSWwd+4WNbF/ri9KqnYkOTzN7wwRndyDAS9Mj58wnXOzDgq
eb4yLmKZFq0UdtWXtJms5+Snpm8wDhGGtPZMkw//rKne7XvNf0ObxRqO93gkkUFH
srmVigrMhtYpEkAY19m5+fHsY/2e5fQAZk09NVwyw03yH2zXUKxIGn0vyyrAriQX
pf6nwpP9KPwhromikm2xnBij3rGH7FC9OLSfcbbSzYfER9tzJ6vJZjzcRKKCIAyA
B03qp40uW9QfUObjHs+EkZGB0tUiRQggfRAsx3qmG/tu+gICn9ShUBCrENNhp3Fu
Vwwy5BGrCBTcg7d/gZpAuUrLqehhtv8kbYD4v/1aNlFivVTXLe5vqXs1O5VwQR7p
w+u6OFphtsG0FlBG+szMIw3T9a7qupb9FTjRZdAViuEtnYBxowv/Y0tA2UZyIMEE
wBMb5OCSDfH2AsrEaWo/ksVa+2oy2xHI7XBTZL+2AIPjtpUCqV6S/f86kTaBGqox
pNgbYOqNIyHYb6Kuu7r1ugBKeBL1o7zOFmeNLs37EEYQ0L/E4xPbANQgd3MWKh/L
HDum+tsaoyxGPM0Z7E5PjvqasqkOSEJvo/FDrepkUJSFgmK9jfzU6Z677LakgX6E
IaainatDn701QGnNrR+rcqbWqTKADoPvx3tdFaViu/zqqDmEvDYtGFYyErxM18Y1
ggezUv/nam4kFqatG1z9F9kt+OUWUBk7B2PB613Ykky0Ca20JATbLJX+gaOYnUd1
+ZIIbrH1o04+xRLzzY+QfmTMf+t3SHR5WbpZGAd1Ws+eAj6NK0JZC0SbDY6Cwk1t
JjpAf4zw43U1tI9ERDLpStv8PlDRydtsPyiksJtFzEvqu0mFOtGhw1otq5Q8yMs2
jF9/TmCXAMlWiZnmeK/ON8OgW9y2SrDndV2ajZCevKuqSlt9Nu6aBZpgDJufAnN/
ficbsqo6LlpYt8hDrVROkFrHzmoy6I06vMkNvIGJdBC0nh1x2OrZPFFP31DOmBh3
OAMeYXtePmX1m1ZzVi0mAzXWrZVL2NP2U32uOjAElJHxTEfHqirwXH0HR3kqVzf3
tBFvXoBszGUPmtrKuwBwpVXx2leb02hNDtaqWBwKIno4A2MxnSmdxS1nqCQ2mIsZ
dXY8CrjHqBTdyXpL1h88ycUrN/dSMg0dhgQVIUfT6iY2gQZywr7AGU+sbYx7lcJj
CZRVrKvqcShFjjj3TOtcuS8CQeDMXoZUhw5IK9Z3YuXoK+GOX4o6MMWo10SyvjBH
zyVg3KAALQItUgwwtb5wjyrEF435GvtkVXBMzSyc5TwRozK3Eq1rzZksmXm5FWQl
liDX2RTp1RzIdn08UhQJUjhdrulNIADmgdfmC2PnMjyzlqZc3NU5AIw1mpm9crxl
2d1NmjBvw1E5x8llrUOY9qtkXw4JYTCetpKyp1rjtZ6K5rYzNQpyb8C8fsbf4fCg
fveQmJMmq6DgGCJkfEcrTw4wwx9ZCl7imUAhABBHYYnc82rj8xuLluCb4nVdIWIl
6lc/eSZ5qVQNXFf5a+90eJTVWPtX/bO91h+RhWu+Ff9JaaMQBXu0qgjWEia0vHii
sMDXV3KaFDjGpBP6Rka8aopgBcfBG/dcyw2okFw9NbXshuTw0biq2FM5gQE1QQMd
ykC9hgf89YCA6+lhZZyThtlyHVwAAXKYMxAhvHjcm+BOlEKx0xhlZ/NuHHMYrykx
QxeMrVRkH/6Gr9mXeocHhJnnkltfC9/zubdTWVSWQRl3QIOFXvgisDZy74eJtLTf
5vpXZBgW/3v1Ml7ALZC5LkM9WtZ5Sqfru75EXKw4QCxom24HQYdE9aui6+U7JJ6L
7TYZZjRCDeDQMsBYBIsi+JaZv0YFYOMXhDoybdmliW6/hbmilFR67rNHvTHdQ6jK
MIWe+0IjulfZ17KCUFCO90Y4exhM3HrCM+WKbHFuq4X6mMX5oDluKFxja+dHj49z
FRximDWA+Tu+3xuE6eAPOKgQvsyCvFbbkuYCDR9NNwtZxPu/sF1S0wt2oY4ndHU7
vqlsexfqfnMymnv1v23J/NqwZv1qXCLhQMAMT+Z06l/35U5Cllvqv8V/fREpiXoV
cbEbPqzDaGHEXhVowAaIscGI8Ek1hJIHRTqYkvFVH6rsIgwbdPFbc5FppqSwbaLT
apY3Vq1ht+Dk6WCA6kN7R8SKaUbIjqKAdGFUahhG2qYxyVpMoG53aCKv/JA1f2sf
D3kEr7XAL/VwUW8U8bIBTaIqb4mAv05dSk6ATEpbSVea7bOsB6c/HNfXEotN2fi/
dqhZbiLYvgmN0LPBZvpMbS26dVbgz/1BVFBfAuFfK5VBaOvVhKdY0QNFLgiyL6qw
L1BIxfxzXVdnfvIlPA2RX4AuJexWGeaPiZgl7KpVTuQ3r8znDtZKj0iDGEowPsvV
6ZlozmzuBnCDT4UUAbCsSpwGdkJlqtmnXApuqsbLsteW55eZA2P0yaSdJQ4OAOQp
dCwKIS3G0iLFEKO+geV0h3/7SnUoacKJrdsNU4Fp6+vXw2R05vx4i2jerH1df1zl
uuwD3z63/TRdz9fBcFhi3viPbxIYgSB9ArKjne5M/q8leyuqYgD6qqRl3/Ki2Mu3
iNibbFEkEm3H4YGwth18WPXGQF7iZqAurb91/8Wrw/vOcxokItaT/1mA6EKZAm/Z
fhInTyieK3O3vFqJolM+2xeH9gGpxg7+bgULCbuNfXNNCLawjJnUKYsdvcf2Mo7h
B/I5l/TCfwM6mthXbEpfcuKuiyo6oRtjkb30Kll4/1MCyqcJcPn0t3jgntXdouAP
WQSRWgzFAAM1ezcxQ+Kp3mQWV5y3jDrvYZSq6HoEg3RFVIJy29n9BwpA42i+UKx0
xKCoSgdrWeaNU/S+GztVKOB0+slWd5yy43InfoBhXDPXSuRaY6nivn+qxOXVlkw+
VE1+GwsoJLD2YiLsP5eXhochlHZGqEwD4pL02kBvXZy9CdGyHA6LrqI8YwPlrcAl
pKzagbBl20pP0HSi5pIZxYyBzgXGj423bNmO/taQO84wYz4ES8Eece4X3Af3tZ7s
IKnzllKOa6ySUWCRopDUQFX2yLN+lEV9Wy1bX6xgQ7XTqTz5svhkt90AMoeqb0TN
fAjdQ3qmnoJrntd1VIAURW3zRijen7lERV7cUtSoM+JlDbcNO+uQEHZ7nZzWkMHO
3QO2GDplWy2I4/uzeYRwv8VjNlJHGCwUcBjal1fMD4dLAkOMP2LRj0nnB7mcG6EF
btyADiZ6ebRwSKcyfNDTt0jRtPpnyS2W9rpDd6ndGdjtOABjvS71SQmzK4ArKlCq
DrAbnMBe8JIPE9Yi8Tp1/i2JOWGyq2JtHtXC4D6UabAPjLwY52Yw2YaMlTyp1IiL
9gJyHmtp1gVH71ns/y1qjsF8HKAONFqfZbm3PaapIlCGffIFPwLux/Zxh0tc7vB/
HwnfVtNRTphKk77Guf3p8y4an7vTP+gVD3SoV6XeSzhu0AmCIhddKMzbrj/qfNs1
rc/4g3FjjHK2smVHv0r9Vafej0xspZZJgqjupHiC+VPuuR03K650XPb0FLMmMsEv
lnFAAakA2EWqYhteW7tt2W8DsqMxLtMWylZpe9HiFbvbp/vhZ5y/5cEYlwEp8DK/
S8JyhvdroCY9mHiftLl5Medu7RneEmNgYXdKUwBf5pSlEFv3Xdhv/RIdO7C72KAi
UNYlVCeMiT7Lf/80iJ8ywWxX1DqS57KCvCBc+dfBa2v3ojAwgnIRXzA7VlWDT1DR
Or/4x+jMDMqXqvGptlijXaA5gN5cv9qRglWr2npfo/iFKaayDRgBmyQfXM2rv5TD
FFsNkmQhbmeAJ73NYIbmgywjNgJE3UgqsPY2deJNHyCE3PT0EGdBb8KbyvrYWYtZ
gYXtE2V812gpswLtfbT0GbYdyGWzrK8Y/wmmCbdcsmEjRyVcEb74K58U74iyhKbd
ByOoNM0cmwsBpmaMJ46OpTPZ615ZA1jUHebqSrUhuVfdQ/zgLprzwc2vmpznNfGN
Wy23aKj4n2yYmdXQpCHmSqN2QL5SY/HV1cEqzccmCXOfuwppbKQhGkvaaN3sizE8
r8FZ5VRweoXuBTONrj+K8aVh/M8xHKiUsl39aTfRFt00TpwQpAOBTJuLIZ74u826
Mf/lWKLMNS1kh4bo0NroIjaGkWTBgFJ/1q2LdW+h2rmNrPHAbVqiFB76NAhkCUbw
Cx47RwU3YRDYRXDLPC37Wm6mOfs6rdG6pgzNRQ1EvifZiPCUzPaqgI3VKOtoB0ny
7rODg4UZXzZQr1yi9ZdoFtChvLcfJD23vgMZSjm1jvaFZm1FAhPB2dTHX7dsmy4W
BInkSfwWwIerXWHFyX02URVnO154GI9uMM1B/o6dAKsS/uYASxI0N6AfpjcNhTku
Ib152Egrn1R2ftJqTo6ECyl/8hlDsQhVmZyoqTSS2rUi/zH9Qmbdp/6G8Rap+w7R
CGmE6F12Za28fn/o4hFx/AoBhmGEEmYBS8qT9Vzqd/CSQ8syKZ4ziso1OV5fpQ8h
OyByLgeQkb3jpte1ObdeKomBU03Ow5sZesOzhNAHm9FsRfVuYsnDhO3piStO/NoK
SQjp+C+A4vA1l+vcWyqIwckXXDu/UUaN5nedCCKWUyEdUgzna61pcNb+FtE5I0Zp
YXbJlew1A5ULpNBSMd1Zet1K8qtYnQshAnBA8L3mtC1BOKLvdmpx0q4HjbF+1pXR
oIbr3FIG3DD9Mx46YCW680nStB84syQEAqyx834CdSImYdNTQV8xmRPr1Gs6w7rt
0M6d9IkSsYsZtpOUP9F9JFMV7MEoo1mBGGgqjGIl3yAvu8otvhrnRznnnftz5a+s
WVCcfF4CdljA9qZwTBWF6AXZO53ZBpHRBhV9H5jMCDCFyPMjofKyclwgLA43/QML
Sl7IyxkBQTzohQ9XRgbyy8Hl0q5bTpxZvMQSVnPgm+YXQlGUc6R1OcH/aJXXq5r3
V/4kjYOb93v9p7UUL/M/LRD8uPM0xGSMteRFqVWljlxH6GhhYC1VbrLUYLXwwVc6
tG/tMCzcYDOEDaovknfHP8qH04qL/iBeKg4lgOJGWFgh0V9pdAm2xwQjsDUQ74N2
JygiEGVSNR8O1ejVxHp9Lujtx8852G70s5o3WCljNJOotLOAJsgm7+XGInHWQffP
RQUxaKqgM1+9DEGY1iggjaU1miwkh00AUHe9OX7JMD+t2zggs+glZE1t+feVmqbd
lJ2dJgJHEJT2NDQOambEK7tXDGU/dvcPIy2rEIJb62rLAm7Q4+owgODtDZqaAUwV
wRenwYSzanrbkUkrEot4OG2QwDvvHmcv8T3OEUN5E9gLKgCoSTL7lm5OSeUMatZT
v9uc5E84ouwqPbMHlRrgPIx+rztRNCOHsUsD3WaRorT3n6lLbuRzLWTfIUzSV9UF
mwapJH+62Ta8QihqqM7HMLkmx52/FRwyhTu9ch96i5aXskSsGFGTVOxEt0xuKcBG
7SlX1PMIcolh6qiwvMP9Apg8+Zex+SaxW+D5Fcd6K7ZoxQPmYZ2twLSUxok6Wy6Q
9kq4xe5e9K+syedlONrErFooUWsTXx3ir/qBrL2Lwh1gL9TcQh2pL87bPbWtAZAu
V+PXoCEL9visV1kptMqUKVocUEbUo2iDz9jtNHWKCWDKW0Wy4HSCG/O0P/o06eoi
78CPL6pX6VC2vJd1tAb9M4IwqCGuLIdpEdwmCiCbLcOetJ53dSgOJYze/1x5hXGL
LLFWs4rVVL+CGLZa6W3S1shuFAsacmSdona3HsG22VoaDVp6D92Dp3LIv1SGMtA+
JrEg7jfiqBtFC7D4gknB/+dKJh9k5lQcEV69stVZZDLoMScvoMsPpLXkNr79M4Ny
v8FcfgBCaqvc1qzNCMgIKFJ9ruYVqkWQQFf1eDLXp5UxaTZA4FmXLGwoU3hbfDXV
iVVWGTNrBQSl3fZIAx2JnbfJyqXxPjUaPwWiA65QL783SU+fOPBqgH+bro9oATiD
kASKaLgF/o0Lkt0y3N+tafsS7+NcdLe6uLLGhA8rMR4NRT4XNzhe317U17z78xL2
jaYs5xSu/48kVFH7rU66waSiY7z/hDC1o1289jdEZSDF5vfobq+7QZwdSJJRcOt6
37+ofogPIgOS9alirjbviuyW7y9/ElEERuAAs6+meSprwshvEAxWyQxYDEAdqKrG
71L8jzvYBEssvPshsdCtrPs91FtjQsWeMdTK4foKou4YR9e/ECDI7IZ2hhe8mfJr
WKhjzJPu75eJLFqlGkIeKQTj8J3v8UTEjuDI57SPWbotSjhRL/WWIg4ajKjZwhIt
cUST9EhWIxtjXW8Wo04y/k6rlUpCvp7WrUWupgMAhbg/vcJ+aJUJcSo0dNLsaWJu
LXnGfU15qh9qUNXOt9c5eWQBkptECunZTnh1k+eDYu456iHRgafEJmd8mro4aiRD
q8df1k4944yTCBEko6faecrtvOu3d9a46X68pPt5+v976d7ZdJAnPf3M/oCxkJ4A
pZjMMCZwcY/E0Ae5aDQKAgvLHUCugCwo8CAsfE8zgkzidofTliO+TNHJuA3kT/Yo
tsni1+RPd6kzOygfJEWxxUUEuLEjedeqKJzNHYHB1pIK/Wi4FIs7kVIjjM5ZaY6E
fN+uqZUPXJ7JAUr70mg6WtcxRyfy99EnwC969rD/fbxcNbvoR4OTvir5Gdn8aZp2
zGcZdHHSUllzCKMqUksdz3a9mCbZ9rJ/lkS5s2O2elz4DrexqvRyoApPUH6YE3FW
3HhheCbehAUeMI5g+xHLnnVISLRqpn9dDa8gVPcXp81BrvlOFCaunOQAT+k1m/SY
A9vv1wnBHm9X09FC/3DWFdQT/6I0R8SJD2JX3fY9rkBS6kQffKiwNj0FUQ0E8i9f
begmZ365jVSTJe9DuCrR+UYGgPWItIQx+Bt+HqVFR0eHu/TQX2bPizozxmN7Mpnx
pn3oeiZDIxsEm5WwbzKnU/c2XRchaL3Kok1al5o7aSKixmPZo+jWvThNPvc1jEeK
JEUWimZ2cfbzo2eEt/Wy/ybxl+iU1NbEUTjOI8IMDYllJi00SBVl+plLK6udIwY/
R2zAY4d47kwhsZ0RMh5g31cBXQEzKirYoXfGjbcwkBncdyqXmAazdJLDmIvUdUUz
nyyd8m9H4kZp2qJKHPmyw2BxYGTqOYBoxz4p1rU+m7JH6MC25r4zkRdG3rxpdZWf
/vme/YRwwvQG3fbXHgicXvtzmR9egwAd2SDIIVsItqlqYxO7PHBpa/ZDeeXCnbBD
JXPDxZmnUF9QcoWUw0J7uyZqgVFaeWNccEIhaKuCRiPc0XG1shWmI7F+dhhtB6JE
4MvXjPzrKMXLAAebRv/dT8rRZclcq35ebjdqm4oy3bkbDvVMk+li7fAskiMPAfSU
TUSO9Y/vGHmxjyDnSYqCxGkxCq5hrWHmWkeXTb4VYjpQcoZbUXhKgizT52NCGT40
2boSBCFPAUuRbwK7ZuEND9xTiwxcc00OUC5Lcu8kZUT/hue3y50brqDjZUuFq5bw
dBibgKR/X8wb4/Gz5sKMjl02k7m1OdO4c0WuDXcKa2VFXuA6/09ZbkaMRhyI9TRl
8h8L7Dc0YDzQwi6DXGAyyhxpHfzuIW2SVSempi8P2i75Hf8hdMBag4Rg7kMoJnBS
KhH6Wnwc72NS9r0Q9ROcDUT41zILJoK45AfsASuBLDQHycCSi41F2Rw/GyurE1ef
Y+QJk/wUuA1PTUnYOhJYL9o/x8YGNn8msK1q60ip4k4MyWS8T7pTwWhhwuchB8Dd
k6iTe70GGPeTfN8qvQYke/n7LDnFPbyLFvgT853Na8Yf+lXlbLpTUEexYd/FxaC5
/YaTzx2U5/WHGnsYEY90Z8bQZEtcAoF40gsOBBnppJCj+UOBEwgK+mR5ATFrd8nl
Hs0Gdy27NSDIxpj0hRLCoE6ZozsrNFhMzIc84DYg5uPgS/QwAP5PWCLmnC+E72om
WcraJl0w7NRyzIe87xFv9CGgxkjz4OsxmNTNGmFuHu6aGmom5m9SQ0p5XgV4Fl30
J7XX8oeywcr4iZ5W3RnsCXBWgTQ93msfMBBbol+4HZvKVtCe66JfssyNNcth0FOI
z70IRvmfR1OkIveBjU6LeHjvxP1EDWVQ9E+rrXiLv8jvONZKhPV4IWeTuiCcdDcC
GiC8KWLzPVGGKpuaovF469EOH5z8AcDy2LIAMzBPl9t15jtZqUgGUJnh205yaOIG
OpiuCj0Xt8i1NsVDKgCa5MoXCO6K0CcKvrFTbRkaoBKGbAWODatxUvtDKP4l2x4r
VcLvIfH9i9kHpNDq8IbjmkW7H4Tz2SPS6+G1DYzsYXBFlljhwz+JTqhNEEBhVo+c
HXS+RQDN3U3QnW11V3PX1s4zr84LShB7vITlChb5tj3UuQ+AleZnnugOqnIYPYof
Cvit3bfeAFkiQz1fVLXd50d9NplwMmqLOQtoYaY+vDSs3BSkHneRohxJFPPE2ZaM
r+qLLCZ0+DQM0kDIIcoAXCMQnonnr2m99HQQ+mlrQ3N/iFk6zq1e35VDTo+LOMEe
IxDAOGrVvW/FOGAi/NKU9SSFfuSt4ZNTLDi/4kyLOdj9uaaDh0riW66f1+/UXBKl
l47wNTfsSOtY5pCa35NEtGecRBfWLNn+K33un1w9FiXRX/xAzqKWhORw6IO+KoO1
94e/+Twr1ANrteHuzNKCsVmyN50JCl3Xu+fiVpdLKBCg8HBj6cDg5eLhtCYoaeOD
QSPHoKvr9fVoQoCw2QaaSYb2yzpZXH1GxYvNHhl3ThvclyNOd9nz0ahKVQvhrdLn
/TrHcekO25XEHka6bFbrDzV3BTDtGMyLzo9fkqQTwOzBrTk7ChJbQ4xarU0jMQwB
himA5eblVQvSOFbs+ntnkMmeHI9AXu5o8g6wTXQ6JLumRXSZ1k8KSEWfSGXcVsM9
BHKT7kIy1iuAPxQCWjhK7A0bUXrBJTtJ3bONwAyF2Z0sIKy1Tynrkbz5npe5xNZA
Q12TgKVac2rmvEezPYcN740CURPLScO96QJpY1H6cVY8M1ZoqTEDzog3LmNH/wqr
sHK5+TrPFDLYmOnGg325Fxe0IFbXQRpabHcQ6miLA9JnqmFzwEuOBGZnFKRxq4Uz
PnF8m8e6XXp+LFLu7cNSm8dAauywtODKYkT/EgvXdvR5I/VhN8/mvCLYO/6/9jIb
79WfH/cdjklIpmkNaI2RRggZ698fDMXlRw/0wsSyrABwqEy9XFCL7tsZyHadIkV+
W8oTfEEaJOsVi6Jk9IFGXTw6576lUj0N/yrWIZOqTSzUXrU8+MHFFLbK6WA58pZT
hav/hIQLcXEbg8sP3oUAggIXD+XWGBHFXkDO2v7JFKqm0ddtf0e5uMjUjdpg2MfI
F9qYlnR19JDNXuVDNkih/EYvU2/o++9XIQBm36R8vqwNxVV5tvkaA1UkL3Wpr/F+
glEIdn2SMuGa3N4VpcarJTppyw4QlNmtb4irlyAioEKie0ADQhq9nnsLcnkkPbVE
2Nz71qxZUo5IhSRrBBxqLlExyh/cmIj7XACln7AM3pkWU1qJ1AX8OPL2qRPe1ugJ
d4GxFIDwgfZ4wjOWn7TlKkqMe5K1Vb/Mavdmnl7dmk/8NXg8heay7H6L1jUFAeWT
Gq1gSXNxJnKqMsHsyHcZJTbvnO7b8Mrq6Qxcuk9/sPhb9GMjoAPcl68sIr47zFHS
xyZPTduhCDfEek1xb6MSbsrhQK15Ik8bXib13ot+QrYCR0S652n+sMt0sExfRI3K
pUAA4abZNmiK7p5xshAhvonPkdgQCY7xx13IjIH3GCnEol4SEVZOztG8D7VLBUTt
Dl4vbGCXTHcTWpVHtGVKalNFXh0WgQNQFNfR1gC3nc6xmzSzLCDe8xLGJ/olcA47
IBcA1wAeXMnvHSZ0eipUjeGrGA6mrAtppbc9HoCx4lH+IeldrgBAazJxBUu1DQ6E
BOnHaimLg1oPCavBFPBfTz0eI4BpiICXAoERcCRikOUUTl1FJOCfqvhnY3KtSxcF
1iwEB2YWIqYNmTuZDLCEYAg5mbbUsyJtlSrCHyuXpA4ag1t1RTZcw7c13/HDXaSG
OUf7i9FOtOD9De6KxHp/aNMVsDp3MLOkx/bH3+L2Ky5sF3WEyqGlfykF2mc2WFCj
q7n+iAQ0xxFiL7AChuw/aEIu68L9nbxQ7bQ1J3ajHBnrtqTY9NpkM+eOblDK3FUg
ANkyYnooX2L0+pnn48eDjeK+r9qpELmWhbzZOsB/OyJaY8cRwvdzQubAx6H1M79T
yRMW25d1pii8NzSHEYJRGz/dJF2dhGvipcfAKo4XHbfhF7oCndfNZTQVV03xqCl2
g7zvj7WwA/wL+tK994cLfseF4dMVRCL3JjRVlj1j6ZNznv9d7i9aBj7+tibymU/r
dn9B+CVJuOwWpxE4p6+CftrBONUloVKAmdCwaleYPOY2hmYJ4nTZ55aSbGfu5rWg
9/jswn29QYIRuDZgm+k5B97ZL2K8DakuKsP2Yz97zY0dM3sUK+j3kqM6UfCgOJ55
NIk1WLiQ9f5pn1wDnWS6hSJPvMZQ6yEWGlOK3SnoeYoTNJo7r/+PIAqyX2KB/kPz
6HOBqVSeDyfl87Fd+XVYYXycWOfuhfTa2s1QeBBdmHlLv9r6U7q3m3aLvO0dJ3QQ
iV3SE+LYoVBxBgEoLVSVgiXms7qzXh4BbCeVVlQMhxYvAL6k9cuZMq1371CNIPwa
vnejE6oV6UJItNqvUTSbWvKfK2zn+G58jEKcKK8jA0oRpB23+G2nLRYjmK/wugH3
7j1dg4T94IqGiVNP05BvNQKi1YecUh5kvmyNc/8DDRTrPNhWuVa7YvYS7MfhUt7j
GvDIoRYT0TSS1OQ9vrnasTXaF4wOBYXrDea4GIb3N6mnItHnhVUl2/Rcm5lxn+lV
BxFm5jEUslHGMWuKrhad6Hw3B0G/YR3JPDF8b8tm8PtrAHA7kU2aYBQ+BwtkYHLL
jqUnshcnu0tkVKK6c1y1y8G/VyzqV5HDI4wtgb2rZxXCIFRb3fpMhh9HQdymmVro
AkseooF2xNFsglxiWiiJ/bt8xKKEwQWDvAk3kTMtmn7w1FGlkJlHS4FC2/uYee6i
dkBAuZ+gTeCJ2Gc7cMNhAEme3whmioBPn2MPWmky3ZpUj01ljFpmQ4HA1Qt1SZmp
v9zlhtx3lBwEN2tpekVX7X1KofOqPNcohbCllK5SeK2yHsMXISAhoB6BjtZ2aIPB
MouialsVVt0CJcbVrRcxueR+ainWHEQWCgo64JuzaYNrYHMAfadGAVD/rvkx7xo5
x3IvECFsQffJ4w7vYtXxX93u22snXJpVCEUs1FtKjEZmrUnfOThYjSbRnPO5IAcQ
/hDUtx4ZXgXJ/zZqjx0fuXXxuupx8X06rGqCXVAzRGhuSmfUiwbPKCv67swVcBPH
d5+ntiCdNqmVVuopmrnBH7/YRZPcd6zxkKkqnwkwyY9Hrm0PG0OXdgMZLk0wuqH2
Ct9L2p9FJh2Y1eCrFdaWn/9OdRQhfkBK1zxCxDl3YgnEhkE6ZmxvWVbdiKc5/9Fq
VlZRhzS9d7w31TEk2+T9b8v/YJdwsSYdNZ6bTDULoFueqYTV+qAX7gOQRMEHUraw
MlGNfPblRNADaYFaURJJKDKvmSMcAepiuAmGWeQGwFCwIbmPMZxNAQPn7z+N5ICa
p/daBHuB8ohVw4a/X4BDOHgakZQqFnhQaZuXDuUcpC0uNzJ0cA0t3yDAq7Say8Sh
0RWVofhlMfru+5Rc5cf7zXlMMwuv79rf+UAmquI6L19yiij03lxL6Hj2bkH/FXNl
e45SPcBC3IaC4fGcPyWhxZd2lY57nSA8vsCEgSk5Ky/HxiBcNYkwR8Msp1EgfLxZ
F4GbTjxdNHYhiZ/WEctucHZgAx7mMxEOXWFywY507RahCQAFdn6BSBxDWKo4YJ6F
tp5cFAJb/F6zP+CK4fcpPhJmj+aqzSkUMZDz3N6TFVXCyaDW0GiXMk4F0I0fhFTA
krWNzqNt6at2xjDQsEkiS+e4KHLJv+efVS/dunbtij9kjLqkEXBnJSWsKMz1UnM8
BjOrhZmhYSlvgyPSDloxCs9bsqteAkkiqrsWjzLF7aOAXsYvt6ewMoHdZSselPtC
N4+qKO1BHpmD2GqEWUsHwo8loTUxf0fwJwKs+Q4/g2ravQMI9B+J1SGZH+gnq+Ej
t7tgtFjxW0MqGMnbituc/fT50KQCQZeAr+2fD5Tsz8u3iRhQmBMCY0VZKhffMrXn
pAHEo4EGIxM8yd6WedLyirk3GtHfRpQWr3Il47IivuLMA6InMri3FcNpn9XBQK76
JgyW7toPr7/vmrr0kFi7VvXSUKi+ISaoqMRsWUpieNLlw3PkSuAM3xXrd2mLNF7a
kl1Bl2h/b+TMTgP8MrrQzH9J0B6Em0Jgo4ywnlXT9TkRFW5SHL4EvTrI7szmaKm/
BpUeha+R6nN7RFdHsR9K+sONUlM/UCN42emTUF3seivet6I3g16cpfjBRYqEHxkb
fR64OkH99mEnylhZZGu1/90rMtOj40aikGyV0iqUaeMkFiSA0ENlo9N3I6aYcA1l
uIgq9cpDxS6J9C4I0IMy7PEXhu0Eh3htkvo2A3yo3DzEzc9Ay173m8WZNvNgvD2G
4Orar3n5e4wNxHUM2nys9kdxMOkFISkqfiLByZ2Q4ofKjLPQ2IDlyKKVeCNkubIs
IzIW29Rmyr89DMz24hJySZuv+AqhlPWGe2all31RgX39ajXP94GbbXhCcd/t3JHG
AtATgBRXORMfG91Bz05J876ce78wNz+9EkQKSbnuwTt10g2J4mU6AZYE7y28qAA1
FF+FDJRDFO+s5HlU/pcVrFgJaLVu+b5eFnD/trzG8DP1JGFZtjWX6nD+1sZZTLgq
dkHdxLJDhtb40DeC8oFIT8Y5euQDAq+6rmU2BehIhwuHTWHZqncxqDmVp8abhL8X
mA1c15ODJMeDodHXc6VxrHhO4r7Bwa75i2rh1egU4IV6Mmk09cdfxXSu8HhacrTG
C1mb72RyEGNTcY8vO2+BpgqR3a/Ksv3c02upf/JPPi2jr1IlCX/DOwEGxKugp/cM
ahbShIlk/NeD7YMQiC/8FHuQKxVL9d009BrEzKuDW+7fCisspeBKsTrU3q3RoUUC
0Od4Bz6MdFe71RiYiPR1e1hx3WTPOgIlwr/8vAF6H5ueUj3eyzFZXy9KovfSMsZj
dIJcFd+vMQqE3LQNb0759vlgXWXdYIOvb95QVwtllc87tycdzNnTKFBMwmICAHx2
hupeKG9YfhGmL8TDmKAV+L5i5pqj3vCUxkIIVntxkBrdvho41uS/JLIw3HET0g5/
pI6fCYKbR66fILiPvzSE3BRXIziWrDdQ/QhKjvsnZ5EGLQ6AM2WH/+mdbZhZm1Ts
wuP4T2F8crtJT4T+20lKMKyfZbFhNtl4xzWI3ZhqFHbL8g0Dsm5f9F/KwhGwGfQL
lNHJmxwCzd8ei8Dw8+cR8BZmDb4xk7Qb6Hy1JFLH3n2lXNQjREFBEs/GxUqxHuSh
iJ9EEVhRgxiycMLIDmw0J/BT2j4hBIonU3oEMnVWn2i+9n1a335jwR8XxEOuUgcl
d/j35eWGA9FBdvkvHnmZjeRgRqnIFtimZiY4hgSLjrdqU2nNML7SBBfdTgw4gIM/
eCF+Y1+zcDSqycn3t6ykJLR4s+T/iKIv+bMwlm1TWZCX0ERfrd5ob7Ai2AJMFiog
UDuz2Q0E8pAwh7G+uaKCxMfFBVcEaMhY9+PlaSpHpNEPUiCt4jam5v2Yuna5/NMY
RKnv7P7/fBgMETo83tPiRNwRFzeSMTkFhAVvuVwKBEsMBdcs38bTZw7p7OtTpUdM
0N/NnvlLQbSiH25CWRwjC4gPZBJgmYxNYRMx2DiqcAm1lYcWQr7DOt5qtAVoGi0y
8Wc3rZkwzHeGuVbrvDmEpjhHj4HWUp7nDfx3wYdI5Jc4jtntrv3o3JAWfOh5fekk
H3Qq2CWOtWTBV36aQLG8aiKy1FbECqUfdyZ7JdlRAQD+7K7Z2v2mHLGvKS9PWAl+
6t6kxqt+6ekBV38+muVGNwaWMsAvTcndneNbohTHfzFkLJWRTdXYVj3dYLiwrnNi
l/67qjdxxsLBC397MWGcoAXCASGMxgWhozXk2KsLqMP81et26EGvnX9mNBm4t4ja
i8DVfmvMYYlzHaWECDx1NHBg5Yeun4GCPhsaTXanGere/SckFMXAm/zzlLdugkOd
JbHhpibG/GXSECPq5JUh0vhGTXhNEnXpRseARdAA6j4cZ3KBrhSel6cFPJESm7y7
OFWSWZMA4xzSHCF962nKgE6WoZfJR903deo5LhAyO87PAWtFGlzXmMsHfs8D/MR4
zsYLV2w6B5x+nfGCUbB4SOAlCS9i02iFOKDqCDp2SiVIOFA3vSEZ7CWOyVz0fKgD
50VpsBl3Rv7efylGJfiswwRgN20mSevmZq1t/eTkISZ0h6Kc2sNXF1J6saqWv8r/
QMxZhYfEtXhl0bTmICV8SFbFfj7Q6WHlhj+xxDHA4lO6/epZHnvFgJpNuy5GUWK3
gLD1Sep17xsHysT4eI0Orlbfsb1tD9SJADp4672jVof+ZH1M5u9tXOs4aALramzS
WcjOcg6YOyoRdb6kc+sjt75g5zlv3JYpeqGQ7zZhm8N7WG9WhcfK4zKYsnXvJXv6
voakO++RVaJDgf00tOhYU1+H0oA55vx5GEawS1wXx+7cZ19wO1Ue65z4rSLMj1sS
X5OEjOWa1afdsUjhee3m5P267KM7nrlTQpvIxfQePwwtTbEaEXjykU4VnRDxsUOf
KMOgiAMPoUB2atP2xuqBf0fcz1H/9Vosqur+A2XsnPN7x/jf81LIUkgKDlmH3e85
YHlrqeaSOGOmup+HKeYIgq1GV6oSBxEdaYPeN3bqV9kuWKzZytrizXuhSu47ol4S
9yQI17hDJeUpdiwBsaHe8KoYx0seZR/NXCd8X+1bQcMqMiVB6lKhS7o0v/Rezbqj
RRq64QR3XcnLfAwHc4A2WO977GmcHQom564DGL3WGRgJ+5aVnBV2VkNkLFHZNr5N
wDqpsYs8NtnZQ6J/MoiG3zuLvcDRmqnDdQJfOC+XPneOYJNtk6wYqRqMYceBsQcy
D4kbG4GfzX7GItp8KhY3Q2zeWJmBnU3FZHqEnrtEag13+M8K+zBH9Qf1zMmLzxh7
M1ccTK0XSYfA1nqTc/aDHzxzM4ZC6oq7wxeNCp3n/c6TE+las54EZze2xwB1stT0
SfIlvOaPbwV8qkTud4MXgmEAntc3bfFg1Rik8II5P8i1x9zJPgjv9Oi3dZZ47Fim
EYmu94CdsYA+jYNMAF3oD4TVLsgi71lyuX+zzMiZZvUoEt8mwVFFSM+F5Y9/ipwn
AqGjnDEt0y8brYL+TBJXUo2ogxW+BbjgsDCllv3rXZI94odDbMupoB4qyK0dNw5y
iXXbyUroEoGx9SD2NAeN0/ZDWmqnfBgfXgCra/xWiI5JOCS+JaYWJd2wFKx3MzJe
RHZOlecPMwmOk0C2uDa8+UqYxFuKgsfs3mTKf7rmzfiC6IC2Whs55IEUk/wGS5L7
u3Efj17X7g8MdUcYTmnQQR+x3ups8QGA2osVh9sFipkmuc8VsrbG4ynQ66NXNBHb
+1QFwPn6Kre5xzvG8HbZmL4vADUaT8ZIpBbVvMPqS9lx3uZ1Hw21bOEaYzmu+2fx
JsJiyEq2yHJ/RJXC2gkPrOSQOW4cEdFHPK/MjjWZ5vfKGe4F7BgYzG926Yu9AMT/
LJGtsX2fKepHNq5r7skLHZHfuVQNrVA/Pcr383x52BrF2JZeGTOPCX1mfmPZo8tL
YUAFzK2SlI9MjZ33YlHXPQnColtmCfJqhzfg1Qr/F/sPk7XBltSCJPjHYLmX1hOw
ymuGSbgMdjC07kUAjyE8gcSzq+0efC4tmRBJAE85P2xsrLgeH744Uv+oA8upWzEI
0PbbTNY+W6eJcznN+/Z354DIt4y5SUFudaN1vYimwvwN/tjs6nPJJ4EW8RJ/R3Qc
wbo7nQYpvMQi6mdrBjj8bsKz0J0h38kPMJjDbrKntZsi6Mb5DsRkAGeZAHIIRkdM
z79OkLqps0qBq6X6IMczuAIVx6Vwcccd25H00IZSwESmzuaA8rTG/VnMTXPWJarw
je2JTsf4CqF6D8lJH9oZE2Kf2kqW2hwcNXVffT5fSof7kL699MMCKa+msazjQf4d
odQF1M4daCBsggw678zdQqlrbiDKpgbwc/t/FB3YM/K4bhnO9ysQy8HPj27Hca/E
QkS2TEzDt7DTQ+UsIVcPSXPQJ1jHALgTu3erF57s+pSEp6UJTN2leZywe8F09k/+
Zo3m0DscFgAe+/lReao0yOnRaCFHDKT0c/BdJ7Rl9EptSbC9f8twcyg0pFUlNmYp
QT5rR3rEM8l/51BND5e3e7LxB32kxprfgu4Qzk0rXYPuOxYL8DQceWUns2Itl1pG
+/5Ldz0NcxpfUzXbPa1v48W6DwmsgQ0ovchK0DNXRMwqu3FfKY4mTNFPmE8WVPNh
XaEL8o4zwMDmtGgsZ8wxNDYpxl3N93/JX4vxY2oGmaSwAaZ1KHo+xTSngiXeoop1
CZPHTX4DLc6QA3segfouI3tguSOBFh7U6i0938xCvKlwmUlzpkKclocdHd0+cBBi
C6PtFGHVv/q/MZedFBxmSXBcEWmJZCDFvR1uciGIwPV01gVFxj1P39lmIMy/zZ2P
MFMChJ/KJ2GmTLSkGDBve84e+ue3cXKnYz9H9qSpTtLeDZPhBXQaGyl1aoAoYwQP
ImZCMjsiQW4HjzUDbPfx4ZIRmWnTNibb6k0/02aNcsghqGmXUGeD3RQ8ls0SWzis
7LyjjEJ6lGaSoGsY0x8UCpi53xdNAzbZ4uqY795d+LQiRK7V7AjwKP50+EGk605P
PRgU1D8vBn5qHftNlH2L73seL9HNk9+sbO+BidtJ3l6yjRygcqUC/AyIR1wVgA4T
WTFIutMC4EDRkUuJeehjxiLO79Lo03uq/uEWT06eFmve9RLwqCXyck4E4TVI9lLv
vw6PDpC204RgYAYsYKP2yxspjNn+H2a34c8Yyz+n+01vS9oSbx9F0mAO8/Or4Kff
ev47pLkrZ8uSLV6YfkkQEdomOV/SyztYTLbOg1dP/uqtTybTjjyirx06uvKhGfWV
5idxlO2ccE+N0DHMVcf4T2fjlYslXrzRY3YAtRdw/oPJ+1zja2RJjiNzGUj2xfDM
h1XM//JBA1eQzgd/0GkVMS0gz1v6xx+FBQiEmXc7CSM0pTcB9S/aPh6S78Hbj2OA
xvyiVXq6fLYitnH5lHMDjsJ1lRcCp+jDmXYCX7HrlRRj6WUG0I4MC4IAd92JqvQL
zn1gHf5Wl4ayg075PnZOhITffmv5VYTxyAWxFVyJ1a+JmOT/qyCnzr+CjWurs0iF
1BP3YzHqh3SXrWXfz1sAc8ECDYnraqhR7E04tGcWjo90b2RPCL8FfGh3qCfnUOIH
Qkc0Cvxx0ySDMdKF2BzQ9Us1RpKQR9pGO7RIG8q3tRTiO6VCB4FzzaJPvfKFVp0Q
5TX5pAM9Db7+D45NemPN5m6RWqnxNCcRjOj2L6zKR9wEiOhIe5PU+M8h56nfEUV2
Lr3NlGh+Q5cd5cZgBVex67SLVVL2ZtME53Zks8kTOG4D4ELgk3uCKgDI2i+wTPoc
Cwr2lb5KvBPTbDO8gU/7Iiv9Mp1t9lg6+ncSEK2RSM7dprUS2IblCReUALhFnUOz
h14VhceIgKG+mswTr8KCOEhYF0q4aDSo1lNG1TCmom+YMZU3fSgeMLWgLzcB+DHc
YjbmsVBVjAShZvACYcZavgv8maMvzLpeFdD1/gLHTxw5Za54emL9H1WGXBiparEt
HCKCa/rtJ695pMKPD7NqdqDzTByYLYAk4eIzM0m76oaHGr80Q9IeyUgeTbxKG0bH
sW4Z9j2GATdM7VXbKcuTj1DfSe2yBE22eeGRPM442wR5OfBvE4bK67izuHz3QtFx
KgDJdcPcS+MP3t1VH8jA6lOA0s0NYe87T2kqOFasxPe8g1Vgkax3STRekkL0+hBm
RoxQ096hOnn/ylgfFU9XNJL1t+rBXRBu+GntJI8AqomVDno7GyQN1ov4POHmgYL5
a6lIgoqCJg+WwqzsqvIMZYX+jY0EaZ0t8PcOap6y9AMIBGDGwyHG9ePT4CXr3AmI
3vvUROzmnoIT/wyaqwgtZevlzDJvJPozS06E7XyL+TlJ5biWf1lFJpEf6A1ur+U/
omIDCOqxrsUEEFdrQYhJjQdvp+KEU/hzi0TvxnPc86PTzDj7akADfVgDwuAjEAlq
3rvZUzYIDkKKSVGlZdIOyTV0d4CBXOzNnRnKMH3R8WPZVorwKwO0EHS426WPb0SA
foZ9cOQxA8v6EUW3wAcz9DuCruDF3Rc2NdskVxulh3oqACxBWnIwe/846l+Pr40U
Bu8skI522LwgQHq6vEtl9Xn9e+/glMIXe4Jt1Syc1pPnXLAcGWY9jv3/nAYB+Wii
8RZ/ZYYSi3Y2b7c0owZtx3NZGwmTum+Yj2/kxhhJj4LmNGfnJCO8g6s2jNweFvH2
eMs7/IuC026TjaHdod2XO0r2KN4Rn/iHkWDcH+TzvVxahcmC0RrlEga8zmFTy43P
oQbaC1R10gnymRmKA6lYEmMSlwUVbeLXXkt+/1PnYYNWS6eSfx1Yo+Jb4NpkA7ha
U/SL2CVa2rip74dC0pdITiMp+IrVfm/+GnJWEakoiDZeYXUJZRt4TVgq9UkX10ao
d2KOX0xzk7nvq3gBS2Sb48Vage7kATFoWGxONJkkd76KG6QsJlQ8hf3mUARhlHc5
xwGEjw8Mm4g9ffsSuJcmg+k/1uZLPhHpRuJQjUwKTgjYDnvrNWQojrCiyF7kaoo6
ARCrjUD7Bmn3ETE/AYCoIaQb3LIpeoVrwpHQck1Xc/wN+WamrDZ8OSV2tzYhUKeO
Sh7Z6TI5YtAgLVdouyR1zEdEIcw1DWpOAitO8DdkEqVBSwX4gMG8v8xBjxVSthh6
pOeBb6YuzXdhlmN1C4oUmPIwgNlhvSdfgMLcjTrV5IHfpDWiglOgFJg9xoinLbzD
2xNUHxfhX4CFefLd/X4vEV9FkadlK0yutCTKO+a1Wyhb51J7+GTLi/LzQu0XMgTl
xxp6itHM2V6n2j/UeGTENCXAEISAphwtzCPQH2pD05Ti/4aFmBniq1haKU+uDUhg
9FkwNyz9PtyKPBbFRi1xXwcuA+sOlH/1twmbL1yGbyjs35btXmAV4LIae/AgmwS3
l4sNbpp/71y1HoyGKTctUurS6/T2enZ9afFsk2BY8dxvO37Ndk6p9xtTx4N7qqC+
y8V3leat8VVgsEsSAbF+hgcM1u7kmtzJG2bRdqfw2p6FZI3yelj6HfilEjh2pily
l/vYnj+ETzQzsX5C4SOCCYm/N0yvrCdRdtiKQOo4eJFfomd7xWJVaghcwMW1aOOF
Yvya1Wj82mYvoEu9MKBxeXuHJDOwgw+lyMD7sn1+cPPhU7QtdjPpC75ennF2tqsR
wzykDlwkEweCptCI5/TJ+vc55u7Te/J44Tgc4PPWHog9OBm7MFp6GRUOBZHiZJZt
FAggmNwHk14EOqaw2kGB1Hze2/Z1MTRU+2dzcA4q4ZuLA6ptc3STKYLNGYeNvACC
RbsNXfWp0gwoSxmK0bOPrfvwDrJFq0O/9J6LG7VQu4qR/xZnV9jD8Yt0Jh9LlsHt
oKXr47JtPFrMFcWOsi2wcn3YP0W1dyGaKfrBq+bg+Fwr4IaBi+CwnlQ1BVTMfLeB
7DA+VY5xrSvEpu8RLiwNNKpUNVVXVsyncyxhhNG+Lv12IINLsnrfDvPb6zEfaWuf
vFSDrgA4xgiKeTtPUYxL0GlvCA7QWXCcUKly2EUOVMx1vlsZ+KPXa6zWJ5xC2ZIh
HokRmDZflIghXmdJjplLmOcs9abBQuz/qKq77hvIU2o0fFkQPurLxnl9L53gWuUP
1TKbpm63uBoS171I3W6rCeg0/Ck5aMq47UY8LWbFCQMJiMYDXNiqgDfGUTfpTk0J
dnKNKm2/2PeCnvtr4FY07L7euFi944El3WgBqBwDAtFTk4YMmQieFg/cN9A3glcm
SFmFZT+ywyR1IxLbI2pOvwsc9dQ1J37v4xpWWrrFE8tT0w7kc0eqRBnsqBDHsUc1
8dFeOpkWGgyp7sL/WZpEYFzfItYWlwsTmXnRcgyU/lniNE5c7FRV6Q7IJ4nJ6F2G
MSZA6ECU3dKo4Eyj3ithIaZkxe4d7cyB6pkbXfb4YLpz1JEcxQTBLtLdLrtnaSb7
1EZ/y2doMvlogJ0L+Dr29K3SlzeFFnQGrtHqI063G7FX2M0aXuQR3AgfrC2MV358
nd8zdDG46bRvPVhHim+TK0dE5C9lGGcpdRuMnI9hub4N4KSIwhicgvqsZ+KHnU7H
36BeOOsENa8YhVD8QNEDva2rjNi4Tprysfohcj8z7L5Ctgy7jF0F1LVVEElfrF8K
mxIuZgCRT/7IWSwk3MwKvNiEMPKfL6dhUsVrcmIZhL5QHoA/txgmRBcaVQflGe/r
rFsnTAB9mT/0ZbnBPilj13DRKwmjxOq6b9EIjWAl9kpTkUuCnC3z19cgznv+LXYz
eeyIw+dfXLFSaLhtu4HaAk0R1ZAKTNopYEg2D6R+fPo29SoxoZELPMwU4FMxH6ig
0V0SLgx3bxEPbP6/Fp1I96x2zQTnWP7uK0t+isaEaDeOSugFCf3gwQNq8JrVoryL
Udfe4koS296QlHt4pn8/JzL4tH6G7DVZTjyCVA53k7GPodEI4/Cg+nDJUDKjX/Bq
GyFgVwTtZ2MWOJTGa4GMEiXErPWHYbeyliSO/+dsg0R8ya9YnRx2axLyW2ZCDc5b
OhqwRckgy3mcBX7B4FdrqUTOhfpos72CGEIfG5DrbiJ+RMD7y8MZQk3Lo8EVtvil
nzVhMf0zDznvkWGIWninD9irDlu3+AppT9oDA7WIGmR82snyS5BpRl76aakcSOpw
vbQ/sWZgEznEzXtSi6HR5VADk6uAXub6xNAKLHmwBKYiYzWde8vLWwSDVNth3/4G
TTpQXHJgB/WrhJEJc7igCZqnx2t+b12T75UIG4g+M2s0wWmdp0Za32xuRWBouXcf
ZJXze04A1/w3NJxdR5xm5Mvok92803SPTvE3t9Ky75TwFUVf5ryJlly95SVMXBWL
a+5B1uPv0EOKDDMg+BxnwYskGImD1h+uh7Pih3gtPwM7PCcA6r7zmom+z0hgQQK9
aTs8AQogPicSjUJ8pn3rqdYFaG9Kt/xSXhBLD2krjV9u99u37k1ieIyXiN+S2Lbx
7YiqG2a0ivjxOnYl9G/VkHkZc3NSEGbWzgGcC8rBu6JVVjQ7kArtaODirP3JR9CF
/PHxLfsBO2d/9CxgpSn1FFSA0GKMlIT7F4PDPRBXfy2Iusd8n95nnrlVDfHgNLHW
2v2E+9cg8ArUMS1I+sOITOV7ekMWB7yJxfrwdgEbtGLSga5Yd5r9201rloW0EnRv
C5tHCK8WxaWHaEAh+UgJ1GqhpclQ714mhZtSO43W/fRaoaZtAbPqtHEJ81Ai49n9
1ccDr6SrSjGh0BtQxfvSOPkfjsHYb/Jn1LzmcxFk7v9kpVAwqfX0QSpVQiTaP7/p
b6SBSa9ZyovH/EGGiUrdoLOFWYIc850aWhhodaLgnizkjG78V8tj+Nx8XwmHB3G7
hTvB7uvOsMV+d6XbnH4quzjcvy7fk5x0KQprPRM5VZsr9xNnv0tPukK4o/qbXkUq
OVUk7b0Oq511ofl51HZUYdodJrm2goMPACNu1LNAel+auuwthoAFXviGsT+taWsy
W5M+0JlIxYc5YCXtSTB4XJfdvDNILK93+H2WZl6zdlGgDxQsEFprZOxa0CyL/fiU
56iTT/DaWJbTH7VZkEIs7IxKVy5E3xFI+AWJiZrGdJWKZCfuQHd6UJ9tRWBwtcZQ
ZUVcT6/J6Eyr7y7rftIe+SW10ECwrwmgrlEIaVcJ0dVQ02kPW0eGv57ven5eKBJK
2rUDxhUIxbCjQoc6PivxwqoWTshN8/daB6mNMd/7C5w93jMrIt9bA6rxdJIHO7xe
XUdC/VwIMrmBhx/dVDRz27D8RUJZSMBLUwg3KBBa04QgD/fsHNJiBonmwMHjVVk4
nvrhusfnyVqQqU7BU+DzQlUB4/2i+012WrvhJhIBDhicC2aaa4qaJ06p570Ngbz9
b9PuYDr/0KsZykCAFJUv1uCKeQTpU7EUxSf7qyAszOpUPLa24AHfk5lNJbGLniKY
VnprgG4WC0I9Cj9+OenIO6P2rUpx6Qi3yDMbAeDpmcnBkfqpTSyLUP5Udofu5V4u
m2HFaPiK6d6/1J6RpRrTplsOJj58//aHclZqaEoIDE0jzLnw/U22KC19VxZVf0wO
ktCjf46huuSiuF0lwQditvQC+l8vHVqYRDfLe6Tso/lhxGE2qiZhfzz3jJCay/hd
8GZ9Zw8hS/7x7z6tXynCGXqvZZf+R4Ta3AAJGqYLY5/BzTpAo8ku54drmR4J0/Dm
rmr/MK2fGwUrcg0C3luvh1AiPEHe6tPY8fONwLKl/jGu51zf9DK8bFJDEJlmkU0K
xOiI3SP+yhDkW39412hNfNH6knLJGYm8nfQPVsY7QqMyZrXx0Zdge9Z3466pB4av
Md0DX8oaosmWHAivRB0JG/Pu06admXE+BgapOO0YaPoXaFTtx7xczTe8UG6DJyNM
DmW6xATqhrME19A5KNpvwIErMOCW1Z8erGN3wsNMQzw3WczCI/zacHcLONZ1TmBW
f4zClQVzIpSsz8oq8/0i6uTSMOWUh1zSTo4muiCko/EdpPDFGwhgUv2gW31oVc0k
U4WpOR50fG8X6vXkoeB0p6dNcpi3vFy5lAuzVImIJMztzNjGLFkL++TdqggROg6X
BW7sCqhVpY1cl4adAii7GTPjDU1UqzCUm+TzTR2Pl79MpkoiTX+9Ik1Cg+Js8+bM
3VVqdiREdWpPkdzcKg5x2jLWPpQvO5Xl7ifo3Z0NcvKEU1TPwXV491jepAwxOI8N
O61bmk2OgR2wItgfxiPGN7KQzFSxUTDyeJSLDnJzDdAqhe7zB9IrXN8tKkPHWrUa
cGkNZRH17UzLgvNdxYeknesWJOeil5KPR+ZBKfNHw3v8K+oUqedN2jpiyKrnV5T/
zrWVAUHBoaRt2tDGdAGDQKThabDfH69ceD95owqTa4Tr8zzUhAa2PP6UFmOujRmD
U4rZHuyV3RtbQcjnxcNXPohg/anseRvkARN9INz1wcPwe7EcwJEJOlh/UpooBus3
im6WH1XsNnysp1dNLk6i1++m8uJl62/S++o1uJh2rKwVIY6CXeLj9XXfjdSW+P4f
hAGEEZzNG9ls/B2txvA5hefDt0dsRKGicT3QoKlXu+VfJeXLaVoBPYZ3Brl9lK0Y
29RE0ScAqnN+ePU4SDXMox1B3sP3BUOC8MdJBaqmtmqTPFze8w6NkpHLVcYqHwwq
8Vi+a4YPcos/y7IN1qksVn5K2tHcRQSG8yT+EKsHrGfqypHtb4G+rhUBy9xYYOwD
Shda+o6rdyBfF3WRB905LYwj79WS32oAbKTgcuW1dKDkKFPpYLOED0CG5Q7+yjqR
aQkNMGXwiqKEJS8AA2kUyeODPeLueUskqMm5DxZcfD2JIlg3qenqMpzyuR1kcu8p
EF0kupL2wFZTsrr+8vz6cIetctj9JWWSLqu7kDQQ9i5WrlvOjClM+V1ycCQi14Kc
nWdXopg3T9HoLzGXqeD2DCEOPS88ONtQPUUMUp+xdA4djs3VSzyFGymxogP8v2ud
1GshLKc0bPGYLvuIDS1jyRjjOb/BTWVbDxvjF+rs1rjpKMVxuHxaPHYHwMu9/rk8
qJjgfbkCGE21m5Yz/5UPutEKrIHK62d1jbsEUPUjqK34nRR2nBJ9konUZkcvC09q
GiO0XtO2kPXIZ07aMRpgREdtfZ9SMRZulvYXyEOtlGQdcwXDa2ardiYRMEeL7xno
Oeuz2WRIHcwvC3O6M48m6Ptwnf367t5TQdvzYBQA7+T9BmHyxdHjtHEc2vcPAH3m
bRx93wYH/5HsZQnRGQbM7dPjee8NJdbsBooRydSEAn8QIBAhXGkupGCydd2lHFWl
DkTOb89Rw/I4JSCbbLWZ1eP/1iZUjFdCiPJUb/HXoBDadgokaWQobjuUxNAb9mIT
YiNZRdeOlGpBmIhbkKigLl/hi+rwSGE91vcpl1ZmKDl7F3ZkbN+YkiRCegKK8/XX
9lDeqi9Z2PA5lZB8aVpjWJzXJU7olvQQH0Sr7YgtGdQHnuyQ6hhvwjgTdzQIwdzf
AMt3fDMLPs2Fq7KHghTuoQAOhomhVfzDM1QDxAFSQgpCJhvMh5oUcTobJG6TOO84
JSPgzfFuZ3H03E/HCUxJULMtYS+bRLWOF4aYGx9FPg9oaJrZYnXMA+H8Ow7r4k4y
30TmguPhEfl3bVfRojdmseVB6ffmhwfgVi7ekcwGHix2x6wossnxAePGupHgzbYW
ME3UeJezD4IW/czy3cTCJXNPmERwJtoCX60JU8uWEkXr3rE2TMxEM2zedQt/1brW
5YCLdYU0ClPxof9Jv6DH2Rex+kKC5lAfBLH7dzNmX71e9SxRrQeX3220mSvm4DJQ
XJUnCAz+lTmo3OAsyS5iXUnzvBo99PvT/163FE+a/g3BfsCAGYtZ00l41whKCG4x
7gohWlTkCZzzOaVyOLmgpqctrfpx54C6qLklH3ljKvQcwTKEu4QW9Ouv0dyEHTVH
qy+UjRfEnKqKer6QrbCehQYRfBdWTOpclnnTaMrI4D8K4lvC//hHP1+G79nUydA2
e9HQKiEBsIfRmZgODR6OEFt/huf6XEP8MVeutlngufLD8f5RyeuJIwCtZ6G46nYr
NFmXqDYLpC1bBPBitg3yqSgaQJTI2te6pqYOCYtFPQ3KYRS64xHFdlZNwI01D8+L
NVePxaJPoO4sHjeLQjO+/IWRENiTiVtfciYKnGh25x+25LPeUFIhXbDtaq0gTIXp
McJ6wAlvaHfmrEKfWxvhWWKDRZoMqSOXv9uCwIXZ024qOeKMzA12nJKD21p5kIk6
4mvZzmXkvr8GUh1tantx7oqkBE1BixzUXsP9POr2TK56QNw9ONx9YUCLtv3cyNIG
SMpaA8rY9G+elCB8mJW1WH7pTAqQpJ2IZJg9eh4NgC6PX/9OEbwWIgJSKYymvKy+
RcyYzPF/ux+4Hj7th9qJK+kRvnTK7dDirHsYbPzo6zsWGvrNepF79dieTdlYyY04
DifzGIbs7Bxc4/GRIfJo+FKwif2EInjmEMq483Hlimn5wkCtl//VCAJA39L8Kh4t
qzJ5/gh78SwKGZzxZ4ZtN+eWZY59oA+9tf7Jk1av1rJgsgxJ6qdnqcov0aqM2Lu7
Z6aXs6EqTzcxQr2xZjbsfNtyGsJi8SLUNmEbNnVwth+88AeudIrdpHR/LOtIfwtF
aOqbEgxlexsoMvD1KF3O36hu1jjUQVGET7MiyVjjOUbw6vT7zKG1g687lsOYwDAb
m/TjtcPd6GDGaITBg+HUJtYuQEsomDQLXzN/QAgBQUD9GFWl2oWH40LueC1KYbk5
Nc+JyYElt3J5z6oeFyE43UlCKT3z6D8Rw/smRjvzW1x9bXnXkULYaKgBL2Py8XXI
C+opmzJaUcIxN67Rzx5VGiYPYkWcSRjRU1U0MB7CDt+EqeTyhq3E2/a1Lnpq6UHo
jsV8KR130rySKWMygOYFt9WAUoc9dZGTwZGD1UjPt+dGEfRFOtajFuNsISsI5kHq
ePrjQZb3llLO6i3tgc475AxYJHkXkKUF1Lh0m6q1Q2+q1rmW/XPLJCQuyKL8s0jo
s5uk7pHUa+ZLvjGXKt8/foNWOBjxql+AF/2icXZotyQIk4TztWqVPfnLcb3uqkum
yaFy/0Jh+sqMSFtXrah5xKTqWU/iswjl53Eduyy+l3mQDsNghwcKNOzNY1+TUXhz
lVC2m96HqgSfK7yCt1B1VDZ9Vm4LSe+N5/WzwgBuRPS1sODlK3Yo7+qrTmpqgW/c
HdB3ZJbjLR04Syx5aXI97VCL9pmVnLd+NybM/PbN4+Unpb5+01V039goVPb52QFH
5lN4Li9k5b4mlqIeNktfkl/JdWyNn2ceZpLHaO0QBJo7eB3xsMPd14AewknHo/Bt
cDzfvtaT8LTdM8uf1TahJRmM8osljymlDCHMsUwBeWhzSwdT3nxLYr5N0ZOSgRjZ
I1gTZ7XMtkzjAgyg5XsbN43M2q8XVauSDoqGzbm2H6VN2qRSJc8AAihz7kcpEl18
sKJaKbR1/MFUShJ/oRschGevKGZ88fk+ZfXFby/kFDMtRfaDxDAHRR+VJ+Y5PVcB
pVC3Pf8Lj4JMgqCB4FTewUTJAgy+EU542Gf1hkQ4s1a6fATmmS6Z7Le6B+LXNIW/
9h2XPToYiUo4aGdBOTRcn9MuDvinDPTS4OoWTR8Sy0+kY4bcNYFuw0RRkS3eEiw/
BBTOqMKQyXs7VuT5RDYvT1DqIG29x+eDaJSiUHAwdOp+AiuTOEyaUGa8Ox5yhh9S
L83AsBv3v00qi/XAlnFb0u+MIJjwH18iYeLBZjro9GiwNzo4uH9v+vc5sZTlfz+B
K0PuDGlnskmhU8hY3lX+16jNxjbH2N2sQXLLope/gKSqR1d/Qm2RP62zi/2lk+mt
Xy3ljgVFnEZRaWfVtpujataPEY7ZMyOwJ72gpFKjYNTkl9ytjgy1qWe1/TekSQZX
4OVpMgdtHIHo98bp/tDRF7PisHhHBzVKzIAPcIrB+i/EyCfecLr5EcXuXgbIoAJN
49fIj5ETydc5YXkFsf8okzRiV/UEZi9sMTcXBr2ksGa0xh96Ja08MdgASqHpTJzD
hFBKEXS5og14G7qqgYFxHmqiTUF01shFTQzTvIJewqQHXGorWwv8tvsXAvz11doW
iSG9H1//uO94V7kpAqXzUoICP9f52bpuqTspTsCkkvCEdd4LgBrJsQl9mfYiD+yg
Q/x1OSElICNjq6seFx9+FaqQIc02ots5Xvlqdwr/sgF83iJaXn49BozqSLHg/bdi
jAEGyioBxfC3iXRUYHgCKrusLbhH4v8+/vv7xSaoIh5EcgmX4Au1LEjHbhqO+4RL
MZ6TUeiB2opuhMHlWgCDl/dX8D7k0LN9e6nr8J6JeV/RePCD6zBv3FIJkDHwYVel
xbOsHLYTHBLlBVNmHa7CFId2i10Bylp+rJGVzioMf5A6eX+MDgrqex/9gW+nYOmU
iGa5cD2Tt+LuXTezMvVRy6+lCn39n5i7fksOvkhfDxrFN4JPpzQRyz4a6mj4G3uu
FMMFolqOnwShKVeTFoDTLYyvAOh4tp26TwpEYa3NTQYFzG67R0X8dE/YnIz+X5Ib
yKd8Lq+WTdE2GyLKa5CQjVzYX+0oCrWKlw67R76AHhcS604oAMT3qx4djQ5Gp0SG
Koxo0apHJXg4nMUBkC5ZuxzOkNl5Pda71SY5w1ajfrk+X1swU/JuC6W9y+zXLCmL
Vtc+psGyc9RsbrwZcTsRXThW1kUkTnpmoljQR4QhfVqq9q4XPuXMLDhElB32xQA3
ns2qLiIzJsQ/8DRJ+cpuimXfe8GW47KMgf2SGi5yX7u0JS2awClSbYjGoH7h6wVA
mpCaa2OHbaCo4MdMDOkTfQupFTO2zt0Aj8pzBb20wYMc5OoLjr3ZMYief/K8uUOb
fGh0YpLiHVE9634qbH+LyF17F1BipDnXGjlQ7iARGvAoYDbvj27ou4VobuKLSU8k
oDoGxDuRVFy2jJP1403QjF+QbPFL+cVPWZMly5NR0Ki2EtpOtdrkKbCcbG5Z8eK/
aK98I6mHethuOLSw7vkKJvfwv5djZm8R/535NxtyofwIjMcnc5MCiKBI37rYjuMl
AMLopqqdAswXHHIKNqmuAjdRkopPwy/2tHYdHuBGTGc0lwNT71DTUn0zJ6Xm+yPg
1GoviEeh3xsoWWOKKys8XB7DUWKBVwWgWyzakkOObExMIRU/DOqdLq2olN9R2pGZ
y0GC20kTo2lxVDScMycCmGCGzQoyC/KOF9SFu8X+h2dasbUJDSiYgX6ZuLkH1okj
qyYAoedCsRijEE42lba7L6utbYnnHd3l9RUkkyi+1sfZ/Zwg+H5ls5IiDNwIjlqa
dpJFSKwfJ8Swu+D8aATjYIRgkt0y5Ls5j2bgSI+7QTt4Ny8M5UvY74MFvvxz63ZQ
xkc5Urck4HLIwjzAkJWgygHA/H34gW0qkz0wPVRNzwy+NJ+K2DXUuwNqiNDimIeT
VinXZ/L6VYqv38KFlY3jbddPdxC3jygaGCaKA385NTgh5nT8wrbuhZJskQUdhej3
/his2AU0GbPW94ovhSqq4DjOCtVNpaMJfOJ1Dav7RTcBaI9zrbdo36F0+WxVeHbn
08EqbAIbC8l36Afxww3u+cp5be1eYWsUKrSbvtA0IsMAGFZYJAa/8lO/bAGW9LKa
VBl/+5KsNUL/dFTZbDXI6VXwf7gDR2mwMF1z9YB4cK5GXkcllXVkIzTaMg4O3Atw
XiprddVT0EVmZc5I2UlJgBwj//OvBH5TrGI4IlGl6e2jdKXcxInZI8cu3QSYHUv6
4cuCq9xomMZmdHoSwU7ELxUesYXowAtpcCETNMsT+LVlyipyuv+j6b7knmH46imx
9SC1FevxEKycPMIyJ8MJDYRxbWh9b/nBxRgySQ5nL1ha3DABzQbe1l4QcgxrcCBh
KhRFBf9UBfaSgZDNylXHgGEIOoqQ3sglXeeVGkt2QSAQZj5U7aeSGQx2dTyGPcPA
gRGoCGvaUgJ9NggFC3uxk6M+bZcKkGLBuSIaVfnd3RuxiGlJ0MhwxD9UkVo9u3Eg
KqPyqXEgeC0c5Lr3OmWALvEIsCvo+rx6GVY2ayCTCiD4wK8X5TkBMpvy5lrfNcPa
2VhRtyrlRlpHGTZdm7G5n3Go2uqzIe5id5t3X1ykKrOIJtta6+5PCY1mEMrtxquA
o6rPGct2Tcou1MnLzrndJUi9X9nNB9sNhG9/i03sOKsXohqKCpKE+A0HX2pJvvj1
uua9YJSM9ZeI2aAlP6Na4dyo4WhHyx2xqD6CWE6A6027iQ/85s5V2yr54aNQNVpI
BUqnXFTxKn6NRDrfHzCSWPYm/sbWoP90hLXuAbgrs5kzB0qooQJJM8jFagUOznPC
68VYEg971Y06EWxAQu6BgAWADtDLGJoQ6YK8+/vsvJAag1gdrG8PMrnCPF5FXbCN
CEZjsfE0wirrj5trHomRsxiO+yBA9W/82BIFchgbbGtQRhLxXqBspWkMKLAp0v6p
lOs8YcrlehW+5V9YcwApySsIq3wUPEPPuygfaMSpdzy4ZYa9Ucra/OUkxFwlnNPs
lzIvwdRt/8jhjuzN/UnlyC2zRMRFwIGivRfKRS0lh8ui0dUcz/kRcw0PydL4WZg+
XDz1VHwNSNMKpX9JSnnn0qM7OEOf3OO+GS6XUT7Hw4IJwC54muJ5H3z6kaGX++Ne
xg8KvWaZneK9EnRb+YMOAFhU/oulqS9E7Zsw+DID/HOhgcbeI4Nay+fUkJ4ecXnH
Qg6MG1mtO7uBbH+AF6BvhcczD7yYPsPAvbhclN0xhFWHxABWs7U5bWXUl4Gm5Z6H
np4OKPCruJwYnBLTYxhPefBeL7TurU9dqmN2xtjjTCYYMyQpVb7RlAY1qz/CjCf2
NmnVJ3+Z6qxaTSl5GHgJBQWtNh01rcr7+jdKMB+pFTWh1QTMaEHTd/tlsjdIW9Y/
MPNEgbn6YWdohDxNkwigeF87Ke97oqlmJ0NxW5HO6WwGNUERJjsB4TGWSdQPGvgO
B6M0FZuS1wDzMY2ATz9xxEp16Wj0TJrcINdAO1l68BwVh5xOKTuW4fOONvhf4nRt
YtVJYn+QQHmC1xdK1JE7WcOGgeHK7kyIpbGsWTxpQ9qhAb5Gc0iX7pufB0qLajiw
lHe83NVUy5RaKJEFjjV5TkUGn40of/WhCPKQ5CFVqX+hhwrZNHWVlEk2iXJ+sJPy
hEFS8mGMJguqaR8uKc5hYQXM5CBrUbzO3R/nagiQOqFqQzRRL2BSe9gIHINa8ceR
CJCIQJOE53EHmFf2BT2BYw35t3TEJQt1gXYhahRE4KXlwmwTPmVUkSo0XQTmjetW
/pRh6U/3+SaOxBSUkPPJCCT60ZOdjTC2aIwm6VYzowj8OPo1FywzmVyxEEzInqrB
hNlKUGoWQCtgwiZK6bk7nVs/DKJd2vcbl6Dmtuj75KzeXhSZwgeCPJSncHyGW8gV
FVjz6Q7g3gEsrfqDZZ+vmaHZGlW0Ij7xt26ew3WRbiAfrV03Poy7lJtOkOMW2TLi
SKPgM/Vjl+Cq0t56sp2b+ppTZ/8jJ9woH+NDxtAbxWv/O+b0bXjV/Y4Jr+PQsOjw
z/arKSKVhM2L3QpthcutIWOx6DkszSNZUaG8vrAwgl/qkGDDHn6tUXqPEkegFQ5l
RVaWpQPJ7CC0F5ApET8bDb+m4pchEsQxYlivLup4hazZ0dncxa9pc6uElQ6lnHSD
/dIvA5ispqHdzmGON8+mxkpmtU1MdActGl+k1eU7+ux5JJkBkEWI9776XYycQ/qx
dvbvwoBftb9w7c7vXz6Ft8ljF8H4P6CI2DyF+TR7hxryFK7xpU3Chl7KOwnN9K4G
cn9NYPKuxONttoe/FBcXnZKz1FLPna2ZHlHBC5/gPCWQZp9vypSFRsA905/e4KrC
Kyv0MUW2NI3a75bs0eckmuQ/g480/tKKgysOU/AqsrcPOSj/fY05b6jJxkUDHbo4
Ic5fGU9Gd3tSgvUYTFfDnKY9BM7xdUlTV8tWjFVI+hNce6P98st2tkfoBUvSQ1Vf
l3vy96Kotyffw9VddHb1dx9/qWmlmpx7iFmNu1St9LcgIe5wDvDFjn/bMx7UVDRV
RFAqsetQSUxTnZ7vj2rbJBEeKVQXUjSwGtN3zF3mL9FAhWUlS9jBPT1/aSqVdaJ6
+JOS+PvLX/7bduUYhE00kjKEeYSGkqxV1dTFpmhFv9xcqQp4QHOsv9Qt7A93hmc1
zTMhDcyObvPCSdAhD41tJQj3OkmWlCatr3PqfAyZRviCMIypd8MSsAyMTsdgbljf
CKwyPhM4P/SsgyiKUcll74maG746RiSw1IHNaTAktszJP0H+PXzoC2zOWLvt2m2G
jm42w6htZA/0QmPkA97Fc2uglWMBkfNoSEyBlpfA09BByo98kExgnfDExdq1yxrN
nSyyP13Jy/696OCSXYIxw5pjsPX6SbPvskITRCTNCflImCSM6VnGU2y9FewJAnmw
ky8h7GQ6aqDEPnrEiTgK4fznF8H2hs2f2HtFijElvj6mR7dSr2fuHx9qz8hIDlnn
DyzCLJ19BqOVDnlG9p8ho4TgB2bO484gz9SJvWvsqisNUY14JKRJLjatM3k0t4y/
8M0G/uVDG2Bb92Zh4MjHQk6y0+85Gu/5UsD/MOvTILC4/GCvK1BvNzfJ63Omd1rc
Uqt1mvklwTuMmZYDQIlGa+s2FxNBDi3UaOcdSdw1BxBONiUQ9kHMwgCyjil5jt63
FKHcnpcHY5rTJFMbTpVGmb5Ki6zMdQ1AJgbV2ZSwOIymaQ+939k/N/PowGntHduR
vVy9+z5J4C6xSq8NyzbmlVzj2pMIljHiebWMpmhA2L/Vi37HrXeIg00Ky/cJAkuE
BB4XyKotZz5+8+xm2pWEobJgoIunErGpPkJZYu+heWxZLCsO5GD6xPNTNnSTwOCD
7MnQrn+e1iJeU2ev7xPc9cygggJEWyP3NoXgBC4aaiCD0/BHFOQtFGJYXveczP/5
9Eyp+BMERN97sNbZ4I/PPxf2vAwVgE4Fdy6Q6e2lN7caxNfu+4hfjsFyZEmXvhwA
uDo7FqX5K4D0oflKePbj70PKV1+uKDEcBssUSu3TL0/S4YhPAWv3fZrSxKXTEBT+
NB9zTlk46iohIQ9SmXuhBIdbr/M3h+6f0n9jgIpnoIm2OQK6uav7d5uL59XwdQQ6
7f8y8CnLPWeArKbPpeuy8+wrmLEiyrW/xMsANWgdDMe4xQRSS87uMYRl+vVL3Wdt
0Nh1JynQghGWt666p9PV3hYzNVcMBq/5H1chGDmo3EbGayItdDfIWJ/EKpCVcMVu
tUvQTSvkFC3H94ydiVnB6rJBLnv0frOsrfEW71jNKbO8pU0aW9zjIOFYtDHLGERc
fgKyDH07q3NT1KiUseqUKXmKuqS04iteJqnoKnbWzBOnMeJtBjK3yx3AABSpZx7r
REoBOO4FxaofSc3qwVXaJtWSHR/wV51Au22i0JDDNNLkDDYSsdlTe2tqkOxaUDrT
RHNFfsi0CN9QQL5z1EeZgrdpewMchMGuEnKAHWbO6XbNNuwv0nBYO/xAet7tT1s5
29YdWgZ+UKnPmCq/HQwzix7big7G7lK5P4Wv/sHvKh8Zx3aIbZYehOZi0uzJOrcp
o6yHmH32BcIgDi5MlPEkeJ9/2O09pArR47UEnZoeiDCZuW1nl60lHSAHIT5PkUj+
R9VujYSSlNqStTF0bTt7aFMGleoDvy38MpmZPnmMGRiZZ7bN6j0IBr/+KMRLrq1a
cohW+spHr1ZC90IP70LPhxFWVxsICKlMfSHTMWO/LQczZX60IUU0bZ5yFka58BM5
SsBEAHV4EZrC5wTikZiV1gxjz7Hdfr2pHsXZOVcBJYdXMbXVJwRZ2LXRA5UVxTAj
n4D6EJ9Mu9GfMxl6Oz8ERuwXJD55bg45hWw1+aHi1PQ3gcUXeL1DVRIDcjUhSkZt
4PlBX5qf+DjFwBzwelIPz74pvNTCyBWW+Ta7jzWlx+rQmFmrC+/BeQ3vvEZijkTF
Am7SwarO/ZEFERhZ+aPSZ7o2rbV5tnPBlV2E9ol5eEzdlDUcgJhO8bNVCqorkc05
kl4jvqIhPPoK1jMwEEnHltBTUHoG1lonfAPU6CORsg7BeBEu3zZkL1wIX3X24LML
d/AvlT86mVL/R6FTbjUjPFLbxf/VGW/x672Uy/lUNPU0lME+erJAhV36biD3w7yV
hoSctHJiuOqjMqIosNTfWnqVzeo6UhMKXmMmS7IN4TfV2IaZIq5i54bOIf4OQ+X+
sRmuJxMOgv3Fw7JiwWY6fHuZnr4Rbr0oDsI6MjdvUCy1NnmlEySP3ojn0xvwD26g
h+zB/lF7g+7kSho03tUoJ9nVDTkKi7q8qtnTAwebfu3KWtcW1CfULvVhsYaQsthj
09GkwVrc+JJm4zCTAwIU2btjF451wGWDHYpxb8M5it06aXvVdTJStf0U0TgSUkn5
3x956zLp+UU61RmInvsnhacdnIlfPSkYmZs7pQ79DdG4egglrh2dMOHO/7oMhjVU
vRjdeU7NfvMXCzdQDfTKG+bdF+4qpyuKCabcXMpQ98/oQpHGVwX18rT3Xcs4GAVL
b2s1xS6Zup+WT5MX4uTASKWsQlbP96QdW2tQCDP2X1ZJlrRHdv5synMvMugXRfbZ
yjMhraKxjD8zIWbvDlkzERkPXacph4W1oIOqvhIVa7wzxo6D/3Y0u5SQQprpMEAn
3VjrsvFZYAo492Ibejsm81Lw50XwebgBzDI5OqCaM634Z9507m91b1DTBjhStgnm
ZR/bSbQtkkYx3miJYQ6nhG/lkK5uipTe/fnQapxHRf5N37IH8dM4dfszOCKUmKUX
flXqH7CDD3VIiIprNm1Q332ne3Jo9Fy3hpCi+GpyVmgba7UBTZcCk2MnvpdzZPMF
wMe3bQ+P++cL5dXMtSD+JE5J8xyD56Dd7rBtZxNPLKMonwK6d1E+Dts55jGPrSjX
O2uyMR0o9ReUhyyA2qVsTh/6iMAFDwvjeNyxvbu/ZOqoOBc4g8gMOSoZKvVPC+M7
56CR0Q/m5ndOXX9FgfB+YqPwukoBtxeeftpEP0QbUDTyn3r01nCgaLjkcAWWWvhF
hnaWX7JlcCQ/2CCKmWqrT0sRnVShHd7lhQqV6kElFmiGxxKbE544yVXQfzRwLZ5P
U48TS8YZGHprHbS8xAAjfwNPYD94evR2etXXQl/gLFjauwQefSqrUN/9a1n4lQ9T
8wDt2yXudHMisrmgT9ZFAsgkEx9ZPPOK0XqNGLkSLgwyGpfLSDT1vHBXGmldWsyQ
JtUTIBgxRJS8Q0q4R0IWWfWfuO9F25hdk5VSkb/bz5MtP3/8bT+jSj1rMee78uu1
kz8QQNQwd0TwtF/FQaVeZbo0ALAyDvo+OSJE0yQmHOTar/BEckVne+TOnn/WXKUw
aWvCTipX8kLVcsLVYtlaH4BhHoLr5rXYVBJ4RiIav/P8/S+d4122CT6Pyd3X+G6u
X3RXefVfpNLo3cOvssSK0Qenjh5O+rmKm4o+9+Et6lr4EJNrH9s3mKhBwA46jvOx
cobZq/CNQUcP3GnsCYhQDaG1b4jeRZOsfG2qjvOOGIfrlQIwNCIeVh74grvQsUtW
X2242qtLhyPSbHQjXmT1uwMbqw1RC/wK3pND4B+SRQat27xfFZaNS+aZ2oUstQPq
p0OphRPZAqNJ/hgO9HBGAfm1UzSWlBYENN4itJIyALtqFcjaYd/FfHt7pm3KnXvw
i1yIoIVrdzt+r6GXUFPy7LRx27HlsHBHhSmcfZuLiRKxS+mICb9iLDvuFJPDSYju
auGaqdm5j8TdzBO8n16RBVGEY0UiedXKTGVa6jBAlnq3zrzT3eqESVGPfFmxEAB2
HnJqcvBAFRfNk6rqhJzoN3Ss2MgLghMxaGxM+Umt3r9JiusLeOSRAr7SxR2FxCx0
53TRhEOBbGu/gorsh79QIk9Di56/wTtNyAPXzHMioNdXVFODAVApUqjdHXvsY2B5
PN8P+YLgTNtd9fQPQbyCdAA50RC6uV92j1IiqZGDZjHI+rih5ykwTnqcDFy4GDFC
/mKVQshNK9FUYWRTu6WqF7snAOrkdw2JuvSFiBtPgxG5GCjYMR8AjUqQfGLYt32U
dIeC7RlnUrk4SnTM6R9istEGVVHBw2s0hSrU3H+hlzG/htfK1Il0sL8z3dTswoW4
BT5tz07MVa1rQ/rN4qATTI+29eIbVw79MbXj7VQ8PjX+CYSbbgJs4KMsf8D+lXAG
0GNtMPAHespYD93F9m3Uz60Ik37k3X0amlmyfMiLOuf++kq2cO7NQCDSx8XMf6lV
5kk75qpdFClhmW2wkzraE/J6LCw2MwCCcpqKZwGU+2GrpI4Bbs6aDGEWKhc7jNvK
KQbzUfox9c8dNBgxwNKqo3D1/d5dZn110aQuBJEQh08wU5Mbbi3y0giaLeO5U/6A
lu6hi4YYnrCGKr7WVBjFr3PP38LSYTB6Bkcde/51OCZ5MKjL4vHYcXjLhl67Fj6O
/LRksfwIEdOi43RUfWPzkAOT1llKUh8PAiTSn26lyyD0svc93speJM7c0R3oukjm
CKza77JMh0ZxVPt/k+k8H6ypt5VFZJnDz6mWueR6/E4FL3Sclq4HnJRAcb/eVdOe
DqBPWLwrroK/6LsLs8L/XCysmP6L+wYZz/TWI42V+VveUAlQNbTbj3Uo1hzbgEuV
MHNiftggZvjrfX4OwYE2jPslRm9FHtIRNShjN7cSOmSMVvIk/atU+uwFid411n3r
lLPjqQDC/CydWJJChQgjKp2htVRpZSuazutPfXkRY33W280VpPPdma0UwUe6Ge0T
dRwvQdL94cl3nkd7GMxpD+olp6SPOU1TG0iVGAhDp4FO6r4jEV4Jtfy8Iz0UK5Xs
hvGATMBHeBq7Lo+LWSYz5+CljNn//rdY6UeIrh+X3JC6rRDtIRxGN/1q/HNVKP/O
ZEyVif0rzNdoBqlD4YvlxnfcYFswNHacTp8+d3xPmdi2bKrEChlbmhPizkhdbsit
JVZnBiisdmzVc86TJOcx4boUrmuZNNQKe8xjY7rVfnk0smDSg/Pk8CaD9RyTHO9u
+7uqADe5ozjos4WAE5de4D49LW1WqsHqqfRPX6+xdcUj/u7TmK4HaqRaGacktGFY
3ayZP4EA2rfUTBK8nW65G9ojgWBPynFG9pT9dpGJWY6CrzOvzO0GG6eCrD4OhcUK
ICLwk07wM6sJp9eOtLM9S4vNJz/s4A3xnhW08QQeQtEpkbhwSbdK+N6DQJWSJWo6
kFLOStp/8sKmE0IDSBVd61pWQfAWvgkyk/8l/gZG+ndGlA2fz8d0CVCGiCnQqd9F
MHnjc2ms7fm8c/CTsnsIPiaYEdLyn1hWAFtdlZ9FFr0rzLJfcAdo9UWiZ/To23Vp
kSRYGSLKEP56Amq+gFVyaDoWo6TQKzR1eCUn7I4ufetJtUfhaQ/XqMg0X56yQeU0
bDSrPPlQvoStRvuLWMbKdcvXgHfgMIqLJEoaZP3vJmP8s9iHr7kU7f7R/oZRXaPg
TyUNsgcVORGiwAFbGMKAtA6bai0HUcSMI5EoE5EmCeTyBxedo8StWd4skrJiO91P
qaqEiT/x8mv3rfUlTsAuf7mLZATpg7iKMjezzOQMrbXVpgAETVzDO7WAHcqTd+QP
+VrwzAFNvIxlYzQK7zlds0YL4mWy13oEK5zGObh6E67qPL+ExXTV9kzAAw1Lf/Kx
UHmlmcD6AQj7Kdk7d8gji3s8cSrNVF44gZQnnBRGoVLeSwfn2EX2no7LzYwpYZCQ
KaPP2lyw9dXGJUSlr/Cx5HhEbtmAQmW+VZ9BxXlOVo9F+kS7fCamuxXUXZWLqS1Z
JQcLH4P7mIKYQLImW1LEwE++9r4Gf0jknORY5U+Yha02YYTqZB6tbZH6WgB9+HJx
BV2dm+hw2IFCYA6Ifn4DVs9Uq12lIekxgjAMe2R51waeuePalEDrnlmz4rJI0tlB
/COotpR9bE2ueei5GMf5p2+mdz9dM91ZH264twEnQYmK2C+D06bdJY9rITws/4/a
iH1+VMOjyopbsbaPu+4vdjOGBtWb5lbaaa0vFSviy1diFSsnDJ00TIjhRJbKmJOa
zyInIMjtwvD6WWtPLL1oPB0Rf0DiCSgb4bzFXdwok/a9Du7NXFO7QYI2AOVlYGAB
hEvxTCM8lkcrH/+iGc7ESinjGohkbbIKJxKSpMPpxMqM3Ksihu5y+A3q8kcsJi1e
5qMpwb4uQrlF/q4CY/07VVPTsu2qo59hflv9OEb3HPtSzRYkv5nNpITfnsDOWbzX
h/n83tYYRvHmnvc2kWpWeyz4eA1XUfx2aUdqMAJEJPwlwUypcXVeWtsV9hY7EP7T
xMxkF2r9/T93d0tmNPcwUOWvbLYlDuDoMnfRSDidjc8GWMXUXE9N/kpvh9svyNbv
FfpiUGTw05Oo1VBVq/ME3uYwPXPmey9JWRZmWLNIci/RBHr+5omQcJPBpUAjR2P/
uhBntj7FSCW7Kf0wSiCrtWIfCG4H/wpRN/hQ7yDrk/AB3JPlCs0mLoF8sA29ByM8
H69SAa1nyZeirN4CL/uTrQgibUAql36kCaYDV57S49kK8+x8SEIC/0k6MIra7bFW
KNHKgU1Ya7/iy+aYukoaGg6F4fy9TnH7adGLRHZMAa8fj/Q9/dqfGcyQBqyiUh/+
pgc/T1pkH4D4ur+hbJ9P1J4qVGrBRPNsHCYWP5WAhaofE8mrtM+G/7UwM8iLeAQN
MGPwiyenDhRLnYZT4WtGSeEsZ5iJoNz3s94LZxeFiLYvR3KwE6BuvkABpgy7sbIb
1ozul/pxzuBzouqEGErf4sJmGrLDKMiW0soW0oEEGgnYWLeVWy2UJXyDB7KlpgTj
CKII94bMGb4F5nqcGg6/qoEOfwIPKnA/vPqgl7CvhSFu509jbVui2NVpwc+yd6o6
rb1R6miWzSlBctgBIWeCkaag9hyv1874JscO1ylvVobEZoiCZnWAe4BjmqVb5Ccf
ynF95esfcU3UZKXY7M1QBaAbSoVLjUH755S+xH8Udr/teAI80o8wV8jmIYFybK0V
h5R3qh7szyOEhOoa437lAs5L3Qjafj8kea/QEYaSbDYYouCtYCQ+0TJZ3vlX7HHE
CgG/lsvPPDV70Sk9sLyxWQL4GRw3giBekiSn0KGvge1milH6UYbY8aDp4x7iGhg8
Ozboe/Hc3qVOhP+kqOq3mvg4+ua33bant4IlhcUZWtV3nwsvLx5QYh1f5tgnydzO
ERs4o7bQYCs3+C7P4jPULUp6GvP+MF/YzFgcptpHDLSFlmtQQevrBzl0zlgV40di
4qHoEbOhsy3JdGjd3aOSsyV4cGtra1HCY8/r0EcT6AWPG9W04rQN0NVaCMkENmav
8oEDNm/H6hb2upv/JtgOhK/z6WNNofKIYV3ROBaCdl65U/cB0+y9ZiaUd5bwsDoF
kiTfFA01n04bU8h7IYoJ8K8zjIJNOXAfkmQIk9SGCmn8v8jIyW9cCPFvoNbn+uF7
VUbUTjj0ncgORob8Jt7muO2NR4b2zU5DW0aMrze7uFlEKlj+Lk7Le77JjYC4N8UM
kCPluipfLb3zHJsbc0oE19XPJ8+ehUEhnbjYT/2k5MQbWpFW9e8jk8qbDFmofHsm
ey0rkhPJhRMFUBY7ifelhM3e7+Jg7+t2xlVOWJogIirdM3FSQrLukXppGDMrnJGy
uwhvAB1uIAw/VXQkNqAiEOYTwoL484B7aq2++lB0VgfHKPGrswvU74QZJz9H+iCh
v/Rv1QTqBO4thBryR0xiaLoI7DEIlJdDkw8SMWtde81YkDPniOrUUOG+bhOVeZqV
1r5pWbsRJHl4VvpJswz4Kl4RTGyYHlD4pquZqgkvXUltGLaZLN0uZZHIST2WTUwO
IqJe804tbogeehauy1RuIu4nSwXq4JbRGbXkfVBUeJJf8m9E7pwb7IOsLMGyvhQ+
/z1Pp698P7dcAb43IUECig6Z2IQ29F6kkeb6Ik1zuoziIgES8Rxc/+MD84KL2YV2
cGbKM4omsZLcONbNVq7XHiI5YtrDKvWl9EeoY9RCpraNUhSwazW1qopqU7Exvziw
VCQi4VbUagNc0TVaybvbXJvV0YPogy3v/KEsh+qZ4sB/ADxcdwJi+sx0/7r3qBUG
6tpMLBc4GxwsCohmy7W0roFCrKxGy8Ctgc853B2Pa5s0Z9+/4OjC+Kh19OGPdvMA
RH9E3wym6gArHgG8MzRZM56zrFzgDIsMxb1FteUx9m1DWvzCL0HJBPCstuRJTBiu
mxTaB0vPHDS7FnB6r65fezddj6xIaPowrz69lhp3oE+rohdMyD75yDDPeZ8XWMb2
0sID5zDlY/LiWDKJptrMq5hefe0uyY5q4goq3IU2sfA4nW5EqeEo5t3WJYwI/f0b
+q//KglvHOUq2fuOuYKEThWpXcEZXqCwyc8Yq1kKeX2Xc1H6oiDuYharlIhhMyql
t3gg+QGH9Z8P6zNrpZLYD5Vc2tWBsoEd/pg+/HdLwZloWnRg/4D6RD3ZpwQHjPts
twbXpFfl/BMYYWxE87o5iimYJWAHJ3Vy0H4QbNzwkAGwQCmel0NyNJyRGFlgZalR
812qIfsfgLSuIvgjRbVQE6lz2dPzy96CLmpoa/xt6s+qgO8wkBpRDJ9C2t28pWTT
StyccW4OgI6tshmT1xgb0yLp4zf4I1aXVXtns0zGfb+c6HLEZjwq7hRiH8Lw5f19
DYlOrLMr0n1S5Ucnr6ET/sKqlCjQqZeCZpRu/pRlZOrfuX/YeLvjEf3c1XMiT54p
tca2YYFye3U+KKdiN7Uj+4kuEVpOmkM75VAdFNWKzii+KMb29mEB4CvCWvVicojs
wIC/WmjNVIhuMwT+3ZLFMavrF5Rnwv5pRGn0OUeVIfo3XXsiM5EfrifWO1xJwYHJ
u2fhbcmWpv3x0vxr4yWGWvWc7nf/jiO7Pkk6BDgUI+w8msvpDdpVfxIqORZnBBaF
3h47nmQk+AA/VolGi+BS+YCCA7ytZg7Y5Klj6aDjqRGRpfa2CJ4jvRsAIlIN/keB
ISRUDc2JZ4CWi/879r3ZrRZp2FDZR6Nu1nVH3rsowrLDRzI5MdTknXA5CpATT5IQ
HlK3IrgG8YJhk/CFNGb+If7OU83SeZ6WnUbOXuRRl2aRDoOHycyyuCeSjccL+WZN
zQZ86V7kx2C4BjD+qJt4HRpIFSlNKU1aSBLsvD8mlTxEIub3r9cswYkm3tWchUGb
UI2pgSsHYfKbXVANdLpQ0+5MKUGTMMs3e4tY7hNncHKKtmIh6RpSE9pq92iWA1LL
+9t3DUXEFKMnyOWrD0n3BmrelucuZdc7qn0mymH2bP+aBUfZVpoPc5fxkXEwvws6
t66znGScQ+HQiYTcVA8AAJSRG70uQHmF3voxE3X4rBUsJxk8LJGaTjnBgnr8GmMF
M+mShz/r4ch+kx6/VQklgpeY8pkEpi7H4sHDBICPbg7E75nLrSpR24XE+RmbEj3z
tkdPsSAC3bOfe/Uv1a/u39f37N8AlL2LJVW1VKAFLvykET9V+rC+5xGrUPpNIxHn
PnwN1FXPAmJ9t5g9/mZfOCXJ49bNE226lra4oNOy1b/UWp0wPZKGOHohxJOklKyw
QV/x+fGJq8tNjNL9QA93Y/h5Nv8M+0KAxlibFXIrnxuIj3DMbgZbF3AzEMJKcxLs
WhUKOryjIC9zhlLzCyyygSluV+M9GfTDw5m8D+JEil3X818SzJJk8Gin/EP9D4ht
sqF0pgR2hKR0SZjQweEhRlbJJcHyiuUNzLg1AA641n+DerAADG3lsZkNi3es7jYJ
RgvWbN6BESS/77AneooSk868ZsoJal6ZsupcyH9dPsS0tO0A+aoLhWD9iPnq2bPY
HHO+oXmb8c6V53sRo8gNLsjZRJAMYc7HNbhxtJIf61jfk3wl8y3dMB+4NfhSvT9D
jBezhpvpv2GI3V2XZYaeqHXfkJJJ/YVeHY+HIa9zNRuhDjSZJGbrurRP+JZo35z9
km18GpLq64UgxoJYUeHAKiYs02K99NvQbvs2zbln/KIhuhIFBWNKc6teDl7ent15
dBuZfgTPv7d/K/dH8uEjvsDWZcfDZd3Uri2wMLUsPWrABHvy7RPgWRzsAldzfoaf
SSxDrJNWIRroLBdHLEzHzRRbRyuUtvdibKfUrsiwn0d0rpUTyyZbuVOQmutP9ldA
8CBO7PRVPR6/2xFv183AX8QNNQbZK40NBTzxNik30OMZng1D6I9TkZw1hKIG68vd
dT51GFn2ohTeovXR+YcqTqQXA1E7sUxePjOD05RPLF5zitY/KUZs8QPWFu+W0cfz
B8PPqOm4nW/LuBjcOwGAbAhYagnQKAFYPSmchb1XBRs6tGRXsRkaOTtgzXmf4IZa
Bx/qU/FRuzwmq/ZqfEI0YnXv8nivrKgv8Q2G/Mt9DQRLSFNh11nn5Ux3Bpyrd5I+
kGkwQWVSZq9R01oR6FLbGzI56WXrJIxcVoOSg1SZqHcRYFdWTkuQ3+9ccewSRgOx
ZmHBV5fEkWNV8jK6WwxdbhspyKPte1YjDwP7/FqqDrlqwvAO5eVNQqvSNseEWJwH
N49SMeEBh3bH29qxRAIwIlPWQn596hYr5SEyGX8Lbbnem0u7Yura8d8kv1HROWvb
2XR/3FAkdbPAfDaFLRZyh82HR0kSGYQURm0Zju9sQT6a+zRNjIqL1NzNe4VhNVYv
my8Px6K/uEYu4Ec0WnnSRfSlUJrZ8mUgyOGNZPQUZGpxc1Wx8m26UG99MuBwLAC1
axqHkUZLU938mVgp/yB6T/xbu6rYR2oTclEqpexYcyh5Eohmx9E0ckWBymEJWHmQ
S8h27lJOm0eyHlUbqT5x3sp7jb9hBA4ImuL7zoGao3MzcoY8/D+MagB/ey6koZ2b
1ZC0JY4fLaE9p6EfCOmjpc6NS0XypNCmEiWrri4cCxO3HfJJYqZkto+RbixevhbQ
LBvE3bLXBSh+p5uSlaiVDq9hv2hMVndq9qFv0WUnhmIkhr6pmhc/eyBLpYuK1ylJ
MboxBwg0DIaMt7I3MShpUprnIfZ6MlkX3Xw2cB9tjltAMcVZOq/kwbsW/FF9NRKc
4yqjwMJ7RS7hCLdFMfDDKDyTN0OHUzWFst9ac9X8WyR58VZk4Y0VsC0bEpmN8ud+
ICTpIGGCK1+3ZudpjyEgB94SxqR0z+ZW1kMVE1IgKr+y4uxZG9YwToBKLH/XN4/6
jWgwB7U8K9URaffAS5JCrQTBdZqHmoyu930oapUpv9x3PzrcJvRZLB/a6vcEK3hN
X/0tVmPbdO35TYHKTY1ZMyU3i0tI/uPFGZvNvshBw+x1bqGGfjClVtdO4wGqsVFB
kfz8oHphpxzeREUBWkjw3IUSse9V2KnMhsArOeAA0m5u7LGKoZVs9E8m66eqrgtJ
IYl0K2bvVyD4dMOXL2g6TKY4LITv3AHlreBrRbJa+I7dLUYwvffbuXvqI+cCfTJ+
SnbnzVEBpLkpIB+3N7BaNZ8On+grsEyNezKR5LZOFQKf9QIw4ziifkJVuH69F/7L
xvMCc2Oyq98ErcNQBXchpuYOhKDskZdPUXJoywJ5G1ZaS+LzxC4ej1ZN+z6ayqKu
YLHKee7Whc3+vAmnDFsWuZ0t6MwfcoF3TYb/Jb1g9RExGT+3oAxCb7ZW/CP6387W
5yGFwcI7wJV+oioKfqbwKqXOELgSbBpQJ1E7uM3WHMb9AW2Vef7hEiG4b7XGRmTT
48TY5s/mS5X9TWf6e0Mb2qmRffT6k6dSLzunhEGCEtt7wx3XqnJOXJOYnU+I9Vp5
uFHiU3neYLBITVQ6QMLG+ntIHfT3nzDTJ2zoy9piM5Q23Y4LizIV5/OLj66yTjOg
qLxOuKkb8AFdZ8wDYr0EXGggzQm+DPurtV62zJogr9xWrs9HHw4I2sLNJWeWx8Lc
F5NQKSneqWzjIukHkhXTbg+5/gdDFgGF8MOLoHMJ/W92zJ26xDtUUpG+Xl3JUqB0
UN1n3X0U+UZHH0Sr+fc8iE+yZBUPfuPqemPTBaVQHUiI44qIr2jM5UaXbg/Ahx7Z
gBe5jrlfhMq4IjLo+4ELdqd5l87s16QnNy4QOAOCn2BbMih1mrSZmJH5+JKLsuzL
N/ctyy85ofmOyXhK3YONglGKAiFlb7fBVYd8cjrujcK3rKWv8tiD6IqbHKvG8bRl
ghV3jfiEsjpPC96ybfLRcV5O9KhMytOdilVGFvmvcznIe89JHXRzWKxRnQRWoeFO
5E7KGf3qG3QkR+ZkYXeLCZ5J2b5zfybpPNEDmsGiu3TWB8MU/4/DMmRlZEU0hUx2
Vo1a63CDA4VpfDUJSZ0MZge8Gs9XpZWt/EAgvnIRGNceFaJL89muoEGnOq558S3+
eyNjCM1vN7Ogfq5MsMfc8n6k0hzWHjrxcgGqHFNm4hc6f40G+ZdK0qPMxqNBHHy3
zPfWtGcCJdR9CFGlNxUNiAu5sSSIYlNqERxE61PtaRs6WwDp66D7x73I5H5hEVg1
e9LjFVtRx8iOlMGCBNBhQsO511VtWvJbBsHA2fWn4CNUHL7tTIXQdG5yQrQpRLx+
xw9QdorWAECqtmpttOqw6klv5+uksYFhOUr8uR7ENdKOWx01tbq72X5IO+yZ3+l5
NCnWOgwdAqNIUnwy251YgrYhkDQMx2x5rTriQHU7Zz6nZIbElafRBIk+JGT3auUQ
g5r47VkAhf7q50FL1T2QDUhYhF1Xgt3S6E7Utvu6fZyMqvQIedDfRTX57AXWw7+x
s3k4DG5+riZ4LOYyHYOxPEqE/K9t63o4OYzkaXm+cfNTm0R9Vv9Rutx6Cn5KYZhF
3qgHpkiLhoBJSPlxIRY8Fu9bNjOTIl168WdFBSZPh1S+eoFhSjp4qNd51fsp5eKV
QUPMrtGdJDemZhY9MoF8TCIb4LNDOKLUusuEP1f7pxwgmhITofyqZ2cMje13A4Bb
LP8P8gzLNBJe60mP+UqxkO/fJe/G2v2IikN+w5OKcjDL0OoBK5acmqkLVpf4hy+A
CmrZORBphJaEDpsPfha4kRUBF6EgbR1Ccuqg3IfqqjEZj4qz5WPYS/sR1Nppyw7M
U/ROJRdV604cQ3WT2kJwqgZXy1hl/6iflsNrUI6LJXg8+pqokomG8nlqK35M9lpl
42UL8Qd9BlI711MhHMnpmMixvJGZ1rCOhnIVED0LVJzVjCc0yCRhC32ViI+9nFZp
arWjmdTTDsOr7NBmCHpYkCpzYndyZfI0Lz88T9JuS9YkzWLmoqO8RygPUxwL+mya
p/UHWDBwKfPGkBILAVZV0iFu18HkS8FUggSdUvWMYgqbCMDF0Qp0uvSV3+rkJsdU
Rm9L152VeIAWj4HG4VS9Oyt+TsXW/LyFhtpnTTcwsAkJ17GVh0y2x4Xvr3TOCBYr
RlGJc7ydAI9Q0U1Y63OV4zQM1PuzRl50kDgVwgHJiPoEstRwEA9y40XxRjAZUIMA
t3xJoT2Lzm7VyJ7P308p3enp6ZFJyk7/c4nJGoFJRyLRSf65z7ZGfKaEgPZPoqsR
ggtget82CouWdX2SmZq9OqpAV6mIKBNIuqCXYLdFYGGtxLoC81ybbDNbXKc/adZY
Zr7EVX9a3b5Ybs5A7NB5iQLQ2DYdJOWKDtZXUSrWyikeQPxNt+85YyFOF7u9bYSa
++vqqUXwAnE1HHWUSvecRPMT255TSMfxm5vLPduqcJHSOnSW/DHAGO8u7ysLdUFg
Sc0Q/CWAGSPHPkdTBeWhFmGdBXn2nfVReY9fv5Z3u3lptV8DNTYrEraLeG+ADkpz
wJvtEKINghd70ByZGS2ePxTOKJVI4XR9CHYxkhb4zD8bR/3IdI1c0TZG9cnXQWgG
TTxHrN8t5Nkla2O4TSy4anDOalHQj1FeD8xFAABHPmSjNKyJmnkO3RMBQcT1AGWU
xQ2L3MbZUdLhpxIG1KzpYJAhCvba54xXcdpWWsU6nqW15SAJXSZ/cJ1rZegpauiC
nuj7DeYI64ErdPkZU8hycyi5WosqLSwr8VklVVuoTL3ycLkB8T89HI6ywwG1LCrr
R2+SvrNP62eXJa8HNbNhEpfeg4wMEsc9RzGzLxV+c3Z9WYEF+n2/cMlOZ9aqtIQ9
CNSX7DgrTXZ3QdmooQncvs/hDTAANHPnmu0KbsjOfluzbBqTRqzIl6ZQjj4yE6En
KefP7nUaIt/mi9Au/XTh3yAo+M7y2PBGDM2sFq9TSIe/WFMPF2xv1EnfPjz8hq/N
BLO2gkdy05Z4RHDbr1aoZ4BbA36b5xxKRcLTQ0i9HIcNFW9+9brcMI4WYZ/uhIfe
GEpnAbZTxVYSgsXISn/wmA/hporHh90mjGMg6i2uw5F/SiZz0e4SvWBTuaW+RxnO
8lU2IjbAbs2cK3e2SuEcXrQliWxPVv2VBd5i9G/jMJt7vB3ReqT9yjDTlGfQXrtW
rrey9ZuV5x5FLKtC+Jcc+8dtvDO3I0rzb/JoQDXbXaCWrw+AoXN901MOfGYgb6E8
3gIyKo/AxUxCPyfcHZaBy38k415oBeow85B0JNyirVlF3VstSEmUhFMFjDCBkzam
ollE4bi2TLCDGRvEQS+kXIBX8nuEMvkbd8N640trw8AVABslNH6P9ODGN/Q0zqG6
9zQEgqenwqUVGmehZZeNArprpJujCginSPvPVm4kzkVDHbOHy9+cWBcqfnYzppzt
9HupDH0qyiSN/Ajo3/YPU/isGf4b6GP5RXlm9sjlpNn7u4y5evu2m4jQvsqSeWKu
VO0gVnXFOt0krZuk3WLdg0C+mmdqRkd6k3vyW86AXPP6dYWVOTJyUzInXqVhOmk/
DnzTbbZqYCULh/4cYASNHXZmYETLl3ZujtuJrGeqovMFWuaIB1bdGl/QItYthakO
g3USc781elYdh9Jx+lp164UxnmpG0k77UEOKWBdkKbb49opDpNsz01RQUHwWcoao
BHsuVE/F6wgg5H7x1m8gp0jYl43h6hPVv0wriTj7usS3PDYG3GR3waM+OhKnv+NG
oiD7mqyP4+Z43rrp5mxKQeg8DVi38bQ9iEk3/wg61tZ1d5+Dfy7qiobJD70S80fM
7Lif0Es7LrE9O+rUxdd07UmH5MPtddFHN5BP6IJCiqbJpuJct33GVVoAfVgnw17m
YtRjr7KTXOn5ZvHV0rqmCY/nosH8arq37pf7kqffi2zmOaWeWeRfLHjdyqR0YrlK
7N1tx0nopT+tX5WfACqRZ7XfA7RbTpL2v1OUpM2djU0RybwN/q/D5Jgpc2+oILhs
pGPpWXZ/KIEk5mmNf5pI6HgurDfLLm0z693jwfTGc9gmF2lWoA3wrRtBmHptAlmI
C9qpO78eUOf90VGlCw9lEpsZZ0O3D4OI2yRMGvpS49bjdUkCJNBUFtUwfqW+WtRV
0EpZ66papIVGePKHEABIZaHJItT22oYla8W1rHNPmZ6S2izGQ+a+qgtDIobdSQgh
6Bc4Jhrji3xSUKvyfllmCqXlBS4Ae0VkLe0A1BaMZ2J6OtooamCmQJDtlbhhRD8f
+4r+ZBH+GIUzvK+MNUBM3tkxc8Ihy6hMZ9U7zehvM57L/x0A3sV7FuQzOcNW11Q5
feCmhIE2UhMLp591QPuxQV2ZzcqM4B/EOnJzwCz+SmLoG7GInTrbeVNdMjc2DmQY
TFwZUxZufHfwbqhNBLraF74KiQOY9f3sQclg0b2raIZuIKJSohC5XQMeBOkXTi/6
Cao1SyKRvgoLNWyHCUMSA9SAnP7sVyVVXDr7bFUBq5N/0OqBOn/Pake3iz3GajOQ
clrjdnoDDHGyV9z3JqwajDai6H6U8VS9vtpEn6Rh8vlq684rrub4ViGNwd6AGNga
mV/y3nCeqaT8I77LFUZzKi1B13ohCydfGblv2/QOt1kUFhMVsHtP6bDi0GRqe7xw
1qQH/xeetNcb220XNEYeLVV3hAvBYnvHdvYBznoN3CqTNX0o+pMzRZthGmy9HQ7f
Eoe1LabpnkCB1Flek7+84bZDC3/oVyVmiRslnKLlP6+r/76dkDFU54gw1yP4/Wqj
cjeVAzKNaDwyK7XsVe30czs0nJ0UnHDwBW5iIMHO2kYUdKgBIaw2OvS3KtnSqbfg
J3wDSAsljIz/CO/UDiAozYIIZ2y0P2IpeXi9m52uihkQrii/u6stfwesZmi9vCMe
71P+RS+z+m/Y8hYMo2fu8msE+3+7HFd25fzZErZaDIOHKXSC3gxeIMUvwrbjhGB7
QtpjgfNgq7Bt6s3cIbrtzxcJ6XKrwMZxlxOReRW1Js2qO/h65k4BfiNTMLsFTjUw
iw5b2/eAivp2i7riv7j9v7mvgj/1HWYNuGGYN2GqecsWDUR8OguoPaxl7Pm8bgqV
uXiMWb+1si/8/DljwMyP17QwJdLbGmiRiY20BBO0ZcH2v3hZhYJ32JmnWQBubU/l
jCNjH8cFwKKVgyBJOgBpeRLNyfu2fmYcDb6Svsp5YJDL4A5vduF4kSujcrZ9HOh7
IeR9VqfY4MxVsSdRFe2aDoyLgwOMB6Nf+N6lngX3+oJNu9KGpzy7tZTcrtQTwwIZ
TrYoecX78eL3F5s0TT/Rj94GpN0oZFuIBf8TroMse2jPWL5r8EjHybZUwFwL1QaM
RzFwL1WnmJ0cUI1YmryoWH0R21rkd1SQniazn469RVZvSZxFrCRLrFxcLgGpbUwQ
t5z4zfmNwAcEhqodc4v2L+zuvMzpCnQFtA6tTNGqvgxCOM8Evv3SCJZ7V9XLw0vD
YTo75WeAMI67N5rLSxBaKrw548DgAkwL3wP2aiK72u987gSnklWwFsnWoy3tJ7/E
cAG7Tz3bNDvM6IRa4KAWAa2l6AMXLwKogNGoacvT4k37rrmP56wGPNHw95R/ahDa
wUF8xoNUKxqk6bw3E8HBflGSdkaZbabkUy9DNZYTqgi78nQO9JmwHu28JBfN6o1z
wjoKHDd//Ui+ab93qni4PC5JQCqFC99psilsNm3p5DLQl9Ryuc/1pqNr4xyVd+aT
vJcqBr3qJwRYNOsJPRcntqYez9Tgx6GtjwTdO5W8bvmPBacIB1NobnnIxumQI8f+
+Rwo/M0+SLdPJUCKpjtraw4qqUJPvVY6RSs6pii3vHC+xwaPiB7iP+d4NF/fGXdE
yveLIdriDSUoMc48bK6VEpmtyxR8XgX6izVwpc+ity89EiV1du2OzrBW6Lr8Fpis
2YsaksJIyMTj88AaRHOQXBfTMpjd+9TDMKtCTlRUkNrK2KRSRjyYDj+poYpXinBr
L5aA21D+mQWSOh4kNzlblztC1QVIaiP6k6VSuK4mGruNwqyhRy5hbItEvaDJhAIP
Aj0JDra9X4w+MJ/5pOQvVH+EAgmnATS7qpLVhwAWwm+zkZjLkbbEHZ75PCoBydzS
DTWEaQhmwgZ9OoiJWxmsov7yuXx7QU6embrSe3bDw4u9G9SkVngna2v1xjwtxPek
zqY9R/lvhDoKRy6DBHYHHO272jfSXBuFJn71jZitFeqYw4aiW3UZhOX5RDQX+p5L
tOLcYa3L8O+K2TOmz3x2oIC75tKcORRxZitoHUw1KRmCh4jrYyTFRaxrExDc10dM
R1Azxs1gZnf0sWPJNUKUiiD/7NUqXTadc/VnltPgQFC8Qe+7NFYSGsGgiFvNpUwU
kurEajKCBvDCCBgT7xLi5LtGVwaziavuxUDmrWspZGTEz5AsekAEz1BtODjvSKpm
clj1W8XpAGqoYB2IhS76oT3N0UH7AAT3cP7/2RUDdgAfyzgKN8iYKxQpe//YqGHl
XKFnDAXkhOgagpEXiyOPZSarNPwzzPG8L1jezJaWRArBZpGeIkO+uJl/tt2P2Z2O
TRx66GJ0KaIjbv9T3USpB917yJaeRXEEN8ibSpS8bZtybz8u02HsquLMcqXIDbPv
ilaewH/zHThlI4OnBrxMztnKccujKwGyZwe/ds5ZE/3akbbUpc1nOyfeKzTzvi8P
LnNGnRem4j1MERpL1sgACieL5Z/6bJDdBblOqpt5NDotLQ0OrwfA1euZAfkh5gqt
Q4sT1cweoid9cLwSeAXez4kQNymtNWS/yXUb/FfbvMbc17+KuiPGRkcSob4x7+50
Yr6DghfBQXn5lIUYU9rZ6MzwD0rSf/4xqmx3RtD31vIOxrA2Brz/9z3qWIHAvZiA
Bk8CSVO9B4G69h+Pb+Z2C+2RaEXxzJ/r+rPrZmrkY60tnk9w+h2sRSf21ze/+s6N
8Z6qF8XYPFoYzDoiSI9hgSoPaSmGsWaDyGMbM1DYgkb+YVxzK0ATuRFiPVsq76zf
I+/Y/gqnrMz/Lpz0aPe+4/omOJaWlGBlGuniGolDMNKvi9ujGLIflPtaBEqiQRVn
tYZHmPhIqpCH/UstlSkW7CTcZM5qDHFhViYF6YIdH4gcQr16aRQl0JMaFHLfSkJV
tQ8alM/5MNLtCcIbAgJO8mmchwoJ0KD0LvmVKLxD8eWl94nnCM8cmlLqUK18u+II
YvCuWaaKT4rztvoToqfOFFhdK+FXFt2MCD7D2qKevwTGae4GscIf94JlWbpDxXFx
i+eHSoMoUV/9FJfuPJuzrTqAPuuF7bQOgEix67Y3h+Tipp7NQbD7p1ws8g9XSOwF
cwBdP70dKjCjmvTE818mYj7Lvw/cLpS7xH5RibJBTU1gEe20sdAXYSIK6x4yaakv
Tb2x7TI7EgOxdJBb+7pGPFye55EzeUaT+RJCLiAIgw8gXLUm+y5SDir1iODBXGlz
pZ7VR2ODUTTu/UBm75bVzI4ieUfMoBq9WVWHBYhCCYolZk/F6MvW7IYMkk1PY4lx
CyrFfIR7M51+AewpEYrsPfTzBxm43i5f+yiDqbQgos6ZhBSDWgQSVZQBLGliMkBn
prhWc9o5vTlN+W/Vm3l1CJYjwdtSZuPx5vJ7CIoew86Jp74hV3erVTNRo6zsPSCB
lGJk9qsYR5vS9nuYQOY0r96zUsEFXyFnwnmlK6mXvqNuVYbUVXVL2IySaVqNhrxc
3phFPz3BgO03sHKrD/ne5xYr5fc29OvQGMVeV1J9vbDeXEexfRQ2pF0XoeIVeogp
yu8gD6owRPpqPCJL4vYo1IiHl0zt7H1o7I4KctK2ccj8D1K/RIsfD7d6sCgiHcvP
kQP6WmS4xGFNpIRrkpiFZtkenNmGilQyXhAsDw6PVp9XF6Tb6A01P+hkrFPKYcCj
BidyywmT10y2wzfvct1XjAwleTfizfC/xwRniuXysaIeaOq6CuE/vLvxgud/1n4B
baz9PX90kbQx7p6mLGEoOaTkup9Ix3mZ+M1GAz/OgkWnzemBtmwfVwgLCzPYK7Gu
73tpgIPZTPDfFYozgeWnlzlHpcOxm+udqXyy4JC2LHN7v97dpFALbudObbvqyCoU
EK2/73QWRDRQ5qtMk1qW46DNZ8GxavGaN3bjyIjhmkvKXz/bCJO1JxUMBbZCPXRp
l0Lstfs5TBM0I5VHa6jvWAkNUP9+pD2NbB5X0W+uURNgsQ3Ys+HF7hg8Vnmxtu3h
8QCF527OIn8tEaNd2CuPBI1H9Fn8lGWKsIAYlf9mWoZUuYuyI3LpSwFv/V1QbjJJ
vHVkr0S/ZL5ywZaespWboxA4OP9DiPxzULabVmRZHAz/BHYccJ+htpF+PBR3ZdEn
1CjyxwqyiV1wgh+MH6i6ffVvH3X9lo2nUPwVIONj7GdOZPC26fiaB/7OeezSX6Ke
GYIH5QttHBqaOY2cSmVHenZtDcmGfTZ180m1UhLtUfvVoO8GMBkgx5wzMhFjQjT/
gpOg6ha5zc4lKAMg/vgqMx1ugwtR0+8f4UyQ3MUw+N7jKWE4C6wN5bGYQA1EpZE5
Fa8JxrHoJCU45OyxDDXuJASS9wMXpMEsacMl8SL8jbREcVQneQiB0o5dGkRxg9h0
TxS571Sxhl6z31xzqTm6SoNcqFw6TJoDtWYuEN7Asj/NslkUV+23bJvO+L0tsoU2
6t0orrAsYi6zJ2w+40Ey267Q/wmfb1CEDsWboIKWVY8RSgsxfxrVva7jWp20xTmL
nJ6KsBXumyh2oRHcFCrDFmqgOyskOlChT0Zlbhc5LMXmTca2mlGp8U7sqRv9LBpj
uBwbrXWaRMMrb+9rfgT4x/WN5O+ZnVrLcqhyu4MRQb04Jb//QScA3TESba4n+lXD
mG38NTJ5KeF1MdL33WuyT6Phkq1V8+DxiS4ooDVr0X67YbilBUa39WXvJr8NNd9r
d4wxJZmswVkwKOKqBK1rpWzXdH+kBIW2WDVCpBPAqdt1rvaZ875p+f2hWsqJxQeJ
wTaz5ALXh7y6tjlRQDtdNnp5eaSpETrafkEv5w3jIlcl5+TknSXZgwZ9dtZ/rMKo
UtG69Sp/2JfDYwiIyRuDcCxBkIyIm62Bk4A1W5eOqpWaZOO+FzDT3wz2WLEVCvcX
25vt6Vijgo+ukF6rNQr9UaxR2D3qBHUDlLY5hPSL+jAIS7Rnj2pUe7SqB2JA8lcD
o2Yd3MglsBlAEkTC3gUZNRZjo0nJduF/KoiwB5notV05WJuzI+ETUrZsLIHsKiap
tLTBOw5P3TIprX9jR0KwkeTf50axh8VOSYli12Z8zGlBZ4kZG4m/Zggyt/SGPpcY
DqpvY3515y0EjXDTtSNTULak7fzSSwpFoVnxl6vuqX8sroiwdgK6lglMDHae7gq7
xe8hM8Ova0aN77x9n589uiX3SmmmgMYRN2sydRER2CY5NfGnXzMuEBGmfhDkacgz
LleJZgeBwXXqgSb8UnNW3bcOD+jA9ffVppJd4HHLkrg7uONlDzphDaFboa+aESQa
7F35ubAp7bTfEYY6NfD0GIa/e5pBtI5DrrZiPJbzyF8xiNWkR+Mhs4GdPdzV3naC
bBK02scKHyy+5F2Dvh4P400zrZrVvxSvzdz06QsnHgsulOr3P+QODKzj4It6lNaG
1t7XN6Xc8+S5lnGbXJ59RnfEy1OMunaxDx0BK8fwULv2L7eoaxMy+737Nu8i+Z4K
XcSgATeAk9xuaT+pAP3NGC5Jl1lP2U5/Lx/oNyTlkWEV3MyJPChmLn2Pa/3CJJKz
V5aijqT+kUwSqp9ZdwjoY+u1KGdSdc+T1UJ/OMe0W5wahQ+H9rT1/wLgtov32zBP
4lCL621ZdGCnUnnGAdf+in1PpSiW8gCilGpzn0UAPhcJ6+7l2Gu9BQ9LV+m9VZI1
fozqOeJlHSm7KARxuv0tWuRb96scuih0bU2XKOkfe+FTvs8CcyaUSF2KD4eSUVVA
xgYUoegNpPQV+k7YfD+mDep7gTy1FOO3aOqXQvIUuxNkY/vZiBMpaqkyeMPoxosA
AnLLvo7bX2sqPBujn3YRdcqAuF4YsZvh41QzbtvgAEhK99WwKjwtQZbCFLjuB5jF
FZ/6c7ICyQ49hXizKlPRjVrIRaNIt1ZwEo4Dlp0O1QxgSPoAzLWsQ4aKWgVR9cF8
IrStRrIXXxQ7mhfsL4M78LLcpcF+Otn/G5u0B9IqDlEXix7tRROpEjFwNFu7UXwe
eSDczyT0ErxmdLHIHy9VpWpG8QEylrO8mRugdc+l/GxIgKlpdIged9j/D2LtJeXm
LBJXO0xZWstbUHMhDnHUzpA0o3baXaSe63uiIpvme5fE+osGfJnPxmLr+P1bOSyK
4FWLxnIpz8CVTRbbtpfzHN6yQy+6hzP0dFcl8Wbl8FWxfetkPrj6McF83yoGqrpr
kweyoIGnoekYzBeRMtBdMf+j6rioIHqo1jlh/xHCCLSRUSqKr0KNcDxe9SruFgCS
EI5nCekV4JGKrdbaXxR/ZSxlJg2uf3sxL/EzDY8EA2wQtpENyZUE7Dke45keAyBl
dRGi9O7FH941QnouKSYVoHKb/03D9Nurju9icrpzeH7ALMPbH72HJnl+cO2Rhj/f
Lr1yrWPyswBkQjnNAkEkEAMPgIpOLV9zRrRJIm4keIWvnXiBI0c1mWpCS3hfSD/1
Pt6PyqdpH8KyzdBs3zdftYtwdHICih457uVZUd/7EaYudXmxnhKEtW/rE79Yfd/d
A7F/DCgtdJx2zUmTIWY2SwyK/ruB7JTul7rzfPQFNY+93WSFMIXYSvdgYpUc2nlF
CcqPf06za07hgD1M4m5e+IvW7tTmw27TxMPCpwEUbD0A1NFnHLXxmTUsYTbN0HjR
W1I8HxnHKZC/Fme2f3BhK9jtfyWKHU6yblRho5uROg2Z2ng2jYcn87LnyO/ishuY
01Y1hw1NLv3ERtUhN+Aj+YDVm5vRMiENMkm1qIwX80oK5GfsI8J5oGddecTWwySc
cYuLL9fptw3UOKAmlk+H2VegRWsC/lW06bFKXxvZoFarT5KWsWctE8ra7GPOoBt6
ETTrQ0F9n2xFm6TY310udLT/osCPAPwIXUu71C1b905zi9k5JFcwFAUMIAOGELJ5
5X7l8ZJ3xbjUDToHG8cCHp2CWCRyNvZtJhZpPpwDzmEVSla8AwcjMFz5F2U6hHS9
mQY53XsXrmiXldIJKISmunpMrdbid6ME6W+VCptzeylm6ZFAJWIz+j+VFftiKtkW
JZypK/o2W6sCC5F3StPvKlGZE58L4kvt9jzfGIavfLtd6CBz7T5R+dzVz0X+8vzw
1se8Nsv9J7DAT2GPwOUmyQ/Gk2Rl1Q+lrM4YDBv+1ZIaxfIxW5MzMqwkjIB2Y6sm
RyP21dc3dhjsfV0N/IulgCmysW12AMhc29WIlpkzbx2AH/n+i1N7bNOX14vK0K8p
B4RyKknqJuwZEDUlBP7e8CkNGcx+svbNjg7EHkq6bcCuGVsVRi1eDGRFxbDmBKjK
pn3KFjNuDpUIGpOFk7EmvK3kmoDtSZ+/blfDtA8Rj7PuV9pn6cgiy2usceGk81Fr
TjOHAFqhFN1bIzegXHApy7oPLeaD9GGLfn6yTvzKdtQmp5Pr1L2StAeKzFIX+jYj
8wOTBW4FrqVqBEaW6bUaGctO12swQOfeEvYxSHEiS+WdZ+SPk6OtTelfjtot46aY
SRBItS8UbvtJbaO7vrlgO9ii7tAA0d/620GA4sHzX63WUDzyF77Jpn56syAd9aTw
UKaPpYS8qNMcUkT0KJmRbpoTYiUkKQ0AduQIXg3d+1l5UP4hmLbSY4D86ADQkpLU
shVk6W1WNeXDJXWNvqVvcXpWCwEwWcdEp7AGp6ttF+zbzxjH1HXQa2dk+YSHYgBt
HFNDCocKAfA54ED+/2ljTkG42RdKTB8QfjX5iGoYnj1ICF0UtgDlMe8Y16DxGZmV
gInhtOrZLgzKtNcxLn2RPPli3lIyewc6S6CjLbDVxYLLg8l9z1Q+Dzc3SyxYS5W4
u01LQZuAdKNqzsKHyVZ+AGPMkpSFOLdGcGkrwc08HXow6IeNw4iimi/up6iLai1L
gcRHOFHKJ9WUsc2PDnvuKm958kEb/YC3hGVgnoFuYx23jlpcJk06+5ZcEo35f1Xe
WT/XdAN7O6Vd3yW6iU/xibEXEa2fISOntErEGqa5Rb3g7uHHx6IRud1A5yvr33yt
sZNxoeDcZxlLEjxT30IuqQITZ6Hlmgg26bDdy67y4PegkoUgkemxRiFvwMcE0ADc
DNXa+D8eTD0oJZxZ5kp8xlueHL6ZzjxwrDObU2dujprvOlG5kak5SX6hO/VS50uU
JsXiVOUay2Tt5jpXxLGw8VnuB3M4qRfF8aBP7r5kUC1BZEfxu+FG6L7tOak2CQ9H
2V0pQy2mTQZdJBvhsrXh4Agh88Cl8eH7E2pxI8C4caQcHU/NVrezEWoPuZC0T6RV
Y/mQlckuv3ym+HILd1eloU6PsEEzed3WdnvVKDKDOpdAdYynysiYdl5JXQin7zO+
LB2LeAthZAISLioZj6qfszuk3kV39Ik5Io0chxj1721tTGFUWZZKazFeyChotMWt
xqeIaNeJWSw4OPjkil1e0eVs5Tnucq6PNKinNHx4sW22OKoNp68XrwmTyWhNY/0Q
Q8fO43dvYS19g7YCQ3wj66N46mTdw/7eP2U1g7STJaEUg+1QQEksw3bDiHX96RTF
n7URnQ+m2KTzCZid/0a7bqVndou0TV2e25TXkvIjZUXxBoSwjxgi9eqLOEDyxtVV
jBwMTDVufRup1ivEpwaf30AOt8dI2k0CEcY0SUGLkF2rg9L+i5raWJBvIxMiS+Kj
v1tAOe69DD33iW+DFvx0YNsnXUptMY6kxAFPk/mie5biMyFxRfwrsjBABeVLhE+i
AEztIEQB3Fyu1L6no+EkQjnxx1F58CWUSnvEWQXIDEaMQ8D4UCdVgqbbUAjCQm4/
zLAbYUE7zteBmdclRgAFphH32mnXPtthQpQYl5QFbPJ0V//BZr5bAyZ1dC9wJSkl
QIgOZxmpo3DfJX80qmKCmOEjRDf75jDbfuRqLiGeHRHzLaJqKUtUg2StWLm7qnCU
4YiMs1fazRT9cNfFk3Trz84vcQrtH6Njqbbfyc5i1efGlW1rgl9QuhZ4hqME7kZK
rHluTCo8PzQ0qJz1ddyXhARIiQx3mkV+65K/KFYA9Y9FH1UE6cm6Mt0KxiKsTRDu
AQSb08oOA+tBymU0KVuVB6VV59jY9Ft6jbMtNON+VE4M9VWTje5FbOtsd8iJGO2n
E4tXqYiNNR9ph13GWwwSpkjYB5H2JoQxCN8KTGnJaDxCp8P1LAswjgbGRg5ppta4
mMm2uCEVwHmw2BR44x2jHh4X0YbrTl1zKcez2SlYb6MvrdTEXMRBSRYzCo1FROz8
zgR5qhY6dnYbt+ajjS8wHFTEDPiWXawfPtV2idzNBmKIOiLpoLmeFskq1Q9/rr8m
d0yLHy0RGCKY2nCaAmOsmXrKqD2iTUAOe6QF7G01WxV385nRXw7WOaNtN4b63dSb
vvsp3WD1lXvOByYEkKWuUrdkwxeRdoTO29sOwsGN6cERgvgvSyZ8wxOzzUgmjlBq
VtwWEksUAod+gJ8sE9zbMW2GTEfqZFwkKxueRrv8PE3NZep3S2/W4GzmM+gwd74F
x25D5jSgBhOGrAsDcgYwzdgeQ6s8OJbCo1t4VevwALplO0o4XFhaOgdi1fGrxvk/
gtXfMg27WGTZQ8pqmLE+EbQMZFwWduoQv6OArIAVmReBk+IjF47QrwN8AoFUYXXk
54KR+GiwUityQ/Hsm0/PwSIq9RwyMGzQ1ctYGNS8AObMHFsFh7Cbcnu+s/3wV6K1
1ssxkqmMAcc+s2YB2dmWz9mC6qXveiGsXHV1M2TXZmy98isvJQj+2bdTYn0WUz3V
GsA7927fs2o9tPp08SZzXzZIkeLxpRlNFwBTh/GTvn1hBZXuVLzl+z2JRmqaCw3P
FntUT34ZlaQA+p62sNdOU+iPVx3qsD2mVi6nhn88msnHpYL0eciTxT/zSqE/MuYP
U/McTbybBMoehrVJyRqkhijZEjCKHqR/tOuxW1lUIv/XqUm/BLoGG8TbMFLm6KAk
Ikctp7TnGfokUfOD4ypZBTGqlPwRACx/82+pSGCuQC8HfMoY+4UySQJDLMcNJT0c
rsGSWiDTPTvTbHRutuM9W0+NULrMqzI+m1cXIqAbeIR1oDkKW3p3NYlCnMtUkR1E
6LSiq3UMCmbVxhHDagDkgNDkKv5q3oGR7ia8wGz4LtJaDruKh2YEigG7lcX3CgPD
43gazgtWCDMuWrVnGdYh0k+JmRGTgWgdfMg/UbFUDBmirhByUaLNktdsDjTQ4nfX
4hH9VLaUN2jS1urf1WrnxaSQxaxZnvEtkDdVBBfXsMBD69RKCfwmFhyKk2zygHI7
8a9JVa+mM/VPTH1OCgiecJbWrcT/Vg913yuDm9oETsPEkmdeImDPv2dYqvALo25M
tFroNIsNAUOtk95gmvxpJTqPGkYj5EEbXerfRJUZ2C+UWUgpXUkzFRZm+qlG/wTb
0fwasUGIkNMko0kKkIz6AxZ36SG/YPt8x2luvWUv/p6BeeExSKpoo4CF9cBO827N
NgMluYenuEzR8IseMsfjTkEzCdw5aNN4ZwRWPrSoGRyYEFoAxGkyisKZns7kAruM
x4pidp2BdmX14gzZGtwDhWCHGD99eZum9AECWVlWJlirW7anGNtkmhwOAK60lsHL
Db/UymjcrOmteNO5r8dz8Ihe3bVNrFu8pmKXU8b9VqSxJliZ7BeZP76yzZOehVSJ
yvoZHUU2Yflz9/uofpbCcVWbSKihiAR/fSYSChzMlyb2MPz3i/kn3Lkygacf1WwD
cNKiytrOjCBvar1aG6RIQRX9G5MetvMjpxlrYOxtCTSJC5k4/w06QIdAqusuXkUD
giAi/XUnOHxJF//TnmgqPFWXuX2wwZR8R8bpdmoedEwZ6yZA78/SVUGAbbMFfci5
OcJjqVd8q0aZYfeqzmZZK3PHxJzShTzvHhb/XJ9QCBiHsadFz0Kxn/co9NGqaMFC
c7NT78CPrYXzWMemw1pguPoF8GWEci5A7+F/Gg/lsSwn6pLgCrUD1olXlCC6T3L1
2IOR1h9WejPqqa89ugerUGwcdUOMc4yAWsU1XMQzZIKSUqv4YWqSHW+ccTgt5FOG
s6TEjoaCoyn9oDt6yy+15BuxEZbgdAsu+XOT9OCu3OeYYJ/2fAY8dT0L36VxjO7t
6nXUS2cXE/lGdlp4wV+JJ90mDQ0zDNHrApSsUCRh6GHA+ZcV7Y8uv0Urb8nqOY9k
KGTrNdskEkO5fJSbo/uBliKh5dHxdX8zUEJmqKM6lc6WVikKjenN7nkUsh4jSyjE
bw8SlJHpFjJe/YDUhe/0erqICujimyZQ3hYaQl5czqXp3z9pGFXtuwItToaTdbuX
essFWxL4nm2ls7sGpPKN3F2J8vbLhvL7r8xg1Zx5VB8ot3OS8isCYuViVXZYyn80
ot//7cljHZw+ic9G0uNSsY0jdqs/MLB8Ij6EY+/le49PWIUcKknBjeCzbbAAUu30
xqHaXl9B+EkvXn5tagCp/V0objjOpncaqvqFGzk0w1z9aY9pN3DY1uTYxkqF/AK2
KdtMIh3/UbFwnAn07VfAuBRp20hxyn03HL3FZrvkGd35Jo0iOvJrqlAGzQHT+IrW
bzp56D+Au9qr70PfKpSWYMnL8NZJpFE5eFcxyEck3OZjk9n8FL/ekzs5BxIRUNfu
8O1K/uN2Gs2cXs/uH5CQv2E7BRuMaJupUklWtb+A6bo5R+UeW28t5utngAFVqDuL
sYSHf6pyJM1a5Q75mighn07JxlTj+I1Pv1tzs2CJHnvL4gNJ0qPlhGmC0ry6h67z
qYl7YKPho7/pyNyERAOpD6fnSuuHjF55Vddrl6GCDl29kzyX3dF1oJFvqeRtTp7i
isdXaj6879NtiK40HL1BhEEhui7p1ZSSoR1M8HaT/X8WLVxqAI6+yyikgmZnn3+H
VbbIwFBkHJG2tFhUbUCFNJq9U54GYChnkeSJX2PVsUDLO8bbAvJWNtSeXvQZWqGu
RVn+fpMEgjdnnpxBvBDJLdbPmZNBS7uBlpVPuK2lbrKNISINxMCDK7BuLb5iQ8Se
b9Lg5BMVB6BQLKpL5BASCx6TJl3CNptUp85oEgOjSi00t8YltiS0qraizjHhJvW3
9ChM0YSedpQbIAOZrjmBhRQB2luOED4Pm8VQnmtfmxeahbyDED1nzWnzb56KVQgU
hdsY64hjRew2esvrUQkrZ9XURSXUuMz1DV86fbumEqCy4jW8Dg38m/0AZOMTjp6P
RTWjKwj4DtFbOTQRW4IOyxS4v8NA2N7QsKtS9PLLoePMfSbipuzourQhQVOmmwGW
HkvfqTF+oqz9u36VOF/MGOTXmlPXtg7p9twiccQOj89eOqzjLwpUMapyEwgnS3jS
dncsjsVJzcFzouzWNTJeKE56XygpURrUfsFh2ED0dFGHM7+z14xGgqWPAYy+CdsV
1zhr5u++w0T0BrgXBimWxTr3dbS0/G0Q+iG/11jWYkAV7Ymg3ZmDQHqH70S9bWCO
g1p0gaR950px/2H4A7qhyQIt3/i8vuMUyk/YXq6kmAhk6vi1aklkakvsc26gG5MH
Djfei+Ex3kp8RUaex1/0dkK4iXkN4eg5IBKLnavqoAoHmQUFNj4w3B13E6xfCRXe
YtFTvATrZ2pxPZxaV+3lZpI2pAxwEsOwiOFVgKBxg9QH8Daq+c+BU+SdsJHwA01G
f5gqVhLNkRV7zn5v9BIyUEiTBaLCArMjsZvD/OshxjJ1MgXpGn7d5N7lnz37QTWN
bqUrcOgaiF1fKj5I1t1pVKJ+U5/pazdAk5zWGXZtQgregpb2m7bN8nIXFavGhUeh
7dCsq/tmK8nXPOCC/zoG5J58orBwMWc3OvhRheMgYRSpf7uoFnT4pQKDFjfkF4qk
IJyEjGU7F6LOfgvJY2R8YLNM9/PYXBG9ggTIihLTAjpkVkfZesM8XPR7D0u96sOm
PuNlektkNZ/TkqGYjtzY9G30I9B4qqvWusfEWBicFuEEuT9bCfxemAmJgguXbjIU
7PM0O18NMp6W6KYc96hm9A1DZGdtQ3Oh9s7ZDAmPB2Yd72X4EMOpQJwPR4pNYCgr
KVnVrjIyC8c6hr8tmd0MnqQf+pRWLFypN2JMl8DSBtSqvFJIDJul52r9fHF4t05P
11OLYisj2djQbEIJINwF5fKI7vA84+J3lyjqgaLhuEdsvPKBuoYpJbsP7eBIgHqQ
cNnrBZSGD1UOqo+IM8760VoQAV1AEDGENGh5GqDuTIqChHsYr67uavpAIVeXZuZs
M+IrQThm0bqJne+sAJybWTvqfPUG9RKlZ+pIkVSW4Dd0QnWzKG7ak8m3SkHLuz1T
3qFS8rJZcUkSzE42jvQMhEA7axGT+I4B+1v9WLwoI/LKp2Jij04l41x1psqbVykz
QnzYGUNk4fd0gwAa4npqGiTXlpoYx4QTHmnE2LWYFeBcZLlukyVQvn1L0cbqbxfz
8mQ7uB9wgGci5Id6MGRpInzgIMIpBRNhDLPqoU/5hoc7SjYD78zrACNPOUmEOMlS
OxdFJ/0/wBceVZcDYgL/URpeDhqUL6q0bZ8nt4DgmbdHlrp/OmrKYKG70cY9jgt3
HNETmNXtWnedJjjCRgB0HwV5Ng8tMhGTETx1MVaQZgSoTgvBiY7naowKZt9R3PK2
lmrG6dnqoWO2GGmtwW5S06S7/VTaNaJ2608+tlE1lrgvUFykGTdbBx62wuKPT4Ab
NuvQt3eVXH5MZShFj1TR4dJTQL8BaFxNcINeAknAOQF6k6vy/asFluopTB66P4wX
UlSPTA+1O1+FLhSuuCP/4O4dmUCoXo0q7paV5Rx0H4KXOuD0VVf9YvRvmMAMuPlg
fXWmreyfuG30n/3QSJYeI3LOHADVuBoBvaWPnxL1+itgxHDdi3p2HAbXTg3+TjSJ
76bee2BuJEebNOwfhzbhbGZGw95n2kdRY9EkV8DQMFCbADpYjHO/zeEDTQtN88ml
YtEK1Su2OIgT5lOPnqA1rtmjb+p5MnqMj+iR4cyN5jJuWDFnzlh/n8E3n39du4hp
0v1VbH5K1agCo5KYWfN059iXxIK7cekCQ4yA448koMlVtJLGqlt+OcU+hMa2D7Nk
o29si2h+fgMBSEyLMtEytL6ofMCqlIPRya6g7+wWmBZlErJb2353MSKgFzRfEt4T
vCPA2aVdiU3iHHz3KcO2K+zeNrTcfiZQy2QS+HdG1WpZckpSQK7jS8NCT79JdIed
6sMK0b0wq1q9I7axU/uuJELRV0htqmLfqtuf89yKpvSo5bSctcuezXv6Mc9cjQTV
8v1oyDKjd+edi114BxsyRBYFZK9yFf40a5NwagfjQp6Gf1MHzu+2QLCsV0iAadWr
68u4qAn55TwfFYsRJOBju8Jy8Gbf2pEFuWKH4fW0G0cqNv4zteGCgxju7ajvzm0Y
hs1qNsc/x/uhKW3EzMQpzRkKrLUBdHtVbG6/T2keNo8Jifm9a3nzm+k4MDSqvQ1d
GKZd1T5sZzqbHvbAJYohbkFMfBYOmSxPklIMkp4wnJgWuKSGP7QRR/VG0oVxYoQH
QZ6ItHzv5ii0Sujsn5+sUhFA7l3mi/mNC7CovoJHvPupjgmsWnEBQ6kifqgSqWbm
Cfud/DBqjvsdlQmHUAWgRgm+5WsDpPYTG+VJWIhvpy43ZcLEoEys+lNOwdfK12fr
m6IFqPgvsftOYyEWtNV8trvOPaqLHFTrzDyAfxYuB/EzXF/9efPDfcr9j/Q1oBQl
hoEk94oEbY2WtmyrFWwSby5KeNZoV2RnT6EDIDbe80PLML4z7BqUcMdkYcQBZroZ
QFedXNoRcpyAl/PJ1qPHFo20Q0oPdtMjgK9/QacRBc993Bqk+GleUDdjoqxSOcMo
iRkvkFFkhEQSo2Jn/hHKED9fn+VZdfZbKDp7SwoVh2a1JegtQF7T1uraWy1Tvpnk
hgesr4kz/3iGZbNotYNN0QhOdj4yp34/rm82NblfIIGl8UHUqbyNQCG8czhxNo2i
2UQP/+A43XvqFYR9Jic/MGH21Cz5XAf/zbhYaAlwQ6wkyZmOUCxl+vp6eD80jhNR
R+FCD6ZFcKwPHNK0FeHuXuykfXntd101HLErrVMt61CZIc1mLtmwEyA5ubrKb0T0
BtD0Yorz7R4bjhFogh3/XICZHGDIc6w3I1SHYnlMfNxQmPqjpCrFnKdAj4/IC/4q
9UcVKl9jnKchFY5LnPIyfhnWHi2jr63SZ2Pa+ODj39p0US76vehJFmrN+TE1tsTw
8HiGG+4hmkubBsl0rovUQBtOddyzSXzI6oVlmDlE9NgwsZByBqnwsHgCeR6ZxO84
LwIY32jEl68+S5/K8C4vFQqj7LSwu2G/bilDylvD+wosR/x6Xn4I1J2VL2GXWHej
5dGeyhHllMM74lcOxDaZ5hFe5uKAuNAxxgf+gK4cFU/1RDIXWKh9RLkULJYkXaxY
kQ8MzU5xS5goV2+rOw2lsogmjlu+lZ/63Ujl8WJSF5v4bbf0svuSqh7HYdF7irtg
KtRmX9yKpCpahIIZ4SYkRlTkBhc7AThCsCgoHytQdxbCpRraMzpACCPEEKZYNaCa
cPg8XSvdfv+P8PqXBJjyFRqDmunzfz90WzROMQvFuAV1DVOZh0gMxET13idCZW+n
LIpD1bDvxeqnsJnTlUgxveh1q4FAH3Kf2wV9Ek5xX+jEYjBR3WVT2WWpOjTzFthY
Kvbg4NO7tagSToidVZ6pOVLfymECODBbP3HDxfU4bBAgUJICZavxeh0ecCeYrJbp
IWO4ThubzBAKOpjujHPQk+0gAfMD7nMbl87zhtn/s/riaRvYy4rJHIpUOko6RgTk
kOeNdiAhqLpiE52rii1dYeQ3TdJlnnZpdEjw+AOYu7XFUmP0G/K0rXKTDx6B8aeE
gjw7nr/StKb50fv4wQvMXrz6VHYttZuNSdvhaPV3DS+9BwYe22wPI3v9o5lcgm1N
v6L/IULYNE/Glvnloz/QowEe51yxeY/OPaNtb3tUpNZ4Nz/bq6rXL23tPLpApkmi
TVzFk2xvzp+BdEp2mKf/dINlKVtkkeh5wb3sydeev5YHOvevyQXO1UHIRfD2w9LX
QFM1XA03Jev1r1fOF8JaZe8xrYPxCoikLnqMhXtH8LPIC/goy7SnZ1uZQBwipkth
2zP/o1KOG42eBoc7pyix9Iof+XNzJG2S5YhL1QLb6yxfAyKWTMyJNZ//9zTa3ML0
VhbpRASqmbVPglxX+s7fYj3i+1H31aC/U/mC59g3zCyVIsQosPKZdmSVDOx8AptE
+YX5iIjThxvzUp//n2ss932c/CHYj/oUIuT2KBRlBqJmqNvRKxjo+uGV/vNsJ9G+
UYl8oZL9fnkvzX6vLlWuAPDhuN9n3VuB+YAfLsfbsYl/5pGRb3PGWA8kIqWrfYiy
GSQj7/4bgkYaEBqFCQyp3QMBhRZz4y+WNafmSjf8Df2xMzhIG8lVNhdRGWH1dBtm
bZcfudgiu1Gbch8qGmB46k588m4XUN/Xkg4pOHm9a1ZVn0ru/QcuNvNzPAobuLDo
5dTVh1PL7jgL9SkmNE5qaVUQlasrk5V25sj75Zxr6JZZD0cg4Hy5Dv3v0Xbutun2
xGeBD33QslL+3Ahenv7FGWgyA1SHQ8fvhhxnh4bI2XDP1IxmqXuM+cxQqiC8CBYE
lHc+nUBOxvM6A/xnLrUgH9WW+zBYQxbmYW3I5sTuXpgL5GkDC76y2qsRdXISO0/m
Jut8hHp5MjzraDBsn1jA6MG+F6dzGfrxygwtmYj22AH+BABr7+UCss6icLfj6Pu5
s8iTZC5Shr4c8SiWTlsASqSG59ZifqKafc74EU0DiB4BqPWCp/dXSQmmipt4onCR
TkbPt6VJeNXgxyimw+Cf4jlwtrlHsCjJa5qIxKourk6jod9d789RMlSOXvpiu38n
YQ2FYPSERzS+90ItJD9xTmfjUiF4x5yvT7AoCzYHboPqlJ4knVhtvY2qQZnxtF/h
Qkg4aC+ngpHo86eVGXTaHvhky6pMp+gIYgmfpbuwc1bfhA0Vrf7PwR+UQ6PvoruX
2KE2L+PluGSsPEAp/6EX/n/QQv0Y9b1ZbbDet0utW1jWI7AGTQKKqF6CWrPYZ1qf
W9ZbbMtsEuMyYdMVR2eXfxvItHNlIIbGJTGQXU+nfdGz1qvLJ4N1iDBtmsKm1DBW
aIrpel/Ts2jQj9vr1ayk2wpKB+M7aBdRDv6qXx8tmAvkxJccAvZyc1j6IQ/Fvje9
NwP02H1Xy4HNrj7r6T0qX2vUHsRKX3GUUH2UsKPTCRrAKDaMCvCznXcU7sf4kDpj
UVngIG6BEHFdH61OzsdGMsNHqE6OgjpSHiaCR+4B4fd8pYYau5NHMq4aWZTBuNo7
oAt8j5oOcRemIY82K8bFfjMtaIv+Jx8iZC1pFT4UgfTS717bJ2ey+RErwk4m1ybS
/bCJLPtrGcnGX4666tJiLDqf8A08hs1KpoLXswOmv6bCJkB2tuWrnm4eGVzViEtZ
NgQLoHQKmL18p6qp1x+ErKM25CcM/5Do9fN4vfZqr5i/8BeRdz9IF7tQQkKXTbCK
NRbM1qIM8wiWlLsAvQbAI/bwu+PPAv0BSD+WcYArht+xqA7LPFN17u+dOxb1FWeG
Q55NRQTLLm5RT0OH9Uwdwj3e7htsJugfU4ddBBBf8JHab/sGOlFaBK69Lg1G7m3F
5g/K9TPHd4GTiazHEgnPcEZV/ptMUPCupRKboXBZtkRlj9DfzQs6yHJPvkmbMwpp
vQAwJSTD6igVTjyEfnowoxBbxs8kCIw89nArFZorNQcjeyNhd662hYd73EmXu7Vi
FngwLG17YsT1TQuNlBWuzo3h9FLJzwVdgVg3tnGuXtLEjnZp+rurwlIi0U3az3dr
7DxhNb5Nigwu8W2xp37ElL3vsSzW811UQZIAPQgR9fkSaVp3eY+tv0zhbOqmrTVS
J8kEGyv20FyMD/OnCKsoxTOeVDo2OYpDk2CuCvHtlyTHw5XH5pVAKAdITiVGlOgp
B4aCY4KvN0HvLUY43143G6A+JDJ+Le9n6qP43ZUpT3xtlrR6eqJlAkOwwNxkDYQS
7v8a5ilxo+IcaK0Y+1KtMZ0CgvSy1JOm8j11lgMs3AKrSgSXB20sQgMBCIKfSqLu
VF3K088wh5I762NPcY5kTy9YIa47Z+a+JbH3cHUfAr9KWhASRkptR1XCp0FqlI8p
wME++diNYThoG/FNtCpCsWXqgA2xItKvzqoCNQUIf1khS2UfqbZX28HOnUkO+5tG
/fMKnBgzvrg8xpJQd5JqpYiNakG6CigPXqkiMsdKBA2t4ybd8vPSPDuEQ/m7ekR9
apBFdHjl/Na8foiiFsVxZOJhjFq04vt2+JySCsxgirzqzFWqtfvINNaEo3PmNtWb
LYXUZWhM8uvvG0oR4KowiEoPBikEEZkxFNUqkHQJHdd1akoTkqsKElFBd2IASVId
UCBtmBFQ3HRJNJp2b0v4ltt9JY/VxRdOxUFT1RvKk1Km9CwaG4tOghT4Wddi/zSC
QUlib181lJYBPajyqjSmAoBf+zLSK99XVD2Lh8RirDrpjGQE6oVI96tl6GJi67XF
glwPUA8K3rBlu414hhDFZpP7SmNiXoSH0xe4QOOT1VhOVOnCEOK1DDhFvyr+xffS
/cjDOqBQ35mewl/umotM/SItFrGAkuWz72T19A2moOi/BpyaMEnyUroQQp/tAfCp
sgx7NhcKxWgAK0RQkQxW1MQKKjpT23xxXe4nVLsaZr3vRSuFZQbtyF5QVuifdKGL
eBpIxWPI5cg9L2hjDeOxpSvc7RAZj937J1N6ipSLSKbJaXiXRlicudII6vce/WI/
23Xof+/gOMYPnaO91hdHGSdNI3XbwLJS0ssh/Jd6VlDumkWx0/rFUMKy8FjuW7Nh
zzwhrd/hBjAVNWxQLbyQLBFfY53CvNye7x0SLtaGpS26tyS7Z92K50OOQkfeaDN0
IiwQy7L2+/wMpBXhdpmrZyy0aDy2TRgPjNSF/qw/X7rKmkBP3m/8O05mN2CgMzCA
lvRhlxUOwm46QekPd+ktgQHHNZ08C7u5nE66ofR0lFRXakzfj8EsaUBRjnZ3sH/u
GZ1aKFm5fxR5LhLz5DKTEELa354upQeUojXlmx/nG3xQ2PsdBmZqk7NExfErHLz1
lfHcKMmLJ2wg9V7r7bumehMXu4xL5CAKyYEWZtJfBCKi3/6WKx93QCBnN2O16Cll
yfF8hKbsZm77oimHCw7jlY1mJAiEoL1zEqZIlMnUQJYteeeidcZ3/Pqgf5UOCHId
e8rXkkDafIADiHB+3rgSeDve8KXpgjD/U/t36RIwaO5LPDw/UUqvQpYLAiOohHUF
MIFVjC+SL344H1MaowL3lQSk0U7D522HEeJxL4eZgbnKmW2cTIYyUIHBT4Hmv47r
P5mLrXB5dZgDhTy9CYwrCA2vOeYqgn4Lu3I71KvrFw7AeF+UKPJ7jEw9iCtz//dm
92vbte4wu8lKOwQkkTV+eKEO5B0hbGHFbF28AoxZtKk2tt99ZRNgnR3M9Nh9zlAV
PtBn6siyZDlTbob2AuMTO79FL3Xa2rRDsiwH7bN8dPGyvIQ9NNaICTW0SoUTjhX+
gamZutLDuy/1E7gW3ggLVQ7f+pdR0wGbG7qDkF/dreRlWiGRTlJi4Foo8y+H31j7
ipKNoeaqZsVwtG3Gn4YLkvROZLQ39kmNuNnrWeJyRQD2Zip5tFbwgCIcz3gCdcny
O7aABFwHWcpvE4kIyY1yzvpFj014BZ0LP1AZl5cj2syKZKdbnpkOcwcbgcv9xcVH
SaDojwhJqoFmkWW9uImNqbdqeuI3AMhZHQeAaU1damVjtYXCt6Gx4LCgUwXXR7Hk
ztGHtuqrBWBQkWXYPKAIAs7nGhn0E2ICiFQgV1Lxxt7gSQQ6TNbK1Nqrctgj6kfm
S7F1FWR4CrRsqa0WMx+QV2WiL5BaFN88P/eDkQlLlRSlAMdaO9XMKrtnLqNYyIqQ
mytrULAY2iI1AXHUofWkLmNBqp7s+AFla2fzsUTsl90Uw2QGcAqKT+iOJiD9rcNc
LKmHQ/eUBVI5DMHSObWz/G6MxABmiFb4QU/V1W/zt9xfwLhXuAlSBItEOoGfGGJm
oS7FZraS5YQUo35GSwNCF05o3UqmpTz1rem3Xqp9xqglASz/fpPwDk4sSio4EN3c
GJQs7hXZ0MRpDukgmP7PJJpl0/qRvuZIfKMD6CgILGncU3Uewax079rbKfqND+B3
nUO7p+o5oJh3M4kvIZ2lfxeXf8uf0EIqk5+cQww6EL70mOMPG/pUCcYLEz60J2sD
e39jg8tNmD4Wl9IpugCh6uQpW3Fo3+vLbqhE04DCiklecHiN4F6DQYVR1ceBip/2
rwrdNT4lFVmuVpC7H/bKshnedBTBN32MsBsLq2cWWI3IaKzJCuWeBC7oMlOpfJkW
WWxn84vAbuiga7lclCgYBjgO54YhzoT+bjXaeGFVwO3w8UGG7A15iDtK9jknHx7W
d1hF40BGACmX/D/hx2vTUFnM+wuB3KQiwpWD2BP1eYSpdUXAoEYUri0pQxrRd01T
zqMwqO5c/A7ULlOW4wXnpusBzZVcKug3rYyMC1cmOEzYZ0+fX4/+RLqeNgH74DQ4
aHBrl4jund8PVfUMHcYQhAVQzelCetnYIKNz0lXbL8X50jCWWQ/y28cEntcEiEav
aetwP92FZGjs5NYeCB0NlE/Rft3UnLzkFJnxmUhbM1e8UkCtrfpypqupCgT1gQRV
QlxCw++mqotMVyDOPGaoinTCYRJQn3HIH3xBnBRw/3B8j5asEpBj9VvDiiMUyzZh
F0Zy+KDzkQjhY0RnxIqq5oVtpDxfc6ipaMKS621Lrk1536CYXCeZizwzLtRlyMh9
IFt9B1K1kx1nTZNVsc1bBw6J4+gwFX7oumiYkcULkI2C2d2maSYOlXJ9hTZU4m/V
zHjWhw7BAhLXU03w0v1o0hfV1EUQto2yeRbtBSahbCYZniuqxl05E2A8d6RUCgkQ
6ci5nN3BLfJrMDOmnIa9xNpmOgnrgExcoI5RaRvN1EDEIv8g3W1WhUKDTOwzSQty
8EwG7wSmsxYjECN3EpIc6R21PXWD1jP2q4GrjMh7FkpLkRPr5bD15mWYp/IAljuY
IUX6vDBjKQNmX51xgLcBtMJ+/PwA0U6xbiqtsLcInTp12aZHSkzBWRSnaWl2PJxf
ViDzekpmYz4coL7gQlIQ5idi0XZpWy8cJHr6wIiCjv1AJ/kjYoFPJd9j1hI363/W
P5JN3OfX9CmZ3fHPFQHZ3yG0j/2m9Y3dIJuU125IREhtHMqNE2Cw5mwOBaFkVI94
1QkVomcbeSEckz71O2LkYjl2wCYV7kCz4OUgFfPzrnGDVZSkcmHup+NWMJDj5fjO
GMY3Fm4PXmMl//WuOUNFQQMLshqpQkgEiJ8K5MKAKe5LcqzOHNZaa0OAm61xTjkw
I92Osce82m7J/zpCETJm7AE5JavY7C4Hmce/LbFEkUatfPT3I8Fp38D9ym+oDji9
ZLkipNuBVxKSyjAP/5FsUVOwkrAsnK5OFmZ2NWl1tXEouQ23JEKZ6nmBxVeI3LPD
WbK3lKxDdh/00fTMjalREDmkjmGtGBVe6IahGEljuo23dltnShtpAaOfwXB40uWh
KrKCJNSbhTGeN+eGM/KtNzTcAqUfftI6GVeZwqfqT9AwjelVLqSKR7SraEiUcC75
/Lg3q+OjFJAV9+jE8Jf7alTdjT3HfHe2QvTx5TNsZ4QT6i6GKRYPNpZ95pRmT1Tl
5k8QZPX5kWFI+7+n3E8CjuKwSmfh3/ioWokpObpcK3VruFwzIbes1V9AexBx8F7a
w1PUip8Y7Qsrhny7P41rSgm+BKr90taQ9XDzasEEhha8zyUCeWv29XCxneUGDuEO
GtX+qh7xKgrD0QuaJ/T0JVk6anBYm2dR37N5xxbEXaq0l9xtu849Lp7SzvWLO9R+
RPTJuq0LHmhuq26F8sq+fuYRvMO5gKKP47mKBG3yEpxZl4l5QwcTx0J7+BfCDlQM
7Kd8CGB09hIa98JU6UNZ7E+CHBU5//Cx2+qA8+CrxpOLqItzTnU2l6OdvhPXOfEu
bBpeGu0sD5T2rrcU5jks31oDqqAyODzcM4zpdJ92CmeB2qdnp/F9mN24/R9b3cxH
GoKRnfR15D5ErDPR5OwTbJuXYB2RVHBxlpWuLlDOz125+9E0nQ0jaKGJlP681P+y
WtOz1AqrMxf6H0G6nmkE+BrDCFcCToHnaIm0FTQ4FVtVq75N9apI0LUFSojlHlbE
DkGlXWEy5GZLwos80IkORTKdGr8kPoRCIbxkpGdvpmArTS2GZd4sSO4MYFA7pAv1
mTM3Wa/2jRqgBYR/TRZo/q9ep9ucb8cpfWquFkyBND6LcHAqTHo+ORrZCZao1CIw
lw8Rd++fxsJ0NgH/YGtGNVSWzeFSos1c7/L5GZp1s1oJqQ72yWl4IF+IcT5IAd7t
uD490ksvLNfM/Kr14taXS/fSfnauJYzxiGobfJDnB0en2btTehgRY689E7154H/H
1dPqZXUmQO0n7NwCPh6Byjpu3nASoB6stgUNA5T+055Tv56eSVO9PCKRfIPXb4Aq
4CxYQPGu2VW6OXOFnU/az+M7/vE85DPQOxo8tUln1TLRrICdEpM1M1PllhHf885j
ziMasZWgtJXE0wAAGxW++zmaVe349GbljIfSit8AioqUXiIdHOaCm8JqNCISJDCN
+xagyLBwDv+4YEcfHHkJqsxwACoxYhXebpICfHTx1yBwxV7KB6LTVAZjCX670zRP
wH+QNGDZuk6xHbDZq2h7f8g01mS5R6PN8AcWd9ywvstGLUFyAa3MkrrsHWAdoF+3
nXTg/Zn9qOyBoIAX0D+GkeT99sp7Qp+UMz26FCWebeFY+7ggUmL7f6j6cczPJ6dQ
A2VMoDJOCbh91i1sORBq3GLecB3RQbjPHe3lLvdXaU2Wmq3byMAOHaOOxWZIlNVS
4oDN4zNedi6vSwYJDTNsMpInR8xf6YMSZJhmeE2LNs87kVHyCe7W5QTiGjV9aseO
MDGRkV5X5nB+9kZwC8N3FSUgBf9UgjMwRsJtdKg1vVLfx3EHcBd7UMD5dA9KM+AM
q7pn+3w9eqTyhYLlIKGN8Sm776iscChZKXWx2t9HNN84uNRqxoXJ5pvJ0SahgU+j
Cc7D8+vFU+r6FQCNgIWAA2V/oETc5DOHUidbFs/NZjCU13oCtnlBVsReuFQIV133
eptCRRN8yC+R3yMk6Jnb+pzb6hbhCDh5oREP4WwOXFOxen4bRm0B0sPoiwZkHBQG
HmJjBq7Ls1iTM6bl4kFWbscuclmzehLtb48WFFNuM6UR0XRxQwfDMz57jtbFoS+l
xAMV00h2XgUa0K8iIAg2HyMlRhWlE2sTTFi49fe41QLKksFEQkw8IaqgS3xcdVPy
xc5baEqhbGnSCwpl3Vclq+nzYjxlDFzxnnfmV0r+Me/Aco3r2v6H5ELHf1cIBbBq
kTS+r8L6It3o0Em+4h4WmIubT9u6DNQE5/5sblTRbpB1AGKKZm34+xCn5lmFAHAG
1jzOAbgdOD6bWqgxXynFZwRYhPGEyg4+C7tGDtlnWLZ9IKpO58FeOTqsiWR/z7mh
+8WaEyO/g6XrSloMxDkvUIKtG0N4oztKpCqJHnVXHTGuu+oVdGUc7psl9TereU+V
4axxu1tJoNuiKwvH9jZxgw7Ci1Hh3XJWgpcslh7uBjzCJvyw2d6h66i3bu7lYJBm
KwZJKYB8Wbf/WQrzNkmZcfDo6iLyUlsZnr7XRakBYb99xkTheBQMsZBjtPrxGsks
8gREKadRoAV2oDICYCW4aB8ra558R3PL+NRbzf8dZdh6/s1hc1xnVygpIHmcvewH
8+jjHNkmp+g4s4DfGKbtl48cJ5ZIdzX6nlTwC3Wb7GTMx/c5D4alRwLz5UJwzKFB
ii+McVynlnwbaBu6RspvUotKI1sPPfXx8oUaim+OwAU8cHc9yzInwFVDapK1ptNO
dtK4nONOsInR+5tzKHED9gC6HA3FGa+uba+WIae8jF88wOWqbdXInBJP6rc2wIgh
WTr4QolOJEmMKdybR8ztEDN6BZivodwy7t/8EpcpFsfVCrNhIvo9L2AQIojqDsfn
xrTKYaMAzgwnFT9ySZ39z36ZScdSxQgo40gH6R6VKyChflY94to26f8mQWZArQ1K
bFWOqUdByYpnQw6bPa0qnFGH3js5epyW2w1VlONPCN5ilroYBRWaajEdJU9d1AAy
SXC51XNm6hUfXgHKN5LgWH+IcDx0FFW6ULTyDVJYE/Uqru7zUISnCqI5em+dxYor
hMPSw+bzO4p0vT6cGJ6N1p0Jkz+gtfsDh+1PSpO4wwd7oyXl6k3nEfWDG7MX1Apx
pSTR/4DL24PN2yse3T0v+ZgqnNXiRyCwiUqnMI6K2kxdmNb+NaWEEF9xlkL98yKr
e+Nd7mttVQeUp1wxgj/PZFs1Z5c0sSlazIaCJIxAovuYRV6qwBQQqw9McOMqHrXY
frq0L4Zf0aXcBYmKPr6Z95fFT3LUqvs085uNfhCwwIU38renArln0QugTKxn75/M
AkCkj1fjJ26WAfp0HZ9wXp5pGl3uMcEgVZbWdBoZDhOEn3UyOZzdaRH0OxpxwdSr
hjUHEXv0a4+NB3KwUangNXtTVbGg9Zv30v8xdQJzj0cg+JE5NVThbs1UEgypjpXh
ooyagKLfOMHR0ZeIuzlu3FkAzGs9GBqLMEbfG/mnIQdVcCsCvgqfp+5EiX60GPcx
as61Nt+z1iy4AljBmG8B6i/ESx1SXD46+Wv/Krt3ZBOxqz4x+unPlpLsJU2qhIlI
x8pc0MraHmgkawnMKK3d/57nur9iEf204jWAfRcINJB9EGb6nPYZfFKoPFQq+s9k
VtiUlngPMY5VW5ORrJXhv3UTjZLy28ewRF+LerBk5jYv7vLE1TXSoFa/vFEgAXlm
vytt4zJYG0T8w0Lrh0HGHohWlxjdLY63gj40Y7O231BX/vIWyr8eXlRNcaQ3Nq4d
+tffcfPe18j38euVNulJe+NCAsoN5QYwEnQ84Pi4v5ptEnaaIV3zeNNTaMCfm12Q
BSAXgHkT0+Q33g7fkhP3UYDd8UDdCOdpX1vuNPqakjed2moDo3DRgUN5fMRSSTvH
E4F25W1ZabSPG+RGmJyqLgUghjrbWI2gMuIG0WNJ5LTObON3eeILY+SEPf6secBv
+BzR7EmKNVHXM/kHc0cBr98T0GSIUjnp85NxPnCAvsutXuR+ZwA3Uw+on9HwdqQS
GSI3vXcK/yLvqlRzcJJAmm8CIEtqLGV6NRJsDal1Bk2HA9ihLcC/kuyPa3/9Gbkl
VLZC5OaB70XiUXMkdKLZTDIFpFFDdh3HWaJA5SgnOdFdRGR4lPpwnEtPzwTZLpoz
oaxvepfVIwsWoU72sClFJSMVz6m6DSENHskpXV4Ah4oJNCwl5X1ij7i94p7Rs94m
Czay5FOs0begTxNvDpVevOWOlF55RucIezGyFOj+u/k1D0+HpNDohm6bPaUXzvKD
e87UkFytsN/jV88ucWAj57R9Lz5ioJS3JMcrTyB38c7dyX4+KDdPHenCZiBwVgAN
lnH7d111JgtbvLsAu4GPwIPxYPPVQJyfMaN8nSiRgaxSxZYw30Smao3mc5NaMiZQ
Vi+ek8W7JbAplNPKb1EGDkirg19IeelwZD90phtNbaHsFaLYL/hmcZ32iekv5yza
22A0aFVlefEseMh98og4mTtPHnA6UdYQbinkuUW25fQKxXdAnhDExvjj4kLVXPyT
mW+Jb/XKzuicTWbkKll9HW3m/+0O+Q6rn3bXU/Qs5/s2fHqP2UDELGmfBfJvM7vy
xjJdmm/yfw/6hwxHK9ezlSZLQ5+/9fZla9iHAigeLZuvJBSXxx9RXLA36XfTPxA6
P69NkKIxKoGGjmIsbteRxRtIwk9TAhBmtlSY7KVvnXi1BgkiRBah+nCFf1zTYg9H
YVisfltTtzRik5bQGyBthyIoL5jY/+VxA4atlX6PI2DTE40ZmlbowprVguqnrayG
rSV6fgQMNGSBb49kdISDSbZ3ppLlbMqf3najPa9uofF/gS1W/tZ/rOnduucCBdW9
6KDq7fo/aCRBzLAn78iUGrErxJkZPhjeyyJKo5Wtue1oMVGA6zI4jLRPYgPtUmyI
3yWI11VArrijtsp6mTHiY3i+Wf4u77osbf1M+OSnI+sgQeSt/gn+7zftqCW3kyWJ
/418gL2AK1sCr2Rerl4g/eEk117zkVCCTBa1UuwvzQdK7lkIfK+ELeTM38J0SHKW
rLtFqo0X7rpMZAH1gqdD5bl+jFdqMe8xDX6bMa4IAZ0R2Xp8+1RWfBrtvYg6vEfH
Nb5n6MBOgzYhmcPPmvrc1afe6F9G/qyN2r81jmoQm8d0CSHJfBmWkEe9KwHgOBw1
x9+A2k/02WCkmrERxhJE5caTdK7CCQSMWW9AgE3605Pdy0FzzpXC2RCu0aMgRhRc
thqXtcdidy3qsVoX7tPGGH1ZrA2XHooMweJo6z1dyzkMQoBpJRHzCab61MVguNIC
8Kjtj1pSG1z0OUspi1YDghmsbeAoV/XDab5oOKQh2N0mDOrlxx3yq/q22QBMIpj7
fUPHNjXg1UwCiy3T5DdqGe4eI1pms1wkUEGg9/5H8uooBWZiMIjQcgUqJpqxLsZH
Rkfaa2mpBPn6r5T+dQrQfHRgJoiXDZkYlOKDhuHEWazt1X+J4Ww1Ee+o5VY9tuTM
153yYSbjXINOZUgIOhbYBwHRBWoqq8BuwqHYrXslyu68aXCn69Qj1AxPBQngxLiZ
aBnsfNwMG1h0BhSc5eaz0wk3CUBjXIog0n0Lv1+0GbWHH1mATzxPYArxfrY4mwUP
N27U83akUI4uzs1mq8cQWXSUmeFmYyTDrjM+GX+THTAJxOLP0RYquYujT6Psyzp0
FW5IoY+vU9g2NDjzzu1en9AjnN93NWitW1ehIuAoSIk1R710yIoyo0tCWtmmMTGx
00AVNQNBQsrbIcZIOcXKxX0XCRD4OLXLCGOM5ocvNlr09ZKkBs+m7s2R7jEoOU9t
vqfKVwd3fRVxshO8bHUcF4wFrc9Y3lH+opfEiWqmWj9kYJEwK9bWoyP0MIqVyHfd
3aUJSdjTIMzQu+rCsdgQDiHzEhMcug1thCHDyQtkrhlwAnSoZ5yLhYQyvpDlRx/u
ku18T1gBkj1qVRdRP7/gwW2mEdOjlMoVEQ1r7vmM+BpafdaJXjREYu50tfaE3drz
NDx4InLFnx4SCMllWqHvDUeYVkm8/ytTdMtHPwfiBrAUrafANB94RPAeW1H8bUFE
NAOPM8acCAVq5wpZVIhIOxQDVhoLKDb0iPSIigepGxTxKfwl4mPZ+2RQKJ5MC0sy
oxsoR3EPu1z9MtvoMgm2cdYjgES0Qe/4OdfHPVRVPtazorGvqJdJ8ntid8YoRfNl
3hRZBDEBGpXgGWL3v7qfcNlLvAN5ZvBXzU4j+qb8RrKiZ29/2ua3ySZ+SPjzwC2W
BnkP2ga/QqwKh0S8uX5ywRhTB5+SL2QxkEEx1C1giXygHGTKctAoNa9GDGMK3Sg5
1RvtvfpSL0aCjgPeBbfFsspHTTgsni6xbZC5vG1Vnd8FDag+zI1fjbTCq/2jCs1O
8rzUN8bY3sRZnDkIO/gFuYGB/3scC4yPy8gbJJeGwxZNBgMGa8b7yQKTNM9H+NTo
BfC/lY82wxp5Prejw3xAwNssi+5RPLlHN4o6hxyp7mJ8OWWRH9YD9m0b+5mXPwhh
bAareZQ+pbmlbRWoBwSewIj6gNB+QnBASCIjlRx5fXPfdJZLHiNcnLuwNsTDPrQq
jLeC7/1AUi9ZEeqyrdVAxY+afQAoK8X9eUcM71TbwlcBcSq+LonBPYXdVpMraQcR
t1Tui5Mu7FV6OKjmaoHKwy3r22P7x5lUUdv3izdlTqMYdBkG3YAmbRr8eXPDU0Z8
G2rBFsRWxa4j6Ipe89qQC0/s7il2Jv74rx4Bzz0fOFy1CFH2ZxIM59C0kO51Hic8
SFeRzMnz4LjCyPhPMMmnobaCe3eS/aAgoap2U50xf3mTWvwEKtNmiuBSM+MKywwx
6H4VnjhsW3eCTPNRLCPfSlVZAtrphcwgOuNwnjXh+8YYZmCcQSrdOA9Bc1I9lCWc
l+KnSyYABWPfrfny9fYlHCmlASjz/hX3abhKjAOFXGf+HbwrXFnUgjNSch96/e8z
LTXQQZsjxMD8a7yHNKy63O6ONVN/Zb61K67M9hJj+K9O+5bpjrXa2NEcKnk6B0u4
3ID5rPzgOCmvagZAExdhjYu6BeM9yYhm1l4gGaDxfQgrnUolMUInsScNHOuZ1rcG
yRF4zeiw0r990Wttt6+hEFRKL5aY92YyGaFZZJLPGzVqsAmoR8MpbJozMuIzpcf+
DlqYBkZqGX6wBAvIZX9lTgUQ0TTNtxDRjYKe9rFEtRLpYR59myPoyzS8Q/gJSU/0
3fWqDPcNQJbtD1/A95r1JBL2R29Vn0KUwRWHWHHHx08qh2fmPfe64GR+S5LN8X/J
CzYem2LRSNSRNIQ7u2fSw22equZCII49ePdPP2AeSLAZBR1pYW+XAL+naDwAzsGn
IcWoqv8ZoW3xE3tV0a0z6rM5Rfl0F++Q1v9r1hesVHpslvIct7PJ22vc+p1UY1nj
Mg7RSXJ3n8UzS2P5aptAsVUsCbIeQ6gllS0iYLQ1EbajhVBk8uGzPN2uIkYSYEIg
RvEHqASXn9vzczNsvzgpr/c29Caa7rJgFOPc3h/AeAZSpVl7L45xGILuRgM4HD8m
QRdfZVJFmxe1PMDNWZ1vTD8tz7z2JTPaCN6RxUvpcTHd9IJ96JwFOOcrbw/ITGP7
Af4hQXJHe6RaTe04wMQkG/6e2/XKQ3CEhZrKd4aZqfSGoJUD5Xa4qStuU4NkAkNa
ZgQ/6D+g6j4qciWRJDMGsdQE/h3TD06ahVsBOWc+kRijle0Z6N6JtpRLI84cfukm
l6zPbGXUtkm07TnUuo8d9pvSZSEGBqlYcEmviylp7g+xX92yhxaLPkNnnJdVcANn
lMrYYJr9tNt78Phwmt+GZy9IxEfH8BHRAjTuGIbuGKKyGuBrg7gDqc/ngXwLphnt
ZX5EUv3ZTgMn4VNpLJPvPQqROGI8DxnGQvtwhd68YGgxwKBFFAYPVVFJ0tqYpKdL
Hc7m4NiIDMhHyi3fGrDGj2tkPS6NGu7yz06w8qjFR0BPFHgtGGvuEcxBns6CweOF
hVTKZsXP2T5yPA3JZHLIVJpYMD4j9wnIjZoq122ATfVeGU1Lbu895UR7E6Ic7R/v
3MiapUsSPp1ReL2YeS5pFzMZ+BHIuYVHo1k8ygo+fefu13Gf4yfYRBb8lFnGH86V
P4zdUB8IzIFkK+VqdLhjFVUHfWmc+udvZ4HoTwmdlkcoExepBIX5OGBlV10UewDt
xritQ63Uc4REXU+/mjsF83L9ntvGIgmisQHWoLUpaZFDTVyqJtYEZ9Hn4oWBeK1D
VLuQRbnZ/OQ7YOHzerTEEeywcU6mFDUK3/fivCyjeiHJMAsM9OKWvoSCNJd0o8Ub
JtVt2soy8YeEw/AyO2/fads6HkTe30d9uvflWpgJ1GeLlAZsQZ69CLA8R8o+SdOn
W0ICIVc1mOB7o2EM4PBh1XQmFLFtbn15UiKJHCIRQnKYjpcuQcSh9evmuUlfRx6O
PC+r0+CYwkexQT+kxSHAidcK5aT8kDEfRmoT525Jfh0BJ3KtRgTlnkxX6aY0fUrH
CvJe/kT5mrx1K1KHibHVPFEi+fE10xUn564z6eQwOcLB3Y4w6466L35Puwlen+73
GVOpUTKVD3KbPkIlI85D0/kUOHyZty+J0/lyy2jAdA8itAhTMAvAw4BVGv7bFF6V
zIFd906CVHQpMKvfwC28aNOFQfZDFB7Zz8apoJr/tVIUJeDe3KqU7pYuwZnEMdEO
kkdPAIBxv7ViOQYwR/zZpc+s4clQ+pBaeZunpxPbqwP4mIvNqAvKeNXbqgbue0Ne
mDLGgNjblaMSQW9cBFmdUggowre+w6srHM+n43FG2Q9ZGJMlXYsJo0UT4hD4locZ
dCMc5Fg8T2ApHfRRNXbmYaESp18mmnnDLTE1Lu8EJaf4I4a5ZF4iH80i66So9E/W
f/2SnGX8ZuELs2fpqlgPvt9z2BmWYr8u97JebtxJ2RzpGOJYbajI8o15qAmFu6wQ
zgV+a/WMb32VsU0F0H8pBPqq3s6H19Vq0zl51nn/AvWazSzYmpVTny9/idhY4uCg
+PWSuol1Cwuui4oJ9UTg/4RXaRs/nYpU3dj9Tn//VIUCBVweexBUun3ODrp1y0B2
puHtt538o1IL3LPxw3/44P5+7n1vaYWIB+myiUDSGvOE8Ljg/HNfZ11RvwTIP1Bj
O1FDUpRsMx+bxzowowhcZQY8GQRrRRVwpJ+9nVL2u8AhlD7qNeNQPrxw03EGNpTY
HjZDuTBma3+Xl04Ie4bSkFKYH69tM8RzxjwkLjVmgI/+Xcd6S4ZvJ0BbNgmdJdHq
lcRlS5KMhcO4CfsWXNFdbqm4e9x2UXSntNx80gljsppY2juAob4j4Y4CfauKsxCH
RRsKmSnI11AK35stF33K4bIsV9VkfzbQ7FTCdroZZuCyYfLyoauevEMJZIHsNavO
w/7jRut7WPXXm4V2liCr3/ZmrB+yJkIysQUhedt+L22VDFhEZVFnlMy7Q1UO4Hag
BozpBqS3HBEkDkelltDAFXs6oQZoJlD9uMbBSmK57n8riH+1NwIsq3lcth7ZjATc
lfQ1bWlsXE3W1RNejziYAH+JvLR7Il0lX7Qg0JxiLSPQCQpR/nTptG3a+0q61ix8
02vNwcvSqkbq29+zxRdiZItTA/reaikEGXLz69kHlHOhdtg3Jk+iKAWR7yJ7/+bh
CW9k1epv8r13DJpg3OkFsX+QiaZprX6tZKlCR9Hc3PHSme0tmG/Q9MaBKKkaK9fD
QioTR45+HjNESutDH77sXrRRSz0SV5jlPs5T7hm1IDnB6bHTj1+P40VtIH8OVlbc
tx8ETTD3R+rHEl5nIIT8mXhuDUjfLV0w89pFgtzP0ap+jyiAwY0FtadAc27NVQVC
1JZE6OSqZu3sHaBJWTcGYJbP6nayYN1qKcYtWfRCd35aaRy0y/iQuFIhtpuiRVJZ
ailhntpm26DwdPFLgjmfmK9WAy0Op3ocffrQxt8KcSCkZZOyq6aPYD1KNDefj5GH
9wus40O0VZpGt58ZizyPLKUVW63vQQbk1LWHpziGwgqT/tX8PoPu8ysM90+xsQAZ
Fv93Xl+k5l7BJHFo0SX1BdiR8IRBZwbGxAe2PiFpDmhvMaa8hY0EuXK4QY2/yV+5
r1eh+A/B2m65LB/45E7zbsyd8lgC+WmQdP/tXlo4p7GP8Gw0d50g7+pTjMkkL0oO
kkG3gEQv9v7eCj7cha3QO/B8VrkmANdyRWhgCmF+uwYek6EzOC2i3pzotKVThI/i
vuDdyJnpdF37oI3hOSQunl8Xc9GqvaO7IFpvfBN5v8267TC2iLhMJnv4o4FqAv9I
NrKFm1fjm2OyQ87esVNIK56NBCZ4D6k9Am3qSamhoE54TytT+nYB25tsNc2+bhLX
JZLFtBm+fjzhJuW0wP3ZRgJqnF+yRi7FA/F1pcpCQJcnh787mQCe2a9Sr/+so6F5
Lg0ittkwRTSeaAV82o22/zKGp7VVlb5c79AUEXi91vaQu91Y5qtSONpfnEMw1wL/
g8fNJ/ID/oIsqo2/1XUvTZMJ+osfHzal+jrViNNk7sgcmSHP86A+nJLnXjLxM+4R
w7yE117SrFH0o5LhPQsnDUvtNWHhRunbm0HDLpVa3drx/WLQeEjJch07d+3GcHLx
6A05l+xVAqIprYG52DmSzJFKjqWnA4ZKYUKsBfzJ/nIiOugOuxjme4K3xx8GO5tV
Aa1H3ddPp8PjPYquNsyh0x+EQdIzyh/dK8q+KqAYzpHLX2GCWd5HA3a98lF3DS9e
vCarmx+oBUHCBJ5/zSmDispSvuXMToM0Gcxx9/wlO9ckohjz7SPshx0hBh7MmSN7
IPdNWAgQ8+CRa6hxWm2nhbD3RERKkS58ahXeaKYfSlYa6SoPQA6JB8LDk3CZLaTw
EIoJfSqf7Y2+fp7psZrM96bMNS+8xuEe7wcq2+czrLYZiBGUZkoR2cAIBAkUK4M1
0cIc3tyJW0euGBucJte/y4uiisZnXRHbXRWiuSlY+RXNrFHHbngs7FJNRo8wbQJ+
vt6EMAJH53fx0RtcY79gY1cqagOeJEurKgUmMKwaxGMzQGNXS0LbAhd8JZuCsJJF
WZ1+C/UhF5Gy5mQmaFuQdIvw0bJaSymeercuYWX0HSUa0NjKaTQlZl6DmxL+W2nG
jf35K24Wug4wnnigQUxK0kuhNWsH14swXnLgIip7QtdNSyUWuUI2QHc4GG7xs83l
HT6uUWxpClAO1QVr++BT8xgD6XPslF42F02DuaIxTVaVJQ4P49EgZHYrKNdHgrCT
CEsxBpeGIn3yjuuHZ88Un3bp80I7VE7tLQouQDBo2eT/KX1efeU5cQkYSjsv+hbK
d2if2ofnTiZMdZSRKoVmCmFMwTOUvT+ik+S7Ad6FzDMYTMpv9/y9YyjKc7gSATnW
EzhsbNHPhu63TdPP22wkHccMxlwJygT0fnNpRzhn0H1I8RGrlGbNL5E0qpCl6wun
8joYNmOqz9UMv3yxUu7NhYjRU0lcm8vocE4tFWZ7jFrKSIcFFdqyBJ2E9v6xQA/r
wi0uETp+cheuWC/nVFT7TL7Xay8VOWYGmMHdYfgUL7+0ZQ1SRQafPVdA6yGG0qXo
8p7QuM18L34XgRNUm8scBItc06O81TZLk3BlNz/8mPCXXZMOCyncshmpYJfMoo0/
2HfYr29FR2EW4yRiUL5d9zQO9XUBctWPJftI9EopJf7IrM54w4KvCMD7Qwy9ZVld
1B/b/Y07akAIxWUpmjQaeJhabEUCm5rRDWRuLZW5J/jVR9nvMxrgA0coVRQ5S5Cj
on4bn65wHlL8pUtsukLKAE0sJwoczXmDyQkmDnz3iQxM4u2JAifr2sw00LGlkTpy
XCUKESjiXl8lMDmWSXWIv+1aTN7gjMGxA30ZsdZLvH3rhVnpfIHyCT/NHnGVTtRh
ET0ffjAHjkEG8AcMVD/A8QjDqLVgomBooR1YMzre2vPquLQbQ4buTrUMjudsYY8e
oF8U4ojhdTW55HUiDot0q5MB1LKu+j3wXjngR2vQWYel8/6DUwlBcfjnDooWm8oy
S+MSQ0/+D3PUUhb92MQOlasZgJjfvu7DoidU9mOZ7+udISIQ3tHuqjHdmwFQRUpM
ycIsagh5AzqsYy2ayD6eGJU1UevjSQ0TATvbBd8mvIQr4octsWvmOpL/j9VAa/bk
kc6yA0ybGjnm5jqMF7y8lqP2Si+2eZFauur3glYjjlcohe0zKDX9GB3SKoY/FyX7
sHifddd/RZ3xep4DLByg1UHQUU1rHNjPgD6rg7HVfGfRPGdb5X95L+0PKZmp4Eyi
kWQa7QaNDvJ4HAYNcUMnG/YEKSLE6bAKkOEtkkk/3T5Y1e4DNT2ooGuupdxkyINp
TDf45eVNUaAPQkhcDtf/o3/4iNZdK1PeGG7w94Pse+++D3jAs7Nqtoh8Y+x4KMmc
4EMa3v9TSEwTa0y/rpJWnQ73FOie9NULV7v3rjWk7yEtZP6Atbq2u1sI/jSRQwMN
HS6423KKj8etBqgWOm3FTWuvSw2DYTyIO0DytpkUckfFpb92j8HNP2ZlBALg0Qjm
63gduqB2HGoteuFSHffXNXdELArvxTQsMZqeJzSA9XpS4tglZk+C7U8FHiRQyEsh
eYxgORJ8mddNdm9oQujNp7ULilJlpoCI4L0u5f5EOimqMGTUAsi6sdQCdr5j40F3
v/TX2JIrpidKf5ZyWD8ciGA3fySLHlh+zraWmsjkHs+V0tfVo42/aoZtsCud2DD2
/aHexhZLg1vurd9yTHdm19OBQT2cyGBLDvE37yonWLOqR6FsAFmfKAV4IIE1WwzT
QdTTIr90TddkOZ0P71sE/P9aNrvMLOpx5mx66ONTjXHI16wpica3fYW/aZGME/Qj
pgeBTHBjmdRNEqjoHBdFks4FHQh2Dd46GhdcaLhAQuoUUMO9GTC5e99FhhPdMR6J
ImMbJi7w2yGjo0WfkmOYboIkoj+BYGUwDCYLog9gveumD8kcYWNCceLDCxmmeUc6
k05wLVSy084U62IZwg/foA43qDjFndEa9kvoV+ahRSFaFGceJLNHiJ0cBkRBkqiT
reubFO1KpMWUMobsSXteAUOtvlLar2MjoQQTr+gpEXBMmSFkUU1GmG2d3iftKiSH
rwAL0qgzTm1cfYChcTSELfezWK6EJmxzJ25kBR6AzuyqbGA+Iwyxwnn9lyt7tu4F
fITexJLhXT6zH8jr0rF9h+EHrAlJDPTR4CbD0kCGwjF0K402z79H9E7Rg7M4Zzon
C6Xv4ckU4bRlY9CfMjkFZjhwwV4qhZ373nUNhvIeRP0npPGlaCtU2Ce/AajuNNdL
M9At88uJt5NucEO1a7SYrTkscWfNHHCynuAA6bEjFIVeQSyIkWynEme2HSN6rWn5
x2qKc0VJF3Z1c3DgNG/f4ylj8qVfRAjO5lef2BwXA2dRkAogwAx/m02ZmsWEUlwM
qYV/FgV6Up/jbbTJzlov7WKp6WDm7XehP7V4Led5tdeBR4x/XYm+bXfWGRkl+HHt
3uxBrIp75h/9d2lkpWSzcJG8n8ORJDChCZ8Vt89/zPz5M1BMxbxP8XfI3UgPbCrO
PNNbOYvFZNKTKZf54CPly8yu1nhEL7fR8CpkDlEuDN/UMqA2Pxl1Id+WdAd6NIgy
grpYA3pmDHC3XUQagMMZN6YcdK7ztJAyEGnvBW7gVjpdOsKgfsnpP0wCCWSfvzZM
RXXPweU0aAyQbFDsANhYdbMLlUZ5vLx9SsT+HBgdlq6PSSavwvITDputTRhjlcrM
CRrGMtRNy25uVodlSSLxno9C67/ukYJnKwJDd5Aq4HgnjyxUARVQIpkOZpcQkyx6
3C8inX/8VtnNflt7697sXeAdz4e2DBbr9LJ8GTW+KGEb5iPuJfkAgsnd6ZeFUCJg
3E9+racHTGyvk2km/Dee77enKjLHxJ9ZIF0U/Umh/GaQu7YF7JrGe2rsOiLlE3tp
J+juaBYn/REN/jZ4UfjSHKVzYMx8qWjPzjNmJHK5sorhfq/0wmYIy3njA2PefaGq
63/xsSMGSQGFDbKRSg1Tixgt+VoQWqHZ1CZ2642FYL+o3lxURgyarXhukUY3JFkG
upqiXb+eyX6gO64k8fuEyhkPOOlyNUksN9zp2XM5u5xGcxEcjgd8vS1jA/X93tbY
Vbu2W/CLTlzCsWrOZ0wvZUYKQ+zotPTLL75M19PcS49mFaEklKFclX3SLmXp6tjj
4jof88NbhQTK0cOfyCl5im4ydXavL04Ebt+/YAodgPUlhea48/PCuIPSpXUrHRj2
32Hcvu+c//pyEVwADw6wANViRb77Le05qGAcfEvbkUwaGvkPVuzmTLsmuvEnFidn
q/gulZMK7h519aqnG4BKzviRp1ccXoS2xXDIm6dI2Tb3XbZouRTgKQOGO/GmrNvg
Nzp+FFZpPtzfEkxz5ZwttttauO21g8aEosMs3Sdslh7U5VJySuVtWRDjXQmjwsRd
BvoqoIn40sbFFNt7FZaCopVULMxaxPqQ7N9ug4miiVxyWwS7aKi/wye38czoLpx3
AiT6i/IJmUchZncaaTZow7LX3i7p24cpUHHDN/qdYyF6mD/elOWbynYwVLRSeZj8
UXJOzwHbWqoJqVgfOYhzi+uSIU1oelTDxtO3EvUv4DARZP5sP/L9qKcjTHP3JXFA
ruPiGX2XKbTQHLbvxfS+ac7KRXsa1qF0QawAoDEwqw0K5Rsa4rLmjctgHhRJ2CbL
bY6Q/1bDKK/kHON5kWqL0JnBBRnzQPoyg6/W/Oz5bamDfszCSLKuHNYL+L2w1wHn
e/R84GXU0uzmsTcZ961PShmy2om9QChgnaILi/6Y60CPgW+BlENvJoWjOWqMhmL/
QNOmGDXd3Tm6icMsaYz//rFsW4yH1QlAOO5LREaNx3FjjXLKxEl1b2TrQntbzt4W
rmif6jOGQOLElujO/V9ftsDtn3I2C6QMajG6LKdd1uU26Y5eHIxDmKctaqpVQIME
BO71pfX79hTi91DgSjoHCkTO8zK1ZkjGkf7K5PUWLMgSPkZRY+WnrkLPT4nxCs3+
PCxV5sjh5zSENTpYfUOoNbRWVRPnHN/K1F2FuA6e8OVQ9Ya3cVT0ap0nLeGnXAZt
VxDrb440c295/XTgCAuwBzffONLusdH3fnj+77suLOM5I4S3MLsCXNc7JiNU9t1I
u7GXoEe7rOScAKv4SN9F8aZJBpunk4BCUEinlDpDcN2dFPUQe5wuD6KOlUzjQz5H
OL2GWovWP8eHAf9fLtAuCfgoEB2b7RCh4mifh7x9fqzl+uIMYSrmTgaGL8HQcT+Z
ISwdHZaQal1gar/FlxO3orfptJ9IgVpNFJjcW4FyiTsNGTc4KUYtxj1KTVGnRGsn
/BdjTteHFINkZCaDy0wjfe/866NcdnDMdgabcVGhLr7HCQd6t16ZWveNiJH2jWnt
q4NuAJKRsOsIEExGMr/ppwraHhLLhGwycQxHwVwuePLcU+NXK2NAUoDUdFkGNh/f
gyS/mIKvHHHSui8VUQNZtWHgarvPZgSm4B7/QT9c6WQmcGK1SK6gKA5p5nY+VwZv
jOEExzr0WT9nrrXj4YLEHPs3UiURgOcJRKa23T6AJRmKLf/mSBTec0FPaiRfuW39
h9sNFpUjHA4WgUz3ddHf7UTHGGOwr1eWFFvwUnN38PP9TIDoe9FCHUFP1OqkYsd/
dUUhmanp/GVzL3edsd7eoCyI8mPxtjQQzFkl7/GnmzVy1si/OlhTOcjoGAp474C7
tCI+LjLP8SqFF0JXj6Tpl2JDyLWzQzC4XD+dhzUNFl9WAxnLj9cOwmB71pOhy/Bu
v2e5cqRM2Y2Uf4BGQRcZAP5yzar+LC2fDzs+xODiJ5DCLs4P15bZCzJw4G31LfQV
68LScUweN1FvZKS1HBiFOT+wjqVOj0YJRSmzdVivPsam1xX3XlBocyqDKbugb8W6
lK0m1k+C3E6SWRCuH4lwYGF54USkjO0CvXFmQuKbFsJ7KbVJbXfN0/BWtCHhAzHQ
qMiTXdvOfiwKF6EnKY/WmPgC/wmjSA6zSPWMZAtlpX/s4FUtgEw152RJ7Xk/loKi
KZ+u5Q5sIkSQP0LQyzqHq1giY0fU2yALh84oLGv9dG6Ml0Fp1l7pOCU6oHw/VgYg
ZhBLc8k9slejkSxVTgPQfi27Djzl0DD4vJne1RgbOwaM8KlUDCElJwCcWjmcxiOg
M7C/wvpLvxhhdnaRTlDky8jJmfVDl6dIrr9GN+kdt9ClLm9mtCAmIXlgtExpvJKP
TXSv/X5sGeWTSluxj9+oi35Zj0tHg6+IhT/QwhQQ2G/Gpwru0DukS7Lm5iG2nwPe
vyV+/uCMoV7rWlA1wTmGp2zUvi9qqUaSaOhSsVj69KKB/lDDUUUpkHgeRFkzt4zb
KKxSbSECW/PDmhO7UyI4qRF/wCcfBZkQu5/hj3C53tUfpEmha55Z0am80SdDB9CR
qvz9jBp0UjaoaTUhl9VU1jGD6rP5k50cc/4cWaZ6pqFdgRjSkwm34m+Lnfk+CcQ4
/AC/xqdJ75HYr0CheqQ9CtqNK7G9cC01Vv6Fzl17okFFhJl0LEsCe0VVGnWKjYb2
xWveBRpgOrPYX4FxDOVIt3QzP2w6r8SLB5XACquc0CH3g3LmoxrJ3CXslk12bq9T
jWgjb5LqCFucPxmVkFF4bYmrSljXGTxbVMSslxjTJ552TaRP12TpF70zwnx4uAjn
EgdXs+8NdSgkWPPwOXH+gyrqYxa5mHGug6LvWqNZhfKDgGSp2deNkdq1B1+M6ybC
OoLx5keyRF4tI7YmhDmakmdV037sR2BtbynkzrtyihYnkjoyz2M6swTcCP6AoqMR
4/mtGkgsgLgsjWXE3qmlST5bOw9raaQWu8FUpSfL6ebq5kRSFO3Yt59dT6HqAGG6
9oExPs3+sfsdDYZRyj2Klb5vTjvbRhDPnalMKZN5eR0/rMwgUD5bwrBGjPNkzCdX
J5o57DafSIw51jIq3OHdc8RCxOdbC7sUrOTvIJzflhd56Iq/Wj4fPTNbP5LLXE3x
wObzaLjdqAp75ik30R+Q9S00M1Yrp/2JsIZ++xtjbe0622l2AAW/mqpeYQlk+rjL
XFJtJ7xQ3u9hodj4q403SUclhTvVecpsAFEENjAEKFe6FHD+q47IHAZGyUU1MZyd
Yv5Ag/U02J+3qBJvi6pxARNnIlxV2hEHCUSYTD8bL+T4yrZNcCMH5ubCfUwKkywy
CPPVSxpXsMCkdgMbvaSSROST3M1rdQMP67Xy5OQOJptiDtNMFpPqUk61tWoyT0UV
IAXjuNKldrZeqAjISIioxwMd2Z6Sy+nmbKHEd5QehorNhGFewVFsw3zn0bCBVTID
V+Ze/J0K2Cr3QtY3SKoJ/bqYnNXvnWc2vNrw1nAd7nBWyMZ59qbcnCZs/9O82Bv3
9k7Jlda6F3axfbUrsFQlvTHjfH7CLbg386EvMPTf5+L9xb3QC5VNHy2hkmhx5Ncn
1FKbZIGMgG0RTuzvvsSyHjwGJBpcRq+/9ony3Pu+4hSlkE8xU+KynEUHv87f8Olp
JNi9SBw/R99BpFtTQhlfsf/vJWcwGf+6p6Pt9PZigsW4F+qn9U6nH7mHihzo4GjD
xxZ2FyeaJlWYdHfvIL9hMZRPWxqENtomoMUPpTpjo4ka6VkO2nGH65SrhDJ+keNZ
Gs8R8fnPBqjxdlWUgCL/haeAbe2uA4CSpWMOIOQCXa7Z5ZUQpvgyz2IEwuyir0rc
QbWZsZc8FaHcw+p+5VxsoahFdUcx1mDw39uveZhO4MH9FdQWlEcnSfuRWefjeUhp
6cTjQAn0RkvlmdjZpwG0Iq/eAcq4Nue3PuPShw1Hf4nv+84fqtREBoy8XiDXdnRG
pm59lptvvhl+hbAIsANAO4NoZZrbUH7ZvDvZv0Sp38ARb9+7olHE/iTPUzGql9j+
zi3l/5T0KLyKWNkwltL5yuz/xj76BZDXP0qtmtmMsbAjvuCoOCl56Tgx96lcwFLz
uqv1yIqSMd1vxSHtyqB+iVsailnIjgeXk0wylWJgBXMW33jo8L6mySC63gYdbuFd
ij+fqAvoM5bVxp866Lp/aeqGLnkhumgW4ZWs60uWnLJUITNEzDRh/2vYFD+6odND
Jkk47qEBOrMfmDXJ2BdLht12ZCqFLjHz/yMBb1xBQyKRBit/e2K5h/MVw2Q3T5YJ
4/CePcLT4UR5t0+wGYgHA3MbOh63G811T7nPR+jBUTGoH+S5jbA+759Ci1UrHSY+
CZlv1mSj6fxc5icmfZ6lywHhGOxE+Nn1OTQmT5pQix5yCHnqn0fFQlPvkk9g6Oeu
EqOn4K6TFdqfIHmluU9LwWhmUBiIXmNEzW1HafKphJ6SclKBAzqH+ADZA/US0ewa
mIDTsleRKkaNYRSOqYiBzAcz7qO3TvUBAq6qCOKZM3ULem2hixt4shNJKbfXxaS5
HYpBkDpnYortRHCWnnJy9khv/osjhch6Y+hN/BHnO0DVz3tMZ+WvXnbi19y+Z7Wa
v42DYaq/nX7BXz3C8DzOwS+FOo2EYmWMlhOyFhiY+LpkYMMtzCsT3Gix7C71IMXI
/xSrYX/m+KD5S62tRvE1Jdxaf1HNW0qm7Z8ZAOqHUbdwcnlL+lr7v9a/4rFr2+PE
2xxHB/qi1rFMfnLaazwW8nh/Uo9pC5n/7eidxOTYRJOP8+kJWKvgwsPS9QajYQ3v
Z1zbrpDeXYutll4BTQIzK3VCa91dePk1/2S15u+TyPKLH80KzY28XYSLsISgTh53
1z3eRTaJye8DYE6pD+cJB3HKxJMPJ1xx7G+ZLTbJ6l58BNMHECkJkfHCMgVmi2pA
EtEU36CxUyRXUzZ2Q8VYbv9T42U1mBeZ7jjr1Y9GDdcxkGVK+tgrMB1BNXs/ebvc
8cPhONrCcN0nOSV8zWuByPyFLdkSvrhkpbDIMjseajV1rDN0cnbiFhEVCm7vgi+b
xZHtGuOac/KLK5o00gJGroCAtpuMuhQo0HTklfzScvc0u57cNWv7HMqLH7StQHIw
8aQaGad4KKypYS5O1priMMK/2pyhJQ80LViQSbi3Uvd8zirqMBsNtaDKd3rSCQ4e
+2+QxMbHFr6pTJRD77a5kop2vQnBJt65njeheSbA1qGQQkBnvr5ZISoWoNI+6L6J
Z7FWSJZvieluco52FybH3zs5IEdnsPZDpN+7RhcpEeMakiDfV4/78et34RvaY859
AlDB+qTADQ/k3E0R5hfJ0sDse0eEZvE5boXuC+ETnLbuMPJEsTqURnu03rTQunx5
hzJVzY4pYD3dWRAQbydOwWyofEZZtzrib6c4n00Z4YMdkInpVmva4q0submJhgbg
cG3lz4KyrYIarPfC5NO8DIF7FqoHO8F+APfTyF8CJ4wHs4GrLcqhjQO+6Zj4HY3F
0FQp+3vvNv5sdPUrclS2Im73BexhXeISNrieebyX5YBX+Kx1TYYx6sC2PpfNKmVG
qzqrqDYsj8EzQRz7EKtBSupz3werWIobhg7OPuXXX+jcYl8Zibh7AzT/AFSP59gd
WGLVjMxIA0Y1iqh+RkHCNek1bib3MH2friBzV0W21wNxKSDeqJYnyztQ93O8IHvW
vlQPawdgiRWSctLgJkxtukBLn5KgupU4a06p4IN25E4l905dAepi9zvDCz0K+6Eu
VzKPMvwMskhiVRvZwn2JqryC8P0yKY3nnDcS/yqE+fAiLlDwMR7ZXmnP8SXbqMxa
o6n0BqZXYsdbrdva8E3t4hj6v/mz2t8qx36YOl+bALqBI+iQUH3+ZClSmNBWBbQq
86OjZIJwNPbeLMRfYk4rhtU7+BbyqQuC+sGyL3xFhdznY3eNJ8Bx2RXQ13zBrfqW
8k5a+dH4bHye+QkqkhFEV6jDgv65a6FbBrG97Ao+g6oN7uleGPMlCXehbc3+vqwv
zKZjyZ36o5nacyxuSPJdjPfNQ5CcNRU8qrj6Qbviiy9idURQ15111q0kYRHlrxnG
GepuraDLd4wqLdZEgv5IU2E3xKMDThxUP1PsA5OZrey/fQidKogsMf8AKXvRTHo9
AJGfjLNLTYaN5vxfc6GZZ8Ybp5iUMbmA2pAPuiTh5ndT3B2SWyFTHZ8mW4zrz62i
D2lUGISpAZP1HHHKz7LPHMgy7Qfap8YwbAuK9QDwDAUZ/UFPCBKpdyApgs6GT1BJ
u8F4vNuvzOpdNqQxbwqv0KhMZsLypQE1AFjNRzAllzw30EwDsHLxIZp4hpdRGahi
QpXnJIRNW/Nm/5pPph9e+E4uDxkLcSfQ9ZqRv2CzxrBvRlxb6fKWKLvmqc5JnX0B
rsFZ9W7+yAcAT4sLTBLHVrRGMSq6NEukXiaa2LYsY9IF0whA8DiAayrHfyc/7J8X
d4YaGw9B9NTdt0ulxySfgeKLSShRYoCrL5qyt4uE2RdHQWp82B56AgdE/a2hwHzv
32A92TtBcnQRxMhERUAjx/byIHWveMVQGBseSWWNaG2s/2zyZjnG+N8PvQmCj9QL
/7qmk7yzQgEYSQXqKnxEpFQ1d3yWKejPvtZmUlxlVi8oBTBsNzuptieLoQmfsDSH
N2pPbPJoo2QaTd0iSyaL9Rlkrf38Tm3lEl3knzSnOugFJ4kqtW0CKiv1oI86+Gry
62PzHCwrcgI4ZlwfcNgpKeGvXEnmwl5r0AHgusinq0DTcIDgcBLYEkepMTq8fWEA
pngzHdHeRNj5xKXF8bLil42q0jqHHiymrAMlPV3RaCMi2nNRg+VCL6zV05Lt2CIo
LSLXi/JLK1k3AQPngaCPKb4efMvfhKqArzAs+dh5mkjSMNOd7yYSeyfAiODKSp+X
SLSO31VXVVwdLTbnidwHTyWWiOdOnwK7/dfsbKLKY0si/+DOOLpYsmTrGBt7z/E5
ojARUyqM4+dZnByJKRv5kAcqoRkNHkhoMA2zUfTe5m4C55ygCvx26/KtvqoOjNIr
7XvQlb6Ghww66BDHTQjFovFJKJep5/ejuc+6qqdxCKuqkOEL/dHDtD3vAL8dT1/8
0PhXi781FmrTsiP6zJw0BVQcs5dXDb+Eh8FuSXZO0/0Bb0RT0yYNYXw2S5D3W9YZ
wSQbNC2cDc8vwmblMw0bN/80mcJEiPZQSMIS/MqSQ1DibnlLip8CklXgsMx49Kd2
AO7xo41zHSyenIwsU6Qw+Ha0WJ1B7e3lDUKI4uyb02Ic4s1MRaPBRGlQxitKoBb0
QxysdZjDHX3RJNn6PKP7Mt16SP5tZCdx57eGl8dl0TdqJhtj0tEZbn83nX7W2u4/
BxIUa0dPvBwHHDxjmnLTQ+Vd9KAcQ2wtn+97sy4kohZrzzuddmNMmLA7xMxHvDAk
nWO5N224QinDzvZ/7mSR/LOxfHKrxuWk26VvBh08BA59UudLu9Qkt3ljbbLFNzRf
2/nN9A7jC7xVWbr8I/tiU40ORovWC0gHhO+d/Fx+4m7W3CtPYhOhgVxBVJBme9OR
mME6SfuT4hWogav/YVXK+EUnJ1xa45j8klrda5RhPIKFFLpiDAiEmeV5O4nUKztG
qsCV/P9HAbfbFHTkKWjqDq2MkdM2Z9TAUHjipQbEfIqb8j3F0n3/TNGTVr7GQWYY
xSwNDjuE7lZL3Iz7CuauDAv5rEani0AQjVvd14qIDA4tJIuf6S9i7aIFuxyTcqp2
XmewBzPShtVxt1e+tGTKlIBNoLSF1YL558jq6Tkn5bxRdm0x4Td7NBXH37KUnZEp
axO0YfIi4j9m+98j2vr/TkmXDSnDHRS7d+vRarFjAFK+eJoRDs9A+KL3bQw9yTwI
usc5yMC6318nQcYeiU5liKb5gTm8c4MLjjgqnR2UYovCMuSSlPb0POLd3QAiEgYR
LkwozEVzWHHZ9CGLIoFqsp18SrDBy4a6dwCC+w6NMF60hYkI9YFcfMcKrrplkWEj
jL3sqmX3yI3GwTdtsTTo8U4YWEcaSPYt2s6LMZh5SaT0nwJtS+GMs7H/2tLQztM/
w3EUAVSz0cNJjIvfvSvs3pcYH8E37nAYfvMOfFBtFlyaeZnjuCtMLvrtu34wHHeg
Mo2KeyO0lmKb6p6SPU9n9MXFc8MszxAunN3pQNtve7yu+Pq7yO0Gr2WWABkHJPpL
kjFW+5480SMQ9CGhLGQ3h/VQGWO4tGPuNICB3XSslw0uqzwYLAc6P6ImoKsXUhd0
okjqvIzShq/YbaK35z5zrQdgKkEaikrF0I4kT6wKnTotSWIFuUi/es2YH6aHhxs0
AdUMhd88gnc44f5Vu+IiB0cYmG92Ui7k1vuE2FlIeUlI0AEX9T7sL4JjkYY0a08k
zQUSVKVx3V4fd6JPWSDDDX6hHqozsJFuCBpct/mtqewe6c4xUHKXH2nEV3l9cs70
Q92uLn0+qmXTvIpPF0OehfFH8LQaUfNXan/S+qdMkMrtw5H/eeQobgBNKjTN/6R+
BVlQzPnfKOhTsp7dCKQwfQcDXKxdve9ayyJbeLP62smC+A1Qi4nMa4Qgbj5xyQP4
RrLOnvXbDj3Ox+b+y2hU5/mbvPQJ0T8XSPzBXnpsQYy96GtYLwIdt4tF7PGy27xR
FAkmL0rDSVChHGcr8lf/u4sZTFB+oGGoDtq3myygXZifCwlwq2gyWlX5T6xTL91y
X8g/W4cK9y56POi6xclzNxuAndCA0YhTjBlHU19NkOT8SOs9raJniADCKWZvBIJt
wbFCQ1RF45eCreibwQ96Q5lHHTXlUXtpHlbgB6QSsPr11yFv6T+KKZg4mfw/lT3V
Z2lGa1CYCjRmlgy6bMNQLyMNVhhCTNRpdyhUGzG4hCbyGI8/cDGWYTQTTcHh2r2f
Ev0OiJneGNOEaogIsuuxuZ//TONtSO7UFasiPHub0ZF+qJad//RcE7ewD4uYIaMC
XQiOBMLDZl9IFtMYKj9Pz5e2Mj+gl1jitJUyAajVE6uaoVH34vbPjc90WRwARzsC
Lk71R2AM1W81vFWlUnZCW7cmuSCa18mP/1OfgHU7hKnPLV+mlBTT6UbCIarkl7fo
Bv3Ia/IJcr8ZKOefILe4xrsSiQTxa3Jt4jzALa08waeOh0xmdyhx6WNgavYEIp7Y
J0LY8I+dH4tjGDjmvhPD6YaKHZkphKCCm8gCdcYx3jpCOLigiykHfWDyhvELNUAn
A9GGWPc8dwoLLdbdykkFsNNJp4OyjrqNjfP1+WsFsYku7QVWn7XYLmsCXx3CfLvw
4Guo4e+KQrwzAwaFW1Y+YHkkhWaE/+Hehf67Wmqb6byhOSKdYx8uFyNYXiQRJWQx
uEEE1QjKOZYSlCSGmfma4QAVtbPpM320VEgclpELna8adOKAhysC83BYxcIG6Zz1
SY7P7KiWGuo1rRg+SyFVTNvNHG9VIytvY+HUgQSu7oD+yBFc+W9+w/JxYX5x8iIC
2mrvLmm3dg9ROMJebK4OgOXiJ40kWTCJtkd3lvHgjfYUEd1E5ovy91dWsVnpRYFl
XT7ZYTKAUPaPc+nkx3iBnxvYjbWPNO3wB9j4KkgKFIw/AxPUuhOrO7eHhviPFqc3
doH3SnFBszT2D1zgMmDB2jcUgTEaW2V/95DukcwcD+DS687FcpfN9Hl27lYKWbF0
eXArGdTdF2zrv6iSPLCdKNzYMIPuhJC+KT/Ocw9PenROfXQwbyTnutAqUpFlSN1y
GRSMqcXgH2y37alhKaLJsBnMhs1jpwapeshbo6jCx8j++9stf5bEfyATUmHjvMkj
NFmjwCYwebA2KnkHmbEXlvTo1iRk2m+23jb5oG8PAUnDAU0kn0tlBeOVZKQueTuM
Zbl0sa2ieisq4xn45H2WxCqsZ01MQoQn35tjny2E67u06nw15bauFROqrks3DNk5
NP46Jec00yCmS8KkMbnHOXZW7f8miiGHt+qQFe4rG11GmJ/rLsxsE6thC+5k/KWd
1zxvYmqMF2gzgpiLFAzb0v/+c3brePUUSuc0ukUJy0LIOnixm4dmlag094aTps3l
N+T6ITi2nU/igHxhbCKdQZ5IxpP2NdU5fSilxwg3Jom/8d92+tq1AU3p4JB4+gb5
R1bi0f2t6R4odM7FLq28W0qaycY8+ixokS0iH8Tythy+CFjZnBQgdb2J+X1FDhbk
Oce+mSb986W6a0GhqDHEa9OHgslI2PJWHJroL0/UJ4Sf3dF0QMdQIrVwXlGJYLZH
ET07/6Uly5RT0zVVXFpyiqWEYNd4hHGxnpH2fx29s8bZRu13rASyxuR7IimPErZ5
ts2oCzpbKcfwRUnqwWPGz5pRqkGrLMGGBIri8pJ2S2Ofoed4OfvWpEZQpupkxlgS
MQoSAcZzrI8PhF+i/cZewZOHlDS4SxHo8D7+iDL2fAXE7+9XaY1LNDL9wT6REp8R
Qk+PlnXWNog1aX/bRmcViXEjgkrFPzZrlw9CIpQfAYjVao0PYUaSTxJf6Wi7ZjaZ
1DR3FoRMoT3tqOXi1HlkUyCPXi7+hYmrOO+LgZXRcXb5ocKf5yh0OCqIuetO/rqU
k2V27lbVvR7TtJmwL7EHkwCIHFcmBkwEIvbQbaNffUtif0ZIKxCUhxLS6D5DbtM2
4DZINN6vYem5NyhDEFPPv7EAhjlFOiOhOIMzG14ui6hIvXgaH1oiOKW2DKtQJnbp
sYS3WHpKkiufdnZr0e75UvFPWJTByVF7uTWopJFSy1In/37G6vbvsly4Wu35mCrk
W70SFqRP4t1SDc/cNkVh1oYQdIWFXrGEv0fWR5FsDzldph2uZaRbdadEWXq8kqY2
kAkY7gxfcJW8nelUCXoQ0PFUELiEe21agxloTPMf9CQvqpAkJbDhla95LvcrcC64
ndtyKDiFObKnJFnt9pUAs9/f832NtYb5FQ/K3Y48LnFlNK0D0BNvTyqsEpJEDilG
O9PIFW9SviwGkHLBJT89wZTn3HOWkmrtfO3yRg0TxY9Xcd2ZBL3q6MQMZYk9gBIo
XyPLh7bYoGLLeHx03ad41PVUpKVcKGrCMA2UEJeJzfkMXIMArSk3nGf0EwPW6yVy
sfprJh54TgrlI+rAG8rWWh3B0bsnzxvGGfevUZpPiFxWc2WT7jq9MAup6rF1SXk7
RgpSQwOMf1FrNsAEl6ymylkl/I6sBJx6ieFATe6l8MhKE7kLBTrut7sMH+yQh8L4
NH6JQqwVFaah3s3rE7Lku4eoC0ZVQSLIlmjG+cc/pWq3Z0+3PDwN47L5ltJq8VjR
yN4tEq/V+nM6ZcoMEG6JlLuUfNeJpCT2tkLqVP6CliY97c1UXDFmXU7ji69rU3RX
xc8eikfVdBgyKN/jnEDKIvlUiEW7Q/IOlu69R5YA4/GbjA2OTwjeMkyanYM/u8+d
mt1IKxl+GmG8zhSosoad1pPG/atiqjWAE5oaH18i4+wHHMrjXbUiw+UQ+W+5R7eV
HOIPoeBDKevFXWOugW3w5paus/mRi+2+jUfucvem6IxVUFAMxSq8GFxtLfb/uQns
U330NouWbSWOkXlboNaTI0dU8ml9opFe0ZQ+zenQJEOD0sP2S4SjR95R8LPNnoyW
8NoE0foR/OC9u3jEDbx14hjvyobRALlkNv5/KZIGbAgyBgwgwnyT9bqucZhRNmKV
9unY68+gImRV+6LcCgneA6AG9FFNbnh99kVfl8b8mS80FIT+ks3VPfqFH+RMhXzP
w/ksjkGmaIuyUYxj+YxSiKOv9TiEDmersDk4ihqPnxgbQZI+Gbh3SLH1Gn4hkhJC
GVwAuJF79nANuzXVxbf2mV0xVrKfuwBL1AsFpiapICwysmFh8kIdcVcwIER1q7oQ
0YNwziapg+e7uXs6EdHk2VDgAkPh8BZy0R11Rx/P3pjw7jZzlozf50Dca+AQp2y6
x6Ur3pckcImFVCluRxXsP/KkahmERi5z0DYeHJ+Eu8fkgASkCiH/PYGy3G5MxtMm
Y0Ia0a/T7NO0O61a/07M2wqJNajQSVAvTCIUaW8KV+ZMCODRZQYjYFL1yWp4s3LK
wuJgeYH5Krk8HIhFjR8gknFwyLyhR8pU7YTMPS33tW7ExibBhmGZz5mNTHTmu4FG
Fs3VeuIzaKCjkYa4/Vyhq5rbEi8jnikSHBvm8jVmrnrNpZD3kNFUSQQbMu6qAH4p
CQvVu6cH9yEFCtEWQM8VjyJfm9STQLn6m6KzvFX+Mg6qIfl8kYPNQTj7FiAaetzd
qFNtW2zXJjfDY3uMeMZ5yuc01gO+kws9uyTn3haX6cB5IqWIMtC0+CsAiMuJm3a+
hTj9EbgQmUQs8mcHfPhcs76r3Y9kHZftKEZJyEtfpQFFgDkX1Vidmdbs9TsyttF8
cbEqWnItITBScrRyRW8munwBGhfjL6ITH6Wd64N4/QhAQK+iW4fDyqyw4dafdGGw
xefP6Qm/ylCfRgzy+m2XHjJib8Zqzo79Bl2fWshbIgTGgmIIIkB4vXfpMCJ+xoAd
k8yw9TJq0hzF6lt8q4l8R9H9iaUFAMBUxaLbH3GTUhakmIfATQpKbuJhKvoEhLQw
ekgECtNWDUNWb2G2wrLr/VYjgvSU0lT8KY43TUigAN3GJY794NN2S79SknUa2lN0
YlNhQ3maUr8u94qHCCmExrhYHaJKDm01jEPJmeObetaTFZnH+dZnvmXVbAvpxgLm
+jDJ5YUF1A6Pnmi2ZjXoZMszEfkqZ/tt3D+eRYRPAIaNY7F38yHQVOA22shBm9AT
nBFG/qWx2qipnoM0/Ld6Z922eGsltxBbnq6iVJErRfAFe63yYBDQ4LPI7NPXwv+G
iSf31faRrP1ub9eFLPh30hGrIzkVplb/GaO1ZIvtd9BY3fSI1cQ5DXfnC3J1Fo3J
wr4/2mY/kodDMhlASgIhag873KbNXZ+fmIJgQK3WmVQ2uu2DRAB2JfKc4k/njokU
vlkotleQ3GMDNs04VDFwt1SZYT/zApC5mVFRBsfzS1q88nq1buck6kWeav68uCf8
1kmcl6b+ReC7ds5SAf4rDtjzPtnMHD3aIYqGXKBzdk1wJ/nZHEVuDXBI629OPW1D
7s0kiizS6PkGKhBeZB4xdzaLFpG8x3/2YChQ7fwFwusRonNIOHhHcK7KBFtS9xDJ
rPJ4DynIskUgIQz4sy9d06FyK+wJFHvL+uSAQwkjdNVAq+YaqBYdUvqXgXui8KC4
oA906vDpzBj3wei2UjI2iykI0J8I819htZ1ssehyrDiKWKF4Ofa92DQS1qPXloaL
M+yg2wLC8vgVJ9PLhfcaDS20UJYn8TMLvXQC0EBOYTrRM9od1pzIb3ywcfsfk3GQ
7chqEQ8sY5I+m3IfW8/bcdgOVgZyv/J2B3juYOWy0c+/bWUgA2Y10QSQTunUExIh
6oSWH2VOpwf2CSIv5vEjzZ1l5X9pA2kDYuZuxf+3/VqqmnzDKDoFbRhwnXHhDU4p
4v7x08xk3Hua7+RWfSs98f09kf+ATCvRouJiH1LWgQ3IUQxtPKRP+zHT0KioM7oI
1fWaiS48fm62dnA6TTZd7jnekPsQ1rgIBgE3BxPMI+DY2/V9fiWXlZZBsK+7nx9z
NJapiINhQ8vRPv9j7MNkRjHL31kdCpTzSU17KaA+b8WS6VVqn7E8zWZXXg7iMPmA
8VJXqH6aWOlt+rCOgOw3I7ix1FK03ZLOHhYv2snjRQJZViknKETwTPWa58ECJGyB
9OeOrl5jG5/0CaL+NYZZONeabyyeW1jkbPYwBdwni6fFreDy/eGOT1LHWaR80pIq
iyIN6Gl46+LZwgk298EIVQGHU9O2NUq+udwqfDU8lPv+GX9+IooDxDQTtD7nbt6c
2GT/dwvzlwzn48G/ct0Szi8t2spJb7VLhK18H4a2Lz0vuN1q3J8z0rWtVHxxzy+f
iERhfKQLaDOZynQ4BVGvBzTrXroKxEmYwgQkX7C67Z3Hjdj5Yoc6Obx/n++kOcf6
yCLTEfRXbIFWvv8OEKBNeBTh0FKAaMvBoCkDal4tCPc/ONwPPd6h1BO9WlVkbq45
EJWqshf+hJc+0OpSINot1Ghv/DvBuaxV2yUOUyuaaZisJQG3mSc9l6Vj7XVqftQJ
1dOG9Yd+pWbz12+a75pLMS5XovEIlcZNA8uuh73Tqtnl8jexvz0gyOTILLhytwZW
q+92AhyjSngScdznwQQwPhp2TAejLyGPOapA1jvHYQOAWCjEo7/4k55lBIB4zrn1
hGPKEk8HglQTGSA0vs4yF7yYzEZAcojA/plXSoEK7B5ePDE8Rn4nCCUfT+mDnmNH
8EeQXshK5MLRLRZF46odCZi/Kk5UcZUsZgOVII8eNT1kCdugH0Ew39Dy5+xiCmW0
aShsbKTSCbp8HqaM3h2zx0MxTFVe6ziqFEdWs8IGDT5MhOQMndKFz+drETLD8T2R
STdzycruJvgwE7KIkyMSadHJmQJIEmq3XNBduL2awZq4XpqwhuvDYe9MTrG3+e0y
AUfhmyIWwOJs0UfSbHg5Pb8vTMykmcUhYEPDAJsSMnuEIs2HUBpj9qQdgWQIjpDO
6zmU2oad/UkLu7vofNivcJKqVa5WAeKcpY1LWFblnu30j8bNlACxsWbEH6e/ojiR
bVbf4DZZml0SBYOpkOrLb6qgYuGkgqB2OMZBj/PZkWurhyEFQbt3Uz9ZAPCNGOWl
rhoWgwWcUPDyJ6xSRgAEFxDCGlnRrHA7O8ZkJIot6bOsOBLerlsgCY4BZnpr9PgB
nFVvEUafndlRu4JKLECS2HKscZwWT4LCLYu2UHZJqcMn/MHp0ETl/QOi5j25sWdL
wdPVNEgaqxS05km7z+IK7Z9Dfg8U9IGRneed5PQbsk/620oZR6mLhW+PEaWIurGU
iGnAMRMLzRGLVOwpIPTRWgbGx7+VRo9ocGWPvabgtcjM5wDR6AnFYpntgSNMQD4Y
BMJYeHPCwfUSipK5G0VwcYrwwBJhoNaY4/KVOsgh5XGXojaBSgE+AZc9FlUY/bEe
1GCy/mDJ6Vh+kXB6KqP8n6yyd/qN4EatN4JvwRxqJzqLG+kUb7EPq1XnXWrqW8Cs
IZNBqR5IrtGpJWaM7vG+uTjIkJwtUKi5Wmp14LixD0k1Gosbn9zUJ9+ZrGkuVyHZ
B4/QioK8KuK/L4WBHlX8Wjx/VUcMeO4Sxq0Eyn5VbnAi2fid7daL9Vcss0I6aWwg
C+GPStiVYOpHpZjtho290Tb0wKaM2GDYa9B7b+UFrRckGZjGPBz7ouPgIfDWqeZJ
KOx3g37usd2fvKP1b0HlhTd51qU+fRP3GV1jKDz6VRGY6jzoFASYjzviQTI2oBQo
BxznoD5Wz8XlURXYjjH/7nWgdVazzhZza+6k+P7IjcORcEBxamkwmlHefnKagNkm
qmroQ4w26pRyovbLEYznbxkpf+xyGNF/wMsjWU85UHFc4ZWeNp2rn/MKTcmktOuT
lWXypiON9hapaU8gTRk34qzrzvBP7Ngnu+Njw7ec2N0/PKUluYxnZxNG/JQcqdOI
dArX54AuinuMmPAU74GviTAhSBchyiK+j4OhOcLlC0pTF2ks+yFlJLbXiYIghI8b
LtHTFrzsz/jRbMkEL5gtXZJ6oOEeIISsssa8G3f3jJM+GMnfBhqYDAPGe+t9jVM6
utzaBbWjTbXhny+D2/R2QSWsMZ2xx/kCDJruleOAUlGWYXsmTiHvItVNyRxOMUck
aC5U8gfjtepoL3JscAxOykb0ZleVjOslUqW2jDkY5UnahRTXTSY87iMknbEofkf4
83FzD6YIbOQwDdAPVH09GJyY3XrTFjDezplmVs0gYUpbTOAmrxKOSWFDdbWr2bM8
IyP3PHOAsyACFlHFPkNqn1U3ur88HFx2MEpH2qsYxBHYlngpDKk+dyWkdM+mtmxJ
9vOnU7HQ4S0gQe1cTlHpDP5cnNQH2i5q+JBcnUv+4UTBbWRY/iriD6ejPIM6uxVr
mwOfNYy6yRKWMrwizQcrYYvnZS/gy3Yp24ep0Q6kSeECgYhblGPPSQOZLfqbYkAs
hIi5VRlKfG4dmY3Qud5HnKnx7Aa7ZWeKrAuQEKKjGjtg122vKvM8znT+INalob+a
pfqfSowOMi6IN+gsQ+GChkZOlbjOXOCbKaXxqfy8iHkfIyrsqUR9WyMVZ05rGqog
Q2REsmOWglypFAdlccIovoMqdUixFts8QVjMgk/WklbRJHi6sl+aatv84C24alFC
kmqP90bLTvKv3bIc2HwD3yGZ+5xAhFzLZ5trECw/0v8xPf4oN4pHzFXj+OQ+buoB
1ZuAySszzpMTesFA6ADw2Ry+Lte0j9NdV7WNwrNtSuqlD7lZzgUSpGqNG2O1uGBA
xw5FfstKcw/+Ycl0crs4Y9GP5f84oa0k8ZAT/L8ntK5eZE6vRIHoTe1Qi/dyWZXk
iE+0I+eXipxD+ww1e5WBW8Wmx339M6nTdmBO5MkIwMKy2aq5VMZ3DrMSGOkP7EH3
PCYZNgW7g7sGPwfzZ+S/fI3RWNgLZLZZ+uhBES/yjEof5ekRqD1BO/3fkubHI1Sx
DaXuCMU6ul4vqnTtKqMZdHeHqMRqjZDOf1PA6QZMNmq4DHwBlk+burJUoaRYYSW+
ltVzb0eOLitWpnRP7cb0c26K3neCaX5MDOzKmFU9iWhEkqn1T2xaQRwcT5oRC8s5
OgMCY56fCTjlmVaeHxpBS2n1mxccVjry8RBkkV2lWYi5ve3bPSn4CNYhA9165Mdw
JDaBI7uXLYjt+usxEbqLbU7a90mSavEYKOmDawrVqaI6CFdGePZr+C1j9bAVQwQy
W10FVxDfekLp9AWOmyI3fIaU/Syrh1fQ1tJ+OKO8gWccYUKhvBKKty8SKqAg33tG
xTq0XShW2rDHKM2LzHN+PcslRDSIzRJG/VWEFvJGS3G2INlYfFyRy9PIAoPx7wNJ
M/7IyIKv9/KSU2KxHudS6Iu8IEf2z4dl6Icp+yL0klaxw+9CxbLdAJqvmMpqM2lq
xhLV/CV9f0UyEY8/+di/L1MUIruOwMC4QDHuqaB8C+hAY/bp2gBmnISWbZzffCtT
c0N2sZIKISiuPj99h4VASN/rZnrNar4wmUIMkq66N5x5wQM0uN5Z4DVjMxsye+Gq
waWWFAYkcDvPATbLMdFNGpG1/2cMrn/M56G2rzEicqHB5hFxJUfWbo6r2RVxD2WF
0BVhIZER7P1zd90Q1w0l53jkbGlj1tTAJ/ygbALMwi69yoZzYPOnYmpjZIiUD0O7
WhNadLgWVMNwsZimJM/nGX2wvmMmNjjPaX1jYt7r2MuTJ+WZ8Y95kAVf5DtCQ0Za
El33PMJ9FkfCKBREf6GmvxdCEX354E9RtjRinazokFP5vzKYAZyRUqZyI2Py/QYS
aMC4vOFSuXdUWWm8ygxOyi4N6rq5F0g8PsWzsgiyW6zMeaIftIEXvOVgLYHsg1XT
vunhMUxKzl4ptPya9JTPvq0ZqUeC3QTIj2oXvyL9udwlQTigtFn4clcEyJ8McTt3
aBnQjIkWr+Cb32eqoLqCP9RxHaygDiC1ht9VS52ArMoWa6VH5MVoYQIVCsyySJbZ
hSTVkm+1Mp0Q8/5dVvRjPlWJbJuXbt9b0GvNzdtmxHcHiX/z+Y4+qISteiR4IHf7
+lcvlU08mLhXRAHbf9b1QsrMRQkY7nAatNrigjmgJtsH8pHLOnActt9XQrkmbfkH
FTkMQKmpTMzdIYqLgCzCds12hh7MJFG8zwugyllxbqdmjCfAmfObGv5hfS651MuI
2rxw2nkZxHJ2g/8JBDQrGwazSxMOjLhTxXEhvVyYbbioB7ryIWsnOkobL8d/09Uc
fG3B8IIaHfCdjHUodbHhwOg9hdBF7ibK3xu5wrnItFX5CVvIOIIlzG3PETdC+4F2
CEH+i6XR6n/EsJJjpVDOxL3LEFCRQNj+YzCbeT/1AIjZI3kK2HR75Uug5qi9j+Gu
xm+32hBHOLRhGE1HBHzK6Lx9+IDR9PdiWpPEQRFuNZbf5sqq+jOJ6XOjX/Wv1v4j
GhT5UY5tdZErCNf2+7RmdDYQfWQ/Leit5GPWvIuFL2ft3ZbVoeNGmRYcgjACDpD0
TkQodEhfHv04VQ63JmcZYIcaZqwDIQ09br9PBuXAhUt0kjdIFCN36Ehq/DrFmQRt
Y5fdW5A1OcECtukJvHW3+Sk8JqmB6tpLhUYAYL4douS8FVOs4zGovY7TDfUAJ6vP
ALLhlNQV7S0PtKkKfUp8qQFYIZHISadcLjrhZFVG6xbWtyqALhYA4tRTJH6RttlB
D0pVda1km0FZ/2+rX9GdxXN2LNYeGqGY3yZ0H9u0vEHdvEyZgsKudqWxLSVsv/uS
RiWBZpD2bW/Yol/IxPBZXqItiIUOlCDfGttdeMLvoGh5IyB8JhjaRBAdwyqF/5Fa
tzKg4UuI0weWl7nQzhIAakmiLjF0VfRPW0ZRsjWhmKs/XpAiCJimGPCFGRqbFX8O
XxAL+PP7b9PdcRGLmucjRT2F5a3Iy80fHj3+Wz6/ce8vSMm9L9VQma+V1/P3QH0r
+VVuMP+K74Wp0R72WhqT1FUSx/mUG4kaGG9Ex7qPBcU7lBthnFfJowMXcPy9Usr0
rWpUvlDRl0NwcFcFp7Sb4RMg57Wd00KE/HXaf3Zdtt6fF9yIf5jXmtbl8W4wV6h4
tHScwHyDJvsU6VwmXNPTDLsjyjoxY7LPrwN7iwR2M4ciGjSXC+XTqwvF9mNSFhYF
KaddnHCAVcmk/fe+bCG+557D3SV9wvIVvU1FkgLe2mS0Bx8J7QUpqFctJooeu0db
Sjn7C3Qj5D0yexVzbbbdxbHWmEEsqfSBCp2zKP8wAqZJXKoMTQoGjIAiCrx54xWO
DMXbJHw+nZDGJxa4WA+ANKABcE18+ctX5FpidjO/+gZT0YJvnbBNLsal9gDW5+al
Nb19jmYxFFZNM/ie/wt2Yq4PMUn5ScN4Rxj+AVyXPqKWRvtUwTvNNJ1R7jnpPSvQ
qyZ3FOM20Tk35wLmhsJaaVl1rEdvu1vmueOJ0ETiSBaCzOCjJjrVD56Sa+HragKm
8RNPEAAQXLINy8DrKCwEcfuDVWHafObMkGTVC9nqzIf5S2qpv4qACYbrJuCDS0gz
GAtBFEA5KNeH3fEr+4ZNiaVK+TE9cEqcfilSO8en1Emzw5+h3ncZ1V3ksWyQ/Mua
hvj+m4/o5Fc9JSwuR53agal4h95whTI5M1BCOurx5fafbgSdn4I3pkXjPYg1pEdV
CSscrTV9WH4y7jvOC/u2s30+Z/beu4aA/CFJsKmmfZtyikxqhwSZrDWj6MnJYOsK
vXhtelz3U75OiI4o26PMS4mSyjnjECdspJzDrL/DbNXQ6gZnyRuJoFghTqaKaUfk
z9+EksYF2fJQF7gVP1buCcEy8ANYZ9KtNl5FkyF9t0IvQy7nunpctl84Wr+3yo9S
DqlWRc6bDQJRCNtCR9WWT5bUQApmrlXgHtCJkFCdkwoDF58hJi3v1sKi4j7hVkUj
KIHogjaUx3H60NkO1FWaWvhPlXhXf2dYxGvFVSe2P7Tg+oMegPx30RVr4S1o9eer
3SyYRh/4VZulwSuYK209OAzeqn74yXvefoUeY+Gql2eqtU7TWUIsSmxey0lEwdyD
aKNkwFqoYj+XQRRbfpMyAz4da3pq24PufIpKQGD4YrfUEOTvVgRMvGg79FgH5xx5
9SpbXjxDYe2JRabuOdJQ5pXuSyLGV4Iek/KWCc+8h8CZdg0k1mP+td6tqDEAh7cJ
MhP+8kECAPJ8J+Ehw5NM2kzbyL8jJmpROquiYidQ+JHE/hCDfyfuoyd3OKkxWMFd
Z+F0RUqa4tg7V5RgUh2amLpu1qbyIqW1cBqbYqRqUTuOURGBo/JT6Ynnmy0f+xiJ
no1QHZRYNmQ6ez3TKD0GLZAcUkU9anXoaDwkAR8nsln0GZc1Q/hGtpMmVh4EOGNU
C8Cp5ur3dzijuArDAy6Sx25evVtqyS2s97AHYUZHIgBfXg06oaYz0Iu6lIfyRspo
Z6/X9nRGo3p12nWQWcV+r2d/g9QfGMEP8iCFoWHrc+9RUcBYLL0LODxYDUdg53o7
jxGF/mkADD8AbvzBHZ0eIBi+p/UvlulMVtBhc2BzuytfzxGaUJ+ckpi+mYmUSN9J
EcjKvztkHjDPZO2oLSrTePeEGrv17zwsV8kIK5gQs8rPPTDcXiuzISRMiJeQ8ewt
aGQtF2XAz2FrZ4ZsnonpCd3qxZnJSy64ogdlDSO9L1zBL/saBBU5XYUSxjBkO9cy
irtPYAl1gvEE151ZHhe60O1pwcuNBUgSUkBiuKCB7ESO4Qc0hZAjaXDNrpVVVaha
EY4ziuV1WsTEgO6jgAnx8WxXJplan4pO4HouG869tkJRM2+fPbjKFBIHoNIWr/L/
qOIYdesoKG6FWLrfn+zXGve9eVjvfD12AbDL6im7gzQijreqp8XT73tMhligeSwp
35aeh52Jc6Nz5V90x1Hvf/19rW3TU+C1cLkX12TUzFqHgQ5JWNOP7dVflmd6FWVp
THwdDPGkYAOzG79CSO+VYwF3ZMC9dALZn5Qp2wcSpMZgPcbcKwLOnWHgvBIjiCrX
VmLfWWlZTnpDIPK3MvIWa1YNN+G7XcEvpA1qgai/xhrO0Q0iSROwiNqrokQWHKDV
+MPEqhlfrPsENqeAuEYtEI5hbnHnFrX9g+kisuaPl3tcaxf9CLLIS6Y+o/ODRVbl
hb4G8OZoYnPXwk5YYaq1JkUWsOMNiBQuaCpG+Voc7NjK3/cqvUVZBJJTi3g7ugAu
NRQ9CkOvoUlRRHhTr5ftRmtI26m9ipUPxnZYZdcQfrrE3HqBxHlNAsvdPk1zE7wB
1LSwxRrlK3KDVtwmNGRu/wg7Now3oP1fHrONJP1W6g/npCsI3Mptwt7M7FbkncUG
/TDosSOJRHMdthFSP4hbsaFOrib5DV948NEqYtlrWQeGjEdCID4Mctc6+nUvIwA7
kBLhDq94xJffuulccCf/QZpYnnZPD1f/op7AZJc9FNXTPYMNXNUz/OQIzX7J0vBi
MUhgbmn+gvFJIdPrBKbfzRWl6cBTXwNDfJcIRMjKiiYmYl5Gt9PpoJNl027a9F4l
i4bLae6S0h690LgJ/rMNT4IR87Q47dByHZj03IRB17TRQZcm6RFxCCFeH8U+Wa5g
dNEMaYCd0cBK2WqJXmpK5GsIwj2y3jWY7WNbRPur5J63Q0Gp/0Uuicnu7Y5gYsV6
sTjQM/hiJCa5ueP3rRoXpEERLb8O7jVySVPxHzYQW8HSMy45/b5aivmQIo/bTnK9
/EJ2XWEwMaQMYvT0jM77HL8k0m4J0myRKd8IQuo+iP2pZaDEh42akt0V4B9nV4+T
7kUfJ2xafFG1k64svUKhAWku1AiuOYIfRRDJDHCMXxtGj6NH8VzPOf2GqJQ1PEpU
cLOfLzXBHDB2ShH0g8/zVSIH9+/j2VPATD/QyFjuzfjNg0V1VBUzVcI4V3eq1TyU
6OCu3XBugnRUtoVbQVHKhoNW35NvM+3aOuNmVhHhDWfg0jPC5CEksMrySnEKANwn
hLJWNaSSeFA5cFiPRkCaQPaZHR3kPtLg/XyUnOvknRaN2xV6Y4cUnK6Ci3mqfGMF
otsRTDSMC809/DGubB440auvQJASbsmsReF7ZZ5fXBddbKTd2If+nrs3KvUf9Os5
5c0HODQQGK1YZlTxhLlj8HeMdUaRqdv2mKJXJRl2qzM9Wk1kTwStq+KSzIXBQg7L
qCt5utpPTpRsGQBBdmMEjF4K/YaRgm9vXjh2ofLXrTffKn0LqiAw9h+YRkBYyfy2
JKo2YNitCV86jODwLCGmYsjYsCT4yDdVex8w3MwKxR9mhWi89sXfhPMVED4o8Ld7
Q1PNGcyLz826x/ukqWqDzN+5WpsCk14Qn9gEvCiFb07J3jbOYN7X2Hg+7q2DEsLz
y6AsfUcEV+RXhTw0xgxmAS/WwTn5J6YryVfE1//LGZyEDJAWhUCzxcS0bYLEFuhM
ppMnT967wkph4mE7I5w8l/hEwLRPILO6hL+sQmGvQxHWEKsljcnR8r1wmxwkbnfQ
oWt0mGdLE8mjD5Zi2SeHLEB9SX0LgTIuJ2xXaVTaBGiwQYFFAg0jJ5JmbYw0knZv
1iZPelULjaiDM5H5llrKDP6t2/aPX2/xd0ZuzHgcWr3G8YyENgDMcJ01oDEIwTBx
HvhkY4k5SAjzUYAlua8/fJuwEnIYfHrNz42Z57GtB9It1yYDMyFHW2K3+15B0jwi
8XpjdsmTzEP1DYDCSeP15vtbTwa50mWtQV+x1dBwkcOvSXiX5AQ+LiRyatcGEtfW
YDj+q1VwB+nDtZyl8vqROYnnS65gDHWUDtzPy7MjRISA0L9towQjFdUcolqU2SE1
7PIutjMk4vpN8h71hA5Zk6w1WCi0ioFepbSXDC+lQ4JDfY7eRUshl181V2oc9T5i
tAWZmZjLxPki3hS6hTlkYGcJPyrt0aJktaNrYPBeLOAh0EfBrJ/yKd+iWB6Her4Z
7MsKblfzEXyTDR8yzITBrE+B04optmkxkiJWaf28EZfN4jkLrfB0R7JcybkZMYB9
FF+7ljPAtbtk4DZlVo/C7VgONk6otoFm7CYJjQD09TLx0Ystm64sLdeqiNlMl6+D
YeXvqH+Ib1KAuJpNej1lohGSkGODsq538kjb9hMst1FkG4VAGAyRRUP69uBP9TBm
oLXKWke9cjSsr5XjC+LkyjAnCBL12pUZqF1/jZ6WlyGcKRrVNLlR+iOzw6pvDLbf
7dBX/a7P3isbvQNJkEyQBPbjYoFPqsSYDPRYOO0l5BgwggP2pOu2zwqrrHEUcJJ5
osfJsUmZd1k5rD1wZSbJEL93Yog99CmBOi/8ZX3iQtf4vO94p7DO3cTSwRlflTr/
S6SRP0D5WNUAzUg64VIST3BjafGHd3ZzYG3RUQJR8s8It6rbFslG2gkg7Ht/hESB
oodTHT8GoOALIgfk3eBNbN2waFOHSVSOEFZv1Sm2AqpgEzU1zvAafhDIpoWvXUJR
cP2DmdTrv7+XeQA1aS3ryW4pbksoj4tqrFS8onT39mo4obHZ/qA9a0GoEcXuKajc
UR6AmJwMud0g0Js/Jl931a1utRE3xOMFyu/KTBf6pktWNHdEgpUuprctEr28TUOD
HnuMaEeehBH/JiGQVEyBFKDp3JoDj5AuhdKDb7333oonfFoIz0ln0yQUSihUEDRQ
H2H/K8vzqOWpSv1s15o4N2yt1NcwMlsnPPanSKcBzQIYoxh/hv27GrRdL0thhGLY
gyR778f6a4x7icIdESVVMdolC+6MRjQNMKY7AZyMRmDjdhcPa7JuMxcaoyRIvxPZ
5bDA/ZvbFiGAIAVH0W7hSZQ5KuY0JkoHLrlrq4mN6iDB4pQBGqGdPJZTEXvjshUv
RbTPCYQ/yh009q96ag6G/0/IbaZ/P99QzukP7JZV+KrWm9YcZnv4WDR3FrBtMgcZ
gCpLIKkMF4beTCW8p2T6o90g7nYPsQ/ALQsk1bYRvyUSL+AaSovlyAgRybfMzH/4
y71hLGRewFvU/cUVX56pgykxAVG8FeXRAPpffiTQO+30NCXtBC2Q9GaNpap9thPA
ozbq9t/9zgPqtnThBEScQDd6VBePEQVwftQ/DNNxymq/ZFBwvP+YG8E40yi7nitV
U5WueXwfWmGq387rmKxQRICljVIhPnI7AwpPevsFQSfa2OUjJ3+9SV5RC6jsmMG9
ZBE8ZycFVpviRuhFsPGx/ry9eXRx82rfMwvjS+BIJRtFKJW7ksXaWN58QEPdUino
Poj33AWctb2VBcI2pT4Awu96tp+/9t36g4xiSpearsrrlQCkXyW21Y1P8sBjfC3A
i55utXb5tP6xsSoymEqXM1nMi+kjwGOj/wTvo4q/MACKzynllSHdv6/pbYWB2Uh9
NpiTkCXrupuiRRNOu6IHDZwDpm1IitOvJFjzWtM+AJDT1GfIAw1L8bDCosy9fAyR
1jWtVNrMagJ7gf8cTpULM+l9SN6lUUfP35VcfmLjUYPuOiWyChXOOSuiDNNA/HbY
IEL0Xyqu3cWUsYoZYlvbRrhGZY7AyHo+UM/npiV0grpb+1EUM/sIisr3EtmPUTuS
8+S3eAzDLFZ5WAyqAgaUfIHAGLu6JrCZy/rzN/X5PPuz8mhzZZqNq4yQrw6K9DOL
KFs/Q8Zzwg8ShD9Rwh03hBayr1OaHrlULM7r2H8VdxZBc0Tdz9xq+/DFyveNTm2f
3rK90FTSSAPvvxdKXpMgHjGgAgWgmtObd8pDjXeCFBobCQbazoUtzVYXwzV67Pbu
ys24vfspzcj+IzVA819q1CQKR8EAR6te7YdORNQk3F/0FMvKM+uiv068H1Hwq5iv
3VbFVm2fZWC0JM4RvB4uHh/jemQjftBFXNRzn2aV6AXxjDRB5t2ZgfoIinWezBts
pKHZIX99LtJ75Lf7PsHDRsNhLkhNiFlp44mdirNhBy90w1rbDMoZlwETpyUzAq8Z
Buht1to9MDWr2IoH45mbDgcodNk8FVH+kjpKwrexs5+t0lQ/JS/wY8Z+KAY/4cgD
iZXzDZ+ZdUZTG0lRp13DFw6MABsKvze9dK8JahuEvSAhh6PykF6PX7oXrYWTvHhS
tG5mUJzTDcKRTckrjfUB7C8qlCtHJcBjltkk0Rhxipw24x+vhQ4O0oEue1tLpanH
PWAYM2ww52PDDtd3s5+g4IA5aEFLvwTLMJNZ3sxvqT3+/NbNK3FVhuYIxAMUgaO1
zyV5Qz7zPEQO+DbAsm1Ou6291a5mf5EbkCu7diIEFP5fqMy6RBNKQxRl1LcSAc4S
jEhcacTKRax2FXCEk8wDVxRJK5lbBakOl9kxJW9aj07BsNOKqVMVfPAuLM+Oyw7N
4nxmkm+SyLA/gHrr7Zw97kgs/+3KTC9SDHpkIj6VWxH104Cvbpo7NOVLwQ7ikWYd
MhCUnq1sQdrgB5al+jDDf5HJ8bP2dFwGGMcwrdrRkG5CJsBPL1ZVIQMYeTWKrcys
gQ2Kf5nbbJ6W9xRUJ3qUW+WBEtyHQwCCa1tj175zxwIjiJW5AOhhHqKIeCuGvswH
ZC6AJ3ZHaMzk9i1NMropS8v0osD/CCp1iaS9Pvh16J0nQIREIR6hyetCDVnKAmHq
yO0P/WCmmcymGRMn27Mq6C6xoRjAcYKjE65FSD1iObRQjz36QsuizQAlmAFzDU9l
nmf2+ZEUgA8b058xAQI0CcgQ7coBJu6zTDxOqeYHkw4XQwwYa/Niy4ioGzjVf2dR
yJufO2jfm3BHxRCJXD+/gYPC1oEC3gTtGQq/zYHEpLow8pZWcQ5jQ48vFWV00xnb
FdfPFnriT6H+7A0tODvO4sm548VoZLy9xh8VeHWtzKUdYG2Uv8rML7hIWwan9aL9
639/YTjyRpiW53H0OEiDtMypJWOdJqYLuatiXOVdpuGHKoMso2UDAH35xTGw80B6
xz3JLZS9amiE7CEpHxyVAgmdaT5rvEM8K6YOkf7fH6hCwZL68GO3wIRzd09JF5Fm
HqQTRInavGr1Fm2cs4bGmUmcBm5i9q62TqQvAzGcSDJka8U7Rl5flUtG0dDrBuJl
qZQm5c1YyJrcNllG0JtbBa3AccBOXFTtbEgoGSIeogCzt6R5uukyiscJXrUwqwKu
GfQpVaOiUm8Lqlwwtau4i4S0kggRhJNI2GRmn1MLrByitgLUt4hfbK3OonqFupqf
ye2rCp5e63aiK00Tk6BLEpK7DjSPh8FL3D49t3uY8/j5G7yGTriBKvNbZtauQBo2
KY/UgNbjAme2rFahptlPQyMzw0l8qIsHu9iiKYeDLRPkQEzKEFuKcIgpwA/F1h9P
qpXvxVibV/x3+Bfqmc/RhDkQcvvxtMKvID7sZNB1vN6AB+Xpua7Znrd4S4QZ6OF0
fDrXwhxc1+FseMWG2z3EaqneI5Ys7QF90QehRKaidy0WP29chZnXMosY0FFMt1hN
1KZbJCuZnWYJu0AB90SYkN+n+lwLzcSWP1Ql/C1cOvB1SujRdF135ASOXowTG32m
cg49sictj9OVVsfiBU4mW0iFmQilwUpRl1V/O2nJk/FIiWmbbTay0Ebj0YEZrJPH
YOmy2NV0URWJgUyuVCBdgwEoF9TfLc+a+Xfk7qeQ9tHFWbwchlmt5bth8jsfL7jF
Y5cuzK8g7fcY2qmCVcR2ZnfkCZ3VsSFPMChQLF6UFvtku4n4qu0B4fC9EzvMVJX2
91T41jRmTEHtZ/WVAbEX1lOOUP/ZEm01UGoYuleepqy73waaIum0Twt7WnFBCBEK
i2N/e6tRgbOOjBqEgOjggEju8AvAa45vTbAKrTzVyxRX+VrAmP9xwT0OMp4JmBxs
jUw5HyBO2s7KDXxeVI7K5N6DbtT7IqLld/EK5H0eRzwoi6zeSPcQQLwxsBq1jmLK
sn7EBIJYDRaAlH/XULydLZMUvPCt8pXdFX+u+847YOIGDd4txVJUZDQv7FF2WvLo
OsFF0EN6nyyhRy60wTAhkMlrnuXBUzbG/KL1EMYK/pWx6S4qc/eFlTOM347ZLbUy
gq0M0lxUgmsXFH7e2I2C4pZbtyDznAkFN4rrItxfGz5/g58ECJruhZz1VBuIdi8J
4YVrPyW4htIZ7+5esvV9wneA1jjWBT+7d1nhFACX73LV2NWc+jdgbk0lzn1OZe1L
ewSzq1TkP+0TGOZAX6XevZSH0nE1eDKcoQkaw5UndVrBnsHauu5ZqP3DLh4AqLcd
F+GEiatnnkbmHzjniLd5UmYOfWSPtCiWEdur5zjcCm5bxOUMEgchbQN0Y9iEj5KH
9a/YqhLPm6/VuqMhgd3DURBClOJuYArMYzKbTJ66yH9sfEHIk7NnAAdiKj180X1p
k0JJdmdsx9UUyLV5B+KtCBKhdK+kU81+xsPoK11SJ0ZyGd5Nql0OoRFtMMr9Qwe/
jJzw+W5/PjMSacYEE5U9AI7p+Ddmu4rXRQSSYtYal6JJog0cNG4rSfGrNiaifmAP
yMp37J3p9bXi7vmdRphjXvGlm8WweVXxsDq+9skQMQFIwvGAb5rvD0TI4R3e07uB
a3nk65DM1RoHgspDA1/ruleNhDnptXLQ54CxXpfIindFbdsVjn+M/5Xw6Dg2wkp0
piRSvG+VzB8wLiAoV+ENJyaNe9svAsgM2JoIYF++WKQPuXltDDO0ybO2Ru6DUeDx
9fkFYKZFCdFS0y/I4zUVwIjKi+e1EZ+VBa5uOtAWuzKzYdP5Z0eqXQsuGek5IyNA
FqQfUob1H64Jfa0Xa9yekSUlEhMtwQ5Tnzb2JOCULNUmOxEBaYhgJsHYPdwcBO7/
iGl4cc56JcdpFNcKfSYJSvFwLNjYKVGii+Wb+bSn2NDz74VcP5biAbLQbxTD8DIB
j4qJtpb751BiwLsMjC/p0xt+C3qx/QfH6WE9PtyKRJt1v7QE0Bv3GF21GvkYIiGA
mTy6+WWRbLHRNntEzF/bE8LccRAq+XYRMhImtUGZB+VEAWHIqJmwqPqf4ObcrAag
Gf10ATXevYeALXzjNm0hnx/Q1ZoBjtPLMFG1bYRTpEp17AeriYPgXn0Cc3N4pisE
5FH7KlmwtxAd8gBzJKoipcoSVf8nagEcQW+16faX5Iv8+KA7RwlvBCGkbTIoTRKj
jqRo3RBaZzb7gPYvhWmiJn+ckv7LqXOlncSbrZ6oEBjB2gSlkgsNUZ+qwAxgZU9E
nAZ6mSYApSXl+8qxztjKfwIe+FIBnwYBCHZi/o2Zx/QpkLZrTBz8/WLMOZlqGvE/
1dWwgFt3nU/gZmkPQfqkh8jOkPEQnlu0GbTee2jOVdiWKaWHGLiiVI/Q55hy+BOz
f9hpylHk+P6glqjqTL98yN5IrIPnpWzI236Srrq7Z4Av38Hf4riVvG8vN3Zjx6n+
hS+Qbk0RxsBKe4aUBr/9QZxZnm2HUtENyBx8JxnB1JxHE3h+7hhXDiwwmDi2ucTw
RlkvsKR8HeZfZIgUnop/WEHjxXDpIVxKObmPrpCmcubYaUEXKzQr+QLqrUSLsKDk
tK3JAslKNbB8I4EPYOl11oIPspOu54wsURxtRs2O81js5mj+DG9oDTJM3FLmF3+L
CwPr0n1KRv4Q4/TLfw4v0L6yFQfqDZlN8nZjMbj4+WrzQd7KUySDGMGSU79WTD4A
GQDy0Q99PlF58MQZsv5XACzFkfrVwxw7wkCRFCQ+ReMFl8Dp+p3re0W3xOejt4hF
bszIp/i2+Koe0zo+YzpYGMJ1IA31bavvhNgHc4SRrSSpgmD5n5NOe19aNJZEU4YH
6378Jei7T4opWQcS15/J2LUfRBvlhwtwu3W3t2ZDboD5M2IZiK8IAMGkVY0sz3QE
5IPtSfD5MKYtQwcNf+dkFsmb80ZZJAfEF5cYW347u68w36egroMgZzUrqWViZh99
Y2MxD3zC6hHQvTNEaBLegNKVq9ZTFhxIv7YmkBVE4ldTx62hIH9yAWD3Ue/uLVwa
FJC27GUTCTbklA1Icj0iuZ4tiMpu9Ur65zIdKBO70ZQs7Ifb1V7W5O28Mw6MKHtq
UnKM3F8qVPS0YBS2Fg5e3s7e3zWVp0aBaX+9E445/A5nZo35Mxo4GlTe6yRRUr1F
OrBT+7GiR0g9j3GLH3U61oGJMEPgo+IvHK6SRYs0UOnlWzr8sCteeWvgL+CjgJAH
55xYjBNkAdNDhYHMZsQyYjDU7GemA6U9x+1Dchd6+d2UKOSkZ4EKEs6cA8/eMv1E
SLQY5ZWq41Pm+TpX0Wjcl6qR3ccUuFWpt/rA8mNwZPImQKU2JGapzWWffXGUOxGO
AN1IJ5QM4Ut+WaFYzmZJthNCjXttaB4+8E3bym2xKEa7gJ45KenhrqknSgzE56BQ
6go7DyLh2brRK0JrmMmnldVWB4720BDrYHtpH+JIL1LKBNUU5JI34tFhCjem8e1k
9DxSCUmdHulyJRIwxoqgvJDoPhLPoGfLtYYZfcPWcsRppLQwrqk2lwcOff0PumtK
JeHYoQWGCGSDkUsykA0aQHKj1+lvyiGb3nHJbHgIzhFB10WQ8zJ9gulWWwlBsojq
w406bMFIqklPNdt0Vid8QbGz8U9YEIB/7xbk9MDQXlH/nMKhkbZDw+cGepnVJ0wb
S8tZeYtkuzNG5osQJjS5GntbDOXtYggp7NFD4GSsEdP97alaEuYTz1hzsUtoXp0t
ywa2T+15xTnGE8kLPiI2OUlkrrITVcMffsrZovSDgk4qloESrE/aV+Y5jj1drODo
LTJtVib+3uuI21+lcwPv6mhuElnMJj+GyWSdglqEXQkUIv1fjpmS68iR1nrU05Lc
h6T5FYXBM+dGHIzTBA5F3EbvFD7EKL4DzU7OPTLQRwNW8YYPAt0V8N4kWw8VTKJl
OoPFEmnMBnbCvXsbTvb4wMd99I5exkYTGK/hniNFVyhy6uvlPAbryuzmO5nu5B0b
RZwNJY/qVwrNWzZFn716HevAxkvmXaiXUtGRao4KlHDPlpA9DOiHQp7MLaROEDj+
PYFOrG2FFbaNyHq0/Wjt+Y+AKkM/u92Fib+5nLNVXDb2ssWXM9E3we77VmXDr5lQ
JZA53yew+w579Q5ZjwIzz7wO+NgjMOMGnOiB7kYdyleQEj3UedpaTXZhSqIOBz/O
jgixk22qhpQpVhJObdrcGKDmLhjNcFrphcGgU5qEyzzVKIe+luSe6009XUZKscLa
1UrDw618vaT2InpsrsuSEWSrQhe7yrXhzi/HkwN2lbNY0EF4YMxW36tIJHhDosGo
aKf4VLfxd92FwxJLBeef5G6FpTlKITRt2iJ+EmwbjvT7s/Dy/jnW6zmmfNof2jXs
6GtlesBherdQzEH8m0S92rhk2TAfAxVpPYe/mSwgexC9szblqZeF74jax8GCdry2
WTCvFI8PWBvhfFLy/BzaxLXvxXIGS8Vezq4eAShvCzDHMhkKLp1OTFwQ0f2BhyKb
TXwtUbY4h3UkxWdd2YCIW/v3R35uubBnC4eBallHXdSeh7ioO3xS1npINcgFikeJ
9mViluxks3eszkApoEsyZ2ZvUR06j6W+5XUAgeh5jXwtEa+I0BkGMThuY0vKsY6P
PQtH3+/YP517XdhWJIDmOFtIT/xL9hjSgN5r8a2N27otYw03UubHR9LfHLHgoTSW
w1N/b7DtikzapH8m4X5MM+fuETuWGl5qIF4lk4spOMMr2OnusVP95j8vvEsdCucK
qVghdEU1daScsWM1YUhIZ4s+F4+Yd3uzy8FmWEZeAZ9LB+XOjNUP1sge4PWnOiqi
BBvNvnhltMbzcuhbWazxOQ/z9asqiY66PA4fIKz8kTM94DxIPzHy+26KzrixrTeT
g+ZONt8T2g1x5gQqmO6VhDZEFTAngruBbef68Z/pT4yZLj65EqamcsPYdDigu0nx
Pdjd0xWEnTiosXZB71T7h8Q2J5bhHQpMrF9BfVH1oZB9nwRVpP93YcyblK0Mt0tr
2XxKux9Y3o5407pJzWRF+gezuewy6hVvxKdRaffes46pnx5odFViV2J6wF4e2sUR
w2OU8bppO4GgRZaG4BdBAtm2A2n8bn3HUMCyH0yZOGtXhQycAAkoSnHOCQpgz1P6
vFjpmGX0/ni6IRrsl0NjO2yRIZTawY6nC3ZIP2dCM1zazbcCkZ1vaAyr/5ijrOhN
RR95lX0qGtGQf9A5RXVbH8XtHoT3rlVNmlOSASxaL2tTAVNVuea1YlijPAbw/lfP
BsAHKv/pmroroUYLfGr3EF3Ys7BLieGWSFwYYmrA+hRru+a66T5eefNY1Zrn3KsA
ycf165vr4k4ds5OQXzvXttsWQRj6MC3eAdKJzivs4MPeiDJ9B5GVT03ujV+/01Hb
jIBW15fIdl4mKceqvX7An2v6R+GLKcKMBqyuBGpAKhDryOPzLt98eIsEuRgiX+t5
tV1uSr6OMkC8bE6TPWAI1wxJy5/6vUirthPqDibuiPpTPSKahYTKnsXPtd/eal66
Gi8qSDHgplp9VP5VrDDxuSPT4zI4ILmbh0X0agO+dKm+SiMalpmjdfKjuilTF9lK
pD7EwCmaw9qDW199JAmHSK8JrseYv1GhvYMBLfV0wTwOahWFHPbfEj3ErjUi1slY
cXX1tT3mDCWS96W+DDEtpkpfK6eW4+ezp0ZxgnwmPmc94tTObebrMJ3TX3b23Pfe
PhRhfvQ3CX/Lz30x+ByvseWYnCC6U4WXsM37IYtZMaOnKkHwov/AplAnrbrLXRd4
TUvI7G5DBEntIrcRAPQIMWN2jGMI4LYKVdPChyKoQ1qLuMcND4JordrtjhrgveU8
kqFIWUjnJDqTEbk0wAvGyJvi1VBG+LWCdXGk6juTowH6XfVRWWo2CGEg4wvBnqV5
MXuUzTn8HcGnxk+QQLI1z7O0hpn48brlGb+m8G9lBcD4ziiddQteI0C8EXbvM5WS
Vi5qXNuVOpZ+d63V2/XtnKt0873SmtMLCRf6rF+Yelg+aqoYEspRwIH3tjm4mrf0
dpKcIUjCL+1dMyYate8vvUwheUP2uEKMM76phYw1gTyTJaIa9fj80u+5JE23YcPl
P+ZnCSHVVWPSXsK7XZT4dvQmvSzbyszM6L/gGMC+uLw7eDlqQlZJ/asXnURL9+Tw
bqpX1NeiV78Jxpe1Btm4r0jzri6eHEYit+1G6yL2UFuBKMNr410c4gVSDpkvT5Cu
cUIbVfwVT4YWCzkE11I/hx7F/x81J07KbCbT7zBT9995adOXjku/+dxjGRXIC/GY
3VIoZRMp4VSdqHwW+WxyoAaAn6PQZIreBg0Uut4I5AiRRcJbwMsLePJgctEaOliE
dr8XQA3FLxnqFdppuCdzqADo5MmdYzeVdL30OaplANk8EVHDRBlII0xbaEx+TQV4
QGBs7gBVbg2aEJJcnmzTy7SmW0W9MTEEldNYM18cvbDR32W9+kk7v8YyehzpMSrV
ZLwVzutefYuSzxOfYIa/eQAk3q7mOkW8U/OT2MMOCOGwnAgGmMDcI2lzbaY1AFOQ
0rodUxf91UCk/PODe/eL2Dzssg0NYjGzgvEMA2b7Zgxu/9MmYU8XHj2R/pcKKiLH
FnhmPA1n8Gmr6Rf2Nw5b69Ps3SlVW+u+LK4rJLmVi8SotqXgsqMwFjN3EB/CBJs9
Mpc6erJmR7iuZOMC9oVbxqLXqwRg6rWHBfgRjOGO6v0fD7eYYMOb8JASzaqJIb1p
3Y+QmDaJfeyz+Gk7ujucvDF3UVqehbD52f7/Ng4e3oHVIcO5onSvIXdcN/jMgr9N
7VnrFUpDD+l023ZJYnzsswMkNLlsBanOyxIyTPA6+aQCYitLezAIxuNNsbcrKNzw
Z0LVZLPEBBrgCXPanXR1yyeMG5AhbLWybv0ktWtfWKsFAQHIVJfNiEXJozakgnBO
/ntXEaoqSf50CycgsqziuIwYw8tct8OVNBtNQUUpb2OpPhWLCcEDjpv2XxfMXlyp
rbR7uvvG3AuZY+t8dUojIChAltQCXfhyY1l4ceWlbLw9C35aAZ7aRDumTQ4kThZa
d5cIxswHXFxtyQpRMAIFQWcf+2Xx7I2jxAzX13sxeVwxiw1IWti/N+/KtVkdjyRX
Vutk6L/A5MapU6brOsHSlze2yEfreFoSON0AEFzAWcBbS1h0YQjokNB3NP5Ggko0
YsZMyQRUMT7ELKo0fP5UBT55LyIkYvptuos62cEYon6+vDEoH4ox+Qq7jvzUPosq
/UJvi9CZ7iakYOkLhyNl7f09bfp6ciZN/vcQ5V5FdTsc2ulqxDuZlscDtvqTS1ZN
JbIiZXIwpvkrlaEez4QoU10YWDIM73izBuZmmvBtg/nsvQQensNoqsyNYwFiMEdf
Rjcd90z9bAI0VwRrzVXLz/Uip4GFGZI4oUQpvxhqhcEYyADCOXZCLFXclWyQpe6o
iOpdc0PcCUFWczHvDeyJYUuh3SAWLXGoQ/alSNAiiLoKVdQs0DJvy60e84C+wYcS
TZ2UGS9OizujnSScUhhK8AHofZ9ziZsBYAZaA0ZCC0VpcM+6oy+U552LUVGlKSqP
lkiW94n43VfIYJTTNbcNkygwdNPhKxcNxZ7EXrhNw6CwavFw9AkxZN4hVHu5J6Pp
rBYcFIrOcP83wHi7o+MBlf43rvKVCjW/rQgxFciSpYxHQJit7cIMtZtht5qfDh+o
2i7EZiZ0//P0NkmE+wr/7GrgavARERhRs5cj5Rg4S9K6kR+wOBe4pYEeeSxuXaUC
FjvpG1eb5N2TKGu91kjn/pbao4kl4J9V3vDotkiMBwfNbM4IKRpFU4rwGpnW6ETb
s/Vq/srEIYpOJg0qCChnPbB6aUgA/S3CehtbFAm99gDoTssTGF1FqnkQw/HA+KIN
GxWFK/NYsBzukyimjLGBoYNu4G/dBSmp5vLAoIaIGNRTZHA4+a6n+98v2DeLBFc6
a2uLmGUhbIH+QON9aK+8tOVrevx3OMYdq6zy+SG8ZH/5oW4QoZaJ+lmfHj9I138M
kwgHG5Y3Lq0LPjCkLUfTezpvxbiak3ir6mdBUesxCrp/l4TdrOMyb1EpjApTyvg/
uf2cqUxt/+bNK1mivNCOsxpkES0DohV6KCgdYWlm3aiMU8b85uQEoAHKSbcpOKuy
hFRGFZLIkMARAdkZRGFksBSRzE54WkMRtY2gctbcruqFE+pRhmAWhh3z2F2mvLem
u+OtP0/Ow5seNkBCefd20QUG8ZyqB4cmC9dhVkB70uP5EAQBtlQxQ5qWVOprKMG9
gU1e4IZm00ZIvRNmOMveuZZNH75fSXHsh1xEfuaqJIydgTDRwGNlYrCpSQ8y6p3b
q6jloa1/8pY+AsMMfP9ERxlnqB0Uax8J3KbWGk9lr829aFnPHkKAz4eUBdbHvVKN
lMr2cihN9LWHMylKo7ueniD7EBJ1otGCVOfMLZBGLk28jGPbT6P5y+T3MNWZuWgr
KfJ9utBjj3IIMdKAuPXcvI1OPXOfi8YGcD17DFuqbK+mNXLkgntKfDU0E7t9a4hp
BqM0jM3uSe2uhGb63lEpC4bY+FTm7WgIJFRTyuHFddnq9+DeAka4jrV9lcki7/aC
Kt0QkEZu7sK105nir0WAUzshG08w5Aa2FXnntch8GjllzCKnlUFSsd2VamnXhL7s
g6Hi6SQVyVSbcFp9lgREJsOEg3FfKD2q6K3vHwcZs+kPkBVb0WZGg51v6kB5ZcFy
DpUBnP6/+2BSOzWma2u5zTCwppE3GDDaMbK+0IsdcviPsLXh6c/7aosGVnTmjNqc
c4Ty7H4vGtB1WB7F8F8c9AdjMZT1eQNNEEnsODxMgvxXCpk1FdPJX15ifJ9VwPwV
SrM3pX9xhUG8QvWu8i1Q+aCA2+JDA2VZ5y9E+rXdoBEqQUccxKNiJoIQHraYlqy/
eihXBzTOJPdzIiC9Fj6fKc9XoQ6t0Jic3PgyBsdzok3Uu84W5oM/2ptEORavvgyJ
vGmmtHUKDxbZjfM1or4dNwFGT++STkFQCQPLGyW4FM3eJZE0zqNyw/LHFRt4GeV5
fR9I4FoeFYgqRITmDPH41a0d4v19ZnMZeDJBrktMwPA+4GTlB0ddz367+NlIpkVJ
aQf6XWnSqqgoEeWpWUO0gYTruo5k559xjTMLlD6VoToMVP54qyWlvOi5jtgltshp
PtkqO04gbdIor892woPMdeK95w66EEAYItQlT3r0HYRtlra+M3p3mW8cjwWfR9k6
T8eF2CoxV9B8GeqMDfJEDF9Rp4iyXGXJnlzvQTmJWKfZYiWtzn0vHC0MKetQHfYI
KghrvL1Ipnwpn96MyhUGnc0uCBNWAjs50GJ9o8I3jldAN9wGXgMbkCwQmktmlgqV
W6yrx/4QsMkqXKiishUNwqWva9k9b/Mlb56fhUSEH+YO+Z+60oxBG/V0ibic/loq
1kcSn/EHsmOWfthkaKMzAH/WnKArchFYzmvVzL5kbRaIPvXtMw8syrBU5+0ixSbW
qOlkKZ5GNhdpTZDOW1quJbaK3uKn1trUzlyhjWdnE7BQgC8QHwfDIUoLygFkiBFJ
cM4VQZ/8Rf4SUrKKOMdaIlnh+NxA70GpACAfHiyWKQ4bPeDXjvYwtoP1z55C3fID
VBrIM7E4VTYWlg48pqMN5qMvlTFeJiZhWUv2plWef0KtJGyM/o4VwhwMhk8tfjyz
ttycOYNdHhfweRsxeltnsiuvhJyTIdjafpTYKWQ5J0SKnND4G9BO+cM5hyy7eC/U
dyYFMK91LhRsC+EdSSGDODjf4JksAToy0LoYiIwkyTAiY6Tazv93CuGhCTa0BOHS
Wc3Z2nufuIF+BRKx7OfwEgWYsr65Ili3KF2o1ZNSvP8pRtMapgyrrCJvc8tCDNqU
7mV/q3PD4iIZfzzf7QqRun+H7qSBBuT+qRxyaWV8NAVfKkBzsnBRoTEoymjN7qtr
vQYyIPzXx5fnCqP46tp/eg5s6A3ODdN40nqxR8U1YkZuGKxD9le3hFpm4Aw0fGwY
uH9r/ZnBCZQbQP08PY7HuSDzxvqeeaxkZ4j5jeQ9JimLbt8I9nsx8j5NiELkk3xY
r3cA0A5ZushoaEcbVEmX5qQG3jDe2mxhyWb3s55IcDOEjZ/0USW3dwRFZ9MFNAfC
vu09YdmdqjR5bg3V/nYTJXfeNQuf4Q+CGsKAnw+XyDzMjR9PhotbjntHtw1ik9ku
BBYrmqq7soNHTStx62f8Iwl70GiHXHa+XzMMFihUzLU471XKSuk+Qe0bqwvdD7Am
C0jhnRDJ1wagfBf/MHzRrOIIuyzteFMZV+03wG6aE+gZIPeZha9fjLvMFWYadY3K
kV8ulG1DcH6T6+VDz4t39uumLMLwm1059Ysdvl+1Ug2/Qn1F5e8b4Ur1my71b7mh
v2BhRJDaoGBSL9jPzXKg1BSGsUUq+Itz/jG3qo59y4UJoxJtIIm7HJXFKy0Y4YwW
IJtzLFIv3ctlTiydCDTmoUYgXnjTGN62Tpl6fCNWMt7E3KnAEj0MzbSix8K/FFeG
T2b7hhf3deVlyuZ1Te26J2xdwccsVspzk/9wjCuwnczeUcR4J4RmirftsjNcdfnI
Q5FVHoTc3F6y4yz73aEW2MAvCHGaLy2efcnhXZTPdYjGCwSsLRMHHr2IVhE72FDC
o8EqUz/AbVtDJCk6FBN30hg5yFYoQIYockRt1bRPoSSIdeUEEYGSnv9gyBK200Fg
ZnmfAol2dkSE3wTVHcjj36gbQ+aMRKxQJBDez5BVpRV8G8AtZqWWiq3ikAktnFA2
vyOym9ZDAZx12AR2l9HIp7N9LirRvdfFc/cjPAQAZGK0OEjwLUF47yU5TxcnKUup
oPz2w1CKmWYuH6kRAs17ewzb9L+hVpXXCqT8lt46qgXevw8FFLvoLQqALVJrt7vL
nMzBeibnr/e5uaIRHG6zRhksRpKHetd/Ffak9EKta6x/y+eVGHxZyZeVDDJnJFit
sWB31+w0NXWzTvqCX6KDFQcB62ywGciLXCf2ua/YBsbUXAa5rOPxu4VAAFVoWnTK
J/VFmtZf173qWFn6izTgCfw5vnk9Z/HsdDfuvMrm7ERFjrCfhgTWrX67dh7XANhc
VfFemmTOQRIg8YvNpeMcZRC2OLxmDvOeLqO8pwF9y7MXKj3YMa2h+0qs7Mz67WnJ
KpNWIJuiGZREOA7xAeOFogy53wDcZRrebS6+2EYNhhnsekalTWSE0gm5CiFkw8uA
0LlGpZvZIJzsLv14g6e4ZY2ywO/cHPK3vKZChtROVtqDCoTH/1K2M9mX7+FTSXqR
GduSKq9toNUq/xKWaxkLHgBSv/bwHHRA2LGOACofDIPdHSknFxK7AL2pdEsCkois
gKodP7EKqxGBVWKuo5Zg8JM1QbFcgph7W/5uA8oLXVBRCFWqD2NyFlSXTcsVTB2e
WnaAHjQNfezR2xe57oXnb5CXKBqvlnohF36DcuhECiIJFwJFIItAZ+7vMNtLOLxE
iwUxHkH9I8NnOuw7gWVi5397eP1QNEm/+2rJ8+QUydqW2TJecVMfTtDGVM5Qhsqp
2vneMEinaQBqqYjNxFYVqX9zIpUf71qTpdjhFjXqYL6+aaoMy9QEIWhhsL7Wc6yA
nrAh9GEFJSn56eGMDmMlb7k62gZ0sj47OCMd+BCZ+S+zgmcpCTcUEj8tWEP/X+SO
8gdLUAwJgTpDCHNQxczTX6zrWWkd1p4XDxmez1BKh5AIiWKpAgKk4rKxEcDm07lZ
eZCSZI7zydFvhzBfJzC4NnGyQxOeDDNO/rn9AMdNtlm91TJlB70aiVrFaUDLxpb8
CpBLgLwdo/APdYjXpcUqZ94U5SbdAjtY0sOfARkBpm3MvN62WSQbg4s83fY4ZT9m
+BosNen7b2jRoOjdEiLbby/401Nzf80F7xUsCk0PxxubsjbJqr+42e+Iow+o70lz
ucZpRr6m5Mj8IWQWmfFBvn7MGL0miXBCkoECa930YLquO8SWE2J8Q6nUbr2ELyND
xCYuU1GVo+WrySZ3/Z8hvso7RLu3bfrx10LRXotSUUuYhLy3+Vm5n7pfaG6Kd29c
zhUXVg6nIJsiU4sGcOnB+Gmr72OabzIBY7SPI1cxSm8YHuI9z9w9h+o+YbRaHjNB
TEEYOTiM1cES8xjr/QxuOxlpwBghRqMy5UoHOJVJDpviCv+pJ8sJp0Iat4GuTGb1
Ix/t4Ibu96ZE46P7BHSoO6wrVicqFa2D0DL+vuxrYm0EKmjexSLTaSeHPF4qctxy
l6pTy7Lm1KpLQrvj2qgwAFFd/xYLTNpLcZ//ad5vH+qmWRXp/s1bwrrqipqsj5SP
tfh0ABaP7a+rx9LnfGr5HtsB6obPRyCeRfxSg24vxkeL8LNh+hxGTLYm7XxRYXAQ
lMmuPuRoeTi89I8ZgcUR64hUMBo5krs7LIKJuoKPB1u3JO8Su5FR0t3VnUk0jUZw
jLORiPGd6M/V1auV8xe0yZtcr+2AEg6PkUChLWfLapR31FvJx5SD268p1A+hP8ob
qfeSNox5MXQmSP4ZOs36jmhdcspDcsyq0RA2LTnlAour1GnHYej6qmi3Y5O5N0CT
RB8T+KHWJFBK3DD/uA+uUEbY7qBxGWGJ/DD5o+laovRlqSdC08nA0KC+KIm6XuEx
lrJVrBKYbsCTy5hcfDM7VLAmk4+0dlQ+Z/45AOBpPjhCwShvoldgIvCuPqWC0+A+
B6E1+c316sWCYY7t5KuPFuRixjdgZZ85XANYSMova5EPorjg5pu0QmQcPKafTUkE
cCeLd4Fci07KMj+BO/UPOur6x8ayq42tkcLsM5EVTsqGH8RKlrQxw/Toi16aNiTv
GoJDka1kVgHzLMS4i8EIDiw7R2HAerkBaJwDfmgIZg4Aq9Mi6Lug3fmTNsQVzJOE
Wl39rxcAtKPCA75E+MKugCaqgxAB0BqKPcKueQV9R5nCuuDyMh2e3ZEO6o4ejpwB
xSv2EWOloB5CBd6GbMoPui3ZHPUuDScAjC8ebBTkM0VOr6IacX5544EKps/5LvkW
6cWLRHpS6SfT6Cg4YmnWGgAfAu1CdLCRu27096kFuxobbTMeAj6HNwMSD28eTsg/
7o27ZlQYKJo0mbdX29T0cDdI6p1XVU5RM4T/Svky1fl0CqL8JNj1OOo3lJLVgdCc
omgJhnznYDEon2cMDqgRc6nD50nfoYCuRokIBj59HzC+hv3LzVXXgT78llxfgmT1
8hcEzOIemnS5VoU5xaOMwr//MWMiuj7hE7BTTUuKXrMUQ6tqhg/2MEOCIZGjtzUb
ghz7JNXyHIqIndxDvg2LcHUPR/W9pcefthZ5ZucKUpUZPLdDzH5PmKTMnK9Puy2d
R1jZwrPG7/buglfFfUxplt2jNkfQC7zKk5MrrEVYWnGzlP+syVnGbI8OEEdRv7xN
HZuRbKTSbjuU0Gx0fF0McPpDa6ZeH9BCSAbFKHwc9FSa+dg2Vox8ZI1kNEk8PMwo
clhU3eIdDNOapOCul1m2jlMa8Yfv/boPhODWWAbbWc4VuWpCwMdF2kL0blD4j1Fq
YN3BaX3GKRP9bvxqjH+JXkDXoyFVukFB3yFGLbSqmQhPn//7uLQC4sta4HsUj9Si
nELzQGYEJ/CC7C1tW6YH+puis/53R1YO+ZIX8vZ4Roj98RAT3GPRDoWsvXx/LOTd
jNQvrpaehIfaLlp0cI/+giNj33lNgY2HK853fJceeNySEGb5qbteliK4gha0ORyr
+MC8MEuHxC94B/j+rkkkQxFQlSGXX3bXHDEkof6uEe2lSFnvQtUB/IKuSNwv8LqN
4hidAC2RVl8s9A6gU3h5K5EcFx4SBY3a6acJKebTRUm2JYF5FM+VVG0YTVsbeybx
wAKseBVZUp2ysQJkn+oCMwo0Nuh09U6ltL/N+B8hdLphlljFOxSGqI4dOXjyn2Ar
wYyyM+Jv06J/agLII3NCDQMwE0nPnccKVV22bntfslTHAelX708j3Ujqp5QC8Fo7
PfLo98cBNL2JnJCmtdBYwz8JEmfaev0sWob14CJBcaweYgQvwygKZvobu48aGfzS
2Z4a/YL5M3bnj+v5BgFmmFk84wXUgUOXPe+zleRxTxP6M59r1k5g/Rm+s7MrF0CF
HRMzwGZWQQLB76J23KBms3zp/Po+0UHlikOQzkiE7f1P0yQQeq84Rpc5giygniLZ
edfWUCrfXrMMbq42s4c+CAFU86mWITlUO0Tw6FTiImHqrp9ZPZu39wNQGb6bVmri
7Hx83HiLq/kIDSoHz+JZ4AKM42Rs6wlGIXrwTnHBA9PLwZ3wX7kogfjxyYEG0nLI
5mbf1I+HsvOJGlmOcHqGPq5/pgARoCcd2wqePhP1f2I7ksodDoTv0JNq+3QgdF8P
nO7ZdQ2oTC7jvZ/eXxHse9gNqNVmDrvHP3lun60eBf5mXFgZAPWofMTivIHe9oTZ
G3zt+8ELCzopQ+M4YxeJXbqW36tzP5PLTVrc05rFhqYhNlrnOARrPnk1lPic4c6t
ICNHWvuPPYMKO7rCZM8E7C4LqRo0MRpurcJfhrkwkc8+Y60ADCQcGjSGn17ULQ7Z
DyY1my6qdx4jTmdSlcmROohi1gLv7NyRvPvQR0y9bOqD5i5NE5vKcFz/R2nNA24Y
8jJe+QaAAYBU4zRxpzZdC1cWXf8flmm99HHhPvMh9vIsD+g9pOQuwzMuP9DXbr6y
gEZzJDdm/S5py76qifkH4845EAq6LyQzLaG9uV99UGIuabuX7jcH3Gph64IouWPV
OKWH4mQHRGU1BAKkaye+HK+AtjVbpTP56LGnwhl1hHtIdAo2OHyY7UvO+b518s0A
STe6by9f8/0QvDU7OB+A+IucCGwiS1D8+iLDGeUHS3wMBEZXBunD+DNzD2L230Ml
7kc1xsZgZyaB+NOFZ44ALn/O1/+rfehv/piCPWEQbsnh16SRuCalfXAs/yl8IhSE
3Y0zVmZk3PPTiAuzdQ4wwJ+HY/s/jhXBBZmvTEiE+ljEebCDeS/cR0bC2ZzXnjCx
pToz0kKaIf3M48M1r6JX5t41p3CgSV9qHcuNYXfJcJaO856oaKx56VkIBPO0UP9F
ikyTQvBrRHP3vs6qk5pmsmTI8vimWqVtv9xLe1UzdhTCvdRIUhuY5+ximp8Znrdf
SbyqJlm8pfyxbexbneevpi+LQr3zgXNnGSN/vxOnli+RHAr2gOVHsgkVvx9OAU/H
ube/U3wCjPfmnFXH6q0+E22zxrplNFqcYKZAhJ7uX/Heq+/WlFNvMNbqpIwQWUXX
hZSbVuA1QRS9ynU/oEaJ4vipw9jmk2921o+zYcp9d+aFf2LPneULGBQ2I1zwOa8g
aoXT3ZcmOIwzl9Pns31M//YJgLHr1vy1s62MdkfXxFKqlU+U5B4mcnSSVPcwOBZc
sbfN8JEd6zefG1d3+uaOjbKGPo6dG1gui6H+ogofTCfTRzZHeCSg64AfTTEoFamE
JlK9juhXSOLvW+Zx9weqL7K06bjWOx0mmsa9HWfi2FefdCFWvsyTvy+r51hjL7xC
fBTGEYkHu3Ruwdfl9KGj3QoYcA7keAxmInYx4FgoZttDf0Do76PEvsk9mX/QewFO
90OjSsvzmijqOJixEhOUdymbBP2kOc4zpIHQQpdsu/n36SLCHbKfv9jUAjgmpPhM
LOA1vQmKytTLRTvPVT2Che7UI3gR7mcqpKlyIg9LSPmQ5C7HN9/wRVPgVMoHg6Gn
PEYVGZQXmdy2GeyX4g7uOML40F0MtZZ9tXEHeCcnk6c34OHtpsV7xisKgBjVZr/8
H7BNGkwSPDaPe/+jylx/kX3CYZY+ersm6UXD5FbXHzj1EwFQEH4IvOuoOLbW0CPV
o1rKmTeM60ixLrX2RspMdbUFYqdccWkNo5H74prDfEyIvrbMLiZZpQhmydEi1Q++
CCJ5I+puLzuSJOOWhN2D1wIR+Dfrwd06vrjU/8dPXNiCJPFVYK88ud+ySpRCg56+
6498ZrvNGDPBO5UzE+UU3zkw2YdP+ffyTSOm9bqv8rxWf5AYhBuyQZ1gzpiHingP
+hBIPFeY/RFxduroXaPJuSqIvh9OwE+o1xqryvxz3t4kidbTdnvwRueGKPirA7C8
6H+8P6+Owx2TkuRTvcQv1zYp/+mPSZC3jTLvcdT1PUWll1EK4+mBr/8CbLaY7XoK
v3r4xJiUW6n+Wyg4M0sTmwxKzq+KPL4Y6iapvatPWbyctscgFQsAo8vKFJCLbihm
f2rLUgKrOUPAxGZSls01pboGvy4Qifl48TBzxygwLcM3u0+mEgArE9RNuNgqiv2N
kqmHHjuYj4alAxfqIJIV8H87ZSj8ylO8nZ9WAxDaOTeiqqcxfvoFV3VYGp8fNMf0
5lAVwURZ+Z/oxu0QNAFRsW5MBpTJSs1jZA7WlzjjgDrIlljeO0DuFSsFbtKedJUe
IMJD/C8KoHWdESNlkP9kx8nQHOMnSrigmMOBLTCnhPd9srxrgMdGWQ75zZnSGcyy
TpAMlBm6PZallDQgD8JBkLvyTcRGYGXeIQKXOsHr7iJTJt8yPzT3mEp7M9Rvt4xL
coBMxSgOKlArUOf8Jw+5pL6mddgfZISj+dzkrXfbP7STsBgd1S56Mo4On4TvDLhu
g3UNHlULOnJhrHx3vfsFteiVmeVaxVqd4pI/i5jXDsrKNrbGVNlBEf9oJOR8e6FW
39F+9+iRh6XIMPgP+yYM5TDEYJV/kI+PEkwBZdj1CI3v3m4gCvn4Cn9jZHjHFm2x
kB4dyBTl/V0dcLvKG2+O36GMjvBY9bwSOtv9x+CCEnLHOwYoXUrep0hEJ/PI6gSI
L+vJtZGlBIMLqM0g0joGOtdtCdMqjhmOMhnMKlLQ/6aJwbO1FxOUOFLTCuvkNYEu
JBcfpdMn3T9jRzwQEdPCSFFJZO4jNXbG1Qo+m5hxY8rN6dNvokGrVw1P9ifQqCsZ
Zl137K0QiGHmslmD1iyWnAWxZmb3BbCB6tlZmrdOUuYkf8BwsuoaZpcFDnRaGblJ
bOqC4MxRlerAIG1n1IEL2rxQW/3zmbPARHZNHkEIUvivNgBXsFr7LnFQpP523Viv
X+/akFWnUTFE9G6UhetcvSjsMCGlPxqhnA37/4k1VhmE2uz6H3wi0+wtmFBqONv3
gwHZ54k5HTipbCVBtjFLnF4HbpRHO+N5jIG5DhfndBQI6CIL0WFit5KDEJxxmZbw
zINoai/RPqWu5Y76XXXIDF4mrnhGLnHWEMp+IllBfP/5Qe2DF3Bfkc2PTiuJYCOZ
cQ177H1Al+baPN10n54vbqerDP0dMWzFqhQKfT0CEeVZ5B9+jKM6RnytAc/ctfRd
4MGxs9pbKT/WOtSRDAuApR9X0ns3wVwHfDRKeIzwvVD5T6d5MZ9AX450I/it3Ilc
kA/EJ7UUUJuD1i47jWNvtisVCJnomZRRvP91C7wpfm6SkCtYJYjlz+5rG0mtgtGt
DbR2Lw5X8nDS5R8WYzv1+sx9ujMtzCAd8QUkfaCn++bmFQuXzNI86PsqA9Ac3FKO
0SfXse+iev9dMQH4ukipF2F5RIxX+PaB37G4CJwKTLjgdZSHkb87m+jzt4amdIm5
hcn5kGGBIaT49jlfhuXOpq1d6t1/0ZXvWX89X8v7EPJ+Hqs3ubRo1gzzT5Q2YVih
aAWGFDYJr9Myvx7DXz7GYzcbadDOjNWOJOfL6VS9hyfCEYcKeT1Mc0kUHmdTxi4R
YRir5fAXZrMASWZBQQEgcnJxk3/78p8+qhr3qht2pYZCa+0xLBJajLZhTkos8p5A
bFTD1lZ709To3iaB/epCSXjhepbUAIBkx8IHkjaE4aEfO47FKpNTTxy8z48T87U5
bSnQ8MJJrMqEyY1bIqxHC6N1Ljpd0hHwuLpgwPQKoeE9rpN3FL+rdVjzXNwpkA5Q
G7qkWQOpqV7bJ5xll9xzcUgVthorT/6r232OAuFgss49r4hVaKQ2VmPqwqlxTTIT
hcKyQaIQWOAhdMNN9iu+jtJp33WqHt7Frcg3w7UPWuvZEhzDqSiCEw6youQlDEmj
vFTphhkFlH0Jpa+PpdT6XzflRTnDbNzHsFLmv0zK6boBT1TKRHUfbgZCnISQhCt5
P3pBMAROoLXg81e0mPLL94esOKgzcz5WbO5oWKwbmQy79YpBnl1jn1lgotizfPi4
6NZQMWl4gR2dQyxYDxYYcRDYB8dIZlEQwkOJx82e6z+u/3TqKowCEC5PddBJEO/u
rtrY1cAcxbeuo2XPWIpFy2JlwAQWNo+l6XjZCzVIBXSll0vPtfR7Y7ZAA2wZ6yY8
60/xEFdSx9dAxqPYp4CjyXjxMoJKkX3tTh+nMIuQIzHZgpELNK0+gysjhICuX8g+
xNSJUTUz0K8T+G8IOhsOX0P4O6hnvNgGWam4VLTHQtJhdYSp7tBQiOLDUhajSRvh
sWrewzodg1MQ62H2ua2j9y+jB3GnUK+fG3BmRpzxcaT1RvulF2u9RniA3rMp/Uo4
ct+gEcdAjCGJ5NgtxBJGkCQ+XRf+hwpLk028IyDO0GY4T7vIpOgIH8Islh2N30Bs
Zw4KJvNV15JSUhwpK+IERDLAE164S51xcOfem/MvjoRPVY62XaMDR88Llf26B9EZ
Akx22PGD9B9+mCUrWBjIa9JNlsCEdjvGJXtzxJCMHLQSXkIy50Z9Bv7aEJ1OyEII
Se2IPAZe4juZAx+T7xPxRmuPapZ2XTwDjsh8vk4+S2GjWCK4SP6I7Y0XrSuHxoYg
8f9Pm4jl2jQqrRgzdUbq4jPd7d7LyPNLjaSpoOySYQjISFGt5dpzUmUl9R/BeS7j
4fzwdaeDj9V/8D0h3Aq8q4hXUeHNSmpZ1JDQ2sRoHe6L9euw4aqcarjlwkvX+eeV
eLiqeVbNExj5N2zvxIsJ8Rkigdu7xmDENtZndHVaQt84JEMLaqQPNvV/x56EohUn
26Qn3leDXRoclyO/G1eKdxJRiICdNgjWaxBWnwUE99ojA6LTc5oX/paaNTMOjvbf
62An4jSK7WvmHm7xT3xZJTDe0ZHczAAZiSN3qsDIv3fyG+LnZN55LAMgqUTGjfC0
iU0cq5DDkDdNNrpFNGNg3WG5LVogJyiTpeMQnbC3CT7yNssv/BYQtH+T+NMln1Ed
jfCR3nq9Qu7MMcalQspxohsoMWf79OBWHrS501SEOCF0z/IpUbhRsu9ER5w2u4yH
2ROrQhoGIfN63nscUywj2rv1euUO1aqmCghVVQvy36x1R5sOCOYUzeQEZZo1r5yE
rzx8Ddlm1Z+Ww0TI2h0+pohCCd1Rp45LZSbZsA+LUKUVCT4OUU923E/mYwAuuyhD
ZfYP7fiUxtoNL+NhRxmKUFtd0y8DDTs76c+/lVDMT2zbOjVd05sijAdJfaHNbLTv
FPuy6vFBmcKjl0i4icDjRKP9nzklSNfCuImHhh4hWHgo0tq13Db+EwM9uWP87eto
s6v+nbtiZkPhETxLSRs9DZcczVKQd/+NRwKhJKLnxT5yF3BmnKSJK7/Ux9W4ET0q
DDz74CMzLkBOEiZGTiZasrNODep/EiIKE3SdG1I3f88zQPDMoNK/7AQMc0tdvkGn
jOO0HfpRO2PkTUFj1h/9ZlbPD7n6hehUAQOhVSrTZvidMx0G5DcmQqAywhOE72Mw
xWenOF1hq7bLSuWYNMoaYXl1RS22yGHNaqq7J/MMk0t8uPmerhDPHxWqS08fqgHQ
voNqMnmm21mneqFZd1nUIy9qN+mhqdsxx26sWlrwdHuSM37vNMBwR88BiwEPWLaX
7cS3ArQj4T9pfAtPQDMX9ga+EDbnI8xPo28bW4OxBO5Mswr5RDhODqgOPyhDDEkj
ZNl41kP1F159qSRJVcgKyj5dDVwcZXleV4GJpNMHzrpv6Ed4XXNa9CWtHLBmOarG
5WONqru4RC0y550foMmDI+wXMrdNMdM4Z7v1FMFa4yS5I9GxSYjhzVyj79k56RUs
VPE6Z9SWi/akTbu2Ds2bem9sryYQkw8V2+WT/XEEFjayqBxB1k7d3INILDGXG5Fu
RM24PjpOKpXYXtBl4AYb4dvmlV3SqU+a/mQaAivcda+CQpZnn7sL5j2GK2kOzBLe
TqK10JGQQbdu/lQrd/W4KcSpRtIBgjLA9OGqdrSvGblFEJuuCvpHdjXgrn+kpeuO
V8yxCAtst3/YMp3YceOPEnJtYdsN/xyc3H3QMb8kpsqIECJIZninS5RBEdYB252h
v+QhSkoyTrkd5lw2V8naIdXgo/X6wmpfCoBdfdb//kzssq0z/gqZ1b55YTzduUSo
vD9W5mXrDZugGwz1Khb6wdGdnqqEwpVSSVWW48NR7bmmMd211FLyuMmEyZDqEQFr
A/PQg7X7zPzxUkpJl/F0yXgteKeST61SlVOiCkiL2PdmhQLjy427zoM+OiRaeB8l
Ai6iJqu9gp+O2oapKIB713A5YnFrO9Nd3bOZ9GgkbaMQme43nTP6OvS0fJKdn47P
bnaECVx/pxtpexw9N7X3G1f4LYECIAdE6wJvLW0AFr5JwilC1bl0ZK992pc7jXSr
nNDVBIRBVeHOGAa24oH2RElA2h/EXQHzSGehiqiZcPm1183YKjn+0EDfw5trXUD3
UhYr8efaS2loAyF7onvCniG8+2QLyPG2L8+hO8EPuLwWT8z7AUctVH+nSVl0Ghrd
Y9d9lqvkNFpPsveyYOWXeu2T8IQ8uTiIZGE+ESt+GnxCpcca2YunvBbm4LDXXOQM
X8bvH5Hv118T9k0N4LRdxtnHYFeV2D5ESob5H/wJfnoE6idmBjautwJoV+y6xtk7
5e5J7Q/BvYBBzL/e10FrBSc//AJbSSvv4pxmFoDWwRZ6k3JWB5ipqCyYWocdvPjf
iq96xwIRrzyNHahr/VWh5EPJgF9ZtqDs7xeSDIdnbCTjCEdG+ZXnBrGPymLIOKAd
olscwrK0xYwtb+tMuBzkC4fDSonBQeejvzTjMtws4KtPH6hUKmYlOBD9kf4jYlGe
yCgSLoOc5r/pz8XKdWxBuVU9Pro77adsjqSADJdddgCnNj5mMnbtWFbQrwPx/o0r
FAHTqDwNZnC9JQI6yVp9d/RFBLPhzzunUvtP69jQz4DRnKY13bFz+aCcHY/nmHdA
pkpaVc8fE/hgjHZG5g4fmffmTnshDDIFM3yz7hbBGcN87Yg1lxHAtA9g0VHoZ6nG
pFfF0CoTBmT+48LkdjPsITbw/UQzb+wpBimez6six/bWS9oAbZFQPogwPfv4XBSv
JUO7R32tzjyuJ5xTkmYpZPUloUj0ZaxOO0Pw0aZ7ah8khO5bpq3PAz7fsm2hqfD0
lSyiCJQiSVmnvLzWhY8vmRxM4oUW7mWpzG13FlrxaIbA+RUPa+0HsKMKsz7rfAPV
HljiWkSDWqcvH9BHDH5KLEFTRfQOCjBooOlQMu/otQUJf/csSGtZjTIIs8V5f5Xv
jxAiswDp5hwNK79ZFYIA94Xs8uW7VX6EMj9K6E9CxsxZZd+sko+gd1XA4N6dcWN0
RxVEKlQ7Evsk+Fg20j7XPtI5f8H4Uk6vEfyc+SlGnRmZ6P/jofjNzbgpTg3MgCRs
XnHSpLOdMZh0oCqoW1Ntb1oblJ75q+pNl1cCBX9YJxfCSozyDUWASyB5pGmOemyS
h3gDpxhPMeUAryVmLgsVPmUhdnsB3ujfOhaKaa1tHn+V8+ujZi89tHxPpA2kvCiF
f6RSFMFe3p5NvCLa9+XT/Rx/LuPe77BYvJKp5KJVPNqcJMTQM2+XaSZJTrE5DQER
XgbTczi+20Xl2q08k4RyVTUAuiv4PptKoYpY//BfjipO2A8WrfR4R8E3qOb9pcuJ
XEZf1s01duDN4egCtpmtfV4ppMH99wpZ0MmECHQ/IuoQaEE/KPWC65KpNG0Q9A6R
Wm+AxRsxv/lpPR7VuIIYrAeTwNvTGCcxpFCoeRPQzD3Nbu5i3qeDEkyIVt1X8rxc
R7mHxX7WZuTF/oPMHxuhJ5G+TdeWjfffJOMuBe90QZIjpRtyTpq0iJ+wlzg18uFI
rTkT8Ger1dPaewoIWqK1tbmLIqHnE7+hJCjKO8bh00tzclBRJbHiRUQrqf71Oakb
9KQAWVor5XofZN8rb8wHnDt2CHyYKb4qBJhTktixC29hHlftoAaSzjWheD5kcNUQ
U2CBy/arJ7LQEAkj2iXfeXpgP/uE+xMkt8jRZmIZLzrMaKd5OCgmfdflSTrt4kY8
/kh+2eWtLkf8qkQfruZXtsNROXfmYyO8/6kFGHa/wk31MkxEI4F4uXUo1+acAlGy
n4VaQs4womkxELI91MXUIfLejx316du7qMjs6JCDeD6Wz8R0EXy5ZiE05W9bBJ3w
tec1n8pOHADaK8BxF0ReICFoJd+gNKxMPQTL/M1znpyAnaX5/Av5PJ6HC6kCQJTv
CoclSsyuH+suGIK5INSazTa22k2maRXpACSXageFq0ezcSOO9oGbucJksgoGzDen
Hh6rnhrEd7XgWVhfOGFOBBFFoxSwL8lKOHlg/TVAj6d2UARf7Ng3f3GCnxCvDQVI
UE4cdoXADRtaAPbPFIadVZ9B2dv9034YIWep3Ojtr90lUT1pEhQ667EUL/8IWS80
Lrd0g2L3YMLJjIhAHzRWLjek/PHsHHiQW1+cQwdXA5tFLxsCMvvqBUJuZ7iG9re1
BMEUFiOmKOo2KpW0KvaZKUJZ1jx2qPyL8qspq6DLH9HddhDV+97YpMPS+40gZ/43
pTZLsw4RR58Q8a01ikWBRxY588nqBAQmLZv3+sZWUQkPFvego8oGfnH0xNdihV7J
hCvaIG2nXcmUgByi5xrj0n+dWoyweYNj2GlC6OW09tBSAci9tAJeNe5sfyke5rh1
nltQOYpMXqPJFVIL3d8ffr25jqA9o/E1AYl8mESRsL1PvIOQFaBw3DG+k5AGKAf6
IxaAuhMNbTjEquXD4UUvr/9Y+/DZGGS9dL24sqBa1+cEBQvTNtgWFQbNmqJs71Rf
kYfm044aHDRTMt4qqi4BS0lr/VEOnG6omWr0l6qXJBLe+XrwS9wFf1wDVS537R1n
RzQX0EmhQQhnXSs2mgzVS9j+K+UsHyOlQiaPJfKr8PLe0chAkDg5yUimt44AxIOA
cByb6QoZ84aEsq9Q9jZCC6rzYnA+/A1cAytQM1Lhqhz6Z8ztIJ1tt37qfUQHVl/P
MyiOzQMEF4ihieUAGn9lExWDPI5FgOHS7KYt+Ae6OacS0VmjcEvqK5+iVrMohGfA
6TE8ud3dNq46GGGmx5ozU1svys/wKx1CJAIrorRst9uIpZKUbwQewkG7p2EDtQx+
eIRo4PuFORzUXb4KJhRFwvAnREZhTLO/XuPFsij58OzSZS1jAczjoGn61D1sRCcM
CkF8Wh774xqz+zufPX+aGqAKmKb+bRE+gDJhmtXnuOqVGkDgaO9qz/jZSRQbxNqY
4ZmQB9O63etcuDDXs/LASXLoL5d6xtacqHh64yr1CSRfO64gmbjFxV6u31IS2NCo
JhIYp+l0J3BYr9AyIQDkX1WET/N2AMdQnrChIXtzRu3nI+YdAx4NcNU6LVBRAYsW
sW4yABA64Ucn2HRChR1r7KSp214cghI9Tw9p7GgTMQteQ96m081T/fYauhk9VhDC
llLTXa+hZC08mkNEZ82AU/iuC642/Cez1MOVf2klLCvQ44k0b/nDas4IG+pkZfSX
bxKw6w5qRPTwLWySsOfTZpepi/Bpv6t9bmU/OP/g5jAPaNimZ6oBf9Q2gw4kLvhI
E6E76k08CpPzidEK13D26bDNaGNn03wZkZoMVg7vozXHB4TtE1iOpgu+NKHY1VTa
Pu62/YLSj6LQmoY7rfIrJLn4H8I7Je0jYnt9koKoYDtrqKdDWDjF0ZwIa7vAbmyD
xSRQxNMbX9u+CEAnK8LnwDiAYvqxLpHNVlXOfJJTib1fkIU+XJ58wmkT/v/tD4hw
mEWMzM5YWGKn9bJveR0GzM3Ef1smY3zaX+rodivoaR5Rbwm05aLCaYO+5M6nVbqt
HZooQ+ciz144IbVVGBQsTL5mFDlYKzir3utfIkmTOqtU8jDkCD8sanonwrjlNMzj
5C326a+d+4OhWPZ/FRgcLI0NChJm4HLkZ+MxknY1ofPBx+XyX6Nf+Vr5fesVl91b
TlKP35fPHq43+GMHPJIYJ41akvvGtIHyd40K2yuSfjg1s9W219aVL91OiJsOfkVk
tL9dyhwN4Q3wkNKAjnmBFr2udOl+1wDVuw2vCMamUIJAr3sHdm8TBWyCT8nYgZBt
/dB7Pg8ZSOP70OyR82JcvKznPD2Dou/EmQNK7GiKDFGefc52bvQw/f75WCjakWTs
8MwG+qPnATyQL7ee2/7AslTnezf0OyrXQ8gIkmA12iTmNp4/qmSE7M7D6HOKic3D
FJyCw1fOfzLxfuhYYUYEDzsYKN4u1fDibGdRisqXGjpEHmAbAR7IrUaqHYE4aGW6
4ant4n3j/jhrgA2TPCgoVuU6MfVrcNVYsaUYYMHe+wc9Yo+vw9uLYLqbC9EPL5PR
3YOW2Z/Mn4XTmYIdRzJR8WB17zAkoxPXANxobulFkogXiLspOY9GEHrosebuRhyb
PNJJb4UtZFyIvPqo5kZ1zmOmw8P79U/vAz35Eet4dqZMH6CarQS/H9299Z8xeNyQ
zbf0AALDa1eKsRzvBzvc2nqhsbL4osZ4DYfPDkoP7CcbUyjdiHJda4YfVvM65BFL
7oLusFo/76+otM7lkDYzxWmx173xyei0FQmMp5yQWxKggNPApt8ZhLPN4Kome99O
LQD+HUzosaLN2jCYdhUB03C9xphkLykjrXbWwt06lxtGvxeIrOPEMUQF0gcxbbkc
7/QSg/n9aq5DBirk4wi4pagFvKkfW6gr0+Kej9TRutgg1Mm4i0RJkWJ7PQoBEZpd
kQK7BPHMNWKreyuITVK11KW/swpaaHRHLSbjSadJH4xS+F1BGLdRW/Ga+VdWO2y2
hcEa4tN6zhHfOvAEi76yQwaWgxxQIM3t3A5MKnXHGgFprqQPOTDN3ick6JvOItDO
2PQSpVPeTHJlRyoPNnXd5XTiGvNFqCHkV2YjzekKsrhe9qexCZQXNYc2NmP2uyFJ
i2OIVA/WuY7U3H1VVQp/RyKg28SsA3uHEuUfm5qaJdMaZy4VeMW4Qs1AlSLJycyV
/t49aNviMClyv5+JqF3DSG1118iCSfjfObHYEC8wcojJQKlpCNfb0lcBljy6tQQr
g70WV5ZFnLNa+VnO7nbrot8yXy/RHiMvAlIoCXxO9PFD4Qqkfd7u08W1dcY5i2zG
8pAl4P4863QC1awzBbLzf8KePe4yUCybl0KeEs+Vf54gYehYtd7wRCBKu8F2Dxhp
CxmUNsnzbLuDWRq1Ya3IBg54R9RAkrx42nYnyHot4aLjmKTtpIoKIeRSz/JlNaUR
WjhaRuOAICMhk/ONDmIuG8fz8pmgdVEhnbINlsUjOeQVYO1ne45HYZqV0snIlMz4
1a5pWjpAgvibNWhnf3JdtRp8mnsOGOTweKJG+HEzhF4O/ixNkbjKmkTyvo7H8rbH
R0CA1tm9Wqv2R56uqgquboDdrGCpW+TkWGRfqfTly9KgD9RXnCV8ECDGsFM8oOVB
F6JK+1zl232YsmEA1zyHeEc5utlVMTduMFKO6SZZ7ff20FYI7Q9Ro/u/7reYoezv
H1ZlmZ7qg0H4s2RMXjKKgoNELE81XZOtSiyyadhge/uCrWEhvn/kV1XFHWR8ytpk
qer6HlAFoqIVpdL+9OIvCbuOjuebkOmEOgX87y8CyKEdPfQ8lLGLlXV2iSC6igRF
+dIbywpgHoVmbbiIn+uz6UsVC2aZtwN4zYuhhakr2TFgenWZjaWx50YsesfCSGuB
viipUL7ylh5EelfqCI0ZRYYsmG8YvIS65hQJ8tLifw34ULTWV93WOEVYmF0Qrfb3
0GO9uQ0vOA3g0rM1JhALaqY8tKMFZxUL14IRR3Ebw4sX2xnq68xpFcPFaim5kArb
v/N7T4LEXb88daTYQZbIOdqWtkC5Pjs3bnxsWRmtkm8CgcUQDAm2J5qsAVTHdDdl
xj2ROYMKDySnPT01Y3zghv/MIQFp/k1D3DuEnrSeciVHAi2fAUnzjp6orq5BQ8h8
7AQP59qCwiVpLTagIQKf5ntFO0vOehKMVpuATEz4pnCBgqxLj1ZxHnnisKie6Gp3
eZx0vRdDe5vAyrBLHJ7jTuLIVURbJNE2iaUj00Xksy1x9rMxnysLirie3TZFCZX8
cg6S8BSrWpd/b3UGsAkFnmrQJa+/93lYtT9VIFFP1A54R5y6MyFD7Ak7TFiKM1lw
ICsbJHI5o4FtyUKlJ2USmWUdwI1VKpYJythkgVRz+NHR+0fRgBzAJCEEZnycN2yY
vM4ivBjQtuaXVgqWhuMkmsbBTv/jpYxFC8abw6FIRYD9eCmqqSP0wP76Jx1FMH1H
II9HiujsZfCHrSmqtwZOgXMWLwkR809m9wA6JWMNkRuFQEEHRhM3l0aTYe73zKgS
CH3Pn0R/BwEiuN07cC47EQvOq9sS33eLM6YLZ5FjDV/L9+Dy81389iuG7/QDisTw
wapR0x8hF3QTRfPVmz0LeIMMTFH4/2uHqigezqIchTShnl5TnmhDMxTP/upK759/
iPyASoKs0LsRAQnRd/bCjanTYdOs1Dws5tNl0/3xvK5JJsD7ojvnQPQ1UNlC6vB3
KstAbKp2VbGjAkqbSz0oljoyT8a5Sfh9Iv8ENGkclaHH6ol4lnZR3EQT6OyXEcKO
Mzg/zpMV07AXgAly9cQH8GDtU9ABj/l9qoWw4o9UL4jAcwjj3QLRRrMDPsNGQKXJ
N4WJCcHrsSSpaghovDYCzpM5ytgbaoHP+UQaeW8nNjCuncFBQXJPYYalHaUH1P/B
Si+0k4OTiZZIn07HJr1hdN/wRbXce7ZeCBMfTNDq2R++Tpkrsl5H/AgBzk2I/l5V
WB2dkPzn8BRBbE8FI7KwKY+hez7YFqxFQYU3sOtw70bnixS3In71OswDlJPsXcyS
bluVoPpVdpqMMqhke3ovbWQYUNJYAXv/r1GiWgnERc2vosJm2hztvYoHwBGn7ju5
Z+5xMKKrk8ypJZGKX5hjRTYcwN7zRM6J878S6xX4pLR12AG+unZWo1/jObqKXoUu
63m/5jbHfGYHxBVGWPDh93Ftsb2n0ic2CDXlQREvqgd61I5/dzWfUP3jfkBhTN7Q
oXGS02rG1KjLaVAJDfyViiQSB57nCYGmCMFJRt2y8k8/XtXzkynLt1tL181ZA54b
QZSsceLVhu+LN1QjlUfMBd+tNcXUe0asZ0IT2TYdLlQNG85RGM4927OFHVjppEFf
5DTMuXG3Hb0e2UPFYUDs7wfM1OHY8pbmv5k6bGOnZCy/U/+snLMhcAKhoa8BbiAM
qyDvX1Z2eKJJiuNk+FYjdDSzM1JajpHt64fWfcAxJXsawsHaPmP3w9/n07zU6dyu
SBPhRZ2y0OeEC1s0aLz6yU/co0d0h1/NPWG40nDa36CMWAXgQ8D8VVU9EkRW5nE+
Y5cxFWvaVywUw92a99CRvIpKlNt85pj88AwBMH6bZC/LrNQMhZLYiH+caSt0nzia
1V6jykgYaK4AyZffREw/N5x7BiJXT6H6+mUhvvhDKWytGiHVt1QJnZtlsUjQ7jb/
KaSjWg3pnx1eag2cNEIguFsq7pMW3cfoTqRqBT/WMh8bo+82JWQ5OCcoIZIZAFhF
d3TnBktEw0vN4TwXmy+VZ7v8jW8yjDRm8ASaNDcCJ8Y+sfDoxgNB/gHhft/BLLKt
LyfCdIb73YPvrjPdFknH7LWzZUDjDYimoBqbwHqtX+3NqbaLfehb3pBi/RgoPyCR
N67FKn1fSROYSCHClxLzNT+/Vsdle8eUrP7+o6lmEKE9rjo/+8IpVtXOMAv7lZPB
G1d3RCE84BPlRe/P1k2P286MEl4GuvGG1VH+Yc52otJij9Dh1VVOwDOTUrAH9jZ4
7wF9qHMcXyGhySW8hlP5igjqCU9UBYUQt/N4sx+ZWV09yK3iW39wFJORg98KCBXb
953c/oAQa4HFWjCsbUGWAoNZmwgNVBGGf/1sk1OpJR6/gaFQVfCLKYPz7YqHe8sD
tewxEaU69czLdzi86gYowAMAOq+VMFbynNHVfDx7kFEGgt9u2OLOZ+txv72LnJek
X+s5BNA7fevi8/BHMmuAmV5SPqRNM/fqiSU+p/+8G+aKmdE2KA+RexdttxNzvhSf
hDdaop+YaOrvpw3w7qBXIu9ClLvKfwDIHVyHGdzm06EtBakf4dP5H5NNf1svEXKD
hUxzzHw1LBWK8R2MpGHnxReLS6vXhBgvAED0u7dt+DSqR5b9qmbEyuw77SLwgQaL
IjVByLB9iYJLrLNMPE55yzsWj6RFnY9sPuY1iRDmGqra0pgH2iWwuWWx/4i9fMB+
eDSWc3H6rU1AIM3RwaoKYHiE26gfjQsPii6ablezWokvU1AvNCuIh/Lq/2iAwfNc
3hBJl7Rpah1l1eqafLVpEhWlJ50nOYQxnPcp0BTxoEDge5jsLgfjHy61tsH2LQfk
sezimpTLJjMTf34LWi82UX1mflfG4WhDEgZm+beuWWIXzI7I7EGZfI9C3+s8kbtK
rXC27nNYfafCngECbgmHrOXAHBeC1XArdkImaM3co+UVpkDwt/DmvuiTvl44eaik
XvUraOyvDKd3inebUwYw4HNu/RzMWVfrxQh41Je522DZXVBRS+U14UtGoSe2ut4d
3NBLPMnmUfQYpHyQOD9DrJjhIDuE7LNFQG2359V96PMZsIs+uKFI9ZSQjIMkSlAH
7hIxdXJT/AjNcY3lnQSFLk247LWcaoV86qpEqFnb9yK/iXzCwbYfYn66TNP+9mt9
JAKsO9B0F8Ymbd577UCoz/ROTH2jbFzVLUZ7AKzdlENgEa8pGihMKzmYmqCkZo2A
sIhYTxHdgIJF/FVf4iHPcKs0hUB5TAW3cR+CK2MVUD9EzZ56vGoyC6kAEferMgCt
n0H75A8oIuAEWGCkYw5pzc8p9qnIgxRkAz3CApiSS3NZbJHCu+N7+HKWaimzHKuK
B7/I57E94ukgXdBX/y/r1de3k1ga3tfVkzJsxxySGTc9ia+VPzV2HcNYsd0UTc9a
YasWOV+jf1wjPCtluPqaOra/dpgO1NOxbPhyoiT5c6uo6bzMCPztFdMWvVH/yGbp
Ho4OhbAM6aQ/1JDXtWnNCeefkj2yqsnWSq/8qiCEqenkcHFrbGQfHXiVtRKigwh2
GtVzNynagRyMc4QUmgjEmDeN26bZlqAEuioghkZcroqueK7gMvgKK0e9rejIZ8DQ
qarVbIbpGKwsIZi1mIoIIYQjFsQmU0UlkH2NU/NSH0eN81P6nYMm1XxZV61qnnh1
pohueKNYkj/GhBcaxk6AXvKQ9OjBdeS1mrWo/97ruyar7BXFOYcnbjk67fJPjdsy
qTB+J4K7jXuwOp0QjN2uuIRb3DzoAAPQTMCpfjWpTq1jzR2UCRrrWYKL4cEcVE1w
QyypsxROtUlJ1O8xv6qXaALZYwT11fyJCNIqwbOYAE5uM4QSs+OPf3C11eN96CBT
oxIU1lWdCp7zQfotI68aSEitQprzei4YyARHvh4ZQaIqzI6KJhyvSTwNQp6lAoS0
mRe2PkTJYjl/YLuzb+beX092WRA8WtZdce5kmNDFh0bb/JDyjM35oniF24U3rJRF
aLSUw3nr1Cplupj+ZZT+L39UAyq3QGG9kJgjnZnHwQyebEuAKjqEOmtVCmZ72r0z
KFdDmrj0GVgTLtlXVPYrz4TEDda/ENA/EPy3E0tlSLKulSTHIhB2I0i5uDgo07pt
HMmV64M4OfsbJs6j3W8WpndtdiakyCgfoKW//umaUF3RAel4yxbx28aw2q+3SgOd
WbeSB7V5GZzZpM8Q56HxPxTGBu/1U8VJz6EZ6S8I6NYkUhrjx++sxTUEYDoksz0m
42/D1rGN7zVznZGKGtneG6s24xBUpB+oF3arAxBqxUC9U4zAN6WrTCHO8rIt9xod
bG4pimpk/ullTFpR/UPj8LLaJDYb0VafSzO1+r4kCJE9XtPJez8zb3DkkOZe986y
dsms9pcKjXjHRtdTa6BWQIZQbIUgkGuJQYspDjNol6vk/MWKwefaaQwGRf94WH1d
32KMQKWN61TmtbHclYjiLJPyMIG17Jf15fDya/K8iFkEEcx2toAIqKuMlG0PeK5m
R0C90G1sTP/kfVkHcrfhCcLtyB4kwn9xJo+sNIi65nZksJ39Rb8oC88V3lg313YU
EnizQy2Q15CloD+He14U10y9qI5AfuPgZg9cDHKm/IZt/4pyGJWGOWGbGtuZouJl
v/R6luPb2VXjN5K0ts+f/FoOcxrKw7oyei15MCUZiqVE+HDXbxcUEpVYLeHRl+sM
IK2300lVt0ZDA23RVmpQMgcACjyk2OV+0rbBtlRxQ4lu1UZIljCG16ei0ORiIRdu
0uvojOKsx1J5ZI5rfObSpVdKXhh/Lb0zXtoFEikZff5onB/5FZxvTwbvPRlUCOsr
s8K/BK4+QlEBu+O1VAXcS6SCIE+8xrEIWYjVSXsVgBN75/oDTiicUA8L4JsSIhaB
nN//5zIHq9bD0eNwKKrlT2vc68249gnKF09m/0i5vuwe0QSizu+rZQ+/Q0itay3Z
Tty0SAxPMI5JHHlMo1mzwfpZVqA9qUaCbWotsMrxvr/ZIJuByPpTMQKtJuTKZDdc
KlXPlW3ZFGlclpTlOSf2I8FWiAHxOEKA/5vR+DoQy3IEHmkB07HsGaTmiusT3KFz
99Gc6RLvblR4qaFmGjHCiTyv5sdk6mC7WL4Xo/k3D/FEdOpq0v7rI5L1/s9ojT2e
omjQ1fwLPjwGrQIand0Q5faYHVxspenoiJ/gCWqGDS3mgpHXvy/PZy+rsMZckofp
Jy4Jtwihkksnt/H5eAaEFZ21uB7MtsYFud3cXHnqOrBa1SzVNVePfkqOO6uXNEKa
cJfCDMbuCu2hYbMMVe7AJtwyXLesoTLKJf2/rmjmf0Cmkd2wGBBHO06a3H5dO+8+
msFuPNxqX7AwWlT2baYTO+z41ACgB44ezJ2T4c/PAJaROlxoYvGMoGuUMUae28WS
kdfEhP5OW7cOe3H1e+v1c2gONCA0nJtuMv+y1tT37WRKDGlQx/uHRkxzkWznwfIK
LaIpyjYHFNmCP3X4ICTHKHCX3EDXnMsLhhdkEqK8dAmHJPGuRMJgGCjDsKfSfdaL
vGiUtSvwPE2QzPHYrirjA4NY0GP/rKn7W7kFCwmtEJT6ypGUMt4BgdmxIsYiTmI2
613CxQybj2L+KS+GaIvoJK8MAVPpxTRRBfgKzOlgYL3bC0ZWM8zW+UbYtopu/I6B
sB+DU88ymH5pvd/pjn/JooOC/ct1lThAlfeuftMPbmswhZSUqH8/Iv9J9/DFefXA
rK0Ie6DooFSNUecf0mzE87GB7cNAbQ3jhZGenxyYVVtHmRYoq3Pk5fuYRRVcyxBF
/wPv3RB2kbzsmZvBgx5Qp0BjdV8feNKjQT7IyDkJKYFfHsLI6xUPXtudEU4WT+8X
YZuSAmEL0gKYaMFy/mLvCF1gNTxzmvhB/0z5Ot9ONwfMR75X76kBNITZulp7LFUF
CqluqO0P8sNGiRuOHVc6gcA5ozJ2FL6st9i1rDjrDGMHUERQPTsHCXmGnz8LHH+W
Fa46mshogJC8YdUq+6CZA4x+IXO8ZeHgXy+epOKtEr/kneZ79K6l6qP1VtcD1j7V
GAkSwwQQgo8XVslm2U8IVdjMYZM3OAYQL1UjqP86BP7qiiJZT9plrBU3GN9D7UpQ
JOLkMDA97fiQKC77kIxNNF4/id1ShCMihoIcXwUfiUk6nhu6ybtGstpvuwYUbEYw
iW3tZWejplDSEhrzGrCcnUdddAJywI/gb2++3RvNi+1jgxdtLT/Fp243bAx4B4fn
IEa79P6WZhHe7wnRD6DCfqn25ohy4YuCP2Bx3xItn2Qrs3HxgFu/ui+nC6Z4uo+H
tx9WR2j8bZa35namk8OzBFZ2fxElexx1Oc4ZF4Qi4s1PHCezjJGn6CaIjXvCWvkO
Qu9Ir2fzQDBvwHIVU67FR05GitKfDH/pO53qmPEanwjog3VYN9ik2yUNDIi3kpKv
UDDutADjm7GpzXiOWPtRSKJvlhDnCHEjYkuF/5FxvjLhvHYSrDrdWWQPG80GSEgA
/hJbItLlD1p5uO1oaak5dPbdtbWWOJVtQtxBuB01fdBIDiTDOaSC5EJiqGfeoAQS
dSAB4u4BYPNY7xh44JrN+0y82qO9MSZSj6t3h8sDngjGLuEDAzlS4Ra63Hw24S4E
KP6f/F5ygchCOsR0Wi1I2XcZndS4bICuA9eGvJyVSTN94tQm83QaZHnUUElBEZWV
ZGeSai0FCB8sTxVYZM8Prv3jEismiHJ9dst0VL2jzE4x5dhGru8gXw3LY5oIY7P5
LL/+dHZ8F5KdNWXyBOkqb215vgZQ/L3eY+u0JI51MlW+BzVWfYY0V4SC60DxlT+f
LW7Z7b932fZM2nGtjwL+yemrv1seyD4jhDookJGG1nDwWzO/qskteJFQMDWA8ZF7
tL6seWaDkkC8zOCLPbsaGNzQLQto6foz/EuefiXjsdApAA1g86swbW1IPXu83KWr
PRsCFQwkoJ/S5NO7NK2Hmrc1dKszEQJXaLbyxZ3dR2zGvIeNiIMGm3FS0nF8opAf
MuNrNgIkAH3/MccaciYE/0/t59IcGzgPtnBOI/ppIxGNpL9D0r0//Do0i/87oD6/
jvr0ArXlyhJTUaNRU5U45GJHqG1lV/MtsvpSJecJWAWG2xTvitcs01j6xPCxOixa
nOGuolIvq8PSOprjufKiFUgXxJLZogj6JGlkAUQAtms7ZakW8Eb7rooypSDft1qa
iH4KbVIwPhp5k2/mH0YTrro4LU1CDdv/BJAsEwPnA2iVMdwSKd2MRsexA02yb3WP
JL+zX+On5536WrflHxK7Nhs6HR8MMJFWuvqSKxokm9DvfDpYotMHT1wDxl2y+prQ
eB1YHn6NVR9g4JeOlKGE9OAEaFLLzEtBIvX/zEqrHdyXs4cTxAZ+bN7g4GLDZn4t
bo+Jrm8ZbxYdB5i6LwWKiv0QdluxtSL6eA6VSSlDUth6yMNBnYOihef1/QjY22ZW
r/R1DH7N1sDdWcNiiGS4ppOd06/Zg2xOafcP4Y+eCk1uVn7csiD+165p1D51d5gc
OPU0Foyh3NjVvkoSmxrIbUcimverbwOoOUQ58XEMMXolCy2xsgiL+JLef09Bn8r/
iSezk7VFDnwUALoh0qzOK5AM+V1Jv+L+txuWoUhAlI44YkuPOo1RC13cLXy0HAj3
B6/RkL0PLytkhvaQexIGH1euSnx+G62GRwDxyQKASQ9ZW0F4zm5cRKy83XuuJQu1
VX+5qtk8dnYMTm08ritHe/QGWxOLOtLTqsl0m5u8pdnlblGpHV0KBvSFWIkBmgPO
Jf7V2pD5XZQXN+9TMza6RbclEuMMSoqfLNTlkizJuscThwpjHXr7JINZ7hki6nyp
h0jqRSC7VLYeJoNQ24FKoxvw5WNAStdnAG6zVHAZ5eDKmygWwMnonwUGMvG65GYu
ug9UR4Ljgrfxcu7M6KhhtKA2RFbxhpw5Y03ZFwnSfEdiSicW4tpj7gzOR7d39YQs
+o53Ts3ev/5sG1qJ0isvn8VXXZT1VXAh6z9HGXOdzu9eWnxKPSz1g47hDiM0SoWb
F9EDApk1E6cQaCuPvnI76Hd0HmcguKs6h9qyrURk9Qzmm7fyvWBxJgOZsFTRDo+p
tQufw5KDm2ImcHJ3Q00Ej1bfTZNgyX+Wc+d9CEuvI8ZZflxNw0+aPjwv5r0WW6xf
2+VppK5U/yI9o9mG69WVUMEaTnfK59G6V4g39O5AifhbCRfo6/WZpkVzJst1rGJd
GWtido7a9hJ7meqC5roX7/jVV3iTNsuGlrm+nkZRnvPO22Lusv64DgbI749YToiF
B/LfwEPbPuRRVFk5car9SfPId8rjVabSYknV9tkiz0bYdrOfG6eLmi18CRu7pfRW
wPhHFYa5FNpSL+XwnmpQ88vgFtONn0QSckNaDwJA50FWy4FtYcIyKdbdTGu7/53w
BaU7FETsDLpNW3+b+fJ1p81ZpkQCjjtbvpqaR3hyYHGkyBd8UZGG1fVPm9rZ2PLC
n1RlPMyeDD0FGuD/Ja1ysG8zlS3+5B2PHgO0Jm9FsA0JtCflqk57Zc2Zyf+RhDs1
0OEt4m1Hb9ex31INMiMzahlWiSgG7KPrHvL6XvBWD/D6Vin/4Ux3uQ7acNT1FA9R
5fbUGOs21rnpXAxs7p31breUKh8yLCy+3VRKyfnxWpog2VlqCvVwf2UCQuk+4uV9
oqHj5b5TNOlnQCTk57zduu0QPZk9okvNzfpVogkfbhpYxq6RdcT8/dAONeK1+T0G
H8mOSCVses+oDjWqkG98krQuYPcVAIwOabLrfR/6KHVrdxkVy5aCxpF0+r3fu8Ll
j25XKN31jsU4Q/PgF5KhXJXXerFVhVGcjT7kkYpqn5UenNDZjAT2ihunov7Faqmm
6f8ngQfxoxBJrtbDn8M1tFCuHa2NdsJZbiZMSm8Cq6GXPmhrPbuGmG1dU7iTDuxm
GUK8E0wEVBeOoPNpLGuLzIxlX8R6TSmIXGnNvkbQVb1wtZUAdsvxCXODE2aST8v9
b6+1cOfBDBnqBvJLBAMIZkEbtBzP6/3yKzko/jDUVcrinFTyYbf4+44lngcWIY7h
rM2KKex6u4DDSxnu7Y/pEv+UNIkXG9RIEjcZa7n5wh/T6xmsWPDJWjUWA+HNe+Vm
Wt+FcmI1fU4dVPgDoPyPHLqeH4/qt6uT4M5h8yv+n/66KSfJLZc9XmsL1O1q0+aC
QdBcch9O2w0wwkRBtAdjw3dn7SYsyAiHvUvF7jwctEod8oTE3kRx6+ruh7qU3W3p
Jv8miWtPGH+ZsJpVAzYUuXrPKaJoUG8bY1MJez6pRFaqBLLfobcWyXxGg7uKhVtU
QV6PVlUV0kNjFvnFxu1P7/PMtuurOjzsX8dRk6udwbHksTVXkYJU0m2YfumFfyiH
H/oPSpLKFErzpIYTq2br5s/KHOUBWcC3FKsTAxlzoEkNAUR6kYieTQlDHciY8hFy
qOMRqEQG3BCbO620vpmH4YmzWxWugC93EJkUJrNJ+IVi7vjW+oxpADuhUnjF+sWz
JYtmESm09fO8mTrHwRHkfI/C70gZnGsG3o5Wp0tu8lTKUuE86phLiqUUnucOSeVe
/5bctzuj3Ok+7j3E6Nfc705OLYJK2dbs7yvDRwniWBpYX3TigLLyA16if4LSfPu2
QS6HWfJcl9Cb7YzaKRUNyLOFhfjLTKuoSbTEJYjwVDc+lzdu9QYC8zGZPUkJFXQe
oXW3VgceRwBwGEq5MUTW0gFyBky9VOhgGgox1duNcj8p+w6sjTwFr2SP1xVyua6p
1iXozX9u1bKGHDikk0RgYDQOZzhLYoZeFf2zrq/69DV91zMKx4nvm+fKHSwPqVb6
svLgM9WNZY62sjttp/LfhyC/gl8hcCgN5qqZYLuUlwdY6d+lllbFcXxvax2L6wQ3
po8+9FAc2F25TeOC6Zb/y3xYE+Lmi00YVBjFFBpI8MwuGIpfE5QGe+KoP6IcI3WH
TV9knkygpyzZw8XuHEjv6kjkKqfeif74nYI5ogyQUU75+TLW5QEjWTacRJUOsVfo
2p9Th7mQjiPhaFOg+tG+mVtpGU4TGA/r4Jjgxg3nwG4EMjgDgWA4hAyuGTnuV5ex
jTARNTwTl+Nsak88T0p3Qc6URjyO8mGOrdyy0qeqI50BqL8Pcbp5U64kK2lWKfC7
BTQH5wV9Yx1ZiUAmjLim+MWtAhjcBc18HS2p6v/1KHNDXVFdCy6fKWPOwUJVBIFT
fXtTOMad0XylXW4wZmdoFrETm8bCnphzjUt9NGpBCzuXS3JId34ZSogeTyJMLFiO
AuXjVR2UyZOMYZLkeU8+GZyWMsmWazzq+tLB8hC7Y1nPTDBAOQrVITFGQtWqZ8FS
/asgqHGkvb5QKxlbetJ/OJ9BxOId18FTw23GX82xHEX+zaOIBn0OCYxJ++nQJXlx
VBIKZNRtOAGrBQ9IAxhSTM0VaaWH+2JzqeZGNoYKbvrxA6hECvB1jVtqqCejnIUS
atwYTqRLBbzJXg0cgjaqBGpt1+zWHlpKfMTPN6+PCd5IWT/6a46Hav4RsAYa9OOB
2JYq49XhgbgoZ6dB3IpFKLsjK2y6XOPo99Wug07V1TD7UmyMHAwxdvZGh0v5BPhH
6iyGpucmMwjR25rxde9RlAaK4ZxHqJYf+aZaa/6+5qpiSbDxIZeBPIX1OgIkdxbO
f7SfrZOTfwQXxWAT/9WAtNtGA4FO4L99sLl2YcYQFLl8ilBLS/JP9y4JLHzgWtQk
FijHosDIdW+E+9pK54EumRSp6ViyNBJ0Q71OQNU37K7QuTsDCGAWb0FHOSTmqsWZ
3kQ+P3lSeCHwOoFBsvs+KNN1BInWPkvsHrRCNTR0jR3DO4eeI0Xz54u3HbR1VoaM
VpJRxS8RUGC2EuAQEwo4BclBoftQgolyIK0Ty4EZaFPnXjI8SeFVeTmpHg+hUJ+j
SOPuuY82u6fh4TcyV4aKzTPmxufxttY4m9nxEtmF3S7SprddWXr/tD7y1WtF8Xyp
Tap/leL3hLR8/dndosky0I6lLNpBVzP7hR/ovjJ/NoPug7ac7RLR3nk/bTHR1Caz
8AdMkXCImbq/8ZV5J9l51/Y6Yfo1WK6ON+wlSpIqZ+wKBqlCCoToA1NjjbFWZT94
LcJcgyEvsT7Lxoy5ui0ssGx8hi6891GmcTHjgfYL7HYReFfpY9kWNsujeAyX65Xw
eCcEDpMNTgdPf5uadNDp0JTxbX00MANWytvcUUZF3iTEm2xO1sz0iviFHkz/UENT
kNe124b6+y7hbZxcz/WaO19a/fn0unE0UGukm538dYTj8CKlO8EORa6IokTCFt1z
Qci8oN2XOpoi/P5aBzv6xY7B+XDWfX/rxVeUM8n+l6sB9af5ZQBj+RKix8AMbOmh
8sX0RXFXPN4WgF2xcy+JcCer3V6TIrYU4EfE/8m5BINWisbwYAXHrtIfLitfUZx8
2qnueGiZnGsbEgrHVyHCQCn0zFgtX47s3uQxnjo3naoAZk/nwl+hq8rQCScbGZU8
G9LT9DIKaApkCCdB6p6+YADnUhlh4pstK65K4Vz0ltAbWU6YQiwf9PMGlDba3WMs
jYF8Ou0dh48YJvLuJugG4+toNRP4I+ZuxXGltGzFmgEsT/w4p/WvdIbzk+SVb9jN
RnLrMqsUjw1YDAgn4nC7KimFRQX9qLO/gNv1ScjjjUrucAXtw2SGDGLcI9utSWgs
9dgLTVk5vf3mj/PXFd9wOquCn75FaUBt1VmzatFbxlA4gSCfbH9blMVg1Gtj963O
11oOOgFalMZK9xX01ttupQ1IE21kZSNet4xGl7v99w8oy0dMtuLVlzY7+jDveyis
Tq/ij1FMbdz23a+3GBkEkmIkBCMuhC0N1MOLvth9S8nYqP9KFoCwP1/akP6R2AAh
qssNguTl5GfQgsMUZ4G02wmZzLNm4exVOe/8GIVxqmbdvwC4aqQ17ah6NI1gB1E0
OXdujjaopBzpwIjDxU/kUWxZ1iOZPxYjTNbPQV2C3eJnhlcI9am1hFSa+NUSZl8g
kiS3fhJpDEG78iWuPxwRHFjyc8G7EIpl04jWaPhTn0K7Olel/7qB40x8rfc5sWU/
CTnjqfq3WgxZG+JJ0AW8WImE799OLybyGKJGlUI/TWmTjMZEQjrJngX7AyD7hOYa
WOl5wbW7pLrxFb7nVc2a2oXCZxBCVvTXlxx8qU1ZPlF2IWR7L9ti9MMWRltHn5zw
e8/RFzSblerp75FOqjLWNnBk4EYx8EcjK7jiQddHF+bRqnVJB3ExG3Z9QMJAIGdv
Tagh7P2hcvx/tT2T9RdbSa+gBE8cP4KVLGzYk8Lsl2xmhIb2VvpEFNFvjIeWMQFU
MiJrojh0D8VKGlm1IkLhNZcn+8f5lY/dHBp06vQwR82WmpsTsxMZk9aBYiJSdAWk
+aMQ/k/XJUp7Eg/ej+QQ+qSbWdJ6Ja9i5mULIorzTDWw3y5aLNRNgoaKxwMpMSDj
e175zwUaPMFyl8xjRFdCgDI6IMNkh5JV58eT5bNi1A6nRDLW3qgKN0kCRjHz+Q0v
m0OcYzk9kMAzmvr6VZKcoz+xmR8xlfsNh2USx8CxTpsjKwVE8/t2AWF3TBmSC5kQ
NZzjc0KEWhN2gyyCuSwsP0Lem+436Tf1qxAaLRZcRIuWyFOSau3UmFSEnd2hEjJA
pWQfsxdKLchFuXgMveRbbsPYWMJ5gPKs8RGGg9ioYHl6j94iIqZlwGB6sZOtuD+O
Hz4bPCTRk4Wy2MOSzF2MJRSqamXq79ySXaU+NfvPpT2nCWOYOQAFDMD4BUtouPEE
GizSVzY/QauYSfuJPYGWnlMqz66FPQHkgz27GLfpFmIFdGpQ8rriv3EijbDWnsxm
AWFvZNRJFOPAhUTzUEz/TP+ZWJYkNMM1R3Dqswyae6QH5l+xfl6gnje7q5XhH80a
B9zx0D3MWlwYGL90hlHetpls42ik3HFHozJJ0z3SVw4aVTrg3eoZkfPkrfxlHLhW
AoYf+PrWibXyBcwKZikPuvgxtp1RqpvhY8wHady/aXbPyZNNY25ZDvqPb9K/gEro
MmATP1D8ozjkDDYcBlJ5jvhJTQzVg0QHXVbLHo8+sbYlnodSCL17y24J8YNiWCXW
RaUy9zx3qWY41f0ga2jlW3AkkAg2L4+8XcdHaBJlzRMH5ufmyeo2tL6IhT5lkqF8
4rfAHmWMSr8xxP0/0yk/nUM9n0FQgJI4/VO8Me9odop56x6YqPQBB3srQUbkX4MR
rsAxwCnPYUZm3LtfO5ojZmee7LidaW7qaLbQWhiBBmvlD8RHqQEUflkCbFwu/asw
/i3Bgi4eP62xzyXGuCStnjakIBRnFpQ4NNPIK4lr5doYDskq/M2TcGlhlr2VUM5x
r/8613PI5O5MYyepNbluXVYs+CyTMXfPALlcFkWEaAU1YaFOgSMUXZXe6ClBJXHX
+rTZLKZUjpQ7RSSEH4NHNCTn3PCGVgj0tYRYUwmelagxsd1Hl2t9j0SaElCceyLV
T7mXmVZ1KQE9I9/n0wZA2p7zs8iThJFmUhJCymm8aqhpckL/AgmTi9/CYkXwxNMn
Lt9XiwmM4R/V89yNZIfLqqxDHiAq+UVrU+qQy6b9CiaxM2F0ReMYU3/C3CZrVogK
lDyDDYf+Wv8oPfftUIuXEJgTPOIeRxpaZvg1Wvbo/1f5gdmIbRun4FKmrkHpEqKH
rLsUVPmJldrtXRlsThZDrAD+eOXBajSkZ9rBTzeBzTQB5yOke2ud+4IWO9ZS7Cg5
NnykgZYmU2hOGBDkzvk2/OxUEXgyetssTpRuHSkzi9Cnn64VFrJC+hx7O4KxkVTH
YyONa25ZdkuElQr61RQwxyR+//+1VLHWgPI3WrMaoWSxxjH69ptx+7lzoRdOSbw9
hooXVz/beBzkzDm1lHZyZeNUDyH03dwYh5SNloPNyHCJh4k1euf4KshcmrA1zBOY
g09nmDcYpITgf5q67m/C1JFwuSdCSQaAD3yWo8f0g0NjkLkEvmOSTwES5TQV2JSA
I3BHeH++7tq6p6+zf9FsH19ogcdaRyQhojiOoXrDD7PO565imc/ezE4aeWIBOv99
XpWaMgcWrMYFemGYDhTbiPP7RwRDZJDd9VPXM07UYRJhIF3ty8N7PZ4s5d2g0pPQ
AJDbleqcj1ghLoyaupFkmyn1N5vDMilpy2kl/+gQIsYRUG/MWPbj//QuA12enP94
SdTsFWJ9BmUEoELoP4WZCvplr7QTyxCIKp4RW/pWh6eApKRieKX8uakoRgU5mL7l
ojjMtCkLtazYG4EYJy4mSgow3tq6J7V//MetGp/5jt/9GHmfikCI2aJ73zYZPf8Q
MMq9L+NI10TpMlOSm45xHCr6yOtENaX82glfB3l1iI0pNGhxBn8hvSr1bA48HaTP
sACCaTXhzn/k1v9yeiaItIUfuAoqo50pj/W6imhaAwatNCl58JViUIu67ktaD7N6
2aiLsGbPlFvrE5g+6D6U2K/IfXDFsrSSgUa60kjbaPqaNI0vKsYNW0lSi9XEiqh8
Zu99UaZX/ReHmg0iG4PPANdv6shg8FxgA6rn1fHM7NvHRBcIf3UO9esi1K3tgxBM
l6pGcc2slcqCf+PeND5mhpgFtW008Va/Sr3YXvR2T40I3Rzjt3Kg1v7vb62RVF5N
as+zGtt2NxZALiBMEXTUDwOmY9sJDTbtWmyRgw/NVzBHI1fCWoUCAyVdlzQY+i7d
BJplG8kPIfvKbwxv/QgC45XIY9pHA9hjU+fP03iGsfw++cv79s6I4aRe6hPfNO4L
HaIU8Of/iLtTFcQCCWqfFXF4Mu2k5DA9uhMPWOB9jIToiU4yUXhRs8T5gB64g6J5
SfieaoC7sZ0m30Qrn1pGklD4w9wItJ3D1+I0dcC5REckfVLl0F+5OH1Qowc/iuz9
6pb6NVn3PBLSkrXkBe5kW45mfUHzhNvpr0+CPcwx56vnG1vOCGrrDLAvyIIfIoEI
V/u+xBtzlDp8Nh0N7HzjsOyNh2sWR0fBV+ORF4cW0HRQDpNoUPuYNmto7U6bsbEj
/mVMk/4WnnruuZc9WjiLsWGbutEnSeA/zQ6eEPSaTepVqhvNuOEcMqBvSEkoIowj
7LxlJrszV5CgDMnjaTOrTiwOkn538DJcDrlnBLPOA8kTtNuNkOSqaa8Wt5/+wlXr
kAjN5L0NHRPjCoQnW2yU6sSKhyafCYHdDmdUf7GuOGSfkwD0e3LV/9ldD6LMSVkt
PcMn0CYvev+1Tc9p0Ma+lJZElhQf3L48MMmMOl1aXn/UyH9SodQW5wbnF6v3Lcyd
cWo2a7vsMcoMrfqKbRJC/+5bO700pD/bApcPs9T9yUIPP1nND49xhgM5AMk0xCzA
ypuq4nxE3SZP1xRfr2X7R/4Lo+tBrFvsJkg4iDgwMMmf4BN9oIVIMnRJfXfLzx46
bd1CEI88V1qA2Ke+ePo5ptXkfUUgSkpvFBAeXaThf3AF2BdQPQOTkLEFl+EKIg4g
e7LB8HAQ+xinbBBc/BwBQNQTCcdpkIqIEuj31x/yePvwmZhfPEf9wn+57dlFMXeA
uuo4u7v0ZokYJE8YpmzocvKDiecSYqEiD0B5T5pSDCWFGbWZ7rCyHK261FE2CufU
5fy1FhifzcGC0ZHAT+g1cQrTe6RwJNy/H0fCLzo5RDlCifRVo34bRPEwfYdYqKsm
sRjpFjVM1OHbgtoG3VMtv9SXONrDMPdYmZTeym4/ytO4pUwlyuE+hXP24kUAZgwI
gBGwGVZdhlfFy/mlkZbiNSnEpjxuGhpBIrPqHjLAwuFKdDt+8gMJ8+LZzS1/RjD2
KNkoedrTxpwoMixW2V3oFNT9XOo3bF9OxUE4J1ZVDn2kv+fx4H3+ds1Hi34zvQ28
ZbQRuICL+AkEjTxYjPnwVT3bJCeHEO/SXayVRnpqTPsBkr61gwJcTWYmF1exMNNM
a/w8HzOQu/4jcM9i0goAjsOTMHgZdvXU/PeT/x3T/kVfs/PuqPOR83Oa7cFJucP5
Pj31f9NWd939elf9pz34ta72E/tzXc1EOBz8FNrjvWzkrmpfhH/Zpr6IX1MQQ2JZ
cNV4zluERm1RZTQ3SsFCQbmF0oYn5zQKCSq2n6UItzKx9ZS9HHAhLiG2WXJLwywm
yRDG9JbOyZdgt9fKcbQ5DPSZrYijQX5E8kg66moJ0PoO0UdGta3eKJ79a8hW9Ren
TK3Kj3yXCF+vLKzXXh0cm33N6N5FcCv3ERCKbDfv9brsMWks8T+RpMFa9cBhaS5/
UkBx/2y9ohsXE7MAWtc6HV5yTT0i+22sfG/uTZWnNlvb3CtkckoRYabUy2BOQ1ba
x9PzkYuibIWfSpouat6cQ74L/fS5+tQAd0oSaibTiOS/H5KbWzK6MOU4/TmLfDwI
kZDAzTb6JYcl3fC25A3/RIna9YanFlGIib6OVjyghWUA3d9fP9hqicOWa08zRT+b
am/1vceMFYYSYxcRdAKak7NVhrr7CwS/hfwQDzaG/MegqY7BaEYPtfRUj9A85eQ0
wkJiH5cFsqY1w7fo3VqHrnZL7Cz7gGEkkLml9fEyG8+eXXx4WpXbBQ+vZ830QKmE
FCpeRHHN+2x8RA15kDXfAjvXH9tj/xm2WvfT0en79Fe1JTNp17JEjnkcg3aRNmvY
JY+FyGx5MFC3uvGJDVMLTSb7B9yODum6II9ygWsaye+ZmWdvsvzvJkFnAcfoUPiQ
yzwUM2oOTJMVHs2gHgYT7W6TqVXGjzabRaqGyX6TJ0VbLVddAQVEIBBBloKDQlnl
L5cIQX6bvHdVaqF7hFlMWq63yIt7m/qxvmUDhy+GOKkYAaPCaLPfI63xxVCkzqgh
glhuihvkKVD0bRBuRIpObn0o2V3f233drsEsa+IpJuOikUaf724glNcXzittBH1E
MfGWJLqVhGCzwAgY0hUZ3yNVfsdJrEV6DykRIO392V9/QfmbOMO5aWtcWrYssWWR
3rak8G/YbsvB3eI61sMNaDDY81bKe8xad5U++4GBC0nfP1K3G4JNXNTtTaQ/pDX1
CdMLzZadcCn9m9k5xXHp66ghN84ObjJFoWbz9jaUldztsI1AqpBEQz+jJz5d+X8Y
ttGpN0gCO14lDhXZtcgF1lqr7OFn1WV7MdWR6Y9+lTm8ub2Chp0XvT5rVaRZreG+
OSvzYdJHhbzVPUWPpyzv7OkWAP3Or/nVmMt+FSqG2CMo+yh419mosyuQUicDhIgy
sGbnbKG/hsODyrsQpxde9R+GNrKAB0WrMra2y30sIYk7Pv4ONqDfW3omHc5uECEB
dpw/CF8C2UB+i4LEJzsi+v/1ZAlarkPjqS2Hj1VfBUQi07pXM3h5cTtB5n/XXIqE
EbyM2SxmLd7SNqPtXrybRinNvdETEkc8K2Tyf2m5OAW65WjQcv0W4XYEBteeYp4/
Ih7cNx3My7RGHTnWcZ9ez+A8wV0pQTWfk8aUqAKnkFLQuCiHtovIXZsvHsCUkQvI
oF/Crm3lwJf2lGUKuSPQatQr2k8EYtHCO7tcLkBSkWPJz8dimcvOSZx3m2YJxp2y
fsUFrhUU+e5fxwgH/JTGvGZYRgGXHsIDlIHTKQdT9Q7g4Jx/Jvf7MaoqDiP6HmEC
i5O2+EZMZxK2Qo/wPaNRGbnc53AC0POp5OZaUSqybh9ppd15Ut18fg0WZLgQWedA
JDM7dHSyQvpA/qHIClmKTT+mkNgyF17p/oFDhicy3L0GZ912SESE4XzNkEtJNE9K
mejUMRdOQb3cw+OjToMwFovvMojxw+o+70iGkzDCS9/xMVm2oIuA0W8RjDTYK3tG
7YiIkoXE7mgQZt1mLD2EJI1DllPydXTSG0ZO8+Go7w3i01vggqk9FhGBQnzbToo8
7EUt5KbUhv5grLguRZZHcEVzIV/0ge38PnP09oiEqNWHu+bhih0uGXF3IC+3ehZW
HZWWjeV7juC7BOKhZTs7yz/cWlyj1jB+lzPvhvjBHSrvjF+SejLFZUsWRJLK2hT2
TrUlfLv64TqPlATRrCWlKPbwVsLfTLsBszVpY0yOpKFFLctG1TcnYuEnmHqViqOq
P+8GbWEAm7RFeHwt9jLRb2sTyHM86bBFqb+YCKHqLCytS60cxXX/uIGrXcT4xzDz
T0zgx+O1BY+QandP+OqGSxDmTutW0gDeBsKtQc6/JMXUNQYAVEUSx7XFRPgqCyTA
2cbbzK8/JGgifnRCnXhQvNciSRqxk4a7ZlBsWP0RbSuL1GZIFv8ybBKK+Z8FS522
ytCGh9kn5H6RlWabZHCDrfwD4p10JjlOeGn8J8yU9pWsZZMIYfKykjRuMhREWJwr
5siUL1JoLCPb6n+Y2xVzXD+hcFeJkwOGxVaQEzzgsXTnhXX/fSWnaa8nY4ZWCPyd
JKbula+D8PAAsLRIh4UTY+CUNfetvLFOaQnpq3NnMSvqNlUb4xnVbbRD3mqZClfY
870Ijxg1qk67Tgd3d4Ylw9Df4bxHq8+lSxoDeBIhToGbtF5a9Om9LycKHMKCk5d7
CbZn4u3VAEM5GniZH6K0b6UrsOPAenfJJ8QLqBnIEdPrq2eBbdXAUZtrQ79vkXDW
TjODAv0U/EHVBALXPanx+gx6I8yjD+We+S98KrtMP7hm1SPO5OFMV50Qv4zd77NX
KfqB5bFPKiK2IFjUqw5wY+awiOxxvOTpQ987HmLPhx/91YyUJ6BVMdBBUTQpGqQr
sNc9PdTZRO+notXhBqmVEA46U7KNEamtiubMFdhy83r4AJmYkFzzeSBg4OZVTdeK
8Sr4Q44ey9k1gX4l9nsq/WCyMK2vcfgEchPyFuoDZdxRGkIvKxj6JmiDB0CRjWFV
EYO3zfTCU+tpiNeNe3feM34DrSA+ZFtS0pTLbC1vcCFVh8NvVPmk9zh94d57ROLb
++iLEv7nIdlqQA2xUNUEZvZmhfRlESsRqpDZt2I7Lw98UhxYW+9tC1bdiFtatrqm
KG3/J044fgEdXfTDbbSQKWYdyFK0zfA6Xw0RPz3LnUnTYBCJ+KXd/mUYWzNCn9lO
EhNTb6oQO6ZOuaU53+eXMXQ+qkkE4Zy+OFaTA0zcjFNNNn+8yXq8mEBEN5mgM+VC
wggYVYKSgyrWHgicmqJ1inhNXEqwUAf1V0Mwd0+7mox331oV+SnI0joi7mTBl5R+
1LIQ58RxTH8+pAJMTd5yr1tBXlbe9yTXxN6JYzTk8t+PtPaohjFZo9CdE/gQ2q6M
ck14Oo6M4Adl5JjOqRts/8e1Ie2YZqyIWO6sp+u+Af0znQ4/QIkyMN/aU/rCOGxb
R7Yn5bhL1TWIjTpnoVUifaVo5700wxq3Y6BkKdgObgyZV60+TqFqJFHd4ZzOwxTG
dJtcwXHZiIH6werrq6c9X6alRpXLWE9Pl8daQSJzwL0bUSQuddoHrsunIYZDH+tN
4w1VWuY14TSFbQApFd8b4k2agdE+h6SKB8VeDoFfWRxJVhN1o0Q9kxYRlsl7NImF
RXdG/CbMYY/x2xHTwx0MYt5kawmmvsfQbhByjNOl0iUQfF7E0hGanTcyJEQ8AGrs
EoUImr3nRRW2kPyigyLxuoI7lzDwZMIyTnnK8ZDN+U1P1fz02Okdwg6qKPUNiw3o
Sny1SdmHJwFHzzsQWNyB32xHbozFdj2Qq3xnAAUJNIYYc8HYIwlrQx25KciKyMWo
fOcCnhMxNhYpObvzP1fa6I9qIxXzuyHhjDrT2k8IJquB30dRlm2FSJ4cx0ZJ+BJ4
TkJGr4E9iXtfSFkp4JwXMb6Pe8Qk9HxOWC754Ou5Y6crZY6u7gpnNGV7an4EULJv
CZ6TnYsNEPV8c08UD4gUaFzME+b5KyQ2BTKh9xBHIflGmNWHKlb2+muInJcNlyO4
6pegXzAqDWxiBPkcG0GgPdW4Z5LVwkTxlMk2s28Rqe28vjfxstvGXMwrEZ7/CB9t
ZKPCXCAwLN/eOngbmqYLrECOU3uiGKLCFQYMxdQoZFkqkLj5ZcS/IthKAVJpkdaq
NA3BswIkCGH6zqPfy1dhmJHnqIHg7eto++CWp1TbKbgxD3C/jC5ZSqrV0xmANz8R
KeR4VJep+CN5TixrsdJtbnGEFoeQvhGY6zpDg6ibcLgyghPGezTksjX4KLsMRDzH
+wMtMufldq3MskQ2EbMZ6lDvlyNejBJH/jG5tPVWON4mH9nL5ry5633dU5r26glr
wPfw+8CCzZUa2vabf08gc0KQ3m3z5mY7w0OBuwkWNNO66cAzKhofGRsFVorRF2hB
HmK5XYmARCPi87Wp++ggqJVBGmv8JyBZ0Pi60niXDMJv/gWbsZDI6rXGo//pbWTa
v9jCary3quYhuQ+sVQaDh4+7yF6wI7682G57i8wXAsJ7jM7hK0mzqmiyZ7poio/H
i/Vg4ee7BJfCD9TtN11I0EejM5ZsZ2bePEz0EqbwCayXyKazy0uqb6y4dyTm7qZM
wFvBbGI7m7KoZOe4DE86xtVnATCPI+EEkabugpdO2xVFPQLFFg/e/gtLCQDpEkFw
tcWgKwu6BgPhPSQJ+KZ2EmfGseito2+OaNpZofDEfrcEzeePeYBVgCDf/3X+H8Tw
rju7WpPs3hEPefVL3rLN4DkrWD+SK3yZBUjsarECj0s0kdpmMv7CktsQ0M92+gMM
mujLu89sPVCIZfda2KagICUBoZgnyuBVATcJUmy0KmUiecywYUlBBj8eT3M7L6TM
1JWdhccRp3k8UCxCjLStcRubYxgvjcs2j41CG1mEJFHjHcXXOk4ZTSWbVqJfKaWK
xNrWu5K3iL46G9hzPBkPfcaom5qZZOV/kYxUGbJgzasDOUEy3NB1oGLInB4LFOM4
2nLVWuEbhNw3LbndmUxZ1WqIEbr7kAciE+t/9r9hrcXfVE8ShUQtC66Vc+b59Wi3
bKJn3KM0UI2Ve7aAkMv2Suo1/efTWUKGYCAXBAhGZElW8e0bkwzckxpLloMPMu8k
NiZAgDcXE+GPMW7KKsDOUpwRGbyoVXaW/v6qBvpE5fIV1eHvw+YB8pifBbvuHStv
BqNsenKpHW5084etkUI4l5r+KwAn9Ouy4JBJ4O6b1kCqbQNyfLi+yF6FEl5Zfh4u
EPLMnO9qkSdTo+tW39TZcQnEGt0e3Zlbk3tmrkswCBaOESPaNIpQy5WApn68Tvnu
hYuvZVVQH46Nv5948ID7T5H1WwFZ+0tXCimtTdNacC5QlumGQbv123/jtPYLdLcf
2SUTV7ex7IkOUYQSU35X5qJi83AeWKcT9GUZUZPE+FBomv2iv3Um1EdOzwpOXNPo
YHWaNaxjCZTqHlj9OviCUepUR+gR9LaQbw5dX46CJhRc8ElYATiBXzbYSascddjg
Q31ZsToX5O2zoKrqNz0TKtOzx1AIoxNh1JLAK26iVWwxBSLi50+lRjAlHDpKrOfP
rDxJvDrvj9rCc5/GgEmE23O53tP/jU/9qD62vSwcLKe+ZTGn51hlZHg2VQOc71yb
23eJSFwYtj0MM1lkvpWs1iY3BsCueokPsgRFbNzebDev5d1q7S9KOwkWpLijk4YS
ft16iBHUNtt0taiYcnmTZxMsJl8/vD50mky9uZ8l7ZFzYjigzjrwxRkJJrmrAOlD
xOyaMa7nwu4uNgmmKLtvc6T9DtZdwixnY2oGYem1KrD4px9I+WskOeNpENwNaOzz
/Pm+iAU+2AL23Yh4fazis6PJhRjz3K/mzHZyOjW0RSZdrDyx74T3wN42Z6osPWx8
7dABVcItn+Ab8OHoX651YLTs3IGM5+sIoQ8Jz3H9n/PFITXl8zzie3smvmgv63D2
4+FFIyE0SQC9TqZr2zzbI6WR/oAU67ogxnsQcAoWisgiv+PXUiRRCx72GH+XXEv5
hWlYaf4FxnS9/OifQQGg0AQm9WJS1322zH+oOHXTTJo+1WK2tci3fifRmROVOmok
VlWqFuWK2YqSLvHMl5BhU7k5/iR/hkyHgcGcFJyJMzhIig8CHYiwYkbAQL5nvvBo
lrvCAITLnguw7UfJw/jGivjO9Jr3LrBgytsJZDOzGxURhB/WLUO6KMRwub/vBmPa
/oW3/633l7ibdcfx4W40t6+1gV8hDXeQJWIeQUO8bqErDDmXMq41NjgVR0Bq+Ifc
srvWKbTC6YjXIw2FRUQv2DzvhxxCSTGC65Oq1SSk67QJGkJBZRNZ8Va9wh6ryvN4
x4BQ17F+bJ8PJpbvcQcfZQoO1lMEt6kTXP+MOpNF5jFVIefWDdvamD6FoMdDLWfF
TlpUv9uKm9rGLeSbRh+j2NytfYxNN1Gb7/X0QnsMqKMb/sSAWow0iq7JJK1TL41y
6hGpwagL7qR1OH5rn6C8wX8O2yKB1avzugMkmRGEaVs2rRKxft/iw75smIm4npCP
dWRohBmLMLQ7HjJFDgPah61kjP7VkDnB6x9/3SVnvYAVsH4xai6gvWgZoe79wr5H
zU2wFvriDooRTTFF8k0UqMJdRZUAMOVrB73Vm+0XgFXAHZOHcqyAcXwm9P8JF9TZ
sq5sNAnos5LYt8BjeRetR6h+Qe4WLpgCrtaDaqdZN6QI812Y+2X2w5sN2vQ+jPgX
4CfuYycERduCaOXNrMBplLJxAqYPYWIFBhG9IY9rnV5UU8NMkoi2KMTUhrseu31q
NoTauHFqNOMmfKE4sb9MmIJoMvowS6Lc61UweILeF8P5GMMPaUqI/g+XQq4htpJK
WV5Tl6CA4S5iX6WK8C3+GcMQBDihhniNTuIWl4/mR+WX7bEP3tD4LC1dX8Ms38p+
bcHOEL/lf+BqtPhr/U1X6K+hEQ3IMZiB5iSjlrxq3sJ8qyt8nknx/Oo9QuUBLNet
/ICFGDFtLN1qDq6yfdobeLtLUiKRDk95GoCP0H9VYQo50l5s+hmLnUGnVYe2AA6w
3xcOhFb3qn59SKR3C8rXOFUvzL/etrRYUcyNSIqSp+FjHrCRfCMKyQlb5VW1NVUU
3bGsNe67brO9eV5MIXObvY/tGlnD9EI6WA07usmgDh1wC5WI4lLyXn+SpOeaaQDn
tiExYt3SjobwuzH6uQxijefvhEMdLZpn7DkFD3BDbKLs2D3UcJ0VtdYHZOi573NL
GTsP9vFIpYKiEeG4mSUHzLnqPazMkDx6IvpsyxE1yC40KHBf9K4KFzWvgBwic97U
lWAH3h5pHqyLxaxaEkuqLE6fMOz4418m5RjcE8xFrosGinHJVp5duq8D4p+wzbrt
4pZb5AJ+x0Se813f+3bSiFhL8Z6Wi3nGLDA4GEvag4CZ95F8uPknEVDewQWqZ52K
0IU4q0+Idh+mEHu6Qwu3qXCwroIf82o4XtTKZbiXkLjzdIhWCOtWfIWnlJPCK3Az
AGqE/fF7I4kJH1EMkSiZs14jYOzvFmP/VtWIMFrW8oon1Au82J3W8CMjeDKKkJ/3
EAIjWaDFvC66EAzYaxl+jI0AtC2imC+UZCdPM0LRrkllfD8bUle3CANysvBVjC/T
G2Vv+4EhfcNwnLJoZnuc193iEBaLHrwDIh39XAnDoB2eijXJZ7/irV+3Rm8JjnK2
f5UBxu03eOgF6F6NydXrgkhmiEc0xlJkzKj4EsSQLsfGDvRMjxa7NmL5g69mnR/I
PP0zsNlyH0RElZ3vbVgekmhPmZOKdCzm4E9ml5nYJuaLB3Ce83p6OydY6gzoBnB4
8kikKpJmr2A4iriSG5EWTB/E50G6MBgESWfm+zyCS1CRNMd1zO7K/9RbAsFCGGtT
+bNtEuFCQH3ZIpKEJH8rUQJY3CS90awyJilyB6b0PkuyH6J9Y5zHE51IsrzvyIwu
EIQru6zIKNE1sedGYYEswNDO8cpguFsy42uJ0nGSr7jWuuwJ1Z13piDIO+LtrhWS
nU/T7FejBqUoSNOPhtzuY/9xwzgxPowytf5KmrGdHYyovsMaUW5EDVMNQWzqTQ14
yB/KjW/O9/YFOVCmd7auR9B7iBjWGds+YvGxmu+o8WFeGyghTVb7ul7EM+d20z3t
FzaMa4WhVJoivRIFcqM2eM2SGWtX2io2cnB/sbCk7uJOK0XTdXrsS2TiAgnb7KFi
V8tJuB0z38VFLTv01E3cYq6OOHxOVeTxUDfli0HCTB7/t0enJKGF9NWkyT4/2cfF
O3+cXB698UHcVhRQC0MkkZ2/hGnRUZgsU89Qfc1ArDieltqWqR47By0LDgpsDy+Y
oS8EV1r+Oq3aLGyCxxU6bOCQkoxonEzZRAr+Nbago6srnQO8kLWjQn9k2hYTjWKY
+MhwBnFuVXa9N+oAT6+8B16A5HWN2FlNvlmtpW5pTT1WHVsvc2Bb05xDpsOimdYC
dMmSPjAQcoDZMq5vDdla2P891bFepGIXK05wvQA5o/trGae7AGsetVH6jSR+Cz8S
Sb8wOqdYT2k4vOioC+52tYefcFuh+W5daxdRrSVOtSvMB1ujmsyrLndXV+rGnUPE
l6KHt/hVUk631I0I+vAXlsdYHGdL/tyF6OWB2wotkXOMsw2cKAlWQMaV8hLJIfot
QWP4x649n99EadlfKRjOeZDtZDeM5yAEtKGF+cYkb47awP+dJmRcFz8tyECp3xVA
VTq6Ht4gXRFZSlSILbAXCXvOovEo6YJYRRGzDCO/rtvnH4Xrksrab0gVUj7xmkRj
8L3zQLOQZUL0webw9FXkSO1QKNF5rWO1/DYqmSuQWZSq62UcdwVfxfVthL1/sQzp
EVR0p/30dy5BgiyeKZn1hw4nWD6Yn2+abbGJcDfE+4GQzZa3tqckM+h5a0AzIf/v
chH0ihDnNcIvWxCsFfDWWQmeM8pNNkX3ng/INLSCStAeEIN+r54n3ZK9ttrFH9LY
w8FqotWafdgdVOYfARgUYL+6K0sD1NnkZiieLM7B56R62H2bEQYHwqmnKqk75hjb
SbuuxmnZDYpCDrMRJcQGfBKwiPlFY2YaKKHMeGDJSvfwL++1APx1fs/XuXb9ITa8
U5wpQgHLJmBWOKnHq3pcqBbiwoLznmTxsWrcU+b4wyIJ7UAWf22hzbm96V4hw16O
lGkRvCgLKHwh0uvewfbt2pLOtBIXUjKnilBgv7JNZzZ0efvKs6fEx+cq5ovDSYrX
Xz75ETvsZ4KZ8aCegPhzhLKz0/IC4U8p8cSJHud8wQvKWye2EzKsaR5Ju/LlZ5F3
I2JZv9ZAqkT8pBQGieO848Ii6vDswiNCifof8sqe6s2vnqD2xOornaEZCP0NOk4X
h5g9WZjjQRZa4Y17UfQNytjoqS3+t7pO1wSi7XrDoq34cVflYcNdJUivadMGIUZz
eee9n2Fu5q9ec/zJksP5kpepCqHXXsVkXyDPopnuQudmaIk6so1u42Nyx/Pew72v
fVLbd08wiviulXa6sdvONW1JhJZ17MMErNAWSQjAtBuQ/4AQkOq3BTkPgQr+6WnN
fvTxxRASF7j2fvqdJ1mkagdMVgSf+chL90lNbgHiy2pAWVniCwI2a9c82j5V1DUN
tQq4e/GfE5l5hHlxb5VmjOP+AF+FY/hQzv7DEuYLlIdHgdFnMMc78NAjmlryLzJw
NOhfnNJjoBRH7fIiZAgBaYpp+2SyfK4c5I1nVG9Gu14UTwLf1QcCdGMrAL3apEH/
Ow/Co3YyzOPYTWexYatVmXfqZZQyb4EOaiWTvqQRnlCK+SHV95TWDE9FmbXlJkpD
e5gfN7Z+sEMo7jXeNLyHbZBSdgxKk20xwvJh/Gq0SYA/eL/kDFKzuZgTUp2vBE79
zYciTdVmbImX4mbKYFcXeTuxnVnwjOJI1c0aKfyeHze4PiIfb2vTUpvEMRkKIGRH
OGrHaMemPW3Xxm7MDbno4XKxgExsPiBnhWxvI0sgmVTNt5azObCBnoOVUFyDkRXy
Jyj4ekJoDB6BoEeXUBJIawmPVc3Ki+K+qqKwhO5cdtRDipp0YhHbOESDzh7b+Nvr
SDLrF4ovJ0wafVXBWAvs4zZtTiutEBQFDzXG+a2qy+2a66xEQYQdi8LpxRXx4mzk
xNEd+6efkzMZ8Oqk58x3y57fcST/xgIsWBCzETXDTSm9WPdIZYwOa6JGxj6YuTqW
5meTs2nSqD63WZmgIDnITZ3sun8T7l1XKZAkMJQKNMrmR9tUxHWpKT5mGTvV2nxH
yBs5E/ILJQa336G4fTn0bCP4RP7phhe0pXYLkenDwXCQDMAtDTqeS5Zars7pfgIv
BNDaoJPEXoiz0BOmW/pUQcSSnSA3FNekYm2jfvrLKk6oPm7YyY9etRGrVaWItsmB
zksXCCYRDKH5vsAfbZ+Eufr+TbEo/kRrZcGbd6qEouQpJKTdoWsiERXRmxVO4riH
e7HXlJy+lKFMmWIIbssNqOZw+FeDr3X8jsfaYJeNaQuV0B0fO23eL6mjh2fibqNe
htCLDGtEMoqlroHF2mT8ENIWTJvJOTpIyPHk4ppS3MvcMnI1bYP8JmHtySzg3yNd
W1Uv3f+RumqLlmpq9GT4G57jj/2PWcCESMMD+9kedEdBVR+waB/+CuMXevHd57cK
u4gBHhOowONwm2QFRfNX6ND4miQ5jfKAyg2xl2s3gdI/Uxlszpynew4j6ypduGmD
8YRc35xLSedIyB5/33bCQbZm5kwYuKLi737aNES0DeMLUsOdcFUz690cRtcRl5sy
ZZHIua1WcmqjjFL4TiyYM3gpdLLQFtsRbiWCOJ20ylCHDEffBk5EVre/5J/zChaW
Jq8z1DzjclQqsHVW5XqVnDPtd66NCMXEJo0b+bVMeR09DLGzCZEAsqoCksKR8shO
QJRlLtgzERN6UfrEwjs7sqK28XUMe7vwAJGVA0r2X4H+yLoqlL8slGmDwAsEt6fw
ELjeBV/S60GgjrYzHlwHXmNA84+2vlv9gKUQYppdGuBZqKEd8EIWecwe/WSbyWKe
mcMkmR/D+RWaDMXzNRVWVPg9TeX2j+d9Y7GePGTOb/iFdHeoV5fP5QkR/gv729S9
24FkYxAUG32DEdYTZlEpA27Z/ywMCLJVJ64HJE9ybUGPYyXexhwdJwHWBcNX/v7P
J/Bl4mDCpluQuWqQY7JVWnUkVAXHpbNYsGNbfGaa2pzNFMADFQXAf0Zqlg4iElZN
accKiVTgiPiTLdS391pA6ag3D+Ck0OrH3AUvGzqBsjr+p9p2A1h5waqnfPnD2ZsY
/CNTpr1JMMlNJLR1Snrf3BjqolY+QSKdVk7AvQV+Y0p4z15TnNvEqQB0tF8hcBe1
wfGmP/9hl42bDSTx7UX3LiqgT/45+PI5kNpPi/dlKLJ7xE/uh1qW7A5ofVlpu3o/
/ghFxRoTTJWkVKL1vFVVj48Buh1FpZqkR5T9lEhwVTDlMCPb/uouMlQzPE2MAokq
qGwBhtRGlIwJgUk+Yr557RpvYVe1o7KW5DHcqI+C/HSqLICJUSeAzUmNSVi9amIE
Y3ebv5LRBJmE7D7MOp63vy5s80tJn9wJsahzNdeETaoAjfxXpGKRPuLgNgUiKbfP
eNYtXfFNjnJOtff84mUAglyrXY5jxA/GdwTvbrWEKwE8R53tWZIeXKlDVymSRMLD
pTkCY0FMB0epU5JKj7+57nril5IjyhzPRERcpQbldrf7FsPvTSCeuxmRAuZGMFO5
bG4f5LzCoO/w1VhNxxEsG4Ht6tGrn66TTM4YhMYHvEzfWRgkTsLnPijTMY3wtmXC
59dd3HDdG2kVl4W2Y6na26nvVQtRv8kzpuYvZs5dLByPxXzCAc9j1kEQEsxTdc25
MALUEi2wX4LpYcYG+/UoCo9Qh19729QESZrSPHzdnC9Z5bHTa/9MJwGA9RY6pGzp
SAf0LcSCJBpQ7a/lDLywE/ExEa0tgDqv8Bgbp4JEwAgTbX4aYie4CuopVCCf/aAJ
OTKfunP8IVlUQ+PL4ZAxXmpwAbkVtoM2MBgAHzfED5VdoZsfKlHNyHNSHRpqHsjU
JB5vbT52yDXzluavrNdcMCB4cXvft+tBlLiELzI/hEW2Yv+F7kRrmaxv+lRPfcC6
lF3h8p+bQW8a22Jcvnef9vTjmTyjN6LC8/eTdKKYSRusjj8vkHyf8MmgPAEuAUfk
+EHlnvZK/KfNHLJVz47qxWIXFAJfzmPlq/3q52NOfSd+BRW1T3ifO+Nn9DhL+ool
Fpf/SSmqiyNkd0GzeqIIqXcpvfvj+8MWNXTFZC3wFImC8j3vUzi2vzV+dAC44WlQ
aSKNqhlAtNVxJwTuLniklMKusJkGfhY4h4eYCOkP2Uf6Ujgt3tnZ9eS2FlosW4yD
xOZ91ywrUSuAic5RAHHWcQZkC+1MARyBsUKVQq43ThSTDe7H81pOgXwkZ93UpFft
hQ+YAl28ZOllNv3ITjKp7oSOR07E/WpQHGWH25GFeeeRBHXw39rNYXd7+J07vtDi
PegBziZAhg8oSA2/NlcllCPQq71NVbaTMpzH5e1SABMX9xH05/r3eUr5dRx/PAHZ
mr6Roh4PgsgBylnOuPCUgGwpnmQgYG8uZbdv9W+vIzCszv7NcGkFcsdKt5ZFEGak
wluKFQ43tKYenvivJ31yIM9WU1Zs5q6wM/euz7scWwCopBhg3OWNf6GZ3zvJ+zZB
nCLMvWMfPgQKTWUWJmUaZqnuEG7VcSYZhqLYlCwTzsGzwp8y7U+sunySsa7+GF14
n3ZeOL0kpww2fqzEBTtnOnlQi2dL4H4bVmcmUoFkrv5+vRP7AVnPQjZOF5FFTvUW
5jk18SuRnEU/aUKDtXdtOjFBxIcx/mwY9ACOGTfREhvPSGDrQDEWzJjkoUwcJlnV
0YcEt+vx6N5yNb7qwCeD/s/5CjiYLZdx8bto6lvxrzb5ofN6LP/BRlZUhRiJbemB
CTzRTvsdEmb5HUOLm0hN3/hfDrnjOu2de4AADywavD7LE2fJqLuIajj1GhlInwfS
vEFEZ+56gPVJmOTlaXKKennke3E+mZc9xqzx4kEGK34WZ+8su25n+1vL+9BVnHxr
eSa1iHCGEejx3nNpr8F1gXxf0is6u0hlOo8JquAjXHRopkHPRZbZ6av4+GYtsqqD
+LDxVGdEW59jZtHBTrzpXoWwy11q06zqXnlDEwf5MJFohrLCag8RKPoNm2IbUZG8
mK/MVqs8aEw+Dt53JP/mnN7NogGqHoGqUO/u60TBMM/+nV05KY+kmNX+gLj1xFCy
Z1dcH5g/kmQ+zrcIL8Ic+dQ06qj3bUooR5LRjcnnqUFca7l1lPmhvnFuEtepmeHQ
SqyRba5+zBiFYa2UH7ilz8Ay2/BxahXOGChij3SHJKWbsELxyAQUEJO3M3qAU1Ag
hiMz1hdu2tPtXlmLeJccLJ/24k4UXL6yLWj9b101mokoPj/VD5nkkpg4S8OidUQE
KSbdBDG1d8h5yvhX9UgQ9gvBsOB0VVtFlAfeow+5Yp+6Yxszg/MA4qRp90n2nl+B
AcPtC6S4kGKI4M8pd2Al0DgRb/VZLwNBE3sOr6meoD2TdiLDzOwPRCAXfvVYtJ/v
vJqBazj1zKamiTNrQzgf51Qk3u/H20q4+eMc0ubw7lFvAUyHmMD09GDY19WZwP1X
qf3kJANgKgQXGKduA0Rf7KR1BVpa29UzzXhTXrfk1WJ+Kakxhj6uhAj+M3KLOPt7
vUzowUql5i3sMlNPpct56VED8VLl0yRTIfO8R03q5cySnJwQG50AKqlj6K5MOn6O
4ZqDh2Rs/K/JQNB1ZqnuKalM7E7iSJ8VOnGjS+DmAEBTBGEC0i1meLARh9DS35A2
FtLlGgep9s6nLKCJQqPcJz5WL0lzR4AoLZmIovH5XF3/2kFLZvOM0wloLCewfIQw
Hf6OmmizwdbTV+LgzSSRXxwm4CGm/8a5WxIB42f2bxmLvybSuE90uOZAD2zzKbZN
PW1YdKwbHXx3d/mZ61SSVErcOu/2qtBEzL5YNcNrbA4cet2Ekkp12pyWRf8u9UBa
vzZpmdlt00Hu6NmIHPosI/rGHxFAmNC6gruIv56oRyiJrcHs6Vfq+Vx02ZKpX6JN
VX7c8SJi2EqPik0NdnH2V1UH0Gz/islEMn9/lxJGVgRyTZatWlp+fWutTDCMfcDK
EzHEcmkDi2ECu3jFOurn/TU1scoSaZimni5OM/tktOkWZxzi1SoBlRJrYX97tAjW
vX+gyWXiAmEsoiPE4rP99XNki9pliTwtXb31+MFcPpHPq8zTo0YmrclJ2X/2sFgD
/SSwo5GrzV9/zA4RoISd+ioyaNRdozllyK+ZTeQq+Xdy+PdHEE/qtAZSTqG/cClM
8zEdoFRmrKCRoe44GeE/3kPxlsd4vk8uPcSyQ3leytOK2Zeq7oItBRchBkGkrusB
DJNxPthutNl6UpB820cjPMp0q9USV49+qTKTXFTgcWoywZmnTrI3XJmXJI3HEpVl
l4Dxi9bMOyzHMjMsJk6PWJcWjLvOQMeJl/fIWF4n5HgPbkTViBIm2giyWos+Xiy+
4s6HbftBmg0cg7GI5lIfp8gg/EkXrSOSX0eWLzVEvwdlTF3RAnYMgdt7EhqIhJrN
NhwH7hncoau/Pk6IPwI+k1xjFQqJmZAHWU4E+uZmru7hcwT86cEoWQUniSAqrIKC
ip/5S7kTy9t2GVwXZEoztXsaiQcMiKbWw2QjE1x2MD3exB4CsvnYptYNLdKjegl/
MMTY0hEdQEj/kehLW9Bp77p73TavFLbT1g481xgcU2StLRlRc9twRvFCqbQIwG1S
IcW7bZZHZcaj3VboBMMF4cfEaoLqOvU5R7AmAt74LUqnLbTHtNkIWUncPuoGUEzT
XeYmooD6EwKpCkKT/eYWTUh4zj+q+zDA1/SDMmwGrEVmfP342jq68wyenW6RCum4
yn150y49m7pBUmXt3gt0eErv5u5XwD+S5FMxb3nEDnEwjFqtltjtMVGGAdw9bljT
fpeUfvB2oHGP6RO7O6l4Jo4PGiPMJvjKumFugNqKKmntjy0kzS4aD1tP/RjF99qw
2h3By7TBJXCRoqqqMnVtQpNad7AuI6l7oNPkefGdckZcfC2YhsYWPBafnTsQ8gYj
VuZfoz0R3Qm2W1wojCeldPHTaIPBpel8ySSbkU+aMOAW73ctP1mJM+aZLGLFgjl7
GaVndOuJX10p4xZ8zs2vh1YDQ4rbeh6o3q6b+HY76cBLzshtPtN0G2nC/G0X98aR
1spCmjNOp3txZUV0ecC1Le81SJqaXioZ0AQJLPGxs0xRJQ63O0IyOBSOQ55jcdDM
ZrDqF3T3KB0H6zNfucfUZVkuiLOS/1FHeFEZwuUZVOEj0f+d5REl5TQifE9HBY+w
St9HrRsm4hJU8+v2ro2/FOwwvrEpW58noYcyloPG4QSvSac3mKR2WMtcP5dcPqu6
B1MjeJo3sNZcofjbsmF7Ji282Pi3BothUcXfHqikEwbOngcR2FB94R3Q3ZZ9Eo/+
bUsjoTZbd3C5rMGiw2JPCAiymQwX4zXWgla5PAhf6x8U8zms1zgXvOnnqQqS3O3/
7br7zIFZFTF4YEiAbEnz9mN2hAG3+A4EYO7oDIEKxuXH5JcdjnqHdVaK+lUqoxki
/p8wXk82DNq+z6d64yojJIAPKeAnPLnT7Ige+1m09CfR6IaLuf/cUzi/QQ4VCLG0
xiIGD1jKvk7nBhRN/gfFUP9kMNcFhx9KfWQhtcuDAMhXLKtVbxJceGBIbHl6IF3c
SEyivv9dY8PbEX8Lttjb48NKwJ/dzTiLEo02WEOV78b2Jas0NELYZtprg8jfhIz6
tUCygQIHFJ1Qe0VIbpwqtEMPcEma21bheNWPR2gXHaHQaQ+4dcyOu1LDwR0KDw9d
Jf+50Kw33j5nSqaiCH2/PzrQy1XUTpR8TQcwz2dBTR5XEa0xN8G/8QHYxWG4nnLA
j9+rWje7miPSCaH4CIouLmtALjs88iv3VwGMMSIfeFHXOMbnHpIgxWhBiefoA8Zs
iueJghX8PYaguztFpwXwoyyrFNVOSbJwOs5viHLZxkLh4Xcwtt6n7W0HammDYQ9v
m7VDWDGhFp2omhkreMcpMyOy/3A1MDv4ryJAlw7AqWEn6uY0r+xOkXV2t9+SNhGV
uhpWqMB8EbG6bfmrfXgOYw/wUp1Ntb6DUDJS3UChTxc+2Arv4ftU6WcQrdGzz12F
wh+EtjxYogVd9bxhh52+k8UfW+Hgtoh+oH3yxJRk1/lTOBL6uv2JwFJ6Wktu51QF
Drxm+68Th7lNEoTI7HEGIYG+6P/lQlWgDEzZrnHU3HEIs3ISPGP8s3ZxurDubKG/
F7wEdQNJGT5C/khYgcXpasNX+EDTJCID5gvJvWVFWF1etLoaK0BS2RLE6RILJvRj
DZZ1eIKzRnsm2sHuNkAhapiguv2xuqm3BxFikHv6e0SjqzxjzHyrXSAdo5gGmwbA
uFXrPtieDVPa/IJXXSKwGjmdnSitZrZsvIWmhOwEztWjf8cJHBB71Q0u+B61j7T8
8riiQS+loO4350g7+y+WJ1YnN7GD6xHmiWK0NOcqcGotpdLO0Z5mbupzvQHWjRDr
M/TEaEga4Fe/UDwSd+HJbf3LMvqff4sJ9FWea6BB8LlFwubvZ7xs3ejzsmUW+iTn
62Qi7S4yWf2r1Zu6TP7QhnZcGZxQbaqO9niT7kalUS3s4Qiy6dRd4QkvPsfrHBoj
FmTfM1cBQHrzP9wdbF0jMzzimjtZJ2QqsNHtbkVlAqbkDyxXqBNsC98lR/vUmAd/
kAeX/wVUFhpDfbiJ+PYgwTbos8ebVIW4Qf+ZNlq16hZb9LatcHuXJ0q+lKe+R3wq
vPE8ySGPfx8dg0U/ejPwSLxh81mU9NZuogqCREZUsGzztlZAhxL+kn3QCYtwZP/4
+07VHZ34tuE2EpPyaSK18S3rxhHbH93gGkbgdJeuAphmH5IsSpMkPkR0FqcU2beu
Pz1op1aJr79F7OoVP2sQV01wkrnGonFRleUHsTHrer3mpQ66cUoJBNikph+h51Fz
K7ERo/IiBVpAdbmDRwfcmSACjDG8F2NQay4BSdJiP0BN8LukwI2LxcuhTThU67FZ
sLdUD9Bfg4/D1mWc9BsHHKS8u6iVvypRaZHzkImsrkGwqQAteWedyxo85OHmr7tm
nRobk7knVmFgl/QLOD3JemthKXlYSAutXEF6WwUUeAx/VpmYZLd7Mm+jSoHRmK0N
7slHLOjbvOyd6YOe9xcZ3u7w4lzKbL1YM9hJWQ5P8r+nWfiiYoS6PlXEBNyztjJ+
rjnwceWp1xkKRaeQlYkpbanpAbgm8RUQf9gqsYkmNzP6mFBcc6lO6JcALthbtmFZ
arxGIJEzXmySFv1nPIyK4Ui8rny+ap5z5GytALOVFpWdmZk2ckYCzEEcM/9z+1x0
B0ci1/G0d1KMkpdPDtkzS7SPPIkgxYLlc7+pZS1avc6drxOpulDU+KSOOStUUA6J
Ta6WNw8drgu8r7NFyzrk0lq2tpTUotue1yONHTQOEkV+TE8Q/JhGfv7EnSaskgys
AbVKYU4iantun+898lcIY8/oyyviKw8Kjb97ev9ARtmXhxB6vCa8iiB1ga8Tscgr
3Dl5eayYoZEn/Z9bBMg8uPuGYTO5lZ7LVSEWxpQ//zUwTiBBw29Jkw2PhudFIvQv
nYDzvvbsYf+q1C9vmiOIYTsfzxW8/l0PfCyCt53+nBO3WRAfkOIq0Lxbn9v8RHjA
FYCaN4kx6vx5zTgY/wZau2a19fAiGVqE1oad7XF6rE30YlluiSuWYtVQ9+l2osLV
eou62n/MxDBUhH29lE7NqDZ/2dnxEGsMfpAq6uiZfH+q2WhPJlNsGEKdrBnvJeFg
n1ShBLio+KoTm2OoCMWu/+UZSavXvXPVRo3JDBH0W+4ejg9xhhW2fvLNMaLja7kr
4W/sbsIyJtiUOpxaZrrRzMuIIH1WcglMWTiyl1J7RjEfVbYuIkEC9lNFbmzfCMI6
VtI+eHjHkb4WdTIOb9jqvL9D4WslP6izT2OMJeqPGeP8ayDTWeUuMANlq54Ui+zO
LIHoo8XeET1dtosx7UpNXlK3vuHmdlkY1xe6pKlr13YSErjXentXqzD9dspPUK2Z
f5cVDh13GsnPUxnESJEA9lbBGQOb/QrYPHvYjTZ8kkBbArzAQW0Dg3BC/74Y840B
Z9hjo8YqZP0XMEIqOeNh7k/URuBJpyB+ZxU2LXuqw6svFoSyCWhQUQa4WQsp5baY
okjUhLgvuRdZEM61Sci6cRs508ND7O/1syCvauH9sI/9qCcodJ0L2b0uQ1u3CwYB
arvgefqlaVlCQRMK6vmGSHBsO8TDkuqCkxkH3TSvA8fc0duUseFK/MuwbHyt/VDI
tHhHXxSQ2WZHLos1nymG8au6NCAGvK+E3rH5QXWjq8+T8dZ2SSJ6DzPZZI0C+XFk
aZxSDvaOQRkUX7VEPbL9Hfm43LXGb6J8Tg6DLGzawJtVwLUoxloICnt21vTvartJ
snERtekTJIykcVl2+qgw8Q3BWmFQS+Ku7auiDS+oEzkeerPugYH1UcaI+VYCSjSg
5r/+uItbtuOgNOXFxJzjaR7Q6MqQs9gXeUP46o1w9JMtkHRspAwvaYsrQWFStBJW
1w+vT9uI2OzoqGOAhI69CqImhaWTZDxyA0RjQsF74T94JDE32Tp33Iq+TRPP+9Hp
PMzFb4ZEQv2omuyWaF/wcLaEE8FtJi6Fm0thJ6gLyIEn7TcdDzfNd2jAQtKhIYCQ
iKzb/CsWQokzb1QtM8ySsJfafaLQ4SttO1hJ0wPwHXlb0y+VhM3Z4WpqD9pQ3dUo
UmjSwKu1zXxxXAIgDYs0wwwbZHqR8OoNEZ0xAB7pbahBF4jmOGEirIcWSb9CLz1U
+TOI/kAvZqH/l3xH3/ReeGs5t0nRnzrsB7GQkE1CIsb7918tHSvvnSC1EzC87czC
DmtUPceFJqFW52t+d+e8ysDtEdHLXRLYNqAH8KCufAHweys5kLX4gFfgl+mA27d0
i1YcVWuh4ZiT4I9KSg72IVcqU6x9uk4ujV7TAWkg8i+MMYtvvfs/wYnkSblIOtge
teB7SwH3Zdbcks8EWde7jebWklX+OJWdet0vd6a6K/gmkwa1mdw1aPcG9fvE6JRQ
elUdFDS4wtEt7keb0aQBCUmTk9OIl6rZYOGckg+qzleqH/MtVpbM7qd4akX/7L2R
1SDdVu6Ol8VAmtYK1mkAzvtSwtRqzefmJmxChQSRt53vzpHGB8/a6XhJccclKzOS
U4/2tzCZQb0I/Zr6Yh8RN6dnhzvF5AxjZ0ZVzCLSgcY54BNeCbKZdSM5uiZFY4DW
dx+6+yoUWW/cVrCn7uPtC7v6zsdOGIa8Ew1T79u0nqW4/kcukhYdUzx1RbsAy/hg
NQH3AXVqa5zefZ/6vZq4pwA/i5GxyxQBGezDyEeyOAjH/w4XD/fQiu5d7wlz6uK3
y8wZHfVeYg3YXr6mpAq4ZSYMVwZM3fBy0bl4oXvs9S6FMl1eEZ06iweWN+cCBvF5
WVpFDBkr9kD7QfjSorYBsGlJYXMGNFvXs1mO3bZZtEta9O7fvoNNhznODcTDed9R
Qqhb7pDtEo6jHB/T2UtWoPd7mBxYCwaD7QqAdHHh0VpeF6GXnC7BZcmSy0Ye6cV5
oFjM5bhA0jfX5cUnPeCeiyenFAi8VettCi2rgymHYcQzOTMbeJ2tjgusVI1QUnf8
ofaJmcMCzf25xBvGIpkHppjqJ7xTMQkhG9vw/c9JNGi4cI97BXsJYudcRSOxaYwA
deG3vY0fb4yxWGNZ9s5eBT5krJVdKqB8pTKq3AtCUv4wKYoZDh6fzn30KAjU1oTP
+OjXc+7wSW9s75FCv7LKFwVU/oyKVXM3vAWltsyXJS/+rWrybDl2/J/JcO9UvYXB
LZA9pyga0G6HUVtoXP0EK1Dp5Xk09J0H1d8USosBOVM/YzA+id2xgTvZFLzFaItA
LFWmgnqq5IT7Py3/yZFM58t2tgKonPwJfUHEw/SMQPFI/JZI4ykdO3VMfRKxJiSI
b3o11TWIJ54jY57E8TWkfp8T5gkrSq9MZUcVZinIGfyLVhMcleoKqFyoC2SNlAq4
U7jSrvU0zrB6RRGoExjQdbIauZL26wOm0/yQT7XfyStz2hRUZVj6awKy+IwzGFSv
wOAlU3vMA9Wd98MDuJ3dw+Dm2CBuwJMlzCBqTZNMVgsuHguBp1fohfVY+6ezCcMV
5ikFtjVUIf+TDyPU3Vxv2bdR/cpVqzbzW/gSYwPfDH+fVs71ZHMCh+fc/HMYkl4J
6YziU/G3BIOhGL+IshSNJWCkvpUHCR5zKOrAPGMmTL5hHTD/4tj+hHNeXB1xn750
w3V2GgiyTEdFJWNRdyIJWW7JewkWQCH6UfpzX0YllrQewtUHsyfF1nUzo3ITQvSt
a/mt5OAPp9PXztkJAiyr1/iYJP+pVdt1jLW86PWVAkWuAMzrsWhKXYnOIL0Inx/8
W21jZEXY7t8vDhclu+j44QKGCVW7HjRwiL1YdESAru7HVOq3jXYsUclryszGIQng
7Jbn0gSLc3svK1Ay1Z0+FuJJnQitxZu2ntEQH2CvDZNCA/apDOdjm930GYf9O/Xk
vvEyiT8dea4sqIUn5N1WJsTmnDnW6z4zR8laJymZCOsOVw7dTXe2Yp0fnknWIyv0
yrP4/KWzUrl4PAD4s9HKCnsmJ0vcZGWzfv+riGL/AP3xhU/vmXkwJTHw4jagbMOw
UsKAof0YX1In8RE4NE+ac3zhieFeUS96aApWyw7J70RcdCSPfhbNy87n4iUBEJiY
UkSJAymnEEs55Os/neYRNZBS4q85pXpA4QtGJ1sCrHQEfoOt9rH0qYeOEp0QyLr3
iSQFvxCD5f54RzNSzUsGK7EYTLsimW/5LsSEH6Ng2xWj0xd7SGyqGlZcK8FzBcWc
nfCNuEJZlI6OEtQalq1OjQkCzgItKI7Ls1PvBF+FV49HIUw8TybMcfjeg5UCS0/9
gvTRQz8dUX/IraNnJKnkr4X/U/m5gOe0B7PDOaseQr3VptughlN7WBT3RXIVNGqW
6QuRbMhiCbGHg41EL0diI+iFVYPOnZg4tdC7CLVy/9LtQnuI1CXOwM4pklzPP1BG
RRmByh291ZW3rCuDdApfmyfSfkkidbUIcFPFuAvGOwYqfqZmIqeiA7SaGQc7Kpf3
qgyeOfcu3KIKb6TEdb99aK9CqT0IY2SDPM0BRYNL6mQlDPJMooICSmO7/3MnqxLN
xeNpO9C7JZREiWHBq1Olt068Qo/G6vauJQ75ACwRJjLK8Fff4WqinWmX/JWpF0aK
wuqVxN/bDnE7+eo8G+t15KXtTW2viglEqHOt5S0hhM5ipIjZUCcHRn6cyhl/UQgh
iWpQN23zWosia9nU/kemSuZC9E9vrP+/101lnbPwGsvmKbJ9bZGVl+4+RZclc6B0
2xkPRa/vzppLdDlP2A62/8quWLLRl+pSmXb85giRcLjxmsdczlsYmIuIJPLtK98B
AGPrwrcM8PxLk7NjFQHJeS0qTSqmi4FzLjPlh6JRRYV85JUprMK0l3BgbeTD4DeM
sacvAP8tcRRC5uKTZlK52fUm4RUaiPkvRwhZoHxOn5lKPZCiI+D28RhUtz2UHfn7
Jie4htDiYF8RCozcZqNt8sgym1kK4AU/PXPl3fP0kayL/RPT6oosrgtUOhL2YXvt
OGG0H1tTLZnkUATElTxrrJwCvEW6XsFiOtlU8rkCtrwpdf6L79MTzJXYrKG1UOiI
LIdBTtv7HSFpVBlAUnsW4hjQmK6GKl1dg42+HkPKNda6AyXa0Uip5qWGiwFPwXl0
1zJ4AnljqyhU4neWLpeSpKShdqRxdkX5/PrF+dYpKxUdME4HqU2dmaSSyKjLwuyE
6GA9rhGgAqm4IA8O4/l35Q4zdSzEWRDXFNssJuHSo2R0sg59H2+fvzdx63luZmwm
EdLMWEjA47DR2b0NGekSzIFlgLUOGj+TTfthjaK4QBerzStoWVDqfi8J8Um9xeal
pV7bQDneiCRv5bJZnS7PS9GBmY0jBeXqDf2tZmLNzGf5SbKTvDhOLrla/PEdROyc
IXkn2uromSyWLFxkt7SIINfpytyS8BdqEfIrsXSI76rcuMlXbPbDx2lrcHBgubLE
v6kALE9MEh+xKyEmq3Rw2xYWl+iheQ/7dbM4o4oeo8rT0l7f5dackbpSgvxJuH7z
IwTUk1hI80KuqWrH+oT7w1KBzkePSw9+BrR7axISecRmzPs1HFPwE/7ykYBzF8d6
BpLDoyVJGblerpwdBZ+SKKMj3NJW/aeilDDLneUCowvabFm9ig6nWt2Zh8IRH91Y
khSDwxoomFx2sDrHOJfrhQmqbLTa9F8e1s/DuK2Mt6RjxgemI9ckqcrq0nv3aq8K
Wu8dd8+dgw3G6ChxcF1O8ihF/8R1CHJzPT+AUzd1pdL21EFucepyRwNobt7xgnPF
bFXclkmTatqWaafMGZ7gQI02y5J7tzkXtgPALU1O/kM3rEzLgpV7UR/e44nyl6FX
qIrrr02Bwodi5KA02BSc0EfBabxRQAIOACLPacwUL1YhJm0jbS7h0LVfBh0v7dh3
Da5y9F/DNxzRaG8Vz5iu7f3rs+Fef5lHCTb3YEUlnvTZ4LFp1DIeFAxXeAxzyUJU
s8GEuKYOJt8/p53j55AhA4bHXh0TEI/8dXxQEk4VhWpH0cZJNKgdMQuOJes6njLI
6NtBotFNunUlG60di8Z3GsrTOLhCbDhto4txpfKXIxquEg+n4uqD2gPoRnlCfyvU
jq1sT+k+ZQw8yg2idalmp9TTYdKcQQeSneGGs1vudd2bdJ/ScV6EFOBsLAQNhzaY
zC5SK0LH8y5MwbrJdvETTBGkTuUqLkVQdmil6hdsHzCdvB0gmKYHuoUi2uuewMma
Wns+rvby8VpRCP/z8/0q6tdsnRAtOuphkvKdQVdMlGAc1Mj7DW8GI0BVKcLtS/2W
+pIfMsNuAPtLoM3Wrv1msBhR5+/QdVkza6kBmlmZ430++22LUKESs1IEdbopEfUa
nkCRVaIOoQdO63kScNIc1fdnXk2zEjzOtNMYBTxhqCobIeXjNWGq75RWnMZXDHDp
e0OQC5cbxqd6IxYDzJsTmNRF6Mv486zm55C8ipifeHOs+L1rZI0Kns8gg4Eh83yi
BloV9fUH2gGomLgR0FcxuxYsuQlHzXxei2P/3G8JeLs1e3I3+6HDuwPwKsox62CL
AWYks3765qM23D8nH3H55zpFMJIvHPPbBrcnkhrYDjV5CTidsyYNNJhTEnUuICs+
tm4S7gyr+LR1mM2JdoTRi5QGunz+CKTxxPHd11ISi+YKWUtCZTKu0gZgkIK5Z5tY
ht0VDIh1DESqh7v5SDr43+oDP43Z/SqAtQjck7qQIXG+fQ2i4/zigo2O8wAL5bvL
Ol+fhMeyrCa+4kuZVp7oeq19FVM3S7jFw5Old0hsmhQVqOmOwZs5eoVeF7dD5rzi
47Zi2/eLk4vM2CHy1NYifff2e+k4+ZNd9j3iTmt6WGhxDJb1E252Wc971BeU44Yd
TLSNpTb64js9XMexcJsQA+sA2aFALVl0samcDPmOH0VLEId3v3SBHjnY2pmwtOY+
wZU2BiE74JtLwe54VGuzWhZfKBZ5t97eYNpy8wcpt5OFPu4XgCarkSpomtPWTHt+
l95UPo+hzpRkD5jOxDqjS74+MUyunfBIx9LPVws5Ti614vsOBJuiGoXMneVDvUbG
5L5+phGpbpFpmFBe1PMrozRwPB5qPQl6cFbDgJyxl4yZFiYkOpfT8aTfW0n+bhaC
CZ//rFUUxdaUGNOuJWWXEe9GDrvaJdI6UgCf43gV3COQxoe7MOhul5U84iHeRrZg
tEWIk+V/KPA+kvNyXN/YZyitBNNJ/gtzKNERYzFzFWfUH3QFRmAfLp/D8CjhgBTX
F1/fKXpkSQZkmbcgVAoq4OoSWmDG+nXHrbmR+DSPDnTA/8LdVinViBSMLEHlHR3H
wKDFa4rtoh3GydNyQsCkk2bDLUQaEnlPk/9qKigvUNvVLYfzwiUnrQ8C2Q5bxkIm
VQioLr1lxrjhLklM4rpVeUKihonUUiIx7LATV8DrweRJuYUueAg3CLArXLAuCfLD
GB3t7Fom5U/b0YjJzAVsIdIjhTC0yICfo+EMLIDRBuNmMbu65BnPbfFIUxtywFpg
pmJCE8enKjZ5wa5wU0lojuoVmnemyhlctGKejTstsaSe3e59rVd9+iPqJkYOesGi
R5X6n0hFXlk8oM45cxUkJ2JDFhlrrMdNmwu2HN8hoqyTrHm2vljLgTGivVH1l4zH
wKLjF9E2gDrkwwuWYxYsB46BUt0J63qRjuybE7HBEa0+/X1AGbFGM6XnkLe71k4d
Ed2ztRJxrxvwICvE35aYz/boM7ZICsqROoTjQDJjyqd7Yv9FZjd+w6GkwAQgJKRI
YGknzh0trdSMBjRnW2AGYWhiywUymlmfCyJSuj4uJVZp8wGbxdcUm+d7zyvfV/RB
8oOr1Z6QqwCebXjhKcH03IBMllZnoQapOCO2TqV57snMC5RopDBtKYoZF8ckIFl/
+L6Cu8Pmy0wT3siVwSkerLHh9HIzzqJ1BSzO/YjFK2S+F4qNF3roVUyE1JEFF9u9
Ly5h82672nXVWQOMK+cldczs4MBy+6p/wivqcFEKvIY9oYgE3l9lGhZYEtk/LTg2
km1pZwoHjYKX5GCYD6JAEV0EQ+y+elXEFQbuN8xicGoTjavHgNoICb9C9hFGktUR
AZCobIk45hgCAVzZhweFFZXxh8jeV55nVzPtIT1cdq0rKovfx8Xpxzd5QPoEFG+G
JIuDxuXTQK+9+LCtCboDMV6hiW0/Q3rRJXPswTGyu9ydKR4wioiYuuxpSlXvn6sJ
D9D71JDXmrVbKsLBwnaSPjaGvXtbvuTRvpE/7UoQYSAcl2uKGQqLYibrPhNy99Oh
3iZ8yJTxKd8CmMVsJ7U5CznZgjoqihlq6OFgVnbnqB/Kz0RlKx0cEk0NIU2W9BYX
10xayjNgrOOXCtct6B1mDGfot2b9hZPJtnr6Fu0QxWrsepvaMuhmTtighS31m5Cb
MzW79MQZ1V6/1dZDomGFHpKTp63EO8TBYTvXKUVUt5LVliumdGzmo6Ke3UoFG/Hv
izNwxq+4pgYebM0V8gL0ELNEVzrDhIDLh/49MS6FA5qO9DUfI1vRsjsifWbSZDoh
gOVNa1o1ESnh9fYhaDaWnkE/zGP4SU7ogenBidttqA3/tGwKWuFD4oIVx3x1qs1z
1j/yzh22LsxYznNWdUbc9SjHnV/bqErSCZS+Eduo7IH1iNrHXDgBEZZGYMr/hqlz
btHZcIASixKvK1XBldcOnswXmn+jcAqFwLjpzhymYdvi5gsqiO6uvOxx7PlfmLYU
FoyMu3VHYvC2SWV6l0kFgiHLB4kiSWqV0PEvI759vrjJikvjgk+UekRJKIE06Vp+
4T3wgnc7PgqKyojhq08fVAgP+zQLUqWsTGKUQ+TOczLExXzdR9/ClxWyc3htKGGO
badxqCwyOtbnT42I+iNpGs5bd5fpLQVLIw3eet4i8HKS2H+v6bTXwY60TDoErBf4
dzi9CPRvBY+upV3NEBLR2ufXD7WRwNRiqhuYOJbrFhQZ6Wbqu6UW/nDndgsMr9Ts
yyWdEwxvingHGmzj5Uye4rgohOYhS8wIRALFP4BvUmu/TMuNyAmnaXZmy/AvKQfD
t4hzqnnK++UtXlmf36wGr9FmYnUnoUSm680ak9F+J9O80FXJMhFLldJlTW850dhb
LJGSA4vB5GJ5OuZ0ws4H9hswQwQL0JY8ojLaMZuGM6Of3z5BtEX/H21FN+BSevVU
3/xQvSsiKDTayATlcu04PJVgvo+EQzSP9ZWypDRgCro/x6+d7ONxDanOtfD0Vnw9
6F0wX0y4MwtFQ1GuXjgYnBMZvDJgN9pKYqPBUOpoSmyB4b4HxnRIOPAiAMceeVG5
vhFsyIOYOq4bOs2LSted7/7aCqKLs10Zz9KX23fNtD9/pziCf5AFLN0l27hxNJch
svoGBdNUAd1sBN3tU6ClBhLnl7+t6MpLkNdJdzIK/uYLntkz7Cjc+ko1DE/duQE3
ObTgQjpgrJ9iqNJ2MmiHUoQUqE6Uti83FThlokIjo1GNRFjyAblmelyzkTCKC7EH
kTI3eQDCUO2p38PTIHc+5A9SQQq3/rU1ZxtzsFrXc3z5ARs6SgmcFNTVlL8dFEc4
qk9TaCDGz9k09+9FYKfvlnUC3K+XEqD6gdsjXMSOEDGdVXPdJvhe5X9d+28C3a+R
4qkP/WZkQlDAoLejj5faTZsMfAkHenvAHyPWn++VzMf6CbqHfqkmFtJ3+IXPkb6l
K3tLvpQ0cK4OL4AKSowIj6/0pYfRWACC3FpWFQMx7FqQ1C43wGA8n/fqYhD+h8Cf
KXFEy3A2sKeWaHgU/8Tq00SMyf0fkrtXMsAGXten27etS/iCb1SC8zbj3zQvkMVW
k6U9A8RDrzmBlfeZl7TlBhckFDVxf2Js687O4m3yAUrffVa4y7UWv1PFuMM55bmK
nY4AdxTGtagPViOR/DYqD6WRXCQXHH/nmku7/LrU7oaCPw3UlfkBbYCH5/4q+B/D
WegV4NmRbbmUeRCT07zhSZUX1c/GUZvo21zpt66517Qmcf1j6pwREaD7rViXDRiJ
ZhP9vBHtxBQjvVGeYgjNsb8dYGKGHo8SbmfV3qN91xY7uvXjik1WWkxXrfb0LjMs
XavNb2SZNRMxxVaL7YaNQmz4Rd7AzbkiLZbb1zaOE0v4YibzugzXKB8xaKaXXoCU
3iCNv+lpZ5PAscPQqVYKKjJ/iowXAi24jEVz7JAI3g/pVwZZ6rz0B7aOXTmrohgW
zlFBfTinb60uakrQZSVeMyEoCnry1axHQqyDcxLeHS7oVPaGyM8LVv8Fx2RpyPxV
yDRqsbZjgLL6hWqXrtwn3NTWcBlEpEtcRdFTXErx9MHIcjhx/6z9kZ+1UKZNy3i4
nl0s2joBagNQhJ+hZuH6UvD8uv5Cf0eaAEBKAtgtwfF3irfXg9vyPDQ6sr1unrV3
GTSBRGdGIIXVWxqlwOQ33zpwypBPF2bi20O1W2DUuv/xHAcuKx/s6MzxI8x0cjm6
QtFZkXiZCH5prBE/VqeC9alAtc76+yPMXSJl5Ad8IDraEoorX9z7t4IbUuFlkMzW
Kyz/EDBE+8cyhHRX57eAbNV8lMWiedtCwU9XQ5jASxQWb5z0LFbQTDm6RFSq6Dwk
fHkMxyniHVucDU3bG6aJ0Jm81ZHxu4rPgm7NijwTsQXWw78ZPDQxpGHssdhzZfU6
SoTBWrd9ZoWtBgFdJkoYj01BC6UWLw5K+oadjB5HQVYx4hxoMX6wH3MV13DAmUy9
MhkvZffPEkM7orM7OCRQU4YbpyHr2O+gSSzTCuwVKbTKf1wWTPeqTIBsx4TtpW58
1/6/3tN3hgyDm/CPUfJQC2u3ndAl7K+6Cx/IfmtJqtbaD0lqsTsIXA7tkISGWDhp
GAigrdveiu5fibTykK0RY/i9d8KvdGPycnnzwzGFZ232i2/SkwdihUe7ESZ6t0Ng
mym34dciIk8pt8vO1U9KJ+DVSh4gj/TdcxLh0wkEMJR3WYi42cmxJ1xjCuSv1vZ7
OCIo/j+mXBy0keV5zanjVZyuXcM9gwMws/IN71XE4hb698pAuZm4Q0E/Er4AgT+1
yt5jaf3drj7CFBz+0QZHL1aTUyqE63Y4BGnAOWhESMDTbHR93XTf5L7GgkqaUuVo
V81A0JmIGz0gPyzSl8GCQgU33nAYuYhcXJ3+2he1nuIvNwaYojcbFB/K2Sy5Xxgt
kBeyXhOa4YtmPXU8CqaBswSmb1lAFCBveAozjQ+TjeJvYY7HUaFp3ld+ZueXy9bI
08nY6C7i1gMhKAVBzDY230WeL+/BJKNrykm1270oF9IEjQdgPeosQ3yxBFFEunq6
pqMGbf02mRim3AwNmyLa4LGk/woEhTvzDph5++BtmhRUFPufWmXd6ECPCAxuzrVn
QpsbyuS2HtD9u3/cAZQl88Q28SfR+IIlH3hX3/FyjkF+oa4bGQS1fBaoDhgCYHYr
W8LYUnnuowS0nhipEzGU2cCqkWqGm5RCi2aVkPudUuAh89n5/tRqDlxwdVj9tcmd
oR2SPTcgXTtVoa46IKFK7aiU8I23+VwlkZxaRTa6zdnIvaB8Zw/fS5KlHpyjUcbB
PUYVt7SMc9CYr+7KSSm+2Bysy3QamiKUHQkCVjH0ixOSDGzrKdes2OXD6t1ylNbK
cW6WB9tUmd2m6AP8JkIqplQ9mMSM/TlV9Y5422VjeiGQ+L0k4syD56otqKmr7OiU
ZiJR7yJWIIzx9V47GASif7V0bEd+ILBFomTOBhV03+4Eg5qEmp4eg0yBkPtIhVee
lRNIrUzyKZTiLUem8E3Evca9uz3bJQ+PqCXwMseUKtjWflO4BBCGT5pINdNO/IRc
9qpJvayMcf5MT0gsZt4LH3p+6WseKnci996b26I4TYx8FXaEZZSgC6o96wYqVS2r
zSV0euhNPFIpksfEhrdKxQsHqB2mzfRZg47kl4hXSjNJoxlqAt1g0y/krOvbmsGS
0nbOvFKMK5qxwIXxl5rZ7Xb5NgPrgrMcKtdN3TexgmAscGksldK8qNyoLy6bZ8Nb
r74cUwOVmYjo3ZY9fCvR1RuMN2nE4+oo6Lv7bBWmZjnzNBiB9d+bTDL4vUPLxN3+
voDdEmvmWTahvx/CYgL0dlThjj73lvEYtoH9FfSiokkQ5sVQ/Xw9J8bQsXhBVEvz
iqnvi/qrA8+Nzu2XgZrfR5nh6w8ab2dh+uMwvOCg7vhp3zxQDekS3RlvAiR/VJeU
zBrAEO4AwwLbqZ1kRXvt6R6qn+ssbLyioejqwqpu3awZdEYy8G2FN6l1GJ2XPMOu
7L89wKuUKqVtEk0/SoeVAIoXSDkPsGpdm/GDw+yuX1Y/iPb96UbSTiFVuno1QOxj
8mKNU1dTw2ZZMF+nAophmHs1n+/SDh67RrZjGOkHMNA7Z8rlKBB9rqgvvT0EvQXs
R2pgbmt/R/s4xjE/UsYY+J6SlEitvrnw0gGqiYUsdhVsrTZuDE2f+nT84kcT6D4l
KloGsBBrtYuQXhPtut2aVPNwPzRwfJwoiQ8AbDCoun01qpalJqRAnOI0GxFG48ol
MV8Uf0rw6kUGhSNGQ8xeb9Sa8O2RknxRn069R4m/WynmvYg8/zNCCzmFype1A+Rz
7SI43brQubx9jSFmzfOZIl8ATYU7eLbUEXD0YWcABxc0SL4M4kwHoDazUE8iFfP5
o5DwxlyOiunmrPL0KnGBHom5iyPNdI7vHG4J6BJaa4gg0wDJASsBEBq2B9V1RWp6
5gnzZ5DufQ+6I54sdr91VG4TxH9605HJ8e/AVQVILrt8KJatcjMflhCpdc84ZaXA
aGsGGBwfN9JUg2qLmgG0pj+1crQOQtNp9BmqYRuS+7fIHLnvmvF4XVNJJbAhA30h
BZ8kuV6spxgI3WlKP3j5+oy+mp6+sYZVkK3WZo3Y4ndT9phKF6VtKoNKW2lvYCIV
NqrVeyGg/3OZB9QfzAoPHov1+w02trOcLl2TrsG5fbCLNJ5StFYbm8HQvCXn0zUZ
OeFaPT0w5473RC150SqaRlyA+zxsvueps4itGxkxzMkowWRO2xhHZSKFcE2Yy3hq
ulWs2yyYU2rGhVIUISrb/UtXnPM0VbG6jklng+NOtroMccn/dDLtMetTLoRdEH9v
hH/zYwNfqNkYKDaDr0T8Z9FnR7fp+uNB3dzR01aIcpIQ5DboKFfa/vZ01eYYN56b
nFOSoqPAwnY5++MGflHcGlG2Rd8nuzsxNXsdvvB6WBI7ZEG8jO5TTPgzPF3TBRD/
lcbAW6dNSU2DI0zUE30KqjbCBoebeKB6LzZXMLE+wvExGr2RNWGVnYa9UBTErQyg
4y7Im8wxEoZ0UoUC3E9K5v8jSoSYyYiXadSQmAp16t3XjxGrRYt7cISpD4FJOHVR
UKzWiyJYhn4bKD7/L7bt3yTL2r1gzMVNr0G7M35PszHjYt3zlvdDH/nWkSlitKXM
Tilve/ULAFnVYM0g687zN1loKspST2s2hJluWB1knGVoU5SuVuxdDOtFbKs9KSmM
Q7SExpFJY90yNaKzvpJC2G4dWaJqt5+lK7JkBiHHkxzfcOkWZpx9uLKsOWzmtYJm
VYNkkJmXgJtyoIDEz6T3zf5gC5xGOuBA8uDEgA/uKOzouOltMo8uTnEWrEuKC2/B
BS4Z/oWES97f9H9CSAcXQNDvd4Q0oVZwxSc3wmegd2J3ipLu0haZCPJP0ISZQ6yf
t3np5BnsMw1RRSZ0cxtkKgK2VyVMi4CFKjXl3gpV3wj87ajSVqRrWNKZDmiRtQmA
2ZuhPv9VmqGo99eVM4tiXDJLjzuvyZlQHi7qEgZEEm+Mgwk6E7FfoxgL3S1My4bx
yLyiZR6kCRd48Ds+asmf4BR5NytRDr8ETyZgJ1J0ThI0QzWYfzlJK11eUI6JnRtH
7YptjhJFGfrLtHfC7ReIK/haOXTLJBBMwsA+bGnTzRJh6Rfe5vn4UD8vY+hCYImy
WFg9nJ/pS9Ar+IFPZ2G/O33R3oApVzn+7obT2OcS5sceW8n8OcZgxUHxY5c2ciyR
KmcWpcVFHpm4+nDiSQDb0shJDmlufN1yQ7VwVdniGt8/rSUnTZs46sWMrQhv1gt7
rAufEx+NYMr3dhKc4ca8QJkxyzLaVKD84iZOkYX4/FbL5f1cONq5ekOR4hG3EUKo
wyIzwxILN62fqe+OzVZxNoBe/gHeS6aaTQiwXxcN3AyouXAq7nOVI5DJ79fKzUJV
k3PHFoEb8pFTWId0lTV+a+i27SHaH0Vwxps3DLAPir3mtNE8sVyXld53R/Ipq2bu
xSLrAo9fG3RodDvQ605LyyT1z8DlF9EHkeT++qTdAIARfFhUW/gfJt5MXbrDa/Ku
fMKuU70FYxzIl77IDSoLJ1g+scq7wZ88He0h5gs/7ZWyCYqckUY5lVX0tNhduCtc
uC/XHYaAGhqBpJMk+1nbhoiYbYB3toWkeMxvSLZ1zr91qLJmD8VQreSFchy5BqYf
/JnpOhaobcd0kUO2vQxMbgzkK6muGHLQtUIZ3qAaudCSAu2WoZilf9f5/IxLUSzU
qjj7pn5QBzAeXl30eUNq/ciuhqPZ+d7gk0B6cUWaRAKldKQKRTQXPNYOjEa0L5Lz
toa5+PYaWdREozlRbx2IubZlZz5e2J9uCVYbNdHkbAcb0ij+qvUPr1nXhkVl4fNU
9NfSL/gzq1+bxHK6rm4OWm8r5f/ZDvfE78tHuBcClqXyfXD1ZasF7EyKiyc6bxet
YhyHnnif46nkW+T2KF+rVr5l8oqgPu+AxzDL0RtxsxMUf4ar1qN95GO/Dg8N9jKA
FTcjmWomCa6BN4tFv101H+JH8NE3Xr99VAPuFCmQq9tbWXaCNuASSlQjC1g/GWS5
btG3CmLsh8DTP635VtKkHyvlmn7mymzG8sUfRBxJPOiLaoe+tMPdDYvUQ2DPamWQ
T3aEmNbQnx8OTnJVGn0eEDfLVE7lQU2fvkvnOHcF1KH+EXf9MtIkcVkI6dgE0sBM
5CAUfxSOf03gkfVGa3T0Ky1R7o3SRVQCR8FY8m4IPg1OPchojnbzZuHVlYtAtDr9
mALaoNA9RoLJq2CxkODiUchUc5WAZcnLYtq8uGy+E5reIUw5P03R14ZPJu5mwFQT
J8PjJSQLPk0fJeLp2lrOZX9nafbn+PCQwv0aLU7hFAGep1ZnhwYGsM+886gMYueR
ZdJzuu7yYE2W7LZ7Frssch7XGASBmJIZdvFn1k4npABieIFi/sRE906a4FM0ix/J
8HSPiV46143vWsGAPUaIPHRSyvPI5/Un4eJ626JDMtioMLc1UWxLXvhQmti6nkno
cgCCXVF0y5Zd/dFDMlE7nvVBtiHPttg08TPoqFrdy/QSk5+Y34U3rW86kfe4l/t8
WfJ4yIKovi7cp7dPyXssusDzSu7FC1MUBocNMuj9xnBu6dCkk+HPyzDsbHFHQ9vk
r2pD7PpSlLwzWEZIIp99rJ3DG/Qp0B37ZchcJJMxVYhdrtCGtJBurLPz04XbAPjM
KZn1ymeBQnP6n6WLFdvfykUTTWlbETyn79jYplQ4AtXiUDQjUMqgYe04h24pWGqR
OtYZC35qV50p5Se/mezfZ/2JdxGsMbdrAg55z61ArQCYOI559BS55VNnj9SBfEHf
UhB8SrdMZDOHvZ8YNAsXL2FhJ3r6VfUF+YYKunPZK7VpJNt4u0PMpd40kejjR2do
JSzggL1QQRZFR9p0hThX8pwQsOIHN66VZhYN9mhL7wfFruwzA/oisFxkGRA9zRpv
tGicjNDxhH40Cvh1J230zLG03Gh7GiiHR9+sojqVchNHkV71VPtw04O+EFJg1ZRr
l++rSXZdsm9oog0Tx3bBSl1OkK3Fe6H+K1+9pSn2q28CrUPD4lpscVabDs9ZruAt
RK+b2IdQJ5SX3ibRRmSiUxlQt/uFxePDcRCf/G7GLZNahX1yDhODJGLtSnfaeyAk
EeD2gjc0oTr6RHnpOKEknZpOhFz5iKqDVrhCUg3rzn/ZBp+SQhE4DcHDe/oKny3M
H2upxd51qhyE+rxNfgGJEwEVp2DQABxTfKfwdrcfFjjuehrdbw8ZYR4s22NQ/omw
7ZGPX5BdnIxDKIeH+cyLhEc62xRFLkIoUFQ7iocpXL/FGVfR1OHCXkAfKKNIcz67
s/SueBcafNk13vzZ056bNSEfeQa6V9/G8YBDkhcEhxk8YTRew/P7RA47PVUmKtSL
RarB1I2f5XSHMSyhOJNBckZ/Wjm9y3vMcvi05arfp+E1TXO63GyjssWTUifuZCOT
Tl7uxpV/MWbjpL0Y5uaE5ZMlDQ3g5tkksDb7as7DJfHZN+GcYcBtRj/ORbdmgZ09
7BGL8XOv0dchP9cIFwqNiVC5dEZRl8fF6Cu/HZxr4wag9yGaKTL0mcqWVgyWdm6I
ubMiAtu7ZCIF4eOka4PTh2jLa5MLOA6n9yAZ+kGOduAKh1zkrwmulk8MoZwRCT1N
M1tk5YBqAURsiIL9Qw6ahO1a14ghm5lEBzACjpnEe0Uubj4+JT+e+0vSWLtkOaiN
FJZuJRaXUfUkz0cvtdNaC2j6EVgkLhOXlHZn3PmYBaUhQ2nT7EMvPkixUZzJNAMd
m3kztG1WRdxxhPHKkh2cAjU3RFkv0LLwFENvbs8GIe7w0v5T6mrTZQMSd3cRbVBR
8O/C5xFNXWOGU09g1TxI6mOkeWX4hlyijf0X8hIFZoF00fsl4vXewOcb9j38eW9Z
u4bZJsvmnlujtoB2e3qyLtpGid3neXKsfhQOMZUE8mR8pic47Af8geOjI0Ntws+X
Tg/Bcz7jv6fFs2H5kftcqauHD9vrq7b7uIvHJtNHXScxLkc4sqTc5jc7HDSm7Uex
yHpLlkaR4W9lTrN0p+k/oRfRYBkXx/GOzsvT0QoOIIImczCEYBRauJ2Ln6D/RZxz
coQIIEO5avIENaavId7DxPENiMheyv4LRGLkCukpMUwFhPnWrsUGj4s1SzpAPxFL
o0H1WjVmffy4aRqFhMN50grzGGAeYCCoBPulU7zVZaCS4gAKrwbXaHztH1y+WJ0P
1baSSz6BrsEKGpydXgYWn7ZUqky63PfUPFkgxC+wwz75uWcCZ5Z3h80jdDUZ+L4H
hWrZb2v/Lq5TZ0GuFD8XVFPEFYrviv6NWlldf2nsKw3DJ+5FrBucrPcPXxb3n6hh
Zj8crNL5NBzShmmSPUCTCtGlNxV0ccPX6XfK5BUB1egwIweFEiKEUKcfNQNQxcAc
d5Y9a+877lEziwzNNdEGCDLkW+WeAXUW/38PJsnhluItUzfeyAs/I7mB8uz1qdxP
NNzpWPzlEz0nY4rhdLj9udcvw9ISAhARCtZSuwf7+K+MMO78AhsPofWQwFmSaAJb
GUtIlBoW9Qd5Hctl5p8u6hXjmUdm/5VeE1RfzGcoB2tUW3MI7cYtto0Q0xhrVOJq
mQr7oQ7QKfDympx0XNA8EZqgFv01nvJmZy8R0Buh21kgOt8HtZdksqlIZNPZlCtu
FuF/BHvUY/4vBBxvbl7KpUrnOl1nso5l2+/GK+AcxEjT1DmTOn4O8u+Uo4LD8k33
ummYYF5v4nbZL8+d2zy/5XB6wMBlgTdK+gFQljr/tcnd4HkZyPyOkdulWYIoMb/m
EXUDqU4wafD5U6EmzIvJmd+4/hmpPodS+MD0nvXopL0mMI+d9gXFycCCiFbjN5/C
UVTAFqThqGTw86gqJ9XEQShabZbmO7Zje8f2kkhUTXpGlCSrWSmTFxOroi+IXfFy
5FUgi3u3v6QQWUvj/xbhpkhMHF5J/IHhSUafFMpz2ZpvrBDZEzI2mbxiilcOOChh
eap2Nh2KQpJu/t+KDv6mMVAosKkBJ3DOwYE1dOPuhsnWAhxs/oQQTi+fbWrHt43c
WOr1AUy8Gtkz91YmsC1kEtKsFMYEt323hfmIElHrBHFdL/GYw9FKKA6Wq6R/dBgR
1Oeiznx3+34Qn7aa6W8ksnml5xEpcXlvQVskMB83dMC9cSe2xgufXUpG+gWCKFN8
kybDaBuhdQCk5VUjHg/QHGdrrHBtr/RCcdeqIYmS7Iv9cZJnOW5fgWzWRR2e532T
9RicHor/QmRZ61kQpm+lF7GrYIHAUU8E1Uo9XGvWW+HUHGiVFn3YBfGTwFHCijVu
QdOOM69QgQeZddKIIzvjwiCYCXe/4j7aqwIRDpsxKlJ5eY67xm4BsPU8Sw8ihyz6
ua+I1iZr+9eEgHXOM5I+9mY1QJAbhCbSadacTY8vfmpfc98Jchw9wiPkJYDHW8kE
mQorUofURfMJHxEp+aItzIDg73CCGtyIQ/2vkS6Pe1RvKDSUCVVWwA7MzjDR64cd
SnC1borw0A8wSHHULm2caB9GyTfdL3L7hOQhDgtTwogaiuqp1y8/ynNNT/8MeWZB
9Fs3Wt4ImaIRqSttTFYyQwYQZMzZjWqNqHGF4nEdemc98DJ+v6RM3eRsLY7uEE/e
2uZzA6uX6zFV6WSed+hr73yJAH+2h/+V3KarIGfSJCKrimo9PSrsQ0p/l2L6c1yY
YoJ1igZByjV+7y68joKYccn73VjpG9vnyBmVT1Yi6+IpxyJI8fctPj9XR+IY60X/
Ur+xNBN1Lef85UlSiPQ+xLa2Ugk45SvUuQR6EMRrq2pQAClM1NXoZwtwaJx6GaAk
7VplzbuG6RViPinC552BXHiqpD0enzEbC6n/HpJyBim0LftmhwL8F/ne3HHqmaI+
SblwTZNkQzKCaODQRQ36ThU1dswIlBb90I2VRX+WxgJSMDXEH4MtD2nGb5kQnmaD
0Dq/G/vTz07EPnPqP2IIozhfT0lf4IRk+KOqaD9Qqgf5zl7lol4gNDPGli3i2DUf
1ddXDWM2gPOM8yP8kdaEu9E7SUA+SI91k8ot9plzaz3X5dhc+V1Ig49cYsYaqNou
grKZ0DaavlfCyKoEV2gmTAk9z1KQPJ5qkkrDP/g09RO8Zy+P4nlIUOOUbgf6ZRcW
myMp8GzyCKyLbJVx/yoy5sAfQw+fz3ryN3A87d/f7Yvb8iA+5V+ocI7NU66yPyhd
j05qy6396smDoYQefMxxSmcvI/2C5LmoTZSn5SaeqKTKhVjlPq/dErwlvnzbiiXO
7qCQcHh5aGGWD4xNDtJZjpuCP9GoPd1mmqyl2L+a3hRKff4fKlAt4AxYkxQTQX8P
ZAJQCWj5aClo64B87YVuIXBwScZMgTOrxtKqlL+5AvEzCuP1VH0sJ2CkCWienclq
d8e9iW6htfslk8fzKR3MKrsAw4qQtPkIDFVMv9cBKsdQy0i49J1xHwMjA0U0AZTD
pBtPs6ObHmcJnS9rkQLkKL0mpnOg+VIUj7ogOuz8MBl8aV41uZlCcWiK2hBCC0cA
KCgIBS0QIlYz8bqt9LuVZrOfQCoH/GMozz2ExR+vDuaZCO9wy89WPxJOrzwvAb1p
CkOtY9OE2gHiswnJ8pAkVWDOItnw859K/9QUF4U+wo3upzAg22/6JbO1GHFZWzFy
UdfyyqE3GzHIsnaQHKuQvKlnRqT7SJfD0snsx77KQa3jSnxD2AaRd0wKKnloVOri
9X+M4AyeifztzwBpff4w2DvNOK9fPp16mmWiYQ8Uv02JI6oj3VCgzuh7ztDd2pu6
0kJk/IQg8DduNQvMUyIqtS4aOjgv2f5AyZHcLm+verImx2tjlmzfUsBQkF+VU+HQ
FuT4L0COS1SQ1V0jBDrEnsIxWOtbOPmK7zmeKCag7jCmtC0OKzxKGLtAjKBAOpfj
l84DRCHSwKNH6WT8LfkVRlCy3Yx+xP4tb5lxmA+HQcYlolJkcpKlciJxq/UzQDqN
HYu/dTU6PoU4dDupvKufGFpkUHJmw3MrDSc2cH3J8nYWJE6UpPPbw6jl0bVd1Kiq
XJt1fZ6j0rHAOKNSi7vX375oLvld9wJtLmFzl86SbPtMRf8XyTgNhFAoH6ROI3hP
/rFYKenP/WtfmLmvyFFwxcfbH/2mlYgoZzmKZ04SOOq2wTTk+83k9l4psyh0qh+x
NhELnVReHh3M4JRnlv+54oBSqY6fdA/u5382F7pq8nosE3/1YImm+2Kgoy4PWA8C
6mppgY+W2Ctudtu8cvaX2ykqZN8tu/ycA8JejwrMZVk3HNowK8Sh4Pvg9N7OoHv0
tmS3JqYre7SxF9qr20uwbiRslbhn/L3rbI5ay9SNFg4JGqCv7vZwH2o0XMXVxD1j
Hj2LElrDpFhwijCtQc+HXExe2CgcyGCtcksFMcOAsdmKHd7aMo1tjsrWsWDb8qt0
G5MtwaY2iGjVan7zN3k8Q3vO0ari+sFX5rSQl3sWiFTaXOwuKm8qqHS/wnSFsJXX
2xHhTIiQBVR40iGA1bLoFvwqEFK52tOJTCQfnzi5Yn7beK01OuoFo90iZFJxxS2T
fZLzlAhqsVAYAIfAnD+I77cD0BJVtCHq5OUKHsFHn+U+bWDDCT4crigAz7Pp0a+p
lRqB4Ybpj29+hg6jS1ydsEQ4487PIj8vXLcmW+4bwBcIsK4LdFIWgfiVrfligi6C
ty/8PyK6rNnNPRjQA0v3hDCgIvrcYtNKKvrGNKQ1tlr3qRIz8YxgVvbEBTnEf+E+
vpZsWAI0kqdD3AwCNkmEdhrV0DggNhlvFM9wTkGqKTIx30mm4d55K/1XxGAcJ691
8Oziw2Dlj85pez/Ruo4nFnR+u75E2/ZtMSG00PBcjCuWeHBrPgM+uwUm0dNN+QSC
jJTSZp6ZHTvjpPSYpTPGUj+WDLOYaLZxhQZ32lzcmHeEWH7dWvCcqCvrbVIk1J2U
R3ASqJhgVKq8D6oOrhWsBCBvCsnvrkWZF2NwDEkWpU6e3xVLXhMneTvbmaUTJD2u
3vkgVGLyh4LTAFmmDjybkPe4dwfcXSLjrTxRaHi0S3M5spY1HK8JMt7I/nTz8K5W
6jCsvk+l/4rbbFZocBZOKpbnqm+8TPCw7OnRoR1zkHoXOGnG8QEKrFp7BmoazJfz
Ww7ps/kyTg20kQxKkLbUD/uAMtR2p9pMk6uVzV7DewVHeMWcEIwbN3e9+N5Mjxgt
Vft3N3my9QtuRgmo2A6FVCtBlENNInz/4jFv8QGIx7u6ErTI71SZ0W/USkwMTwrF
ZLhCAooKvfOREKKzEPzxQzvfHbbLLwCmKfjBZYd2i0JGkTrboffFNlM0O47wVwhF
mW/gW3LsOyxIA65j6Vnvhg7l53fNYOh9cQ7zfJnIuu9NL/Ztg3PWDs7CHRfLzMmy
d6L1pdPVImoy6sWxBg2j/SW/iUVY9j+D0qR54LxmJRwNVFJzZvSUnIhQI4zG7lKn
/B4AS6aUmYHwOKjadbaYpKatRNXg4zIk79+ugENAQvT39X24pVX3DtHhe2vI+JvZ
wZvuQC5mjZcWcrc1Rv8YbEkP7FDAX4rwzoW3G6ules85L7mIusL35bUu9gcWSX1p
rIbdKYA4g4vxCakOqrTt1fg9suofCtryAxNNKZXeuWLtlYjrI64YsA5HS+woMMq/
u7TGh/pSIUtsfCoXaxp1nwYikD1o6fwxoUEiQ0fUBOLahx4z7opJTsv2FsplY1RF
Vb8bJjyE3tGCKUjrBbcrF8CBaZdRlAsk8OvQrnR8qhfb+LVPrvGdNi8CkpkqxKM2
2FkVLD+XSTlix00rVerz99CocvrwBfQxBYbgdek6KaUc5cklmm6YRIQmJhbwtzot
ZqMJnWro3SWBohdaY2U2UJMGmej4GTtk0fP8k4nGUBj/bBhoc5J0MhzZRo9aSDkK
7E73bve3BwY58Fceae8jOMRBRCFVjQ2/B8yU+EtEdUsURH2twIL2hsdBtWXD1izd
oCz7i8nQriGHICvb+Qq3gkEtTAY/3JluOXc0kea16KWv/grQJ9az/Nl0EV2cR1zO
mAdfWtJ+xPLhT60Wlxr1pi9xCHZQ2LXha9rek393X3qCQ5kGUDF5nGbVOryb22Gw
hCXSZWGpUhjx+77X2RyxgZoKU70uXYpcb30mHO43/KL5pOH4XZPVCOrN3YJfuXhb
UaQAGPe+VTLuQ1+1GdXjmKEJD6JochNxynJgGWroVh6YRwXqddB30NOs2hBsdJ0g
kTxXwy6pT9cLGbY7WauF/sfvvylzgEW4xWR+V8P60TReVadSmRkiY4UKhXuwqiNK
uN5XINg55JvKH3aQWNkqPV4GiRkJu6ojf4fEV1dQLQgVSxAuAJ/qNvTsvjiTInaN
YCKznXNP00CCJGo2ZrMxMBWBbU2+xObabxUyZJXRncf+ARBK7FpetOywCUi7dJ1c
V8RzD2S/erHPOA0Cs+M5fuMcEAOlwC0EtGKicOuGTU2SJWLnCdFqkV4LwtmXE3bG
hQN1BhZUgeC0dFDNP7f3VcP4p1ZhUicZ+Hf/iXgqseYZO/9iFH1GJs/JtYISfEXl
34+uB5Is1Xj+hI3quaR3PvBviOdRr7B9mIKAq1FiIuV6R/KSb0NEM5SWiyUcPJEC
TieyavxUi14d0w96S55OkuXdack+ZyVw8HmkT2dvVQwhjg8rX5G/hr40CNNcHGMV
BF88RrLde3wX66DlKtV6WNvPZXUUE8JphA7PwkmljZ+bYuDhFcSYjUJbp4L9EmE1
WLIHIpEY57E25czw0mnzpVHzMr0OUunb5K/r+Rkm+HaqJi6siNOrW7rZiVgBvfk2
fMB97C27LKBp38odTD+u3s964DHOUiueze2oMbf0ak0DrWlo7H9sK4WEn8ueleU0
Uyy9QP1ih8XV1gWhInZkYh8SXDBJpgaXXQvi6X95SECLZduVxUag6ZvBvG+Zt3oM
cG+9KmZ+iAgpHYUm+t7U8sJEwIAk+ABbrmHlilkljgJIx83aSccidcrdyB6emisg
fqs0fpqtJx+2un1XZjvUieihZEb10DGhT3Z8AvWdnm73dcGAVrZDvXG27DsYjcsg
ZFbkIwaBopyQlijR2AUBibMwkrJ2o7I2XVobyxBzMOvCObg447b9RKhv5tfZuJps
XxjdU+WdptGSKvuGNU4LEBmNcwCqPggx/rIh1V7NsX7FTS1XK3Me1cgOZJkYfd8I
ptg0oN70NGfa4YAIj5qARfri4niACOk1hAo1qJ9VPdfyJAhCPf4qBqWP8AFfrUZP
mzjBLB5ldIHeGtyteirOmlsc8wyEhnIzWY07f0mNsSgafTbLzrqbX9eGP5L8LdNl
3NyI+iZa+qffuCEeB9xgwYMaQZ5TxDe0PQ+nLWSJH77Sm7M9ABTrmekVq+Y73/q6
Ot66NW7emsX3hYzrdys2+R09Hx8APmPX0eb3Zmmf00cFTO/Ssro2sbco2p0qyfMR
4U4NkPVocJF4NOLfQLIMUzbX+EyLExvqB+ZRV2Qn84vRCQUAnrLcV4qkFN0s/ZlQ
L2+tzBShzRC6yBnSk5rWLE76ufOStGW4gVfTMvu2CUOAyC5nVnWjx1IwMI8yGKWj
g4bltLp/Jd/vbwCm3cAKU+loL89nqfOxaNQD8rxuzooCNzwhJ6dS/HPvMXyPOQwB
+buIRvYUcqn5j3cUFOLC0qmNFb1VZEPuFZSC4PDdX5GY57NMOXJqGY08dAf+WasC
dUsQWyWATGNUvZZ6RJHlt8r0cbj6Gwmeg8irLHSBl4LSdYI6fUk2bzNq/WBaBzSW
89VETCJiPX99JlgaooGyXiGt+OvjInajLo1+P1XSRNcuZO4ipX3ZSdNeWryBMaIH
0zlZ+0TPUE5tZe3l3AOCq/3/WYKeZkS0ehvXtdAd/Hbby57dq/AVquxqwvA3T5PG
ckE14fmIuBXPMwW8L3EpVMVbJzk0yCABRgattQagczPYt2IgT+yHhBbQ8GU4wKNS
skOS0u7l6adeKRENiyQ10uL4XO+qoOWw9UIGNZxMyQnYy5lAPysa2sekksjcx1hO
N2hOiRKTrOBV7TS/z3IsE4PyDDYXJV39NFbV2XGc13RnqwBUeG9fRwEcJA+P+0tX
FwFITJD51RZtlrQJzqXnyatjlZd7zdgxjyJhisbaG1hMyPDy5nJzntpRlvhtu/ZN
UPePtZ4KEMAzXBBPgZqnqOdnzk6bZdGAUhoHz8B7sce9aZ3rAjmKe+d1qSiSaYnv
eBwJi0+fSjcWOGkbX43ADo000ectJcQwz05jWlSN7ZM7KSaWi4Bz388LxbvjGEHX
+cGTFJhfEUi6bMApCJN+0PRYAsJg76NuGraEyu2gYKU773VS8irafOwGAvfU0QzT
Hpnom+cUl/QiB/YlAl/gYyZFIF+qeqz0Nh7zvhrk9eiyDB5F5owUqa1QzBkmNPT6
S9oyN/1eoSXPcOjbwJ6UV7PPrzFkRbdIVObTLzy+ybdrIi9XnwtGkj3wa+xY6jrl
ClXfarhVfwOjFT4Zi67YPAT/mrmSMJRWjvrraI192MyiTcxZFb3j3ojNgxgxpd8f
Is1FYrdq/5SpYt5lNLisFj7BsR5TjI5XYQ8yj6AleHZNTRDfnmubk0fjRCTX4isy
YqKkNSDyt4reJ2Eq5cWlyUw5/YoQuX/12TljBsZmdUieQNTCggGozL8QPMHYtKTb
DvJ/J7kCG9erMJFJrPoqoClEnDX72DLeJmS//3PRqh/g4bH1As+fv+AgBLwAHtas
28MKsrAwQMTru93Ahke8FvMp3wRSdDLNVVYfOMBDlCoMF0J7Wb9UuwwST67YRR//
HDwBznds9N6wgm/Gi7+RTGIFk7kGLWx2/+S5N/sdG7wR852kJW+XW3Egb/qe4FT3
fqiDtRGoLy7WpCHhVI7M6ZYXR+DFiPUNKSBuX95zNEQAJ7Vf6J/0VQizWIkrbNKk
6r9YXg+2tA4GsgDVRr1w/X7pIVpGrhRZzTenXVV9ACCBfzbCzRWUxNCw8wp94FOj
isJlJwZfRW38UJKPFSf+n1LR8pTaBEhinm5NReUw6TTz/qETQ/Q+PqCz43CgBeUf
0N0xj93pz3hj2GPCte4svGv3LeZDiVhpjQztWZR1w5TJRO0gFB2lNs1O+LTSZp4w
Z6RzgxtRiIMHGSsnCXllywsbSG7a0ICdPSZd9kO3ftV6mavpFufg8FZKJ+F7wAD1
+P60qddB4lFIx2N+dOTLurtTYYIRgJAGwuTHuHZPdKb8Q6Kxg4wRCoQbX18kHwZ1
6YRTOcI4bK574z+Vof9noh/JSEhY8FZ7p5e0TEp/6J/uMxRpOa2H+HWg0L9lNAba
SmGPQ/mf9qyOLzWM+37IlrwVCxvh02grHdmv3TEnD6EuEF7AaCGxvM/axvGFEhv0
lCwJ/ZisQoYoZ5Bub+vGSjz2Q3hm6SWfayT8TsbEF3RYYXT7JVIqXNjiUDVOKWuk
qo3wNwADiCZA7F9wKJ5WJM9iD1NaLJkrzLJg/iriEpgMcUCxlz/n81SR9iNKxjA7
aIwj7gsheWQVNgBVGYs5QdCsI1GxnMJHgN7ZnLflUvUYqvO91+KB1hNMtirbV9PF
j6HSRp6uROauKTGnRuWGBKCQm3xIlmNAiEGT4ucq9w6bR7lttz1n7itZPGmvEPcS
qhulVO0nsuH5FDphp/0gXtLU7qKc+XmlvOAdt+qy3nrVo70GRovQw5ol+J2fdle8
nmzaDx7/HezMFkW4adKIu8txi5oJtRIGp49czYMT9JDHulXhsm20u+atT3+TpglA
4qrAxEat6NICA6CbHDxRpoYORyTyIyWhJtbj/eF6WTXhbaT54bocXGfzF19d+0x8
ghspmd6PYfW/ScbhO7U/arJUVf6ShsNJLDOVYgSpuXUQPhYo9fcFvrnmonGpMUpS
j+o1PLa0Su2yPr0kp9ocf23FPK6zVrdaYTp+fkYu40XwR+QBjOoTbw/rIM3JbcLL
HyaZGjm0tmF8LqDFU/N0et7fB7jVAs3IAftbHdCKvFsd20FnlW9YWz+M4MEUCiHW
48Z27b+1T8OP3Jv54z7jIdfUm+irgIFZJBwqoAEAEE0e7n4TQ6KedaCkiuu4Bqux
2CHGKg8jrCKcniSDej/73B6VhekKfgKEGyLlItxjahqsH78MeNO9b4YUGjqtt5PK
NU3VnQMSiKBR5unxatZdH2yV0uPo/cW1fFsFREHvRavf41E8fVsn3XKkhaDGJ6cj
Gyvyerx43kJwD0In5afkdEknr8fkL27Eif9tFmEk4Ttd2QdqZkcQV1rdOHTmb4en
NLNScu+GtQDWAbeOuOMDI+w69JkXrweZRqxU4LQAX08ivpfsfF6gO6F0v8p6TCRX
dkN/tRH9fBn3iaeZz/HZTtN22+Klwnzz/EaBF6S6GYV1N7c09XvGLzWKo2p7bRW/
lTxtZbDNpuWCOQuc4zEfeAFsPLDzYR8cFyMYGx/Ji3N7t2H5zN855weTlZGjR69W
hsFYxlE0T1ZlTsfv3YOd3brDVNOudTv16XKu+w4y965lefpEMlgwzDIEhIWOtrJd
1HjA8SkYjYNGdkasLnGw22pBGYQpFi9aGauVyyEucKenntRgMEusqoQQCnul+ZGO
01wPvNKty7EILKY7ImD0JZx/fILW/nK/zUhzbjgnFS6mX5boytVwvoapIOozv2/h
twv8vAqynAj0euqSlYUgdnLz7mDQqSJgjhhaDH28hgIsvACSFujXMm+lH7k8xLTq
kEZafqDGy54zTWRstcRmvhRLRdfna2IM7PHeH/+BUpfHBnew8dpsBVZ3X0ePjxCE
m0tBKn4PsIbfZcHK+7Ls6M8gTJoTm6oXAm35hxb7XOwoKykGec4CPkVUqGBBMhMM
8gnCTDCnlI1xHWdAWZPRpG+hkUQBriS7TBV0VGCiFMaMJ+56BYZIMnlrMTDSRICl
myMZu8m0+x9VxTOck5EAF4E/xBJue5JbnEDuDNapwGt9w5knRhrb0dB9SXlB+Vk4
Y9OBn12fjrQyIDLYMICvUM42j/I5isFvSQinKH0tGoZ6mwvynx8pPmNkWe4/qnGi
t1JBN1BDPMlAqWNnn6ZJQ6Prey4MhTRyElWVcuqilUfPf3KMLQCCiFDOwDYbNVfk
4eFthDFXCPIhEmVgSB6ONEKnOgBjIaqHMixF15efxUmixC8WjaNUrMQPazlZq4x9
ORzKut1dDl0pKxz2bTp6OxpzIgvq8F9ueSKM/+Wj9Hh2x14rRDxlEyDDtTRlq6nq
6d5eQdydwJtZp6YuyZ7o9nSQ0N/AaE+Umppo70X05OBFqdcuYd8mSP/kqN2T+fdM
0TrhW3r41yCAIHVmKhg0Hdiqlmr/mgb1Z9gHJRSDVH5OnpEPhb4xL7BGn1/Nc8yq
B6oDr5W9rpRe7dmNZdaOrE0Rbx2nFSaYKEDxFuDTNZVG70k3zd6HGgWR5ZSj2SrC
RuwdDguBD8I/eQnNkwx3uh5Apx8j70AWWOpUDfzMvvT4YL65xAa8RlMFpNVQyye0
ii79mgzohle7ZpcdPa1SwE/6GsXQuxJHn0ZKrcItUCE1i++Z1WbF3r+R8ErlWRU4
Ujj/RXc2qNu/tD6pk6goBNjt2oQHBFkjPpGvT2d3Z3KYVRe45QFxkIPM9SN4KJeb
gg6w3q62kM5rqF67jmMIXe2RWqYsbvXS8McnBkf9PiogcN6JLQ1j0QKQxqXOZIiC
zPVJvNS3XXi8ORvVjfq56r+lOs4kv3tbomF742gGhtEbBf7QFwctjABHXU4efSqJ
qUaWLAVCuNt3EYci0GfQEney6lJfi+PkXdqoeEvi+m/2R1/XjuooKMJjlpX4ay2l
wS2Vx/I0mJ5CUTfnOU9yRO9lRvYltKEXw2M99LKzvuHnxh01ky/Hjc50NeUbK1W/
5BGcjMHBmB8XujS2fVzX52mR7sjM/fODyoEnx9E6FGdAAzKSpmN2IG8WgUoj7FmV
bDqKeQsFT2AIUyyu670PODV0osmR6P0qqgyJy6UjDkI4UHJhRVY6IhKIfF//x+zN
DO9467/uRW4DzpHjsrTdHqTQ0rIJCGUOcO64cjbrNLUESqzwg2QcP8Q1/u44xhMN
1b6tVLaWuBVnsTTdkieCNyBQu8D6TGuZs/lA79hVHo25e497N2Zx7Tr4Fl6nI+Zo
4ptnj4SOjXw+9Y9ok8Jjx6DhnTZRtuDx+R/Ug+5cTFIPRPr5nvGmfIg0cZe28zyu
zktqP/rg9TK7DfETB6Q5due1dAH8yZTSTrRZRTZrtFAG2ZRtfdv8+K7FLoKhgZNf
m79/JmiXTrYyu6eca97R44SOCJpUHKAOVtc7MTmDUhk0ZGEYSDb6q/lKKIizCag2
gyO9tsiSv4mNxsrTNnzfeOM+oJN1ehQoEcbPWh9R2sCbmD469AC0pkP6aNKrSlnl
vDFlICXl1C/Te+6lZGnUuhrG0isHxUeDqwxhoDAM3gr66YL/kpdYB629H5BbSy0J
hAtA4ww2fsjRuCVadFsVu9f9xXm20MZgRvtk3hOABH0P0ZX4ic8l8WvQcdUQ4i7P
cSedreC6h+Kf2FOHSemqKzY0RoYKLiGDRZJEhj1vxQ2LKAmIEkcZwGsLVtrEyhok
oe573MO0aU39zo/5kXP6zhh4N5AdAqOfSuoTt6UUMI+GsN+HmGRW+NugcHgVxXpB
2tMjGcwJlLiJWlEQHAbBESkqsyQnq3mOxP6hDjW3KrPBJKH92yMYkYXFnEx4K0MJ
BSOCVzBT5ySWCXr1lYjfxovClbY7NfLt26SiM6R8cNCt/4zVI1Qy4/qg5a8K1oSI
2lGajYJtTXjSZwzB/ycNTPHum5GFWfWA2gUtXB0c2HK8Ua9duKnFw8YkumZFUEZm
sowimPHhva6YGx3C+T6ch8Rwt+quisWAHfKE1Ynsw2qKahdfw4uVt3tXYjhJbNR7
x8o5Ul2mJB0hb46K6eMFqpKnL5gOc8On4yZq5GBIV0IjPP9DFdBSvxQP6AHcqjD6
UxaY8X9nOo1EX1f160h6kgs2nZ2yy5dvSMC8QZCskOCS4xCLunqWL39BKOAmF6l7
Wsao3zWc0iXNg4uB8gAR1b+IHh2IKxXenn6LK6krc5T5u8yOtYwROm/el7Dq8kKx
dzup7q3tPO92oTEfg8i6+oGu8km8ZotWx4tIbxjU286zZhqKaHkVWZqEVo5XS2KD
TQvLAtAcV386c0HqiGHJzoKFGJYAssG/nnb9SSdBbZFHguygTgpIp0LrCMK8Z4WQ
g62260ntR070EYIpG8QRX52M/lphEOq7+F9V9rqwJMUZUfKr+T9cyC160hRCmd/Q
dSAEyiNtUE91OTn9vDOgMrCa7n2VK7BYeDMquHQdBg65uDTCRgcKOU00kywwe/t5
fqo1wF8UPxiCWubiExFJd4snPXWdQJAiJSjwUUp4TCahTwaPJkHKkLPzeXIiEYA0
PcofdEpb/IfHedKLWyRaCXxvxw3MjtVfp5DJH6y0a4W8YQDn7+kOcSai/OWt7twT
IVymStm7neemHVuptgtCeHdm0R66xQhXQKVVVSSv68W/6Bqd9Tfck7bgNNy76dRq
zgXjwt6/qN2OefDOp5T6KZqRzdn9UrGALVTKxPllVlBb/33rCVuOOeCuly8nM0qO
Qf0zehDQPqCddadyoPvsuINWomqwAp71bIe6zOb1+LZnTeKlnoepLAgvWnFAxoRw
mypaPndTO+xDhF26/rKQaJ7dwTUap+b4ksj27SHx3yt1Qf9rp7jA4Lee4AglZRv4
ZLqRkMsoxEx9OM1pEa8cRKrUWoSf1uikctw4qU3Nu951fejC36pubSRuvxjNZsIZ
ne4kTgdicVw8OHa2uiKYKqN0BGm6Hua9YAjZwD+gFA27QR7+2VrmCH1TQTc68gzz
iThjU3Tc5aA60C4SB6Kp619wCyaag/4oQ6+csw3Fg1RHrytFX0c+t+vtbSNDxdrX
Ou+TbOKlBbty0F58XYpWOzxUr0WvtHT9Ls/AH2NxL7XyrabpSAuRNHdQVSLhUSMc
2WgzabgBIx1awJEWO3QOQ+gl0m5Rusr5DohnlT/puJd1vtD0MQG2IUqv5FHxKYMS
4Bh3k0QKsZYkkB+MAIOTkyqdTM9VQIIlj29n9FBp+hC4t5Ox3nj7ME0nzfChHSqI
OxdtJwvCkkhgvoTTp2pQGZ332lYEwTUX2US7B/7Zb03om7fp81HpvJ/xEN2d8KfK
uHBZAbND658lWCn2kMbAySJNKBpUlUn1ZLDIPADOwzoSaJxtwSCbPxNpsc2KBvrX
6xoTjLppvcoglt+L6htWEG7B9m1o6AaZcd+dg8BZ2TBjQUfzZjGJ+H94+1nDQO3n
aGI0iBnfcvHVzaaIjCiz98fbIPoIKu8M/VDCvWz/+LxXnAjBwLDjL/t4kh7UdVV2
6PuiwRaBsNtsRiUCzhXnp87Xen/NZHOB/8h1FEwVng3BdnkuylaGW0Szp9Fvhbg1
RxDSwjVCbq5oyoYECaNbs4pdOhNpIwIDqpFXhUcdB/Bb57DIagCmu+wKECwrFTre
hPRnt31Xo053Cs52EOVBrkXQ5AzEbUnY4jQ8GC6RtX6ziH4jdmtcc9EEzlUa5GfK
h+YP2GRZR9RF8z9IRX7uY/lQKmoExomuq/vCj0za2qJxbSTQaIhL44EP2jq/zZrj
fFzxaejm/gBsV7kpHVr6cnzrAETRQtSlIRWXhhAPiOjKWN3/UcnzzLE3INic2DTV
HA9rptyAWep7Yt9EyMXWHIDuRTPGfVnupn2AbyU3eWDslS+lK+4zMoftCynQagKY
4IyzPBTBnnT+ERZw+dFi/mgNVWV121nOb081emNQZTtZfTeJ9dnGTz40GB243rZP
DwuDEBavptsgJDYadgBsY8dKUeEu467DesSCL/RBpb/7nSHeSHpIuGa4eIzUNFWy
x3rChbly0xDfKrfBhzVM/Y0wsU7540IQ/VXEPfvxrUo8xJJ9h8SFy40uxnP3yc+p
DACueEJzGoykqydE6BnID6fVN5o/H0eyNvk2TDltykM/c59oZxh949ngreMZrTNg
oxGx+g+PBu2ajx6wrVo+D7i+MthO20sJs3L9in/DFcwUojDaalkO4NC8zn1RzwCI
wgXaKqnY5D8gSynN3JScGOBY/EJr6VIep0+IQRhSf1Wid7Wcw0MoZ6lceXBcMz7U
AvXCl3C2l/KodlhzDyIclyyvIPbsd0WtRcAVQdcAef5CapUsxCgP/+Pe865vZNC9
qCnPuPaS5uNAqTc2ompqT5Xo0TPT8OEMbl6kOuuKTL148JKSu9tLqzbK/6e3Rq3+
IqtuQO6sIid3ie/T3GS880/VbPSYQCT3EiD9J6C2rvJOdwxtX3ZwCL1CRZyyw/az
AMUHOHyOiP/kUUiI+HiillBNw/dOhDYKSO++suMpRot2lGbjN6uVvDiXKXFE52JX
/D1KoFPxFONaK+FebYUDK8eslOXk3fWvrHPadlaXguSeAqT0uSCVd8xzV5I1GWM+
Iv7K/mohzjqD1E/ogPuQFP025ne1I4jzfNZgCRX2DhTUo0Z8A2DGgnICM2neajsk
6/efTNGEqMhMo+5HkseiXGnXNbLaJAAsDpvhZdJrsU/JOaEN6rYkqNs2lSk/hxhT
NQULypbURajd1bq3WWwhhcXWyfRpoW2nj28uH5XV2CqrZAJcCXctQCKQBXbb1Rzu
Gz+1EmLfvMGjdrF2MtNxEkuj6OY0CR7g4rrC27mBLdV1iiYNpq6tDJBEYdfcdRF9
kk4zvvIPAkxgOBdw8UlimJvHp/Q9troRDhMwzY3RsYjAxvghq8DcZKwm8C/5GAUM
lEF7rq9/FKjehO3YbIr6NBh8PDuH5lG5WrAD7uKXArQXtmtW3BsDQhZ8P0fHdupw
QwW1uHZM3bfD3WcQSEQnAZGMkv3pUqe7MJSaRCAAVTJV0rysZgapXFau4/ykZ5gY
M0EgwA4yTeWB0qQMg+zAqf/4wvvwGYWAFmSiTGh2U8m0Wxovai7lUQfdvXw+I6d1
F7EMBf0+QpjltmrOse7rpsLWaoQK/90Y+iYxEqNAKzxUYy+NvjUhtgFF6hDd9aD6
D1mv9YSGIAGW3eEomW8avroR9oe5MYii7jXmOVSkSml5KqtldudBcV+3HsZvpap6
qpB+3ndWt2lrHhKvYpIxut7Y8zkWMqVd7d1+OQSRcV1VIde+LSa8+Bucpb/gBwvC
EMM/0xzhDIqw+t/N1sgUV+S0d+1HI0n37Jd29GVYDGuYr+VW7jSRsJgqW7E8wCQj
IBYG+TNxDelw8tOyurr6EnMFtzzQ6dhL95W693QMVlDpj1zNRDzD8WS70c9063n+
6eT0oLsN5sEbQMBK4ThgiD0dIjfR7fJtafRWBjnm2thzx5gASc0P0UQKdfIMQqJw
0a+Uq+WTdmbQX0Snb37KumFDxM+WV/nnwXebWbB5qNCmGVUZIPhd/xt4gMmTzNuQ
Mhl2YfRgKAVGG5w4s7/CJOJVZbA0Dq4FOOYBtUOHH8NiWhYr3wrsL0uHXE7Y3oHJ
x7HxwjzMmso1Wjn3N23ZOCZ6Us2HrksqtLHWnEY9Jxz+81G8rPS9ycgAHkGYsgFz
doOMzyJ6LIAw7Dr451KSngLwFltnTb+FXOsSl4Ddgfcql5eb0w5NN3D2V+/db7Mf
PQw2Y+aD4R3V+uYY42CkHyOcaIHNqcUHXRQCsO54VKgtfD8QC3/YxsReJmkR7w3o
qWI4Lf7AyobVDXIsV/prKb59psUZlWY6457hmhnko43Im/fZgyINEu3OUHefB8t1
OJ8LqVpyjmvnvNPQPo2OxjfEsoaRfV4s9YUUsEy5lyWU4Lu0PNEXkDjLWHK10rvC
P0AaJ1+Ww0dkfEUfA49OGkB0FJqz076o0RhwFWkfutIxcwgsehGo6t7gNBTrgizW
JbztIoNUjxPbogwcBU8tiTX+d/9kj3jqYSVbWCAeuhF6c5dlgNTOUKTV2y2q2YlU
tSHU5bTgYC2Yeeim9vZ7JdqgiA7BUSr/Sc/cEAQhzBr9XsMzCz8ofLYrNodZBud0
lVgARB91fnmmlbXkBWXsC4kCEEev2eQg5i1sb6QeNAl5rv7hLzDwU5BQ+0xwJc1B
qex//k9avZb8kbwAtp5DYPl5ekIEM+Qc4h8XRgUqZuzl6QgUOOwXG6fZ6FUwcwKs
rGhi6vQCwar30e81gM8GB6hFyovXzP1XKIqvuOA2gGNiDh1QGCiw3Kki0uTYsDNZ
poIeqqgOWvga5qWrdemF7nzXib99p3kNhcxkzLGQqLkOZSVCuOJw8h5JdvBHqD/U
up+VvAfWSW1njV2LGBidYsTRBKmxHgFO1fngjxXZIClxFequSzi5xfqAsQit1UVU
Ex9f+KSqtXvwLT04kM1x9olDqyzY7WqRm51+yVKqNQICqw1199ZYTRek+td6WTRQ
uZpxfSOj1ClbY4zxhnwMSZSGV98egBbXeeDucDo3eJ7pNic5r+GFIkQlbLv5KFcY
87d0EX3xA72MeCX4tJXhD1lmPjX2qom0Jq0jJht3jzoOlAF+mjH6aIWWiR91aRqA
Ne2h5savBLRAQZPgkZIH9QfXmrC1vqNVNd10JKvJ7x8T+zSM5ISgZqANnAn0q5Da
Y/WoA0HRUPuMJqWOhSNQH5KVzp7cDW9ROhB6j55EgSV3oUoln2ulkdxQvolJrLlw
9RF3TkQeNWLTkQErpcmMKS9gFtP5WxBrTO7RO6gZHCbdetRwtfkm3UJJ8BTr8cN4
hCUINfIXfAjEf4ROLyPH7FH1oTvViQsBTdxBGusmivF8pMq813i10Rpf+I1BujQM
lYrjatTHS5N3Pk+6ki2R0w3cODtHgn/hNLRgXvD1qiK6DbEY3acnKZxcSgKq5D5T
oAyIRiuBv2Cmoan014wHNi9AqxMKz6lLTxiqhJifHKpqgiYkxptJVmVaHAmbhJkD
a7EU8rxFMrF7c4iv5m+MKBuA4SXxL/pdPC/IO/Cx/5wNb+JPOSHApbMNUVoFaEBb
4G85NMQ9CztllHbfDfOuh/FF3Iw1U+UnS3P40QDZ0YCPXkwT4SKV9yLsBtSFKqKI
RmzMX9odD8jdr9UuIgWYnkQw6yY4wPQf9diS1fPsTR3BbiZ+sr1G1H5fnosucdLS
i7YlSsoDwaqFg4Fkz/RSUeD/igDtwBKg8MssDg2ehhw4DKPs7Y9oHMCZ1NzXSnZt
vTKk9PdOKQK3WDrr65O1T9xu1zm6P1adU1Lov6b+yAil+7irDu320xrYegBqDD7h
hHArhaDWgb+0bQhqCRz/Re5McrTs4UipP54QkQUbPpl+RPVjg6VMVkaMG6MkLvnG
4cFt8WqCS/EY8KT7pShReE52owAyI2Z/L5tZAz9Bqw9rUGcS+02JcVeq9xR+ip58
uKT4b9VDhWUB/WA2jZww1rJxDff77xhxoqL2OESWzWOK0CcKHSF0yIDIxJcB/pbH
x06QHXuK8AMst1Xh2QzIhEKkvNKCXNa+7JcemQs44tknzs2e7RV38k3lzy228yL+
uNw46fMoQCBDqBwML0lKQpswzJlg67MWOH86Zl+XlVEC83FuKfoLNFGMpEfEkDNn
UAjzU/Ft8RIQgJUZBxibgSpfHwXRRYsMu7ZPYFf7QWNkKeA/d6h/12VmJ/L5qJmW
sOeo2NCIE++PzJdh0lbrvAEG+l9CoMhHLfFHXr1u+K+Z5O/5sIkojkB95+VeREiv
NAwD6GMSn1iD7fxFKveGjw+zLkEi8ViQEMOiYzu1hR4HRQBSP75kU5d7vbUZslGT
f3n4BuCWI/HvXJ+nFTcLJi/6MK1LwIRUpa7ZEWOgG7exmSl5eWUhfTEEeANgEkte
0yT8PjcsFraF006qMSRQPDXfjCh0wn/HcE+XxTy8UBEOU1ypHjeEyKpEybdbmw/h
dMuSYzbktktg0dYpE8ogOIDeS3iBeBbARxpXbHXjD6T8sXRrqDdQGk2dsJYwbvzK
oyXLgQgslDveCgdo1AciNZlRSfv5rLH9N1+T2rSwkt4sVJ8viF/cGzOI2uLLWQyu
RYdq9tIe9lUYrGztzbid2PESUb+T2YtvIPlFidMHoPObPwQk2/cSGVkflxMijHYt
bKZmt8bepyRa5y7zJvi0tFQe501nVrNDo5pieYcE6k6nieSg/6UFCF3FgcExYtVN
VG5wHR8H6zsada8vytjNdVcn+Rk+HRfseB6pO5pKL5QgMwwZ7+uonL4x0nWKD466
7rEFs9wQoqSp5vXBEzWSvo6CQ0fg20XnlS5eI6EEuShEyB73YcGozL79UZYtgPTC
3dpuuwpf6KnXIOcEADTVmkgEyRDc2LGekmKkFVYnGFfeeFkrBaiXOeJPtIblYXD5
e+Y8WcpFL6UJIVSmVhYHUJCWNDcMN3F5vHnkE7rRV+hYDhRw7SB1kVIEY4Vd2J1I
tWnes1CW4hpyNDYWsRD1f0iwDv0boAL/OdlJowl7H9+HDMluZXetZ+NDHRVEnMpb
KqiCZhwsw5GFd42a5rrNFvb6lmW1UkEZejTqIauvid710DYql+pnrcU2fMfBoZlB
g4HlBKC0O/cbwAMXs6nI+yeVx29h0Hnu+Iyy725VZV2FHQcLq7TSIXuDmWrI0Cq9
QFTv/OniWfHQRYoAs0PtggCXOKRR5FAbwc6Ggznur2i8FBhFbRoLTig6vSwMiYNB
lSTXBRVgIrrL6emmnypn2LrNyhAI4KLkbkcywEltY5EgoLp4Jy6vfbe0vPVug/N8
9pLdNjbO1N4M56VJnpHuhL8If84jSiLEZVbARFEDgx0fQ+vioLuc3kQQYjsVAupm
kQsIZWRBZZr4rIdpw2MahHOWavN0wwBQmoHF5RWFfgmSecYt8aRhqRYxNMZ6JFV2
cTDd07NbsmrlbgymYO8qbhCqD412vJSBl/oa7NBXOQ+77OjnrTHvhY9eW+sJiwFi
6NXNlWPm8e2PdAkHfJnobPiJIvd9Ui9U972iCS+dX8bER2MYeGbVDuRJDPDDPenT
LitOnh4+1TiAbX8HtJS2OCWZ+WO0Cgzsip+tzXwgWP36s6IgH2zDKZ/7KcNg0A1Z
vZG6ENw/OQq8ESKtu4H6NgcLUf9Np6pmL+cYj4YpY3Z4/hrEaTxfyQUVn34fLIWz
msz3IX/fUUqNRF92WXdiuIKQ3CMnhsjnP3G6GuP++mde6XYwaI7/4ta2ET+nTaKX
CCglB1pnNFKMLHFxa8drEXDS845BVx9ubE3Q+x7vkMPFYfv7dfl0wHdAv5QSZjc/
d3P6M/VQHtOP7g+XWRhIfVQzyQxdp1qP4IfP3EdpvMfOReX4fa1Iz5FsMk+JRJtE
xADQohH/1fzEqzg+ktmF4NNOfAvMKbZJD6KdP+TScBpTsQdGtO+ylT/xT4MBJH0A
yEBOGjCmRn6OBeXvhjbVgmRpXO3TIPp6bwGy2Y8t6hCg0EmXW3NBKoyAVWdQz9nB
Nxrq8W8syLMwquv82kvICKIj/zBhuq52eBeBKt2KTwFDnfhjYM4kRD532baqGk8c
iW+2EdgN33DNs1bLM5+9AMhbciylR3RqBqcbpwDDVG61DCqXl7H6R7YydnBIwrc9
OvG/2IAM+9bRVMzT6SeEp9gk7Rs62OX7WTPr5GKh1U0fmZgUkjJK3dq1vGjF9nW2
6aE1d6rzdh83hOpT56McG53wqH6Y7Obcw6XuUpRGtR3YJ22nevRWuftYg9NakWSp
OycWhkFrgZCCNdkt6xhPOpnchP+SDfDU4BDjuHFHx2nGYpnhJnAnWNdtd2FWcoUn
tQ1gN2IdjTAT7xg5p/eXGQL9WEkIUBmT9GINRBc/JilKnDwyq6RLzObidl01mWa0
VcXHetnkCGhiCbSpPS5spvt7dwtEArF9bC2PYOQC/vy3jQ+zxGvP2XJSh7xtDLfq
ukvK5YSh0oJ5GJWf4CGL6Vua1WCXwG7yFcurU+GeOWQPMLqkryWXZVI0eZY65k9y
qkfPiXbKO/E8JaavOtT/AVMmtWCuILgAkfZvTK4bq/0GcPF7efQBspEyidIlljRB
xzjV5Vvgv1VnA4vJIpAgn74Z5zy7carOR2wbOEAN0kU5v1BkjYbos2U3pWVbb4xK
FgdUSgJ6NgLXdxs7zau0arEKCpIhiWoG6iOR8plksVw1QRkifjSOrBxJgZekVQOH
rC24b9Ja32gUr8dkx/JG0vo7/CBpW6p/TX7rxHevGRjPgk1UK7xvntxt7WH7LdO0
OrAiNQUid4gRTSCmTj9VRMJGLnJcV4JsPxAZkBEbTz2w23qzAsUJ5s19giaXw2qQ
h/t5I67G7WkiGwLlpnawy9kNk14nUjvK5mCzZNs5FJkKWiku8qWR2vb0koFT78Zb
jXZNdAGFdlKERVcDHssdwLwrBnWmurKuz4inItW5LzduCYnAj5Gao/yIG6xVVaUG
AHGh9UIUCxnSl4FWD/Hf+Sam+am8p0FgIVQkr5ZoQWAvVxuzWDVZ4EkyN3MCOKCK
Gb6gLB/Oevn7G5J8ZQl+WBcez33GZU4p09Hang1PnEWATA5W3LfdtwfLmtESdMiJ
3btO6i91k/HXo+U/eTaE7Tl2T7tDuPbZQ6cVmY5e4mpSEk6YLlOyX8uwgQEZMXYe
HXM0lCuG1P55nYshdxSYqEnkAeExjhlidOoSvgcFRy1wM7OGe8gDzjvNPzBWVcmZ
NHqD+rb3I+OoynpNltkBoUY3tt3QipF48MpFk2YL3vXCjTM7U60COXp28Mhko1S1
mSCGL9inYH7rk+mWp0/ycJVITmQaJzWoBCmrSrQDpgYBn6UfMx9ot3Iy7CFR8o3Y
5pzCP6s92aDYv7bZo48M1UNPQSxY05w07ZmXERLYQg+9EH58LCyRZSXnSlmgcPA6
WEAq5Rfd4SgTCItjSUG8gDXZaA8yi5j3f9J39bSwsVsRRrs2FkvJAxuKWosk/j02
IZPFZMXFtzSKyS4XKx3LXuZwqRx4FS/pydsfsP/LIPe1M1Kf41Yw2Va2T9PM4C4z
8w7S9/aggkQjdNu5zEtJjM8MJVpToXybVJIJAH1L78TQWpcxm/7BHcaMjEsP/jrQ
ineEf0vUMzoyF0npdk8MrVu9EF1s5/KRGEwrJD3ImUsALCX94C3AWz22se83rquO
BDTQcKgijt+O4+aj9qtUFTT/wxt8Nu25QWzsKRERRKMirhFm1bAwEPUP+iBIQnSg
uvzycnEC5/rQh2AxDwy6o3xURznLqqDJzltOrArAP70sctcx6Q9tjlwu7Ptt+gSN
CFbyJ99bCzsbjk2CA1m9kti3RpdPPgZEXDaiTNA5mta9TKxJ9xgR4nVOaq87iEFc
HJE0y/5EJljXP7m0dCv4PqllRnYt7VFkeEojxJ+DX6z0wtAuYIjkDUPNQ+OwwYjb
6aq+kVUEhYDoi3I+fpEJZTV8UVfTeIsK5nKI7tO6P2w0giN0YxVhc62KBwr1sqAt
7S1MOmoh0bKD1AFoNxXVeLG89a9+gGFuFaIfWVxM3qaCmvZqRiZVGuYl810Lyu2I
MEIqyO+VazFlJn8p7/3gXPN2Vx73m6eAXpmr9NZjw5tV7DxJd5duJz+zOOIgvr0+
FsQUcSMi5eoWZEpGFS9T1++gHjFbsxVDrYA+xTn+Yci54o8LX4VOBW7GRDUzXeBq
6a901ALv0Yp4xCCSN+VL6eVtjMgDIqjr9gOqhWXl5re7eX/hQVRo6YmUnjQkjgSr
JMSzqJtnYBfTa6LkNWUWQFA9wGEWrRyXfhYPLHAdAJp/lYizHtmFX8fp7U3w0i46
5+T/NMf/sQLTvnLtW8u+rAidOz8HqO17122nPNszOtJYLr4Yz3GFF8z1hGmUEqGe
WZEDO5J78zmjNKmejxQrDfyKGL3HigZ4iiVGxPPEJI7Vit62YYsqKKe99cGiYnKe
67S8em0k/nT1UkkaIR0suMQdcLYyWyVNJeuELf0z+Tb8WsZWmo/Z6aaMzWkXWi2A
uT6XkrL/KRNVDIy0mPKR88j/Pa10UQzwEr4KZpqtgFB0Rh9/vZPvYlwn5hRsYhfa
trdgwtnzVQgafz74JNHljQ2uQ9upfENseqD8KwKTja36s6ZSIcoYQ7iA8sdQBvAL
IbFweDRGqkhiDzZtGYyJ3Rc2gVH8iLNdSaYOm4e0tKSfS5InHXpZalZP4juWbXaA
rqJvHkUA9qjso15S3a+47qOjyR6lXpWt/95rOO12mV4fed34vbGuRKM1KOhLqck9
opqjhcO6eD3A0OYgszLK92WGsdhZpyFlPIzeNYWvjAwbvq5eYNUIbMOkqM0UNffl
ivadwg8n/3OdJciDbKkWTanZA8165uNIFOpDiH7iwqhU/2JivM/kQEbpMBrZAif+
GPqE7fpCaCykdpqHdAqvvz3V8kJLf1xPuIJwBktew2RqvdWwO6CtUnQ4FTa4I35P
wEmQlvhtMRkpWSLyWskg/ghFXBU3ndvI1untUVejjcoP3k8C5Xh7VW/rXKroaGn+
qSXIa+anZTDi9sRPzGtR1SlxOqY+tlafxgZnAr5c2WqcMndz5gHcShs/wKlQ29qP
6XJRXG5rGGKoIxLjkoaXBIc05eFLHuXjawhk2as/KUyD7Jl5wX4xnljo9liW2ESw
MMyDDYR/AxeuxvIpjqSvWGiYp3nLRPXbzoqeLyoz0aTcY9EuKHlDS75TLXMdL3bt
6B5bxuFGPlCLxkrtcCj55DbNuGuyOoV/eWy3pf3X/axPFwy/8yQOMCmqcVuSSkiI
iDHRbYBxvxKW4sVDNr5mtmgGrEXrMJt2QEkD7pv9u2j+v0dgJOwfxC5JzGqRmeHz
WCLlnEa5unnGaGzs3OOmeb+OdwopMw4xkcOMruCtWlHiZY0F2lCymBqYPFOVYcr8
8603YyXAC4SV5FwtEThkgaTO/SaEwfMcfPWll+h6TvnMYImbSbRKTlaipSosECYG
HPp5pF8OjIipEvy0qFeFa78bXDnn8e09dtUDIJQ6FXnOQmAD15v/SHxfJn8bZYB6
2sfy4f7Zg5jRNTalJDbeAAwZs3GT3tlCIhR/xahvZ3+SHX2KMBdjL/pq7LnVBeAx
ns//KOtwfZR1wvT1ko/UqZsi16eh4KlY1DcR09FJPurW6kxgXx26lp4eX1IzoQnb
yv+nh0ol3pSnE5Z9SgYzseV9ZLYXSWZf58WOCZcbcKlsRXdH9ReexuL6SBTY5QM0
bXxhRk9blGA+h4DGYhU1/n67lk6Z/oYjJvTmG1qE3/4y2+XeyWOpHLLwXwCpilNU
vv+MXEi7bmluEftDpIa80TkRTYA+y1t7JVheAOqUFylWqClOT6Cv9jXPlAJr4D/u
Ss64Fc6y/mCljaOL+S3u+DQkaxAL/9WaLkt7N9S1GqDEOVhGeSZsdaNdVamVMJGg
9c+EJdTN4nTJil7kNcIIwHxCh44BU6WjkYtKQUpKRTM2xlUMbBbPmtykG2cIYHJm
h8WTjFPWFhf3vfdcYSiFXIlMdIIytlO55F3lE38H7SeDtm/snlDbIuLxZKoIgHOF
NQv/iyJkPH5en0icL60m557GzmBMvBvQzDPVnH4FgdGGGxNO78PtTm7NveDUhXTI
ry9Kf4UEvIML9KT60X30oVlfqLArukL4qIfumJO4WiQLvRDyVBg0d7w6ehC8KS7u
GShzW1oq44TxglNmgvbYyYFKvcFNTI/GRb+GAXAqcbl24uASv0053NWVLO9RhYAp
PD1foCphl1gt7HxtbluppcFMoN6YUoVuMq+4iQyux4+14bRaIeR29E2ISXSCs5Ph
F/y73FsXJ1jXX7LHgtJdeh21HJ3x0fjDJuLRPKOtEdNE0JKSUTZLZDzelZaVWOIT
2p/7U/zzg3yXjHostDBdkjv7Df+MrdbZpfQ2adMxTk6zGB0AUE3TkAXNRsc4ky8G
e3MLWk7CO1H5uQny96IVj3HHyTiEed+5FpcSyr4aifSQ6mYupmmKiyzTpUg44pjG
icBHvpVtxHNud5vO/Cc//nJdU0ojHGxzDQ6jDm9tyOf3RS9wbne0yRYWp9ctBgpk
WVfgoBOWztbFwfxEj91My2j0pdJjlT8jRc3252TvniEACAn1jqxWEJg4F9f5pKWQ
rwvJ/zqm8WbitQ0f53P5jCy/QxPF2CFnzTbEDTvqyFe+vBGe3AZGe5yXZuPKm+ly
clzxev1cZm1EY9MKiryvxL8zyHIKdgHErMonYBwkYLn5CYn7g4sXUigCmlH8xgCV
Hs+Pc8WsYi+1GpWf5Ne7BAeUKJYCyT+jHhNCmw9LQY1PaaZKGN49kn5YBJemte9l
ah/8vHXejJ85667WyZWpzlMCNMMPzWTCyxsYvNQh2ckN+OOM3HUulP8ZEGTUMd5p
cv8FmSYKmRDvndnQtWQtcmpszGbMhikTVS/CqwohThjpbne9s4+bbzHVfJK8DEBB
wsy1SIbPO2mqJLlKp4liy+HaDHPKEZK1SxpnIsTRKgppPzJT4pigURMNsg6eqldB
UjZ3oEwo1EhTA7trdTOYRC1g/eyG/LEt+NyHevSn7ng+pIrQhkcT5JZi91qT4Amb
UpKkogGwJhJDPVb2aUuikTiRzm3JE3FXJSywp2rkoAQEEGkQf8FDH94ESXO6hxnY
LvDf/YkpPPQq6O/wBPJVY1o9lVwEo3WicmBzT7qdl7jcAT3GrwvQHqmIqOom88Cr
La25w+F19Nr7cqqzZgtbeSpygK7b4qINTvO1BZAv+UwYHxEUPY9n/uJKB1MrgGlB
RffcyIqTiZuk8/qmbuuhQyM2ZcYRNSc/fT4oSsHc2fpMykyHXfaO+ywtPVxn94yc
ID17eM8jgx8cV2CDjlrx4IYY/Jg2vMCA8fzB7O6ZJ2GhHt2pKFH3mvlcJBWgR/G3
dCqchzwKM5i+0l7c2B83TGi+lk9MxQKzNwAgX4DcY50ej4HMSJVJZfhvzGQbfy5q
7LiYotnW0Q9lPEpsg7wNDapHqj4yIF0dBIQte8EiLzzEP5urBaBd/aZOudLC/pvM
2u0DOJ60vy630k2Uda96pSswnpUXVtI9VYoqdfFlBy+6B3vcFyV7UgZrZXFi6W0w
JvyWX1cv7bvTnJm1gUkN/zDMDVGegtpaaK4pCk6BIait/sn4OBzJXxPQrfGu6AAe
9ShxI9DgSoZyXrWn6vys8kSde8AbUSrhCM7nVu5YZ3FRL7C1oYxjXnt2xTRtIf3M
lVp4r4k/bXj/dpqk+SsG9jC128THXJahqBXfdGYoUjHtl5EufEsrAh6UeR5SKwy4
FAkeIzpJnhpzIkr3QuqtHq8J4N/5Sra1N8NINosgK8I+sBTZq6762ZvjOJcPXSvC
5ITKp+MSVyaPgVhvGgK7vm1SkqUj8PMKNWKPoocowKnlzQlGxE6B2JnMkLWCcxDK
BUeHJpYk6TnQRSmb+nkvA9SmdCjpcFIgI9YRK3QvRHj0ahb5wCN+lGuCnKOONcqv
LwLcM0z7AZ0NlWLJxiP8bP9EmkTWls/PlewyZcF6+AC0oMxFhDc6UAYEQOrhpwDR
A78nnyprFAkWmObsgW6WoKQWn4ltoXSxn7rS8cJaYS6DMldbHayrakAvSCzFA35Y
4C2roPaa01P2JzSWwoRquHkpdGk0HplWUB9JLzg/CH0UQB+9jnxSb5ZzeiTdm9b8
z51dghTvBHPbqDG9+UijAY6WQe9nmZ04w6klQLF+4/aqsAJVFv9oQE8oav4n2uI8
EPued3BM5ppCO2JPz2U0X91kSI5JR5lJ/+DneGCDMSUIF+qSiLHRVjFJi1Xql7x7
Cj8weaB4Nv5s0y33l2LS2dJwVemOGUI8JR5Ise8OJOi0lJqE/BcOo5/sRtsHgz9x
79Jvjw0uqSyldJjI3Q+3zeSanUDD5CX1WdsPqok5T6C3cWu25R6deKngNDtaJSbz
KrOKkN4wXoLx3VTZXeT6bTPf99FMMIvMv/pB23kjk/yJF/4oUNiwd6sjvkm4Zh+D
8aI35hoeiYtUtb0ckni3x+ARXw9Y4WkLCjpoSPGgZxT/rCr9pPaly+xZHCh2c3f9
vd6E4H+loEfsUQUEm20QsACRD40X4vO6eVwlHCkFVyjuE+zsxDaGiHJEf0WusjRY
nNb9BhqpTj8ggKKCJZMFMn5ATPiEdHbnyK1qtcEzfOZiwg9rSISCa8GuJzKJRf4a
QETfBLtMF63xKWCPUZV9UylTpotHEWSmjjnG15b1I30Ju8TM7W2BBHgYnASTG7g2
niyaH1UPJx3S81oZmZO+5XhYGOtHRw+KWmoM0skABG3w1vi0lBQ2kZ9bUO84D3pZ
50OjhrEUV1LGH7/gLfK1rQOgJcLJTaHL5/hI6uhQsniTqCoCbvTRK1N9fTzOIlS9
Fjwu+t8qP2lTrmuYc15Ucrr/nafUsGf9ESwWtoVCCkZ7cGQ4Idcm23DMCIcjlLSG
f+hHYynxUF5drHOn4anOB8goebNijxjXHoz2kkG/fK7Uo5GlU0QCd7LI2iVXhKXk
bbSTXtNaPiHoqOb+nhFuFTszVONH+PgYlVZKEn0WySjrwyP2df84eayxRY0BurUh
X90be6R7g4s0+HUSsaWT4kEnuNWD+/0c1Ug9W1RfaBxt3zqpV+hgiKZ26Ly6EmyR
X6iPfQNnInvMCDgwsOc0LCKXtSidU/lLaRd5lw8LonSnvs4+5EAq2F9zxQDeOum/
c71elYHbHtMuxpaltOv3e11YviQglaWx2araN3L/ZdyOGvv27A8AAT29uFnW9ORy
qO5UEqpn3gy2o/ISZwmsWmDx1vdzNdQrFbFjI2em0yxxvZQOb19ElvDA1avsurgQ
9RJgJeJuOmFTlX5V/cns0ghJXdTZxwNPg6MRSsf053mhsqBDjKJ+EmZLQDVexdkM
oiKM8zXyjgXRIEWGOPvoHQEYoe/YAqjRUawDRVSfJHJTGUB0sJzteXT1loL8jnBN
+DUvxAEFkQAd9QZeKi4+f052Qa5l84TiqoOyXXy+iv2q60oke5Srnc00yqM28WT/
ciySxl9QGkGWcDzWnqaNObxXMcrIlTsdACiiKx94LeS8ztznREOH/nhuS4ljRQon
/Lti9n+82fWSfvI4NEvP4kU5sDkEtzmw3Q6SO4qn1AUu8cS2bVnljqhrf95FwO5H
kisfpvWT3adaIc5WA8VmWa2JswPxBuchyNv8ZdDzvR1m2E36eezIGBwPW3PzAP3r
wnpaTN0u7LKZsciaUlGCQbEqHBDGK1KQ1LCtI2cE+up5wWLk2PpkkJAsqIfVVWf9
NuoybZvnLG7y86arLUeTFVArGMSe+sxYcQkG1V83oWMpCo0hTDEWSUhKLCPzeL+R
EBDAgUju5JoU0M63dEdbYtdMord/kw8UxOQDJoVisQnKqy0KYSIiYtVuAHg2Xm+k
FjQugeXoNaT5i5/C09VEGDb/dcYMqb1bHf0Jm75CQz1QG2QtLZIJtkAeFO2aqf3U
qsc3hvB1B9C4Ia56OU+p5rP0BOTlaarvvmw/fMYeix/jgXTkwxH0DvZHDxnxNQ/i
glRD9p8Mm47bbS74QUF4GkpEae+uj/UUlCDZHoiIohJi5KSNSucjUIFb7zXajtfs
fTsnmooqZs69rFtdYgPrKEVAijLWVboJkwAcn6RY0fmg/R6WEpNB2DS83keFvHRU
AXt0zDkRme2kLt8mJxoVX/YsA3UZwaqlhAlQRTXfBpIcBXODpNhnoEzpfKseynIw
Zkf7S/UzqQ45gcptFGEbfGEVH3AytZyVfaR9NvR6BFaKX+cZjZeK02XyS3IxMAM8
4A/Kx6meuTChomjkotNQNTuxgU8G5o4DuW/HFg15/MkmYaduXqe2/xoSQ+R23koK
XOmW3E3MK/YCpTw6UGuoaJiOjFpd+MaHvJnzrVvoGE12aLGI2ioZyeCrovkXpOFh
xdxaEnXn8FEwlfPZiit8OTL2fXh6XO18SXDGDcD7bOjQIG3J2aCrCRyekW+Bvw2H
f+/GL2ZW3lCu0VX2b0+qP2SH38VRFnj+1nN3i0zDl3a7oTsSLYwxCMdUFKP+Y242
T5N/FFE/DW/V53So00SxzESZNasM3XbI7ej8AbNwdmNmxOVEKQ4joPO+SJrq3f8f
qM0bHQo+0R1Pdc8iHgpvr3bniZiaqxXx9z0VVSp1NqNDzhQKFNiF4WGn8B3rJBhQ
RKuj0kiu4zekdZ70+yfCfJ4lnQxIzDDXPymHa9P3ghzwwU8EDg8wrHeQ+twV+2YL
SZALQVc3L56IsX2tOcC4qYxWC10TqyVdTM4RK+H8FBkqfGYBCtXpvz0rSVUh4XqL
ROyu1EAcLo2LsoBEizq7xerdlg98zJulGkaAzdCcFH1hQY1ku1Ad+sfmBH9aQsNJ
NF63FSQzqdfpWt7XRVVWIUAIcHeGspzsck1fGxc7/kR8H2LxI80xg1j7X2+on59f
puHtd9to7Yd8hsqQJclsudTqgg0o9n6wR9cxQdbxXvbrLaZanW1l3nODB7IYB3Mw
hiochuXY+mvkS34d999+tCW04Twyz5QZbjWDueLbERVFncYd+eJETqa2BS0zVgcG
wUK91bLwPLOLCDPLLIJQKJt41hlY+Y6Si/Gn0KrZmCBLBiF++O8BKi3Mdv5Dq6CZ
aIExrn4iWO0VW/1YGKuM7HAGJGQgQTSxckwC4VDoemuOybbqYUgPjHJIp5PYFMzn
U/NQs3vWYjK+26EiI1chMgJcoXLonT0dBXZfZF4sF1Osj2aIn458wu9c7Ru4ar5C
GxXwehdz9ydywpzQGuX1mIa1tTLrcfdn+iqmDl2h3BfcDK2T/tLHk5t03EfQxiLI
bSPagiaVagJawEL6PScCwDC0wI1hGrtxXcghHpGLlCPhsvZO9blxobhjAUvDh9qR
4KUmZ3ZRyho9Pj9ZQ+C4xRf+UkoIP645Thm38CIWGppRjJiDZzxVxSKOpMLSFjYh
3typNofRtdeonMzXYAnUzmi9BQKpX09VQV68NRvdRqww72c3vC9+iE+8smcltu09
lHTjQrUmxjlROeKAG529kbZVExzWIceT/DZfOG6IMdklsBr+ZBXKm6zHE6cfWly0
xvP8dhKjjya7I60DVbaK9Hg2i7xt0hJx5b8QD1f0qT5xdfRU3ZXtx2d/BVEO9AqM
WbY+62IIbwXDrBz3mGPkg0Rc+NIH5oCKg65HE37ces9bqMmYsxCwDuRUmIufaYCj
DdjF/rBz3b2Z0dwohpSe482i9VzdMoRsbfxbi2WyjtGY/5zmY9BTnZZZ/YIn31xD
1bTxJsOjIHFJrrZqem5Gd2rRWByxOxdT5DXIsZ2+4jGQUG3VJip0fn6EWMe0XYfR
OVyerGvWXPZUB+D3C+IQJDIVV91RoOnkV28p/tkjKjZrqwgdyII4L3RmKQB2lUfX
8dPkn4WStP3Z/wvA0lUK+kUH+z5Yx7pQ3627rOlgCEMmyzotNEdaNf14Mwjy/twR
5PqAoRp86pdJaY07j3QU+varFKiibs/Dk5UMXgqDUGfHNj260+4XlfyED+4yLjzS
ws5V9+ibGyUme6yRGhxpR0KKnhqFKitZH2qt8UBZt0ptPC9uNJIk7czs4lb97/Oe
t1c2py79gVtTNruj3rWSj0GqvY8+zbGAxoPSz6YUYeknSjIccRdgigF4Mvr5I6ad
BN+alTwlpXJmwvX78/Mw3HqiR1yYeobgijgY03W2WXS+CljcpmN3CWFhKs0HNyQm
tfV43/RKcnKrJWUqL20XeCLUubTqEJq1J7ix+NEiKk+CPgUHebn5LCelNbOSjg6a
cYVs7ycOQ1H+S7SLP5fr7pY9y5f/+dlzD6PdiFE5N0c//V36d6FcKBAvO8NnWnS7
9OR+4dMjdsxz1EpDlYx+DlCOSyfNZhCNUXU4wt5vMnQuR8dQo8XTqesgVVP8hXPK
uFDXbU4Jf7PncSs3ztepQBR3f/zeC72qrOuHZ9b2aIEDMPt4RBFQNeDgB4yOAvD7
FEhKbGXpOoQXeC9XHG4KzO7WGSXtxt9l7/UWNYNCWV7FEHf9FuSizwagW9hVJfba
n5pJmcwZWZQ8EoQhLm/slJIyddGH9H7N83MtISid/K/tZgn3qVeMtZnZt1+xVLaL
IFHgLKh91hox+b+AteNtLvJDBJ9sm7Tv7v2+mUiawyixqljS3mKmOrUCDfRxzWOM
dcB49Vt4XQAuX1rWWXxHWSbwr2PXwYa6ejpX1uPLYhUykNK5muXz64/h4Fk4s0bD
3EDy3uNaItQxWozXtHhv3EUbjEX8aVXIJ+PS0AtUypGXP2ppBQJPV4egbbBK+ygW
TZOnknO+SUdnbKuB/LgeVJumVyR7b/5RiFLnIGcfZPAAa+adc0Zi8NRBPmCu2H8t
wwwGP9NlpVQI9LAdf8r48BIIjvWAsvwFNVxvRDR6GF2Rrzvuig6J3SX6iXs0Pt1z
VAz8xWAWYs0tnuicIUU1i0Ya+Fi81bVw6FIvWXLeJJxm4J4y3ChtUoJZrOaneY5p
ohSXCShbq8+xuVQ1XXHPLlqwGA0h8TfPYovphjEkNO6cW3dimf+CiToSUJArEPZa
1Sghyw04f2xgqFlDPhwKUxclZJifUol13qUzixjoM5KbDw+7zCCK+m4Pso9Xhbdt
rPKgjImK/bAZy3kZwHZtXYgaaHphfdzxFr1UMffCxDjjdpTF1sHLrEOTTy1TovdQ
rICN5nf1YG6n7sBtGsueDWncSc+pAhh69KTrP5EoryO2FL/ixWhjmFVsRJQJ1yLs
W2PjWiAoc30y9lxOaxuKI7WEVxfKcENdHpEl8FFjUAhA0Gi5knZr/tt95of83Q/P
bAx49oPLW/4RfB/xF3oOhIB5kg7lw8eMA3asASGA8vfPz31oOGZOQozvS4kPeo0m
BoDKxMaxjyKl6om4fCni0Ecklb5u+W7E4osSi1GuKGoXMl+GRs0+c8cfOZg82OjQ
Z+Jte7CKyf/lo4UFQqDyRbRmDzt9VjZMdh5qrHDm0xj9hcl2OkqXhmCOGIaOxMFV
ckCgsNQrAQ4MGSd3cDpvtIxC1U8WFkZrmibZ1DdM4ZrYsGAYlitGClQSpjJBOLZb
u+1mi2odUaqD0LtwRYtDFwpwkaTnMEfCGtJzIcb1L71ri4fr9tyvAt/vMBhxJUVD
r5dK5Tm1G/IJtkFwzJPVRQFDcs7tFi/xnEVnkqPrXGizBUk1ygCUpIE1mYHGy0Jn
fePjFsHvp1wHXfZqSNyXJ5nIPHutSo4vtkCDza480TB2es0+q7D1tmUGi1wikXxv
V7Dv7sTpjpIlY2edn3ozI3N23A/fbmSeM5HzpP+lnV7A2NeqglHKk5bMKacrKNIN
DJRp6mwPhA0NBT5DEsgF2Q3RZkZLgAZomdE2t5ba7Qe30mnBN1Xc7UeWOKal6g/f
YNjmrvMEk4XhVOabPPqdPnpgEoiBTM0q6L31O9SQ95L0bDTeH2aERPl6+2UpG4EB
rMatF+8hFXZTUuZZUAIipebfhS/6jeTJw8H9Ps2vaYeyPM1a5GosZuvi5A+qi3aE
Rm1CvE+DLxNphHdwmDDMdJRwfnk20wXcG5ACpCIU+Eya+/IFEVihQDNtfUf9jWcz
b9lKvzul0Xe3qdio7rHmCyRAaSwh2qYjyMUB5Lbe4l/fKLPOuiSO4M7Hk8FP/8s6
lUNPh2Zgnz1yK63yPz8HlxPYOF4jbTynwls4dMmlyKbJZmGtvz6a4OqfrCNO8zWr
eOcU8HzsoePOp9Ds1ef/wj0uBgnvI1oAvPTS2UDDbdtrA0TWn17zzHBICaswi6WU
hdzPoK4iPipIzbCAHY7yDoZL7VyeQc6OKdMaBWdnmjzB/Gpjcl+LOLa9HPr5flL6
ZvlnpRtJlysBc9aW5r+Okxm5MkyFdCPcQNYOUe36dvfKdJAJnjKQ61ZfrWwlbowd
lj6F18GEquMjhE8DpM+Hhlxsk4o3I1pKPy1uio/hNpxRIv0kGrAmMS0mPCQwyLvb
WSl5nQzF8aKpTnlCUulTAFsX8hYkWX6nupvZNNN8eE2+n6ZIu9AfVrOPDT91t4Ki
smbmd6gQSvgWL87vzXSiyc55SmX0BMsJeXh/LCRmIfkwAzY6FxiH/dPFlP3yRWHa
TjjTxfkbYKDlGxLnuR48ENqoiwyf8bsq8R+PDHotlydiDO2yfYBSr1lMGrSYA47R
lZgVpRKK2PbvJ0GWYM11ogwF4ahZp2VjouOND6EWEbmvaE0fchaz/18YqBh3YCGe
IB2QBwnHApNt8GKJBncY3wrRex7s4SCbGZp/II2q4HFWkYCmZFeDYube07iGVNz2
k8QJcxcxPyMYjai3z6pv/pyldMS/AtIT01g5DRAgpOC/rAXQAZ++I4Pek7SF+5o5
g7G+5KQkfFRET+xw03/hwtajA0sZUCybq+PxnFtDh2ymJKI7tSVAuE/W0/xDhZmt
mPJ18mJeQktowzI/Fx/J9XDNHgosxlj0oNwjqwufkPhgAEnWDihL0O+xnadlrIAV
3t/NiUm72NAwdytsCneER/uVh3X6By64/VNZsVJ2egwflxRJm0d6tvhEGlsSfeRe
PGccb4PsZ46TJDKNJTHV+oVz4DgMFe9LQOtVGRuMlGfsCmRuLR6pRC4NVHmXarKm
FQY4MNolYH25aHkr1jstp5m+8QTFS6Kji7fte/Ritn4tFHH18Rt1SBuaFzYEjl6F
P7yYQ6FfPXvx+zYHypwDrS9CXXh4nopTHPO6U19+bLf+ngWVzWeewGXNY1AjM9NK
HyjAGIvaycg4Xxv60I/1Ag9xpSH+QEmVYn9Pl7OSJwI+pcHcoD34jhilzjyf2Qop
RUTj9top4IAH0GiFDRNrNVxPpcaqH4WRsFJtV7FO72TtvnBpmkjRWBKncjXS3+p7
U6O2oAHWR5bTEJW6NaOsKnMxwoeFF0iY9eybpPuMDiF84HX3jM6e5nJxBQF3faR5
98joS5COzQ6M3TOdJyW46pwyWynodeye7Xjo4qFv7o54W5Pe7OyI2VBneyRV5gpI
jzRSbFkGyPnq86mKtyDCmO0CNuwS6gJt7YokrKSJ50GOEDZFae2eyo32Sgke2WLM
ah3V/q0BxR5tDLcJvr4ed2t4V1bet1gCZZcU8UGgO1ysKscRpvpTOWmToC+oMZdl
hgSDkaMFmrKlZBMkRD55gTAl1Yf9M6eGbf9YBreEiNOQ93qjED8QaCHmuAJnlW9O
p1o2DbJrK0z9zJjLv74VR5LfMb5ouqZl8neZ1uZuv1zMx+40EZ0yj1M8L+vBNnPB
IVQjEh/naj+ybnuVv690z+YYJP29xO/JPMQn9iG+h+hv67NyVi4sBKelDRcQNg0Y
cGc6WapWlBgqG0UEM916GHxXqxKd+kEvDvtVBgaV3kDAq3RnXjDQ9JI3/DdwOHGW
GbW1BNYv3FofZ156spuPtQYdmrP7Ozw9j3RLcP4vyQHSBe6v9t0IdwOXGwftmhS0
VFSi5iA8s+ScbmLWnwFiTapxQYqiXfi7A+g3rqH5bk+9m8Ad6rCxL/nr0EJvsVEG
44K5lJHUe5QWLpeIffZ5YVC/wb3tS6iDrES+OKSRXMp6J1kFlUpdLs+e38cGqLNM
ec9a9IYHjvT+jmZsPKvRa6VNpCGEqjAtU0z+5VlI6ru+XkkjsplK5Ra+bRaAYfxk
LFbPCUxukt7tz1sV6TxCgIYRS9laDO8FGJyhEiSlYzoeEorQMdl6rYvGTpiTTpoT
jn4NYmxCciRePe0dIuwTi58ltJuqTvknSiFnOFVurYUW5KRr5H0jvQSWbdKDNCAv
RYdDBSZnkDxr7TunsOxaEIYCVOWohFsbrhnlhoGE+W6fQoRMpQ/pF7HvLPOpD4CF
9ukUzm9SGRfaxnJbhNfGbRkO0bLHeaZQBbu8gq/9xWaEMJ3UFgzzh4slzXmm0eks
hpOcLQQm4y3/GTPd3HxpDFjBs9hqXvd+0HKqAj+b+TIQAIt7QqEM8cdDCo5n6vW1
ptJ5R0C9l/0Cvw9dX9Hv4/N/hgkzhT9ckvHZsz1krgnlwkcwmyBrbHxsnGuNCdRc
4U+RH7ACzDXJ6DRvIQE5eCvLZK6/ctnEdBOkvVodA3YmAOh9sgpcnuxZSbFvwtbA
sEG/1C258CXHLXRs28vD1O4EI+IjJNKsJV7JaRhe60K1spLijatn5FJvt8C5Cfv3
rTIGq82VLBwJSTvcinFqogFKg03VWjq3HBZ/jtE36TQ36xl5VSEQjWN0F2Jg9KLM
0RqJ/yFzgSLTVFf67R6JO0pcPiVbJvOVDfAklKZWcw88XBW1aHfIA3QJs2OeFoPy
FTT+jACyK4EIrn9Xrql1GYjEYsNtyZATs4bpdbRmWu4VuuTVVc7veBbUcCh8E8XO
fQq2UNxXDY6T6Pasqm5Cj+Ubh6xSHeFzIEoBBw+SUhrSLMAHT8ozWVI3K3LthmiR
+jnyXUXCC3ORtJ0Gnz7btqQ0WyGFInwdgMoDIUsJytPM2lNprqoFAgo9wvvi6nKI
o5CP9oE+/VCmrvXudV4h3RTOx0D0yUCVb5eSR2WzG68PfkH2Mo3pQelgP2DyiEUR
FxsamSEoBmMDxu/oVj8XNDmAXhenOMdhn8qGR6BUZJ0MeEeWwSVmFdLvMcigqJsf
kav0wjaseeUOM4GK/ZHPMtOYoLPWYA2r+fzT6TuYcmt5LqXbuGnIIgbqgSNU3kNI
BJNjgVnFJQ14Lip9blZPdkZbaXYrLPHLdNFP0SH6I8FQK9iLVUOFcnLHtml8BZ55
bBWoKWWemVAEw6RUv5C6pvP//x9Iduptzx3udMe/AQEVxUx/rfCe/5kaC4+5/047
QLtaSY9OELp/rs/dBhCLVWybpEMC6rkZwtlp3Jfrd1b7Uq1xtl2DR9PUtL+EWnOs
hRX4L098d3RqG96T7pocYuklpCyWjH842etJO8iHQ/rLMZG+EgF1YXa2/DTCBfDg
SJ2VmudS46cFgUE05HmSgKmjpy+K2WrkJ0oS95hCbC3JShYZ1rwX6dxja8M444p1
G+hvw7LUb4Mkr0qQqwy94y12e+LRNnqfessfImBoob/dz0S7P+xQminZQMSCE1A0
Ayi+mT3AVf4pc9ecPgepbp2PjnV06QfAbioHLL8LHUoNbW61x2Sja4fGYusJTNYt
Rk6QQ5v99Si3GIfKwUy67dHJLmN8jX+mZDr6AC9GPOVF5t8AIxnB8n+EvUh5WvbI
iSKfPTWJr4RPdkOvaO0knWL5/eGSTzKCxZeu/iOxlOpaUEv+p3yHIhrgYvzsD4db
N67DV1WMiIQ22C5HJkygXvGCgI3XWuafESC+hDlKCMQBsyBOMlul57Kka1XLPCBL
VOa9rK5GGdURwmYiF5ffIj2/nXv3bky0fBJqI9+9XL/GFIRsxk/MkD1W/fh9tSV4
Jz+V+5oX0ehnxIbvc5U8mnRR8sG32sQUajUR7FAUjREDldRR29prOVJjLx/y5dJM
CgTw3t5v5gMGkPZqV2w3RxY94tUUUZi6qk9UJSyfrbwDUERZE9kb5jkyLND1Ql37
LRkCxMIN2JAomEReX5I14GZbxyyzEE7h+nOP/1wpNwPgPMbwyfxWhXEJ2BciBvCP
Icyel2BhFS85jKV0CAv5Ik5VkU20odV1SUnVZsLrof/WJrX7sNSI9H9VJPzQLLet
PVNVN1UmwINJuyqm5wcAI6EEukKafMBHHo5K/GugS6QTgfhLt+u46VmlCinPDmOV
AZHdpQEUxP2H0BUHBBmOFQjD2Yl+KTemKjBmY8CW9RRRfcd6fM4IeFIGrSnKWX7b
c0nR9dt+DHrSplmn3Qlyob0ei85UepZteNgnvmHOooUlu3Zo6QKVpanonEP9RggQ
wcnV6T7niFV/GF4EyujtpVdEXIr9H03Z7gwHGsoye2yGvsGqK+JI36c+SmkpOIoZ
IIrIb3ldSRSUN8gZJ7rhZ5wuVicNJD8RskH131EkPvUnIuNckh/DBnR6voaqJVIt
tEpuXfuHFlBtOqRAq+FLonNUMaCeYLZH6DjaSzH1mp20qyM5KBkX4FhBsKaqvYYD
BYV3eyTVWhSYqvxMLhnkS1mW6O11gDm/4S96vgjgqn4D6waMOuQ/T8pNdlWOxrMQ
pGLXrBJ9nLfJv+HCnmYecrvX6Se0m19vPlhVvrVi1B6AtCUZG/V8cXBARa8IdvYm
S9TgqfK86pden6xd1KiR2Xojvz3W/6qGOxxFRushuRN+TFbFcPRebHhgMc2BpQCK
YqSnUL3kfUWPR5x/tlEdUNvFng0cmRXxhFI4NcDbFpOlD59koUTFhbQK/3jdI88A
P5DHe+d6YdjqrDa8Tdh79Re5cUmC1Xt8OdW2cJ7P+IBtS5qIvX6vWvganjBtjDN7
Y0ZZDtzbD4Q0HaKSPhMoDar7gFKyrs11DJ5GWRUnMHl888TpGPTPDRlEOWtB1nJg
cHIQJegf0dl1FlWnw9qubJf1do7XmpvS9TKJ0pEXshq9IoxWUhK5jpojRkbf7NXS
UgQbf/fommPSpOspL05T3clcF4j3cdB0WmbE5zXTScVeKA1jidVjiHVI6HEMFMDs
jVUDBIZ/UM619jVJHTTx9Ln7ylk15pCW7y3YgM3qDJaM79kbLZOAnoDaTvxwdKf+
FI7AkdvAqgz5lOGEoXUPu9ST5t+PO0/fzyLbtatrQYToAvOtbJUaZIgnq09hvtMS
eOVsHuktUSMdu0snHivcz/dh3xb/lvxFnUYkn33hWN6tDneHImk7d88jPMYLQoI7
hJ7taYDAbdAqsK/dActDSXLY16rmXL55sTrKrk3/Vq1Ueca/oOL8aCXExMvMl296
cdYhbvd0RG/CjImTqzdSiMInI+SwgyMJYM6eeeI/L1Q7zYO2ma8Hdpnv6zE0Xqbl
exwHhvouKZo7NX3lw4/lk3giE29uNo3+oVJZpHF4Jn5ixvG5wCI7o3QOxNt2meEo
xrTTswg++b7XO563q4lgX2FpDBpTbjTRLjIDekJo9qnsitIYZHA0JznNie0kFZbg
+GrNngTjbJKjbue2965TfzuXsPx5gbB9HxScD61pLgSmA2aET3mOkxjOVb0b0ehF
lusjQrfi5K2ZcGDg29dMIFyfaIvaxZveuEVo37eUYKf2ux08JZvQCPrTL1dW1Vau
5TfChRXefYspwGy9Oj8cLHPyA3P7ckC3S2ASMCzY5XALaaCXqXS7if2uwxgG9F64
b/gnbTSyqZuYG6LBu+T+4YAzlfDpmmg+BopsqZJyvIsYLePcQE3W+IHVYBI3jjRT
rgFWktpD/QeQ6ElRScQlrReWOVncc+C7fLg17gFQ30ixIqA9TpbvbiVaOwr9cgM9
Jdo5kmZaKz8B1p/cekHAbo68GNrU7p+s42e/8Sp/yOeIHDdfJBdWEGSfxR0quMg7
o9ZNZ+AG8G9w+V9zGLxlx0DIJlgD1fEqI8SQvO7Ko34kGm8s1N2uM4+FSui8HMq4
d0TXZ89X6B6a9YgsKaRIodMd64zzlVG9PCHsKqbEjVS2edVfSglqlheNi6/q2ZT1
8TPfryZoWXHo8vyfydHKfmz77Ptlcvwa6RIy5lSZYmKAKvF1KPaI3FH6ClTFMRXg
gXG10S9R6irPZrDhoPIxIZM1JoeVJRin+WIBwgQbbdJLaocEacjRSgbK7eI9S9oO
YKO0Hqbdci3hs+85eacB13QhEATdj/thxur65HMu2Pw6qfs+4wHzoxNrpF1uPTYy
4XqVuzOh/F/8mzrXcGagMJG2Jeoeq+YqXx7QPwXYQ4A/2Q+P3jM7pHB4ZypbVuGR
ZZyTSTTh8FLYR7pACqV4IVvMc0YVO5fbHMXUx/zpVChhjGxASly1jphU+CL1ff4+
e89WhNyvIWuNQAs6aC9bZT1Y1MV5i3vBYk628rMYnZuuFBV/GNokVeH5sGCYLU7X
6a7vqkOSR3zwavzdKb6hV57txKunmC21qbn7MRF4bV2O6sFNLpFrLsLb5ZSesSes
7Q3r5zo7MrjAFRCsddtPgPY+koqfy9mfqq7e/cebXgrYYoVyUuxtucyK5xWuoF4M
i0Xz0mJkpdyBGjLFzVQfmDl3Np6jkJax6XcCETNuGIiushl4EH7ExlGJdo/nXQ9l
xttSqDl89k6GcwefhSIf0TM4uURcYw3BHsuyWJ1ImoGKtlBFMzJBIjGBMRDFwyCk
uNso/GRKrbjvF9VhqUB99VeZkjStW5ab9N0QH80IPKv2p28IweSjzgfmbeNdfxgB
8kB8hyl8UsXrABmtl1ipNHaSe9hnOAplVDb3/SPpWf0bLu/LdiFQUU3G1RXczp+B
91MCZrJBD0E+MA5kmhfIzUVAGkELT0YIT46jns6xHr+8aRmT4lmYKT8BYyNwzr6x
COJTVOlWfd0YP4mHfXfPRFwgaqesGbUCenGeitCqpFifR7gJlczVuoPPulum4rCw
OvhzDbIa58LCwxkjvZe0g3PCY+1xzE2KU4A8PACQUX8ic//mq9XlolhKpXulDubz
trMKj/+XEAPnlPYUaViDlAXsttW/WrxD+SYrD2EGnhgSiJe58Tl4XW7CEN9jSt9I
XwIPnlgHDnLi90/lIyijWjR/Tsyqfoh2ieqTy0Sno2pWHSfXfn5ol+sLkzCNBMnx
xC2f6lFiEFOm6YypTl+7JKI04p540orZ/jChZai3Umyo8LiFTntSQlMkY37MUK2b
jHTxtNcKHXHigVC0wPdboMDcMCqOc8PoHpHf+GgBUMvv/r9FaQFhGUoisunrUUEF
cB136mVsjsrP074tOsS/svOT8Rmw37fZ9UUwei4TUv8jRAUzRO4QuyCfPZDI8cAm
sW/NgSdqRwZ+OTV2U0+2xotnmtrMd8hz7HDSvc0meA1Dah5cyFeowCqc/gZq4Q1o
PJGvzoaIlT2B7P6GVVyOTy3CVUvnOsE/JCO0dJQ32CYC7MGrakszdMGmu47t5OLF
E95E7hYjpn7c5gGaulPRqejSLp1D2+DBHYMy6tZ8yVg+sK7j4/FThfQ6hRhPw5bj
OMSaNzoofulqOCDBAu3X60BRf8Fg8bkfSPfmWj9ylejDr7847D5/HM6T+uuTaJGr
sJWrkHlYHYyvMK8/wvbyfyqMidpYxQUpONZIpcxGAxlMpYPDCYvXpBF6TbjS6o/f
euJ+IOUuMPNgU7vkt7jEIXjMekNbbJ+gOc4JqyJ8Qh3TR/+P5TdSVzDZ5gsb1tcy
g5aI6k7S11TFotFKkB0sL3fqx3LsAmt+oukNzApJWu0739cvFX5k20Xfy6Y/RrlJ
dQsLgfXu1O9Z5JXLDK5zu422A9oA1qb5rEBYxoMA/ntAeMj/FxPG1D3U1tm1h5P+
sv8Bw1v80wdN72rlklFeNqoO9xoqn+iAZikYAR1VI8p3xsHx9hMiVPsEy9gPW5Ir
4OTtJsq+XIjHE68zCGeM0aKKaehg5OMSjRQWncv+DdSm2mDM76vjldjczOf6AgaF
mkpjL6J2CojH17xpOXErP9Jb0eyTYzlCjjUtT8+0b+KzUyaiky/WPAxeF++nHITT
mKClIXFIGulz70Lg/gRW6UptOzTLiUn1KR5b1nEN+x4TZxgWlEkzxuTkrvOqSMv1
2A2HmVeMA1jHnfpLfDBtooYS6rTUkFkgLjNnS7xUrN/nUcnlAeXl9jsEqIRyL3b6
HpxPplj/XgDApXuaKdM5QyzclRRW8D6rxLPf/kxkXvY3eA7FTWB3lEmAmFyU4lni
kxTj6jb/cBRfeTpTWYRC5B9g6pmW0sfJbc59zVYTtU/TcojlrnZk7Gr1NbxGJm+9
AwuC8r7AsWJUGpvffdnX3xLSdzxtchWlcdVRWcoshgZIc9Dy+dkDxJoyomoxjOJw
jC1C3ybu9YWH+/mCkUNKl2LdX8h4x1axFWXOIIMAg5UAjoN4KQAWsB0mzEQp75QU
UNsbXgg53yEqWg1ru1GmBgz8zpmVtKQqLBMz6TxVJHaGPykWSrKpbfEEppyxUQih
vLQY6Sf9POHYbpwQ6rH+j8eBl02aNW6P/sZHD5ed36V6RsyYy7igsNVTpCOwpbZK
IdPpdmO3ZCjKf0xmx0KrMLctDY4gKaBtGHnwcji7rOypLHALSyEQBBYZQKKbB5gX
kIZhtvFGvneGds2xkTFIr3zYLECHT2JqjHPEzvyKsXHCHbXvqQZytf8QcZjVo9EA
dy1RxKrCT/4cR6/IxPHzLk4m75roGmUKT8Nihhjnfldl5rfpfzCwtnsDkr6AlJdd
W1wnLMzrPM+hYVYuWJLYHisQYkakVYAcoaiEUsEUKawTaOJTulJm3BXVaUaN8vcZ
UKUHO93EMZLLGKLOGUJEfsUFhs1yYO9GYewKQG8HuwQnjqh8SjrGckQ8/DgTL/La
CSr3DBPCD0MnMuQC5vIBm22qcGIS8GADqEKrqdV8uIn6+M/7I/tCfBxNz3gIsL1B
gWcFHTW+eYT+NMgdj2nTyGaVuXDwK7z8t2pxzvBATYfKBbK/5XHRuehGrTwYZxxK
2PS3d7EG6TyDpkP0I6I0iRg3dhXWG+O8moWiuxSEaVX8//IQB/exttwnyP3rpXTJ
mWqIgmP5g7SC69O5h2/oDzH72Uy8u4P0fQeXZWKXcF980dMvWKAKY9uS1Amax/RV
9TgfTg1oRaXhaC9FS4ZweUCZCKStU+RG6/0+w7U3Pm3xVkIFqHHBduaWXd0RhhgW
EMz5G5emHTvTX1caTsM+x3njPRj0NKiH6z3JxUHdv8MNWx2yfoZpwLXX8NwUcNTL
/nNJ8l9bNam/vlnZW4DbuMW84pE8P6ScYPp8S3QR43IDZxj+WDuaMNkFaCFWAJGq
mBtaoplW/X85AJ9XPiGGXDIQR1hmlaDfLcPebTMt4cPJ39D1BSKPAXFr++lVGJcm
ElATIqECfw6S/Cyasg2Yo/W//r1mRAsdW1qMugEbh0RZKTjQLXyrtW997FJTPPMo
h44zK+fvLd39SBdH0hBjpxf+yCD/Gq+aE7otTK5fJdqyeWDOeRaB5ubIAaVXrn4N
Da2sz6nHAGoEWQmGupVsHNV5JH+Qp0gp5DKgXCYopyaw1J+oNjSOFx0QNJW0u3jk
bW1KHewiJpkj/7an0ejtXwG9gIkoERvYMk2bgbliSptM+zFD83LYJCI4mWh3Gbs4
1EL0ekIrteT7q88nHPtrCNUzF0Y0lZl8lXf1htiwwpgIs+npaY6RYCWKugxJOStF
64LecVnCXHWFtw29wK+dgOPqkwzbC+a590Yh17CQ9JDrobPl4j5x0Q48fnHz3PbN
BzJnaBPZyAEPmilifEZoARqQw8DN1w96BIZ9cORyGrr6hoYbjFnFxOmgzmS0RXTm
B7hDE24m4XJp9FgJ7ra04JlQq9B7QNmsIHSKIlM3rBva9Ol+wKz6YNG3PqLriLa3
Fm021TBcF7/PX7GAhzXPqAkbZPHMGohFufJR62iTz+jQ8QIW+FMCmGYcPyrkZwJl
zbLOYFwvRhD65p5YcUdKbWBrI96n9sRMznPQHOEFEDMmbrJ/Sxmzo4OrhJHhYBCo
nSY92RXD2oph1fLYbaqUc0zOoxTrTUzAIJpGdd8D5pR5HO9AfIYEtpcnu1eYH62p
3CnXkL4b51523QxWVaDAXPrbhpk9uWt7AHwKH6TactRvtXASmAvuX1kTaK2vJNrE
uqpbG4i2RQnegP/neE3l08uXUyH1PqSR80DDC4En49H7YtWg/BFxdxOM+85c2qCc
LHL3B40np9Jsdph30+yOGElMf/gR3GeazPJDfVPvzSwEy+R3uFKtLTqZWlLO+YoW
88sDXLZhwVWrKkt4Q9JQeSqpCK01EW/994jfAtA3iSYdmbwISJRx4h/1B7NVC/xB
z9E/5vb1D4yoTOdDHfG7JgR+/EN3iyeWVRNvaRhXXbYIDiz4pjRLjFwizxFBjtjv
8thxehl1mSkKeXc2dm4xigDc99R7shZmRtzaejMJmo54k/p6wVvZ4o6D4cmiXm48
Pd/adZzm0iOdac6UjxjfU6VN5yVyrVBKMAT2+sNpT7W81TLedPHSfbzGyK+Xwvty
T9wgLj5FB5YobaWzVLTCK6w5rQluVG+HpTTfHqyDIejolfmsI071x3JUbTeNMjEV
U0JAMAD7LPHZA62UNuYuhoatb1YCh25pLhlDZz2MEVpMfY0AbYL8MQNeh/wVNyyX
FAKP87wa5ChSMMSqxuSqsXp2aHUbCWoVIFgsVZQqMebYP8TLGxKxXzdjOJWBgYdx
e07reuTpqGtj0jQkmavc/U/8UCb3V+7KdA595zjDdOa0aVkGElOw5dBgN3Ue5/Mj
zypo8VYVmyEUznilvGTTL5ixK2fsxI3DicVb8PPj72NgBJmwKsPauwXuuR4vcUg+
LXoFQpApv4dkm3EVTZ6HuTiDr4IOvNLsyMhKZ2xOjUThvf/7aNzhwvoTsXK+d1cf
GGJNSKd62BrgkufLFZsTgZ4F5ME3EitkLaNqzfdGAsXKWGWMaDYR0Zo41R76DFoV
hK4MnOs0DF2ruj96VJrzF+qEpLwN6lqDsHpXGo1lUGhKfrylVFQ1Skil1rsuiDLJ
pCD43Xi9SC9oKWvQqssgi3rsB+hgNmb3JLUzsuhTGVtoS2kVV3A9F1TBioiRzeEc
XCIP/BL7nzjO5GYbwjcDmteXRJCaEfyy8ShfGA11isqmo/dQhrJ4d7SftCcdHSHq
IFDgtC9nm1sWEOc5C5oXMvgcCoHsDD72PyqE6w6sWBhRqisC2V4ch3O7HneQcAmg
MU11ZJ2MxFj3DqAigDcpKiiEPAJwJSgfF6KiVzl0n8hWhD6TgxguEraTfauqVXsF
7um/ikv3IAdT8Ub2HWVxafhGQwc1jlMc0D1roAE3wLVtg8Zwlb8nGuvqMlD2hmzl
B+GDLmsTvK78HQOa7jXLCXJyw/PumsjMiLWTONUVJbZow5HfBLRWUSYbdTrClyaH
hE7TDxwJUKcgqKsZCsjKIl8Y0KV6GhsTtrHa1SDuLe3NlssF4sk5sjIXCczThJ3O
yo5A2t9qbC1u9cJc8Z1exmov33p4tGqBCh8p/qV9R9gN8ThpOoqtiYC4Lqh/5i4P
5rt4KAwmvW5w2J9JMm6QNrdj5NZt64x3bLCFCxfBjEgynsGku++IKubyNO8ijgDF
Rj2trmO8FvEVi8JasNDWEgaUlP3GVkpasc1uzWKJrKqHAltiuIKPApsnO6geFDz3
efb7ucBqruJPGug3G5EzROHmKACFHVS5A39jwdoZMZnoj7Mw37lcFDmYx12Zkst7
W2I+/CWpTb8ps2oHwIAGlj71nkWCLZJDmIF/IQ3CpSL83zExlvNtTIGzNDAt7E0K
JIc2Q8FLijSh5hT92ohyh7lWN0/zUZC5Qi8bMl3PZ2aLw8ikFYWfvnKxbFJbcKc/
/1hUX0zBiCHs1uKOOvAR5ZcGwl1h+nj3KkILo5XF2kD4lWwz0otMSYciwly/55bG
vU/bp7ICyoIBGQjqKAlVetuo8+YEBdnX8B/fCxdgIG3z2eW2F8DeoR5xkUMW+GoC
9scJ/Ly+viFHcDZLIrlFTHR16S+Kz6I70AFGp4qXi5KunVR4S9zWZPnl2C3OOrnd
V9k/82bdyvzw7muKsvijfc3yePqeJkGIOx9YUdLdWOKStWoGg7kIAHRYI/rje9+G
XaGaRBYrrh343BrrPSvRjoKWkBIHRpjpVCaXtcyo8pkzL7oiL4ZSnRXr9FrMV35d
joEnGBnlvlM3ali/qn9mGVYFht1pO6LQYREF4hdcuqLHszbggO+EB0KSwKYS+VUH
sYBDS7od0dTOTy85PS1uq8Zxh83mcpnaVGJpDlGUnPtjWW40anWYwKXfmvvG9MzH
g+FipCx32JfPD3HAlbhgpXFMEryytkqPsRdkVRS/jY78FJBWAF01IOr/YdqP8Ix5
99loc9z8QO+9JY1Qfmlv/pKW0cG/knVDHb05TitDaObEAK6WyCg5xs6g1zL1UOIu
NADHaoEa3Ce99p7UvDv0X3Hg93UaKbHyIiEdtdex1RCaZgJ+czYabQlPEgVvJLeF
SaYuTrfnK8jzi18cThQUslpfCadGMeLBEcksBTk8+/FfrcFnNZosSXTyKv+prD8g
ioRMT1WC8etP3f79Xz/uU2h/52GsQs147flQZAVu5bDWpEDMf1ld/3bsAyJ0I4ZC
vVwPN90gr3bFzufbjxaTntJA+RdHRrrVdbmJDbqUXiB9BIJdHGW6UPU1YD8kt55K
QBj/D7sA575h54sIDcOcxwxlrQdf9cGmwO+hSzteZQEEQue0J0TRHuyb9w9VN8iL
KHy2KlIkzvMoQBLkg4ppt2+D9iSt5WdCDliLqKykaOendwaXJiFp8RpEgZxKs2Ny
k3vCrwA6s/xsSnwNqByL9jqIrRB3DlAwfl3uHGA/5x5PjhOiNLcgMUyPBqGbA1rX
QhL5tN2ull5shmXc8jZqqeOKIji02BYi71W4dwr6+n2lW5IwcNGECc5dzLhm/Cbv
foppNL8WP0/C4jcKFu/PL6rFMobAIhhPWiVmnRMSzVwmIvQRm9D7LO4DFnojrxNF
pVDylQL6ZcpqkOFNACdyqqml/U+YNLJpcF3bsM0RT+nylxNdfIF4gQAnIjfrQBmg
Tg/Os3VTJxoDBg7bnj2vONglmXrWvUmUwK4CrxQs/kop9OiT8sUbWHI0GGPA5KDE
nwFV+b9bKi86tWZIhIqKy/SBVWGoaV82n0Jr63XE5uz3qIAGtiI3Hd10nI8zUb/U
wRVJHkQVFG8U/HmHTAh9ajmHMvdMMlQI/3soKLXpOMQ5iH7FhLlV58lZ3yInuqzn
swnzPbxIhmXprdvycJZ/p+paZjrR7Qa76JdpIlD1B1UkGqnloDRY5CC4Hj2tbeuy
qlB+GKJiXv41+2ZUQjmWxzejic2tf8keWsWlW5s1jR/ahAgWUL9csu6EiB4XtOK8
T8q6601SoQ/PbM/TOQYmYGc1t9VCP4a1KLQrXQlc9kIhaFtnkJDasg/uU+mkotu+
voaD2BoGlNdN+Jdb6yQ7Y5qjNt/YpyQO885Hh2CGpA1ubbnmOHD4+tcakUsb7EBY
QB7AmKaR1qLdFdhIypGIelxzq5KLqAg+oxVeu5BTLauiQZ/BCpaDy8ts9e0QRF32
9Qj9ImoarLJxcQPQiJahYA0otmAWnylqN6ayatC62SQqRsY5XKcpeS7VFUAhi098
jNQi123yWS6J1oAtEAcyKn2Z38lutSM2iHeCZgXoDhLeW4cLoh8rtLyHo+Fu6cM5
gh7uGT+xx4t9iCzRLDX/Sg4bFry8K5//VruvNi0049vQ2piMm1Uw7SEo/AcIcyU+
cqO17jrWXq+AthFml90ISJ63xnIn40lpQpbK2oQxUPxaXn0GkNK9/qVsiGt5ZhEx
I+tcbPU2Q5+WEV7rcXDQ4Z5KWXwym2n4BI4NwbKli0OjCMdVIP48F07WOXSWPXuf
GnWwdxG/Jk6NHSIKeTQkWKci8Quk2eo8MLnwK6J3xkHd+D4yGSz3r9k1muE/Dodf
XXuJCeKjENFJpN0hEaB+KCul2MKy7CWGHot6GWrgMYyc3fmzee7VjEWVgLn9zAq+
vNIZ97BdWN6wYjLkQjyhvyDcwrgPGPLzSvkJbsXdSVWAdQ4qIu61fzj83IOOXxyg
+j7Tfasc7lzg+1uotuLQQ45Q/jw56fC27+84s/xKxznih67gHaVyvdKwwbzKRUpk
a0PgoSuhnOUTIz4gPMZLPGG4FpMuo8TAENpxZ4f+oJlrWvrgOKsLR7Eg7LKP290t
Nh9Ci653ILD0kgda/u1nbFZvO5cBQQ/opZnZpRT2dQZkZCNIHMcID6SefJM+DubT
92yIirpeOBBM2pZUuo/q/9uzJfjaSz3VAldDJC8q1fR/LUzWkrFhyFIyWdPM6/d6
Mg7KFsmPSiLD0vvkx+JSnrfS6yFiVrsZMt5ROhNF72OXtUmKOQ4EzgN8ecZaCL26
h+utkglZCO2r4SxTc9hJLAtMXkuI6Aew4RcqGjRLP6qDp/XicOUkvOXT7vo8kcnJ
osJZ8X+uEYC2fViL+tPGwVdRRfAkmognlkXoSaKuqyNtk8EIPQDrv7mDu+UeI29u
qbct1Y1Pdwk08/v4BSiAM7KsE9g8zbbHXtqdLGFRGCsZ2wad5ipL3reytpCRZwhV
IzTx0ssda9ITG03ZmFEfQcK3ZNZFzDEn+vNYvWt1tLYhZ889kZhkGUl+zhp2dfW4
xCu/1kvGGAHW0hcAirAomLkhKyjeu3mrkJrFPvXG9xcnxGTPF6jDeqb7vFrF0jjq
uC/p2p0OnPSxZaAkBzxiVmRW+Ha67O3tfFcc22FCzkBSnAZk2M+zkyRV3Hi8G7p5
TZoT7xEfv30mL5g3vkiBHCinSfq7NjcIgP/yYibSUEfNkV89a3RCsqhdW59Anxxf
5DvWJa5cJGlEOSHcoPa5iW6jYFtVErPdDDuR7WCeimmGx09aNTck0iwBbr8iOC/J
ITJ3skOcdD2EFh/Q0Af2+JxINiOqT32asKXOBJvBk+/gF0h9E/e6ORJEBBcpdxPm
imUnhRnNxClb9Rf/0w0DzODCRj+A8wCKzXVkNfmFxdSzar5+vaAavAXG8QT0olx7
3B8MAVeyUSdl3xvBd3ocSdSHUNrmTaR93pwD4OnfYQUXZL8SNMOTK2KUVb5PQ6kp
WzRw9LBs+ksHJauHAa/RAScbSzbvJ4az1LH87RsxSnxSID3SfF1u2X83EzXhxhDs
YJ+VGJ/lk91/valeKFtSLws1r60LqfTVjlEOC/CWWoJ+l7DWhRWcbM9ZGLGPYVHq
pDjkcm0u4l2P+5SnVyBufpDJwTPUik3w+3ZEsVd7k4aqAjeCq26O+JSe/0To+JrY
V2MnAu8Q/G5YHlz9HnkwHs0XwiD9oR+jMkdaEV5UwzMzSXIf/A+DH7axT+j5kgCW
FSUWGE4V5alEbr9Kbi9SqLm9D4bfScirMm6rq4rgg8FmrMXJAfWobuhNeCBG25tb
RhZayYe9owO6WtoaBq21w+jek68oMhmOGOXu2AW8SMWnW3sJcq5zn9/62umpTXPt
/kaNg5d0nYPVxnseG1mGMsC7V+dBFHrYaoxrqiV0JQvdYvL3OdirAZbGKYZw+nKB
ouSYNnNOZfxLV6wwSrplIQM9Dj4cNPuK+fnxFUl6Kg3QBCbgJRnpfFRFmnGpGKKY
/G8waMhlrTuHu0ZPfK8RDQgJ8FfPaH91bj/QBolYitOCrIFayAU7Xs+t3bi+Y97U
0Uzn8+ITAtunWkY6cPkErCRrgHfcqHTMgf0leGLjXoRRXmh4GyBCSOMhfR74HF1g
cXdU4S94ITbbcIaHXZKoPorH6zzd5LsjqPgPiuN0ah6JTBADTLUqkp97e6+hU4k1
SVHcfBbKubOeQqeQt+pHtkFgH4LwkaI3QjmBix3v9PEypRSkTy9GazWvLojzrVSk
Ek3YRia+Nz7Do+2Fw7Mq1+tmwhcAYCXns2EoPva9hP4jQyqo9M1RguVJ/QDAxB74
lpo67PCeVPfOA06teK0QIn6YEqFL7i5Yvo8Tf7NC1aOKUuS4YrsciyZceFocHnOz
ag7K3nl5E7Uwe+NTkI8S0MMIq8QqqSGQKNuEvuFaXR0of8AWZQhmy11O0xd30fRR
hqkgY3tgnlVMB/PgWWUt+pyd2dThaheS7vA1j9qJacl1X0Tsd8FbLe1YW6w81dtO
Nc7U9aQ4QsSYWKqKGd2ckyQ7qnGneKee+MbUNj9AAT+EFgKV8/zPGd7hELaPagGW
vFOth67X9jDJLCgw1FGwtqnZvox58fO94BspLQm47G7W+XWTirpXyQNf2MNdIt2Q
RV6raiFd5Y/Gwx9xwRO1x0FiNJiBxkBlEyaTb3cpdEgk9P5qENnoEIdYZ7/JXz0r
IKZr9MQQp8U32HMgZCTzkKZiGtN5JUjn9jMJpaaal9GFkhlfAQHYGK+5Nm6ZdRqo
n/EQugyji/DCmb4s30M+Y/daCWNAkk8xZtHWT/YKGdiNh8wkIm/+lj8nJ4lUxgfz
G1F20DgOOiPgOZH9Oqamf55SGjXVbJopWk/Dh/caFbB7Xue2ofDeBvW1UFkLdM2S
f3E+BiwHgiDsCXdQXoBNvREZhb79UEJKNcTaucribevy7BxYE61DRL9hNLO8upkG
eGz3XTYPM4USZFz2q6cVOto1VOOYP6GSks09EkiBoPfVNfK4RqKwO2GoECsC/b2S
TlmutpfXiDdGJkAZ4yUo+fffgaJMDO+PW+IpDE3e3l6UttUBe6wXZzXZWge0Tubb
8ddHfQrX53uzKt7R0olL1pH4na5TkzHOOmuhcfTsn6fJGlS2eeHyBXam0uTKGLHg
Xi6qig9lp6RYGDoKRZa4qGzzURL2aGxwtVYF3pwAF3PNu9+yf0DQDAGz9I+hM+m/
BzTBNICx+Qpeg3Tn16lqX19lLK6XVQRSbqo+pqQDkk6IYHXtTYlzLQTUKq69yGzH
PNibP5/j21xggzL1j4Dfx1e9mSKY0Q1JhH+gXC4mLacmgWUoEJeKA25VRzwbgBK2
ZMffXRXJqxEHFaXYWO2a0euJx29rjKuEjkF64FjSGSS3mh3UpXxx+H5hrCQn3fHC
2Okw87sAc1B3pjW8WK34BIJeyVTpEyGE/J8C+J3ye8Xem0AFAa3IrzQUjJaiT/Kz
F5EKCHleFtittLUnh+eCxiudoib9guQl4vCy73lNwVc1YZbcvlF90IqzOhMcSUHE
pTa9FvuHqYDlllLoGxCSfTWmcNE/7T4CG1RkXcyu2yunMeEZ7PPHts5+hkHJ2BCJ
bZZOODQAPc3FIA9v3u+Xow/1eg005MNTVmY9KUDt9SPMjSu8E8gdNYbfYSIPURc0
L/mhn/5ttwOxpz+iCiQhbUS11EKH1roT0wPcS/t17cP4T6DjkauAkhqWzXz/3QI3
TJutfgR/e3MQ5RxXLYF3Yms5/6v6uCmddeoroD/MDoblhS57ZHjOpNQeEg49jk1u
Nj5C+OR1pqBGb59pBLtNUoMAVAs+YYeqhIcwa5SuH2Glc0K4DObPpvM0QljIT5Jx
vWTKj+pJMASK5k1PAGu4b6b5f7awBiO5uOZgyFXARc+4550GsxnJCLz3u8rKuxl1
dhCXmtpHrY6/4CC/NV7CuIWhgUdDSuDpSj4j+6CnHMVl+jVtirLuB2Nuy5QfbHCj
dLKhTVhqqa5KCmbGyCFnompqNmg4mumUWoDBNKQ1gwLb6faEjQ+CYmVVE5Hc//A7
6oAVHkn+YD5b0SRTdtKccL/3SlrG4kGioMi6xz//HGo3lVAxc2plou/Gwk27ab8N
OybUgVJMnbzkPnhykFLJDPgv4A4qyXcDcgupBUidWtIPBJtU9wSmw30+rzqhQzSi
yhXsfvlbOICRbZH7udXNmVTf4o50Fvg9DnPd2HjRnjFRIIluGtxJXY9Zvb5Rx7gT
CtqD4O6mTdSySLoT9xEzOcniz83wytL/Q12hdjJlz1vGiHfebUJbZG1OwA6H0+Zq
xAwvtjA0WZ7RCHqYxfmUjRgC0xVzJl6B+giZTy6s9LQXrr3bIx4uDjGM7N1Qwzr3
PCjQdctL67FyGH1DdlB3KwXp9cqZcbcF+E1ElxUWyQsSMBqw6lHbgCaDbx9lAEFi
nWhT9HkMrDqiYynKHTcbjQG2/lKPlXygZGWDXyfGOb730iwtxk8oxSS1KUoDftlw
wW/kKeeHCp6MAD9+qVuCAsl5c03JHr1oRStq/wgAFswlap30UAvHlY8OhargQcby
BWBCSa8dBUVjBIGPhgk6UUswWZjSgc4K2DF0jwXN1PWnESMl2H4rMZK1Ink8CsCe
2e3xQgasWvS38C1lQwwIs1AX2/ROZF6jdTBv93nAFlMHIUrsXovRkzXRDF5oXFoN
+CBUlbfaGSGSIFsQapdDyicGiI0wGQPTiF74GNu1TQIovmKIssUIhWDARBRoEY+4
dX16/e7w/uPa8qxAw2sEUI26vlFIa+WlQ4CTc7QIWWpNCAEwuVGRIh/cgGCxWUN9
K42LucSBhUNSrwbz5NSXpaT92c/GJB4MWcaiKWcGcqxqduE/4LjxWRdVvly5i+/p
dh77DKjBYeovqi6ApW/2HwIPHUB3jFl7a7MMCUfEuMGnOx9kLuTyNibjnIA+UYmT
Ud8Y/d2bbtOyRiyPDHyvWqRMEYtT89PhzmsXM/2nYl0OMhflbtltFuwIsD9PVUzk
q4RbSi9vdBFmzRxzBKm6Cl44EU75cTp5aMSa1N8yw6qeOvS+M5owdUmut45FjvcK
3fSsDv5o2LjsSX5KYlnTfoECIziGmMJ480etbLUMkGq5EUGKrsHidBfltLTMin86
aADc5ve72Wu4ZIu+QGhUKr/gA5e5NJcRYeUdVRPOQSfnIPQnV++yT/a1xcmh6yHP
y5fgULJ1JLVsUdPAbOtPWpCFHrG/Aqw0YtH+2nnjjW/MDdt5mqyE0hwZywpVCWKA
vFxH+PRtILLP0ig3KtMwIR6Kj7F4Ptu6OS87Pt9oDFLuNVfV+ZyOEb1KkAR/dbqe
+IiqaOXbAxvX7lmxUQmrwImn1aZdELH8+jNqZhWIt4LuCAVPSoKTGAlWfOQoqcED
I33OiUx+kULFuq+WRrjk8qRsJcM4r2ZuSXpM3wutVJTthF3Pab9vuiCPf6axB1rA
5RHQhijNqXpwZWsc2IDMBIf4Rh9rY3o3Zi2h3tn490F7w+Im6M7r+75fcav3uyUE
VKLc6FcavR7dZVy7vYSkgu7V1bhhSs2VNeVPmbdFOfeXlptrrjtISNI+9PMGMB9w
mSftGPzj5Hk3EDiOOMRlCXAC/rSL7DCPtlWbH0IyTXflkhNaPOAfi5V4CyUxdlZE
w4QsAwyuV+MJUoKcinGOkbk1pahqlCWUpEP6gxcGdtY1GC5CWKVilTNv2kAg0NJX
aNoFAbRx5XDV7j8+Pc5N1eXd4+OYO6QcIzUwWtN6V+6KIpzZ95/IMgrAvuGaeTs9
dAFh3XimVOQrTp4Sg8b4KsswoxbF2E1AoqGtMX0LD+hzwfkQ2rfMBbO8uJL+vQaG
oJ5aTOKT7JWQeBQMVqNRuyPQ6o02/5sM7Zi3k3n7ZJMNurdzCvrbRZuZljmF3cLY
jmNVYj58A9zwnRVamif1V6z2CpCa12InLNbyhAjt9jK7LaphwtL4KZQ8gM1QOQ1o
cFWo1bC9NXOcCzcFJm4KrUdGQ7831/6OOz3jJet/VK2QFrW6kyugTdZm3dTyvxEv
/A0bQw1SS1O361XWMxLeFvVCDNTnFdcEYg6+i9qsfO2hkTOORV0S5VfEm0JVwG2F
3UWeGcE1jSfUiu4PFSbREv2EfYuD4NPaqLSSyKzlazdmGgsEtHGHy76nNl83ieNS
mF1fanCZGHqA+yXbvTPqdDnQMSHhHXmNceoKAfyT+fSFP9m055JCMOB4b6RHcTNW
R2VoPOfb6qUs775k2OLsKTahHg5A2gi5oHBmSj5EDhK5bUJmUDPUoe9wVCojuzZg
NTqlwOz8K5ahjqzdPkJ54XfIAkVZHYspaGgIkhgwvl4DSFznks6L08TNTt+oC1HO
KWnmYOIF3av1PmLIubazIWVM8miYhhJuCp3MyzTVucwvu2Ag4xQ0q1NA0kEyynmQ
A8SkHM2WaV5FAT/g/8+RHIIxJb2ZL0Kllmhcx2HeZf4beaYB2+iFGPk500oaHVwV
P/4nHJjrfShnJx4jjEpbq0hiNgYFRX9UEZxSuQW5DwzUO49nmuyMCmSogWtLp9yZ
ToESir54Upo4d7hX9w3iAT/ioCx5j6KuR+NnLiyY17LVvDnp6cgJC4ZcMxNCktIp
qj5PUp98mpFYpEd9Ui1eeOWErEdqUziPLCzXl23NAEmFHS+HVL6cJPUvyud2Q+km
9o49LQGwpHP+YxK8LV98f9EuXwn9ywV7iRJR45VkfkD9H4yRzNZgCK9x2xqiY2P8
yoEDB3tqCgNjmbTl4yKk4MOcBJkAzC0rwIsk0WarIOtA0R+1Gxdsiw3FWf6s8ycx
q8VrZiNR09IhYS+0LOzDMzb8nRl8V1mlzjYmI8Xokg8eLHwXIbd9UF8PvBfTIout
RrBehvRkrShwLLCtyR7ZGCBXhkxjbS4KbMmgortkWbwsfVT/y1c9TcuZvYuyXB5h
YpMzKJ9mFZ3bkeeZPL4pWR+UOL/ge7EbLCIL3/xSnm/pTzDy/44Wwr1z6I+P2wsd
vqcVuiupipVcnAMWHeVOw2PXolv16XKAQCxAwaY4f+u4KC94oKjSmd3J8p0+pdA/
ei7koT4VERXY4p4cirUvLrWGEq70/y57TKGIUXizDrYeraMjkkIvL19KjRj+PTAS
GC7aHYYswxGxKBrrxGiDgFzmySpTD8phLvXC8NbpfeOIVTmB2GALNQ8e0z+mor2S
NTtH+NhscmFPbC4mLdzc1EkcsLsjjhDMPiTFXkztMwv1Dau55lJqQKTlDLK4GwMO
3SI1imRbZmFI7256d3U2W7VFwABgiRigFLTAM/cmHnRgI2E8fHDa2BEs2TRnuyFX
XPfDr2Dkfs6Op/0hPPY56K4R4WTVP4T+V0aLIzlnQhofH5npVIGqZNCf0TcAgWOz
xxrLbc+/R/Q9EaXwaIYj4Ph8AiAOUpJWdLaAQE1Xk76GJ7yr48kdKGFwbtifieEh
vC2OEjlgn7kGak7truzBNOZvfHQ6vBkK3maJ+B5nUXNHnJytTlQLBCtR5an4NVjg
xpRuIQg4T5HOBsBtqfzs+GI0R/4UPuBHO5BsjOyIPUnDZ/4FfOUx1g8qOpPGSFit
kqQZ2nhLebcD2kJOBwHTp2UlDlkkqaTvwEfbU3dqpzHpVlkizvucm++MBJ6BkX2q
1lUQrEvW21bHrhKX3LB9OAeV/T2uO2j8PnA4cVH0ctXSDi/GjqtjX9GfQX8cQtE8
tRPQFdrKcZoJa2k2hTLk04dZzChnzYpNR8xFbuUqPkq2VT4tb4KwSP7+rXmm7yfV
vL96Mw/cqSHd4ItdAjVCKnrV2inAqu58ONbRgXi8w88smiR3/05AGdHBZinfRfQh
95iXq9te5Ku0mx4qGwZRPAc9d6zVFaoYv8gBG8UkBTTz3vSgPBaVewtWrCclDLtI
RaGZWPj5rYtrfMeD5EE9UTCNXt8emw24z47dpPA9UiuAysxY8ikbC+lZst+avmWf
S5Z1xj1MFzzTZWCVdiz8hQTcv6iDP4N+F9QpVuw6+t0rq6npqpxRKpag7exb+CL8
vqSO5sV72Qnj/GlPVl28Tv2RHjhoSQl5hrnRoarcO1oVomGTdVKTelBn0CHI4EUm
RasLeeusrC1gD/8gS+4ipzs9ZyVM7RVpRumffOlZZa5REe78FHskrO7nLDTP/f5L
R5+uJnjHWvr5YAAGn4+zWo6EjtHPXBeGJ/vjA/pcEwcVMrNRNaog5Vc5amHKphYv
2sFFtqSV7FIseUXWVktRAJBDzkPSp7Ka6NGE6Rq7biltkQah7qaN7S2rME940wEJ
DF1yblRHUW3dPJrBG5iFDLghN6UfXbQsNxtOz62rJAKoMy7PY0YSaTlnS4bMmI8m
ErE1SEcaVS6ZatZpQUzrfSmc8EKArWROlJ0xvIF1Mmrr1A/eaWdeIzDbkyuyV1RF
/+GduRNXpOFB/ZhWjWn/UUKhellAVOr3H24jH4650AI4FaoZL/2hnWdY4JUdk+TJ
epMDyU6HFpVeeGVgUt60p3iCMeVn5kQGbzLgR0/H5NgTZ0m59W3onyEe43ixxdbN
0YYJp/bpbQhiFGACijUwQdBBqgfB+DedBLU55VMyg3n/YRZfNJ/NG4ivvMZ0vysp
xuNJqeGJe9G3VG7wdWvxXUkfnPnFoddOoTnKAnXd+fLTREXyeKIUp09n5D6ERzN/
ejsyzaBAJtsJTh1Ur3ba+Rsk7YNapk23a7MrBaVAr+TeXQOdWdPFy21+5JXB0NoJ
IeESXJyaTKCftW/ZElhWx9Dd79CL+C0Sdsxk4ydpA1YyRYl313NCCwuOMJH8AtqL
WSJiwHaL75MQriseWXdeP/sFSj+D2QujG7iZX1MbxXPhATwYu18QxUzWhVmq5GSj
jtW5zaQxLuIHp7i82PaesGzK70By8p0NrP2yL/Nwl0+pus40esHpgZSQ71tD4+Tu
k6d4cTgtac6wre9oT0uwu4PbvsbcwVUmGHra5XhCaqRtvAHPdZHNg4qo+54Zmqdp
l3i43oqbQHAZHg12r77G2VA9AMxr0iRyGRXW4LORzyYglC+CccHWPUVFjyGGiyQV
CImPFrvNbcAEEnO+0JTe+h/E0HFAWdqZWS79tl90u2cnF2CMIt9V5Ao+66p2dJPM
StKDprqiBIReSwear3ne+yghQCF37953yuIQE3YHSVDXg5vOhAEoXUKnKJrNueAU
qPslaXzvsIAcmtLAShP4FQ6h8YI8EUI3enWDrXJ+jDwMesBooriRspxsRar4AGEh
YqYRBYcOpOCGa+M6CCsiHXy4GMujiyO6xc3lN/mCyL95ELigF7jXgnFUIq5jmWPN
wJHzjlGSx9bVYpMOHBuG4OkCRnZ44PW2ePlEjtR6avDIkM/iZGQwEGewQmo+F5jT
ovPW+Da9qXuf4G9hGYFy/GkHAnAzhjGJZJN1skTaxgVHJhheblF06XO3UgRHNORx
KLmXVmAx/gJy0+Hv69IxpYr5UdnDCDUZJwYbljGvrFHh+3G9hGKqcuuE0SfxtSW5
JWD1ljamNxps1XtZy8Aw6zv0rpyBu1y3W8wbaH5Tffn9WcA/7J4SyFkT6hK9ieJA
+9s7OY9OEDhqgSy239OR/koCuIsqnnyG8eQ6CwXbUGTiLmsyvvcRkzajdjl/zYyH
euaRWjGbZElmNlkZyP5aqiDGum5ETPlZnH0AkEpUJ9IshIXF5SqjIEJqSRTGTeE0
JjiujkNV2A4iwl6KaXfAHOxIstEfcXwMK4Wu0YcnS4XqN3TKVsOy4/Fz9qazR2sP
J4VE+w+hs2GtAraMtRNjWcr8GtUbCYNDflFqygh+g1m3SkN3u1tgeiSH4bArOYCX
4XTw7UvyX9YW+dlhuGHTF5WUCzivTuac5DOiJEV46881L2Ahx/3tVe3RKqdGRU9W
bcYy/GEeA/rRSHRVOJWMph/e+qiheO3Fr2MhYAZmfFHvC9XNCryN71fe/wb0IXWR
0+cZkAKQff+eil92rySkUfCJqmEf1dETMAqfowR6oLeGlTr8QWaP99NZgnXd5Pgs
+a9DmkeWAWcZkuimdKmQTbP52uhpGFNSMz8UkA2jF5rhsBfUzDufbXKM70t9NQWB
darLMqDGqf2B8T8+jSas78XLWYWVDRCx0v4SKTupRZP3d9Zccbo93h5Av0A2mZfk
2/+ql86Kor3NK3nDEWLMe4Xca/gQAaYmkkemRGb3vINk9+S26BJeMDe/m+Q0jNl3
yZ8qXSKMr2gUIex79xi9meo8I36/mHOWlzLpV6RNOnpMlxYmWjc3lvzPbDFfn5WW
N327I7TaAK/g/OGmA/VHFRGXdu+DEUUCDwo4FMKvyWRAZW2Q2eh6aTqoXE+LOL6U
s02G7EmSrqFj+T+rJQwX0u9lhsIA2Q8eRr727rHN3vRWTJQDc0mN58qlLDoR7bxk
fEtmyAACaUowGdSzRZTO1eAXVmPtk3czwLnvdeDq6RgX3v2YvK9S1fdU93LhLQy9
hCZM4se3bkA8lcG+OmmNlAseTps+/ZaoJzGsSk+lQdvEFYsWosseouEp/O0SNpoK
nrnP2f8f+8xvL118JGlCOAfcEq2RO1HrvTj4LFqDldxt+eeJ9YyFhVZB+vaR3h4n
4knUZJ/re3fZJQFzvbeHrvKabKb3vdHoYC0yobSVi/uigeoyfFSCRqXq4oTa4k9t
cirH6ORlU0auRmG3g7GshnHMOkL53iVqv+2/oFWQ4HwcUkl1y/iA7b3zI57QGqQs
IlzWno1WLf96tm+KCy5eDUwo8SmAX2pyJho2o/S3B/K6hy+M8OLpd0Qk27rhPaG0
A5p09NQx+SZOgF9uKRF6/a7H2dzTcLvWNiZzFCHdFg/fRK4LXPUKWFpAkks5ATCA
jjK/3tuXOgU8YW9/B4FEVpW7a6UDePyJTzQSjQG2sD9Kr/2vTCrC2LlK931RbY6j
v2tn+G9JWMFDlWV58L9REkfIEpD601J7y+1WGhmSM8U2i+s9xndphVXU8qwRgcdA
r4TQ5qSuQiuYbdhmNQxirIcD17G0XFM6AqNOgSjnNRYvhuGqCqoTI2EhVdVs5W4W
GKq3SjEXKeT9nDaT0mH1LcamB+mXA/WKVqMl8t9y/aXXNEjqRVj0c7mxJG0kGGuc
MDiLkagRjOixRzAMMidvSxuJLuad0W6Oox2GWogDPNnIGYYRjZohOgZkMpVO1LHZ
nSYpUwpMsUqv2ywRvP+sUwLfHXPjc/tra3LR/hM1mzejfHy2+Jco/Kr0Yc8EWnXi
N/lTPh1ssFMdmSiz3gyCmw3t9VZdz5DJLhQVDJe6bStouHf0TTCB1VPVL3+/Ghk5
Uy1JydNO49NoyKpJK6OLZMz5iO0MOGfu7UKLJBrBnz/7sNaXQ5NmPaGME7VdQVsy
PsMEYg7hVKGzyjc7HN4VbRFcWydIlOWakPok6kKeI7e24EyBCpY/sy1rTyHcI+OO
H67xWGX3H9Mx2/dudrqX11qvbqs6rli6i7x74szmheg6Ynn/vH7HbyqKgy86LrV0
B8s3Rp9SOYJy/18u5QtmEG1U8MgBlDV4a9H+eOPuIzqfkkq9K2IIisf1Kyc0JKLE
N+zgMp1zRs3IRVj9MNj+sIAjNuIwlAmS65S6AfENwH9V6z8IAwwVbDBiJj7vYbtO
z6XQX1FzlEsDBXqoIdMPsZ+zyB+nlEWENzeOTmfrHdaoGxHY1CHM90IMQbjMkLIp
d8GhvyFtU4zw/Z90XMchIEZqkLYNguZLJiHRb0WXB4K1o8AgBbTfCCQ3it9cMuHN
8QQiXRAUHO9lkYbGLiejNoHZkRw+yssF3Ni0U43Wg6NvUL/LhRp9j/o9ow7DLdfn
d+yLuVJ5SgwNNfkbx9DfNxm5k2Kq3+xazqYNF6C4FNdekzLJS/haRYqmorjLxlCu
Hsb21l9ZmY8y0qfAaqvfkr8C0nEdxOfeXWAIvwdfjcdk9HHxdumAoSlcMeb/Mgm3
HmTkRnA5K2pGNSS6d3P/WM5AnXPetd1dM4tPlpskZ+qioHn+yN0cJFeXFqDWBAiH
XoEJ/SW0Y0ubKV3boOd2+L6BpDdwjmTxcK8c7gHM2xDAjKWUbpnH6ZM/8H3ppUTO
QbO1iNZTvJpOoWjAHpr7LeekfdMR96OsPhf/hNQApfBqHFKHEKmBwdFcSk+n/fRr
iEGReMlLAvjW+2hu0hS7pzAxp5xRLSQS2wNkxGoxk3Ne39XCgQDChYeAGsWRn7pj
rw1zEejKRKxQQFhYAdEaYyuQOS5XNgfAWsAzBcocbQjQu7h6llk8H2If5PiLYAxZ
ShTmqdNDBV+fQELwDC4XG9PrDpJBX7SD8L8C2YHlPKCjyBtbfIRaiWP2d1MqaDbe
Y5vZuhQPUBmKPBuM7mQujb+rS9vp+3T4xa4PyN1WCiKuz40YY46bwp27QAt99HbV
DWTgLe79G4X0pYN72R98wOZE0KIcrIG9F6mn8RsjidyfJBiYfwnPhQDMwx3bqU+E
iNSi6ED6OZO6E1PmhztiqJrJinrvUy1dz8Lqg2MxunxQ/R19uHZug6nvN5uQuj/S
hX0uPmP8XQdxo3MoTNloP9gKEixQnldTLeMYL+MM9FPsqt5G+hfR6BgC+JyPZm0X
VEwAVMW5NM0164UvdrcqMa6kIPT9w0LtynALJolFJ7oTuNfNqez1Nk5kzCIcfN+l
tyUoiDefc1qtYfdUs28dfH9c9RYGPcFKiPCVft2s6NK02bNFjG5XX+OXA+5phQ8V
bV3LCEZPmAL2kFxc59lHP6Nbe3/SYSWoKrM/3bKajQs2k/w4XEHEwX8TKZCwWSgN
dfGkh4nR/AM+iiOWOrDnJ+ZhGYnpRTCSKtvBseclWbICA8/0Qdx0WEMtPa+Z/q2d
ma2yC2Ia78ZTrjrXosKrVnveZtjOorRGF6rIkPz3HTovJfSdu0kU37eHKTVO8Kjo
zyujkx7QS++Lro8nKtNhL6iy3xGTnBnIDh1ipKIkm6zv5St6kUdvqoelk9Z/Z3aS
L73++cI+ww2HBdv+3hIJx+lHibmlnolGRIGS+zL67tzvf6HfQqJq54AEQArYsoTv
aik4c0/Tw+U/wi65YDfYFb3eNmg7ShquB37CsgFUfN+4iK0kQJJtYbK2OdjQpuum
ulS0V635v1QwwKd2qfvuwLYoEudJYvcWA3L0fHD4ehvcIAPUEOXz7lVaRMO6ih1B
LX/f1XeGMwORSey0RV8avPmnG8yUEt5gb1OGYT2xOJ8DyWs1764WNPm2KCqkDyRc
m0mjm4xOPKODZp2nELh+u4BfMx3b4cIFyBYiaLmL/98XmCK+fFduRAAvh/YNoVGI
lDLXLq6PnEafSBvFxsG95mJDbhhT0v3+PXTbxSIOL16gImjlqi439zPalH/jABFf
X1b5f18b44nE3JmRcMF9SRo9W32DxWhWxl0T/mHeQWAX03rUSgDg4KMH+nY4Pzuf
YtcgeG8kIY5zlwUQdcf+I4u1D2ktS7s+G0j9PKUn4HtjN47DfeJDNbshHMra9Sjb
v6FNHWPqB6puqlYmg2POdRfExZda2SU/h436ZOR7X5HR/zWPaNd53M1zWb9PSdSk
A1s7CM0HH+KaZuugW+Ih0zSxk5pmVn3PFmmyA57qXu7fFgxLD8zwR54yMjeJsJZ9
zYITjf0h39B3O0CfVpKRyd9I6P/Oh1d0vaMKScfTXYlnkO0mIX2HvSJdBk6Tjhh9
REjJ3eCgamFMW32MMOJTx1BJ1FKE6iDu8x5+ephIv66s6ExiEq0ByrWp6FC2ERAU
8AmjW+XIjLgod7ghOlMVHTYSTSdDV5q4meyYSvKpEsu7aIZhsUN5IhvTRbU9zSBD
KStgjP7c1n6MqDt3jggvtloj6XzwlrrjoCWhvShJEpg+5I7C9gKwu4hf+gKzpojt
ujzAQZ7CxX/2xFKUNrbtTX8TIJbtrFkD8EaLupacVwp/iBo/hJeUWJpKApi3t8lz
JoCB1ca89g/Bnqc++anNSS2DMMiI9EBJ6WI0+cjYLYBJLwj+/VvmvZalTwFQEMel
MtnGHIiDaZwuepqWCvph7hfBGRu3iu3Zkma6H477eyhcjvZTL4E/Xv9FvOKTQOi7
b9Dj64fKA/ZWOgXlAwloq86446EHq9yblqAP1B9QooXAMzJxCybEg9rT+gz0G1b/
v/BLCMboNu2zl6DBiUzY6z0jbGYr7CnIo9SxDUmwGM5hrRL7cJ0ivvy6PmHrWjlN
0lqS3GcMAZQM3+w59mHDjocUHvzTKnge9DSdmEqIvtiXqVWFH2T4k17VrlydiNyQ
BMBqE8FoozpVw01pb6ogSQgiHxev5PnBy0fXruzD/A9dsP/EaDfdcFGlUbXvQc5z
zJ06JN66yRmCbUUSDFf6gmlCPziVgxtBbHOmSXorkuALsfnHJioD+8Wpx3MSnZVP
qSylbGjMFQWVfzbN55Jepp+x4nZLRZN5zvKekQwAavyNFIrKYTICfZuUK9RLaKQ+
ScrmwmvHbxRfTyJcBVAHI+qITKd9CWz2YN+oj4KP1zMmyBja4oalnfLrno/bYXFL
cS+DhuR6vWkvWSdLgECexhrSwtav9imARENEIkkejEiA5ZWH1AQNXIJJw9shXXtQ
yknmeaMttckbUHMWjOcHHk/odGSIsp/zc1GcvJppqk1ZBV+1ETcamnGa3jHIYZGr
ks4c1ITN3iadS8XGzhTVDsbJyhL8i/p0PYyPmybneFVjCdm8htek1Yqg+oa8NAPX
LtO9m31Yk7hUDkgzxLos1s+UXHSxKanhAOEIsoK2NkhpybW+SWtUE+yVY7TBdkpW
nExjBBIYppJdzof22twA7B21PUiOPWFuAl0MKxMn+br41omVfDJ9x3d5nO9Scu5h
JE2vlaKFekOJ7HHbhoVPEE4Lban4eBdoxhQpyx/9ZMK1kalBZu8u9ylUyy6VyaaT
tc+ENPp8F3uNv+2YORc3LsBkWiuJ62QhZ0jfKsYOwQa2BXXUX09cirk0+CeZZ1vT
W5SvRwRJO4hhe30wCX7zg28WV3vdONfOpl87arZbJJQ/Vi0HW1YS1E8Sobuf501Z
NFhv6P0SvY0EGNMNex2xdxXiG274Nm/2FEBWSW0D8dmMQfXwK91KtceEeXPSq84q
OpEOGaTlgHrQJ+Ka5hC3h2vJecJkkRtWHj2OkNTrWdtiMFnsiCPm7CGS0c7UQEYn
hqJwbsaflDZH9NlMmHQY4kjWbpTGnQ/cffZmo96h/SzTR5agtdl3doxk78RdTZnM
nfZBa9EGAPssEnZX0ZN4Q3Hu+m0AbO7cgkOAlwdYsEFoDrLqov8IXKhQlcy2NuPb
2LiekVrUUylZnDkVB1DCjaZYODt+aIIl+2RtcVBOaKdCxVFAhBrI8Qd9Q83WROIN
S1IHBNYuXl1G5B+Sw74xBd+lN038vhFTicrfXZlAxF4JDI6jSKRPuat9f2i4m6OY
uvi+M0t+osHI9qJLeiea4O7R5jUnQpi+ekVcROjhglZkWyAdTjk72qkv74rJ81Sb
THYXbh6w4Rz4v4D1dwtC8cEsjQwk78KpAywiQPGoo3ma6Yk90zQW2oYtghQhLYTx
oU7ZthVgRJP8G6xRibOX/NlyaseGeogBe7B/alXCSZurdtTZJy9b/lv055ey/p1l
TFAI1L/oPU5/NT8mqG+K961huRo03PDmXIBgjeKGIbNia/NT5SHF/S9q+KJinpDa
wao43aKNJ+wdBoc37jTWX4SPe2+0gyLCoX86MPz5KdYjKkT0G4y8POvKovLbiIr8
sDxbpZ+uC7/MUODIf9Z7W1i5+FmpulDVhtMsNycspLMRAAz8jFTE7RCGl2mhipsh
s6qfmOWvvFZ+h9C8yxWdy/+0Q2QLGbWQeaPlXHGApdK444KauPSRpuvGI4vkyrpB
ggME05sVK8KdPoWEbzrLJrOxkqxJkxMGT2w2V2iNOyc5wET5x1NNbYk+pdbWUmn4
7Kqr1/IO+x/mUek4fbijsC4hIcdYOY/7GBHbPJjKYW2H05fS+qKEaf48pLxANo71
8cXN6sg0bseTvAAL2LK9wlioZjkjJMKrCrG15YkFie6bRg+PonMFLYtEAeI7GUgM
rYGXae2wOFPvzO5kDucEFOHJSeNEJkEhMgVpEb8gGhAnxDj2SU9OFmrcgfzHFInd
uInKBmZYEb/kz8aOq3BV96LFd4YiMxdrltELHiPTW7/LJal52idJTJw7ClPXdiU9
M29TxW1e/PLUXgpWQLEtSvETADxVepTPBIyBdLfc+RrJdqidbDFTYJ+5fiQdM6XQ
A8BdnomKVzyUaEWs+A/MJcfff7Iqml5ifY5WcNtmz7poH8kpWJtuenf3dGWSKN4z
aIyAG8nvw9UIF8oc3wKdyEjVghblYQl9rIFtj10suFhPoT3b7NX8XCLVlOGY9B5U
E6N0/fsqtxAITE8UpHcsQY1ZSrC2CYJWKv3LeOZjBQlUbNxbPMo0tkSfo5DKW6Xa
LgmetVpXicb8Ddj7keE6+wnXSD1MY9kngUCGfe9p+8Gs9sFSmnoI1LYbb8pUmvI5
QG/fzh6nS2c9F556rjiRnbAD5lUDrifgkvSXp+mtaBxNUv/1R2fvv6IdAYj0kZwo
6n6+ZEurNBYgrz9lkZEYeUGA+E3KsNmf9YZq5z1Gz4nLk1VsbgZ/qb3vGlc0WkGu
fxkAbiDITVzC1At9VXzO112c+4CinbDNUthSNTs/YMYCVhbJRfxYz4hox6P+AdgW
lPGUv2AwLcbXiypvAGzld0+HFB5kJ7GXAij5UVTEv/0Np0rYxTKnmOvBPh6yTOUW
gb+eToXo9CPojYRWXa2Wq30fkSwGqQhHin7If4bzcP0AO9eIvYwOk9Pm8UKDIvmC
vfMjjllSFhENLj8uUSmH3SznFZfKlOWE1GeoeFr6CPSowb53ci8sqTF4EILw5zFs
nZ+XL4HzDasZH1K+vHjEyMDV7eW2EsJGTvXNJyav3z1DjB1KnzhqjSztf84PFd7z
mUyIMWQwoEkepGigrCM+XMjyF0zeHsAaS+HEmgfSAi18IWcMim0TASW+P8dcNep8
0M6PL48oNmUztde1TAplefL7NSWxOrAWjfIBLuJoIi21HtzuohpDqCIAeI5Eew67
OeHpH7njV1eC1u5z7+fj6JnMEYcyNqUPSR7N4v3sIhIkllRZ6YUyip3qbzWYBG2U
iixV9v5YMOtxyjFiCUr1razfgApuQux78Kew6zBedx6JwvUQgryfRGAB2MP6sS1O
KXkIiWqHvXoipzbEMDTO8XKJbPhZK6q+5f5mvM1K/bUuBl5fZ3PMn0VIi7tVqsES
oBtasBOBy+pxkJoTJ5gIXeh2uc64wnbHIv3g9OXG3klFnMkv3c1uh+a/Lwve9DHD
DwnnzEC/N1NDfBqjuM1ldG8SnKODkctQEYZ9txFQmVqHnCCdhjKMBwigC3ldtTkJ
PQm7VJ3hNGONGWQi2lz9uxdK5rcbCRwarCtG+jPHYv9OCoa/Kac59TdDpQuwc6jD
G+2S0xNO4HmYnGHKufbEVfdboX79mdBEok+sEp/indTcySI+sNXqUbtWk0dr/CQf
Spfxy4ZsdfQXItLtVXzijAAOqWFOe01lhTaj6iDSFQ6g01iz+ItJEoXwtMJX1mb2
KKlPhEtGshlMP6CBj0rAYD/my/34veYu3QLVZm7NCm4haki2XBR4K6kDse9923Ue
t1+QUBg4JaZH/RTJagBC8JObYT8DAq+pQuW3q81TETQqamHCkqahDIyZfWT+h+h3
SESFyrtGbOElXCwnehX8vxxXvS6TgNaWrEjfXZN3lKtAvmK+n+7K9VbbtCwbaDRK
HBVFN7nbyqwK36mI3wt7coT431krF2bpleKNok77W2KbjEiDqf7bj/ZNiuVfTpku
FZHlCc5R9/y9SJJzMqJXsS09Bs4IfzC73aitbTEQt85FrcoDEfPcmCR8v5DlZvMd
jQSZI8ELj/MsT/gA7MHVVdGBStPBAZ22NmRM5zaA1nP7RxJaNGqAaShSAOEHYcpp
irWSFeDodwPiQFB8/ObUl6/5USDBr5XPgY77sizFxClP7uJaQ1X1P3TAAce7cyyM
J7jtkOa/+Gp6K6MxPYoDEPrLp1AHHVpUiwog4Ryb25Ed/WVgAiba67NBJ+buZwoV
YLQd83q4HXqyjyqNg7DfNoRhYh+ae+vxwDd1bPt/tL5sEzc81rTTdQ6wzMz+4dUF
TM7HC394wbSxcyM8D8IBTd7Je96SdYMRbRfKA5sNkOVPHn9TAOqkllUQshiNr0j3
CZb/HfVwOpApHmO00KWV5mF2CkMIYUN3N0G1Eh9X8NxueFRVBEDvI08twZGBWL2y
XcAZaTf2LV8peXoltO2ZyzFHaZt3fVAGdax22jr123/MYb91jtuCRA0bYdpPfFUk
gquZj4eNaZ6mOkcgtc6CXOVIrGr4+OfGvmbaxhbj28i78Ugtpwt+tRZ/v934Dlu/
P59FUJTkJHjfH07s7hbtHgEpTcp4f2UVa5VIvQg87efiMtEyrOroPwlI0/XTXwav
oSgBu91AKH1DF6Q0OmZhH4Vx+X+LAeUiUPxu2A5OSGDYuUuEtt1GXoWHzdoKUQsC
DKyVmvcAQXh/oVZ2HLj6FBtCRk+4Nmyl/P1WnLuRjVGS2JUvN6FWQW3J/XgM0lfp
mIzLFfY7tilVycyTOTt1zD9bHoHIJpfBoeZU+HUQPrUDnI77drWpLOtEG0fyQxX/
wbM/q7uOpkrCaFX4pwFXZbB+FAKEh/W6a4Ur5H4x/xcxdSouDEqUwtDQd9S2QXkF
8RyC4oaLJCye0HW9zRzyxVJy0rPMIEADesUeJbxFMEIr/IuSdIasofBhZR3+UWRg
mNQbXddMygqnEJ9Ze/FS5faMSFzVGWNLvZAEfhJeSaaWk3SkLdrZ5EBF5kgCeTrV
m3SIEwMvY/bwXfUcRuvRhwsoqYJo2NMyAka2m2YvzQRDdbApLYBFtxAbnuXIkGF/
UE6XPnNfEHdvXGsQXvDrLCQN6BA1zqq/MGPlNgYN+z2BrWbnpkOI3dPwPTZRpaKJ
XTWkuFJJET4j5hfftJUu46N85gtOwn5EFy/q+S0a7cLZOtDUuyiiDwzad59f7Cpz
h0NcocFber9XIIATg98/G9Dr8uxx1EmLrMljZOCy+OF2s4m6vHglGNKUwsmJrHZW
DCTZCYfr0ZHENhOujAOQtY0bFulwW7+6uUyHgPplF2rvRrjoPjTTo6fuh9YO0dM9
kUYMmHIEBL7GoO4vqVjGnoQ4I+mEmnCaglDMdjH6qEStINdS1xjMIomCLNQi1vi+
sk0gBu1yiaTNvEnhHQkmvb0bB4Rqtp6QbmPOd3Sgxl4tmK4zF2pmjDDDeq5PAZ4e
GcAL51rd7U0cGu8hn/MuyygkDvb0fRwHY0H/E/YcEzs6rB0XrHgXroNzn4EDtJYq
9NtMsVMnzFso0JqQzGYg4tDZRWAh0OpbAZluoWzw0D6Mjh3nA6dp8pi/FXR0qNIt
KMCF3NUcU3ow9MgZXRqKX6Ml+wNpMua3LeuiygA3xJGZw0lZClcgUCkAfCU0ofYq
GJr/bGvYZJci8PulbzGzYig6O+toklK/Nsx2JhmyVViVZNDPv1q23PObHfF/D3Bw
cTZBmL6TQs6J604OOc1YXbbMLzkoXcds6L1UqfDCMMNWTSSLmxiK0wujGe6PJOin
2xSj9Ui5im/SSB2q5v5LrOYIh/mbkiOa1zWCPbF+Bh2BBenJ/d83v/XvmrB8jm0i
EdaUVmJalZQDMg9yxJlmSsyB+5MR4Y3L394h60th9PFzSOn+OZEmmxTdxD9d0/GF
ObGGnP4XGQ28yzVHJMrA77D/Xg/yvFQ/qRz/q+jMUqhdQCFSCk1vBpWaXOqpSCAm
NYaf4dc1OyXxf02zudDxbsSKwYVSRqLGlBzvoixJJU4Wa8//cPFEryoVZdyhUvx1
g5u4CUSVStn4H/yFJ3J1cTOR+CdVe7/QgS+yTAH4N/ErlfSWwNChLTPHDNJ9YqIt
4jgYQTo5RAck+jLkidMP5KC1XPm85aXGlj1lV7PYaK8EPy3O6+BtfHHAbpZeX8l5
ldxAPx1IAbqOcktqMHh4Hso4aHDW0HBWaXoV0rPOw9J3WQrdhuaC3ihuWrgoEvLc
K1LaRss/z2Fcqt1wBiKAFzDeOGtrEHhBt+vWj2rdtmysKcRrwlQQ6tFMvUCLgVAF
b9ICP9dgTEC9uLmNFaB0QblVxp/BOEIFSEwi6wPgjPHWd7MukT1DxqAVso3EBS4S
mNGMgrL4jAieYBdFMzIRudhQe02egwWAjnNLOpcvgDosMQhu2N7nejdiZmwSNQlr
DssI5+8f9/DQ1sAnICK2Eijz2tfKty69kqjGSgemf+PRB0xiD73jkFX1lD6D8wAP
9h6OtDyzi4JqLYd4w+JeFJGAnfySkq3PkQM+NMZAi1qD3TfIkhPX6MksI/tiKJYL
aqwNo0gFcmA28nX26CqSQwNEDY4OPgAw1oc/8Hpll8yDsbTAggckDrTCBH+X4FdD
xP6TPDZzl1ml0zz2YowoqHiZsUfZcWBrABqec5QrQjwrtXCCKUqehVZeIfePh8x7
1AmdfPjuJi4YTQvm2J5/RXlOkpulB90cCYyOJyOJ2GFx2T01GUuWhZ0PnzAqKR6B
rcPklH1YQfZf/NJuA7srpugZ7ojmZLivdyLUtyJ/+gHmYPxs8eVvn2vu96M5BoSE
vNTtTSLi80H/AfuKvas72rJxcFGtYLpYWKmy/o6GIQlSLG10YCosJ3hUwIcx9k0p
6nz0HxcrtvbIj5rPfb8OWEBpob4CW1h/3z/3r0N6DIgeyeTIeavtUePfmxojWpJy
uUIApH8d/6L8pDc+NPfU6BD7IsiotHfY0K/xxWbvTXPT5VBpfjhIQ/sY4QaGd8pm
PS4UFf47oTZUuX0eTWKOz2aVdxIR3V879IkUCT9kaC6wgXrFonWpZWw5yh2WUaGv
XmKzVWp5fuhFMAaEMhkHWoAf70x1EDFTz7yZE1E58CgP/p33OcAwGs1NVREcFSet
ZYg1SScZqnntBx65/gXwIcghzNrITrRqpnAz6rZuPsD3OteEsQ6TkTPCxjyBkfG5
nGFWi7RnLQZ01GZfic8qpvOJ60abcTn4i17gb9uoJ0maS3+7rPTcAcYfdqDtLcHH
SG1IVcns8uXthF7tbCryNZwXRq1Rv/N+65GZZcONfHXcE7Ze5AUYUMOieJVadduS
sRQHXXw67Gf7MDsofrRDQiSWCDsn5jAU1d+hEBCGNfrcnx5BnxN1d2n0KyZCjfGu
+/Z4JiTjJJACGS3Nz6ZFk0Sf1B6Uf0MVTqdKydBpshGjfu/tI1CndQbdTKFUEJyf
NkNEeIDwcTQsmRgQCjWtO2SjGnMlutlrDPPCpRnWgwDdZX29fP1X/4S/8nEKePUC
BZEyHLRL9RY/5BZ7Z6i9RIY3mEmh8s2CRzpYwPSdJldr7OPM0lo7c3SQzz8QfsZb
ygeSChtAlj71SyGtOitkG899zAp8pOy4QD9UllZAHOdeAbWl32wUC21WIqt80il2
q2MDYstU+ZM04VCe/LL/zPSb/4iSRm/a4PuNx9t1cm7ZbcnJ5eSSuFWYDg6etmRg
1LIwoXODJ6ROAN2I/RMbQUzwwHf1SNefLVu1svO9Slum+dpz3FIAs5zFWh0uyyfz
lhzUUcApjSOpMzl8tPvMD86Pw8rUl7MFuH0Sh6g6ODPHzu25nPVlmvtc77ZER8xI
ythk0Np0KokAH2FttnLqWZm9JY4RIza+JjJKwv+3JL6YS9GYo0tmvHU7pNxdw9lD
9Vwp5VVUQAFFPC/XRXcSdNUEBllfwC7KfA8ZnoaGGatLSDJ1Az8xbZtMijMQD+4I
nqaVknfDHZkp28cQvUlKI/yCi5K65G1wu2oxYa8vGo9gTXDP9DDh/3jXwMWKduH2
NKwzoOApCjNc2ajKREf+8DYe7gftIOdCkMOnKlb4DzyuHxwGbg7du2rQlxE9Bv4V
OmgoWVbMoGiYsywi0u8ls1/Jw+dB1pqWAdE8Xkdk5zGNIeFjWwDS7CCj94pcaToV
h3mDdkPCyOWc39n80AzMvLZoxkRNsYSgMMbU+uc5++l9XDKtQFEP9mMUh/sZVnZq
Zq/tHC2jc5fVebkvUnS7CJ3SrTNsMaBdatXhkGtqshFxCMH9nXM2EfOvVj9WktQQ
2KVhuFRCZNB4du/GImKifAJexjs192Zk+HNir6tGAGhlzNSxcNh9ObRN10JIUYP4
cs9UkN+/5RXw3zeD40R6DRaygCDZDQpw+5gDq62BuLIYRMis9K1UoOe6Xp6h62ik
NrJwnKAx0COl7OoGXKMxfkmQi5UfcoO2YERCwad6OVHuZ9RihI/Dm/QZX/AmUATC
Xhw7Dtiao9mbFZvZ8nnYyy7XYDeGXe/T9ImXVWU1lx0Sv7Sd8QVWIpGCClqZADsl
0ItS8hInkYSeliPt4/avWjTCqG2Ps9teiJZCJwIQnuA3sRP7Cvdf7VbxN+CenAvA
QTX9YIs1AJFwoQXr8kEKSkHOD7XOlu4wvz9Rn9cH//PIw82pxmTsJUAIrTyAl02m
ypwUNlOn4Ua145m5+CTOgwvO8z+gayqnDgty0uqgZZN5zbWepPiMPcE2+iVla+hl
CPhQ7IAiAP2PfWrWYwtxz2rcDJ2Btjve5kcDYggYxXEFidRZhSYNUioSFUoh8Gpr
UuIxanlel0MgdA/XmQaVIRAW1F4sYHADxdtP8osJzGiO8mX1xiOni/lMdunICNUp
kR0CfhrxjftFgP3EcKR+M8Pd6+nwXECJ8fJncNhyAuvSy14DYhghl1xsy2KI6+xC
2glWDg2hEbq8dnfYUZQ66jSzi45UsFE3uuebMDQbj59GS1/DGGoF79CNjfycolvt
yRZvJ7Y2mlAJlMZLtKO6uOS7lP+blN5ocx3QldFj0SjHH7b1yEnIqfyjONxzSknq
mSMvYyX5Dg1J3G0uywlp1UL9VdyZojVdDIH561QzBKG8082oikK95c8D0D1b4QvZ
+y4+03hxU0GMtYRCYn4pmLBlXN4kfDq1Fua4ltwBpYF20IUUrIDlkVjwxsLO7/r3
A7wyi6NC8xNwfxeYr2k9U9PY3aRRoaiCQQOS3CUDffjM5FJBvmhu3h1PdjvbUjU8
7PaXgRqnlHiNPvfzKe1FtnUBDriEL5EQB4w9BerIJXQttFgZu3ZtfCq5ZvDEoChJ
7rWktsKSjhbniMzezPEcp4Y/ontVej3uBSgCBWuhdScR6JfPhKoEAlqiI7xOznGT
mMUeNOMhiMhRGHH14Eo3oKWoQ3XgkCCN5+N7YlXA7GEtH6qL3BMdTPr0E7AP41ey
3u//17fIZBqygEkJGqmcpEna/Q54SpZOznQzoYBTnUb0jA0lXfhxuefuL+U9exzw
HG3/eiBiFad8AdhmZaI737rvSUBmS3Nprh7wNeSs55C15CF0fk+ifs7ulE/fEFAZ
OgRM7BSXrXH/pUrxumpYNkl9jXqPwEU6v1m1Z249u91uP4N63Bo4u8rveH9mWSHm
p6XOFqWUdpat0EI6IyE5WeGy0jrnKmeh27BpzD382lSh7PAfcCUdlEuqPothiUNS
3jj7ihPMVC2E7ieGyoVnwS6dWGSgyg8/iK+dO1Udzz7MeyHDP7IZmE2TpjzrNccz
pI5x0qGgdDdDKRe6QD15jl4sU677/5OPimqkwdIUKh3nSQ77DJt8SrrfXvbMeFfQ
Wuzbc8hlqYh541SEofQeO33HAuKR2GoRqKsQPhSpChhweLWHoxrTkpNFFZswAUgA
BlMsOhmdD4exu64eR4qPoXUx41fZaNlLJJfhUJSPXl8pZ23XdYaM7a4YjWTlOXeS
2K2R6U++QK2DLiwiEnMHE97QcHxBlSAhl0fE5Un/7C80cHgWJIzXu+Ub+dW9cx3q
nUg3AB30qp4hrfjrQNeivPyBnTh7VcC/gnsL0zwStE861bs85UKZYHF4Yx9wE8DW
H88G8xa/uBeN8sC0jFJdchnCjkX0JVJcpC1+LgvQQUO1tQWpOh/6K47V6aHzeTit
bbwgTPlLh3zOoLaeJiOlQnpT9oKLr34hhs0yAi3OihtNyWbnhOz3gMKDiSqENGL4
Ycd0/2O2agt0DYKSZZcLJrxEvGrVTMV2vuPU5oGdKoN6t2a3Xv/OxH9G5ytWYOW5
xLhIp0Vt8HhOku+UbcRLWsWoI7mp1zKO4KIZDwNHmgOQlAPLANL95H5v0lWEzsa1
dDFI+dCpGGyhped0MVTm5xwnM8l89pKYIJSxongDllxozhG/P8YzqbrmnIY3elv6
qqVlZNQHh7QFHMzpC0KT9Y47SuH/gIwRfaDvgaquBdvFfZtSG2IxDbc5QaDQkp1j
rQsT6+Y1jgdOHRf7i5Z4R9ugS9FsuAYrF69BPSdDxMTjEvUaX1BTSKIp//L9XfSs
YLS6v6VTge2/lk7D3vMABxya30Gvg8zRP1Ybz26FxlEVrNq4VvuwXWhL2CYoQE92
W93WfX7PwYeFmlfjrOK/iPJzFjnb9tv+GsidlnJqRL2x3BPCKMAsBZ7+/vHDJ2jU
LZ8VzEvMFmuP+Zx6xvXeX42WYMFkLxgMcOkxrjD5HyVbPs+NPPTPuQy4VEgRnpwy
5WargjBaslXcqyVig+ATs+vRZsT3kxEVqjlXeNX8CxFTGkjyndSQ3NzetCAZjsaS
VsQHSGJVNHJ07YqGCeBShKva0KFIsZ0OxLirNxXeo5nq+ZloAJznfUvXNIPEpEBm
odikA7myE/4d/z7cbN/7kisTxcYP36uSg151hiqpgEJTzFlFFRAZ2YJfGodeIwg7
rwJGvS3lTfwCIky2vD+K9YdpoOHcbiFcdJ1vvOpERdDAer9FJDfhtQ1kju1QwUX1
sHOmmT0yTbz67VZrc0ZJFoEEQlTbFBvajlg1uKjm+Vtox34/sA8YmpRa3X4Sz+PN
BdWDxevcI7Su+TFlhDjnhqK2QTBe4agyRlrab+LySodEpC9GahNOCQSpAWkJ3ZK+
0JuuEhc5rIfJV7QAKKmF/qYH8p4kkwcZpVxL/q6YMns7EUg3bWb0LcMpd/c0zMsF
iQlLB1JLQXN0YSyXORautHmUi2toJuDZN6tEANppD/34VXi+UCr0dUvnISU3LhY8
AntAy/CIhG/SlKHO5faHEEcp53A5r/Byyd5X3B4SDMhmhoJDmfyMV5W1HtLBZ4sR
vzve7KBMqBl9wsnIZ78C8Mk0Hg+H1r8+jb/SYkq81/IMjGYYz3OPcLu2SSps6C+B
9h2KikOxmTxU3CoENlwIeU8oHee3EHbAH3oDDUB9GZ33pWbiTsu8tTWhaEaUv6JO
DnQcdCnkJtq4q8aU+MR9yhVBFhDyeK1Lkdik57ZqLKrn3ThxpHtlVe/sJMV2kA5w
EzQyJ9IQiDfBJngZ3KIE0Z1X0twYsrfahT1mpQOFPFtb/MGU7ZpcLqbU8Z+kQk+L
mspEJtXeob0o/KR991T7ekcA1tuTgtqce2W5CBS+T0/aQ0mVBgGrZ06CHGHsnnwg
7ayYw2nNEcONgLAbQLogCsDw5tE9gCCfHShoCbjHIXEgvZXxrujq6ESxErsI7peU
lmm6eYeTy8ysR+SfHbYDEwF88zp/3RWC0xJ9qy/uv4Hd1zDT2NYwPiLiFeQcN+97
ydg56Cuq4+0X5vyJVA2jHmy9onfxz3ZO/Cqv+j+TKrYcx/eAbYhvpBVnmX4dBB3J
k+UauoiKUm9LGPTllXuEaRJ815LpO4f2cmnjz0fv9xU8LQNVsXz+Os0CtgHMKbr0
+9/qy9QG4ZATzahZ6sEks2aijWwJ0EXvA0VqTSVoNp9CEaBItH4JEDjGNEgpRHj4
VHKdBQpeey1LL0TmDhw6V0Dplw3nlaUMiC+e5zZ0fuFQm1bugOe8x92MWfi380Vc
HSpLzW1gFWE9bhS3ERo0om7qrVR/0MnXP0nixnNuh6XcCVj9GkWQfCzH6QBLkVgl
Lv1PkzEpeNAdi8CE6QRZ1zeD/YznzA7OxUOKdbo5AXjWfWHlVxuApNhILrQ09Vzq
3VeCvCzA5eRNgLj0IOX6cV7XsmpV6H+eAde4uosPWgoxw5F7wtTThIE44GyfwH6s
5LLUnlVCMBUtFTi1Y/aGoM3yC6iuP/QIpDET7QPCK2IWFswEb48Tqi3xydwWn163
gXRugc4ftrLkf90R3ASYch5+eX/RcdaQiJL0J4PXL8LdoSyxHTRlrEicQZcpgxdl
eWiaXW8Zkqf6ieuzScKlYU450Tj9gAG38wMVTN7M7Epo1OjGyzguOfi9GklS0ef1
ETMLNovELeNJ/X83qx68HEqDxugyG67+i054qrAQXK5xfy/4SWGMogkeVWhcf90z
Sbkbnh8Yx6f7wk1KR0DSkeLGOmW2MHaRQldu68qVM8LJQiBUFPYNZfgJOLj9Ufmc
o1705tNuMeTo4bn5O0IAzvXq1pg+W0UG8xw78dckw2H+IiFJ2kZUygLvVstEpuRC
jjq1Hq3OadYPUyrriV34hXQ7faX7YJZz9FBb0X9zD1MaMyYzVFjWuywK8BE1YKRq
9x+C8EryS9IPJCvcMK9RrtAhC0rjHp4Q5Vlq/xH83jRvgYa897imvNzdslzu6Im4
ZeEzO4w9sbEBW5+qPPIzp/92xCRgcTu/25nhp1uZGqDw4PjFuTOeGG2PcNWNVc2+
Pb7rN15RmB9+hKCLP3agj5m2Iz1b25nDs9Fi5q3t4eOJ4HgBhX2fbwTquaYNt19p
dUZb5kAvW44/VOwq9jy3wOGdDEMAaA1W9MKd77nTxs2zGbuE0kq6aVMDJVlK/Z0j
k0eawIKZPsI/gWx2OFfJOXkMWVyUQ1c2C8qsoBkeL797iHIezWjMaZYG/I9tgKfp
w9WdNTq9KdU7fcazjkDulUxgZH9MvvKKik4gIJCf/cgl3mu3v73y44CV6XcIT2Qu
94zKXXoyyAqHevURpzfWe7bN8K+BJ0B6Lht0v9UrA3pksM1TD3FJ4iXVkA1u+8nL
kNwaM3OMZ53pwRggQDP6pW0MEXabcWL1CUKVukgYb1izGCTb5JxHW9KD0k1XPfe8
6huDJtghMX3REwivlDoN9YYEcFNMscBGlU3mKx5mmHEPbPdaOI+Kx4XOzy8BiHAj
jCcSfB8C4YnDfhvVYlety0T+gJQoUMn51C/ppj6Z8gqEyE6CB/Zl8C3FXU/xEHh1
JfwEDpc+OfcJP75rbOeHdhdv6rlpq24r985gyWc3/2RTtw9Fa57TaEAXjuwPTQyW
6Cy6k3yNywjQVKVtxvZl5A6BojmWASHw3Q4dOAMV8HFQGwqf2XgrNdoylb/PTlWl
papVZS90FgdolZAWR5to1dXlLr/ZJEGZZ4WlGTJq6DInS2+5ZiewDHzr27n7u9CB
oIuZSsi5eRgEgvG1yhSC3436+V8VLYXP/AP4QW60IY1dszLhvLiA4jx8KvB8muyE
Y/Ucgv0N20eDgEql/NlDomyV5NizTKYj4gD4SQ3lHmldewZHmFZ3PTGduqOgm/lB
6fNxhuj5X8WvEvo+05x0gy9qnJhDcbLe+jPTaFq+uEJ/OdGjRToNkcDFfb/HNaR0
4HKySq7h9WJeHO49dlZN9sujNeAHijoSJKxQDZfcyFzGC+V4DUqPqLwf8llEv+5e
Dyrb4le52N2zQLzhJJ4nJdbCoYnmRQT7GzrLz0gO8aSJo0FqqbOCCD2eT5a0jtf3
v71ajXG6JkH0hTId0Dyc5iMTs2giYJN6wGWr2qDQA4LvnFZ9aQdhpS602vqgSipB
IYWj9lKGzabdVlh7bLPbuLq0Q/bgHDJh25xAUI7PihPpcZeRhIaPiKOgcb9mJlRG
2WDiHzPXqc9cePrvLjJOjdg7KnJunrK8BNytLpZS/nnQK+D1rCozPTbsIYufKWG5
Z0FbD09JUxSA+HwkxdyEZyvQyRvQn349GT3hEtUb9xmzoDJiliuamEOibbvkWTO1
SlDKf5DFTl3wlR4bwupRzvsZKHrlbC54zDfmnkJLtf0RJVEguf67oCnG6UTWA5oV
Wloa7B0/2wezTyv0iDcWDVYl/e1Lj9aMhieO0L6cZeZAp4VlrHdTLjdUfIahDRgd
zUf0Eg5ovVIu3Yit+M9qhufmYX5TfaDAy8ecE4HJYHAqzmyCYP2LA5PgYVe/sOzh
9ZI4bxP3pWDa94nQTOnnzAWEfi5J1MdzgT2+1UW3R0hZHYX8FMur749d/hrlaYH9
dwlOyx+l4m8Nm5aksSXpaQUpfKYdhkDOQBSP3Kw4HXTowhH4EWNYd/xpRGNV9hR5
eKFQq2Q5n3VtsCAQ9npqsIhlx+qj4RPoCg6U7S7kuRP/B/RfJxYu4gXg7itNgFWj
d2TmzLYUcPFilq/e/D8Mv6NDr3lY4TrbpFbyyd6yB+inn6N1+LE13aiOdpZ7RUi3
yvarFOXPxyIujsL/Qd/qkSEzkM0jetLlQK3BndRETzWbTe8XAXmd5UryFI+DJ5MJ
PWz6EvOQkpp7/2xMCajxcySLZgDthkU3E5MzSWuWmKHDxLlqk8lxxhrDA6FSzJW1
9Nda2wTnBQ/9gm9cdGQnMvqe/Vrl7Vk9s0cqPJy2yBwlnlqgc1+S3YYBRRI3CJLY
ej/wDx6kgseOB2PNO/vWjM+45seGwwVEWsuQX1fVaBurZlvDz46omTXn6PQlE9n4
gXOvhxFQVDl3DHaB3yUJnYTOJwflnBGn9/u7mIYsx3Lt/57O5CMcIeYd/jAtDoKj
3zHV6ZE0d96ipVhM8xvS+lXOXGApuGclqmecBiy5cc+wS7jW0Ymjn3AtHxRaQ9MQ
j7S4B4Ymr9i9AIglRoGjQaWbQMhak7m1/alDqYqHc6nL8imKsPLO2xw9Uxeat+rL
xBemiRpxlXiobyBshY+0z5u0VwqhsuFyKqrkytHfhHinGed5AOLMUdtNM/NERJZa
T1wdzOzsJtj1npmkQkeuXpuPp6FvOZPJOiBSmUgIARB1ac9c2OzcyCkzHPW6W/Og
BqOM+Z/8fO3WdsO7xfJhQqYtroLjK57UmracwYXLQfsPI2l/ujz/pPbDuSWhU94n
O8+4xP5KPMJi43jS1QSuNTfOAaSqtkn4XJNMceqYx8i3aM51sGNcE8ZLaAkJdSh5
q+Coa1Xpbdm8ppc3dVJqDEXJTe48AwI8CsCpHdBaixjTZKOjb3xBm4xg1tIdP7G/
H8EQXY7Wwtr10CXV9F0Pr1zE5EWv/IC+lw08pn2O/FFz98r0j68P2KXH/yJEJAfX
+vFmFWlylnDnMRIsFMdoJ83oyT7RsJe0gic+VNtq8YnsuKQKprOE9hmhRX7n7pKK
MyLsSRIcn3ufs18kBLcX0Oog/0zODkP6K7MKAQau1iD/6Vveuf3z3PsxPU2lxBd2
5hQ5N9zTAvZAXg4tvzWppm1UyseGfBYbdS3QdxBM487MOeqh8i+wUvsBCG6Hr8AV
yhXuuwN2EJCO3LQgZSlilr3dsNx0ZNUI0CHPYAp+5Sj+5ClHg5m7tATqQkvJN5pV
a2uNh4tHB/FFQ1CYY7UvMjPBiQJH9hlakHfh4qPgMlHVLRtEhoxvDXv9qx0ghNal
YtRy/S7DNTfpuhXucG//pAUY0qkq3HLiZ5mkBbpwkQQ9kX0xaCLERnigFXIp/hyU
bBZWBpb66rZEhNDFepRg2giCsCmB/BcuRUuqecMulE+69UAEcLa8URI7PTxXvPBo
RdL6QsDVRZbsxPi5Olm/UvtqrY9hOFIj79AeE418JKnPz+GC6xFI6O2nQ1tmSJBh
VRw8n3zX12tISJ0f4qS2YSjyfAY7FZbhBd0o4PwPGFNpGj753RTn1c1iD+5uhGwQ
dbmzUxQLVOwJUYx7s4cgIiaYouYXpCHDrusihHbOHnQ3r0uN8ojZXQz1PCLLlopW
7DfQif08GOI9vPH3IbfWwnvxJZh8jhmrXwdrLjFLcWu04OU5QdJLthgOBQyaCyza
m2QWWylMmCLdtDDsyGRFYuFYgsoWtHEg2QaRPfiPSsFe4ydeP1fmER4fCXYsZ9FS
6GEvR8WvBXRzVg3CMfUZX9xs6EFTugxfzB2lmBKFdfIgCq+UBymlvr0JuDfeIyKI
coPjsn+P5bNNqIzIht64MnN6h+R+Zm8OsvmtLlyxi3oX170cqpg0xRmxLxdSniEW
26zteaiGY2cC4WCN6fKHPYhWDHJlMfFlwC802i3bdRQbnbLz9RU+lUTqmTe82oju
bRHGY/ywRDq11C10M5w3OFfSm3ZtLCG4QptUY5R18p9fpmwGpyDPoklC5LpZZeK5
e0Hc4Fk/aBZ8jKTbO2zbI2MMXvZ0Ph/cW7ZgPRXMvDeslENOut1Uul3JXxiyPEwA
MsY9hAdteXhKYHBumpop7p7HXhIQpdMow5csxOk/j02ZrMQQpT1+4B10upqLJeSI
JDRQte3Wx1Mchf/rZg7LyhQKYp4HMKs/YYu8RO2Yom1Z5SUDSTgvKOO1uuyTiNfg
E2KW9DPuiILcMY2zF9hoOkw+1ow79ZG2imka7GDj+sRjQbN6X0g6bo2WvV84wL7o
JIhJ0miecQN/kwqiCTWp4ZUZE10QrkLaydJdrFjbX2i40tyEP/vWdtgga5j0aEWd
G7+Cm10o9Rlp8MrW0uwQD8R3LXPZ6RCgmTdYSQOiJma+2bh2nZvxKi0ulZErvfUs
tw/GDJDunpwsCJfbkG2D/w6SUsqpEfNqZQRy6gBrsj9gczvAX53S4Dki/HrmAS0b
UwDnBWUHGvLzED7bgf4Vvr7Ogouo0NIMTZZI2F6BqqREWVasjKxwViqg0BCZlYAE
ZQgWUHvsd0bHY9XczcYKwg5wfiRmycQH+4CNXQw/+ePuPS6v+l1pHgO+Y2x4UzMq
emjL6dezcACK4j64vKMVGtI1GNWAaFQrm7WaO0QcgO1LXpFqKT2nt/VL1EOSt9GW
8cTegmDQQhOlhEr7EosyD80hGIgv/wqMAKXyfmLvowslhxStJuL7VizANmJKsWZK
jPsmgI127Bq62PO1Va+Wm4qQo8Q+fcFQgGh9QC0QkYwfzmX1eHtDlhtSBNOsZa/g
mqERgs3hK2UflpAvYoYeQIQr8EaoIfxglBK/fClDjcm8xrc+OnsiC4QpKtXjCHaw
5rnJcvyN1CPle421MqzRs8za5ejXd0R+uO62FUxP/tqe9JSSmNBi86Ntl5yrnicd
TTFg2s+VMDEjE6dg/VZN3Qn3yeglCVh4BiuskBO/POUofAYsyicEKngYf/oofWLl
a6HwpncVxEjDydo6KSVOrQjf10T6p1bppyPKEKmOrNK7GwTFkHdArwpthquxxvcA
A6x6W6ZRnt3y8w9SfZCp/uB4bZEOf5KqYdrfwiRF1M3QctSjRDC6180GZD8MtLeS
P5OEK1wpFKCUN39MTTHmbrLyd6sS9HC65xqMd4vDEHvzK5YyWP57RgqXnUYEWQvB
AJwsWw71y+OvfrVI+1gQxOZJQjgDoqIbRANVgfP0ixQCBFmt2F3aRX6VjP2khJgU
j2VOoWFLf3BYOtIvVs0CHZUJO/NiRbWytu3y8LkEX5fsU3ha+SpPPP9bLB4bUTOq
RCthqEL+8Mhpbv92P05sfevDdsef+hGf92DeoaTb3L5GhG3fWm2XX2dA7lKDCD8d
EUUoD43XLEqGwRucIlht+NPv0kgKi9/Clo16w7MKW1LZC6DipF/hzkgPwWhYGbh2
oRLhk9i1WF99m1Ayyo5/cd4VuzXybx6ZlyEOmh42hKJGF16bt12hwPUM/C0Q2VX0
A2PUQ9iKIVHrArHQR4T4FsLIKeIatMImUjAn5kPFUVKFpNtA4NUkhw+8KsIPiHPi
tsXj7tD8FuoVUv2pS9RNAFYp6MRh6Jt2GnDw5Dz4+tXqSzqwDIf+E8AjV4iR3/EC
JEfV4RNjPB7RH84DYKBOCn9bIMNFQzwTTkEoR+0+SPZwI4O0SZ51vjTAI68J4jve
E17IYDThDb8Zm+gEwwRgQ1WIHV0dx4yz7NZDRaejFo+p68+Kyu/Umi7W07nuOtmn
12Owd1gSQtWf99uMoDneIRoczKTvfYYMRzmYz/81QzxFsRRL/nWARtJDi2LMA/Z4
gx7Ih1Z2LlSjt8Z9F6EvqqlgRVaJq63w2VBmeMFRgStFJob7dwDGRhcFbcGkFBG5
yrfsWjUZxoFFfcyZ/KdF46mG1u+AOGco3wL36/defNgIgRHtTH9oZGe5cSr+BDlc
w64Z2G6Bx5J54N3izuJwEx9oDNkukrBB+6w+rpY26+XHUllcwRTIv+WGeWRq/vL+
/NFj022wjruualqeGDfijFDoatoNcx3EFlt+ANCCeUu0EWDPYSMMEpcBjL/o6rEe
J1iB2afTjYYGm2MqL1+P2FqJisBpZugqH0QZFoHiGQhKx2HEp5etdFIh84roUy2Y
m6NM46a/94zC5luQ1wWhNkBFcA8+3gb2Lg74NVFLMyQ+OUM+5et2Vbp1MvfBR4nr
SpsDBBoOqnzahOgd9bKAHig8iqjCnS3uZKHysJCg4iL/mghf6S5tlSkU2lsxXjd5
mU+WlWHatc0fDxy4TWcRDibzn7aALdlep2g3gYCEwclP/Fda/HCAxp3y3slCX9vh
8qtbwUMz4wrAM8WAlqK/MoQSMFYv/1Y0iOPGMm22H7Hr8bzV0tpoK6a4B7yXWI5c
RcWnrxHZa5DO7CI19nIOSrF8TutbtLYGvxfR+vHnPaS8SBvyYVUuMxKE3tA4l7Qn
dMj3xAsr1y2PbE7Qn/1UU8R8i40dLcGAbGqfPYZ8MVAER133qHEptQ7yU5DD12OZ
LEFtZKdgv6LykJjs9peVeYWw+yBCASU4AsLLL3d9LKp7cMADvwL0Jyi2QUZn6DW3
WEd7lelcAf3AJDRGjl0XdEl4qf07NcCzP4vmijFw6OLR3EJIfeEYkboXimsre6Ux
e3xZ5eNkNTFz8x67CWzzx0/sp/9OZPFoPzXh6YPe2U7p72aHCaNU0X/fKVjvBnpj
Uoyofy9UfbZ67M4xbBrkNjnmXwJUCNgggdOi/tbz037Rm6lUrNP+w70C30P0uwu+
RmnsWXwhEVLlZWu70bwbNLXhW4bxlgIKBBr/oHm5gN4E6MVOwMp9/7giznPXB+bq
q1GaJ+L1Y+pbYiISgTNbTRwMfsK5CAiUXsfWJhr2DwDun7Zs5cUVAImwyf7H2sdw
kAp9TKnKL83r2QWwDcScp20e63MbqPx5OGt5EfxixnUM+eqXWcwfoofq6qISsd4/
Mz+4gumrREN/60qPRBWxuuqf64qIC/WxmJSgoQThGX/Isqzt9DXQl1a8+E4foOwh
hrNa9O7IyEc00eWIe7nN2CBJHQiBWrgxQcqrwfNGQD/JX1NDxuDc/vVSlWjFB3zr
McGnSkNs6pnug1ytrYSOxuGmLIfhj/TdM64eL0Wu3hSp+9EGQWORj7wsWF2VxmhY
QreXjTsKKYoJnoMrHqsuk+yQ25hEsduJiKan4TEGSR8ha6hrdXpqn8WmuAnFRS8p
0w4Felw9MBIqcGMQ4tSGYCr2DmoZ9hSL6cBQj63+o1Lfv1lX0ySM0gag/eOw3rt7
KLPHGUNiHW4WN5K+EnGfp8zOhX/1u1TAQ+LysTLWy0/LVZCuWJVvCtA9VfvkzL2W
Psk0+xI3aQSoNQlHo+dwVX0A8Uxd2PgRfPRplw5Zmr/nF8JqnWffhZ3B8i25SriW
AaE9w9lt5zI4D2tSsodtUrs17bsA32Lh5CvgQ95uZzbgKO+WFWWxPDflE/1M0Pe1
BumShwlm0+z11iHbwb8ULgLnlStCx1r4aw6eIvBrG8hGJUnhSEQAoZQWL5+2xsQ4
f+LHkUHXy2SNWLFyj2Yk2ayXSJJbqDoKWwiN4K0cR/q4kAYqs6Vck3k13VtXmj6X
cg4Om10mwwqczD0WrBqwaKD73cfHLw0JbjXt4qtNfWRTJhfxWWmjDLokmb0eip8P
70Q6dSAfh4InYWGkZthCigHO92pKyL6u8FD59yS11RhQadZtMZeapXSdbOOEqLQC
rLsfXca/KLKUF7dO94rwc6td/3vDWb1rrWkeNwLhHRBCw1b7//ejibNagjvVZSff
NetxSTysQzsN+EkSzAj0PSzYd0AMu7kWTzPpF+TDIE9WeDPBqVOUAvAhn8lnZ/7J
TTpTsUi/VZtHyzGP9SlOsXYJgb2wQQCjOmrkhFlFUcyQxfdfZYypi6XtIvuJwbtV
xlWBb9dMo+jFRrTDgEE4mLxeahf2hZbNwalku/bxx18+iVdfVl5Xl7+KWG5kfziM
VOrh2mev8cc64ksgEbmFSZcPhmxHObX5aoBRj6FuULfvcEGK4jCG2op5QNlCBIYu
WcAtL3Q5rGplF8KMdW8D3dOib+LmMaL7uydRez3CSRp4ciFrEwIb1Hjxs8JQb3rC
PtqXFICM/yNG5RHdVpHk7XcT3Qclfdc2IBjdnVv6/N9d+CYFkWxjmhbzx1dvGGTH
G+Jag69Q1k2k2qpOb3DZdW/nfS0CY7ilYgW2oxHV2hUZh/On+Pzc43F3iWVJAZyf
QGmoR2fyp389nddoPdHPanepj0X1EDVHD0ukE2/z1DjHMgDXOAHJ+AHTabuoBZDb
Ho8J8WI5fvxp8OoTdP6K9if+mB9vqO0ApjvQi2Ae/t9Yaf00nXt6vI6Hq3MHWDef
L264eVj4DcNBwEfzGWGgDZkVjU6GgCyUEX4sDHmeFi7jhhtIz2S2o2PW1uPnjzeq
FbV2N5qtErwS3Obsupo/iC3+E6bB/R6kpDOfUEMOtVDjrnR1iT9Fmj0Q4KLZdOc/
CyXtqrp0odjxAvEJyG/gdcQjpm6Cbz7kpLzT2TI6kCP8OCcRPbUaOpUSXUj4f8b7
xnyLgOwCBKWyhqXi7kAogbj0HjN5rgGd2GD3xbmSlJKPXzxDjJJq0PjYSpdIpZ+C
qgx2ZXrHdrMQfjM3nfE3RyUF0UnXLS5CnhNRxNtuAiNI7RyPpzQD/4Tp4JZC3xxY
+0kFuQpYPSRYrPxpKzYQtECr4QvOGQb7swHCHBVLx9nJlQrbxFZZ61TtleFCxN2N
6f9ZKsB5kQ81CNjDKDvaddfTrmH2N3TL8TItFoC2wX5iWcziAqQAQ9LKEJruwsgs
dNoiBHkySYQdwllUuzBYdXFOAZADxvI0gtvR6/n7lpR0pm+Gd85nfv6AHIHBqlna
DtEN0sKIhjx0LmlEKNs8uXCOIhC/meagvESTSzpKrJNKf+ompfSNrtEa++LzHmOU
pLGvpLtlOJnVA0Rh5/0CMHR9yK/CXAgdl8BhvuiorzxdrlU23o5UKcm5wq74n+9i
lSQOewLjK5glMaSma2qZWvt3Ruue+CH2iPcbg/y9EOWXdJdTXIXYk1UO9z4ENMHw
2exg2HQxZfehTi3k+1G/LuXpgW2h5z+fst/Kv6e1N0WjQsdzY9VktD92Xjc7nBmJ
1T0jW/W7dC0AzvEfwHE3g6lOvhaGY0lKFxzbCjFIxfj+UTXu/ufgfophjb6bjwef
QPYJr90hYvKJ6ryfXvPYHn0sZ5HC4YCNvQmaxxC/d6m+31MGs06+9jkLBOmypVKY
xTFmlCytN2NHL5PrjFegi2gVnRMTgXZoxG+lg8FNcNwRiHKxGNwlH4bRbJOElbnt
Q3rdRMV/XaOYBcgWn4mVOG9wW7fJLRtCg0JoDsd2Oje2sgPJuZA4T1A9ZUUnAo1n
gCdui4HYQO8Lk0r6yWGvGXFAjEalQX1UbcpZOvQQA+OvJk7KLX9XvQn0TCy1Endb
ZBw+fHpvYE3Wn86C/XR34+5EYNF/Do2cmyec2mJt3Uw2mEXY+qnVJZV0gyrIou4r
dAnj6eAOZ+HLsOXqpwIT3oKl0WM4kSbVVVS7yJVPtL+ldyndO+1vFh/zzvSqsFAe
ptzL2F9gs3sUZQVaODxa4iqHgFxBFSQ8zqw1//xR/aZR9GyN+GL1KWgdEKq8V61z
1XXIaQv+cIxueqD36gNnYsBoEpu8+CRkPH4eGjl4aeftTu3wElVOwEeebUVeMG0q
2flwRU8pJd1gAiCHeFB/Kh5UMIgnafN9Rqgs3cUU0qBhtcuGnadyLyhtqLnfn/Uy
RmsyP7VJZwyiR2EnNAw2r9yT1td/kQqW+ZyLBIyuR+ENVUjYxvrFAqd4j03FrKIN
pYHtuKEAf0GR5tgvcd367M/opOMMPZOB+RYI1FyfZzpgSzZZI8zEQHiafeCG5yFh
nZiEEWCb9xe9+YMyVq2bcRiWSZ5lPAK1PL9fLapg4T8+CKZAKsVI3sxUAnY/6uEj
6lwlXmh3Hw9l9hyArfRZSaY5ihALv9B/NHRdYznR8A//sZJQMsA4wJ4GYYXHKC/u
9yB+W3eZs6wcPbd3Xcw90lKAX6cWmI+zoXhb3IANiGvvMOZSgqNZmgAkm3znKnO3
vuvtGIiSsCeInQZfA9sNXX1n/w+lcW2fPWXl8SqD+aZMTL+fjbZtx/mRay3nLty6
61GCbyXKXr7AUWHGvbrvuncMGM2Ml4lPpS0ltd60kOE8EzE+x2XaWOlOxj4h6gze
N3mG6o1Gr1ALmVepWkZ+6vniIUXsxVbrH6YWbItxiafiTh/Md+Xj0J9ebCQxuu1L
5dkkn1m9R1om22sqHfwg/sncHHmdhDYIAAG1j19beCfibRYhJDauMzvg1O+rU1at
x1sk5EvrAfMlMfflqE15NFQ4kpubZ+IcLOXZvWoXo6EWIll8XvTW8qwMfyFMSmOB
1iRTk8ybtNsu65uZVilT9BgALsszXW6wHx/b/Wy5rT3Dfqe8KzcEP/6YJfZP1KpY
fNRN2Q4pnKQm5joagJFAlNx/kjN6xwTmHpZ66XxqAOFuL35MDc+nlQG+gI2FB8U7
wLjXEDJo1vc7o/KznH1iH5uofGMduqlIiUg1N2aan9taEsX9/ntlQ79xJBBOkAih
Awjz7iPO2ID1LB53L9gKf9TTNgTqaa/U3XBm1lajqaLfjLDzAAA4wC0GsXfKkLiU
jX3/pCq+5PWRCnFhB3LmVUO0SJQ1pPyUbJ/ad+O6kZQZfm+ZrNbiN2eLy/PsrDMK
bNlPqJjWo/MypS/u1bkCyVJHenplZGVF99maUr573HgM/592fLHfSuOB5o1fypYe
QQvsV2OEEfoeioNbqw2WYnhGMzn8imHULOScvdr5WteE03vUBLhP6LxjnWwVzs/J
bTOxU6wCcad7NEp2UhZBtMm1W+LtIhIvnu1Wp9bSTUdL1la9JuPAwXGXsP68Zk1A
I6N7JOW0qASzYDagO7P/lwhCV8C6rH3HHX+F0Lex+ITt1i47m6UnuH4d47T3t1KC
ZZBp6Z3k7pKCR8+Cu6nztuhBuSewoc/5SkwqUzJtUFz11bpw+exNn31YbemzpRvb
tM7NSKANfafIU7OPa5N/BHi2civOqSIOaV+R9MAlAZ0QPE9C/oy7lCiJGPOeXrco
k4lBeJtRWcWOuTUCfH7gmYmQmGYbRFMAa8+x1qxtF7xnkCTdaBeuFwkHfIPkepmM
nX/Q/2BGIKelBwxesiCL6kfBX3Nts8d2RzODGE48r8Xu6xTl2B0IjFdA87+JHEO2
FasKIaOMPv78VeomSNKjGANGNPk9+7QXHYd9YWsXlqn8+/jFpU8xZL7OwY7Ijdcb
UgQWmB9R3/9oFWTC2Qg7dw/Us45VcBkYfOL3lvxyIzj8sBDYNCeiKFaSntqwucgb
QYZlY2QmhEmhedmp7uYFFeKgYE9MTS/d6y7U+9ZYGT7bmGUGFmn8JT2CUbyA/g1q
0QsedoB2UU8Po+4/tMeUPerU3U2f7vMvnpy1TBOkH6RGg2BSzMaRWraIDDVRRxmG
L5vm69VSpIPDY6raHD9BO88PhugsfC64dmBIMclcdCPIHJvqetcNIqQ/GsQRJ4nB
Jt5IZ0Uv78kB89NEePNwTGjxWBqC/ITwlDTyTc95C8L2p9wY6JGlf52/AYvV2fKp
0tyGPiD9p2xiiyqFiVdllibGJttyUHRjBzdWwrthlQwU44z+XUUJKWDso9uJw5Tq
Vd9Q9pZY66NM7utveea9PkqrUfbqj+GImUjG4S3Lktlp/1IfPQPBMtCPVHnZU25Z
+1ur/nBmnfZJhfBUSfEozhSsmUrp7hxTIae+h7wpCh8fKBVPRIV+YXoN1ZYU70HU
OnxgrwRInpbSOL9PR3dKusu+SySNUCYH+ioFKtPMaH6HTpiJkO5WguPbubawklrH
R9SrI+JfUF9oF+5PdedEStLrFy43WWrFWRdnV9t/NBDFzg0FLyqeNrSkyQcjy2wm
FIbQ6w6Bjy7dDwCjNSXUEMTwE64cgYYOHm4INy3Gx+UGvA6P7tX2AQ73ke7/LnIN
p2O5ENr5SZ1OgPlLbcPvyMM5ZRHLzOrV65uNUeFk2fY3SaEQdVgIlgvQC9n1o1r0
5YjwHTYYggz96bIrrcipQTQvEZz4x8dvCOf5KOH+zyDrsnoJFMcRCNIwAonvYsXZ
mfrbISWeWtSRBp0c3f4Uzffp64+0ZFcWCLJAwraMQTBbWcOwxiFRo+Z+3ICM+lQW
OMlXBTFe7DwdU6BqLzx6v9bLnTfWttkMWy2o6kS3ovMLbULUrqa97ImmKFqKhg61
0k42WX3QAKk5ZYR4E2oiLLEDB3FS5UO58zYRFwx43GaukytTers0meCboG4D6tCr
SkwrJp/cB5l8rG35FjeMgnUDsZ+pvztHAvvgbJVPWfBK7MQnw5nXGe4JFAt1vWKQ
ppjwuSK272oDsqbw3C1vzdEWJADZyn6ocvaBFdjKO/NF0ZDda7EYBueDp81jl/fC
hmTBUKqP4/cPADODv2gCY2GW6ma8NDCtGkjkQ04JpixgKAKULALr1c5HlaxgT5sO
MEsXlpuY11/L8TzOoXpWD1U7UYTGOGMlPevTO50GB+90eY75tPOTrc4grbrlePEW
+V6Pn/yYkxCrDD/2qYegDV7R+hasHFuaPdePY2OhCF1jq27emxPPvU1i+qp7UYV9
GUtRB/XTUOnrqtDlwRnYUh+AHSJI8Mi0X+O+7k4Wj94WaquZezlfjh8mgWBXtLLv
bUYtPSUHqr4Ml3rMzcoum7GP0LVHASwN62yjNaDUxkK7btZncWyY7mf/m2CoeCBD
aL3ytazjGySP9w2hqt1A36yWnbMPNACav5/2U13eUOYJ52nX+Yn2lTuiGMnj7mvM
g8pKq4uzZ2U+1qSRxjzzmjpvaViB6AKLatuhPyOhvMUlqvBd+oc7GT/AyE9uBO/d
cck1n3I0u/783wFV9WyN9dsFSAEt6RX7mUg9+Zu5b7HXE8Z54Tzp0x6zGB2cp6ak
bIVkf1vAZ7JTurKK61nrUf2cUwZ0SX9dwlVDjCNP+AtCy3mxslNViV92u0Bv8OyX
drVDkwR5eZ6ipHOyox4e8sA1aVACrKePz7MBBobcHXYb5eGQA6vOau8FqkCoQul4
u2zr5smBm+5X8D2GBw2Oa0H5+0ES4DNvesKOmOcjI3gVD6/rwlzl0GDHGMpC1GGs
TF+WJqRtXcQljAfg8m0AbRH37qe478G2t3W6kK5J7JURFXYwUlwErexCXcolggHn
knaPpn85b1WAvfxGWYnFtsbLm+kmYB8VTiU7a7Gq4jnQWFKoH7ZWPyd3nOutJFCQ
dBLoXs1s5oLHhPkB1bo4sFeHoBoyJ6bciGWECRscMPRo36eoNR76VWUjslzb9siR
wZPipkJKyW5ZI3kSnorWv32J9FxGx7Xboo5o6VaGkcQzhQD6x18O2Ntabsje8h6b
TlMO9Mkf4ou5Qy+sqvnShwPivyKUU0h3m4qYqH1xqoEaKWGfaIDZDi9+0sBfSxLi
jBoLY3gQ3b0RVEDPLot6l7Ku58Lts9/WzpZwHCJ4b0l69siVTYSnVRK24tOCMgSJ
BIQACTBPet4QrkRCT+T3zkspJdbt5v1n0MnMaj+VR+FSInf079VejJJDCDAxsGtN
NELexVQhS/ofFWfq8r1s5e3Nv4ELMIc1RWwBJtdVzjMmquddDrySGmYXR8QQX2v9
BrbbfoZ7KTl04PRPjCKdjuEhD7x610NrkhQcgBDLuH6REdDr8Upd0dNmBnYiYAO3
9+SjQ4lS+5ZDylBKayUzHViJDp03S9KssqizPDwLlMO64b/6n7GJfHAxVyY9vdKl
yC0IAxHQ9MvXWX+c/BgNo9/ep4ZRk0yjMWbiFjr4Z77PNa9uL8Gx5L58eOyZVUZy
x0y/xciZo57lPA/3uTINltMXxgkimFlswYU/+wd/+higtyOBG/hNBpFgYPdNWVh0
6HAdwiUWMaUZ7bSQ8GzgjLWQswXXiciyUptGwacjFwd4hrZBip/qdv1NfOv4aSsM
LOZk1TcrghT6Ft57LlGNXH3lmLqntqZ0kHuZ5whoBtO4sG8GXeq5YNz6O06S1S4R
NG1Dpcx2GL02ecmNTex2Y9A+IjpZv09MDhU9Emwxhuw6H8jX6yXppkdvfSyPxoKq
f0cAj7M6fltbh0GAbeIrHeIkz+lic2E2rWOCGW5Rbvxgaz/DtSUd/37KDJslxaje
0qOw06SJD2F8JYaimjKdQKa3P0jUNz5My9ljSQUD2olJlkrlIEANAQ2Bq6Mw4V6o
c6gQO2IjMFzloyvfcfPA3VbH4vakW9a3tGBiITwwE/NN92BgQEZQN+s+a3ehOAQl
qYhvQhH581yutIBkCd6x71o+sONeEhy6GbKhiT6pvgGLFFzj8rHjFamTHhNpHoR+
kNrM8gZe4/RfZJ278qpjVuivG+3WpBbd/Rf0Hp52FAC1V3CEASrqSArpFbYTkjpK
iAc152n70BfHbzxRcNMytKPa2xUFEj31XfLfzU4LyIxhvLaGjUbhVPzBVgK0GXCH
jjTQGfQE7mhVY2QgmuqxAJhlv9aP+5ckysxJVJADCTyAJRVDPQGeihcTH4ro/WW4
QLlS9KWY1ehUcZI9M5u1OB/4oVJEj5bdpzuOH7gGgK98fIeYsKLxf8zkXqk2zg2x
ktNhF9ee/V8ROAJlViOYkgRbg8R06nRtoJlclxKKYx/KzmBbvuij0tCl5hcijwch
BTDtcAwFbnPlsX4e3UF5cLGkbjUiwOeWxr66jm2L2wrKwmGZHPJBXl3HWr2wHiqv
G+PqaBLOwcuA3lfhysTPSPIyqHeHK7FmJUEw9/UuKiD7z3aGSZM0vkSzI+6RZNA5
E/IkTz9RKBxMTMEj4+nlJOojLN6NQzLjeGZnjpElVbEus33/484tqawzu2a0IFdD
HyE7vOhQDsGOK202e1o9c1zFvMTX+oUGForDCvFJ1f4WIapqQufyBIlHIZTudEw3
r9D+SxDO/MqdmSXj+pbgpZaMzyDOClcx/SFTeDbhEshkjTSz3xkLkdQJQC9IBkHh
zObBEofWHgcS+oyuoQGiHIHQ9D8f4X/cdtuwtzRrsKk9YxPund8oU54eLbMCHlkl
LNZn/p7B1RXBKmS1uTwI3UgTEJCJbZ7K0FiWCoB5U5v232hU6ZsBCVh9NhtV1aYQ
ZlPRz8AqLHikm9KccIhS0Pb0mGCjcphXIcuQ8oCsbtsLXHvxvl+z4VnoBDVKApm+
eZ9kzWhYFAeP99DZtUruwfzUcj6FlXZ/VGo2Tuc83MyK73p7pmyJn4EuKed2B6fH
YiSNgh5kyRt1ccOHKuLQ9JISJSZ+9Om9VcJ4YIPIJnnrFgmMRHtVx7uk4Gx9a0fa
yxuAXITNr47/FJsg6VRKRkh/5YTEvMx51OOuUMokhGtf9tZvBaSis5vwTXAWBcCQ
jfyQJ9+0bT59s4ZKyp40bstbr1ylQy6QoFYCj7b8anfVUodv2U5EuHYUEt1SYASF
IXFeqgNd0miBjBG8TV89mV4BD06lgKC1z74fsT22JAfZTF8tXc857xKvDqo7Zfum
7ncKvbpgQkdDvJAae1tBAhD+YqWdcJeXMlKv01+UEgLNHb00Asxyqr0oq6/IkaWg
wGnCXyfCO9o4FcqgRht2J2RSGBCrg+SFalZsGDVaaGqI1xpWeOHq/u35vZtSV/ig
/8pfnezKxK0BtvdivpfvXrxrj0sYWjz5IaGcC3kQI3tUF99LEle9K8Erw45NKin7
9lEh7zCotvEXArlLn5xjbG5/RNzBDESe05n+H7R5J8yFS/xUvbKIElYoj8UD9uLI
PORCtAbSuA5nNlLjVBB9cIUpftXNourxuVFFdR1aCBxWF/IVYt0gGjTlMUGUZLO3
3IX20W1SifaiAG3KiMiYSLdCNWoFR3YDpPeNAAUV9ePPXr7QaEaxI5WP/fJ0oPmT
qT47D6ksfHIib1utmDEumBKUHnfw0P1qjrusHWhbV0uHfeqo1exty+W7qUlFJAj1
SY7JI60o6IAC76QKOxt+x992NXyk0xoWC4wHA0OyJP+vLDGJdWd3vYSThi9d8DP2
m/r066AOsUo+pejQFguwMP83Uwh98q5kWDtqJOln1f/afovjbnloDmmt4HBlyoTG
4NaZLWxIwmP/gFB4NjOX8kPazhP5HwQdVyPD3KYPKq6M9BxmTf4proatd/G+o/J+
lay8cMn8M3LJEjaUchKiuNZDppUZt4IJbGAhXYPEwwdWPy5GwqcXmOCskp++WbiB
r68TnhONTDZxBlseFQdTUyTYJHWZ/h/UU4yt+G1FwUbX2d0A14PI6IZU7xgntuUh
byXkSPMvdl3V4s42YN+OXUu2TTE8wBrsa0NwOrQXI0CX+NdKvuKjr8kxELOT5HAG
FPfP4na1zBG02TvrqBPb/bmTe4FBa6ffLJHz+3WyQUAXAeGoUrqMCWRJCVUOMkht
mOcL863U2A8lS6bTw3227YvBS2VG8LfIjWFU6fenT9iHo7iTSx7Jqkp5UD+0v16m
obwUgiU7deh2FO3wu3oAnLT/+TaNchhYU4E9rhfpgL5tvSAolDpU6yjDK6fD3e8t
AhhKPiJKM26KYFwd2t8ij34e9X0+OBlrKY3u4BNM6Ig2CSUlYrDIhe/XtPihPoy/
j3YAI1Bn1s+UswkycRU4OUb/dbcgndCCqpYpp6VGkWwXKpUjlC5B1oMv8RoHiSmf
zxe0IIXdSbTidGaIHEVotSFzqTpClAzvtT8lv2HSdNVX0rMJySPqhvcArABlfZ8e
8N+sknH4MmuEOR4YIy9walE7MaBl8Cyp+ANhb8ncyGoIsg8AtTFKvDTO38ldPYr4
d2FOTXMcomBC0o7zcL0K1mnBInsysG0EM9a7O+ok+ecSXHIzvwa6YxHIzuOduvId
XBMj4rF08BdnwKQKuhpheX7MbaTOKfDuRqd+2tJdj6MHHCBsppkMvsc9Qnj/Mt/Q
2cboUNgKypv2REVPh+P5FhEXTsucKbc1+nWfrQEQf8nly6AXwgrVYZGfHxeKEyXc
BF94UMLM5ZiH5gxRdePJmGw4R75DC33Ws/sk30bi2BJApBhYKI43vfYlGDKJPhA7
65KbNMDVD6vNuNg1nP4oZg6CLfgKpHnmAEhaVATQukCItISAqXLQnnMeLY3yvCnr
mj7ClG4udAqV46eoF3Y9/A7CXW0I7sv7M6W/bGGN4ZpHGlBVcc5kfKqYxMkRxO0c
O3WspX2xDfbz939S8eZYWrbYVnfV/ALCxAYR5ZVa8+h48icwUPN4aYxu8RZEcEgH
rIpi5xw48wqA15y7/H3nKzNETdv3omVSU7V3Fp3fe7viHu3cOVfVeEhPcfoccRik
I+/34gcb/v2tDrQUuRR19d3THaOMJ39juxLYNTnXkXwY8fkuB4g6SK2/ZSSDEnDW
pbrFfiQl/0DzhMEHSsRFvYJhsQzMExpDNig4ORY4Thv6wq0kCS1iUspl5AVY+zV9
9D8hARFEDmqaVvEl1/QiRXEiMq32U4JGdiUPXDDFaMJZz+HiBv6AaksQJ6CZjGtx
AdRXTdXHZsAAZL/wH1Ef2tMEPmDjl3eqOyfjrCJyrs3Ot8ateBnW6yoSp4YnepAD
PCl2THjC0//jQiu4Shr7AdXyF2rlLHJR8PbU9TWzyKP4T77twf6x0ExjzT5a6bl/
/PIzOxk3g0Z1kw9PCOIcCp/lwqoMVmycD/94+vz7oJp7htL8DSA6qllNgu7v4zOS
Omlo870LGeugkjPbUtZcY0IlvKH1ByR4pFLE+HHpYNB0+ySuJPRqCDUeNSrv0qLm
HTZ2wQMlJ44l6WBkARnV+nmenOz7nkIoUOH+1ObZ2i5WiwRDuf30qLYPuBFgMGzB
QBMHQkEakDCbf2ygf4URMY3jBR+fNnzpfe8pzcqJcVMt/JMtqL0lG24inOnYeqVe
Z+aIORyccvYn3SouAnmDO5416iDDc7M5QqXRFM7oHuHh6WU0ccAtoeo7fvjfyo1U
ZLrc+y+rZb31oGxETrzSrc14BmcVYdAgEyw0od8pl8csPDCzsOBKwsPjC2JgQwan
ec/c8R5VIpgvRCUvAZNEenk9/YTUimUnaKHDhg3PH7Qyac6a33LlI5zCT8dFUNaj
vinWG9Kh1AsV58z5T11tfKkM8qZEOem876EsuPDa0Cny5LDeRTcAjxTomXDJBGqq
P6UAXXXU9l+WNOBA0c7/+nvDSODR2Gv4AjBRQnfaG9adsH0NV17NXsVId7tApvQ8
HXUPn1al8TYdbXLrRToCn0i43c/YcCqy3kEFDemIQCxLhdQU4I3KSz67x0+NuhMj
AjKm4Z5Xam1AvHeMSaagjJZgN9AWlOJqMCDf2HVL6jEf4bUepx1KuCuOnp5KjDB3
n/DkP99uMsuqqz0eqbluKK+I8PsBovoYvELFLjfx9V8zsJe0koFGQucKKq05CZ6z
2a7f+RW05g3Fx5dbMrYuvf5IUNgNosQAH85c5v6rbO/86UKo3sADlE9UNaasMfmP
mIpYFefLrBWoOhYUpzF04zMuJjwJ3uYzr5cWCgH4amd9z9kP9s3+b6XNwjbAlL3u
z1ctNcPfJDoEkq219OVck1f88LcCGGa2dF25WVX/niUq8xaMU/uhuBewZlxFaUx5
aHjIClUTGZlmWNStUvXzS3MGy6TzXW0ZIs31ZDS9ZLVmhGI5VZTxs6dCdn71GrKc
IUQY9gwrk+eHGBE9CZ4q/bY7RAHW5taA7no48CGCZo2Q613HASAVmT27TF1cmQtM
VMhkDZuuI9E8cniP7Uu9kifyjbeq8DPw/esdiwDt347GnmyXuYsB6uK+wiXSdPFI
b8sbfRjKZmVW4NrG7EOd6xoZ2OtN+UeP26PAJ4RoMDgL71+TX1rqE9pfdLtFS8ck
qEpFGF00HcJutVGwbuiH87V8le0k7SNikMcTO2hNBtJEWCN3x61Fuw3HQ+k5rM59
vLQysM/qaDRl1ndDOQcKM1DfNvTvTIaC2MFFSZXTPDCPAI+bNYgkIsPtx3cEkR/F
1KArnhDZxcQKB4eDJV7TFJ+yaf7cumvuYHuH0lU+QNmP//0sA5xQYuVvkjYv5rkM
ub0XL2detb23rgA0SWq9e/eI2/E6Wg6srWSfIvwxTT0slDsyKXsZym79oWlfnvZE
KEraj07dygUbgFi4ECzKyxLs0ucKZeKYQBJ2aktnEZUJbSEidiuhXtVfWn0pbl8d
eIkl5uaDIrrd2XmQphKFNex2XMhOfSeUXxFogvmb3+LCK/apiMwvCmlKuvimsM0S
JMAAyy+uz/3NMf01vRgfKg5h6O+tp2/fdcT0eL1QhEVb22Jk4plCnDT6JKS++bOT
gLI5FIip5Gjfaad0pCNQFbWFM+0nSbj08M/fFTudgDvL/qdk/hJjpLU7UF60Zzl7
ETAybFYOYeQk8lfiPUNKC74tbysKROiz45sHPTcYMXrtNlVZTRz2I47Bpef7KTPa
a7v9ulaDZ+jTjEpOU+o/mVFTe2q9cx0X2eB/YFl/2Gc7n6omoEnj2MOwvEeMIV5h
BYLom4Wkz3a8NvbVnqUnjAgbmSDqpY5IVyLyqXn/lyQc3ddJqLeIfrGGdlnKa4U6
N1BOXCtJCC3zoTfEniw0d7JRPC+oorasXM4W2hdHG8jWEzNOZTAbKiw4po4P3VkO
f+a4wMrcpBPBZEewqwNs1qHtGHZprhACzytVGHxnzEN7PFaeE6+IUabpRH10OvAl
eCdEIGEPL4v1mJ8gJ1TbhiTfmcc1pBGPKvNh8IJm1shuqMT1tdTZAMb4+YePm/h+
uuKCZNDdCKbiqmONh+0KuAdQVzK2JsIztcQkUvOPww/Wx7JrcdW6iNAJEFwGronh
36vLXTNqG3DL+9OZToJbwcE7stmlDQfRB179qIjjJq6/97Zfp1A27YoJqad1QaFO
zrnmb/0x0YqC7jpuP8Sf9vdlU+bqADBw7X9WItEdzoZDidnlGUNipCAKVy1SGQMu
8JFAEupof7HNyWnKCdC7pn354NIGQHL7CoRUVSkeBCBOMfnufM8IAJo0mMg+sLb2
DLIFA9r/AI2C4apVhWqXbk/GMStJ15Dj6t0ED6bwIz8GFvnSDdsUCjwOiwLcJt1x
kdJy0O6JujjB8BWwULrbGsREM5hmS22GlE6konVg7CYre0GRsylyDueEzqE4hkgV
NjrJZx0XGoouEinsW1/fBN/6H0djQQE3EZQkJyURgK9+VHuuP/eOQj+uC1HRzag6
TPzVO5Phyh+FtIi1jS1gD5IKXWhjqRzGz/KPnNawH8FsFeivwAWRZ4WzJPA6kg95
jXfqsvorLR1VbNt9gMxkvbMhRSiwAVcYwmzrPUPhfROW84QVF1uJW/CYarL9NMtF
3nBIV7MbKwZXhi24jIJsMSTpZHfG1Yi77Vk7v/3Lu/0slR/w3yN9jGM0nkFXfT6W
o30fsiSpWNxMo5dCxw1IvcnJQTMkKovh+0yt63zFbKNYIVTo2LuZ4sAd0kKZcJXH
9Xn+vIaDhFi0MYiXUrvedFWKTNQz21TVi0Vv5hkuOHD8nbOVm2VJwzFMcoF2Icx5
i3/Wqf0Wfx/UzIc0zuCIWtiPmFsoHTRqO2rrm/TkwN2pnE3n7X9ml8fLthv5bET+
b2vqTptWQTSpF5UnUpsH+zvC7eKP0e0PR5DngNl7F2Pxbo7T/6fJCibO+fTP5Cym
DTtEiVEu+cX+5t86s5Lditr8MizZLcZ5/i8OzkmA3Tpym19ye8OL1/cScNwcpOxB
PQRNTgSxJ7QtrtfuXwIefACd0IfDqbrv6iXC70vPs/1nwk9SNvcQnqx4H+MUwkOQ
J659cbd95c5pHWrSNavLh/Tsu2PKQ5FaqHa6mZhBCxahJEAZLfIrEp5/PEjkbrXP
Clcvw2B6UO7bk7snRxWBit18/pCCR3RzNyW9BeBJikPV/8MW0UcU0i9eXMTF02ts
+2SDdAGQYBERBOom/urd4caldSlwjM8LScLrEG2CB/GO8fk9HOkkmsyH4MFPfVKZ
tq+qd+463jhLSGqihXxyLs0OCBkW+5Y/YUGJdajBZSmWeyrR6bnkCVMc8FHoO62o
62WS5Apm+xTQY51kqT3CLRwYEjmBDL3UDmklw2Obw6HVe7c2lmJ1hkLA6rLtCJLb
/wtVImeLsCIqjZsq5FlwMLWjF5x/8xCK+I6++PB8C45UCPsygs3D6Wu3iBGBeWzd
28KqA11YdUSAd6AN+rYKPO9aPcfvLvDjc2gtr3o315H541JLfBkbR1AaqMxEq6sF
SvtJojkcFqSSJZuzmpj5Y9SOhU7QMaGNLJUZ8QSah+J/wsZQcPNCTkuUN8njP72g
2ds/ZwqDdePVKoh9h9jNLvQJylhpDB9EJogMG4nReKKT7HnByksRsVKOqwRS8Fc0
Bwl01JmEykWvOv9lcMxvvVi2oeGcNJ1tqg85YOo/fZlRaFIBKkkw3nQBHyWkg39/
a+pBbVGdvUFR3geY8Zif/tIksjF4hcQeRYPx+AqhP+pBdx6GLmzMOYpb+XV2z8wU
iJXFKe3dLQZy0Npj8qbf4nJ84l0pUi6QcuWcEnvF7krqcVNJYbmviYG77zKnFf9i
HviyHXqEUa2cYv0HLQQqH27j7b/GeUvMHY8iTdi9zJFu9uW+lJLPWnJaIHwjD3BA
zi1ijVTPnthsUSGbrSUR52WMmjlMq93cZF+YDiKoMg7fK3HIPf45DJ6Fl9zNmpet
C+y7kwL6WU8kmuM7P+gXEkGCU/BcgMhrHgKAIw/NnsRsMoIjTdmNPqUlF9cAtnRu
GWNj0jm/z1mCupvU2A6+LYAjhprMUiznF5cT0YVE7Zmue2f32CbDol4Pkv7/AOiC
Kt8hDDT8ysz90OiMziRiZh+bJoxZdWiPsVs2sQs2GfcQWWbN9/3yknUHfO8qdlmg
MAIZHC0At6O59NA2eWG9YMiw+l+mYRu/zurah+DEaGbKHj1jrDec4+CC6D2cLGPP
N+ODUJf2ND5zYnfHyOfubQBbm+Qff18hbFrMAlpBCNKFisfOZVkn/RYRobXlzIjY
sI+wc7iLN1YQ39qAwiOBd/nh6zk52SjJ9n99427z5pCkbFpNJalC+/Ts3wB8AqLS
GH2L7q4MRNbicD/vpQ++fgi31LSX+huk7B5x9aIPs/jRcpRNR8MbMDW9HFsmxLUM
7NKjljNFHUTLcMkPp4D/RtW5g6KEuYCWjvs1cA0XWIVRmbk5W1bnLFFH9QGSpn5n
KvGbNeFK82s8RU8rIpnsKHx1h0dPg/Gg+Q8eFm3LjMc9kl+eKseoltzaBU8lohJD
ygX08PwmuS9ZmC70SBPB1Q6jVgxU8yAVjj4RJLhtn0bWzkB9yoZ6+jtmnPB/1g02
pGNBQ2BQ6yKAkjL9ufH+t+sloP9Sm/QmD/BcIaJCbvzbxESFuBCaCcIXY1VNSnz+
NTqR7WSdLvasAReMj4bZvE4nofkluTcB5lZXk13WuQ2+OqvoD9xg17Pt7eXUWvCj
rK4gxhAG/cajJKLObYwpp+OvsdG4YRAHJEOsJhuvrHbBR8xmXlwQ8H6Vx5Uh+36Z
xgEcWoNFvaE93fSRTP9WQmZNbtbVXsLRZxJrBg1uiUtMvGNA2QAqmnpM74PYc0/T
UaLj8Y9wbPOnNouYxvX2f9Cp5QyYylwCLhciNKPDZwASqSEHCVFnhNrR4eW9h2m4
eOm24VVH4sDJxjyEXGcnS4zpb2a6Y6BHLNrPZVE8Rm1V7WsMxyOCp48p8kfT2CO1
U2EjL5WMhlw4PEvpErVUZsay8Yrvj//uEBQ/VHx81aDlwpmBLgGasmEWVKmSUuZb
Q1csbY3uwT252DLWuC55SEadjAWDbh29RWRrD68Av58jRbfVnSqc6LxsqeQY1iqw
GW25TXnvkZ7mld/izMoL4fJKySKaZuA5ldYvSA5TypMlkZgLJKyrjMRR5nzLS69Z
W7Ww/GQodUlxHoX8yMmw86hzliOZeQj4JAuhvwJU7gBpN0JA2tKecijIwtScYuQp
ginJbn7Kpoj6Hu6TitQDdA2BqfgkefR14TMNNyjBdbEx9e8/xteo8oqRum1Eayvu
PlqtqtZpdHRyCXCkme0+uCMoF3A/iRkhJ7rTDKJGFb9Wh2Gj+kNBcP7+V3+trPeL
ZIRg3/6Z52avWFKlABn3jM3B5/txwBOXpdr4pncWxzwx69H6nxRD69ZdXDxdupOS
lyvi41IMx9fQSTkaEsWG1AbVMp8H9jm9HSHEKwZv9dFluNdJcWbv/PcutEHF19JV
B9+pua+vcKVbGirlBwTjO4Mub3sTMu+EXFTLtOCdm79PmUCOEoG+yYU3T35N+aOf
rRR+4+ceKyN34Q3h02bVZfwx6fTWKo/b5SNdxNq3QHjRn1tEXLdPAR7yxpC7Jn0g
Ozxxr7ZZA8DS18i0gupL/KtMATPMSvLrfYwAw8qSLKXYolRNX4uNm9CVtRO3T6P4
K5ZfHILGti0MUOdprHVXAhAVKlXIbUUxGqwdo9PNoPQnqI4UdOcqwOQO0O63tMrv
qI0851uxXYnTfzIZyp+EIMGYqosrUP1U20VR78kFR9yzhSc6ZvCwM2gO7mhFCLtY
O2Tc/WWPFC/tBugh8VsYsycHlDXD7pofPGI8Fxh11dxIYIIkZ9gZUjk/X/b+54z1
40qefLbqLlUFIhtzVZUnd3yZSOD1lkmwXO9ISK7Of9WgTo6cDiS1ImpXZ435JnXX
C3n9pkrx7r41Q95MutsjUA7MJyFF/kUIqWYqeBBVcIGPY6s4t71vhRtdPN5YLBen
Cih+PwH5xLHT1pSx9ryBVNuk/x4hNrQ3hQ5NaJV891vU2RgIqXaycZ+dfblfiewK
v7uLuxy8uKxIz9Y4a6pjHQ8lHWxD/yODVVp4po9wLpYh3gEa9VHvGpRVESVCQIH0
Xeln13rkshAdSwR+yBXZSC1lnJKxxL88vfvU9QUWuul2E/HRMr90MC3xsBvN1tnb
TJBIysRY/v40/i6R7O1TGNx+9ObHnxMvWsZ85YXR9IDvjIxADeJCvCCtCkzqZfq6
ROa1vOHZoE1mk16423qOuDKJLje/AeFWlxnShteZl1IS7QfPARKn1RCUBHkv3Nu8
SDjidyqRPm4hvRX/LkWclK2rgOgsqdisoW/Q1/BCvsX+QG3A2yIRyMSBS8oC55Si
rp0uAyGyd2eJPhhm6RKZBPzJTHFooF8OYlwMlV6qRUZqjTMgMI0J2UaJcnD6aIiF
Ya0FzkV4qojwzayn6NDnouIiiSaQ0ts9QUgKjpK3Hz1eAPbJ06rVUhpOfsbAv2Hu
6xItzxy+ShUZ0Og/berbJp0meBJwFn2qdN6MrczvrBZX/QEfZG7gZ6K7sHAE6sBM
qODQBlRplaBhXMvwsthViCV9fRbL7mhofhf2Fk/HM6UuRCFHRKZ6+2v7FQ6FVwIM
ONxcVl0Hu7Sv9BTNoiujP6fpTxVueneJ7QOtwRkKyjLKnvI0smre7ZX0e+IKPGB5
m50l4tDd2Yphw9icAI//8YTcd5v71SY9ruuHGLMCTRNp+tbhhibE99YEGwwIh8Tk
2KBQ4ckb0jvDfvwN4y1jO7Hztnl0unXaWXzBhcKoXyIJVIduAJB6EEKPn3yHrcEt
exM7OY0xcZEBzTAtQ6I7/Xhd26qtnCQHbw116rIMUcKSHljVR9nDpFDxQU4srsNp
t+R5qN6dADC15a2FoECkUpr1X4Um0K+xctG3ZC2NPeuaD+cmuL1/+kzIGTn6tbIq
ZHiaclrc5lj1fE+i+hYgVZJ9lzXXGVIIdZY74oyN7szD+YZGgntuX9BDia3H7q33
kPOFSD3PnYZIlN95DFqHKTNrf4+mfr0vpX1RDWOrbH46+wWQykg4zgEcqwz6iiHI
GelcOc246PeTuA9GD4mDWmcIovjsqbSXsi6iFPkcOK7fkm/fdkM3YfHS1gJX3Djc
fSy8HGSGCb/L39PjlMtSwscMgjueOo7wHjvK7JAbFhjtL7ByNabrac3k5Fnv9J7E
KI3pJ186UV2WEYFwVKcSTaUeqocB3GUzKysaK7iUUJAmfZptwmm0MQAl6nNOWXX7
R+FldaQ5NPcv4K2H8f3LtMSaCf0LyD9GviwOaD0mBsWG7Mza5L8OX64YmYvsyfYG
sSFSZpEjE3/l0dT6KO81cgcg82fO8BUxjU7U6TLcWYp6ZuPBPOEf+kSZDu7IE75d
/MZCsWi2KFBj2t9IARWagLYvW1iTz36+RGXDU0McvzKWYWN4ttfdVlIzFNPv+9aS
tWuHKSDLlxa4hl+WYJcxlNGvMsPSJboQkLpcXEPwzuDQAyY2S6qWEE6KsxGJYhBB
gZPmXN48C3wW8TJvRylnUKraqFYwUeRG5yX75p029DV84vm7yyzU5qT50rowm4uT
xSfeN+SCPSgiaY0HXK4N0rRqhsz60rEKSeVlYSZPYsLZTIG/4DoZIwCEPCCjTSpQ
gaKgSAmjKS61LyqkInQOnHlxVPm4zQkgDzBwxYFg+Vdslpaw/tJq1eF/lzi2/Abg
gsJGm/dNMg8H3pbCaL9N6ofzaYjacCx6hcoMyllW3GEz0P0fd+5Z4Se+a7SjszwO
vVnxIyD2QJSFWvwp7Tg3KsQhU3RdBojSabCOPzgwzPa0AbIw5HHPLjMlDF67FAlS
WfmRjAQPv9ZUltycIQkXy7Je+ygDkSaYshGN2v/RX9E/5nV9vvzmFTaDzvRBB2LS
/cn4JIBGUDerz++w9zgW9Ut4aSKXwH9bkOruxCcD3Q5haK88YaMx7iUZUDFUz9ks
TT25F9WzaKWRT9Tjcd8QiFNCMpZFMOFuBHHwFP7+V6umKlzDWLCLqa9LXnoUBnTC
DdZRehbigVzn+uk8xeOO5VKM27q35EGgf7cdMj3jWabvVobW2s8sFdyGwvlfbSt1
IpSSmUK3tkuqlE3R9LkZpS7Nhc6bJVmz2EbM0rhUJxYFOLfRQN84+t3qx9CN4wyE
2o4pfZMCyM/zRYhlp6Rta5ppAtkO0VwLVWFEoxaSvpccYE0JoN35I2A1xpOiaUSb
3LKiNb3kbXTt+FjXM80vBfMUA94mQhfdqsNcPNwPykrU9CRa4OZfyJPgrugv/6mF
57F6YrudqXsB9XlmKPErwh1S0qXSB7HHqtPjisgBf8gI8cxyWllNMXwVGGH/uAJI
+9uxxZdV/nNo4cQGZkBAUt7d4MJn4euhQG33zZHsit83/A4l40Aow5lKz6L27Ehg
47cqFth3BjthPKVEvGKcLJFaaszFlDGPgO7feUVHkHtUi643z1YaR4ODauBwyp/E
jYRGeGZ0EmfkWKOT96ObCoPVXLY9oYnxNx70tppqaBk/kKNNM7ESQrGCBuwLQiJN
iAcKow2tnrJgYdWsyyzLAWz2n+n02RhiXExWml0w4h53+sF40K27Kq6kk8vl9LdT
VmpuuMI7fnLDOioXV3YMSQAzzTI/g96LmDcOJ5d9ES/6imZDe4b6Bm9jicwdOPO8
bA8UcHHY3DVf5zXttugfjU67aKUFNM0wOeB1cxg8Y0r2ez83ijjspRanK+mlfFWK
NF9PlGjlzuK2Myu/x9+fQwz0Sv8nA6NC0ban5+lJtISX0xjwrTtb2Sh9EjCDxR40
iTW5jnRnXJ4P3NvZtm0d9FyGBGRQGb0ws8spdMNt0BZHaK9iS71q77CsCym0Iq6f
DyKxHGY0FPXgHBV6Mky2pv/rh5xSE4i9GEqX3bUl87yBBSCxwZfF8rI7gp43fz9b
zfA7ZIsswRqbsOblgZYpHAi2oDDWdO381VbUHp9rtzb3+bUWz0J/z/85oFcnYWjk
to0YarQqieij07/vSgrjx45N9fjNUlEl2wbBaAViWZ356T/UkYgV/QFOlfRpSuSI
NSqCjnv2QTBfQWmLn8KWMRwGaJ6XMmGjZ1OA0jI2TlRnSi/KM5wARJQjFUCzZcXJ
Gs6VdB0+PZS9wDaAGyj1OuZfL8fD8AAHUUN53ErvB+XiLNfEO3IaIeDbMMe4e7W6
Oyn3vKdN+yLuuGw2VYlID7ABq8ybs1BQy2Ows8sT3fd/bZNa5PEOtAGyP0HLVhYs
pPClF5zFiYWKMFxA5RHCbfKPhm2rGyEBgHcpnBo/v5C+8jxKYJgCIpXsNrUWHEJ/
Sn70X9JKKOmLyNkewIgpLAPF/eTmXNJ/9w/xIMFBJSnPYyBCCJ254SUy7VJqWDBB
0m5J6M1mFdv5UbhBaT4vtuaQqvK+ZrQJOCl4XUiKcfuBe7Ya6h/EI02t3vki9AP0
ZScqyh3T1qyYYAG4EEP3/z66H2LeFmE8ooLJkE1SSm4l4E5C5LaBLrAhL6p8B2mq
QVOxYKEFby1AFNYFf+wzzqHIOYCWRBFWrhKga8x0I6c/DgYGsgRkb47yj0+vdo4f
vF6crTVRjL2G1xV+OgYmK7GeY795hDVqeUA3SmBp/JtLBUfIAjaQ8mEHX7NT/in3
AHE2nkB4VzS8nWjcBaLIdj+ELl7Gv35bOPmZH4T9U5MprU1SjdKxJ7Wc16Ue0mer
aFZz/u9EDc9YwWkXijmw0+C4NPwxZQa9L4LWzA1W7EnJi75vibX0NwVW12dS50ZH
Q130PEc+ZmbEpUZ6rRF7qbHajCj6MNY0XHs0uWYzI9p6Qn0VQVHcdwA1jGjz0LAI
s+5Y1QnhUXzH7gEdaec2WCiH5VDEvbj6WCwrPF9tGDUtX3dH9G39KmQgDBwAHIEQ
zsthHCRMv/0JrctEM9fq50kQRzqMqZMJWUmAoa2YfnMlbuS19sFIj0nocbvQZsVX
FJJ/4gmygY51bUvoVwXkFPBWfVZRlb2y2ACToVvGuPYsNaNTF7bB4xdjsTl1Fg35
v1HPY2GBgO7PDggFsTI5MLuGbdKYpy74npfwqz8FoJZnheLfc/WCxjQnRNQpssLQ
Jsl5SQD6Mf3S6qCGV4Ub0w6FKfCZkdfPsQ8iEaPbSpR4u7fv4vp6VmotDPJ0qaC4
wOItpVleQYimEV00+dwDJCTd4fETiT6dYt18zvF0hFJafVlkZIv6w6pufOzKVHDh
Y1kqH5vwa4BtBBI9NBHwpDxof/0nwxhSWxfbGpwR3KNfdUUtjQ4wXm9XFR8czBLw
i1MNitmUHPDA0liLr+s1kVfgvMQXwazfl8NEdtPKM0RBEOCwS5I0UUEAr6mODPob
vKFVBMwrT8abLCuEjD9wbWohMHEkoCyZymMyGENGZAHlGiJn9vSlhPpUtqWIcg9L
uO33iGcb0eDJQXQ7d8PSNUsfAIvyN3jVdwFYcBsw29A+PEIm9OsUo+IMUNvA0j22
KP40Fgs5nyYLy7LCxAUIc6cSVi21Nfoa/tGqq4+JtTCex8OvEdJkviHKCdcYiwUT
PE/zS6Ioj3dS0DgdgZfc0Miqc/Smq5aEyk0rffBpA/86wqEiDiybCoyGJ67tcdD9
KsDH7THWUX9iH2IO9hxsmoqnKV4xLuMR6uC7PfkDrrDdCb2opOwpgnkFfXpLyett
yDETObIMHMhdUnXxPbkWSa95DgejLi9Dguu/qHESKmUxEDrJmkQaquOwTP2FaU3t
T8EKaT15nNgXLCG6EG9LijU9cSW/TWG8KlI2EGsIynP4UcV2vh83NEEOLFZ703kk
Vs7ylyvF//rS5WnlEprO53esECWOZhF+4yS3cCjlQPEqx1vhgzFW51LgsI/L4d89
fTBWJ4lWvWBkvjx21+CFhYQa0ImcCKyz50auHQFNZ5he5rAhScang8dbyhWOVDeJ
ISe4/kw/MrUHed1GexjM2xxfMr+9cfgUQI6+U64C5VFxRqgPQxuIGoT6scEC/fLZ
rcMywbJVWQlPI5hiKmUJc0/6idMwU6GLiyeW/5bU8pJKBrgbv2rw0kMLFMTFx/JZ
gCX/E5OXiPv3kkX6BmsY7CPPn4s0B9dFNjMHZwx3ndb52vjOKkouzLesJs3kCmiF
9aT4ZT/L2GF8uNLhzJ4Odxl0MIq6tlm5Zx1OVSSglOVbpRIAdaRkPPSTx3bpQDE2
7SHgepOqzm0QdqyLRqXfkJwMGwUi2s8fwAoichXNxLcqcNsqkhvWaOoK5talOF5l
XQafWxKmBORoNs8AFCS9ymBW0Mt5Y11pcht6oxHIoQ1t5NGi4uj7e7YVRRqS+MlI
IWIaDSpCtrd64LboDf4YYYbj/sK3phtX9+dqLEQvW9Voh3ZopHPVQlGiIiYMcshx
vc/w8fGp2A5Ilb8poAC/wr9Xb4H/hbnDZcOYon02Hk29KEV4rjI7gYnNKVwW4Dyc
kjGdIqAg2chOY1kCADgl6qbqm7KFjyjBGGEh9UuXLmxNBmyTbmXVse4b1413XuQ1
QFqgBMPVVRMr6jk6Et65lGQYsSqnzroW/itqvVqWknjG8GkB3MiCwkhVLvVK2UoG
xCCkR+ffzRMBqwswekIy6QpSa+qLEC9Wk6L4ipfcFBRsQuOvfl+aaRBLd+zMD09I
fyeSiWnIUZb0NVmux3eUK5oeTQHLGJoCwAa03S+4X2pnXIDznrSTtE9egnz4sbmp
OXGjaHW4VSql/o2oxTjVqLb2rwSVwq39CvbnVrp8lBGApRmtuCqGp6/dT0l1Mfl9
06CsPMASZmjeiHBTiPNXlCFd9fARc1BksCqBEt4VGsjnzmvY+p01rXShl+kOiHUj
8Vgx8Mwm4mPAk2RpHFroLOSOegL98kaQ+4x/Nh9nxxN+XeValqgDajPDWHVWPQBD
NG01Et4Fy490ECcwr+C41Pkp40xdwwqgY12YwCq02WkZA8t4R07WJ4cCwL5Gs4Td
lTcYLkJgAYJNhP+dlznzAH9UQLZtLSp33K4GPCLm9EA3VM9U5nN+I/tQx+rhb2TS
dbdPgsIm1GbWhk4nj8pe74LRokob0cKdnel68PkEigQmLrnw1J0GDHs9huBLlA+/
mxdprHDIzl4EA29rlMK2GhQI870ql+RjvmJolmPBqmSr3fQznIVgf7zdFmarTJrd
9jlgY/UaCk0vGXUWbIflhjtKY7y9wqRHzB7tVEQaJrdEHKkTBGK0Qqc+4EG2FH/u
XnMrSNR5NRkD93xqgH3o8MU5EisrBBRTdRx6jGaQhTRs7G4gXaMgQ0/5QPPJ+05A
cbLO7BR/ZmXM3DzGF5yV4xR/BUOHxs9yqwF1TDyqMNk9wpouQ+4wDESlhSNICTbD
YN6j9adBByVWlfzpBU9L/4pGHVRHX0Mj1bzCzQRF/qNOjVIV4LUJwxcufRUcGDQ/
GqKSIqmr1J/lG/AyFpaJwDW1EXn3aPwQrsf3y8eSRYvuANWmFYG3PTQaAc+wbec2
mmpmCJwNjKii6NAxcseEuTWxgYEzqQb528yik3zF4/RBN62YCe8i8yDFwINa9vaQ
A0XufXzXzg7JFNvNAZJqhVh5xHAWDIsGZgzpwLZ/gEXEd3+beOoGKafB/Zv3LNOi
wV3Sci3ZH4tByzHkn/Ey4CEjJDX1AlGW+l14N33meEeKi/UuFtWk8DrIs9tCSBu3
/lDHXgglg2KGsTCBJYE0I6d8Io6FaXTTERcLWLFfYPsY0NpoBdCFhZGL5zH+Q2er
xe5fzuWY+0hcbdsEKeKdLMMkcRJEkSnEAumhuIWhl8DoT6RYS2TnWIhlM+KRJSKL
ALU3MBZXho/sk/vJjD7lP2Pa70OXOGvHwkg0e0+HG9fcecOZBy0hgwOl67Im96xc
J6X4soCbuYzXTuOc2+GG+7h0ZL5Mqk/7henJTUTmZzY533PyqIoYWhqAC067DvEC
fj8oe8KrifBzqqfPSlc98nmPXxuEJ9iAtfH7agyTVDRYaSRVNkaYmqHeHpOH5W+O
FMNp3UOEf1d/fSwCMas66iWb3VYZ9BXsZoi21xjY+/e7WrKVP15EswhZgk2rqZsz
2yH/9Uk4p+5ihV4zT19mBcb31c1g8aADVAlf3L+A9L6jNdVWQm+zZPi83jCX0VzE
yzlumGzQb2PzJIxCq+CMpe1hEo6u9Pgra6X1tA81B0vfUaPHej2SKjeb1JShWOjz
opSp8lQZFOUvR1UKqC2gFYFaiovkX1i8S3jn6nIu4jdXzlwxVvFGbrNg/x/vXkce
UghY9aMZru4xNAlMqiSpY1fXVsxTuJ/sge9QZTyxOoVtGEwh98Qlh/Klw07dDC4h
GOxubbYREu7iI5yyC74aNKwDMCPeCd2qZDi4XsseGhv2Bcri4qczKHCgtfDdy/LW
+vIALh07C+jwqEkYJ4aTocSRwhWr43l4ILmwl0mmxDfrAkR4Dq1NNWF2JikL5BtD
UEuq8XTtws0h+DPjKh3CpLStApu+kUdQjkvDdfslhleELbZmXVxyAF/7QJ3a2Avi
IuNPrTrdr1ErSNrUQba1G+R3HZ8KPOE71q4OaQgkPRmuPpLuIQogSk69P/HgTx6D
3vFY8l0+GvstNQWL4ZDumJnyVx24aozARk7SrbwkPcbqbM7ogyVBet42oSuspelG
wZSNmdn/pHh8f8gT6tD+2nmQBtxICXQxTQXdxZidX5uv/Sr5DDTJXAs4uVp1GcBO
SPENTgUIbhANAlhUtSaV1B20p8G1Zq+pmM8zGl4cpg2JnoUM1qUu8iAA531BK6Sm
YOo8VL0TWYTsPcpdQ6FNKhnIrdhXq8BDjiFrKPHokR0tlf/td2Xj/FdT9epKD7Qf
aFlbfBxqSy5WbRA/us9snPexuH72TTUky1rFUYbGSGj/nnyXNC/AELSuxGC1KVRT
FUOg+bAaN57CbojFcfD3mzXQ37hTKtJ3GDUYl2izlBZ5L23RnciBV1W88gyzfopi
rJapoUTj6bcQ3G2VZ1f+IbPo4CJL9ump+odNmwCUxbqkbtQowwigjVtMAKN5zvdG
PnH9Urbr9/RRQJHQAc07/70ymnsQ0JuaJUK+/xCFPOijVVascocgAVfBUlTjzi99
7nagvga/ZiLfT9KUlOdH2wCqxFhptI4HPTrqocFXGvrApD2vPaJRlydH1T40X1mb
gkRSr7lZV8ulCDNpnEOwfQT4Kfu0R6vZU1c+DZZVeZnU6ys2RIB7GElS1rOZHnXB
HTNIU6gywz03ZZK/FY8k4EsxszSUHC4iqqN9gKur7iPGdAoQ0fMtUG59Nn5YbA5f
PgiWGHU1Ylfd8X6JidZYhP/c9+sH/7VoQAnn7hL2mYIldKHrkgWxlyZQ1JGYJkNh
KckXIwHQ4U4jsbiN6CUvcPSQAEdBzeEJetdTwXzvB3mH79C1/zxGEUvxEp1E8RtC
dmXURcoqhE8ii5oilR7tcKvc2arl09BTKt16PtkUncPwfMpvsGEBZKPBn4FlYLxw
pnyZL7ag/WXs5B1BQMFwMeFtsg7nxPCE6EdZWfdHBCnGGIGjTijCNY8G80sELH2e
5n1xevyUOLbDnYLXvPQeDlIUgIQZ8I0w8JENzYLQELCxKW3U60TAAMopgm6HXhfo
Bq3qJjbkkKFGG6GZ3vFiA25emsialuubSy7hLcV896MgIXfWTbRelBf1s+UfBT98
Y8Rbmr8gCLwJWqaOy8c/Lqw6qYC1hlgVleSCVoCGtI2KCfk8RYUExBEJigkS9+VY
FVlnSGdraD1RcbrSZvzgVH6WQhvDKh3A2xxqXgqFafh3j0FAS5PL3xiOQHh5hCP3
zBZ1kFaUVM9S2ArIOiLqrpaQBAdmHoYgYCgFTDy9ONgC2j526jB/u8PZsRQ6kmQP
IBfQCu1zim2fc4U3572/FKWtJMIqvz8SiJ7QnBOFdg2sPLOidW2yOD46YtQ1ERPk
y7rx3t2dFYTdA18kBcqAVdvUyjFQJlg7KeEEeKjsC7tRNvwezKN8jsI+mIcuXRWX
IgU6xVZe+eEZKrQRayIg4d45FhUnMptCTihr8JRI/kih4lnASHWnT4kjnWO+l0qt
YVqMCaijLM3CQZ/CDjdElNcaqGJjFB3oAjbE7zW6R13tRrN4Bg+WuP2ENZT5+XrE
vMKI352sKI6iN4heYV0W97hXWFTc799wZALc5mw9dJYWuRoPIqPWqbNgpEChUWpJ
C28YH8ksRucRTrCwbAEu5B5Jw6bUp7JPs008o6P6ZvIkYN9viXJ09tQ/n+Jqsl22
vVtbzdchtx8dBQgSxxYN3arHFjUClTU5Wl77N2bGV8wJP/Zvlh4Lqu8hG3HJ1pHJ
n6nJaqv3PCqQyXbxMgrdMsW3/8dSQq9ni+xuEM1OrFCGqaCkXgXbqHVPruN40HPk
nut6te2YijT4ImuO6SNL9I9F4z3czZmv2SQqoMD4+NlSCZ3GAXo8fHUWvQ4r784z
iBHmbjeG7q5KmEj+pKxsTR0B4D6qymKU9d6ZpfWqD0I8DVnfh91mmPr/lsSICgPE
p6JUMy9Ol7mMLGCXsSmELhS54sVBuuGfg7wtWTfUUXSOW8rnutXKQYt36DulkpO3
NqxdaIOK81P17sKQaSVn2+PYIQIdGfndx5NClu/6aStoT+WWjkBRZ6b6fWOCyXtk
bTlhNAIZc3D8vj7VQn2idAu+rqkl9L6VdWVD08c1W/EEbwkjFC4EyK1qG/94bWHt
5AU3ykwdioFhcmYOMxrghcrg58xINa6s430zNcIjt4vFlu3mWDzrWUspGTL/67Cu
5935OMcqYDhnUXZ5dE+Kapcdh0Nkl57jv/dw0imXTN1j8r1Mi0FCTa2YoYIC65FR
lAR1jDixzKDYJ2c4vqztPgKIsS5PofHoyoQ4ssIO4bdTBlczLa977U3ilnJSPQnb
vU/+DVL/dctBRlnK4vLTYtFYZ6NjEEmRymUydaCS7CIW1e8DK5Q/0HrfQtYFIrXx
Evjl4mI4RAhqBuwWYYqnpLIzaf0QtJ9LMQm/DJWnoYDVLPodwa/K0mhP7IE2wTU/
SuMSMjQvn8pLsq5V0JSaVQts6VdUI+kccV21tvhRlfl/tzBIip9zRa0vTR5HPtsz
e7zZRUHDMLCa+ZNw8bxxxQ0XcDjuZmoVD8BAacdGyjnKLCqoMm605buTphEivnJ7
t0VsH4noHWFWlZm53JkyVvHgUjzip2dx92WLicc0YRFOFc/sj7DiGxQdrZTq0Y8Y
nHbdiqfxH/qApsm08k04GPoU7k3mjfih1Zd0NR27Pt2yl3sJT9qaCHN8+0AwvhyJ
VTdpHi6EgUej0rQNvbKbzs0iHUKwOgKFtHPfEodq+vGmM+Y0tPLDULkK36ognhGB
OJvTn+dcpsVEKNpLX+GQj5JvfU6NbRNXqhBiZbRx+w1CXxXdqORxtmdwggK828rP
vBOa8ScXLF7X43pHvpNryzlu6vAsRvieVjhURGGJVEEQhiNrdBMIAD0PiGCkW74s
5Nblf1GJb8jfzW4hnAht7tFrWbAQ8MOfBWN4Hq5SIFMMfN89i5YQ08o67v3tN/4N
E6dmDJdw+f9JVclCxmxJUhuOZRtJJmt/bkKp0gdj/SOmUEooJK9+5rXT7FRpc5YJ
dTX2mHzYbLSCDc96+PZ4ETFqapzRuw1ijTgv8HtqgjHbt3ypaavF5dnEO0OkCM4F
QMfIPBhe5sakZqjSRr5PjeWHEPacbVMGLc22y18a1wrqrLmQ2aDMXrhO8xt33LXk
lemxJC2e/j7YRuY8yMC48O+UVT+i/DSSTkDMz/zKOaG99Fw+aG7F9QTEre1UrLSZ
mh+oiZJO/tkLT+4tl3uRQ2uoy2/aO91b2Vw0RfPfAVsjOZ2fQfhhYh+kAxeq5LqP
w7hPWZDXGCrq5pa9T8AQrstGwLllJjCFfuJYHR92WYkvmdvLcGiy6uRbYz3+JQPN
0mTu6+Q02U2HnsDTXauapIjjnCGVQLaBUatjUAIQ+O6qg/qq3XG/ru7A/8e3CUXf
rUu5UqChpxTwimQTc12eKA5ZJv4nmlfddYXmJe4ZTHBkhKFZuetDlibSSRixcaDd
0gzlKVU+tM/Z4ozbgMVmJEpPwzUueDHOoA6pDnbT7yysCjxNTw/OHNjsm14HxC70
bbebc90FZ2cZXs6p5ems+c7MhTpz3Llm7HeXMfbdcVdPkwZXE6fYYnUpTTCWqJyb
SVB2rxzHuigOUIEsrSrfPDUeXe4TU42UqCLSiRV4A8T5qKRpmrX1rEPxsdLsGQCJ
u9TZO7nO5u0WFXOXW+zPHNDmqs8dy7OUboSMB/i8SVN1Mzy6xiei5SuZU6WHxvn9
XgL2z+kQMaX0Y2ykj2dwqSPYlB6W8PdfxOFsGHIaTtGhljH80dgyY8YylqKhwfvR
snp+LvagT78gVFuG7T7iJbZhVitu/FMGf1n9bda7QRRQvH5FDR+tfDnwdjwDvDeM
3v8PsZeSugahtFd5LV7ln9QY63HQKa31lz1UVYMEfDeJ+16ZIRGe/S64yUunruZC
zR9ICzUopOEwbIBFWP4IkPxDfdD/zzkNaA7IfHapwBeeSzqp08U8CbXgJqWGhRx1
ZQ2dfR/tZLOGxI46HR2H2cqT7PZ3oeUIhzspia+/gWC7TZtopVjny9xMWehrcZVJ
gbFfzLs+UZ1L/5cKojz4YVezObTwYu+qbFw4fgYAtcCHiooc8ywHQ911Z/3wPmFj
E1ZqmGWgrxzdy5TM7i38Y0jWmR0ClQMg4pEgi/z7ZuUrxEK2fHn5ufw6MHw6wpVb
aRqIlg7qU2I1X56Gus8CAIApqdJy106D4ZDQ3lBMfF9TB+6PJV69Dnc8q7CrON1u
MBOyRUxk5SJrPR5QevtNq9CrRV0sjaA/ylVbcHMXtabFK6fhKIa+7e/xGt2t437o
35kCrSe8XtCSb9SsUnXe89obNVQG96kyP0Gas5FaY5c2JS7fpHZ7bFy14FBgHgTS
a8sQLbT3791iFCMV9/8h57jJ7SfnWdnsy36G6YvFSzc26S32lrVJhBcxjc0OgLAK
BW0wLv757xNvOGp6svvd2sJecaNrDeIUvppNwfKi6bKVhr9QymbGIwf3zz5bbnqt
K6Xs1v38LffxN2bqVmOhe72+gAJaQtW5+b/rGzdbIwT7y6xOzTvR/Mrxv9M+WYzV
2ThVzgJuG5B0uaQtxB8LLz0gkTPG5M0yCaQ8vBwsas0QgywQHmwF8k2n0Gi8TwZ4
+UCASBesq4jL7nHEQnZ5RkkC9GGsO892wMVO7r86aa2kIvoYkNcZgXQiGmSpgkbz
WKf7lppzZcROdIKHuSgxa/Z6eNExmWW5jq12bzdH6eW3Kbz37/aHvkId/T/JV7G7
c2edHzF8u0QRPF2vrl/XOtQuOAgrFGoXA4oC/5WZLxv3RjMS3sDbChj9brItEn8P
3frnFqkLvzvu6z8OxjMPc0ZR/IzB4iwqyQ0glx8HurPMswjzV0w4fHzeI9a5WDml
6pqi6LGnlG8B3wsTv+Y2BG0FUPS0pq2YvkHOT/W3CZeqmtcv69GO/W1EL7rsYVgV
iXhhrkidHwGGNap2Mw1QKF3cKHknO2K95PqJraou00imDZpxYOhlAAsQzMe5TqS3
GuZBu/c9nXnxlEX2SouXLFe8bbsD/fNTelcdT5DIladG0mIBTrlUxafiWYTWaVuk
EKGT7Xm05kximSQvl5liVRcmbVHqvnini9NlvaBiZvcnLmI2OIxCYzD3C1V8jAHG
iR+3YMTJzDfbvAA0fruzvrAYHdIJo32UWIhsK9l1wQaAxTSM73B7FQ4I16O1JMte
R7EWoOBJvwKVHuI+R6ZOEutwu7Z/kmKClp86c2lX//2tfgyj30SbvgTfmDukHb10
58IvytQyw/sbhbcJD4yx0KtJ2Vojt4SXxTv96SP1FGOy4EOlAQPNeSDJm1XlDQOH
EJ/GeP1vWrurvBL1cHWQP/O3hOQVxUMkdLr/xfbZDTOt7EhRCXAtISCoCrrfI9AZ
/rG1Qf7HS61gdHEKnIzuwNgySgk2kncMo1A7JgVn2hc9CWmHFchikqmpGcKU7cxv
rB8LmqF2jiPQpNj7RXx8KDgb7UAON2mAMZnYotsl7Wkq1bA1B+RNEzWxcUfhjkRO
AX7uXTJFj1/pzQRwSTCizGoiO+UW46eGUXPBJXQez8VvrvuTu46FD5T9fmS1mLqG
lz2YkiTzaLCoM9YeOJ6wZNS41o1LNLzZJzdeBW0mX4ef/wx1dfRQmXhpWfvA4vTb
3054sw38pvvhnzDF8R8yw3WlAoJ15kRaZGbXazuW7uRzu5EYD38AB+mkIHdjYvMG
UXFH1JuYXCKVgsn7KGlKErxTOFFRc/a/wqO6ptTsmM60GlX95921CToyVG8pOhYA
u9zoeER/Z+VOhfoeaN3nmpZ5dO+dgPiSCJNu0wmrm0XlqZ3W36ewfkSwd36wR38J
A8apYVCPxnRKVsRxIAIWQLSnq1wH4uE6JK07dPsQU8BVquJj/coVbxLj3EVl++8H
Rv6aCeDYDW2rGQRC1wPxyoOl08WSUr8U6nRPlnAwR/H5kfXzAes0U+u9GMcGo5ko
gw3hm9eXN1JKfqsRe2Jz9Hxqp+q4kfgGCTw5ZW866bFg7pIat8Y0OIcGInsmSiU3
fl1DdiUZiYxR57DKnHS38FM+qSDsAfynvlwqnUv5x3C/qywZIyYouWO7pfcXKYV+
e8GbiuPmxuQRlzff9BJVHBm6RttTFQWkSjY7e7colnkg9j4E55+RA8BmtJ7g6P5R
/0qQ+RNZjSEEudQo0AS1tmk4pKK4A3KqtUECBALMqXQJtHnUVxp55kUCJnj8bQiA
Hxsyag51pvup7NrZ1mKCbHhrEe+gEeKT6gbVtomD2EP1viowwAigupO+PVHHAYta
TVabCjnOQu/QmbSnACnOojJKYNam+UtBG5RXqVZDUvBUQRo81RVc+0DjRPtuaoXB
gtBMKh2YUXUnCZJ21PxpiIUyD9IPpJF7Xc/tyPvcTgorDcd8d1wwFDfqEsTv8Rkc
/NIlwA2kmmwlAAvHgtMJFCRW//d4u8bK+BK5SIu1Ck2deJc35BSGZxx+8FShrbHM
/c35PXBw9FVWDdqfOH2gyMMYs6T9r6nOAr7PYJB6N5HwfE37wV40WgX5L9pISUYn
w1+BhCEENK58Uj+EuGfnl8J430FTR5xx/Op/jvql7PxOQFPWYSqScuL8jsTNnX8c
lABpaM0d7tYH4UYJMv/VjiV+H8OEV+bB0iQYiGHOLzzeaEZdNEi6tbPtKEGQCHVg
csLkcoAyyMCo6cDCx7YxWB8c1NnMj+OR4LEnYLcoc1UJGi37oyCnaQxM+S40fn4D
pAyksnpFH6fYnP7nXqJKhlSXZJUo2Z88C8l/taTKusu57pa8CRHN924TxMWXImuU
vGqM0XRJq2Zf+7bRFyrPCWvLGMrCuTL3+CeB4kcuaQJuyiFK2lK/e2/A9bNwIrKP
QwlpCKv7BrydYF//qfdfT/ZmIX1vsCY+fqK+nTld83ziKHLgVvQ/RjKAIhQjbUXx
gmolIceNRC4UFn4DyJ97I5zaiyWUAIFDPdh5PcKKINTlsR8fowJFur//si/aBwth
eUvLhqc9L+p7QzYG3vqSl3DRbCQW02xvTpP75C59sd6r5efi9zK4QYgQVzBvSRyE
ozb8RzqCXkcYjTA6VzTFSOjB8xcVQKp0kWdIyherehz/L2fHQQSJSxwwVRqabwck
Ra1ejlRh1DQlcACF4hv/JU3v1qg7PNP9qfda+xHwcuJqxZlhaxNeqIGZv3bO+vAv
81PZ5eOp43fsBtLevU0AW9zpmoj88B9cs/OjUsNu9/x2jc+lsySpQ9K1j1B1Y/28
TspO0EyJ6r2X/9STnB9iEBFu9QAJUWEsJ7KftVAQxuRNxlFcvN4DG7N4L/o4Bkao
t5/Yqq3V2QWFRMGWgl6FVPuqbP6mTtCvx10bQxAD4Ox+S7QRrn/e7DKjCPzziZah
vAWhFvMSJsl+KYndIm0ErCbZKTzY+9+eBrhExiXWY0simwqUbHQQNO502dOdKXK7
Ths0bmYUpbdjKy0BxgJ6VdczwUh+lVozabSMSeHfuRkblb2Rxy3zvS+EtF9gfl3M
RYMaFE5qbB2ZKcVkJVQMFQAGViImlPD6kjHYJ8+EYnwKVPk87nOdxPPuGvcyH4Ik
mnJtCid7RLzTZyvXLCJb6EcAxYOVgUgX1KclktzkEghwkU0xYqtDRw7Pje/1Tnid
RqGrFgxlog2uEg4xADPetz4p300WJlvzyd11Nc43do2DpfNZ3bzQLArmltk6++zw
OJUcGGyWmUqbrf0WIGEGNqQIQMo5G7Ys1d+iIUHobBnG+Czblo7vgeyPJVA3qULf
6+dMjq+g98GbN9D4An4HAac9R1JTRJtu44KFp5pkN3ngYNo4/W6xUm7DboLAhhhb
1VqkcOoNdYNhHGgxD//bH7oq53ziNMfvDeiAiSxaVGTrUSRSVdcowEkfkQcPANij
remJnXdw0uBUJhzhOkQcFwwxhv8XIyFrvyrnJ6Evpzcwm5c20xqpDp2kUj0WwS5D
C+abxlSDGc7MdVsQzGM+FTVwn9L6asWuFBz5pXm95yZjH083Uz+eoiRFClG/BdQm
gn1WE5ZMlcJ47z8E0UsDfsotIB5uv0c2CQRT6DHEO3SgQW6RdJlYZUn7gp0WxTHW
ZqnMfFnV9s/tEwfqXN9CykwNWpVqnWU2xkuqA8Z270lyKYzJ6x3W4GefuVjG9Ea+
rwHQqUru9BOZWoZxbMOuf4QP7xSflRY63g9DzuqMr1k1FsKrYnieJEoEhsj1J5An
qRoBkrPbT3gJLjEPlya0tUwmiEYv4Djo7C9orGn7N1imW7O/PtTBx0wpIF1EEZd6
bDPDuWQE2SGftSBa2uZgpGTaOK7ZSOKLWoowvumrmQYSja1+tc/JfailnWf4urpR
4kO1NV10hOaW+b4q33onTK0vKVn7/8uZP+yx/95pfUfCJtjE/bJJxhaK+Za4UCTW
xSNgtGrlVBWtLMJ9rJ23hTCOAq/GX+cZ2mGfY5ZdUrpQ/ZaWcYtM9tSx3dX8qtw6
h332Teox+L4HOGy0t27RJbb73oVKRxIADsteaMsVGjf+WbO9l6j8nfKrJjC3110A
3znNFlBWll+2fZ1ifJ5a7WgqoPMEKU+lmLS6U+FBttgAAo1l0hqKlh3rhTcq3oPs
jyYv7K7HXmjN1XXO2cNoAj8bG1kJHHIsh8bRWV9c4HlqO2+y3qPlGTU4VkG8doI4
rBHWM1WwBjsMK6cbdrf3EnT1qqFJRUZgmXkioN0zJvdmP35ti3bmh/Fg0/byMoUD
u4zox+zf8/ubi2h4GvAjH+6ygh43V2MBjZ8JFrqMjvc7bqoebeTP1SvdVQOYtLD0
fFK6kexekPXa2+VwVamViRwyuSGBG7Qj76IeaB2a5DV2o8IC2bqj3mg6HD1S1ALp
7d0ANZFlnVYVpyD35UyIhPPIJsyUrUAhW/zPcsuxnQ+W6wOEcLErzSdDSz6j4DtP
dDR3cgOaLClF2qaG3zWeCNDfOCoX55v701LRQOii9nUf6tPqO3qB3iHuji/rQJqz
ffGbGAHssSuXceQQdqO/CENVHIK6AzT6uiteNcR6A84ds2qJDcBQ9Jez13EFiiGp
fgn1j62adM8lxauEbbNvlVuOy+UKlAjRGkuCJxOUP20QvEXgVLPRFCYcWAA37Dmh
KgslVMtVcKY/wtYC9qPb+TBBXH5DYeRo/1ZGalJ5VogaTqdIW2loovfFaCuXPWwY
PaYDI5cMQk6XGp4y4ZfUMIDziUF2zIFQ1PMc4voY182hklPOTWslQb91dJQYGKeb
UQyOf3/0aNLgGhgim2+tcaNbFx7LlItllX8gbmaNkd2Mv10ekRxo/t7rjsixWZpf
kthj3xsiYz3ppmzQMjjoV/pC7HpHp3ZLvV58ZbLbHJ2pyAtZ8HVjg7Ao2FkCCn4v
H1SDRFOwaQWnaCJrYklaISCUmGmfscjfYXtXrld7yKoQXBh0zxYsH3K2oSdSItze
y/zJ+jE4KacF3bi/DhprBAkD8bfE6o7/0TNMOPF+nbtZYcjvxpX6cf3pVsgJI8bJ
WYCTUeUemQRJ/dOlZu0YNZPv5iX5IFGrFIjxqjMPpWlPmEDYfkbbk+AEm8dB4ka9
6vE5gJ5zi1l2l5rkFaNzAkmsj47ushEr+qSSePp+xiZIeBrkHR0qoI8enzufw6au
vTSH9CIKMs2s/fe0TBxWGyjSnw6NxM6qwEAk07FNlDogKLMPRTKpe8lVQxJoU+wQ
Pr8s/HqdygoVkgtF/RO8yQRho9klCTeUI9NObqAISDMN611ASi60LRdC8VCZqNvr
EVHX3xPIJafxDytuCWsJOHLPVawJgTL/lMk++D3fr4JsoF6HDMYpQnB6rWm4WRRA
9F98HzhqwMHj3IdWMqTMX5byyBuFvhU/+y0Lz9L89TGg/xsDlZxkxRCeikSQhKoJ
JPjDnidVfEkILIlOvqu1Al0R+P1gYM+nBlcwFub8AlXl5WAWyq8dDNJA9cW+HklD
1ulxuOISzjI19aJ/d0AQpl7PZIVGTVX9SNysZGft85bTVP5GvF+B4xdkBj0cpFGs
7V1MFXurC1ywpPWyEkP+SjKk1/RvV5bppqzEj0eCFqJ776uxw0/O+FgkyWc110/3
baOS5EtviI2CmVLlTFoPP8qbqckfRRbNZAQ+E64Kf0HuTAMgKy5qRw6IHI3mz6hB
S7vLuFdYsW/7EtBjHgU+Eg0alHK72BiUkTludGZdvMoXZrh+bp5/E8LTqBLL+YjF
OKqZzsxa0A4Dk4PGLK2McOkV09/4fi12cxN8aLlRi/ov4Z8xxOIfcTUvyIt7816Y
XpMplyGY9EHmSZ+f+77ipTUDsozYrfVmnKIR5vo0+DA1LkmrurYBRfzFHeI2C2wM
rJG28nTM/KJrllZNrNfXi/IpN3aVpb1O/XHxUry6BL9eb6MIcCR5jyPJJgZ5BnZg
CqQ/3i+anUCI11lb4Ma+K9+VV6qgx5ElZdL6IaEV1K2SfPcX7fnI29t+X8gVWe6v
Bx+8HXJ4KJvqfb09OJgbbi1f3Icx5hnv1kRVV0F0gam3bYhrLPhbhHNChL68BKfC
93FSUpp0/oOJrKUcIH9TXSKYqYIyun5ZeYkfe89SVi0liGm8EDY7ipyjwRSRlCeR
Vl6c+Y/Mk3Pyrb/zLuKQTtYZ323R3lfR1/EGRnfnGCgwZnfJLgoNbwdg3Kf7jP9x
NiElw1MIVGoo7oBGN2JlHtMo9qXHfiG9czqGjuGwtpLJBkY8mNV8zxRIA06Pe5im
lArg6S1c6bURiQlv6Rw2nL4o0hY+WY+noaZdY+KDA63quPvC5pItIbd2xic5zEel
s2/EFQoAcNYynfhetDJ5Ol6IghGgMwccT4Kk5zI85SgYpzciueR1WpRa6o4m6Sjz
RC0juuAvHsKr4jwioYCd8jg/rgrbOdcufL6bHtVOf11crA11mTdfo8OBJUgdxpEi
QaAnkyBsxP3QxzVQZMkCHxlDyHOQh4eYll44sPeb18Opr6v5z/N3PpEVBuiOylUu
pKFKHCxQgs0ALr5XHEYFYr9y2jUzC1gfdSQL4q7duUKltBxaExVrDF/Ft1NThTXt
jPObGjGoGOyY9ojl3fS52tSN8ldirUt5P85DyYIrtnoY3nTglER7AZPKErDvOVKt
q+NeQtCBYqujbwFEo02KlgGEycKNwwcHaKnw6JgcnUtJIsmeINNpbBvUr6FJQHi1
PSQeLR9d60s6/YYLyyjJaEbmuy5e77RqTVgvKZzeBxLFyKmseLq1hG8mNq5r1pul
Yzn1+6WeuJyG2txoZUJV+s/t81k95vDTGJaJYwjD8WUItSU24CTm1HTSssc31cj5
aWIhdqI6dwRuN37W4m61sct3C1UlYEnY9j5aSi4bnnw7vtj+xroclfmfLdnwPD9q
8KaU2V1fLXXfpIxCVktQV21uEuGoNmriWBubEh74iF8JQ2YJGDdtBWXhkPsbrrW+
uv6Au3mJ8VKuM9ayzlcEDZVkD5EjbBYeVPl4tCsdeqrWkhHSTS1T3xY7zo4EHLWy
arA73UsbiH46F0s5Oc36qECwL8v/D57vumDzuBWO64PHn/bvLPGhNmOagClErk3R
oA79SdOd6BGuoqnSxQ4eaOz/GSnKwtAc4KwcubppwaaosLWjZOUUtQ9jxaCEN0JM
j5ViLQTt9gIkEzpSn9yD7tQTklkeXe6qdJlkTXAvv+tvHqp9nsDYZNSG5ambA3ZP
HcTSXLqJPOvrYZI0J9XpiCpM5i4GAm28v+H3cuP6lnBVJuQR4r0En2Q4t4AEWRfA
SQUcPtp1Gu/hKZmJVIoFts6bzPc9/HhzNIOTapn2AcirSbelE5B/qiN/I69BJQ8p
7bgZD1IQ59mymboIO+JYEtb6pWgfEYX2AEjxFEYuk20/nIDaXpjPCegJoUGs80ww
UoS78OCtTj1Swb+Ml5EHUr12RljKhFf/rkINh4bbAopSkc3rde+uJGdkppyq7ZVC
JTMjfWYLqcg3pNGVT1/S0q4dwtIchB89msdbNi4IvaNvGkL6ePOQS91wksFwvq86
3BnMFpYBALniFadWF4ekmRbCgHqBD/gIngc6udIMbd25XhetRut6CTpO6s6r7L/G
XM+xpYnKYBh1GQLxK3rK3R6mb4o4OGqujWYTrExn0+zgvwucpfpcTNIse8Q3QEBB
RR+dYz380vkBVSi0H14rL5D/qC+qpC5uiYIqMoUkl9C8tUbUjOvMWZwUeGxOKJWA
RYbI0k5wSJvqVUoDsGTNmfzhPGwu9b4ILdT6KQcGlmfls3WayuLPr9MdOfMkwslc
0R++OTwdxwWgG6VSJSLuYdm4fkEsSUNY8KfsJEo53Wzm3dnK1EizuRnwJiZMmjVH
+M5zkjgk0FFIewAILp96kOixtZUST1FHO9jAvrzwuAv8S16AEW3eTaluxK7ooM0M
FePTnp9w6lBRYHFPbUjEFQlQYe39iVcRmG/1bLA53gEdWjoVZhgD1HQquEoae/c0
n4DOvHF2UawinfMy8k0J0iePLWpkKoYUQHoSkyWHt54iYVOEFGM+e13PsBTI2g06
Arz6g7vNsXIc8wuqPzu2RgWEXb40qo02MsgvL7AoZD7uGQBcCv5fbX1P8waYx4uP
TMj3Yd6mJGvNt5vw/cjWvkUqfj0R1jX73/c/T3SCAEgEALWQOjmY0egdP9Q5dOQj
qybQyqMJbLvmVpwgPuGw3QBeLnXCVC4NtsQLWgBNeoM9GjGzU01XO0qUXI4yPfA9
vyb2pVsj4Z3+86Q5pZc9vikX7C24bqxnjNfmjz+/QqskLBwfsLJ0AQTZmkyUbyg/
0kReHLVXsCmFBzUM2kVLFfutHzKyMiget2nfxmMP2BRoxoYTIm0ay8YMb17TjrHt
X16E3rhoTc24ryoSWzncxT2NrVgQJEj8vlBJtPu8X8LzJzIVFxbyMT3aUSMxeaZ4
LSN8ae8yU25HVcjP5BsmZeTIajJIfv9HZPuP89NgIKQcykbFC0GdKyjjU0rMORU3
HUO+EPRqo2DWLZ+4jka34u2MxuVLmDCoApjkjTtYtupoA89qCB59DZQhMhLM3ZJU
na3sxFavWhtA+ixLYg9xN3sn3u+myXNukVFWfT6XdKWdas9bPwC+CFNJqqWqkP7Q
ROZoko+uEYl+QAt580rD+A+ssG3ZZ9w7jqGh6bCvBtjQZA8tQuKBUF4nHL3q4tI1
g/r45bVocxDn9rGCIu9CgOvNUKT4/cDae31kO6KtaczX0CMMUJOEKNUFIN/2i1W6
un2vdOBAb3i28bfkFRuN+TRFGm0/+U2m3yVlcEfkBeFsXPnPQN4QcRklodkFaucI
CMVmIip0jxOTNhzJAHV3WE1I47gdeORR9QWtUdS9WqctbPFMD4XCoVLKYrY1HjRx
8Ma+oB9599NzIoHBbVYW/DWE0FgS/X5cJifPTKYDfFkGb7M0PDVLcJU6DBgWT4NZ
a0grFdfkaT9ZcMXMhBBAQZF4naqjhPwQ8QhZxWp2WP30wpG7FHPUOglPQ6AtMJsQ
eMQNHSOGs+29Ho38J8jQ2TI+Zb+rSh62fFPCE4m4lA6zjlrZcDd1kr+G/JWRf3b7
UI0QfPxjMTGl6dsjatsO1wxpJ3BriHAA9lm1LSCrjQQ2Ns4s5bOyJrRnmhh6/k1O
rnrMTOYI1qDTWWnKdI86RXGh8Es9aqIfjzE4HK7coc5q90Y1DUTW9bDlnaN0cHOb
J1pBBwWWzG9fxHhvdaqX8uGldrVE5Xl+LJA0UIErf7jG+/HtQDqXGyWAAeyppdrN
hDqYkOkJsLgU5hkdqrQguqaf4eKyh6pPIj3kAWyvCNcmI+9nprTOPavrLQyGQ46m
vtDvc76MS8hQZK+AMcSmIiyThSsuQw2s6El0I++rm5kQOzLT7Zr/vrDmWec5DN3e
Uk6k03bZx1fAHD3ekiLRJ0qq4hISUihQ+VKNXG4/Yp0k3WB2lYy0/9snfkYgWxKn
cq1WjRvvltfkWd9RJs1xDHFGuTcDuQXgSsV4GvoF/JjrTNgYEKJo40GSdDO0xbqC
lHqmvzgtj2JELv/ZILurJO6mXpDQa3gUFubqByqxXD+rHmVSu1Vk7XyF9kEkbfXi
fyNy8iisZOXMZ3gkg2WPw/tKLPXlPDhIEnQBc/ehJkw+13z4pT0k+uVrSowBOTgK
LrlltkYWwiLSoC/VR/mX+8u/VNlsfu4YNb/IU3EEc7n/O0bZdzb7/4apBwMs4zaF
rLnKpS2GhrUIW0DZiR+WxEmsGoJg/l1WTes6SCqcOJb0/KYXSpfbZAsQubhl1aCC
z19dw+F5KH1rDAmJ9/2jLLjXBNLk3yBbRObshprSlG/fcRWig/45BrnBV97I/nO+
nKSu0OSZznMPvbelW08zIuKx2mCzCR+JAivLvwaFgA1Z9A4adxUNp1XbDD1yzi4p
v1rPM8IshnGKlBKGj6McZ0KjURU8vrqAleH5AmxFGHvy9brO3ubiN0IGjjaNwVPB
r2j+m6QKj09o+kUjITq4sPpL0pML/G/T/xlsSZJVSEIN5+xM31aWLgDPaTV9OQY5
wNkAKcv58lGkw2N/H43z0AuVfRPtjyMwZL/1eLQGaWu8VwXy4u8fNh6I09pcWRje
fh2J3VbzzvsnqSary6MmR2TWTskB/0qoPwGKddUwSRcdA02XPo9mRV8liGqNXVoP
yJgeIRCSneeuSLZWh4Jv3QQP9B8YTWHaX6qWIQK+3o+I5QbH6HT6wwzh1pwIZzP8
wWNVav03n+vV9P3iRvNFZYLJTH0LwPTKJXnm3ssGhSmyuj/u0nPnIHpi8gHlpO0O
uD0N6w4gzZCNKmO4d+KWJn9bUEACSs7IX3wez+PVPPXITaT2sjkSaoFCWnsmtUwD
x+OynuHVuz973vvZ9yClb9zHq+scuiB/cxPG4e67qcK6CanvC0KdGthT6LRDU6xG
EZsuhidRpHeLY+0cnoo2UNRTu3ctV5PyirSWPAX0iYDQ/+6PwbZ/AP7o/moiZk8m
smgBh5ejZTNBASLyneVC9rS52ZqpeZdBjI5GHRB9MI0pQz3YHT4gUOkSb3W1xgD3
vS3rY9S2TgClaI8sSvvN7b1AliyfZOH3sPazhEkDFt2oJGRnktit/diMbd3p39dO
rS8/be1oT8qAMBMuyx8cRtcrm+b65Cb73oLxUUpKIPjc5s3u/7onszvYusMHOMDA
mNk5RsuHIa2iEx8TKo+WuMNOZYTUs+vT4BWXEeRKF1/xyTB6P5IBnBvNijqBYIGY
L0bhMsmGBC9L7VVbrfM3aXtcJ5Kv23dhLrtSsM+b4rg7MGaODAyHQJydo9fyeznE
KCbR4J/tyA72heA0/nXM5il8JEsnXfUq3Q6BujgnP4obgxRPzzGcGtQhgBExd0a4
tMIqNvFSI1tG5UB8UNCuemFthCYAC7jbA7bcsFaMz5kisjuRBgCieKtSwuh7Ao/w
p8opmXXnwBA+2zbgJ3DYFXr/GVpbr3vbGY8EBZi0j5hL0AWYB8BE4lY+PUwiddhu
2WZzK6yxz1V/qGMTKbAKDIb/9QL8Ag3isSs6utIwrWRYAPr7nHljrXCU0R+YADVM
QoCzJdGFwyoXe2gMqXfGxkBziKTCvhieEpUdbn9VcF4L88J/rSE82zHNHCVBTwf5
4B9OKI3m7exErL+cvLzeOqaQ4TPaGfa0EpsLOkMT4ecGAKn9gd882oQ956y9aDYC
hn/puPqgMvv4G6BkT3wXz1k5t4MoMglZlMYRlVBeoI6kcm8gxAl42WOjUQrtvq/Y
5mRla99IZtM0wLvnOQpcNv9Qh3YrY40phi0lPKMA2vk5Lhvd0J6zxdX/eo13AqnE
ppM80ruhFQExE8PLErzXy9wiigwt3IxkPQkt+WUW2trRR/JJZNIk36zr6A84DjiO
5cVdS9288NY7MqXbfW6IJu5JLWg7dQW7TlBaPspIa3SdWTCFGixiiyoRhhTtX5QG
og1oWYCeorJj5ZfykQP0n61sRyFGn3s5xEFe8SxVcq7Un4A1AWN/hmx5tE4SC8Mc
vyVsLZmJV5sdNu8DI0R6lUZfITowIhvsasZd5r5k5L0UBwGEsKImo9+sAKa9CXwC
3Jb3raZ1rNPfvvpitAqdBaa8xP6RONtO7ghJzrhCGLSQ29daP6BKwRGW7MYzDDfR
GEt6u4KhDnBM1qZoO2ndj5pkkjDo/kthno9Om0Y6/t3gbE9yajJWDPnGWU5ftRpe
/gw6WGmkihuuMpT09RMNXEB73vSuUJcCl63FE6PpApJWrtrqgtew376+ZQTKQ92Q
EnAMulGRg8bhCuvOt7lyu42k1DFe8JPCcSRn8LauYEdvWO8WkNE66CqI89QdDTfF
WCQlQLwDbP//3huuo0NyGnwNDjVCp4P4RDPXBDnEv5kHCQ93DhQT6+jzzyKNYQO+
9xZTH/IJuZL3tcsTNtvNmJCZ7tOlOYr9Bxolg6pccv4rXZQaWynlNTkZRvadmxWA
RtX+xES206ZHMIbCkLzaTPHbbVHBSsSlgArIsz6acSL4IQhahxxzwNgohAYjFpQN
bGc/EOxH0Y8PLG3w92mBcAw+NwP4xpOcZeQ3FH1Tg1W5ThIvSJRqIZRRA8lKMFsX
yox4oe53JVZu/gCpf1MKcxhnGndm+9lWg9+YADR7/DC4eE2KPdlvurhla+ac7aAm
28m86tU4L3aG0jOeyIjpdmW0l6BggnHZ67+PsB8uAGJisxIbkhAk3JITSgnCUEDP
vQJSdRPSeNfdVY+Os/4S7e0FSHUAO6QaiHdt4JQk+PapG1xe1MfCozmQGdoiD+IT
x2L7d8EXRppr8YLY6cHLNHBORVvqrH44YhUdNGTw2Wuz3YFt15SJRXTQSqllKiRH
6Y+iM9tuwOuQ+rRRDbsy/MNU7L6IPcnrFavz28/YHE5OdIYhyvjkcmA/Mt+IP6ki
zCK2JvmSP40QZNUx244qbW3cB4o9UGaLwrYLNmMG+0e8t9ZfuKKa4AsQ/s6WKO8m
rplkG7uhgzeq5TjlVZyHxNw5N7cpDDpwHOWiXm30uwYE4W2QAcwy3US+8YebSUmL
v1Tzle0A1MabdjYpQnhJUf1b60mn3CWGtjSEvjkt7a1qaUuY5ljuhNRiN2Rrk8ES
D0ti95Ol29addswmPPSocw8ATYaFBKQ6EhpOu44/S3EzGPmmnIONTrQT7tS56Nar
8zdIYZMtkGYp3ni0RyBxVzwlFlIRWK98Ztw1abjKNY2CcwWpF5zRfA80hH7h6oz1
YEPHzps7NyPcShtVVCll2TvEnYU1vE/hm1rosW3a9Ht1Z9CWWUwyQddNI/EGE6fP
cBMD1eQ59VRL480Q0iCDjwtMTjrg4zaVzEKRGYymy11oCyh+tBJAiBNrIWsv+pMc
CGK/vNAAoNmjzDxJ98dXlyiFGXTCJjI2nYxNTRTqg1xjEJlXyn+STNENnwdZ3lhf
k7Xuc98D0dpMEPa0w8jObnaloFoRk8WtfauIz8MHzx+n461f53Po65/RX0HmiMld
0LVOW5q6hAmm9BGG3fSXyqdM/qL8eO/eYJ/d0zikj6agYBAcb7BMlJhaK/4trdic
kiLagyZ/xFSsH23f2X6mum5VCxIVlcTCcTXrZDY/cuOqmFwpfO5oVKfqfb6M6i4N
4Fyjd2sbDDlTBczs9BhHIwWrGfkOyHKNr2blymODC4z1hfKiIbjDvS+GRl+YnUkv
UcrKySPCnjPwT3koz2DunsMdCuSmO8dTDUwCaWt0UyPo6ApZLLOvxphc6mb+dsRQ
prjHdkib2Ny0abWJb31fgCbSHbueLT4RsxZ7dT1ukxUXM6yXyjbDJohY8hY/m9MI
FuF0crCZ/MxHrlOD4+Iw9j3JJyyX9CWnycsznowM/gLNeSqqom5RM7Fm39yLji9p
j4XS2dxiQyrzt6EiQKPnpcKYuqSHojxUHgRtHfng3kuXvobN1PUJ6SRKPrrxa3iG
4A95PwiId6MouQG5mabDjtxk6zFq90/TmhUJ+TgVH9QY48xzyruTXRueNihUSgDy
gzDp/sCWaUEZuFIYK9dp8ZUYKdLdPMQdBZ4QfLIg7YvXOZx4eHXSUJzw+0RLaJFa
ZqFGPgcjf0A2rJOQVa0iX8nEzdzqAoAnxkq419zh1HvQk3dVWUObydjvidEMMp21
a//KRFwuSJWLT2ulKJryBOB95xmT8gWA9ndTdR86t1UfNhPHZ9fZ/rPt6W+szTKt
Rf4PyFT/2gTwp/TGZvzh4MjyIetTsKm1PlP+dURJzO0Ulyctv/8WBiJ2ar7zf08h
4mtzyAUm/vYpwSdZZGKkh3OWO9qafVJoBYNhl/EFU7rL1xRe5FBmk4NqiOGftcsH
XNiLek6fUYful/g5lp4IvBbkRGaYLYQISMYHQzWIyq/wwI5cElWLYwDrPiWLy+Vm
HcxV10RrcG6ITLtLaf1IP69C1LBTFTkZeNpo9VpIZH5B/Gtw8hqptGdPTCACHmrb
EvX94BvapqyRr+ildWnpi3VKtsB41A6XO39w0ZlCFJaAN47e2u7tjgoEXu5e5Vib
hAHwdBluJJwKP4bBXUQTErTKu4hCdzcr1ogbP5G62OwV/Xv1NoQjSxLB7fkAnrJE
jF8KAUbojpn9vBuFcz5rRriyxUmZYSpysBe5hZvSNn6hK3oL2C9FvQ8yJbY8UlA2
nEs+uywOQdMiEVVdGKbUDBMJc2i0OPXotr8rIhn8VcbXS4q9XS7HYLo7irjLJ0UE
0Cbyebno7o17Fw9O6025ErEc2n3m9eL5T07C/Xoy2OW5JTL9fWaqymbdhCF/1JXe
gOwBNI38jvbj8xNOycdGQS3nksPg8uLuSwh1OPYuXBY2sjKiFfzg1QRZY3HsACmP
WUV+ej4hWkiDuButy/eTtbW7uAn152cOR7YquAi3m/SSEr11mmgGmRmx3U6fzgeY
ByW/C+Fktoac6pVs08zjctHip505piurEUYUBR1fM2ZdGvZAVvsEzyYPyP+EC/aG
Pl3Fp/ky33LzAJPzJZUddpp3hCrncRFUySsetPqxa6mUQZFWCjQeKKKns5e0yPBT
JahpSyo4DmRes5qLmHNJgk4GR35lDirn04Vo5sgkDCt+MZ0JyzykqEAicXhnIhuD
DVgjJH9N6hC7ogZ5VmMTKaszgy9xd1Qt9irlAf/njCDAMif62jfO+kik87KJmIex
Dj4/wlMUBhxy7Q3GSUaILhdqSFMZz6C5UmhWsq5B6D3Q7Vtfw/ORvzEJUUDAC4qX
1HJ8EDIEWWco4W7DXkrTp8b+YVC32af0of+Xe0AbsRWIzzsVmX3jXEjnqkvSa+Qu
cgwgDVhzKL/KHNHiF1Z9aZ8XyVXZMt6jt58VNMvd9PJnbuS6gU2qOdY4ob0PpwIb
BML004n6CkqCLeyuYY8z4rlFttjYPd0gF7xMnPP5Uin82utmzU8LyKSpKpoy8yAP
BmCby0V0bpFSpJ2/eukScrE0WYJJfRrVMuwVlWV8m86YeWOFYJPki5LsUXC+KERx
MfkdD37MjTCyYaZ+vvC4usL2uM8MzpDh2uVXl6rigSfwv8AJi8kqbD9uywunDGj6
QOQw51VDZyaZa5K95BKEwitn5fpEycGJ11npup9ROecTOri/UigyUBWDMWi3jaI8
X+pNT2V3oo29uQLZeXDCbJBGffvCvYPSqx2/PCELu+lixYNm4SKQO2uNr9ya/AhF
3Jc5dvH7klILYRoSFpVmydouxdDUtRtRX4vVY3ei5GUxO5ztmkS3rD31rytfabdk
N3HCoOLj+R75bsJZXHni4xh9mfTAtTGARhc/PuKV7YO7ypE4fk+axecwStOK3IYr
iWELB6UaOz8TRi/rREsjUjQ0YHuxCIITXCPYMLgTWBQlT2F/kYGs+N9NzzjZf3vl
e1FBNamk/qJCZYbJOb7zZwCK6PwicH/a4bnNPWW06wDq1zVo0H3T6gL19pEvQbbA
xEFDox0C3voFI48OnlG610AxwifyA1g/WZSrOU47CUaOpSNJULcnicha+OWaVL9s
WXfdYQ+6j17svJ4QEyWc0TwfQeoyIvcgG0pLWrRzYv1xM1CApDb/QZtW2My7mN8G
TweMWXnxFUYQI6K1K3FlTrrPeyKAhwYoKBDobht1OC216RoDMNB802lPplWIZY4J
4VjV+ueUsk0xSdBbqfz0qHlG19wj1NhqVXFxmpkwhj0gZhYSBsGRPqkgWgdhf68k
nIU+AsBdHnHAhgvvmqboFVD0XEPblm43ZP55Ren1CbJhHxiRFHb8rgYhq6K5W6mt
AnqEMtQQzj91HBS1E42F1f8ZGgum/F3PXS29YSr3EBQOU4bho3ziK2QDHomLRryU
6SVWzVw714r7pG3uqIfMrtuZZkgH3palcZZCglUkood9/0l/JBlvsVxbAowGVRHo
hApIGvlZ+pauWFeQZ9wEDYxUmQsDMZ7Ot807JCDhFGnklcgfF/y9rF6Z8l4Sb87z
EccJRuSqoR1MIyeqLQyLKP3VDR77W7hKsHsTSSgYN267soCmHuxTtSJshypY4pjZ
9A29fusjBY8dOBW/QK7aA0fITIE5+173H+SuiKpQD52lw2iOSBzSJQ7p9pXHzDOt
w6zEkeIBqgNjO9tJ18ZaLUgU1G43pja8Pfl9Ru8R7WHaWb5oKjPoGH3dXrH6+wie
p9M/qLCbgG42dExtTBa+V+7dNhS31Hsvk6+XsPRsQHUnYk9hsi0MWrl8vRAeYQaL
yMMcuHOkZssUS2Ke9xpCkjFIq7j0PraxhfhJpf4HxyHCbOWiGYyXvwRR2T4e9vfR
nSyJFIb+OhG0ik+eELUt+5IFOojbwUQrzvp2r+tQVlZ57gqqKkr4Ce6761Pb51l+
DBOOea3W9T3uDdeTwSipyRpa0shcxl0teC9hVgcOFyIPuNHssmErkycIZj/iNhyi
S2JdEUqdEgYat/d+mjEYLqOVFufymZEIcYiqkEjGgaX2rFFQ/1I3cJ0p3VEESDNR
Pv42142BNidzfb10Fp74m8uzBn3bT4ltzFNx3CTjdIYuINxwEgGZGeZogm+VF/DI
G8QFNpbxjp4jp/Fi4binjYLyZ53Sc4kBmEaTinnF8GRcsBtzvaqOtFmaB63sqxfR
s1RrN2fIlmEgRnb3pz8nKDhDS4sFlS57IBtAGBQ7eYYRkF7DhY72YYWE9ugxOUEf
AHdP5YTWjlxEXuhUl1xvUkE7YK69XaGmwg/KV58ePuDVJwDOEMbHXLq0ahx8r1uK
fWqhsy7w/ZNqc/waTG6mGi8U6bgQAAr1dxdLUMLQc5UfInxvzlKA5FyC4CojAXPw
1Qb3twD3mSCD3v4NCkN2TAW7M5QFYL9B9JabXvEKJfpmTbrWYMcjmOTIC1A8nBMW
EQmW9H6lApMNGP6WEAc9C/utORQ7S+w+kSRbWhrpwRHFVmuq4Xe+fX3qcMydCmKq
OCuxiFJWVB9YMj05W/lxGOweHd36CjQtHwHunOql49d2yy+uA4sKwR97fzMjUnjS
x5sh5Ru5CNboOkUdAR8Vfadk7a3fysEmCLG/aQWUbx5pwD/sU4OKzmWrhtJN62bU
6QVCntEhED/Nnppa+AZcBhVoMu6XOJGaBjdZm242rtHct0q8bzIDODwF/YCRJ57+
x79D53mAHqjrMfvhswsfpulCyju29bSrAf2usbpwwLB0a+LERjY+Op6B+Ct9SEoh
ncFt/8kSyDo8w60GdiTNSDu9HIIRqgmWGaKdAlEiJC8amNRzbWjpZzQk7yQWdGmH
985uI9Tg7+VorvJgXMFsFkmV89VQ4t+mWuszgllUc47VQBCdcF9R/4f1ZKIyjmSF
bLpSiEWyP/aj/hjsJWGOPjmGWUrWkFW/sHt0bNC0C9ZMxoct9CgrCdh7wGFRpfSl
wa8KAwT+cjr+3CoDJyOD6FQwapF8AfS+wvdaEWUg0o341o7eZ/rgdTnI5a4bpJpx
aYUb+q9u7fetx6nBiShVyzfdp3FGf2SwMJ+1wfXFY0zsuGatu1FyAbQlqHnRTVTw
n3c8PTj7z2Q2azw/uYSAKIG4dPxQms8us70AJsDMwbllny/9Hdnn8NkA2oArzIeh
0DVeyodujbs7c3IcWonVJnLci/PW/ZDbjW2gQPuQpPbeVMWEezWCXZST/49HqVfC
u5ooz1mJv7kKIFHDEpPL4LoWQzv6ezU8pH5aHfP5rTZ853CIlIetgTgoMXZRwAF3
+8jcaSJ58JjZ7qCVq91rnnrUNihyPcGb9LEmCj1yYrVx94kq0iEAVXiSk6LEvtZv
OyeArCHtyHFNJ1XbvNKEkg7jbAVgNEN37jdRMncaICGbtl3wfYqwI13JVrgw5kLR
+96WG46UcEKDx1ntSrrnaIoLkHOc6WoX41nTTfJR1zGX2XIF/Uz323lWzTiqN8Zm
7cFv/xZYKQOnLr+zOulRa0M/XfKOXQyFmhgd5RgR76BYjXdTPWVSUNj21ZeFhq3H
wSnwGk7DWKd2rGDTuwLVbssepTHl/fLojM/qlwkd60FOhsUQWs9P+rIWUIfuPuwV
PWwPAlbu6W8osX3aNm2XNUKfijUVkPPwsuAWEk55XsjuNSOHg1tv7I3Bq7ERhsYT
dkI4DKCF6nts+K4eDJ83NijeryT3YGZLQckzqKcp+bP/fLDE3R8C3/BRKinIjdX7
daDzBVcibJ3k6LvdTmAWgfx0l5CU19zGdmulrOgVkOSxVNv++4BqC41kr+8w3KWf
ETITSkup0nCgQNBNdmHwcXDgb1YYmnYc7YlHstH0Uo3Da/UvmMTAzcutGuXjvKMP
xhztyP72lsSHOGmklVERRhHe6K7EdW94MdF1UVbXLH+is2qYsIljDjQ0Qyjcqvap
+HvgkOxIOCZIvMgFTIUAeoDPWNLduqZJAqQwzUBm0pu3qZWcqGutvdh8rfbW1sD7
0tFtrg+mwdEV6lGZF+iDG+492udOnw+4XFkTrFUAL4ONJ0/hUQKYjkRwErESJmbC
2CWezs3AC9amkjsSRoEJ+cXYx3PUJ6VgcmQbPonODo5XAAz4sPGGvmHAE8ovfIWs
YXMmDKIjiGFUFlWsku/4DcJtOdnP/6MdUlWuw1ZH4oyon114B7RYB3FN3bQA33p1
XdWOFV9DynrE6ea4pRwuUl1oEvchl4VqzASZ88SgYBgZDpduaPjgvRDbGt+IeMtS
QieD54MwueRgec1egNvI++XhR8tqULo0Ov1A6kPFmv7K/QXplyhLB3lXrf0f2Ttu
ljaUTjDlmmdrpmrO586DTqKxv1+marztkDAS5PtbmW70GdOVV8ZcNkhf9U42rPGY
cHGcLy/FiVpm53XvShc2FNUVkVz+3ezpjGzWJxgLpLTmij5mTNRCRm94TZ54p+/u
dA59gdA0HQhsgjEC17s7oT4VFhxhrtmglXj5Ksh1qhHvnbc8RIWpaQDS6DskYE0V
nxjUtvXRjuPvqm5byX11OEda6rhUXT11duA9rvWa2oq2mN3FEKqgLMNOr7GryWjx
pD3slZhsoYB0CFZ8wU+q+kl89LzSrxFQB7u6nJE2cIPl5HGjjo5K/DhrlR0IH3Yb
BeQl2t6Aw6MNnnL9a6aFLhHfGo49gPGObxTWkLNFQlZgGPw85YmEgK+FcsOJEnRS
LMX9IkBckPcKqv+ut7js78j9CM3RvokY5Vyhk50lpXQ6OixRO3HHgYeP0aodo6oB
r+Vu2tLt//KgAARNRiBV7W5M2QmQ9hmz6wXZYz7Rib0sNbYjxJxKWXhTbyAyVPF2
QFRfFNRCeu9Lk/Vebk42VbX7VUeb1KhsaHnR1eTr/JYXpLBEExamBCZ0YU/uc4y2
Oq324agS3mhL9UPkyjNc6Astbl1vlnc6pa6zt/FOVCsjCG4XxwkOVaXwlRoChhTU
A4ZhJMBmv6jMzp2snklxWt+y9Tr8oUKNcgpuVJF7WgZlG66wDjcO8kPHc1m/Edu2
o9/qx/itAZECAQLrW5wDk2zs9bHEg0qFPiEEYtTbz06YKqTBa36JclXf8E4Zrsus
2zXdydiVKYJ11AEVL7mXaFgg+HUv8HPPZBdhEU4wSP/rQ1Yd+eO/zoBNkU79tbpF
Hs8Wf1J3EtvH87Z0CIlaivtNrXFwl89f3+WMo+Ym18yD+pH2d1hchRq2jXbvG/I0
wwmiX2SV5TfYz2eWBemC50Ky+h3yx/rCuOGP4wgsNQuFlDHjcJIFEfkYNfdMt2oN
otc2tj8wHSywDYpI2YCnQB1VPMHWfkQyMQ6Y9udPqZRuCwvvQNDoKm+FjbQ42KAo
4O3l8ZVuPyKWyTjyNeeN0HcV7hYuFbir2tqe8sqJwwDmQzQgyB7uDw2Hhl7me3+N
5NYl5efmFiXTis/cSn/6nRSm8B9Ucldt9MDT24dTb+yiRIVVmwAX9a6te/kzBfB7
gTEWq66qQZDT4Wpgxq5leTwqOKK6N8L5n1A5nVI0xTu3rz98gsHkKwZ0LoT8ko82
5VQ4MDs+DdV/S/Sm0eUpudPr+2uG8UtX02tG2bOEXg0KQ8PbF5tLJ+pZ1Fk4AFmA
QK2ku4JetnFMJF5cCgtuiqabtePbbDrQjTtBdlFYbqDir41AM3XjYz6LRV7i0TrA
u34KRDsmO9O06VHkzZeDnY0+yQuDhcNSnYnOrZ+85CGOn03UJfI2Qxt4bYvaUJX/
XXo3n0WQKOX8xrmDCol3+3fTfGPcvixpXqU3dK+Zh3+wrs6kSb1gWUssgCR6UUQY
/RPW6vJypcf85aSSVNaNQ8n/kpjIRT5jSH43PWZ5+Bwez6Jd3X6Cjq0jNrkkJo3m
eysV3J0WNjN2jls83DCXU3Lm5xpBQbLxxhHvmevdTsPAaX/7ic/KJaxMoDoKEAbF
F2V2NsKtTsiZuiWLiJLB/54Up3X/aN/GHGcX8BSyz6/5+NmggOIHl87oeGrQZVjF
FV7T+mPu7PBgd5Eh+2IRZpEEXebtry/9MQ3Aq53aDkalzhNYGjeD7/S7BGra1N0k
RkkVaf4BAgcQbVQJgpLQLoGHUFuPdMiZp6w1jo5FnKVUWba3npmQ8IBdYgzTDiwQ
vCvqGW+PmC2lbyO+qW1dTDtvUG1cRS2b67GuN2n3eGDO5/IKwO3hYkTgQ0iaSV0B
K37yKl2sQXtOTXgB7Whd4fmHRQg3pU+glwCZ+uzaBQA6tmZnCt2xDMFIrM86BQzq
b+txjIndrsJUnuoCqeKdxrKW+1AsniM+30LzSmbs/vbAGHX/J2v+7ruogkREdzYr
Tz7zvnLSFTeY3VvB3YaYu58+UgGSIVBnwpHHk2lGGuZ3VHOeZ81qusykNTRyrrqM
9nYt2KKUgdPiPG1E/G16WcnaNT0dDC/ktgCUaM9lsiy3eg1GquA2xG03qj4fb1Zl
HLKxnMoqUa/CN28PjKGJM6LSfQjesan+jA5Q8QehBZnuoU9Xa79LPCXA7HqlxWD0
Vy7sfXpFkoujKyh2+gk2dURivpGHIHTNGGT5awXEfiYb3Hl8BqTr96HP7p8VXJEP
BE2NYrn+ftfvUmPkr0Af6SOW6HTjbJbpdb10uzPaVVAPYPQh0JqdPpzC9Bep00TC
kOHJWrI767o5Sxrsy/DMsD0rcFeLl5Ild3D9z5hvz6WjhB3J7Ee/gM+AJe4Katx3
Fyj8RnDrXrhFZgeV6H68D9imLH0LVZoj46ak96KdWn1hofoQWJsWxq1l2YrQlg5G
jANM/2p+bOlv18DwIl7yEObrZP5d4/faDAB1/+q21+yjDuhxDRT1KJp6EsWbb9Z3
7NPGdKLvDyY8Nh8kU67MjUzrn12jHlRrgRIxtwn6efKufy+a9ebSm3r4HIIim0oX
+jcVoUWBJA0sUBqfMQWA6XMUqxGNQI/x+NVgy4oCqUbyLRbJNN/lS7X9c+SR04Ae
0l3xilh+9hqnS5D6YUX4WAz/dEpupNQgzSuTWb22eScc8Ud8GrvkpiG9uxXRNYz1
TnPysJhOvjeP9iAMbz+lXCXwPrANJlGOx5KVixXFOAedetq2wT4PMNjSo7o/9kM3
UF3ksC+y21kyJr+fqDpS3nljIVcOgFq5RYd+t67900uU32jT/MW4wt0A/FyJAT+E
ODesMXOl/0T4F1LyM4QhtwPGRJOOSI3W1MiwQCIVybyHgseXdbQYxF34UDC1vdnv
lz1/Bro0Lnwc/i4C2/GBCZXCddxfeN0FH7pZJNIk+2MlhWcV/umLNaP/TD0QE13S
cCIx/wV+nRoeMbo2HO1vMcrIGMdhu4hl0KPKE0xIx5991iYfqX+v1Iy6g3Mp5pdV
yoxm7l7A2OKZaPIHxHhg8sUDNdNLIXIg4Mfe56jn+NgtDutG2JBGobHvCuiczHOA
cF23PQgwWGeR5wjmpcD3Eck6Umfaz7osTE97rG0caNmEQQVkc8vOKAgdbdOI5ZxC
K1U/GKat4PL4CLsqsupq6wql/FDvzw8S1wmVh/FwL+w1FdSETzHo641GzThPjUmK
WxI8wumQVON70HEt81cOtsGTPA2y6ZVarFk/AG/cLaLaTaKddnJV9fUOKj4s6S/i
3rr+Ik0YjLtztsjMxL0j9j8Eoq4TyINrnmPsjOvssXMr2YNFdOHapkFmR1vPmjGj
i7Mo2qUfBh/ESY4Msb3wBMvXKTV4PxTMzeLQV/M1wdXb1uhoWuKe5pLvcIsmkDbg
6KHnDIaUikXxVXCREQBkdhghtmEBp+jIcKQ0GE4y7QSZDkUa19WBf1JiItEXFKgf
cDiaUzXMqJUzsmiMtPZqs8YNpEG/O9BZXO7i1HdzSVSRkbNGX0CdipNKLHDcsDYu
nYyWOSCRLZ9tCuqmjF+iBnUvTq+Va67MqWdqyz+QBXtOYopu75dAvlfPZcPYyBGF
NFqpKExGerdA7xS3e2PiGWykQD/lvl9Ldt0+CNUurFMT8NSFJ/V7UxMEz/4D1/nh
bfXaFUjtW52V+jIFeyO6m1kgzbnLdCtxb+TLvVlpoj5bNTwsVQ7cl/TvinoFDKw+
AW/L+f60hhVPvSTAu30xbdc72EgWzCB4P9MGF2jogkasbbIFHNz4PqzlAIbbLGv0
2YwAunF8cgvtCqJzkgYZ9dB4xL7aau2OUezSUZyelAA1sHjyrmp8SxoPjGXkgVzD
NG9/mQLhWlN6bL+Q3hvc46YId6oZmjOFt1gnfPCINlKzUhgqw6pK3HwD9lSNgmL+
ELuLtXtljmSXgrZLzqRhXQBoFzydogRIodwr8yjdOttkHo9E7Ysh00tTfHgR0gvk
D8jlvZFwWOE2gTnptNrWLYPyLjFGOaPx+aRx9phLLbye7S6fMVi3+5fPrP/ZcYey
bz9atgFMW73kuhbbwoN7/lzvR2Bb7S7iS7En2Ol7Vp1Tn0n6yoTO+w2WWuiXENHN
6B/it4+/w6yNiuaN36OzUuS44QwHjcvCMUv8hKEjhDydvcoELpnXyy54+HKDXxdT
kzeC8g8jR8sSCiOSLzdj3pt3PxRTxYVykrRa+isImxbIhzpa378l8/HAQbwOTLUh
WRUcG3LWe9lOdq278DZzOg7ovEDln72DkxG88nGBqTdDgdELAYYCVkXaivEn/MTu
l69PGhpA/sRX0e/7xCnfICtnEpqTHWsxKE3oUbaD8YTYbk8Tux4GMek51Md0C1g1
Qxk/fK+kAbthSVrt3gFXChgZWhIS3ccHdNkYsT8EcvIQPfRQNKBCmkZc0wMAZH7F
qqnLHkrUIsXmdXz27FADxCOrR8db8SIMAPSAUCniM9Q7WkWISTYcaaDzmz7yeIx1
2YFVclTKSIwwkK68GYZYC7p6jv/NsFqS709KjOJU54k4DSexh/EVIuewgbDzoAC5
V6r8dVv82GmEIlObIr5IUEnUmOYy1GXR7wIvfM2MplqRdrLd44Xu6znL8ZEXy+Bq
EocHxKp8NFPqGggLOjADvoXvo2WFwZQ5u4zB3kNoIhrW5hgfNA5qMN9F1So6sdd2
p8RQGit9DVxQ9xpNEe8XToAeruoCGxTse2UaPMdOalK1chQBTPxDSQio2xUSb9VX
9a4avvr/4IZsmaY/Xi3gzuUVgsqF3dFiodJfWQqYYKjNuUxQgz1Jdp6C/ysnZByk
f4cVkOHJhkWbzr45XTlX124MzALLS1Spun9Yp7tZJmv1l3ovsEFr9Tp3Kfq0E7Ug
cxa9P4Ndue/t7oMM022zOUMiEJB7y677F3yOZ2/qPFkFFbQp1mclVSAXTYkE+6BY
olFCro1c/63p2TWMbT1B7Eza9LnkainsnqnkTndOhDnzklPv6nGDM2u2k44+i5Cf
QSxzAFwb+hrGAzB3P6mR9uhyxaAtuuEzLlV6uKNgsGgGUb647vJ4JXXuR+cqt72l
v8JlNBiX/kDtyykTBoT8aMvv+8lYhHH5JAFKHaOZ89ilqf4afkO2xz1IlBVP3eI4
4N+yV+2aub5y1WRPTpvYD6sYw9NA/JN5ej2QUMy+Uz7xO3iE9sGICZXWW9iSmiLq
fVwewFYnWdIrsszrH4xJZIzf5UJH0n0+nrqkN/bY4OuzUQTiSg54yA4BrcXYKVSW
8el4UkyN+J+qdeTFhRIoXk0h0jNsBJAD9+6uy5HSz7ZXcYLoKVzG5YdotWKst2Dj
ASfsNCOwBVwUrnd5MmA66ptQ655OsRt8Vfax7kIDWwHMjFRKPH7eO9xYNMzgxX2s
rgtUE4mOWOS/g5Baf/kJu0Hbq0f2LP+oj3TiEGJ1zGfbNhRpF+UdcG6gDHWky3Gr
Md6JhZyyfqiHT3+U7vBp2bJAd6K/1UdyvTA8AiTupb1Krapt7il+ws0w2GBTVbSM
g7CPRKP9F6h62m20k6AHpmTvCl6nrWlQBbAOo//CzfAAdGl8oha8XWvSKnDGGlTz
MeRBeJdrpc2vjqBCgp7E/584B/lGYsNjbcytdDqo9Vko2qEDQOITmZc0KO/QFDCC
RArfO85LPfLV8KGPZHurq4iqgIxcmleR3L9Kl02BjaPmSxz17Epitbx6I7Xk0Fkb
XJunXeyIZ0u/eevj8ebxzkySLqva16J43J78TRv9sm0/nc5YtAplwrxz0PHnkWga
1PkY2nN2YO/r4olFbXuwhy6Dg8OkPq1OK8x/AhWui1pm8cFiRabds2U9yFnFrP/n
ZXTOriiaE9DGRFXjdM2EjpROLiSAwlCrLQ2hJJlWO6R2vf3htDa7Tbes1r7jUxya
1RLYDVSgKuOxeVxeHifRLf2YhVVGmX/web8R+o3R+zWpZo/mLmX9eS/9OGKE2LS1
se8asMoTB9wFmprwkle/Q97i+07alTU63mFYtwaBpMSnjsPZMSJuXcqfak4fj4hu
O0Zww48aQgd1eXDo3rQew7FMnnUS8b49VqI93tbkjWjTcNUOOFgnA04FjVG4f+YQ
44qX8L0zJCmI3JVmBBSPSzlOpBs3Q64FxpNScQj0jvfomkBSNpDsLDnhdiuzE10I
6F18btzCG3w3MwwMsF6l0Cbh6gJYxT1oC4PEeiYs7VgQqS8DApyz6BLpSaVreix/
djzPDwmvCIFntsT/UE7ddoIx5LsEs5FJZKmzmhbjgWzuGBIApfqn/Ef73b38Z8S8
7JXs/xMuSp2+tRIsT9B4K94iTMamazBKu8bC1tclRtkLDPFTv806XCYMmcbsxORw
juFFLjcBKa0ulq9Q5O0rSHymn43KnQ5lB6/1svjjbUC8a8YhAPK5oKiH6RZ2wahb
GUI9ATc2vyECtIMOF4kziR5lmanwfvUBu0xE1GWa9skRXYzOS47pE7htnem2KNdj
49IOpjaLvMYyimTf2nnBO24UqPG8T1qSbfyrihWVeLl9EwrEoyE1vdCyrJS+oHLP
z0qRHu2Ey2fSSmEk3C/M784EAjxMz7f1yExM9/QthbCbjAjBRXlOX0qVPt8iOnJ4
vuNRi2WUZHM8LCQmzSvqGYvWZmYtcRhQA8aQyvP46ctfGdKR9E/pnOJH7gHS7j5a
hquWR5zNnPvyeAKiPNyPkDbQaZVm9sEBo0rcGMUBzpRt4twMDv1NTa9dlgYExmvR
M3OxgaidSrTZpswcv3Y8ugIP/xhUAeJ4lsrrTs0vYHcQwhNLsxeKU6ukhhke/UHO
PD+inx+1TIJFFo5CWS1UMF/PJU8LTCr7U/S+2zlByRnkGnICaq4Ddaa5oI6QFYPe
CK/LDsJfHRGeo2LqdT3ElFgrNZHFzNMQy9QqOk4fYWXmYRdVAQHGjaCFdkZQZw6O
p4b1yjsQGEmouWPB23Q6njwYcNFa5340uB1qys2ThIefH8JCKMyM1clIg11+layO
wS8y6+ziHNWC1Hu4Q8TnSnp/r0E/+vFKC6Rc/Hn02UIJC4/BMsGoBIFqrDWBmGRv
UhtFNp9b2WjR3r4NgdgiCoD4TWZ/6ZFsvpSVUElovz6FcFQnzebamdui2+AWDLKA
UIGpytvoMUxC9LK9b/XpGt/8Nvh6/qZQTWkprTECFgfZI/MHNrjyJzDeF45JnpIe
eGITlOGJaEu7H1/oVXBFOdrQrUzUGyqXgp+XUnKgLo1AFue8X6cZ2NPWxOs5WI8m
etUcxu14ejpCOrTh61qmaiLcOO8u/zxfbCK0e89zXdxX4yhTQgq7mVV0bo3KKUq4
0h0p88ZUaXqYgw1T5jMsTMwaX8WYlPyT5EkX80pNEzeDIShTW5DQ4PHwH3XQJgY1
YK/+emHvjDQe8tCFOWsoa/0iO1ptJS1yxaqtlaRuU5s/ooS9H1GE8ycbOxvGOb7J
nlxI7utEl8o3PTiysLpGRUhnaIoKNyRI1Sj0WDo0mpLlJJS5S9Jr0QPTS7hpRFu3
qa2HUS6214OQM+113krHFI2lBDRLgWIclEYkNjKysFOyPf935+z3VCr8EQi+Sor3
ijaOwRR/yl1fKH+1Bfwf+m/w5VVF+hHzyVl0Lvtd0PCS18nq8//xdkpsyUTTpJJe
QMl7sc87JydoTCD5AyQlj/LjvMTzLwuoZJpWArXH903BOY31lyl8XznqZZzZFT0u
H0K/7c8GEiw+xXPNzhAL+RtXhwzXi2hF7Y6rLXrBcH7H7QqGIggIo7jBezVEC/KS
fHurUSVZ37Cq41DUaiv1g3ljOlS05qWOPR0A9F6iFDaTBu5jJEfUAVEBQFFeHqFc
fqhjQL8jfvhsqhfPY4LFWfwrU4VuRbLWzx+HbvfDP923/B1VWGECOS1NvIPUmdal
kfb3P5x8B6iCGk2Sx9l2dQg+9Ht0v/jsNX41AOlJG5fIlnWF4ZbnoXI6QmK4hPK7
VqHkjoXxBMcrfJIZKobmXQ4w8Ci5t+Bc7XdrwpIZdbIBMW1Vi+glCXxgEDJPmL+C
O0P4I8jo4qkLOC2GlXe3tZuLi+3fHuSzPjKiteTNqVDe+NZ7iRbdNS7Bbv2NgJvA
6Jq7eTeLofftPaloI/H+nviNNvZUtvtw5RumF+8lSfR2PEd5tOixPBLjpZOu9joK
oi9k+3rYvmqJFn/+OJE9QuivxRUaGBGrPyKWexaa831SHAPIwrQ0Gt8drbJkr8eT
pl12wnm8boE9m7bGlcU1Mj1CHBYz1SpcCwFPsHZLo5dLrJm2xTUyfbXjOBCnyqrn
LMkbrPq+yvc9xKyreMXhz4q3vGvt3ECGqKSgFLVOFAQL6l/ziUFNm/N0rHl0n3Tm
+WUiP8Oqpw25bhdocUZ/1jLMgrTzfsxuGqJr8yLCRLEDnRWOa/nmU/pRerVKMcxt
UofW7r00Cg7vVLpvItCoZoXLG0rn/PcmIo7Kp7KrkMTRT10kQOnD6c8Y1T4Upjv7
Yo6UWQjGsSCbIAz+DYbxbe40qKF46uDQpMPs1lgUsK82Y4Nk4Iec+BzytqwciyVb
lKyBCIQoU9ByuU+9Jafd6sIL6oJ/RDuhlVoDkQ7ehMF3uaNAJTJUjIwDVs/1ZJua
UovPkqkiSIl0Z18Eg4/YoCK4kT76fFwUEUtXiuqAVTAsman9gJ27f/khmTkK9zif
Qg0c4b0IUq9DHywMDokN/yD0SBzOrFWgkbf7Az/uPVUGZFhh++0mpZQYHC2wisxH
dZxMig16kuVeFUbWPwt9O+7SWSVU3eVRkADQztp8f8YhVwyHiDw58kSZHiZzyN8j
9s8jbfd3yVMFjOCmTJmffHcpibBAo9JzZ7G3OOBS/Fjpi/8mK/O4C/3lgEcL1WhE
7ScGjRWMEZtyrDL4qH+JqITdaxnwiL1L6vglQq6XsmpsOf9EEYEb9ghb8CtutNJB
QDgOp2wB5bBQ47i+XUHLpK1PZi8gHWU0Lv1YA9/f6SY+GK3K8xd2qQ71vJhl/6vl
d5qmgpXMq6dsc/2WwqI66QreSW8MB5U+2gRE9LyYcpWng6QANF6HqivSxdRbxMG2
HJw58SSKrIqL4KU5VkS9/voTxy78TPxN/6lbgpSbo3MowKT1YIH2FELCH42hMygE
cYgII7gT3W2SgrOyFCg7v7BAVp+lvf9MAxuO+fUZgcFkGG6J03D4Cl11yjWaZgMj
WRBz6eRmm5PR/bI9DxnI3IUTB+CNgWrhcdEYdy2mEJeRG8oF4/bTxiF2unvOvnnY
PTztxhBrIdQR1QDCmcsfLsxDKqHzlMbXi2Uk45o4SYO0ktfJN5YmTvGUlraQtv9o
nKJfVGLghSafKtSQ1qg9TfuZiCYuCTkryjORGSrLCXZ3ahix0sDc7NmsDzlc2IAU
giwD3nDdmawlR78W7g/0/fLRY9ryKdwwHFaDVI5Ib3ODRHgaoFmXhOj9oZEvJnKF
Sc3NqG1N66E7cqVPBFKvOerIEop2aTMPFWPJiFXNxWpBXSuBa87fwhORoDQr136c
NmkEGCaTQq5Y731TbezeE6EYqYl/U0zmIjm/MSvTzFqmenJ0TJsr+BGIWazC5Y+5
ZIKwxhykCKTJOggysO1w00cH0vS8g0VSuijrl8GeyFi9RccWrqgDZsMVNM/lya33
FlvtBpWiJZbFxKLzVYmho/heMKHCqb5Qvv1A/DozG382cvYibKhZa1+dbY2JY7s2
GUCFG6ogLRPcz1TGGyFWV7wcWSLMmjkiogSW01LAlyA0A2yy4Y6zabVfFIfjJ2Pt
kbJvN7gcMfHdZyiV9TdViTfygPfJB3XDk8ZbjbqLZkD5DkYbhPu1I9ITR7YpBO8H
yqD+CYFlMm6tYae8sZyqKdahmaLg0QpHifea/4aRPt6khtDF5nYvxo8SyIyYXJf0
Xxx439kCjWAJzgzVeJFN6d8BtCqJ4Lb3xAQNa4P/ZEyGmlWlDlR7J9PRw0Q55Xjr
jCrRnpdUtC0ECDWUtERkHWpaBnGl1CabfrrnGmbwkRw0pHoGgeehNGzUbfs2gIkS
Uo42WtRL6RqrYzSh1rzIM2twmF63n3mdNfX51O6zLPODY1h0tC+Iu4IZGnAAlRpE
xcOXpS73zkfjt7X7cAFX0CCqfO1HwYCZgKOUqGBKlfK4TADoIDXvx1PYtDuFKZaJ
bd1vhHDRy2h9jSK72QUR1l9xsN805MGtBLaBFQI+0lABn49zSiygf+osn/OSLXih
GL4uJ3LpRSUpfeVlsrk4oXmU6hZdtsju9TRlnpCSs2d2isxt14rN1ytS2TALpqLu
hvDpIoYGkXU9I1e+LBvUyKniPuaQGTbuJ6DmdcqGQxY+75a+gIW8oaoCrGOk9wrw
7Rz7PPoCzQ+Ll+VNfg9AUSyL1WUmJzy2XqXzFtw/8Jbj4NOL2r10z8vw+AIdU1YG
JSCgcHba4vrxUXjTdCDmzu3265haehp3zRKA85Hv9461NyPyGGJ/wXL4Ujn8n0iU
F5bAYiyCDjjuSxe9G8fdbNerkAFlqUqDFnmUEjFnjKF+f471bFhWL1SVHd83jV7p
CkJsltB06i1gnDWissqjXh4JbKT5XSxGWVPyExVHISjYXGPHX6z/Z00V9/eFUVqW
0HeHraE9uAHf8nrdjHeu66CgkWOzbmyWfVtHvZTpk8IdQbahAVTzsNxYKbzFOmQO
Sp5FYmpCcOBFXwli/XCRN5JF92UsnxCHlW4PrW9EdeuuOWlEOK9aj5FqACvnB8OL
YWNDxuKmF+O4KGI2/2na8uBmCPywg65gp+26gMqohZ5uQS7GehzosDAA/zPw3sbl
PipHotXa2AB4XdWVon91URNzvyphicQqKmU1yg0SMrBMbtaStDzCS6CgYoWJiHyx
fjF2+Os8hxlGOloC0pP26i+1TbBoFXlZpKvVnV01bLmkCmkV9gfdRusgES32PS/U
dWedsREvxG514ACKApsBhO+jOcMXUhkMXj/XVmv3JnGKNtfuJlSCAROnTAVkSPdp
29LETId61Dt5Ltuzswx1ZJ3jHqj0d+7qiSaFef0yIdGBmxznH9d+Z+DSavCfYJg5
g2yVz+0WMw00ObxUgrwt2z36l8jA45V/rmir+q4HegRz1rSUSXt4+FIpNduZABR4
p7dIEbKcazSE8eSecKybpWpijqIDKbrNAn9avOhdH3R+gRO9yNu3I2FAL8jV4Psv
Qlwk6zJnhkaRR76ayiT+s+9BeUtTERpIkt8HlhyTI9+wuDCsez3EpQ+uCsBTrWiN
C+U8pwmyNzX3s0lsms9mpdobKHBorHqlTfDF1y6ND+OqeXwX2+4rtaCv4yvNvsVP
4N/DRQRxVQ4VJhLOkq6sDKcqIHg2i3p6SJQ7pU/j+9LfMg4bgV7PtiqqBty7mFOS
FSVM1wpzbc+QVuf+W8gbOx+r/L5+MGL2TSXMkmVsW0k3K7V9saV0yZELx0ljcX3F
eAd2NNozzl5Y7hapZOaoOO/+qX5ReztNSjgxhhHoEfodzizPGUNy5ROf6utxS0Pq
WOorjWuHiipaYchvQitusC7OGu9aMIvNsQtYUUT02X04pio8yIwN7zVCCMZPlGsy
87gYYt53+Qzjs3D27DcgZL9YU6898l8QrVm3G6i2qUzi44KtglSJgb5f3oTYKec6
nXsifXtF/qJGTD7cNskdIhX7qxJG0Ackh/ZbPEnxLL6j+82NDnSSWr4RuXqpDkGn
PBM9bvMH39kF/uUy0Mp4ZieqdfCcn1Ca1V7IQyd+bKP4M8UjWyFBLQuTCHEm1POB
PFSUtouZD7oPIl/7jRq2KyXQQE/WlKgHn8JwWm5YMJEvQS4Ru/gNQBtmrieOWng7
K0GzcFsx5Ow/elkHRORNH+YBFub/wHnK8+x2siTFyhoUfecy+wAL5IN2bHGJJ6iT
DKQ5XxzfRt9nTg0sBT5pF0BTgdXTfJqTehB/qg7xrxuv5bZoPOHm1h4DdnsbZkxH
M0v0+McreIMj3ovt1eLToaPrDUWzAEcQyOsO5lOrZA8gtdBKWDOWibI3CsG6MtBl
fE8SzqzDsaK+7/O37AVQGOmuaR47kHY8aDQ5laxozR9qNTfkASazdYrmaWMpSRTw
7wuw0qrF+c0swErSTTj0gOBnJI4pAQbqwyIkLkZnaobaL4idibBfFPVx28p9bNI4
QFC2/LJJgf72NYf6ZC7b11lD4kSdXmrDZJBIcgs2mZm5aUhxLaZjleZ9a6KQEtIU
9pkFg/uvMLdSLoOp3PCbLXlUbSIiYL7ahIDOyue7ssnhlxmO/3eNGiWfrq3DBERX
5dcicWL/rYX/buewFqiGyHlGhty2RezIgqlEL5NfLK8ZGSmhBVRXMlQjDscUMsqm
oszNMlox9+vtZyeeUKuG4l/yd+jE/jTerqD3BloFd2jPqMkG3iVzKbERY1STwB6Z
nC1czAQX1DGtsTk0iJLJeDr2eGsl7/Wsmhx+JRELEcz4Ea3/yb7R8z7LGivJyaxU
ZGMeqeskq/JyJ/ayaHLGWBQTMnSRXPMxOp3bam9SNYmDwFAgFg0og0fviMomBovW
j+C8N+c30HqRVkU5UlGo1Em6IRkUI46W98DKVLri3ml7xHYA82vwXoSk3FY8Q5ws
x9EeTkn0uK4D/WS/RTAbqvsHjtXPCdoz9siynpH2ycFsz9r4/csIcf6yvCr0/DgZ
VqAELKSgTRIQpogwspGDNfFZVbFq98QuC8Z4+4PIzm3jxLCBgEYWveeswdKZJj2v
B50CV17wf+ZvbYViE5pcEcsz81i5n6EouL4+hopAMB7hrRKt+QfITkTTWAXIF2MK
Z73o0Oj27nncO9SEVZj+EZaKi2y+qL+0320s9BiCCn+UZslopQGBPI1Oa0KKBq6Y
UeY9xSOBHga3V7WHODbkPmhEvbaNrKwvYn+/uU34vxJmMD4/S+y32AIPl81D8k9J
KrAO9257M9CYXQr6jsvlB8Cpj459NY1vKPMJ9u8UwZIL2ePB5n6J2bDZEZDNP+jc
B662lUTCxXgFb9pCTnCyvlfYrvYHOL84DXI2J6Fr6RhhlJYn92ZVkQdfKLB5SU3j
JtBmVfOY1AwJZPcj//bveBnm2wpO6IKJ/YXkDOGGl6xF1DpRcgo+CoeVd6lRjy8A
eiFzxAOMY699ZB2IcD4CVLJVdYN0tobk4z9yLEs2a9uGYlueI654IBX+dxOoy/rJ
4XhE2ghZ0VwUrzhczjdrVg+0s1YoU3auKcW5DWzs7FVemhUJ6b56giHLKib+pByM
euPOsSEAHcSSXSx0e3Ckl9ndDc8nUkmB348R72Eaz7Yv5E9HQdWPZ2R1eDzT7Rl4
5azVInuo389l9KJ1DP/uNV0IwMMblhrQ1aXaYIXwmzZ2OB6fFKM93mkgSVm5TyTr
pwSlQSGKmpdkG2jZtgj2JFz4S9AfZtv3BlfeW/+FU9wzxTNkeoMkfdZosxH7aROj
QDr79p0KcO+KmkhIuW8o5hlGHn22xTyyxFug5ErPgSgO0vkBR97B2gcpjbhWel2m
7JSPU0/prFLb/7qwJ1bMHI9ce11/onUlossJ3uVlexnTqVi1aRxnbgapWqmBvCRH
J9fs9rZ4dJ3cfdu6FV8LoVXgOrBN8DhHOBvbsJKRwJmrS9Hd5+7gZOOfBEdfsTcp
4fHGJ9ZR+O805oHJzu5qsxe6LZPDDu3z48QLzjscuXlF7Ny1eJhAUzC3x1MpxbhR
mTOUkXs/TcYZSFOGMaZBCr8n+FFhhsl4wqi8J+74zQAN2OziBJlFh8NVoyGLpa2G
uEkC1Mxo3isnU3YXCnlSd2BBLQ0b/KJLDFHktJR9sz/sru6375y8bmcMlF8f29d8
zWC5XnSYWDn3FyasMub140BVuQ2O0iAiZrU4oQMPJpGanf1VZB/zaw8FCKJfOwB7
zfLrvuiOGMZAnEembBhXdZOE7exIwke+ExQyHyA+Xcmu1qy27Kqn6xEhzer/afNS
TWc/0JWEZowoBvyVKwYgaIQw4OviATBQoMPYXr0zuirXiQcW7fCWvT29jB3CjvkN
x+ZKZZRlbBnweCRbThi9d5OLT0ndxIHrAgDuP5Wt1UgbOEfOa6JQqWI24euLCOFP
kmruFYR0OdP1DQdGGs8Nr3Ddh4EsxnYsHEHVuKHcmo/77sUfweLU22WBg2DXnVo1
Bx6QV2wC3uAQuTzjYsnNmn+4/BlkY79wyZfaJw3nZjTztKiuEJ9I7XCt0ASSfPXh
6lCVDCvzotKS3lUsB/JpRZmnYQ3UEuj8QBfJjIu5YZlYWY5bVsr4DduCbEgQ21L/
F6aP0OAh85WYrjPLBg42snJHIFa+RTxaxGiW5k7spQ7kLxqjBV4xwxNLncZH6iVH
/PRYCmwau9L08/5QhH8QPad2bXvklF3HitS4cZZRw2VcJoTplMONzTXtYf7C0hZw
+vyejps/7+EP9TeBQIjYpQ4jkz/8EKBmD7PLteeMzaDTStvxRhL/0tEsVteYPsLu
PaHN1n5hKO2lS9GSxhMpz+6ImdKAZmDvsDHTbAjxMwaYieoP7mMLWOaQSYNiF4ja
P127GElE5BmjUjH+L0oUmvRyReLG17MAoywfTc7myJSONOeLJLdt2LPkl5Fs8xG+
soy7f8zongCgrNpiK/y8EriztjJ9vXz7M2TW7XZNLbS63dJQQGhPZzVMMAxxaLfA
ZfRbwSx/x/iXt5jiNdRpOS4XJiP174+PscVBWyq9GJJBSX5V7bEPu+04Fu1iuZd9
C9j738/rQgQYwZbg+pmvaG4x1tiNXA2o0uSj32UDz00IAmE/+jHUZ1ayoeMXxJT6
rrQdDdFoT0QLP1EDKNtAm34FVyw+lNLXs1BkOH5rT3jLk1KOeOwjLDRvj9dX8e34
hmxQaM5lgkRO2RwvmBAIUQFdA/0smfigtQBCNxlsCcQDdNNRehOdcxH9kVBvsj73
GCD1Ue0ZvTv/WUIxlnmkPSIAejClGUrRPFm4ebiOG3wqKxb0OgKMVJpjg0MgLj8j
9Mu7jiZI9+FDjskSaaegbJVvOxdlCy0+MTUprlDyaIU0Qnk403ndDrhfq+4vg7fc
SZqsygGiBp26ZnMlCAOZBnBbqqA80M9XtuEsAoDy7dgPx1a/TGDdM/EIeRj9LzX4
TozAoiASokxSPw/4wMukNRMqy38ZRxizoZLBrr/T4jN6LVUtMqd60VbIJhjLIzAw
bbUt5fBqLwRo1z0uT1eNOgFyRa+tU9BwpLimJloK3je9B82P8M5dWdj/vD9UT8Uz
VEBKJyjfENMES3+oC7yLCALs0DXZJ5hPvn3Ml1niNfay69RZDoRrkTErQVkhsyln
VkmbJZ3kGUJ3EDE0D5Nrbds2mBicBv1rtvprSxEmlnHNCuVzxBfEmf5ka6LDRilp
/5AeP+cEr/RwNLeIpKeeL22tZzrJ3WDc/Y+Q6MgG893KXSx/ql4k2nYIZRydr9IE
3YmnREiEcL+NloUDerFtSPsAdwGXtS8Zk4mwS7Q0cATRS0uUa2cZt1B6WhD5AoK3
ma9Qd1ah13Cji878w/xcjCHzYUcb59VBDbwwIcdk8+ZPCVF9ucCw9xDK+wTo73kq
dDKA/bC+yEFYuobZtZe76wJ0GSLAXsgdgbSc2UzkIOfSUrjflKfxOf/EsTIM5D/z
i/ykUt8l6LsrxW/w7iMC/JmrqrIhe0NoQDWPWUFjK1RjHGco3ZAn6sR5RNB95JvJ
VomvMkLNbphGOpSXLhtiWDuJ2y5zp4jqOA5df/SRdADo811/hq5YN2OoGILJGHPv
jClM6+VJVbqpRCZ70g6m83X0DON4X+EjeJwJYa/vlao20NCsfnyynKD+NTpl37zh
wUW1QRSStRIdzmRfqge420sXGQToAy8mi4mrNhqOX33PUjU3Jfzj1I9a5MswFpG2
CQ7accvINLYYvxgJIJQt7fOxCApMMEv6KCUChen1ueXNji6u1P2VAuq3uVUjtVFf
9z3UYJwRpdX2ZHgFIbHRcmHnMtq3QjuDl93TqZRscG01YDtCJrKmq36bpqaWPryr
wUHt12kFcPWbIbjFJF5yH8YdWvIsWBswunWit1wkP0nnbIVpDFNyC47KzQJOdDJg
xasbQdDX3YhNmbcjRS9jMaWMfW85/K1FJoWuczgD/hq4l1K0IHpGd70iwP1W2RCi
ouPb9yH7H19luPLqTx9zA2hFOkZWw8EGJSHSIbF9mHq95J5omWfG01F405rx4c/o
Ej+6y+hyhv6hOvf7UsnbOBwvYXjE2MQ90Xg09SA8rJG8em0RP73ZcrJRZn4u79SJ
aPrqiHzBgUfYPQYbZqbTX0r14sgl7SX8Rc8HrcrrUL/+QkwaJIpuHbdl+EWjBmk3
Mk53pIGVv0FCzXUNv4dCn4DqyJcCUATF54IRmnPty6WO1baDUqWMypa+jtv/0Dx/
MPrHUPMdWfhrsxuyyPBidUqO7szvPZkzpNJa3FT2X63Be+KeIrJtBgS2ZxmKb3PW
rTolIxQ3nsMIFWx+/Mp3a3vMub6ifFLkZDBukOfnogdITGCGcoCyLTEli9Ag3gpd
hW6DSX0agNY1crA9BkHJRwoAE+8MA2rC3BUo2Q3SS4qdcTOWyh8fkkNwLuI21PZX
P4SDDsCeFX3QBqVi1Y+kIT8scLkot+GwanbloWWFObwJXlJvh+Ato99KN8HZA0Sj
mO9vYEXmRGXsCuOP26TP6/VQL6Fy/3KfvFW0x51SBbQQ7u+tJkYKz8wU/EigZtOS
Y+w9IKYXN+cs43ZjMe6oYvm6zcGYNm14RQrGkMmkJVv34mRlFluNBZcHR6SMr40e
g05C/VKPAzurV0vbpxeLmuunBWRYs+ULJiTwGQgMWg+W4P551bCYaNfzWnUL08J/
f/6k58Gch48q9faNQEb7/fAXAKqKIAUqpYxPnCXyT9Uygq2uixTQSA7hJF9jc408
yIqphxp0b2EM9cl2B72EjFoG1G0kMgxmM/R1qX9eLlTxJkye1PloVMGQpXThqAmI
1+WOz+ds66JdxuEa2I/qgyi9wNDFauLCzWL+JdYFaNG3fBvaxFEBiwo4GDo8Wa7t
KKSCpYT/JsNWijgpABLbstub+kpBys1OWkIw9jOSk17LHKkOLyz7Igs3AbEYLfqM
Qvib9t3iAdt5MqitTXX+neyTAnC6glRWLXgsgzVPAg17UWIJs+C9rw4qQuBZJ3Xy
vCoQmf56Lar7rRzWztIq8P/X6T6U6yfIVwU8H1xtWO2PtM6hMyqZE2zlYfAHEXbM
DyMp7yRY8O2+Zu5QIZtVDTFCPunuiC4nBDr8aO0foNQrEtdZsPziCJYO0TZJTNT1
d1Ela+TS109yNprzKfPlp4liTqDfISFqzM9Xujiczhe3ZMWNSAGitNbhzV/ae9JR
QCv09nMEhbfE5Sl/vppf+d6NuGzfXjlZGQVgrZxCW/f4Vd+OMzc6jTZFqjaftz+S
wqAyM+aGrlBdOO/2lc0AWlZ1uA6PcMjkhb0/6tKLKZltP8rPJTgVBfqjgjI+Dnob
/Wv6WfTlvrU1I8luKjXP87GNmZCqV719/tMnMDBoLx2Zzx2ij7DsuXhXRz7bEUIV
VlHK35gmmuvLBIPn5FXvsu0zvhpRGjCMQ3ZoQYuS1NyRdDqQO2VO/H3LvvZXF/P+
1oNwr6FPm2Ib1VPHMoPBB9XbERfDCY1homtw30fdZoUIZPK92kjF42Vmx9BGDQbA
kztFT3EedE014sUUWJ90SwN1LZKyD1faa8UtpzqMRy16BwUEoHe1e6QkoGjAfE4n
pvuoK90TvIghpS0+wsclSKep1delFjU2vqDypoIcuCJ8v7cw03ads6W8rchtgtOk
m8cSf7BXNqplomJgMbSQFJHNb385jqCZzhH1sZrc6SI6rJnt3SDXn9fgUkyjpwEt
MiZ6+D5ILlRMM5dR6R5VIJXnrk9jTyX9QOOpi7eF6+pSZRUOr1h34k1nlEOvNo6M
4Exj3tc1UhafY0Fkqy6RnHPMa8XFP3eCTzaBe6kDzaiAwG46FYf+duk5C1UPA/Af
tm8g7TYfnG46IiXrtAyoxkJOblk6EuWqXmUDOw0PMhNdn2hRsoQhao2CPNqRuhZD
oP9E3+Pz6/OKAi+CpzzdJRlemcfcM7DTJxhpH2FaR2/DMCN8NrZEQeGfrlOqQERW
OMJCtgqbD1N6YYVP4xi8Jf8ygxrm/hb1Ur48bCo1ff3HnCTfCD7j+aVPktgt4rak
sUfbOh0mYBIWyPKf1/LuJeXoeFR4s+hTkcWtQrx62wNT9KkO3OOaSqGKuUmInB99
LWHsdK7sxPHZZ8ez/6Sgy1XjMK7JbvnrNtSUaMnjicA1+otA0VVLbimg1hVgRGhh
0sN6ZGWXsM9g6p09omAq61iAfUKfj8+F5EoeSp8BV5QGenBhIW4HGRGnD9tA3mKk
vh/Ri8Axrwcn7Ge3GWu9Dv7w7vFLVDSMp8m/j1SHkgXU5fQmgDvXW/PACUowg9Q/
0/SP1w/gkANPOcEfKLI1BwCC8vmMLjMZYuk3XhF9Al1JvEQNfrZFN6qMYETj+8Uz
ui/GFkvlDHmom9lcl33k8u9FE6zxanl0eMPigKu8Rr619yNmzbQ/N0+6TFJDms06
AdAaXK46ITXK6KuJlCA4QA6c6JKFLhuc5uYUzWLQI1bKV9Q6FifbDIocPd2CEXDl
iL9NPX8o88grK+eAwHulprQOF3sH2t/TVU72isM9dHDIWVpxQofXwRb8Kvh0wrod
OOv20F2BbY4B2i1PQoVkgzaM4WCIssSPCxiGpvgcHIBolfbM6dlVZhNNnuQsaiiM
LuM75Lpoeswkz+s3BXsKsQeEYoioQoDn0P7sHEW4o154rG9dn6gjsuwlsk46Jx23
3g1sFZlsnnVtVKZpRci2xzzpGm8ywk5UF/yR19q/0z2LDpz8qk97TITC8zBwhaeL
mbmz9+X2sOaqH/9b5lbwn+RnTK8yhY3XfWFYhUFDkYToiNEJxR5+qNOiqkUwiY1X
n2M90OieI8fZ5ZvRJ8UH7WhRZ5GkeTjM2VyvRJMaub4jGx0QNW+IMTYVPQQWvJc0
vsIhLOEKL+/ttWXmn+RDcBNBhYIKFe5DAMvDG9fyuWs+e0wSbVxuy1KllL+zUVax
VdDGMUHfE6WErExRjGgDv+HvbEYm5tX/ZCQqIdVnOuVPAkjYVg6gf+DVzxH8pMic
rvS41QVfwSk2hrghQ6GVWfTk5qNWWs5reofoCc1dDpbhjGqm2YPWtOwUM33HN84D
i8yT88mBL5YFZibXzEh82f+ziMgFCswuzIkBR4dP8mdIAk29VBsc2HUNFHDVKrGU
2aETHQrvxevQ2IKL/VH0Gk8UXU4tp2nMXGzUfSMvZ9w8ep2OMH1i4KcF3E1UwGm0
IXO2vSgsTSryccu5vmXd+rC1BqFE+zJPTrYnxbHLrmaqoxhOAIjS2aNsZjyJQB/h
0WsbfKwbOt9/6cCVbfalGIY/B8RWq2OtemiDIccnurUgIpV+HgCFlY0M8ulkHRzR
z8Te/bEYtQVHTRnglgax7gkw6OKXWbZuXnnPe74jPMLAX/XcRiyIEiJyr9NGHVDk
2irrYgbFHUeMRvUbVf3Mzb2Uo7O5Qaupf7VkYH8LEbotqQuGMvf4dyIwHLEGzW6b
IpakaYF4hhUegWu6cj6gCpoZs0SEDBgi2MrgSCm6wsJfaUXxYtmXC/T8h2J4S5HZ
QVAuOohsI72taMG9v8q/FFkWf49I5pM8iY3zXOKi83CQOq/Iy+2tJ53f7Bvm47Q4
4686N1/yrugKr6IXl0pMProUxfUsHHlZYc6jQ5/KepJVi7WLN773mOzSZD4H8AXM
qPAem9gkVi1i0bPcybinN+gJhzpk89lM5VuN1lDfJPJ+XRGh8G6ynbNmnPiX7KpQ
ddxpDaYhnrAldQe8+EMGXDtOUi6DHzA+Pg6nbN9gnAZCLDGsiDT4tGkiCZ4qakVt
Gkuxt+xWpuXhSwSUIMotZsm5ObNbyg1DlQSBl3EENSZVrr4uDKZEIUqz8xcyVQ70
Q6xga0BZeHbhgHkyFsRMK0rhjUwSSsk9BmLr51MweNSX4GOzxsm5W5nyP43y6Fjb
+ztxbMHcij5ewiemgnJ5I/Nr1MdLtPVgep5FYJeGJQwnbAdwFHpTUueT4RsrdQOu
ZC+pKSUKQH9fzH//RmJ/AVnvXpBL+P/Im9ITg/OY/dK4LlxG5ePvFqVA2iGP3Nod
qjUzP8WuJcFPmjll3pttrnRhWpKFQFoONxKCEJWfMtBE27EJY0MsLH1KhtSC4TGt
QG1WuusnRCTmCCte2eGbg5c/Q/YZlKyeq/RA5r594XNV00erzL2k+3BjhZQkX0im
us1oLwtjkGNLe1tOL7rflYK/d2bA/eGKUppMU0gAOyKFhAlpqa2lE1/RITfm9+kl
RnPG+HUhaPAvP2epH+SRUBXpr/0vTlgUTkp2oXcjjZUXvNhaTDc2ytIFhbVVb2C3
cNRL0w7SF92Udw2kVIsv33tP4U5vyiIsXOuZAl70j8DOXKK13wRhYbLZw4cwXqYm
R+N1nOnryNgSWvEZFY4vGK5PTNiBsjNvGEqph3TrneuPmphdm2HFvx4M3VU4Cp2i
a3Z+tHirsYuupaIKMQCpGBTzYhhWtpd7Ehjou/EWE/aVhFQRE1NbI+QQsoRArisi
2AET2U7OxQ0dK7zsu8yw48+l4XtolXllucakyIN20OPnS4p1Q0z7AoUI0A1+FP29
8rllX2TmR2J2nPeZZErMY1UmuBh1cVuFAPsI9DwGb/mjteiD2U1ngfqgG8acKngm
bjH+rfzFxjGdaOjzI9rYCMo2V/WU6Ra81SJGvqK0eUymm2TpzZ11INVBffWIZNpb
IHSKdi/HQEjWJhaedMYEmlG2P+Ntc2O8R4pOCT0/EsHn/0netIJlGfBeldeoD08M
ijjrxtsn2/k1xLoORZKCnerA30Q7unhrfkuDhL0sMZX/Eeeq7KyOcv6JQTPlA+u2
fUvdumzV0M/OpimLEkOuw3vvhvYCvsGsTx7bHH1+KxI0ULRDpzSe4k+tAvtisSaV
u6rNKoCWuPyaLyUw6NEJSdsl53Ue3wrOuewYm32HoIz4wxYDur0yZaVLyD2IbqD7
rb7rmD9v9mz+jeh+YPtt86F/7jTrm+/aYVnVQBXGm2ypbTVCs6B3K7+Hez39f9MU
3tJm4dlwmpPB84foBAAaAdz0DVip3HGHBKoIYvd4H3bgK6gjPw3POWcTqxIgDk/O
IgiI/OUAi49Qah1VApMX7zCjZayiKb84fG2JUiSvpWfBGnaA/cvFNR7iCWlc618m
PZG2lLiW73lI0kSLRJ+VFrBR07tSWxr9ZqVPfQfWOo6OZe+hKQeH87hFAt9VY1LD
iyypDCNTgOjn40L59Sdrc3q9cY3w6O0wl/XhcRoclaSrEcgEkMPfdZY/Ep2+bNB8
doQU5b3UU4ikM4upbl7BFy/l0kiGIlaxABG0j6fE3E7SbLiPeJc2MUg8vDy4mQ4+
HUYQMFII0y7gJ7mmo/FhHLxzzwL5Aq2qR94XK/LrrlpGDjCXfIYmTQgaA5P1uzwu
Yww3U+EZNggpktrF6UTYxlORta+N6dq6h4mmQO+U9btj5d6IeKo7ikBa4ncgc4nZ
+xkeVG57zhy33ohlZlDvH675BggKzBoYcJWy3dHOlCjrFcx5woOc2UZDd1tiM6th
cMgzO3L0OWjQ9jWQthv7M1+/GEFklLCxOzYVyWCo7zpHh2n36hGPQCedGSyhABaG
logQUfvLy92lEjLhafqYaHvICFvotGRMykbo7REXYf+3CiPN3Zf0ODdoc0Ar2yN9
Ay+RdtAp7JE6if/coUszKyQGL32i+YET/g+fQsC+FZD8ze7Qn3cW4xomkfs/RvNN
Gsm/wyfbpKiBF+NEJo7jfP0YnpuQQPIBRpcJamO4+f5f3yyOvQhpqhiI4X7ZUsXs
+jarGwat1A5TbuMQSsH+qOxDBoqc8UEfbIDOdh0PKbsqX3w+C0sXgin9Se3lInUy
PRYOgNKHGoy4NDZzps8A5aIPr69DfFofOGp0xTrldescBFaGKy1s5a8iANLRTzHr
szXgu+2V/+frLGT/56SaidWvMmYWWugrTxrtcGON8c0e9/pcQ7e1ymL+LOMepE1L
7X7nrHqp0rgUM0sGjSXrI5vcAha24/psqKKE5PEnN+bWdvDxef+wePJQpHUx7SDi
8+dMvfH25w6RsWytCkJsi990J6ictFZTxCJYaRFKzTh5j17Kr0fJwcELpkyfVGcT
6RS6hhejSoaqe+HRBDvYeMso9ij3Ht++Xmml8eqlon5vitJwnkd04tDHg4CRxowQ
7sPIUxMULg+GDbAVSobdnOA+8xDXgA38inlZjOxIQvffaWpcFbV6n7mWS22kFbQC
qx1jgfOlpzYp8jQ2v5m+pQgP/pEl7MQiP5luzq8yf39e+x6NZbCxFODIf7rdFKMi
Emry0Qc6xmthdA5PtisfoTbxwiOsrBpiau+VuhsfNmKsgCfkZQqjXirSAM5N1XVg
KShKdSapSXvj0sqQgJ7SFK0iew0lZLBFExdRbypFhiJD1m/TXMijQV7HXXPuY8jn
jqaZPsQJ4TxLQmEM557Zy935jb1Hc+V8M57hl8vdwIlyiM+4DRXL7pBeJ7iEg7+h
+dQSX98mgSguGQa43Di59Sz5fsEpgz5x5Fk5yWuD4v64blpvIWoPvV52rNtw2ocT
R0VGZOu7laP6B+2f9AZ/GRgEnoCUBAhhB5BkcOx89J/cdRKq1Bj13nvqljLE3HDp
7AamdqYnuOpRa25Y9lOoFglDsk9kMTh1DB1FBLNwRn6huBiwY8qcUIpD5gI1sDEa
v8+C8zizjkaBcNJji4JHla0W3IDfxlrxvAv/xyymkdnFJ8VgjKnD+eru+gAuHdUt
uZFV6iHMTTXZbo2NaSoEnwkPC1kZ+6yqtKEnGz/R2LQY8Dn37t256bEQvxEotk4F
AIyh1IqEuVGTxZI6oU3iZcNVJ6leckuyuk6EXePWDqjL7Qe6hzhUXqYainPsmvh8
o97Dn4JnTG+xHNn/VDpl2xIbvYwQLv8FJBCA24Q7YckR7qhqlC5t6uvJnTlm7RNh
cr2llzQixTYfJmUIq5kQJcWPy0+kun9/fJrR+GIE0+5gOf2f3k2+3BBoC5Vq+ybJ
+6buCby0ZDiMxoBEp+i7ksKBxzgZ6DqpLRChmZGQxZxRm/evVXnU8rsUca5WL+bD
2VgzC/dlis5X3mIbU1P+k9gN1DGrY4hkH4xkNW36t6WxMbGIr8YXiuPDXVKzkRdm
9oGMBkr3KQcVc16JnXZz8fi/vIzMNv/DeXPr57/ORkXq55ifEpVmzsSufFZyLsSz
mQfGnLYudpFHpd/KLLUOg38mLl61qK5qBQR0b91cd0V4G3dtaZyEcWcVCxLyUuAh
CEnMDTHY6ZNac2tHQIMLweY3n0iHzXGi/kBB/aHWxErdJqes4gnwxuXf8jUpnh7W
1MAz7Bi4VT+l99Y3O9XAL/6H03mUZuetntxkFs6VYTLnLfBdgX/oC+wNbrfBPB1u
HudzSTNU8DwJcbgWMC5Ngb7jBA2Cr+7cSWR7O62YLVBqI10AMC4viixKuBZq9b5R
E7ul8YTQI4Npm0QhvpCBERsqWzFylfvnmHeP0cq4Y+neDKmHN1dhsj+yb/bo5qsL
7qOi8KywaZrFc4S40yZCHLdmxuOjNj7ryhuIHCX0V8YoWHPXMXsYyAsUCxvjvEl2
5oRwadCo7O0whdVNxL3VvM8ApU9qywjoYXEQ31vbIqlp1FP1J1dyHp5Hg3h1YT/U
1Pri1IDb6RCW8LpG9NZX1/+YOCFolRSCS0sD308UfBmlmxs2po5DmOmKMohABriq
svezcOz/eVmieT4p8qeAmHyFCejmOxYsZiWtoIZLjXlhdQ1Q/GYGGmD4GN9Dfi22
x8+sW7gSFw8G3PcPHXsZI6aRH+55DCMNWq0Tio2s7IxZS6rvsapRZwG6XS8YRgBO
tktkzPK4ZWzjoLJ1Mb1/LGPxhG7j0EpjF7Audb/WIVDKAGhdaXt+1TsHARy+pmXo
I5eOWqdtxhgSIuchDkot6aJWl9L6S02BYZKx2j2a8jgS2BUTQWtfi9RNtOc2s83F
UzNVKyTQ0jfr8RUORWmBXpmN8UtIGembFSBZRslFuAHfLJTZSkCsYCROo9qg2Sgk
QbqPWTTDPFEA8e9ao5+KVcFICOIvquXfm217D8MnSX8gE84aFtR4kfFmJv5HtqD+
5InXdn6oTwUKqJnslQ2tGSEvNYHBJ8jZ4GZBHg6c7Txw7wnQZ+BkLwM2uVfe77lW
xHz2cniOmfUJr9D3UMpqmQ4UJwvzOUx/K9wfa6K0np6x9JL6CF4VP3thk5lY4/xf
HGgLP93Y77v2sBS1ydX4uUgokPqP8ZZlllYR1oHVacsL6ouGIFTdE88gqMbB0E03
KhlgDTPrEgPpG8KqZJHORMZEii6jcVg8wqjcAiMU80ScQP5Z6hzQ1pVVI3hzyCQ5
d4tlCwh6C0ADTx2gqWnVzGtD4lnf6R7E4p0Md3BxhRSjcbSqvMJh6cBjqgPdtQM1
rY2bFoi55XxFTRD9Oj6opIW8LVt/vFQ8k18lXoU6diLTylVqmZblS+SxnPxAXwnl
vfTi+j1nXlhAWEznZdZMi4sUXuPWvUCepS2QBbGBdaIb8smn7y8wdY3bBpBDpydA
OfCziAMUnOb/jpOCDoVTOS7CuoUtZ+eApcn9qrfEMc00HKFTkgoY4emGP8cJwryd
OLrI8kmRClyyBA6CqLzM8B/zysxbA+o/LkIhP5S34XAa6n8kSgJTRTLDBpDcm4Tf
QrIg4WRCO6qbV8zWZfMEFdE4sQSasKmb0i5kL2VVWk46C1NVWTPWW2K9zMiJuiLT
xnAhWjLoPabo+FPQzWSRP27RzM1VSFDo8SSWj1m5N8a3isiYtBi6nlqtC6Y9o/UT
o8+Dm6FiwOpC6WI+qqwllfL9ePDdCTh+9ofYNNN6l75wdgZ8Q+WN3j6emlE7nK/1
L6FGzEggXnoCaysgvcjRwzFR2zL0p8eg75bisWj1b/LB4ed7cNCGmNPuIX/KiKiJ
sd/Slf0vf5R47M9tJ4yqUx663bxnRgIuMfrXMYg1T4vCHHztcz7jEsLQ3rpnJIdV
MUN1TbzQ1JnQWYqhqxizxW+AWG/wlMmvhL9ZAusJGvpzEGoexjUpNB/aIvgZ9Yh7
pHkpiglmEPWef7vNf1bx0xOHZfcRscjqxkwafdI1jTkgMLpdnoefjPpXoG1TYyxV
2Vto0ccJALRg9Ivrb4ZNeQvTPqTucKKMOpZA3S54l0Tm/XEorD/YpQaLRMobsCeU
V+R2+PCQqiUduZavWaWxE2QsLhPBiMF4K+tq8/sHwZISsAHUjljuq31lnwnV4/65
ic9V7lvcrlezTT7tEWwpCQAgblEZRVB1j61FJO40CnUWRaQaeXZGAQnrjVRS74H1
79A18ZXQBwQBe/gQ9tY8alT4XhRikRLfZ20RMgTNAahPYM+1oIiO04C8Bg4fCERj
hd4vTlD251aXJyFFT5Zekp8bhe4UsCOxq+EbjugHYsDiP7LxOxrp3LqXrZQeUmoy
II9L/GALF0p1IV8Dtu1QZIJ454fHcQgE0zwTjTNvQmXZW+INCIVvUHumksJnlq+q
F6ciq0fXGJP0y9/QopFZsdQ+fpcNsJDOWSa1uK+t6FCt6plNfwz3o4J6nwBR4qnH
ZwuTsCO9w6prBerXvV5qQBHzZTfRlnb704J8WAtduUY8TIMr12oCdUpRXvC4hTL5
Z3NtW2IWvr76IRaqUkpwYcenNBxrq30i/D5K9VJ/hM+ux1uMb+QgBNdJCD1+KBSJ
S56EA8a5690Fdx+kgKPzXhgBlo0SPtvlCLw8RNZ6wNj3XeVcZ8RYgXh3Qe+Ld5Jw
JG3lnuJVOMkt5AFdYrPi+xywFJxgZrswICghIvX2oYGuOZC0FIiP0ez3zgCAmis0
y7jnDwWP4LbQhGV1V2aPrlrrafvc2ihwJJy0QfhZA21fwXiBxJ4UKtAwwkTfzxFB
fupV/4GfRKqcTweZ1jtUWrdYvfpmsNInDTWh+L7JbkDLgOV7Ew64FYefH3lJ0QFx
gzPwXWo9xm4zAnJP6ZU5PKAMC0Wusb37hQdM+nyuS5iUJq8z2gXHvnMl4gdYNN4X
40gRbXzmexgebg+uwAdbV08vDNd9V3W2wNq8pVtygDPnPyyTCPHKx75nG4qgxO1R
pfN+w8ja7cGMq9XfFy0mDbVrqz0l5ll3Bu0RfXTY4L9MN0WFZbGL3QdbaUoyudZG
ybLQZwyQr7K/ie6yZD/kdwdGIN9zk63bKEOG6dpTYbk9jFvVio0HCmuGj6JlKlW0
LQMPQXg7Dft3ao3bWvUT/WKr0bWFr777B0oSdWzqn1XQFLHwXITT201kWlwRzrOv
UB2CWC/cA2QXEo1WFdcZQRGaKAQs/DsiTadwrjy+YlVFs+mccgwroVtkakPGdHLV
SzUJXroKv/gfurXoNqZkmtrzMr5EsbaKrSmit4PX9oVyOi1/5O/WwCk7eAQ6S7/j
IU99ObTZ2HyrnPB+udKley1+yNuU0WmNlBypbsrTohkO8Iyz7NNIWd4331yI6gEs
BjIxSvsuek9GAVX3cRvMaj/qMM+6pP2nl4jWYeOfYn75AeHuW7nayCzPXG+erwDy
yWJeM9B2zshzB+oM0bYDaP+PLfuiTEr6U+mqqeRf4bNfFs/uZpO/qBAk7UtC3tSb
XaO3AVGRkKgGgujKouZYLNsFa4G9Tmgz8J55IVzqfLrn64xctvnQtGD7O7rkyPZ5
RzAZ6Jykk9T9RcXc7lqVcreYWyWMFJ6VjB54kyP+faoNk/2KLnhMSaeCch2st34D
EN8Yy+VyqmcG7III9pmdV3v58zQ60IXz/QjVEd39+o6bdsbo0CRRIr8r1xo0fKnd
HSLLrZtQY30hDQXStlUxwc3J3Fw+OwLyR5voJYi6xqoFCpDWrSMktuvjyBwlwC8d
WunexZZit1feXFboy7twEUrwzWmp/U24Tj3njmzXueICTVFm3ecpiCXmquvcvcJD
GazFdcpndwdRldVrzqhxJtbDFJwtOQVlXCr6316rsCHoDTBxWXO13qY6+/WuTMah
Hemo0r26Ei84miju9z9B/F8XrMEJSWs7SF+8EJF7OrF3LxYqoUPvb5yjOoMYgQu8
+G2AyJX+bZldG3hY0MZ1YfGoR7JkCKW6I0DNvDstMzA1vLy3IrHUT9YDaRkFeQV5
8bAv0REFf4Bix8VmciY8wX0JppFQhrGY8ds1Q0YAQGEWuqQF+cHrjC71MfZNY9CW
U7B4OIS08V7C9gJZhPruvT3c9ex8XxKxQMfMbP5rt0YFZ/HHUuuC4x/Sl6pqDMfI
Gc1q6dBopioineeDt4lfWfT6bGUw60W2tqa90PA8vyimb7jsSL6GGJ7HvgND4Zzf
CuBW2mROeJFgLT2ZP/nNipvPXwRIz/P7j2ZRhnn3rUu5uu8X8gqvPb2558jlDWib
Dir2f3QwHG/b9q6rSUnLURaRMNQCRFlQb3R/22ZjvLrU/yBHhjhIwglVWZzSodhf
/c9Yd63Ug4Hx2jQbGjeAFjMPFLDiGl6EzdVnl25AhmmbFropOzbq24Ko6RdhPQgT
R2fKLnrJNECSoV1KQmBrauBO+iY8gGt1KGDgAqctTleWZw2PyiLVfTR7Rw4pPHBv
durLjxvtrDeT7tgk+SdJug/eo+ncD+sSXkRBkCn/0v0/mvmVbL/hrNo3WWM5G8cU
PI7MzvoHPpV6yNhO775QEwErpZbnLXmMC2Qgv2KOimKtNHZ8zUn2npC0husipl+T
LkajlAlLzTTp2y6Q8ROddo1GwJK5PUKi2O6SqfPT3EyMkGqufVjBDeeEr+NHQvdm
DgsTQ8bzNzsgFODRMbkc0Vsnth1qxmKgErLBcDMcybQSAM7dlacTHlCCTukldU9W
dyOI6RbWWOZSY6LSbONtW0glsK8Fz6hAPyKQVj2KmNl9wXW3zvqiYOJpARL6kOFC
F4Ou8mHlTyCtxjYGFE3s4vDwBrVHa8gbUVpWos555zEffPyvjF6FThpuWz14HVVa
GpKNMZiAGlTioK+XcmD0p4Kh5MnSVQMDfvq+UclkkiY16FPRnTSO6ocF5iYzdLVH
SGhyLQQxxpipJ5snKicWvhV8Lrs97/eIN/D02T4wvGgbdnxCXzxDcm0XSg2off8I
BsW3GMdUOo+XxDTHgIDypA4NWagOfLH6HBUJLslV524bfMiyDDKyrqWbjlaaQXC+
Mh2N9zahGi9OKn0xJi6Vkt16pjPvTSSl+RC8F2MrrTEEO0p8FwED3GKM+HJSHwFs
6zcLwJmAyXKJsgq/vPZH3B7mEfaURvr678EG4l0PwVMMXNTw2o9na8CeHbj0P0fy
RG438VSx9bzcoDVuzLGEuO3oO/+yY2k+ZZzAHJHzZLfDcGcr+Z5Tn4rl3tAcCsRd
RYj2a2DthCDATSOqmV1E7VoWOAOpIREm/X9NMHzrxKFSWk+wHmZnIa7MVDhbc1Pw
fnkTMQC6Bs2+gTLvPkOSNjJ/8YdDnXEcwyMAWcE9YA+3HGZIrlWMJaob9z6kNdvV
e0wDas9LmyMYQRXe0OrFVo+sjEMxiOF/0efrO7GWIvr99l4pUc7/kaMvlUszIikb
7y53N+i5reuzZ5PoewcAb4Mh6UVN8SxeU9leJThCj5a/NtnHx7ZvdMZvy1lQhQAW
JhDZYY5pnzH3ElJCQ9Tt79Qs4AE0lNYCrcVRB0siwF1o6/7PlDKYIN1uy5zAwvnt
lKJDk+KGsPV64KGGgeXYivFA9vPklVjqUa8Z5AG/zleAVy+tdAkYwaBCxx+fTNRF
Tc/aMeFFj1lMRM47OGjD7Z7wjAR2VD2cB54+QOifN3zfERco9rdMtND0MpqSqZsV
PlTxKtUf0Wok/CZj2k9d1i54wfna3QLgiQRMZj6BSsCYHFbzpOK42a/lzWzUPU2g
3rcBPmiQgmFaUjj+ighUUkB18zz5vt8z4KaEWJTKzdJXfD//+aLyRehXPcmwOeSa
uuAic8LS0cc9QhBlH3yof98yDtvUXSAl+HPAjwwS4Zais5hdbkGliYbGzUiLW064
eFhLER68lKdpdzmUJQLHl27irpZp9JiebHT3KK6OhRSV89bcXOZPCHvR1jqL5Rnk
s3q+L9EloXKvr9lVKOixwTclFUbGGP6uI/ke+8EpWXMNX+kjxgM6JLKAPFSH8mZL
s0zeSlFA+p0r8MtVnnkuVPiGIbR+VfdquGOdMegYghJgjLsAR2bRZpJAOjIMiJXs
jUsp6mgHD3Br5YKm4TCey2Ch+yUAif/EZZ3ygE0UcIRw2IHOngKiockNoMcfF/7T
AMphorctp+VWsRm+uDJhG5eyk+O/cEKnFP3e28KIO+pLcb3OtovzzozaojQlhjKL
fRvXtsANbhvK3z7PkGds5AD1lsV1Sa8Var/OHG/eK/c+EpVu7qG8nL69nrK8Cm3A
p3Am5GO0tcBy8IUEzdzkSu8DdtD3TeMDa05/PJovVr2yXhKuYBiFuLH8E9aJAYOK
/Y5YRl7Gojzo5p1B44Qw98LODV/L6JWd5KzlqZpVnAMeyIX0YtWcW7AQ1WeOPOdD
5YxDrxWrKlqBHVcP4j46O4Sh436GQuXckCaW3VdJpVDukqoMGRDqWV6XehMgdpvj
aFRGfhITsyepONiGDAvCisBOVN/7L3r+NxK46WK4qSd3LqJCODCP4ZbVZBzDE+gD
7yXJOIW7t2GZxXlsUVhC1g0Uj8eypWbw3JBql9xbZzAsdlFpZzG4dFz/QoakDelk
8QzitdkScRgQE+cUhY47jijRHuX8vPiJ7zA7pTp5f4I0GDaDDsmt52Zv4ZX1j9ck
Uh+/GN3CYkusku28oydF65V8rO8eT4hV4Cc8zHqBlSzZ0V5t2dIcZh7HTRdgHS7+
7XgZ9duqF4GBZPI7NSJaRcOkMfUFxInrnb87Bmb/SvyaBgmVCTQ/4GdvOYbIFb3o
pAGjBxO7bvMwkrKhKM4j03LudVhszLGUchhMWs3LZAetCAHgiq0HQPPcRVZm0itq
S3Cdso63KrbC8u1YW3YXXgZES9zbTYd+E0R4RUBo7OldT1SOcEG8gc3sTNINvHk8
9D3Y1XxLL+NPlgzCcNqXvyVQiguqKRLnlDEqv4WbUY72SUObM0WHFl9wN/D08erq
bOLv9Lzv889aMbk8qvGgSx46XIMc55pbKobDec3Ix07wkjKPh7QTvKtXuGeJ94CI
uJDGGnmKCwfoiDa2VnVRW1K7ciCc6RAHhfRGIQg/d3xrXz3rbvQtGejSg2VrKNAD
NInTUP2IUUEOMpkfLh7XhFgP5RrPZcnGaVCRWtz8orRjvcEoB0UtmmzCSxPia56+
3ec31JTAvaGUTzPUZYbfXvPY9yNI7eVdZNtR5Q+K5yomi1vpTMXBXe0sHUyjitrr
YmRzcPv47hUg5NwJ+e+bJkX39gtxlNrj0pFLR06hPWxc9QcnUuK0T1D5Z539D9RN
SMVr+h/SMMOMDvld4InXqfoST7SEmywLIjtKyCWb8gXqqlTMrZdeufgIF6Hd7hWu
bCdSHDjOfrGcCSYpFuQ2yPWfmVImIzpNhDFfRlotMUfPbnjkdMeUNyeq0yavYbea
gEt+tIMmcPBv/myAvW17eJ48XKYOrt1Qd9N3vrEYx/ZnJIBUxK6eTNGEKboQ4zPL
Ljc0Ee1ThFDtrFjvI6083sAicejlmKJM+7uCvskgpsop8VB/x0nJJejOJd89HrH1
7GxN31Qo88W26Peqv5bjJb4ykBkNh7t1V2N6ldH09n/7fG3PdZNVpUQDiWM45BwG
DxfWHufycIlguZf4YGrvAPV9tukakoGw43aiFr9Bo77Z8x32AIY3XpWkQrpZH5kN
ToBMYZy3Z/Y4mKWKb1q5vjp3aeJUeiaR+ky2G1FbhszkYYYSNKYreP6hva3KUM6i
1WlumKTHK9KXvNQMdh1xEkC/zCBLbncnR2m3hjzZDTAA/Psbn0M9WkrOWLJC2IiS
lt5fw9pzlesu67cVRXrEJuGkKHRFZOpgpyQzYy/LkejOxbXAomLc5oR5cgd1HlXq
rFdAby69yPTlflw+yeyZaRMzskB2pJS2O7XEM45ZBhCM8mrYb9eclkxd4PzPmUUV
F1ByRupVJhl4I4swEc5hJWZrhhA7O8M2brPHEvRoLnS6rzmD6flaQyI0rGTHsGmZ
Oz+VA2VhAUGavZeNAwK1lo/GEAL247BwyG+IZrbAp3NLuR9xA9q6gjFpA2RTOxFn
SqX/gHprYzQ0pPnmKewviz3Sx6CaX+wYVnqalNorM86Sw3lTLjmkDEJwCrf54cpH
XaEt7p2WVJE2PucDzxkGw7rm3WGEA6XkaErvTXE2tJvEuofcdA+jwBQNGHLd487D
O7AvHGkx/V47jnCq9W6modZMCkZTteGyYyIAW3k1pi4bEcYV1GGkuGOExGwM7kdK
yHo/EExgf0mI3dpWlrIRQWgEf2L6UvQpv460it/AJe8n+0ooHyMq/wVmi+BU6k+7
bxNep3UNVeqUl6OODr3Uje0yErQwEfKMf5PRZUu5RCmIVKdh9qKzmDiPBHqAZaUf
fOheJKEOFVzIDy/7oNk6d+Lj/U84asLsIsKBP66juNPgJbcF+I4828ybTl2BtUxN
UZe/zUrAEloJS6b/fmXBnpPwq8CHdQhrCq3WxDbyYOf674oypCL+BgQSBtPYZN/L
UcvrEoF+O4b2e4ZQKTCGjnp+1ZQ/IlE6aGKVPAUJJAQL8BkOX9vBrut4XgggLxmx
vmM4XpBc62H28SjOTW0k5Ly1glnGTKpJKyk02afpFM0HMHo50z+/SHVu5skyu4iI
WxGOwM+EoeLIqsKGO88G/2kZ+VuvVD0Q+5uHXezmoKHeivxwWV2gHbbdJV82VOJt
XvYOz1535lMMaO2NVrk5KxvhJo000cf9zSW9psCYqMUVuDq0hVM4qZpVG6GEdHuK
SNJ/3+gUWRy+hydPG1amHk1MQwTpvaOPWelLpU7EzoUy7CdOw46/nIDpmf9FEX9c
Mi4mxDf5T/gj7TllDbWrdZEQAwz4inmUEHtusStvfcXfJ/Iy4M+cw4Xf12xHADrm
OktIB39gaGJmiXJTUcUbWWhBiBWpLG/w13cDdZT1aaeb5atTgVx1YyBKMWtqqv/Y
tbVcVQZZ7GfyB4Lg5kqSFdz2C+Q/omcX47HQrUMvHRnVEl+LtrAWLM4yFtdWMy7z
r9jrwJsTYndrdrQFn0D/Dk84VFoamFulZUcPLipcKNdN8JnmupuRe2VP+FkLk9aU
AzGdLTNnqJ22Kpkf0okt8fkyphXEWWLAsd7pnrjKWeSVWZJd0usGGyD1c9zEG935
2SgqvrwWtpid64JLIEZmFIQSYYMJt04m7KcNn26EaAubGWyVvpjtVE7f4omtdJRE
/dmvyW89OtMu/0D1dJPgvEn9xEKczYeLGVHtTGJFHlbwG7VFZGRrdMDYeH0ks5u1
OndQ9m9lgG5Kbs9nj4ElriYJr5zGVclFalnG3VHFIX4DoMRYFWhkgmfkzyr4m/nm
xJDNyukh14eFQInIg0OtIAqL/RzWiOls1eaMsUtkIvRPsIXF+cZXj2ZfB5NSmeLC
GVA1e6JLmw/rPvtzq+YZejwb9MyuhsS1k0cMKtWS05ocjeEictCtnp2iUry3IDcR
L1RDsdx1zzsORsipqJBbvyjiLVV/mm177edr1U6uxuAGFGBT6tex54B5bVJBTa3C
7DnpAVeIaGdfYIE9bL3kINmnSHPqLceAfVTMRQn9/0OEfSSXHEHQIsyRehxt0QJp
DduAbZWNlX3Hv5ciT/cxrvnKIwGm3lOT825PAO9gVrCHCGUOX5PeLQ7tFXrAyO2H
IR+CfRSjrZiOP566ghgWNWK3R9W9jzfIqrTE/wUq3CmrNBexjikKeEo2vcSB/yKE
r7frNI7gIvW6f2ldU0TaBQJHEwUP9Mb0Bq/QyOu2dEXMFobkjC6PAdc66Kea88hX
VRR3KpkpdmMIi78Vp5p3UKs6BjPUOulnGYvBjhtjDAZ1ATyl1yiNj1jdxiNCF4pe
aBBL3+SpKHGVJpSkU7ql1kUQnv3mbJynhi//IvWTLPnn/R3UzQPdn9/tzPKjNLb4
XRMoWPFI3raR2JQlDX0ZLgNixo81F+FejxvPoRgRHGhwLX8HiLswrSGizQCbDlG8
ybzyA+ZfVIulxjLiFosPgM762DlAZRaK/g3ODPnvvgd65mEbRbT5kuVqdVvGgKYQ
6Dl3jwFU4x6NHM0LFwnYBI6h8EWeLcF7MvPo9QIrBkx7SSWL4gRIHVIgMFgd1xty
r070YhHulNGNLnBhKHSeZadFWZ0G28zIu6J1rHl3HyEmO3/7bOqX0YS6iI//qZOz
tQu9U0MsGghPdPw1jEq0JD5EYSNdcV8EQMitcNq1isDpmSEMZyXQ2EWpOn5yseSF
KSDU/qMNxW9wKD3Cg7A5wiqUVfU1RzDcaOBsSyV+qVs8Vwrn+nJydEbiZBcRZ8AJ
8B/+vd4hFcLXrqNOAMlL0bGbNH9sMLIhLvWEx25ud72zkpf6khqv4SAJ4+tX93GU
/zbepQpeRaGKz3OieAIxguHoJwZCuISYMcFQwpmRfwHJHaXuzx25VEAmxKQoyZvZ
kAwB2fqIaylPjai9D9pxbw7PpJCSAfylmDz3xn7GO2sOvE6TdYglLVZ08Xnf2A5X
dex8/gSI3TqPRycoSH7B3E4ieJ5fIEqRze7Yj5l/tLhaA/JlwgarIA+5he5UE/3Y
NvezOqfYTDZcCJtktwauyWA2F1KdqSJEsqtw098eh0I/sTtEBKrkj4i5IK5O0Rrv
ffrKPgyU8RhRfRaYfNOPHi8kml7kg+x1Vg5LG1WosLCd20t6lKcklo7nrg8am3MJ
p0AekRv0MzEKgDqU3lMlcvlfZdK0Exqe5PV2oCmTRtK4mU4RNNypXELjanYzrtoy
t9S0qUgKyLCzT3ON77RBur3GceuQyZl7YvLcmxTzm4yTdSq/u8+vWzHfWqORTHQs
jf91A/W0483TMe/6sijw/rPFd52X1SR3wMf+TblYlgIWRqE25ds75g3uw4hMdk5X
ah2LMPkU3qvYJooFx9uQ7+LpgLDGYkCiLRyh34WiOOJAyJ5FFXCIt6O0KqDOfjHZ
hRCecIc7WDj7aFLP+47Yktz3n7oJPXhOZicqF86RcIusDcxhF5ybnGP3N2aDFc8m
CUt+J3YfXoeVEEGq3koj6Jy0yoMTKpX9d/xNeFZL+W18PFwZOnB/OFwDj7Xetic7
Fn7fG1iZY0vDmOVRVlG4//3nfOVH7WVWKbXxnNBR8t/0/NcQoIOslen9JGQOPWtP
yl7FU4AWBrhTQC6OPowxAe0j2CoDdonYDXa0a7komL8czYnLTj7XkP0zH6l7eB8W
kveCQBlh5lWpK75UqnMZ8R2zuDhHbx4j3PUxjVNEbUcUQo31kXZ3hf3v4Eb9Ymdh
x4DNMmFo8BbDHNyBEV1acDg8dFMJ+2e2LMOL6djD7DyRaEm9pg24NJ0+dxrPn0gj
6b2hIGkMQVBdkeXnTs7oP08LHj6Bd68bCQ/PGQTxW2KQz7ezRMlhLUQtYBjtKRXq
zpTfSQ+qV+rz5pdgX8mcuKaOQ6iTo7sTb7CHiPypHXRgkE4ECcuxYwxa6c5fTyq4
R77hnqgHvY4s4F2sW+elIlH4NNygtXp9OF0VERTaUdTVTQUw1/np+JgprNJfJfxj
Wr+SBYpBlHPwb8FWlCt5UNQT0xillLObH5QwbQh8QNonHnEoBjDOVKRuSBX3WV0P
Kh7ifeGOoizMY/69d/4le5GpgAm4nN4AJv5ZQs2yfznyTKouoYH5njGs/UmyDQfy
LhtMdDxwpbEOJoq0o27J0Ihtn2SdqftVc9h68IHj21JpqgACwUQnV7cJao6McuoX
AaxZPc0kUvdNPO5vfEj1m7jQf/u0rHUaXZv5+hVYCHRllz9rSyxgeAtgSzMjwlzf
RU4N4ssZcmiJvtausZxzenDiERXBYzPB+jWhTzttei27H/9qSFGa7CYCNuNTEf8K
zuGfDNZxmDKtQFoUQoWb1+a5oHnQCW/IHcI6rJh3Ylwove9zwUV0aDxe0l+s6TLy
sXkvLky343fL41+KOwjRkbr/4c5qg4BL7vNPvwPy8jMe2IxrosyiTOC8MXT65iys
iCwZ7NCRyH2ezaf/XI0m1sCLeYC85NVFW3c4fV/Ib1kHrkAAwlODHkdSGsBtDPCb
86Mxa/owXo44WHfIYxOZuA4gVKJXzNRrbZJnV9Bjl6E0vgBdkdXAn6LKpbMypxw2
fS3rmVuDqHno+TNTe5oXvC5lfa5yzsjc7YNkFGuzyUaILSh1u/YbefzWPpWRUfKO
s4jw37HPb5n0+P8KmU4T4tQ6Ynz8OCUBybURWedpRPoDpmge6j50A/PrHI1fGg0u
8gs8XfKPYwBn/1w2Q4Bjgp8v1+5/F0uwfNZfQq7aXBoKDY+zCoYdf/PN4Q6XKUgD
F/54k1yp6Q0bJh2x3ZGsOOuMCgCR5vRoWcObyxR6RK5WrhakIMuzuF8s/SvUa1NV
DgxW9Ff2M0EJxrVMJ5f32Uaysgg380o+F6xFolWMBK1twkXGNUH2jO17GNbDpzyi
ygT057qwRCDvnKCgG2sY5J1HQxflpGvyFhAxijFCuKF4hdBasiT7rHK0dxmpqGzV
G9m1jOG8oCnWv7nAzmShoEHu670RmrcvNY5nSpccn2gAbYZ0rp2OVA29HYXW2jyf
DkQe75ZJ2NBuwiSH3IjV/210a2DbNv2ro3iTGQlUB5mbGxkoDTZIENvEFAp4kIsG
9aI/bEF+OLC/ZeTnJtCZgzhOiDlYNKs0l+4qJseVOBCSyJBKsRsxtL32H0HmDOzK
TFny8IszbmEN+HE5j9E55QICN0RalEpHdIpEoRhsQOh9fwQAVCwTtRZLb+pEb1pD
LZ/48I5c53Zv3HEYgo7o/pnXqaZIpoKvshEIMpEdu4v5Qd8oYtaOmKntHdRd7m43
dPNzJKiLqwLErOGAVJ3vQOHWvvZ6pXLAPEnmtHJkOxJmAhhL67xARolZE/d90P9A
Z34GWOQOCagyEQGV7J0kRHsvhhkQQXqXI5s8SS/8Amm1XXOO4SbRdJ9LQSalPoAu
y375efu5shWrlP8YLAFhQxxffoiyc6Qi3x8CfwdoUGsIykY/6wqQ1oYm+Zt/xhPv
eaoAjOGXQs8BezFGCPvYd+MXDAvFT0EPU80ApYgF1y+sUXsrPphENqtxn3zsumFR
pIE+GNRmn9+OrGVZ7RFKa4NqnGvFhHRTx3RuA6gtsq3ksEtEN2pscQBHLKR6B80H
PCi99OCPUV7ESnvPHLWWuCcRN2GabigPCm9YDIASATBuUXbUQjprqNeb1QVVHtNa
SjNf71mmkZlBevQhgLXLGjfyuvm2Kjp9tIwqSvE3/1Y6kOmfwKVYheeaFyWXUWjX
GpRjcZBHHQNib+chB15GW4z8rZJO55faoHx7uD8jlXMnNSoVTHciholRa53fkQeP
L7xAH1Oh8kPdl0LjK5h3G9YPAjbdE41zyW8FIPjdp4XhMoj71kUrwsq8lDKU98ma
7MrsreoVmtxJn433ukT8sDG7Gs40q3Ed1XUeC0ZKod3rQaGMgCEjnswPk2wVMTFo
nDDkKQAhwxxY8Dgrazcf/nEcsBxgwcso4sNqaHQJbDH7yq6c6RXXZVNOCrmH9gnA
/yhbord/dgM08gkLO0tLsJEFojI5gvunP/zpmljRZDZa7EaTsppG0vk6/OZFKbFx
UuyD1VOSjsiSiH2XKmqTADG+9DCZzbeuYj/UvBTkjvP8+w/208G5svNkuE7zDCLG
Rvi00F7BfWL58bF6Z6WYX1a9XZXRnJwBc5W/xI7V3N03ab6ziJY8piVyu0xpmJDS
ucvWKgCewXalpKN7gPTz99tU4zzp6Y3KcHJTibRJuMzOrmvXbCrkyzpLTCbzy6Oz
t5gW/bSxT24gZKOxaDi9GSlJpo68gC9RtUkv3gO+iJqwRD+XNxYxOByv2qqSt5+J
1VneBVeytw5icU1IURNcRfYR6ZIE5AX3biXMSVdk8Wu04jpYdkK/l7Af76KdufUP
2UErbENo7G/MeQmJ6cpQ5QS+OaQncImnw3/2QJO98ar52NkPz9I5YY52jXbDUTnB
11m4sNMS7t0DPrONJtQ3OF7NzkzjC0faA3bCu+9+dnoPd9pLgOK6vzpOIsUcH7kx
3jYq5JxKtzUkWBUd6Puv3nw4I8aI6Zgild1ALTPYh+URPJ/OR/Nsff3oEHabNMWE
RdwVbzylQC9f462Kjn53yDWgG7DSWlSN/WyeY+G0oCj2zxG9u017Br2UC6HpuIuY
6DjQHC/Uf/hpx/P/ZMOZi1eWaWGWLNzR4DE7MBilN56wVGGQWWXYSKyUahGOoLUC
A0hwr55spr/OMkWHZw9aDyTY6mvrvgwSCUMxsqQny/KPR4YNtppaYblu0Ga7ICcQ
pNHvwZ3GgklS1J1ZnyVqXLAvVe0qEzktd5JGi20hSZR6xWCbRlKxTR8MgASbKCp4
u2aROTwTIiC/usjUrFClT288s4D7WJpL7z56+QZBwk/pcgn7w1FU5/mc8racB/R2
imVPI+22znmzeS27LvyQxxUoqcVhg/Jk1sAfrX2gwg1ogxZ23AVOh9Gbu5Q136Gr
PmMgyH2xMfNkzydlOxflnhc78KH01/6F5affnLoCyTvnXBNw/u7MSb1lSYhW0lRH
r31LHG9IldwuO47jAr17HKltE/99Ck2UNKYdtB47rth31dJjJYqQ5nVQGpBhM0Ed
T31B8Rts59BUXnC5ElkNESWYAOb7r98axan+H1XbTOIuhSDUXd2I56EBB6kqGE8u
t67d8/UGI6/IqVMxoRd5jLF37n6tAT2xqE4w+oi0nqu2O3bVH1xNvBeuOnV+FPSl
5qxKnciKUTX18JtwGzD/NyWeNrNybLSsWozwnzt5OTIqI6KouAIAt04mnbn2efLq
a46nlf4oTTzQWe8xzrVpwMBJhfxR9HAZ4gHwy9UF/7n3W5vodeTLt3AY8pIGfbG/
CSW8ICYqZP/IVCZCsaz8mcX6JG/BGKpuXzc1+aHRvxhRyFcqIyXOSG+Rm9FI5AIN
A4tURQkr10+leG138opCh2OxwOPRMsp79GV7huhhgfUdLMAYU9LpTIir9aH4dhno
EoVwAqWOsTDHTcnHlrkyg8KWW5KGawotqof7b8iW2vllD3Q6BXmdiSpmaMcgHg3q
yTzb+Ph33yiZ4qjxpRSsVbkQuevhLol5r4o11heGMff3fvehD/Co/HbnDL7TO1gX
GppJMrffKG+oVBUEhyspNjcLq/nPWFwE2OoWkOKHAC9me3z2rYq1AZmTG2UAP+n7
X+oJdqiL8BTivsRBB1Lmpr+Nb0KXvT5m9oespMfEHf7dKumpgB3S+0CcBYYCOWda
BcFMm1kNvCBEMUfkQjCEgQXx9fNCMMih4lcBLe5e5a6LNalkm4s33GpzEvAnVjIA
RLqIHVwyQj88I0IOfwx/jWpOX7XT1Z4JCYeBHdXrJFOorP8k7PTGg/dyvROiRxqa
mu/J6A1RZoAg+1yK6MLpI4j2AEcs3m2NIO/OlSR8fZDU0WiB6aXMWjnLKlEqvLgc
EbXyqeXkbSt327YYTvrqABb3VvJeLpx66xkwUEe2WFtD8LYYSwMuSqPi8jFeMtgJ
eXI+v5L2pxzaR4PIFqxYXzE9V+qTh/Z1B62SczMJsgXoO0zpFvQmzfTIvKxHs3Aa
hbjc9OCc5P2J8vSToWfDskJ+tgqUSRbuh013sVxEtsCCXuKpWXS25te0BGcQl2F6
XXnMoNPJCj+iy439lz53g2OalymyHvvyvup2f9B1ISywnQSsKJt9YqfZtOrYvchD
lGu4kp4Dm4maF+er2f853oid0Ucsa6rJGmnUghYW8FHBda824BTt4J0RS77iCCV4
u5QkYIy1w7uqlVow1B50n8oDcQvzU3KBhv00KmKoTvkYbhGHUZAoBVcY17dm+TRA
URFinRKd1LaOfwjtIjqHDY3V5KnoTqgg0aUJKZ88u/VIJ9L7+w23rGBqzAk9cl5W
tpLPK717bWZBCVl/PIfsux9euO80Zz5NXhy7Z/fY607ry3LvcviTmOZce0rAagD0
a3pM+i7BsOjxSNcV4CqBQmxkoAU3jX2KuQKCpQ0WFrOPnfa2F79BIJ5CoCHHz7rW
Qd/zSPTlpK2Zs/BL5uLnPtudob0hgyYpWpwgVLwCqI8aqO1QnA3P7BZXQvg3Xdu8
Au6fxCoOuB+foJR8fwSHQRRIHJ5etnCupvGTdCgYsSt4jlvv2Eo3q9GqTQ7cGEsQ
IiLEuxopWqxEFijOjsB8/LzExx4EmWgipDGC2Fl4ob5aEUqw1awsLnMSojf/vr7f
GPT0qA09o+oGZr8DqiLAdxCHPwbK7BVhtIviKlErCcNHzvQX27Xz2fGG2I1MdVhM
lrMicHXdLfE8QHE1qoxkwKIUHuTnAXqO7Zxd4BD+W9XfOXS1sZrSk8RcnFM6e7eZ
tXQdH9ocmACUhoO3q3EDhMpu8/zn/cLZyOEvYoqIsb36IjrOeaVnj36LmpNTqCGk
itN6KWau9SajmKhlyl9sx9NCnP+JHYRK33DINuo33sAm4pEh6kaD4TknPC9x4kAy
c+Zr6b9jkiseVyQkccecBTFYau2xsLtTFFDBtQuSb95NLBBuFd8Ti+OcfMq12oM4
2mLerIBc9/p8aUwSMxxyK/lF+D1xEEcpJHGfDdgwHKSVMDUYeBAlXG79s2XAei4O
ErPXrkfUwExHIkPBh9O3YYcqdEu8nr8LgeA9Jzr0Xso1iPxJe127R57M7jbBdxo1
diJ1eiFsaRb5bFcaAi00pkCABBYszd1KOrjAyZkluyeDFL98NKTwTkLUJJ6C3Edl
fZxcA4lcX3SRDe37q7Lmc0DRzNNDLX5tLu8hLwaxcNrPmSxqdpL+6QtbWlUnyVzj
e4dIj/bRa4AiuaQQgIYJGE1BED5b3CNpYBuK3+DYliRUvVuWISRX94Q2t8ye+Vrs
8mwJWZGEhkErQGh904eQk4KNjfzqx6v9PqDY4iF06nsVDefo94h0lXqPQtj8wuo1
AYX0OAyTUVTB0mstU2V6sh6kR3Kq6fPr58nCPdPkUtY5NTl1Bc6hDJz9ObXayHwS
codHi1pxgsCqJXz5aW4184HfOjFsWtvB3D3d/3k9Fqj6oBqYN1AXnwTm1aE3Ve9K
hBNtAHfuOK7D7apA7PtVAHo/6fRw2Zm2pu943Utyh8XTuY8Y8WQ2AYNwDN2hX1SU
2jTBtbeQfKSkI/z5jCskhIOBwQkMCKWmf36pvWKNnBOMujix4PKUFg8DDQKhpwIt
p7PiuEdPudZ9AQ+skmjXhdmbb8Q4WhpQxBg45O7Bzx1HmxiS99MtjvajdV22oSy5
jOx2hg0agnMJpH3hLDXgw18LEiTg3bMA3Vbz0VhK+rghLcbmJc4AJd3drenEcLUF
jzgh2WVGBXLtHKV3g60BqSYPkuP1lfeW1wDJ1VdUU4UwXMd/I/qM3dp7RLKxSekv
f5aQExuLy4h0gdVDqI2RPbC/pTAl75KIJoUcXjArCWx9FRxUJ2fgc0OgmShz7EsW
ywifnFyuq/n3X5zEA6LKsRqkuWC//zLSyl0Ryu5EZ/S05pe5T/9gKwOldsjtdkWm
e84aQTB8K/vNJtAYDGOavFDlnh6NZU/w4A4kF5+mkXgwenO/pGjdAq6MUlXuUMaG
xbInhHMQv/ZkdQC0ZPAWLJfAxYlGkB66FM4mj2Hnr8YtqUkj/z6QJ3KkkxB03ZOL
NoO1kTx/0CnxOOOw3++yXn1y3rr3P/gsZW4n4lIzNUXwAwDrqtK+syl8NK56HER0
07S4VZ1e6f0+KfYD88XUy0CJ5GDlnIn0EqXCIYMILJwjXPXnyXUYvkBDOIl5OB+D
1pgd3V1rGLXBrgOK5JXutZNHgXotPrr1ujbWcZvYkDi0+WIX6WZTmNuUqDsEiEdk
z814kScu8/oqc5T6f6Qk/842m6qY4ME9KfWE9wpWCnbAuODzf5tjPKJltxbwtbxI
HpobZpUPDgNEtWVhX3VR7dXeIJP64O4yLT1+xsrXoyfCVSC13krsgvOc9kYOe/dY
BSc2ED8vu22D+WKzwSA3PqYySvik+fn8kgjZU61vOm6tVU437viOY9IsdwJUzLig
K4HYYOKP+56Ken0jUipRpuShXTeHMxDD9OiTDXa4Da9Bs7fiYR1IsYoRbLCZJkQD
Q75gYe3IPqkJtitdNhCnXxhF4Xke0SJR+TDclNRa8Z8wuJAbUHXuvAwsllxd3UEt
cg2ljWtbjSN3Px2EQqMrVADgquWEUlGL3IT3dZq9IzjJyGv3hNeUpFXFdLTiwkzX
blv369pjd3PjifU20oJS4Xuy80bASBT9wDrdCA4OuL48RGllLxY2jRfoj90mUxWi
l2G/7xhyGOkL+/v8WORED7NCboHR/gPCTVIa9lTsyANHh8TpmcAq3Kym33t+8Uo/
4RUXVNGQvRQdXQidaf/dlZMoWDFMyNzAKhn/cAEJWPyuUgsa0h8+a8FlGzkS0ve/
++TsbphSjbRLuoVae5HuIt7iA8oIvV9QQqlChIdknSJxZmfcGatsA/J8QgJyHGIO
G8QkKTmmVRBcJTw9CT1YOMbUeHJ/t4NUlkzSM9mcaox1w0sRKezD5XlKQV0Xv75H
6G3U8WMZCLVLMtdItOFYCCd0CSE2389yiA4vLXazhu4HFiUkMql+0JhdCPxRDatB
BmFAniXgYHVUW0B4uLzcIjqy0XdFOP0yRW/3fVfKYl9dm8BMbwpBlm1ixEmZme44
1Bmj/6Zqw6V6/yyO7+03CHIz7rcn6EFOZV50VQTCxSbjsexpMVKN3yzJc9v4waVo
Iu5bWWMlVKE2upzclw+WJMKf+XwHAO9xgXo/9MDwWu1fcm7rCS/z3Cs/jIBbRXrz
bOj8GjWGfsHfHNMc4hV85OSinKU7eT9LYvDn+uEBGotSn+rLdWQkqUj+YNRyzMmM
xNLHs51p8X79IgM14WZAdJEvV0xgvC9Z78hdWwQP2o87kbHmYDk/qRwgKMh10V23
FgQQ/5lbwOzYSgIPi0RThqpp92YQfIBw3yjz0RSC7Qvlt95G5datK3j5D3orj/0m
TGxOkq6KTMrp539JmWK1VODRNTiHvu65tJOPMf3jVc7WZHd1rg8z+G59V//PbR5Q
wiB5pFvEuzLEI97pNhr8IFKmOH/+XyYTlwhvNWtMWpxC+e4qjGY4QViQIH++S9gD
i+yAhvwL/VoXCDY20DTThEg4t6qNGT+rKFxcah491K9w0Lgj0W30oFT5a+CcgNGh
tTtn7iBrDr3yygOBaxawI8/DSoflW5xCE8axoXkTQuN+o0EdLeIqr0XYFwRuQOqf
iD4VrQ+Tp71WdwsqoCULe0paD+/pZpK6UuVU65+Lu4HjhYhr0FI5KjNBRL9I8WW+
FAxvrwGCTlmYE3HTRrn/VjHKAwvP9MXdIG97mk6qvXwBUs4ae2cMolF//Lsnzbl6
6qWrWzJFTbyZMDeMwVvPvqh+CCojp7I/oBffDq5anu0VYefumMdDaTMqV7swc/5W
7JqcK2q0bbRfLYdohC+58VI7bO89Thxf6B000Ptv+Y4CAuvFggf4lnYasiGOmKJg
K+XEY8tztpSdhhPa0oT0QFrED9ykzqx26UoIbpX7h32CwzrROGxtGJcvVMzowzq+
4YtQC07fGyEItLBUzaV2qS5Uf18O578LbQEoguYPdqRk7utjDlT7mYxCgHuhFlvR
J5adzE/nG6CxwS81ro98gYNQnkfcrkc0ZLkbd89swzWPpUb2xf7sGXRemqYLChz5
5gSP1i8EWUe03g7tTVcXpAmbdCJDzS5Nne1QWTV0OatvAU7fdCubITwij6CeTylP
ofjjM/GnsZMwgJ+LrruovUzJQ6SOf1SF10A8qvoHve/Quf5Hz2RKI86EE0iyDf/V
4OrdHnVbxE7Q39XgubUwigDjXxgb3yX9xIqZ0u3/tIe++rXU5g8CnJTuDYTHeWiT
N29fxlhn1u1InnffrSq1v5tZ3b8tDqR90vc2J84Y35ndWdS+vir9JSkc48/GCn3I
UDdNsoVEe6A9YG0Onjd8fW6UFIdcCVqgyxATzK+OsEo+oja+JDQcei4A1P2OTI7M
8UBoQw/DMUFGYg0ALzftYF6yBAssvKSZoyO3qPygPHRlALNq45RGZtN82VZsRWH6
z0muu/3xRQC/8eQI0f0hCeb+j/ucDjm3eRmz5FVVNVozVL96QwagER9ud7a+uiT7
pA23BcQXYkEA7x/LL6U6hiPXBkkdG6T/rsEqI/XjIo04PFo331DM3zRmRtKI9EgM
6HvSIhzwpEfsMAzGzoWH1Lc93EeT/xYp2VTg/k3oYy0HeT5iUvKJw8eIekB2UID0
Yh/jenNV3i1xBn30/Y6uuFT+5s1pILWVYjx/EtmejvIEvIH3CYw9dmFgm8riPIGX
VvnjkCiaHU/vm2oQ736BmtOqjJd86fdQwmPa4pbWZcWKPh7skYuzkQon2VVLQJDA
hnKLpgcoMnDwe8uOvAtpETQ6SPf8PT30PpU/8KQsk7eyeFwVl/0ZE3iNDifLp1w2
Ztf5SqkzFdnuHSHomzMSeAtqcLuX5hNnFVgDvU3wXlajyAnBdKa0EXUvFN/9DXSr
WFo3eJxId/o7SlQGZ7p3WttD14G05NqJIzhztibCK6LviRY4HcXsAHPEHLx6qxa+
z5utWWo53XpO3IhBKskt0TT3rJIj7W4ijCIPvhkOLIAgE2aRJFM9zEw63tLNndMu
CHAd51k160ZXtyenEHqMyLcrEGRCXkQLnd13mgzOubN45qQWJVu3/NB4dNjhBm3S
Nrd854uRPRksn/MG65BgRalxu7gYzIDu/TofPTFizilzgkAEupo75dZitr+VBcqT
A8E9l94kjFR6UN+GY2TIc9ZfyT0nHgDsuXfb6TdohieQ1tik/FkMM5t9PZY1HWnl
Ob1oNpFvhfitXOkEvGYvk7PjEorV4Sz5+VE8cDluW+TQNkiHFI2TJ95cq8gD913Q
MSvGc9xLoJIgmeYJ1bjixWKgd6I+L4/aggS24wka99IWZG3a6N6nCRrjM5d4gB5c
FdbZGddm4KWUeO1h5qljNAX1oIMSY9DrpKYfDj+Chiv7Ym6FXQ7qXWXTFpGiNc3l
kR2iJahsY999WDSLwiOJbUCKs8xQNAH/FBuGa4HV9Db/E8f6IxPV83HYGEqRr6mL
xT5IacD7qm9ztavmM80P39GUzE5g59+urV02kkUJZ7LKiBZsg8JEVLkdgEaC4Ell
4mgc7KySrQsCZYWDnazKot+NYYpxvR2tU92FS7RQuknv6KIBTzSR1Xz20XIQc9i+
cLtvxMBQkWyIrZFY0ZE4sYw1ZIgHHhtnQzglX8g/MV99dt+frYENdImnEXLoSGda
5/uPCQNh9fwzLdJ+OOoOgG6mEAgTVBQWR0hdtmw6ertohn02r9GxbMWZPtQ86gDJ
iWorliPWiENAcwcipIEa1GtuIPGVFMqb4NA19W3gE5grlkJ0zkLYm6UzMucoknzH
Ez0lHT4Dk4mbN7IVYqq0QetjuSu19nsbnkQmEQwmf3sAve1SpOfXVp1RlW6Q0R62
qnLmfF6Vnfs+dYN0c6PGedMb2gz4vpVwl5bYYIQnr4m84pWx+mAIA2D+KilhJZZ0
TxTU5P3aU1TkkfpUAuZiMpRB88IHFCRYuG0UDFjnqeq1DeG0qDtyLr4QCD5HCKG+
bVpG8XmJXlhV5QJirU+y1dtQdxI9roTSEOa6yJpSf/G70gs8ukInxi7oCDs3Xv6Z
8A/oDwKrPuifTWflzcoj8LS2VtxPLx/js9M0eWEOVhZS0iIejytIwqB3NkefQmWu
nxUfKVC0zR18y/MmwX39hNSr8Zb4K4X7FFLNCP8mvgVEBFLdhJiEstdfTGZSZDQt
XIRbdo+pojLGtr4tjlugrrDO+eFCiXp9D5OWypxH9aVmK+QyQMKmSZqN896o+3t+
XRu28+9COfHtTjvi07XbHR2fdnNX1SueHe18ZsZzkWZcThLueOuEhYrFSv4BgcUO
4D92LAM24cLAZzQRoxJLjpDXQYXkSZMuM42bJeZHCHZGGDDalx6Pg40srsy3/O6U
yop9TpSpSZoRf/mFVv08oiTZWQMAFK0eHolOiqzL4Wd6Viivm/QwO2m5AyjG9WQE
RozKZgmXxGht0Cr2s3SmqJt63YJR3bfbAfVzIVfhERbJKnc+VxE4NJ2XCGy/Yr7C
Ajd60djdQCxD3IGaKWjQ1Png7b9OiAvFUl+wCB1UjugvirDbVfaLMCfogvo8pYRt
a/LppRTDIYW3jjwFWWaV7I6u78R1u1QZ/g5uG3nHN4IGxNjpvB5blOYDnbNPQ2+G
CoPgKUj517htdiZtbxySHLjgqcLnbd4BQ2Aqa4+z6v2JMBGTOjBf+RZnjiSDa+XE
AXArpXHwlSCTcqXRa5z0hmgh/UZCNsnz8Am4SimeOxmylW9d97Hkek/dlHrnDQx7
B6mE3Uy3I3umnwC6kEvqjimpSsDEc7fMIgTFIN94lonqieKzVg1F+rzcAFbkNSU4
Tbdrf5G5Imj9J1b/dwQXTG9+Zg0IBemsp3xOBFF/de4LV/uk+s7nKPXmD9PhQV+i
Tbo0LGgCqDUx1acwH8/TdCwMdDEEUTo46WgtJOESI5M6aY2Zsp7puNxGF1bipGkA
MDk2JoTRUrKlIGI/c/OiEuRezyZy/I2fcX/pfIQgep9fDxNVTNV6T/RVAq/o90I9
VvAWDr2cBbuhmstgtxBw7+N0Rnrdny/46y81yrXCMzrSSm1HkI958rxW50F9Wdd9
/jVEarlxCRrBTJDV+XcCPGO9PvRXOhFt3svXfqTsVFcbnjsNKZfA+TEOlCgJ7rKT
pdGD4lZhmR9FPahfmGfAN5Eapk25c4sw61pbCfq+ZJgm0OS2mw2XWjGZE03vONVW
kESVS4zC1fSODbVPeiYSl8L0Cf4WO0rBlQxWzO8/6aeEf1L9Ds5JOVm/7gaxlj0c
SDdx+cFb1TQfcLO2eIYEPiDoelnmivov7Z0n20xsdq1cZG87ln1AFRh7lI2NujnC
mLHpMdbsUikwUw8r0siI4G3uRVnYg8EZVMsfGDbpZNsl+mVBSTuwoCxSNjV+1JOf
1AB+iD56kKIaKC1PAP0SodyfNGdVeFFmuD/CAY/nfZRe3qs1Dcf4t3HCT3jyu+Bk
Yr8m0a9/RB8wDsGR7E5VLCR7CMAmqkHtmLg9/tt76ECXjYxcIiujGfjC+NER4CWe
hFxQyUwlXYkiNAjKCU7A/Q21ZrB0cgJRmM85KgfNJe2Obi+lfSC2MlR0ieV/UwXy
huu6TZyrC/A5JLOr7vHFyz4DH72phs1ImAiEH+RKaZ6zkWf5yv1XE5m1ZWTTldO1
g5miiLQK1ooEC/Me+iu+r92FhZif/VOKVQzdSq2BDiWNgzRh+igDv4PDpY6Y9k+u
GDA3vrI//6xGCoDZWyzmUgc67nMDEXfJIaPivED1mSHUumUM6Ax4Lhtkl0hnVZRS
378NM0ScIIH7rMQNDbXLnoRuo2OhFOFIkTVq6aDtfZj7UrIX+WgIiB6j9M2o93OM
UaYwzkMxajiL9bs/1bvEx4I9aQSpdAWyjhhCyDVqN1le07Y40awWhXQJijhRRdB+
Pd75iKboxOgx8ckCXemCqWxUgqPYUG6KZwYsU/M11dZRrb7EmtHFn1tLJF/CgCal
SY/d495CfqJWd8lyMwIyyuN/Mon1U86dbzwIrLTACngCPUTZnSJ2TkSqGGnCQ0rv
1upbpb1yPjAQV2bmB+qjvAw2fNCr3vz2jQgfrXZ2h+vGHbyMG3Yb+HqxU603WiMx
n0yiNQzbE7OaQLfaJzrY58qJK/Ap2RttDMFt4QI2Vzc8bwJe9UlYVi8atze3vq4O
VC+4SGPkux6CRlneCPXs1OX6hCT9HDZG44iq4No/Q2KQSKs0RPPZju03Eryk3fmh
54FALe8i7G0qlFCuVevXRBtwFMf9cnKYd34XCbkhTxdYMIbPLxFVd4naEryOB2yy
8KfO0WMWaNNL5XBQ9vUCeE+gvXkmTAabQKFjxi796pAmhKFwESUle1JRX/x+YnbZ
r6O41wrsflU073n4KHP8a3HzrqjD7l7qntRh3yjdIOV4HNA+d2rFVj54UFL5UAbr
GNFO8fSIRgAMzpKKvuIG65Qip9oIIknod6XjqSM2BVa4HiCFutb0Sq82jN2+DgZ5
hQXfpb1WE9EGDZq1l9KoruiMFHjxY8/FiUsZXGH2F94Rxy4AbKuviodkrKfphX6L
FuJxSIvcEftojpKnHhw+wbRw/qTvDa/qryqhm1LoVd+Bsz95LyRTrmpmOtbgHCKt
iaV6CtiBiZ0cYN9Bxx8j0iaOGG3gGcYs6RG/WdCeo8+KJ/ZsBq6Z7BmPg5pUSROM
kQJ822s6hGisvLomSInuf9CLrIKrBp+1hghb/5n2Jeg5SjvRS1f8/9+GfMTe464u
YOFfJsnXLN+lr8kIVhEIEHe5vSV/LeqlNAvOScWhIDUb43Ho5hXGLFxBI4I2gu+q
JOcGyD7BvkIlw8JAnSsblzoyzvvQjETC/+Fgk2l8+axwHbAOvjWvHFBlhWqBmt16
ilCVS9C2sgTpJrZCJenr/UN3cHBTPDbjioLbdV6rRYbgPPqDAyWOcZg6dlrhD4Jv
bny/GfcdOHxM5rOIBozBGx9XZyKpefjYseAd3DfnYzyg3s2wCnxjHcZO0l3R482g
eyfG1cavlfdhNqmop4HtdDeoieE7cqWwp7WTjYCiATJGx9rHWaljlM0SUhppiTwD
dJ0dCszSvsMMBlJXY13rFGH3fBM/x4eaR1S0mUkk1V73rQCvZvu4Nk0KXluS/HAz
3NACiZ5AIRjOEGeqpbZF9vBAmT7vOWMlLrPo1SGkxvtctvak40mFaAVNx4UEVSNZ
uaAjsIxMJ5iaNaI6bq1FUCsZpoGgWdR2ZinXt0zkcRiG27epZbSpeHmBYbQMnuuK
mOBQLqCLqUW5wUJ/gk+XpYE10DctVH2o0IpY8tPAJqmZi0LFm+mNGa8mky5XJ3h1
khzP4VS1yZRD3bQXTy3oFYIXIeI6fnGKxzCMnh4N44LAzFy2aLUwfwd0mnVVUFGy
fqDpRBMapKZ/CJsp7DIKFJNBXRdnAME5lD2W81YvVbDRK9UrBBIqmCqgUIg0IOWk
UTcdkRKMcHe/4GK5u/m+d1Aj7BLs97TBPun8DEZIxFZunn/nUy1EItmeeas/eWtj
igTliWebVSf3KkwnpWiVZLjZoOyc/EELdHQZXQ3fhVjVcdixzy1lnvhIlIkQBzjZ
avIA1+nSzzwDh6x4kl5QB5kosXzyClcV15c+n4L4nD6WLrH0L/VQCVyTJtNyyPDO
Ax6EnnM4lxZFn4N/NP8qmPukEn0j7uEqpFKZXDFN3HPFMLOlBWeEuUq1QmlhcoN4
rGt5LYc3W1ZfmdM7wgTRI0PWhGmyjPWVzoKEY0cd70ds9yRuezVerpNiHZ7z63JJ
+UniiI/Erhrs4jyD0LBGGFo2cZ7tAh9eC1cybycmnfp9oe9pXHlQ0Nj+kfd90Q8o
8saR5wJfxToyXKvREnPojk6wUqXrdmy2FcdHj+ukcBV7mln+ijXegz4Pn+xSDBUm
fp5h6cuGeanAeojV4Gy/CQjkD+2/DcLmBX/Krn1xLX8EZn5Nj6L48gpzoXq86dwH
HuP/22Hx6awzDYYJ8x3+EmggMzR34Sega0PstxmRyw5iZkz36DgppzKrPSqhZJxp
ZkdHNfJTkhtFv6yWYmfWkV9eBnBr+r8QyzFShu+86nTGhUXgYACF9doacW9o3hdT
ytEez0F4lU6XgVeUDXuMWDput4j/OCUex/a3VMDmnrn0NeILZIk5LLxThwXkNP2E
nXntNvPTFnHDR/X/aUxyRjD6SUm+UMCNjmMx11Vr1kLQYsgMshhD/iTH7yZO9dn5
QaNA/q5crKAEG3dtFe1JhnF7FHK/xBwiD6G+fUmxFuu+uL6Fsgdlif1oUf1X5Jaj
Ke9AJlFyfYJ5Sh/INf0F17DwyU99xoDBH9FlKSF5Tch3+FpWNHVX/GlEtmKUxMK+
O2gLtjTDLDvRQ2Es3VLyEYNO+CGCHhlLu8s2Wx+gXDD4i4cFyRzF0PMyJommiH+q
095LErHQzZPCPskblz90SMLMvWUAkvJT3SAGuT9B1beH4OiFAMats8B7hB5lgQ18
OFAS/rqqvLqOeNOcWNLNxxT/+qLBqKSJFpTND0Ye8Wa6RosTatIJWZVz46dPBvy/
Z1ax7SmQ40K68O4JV4fPMB0l+tKk8B7nXMcBMhFJPsC3d7F3tieGNyBZWxb68T44
dyyojJvXns4uhPtQaFUMqZvdpV8T1FXO0a6+UxmlfFc/FU94z1dlE2WHMt3zWfTN
jMith3iFU/reu1iVhmfTH5JI0yyha3nkOAkF5EgzBHaT/gQNnhdIEYs+sfVKqojL
xrr/o/TVIZQGPQPcaeTaE/dp6yZHAgXbImTJsciQtmAjtwUIu9obKCKLSD4hK5Vf
ij403splZIfizELGrmo/J/vSzMEGJcZkhRaZVfCfswcasz0RFDWwWHHjygzPbtOR
dUUWh3yt+ZfhMqJDn34iCJd4E1D2CuwBMKilgtbg+7YdbYHYfdNjJJqxTYRkYtvv
yZxV9TP2LlW3TK88FdG2T5mA0i4+Upc8KYJfKPH+fyY9KgOUcgDbmiwHDrfB5BRc
G2zkLp3VNPbNybl8UdKhdci7t1pLc1001kKL+2K3gPb5AZCWt9bb56ql9lUWAe5c
2eWKtZS+A3dbwp3DJJjLiuTWWiUZFciAZuP60scuXqjLPa1saV5QGfZk1k6q2CCw
WWGjKPF+Blxb4zCfJsaNTL1d/FqNQicljqXLG9+wzHyxOZjt/+p+o63zo1nkdKfC
FA9b9kXcz82FeGJ4z8FdtMVz91aVhHxeGA/RyScIJXFyaD9Chd3Svbxg9uwBq1Dy
jTOG8RAkPQTqo3By+A5C9MzrCMrR/kz6MuJGewbhuAmV77U6hDSwAu+7rd4PT1lc
IO6FroMLQLuoeO5Oy9Ls9NX6S2zcBSWZzWAYh7z0448YvcmDRjwim/ww/pKuNsh1
UMX56iRdVHqHUgH4XOgXFHCuELAN+y7chx5qy/kqM164YMI9kZNxRvBO3H4Ly/i/
jOD63r8qikBb35uAQLbl4sco11p8vtlwhKVGxfJuC/poWinyfq/syQBtarGT5z4z
AcDaI+rz0XB1w2+65IYhhscJRmF3X35GgsbMKSdPFlPXPEkEty853tmegiGfZav5
iIXh+ZqQVTek67M6Hj+9HfYcpxT1ZCbDakz8XWywdkfuekhnCtYDCjsg2mG0tX5j
UWDrxnCNvXLm/1eZOjaRdb6ric5+D9dZb9zKw0/dctFPVsVR8hFQYr5xMDwBtorh
VAH01dPkJ3DBSLlFVXTrJBvwZj15tt6qgus4o/2SlDcwdMNtFGI7oA9xGoAq+UzQ
ay0s4R+zGk1MUpxohbA9v8g7PVk7Mv6KjLR5jRoV4cQajNclNIFhlabJVu6Tc5v8
YsyyNz7qhINnq5eijeLvCCI0ZxfEOYYAO2g95TCgoS2ukqtFucgvYR8ogGYUsa7p
dviIYyu5Rv/m9nVbZc3xXZcIu/mgSV3hDjw7r9s6VNFm34TAQ943Xp1KoQaD3RGg
OXzeRZktDbx7Y33lqFMfP+t+2upyQ9HDS2NKY4NsFZPtsYW9/KcOODqxs5KaqQBQ
Sz7Ev+SH4vO4i1d5cNSKYeBPvO41bzvSWVBl9kz7dZsy5WyiL9ot2Mruttbl9LZS
hz0fPzrNgd8a5m+XLUH8n8S3CUEBm0IQ2MDKPxRdXzxHGUM9ZedqQq5qY0bXKciE
tBP3pJavThEPVCaZT2wOZqOAkSySGfGmjqCA4X9lgXVcyXbUpOGQy0pp2rWXq7tl
vEcvQbSuCy8FbD1kuepyJ29pbTe8TjGQcq2sXnVtZEKPYYcxJxxaSz0Nu85o/kTs
1b0AKizFJegmWvDqd2+D3k53ozV/+IaO9jHTxOwfW2fpX67Z1icL//5T51U5GQBx
BMFTXkjAjPHC55EU+xmku3VTYB+/m1UbvwY7QZjf0+lqlqjXXP3wkOFWA+DQpuyV
EFnrHPClq8yO0urtTqqiU1qJZr1mXIq6XEW/uW0cQjDlCs8SqZZk9SYiPV9Wu9KV
oAb+Z3JFoL0txCsla1mRqovu86dD5z/KpYeStkBcdvPqMzziqL0qPagDo/lLkxoA
qV2j6zN65eYtr0Oiv2Ry3WUiKmz7qPty/f+3DDE443pmJhV+CSyWmU3s1cRjPgsa
mXqpr9mZls6tERmRNPVP161oc4Z6ldSls076Rfar+iJHWPxvK/WzoAaZOICRkQst
mJMXmUgrOeoMQa3tMjk9co003JAMsF5fio9fzkUw+3U66ANC3Rn1JoYO9M6I7t1W
oaxugDvQFCnpvoXtILsIehyAOUERmAPlgdld9BKIzTUp8rSE/u+mMJPoxqQV9r3Z
b6mDAZ4wBeT3TkvE2DxG+gkQJFplZY3oGjvRSwgwm1B22yVdFc48lx3mTjZtOmHn
7FAdwJ6/7TfJ/noDLFcPUrvXg1+iEHyVG31mAvnizVN/8jz4N0+AKb+mzn/TTtS2
8qsz9td5sPTo7Naj4Xs3e7HBOZX2qyTup/YiJfwRY+k7ONwDJ2QA2F0a/kSWlpXW
ST7n4KneDTSmo5VLtf1cUvvJ6jzSGApKd0G8Ppj1pjXJbrkqYSXzxT6a360chD+F
QKgEbl8dkckKTnrHh96mt6xBR60a5IemgltKuevswYJX0FrfFmsDCyPUXf/tFfu6
D4pQWzyNtqLeKFzDEZ91ton7UtI+rsgXAKCkjbkvRF1l6/jgYAzmZtsPz0XCRQiV
m2BiDoRGr9rOlvn1TgKY3MxRZ04A8am0G2mqHWXoOrioE8gNXwlQEHddozADmlVn
T2OG2BXHojQB6onpwdqFP3lAalKIvBUY2SGo0dnMRIWmzPosBMapOzzpmPJCBOzj
Eia6cdywwO32S34YTBuhDJR43LO5ngUq9YSeuUwkKKzLe99H72DI7ElLNOO+MuS1
mQupIGS/KH/E7qJke5ZdjApB3M6biMUslkizKry4iM/XmJTdW37sLQyLf1dbPZCY
cVOboJH9QJW2BF05jefiu0LGFf39A0e9oivQ8ZSIifr7Sb7ClObtvNoYwla3mrh2
8LZEaTP951X+LyHIq1Xs3HMxozy96ojDxGf6yQr/RJ+fYS3Uq9ZvVYN17PlaH1TU
E+CKkHhNZwjQCLZb/In4Sq9I/gdkBfDV3fMYXO/TpUH+c5KHxq9K0+zKYX/XDmpS
DPitXZ3cneMg5thMe8X9gmMRgxhvBHvpvXZywh3NL/KukhBIeJhnAs0sVezyTugY
UuEFy+lF3kST2JjzBHS5s2wVbt6X+AbGMvupJlZHj0oof8VN6GlEmF4FZBzO0DlN
799xaiyeMyDLU0YOc2Msl8UHT4og28KkUvQPqmi7XHtZ0U/ctqYRpbpilxdqkBie
pMqX24wlDLETGM5OBE0ztNNlKQUroqswTFiT5tp9d7c+jTVwgSI1P134d9+sAg9C
RWRk9MuhhzHSCFnV+f6bFWlTCvkTqHjjmapPIGZa6orqaWM/jsAbRkALnrOYwQD3
jALhI7z+e3Gv+ySlmEtDFmZxsyzwVhHTk3VzoEgUNLCTrn4gWKewtnyV3O2c4G/3
WeT9byJOZFcRHnYkyeksIkfqRGxLrW1zX5uKJPkKmuIRJeTmroeN3CqFYH273lFd
hiAoelQuPcu2hMKcjqE1pLH9CgwY976cnGbL1/p80ildrAkKL3eEr5qlEeVqMtlI
r+0Q/SkLM2nWwi3dcO94IXhmf/VpgmCMJaFokOaquhBIvXWfAyj7wQXbsEosg7ad
xKos8Hdp+FM0zmgjSxhXsvMBVfazdUTcqYnhaS1Q7MIgYa3TdzJU5VaSTCmBFsO+
vyJWBE1HoZ36IjNOdXiaRg/Er0LC/GiKzOWWpeR+rqh+0zxJYsD6/fZTCQxSTe0y
nudv3opx3DJOTTeFh9ioP/lAEXwNR4y/CUCq9Yeb4bPYrjDhniRpXzTDPk0Y55oU
o6M+AZhrhv3Aj4vfxBuOD6Jo/L2Y7l77WxCEG0WI8XWDZ2g/ewJfbZXtEOxxt6tE
5OM4NxHqHQ9mNxAyGlwsi897fpDajpoojpHsgsqr0ph+zs1y4ecYB8CMvqfLQnzB
vK7fWjGSlwrYaSftObZvt1AowTbpefn+UamTTRkINmy/G4kyddYarWpjbX0+6raN
SQbgb/qAKgt1IVrgF0f94y7Rf4Hh/GTVxRRTnaBuWeVBcqO1O5A/lkObJWh9lqLH
aa12swi0px/ItoFk9pr0rBG0U/rw0EF05Q07PodMpKvBkdr8zVo7WsZLTbDLpp/J
0pb0WC8OdkqK8EvoBQz4i0epIj3jjIhWUj+OVOOUXrgJcMrmKeSe0rxVsKMWPtRO
xuzwIDDZrTBHi0nMxeZFKdsioilAeNOZVSk65+gYahuMHx64xpJBvfZ8v7py5l6Z
bDzoyzqITU3VP08ov+RWu40g3G2cn2i+0vs7Eq9ggPc9IE517G0euvKIkZKtge8e
aQgR0dupZgptF0U8jzHyiNbREiaCPeCGosHDAi3DcqMOGC2PlhmAH+kp5WqClB4i
921ErwjApaGDGn+0lRlL7ELyZWc5ylLqLZi4iDUMYcyP7SaRiwpzHTA5K4xezphM
YClT6Q+alsjz0vQjNPJtuk1cG6fFQkH+G4efMpek8mkQUWemnsG4WoGxopyOKmlP
ox/nR2L2jb8HrPVXDSIkgxa8/Dd2/h7lxxnFnm80YttOWWtdoQuCfPsFSL9NyKfE
j+RbcnrF+PsqaOOF+9SOR+0YrHlwHvOs5AJTHKST1hDnw9kjxiHC1Cnkeu20acBY
6iDjnLc5QnF/pG18gKN9BNCF7lmIlmnbYcMIRQ1oC8cNNfeVCBYVXeAEtBpdtDyf
BMPpKx2ICW+RKbkkYcfk1dLunHP7Lo82R+531fHaPSqvzk6hXXvfjuQ82H/9/zrG
Glb1JVOv4gR5HFnuWUb7Brjvk1ujZjsf5n4WBw7qUzzNbWJ7nxosoTu93zINjX/+
PWcgQB2x2vPbENm2kq180Oea3CSWE1n5XtrBOK59zqpeDFB9lt6+N5qJ+hk/Cb1t
XF/6nBMnqAE/LrXDpm0h7hcLAz4fSYqzeUbrOsTJH+V3ra0SWMpv8dW8s5sFQd9E
5hQUh08C1yxb+FBTq2/w1VvJ1L8GYN/t3GNDux8y0KPZ5vfQar21WcqSi+zGVBpj
3hh3kzT+H3dg5jxYGFOqRoPlOvEGR5jqWlWG/dnPLgmKlXi96HPSkhGkzUL2O0er
gj5bts5iZ1YuBk/XqKmonGJvbUq4l25PwPJVtNKpL7blDlo4pAxziUmXU5jHZ/cx
74Kz5ujWvzaVqCGq6pSeSLGfzRdJbCnHJ9jDYXtVWBZIMnkpTpYWRIRiRJIB9GaP
4RNElk/tLuyRGCTSNflBfbFVYGnNfr8zTM+7rZBuL3vL4hd2VWW12uxKekCfzx1/
HEIfAiwXgqz7B6sbxHAK741la9ulCrRfwzNb1IZtVXJALAHSY41VrwLL2lmfaHxx
ioV1/itccXL4eNtDctVzeOHdaGx7PWFpy51NJ9TqiW3uEai6LqP18baPAfPIKL2k
Ir0PzyyAHOJF3DLK0ts7UbmA8JG7c2rKukRTnsgQ57hD3Q1IoCOPqFDTX4mmEhlB
A3guksX+a+Y6pypXfsjBtzY56Ydle7igC/APY6e/94U0CUvYD8yiDErDVZi1zgeA
vfO9lTIHuplWQ+nA0HaOga5ITG3g+3S1/WzCHxGHlclan8D4NvlBLJT8yinpDn+Z
8wyUvnfcjytPlBvEs16JzMdgLZgm27n1oa+B0VMsPdBe9bSmOF1Ymvc74/ureZ1T
Bnjl0K1wGgmKbZcbxaA+PFepxe6rK1k9cuOAqUnmwvlGs3Om+kGSZHRJTjOboxEi
qtQNjuZUDWQ4UEB8+SLyOe54a70c392Fd6h8iviQqY1NqyIzMq19nalcYGxNuSAE
ZhZ5dVDXeiXTgPopt/XratCW1UEc3fMowjMDyEq4X31hAYm8dAounS/NgU5k5kHW
Yjgtu1Ogl8BXFrVWY3B6lNbDSxgm04JNi0bmk/PlZ+NoCG341q7scYeMrEZk+tjl
aq/H3a5ejMZM5TTmw0IsiaeWHl2X4ccxJ9C5Bt9SE6qR9RMA01p7R8DpDfk/l/SI
4kmqJ/Q2C0jysMVpJ4tod0lGz2ZAu+4AXoxnvRZb1/ObIpQkWjkVK0SASHrLuS/r
iE4JoO7YiPI8K42nSGfj6KodSSxAOh04YxUDsHG2Mvy7B5IgGgR5H0rv8DHa6Ih2
5+5xrh/3y0+vXiPHFQZ7qSY1OZpk5+WYIFUoZBHUxUHRjHhdymK25fostFelHUXs
oVP4BgmBoxtZzPljluHQGEtkMRLL5Kg6h6TsYw5eB/P3AOfgDHpnQDDzzk5tBBGP
EhjzkU0eQ9Hhf/FjJscrG4oWJ5mO7sQLHHPg2iOSMgOGC06xRg4KqtanTS9BIVO5
DZCAPls5Xs/z84iG7XYpcw8HL0SPVfQfFaUNVfeX4Q5/AfcUqbotaFha5fdUU0ga
rIX0hhY3kWt3XyvvMoBcbWlo+hYT7ik+QGbpocB20RIuHetXiajg+q6YUQOXiiug
T0BtoHaP0xVqiNPrDnc5In3zX4wQ7FiS2DTBIqYzo+SArJRUwWK25FLaQMPVkENq
fsoRzWi4IVkdFjgRTPa5pE7Oh7521gYshckRO+oGR0p9LF7fPTkLBIqkvSZeuD42
GrUx5sntF32xjMeavW77IyVDtCQm587IyGvn4oVCokt7Aozb1lUfiKq0EdPRreOj
bst61he6Ms58M740veFpZa45TE6SnTdenYzj+/PD2z3i83EfpTJUdbGLBEPoXySm
KmvYiaY5PsX5iQXypqkixbuhmPXuWwZwIMUD5Fjts0LipXhWsxZUHuPg8aiAjVjR
Qx2S8ekzCCrZXG0UG7AFBdF4IEMAnUxSWcT6wiOzqLsNjJtpRCMqoV6pVFZmnS+3
83IPyWhzgqftgbdxt1dYjedIR0YKm22YRZxpViMNC9GbqivcbAkmku1jDy+HX3Sb
r1+ZDpbfAl9+273kzeKDdk41uu7sLpYlg0DhWN4y8CJovcO6pJLVTXn1U82+xAtL
Tv2Rr7fJO56ulPtIKsl/rznwcrZTs3Dt01KL+LC+0RIVLq28DruGev8urp5sTzn+
YqVnQBEDUHb25/eEvN/OfmVRVlxd9ET+aZXA/ZDGhY/nwoEF49O8L5OHuN7QiIFd
BTMfgmTxBSd/PQN7kfk+CqjVKUT+PWqiPBzyxlPVB87Ro3L8YpXw8e9+4/a/aPpf
l5a1f/yObGj+hljGGwgC/jGffggf3D8UuyrOLvYvuVecc0QVWjThh+NHmFUjM0sk
Aj6xPtxobWdq1mYAXZ17C8KYwdKPBHHK8UtGsNoV1CUIoXFcqRhz1OqwNyxerzku
hGksgYZPmWfh7736YAejEvRL0WTVgr7Ebx3qjdGq8MK2kuG257tIYxMACibRdaXX
/6DhOSgKlvWCvbB7ln377oO2wU8FhjDyPor1lFbUvpMbL/uSlUODjZajxR25FJs6
LPRKkWmRrp5HSSfgcKNJe+C/dUMcDx5fxCq6s2o6k6cSmz26t8tDBmteHelRfM+i
awX8VcA8pS+KzeoZebDIIQPAIWa2M8dbeG7T0lqkmNmxlGzYzQly6YYqnfPfEz0e
+yOLUUcTc9ZV2l7r+B0iI3JjN/g2SaRkt43R1fM4rPcoVBaRf+Zjhg3L1QBENYW5
XH1X0yHZxEaEHyH0h2U4kGZC2xzJhqdrnDWPehq4XAjiqCCCxSwgtGWSDTZ/8fcD
V5yvoGWCtrQgw0+Z+8V/ls0xy1TbbLy1XFMQOkyjzGZNabhCy1pRl+Z+tqtfFQwP
w2Y/dgcRMyRrZNfMl2uob2aSKEjCSS1QLa5NLCNU8XfKcomP58HYwLLcyCFIbkjH
uXgqhWGINB32U11SltGfwdmzdwFRV7Um1IGuQCDmzhciHmclOTD85ZAhqdl4yJvy
XdmyJd4DvLOdffkSaWnauSlwIjk/BrlEYsVi105P/I9B1ljF95Ef1KhmDtdAcB26
JESAHnJMURQxCzW2JdDoECBJ8jatZ4l95858yPo5ZFbZKHev6Aukmn9Lr3gseTHM
ftAfD1Iso1Qu3HLrtOQl/g8J+rGMVh1sIs3NMsUBmpXYQxnqSO/qcVHDsv7XGwQm
KzjIqn0vQdVRtwaUXEUOQN8jCiOOqP5DkGhrYcigw9+7AEo19g31Iml0wsql7nbI
d8Je7qQoSwuEmoimtBXYTx6gthF8XFdJl1iDPSS2+eLz8Vji78l8e66V211kgJmm
EU+iwwVOb2+Q2JKlc1+gz88th7wQm+tO0h+nkKypxZCqLfCOXxxCrsC1bP4EfwNx
mRKglkGlXswQDqoWEIhP7HU8nSvjeYe6Za+RHkqvGodUcLrWVdhC+MdYW369cguO
+f2Jg0VYw7T5hohb915k+n/KGSoIqvDGqAokKWJqQfZSQQOe81fOdysbr3crBgay
G9sfNoWOMBCm9Z/cVK6yhMPQ0+4GWX0mRFP8zl1jZBdu1pgEgRE34ULi2/rh3LbD
yIncn9a5rTKiyVHRDCSWKtQ5F6u3grLu8W+8u3xeoQBWoffQ7Glwpr7KcQbwJDb+
oND1CslHjmk9efhY7FoIi7MX7/H0vQTSZaDL4IofWLqVC8Jpuad78Y/BzFdYQRBC
b+1nwwLDFQ05cPnNKCQRNtuU8JX7JhGADran7sOV/46XWPHol1mPfoAjgNTpPvv+
7g2sf7l5EyAS4jsTC24n+OgSbW/hSg5jr7L/PK85t1/z4wA34mFktS1D/8i2nL+B
2KW9NiDEG7KBvciknD4IPjd23c4AaKicvD8nRZLuzLXcJ1sX5IUm17XqvAYg/nol
y9fuiEsdD7+A42WQx/7fib5OUKfGfvHtDb91Rcw1b1lD/LZs+sXCY4kx3JYRmiji
Bwu583g+DGqaABKLxWO3DKVPD2rLQlhKrHpHAhT85auATeAavgp+PydMOAmRIOPy
+f/vNKC17fXJfghTw2y9RUxiDOKax512f3+YdwAaQicEAJMqGI2veuEBBu1MiiA3
U3baP9aqFIaftb1YGW1o4i9PmwELLv+sgI4UhTpV6VkwzXsjrGGEAQzj56gjfPjQ
q0hEhGJDppkJzLureYzGhQhtOcMvRRIpnCec1c4tQ8Zqukw7N8+PR0ksVIFif2sT
OH0ElH0BvCJn36pzc/7WUGH6lH342HXdBEaAnKOJGUpXHuyxn7OI6HrZK3J6LXRp
TRbs5TDuDfXiaIwBqMfsaHlnAr+NVI7sn5p9DIHLyQMaaS6wTPp++Swk34Lw2s3S
VbLNq99OHdKkUsQRt4+fMFtOk+KtnP45DrraKShL1yywt+4fzJNczrrG2hsl+Lbs
n1wlU+J82MoqAMQLpN4SfutGfFt0lFqMfBgFAue///Q2w3wWiD+0Byap2JoaXGL/
VDvg/dfrYYnlSCzKGuLvzN44msIvfqHrUn84egBCYkaNTDP4aNZP6B7j075qC4d2
jLt9QKnI6nEq9PC+dDk4ydHGBSv804SOyp+g/5MmGoBQnHUBD2sSjIK8knR79xgc
rUZDOeGn1FpevEUYs9423XYiyL02ZBcZyXVeiEm9yogOQsXgAkj4+m3pbqfW2yGY
QAy3BOcJZgeNCuQI1LD11Iee5xc7yFobj4L5E/W24314xJGt1Eq6jUHd5wYqLVwK
ZAfA15ISbH71lJe7VFZtRdvyydrUfO4yxV0bFC3Ie06wV/1C41N0H8jv0lSpw4t+
HXlfllTWfCh4PNWvKNHeQz2p9lEF00hZnOfCVjuViKZ7MlYP1RgDDHm84CZsdBcI
bF2R90JwVG7SOptoZyzKdS4lOzsUqw2HfXy34RMqGX3YI3P7pGb/EMTGl7zyJtXN
aygmfiYug5M2z8oUQ2Srypi7f15txU3b1l5jD332taZsixHSo/o7necRFD+XiafX
3TDCmNw3ZPP/Wtxgw9/iqrOYlUS2jr8g0W/bBboSWSi0LJjFWg97hRsQXXA/5o6X
KkBc15RPtetLOsSk/eOct9hjgCSQxkTKo74A/LKFRVvcOEVRW/Izl38eFsin51oB
/3Amz6IXt9lirMrjfH0OcJZLAmrG4CPLatR655lZvuGQpwyckNOz3gDWX82Wb8VF
eO9i2DE11tVPT85/8Jv54GlGvbFxjV9mcvfgATGkvVICE1L5LnBEV4nI1jAHGvJE
CnbEZZcKl8FRUssaDM4Sr5b2o0jspSyHba9dSbDhNOF7xhQSEScmGx558gqYF979
nLs/2y+52WATnOtdZp0YgaAexLupCKazpkpdxMvLpLDgGE8ZA2pUG+4lI292ZPkt
ClGC0Z54205UcwrZ3aidRF+6LaQqL443zcGG5A24BYDoGm2IJuTTfkD1fxRveIRU
Kc7jj2XWXkppc/TwyqcBZDRQpEVUp+REjlJKU73Gh8HVLmToBF+3KE4PMs5kZv3K
Fiz+4uRUTjX4im5Lg+fbPy3OkIpTj2Pzxfd9n6q2ANQZAZuS8cl3kThW6MWmub3K
XN0kwRk9kpT95keg5rQOQO3DTpK8iduuqE48djJy9DDQZi8eXoYSPF3aqefBHN1k
e6cJLvbiA5vsmz2K7D2BqcDnAyjw2ktLh3S0fSCIOcUYrtft21sOL12c6WRd/GHI
4hEJlLB65PXbjbFuUGtGGd7hQXe19Helb2NmrgeVpnEKDV+uTgp32Ct4lAdPhtfk
hn99V+aq4RkgYMsB/wg0s9QNN/U4WK/lNY2HnxiC0jKgcux3TJ0rStjHBnuO9DTV
njYgHvbifEix9dPZuuzGV+egW2N4rk6d3GmRF2SdZ/vtovhx33SqCBqhEl8sFPFj
0ysqJG38MQSD4orGvdgamx2E1bP9vNIZV4jMPvrbZL1zQaL4aZGnIVPP0nkHjSxA
SCGHJ/pZYuszSMiZVL77vPncBwy8xX/eW6b69VtXBlOQ5Yh33jCAq12uHCe9TQw1
w6/mJ8IV4uBRE8+D5SYTJDnoc2Olyq8EjurmjkdikWHCvRDU13zNWd7nfu8KEljp
oKLCHYm1De/8ozzIm5WpZ6oOtLqtrUnB1/2P2koPoE3qmYmdUt331CdQJWNJDmkd
+fxVKkoQRHKdluiWWU9B4Z/QlcSk5TuReoqRId82ohzmjzkGjk84qERjP2YGKK7P
8g3G71/t1nqFh8Qz4dkFExeQfDAdSJi8UyGihT0NbF0LkllMgyiQ6hN39P1xSqYq
rfqZ20G44qOFr9waGNn9+rqHl0/t599OD3uKtaPaWjbmratFNAR3x7f27+F+BWlZ
hwSgRCmTTnPD/o7jACkr4rJjTJsuEsrGNUHK46vQZDzYTDg/1JSbbbcZExXB+g6l
5198erzryL13nAcbhRf/C4zLMurQSSNStmJWR9hi16pXYdRZiyTLfxlDZ5XaVWCW
56yJykWGYOlbLwUeIPLW+ac9pxRCWd/fP5atXIYynie7JIy2slXhZ0Dafssah/3z
9+wm7y8md26N4+K7/MMrwyH6H4ev2f9EQCsjF5r9Tul9IViiIOgttzWkOk44NYG2
cC++lAB0OgiZ6b2XnAPHbv1E1KpbcheVJ62bhmAj6vLvRitj2BSnmxDHMXyWIVmw
ql8TFprJ2bDEuIEzlB4PPMcN40h1h4kLPtPOCHE01dXz10JYfDhmbuogCK2OQL3N
aNoE3RmXwzGo2005luDbirEMKjA0b6CGvXXgPtMwp5iSjmWn9qAJlJB+hxReMjO8
vNreLhtq/Nx37wfRRupEv8ZD6bLMmBqJAuoz6i7hVxuXkfeYMe+CtxcjvDx1ta1/
Nv8f1xu/PwY9F1bXtAoaevqr2b88K9w70N5mDNTdntdH9+hxFNMxPONCIggRs2FF
ZRYQNQHgN4pS03p/g2vaEul2+V2ydM/egd1YZrFBOzq8V+V+a3Erc0zwPx3PcJg4
5/nkxTnfXH3SQ6cwOA70waChvNXYU5fu7E1tHGnmikhx1fJtN2cPMzYwSNmpQHAE
QSu4bughbv72OS/hJhsfJFAwcJju56eJ4/GMyh14v6CvQUnv0qhLY+dsM/W2bKdl
ftJda9U570IgLw4KeJymRnR1RTNRhCiy02GIXCHgWlvZ9lI6P+CBPTF9M7b+wbBj
hBpD0tCFZ6/EMxG/MvGWcW88W8+B/q21I0d00+xtomj05x5yPxX17TYvYwsVWoYH
L4gExKE3TZoaMh3jx351Io7hkHNGJlE7WBXEDHrmT5JlvpPs4+9ORp+S9jWFJDqD
0gjQuClVgKI9NtShh3IuFx5mE73WYd6JgqLlDU1yYknNOKOWbshnvyKte+YzmOC4
Ux7Yno0aUyS0DW4UefOaPvcjN9Ut5zaHP1K35DcxNwo+RZFK0xMyhw12qsSgcwWI
GzRWLXWrGeVQ0NVbYdM/PZ+lYYgssmz2Ipmo8em4+Cxi89gDrYVam0lZVMgwMWlN
8l3wUCXqOdPcybD6Yso25/+/tmjCFlQ9BcRoyOcOl/waAFzO/RJ2I5LO3rVvsCwr
nFcOGQhtFUF6AJkaeUh9ufLHBGoIBJII1v25bZ9dyLlR6dOt62Vbl00N9lBGMB1Z
g7VwiZPZS+59Ijwzo0rnui7C+6cUVBaFP9xrTtkWgTsHdsB1mMrkEcUAUgZtoCqw
n/m75R7GM9vDus/2M7249/coOSc++c7WEH5XrCWPMzDmMbtvaXL7yvdH7z05GTNx
9dvcYXANw7mNAkOChmpQoIhb8cmVqpE7WYSwlArgkAD8E6sVeiQxEOmVMQYg1NjS
XFQDfvbX9F/pXEq2zXAfyPO/N7lyYZ0e+dbelYnQRiQtN7ynhpnI5bgu2tY8Gcuk
7H2QmViMAHW9NsloC/C+JwjujP6AH4RzZFPuT+rqElG7aT8qXxU8YP/B8bSUJRh6
nrRI+EgAO2pHaQScLE+qRyGtVus6YqDRZrPYPJTYjx7Q/goaa3g5z0o3KQz8fgQz
zsCKIHJ7iuXOaRHKG25U0e2nSIAENZag92GhPoJD3EevXybqkx9AlyJjo1nov+pU
/7So2qe1SWIq7rCKgQXBAgGvLf1Rwz964dvhd1pD5UsTd7FgyDje6OoLvkCL1pTL
FOxF2AxVjjSgdKX8IwptjUcGMcamiRSANfNb0N9WYvWiMm9mf9hbKoJ77pFF3vt6
zLjsDCV9+7E70xO0rV371HxJn33QFaJGw3iZMgTG82CHBZTfqExz5Fx2GnAIjBPb
UPIh32zRTxThSRwJqQqzV7qm5Dc9cKO8QMypJrhIgRKX9wr7Bx+4n3a260euv/v8
X3celce/Jud3mj1HaOIwX2/GAh4PER6HCO6IWXkZ6/P9+V1XqKnsr/8X/D7CYUij
Dc7OhXSQ3RxZWHfNTl6kHta1uIdU0oqrzKT3hr+m82SNIBWJHve75fM0g0IpU5bY
0hHv0mIIzITcCpGDfErCp/9oybjau+DetGBshG7O37GjaL8MJkC4SzdlQMSotCkp
YMY9zYgTF7WFJQEuToKG0lYn5By7iUPFCMAwK7rjlr/1X262Qh9UjUQJwOmj/oSL
PmJ9YXivlOMN6AYJc5Xcyc1k5ZEgH0UtI+fIBw56y9gqB1RPS24QWeh6iY4e6jYP
o14r0Iq7oqGZqL9blf+285Ey42nB2dXloMVHPKCDpaLVqo+H+N91HjM7Czi0lgrU
pwTUqWTG0ehx/myMwqTEA3hQQL2vjpWshyoQIsOUOfhLUActWNdzZqFo8E63DnKT
zIhT2/gazwJFTB+wr9igGWH/Vhj4OLVEailD7iocyXwAPQZQQ9Dt98UgRFqFqdAO
OSzOHK0+0PDpSJBqVLn3u7GuwlVa9EBYDEjFWKigxYyT2se05ZnHP+9zW8sawSjJ
laEeZomWUXGEmmAarl2p2ZYXxie2439py+hm5bikD33HDyg/xn+lSVT2i1MFMEyN
iUOA/YCLiW8VwFTYgqId5PvoUXqM6vI82aCO0Or8icLz81N11bmtV8AkPV0Q83e6
9/0SrPIetCNeOSlB2RE9PLPea6xV1tw4Z6NfjpdPzmb5U2U064w/bvaMa6FB0sEn
YkjtvkLfJfygLKjCT0LELQ3PGCKCpxPSnrijKIyKLmO2BmPTMA+KPV9pyZYh/61F
oTYR41G7KrdHGvxM4RTK81J8VHcc1V71/VDsVT5p/VVNlWHP2N4MTH5Le60KIso1
Symf+I5Jw86xEIGMgCTfGzWiP4KUfb1PI+VlXbpUinMMeYrm6e2RJ/QUfhyDtOzA
rnqrbXOE1kMmBB/kbA+Tq7sraVu/tseqvXU207RSXsRxaV4c/i4S3ZAGe3GKI2zg
0vkcXpfarqf92GTzEmDfMTc/hoaL3cB/cuudgCFYm0L1kB/qmVrVj52bT11xdb8Y
C6AIUBpDNPk3XccZu/wRd7buoVrU7d39yo+QihgU01QFKxMC1Mz3+pvSnIyDGZzd
9IbxUpMeRag+drfYIUuIpAnS9UvDJDBlWQgDk2CwRwK1iGLlZutQMbP4bAJ3T+m1
B/B10Q0fatb80izTst8vGFTOBEp05TskF8ShP4ZffqbLLgFv8J28HP7Tc8cBeF0T
2+cr6J2FMYyTBCcAMECy31vlb/oix0/HnTF+FidPHlHrIhRV/VZrplbDU9hYTzx/
og81+NeFoSkAo2KKY7EWN2gzwfn+/HgP+03C1Okr4+BkZme9kJxAhkQQ9EULitds
Wi48V+PttoWLcFI7kP3hgVNL44VBDB1vh2vWTQHeVV0oOWocymPYrGW5osPgTSnb
w9XcckkDghDTqQlNQGCJ5iKwOWgJlN0ShXaokWmbHZBL25aPFmkaLkLlYTEkNtfa
PmkUW2A5I//FNJ/EHvnVbFYaAaOmnIiTPB/5EtYlbUQbtSrZU5Q+LM3xNrjpZf1R
6mF9c7wAtCDRsAgZsWwwj0Z4TlBAV5a41lh9m1nU7L8daPq5tV1ZYR6aOQ9JzXWh
WnQFjqmXduC1tLcTDbhHg0zHZVAl3Xv15HHSbg+Hk8qmWZT2nSmP/9ko6eLeA64A
u4PGyCGya14uMZ8h05zusHdI4AMmyrxwFyDRx5lkQNgl/i2DXBwmiOPTJpGG1uVh
e8dhOWYq84zsc6nhWXyjTBEh/2SbqHF7d3Yye+q+XmoE2FMECwvE5Wb7Ej233Z42
sHF7oY/LL7GODt0S9WLzTSARBhJTdJL7QjZTVtLllfOTrIuzXoImibwd+ZmtC9m5
KUfjDAeNT3BHUS97zLFAUqa4F1Icvy1n2G7tFFBJA1EWA/LWOhGssf8D/VuWEYBa
itSn2qe2107jQHxAId2DAb0OswQcIBnjwDv+c/+U4Wtj9dNTnG21YyTn7cbFbPTu
1k0Ck9tgFQxjwfN0Gzm/U/Lqejq595DKWGEm5ZgozjWEjqyN59GTfsPnwAHNfA1x
pvsxnq6T5IvLpPSv1X3sh4ev7TZDlQPdgvyaJKfZBj9svwd+3/2RqyeceQwvueOd
q7cMUDpB9KVhXpUNvmOgsZUE0mRQem7UD1LM3r66kBfYXjh3o/B7a3E+BOxgfthN
NQqHpKzsfnE2MPESMQBinInXkVFnRBbZqeIVwpUwlSKZny7ONLrpr12ff/s9Y9oZ
vZ4bCka07C4TinhDsKoyQ3pkT4DZuRJ43UfUjZj88mNN5+O5VrutmLqVC+26ieQU
27i0uTPwHFVtIXKg2hbGJ4YmnPVK6QntZO5+p6T9VjYYko99kQArg5lBJt/mqlK5
sOuQHsBk5CbtaBTcwCEHwzvCyzzTTTvFdW8z1ctdaRCNDuqP0+JtCzkUm94CiJAY
dsEQ7Z891QpxBZbyNFgaXGdyhrg9eCjSx5ZQCW1bKZYvnNFczKJRNNKOGSVRosKd
0NhXCVhst5oSwQ62Okwr3IStUia9xR/qurEPO6dq7/qUDhfx6q+kO2zY86Dr+wAS
bN7vhKOSxk5NHP0R5LO/L/GOSwnjBt2wYVYpGgZ1cGJrZwzDSS4ZWmoJOr+Y86yv
dqhTrkQNOihMhZOv591qGUI9rU/JSKX/sbJkaf/PYzFHo97ML3+Tui5mpHs05do5
3pXofd/ZcUMtgduabtf0jlQlorQyGg76ptI7JJ4Je4faOL9cwlR/Pu3ljivCcHBQ
JV/hrarYq4m727hXKRI3So5nVubTlspVpcaX9xZ9nqbz9uLUMpmG0EjFHHrtjmc1
8EUpas6IdGN58rdhY4WmM3GZlO5Xx0nlINwDXHxIvF5b4G+F10TSyr8A2mz0MOn3
lATeBfbCh04REDm4g7x8YjA47+a8cn0sOc5/GKoJyHv4oUKqgFG0EBV5ihvzviMG
3f70xbQMyVr8dZF3f8xrcABj7jerZfBFNl8duhzAFUKfS6Ul5katVtbD0OOtcy7q
5h8obTmeIIyYgWM2vjnGDHNCMKSD/IK3BvnFhs7Va3JDgeWJvkJqqFMXh3CfVWv3
C8cmVgUamEyoDAXy9Mkvf4jJXtcU7WKtwYPKQbdK5SLG0DmlX2/VitpsqgoxVa8o
PArQCTIPEp5AC/GtJ2cqJ6QD5zNAp+ziBYfMPqiVr7sbnphNx7ERBEWfK+FupV6T
J6orj369zRs3dSkhNv4lKE5Ru6I3hgIlnQj5sm0luI+4Ww9lPqt3yP/xxxdJGUhR
aR/UbfuFbiKafRvylPldYuUdXud56MjUj+obLs4TDLk2l9ghtlW5ipK61depdnfV
K0YExh5YTibSD08+PSBOKMs1fRoP9hVzb3nYe3Of+E3XSv8X/1NQaZJqdwubZlh0
/4LxtARyhviHxaNQ/8YbWr74HxqR9LyiDnyY6LnX6Zi+hNyJAS2DnS8DXnCtwk6L
8frHId5HIVnKwrsBx060Hv9AqBnNLrqVoXtlUCzEp94XKxNbDjid0VuT8EDC6wSe
+dd7ALjQwG09Ckad+8UMUlpd4XO1YjdlQy+WzZFy5sFaR3WFzCYQzWtw3oefdxtk
KOJayujInxq6R4wEKAfUHY883H3yWiftc+wZI+gMPZ9hXjCcatg6zfAls53+cBKG
/8po1+7YRTLYbK3+XuUfGqHPfjh9BdXKeW4Zhny1MIv7/zGvbE9qICkhCNIvgNy9
K0QJP/zK6D/k4CX5/qPQDYa/MlbE+g3CSM4462lLWkntPXoC5GhY05dY7T+C0TSy
GlW+MtFwwMW+JY8hHI2ilRQ4XPJYF/nv5wvdhgqNp7eZS2PSq9X3mpydtrGSI3IX
ljKdp9Zz4j4hzhR4aY6dYJYtARO759EslK6xGu3Ivph0OPb9GGOeeZEc+vo30U9L
bUGd9A6ZC7c1kn0zV2tcU/Ak0ugUtCGM4RuX4OnHiB6WmZ79uo/hwUPm99gLIgxy
By96m3oy3r7AB4YZCprFhiC0Ou9oRdwbzjqZHqnYiDhdKBchRedDdsMrshoUNDQX
juVaE90i478sgqVqktalWpt1evwUO9WD3ImdrV0aBfsOtfUw3xuQtIDH/g2oTofK
Rl4NhuOI3mKdwqIPdh5dyU8JKIWt8GAH2VWAFO08iru45NsX9m1o2NwZFLSzYpaz
sBD5IBNWuQCFxg+yejUKXN9644JEMKngNtK7edMfU58RA4jhUcSOoQPlF5r6fGED
QAAmQQCLk/mrioopPjCkoRGs4SYSmunT2MvebxEG19ztiZC+nte4IW/9uPjfOUyK
wujGMnoh6Wnr5ebQlBiyZ1WbnCrmNADHVu70OBFN/2/CJUWw/CVN2P/I6fpduBmP
xaxjWu6cxMR1iwS+1AWfXLlkLG49Z4hqkZX/RjtojJzdblEOFZe33pvJ78wrnewI
SPhyJqCV/Jyj3DFhDxrVnZiqXPzlsv82iebYThvgeOK7QtBxudB2pK5jEL0n4NU3
jGeSZ+2gIqUk8fbcrIriDc+WoYVqMiUbfhwd2Gkuk4Y3/b845Tm/D9W2JkFJmarb
YJqsMl1s+vVT4gfehSwgASmh2yur0USrpgb686yn2mkBBuMFIuvwJzfJcnY/DH5K
bcLmOxZJGhtMlGyYn2Khicv4VRAi1RwJGmtVJYbseoriEJAyT1wcnACNMRlZ4/tR
Y79fJS/2DFi3q7NszxqqPIBSLrgsN2f1f+WzK7UjIqlE+86xg9lr+eLHaX7Px0Bo
lkauThe1DwRzjeigXHd34mBp6lnpbvbncMe4QUseDSsdBUzyHOC+Vp6ieoNPgl5y
WemQHkqcoMq3Peycif6VwNwPUVEoup4ghVwBzv59pYSO3td/zbAwEv4e8E+wGAGm
RcIsbA4X/8mvTVFYHKr/PObI5qKP2S4J78v6MeAmWsPl/4TctZpJfEVOWI0cj6Pr
hoxQF+cfQQLSRbZnMaIYCW8PFsC3+Vtz978A/M6u3zOg3JuWerw6DIlt0PcRu6xX
f8fj7PneHra2yZu91aj5/R1fZdNhoftDPZ/4Xcrgh0GddsdbDs5B/6CZJuup1/60
DCg/B+kADX2rztExBi9U+El4pTYBxLMVuc2i9PYshn+msNRjvE89Tyc0tGRnU0CM
7srFhdQx08aXu5DhjyzzvCSBm63uTibMO3KE7bjh3x9HpyPid1OtY/B0iJBQMOpA
7RnLk8SoHpwdYkVNQBmK9qLVXlZOBlBdFAcw1hP5pG9qLSaO++L9OyRSdZQhLa/b
8dTU2u5++PmYqz7a5bCgG/NfSN6cvk68+U+tgBYFV3JgJszQpU8A3KQ7X8jZ71F5
HIiGiwnM91QNSoxzB6chw48oQQIlr86WiwT8HFa5KCXfZwfzdRzd4ybHoSFZSiaV
IQ91dQX4QKFQFlo5/URgwOFREikksf77xc3WaVGIsodMQ1hqw1VyHKBZA78H6ZMM
11B/EGV+EZZfx8/1dH5dm32PlIqKJjZiG/zW/hwefILxzBoCCAUXOalV+b2qPg+2
IOobU4AQat1lqs9UvT7Zw+zbpW2CEUnKdmaVEb4Oda+x8N9dnqC8hXnTUXZIY1FR
ADvjbxYsBUYj7e2kJQjp5Qh7lpd43IQe1VGwQXEndaCUK2Y5K9L7RW8YyHvPtbry
iJiQUYOebTqzm9xUbJdDf3QdUuJujhnW+tEkot93yp3tXleYLbrcgr6f9rDHUJQT
2smBSoGVfF5EgFyl6I+9Le4h9Bq0q9ZGMxvWNzQ0Zi7u9SDEOqmrfqckdKDi60Zo
KyUtUPlS+SdjugapyC0oKXLB6ZlVRmXv8ieyieuZ1CIThHYvzC6Cq4dl5guh/lb/
Bb2UwNA5oVPD81lHjAhpL/CrwsP7R7ibjqTCfarrnYft26sXA3Ee59GA28qnxqBn
6krSzfEVxH2tO6EYQKLbOUEyPHgtnmSNs+UZBF/4oOFUaTqs37xeG+09klyRZ9iC
58J9JAsqpSlAPgTDqxK3fY0rdEmE5DCpecQQyChIsHr66mH5cFwuA6aUc9Ze9Ll8
IT9zR+tsRTZCy1VE2Xih5u0AePx2xIk29LhFA8M8OLC8VcKMfxyuB652v9nmAPo+
xh3mOs4cYflwktu1e5MioP6AoAzGw6TX2YrDVSXqzgGiCC3lbV4xA5s/9sPNTuL1
1zMNZdB2M3nKUlg2vof0YGXpA9IYvYXtMtrTSaQSBwiC3P08VE5eNCZ3EzhHiip4
axkknbHbu26Ulh0NtNBkKvRjJicRZ2GEEOvSDKUYFC8rYaXlCbxcGV5UfYHSy7Uc
noD/TZ3GmXlzRdJ41CTDPDK+EbHutIOcL+zFm4qj2TBFYzWsKwZjcL706MoyFusL
GQ/oibbcZIke9ccMK/eK+plpsbvrzQ/EKqFhEalpnKlvnidq5197xDHtmEdiwhLM
ji5/Kc6sLW/CiZ32ysA3iBCQnnBJnvBVNC2rIlyscHdLXleWHe7c0wsVQYUqIT5r
Z/uWxDG2QgQmVjY49ihuPuVgE5+Ht8XheNFPyBhgs0gsdDL2M1cmX/HMNz2dfKGe
4fprOGWamnJ5IeQIG2OhKt2RmcVxRap/9AKC33KnoTwLyGmbX45WEVIJa/wVmPtu
B0uD32mNZjAJEwRXebNQBW8pgdy6lK1J5lYTTTAphGrEgz1/kJuEAEn05nbRtuXD
H2skRDXvs4ppfWWUAc4KXFV7YhyASllgz6gQP4zbHQbAGc8UBxVJaiXQhQQ70psK
nJd2OMiUNUQ66BEzvDse3sJiBHq5NEHQBj60JZfWqxx61jE17jalc+WjI2M7CsMN
PiT5xKdb5byNxNAqq9O4k2PzSAIQzsZblulER9nDMUzOGz2onePRj4zC1lddcaPJ
c56RDd8pSIA0jj2kGQKEbSPVYYQE4SeBSn4rMhpihwFLEqF0EQsnsGRpJLRhDNO5
wEbCbSFG+S7/P6DYc5U+XiinzODMj9a0kijsYmR9Q4XrrGOutuKQRLQhqVLF1aGn
bgXdfAsd2Qx4iNC2NcMzTzXBgczuC2VO8SKy3IKSO2LvUylomcYKgUZYJ9vGiNfS
9pc0kVjGigClc7NgdduhpizchaNtCFzxtSmbMme4RVzzfpM0u5HOQfG3lw+qP0w9
a+xMI2wFLv+0WWxPg7BOMN3Z40RW5lJcXSjzbNhttQuBs5eOWTE/prhRa481wIuW
v2x3XI+UcivoUt1WBeIWC7Bxo2fvdVCrzo2IoDiI9mV7J5WQL90r1fRvU2pP1RXJ
1Jerak06T6fby13yTTgEgTXO4b2qJ2HL0ND1clRWzkTQ1voCoqhGTVEUtBYzArbs
Z9uy1U2pF3iIzhxF083RTQ0obg+RY49h9VeGoIRholz29psMYIPMmeKgWBjQRXmO
pgvB+tXHTN+/VcuZlpZ+HAWYsclKxLffCj7tLhz+VjSWcWY4FTcJ1OgaonRJIef0
eaic3dRv3UXLG2R+ozspffIVImR9UjKfj5PFHk4LI5lWVIHz7o5ivWZ0WVfKKXPk
BpiOH+xVatWQp6CY1H8uPJuMCjakvkeeJeB0GGRZ3jPf1+pORUjmPq2XC7t/atdZ
o+rFK7xk5FRCQzs0e0tA+AWZ8wRlyYm2QOahXapDTummHet2tJz8I+fxg96I5b5v
6V8ZF4Er3Bss7lM0YkFi1ZoP0B8YeKQ1knddK3TAKWsaBrr6pD9yxj7bSqQEkOvd
RHPMnyrDbTr8h8QNh2D3EbMn5yxnTwX3wYoEXJmWMJlHTkiatp4Ig7LR0w6IYwVs
z4gYoAWaaNl213u2wGMq02DGgy2lEQRHXaVKUTOELJI4vBicPTYE+/lCcxeD7X5A
JR6WBuktEimCbBQAZ2ch4QwZ5INkeqiO8PSb8JNchVYZOIhwvAvcAm6mhCxKn4I4
uXDUH1N3ygPulxVkO4O3uno4+n8ztozxwVVTDjYF8l47OnZT1qDaum0XyecKeYs5
lBHmHA0xfEWnO1XDuo45rpGP3jwYcWqxZqGPrLNI+hyxc7O+Rn6ZxZ6AKyGp5cWV
LDeNbSb74N77Vhe9dmPEkA0gPYntpZQAzWnNDGgA2HAs+b+0S4rTgkJ8uGzr21/g
PiHJiVmYwN/CN7K5snkGO87kw8ECh3LUxnWflYdOgElPSr5hgPz7ZoX3sG6xLkaT
6Igk+jidsKC7lzY0Cg+pBAPzd8uylgGWoqh/PpfRN0LSAEJL3mkZ9y0htL+/F8aY
tJlTKyD/atRSV9VeFg9kkbhqR4Q922KP26MdJGsR3eW67xqCHN19zd64Y/Sdc/wV
r+NNbd4jBBI6qNursoN4l2BCKX1OV2gdE44Ck38Lbaqj28B8EJvuI6OEnNajLS2A
/QsK8ZRU4RikoIEeQby472q8Kk2g1oULoPN3NuxP5N4WLm+30bY6Ne+E9Bilp215
WnMnUlvM3I8T+STSkFryXdMaOkOiR7pqNnk/W70heDO7rNEKajXR6a/FBNaIU/1l
SOyL6WCMYbeFBMmzmc384bBrT+8SnNByVjGuFeZcpSSR1xMuAEAWTzy7xgjE1J19
7dCh8kc0CwjdoRaXceTb06j2zrZG2Ol1LnJnOiid0BSFikb0h8NeJ2/r2Uyvv3LZ
pVQV/jx1aKohk2qd23PVlnAnZarBCIr/Fpb+CD0uHEyTtwLbYZ3//WJGTAgKZfAb
lM1DigZb2uJK8Ng+ZiFicnqgc98boQkCnRQcEaCdoOesrCdOLZ12GX78r3OoVdCx
jJarC5TmViG2zAKlqjtMYuLYwcaypF8QRvQtVRFBu9JRe6YAGbg+MvV1+0yiKt73
4DK1YZ73sKrXgpguj4mpnyV1kI8n0JKK8m9a22v5RJnnyMRr2P4samIykZTNhT1I
hafvsV29yLiXOAdjZmsI7bvFWU4qAHiSlJDCfYkilTioe95hrfosUwqtF6CJZC6q
qC6rceQUrkqhRdv7kP8t43W8IxXFEa1NDOOj2II7RXbRyagmelh+qEABiXwjoQJ9
gnPnzGPeKHSHlVMEV3XqBaxFgku4rQAEEVL+VUCQkPuHmYcBhMrVY2ibt2pUnTEF
Z4sW6P3z8/xMaPKHnPvcKGkxC/OxLM1s5M6IvbcRdNf9KXzf88DB2DnFTUpWuWAr
KhV5Xj/acmI07GkUiog/EFjpboT7JnKa1fH8GF3FnpFIZxONuZkJBOVgniiuAt51
ZyU0cxWTe/Bce53o3yxY0G8W5I6gb7wB8hZQ8hSagiPJe8L7+bxWB7DqUTP1s95Y
mm2vSLMVaPArzr8k4RArdUfNQYQSbOTiJDwwRcPvAV2pFWGs4oPJkNb9iw4gM3Nw
coc0vvdeIHR5/CAgw5PPCFG6LoSH4TwtcgDo+2MfAgRiVztXvbuCKFremqXjNs1O
j5zTGqgDAqbGPS83qDWGZEASPiU6JC9RKVms6AShJugwISOGS5J8ML0DvKPhwIUc
v3Jln/5a49Q5luPK7ocTBqFCygbqZpO5/CdWX7T7mPeH+kM/l+jQkzb3uRkENv6a
8bWP5lR+zbgbcEzkhJIDIcMONwhKbhZjpTGpIjHI/Z7vDJ0iIZ648sStSNs9Ktw9
UJ4iDkCSf0W/1y1r7gmSzYm6FqwaEqdJ0q+Qh5dpUZaBmxk+nMEJVRjELv4EfT8q
25g0xpe8KPkDuWA0VziuiCf2XrcMmOBNbfMwhXbqTbqYrd10+tcD5BCCV4NfkKmx
Jo/oMxItN9VRD4kNC6Kpc0aReBe/mjO5vOL3J7pkzCKQdRUM9bBoFeK9oRizQDUX
WINLaSkPnPi51DVpSBED1xalqHJPhp5wWhCNu1ateFYhXJ8PGcd39BB9hBNwSF+A
7f5pKT5jyCL3hDheKdUmewcTfZrwaa56cMBLsyQ/07pb8e7d2ZtArmfiAA/whnwo
F7PLz0fP7rU4EzY0wrCP7hk9I1a/kh+Eq+pK6bw0fA6d+a0sTXM1WgxTQquwK3ib
An3miZkJouta83372srwRSAOS6KxXb6gNleZ7q+zUXVBxsGcA1BnVRNpkwRxy4qi
GZG90Udju3M4QfEFUZjdDb5HTk/ZQVTmtz/2EpzZ+s9bpBPjt4GxOmfdIDQms1SW
veUdChQztBhXB3AWuziSH8QNvO3NKYnCjPy6vQ+h7+3Xpi+CXmM1yCC/1l2/JrJc
vmfTvU4bf1fMxkZPrp0rNPcQo/yVCAnFZJslmy2lGN8uR7DbNap2cEy7zKZbzaXJ
WXkZ2wWVIgwKFSQCEhWrIgC8eZNas2k9+9qI4IqDLT5fD1FDkcHHcC/vhc3sGOCO
DxIE6XQeJkRg1kluf+KCi6rQ3FxiPyKVHuqIlWz7ZJb8DpbPP+jkEr3xWc1RtYSD
kc38ivpzxqeNwZl2uH3qKOm40N+d663i74ODCoRXh6lzZExVWJHBstrawJSQ0gRU
FTykHsBZ15Tjfc9ByvhdDxTmXyQu9zBKTJbIvCd1kjIcKr9uDss+6Z4aIuIf41nn
kVsBx1BuoHfpN+utC3vi0dWS5JM3zYm2RXNBXww0JcAbqKVmpnsP+UmaXEoFEsih
W/tWD9RpzxZfSfinyDrwUV8fzlpP5RnfMuzUYC/J6nnQLs5xxfQx/0AWEqUkw4li
cXrLYTW1I9COYogGsT1UeDcODGLcydQZqDw6DeOCsKvCKQgsedjL4Cdaef58cSqI
SkfniEhLcw/018CB5hdksV+DqNRHgGVyQA17rQGBu6DvQl2JlL0EvCpUub8sW+TN
xbFbdV+5AECsMCB013fm3N0Tmpmnn+tqOOxTfELJUOENUMUjIv5MF0a7FY+lfxd6
0i91ljgV/Aypk4dWbbZMoiNKdTLORjAMFfzJ1UN6eQbasigIsDXQSIJw3f5ICvwr
QSC3O1WfixynUfoQ9vHrikZ8/PU5bTphRYs+QuJUmFg+ZGMUY9P8HHyU7n63nqCi
xUE2ppG2MHu1Q3gZ+FzncX/pV3uzED6DyceXAK/fIalphq0RcYiobp7D5hGI+Mn3
5D87XyvuQKC1s+eoCuDi1T2woyWZnzkT/cn67P9Ek5IEJZuBVDEeq7R73mqwvoVO
SA1T2A3YIF4sjODJGtYWfnt1tZjLDsZriLcxHTiaWDDjqSK4eSW488ZJgtoYBqAd
A/djPX9zET6Jg/D/VeUmX62RAORr3isnXy6AkRSwkx+JxS72x7x1dH2TURX+RJlC
Ev3DotGkmIrm9KHA8qsE77UMroCU5pwCJc9taIr2NcexHSv99+Nff8Bq4lg/ESob
aO03dc1qN3+jBp7k5J0HEFo4MbDAlh7RkqnGvqUTBVyOxdib1NC3vg2VSDmvd8Vs
PKBRp2SH1oeFHlHQkJbx14hIcz03F8PklYbrhPmIB8k/WZWNrwspdp6gO++uHp7u
0vsFu514IKvCrXr+RMiQ9yFIkZIk8lv8yXhZP0svxxNZqxEG4G6lqrI+UNtsm2cx
3NeG36vpK0rUFPNWIqBQLBisEN1I+a5kMVfw6Iok9xqLacpEuQoTr08EC+PSi5ZO
m1k4mpCqbZbP26TSh6QouPoWIk5ATJb+lXkpILXg7+0wkLtHUe0asVAbuH27rzBK
49qbTV3eSwfEeiKnliXcqFTjYldciQfiGQHK0VfflBHp8gcT+2+ySHo7EtXiwYNl
kRGEDj39V2iHQ/fYv69LMP1o7P2gaYvmAkyLKTxhvPlvGbkTa30b6E3BAFisLKW2
eBWcjWYA4QefKUBk45EDHndCgkUq5mkjMuJ8C8KfUoMipYAgqIp8gmcN5Q0VL7Te
T/MqiFWjxD0QRKRPXg1Tc2ibhP+1yN9I1xuA3ctbLFt8Go1N3ld4v3D85aOGRo6x
Z/s5dRmdEcN57NUbEKBSvsb8nYLuDoWYaXxfNnJbRIknriEz437x4MdcAQWa8Mx6
zP0gboYPD5OQzdVyQhW6CQuf7QCRli4sB9TSxWumYBZVQPpq6iH6dAzcFmCFAvx0
JEPPnDiyJL8hQQ/c8t/XjHKsPpHlEcVW2RYWbocwQzTcNf1Upcn7y0f0hyaIg45Y
fSIbo8JpE2u5B0RIvmBwaeb6tLN/Capj/V7ZYLaWj4KG78jsR4OdoMmZGeIQZbk5
PsrrZZxFRGU1gibV26hAjS2pORgbDeitG96LTgJ6WBfGObq20euSr44TdJyURGo4
FP47Ac1aN9vItTcLTj1L9omN18Yc/7aquRCy/Pvda6g9i0zemVvBLW5IGSs43S3p
uGxu6lt6Zu75q39yQh+ZM/jDdZXCzWRdNX6qN44fG/VH/KmB+JyqOw1DBVHP/kV8
t1jZgbGIEr6dZvYYsiGPO5CNBQ6c01mjLNz3nNJqv5O0X092GX+210NQwZ+m0jpC
17E7wPl8v3Yz8VCxuKC2QqMbJkL2H5wk6xhy+HCZsCCTQOi950M+UUfyCKKlTHsT
w0rORE56EUTn/bSWN2FHp9muXCjE2rNVq+yyOlYX4U6wI1DNy0D3JtvUosxles39
Rj4/7LiOill7tmckA6qIUarT1OxSLmDYOzXEUAyVjeKOYaIqljvdC4E0QwL4mrTh
Iuh8SODwg+m9gH97NscH4venH/vJ4Go7fbywQ/LvXHyEXjmBYlqWRc5IXuYu8DF1
sEHLjZyVaJ+5jydpAsY34vsIotk7YNRFGfBCl1S4eQYtUKWsFRrpuslRC5HPALG6
uF8Hqzw6ntNDihLhR3DBgDikhZFpsg4y6tosaBCUvQWqua7o2oTS9rOVdVymLfqQ
wsnqG04PMhoOC4K2NM2jnfCHrmfXsU0eNgn5Sd4m6QgqKdHMr142LVRwilvhs8Y6
U/PxzFi7lJ+Y0Ur0N3d9Ot3culPRr9S49SKo/33RklXfHFM2wWALRuk2YnGtNkbc
1XYuw2QYU+6enAkvrsX7FpLpB1mpWpMBCwSD+DmJdHLcf+gYl+PpBY1r3SsWyPth
7i6suEf2LcJpxTQv/MpAaDN5P63ta81wm752lsI9hvEFclmdpS6aglur3ywoqk+E
MLV2cB3GWLLRVD5r6zsjrsqikddbfREZwY6jWAI29lKOzFk4snh9D8ZetmVxF9r9
3rHHplJTcU1d1mAPMXzVzHoTtRa30A+KCXiM+GYpr+RsxAvXWmv8Qr1oAnW6lfxB
8kAqJxbN6XNc7Dd4s6n/h4c61G8g9OVVkduqvgusSggGGDBkWHREgEDokZXQTps7
ju34aVJ9PsZu+MtwvKMmOnyaDwWM3WieohaMCD5yxSVP3e+4qw6wVXH8zA2nzpOq
0/u7XmUugctBXt7CIYKcO9dDLXl/SfDfNZR2JczWFnV0nEEEdijAq55/R/5U5Ft2
Z7vB+RUPH8T/gLKNtwFa9LZ4T+l73yw0SdBpRPFyjkEZ6FjZdLjyH5wz/AylrczA
UdFUuk06Qg8+Q92FI1LlMgSqozciM4cfm9zcUHbmKgqkcmv0HObYA9yNnqsoBonC
zsX6PIPEhPYVG98xR6D+spitaROljfljlGh3TlYtlmgY2wlMZ2bTR8wwEShJfKx0
A9ZVWgH81/u6D/OZxEc4JdM3F81FWxqUlCD2UbM1c5TbsZBPvxH6U2vbRK5kmZ2r
yXFbyiNZBqLYs2vvc7Xefqqef6MlkWZCpYKuny5jXFVPohuIQIrB+IPj/B7ueylV
fOYi6szzxPUkK1AoSxH7ok20CySxZfCmd6VMEZ32s4vvUhJ6tbsfHhZTnvzt5VyD
yTkz8DsfVTY3ayKiwqhueMNCSFEytJhXMVc+w93rmY06Gu8Wj+XktThyzDEUWcAb
BkATosSS7a8+bSBv7wIHCez1lv4f7+4lX4KFJLBK4ITI66wbRthhlK5QKLThNRxe
xWXJYTZ4te2qQRXN90HbOTUh+TM1OptC/0yEqixVJHuMn6QdxQykUZWfgUuVx64L
5Y9m7bmRdPCE6M2L6lUhX6ZGClygeiopwLkZVyEIu0/6I5aIlWNL7fyGS0zZxqNR
iWLuL+jfyyhLT7zZXEqjyzwGFulL1z5btHKk2NTcBhwK3vkvFYzE0dDmHsNYiUBa
D4+9MGm9udehjfJ+kxRyeBZOug0LDBlTwqsFAPpux3Rp+kAlksPnPf+/BZZvfHi2
GtsHab8/2dmHk3PGpsD3TPBj0W6AaFU4ie81SiODCf+DvweVaPR4DJGI1bBCdom0
UVlZgc0G4zOtamllgOn+t2uA9w7XBFv+wxQQL6RFpatUMWuUJ2advgVY7qBD0nV7
JMasYg2MPdqb4svqKETD1coGZblPI8/bbZe+oRdQUAu3cCDCjQlR1Y+nHwyOlRwf
f0OwzSThDToNjQsNmwl9eq0rEHOeDfH1utF8m6L7YRUPiWpoPhyq5XFTPJ2C9Yyj
wXCnrD00yZq5+yTE2w9Q3uoAyXpRDJRai9N5ZA53GKvIQEhOuQvdEA/kWaz6SoyP
8tyscK+5Csb0mg62jO5zl2QW9vXx6GLRDlM2G41QAdmmBQP/Vj2xwpjQ3vqW6IKA
NJGpEz12v4R/hjAit3wBMS+jDKoa/hGsPswLn0MU2TIo6FjBdROKVP8C/BZnM/+/
RNiPCS6lcECp4hFQHLPB7n+lLoI+XVN2OariQumZRXDzQFl7BchNaDTRdjhPCDh2
kc81gsO1vpwhR4f0j/1XjkVDomrDkaYLl3IHNA28t+TzaCbrcuu+32SVejFmhvJW
qeWkG17YX5jPmqHEMCCOR82+ctKQSaReFBFbPlEVuaZTA359Ztq4uMfEXiXK9ZFj
NuCSijIc3blfhxFl7dI2mUVrnYPJwwKYwuNphT8ZBMK2OfR3AAc6ntwDMya4ueux
7M0ekHPz5AfecsHX7foFeIpbwG/KZDAc0MPyjvuAuSgbhth4ZJmd9D0gBp0175B7
q2jWJBTadBRwiLNXFpcZeJ3ZC4/VybHAaXrNWR5LJ0cXuVBz4A7BdJMmSMshTSIV
gEd3quVoGslsaEa2p2EdTeEKeQwP7IAA9ewwRTGflZF9KL85kaxwqNR/XW47jn8Y
SCwrvdlGluULXbC5jvbzpwHtft+wC8LbD2Rv5cKp78YpuapfzwxGYeiC+Z/gPysJ
EGFkeYP1InI9pJ+6QOWMMNyMCw8cMuzjp6hsgWxauEp+NjtMWBKStALQYmC9CZ0k
MlQsXaaZVvOJ0xJtqyWVnxAI1wdgarP4N6GIbiM8yqGFjy8a8nujXVwttrvVZgan
jd2X7QBSL4mTE2p4OexSPFKoegyv7Z+pW+FTfE9ieGOHYiVtbygBR0oFaFezEhhm
jBPmzx0fTgxlhbxf55jQQ2eI6e9YHtKaxvsLK9wr262fy9qbqBy2lnd6n1pYMD29
I0CRflGeV7Ti39kR79Ovmkat3qCEatNqQav/RHoQ5uVOPxG2MaTG4LEWUz+SWI0F
86eVH6ldR/8ZhjWL0Z3QoSz/u0/y9l9tuc08ARZ/5NmjRKrHuNX178sfDlNxxHlw
qgJeaAFwrtLl+9BhNblg6zrP/nQGFsXaF7NGIfHEKx3RrecO6hgFUkYcY927d412
yrK9YPKEkQ9l2cnJ+GGCRkepeyyvDW8yjQC4QVk8dQEZj8YetF35oySCpN82EmWP
huIVEf2VWnTmPoLN7AD7tmXibHEjgC3kl4xm4o0WJ0/x/mJUy85qGdbMjXwjMo4+
DaI1x2f99M/Lgzz0T22PXlH2CknrqlK25QbAGdUuJxBtsP7SyV0sEE83S8exi0nh
lJT24TaVfa5BPGmtsP5ZcfH2otNsGLYHHRtbGhm2aLhGkGtyLBCxjHkj6AqhQC5C
AJqFPTFEz8fLGrW8RbJjCmBY+NfqPWpMfDgiZ0gO81RJs4+MY2FepVib9oW4l8N6
rUZDrOquK8D/oeS3RCL9hu12L0cyiG41COYwPsxKew4xCZwpvVzDnteE+irKjPDI
qtul9EG3XVXGzyEqELo51FDyWhlUm98pxbmWtU0ysxI+WmAgk2d3P5WRn/SciVWH
rAf4uoeb0rsyWVfuK/wEnB4tQIwosRwqujA3Yf/pRoBceb5fQ//esB/Zx39AoKjj
JfO/Bdh6Om9IOKm+ByiNQhMhCEsy6TsQKrc0KrQx7JIEzE4U0knGetWjyU22N+hA
0xDjeK8Fr2hHiiS1/A782hb7ZAeJ7v34SSh3MOW3fWKZEI01Tt49b9HKHphiC/UE
s16xBwPASJtx5sV9IGYA6daiYeBF4Y+vfeGTh//LpwTJq1HvEvg8AkwnceGAwHNB
QKisLdQHIROnZuc9cKwQ42mI7hVMD5brhizMrPebF147T/0aR0tCf3Fd3Rg/ARN/
C0QzXkz4gqTLKxF6L6phRVwrMlYrkSXbnJfSfJbBE8wiJm+0DtXQvlSNjc5CEDRl
34z1gvCs1SR5fnYGHOcQsBWzQLlivtA6lrjbNs6CLfYuzuGSGuZ0yQMmh1Sz5b4I
WvMyKxD9DXdRzvSmP1ecOnMXX5zfuoBYDyqB1fRup0KDSCyh0Bjdge1w6aRipD+p
ze5dALL9toEswUpi7h7X0Qeycbpmeq3nalxxf+jN+zm418mjgqtObusQTDR+ytxB
1Yl5kMUkfnlyWZbXajIYn38NlcXGD7gzvQreqeC73cpCoxUi3TqYeVE4WsBLF33c
V4V2MH0M97gY/zbMvUaNWycGflKZHGcfWB8OR9HZu2lwUVNnz7uXCLuCIp2Xl1Ls
fwHCtYdQv2JR8LpaQmQchsiS/Ou2MDvEHZJDYfu5EoUrFh68XNEsWR96T3MYAoTj
l/wBb3lCzgGlwxQpz753W41pQVeq6OuC2OjWxp4H/rjusjqomohuCAJrYcaU/SP9
o5weuVTk9QK5rkUOysObZU2UtDyMo8pTx9CNOwavP5JaKWKBGtsw9gnGXByG6Dnq
18iR7e6l9/Z2jwBR8e22OPnLubmViOB6jwoZ98fWADOqPlZ05mpEajEyFRpauqlF
4KRYREPayrd1pGyoDTjKxTMeFOz2jXMJXFQqiqGfiVBW91/pIIMBuu7QKP+FMzUl
OGlVSz97EFURZCsWjmeUOJHJU8w1Gfpxs65Nz1kX90i5YodUyaFHnfJQQdV7rGxA
sqFcx8wN39gXAwazFdhlD5+UStFZI+THpf9JtThdSNAsBtYBToWSp4e12ViZKVf9
fTJqBB2sO4Kfvq25s8TP3YQ0fz3iUiQHuOzBbxwImT1Vq4mu96dKgOQ0wJcV2r5h
CjGhIIE0uSY6jm0T1atqqNY05Gz3yYjc50xPwcFhBaJ4loNHP2jeZJvIUl/PwxmL
qlQNtHc0Q1rw99fROyENu+1vHHNwM1nWqki+H9Lx+atJqH+FkmL8SRkD14abFbU7
TmOKB9C8gGXM4hSeuVXoen5JDxRCcHJQIoshP9vM7eEHelAcmnn7mgpmBBOX8JLC
R+Nedj2kbiFFjv08MKuPQSiCkYWYliE8ofkhSQ5wfiGjEIyZfPsFkeQF5VQX9AFf
Nriq9gKjlLK4c0T9AJ6rr5pntlLzsIq928LhjArEu88pNtw0R8DhKo4cdSFqAnZW
RHGLuMnsAG4deoeP0wLGPdBsQLPYEQZvMyC6rYhC7dSSImMacf6U/XcUeyKnPgFK
mdr1XoDY43avh9hX5RsyrTcrOtYWCGkS40gW0IfQMp8v8LxsyzBFL/ybb5Swj28B
r/vSCus/zfe0bA+u5hiaELL80IlYIF6uxV9M6Whh4Ms2xNnSyHWd8MjAA2I4227B
jnh6ocz0t4ju7IN6LO5lsyB5QXt5BVDrL4U+JrU+l5/eXihjASrCrRgzmgoJFBAb
CpMOgBabPYSnZJKuH4OX7y6ijdz3HXqGcv6KjDtdID5MHFWqL7Gb9Y++QwypGsFF
NRMABnvSm4xmT7qcDJ+jNUBZfnmsXh05ijnGgGT1pyg7/STC1nO52QxBGIzrKtCJ
QhRSh8ecepRTCXS5rImLc1iMXWnvzbArtuSx+yLqzTUEbPIJ6+PpP8/y8uIsh69Q
UHf3fX4HicYFgcXQEN2XffkVJ6rbDiHRb0gaHaruTcZif5w0jmkImikm1wR8Vacl
hGRnRPvpv63bdVo8oeiell4B06+IHpj7jLqjnWIer03AVr/Co/ff6dnQ43WBTTTZ
W+D/zdr/wqjbsLc+gNWDjrGRXFy96+sxGpA43fgTeZYJdnz+W/9YLFZyNkFdhchL
156cYy71XPGRGVt7dz491+YOUFfTNwBfYTjuI77rghcQbJ//IiPZMEJla4oKZTgC
t/OJXpkKj0CjwUS4U2N3hD1vkMzj5Hz+1xwVdACOGJj4Gte6f19WCghdUdfa6lvk
COiGD4CZzTV5JuFrHpfn6dWWUIDx3nWGuIdb3kKlXBBumohYJzLTeBzOv1y5xpjr
l+i3pfJ1+rudlBPRVT0BVK502Dwwu6DxT0gZPE/+JxFnD8pDu+GAgBNrnkZGio2o
1vbq9y2Z9yGX958ZmJO6yJAClV+peuyBxkYlIj6eb2wnodklnAD+wpRybqEbMdyK
tJHuckpAre8HG73Hcp4NUqo+wJ+uYGJTXgq4ol6YgoQRDqDoBxr0xLwy8UzjVaSN
dtM5OWxtcFvucKVC3Ba+l0Qxe2201TAIQTOQRyG3RDrpOvEB1zDyRQps7sKFhP+b
Ho57ZDvQx8toOKTCNtfNeaoPEqyoHrleq4Xhi8Z9h8ILIvEtVOd6zhqtZ41gmPUm
EwqpoX8JwDyY5fBXFNandmQr+ExS73QNF1A6UESHlR1E8VMmSrzVwJ0/aBLu6r1l
tf42LuftdV+5qsNEPWCijjf9katAvIH5wsvQDO2ffVddFkAkyLU3vJCakjdSx0XR
GGp8BZVXr9raugh2U8lVfMy+MZ2YqLYQJedIP//iPkyiYAT5jPIqsZNiaqmpD8fE
dCmfGeepBfH8+1sgv8s/STYzwINvrlvIYfcxr93NirkMOY26yzU+hPc2Zz5O2loy
5CDnZX2GW6Whm4wMe7je44QTn3hOF+hhYAe3xsS47+khjKpdVgvlAiP8ryEFitJZ
42L8ttmPUhC599CLyJMgvzHGolaw2N8qJZf/+5gpIWHucsOn0vdKoNCki75jH5tw
8W4jnkPnDFeL2F4Bw4bj9zE2ihn1efsq39XJWF901mvpoMYBZFCOQfIlk+2XDuyM
z/lna202DOU17faqU7ABOoI0yqY2qTAtgkXb7CbsdMgHe1Y2UuE032WYBhH0nNZI
3HcNvKinG8z9Fby6ulcny4tQn9ev05k9GkGmWdnR+BO8pUq0bxhdY8vlw8A/hGaD
uSZkGwIU3xgLmfknI+RlnxFRsppAwRkJmmxnaCssUzJR/xNcmclC5Tt7oFDo83Gz
k/ye6uUzF+8b8PSrLNF9cMK5UrMpoPUa22c11/nKCbJULmimO6MLvaA/iA80cTeq
nQjqHcmi14U7F/1bfOFMJ5DNCvSRsxPkNt/8ITRrO1fHvCTi7G6qVjKD210PHXHy
MeemuidTcSvjZ5O5Ut1iIwjfiJtPyreEOSbeeCxx9tnl1C33xP9UwkO9KQeL+NI/
DblLyjNJL2qygs2sUZbS7rJ6biGVkTh+Tsi8Mejv0r6slEv3gYtVqHo9uJb10fWB
Z4g04P7skLavDC6o09ylBOtbZASU9wu/37w9GleN8addXk+OZemKM8IbpyLa4qzj
V/63LZvVAVPO3THN88psu9LyYXnv2C1zTVPQb7x8lQaqyBBu259iEW8VmSstHcHA
cA/cGicSf+oxeJbuCj9ulfYt0rkd3WtOfkSLdwsAyFiAHRipqczszf43Mqb5pYe3
TqXSJTU7xZwWImDjp6/+mWyby10Vdoii7vwtWfTV+ZNRxssKLx+Vg+dULq1YNzKB
8GralLbxsrYisgtK01bP0R9LoP3zlXw/Whk7x+qJB6Ri+s7Y3OW2Vlu3wZi8312s
zLjVG1jJTd1gv5XId4g/8mEW77KfOo3sNQ1nmFwnH+6/zmazH7kjG30HTNeivlrR
rQjH0NDmaqQcN71hqD67TyKMBcNKyxYLIq/OW/E2vrNK7zpDtPKc1VenGaDemT7l
FBFCHtP0R+SNEuYXT4m5w9bE+wtlUYPwBVELqOK3FfLXCGJB/6/kJ5ynBW4YVF1n
YRouM15iFY9ObfBz85MSuVyTKwGnfg7sjU74qe2hMpJVgbz3rXBlDNuT83gaDIiu
2ev4hxjiad+WcBEjXi/2QoXfNKhkxi/dt6LcRyxTwXYEeTQmdeDBH41CoHZKij5n
e0IeW+vf2A6qinuKJKSRxpuH/zl8zgIfyN14NhJqpcMvjElfYMfqPdPLpRz4+Vod
VZ/rsEFqQnCXUQlqatMQj65SuSNCT5AZGWDInfJlY7kt4CuDl/gK10g4bZLVNpAJ
cQv4fO9h4GhoW6j9M0hBS3UE720iGnR3oDIliC+qGe8IC6AblbDOKzYI+8YCyVvn
ZljMAEMurcl4f35MwAYUVTxlc4rAA4H5v9k/H38kJUiXG3xDhj/aB9+bk8IlIiXr
71Zu1PobAXNk4FMS72KE+X5g9+PpvgxPyp1NXptCPlnwKXRi85/XVYOY9kXQjTKm
Eb7xxosQs9SDkML5lgN57Zgrx6qP8qohy4zY9QnV/ctYtp1ag/XFlB+RzDJhwjvw
yE4aTdWej/2WwxFXSc/akIva4ulRjbv/Ovg5Qgig93k/fw5wR8c0eD/BNF4UaTOG
wnRv2dK005rZSBLobT+UBGHz3Xqz1ZbQkgspVgvZ8Q+/J64qbUnhhuin90IffzMn
BUmy1L/Hyym+mKXvyvwsU3SUWfqaqG1lKXkRiBaX3A3pUS93Xzwz4tk3uMaSkJiW
dADaftLc1cT1lSLXU5/ZymgRCCCaiK+0mg6lGZ6faeCg3irRgFA8+sL7M2ys0bMM
p+1pb1aF1C9hirN4ZPqLG60PjdpgbK0oo93O2HugvUO/iv8n5gz05rgRrm2DBLeN
sNZH7Yw+NJ9CGjvJYuc1o4m75XyIQNWqD1sGquzkiySjQXmwNq032jdLXyvs8+7/
V4aEV2tRsSmK/a5nBgqRgIMiLEAR6GTxYVX72Q24QZo9A3zHB2qlaO9A8h6Cnw/O
RyrbAuYBfw5lNPj6SY/HWzLb1WjuZ2d5EAhcL2tSeVoVWbKuBPza+WWTnvN5S/Un
C/tKtsoSpScD39NmWR7QW/hegJkTJYymcuUi9O1KRu+6i/d1hnofIx1EIEUSBmkg
Y/0Ad8FmAhejw813m2tn/6zA/ot+QbjF/eqvBz6UXMYTrWyxQcHFKqH2T3RCITJD
ZsjkbPFHKtImoFBJgHDLM2xNUa++8wMON5b8TcEqOyMKWR4xgw/HOahxFfCzQHpw
sOqKtcOWO/+FbBOzG+K7AeHOaE0HZFvd8B7z5u33dgWrQavzHSOoWm6EKWmI/ZaF
LSidKcbfm4ouMakOiAIQGS0AHl5ckp8iE485e2LDJ3wcfCdG6PQl2pnJwrYmtY/B
v020VSK5g7axKr4lhhVPvU0S56eHCWdF5sIbxVa2SS9s5euDlJ/tzlqcPjrQ8duw
W5A4kZkgAgTn93whHkkvaUD8+tXiIzboB3WSY0UAsdMM/1lWMNk0HR1MK8Ja5dCs
usv/Tn6Qg3uJCDodfzse9H5KBTQLe5C0FfJmHHHmYvjruHax37l/DoXQ7SLlGZoJ
1U/AYVoT72WRimK0rkh7iOBg2e5tgfpvHldwFAqS0s4cfGWdi3Hkwy1NkdHPwSef
V0/VqIkL266yHEowu4do5/b1nx5y4Uiu7aK1VpFSRCdhQCZtZPDhP7ifCyFwxrd3
IvIsvoY9RrTVcbmD+om0PYOZH/VY0UlTbLAQCSNEH7N6OyWbDCv40LSOYwy21mOW
jcF9S6GiIW7UiI1T7Ku9yJckCHNi7T+Cyzu9MY7XZVtbNwY+VuC52l9Bc3Y8zwHE
r19fK9P9evaSMNx4NG/8k/63NeJQGQWSwpBGB0gC2Z43fhnSA5ewDAVktVUibFt/
wujiFVAmkb5Rby4giLa7H8KbmwXSumaYck2wh/rOWnI8tR39nPOQ9WiDMXhfer9n
R7Uh229AwVpIf7PlESLht0q2RS6YqFABOoSoiY3bE4rZVp3b/RjNwdAVW0aN3ZlE
uSNS6CpWDtCk/7m64MFKACKG0iKVtr1GMCF6P39zuRcDFKRulwtEvq7Ne9gg21S+
SyN7mIpO+BV1pYX99MgYGd2xbcuE2U2ftgYmnCgN24BhR/BQGF5cEvTNZqcRJvKv
UMeTtWA2BhB6MIE7oUe9cizr0/bGp+5alWI4u2aFcsmzE6FT06FTFGKDv5DagiX7
/SsSI7zk7sGpNpsA9EUYdoSIGu33cqIQDb06w+fTi0iNoTeWNlBh+mpCrmaCvlIq
IKwDCkfDOUc7SRNHxrGYfQh6OYnkxk/dnqX9PHedAptz/Erw8Ja3e2v4IIgtjGLr
wArNiSBuLBvGhGzKufrimuDh6OFqXLRYJw9e9zL4tBjNFRli7jsYnS4Mumu+tdCw
qh7kdcdUgqZtPiGZ/+YEa7b+HeJFCQ3DZtsVannd0OogY92+FNxVLQi3U9XQJe7g
62uERcQzivtEfNsSswW2/IYx4VgcMkyIFshmflr1XdH7g91JnZJuJt1E+ui6yyjt
fo5mA7jsb6KVzquDAoZeeuTnMRJ3imrgo+YzDjwJv4GHKaPeSeOES3lvwNCg38Z7
q3kh7G42Z6FZ3SYwhrL1RScRX/Rc7cBxgnRAgMfMcwGMK9r02ns77JdQDJgRgjiW
StcgTsk0BzlVNRrOR4OTX/j8Zf5wEn1Up+bQcFbcKXN9CbmDhYJ2c/HODOhBAJTI
xHdrJBzvYQef5/tVNQQULd008QTKOqACHqYSq8LhqoikbCar3epI9Fe76pQGh+fF
xcuimSIrfgKplebFBEyruOBtaicIa26Zmo9MGsXAJldlRruA7IipVqCQ86Szzw8a
My/FLyrGtpWucIlWZReoFeSYinRK42f4eXPBCol80RnZGw6ybmmzaFerUJDxSAEY
EA94QFTXF0ccAql5fTIlKffHjktyXi0JeE1tTSUJ7rz+3wzP7IIqG00uQWWiq5zI
IE28aMB9mldWaT1OU0gL97pRyH3LzEKAQ/5hbMdTwDwfbairrQXaDgNY8VfhKGnL
UH77Lqub/jt/b3oVQrd51uw+ApNgDuE3n2J/RXf5DrBmnBf4x437rwSt4Np297qO
HrnOLfi4uZMCpC4XV2apw4EGqvrgZbUb3l4dzcrxHuGAif//QDamRmhM8BzYeEwB
Le3RQ64+/MtzgvsZdUSfNxjmmhm5vIlTEOUqea4pfm7cF8ol+x/Er2Uuz4L48RwH
QCNUPUOqzbbOjvXRG7WVveBTKlDt/rpb5WK0iUnnNVCKNua06Ud3xxt+DWXlCyFL
7BPwspMUSMwZyEY0puShCgaHDphqEkdZtKv1erW4x9M8qkU1e8IH/pwQ0APYmooQ
4cdK3DCOy+N8IEuwRCq5s8UMIVkaGqmC6IwSG3S0tWuaE3pTeL/maygkor4x98Iz
sC13DbXxtez1ce0OVU5PtGbw3Ka/bduhSf2fKkNsQj+6QrQ/wHKo21+ZkMt7TY1Q
lBKNnjUGTqIZkk+OYH2eBb5NmQP1mjuBjXCvRcY/vEBbKiu71W0DUD2Oxe91TVOA
DpWoLQJNfe0WTnJX8qPaAFmUjSnT0rFb8S0B/1w7W7TSWZ8yYjgysAXQUPOGfbOO
a5mASMvViNW7PWnH73+wp9xBWmqB5bhjtOxu/mKXqZIEy2KxuRdgrtGNHZnAYyAo
NYYJURW/WGkmRCR+T1CaQCUERQvyym0oAitSAsQ4bVpTXFSaKeuGf1Z9P7x1T+BX
kxU1lBfayXURQK6lgArLqv+FUlKd61oUFbv194uwCZP9Te5J48PW4wlCxLMsik70
8iYDFwXC0Y//b5DUXTbpyInk8forUo8xTbsf/hpNEBh8pSU23ifmCmveM/Iyk7Rp
8ASUTFzUU54lxXjbHluWIC4Ndc/IPrf7qCI8kD4llYX4+Tk5gbBHoBZzSPDM6rg+
w86QfIb1BN6gyZgDzHcu6vp+z52Ij7KHbUw9kZBJ3SFsSdGS3shSMB3QyhEQZXtN
z9ATrzWlp2fZvaCPWaUp1XoLTIczVsaXIIGHLJudJbLs6XZZGNTIV1erpWOaobJz
wrCNQaf8eeYDnpeHHPDqU7wCa6w809b65PAV7lz8YyDUEdLVWukSbKRQgH1vzeao
6lVghke8IVKnKU4SsERPmnOIOHLNy7KBk+VVJED+COtSzsaiqrUm0yFdy7iZNZ1V
RKjSSYEWXP9p575imUcZVGQOjYkU2fsAyr+JkmzREpb7/2fpTqbrOJITLoyGY8/k
gbvXXLuTJvG1WkW9pfSFfqCn6wozRXn+lps/3ZLgJd4dY/g7Kr8onbBZcDUBHtMN
9ac8i0kMgRjRgSK7ZNHUyik0DWWgcj6Ktq0pfwuDqABTylXLVqlnMQUIQ/AGcLz4
WatiWZme1BblN65n6N7wi2LkdZvVwdBiXCmutLgidHRd2Ydkk1RZcqD/LtzF4KsG
IC4oBO7Yl3dS6LRRWpvsWhb5QmIsR6FMeEt7/5yfUBTW4JgTLa4pMF/jfstV03LZ
IZimpAF9VulbsN0Acto6iotcVd8/eSUyD8ucFoSfZQCu3mxHl7hFRpQMe+aPzzZk
t+H01un3RWaILkjaD1q42ohXBAB2clK1Wbj8Nmf5PuM4iVOLvoYa5/rV8apD+ifZ
qTK4DOYg1bDbD/FQY0c1ohDzEF9mljh0TggjBDh9mmt1W8Y1jWhg0j522Hfn5k6r
lb8xZDRLQZQRNFldzoKHu9F80ZQ4/mXBhCLRgNrESr8L9Dy/VQ0jXQ37f88X2Ipk
2SXV19fPcl3xt310DyL/SAU2dREe6RW2U0YDBqyJrAXrD2WBMMfT2vnyJOEJr6EB
1jVoDg3rrDPzM9TWecdurzxHY9f0/KOXHb9AipM+s/GcFqdMSjDIImgO8R+JezUr
9+sg+XvN8WJsGH6Me0wA7utWjvceUmv19CfxY05gxXXTXzAj4ZC2cJqzzhNEx5Nu
23/lSQZPqUepF42Xt5oxaUYzgDoOS8cV/LQ40ptyzs7p2emJbH7fKpYxD7hYb6to
+sbQ40Btsy6sXh84MP+pLYOrFsoewNS9csorxIY67mdyAo3SYpFSNP5wLnc1VuQ+
vUsmXQNo9tr3xruOc1pKOkyvi1ltZzkClD4gyTNaCStZS7WYcRq5cNPG9Q4lkOh9
3N2RFuizZBOASBOUZyiY7kPXSzPhe8frIRw2HcjPpOgT32WrGZmb4gJnYxxbDYvM
WoWdDZOQJxUrpwn7te2bCMdnBbpxH0UKCMqeXi310qM/MoC+UFK15Fdimi9MOkZY
ZjHDSo4wY1GCF/o50MQtzdVPr3rxTSB+MUvrHG4BxiOTaVgOYuebqvyqR1Dnkuuw
tTBWSvEaKE7MiBFUEVnAiA+CG+e+IbQkAwWzVeInygIvB7aBfS0Inc/HgHpehspF
UC7Y2FDNXQOjW7GwHY2RFk+AW6y3DbRisn8NYY13UBejU6r4W5aRMDHc2fzg/+QI
UWS1AtCrB31bAyUVzgBz3KHpKXNKyvvDsCdQ62DMm6fcrtFGSPMBAMqknmMZCV1z
cObrozhQA+/fGTaUEXrgafrkSPQT5HMTG8Yli8q65jvRkXPlbbIbRsbdDBR/lAWo
nJlBxNAlLu7TF1yjqManryOJgX5HIulUGSjIwzS6fgaWW3JpQo84o3v06o7y/zsD
StApa3VdXxI2ZTyy78ANJ9tM6buzkErJp6uSau/WMnREiRuzJ1UXSJYwC2FQoHg+
gojY6aYcPas/Du92+3slkNyeZTQLIxtDvDvgIX/53HDFb/CupJPnwMxlso7DNd40
A8LE+uhJssq/Gt+wrMTEMtBZAsA8krVSFXdlIZiA4EC3nqPBk8hwXv1fPBee9iOn
+vrr7OeNJvS4Jrtpv19Pke4j9ACuBoyR6gHAOTpdCpZf8X4GZzXuLLQA6HdF6D1s
hxCwCd8Gngt6j96i/MZY8COirC51q3pR1/kVHa6NOwNtyKBLMHF6Fr97rcRJQugk
NHPvVfcJmlUnS4lPiXO+ZRF1jizk2go+A8kpaKLlmbFNMvYXbRnlqT4uIh0gCZUH
9ksnbifNBNWUs3JhrByku09CWtR+fTMtGeBsg9SmpMJr0WFUL9QQ+TdrjupANZye
FC5MW8P6+nuzLUP9oB2VPdyeoweJKESuRTcDgfp1gp1qBt3arjjER6QSPLUlmJ01
xWb8OboOYtTLrjVlmAVXg2GtIPQNvjIffhoygH86TNpVqGXeMNRu2pqKuY7gcj2R
784iTN0fkbSK63/7at2a1lg5dYgGw8SlE2yxAQLoIJ8kkkplSTCwT3ydVj3sZUDo
bIjgBQFPer6MSKUmWU1pkhHq7GlGPedIGyNh2Hwx8yUZiyD6Ly6RWCjkqbz2a+G2
53Xa+0uQ6U1M1xwNydRL5HhJGtzx5CKVN8t3YLYiAoWiPISBu8qvToK4UcEkuPot
6cA8gI++yafxBiZ+7VvDm87VX/y1E72aM5Qd+3hSuSgv4uqPtqF4+fNkDmU30jSH
iLNJ7Fcuf6f/q3CUAtoFLvmuM/en0+yOQ62J1SxgXYkfzp3YMl7jHlxkvTiYAQ3v
Po5lc2/3sUGSpYS95xJj5+5lb7YWxoYGkq7HC6wtMmhUU/3K2HYIjRSdCNvWSIBd
FcPPTn96yiBWhq218SWuiBRlp4yxRDKOgyRQIZhAqUUOutLWg10ZAgXEmHPhbhz1
9BfjxS4TovAGuELuFnEBmZDOLplU2JfD+KH9b0Zv4GvynEGfGsiTN21oIDnr8wIE
ELgjN7ayh1o7D3p29Woofzc8JtFNQwze3WyAaUCNYYiX9FaJKxpfr8CKKQsAbLUm
4MNjhoa98i7/uPO39+3SK2yELoPFsCG0k+LNv0bv1q/Fy2YVSHMXModsdjBuQGZb
PXL+mySnWMoF/si8IyCF4XxkP8isPEuBC5mDUpEPyaac9e+UJFZp8tnc6Kqd7kuI
mkMLc3/LmsVqe6QAduHh5K3Wgysa77ZbijXSboCUvRLSZDmdrINmzJ9JgvJwDpkt
XNmsqSZgL9gP3ZrPLHVl1gARVKKTdFiY5zg+MltxnXgXYoyv3mxjXyzEvQA2Yy7h
fx9tOXkwZo4XTaFknnxNq0Zf1NzfMDk+bWz6DCxw40L8RAG8hNM6m0Hr1OwtT5io
oREfPuPjN4HMy4iykkajdIuQK6xvDm0+wOE52AOAxauJrzu42cI8+e1qxqp/LFin
C8KkcJ39Ztq0WVYJEyxgqP/ChZZEiAjw8A8M7enAKF52aRn/UVaDzyZY1Tl94Gj1
LG6x7O1mHjAd5fcKCuqpSSc1k8hkOEYb968HUcYuQqWmAK65x84JiM/62PnSVxrA
E9y1K9zZoXO48Q5OZ1ljhJri5MynwoZlcLP4IUry7PQkRfmytf9sqe9+dF86r49C
scdJeR7zZ9V9euVcOvtnIdSCf8U6ar4sYKO4OkszivhzPNQJyZYqK1OcXjWTOK6t
emOFZMOm3cwTG6iNLhgbFECH1xw359UgQD59N9tIwpvjPgcZYPfiAqKGbY97pDWZ
5rnoBOwiPY3npt+ntyoIX5TanqZMwxa9MF5vR4G7xdTG+vUo1yb+8pIo/kzobe9j
LBL+0286j+6azUTObVfgNeul7M4I6vnqzqf+xBzfzQh8Xm0YZzCKZyAl00ce2Sm7
LAjWj3A+ZODM3cYCnNGcOg/W0aOmytSiPW/Ry9ZQwypFdl/qXwwiCmlccemWbXn7
d1S+tqmWw7Od/M8ZOQQq+bPB04Xp9402CQcEKGkTMGWFQcQl/eNzW0nu8LFETvWR
oMwNDh2jEn0awgPjCubkP716YFVqLsPaCQnz1L4aE7fRh73jZ1inlBJ3y5h1xf1T
0GhHNP1t9vkocRi+IOWy/kXSmbtZGfxCaSkP9i3W9B8sc+JLxZWnxAhzrypliHSK
0YSmaJT+dVQWOn4175VXn4PboEPycEfYaEuOXXUC+IsFalw/+R1IoWEQeE+wc6NO
K5RYBEeeYdREXsMjg1Grx6aiBwFtD0f36YE2+bNYqjp2V6KJ/HmNIXopYXHsIeI6
aJhEh0k70LjbffvQbsakJwjgwCu/jBxE7N6mmkl2VokFnVkqY2W2d9RxnPm4K/6+
GKuHhhtrYZx2hZGBXNCIVZctavunTW3keAmT0KF1ZtpbnEtSMo1ZjN5j2dnJh6R3
GOBfhbTipa3vCOuR9o27DKdO4zF6KhpATArinsl06aMVmTbUqhPiokwOkRhR5ox1
hR7+zM57VzP1jqrY6jALWpAXeY+kJFmtzU3npghEHba3qs8p3hi7Q3FMxZsaX1W2
MMATGG3B7JIfOuKgKn3b9EAUWADADSciLCalFo8tBMdVojiJy6Br89RTiNVzZXaY
cnKl0PG5Jdz8bwDCyGsRLXlvs1cBq2ABr/lLnVC8wn3ay58tNv7bsVaOxdmWnoCC
Hc9vzaZSCPZG2N1FcnqWyhwqYWKCPNcjIW8ugSzaFCEIKD7wEmNy49Z0/5+BdH6z
DFlHKltXyW+fthNeWayolt7/bF7gevD0hZK3HZDI5Ft42Jkn7wnpH7nKFT/+PN8i
nlkQt8R/tM66xni15T77rgIyxndFzDj1TYCu2R44y5jebKEVnUQBSQZhqPkyvWmC
znB2V8fX1id93w9fi1tnKIdy5lPhh2sovOGLcwKoD+sFCZ8t/k13NcOeL8CRlMLi
1sxNaaHGipzU5Ge9IEexoAlfieEvb3fUL1+8s3U0ljFFmTedmlDNQIrLhNFn1DKJ
ObdTPlhNoHqZPqKOM3PBqWmNxy4qfrgcv3t/wlfTADGgNgx70fBjEVGpjntvx2TJ
nkE0EGrsUD7cR9sPqKJIF70X/mr/2KsP0qp+NqrQFZchAE3JV4YKzAwt/QjDjH9r
1pW8DiCVkpk4/Yvam9SEk4qInlFFp4xpLtsijyPLW7Tk1wlF6XyLM8tj8R5faO2P
R1TJEZwVhDuJ29J1g4j76jno9Ji/T4ocr3Tw3KPpBcAQZUDIG2gaoUcHAXT7f7GA
6gP1ZbpLh2z+5RXqS+klfP8Bx+La6m0Q8TO2NlFv8lT/QHPFAEYw/fU+FCYK7eML
ED+VDzJGCpV9uNomcXuY1GQgPxYno8HswwIwCjRGzS58c00Wkek0rmDAGr0lAVPp
QolHcSKUAIYWDjFNUgtW+eh7mOOH2x+yrAh9Q6yHpHSvn8TxR+3/KR5qP4L+zykI
0oiUjWJciMYvFQUc6HhFeKNhvgMV1F3LSxAuRN/dJRZorXpWK/a6eizXCa+OHDCW
J4oXE7+ldrMJM8L02ynfKvdMwkcp4miKN9JVq0RJRRuj8i7ghuQKF+fMziv+J0q7
C8V6B9Llu6ozUhz3LYc8wMh/5QUSxx1n0gtSE7TcAweOYaoC9J6u6lYMpZSdmd7V
kJt/uEn9FaqyqDtFSsebWDCWy+umThXh4DncxclpbejnzMDyFI1LD9AxuzaGYSmj
19T3POvVjZmu1Gdsqnqn0dkufE+ApNnXW5RFPqrswYYho5jjSg2PquA77UhRjKHr
/jrNCnvvz4FVPJTG1CDF0Bgd1S+YOXTPyyCNAt++rBBxkHgTB84NmtAwnuSgOEXI
eB0GOpPDpP5pVrpbfNM8ib/ss8/EAFmu8J3wehRVsjyUImiwv8oCW71PDWsiPEyR
8wb3zSGt43NgL4ZQXkd0ykoXoHivt56vqSdzmgXvlZxFNwWh3L1QeZTIFDeoaTGi
5rE37H7/J3RgQw4b5HH4zbxeHUvdNqrjERF8vLBkl0KAmBfSeMmyDEj+FG/jnM2W
IjtkcYoPggpL/dP/9goR91NKMn/Jm/Px/K3ukY7YAEr73UsnDbwt0kXRBlTd2fam
n8tOVKol4zuccXHYULQFSbJEsBWZfJ4mAx7w8StA0ghpBWJ6+udb2ybBjcmI7JpD
UFh+sQPiy3wsrKScu+fw5qn1asor+g+Ep8FRZrum7j9cweY9Xkf4gvDNDYjnPEvr
ide86JYDXYpGhWff6xxSmmBKAwC6Bx//zgStLn2gtSJknMqpEpe3ZBGiAcjM0KfV
pwCewBtGp6VdDgveXnbXmTFKFxa9hM2yiTQfZ6e4lIf6Lv5n1guyTQUP86fNs52G
h1m3onbo5R+Prr14GlY9iHqVRKMgB8/5AUJupgMgkuvPZUouLd+k1LEw7SMsB+ZQ
FfwHR/bHoGh1JhCh+zJ5KllnORCktf8gCFILgo3W1Z7uiIpw8q24+uRMgn5UIfMd
ASvOOG9ULzfI08zb3wR2k/oVPZZEXbySzcKcy5+JB2IaPsSNoVjDGSUAsW4v8t5n
/ejdEHaEnzrH0OYmAweOQfixrl4gcDqaL/GWZhPsCp5Az6sOuVORcNkg78P827yQ
T5KSC9iNja6wxKwrzl7YeXKILbH8oq1TqZzjbVVPuOJIEjuMszYxzt7A2r5hRIXT
FCdkDuZUxzmHTSiDuD1QMosdaQUM1q/+6BSeuUM4auey9pLrHj7FwPcKCnyg/cl1
qTOMJqynfpB5q1/rKx1kuNGCPpD+aD1bslMTaYURuawvFCTmNnndJscUyBqeVA7I
mCq3cIuELAHpiTm62TL8KsiWD88LghLu07CCS7j3RnRmSRwEbt5tDEv3XTE/S6qv
46TevUPioH6oMWKU0tcGUsVEkeUUqttxEF/niEhu8fqgta89FA+ViCruzMXIqDA4
VTSUz5hYYhv4GMxboF1UsNv3yyjBCa7i8vWyKQB8DB68uyJhuwVfziAkZpFALUCF
mP4lqAQ1SLtYVYBo4lMoH2Yr2UbvOOKsCl1I2m/n8ZiLLvmQsATUCs/YIqq4si+O
IZnubQIBo8gz3x8rQU9rwivsPsOBOJOfFghdeDNfRIbwweY9wy/vMG10yv4Wbec0
hSWsZj8BwfuK+Cj9hj+ewtVDZqqhi+4qOzmXvSpUocgpAZQZdMIXVB3q06OBvt0a
WdjuiZwWboJt7A57Sdlb1SGDRE7oykyptCrvyk0kLwP89Mrag2Uj7lC7Pez9OcYb
XS+6WD5V/Yy+Umb/c1FTCHCgI05CssvCJ9upwE9XnP5tRatsRP/5om29JZHApeTn
Dmjt4xESqw/8N2iqZDX8pFuJnVXY2g5SZvOqLX8Chf+VtoZF09B/alu8rGG5xOAS
x+YCiSY98O446r1nE9CzitEGzOQHUINORmNOnOYNP2d4okaPs1r+xjyrgdTZk0Si
WLkvLekrd9FBpevtpvbDuWCAkZpK+F6hzUT7dvN613v4Ho9oTl8shpwdLbroTF9+
Vhn4+RqMOKhEU8AqqXrhwRMrwr3WVrNUTIPNdlyCmsQG2zEG8qksoSkCa8tkrjLy
QFmu+yDZeCLvDYv2FojUfMMk+rqW0KQaDAJydY7NSp2oh4AhHBcfgusAcxqtPMvC
SNITV6zDzd7UBZZxQoKuEuoRN6+6AIvLUjgUmQv2YjiqUPybdmOvQNiECeR2Z3cf
eIn2M04l3wgFYQt+Vsrsu5Ov7Bt/RlL+YzwP0FjvcWiQ0id56zfmN2T7me8aYwfH
Rfaed+mNXLoIdB6JASEb/93iiUreqrv827sMh9JbSky3fiXH5KqfaF27PyiZgZ0/
50Zztyt/lisd/Yuddrx7Q08Q9D01e7PnJngWzCGieVg9fHwEc3zjhvJGplLHhklO
wbsJ/a2SsyTkvTDiJJpSKD+26vIpziri/NCREZk2po/24UhiPhrldA9Fl+77WTbS
uT9HcOtoPptADl3LkZlvqLaZyImKEULspGj0g2jxKj5QF/yyg2ZcjKG3ICdDlD4K
Gt1fBhugg6+D1CZsdm1K6jzI6fN/O80r3tygQVetDjsK4DQjPNLwbAhTIEh0lzw7
BQ8fAjwDXnqulNhISb6Z8dCfRvJne2xOylswpuf+m3YrkhWhv6UhKTpAwt3VchiE
ppIa7/aKpDhz+zn/phcM8Pi5NQ7hGhTAMOjWboLyrFb1bGeRNPD+30vHEYQouqN+
bd1shSXJlczQh35xYqhxQq0dCMBhNYGbz4qhqtHW0U6Q/H+4CY47YONfCAHs/Pcs
/sHcGbkuJAydhtqON96Q2uzahI1bQGh1bN4E1OGYXPOqyPmD6UdqoYPy0XoqnqdL
71t98FqxsEMTMuXppvvC0fR1LA3hxf3vyAdS7YBiwsYMXulBGaEZxowFd/Z80fRk
wDmz+MC0zKCHe98p7MtWgJQAtE66XTnUpqnEbDaxJ+QYvMh3YfrNIIRitBm1emmH
am18P2moz1kUg3ifpytH963YDlrbqGcgInuGI3AK57JDaEUtDNp2Q4MBC6HGmlV4
2yJk/WMiYnEk/nbTwKJIQFjOunNTj8a2Kr/jBPXPkPedFKwVQfzYIt0Jn5SGfN3n
igNJgikttihJ4+JOsH0b9atUQa7wkp2hVM0ZYHj7mSGuHsthqMVPGkITqCHvG32+
rBwCyqRY8cpQA067XGs1GYx344fS8RHdpl5SnvatW1g6ptBVcWwPTQphEcES+SIP
gb1LofWL/GLSE6NqBA6imOqHryITLGfGBwl13SJ+EDR+WmPiDr9B3e8Hnm/mx9nB
tKSztdG0FdK2IgtZRI0Nd+x57XJJiKtprKU+i2+gjO9zKdUUvM+yIDJ04f+bgmuF
06q2vH3ZL6fG6oVA2sISyz/aDqcYBXoVOCTkUpT0EKnquj7z/1sqUq6FsKg6xQau
nO0169Jz04TxuO18pl57nHD7lxnffEGaKEM9X8tIuAb9WkDJcJd3ZRhCBYMuHvwz
wFhdIreXUDeJv6y8X3Xzl8oVgzfFz9o2gp63h2YuN6/ByH66+WdGp3ekSzeiFM1q
UFCYBM/3nPrDDBPB/ZSqmy91tGTLP8OzH+PKvfGy693FBmXordjOfReBbSFl3Twt
MwXrBvMG0R9QmoI+RC05Q46e6HFVHb9vC5h5h/0y9/jkel0rzYfTzP6yTpzdm0sh
fZCkJK3WsHbUGqShKS42RAOUOT+2KCr3It8fjtjbNDRxmNn/NKkJbQiak3i4v5jE
D1y+WMQQoxCUivZt72yOR5/Ifj+vKQKB8yl1xbkUf7KuNo+gRCIx/K4etrqSq2Js
v39c0tLfbsoZ9OK3eUrheDyF72y2YUdsxwbF/QkO2R4ZxFFEGfzgXp685UGibMB7
kpOKM9oYgTKboKt0yNxRkYZPJc97gBTithG3/vwhKyWn9i/Bd3LgjZZv822rxpMj
YOFidGSqxFJizdYl6Vbjz4S53OuLyxajTrcMB3wb0AgYBuhmmYqVVJIlgmbjNCMB
5jYx4LRsFKLWsvzXeOiz94jeeX0z/NUfW7Lla1HZWfyjJ6zg7t7e18L3T4T+xA/L
WKHyGN2kJx/mc+gyMG97L3t308VOtuCfFt9MvFO2lt2aPHZZM1jAj2/48O4xyqL5
soWBLEfKsXC6b2aIlLsOTMmRBVTW6GueRbscr+Rw+kAzYo8rKDkIswOi0yG4y1Mq
adyDlO25X8xawdv5gyBVch34Q0LXLJ/jXrlBumfMNn/T56We0ALVhC12EjDehoQv
RMC4up9pgK4bBTtOh052yGcRxUShJfu8NfT9jAGI7Z5jESGBNwyFVzsqZRARFiSm
KVEIUFFFcNqJJltmWxIPAp/VDJ4Wm8OFkYgFUq8Yk9pLdnPvOdAQY8By7ZSTv6yY
27WpYDhK1inJjDSWDZ+zWPt2qrIVIAwMzl+jxS8pCjSOUAPrzAdG3lTeoKgsoSe9
oYXnGcUTYHQgYpj4LqWkHnN3bTHxMXbWNu4u+be+Du4GjV6qEkFgZfzLzBklU1NN
jSZdUj9H5QKNw+k9sukkJHCxvD01tAiNkKKpobwnQ/iivmbcwJEARbQ5glBjL9q5
ddBcDtzLB8lVaGQedKH5L4iQyIrYlxKTAr36DUQ53Kyp1ZdsssjVyDKWkuwtTLKv
2A1MsJldWNVjbT6tg8p55u/X+tE1MMAu7qNwAD4uSRWP4I3RJCyhGYdEYlsmY3lB
ly87Q7100+x6QFADDC3JV7PI/5hIqA2Qk50biJrdbNEhzuE2x1KoRr+iHBI4yKJn
0KV8rp6SFqhPOsmNliqIxw/VuPzs4oO1q0bwBntYXD5FN9AFb1cAyt4iAts5wBDi
S4ulGvBhWvje3Ye2YBcajA1GqMoUz2ml+3NOn0IM7GgkMUlSlnweog6yvCgrNoNO
BbuGwf7+ik+8ZQEAzpKK1E/0zeuDglJiEBfNVZwO4HIKpZtrd/d449rbhFRX6+Pu
3iCCqR+7gKYmbNgtJKvlKM9Uzy4hUgPF1tt3Jgqj1/Bfr5CYuJ9N6f5XeizRVCPG
Z1NgqT5kiutTRGlGc3BDJ6c8kT4bjhFcZvlISE1BMlz4xru4OC6Fmg+4r4mWz9t7
mtfcnAhjGlLklNlTyzHibAmsLxOT/wUKCBc+hsYJQqwzvJbOWJHd/2rn4kWCH8Au
XbGARFX7YvNUPL7EWa+bTun63mc0s1aPO+TW0bPvG1x9vgfrwKJhq73MgiqQ4Ae8
IPTaYUcfnbJETiPdQKDQjscWQil0PH++q9NJu9hOnjB1FXIB4lCS4h23xuPpTc4U
uRphrzukzUa3jafuuE9ODJ5RKX+Yoqu8N0MAGn0ALbNR7pRqmpKsDQhFgaYkOqJl
237KzojfBnak1G14BCCXEIxgBf/Biy8I3v1Q5kh39s+TvLPyGisrOPvrUjsf/g0C
pcv7ghCIkbRf8kL9ohJul2T+yQxIwXR1+1mmUfyxCuUiMXRj58jPfGp8jCa6WQ57
A9V3+42HQ0c12M6eSnouKOkrQItGgAGnWKz6PS6LXUcPn8ZQ00lVob+LPoWbb62j
ebjgD11JCT1XxsF7QE+TIXWagl+zmO1rnhEmu++7FPdCTVa7Aq5t5f8y8cLhzdCA
TJHIQ/KXtORYgcNMbYTg5wSNoUCA95NTUa16OJszop+NCCVQMBKjpVVn9OYC/S6L
aPCIb/8V60+vqDznMr17EQq4PvAGJIrAYvd5OdrSwfEjuqkvQylPuo/cM+amWk0L
vBfWs0xXNluj1qKmTLbjLzhfMVBKd2szDXOoYWLam5aj6VmmHzWidpaYK929xuf6
3vud4uBqbS9MPu6kSE0ehDwfGAa+GKTChjciiqVbx8EdQktIZUT0BGE9CY5inggk
Ihp3RWSGpWxhNN9SpVqwRCVxUpMKapJiwy46eFl/nPECmFOJikfXmbG9Sf/Q5zkJ
a8gYy353ryiwUBk4c8vOM6Jh2JXumy3NLc25xKBa3XiiSwxo/RpL5hy31/yat4Pe
qwriUvnSZgLWaIgXVThKgGa1lSO6yM7vJdCi8mNhFBfRbZK253Hghji3Btx0jfqL
ywKJu34/3g3wRZ9IDbKQCmgpZh437R7kUO+MeF0NqtNWOGBP/kRG4N9FVQMnAE4H
n0rFzhQvgLJFG8f9nVZpk84P8au5YC4bQRYZrrGAeJCRPJHGQWEj1ANSP+q7Uq4i
CyW5COB9DJTSZGaoDYLo22XmrcztrbTUVt2wShyvShXbQe0bqtDyV4EnBViRqANs
Gub0oqFPkHzJREIN5wuNKdQfwiR3VEc0n/HBUzjLeDxz+f2cZCB2GiC5l7VjKO3d
LwA6W8n0xtt4/AsLsJh6KhrPftxRKwWPq8zxu6AN5vVX6dI0i3vtZQLgW+IrTvXm
f1hbQU2zxhRjaj0bGBjl9SaPp38j+e6sL1xcC07Q8Xxyqx7OPlrSVrgH74/2UlEK
cYsj06Y68E98r18Hj1k73KUxv6x0HMmRjylViHAauklUYnopMsPKu6+63sQyaNY7
t3Q6wClsGVJ3x/ZCCLLa7KeaqkIFggVLK9ctieSfUdONWHsaQ1h46HeVDyRIgodB
Fk1abW8jdkWb8EnIywMOVIVLd89iwQzMpOKyEopEydYTsIyKrY7xFR1q7utOCQpV
oMazVfeOKCsOB1WiUVNnkWN2M0sftAL8RO0UXe9zDnh2HuoRE2R1FUWxUHc5D12w
Rj1N2DErRgZNG22reiCRKG750F8o5cm9Jc6Jvq4bVo7btSosIvOFNrc5Rku6n3Eb
7jO3gzV2Y9R0acVQz4zObldH+VjFTUx5ip2c/jzOSywkcBiX1wxEN5adqQxRxqFQ
4BBS+rxy4WiQxBrigX7ZHfSwfyM1K1Qj/K3WmPGB7gEllNIW73njrPxPncvcANWL
slzVtqqipJM0JKnCbrZlRFiivWiFSNPPv+OJ0heP55WQ7ODlFJ5+RUJI96f4jINM
LfFC7WMryTqwqnzFduHyEQl/E6Rb2Qfc9jbeif++sUqXwwR0tGWyHTJZOkKnD+hZ
kKgZOq1VxSHDw2bbvXTZKlYqZ+kOCqrxhM5xW73LFph4h4I3uJcpEr2lSVIY7lmH
hqkY/6e7GN0X4ble9aG1hc1jsKeLbMRELUYJdQ95nmshUprUipde8U7MNEQfVBj7
ocTnlwfdKojzKXo8pX41MQISXaL8Ops9S29xOKjLO2Wq2H8xV1aQZoHZdqqRyiO2
PrMnCjecycKjbSk2rYcsf9bHKbn7T9huu78pYPa9nrHbfT2hxGNTrEW9GwaX5a7b
8YQy+pz7A291xF8/NJ2Bc0dOKb39p6h+PzMOKVYoZfqmH2D1gBbZCm3FziNMaFEM
ldwK0arV9opufRz7bEwvNucfC74np47bSLSZ8nniVVeG+yT1UMJUj2lSWGKoxQvM
mspiMesv3eoT0Fxkvs7BctyoIG8IbrD1ZfdtgEuJXWvzKvUB8Sp28iDBoWZdpDRi
+ymZe185tCODM8vT5B5K+nxtQIGOGhbbXEV7gAPkVVVNQXGBQqaD0rE95jg0T7/P
9CYny7eq/597ZBaOCISQrzPrlAT8H4pHZJNXfXBfDpysNlQNpIMbmDIC5bRSGp03
BU8H47ZcCPH8RGxWQoaoitR/+Z1rNUs9tiM+ZTPOQuiMF3PlGufpGkb7x8rl2k48
rwsci9cr8OfP5kyutnXdu3x7O1mWJd8r1Y0rbbtaFlZbNivtm8JmRcPI0qYiWB3l
gjE25Gdchmnu8v2RYrupbLQIoSDqo5GJkQWzjfC5b8u809n9Cl1ZwVVjgZLApFIB
bNyqfP7p/10o2US/cGdQ4zdtY9wWpn/jCXFxCol2iIFmMAmrWWFuJirjNjz0OhRL
TCw080juuLW6lvlOUpsuGvMt1skD7X289UzrOFTXsdSnFdgWVcoJGUYxvj0joB3+
+nqWWPy8amtxXHpTjHAIUTts5jdGTkOSpi6qIc9pYozUYB3nWFeziDyNvLpaamSd
ZR4tnz0in8GvXqWOfPawN6K8/Keb/T73UPJ6nVZgBwoCiAEah1S5JmO6JA26Dh3B
esxuApgiTDXk7aamscX6ibpQenPSSxudzUJfwYcfFWUl4KmOgFTWbDFdnynQZPhv
3hY1+8p0Fd2MC46IktGvNn/za4bfq4cbtvKIiXPZ2uoeobb0HGMChqvwByiBHNS+
jiAHRH0QVZ8F+Gy+o9AkTciWmZcHNRl+oh1GKbRjLvELQh6ggVatmPnxa4GP28f8
M955KkzKQGBMinBZ+VaM3mHRvxCavNk1Jz34nXNBhHTdf38XJYNxJeBiAAN2hcfe
3Wm0gLGrQFjem4Q+ShtogbLqwarchTmnM+E7xqjB/GUEObIvMuvdes7MhNOtzzGE
KOdlKaSv6QPebFyv5m4aPlq6o7nCnEwOLnzWOOuoSO8TauDF6lvIPaAJwzuDEB8Y
IaIhVHoQjirYy3cQjn1ELVRbyq8P+LhZ7wKCBfP/u479ZdG8OUVDeODq4FOkTb+w
8saXGN/ivJwQ9sGG9EbtSyXRZ55rDEMEycbB9+TYwhacRyNNbVIc6xVqD2ZqW02d
YO/UbwpJ2EfPQzkjqIEyTqszfEae6AzvLUc8jbdMBjGNpcAVhj+oFHVKKcS8HVA8
NURz7KnMtyOrDq9Rki333pojUHHps9O786cQ6NaWNp29S7ixPwBGdcIL+I72txRG
zDhG8KoqBWLH5Xs3gswb9Deaj2BqXrzuJNGYxXEDUNizqQyn/L0foJn/sCR94alB
WndYpFNFVj0fLIVL3MeGgWdDukJlsuaqpOXzPx5x7HV0mV+gUU2Eq4Gr7WJ+vlRJ
lS6lfwH1NCGDIwXJdg1qNDeR3S5Nzvx8kss49NSWH3exzv5EwQj1m9A3b5UykhX0
C4UxSohBMwrvbT5k+mSG8e+WLoPinhSCumlRCGAjb+FDw6tNO8CTqzghhqrWE6nN
gwtXHesXv9fvdyTABHWXA8QyrRdrWBhqzTvxdZ1t5Cma13vXGQybv0ETDEgYwQ5Z
nrL3V8qdl2Xgs4oCEHO9H65Lzsu387CD+zCRKpWS4/GwPzIrZle9WOERMp18OKBO
VAR1RKs7+JyVAlykjxUNLGzJ8/LRvYJCOr2qn7sTMw3S9x5ThAUSV4oXiVO9C8ZH
O2AoeHwsyAjY0n7t6/bvFuzaVcdHfX6fjvqU42xWLKDzFI1UCN+jRjjDmRwbiAPS
dIx8Mw8J0XzE/KMxATp4AP2cQqw/J2Jwg+jtDeNwWiNBCFQ+efZN9+5AOlZNEkP4
DbUEKq7vT5cb1MYPCgggtr8B4RPHjCyAKpj+IDo6HzRtziiGVpbrW8Fj5KMA1bz1
wXQE9GHssv7+MSXozfXeUQDWzYUBpF8kloNZk35GExVTikVlGfjr/wetr51GR8Vt
bg/9oQffOdgebybHfOMcjnsDkBCIOqYzCYy3zO2WIG+ukeHmexrEZJeElu+pSCbn
qvx5fWfCDZcDcZgFwmku/rc9+hh8PI6oeN32GY9Aev3G07up4nvr5WJ6hxkpNHC7
/1tCUayMIfRnDLXp+kWXfnrOEgreZxp96hW2BqZHEcfLuqoa8Kya0BsMbpAgb2DG
5BWJzbLSxYRq+iatNmnbW1bL2dBFfqzaVPMTx7aWqOIL2h7yyYjZ7o4Am3IVLJEb
8u1F2dvLV9pXKTmfi4X/gXpwnxs7+Jj36UOwXvWjetTDEsEDNlBMifhf4qV+f/lG
oAIRRezlE1FN6BnVEWF+ZzzC9MdVHZ8N3ww8wK2CusWNi1MOOM2BNPoWrjXuRu4p
hq/piRkkqcWZwCV8CS4ZkOanY9NiBXjAyScQs0fdBgF8SieWM0towqO0n5UrnJVo
TGiGgZIjYli7wRymkscgLd6d5hJ0J8D2xQV4MnA6ASy0RkwQ1fzbPScKV4HdOtCH
D400Zq9Fg8qQvTtDEpY160MYZqXyfW78vXXvduwIUkPFAwMSMLWwe5kU3AOFYd7F
/WPWiMS4qCuUtP5ra5FGeL/rgYKQrdrCvm9he8U8WU/wQYSs4N41zksVTxAwWXIn
JtCOBuOFjRbrCZHY8ll0Qjli26ko/O+347lIpqtk0l+yFc2i7Nf8QnAk7kM6zpMj
2SZQVLhrGEIMYVPlgkeZaU0PVmNDZCuYSF/LuYPngdHXljoAzGIFgf4Bho0WOFJE
enISDDn8YwycOQE043Dc7Pu9KZW5TnAgwjaDyXHDR7wVfn5TEz9zAgxCsBtfX/Z7
5bqPsvp1u37/gEJvM/zYwRXLcLIGffpRjIQDMN2b0HQX14CYzRyS2ApZ4sBMpRtI
6nq8qfFmPlanYr/SI+E9uVyPlbWfYvWvpUsrQuHsUQTSSiezcelk2Eqiq8Kh+BVj
aqrvMUg2XVzg+mHOtuurIL3FFNWwENM3AFMAovoo68i4IWMwMaUTr0vkX4kVub6/
c5xkv+SXO92M59BOSLmOC3GSdQbEIrXGr98VcoHIJAt8RdnAL8YIoSwqkp3+ketX
alPYbh5XKz8kyRQkhds6zsPMvdNuOeC7KbVf6lnkOmDNSb+CtI/dHl93e6ajJIWO
y8j26giyD7+EIIq6pq2UXu6/eVztH5kcOx4/kwxeVn1NCG1SBqFQLs6jfzOqogP0
Tw3tc4CU2cmA4oHzM3OaLQ45UVpg4ohpHRUy32JDu3u8fRpfnLh3oVppSMeS3PJS
fFhkWrOFMC+dVVGqKJw6bnQOWbzfPsJf1gxmZkDo2CSZrEmGT04nQBqZYhsS/Lrj
OulZS+mbTNMLsg7BSfunixOPv0yYFBSH6N4mfOefp/LmAVMTdAbeDqG84IKz2RLw
aVpmI6mnHOdgH7CrhFl6X2mlJD5Gg7TJ/fUo+3JGWMV0Mq81eTU95QM/ZgmbgJZH
mjUJr3AJRabtSGXWaSaGZKS7DDY09Y5rTNvXb3mbYWRyXvAEBnEbaW3b0Zq0hSdG
+baU/V9OAydZLSMQ26FNypB/HCjgkNd4ZYEAbzDC0s/lK4Y7SF1s+hXr454hFp8/
w7rU9ffslAaDehXV6oCzvS0ZDJuFyRqvbNGRwV8zhSi8tuaedcjYUAyivRVFrzy5
TUJW0GHIqh5tTZaXHyRHhk18rknFc4oG8XacJLJ3XVRDd5owANX8l6w1xTRRHJYn
FZNTbBgyIZXwA/wb1+QdlUmuZ8KSOR8pKn1O9/BVXJnGG1yD9mJg17IWpoLf7F1o
Nz42jF3wyfu8Ew5+qAxWkk2cm/BCSHDAkKQrymTWnXsagUCxAd3dJKstv655OiAJ
eBp8cqNCYld8JK8xNcOGhVHpnPY2z9wSMqRS4eaxRkmnjtWgiZaKPsd6URMt/CBc
ct7lUHADDqVCXouv0ESLujq+AtM+RztMe1Y02Uq+W5dZncLErVKUAu+nZrcZOn8D
RixCwn3Xqf8nPuKXn41Yybj4EeUpC0AOV7CGXX8vgxbGT7/b0V0RzSKcWJhtE+NU
qavgTHxrbryJJLWNR/0pTqodB1vL/ESOfBa0fwTs0YHzoikfAutY+4nArRITcwWm
tSOQZJe2qrvALtyUytBAN458Nub8s+radUpvMR9Uks6y0THZX5NWeMEjcSb2JDSy
OM68y6CqA9WWWYLJ6rYReTLJNdkKouFFjTbVQxnSof41dnGkQT+SIrbfgRvMgZCR
KF6K9udxuuCwVBLoOHLCPFWw0b4jn0xLCP8B7eROQpdWjYbfxiwn2a12yBg6794G
zSieiKDc28Jv0Mh/2Y8NJBp18y1N67KgGAHiffgZ6e+lz8oBY1J60xdFMXRXgArS
uye5JgKvR3VJwFvuTZqI4hqQd7SkfpLaKfI6d96vMvtYy8+5I0c41JwKedyFXeGi
/PF5pp4fGEuW78d6QbcjpY4enHCy/fVgYOfCOqAUHAltPpNI+vFGJJyudsd3nx9j
6Eh1NyNzAM2KwEf1+O1WEZVp+zLSYFaCQq3uZsyxMomv/U5NlOu74CyQZzVb1Ylh
a+8+8pFQnFTDZSA0PlwLGZJIMhmqylbLEfcwJ4nGhMxLq6CkeF+ZHuepcnmP9LNN
nuMySy6Cr1+KuFdMLKWSs2RQs7fEBTA/3t259SoumAElAhcyVJrKZwNEHHV3+09c
84MB+AIZnq0P/L0OK7B1j+vPkvdDgvFEWVAiQxEJvTc0ZkyzFpOS32ysepJV5IFW
e22+AMJHGBpxfIsOI6jB9HNCXv9xDKhX5FBkT0KMalCAsmrb9r5Dpv/kPh84nvLG
vLYQe5Oo78HJe9KdbzEE1iAcApqge6e2GkllhcHdv4h98WNStXefzlUlzIVPyV+o
oZwangMXix6LQPIR+21Uh7gK2J4rf9HbMOV/tbJ6zmZ3UAJuZHhQmAeOt91OEr2v
Nbcgcv6UPpvf6GuFzJwupPSmbD6BctE4vK/7oqxPVHPmzQJMNJ956SEzwYVGKylE
QNyRSbp31OKs90yzegHjSUjaSM7KtCZhUZnNOvrbnIWl5gypC/QSCPW/V5r1I7dD
GB4wvIE96izf+Horz1giG7Zw5eklgu9HrzF7y9szrtw9E5vyhqpQRI3ZUVugy1Et
KgK9mQD/+5k4OnWOo0oDts8ts0wwRVntcErRsNSUdAZCLU5stQ4Q9Q1EWyA3v/oV
l2+9wrOGVb7m/opiuwLR8+DpL3aYUBtIMnGe6yUEf/mBDxuNrEe+2EmrR1jSBIO5
rKJdmgSzfoL5pfgIBBkzJC+A8Rh7QtNC4i5NZamLd1o1HZPwSM2I0yJSt8VRDLto
JQEV8bRlI2Dq9Jy3FurZeiHL2Hutz3Q8mAcYu2GhGmAL4wktucxy/XUw4mtxdI3/
4LcjO9tVX2gaGMw2DzD1skWOqAKPs9C5ADo42Y245C79cgXJT5Z4MQtHY8t11nvp
jQK71YKKfqFEDvvO/9WR365z4H0fY+Fg9Rh/WXfo/2lgz2DYCnflJO17sFsBM4I/
4JYDji7843+K7+7Kav9fG7QfO9/i59PXQZ5q0JgXnWLMAFUgrsKHM6j0td2edcgR
EYZpK20rfHIDsVbCj98xDBCtxCRx58FTCRQOBMQ0KcUQ1VRYJAZGyakyqmY+eK3I
kNaQcnxBBrcfUbiNvFUmkS1E8gHNtsktUSDMDwfZtx+vQ+Y+diQ24Vhd7Q8naPty
cmHvZ8qKkBsb1Rt7jh2z8D56AV5Uywrkq6BmdTexBq5SZ3Xzqf+uTp8ftuOXhvNT
ipv9iW9odL4FBnsnMutX9OTsHTLz7dTv9IQ9piMlsJC/2URVVOvL3vwfIzsCBg0k
tMhV0GCwH6nHHXDY27j9v0I+T3MTUaeu7PMRCChPJoIRkVHcrY4jYtJN7YKnJNcI
jpSyu3HbQKab1a4Ka8yAjVOpHyItovQd5wMi7h9LKfrKGA+ZJ31m2Pa8g/llcAGZ
fWe5382EPIdFxeR3v0Tbcv3grxDlRmxYhDjiuTPOxd7puO07GKRna+TISph3Chg7
rF7L1Smurx/Y/0UyBRVgmetOQMn9hyPt31IQ5neCcBNob1IednR0XqO3C7i0kfrL
l8pN/XH+jobXtaEjdcueytOT+vkpMwSNCSDVjDFkPaepUef7UprmV9oYyifSIx02
boLrdZtfj6yj6OwbdZ/BsrOrty5l9aQQ9Pf1uCWNiYvxN+cTURXfbqdXVKzNIwnG
XSdfVaD9hPBxu59TCgr8xQ5VRfokelRQODMOCILG0KeijpknYe+V3XMU6+Ex1sTB
mjxiUwyLy3ZfEVAWhehkATsvKdN8fBKT+TUdL0hhqKNWioG7jLl0Vhrr2mb+WGo/
pRnVJ3A6Up71dvTH4GUSUNgMARtcpwjaJAR4GKHBS5W0nOQnOeN+hfSaQqwzOYEd
E+JFGsAUAfPe8bk8pmXMSxPTc5kN4wM60IEz4gBgUzY0kfLtze4hR5BW9lPwXTTH
wm6BC5MazmuCqW4pYX/hMWs5Mj4MFLTqYOv6LWhxi3A6kSRn2w+W+m8E7aOhtOHa
AHGDdEIv2IzQVEGptHgW6Z9JmZSEvMz/7QNp7+wJ0/ZCrfRUcCXAOCTxDhWqW6UY
NaMWv70JyB0w05ozmUhfTlmPkmoG4PxIWQ0Dt+Lmoj7Z2z8XF4h+g0DoI0yFfDbS
oJ9rNe4oNToIXFQBaC7LBik49aVrp3bkI+5g885bdEr8gxJ0nMKFqfq8iFJOLtlp
USOVhgg9C6TZAGY1LuD/fUluXYZ8lgWMMa5I4frnstg1EQXy87xksLpu1R0iYoyn
4slBJbXuLgJePrpHHTL4hpKKYJOx5/8kNndsij1FOq15zrIJvn3NlUigHOVi+SmQ
UThKeV8/MkgL98Lgj7joiD4qKr1O0HVWPgd3rvRwlNMQdpz8HM1PyVWhtqNzXQeC
YXwcrqdpW6d1g2JTMT34V83QeL/JSF8LWSgygRMkiYlEsOJwXPpeUuCcfhqTqeT0
HYuzBJtYNEqKmr+cQOdRoyaW/a7OTVKS89A5IUJ1sF7/H5sIF8nq7uibF7jj/1fy
H4714jVFKXHWEzJ/bpc/ttrHga4xQmgGkbRssPC7xFZoScTsHvnEOKU+7UdqleK4
lVGiLIisxWbanM1BXnS3VhH9kqxGrH5zk61XU4WUihd2PMAPihYYQkpvRlGU2AQ3
kRoYi33higMncX+j3A7NK55r0TX/EHb1W7u6UoiK143RjwMhkaoGdjF+adM0+HaH
mp1qFjQjW50Vxpc79pZqo/5BXR8vuwQIxXb7nvYdz3K8gmEOMfB1Xz8gxLgNGtzB
KNvqTTbryFrlGBJ033liBSHNl5sxS58tEqpcCTK+lv70G4p+QZnlPHTt+cNpk2WU
VhKWEPcX/s5FEw6AF5VCl6W02jKjCX0X/16pOllntr9cic9Epz8QC3cvAQmI0qwA
SXGCsvIDNechqa7DxWoJL+cWDnCOG+1A1K4ESslesfrgVpcZrol+1iAbFwrTPcsL
ySGLqxkU9M/DqbhTX+fH5Mty9hDAYyNtrE035anmGkZSDASJupJ8h49V9zaRdm+f
evqtGQsaN/QcfpVHqPxubPABUADAoBoTSX+3E8OwqhnRgJiJUeNAo3IdEWnC/VbT
dRDHVm2fiXlyQdDk2LTEsKkRaz2+kzt2nBJ100LIID5ypVFWMomIOeQViV/Zd/yU
saW1JQrNtPzPnBS/ibcbGvdazmON+dVo1eNBqP4cD3vVXGUzbGvkAdPlfmRV/UVY
OM5h5mEkpSdmQViqjt3QB95VmTAArZmt4ZV64+7+9Bla3G0k5ADAI2yyiB1bCJLJ
YEO+k78lk5JYwtSmLamo9DGLKhMNSuV6KF2Am3WC/hDEC8/4g924xxh/cz/wD1qC
Wlxuj/D5+WvnvH/clGmctYW2erWhNrDJSb9K+5nfcP1VHMTPaHsxR5aZjcFdvvuv
LeSmXhD2e7Hg7LVOj3xnXU+AS8+QYR7FyEh7hm0idMNMpDzV2RD+pRdI/LXcGSTI
p+O6UjXCXHchtlukNsfEiKTT0nacVKUIYwb86BWc7E4TrZfKQBzOHVhCKqM9C2qz
+Rd1AB9WGvr6SqsfJv2Py3goeDHM8M9udVDJbMBCDOR6C4mSh8cMcYbnCjipl4BX
9YqCmkYXQUoXk2HD+YiAbpaFz3/bvuzudtbqpPfcrx6DKYN1T2sdbwam3qFfk4IO
LEtao420zVzoD7peuaeu2BX33vB8Nt0AvU5Vtv1QyjIiawv2pxgIa0FyPzWiDDlb
rI5UZc7exJ3mmuq48cV/NPUUhLGjU9gFRN7NCdpeAuIy2rxjM3Cgtx4rmKKj4H6/
7nEDl4G7JVYKPpc2oqSyXifxN6C3nBNwXqScbMY7fg5stWD5LEzzZ1J7wtqxL0Gn
uIUhjqXSj2fD1tgtgu97nSK8+pPLHID93zi8Xv53yZdWFmH+OjpuJbMLwAVgcNmb
r43Hr5BZXq0qpQj7QsU1n/oDHNxt8Mcsl1TX23pMFQO4wttVawz0R76XHTK0dBhC
5Do8ikatGBmhXO4XZvOeYD3QpcnANmR9uLCf/3/aMpa5yAzxk95PmjtXhUb7o6ux
0rDTqvgdcynTZ+jbQrZPWSTbDLQaaCwJzR8uGiEU5KnZ8TN6Jm/yZpylfhmys9xw
LeRMYZZVqpyAQOAokT2iptPeGTeWQW9gBNWnn1vzIzU04RTuYvQyFNQJRnGGuzaI
lw5qRBML0AIPiJlCr9iyTUich2LT8+sRlA0VAfulLprMOG98MkqyiF0lDraeo2N/
fsxrCdeRnWMEZZzucwMSEgTE6ew0jMT6RUXInTpjhCHXndq/HOdzHwUpLl0VMIrM
ybsWWt0m2mCKRl3Ht4ElYMYJBNRbj1alOTU+k5U7ZoonNEseJylPKbaNqiNiFYa6
IFmCdOfN7dLPBbZ/siLd06SYoPYAfugfX6uJbIvs4eGn3AEwoi6ssEFVCjYmGUfk
MsN4zuOO3BEO7+XcpBTI2fRwCh/ux28V37FWozHUqI232eTRQ0em/kMY2JYEkygP
NjLbfydEaLGGA4aWf4wC5xCBgxMnVzjOo0994bJ6ZNNX0wiufOppe75bJyA0eeA6
EMHbPr3H04xxaDojSoknGaZMSE4N//B5jxeHoJ/Odt6XLg/J3ryYB4KWXAW0wJ5y
xaVWnBujb7o1mAmtGDTRABWfNK3FGTZ/b/6YkrI5qXUQ2diIKWmUBeJMLUuKpBOV
y59Hzqb9iJ/nSXPGBazVd6l/kuvt5Hd1Fa0ze25lFLnOgS0/+Xe3LPkM8gp/5bm9
EzNIaSBcBHkwnydrExaVQ/znfd948bO/7obQWMMzP0bgw1pVqY/lXLNtyjNLUcDx
hqp9jkAtwa4lPhHs3BNfYn+3yGsW1qOnWojnjQbgtZDKzoPl1HlW7K8vLzRfpOH6
08eNdS7mTOX6dUw4VJNs+8G+uGuaEw2CWuGNx8vtEfjhhhdvLVaShINXyWtOlfI7
OyKgWyVjV/WJFR+In5f+L8H7AYL9zj8lJeifU5OhIQypHO7glfNfxXqLB0kY90pV
/LTdaUHmAb8I/aeKIjlr77k6UzrvGsZ4VUA/Uq+Cu28w0xKWIvHGoeBRwS8vzaVq
4piIWgIbMuTKRvGfMXS5P9XtsltzirtqD5rSJ8CWQOX7FNmygk4aKkZ6YtPe1H3k
qICr45Qye/G5tA1cnPj2CMjZMCvpja42boo2rkz47WWNZneIvwnrvK672inXgFtK
mAtvRZu17k2cWBZPUgf4ssd1+5kxlQjqGdkwiKaJVWkkn5KhrehmcjyQaBQt8nR7
/NK9ZlbYMqGZBFYZ0jwS7yBk7iKR2VsnKSW/oy7JRthNw0MEfJ6vGXCLHrBrJBxp
8zqwYXpgm6AAAOgknoih3j1gHlh1eEogbG3DNXwah+PxjHvVtQqVpl/T4XHodejZ
TDxa/PbcxAcx5zjF+UFauCJp9SpnqyTO6tZG5LWWoYGVjY8zy4Fj8nH3GWif4J45
qxF5ekcAkCPCT3vYsts+kriuNndrX6nrSnNv8VQt0fNi05ew/2QgexGiv6ZinukI
+7xpwu/uo/6p63yCSt2L/yAnKt3s2/t0iCW8MXozogJPi3GCdTWHLwSxLgAdp0jP
QGLE0ZVTNnILAhHTAZHADPb5EKi1FLAirciTbddF73q4Uv8afzMpm9W/CoWRlkEV
PyLxmWo67yq13wMLGD4uz4ku3nU++d0o6xsgjMIVdV9XOcSResYcv+z9aQSQ5kje
z2fHjCB45mYsl2y6jgaRYUKhW9xtaPCusYYNuMBMgRSTYjc5FKt/8eQal1+yA7jH
MaM/4S0D0miFhXPrMAPp//RfJlEsbGfvBmfoarTRqokO96/KMORUIQGuCd0J+LLZ
jf5lsO+9jbdvsZcxFb+defRLg3Zwy/hW8/o+6hM/Wt+tv626X9Cn3ITJdc4Ulhgm
EtzmsClFnB2+Eyhz5iPgZ4nuI6euQvp8h5MxFpkIOJymZ85AH6flqsUyM5YVhKwk
nZyLiBcnf5gjRdiKEVZ818qbaCd3xg758RJAt/LTiRN5LLZ2lspdglZcTRDYV59H
MzHHJEy22e92NzhlQ1oAtv/J9VAJOIR3EI5kxuPisQIui/CoU9AKm860bucWkGp2
lB1zuxuTXqpWJfRpyrsEInWw/WwKM2KP9wRXxaPxWTfwJ+Gg8Uo7bh2xWp1KkvER
HNB4ZeeXddCYNfFj1jaGz5HaY76fSmUCmRxOX9tslg59TjLf2z9cyEhCn2gobcsr
9a/Gb5czGNmcHLqktGzZZqlVAMuk+7HjrVsR6gRT4wDE8q+8YgrtZe8HtHr8KIpV
dBJYpS+xp9D6fXUrTgJr9jBc1RfKWTTrtVIf96QXWNKFy+Fn5csx7dJPrV8kunbr
h1T1K1b+B8XSSP2NU1dd1UFaONxfgT4g74gCreafeDFVtTAMlPJJ/MtvrClPcbnX
YXuNbX2hhztrK/zeSc7pvkqlokP5rDrAjlaI5wSXxaYBfOLg28RNIUgW8BLvPK8N
vgj6frmj+WX5oYqX85zsuhoIwICiYgUOmNcgN9w5JqLXcytFTf584Txji2nfy5g0
C/b3LLVt8Y31qPdYkPDMIHduYHhaSN8zeQbcc9bcNdLKnXkrpkL90e/v8aLhXjv1
Vq89EOTnL4AcoUtSeSz9lWDfh/ukMjxMfGzanYtvDNVTZD379X44UxEofJZs9uiJ
9ZePZm7t9dCrlS4Jxg0m4rAqjknn/Hm/OTWZzHxsWksLH4jqVvZ1uJV/yJbrykIq
aBf9StsCsaWAJq8zZMU6WK4n7Dzoo4gVLBoPd6xT7WWnvibC83ha7ssQA+eQqVVt
/MldeHmamKJyx2tGoVj9YKSH9sOl2XRnv+CFPKoskyCcqI55+KIXBXJADC4vQigF
e9u9d6Y6v7HC2NNB1qTy/opCRm0fAwr+4dRGovaDkb22w7yyOyf0FCv6AfGuhT8i
xOWBxTJHToYxgWwk0lXeTESjZb6AD76w6AkKcBHo0TplRixPQ8sopXTy66syqIKC
QoYbQ5VRK1sjk0XfYCq2fzJg65+wBK+uPYEusmelnMDzmb6OjT9JmpY4duz4T2cj
NaeZA/BLKcqFYCXuAZQcm4tF9hRqVkrHQE/pG+DXmYXn94Lbfjp0Q61keoVIj5vC
MEpPJZ7Ay5hpjUZtBsjU6KvzqIdjKW4DrBRuG89xsUAnFjLUCU4sUxN9FRWefcfU
XPtKgec0d98OCyvZWWhcVTjO1TL+7UTiYBZ9as0v/nh8sBNnDVqUArGnyAZgB5cy
VSPfCuUv2PnjccU2aSDibZPiL5YqNEptafrEKiO/RdEOHvR36PPmOMwgsPDpa/M1
UUDmvp8HvWFxlkZxFI9liq4LqrqNReEFZf05K96waeUokdyCATlXcKhI4OsVRkT/
CXg0CilE4J/dDQBk9zvJGL5XnOvc2TZN8U5MAt//WBZ54AVZBeK+NbHxQoI6qk39
LbOWLyzGoAKvNmReUxHykuVkk6OC4OVXvD/3L6VS6J3HvgLFd2PoxJkQ7TdY9h2t
OnqLKKQQ5HxT1GOMVYy1LC4KRqprRyqDaVaHXimau1rWce/C6r8bx/gkxeEgYx9A
27YbM7duwSze25CX8UkqFWAuDZ6RbjKi8mDGUPl4IUfDgdZmrtZTAOfXqXdOibPQ
kKeWGdSa3Q3uPSrY9Zoyx/knlJd7kKJ3knerYwLdqDiz9c6dtSkKeeq9SWJ5fzOo
OFPv0KBYTWoMrnigcWfMje3uiigxSdk9GDe8P74x1LQ0TgfCLYWkLFm4sr6sVx2R
Yo8GKSv+uWHbsVz6O7kIjf2nlr8yp3nG8+ut1RTP5zK0j61l+2BBrKeaE1acf5qL
sFSlT99DoLXncX+RSIvP1Z2t2AE0LxGrooIebQlv2IqnV/75TJe0FWkoQdx//Zlm
xgR1w47pao9GVMmNmqLuC6O2O4hTfdGxRZkh3rzI9Dcisu6YDx6WxMCQtwwy3jLH
YVBBqvOFKpUKISpDAdFXtsIqCwJ103bE0nndcHFdgC166zSu+az5qZ4aAEy5XJ/P
OoCkeweIx6gVUYkFOC8Q9nXGJMj+qz5vQMRZltNURImXU2GYSkpPH54tC2OuGS0k
mBbKQB7tpEghTQKQFuK1r7XFTTcaH+K5c36SVvgYRakeIzE30JDUu5Y/KvNniGLv
gi4G5z1FHUkNm0iy4igznUXlt4VkERl2cmiUkgwNEowNCnlPwK9r8/PlbOlFudKY
6yHuqF+M3sEpflM3a7VmZzs8eO7eTf8BdE7ppmymxceJWpCao1aYSrfk7QRvwe7q
/H76gCAU2IRau90BtEMOvpyn5tC1RKM0ZWBvEniO1KvZz2CAUhNTwLryB6Ao2I5k
Cly+tWUlJy7QN3EmwCa7D8P7FEAhGQPwu2WoWrLiyynjGNgRUHp0o5efIZqGXQTT
FGygT6f9W8biehd5hSXMTMBIZ7RW3VBFJJKtjj8JsiO6Op4mEjNVeJw7XYVn0B6m
yC9sEr8/qaj6orllCWGSVjGyLFyJRWoX5bfyt2RqrfzWFwt7nDq8ZvuuacVTfdxy
uCf93umxBAAj+rGaTMGL0Mu5krAngZ2p/PcWlkoK7HqLyuLvyZ4HYzZVJhTxwBRA
BhhF+LKYNVywHDzY9jfWZSfmCTOZmaVl0+CxGfCYM9gtI6AL7JLFtFXtBSBjL2na
a21hQd0ZA7J02qFXpbE/vPiOZg9Dt/19f+L3Nd12F52AkZBw2RzDHBNph8sjE28N
xSJ2MUJWi9D8TE6ph6JmkaNAZieVowJYeIzMSTYqcimtKdvT2CSH3e/+oswNVHaD
xwdPNYyzuM4vV7aYfOwAkzhmkmEGZnNHEAJoM2bxrbzOdBIbNiyzBFLYWRgi/5h6
eaZLAJp7kjGVhVX1XlVJiv+UHnOsI6OzxNC2Oi0Ktr5Cv4Uuz59Tn/xeE1hUyNBV
CJ+y6iqCG9bJ4qgPziOK6wsFJa+M9i9p5k0ikwoE2tu+78GJfre0+CuFeok9gaMe
Ha6iAVLphgVAnvN1zZnjYUlPMLJl1Oc/yT3nled00HsauzRMoWi0b7E77xEQqSGo
obTNDsxJ4QMUVYlGHc8ZFFD/cHa8KjJMmO7hH/HVpw63v1B2j4e5O/63pzA9+n3C
oJrzMnc6BllI5OaInSUaXRr5W19jLlZzRqNQM2PD9kytld1gBWPvffkSWhxCFQXO
HfDMU3mnChIiuxioSIC+t9ipb+mtzYrGBBZvi68KJOGO+xMN5NBoi5lrLgvK7AF2
eKF0rimjdgHpsxZwmQd2ynfISA35t9h85mtfQ0rrg/AQABEUiyfIP8FsZQEFB/15
+ptKCIhn64O1Pe0V0/uqU+UG7286Zdit6I8jVOGF2GcVd+KvKCghkiD74BjrX43P
mp4thzTKaFALRAPWs4JfEojBDVmJdqn/2R3JcGJ6bNd3miyi6YHGW34lMXlzJ8Gn
tsM0lu/hzUQydWInVhMUR4DdwICbZCSh981VJuo/AnEi3KPSQhLx1W5rdJbFKm6/
cc4xLUwZD40Cgm9S3+4PtPF1dsfZdAcTjLW5xFg/eKpAj3m2eLPyRXOzS0yFmfig
nBcnglfGk7qcRxjhSEfIMazvx/29exwRp2qNOLLcyE3vPG5ZCLMiv+j4J5aKUmAJ
JHbCkMJFhIsi1Ncswf7WzHhCBMctAVQwpl4ndjnGWxptJwmrbewFtBBQBq/9RKVV
RBDxAItbGF6WyMposNtbeC/okXmnA5Ttrbq4TObMcQcS+H4z/UINY3cnE2td2fUE
Y40Wlse/0J0tge0cePWKzIr8B1mSzGaqP7Yhc/wogGvRH3p0oZn1MOV11FA3hnVw
2xlwznQ+Uid4jNRrNBa+7WVb8erpzzKbVQfI9oSYdxOLerzsFMlbVb/284Z3RXOg
BCqAb21HwA3u4aYY3iXhRA4KJPE61jl+5Y4jGfK0D8oBvJVH2S6BEUa1U5/CbfEZ
GRU4fHfjl3XyFDAyF6yzopaEssfAx84xs5h/w4eCfjTAeJPKKPTSzBYXx1dgBTem
CIduNQGD/PN2MPYvzcnvl2tXwPYFEFjGzd2r+lGS7v63DEm7Hw44mVlYvCE/THc3
7TW9aApTIT1v2sT2Khnaz+/hM5R0vYtS4ChNyxxfBpV3Yz27F7s7c0MLCynz/W1X
OlGnBRL1uh6tjiIJmwG5ZzQNtgdHN9uDL6/6L+PvrtfRXBK19it7zDchWmTLf1DD
R39o7KpKcSLbY+2f4gez71e9fUeLSokMBLp82XhBNmdwNtLwWluqY1Sn01gAFaqm
pxAW63A6CoFi078r/g8D79wW/uIyHVfL4lYmK5PY2fDMUrH/4GGamvKBL7W3S/lW
OaP4/5rRsEiJkqB3g2pxDUgYs+xhhkwpTaJHDuBXIr5XIekZb+PDnjtF4r12ybp8
2qu7T4L7BlskhAe1UTlrt1WzqFSV+RaKOAmvLWc2/JK47nLKZG+0GPNevc2w3bQO
lUg+rhS+9p07A4KGFy95nKFAvuyrYU2sUozhWk3e6La6mEMcfhsVoijPvvqGXsvR
iXcotEPGC64yC3SGgusRylbQvLmoL43DnDSucDX/oIXkh03wh/UtF24j4gsftOgc
wM0gDTVB84m7GvuHU8i9aT1lXRVYOIYxYP2lxsoYm+8xB1VRgeP2zShJ/HQVY2uG
dfT6PUJi7TcDETzZ8KRHC+PZsKOP8n1AWiyNbB4In3gK8FAPWNsM08MphVjhkCF7
gW6wSgx5QO7F6eGy6gRpRabCblN/LByzN9MeWr/cubGUDc35fqxdPOhL5LwTGm3M
FOapJ9uylNwX4m1SWNoVtweGZjUXeglxyv5NOe5uoGick4qkqHIvu1xcaC14qzHT
y+1UzyGIVUCAXDlua0o3vEr6WV/v6c8n8ewpp7ThqP52uvNK0z2fd7eZ8SPNFHn/
aLy74BnhXT+18joUh7WA365tjlr52ZffC20gTroE2UisQwqBNRjSDD7F9D6Xqxj4
O/H9Ln4DSDWz0Omyq/QY5nDR9YvXf14RkxRkJgfvUjYW//P+XClHKHtTT70oLtw4
8Oe1rZLQlqq9/k8Amn8lhphCIeKYOZO8DS8h1AquqBBgInrZ+Q5ROO7NTxDEZzYj
h1mg44Z/MsDs+vqWn8JBlbNx4PNlb9YPgX/uHhIYr+USafPqL0QGQebLouujNldY
Y22hM5fO7FGy9yZYDBiMQBJOLEyCqR5Z/mrxLypRsNuH/NdyqUosg7YRLus2HmAc
oVGTtbDFpoCxk22XBjIe9H2L/e/Cs/qH5d59p58sU+cpus9M8uDsdXd3L5pLNeCC
3+uaHZMebOnSYtoyprx31dzr0PWKFjOytCSvV953tIPzn6SC/TNj+PhwjTF5g1Az
81cuh8EzenZzicajLH/DmaVhUO68BZeEGBXD9Zk1rCanDtryoiYoULTaqyBaGPzK
CrY2TmEM9P2lJDKdIKqATlklzHdooxF70jD0reqH7WuMZgHT9Zz6/lCvTkq2fuo6
mmda2rUDeLKaj3iZHJm+yONasOF+6K6A9B72Amgw8Mettw+1XYoKf7VUXPBQmmG/
FL0hwjIZF3lcX4MJ4g9mv1jyiYsmeRya4v1wB4QbZxqsAjDCNYDevXaVCHWb5u9u
eEMj0U9fWNOR1HRck6YqwUiQwSeBPmz1zg+eX6wAwTLlUzufqB5pbvbqnmButvB0
UMt+8ZBoQVlVJ0dqWUERD59KcbvAk1haOdjnA2Rpi+vhNHMDo5iqVP/wiMHsXQ6Q
gWEqwXPKuu0ge5ovhT1bLLH6gayDLPatKLYEYnk6NTMU+qrdiKvwOch/fJMtspdC
CTDSrD3xMGhI8q2Nls/9PtvEo0ZPNpYJ/mkuBltEKL3z4ngyywlcnGfThf1thiR6
cSyrzgDVkZJP5ZRkv/XOomdqnAwAEsnxQuSpcszUzO+BSvXLOurIZNiJVD9i/neb
TaDTQjBXGm6DYDR7je9pbHLV+qNXQTXoubkn3CN2KM9pa+hPVxrx+WgOeEj805jR
onDJ8Gb748O4PyRu76wJMJm2mFrWGB7Lwgj5jUCFVx8claDvV5n+bgPcR4Ufxxl8
JodyFfCMBeVvfVCRAjICDRtZtP9vospbPbfgRBNtXXYSece+/kuJRnWxEbQ8DMq2
DM7jPeZ4Cwgr54tEGFoTZnArG+yQYAjjRkovuYC49RFIx0Om1p5OcUlFbZd2jPn4
FwS6tbgs3CxjblceBqJLCMlXYMqnIEnMcDRh/GCTyBWqwPCmzBFn5Kgh8N6Fhur8
NpjcmNpjovRmzmu8bOc4DBGaW2tnxuNGshhopqwrc1yBKUE7zn2RA8BXlilf6MJn
ICj2sZFLzggDQ+0oYL5fwsXrWOopMpm5O6CAi+Ubx8VeVIJtJnuP+TEkk04gjYah
/l4ML5HoY2Kf88QV6txqKti4+6MHerksEfsL7acehYdhaRRY4bCnuYvmtnSzdqaJ
ZKRx9MpfgoNUp6KAyafuteqIqW4vaZKYjLR/6j/G154qMfdlU9mrjQtCjwtIb/UZ
3QlAPNEgR5DI5KRQ9aTJKwAVYg9fcwDm+F2TFadqQm9eMnpeVEsaGx1o22L8lZun
3TvfvAN9o16q1j9aOec8bl3GMCbkNW36+l4Cu8WreQMA8q8Gb4k0mv3n5N7+pL4k
FPw0AiY1BjH/vj0wGmxrTKC0vNiSVs8Lpu2AN3MA42gEy8P8Rs8WX/QQn9KR5qS4
r8ZnCAgQlTIgV+k+iXn/86BlmQ+uDZf6ENu2vVRTeCxxus4VwaM0KrXfzzgcfKNz
n7TbEBUG4REKWQ7PfQsQ/RXbiPExjoE3B31/GhhGFgRmKJ3INXEDa39+TUxT3X76
sEFRv3OC5y7P1x0rlF/aLi0t3vF1ioocSrXEZxrxbVE3O2l45y+75YV65PN42688
5v3RPVAgStR70xSRw49mac6SKAFK0qJmNS1TnkumC4xiuXUbA54Z10v7dhwlCsrJ
7XpNTmUvsP970K432rP/H1Bo9PpF6zw/z1h8tCyhPzwlOeN7dLDr7LyU6AfD9pLH
gZAAstYrZa2lhwNIoZfPC5Wfeg2deY7sCJBkWfCvSObS6CpAiBNhPzdIKrVUbLfb
XT7IVHn7sWPIb5vQUk2UVFwe0lR4793svOkopjDpAiR8KHO8pMROJGrQyK3vtg7f
PFh7PQ9lpolCUsp0lrPnPwfdNfxO2tReboRkF1OoWg/3pxqaRQI7heBRucQweTuA
/Zuzbp36CvOzlWmn7uJAJw0UobA/z+0lDgTaz7JAVThLfpuZUNfNUQZQK5XiUKst
hVd2pN4F8n04D4gx2iCMa766sZ1c4geQQRzGTYPVlFWKB5ocMEgw1EMvrqQbzsBy
1xlKwbPm1JE04hxDuF29DuWIv57BRKE2d72Vo1bJE5eAx3L3pHg/SmvxMOTBBIRC
kGbiW+d3gEoyc1d7Y9Irynai73TFxIF59ayRBvxXRlGhzFcBZikmQeBXWxfM2mIH
yo6xpkfJLqC06ns5SIr2O9aGrFQ/sG/qNMtSsnIuIJzXV2prMj96cnHAeKmtxFGx
NHNm+wl7HwXAcp5UTT2Z7TcmYy6azI4ToOM2DiWFZJjdiyc2CKq5gxHEEeD8l/kJ
g29omTOY2W5Tp9LuG0UBbTc75Zn82Auedf8UJ6E7hidZqXrVDEj52rAaT8i6bzLG
MYA9inxABnN4FU+RhwDuZmdP8e4uQe0dHotWWQlaXTlyxUyV/v4029QoVQSIXCrx
R1w7e1PBYOdvqjGQR51z5COL5Q1mqy8/pztK7jb0M1SphtKH4z+kIPgSyWbh2AqW
IyCW+6N6aHfgee/J4h7B1qUxo+5So6PvokfjWw5Qre1Lud/uQWrLE2nCO7xxfScy
E4VO4EwXfeXUW4yZHzUVlKWgpPd4Ssjtk+CVHndKr3XkD9znRen1MyRFbwCh9edi
oxqZ9WcaZCLPF5iMDZbXGucM0TkyblLvtcb0593WudeWhC0VHNRR+Dpz0vMwKwW8
WENtMJz8qN+nX9zdoQk82FFKjdkxAGfxHnEGcwBuWpIMw7XUKs25AkJn7kLBGtEZ
HniJOoHRGXd5ky/33GMgTBhPUfId4H3QNCFuLJLr0aKEIIIoqCwJ+7FPdyMXSx/L
uVEtxC1IhJ9XNN6s+BhFM+gETsJxXC34EhuRihg9Qgd2pWYVzyeepHEmAUt3OObs
kXHMWvs/uojEXD+5qYMEACeVYVJmyfihf6p8R0UpgNiyjPrLnuWfsHZ+9q9VVZPE
gMPZT4By2LDdFODd1uSMmtKWcxYfrSY4EMekfUCBDQuBHu8DTtakqd8/HcjtMORa
PTYOY8Jb3EKEZenZCDAe61eZixniBsRY3+/pRMz+VFvMs/bU8HVyngMyqLbcMM6A
CEaMa54EinGwNQLzTPaFhPIupS8iR3Lt6R1OdZgTE17gRsFeL3RYEmiwBOAl+pxt
bgzQGUFaCz7ck3SKv4TUfjvf7jOvzdJxiw4hm2zbs+ZBZjCc6l7qowNohw7gEdTX
c6p3dTq88/XhCq3WXxoxmQpYLTCI2v50ee5d79WjrUHFoh+6s3YQPdboyrZxZ2l5
MRIjWNu84X+/8qbldvdzto2yHKPdFxXBK3mwU7J1s+O4x5mzz2wchn2ka9mV8Fqw
XNaD9mvR5U3w4TRJSVbmVzEan9qxS+iSTVoZ26aiJU3jzYpPFYKrVTapzLz88orW
4GrNDK2gSKAMqSLTMZWwjz9BXUHeIChLMmD/8aAMZyVmaAYrZpAHzHtcXkX8Ox7d
EquJ53ImfsFJmabFHVn+SJkpW9SQgsUI/ujGPa4PlqKUFuR1fds7RRyJSaeV6vf6
2mPAh8bzofkasu78+B/lGHKQOCdQ/4vPnkn2/z5qI7LmnMhDXH5EwYetjQAW33Nw
O2VI+dSYUyrXc27GjoSgTAsycEKaLywK0nTQ/+BjGxOU2bGJ39prbbd6XNuRCZyz
5CQBrY12dqu+ztoTsG63dnLZeApwZ2j8rHPjJ5bNd5T6Xj9oNjA3uLXzjVxH2foJ
bRNFnaS4AOf0C8xjf2wIssOR47JJGnhzAdf2uNenL/JzsVUdVPaNjzOGaaj9oMVr
m0Zr+a302Pa9yXDAlSKqZCCs4owX8FNSEYyvlxHKLiV1ISLi42Pwm3PiNchU7OIJ
sLhrQTQObB3fpQcB2MvdaFwE7DWkyEhaqfN3saQG9Y0UOiBzuvxIv86p3cGC4Hrn
DyWmzrZ2OepN3mkS8RLnUT05Qzic1dNjf9u+mcG91QrPYY1jerEjuZrkdhH4cJi4
dsFXQ+qgm0orLXSihMyNmt/HAVBpSg2e6mekMsuNzssJ8H2WdsOZyC9MXUjyGwWu
te5d5XtNadHrmMtbs2NQvjYGq0XOBR/QBalsH2MKtD2JEfuZtt6GZwK3FXGA9uWb
nMTmyjyR1+7q4N2bpYCW3XjV4lvs4c+SJX7a/6/iejNyhP6fsiAYfhznUnklkTOc
C8ivyFOI7qwXio4svlCjDgkLiimMc+0fdUzhJS8BqKYOLtVcMpCTVeSF4Ma6iUup
z7URsxt1oYl23fuxnm1zCrUNM745f5GFOHjv95WDWsgPIaiv4sYkUeMBthoLhTM8
yZF4r0eIrotAC0j+Mh5T4oBZ5Oint20n3fbZduIb3VUahhLQ2uSJ1OVZhCyAf79R
R5hSGpJLWn44K3tm8skLJoCoviPpIXOWhUrIUH9EtsTBBELZlKXRlZuTUTPdVLdD
wn4u2hKI8njw+YeFBYAKWa7gkJs63DqXMeuQmLsiLdZqO1tR3KQpYTHpI/0rqYBM
FeKsBiMkcQFJCCi/PyIQSCqcMJfFdka8GnV/FebwkUZGfVqTixeyRWmrnRlBEa0+
/dtLIEFmAmWQrYebik5wKzXr2EXpp8QHxPtQS+2pPZ/zELg0L7sQN7e9tNeuYBB4
leys6nuGA0PV55Dzj8ufacz/WAAzx0bi8S3Q+iPZAq+zh7U3t3i2vdmXmbOe9vDV
62tLPYGEsWu095MbAj/3EGlHqC9vmNa33+GD7jNoUnHhFBo9a95PuEGN9SKgAe1g
Bh/UeLaH7sml2qYOrAUYILYF23x8lNLw002havMbdWNnCJwqC4Megq8CBpJ8bV1r
96cy2CSEurJ7jvpmKg619I+7nTcOadKGPZtEKeEBpqp9KwXMJ1w5mMHaW768mS6m
DmKRCkZRmXkNbrBEBHZ5vHIqtfuz0948EZqermw38EIldXEqGZKjjKiiJXMOBN3s
ut7eClwbAs+gsEvVnFRMMu+KDhgBa/ieWkHN8lnU9G+oBg5Ra/e1ZilBUkEmleBN
0+1kTknvBapsX5/V2uyPrCxbb5Ee1WkVltK4ivt+bTEc/bO53zoHPxUOkFw0RY8+
7vAvBDI+CsscSDUjnlmhiwVARpdupwcaejxZS5KVnAgN9xRmR7DZFMh60ny3zMRz
/dps5DLcDGFwcGfqIEzCVV3ivYaRcxEOkY8jyOq5Tcl5uWFMcrS2pwbozdGMnLho
Tfe2LW97V+oQyF27PZn6fFz4QXlVxUiRNHTESTCOf5SPTHwjF30NTzOk/6V+2JF0
+o3fOlFPcgWPdFMCYi5WDriQdc9Qud8jcAqtBybUDsIe9WAQHZap2kpUlxSz+QW7
BS2pIew5BCURkR+Bf378ek6e6r3PrvWl0CueiVn4ZqKQpsVFIQs6qcBG8qAtHBp0
NFI5YgGV72VBfrZcllM+DRZSWfjFIcMGZDtXc52B2RhB3iPl1l12//Seb6Lpalfc
kkUqQg6GkkS92Skgy7e9yOmy5hiXjWnTYDPhWNQDJewYvrIfCbre9xDIuU+KCViB
mBtAr3VBkMmNiUdsoqJBfSmKJRyHWJKOPWycRyrGSvX/A0b7SOd4pm1uKjdpG8E5
T4tX1AmCz1oVhmJvTm9SGmF9JmJ/3UQMxobdLm5sN1LQgcYaSULBA2bmyFeny3Tz
GxsmnjUBhnXmfnAyo6x2lM+AK6EybBIW91oOt/QW8MReY91J0qMzyjINmZN6nMLy
qexlcj1ga5P7Q+LkRGVRlF4U4deVNywlBNiTsPryCIBDq8AZn4pT5WDQVRCMbYKL
3pCynHJWNCtzXhyO6IfXwQb9UbMU32KoJoNYlAlc5pCHn8pJ95DGN7L6gOAVlxTj
pj40iHT/VPDYTV99tO3ceVLzkeZI4AJbyaO/0W1wqXTQzce3DVfHhKtK3eJ72DiE
8wC3nVSbwrPVrPnOtcCbAvJiogiDSJy2z7ql7WIKiJymq7lcMOMkfFDbWVmyKNqN
Cz7X1Zb9m3gnxGLHUmpSdP+QNIOpQsh0us013uMh85AaaQkBmYCL2ADu4Awd2sCB
pgbeVmYgTL1KW6hX3LqsyBR6nWXiQctmRAXDVBi16+TrA6lX2uzjNk/1ECCuThJ7
PJV2zuIUNf8sNhvsBKPkMkylLUQod+Ru6lncvsIP1y2PoJ8OBg/4ai4MjJnKg8LE
chraIwomMsJUgV6aC+O0vXJntWcE6NPHuz7QqVT/l2xm0n5xJ/3tCabvBqy1tye1
+nD/0uBksI4zx21Gc4bvHAruAsfECHwXiI+He0c5wjXy6RLWqn3Pw7omwODey2I6
mLHl9bm5mkVsYvXWK3xYCbRWhCb/C+J7ckpM3hLwnRMFh/tq3pkkl03mQdCDlUc4
lcJG2Aq66MGNsKE5D8nng/21fa+gUdd65D4nKQ/FTwMAfHEtxcUH2v1MFrT5ohOW
p35wQOaBI5r/6cX/SLaOf9+5jgepaYCc/u7BNw75jn98XaixrkiNG51Z0IsxEIsj
shyfGSdcyFQz9B+TwO/eh+MNm6OWEwrLkufFdGmhf7kmdnQLVM0XllWQJEGmIukX
CGN0FUVu3iVtpnnjPjw8d4xm8oDVv8QKiyNCto4KN1wsKcYLkWSz99eYBRzwn4/x
9CER6TLQNdFts6vA49kSPm6a/QUlNcMt6joHWPDgNcf1ZCC3oXlQq6BRq1QUCrtc
qGJezT4TyDym58iT2BZp+k1rfv8dUt3menUwzbB/BKeD61XteqFXSo5MmbwnabKo
77Ha0izmaUcDyqp4hCOXdP/t3Oqi8az4sRMI1NOYkb9R12smFxK0aOckw/TO2T6A
bCfNBdncJF5So3Z0TzhHoS8ydT8GPJU7/xSc/zlC8NqAt7aLdFvXeLmaNaR9TYmK
msNIfXr4Yv2VP+k1andRRfcoKnIM7dfiCfAYPoB2c5ISRfRkO4NHd7WOS01j9/9t
Vu7JQ6x3aGokrIJhM5bk5zaC/tuNF1mPNUszPWCUBjO13VaVJOOOOBCn1vD07N6Z
NN52tEF1eDk0PhpGgNo86+D8mFITIuFfA9xdJ0J5Rru/JM6b5jv/NVmL/kU0+2Wv
bQXr9sHPNJr5Cf7IN/jXrSHMQ/VB8YcMry+Iu0921w7rq0t8L2Uhz3YrScVCrY36
+Wei+uiHBEk80OCMxzjWP9RJVFImz+PbImbXEhwqk7tM045NEkcHPitWBYbE/prO
BUWm2rr8UAhnLS0cOcAGoCrQU/bHUtgG7v+9qE+WmnlDGGE5kWueQv3P/3TS9uEF
M2URpfQyy48bPLM1GP5EKJqNkRaXdXyllBoBCAFhOfKwz3Wnx/EYPk4baLX6AMZI
5hAeLwil+goIeHc7QTVIuRF/+VHOZJtqZ+gefJtzKF0+dOP/dPqv82vCAzYZuREM
uFELDBhbjomAvmikotqxtE9qzaA6SmCd++qI+bTLoaK940C6VxN+37G0Gh81vXUx
S3Xul96AqraB/HOvkKlNhOJxMkFy1UOE63zEjZW6jkA9lgmXO+cBap77Jjsp3FlW
B/No6QLaI/VdP+JS7tAo8AFoDB7L5MJ9aqtYOos5FaLHTaY7Uf3x9ebFF1a9mw7N
6YT3LDZzanJqLG0qar/3amf2ZV/ncvUDt3UvC0NVRWPsm5d+4QNe8dt9vS4AfRzb
xUGcA55B9xlJnlOESWbYXMAUS2fBSoH4fZrlSaCX8lIdLgiXGiShqj35sxXCqR+D
ndTYZF6bnRtcsptC5mm44x6AAFdvNBS7c6jD7zaJx4irZWeCS3IS8pTOCblAEhka
KeTAU7hIFAtGY78Ft462Tg06g3Sv7qKnKy8rPw7dkJDxjHiOoMAK1M5CsbanF7jP
Q4vwknGzSh/Nm1oNB47br+6Najax7fIg0LnGWsB9klxEIgvHng0oolIcUwNL0x0z
kzhsSoR6v3ZA+XqvPRGzPK1xeZ1EiEJgGOqBx8iW3TFmPkAdK/YbeB6RMgpDclRE
AQ1OZ8R8ySnWrQFpxB0D09bBF7jkmOt4zw9NeZvXB0yobcfiS7JKyR4kPI3OBGBX
lCMEeNGXBp/Ea8EpCLCrgDPTeL/lK1ZgyIRNClAMGPhPkDVmXptYQWJZ4cGEBheF
TqdrtOFdtJqyztI7kPWwGr6RD4WgLt1OMlVCVY6TcTM/d+BmAx9KzFumGvFgK2Vq
GdjkoXSvrQcKqZk+Drh6RyrwCY7WN5kpx6cK50WjB/wC2FBCJR6iFDGWHJmlLaGi
/9ov4ZO/7hSkK79HmG6KQJP0kL5SOh8OLTy8peDTHmqE6wkMFBc+Uw82tHQObuda
DiiCPHVUl/whIR/OhQAprIM+Wx5ChlZyS3+Qfj6vq/LufSs6yWqI5u1KYdwtTblM
41wrlFuh97JVnq42U4bsMnUQoV67+X8QtNA+kjZXr7JGnmssLukSWB99LvQzrVlp
QctuupGNDcMbsnlPNy7PU9nTdUmdZRgmgDO6+UdzJYBHi0wTWpQp9EgqejgfE1S3
kMLH5ZaeRjtFxj6UZIfLknZreEy7WLzMOAHLqaCdniCp5mUqn48ATFaDfbtjjFsf
wSulgbvHneDQtn6L8r03JOP3kBPn68fpxOMaKbxpdQvUHcV+qq+sBAqjkylGch9W
Oi5dMRbnVAPuiuoV+LWYasUxFGvSehsFnmiUp/Dfv+gUvT9zh6F3WGkpoTctY0VY
wBzh76zBMU/8wSj4QIOCzvOFtbCO8d45c2JXXQ8duSt0JjNpbu1BdYbbfelLocNv
HOOCqz9w1g0A3s64MMfFAZuixNwoSiudtX788fOTid+wt6JZhOII1N1y5LEkTu2E
E9NbTGrAvOstd0XKJVeEUAk7VxJPJW4URtQJqEaaFBB14XMpwYWYv1jzn4C7LRcT
u39Hs7bUYKumsBzrKKVni092hNmPvTxoYN5oJ+y/lnf/9X1kmXGK2xv/wvgcV32k
YigQnd0eqf783I4kuhFMOubqxvvUAJw6b3cR1CKcqafLr16ScE1D7Qfx9ujsa5XP
ivn6pqBE7pg77fPlK046Yu3tywGDDOLZ/pQ9jtNCWl9beOQZgr3uYZCtJBZau8tU
aejg0e1c0Z3upks6KdPU/1b3Z+PM5XYbWe0wvXwJ43Fia+08mzttkbzxxXyfAhau
TrAlEgEHc5w32YCKQlw+UfKpGiRhftHWo2x/2FDNu4xpJq44V7KNxQzfz60mJH7i
wTgsWUG76UU6IHW7MVyZ/y50gbf0WPWSz599t97h6oVBdieEqJsMzaZGe/Yj40QB
62fCUboQolvYskxKS8U7PiQlq0pNKhRf5FKbATq72TNsFuY8RGUk2vIn6yNqju/E
dNBVY2q5Vp1ZMn+KsDK0y03HRHD93faGb+t+cA264JR9nsZL3Pit2XU5jEQrhDjd
ao8Cum5+FM3b6j/b22sXCtz2xCfWFN0wMpUnlq0+FuAlvyNsF8eRAnq0XLRmNOpZ
Ql5dS1+ATJ+g6k1lVTPR6ya9YSFD6NaZphDXnjstoL93AscoDl84zJovw8kLSWa3
i3r18TBb7SEsLnSHObUw6pE+xZFfsl4aWNEGwbXoeYoxAZs160lRG8/X01NTHOWX
scd5/DeoV77MWMGbW8ubn4IDaXUtbp04xIDFpRJPh9IeYGv1ca2941ekJ7MkVVY+
LIimVBJ6s8jeM1UpTZihPLMUfj8gry31l0vkpWvu8Zav2eO+P03lwQ9ohGmlRQNT
5hmIn11GLCrWlZvlmBuYTYV7qJH4Qtq2qVle+gwtUhkrwTAwWmaosbru2gg8UT1h
nWcHidakHSWOtz+A930bf++LfWw6sUzUiu2x2SFSZQirWRe0+vLl6503DBqx031I
xdwX0GFRKvN1qp6xOMTOtWLb2whN5E4rjMTH1motIc/s6tyFQb+gNbvkGaJvbWJP
UZyZR9HBkrQ11Q1+bI5my6uURteGZvz0gIoRkMxIBm4DW2diijbZYBusZyR1v/FH
Mx6v8gzkGixFi/f8xiQd96Scb7doVq3NzAiD0LyZFI8Mans4zoxvKYKKEGCIcWbh
U2pvmnJkYPcRDTkzumcquPFN+IjC5RvIy/07NAPREC3u+PPZJB/2VrfWCnG8W+Lo
c8QLTQaBcqdDQBTyQrFN4fgPdZdZ4w/smuMu6Pwhl9CaBJQg+jWjcXlC47yTumE4
NAPAtHW4vt+7VT6WFs5ZRIJYETI3bkm95a3LLEeiCtWq7hzVEekp1Vxq1bhKPAKj
7a96LsRnIX8cRGsrSyWz/viDNshmr+7lO/gEGeX6AfuObHm202GpSVVbmR8fHT/M
rriiLOkPIZbnTTc0a62I6Jt4DTJQXugXZ96TYydyuxUpP+mpPtHonvgJmd/jBkVg
Q/fVy5pfK73i3s1r8VY0/0/oCu/q6KV8sU1meejluCH6MYa+SKWIFucy8DYnfi/T
GwwLxloUvQpOwej0i3HNHlV5Lsw1CSikaxOTUORPqE65FdgMjCvqUXvMssf5pIOS
S/fOl6GdZXA/SWS3ueHr7YvLh0WnLiK+H7U4vVi/GSo7xxTNiwshOHb2WjtG9+o6
GZaJeFS/dZxzaVfioMHqaYtkMBtrupZ3Z7sbWmO1Zsaw7v/k1aZLV1BnM5o0DZZA
3aLWyC09p4y/gQm072lG6BgjLxyY1rWZ1gawGNk1EPUe66mmBjURftGXMLZCNtyh
6QEK/f/r/MSFu1QpMQRPxT4IAqF2FKnXFK3QlLGZsVALYhE2AhNcu9qxHqOnHwSK
eCdfup+ZxbHHmOE4Gs/XDPD679UZZJvDLx10yAtpzKsMc24aZ8vyCw5IRdE7n7Qe
Sqa4DXvg0njdajO31e9g5isMdjiuCNmuxaWXvzJwC/854qYSnmEtvacQA0k+bjsP
XvNZ9gN2jezaUbyAd8h0+NN8R4vgGXjLxWDfdMf/6xJpPvWXMnOnzZLDA7C1D5xi
NfukICG0C3aHi3NIRR0FWeV1TAq0KUnVcF+vEmubGXhJGTkyZtUXWiYyHZP6ivVH
ZpMy28AW2qKJ2g/T9ZTi+CDEMI+O5PuBLRABgMAobzJ0pRENyyb8TRwDkZKa75qd
9acZo2Bvg+b7p1UtDHhbYF6PLzoW38xOqTdiJ+gRu1uvykyugxhz1POLDkS7o5qj
CFRwP8fptYL8F91xQ5Gihg4uNWlMW3uVF90x3yyoU6+HD/iuGETdoyX1fUzzfScV
4lv2MQZfMsPSXYavx+9An9K2PvSE3v75Ym9X+r5AOZObg0DIuMM2wwogbxQ0TyJk
XXYNoGwYEaKGpZJ7SzVE7SO8jCHIYflV0ZAVPAytwaXnuVVrG4EQVDg1kFDXHZ+X
OBmb6F4irkJGkYPYLdMZGU4hlrbaXRW8bU9wP+Jq+UlRs7pkMXUTuuzSwqrGeHlY
cbM/ObyOEKPvLvoXgSnbasoW5ajyjq+BfIXBuCSj59IhVUqzXPTG1rH1m4vZbFnX
O4xDW1urxceJFve5V3RqUyXa8Nha/3QJcY4EqVZBvJTeZbRkWKJjgQCkBRnK/aKC
DVNOv2+McbHEocHv9Fxg+V7w4Sn8y8FjCgiMFwAUlIIm1pA85NFEypJoO/OxpNm5
i0joaVw+3/dmmVx4vseJcL/T69D/1I/ir5RzQASIe5loJVqaOeqlZTP5VHgvSEyJ
8wQRHkll5jTaHR1W6NQxfk2/2wSHJFF3JLDmCqZMHqYaz4ZS2sH9ulNJDzgqcF2h
K6JCj5T0tLcPjea2OdugMI1JGK3YPbyfWyrljVVsBKnvc+yTMErlO0nFOtBaTBkd
Dpw06MtSBvAxBfz9x1YsadHJJMOohasUllgydATY8O6j781Knr5DYVTGNs2lgAlz
9gSzfRx2M1+GWuGsXE3BJPQB1iJL5LxEIkmPrB1Vgkgic1jaqJ9exyyqdXkFL33H
P5vq9I4hdfl7pKA6jCA/QQwMkkIfK9ky/HrNs35RBnqHBMfd74WMbr+OD0g6+ekH
jVBrAWikQD+dmbcRBu7Sdn4m1qrH9YRghNuioUuADK+jH3Ay8UFU4aSdRjcyfECG
15qwSwdgIeFujAX7j4OwmcfP0e6LUaKU47jKPF6qZLdb0onL3LkcbvF4OZfF0kpz
cqmPe2wkK0kdSBnZrMj6vdycCu32qfcdsOi8mCBDCdMz23Lne2BqGiXViupJWwZ+
GKYPTdcTvnx39jb1YeUXJ8EdMdcWUxAqKXblD+DEpUfHttMx/hRv7hMyBE5f3ebJ
qYM9hTrwD8Q6jlsXPt3vAH/Qxbwj4bl/uy66Wb+TD0FPBPa1lGtoJbUwMPusIIo0
khLH6lI1K2SHVdAW0BWdIyXX3f5nGyilhyUS9CiUPt9MweVkhop8n8Bpp8eOElHM
t31bnG80r6jASHvBy69xuUSHfJz8NjvzBotHpvJm7dsY56CaO73TFTCtM3lASIjY
eZNN2pqLn9zARNG4Y4K6i9osFcJc3HOBXtUA+0018qcP/Wfefm/q3NqzfzDH8VP+
uUxWH8yMHAaLVilRBa3WgqcaDUlu5bDuGXDwKcrI4M94A1UdcFr9k8n7ziHbicTp
Aa7+foq5ASaLU6EN2PUAUGMfmpNMdYKL+KH1j870SWe3C06Nx0Cqk6EAhvya/rwV
LyYLFsmjtYpeqmrUeFj42sUm2nKQtNuSu8eLTkitlGIRqA1Aui8ypgVRVi1+n+Fe
GBRT5LE+I/qkX6H8Ts1tpV0LVP0eoa6vOzz/3H1QGuIXEgTocFDWah2M8Fi89IOr
wId2eSsE37o5jSEnp/dcfdTVEqd5ytt3z3Euv/RtCb4/SusgjXN8XbmaqjQC7fwj
KyuN5ylQruK+3eZENM0AlhBxbyx5A2+W6Rol9JeRIxBA6+LIW5/npwPgB0to2RxU
DIzUMZJz5b745iZMRG+lcdtoVK6VuykixeboFuIKFh0aUocxVzn/XRDhl59kqjQ2
CLQe0zAStiCM3zJIvRSHeD9tp2ed33yFfBLIlc7EQArNEwrT2rzXiHBQcGiD3QiE
XmEoNrhqSUTvZlaW5bdQX81HBOSqAFfnmf1lNPYUXomgk4YJqrUe5leFhmw+pE7y
FBitF/urARC8gOhbrgD5Pb2LbeJ15+ShazInZ+6ATHdZHLBSjY/jEEAdp6gCpjze
dHuhO/sSVdAjz6ah4AGL+YdwufLIFrBUOIXKraUfIT6TRLckseXgBibaG8sKCTZs
DtPFGl+UO51npzRmBMyQ9vXHttoAa4jcOoyWzJjR+rnHr00xNb9DEOwwuKPLT1iF
zDHZBlt8NO/7eeGGdsoz0GfQpEShv5ucNkUjVRr3QgekXmdayFdQcDi3kUMFfGU+
0RiqgkgeGZPNgfpX1ZraHddEySFpd/fzQCFZOAEF+sPbixAD7yABpG83B9qmxDOi
7WlcUNEGIg4xiwZBHroY+EmQsChPn3AzSNsdhSJJxXmOmpAZuLTW+FS/ch0QWaip
sdZbZSxMoNOZ2TfDrIG21j3XawmVSg3wUAM+hzDLdAlfwawyKakmrAzc/4UGefv2
y58VGKz7obE7not0BortMw5rjjIn/AkEzRW1DmsnuuNu74w9+D7ZOYwJp7tSG7LE
kvVO748ZgJWXLcyeWFl0D5Mdo/v3+JsghDtJVrFDtJpRHqGJYvpwc3t/IDiLdp77
RDaK+KbewHV9BZLMIuePvHna6N5IbRvO7h7YGHFPBTmbu3nBSrZHeDwddm98CJsn
y6/GkZdNIyKOlJZAfnsPpIuDoA+nVWDxqAaenMI5dYoZk66JF/oHSSj2RpKYjioG
92fPjt9Xngk8oEs2Ld7+W2nzn6NcRgZkdXL1KeiV6WdRdgYvqVuxH4Ofc0i5chDl
0nThhB1mRKBGTmkJHdiXVVdXFVucd69VZyU/+s1z35Xr3W7QEuFJhH1Ej1mixpT3
MTTnR2Ak/NeS63CTrIbMq603iJL1/9FY9QbViap5KCf+7xHur7UAU9DyVxMeWX9d
f3Khe2hXMojOWfjCNdfxFICLPMF6DtYmyWHAX08vtmPC9l9GLjSkCg85OtnSCBuy
ogRiZgXqoZFqfyT2NQX5tvO++L7A6ffrKuFUnkwQ7AVOR2qMZJpMnESV3BKVYUkG
yA2SQskwMOcUTofLj5HLpk7xEyiFwY5ShU3fTtUwtzCT42sBzsPUmyY+U4sPQ9mo
RYyjFI861pEzMR5OhH3oKsrqmerCvfzHN8xSkedjsHufvDXuZdb9MFXd3ocFZNI5
J/uyyRs/nijvV2CwReKrbY6/N9Bnmzw/IXlYG1yO0qzWDTn8yvjrtXIeAj6DfYoX
LrYjrk3K9Q3fU940GFbDVMoHfKDjaZzNnQyn4K1NdfAKInhtgclcgBkWkK3ZRkES
aJe+OrpMPW/NZo/voT8wTKXi3/bmExmd37e4OHPTZorrrn4AZEbvAjMXi+DtL9tH
tYg9aOPGDWp/8lJ4sQS4wNA5DZmfysfuOigLZpKh0iasOGslFRQjANpxeTpcmZsC
uZdqlJO4+Jd6fVwXRfxpl/wO0ByOOwpjiRJWUl4NaNfrGvgvEh40/jv77nxZT9IQ
iCfvf1RTjpk57rEXPJMB4XWJdhQ2rZuENhtSpGKmA4OwLJlycZaHKOEQKcU3pPVa
7vp0IAtYYJpOPH4gz667BW/649QrR8N+pKiJ7BqhiQd6VMQZrXPRFNjCFusNxuQQ
w+GRZ7sx4xa8vgV3WYD73qgmRNpSU8Obw+VVOPXSr59dNmXwq8tWVaCGlFUPtV0h
znfhWqMgBwTf1pFzjGvAaKHOKGdgnqTP3CiYaOaQdSWpol7iP//U6rr8LHarGbuX
AhgEpc9iAAPLI6Gy0tI2oFoi0lERHkuezL35B/rsdPjUjhhhwJsRUlUm4nQdLQnd
PSOA+XQUj/fxGSBCwy2u1fM90dHiFiSLDm8FvkLV4O2OWBLcjTUAPZohu12NBaHC
gKcS4cOVbMo+tya9fSUwuJPymvonqs3hyCNCdSlUgX0AdVHqDKijClk08PDWn+rl
zWQjxpWoE/Qkuijb8xKIVz8pEQXPcuVZigfKLEwPrnmXh07/8VvgVaf2GeyTgI7X
csgV2dYo2aKiKTPqNGGyK+YjC3mGhY+n91xGvCrUe1ycfXCeesAXt0EdSDibM00K
PSRf9ihFZWi2iCqeaf1ilS5PWHIdZncJSOhoguKthEX8a2BbBHrIO/5802q0iliX
4uTF2V+WiExz4X59ARShM9lOrY8eXMY+RO4E3k0VMYDduq23asu/bvkAtGePtoOy
qjUSgCkqGekDUSjEoZY04ZcIdKCf8IIQZ7rjVrxSzhqkpFsoaTmX4aC8eavy3+1h
Jj1bUeTYqHPdQ83rlse+fGHGBT6YgLsz6wmBFJ4rrGkNcumXgp6gThtxOv2B0R7a
JVH31xQJ4v4RDOuhK74/WQwQdczwxclN0u/PNxvNjUxTYTq7iUg7G5Bf/DaZmkiK
FbkfqOtmwxLYOWKIQskJMXn2w4+bVQG2bzI45GHGbpW3qYIKPVDDogcjY21Diztu
d5vAUW10BI/cVCuKSrlaAxN2uSDdgZvlfryHS7JupdG4D8NLnspXOSBFr1xHjc+U
tS8aUZJTVJR8Wiit6To4Z0CuOuIsi0JU9iY35SllgTBez1JnPEOZrQLyJm1TJyMh
b9UDh154NEmBeLh0Vd37ELt+6EGcofFcgtIQ8H+ymPxLrhKkwMCRI9o3W2l2nuq+
wCCnNmUL25j1/NhAJflE4qT6mUdsUqWtdrnHuzHnOje3Vgpv56Jta7oujh9Ig8B2
6En0QEP+lPczs0N3AbDmOP5wb44xJ/w3yjqbYDqLtaVlPKWh14IJHztOQNx2ncxM
115JAdc0GSPfnB3wttGfGjKqvpKpxk/TILTGtVIY17UJq6BaWYiTSOm3gkADB+JX
Cdu/o2WbmYARTN6uTWZgqwUQhj9EpUqV7d6+Mkiz974ullVkFRL0LfPK+bAiTGFh
fdhfL9lV7jaikkrFXmWDxeO9h1KScEj/YAm7SERPGu6Hm+j7c2s/ye1MGbP+szyT
AFGZzdkwFnoMXkG27UXEB7P7iE3TE6Lzl6m1+L2G0jegIH7MLNjkYPq7toQEta6C
AewK6qWFYnMxwlkVYV03G39jTqNlVoMU+dFbxxaGXWjeZ4O0FvteZF2tbczy1Kf2
hTObpLBt864wWmByGbbd2FH2LzszMx6JUnWn8ISvgwaW9F3hrxkWRjcDsfLrygG6
vCX9IKxWULhYDA700yK5odQToH0kkMeviIvz4k5Ih+JPyCETq2HF71dSFuRqPR+j
g3pQOq8bZkeKWSiNW68/ap1frKKVP4Jkaj7ZinHtePQXhbuWM2AJS8MvBuG0s6NR
nD20zm07HR2AZ5WStu/A3DXYSTPShUAtmR8ww/8rHXzZEgPg6HOjKeZdxv39g+jY
Uu5WMizsFWc8eygGfan996DG8e54NzCv+VT4zrUdyDn0mpJJCb5cwWJyiRLmOYkV
oUBrXJupZdpOAa2X8bM/a6f1M+FDw12AyC6CD0mNYtzK44dZQGPhIOlt3Qrl4Xa7
zx9EBZe6YP1cdk5GGukXgEPNaLaDoG24fdW7kxMxuF8rgBd/n3v/xfHoCFOL+Kqm
w811jfqaLqjuR9efz/sBVPJsg60FgF3gR93NXkbrp8NGqrIaeFCOFoendD7tFczt
c1GxCZY6nlPkfjlYRxTvrbQrP3W7EtO+3AscUOo0d9B9XpB2C2T1mmrMYznVcPa6
Mejc1nhin67/TbskgyVEDxwd2g0iyMIDX+AJxmFjV7BUsDxs35FjQZHUKl/JR1fK
57GJZ13AWSPKLqxCFAUyPmzjHq4LaVDtHCcxu/gecPE4eXeWeyk+x3g30z5uBLhQ
QbLcAYphVjxk0E23GBMZ2KtvYcG9p6bIrOdjwZhb3YccdEcdFkA/auAAcD0oDS/z
0pVjUkj4mSeKzjEkbwSHm8WGNCF3zgQz+UaQkRL2uPo4iIUKTMTZZj3qrnR/72JP
SNrYq79EYYS9Vj6ggxZeH3Z2QKVSZSuNA9BVBo8yU4P+M+urTvkHVXYGiUnKjoR0
8p7q1qz8XapjH8ri4GfKwHa0VSI5YnksFGjGMuYD04xOm9F0y0ToOY4bEwrpumNh
e6McF1ZoQhk33cC1SIrbehxSfVKTJAwWNGGlseC9Jv63YTvvoTtwxwBqxTCu58yx
sTT7wHWqCP5NukpncPEt5tWJgsrhXyeLK1Dh8Y/R5ZtRl64Mh/tdDpOJuSr5U368
q6wf3AFTRnFa9EyH/N3z6pTKfUVay6Q/RjTJ0snA37+1HHDvgg7zaWRQGmZkkZKu
kptGdkYtQTYj9/ASrQmsTcdW7Ip3vqk3UliJ36Ygh8IiR48IbX9/8NVex1WuNjR3
aeA0x+OqFP2OT+/JuyDU7qIiVCn+w4y07uJWqjMf6DPQmBEQJXbburBZRBMgju+r
qV+B1m/VpQi/KilGyse2B/lxyAwtb1Jm3w+3bLMFfVzYows+Grt2pQU9lit72cAi
y0/DgVOCSSB4jtYFaHvpwRaLixD404eUFl+6viblRPjLeBULXD7nkr8nlMPkZvp8
SHmqs6eGY0rjtQ/kMMeIU24RrguOZuN+ICui8xpiJYhMHIGYvDcIjzc8cW/RTYLt
kDi5BJCOrM98ycAMLdFEwuueAbtMl3o4Eec2VwA9sV5n8x3YcXUto2b1YuwZ0jUP
3N69WRty+jhFv8NOFuQQetueHK24hyl3xq3CZel9HouoY8KFJklP94ihKnusI1Tl
wFnuldrBcQ7pUzAqzeA/RReZUy2XKzgTPBl4l1O3NrEFqr0BT7BPxEq5ezJeTum/
2jKh21VmHpOYQ9yI944lj+g9u3ElUsEM7p1dPrQowmhWitRF35v1bh6HmOcoxKS0
EnAUYRJKGfFpu32mNbqXRW/XIKVEY9BX24GU81Ck8413+qusoYtVm4DRG9qLljjT
XbJw83du/SWUUznymP0gX/6wElk5DJOgcfUZ4wQP8YW4h8b1Rcol3sxdnvXDYR8f
EqPA4G9oKxiIIzhkogSWwb5sB/fH4pCdWoxuHqromgzgQZwXf2drP2luxS2jYzDR
Dgg2s3FCYoM2K7eb/YK/0wK0A08OgPwq9bUmjP7M7tF3zcRl5Y7W8W39XEEsYKVU
2OqUMG/db2eiHahBHrb0R+dbTJaCIr684poKlc+ImlM7G+i87m5raDtCNhWSHel7
EzXCL3W9IkKtpy0DLbDdrg86y/Psbva7KAWOOCtigEo3hqC+/oEbbU+CyE1peH3H
Aa6zmIT/3z9Y8JBrZAqzkI7zS/kQArOJyq8NK8VA5ZX379owvUDSG2MGBLc6LpvN
fnJexJ6h9cKv7yTAzSXvVl3W5Y6UkW5QDV9KlNl3rie9ov5I42mofI/dlHCcDNUH
59JxF58ob5wDXsJqWuLys8ozQgUzK0nsMtZWAritd4ylMkAIb7xu7CpcGiSEBWn7
jW/16wyvjMczPU9AuhC/5YA3mugEX6hytrlG3OsxiyY79cOBq0OJ4HkbSvqyd1UZ
4LxtDeGE4eoVwUAfbLT+uBsH+9Xf67dcmKJKAWPafS6Zy9t54J7kSilURMZmYglq
M+QQgUyAaQ6Imgp4sXKV4DSALtaLG22i2HJV8k0BmWMqPbcMlpZN5eHmXGLcQdC/
Fuxf6Nxh21ogR9RStXCk2o/IPCTNdlLrPM9FxAcCqOjmDTnhuyEdaZjiE5z8NcWE
9x2qNtJSoekkeTlGOzYjjryOwrtMGoIlBpnegwA8vEQ4brOQ4GqTjzkOvWoPJ4Al
8zfPvkzKRcWqg7L49PKIPPqp//m3GwJyQQkPLQW3P6IT1wZHkT7t2RpfFEjbxPsF
/fR4QdLxk60bZPL3xXuYkJVJ3xaLGgKWxGLLUOZBBSPosQJQUrXtbyuuZQFvwNgW
9vaqMErv1fTsW6/8BFZe+OjIzD1TUvZZZEnZ2u3823KqcCzIHpM2+Sstxprp/tmx
5gIOlHnecErENfDfzn6jbkxNNROaVwyfQ7tpL4NfNNl7+ps/Bw3n7hezSMYTfy1e
s4AjPCsdSQM7H5ztUAXXUb6Bk+0dBwONpoBiZEGY3L5oq7TmOIpRLIiyxSETmZzH
xHzkBPJ0j2WCjAyKdT+WDUsD35cI/vV8dHnOcy3XYkUq+HRyYbq8E+M4UDUR6Ulo
MqAUaCONaM8u/L3ppSclqI2i69Q5+tdqgy1pTFn9PHzDHV41KOHhTeZNFJqrsy79
7eVa2o1xN23CC+/dg++c1Sk9w89X8FljZsLQfW/qhzO+geXUgAefAwQ3loFxJsB2
z11ZMIa4odnOu4V5vhHds4Q1GtM3G1lmxHHH4Qay5L6Z85fg4GXSsEbDFRJqDNep
ypLir6fYLvkXjCFgfmomeoSzD1pQnxqlasF8uIGqtMzsUFtnDDKPYyLPPD1UWI7P
z6x24l/VtZHT0es7z0JEZOc0APDDJWHakkrO1j8vPNN3xs2DAVlJ4f2fX8TQf5+F
DUoryEdX4zRO4yxuEeb/XG9z6PeJza3Vazr+9l/NbIN6belxEPDivlQ2nx8p5gX/
U9uJDr4cGVQG8jucOMRP1jV8Au0G2ouIgtXyMn4L/k7wNnHD02YQ+a2h12pBEWpN
9PUfn2DY8jw4LjiSeuanQ900I6Fv3Grd1WIR6+23yJSzQVabeNTvzVkaycQbaKv0
r2TLFlsz+qflFGUG/zhnrQGv/GRwKMrFTOcs3Hdc41POL4w/bmvd/OPrpqNnJaue
sRjPEKMPD2yxjBLleZwDi8kiXP8xIPG8PkMrzv0KjJ+OpZXkCyWBSrn8iodU15uq
0Fk9F0akX+bEapvceFzDV2E/L3aM6kAm7rgkpnc7kRIv82WI/6d9T1xKi+mmlcF4
dJDWYwp61QuDFnQ/OyF54EzivNiVKwafoW3kYSipSCkb/Ce/eMIu3eCj7XZ0U8jb
5U8U4rZNTVVw7xjecM0XgjhLjTpsaPlL1GtGuyn5WjOEZ6vZqFFTgbX5lWr1xvZL
nbXjLYwUU9UtfY0j6fQURjojNjO0I525Fm66jhoI1pWEEaqcuORuvdGToQ2SELC/
5Nv3qIP/OU1LNQV9zmijnUatEwEz0GMNPgpMMzjhULybIh5nSOZdAunAQj2U7nta
PR1Hck0xBTmyBQi1Th7cchmFgc/DL+UlyFDOpgxBx2GImUjQKHezR0Pp/m9B7uyb
xfZOHCNUzNF7iSf0L9BeURXAtcAtn1Qru+52LNdlj0cOzxe+8h2VKT0WOTM4q11n
mjFrU1sdRwGqJT+piaamYjX75YCIWcY2OtFa+JgjYs/83fuSiPh+7n/370ed5BYz
yAAHrB1RuLIpPwvX0+fYywpD6CuF27MpJCpBjbWh43PoALu8+YR73+76tcyt4Dyo
r0zrDgHfv+tgxTKWpXKEoF7qmh//dOl/YJvlNEvui4LkWyhHWBK3/ZKEM5FA8798
YYeb6Rvcg+iEspHeEtbCgj/yER+wlTZNs2/Bh88jq9ZshF29+BxEOGIdyVRcuNav
eQMqoK2EzEZtE9K/vbzp3EB1rwsUgqanGN3mznSMXPX3Pq9AqFwvwqgilnRZOe8w
uGD5Wv6M1hv3qVy7+Juw6O/VOS3yDUk8mpwhdLfCndx+Xxud22ePEKrmDgUOY+c3
/huZ06/fTYFZB4pLVoqGA5e1Zs8yAALhJpweZ2WIxl5XFr7+kdW7hStsSkvX3tUl
y++e8/HBK34Kfe1EvnGiZG3412lI7fwZBg7s6IFWpU2ctS2M53kIS+chFLe3J3Vq
D/tj683KCp7Baob76BSEsjbDM6Er1yWlDPmse+Hw7slb5BaDZQ+DconOxImB36K5
OkWuJYEPvZ2/h7Z6uItsn/Drk2MKbKhwoD6LIZsj3tWa3enTPxrWYTSIf7/bWHVC
AzMKOkz1FACRfOSXjlX4Bv7w2cq6IxO5lYiPpMTC0dxSnlcWVgw4cbnMN6mt2p++
nbSBa8lgmV8dxnGmOpKrO6wp85luM5oSy7puhiDEBO6tc65bdXhRV3s5elLvlWco
x4zE0CEXMxDeqK9HOP7KgzqoMgzt+VGiulT9lWq0oCKXUPoUc6OjApiLjO966Zzd
mP6T99Y2dxYFkWU5DWMfI1CT4gv8AG+wmgi75irdOZXpD1ZerPOGmSOdK/e77DZt
QHQaIz/eeuZDWYGz7grzjdYdJZ9szqQNphnSXAU72kh5x6o0Tib9xBhhMOtFM1zK
0GdcLGwJ/ZIUFXjA9f0odlufh/Rt7RDleaj0UAwhyLEMGYzILb0xr1i5jhqKilPK
r6CnaLfS9s5YcYuKNZ+GgzxHQQcQLtqi37cd0Y0GfYu2fbaOP/C11WxEuPdyR1Ot
Z/n7QcBvwc2rEt9mxLUZuPqZE18ncPNb0p38Zy3NgAP+Ve1Ds23QpPk99src+t9W
KxJi3g3kSKyx0vy5c6Q+17qr0H/usxVh5tmMSzwOr/WVCz4U9M1nZvO/hpCXrFEl
djBnFoEHxh/E0Hwr3DQmw0uVyTedq6WiUBQBLO6D4HOelsi8E9A2sOczHzAy6kJ6
XB6p/T8AIGoM1dNs8YGQ3NcKzOQ5EIduk715fd5amDPd6Rujb6UEy13orr/lARop
xV0y/1jewKI0yXbmijpqOjFTGTqYlKPKo4wdqsxxyMVIP+H4DpsC5pP9h7Gnws7x
not9sPbpmA4jGhMlf8CzAB0h2Asfem3TKgqxPzBokw2UgkJYUx4hV7vdzktGRSNP
q01HqxV8u1X4Re+OiByufrGXTIzad//CCFu5u8BGQay/2D2V6a9yHJ7Tp8Jaq/f9
lSgtj/bzV1pLeH5XDKKL+x+r9Yg+BbcXCEpzWFnr0r4nUZKumY7oIeNUN2zlC/br
ARU7m2peWLXfQQd+sxpgLA4jckvW8AJyRAY7yw1ScAKytyASl0aM+PVpC4KvajBO
t59Bzz6MujLHG/wG6u6xEkQR81y87KdGbSSzVQw4lLWm2Ew/0bzmvz2LCUxXo5rC
JtdpBnsI/aVkmq7RROiZ9XkO/ZgdYzfkNZYO3debGGVZcqCzNNH+MaqXQf+PAxBA
GjMaW1NxaYtMtwBWkuHbMepc0UTf3578c5qBhiD6l0qUsME0fkGey2h9eCjerRrM
kuKjNilvwU8iNsGZTequqLuAlvx4ekmANO4uGRpv2ZNAUOBK1kyAQRJgYo44xogw
fNhnvEuAC4ML6p0BdIld6UqH9ZOH+Qlf/JHBJ8U1YOmO4UQbuBS46oUG1VyjwcGm
J9BlBxKGHljFnuQe7HC9h3gLckmt257vlNm2RQFxglS/lhNwx5E8Oy+/WCphMxaD
khAUuAmMsdMapTMFtdGJ7O52UrFiDBiHD6IZJmtZeufpw9h9nM4+Dk4wL4Pgz6tX
4Yoba+8kIj9moBLAPbsdX9B16lX7CpX5SHnIXdUcGHpa9KSLVBQk8mqh6OzyleYI
Kepop3Z9r+fUJXbaDp/bVMNH2QqszyudU8sPbfNwbFTt8UoJlSEDZCsAi9XuFc+1
lZuKNejxbkc7R+v1IM9XBJpfZcDzZSsBAXYECb7+SM366HpdduqS3tid7iiIOt4l
BT7ZFPPfESwpEhh229xv4Spro2oXErlso7l8BpiCvBB6JMSbmHFOiGPOKfcTOIi8
iHMCP7LrGxOfGoCw3KZODZDfB8TYVjvuqwmHEALZhiR8oOJz4HtuSb3aqay2xGqi
D+bIYBarrg7oc5dC/53ynjKWaJG0LIGYlHPChXeuhkN8osdp32riiKDcEVph/wiG
9Eb15BUgWonqA/+O/yHUuBkCpVZq7tLNkxxklquGncpoj+EAUIPt58nZqM3p6Mcg
s+NZzggUP2WH641h/VEI/UIPUm2h/VBMPePmEKwmsaHSKlDfJR4NU2vN1iCxVQah
qAnaCTuKQ/RlJcalW7yJZMJjern8gj46Amc0/P70TwBHv1Mqm/HBhjP0YQlrUq/v
PPmSGmaeTe0PwSvEp8xeDrrm6Vk7KxRJ8K6sCQ+XCnAa7BAMmmX7I2Z0ynKs8AK1
lp3lvlg8YIcjQ0ROxxWSJwyX6UyhAgDqkvKAB6YN1IoYA4fqO7Xju3VxBrGELPZo
4NGFb8ym30lu2gljcXNoSBKHjfKxjrAsHANN1zqV6lDhmQOgRCuWUS6RjqSYcXWt
4yHv1CxZwiYuXHQnmi1G0na9J1Nej8DmUlfdmQDsvUIbU68iDf2uUdECoGPS3rFl
71oFuIMsuwgBgthMcwgkd4Wrb16UpujqD4RGi/CFaLW9L3F5oOM3OkW2BBE17J2c
8H79Q+N0kWYUYo7JV3U8Iw+wNPuDSCaI/SGjx+ANd+S04FAVTnAuo6qdU1Tp2TpS
B8lImTJDCQe3tNxGPhj5hHD2LOue5pQlGRgbsvu+tl1bVGHpJaZXkuGILZi0XkAP
hwVPw19NU5+vQ1TKWnagQJnUifc5dKmX/DjcRA03IGVl5GGNuZQ48L8G/NdRV5w1
VBlvRMwJKGri2E4+QEDZnEj/J6LbWqlVG0slun143bRP8xlOvZN+DD/fXu6Vuhqs
gI6fTQVJUvQEUIwi0miBUQLTz5Y3KjNpm0uRKU7Vcq/6iclA2ecgaXOEvKrRKtsV
O4wrbj5uDBGKRdcVD/I+YuDFBdC8+dLHN6wwPqn9EMVxiap8K/XKolR1p1MEuClu
8Jyivrzwq6rko56sMCoAdqiIX6It6RiaqYgXmJdg1XXi0+Rio3bFV04v3mxQItda
wBVgsyoynrGu/731pT1If6RnY5zQo91VedRtYxMbhFpRdnYBN8EudNbCAnylFeQF
2fe/p+9twZMEQoNtR8lsRCL7pPEeQdeMPIoqd3o1gBosITN7RLs6DYp1NSSDxcB1
rH7AMvMmTH7tatIxeZaYUYDpHjIqwem0YJ/eAOdpSG8x4B+NHcdl9d8yslXaGXk9
MG+lyU9Tt8PKAMfJyJo18Z/lcRu/zXZB8wdJJ8m8BdGJqZpjhVX7T+hAaPStSqlJ
+HAq/+CuvetEA9yxuSZ9rhjRcKii2Ylr6cPHXGkbTLg4A/g6yV7JEoVwDooj5VAd
ELOv+JUi8HupkulrtZuaEN0kOxZiah5ESvbX9wTmPFas/HMmmNFz1/J7qq2/x8je
3wdVmC+YxId9p7kI5JOHvPngpxb8kXQx/xzrpNgGG2QQOPvVIee2b1ZHd7WmzcAN
sb4nGR0LP0/0Oh+dlvmdOiQpGDZstVwQPyv6UdQUpklppt2FAnffyhgyhFFfhPDA
XAeKVbenuNGBRLSsQPTvq2tc/l6r2k1jDDwplDGy3TjqIm97NDSwZMTOCNz7AJ0Q
OFFejFjfVR5Fzmfaz+yIqokIJ0HUJHA52NuoLWsRWYl0Hf0MKsp+YJCfbtgga1pD
WfD73/Y8fyQHixIopLzIANRgAjwklq970RDVFffbwehBvbRrqlU0Y6wvM4GeTSp5
MXqkZ0441lvmceZa3SkeluxFeOiVx7H0XHyxw3But+3LMilYGQTC/WzcZBZI0OF7
VuVb74zgw4M6AEhglUt95qXw7tG6FqqEeuQ+rfYE15rcMwPDbr2AlNIrHlUcIEqO
WTzC0GZWN8tvgT4PsxzJeHcHpLVycDVLWjoWrZRLMVnwrBvQ+O+EEgJdCIT+IryH
zuYLAKWGIaip5Fs8LbMguFg3Nn7NPT39EfbXkqwolrbTMwzarE6pLuU+YIh6Krzq
Y1np0SMUoIImU6Cs/0ryzYID2+13Zrmbx+JofkbE1dqC46omF3jaM9MtgvmN8SW7
H3uru8PKMLEe+wzJj9xc9PbhwZ/loRq0IIegA8CGzqB/o3Kg6g5rwLxe/epVnTBU
J8XBCRf0fMSJrzovNeIVrkDNm2HFsvYuJVM28uzMmjYZH0xspbbATh+z7DAtsuZ7
8Wkox5Csj/uI08x5AMVMhW/faIC+mAykuiX5Se7RIeLyV/kY+dFMoG8EZH3jDJG+
YMPL1+T4h5fvmxvbrslAyNm5xT/yfuRdJEfHyUFW6FqGq+Lfc1VhnHbBQmO/fsVc
0u9iHs3h7evmsVPnTDiOC09/AKTVkNv+zLmMfXyRqcB10lAEt2+dWN4rrLOTn1Em
X1crvdjb50YJcxNFPD56LdMUAZCv3X6so2kFPsZTZWvEqnkgiAJyZP/VcwOkdVJu
XZ2cWj5c3s/gwf54a9HRKzzwIEhhmROC8oFX2JPjTQA8aohtq7PhiuquR07L5sPW
wELrY891kgwNOPHJm167IsyYV6D/4qKR/WYc566XYjtslQdw5+ZTlWIlCJK2RDGc
EGIRqcBP7Em3q9WWKCY3Yw20JdCuylGhMWpRJE1edzUK8nMFBVjGboobdcuTTsGO
8doHmfeCu8IGpfPlpCIAHtQ4Ozkil1BMjAvR5QV8hW1Tune+ry9QCrA/1miH/YMu
6Rer1UB0V8ce05cwiiuiiWOdiEu7+wodHm61lHicT5mupZ3ih+hHbsCKWrLAvEVn
lumApBpP6D88R4qKPw8svd5KqG/ybR/P2TGIDWFYZrxUgILw0MHa9/XNUSJRdfNO
hKs6DNPgPmD6tiE+W2Fip6Tq8MXizoKoe0hMjzgr5mBhyaVF+PMF+C3Obn34YrVS
tnzfxitEqljidME667HNyErIKJiY6pwThSoJQ/BBYQ+sTmhIAeqF1ck8QPydFMB+
SvSg4Do386PKwfleNt5mD3dMK3ZZu3HOluKLd3lwECbHRG4rjYspTGXbRWHJXjDG
8XxsdEDDKx85RKC7BJpcau70BNBdjS1FodajsMZI5kw6x07zq2xGny04cmLZ/13V
kjerG15+Thwmj6Cd9HpwsPyihqtNERcR4n8l1oeZTyLq02mj5Bzx3fkko7054ZKy
YO7RXEjox5spXZFo70CaR1zgpdmvTIupN1RxAl3/+tj0qLH0VMr34bmTvKCNIDy0
XY5uyCRDK+hAw8TEp1pSxGgH63pCxVLJQnoxWEIh+a/x4ffVl+/v8QKwvMKnwqgs
GX2NWo5L8AxI0VEXdStsyhllNaiOF7SaBIhh43T+cLZ0VJHx4N5C6lCYcRovJwnv
t3cCbgqw4n/Ta+Z3Ie4V52Ivk8O8BHcE+bm6YCrITrk+F2QO97ABFBfUm5Q6Hlmr
mnvHZw2NPuQkzGXpgjvHurxDx3TGut2lTTeyF0Atj8Ixv8+0cIiOyTLZvwyPThVK
DRFu+C2/eYOr6GIxJvsbuxOV+hgUA1BJyYyaCDofDhsuKq9Dr/aA4x/Nr+xjvynN
DNXnhVIdFoc7E3fS/S9F9TPJyDmHwZubWVS2oGKFO4P8SpmGB4lnS6qCyG6vhGcR
ji0lWqpO8qncGLCRWIJzQ5e/EK5qCjaQhXJsOeWqtsZR9KIcAhqgcUXld1paa0ig
4aT2qwYJwyZGGQPVzGhcpMywy0jfXh5e+YhiKaBJQlAjOyvbgihqMMRoBXA5DO+o
8I+neQCRlaZOUhTrV494h9Y0ZJTBv4v1/jml0COb5FN2SM0F9kJgrTL4HSvB5wv8
Y3AzRT5VGxIXb0yUdYcYG44nhFldRmlbyF1dh40slOhfEAYLp5kL84K0iJ5CDlVd
5jzcBZnvwU5TsWKL1JFZT9FBFBlcZDEo+dOG4asYToKFs5qSLiMwtxpXpEt63mGy
k8l8QoRkMKFz8gkT8g9Ys6SZSmuK2ofdZdclgCC4CdhwpZZVLLt0WQEZA46Jm8OF
PjCYfi//CTpxBk+bsz/y+A+qeug1jmwr5yd1BUjWg00pgI/rADOxrh2ehaCbDwR1
y3HtSw8If5Y1U3tblf2ZP6J30p4H+5is1LhVCzJ5c/a1Fvi6n45ayUUc5lf/oj2I
zoAXzDTTpvAVs4DXsncQMk8djPkNx64vcCdygI3NzB5GwGlFyXcLP8mb0jotGMHm
gnINrd71c7l6A1xfQPCfnr6PF/hn3JyxH4/L0rTdaZ9kfn2B+zjeOFATQiWQ6x/9
GHpNP0gYhI3EThXzPXq3IVbaDCAZLbFaCj7CwP6y/3Uj9eZv3zOsnSzzCUOapbFr
E/EfNkBpcGAVNpqDDYC3I94P5RwRVs2lXRVNEQDcDnxzmiz2OSDh1boyGSpN7ajF
irkSCN8U/HeCxwQDz5bUVV8HxVzN752deAflxGPtjBOAuFbi9KG+WEwVnlDTYlRx
OMdx+N4ITcDGZXjjKi9+BUzvpcO4h3k/mbR/4EsCRlYZA1ptxk2ZjvQ/pP/S2Bt3
RJ3mrJ08AW/HC0XqXapc8OipDg2h0d0W+/TlzK6cyMGnhMJdUta8GYSer99HCkWR
VvmKVRYDWEMAFHvKhC5P88JACbq3Fpu1CoDpjEMhD8EUVyST7ocrejqA891LwIL9
lH6LK5Cw10Zj28SJzH6wSSKFZBJENQCqzu66q8fQb4G09y/+m+wBTSAjDJCcsyLQ
Bct9CmXdxYrWRL6REdyr3ay2xxbO+VQ2+DcKPfrjeciutdqaa7JUZBQK/6ZAr4yS
Dx7qFwMBFrVsq6CNH9iMTt9d28GvTCw+Dr3tEqZQPEZn0QHGxiEtuxAqZFIXk5hl
wJqldFveMFPKIs6iIqzwHcoCFZgP+shfFQHjjC+1QtWe1VokK1tBESSJjymHXSxh
En4wdVmJYXWBiZPy26AwCLFmbPuT9O4JSvL1kR+fr9HC5olvqh3xbo8gu8tUj2ej
+L2B2aRcjuWUdpZZI+EUUTJ3ikoR7isMqd5bT3v7R0sJU6v7v1GkTnXka/0GxJvM
89PQGNDXgdFM/G9Ghnu7jnke10New1d7O+vUIlLJhe4lJHuayo1z4Am1nZ++VUMu
TuHCwRcZSi857/FizeObUK5T+iilOxyGyX3+06YBGpEXMOiIOb/zyXcFJtErBDiN
qeGaiOgK3dq+9aHLA4Vg/2Hadn/Mo1GPXELIK3bhodwAfKkGCQzhOVhqKBd6W33Z
cq47/EPiD2jKNk+MX4fM75IQ2WILH1rIBA4caL/cl8JScpxerdCUsT0Rxl/kae1+
vx6vwsp0ki5Hdzm/qzFD0BBxjJmk5KWRh13cim9wgEAvttZx6NSM00ZVozHQJP7K
6oRk8Khdaq5KuUJVgHmpfmlRDOWcagXi9lB8x4EgteckBG6N2lB8LTOizF0CFlrA
3RXwk0ZTQx20Z0CmtsNOduKcqO1z1FCI3acR8Q6r/UiLM/HrWX+nPW6Ju9up5v6+
SBgBMAriWttQwxeu9exCeUW02lOYHQHsGwpQaka/bUCLpjM7HHYFKPtk9RKem/hT
pSGOsx0T38EJvCrimsrxiplCq5Q1Hg1dS8fpaVKCEDAkWmaI89dWr47R+uIxLENY
hTOCgNhKehUaBH+/TiesFMutbrw7Mp9S/iFKTPLQyw1uxBOXYsFVQ6kky7eAQ/lV
ZKgS0zbKTZTPhNA43oArw4gwsgKRUGuzSYfab3oCXcB7wtlNb1fV/N3tGXE2k9jJ
WYwaVbnQFhlfRCMMd+c7DK0MmDEx6arU5YTts8VFv4IqFS/TcPMyAGi8IQa8oQai
Qk5ybPqq+hGccIHad9xIEEAMGYcyU1BidZDiWefb8hcCLmqRpSMW7tfwZUiT1Ws5
AyWpMVh5cmWRJVus6I+Nei+ThcCJVJdxgBoZyv4GJ6Z/oB59DsBCE9KV0fdubo0S
7/gwUKQfv7SK6AJyMu1PAOWLejNgSlNgJMRytx70xSfSgMETnTDHaPQg/fgTJC6o
DsQWFO5+Nv34sKX/HqDV/lJL0JPDYdHI6yxMjxhfldl7D+n8mncJn5D3uPAotDAJ
5SmQ6hyiX0rdOpMUatnD28NbmvYmk0QyXxNPEL895g/3U0jJ6XgMkEVFQwWK0gA5
MC3O6GEx302VgFCssk4dLLgfGwhrNdaYmLAu3vdkl1X7b61A94bX4gBZzeFej7v6
N9lccFQMfips4AX15dSUB/RcPmIzTgHJx/ir20kMcV0vfnThtOBEFQ4qqLUXthRR
pbPatG6FbE1pWB+vCMzg2vvUR4b+iLGmzQOhFq1E0LoseEdjU65CqdknFBq/gaqQ
SNKUixu5M8oHnfy4OLbyk3bdIdZQEsvj7cRUuG2EVTAKx8DXOHXSfx/42SUxMFij
8YxsIjw2X1+fwYfUUQSj43+wAiYsrvWi45DcEcqLnNDNmz7FhuWfzeS0jUucPuwK
U7S9xL+OnmWJzuGuuyPQaJSGxobZj2mOpYNu3gKSp5Wddo/JuEmHDLTkWYXWy/4g
aKbcAjKnc8ukPsgh5H3UsA6us9AWsNF4+kqJgUOLVl+zIO/uBz1ml78WPErbA+NG
+VPxMgb2HN0vKKdUwr09U0Pyvw6lkiwJ6Ol/+4C8pg1A7S9zag+vBPPJDHzs6jVK
N9ZqOHfZhqIiVxtPrcdS/YBw85UJzLtKxm6T1kweNntdWkp7KAU841pHApa+H7qK
WdX+nRQC4iere/CxDbH1GaIx9//ChemIPVnrbQBKKwpKn/6up+yCseoB6m6SfY+S
czJ/W+5lIAmzBKnnsjj6fyiclZJFwAScQZU5CvPoQxAhHdS1qVoEecqe9f2CKQMq
w4Ku9YRKFJ4IbpxjNoVE1lciYpJUatXXyLlb1b+7e76uAHz6nXMZgdfmSfxTwNb9
tO/w0c0yYABcM1qTqNULiBbnpmhiRUeLGuXsrLx7cqUI9r7RYfinMA0TkYp4U3w7
289sydnYjRB7BxoNNQWJOIN8HGnD4pYUPhK/jRzPX1zlHOHM6TjF9zTIY2NFaT3c
wn9PkKkwrkuj/WZ8v9N06Ct4ltRgBAnM7j72bD26B4Yn/vGCzLFveqMLVwrkyyHX
UKyvY3l5tsQ4OFfxWJbsCdogO+YSzoTIBCkOCa/o11XgV9T/50W4qqVZCTozQSwf
WZOGglXVo9xpPRd3H71c+ny0NY70KzEVNPAgu76U7TK5vU+0CyKAyep0jkuLQ7N1
+j74yeqXqS9gX5CT9Ri4d4ZQtjKTJfvJaBwxvIdE/ILiE3LQqZHgfM9TwyCfcydJ
rGcrF/Vg8QEcgbvzRMGyldZMJPHmMyTsPcrqWc948w2V+i1UJNpj+gHGlKonaP9o
7aLjSYNzMDjWQfxNcfr6SHgXhgQfRNjjaJsE7zhQuaDfzwF8DKRcFmVrcXnZftCw
jJ/z8dobbAcGITTt3zHK/pEQ4ynH/Cfolgt4p9GddSR0z5SNkFDb6vtpEILsyzrE
3B/Vr/JWzxN3THkziHocidsmmlzV0e+hY7OhXywxn5tZQlC4MGIu4LoBPq2i6W+U
Vpni36HhPud5zDDeptlgREDXs57E3fP72ptLA/JpSg3/ZrmHJLcVCPxi9dWq3qCk
GSBqlP4MRIkcpHLX2mzMqfcASMguMru93cw467AclJ1P6Q2t7B6Qqz6975K8IpDn
DsDxCMlacyf8RPuWRcAu6SV4yhJ01DBSRxLxgbWyKTRo05L+C+1W8u4KXEV2Gges
ztQvK3B+WSriYTrsVauO0Yezd7o8LgaPaDIgAenlqZcixezDHhmORUhqNWtjuqGs
J+yXk8FCdRuUgGAIMLEEF5w1+Pl4rFu26HaCi4JLtzdFPgz+Gd8SljVuMLz/XN21
eqw7U/TXT4+cJLUY65MwezSJQ4jmIr3FYeU2cwDygGW8NJOMKaytrIanQ5zNDc9v
tSdaWe/KMsw6pIFRTUwWe/ZFLQwLzJ+pIWIJMhxM/v1CXeZvdr0tPEkZSvpxKORp
Kzdqd3oFmnr6qwzEuzN12g9HI44cCTu5pbqx5eZrAln6kMnXMNcSKMemyUi1MaWu
m7g/FAu/cOlVfCXEy05zHqYpFohr7iXucsAdGFhUOJ21ODj93VdHacE8miOwI51p
jD8y7fs4EbQj92bai7aj4VMADI+rd/5h+uv7aZ2wAmUgvSbpSj2+hhwaXlnVF6b+
AW5d4KB+HAWvAaGL8KreL9DWa4uWGp36Utvj14ryC6y7Rll53uuyMWNIomWqw/Xv
nw6siO3qG8HYGwRjE+UbUaNdAyHCCKI03MqSKo0euZ4bKu5PCWZZtpshnYI/pv6W
ijTTFnL7r8YvGf4/qOZPQsOpZ6Ob+H6evKwAhMl1XlcaMzvAC4bDdwMAmoZVF6YR
TfGISNwDrIjV5HWXzbwbwlcWXAlHuwc4MeYyydI7l7TyAjjmyBE8upmTjrRrDAFL
6VbtnGCdWdY6VG10sHsUlOl0EM5a1wVDgutn9AUWKEixbLmiuYgrWhyMxwInv23Z
0GAEmCGGWgLihKXKLVTVugjf2A9mJx/uf/hW6voOg8r7bH8Bc7eNnH/SJRkB6j4B
CuI1rY8X+4smv8CK3KZbEILRTt3vOyZU91SQrRH/zyG3dbZYGfZCOGhcwfV048ga
eUiJlkCAmcnc9yKoAaLj3g3x3Q5fUtKhnhhFdnWWfm3UjqRSy8bjNOlOeg0ymMY+
SRXQ3buMgcl3lKGTpRvZ4QD1oGFIWYHyxfh15lYfWVYB9P4vF3QtMc2GYpfysDQm
if+4MQiYp0zU60a3LFEW2/ds47EXALELi4NMlNjmPFiwpRl5vwH7tOcnZ6mi3Wqq
v9YRBnFVSYDxZqZloy+sYfg3uZPc+UH4EP1dphFfBIPGjDYD0l38l8GOAOZQJz5i
z/YbHvhvw6Q/qQTAMWQZv5pRreHWpNDE+GAbNT1TBv0tz4+drATtJ4xwLyASicap
TaWt93BqLgqKG2wzA0KTv+Q27y64kBdqbO19Vr0DZCessXJi18L2M3kPcIxLMTPF
2NGPMInEQ2F1+MusTtdeUDF1vHRFseQabdf1Gmxpem7jTr1SyWCR1AVFzI/TkAlR
plXmRaf1XeGPmJDYAWiDd/FdNl/N/XS1OeNvMN67KIk3JLAbYtRMUR0EWivFnsbn
R5hNvRg0lDWnqRUosvf5f1E78DN/6MnwbFTAFYyPLx5Dhjv3dpiW44L5N0UKVwTF
mcGGM4FpDBI4Cy92uQpy0YXEXjMzAa3JlE9bfDeow0K3m9/oHzOLohANu9TKOGEh
dzWDnbpu0P2Tqz16S4WGEpIZKdp2yQ+tAiBFPyk1U2uNaLiR0Ir5phUT4OqUSevr
m+WsZX8f1IbqZzrC1NihsOZ10RoIokixtx0es7ctulXGpYzVqo5kb3O8lnRZA7IR
nwbjUK99zMBdISaMRtTPeID7Lyo16724VdOb/Gqy4aTGMgTECmHMjucLe0gz+rUZ
h0FPxKGSPzvFmE/jUQUEsvEwqwr0YCPlpksK5mRDmy2Th8pAsSN9NcoU2h4jk4mB
JM9yenhJGa9FU7OXBZpMVI1khqeNsrlgX1KZpJzjApg4qDvHvhppkRfTsbK2Lfk4
tF0lqKBeM+03pWnl8iZikzIGwVBC5IzznOHKFvSZjlA5BDX2McMpatF7CQKleLiP
bhvsjqo0kpNyvTAVDPgfUNQ0Yflj1/K/jFoie44/PKGtn2r8NGLrgKorJGw+HQok
7nEH2NaZZpH+uGxtXr2kJWpTndfaAUmb5AoVba73lMMVMqR1paMJvpX+dKMQouqC
fwlb51k5pCKJNS4v9gnrxvopeJOjhkUGd/+ua0/RB50qf/kumA6yY8/u1I11MRE9
MBIyiQCdfmPoiTbxh0xUOF88f5qa7keRkhNETCmTw/F1CIWF6oVSotlnG4dpqGlW
iTuiHdA+U6PpS9+rhlV7JsDoCf2/TfJ1taOfEwNbjdFtkz2jl7NvSSjbZzcIqx+Y
meyXcCF46RfKA5hCsn0YD+SjjZJjxCde5FULFYxPLxoHpHL+ybtxh4jzJ3Up8XlL
QrQ6XB/ptCTGRsT6Bl71BA41o8621qqJCnNb7FlfgZF5ImRRnWXjoQZEw++ZCItq
aakFwTqtZYtMZEETljzNrcG7wh6HBLtClrnby+KpGtxUUzjCxddyQ4+3iQFV4urG
Y7MDRqoxVMRbF4tPiyOFBeGBO6hGvDUrGWV7RRbxN0fl+6t72FDW+0JrW1Upb0uI
KnZ+CJyA2gmcqaUXvyxeDKtNv6l+klI3hpKuuoydO1tXPy4giiXTLrvg0ZZ15Ovd
vvUMVj7rDU/TN2qd7PpnN329dMp4oY+0C+1//xkgbt4QlmHyWQjdqOC8q2i9zgUb
t/htqFYxii0sTO/WTxhijoQfFBNaKj8l7CLwrX19Vb0FGFti6UV4n/oiVkWEL9w7
++Z5wG3VhlqZI589R2fotVbCCLiY0rvxOdZdtzVVYMA826g22kCn0F8B9zepK7B0
Vb6b/FfBv5ycCavWrpuADlOwYlLYkNhiDn0CeJlvq3PeYVR+DUrUReXXOLqg9D46
NqZ65GkOTAfE/0dPbTEeEmqNmni+88bYQ+jwAJ61rsy44Fpb3DVAvBJeeHSKTlT3
wBQPMCPAQohk3+eS9pYwB/jGhlRAs+vac/aR39HJvTVmn+JvUSKlhUnPCZ9CYROD
eXO/hKc3rDRRH6eilXd2mvGSlT47Z8xyr8Y4/4OJraQE1gEw5y1KqvDv1U6fcm5v
RNmFA6SytOcMQz2PpWNWhSTnQfPwuwthA4d3yQ648X+iB0uMjjo4LomLdGxhZ8ka
yAkzPpmnEa/yBsxydGW9Sz5Q/01UJdAXhEuW9yxSj2ixRaV+yBzqS4jzAT5ZIAOH
S7AiW+wPH2RS3fQW1rg0NUJZuqzmJpG/EczjrsCxj18c5iylToWsUyKOwjesLGJ9
gb1gjNq3ei6ukGIUvOyJ5ebzCIT0oTkXfxKuqEOtJM4nji5k/7xadpJrg4QJMwHD
8OT0SZ/+xprTHAp6kg6S1H16so5w2YqUKB6zumhgsbJjPpCyBuIGNLOC5C6GXWoe
LG+qefAj3zjm7KgRm57QVEJr3wXQb10qv3q6xydNJeG2ysnId0dM0QymSGV9yhh+
IDIRhVHdIAmBFlkZLgw6yvBrUahmjZonpbNNKdWwkjguFjvFht8jHLWSL4WUOQRh
4fwzg2wWxe5PGwdRPL8OhZdLTn5VkLebS3K8dxT1Jj4F1AUmBt8DzfuDQn/oqmW1
IBbjH9Bvu9k6hKP58muJmvQ2m41i2R18NGCTNbOjdLzqjsYIvPjYMS3BhgCpB2Ac
1KLjvymlfqA5i9f30GIzIbjad5ksUoPfAzIObvSRLSxJT0Hmk5BTIJ8vuJvjF016
uriKQoml33uNtmi6fxH1TpHtAW+w5i3BwA02MeCDU6mq9qjR0zM38W0HVxk22TWr
KJa8mHhsKknngoPMoXlDvX6A1xAXfXcLN5MrjhLq7D+L7h+j7mPkgCjIXEwcLD1N
IxGVDeiE90QOofjjqKYEcNLOA3RstLaHO4mn1F5d87Uc/7Bvi8u2w+shABTBouvI
ExL8JDdF//cVToVU2lb0SdRFo9tv0IWppU8E8ogl7P/d2qiNBjwZ7auhKUvvUU+k
/ymvc9Evu/C1hntb91RMtXKQ3Wyed9Bnvqcl8dHfR//lwa8XcWWBJRapYK5l9/kP
1YIRxflZLtuuDGAymP3QcO6LlFa3qPOC4ycJNwzqHluP63bBV/Mf7jyDUIRDG9Y8
FeaJ04sRJi7lEiCBEvU4KLQ1VUrih9+8XTWJasZSdkCqJbp/quqvj074t+gMyBOk
0xWI5wHSML2huil3DSbZ02DHrZHC5wjPqIaTF50EdyBTsMpVW06liDHNCn/5Ysdx
lMuF/cE13nSsgBGhvoRucyOGEAOykgwQNCM7fCJjMLgGa3Sxd3BXMkkV3gf67C7s
s1CoIwalcpT4xWRxBPnF5+VzNoB20FcMRUXw6B0bkxrJgYK6p3KqnwzQNpSxI5WK
Xw2NgBWU5+AeTeK+oYMS/csOvJ1CQ6ruClbVXmBXIs2JdOxsgqeZiBzLetOX9ErK
bwzLabsNzNLTD/xdpFFUu8zTsRQJRoBbEAgt17fusEooAuush5aoA4jYkZxA22zu
bfuSkoTWSw3v2NlypO5Kk7xbE1LPNDX4zmxHSlf3Mbqm92vqXAVm7Rh380ZWj1iu
LufimE8+pj0OI3YGXOVLzGVFteUnI2dQ5D0EUJ4I1Ih9mWRTJkFrSrVG4RdulfG0
rMx21Mw4dK7aLKt/H7YOauNnMpecffrscFw7AUQzElUMRRH1l4mVrI+NM9jFKeGG
I4B7dtgVxIJmQn+1MsH6NoOW8u6u44FvsYND4Rp2xCpIwfe1nVZ1HSZD9qcxK/fU
8X9/SyHK6YSazj+UP0bK5qT1X9EoB76tfFzOZDg87lBDHRSmfKrtFqAvbmLKtQ59
BPkIMZ4dDqCbXLeSkDqdGSx2jQhPKySYQ9N246V7bPQJZh44xQcrLsjvjPVwzkOZ
0QfzcEmEmTMYrxAaY5IRrKVBrl3HgHActwmTW76rXG5zLyV52cg/+AjzxCSHA0wb
y5T+LW3KRhqxODkZ3Sy4XFD/7+I22as7dZjhP9/wF2tMIiBE7rNJfhsoQqrMBlAL
pNYYMwP7XTMnZpr1dn48I8SuiAaEj4kRxa1DEHpPWAUTJ5QWlmE+Vg4wsO3QtL/Q
t2DgFP1SqT9r59hGt5yAaZ1TXBTHPyISdc5JzNZkVZuJJY6O1hJj6PxbEdfn6wHy
3EsU7iv3najYScfah0mujDLP6MEllGEm8GQrKlXGSh2PbuaqKoonuDddx1NSFJfZ
z2fp4WBU04NdVmZXI5+5Z6HYRpCJ+URFTn5Tch6rHo/L3fQcKNKQS+BOnA64dxHj
dE1en6G8vKEP867T5ydMpbGF7Vco6PVc6tX3SKIguVZDOsoyU5M/+dueyggO76DP
0910RhnBVtsPSOLFKtHjhgFYumH9AmYvgtvv0y1BeqnG4fBXnsMOuXid2wYuBieI
A1VwdNDoPC3aLxnjJsQKxwgtxJQ9iJMOr1tiOZyxZ/6OF4SKycUwfK7XH84gZpd6
3BkVNeWh+MRtasR3RTxsVhEbBWSmP2VswwPVF0PhhGm45hgIzXPD8hPAShmG63/h
E6cmigYDbr7ZvTkzdLq08RT/cEZ6oeej8edSRjZCJNQdAx5zH7gWAwbU9ROjEC9J
3PalFvTbKarrZTzY8Fvvjd34sSg6Z85KK+ah7mSGV8fak0p71uN/zvCyRtU+8Y6u
7Z/UaWGPuZiJzUySFJxSwp62yJLXX6jZ6PIcWGRlrQv9lyPaUrx4T9sOtbyhW4MY
Ea6UrT/9+YJSBbNwN7Kjht0R0ovJ55xExLFFXG73+7J1Z0v/1TJNtLPLg56FNp8D
Gi9u/AFA69txML7lsiRP/6VbVXXqv565yLadFM2tBga4QjRz0AIdHTXO2WCc/nYx
R2P+l0FPwtdaYtKyrbSxfgkQNJE+T5QpfoGJ2px2vvbfv8+ZVxU0ID6zbIdt49nq
LE+9HWcI10luX7F92KNsD1rCl1htIwJ+1r2tnHfeZQbJ1H5ii/Bu+GHrVUQEWbQx
nZW0yGSNaQtUmt1MZkzYn08iApKmUqcsjZaBS9XVDcR4gZ9ZEhWyRW3IuqZ05Seu
sB2Hl9L3b9HscjIfrd+WYDtII0XkNX2uxfXBOWwU1s8Xg+trne6JXkylnJ2ZVf4E
Ugacj2YANuVwNMHnmNwLLffJ4txGX/Z8mYxx3igC4iwPYuejryquUilscofTArFg
JdkxOeG1EDgMCUBPtvRxtLkXAOWvP5XudQ4nERpYAVtweiANg/sjVf5i+LllZd82
EZT7vhCS1Yu4q1mOCmMNHoNE09FTPIDOIs9EH5Zbg8ZqvWf6w1aaYMmriiJZuwoX
ljsE++FqWyE8vcdq7s9iYoCRqOzCzlWD0kb4c1pnO33jzt8IzAMpsIdMKn9J7WUN
ZKKAJGpy8U8b3KSD7QncCyHZ1Bc7ZUbSfefG20J9QinISTCF3QtVgN009nRaj5SA
eqfjKK2SaEFDfljFu0aLq8MaxfGAR1LVHZ5qyiNOiHscJdni+sBL6rE7UPvlyhx1
qdJIxQxlX5EJisPOC+GmiQq8sCqOB9msX6TrB+SAWiGJuXxO9EF+WmJ7Crn62jRy
MCtDk/UZy8OpAy7o5gaclvUcwJcmiRx3ttwpjDl5qkn6NWa9N+UaEf2mWkHqTvE+
zK03akhPpMOCa1HatMVzb9Lf6JzPmOzA6Y9JG2hutYgfnN8HO/K1mh8z4mbeajt6
hcU/MX91E2G42XZ2h7rrRqq2guM5dHxUX+B3z7xs97dr3VRw86gJu+x9eF2fhs7V
6lJ+uCtFCk8o3j5Z6tLgG98MHWm3b1SGSIlL2RvOf0SPN5EfosWCpn3tJ58b6JJz
MOwEWKEKajXdSzEvnf34BU+E4vSqb/qhJxZxt0bS6nwPPgEohBiesPP8dlu4uM3l
1/xPxd9zx5M6u9zCZWhuPgagxmu8dCnx0/csdMlkKVD4HiV7u3+Ytmz5lMmmDhWX
7iifh9QoKQRD58/9DNcS5lOk3r94fj8p245JlpAMY3sD7pd0/R+e7PM+gr+evFIN
itVBCzaFZFDbRJbQ55K7ooh9rZtx15UmSx50yA51XfjCbS2puBKqwZ7tOl72AUFk
/m7DrONiBinPOFZppyti2Q+ZX2hT4gB7RDs5okF5XnQDFlGXrgoaBSVwmRAZG2pq
tffv0xbab7nev4DnkR9rgh8al6oSvwUE1sMi+9TMkFfQTUT+CjA4xffMimqSGIKT
3jjejZhts2TCYPmNWIUkahjKypWClLRD3lzGTEhcN+hytzoV5zQFV1VkVNky4AdX
J0e/sk6YKDEr8iN1GiK3JbPV30ojO4kOkYd/rAkPGQK7KUWWZxalQefWxEv8QDvq
GciMDpjDX0u6hPRUwKbZ+aT6nxYbQG62keW08etNhRiYjZHXtjZ2aLmbvjj8WPcT
XDCUW3YgSV4ff/5P7+FqA5wg9JdEi7dqKhj1EPh/AKbOneOsbfdEwYcYu95Fjg6s
kqAp/DjJdpITsp/rjGrG58F5I8NfPQ7U34i4KjUrFeybgYhyOSnbjYqDGNy/hEUJ
CxOkRURGkxMo5tuPGqCmvb8TETDNgOPAZYunmrPNV9zts28xNkKHZs9fqLtC9p/f
Qe1sf8jHmddQNnQM5tgN+UoyCbwoAG9JdcdYC/kdUmM14yylHVxteAqVWnmCOOy2
7L3zC+gt5Uh3DVyxn0Ny5k7t4R/+/MuSh8AIg+61+GjUz5UKTmZAlHlfQCG0TFiK
a+3+EgB8UZIkYJJ2Zi3fN12pf3WGtUTeyZlp9ozIH4MvQchHdImSR0XEToG18HSA
TF9SYuNaLcgF3QKwa4c5d04cNKourbTAsh0F1QU3tORq9NHoKYs95s+u38pcxCy5
8S1unB0LG7yJHMAwPmtQ8syWXKcjok2JRTe1r3VaBaJRZvH4ULqr9SFQ5mL3fPLr
26MuMnHPIZfPovxWcjPPGT24GLVi3fh+1QAEyTwYDlXgsL1yrQF4MdmJlVX+RqZK
7h2CccwdahQdtcCh6XAh23M5TOhgcWhYTe5FkbY1l0tJeFqSh4Us9BuX2SjMqPxC
fdmIbdSwsWOAP3MVK45lUf03U/N6Zem+YigLjVVhSOXor0QcZ3Uwu+vINk9nD3LL
MX8gQIQs9CmZUTDFrdf6uy0buFnKIcOfXFRynd/WvKblCdlfK8MWGTxuhYl+6Uam
YyQaAc6ch4/w8IYM6/pWwGDK6U7P/QdYspNHVyIy9nI903EoSa5eQ6aATT3o5Yf5
RzimzDrdDb21KNTc6YcWK7UkqF+oLSpISpG9Pvb1oXrTkbkSoITFUXgEUpPWMYMO
vFDovaJcKdoRubMJLj1W1G4i508kH08D30Q338tqkCWXOrOhFdOOTUmNJvg+U/rK
SIXi0cLMJ7Igy6gX/At12Nykzp+qXsnFF1PRKQRtjo51etz7fBg+mxo9XRTTbJOo
Ogr17C+13pV9CdfqmVw8m0xb7e8xvvtFSWgVcshxij7CQqAh3uW8I+Qj76Z9XWWt
Wvs5jibUfITuFFAXKpB69nac/NhUN6eIPPCuhyQDS/Gi5z+NxmpLGu6iGO45I2Fn
+XTcDsdqlsNtQ4A0B/cSlF/gOBAMeXnyjCbD0OPwdLUjG6NrYj/dd+ji8PVCS/QV
mLNTR+zobNZMaPpLN/2ws661eBqFdWmduftJJkhBMgpnjFal62IwYOwdjFjo6oy4
lcG5/4QyV3PWdlZB/l7OWUoT82RWiMbVGoOPPZEMahJxedjQ6Z7HDm61Un04nyr2
f6e6SkBLiYrkf7LSiuLy+Tn5u+M6xvKnisKpcxRA0mJu6GGsasXg4rcrrTggPetJ
09/dJr/d1r5el8RfJoEerVNVofvWdT6NmA+sSyx4hxdi6xaVxziU5NekS+f8fikw
sRgbR1rsOfej89SMof8iWj7ilu5r8dllRzWuz3OnVLZDM7wvpX9N6fVqP+oo7pZI
1Itjac3zDSuejD6UKOCb3LkbXOnWuHA/sbgNTpn4y5/dQsZarIo4ERy/TgvTrWGx
k3QJxjutcyrkZMoaAn2xSBZ2bLleomNEpW3C7lTZhgkDkPH0flgSbEvpns7zfOYr
+VRrz7Y04UOf7QxwbN2pv4BpmDPwtsQXd3prfrExD1SOI+QK+uHU2gJwCnt7AWxM
DvoaQb74TXTmSl0xOFlv8iOYWftBTICAiJyZG61NAzqS8UsvUO6vd77D5Nl0NAHA
1YueqTZT2DoN407C1krqu5SSf2sakcTY1a3m1yd/AxaPXrl71ToDJLZ0zsYS31Uu
41+gZYDvEQSLIazAirBV2OglEG2BfuMUrlAmN3MFTZNVs9rQe+zXWP0m4NP4cnlB
9yzYYkrFbcFVJ9wGR3aQHxVhqkhxRobLXqn/sUcSRKROWr4EW41GhO7TiNGXugZ0
049I7xR2xUPRfHa3w+3AJYU2tWThHx+TBTJva3HFXRGDWXQlh9cgUOhpS/QBRHiE
3sGe8LpSb6R29WVeZvZlyzK7gm/1msjkSxpVT+6qEW3iwTl9bkebAjEx/OBHboW8
Jqysu1+Ym+jdVRdPppD/hAjiK2A3eAQQobh4q4SZ/eijLT9cNsXufotOhlRMXp7o
obRm4nY/szGeMoKIfs4D01TC2T7/f7ZyDR4Lg9UnJ7P5GmRG+blNp4xrjy8K7xtI
pn9LCirWZl1ItENH4u4raJn89qRNfop/FeP+3005rVVyFv92/x6rIswqDJtMAt4u
TFtOAB1rjSELm3JKCsk56HDiy46BOnkfqSCz0SkG/9gAtewXIXXwlvoEEExfLddl
IG7c+fX3/y9LXEFjyiSRChgIEC/nN1t2a0n12qwFQs0NYmRPYbOL8htWw5o2S8/9
fkauL2kKzwwKCOz9tVoQGPSXR9/aks0T+pakelKNidQi/MUvCxQu9ZtjJW6VCcN6
nPjNaYpkTS6SHVG4rLIlj1cm893Ta50HvIHXl0kdC8+2/T4x3msLhPR0krRAQzK/
EeMH6lw9Sa4ELTy/zlz7t/poxln0TBYTcsqQPyQNutTeafTOGdFAwuV2SC3VRncn
V5Ra99DKsKqrgEn5fxLkDncUiYl4h9aPjd0m3cWZVd1wnDH0Jsz7++UaUstXstyZ
jyt+e8DJL68l6zryWCq6PWW5cafzYNQn48hBbppTDtley1u+hlTxwtHki/1hofQn
duaDkrPVTjpJZ0ym0p1jIbGo7ZBBTZe1MccT9H+CJp8km+36VtQi3NKAEqdhWtRD
gX5Vg6g3CQ9DBQQbgO6Di6gcdDziVHyqyCHgFb29HZe8vN/5+2pEi5y1Qvm2z39E
2m8SMgicEP4MIKXguPkOo7sNrMBCv9NEl9+NsNSE126nVZprP9z+LnadcqQ0E+Ls
/TBzCXvtbcCyHooud/kwJQ1lh//iRPedd7SKlVAz/07wyB9mF2B0vT+2pRQpLT8o
yapp9XkAoeCUvi9hj6L+snZB2MNvgbVSBQ7wnQRF+qVDYxtzAnZWmV1V69Mxqcks
IcR/I+nWvhyxj10tCK9Ub6B1zMDXNWgOL9AGEguLck988CvEg+1/xdGdqqfJnZ41
MgByzZsFtjrXxtMNu+tD4crBqMLrkzudaFVLdpx5sNQ3x3wfw/H2w9HWc9ND+3ug
TgXWUgsTBL20l0AQ9Dn5M6DEfTE5cIrhBM0Jr47rf133nN2yACrKfSMkc0S1ZtQ9
Dglg0X0uI85LA83+LEGDOJMjEqEUU9qL4EXWNy/t2RCQIJ5L5XpP6HHKaTD9YSh2
iVFB1/x/cwbP8afwvzvKB+sfU3ZDtQsk2mGLdubHcdwYhUbF89RAlqrKJIYaXXi6
P96TxpHgw3g+KJYVa20/radw2Zkete1vOj20f4ZeVHFUiIM8fBUWsfD8GI78FBna
nq+uJOvhxf8av0JiFPen0zawf1kJdgEnndihLGclcb2Ewzaa2WT8d1+oCT73KnIH
FVHwbCwChGqY3FE9n7/FjEDeYha5qCRoDpCknUUL0JG3zAgzK7SJBhieQfN0Tn3V
BfVmHCPCOVEoxV7i79YON8YveYlIQV3SVxe0BqUBNEyfS7Kt59WFViH6mb/vhji1
zKhbSyH+O6sjFaE0Qf6ZqevTsoGucW11HWV3YeQPg535yzctwQHMJ96/NBRmzV3t
V8sTG4lfQIZdYZA+srUN0YRbEu+HAO/w1wYRE9DOXo3L7wYVaI3j6O8Gi2fsDfag
dnMw+YNfBgQOjT3Fp8URdEcz2LLUB2z85AvEfr5265qddhGZefAk4EIHDrpsDW8H
DM8ARc2POgnatuPMU8pRWwNYEFdPFIAGW+1QQc5TxI9i8BP4bwhpHvEQ5+A9MAWU
PRWkM6yTEt9sLkCQj9on08AVxAR+8N4IjcfgTDwT/X4xZiRr3HoO8TGcOwbOwZx9
cU0UlpxR2SG3ecXKfNt39FHXhtSftxdURFsJNJMB+vWClPri8sN5aTIwZ6pIZdJX
bOCxX+XV3eMnLUda+j73PG2dBELwJoqyXwLAoafdI9Dme3279d3n/P7eJCeNVy1/
UK+D4KJgqZYAFPiMm4xT7xjhdoFRu1WC9WAWXYRqnp/eE8+dSdm8SbcsQSwGIfCe
x7WniWf68dUWjSny5MY7dfs7H1nwwvQcL0/ioSKwSLHMN579YP/l/q6pDAnAJkxx
rFln5Az1sxOxwHCh5UA3F7XjwUIFenwqFfglMYnmwPurmzY4lfzkNlvyuVIZSDGB
CQq45wrnNTuI/fskW3x7RLyyEfMWW6U3b90yMx7Oa23Zcqk45h4Cvaxb1JP/Zz2M
JrEbqhH+rOREitP3XS+Woyl/1OdOeQ9dhq6vImzeL1uTS+KeRbqMD0AdnDGt3l1+
Lvb4BrcVYFkpLc4njjXpKdNeFlTd+PMz5P2KjewSPGCFdxElvuaeT5wxAeatHK/g
IL0QYEP/VYbZfmsK37234W17ITIJlQ6BDuxucR4oz9zwKNAwimS5xKLxJ9ZYMJFJ
IrEwzZZ28bvsSwzTgEAeSObPpoldYL+KnB4ZMs1vW87ag6ZXT/uTAScpUC4fYftb
E3fH8bdG1uoP6Z4+y1t8c8c0MyswZpaFMaF7uoVm4EsBKDM8W9ao5hKPB8qGrVw/
J/81uGSQXJRgZ7lJlESaxQltnzmrab4yqBnnoGYW9/G3RwUGYNPrPDUIFwMkQ10W
T1mvneoB2hdqMRexWU78B+anp+kP1xKvPev4stz13EPHWRKFGoBfjNd+OP4bqN/K
wxG47ptUgP+fGCBVYHnorNO/ctLDZf3YYD/r+FEWiVD57YRTFeAnENpY5HORveR+
Lxq5+2nMdqLw89n6hzuw+p2P3TQ2IECIwJ72KWgEo4zrDFnrTZFnW9OeBctqtgfD
FBxjTJGBcXggnR3GNCzPtmMbCKQRlTVRFR8PjHgshr9g07KUBgN/SrYS3wNoqybj
TWIVCplp/fwFPygvqwtDmQaaLy08/eGpSpAZBrUN/dYxUmZAV0BL/uVrQluvqfEa
5QEsXWEWOvrXupWy/W3EjvVYumOHc79ZAbiWxx3Re8prrmU+p3rbbe3JC+X7jxr4
rDgN2aw01n3s0XSWqp8jIN9StU6c9E5rJ27fk/HySsnUBVjYJyUXZmboYFUEygfU
CYL9BfayKmJq2qLzY4QVmDUdqcpu1kDuAUpgQWNKEZ/5j7gWzZruZmKKlbCup5ui
Vpd2RzJBXwbIdD3oGXCnRk298eBjzmuuPl34vDE0UB952iGhgitkiBd47XjOqLik
MTdGJhjA33TWEi5EMw5LaaSxE94Kt1cfWznMvbN5jiCPqmoAQwDxDs3e6TbTa5cg
TBBi4LXh0WALj1cEc6o3uzRhzLL9pYyNf8sbJUkTh9otXinm6m4nuoljzwUzlw5j
FiBOvOX5xXBd8BQKcFVWbLjXQxQuEHOOZKLz49hwqsAfoTCPcJbJQ1niYLVShTiB
hriAMkueUprUNoTtTDEdCRIuiUTj86pUx0jouPZqbsUWF3tgZWM/21OeVY8+CTAe
gSGZhEgfK8eyPniE2nnHf36hfRKeOky0OQN421SBlq7vZblTKRPV6x3o773rHTcD
5lJ1ITgTWNQ5xWrTIiatoAnThz2BpRWJt2HhGSiTqV4wuyAqm9Y8+nu7+EehtfVU
zHBd//B/9jgRu8lm1gGjrUTSZ8pfyq08LM9z0fP4mhSf1k9FSS+9WYfwHm5S+GNa
c0Y7zyAXM4on01lrZ+jucX6tprLEmjSgblBkSij6pF0ksM7QH0Id9wyV2ELKC2GQ
UWGEAZfsPNEumVxPSi0CueYM/wCtRReZx6nfdJMlxpPQhcORid1uGv/CtVssTodG
JkkZr7MaKLNp3VylNrnJoHI748qM2vA0qz2T1AVz++4PfMiEIZP9rE2YQTblWk7e
Ifnewhm1dJPj+NQU2tEoUELTxW06Fg+8XM0VrlAUoOLoIE2JBTGN7GLcGoBYZv71
vKBWKtFrLrXRcjBIFT3N/5iLs7UokaFBEtLPrpBxHpPGQsdwmrft6b9eAcR0qyu9
pgCmvIi6ALRMjf9aRts0+PPIMhoEjazGQsYHyBHL9tVXVm5UUgCfxTTR2acIisEi
gyk1biYvzeZbvTvKMMt+ZVvqflVxWdDSDrqOz8DJ0eYP99rMIFUdOGvVFK4sj/dM
+Ayzsjx1iIV1hDQAy/mDo/rDFrlsfGicMWbpKQWWEeFNQ86ha6abzM5v5NOKVdMf
V26+YQT1ZEsnsS8/p0Um60YP22pxUdd6JbHDzJudgbQDDkZJLg5x0az/wVgL5ZAp
A6kpzZW0iaHa+jn7BBhcUYNQud1U68wBnzCobQYjNNKpNMxOKVe0sdG9HIiHyRSA
uh1T169ROiqzIbhO2x//lJS8SoufSz5ZLJWOrwDoc5Wj8UWM9cIsTPO/O5uylPmc
FPJTfWI/TJvNrCVkQKe3Gw+DHBHDjnNl2ctp2m8v24C3XJBMi5jqUGFisIFrEy+O
X7WWR2iJZlXUWawSdqwUOrOWh3iScLt3YaJnY54Jb9dbgi6mJ0IKUXp1NYJuv1rH
VsdLd6GtsvI8I1OH8/JVQf7hDNln7Daq8exdwGfgGX+Ai6Xaw1nCeISMFa+jzX6D
gsBugG/rAnKNk8jnKTyP/DpTfiyNm+cNYorv0rtlwzi59JN4BQvep0SChBp7Y31d
D4Izzh4fxHw8ZJjyvVbiQsjvd7SBsE+M7q8OH5RapHI4fkCqaGxK//60sKF57p+u
F1at1p1e6TUEPUkaeX7Ue224zczyMg0IVo+/jVCCzrVLYrtE+jU8VezH2STw28Ac
CLZfnvYRtVhKhHpdxO0rnDC5YFv/QoMdNHWyzEwOcWVe+EfPJVF6JqDrpWCvmAAr
Iy7mWlNyvogpTHrmhmAlgcODEjemqeDDFjaXJq3Mc47tTEuLEcK+qyhg6Sj/Kq4R
FxcJ3Dw3FG9U2bnEd1ofxyEi4BsDLy6ocMYPUAtn3hBRrt+CMLpWnRXHRfIURe9S
nJh50JX7hO2l57CwsuZPKKlTZ1L9vDrqYhkGG3lCRhx3paGQ1AgdyDBGPG5XUilK
ztTysy2kSM0563CdpjvnSrt7PCtiTF/J5n+PltDNz9BFv09lYsc8JCDk3ddbUcGf
5UrpQJVIIf7X/H9XpUA3f7OBBC0RTvs1wuRIkoT8VcH+ivjlxurmegqzTqmPJFOa
mpOoEbEGqfnUdjkGzpe26kCLvW1aKrfeoh1/VDpv9/6Kbqj0wBJL4mfhcRYbGMjy
2dajm5r47RcbSx+1sHBR+9Klk0rt7qLusT9urv8JxqU9C38xNm8jZnYCUJj6jYh7
Ilp6B7QevdHScXnMGrl5bGfJA1tPzM3cOthkKJaiUHtQuE1Fk4lJwjuYbC911Fj4
hc2uVUc7jF8Vond7wp1mUx/l/WVeuQDXiPsL0MzsaAWJsGXox9HwUx2OXE5o+RTA
gDmbZCfbzmAHUTs1yUhUQEQO7ytoltbq8lesPBdvmmLrgQUMs9HmSjKX3GdjCxzh
myHbzIDmJfrqYI6/JYruhjah9aycYadZzSKcI2cwSjh2O47HoRzVVexC5fYnr8da
i/jDp47Qxr6rfdkWIFLATBj1eDs6LBEdJrQDtFB+beVmmzbpGkbrleGOTjfjfcTn
9smNojCsDqGIM+I6smveMYqCM6CoLCDGz6NtjT9AN389YHMRAYB68G+fbNLBRprf
elyV3zrEVtmlSnJwEkf+KGluQNdv2jynMRa9aaeE0I3X9DDYu5elURpUy5hEtq5K
sdO4vCqX+bLYGFWtrlrngDAn0+l3vpIJmKP02BL32XqUQvWaGsGjcwTQsvZcwWNa
2bU9Dv4MSM2/mKAO0ZXQAn5G7CX0jyPyDrbTC7IZkrpXVK/nA4fVbh2IiWbGh3+V
7Bl7ARdFl04zP0fQ+HdCUZ77xgrg+K/PUw0MsEveJkf5TAuXJk1IM1HRSsur7hLS
o0YGymIvMVhSPokvcUdzWCWHbat67PKnfEjyzTAEtM6nJkfQLEw6fVTAl3QT7qkQ
9m69Qsa4zx5yklUyPeJFXxQvqkUQZKNl4yKuorhNQLd3BIueEy/TcSlycEmBWjst
qNd81oWgfN3WCDyPHmriEP33Hk/eLjMtXpXr+aU3OvwccCSZ+/U8/VAxwDxz5ZQ3
Aye2vg32ZGSmXBdQbYXmHC/4Tm3WvcwksyNUIEJEailLkIY1ZKPIh1Rng1srp4of
Vbc3Q1k7OGu2i2/fuyQEsIrOapSjrXRpp244jvzzo4piacfNjBlnHmwMZCkzpGUr
Synq8ueCrMlw07JvqOaNme7btTvpGo4gEaWp0yXeJElsTgKvGvi+TxptVho8Z9YG
dgKP5Sa8U/b8ZdsYf8E2EkXCuJt1b00HqLDYCrBMg8/MBN9utwzugNpPy7bX/H3z
mXjUnsE7zDh52aMIN/4xvc/khrS0iz+IBCZkc+jXjvEM5VGkOdYmSZYnUScCMrcj
tPIj14fNHMoVsrXgidmFLr6fMFmncX36RlmjtKaasFh9AjsD4ian0CVHFwABDDpW
GqJM1NZYghgBdXx9tff8RQN9LkK57k1kfZSxT0Dx4rt4ee5zy6YhmDHM7nxg5Q/4
fcCAEzkvmXQNGnt1a68KuNtxL18Odpn89IQU6VB1QNdHEFKleOlKkkaL8g9A2Kj+
BuIpCNai5EkdhYW2Jk/vTJJHB3BNbhmJsk90YSvlwrqO99NIUWpZplmGy/utRkxM
nQCm8swUhPBzCC619i2a9TRmfKC6x1bZbrY4p2Q7LbTtaPbCG7hG11T+YoS8i7/A
KiLTv0iD0cpxyAhQuyGcvHznfptRM51X51vWaW0ZBTxcSlHJ9IFKy+lxdUdFmzX6
pRS8uWaUrQ9LbqmOTmQDB4aLzwxVYiRI0OoGttK6Yx8QoCxzrPqJt6IFUi471dX4
wy4YMvT/1CnICZgeZxZlAGhgzYg9SKDCpjEFmO9O3vwCnAAhJggVSeh/MSDRw0Tk
trLZQEDkaPck+Ezr7S/wR8SgauUJK/MLzIYEI2DcensCLQVC0LXPFAEcrqTfl82f
Ao2ZpqRAc2owRSmK2XT9zMA0XS00P8zf+frb+YBfkqSusjRWqUIBu/Jr+E7c0C1q
LXazfDhgpbxHoTy6CDJVqLJ+hitCSA6e/86q2EA1ywAaAwxKKo9w7MOHR7e9l63/
2Szf7esg71SY0afNZ+MkazlyUjyTySvOlEO2PIt/01hS2HjlQx/CWB/cNkO9FW4R
FcfdCYQcTRcgIDDvCHeF9JXLndSVOYKAmJVYa7ASGWkrN01BQxL9vpvL/xEsjIQD
0dmCAq7xTIPY1rBlOs2tS8x1Joc9jZ3XEjAQeCTnLyGW7A6yvT+VTTPuUNKdM055
CttZfCZ7sQP5mqSQ8c36PrDg1sTHfnUPaPftMN1xRvxDrs7ss07TBhNh1MnGLefR
9WZ7EL4+EiuemPJLreJUaSlomUIIaHB3wxyGWvzX46HJPQVvaO94idDZCUpHooEh
ymInhemjvOHMU07oIQmLA8+beY/+C6E5CPmqp0kA7lAZWC2WPbaEVFFOZhlcVhM5
5NH80+U78dVtZdhvKg49TpsUF9/OSrB/vYKURIv6ilMF78T/vuh5EhKPUYP4BBaM
1zVg15uYt+mXuNmCYt/0xK/GTTgupqYGS783v0o3oZGni4Msnh4UPFqc3g0UH/dw
rS3F5muCEQXEynFuTx9xcefeLQ/1Is+VtRohvp9MUH3Ugic3u7KjnS8X+Xp0L8Ir
Q55iS8xWQ/mSj4bRldNvkxzJ1/Zke3vtO11blJthzm3tTnJFYNY5RKR3WywSpRho
AITMmnkwCM70CQHcujG00fxHddXTDWHO+g8Cp4dCmh15SFCFSyqsYeUslm5S8ITq
gm8u0zo1Hj7JgIyzDkfaNX45xj1qW6UcT/R9B1Qwbj537vEct3gNho2glSBbs1C6
iq+ipxrKLb+Hc7bILlFM928ORwLXgU2KCVoyfwqOENtOYXKigcu9KWDfOdiVhZB/
gI1lA1DpO2sJK9buDMscHgi4XaPcdjxkunGg1O+JKS3SFUlSQdm1qYC6SfW7FcPq
ZiDdxBlSpoFVyawGdd+5t1la50jAZaYRZNnbxpEjAof2YobwVuU5l0syI+vBz22e
buhSqnXxnpxkWmvY/kLILEGZxHNX+UnvqsWJ9mbYs+/FmJOD9PKkuSEhXE3CKmhw
jiF2FTY9zucaxVFjMdaX+vBKtrAxec1dtIZCRx2cLowDVlEHGGgCzzODglCQ9L9V
p/BK96xzSxxafQF/AvS9oef7UWAGx/dMaldL9Dg8MCuUIDzGhtFEH6IafYSKyyio
bjaiAeg62xdaC6FZ9uDDFKMImfh+Ky6iouT4j7QZa3pEjLWiFhyhp2xnHjjW6T7N
yj9V4zwdyZOJVQ+lasVKnmFlUxelZmxD1XT6xBEoIYAVuVcz/q+JSW49WsK+dqd7
3HRkPevm5G5cvNadXQR0alGzebRQr2ojoQaqgWe9sZFVG6G2vWudbBg8gm0ntvsc
5RsucMGRW7hxe3nxILOKI8VY7gSjCAEMQeN6cFbamfYmsiHNFYLMn+xbmJRcOxBj
EIN0v3kcqgCu5bnPkH9BmIFYrbT/c++1DgNrpkgTQ+HepfKIbezTibGAl9FBVUZl
0nfQT8/Bnz41RlIk1dKYsHNqXYZz+19l+7P1JiG58C4vJhqavWs5SNiszh9KfYaQ
3vQ+mxFJHX8DAd2PuW5hQNxHYrHIiqK94HgzF6kwMer1rnVzW7ixJ5S2fAYU5BAi
hHZVX1qlYD6dak0AHq5159VKpMHS4poTF7uz5rmdlPoLYZpzNh3YOz7schMAvCnf
FyNRaySoGWOQ64aP3sawwSY4BCO6affKcjryX0ctgpzy5/FH/M5QrYgLBGYW10rl
NkjfvXiL2ywN1q5aP2JNhZBd4C0tnfdVs+8+0wFFo6KgDKTVyheXW1SZ2O53NMD/
EiZaWJkpNDOhmsw2FwxHttR8EgkVikGx1q2rfVgdagVNsPFslX/bEbo+/VHesPXJ
zJC36GZla6ZS2azScT+scTV8C2C4xw9Z7zttIb019va2U2dBDziNiClB5xDh0LMR
zo+qHgZh9u3QjcgNLrZCqxGdvEtqzPeHjDUCaZhjjglnZd88TkecfsyXpDtfU78K
CB7+/YF5kZjf5f+i1cskZG8KNvyEoqFOi0aw5E9cZjrvHw+CW7GsYAzVPp3pSMp5
nBEN3LGn0fSRiiBEzYRF0KdNXgds20R23ZTv6MVbma887dnXkVKHWstj6/2APMB/
8UMoQVfbUJvL51vnvPDLeR4w6QH9R6w3vm16FKclsEI00hp47oiUXl6mBL9M7jPR
5mZquh4rxBEfhIiczKbH6DXU4KxTQikayq8+szTDBjL8ra9sDOCMMR+no1td+RQw
7UUEC6Gg5sjnghsr2dwykKFskpbsJT/jIFeRwjnH8j4SrmFUuR+927zUOR3eCzIt
kTYtbFb20+vKzceFVnvRWMoMjJ2hh6Ga+OONStqV5qUGmoIzUUlGXavVqAsy6xD6
ta/drOPCaWFlKoMDoyfXr88yEQqMxbpkBVjvWnuY/oCgDh+tMGbP9bnLsKq1l2JZ
R42/Lf/DQjD1fqI1BfMtoKope2wmS3PCDGMXIxbH1nrq8LRNuM8jnTCfM8f5IVeJ
00lfJtAiS5IivlP4Pllh1qYj0cTmzDb5ltfzf7SomCX517D7N0RMOqUPPXIHc8GY
9xrmZypLeet5PkEm5X7fhEDEVePXDW/AUOrFT6zFj/Y+6WULb3o/q+aNcJVbZ4/4
fOKmcSO/Y4yuzMiQvkarskvmHZ4pr8C6P4ORAoXviSGAgYSPHzH0b6HL1OEufs8w
zJZSr54bXuG9jEX3wBpYZvPsGGeHDuZjhlPFaVDYaA0qgMmzf78Bm97udh6qrkf1
9SX1MDnQeosuslb2pt0/FVAT4ivy9w8EJqqfh9TyBS3OYxi7C4ZNUiUNTLtd57Rs
qZSO8nFgojQBwEL+BdtJB1Gg/drp5rhdDQnXJl/IySqeSVc0T92Llj80g2YDcc06
FpHOqBagAeYObrbVdG0ioF3Np8yofgBU82fsPDQ+yG0Rd3lFtuUh/Zlx8uDxmMyR
yNkPXd2pTLGaBJqgpF/XA3/Y5UoDRKjLQxcUiPR9z2KYdfo1/fB3rvqkuOntnMt0
KeDz+lREqqTb2O+rYp/WpMgjZSvKo3MsqmCtM7mcq7X3YFMhYpA/maFGV4l4Q7CW
9Z/rP6wiW7X0xwo/Ut/MsEXYmxWJnPvzYtw7BMH9iJmC3ZjS3NkQFZ6kqcDzFqM9
SCh/nb7iJrS4lBFWdYsoGLYPPekq0/TWE+RwkZYBJQBNS2RcTRmNqkjFiC1iJtaX
5fvtLty9EOEsUNADxOLLxV30sXdo3X8LIEIVsSSYNhmPvtm4tGUOYzwQCzjdzDgQ
d39hssM08jxRVRCBlrbVjzlrkQRXaSjUqb3sLj/Q8Kux4krYc0dt/pEKFS6W+cX1
fznJPaenVHUwSZTJfv3yOmFFCArKm62B1dh/7DfFsw0PlvmzXXQNQNW9/GSFlgEN
Stdu81s/4dx3qT27O0UljD9vddbuYVHXj18j+7NRhMIxpdu/y8NmYadP5x30cU0b
xXclNKiqe+CI53EYqIXptbYWkbWRDWIvSgIrhJTSS3u+/XiqGu0zt8CGestP4oed
9pzu9PD6ULrAii22fZdmdIhyS5BDeDMdrNLHalhXcPmiaxf+66He9NBxQu9XaFrc
a/Xz9JdfpdHVP+/8B+FBuXdWXXnqNuPVZpl4lvySmbrXUhrwrMqLIh3P8miBSWBO
xHpocMCVYUEhmEBC7Gfe+X9GvIPmSQv+rPECZMX5rhUL/BvTOSBSPO3X03ZmBz3I
FjRXvQC3uKHVcL5uhfV/uY0hT+q2B0b6f5nSbMvEb8JkfvA+nbyzxZz3+X3gDcBC
5n2VI9PpUElU5mB4jpqaoxBC5E/Z7BpMExqPqa9GbHA8kfukAxKqjXM/zln5dg3S
MvsVBMt5GPr4gYy+wN4raXs7CYMqfkDuzSy9cxbo/tWCBheYv5J+aMqflpf2mEAT
lP43TF7AjI5xgUd94DxCsL1SygjZ0xMxymoD/wOiZE7L6uLjr3AW/V1zAqMQ0Akf
DLJY+a7gmvzl57FQh7Y6PisgNRs3qg/dcGnoR7eEHMNkoQzHZe82g3O9VOrhWZ7i
DMgTg8FNaKJiAbfZlalpa9PLWsVWDOqaAhnXg+PYL4GS/J73wGqO9caGPqcFzDIF
f0eLXycFT8fHub3ulLj9tB/l9eRmG4GCVoplWDfzZpTrY4gf9kcLW5PoKiWgCzdv
2tS6Gdyx4dKzw32oSb8Wd289rax0eIr1X91fmnmS06BfqIUWN8V9fWNMJfiD9xsQ
mSLpKfe2feuv1wUMwehP8hbCETT9NyXrd0XFpY4/Bg7yGMP9fcq8NRX3VxniZCPq
U1yXxqkRAqOQmdb2LY9XYQAB5MaX0thE+XcsjCWPmjGy7tePT88FnpW3HTds/ysx
7ouLyJgJpZUazQtCxMYYeLNvTjLxSLsNEGVNmjYJ1FHByLm9vEoXkkME36p9nQl8
dZwjANv2OXJQmwC53YpIiwvP8grr4oM8cE621A0ir3Vg5Q28HunolhwNlxayLJq9
KNlL6vGuGSmxTBg8V3tJMq/LeDzJkjnQu4mPFFE6VA+rjHMGH70ksqrwjiktO5DA
gAxDl5JXgejuUUBwI4sahLVCgOs1WXHAQU/UXqRCWQLhPXvYlwgI9rF//PQlhFof
iaM+9P2YEYCwi2AMlYWPNrrLTynsPSkFZjDuA/voQgGhb/82IFZ3d5eOO7Dpi1g4
UxOyJZ3Ahd5H3l6kkDxxZrhjtdqM2E+/oe5CZeNNpVD/FqbkLlR6lqiU6sV4BjNg
k54Luubfp3tNEy4pzau6PMTRMj8gsaKcg6nCXLJ4yG4zrGRQc2l4tSmkwoVopOvh
QtGvJG9VCgGdSa0Tldo/vFN0GgnguexNoTqUaO2wcWSM3ZKN9h+ZRmDO9vCToXcC
tDaw5sXxBwPdZNcfx5zbmjmZUgCeWMgtuGlvBpspDVZsPw+zXSeeBpdJv2qlOZfb
2nFNKVDsKcozoJw2DXEkPZed18iYavZKCXNONMxdtuZ2gp19ctLl1lYPzWgrhR2j
G4pox5G70T8EFRi0onfWO5fKt3s4r9CsMadXviOAe7aVZ2crtGPvc3W50XGijn3R
BGT+XhpcRJfDDwXI/mE0i2JXLjFL5gtr7HvfvOWOxGg+Wc5nwsmi0f6c8BXFD0Wl
8ICSXVriprTcWkpwAIvJ0okeaB0dlqdNIyzhMiwAkRXntSMOPMLVtuecRpS8ISZk
hGLdlW9F4DRhJ7dwzP+1YHj7bkkWVN86o21zW45POq6yJPdoXepdIuk97c6PH6Qz
x9TEwLA5MjXFGRNoIGRFvcuu6IIHGuExd84yf7bcHZrwsFmbufo5Br6WjWY8FfYx
2rmpn6CQGLclHJ+RcUgNIwtTADxtd/lX3YMfVlfebETa3giAtbnz38A1mA+Exob5
ZK4C4aW+kdVmfHIyi3VhBFPsudHHkOb3ufmO8yCDfkh+i+q3oNKQzxaLnraUDH53
uEfVOmvO6RZVrUDVeex2nKB+oJD0YzbpM8spzzOYs20rqvgm9mWAaGwWOtg1XT25
BQgKTVPmuUjQW02GoOpVFKxNSfyqKhvFFVF3RlvrkGDBxAdXjl6Qf/laQ9OHvPLx
q7YgRTAtCx8XAJHjBDnUjI2BfEW/B2QV/uIqMJ1/dIl0v4buMWN/Hc3yELhWL+ML
vmPObRZAs53p24r7LayomeP4YSj6kE+A47TJN9j9hVUjlZaybXaXNMqMk/xjobv+
87SWFZsbobmNQgblpKbomQ1pXs7XJPZ+1h/M7fdkE0xM0E2qgef1cHFup3aw4ZhT
TMmvsfM9WuIUJ+4eJfTImMCl9BWLKrfYWHe+7O9koS8yT2C6pOcrF+ROOcuh5zHO
O5m/qRETXmdZvmUTeS2CWO9+PfALM55Jt1fSoEq2FJAJ75Libr1Ye+/R3vPP+a7f
LmpLxqaeKsYpB2PyE5kewtmohl/mRh4a0rdZ4MF27LyLn2m5XkfOPF6/WD7i55tp
A+2+ywh3Ebnsv+8McUdCrvAwLvuSgaw7h4zAIrDXjWjLF1dmCW4czh3o+pXDkZnv
xtj46t2zLbob9sWar2nJeL+2m+E6CnmnFkYChDdZNc7jR8dJB69D9SLc5k+Esk2i
UAAojSAjVRkNW7wjT08urm1QJX2A1BZ9CM4b5841XBscoUx1KMvVqlBrjzOVehT/
oqK620A1IJ30ts73KJyIwi1Op4oYkRvgYVAn3gNzHljjTC0SSnAc+aH2eH/LotY+
I8/BJBivN1yvkooCut440Cymiz4zedZfqVZHuob5lTEV4z1nIO/gjg8UjOLCIaCy
PjAFw/RKT49jV8AW5yyL0HHdQ5jF2ThR4SsIYl6MH3DwqXEJqlRwY7qXQWDjvIsD
XWoKPyq7Jzvqag/RrYI1qE5x1L2fR5Z0LzEpDkeyNOI8957VMDjY4JRHpVQMNtPf
OBAaCdaKYw7FxacMDanU/UNz1z18SCMNiPfUrY46QFafE2uoJKAZtEPYTX531YzU
9IjsMEe0xfe60SGl+dub0G6H9q6KU5iQ1HtXeRO96RfELdJm3iCpPX78d//Uvzs6
pbMzh2gz2RERcAshh2FvodvpU0r3XukqvdE35+Ygm3Dw5WGxdmDTV05Dc/lsFj79
53EPe1vAEn3BJK1HxWzwxe1b6mi1cW/20I6hTf/74svz+XIOH8guLgdIRcS0kE2E
bH8OzjLVTky5GNyo34LwvDjwETMrATE8KCWBNMldduko7J0LYkz+heiwUeL9YZye
8tQpqbHRppeJSnN6VFRQ42n5G4M8c3i7FzDIL4CA/CVw0z5SUKYoGlewUCpEoL9P
vqIxs0HVP3/K8e3OtRAk6gsLCmTfsn5Dqc8t8fgDOK4UFPf3p7jcr2/j7rAtBKB/
Dva/tiUjXVOmuy7+I4xyjpCiGDT8GD5kDnaEiiTuOa1ycCMENSdD6VViwnOTbeut
+hGr7SSNgSUs+LrhWfrXKqsRT4/RxhkRywSyjCRNs+BL44n2Fn1eHquLsFSRJUmS
Nl/gSfiI7xGPsDl9E1Q8dLVnF0mXQ5H7F01Cn0EmjpSLQqfQfg7aqiFXAmW5pcnd
O10SQ6Mfbz7P3co+doHJILdaqB0w0o9R0yGDzNSwHOYD57yg7CWPFgWi84Z5pWf+
ecjfkOu26aHEttYnbfMgt4SQwlY8PAiHKNGnyYe2tyqkifB2tipVXSUig99BP62N
zwOfH57PlDmVEQ0AxgBKlTGPSRjyuWiupJg3n85Nr5xSYK1TcNhNIngfHmNJQWix
002mxbNt4roHLnUZPTDjd1K+OhkMv8O+HhIer8D5+9rFEzLg8n5NFYacwLPsxkl3
wYH/OwhXgBpbABTOq54G+gKAd7vhJJKUkAgSJ3QiYPUnfqSosGLauQuvof5jGbrJ
ubEoO8m8m+8thtig4XYcVL0erqV1M8J2L2iroqcXtg+mpuInbOp1AsnkPhrwMGxM
A3pDOJaC+N/CkWrN3w6ePM+3j8IBg6WLg5LcRv6DH1OH4CUKI3IxoBvZQoJ1XiBy
+J/f53htWLsfKftCx4aoqtpqL4dO/SOCbctOnAhMB2oOlsqf/Nom9U8cCNF/zLfj
h6HM1Q9mgpGU/7MBr519F0AW5DbLK0OEnSohrSbk4Oh8XAmhyQupg6pZpdNFnroz
KCsQqwUJV1zDgWKR5X/onbosiaSatIUvlPvxNZ1swI8wfyB3FEbLYAzzLkZKht9I
tbszFLsTQ7ZJHa8qvPmTpTt6aqKKTi+UYdvtBL/KK1V9yPTjpqZhvW5nQIEHC3M4
Z3Da7Fry3Cztpq5O94lgSRd2UCsKmQ3U694gXEjYLZcYmVEU25JVBg2mCovrPufr
oTOq5SAz6Y2WKSczq1moE1QVSOSk612r+uPLim15LAkjUGDwvfgfb6X+aqjr7Nsh
nXQaugSqNHrNJXEbjsypyjgR+LHspUWn/VKvHcugOl9s+zlAcWH3h2yvCcxNmWNF
5M6M5ziR0A9NdeRB5Mha9tEN0EYvKbYTzePNs1lvLeloXityyz1BdF3UShNgyw4d
fHvwGRLgx0CM/JtID8N6GmnRn38MV8i0wPweGeKpy8c9TSxKF7MZ2afPk2cF1Cj6
+rptVoSTPaXv2hDA+0/zJQCM/xI9Y2cleJpSMlS+x3eeo8GAVAiDxxIkSG+pRyKg
rfwWB1S9xhb+90tqXR1AfHhwyRkM9moOCuLU1gPb4h/5yMFjMrIR3v5/wTzHc26a
bNxq1vAuBdjgDu0NI/VwD75dTCW2Qkr/k5bGaNIJ5HKcf4zG7OXPYkX6R0R4yynT
Qedyb9AqdEc38BD6ELuXBSjdXM4ruMndJrxffPT5G5h3gf1MEsGQSA9mv1p2hcl1
T2qtYUkRotf74LARwkKAWVB8qusuKVgChPsrHGRussna2DgI2yoE66hvSH1VVuSV
Dswfp1i9uc9D2eFZvelzwC1tA7KLtA2rNH1S6VcWLpBHLcbiOvUpkoOGge0JEmot
+TzK8k7Aibf8O8oREhRGbHfqtB/5mcisOfKV8I0scc9/CqVPIisKk6ayLy3umwAB
ZYiIH18gp5uYrruzfg8H5NT51MhiU6LpHl+e0IEsOOc4x8h3MAFk2pOXZOvZdkHo
AvNSWpRyrkziO7i5s/tM1f8lkaAQOKcOrAxSltSuwU/m8ZCNuy7gfx3Y9Kv1V30l
k9M+TU5XulIqjJhyzIbtQZPd3YuA1OA4LL040zekD8p48JjTrbJIO86tuX6t7AMk
eFOWg5CGArcH80amh55BJG19JxlicSlULzNJsHuYVDWu9JCGlOz5K+vHW3eVyBxU
AsRwiTI/Ts56aaWIii/gGQn7HG9JJGBGo6x0LWOZ8QUrZQbWUnodfSjergvK9MDP
g3bC+NlKmPlTmJCdVUKdgkhZZyvEQJIA2XX9DuehnRBW2yAmCWxuEnxPX4VMLNbN
L4+Mq+vahTQ/ay5yxHR+5bK8Tw2pRXJ2wC0UWAIxJS+BBjL4mjsGkqY83st4gIAs
eFuPSEtwBbB8XxQHl7FAEHEVgZNiLbtcoNZrcj7DEEoGNFBtV7hbpECmnLVNAGuD
EmiglD3GTQkuMIuvOY6gO/r+Nauy6k8X9omNwIf0DGknXQ1nleyfTAQkoWFfYZiP
1teQmk6E08Z2pGj5eWo/vSe87hOMvDFZZcU65xX/sZu7eIq+LLmSh3xE4qMJ58oM
vq8tAQvw2wemsqUJNBrnivjnJlCRBR8fS0RkM/wyksb31S/GG+AAwWLXYddF3ntO
DlWkh4QMA4ocemce1VV/sMUYZM4r1mmGF/22j2VvhAZzKtCDQfsTHRp5GvkMURqJ
ADQox+c414cTA/EJOlzGmf4tKR/Q9tFi6WTPqT7x+wGfsUux5kob5OS7O4OTrN4R
BbJKbFkkSj38SYu7zsqR7iBM9/P0EbDA+ZyeX3ZypH3GjAJpV/wllVWWJXJNJydZ
E8epopUyG83hnwDle3tfFuqKjDwd0FhykmFWjLkSg62Zg9EPRv08Gu3lak4JIWPI
NNW1Z2I44QFGowQrRB5QOZF3XQTwUWFqtkPhAYy9STc3JSb0ecgXUlMK0D6CO+p5
w6Cbda67Fnc5cjSWCR1DtjbKpMwcIyGH+rh7PlfvO5pekDIlmGv0wa3BmfLWk64f
5/ZSrXUb7Ply7oGDUXY7XlWv2uMVgSxrfp9MQ3PpbvUdUpTsRToK/6jM5VtDBtYH
YemlEjK0r55rmhdHhif++sn3GxvxZjwHEJlfCM59e0ogRsfR3u2Pz3FfhI2eHg9+
oxZlZTsWFVWmhVaFYzmHJ/smXjjNp4jG37nejXgk8IdpzplWlZYy3u25DRxYMgsw
lY9dy1zOH/douqh4ESmf0UbxhQ5itCvdK2uss1y7ti0OzLmXwnLn8P+HKlijv97H
tx+HMOoDyax9ILP9qS3gzbFU5klXhZ5NvGtVc0nI9kOVSL4D0wBIf17l5cBi5Yoc
QzDTmVxoB6D/J/PZusztHo03G1rIGEyz1gvAOSu0zyo8xhz2OpeYEAA1FTYsesV7
Onv87qeiEhzlXXipzidzEuLjekXiXSyfVU1OmhdBF9SjFJOxZuUesDh3QxEa46rV
P04RmJB03E5UGpZA01MV+IRSsVwYOcFrUV2dUpMDxEDrrf6+tFOsskTu1r2vKpkd
0Q3TNCJiUYrXrdRDIPFGepOsddLi0MNX7Fg0aJ5y0RKBdn0o7XabnNKyiwXtr/eH
r0pPI2qzOjxyTs4+IpmUdRFPlZ5TSezXajPtUvWGsX9KV6f6B0Du5YtR0wEfZhtu
mhqn/f8W+nqYDMzkRkSS/Ge2VL5wpG69FFFNBmTQgAMtHRePJCQp4/BNvJPfA27q
w7TFJHl/imMlEKlKML51GMXHX0CrqbYq8S+zgwajSotaYCvklVr/3cNdpvpwzgHw
HAh05noaWIh3sYEI1FELp5EPOnFBiLOJ1YkQvGurCzo0LWtESQ0fZ0/nO3Yxx9Na
xcGs44I8r2PyVWYM3XQ6jxJ6DcHzB/kEwakSxjjIqK2kTJW5oZ6ppmc8CqxOYM/1
qrkOONIhrlH+LgH6B247hrR7xx6BXq9rDJBOvewncw+3KHhWfBATTnDOawsV+cfJ
EJqMvwf5A/FDAud7DPY7Np2Wh2j95MVC5W29bxOXtEwmcjqB+KE0kb9rBxcm6Zes
ZGAg+Yoz6KHtGa3aS5wgVRbBhNdsxvFyeE8N3gzgHmcKSd3J3qZpp1nQB4ZIowIV
qqEJRv4rA7yynXTeEXfxUJrH1qzNIZNcIVxyhvIFNuk44W65m9Qq6huJGV3kt5Cz
ULwBZW1xfWwbPs1Fi73yLSRTTeC5rTfvkotiUNlYIWUtObLalAK9rEail0R3uDEO
XGMzKJif59NuIvoQmM8XfAxYWZehijK9kpY4eTpjEnt4b8vpcLMhidTWqxFw4IIP
cBPHyjGbWldeZpj4SwC1OaykTZPekhQyumGfKjdsVQIxSrcE2r1K86CGCarW2msv
bJvWLPkysAr/GF6poEZnehYFNKlpSacVTUDOAZCz5sJcnANwcJD8Jrh3NC9FSsOu
jjzLMoOl/4uMIhdKOA6d0teN4V6CPpek7zx0UBRHTwGAzLFU6gcIfJm2SPRu4g6f
cn6fLhWNdht6xtnrZQdGm//FihatcxVbYoGoyLYYBra1VJvrP4EMipuPRJuRY/qB
Ap6KK9E72KGKT/L3fS6x4nBhZ4Z9FDIiUrErUNgnb5EDWm3AcOd3hOmn184m1vnh
CLyueW5JcWE4aTmygo++gAhlnVQ6kP6nscJB7/O0Zeo6WL8+zFleTo7m0EnO0w6H
RTcP54JxYS634Lc/nbfi0TCN58JM4xGtKtclY+d/2IMQvh/46PxVn6cpF6X4/l76
5htRKU6zFscwzai7RuqEoFR0ZgRCNy1rY7goIqNaAL2+v3ibX/2muhXCedSNrWyG
fiJPsGO+xl8HtBN4kSXEa0PCJ3C8mCDY/RMWhU95buLKneZAhdqUX19v+Xe7ii3T
4TZuX6SoYikpr7+QK8q8WxoUIAiUnE45CHgzMiRULmOvGdFjrgJPet80fMrPUMxN
LxWWkA8aatKYlNK1HtUwW46HmpcWAXF5y5WrHY2vkihMymZ7JaouODccU4+OygBv
KHwQoEIFSmGAPB0TqT0nF5FsFeuWQ7NZ8FnklFSP0uGcsVn62utbdWu6b0QZmNXp
5373ld2YHYbzPPLdpKRf1vByRaF2+IQDeH130C2rERf92ddgFhk4lmiDJm7IBj/y
pz5EOrylbgyH8Jw4E+ojqCX/eJQKJNZC83KQLRCjk6gvvsjo0jU5FZNxJnX9WZwS
Yr8hO9MZkZdqo/nDUx8hcl38bB48/mM4rP++LXs6v8Ii6spBj1vZruOZHja7G0Yc
JEBMjXU+R6gzAX0eyXYCOIDI3qYuiWnhAZBYIJNfWz+8mCNc7ZpKPhDvxij7i7nD
oy1F3iZ5tKzm99uqfa+eK/hvay4ZygA6ITASt/WFE/PYLJlcZb6paFwwQ/sWSXwQ
2+7y8ce7dLNEzYnUQxcrqkSjQalmaORrmRWJREDtoC9/7Cxn8Hi081LyYV6kYJWu
wYpCujr7ktXRPf9DuoMZEGLuyD8YHqmk57d/zWT5Y5xKfuRq8pOz8blHqvX6M//Q
OOHbIs+mbsDNjiWCtGjfcXYbzUfuZfwSaSelTitVXB13BYAHN6KyldzsiON6R19T
zk6TD/rdcB17uMIjDQN8XbT9k69umR2cgqPtvP0tDHHqGC5qfF7fCirkrq4Jz6i0
kqV8FNpGBqtpmm1Zecif3tbYYAcLs7/VFDVfyn3flCujUnpSCYqyYAJD/BESZz3D
6PXuiK2aWDdQlqMzdogLuq0V5wTYYrT7z0hFZwXOL/VlFO1dKleVdhrA1g/+sqiI
vWPicrOiVc6dJIkz13Jb9oU+zjdYorI90nKtnGicNZlk5ojboVXGDdwHTEJft2ar
ddTkLkRZ0qKiDfVnJg0ztXjp1JcuEPfyRHeXHIfiAVWWi8824CSY/FvnuBRW8+N5
DwwhFXmN4qFLZfz2mxaMds6LFMtdC4A8YFgoSkute4SEBYt1b9UVeNTwdk/JHYgw
rcQ6Xn4e9WmQ6cfnvKXciwdowIpRKHu6OVbwtmfueGfZrEXSNAW6gfFvuCiK9XFD
w3V81MMaEs5LC1fn9OANEF1Rdxyj8Z/obP3zURF5U3hHFPGAEINvdgkpa3jyHwN4
OWpfMsgBDz9b1ifq2vobVfU9ZTlz6vkd3B1a4Ku6q1uD27aosuQJ9HN81gcDtH/j
8dd2lJgtpKsg6VxYsB/5ruK1jNoNFioJ6kSiH3B7H9lGD6r/hJ3uWTrLQ5y2m6ze
xJ0YGueG1zV55vQL3EhzcpDh19XtFv8Qjfto9DOZLmIDAa/BC23hbaY9eXnMaImF
bCe7ETMGYUZ3XUIZh9c+ZslAjn0mS4Pg9NBdMsym/1WriWN814XWoBnHfhhXUU4r
edL6CBo2S6nXtTtmTPYC5S/yN66wlGUsl7TgcTqPW872Vk28Tdm9Tbr6bkEIDO9B
BPUNkBpJ0gfgo5bEu9sT8RAwp+hqsQCr3qf+stV6f2t0oqPaXVk6T8IYf6rt7lD6
I17hxkZmx5lUttMpVNZ2iwryrLvu+gStYxeTzXlAdnrJBgJpa2/h4eHJ2c+5L0sj
lTKM6/wSYeJ5rtN2JTAW/tk8XAxiFUO3a0gS0UHlzKU3gvcbKiUYakdGrKttk6XD
0q4XoYZpwCC+oR/tirkfx6JSYL1hczDhqF/esb2txwTUNHhZev/EStHfX6QqdRhc
KPymxoMaUM4KvIWYwQb4AE9AtzCbKeScODj9sKkyI3OOWIw/sHiTGzBPuYvnckb9
jrY/sObJWQ0DzRCKm0/mFum5ckSHvE4oSb9D5rHTgqsFl3IpjuU/bQ4l7WgIB9d6
BGzhQd693GXFYx2VUj1gergdkvWl7oD1YttXNt0zk+XY1kIjc4QFrjrUleuaDAMP
MkNelloHGZBKMXodIs0Rmy82LDGfZseCoMOiDsMQEbABpgwaqJvlYsb/SsuAaERt
ghhfBfXH0oTNPgp4ucc5XN1qP1XqsdOO8WuksI1wzwcRfE9gforZ+nr5csLL9UhF
C7/Wbxcxb2KzKF3gwpaYOSSQEFv3EjGlwSzNj8pnKVj3Mx0oi40l6NJSS6ht8wJf
teuw4XS2DYEyUAP44bARHtmTFULw+J7bWADr6gFeDsrbhA3nPlltDSXD674ibSzz
ul7rVJ4IXu3WolBfUUnuqgCaHi6M9uzliHDglPyYDhZ7JpgOddDBSml0PGZa1Z2s
xP/hpJV9v5uDzv4F4WfkJbnirLvBDJRf4o+rumyx2yyIltCdAyvikAHV9cLqrdYG
dGcmGByH2O36Rk7X7gJ4XZmpSp374XsRACjzFuXj9D6pefKzHHtWv8o7avByl+1E
U/Z8oe1YoYS6iAnMp9SXRjErBx6nhdRWZKTv8a3/r2mB2R0zpPcUYLxyvJJ18Wdt
f8PwPnFuSxP8gt/ruYd7Jfp7hkRg2yauGB2ylElcG2bBltXtp3fgCGK6l5ckyltW
omr7O6EOydAqtT6eL7VxEMm5ND4Ykrp9PtUVRhbVTWE6zeCmHxWUBNjKSQoB/5eR
5oNrMEqRkzhGM3dLGHzTlyZ9DEkk0EpINZV9hU6Rmp0EVqSj9X80rZl2KkJ9ei5U
SgcgNxT5luT9ZgShI+RjmUTVWT8wI9D9HEi34xtiHdLtgf1SwjoNR1OgjMzfH9Vb
6BFUE7ZCzM7Wm8L2INkhJ8hV02B4huY/d+qnPStOCjylrbnyLJAX7F9H5emHiboE
ax62eHaf6Z5v/v3at7pubUgR/Uhwdu2vxvTXjvvYarG750mumCvxnLWLOlZIJ3W5
+NNrN/ttvj6FVPXh1d+U4d5QOCOczBr6h1hs3Q1lYscUdUqLHmxeKDS4r6VLZzhe
beJ0f9/Mf0QQdDMYg25ZKMPaQler6I7Ecy2KBEt3w5lXmg3Xza8WbNUwT91N8VL6
ARRGntDuBcdygnZI8xcpYSrff//xVWbYHSqJSxWFHCKCXg7GziQvbR8a/Zyw0bqg
lZGA+nLVOuPh5ED6IN8+UXFTmty6q7q25cbrTTOJOFssFxwEHu9d93emifGdLe9J
0Lc/GAr5phzuRilzIGi0tsjzdtyC4xiqTcevuA9RJAk/TPlmn1/TGfiJ8Qspi71F
gM6tSIUOtkZUzp5E17cF5CPtripiRzDANJkin+W358Qo+cOiWHmllfdOF1sqNGDe
rqkau0YH32DgRNQR3vRYiNTlmNP+xXB0Uxt5r0dWxe6mBkDMiRaPY1TBWoNStOIv
IhZSFcbwU4G+uofQzsg2wojk9D5lhgciXCvRbPsC09D8KwyQ/gQ1Xyz6zKEEfbZZ
u0gdZUobZf25yX2JIWLTeMnf47uHqLsYTWxTHmIXFhE1e2bdurfqNIE2HGxA3RVS
oeMr9NlRBrz7bg3l3BPW+C45U6eUtNdv5QLlLRGVo4Hmll0j2eQbmAQtogoaNPPR
VUCRjJTkIZYCJmLRFRjKFyVs9jP4KW2t+FVfF1GMn89lYgZg+JhdHmzWX+QI+Zmd
nfuCYU0UzEirZnwMlPhwJ/ku5Z+BA6ILCd02HWbiEpNI9kQGP9tMeRY51DZo3cFl
UGi4f6R6d6N/fBn7DsYkwu/JhztEosGXpGOcUR7KGQrZ3ygUc8FYLH6JK6Eh0NZh
eg9/GmfPpKihMRFNHozaGWBva50aLMf+HSvEl1JZesOmrfzc/Y18kEWwnfScJAJj
WY5OGNLt8ri5LBvEwXjv3cDMBJPAmTFllVyTh5asNziuRQSOU5lkCjhkhr/ghqjR
DKrTRQ/tCGUaC+EcD48p7TlI/otJEB3FXSLjD9CeOxSPLnCFgRwdKmx68mXzq8Nk
jRdJvoD19z/hUM9++Sj7nwNxmnh6KByEqwfL0zDFztIVDpmW5FIC8k2xrhOcN0Jy
WR22XdSFY23fAsnQlvQwM4teFBM2qZugRb1Wteeckf3gLvN1mrpsgaGb9SsYMiVt
98jlESgANnmAZtJ4x/23lgts5JLKkdhR/4/KrgVrOfsIKRLkZoLoLuZnWUPNCjDO
pmXoiM7GtbTQ6jtVq2V6MvyEnxREKP5v/1RD+OKqqkT3594H/IM5ArHJldKNOGvD
vKUrfKkPmP6Wv65aFXy0r5yQ/Nqf5F0jix3J6+/Ek6+OHIbb0qTd1EmhmDVLfcp1
K2ofQuxTmol+1DM9oogXRyJOZiG8rSpuwZEvGCJPhbSihDFj1LwudlLtUEoDDg5B
ifvlll1wHtbz8XksOQ/qm3h8y85S7muObuTlO8ORyopAEeZpPiZ/XFNa4O47pAFJ
WGEZYpoQ1RsR0ao/95W/UMUOC8OBL05FdEqJ4hCocN0zA9LxWGlrVf5JUKbTXJHt
MGZx9scZ5fQpMqI8usuBKleAfbbd5+vBerQqsw2FkZpenBXoDiLhBULLf0Vv/pAU
1FShYOJ8HmWYvbrGGUBjOR74HpPLi3n1TKD22m0fikiU0+2dxGPecBG6YsYi7TqS
HTTRncfVATPsspURXO33GrSo+9H7OcRwoUI+FXSLlzLjIe7EYV/71yymL5uXKCs9
uMgmB6Iq2vrY0xh/+E+lZnASjnJ9P5Uq87be9cwY6YQzaks5K0ZTOGGmZp+o2LxZ
zC135raO/Uu4Fl5cknZ+RRTDHJukb/h7ybX1hm46kVSTTkvUkOXXCHjnpWQoo+MY
+wcf+pkaHVfOpjUuPTrjt8GNZfkiUiN8R7aPxg9pUMGZtcdOxCX1GpffBbNhkqMr
Y76CXYXvZOTTwXzHXWqVXLW7w9k5AUgYYe/FuKw8qTcOYcljMKGLzQPp8s2Vfz5q
OJXKXDic3u2tffxl24j/mDhlE1BK27e1n/C4iwRfG1aW7MeXG+7WMoGrAz3rZSz7
GFkzZc7X5MVhgurA2sBzujdwVxS9f+6rN+wzqUUMC7mxhbm/KTU3i91E1jRMBjHt
xgDksuPB6k7iD32Pcxa9iayJlV6yrx01iykVtHu4kjC1XxuiPxJC8v2x1lhcNccX
BjMCTNKMUH59IBw8XeKqGcB+iI9de2EVQORasUDY/1zzZ7TbruxAYKkIM0fGAoIQ
CZULcnn3zVWAX1jnx4wUX9evMla9UjDlX8XGnaHc8ZV6Gkn2AdDmjzQK7Juo+Yox
Q/hoIMPoUFe3RLMOJeSk51n4gYVCM883n0t/bbl2YHN6FLiJYbYpjSXmCsVcmc+s
NxXiVOtVOdVkmX7kRYlKi2hT9Vhdnay1Rhs2D6AjXGNKvXxgmZVMIVAE+KsUDRvv
qznS4bTYg9B+jy4QWKXx1NtPxoYwpm/oAVHtG7Ti+0o+z9ADPlmPeWaFVs3eHXpL
hGZef1NzSsEmljGnnLQMGHO7UThJQ/HHvs4z9lOr/79v8zVVg51hPIL1sXNyKyV0
antVfiJrr4NeHZUPVys2XDj6cx1AIBG9puFhXC8Xcs93+afDup9K87PBHXrzzpqO
vxjKkOFV2NrUBPoFIY2/t2NT2l4OUG4/br4QqyTegtO7dNbBzZbMoSCVdpqXw7Lg
yCtPNfkATWHAO5NvHG+V7KLcHpow14EfSBPPlWTHAlfGQnFZg31Yp+z/sPdFekUB
D98qCfpuIRS7cf3KfcoRqhKFh/UrH5B2tvgLnmXNOEWGmQHFVvyNKrIf8ruo1v9v
ZVYA8t3BBQqc9XKUxGRQHoAWVts/BB2afjdUfAe+Xo0MLBxEvgRvomdKfXjSx09j
pTP4Hi9i/SyR+UwaHenXmHCJAh06G+nqvajHMGSHz7E03AURuLfyaAwhdDYw3CCS
IYIUel7+9VeS6tMtn60wWVbEcyRvCNWla1rcBea3rYKKhZteAADOIfiRyEoACo4V
1FSg3WkMg4w8mYGhFbz1hpu4G0G/r6X26LozZ3VS56iaegMDglEt60HBoQEw4qhU
qaQhksv0pnccPjav1gjCDCZCQ1IzJyr48lfpYDTcdrnQhgub8JdtQ8Vun+V4Qnuo
VBkLm+MubQJRn2VRk+AuTFyL/nfavl3bg2pl2KttTziJc8YWEGE2q0U9M/dulYOe
JSYuuguywms+eaRgFzYLULp9Q5xzZfp0DUPtZL4hOf4g7uvTOe5aNLipt3eUen9W
3lL4IK0Md64zlwqAkoP35+SAOng908Txd8nQWg4iZVed/W7zwc0tJdD6xFWaLaHP
yQsk2IQ6yJwqzeH5YZj9wTkZmS8oW7WZHd4F6/zRl7Z/d2DGEQD6YbrjztEFmcmR
AVD9gmNXptbInoB80T0lsGrNBWA2oRi82VjDLOnmF+EfIBHX9erzUlmfzMBhwAw5
Eqx+2rnPMzyhnlkLj917msmosMwIrhFnv6YypAoLylV66ZyDrv9JkVd2NA8Wt/im
egAYUOeQW5Suw11zlxWOeO1Q0/1D17tYK3e7I2O45rfIhbw8aBDOGSPcNrPiQVVb
ujK9lG52Gd4Fud58y9tkWuH/TO/ezRyo2614KeVktDw3tr2oX8Xulo48A0fiXdfd
0bU1QS3Kcu25KquGBx+SfYjDLEF6u2A6lgVssDt11cXpagXo74xh1ScB9ITWknnc
hIfzU9b7xTYe1k19P2If55ZY5Fl2qlWlbZAm6co5ORbKsJQs11JPHbO+og4iPOEM
K3ziWZCphiTSo2dmG9m/K1QOq3a+GbGFcm3jHzNoGps2DiM7q/CvZV3mitZrvInS
PhsNMrd2lPOJk6zkXhjqLTOhMWnueYsgsk1hUNAtg0WUAnah2jO9EGbewpRxqKTo
SBVtOGAWTGMuHJwIyZ1V9ugDTFDojTah0QpYFF4n+8M6yODdImZYp0cbBcigeE3q
yki8790xIM56PIiJRF1CfDgAw3d9R/yqd1tI6IcSS8X5qpz2juSq3T/AoBivx35G
OridCec7i4LiarsLDGtlgc1V3m1x/+jmHh49VMuKZVfdcxTkymzr9anooSVDskR1
zOHSKC0fFW2xQ42te7D87KuyXxdR5MP7NhrvPWvVO85/vLPXt/ZZZtZM+JaBLS2F
tBnL3XwPa2mcyfkqZm7XBHP1lWbKIWHH3Y57Bp7jvYx5whT4zSegeA1vLNJXHucu
pQW9MG5hNC3et4R80zDRUO04STEZV6U99cG1jN0dacClOHBwwok6ERERvd2eZEns
OospuiF92vdqEYMhzEiBhFfV654ojku5+ECYYPmR/ewbTWzhbUdLVrQAqK534cE1
MMtB4v3Obrr+qbd6izwITyFUnW6oWd+2ZL/djtU6pDd3uPkMpmigWiRdzbDZ4K7R
zN7+tQ3ZjO9+FkzwAlvh947NYnKEuS+juhqTJeTahPl7hk0YJX5Q9oVpjIb4fx1h
tv/2y957HcHaZsTKLHqLe5xbSNZ5IeVQj1Q2q91uqd9aDm2tpLidQ1r5pAiWDIQ/
+nAP0Y+bVpIwGEVFFL2rygzK5UA/iDvAzop6YAZf8XL1SRQFBziYBWS2ggcBpxdF
Pwax0WjyDCS6ez5uJWjFvACdT+5cav1S6Pk2hofG+L+hJTwHVcpu50XJACb4yBVH
Kvz1r2AnK5htKUC2WU249ySfB7zANQ7/DCmOnEFJLll9zL5AjeBKjwTv/sIcpG25
+juAYehITOODrujBZoUPuL6SUSvpcR7bPy+vk07b5a6cHUXbE7NjVNi7QnZ0hjeU
bzr0iEsMHhdPLMbFipfs8ibVR18E/SEFLdlb4RWZnUHb9ok+oH+7cnuRgeukCtZx
G6qBwt25wbgW4EN2Fg2LdxX4dfgnCMfZvxD1JYaWKoYW9g4NM5Np0kNnoMNE3kDO
cz6q71InLDoQjXiY6FSI12gXhMcLT+bsZQoPjeF29ZhQ26nXQYsM0hzLvAJhSG73
AM2Owz9VixSUrQnPKYWB2vb1W7Gxt1jDYkai1lKifTJlKCfx5DoE/ATxTGkvPXsU
4KlgL5N4TDb78tmNESU+r3VkV7LZBayq2UHur6tniWXmoAOKX9r8HGVHnkwMnyhf
kb49WifR23dzzBlWgo5JnxMc3aVn8yNvpk3GxdltoXWBtOjZ+spJkKm1xYx0qzqf
5Jz/YV/hPBX3mwGDxHlMM3/gYmPFFGCMB8ieG8T+iy1DuRJRutfAsgo01mKTvU32
XXZ1PO6hVBw50e5gX8vptQrkHvN225ojHAICgp4Hg6JkxId9E/8B2xRdnZllnqE7
LsMx8RD0euHE5QiaArhKlLxjFO5kLaUsOMCy5x3C7OG05faj+B8bwt6X68gLWnsR
TDbqO5B2E2mKjOsK9raVNaEM3OE4LdsK/0hbGXZY4vGp3JJB8xGJekdH04o6Gj2X
tlfHQK2ry04LZZf1U0xmUlWtJbg6sRkasaExuYsp8aIV6gAqyeKSzBgFIgY3PM3B
9jEJpzIJlm3FrpItAUOtaK2RVu7Z3Rczk7EqaobZAPoT+s3XyfuWW8RlirOov8/M
4EXkFWFB87SsITkNsUwhTz3KjhRBMftwGMvr//SBEIklL/GtocwigPeJbmkyLVzH
c7oc0mASsPO7wNdOuCooKWnXTVScTNofVE94VCE8ruj/75j278xaLSDhZeqqjtK0
syTeO3H9e6mnwwVS/WYBbQ3lI7UML07eXKJ9/ZM7Du6qKW57uKiLzjeLORMRSkh8
dDzTWPgKStw5ZuRkljNJA2qLLJz90Cy2azbcx/Ow0DlkawnRn4jX/kNhbiHaPJGR
HzPHLpMGV2GLznCMOVPlbAm2GtwMXG1aCEfNp+UPxt+1mQovUh+pQX4eWQDDKZRt
dO6jo8FG1gPj97+meLCrSbDLBA1YUK3uMImFvr7/Cc+zoaBUMEERV1WM9KauGwXg
AmUuIU2CuRDijr1PZYNBUQPR8E72yw77SxvWpG0LpZTZwx7dv7ridr6XYIpVpwmm
2vf3mwr0zcNVO/ZMxCAIbsIMOzfBLN39rNvGzai5zdHGpmNJyDd0PyPPmnG/GK9V
znc5Fb6hNIu/yfX//h1gBzepmzdxZWMmLEng8rgSLIR116XinE0CWRTYWdKeeBgo
ZEIMuv74C7XdeeROdVGwzBTFaRoJhBmrTFBG3O4zRu6aNdM8b8TxGXExB6+39oE5
l9ZmhchimQ1JI/CXIQhi2u8unObXwh5QdfENNE5wVWb7KzhpSF5HBVBNnAAT6AiP
AwvcJWt9ujM3rg5aXoyww4NNteMurkKS7Hu1l1kycJg6k0FR1eipraEiTMYhxdSV
7DGFvUbq4NYKUEHSMKJiGgbvPJLkS6Qgo75csOaj0j65jM7ThuRe++PGPx6qPMim
ugyARR3GcTbbSk9CfPO89aJaZMrpLoZLqPCw3EE3Lhk6jvAEHN2ePXA7uX0MUp2T
PVZR7jBATCQQ5rIrfFl4eHL7ED1GCCQSxiIPmwCyDc62WGOl6fp+tihWrMaaEy08
IfQpIXkQHNylJ4wg+bAdicOUOEigUNC2OWQxdCL9Zq/aR46Mcj+vhyuCs06xeB1e
3YlmTIZ5rDiDCbfH1D5L0w5opVtvH60G9jvPOavt/eOONxjVrO6DYZVlf0kIW7bO
69QJBAvh4ryJkDwm2luu72k6Yvc2WEXODMcr8S+TS7eY3vdCOdvCgncjEl29cWOC
QA6ALkL9wwZ6UuBaD8N7/mEFf/m6v3uZV/UnO5nyrx5dgh4atD8VbnAOOOSXdURU
MeXSdpEhdOK0rREYVyEpPDgYAwzvacY7U4PJrAzTxCD4xjGqcS7pn+z7V+aVphmj
6FOB6Gpe4MDhCuSb559oPxk+C7VjFN4dP2BKcvgOj1VMK2fGGiYz49o9hwArUWwg
9T0oW0nQL7e13cSJSM1aeXXOcgOBquQw+m8AbpLry8SCwre1ZD75YgFutiAAg0BF
BfHRRzFtY95MXKeuoSF8hXH3wrxzsbJ1/QPY7PMwBcxmdXgnuiuMdl6n/CETv1aA
ChMQ2coajGAF2KJa0DMy7vngY1XdIWSS4jTkElUloCRK/W+TGUzjX4j0rO3Yi6Bv
Om7TfJNK+kbn51AtQ4eZbjWqFHPIYKYlUePCEAA+SHwNbfqZrIt9/919CZVjnrDn
As5JrgF+kaXQFibm1gGtog1yxP+yhWsWDrL1RLndkdtBKbXLsT19ovnzTcUryhu2
8Mb4yzX8FEW37NRPd+nG4i50N2EdfzPzNIS94C0OMdbfX87VRPQOlEzVi+TNIVmG
9AqG9jlT8N1Oe2a5Pp6wCpGYogjKed1lMEHMjQCiu3N60V7EpTJvGKfR6BIaIo64
f5YvJPIVTiQFlBCyhHTwkFYNvId0y0CtItdguipezICfxe0f2ZbZGpLD71GXkCuB
sTuhm19Xr912TPJd8+50PibsGj89mVbYtjk26AezVpdMSInkSNelnUyxfl01F4DS
7ln5ajhvxPheczMmUv3fu+0iwASJPEaBnZt9Kpf0k1MDw4doEF7ixVVjapF/dTu1
dODOnCXRSXhdmq5TuBMOoI0IuPM4+z/HPrHs64xnaF9FgKTrFf46scIKiA0Eb31c
k+VbBvC5aKQazBX5zerz2coZcx4kv8Xwf/2wrb0giMmVIcZiSd4v5IbkU3OTb/9U
QcIwyc6p5FnhRqr/CCwvSzTL5DRtyvW5NnJYnFwX5pzoICfgyZHJUWoIGDu4aIPS
/3b2hKEh4J6e6r+WXiqZDe7q0tK0WqmhMrV9MAl+Ie0HnPNkTfoavcXD0+WrF9Mb
dkKweiHLFxs91fW/eylIHnYIcC8K7sdU+Sq0GPiGdamv7LLDddk0TIEU80wlx/l+
xaY2JmabiSVb+KzvnY/M5CcmggPCLTkv0AAiDXp7oEyd1dKJFF0Qh5JgFMAQTuEX
v7TRf/7SN5CFD7aDxGRxefqsniNp8FkVQloYmZyY4iwMqGSNx2uNy9ldpNxqmNQ8
sYl8nrFA+kqUWDMcW0MgmclHB2f7NsX55R6ccxFuDu+irpM/5E/sbpB/Y7yPT0Nj
OV6I5B2URtdFkE9goAJRSuxg7kZ32fkz/mfLQLjCTTBfVlO46TXGQEA8/kxTMwtM
CPwSw/Qnl6gYpnsgNX7gYuaZmjXwzMKgVJ5Z8tyxw/n3CCiWLYrmTiRo19EIJG49
ECMlaboV+zIS2iq7aNR+erF4M+9A4bNjOe8/+r7kfCmDJkWK/cihhddTjms55J/N
oo4cfIJT2zJZ9K1p6Yxa5P4UZEoVTyE/fDiw7g0U9vJEpE1Da4w+ehoiBsBV0GLz
Wpa/cCoWaBucVTbKyj59Mb1PWIG02rx+mH4kEeBw1mk8lLOlSTTNieMEehbeH77M
2+Ourdxu12ACpQf2vusHNBgx4s/p1m2Pi/yEpdYTf6aHLSnM1NJ8ZZmHK3YO8l2B
hazy95bymf+8Qqy4Vlr1gGUUr4a0+XZZ6YQDSYEAHYfLcOtW/MYCBWR+41Yed/W9
9HMT18AQ1X8TNn69LrXP1xkoJYzPbatKFnrgzP3Qu5jZGOxd4j67OqQt5gpYPjNE
TX9eFtZmq/0lNFiO5IRA2R5kygmQwa6Y7EDs5/oYMZWmBAfy8qweEE3u5BVAAPOh
QtKL8kDAfa2+1LAJbZXiy5/B05++dbbUQ5CMRB/09BT3hl1xzKZadqR/6HCs+GrW
CibEVJeasL55VDoriTnCMCw4gD59ZGpbBMyzlTPYWMMTmVtjf7BsfVW8mhO7JQZS
jKwF31rFhiRGoOoMqUYpw6cWjyJnt+wngcYPwWLVokE+CaLBlmfjFXAK6JkUflHO
Aye+ItJxmVOFViWhUVWNshg5wYht2HJ6BJY0E7h4EHFkKe3ft2oFJtXhhLGTuUuJ
TopmnuakhffjtDE4oc7rH8YmzIvy/WR6E1WAmzrTla9L+S1pczfjFSAAxWSalism
ci0YO4KSuhRPfvtQCKRrJuJXURcZGu1QKu0ATZmRLQNZDX9fzS2413Lm6c9WdaG/
B55kPJhgcJJFcgfuA++PEPqkfWkMoq+KFYVGgjqAV20pC9EOW+Umv9IkqM/Z3eZs
kYPtz5/HSH1S0CbLZpyAF6IMd2mmUf4Nz1jFJfY+AdUYp7JUdrwjIaUWESPZ86WX
HRoBHvQ+CrNSjqzCtQwzL7sJHRKFAuXYXEBDo4x5i2TQFt69GVVvOvLI75Ho3KFl
l+kPUPBc5M8Z4cqCgPMKnpCCLOSy9uPJ9s8mUF/bAYgMYt1WsyFuW1TEVGXyMWGi
+Z0MYylKxp8f4RVhtzXYItBp/5QwA6x+xKLP965eifauGix5J0uRs/ZtfQdwvKmS
Bqg1aVwOhplW7gQCMxn2qa1Bg0kYTiHjdAPEsHQ2E03HihLM2AJKLl/hB+4aftwV
3PEbhs+zkh9CUBFALH3NVgmd3Y4/YXB8WTNkUo6/jcRpZo2cK9cAOu6zRpV3YbxE
wNcp25XCxplOCVl7ZBgdsu9/Gaf2HeBzIlOCtX/LvETtArRp2HCrMu11W7ss7RWY
Dt+9wTAbo8UkzNDnEqUoK/gt90AEebAlVZMLRz4YrkZWZ6301ssciSp//OAtl8U0
3OS8rxp9ZjIvbGcShjGV1y1uDGz+kYV7u107+13+0zHwMdw4u30645iDWOHpLLYk
pjU2HuP0zwKXKbooUSeqFDTKodO/Tr5k9PLfGsEj+jGl3L2D3cjHyZXaRIwWkazv
DBgyzda1Dg6FnM7ROBgPIIbOapJMVtl7hnv/FeO16TbviS/pOCp8GgFkl9elW/WM
5jn7e+IISMEXxrpgeGvtCFG2aNk6NyI55R1yclmDSS74KxN6Idb36pvuRv8Q6DRG
NDS0jG0qbcUovqlXYJSFNechWwxcjq9A317FYOaI3dfS9Jm3ejxPat7bsDIHttEe
Sm+ag9C8Yq4GxNPhr4fRKtqAFgk9l1Klm1bugdyuY3U/VAaQFaIFdj4CgGXuwRHT
lJFuwcieAnsCr8Uwpa17ms8MG7Gl1BHuwe/UAFrVhvzizDs4uQXUlljYqN9cqwmR
aKRR2nQ2kSy50dWWy0Wce7odoc2nr+JnLKAJxL68J2VHoGKMM2TVuv+A+Q2FZNGi
/L60jvSuM8tObNz/Cvp+nYSC4AjUEFoFf8OdcteDxActVeRvvfQU71yzQvkSlfz+
/e36OAyr8uSH9Hl19DCxSps1MO9lpAUfL9O0mCAggpJ/A1ZApxPYNjNC934dd+0B
UBOeFktGXW4X6ugqMGwuNw7f2gesdaqTUyP7wikDTycjFsuaWpXxZ4iHmfMvqeyM
PrRrRpme2E788+tztrHFBKTeh7f0i5pmNtz1GpHttlZrB2DflZywk3EBUg3o3Cuv
sjtipa8GyVZriOMPfL8j6aNgHxfltZ9rIi6AXZrowRfe3n+hzQyaOLRgyNIMv5+d
ZDIshB5D6nzk123WFgc/f+ivqX0UPCQiQ6KSvJDTNso5o7nWgveByo0CG2tbLsRU
R5Ul68Cg5vbm2JCEKgLPxJeLedF0L7g7LnHHR/TAnIdZzQLbeIoVf4/lPnw9QZnE
J2npocMotcArHBm2sE7t1+yfsmXLZcImMoGAXzOFmJRdRwd0Jo7+qYypuoLzI3kc
dLBqcuyPQAaNNB220fETReS6szcr7Wtn2tFcHhLYjoKAkL7hTbVFnrLN+wNkI2on
0ed5MGGqxFE8F6944gaK8cv6UQaHh/zq/ipqeT8FWWnJz6dtxsnJGoyu3ulRnzOT
UgH4hdQ0bNoJEYJpcSHdMGW+WG/vJc2FZCaKTtr5cnDhSgHaZTaZ7jLkPn3XOmF+
d4fPOlKd2ErzZEK6bB2z5nq0lhIHxi7usSWgt6zwmJfbPMSjcE37O3ijHCLVkoLQ
m6xyyRBvsLYF7z85RhWG/CQAo+X2XhQjeyAuMrNax3COqzkIMr2Pgo1GWREW30G6
vh3xuJbFojbH9RGQp4QaBczXpLlKpk2d2ADjIWF72qDfOnx2TZusfD8LSdT+4mF0
8vX4/DvSknsRVgyjzCwP/K/XUFyjZZZEItuaQg1SmkByJq89bioARsD1cvA6d1rV
NW4I/hek51SPINf3SPC5h7euLylBRIKFDABdwY6tfR4KQ78yBgyIN7SGC2bRLmVz
In76fftF9HelR92t4qlc2Bw17hVLZhfNiCRNlT22q2Ir/sCJJ/paH8DCnEf2pnsN
XcBxbeUJSmyvwUfi7bF09W4V/c9lhJLH+rqrYIhSaxP4BNPjWlRd27rB8rrMXSw4
fxmOSF3n46plYfo/yWy9Tmmyu9P3FON7OKY2/KbPqUukHudB9pK8Iz3VcqDsvN+M
OHCp1vQE3xDRY6LCcN4w0SNTIxtxHlWIRWWZRAZBaxeS28IZ+32AdWrDDP5GYi9t
Iq41mxhD23jzEKLywLz7WSi05rPq9TuZ9cORfuH8xomYSmCiq4PGa1Kd4fJTd/+o
FWjOYtoWHt1mdL/vvG3WXarEgm7hzcjGLI4fgGWpdIWf9HhQgd1drB3W3/46vJJy
c96LWeEzCHnne7/6cuIws7p1JrscYVFyluLoPlhsWAMC93lSuHgNUnLmchQEgYuJ
dEIl927+uzUSZjJ2qI1iXVLwJfbV5Iq/ejMS3MqJB7WYGOkA/4frfWvKiCGrBkOU
a2v51K8VFswn7RDmFaaT/Ri4lLzmeR+J4k16i3ymyUAipDs7CmKJ3lO9pqAmOQLG
6vL6HL5bkmCh/ypAftP1KR6jDW7QZb+jN2diVsVpcaD96YPP5HHojFBrXTjRrvw4
ddsCqPrHN4HBrwhTkoanP9isAE1/wlxZP7oqBLP8CDSQhurQBorukxX3fDcShRXS
mMqTdVvyFTWpBoQN9xdqwOrX925G8qw2JAxR6FdyUdUZacmcUd4yFspOaNdUCZqb
kiNbtYHJb+153b4svHbZaCV3R1i2YjF49WCRtH1fnPjgUXuP4ihEG4UHI/t+nB82
cFJyINzwNnmK3QPPkAbaKv1TEQisPxiRF0aoAkR56imCNHiPYnGeuhHrelSSTwZB
uRGJ1stWIfEC7ZN7KZ9larvhm2+VBfXpvLHZ4j3Rpw8RshRbmPqyAiggLIFWCO4n
Ca7WOiV9UqlzlaH8iWw/FwIiH83PESFsX1WSLWyuY99yCmsGfwqxXLvkHSUJaST3
OrVOE1O26gtjnlKrclvW2Azvv2v7142uES6KVXbHl/olQHRvuCRdvUtNV61mMKGk
2JLP5yWoutdjdia+NLmnrH5kTFyA0RfePrr+fi2FJNCjFZnNtjDvvi/fe7/GVwWO
yMdE/j+la4z+AboJCzeS3oC0dyfwlOAOJX97q5Xk14jy12qhp9oV3cmEqz6m+LhO
BAZZi38xIDjU2Vhx3MG7fbzh0DQSf2NtjeRWLockc61ydcE3CXupUt+mWbNTnqf0
SplrjU5YQfWgzq8TCkCk+3IRcPzhY9fVXjXF+Whc2d6Bq+XPgWC1HVPZIf5qDWTd
vAUZM5vjfAtXW9xSygML6FOV9LrIVQ5Duh6zElurq9RHzo9BVBj+NJOq3zRLTH4r
IJylHYeFCTuBju/2EnW76nF62Qx6ATAyilb7D5TKdatyuJC0e8vJkW3OitOvqqxn
527x3/l2Clo9lR+wmbXZyoV6RFNjoBgGR8Fnr+hQ64BiudlYfBOAK4LW6CUkOiKY
JaH883sGYPhb/WXj7WyFoiILet/v/077/wQuR9WDQMBJ9fSv9bcpQ3oXlKA8tzFy
Y3v2D5+7LJkre2yYYoV+Ff9lYkjBswW3uLmWETeRk6HcueIsRIxyoMXULIuim+U8
yj4gqcsjf1436g+erKPSZDgJFzWlElUtIAx3dFmQT8zsqjC3Rj5stTpdvo6I2tQ3
MUQ4fUZ8006ZuY0jyq4FSTp8FAjMKELm3AbJ0pczynTqOoXUyhpSu/3dPt6oPyJs
93IKwsF8tMtzLi3BYJyWI2+aX0br6L/6mCr3TFHd0as7XFJf/5IjmP5Qgev9j10t
wf00EHqZwrWjg1Hcfv2W7uwmMcN6e1zchsTrcbtKzACV8hS4ZtGMF9HkPUe2VDa+
aeRH5huYFhXrA+ox1xqXUJm9z7ZP3sY7/8vWNVZE6HiRIlEzcbRNRprRq7rwrUMb
Mpk0IAIZ9LcfliqsHlEhCKyAIMFG/qJjj+KEQvk/YG5bGmWSsgydJaNn6atCSb+Y
I44HEGzs95k34z5/wiPJztpW6m/vCt3KBKi3/hjwLcLEuzR324dtT4F72T6aG047
sBlvQV0CPmJASyHlUTNh+lkgOObszLQxRVn5lrGd4Ba0WUUkOIqDPLC8ZCJh9XUy
VxahWKkAe+ri/0QeXHod3CC/RTiJH9y+PeqZBHxKVikoTGw3oi2irt741tB2HQO5
B5pJtLnGu9lOj6cu2af7L46xumc2wH+UTtUs5BCR6O0Y9+WdQqk2DtWkcG8XOuV3
LXbjd0TWoKcDVaZNzGXO1WZpkSZlzbBuJ5rJpF2GaaUKYPiSNpDvbkrAyZ6pUg/y
WmW/vH/1/WwrJpo45Cr6SjzARIFYxKyL5y0IziAlkXhkg6391nequhqBUgl20E4Q
Oo66x66aCDOPOknSo4mQviRMEsn7lpqwXyIYqbCrCGKEevc/lDM2kzOldJ0KUjo6
kfgaYO8GAsrfW9PEmsUOCBKFdZOJVD3VIifDYBckZmt9zOJBLU10IoztFs5n5RHv
ug7RLurGKa4kVzeJlxF3u7ldkbosB3nrGLZNmW7XIFrAx6PoyZ7Y2lvMOiipAwQw
MsCWCrXthX9OQMihIcq957FQiV/mAkJBuLY+9YUWJUKaF2ljY2L0G5i8DbSowejB
hAVc1pK1B25suMyV95F+OpEE6JHwQDN8wuk9latcMv7TjX5UA4gSh9SHeZ1JfmeD
Gb397IG796B5dlYwAkqFZl5fGdAdT1PlHM2Np9DtqedBcQwbn41RgI2R/LBK2JW7
mibdkPozV3qvZTYmsQjNgW0iuGcRlriUnt0aW81YF4Ve8wMsTqsTX4amR4jMu1Cl
9zih5gaD/AErmmG1V2QBUfeeZovGs4vCuaq3na38oEhkb/dE6771XCnRjpPXjE4k
FC3qQnb5tnbcDAxyHcSqYSF2LKgwu7azxMoHd5g+Y9ZbbyY6mpgDwqP1mRH9iFvn
tgXr1Q14r/lfR71stMfb86lisULPmakSXZU3hcjfcRVP/3vq93oM1pI1Lp3oByrh
9vsuVgg6kVGqDOYlptYIkShAobpKY5NOBLLJgJ2ICKJDp7w/cdXvFAl2Jjx+W9DI
+lh0YLbdQhIbDxAoBQg5zJMWPW95uftW+58UFxqG8jvfCMviYwf1YBT5lNQeoZ56
tK1yzHrMhDgmkKepzlBB31JguQ57bKxB6QOHBRi2Z/SIR1Q5Fg0jIT8nV2QEeaS6
jwhgYYmP4B9Aixz4Lp2xMhx+vDGUDjSTMO00GS49nN4B/ruaM1rvshbWtdTfO5Jm
Fj+7F7qjKRi4brhoCZSlt5Fw7x9QbP3AjWqy9AhUTBGwD3Z7EKG1Fv9FHaKbyJBn
smGg3sAblB/3Jj4KXeaWLiNxdVpfInK6dMINjoWzq1JeTlWUlgrStqG3Bg9ct7WE
ofrm6YOeUfbzRKAcZ3xA+u4UaTHjV3WCtaaCQDmSls2jV9VlpYPD58JPpZgHoLgq
Hqj1jGjsGn6zT9fVRPgNPvsGegOsWSuHHrhHl8TykCfdfZLoFb8rfq5ANs0QVl/k
RJ1UXftUMaVOiLDucCOPetmpUHlV4VKReqa0gBoRi/IDQ94SZEqRQy9EDMAlxfaR
EOLmM4scNoG+TbnEjclhFUr3Hh9vXdHzSsSu087LoNQpcm7iSPWMPVVQiUQxZeM0
vvUjfLHVmI6ojo/xshUddJcM9zz/pG5VepqMnUM5XLM/7vjzRksy+XyHx1vPHrVE
eW91DoGagrhHJcVAP75mjSreBRukY/R8cXyFUyb5WQK2167SnM1V1bYvbXsJCoUe
47LjMTePARGQPDVEvwKnxJFLTSLHq+8qj1yxJ7RK53cnPcSrb9vXIkLoanbJXUPb
rJoYwevK8yQW0dSV4qb6aNMFUAxBLQ4ZhvmGVoZAJIrfkvDaqpTctxbeo1zWyrb2
VNEf8mlQiEVr9Aqa/yFRzXmV/rt1n7GJw/MBjIdzKSyUACSmcSCuJlBOoKAFtPAg
R1+RiSuONrpifalhSdIxq6dOUM5UnPK8Y3OBnFvQA3fk9Z7yEBeKWWVZQOeHxZmC
MIvOetRPQ0W2HDGlUOkTu1gof5CkGRok4lj9rYyftLrS5IHbwo3UYtd1YcqOjpfp
TJnDdX098epH8NRPpEQhUorL1pI6S4YOBC/r/D6o4bprZrcVoTzVBAVeH/Knzr92
dZBzOCEs5nU154SW+sNVKCcZZKAjBqlG9+rKaVwOrShkIhfSqTfpD7m9L+L8qqL8
Xlr/4CGlIXKW1clRMSFMBPWua4of3JQ+2SNBMmBxto0YHwyIT2WkOpLZ9Jx4Hrrs
2sAqdLnnykSebXvZZcDKpkRVOPnpMAUTeghWGlnSFzMnyddUw051bI4bD6MmlK5o
En4yXghxrRCdWZPfWfZDpy1VbcYFbMtYTwW+zjUITdo/gYU48FJBy2kFBmRWpxeH
dsP9lDiu9FhehciVZ4H3Tt1/yinP7wpF50o3hGeEtA2CCFeRllKPvl/uM+z5dKu+
uroK8wcCi+NGenQR8146wgXyu2RRGtycuIBapW45WivzRxirUo9Qs4fIRxagLHk0
h1Fv4VSdRIB6X3g3i0PXEi0qqSbSDNRxz5fzNQeIjkusWf52nPMq/veqTCrJPsoJ
+Da19aDW+jLsqhb6nYUCg4ldJQdZRAYVuVwo4rr2mtyLMS73Q1aBsoSgGfnzWI0j
99GApD4CXguDJgvc/KSyAjCN706SW0rxLfJb4XdykiLFqVeXLZXVvuZZd3jKksJ2
MlCGNyzWhJlxXTeJX88FBDRJ9iRQuiQgX21zeSGaeO7tOZX3tLkh9C5reRdByfp9
XUYLXsiFYTwOU2PFdBt84jc24GE5wD7pZEWVBkHkc2Kqt451p5C5Roye2PDsgr+2
ico4wN9ad2DRh0KAZQZ0oyXAqEIencATfl74zGJlLvu6Li6QUO0Gh+Wj3u3wb6QN
0Bzlfns/kyoNoiIe6KJxqMWDJw3z//rv+5QhP7MbKYA/R/T92ktOuE+PK4fN9X7r
haHArO/PaQsBwFBmaEWSf1e2HjdI3Oda7H2QEvMsbaPQf3E/LvitI7mh+8JIXjzc
c6jns9UQkwvILDkgvQIALeEBI3daYYmt1ji+5TrWVSG99WlK50Dh11r8ikEJLgIo
ZBMNhNtubjR3TUPp+3LYiILqPs09Gj9y80SXmhBJPi56owbldxmgkNZUsjAGEkdm
y2kam30YX4frReexqIP5wgSIgMWFvwlgPU5mtI9klR4uZeevRsQbllwfejEPNZ2r
XYsxwOU3YQxDbzRZ2RpbkSNJgyDgL0o5lJ26q/1Pc0qcu8IiH4bMXwFr2yzn/qVj
kA9F0XxXetlpbxBDWxpfv/5q4I8bImqOhA/sA07FaoEssC8Z5iAjLKDEp/XdlE4v
R8ZVxUMrphvjIrbkICQtGGWGjwXGg2us7FYWmbS1C3yLfYkJH3QiGp15tKt6rBbO
1Mx3928e3R7jkc5URos85+aqZKOC4x/BNQC0goCv/KURsM98DdjiqQjTqq+EcdW7
niv8W/BsO82y5RgoO1cGf4hOze6sCReauDMVhVVU+c7QfjfO0GElhu25kCopo/nC
o3VmD0MJ0gwRJs2nmVWYkgupu8o/q/UtuzNPZ3jObuuhm3kLZWO4w+6Z1uwH1jqS
iY9GdM1+wrSm6EmS/yszwbuy8mNP7Sl0QKnzxueYURLpMSbqSCRyO3iM8q5/PUO2
dXIKKnVvNNZrLphRKKPHuoUoJh1pxkAROF9c18Wg5yp9UwtQIUCk97bkWIQ9s3ew
pEPDFxM28tx0hvNZsbksCN60vYLwX9qB7FDTCIBaTfiU1zUlLy05NTllx28Sytol
sPSIFXppQVQm7x/wXmTt7DV7yC71q5nIU39MnhPp0ut+3PcB09EsDdaI2aGnXqFn
0IutH8esm9a6J0cNpvHN+kIFcSPG9LE33VbvZlhAD5rNpfIRKIOMkambKanQmnmI
wTIBuiHupTtGWZE9Rjzyrnzw6foTVtFr5B2JmlmLIxJaMQ+o+i4JYUnpKVn1urWt
0KqTGAVi9Z93ruPF7w7lTmuo3tOZ2KSHgv8n8g1nuOfbHiee3/z3JwCPGQkkpmPv
3CunBrhbautD9FzJgqfZbtbQ0uCv24U1yyTgrac/laxztxARcLeYYjZd5+cHuQPq
Tp9gZ//JzzP7Ze5c0eIxnsADPH7GUCXc+aqR0E3gpkh0RiHP2ioxpBqO8DY9jzGL
HN5disjm+LhHmys0R67w+AmpgY8MFKhS5Tlf1pyJ9e+2OEPionP3D/bdjPsNEeVy
pXfsnyfCB6nVqyhHNp+f4IkwdNVozs14rHs4X6LbLToMZoNu5LPqXKEWVBuZ7ZZM
2E+m5Zn/SM3O4kHw2nUixfFjWEbXhfIi1UW0bcH/f+Hn49WnGT4JMSRaWpxBJPsb
sLZVjiCBIHLXSkmUoASuppWAqe8lleGYF2PydiVoQLmANOA8y1BBf4IKjKOHgNLT
rLj4Q9/V+j/9KJ1fE3R+jieFbPDEKsyPUBtMXIEY9p8W7BK8dPnMzVOlIAPdow5h
JFtwE5xgjbLtbvpR/9P3LmiI2VgRi+VGTmr36ema2khvkFS8P6uG795EY+TG7EZV
anJ+gwMyQGKLps/e0MNW5sOQplSPdvdTAw95PtqRrDAHVX02hRunP5SNNdZiPZH3
vYuPWQe+om9oOKwjKvYg1gqmoTJZkRMjdnAzJa0FhakrXFA/v80OZBdaMyIVFJDd
zlBpbj4rwmmy+YH+Q+w7WNVQNgqaB9nn2W9eEYncrk6TM1TvaELmcPLdHgVkKhdW
UH5PNTIGubPWXbLS7HwgISPwSFsBJhGoJexJW45uWhNmdyHA7IoVtHQ3hqHm5OLr
vfOFbF1G6+Sj1OhS2fGWM+aqH/nuKtHxI/uWtJZhCkE5L9rRSRIgRTurgg8k8SZj
GDJCIGZ39eiuo+LHGWQbVQ3K8zQ8UNTijpRbycjSx9H9U0rwR3UypwZR6330MP1e
iFZMTvhD14bS2aZzdr8ZvPMM6jIME2jM08NpurBjEM3js676P+nn51+jSUgqFdfh
xU+UG8U3p1PXBwGJWYLMyDVZDnW8mDshR8lZ+/ExwSwkE7M7enMqwOu1u+NlYSpo
AJazGt1BegKE+6hymmmlFhW/sE1vaig33/iJhmXxgGAyuHz06mbCPizSujG9Ve12
+aucfNtJnIw8+dPTH9ZxjHbGV306DmBexLQPHE6zBtqbIUyN4DW7ghOdImdHerTW
iGxR8anymHhSosb/qYxxCyEoNN/oO2OnQR/TdF2w2RXb5peKzhMCK0QgMERg4k6H
Iu5q9+dh3Ogh3JnVUZRWza7MYLxlufv7xeHGA6A77N3BtA1WP9rfInqjw4wNvFGi
lloB0MhzuvuG2KNcyrAa3Sgoum3KBkvd2EthCvba141+eKhST5THp2YnqhA8OoDk
v84Pu2PHRmSlSPHPaBAFVoXnSz0eEslRP0Rqb4rNXDqqi1DUAMhx+XClmY6/sBF4
gYOnomoIrbERmxkLyRISaVRl+Ea49RFTNVasgMq3rv3v3NlA4O95xE9murebmBy+
JsPZ5DG1N10JOtPGLxXafnl7yTdaPmEuOPedEWUbbqV5ZMRLc7wa7kCnlJcbY1CS
uxF8GoRH4g/w3j0op/OqOm1x236rFpR0szU15nCI9SfFlfsQttj6jiHBfz0yho9d
6k0ys41pARk4cHXwViAzzibwqhzD+HMPkp5Rb56aqGJs1TMEIQeMrMq+NM41xOwJ
5DOAebjXQmPc6ZgtwDxoEShl1xXLDF5DJocb73K9MRZuLpM368X3TfNt9mDnhYKp
tnjObM6iZOl/p3nxvPl3rixP3OoabMwngq/2t9HAHCIKvQhxufTPmmonzB/YLPkW
2CaxpDrmOOUlZSh3iZtpgJ8AmmMR9ULmzr0efziUjJJWAAQlX/t+mU/XXlryadfJ
PgY1GnqtfqwxKjNWT4DnmXGj99jzqpMapdOJwTToMm22E/+L898500VgZnG0n/9w
ud31Y7zM+avdDFSx+UakZjYda0BBJZJQv3d9BlevHxKMGA+Pgg/6fagsMAV4zQaX
LkQ4b6gJsWCEnrbcSxp2p3VHlrL8V+ByTjxmah2KfayajF2T94nvBqcZKGUE7N3A
JrN5DKCWTamdlUw5kogTpNFOgxUCWnF+BLi0OL2NCNGa6oa/Xg9YqbElYW3HZ39v
wM3qhVHt2DnTGCbhmRTwlkRrpu0+HjQK2AYwJN9jel1TBTX/IunxBwhpukx4BtMB
witN8RZP6MlU4HRUKlrKUws4d7d19tuMK6x6EQI+wrYDiRKAbESNDcY9HzB6mszk
TquqPAuSURsYlBSKuxqjw/Y0Dja0pxtyMsBfGhLS6lVIpMXeq8tKOuFBRkKjgmK2
yuz+u28I7YKa/Eyf5N5dHrLhkgmho4FUj3i2x2koyDvj8XbOP+EHeoOzYMa7/shc
8fauwmpTuooQFopopM3F7yckjyRLDkH5gb1LLJB38IHcpBd3aEkzXPm+5J5VilNQ
Ih/YFQD7sEnkFwywkUW4RyDD//2E6xiDe9XpcydI3IlJYw3ycwaIcCKtLeLbWCVM
8xds8cLau3vgOijm8tU31UnFkWyiqVTOdyY5NC4Cyb/hmPz6Ydk88qqLfDKcbSMe
wZvVyV8wm+ltAMfF6zgCADccVsszAZq961ZiL5ZT5fuyJgda+K87+HfPUvHxiCw1
/UaWcbQrFhKiRY0b0ut+dW/t+0bS27+qKGzM304myKst79FVDKRJSZU8MyVMVHAi
EcQwvuq2vuOx9l3SRaMQcjISlDb7Z235FJT0UsCUKoPVwBrUr62z8yKg3hQt+NBJ
WyI48hYpEMt6R6usVjytU6VwibUdVlveorArEGTlhv/VAcdqXNVMCk0Thc1PbClJ
UFnarxVtW1A0VYtp5f5PrgOv6gla92Q495Dm1veukYxVAIJqdBvqMUl7DEbuaCsk
42WkWqlbOszG7lrrfioYlSDS72KweHdDADEPui1w1mpLnMSKkb2T8/AYvQC36Pt9
IEvrBdDBPWDWCEQvEJLoiI+AbYD8lcK4Vk6Tffl5sqDXntSJSXa1C41g5jq0esj/
DOi0SGCtyCTbEGIMQ9f8bz410E1jKiRe/YojzmPp/fmbPIr8d0m5KEC8SR48Ffvc
7PwuFAT8rFZ3NYVkDmAKi8tp6RQy2pzLni0orBtloMo8mM0//PJN+9bNKD6M/xRk
gCEVAkyL032N+y4xGIDZmO0PVkg7V/bg1oxlWGjMjEITYLlkZXg6Uc3isRkpynFI
c9XqkzUFW7wGm/ejHCdSnU5zgEaN08NUKkzvrX/WenIEHvhZqnvIZU7Ke3W5YTsi
ZtRc9QUkmwa6NoNUW2EdR2i8zQKABnSsWxephtPnQH2yo7+cqSZ+JNnz6nQsku5X
fB3xg5+cxYCj6GWIivoYjtzTLU/Ks4JUEQRUKPaxl07KrlVU1SilwLqf3znziqqU
0fzs/CtQnWBPwpA5MU41KtyzRHUaurujJliZJOrxhheZy6MwkgzCR/C6FLOwb/+E
CTCLePank3fe/xhLL/D3qAlTzyIPPBszdMm2W6rP1kxAP+0T6fPuTgUT8OUPaRHG
ITYFLkdnhe5OiIy9U7UP0zb/V5787HRPvviBtGrnXq447iiUF5OHSKobl4w5f3GX
4e0tP1Boqi1hv8G0bSKwSEfzsI9xeVufjxRklGZDMHhl2h7izFSVGkli4IVtt54L
UK2YlQXHJEIIU2BcBctFByjQM+N37XQWMEDL6yBzJSZSpjqcj1hhrxLHzreDH0QH
Sc+TO7ufON7ir08gyvurlunqPGFuiCLtnpoKxwN7+FvC3x5SpguJmeBjmkCco/ho
Xgo/ecb66PtU4oQC7E6nXcSiZYsEh1/yOYraIcjcH5MYoGl29Y+2Pon/MhfZ+DeG
eOOEBVNI1dMJoYP2PNRB2Al+Ocd2mgSeusLAU48T4ffmJZJOMbICeD/BM6wrG+wI
4dIJNE98NlN9CKqSGhTR1kVcFbF1pPPn36TaZmQa1hRPeHVSqYqQg3exFsW1+a/V
J7Cscm1KVl734292gN7BjN+nda3JJ2QcEB3/KRynEay+RumfAKWTDB3UDBa6YnED
/Dhn6sfksdaG2kkH52ayAVQoblPG/xYbhNKSfMPk/uEyRZKgkWTSo2c8BtEdaX0g
9dEKgzwayBA4gp1YUAYHgC23nEKFSWrgmK/4XrYk4D4tjKDA7eb8WJk8YCdSrO9h
0PI4h87jvWyj9MoWA6NdIDow6+Tzn+7Xmg0RXAZigYJkqrxMsQh1zpCp+VnY+3KD
9tP39X6jmEg3jo7kEC5nexqIaAEm4lszCSNUlLMJRCOJ/NJUqknz11TaShE4H078
uxfL00pd6ZBf9FP2DtVex8W3e7URoUARUF3sNdbPuLNTusUvkPWhSjIqr0e1tIZt
lUpOTTXiZSFGDPTsxgjoQuA6TN+ti1LF+dIB2L3x2NrLl3t186Fv73yU/4/kokCn
u6jmA246PdMFrb5UZmFdUdkTLri28SlRiWY+D10uaSueQoOdlMhb5U8HtR4pXS0P
hwxTvlv+O6/BVKBKmZzd3aQFXDgoBIgO/IEA4yTx7eSa5Ai/MDxt1ZEur8TVLdrE
/CLpHB3RiI0Cwp9+AVLxCbzSfOLWiei2dTEzZq2pLAKFzXTLlB+98xWInLlPr4KM
MHINTDICDnhQewt3KTgbWzqG3FxvUsbAD6yBt3aDm9i1IH/2r0Yjf+B7i/T4AbST
JyZ36oNlZE/nx5m07kinLNBE9UrChUDfuHCymxL1UtNmpFglJETdWr2dq6xrRFsH
8Tad2RESftCbgG7CyCGCjGpHQNByX/XB4AdlTvl0n31kIwrSs/g3f8imjdqd1Cw3
0iCyN0+4m8BC1dDGzfkcCuNkiWYdiVHPAlNrLeciN+Kwy+yEfiMiYLl6xOQRHMH+
M5WUop/O0NATQOIwUsCmbU/jEZTtnavke6q/Xbsp2UGIruRcZOMDy4ZV+DrJ1K2/
vYQUyfwnl0uKydJUsxKhl1tqAGl1NWZxHf9WkR260879xhUFbiCEuznVmJlDy0oP
BTeX7YdqAu7P2LXr+mqsqph9Bgyh60FQpWdjzrh33pubEQY3xD3b4/YwsNIgivRT
N3y1OntZgd8twTHx3lm2cZIfJxi7uTTj3/sxNkAJLNetADBA1UbPvnaqi5JCLB1o
p5rzvCWY9CIQV6WIgBxfH+VB2ruOXQKT9giiR3ipIi+aGhMaLy5Fij1QlhXjNZWv
B0sbhDlBEkwn6f7v6Wr4W/xa9h1kPez4XFwU+kVf5hc4i5aqwC+hXyjDKCHYW3LS
x7jGcK3eZ/Ujv7ZfQ2UM7XV+m3asrd/4RAY/Pc2p26eZ94imVL9rdxgtbYI+EXOr
X1Z6S8sP4h0RtmId1i5MerreLP2FMW+Gr55tEuKeo7qv3xuTEZw4BRI0FJdM9rJf
QZ2ev/0r5T1IlDeqzzH/X4yeVAxxhW9lN7ZIDa3JRAuBtrT2cJzKVu9tRcmg4rXj
u7++vdLtHj/6KJjLFP95JjQelvLmNZThvpnMjoCes34lEljtyeesi/a+hz+WYXzO
ifXMciXuV/rlHqGEpLjmnvlMPKWhIB2bcR31Z5CxmmXFZNjC5WO0kqpXYtTT5Bif
WSnsQT/IX4OT/k/JctgZVmZf/gbWJ0IEXeAI7A3cDf4EVofenAG/hBBUGbXJ6mR0
Xb7teqMIHQtQyvIzCLMaIRTLWz/AoBQhCPhCr4h/bp1Y3Ub389xPV6REM3oHN2cY
o+wJpjQQd7QgadNOc7CSa+6dSvaxDu5WE23Wx9lQNWPqHPgdDmKJLV/V6LgYMVZj
w9nJGgRRwP9lxYuzTuvzAkmjVgF+ijawusZTnvDcFHjDbbazZvFEU/RL8jBGYBep
2Z1FkJ6KU6pxKG0+uipoTGV3N3vsFv1rzhT8iLvVAN+ATwdW3FnxhdO5gSgARfVp
NtPmY7T2YhOSbOOS7lxQNy6gjJ/2E2A2qzz1zx/defF0vzsdViCD5eWb7827MA08
AwMpvWQfvZVsz4gHBto2cwdKg5axNqnGKg5p2PX45NbPAkJxmUCACKY6+qB/M2mM
wOk8UmiF+apPitvXKCgx7Z/ZtM75DCupka4PNtD0iLRMn3dh3YbfypfO3k3MsWYi
26l5hJhmxmLSmO7mo8NAn5zJ/Bn5QMvz7aQP2f+CvShLVMXTKRUnsaF5b6UnAX3Q
0/5cfjS1SNidjJOkAk+jjkp4zwkFOSv82wo54o8Jvo4pIcGHfGOJVOSI79JW7Qh3
6m8xVFKSJLJDg43PiW03WlxMSGnIxsV0GCS9cP7/SGYCYxuMsTnBZv0Plxl8mKyi
0Vwfp4/sbrX5Q6I08l8OLdYbtNse3sI1rEmvRDaz1qlks1FEjNomJj8C3JoYY9jM
d5EAsyY1JN6ZiKJ66cs+4JpvTp1WBI0I9LyK1U+cEXFkEqOTM9S+ql21A9UpOJym
BqGIIqEapohtrLrBz9L2ivWdyJAm5FIriXcGrxy650v5L/8KQsgrQ0ctN/1Rp6/i
3v1vOAxBmLKr2zXcXR8PeOkZ9jO8w/OiTTByA5P7G549I+NTfo1wnhGGrI+pxA82
nSYilPNds9HPbU1Ys4vNuY8ERNpscNKp/lOs1XE51wCA/PP96jf9nVZvcbr+x7zv
PFM3Hz3nGXs0ZSIJlYGhqSmzq1H8UETDDj3/9b0QeD3Rz391FNaZhBhOXcxHSRMU
4bjsV+gTWD1MhBDfwnNXplTTFTV2F7lMZvfO7S9wVNtj/bPkGyPwZxCyTvVSCsxc
zNWX9UD2GyhlyY22gO/zPo7AwrUXgYRfyLxtaOEsC3W1V+tcqFqByBvPPwOFvhEp
0K7Woy+Fk5RJpnX7pmLYEOYVDs4ShClh7Sg5T7cOw1ck8bZHEnSmvikf5omfYwjX
Wxv3hMnaX+96ASqln7BWCRRxTG+xlbfBpIOLK+VafO3bW88GoIVdZgYzI0ib3e7C
faVToxteYXGqpeCXnl6rb8VcpqhTDRX2uSth21LXvR+dUFPTBJ0XR3bcAFluuKFC
5UWnMjYeZiko+UT2sJskITdBDJhEj+wG7o1c3lnXalnJs29kQ/fvurzhB0qp9vYd
T95GFwsvYChjNZhj4xEKtS4ylSiGgiZTq8YbHvDh9BR3Js/m/qugJmoFfd2R8kWw
tC0wEPMBBgd32/c9WGTVGc06m7bSnF4YZVIx10aR6Idx37LnmHNz8A0E0hPYxwdo
PJ8lwZy2JB0qgeUr0rNUBLf5BUhcZqxl1ufhswONqMTJhtodke7j6ZlOoQwcrQRA
70vtTryYyYO2BSPcwoBAQJyjKllbUIiqKoYBe24NRzb4hRYmKpGDcMgHXfiGvxdq
VeYzBNN0iFxBBizdfZqjy/x3I1T+K2XOW1ymmql6MQy9qxhkJZ+r5fInsw0vosMp
VMBdct0QOOFnyEtYb9FSL8lJUFCGusgOPzIcefpVpj8kdcHweY69PPK02hJXkeqw
SFGMAwoT3ICjdgTYZrT0QIQoQz6TShoixCh+MnezfVg0JoE0E6adp1DItcLHJaPW
/L0/RCxB8MvnKP7Bi18u/C2iayR9P+DIDQxXLe8zurCLSJHg08P5oU1Fe4W/4OZC
865TBIpW1oYMlcfnb7rcsKoRRCMUr1fTsjZYKqoQEEUu4EXGgx2w+SZk+nKid1ef
IB+agFHkgaXEQzo6UMCjmsgQnvdsWNnVv3q3vpnUhP1TGkkrtjLk8/EyTsgD0CmW
fdrNon3bE0tiKqLwju/m1DR38T2q3h1JLpg7iTeS5vfkRQhuf3+1PSIsTZLxhQM0
j47qoHXYutKnGX5ZviVKE7pibgrvUSfrE1PxiC/dbgsaLmjF9GyEfkIAlJUsO2bW
29B3zTzRq8w1ooMnf6J/zVmYzyGh3k42zP/77wO0oBQAVBhPnfaGqpHVIuxH/nx6
isYwdTS96W4fiEb6PjoBi5gw5vQZLBRW9h4WzKyC2VGQyAXK/C/wV9gsNv03G5B2
2xYw+cSlgq1e5ZKxHskyd2YR9jUks/4yY0XHYWlRjDl29gvYQbguHu+7TD02xW4v
pfh5NHAF/3oZIfdwnj76EciP9np1rELelMSVvOBiBLt2Dp5jwFTIOU0VD1ZKdXsn
To9QfdvC440TgnbhwmMV+/PXTjJQPnZP/mXg6SmIMgfWF/KnIREyJY2YZ574rmXe
5dn6At8GMALA32LTrl5I50bfGJwnoUnPFJXMU5fUnmczdJC3foole2ZH9ira45gW
3mEzjceF9byM4AW71WLSd0zMo+e56ApqI6R+ltZZ6BkpZk8RWlWiauDmkUNhTIEh
eI3Es9sEvdSSCifjoPgo5T0K6IYqKBkAVP26uS2p8N228wMBHwbLfE/EM8shvWIp
oc9NJgjbpCffap8iz7g05vbVkE96DUpbE/lBqVKbIiSybd4MdULYW/RPYpP5ZeSS
LrPBr6gE0JGTs/+kCv6X9I3WSFg8MAnSLbjgnvf/Db52Np2gPSlQTmmWJAEWXDlw
Y1xPU9wDiNYvBR9/ZHmXESk6GJA7hjfWPUUjl9RdXnN6xVYyN8QsmB1PIOCD+/Dv
9Pv9rf2eh/UqcilJeO4U3vya9NwKtAtyjZiwg9CaAPFy9iWSFnm8QNmtodlBNW2p
5NxY2GPLjAfqsPKJa3nz/87NDVK/rrA93jdC3ce1gaG/1iIDB4dEnrJZ7g+8IK0T
C1EBwJnof/Ge57G6uVuKsRixwaH9qD8r+lCs+iFg4HgCUlQ4pUEJZJVyE81NI+5t
IegjVs7n+sz3oFrH25ukQlVPDTIumAeKrU/Oy+1X0HkeNX+9REijjZy2BjjIzfM4
sn9ShqIKCdjRxvp2b5wmNDdN7uUW7QqQ/cIT13lEW1RU14MTuI87qlmP+GhviUfO
mwhcNDLVKZBAkJ3MpkriloWr5FsM0d6JZJtsPL8G7gDeEqhCigEUvfdOLftg9wDe
81lZFzg2WxjkGWNRoZHW7OjAGZnXWPFdzQfpIok9FruFVn52UDThCB+Ictxs7gV1
w546/UU9nKhBY0+OFgEVYFtyaYDI4XGkHgd/cwfTb8L65IWcI+CaB4w5qIrxs5EQ
80+GNUd1HUjMx5iKLorzVggmNXr7JooXLShsT8wPMfkzpxdQe882dxMStWL0vjPd
bd6SIU4Gt6fLt+ECGF2Z4TbZuao8XDzYIhV90Ch3TcrjDcbm/r9XcWwt7B4JVsGF
7CxtXWGnGrVzuxBkjk+3jlPH22GzNPiYIZYmVMiN/myc/+wWIqqrGQf8O1dYZT/g
3+u8+uaHFijRQ99WCM9QLALQW2ckKmAkSQikG27ybnWOCOeCKcv+jBilONKcmGdO
JK/givb2XydqBsknLmr/flX3X3TglWbnUKRBVvh/D9htJGYsybc0NdjHs/YvF/tx
vWGf79kCrI0M5LY4KYjKVMEXkH3abXe7Doh219/f2vKoCx1iNHuJQD8zXbXB6MEI
+IzsIvlRRRvZQnChVBtXcZ90xQPjB+Inbkw4L4amYhONqGsZTDgQ5bhHRs0b+KaW
BIPCbK5iLornncvpKZ1wkE5uWnbwNPXwvNc/7FF1oD3eKbUdy9dEQVNeIO35Gxgu
WDmRLWKL/2ickr3lmDgCC5z4w32zFwpzP7jQQ8Y1dIACswCWCeoTah1osamZW/UT
1zM0woWEhwWoyuIXVMB/pb+uSkNkrJ0igKqeRAFFxLWpD7451E6sWQjqugXYJU7z
k7x4vBjhNkZosb2EZ5DS0FWr/AgBLdk7c0+vfDGzz5MEI61I6mDt0CjCxvwc/5cQ
lyV8/T//HHnXu0Phpl0XeliuwQjUkIvPnC2+C7AnxOhCPAK8/9zohYA5VDCxcJyz
YQFrlGHeIsI+ymry6RAeTMyp00mlOY55wi+i7XTBZOWPD5zMtXhgpT732MtIijRh
WJ6XWRVGh827pUHUN2jGGqvDuvNwmo89wqg+7N8D5VRTD5bUa/NxRhHObVQ68xEz
SjKHJH+7NCvQMElIY8sL5FSY00ThdSHzWbTRRrNFP0nMIpYA3rwBsVJZdCousA7y
YXeMTrFdfRfOsuItBkAuejVeUXk7KKsB1T5XG7PatyBJWh59D+WO0ZG8YZ6sSFAG
PFYlVwo3a1z1TvjwueKRZa+oEEKglmlElccfBiAbWe+AzqZp1uIIhbOraFSAtG0q
epvHEoAP7s/Bi2xobB8dJ+Ly5ojRnKDc4MxRM+ooRYkTpCASbsA2R8jJezKynFyJ
FhXjEzCmeIUUpyNqLOpoQ7hmhqQgFPKwoX3giF+Bs9C1C6EMP2gbfFCrDOq1DWiO
n7Y/WrD8D8OxMyP1vunwbNZh/JOYVHJybXe1kSVFpexfTZlx1QELwAKOcg5z7cyX
Iz0yAjV/rEMVkaAWYmuY2jMG+6yD7kDhIMSKuC9JxulOuLVIYjdveBCFZ95eoduO
ZoJhafdozg/+DAO4jlYV9gIBxQ/YDIy1VNTTfvEnuknmrkPzeGv0BLx53PlpJRoe
fFk86koo38Lrz7+Hy08oBy2LydLw2jOqjno2P6BQozx7TxFFc3fSY9xhxf2Sjcge
RaCNCSjaKDe6I8anyguRi4aK/WfY65alG9kHVDYwv3+UwQJN0/HfJh0HFvXisoGL
JtFCfYvtYUvT6Q4FAw4Muuil/RJ788pfHEqkCw2HwA73zktPxo4R7WH2IZTcrLjU
2kVIEu+ltNRUTr3mWSylV4oXA6cCtgvMduo+32kdlHNTJh8zxosiPPZRuQDXHHqn
79tEwgGTQAsynmpBu6OxaC3Tut3HiGg5nsMJMCG/MOwrJB/F82eFxRmuxfXgtffR
D/lap46eSiOzWhWu+bDc+xdLv5yoYVJXoy4FvqgbtNTUD4Q1A7Zc3YM2YcurDxtY
X02mS5ZQg8Ri2H4Rm1MIpoYCPB5fPRsISUhOtp4u5YFDfeLUao5WurFZddIia0di
32bzq795QxnPPrciAy/GhBuxdrb/mRhR+swyl/3kTh+AsLPhRhR8Gk5UGj/ZpV09
U0RvSQQbk32KbXINP8KJRRMZzk0tqPPl2aDj9I5TkzRAr85XbThbU3fzPe3RnM5U
WC8OLCTZP+4L7SEIpjwal7SWRbDl/moGRPousQd97iqP2916zfmtgjnyi40DopdH
ByNNOiXW1KuTKLSINP3dpdo8WYrNYyz2KNCzVpwM6uLjANX539dzrplaDYypwnAA
SKVXbEC4PXX1fQ6hU5OYGgGe4Nv93EfoPD6YIDwIN75flFCOP0ljfsAqBJdyjdP0
Bhu+Gs5Bl/0ZRdPIqrUN50X6c8dbgVCFwH1mO6O9dVqqk26UUlYk2noz5vzXryB/
9otvLXttVuVvwHACndmvyNdrykev1ywIwM4bMugiak9DnLTPIHRqWkOb2O2CE3sl
5f1BkQSfIfbDR+JBO0SPK+gQUrqBjpi1HUK+yYiLIktdMxVPW1b7ap4NR/WCUtOY
gMMIGkhMS7bNFOYhhAJ9oeLNNgN4Qfe3AV2y0uK3YZRE2RHpmXrt/8lN/LQ7hVPG
R1dNUn9O3BtEJxitygmx3z1oi7QU+/D42Gkc/bnqalM1e+1G1n201AX9zKro4jUi
ELpteP5NFMJrPpT+dEwfqgG1cWcJvUbrIFt0AYPUe/I0PNEX06Vm4Z1o+P3vyoc5
WB+eCKSl27gNDYVIBBuiRMXa3ipOQJqw1+trYyUp4agUS/bHuhv+CL0xnKjyazQy
NVYdI/vHEDifOs/bL0SXsgyKry4TtvIyqMki4Yk0eIXqj4haHsuFn5NGVdP/lcMO
5k+tiv8gs6VpzXiO5cb4PsDmBmOSs03nUPhTDv9RX3+rOmJV4nd9I9hHy4WBu41p
mkCdLeLs9NZ1jSJA30xtQnu4b3o9oIuH8UUr5c3r826i0HzXFTT/i3qdFPNcdOEz
7DhGkXurjrKLlIp26w7bYDu5SDAfI8BmKj1emV7d0DlyB6BzNG2pPaFm7vN/jMSE
2o4Wg/n/fDbu+3BthfckA5KKA47bqapdGGKA6GIP1TGhdksmprqI3MPWGH7qSmCf
94PglMq3fNi6n+5e2LIGZUOnhoeIfMy4X4QGVFDhv5qW86PCkNzutr9aXZ4cTcf9
6UEIvkWoqPgEtdUH1D0/AAXpcDtwiTnDKjlqwfZ2L30EDuApvmve/EKuOWj63QJN
NTPdPTdbosgJOD1G9/gVlSdKYYW6SOqT3X3vVr90QWEOv42hGzCtTpdmz279Rmxg
SJA84OxkeKICpEhkz3xsYmEhzrU0LfLe90or1xbnygmHEPPB1qOnuFOPC6i3yBZr
ndIL/Tl1JhVfeLhiIIc5X73AdeNg16kzHAhSG1xt6gMwiEjULmPQg9l2CD2fhNVg
05XcKFdf1grCKaAeAtSPASWfWUUj2CjkeqNEQ1S6yCsEK/WgB/c3dU6XE/9RhM65
ix4FtW9i/8eaiE1p1Hwdttjun+wU/Cs2X2HTAf1lN/FRCbgeBVrM0486YYiH71WI
ZqMKm7nRZzubyzJzStWteg4C8y+fb/dpFnTfWsRImTUkqMRg+Y85RlX3uenMwe5d
PoVXsLJEn4G9JAoZfMsEzNeyLQOl/Vblis8gIjMEaCrXBpkDzwlP00DnqyOjeIsG
63r++UglqPgbdmuFKZ91ibSo5kYsrDRr6qldez3wTdck+SjezXolh/AsTlQVCFh/
QY86i6DTF3miFZPOBGWBwEsuOEjIy4gk8WfqlPAnRWqyzeC1DS/zbryT7EAYbz6I
qGMqi7gQgreR1S1KizgkIcwHQfTx7hCTT1KssbLSyJV4RG2hKqyrV14jhIm5MB2h
N5STJowK69qE2G3CSBaHnt4ngB/gAQ77AeJoVbfwIAuLW+zaaJcY5dmM/1uQ5J7s
lqJU1lacexake4jlO6dSuRUfkw04Bsn2Y7g5tvlP8zExDZ0dzfFjMxNLRRZ8tHUS
lW68ZVixb6Ps8XTG59Nh0+c94m30KjWlVOj0pXfPSIjcODRcHnQr04vVSSZhszM7
2uXIdOve4M/w11Z6RJ8XkrJQemGOCqdUPMHIr9G/HVSXJw5nDDvauHg4VP19n4AE
pIEhLVcYMNYRp++DriacxXVV7UQhmvHbKCesg3GmWACpg5N2fFsTkXzVbNPRDbSq
0eHV+OsKj55td+r0SzK5aJOWIT0o8X+IQssM4xlKlqssWnx5soe62EZXI9mNWKwK
vMRChcALft0kTu0cy7ao3HBykBy2uLMkOk86EQ71KqBMaL1aTx+JvCvHMeP4J0rm
kVjQPkYZuAlzo1g4TG/dJQdmhoIcchWX4l8sM/Cds59XPF+JcE2MMAr//rKLix4Q
wBLseXDRB1k9R1ZfwjO4K8aMP9JRq9kccCOUtrfSjoP/4ImFzLrFM1mI43b5sQFr
lTiGq0BiDQ98oLHu+ALiYNuf5iw0ZwoozL1kS0oi3hcB0QdFpCAVodGbMAL2GYso
KgUumopRI9nNMdG6hBj4SGHxEPom44Q971szO5rd02H52oHacLRuNC4G+G8PEbdW
M7gUwnBXiTRnchsIl9VjtJ1liyvA1ysOdg2RG5EIdsqbmQ+pZYdJf5QJW50GksYL
wPASRlKkZ+UnHuYNGWxwHliGRmTKqYZvplKd7NG0RnG4dscA+0dZht51jXxZQuBB
4msgbXPLq815MYtfVXF1/UaTqL6/iWCfvSHTo1uhxESY6ufz8OioTNvgMYAl9PMz
QjzxKRDK9ad7koTF/fvBMTwe6ibwljVZ9WakUrZHuVDHNTieTskezHUK9R6Idjov
W0HGTGU2v3xtaUpxmA/kY053qhoWzaRNLuHmQ8QE7g/BcV28Gb6pxwknMZjCRJ1g
mfnn1YLHWPAGhJ1sORx4NVppAlBPWp3YIieKnnmHkHUgZHugRlfi5/fmQ9ALTAFT
hwQwjJsLzP/lj0AEsRi5NrEfTny/2HvJ4Emets20BzgB8ZDZa96seYUwqouHmxqX
3DXIqnebgaiQakTaMnVKqlXyrTGsBAaWhRtu/819p512CgVFQCDMlwoqTaKJTTi0
rFbN9HtSH1EQKrsrJqMvwYBTuScoh4p9PNCUVPN5cFTMW/0ds1GYRMnOCHvYBx8D
bCivLe9s8fvsf8zWUGWnNNrbFGVRPhQ8TxAsJ5CPrvq3jmZ7mx6kWMuVVlfkpqql
VM7gDBrO41uYYbExswNRh+BRyDbQRgkNGMYaRpnLdAZYyAEd66X0MJYN+KoPwoQo
e01lSnY8WgN1Jb8YA+7R6jM7rdL2+N+b3sejc0gKPpsMgEyGXoTq7cQpgpAEcf6Q
5Q2TpXa7gMHi2ea9iEyNP+x9KmnvOHUxlNknnHioDQDdVLgISw3EPaNCps9tpPG6
Y7Uyb30DvHgDCQFMxcCqrAjpau6WDOrqhUHXQg/DtuaGpi4Asd7Oj3xTmZYCibob
nJRipCfzcRqYSElQBtP9d5z6VC+JD1ntlPk9Dcpwfzurptoj0EHgJaVgJidmpN7F
nAREySAZqbwPwCiObF3lm6z87cHpJvhcaDdJqHw8L0xH5We75JYKjPb9oXO469fi
1NztDcaTX123aoNQmiacDTenLJIyPNLOBo+ABmHj2I0aWAF4lFFhlYAPjVYC2djC
T/3h4eGQa6DPcJinSnjvNge1IkG1e0JL41o65FgoyjZ/NfIh7N4sKpjk9r1BuV+Q
AXJ50wFQL9opEu7q0d+7HDwTcSDIhyCWsytwoc5+5fqtaLQR9hx75hE9Lu+uz0O6
xUzgF6rX0T4r95Zn87dqj5F0CH98dNuUMOzn3Cq/+FzmxZG9EvgvoaLBYBSYDzen
MoCYIjqjhR+1gOlNY0w7JwYCUGH/aC9itVlQgPlPfL+Q0YFgQ438uM/TOpK3ciqW
8XhhgYjfMgfsTESBS3g/Ng8BNuqBPO3OSDbF2TeQT6QEA6jAtIGt9feEVwyJSEQ2
wSt7RMzB0Rz+kSpVM02LlHZPu7kakIWLoejelgJNhOerGAW2lG7CzzWC47CX5PWU
I1HgAj8uXyYammdqLJAIOj4FtiIpS4PzkmpCJusww4oskl6+cqf4Trdbh+qzQ2nS
EW+r9sfvCiuMR9VIMrxRRMOjl99XV5lN1XbcdpnIBkhG0wRRgULJrMBrTCKwZcMT
0CjSSJ1icB85b5VNu9mHYD5Mxy4FswSOo1iJda7GQN2Vbqg8TtIolWJvMiA6y4b1
/JFHKBbxmDP8Zq6VTIJXD+QOB8Oq2jSyEmGPy3NJpu163tNHJlUmLTBM3YXVz790
SoFXr48SydeBOU0aqPEii+oXS3JxUAISGmRxSlyUS8KbjkJGCQCumZRaRsI3IEuh
2tgVSr8SuxSgzx2hUvwIivybJZ71bJO8jr6dJOG5GCewa0d1hfxyRROlYgh/957N
goJbXbB9yv3PtFg8/0ol7neNPQf/TwZlBXUtW4vWwyQ/3YOuUtYbVUDPO1RQ5b4s
0ehy6hNRRAbWVeYDg5iElqcIHwHL1xWTtcO+By8Y9jV2ugAe2CoYK/GrhyzHcjnY
NQi13gtmFmxJW79sLhCqFrYj4Qr50NLBt1dte7cW5zJ0Q/3Jey/FqUCDOsQz9MT3
NVbp6LoA4i0YKn7pfKF6tel/TnHsxIseyCN67ykLkb23gy/MGeZxYxhfFPktzkPA
Lpm10EW6Y1EkKwrB3vkx1TMBYdOP7h6J4xXgDjvs/kLHzZ7104nG1iBxH+5ARWxl
G5qYFlfYC1FK+seKxxQv6OMWf5u+epIGpiMBgJe1Ffl/i96Gdk8hxq8O2z8bvAb9
cmqJu8e9XsUYrfjM35eXd/tBklL/n9R/DLXxvhENNsaZB1uqadEC3CB6fJbVj2lV
a2tOTMxSNigsQ59adgeDcBtIIaOTEW4IOY5AlQND4Ye7WOhDnhribZH+h+z9X//l
fm04XiGr9CRTZwJp2DRLuFpdc3Q2E/HiOkuxyI43xu7w6SrNpKnbQcpKF6cidaur
JdZrcpB9t0yy5V0e55xlSuCDCPP6i4dvPmbTcUWbuVZg7N6p2X4l+vDkszZ2wpb7
1VKVZnAMUPtwWZTyzJ+2udDH0iFHnfu4ZmqVbtwqRmxFBERa6czKTDLqIBw0078h
cv8Kny/FPyhZDZBGmYkPDKY/55ABnGTM17J5eBrZ42B3I3Iqb95hy6OPdBk+2UOm
Jstk8YJ4TNJlAXZshh5XL3npYtVvfgnBHcNzERS+pmmGVYFITWqJsPKiP4sxwWCn
tGT+upV4G9zBgz+763d9MfX1XdaIIWE0uDbryqINPBCCH8GmznwUYyiXK88Ry13G
Ov8Y2EoukH8EoLCE1wqu2EZ+WNij5FKecmIKRSO8NrGK3xHgnhRwJ7BEwQIIBe4J
BYzizcbWjqenJI3g5aowdtebqAEI2avye95daVeS7ES9Q8sAuz/yUf+DmNCvHOZ6
nk9qkoo1Vf0jxTiS27xH6GKyB4UQGlgKgFjE4QmrEnQ5ht7i7kq9oqVNurYXESg+
S5UJYdQ5e7oXl+KP7suK0VxIZlntxPkMOqKKWuKoRGP3JtMpEnrwOefwyfSWYpy2
XsD4MPnMh3+MFKrnXa3Q4B62cYFLGOtuVmxkQIhUcwrSh09+f7O8VBRJBqg1o0GS
RhnQwTKMSsWjXwT35plkuNfiyeuHCMidFn9i/b0H5p7woBGVghM1WNJ5g1U2OIQ7
0zQwhzyQ8d7VMKfFmhU5b+1RaO4in9RPPhwT9g2MmA2YJqfByfwS70NxITgjH84G
cnPwTATegCRy2BEpTtJyTVZnqnd04nkDgs53G1AuzpCn2ATZJzniy+x9+f4YQL+9
bc6TuIkNdnuFyqc/RDgHd5iGyQoOAU/gJ6zt2JR4HBRd/7zkMGL0gkCX8fzxG6uN
OBgDL4fL3dC7T2pVFbXLtqyRfu/FDTO+BD6DQ/iKzyYCtaKCgzje+tBwHXe2C7AD
H9DSESqNkQvUupplsuEXAzxABJ+QT/oHCBn4A4jTVL4TuSwiYt1+LOLBAbwfczeD
YUJJTcjgKWbwYikNr1+7LDmXcDr2U3RV4iotDz80T5LTxFV9MOSsi2E9WguMPKWt
e4q2h5zTJgceix1DQXtdDRpb+3tyvzqrXQG/O6HEF+FeXKSTDOe7KSAV31UPHUCo
pPTsYBjesLEDJuveRYvGVjaTOP6LK9bO299JtAhaJfKfDIATOuLylCNKbdznr8p+
pzexK3Cm/b6xZ+Vvt1g8RSx+mGzBjd3RZoE439cz9vS9HYAY/7nkPFZrwtbmELSz
nWc29Z+4XQG9yceX8qrp1NJWcXZ7Cs6zUQpV9SkCojrjlBagA13zLI3eohNlUxH2
gfAOdvmJAtOO+w16kNSOu0QMbQEtQ4ENGmxH1z3eV5VuoEIsgdClYfWZyCAZfwNz
H1A+0xNQQVoIEXUzI+OByjULaEEeCIYe/TDUj2VDNOBLnDAJ+TGCa/K2l9kp86Qs
rkqTYuR4uitVA88723WbdAIDb4cKUhZgKRrAtkfpBF2/kcStyqkXDKU4uDlD/4Wt
q8YoEYh0IdW2Uoh22lSVpg3BytEbzUa2n8cpPKjQ6h4L3pVLa+uZQjpfzA84Jp/u
wN0VFykS9STr8dnViZsBP13NxwQ1B1fyiqS+4+ffWj88w9Xlg+cAwhQepTk5Qs01
hatRNcI/FlZUhybFF6HR/dNGm9aApnKkk3fLa24zyKthenmsEyV43TVyd8qJcvmF
KjNr94tZyZHvdB966C0utRYylW2hQNzMQ1oJ4B1VPn/82zyNi8x8q6TOeVZr2+I4
HvfmDRMLpJjrpi2cr2ZjYk/N6XSYEV2B4WPXWRBkYT1Bo/sFUmVXzJK90l9QMI7R
TFdktp61fIBGYxdrVRIw5BRUf8rHEodv6Yjf+P6/CtevJHxNoV3fvwvBOTgbq3/I
UbxavNgrsErQsTT1vH4Cfa6BLGO/7PgSs6LWR8AtHpE+/ZivvLbzNyEtgsxDU32Q
Ev6cpLkXvfgo/C/wSPFDHVGIr2h4ApFQLXUKp87r8FBEazq3bzaUvUMr5hYNVwBI
Ox5MmysQ5c5g3tm7AUQ2Rr2l0UO6ZVoQ+YSnY3JKYLGd7TqV7ZAGhLSnx0riIb9Z
YvslSHRrjdeBm1kngBRftZrTZMFFVq1jsT6SJfDz8hkEB4EErUwM9kiJaugk5oD6
ZIOIlHIYOMhw1mxWL8FXCrt+8ecjZat7z2doVoGzeAGVTw7pSln80DHhLKrtZhk4
VWtuI3ievrVKHGJUT0SFBHkkWYN6AyRk4n+/Fs6bXtH6nP/uJK6D4uC/C8eGFAf8
UVESYlSjLOspiBzIq/DmT6UGVCEM+0qNfkwYI3cHhNGgwoPs23QtSmGICpfT4n7M
BgXi5JY8+jYGas25FgAQUtFtBG0stjtbBozVSGMJQolu4GA+oEzKt5Wc1vSRUmC9
Boq0l266Zn8KuwX/r1PxCXGIz0rzFgpUPQTBrK9b0eYLkw0lu1m0hP7ZfK8pA8Mf
QgTlWiOc91pfH5LCp/nbRvmsZJUJt5EqQgJcT98Cepg0P1S6fDR+bZB0xC2+FusI
L2Stv8BNa89BHa2jHz0D9ElkRvuV/cv6mu8GOqIpG/hewJWfLS1aKqop3iacvLas
GVi/t5PQTyoZKGbGwncyECCEBg8Hh01CJ0esdyMGc5w0jMk6wM4GzqlNp95sK2en
OISxDOoG+N3RgPisK2VuvL/2Y0/NhH9EGS+kqNnapzVkWavugAE/hllbFdG+uyb+
24HDuag/4EuDrXsYLTq36kWAxZZuvTNo19+uYw78bJWh7Lh1Tk/4oIHW/Zbh0m1k
7ap1IbvQdcF4hnNnjufKFY97DZwgP+30e0NT5Vin3BC2e5ou7STQh5IYLv3TaVRP
vSlJ7GCvsl6OxmSuzBopP/JUgQsxeYH4dvZ372yDiF1ODrG4cfyLqkaVgHus+rgA
g5m98A3z0Y90Uuya7z0sjQtbXO1SRMCau3fEkkShPCsp9N30gQZoqXBo9zBjmnvZ
KSRVWSqzCUYOGmT4m4rw13exo/cHkJ/wcZhA1XVeAleORPSu2OHRtzuYyNQ4eSzY
hjGvHjuZS12jA1e5HRE2lysYwvi5S0u/ud0BaMpo0vQSN2fE4OG711bRlsowsnWX
CV/G3VgbyEiUwmbo54Er+BSWmHaQxiB/r1icg7KCJUPET7UHIfVML1owqe5G9JBL
I8+jshIRK7NhEFJcm0Czxh3LY26zhGIOvlDzNITdQEXkZX3FfYjKLbFpz2r47E1P
foX+yrwQfPOFE9ilQK37pa3jnv7LpE/QHPdwEZiqSVfwkpjtA5BXanIYGffuvcN7
XuSaLIwEfiM3cJFOlndjdvR9Zft/31A4dDOh1CWyJpTJm8FdGEWvo9scWM1SR6Zk
VKSRJ7cUD7pmQkw37RShnWyIjdZXviO9Gi+NcS1Nub/p6/Zo9ELz5mz3UWB+tr6h
iXqeVEgdf9BFH4Qv9xogl+23vpo/KIpTY5qFWpgFPVzJVBTECs8KVU/ieXrYPXfa
IgVmRZFD/XJvgboRQoVCRVxMx4tB1BWSDfCI3X+WoZw2J6GAEmaZa0KRwrNOGxWY
8Oer2z2cvhd5ib1Gh+gFwfTLqoXn4338sHSYHAWImOsLrRnGnHy+P/PbrFimYmGI
B2ZTjvo5LgjXUWmHa5dj6vF+xmwdWNyNivSnm/FlH6GMJAfadxspVRciUgq9QB9b
83YQquRDtywV5pDptV5zR8lnDXgNE982IhDwgwerTaDzirBPd3NXpgGk6XJTrThQ
dvvAFJjgNPZtv8MfkDnqGrY3RXBySj+ln2zURGcS1gbKDzQZlpk2t/V6YykYvKZ7
w0CjY58nFyCRpLA983n2Yv1DI+lHuZncH8AKvhIxOErijRM+f1BTB20OpOwINz9C
qu/aUMGTGAkiNlgz88d7vV1z3DFMDfrVLuJw+dL38RR609lte1CF6wZR/Yg5SUCt
iFNEAHuegd4jjqheTaj7agxtogKP2Ny0I9EDx5AaeRjjFPYN14Zg/QaiYGQa5HgV
d5OSAoCFb2c7MNX2xH76sXjK+1AM86/TE5GQROnazGU3J024RwtSGs5dfdrjS6EP
Lk8qeWwsk56BJ2r7Mxl/k0x0EDOA26bL1UmLlsrBD+4PE6QPcjDCCEpgu9Y4bNi3
auI86m23l7kQf18Ojev524FLrKYBGD67NPxKTcS3X1zSo9jWfoweJ64VxT+RrHmt
z3Mthg6O7DhChpWzPmvN2V+4uS8torr/kzl5vx5QdB6lUCiSAp6X2R3eZSJ1P2Xa
XpBTI3GtkGM1g5pG1q/u2Xi9OlJr4K0V1mY/Z/pqipIL2xJCMbcsQPuY5I/5vNvu
35gbunyt7dsmkmZAcigITfc1dzFmOf5ieZm6scTRD91htdc7aILzqdHZNf6yfmdv
b3iCw1gec1MecgHonXK0KjV6snycqcp7asJfG25MwGMmdOtYTsf1YT4fGbD+NTpW
tf/JHBJtvzHeUkWgV/bYMfdYHg53v4QliOy6vtoD8a+HDvZuY6t2CEbCRgHZKoRq
LOWLHk8AtDN30XYic5rTCLcJkq+6NEjmJMnTETqMMmIazcEsYe882n6ynQTt27Uh
zmc3JEL16Nu8Nh6li1+s3CRIUGyQ/oOgi5JvusQ5fLOmj55cWjdmNAzJpbOBbx4e
EfVJ7eKCU28AyxukjyAGWoc/eaeQhXN4Ye+HPpjnbL6kB7cRN5zUvVfScrv63Nny
Hzp9egESdBmjcNaJ1lvmZ3rwOfA4tmUaVcEQwSZi0OZhbAIiV/xYzKzt0LgL5QK+
DyvhDF2FUUEh3ay6SXy3in/O5kasMP3boZnklR/bSuoaOFmljXpfah7VqyiiZ6JY
UxypZBJBbxLe2/jGg+aTpwGg0B6opEHDdzcYlixweJ2pDUErm2bJBRRBoVbTvYQf
JL1tQbmxqYcEuwSu7RibZYxmVk+XudE9Y9Yc7z9rNf2Z//q93/aSBXHYJjDOsl5a
CJI9kvO595EePUbjBeKTiR1sN6v5SAT7MT3f4Gg//iMcOFWBWK+wdPqmER3TaXon
oAPOMyeo55Yz7dc379It4vBsffeG9hsquDEJqWWIND4oMuxBuXkgvie+UUjznR+K
PDNgRZR+b2D6Tv1rXqinbXbhulryem9P0k6l7l6RWVxw0j9lBi78tofyeICXzEhf
WQdWqnst43Xv0SamDCN0JLlR0tufw1BdXixvSPAx1SgqSF78yGYBb0xBltwCLTrY
I+ll4tqi5ay7mk/idqmm8JXp0si5x2OkPBYa/DOjbSC6hghJrAepWtgm55oD0xTO
jeX/8kdqD5LPCmzp50CxdRJWGo6r/Q01yRoOeXlaYSMUd+wsGxAkBX0wJqmml99g
n8+qyimcTVwgTqBokJFMUZS9JkJE466mPBd9616R+HIVnsg4g662T+PZ18P8EC++
prBpYjypNdfDeCJXUao/mmsjuTVFxY77nMllcYsbqtk6cNZxLKQpRkZgVhvoZqHn
7KmizECVzS/PDYaPVzhECTzRA1FAuScjyn86JTUWSuoM83mvRPhJX+IGhXrIR+Ad
NQkSstu1w6gfAJQdWXV9stRjAxy8aZ+5BeLDTJC1MxCc/keyOCox4k7znSjhGm0w
qQk0y+4kh2XkYkABn1zO9CA05DJWvXzJcYQob2GkAupEC6zu84F3DDMNPcc/Rj7E
erqoqI1oFmFkUzJC0qODDUOIIsxSPlUMsEq9b/R02xxwHTxNUbo46EKRx++SWlgG
BZip3A2QgeHAnfzynZ3uKlK3zm6KVFLfgHoFUtiB54JKtw2D18hxMAzIabwHvmLO
WM94J0GuC61rHeBQG/7VS8FCnPin6NYGoiXKT4jsGwAPAZ2INZ+ODXz77WW0UniM
mNNacLrKnq0ejWUIz5j5ZiJsSr7RijjI+E/zmoGXrI/iNmdpXtqKoD7eORxDMYoz
EcF45S5c7cJdkhFl0HVHf6iP9vyrSy6CTWZwNMEMfjaTf0B+fQfHoVzh+Fc8Uw/2
k9NsXN2s3MN2lUPMVLDodY++f3/mpYpUXnaBle7tXU/xFDkMybEDTLbw05KPTl4h
Zzti9HzXKWzEEXncPWscZFh9u1YqnSiw4s6SlNcMsrF5vDwD/AMCKYRRLweg21Gh
XczU2knUOL5Grr+wuD8J2/Id0bbga2M7py91SOEiy852IfYhL7bt8MrJT8FkswtI
8R0i4nhFPLy0KDFRbtnmHpylsJSxaDdXgSO9Mp5T+mehI876lWpfcbeQzR+oUNNu
64DiG2UVmO9YDk4EusJLl+GtwKep7OFcEs3op9Sv6++x3GmX2dfp0HeJcyTPuBNQ
uZ9bDdMPGV+QizDU4Zdz7CpA4Nf03ywsWUPc2sRuyylltT/UlZ3bvYf4tOQ7TCvF
uw/I+xnt8p9Z+/9MkkIz2zmYcKRbrU0qX5Zyn9ZZGmIVysvbClg4qsE04l4/QX/e
jAGHe1VDs1gey7r1KIwf7TupL5f0+A7PS/O7D0eVU0kF0MarJNbBj2E8vzHb9tzW
a7nbSEbAzB4O8Y06yPl3k5eFeSX9ca2LftMkhbME8wB2pz37/WnIgVRZLOa+efkF
Md81XQmr1u342eghcil404AYgbKhcW6OfW228FqhiLW0p3YMGkJnn32u2atJLgN5
Fi545sPN1GHDesUk31aqQCSq1lMaQwZpLLSbqj5X1xOgaSUqDu17+lh8I6YnbaYA
Givg7gkj5JG1RKoQtVjr+BGV391ZUg1vZAEq65O8/d22+LhYQPmkSEzsZIjj5PKL
eB1QqS958wHtRwRSwTH8A+De9Tsq2c/EqVK7a7bd8/o97j6c+kWaq5QjOk7mWFZY
dvRxmoUmQmCGOxmsqMPtuFtHlYYyUKLt80fh5IiEKzz6IrcW5VghYzL8iYrmilwy
alAzE2FpiXqQsonVzlDEao7vtn52yJ4blHrFHyDvSU6c6RszdS48HOfOeLE6njsM
QoKY9dtVh68RLqnlq27R7Cg2rUyLSg5jM7y99tyfJAAIpM43dOhHGlp4jrgWP6/i
udJ4jwv0Ekr7KcN19qIuuWKgZ8FTD3sn5t+tQUbT10tWYUal2RWyj71eNZN5iymP
xYMZTqOyKNV6zwULOdbw4EU9XQVN6zgQdCWL448liBH0BrHd8DQVMHN3v03joqJx
e5vTIGL74uQ66P6UjQmhy3CdPBaeXJuHlElGODsliCXKDYB79L/2vwI9lP2tWlAV
k4ftSxz6dGSEy0EW2l5nGEx8PtWfDDZfO2U9h2elY+xxa9Hln4jrbnhEqyym/94S
4r77KJu83YsK/i/4RkQEhAWJGUpxsN+i2QgFbOVzhtNoRYX36fO0eNqq3I5hizMH
CGsNHRxLI0FMUMH1v1BS6KgnbZJK4iSDqpiIcuuLHvP0DbbZ6PJ6bcuh+MQ9d2VN
KRmuwB69LSMPDb+GeVwE9NXu7Ui/adoC6FjcW7uffGEdo2Pw6zKX3LOrQ456oK/9
HVm3ZyxVv49abKlPgcMqhEkitpB71MpJj4CGWmyecgE3ObcsRmdnXYkXJV6KrhRE
GbpFO+Rz5pPFGwZOfhGUAfDgIge/mjnW6HMlsi9UxPB4vZd1/k2JKi1ZF5bQgWLJ
qnnfA7PDiifT2vtbP1Z1+CUO3baC1q+nyV7t6Ha5Qj3uBY0iR8PLOH9bxF2Vn6cE
MtxWQT4+atKSTPx9jh+8K8Tz8xeoHIwm6crd+Rv0nXnFK4VzWkr411zXYJMH5g+n
o+iJ6myiQiZYAj8WXahFfAIGmEWfhd25bDIugRxilvyyK2eLROhtJkuVLSow0r5+
PWK6V+oUKJpyPDtbBZPaQ9+EN/3yXCoV+Za61DKStF2DPDmhX/o5258mrsPy6OVc
sFzIBkDfHD4V3f/Uu4++XeyvAYar7CJkjJyLsxhHelu0cnCXU8e0G1+xDFKEAp9n
Cd/4IT4XAMxZKDtyiFdCITdGe9X7iMOn8uwYPFPGP7H6Dzib9r8t/+sik/Hg/oyk
XQemmNBzBUV0FbVqMjvKWtVoYPrrxRyWfgZzvH1texd4jHtQ12gG50kyBYVzMtDr
xrDNT92WqliIN6kgmguW78Na++Kjgfltq0Muo9KAIu406eYtbeAlmi32iuT86b1o
vFgVqXDX6TrCqu8bV9IGy/vxUkUTpDVc3SZrpjTcmk6q3L3PWvKzaDlwqxS09Aq5
KsJH9PH7B/flLaYWxIgXREhp8J+sk+zzWPpsxBiOj4ycxrYY8G21bKbkglYyoCKh
gN9O0vI7etqiaD0BP51nHHtZnppSRgh9XOgAkgYPuGVmO8J4xTTGaYHUMJig0gDb
/FUNMzJLaV4K5L4dRy3RwPybw866jm0mBUAq056dPn+RYFbFvtmFVmcw1Eir/PrK
Yc+QSwPkJIYGDAkqASoBcDto381VW1a6Mb5O4XAc0qFDfDzh/7fjhGaR/AEX2Nlb
6Lg74l8nGR6OJkhpdxe+9GxFvGK+8cctStpCNI3CBHTEojsy6xu/aNlseQGe2RTb
fwUjJe/jWGWyhaJrMD2aMC6Ftob92mEThaU7vDPY0StH9nct0xtTvBWwbI2ZpnaZ
1P+wfTNsvXUZtC6YNARR95dfAPK57A3kuH0mcvnVcSnLfq9ZsDlepfczqv53XoV6
yV6YozD4j+vjZOsKhy8QaLrQiP2/s5ko8pVGSVYftO+kMr/teWD3wPuUF++Rlykl
w2NCwN57oZ4UWLleoeq+BTQ53cjomXRnygYuHJwj4AA2qRQi8rMHygKj2bLvPABJ
TlWv43G25PC8tCRZbeadYQsYENZrcfWqFME4m2cm21rojbHwiciq5u4zYI+VEsBA
fc/ayMdZuv/EySE/YIwi4mqja95oz7TpPEzTRQjlMtmfcEPL+izLJEVbbS+pEVBq
qbDsaCm4yDju0HOOhZoZYQNsGl9r4SfcYqzeSBvrTeSm3Q85Vnux4CpM4pCOyVXn
9aKKgibmwk+9hr+nMW+SHmIH7bJkvt2PACO8e0u5uhG+o+wcqB/8G2pE3eduFmqm
o9egxTCbrueqpeDiY7StegGa3p3E6BMHQNW8HWPjw+lQc9qedI2RPJD+RrAGW2D0
jVcG/uYUgbKBxMvImA/j1onwajQEefgDr6e28QYUawvXl8VNQut/6M0cbdNgpDZe
7IpMmfzIeh+GuIqJQ+IRLLWnjOt2nNnQom9s4kuf9lsjSjrKS7U2vZa8NP+ZWSQV
IXrFLo63ut10L7yqBlrT+bS7gX0HO0U5V3zc/b5MJG2iP079uIf3bcBI5eFpV+f1
/f/3aN1SskxgEUgYwRKmAyaDycNYM8aMUnH+eGpWEA/b0vuMYeXpZr0ti/nPHqHf
Ivdr8w52P/RsEjeAHwuP20j0du6eRaQN6IcGwk1xXKm7FhlpnbYmuaK/ScbpZ5VC
ST8c8aBCmZvoX61+Y6oXhSHgdxhLfT1NFAfCV4Ph/q2TQxjtje3xgPl13vqRWOMH
/YIZghHzkeqwVOA/xE4Kre1S4V6MYotnUT8+guunOfJKyo695XqnOKHaASTsT2s8
4tYY6SXMyGC4uDRTp6k/eStDgBpSnKGIVIB0XHsht2JlgyjPHaEaXm/GINPBymNa
4OuPD8MoB4jwGd03EE4knbNZ2pVjEsUwVkyBB/lUV+iQf3Rxhk9dqjfmt8y1hkxK
Oh/QKazPEoG7TBRiapfkgRFPoT6qg/hZE2ImcgCSCThVlmeriUAKmYP+K6e6eRub
KLfc1VQXUiycd6cWBdVfrcyyq0/YGMWA20IksPKZOkhsZadefKmUragF+Y8BG41R
cKEFSKet3mV1mLV45BWmfbZT01mrT8ztfwfX6yoJOyARYRwcWsNJuXeR4rxwhW1z
QDW+LpccjIZdLGbxcWkLLCvGuTZY68In69AsU6tbObygo7YuHw6vTk6fEiHDzFHg
sUTuE8NUPpfzTbNHR3gdzOpqwh02uGzwk3Cmd55XgsI4RVqngvYB+HtJE9Tzp01d
cMZMHG73sIMmOemOp/hCe/8E/D82UTwjfblzL82jqL2q5QcxKxrc7f8H3XiEwzOE
81DV8Hru0O9aaS8VLFEGRWnu13hH1lsMFrhayYt9qcY2oA/x5d5XgAFheolpWJTW
rm1YWPpDzyIBQQ5COBHT+iPPRpQSQ1HxgrrXF0bsAnoNQvNeyelWw6hFRiHPdba0
95/ChbewfGJniFTZ8GOh7L7JjgTHEVl5kAmEu4K+eSiMAdFEaM3nivHYJum71s8K
rrieZygBPgKM5qo9TvHgNKKfsqTQeztXEVWMyTjfILAdVNlI9FBXbaFkfAbbYNEN
QAEHAfv1Ue1Zw4LMHL+7FLKzCXOdiUWEeVnJ2m3J/4VjnItUE5r9Dv8wPBD/3g10
YBU7tA7zzmQz7j+d1c343/W2ZVS9YwundZMQNzS+UOzrsyjaBESMea/26WBuX7sR
e2eIWpO1GbfsJ2LZOYGkWjomlzBcBIBCOpEtxDnAV2CymGEfuHx/UueceVfeo+di
GF4K1hoYqE1Uio/CVTSBs/2RTewzEeT3jHLXUzsOxXd1ypp80VA18t51QqK/n+4p
iSf4pEpuRUz5MQ53wkI1KSmIoMY08/9pr1yg5qUO5+sQ3mYSwgfNhaa0IFlxgJNE
2lNp1ZyBj1LbywIiWH6RolX0i4Ewf8CQlbUVgieCa2d6QYlIoM/tmVjmFRgHdf3n
PcHEmiWtpvWKZ50OA5a2TvDHCvszcoQrkMQEJXX0kW3Y4ThaAZIcpdzTdpmYiwbm
vrYtKElzUZ14KopRFOIpZoGzcLrAjY9FFLk1jiIKeul3jlQ/BB1QhX77cfBGB06y
qdaPQfEJpXjypBvp+h806bjmw9ILHTUI7XbwatyAXtobSnCCreZ5XqFl5BTWtqIf
GHU73XKURH04XZ/xXkrqe2JNjDeZS5x4VZi2g6yl2do9Ql2+/BHjFdBnUGHZ39oU
3a4Hv5wTgtjEZtG/B2fFIt8eW33t6fP+gF9L/PHmRKo37qQLOSlWIA5nNKhEUYWY
eJsRIvoK7frTY+vdKUKzfcEsLkuxDgmlA+TRVVUWA3zDPL3BDU5Uh+tISYo/HLCe
F5xzYeVTkKkbeu2jOFJKK+ZOdS1WZh+ghVjIZfFOflAlPj4LE65tP/U342KGuCRa
3WJJMoiuWRFULtlmqfl4ucYgWSfgGFmdt2rgiDb/RGgpXQdkPUOZcNbSdiEVoyyg
weSIKH+iZayOkN3sQEMdOu53OnO/cLeraUJoqeJJO/9YOsfsJzFDKdLOH2SNMa/d
mgWYjnw/ihjNrP2JUH0+BdvAHeLqXK3xkff9+QcpOL3M0bBwnL5tEK0k2oQxkxrp
OtlVh980tb2yWZgrpXZcgqzg6rv24LenFidDjBfxWF4r5nVKNgh7RfM5yhYJ5t5A
FbdM9dX44RpvPoZL/ImXHz+BOYzKFoYbm1aLh0ZoP8JTyGNLTWEFRpXKE6cwdMif
8VwZ22ALtR/CahdMHGWhyfE4qkwxnvN6X8ibfCOIBLQey+fbUC0WiQyP3GbLz52a
Q0g2wEsY+IoZth5DrDm9pCpPy1yGLAiv950k2R9P8wVjL9Cm620QSkEh4kmMwT43
6CSFIkibqfGxIZnBWvd5eUsmZfnIYHWXkXiX4rZYhKvSsO957q3KglSM393X5Brk
mCJ13H+g1/wW/VgZxYxEvoa6RA+4fbCSGfGQ2SknriztWvMC7Q9AHonvc7Rc5v+H
HoOJ70/0zylJ4a3PMRMVn6ohHDtFZmTVxpqSa+uXUb7oQGtAAc2Rq3JccP/e98HP
u3u/84Rd/WVvCqocB0G/8089/LRYe4eZ+jNqgIxGwVZeyjQaNPcsGoJAEfXCW0pl
ve/FwLeJgoYbUcYJJBdu0K2TMWB2gas1VOFjg6+mGj3O09WN/pP/t81ofLil1Co+
1HYs06+7bTx+oI71SePjG/ZdkkUC+R7U5Qn6EohLpmJl1yNpwlMvVS3gwTlfB4PI
l/IQvXmwS5pIyiD/fhpZ8/nQXBQprUdNo29HWb4qTqSdPJRR3/5n7hJRs1+6cTkz
6xvE+uFpbpYBslW3fdErdQJG6c/kDwcr4qGhEo/zfkDw8TGBW/xyRUBP/gtmjZya
ET+yFwrE0V4elc9pdeRO9AR26buDKhI1vUm1dKdm20zZIHa8fPI9DWlwq2FWrz5a
B0hRH9mVzQMAvpchdXfgw3n5YqySDPrNW5PS87GT8LD0K9whyJWxbGDcY9FNsuRU
ATO17Lj4KcTtSdAaU3HeuMlAJzMHevGnQ20ETtKFPDIX9F7nYNE0tIC+o4LMXerg
0LaQFTQSmZbVNiidWwmuwlnpPBc3SaVSnCjPDt8KPefR8RNFffAaxdPGsX5l3AQm
Z4j0YGAdB8qSyBm9TS88ps+Vre14/0MkIIfTeI/1n24u7ghaEbzF3wV/l1AzfKmO
0LX3780WqZhZjSBwGHgyKf6JF90IQegy69x3oPf3Pe7NcdqxPjkJPeKx8wgXIW2V
WTAWPIC7+K0fF/SOwbikjrRDCuVZFfIQPPWj1wSYYnsGVTLqanyFizAxiVTEk/3h
Y7LupIB15MfNPvTdH1sqPi0GSwoisRPxnEiuPN2gSzZFcNMbIETmRCEuF8PJ5tPN
wR76oY0awQJCdSyO+aR5lB4tfJQBeSLFAA9iDGrAXCUW9Gec+QRZYj8Yy/qj3tlA
FpFDCBey1LZZwD3lcEZ49RPI7pfou4sCcZE1S8O8XLHSLauSPYEZBqL2FdmMGgZm
t5s7ataRZd8U2ypd7ea7oNMMLIkJ8SA4n1hGx/BD6laWEHVMabTVYHcjn2qzSUSo
RdpTzM0XMPMbHb6iQTm7W9t0LgsC/gHdCUJ0zU8v4IlGdOtheYIrpVf97HkNfuad
5xbQP47PBC98H6Jo+SshZLYr4D/7uIqCx1myQ0mT4TqPlFDcXbJS/f52EiaG+Eqz
U9dUarCdJMyuceUFdrPMj5EyLmCWO0MuVYmALQziEg771bk3B7/IQlQQTmijDVVE
LVcpyiYekKZTsgstz/FkgfGeWjJC+hsi+6v8bThxUZOyVZI6buIsobd6lOrvZiok
vg/sNnHCzGzpEn7Z2k1/VhIS/aCHgOzP4hHhKjJi5Y+QCaLiEoEBSR800HXpzsyD
cx/hyYqupQYvRZlISLvXiDsdoE4RrCfxniv29kXPUKalBybgwwGyASohNyUDqRFd
OUmx+qDwS+znTmoVm2yESLkYiPMa5J2+pswU3x5PQDe6TR2NzXaNsErkNvC1sAtz
S+AevfApVcrX7MOn15aVZOv88OgYcPfXfHoDP1fsjrXD5mHh1scpOUTc9txZ+lMW
XzA2atU9QFpLqIOlVCg2LmZTsvYyxPR481sU3g7C7hOGfVnPso3IvYjEBSbC2OC7
YrLUPPy8IOMzpYSE9dAyw1UQpeEOHihIOyW0SSUuAhvumxyKIQs8ypNkkofEi5mf
PQc/k0MvgJKywL60+3ZfLDQdQPVXJNLcrf0b954z008N4/B+UrphVg2DH6WXeZsR
XCMeo/Gztzy0jSLdxWYPOF5APZoDmUCinR5iZbHzgiOciw45Hmk6V2nGJcVAN6bl
1ULMAquTV7XsU8M0p+mQ294EZkl08h1mT6rJdGjIP7akz9+naTnhNCDWUxugpgrE
g7c/KSrSbI7qJzr5r4pAZU4HG0H0ud1IFkqrAN9G/raXGKcU7G8xvJnmaKqCb6qK
m8fHhzeP4VfVDOpsgCRH1g3ORpxBFCJ1a4OhdHd2u6UX5UkgWR5SeKUMrzcsCzKu
4Ly8EegWEO5f9P4Js3VcuSb7JUGDBCf/PRFVoOqRaBhJV91BetuNe2xLgqEkJiVF
sSWMgBTshr25okWzkRaIVQXg94D8al19Nkdmm8qU4Ky1L9QDVpIfttI8MWwnBG6u
fMZVyt1hAbkI5QVB0uCCJKfQluLWY8ZxWI3vYXf5Df/ScfoFtYHwgS4g6V5t8pvT
X6y7zTH5enkFWWS7eRz4xCCjHVxxwKpmH0VIpH2q8KVlrp1EgleEFCfmEkBt7xIz
JT/JsLcB+ESVtScr+0WYzBseUVbsiq3vDz6PvpgheCqBxvxGU0FdXBf3A1AEatp6
wf/jTkd/AzlbU2gM2tas5+CQ5UZNjz6+XKyxRVySLCPXBmQ8pVPnvvQ3Ui9bFGjE
+ZDsb9ASKoZeReuADtNfFWOSMcwSxwPXSiTvSlV9uJcaPZVjodRS7bZ6hD8DbY+l
FKUQRObehIWtlz+VZIlgALAkyC9FTpEYbolEfAjLbABo9bGxfhb4HbQXYiBuo25h
51o0LgNLYuys4hmgGDzIl3RIzYjAyRy0RivqY2VgO/RoncmYXHPKa8OdZgjc4B85
q3k9KBttGQ0qpmSTKkt+iyJbMrtM7nokCIhA8fzLJTzD5K9+I+48c8h79WqLsCSM
v68rnYjAqAukuG9mKBNyRfHEwNipGxGyGRtphACiPIyqCrBsKytALBdEU2pitqzt
FC6SoytZN/WQ4Udg3U2L0s1+jIexCNfQ7VDEo7+pI47jRWDJjowZ9cH4Tm2WOE8B
Qic1cGZQsyL27pdmm24fzvECvfDfdwsYhzZ7ZnJ+lkqvbjMbmCxVBvzmhRChx208
/ZvfuZN1ijQCPr/03i9+v2EtxFfgj/BzPresPH8FiwKDn+O9oR6GpndR1UpZBZzf
9WWChWq6Ht/hEDX6Wdh6/LSUbZZu5ocGlpO4VBnc18q7XHXKD1/wlf1GZcEgslYI
aaTpuo1zH82K4vCmEbuFgP2ZRvov1lc3vyAjwYcjl9N4i86uFhZkTY9jctMWykZB
bYWZUBqxW8XGwf9pGPSHu7wICSnwhuvSFwdGteXkNvMG0gfPUNvuKwDDmLEAd4ce
iBf6x35ITT+cktaMOnRtOsXwmEo9gMPdRvrZLgi30NCx2YBvMdGvYR9lis7K5VJq
P7wNAOF5cx+Z0wQc1F72/vmh1kW5LncR0T3ngvzXuWnIY2p4dUN5eGZtXKLH9mp8
pG2j+RzE2tS1SljCmTp7WE0tHM15MVVnY5IFHKlwrcmjYEmMgwd5fMG7k0drSM2m
R51+Meq0P0FJuZAAJRmyNjddvrWFurR//7zmJwJ2tcxfAxsJwiwwCNxF1+U0u/g4
9du+tANnFz7rdd+3VDPV4tOn6mtnWvyUFV5buhHh7C0Qz1oiR6i34JRWF7ITWfMH
uEzMWVKZiUEWUHiaOKHnacKDST7xsiDOvOfOTMPmGwK1pZhY4nYraTgJBlOKASEL
koKTkhlZbPi8+vgJcro3Ij8x7PpA/dcukTpS+DRveBgbrNj8YLSwBls4G5nJN8yp
ZaoOymsX1efRGJBkH5UrvaGrB/MZaRY4Ce/O9DinDmBN6aQhFatVRjMX6AupzfX9
V0pmpfyhCHyHcA5bxGHaXeBwHB/hi2PYcymdl03KoZcKNDZ7wt8s9CWM58XFLpVu
8hdSjhgO0v6f6seK4yBr2CAllklc9bL/x7xoCtO7PgV5LUbD1QYwdKHht3d39rxi
R7WZCvChgP8gJMgs3ce1jQSondEsWqznJjmJWI/DRwrzFf+eUKGzF56YN47HGYLK
hJR13Jc+ud2aKodApT3Q//W41d+Lum21nY6KNwpyo58y6tO0kFaD4llASI21Imbt
RCxZaCfljIe2YLXQ0nMz6VzHBJDO3DPP18TOAoBeA3/TW1PMMzBM3skKqhDgARsC
J/V/0GwrP6x5T3tyunMNZtiztBK5OgbXEEP53J4u2THK9bFV7cg5J5ZPOT++BYFZ
r8jCN/S6pTCUoAqwCeMW19QxZ782aCxXAIazK9kPFLEaUcMZaXSMfNoINrklPdzJ
V7JmSS5sJsUYW98YI+SV7baaj0V9McdaPacw/ISW5KiZRjF482U3xzI0nvkPgaZt
ZcX10B1xglifyOUGAnJ0i8DtNvRXieP4SdQhTDlLGN+zDqzlIMXh60tt8xuIMBIN
9z4oLDrXNKd6xhCfd+Ve+qIi/mJjVR/ZKyouxkqbb6GVn6dhRsNmyCUWwk/IdLE6
lBPQxLJJEfhdj308UvP6El7g63ihupohfJ3PGY9z3YsPalTMDu5oO2wKGJh5hAAP
dIjy/JGTDLWqX4RTW64iSaCJx2FcLQgRBRWvKoaY65F/AsNTIKv+VZSC8gYDqdmD
xwcZ+qu311mQs8G0GKhQ8+zsS3O8O2nJfWuutx+CbvhD6+g7F7LtzDqmF3A7w2im
1J1Fs819mO4820s/dpN1LKoZFldNspp3+xazDJNFNlpDBsWNuYzTFmxw+6Oq50MJ
XuODHMjfWff0R/y5k86auQ66EDsDkccmyTrJYgNsXTy2CyAWZnuN9E7m5yfDxzd/
cx3XcTSQwt08uNx9aSLti6semeygvwEn4Dbn8p6kJZo/RhTJLPll44xXWdvPSD1l
PFyKJXXvIyosMq7qh4pg8X9+wLh1gojQW5HKBJZ6frBSjdaX1nEryQ8keJ3vXQi7
ro/cpjB25FCz8JiVQYwlOU5hasX0elWfiwdRQZmSzUFv2dfiTPjSE3DxkCNEkHWI
21iLX+08s2m3dlzvTOP/6u6+eZw3Ho3nLTkLAAK1T2VJkvi5vc7SVcvrBIpVDWvB
nBtREJ3HMjTUVPzh59T38IhP7MfRf0b2SPHuW51Xd2zIW3uE3Whob6/pC7BpH14+
IwAHN2rfACsrpuUdyMK5pY8uCOgG57IbzxXh6lcuq2UCkJ3V4rCcWmyvFm1xK0aV
4lGYAgqdaeuThGjGg9/7CYpFUHDsOgB9RI+9AjA+EngrziPSPnzEnawMyWLsRH8/
ljMirGxLpzh9EdqSple3yyv7sTuOWekJ7Jt+sdN2UDnX8bErH00i/Tg8ueNM0gBk
fM5FxfE4n0tcoog5RvgwyLzSSV9jEFariTY2uZuyUcnHtf+Xkmm4BnLmY/eGMxyW
vPAtAX0oOroyeGez4eqGJXmLUE+YaBFfBPaxA8mu8aZo0B96rnfo056odU5giaZt
n0GoyU9SfeG/5Wa8OC3tG7zqxnd84zYFLMD2nIkOGFgoRcU+dWS1MgpA29/6RuBq
BpHxsGULHPJcMzPkyhF2+EGiQnBulISuIhdeaD9ZxjhP70gdltSH5eQMOJHV7Uuc
VaO8Z04hpJTsssuMmTYsUk7Gvw6H81pSWQgM+Knw2GKRREWPZ1Kes+qDZQikdmbG
BJkk9MvBRnAhAR2AmwG28SmR8iWKh1vv5+WE8MyzKGMZpMGqu0sUYn6GIaYz3zBg
ziXwFDR09MrOEyGvb7M+ZyX+riQYodF6kR6Ys9KJJHwgJyZTeavulWEYOkpfUftP
6LihFFIP9chjVmnlHYtS5D/diPHaj4AfGMhhK6WwMX6yG0Z2LBVtN7n9SiMUS9Kk
uN1blA71C6besTDLmaCOfviNuSgwKCtNOvJzEIT3c7gGS/eE0DVZ1K32ullfzubZ
ZV5hk4bbH4bGggUa8u9Cu6DbXbjtxP7Zvkk2ZeTmIGeS1CNrX98b2Ys50da/1zf3
nf+gAcJAKQEdF0+yOVZuI4wEbRLpON7naoj/sFNQTX4ZUSnOdXhbhgyvi421JMfW
PMUBYZ7GvXe6jKmlB7MU14+5VuojrvUbjIsbLKB0thwQ+P/z/Skj3H6XM157GzOt
YZhV9OOh6BWVOpVy91BMcGdPiguO96gcuh5BZJVM3froxHUaKOSzVIlCIUrM2isS
H0mi9qT9G9rVwvUA5Dc6jBmQxIRSATk9HUj6zHswhXz98k+7uRIm+hjuJVeB3BsS
7+T8k+5xTWrC4oJqwvFUxJqAz/2MD3wAMUPMICUYgrX6zRAfJKUQTFhgrid5U/R9
xkWhnbKepcXtpB39HO459wV4MKsLA91aX9x4/ZvPCLv0Z6p5pnLLT0VHWSEad/GR
cS21OHFFxxY+TVSOyaCwToaGw/aFUWaiyrkQzK29k01XmyAHk9ahvQhF06BgjrMb
t8h3So8bxG/Q/Y1E2M1LAfGkHSv/aoWnxduKdB31oevhzdJB87ut9fofy3aAwugt
VeZkMdx8FOO1oZ/3fu9ZJH+/cA8zWMAo7VrghY25apl9ybEbjN6VAUbrG1CjhEwi
Hd9NCGJiNT7kN8A/1VJfW+0KkScjYIEbFURzSFYG914ZM85sSaNII+5EfTArCDcV
a73fjKRKX6dG+o/x3XWy5mLfNLOQmvWujru/lyXwItgSJpJXCNvF2obSv9Opq1e2
vtPvphB3gvfzUwN2RJk84+lRUXGVS2Mv2pTbaHToP3Aj70k/t+BjwjclX5omPdXt
aH0YsEElWlpHn4H4gprvu18tWWD9Q9kqMif3QAZH5ap64UHUrathZ0FTM3IfB+xA
ftOjHQQppNRUnK3rQvRMElzw5S0fvknUKKENpwUuJELrasCllk3C+rbj6/nfCxnz
ucFcW08XtxhwzkfqmW/WUuj08ATSbWu1uo0lJ2PKx7H5ez/T4MUnVvDnjWoTd81t
Nl5dUeUSNQWC6W9zpxtU+1rtkJiwTnBeZ/K2NhKxXxoBiOhbu7y+t6wMRxWHhHnI
4ES8dc1kiHH979nF23qLISI8LcqL8GXibGJMt5LU3enk0zxCJVzQ2aVkN9gTQp7w
YwvqP7jARM/oRaqKquRPCpJWImux6rDgtB/pGoniF4A1cKXke6stXc9e1cE7Ziah
39IRlDioxnahGnAN35CEkQkW06nbQ5xWtjI046li6xLsJiAoQcW1O5Iv2tS/QsXs
WzWfmwAFKS2DRbRrXqJhWfWOTRbx6VGILagWzwyTF4jk542wBCpGKyB/4lAw/CoV
288HpzKLmao/0OiLDtDvxMDDhbdAcNyGU18gD8l4qlzb67uEzNL/NEzDrzIFkdJr
fqViySNAAW66RJNxS4ka9DV5GVIpEC3RcRXwOOyC/3svtup5dgOsGYQTw6hxDkCy
wFuvwo4tBr70txQkJav8Mwy/+x1761gdp6w5+DIoJSOikioN2zx7qm5lgPpP0jfP
PXRVFE+B+irwa3LbqJh7NaApULzoR4AeNduVLI9jV+kHmbAuv0/YYvJuXk7yucMd
nO1hGPL3YOaiAc6B5Y7zlIYCvhM3+gNnpIyBos50osoFY3kJrq742VLNt4qo6pvz
YJzI+6qLw2PIg4+Cqq2xEdUlwoq4lxu6+C9f3dlBuidI8LC9mWjI1ixkds10+yHv
34ZklqvJwrf2FWWWn9sIngCGLdEVjbAM1RtdTz0DFjprPsmEfw6GjpPXSaD3svUP
U5eaufrPoPQOjRDmlj004XWjmKxICvvs4GNoxg56qpn9tboxrhChkxbLddJNQB35
OYKBZ24C6zuj4KC2B9Dd5glAu8DbUgkHt/t/B7tf2mN28sWcj5HtPSB4NQ0xOh7l
3YAkNBWkkffwlglWqLryTesxGem+Uvm76gaAxjcZHdv+BFf60T65DOnc4zzQ1j29
sacyAO56NOXbgiliZ7cRQzMjDQMm+hWACEd0SFJ7cP44R5+J3ts1PMXHGbaH1u1M
9DpJTp/RkPkboZ4/d0ArvUhe2OaHGw/FkDW2PtNAYMXlRswdBB0thxbM8/E3tA/v
jA1OY75aLmSp9mucTZx4A308apQ8dyisWJlvRNIulY3MmqPqhvEI2HfBJHd7BEiV
eIFzvOak9EqI47oIkh65dbM8YLQGE2mOh9S3oiHNSW19fywi8OlrAIwvd2AmxFOt
QjWsvvZGrMsgLScQKKr6W9Gwb43PkWZKSBQCnq0QVedDuddUltVjijSDQH+RjHQY
6bNrr+QQijFju1Vc+QtoGWeMQeZs2fSSRhYwwLAsfSMaK5w7xoQ72is3a1zmvn5E
6ucfqF7KArJu+02hDuAAHXYo69re5p4ihqKodJPSgzsI2RhwhO0Hj9x3mys+XeaA
fLPP/RCycU35c+9ICbAiNJ4rlxBostgcUW51qfBY0OnLCwPwMAtrkuh0sa0af6G1
7JuXzvJOqJu1wlIg9lWeq698+ICf5/brJmtnnw1V2l0iRro3aB8VqdLUPcViD9mc
w9VN1OF+wdcCFyedVgp6moffvkqOsMOblohqOYu9/FGFBDllEQlAILisp4ryGp/R
0oCg0F8/RHUYLvWADNp5LQ4MvM75JJSr4m1HUUTwFKsinjw6pgRNjY/dYRodW8BK
rU+S5XGrdDvNDAmpuuQOuK70YT5KFkEvOjj84l06i2fy/e5tg70Jb3rL7jIPUiAb
B6yq2qW5RtjjVrg8kv4XHE808DQJ2xv8vv9mLPo8qbgydH2Tsax82yf6cnmAaaDd
g7RQ5lpJqUzYliIFXfxwgZ8/V04LX8h8lX+kDBOj2Pz1z73cMZ93LZLo6AqJA3Yb
Bv6D/3L1qTDfmbmXFizpiis9CUmld/FKUhpuTPq1pxL13vhb+Xqc6MN3kUxYZ5w3
bsXqGRhi4ZHIL/03beTiSjlKdodCmj/FWFLSEmFTZ0CQaD8vBnmGnrB+ibl1dD0M
XUYvl0kW+HliSjtvxPEnyZDR680nj446kF+VdAhSgU9WIR8Xq5RhflLYpqUczRcd
fYWFBBg2t4PuV4PornkKm004x64WfRZN3Afm6lR079Gb/VGPCNiLAaT5kRuxDFjD
6Mj4qwRmoArb4dzIzqNEJo1rWWhkK/mKN8bIO72DaSumZJ5iXw7roRnIFUs4+49h
SPp1h56+lMiAgwEjy9WZOyqwF7rqg47sP8C5Fk36JWlhInYKgEA5mBb+RgEp6cEz
J4MaXihRO8ntmbmTzz2+IUKygWb0Dz3ZTyJoVRh/oTlqtJMfx9HvCH1UQY0JzFNx
xpK9+7yOZjPIO/VKAOf5zpW+4fzIcGFtjq430AjtASxGDOIXZdGTA8mn8aRC1Di6
yYqDIBDNlPPbEGKa19T507xEGwlixFuIJIAwfdwcyX8r/AenwYJ5uksm5bQw3gaR
HFr9cztlbKAG59HW5NmbjEfsAZQtvpb7QENKnfNWJsUH3kzAj+4K4hLVcI0JL245
sXMI/m4MUiNvnd/Y6zZENMrTSyZcla0u25Iecjg1bQEASVEk3faLph4kRZXKjItj
OOXDFTOiFr+UgpdeQsxJ/FPYuVwo/7AmByKsFgDTZo1h+DHIe5jE3N30MU6c9TDy
KlwqFbFwFU5x5u/7xDmm7b2pVR85ReiwlKiKw85JvmdCsVaTYAbeelBwuZUq1WHY
BU38x09PjCWeJZB9t1shdpDUhO/Iny5bknr5Ju5L9J1YawjYkIrwr0drCF0HMAuJ
CfTlHbSFE+KlIascP5sOxSG2tGKsOakg4BZRrPQcJ55Z7EDNk92haMzSKj3JxB/7
bo7ZxTF14fsYjmU5aDsn47QVVdGWnwR9lJzrJJd69EmT61lAwcMvvcq9+N7XyB3R
a5iFOVrWXz4TRjFMTXu37gTOC1KK4nnxi9k4MKdFmiwy8ApGRXIbk9e475LSdIQd
NikxYuLtFLqjvq2P6Qeoi1Ip/xkFPRUcLrf4GE3NSX/jYCVQBpxLxEYa++z67L/v
P5Zq+wm9fsr9wgLnLSM09DNQiqE0m6uw0dkdSoYlG36rNsfU6QT6Rt8N8DLK9g4I
KkLsF/27Xux4Ik/uaDtqBbN/ePHz5VipYUs1/1hNN0aayJJRxCQQEHyU7B7FRI0c
IJP+ExSq/pifU9GK+LpsfRo/aVqqEPnEHaoHm9HaxB5x5xqNbr0ol4J9otNwxpFj
V8Qx8YxUljyS/+6JjWAraNSnicJCrDOS/pA8OPMKIlwx5enOuS2h9YTO7M5LPFl2
Vb8hInhGBSCQAcwGzyQNY8chUH8BJWqZjTzbE+z2HXUsDSVlWbPoGeZwriO8wbZz
qWEtaueWMrWUHiy7Jq22aQs91Rz/J1iwbIaeusImH/jy1W+dXOSFlGtz0/iEA8nk
nTQYeSGHMyv6qIKhXuvTjcLly1mUUxrda/2gxaIvcv11OklkZ3zJKpuigGiDDqlh
ti4tOZtQ49mlCY0zJTi4Qx4MkW2jjSe/0pwEFaeECvoTOabeDPy0Tm31ebDwhE28
PpL9kVaBOeriIE2PTzM2ONo8TdeRWt3Mx2pwPda85T8p2JgIq3/ZwyW/ZmLXh640
UXWKtyh6F6yrjzpEECNuGR5wopbnkYx3A8GxAUZjB4lcBkTdkh4C2QmSr0WZ+4PA
7qfwkHTaKDIbexFi1VZI7PDm/ngqugBFdPTFHfimE9vj53BpPMoYjP22Rqo+H8HC
bfY/Tb/uFzbIwCemHzjeA2H4Tel6AReHOhWLaRyBKOUIrosxNkBW2H7/oytCHfdP
/gFJEIUvuxafWneOJsEjqqh9nQPk7Y/7hxM3Q9zg71VsB7bVUWrkjfzWK69BiDLe
puU9XBCBavzHS7f94RE+WvsDDOLr78kgwJxAq5SOCgr8wDh/vV8xYKs+ZyicZDpl
kK1fRorMAoaRTuj01+MavZmpNXldUbZaMt20ezX4rSacDQfTl9D6TZ0I1Nv5O8EK
7k1PxqcUUXo83hoqIH0tzLMnwQ3h7Z493zTkePMIgko/tUqCDHiz6X2fRnWqWI6q
pzuzuxo7I14yv4wZdUC2GVZ9ni3AJ8+0Q6L0Ts5Nh+Hx/aYuWTrucMkbpXfLXVSz
ykTp4GWGfpsGdLquExdcD4Gl49ZBF+hgMbIXRqdK/HFtzfrKp4m5/mZfhkucXTU3
cCxBscm7H3k7PsnnZ0oG2c0A2/Nz6HR7GpdWAggqW0WG++Ig9lBsHkSaZOOHU0Cn
70RxowGDpz+PG7Yf86dNMcM6R4RfOToPjQaSuFX5JPZtISBDh0/csxIABKWz03y+
/DTM9jLrFp4kK+I/mKGgbE/sZjrrAZ/r/sqJDadSIHTfSBi8/EYxG107wlla9qzF
0wrJZIlhrOCggTto+cozti6qDdsTtYs+wWvi2KFeRRYR4saZG7bQ5TKDty2QKqpJ
pwTE/45o8bdkCkVhCC6lG3sx8P7+X/wtY0OifhzcFqKwsTJWGcTxu9Zjr7bc0owt
AXiR7aroBsooYNkI5NbI7+e8blG4sJGcwf60cOkNyVJCxFzKZqR3XkjXWA+k38Jk
sCe0jdOS5PCJjRYeEP4XEacdpdqahkfqwKV/rdxASWL2KEwDBA7bAKs/F1quWk78
FDY+MEvnlefFVb3UKujeX9ZYblWP6QNchq1+LS/PYT/1ld/jBuPY8/sFIy9g9N6m
g6MavhOKDmp7jeEqw1tp2cFWOMmLNG/Cy9vIwX9XudPh24AwY8/FlKm5P8uq8riM
bgQmfYo9LmAwwUebwJ6fhahYzETrnCxzqe0u7rCRTDpo/XEosYWaPM0PkTGU9cZT
3ocogffnEjuPX1sZmzLfKWySpVTSl5VRRerXh43swtHX5GSZff6cjEGCRxRD3sN1
CwrUlnA3biOccoLkGHatEr9PxxGHyolzRnbzS314MdeNMyMkFnsJBlR9wbn3RzV0
wyXw7bspWq+ACtgijU3DKjMN6nNKW73GT3tpNqKJV1FcIlCe6sCNo4woW14stoM/
bTDKoAMfPVx37LoR2wnPGyD1kxCwEdDTYeZnWMvbqSSkqDjAY+LWIbf7oddxvnb9
WqSCq2ACnxop9BY1TfYjB50HUGxlndZ+XcFbyUFoUzvKiPIjNG3/hzIo0eS/mbiA
G1zcJCshm0dlibRCzQy1sGZQcVj2QHXajPPw8uGQbxXkkt42U1ZXtfs8jzN2k77n
hiKLzPP6Dv3nxGIMeAyW+vft7x4v0ibr7pBCiiEjsk17TWDuaBixdVHVyLaYABqF
1+T+1Sj+B/OXu6p5puT/fBeE+/yMsywq9sz3s2FOuf0+AS5sE4kLKF6Wc015L237
vHxfaMr7SZcuJalWkWf7EgJjdnMKqL3fg1e1BTmJXhbFE/Hs4a3xaFlYFiw3BJiv
1+QBcFO4YfO0UJ/7Zs2trCvKZCXF8t4IQBvd/2w+Clt5EhLbGPpdT9oaMiscwGdT
VqKUecliy9BaBvtRdDAyuHzdFfueffx7qX8JmqUfAPOC82AeVBVpfics4k8ztkfz
rdy8EBB0jqJvheX6eSNJbMFZJHoJaFZjdICSVTlrO5Y1eiWt9C7udeXizTVPwsWY
9/P1byWGFSXAqnNNYWGr1YPGBkIfLYphGKmdplza8GVSMrtm64WDhRYQLgphvBEn
AfZQ1PqgnXc7d71d0A6uKonwFWJ3gsOVG9w/1E6YLHauhIRD7+dKUwkZGYPskhay
IhWTY2IRZNgm+sC/mQ3uqAMpLUs29g0zE6044exUcY8ITmnXjpw5C7ybkBbJcvYa
OA8HVzR3Ei4E4nSs7lO79hcST7J9uWUwa7XvXR9nqteWvfef4ya03p+lM1ixmcSW
A3bStR+tXEUmUaRr0L0YDRxFgWoBKJjcj78FowB113NeZcDd447SHtEXesHxCXk6
gGUoFNf2KSEtpBVntIU31OuJEo16Bwwblcxm5cisUWBBFXAoPfu+xaihHRGt8ky2
Mh5rpGzPidxdHuAbYvdIy0w/ILYrOEdLV9FcmPi/jt+/LfQ3BTCV7+VLNcdnHxt1
dup3/VjZ+ftirKoXZgtWi+VOLpDoDljQCVM5EFKyBDGDhXP33iqpeKeWNDAPqcFS
ihGsEo9HNoEuu+x/JbLDbAoYZkAaN1sqKSlIGLPMTulhETQiQcxvKCnloD+LhbNN
FV2FeI+zl3Jq2fvn3sCxJ+LwTRxJhBoSvQ/n2G1IIi1/DXZvUtd2pHiP/bo4Nqco
1TV6Jecs+g06tCR8qhKD9RYG9AoWsu5qBLzdtb8pMuSp6Z8srmOOMlt7R3il8arc
VnKoFafZkdTzDw34bFL0IUI52CodaSmQuRzjcOOc0SjkVIFQDXSr3R5SQpnw4XH4
oMJQWbHBYUrIO/Sezf6C8QJNVqECTYYEsBC5LSmst0e0UbXghtFxav1jwzgjDD2Q
T1TCqH3gWir1wNZ4UgLIx3EsfkZrnkL+kXL/o/+CVfoInCOYuTv4lCKIJ9RzciWB
YbThaihNac3ZLPbZEfex8bkRUu+MVx7VWhFlS8NtTQl88CE+3p8LhBbASuYtOEIA
wdZRPsa4Ho4ozujLRWcTr7EA0eU0AjouiMJGZa67WdAm2KkMhJ0g6BuxSM/lETBI
xWtDTEA0Rr+6Ix/XQqtVAiVMxmjhXpcbHQMBTxLxStKQJw/5tXiraPe8+xby6bb5
6K4346/rVDVsQG8tCZxSpgVeQAnIKvP4CvCOgkhoOTMsvVHiNrqWfUKioqP+gM/+
vdiPL46W49JpLxTg8djy5yffcwEbIO3Irn5Yu3WPMwVGlMOXzKWnX1ek+goD1vFX
AEyqv2NY9PHRxPChtZOvFkS2ZbKdTsbmEYQgK3ZAxWm7udPwWOZaZwRc8RL9W9TC
2092LBs+bc7GIpGGpzTAKAp6RR+070XUO3h9IBT+7C+e6ou0Ka1L881iP2bgHvcq
LGhcHlJivl8IqC7SGn0FSjRRvmzq4nfBSNfk9m+TPzEr2tDS675z6dyEIngUgUlB
cwF64zPW+QffcAzCISrHxB8NwZ0ylas3e6Bwl2ZWQeOLSH2cSTrSKbzKJTgIiuk7
j1shofYee1craxN0TLzRyyrqSsMFSOxVfBkpX9F9Ga4EFkbKCs4/U7P7HzN87EAg
WonCpkeDQN8Gwpv+bYiWiZAFgEHCTSOEtQiB76FXo8TfAB/wQPoN6M4AJpFVpsaL
CaW/e5kPEfeWCaw/xHuI3ArKMLP6EF4dfxC4yFObGa1G7MGg3ReWyXXsxYW5OfZ1
i21jMqrflfuqRX+v9dN72YpNC1Thp9Zb8mGUw6rQEOIURvi83nX9zee3y9m+7fN5
q6BowiH/u4WuWQkyAKz3DJ9Sw5WkXaqJCV2+k5PgntMzrXAAOb690RkaK2X7v2N7
64M45yHqq2p/hrs3gjZuv1pR80E7ZZV3YzJIrtq5n5wPDUaogCcUAxTK5njeCiWw
hzBr+5rmiU3dZLcA7dnqVSSsWudPoFMznXAa74V6E6wyAWwmdcTh+Tv2sgG6YeYc
A3j5Hyxl9agn0BOIeWnyMvTLk3D/2ac1P+D2r5+rFDR5jbjElS3gKoPt6NMK4vet
YAIU5GyrhUrmEdxv5V2vWaJGT9HLgewjx95jID6m3nZsQRR9V83ny07OU17FAr9Q
fe91kQH6s9kOd5IAwZqPbXHqTfNT5lnap3OLxrxCOliONa0y3Y98bddgcOPDIOdv
up3bTcL00KmRllRIVoPwuBA7fiCXdgDmPmrwQHCdi9cRg3jtPvk6fJ4NfcxSJfmB
H9WmroIXFXuzZvPmd4p+0yZyLiYIQAILTuPeOoF86DktLZlNThobXgU683cqDG2I
FVkVc6yPqzEnnPpXg/IoTUrYT04MCs9ELBpFvz1SkNmlyvHQrD6FORxvl/NLdRBl
jNSGc77zMOBD2HFOBbJa10j6B2vaZmGBllgP+pXKWFu2LO3r0hD4rhBr+1JPeAKM
69CjcW/j4tcGGpSyPWuHoPJH8BJmfNnzBGl18w1O/N9suBtwBCq0sLsoqMtCyyZU
wXQQBH7/Lbjdgk3Q/zCjmVs4T9tmqQdBFS+cZm1fosjqHU/qyR6INWVrG5Wyu+ES
p1s5DAVazqQLxZSQf7pJ1wl2kd0bRFVBcLuQnjEc7qDGCWgndUwvls9xcpkc8L3C
/S8aHuF7BLi9QdtZ/uB4kHzP/TNF4kWZsKGXpLfQ382wNXVKlLtSG0d18zkcG4p5
zGxDyBmPjX03VzaIZ8/FksELiouZj9x/W3h/mwc2Swp5dQgKdcuzoxSh4GzZpmKr
scOIPD4Qi+0R8iewO+3JcAP7Q9NUH/OiHl64QPvjGbH6oaQTUcqQl0gNn11zUjHz
jxHrhKnKW0N693zikPgX15mTtmCiZI42A+gmKx++OtKfJId6V9KfQ4LxyralcR/i
q2MLgvsB4xKf0YMcX6m30DzTMavEvSC9aSkrPV2yipu8nKv1Mvz1sX+bhMd1rF/V
BLDOzdoxe/Geo7DvDI2FZJyaD/SdryXQHFRYyDrH7G2H3N9aCE1719eDFHFqLrbP
2ViRmHMcgU1VwJfH+ifYM4GXc7V424sGSUP7R2E4f5qJY2mjNl++SYNxRNO3sUb9
nf4v45tKK4aZ2V9/hzbO0gq+2+Yeqqqte7krZ+W+T1kQzF45Ek4q9U6GZ3VpYtDy
QVdc/lCxbn/oI/99VbWBbcaT+T+FB+39G9iIgkd9p1W38ekOpcnIMLvpfmbx1nEx
rwYCD4+TibvlYmR8YLaznFERY6U3bQzbCztaSpOQf5wp2+Z8dJXKIdc9nMu/oi4+
mjOBtJOF7sxb1MsmlNzJqCYF72iwS+ezI6pW6RwW4+YPBic5USGq5rBA1cHen34f
4o1+o33pHwFvO0IQV46jTb59wlP7Gs6LnEUiWhOf7flmKcnB0sDffOvrq257eI9G
/v2wyPXKy0ERbUwtSAX2fy2m2bk/tYDtyhEO5WR5a4R5x1SPErdQRhbCxHmzj9sE
e3wQtJqoujVP0xLqlaM8gI4J5WXA5OuUglnLXYVxabsd3CQqd54+1enqTccpjeSE
dIG3EblrTjO0KAHzqLqfUB6SetAYY+5KqK2GUrb1Z96PC69pvZVrBNtNsnX1i4lN
5VXz+6CxYx2b9Fr5cqc6rOwZJfxk0JYTdPlPZGd4iMityP2/rsUYRbLB9AlLIZ4A
FZWSNDmRP0xg4n4084Zz8Midq4ifToIr4TsBUF07W6AXI7HufZtHLcsat/HubfBD
4dBzRKCea58/hvSE8NKY+G/m85TPYCkSHl2odZA72hxR7+aZxfE/y8phOo6UD+sT
bcmBD+PeOJ/kdYaJdSBd5tkI1qxD/u1X4yegN6+pu12BGT96trq7hKUpiWN4GIFK
pBnl+TVLQsbna1Vcb0XH5BtezyPPjDwhxZCDU4CyH18KlpDJc+B0nHBlc5iKlgct
gKrU9r5AiyucgiZ5JuCiasfX/L4oQK49JcH04HQsQYVNG2ojkJpZW3DG/m29utlP
9Nzvqmpfiy0sGwcGVrocwcN6uLLeO6X5iB+wsNRoD+iKPNDXFFHZWc7VI8Oc+hnT
vMFxcGBPlEUqdVJ/Qj68mMUi0Fmutt31CTPTPcW8Gj+/XKHSh6xUkZ+ElQXb4qmv
7X+HZQiEj+yOVM1MP8uREglpIF5pCqXMNycunRWKTDZnFw1Sw3j12hO18jOOKkje
Z/JMOCQO9wNfNNl85Iyv0FeBqGDcalQmOjqo8aZbBNwL+gABgWgGYbv886bBrl/F
djRA2YKZfGMt4Wffb4GuZW7PqRAz6CxXo4QdhhZuxWo9J0eCXkhWM1U+goWv1Nsw
4CLE9IHbex5pnLXxe80SJqjO61exAEqcImx+T1RGNm/1Jc8Xv7hSYthwB0qnIO9M
QlhNakIMZIaX6UEnTUxv3eaPAM+9VkjuqQFDjPOxc34jUtCFEU5KikRCpQJPTAi0
ADZFKzXg/rB9nprO3v5CC3x1EwY4L8wJwACIkRjQFyofh/OGfbpD3ZsdmBl22e0Y
V+LFRrcPUj7FBS8igMS0kqi7/t+RNYcedZajP7u69Fv1ehI35c8r5MYJgY6zDkFM
oAbLJdQVqLiouRjmJK2llK7QGD3SZPDwSxrbxLsWakjPOS55VNfgxrcRKAKHr3DI
oFBY5l1uqLjpNsp7JjKcP8mQfotiUvajjI/zzfCj0dI+aK9MorX5qTBvOgE7kXTn
8wgdr9zMm94JhhO3f9jcLPiO/MdXNeWGxVArIlKNXx8HrhiT5n2T50zaY0SfB+WH
253RF3oXn34rgu16Hjk9rFrcd4guj/rBKXsiWBz+WOPrTawpTIyZ0F0F1TY+yAbD
NM8AN2imeUjAKrkwwmd1Y9kGeiJXWj9IOtJcsttTAQXEhF92sPbjRRqytsWVEAR4
7rYH41iUJ0VBKtbtTj0lVFv9ZNS2NpiVP4xrUTgKc74/+TLmarB7bQj++hkk1NHU
t79VQeJVMzQKeu1goIq68zVbX+Q3PH4jD5oxJQfMBPMB+Qqfttb2+3bexkqjMoTp
g1T1wfXCkYdjKzHmWCDD4tb6c1Omd8QKqyj2eZQrgaJBRGkTyXn+OqhINQaM1SLU
f/Lm/jdv3THHn80oVg1kI/yF/7ypLmRgrSdwxCnrTbrBSCjM9sxFg3/EeJcl5u5C
7fycgwbRMkkZCxWxVdqiArYv+lDgcjDmTouJHwmF3pdpZGdulM352kEmLpqDT4tk
foP9n/MOzelF430nnpFw9VrDcPSgmuWeC3piFpK+B0PXa1MjGRbfgMezsD6bz5iO
cNdk+ZLZrNZp6soK8I9B26skXOteqnXemveHeLzSkfYX9SE2RJAf7RViFM8i+Ym2
po9DazCRBtm7ZsYZnuNymsCKOq93q7tO43f8B0x/SQ5r1MxQaGT6HE/V+Y9ezuAZ
jrkzVmRsgjZS+lenExY53rmMfnYH4l+dLH4dHrP6aTdKFutYjGSPj8COefqEXY9U
lwzSS4uyF5BySi185o/0NdjIsWGHFU6BSNJMOvz+oVrX8Chnk2l5JCHbZ0/MhhDT
ObTYGUTgGTO5CyOaNYY1jVi0rUiFqa5KF8qMrnTX0EBGpwFXiDBeHda7LnzBySe2
8F2GXrjxGrVC2X2EkxI5DWuqVM78hY6r87jvRhIsu26xclBxqZnt2cc6Bylejuao
M19HNFMHieOGOcdsLpiVyyeBHLqlemNz7KktYpjKvCSg1LpbsLtt+iWeyssizf/g
lmhMNGrm2J7JkT138wumwg7tVkv106E/wc7I780zXoGnY9APVGD+kUQBc2+bpU6d
b9evKMzHJeQx7lZw26q0gXWOL1OCJIV3/n75j4fOGmb8Jg3znbu7MiRcpo0FT2U8
NiRfzCqecX4WagRS3HMhYzmhuo3TPJ/VpMIJwSaQ9XjZPjNF/7kd/8Q0Sedyz3lx
ZnMF/g3J9F5F8H3qU4oBWOthSRxXvWo/XxwM3/iCvdh00BEGjw2Sqq4XH9tBognX
IdJgDxpCVDNRr+snFoNm5zE7NLL8h5rjNVqgrfNh+aASlZvKwFFMT9zq5Gg4DwRd
tV6rX8hYEgtMpjnYZaRTFI0DJXZ/lh8UQbHMk0wvu92ATgSx46Jr+R7QAtGkZP7v
AD3ln3ZsQ/DCPlbuX7NeqViYDrq8F4Yt6IP0W2K0zINkUncOF6jHrA+pS+qAYM4T
u9gmrmbk+BqQdQWuXpnOi2yx+HXK7z1Ln7TKpGzFQtcWMYWO4i/MHZgfPc6C1PtV
PT4qo5P8er+fTreoW0Ef+TXYdTD33gog71ECU1MO7jkNgT6+ssj/RTT1u984BKAq
HYKGaFlL8o/AoNeBM2FaZfEzwlrD+UI0Bl57r3DzVewu83bJWOVVTwhc0AR9O94E
y6PfFW1+AE5wMGB/evLlMVEWdOYZimvN7aRACZ4k1nSO/kMfiSjSV5Z2dBhqKUar
043wCckWhGitZhDeQSbH0HK8WnzSQRz94F7BBcJxaFAUylijp0189JfceooPEKQ1
GKj6jmJ9wPs2IU8LidApTPfQfafGs/Z061ONxiqTZM0WU7bcOQb1TCThj30HX7Sw
e4u5TvV83W0GFNdPf9CvyuAg8DB932N+wOY2rLmcUz5+rPv47pgID5dE7lIW431o
AIibSHwFX054kyOxHUx8UAd/8lr9b1tBCKV+33gaKuvkb1hTJ6hGgaBW7YLbrTuy
siggCNRphjRulCQhW54LnleEuVwhWVh2Z2pkiydt1xDmr+YCqWOStln61/xpjsiO
JSJImfl3TvBD5bOG/FrNkXrX+nDdNReK+IOVVYFptSpzVzgHWMvhyn3wzKASF+z/
xzjTjEWx6b6NM2p/lG+QuTwgoXrbBCh6d6JqparKZin4X51Auc2y7NEUhPXlY9Dw
d1nlrVRFpCOWPOjWBpAvI9BDFQVnqdD9eJktjAtT41VZb6vNJE3sPpfcCjWsUzJ8
+cqcrkrR1eP+6TvSk/YEC8RHDG4WrgME9nQ6Hg5qZe78IP9xNJ4jOoyEaiO1r6oE
fLtrRBIOHyODjwnhnTZqlLYO3fZXXP2+nGddO0gqpV/w/y3ZY7xJszi1rVDpafPh
EesusYGHrjB2Xo4xI9YoMGuJEXb1YYQLRdosI23SZk1SdLqZOwewgN73ZG6zNfFx
CbexzPKPZbClPYcBuEosJbRLcoKPBntnQgdNFP3Fvxv3oSXXrAqtBRIw5ghlqTuF
A6PKSsV3K08i0tfoiGa+CEJEryS1P/W5FPQhbJqymUdUdEzxoNCQAvtJMakOz4y/
YdGmKc3TgcqqZLdZ6dULxKzIfDfnEu5uTiMxDA52zxNVRAg9M3Sy7Y75mbxv9sX+
EjDJvqrQjHo+dru2PCNK3wn2LmqQ3PuUm+lh+Rmq2QmRwNs6kTaNFm3Oz/G34IuG
2rFMK5HTWAgfWygxWNGTDSAiTfogcNzyAJiuk6cEi77VtpOTD+mzjdNNQ7PTZlKP
GhY1/N8ulzDBcQPf/hrSvRD/zFAYqgYpFAoG9qlLLWpUMT1WFnT6z8JDKP3ywJo4
ibTUfbm4eeQCk/y/uoeFkRgG370w7Z/BdCCG3ITf9LjPRjv+lGHAgkjmdQF+V8Z8
+sdwX9wwtT+c/9msz5yIJexh2yQcfiVKRayCs8VECPAAfJ2kRZzM8uiwXc9Tq5HL
Wy1L1JGIICu4P/ncD5m8lKVZ9Hyv1c1KDcyoUYwSEZ0RZgC5mYvCNIHCX2EiX6R1
2tPEZXGs/DZ2DVFhKLv5s11NAm9WgNMaYW4tSQCakMsVURKPaQOKduvlDDcohOYg
KD9gtZUY6O3sptkoI2rSjQ/uA0U0WvfM76yULi674JFUNiB1AREqpL9hBUcDzEu0
rrVnmrczTdNVTED+VrFsICZWakh9McEsexgW4la7rnzgEiQh+OexDV1nTLBEC9tG
bdEk/q8S9E3ffJE9myBPAVfg+SoGLwZwuIf5BlMb1UQj//EmgWt2pORJY3EVPr3u
/19dOmYW9HLDjhr1cMNiG7cVE7JZeX1+7+mwEgM0XFbGQktAJcNnZvEPZ26T0ho0
y1+eCw1bAeXDyVzN15vzRi7fOtGwPlB4mbO/OKpipLUFr/yoRhmG4bcfCnEeGzXL
9m1QbRQf0kVPOEniLGiTM/qlA3NsKHGV0Im+tEaURxyH0xj/ThGK6u2IqqtaMEpl
04g0b5Mg/CGfgQ3u9R/7u0/5Og29zyinz5fJ2BOuPusWlr9gayr8HCPhWF/SZV5Z
s0/pcqKNAKg0IQOeahRw9sUhQL7sl8j7BMshQ+/wOObACLI+mYdfl7uhw6Pb4cu+
H1Tcrwr1cr6j3RAOkHPrAjmFZqB0Tpuk7WckhRLtE8ml4Z238Yas3zJPp+4hcTjx
ETWHecaB8d9lBL7u6l4B6bIXUrimsYryVy7iv3sR80iOBU4Lyk5RFnIE7LlPOJrp
8FmJpZpxv/Ct1y7vOWaNGvXNL5EwglUoZDUg9R+hBU1mopsTfLW2ytlpWN/yL71v
ufV36uEEINeg4XqgM32V+jCDDymU4ek+1SYXtDz2whcThGjyY2gmks86G+JMeoZn
/c3Ay7wCWI1KUFUafMTLlQqtbQkcTlkhJ/MPdWjwpmVpVIgtH6Y37H/d/hurkcUP
/0ZZYT4uMGJjrZLiuI8klRMItfi6QcMWwCdNkUss6FAr/pCSfr/badBat7rs7cC9
cq8WyWrUNDkKyxsLyZsPC9VUcuB80jopiggaActGeVHLtg5J6X0kUIR5844dSm0s
CbQpgZ68wqATwq6nxBn8ox8iEx3daXruGByM/YEBGcKZr0EdUjzQJToC+f0NDaEs
2TyGxTtbKhDn9xik0+JK/WVReCfnRvQS7zIFOpzXfVdjAyBzIOZoHgLGxoshubXT
C1bsfruCwXhpmCRnybh8gubNyLhnp9SRM/aH5EieydB8ol7Z0yTuTHd2qos+vjUm
TDgZfMqdak5HBaw+vWT6FsYYbKtU5Vu5tValcOfcTWqFycf8Dsbhr48HowpvIcv0
SKTJLkyhbPaWnTV202WAFPjnMpP1F7JmEgkqCZ4kgEiuAuwQPFoj6wU2eQIaET1a
FFj+urnTQq9kxbj2WB3Jcx81l0W2nrfHu9Z9t3WBSb0+44NqBAkNvSsNw++GIkj+
qg6o2rPs7gf7lH6TDtin/BBQjRUuDwOhgzCtiD8ypPeUZtfmvd2SPOGDqm40ZG0O
w/TraC7f4puLnbz4WoU/NsysY2vhLOsvRL9NyWR7KyTWG1WrLrXQPZNu3dlLgIoJ
8CBP1ZwawdLanlvxZPKsUahWhscQoOzgjEmWOso612arz5f3Gvq2vN6aX1NOGWS/
MG9Ulfvlpfi9M5RwladkhyDVmrEUH2oy5A1hh86SFmERx0aygWqhG4CNsN3acdGw
JzgtBkYEY39kesP8XBvzPCTJc4X/X1MvjF0qAubdmuthG5tfiOwmJEsOH2wDFAGM
ZMO4AbJA31o7C+kAoGlgOocR8QOeAjAL6lpvv4ueDAUIssK6ZW8ZkbKXMzh3hBWz
+FYaOirbPuVyAXwm6Guzm94XLWzGrAf/iWwk+7Re0QrolaV80Nia5Ie3PZaIFFuI
1fdS0EROWCy+ANKyA23D8tA1BQtP3+GjKYSrDHTUE9qsZyqPCf5zksEhDufji6Eu
ledNt9ibPeXy6gbytN5luSC5jUIy+dajNzul+d/kIxlgodiUODuON1wieRMVLWJw
O8py57Qw1ED0GCbkJQG8g97iOjMRMD5A8q5qJ5WCdhGv+9RxUrtwmvS7WRuC5mTI
p1MYblYxMq5e7oHVhDC42QepIuw4AHcPNQEurYw7rX5Sk4+k83hu2czAgelrtk8x
/W6Wsssiu0av4T256l9ol5689n2CsEOFBmtzU3EbFVV7zihkbVG7cPDS24/cjdkh
HG+qIbD5pbY90wF3EzKK2pLMqXxHfiVuWojCxDgdqgOxPHbeFa9Sr4OA+dOEXZAz
qoRItUE4msXD1hReDVP5q/GT/92So/+ow3sbkKDCJnbw2jZp3mY/c/Mm1DPNzyIJ
VMiI5dSDxwawmPfIkayqeyeP6IOJ9Kyj+lf0ThbkcMpbNioHO3yUnYCKqH6vSkcR
371oklHLR+X3tDeEktBN9LXUgD63ROV4H1d5YA6i1XXKNAVhm77z04ybRYB9gSuc
fYU4tVmWp1wXjCCSpshETBWdpe4QBtI2VSnvx+CZSK64aDrtiNPjws1IUXfMwfFy
ZhYc5gjy8bZynbzaHRx/gXrjyjuK2eV1HWx2qRHso4so5QFCPoHtJAdiHtx4w/cM
IOknAxafWIbdtw5kQG2y54a8SvNL7Xy06bc19C7WUcdo94ASqLN5I+cZJsQm5RVI
LDiHgG46x3YYDiCUW80dusxzE/UxrMmyHXGaCnByAPUjGVhmnjjnFVdB+aQoHXzw
B9NRzcRzQ150JMeN+rX7ybvhEpo0WcAjYh7PzzveQdedoJZMlISEgUlxd+nV79cI
DGCbqKaUTrzfcJcbFInpvNqD1GAAqs61AVpqnORuTBuwHCIuiEmafTg8nVVPMIV6
zKs7xSbdz9/nZ9rTtAZ8FVb8d3/cb7sdqBpZ6q/dsbaBcptBb4dFqeVuz1lOQ8NU
PR863qIOqzpX90a8PSpZXBoquJPcI5Q7ANSXZ9/Vi/+71j/5jRBjx05eaPkH/mcc
T7ZY0u2BVDsxr26nVO42mGy3hNvSHmg5G+FgX1642TZlEGzSuPbJcwkWtX/fhEFf
7oAvnVdhvvR5JWKbtA8FAucgdZvf932Sz+07TskiwUMxfHs/0IKewNuqw0jM6GOu
T7kM51UGvFI4osSwq5zvpMWsmqdKnFRt7oE+XQ7412X+1NqS3E3fe+kWvwHv6O84
oDWzO8NvlkiCMouWZdAO2nPFHEXmnzXTS5oK8k6JYTbfiXGIYhsje4SS6sFgYooc
jiUEr1aDphMFVZivraGPni0IpDzB3JUmQN1JL4baVXT4T4p14F/g7t9wCvsQHKRA
pqKc1SDA24B5rrdamVap5Z0mtyokfidunq86Xoqi9dn8EnReWuYrr99/egI1BRTO
w2//bStIHlF8N+fPDwnil7DRE5CUy2PWtPceALz/xB46/63hZCbY+WEsyVQhqSMO
xDOue7M/d1dpqL4TLbCkARgNW7hsCozajNYQ0tbH/jdBrh/N83rpjqpC9PMMX/61
ml89+eaa0A6lTF60jkWwwETQx94OSk/5ZnX2K9pJBYd3FeBgB1p30065cL1NnrSF
hpMLtitG2djrRJYafG+jXlm05tkol5+vDcQitj2qmf0evlbTtFBs1e3gqc6WWbjo
XQhNeEHwUIOVxdh6VxzHq06v1umcRilb8mP9aNX49cu5Gmk4Tat5Vnne49lTHW8p
bBxlJ2eWXTyT9jSDKTnR34yg/bt98feFz3s0Njsa7/VdsLKo9itD9HkD64gOFirz
zLU+HZoZFVrYXtVBdbbO9B/sACT4vb/7HuhAY2U17Fxx/PKkUa1otinQj/mVHp0T
/HyeTJUNEp95uhdmE7mBtdUdXAFMbrn4J+5efl5MZDGXLRBNgWe+wdb8EL+/KHTb
FPl/5iJ/pxI3tGfLEidH1FqcfTobROIUZduuoWEC0Sfi8IexY4c3VXvdpy1QYd4L
zHwEqGjj+XFVRU4SckgjirPPSXQwSR+FVItIDc5+4NWkaGQeRFqBGro7eawihmIk
Ec4LA74quZNH7XgnO39XwsRCBG0u9O5smS/xk9q2OXDj8W3SJfDAHUGTIORcKnXW
gI/L1jHCFA3bpBFkaRaHzWdSliQPan7rUt5zPITOJWbPaGWRYEPg2ZRwCnTx7m8V
UpF7Bgo6GT1JA/SSEpjL8dV0OWLbU7d0DlJSNkbECurNx9feJzHykgbGKKE6nVTH
0EBIj/al44gNy49ERmSOnuUcs5twrPqO8cpZjzO516Tz4qbqAScMlwxnJjwrscNK
532wU5dl+hzOGBYwvzGrmuPd80Yz6eZA9YC/OB6JIGROdyEObJLIEbDlO0H7LsLf
H4Xe0rhVGTYGTa2bmjntRiC6P1c24hbk0HaivmqEOCyBZ/SDcprc7+CPfojOyd3E
YYcuseirZjt2Da4H3UwP/1BO61vkBVnCUEjMLgG05va9Zl5x8ab4ZD3COmUdCpNc
SU2RhgdSf0c0+wqmL6CJ2e+JMoBesy5I8a3u65xo1iEBoOYjOdmT5gKqiSYNYbtb
xpWWUIxLOXxjEbU9HI3QK44ElqfSjw7sYXMxpLtD64rqSgrOka8VA+zVbbCwGOQi
muNABi0RxhQAnFWWCKZuFiAxj6JLX+yVGKj+n81X8DwFXU/Cdjg3AxoVh0a21gPR
PcEhm1E4YJES+fae+fclXSh+zTWaNyvJ5FYFAxVNa1vjjIhFmwc393nwZGjO0hk5
bYFX4o8r8ySL9J3GJGucG4Dfcxe6Y4iTv4HMlQNa3riGB+ULKs4Lnv97t/o3TpTa
9MgwXzUJsfuQXwpiqDxrbryfz7f9KCAUcJNronqRCoP1pbc/3RVmgYg7u9MwSbge
M/0U34akhssTjiA+HV1l2NdIN4yAXc9m+3xTc15tcGMgIxP+T97+9QUInZAntr5o
mRgrL1hU6jRrhbVxN1Gxxy1cgGxInAYsbnx04aCqcONDL7uAN6jsHpbcCW7cOgpV
BHRYhOslm6gemjO7jyOyIyPYwp1oPCVYLw3zj4rAuYnOWTRtKoK651rHJxa9AF5r
XpQl4hGIMzMqXBZHbFfLfuPizVHJcH2iUvfddUhlILHUhUmylMqP2xx5YBiisNpg
8UVz9jJixPjLVLOx/nOR/iwckMCUiDPBUGTcHix7UWv/8nL9j7dWJpy4CsqUvTb9
gVbvP/d1kSLxv9paKxJM0KEpZPEi2dCk1cFq8gEUTZt+x5BmkEcql7huwToahQQ3
Avp6xyymR641HOS0/sIpD63B2Rt2nQvrIs+qNA1ph28Pb94EUmwcIRBLggNWPZ3n
SVHY3wTOZgvOWLS6wJuITAFmGWthE3KkMPLO2tCzMjKQe1o94agMYqxBbfktqXKt
mA25Ugam19tWPTel57DaIwNKoooYdxZaRBFFGRu+2TY7EZDJ6/qUGDHew16ACrpb
WmCMF6T0QDRAbqirlPio3IvE4I16WCXM1KmqxPBGI7UQrudNLUWXAbB5aWoKd6Ta
0TPBaC668Fv85Jbutzpoknw7Ac9j4YeSj4dT7rst9jc6J4Uosy+YS+h2c/4V2H95
KINOtFw4cPG6zAWyHFd22VUZhMSWkTbEJZkF2Dh1Jz55A3vp1UzsfYYvQZ1GQ5IJ
5zHJgQ3hucKp/neV/inVw+s/KG3s0aSYqsRY5yY0nx7IzT/7fpFaI0Qw37YxFmM4
zAxi2LWxlH/z5P04WDRyG1o5cYQPLo5Iw8dnxzU1G4zJ2cotwLIjsLqoe4YLRHWb
BqHAjTNDhbrK4RAUVO2QO6NHaAeVc3OnrJgdqDMN6Dws2uQzB8fTUVaN6hnvbK5E
gFwjm1dF/q6qvgvUaCIjdcR3Ba3IviolJhU62SRjZUW5whvq7/FU8DJsJuWO+o68
3mvMqYLQZQc0OEdRxAkLOdBJfUKZmObJgd6WzCPgHNQBWLnGtAPJIlzjjRDoYqJo
WJCLrvF5wMBucB2QBM8+5Qxk1jsJbv7K9Wl4jOiQF+YdSzoJZN8I4pI5FjtSlMni
QqZMctmWRRCEdhiQRGsMeko8pM7B2cSnhS6r97/lCeKbAJ7DoPqOlB5IambNHjKe
IUPvJjkFZj1A4urDbMhybbcuwJnn4rzD+aZA/ItZhk4GqpkZaNkdz45XHYzPWVAs
qkH1RvSStv2253qBKUcxt224U0u/zYE5wTSLrQbnOIsa8/kJ0vriGlFYVmV7HMKw
L625lWY66uaqEusWh2wPivbwhkaPR7wg5Dv9R4gmAa4KWFaPkiwgpXGxxmp7p5NT
LcRGncRsuTgvBDZqMsfqlPOqCowejqxddMUuvflkmqzwOjbrepYI4kjsYfWlSO6k
iL3+hRtiLo0JEjcRhwV1hLU4QzNGA6ovWumeAryofKvSIZiQ6MMTs22wxe7ylUBA
FJe365m/CmrL64ZlU0R0RnLTfIAMT3R3fg+MAuHh1eIGn+11duvw8d3vuo8mAYqI
5GcdxKGIpvIw311T/FCUDJKCM4+4v7zTO63w+3movxBbsAfhrbASPNrs0V8OJdE5
XxEi9QpGMJiGhvjlFPGuVD6WfGMjsJdfXR2mLoHCRFTZa6Ay16HM32MYoUd4F1Lo
B50DwcauqlhaNBmi8d/hYdVrrWvC0789tbW8lRaoMgBKXbL6HlVco1J3lbS6U6Ss
UIy13CNYXCke3M0W/vIX3zliQ6LEBONP4aPJOtx2zf+jHEkvb6ZRMBIBrdtkM/4z
8wtuuWCeR/46ABTHXlcsnIFMbY4e8Jms85Q+pRjbk8f6HDkujNXme25SoU/RORlg
8v7wng4yJpPRgNOpNpnHRn5CGIjLid8PJaM3PFZUO6D85GEtIOVFFXULCz7piTbe
IVJkIoInm89N/s6ocR+rG62HxtdChrwqR6UK8nmMyawCfYWyMzur/QgdNLe0UlTe
WPezI90sm7wfDk7g6nUF8sVaCPW9OMxP+M7zLbPx8QbrG7rwURkMBS0WPvBZAYx8
FI/bUzY2AzsIhhRGfjvVjg4afgwaD9PziVOOXvW++RwvYNdB/y8kd73Pji0yhv8j
Dgy9m0NFr5Y5MrBSySZxGIU3nbyzp6OiAt7d+o4wRx/ruyxyU0lPnJJJgV1agFoU
gFyGuqDwiueF8V4H0U31AuG0ei7V5YVVh78zURhBrMeVlKN4SdAxFL9gJ3Sk2X2v
D/BFbGYtQyvmU9OVNN4zx1A4GIqHkpQx7mdF5GVT3xErwx2UjfYIe+CuPQiQIp4G
NgPsgvTFwTFNVAiXqa5O/viGJMuuywDv0O6RieMm37Zwl1V8GNwFPuxC9IayQEve
vebHKDRhzftfjO1IIsv6z3ku+xHvSa/A/R+48AoAUNIkUpBP5Tq6y3n65aLARAdV
lH7lxgMugi5vvkxD78mXqa9fufgBiNd5RkEZH2Dhko6hHcaj9C6K3KwY1f6KTjje
a6/ksslR8PNgTcFwWOkISmXip/8pOtD0S/1P52YjVDK+F55y6x0VcZOBwoc9nQoo
xVqAb2gW0U8gfIaWvFFy1d9XSw+zuBZS/AiZF3xcHSMEisrmK3xEqIQRxBySRoVk
ePlcZCaQQbnIRwnPm7PmOfN68uyFUiPNQVibPDsIa9w4NuTBf6pZD4YJa3R0NzQf
lapO/BnzbjjnR7Ua926rsjE3Kcc9Q1lfQmSkAmr5yl5koPS4I/bJO9bjCHX8LewW
a6hja1UbjMBpBLhwc3SpkQxIjS/esIumq5+tOYui5A7RCauwJHMlw6KugLXj/525
Umufcr3k4tJCnCCuDnb3gsnNBL+YbERzrOQr4k0RQlijVW3nWkvvy4eLqQUfKddP
Q/TGLBfApke1BpqxmvLgTKxW+wSCNtzyv7V5acmE/c7R2tfY20/MS+OBMXsUhwnU
+hL0aJ/JynnPQiMMuAmzYsRk7/D/7c7lhaX2ooG7zy9KEWOzUKqqJF1iR0If/nqh
DNczf451gCHdyj8DCPebJJxvkMUA4EzymLh7N/wTkTfG0LXP0QXSBfyWpTBnn6zT
y/CBtAHAroi4s35ZQNiNttj1vqW0e/vXcfTCCgqE015xCP4qmNzRO4686qmadWcE
xeEbf92rI9n8A7MEgb8Y2uyEaJF/poWpzWqOWJmcYTHtS2WxcCZ64WP77ZrVXKjg
FmygGvjhqWtBnirS5ate2baft/GoYM92/XYLWNVyvgYv6ZFFRpIRd1TMTxOv9eFM
NXCM1dog66U4Ory+EnCaMFQ671ehfQZxVg3Nlea5sOtO6xfeM2dMPuE34NcY3oc8
AJDp5OdtfCZYc4ciq1XwLi4Tgldoc1AgZfhEHFu+XqThjrZrciiEA/s7MJrWwfUO
6JhpeG6I8iUwrT8Nnj6SeU5osZOpuH7mq7yp1WvaD0QrOFKcyR8g8wCuJ2geUvWO
IiscoNEIYH+aHjNPPzOfV/BAVp/OJaBNLK2Nvoraoi5mamVqESvji0qTS0myFAgJ
89LEmhMJSKbullmUfcM1TzsZMNoeFLPCL0Wq6/Ah+Z62lQnzxRiJjtkUgjwJxr37
YkbS7q9ZB6ERlOYm9j1gfbElVYqzgMBHmd41Rs4ym81Rjn8Swdqf1rhQaFBUP6Qa
fUNK+XYflr6nKYgu35S5EFmoxXqA6ozIIowuACtsvJKY/BtdToQjGilxP8a7M6hU
Z5ppreluiT1y+iTg8bZFLXvdXx49BZPSipwS8RV8KmJ1WEjuC9vAYyjev7CV3Z55
yDNjfocz8UJr2GOxBM39ccvrK/CKznQb6XncQPk36JCbLHCI/9vsuhVwv/X5Cn2T
elwIt56y3J+QadwhAOby96fGlcmke4qrbLqD4WTngpfnFGtMTj26m7IW3k9cn26a
HRJqpzd4v+JsDfrlz8yJqtcOpk4o8CaomD8Scis1S1CKlsacqV9dXQsxb/LFmH/X
YzB7jk8NP5wjTy8i47daz8BgmXkJslVY/87fPuYC5RSj1GOErTUIxKuUYlKb7emt
NGT9pcoYdJAaUte1b4kwVz3MrlgEBhmrJsIYcpcXgfrC8YmU3tPhJyqBAGhX4xB7
/pgpz6KVWiJgY807pMxZhm+3gtHEFuWpGIyOQvpR8SDNpTY53YRuD5HTbV1URR8L
9YQcFdph3N1UpiLRGv0WjKvMfjcQYE0wzeUY5kI1YvsU7yhlqfjbQx0Xj+9wb0vC
y1RK8sToaDqpMvZyBZL7BZH2Hmq+paaIxaYPHyVyQPZsVeFcWSDA0JJ84olll9I/
WhWY1VcDmLWmAlwROEifo6tvW9u8voj2YIDD7MYS+iucKeC2CAFesEraB82h3Huq
8dBc9Bt7qlT7Cru1DUmMuEHS5HPjzzVac1kjULrNVu4c4K3uchEFevOheNa1goec
nYJeiGge14uAAkJ+nPKjBZ7IgzuZtxMKT9oy72VSrPfWikKQDEidsZ7VxI256vES
8K3DWi8Va8e30ksKts0wQFMa1Jsi/8/GJ0CdU5d3lAR/dOVoFAksB1Y/zVbgfS64
kBLF1WO4K389CO23s0EPVyN2bgirJk9LjHYc7dPaS6iV/kJp4q6hdlSuvbmPMOW/
nWCRSA09DO5rFIb/91WlhX77rDBDvvt0+fyvv/HLhVRJ7D7H4a9wXzm/ZUEB2vf1
lX7/4gAKfei0gxO3YARd09MkVVrJsQZCsJztwxihlLfSRPN4ExXsP0ZJqOe0xGzT
wwOOZ09SFaVxULp3bsFtKhOlynkrNAVmuzoV4Al+qMC/Vgkdj2b2j0nIyioj+wtK
XovamG4OEoBQOoBVRLA/5BpKuVzukSfj+6MF0x+Ex6XiY9hpq2chXKfjB+rEFgQQ
g5NZqO0/PPlM5HjcNzC1c7mzhWXYR/o4TxyvqNORoSmWGc9arxVo32hxLoeDm15I
7PNqMDHql3yne2AWhcQJ8Qkaeh0ftaCnRAmnRK9NQo4GLqnOu3IgEqbExyisVsDz
8YrDpEHVmSaksfEpdIeP8lJqRVit2vyHByeNuosDRgfhrrXXDYhOZqSvccE7aNDs
jEB/bAJai71LrTWAa5/k/EvUP3yxleW2fysRuAQ460+i2BNriY0+i2Vs42MLSaNd
5kGpb/aoMjCszya2V0ys0NX1i+pggBQZUcQNLH6Tr0MLvybBpIBpsQ9iiywqOY/t
nkdtNcJMa8EoF9GdFYwQGakYlKdb2hPrrPGxJhcs4xKsd1ybD5MEFcrNaePmoM+C
2Ax7sbPumxKChS4RK8HPGdqfxmJZuvi1S6esu6TbvPmemln5/lBBw81su+NQd6Pm
yDD9KxyTkl6fSEXkOzOqcEyULakt5DUsszoPEVU0HZiharYb24xQGEi/OrU2s/8r
xZmX3kdB8uxwJeAq7Nwm4EUEVSbiLKgK0w6WOLBVW1YUax7Iv66ytA5udLDZDPOW
6yB8fAPkC4sr5iTFSwGM1N//olvYhEtvm9XSJ7jUeQKia+r3L6hYX+DCITpLb4oa
ZUiXZECA6Lz3gja1a+vC+Md6hJdBOem8qlowwCtq7KePIjIMxNiXHusR9rwRaI/z
9Pkz92QC6nVXPxJPUdeJFNvArYxfUTxmjKLexMa12kK9bMNu/H0t0i26kZcioE/T
21sN7SpUUMHPjEO0ju9ehxzNWqg0HAbnzFLJASyd6prKBjdVIx7pQd5DyH+kMsrr
WOyurCgyYm+2UU+zwaAe4Nzm0vC67nuLuGOem4DPZTqMCkohiTEJhXaHaMXIKssW
SPuDK6MHF/oqqtMX7uPm063AtvRenXBvAsmFlesgmzvi1bRLFQd5GgELXMMzNY5z
EuYVySg42gO1JZQzKHiWnT2Eg9j3UQmRTstKj4P1EktgumBEm2VSlI49BqISjeaq
kZrvgXm8VGpCdlxy3aYvMKC4IE7qL1wnABvKzGUvh+9ShlqJ3jGKJFUMU2gZBGbK
+UkmSpzUz0qCMwko4mLTEj8Bby3LhnhCilY7B/hN3mFgFpG5XfEy3VWFj+Rz2doW
uKSeJltWz8UwA6qLjih4nTXi7XpTL//l3syYt8z1muhiB2c8tlw6Wv0yX2N3lhEv
eXV6L7OFUWfD2moRq05aAonfXnpvxu/Xj/J2PlisgixffQZZ0FyiSqT6U08aRjwh
zbtIdO7eObN63xStFMr7MsC52CQxvDdJTUFL8Herrsmd4tSGVdlhLvCT18wYDPlz
mIzl3hmuNJT2k0oMKfapFpkQGh+fYV0c8CjZ+kxy2H3X4HdwU2wJHS7HubauGOrl
r8wp4WbF4vVlgoo6DEijUraFY3a3KSqgLI7n6wceHLPePkcwCLy+NmM94ebeTVp9
w6jwUsd4LGx9HJR4BeXn74DqUyAv132uwYcUuihYxuCYweqHF8JhQyC8jXCaFBCx
BJTbqHJW2zP7chMFMF4UC9Jnzu/Za+yMFcfl7d6ysdZDrI/MWv+rKzulZ1Z3PqXV
WhGKtq3ARl8c7J7SZFWeceBYQDXXHmAaY7zH3RP91E0d4YL3MSmm715VSsOzDzLA
6eXQA/NLbadiDyr3g9a/h8DBEWJfDrBTJNT8MBPTUzQATLADIk2YO6fiQqNmidFh
/PXF5rv5ZqgY65FD5ZHi6dzmC4mssUkYh0sD1D7IXn/ru+YVnT/Dr28jL73gqlaQ
unDig5a+LE8b5PWY8Q3nkodjrBNcWSNq9jkjhvbRvrKc+4OAEJAxLkmW2OZHhio1
q/fMuDE3I8RNAhKWGcSui8uvzwHj+aR2FtJWogF7PRb1O2oDfMdX/WGafHsZLxZK
Nyv4hxWI7qmziCN85pA1r0J02zfVQZXfCiiduepGqnTown5M8cXggpyEB3tkZc/1
anakcrnGr1BKzfzvbZFsjwQF4jaZRhqs1e+aL67kSpMovTX5KIYU79zjaEh7KOK3
xIk95vOkK2+Ew26YiQWIRdSIIt4KzbbgtTB6PhRvYID2FPx0hd8IgokgJOjKPATD
OEd3vvOasI7DMl1xOhJ2HrJjJsBo29s5RnFyeU7jNd003TH3V8ZB/wIraKPCcqkc
TwyalpzLyQd1ttnEpX56oBIr/vvPoUU18NwCD+0zAYYRxQ2wI4xFhz46q3i1iBEt
XNEGsPC7uwEBUKJZekLuFPygoqz8SwWicVoIwNYAt4yX7j9ef7+6D2nInL9X5cD0
Ia/UnKNSTu9B9Y93B6SrIQqoHxmhz4EUao6Y/v6IS6M+M5XTvh+GFmBLwEm/mj5N
ygQYg4UhYka75S0H/HO9ZMUJ041MmRHzlypl02yLdbim67XTUb8MtyzuMmEAxvGR
nZ1r5OOQKQtip4P8F3VIZOclmFnCKiG+CcxesbmCw46qQX5nvz3CWH84zaHWkzzf
JhdmKM72LL9zskJJ6UalU8rc+WzclgJ242nZ9VMA7bjUXtcl2kaSPrO9EL4wc+WZ
Yv6Ysqm7kkAvS4G8XsjhcmHPTKUZdlFN6ODz+OZdCdmU8dwFimpuuwwLYTreOHm9
tpxfgIKVg/C2oDQbJHbGpJUqGIIGiSS/Q8BnRYlUKAIFbJcmBZl6DG6/gSQFfVrQ
Yl6R20gAcwJ00KvQBzu0C1q6tN3eg3FnbAa5tnRSCiluqb7aGPR/jUWIG5PkV0hn
9kVSwz9SGvfL8eGs/YCBE6hdC92XwGy1ri7stPuCIStntqaTNRa6LO4GioAO2oJc
sP+okuqxbLPuUCcyAVKa7gpDdbvkJp8GzPPJOac23TlMbYvrwI8z3kgf5bdFG0d0
bH7Ab12OPzV8AYpku0b6m5WJkWC6j4r1WjhX3bSjnxafUGUc55j+AElzCziX71/B
FFBcFsZ/k+bX2lmBnDBGuqjqGdU7+6HvSU+rWrbIN6DCleSAiFLV/uWRCwjBdy0i
KuvholgzVrY8810CsxTTp8FE6W0q1A3fyPOaFRWcyU8RIZUywQwU2xuQC73oXagy
TBC49ZiTOr8UdBMgZ42xsam4OIGLUF5lRyeOLIkg49WzOGzA6gxRhupJ/F6ExyhH
oORmxKrKGplL6l4PPsxBBcQaBGjtHJOFoXKtpdOwPr3JuGcsivxYb5VgP5e+KVjH
mBgg9kKZgXDMeul1R3QdizvT53+0wiy5OFjFlOYQM+r/Fr7O5p+Qt/tV7R8cFvvm
r4VfgP/lq2BF0bTsuF8fNxv1qLU1fR4lp3t/s5NLdpiMJYJNIH5ickXIj4pBicF0
xMhB2qzJhd2BZ/0e3N8ZrVF/RF5bgsojhDM99HJPHIh3tXFItduNGoopU8cvCiZP
lzeCxQByseShZKz9AcOi/cEZZko3K8ykq9Qjc+bsvGFX3S/yEkWjim0ohjnHBnnl
j4ZS/kZGFcN5APGm0EdRc8SLZTcPzyqGysagfE6B0+gUBi1DvcFL1UX2CI05ovkg
YmielTkWYgcD0nCFOJTaixMW/ZjSWCuQMuX7EYgpbvJb1fKLMTuYjAjBoyM5DVOf
owdGYytf47eor218zMgSGCuJ32+Hq2nfnEKiuXodoN8G4X6iiAEtkpde9lWawP31
/gC2ZgRDI4/EBW3E6rmVPySJQIp52VKoNh/Il9hcEV3rzlnjqR4vTREN7jVzFmuJ
qRyqILaEhWCkyF8W4mSak17sMLZQ/v2l8S/fyh2+0v5wQfZRhZ02Ke5OdJtGjJa8
tzyTHKc6l6gD90+QCrsdHLoCNA1IRkge/q398+GD/jxAnzIgDuL9Fll23D8Sq3jM
tIMydX8nonyCE7dY1I166M2I+VsbaNb9VmKLTW+LUXIq6oFb7bi28HHfo6h/Y5YE
53jho40lHhHwcVIsbNwioled5v1DDWhXoTMs7Wyzg43FjYUjcpo7VSlJH/2y/wmu
WQvoj13kWhyjc+Mq0AD6zQGECfKG9f2oKjX7APrXJN4KY3e5dqGPJEaGAr8ztXFw
Ll16BZ3WgrQz1/8PMVcfwAGpbOcdjciW9OPrw0pU0GzrInt6l7415O1KudKoEh3k
LuCulhy11oQ3i8mC0wRW3zVsm7zNGVPsGImzgUllcactTaoYhwm3N14lZ0hu5ghA
IUcyFJms9C2faO9adL4NcuK0RoMpPVmaWz5Si9LnrilWfDGVWV5j0IWSJScyKdVF
iS3+O9zxU7XrSlOGi/CAoWpjJU61jVJTelE38atln7nV3Huu6A/603j1w/JpAFeV
YEtjTJg91LizJG2rQMGLV7uTFNv2AFXX7GEyxzgYSs9nCKPyp37QSOTZ094kZ1R+
feHcyt7jg50mwdsEGU0O4f2jXliYwnUgb2TfyNKXc0ewirpUj+16084lcCEhd0bg
J0rfe0qL18gN0AZoaOtlgTuRuZR8kOb/JdilWdZHUPcvpoV9u3RM4IswwngIg+dS
kgzMzeDR6KmVh5wc0bMRNUdOKncf1kwTEC2tSR8LHvaDQ7DF+bzo5eTn+gjkbn3o
ojocYuIjLnwDjAwjBsvAw8o8zPPQr1lULKZIP7tei7DjAqZA/LfiP9pMd+eh+kgk
Ykf/uXEfbp34vwS/opvgy4QQKTk+vqX6oudJO4zKoPZlyb6dQ/YyNhZeB9b+NeYg
APK2xYxmo+qWHJ8NmSUXrC68CfbrH9vE/zIyWoVIDj3TirTsX/CGIWNW1Uo0hn5K
ZDISLau3Jxw1n2AcbW2i61bWsIFJjaWaYm/Luv0klmku7YztvXH2ivs3SrBwsRp+
W85fr7E2mjWTc1BmqFtlMEIk+U9O+bU+Ai1rNtBBB0cSulVPPv0SVuBtEqzctCkQ
NqpEq/KGq7ab3LsKYjDFIUDCDyASindukRiLAvVooV4eFkdDBCL/076i4K2BCJFq
4wQHjjVHNXc3Ey9HcD8XiUxEvxCeRF2TW8sYiOWJ+ROyNJWKua/+80HAVu2N4AX4
yv4K+aRy7ZleGWBYRm+89RXt2LayZewXpQht87G/vaHhVsSv/SamlXDwYi+hKxtj
kQtR4FGlMCd4DWerTH2yRhVq3G1ISjqnuvcgJ/5WgaaApNsue45yg1wunT1Ee4yR
9HSX1//uczI+LxASA8Ej2fhkQuqwc67TxaVXdGNSBnOMOij05FmER64TmbCNFV/p
rz+ZHxBaS5WZXNgxALkpNmU/lnyp5n0DPdl/de0VmnyE6v7abIAmAjOlIJWB5mNu
yHHoGvOqvJGXJPYwD0qt+oIF5PjYnope/6WZrxxq5t9Bk/mTkIGupKd+WCESU1YA
/dXJD1t7vzvxQtcYA3bXJHAEuKbJ7ehfasTkxj/1lsDHa8Ogmfs9KlBSwlQv83wK
TxUyf7kh2JXZQ+4W85pDN3oE7ZImDVsOMWh49oddNljhs8hBMc223UT9Th1n6lb+
APn3v5FdQzQ0QINriUZ1Fp50ZE9AqluxknDe78X8vLrWGaCcG2ebqGftFdvKxKiO
4uqTG6gWnUxTKBGYA9o8x4ACVt4RoHPyu1UvdQcF0cB9hf8BrLTNFx7f0HsOc0l3
GQVPj5Zd0G49bwx5eB/7IK49riEfzx/wn2GbQGY3SNZjqUIRZdjK7xVdoO370bR4
4HjV12pjtFIioDLJyUnD8mNZEpKpX4JEUVHsR0w7k3cIBfAIN16h929XA3+5TyM8
T+yzGJlr3TTkka27pVNTMBCCskCHAMHRKTwzeKPJPp17QvwjBAul0DGnDk/twrW/
nlKw/i2OvezBrX8xv1XdbSg6QITZ92wuSstN3YedeB0RXLjMBkH/3SXVV/SfcHNn
9VQl1XSlMxjOy1spWpN71nL5ernBAvz43EjPzkxZWaWxoCOI3opgR6XfjR6CmS6b
gdvEncG1iiRLM3EAUziEUlXs/iuWf0MEZH7sQ+opwjoqrQxicAZSc6tkuwEcoCck
xERKHn4A+NcX/RYPxPm8CtUu9sNnU9I7WeJRoOE1hVNn7gVT6DVPZ/rQvK0Zzq3i
G+tUZqMQKK26uSzByNj+UhBp/nNCj0WLnUmjK075vgzmCFOxTL5dvTwrP4sCGKPS
W5EDDSPgfLjmclPUmmEq5cmtv4ti2iBr8EKHRc4E+C+gyWNhJ371Qbv9E0Ds31MH
3sqDMfBv43V9wePZ0CA7bnt/aPLuVIyjU6nbKAvCxLXpTJhC5KzeXdVQlSdbSmZe
+YBq6xmq9aQp47sAFW30TPh1LfFxFSzU/M9V8pJx7f0/1/8jWfvkqh96w1RKpu78
2/gmUVeHBVY++cj33otFAxh+0jSwrI1dB7wwMMh1XTHlHwBn9zmm61uPCvE5dfky
9ZpIf3s2RjyaI5J08tyKHPG5TVPB3NeCS35/KyM3SNG8Dp38skJwnF1Gw4Fnk8BU
GjA1H6BGOYp+9+k+umQLhc0TE986NJblCOW4pAQXL36TvnefnO7YNVPg9QmRJMtX
lcJVmLysoauMr07od8+NrXrDRxe/yQkeGf0mDbmp2fFuxIFJm+Z8a3u9e1D9Kt6S
PnLthPaVAwXnzdsdU9RORTf8pNjPq6CZk51E9d4qerl49GQ8thEIta73cKc90Gq1
dvY9BUXJc22IIjV7af+69FztAV1ljo0+DukeCwW4sywZpIwgAXPu9oCuTa7IuVhU
x0PpwJEIT6TE/zDyMIq5xAGjl527xSuopiiT2NjK7Ck9Eq4ab7dF4WHVTM2Zh3c6
gatXTnqkL2A1gsPr4dTNRt832vojGiLFo1394ricMyUp68tNWwgxww96Sbn2/I50
U8lf/O3aT5MZYbs2RrUvp0ARnzAY7f5+IFJiDu7ws5610wHjzoYSsDz/mgp9qOz7
8J3LkdRZpAs/UE5L6BK/GVqRjYw/ztxFBtyYoYqs00sqWsm6sWnPvEYAKD0FYeVW
Z7IrpwrJo0fvBq3NdRZ/vuxvdvC0jch12rGAL98uHh9wW7CHO6YGnjM+c23lVASy
V50inbRlUwRojGk93AEt7S0nvQboJ/DUpoUjtYJNkdntGUwFHUZIWERdxNfE5rBC
MArOQs3uhwxzJGhY6LdME+yIkO4xsod4ZfEHMz6TtjWD9UEqN91VEB9BNEngJjUy
TUQiLC/DAsUjwSmgeR2JwfrWVa/IJ+3yxOq3WAn7GQP7WA78CSZRhSCw/LV5NvnA
l1jDXYSAhEf2Km1uI1Xwk9tZtX61NdrOdmYp084JPOqtaV6GiB3xlvZor3jrYiDQ
A7xpnY0vcKxECQhYx//ggWslnitJWjXQOCB5Dwn4BHZPVUNugxK/zRmxORtDU84h
k9gyz3siYt1fKJXPa02ojzH+raGOuoREYtYxQhq2ThONGzfxkL6cqvhjvhHiUsHP
ayOngf/QLUiOPtXk9nYrdQWObM1EzmE/glKCmxQXFhQ/zPf7JEDDvHvNdGEIU3gF
8Xe6n+IDYB7MZa5JZQkJXMTj6H/+UuAU7qbpj6Wx1Op5BHmJuMjdygtzxqTEIJ/t
pVRoS4vYI9PhS+l2QG31o8waEGIqBK7LTZeCcRtHVuLv6ZFtOe1MMQZpk1Amss8N
xnIx/vKmMJ1QzRstyfiGzvXfeDwAoHU896C0rkyU1qOf1qxSeTuxX/ZGO3HctQ8D
zjrDdrIcPyy5ryCawV8sy2y/oGw5N6qUP0XjYhBxSY6uG6J5jVlHQq6GQLxxP2IR
AKZx2hCaFCOmOF5dKUVRqeqGrLgauKT3HF59h5WcNzHEfWtF9mZ3ah6yWPBIGIXn
WqcLWTaLfR2zGUGdED7p+a2bm1eWD9xggOkU3y0RDhEtWC/gbn20F7PDzNuCWx47
OSBQeT72LET2jLXXiRNcOk4FHYuAVPAhf6A8VqulQk3yCIHKG1gXItmV2xD3+PY6
/ydIVgt3ldkw+4gfXq9iQALrQZAlIXbaFCzMK4KZEF6b4Mdz7I57Ly3M2VKnpfQD
Gk2O/82HYQiWBOCwSTAT+JjqH4Beh4ctgenpEbVL+rHkN5lWWMCU3fCUVvoq5gh4
wcNOA/ToolxXhWINKhZSdgyMeX2OyKH/pudfJS8OSHawXQPya86+H2yFdJB1i3Vj
wcMlFRrv+93ij1okKvPkwYCZTugejK8EEtpXHozxtXpLKAprAw1Dzjb4we8GEZtk
/NjXzxeUSCMSKhvt7KkinBYZhkOGbDwqgWcc2eDVddXG2BxMBGtzksy1P5WzgOyL
65TE1UodIZRB1Tc9mdLB5CokN4BUkIj7wnHSYxzVrqIofQ2HnU1MbfFa+B5hGemK
HgQUipnfhGFmFk7oDc8nugXZbZg3dT/VLSZXBMPkGgTjAHdun7T9oqoSvJx/DrNT
X9XoXTCSoD5hm/UUHtOtqoHPtkokGGs2S7R+mRPUuF6M+HkwyEVAZ0RZRTWg8xep
UlZzKZ/KWHKx9G7cLL0008z7IiE72cegbHRbeFwprgGLAr4nNq1OaH9J8YH9N0Sy
ad6kCB2SoBKuDdnyruVeAP5zL0FejQbOyT9Ours88Dtv+wZogdkiqaY45LxJCcTz
Z3yfePd1r8SSBQuIA1i4eRbMCpsrybIhjOXA6GQri46P1Y9n2/zvS/qGgp+PnkVn
rYmQ+XsOcSP/FH0U4ruw+MrC98jAfXqpe4eghxhuz0ThJMhrUT4I3Y3e2MK/vfh1
VPOBtLguBIp+MeJsG8ktoooM1v86Sg54a44LUmjglAgYJHBWr1AfFU7x2pITpukQ
9DNfwyEz6fd8NDBFiJmLDq7REV0xiOKWamWE/lljTpl74T/qTKtF4ozMYRyqpEFB
2VJbDOEPv7URaBt902v9+Y9KiwahxxE9qDrxnWptbPXbgkhwLGalv2anrDgNciwH
3anVx3xZxHyKw8oPsNGgQoI1YmjbpspvdjXKAn9Ss7ZZmhg8o4XYADaDFHFhfLho
K9aZvX2klrdwxnKpXxQ2IilpDZ33P+qo4wQSG78UbiEZPl90fms2xBPpA6X4ERU3
DB+AqwGir32OzvZjNyjIFCZ+bpM91yu+t4NPCPz9MnqreZaeVf7AbgVVjifqkyC+
SF6BbjaFxv8tVlcKxARMIoULVs7lqmtNbdUNsxXz+FjeHRN3ILxYLl2TFkfjAC1V
2TXPsOigLJ+dHcA0MuW2S1tbpCI4pmf7goHsu3wa99gSR7vHxkZMJci41IEsSsXY
f7ZJ/1ANohFndE4gpj+7SH+AmvfruoCfjZqd+X/+p4IybHxpDRsmVcFtq5s9uJg2
mR/f8UsJEMv0OGCmvKINBLYPjXdJ0CnmDzoX0YdM6qjHxy7ISzkZ3IHYCaq+AuGN
Gu0phO0bDuZO4bDYOBdze6XYCRfxp5NyP1ub4Hpbnbuhb3CKOm9HwrGCvqnDeBtt
Df7HBPLmuVPgjitByThwE4jOX5ByghkB0q/0EGgCfe4pKZcTeV+a5gsPFjaablOk
UvwbomdGKJ7exOPJhkGcFiXxO1PHKupuUtUB5FRYQ8e+f7Y495zpiSBkcFwtvjOL
9R3iVzS3JfTu1hdyVNmSvC61DCAhpkti4pSIzBKB8PzaGF3gpVCYBRRr1hvDfGR/
O+UMmF5/D6+S2V2q1EUlQlFNZkwTVBQEFKB7WCASfkCDOjZEBagvCfo28f6Zor7q
t84KsP7rNYXt6PKozBQPJF1s5/UnxYp7Nlfn7C4OFsQ6rdgb9nW+HlrBoDHohYLB
oBtQ5d2fl70IlG9HCwzh75b22keDWC8+AwR+Kmct/SK79VScEUdnG1hhy9nJpp7a
ls0h6JlAwm6SVYJVnN2c1ayVvwEf0omNJ9WU5Ef47onpMwC72/nFfdPMoMS7aREt
HpVV2swPd8dxj9CnI62fwNBNXo0ZxN92LLXF+zZQ1tz8ugZHObn19hGJYHwbrzwI
LBMKgCrh4J4NHKKrrWPi3GGgZoRIcz9evGVT2/qexMCLbB31sxuPUTSjI9jbrZdg
HsjDfrfxLKvVoU8FUBzkvKQL3HJ/vlZoICmf0VkAG0Z/nPh1wT26rFbB7Pzk5Xkm
fNrt52a7YXAzZQZS2k/UZS4m5pk680TyKmi8FmREL/HHnK0X+ws9uKXSWGi4Qqpe
DvoGCm6b/VfYOCJSQVlbPGCDCbpj/J9d1izBNSQb89GRlWutVYbmD+opnJlNKOq2
OliFVQ8uLF8Tp2+18YwwqpesnWStkCUvVipGgaz0uJpRptCBqCB3c96Evcrx2Vt6
eYzWAxQpK1vbeC0wszej1Y6sX9jbUI1HbCq866ZrZ0qi3pe0NO/7e64qWrEHAwMU
1u0JPUSCrB3wEsUsASmu0aPzDK1X7wSoodekgS+W8VysgfnKugMcN1Ba+UkdAMax
f2cmdXj4LACg/vAdjOa9V1gNwYwvhSPzBfLOmWO4UTaxd5XtzTNJvt4YeGkxyZjv
4XAV+SVcM+cc1o1OFusO4lSMxGXOwlBXVhVCgUGw8FuI3zn9YeqFh76UgsFMg+Nh
u5ryLEQ0u7Mc3VvuMH4x4YNZXGtRPsLRtxws/ztDpb0gXk1OIFKQMcZolNsscfg1
AEkR9TGvV3V0skDYRRTYDYYGWB1Mpig4IEZknkXBnbdH6dGUJv1L4I4/r53P6JZ5
AGGzkyPHL1dwN0ZefLOGjZrc0USa2cWhBGdd/5QcJpeDkMVqehPNwZshUEYiBe+Y
jY8LpLbLWSk8xSvFeYZb3OrYZk5EnV45YWgHVPFwWz+bWzmuZfEbohhAB7Bbyhr9
B+DoB2AC3nooFu6iRUkJ+Jp2kbjrMlZJTM0Rc5duiGLk1H77OolHUZMvuFyJ68oq
FfVDZghXepxXwUb3oNSzGY1TdQjQ4ze+BXbA0yWmSib4eP6oqcOjwnt5CD6KBZ3N
VWOp6NuLzv/2NzLbQBJjbRRr2KAUYDTYNcFo9AJok9xPKAziw4fXJuetTevkIIMF
JZr5t0GSIbUpNXUprMQBxZKfayJV66+SM8i2s8Evhivsq51QLeA8l6QpXUyW3zN/
6BCP7lLgpC0eSnss9jFrjcTILShB9XRVSfZtkzZYNN6FVvTgIpOhZ1qzAWmbDC0G
e4H3wVmfCkLYrJ1XihVg23cCInzcPo8ZrEq+l/E46/bs0DBZvRkT1bkiASW0joqD
yYMvjdploXajXs5O2kiXOgJ3O+xCifgetC1Gpb/59fLq/xmAmwCPQRKlN+7oevoq
HyvY6MYV0n04+0RPU5QIHbX/0jYUUQGdVFX1FWDSJfSvSqkJ6fu/rfGWoNGxEWjr
b2NfWkWCOmctkU/itQNe0xZtYrtxBBfBuDYgGwxWQHUdcAUjpxoz6xS7lsrxnpNg
dhf74XnPSM5xcVnusbWCSp/t0nI5Nq+NovR0D6tmsHKsgp4jO8jOFM4P/Z+jfh5G
XozgDnQ/9evbQ/Cc8SPlr1ucZXXaS+BbgeMwXTkyYkmgEoPeU5koO5/R8XWl9Hvs
tEaIS1hCuqO3ivTQZOGDsmWSHrJRA8zlHeywVQrt8BElzKcofkXNra2SAOeGkiVz
oIyG88Z1c4kgPA1sHCp3pNzbF3y2gAJVRwvh4kPkCBojVEAtAaswYvKSXeBo5cSz
CVsZ9VxH8bkT62jRrwsBWXvbuXRMQV+5lhkVC+MV2IQ308q5p1jBbSJtIxWXLBRR
JTj5tS8wR9WkuzCea+qPns3XHxic0fGiJ4RwQLwOYVQIaV3h2c//mzmRcXG5fbVM
5GMtQyugSRZze7P1EAOndFgOynAHtTunC+BXeRZw6PrzY0CPMyXSiWJXWjCm59Ll
D8C0RxlgGzbJwoBraqDmbOTgOVPp9G36m1bAvE621CCE5g8nudn0qJQ99/6XcLgH
cbsIZ9g/9B9nXIIlu7l1tiTy7UaXVV++Ziyx3J4Q4vvOUhl005BAjkQATXaaQ87A
MEdLDbbfRLXBZo/iI87jU1ZuBx9zHNu99v8JQ/IgNtGzgMQU6K26qbHj3PdLeg+Z
8ZJoNZcrFLlO7fclN7OjG6J9gB3w33zudo3BrLYf93Tl2nl/grhLNsiEpr6WQFTm
v0fTKkWNTZ1AEsCpZsz/QMfiowqIvyRMtOAAzzQzHHeTb2vgl5eJ7uw1XwM2LRHQ
u77VXdaNCUZSDN3Kyvjh3MrPUXB5J8WYGH9toHCw3HgTKSEq3Z6Z52c65vTETf9o
EIUeamN77iSe0zzTV8QJx26lkCdqFtHuv26VRNbfkz7C3xkIzstW+I+00jKa2hYa
Zx8L4QFN/8BPooG9nLRnPUfhzCSFeqkTrmL8b3+aly/fsmYCvS3mLoivduik/bcp
DUsDWBiLSZnTcReeiuJb+Nx5U4+DwBROunEmNxpnPGYGiugDakmzzX1tbW8waGjw
RIWdwyEBHm0Kl8H4I9Q5D/VsvVvYue6ySHcUfwMBlRZjkG/UVgPMp4BQL7kNi2w9
SdiEpBnByGxHLfQHK1DPi+0m0fRyUPhkb/XLsxT1+yavgtPjKNE8DTYdW6vf0F+C
riebI5ZMw+7cg9aX3GWDXTyHm9SghoUcFDEa59Mbl1P7nr53i0HxxoxOZ5Pe44ql
nG/DH2njRN5IL2jyhhYXVYZF2jy8KQdNALxVRvNEPEk9bNT5rAQ8x+a/nxg0eG4b
+MjYZaHo7xNQXbqsPyvY+/sO1AUXJJKzHS5gy3LPQ6Ls9gnqxKBNhR2BUbxozqQo
ymu3fHwXNoH+TWpri0Ydv5eogqsyhiDbEfHHgbDUXiPtsDxFW3z0xqbWLUqU7k/8
/E6WLIO5pvGYNu9Fi8HL+I2fUONgskzPN9xmNRJ5UvpjALBA88eUCd70nTIyUxQT
7KSWQPVHEFlm1KXio7t4n5MfDN5gUBtw96Bcp0r4rNUdRn6fsLUu+uv5co5VS4LK
ld3I8UnYfD9yYQ3X6zzmjUdjlRzxnsZk8NHHdh8irKtcRFenfT1VLTepEXz+jI1i
oT/W/w1d5QLB7jIVIOBGYk8sCTTq4YBD/qqn2Ffsyy6XdGDoKjhsbdhBV3rq4g7r
3XU6rnnmVvogJL4HBB11D/XWv4z9340LNki1YOOmlEW3C5dy6AlrPhCuBXRonHOe
tPZYinV3XET9qNRtNKuN4Kt3XgM/5I4q3V4IhiiB07DQq/zCZJ8cdzkHvFULO/NC
QEYmtbdZBtbf1Wk1KynnbEUQGesxXhZ0n6r0SUuyrORjZFTJXsrj5hoRc9uIjWw3
alH1FvCEBtzuGStzB4jf/1XUPezUg342I60U2o6zrPpVFAAEduAKKttf5/CkK27H
+E7Td/gOYg/UM1AtNWriPISP3HetjujCMg4e/PaWG6ELGlubV+Vdd4KQX7FDyezX
axAt0Cs3ly+ocpRCRmJ/cMxU9rREzejY5GsKhgujRk4l44oPzXKUQ5pbCQ3B2aUh
PksoxprPNnVjD5791S9cMlUpk1H9qJFDrEbtvZHztHYLxZ0OYVYIJRzE1f20wuUI
PxlLAuNIU3MucFArYaxKAzzb2uVhjzXNZGuohFJ/JOq4Az5j2FcQAw8Hfj2iW/2l
xdyCo4S1R+NjvW6ir56Z3XK7eGL3O9sh9nNT7dfGhvanNtrXIXUQ0zsWuVsmG3Qx
5goCtKUBiuo0CmiEA+I981udQkjqR5IJTpYPSxqm1kzI4tKyCrw3sVm/9ol0p4V0
8WM1yVjLg5N0C71lA8xap7l5kWnNZT3a0cmxFnMsa76yqRgCOz0NdaXoCx6YhcXV
ZeviZvOjstoitY5YjBsjAS6zYKR2skobWdLkpVX0DVFyniy5xrqlI0t1JrhiShxn
zL0yJzPSLPyVLIIN/ZysPJY65+0zdJnLOG39NF9g1luJOaw3CTVvXgTjrtpYQqHX
4+NahO1GQZoQ6rN8Rg65YSa7p3Pv75QcxQLIn1237O5cZ++6thNvhGjJ0zwSEnPA
e/j3SCzf/4n60dnyfOmcK/cSpMeOud6J2X6YGUzK+2sCnAZtAAw4OyUaN4bMyycA
tM8yzCr115K93rVjTK6GadgHt5sIvdWNBLD8PxgJnUCXrqBQKsL6AUKTdiYjIzqe
LHGpkpQQB2AXmmE8IitPVsRllEfNvZlMBpCRNzXXn1BWkSjJmmd1yp6vc6mC9U5f
TG2COETiIVCirpm313v6iyjNDPGelRHmKOzOsv++8Zai71GPaGd9VMCY+Q9qddZS
tbkd3cuKKPfBgStK8ep2dBJoknJLe1j0vHaG4LvJaXl4VEQLptj8DRxAQt5a+Lt/
qzF1lYY5azS9IEIOVsjxXC6XlGUSbDU3bnfykx4l8rXgy0hAtleCWbGHGvPLVL0H
cTtXuAJ8jViE5rEcbaRhfa8FEQ3ydAEarfJVyTNl6BOUxPFmKzCAr+5MRcRk6KFM
OxAr+ooBO9rPoDLgFD+3lmx2AOHiO8Lp2Mtiundd8DF3uS10gihVlabAePtBgYDO
Ta37EO6gRjG5BsVnpsJMf3yYDfSi81K8D27jA8hCeiVNpcVGERsgK1bn+6TskwoQ
St4GUlKfHjpscJx9dHgUHcKxKN2L//f9rEvIHhKvbo7CJg+vssWBrjfJNq10/ekK
qE3ySGv3Kl2ktKf5CpHTgd/jUKVo+jjdxyQqs/ZRKRuEmQKXtWc0CYQqZ6cvkBOH
F0fA6oPUU9bEkKvqMDVlijpRgEd0M3Gsu7+bkRqbCvtAvwvfbiTC+pgOp++hKgwk
/HJKmEzCeVWBvk3VYxdRsAjNCJHne6RiBSijb8id/SALDIrpXWp5QN9tdrskUeo2
mbuUivE/vnXBsW1y2+4jMMsoarFDZCP7qneX4pMAsctIn3mMSy4pOLVU9R16C7rt
m2FIUBJVyWfLjztgyBuq9MGUVdwtkJ/bz1uvsxnPLe7Z10HDem5ouEdw+1yhFzWc
cOlevO2g7x8Jg7j/zERXha/g2CYRliQbqEw9js4oOc22QzzsIjg5/zUe/qsVlFgD
NhoedCZ5L+aapnfAhj1Xj4+ZQYsmdE7NSEw0pTYsy1SApW6AFEmcAf9AMpvxSPE+
1ptlJbtWGpeZEw3Ax1HWdqDAjLEwkEb7ON8H31Gyi5CAB0+hx5jXZ4JdpDfjn/7L
1q4ZFnr9qB5pc62O7ZmYimOpmm/3zcdKi91KnSB8mLQun23YMgQTntexr1SxPoDg
zcjCD9Xl3uATYpLeNbKu7px375+O6kgkORM8pG2FraNZBhHaqWA3hzKZ8dFjE1U/
O4RWNAROwnw0zcDNJuTdH6larCxDZUHKDI/D6JGwMkzduGzt1SyUjjt5fh19AvPh
VwQKXG34A2UsTd+IzCY45OBLtIJuVOTA6qDkOkCplKCUqe/P1dPqZR6ZmgE6OLfG
u9lxHDC3iK37H6hrJICnjWwPqv3fB+A3FnwlVew0yd18550B+5amCABKt1+N3GV3
oulUHalPVA9TSxxREPhpS36m1GygPAV08zZpd+BOzHnmJwSiF/9UBA04BKt7ltVL
deO+ejG8QCO9O5Ptb0wTwNrFWXGnlUEAiTrbzgyfNMIZEmbRRNt9aJini9+Hdt0E
NzaF1Tzd/HMmOut6IKhy7Vz0Ex/OQFs3oqpeCSd+aqCST1O3hDZyIo7BZqO5+uFo
A6F1Ay0bp3uq4totBewY9FYdw8t5VZhE+8V6o7HbFz9vSQ2/v13sjwbGwkrEJbJs
RRP6soGvCzmpntV5oVsmVqt/DV2w2bcHsDwSJDVgOhL7SNE+z4ltmeATS2b2EOHQ
iGKnQIPg0VwdEaUtWdGYbpx9kLcJmCQeMdM3fHX6cJtLA46WqwIjGz72GllHGwn+
xaMJKPZdHTD9+DOGxD364i6CZ+UewqRV3FURWeqNo86ZNdTf9/hscTo6HwOtZOsw
329QmXV7GimuY1KLrGhECkExgb1OvlI8qWBw95REEEtDN1zpgho54VGFoOK4cXIM
6TRjPj3vUbkaqL8BzHwW8iSYzQ28Ep5XwkUDVMK/r+TLVEnDBlHPVdXcawUqi+jV
uS3KeLUwCmQpY/jeVjXMYooz6Usjp7PhPY/bncX+CYOstTdFLtModR0ff7d9sJLf
dqvWCA9xb+aeogWhagW4/QRlvyVEkOPPPRZyKH8P3ShJZTgc426PYTnLPZv5krIo
mnViw2WNMyjgxd8R/hw++f02wpk2rwqOjKojOqXgKTDQyIKPeP3YuB4+l7vh+cpW
OWpfMG6M9Sy3gtQlphyueqXS5cHTRh42LEdjQw67EENppWSjT7iCxdbKvd3H/Zc7
9gm1QCwEhJw1w+VcaPLby+GDQaHs45LLSs9sTbRrzg6Y2xIr2/i5Ngp7aa58CreB
XAcRzWrk8F13mrxBMnY2VFFxTBnTc87rQI1I7jU0cwyXu+WSqywnSsU1jG+FVk4i
onJZNWo9K0PZCZc5fJlQiHn/zK7BOoV71MIiw1kTtHM3bnfJd0pmD4i1Eq8X/Udj
WZeXlo3IhVKo++r+xUvtjuwMC//LUcOD4gaFY4dfqmP6gfAe2IXlDVfDU/Z5y9xI
fPV8SI2p8DhfYyuxDv6V2JyUuebTHP707Ch2zmplYRHDADnVknTFjf2EGjBO2VTJ
78rMZhFM+e3jBFqB89uG9qvbYj35V03kErS+AoCGRXvV0mSA7jkudiWqr3JvVKym
FBocusy91Te3AffyTm75XOCO9AdSDKjURnd++iu33cuRlzFmkotQfnRFaoblQYG+
+fMKutyhHudPM0B+snc/RAARujarRG3/uh+48GyvjUBtmvxkK97HFdKz3s7lvPRY
QIiw87YEsrzyr2qGIh1PBOuzDS/Uu0NHtK/r/7f5l+Te7EuomMUxxjFXtRFhXtb7
CrjcpQwfMltYOiQrKtghuSd9p/cm/RKtZvh7TXj8dJFPKYe9sLugxBpj8iTess/+
ENsJJYdzN2cJVCku7sUPRepQbf36p0mTw14VRK+pwZEskUhxf++2Rt8CWvJc+C44
1u9pCGcmUD/SZPPbV8w5sy3mrQeIG47hZrO3dA5ojPr81MJQLC2XKvOeM/ueCGoS
CmKyKTYvZ+Uwls2JjIR/ZLoArEONLmuuSpacwFh0vIpb84iAoKm6P//4jtx0y7x4
/Y37EGcOpbYGC7uZ8qJWznT5MlmPBCR/LVoScg65IU0EvTPm2z6vTdGUjI8QekkQ
QFTfrHPa1HMTZ68vpd8nfqBqO7Mosyam0N6H4VijLAQ5e5OlMsV8damThd+k9F4M
H7SfAl/IECJKdYm0EBCWU0AjBy5bkFe0qW5SeRbzfxKN3zxCuzOdDytzegeV4AxO
mAkbKUIEcWkSetdAAPD5bZ5g/pdtAaQU3kZu831HQ7aELhfKClj0S8X+fQVqLFzq
bFcgfVCNgkGaND7EhAchsXdrv1vBKYYxMSEljo4S1X9SSptGid2Z5ZKmjIpkS3BB
/JTqVwIHexJKPHVdGIL9t2InBjHwkRcMnfoirbtyN0gPYrFABy1iUrsR10i08/h8
5jCso1Uj9ZG2A8uIbHZMDRqelTsRFzi+zpDWPYG1rU/MY21Uxt1tX3mL5XLYgN1J
m47+SDaMubonRiDNNVrayu3NC6tJdxvnNuSzSKhFlAWxZwwMRcFdo9aqmtDDE2NT
ka0cZDOFMo5pqa/3DoeTrfDAzNkX1lzwlUROD0GdHoalbYQ8hx2kbuF4TrhJDMqK
kG2k7KoVI0OafCIi3cJKhjeGcT/ik8YStcW/ubKqvDKFx8y4cdds5jTDXJ3nVrxt
avJ1Tzqk5omOrGL1d/m4ico+NyH6kqb600mwzE4C6zO9VC8NrNDjw7o3ji/cxImu
9EI53cI9T2RnMBWy6KfUCozhT66jPshd1GGI458YizlChArBv1zerKxKLzGdIj7U
xuZipewzrSB39Mc3R7cOy0f51UEufceAVl9lgTIIEZj+cJUBVT2C39ZXuUBa/nld
qlJ/x6lzuQHAu2YsoJVbZ9e57+7L7TJ5uBR/6DFjYHMXj6fK3fBNHw3XoaK18kIY
coUYnZ5mre2+apowq41f3zUx47IyvkY2mRPcKS5WoKwtMYcvs8DhwZRK8u1obRYO
F4tYGVhcqEjL+dLQbkVzQJ3s4yR/kR/s/+thvPXPQBAaxOF0JOJs0VoTCDpT4HuX
7jlgclVRzduoCCGzJlbxxZ+/1sCymzPV7H5ucP/x3kECaTZkhQ8t7Ptpub5yU3Zo
ubHlhCE/Z2wVO7mWVduBXrhQ8XiFVnX9B8kou5l9eNPr7+Z/vd/iP64I+xywRWIy
kxnyfDXPWYes4o98g3iUa3Q+fbvFudlWu3Y3mJF/xB5apC1pAhrB/xwEWq62dP0m
pqUnMbwcMDrCgiTqerIs72GoA25k6JyFBdKYMAkpz6p0NJsA1RJI34Up5wfiIWkJ
yjTyUi3bnBHKs+SDFtv2dKU62dALbkkLxGO9cgB1yRREeJB1qJLyyM24GkLHtu72
brJD1FdjdCwjkOjAGVdQYA0aRP1iAJMeFlTdXYQ/R4ov8P3GaJNIxh26g1LN5T7v
kF2EcSMiyl/mypeQkdr3nBiOqyiZiovPqwwH4aY5PuPzb7cKKrJ7AvNHfzjexbl9
JJX6XifFGFl4AIT0BB6FeLfQFiKMGRMCAZ23divWbWA5zm2smbwbZh/98pSgSGzm
Rai7V4v5WR+D1ojHWMSqAriEfrfSGruClT2Qp5GO2oDhzM4vyB+o9rkdOZ8AbIrm
hTOUBinPAJL22VvsHL3Jto/Kl/kxjZyRheg0zsqYFl1MoDykcEqzm1yAf9XMva2z
FZKTbQsWYDHHUc+aqFKL1xIFX4sNialjn2VMCQVq9Mo3XCTuCqs5pNQ8M3gr7fjT
guBlWzwCyFyW5lTZ6JyvYkut4J32oK/RD6V1gFSQdiQycRPzd3ol1WpHKDbYBiSc
aNujnNRg+eRNwoD8CTrVAmsTucL9KtyQ6B3MFx1KzSX/7nQS1qZL+/gpY6yNdM6A
5L/3g5Dfj0mSJv2Fsen2aRQzZFKtid7W3o15dUlRFUmGPl6f8vkbRqcKw3pyMxvD
+I0IGclRnJHGfnW6POSa1gUzSyf7y14xgXC13AfaleT5cm77aeLIgxT5B68fpPMm
OPxcRHyOm7xaJWX0f/alDyFq96tZg/x7wgRHjTPhAhUWt8lctKIYgoyh8qNk4zu6
mMV09D93+R+6a+1JEyzBubHllKag+U7TErUjQ5Ea1f9Yp5WOwrUrcLj3T7UHdb4o
0ar5LB1Fgkrn5qM7ZrV+Xgpws/+cMKSZPjuWOVSbYk23gcgarmjIgHhWflQDnPq4
IwZYH32Xy0xMfN+wfzHo70Q8KfdGkzlXFKxi1ANGP0u6GB4RqwoEbrYEj8vWye0X
Ek66f95RSoE49cDHiq62NbVtcov/4ZfW0yG12qYNUHpOjkgg98ZQ37SZaqW25Wvo
IX0TZgXmfUDr9K978kLKh7fuDZD64hCm1FpP1+z7NDLCLCMb9zP4v4eY6Z2ATLeK
M8MSBmJfpSOQClRpQ7Zm1FAgdgD+9TxbcrmmnhlWGAX/PLylwMsxDZX7Zvq7bKtq
eihFTOayrjFfIxV2skfAqoiz160jgg6ggtKIuxXEsxmF/TfS+t2Hl9M4wNI+CLfr
pzQdueMTsVI5mT8gdrramuQV5uV62Gmp0gYvhRnxZNGYLl2ZPTmJBqkbntBGV7eC
rNltZ4O24SqKRpB5wZoEkb4NJ2IHVnaR4fxHPaSoHLY0+OLrnq9QxIxXhwPDKj99
ebqDJpW2ZZwhyiIuqJbzVEvt3HV7b99SFShNGUSnPC6vxycOCXlROZlX5l8w141K
q4Y0Kjr6va3qU34uSIdy84Qa6YbmGTze/RJPENzaRsx/fW4yq38wa/Xkx9FYcwK9
Z46nh/U4EZibrutoIz43B93oYZuS+1QP91GpQKJR8HPBOh5JVFeUsB+4qWD3igCH
5xa3N11w0Lpzk+5d9NwIc9/a83QkUKGnTou/GHEOwr8jDJXrKm8+fLolZuWjPSRG
t2zGzXzOoH8xvfEfmFwu75ty76+ACNTBBCWx0UXEZcFLvwLrTpdDAkgvHsiqZR8C
l+pnDMBQK6EQY9tirSsMHUmmqKIEm90FUAwyDc9eXrOG7SVojMI+/ZvYZF49yMJu
D1/1RgvMN8MPP9+6fujIY9DjMppaFhxz/euocdv/Jh6k0iGLc9IxwkiEGIfmNoWp
bJN47JPvrfUnMAUqsHF0MUDwufM1Jrv/1xQfRfji6UZSwARh45gtczttW3SosDDP
EyUk1HBfm+8TvLol2nSnOothFVx0Rk5E1IXOeIugbW3yDAExki7lP5ZUt5uK/HK6
K9Wf2BhaQWVcErnjo5HZjM1s20sTONvgLvNtDG1LGtOhWmYnjsX9Tz832Mv3JzfZ
OXny0cqjhWMkk3Qc8xBkkSTJItvbPYLrU2rlUUzYxJ3UrybgxeW8XlAyjIdnNsFK
Nd6V+iqepMXGc/Ekyxw+i7KH8uKu4yQtddKjVWH1cOI0Gni4tvCvncWaPfC7Jxd6
awgVPNB1m+HpEabtkAzmJHp0DfmCYeUmMojRo0HjWynz0WVsv6R69Osh1L4LUo08
CnYBzk93lwYYZ/OY9cLc38CP2lg6noV4D+2/lIzUQpk0fYKpVibvjUH1bmkFIOEx
+Bsl6jEw+SNT5TDBnnZ8gYrYzeLoRZ2ILYC3gOeIi4F8mkQAEBsFHonNbL8JnFGL
7FQRQyXCTz/TV6T1XtihyyEIwJzfZkRGu4DnYtNTH6cgk6+DCz9W1gMwxRAGllJl
kK4hLUrGvmgYeJaAPCLXyB5dL5uGbykBtkIwdXMGF5LJPLjMUO7GUcZdtMgz1P7S
hxGzKZtypthIqZ2Cf+ZdUivVl6HdWIKFUQgO7Jym/1z8lwUAIK9ln5PR00xZpzi0
tc7WHhMnteN/npEtnot4D8f4+4GtDDCMvPkyU56OcbU3f+KO3O/oX0s4Xj/64c+A
3GqBk8/uTWCGcup/hwuln2P8Wi7VCKLjLH3a2cNxD0bFRWR221RIXIywUSL2DnPl
We9cVG04/eFe0IBl7ZiWR5kmHqpM/cXQVQMP147GX6UpC8Z1pp22e4/xzuDgHHHI
AKFhtQI++vy6irlzD0vRECinJCMNWAy5At59CDsOUKdtBHIh5nUKZ53/g+3cfHtN
krOoZF50hhXavE38V4cTkeC2xHVTSYuN3MjtJGESHDJsdR9/hLgPJiqwGDO9OEqS
WQjuFMIqhYKza/8hfChPcg40Ptf+47uQ2X4WCDsdETyE5pJ4oFel6NbZSSSimibC
1ucYzpnk+V8DBxmoP7uKzQf3317bN25NBYkvhXBSt7mnhKet9ZsYhbTLns1mdl0N
rOd605OhjDh6vIioR8WEnelqb8gtyGsmF1KTmwhdpftE45din1AxPdiIeNaNJ9su
v5z8polFvsa2aPE6p22L02m+kgDKqfvbpAnFhnZRbl5pdPvHzwbtsIP7eF0103Yc
znNgvTXwKRgxU1H8a94t5+StQXgSgcebWpq2kkLgEEdQGfwo9lwgP9DeFCv/MBIx
8TrLM4AuREFYE9GF0WPBYN1JQjhqeQIjSDw9t6D0VBcT21Mchc5Tl1LXv1PsMAdx
vD/KBVv9Yi4fZUFOyEMIWg2IYoCb99+Mi823bsezXgtFMqMSOaNj7Psg+sY3kTA7
yEifrm/O/8ZbO2pDjgQ/NiTx9BHF6Opbex4V9pgubp26HEF+3B57GZpxOgKeP+n/
TtBwLaOrw+XGopWm42XUIGZiUJx+OSbfCr3TDQfrM5jYj8Gmli4rDLs4gXsZuOlC
ryTU8ZvmC2QnRGanIvYyG7NbAjLyWO9+rqIr2+36JhYRQ0WyfmjcJH92Q/dpCv7N
+DZA8VQmqRadAQhGbyxG1Ma6nXN9dpnDmAveInqFOqa9cg9EfCgbwM9o4pcL1dwk
z8guYHWaf3Tq7OqMnoJKupP7QE2z9BT68B0ee//ebbZU48+A5N012YoMfmbpsXGL
W2/QaR98tY49ZNp4IQFAykYwcE+3b7UPXkc5ZFbDUJPOzRMjedVR7WY4MasMwi9D
yRu8RD2LocoImqoSpifojyyK7xm/7Y1lUvwm+r/ULynwCKt9aaQBNhS3abmqlarX
9E0UOO9OMiX+vAUIY1tYxuMlw+qTQzUAZzj3Uxv47e1BJlYeCJ4LvD6r6tJXMCbO
rv7pOcnfnsnltJdMyosivNfYSgREYBQcO3A3GA33TXtF+UP59dWKQV8Mmy9BuX36
P5FR+0fLJTnWncomW3kwNiiBDL5upYcKrydlzhtWUoCxlhLdNlmwZojnpZoONsUw
unuz0iHqbk42dyf+yq6NSgo5H6GqxoBv0MOlEcR7Mae1rSS+m0pKNhJujFG2yxIB
jPoWTL3lw200xWxHGPZJYysCx8Tqo4IZ/xukQMR8Osi6Y9YIkvnxMr1/a55Mv1+n
Ena7z05rEdnpwy0eiGpBtcjfVRCW3E0pBqdkD8jOhskT9FniekWl28BGqJoXi/ZF
28gLDG4GKPQjSCiC1I79yk5tyCmD1kpeGWyJtxFWvQMKTjQr7MZxVp4ufcjbNtZQ
F55+FTi8T6n1S6C18bqK5ssm5d81tF/YyoTl74L7mRX0YkFJrQUgSW6p6rYmhVed
0BsgEeyGs8PY5ikGezHbxDO6VzkWsRLkpkmiuoCPlm447/5u8ZSwRFeT/VmKf7qp
eXtNtskMRzGQ2lTgvCB2AoBNXk+fgrs/Z7o5STAfqSGr8EWiwoL3RD2oTuxtWbJG
txILlwiLsEBXr7xyYfLw8ydiWpBoobBa865vaxbBmW5j/O9bvWJZvbcmfVlMjQ90
LKNVzVuBDHTLq4N87md7RMzc2HEE9Y07k2XJPU5B7SjRSmGISB/C8FnhRoEPNnnt
i1RIpnAdWejMQlUYx6FUvusZHj8dmwD4xJklTJ/og9UYQ00QASnT0yswtjIZNWtT
rAA4V1UVGMW6ZzZ2zrP/iFauI5+JTfonQDVCAALzoCnypSZa626oRv3eJLOskxHW
R31SQYwN5myDa8136/JRYpySyj1OBjx7za560TEF6l/0bcDT9v/A1VWR5WQJDQaN
9BkEmqJqfZFq5sJQu3dSIC0qLKhogmolljKyFqHcGMtrt/GqyAJgoj0MvHfoSz7J
bct838NeJsr78WgBFnqwJtFFpUluimwfzXbdPNKdufKxNmLNL7Q3Np4eSq5HFkXX
U38Pq1Nd8c5Y/7LojlrtfZJp5yYG8xEkQSfwb2WnWw9tggawsQRKTygfbJTKF4gs
FAvVMnG5nKOXYi5HTIimhoTbUuC316dJG/pzCyHjyU93Fv+n1tFQ5CDVczVeV37e
RajUXlGcfdlA4siFzrm3RxRkrY/RXa+F3TXJfoHgNP8b/t1gqdBWeccU+nz96RaH
UEOP3udhn7oXu90sNm8SCsx1okRHqpqA+dKrHuGP0nWUwbk06MI/CPXYu6qWSaZV
VpF4jWdunxRgzm3dwZuLl4o6ywRmV6oLC2681umG/F4QjJTMwd/EEO1ykWbaHGIB
phCIDlR3xz7wPsDlobHtCnO33tXAMCQL7OhoAKiBG5XiCaQ62A+wssQ/mJO+azB7
cdOJcXIcW3wa2EX/JqaG+xb6TKWCLwn4sh069EJqvINkNS4v1tZbXW1NXN5QZ/m6
hEYE1CKJbIeX49aplvCY/WJWcBKBBjgAT6KuUzDdGopBepqHtiA2QHYG1idsKMLQ
tlQaMZc7Adq+J1kaSWZcQWw2C+vKa7B9fDEdn0KEGcwFlDiKRbakU6j7OTAkygLU
6JVF4ng+k28Z+iqTDx8CdkMMzJQDr7UNx3efKU4tQOqP52cl14eVMUmepFifUHHq
cczsMo9X566PEbemyPwXvk5t4syiItnUp0P+WTKjJLJvqmtkvVbLRgtSNwUAD9AW
ndE+2l0/t+69SuI9jtgwHLkPyuWpPz5w0/vSCwUI9JLEEOPtN7Dfvhasf4NvJDpV
qxr/1H4jeBFCaPjSRHx0CfHBWbGx5j+893ABXTt4c4/sh88+1TDBN7KsPDrzCZUu
I5SrTfAyW/WZMGWPKfxhL0ibPTxGS2iVh9b6VL0iJ6y8xjbnfV9Xy6ftoZrjY0gd
wEf3I0twkM/EC60Zma+Erl/nD/Fa5FHS8lI2AJSWI5Qain5vRNlL590SpCHL6pOc
Z5KQUb9LQ70UrDM37drNFTf13zIKeCcxk5CTmEYOAq3AID+V94yHX0XaAE+mh/i/
W7FlFI6y33WNUpUJ5w2cJnNOqRP254/rXSglSh8Gdb7OB4nGK3jplVoebxuYZM9e
bkJYQzXtXZqfsBbV0Yd0Pd53cF8f8mzPuprvvB1sRBiy0e0Z/penVHhCTdbPvxCF
265WwyuOIN8aupzea9QYhaAPgqmdIWd3iSIw29Yq2ym0FZ0k3y/sOU3LaGJ1w2Kh
wnzcqlM+9CADC/k/+tB1D+gIfN/5LV3Mgr6MQnkgGOizj/3QVsC84BMsRXqM+dFd
z54ytUkccYML+NcVUSJl+XHH0CT4Czu26pA4bx0vGiwaLhFQDJbYtXe/kQ0D+9Gu
3BteGE1EXF8XyGh8ejdTtVRu4P95JyPJLohUJo8dewYvxHxae0x/Y7WGZs1yGfWN
q5UkU4rXqWIsgje29PYZqVl2YeFHTF2rw1E0NIIWIuJUzOzjneNb87OBshjRbx/x
PxBeQ/GSEpaGAgh+Gc6G6QllSc380HHAmCUoDRr8bPBoHDGbY8g4CimLdNY3wKT8
TCqDjFPPFqfVwwB9zEKOaCSq7gKvm4AQiwrRHO7uMegzbfA9RIrBE+xzhMTeOOZ+
dD5PEhbnzmfX5lV2h6B4NasgDUL+oZVSl1QNBDHaWmh1HSU4JQioI2dV1NeXEomS
u593WtE+pvVyUuLbbFg6m/vNqRbYGw/aMUZLc/7F9QLeks4nwzvZ1Qt1TFb3mt4r
q6yyDsoeXwe18YwcbQYnHhsovikP7RkxOBnkbUYDbKyyTmS7uKhcDQ/WE1vCWPyV
IO2sNB3Pheu8vCWEPRA9PKwN7CzXtiP0Q2xz3due20zzbp+ohsKx/oIc+n+EsrdX
uX49reJuUTvGXO2h5IRHsPW+CWCqDF7DgjwfqEJNVX2xj11CGw+NfMv+i4CL5WXw
L1U2i3EspE8XKj3PxFDSc4odpBrWN9iLVVVAYxuf3Hnbopx7ajGuVyONtNMM4aRw
9j6gHSsdG9i+fCPlBNHsStrNZKMS0aMuWffyH2tlldehbytxDb21eAMgMInVmBmq
+H6ddQAvVlNnAVdw0jr3e7k5glCjYnn2bfiNBQzk92uXRib1zBChROsNAmNzQnek
g2ZIze+A9ssZ6PkkWo8cMzwBIr8l4ijGaObTXyV2Z12w4jt9vAm9JhX5vl371Dvf
lsYyTXUGqhU2Y6/ZTHNCXmrZahX1MhiQH3QK09PL/kj66bkdGZZmEphKSbNn4B1K
KNzbCAX2skV9v/l/qs4EeimIQA5+vMnkPFdlw8BLEF+8WKL/qh0jiEwt1jMyOomt
hVYLkUp5LoHZyrdJGxQZR0P2Tywxd+exrQx5XtlGAgzTv5+bzyFwgm/6XvtO93mx
U6jC373xjxki31iu4VHaUQh7PEgIeNALCBJJlQl3SSIUmXf6zG+gLaLJ3f6nlv+X
P9hK1WpxcBdpUGFOVXkLavliGsbwdZTcdBzkw3uP5krS/Anlkt2noy9vPHOjRjJK
r0S0Zo71uZyTSXDg6YZjBO3JkyTEBpKW6s6iUogPffiLAokJm8V2W1R0gtCN5XIH
lZmyIM+9XehUiGQM5cKLx8z8dHizun0JRIuYONHqt4K/sPuVLIPsDe0y802qA0/M
EL8qlNH59/w7KqxtFjjspwzSGp65eDQT+nDFInhg7uAqFMx6cA1eUrSpS2J2h+yD
P6zuUmuXwA6Fr5guKrJSxJNc84NCkhuiuYa6bqku/T2Z3BIGjaFn2vp71A5vK7wd
qNkqKCQpYKCKv70nbc9Xcr0mb8PBzv3LPY5APiRvsX5/eewByn43JpDb9NFuY3Jl
POpnXt2q2wy2QkK+rhhEj9orRrAbpgHJ8UHAGIBC+n0bTtjh7d6FkL4ba3KCLXM7
R0zGsa6AFCfY1k5m6opE01BuPx8DDcSjmtGRv5wzv8zFKx5WK6q8aWfCJMyywFGZ
iLVhEgwpQ08G5gZZQR6qrJn84yz9cyQZpLG1yC91L97SWMhuVmTUlVuM/cZKpv4W
SGGwI2lffhrEGrNtmY7XpOjTLFz0mQur75MDbQAqhFNkxHkPUxYya+syW5SUomJ4
zcQY1nl4O1MsGroKRuvqosQQp69OpDrzsKzN3OpFM1Eym+FSYr2pEHebRPEprVkG
+pNUadwq1oqmHG0PKbos+CimbX708xfrpP8P6ViqeJDMXFPuhh02gT0EnuUwL9mB
0Gu4c5teJe8aGlb3MdkhL1GKPPFd9kY+XLC2HNHFVd5IUZJXxmEwAUyZWD0LaEcf
ZI+qKFF+uYvLmP9Jsh5/fADT4LnrCj1XEXfhcYEVzOsVuSFwuCF0FAH/AKV66zHe
3TkjVqJNEjeLGr8MrY9KGixOL2AUwi9N4gbvWcf21DtmpwBqL6KsnbQAlai1V/Ow
ieBEsXVz1kMTfe183cms73jrcuhFrGy0rHjs82RuJxgzUGFfBSFXtj89E8G86cPk
nyuxZrOiFVu4ZxS31JzbveWdB6W8q3DKjVfuTCF1gUL8Y1OAE8BhcE29lsCyfGuh
g1hxDqRRXdi7o06PtAcT4cHc3pEjewNiaj8Twq1dpREkaAspMXa2usuah7p7fTi/
CJ2io4CHVw8jEeY1LX/rJ1yMrP2DzEQ4zIxNj6QnHnOuoFSCHSkKjaTdai1fvzZo
RFGtVleVeQV9KSkUxWPvEhqV2Q2Q3yoVr4S3NzfSgWlGh8l740cTdOT3t70JAQ5p
8L5kk+AQ9P862Kmt+KWATi/npLAtw6FOPw6hROMjA8YLqKhIy2AyB/fWI4afIBU4
MJNMA+bk15zd5YuKWubwimffcdMjitgNdhjeWJ3e/R4qExSYlHQRQg7ySPiEizAE
KQpriqYb5RJw+k0ZyhCKyH/kwzw4+/hqZC64KQeQbDbA6CRgMKO7qgrbu+sd45F/
8GMsLjCZsRDDnFAzPdzyBbSE3jFVr7Mn53F3bns47s3p2DPLvyK+olhIfR5egpqP
4qm3np9SkU3Bp0g2ZnLhOkp8e5M8+qjzchYQxCO3lretSzCdcAkcRoNwnyl5nma6
7308yzFCJNaVAJEjB8fpjTe9wZdLSUNrBnQJk8HpMCkIOYVQAh+jLNyM0Un6Ir60
hLm2CXB9D/TSFE7UWHEKNKzLQKbFP0zZcT2J+D1dRAHF+8DLBkM1bYIRiW8JTdT3
zHPq3zrAlxILowzX2Uqg1DyMdFlIrLhYNsZwz2WDI2wJ8/hNGwkNegDXwoAIOmJV
6pnumQ1r5yGpHfriY0kD8ShZ6kOH4eM4vlkzo6HIKx3+fMja0JU0pzLQX5C5mc5Z
7ssX9F9COBb5156P+XOFoafOEypkjBZEEDsJZPqucmSjgvU68SBA/Ra0scVAxXJZ
4g0AVP48YRlJzBg6oQ5PvCbAfSvnjqbmFXlGraf+I7JUp8/+gvN2Oikaj6NtXLnW
RB2X/dHaT22z1uPNEjcaUtwpw6SBQXNRMQSTl6+xAs+ZUGlNPTtn2AU/datKJoPj
+OxqnicGsiZuO4jILgem0OYd2UPT0PJjFmegxWgd+7IHyfgpPycgwsFzg83tKWAp
VSt+G3Y2anmteKD3XwXP7tv4RuqP/nRPJqpNusxiLuySFjg/kWE+K2f/GSGSz5eR
5qyqkK9Z2abwU662Q6bQqgL0CCgrbTqnnkvUp0y19AdXftN0ChENypUfSQRDVRXT
Fri0/1r/pZAYNhVzHmiwdJVkpTuVtMRccHFI3WLPfExwsA5TBH0tScy0XQWnQrrn
AY8O5BGn3GtCfwfl9lBcA9kUAmqUuIrlPZm8lxisuTWYvXmb3JcnNmKoRTnth77l
Tkj6w0HVbk4GnC7vL6QQsrvgu0sZpykdVGK1u4sh5pbmHg+YlQLkAU3Sj+16ORtW
CzBPbuKnSc0evMjKbiBrr/X7JVt39t1b9+oFas6Er7KdZHn4PnZyoM1TmW4QJFOi
9E18TX/1fzvdSgAliMdjoBD8VmU/0yDfv0MkwE0/wpfIyZnaS+vUt+Ahjv2StrKP
NJUzsFQg56AbOhO8NSw3mkooQmswMBRiRMDGU7r53E8ET7bUFMppMmOawgtF5RRF
NfPiDtx5TuXNEZa++SUxzQJxAt87ulqhKcHyW0f4eHgPEr6hZEFVg4Yd9Q0tI5/r
C/eqeIx0bjJi1OAplWVhe9H6/q+r0GcrjmYjCACl/+175IhGxsCDw3bODi7+j1XF
6JgH+CtLwv6a92KyxZE9dckQbQt6AQura9gtZ+N2JUronwAnyiWmCRGcZbgHzpp4
GGh7BTfsLJD0nRGuUScfxBwBPoGEug5GY2DPupwJP0iH2PNELKNP03F3jpsl+nrg
oGNFO5mYhVvvCAsX6peZF6ZqqDlSUIYDWbASqgFBpEeARcFW5AHgRrshXFJ6DK/K
dPPZKhQmPVjG+4LkFqGzd21/jbfPPLPWnWYbC1gOodfLWSoXutsNMuzxTfN/NpxH
JlQo44FoQvUUwpyrcGpwftpj1RxH2qDGeScudLxKMtneFr9XE/wukmggWWBIh1vi
nZ2B+eykUI8JigszpMW6dzQz+XAJd0aFbSwYWI8H0aOMBykaYsZZvCfXJwJvYAlx
H01l5TtX+MNz/8IzSbeh6mXk6OUW4gI/UK6di6jxeBTD6PmBeQ0VwOCtyNgPFrI/
X7GA0o+xcmgQ04djokg1XlZAZObILdlFCk8Jw3l0p83W7ou9KvIZdyIiumdXaPq1
XC00xLPSe70eT9jyjzxJxpm44a3xGJuYssNlnLGIvAdaVqgRl3Uh8l6Fl9sU+omV
RGFLGNwJ0WGSGf+y/2Df142TITmBwGvZjxj5wtrqRsfMFuUk3JA75LX0yBupCKMj
ajhCxlrJGLb4H1CKqypEMPPr/liLs++37gBqDeQXO6T9WMta1m7C2LhXeoSxTT8X
O2mxElIwJdM7yu585WZw92anq/CYfQeAXZGilyv8L8B3eCm4yO732foGgVBQYfk0
gRosA9uUNdUhjcC0tEU/ZCm4LD7Ey6NUFEwgapBJ3LH/FRQ8Iy43oaTbgfM2k+ix
0F7PtNnf/0o7HAoTsDM4N4qtn2AXDR7SVXSukjaTcP93JkAPXU5Dp6Ahoy6669Uk
6bxXe74Le9fWMr2m3oI7MLXHe9FxqxqQ8qctgUEHKx+orgd6+8E6CO91divZsqd6
SKu/AU9ITDZEEc40APjO6pIUZHs1QKf/QjGPF+33A3zHSuh1UvQN9a0dsyB88Y+g
xHquAUqCXvheCM4j+n19hOtayc0wG4PIWQIXtpFDD0vlu5DxAYDkofNg+vDWlHbR
lrLvLvP2NpJW3HDjGa5PnQrS2GRKzFVzFOu1MxyCiKljBC7a9nvtuaog8k53ge+v
Z70+WXzAEbQFKucaNA70KAVfsHHi9/72p1G1QGPuu7jqcBLhMOEar3IjTYEChJPx
/EBhwc5XrMVTO5ZfdlvkNaLt5z/++eVOjcX4Q+FO/M7weQExYZPSK/VrQ4b+VDYD
wnrgsfQA5XjzYFo4lJLtuPhCmSaFEkYDOdH8VEVxKy+F4edT7dwU6ty6cALDCUAl
qn3yxfdba3hpSxltt4cCu2UysLWtguaaD6umoSqKn4RhSISrQGwpKaWCSRIGx9Nt
SOkHDGG0zX13HPgA5/kLyZK3BBDWBiF22ng/iEL/YX/nZKe0Uaz0HCGajyOtN08/
/QxFDUj/yqfZwWUWZEAoFc3vQA2E4VX0M5DTV5fc2mHM6mb1aVTtLR4kPC37352R
ArqtROtvTcHJCTt7I3iPgj24piKpvhbBTLTdQMf+Xa3DDNYQM6/pHnwNGNlvGzEJ
3z6u+jJRg4nwFsafVtcGfN3mEdC5FVscwX9fwS7sDQthSmJcl888uhKFe3CSf/Tt
nmftzRlhxQTvl2R7nGLkKclFzmT60Gih8LqtgH+gwvydSioPS6jNL6i6f4w+pVHX
8EDWl/7BsPasWJYg0xcjLPiq8DN5AT/EU8kfmuOOImamt1NmSoV6T5Ua0pYM07kL
BdRaXLu66DNsWdoBLYl8eIhjMfnw6sySt1m6qaIXlFeh6Xbyh6O8tkd+DDKHk+9h
+DelNW+NvENGZcji8tzbQmx6XnmFnEmLSeROdwZV6icU6jKRQKaYQ5oN1VPowbN7
akkFrNYglS+1D/h61Fe200rD3r04Y8NVOVh/hU+ZBOiL3O2CySI6CURNt6SQALws
ll8pmWEMzuy+ewTDC0b4zdtvfiZ5WuL5EWIIDZW+zHon4UABeKqZG7OcIQQKfafV
rak53WQMdIzsc19mzN6oSqOfMwcs+KBwU+fsgkiIbacqh4KBcAJum9H+j0ucAmyZ
rhBUeWgxO4oHqxq7IZa3shBbVww4MNf0aDhqg8/2kDbx3fZ56XsNHjygs8BcyiO7
kU45yZFtg8epGj3PxwlZDSs4Q9AGCK/pCAvvELzPAMzmmqbXXhtF57mnbju5u5wa
c3rv9/DIE0o9Sy6/EUCTRIH/t5qZzmCuKYh0ixPOV26ikB0iqLdDetD/JzZNy8md
TrCa+rSjKgykIwpn+Z5q3IVWu9KmtIO+iafdciyTNwW/1yOGoT2CTr4ucPwPRDfg
/U6HoJ6qi6o68UABSiYNOg4lfmUL3VoH449c+d4KBtg+gpgK2njP1KjAqN5t4c+Y
ffwV/Lw6n3yEZE0Lv0vQH7h8L8I1A/n750BZAbuJzK7+XXICGvKYc1yLz2CHKM1Q
39qAp2GaoW0shjCSukvCrD1JeRlPriPA0pzUs4Az4JlG7Mpp7InwmgN29tPblNWi
ePcy7m2PBH8elQ1e16XJdmJ0wDFjt9t2AB2zu+03p3eFubvfk6ryNzsfgcV9ZZzO
RJU5Lha9rrr/8rxtoTJ7okhqMbfxNtjLX1ashHEHFcLgf/4Kmrei76IYJKivssI/
H86ashn0joQ0E2cLBuQof0rekC2ze7IwB2Vqy9o/IJD9jzHu59JM/64X06Bx50B0
PglZo0tFcqadRbl7/lrnGqMpCFmfN9aRNve7rFgVVeFlzOKmR4UsMI+od8UyQra+
AWmufHmelJtdtuMWh2juA3X21PiDIkaWtRAotxsXy8afRWgyoyRk4eMlL+1uYic6
FExesc6Q4HuCIJe7tgvJT0z4T9FLuY9fKPa6FyNllaI/3R+Un41h/7bSJOrh03rc
kPWlb5a8IeG2k9xiAFcFQc93o3Dez9XvZOuXYWkIxLiMp4/A1GRGCuyzp1EgzkC+
BODeq4UgaO0HBz548ypWcHjltBK3NsoKZ6QQiTFeYKUAfD4SqtRGgpX0jwQMVFf9
ZWhkDz3NuiBwnSjXzfnyhCXA1K2QZYKuRBgdWcWPJqiXMkeCrkRiQeaaOEvjOa1L
K16BncWA8HY8Pr2HbTUlwicpM6SvWam7/NfvAiCvO+m1pla9U8MCi8OEVYyy5hwt
Urtwm1APOMThaGPT0VrA+wdFcyz0wonKA0rjMMcp9VShn5YLenFn+NaiKsdCGKA9
h4PlT79vn33ai63AdqpjHxXZeiIlsfkED8PU+dtBW8RTKeq5iT5mzVQSzzTVg3cT
lFjAXrrGnDPVY5GzXBSfqj39u8n2DthJ1OWqydItRFjifEmvHfJIKeA/8yYWWxp/
qygH5VWHQPNsYPT8Rtx2BDHsWJmvHbDcP1KhHVBKbY5C3PqCvq2zPYUNYMxZPTP5
qQnoERKFPdbtoXZRPFpFMHx84fgo8zoC52BwqRfFuBLIysvaVBZcZiUz7R8ajphB
pD27XP0NpYe68YmabgwK/4scbCt0RVi0W6L7Ex080L2d4Kf5nFDtGcaaocyf4/2F
iKWyxOMM6KBjSXzduC1cr9vJlfwW+FX23XQLyU2co6CGjwahMmi6QJPAIER5yOzj
zOB0U71++xBI7ufawtYUDyJC4xpxofZBAUX0PqdkGcSvT+6StA9f4kR/lGMkWJYj
9e1fCT+5erFgwAoND+feS6L77GrePlY2QHG3WxkhTaGsWKRUDsHqrMbSNJDBju7A
3IPZzqUZDAMjMkzcV7pI+KVkG4nl7tjFkzJ0QexGkJRVNR9/bZ8nfdUyrN+GaVvB
lCX7J2HwLVK+8EoK6Jr4gNvOPNnMyT8DXnq3XX08ET/HkqSXinTMSAjCxW3urIb+
9avAecHK4RkLweaBSVff0p+vNq4MuBHgXMF5QsAUPXSa2OtdfP8N/eMwZqhMc06j
sW1jACuGfTPQn3xXwuEtvY6NlDitaq52ThKZ2A6B/fL94fg4H2vcipJJJxcKxsw8
AussjfQaFHdkp8p1LAH/gXPGAtjEqQGRwB2+PInrkLWexzETVRA1L5G32hBATEzL
1HvaqfRhcEcCbbqK58m8yUt758RPGk7vl6fZ2r/DUlpOcryGAUJZqPkiMfCXUE4V
DMJ8qz8hyuYsx0hiYZxbjUKDcYUyYFHg+U5zfB5Ms7OjPA1kN6ajzBFzWoKxisn0
rCoyA9ghUeqSEon+WhfJkqO55Dorzi0DMdHarLoMvGFoyeNGqQivlMOnIovurr2S
FmYW04LzWuOPgzMXCbUFJaO5SEoE+asn5hdZJ0QxGtrYqxMLwj7VRPqNTGl1HF78
94MsL0vekg7vzuxeUb8Exv8m9+LTDKE8Ch18cFP2yMhYt65y2uhnY3g4kP3TxPyj
yyj3z0k8lqy9jcz22yRB+V6i8b5PgiGV0Ructd019yv4mO3z9gB/Gqlm6WsfCGqt
vIMSpqxv++H/rasO6AyGJL7faW4B84uJur0NvRVzryVurBLYBU286XGEPeEO5IGR
rJxi46fmiI5epsmKT33LY//kIEhQeIw0/9rHrMlHYS0u8rAbd0yCNBDZ2a75NU/o
7EMR8jashQNtuP+LyTAXtHLe13tyrcNP1mbEykq4yZqUOCrsetMZ1jQOW0yTrMOC
rHjTXxn5rYVvv+Le/9IcYCvRfU/A+NZMZpXG5mgxaHZ/uZda0Mj99f9H+xgErWVw
aDEB/olvGgHUzksoZsHfzWGsFX16qv2WopdqHpyXPqlvVC97JlVA8HnAD0evDk1u
tHuG3nhh7wCT4N3bHxkae3SiDwmmAVLfimwlwuNKZtu4FJR7T1DtaGdyf9vbPx4X
P6kcECUPEll9dX+XNwhPhblIQjpIPnhL5wLDyPqdluvnPWVuUqjS5kFnfUoMLWPM
rBBjx2VmsR2wW0KJm+Ks+sQrz7YjsvQiSR8cWmY3DJowSsEQkwr+6FhmByVXG3Kr
mQp3vn08vAvxuHKEqSGxcKcjLWtH1yQxVihid6ZRtEpHBJDj6H6hIa/62VJ5zVb0
Mz8hiyMvMdQtzSRpMg0oeoLhqin0ETkqO59QhGaVbMwOo4cnR62KnwRkH3tbi0Ew
lcnUVYN5bHBZsnYXnPiV2T8pChjgimo8x0O77Kza7j0DI+a8PmAqYsxQVUKvYDKP
KNp+/M6PoTyqbbLmYishsizH/I/TiKWr75ApKtF/9m4IeqGI3XBCOan4RpkADaXU
4PCYXExIxQtyowZ54hpnQ2LDM5zZT0IVZWX45Z3XxR5GkfwpO9hwBvjB9ZvFKpqg
INY7RQ+Hh+M5cbR4v4PRtKrGK+NIAJRH2mOXj4MoHv9AjdbnaX8+bJBW2lfYuZrR
mlr52ei7D3YIaQi/RzK5yyFpz71uKRoZ/7bgpgWbJisSfTqG7HVKfV5B0Z8MrVHq
zA9ovXJCwhnSIcuQoucLBdIcBb51BRbyK2dTn4emUCM8ucYrytC8x0OOeqBsfJXo
l613FI8s9qhQoyR//2J1SvL3rxKKlYFaYeAIDLC5QPYwX/WhJHzDNl5zM/AK95xN
MkOW4YgmoLgf8G+El/fR60bQ8e+/5YOTbxUw6PhvoXOKVWI1um0HdV/zy3YHPPcx
/xKO4lMG2UZTH9ISgwFJdTcamJxRmz4L387rOxRTUsbVuNxDhrZLh3UkDD26K3Qi
oqOgGkNJ5jbMRxo/sCPfbLu9QyHpOfZoUhBTtBj9FCcgmc1nysst+PpA7uG8WT5C
0rKKIwQU64VbdmQD66GnOMsjPrnbMADWwP8dlQsMjaq/ODtwmkc4iBWpKCyo9b2U
7rQrIPmnjk5sGyEoPatDfWH6OTMZ/FhfUZg8aHWvbNtMU4rnYXT9QghWgrguJg8x
8oxo+n+zaOzuBhD8IIh0N25j9EhUNnWuKLDwiRo/wYtnhMN/xk0a+8Yl6y9b4w4Y
Pu3b1QpfV9ylfUobGkNeAzWlSV9Z0AG1kFNglreUQlEzRj56RwIhB6/RgebjME/t
Qtjrt3Gf+7KToUTcEFbFA7ywxdyrZ02V/S2jLslVUU374kkCFqRMN9BGgyPMdfkZ
qvkvJ6HF0VBgpZ+B1IXZHhk2C7F0292l4EQtWMqZKvF8cpu4gIaazSStNVyIQkp/
FJQxMQRr2FJ6V2RAQVv1aElpEISILOS2+W+IWeRVUPUk83czWht02eBL/2vNH2NA
Ifu0pYG3iNcmOUaSqLla+sViqzR0PulCnlAi0MmPHVHLT77ZtbGwu5TnhIlPk3th
kzeUkRZIUihrionFt9xjkRAEJDCtCFn84Fqjsdvvahmh2+wM4kLY9+I13yKpmPT/
OVOIj+EBE5ZtpJEJ4TgRAoGM+03Ys3itQkcUCkG+qBnUafyfDNV7l3rXNfDTYTCV
Zk5zn1QRxfYZVt0LC54SrVty02P62SN8Rq+OBa55K2Sl/fPgTCZ11Tp/Qd9nXmgZ
caFKkExXlpsV1GOoizh2jW+QKHyYTXLp4Se/GXOM2B68ufuYp04Ea1gpkg4YXZMA
MLsVkM3ybC+4y0VUKZos9b5ZTkQ/3v9TtqMMd/TUrsNe7x2TQ7TWGDLEccSEcwlq
bbxtzEpw81WhOh4MNujJ8svlTHoy/Go3miPR0SfGw9QmcVtZqutZV5O7H+kyMTgT
LAg7qJ5CalSA/mOYZTjhpfy8IuyDx1IenHfLfTsEfQ8zpbW9yafKagVHyEJMFAbZ
dRu3oUi72lovZT/fknSKDVXzRpKPI2/+Rl8MykYBek2kRioV5UEefnPYkqbzz+hG
NoHy2OU0Z6BQfqeXK4RwAWFN4Sn5yyAA0ezE9E8spYf3sGQIgpdGjkRgmws4/jMY
aBJKlp8THe7J8qjJmpT5WPGAClJTwIirSzfVMK3XX2R9EcgioozVdMblJwB8zbFK
MguBiaFk0hx3X8Sm+m4v7lrGFQPvaML1Gwv57//rOGEPa3x3IkcieUwMW8GIkfcD
kdgcnhX80FX7udR5mdfxOD1/tdqmN7s4hKudA0lE5xAKom4r3i37Oxegof+E7dIK
nJwmEhpCssq1H7///qhUMbsYB1KP50GlL1hZmDPUMISxsW9qiVYSdLT5Gn7YWTuW
SW/jmxnHuQvUnXtqESDxBV7qmlNpaUVET5sGIsELjcJCqlZenadHYWdBM77+uTvH
6SPJyPv2oWzjFL/BnpMMBjgtI7aUUVErlSqLY2434ieCqkJk5+XLgQSSRhYc9ThF
CNKON0Wu8wIvZGU7nGSUmQQroZ0Vg0hWd7TSuuq2JBgiH61u6ewIDIrQnB9JTmdL
4OiTuyv4WNftwIdvRbMFt8JsX7+ZoJFgWJA7kaRMA6B1F/enU112S7f1TNx+2FlG
mxQt54hOLwyLgaoKIN2BSPCgMv2Vk1jE04iAhCiMNulW4oWVanntI5wrilXiTP0U
cCW44eNXb6JQkGsGzbeO3YWy9i1OCmF9ZeAJ8923SZKVW+uIXOvV/QsI+9oUWuZX
apKD0dDrFBTmlVdsIdc2nYWX4yp/KhvMhZeSymzkdtQ0xGkWqGvnsD2HwD27EMNi
xCdr8zoGUa0C6N5UFQVGdvJAKu9c4g4hKV4ygPOU85vAkg4SgvdhkXhmiTHTAGcO
lY1FYUwdfXsqfqXOqBCMvGo9ViyrgatJD95csqHoc2MypnkZM6UneqiEXN7SnKug
YmhZqJVLS36QSKzjYZN+uUEvOxtA+QkuA0SWJMj0+tJJbRZTze3TPI53WY1E9F2s
OuDkZHh+C0Yj3hjRtr+tUxxwUY8SxuQTmBOCqGf8ZG7SlAnERXyKW15Q+7B4hvrL
fYhZnRkH9u5h9CccIbzwvLdIEvJv7W/6GA5xBrcWDuQv3TeatTETwOGmR81hqhEQ
RlIEEqMdzQy1YcHg7lrlLi9kMCX/E/MoRxpByWs1tBBKvnCMun6LiFjom0m8papm
xNwDZgN+mH4q1cJHSTlzUQvU4EQh5e4A7Kchg56jtbaStVtbk45q242yJtlxCMsJ
RKi7i5HGKoqAmG3WYKGHfoj3wwRSS1h7ISd7D0Hx4avn1pFElPxBw94gYpO9O5+V
+WHVI5VdqvZ8L+a7jeTTZNd8pBdhIiCtczYd5W5OdMJODz/mGmaGpzs9HLx2gAF1
u+igQQnAoCsXd4az6Py9+x41WCC2SAm1g6wvOKRtCJ76hnPkdvpx8RZXRTs9znRk
Zg1Fb+e9REOXlVpPEtgMkiY2b+jeofmTmekT0VEQsf/ZbiiDP4KxgzqWymcxIUXI
txEr7pyjwpYZciFZtSFyyJti2dQQs7gLDTDU2LqGT/K9dXX3bxnkwPV7tuz5TPrA
AKO7RaSSep2xJFQGIRCa2B6KmUP/NcEzVwACxml1qqab54+k0RgHEn/9tuBEVtol
gdlZysw/A1UXnl5RtnWLGF8PwCOWn+Oab0pQ0n2PXTLRA+dYGAHEYGgssiL+3eAd
JDgnM62jQl1PX01tu3F7lYED6FBjNlZ1gwkYVnMaEBs9qbItD4Uf//tJottFj0QL
WibqYVmRsY9jSLQGtZm7uu+tL/ACCaSsABzy4k0OuscnGYdZPqeDz5QR9cAhAsC8
Q1YgE82b5J5uEMfy3bjTO7Y5H7L0IFbrkaGDGeszQl2lty7dtbMk1d/EPCfd76fB
/C0Bo13JEE2iJb/aE5WxTqjrZGjfMSxCVXqJE9IONHtsAFE/UYy9qxs2zxHhmK3+
J/Uj2RGhPlA5NBdRkq/ko6O0cCgoDxSYBIbJ4dk758AgI/oYjUMclhHSiER9NV4s
9DbTfjmQIw6Q90pTSzm74aiY0ai4pAIg7Gig0g7k9Qon3cDXfdFsJ6omhSsEQTxp
U9g6v+LH9v4mXwiq77rIS/hikboBqHd07Ih1YQ9TRg6P0FVVGAQ6W/eRqeIm71zQ
EKHVhjnbwcytCgzHvEg/qPrAMQZ/E/v3HXVqZ330tSdy7ronSnSUIlkOopLUdpxU
qIUffxNqjHxvr7TxPeZ8uexuvzuXzLTjkZnhzVQECnN/bA9IJsTNx9lmzqzHhWSC
Y5cGzjx07weIu6GHLz/Geu7DSUg4kZVsifqWnysh2uf1niZRKbvvqa6g1gKe9Tlz
Wxbzk7+HsP40Jm3luPkD0KvkQ72+9L75lK+a9HBhTd6QbJK7bIQLcd1/+blmm4xa
J6FEegI9CjoF40hE/r2anObWLPFdeOOY3kIhXMxuigGI+DJjbNNijIbxaYq7tIv5
NmabI/so5+IMk3nnOJ6s0Xk5hEGrQqxXXYNuAMdQZj8nqH+O59U6RhhchlZrhoqx
/ADVIvj8SXf0ZKmrgNygTo8mUtoQ+98dyrMEuYKY7ngYJ2zXhzp5l7uPOm6B49YX
gF3iNJFhehl9nltgQoqSj5sOblINfUi2HOntWqDrAFQ1YVjNZfclivpCWNvjp1Cj
dpbli2s/A10EwZgngvBcHv9JIbDf8EGN/kbt7pys9squTdaIR/fORl/IebdKjwnF
h+R7+6GLCU5m9uWAaT95XHRJeJKVWdQiu9mksNGTQoN3pf4A2e/oVUz/CDYKvXjN
KcLok30+kTgzuLhJELJDL+fFc7wK7wqEO2RYrw2Lsad8xfw12+ThJkcjKR/0f8lz
PYRG27lHV1dfQ97T0+QsHWc0APeIOqVuwqPuM2pQthrkQcjXAvDLxbP1G7yltqQI
oJ9MssM0pCPyQ7BKZaC5/MOW1bgt3QmTfJvf3PZdbHJvsnZstBDWrB9L2hM4YR8Z
jjl3eDM9ok4SL/hLuGihNsaQP/sLhGdrTjkxTTC6hH98sGqFuXbqPEkLwaba7aZO
zq5fuFjudlueOYwDVuWd8b8z98aEipWZwYk4i0Xxz5wpCNCX69xkO6P8s5HvtW5d
EyDzI9BVIIuNpsJhXcqvBhMNiOZjdyr+n9rA/cyUnpj0NuvA6EuhqeE9yiwAAbco
d9a0uvC6uU6FWEymFG2X/WNJM29DRb3xCQ+dgmPU8mR3bi8BnX+01v1IH6kAx/7U
t8acLthOQjvjiaRnXJZFa/kP3sqtxU27O0Jrbz81/ltCqOuc72dfhpHkeuPVs+Xn
DEvilowLEFk0j5X/Rf/wefYhKB+YNLujIG+Aw34ESMuGagAd3sUXPtrzXXZR5xyW
KMQVJM318TCEXE1PhSHX1HIEUGMU8oAmWLYt50S2Jfto+x+VLFInkYwmiYdp10+k
ZXQi/Lpo/YJaR1fXbMiCXoJJNtNTZloOTSnA4JYofABreMMKSl7QnT70IXKA1JEO
uxNQ/pK1FZfJ6yUbsj+lR6ovvR9R3arIutuvG5zDKunrweoodBpybydCZjwd0a/e
nEajO0obHKHbDth5eS9gV8Iz4nehzN68aUaQV40EiN3HNXsHwNnKaVx1c9v7Cuwq
bbui1Ee/xYHDVra059KL4M29FFGkqsr5gvFWylz90h62JqY0jfQ/gB5m+CX17Vu9
aHrmkEO7Uk/zWBiVmVcarM661kjCv5n3OV2BtfnHEVk6LfhV0HIlG+nuHuKLHZqw
m7teU32zZLs8OZZVGz1mAcN77TUsVfmvtzG11XSfeqRa7aZdyNZD1EQDZtWNR+nA
ym2nd/yj6lhfgNh/SBfmlMHn10Tjr+1LvG2Zm1xtD5dlOCCTVbMYLRr0flNBl5qv
Mh+R/25aD2Oez7yYNF7VRP1k5zPgBMUdLq90/pJqGJ5s4LkjUNijEf3VbNVjkQTU
AU6Mcoim6Hcn5C5f4zIfCjFPKR/naWh1gGprcVWu3lozgHL/z0QrSEjlF7cd6wBC
4TWgNBguXm+9HpHJtLZn1hdYelUUCEaS1U7+lkOEOXHU0jRgqKQPWy88elAlSFYQ
yFbuuO0P83SMwu/Z0DH++wLI98TKxTpcuFF58BXALEBZIFjvPBAyvIFCO4dU93Ym
QdlSG4tRuYAu2sY/ZCT8RGXkYjXMmJbrjq85G2Pi0WFLBtTnQRVu9nQ9LsFOhbxi
imo+LPda4GSZVBhRzwdXcBnLq+e0qyxQQj68lSYp9a/XY0tqVU9uHFBVP50Xef70
meykY8JWn+J8HEhBWzv28Y+E0tlqSYNM7NqTIRlbiuST08IKOrXnhfk6+l/bzhY7
1wHMVi123liIeP63PiTGyXubf9Uh4IIA3+yZqLUHDOJ/Fp2z5U8xAxzUFcF+konP
Lq/e/CkU+iRKCAsBIpDaCox9gL9eYQGYTbQdoS3xVAafKk2YpgTJpvNRAjZPEfgf
DukpCmX6Xdkqhw3/d/NuBqnlNioABrY6U8UiCI8ZHH2I9BjRfp9LRJVffoVyaE6I
c6HwYrLo/foVTVagMxyW1LslkEM7rbQkhpNoTo1zUUB48uKPvrCHLxzVaTgL+jAp
PorohJjtqss5eVyoxzB5Wx6vo4MRLt4jMrUAgq0F1UdUXfBFk/zU/GY0zR76hd5b
h0eBItgnihvDGudtSS4tsWYJcr9chKw72UEsIYU6CQ1mNjCGSOlrimSIiVGUligW
Vl6A/1fKrRUpOezntUnrYZBcxkDaC3AgcGPITzW2P/yxloa8D1Gkhgz1oBbyYX97
/M+b/DggrluEzcOIEulcxQMDo0HbKetwcy/4XxzKBKoVmvxtIDpVcGot9K0mI5po
EdsA3xO5QKzZUaZfo9B6jdxDBpWrrwYZoDXgA5ce/Mv5kBUvC7GLTpv1g93m77aC
wKg0qqWZE1SAsw8cBVatNeDi5z3G9fX1NGEeR2N8GB9kDatHjlHwPRVjeVi9645A
2FnkZi1OKn6OZ77LPJoLwNTAP3MwVJVJtGnm//GmZ54Yij9PCdxGmZ0JE67+TzVl
NensBqCpRcLymNBnam4maJvwRwjJK7iqIdrAtZCnuEV3DuoEVL1HnkiY2lDygCO4
MYrkdRhweVGA4gImq9VEMuOTmFTzZIax3RkUM33nsv9NzOGO3lgCSYM/xUC/N/qK
EgHufZ7Y0Op23vI278K/uvA0PYXltECbUTHIPFaWlTvZxkDU2RZjekH3rPez2Eg/
l+/xd9pZkCnP2WMSlkpJM4lMsQ4Zz/HXf3whmxdBJzc27G2OZggM2eGpgd+lYmu7
sM6xFzEqgjb2SzUoFyKhgvd1m0bOxzlRIj3HaEcshb6aPO55Rm2C0G1XS0Vn9FTe
o52lklrk+RtRGhSOk2i5MfyH1kvUdDZOJuXT1PpPL7oBhLQeXe3HGUqxWBydKR8q
StR0gWXcHiTIfadAEuA6vv6Q9ebaSdxhML651HjZjDTb7B15uBl4upgySmJRojHO
aRLK5xINhZtzZ457fKegn4iEbOUb6BDMwB5n0SZdjMQwfapn4vScq+bx76Qfz4yR
QNyIaE7BaG9wD8GJhL2PxloWDikR08eaCDYepq/LXUW48kqA8hGf+k0hiSyFQ4bR
Op6QeUuGpFgDJnw1jhIBJwPWqBiyRZ6D/kEBaMmc+ls5WEE1+QBC4g2ZvDZgbH47
DzyxtowTXr4WdTuuAqznoJBIqp/5oy/M+j/fctPm/v2JS3sCgDMWryviMevfh22N
jrkq5oV5FR1jRFEl1K3t9WVntyB/mfRnIhNSQNgq2Kc+5pa7++AD5/sl5yrA0/Pt
adbkzTtuQ9FEIXuO/zw6x2JwBgB2T2CR9jw0nurFDjVo4/EnuEezACsY6a6SujOj
+bI6B6R1VeBjUlKIH6/fjhA3EtdSfd08nC8Vw2/9AcDqd64U9mk9JyJ9N+oDv/y4
J3p6mShdqHBBRcC6cZKFwH/ltNjFNb6pe+6iVEmI7lWoLUQsreZRfH26EXqulGmd
mmSEE9H4/ZbhLmzivzhG+ZOf37Yy7sUOuT7NszqAIHKTV4SGNBXuMHfZjGSqIKhR
+lY70vB746VA9xTBWKN7VmRlEstWFcWDMWPe5x18DAJTTgfaxdyxul21OKk7YH7/
kt5bHgFyZ+SqQyVcnrCeVT0pJP1Fwbq1vw9D8kTM2u0I2DDvyKKszBcBaOfMHjZn
Xs7m6TFry/yrQ1xHQ3GDMkXBvWhwKP/A2x5OD1Er584pBZ8QS0CMCgY1ozF+Pp/F
x1xQVKkxtJKfJbHR4JtSDd2xKkzxd5nCG63u/FB34bnS5+XY0HqE500/BpFWLi8w
PP9V9DR0mkd+G2b09Y/7iz71aGMgF9Ynkq8jQ1/9eV2+GNsyBeFHTxNqpEE+6WhX
VTJ6NRbewRslmJcJy8i4rGmcCxZiWJDbVpm9bh9a+85UFakF9YkwFXGI/H2D2SlZ
RSc4r1E8wfA+o7/HdJA16tjZ5DGzQvF+H+I7LX7TQVcf+1IYx/5A0iBoSX5d00Q/
EVk3zL2TLJ7NzVpHibyhxGCiNzGU7iW2uc9WwZf6yDHxjk9XjTthk9SqjWQMemR+
J8NVAlg0bLay6AeZHn11QhU12hpgmlJ15QFK1jQ4jGZzHvDJ+VO6yqER7v+fgQSW
1fvY2AwMp3Ka357/4o5Vp6Gg6t+Cc/JgU+LFBw/oyLWFXZ0VzmUMYr8CxOfEuuyl
6JUkzT9KiNsFLvNM/E75GARYzEBNusDphdUwHIxVNgVYAwwu4Dq7ARc7L5/iTt6o
VNAMFbrUXEh9M0XJQ/yOg2LKZZOtdUdq5t3AuX0bJT+khJNCndkoM4+7xyBKPK8U
e91ff7R2IfdnHQF/5o2K30+Bg8mg6+Q4zsnT4TnCjFwKJBgww1BWTDSoGa1QueS/
VbHTHdHfHO2XAnMbWrh1FI74k5ZA5KIIc+ORrzcGxWphlxSqewxgSqJUGTHdeMO0
iT/72lw3y0F6hgioe6r2t0YoCmvt2FtyFJlbJD92d+F+UQHcmzrPVf0DKCof0ObY
l5epMI0aY+bPeG9z4tVQkdXEb1c9kwFIGG80k5rSXGu8uH9KUXwp6CApYmykML/R
lFeQcV4O55kRTSxCeV9tsTMc2eeBUN0gqcY4P5RWektI2C70cnv1yupQoSYaYi+b
vuaJNlq6OfAaDhpDWpdK7Sxxkm/A4T9XppRRiwkr99T3QMJFs3BN9NhzZtIYjxvd
gCnEneBIqPXsfCP9pxDfFM8zfe7DcTKswEKyTh8plXZujM3YeeTsyF77UbFQCoEp
mAe88t0rsjCDhq0ZgR+mKKRI2x+LuD67vXUbFRsdn1f20icxlR6UDSdh+kQcWna2
6cmDjS3aoqk6NMmDa3cFBzkivMCGLTXQGLSb6LGGExSR3+47fjJHanPnI7f5TLVK
3QNaCSLteYiLAU/sWggp2uHkXfl7XgrNYHTEQCiSQ9d4ZtcjcwzxajKSHolVyR5V
ahggpThYjDw5BnzO30AF2IGpAZQ8WQn8I+zofF+Ka8aGHUliJ34zNjX9oNH3rQCD
P07MKDwFblxnDOoJHjKgiPlsuSNJjCug3hGX1oHLRv1HQ3m7MdwtJIdMWwKjL8Rq
8xzKC6ZLeQOZbIECD8D41UMC6dJ9Q/KcCErQEZ0nxPDn9oa+jf+tSmwiidhL9SnV
QZAZStPXls/CS6+UE92eg/ViEyvxEny+4jpaAHNjSGrE0E6TKu5HEoEY5897YOAI
zBk4R26A84S6W2Ih/s27HnwAL+ngTfoH70OtLtVAeTxKrbMr+fDLXLxcE5pKF+dn
ini4QevxkxVFwD1O8dcKoMS59dlCZeL431PGGlHBatJ4Vn0GRfLvHjDnSiApICN1
V/xzh1/Ww9uxVZffphMyyIda2aLIggek+hl+mhXplRF7j+clvYt5s3AUlwbtQjiD
Z/bLkxL1OP8rC2NKqJvGsYd00QcHv4NUDkGmJ9u304LGxR5/b7nCVYlMi0uJgx9H
ML+qlEZj+bik0K5U0YBwRNzO45bk2pQRVrWjVrj01tXNZWgIJRo0d1VVRMXtgzQJ
akym6rO/32OKhqptfncSq5Z35pfVhigskDCBaknw9AjH+Xvzp1h1MIgRacEMgAJM
aVKhibg6jkBCkORAvMBaL6ur+yl1HNajQhhKFc70MlZRqVwWQiUTEg7HRJwcCm4Q
m/U3AM5t17uSOMde1cFc+xCEfq25ol4f3O4cjSlKlUgSOHmzp2gXhxX2SMa7NwSy
rDbBBHkyfZCAQN8OTewYEqJLL9ghD2+m5NQGWBEb/d/wiRtEYe2bjwwxBqO+uAdI
U0XH9MZdv9X5aqdMsPUmB89ksoEdZ81r/Q6GG+pVfVdOM38mYifs7VcXl7VpYbT+
YZU+9NheChO0J5nhXRAXflptFFw3Apxcz1ihgcdoNkHIFr27XMOVNnI5DdnMwtu0
cWFmQOMy0d6DyGOZQBZtfxRt7hQXnfk8/eXO+1uLEMSyj1m/VklYiYwu+JNuDHMJ
1O6f7rcHeEW1abHGNiwXEWvV+uoY53BwKRYXoufZbuqL2mlb/vCUaW4UyO15RJ8m
SW7iADSGUH09/mH598Ue9hEmD8ZGWKXKwndiPCDdceAN5/390+S7Axeyqj8YMQAX
MjeF+DVQBX3AuxOQGOroUQ9KFfCsqe6GmvkVcJSXuCFhqaaBfHQjiw9SBBnz+0zr
R8gMlBV9QOxB/3ZWK2qiI+5J/6Jic0Pd8EktMBW6wqcKX9OCkxfSPU1FODz95eXF
0Vrwa43AnPYD5r01HgJPar8X8tbUiX59qdIaAq7kjpfiBfi7LjfJ/r0RtgOBXoec
asMkuSJGtBnAL0H1XEVViKVd+Kc4IfnlCWjqr64xqxdmQRYakKfll3L1sTOxCNvM
Dh9CKrVm32E3ycmOhrbFDVd+NAsl9MVNSmDThGpNINS/n3UPdOUBaEXlY6/6HVML
a5LxDqaqYCuaaDABgaLTHUEEGNvqPqC8OOgwRKvqlkV8F++8h/h/Agbn4kaXqsI5
mI1CrB0ZIxQCI7AFCv+Q5ke48LKdEFUKGYm38fkuUpu6Wvv5/844kOZUzzogzwzj
n3Y0fmCMnNGBI2OfOuOExV/xWk2ZILHOlexy4CJ8evCEsHP45+IfSMFBywvWAo+Z
xzw4FTWF1NOYCRQYdkZ91bHPnA51O/dgFmLwcKtATSOa6LumXdyBdD23wrbCSyQI
ItX/9HJmHHGNj81EvVF/pLSGP2qf68qMrLzdA73qttU2PryQ4EzvRVwflSRGjB1p
719qTI6lHWjuMvO7eQ8YacjWz/5kZGlcfdtutw0gVYO4+o+9CrCuqtv7yknVEy74
9rNWxhhsEAqBzCfkbeXuWTjoDnx0KlmkgfmuqdX+79+J21BKGQdY+iDQFugmxYZu
7UQWG7d/Gc0qywinrZe2rztcPrX163+2+KcExFgH6vfykm//Oh5WgbvQZOTutXBh
CGCYT6E76znOlQbDApvARio96dXovUZCAsWPfc2Ml3ELQBOp/vXJb3B61dV9RQxT
4Ou5CdRm67mims8WBfCrIigPduuDHzlWpO2Hp9n0Tg6+zUNec83/DASO+Ok3eP/c
O/vKHdV2X/C49yDYHGGT3Tmlup4zC3h+5Pp2uKZS/AylKoz49byfhCT+Czx1RVgV
ZuCx7A5X9iqpivINrPppsWYYDQcV1yL5hI2b77CWpTwFY8UfBOFxhmaTsJ5otWh3
KkYg7SdTEBsIVOCUk56oPxQNlES+lit5xG007wYYylSRHjeOgNW9SfEEJJ3tEnk+
2XFBYqir3NOAinMnhgP0coTFqb8jy3IYhjvGGtk55Wtp7zSTSj/fmZiFkCYsPg2t
dqocVCSfObTMTmWRE1LCi5gcOz3A2/6BEdHl/gvp4sHYyAPQQIQento98r4t+eUD
Lzljl+/RB0IaTj611jfz5I2woyKpR2FvKCG4HkUmC2BwzVrZXm1BR5PONg4PqfOV
Ki3Je17mPGv4oBfKaDAmIfTGArURnWCcAfczB76df7hMIeacGE2oPru62K6y79lu
W91O30fo0QSs54cKHeaDKOgza+dNneyDc4LypPb/+xiiDZd27tjePKT1UcASKelZ
t4FQQoNbrz8pFhV4UL12XrmcVIYjrmxD2mhR5xje2F+6J8oWAS9Nf3F3gwv2Q6lO
ls99y4/hBRvngqQKily3+84PMwF7fdcr+S/YWq0/DqUFkdNNXeaLCwAsjOxVn3AH
iH77tCJ+bwCo4oTAW6F7mFkVjzeqqQeGYPsTfMH7l2mnf2DvlHIoj+WPLRH8ozSi
LWUAacrLlxb0IRHcsOGnedtgXK4O9F9eGN3sNDp0++68lRT+PHtL7IYW3O7GZP8J
vGb9OUAEol0v6nK1bVAmsOcgHxYBnbBcB1SWl4PrmMtlJbxKFoinJHlAUX3Z3Noz
R3LQddwfSyoIoJj7Z9i3Oe/hrYWHzTOTQi8Rx2h1aLXucBmiI1G3ruwytBwOsqD5
v2hWBqLOlghnlse3H5oLitLz4anLH2a0Yppk2AVih4C+HWVtVMqdPNgyYXGqtSck
5y3g8/rW2xE6uSW0mb0ojsYQY5HlPvAIhWU+StCnySbRlMF76CUlk0oplA38F8cX
/FhGlOhlS92QQCaiSO6TfPB7qrKTcljDR3SlNIMM3nnV52e+Ysd4Qzoi6PUG5Cex
qweIq6b/71DfnIObXyDtvrtCjq6CyA5vL7exxtv13RiWbNUSbG3br2N3gpx9GcS5
6AXXNs1S+jjwhxlrQDcKedq0b24oNAxfVpC6ztPAq5Y7B46CXmbNFsTu4MpLLjOw
auwRIAA0RvbHrCtwT6neZhxhHN6wl7xpBUhV28j9gYSMvctulnOoSoaNkGlXLFhJ
swfFnqEnULf6l3vRhgw+/p6vQkfFpZd5Qu43nFf82rkkr7BlHeKrrVN8ARYYLVBx
PsnW/4EYnnU1J/lG5W9vn1fa0gAuAQype7c9EUn0AwG2XTmFnWKbd9S+msHToJD2
X7edmavkIHFgNlOAKl33n1bNe5aoM/2GiZEbYlogowTFsyFHaBA2BtAQvs82gGuz
+OsQapec9k2j4Aq6fH0u/igNiGyFQxNWOePTiAzseoPFPbGC+Y6PoT6ayNUcGEwx
x7QpY7ro+VFlSsvTkKcKdTg06ZzHXaxX4J755SNtsELbVGoMOWYinA0yuJHFF6I1
tMZPVBaE9bYiB1vOWmyiTx61EwbEAonLb33vXqpnzpHoQ1mYIj2wJ5WgkmAKDJYY
Rn5v128K399wi8jyxNxnQAMjQF0Jx2yigjAWA6mPvJPTmqKHVUfsrg6byJwuTJM/
o0fvUMPj2eBT2FHyBoiwgiLb0I4upsevvBhgpRtrxPqpkYNPo/CX8i3U4MzbFjRu
Wx2VPr0gEgNj3AJS1Tzqa/rGcPgGKgVsd7sEfHST4UuVDhNBwXd3/9psyDix51AY
pKe0uCRrN0FKet7chdCgKk014cHSB3lULe59KWIvKfu99NTNEU8WJnx6WfeKS/fy
YFpCdWQVJECErG4G6uUFiPJ37Z8u5d6a2OJRhUSB1I4KzdHWQxReuejzvg+iJRxt
FO+4fGn7WgGVjfS84+CHGiCEIQLjjF1mHU6mb+k8nc25lEsEMYKiMdfabXx1ZIAm
o4+XGRNcyU56YFST2/1/mXkDiXckz9LFYb+KX9+qH352T7CUA/SmvnMFdnlzsPOW
jEIwLY9wXAvIzV9/8wm/1C7DUW5FQW1C6Oe0qi6b9ao35lS5UYnXH5sNR8AWT0m0
jOiBzV+mTAmgGQvuw3+RWXXV1LgMwAydUY1vH8zsGpr+N5/uzi8n3KUujUNhvjZR
xDa+jTxEhbYPRvrQdmUfRAMdib0ijfYPWjc7/ApptfQNWPZYCttk6xVzurT4cuQn
8KHfGevAQ75NLAsTuawmbS42v3gIOFiTSAXfsvNgKmwcnKwCqAmmwl/vRQcE3n0m
vZDeLIzb0iC+uZc2j11UlzZzsNkxlh4rd7Yx360YWO/9YHmMQXhxVTvDX/KIypAR
U3LWPs76KEcpzBbSyWYIloXYzETqEXgFs1kYrg0T+wmQX1m/SKn1U1jYZqfOGIPZ
qvd1TjSBohxPojwnIIe67KWg8v5ZjacMi5C3NVxd6DYXQhQfy+BRkIgxz9+Qu7GX
nlhnLlruNf49vEvXVRFAnTA4ZCId9raJc0ij3TrKqR9pP6qqCHr9hKRKuIvOsh62
EAzpmBccWOLX563CYQdANnS5GpP8zXn6b4uqv6byju/9TCjh3Uxia9OH7pc7mdZH
eHNmU6DKnk/K8TOS8ZTSEF39h4MHiCC5EggPV7qAgC2vlG5WzPCnCwgS9JxlT9Rj
nMj8vjPHo03qsBGZeOGmJUq6zE64sfZ2xJZFlG/hkyITF7giHXhol0oom31NEDkN
HFYQW0nI4s5aJgfzzP1O8pl22UdrTTRUCdVHj7+a4U+Rl1DhzX01mUFQZT59rI9r
+RW+k4HSVyugtGinSgtLzT0NeQjDvnwBGQ8R3LfjKZn+JmiwLqFKmPSLlg22Cwiw
Xg+sAyxBYRRdz3EOR9ewAeI7tFnx6RLB35I83y/jRgnQg8cxjrwwcOdbVuxv05A4
rU5yl4m4zFlMKVtAlveFuuXDDSRpchHaTqPBtHM0oYegZvaXAIOI1UQku63xq6rR
a3hRAvJNcUbsVu7GHbmebNRLxwP61R+LxsdM8voXDVCFNYEL516qKMWXpMPLiLk/
jZY+9CWsOFiTQHQT17/hJQnwU7FPsBK2i6c72WFe+IPV10z8pf474o3yeCrboTcf
YorAP3QbX3Sg5JDhEHXXHnbB635gsRCv+DUkvaTTq8HfbhDrx+RMCHOZtYiG82YA
K+5xOtPgUUGrD3s9XScXYsZ5avmNGBTkS+aHT3DL/92uWP9AO9aXHvgDPGk3al+K
l0Igb3vCYK2ozhoG+zoWRN1fnLc1nVGedwl/dnrJt3jay6aJeUmi9/1Qimq2d15N
seHWCFvyQZz4W0uyoom1GMPxBnqp9lprRRRb7wgeoIie4oABwv/Udo3QYtI9UeR9
aHDmN1GthQDUClQhT4xJQP9HILa0PBgWG9a/OdFFtlpf7tpbxv1SH4SdDI3YwQa0
u53RirL2yUI1RcjVvMQ+daMZjMx3hwdBW0e3rYedL00DhEUf8i7MKNlyLDZ36nUR
XpUv2aRoJL0zoG4ld7KLNuJm5GEL5WYQtW4qgg3mmfMCoZXk8HIXIgB/EH+d3j/z
HYPf8S3Y3/cCj3V1y6q1uKGGcuVuRzFfg+D61PGMxFkq5HOFXNBH4wmDHluaz1sr
jVKc74Opqsmj7miMkhJF+vJEuiFyUB1RcV4iUIof8MDxyOVr3BqTP1Ukjj6bAkfd
Jd5GPDWPEf+UizkIN097yKWTaMsOq6ygo1N+MK78xthDEtbzBAoUGBVXoGVy4Ro/
HS0krIhGNY9qxDozK/RmBhJudDjYvTzS5DhX526UMBbkhR7vPHqohTjiwghLqAxE
8Gp8BBW7yw/h8WVxh/xZMZEtnGyoZ82L0frm9GXlr9eXqBLIs+XfhhAFjjNpZws8
UXu2yBv/8AhinG2xwN0ULsQwlhtWuZ3+ajQYHH4TID9dV8sF/EbhJs7YRdioLoaU
yn1ckVbJeLOxH73zc/fELh6Egn49T3jIPhoe8SfmIb2iSopZiv0Ur2BvDWPMVHsm
0N1TfPRqaeODEwMtasKSPKp/e9amWZFke0hPURfpAPgE9vTn4YHB0Aj94UpFtwDD
f6k/5mjNByh1XnpQ3Aufcy8b2dkylkls5nWOQ+8W3BwI9sNrXYHkxlmXwxVUBlaV
Buy42y2NGYz890vzKbZJUBEV2Nfvxhgl8/bUcsBPUEMOeQ3OZ3yLIbuUWpxhEIAh
zbvtGz+uiTGFFN/2tVMlUKoFrZdGDs0Mi4uRmEblqFgwNND1fgiYYkBXhjSQH4x4
0aXBvY/RT6oURXevs3OulWPsllRuoUT/cEnXPngIkW5laJPnYOoYKZgJ/dT1y7uX
ura3C6RveUIR0S+oE++E57zJtQph1Bc79x6DGhvN3yPErKL7zvFO8ph25nIVQomM
AUoqM86gP+20KnNdqcdT+M8/qCLKXCaXa9OoehUs7jlNUw08k64WqUma45US1ty0
pe1oFYxGLxHwkzj7gLmUkFIAaUs8EYKCY22aIJEpIG7gMgrrmm2PNI+BzW/Upc4W
ED9aieSLM8JxJpMRO2icRHXmWP8ZxR4JxQMfrknb5gyJt+nmPP0379sSo6ZPlvQ7
gCZGApxcygU/lLSWGaJYoojDFyl77ZgsejXU3lSJIAf2y5zpbbKRgeLBJu/u+/04
H+bRY4lWINdsIQn62gDMVxmfbLxoD+LULk8hPZTwcbEsFYdlqnTJk+HXR+LZfsQL
bvMupoDZYs6j/Ao3wdz4E2uR7LCPDiz98nnyxxZs012KGo8/ePEPu2o8spDIdeig
dHqR9obwoy1cHq7tG/OLUBUjmUfWH5QYElSh7qSURbE6vzF8ZyLVucZqNGZqY5ZE
LikRxMA7s65/cB/wTK42+71sNi4yM4MLGeH3zPb1PHm0uH528sBKb9OHE6bav8He
dzK/TXuZnZD3/ytLXbs6zk+FneahLdXFS1JpZF5xOfzhm61QWDkLU9GQcHpAQNpR
yhYu7HdZ5aserVPDMMZz3mrLuUKmnIhaSuxYdofH49mP911tQOFfwGos9uQ10hVW
To2Q4D5k0ZHgAoYrWdD2wxxND4BChhGM7tJmBWcUfOb58lrh+qWjbwWylD6id3kY
tYn1QaHCLsLQGrMljj2O1obDWBLgWjqzWfnFB5zK1a/cncLqBAQZpxzjYpyFK86k
huVrnwq24ft7vwchS+W8fM65bYaIym+mNaN4Rn++jyYxRkvPxmJQzX9e9CzbEOp/
tkhNxVcB4R803YzX/VMAEeo5Ha42ZjoVuQpk9lzJ96AH3fWFgNqTZupD1el5Wt+C
tohCeKj2OyA5VdobumIFaOPVkdUjFFHnXobAJ9W3cl9DKzaWyDpEHwHDLnPZ1gU1
F1L1Acie5UxLx+Io4lXc00+FGuMdqMlrqOIeQAqJOuhTOegDfQyFWfWZsBzAy037
s6ip1jCXGp7FNXbJy/iIset5WREhHzrFRi+EMwZOc4750XP25IGLbSPlfufraANk
g1Axkm3GF/b7MTR6qo2QSLYFz8eftgdQX+fTDsoYSOUOVe9sGlsLQmx1+FhZ/vmw
QE1sTDBlIoagTAHVUJNn+/zkrMbDOd3RpizH6XrpQyVdqZARbbDK+/19OefxG3J4
BtvQH0gZUBwRFg6vbd/BqvGuwrBv7SDo3QshvjdJmAoiyH8WWWPe9yk5jc+pdk0Z
o7B65Clby0zhMtJVussV2aCUDYZcqzCQ6s5XJGV3GKoPMa+U9+rOZIG1VTf42u/j
JF1RCOtcTZlM7EFpA9R3GZy3qGLu5rdClKa+3nltwj+2PKVPBOeraSEQ5Z3Ko/CR
QqAKeDuZpq0NQBXgB6mP3iABNdJdKbxNsMHeSRGykMTxwL3WdIdD3tMpxVr6Kub5
ZNeTTXmexwsmYbbsHayFF5UBut+uA3dfurkwEERvZInnIJ/2nxt9VvT0kjPKBfJc
7ifzfeK19mlAnhGmSg0+/PeYivpQ4Wq4434z1A7Q+TSCDec5u+H6nG1Gj811KT4o
+0pbXYuHgYJYyX5/bpsHm+gQ+psOAOF5KcVVKMyAeU1Tuv2XwYhE+yU3A2VtSiAY
HUvmKtbXOTLe6J9Pkf5PeQhWP/u/m1OsyPRCNpza6aewfRlILOmzZRSL/QOzUbzH
QpLPLvJNuyk8/6Oglfoc3EKn+Mqbn15Q8UgsYob3Fh+3B1xS0FaT/XyDXZ3nuSLU
A+ZfGgUiXXiSLWhZlwjPttGFvUW38+EXBTP/cs8O78x1m+29NU7UZ5Ft+Jrv8ddf
KAdeI5t44q/Tw1jGNz9BS7qFGWpAky9NnL6ub3ba1VxvPO3NrrmkrBDrbbKyby3c
K2/lVRP+8oElxl9LK13anueXSr+yx/IPJ0FdwlT7swBh2Fd0IeNJduI3aSJwW4IK
O19r7DutYLtSHXKanO8f/kLoHCLojgrYMWYOcmW7PmqS2LjeF35Ue0pbkhDwH2ep
TsUAsqXFiNwUWi9GcoKkmbnN+KAOYrQR6/KqDEq3rFtIfH6eJqB7kNOU+YEC4biB
nyQRVB8mZ8mGm+pJTyv3HO0eJoxzjesRkSvhCU9jygd8zksq10aAqlBjRsdOBOqP
TIV1vxNVc5FPVOIXs4DgTSET6OiXkzpbOt7ie6KpLa57i2lziMpd9fg+dS25VQD8
bTUo6Thotq/N3rOzWgtDLFcqJeGzuYKsRdcsoUXNOjVyGAJli4ZPbFL1I68N1/tC
qeCH169yShkjNTTXO+4S7rnEbQo9Hon8eDtu8rofafInQgQT9TWkAwLNIA1QDZjF
rA6y7K5X7Zel/BCHLUw+b0rp6twlvJsywKJxnqFNaxZx4YZlizQIYUZxoqD2OLhI
2Irs3xhb3A33hhYfy2SMOcyk+o8suFLW/JYbm8/1DWJRj6EiOP+IN3OoX+hjm9GF
pBPChQfplUzUv45K8fs+52SsHyHNzWXMqB6yDNgYm+ARbRYNUaLABWElx0Dm7rWc
bJfgvsUBzsr3lX9Aoe0aB6J5kJ1xjKGaDHYlWGNYOEWtr/VxrtocpOkpk+2xUwYk
bYJfmDBReE9/fAdAbQj+3n8tjvudQV6DiRF0SJXAo+Y3U1f//hfI7Z0VklPmsRBg
Q6ooHNxjt01y5jltqWkDJ1b7Vuv0vgL/DKpbmrsu3kQ2zMdSeP1MhrGLxB2DAvhz
MieYQsA02LGfKyWTCvjDTzGMhtcUtihvqo11Fc1YVj3kx2xlD4UF59A7KKZW2dal
R0J/QoyvbYrvwlO0PMS0vD9m/NYJ35YE6PDdy5FkD/p8Y9kYO09SRclDzDf6Zr5d
qX/p+QFSCsEcDfZccXud0CYupmU/DbXd2S12qxwU4+42/cYwkjgKWimLnNcz0K0Y
w14FttgGP6UnpUwMQyrzVOr29vRHtzWnAkbqSQM0RsQ6d6f2hB/Y6/7RFHHdtuxU
5N/ZeLqtMhqeRUbyJ53b6Qc47Phid2LRJhFAenDe0AcQQwEykS/RvZc38KzMRW3A
RjQMS2kuHQKO0rkHN5APNvHLtxQf5EQR2yv0zjTFZU9qf7vrhsjvFyZqhwEAGLXt
9hOt5DUSf0/9fzOtTHCywinmQ5GJqV5zjk+L6xq9D4zanhFvCpVIa+b5VGWqWJnb
ZF7q4moBgw4i607Lts1IJQ1Q+C4kKOJ3S5ksaKgylxdNzooKh3jtrTq5vQd/Q/q6
YavouZBdlWIv5Yui49/NPHE/v4vQEwl+mbXGNyISP2fpXMmg+aqgfuw8t6j7Cko6
HrQKGunj53U46EhoEFeqWcOENZHrBd/l5bFXbHH7sbi0T0lVW/yYMxjBJqEHerjx
IdDE00kNBkL6ZgnQZFHFLTjGfrtqKntsvBdwBe8k+/cPUomtHxoW3JbQLbx0TnV9
EA+++wYi+WSg/WNYASHm96EyJ+W2BXZpIjX+v9I058cNRXVxetoU81Zv94z8OvOF
kX8l423a+V9t6Zg3D3O+8X26A/zeLVw6KoIUJ3CTJ3AwyK5BevtxT8wAiKBYBvHS
5RZb7sO1Au4Ie8Y+4VqNcdVWETIIehZHTCzRt7WBQ+Yf03IUz5Ovs+YTH7k7KUWL
gFhHQKkViVu6TQhBIyDhhKpr5vcBd6IYXm/YHL5+GXONNEH0anOkWqe+ZadjIcfX
eX2PQPUb2QTB0Ae028cjng5Oyn7jq1Gno0hBHyUAX0cxW9RweN+SyuTjREM/Mw3L
mlM3+MQFqP/KC9BhzAe+h22eLOh3tr/jNyLMbxUKFYmLhcmNJ5tMpRKzmes3rIWQ
DsC31OzzOfvA2j0sxgQNfxOiPBMovs4MMs+Uly2Vwsc7qhHG3y36fvW7yoc5awnR
GQslxtTXfPsto1EL1xKPCJ83OONmXfAMsVQCErU6KsAtV/A8RUSYfnEQsQfMj1Y8
pQcyRlXyh0ZUOsm7KzuN8it4YLkRNHtGrkA4rl/iN2DYMaux9hSI+sJYCIbvqJbs
sqT7ZpR/OQd6iTsa2TYsshugO3nj9CN107uJxj/kBkyHtj1jO/wZS5ek5cDj4z2F
5mfUP/rjN5wu/NQpqDH+3R1PqXvPPNUkvRb7SNaKLkplU8KpwbKtzCYRicP14AM4
HDavvQy822dnpa5Aq93amray23MHMnxRdWQe1tKN68X5ynLuvqIMHBPbUfdOJWma
LPQ7b2H1ZUF43cXYHiN3NgkY2sFHWGk/A2pkZU/r7LLNzPHYkLczrKhVApHJ8mTv
JQIIYVNyduKuLzzoWjoqdG7MbXdhkfKuxXmEz5EaOCh0Ned0/k6VPzluiGPNcRR6
Dr7OBoEpvZvw9NjWftyItrGiADi+iUToOW6Y0YrbfvIKIlCy2LmXIVIcG+KoppKZ
RcoMx9lK6Kxs8LO7Ply9MDfcuqoktKlXQ/YfzEsjC5+QbAavpEs4tMqkr6lIH1qQ
44V77Ef0EUkzUWjaknoLTLswIr6Lb0dDzd0kfe5eLToNSnNnqZAAkyjt2JoMetg6
75NMDUfKpnbH267pvmvqNQ4EOefmIfLmUsxE082PfgZXNptUV9p91GgSGwqlfJMW
PD94kNjt+4qQ8KKFWQZ0Tj1F5EUHcQ08g6vMThtIaEg++X+WOArooJyF5hMExgml
srMY5ZsQO3yqnl1UNtzK5oKS8LfhKfrjqlDbV2gEssz5sOXJTpC3dTJcUn5dDGru
e5AWMwZbrrXUcYR7s7rDbk/T3l+P7IAbbVV2s6/YEdB1u9jPNKHjH6kqlWDhj8k3
FKmho7YHJ4fNQmT5Pnn5Qlo7f8WaPFYDEig8YdVKXtWPQ9KE60sYMDClQsqB0doM
H+gh5my9gQkU+JwSZy5gM2WnRHMvsm2TzBH9XuPqWMTk/p+KvNomoyg0TgCuLEyX
Iegndws0unv1NoJkTg3tVkFuK/nrvY7gqI+OiHNaEvsbYFuZuw7OdXqjJxX+wgQm
0O/znpFMIgY3gVxllD35rXNjf6lLaTPVeVeRZhs7TfiZcSLW7Chnxd8UZ0qcbUaP
pqEheKzF/3SXX6kAIXSfdSMJWILx9dRg7IQ6hpxufD+HRYA3L2s+8CKxIZSwgydX
UdRD9ruzr2z6HkfbM+JIRmBYb7DHGAEyjhVN3+o99IocjhIOxEJ4DlvnoxOW4rNQ
D4udz2jpVocK4oJYjYuDD72eN/mb7nY0xEjgoa1umoZ6c7JMgIK+uyvzAf9gBgv1
FZjoBjhN2QcYNS15bDjl2Ryh0fJW4KcPvycDZk+ii7ThLfMDzbvutvTi7a2olPtE
ojR7mrcWMwGUdraB5TASYJz84iJYWBx+T2MRvVHuliwzI+QZrGiWpUPrP61xacC/
GvgbamLx37i3QZZgXAEMLWEWSBcS0kTlEtYxjriX2IfnfaYeNsrULG9XwGlBlFl/
9HfViAKQTCOH+MVdHa2wJIjcGYFrQJ/SnJ4GK53pLuEris56fI2pbap/8kArlIF+
zoGuxAX8F6iLWGJZWztvR3p2EStAjSBc2zqeynFVXSpld3xy4nvo695CEMF0DQN8
ofbJRyy+0pjq/PzNQa2hp/z/TKFBWfdkHi3gAgADX2tw5GZlDMaowCVOdAbf5601
kPMstnJ0wQlbGSD+jo2U6ORt9k7qK7UlLC5hXYEkjAgW4pGSwvq7/+Vp8WXof39L
jqbGvHYOTmIo72vnkmxTMVACeghmYUCyZP+UMkTMQfb8MpU1sxr9t7SLwFOVjQWO
GuPxLDwo1NDl2q2I8y8e7FHXxYxL+NckPV+rQT7LGOcs9AC+AwYitCFlajm0iRp5
QhOteWLvI4kyBYrEbWgDloK6xX1QTajKJDMvxvUJAHdWORGmU8+O3FTdo2hPq94e
1GASmgHcEe7RTsuo0+8oEA6WLPq7RDExffwIrHvkqEEeXdNr2OLVJHYzrPXj/JHq
+rfgtuiYUMCji+kbm2dmr/n6NHZiic9hoJ6TkgXYHSz6/P4/io7sIIKZwkgA2Blp
grdcLuJNSm1LL1RJYk+JES7t5VAqG2ZfG+ASxMBO/p3WbGn50mOuGaDzFly/4pdR
QZIuL7ep/WxkHq33H6J2Ny0L4OfOGL09uVSMntq1ztNiGJleMRquUBcgeCnk41ZD
wWOmKkiXPjzEubIrV8Q/9JyBHXkPpNGyJG3T9exEfPd08i0/G6PL+VLsQ1/Kbtoz
GyqVcPPS3J8uta/LPmVcAwtoTVVgCTW2nGa5zZtkYwvHI8k+BUZ9BWRNkUsaectq
UXMS6PIP1kAHN1emfO4UclB8+gKqMKiPfy8ZkY5u5TS5u49lPDdj0mbvW1/fpvhR
hqhRPoxNZxMz202R9abrPi8D2sudIdSivi7M+EIzlTWp2LiZoc8D7kJ9vpVFNErG
nFUbMkUESOBVMcvc/hFep/hf+iil5FiCxro6aPB2rOymyRKqMwqhPkMAXWNWhpOz
Wo0fwHkTvoQ2EU0aiwU8RiYoXDIFzRJZtad6EiWIFtUXYJB1mN9Thm6uiJQVcytz
AnsD9zVRXB9C3uuQZVBDd4YyW0m9WkN7hMLXuIG14T//L9bQ+4MRdA8W/9co8PUx
mAJ/kA1EUJzs37ObBk6TI2VKwxI2guQwCKAaxWReGz0M4GHLDUBeiQ/1sILzhlr/
AikphV3iAmEcI9v3GsnyimWK0tgSF+p0TaXLOZZAynNDtRgyUJ+kC+HL/YyVPO65
7y6ivACXjlbhEDTWDMj93TvfflORqkp1zcvaS6iP4xlx4QXEvVGpkdu7M3dANXXN
EbTZCdvMdDszzeyITzVEYouPhEdR/dMocuzTkzdf0R6ftSGrg6Svnzxdd0QNNN8V
LNioAJD3y4ffxbuHakzcAQSkOpLF+uggs6ZYFkflCUjIXXwMESGK14lqgFM/NBh7
nlPFkd38Xsb7bcTjjm6mVDjWDrR0PhULq9p2Rvd88d2ubMFLJujcbu+uJ15Dfmqq
YqRl0dgQ5b+SX5/kL00raxUogtvRDhulIFNYXzdBTf6aC9SCOG+DgdljDASIvZcO
jQN/pxZCZvWFFGGmxs4TYA4yPnID1nz8fZx5CiKRnBPr9M2sNNVl+G5+wxtB5XVF
hGhVujYX3GDGlJKxMVlbBBPsqCp8bVxo2LGDfnpKup8YB6ELMGvMnxbbNwXte44N
VjUh1nRan/eK35Y3JPcR2mgcqV5VBPqZeWun/RTP3dWXAqq/2TYAmDLZ+YBgZYWm
8wGYIfCAYrUmpgCYHcjo06Sf73mSzM7PAZro4iMadKhkXtfEV6lmf+uhhzmA+RKm
ySi1OPFPaYEzAgoqDZF1Eb9Wdoq3++I36QaflO78bO4MPuR0HfpAKAeEC5vQ9kFE
DK6O4rVjaEiPbpeD3Halo4Ye9QLtd6ja0WtYxgmCS9dFcqtJOqdLJUZt1N1AqKVG
iv3YSt95Hq1wSm6SWZwJX5nNvLnivhkwzE8oVKK57MrEoip6m7cdccDPdWo2KDgT
WiidORJqW5PWUaHi7a89LUOD0tfsHgDqFs3tRJmg7nwq2KnWqquAzO8+J56A5fpI
Sn6QpQnYkuqscUmNsSbU9x7+ibNkJQ2Z7+j7DTDFmioiP+GCwnWITi1Eru0Qtw52
3jW9I+gSrAIp9P48aRv4m9XHNIKFhgEwzlM8SZEreAsMTjlXaLMvtWqlJt9tyma2
vK8T78ApTWhEaj3BERfu7De1wRjqpktHos/YzCurgxOE/4MTk/b95NblKRQU52zc
pUxwiBovSxTo7t3MQZHnylHBmeUyrtb/O9MhNOrpO64imK2vtgvHaAugsMXd4Biq
T2usCWvb2sqtIv3IcqGMBIfQoBqyIpf3sdySqHKiSbSITou0dNF4B1QUoaG+wdsP
IbII/bAs4F6sEVSuc3Wx7G3tlOfIRF+hXMqsOFL/+W9QeG53F4G99l9KpQ/YBDnN
colG5Tt1C9nzn71aZWsbFKQpLq2MxndgaHKSh9ey5KOCwNNBpZkGKQe8MhNigE8a
ieF+pwnIicfo7g8reESKFJKWjd/D9m67PbBjhbqdS+wPecni51XT0dnfu40J9wxA
K8/QLiCnJD9ICtyTs3mpLK48IzUeY8OpgP5rViwZ8w8fidHYecgnaIxxdL651/cP
Bcd1w4nZummsq5DlthuVcl5mynqeo9C5Y5PrmSpFQBcCkNeaCaLlSx4NaiFieXa1
8ttyAqh4PVGlU8OulQuAFv6vIoxsbSd3J5r8wnqt0pUCGmMkfucY/8f7m7O35jue
P45t+GjzZw0Ci5QkVcK9PWFkTVUoHrBsNd1wq8WQ1hfMGdWSRfUZrZ8JSXl6LLPd
XcFBplqbHM0qW1MpYegGfvMEvZrVLpQUygZNWzDo4GiEE8NqVx0wACQPTExNsxFG
HwjPNjrcL7rF+HZ14vSezxlG2xSIfKQGrf/YGQ3DCj4UYChIJoV7p0utpzyQtbs/
AgvDd5Lr5wr5/k3XvH2up7LSIn327xd2J2NEIcfPVlxqc0ImcMQPHbTz94M8jorz
TsPrpxEef63XykBjhd83x6uDRRO6B01ZuGyl7PAt+oaleZrzD0WLWwolaJLUWPmy
jLyoYzZTl56E3RRTHshvGo6AEvGhgXQpRspEB/IoI0Qq58a4dz29jtWD9U17vhrg
YezDfy4kEGMpgC+m4BeHbxZiS6y7TXIb2A10KImUXR1SXm5eYlWHBXOBu/ntqqH2
cwtNqQnVKE9dkzt/t9dw0tr4sDst3WpiVMskzP9aRN4JfrDzDHoQ1CE2g/km5v+w
ah5XLdGBh5heJjkQdJKsHwexPMfSDJVkNUse7K/0/hiQZiHOvtoRiGxUPYXdyYQn
lDA1PyPrEG7kM1UNHxVBXABaE+H5ABC5L7DnsBAUUm0mrbuf1PJz3nG3UZ7AdL8h
KXxJT2OMf2YTG3R9Had2DEvXE6S7SypKI9Lc/uUoEaLuSIIzR9+K0nw/KP3D/zVL
gmLZELFZ+/mTplzuJLLaurzOcpXoKeX6Uq2+syHLDHikIlXQXDU6TZ8TQCKJ64Q7
ynJApQ3rwBMiDpI/AWThzIxaQnMemFJRefQLT3oe62s/PsX7s/3IYhPXEdNHpMsI
ts+7XMhNRCQ2um7V79TYFmiPR5V0hF4ybzogfCW6SgeOuwdEm58AvZSebeVmiNal
8RtMjO7ZswJjulywixq+VMANc2UDm50uJE3fzHYnhjXvAhKfCbQYmw48xrmKGX2x
zc82A1OwFgqibvpkB/0AAWYHlG/c2f8EOD5B8NNd6ACH4r33LTugCrNYtUdU68bV
S6hLHOZOrlmmeCI77OYMLKo+e6WxdY95lJAZKN+lyMsl07GFIJ/Voq3rGzKrB9gp
Ks2h7q8zl0Hll947UOkmtYn2puzEg5Q0HHVkjOjMuyYD0MEBHhvss3F39pHoeDPw
a2CG24BfflvYgW80F8z+9cHw1b9/Fg3qk1b0+OHpEgGw5FgOH2X8YsXhXCEs+dVQ
qvWWBpBH2oFoWCaD0UdAIQ64Wk/RbWm/9k/fkrOMxx2BQu9kyWoe6rdGzpmOCmfR
Pus6HLRwAAuEBjZWFIkErSvRW46f+fyQQqEGBxwdCQOGWneo/wKtbJ7AfS05YtD1
yT3lCdLTHA5dTp8haqe5phNOHKumWHKptGI+k45DUe0kEfIA4t8jYOIFSDcFQObv
zfCGt36mSfFqhrz8AFjvXff5NkimIZfrXT6efMeMdrtG38BWLCWxBU0lqe7a3qR3
TBU9JMpMXK5/oUhAHXZ8LQ9erMrvhBeuWAkQFFknVaJcd8e5rRrbUZXR6+UXlS4I
0b50pu70BiBg881SAmgjNwnOTkx7opG0lfymt2rTKyV/IfH6o1Wb9qVlXPnpjrvM
zqD+kP0UmKp/mdurdI9V7M7Yj5z4/UIKfq4xo0+akANj+lEQ0uymhbukGI0i4po/
RH+pFdDuYtowiLAhVPhECDAL5H8xDPsnb+75dHG0/zOz6flnYO99PSnDVTc9r35G
zh7McRvlrfmz98tTy/yIzydYGjwbHDZymUgGdmirQScybQY4sI9Nuf7+fIqDgHcL
cXKTDKSj6lrwnI+F+UrAXzBj0CACFtWwzw0/4RC25U8e95mCakDqbtKONN6QAgDf
buLRzT4/q57z1PCRr3Af1YKCjsBEncqzi5bhEHHozE2w9AlL7pe9iqQrFG48iDo2
MMTRnkS+hdL1TQxW/zeEJQSq+QcrPyeuax7IwzCjoLybYbIjudxamTy8MjQnjrZh
2d94+t6ob6o3NMyH4g498zvWENC4/ZrsEiC0IBlRr+coE7Rp8w/Ozzp6JA38pQ/R
c74VdoZoWPl40vnjQtgFtrkJUNfE2bPItNc/kLPm0MQH0CreHsb82S+iyhgKdjar
tO7tPlPTNM+R12qs2qaIfl+VLw11S/njR+nbwtwICLVVYFx0jbVLimdHQiYqvMW8
8j+/OlbSZp6OY3RFAiqwC5zWpuEjJFVe1O1o9GkQlDAy17t5/fZDaH3PLkERGJ5N
3kn6K8WF3bdyE2VdQoXOKntVxxUZaqzBNldbeZWRrCQsfDUEehszkN4g+SrX+MEw
rCvCpOHgySdPN/Eb5jZ9qMLMCnAnQGJAHKsbrR1CVZcuCmEeDVxAoABxJNep6fZd
YvX93loMnVP8QLWW0ACFdNEE3kAO90MVNOskqmnF7a6wCSSwnpVOxn6w9y2o95fJ
kksarDLUDCi6d1uMfJRdU6dgcCGU7rru2BHJkP1notTEjuz2c2ICSZktB6oohddC
hakRpwE00s0rtYUGBJwRSsaS5NRDorNeg2jNveCIPIVjEQM5Ikb+zfzRd+/3fPGh
vk7Ph5Ji8QimGzKkO3FbhbsMY+WxIXrBX+geSDtgVCdzPAADRoujsng8AdUmqazw
uegzadOctNKQNHof5j2isNmbSm5GEutsnyVlhlavrJjlIvTxQdcBIp+AB+U/B+El
q054l50c/7H9Aj7+hSMrUqrn9mBGhgObG1XIhknRsw828+ejVV3mbwQk5ONm/Qp0
qeAFEpRh8ZJikBnKykXfTOxbS0B8smZLFiQioRC00R1wqUaktJ2X1OvTeB1ksiz0
UUW730QezBnbDB9P7sxOiMnHkTQWT7KlrbaAJJ0Qp3lzGUHjVo7l+fjyghAeK1kF
tlB765BeS5fcJfOVJFBe3ivS0qPXT4vkiyvU24HE1dUG0C2Nu3VyjwUvFO137wlJ
L75HbJGjw3hhL4zC6byrCKCNd9GYnaeYupmwy21ymn6kgic+M9P6zwYWhzRY1rrt
yT/5N8WfXA3GD8ntDlhj9oBaGIsvT9LEdktlE88L4qYgbYs2iLSX08hrdsiCBoI/
iKXFIkOhaXd5dG4LStuSQ/Mz8nmEqnk3ZyUMcwHYJb9EWiJjdsZavsQwlmeexT7S
P/dUSRbTqChccMvVzH09gHP+wN3dm7FP95VfnyGyVZkY78RtyN1Fivr55+iSqGnb
WEbYZyisEgyaO6eMocyQZsLHTRgw2vSKhgf+7qq4pBDd9DKQQT+cftb9avo71VX/
+vRjqLUua8gScT8nAlHnGteeWSYywr6Xi5RWMQnueQI/V1m1nBvJAaWQovfn8dWF
XN1DNDDNowO4Yq+B+zw/JFgB55Pvm1CYXPQ0I9Cwmr4mmHVw7Ed6841GZalEghMl
3B62nCXNciKZk5RGay/nqBOc2tmz1Mk5Kbg/2N2dva+dJ+0a7QZvsTEcO5PeYLWQ
25bhQW0n8pjmLR7X1w65zxccVO5BSEl4feI2cl9W7edJy4fC/IhQPX6jHKmL2vvq
3YB3gpWFkWOiZwzVKkRgvk69ghjIZ5JpZXVyhZT0l4FRuxf4TZTZFcPX+kZubzUM
YDO9apUMlzJncjBUjoOT6+9pQVzMD4YYclLS2+8yBzBiIUH2dsfBHAi286N1dM9B
/+YPMobbNEheF9Gci4LZQF7rf/G7K6zIf3h/1ZFqPZ/VHdw66x2MbqZLH1n/m9uN
Sr6OaAtZWUQyq24LbvJZ9fqkWE5J5vnBS6PzhPqXoYn7wJg/vBt9lEr64OsXJW2K
5G5hVZOI77/EREoQ8wNA0lDQsZ3Bg3SazNVjbkyYJeL+2us19QI9lYwLKm9YOO0J
UYh9dhBhnh9uRqMaz1H3N1M5iymbFJgocEJKqw1aeYUmnxnWafxIJXPIVXUpbZZv
w5tZrgu0R6IVWb01HiHhs4B6X1thwPHKzN9UTwQaiMUWVAcErqnK8JbkNhASHSbN
CbqQpP2kOqPnZETdzx+X0dnVrh4gY4S8GDXXCD4TxkJBh8mH8LtTvO26mHIPrAPu
e68A3VMP+SeHcCs+cQdgG86nXeniKLQgI/+6sxQrzHbHrQdozgFaDS9ju9txr6+y
H+Go5tzsTOD1uL/+g1PcyycntDO58SnngUnS/hm6VEYMC+yv4rcSoZY38DKiDflA
teHPVm+yP7lVWvp5dwycOZGX4snS3q3mkOsBxRY4o/XIz0CwCeLH5xtBG3jdjQMR
VCdTt7K7M+nzztmAWcMwZ3DQw8Vtdl65NByYvM9hQIpxQ/xHe6nOdzbf0gYhidSj
Db+ZFHme5IosCGy4oxK2XHUtbCNhngzBt5kSk02nljxEiPUnefD+8qadUwyGqMGH
uIya9JGdj57FNH+BiYdjf3/shU+y0IC27/p+n4HFRSkX32NB4aWZrGw5dnTNmNJg
sljJgjGEWKT38+oPACsNIpM+r73qN7yNa5hqp7efu72nObWzWMx/jAuRyVcgq3sY
roypNsa2TDgNWQSsAhnYGkwI7kWMWiqRQctP4WZn6UjAXgK2U4JIFEFTrmzdCia5
+XvQe3o48JrbUth1zeNmjGMjLQWXlSi8ZCpa67UWSXKXub8NvKiLozyTuy/fjL72
WqHTgkRWJwxcPHPxfUIQoGKEz2Cpf/W67YnZjhHg5m44nr0nY2pps+Zcvow5vvqo
ETahFHnmyrOWGF8mg+qTO1C81p7SlpshpFt5CSfbc7YsgP2tllDE955OQVlFMv3R
o+2gcBp7ZcTufiX2FMVEjckPFheWI9HLIV+2LPGy5tl0qjmQpb/wcyhfk+6c8FCk
a00oDTwmdP+AGueGEaWPA4GODAeqwYYIcXvs09Sp2L4OJ8ZgSwpVPHdF2wdhfbua
Qz1x82GwsBhpynN2vJ2M37BRfvho7njCQ1lOk4FUJCfuVOBall5K4a/31PhUEpwP
nuUE+RnM+Cwbg/w6cZipMYDTzl6cKUlg7M4e5o+1YZz2cbG4Tn1whOJtiGlC2Eiy
bS7xU4/8MXTIuJ3RMCw4uIlWG2S7fZoolIy7owpbDB2H9+Wt9MX3PM5HftxP30GB
zMm8yDQ5F2L3ZJtC/wAvgiRCi1G5j0D9WwhGzJj9QOO67dFI4+XmWauoLC6zUiHk
6mqxM1AhCP14/7a74Ks9mYPFriTcqGSjR47G8O6lNWLcj03+8SGFDvB0YWK5qXwb
UMvgYDt5kN6z1EznZFRwvjIwDboS3wFf0p46aaWBe1tTvvJkAYpLEBsvFbE18tMY
cCFtkG3A+2+ADsF1j8dlRzJwMt11xQeUoZZchY6CpLtG5Ue3MTJFjnfiXFyT6pO6
Ou7c+wTGAhJF2tjbKeyL62ff+nPF5R29TmWF0Ol1zLtnCFKglaGMHRD6kfrfI5Wf
EIfe/VnkLId/KjR/xJ7A0SSyH17RBO4cblqBWRowS5IySO4b1D2+0E6IOFVNlTqj
jHsKoHuchT0pPMXQJ6pb6Xs+qbSNTanOOTBFxyZx41XWU9ABkWFv37XnHACCqdMO
tFABslIT5F25QF2fl6A+dE4TrskG7tmjUyDxiVPXRcFDOawx13KLYwLQdBOo57uc
CUABzhhH3XT6NPRrduyeLldjz4aivMqBHwJaw6BIHlkiCzRQwzaA2fBgBbRb91Nq
/NZEl0ovPc3YBx7omuakjejyK2+fSGgM1S4xvHbeRx3gXjFz7cfCOTMJzZzzDBqm
iIYzhS/tdum40I+Y+6BlkJOR+m01wINmAwRq9kc6LtKVWh3w0rsNvAcY3UWN7RSV
BJbG0I0xbf+1ta50O7ekNZkZR9ehnAAmdON6V4zLcGecILhAfJs2atmzDDrJ3CAN
LoViCE/NHR0NOGP+I4gfUhgjIcR3Gf31Hipr0bWOovs7IS2jFUGNVvBLqfndrrB2
7QJXsjZYXrQORfZ4+0YThzTwVunklUSNTpu5qpFy5awSGDIJKHz523uNrWXTt6IJ
2F+aYtod335YQn2giB6YpD4f6BlrIpGymbQi2JQBgABhG0Ee+b5zch8576wANu4E
WQknJAGbY5Z/7ktA+LRWjMLPrkj5NtQEBaqF0pDudFc65NZe251N/MHVKO9D4Pxb
meMp87WDljxLhhDq6tj1Ep/MWMkZ2bsFX8b4N2JKuBB0cIjRykP8XE0NH9J+k/KH
IguoH8oD9jwMapWgVoaBPxfWIDd9rXVMU6RIMEhfGH5vBQoy1b6+SGrrkGTyrcIZ
I+MG8+y8onQqv2ydSjhxmJ2VIGrPmuZlTkaTO4sZEIuOQO4PHBp8aad5KJ0MBa/H
abc1o+YBfzbTnwdD9XD2u9uAGlmBxLAH82lfS8AN0nGbqLAFDkuPRaiJ0MwcE1LO
qQTlONLqFZZ2phUdFYO4UdREMiDIrZuD0BsyJQ0dXArhl2mkZbNSKV6ATGkGD3Q3
hDi/gL6e8kG2GBJlC9Gu335lHkBYZFxBVELBKGMojNwD5uWZnCrQ+nsgzpp+Hmwd
m7+cIdTtuUzjngkkAzezyulQ85z3j0HcNbyiCZJ+tvejcCMJ/TUDgbsWNy/3dgSs
6GgpY38ga9xVHsy1QiGdEP0FYH6Yb9Fk4h+7iROgNV4lbrhqpPrKg8fQn4xnxrzr
sm2uRlcN4OtqmgqZgAMWSQC2cj1qgqZon3LJGiwngnPIvTJUgwDi5LpQhKuggWR5
sgZoW5LxyIxOfEXeBkNvODJpFI+XAFIH8woOyl9tFrM0yE3PzggUNBIkdjIgIX73
61o0Kf5RlBGugruCSCb7V4aOr5vLJe/8+9XhwcNJLaTkSchO7VbRWxv0j0s78Cmv
UT08ZloBZz/+Z/fbcXzFb8VdsZ9XwpfYJyAj2o7N654aDSLgv1Hb1V2fONI04/NG
YEIuEDOWF2heqwG5q51it6xXqgDpUZ9VFRZpjPfwxTko/BoENR0dcmjmzDZEiJCA
yR5RsvKTuYGaLcjcm4sam7cRfNGVOdEigttDij++96U0lUIbc6KgLkAVqy9q2n1T
3gn3m+8e4ov5KWxihiTVS7ddrUf0WuTZJSV/0V5k/Dipc5/luyjoGjP69jgQFkE3
DQOsVjZ6HOHt+6iy5oIpmf0TBaDjK/nSvUWfF/NzBDaIOkjo1Bv9jjOzvX/DBxDE
Dqxbf1SQh6um7Rdga4qD3wvzAgT1bUNAgnWIs/oRMIyPHasn1zsBMafCynlhC3gM
RC9sru4f3EEY3yRAR+d+AtUM0zJqKSr7OhA79uTzztQHvkjG8ZLgN+xUUn6+Eodb
IOjILHn47AQ78Ha2ezf0w3sTmt1dwW3BRgnq3e/OYbZVdjVg3hKk6k90e+EgYtCA
/lNp7XVTMyoZBkb+h3gDy+0175jo6kgnetHiJGn0ZZv+XfZWX2PXa6m5U4RCOJx4
ju2E8KlvCQA53MMJhBlkXY9JUC6hXDczVIz82ovcsh3hOyJJy/eO9AhWwkx5uRar
Hqv0Sz5Z9DLKYnWroSxMf/9p+9r6fwHBLdfCOOSrrtC8HDzQke1WIffdbne31Pv3
3NiHkj6464yDIoUpAh16SGaUdux2nGOmwce9T1PWiWaxTJX2vNS9ZGfCoTnTWuzZ
B37596nKaue5XTK8fvBhhHdmlAAcIGUqc6ldBxVY19S2Mh4Lq2DjzvAxs2uqtXzu
MmF7VixbyyZWYYyEVCG4fTl2MGMKVxCr5uGo0pPhMUAuRhwcR9+iWPHCKuMea121
U1Hhi1YzCqagDPaubOqE3JmIjcF6OgxKfE7wvbrDiNCOlriTCnd/WduGHUZcOiG2
hAYH/XJqXPE0l3azsMq7gIGyVD8V+Ib/GOYVPGVNhX66HmtqX+S0C7j8KBk23Z1w
1YXHIlyKgjEoZo/I5rM3iPio83/U/01dEyX+0Czmub6Kp3oIA7zcbxyxGOyamfYA
yDmlraJKxonp0eK1L5FU4ioTM1VZoC1OJZYxoAay3Oj7zkHhS8ctwaA8UPw41GgF
X4OPflOzcyl6cTctkTLjiV/Hn5t1CmNS3yfuMb+5Sqc1sjlodWlmqbN1u6Ng0CBT
AxjLOt/4FxGI+yCwxgJdjLLTO7DzjVu/GY4nMCBdFuop0Qlmqcy2Kf0EPs/XILfh
w4VZIODW+LGSCXqVbxelw9UMpSbf+XWYdZtMJYIxeRPB7oXzBFEHpwv0ZoB7Z7Nm
bTmCfveAheuv3e8zLvihkTQwuK4H3Vhqi2FCsdcPHU8tVWxC11fjviMw90a8sodY
MGoD3Qkun2sDXJ74DBPViEpXGz8R93jnva0nsAEYY6hqfH5caBAG+oo5BPjHC4Jn
X9TW37cFfkUpEZdZB3BVPyeXRdWUhYg8c/9HoHWJKQduHn8J6iXH+vzChwGAYeNg
UejgFGF+a3uZCj1xBAB+vLdmEFFJZ4vJArCuLHMCZePJj0Hn9ZrgZ/dq1IohduoR
FRJgWYowS+ZckDAiWQFcLQOec1eHhisEIWprvhshLj3ah8l6eSaekjBWEvpUNf44
tosUaPura6W3fONxkK/NVzeSrryp8BOvw09sPM5kNrEkWTuntRDKaJwbuEeCb9ss
XYqR6QvZyUAH0JJtoCKLhT9z9DrZX4Mb/dUEEFr7rSRQbllooloQuP0CupBYCGcA
0S3JYByN7Wcbh0zS8b5VNxdm+xzMJfkf40CdiMbeE2sgkCtaXYbeTbf7+qYbh0Qu
yFe43WfB6f3/AG78LDyMPB5eCMoZ9hnEXDVFDJKyjjnX9Nc+/rlI/qwCKRqTNj8w
CzGn+BJ+Q+w5wcMY7MhaIXtr5zMLMQhKbQi0PWaWQDbjLJZxctsCIBj1+S1CIRDQ
vRIiL9/E1vRt1BHE3AM74uLqbQzO3gdtLmeULl56z5PikqyWFQJ3aWXZ14ZuN3MY
aQD++BIHTkca2m3UhNRAAK8xJn705WdPOG3zSJRs2zpWKYZkHjfzgrnZUZJ0XX1s
I2+KgUwEvsqnPZpSWXgjYPl3MCnPZInbJArRdaQNaPIBRHT8owoSvVoZ3PEhnJVd
0IXREa2aA36iNbrhTKGFJ9W74nRp32+Axj5QkOQzyM4oszI5Esd8Vc7EHnfM0r3Z
XTRulfiS+Tp6QvNHw3QbsmOLrOEXntVT4PMzJQbZoFmIgBd8f+gbi03ArfwGWmgp
0tcFiXSi1yQZyp1CmyQ2y/csmR9z+PUBbFrS60RbZiA0Xpl7IJx6k7QvVMrz6aLb
ts62ul6a2WXoZOi5gOR8fYEQCld+7Pqa4oDEeAIx4cVTDEi7ZPTbK6MyjWt1HQpi
lagglUxtOMdGb60OmGDf4ol2McXISyO1KU5ytrpYQJMeK/IsWzofP3Yzhfd3aQVr
UqpKng5x5jUxX8fD64wDA2Ph9zZ0V9jRLEE6RFgVtLQxBmz0Ar+lZXau8CciATCt
RWgrawr5pKwTEPZpXELyLqKkXmldLkiBOq+VXy0qfaqskOqc1RdoD7yFYCOrhKED
iSsVgZPiCFp1cFHQdnxeeN2u/Kos5dkr/K9D9stFmhJZxM9RYZYQWOXcL5qgFQxt
+FD7DxyO+4kiYRY5pH6TAXhaTxko/bkgks9iVpmUeGsqyCCab/QVc+iDKfYPkWlF
wQHowNxSSxxx7rExiD25T8jd/EXK33jL5YfQND0pWo86roXMfro1JLJrXjDjvOWr
fV9wqzQ1ycHncOMuQtna106NHLWmAjtCdIJ9IDNF2ASbM2oT5E7Lf5idIosMIC8/
Zail14W5KYqbhdWWQMLUZQSI1f6OyXooZMP8vnjB2+9bkxlDM4K5UE7P5Rbo00fs
uqCBJFeWIiv/EPRiBcqztuF6Ojoq/SwO18P1V7032QMYo2yc18u9ROEKZ0Iki+JT
R+8UAfdQ8lY5CRAYkGKFQFNa4wmJ0bVlSBsfTl4NfC8zYREkDx3alE56wIX8kDzE
QZvPq/u4pfFKYJlnDz/KZBmM6eegfKeD7YFILVMtY3Qi69bmKCpMR+GQaEWTtLtt
KD86yHMYOH847PwKp+RK/8FfOPbD0ZE6cfeGeyl+8UcqXyDIslwQ6qu7dcX7KEgw
1Hvgn2fvZ3dXolS/WkffFHpp5TrOtcourSmw7ZNv3tvLQfehIm8JjrleeCzAwKC/
5vnhaG9hZ8DbHuyKlBO6y3hBk4ZFWyddrI7+moQwKrqbhDbEzTk9IlUhMNW29MIC
6WVMjUH8KSYRc4rrE/Tuum5iKsU/699SlSWSc1DwoALb4NJ7SdlmCsqk+MEFWeSV
QlPycderyEZBUxtAbtUAEo6Sv5xv5XT7p1WTZEM0gsjDfY0E/lZd1UHObL9F50Xr
rXBDj5Zmi4Z9LJHdLZv6MIVs+TaEVDNA2R0ImpjwxjTbAOOKps0IeZmsAwNQIDMY
v8Gme1qzpSqd21YVbpcXMWbM+TLFG6iDwAiX7ztJzr0zHwuQ0XlIK5/lbdpTjo4P
75x8UtYXDYBB3WdC6DBCrUWq421RnPniHS5rDXVyWoSRcfi9L+Ocw+Dlt5Q7CMut
XVUJPIbdoOyfrTb2sh5I4UM+HcqFzp2+DGo7XYsvrabyvuznf54ko2D0pMw5boyz
9pOmn2FiTyN04mzBui8iqg3tfoQCWfpqPOAV35eBpRDnE0JZ3RnGt6T0LmM8G8p7
+/oeP96Ngv3NzNXIrOQgpL6ISBYGxdBpQm5gYeN6jF9TEHT6kz6KMw0Mj+5DSQJw
JfSf8IrljbZNUIvyhIefGsgfj/eYWk9M5nArkih7LHhfR00XURS8qmLkmzU6lHRJ
995V8YSt0WOodP1Ml4jAwKn1y3vl1k6n9PIIt0o9NTdj6t0XxE3b+oh5a2dCSBmL
/X9/b6DqR6trLbe0VeI5omPAdb4jSyWmuod+ApAmmvVpQs/IykJLEHiW5hroJKrv
zTT1cfrHYJU6OnY4W48tEl3aD5GSxAo5tXJ7WHVsl6Jj5ucEGAKcXdbBqujXLpzD
lMQin3FG1vKkkcvuWx9xgnWL2DQRb1twHKAOJc56IXZVjOYB4c8hn84q24lsiSwG
okyKH2xk3pK5EtiQxKRFSC/Q5xBvLhLPLNhQem/N+VGJY5RDPdDce04aIfYQfBnF
ubPNzeap1eLPSkXwVr0ykhS/GuNQumYlioEUDnco/LJiuyR4uMjdLXVWPyAxLKhE
mwmG0DO4gMkx8V1Esc7juaSXRftStnmbKa3nXRzLmQBet16KOqfCuoZYm+PmgRlt
LPVYW1LTP5Cmyyl2ZQOvXGKpvR242ICQdDP2OFj9GIl34dk/j8FxtJvBmmWX6Rb1
EI2tHqKFXVRu0+xi80DXfU9hFSQW6JGq95pR+X6D2+QAlPbEcwsJV+cBI8WYfTIb
KJXuWol4rxmOAqlpOerujAlP/kSMjsVEShTRZpZ3gTmMECVuqWygGdOKPYUko2vd
12Jcy2MmevzYyf4g6pxN8ZU6fGiCprq20f9Pe4CD64I+i7rl8QXaU2Kw9Geos1Mi
FCZnlfZObmTY0XsNnIY9DAB2VZV4l8cwcPC1j4fUE1rhrH1ZdR0tX5ASlK02zPSB
3eCBJSfIKJNvxSJijk4rMy0m6LMhNQ7FF4vuV0pnPf7cyOu9I27G/Ww6ngfWkrWq
LXbuovl3uqjSWGcf0BE+DRGntZbcp3vieRE2l4r8E2h/GIdQhUJhybqOC/Vt0WMF
83v+sQYRFt4LjWSgxWOisk1TuvLELZxSsJ2FrFQJ42wXdAmGkfw/iJTmDAJBJjTx
ThMX4ebBTuRAj9PJh5tGlNVWJcdQaRJmhRXHlQQSVOBWA10iuuDORUdvdOrh/cjZ
ujEUISPc6x27cwlzlTm+iUAJJ2Dz+CMSl4xJUPS+vRoC6ddGnHhy4aeeo3kDUeg5
mO52b3IHJsgWsHuYxEAebp+p0CgB+P6lWI+VMd31qW+TqHGKt1oe9rgxL4wAlUbC
PJ64ddIMI+QBBacIGsdWT/npGmqlIXSzKeRr68/C0CMZKSEOj9IecEB/70sQrJE5
1QNnCey4jAezg4CcuBN4SwjVzlfPxeove0jWr2YHgFz6j4MI13grn+aZBjFYjsah
j/YaVtfZYalL8loKd0It+NKYPejrB6oJVCeZZFTSWYvz8I40Rc5qDiAnjtrM35R9
7hyS46J5UIoul+fnsaJg0aXCeB58rYnE0PweZfleXSY6TOtaCDxpvk7QEvp6C2uP
nFjFjSmVuf63gkoWg+ZzOp4MUtqx6kLsbg4VK09tm2aNKEC9RaKJe+9VlL1wflu6
Wx9GSEKFr7NwIepavOYFuH1g3mPrSTah8s8ZINhlTYc0JnPAX/EGuO8yn68+pXk8
j1/Ej6DeoZI7DETDE+sD7PAjg4ouctChfSTbygPubWBAKKpbU1Wlf1riEQ4LtqpW
E/SsqdBpn7r8RfJQzwgri6e/bjYnxrB5zNCt2ZRfc/7MCc6IGTRLwfbyjbOwgdkB
63EdmSJiS5BNxgm6XyZaGjlnwuIjQ41xOwiQdgVF5N+mCpIllzwVxZ44zYHI555N
js7DKvM4XSzIjec9G5XuoQlKCkO2eA09eCAxNVjgfgda6QoUeIKWUGbKyi61oC7s
PgEn0cT5DcL7jT8Mn4mbUVWyb5ZF5sQ8mEn2hlL5tJlpZUT6SDlJkFgplDtkJ51h
UUfjQPe+aT/6pJ2Eku9pLmqeD29fz4qY5YBao4wfqmO+XIuYNGNt/MCT3ySgjEwn
WVxp+Po//o1NUCoFg3Nqh0tZ/sO4OjUS3yPH5lvX50udQWdkfLVFfydTuXgaWdyX
5Tw5IfTtFNPGgiCUOeD4YzVHg99tMEgnbMgmVcnN0woIEAU4BMjSvb9GovbuJepO
cN0ffFSWYrvXb3NjcwYdvEtuCZj46tCPrxMgko2kxGweGF4JQcqE6CyeMfwgIXlK
OTgmC3tRblHGRRBBcaQ2R7ioLb406Vh/5X4Goc/gLuUM4zkP3BXUsTQ87OsTWfFa
cB+hLmaWSg0Gdyn6e9HiyXfOSNYiNVJLPtuaNTLCWd5L3yGfYrUbZdMAH4QqHoH7
XLU1bMr5H6fQhyVl/jVIdGJ18ny4myCMuZm95hjZYm6Q4Coj0WOe0yNwZdOJt6cj
EjYgBpBgNn4HI1GdXVSCzaKqy9ZO6/lIsATlvByyqXqnQ91NcqvIQuuMS2znCkDR
eiztz+HYOJ/ZQI/FbP5og1+5WeJSlok+Jr73G10nflBOwK3aykdT3Gqt/7fjS+kb
LBnZeIUxorQyJefE6UQBHwF+Bxm4goi/jgvCXnnJYdU/MV8zrK4DybpxzRoV0cnN
bf5lSqGtKUj5xf7IdDAtegpuJqYygebExiIuELjp+KHIzwyfWBUq3o/B2bYJ4Slw
ZrTm4BQkEOz910ZDmnly6oobP7v9t0Em8lo26hdY9SLkcmasNLcD2OHxad1LLG+c
5qsxMadKO3jL9CU38DFq6U7aJ5vOYHziHmQGCGdlx0ZewuiS1zpE5B0zDV9vbuvY
h59+Mv9/hywB4tHVsivG30rNlE4jGGqE1RzdR37g8lYpNmklHLtiGT83pH51lPEd
5b7ANfB8xeaAjiTRlDg3aZ3uo/j9c829CvfCC2TMAA9TVfPTBmfdoyGuWskN3HHE
BWxQuZySc2m1CKwG1XgRb+o9jwtL2I5mCcs1NC1k4DgUf2qd3jqtrkdsaktWMnbS
l24ov+DAUHtG/A60JkZFn5OOahVUaTsc+RXqqWmNVKkt3vSCzF3oF2TBLN1C1G/Z
XMxIW6z98jCGXfVwjWXkzjTthkHG3s+2UUCKY+kXINeCMl8GGahlcbzfD6lXVGp3
Ray5tZkMhLbe5xjBt5MHbwp1su6s3+OEP4eEfqJ6WpDQhMn+uOymj31Uii75yT8l
WiTpJXVgwxvIfjbRHH6qWO9a+duggn9M8GHzJoHyuSTc6Ld+2NMg1wh9roWuVCbk
vw4r48GoFDC5d/EKvrBP/UCrjpWFjDuirpbfx4F4lu+Z1f72toVudzT1CO9AapmH
Jb1rJpHgjgOrpLcCvYxQjM+nzJjR7016QXnatqTKq/vQBbdDMca21dSZzBC0fPSj
21o7GXcAygcOqQe2/U7JXjviRWsK7xDEYdfUNqV6RBRbUJFXfXAh2AgxgAVm08o1
ZvFvzytHVJPpLGnGq3WzUk8GfvKoHFRgqRjC5fGON4IvQXcgqBQ/pd2DPHpT3iK4
CKwAtlBIs6mAJS4+/yflGN9DnAnSNQTGTKHMrCCxt7RUloM3nanO3HUXRa+uzl13
my6Rbu+f/qEojKSBfFZWsIj7550Zu7zyrpV0iiqdiFDrb4SgAJu+HJ2su1hHfeYT
bH43INw8RVR0opnXmr2F0CU/eiqShyVFjAyIUrPbFekLlf7OXwxRvwAkTvkNmkzr
Fz9/zbBz9ObafsTxMYw9voBGWkQwGQBj8P0smyAAXOgCyNjLxaFXOYXk+pbsVVG8
Pzy8iksHeXY3uTmM72KmhbvkOvEjHl/rYEJCNve9NXT3karW2If0w5JQzxs7bT1r
kWM9qb/GFFC69RVGq5YwXfYy2eBzr7e8Pb5Tlsep0Hl/u8p5dDEcHJ2/r1jKhgAI
h6srTJGBAtLVa0bSat972Y/q3NXh88J0d9kOsTi31DTKF/oy2vNLXeZFV5hNDgw5
SNFGC7mVTPR+rHveLhfvMw/0SQ5V4ej2vQig/RJWkr2QjIxGkIFU8B3VXyiewvku
Zb8hK0f/uV1ezfKDygCy8OMpZDHgyyq3ARRrHLtg0TN/aDrlciSVYDaDxi8Ttl/B
qiG50i2Ljrk6wfP6gG7uv25lf4b0wKVb3itl4gHqmMXFj/xYtIUcK3G70vvokF+e
Kh5BupT9CpgTWyT/twFB8rrP0DuHe3+9qX/x/w5vDEqkE5C6NsyhhetY5YXevNkQ
ZGtL38EuNly2yp/rvSl1gMPMoUDuXbkw7Ks/2NP+vy8jnqEEvw6GTVviIU4IHIMU
RkuTY7IyQ9v7A8+Hg7RhMBsxvT6fMccqK+/LHADc7nn5MuKep4rZV3Vw3nc8hZcR
AtHZrV/EbQ4tV7gjqMwZphxWNmiLV+H7bXDuK8O6PZ5aT5obyyL/OxiKWpfwllne
nwHhxzV7ktjsOtfQwYFB5jvZWa05crVfKrT1hJbjvtti8Nds9z9hvDmmfjDkvkvI
7prVlvkz4fEU33TRlkRxB8Elx5yoqD+4HQZPpEWvRr7bJvW47N4Oxe96wIic0hyF
wgHkOQGnwZHRPjRH/afCgEHuio/L73bFlHEONiA39C9YQ1WZ8gslqqQUm2HimFbg
Hydxpn4OkRubm/1jvsbBVQ5XUwielztQHEmPcUWtwOguy61d7u/XZLNXWpS6txqd
SHZDaBWVBJSlguH6pHJ78/rdHFlYLIiSc1T9rf3BB0i1fkl+BFq0I855nOrm/O+n
axNJsCN6SMmPT7EHXW2Ww62kDALxEIWfVxBgEGPMxKpwQZ4tzfGOiURM8JxwapC4
KQEpZV1Z1kX5duq5vXFSp3OsEtZIzVMstwhIEzoBigJ1/KdOWRjn2S38TvxOon4L
B2/jVhr7gm+c4Alh3pEAodJd5CgYIgLZ7MMg9ax8Ia3GWIPa49eNgOtdSkShsPiX
I7XjmOZlp0dZ6IqCq5cigLlWPqxQglfH7Et286hlmdDCHNm7Ofw4szWcznFUmvHn
J9Y1t9ohaIdZVCYYZq4cJdjx8fOMcG41jmeiLFW4BolhLVKr/nSugQuzvWvJ3edJ
QWlA3D7BPhpCoHJklf/sfjAeYr3dLmyx4AvjxCiG+3uZ8+ddYuJcDZ/JPrJJXKpg
7r2iG+YHH0EPwuX5EQzEuEtGh6TOnSF9OpOGzmqsB1bBBdl/WPjfSKShnhNRtIyK
ys06dX4hj5VzHMpfPmV33YsE4g1xwCGbBdkHFGHVo+Lp4H5u36b9adtoP4EkXiPE
ICo3kiy6Z06rPcpV3wGROoJ37QS/Xs9zKDyLBNMngQODuQVmzdOqdHGNecvP6Ama
mpNGORzXRlYa0zIR5gpgaZKC2s6X0fWjq8Sf3c7yNQqBxyuRBGDroTlgXfFPN2DK
aHQ1hc4I4VhDCPldVGMOgOwkPEeLmcJhnLhMQUwpcqPTXqEqpkPo4do0hdkRuoR0
3Zca4zjrAxxg60DJuNTjqXIY1bITI+D3F7pv7YVFIjUhwymy2sdsRI2B/jSQGaQ3
uW5xsj4aKb20HKg5oYpjKXnxYRg4jpmuj3GCPeKuJZCtPfUPvrENry3MjCpQzC7x
AbbcPrfdbrHToimZl2CAzHR9JgBYzMTLMSBWqvTLiS+0M1wWY9kGunm7eat1XYoE
cnvu26FtfJ2lh3jiErO8ibMSXlxpgFuhoMfha2r80eMmCkx9h4PfGKL05StsVh1N
TGVy/UsTUymtiuPMlgIV61jFyLb3H0HSR8fvt+TWy/GAcM6KhJuFhUvKZKny6fba
yfExRMIC7tuzY3+BSDJ1jiEoZE8NG/wi7DXn684peWrXv4zb9+SCFMsAgcAS4iWv
5R6PoQ4jcwCCGeAKYrwkSqMKd1RZaita1HdvkryIRTGDWek/egiP/dp0G1QSjnBQ
xQHVQXQNffeIQ8Z/15S+fDDkvqFMaC4PyI/XsSATFJH+0jhvS0FJSgFJ/X4NudYH
vRlTsUNvIx5MPQjyBEh3c5kvGBHBDwFgZbxB4iDUggQjA3Fn2GdeRPzBqrzA0gV7
JUbsoR2x4629ywc0WsfJyzLRKhhKW1a8+45nmK6ohtL9FwHG3xph19hyMYk2IF3H
rWec5dzXItmKfRPvbn0eNLiZE/Tfk3X3mnQfvXxNa4UnPpGko87Bn28m3bXaZ7OF
1+uFmv/gF/xtAsgnQLLTL38NdaA54DkNl2XNWsPvM7BAe3EmbfxtNLfzb5rS3tQS
G2M4H6Jto3w56QAhO3PhAW/kRo1ly3i1ZDInEHRgQ3Xmfm0+8KBpgX5KRuDObCFF
E7PIjUgD1+9bh7MAZEesMSanRC3+ulTf0Mi7wDePiQ3MhH0CgkAfnIgbOXQqIDYy
BZm8HVu6oAuUvqDi9sY8ve7gGwFjUKyoYJoMDVMTy/xAK/SlLZ9cCZo01gyg9SMz
JUs1b0WrcFT5QwcKFA6YFh1rpHnfE5W3hlx6s7OtyZwBGydTabG8KHGPV+0161z3
ufmtMgT5UCFAYQxSyN1TUiiwZiQAoG4HFGT3OKF5a0Lc4dsQIe8EvPu+CdlzPimZ
lEu5ux2qWavdgZup7knAUjmKk+WgT8mmLX/s7UNlyCJsw+YE87wVTflHg4+mp8Ck
4kJjwS4Vq8OcgvyXwS9bsRlfPDtF8vbTo3Ou5x44cADtw5TDhmyl0QS8NZe4e5EN
lX9ZR9HEfFF8WzHlp9VsGaPCCSlX5WSpfsYpBseEsePP6Nf4n1YGvbUJ5eSbYVCy
oofNjcyfEni0HdX6oJ3tNycehjYahGl6XB4D6H9KqOVf5S++MLRdckKHr4aasbK7
NQP7GyqFtZSyWUbEpye+rKRQuA3za9OWshCeW+foBkUfLq2FjGoK1oOnmrXvFvle
dUBHN0tU9DAdpqAMGo/kD2mshV8AZ2EA8NYUuHaPVVBON1ngJrtmgRXKWPQlHVMw
8dfRkR9oECLWgyDZOD6Rl8hWYJRGOGZI9GpF/WnQhUAmsvu1I2JGsxrG4HCSVZzA
umhEme7LES+x8ZcEVt6Yv28GbuN+DUGrDxsZaIh64glgSplxBRt4InZaezzjcbDg
aNqyyHmrD3Bb2kNhzeK6yZciJkLk8cJHQJ7vmhgseEVHb6mXz/O/5TZHrPPXSmQr
LYvaO1+OgCDkaSWc6gtrdVUtlLfwSRXaL5Mbj6ONMgkDZIfKLDfacBoczkKopRYD
ZGPFBvFvsnpYruD20/9YuzGFbWymMsP+lYEMWnkkcf3pH4VfxmOAN+EktM+CRn5a
UQ6V2crFy5g711ivCP44A3YHSrBQyF0fCGBkGfHc4qkJIkTwTTcsPdkox8Ymt7AN
0mPbwH4Px/gZUVehJ+fgor9hgjCF7GT74B4BpLF7l6KgRhx4IPvUhh36JN77W5lD
Q2hVXmb/raNXDmUH2XU9VRH8SMR9oM7lVuyThKOHJ63d+mE/WEVNqTZIVEF6KFgr
56aqB/h6jrq3vKWzbKINR3BXET2lOw6ZTzs3N/edsIkAU0PYlxFxyxC/3p5t8c5b
c8dsVCK4pbOPEwAXTr+URrh5IDDOb4wUzJoj0L02cEyUzRGn5BUFYMdEr4RvTofE
B+LVErxLt+xWZCGVFhpLyT/VTRpWnf6Jve6nRBU0qukvqrLjjknFwJCllDhEOwwA
jcMWXvuzNJtGqlqjJ/RA8QhpUrru09rjB2Fov/bA19q/+1dHufUf0fdMwJ2w5Nyc
eJR7zHkIorEbCvvHeeHNeK2fYgv8fA4jBXzS5ZVgOXFwvb047SJ3UaytpKKabGB/
uhG0lGUcbIZJRokiCUAWVNYx7i32unJebAVYIzE0MMnFayfQjAUeLRry76Uf6EYO
z524EDwChhVb6IPJye/YrAEw5tuzaSvHc5EfA6Ew2P6NXECNyJmVkk/LIpBtx0pu
rAKdj3eHS64Ij9FgQZcxu4jDxdamMjPQdvqWxv7cT2bJ5dW5ByoZPDbpg10seLkX
KWpGOAUXAhj8QIimQ2ZpJKnL+GCja82f7JpqO7aqf1xL37cNFAgdh3/mOPVG6ysk
ozkXrHvFgw6jth6wY11brOnwLygcQYIGukG4XiCsXLVPZ6jMonRXktp3FMqpRl5/
eFfd9pPnrMpSW66fUinRzJAFnQGzo7dK5eNkqxIRLC/UKELJhjkhMHprlhXr7FWt
WFPCO98UPCHKxT8SFuIICqgp32Cf+C6wcI/JKIts1IP63CJPJK1AxlLspQ/Y9fGs
wSphawvIivc6mz4oaSKh35OMeSYpCKKn3BG8/xQH/p1Vxd7uIZaXnQgdnTukBXQd
fZXrX7DFFMD+JdksSKd1KEchTW4MLUZxbNpXY75PPLpcX/CnTfR42IHAePV7Gckz
Q3xdSmbSpi4zYDBpzdpxquPJdu2hsKQSOy8yjODNEamwmWbecI6Zx9UFE27/qSh0
r1UMO7Znm8f5cICE9V2YfM2Q6k5X01Vb3cN6iwEHoAGuWHrb5NAr4CQh5rdlP+zB
77Msn2t79T1nQCN58/rZwMzdBhygVJFKmbrm9EOSb8s2rJwhkOWpUFu4mYEJUSog
ONFBlj5BTDN4DI1FtdOLhn/WrM6sA/4qfW2ecYnl4IHFkX/K9HdpLz2CfPT8gt8n
SSivmq0apw4aeHwzCyuxw6fx9hUv92LsTtapWgeKmXfDlGpnupj09D6licI+u+H2
lxcJIluj23v80ddsYZDF9zOn/+5AAaiKO0K6u1Co9XzQ8h1owLsOdVIV6I4I/VyK
C2TowxY0lrTpvD3s2u+7Y8bdGfDpEymkWq5pm2PJk2bj+DZn4ZTJB1TaSbrcaE7B
wn4mpBbsPkjZh50etCB1isasAF9scDO1a8nXxKLB7L41pYR9UQ4bLLst9tQ07VQY
BZzZT0ZUbpkzL7fgB55IneVVrH3LS0JD1NJYc7BZ0EAHR/zDD3OFCsFmLM+wp3CY
0FaZKEVHlAcWNBEnoaky4zinU7hNTxmz9AI5GAG0E9JiQTH77VvC6HbWIdOoWAVm
nkAMUi4hjkyW4K+URd6MJoaIXyZgoEIItrxptdE5iq8nNi5SbqmhqlnmTxnyddXr
uBvNyn2SZ5y00QAwgm8kB1ruLmustjJ1BPWNO1xGsv8nEMWB2UxzCWPojutoLhzs
6pPdTpBdF390vULORoYLd6X6qEoLvOnl69GNn9uGICXs2Q/C4AKAd5sryYR0PNlg
wVOnsKqaI7ZAePLGpK4Yiq8ziKreHTqhfmzN1b3EB+NMXnCrcbkYX9zPKBCAebkh
PFK+0BcMZ8s8LdntOcB16Q2vRYvDW8EK+REnZFqg6vg0UBW4Y6+l7SGN8atdig2Y
k60GFIDUHrA8uCnzE8Nn7C8P+rcKPjsdUA9hs+aT4wquzbAFbZ/MfT3d5b/jPzB7
9L5MVjX4nIy75VP5IIF50LQdx4UoHgshHiP+2AJD2Ejs7b+3MB9/68r74hyYvnKK
PUbL+Y5Tn3munlQj0NVtReVQNyImG89NvPcp8kx1ZQMBpxobWAUN9JxVUx08ehmn
OGqztEYLWGnXfirAhT+PalFR+oh90JajIsPrw+7k/7vvFSUTtRT7qfgDxp18Z7Eu
XNu0u3d4+0Jzg48Xkham4EoN265iGdi+BPGEq4OMkgcpxDky5+weulng56kqz4ss
/08KghcrM+AIVIUidk+Wmi9Vm2KhmMyytm2l3AnV4XmEMrwbdm+3dlMD4f471OI2
vydt6dV/s1weMNtjueuH403NjEVfIUDd3yrL+Ezh4zOnwKSF5eds3QMysqVjSJiJ
beJIrNguARvdynLEi7DCL1p8vKrD5iX6XMcsfpJhFxX8KFbXGfx6l2wznDEjLGCr
edxvMEsNKFZSi8yCof6obvORhLtr7jqzJ712iXGc32RE4xMTCly19qDYZpt3ancS
pawI0ZSIQrjrWfjJYYbM8bNIsrYR9Zbl7qr5T+kzFjQJBTb+KpRHmTZpHL59mdMM
EKlT+hU284fOq9Hl/6Aepd1YH9PN9vGdFiejKCB2x9TWzjQhcEtlgXgYsc5WsS/j
GKKr2x1itapwjQP2FrlJzUbizqYGPTxKRGXzq7MkG+uzuVotRmWNX9Ha/LR51J6q
viCRmDV9yjPYbKkC90oJCKS53rHmzci41r1xFwBq+TXcMjoq/E9Kp5Y+DdHHrBTW
AHlkiFoUKlziRFR3FbE/j+Qrqc1GRrBF0GBhPZeaNxovKOK6/6ORa/MF7hDqlS5Y
xlY3GWH1otl6kxazX8MPwcqnwbn6KGDIQwPtp1u/GCQ7bXUGjj7zBMjhHsoI3BnC
6MEnzkdOjOqJ1oeV6GqyzYkDUFbJL+sKClT6JMIdyVbkrOYCNDrEm6I1s+FivxCx
dmswGfiIG4DntL+vpC2jTZ1MtAya0tax6LtqTVXuwoQqiHEfUigiulvYEby4ZmHi
nwDbMSFDPyEvNbSyOIM2RWjIYl0prKdgSuXtpx8O7zO+mg9vd7fRR6Ohf1Knd5jF
Zf0SL8VreVV3Qadfvlrms3cZv72URht2PIan7xAYXkUYTql9ub/Ndl/Pbt5h66lb
GLTk289JX6q3DyNFB0Yhi6BlsBpxkZLvLoW0ngJkZjeGMAGTTcXdwrx/DLmPRwTh
VHaXrq2FX0hIjILd7dueAr3Ksetp+rNLrshg05em6YQFRGR2V+GYp++VkAs0MVi0
A8vcv3mQNSBqfsQoRecR0htKAn8tP7L8pxQlCHX6+WXqT/zfyxdRWDHg02veFibI
wcR99lvn4bpH0vJg4ApIWdPA0S+qJ6e8vcANBT5KBYtphe3Mec5mZFBL6f+Qtk/y
jVpp9FZ7Wzeq7UVFXC2EzQppgm+ozfS328JynGiADrpdkBzeIhk5PhunTZ0SdYtO
xBRDYQRRsgJ6i9swGfgcsyXVnLPgy40EXSouLyrfmISxRHVoNgrkQ3TW62ngHq8Q
aXDXQDoh8Zy3xZqBU/8oLMlxJ1fak6y5J4mrO/7jmi9jDGTfhBGT4WMyANxX3MVC
t1jzIOWERfO1gC5NovjDsk4306ydswJ2OqBnSlx8aCxU27vLWwkMxP1iNxKAQ+OW
EIYTe/sI570BIzKEC35GtgnGh6rpaGvU1hs80YjKHUWXOHYT5q3iE9nQMDBRLbSG
TrX/fKcvPLShg3ygAUZLDGVzLvHHiv8sWvWJLFXU9aD9zQmZ73Hqw8BLBkduydu8
p5vTPZ0NMoKfJECQrTzQbn1O43hE8wG6yWi2lqRM+ektDePjUqWmBoXgXHfDLsRk
x9hzXjUUBeFYBXQQJX9KvobImSVuKKZxQa+buM2rkiLAUuqYr+VeHmoeEAjN4RcJ
RGd+NEkPpRkbo3ZE+vpc13XfhmcyH6OBhBg8Q99ybUCSc1nWFwoKkw6lv4zNWy06
y+fBe2dxpx5jxZfS0MoWXzpgEwsDZBNsN88tgSIlSr5k+J5qJHW8s1dFUmPjeFQL
1AwiZdWwWoOCvg9thVEhNA4wo39M8rrNdHJNrfe/2w26LZfpLPCSeu3dLk/5s2aE
Zv7TdMfgHQOV4icqVyCK3LbuLPCKs0lCjYdYCf6s/kuWF2yyC33nk1cD+dBCD+b4
BUp2AHZBHD294UihYPN+5YRYi6nTH6GZ2170F6dozW6+121XCFUAFMb52kmIkDc6
uDTkJJDEsYkgKzqK4M2yrHu4Qvqv4OIFbdcTNMsA8hzz6AHyjFKYXOom4wIXCiYM
ui5rgaMbcJefVyM9RGjdSJvwZyFn+h/FvyMUYTQ4G3YiIdJompk/qEbSsuv2Vjae
9sxgLI2ZgyXiQoXHbE7fTJDpJiAPFGD8vgrXIqFaAEVcP9SoP2EDrZIJOG3F4yV2
Y1CKkFS0IkSPROthLD+X32PnT/Bos+O8Mix+YDsJEwrJ1tHB2lR596YUiFRBw3cC
B5ckQQOm4s0hmT2ift13JJUPntzaE3MFa7wxExSrW+y13c4PKxwy6fTcI6UuzvM/
TxA6ks4HNs1/uFszGd6jHn2WQs1nnJY48MDJ3FM9g6wAjpSGXyLdEQkB09mxXZFA
a/3tu8cscv5f3qNoMChNNKGSSgAmb52JsZEqFJZuLUi7WNsFhVIsQj6td1Zhsd3o
+aZpSHWFf7VCyWtL8eIIEInYYYe0CQ5cRqqnhXZDStuklGjPixEJppUm21R3B/KX
68wKkxZ9Db+Bf+H0OOTfSMcxVrV9BFPWfhcobAEwktsCnkldCl3LrV7/KKrlJUQh
XcwPZEB5n0FdpNcBSwQpp2PqiRk0/KY0kf38rTmZHRt5TNKY4ucKCDotLnR636KB
nnTE7uitupxdtWmds8PJcXyDq2QfOROScJe85MBjpelT7YGUgBi8EjvuWVyg+is2
cD3p1eNo45a/bwRRyFOCefPsFGRoER9kOXR/Ln1vwTwy7QKO7dTsMHcW4QHvFbNd
5SQzdwNP2swdXA1aH4cP/xc7P9QLUUBbYS9vLnzKucWNGu4PyE6UPjALC7X8jcf3
YZ3UfGFrA/os56YbCnHEs5oq6CJxjoTog+7Emc09s/AVao4++bQlAScwIEwgMqD0
27c+tFmdxvCHloWofh1zd8PElkAyHzj7WCB5xrwxDtm46C0ZiWIXDgw8zDyIUn98
qXg8XdJawXqv4Fs9ac+oAw0EDBD+CbF43pAQbLk2nTA/1Y3ZTVMe79Qoh56JcHjt
cufb6S4heZ2jZ8SLv84O1tXVx9qkSE7inALwpSbl55ETfLDOz+OLa7kCgmpFNQQi
/39QFkTjwH9hEh+pn3SVAHxUJtJaDjv9XbqJa5kLWav2vcAsm9f+WFPW9Q0ZZ0Qi
wLyNOaK8IWuvb8M2xw94cvL32n35bdYZYhGooZqDzLH/60DKhdOQwpLS+1LNduOl
aseFzWMDsmwOcAF6lHP7dW9vZ8tkP/ugEl0W5092uApx/m+cfBVCP0+ySuYy6mre
AeoLNwDz1mXO4Y65c/Uih1eCj2vhJmJp5huJTgLSmAUAzcpg+pON5sS1dQdP8id0
NzAhNGbtlg4Wr/YfAK7S/O6sDhI4AZToL4hGZzo3AckUUHiNo+qGlQAD2zT6rpcY
C2WLzkX1soHsUl0h/vsQYfpsWK0wMES/dIda8aoXvQMFB/LM4Ew61iOlO2iNumHw
OawMj7wdABGSHp5JHV3bEcbkiTbeRmbjuO5Ld8sUF/o+PRXzfb9RI6SomaIf3CKD
MayAHvHHQZL2sHypbjlp+CL9PHZWGMBN1zHnwNL4RyYcH0iAG4p/IA1fUnBxLh1Y
ao9Xfnr2062v5DlW0ibrnJEwLidAJ6wRN8sZ1Gja+GbPJhTyEKWbwfaEwXnIoGMt
3X6vvudFtV4IjljIRxcF4lDWykGi4EtcWZBK272svFndVspl4Wlrgal1PiraDSK5
Pc1Fqb1VYjmlQPkon1/JOMt1Tbvwo9c6vFwsUSMUyE3cVZBWf0SJfyomc1FIuWWb
dWdNS+tExvDqy3mGP3fHiG28avELSKUPNcIOAyDKsUidyaC2052V2336hxI/DS9l
ma8bZdtXj7XYl0NjI3YN8M2VezklgRyTA+YbqCUemSHfFQp+heJVr/obvB8jA4kl
Z/GX6PJdm9QH1JFUGWIM2f3ZrHI9ttceA0QKLZ91Q1Qoc6lk4EnDG05JvBg0ppHb
xk/RYriXAeVzkuYoPiGMrZ5baKfLnjlWL8VxqA+sh4NRF3+HoQPK0zIa3w0IJygY
AuxZV+x5m9QivPc7RN5OLLWgDCkVcW7Wckw2VVXEshi7L8NwZJAbPq1sUQocyrwO
YiHHKSuQ3I1J3URfCnFmhoPIiWdIFDaZip9g9lvNgHz0cT35f6jr311SDZGDQFO0
Yc4w8aSmdXHdjX10Q+KFFu6LtSc7dxQQo0uk29P80Li+nBxeWCTYGSZZ/ZtkJx7p
TrYKzwYI6ue5+CeDVc4odlOGLBCAytIIvWefe4u3zNeiURYgX0BdiD6phSoze5n/
h2VR2MbCrXo8z3xD5PKWYNHFZsFdqTqSweAzg6FJJGsPmFyDNBBQXhOrqmE35ScT
Ize8OxfTxVqdIIqZ530zQU870Dt+BqaADzmwZzkZ9ATCIpV15sQjDZOo/QrPVGKC
rAl0iZvmhF9uad7IU8q2te30u4kD/3uFTl3M5bEyHBQYjxgQjw+Ty2wNExtMAnYM
au4mridk8owFvxsOuT5fbQvPqxOHOLsRnRrrZlVPxpl8nMCjixjGML0x1+KR9XoN
xO8uJ4kYpSYrlsHZYJ6CB1iQtpbtyRwG2O3I2apseGTJPFlJHedxhMBGKYbraFvD
hPY39y56YAhwnsaeOBlupptCh0CSB07fatdlyWICe5zu24vj3+6zcJahL4dhfyGS
Gy0sW6SL2Kl1nqqQbqTbFvEggmhpHGPZNNLQ1c/ItIt4FrJ0IF8RgE598cu4wk+J
l6vJW9C1GSvj25uTeEtP1BvlWsXFa7tanZSaxgnkQWaitmoyZd0Xq/BU+BtVDnVO
mIDpHDDpW0mHyhxqGHFovDH/UGmoLB74OW+B40h6q6j5XBNTQIb/G3/f7a3jvRcq
SBszsybqnO9dHEHntbZXTrCsXEq1CyhjozBz5hrIqD2oZ997szboHCJ25xmKXXj0
kH+ZdG38C9ouX6rF3p40iwZ7fZwvosuSA8N37Fd+aYKqVzN9HSJfJAbYhXgc89hY
afM2sswusGS+G+O0aiMND58m5pnS56bRCth1bOUPyTKO3g5WCrN4az5q5aC6vusn
JTAtEqVdUrVdAV/d6g6uv9cOdwL/AkpvdQOANul9NT4Z7l2ScP5t7oiortI+8F+7
0PuKRu0ajW2A2lnwS8JVypKPShvrdyb1pBTZ9b7wyuWDPvgbh1Ji7GrubBH+tn9b
N12LeW/rnbDVJ8wOyBZZaOqO2e0CdA7jaHEvOh57BANX+VpfJpee5tyL8S1uv7FX
3DYp2NCJGYgBzj3w0UA2w2TSeN8bTmQPCejBKUsgcIepGFydmYb4H20usEHJbKRG
oWN+66vQiOSv9EU6Vz6UkG4iHR8HuKDBsN0SG6JGeiYg/fqgRnLKMv4YW4zIlGAN
+QJQP/rsIjLbYXJT9TzXNW8sQHBqOS9bLcPktaP+w+a0s6hFLZSvNtzvfMm31kPQ
q/aGXdMvoB2DAHjrSAhqMVgScAfJ3Fa2bfDpNx5v8aa+iCeAs37fAX8kgAnJntcm
R3kMmM6RAQteUoGc/5bTzoCsgA5ESoMhrmNS5qZkDOOD3CKks/gWAI/Ga51/9eDg
H3lZ0YJeOGgtvZXJNRjBmgryG1MToIIzKxk+NzHGOrp8L5QNgdpqzNI3ecClxyf5
HX2wdBaenc1n4ISWy91quGFRzbH3Yw0a+2PwwKjl01O2TGIcuAYtof2YWwDOF6v/
2UEEcRAZiOXqtiZIUETRlUmi7qtJs8o5pGeJvLVlZziHpHZY9yFjHEWiNWQLCHQ8
UX7Rr/XvLoiVmVIt02i3m6pnR9TnrTvRcgvUWlPFa92maLld/Pr5Yqdu3qpbRFX7
/chQRm4HrvV6gjCnDfM1gbbmadUXovMkqAm56RtLDca8MX34maz5EXpJRTA4UWN/
SMZiVGSSiIKWS4sCALU28YQQkrpi4OxaJff72zOi1rW+IF0xkF893jfwmNGQinqJ
bfz44b6reI3GdumQwyCjm3zWB0VF+QaICsoGn4A9vW5hN32K+Hyl9jXCwS7ZKz/x
YORuQ1ygUjxgE1BszsMduuEvWeeuN+5vn93uBDXMzA69gjlgnm687mVkNzWyajLn
RFtArW5ZWxVxbkznho5xgbm+AnBZBURrhvAWFusHLRglxP4uDUv4gnWXPZxhllec
8N/YJ+Do+M//mK+SuWyVY07+9dkmYMsdcIj2G7NFJQ7X0kKcMFYg52ulNBXdTHlV
wsWKJUkfBOJo2onpAKml3lUY8xgf3OHegAvHVSEDvSi4upnsY7Oj+omAqG5wpAEQ
vcXqzvr7ZxEuvtssQTuAyeMPA8SxqzNJ1bHR5pFPLQSalOVGNjJs1RimjCghWuX2
dI0jM6XkJgyzFdXKW9WKlUnx4ec1fdLPihC23/OS9mwcsGnIMuCY+F7W8MEigDDy
0DBqbExZAOm3AR4Wk6MAsk06VjcEz2aYbLHG3QAgLuxgR3T9W/GoVxXkvRa/brLn
0tBxSRDV1zTFsrJPSa3MNfM4D3beUB/VrWBBvKNopSeP4KwweXgnC/oWLTpHQ6po
PiV/S0O6r7dqw+d+r5TyReUlnQSM89nBdFYdrPHdBn/7bbhJfwe8UVShrVNc3t7L
dD+wkUW/z5zyWOi+lN/1AOQX92+KfWs5WcyDG7iB1KqSD/3bFXAEq6YdGNlZeUNc
b3tDWq+DR5pJxawltZ6V38sk36VXCPfGd5jzjoL2J81ylVhqEsQNLiCSN2L8HLyS
NX+NTEO1GOYItbDSircWjodXlrE8e8ItvsT0Dt17/nWejXjVmG+Jd8AfCfLDlH1/
V+v8qX/MfY+iaQuATStJfFu3qlgJjumG4xGxQjonQHpLpxdKrox6MOj+zjmLgsHH
Mvke0FjyWoz5b2uJ2r0TzViS7o8MGTuyIpYJABCq/zITv9Med4EtN5zG3i8hi0vt
QZMAlo//YygoJSkau28eQMJTj/jc5oCMCR2rck8T5Uam3ijdNBt/lJb1GaUX1oHG
d1zOg9nWW0jMYACsp1GVsL3agERchOD8hUO3sGyp9nZKPNv6SIWfYynpJ9Rg6nIR
0O8CpdQlfN2/3OXer0zNt5ztkrWVd/MSUYdVRrs8BHrZWTeMtGVO7jBdiBBNkIFv
z+Afu519XvDyFgF4++OC6GMk8LDVN+bUgBBb3JQzSph+g93aYHsKbHWxW5SEeT98
A18/7Dcc5vZm2EAgy3Epf71Hvtg2R8XhuzK4n208dL37FhIYpSmabOnk7VFKNXnT
dm+JPvm5197y8BZrbu77CIiRii4KM9pVRdq0cQFzcIbaqD5ohwE7FMtpxzGGamN/
Uv2gz4OWMstUaIc1V/f26lBDbfZZwik/ajja/k/WkxxJsR7on6SvK5RrfHNOgFC1
nnRDyFJvCwERdT5JTb7fI/uTku5k//S8/8jogxdiL88flom80XQO3G/WHgyJgK1n
KuVeKo04tHDCLe6spUD05vOyW010hBd1EZsN3dIzsopPtyGnX6URdW7SpFd+wV5v
ElGVpLQ9AYRHtTN7gbc2bAdE9y599lcdoTKepePl1Bf8NFF7koxZYKx1fMlYCJiq
lrhMXJgBmVvND90LssU0I77dtF1miuijQXLmWO91Gzj1ouT71u0oOEbcOGT7MrJr
/4KtrfIIVBpMEcP+n/seeTHlIEpduHoijxZt796W9XTa0ZkDBYKClhTxSfgE47wQ
xMaNKT07EtOIhZB2kRmk4OYrW5lZcGOqHSlKgYpjpSi8/CAOmWxPu9cXT3I8EW1D
haNhjIzmxqeRrDBMWSlYSJtyM3gRGXJGrWRraVZIavupEHHeGW6pRto+ASw2ed8P
w/ZU3qCqSAw6VIyJVrTxdh85FYZbyem/mqNp54pjoPeVx3pz25asRHkycn/eTkEN
wlIV8f3IvC7vI07jz2QnEv3E6BpAW0FWrhIO3AQg2nI3g/rKNyWlWPoGtv28JQYs
xwkqK/t5o/OVLSgBrudZlJeeKepH0WjguR8COyRI8qKm+rSl3/GORnA1a3bvUYZW
9aHS8MziZnzYoFPpIkS8QI+UyEvJYyNIkQ+KSnjGksNHsReW4OXURbhhRzLS8e9a
TA0LA4yMPTfaSp0et3eelNVJKyrXJfLWqTUtbJ3dPaKZQhd5mevJ9HtHU7vbkcxw
cASHET7lY0LdQrtmZgsJbebqqBqEtEJiPz4Rsbu/Wdfqn874so6edz8oXEtM2VXV
xZf5Z1ShfUswXqai6w+e+4dd0pyaRQk7LxPLsMZn8cdQtKSMHQzLWtxPvNTf52k7
xOUazvuGGOsAJvmpPeT7R2CvWLkn9s/eSflLggnNio/Sdvoa1ZhQ1Xaa60FiGeXR
VpfjewHaXv4E+EEFWSfZwUfxw/6R1Z/8qRfnzk9h6xBCXNONTcIynoiUlMJ87RzF
nRvbYm02i1g7qN+7ES0ubbBM++6/lAsASP+cmEa2zYd+/3SNptv5Lcj0+cr5lzm+
M3IdAK3OdQvT0W9Bw0LmAcA9VZznM4MjitsqP7tZijoz9LsjGnSU4EJIEu+MbrBU
rdZZC/9VLLF4EAk3m4WM8FBq8dVsUWTPvsw4JEikrMSpajXZ0e0H3ar+1iR55bct
KZiJgkun74f7r3AOuXMY1QvVOc0UMlXy4lFSwk19FwKYF9U+mr61zHtktp8zlohM
Z8kYmauKZJ549j0FD1j/RrLS+zL2eQCPMqVdYybwHIPRcPFo/W5s7MWm1ROxrcjk
imwTZmgEc0LjkNjBEFupeSoj8GwHv0T+FXQ0l+VpKlurBTLeiBlTw2YoHHVCrBpE
PapndYus3GN9i9ZD5lUdCcyoPJpF1u+olqB5/XzQDvjopasqpqau4c89Ch1TbRXd
ODDfIkCQ7haJxn25JxRP8jxe0Ev/hoQeM7VPW0Nh8tN7IdfLM7vhZaVwzXZeqxDn
je4daslRcUo0XISAtj0xX86Pz6O45+9WS4MUfsePogpvzxsQZTMM+5xgec9WE62b
UPsfDWOiSI5KeFotRunIh7v1GWw/HhgbGhYnKMId3YXrheLlCGN4on679cAvyn6a
T5X4YbtrB7V8Zsd/8z50HQ8aE6SqjAoWWe7FM8ZW7fpJyETLR0d3zsJgcecSXd9f
cGhXUhJE5LbMk3na7FRDZnE1jRQj/wJx1J5/3bIcGBCM55/le+SKjFDx+1wPgkvn
8eWiU2TBIXqsmOivt1EhTwrnAVke8glW4y+6sluRegP/LdJdhuEK5WhxtnZr8ZGW
1DfcfqfaXPcbFw4caOczjyhdaDQTT23NCt1UVzlmAcBNLwgY5H1ILtKmHqCf/qwX
Tnv3hqDAs4K4ZFh0RxVB1Kap4zZ4gMq7EBMS82pkaBU76zpYTe5Km1OvIJWF2Ves
aDbOdGu7qjRv5SCX2u6emhj4KtviZEN70tUyvPir9JbeE5wgg8XJqx6lnQ099bXX
YyvtixKvzsB1zUDzHq68jDLcItdTh7pAuKJqLXWthRFI2PkkbgtwoBSC8IRGWxAa
kjEjb4Tr1BiosdL3Kb6v8FccWpLYq40kMF+umOObnMrqaOfur73xpUYyFUYw01dB
Ruwujk/A9C6gNkSIGVke687tyddJ1Mb/nQfaW11yLW8KhzGYPzfL8RvjOO5Hx3dV
uTzHjf80kfrf06BaERvYNGPJW+EFUdpCqxPI7NJUs2DJP12nUwa+Dtw/yjGS3GqP
f4BWnE8J0NeH1eIL0KNLvKgjjsuYvw3pFERh+OmVSRAa9s3S+RYwS1Yh2g6bHOuo
DuxWx1Xay5w7u58nof2fX5BiWKfhek+91uU2nrieJYkFBG9YK54vY0cqJbQ8Dnnx
xjHvNyuiF1Q8YiAOb8ZiM2Oc9gFlo4uZDP7IWKqdUng7humK+LbNuJlNk64MC2Qx
9GIp+YyEmfx+qVxYwvFeR1aqpArKRgAaXB8fv0bNceoof4l+oEQFWOKk0qXZWw5/
qe8MkxeD0NwU7lWi/FycJzfnMtxwPMpq2riNiCEPwiWkwYG6VLym413mzTGx9G4I
EzfrQWMmQSHayWwpBTxEg/5vqFJC/V4XExdW/QEfWDBXQfkrnKcvffupqU/0N5wZ
iyCs46pZQqLtj6gQB8fvw5JSmshnqkbDanyjAnaGHXNoAeCsQb9eRCgc+aMJfJIa
mUZkMJO2PosMPWJg1HxLoG+UGzC5AAQAx2HcgiVrj6gMZRvHJj6r/uS68nvihBCj
xSF3KH6uK7xxzAz7JmWYTFzHVe1oKju6Kkq2T27C8KBqJG6rawbIZRaq+p4ZtW2Z
PFRDCBtJL42LL+h2HE8yYsiL+oUcAwSx57/1Hz2er12QJcaB0jcHjoLbtpJf8fzG
KxtToZ8VfyKww85G5HaltW0dayHS3eL7tlY3QTt8l6AqZt2ti3Nikvpo0AwtlPGk
1gakux13QDbVBbC+Y8jT2Zh18QZKvJc5nUqowltTWOBIyChi2A2vdjvw2RFLXJuy
oyxpJnAQa2kOXhk+9kyTMS3RVkB7LX+bYY1IE6khCohNUQwdT6GAzhnjEZh4+g5/
Q6S+dB9mWqynIEGsMXnp4mV3RjOqTjKPGtC2BYEcdKcJWZPz6OyD0OVktLPdl80K
0sT8EuPH7Q/KxQ8h6nr9OBvVyFYPY44mAeijbK9RtNDdG6ZJZfxI16NjN8nwSvSM
OU0+lT3gLz9p8UR47X/Il84noIzspDdifcKxvvJ/2f9ixTMTOz0EoYBv8dH9YyhS
AZcX4Z7dMMIY5HCe1tO0Ir4BSKiAfN2fbv291ga2WdrSfcIKQDU7oZz7TymxqpfV
HnWvtFUJLFKWDEmAFLB/TcGlOFFvbL3s8hCaMLAh99FGIEZlQ9JLeuq7GA9MhGaB
ddF8m/9POe0t4oJd+egqd5cX6p+rzxXUpYBN29wZ4NN9xPD0uXdd1ER7TeP3lnZG
joTB7baF6XAN6ycC0Y4yh/NqVjBCdaYSg5hO8Rn/u1QX5LXOqEIt1einULoeipHB
2MjudwRuMTabkH9lWIaavy4R2sbhK0+Y9/nRefX/Q69hvUeHqc3XD15fL2L5bEYB
tyxj7Vd95DY4xITurGP+Ycm3JYPdl48Y4KpSR8PXGHeO5JhEijRe/aUuoUii3njV
+HelfHBtDQDK6eKoLJ7Cdspf4U+18BPHLBQYZjHRKiQ/zoCz+Jez5VIsO55kWpf/
76m9Wv6dwJ0xG1zo3sDNPf8MRm1qvhUU7S7fRn85GieOGAz6JsfaE57qBxoNFNSc
pN1tI/Qmz679klSp188Y3ogVLMjtUu+WXTsXtuol5t4zIQxEejjxz7Nr1R04NYZ9
jskEmompHLWDe9K2MG+r3DWjloIowo2zlX+2pa6viWZPT9umRJuMB02lFpeEQCkv
37E7zTWFlw3DrFVBUPXNIxJyoMPVi9bbIlatuVl8Nt+mC7UZRV7OVUWyTip2UbA+
jh3pCWl/1iFe92EvBL+afyv+5YT8MReDLNPgn8ZAB6tU7OfBbUxLsdf+lRf2BBXe
+rmnS95cxEoZtfpRjXsw79urRH/gtv8VVXDPqcZ6G2nS3Dm8CUisaQWiUAdVBic5
JzAcxjLAIZ4oN7OUD5M1q5x5tJ+H72TNqcpI+Y1VlDWDsgbYNZg3JV0WiQaRJeZS
EAIRgK2+KaGetIHWZVorZ3RTKrLqbcRqwZ2HrLDwri9+BvO6WbtuE6/W3yLntKGj
/sjCGgA2kNu68kVegBd5kYB6TTmwJ2ULRk2gvNybpEFTyNDOTG+y0VERd6wqyBqX
XJrcoxRjonvkVez7NoetHlsfMhPS4ez6jPp4J7PRqY0SVv24xcWXaXXZXWUP5Gho
u+AP/xPWxEScsgXSK4lKzveZrTv96SC9e1Xp5K9LIBlzSovDU4T4XB5XWL9Mb4qq
i9fJk9YEAtd1GYUEucJqdGqui0HP9734AZqnrOSTNRzEqf/nC4BFD7ovk1s7ERnm
lDRHG+AFcnPekYx+3vqPyFPaPwsNZtAxiPE+Jhwr7kTNhCdXJ6pbK/fXy19RBgr3
2R1mo5kfPgw/ercwikdZ19bKREnOjnPjeEcP0woUCuGf80lpLk4PhzF1ZgGmduBE
Zd1hTwq6igKhDlVSngz5OgezgQJZ9yZzxZOUX12zY8ZV7Hrhk6Frzd53qlZMDcvz
hK8Mc6Zhz5+mhpMexPgnUy9G1FJfBAoXhUI/PGMYDDKQ6Q0HSFkgRs1EEMfkcsVH
8ReUFGE186K86LeF/BD9obumtvwrnPsr5YAfKNjJ7wzXv50qHLfY6SD05eBjbZfB
3qFBQmOPVwjZRa6RxncAGCsvLOovl0prnUpizRn0/vy/9XxjKUgjou19p8+cN0Sc
Re5/Gjvp0SmBptVNaWC3ob6SSZswxH4Tx57iiAT7NeMdsqrziKJoOWhquOIgP7rh
f2gio4ADLxqHVSC9E+AX5omJKd5ltcMS9hG06nrtf1C8IaB1lY46mfTo4DxFwkbO
fpUDiRGXo+HncJXdhI1rq1nZACHVHYvdqcbkQ0ilHfOnRkV1qp9NJlprTZfdLPjX
Yseu7R/ezx+pC8FByb+DYoRjjI4h6UGA6xXLIbmtvAr+yI5+7800H0RGYuiiYVff
YU3vUvx3YSLMc6dpLVn0HqnDf9UqHresoLSEPUkCObOiddnXjO+IYDFmO+samrFD
uWX7Vv9szWL3Ui/OyPrWLPY7ReEKGG2SYz3JYG7lPUymEhungAp2KVbnCpUKI14b
65F+/gbiUlNnJNm/SapfM3HtWnjm0r3BdiQ9nFjw0+F/rwVkJkLBsVJKyVCSjMQA
qxMc2wRD1ZfXn65PEyDY+NfVLWqSMaKYGuj5d8J3pbgKtuSzoBxm6hUJHQxWu53j
WVtYx/t5cnwJqww2gzcycA9R0oOTU5JdjXBN1ePLB7IHtUs63Fruvi8USalVGaTd
9kA+6ljPzy96Lj/70H5YvT8zrvDBhdmT3cJ69JgU4BjjpwvS8BH0in89A4AkPhPy
dWw/pmPb5Hsm0jBMcnLp2UZgWEQE7YVIUwVi/GVay2FcPvxlTCU4LjD+VicUpzpJ
1RYEdSkNJNxg5VPXWyz6NMvhhhW0C2CJovJUVqVe90HrIQMJdjcxqV4QvYMlkMLm
FCultAuQ6EMjt6xfndgJkbs1B262ZvBXhTqlWT9e03/c5kKXCxMTZmUPxnfX8UWx
9dMRcgyLqnQH7SigzXIlQkAzcHG/vFyvREEBdJGNkw+JKsZAEHoAE214ZghScjQJ
D9oJ6zgMbnUfcsJChZ4YOWi3iJd2FiUfKMRtU3SklKWNwwASCu+k0j5ollrIYH5x
V9H06Jl0TGeWs8q/7CI4g1z+o3qwmANhq6WTGyLQ80J2P9XYbSX+Wb6Rcf+KcwTC
mq8WLh99IFtkg7J+VIuut1y7Rn71CPWPhiWyoIoPzNjWx8uxL+tllb5YgmXvsQHQ
JNuyr/97v+3ow4zlWnYF41FHj1BZGpWZ4Z5WK+e42xztWW6xGaZrJyKoSlk9L1Tq
bg/t/IFymduosThV8dXpiyJMIC0pKx5ZVm5pA4G/iAzYHpu+/wrHAGZ2s4SaKCZP
99C/2Q9WAgTdg6bqwzHAo+HgbOEfWWJKnxtXhvJWzr7n7jz4/yF9cAdeA2pBFR1D
39+u0TZnHlt5W71qlnP8n7OVadn1r/EICmiLuUumoRoNnwp+rN0FUDLlxlp01Pp+
7benq5PPsrQttEwCFwUQiGrbVzBeBEiS0qA0Nw5kP5I0QztxhBxhjdvaxZtAhKwU
H2VQ74CALbCXSZziN4/WDjxCHsMWQwFcuKogrZk8KRV1+eMYakXaKJaeZ59MLT8g
tQv9qjCxhkMCRPeuWiKJGhK0jIZs7grmg9+TOZclHPEvyLfEyyr6ExD+CwiuWL2u
tE2I4zo187SS75D8OMemhbnm0kgf2NasBk5cxvw371V6fo6VzWVa96wx+5Tn7Ar7
Hx3tQQHlBJQEqd/FSTvS8unDzPIfgrOiABCv+vCC3o6A8NL2NidZtgACKfC4S5iV
w+B+U6ewwi1eijetdajNPpbK4IlPg/pWbs/pTcwvc30YOZk3IIclRHO+CsTkZCPB
fL7cRf6xALmEhKYyBUQWKef3RxHkk+9DVgnBfeWU/SvG4lcPRYVrcJBhrzStyyIP
DOlkUjRkII8amcVN6ZlFsLd6FVQY/G0IH9f0NwzmweJRVzCVAzNyTWFA0Sm37COS
aKZE3CnRgAKfayvUuIukCZhRiMufxSrRD3NSh7uzXlcgGFqz1NIQ8KhDIwjpe8O6
L1qS6+qW4dvqFj3fOsZoWruZrNoLl2gQwNmRC0/LV1yZ73irXecy3ETU05cdqvnh
ZkVVXPmE9uXJJR5Ho44nGe1dOx+zeeP9QGdFhN14eTu1RukKc+1KGIxAQxRGZWV2
YU4FlvkvdMeygAykB+yWTyhtggnkkCiiCNjVgpylgKt3VFYa87iYqq0wDfp80zkj
2QXYfivqRntBBiRVg87rmIMmWoYvJ5tn2TnRlwKhvzBiwLP+UrRX2Va6IhKleFcW
cSGFI/6Rp7z3staxhHl590OqgfXD57FbgQud5HSidEPA5atagq6daQwq7TWuoNf6
GTmD2jioOWQoDDNJJVMQCLUXeiIwI/r4vx7L+8fZwDPL2Vc3y3kIkYFQDvZp+JK1
qjoXQUjzZ0LqNgGP+DQqiCIT08p/pcvfOSnOSAtyInlBKIwAdnpA6NKTtzZHCyEo
w5BPIBKupOuLcLafVyD16gpM+OA9nsf1ta90XksddNJhRji8BCpaTJ/Ql58YrWou
xvDyMkYERQhH19MvYrpBf/gSF3V9uvOzGzyQskWNhFj9mW0KWj2Eu0nTbECxYbH4
zKpVgXomI1oVL/i96otJoSjH4u2m4OfEqQAbYYlzPDsJoyPkqtxLyN/u+9PrPEqK
5R+tIzAPMi6pnSSGr7SdnAe3KET/duH+Fj0j3UDhb3YMdScvQEbFynNevpgvns7y
1d3oapwibag9xbTSqKMnxYppRcmCODJsPgwbEXc7i1TE5fAFdnSdW1g0/3FFBiTO
xmDhC0UEeircAN+OpQB7Ir8IPI6OEzGFc9qQoxLdWvvT6QtuKFnyg3p6tqz6o184
aDEZxLH04ZCNFH2sh0Uc08aBNIRljuY1gvunlsHyURP9ghbeAFTfeVhU1pnblx7K
mnJD4qB5aLCLjNFsfQMtIFMH5CfUe3ETyLc+tDuLuUGtD+NlAL2S5B5I8aeaRxYn
6c319SGiRnlMYldugRjXITkCtpRaT2V8Qgrwp08AO14vasjrVHcnjsnIkOuX4L2Z
PrDpiaMAN5Dg2cwIkLzlDvY8hgUyRhYNZ03a97G9S7Ppsk3nDu+7/g0FVAcymFHv
e3VUucWxuwM0eqw8hsq4u+14ApOUC8Io2VBFXmFf9SgNUA+MwhHOTsXIJ0+1Hy8M
2QBXYAHKrJO/k8MC9MU/VKPieDxEhyR5sYzg63kL/kbZYrShYWRh3OZZR84r0UQQ
3P4CtxQJ2KTRIP4PhgYld+qjoCHeWlJHphv7sE1+UBooUuIrEWg36Yd+0RnmpDlp
t5hvxKPMxQej11Hp+dub591wSsfhioVJzCkWCDe0vmRbgaDaFAp0hmQcYZahDZig
CmRli0PaPli9T1UGqu2eYWIouAu4Y6Hx/Gs7/YNbykfg6T+FLqMYfZDuL0ct+X/q
GL/jEdQCjX38b0pp2mDKyl0zHppDYGmzyfVSsNOjMnkOoiQAMRyIZJDUcxOR2zK7
D16R8QSsHT/iWrOfOFLhikwDfvEpsv7dtCBy27km2AbwY7CSUTbbXyfC7A+Fevb0
pF05eYchABU/O7j9tLhy6U/CNJyCu3m42uwP7bAiK33sMLQyMBXqEZqoMw6FMVbN
yDRqAIqdNOiewlAHt/LmxLSRLPEM5ht1Jb5Eq4nJgYXJJal9V/Y30HFy1HKdBuUB
QcgAUk13HsoMvLwd1WQeoFebDWwp91dfann+SgYu8J6QAJsma//mLUosEGis5XdC
/UanbveBNUtYtP10g6XXuW9kFN/AsLKj/Y8H6HnJIChDa5LdW3NKpH7Nuq1TtFE1
Wp9k4CEUl4BNbOpnAg2c4eox7NNz+uopczjPKSDTyrgJN3h+59i13p+eE6xs8698
82izR+ipsWKhZvRF563kgxNLF8DVgPeW6j71wUHbIa757EpTyDKGsxTliNp2A2N+
zqXaumln6o5q64Tm3/yZ6FE87Mlq9NKjI9YzH4pUe1whbQ0WS0CW8rrLbihlSKX2
j+BI7/r4MMfLo4cFg/vjq2/fKv3u/9txGudEdaCV0VjiVV6Rk0+1ngOf46Wm0dPo
51QjSb1sTdC1Zsg/I8K1stvQGVtjOZOgAFxQkM4SIk4YYob1sk8PlcL8sgjNJVqX
W4/q1jbZ4Wi51mhHDQHM7SPdlCN3L5wCVKpvaDrW0Wer7VocATVUgx1/zrFZhQwi
rkwiu4uet6AX3NS01dE8HeiB26OSNYR3Ur7UcU18c8PTPhHLAuEL4qiwU1UmwOjp
t4qCG2eCroME1QWpB5ZQmM1oCbww1vXz+d7JC70wQkH5OsiyeLNi+oxzs1GVlafk
MdUWVKq/kp9MQBg7a2D0BFQFE512ZSqEy1ubOwW4Du8Wj/PsQYzCdroK72Jz/Ngj
NRfd1PHfeiUfmJX05yWxhcawjVKySP6jB4efEiDA081fk8JlfyaR664J8+iPYNti
6XAaGxlsZ+L+0orjYM6lSoG+jAJUUI9MjSIYTXlNjHi99bvE3TRU0e5vKgmvXJ4S
TqeC4AobXPdKNTKPlFE3pptywGhkK2R8wt/CrzBazm7aakdRfCRbrQYbhzqvqM63
RfI1WElEjL6NztRwnEhYqtPLuDqeXUv9zIPKW+RKn/xEfC0yRv5X/raOcrjPROSk
S5iFg79EJSybX/bvhYvAbG+nYoaUZVe4pz+lyVljriDm307152URhQf53MN8hjsv
tBl8rRPZfq9z/M+i2cMDpq6CgtUqUdlNh146oRucx85Yflht/XnN6JHjIr9oesDb
01x9hhaXMct+ZDzOqEF3LQHhh4OX7tU8D9usBCPFWq7ODZceeF74RQcGcnHB8YIA
6c8DbPoQcPLVQIoSrVEpOQ2rlGxRfyhF/EiE6Xxd6LrwFJyJsQY3jimS4UEL/O2A
Iy01a0sDlb2rh/8fX6q/l3OZV8+73lFaNAjIjut4RjY66D5jQZzgIbLPjNBOM1ZY
H0ivIsK6Y6vSY5sWZQAug5UYgp/9mZje3W0b0N0YA1R8fVqdvus4sWTxkbJNNX4q
Eemwj+T8Lcw/6ugi5CkQ9K5CwZDrV5i57NAfmNLDsKwsFH8H/cRTFNfjAreEfKdx
sM1RqfAxyckDfzBgnIf40DD+clv9dc/NT/sH0AubtOHhpcvwChVGFa/YjhzaEGft
93hacLVNHP9bOOpEBKlTecnd6ZdO2Chp64NuVY3wWXrHckiEg2w/jxSCBt6IWCN+
Jqv+lK1Cq8IDcSQCs1kku4UmcXkQyVanbLw3//QGbazCOhfT6GWbnzaPFhAJQ3hO
syaNuHU650KqeU/y9e+YeCOQPHJOLnZsHwCGSEyK0IowA1EB19gAetUMQXLaUAQh
cSHOK5lNNBRdeO3Ts1Z6HA+L/gJFcrSv8hKBLmPm9h/Vs0IwMsEcPWo3MsvCuc9B
84Mzz0XbZaxFFGYhx8NWbjpWdPkGEvDeUcoobX9bTytwjGAcd8RrFR3yi0/5Wsy6
4Oh0739GeChoIWvx+il9JAHzFdN55o1uwoQA+jWdjVcQMbXA6rySMyHTrNH8y73Y
mCXHkfwurFXtaTCLC4EKo+LrbZzMH4jNuOLhHLt/zO4+wtL3+cjH064sVNobCXpc
iEPz61VN3sucgt97sPdYmq/NRqZgyL5s0UHwikq4o2KDXRfAMA0kjSwjw0Mq3Z/8
GYdlSz78YBhN1HZyvxhtsV06pfqVefuhAtJF/C1VM6XMIYIJPN7IkYRRfqZs5/Zc
hMoZM4Ur+JQUcjeODgSqfSqyItnsHVFrZJuGB3tcf96horkygHyqvzNhMs98MKgu
qUnY4CdD5OtK+9aT3gSgourJBXIoC4YjgkNjjYMaRryFIve9WgFqC67G3Q+j8y4D
Fc5gWySONHU8G8O75l8z92eMsRcNIAO1BbIz0VktOoJQAgPHpnxBOR9uYrO8w6tN
WxILA/tcSodDvObacKdXY+/w4sueIvXEbwutV6nLSRXj7X6TINdOpl/6GMkhZJEx
zXnZAKCh8qwnAjWRCfjnKVmkW4F88/r1br0dsOLxY1Bxh221P15/kM2uUYzLh1bX
tkDc81L/+d7JJuBii1txEGir8La56V1Kz7hPDSD5cK2WBIME5PXTjWvAu46rDHq9
/2Oc0cJ0c74Fc6vnelUAnPBa4Og7WQ4rXvv7N3iEBYtWvga8XuVxpeUVjMExUaoE
2ucTUTAskxEbjxKvqVhJShPc7Z9Mr7U6g04iVV+QA2qSxXcOW/xmqn9w/Fh19ri1
qvSrGp26vSn6Ec7pFl1UUqZsZv3GgKiu03k/K2X3cq3+Org7Dd1X6MrBlbIl+Dza
FVd82zQwr0PtuPZiO4MchrxUXglOSwepoer6YXttg1qTpx1EX591llfDwZPK6yLe
3OITI9dB4oRCWB4y8jDAP2gl4usY9Bd6OkQ5ZRvM+V8lFMnUZbTTnG73IIXTG9eJ
cgIOZoWhMRyGkWgkJFfasLI9cIYIIeFcQxWHJPFIUjYWl0z5A9mkLdZrFsc+Db3q
ocAHb3+wzYjjUrzKbiNT+PQwJseGYg5QUQXJWuOJcp/393T0YRmIgFz3ulvFTgTO
t1NV1j29GI1M0UalIqqNIMcWTIVo7xNDhJoT8/GXWMzqY8OExzvQsX8P4nVbG6HV
jmCrBR67LvmlANN86H5qzKZpFRCdSdaqhm6pKXM7b0k7A6ytQAnZEP+fmqDR6ru0
hNLZRbiQ8sJh2QywVw+KvoSc+YL9YvKGjYwod45xdaBR4M2l7KdIc4HJjAjBJwVw
giF9lnR9PgsJ+WWv9Z4tEm0c7TQDglH/9+us0Br77Gwn1c7fXJXx4cBHDYKFzq3b
nyMVabmVdB4D611v0OGPo+kQgbviBTfbMqk2eCsQiZ923VRzxQMU+2XlSbzDyPIV
Mz/9g2wAjkJsBmwLN3d70W5b+kIPO/lT+0wmzao7zxmH3SMGqoiVhBld+4TYDfQG
DBYYfhbZQX5m0mqWX0G2vizoBa8+eGQLD8WO+OCmQOMrKs9EjpO5TsuM5Bl3h0gt
adnCyQHu7QOhEyqsxa28pJ70APVuL0eSyX6VXrPGWd8ZxCFz749akxTXQPU8ltyP
mZlG8csahJCy1yyc/IqsDEd/y8iuxI0g511+JfHXP8UX33gJp8jaqeqsiCOHQft2
96/wIVPbKUlaB8lbBmmQ733P/J94iZUNQR54LJTa/5eDT2gUMaAe/70onxBURbdj
iacT2Zu9OdI7TL1EMXP+m6TFUlkiGnGv09CUsiRf0YvvH0/+gftcQ+upQum5/6/o
wMXRWfBP1ZNOeOWixUCgc3bpM5a3vEwMvselG05hM1KpCv1nhicc6XZFKO++dv7V
FgC+tNcQlgKoMi5LeB9+5pfwVnAaZVSkFLhoBgG1RMsWS8dDzu8r7aEhwU6eFaSY
ye+EkbXYO+IGjOl+6ihjpiZ0lZfYtxGDnoMDMmxoNenYY2aiZ7QvCN6CMr9H/Pkj
yZMtS1mzN/trqNqYkjOclQWxgB/2eetM/+aX5lOUM3IljcOeYBR2JTSeTxWkv98S
Hl2x8OZG5xTt6p/Yhd/SemPtQNuJdicCWv30YlVm4zzk3AsSe6/J4AtTbZV+314m
NumXnTRLpzDnApYrQ+tAgIsjN7XLaEYjFpSQTDpmyehaxAHeHHyiFSCTPfXAIC6O
vTYCw5Zwkg/cmTZ26kZ6h9hVG2R6bxKRelwaUPcPYYrkqoxhfXwzqmP70Sstwvug
5BzpGbiC03jgmaCPUa79RLeoUKL+BZf04JKJ6ACCut+EAhnSIy9tA0S1Savn9aMt
3xEU6qq2K+UJMJdwaeUNUOk/5Iqh7BNp2KuM8p9fIuTJUwls23YqZsnp0fIaI3rN
kv0P/pxIta/erH+v4Hf7lb4dZGZYzM1OiCTuuBmVwBE5zviFJYFBIQpul7gfrEzE
Zisj46qzyxIQh4K3VMOmJC/xXAAIj6zG56gb101rzYirbvFEYJHilFqnhtZpwxJd
jOkXm69sr/D22TVo6riyoZGjur8cEy98mEoHQnmWwqYeSKfSF11tpFte9RwNnlZG
peqQBsmlMmup7WNGseGMSTtJ83JY7Yt+mCUnT48wzectNa8llUIY0/ls2YBBd7Rn
LC0K0pKcfwkL9qq6bPg0ZayubPgp1YW32AQT+iXCJzH/Otsr8COQRvL7dQSD1Lc1
XBZK542cuLJJHqJI6dm7wvwnWfmBTyOj0SwlPVmdugR3ENabd0o69eLVRHz/wxr9
ClJjGCx+N3C/8S/auZ7LwUSRktvdMnEINXl6CEvN+Dm5rjUK7JLWGh0/mU7we9wC
qYeneFlVebQp8qhc74EkklspgpNu9/wKWS/d6dI5t4X+rxFrVjrvGGHb6pcwbcZR
lCSqlWziypp2An3HFY1KazUy4plM3fjSNHJpm8khRI+hE+qeFzmGPpZSsM7QV5ln
iD3HzvptLNDyyZ1tjCYMQpdxsKTTvESk7HJe43fn+P+p0dEGCDxGOzeWDkymjKNK
JTWDzGco4kcyPDQjGiH3N80YqVm3gQ4NV+9jMIj/pzpp99LMdID1w1/V+D4PiNTq
kdYhPtFq+H5VDm2C8nFTW24f+dctB9qHXY0PYXMJcfNTAJ2LPZximKR0//dMkOCJ
NdPQqAhM21W6nKpCs41ECE60enIM+xBlnRyyotgvCsyBDr0PijlkTnLvehs2elX/
Vg3iWH2XVrPjgQH9tz2gPN7N4tKOflysAXataU3z2Zr3ZEbw9Ua4rMWW7Hs510QU
08XltOZUx0XkQn86RY9gK6OEMyDxzHXULODaxOfmBAa2QIBbqSsiydwy23cBwR+C
ePVeSQRK0u3L28sj/9AdLhRIsSchVBEqltgVg7fOOVZIl198dzd2j9rN1RJ0nyYy
1TrHwPo3i4oPDoAhXjfECmJ773o+ardC+bSes2PZLX1eIlAGz+6mvjteN8qxGgER
uYY9zH9azQ7TOzgrNBRzwLJzXkR1CYUVnTwWG8rKn0PAYJ6waaP0kpHa6YJBwYRj
TTz7jdhuUU5CzuPSz8LJt3IBWQse93jAiNaQlhVHBcX4L5KtR7YUU7TQ2X9kyI8O
G5QMy8IXVc2udfVDtjx3HZyYnS0SFvpEDK9BLh8mDXvfCWa5yE72hLZwkU9UmQ37
w9+e5CUgjORimiHbDrYUJsPW8uGMWB4s84E63DBqAHTnx6XksJE+G6VmwSJbM3CE
AvC80bZbzAbFW9Gxd9tk7Z4ABqLPxRI7sABCPkzzasZF/xy+JfH1hghM9qZz3BS9
mhMLGbHujnDX8unhLKvov7gCbnan1ozs7mGoPq45mF80VYrK8F0WHmexrMJLs+3o
ri7W5exRMPy3RXyiPnRUoh+sWuT4qq74GwQL0xbIWEDQgyuDEucJ0km0TTPsuX9z
NciWlO3dd8BQqaPElTL/eUOV/FFUfdfG8uTqo+m6zUWu2w7PBSdk9y5Vr4hGV0FC
csuuvr1RLjSygn9Z78Qjgz6uc3l/diqn0b5qq1zPBPjdpeJP7UPPuXmGlWlyc1ZD
N1cvGJi7ONhBE3EQpARy0VqMNW/5aecCR0NXUNBDInXfMBoF66rlnrBATGZr/54N
vQPcWKGl9YjOCdOm4/KMfPSEfFUCf04ANMAj8+7UyeWqG6l9MmoUdyyx3nedprU7
a3O2/IB3PXADJ/wgUHu4nMnRPhwMfeMQr+2rk1ik3ApyR9KOVbkoGIz3X/rLul+S
97NHhdY6tv0oq5C+bdj7fU9C6lAJoWLKRffijHVMIDjei8VcozPcMCKotgHil6eV
7jg+//V3Zh74OuKQiDLecxojmHa3kea/ql9k40yvtgmAiZ/iDOFTt58CLNh7m1RC
PSKR8PBjjHJJf6wQveQ9XpkVpRNt1x/HEAcovZwAvnaLWYMkB1Tqu3Dxs3AKAqCA
KZnW9mayosRCHYbbs+BJ80w9Yrm0qbage8R3pKwuXAbSpHGLbDCDpamZ7jc9tWvD
xNUZuJOTpmaGOpv2dF+uG3KwR5N4P4RcK/Sluul7Ejec/PLlH/emSewTM7XgELRM
3pM0VxqJUdEoGKOi217m2qPdrzsxXjuzI/qXzezzC1MloCN/kmHEeim26yxThT73
UyIpkWCHO29WVMbXBMOGx1CbHA62GG5SEdTCa3toY9ZoJ5STwF8om9gilDEdVfT/
lmaVTKu7oyNKtI9GBcHphzPJ6hIiSHjHLtmRbAZlcP3KeWfTyd2kvgYobN7HNs/N
2wxg+es2NWtMznvg3krLAudffgI7Qr9RzH8ZGWoel5ddBstKzSYHLDVhdnBaRcXt
mS7epu7kehqF5mVmA1gokKKjhnZcBu9O4LCaB3le45uvHNu2+FdvPNf4bVZlPgr0
fJvkQhZrBeR6nwYWrJUQkE4Z1d6I4lu1Q1tXsHS0Wm83YdzV8PuoE/g5yp4I7Tyk
liFlpWsEN5OP0zXpTx2YdgveFcgGFBQs/4CY9PihCU0o6i9Lk61ppgSP8+5Vcuxk
+W0bTBstAmE/F+x9PMmzAOF2meF7cEl2zEI6NlVX8U07eh40iGYjE/ifj1cZHY5B
4mhWONNP2eqGnk8KgBbequgI6M0udk5a9fFlYmVbxYMZRQ3A7ULfx3/tGLHKpAbT
30N0whvuc9cT5mHGaw0rXUUUCC5WjKLXk19AGlnl0vjPkPD+teeN6haFSWOBKiAW
tmELiRyI6qt3iDlrhX1on0yfPIH48iGOEkS2UXrvrBksTqhGju4rP4dqalg/c/gT
fTIUDbdYZgFfXsXVJQTdXje5Tv4r9kKpE5xH5ZzAeZzKWDMc0zRAjliErkYsDUHG
1opllERVedyAT4naAFt/Uko83CC+iXEPHs4xpQiS9To6vqww3NosBLxhzTMQDUJA
UDdfvungwXf4G36kFL0vksjAGbJzJGTC6vaO4xW7z/AfbZ9+rETIkjX0E9SPOmKh
N9T9UJ1Tzd4zgN4R63cl+euMwqPMjBP9INAbtmsXsHdsKM1i63iHyH14xghU+Dpd
VSsSCxv/K+KvauPol9J+YacibpR3KIanRMsS+/uw3l1we4SDU4/Rx8fw1Sw1bMo5
mUxqrq6o7W3TpLjGLyLKB8xHY3yjg5PDzbSPtHj22FBtVHGAdiMcDbVbj2PzUKks
eprHTh8s/wXpiif/8HA9bbuRS9wt3kDRGoTbZ6VIK6I87RopKBdtzbqnq73lBDHB
TJ4F84nXm4VQhbprcoUkbN2wOfQ7Xjn18nCqHxfDGUpbJok/Ck7A1oN/CsoUjtlv
tAAW672ILxQtVh8Ioc2levyLvRN1fxBc0qHZg0ej/S+5LCuNTcpT5Y2mEnIxFKRs
DYTxuRsKVBPYgOgTehH2FtljicyZ8ILFMffc91pkhOxi2KKzrqUP5+Mldwfq5fw3
BJI4696iBfTuuql1/4NhKcP1mx5ZdO3oLN2m8w+8ZfV6nHEInT991ZdILGryDIDo
U7XKI4jdPUaojTnnMoAkws1huCYpphT/W7fClRWTqnnCydP7I72aBAR5PbOvCtoY
LNOcE9AsuoZv+AAN2JmnwaGM5hvUybq0KUnj0ZMCGk0m+VGMawCONp+rqjJjOLGz
bFBVpmnT+a3DQTNY8IXSCFxQ1cU7A1mov+C9ToeOYgHOjll0vTDJx06962KUDHq3
cKlNpexhsMOeto7fR4jnUPZ+s37xSTnbXa0/hiT9jbjg/ev93t+xpKG7BOSEoo3/
yuEucT4wz/4p4rwGZOKuGVWml1nGmi5xfPZvWyiTokxQMoeSwxG7uUuTnaUOF16O
DguGfPgrESp9WgvcQnPoEKuSEswYkQg/8Pur+AOz9iBxEa/aNgUr7pTv7OdoRNMo
1M5/RI6JtsX9HkEI7lmA8IFT5/bLOJBfHoDuJHXi2g/HzXHcS5oo1gPFsZHWRYss
d5R4GTiebAf9HdeQsoonX/pSc6rNBkkPxjX8jrhyp2zcBvBCYmXhng5Ub1zy2f9W
LsBSeqhwxyz28reQcpembouT1nLGHOMM/YhF5GSPLLhr+sHG85LZpNHQ+DQ3WerI
VEmeWQUA2Tmi1yODVyThWAv01cbLPX2lD+0ZCACVdG4WxpzP5Ipk/Z1s5wX5YuMB
O8jxT6vzfPmnYyICGG/f7HKoMGNhTSUD2Vi9g6quErjKJmETvvrWZ231yyDpshvg
HBt+/B9bAe6t52cvt+BmclINPNX339dHZm1KJSGLHvkpZBpKJ3ZQOo9WagnLjPMc
OfzKlGo70lkxUhj2LfzJPQWWPdAN82+QZ7Cyz97KQ6qYWKHR6gnj+LfvHDSHL+7U
81f7iagOFGKXQV7dI+WgWtbG2AKFMqWPkXUYi2ol0+Hx9lLz3JwCR2GrZ/02E7Jz
Cw7HCsD6nNWXLJj242JT8LTNi+QqaeycQzzqaA4qaHl2P23BttD3+3qjhyN+Wc7g
n91acXzp1jaPFc4/QCAkkPz0lccFDJpB8ljWY26oUME6y/iUWxYIL9fd6JBTVQpW
UlUjSiNACJEUGnUsT/7XZl2+3Yxi1hr0LZWs4cgBZkDYVdzy//RuYZYXM83k8t6w
PTl5cmHoIXPDpWvp1zHy4ub1bDoAXq1ZEYU58nShO61UTbYh+2rRin2ssg4V6lvf
fzEQjznkXtdmajgWil1vMtDp2VizHhSNtxFXlIUv1kmuPhqSAydgGZaEInh3oG2n
alTy8vMM8/nsgpb5XqB/twIO2jyYh2jVKnj+S+eY22JYKJ5SIXSqj3tx8fTPxbD8
tjdTHC5Ln8xeO4yCtV+x4D5JQJotqNeoX9JohmH0EPw2h2HPa8wOKZqXE/pbz02Z
I+5Ae1XYxWABaqc7hHx+6bHbT4IxKDjGVB2Z/cXD23egXIJk0SX9qn6PeaHtWkvg
T3jkydsGhybCzrJ0ZCUH//VktDLB4+GTwREcRKo9Xgfj476qQcMDKdjD/pGM8q0m
YSsnbAdhY01DKdccdkoCYtEafBXE9ApsCOckd8phRIC1Ec4MFCT8gUdWUP30DXWS
Ej3AOldxPl7l9bJ90YonBAr5cWtqOZkvAIW9/5kUztqqIUfIkIgqh33t1BTVOrpo
KWPvOpaUvLQpSK5sdSPiuswMlfS/N0cz/y6vqQtVf0DOH35VEMTYdcOhxtdzQ9c2
et+b6rYxiG2/LEeq2MwpeaaWSOoZRRv5dLSwYyaqHr0qVSRZjED9fJ4z2fy6eR5H
ltcljSO2mIWWpPzQlDbuv/AuJ/atSJv+N3W6S5YBEJ7cv8t6xeBA9mSK8SkzIK6l
u4DsD551MOuxuBkp1fs8hI/icCT7Dm+D1aBOSXZjZvf8diz+uA7NmZJ9wVOaESP5
tRBV1L8Kr0uZNDQFz+pkforsVpoBpvWh1l6/nNFnMeSAeVGpAYo0gKDnXg8C39aL
vBDtffqtQonfnbx60fhCXOvCfSMwCVOedCqg+BnY/M6Vvi80F0HtCoqQFJdADVe0
91Zg9QCHV5gaFneNUhmeMDEqPwmLrK+950dcZMihyTaP4qCbKKdfWghJpjiZLN7p
0eWTfvAm3xFpRfH6r/mQuBi+2oQHpesaHZ1sEQbCBG1xQs68Ys6iz+G2x7FIhevW
j0xswowh4FDEPIT2tvytI+BdHkrrPuu02Pbaz6dOCbmqdR+4OJE+F/eKTE3GuZ+F
3oZ9GoJNH4nQNL5VFaXwj9K5Z1P2CCb1R7moGgXcJ92b5SCUMCEdGr1KZHQZsD+p
Wz/+MWK/qJK0+E2qLE0KV7UJkCOqcySfm7B55VctG1XNMW2Ow5ban/XYwDQp6fg1
W3PptpHnpivG4oFPsx5R4McNCSIQ+vNWSE5j0zQ4FxO9uYqgz3SoiW8Q7aGWRpTB
HAk4PLZ+5z0bHkZ8juNvnhBd8NlRvReClDPmPmFbBWdBSQXHKfQl3cLW9ZKa5Y16
G9s6YuPLRUNsxZo1vATdkqZQRc+qJzeaXX9z/vmL5lnkjiLgZwD3sSlRuThdLTh4
JT+lZzRHquLUlqdwqZOFfmEg3AG3wkx+QOiBqgu+XhzrXerRvXCo5cipivzY5s8m
fGgh68hBtYlFAgJyzldYdgBeoqQ0mfu/jRBwZ7OoYtORiS6H12nHjfAgTGoxNR3P
0keSPEpj3LJYyiRIpc98juvFF7nUjLjyHpNDlCyeaRQ4fbjKJk3DNsYP3XksLlBv
bu10n26J41NPccKTWftkCZ9A3u8K9lWRL5uzrbLRs8A8RRrIsfIy+q2IwAfWSEoD
cSSiTWIbHiI0BxR23Uje3b0B/0HDe6zvEPu1KC22m0YNzNn/RDUn4WkmzyIPU3Vr
3tXsvTS3+d4swwvUX3ady76mVXiXKAg6Ibeb5DsppZ5bWlULhxa+wn8ZCYBYQGaP
jvwWD43cl3L+RQ4wPoW2ifu4t3kbTN8OfKrLq1XDN+JWu6Sf9NJak6SJxr+XId8t
bnhvaGKJ51a2Z5HnRWgPgSOLlLoGrimbx3enisJ5rVXAdtrGCbP/w/PFaM8dY1qt
2AJUg4gLRuXGXRVaqKvahWWTWQ6qq1Cb3emowiG8IXFe6lCcihPdL+vi3m92lZw8
CEmRY7/RYq8cqdGcihhsf5YzMjrBVhQdPkI63Ev3M+paam8zEy7hWJFWPa20S5fN
5N/qooeQiVHPCHB2AWMr3kNg3Y+H98a6Mb6pToPK2J70aqno8EZDWiilNKozX9kv
PVDx2zKraYF+CMDtU6jmAUU8+Pl1YuEPiUOXn4ACITLydUecRlACMt4jLd3J+RhQ
DMWkeUvYU1rk+Dwqdz+UZAnHCSeTQFb0Xp+jV4eocZCigs29DDDrOGT1Lb5FjwFp
rdAUUyzdKDGqAbuW+0w1MwVJZ1kpBYpx7llhMpGLgkNfSITB3hqO7GCGSF6z8zb8
fuitv2jMIM1PaYGKoUtHddgHGalRx74njvi2Nf6f8Yt8LtDXuF10eQAmki8aOD4w
1bH5WlPPd+KN2tbJZnEp3Q11GyFFKps3CtXL1oiX9zN+oJgKIrCg9rcYrjvytWHY
K52hxHF4jsqdDqC9j2ppVkid2PZg9Tf2j2exLiEcMNeE3dy9THON6go4hfWGV0aT
LN4pzDaffQTukGZYqRNIwvRp7uYZbuv1Wd/0mquEpgPwvw1ZICV8dqmszUCEpG8o
2iL+Lj3GkHKWyawXv6v5EOzjGB3SxzLPSg2BBGuPCvWY5814t8MWCUaLe5EJRiLZ
PvAZj7SWCot1SqjBRuaUsOo6/g8Qadp9eBhf9eD4UW+xkPsSazRl3NzPiPzb3K7V
y5LzbiL+4yNn+QJRCn5rMgwH/RDqa3mcMhFhqbROGbXdEUumjSRvR5hTzI/Hu0rC
7u57xAl4847SSUQo3HVnFfDAfIaJaKx69IKkJ+dRn4ohqNEMpmgJTxLe8KlDOzZy
KGNsRDiHDWmd+XHtW3X4f/Hk8G/ce1sjU2R+8PzbNeD2R1WZKmBwS2KyJc/huPhp
HXNH+djtr2QHGe7Ira3dOimRbF09JOT71qn357YcErLJ7znGoZFT4vIMDxr/pe9G
3ycTdTc0pG4OnXtu8gS/+mI/1k0AWgxHfCGMJt5Jx65WJ3ea269J7OAO96xzBBQo
i5SP1YfbHnj5rS0Q2f8/wTNb1hXB1Gl0kgU9xbDAWsNKOrMGUAQkw9RKMkmDx9jF
epjG4J5uA01qh0CNOcxdzb4PtV5eFBlVekUkm9Qe4czOv2hkU5cgJ0traqPc4R5m
C8GrLqP6neXVmnDqsqjw7hvIFZz3XxMGQ417hIq/r0o0gWSoSqSGQN0v+nQYFoDz
nxoNbl/y+a2Jz9DxsfqTSSEmaCHL73mQ6ylY0SRo/1RXC/i0GJJI/iMqwHaGD4k7
UgXcBP3d4HHsyN1xXoyYgah5MnrOn1YtqsFBnjUsM5hqZfSajHDlyhp282cBeUQU
iqqUdoXeJsaZ2FPljD5WndRgMGC4RqHCLLwGjLhI09WjVVPWYslV4DbK7GXgmPX6
heVB1uXphxIkGoQyx19X8Ak1GOR/eImrQRiammcXAgwCLK6nH6sxJiu9k/rkVR5w
1WBi1sdOmVMvPeeKKJaEZTfJFeJS9wRJeamE1pBWku4RBHWTrzoTpvtk9/spyeY1
6KRntUu7VokkixYkhy+gKsHGqdUUZtkzV4J9uBvXz3uGM7/lgGyQuhnuFaCKGORl
Lql6UeOcWeaGLUXBW/X7muZan7N0h2vpNeCHUWem3+8JiXryUv6ii6wSG/KFY+hC
hR+AYoplbXt4RG850wZIv6VO4P1goH29BrsWmtjd5otmdAqSlXUWpxCQ5kACo4nf
/ZNd9vXGNk27ZOCl20AlC9zBynAx1JRPPT42wb+n+hB9qXonwXWEQSdh7KO3ZAGD
Y7rk+gBGgfXluMPd4kaGcR8oLrZTHvTou/EsBNeT5JJcw36SwfE0FGMdCiruV3yQ
ru0oQeuvQtEVRdL8jhYxoo8ATIaHnw5RKdGnpuSPZWbxOkDGCiMOewYp1JVGVSD4
7QSBx7hr6marzbLZEkbUMucrJdXMrrSi9LfwjVKHG36YP/a/iuSf9oelVXX+rOJY
qZbWTpQDxfUcPPl3NPrv1SJP0/T2SvmXov//n3BybT4o5CexQKwZJu6bGSoPLEyk
/3q2tQyF3pTnlrNGNPOEJ31pnBnJIxSdeCXNu2nFueseFOc6dF4Evn+6UkVuItS3
SYGC4azvaAqibkQin3FKQOci/3rrGWSBefYQLJ43BBJji8ODu+T9z3Lf0MJ50wl9
QHnXkWzf03xQ7ZC5hpYQzw0HsrQqV1+MObXKOaq4UfvbRONnll18K7pyWAA1Gz30
GNqC70AVsAnvJMAWeokq5N1O/8BfySOhWtMVt3HjxpW1ZFS9l/J+TR0CFqY3BPVm
qiUZIV2AocYt5yIKvJJgZje55UxVvYjJbpIUJEvIUPb6573+uFPAm9Q8YOoTQMTF
5NCYLofe3QRV3x5YurOubTQ9rIyWrWr7kgLm+S7edadDBrA5Q4a2+Jc+8v3rpMEP
ih3GA7puN2x++hbrfT3MwIR8s5kto2J23U9lqTVK8RiaGLkOSYGXwxWxjliQoax0
TeO0FWgBArKATtFR/2oH/iy3lJzQe+c2xKzLEI3bkLYyrFAePNZ/RUIwygKNeiTS
06D1CPisL85qnsdkEb/C+QlDXj06NyXGcx26EZ/WurQlU+nnK+sZXUrpv3jkcYgR
VbIGF2SyrlXGCrR3DuQaKMAzrROBcHdsMHXc4SpOYN22SFANWZQZNvl7BvNWn7Ly
QJdSIzpI6Sjx6MhqQOmP0bGVPmOSvLPOVgWi+9d9mFRsb2DJ6v2PAEPfBGs8E9Fl
9JSPeZ1Lv2AHJKp/33laLtgZ1PK8/TlxiL8UlA4urxnaoDgkLrX5p668gfGuRfHK
5SOc3j6/+V3dEWRzzPAurqLilgHYRPNWmhyx+/HEfH2TziTUROZ9RW8bsACHEbAm
KB/4i55ejWd9zL5bWf/w5YcLrg5bzGoTUMgDkaC/LtF63VcCS7KpkyWrPIenUzQf
34zIRv3vlwR+bfmp/aB4VgxfLv+o2fF+yXu4YGXh3nBpM0IQlrMRqPqQm3kGJvbA
67wOK0RH9lcS6E30QINGfH/Sa6thBE1sFv67Cd+gQ5Wwok+WMmbQB1XWQaQFzBu6
BOaRd+q8QRuiI5RxMBPya8wdR9S5l1+QRNWBjY0UW94t6uWc9kLXzVQhsBU/VTGF
W1k4y50zt/WFNRjqFwLR/CTZuFerSDO3ak7+JCEXZCiwR3BpM8cdSJHbRGeQ4qKM
/g90KR+HgWh1FJcFHmdkj5IE+fkYcYcv6n0NYZb/gXKfyzGIahoYPAHPjx7qKVss
aQUkluRNtjIt33ZNJsTcN6JhEpBA3iCe8n0LCFmrrdTRwH2MZrUoJIIiKB7l92sp
X94pbE1apKPOFcTC1Hs5Va+7jJrMevF1+og+ZdFIRvZOuzWio4QnNjELt8C3CvQZ
ghK2t+E2pxVAXbZdRCIczsMANkOQPwBh4Qp3XGyDxYB+D01sqJh/tbEb6q4XwxRB
q30Ih06sf967tz0LqFmaEY1sxe+z8JOR1wbWqJrZrVV9Sz0dM1VMVo6fu6hGx/6U
yE2fd4TOK9Q41hsUEZjPniosjL9SiaBO56GR1BeYyo19y+1ttiiyY5R2TB587rD0
5CPtD8gbq/y03Dy5xXjfZqCJ3OYH3kSer1oURbrGjTpTWe6e6npXa92OzIn+j4pF
7KQzmW1KKPM23jSr4cGkT+YuyLJieypA5hL6J0O4a3UhmGX7BN91Wxmhg9VAQhv/
oAT/70FD2EX2KvqTTUzyCLKJ6hfWzYAK+4Bm/n0z5o2w3iplyTq/6rE28cm5LQQ9
SZbGpmW1Fli/j8B1sFHqrj3BPoL/vb2DUaSrzoTzvN0gUQaWM56TmjK1L2VsQ4eA
kD3GZf7MxwpVfioeUD71enFNuhP1mS5W6K3TMZAgyftucaI6hC++zJtufa/fIuFm
Q1z8Iu5X5tOFI1Mtbfd3/gdq0WjeMoGkr/+SzbaL9ljdlnjID7gbh5bd568HUhMp
R5wFWO4aYxOpYsf1QrYmd+kiVt+EK4qCGA/zpXWDX/nqcF38uudwl2gWkFt3AzX0
HF5DdzReerLCqkYcQEH8stxiD1hGDFakpXtfHq+4ZSI8CFYrWf87mYzuYok7u0bI
tyPbxHGnAA5149/7ZIV9/tyXvnoyeXoMG4j+KLzsPGfHTsFt91tGMrWUKcnvAp15
p1i6pCVsBnauRTF935sHlQOWN3ir0VDeUigZXRxXfTHU7fUhDQCpyObuAfmxm+HN
KXYSxKnhAzZqArxXhk+NZDXg+cu4KTjcxS8chS0c+8+aP3v8X6frcGT0bWPgejay
uFcLSW+XoWHA7isg+psEXflvGLWrkIpOIdL2NAV783Upe7ODlK0w57qyZK5Orfi9
j9xlaWRwpD3wWOhvogfQEdZd7USf+8VB0D8Hx/G+KVZVq13ihIt7XYepVB2zAr9k
pC57zCJxLEKjHVO8CyIUwswgxEN/vH7UeOzmdN5dX7u3W3c7oXyFx7viGaXc0VjH
88bUt6OTyTish86GvZZ1r91BuOE24NLmfm71vaAK4T1IZnT9pcHfI+8qbwWyfhBH
gJYj1jdOx597P0zpJKC0YiMG04OxvctyUHXNEVLB6k4FmUwZN/NHXy56J7YpObH+
NjTpdcjz2ERTk7LcmtKS9tzEvp3CdyAT3yFeBeM5aMyU2QJMgfM79WDgt4Qhgnv2
qypJYI+9+FF/VylSfSGl4MAq47BshQhYZYvqUOJIZk83jhDZPRKU+r7HdDt+gA1y
aekwMeIolbb7YWkIh2AQboRi7PoORV+fPwjlALV90zeHREzfGZ+U1bjWMfHgmQ/4
Vaxl/nBwvYsb5/zH4JHHM+6u8fVHIrVe8y3J35BXRYjiN1MUMnHbz/SHeiU8wwA2
bvOMtj3ZlV+lkjdpDfyKCLgKd4IagJAzNhSGn4lZ2bj3cmwiO3HSsNcXPd6NKdW5
rrgbPYtnuU2v8a6okaylxIGQn7MdSYwS7XYIzIN08Ig1FJYFIS7pqh9jZKzpRyEw
SujcHbjIg4mwEW1J16M656n9PWCBD9iLp4BcJQ3F59wAqz5ZMaLFQxwK5HsnJQrs
UaEuA4qBzLBGATeNceA8Z34+vBvW5XmDK8SSYh1oDYiRiPgbSzotgjWLfXfSW7Mi
Jrz1AgwSlzmq1OsuSLAxkfqKhZvA61h3bmo/Fm/reZ3n8DAt+2p+6b5SVtyfiEhE
S0Qn7SzijvPxAvWFJB4kz1CyULdcm8fTE/UGuMSlO5WeWKU8p/gfqo2zMZFhAHBN
V/V9m1mCfDeHBoCK4QbPVks1+FkNuh445yrXz+NHxuIoLxu2+Bh1+pKLgMHr9R0t
5f2RPyd9z1OgBEqYQu5EpqxwYb5CsFR0mFISHVYZ9YLOp9CnImY9vKM5RP06p7xz
Uzfl9FOJ30wcx3oWsHaHnRJeF60SlxBp5/ziYw+YxmOfzPvQ7h5W4j3KXtFreztv
M17VbKD29RzRn5lfq5bXcG7Vf1qPxEKORtD96RIgI7s7yOCjGWuNjz72JBC/0028
NjhXbD4+QXJOlH0wOUShRMl4Xp26j5TuNsaWB2FRx/2lF+XtHxZWuOHAg2IT3MLg
JVjlRIOuYEEXQOHAknYHvbXKHBeI3RMWg6zXUBsHKy5/U72wu2v8vzzqTxgXyzK1
+cmSBSv5F9mseBTo0vOvT+hzU5q3NydTTliT1U/21HtE3/n9lumJP0ABNbEdVkDH
sQyvaKzezHoOE/4Lp/vO71Q0pEsHm1LRLShHGJY04OwBU+PW4ymPVUBn7SZ3JaU9
WpmNc+X4nh0OvhfJV/JrWofdBTj8esKWSeOaAH9Up2o0HiWECYia00Kyf+O7MR7d
g1e19A5wh8CFKbUnuR61ZAFmRkfwv94NCO170vydU338w+3pJM5RJHRoqsEbmMnb
fLm4OKkl9ksiYjvpKFo51uUbvrE490mnvU4BJOA10CS9trFqTy7ZgBcQxBd1ctb5
HDRZfaMX8M+isXxFYDmmXZ1OLh7D7eOTj9nATCobmE3J5z9QezfgZs1NY5la29Fo
yVRT1i7h9A2mjNhKQWLZJooCLjANuvcvw0ZdPa/eJpkgTPuYXepmE7hMCU1UP5FA
loXPDI9Hw4LNSkYi2n1CLWodbHfA7IihA2E54lkJO6sRiz4q3oi+IwZxZ/Tj0TpG
1vVhE9lKH70GA6audtEr9JxrXqwFnrOlm/LE0cJO2OGa8tovnlZTPBXiuuIgzm3a
svGUBccvkj956FspjnCKwMDrJrPY6RyOL5XtRCj9FyUD1JQUdobBCwuViIX6iCZ9
0CP8cK7FcvklZicptcf6xblDvGIIJQX+fO65OuViLeDIuNtCwpbQcu7Kukx20OU/
t1q9vmeJlkbg/vS+34oqMLlmNHWLbk459lgesMRRIiFdyg2iAbkQxpjoSP32bYwj
2euNjnyXros223p5oHRr1did1pYAh5VLrMYHyQQOcGEt6MzVHAJAoSd+atC3jBQj
fmIqcF23CDPIHyb3vHgzrS8qKVpbOSgfwokW4zEU7sXpNlgtNM5p8Vlk3Plne01u
AkDPhxMQB3BGzJAsj/z2rhB70H6PRayefW+KalD3oOB3+M9XZJOrwrBvKSAZ4fxa
Bw4OWiJtvOULSf6ZAzivsa8rH0Gt8gPGIa6e9h922TrTYoSdFN10WJ6RE/BqAxRe
Nfz6P9c7ayy8K9KGAs9JzPhWAsMRYe3UsRDexHKYvuzu31kZOJJgXFnEEZJSUpOG
nj182omTDrr1fCZfCsZE2LMzAuVEwZK25sd0ZOEnd1flXy4RrG6FAlkymTUw7Zw1
WSumNIcdsJIc7T6m0DXIOUBw8af4j7AhDyiPaoAslAQxO1d2NtZfzqNtlYNJvrpO
BTzZgkOYej2XEzPV4iF3LSQoAnEdTrMptBPovV/CxPEynUV7xBCqB4N3B5dtewDT
xx5VPbg0z6GVkEycm2zag426UMPbn0pfdUxGnmOzZKNHfGqqwZjv86Oak8vz+9tN
HVKKMJGfeU0B/nGk64DX7ckUavX/tKGpKcN9iVCOTLYtOg1bUUJ3RqkVvbSk93gS
wyNfU7xszJve6AaXbFzcceSQT0b96zv48bQ20o9PM1k+M5Q+A6KgpEf56bpAq9Fx
uU0/9X6INluAKHpCRwbP0COUW1DDVbJH2MMWl+wJR6kUqyNd6CQ5sVVD5zdn4y+F
I9HOQZoSi5CtUyu1qIZrDHyILzSbpebb6ipfJNPqk+iUiE55KEGkCIGg3+n17Q9z
Yy4miPV16sgJ23EFsWqf8NwblK13gEcgPeekrOXBdalw/dAvcZFXnmlu3+2ft9CI
3AD8x7WJl4BKWSP9lAKJdFX282EbIgnbXe6ZwyDn7bHX0LqiPIpYQmStl35FCjIq
xcuv0BKJE2v9GaKzSZmgoLAEzIXtZauShQALm5Fwl03GFQJzSCkHKi9d3AmwwWhN
7cqqt/YkVxRUqgSXZYaV73xxtlWy2YjpjUFHQudCb2gtPT2IVC95ZbzRxjQHh61J
HuFu/HVpTaMX3rvF7vkAMoDTu2NL1ymxkwi2Rqk5Vxtv2QyxS8GhDNGpadD0fVAU
O+39RJLoGEQ4OK7KudssokYSrAFTqGctVjUi5BR8rEDydVbOluA3ffAO+Mvvf0yQ
bhWPRCqHpWwdRZveYMSvgG0ifPPfEb59UmUHeEH5dgYO2yuCPbh4CWhpnVdxn82Q
ITdaHeTyar7oeKODbKFEYhnSm6WUPHcgn+b5PeycrUb8Iybyd3BQqT3V4J3e/chH
2BcyppOkib7pIVhY7HGPgCkVwUcGvwdjMYHJfqe12uS9/ULYr0gNU28O86EuD7R+
GoKDH7lJ2RjgPbm6qaHmpdIAEFxz9rAF9vZEuU8D6lKhJdzVGZMM/UovwuckNnP/
DfxYBkvDoKLBVz8lBla4n0AatIUPmwOMwAKKkp2JjX+sln5JlLY8jybIL16oYPtt
W0JeNMrT/BMw2WNhixajnK6NGqffY2oNt38Wi0rywFNiNRTD9ya9J2udYzUw4cFQ
fTTuPE1YhESHCBU6kBx9eXLhOclIgsetaoXzc1n9nyQHX0ekG1y0yIyV06rZvS6Y
+qd1yfXfPDK8uODnvTin8Ca7YN8V9g0eDCjvE06YsvHx5fp91OZOEqO9ap/XC/VF
60am2bccb3ZnhqHuGf35sBL5E7bKQk/PDFd8BWuaDevUejk6hyL0ZuZpKQ5knZqd
S8/PyJresKAOZPafNI8n+m4Zo/fcToh56F88zyUc2OfpJVb30M/Nfexla2o//A47
b3W0giFMnli7uTblwx0eUu9YpRTJTyPQ6Zv/TnaKQrWCuwcnLWzZ5KG/VHHE953x
AHZCfkZre3oBgl49fX670YzlACzu/jFrnidwS4OYDDoErC6o5CA+klUCTWXkvSn2
Wwexpd1BFu5vIlJWI5kxFlL9fHnNVcqUJ1e3fU8NkxbZhnIpnO/IlMsMF1eijR/l
L18l+K0Wniw4VQ2y1DLCe2WlH0p2+IC6/2SiRWIUNYZ6rJvLaAlyxxsrzWgbIklN
K4BrTOblRYj2Gnja0NWKeO0kbHUc5vXM/eE3pDYN6GX2d1/rOs+FbN2abtFDycKx
mX9t+tMdmZCPcMlDHE5mhAFS0yxb7FcPKCcRPuBkpJ/pzGUOhS6BTka58zQBg6Fp
uPP+8Fhs2M9Rv8VYGL7YtPb40e1ddvAFG0I/BkmpKHsqwHVCrr+omP7boJHOpVa7
4tkNIdr7V/9rHeCHKLRc8mfs/MmfHIr0/3KbfdgHYjBqsGL/J4yXZ7H4rfHVj6th
+7xXDHs1mLSrrHahiizYgaE0fEPcfp1vh+2WbsHUGUueEjWh93jUzUPbCz7Vpjji
vvjos2ZTZH07OaF13vv40By1AkmLLvcgwKjEKyvk8EsbFX18ImTEzl4yG3NTQn4j
kB0LT9BMZCgcIDzJzAYO2XDV/tu9DQXYzLuixVlW7FwMxs1CmfjjEunHBmNa1k5S
fDyX/+9z+27Tvo3SX9ArkkssfQAzSr9B/t5ToGks4T+/h52aqSn0ROwP5jE8VDi5
vivOefMtVY0PGejY1Bq48bUSNAH0wpStIDiKAfR2YPTB/8hXCneHm15lB0RUZ3ob
MfUL1w2u5LB7T+bys/F5re6+bd69twG+KeIHuSvNro1Ig7vc9tsO4RV/Pk6zf2ry
6SuHP7GI7q7vRtqDTZYDZOUcE4t/W7ImgwOeGfLy23+32YQ7h+bIqGrtfOlTnbtA
7VYX1zyT49rqmiB9JhLDeSGJcELu70g9Ls0YxzkH4H4LiNR9RyQbhXLX0P/MrtvF
XAGZs5ELy1EURBQuXGuncNkcuZqtLiL5N0ogNkQyC9D6ImF6ttGzMmcbeyAbprmW
hE15iW9EiggDEvqZwPZb8pFXwow2EFiFQNjSazdbAlI5tZl44fnN9DUZOFRH8UN5
mFwRPZU6rIpJcmYRESxCK9cSkEaWC8c19/bdaEFVsnDQRBn6vHwHr+DfO4f9ARsM
FztmTYmIBR5Gbth4BrjxFjwRjlsNLQdcLR/GQBxwinUFY0hz5g9Ei20QfBB0/2y4
TG5uZSI1xiqWinpfRiOZmU247xQdm8Ti2+gltUuCAoNnTLeNIjgZUcQGAVXchNDC
FES4A9dGrWqnFOXnfMpX4R2onAhqSTAEPo+IXx4eQ1yTMrSfOYJrXKO76kfnhxR6
eUKpUdnX/sl7E0xm3sIs9z07wz5HCfD9HeM6XRAQo/IgnJUQiE19Wz1QWfJDOEeZ
sK289Zzxobi1ic4L/iBKTBlTEn/ZhNFodn+fC/LkWXclzuWlMl1ZiRUKLuJ+guAw
ITyJM3Ygm8FFHOwHbiZsJXbwvMKbX2TyTsaYjUNsV3rN43oUh2X0NZnQvf6r91HG
CG3MM6kBQhS0BCHWK8DdvdizhLYpcOvlGkyqVasqQjTzBhBvALW2khB5P4MoLkQ8
up6G2Yxw3TGfZrtfsthpEorwxqyfvEgBqh+yR1p9M0nGnMJxlfIfcgDAUOOw0+uT
TntYBEMYEtmjakO5J32MLBJBJB+Sx5T/eAHpBH0PqAytVsejHT+pbi27eQNtfkCw
xKrqroViDZ+qM4ZTfN0+o8dzG+17yU9SY9aSlUULxfcxE2bKc6Mw6obeRT0PJ3a3
nMcu7a33kf4o3zjo/sD40IQ9OETFBp5IcCLAXiVAfQqEIuy90SX257D0wk5Vhrdx
bvDnPqu2ha48G2/6GzDDyWanyCHUdTFeSqjz6b0Z7kkcD8wGdNa1bIoCJCzrHIwv
oBlqTvPWozNX79oYrAt+ISClhbhxwGlrEENBjAOPM6OzbxxUi7O5ZXfa7OKfx4bw
Dctg5NTtNOrIGBw2KDjOwln1h7euYHFUM7ETfkEkyYws0ND2RHuTe7BejwHETY2k
pkZ3LW/ZGxSMQVIQ+Om/gkW72lKuL2UBAlLVo03bG9DnTD92e/m77uvPFXF2R1/F
eDhNlL2o1tGLH7pTQ5xlHwaqYFYmv19vZjroKftqs3tUbyLkcLh1nFWLx3VrgdqH
O4bfs/A/F1mUY9vpg3HTor+dEd9u4Pg9eeI3Cb8lmrSghtWBJNvikrmDuQ2edWGA
hHjpf/HLrzwrwfU/JQIhD2gtflI7y3QtV3DbzR054UIxk/y/j389mlPbDv50bwFJ
iQMrfXss24fwtWLRUVbeCGdPX7x2TBxAAB/mlb1yfZ5kKuLihjY/C0ZhKevNvNfb
osl0N8R9vGeXWt5+cBmvMBEFCDMJRMU2tG+pjrZAq+WfJBtlsFI2Vmc6ZL5P8v0N
kpD9ofO/vUmkD1q6YOg0dfPiA+CE12GLA5/ThpBCPkPT+5MkFkrL2I2khRFLFV2T
iysCB13kv8iHdnL0qEo+nAF9lfBn1+RFMUHR/a1b9TLlJvUi7IwklK2v0vgkGYT2
CnvNYHSVukeJuSoJTxkFWp1R3JFS5qxKzSvC4SYEqM/mbLuUnul/gmwyHNky0B3W
vnSjoadyqd7AdkxmfIdfoU/DkfdzmPpUsMpsgnU240t491aMtLTjxcEHJCbBIxkc
1JmrcZkUtdWqw6+OV1FrgRDeTO6z1FblbeKCq5+EJjGJq6LWP6uKbrCduNtwlZh8
4Y4NwnWx2+fhCO/ySMebFG/yTHyUkyxvAXjT24M6Dn3MZawVqi5Roxwk036UkinX
SOZEKjxq6VHnojax8YNx1hUUAgKRt+rMSkIhf+VwTtP3o4L8ghikWhLjv1GwJJzB
4bAa3NidCvUM2SDJy+diOfY8DuQk/m726GrtcPEDK4AWiH24tBBeNCl2SSSLV5pn
IGuiW4fFzM87k/6pO3H4v+37HZruO3bpu38Ki8Y9u7N45/XERzv8bHnKBHrdZpP9
NMMPeu5bCYbHmo32z3GSsjn6BvmIfIM9xQ3AB+NgNqDA4KsUV9MhN6CDMj26S5n6
zN0zW90p2FZxQHJZ4oJSbZoWmBZ4lwGcbUfdcx/5gdluNkrVDP3AxDfXGKtqTMQY
gO/gMIevWAUKuCQnteKAtilT43al5/0hj7x7VWmBEb9MIfP6PZU/nsQPGC8WKpoI
axhujNK6qp1Zk7tN6wtGiBJP5QQCJro+dsNKKr5VQLyK0ag6AnRopYYuWpnF8Epv
wi7Z84IOiHeIkuZB8cYVLXoxGGjWvU32rTpLk5UAK8DeJb4tEcnFqTKOmpXjIy/A
rE//lVpmoRHXVWvHoHM7ikBgw633sG7IhNP5lgPDA23HPzvZBnEmjhjUatS6Mavh
247szgpl9JEV6oY2vTLm6M+YnziU8IMdghzKkajpMkAC6UwBMUAjI5BJHsf7OHqp
hs/A3aR7tl1yoemGUqO+/kr5G1hxhuetxZ0ebPCa6aHfOsxE1tegFGkEnq/Ajnyx
SxGS0ddIi1au6hqmVjY4UpfllfHaoM0+heqKzmhjnK39qYpeN/J2roObWlPhztHd
C2+hZYKQZMmLNGYYw/5/+bw5EM1x20e2oIum0gwPeDKnuV4zH2TiZ/cOR5FgG7yr
Gn1PxR00vh3e0M/E4bZZza2sqVX/PMSh0JPeyieJd6Zg2EB12fwWtJvfeaGi5zte
k7tl3hPPPOaVkW+kez9hSKQOZZGIPuXpKF+XrNmFYoy4l1ztoB32Dz2xYhyKBSPz
RBHzCDxs2Av/QUwqfmIvjU4hojeOeH/KqZgcWbcppm7Ry9fmZEk/el3NQ+uKKsQn
JbFD+d059xpkNPmUGqnwjx55BmPOBTJ97+8o1uHTSikQhS38YWIVhGxG6qjScU5O
EqhgQhC+eQsn1QjDYvodW/d8bPu1Wc+iXvpt8E7iY8X0YJvwfAiuWDDP48s3LYFn
F4hgVf2uMMh3hIOdRrOQIILwqxWk+9frKN0yUe5IZkA4xiehtZjyqLfXZaSyqlnQ
a1qC+4vcW8NPov785c8ViPIE5dBGM6UoJd7hhGRzyvdWUUfRcejCvHLS7FP9gUK+
j8FTcax8ZzwYmnqXqyRKhdUmuQje0v4H389SaL5AqYd0zhZVzYLf292IqrI2cXVo
b1hC8BBE8JMLbbQV1yvI/5h4iR24QWvOUVyHfD6t5G4Z+v+Wj/c+zhdlctb6oq9F
hq8XdQzPJhkXTLK0/igFb58By97aH2LrzhZDEm3SlLMSbg+y4WXShgDqvyNNeL48
gevzyQ/KsXJuR7cjGCt08mW6woliDfoF038nv2+NcgktuFYbvz4RvSwvJdrV9qy7
zCcSfa4/hzRgVuzgO8Zh1m7sTDH90qs/0p6OLXW3b0XUud5SsKAxcDxN6OZIoJXa
7hg1P5a4zhr6P6jE8EdmBkEB2EQbNbILoWr3BOylPIKh+vcRxZhSFwSIRmm526Q4
52SJWXwvMm64aMLCmkEJX7kcXK1F4LNa9xj2BE+sksiG5UYf0QH2+Onb1cGEP7JZ
bQxayp8fa7KojbHk3pPsaS/HilCdRDmJhcVAqMqUcR+030lbdF9+UL2IVvDoVCAE
IvWJSID4jLJsanQSFbB0N+8wpEqkGQloHeU+/a2+dxgfb1GphCpxHvItxA7H8dtV
mQGMpBjwBFT3mnejIgabWuGUqVkNCvpwhMBLOQaH4lEFIcz+9t6Q+TMNPswGP4K4
ToNVYgA+Z9I83WfPN9rLq0XadXScwO8O5djPtm/1Kcg2mRTz0KY1ARRXbk5xtx8Q
YYkxQAvo1EQME/UARZ1gqq67GGSO4+FpIuFKeUiFNH1QRfHHEuZ9Z+DKSwwhAtIL
d49enPjk0HlkXrJcUML852dwJMZAPHaRIkeQLm7ipguetfkhplzzEuw8f2aZEZwG
ln9zOtSwIPNbIQuOM3dgtcIrA0nJhhQunQTflY7uPM5Ndh8EApEPDLiPbmTTjEG5
juYdRcDOwl6yvXyWb2J+HkCNb1t0o7pE2CruxdQXv6k6ca67tfETGXKxkXHTAVII
O2AGJEXMgarY62NWuu6PYhjnU50VbzGZGsR8FDvrI+TSwd8iw5Fkc4A8lGaxrFol
y6LEUq6SUgtBfKtvbHhYjDhEqMHJ8T/tH14mAzYOHvffqVAkXREJy9munVI6oMqK
dVJ/EOKNJ0F36kDWCPj3zxFxvEFihPvJk2s0gDJC1fp9zSg+t2sQoqDPoNx7xxSQ
1ZCG7Y8t2xZHGqkQ6DQdvY5uKTfMiIyM0CBKdnOG/VMB7lriU21Lszvczo6gSCAK
3YKUVEQCR8OdUr5EpWWopjJ4sRo8fDmYE8k0B9xatXlwVs5rSiqjSJ0w6o45MIBX
3Q+sLUgZRFSv26KtCrZSoBHLnifSIrj4rGK0p0uJX5rDOccWkWVTVLrwm2Ed92D7
OcyBpGsuqjnhg0uGtSyEE5kUihdMshKtvzoT7DdYRPosbWIKyww0ig5c2bqdXRSx
efmyzYRCkm413Whe7ThHUBS4fajotHQzPGFrA1R+GwDeJIk15ttVWTpu0dMwlSzW
aWn30ab5CgPyQ573ile4KZ4KLhjigN1RbcnpwgPWRyxu48+2KAXj8eWQUYryoszc
oMeMOYt9MCUr4RP6BVexSYwWFmlNaMBcV6ZfIlOlnI5SRXWNtvFCHVRI3MTuDtWP
+r8vlPFEAj1sALfNOZj+SBbjY3jUHqI6H6vdzYzdxiOWpGWQxoZxeD/6aaDRP4SM
CgAWv737+cCUPowXBUnIgHSHLSuj7zp7bn//fu4rsAA1YzWrychQFHN/oFdrI3eq
D6AstAtdz6s0CaqnADJZP5rsYzoftDIkuq4wYLzHi39W4oyFM7x/NNZA7rRLdFZ9
2+bznr4vS/TL3Tl0XvH7/0Mi2RNCtMlT9JTSucvcT+5Gg2WMHK3LYxY2Mn/EVV1P
1+EzO+PbSBHFm9MhRTq3zoa6qHyhqXRuIS0LJuYZDdCZytvWpvg0Qlq2bhmti//1
ip1qtgHPyleWc7dQX9yJavAoSCPXk1Isoo8sR6u0mMG9e5FhVGvfF6qLDWMYlp+a
ibUj+p2pxc81Of9PWqdnOcrAaQFR0ME4YrBEGGwXPbPxpZWYhcnrC6R1xUTnhZak
0qZ7e2HGbRCtsWDGWf2v6QOOC3AeMQy6rrkITXloyByz5OrPTl+AuFhgUZElZ/va
iS6IyYV9fh9EvhTYhNxlV4g1D2H91cKfI5UPNANH3ZeX3t0PYvwDUoV0PuBJmsYb
Mv3qZMWCr9A7c6k8/9NY3WBPU/8gDG0NsiKkoiwDCM/SubrwQtS6WSUCE0HbZa8b
myE0P3a1hE6/2cp0CnszlEDH6BEGQDDiRBCvCL8QndOmt0jkldCCfZxdSfW5LCBy
ptUGF9EQnl0s5seIwzaZeFO9H/0jMo8nKYBplwrQVj8VwSEbod/fwsDSEyduIijm
/9J5toWpdr7YCnTrT7obyUwSHpdYrvKSYZ15pkwneZuJxqaWE+VijsFU+KRbcWVI
vvAnljZjWXZsFj0ms0K4hVmkPLjkIYfmWFzulxAXdmJzAYiK3W0SQA7enYgy3mj4
4rlFOKngOUlE0D4WS8E4G1H4HAOWW76EB5K7DtMgjfTOe4ZFevwHkJjTk9W01gei
DHSIK9tj3d2Szj8w9PnvYJwxPmeMOm2MFrpU8CRnKYMba6SAkxn1NkQtyCXEb+sN
cjkcP6F5JLMIFw7aS6l64R6PsvBK9A5UGz3aQ62ccirQtIAuIwhlWxxUXuyT8AXe
IkfevZojel8SuOCIsRLtQyUN78rrLS70IolFcaJxbEUIQtT47gU6VAwAjI84RZ+m
xXcbv9uOdNmafzMNrZ6GQAhxXjZZpMyNVEzemHRFHUqf5KUzsN8t+yMqUVqhZlF3
Q39gLuSx9g0BiZi1A85Q7c7MAB0VpM4/B+1cmJH3Gk1FRhSVbmjCW1ucihHSkhNu
RfheWOGTidLXIlJy6QzsHn0yQs7B0GIlMAoGSLvXOrsn2/GTBpUaIRYermH/HnTZ
BInUGDpBZA/JQNUNkJRshzcJ33zJfBjj/1seMSuj2ncHXkVF9+JznMZ4aFJuNOFo
W0YmsvHi742wmoOnviWFCakVExp8rgJ8+4JyG22re5UDPKao9t1pBcywRUwxjGX9
XL3FWlWCC8EXQi9iApTIZkQhFtaPcthUC2Oj08lI5PIH4AoCDTiyHfED/6yZM6Uv
G23DAmoVZcQD9Z7SF+xso44nRPO/9EuhUGZfR49l9hY/LhbF2BN/1BBgvYlg8Vou
b6ppOGD3ZeaSgdd4iKmKgEYFYmfe8XCE0Jzbk7lOUZsc3P+p7P4bRXByaOU3q9wH
mAiPPsr/8zLzyHNPZjSPjS4eP2qCNJ2jYYG9RPU5+obYvMLqFTP5z9XUyqaIaXZ4
UT4NA3yXHoASELdyASIMup9MDNudIN3kcO122F06516efpPn1IdBhv0bK+x5+Kql
DG0kAubQIxJyYPXCU42fXWUTaMLR3OQvVckFR5wQi/F1pc0WWQlngZlAlX1F5zn/
LeWy+BzSOGkaZJ4FzmvxRGjwX/pO+3xUcd2UrW4Mb1vc9oFun72zbvReWPUVclam
UO4jWHw5ea0n+1MhTWyvXXbcwR4DIjSNKjaG9rihYTTf9Ird1drqHXyA1gfvfAyi
VpI8uT0l/5EUAfeSs4leZkd8Zb95Hm6JFkTt1pjUs0QMu7/ZDu7DorMrcwddhSR7
er8Wh8Dg9dhiSF1kGWnDd2QE/9L63MzpT5VFUEyC9Bby/eZIpQp3xqtqJlAJkuA+
7AikMlWdQfoxQhCu7Lvbp9W2TsAy+FKSI5Y+f7EDM2iB9kWncMGGiwjaL1QciDhB
hVIBS3LpvYn3+hT8hKqpUME9bgMB/QeaH2B0MRHAmVN2vWNEfOz1x4WK0S+kgWgB
CfLUZyXcjKnGUMWx0aAZiWnN3ieGy2hFht+yPycflB3ZwOp37IdHaht1wRnuefVw
0Jre8ZiqlYnMn/wl+keXyEdp7f5WdwpNpV6iOVjLZ16uxecbc2jjNnnm8IwOXBu7
sje98YOnOEuZptdSOGq54QGkV+T+qVhZrhYyacrfnSU0OZTCw74eiebyWtuaEcRI
nLojSAU+KD68MdFkpamiyJkaBuNVlKiyLKAY5qRMnMse7h6T4CuBEwRbrm8dL5+R
NSemrqRzk6/4/m+KsTX3o0qDHJzmO8+xNOna3lhzSMCZZIwfb3H682/dDIawYk5D
e5Rl6yKArpaLZKnqSQMtaLMdFVNijnXjHfSRH0BfX3QASR1XRsLiceGQyFKyxINn
z5jDlCsM0efDgycuzK4W/EVHWI8IziCwgQ+HRj24L0SGYm0omnHcghZVwoM8XHtr
Y6C7D3qDHchctsoQis7ZSIkthJg1/3P8aN1c0HgxFM6x/QvvqfUDhzpUCUPwFCyo
g6pKXV4xas7nMBPTh1eU1+3hXB8ck2ofh79w4nR9fjJ7bpPs8pHBgfc/wHjt0LFo
GR3yzZv7JsOVJ2O+LEMKaCZlsqJ5YmGvPMgOvnqDDVzkHvHOo1R+mNNBLzr0NGW9
vp2IE7cZtJ7IjbwZjW4WIDZ0hHm8SN5rXFU+eNV8k6tWaHBG84U+nEHGRNujhB/Q
mZqVaSjS65ahAygx0sZkHJ/ktPkhPEqLakwoOm2TH5eNn8vukITXjP//jWIbktQV
iHZEspr0s56Iv/8P69AUGyJBwVZ03DiG7dwTKF1SOlMC6RGz6sGRDCJmQIwcpMqq
n47rt/PCjCjNG3LRMGd34B0LmCMOAnVfRttRgbAdTMrK5jNc21PCMCSKVnIvsUIt
KzooZgLw5HDkc18qyLln4OkhigRiMAQkromA5jhtoCq/z7/aSU6kSNFRxvz9YKwF
cln9VTqWaJtwfUCYcs27RR8YrPU3/42LXqrk/0j6uiN33TJ31L2QXFdnKG1uPj/j
98jPhrOMgfe0e8VVXQfDtbSVSZ3HEl5qSYKcXcBbz5R0Ys0mDrkkqDJCkJOMw7uu
3EuuFxXvRwmYw6V+dNLzCgSiaQY/Dpn5W9L779yFf6eWtcT2WW60e80ulV3KBwK+
Jr28lbLaSbjpzhxBdWJwxlakKulCiTk1bWKc493ok+vlRlGkFa5T8k9kTGAyLtOU
iAlBUuWnw02FK6CP28gsROg4ScviDiX/9XbPGyjGx7xNjBZ+N+LJjbczzD4w+F9h
bSYfJGPYxdPMWb8bCqi1hBLjqOBeSDfZzbD0vrkoF+FNUvRULZU7ope6lI9ft37C
xLP2rvFsHyb9Ek/g4C0PVxnQt/OFt4i6M3p7Te/oLvTwpQMIvdUvm2VFpWP94ZqT
k27F/D8mg68ehz3jKNdy3MBQAGiCUzBBRIOMg6VK+RJtbnQZfqR0AVeAGOYO+2Br
gEzcKCAvGDRnc6bF9esYxjjDR6MWdAc8QbqwCUXIxAnnwklrcCQgcUx9sTMYCOJ9
3x/ZCICgJRuSk6JOKqZ1F51Xs0GDc4hlE49jliqorRtU0tt1NoONVf1rwUn9BJlE
twe++SKtdo8dsGeIonlM4YDjtUVlxRgd+L7knqKG2bTlYRYqbkjocVVY97rZYUFn
7IAnqiMIOv5EN7KxzxOk4rDNTL9cG75XTKPGP2oVeh8o2ilA06LgKHXsB+ZGlAof
hdcpMs7QygtmO60fnq005MJGOaUkE0UK9qg8BH4ASrQa7s1Zpxg8/kYfLDaAI7zc
4Gsh3jPGWmKqXRhuN0hFcbo5FblD2LVPmYEiUuy8wbup+0qC7g605jMgtU51isPZ
0VfTmAdR7gndaYfrWTtcRj2VDNIHoW4VUFRFot7UU1NqUgDSwurVJg9qhery5rDw
cR+VWK6W15LqM2cKthgTuktxd6h17Nqmwik137qBm2zStyK/WdRu/0JLHinI4pmj
2w6N8D6Q8Uqar13/hR3Un/jqXBcp/qUzh2Mfuk2X3Xc5XXmQfhbEAXCoW9JDBfwe
Nh59NKMNCrGuqib1RyhEKGTV8XZucxD7ndOY909eyvO/EguK5CRTMUomx8TB5zNI
TzQFN3ygo7ReS/cAEA/YRwjsU7lvcQmTlxJrBAkP/8BjZk6hDa2Zuzns77AIW8KC
V8jNreMfjXcG9ooPMDANgMemSVuVVgCfXlsoN6Rv3eVygjMR22Hvho1fQm0HICyw
SE5OWNyNyOvZJKNcX1P2IxI9RdCQH7nMmByfqGejwubnDYzGFK6BQjy25asDGFiu
QHABzpugs6PQXZerA3pHUequ9I6MJnaB00EGZfvtxokyPSpv421tUYAGE7Wx3kRi
NSfdI2ZkNLKFQb2cQGKclWI2sNDyZLMJJE1tyr11SVbFlnI6P2wRduiO2+Jc7G2o
JXHBHrKPT/Jip+H5gaujDk4Rg1KUsPnqDSo5w06Cs8DHxeBkGEQmuVUobfrKdyXT
uNPkzyULBNCFhAGOAK004aX+5pZ50V3mOsv5zl3rGFHApBMUr8W3NN/fLqs2RvbU
Stqamfh4T++iKb+pk0AJv0kYu5IHHuewZFxAP4X73+28TALzdaxJ/NpX6ZQ889hn
kkFukOxOeLowgQmkzm+gM5xkel2QAsmlymfWoRoDlxBvPOBFg9Ru6f4GVNkhzYye
7q/IOO+ZgI3h+Zgb480nAE0h0IqLUeem6TpLTP2slVjHM0bbZerYVGpO/7Oe5tm7
H/fYVEZwS37WTT6jlNiq0VLqJnVgW5iiENOnX8Kaltr0SIG/OI2MoBw0spGo0fWX
pms2kpELVd/WQC9e9hTGgVf9Xx+VnSB5LJWylB1/MQ+gPoItwXPC9tmaMO+hB6x+
HwibIffaLiF2XksAA3pkuksi3OVdhkPoVgVWMoz7h2dBjAppqP85TOu8aDr3DQb1
E68JRWPkZkDbaGn3vQmrawtIHOpNVrl0CMSoq18tjLMIIStkgAGygw7HiPH/EK9q
VtbvnvV9Oj1trnNQDGCRqBDUoWV4/R042m6l8Xk3Suwb7Vi97jyWLBRYjL8m2tsn
azGRV+n+yEt4lnSQQe8R8zMD6EsLoR4PRgApksCdffHP/MMQhMWj7bNtcpZ7ioFL
++SnjkGTpI75J1F6hHZZrD8s5BW3LCP8uSK4BOmoN4017cjX3Ld2oREltQ7wfSf2
T45hoJsEDbnwAPtU48fA2JHUFD2GSMVZvIPuZHaRGG8JrbDq6ngSqO85Ip1+LaRd
cx9XR93bRwgyHiJztiQ65shUB2Gwb+R1Rj6Gg4PCvXK19Uq/he0sX1d+wISP8/cm
XoEG4oXSvmbEZZ3pw62PHZmmL+AMZDGiXIhoGHL0tY85F3t+mw8Qku4jW6EzsoZy
/5AmJ+yVYTbEhiXF4xmIQCJJns2ynv0Tx/oimhbGinAmESFJGGnsK5GjzwiD468j
dHlBgAdF/BldU19YlQ8KGxa7DzYyQt5vbv0SG6Cmc7wgR+YFLeAMqeHDCtZkzWzb
+8FC0VXysgQz9lIOSMNmC95CNFMvqz1cJ9owzliKtcij8jOqPz8Mul10DmmXDML+
N7O74a377V5Tha+8MYT2aPeEJZ8qQ4DFezS7hW9J6WdrPqhHn5e5Wdxta17qk6D5
ui8U04dtjnb+eviKWu8uKK/ki453KBeMZs44srO1Tm3D7e0wgljBRqojbVDqgjEE
RN0L+OnSLFAuvYRETV4M/Dfj9jDeXRhZw0mlmH6yG3e7ebpzM+0QjXHUwYk+U17E
wtbjPij3VXjxXtAp1dxx5ASpb8Nzp8dX1Thwq2WMBBT451AKLyvOt/tbqC7S8N7c
MaxnhdbPo8yld3Il9g/1u1cPsqbNEOewJCX38csrL8ZYcxn7nZkqFjLcVCZbCqJo
21N9oiWXpERGmbGDSa5scTc9mYT+HrBi8fvXE6dwkIEe+Pzbs0m9B84lDbYk9uBv
VJuQITOmlVKAjHKd2KD5zERbv3uOL9jtTg2lpWa1wupmKgP3qL5GXrZjm3kuyn2+
QCrc+GGdu/+G3J6hRtt/Q4yISLLU3wsXZjoK5GGDiNy8sj9kposzaTDks7TTTckU
a4q+gofMu6+n3JN63hSH9jx6vlzbFhhlXDwnq68EY0ei+VMSMOeJEhUa0XFms26h
qlynadEWRZJhojzb/g8mgPFt2Pb1RmHeXOyaQ7XaRNYAhJw+fudO3Un6+A8DSPi9
Kg70DuVQhCbGQCV642VGAfkMZxNMM/5MYnUSxXctHEC7AC/2HwAUpoHqVOeKozh2
oIuHvhYUmeSYi5czDfc5BHUwZVyxIGiMxlnB39WFEFr5KKFvdM43Ls3524G6b3S0
XvU+//EA/3xcc0OyqSEElBGDJ9n+cZBOztmiULwq1Mwvt1bfMJJ8N0Lkz14kBoeH
kBTaHi0fs1qMLOJevdGGUVZAWv7EWoRUAQMIHpZt5BbycRNAwEzvFsUwlNmRsXPA
bhSS+sHtFipFwg5O+VLJB9ABOjUFKf2rl60guT+pEVimT3ZvfYXyFgolQyB8bUb+
iXOm3r6djkMlVaJliUqNTN1N2mZI5klGhOB6EM9k7HlDkFL4686w1QGh+AlorVcw
Z1ja8yiFT0t0HVIxtVmZMXKIgQxjm0Qm+sQpibdemRRXwBzlNjcj5tRjmL3izX/d
Gpdl4d5e3J4kaOJbZ0VXlBwjPhqER9pm1JcXFj1/QsliYcujJlTodkKxCNcYw/F7
cMcV9hH5YQRDCWXF971pkYPLedWX+Nc7MCE3V7YzZs6gs+iPc+Bfu3Dljqcv8J9T
Ey/kJW3kszAnyv4IVY6HSCSIn/IEOShw2404X7gpnfmvHWYEgNSTUZW2Aka/O3Cy
F+MT9lPt+k87OUyo1yoMpJmkdxw7YIL+wH6TbkC+1pjTwGg3DZ1Q+p/VtKA2v6+F
jahnpGW3T8JF86jeml02DF1BHTIjir9dC2LV6VrCKESVh+AZxN7I6YnFDf78rb1U
Jdj7gYb3rj7uj1E4U6lJ1JgxHSgC/BIoAs7evDaMIDZPX3E1rLFpQ/9LZcChwKHX
TyHb1HMLTzsLPox7KYOXXQvVP8OxfUq+nSRhIxMxl8VhtFDhDe7zqsffTlxRm/uh
vzHkhuMOgFKJUBj7pB27dQpDXNlHSTd4uxPR8BJzOCIixxsqomY5kMuECzUWJ8Cj
+ZjeDJViNqiwRtuMgu+5oBN1KFpDvKva84F7DwYTUQGRxta+y5IObztXNYCYxJpI
tsNJnLLAIT7QR/ERvdNVPWe4Mp+U/P19zvqfaxNDco4eN3AIcjL79lXPdxsak4OB
Jyhi88+Qe2kEBFcq/L7Ko/ZM8gJPAl9Ak6qqi2mrQGVTZWrOl/JmwAaOb04+DyBB
TYQpSvx3JVRjbQPxHP8XJCzRWv4baOXcQQJ5GEm/FRDSJ3EZHkZrEJ5MSVYeEGca
sNpjcwcsH0crjIv5E9iOaKtib8bClyAoWzBUJ7iM6NoSvDUNuJdPU1SCbA1r5uP6
QYciKwHDlnBbzOJyuKh8Am+vNZ/poBq3Oh6LfKPqKcu5MIw6VLmP9/jJ9gg7Uwtk
Lep2XL9w9dKZXL2prsPFDlIFHLIY/NiDcSLNague1kFmKw5GRPjDzuWFknlmFQXq
cPBIjemah8fX0s53Cd3L0uRrlaZLJQ+6g1SKC0ZyD4u3fzir4ZbLpsvR5N6SPPkD
xtjquOA5sofvwzNDyntPR2haYrGI5mzRruSO/BViJhDis49/4wGuLWdWXLKDHbPY
KQum1Rvd8EJHuexkQBF6VyES2TBbUZvh9cW4nOGOWUg0DHnVzI2EScFWTZ606xuN
UgBiHeFi1Xq//LXgQFj6rgulXs7yiTIBVDcIgJ3/ZNMq/4tpGdcGd6wg3Yjmf704
aSoyeKyedZuvWn98gVsXL1ChOBLu8ZfCNn6dKNfoj+ZbL5xGVVejnh5T+6bpXt1w
0Leu39Ktj6Bc/XRY/VKTrV7XZTd10jt8TkT2dUwJVzaZwroXsCHOxPNJbFtC+28W
jdERjU/PzRyCNlqozS+R21Md+4whNiPqpkTclKyIDsM2a0Cx8+2SVONVS1YxqczD
k9IB0nGwsol2AHx2oDjc9Bn4nCd9xnQcnuramH8iAb2lTkFrdMgiKv32RZJX1TG1
KbHBmIk620dNxH/1ca1wMyWeBobK555N6H7Ox4SiV/441fR6r0A3OHgy4VP7I58k
mk8vSHUAzmVtUEUU0D7K7zSX17fqlvapDT9qpgWcn+CrSwErcfzRu9WEkTWGITIZ
3zob4lQuBrUvN0g2rQyCoV3Akw/vNYyNZyAIsvhlKnkOZwltEM41X4uK+K4RU0Nb
LjHdyh1CBF2UuwcF/z0rLPFu1Tor7nB+SzakU7JxysSvYzE5f0SfF2Oi/aG0I88Z
lTLh5bcQfTZSrYHwo+8wryrsROr5nqWnsiFkhv8c/egt3cEZIva4G8vw3yx7IT63
dPAd0rDgykwcGIy3XpSQ6TdlqmhSo4+BjsziOr+r0TnKG3FH6TBu13yoo0fheXqJ
bwtjEtLD7OWkUhk6h9c67bjzn/1A1lKLerSwYsKd9VenzpkXv1ClIiyQ68ezEO7E
xGzyMNT2tcBQodmnawLp8htL5BIU3UUwfGkGATqWqGQ0hgv/WCHrkXBj5kLtS7hm
qVc/dUr5tXEApFpIZV+XTNmjchsCxwqZ6q3oDpfvk52CfdGOBjytSZUHPZjzgbMz
zSR9bYTspTJYevFNryDFEzd430OozmanayWfxNzAoIFq1YkdEvqjSxRX0VuybpF6
fGkgoctRFUIm/uq7FQZqAX6YMtPYWLvXfTDJCFo9yaDeKrXMcKb79jOHbOntgAIM
wDyjguyFQYzjPigKlxKlxS+fVXFAB4NEEFrTzO28T+CbfrSXq9ujHV+OUJ8VMoV0
Fq4C7918T2JZ48DWzsrcdXxerq3vAXn00bme+jjPl/G63PhO4ArrqPM05osfq1nu
/tk/Evrjo/cVIUG7sQ+KbX2Lnpb4Ps4GGV6hz6e45wHe4HVZRdLycAfL1PnOnvq2
zLX8PyzMocTJv+/7vsKOnl5n7Dx4AZwt2+97JbcsyvSZIwfvogCWJGQVWAC2AQNC
grfXLplaVLvu2hEZyV0WME1/ocDqqrb9a5XYbU5tCSc6gLHNiJ3EOrcJAFyxKzSt
Kq0b61ij6vq07GGFpL5rGaNGXf+UFF8sP3dZ/eHYycUPppySgmQ5O7tdasqObcW4
qi8EYXl/Laxx2P1RrX9vFaGhe24GBNCRFVZAw7jz46V16G7CK44hprrZgCwmYgp8
coRkSlxEcor/QaITnNIh8kH134tPFXkejBSNdNGfp/rTrA+ofXyImwyVZYi0dzIA
XL3OHLmHR3VyHJURWPm1paBwVvf+fFVMvg2SRYl9vYvGxZptpXDX62Op0nG9ua1Y
Ygl3v21j60Vt00ShKFMXGDD8NoQD6bdG4bvUoP+Et0sDnyjcNlC/IKoOhoi3I+cu
d/t0Dc4vmOx5NyHeG2jp4y82hmKdbh29tiB95kseTkF2jZ1oPY5D3bBZT4Kbj2/E
/bjIKrY9zLD3WgX73ZX22rospCXyyExJD+UraHfE/3FWortd7Bcn1cnNUj9pbqkJ
EGqG1mB0eLwVlzmZRTfG6+iBnXZex00giXui+W8vGk4Nv95dig0NgBUnbmPiMdSD
2uRgiOqnDLg1+XXDg6u9vSIGqkCloPl40v2OboFlEAEXanIHpK0rUMPcgdT59yfe
bqN5o+6kHwwAHEp/a4etYc9mDi37crEL1KRW3X35iZt3RBSSL0mmbCBHqY5j49qJ
wDnfg8EdQkDr/PdRAAvf8eyuQPRXz9UaZ4bd3bv/AKGtK7U7HqIvjS3Y5qjAv6ma
jRYOTkUlAYTFb1/Q5IJC/LPBfPSQwjkWQZmoQt8FjvpolRrrPugrI+YDk4HBIjGm
cUmFUbGVEvB2tekLcV50IPIJ9KvkN6zAy3bezJsCzEFHewnpCTrHroBEpGGE6NRO
PwH9pXv4xm6MhTTfGoDrIAkjBZszMythcst1LDG7YLn5eLvb+nB+nuYl74Am3ojU
IQvxzGTm1jNEn5LMJJzoHPZr5hPeRE/KFTP8VG2e1vTkMz9mQhqr1iXk5GST86z0
sMlj9UQxkCksmcRouAO87uqQYVFlMWIx8W45JNt28CacaBOlNzsnaDPWnEEc6dQ7
ZuaLEOQnAaCKeuFp1vvYCRHd7hliqx6UZG0T/42GAwvVwKDgRF13dbuwOqw6QnPO
12fx2/vVROcD7+ik0lnd3yW0VsLX4rCBZe45Z/tNzxtrvDI4poe3QKfleEcy09Fr
3+ZeQ6B9gpklGuDgRU5IpGCM5TZmYGZro/ugGllI8go98afTeRaRGTGMJ+TJy1wx
X2xrR+Jjlu97U89/29rfmPmNIkBeHWHC49qWEiib75g/mTJwbwTF2SH39qKdU3Kc
p0qtLIF/cQXfQtnttPyHt0JT8Kmv4cKkckYnIfIu4flwDawpTF+eDv+Zq8ab81zs
k6QUftLlrFz92XA8HOTFwFG5YfbTSwz5G2MS5U7ojcvNa0eB1cHn9hoPLCsp4BF1
h5La5tduoz5txm+3FcVLBr5lfN9w4eEjC3FoIc92x8QQIWo4CX/j70aejCnCMvFq
zsxXIjmOhTkDBgTQifknhTYmqjLdI+bXdiE/I8tCIM0skRntrochwdOm3B0N1DbV
RzuuD1NwuFOaq6rhHE1o8aD2GmNgaxospeMm3kZ7XUcXH2sK3ZcRzkpHd6Iy1bBx
/Ib5EQhEHVefE9kp0TFzpvUhzN6d2GIdHe4IamcoFCf4cG297/ocXzTVpbVrPpVc
c0QFeLXqE1/QT0Dh3yDCtgcxSzw08rszlhL+3Drp2XiUDz/m/5RDVtzIkhh2dtge
EtcLT1n5pKpkt22pDfleU9Khw3jYuWFN5cbGJlDBHjcwSACOhLkaqwjNIhP0Ev7v
Thn4RTp41w+KO7QSUr6nZNRrHfkhT1zdjOWEYB6HzkYw55gX7fJZjh/M/zxnzn6V
dyyQoGnUZ60f9YoQ+AwHCiVvQSytHKILiqZOhX3MV96s4skF2L0r33Os09zcx+BI
voz7FsMudaeFCOhP9+SuanSO09cZJwdZIiHu4Bm5PlYwE+xWWydF1x/w2KSJQ0HA
g7MGniIhsTfEqcL4BDOIYt87K2TWrMqp0XUByrnqk0xemuv+mUZdWthPNj4yQej4
d9Bylx9iK16HqK7gwFPeqUzPXPmhrlbkuTYxvCly5qXxmV/WEOkH87y6hFmF1JjI
qmIDObKy5l7+NrM35uhKoDu+lgpBsDz7IzRWN+NBYtp1uNklw2i4L+kb94BFndxm
OYcHCC4oRtorrRNDyg4BhUA07mE9ByGuemIntpUSIwYyFDeFF3cbc3fFMw5eEWsN
uyYle9GUvf2IV8JV12BVPpHFFLr9wnOE3aOw45BjAxnvdKSlEK2r52OQhjI9XNgz
aOOWzm7Eu3IWgjK7CkW4nKug+LN+yj69g1glYlEX+I765tHgaPciudJQ3FskHc+5
W7LxX/zWIzrhc9D40wecM8KG1C7a8Sy7NkCBYYh4ng8zJ6+vTIS/86Dcya9Mg7Na
y/QGoK8Z3KH1XuFPbldcAhJN77Ovd7+B3xmmmTpNAZWByoVwF8bdVzAc0uOJEcrQ
2RVADQx2r5Rb5lWWr/uzbmmxDHukyltL0GFuwH/fXsEyu738IwXpOjdtFxpfE4zt
ElyHJevRpAufgSKNquIWKRLO86Tc1YGc7ZKbQfUSmOL2d6CbqEs7I4M2iHgR05MY
RIpxynIGvuEnLA5RZLM9eyDo8AAJj7NnFizEcVD7piFnzcrGUhlLjENkdHuBPna/
Yl01sxsHypou+vjQDp8h03cPUck7/H4MLYZCzVXaWuCTovRkcSIRp+LUKIja4j7O
8Qo3uHYLd+AiaDTMn4hbh/aO1sI+NBIjelCOvUyK4JocQCM2KcoxgV7oIQW6PuN3
eokJwJ43ePK4AkVTqfbo6ibylrTyA/RnzAtkarDrrPrAMH2GHEEL0t7REsTurpt2
XeUiQsVgmG+Tdn7eDh1kyDzgptsypriAo6JU4gmsiQRtzldX5Z2nqZHg2HdEj8cL
hFP0kwil/QzaL2PMAhk0/InpS1ldLQLXhfBgsmdpYhLqfEUZ3Ef0uFJwCIpU2vqR
ZFgk+g5zBc6cni9qbs+KAz9khCufXTVbb215fqBy4VYDkpfd/cZsJaLEBLDNOswF
Ijsk/kATSLtlA5/Xn8aubK6DEhWL7iYdYWOOU9fiElD3F8jNhLyDd0pmwJO5Dub3
GaofeWWCM0On/6jtoYWcvasxJ1FRbZXv9osDhCAl4XhQryRt77yMGeQxAuZxZmkg
f9vfjavMv5dfsHwwrxwLGiI4Mat4wqzBzJsQS/rRorxNm4Ru/72dntjq/1P862nj
Th+aEnTBmtT+K5sM50DrfH/HIQGhKUineZjveNYC0YCTp2tIThM3ofnSfxl7PLdV
QcoXKeHGIKSX1x2I9BMeB8HVx0SXsFvgBWfnUHZ8bDGNGNcxEthBZm1aRynllGo6
QB6BSGJyH3m5/YJ5kk+CdwqtMyQhDMmU7WeIE2Nbt5Qm9/QXe9gIHU4P/llSuGeG
BiNYTwFznronzYpxKETO/wBuP4TBbr9WqVIF3+Z/R2sO5P4hh3dg6VI6XF+q73M3
T9PW3UP5JDbsnMjsN3K4bSmAbCSDC2uCUyM+d10ynlVRl9lOGDxsJqwQGWHv7Ni0
r2vqnP+aIRE0Ui8SCvT7SV4OpQW1fEiWxZFV9RtxK1JZI9dTS89qMaxXitVWItbu
GlVmb7wz2t0J5dC8ZCdnHdCQh67jPoGYWD/I8bBfSFgP4xpyXio2o/QH7ndNtmJ3
lfE6CmCCWzD6Uk1qgxsOtq/Z6HEu1CPIBxr0DwqtcMMAG2f2KSz8QBGq58P0fS/i
J0RNq8L9I9aPxTtMod0kB0QABFcb1FYII/c2vpO6QOJ7zxB6ROKppi6UaqBN1/tu
Qjqunuzaz/zLop+b2IxUvwahACApW6yEuxnExIX5zOKR0LfiAjJMMQUSU6AbySId
4vgIIDJhaxXfXoWPeMUkt1MyZsHZenFbNcX9c+lgIbWmOqOyy+A+D8oUx4XYnhR4
mzBVB0NPVJjtOER1umOiGLWaouZh9UrbAtaA7eTzbuALTRrNC0VYUOSgjSbAWsHr
EymiUuAgSTK0sFKdJuBkJMKqV9zJgEdzLE2V2HJmmWi33v19HGz1prgwIm4QOFT6
punVIBbQxE0PYbKIcM1erLnzwVmSpHNoby7RmEbo1cG473ynnpJEOL1C3U0L1qtt
c2JRJbT5mKGXWzu60FSkFReoY9KPpK8zOkQMjtugQl7y9kNha81+2tVEHrP/xn7E
KseJPmmDfypapJIEbeEWpZvCWesFAchRh8cv5KeOZw73+2XJ5+W+IWyc5e+4OC29
q/J8Hf7nzoWpF9+JYlDeOOIvuLyWNLcrCOOpesAGkBZugZAyqtLdz3VEWUr+IbpN
i6JR5YjSqXDVbiq3KQoZclFMIFzN7vnpvarZbnrcSLdBW0id1y70e+QDO7/SFOuU
X9bu95jW5hMr5V1IAh9Ps62jq+7fqBFPZy/HWAIhNyq2sfmsGfaFbwEE841A44NE
6vHLeyWbFEShgmOXHcYVaj1hQNPa91I+Ljj3vAOEcHcx7uSMpam7lxiogiqWjBjr
XkwrlpHMPHu8xAgh8BtrnkzMGrHYUHbfQk797Skfv9mjuUwjyQSxIuYzGu8jhw7p
TCUaFotZu8YcWHnEynHVx7TBdqOayzEoW/5kbUs98TClNvQD0NYxRXn49GY5TQeU
LOLNjkU9zdYfQHuKP6O9NumVW5IwUieAPTrMzDgohiEFNjF6IDwoXAEaBwBTsrDR
TzpwpVigjqUxlxmcyo5kDsBqZ8zG6DAEDcFTQQCn6T/mlS6m+2ou19wqdTS6xQdB
BmortFzpkB4cJkjXQabdihOrl1qTea9ZI5/s+iJ1w9Pd8gi2wbfYb5neuz9eYs5L
tX73Vucz0Mbj+0ANa9xxjIEemQy7LO+AoGsht42uIIjJNt6pwCg5Ngcw5DUqd/06
fBfVVx0TaTn1g81Ki4XVAnl2KCfqLhG0n7xvERXa73GYx/RzB4rRxp/XgHATN8SS
fgzSMJajyiySE2h7bgL7QvuF1vR/4BBA3d0y/Omo5Z7CGRiAeY789sKBE96sfHUe
vU7zxX2KV/icW+MSRBpk0M5DXx3P1Kgflr471G1vvww4826Wyuxh4yK2W7bVry1u
cxi5pNea0S8dNv5cMtOM4KSf4YNuUcekwEqoSVVTqV9MbBtYsS8/M6Q90Pf9/jhh
ypKdRAHoIt3OHMb1KYZEzZxfftMueNWcN5rOSNzHiJURQ+q5KO7HDYVLQXAl+06w
EiekfpaE+Bert/EnTLOemUI3/w4wg9jDiNj9NLCnwARHmtgsUAdUhgeET7jIvkYx
WQxcopa8kBFAn5v8Y2ZDg0Xiyi/RD8G+BwML+fQPvNvGw20h6a4uVxKOE5RHMvj1
1blPuVCaIc+IKIViipcy9ULFxH9OgCjYQDD1adaOdRfT5Rbwsq/NAUubvozIIeCS
cU3qQZ7nmjJo0ssR037an7ZUl7Nsljid/Bo0YCHV/i9bpyRhQhfjpmqKUMV8CU+s
Sy/59DPh+gT2QDe8+Vs8ZoU7Qb5iuRma1PtNCIVDvH6nPNaAvUegy5JsQUW5iXxr
CSmSW09jWMyAov7/ikAHIpErmn+JenrLssf3FNgXQuU0jt4cMXeAltAeZBQHmsAi
s2bfZgkPOibRVGO5ovYlgsB27M4L/DF7NygHslAyUsEyN7QJAtcrzwHjv6xCi90O
ENjARj0LHKpsFMmVxQArRc9wobWug2E5tTi5mTiTf0ql9kuhQ2xnGSpR645/7u9x
GLFbjEtodj5SBUo49scK2pa5rSJLxmC9FK7Rolq29uFa4R3esCjY7GusHOjwhbg3
VydtxFSphUPP9ZkN04pg8iZCdcNkGEPsn5yM1l4dH4EPMO5dGQyY0P745d/TkrPa
rplVFNT5bohWMEZGH5ywJsyVaFAFkmkSGoqqEb1ZdjbY2FK3XmsivdBbE2dBmvyd
cEfYHC5k2sJ2fzkLoCLKensmbwVls3h8c1TwAAcage5F76Rs9sBQMufa2eXbtCV5
VvnLeI28cqr1mqcxsoaqBrTE6TEqvM654hn1PT6OKbyyz1z9gXU4QGmww+f7+GK9
DjhaAFHtSMgZ1DHHHndFIunIdQqWIMXbJhLr+djd30YlQgK4OmpbFdkytEyAJQ9r
HUxILE+WRs+Mwuk9rh3OaeMQK5jfD+5XnZW0cX3dU/QtAOY+4O425g8Wcmgku+u7
U9Nl5uxYBDLwZhKZG27mXww9/DoB0WYXe7R3q+iSPZFsIta/jiuHiFtHul9hHNSJ
vHduG2YGboGY8GH87ODDP/cKflVaGjHMEbzCyvu2MYUpTWWAgQNwrmtYBKckNY9i
o6Oz+ploBLLDbTnspmJpMOATcOwOGrvZ2GmvuaVhBHgt87+wOz3weQt5SGNNKtCC
eBkBUvtxPRFuTBEKF/EZFMlDYZwI/lgXIDNCszKz1dDFiAA6StXBM71BeLX+iGJ4
CCuu8HkqiRNEt28e8OXHObP4oQH5oJukdJNmXuohe8OflCv7jI4VWLjRQnVGqteo
PtOi2rueesogboHxqUKEyTwwLYHtLcd1qWKzj6WkxYMZMRAj7yWbC2I35tGE6ZQf
o10DFxsmPM0i8o358wwMje2n6n1NXrilpYb9xovzUvuQTv5GWFDkQC7PgGTj6acn
wamEVUeA5Ybwp2mmrgPHspcUD8FmKPSUj7VLlm0/g1bMXjq0engVOdEjP+YUB2Bp
Eb6MBXOr2tAP5NUre20MmJ8KUExhov4j74/YY589aZ8KYa9v5YW1FVlPR/XYeRgN
4n58lYW/eK1PTgUINlviS8xzPGPSbtlyxUCq4LFqbCCW5dGTpJUdjqiQAyUrp6YA
VkWcpluUARDCbhQBijFpXZOEOBYtQmCgBf1ZwNJheMi2MNFh9Lm4r5Mb5oankyRM
kHO9rwDtV2DmSGWu4vcgsh8p4QcJJeQ6W35N5w3ttTwP72qb1ka3wQjFadxw67qa
BXzHsiIs6BJ/w9Cdk0DJzlaown8aXqdx9h6LdW/RgMciOkcTkvVSJHRDk8PHHNPu
i9nl8sPzREVripJ0r8I7NTcylLaSfP0rLNwVWCm90j7DXu+ZHqw1m1oZFjD2pY9B
blOjU2lO8IvixrJNjFHLar56rgA2wG+P9k7u/yO8V3czO7jM4cKPwoZIJvOuXzxd
d3GQdw8qDZXcR9R/QfcYbXA4jozY/mK0sgi0o3lzg/iclQeAf5XNpg9Aq7Q6sg6W
f+H0tINjZraq+GU5y5ViGOtjnLabKQOy8qDuqeDJsM4CYB39gsNmQJtCZBpV8asi
ly+GjSqczVKpS2J7nfNKcFh+fSJJFYXI2vZi/0Vk72QFyQD7uKTsD8gTbbMRk/pJ
EkIBVFJ5Xcrpyj6TiCkR+CurMmszMBkmvKfUH50NL0GkPIJP1zXlp1f7lx7RnlVv
3DuKtQVHHH1nbMaJLttPe72+w0HQ7YF6bmucd1f7wV57RCUdD8viu6COK4AvFP5u
bSHiK+lT2PV6JBTRQzZw5vXWL7rFxnIncTTehA+UPguZ5l/CqhRGUAa+A0M3iDBW
O5DBaOVcDFTR90EBJ/RVYDNRxgYU0z2uRF0ChlEpJX68DbrBANIwQ4tQLZMNawTT
NvwDvbGCEuGNvMuFA906wycl/W7vv8yLWi6ebOecgzeUFCofJlFORFoQPYCUnZFm
8zL028T6SYDx9RzjhNpZAO8iDh5bbq8fB7H96cXNmUcBrxcK0WHIM5rGu8zWw/Nh
2/+E1mIFcuCRiokz7xnx0NeKDsKE5AcKSvL12pX2lRD2/kv6QKloIeMveBzFJsgF
py0tXgBbPA4/pZrSIx/hLjd7iJfPKl4C4Dw93Dnep6pAFcs6YB+cf5//FR+K9HtU
lUjjPDZNdL6FXBUmjF3kxOqvXuFgxxg4+rDAnDV0cF3X/V4bJ9OWY5vA1Mjy049X
c17o1GTXmMrdpxjymomhTA9zOBHxUnP0JStXhFyAP220TRsQ7LhUG52/n22OGHEr
UvighJSO2WJzeNmTVq0tbZjVXdLu7dsKb2PY6uNhFuO8aBNghxYeHbc4CvWRBQ8O
GYyn0VZgdVS27QKkIWf2UPsi2Rob7cMzwtHF00bsFqlxyrVB2HQSA64Oc0zc8+xs
+uLjaffFJ8vqCz/1Yg+KiXx6bvM4RmPb9JX5IGvNR4+SaWzwzXLonMoU/E/Z99PY
JEIpx/kg3qto9fCWvhMiowiJylI3yHbMa0RV7DJG56AAQPbNjDaBoXtTA/lA/1Dn
xEErCCvGogyKG3nVWRgS8eo4qR6yRCthFXZwL/2Dt1O0PkOs/lqpYOKcZ5Y/3WTp
v2sS1bRhpBLkuiJlgnNhZ2oXToATo6coVj5gOHYnKU35EwOuxfHJqUkEn87rvdgR
+mQeTx95cUJfgzqMuZw3aWFk4LdPMs6TEt8JIJ6Qf2xRTb9nZJNGojmV/unapae2
Q7mrR6GfBMjbh7BWJ7lUoRAPxRX8XvsvxwqaGvd4RKtJG4vHRStNi6gic/eZqcPo
H33QUezxj0S+NlIQrgknqLgDFaITOxGEPhh3eyU7RzmLhMOOEmmRzJXGjvVV4G8t
RZeXuJrJRRxRqI5d5J9V1FJBRA471DLFifU8xLfKaH8zaI0wqKIvc42sT/sS6pP+
GXDL9y//5flRjIIGvy8qNkt1czIHyjeLBq68Iy57seYMILiiglYjrewoV8vbQpvy
/p9TA0SSzMGrNeT9JZuaw7Y1XROhbGQuAELxsxSwvYgUCseQFHePE8C7mRrWnqvd
2RVaP4emhlxWSEv9oORlBoPdSOVkfZ2O+7iQs6HijsvKXyJkyK7BtZq/MK6AcY62
11ra/5wxDpC4LuMn713kntPiTccRS2Qx8q5tU07rQrfAIBFJO9jd3+WXHb47K9jN
tUS8MaXYbqlQ9foXE5BuYPl5dRv/l6X82gs7SOwc8YbljA2/aPMSUgzrAGZZhmhU
/EEYzIR0Rs4S5gyovMJdVry/VqCBym3y+FWdD2PWbC64CmW5Y+6E4ZxwmmyybGPw
JcSRTeJk+LxqYy1P2j2bxlO5+2gxHZ8YZQwyszOGVIa75p/WOISBZ6vZDSQYxQsb
xvjsd4lL29dfIyiQTSnZIxCq5cKVf2HbsYbbCfNlVWuv65scz31ZTPsl1A55N3eK
pTP5IvwxF91uc3xTRPYwYSZ+wFlEwYAJeeaaoeKG2OozmRDaZG4cTNy1tXBqZFOY
uZqE/+n+N0ug8IXUnWJ4zp4CB2EIb7g8dVAmRcjkjLMtAwnXR+iDFUZZBIcBLGvZ
tSlBQBTfI7kim1NOis3sTHav4M0iq2Gj3M9rta1eH5kPL2ZNUlgMqEkzwub3Kao3
VqL0Y4IXQTbxcFrAO55FYRu4JCQdf2hGBLcNAqXOAW1lhYHMDhyuI6vJOdacihDw
5qqdSl4/EfedqpLYB0UHJDbSlP0P4Z20OOzmTsK1f/xn+X1D/4RktXexWRCybRVg
Q8MkqRx675aBpy9I07Z1b6NXahr2JoS3e1v13I6btRJs9hJZ9oyQ4QWjqJs9fPPC
7nLPbJsvz13HZpoy9tmbyI/jyhR9v+z6TStjBkGif0rlgRI8FGK6F4XatNher3XB
rVl1Lrl8ExzhdS8VpuEniZEkQs6DBqPgldGIieB4My75JBGzI3qjSG6N+yhumk9C
s8RVD+ki4GhtGVeo/xmFeJbcUQIF1juEmuDBkBJF2OjK+4XQToru48N/taz/uDxs
GeHIhhrlaXO//j7HjdFzpfqdLf7w0ZY8v7TIW3MPqFHh5xw52cWFYQCJ6627Urm0
sy+0ziOusBHDHklnmnV8gMLSGGfPYtIr6ue7K8JFTv7+7oFE0cDvmswY41o/PPhY
UWXDUyirWWzWCFPiIeao8SQgPMHK2AEBRXQw3slqhGbAGwx5AmmLbNa0h5lrOwGr
DQXSz8vIRgJK1HZrOAyjzXuqCUm0OZ9+cQ7fYSTPdmxNZa/2z53VhBSZLpkMXOPt
3+H8M4brnzIWkWNlQRuHFJWgDNqXmdzFcFZP/zYLkPBKwPuuh84WPQHJCfr8gFPq
LwYh1GRoNHn+j2DyVDiAZdRZwrEE9f58Y+BYH+q5ghtTL7VaLWVsTjTg8wvZg+Zs
fi7A31P7o0ro/D4vJdUZ/R2z+svwO4Saju+ub0Py6MXDIWT7pmAJIesn0qP8jv3a
h3+ZQpJ2H3vU19PKWMGvoR9K294ImrWDHnjZccdEvvoMFMyOlBLQkdl2z1s8tgtl
rv1kgBbi23clI7b3Dz1Qk58nF+NN480XTMVvlgIZ9xKuoaS1TyVZAbUxjha/Qohd
azmeXyss7XTx/hsBweYnJeS5yKCI8Q/Hv+1cZtNIsivh2KuTlHYiNYH1N677/VIH
bGZ6vWmtQRX4a7CjPxHJbvl+6tZYLa5nJq4EEnVgCVrZdsx5j882Q4u2qsy4RRdI
cPcu+amp2YJIuRSsiTqD8R9c5EvxBA0E8zgT5T8+6sJgLoGFUd13R+BDbjXq3uuU
kxGds4eaT5VwuhL3QmibP6jdabiXY86gSlYFbj9x1wm/qkb9mK85NTo98y+Iikqv
Vf/Jiomrv5YHxZJNLaoyR7fc+dQw5R3K4rYclPwPA6lpKFP0vvMm/EhHYZdRXb7b
uZiFNdrN817w1FkzNgqUDIsUh11xh1/nhyL/IvZNWdHLecG8GYFqrVrNWxSnf1f/
Gj60lSC/mBqDnIiAAmumqrkbhsd3UbdlhbfcbxnaVkAEuW+1+YavoAGbLJkXvHmc
pdQf+q30EmGT6GRv58LaItWYTqZTbAF76LsccB7zAcGXdQ6hPy0IwxjUSwAAMbAC
G5iEWepYgBXePOlPechikbFIAGo0tinvdvQcmrmjPBwJYbAzjzE+gKYGwbTBq83V
QW+vCU3pc+/B2tlafR5uH/VExjfMuljaHLvYbuQID0jZSCHXQUqJestlp5ppScoQ
v+d31vrHoSTDTOUGozRtx3NX3ZIBpCxb7LIzAwLd8zF6+1HukgwOeDfrF0XuonAg
72Ic9oICFFeNn58dAlnn1Tq9XiRgQHZHzB+nuNxz8XgfTTa5VouuR56TYYfE9W1D
bufxWuX05TgbHGr7snkQGcDHgH3ry+ImjKByqCK1uRxiAfTpysJ5p8xzJK83dOK8
DrlnrMfB6he+gd7JCDVo6P6vLPd7woeQTzf1JhnluVMCmsWmbMco/UV2nqM8EhTE
dYV2RNYX8EV0MLZ3a8eVFOXNta39NxuKeRMQN5ht+SFYb5ZvO4E/Hcpr14cp/GJs
FwYVml+cwzsk1G4FbYMrCFgFWMbS0B0FFan4AknArXiIXqWfuSr0uWDPIAVCHmN6
mAc7jJlp/rUpP/0z0fV2BiEWZALmcymVuuVYxiPNkOiCJEIEkvv6GM3qM2CbCGHN
TWoodQYZ/NbBjI0SIpqJd5bJpUOxaIv+aVOPZfjFCx8/tZqLLH/AxZVT1buiuFXR
rrbeW5utn/j5Rtf7I3rLfYgVWUpuVDODpdmdCIOp2NrcGyTEfKHYz0a156hEmLiU
bOp+QWvLwHZMPscUcUt7Cs8J5/n4OeR1m3olQavm+Jz31MPCatV6B7zobx4UADb4
kBRcExGJa9R1KkO/9thEzsjOBWWjcA/faq8KotbNsoO9HlPWb782JOh+FNmHwipz
08zK5o95o6rKRiwJAKjl5wEXt4Z2WE9phh8JP28BgYYLpVBJ104S479FSXmOOhHT
SYLDsFwZ77u3/8X/X4Uc1KrqZL1whHBFeurAkMELTTex9kX5JaNnVI4J5jtppkvJ
l8NfXxitJ9g7RrTMp6LHTY8/LrSABInc7sXuJhuCR/z7LQmYOgQnRpftKx8Dkdix
PJIyDQ7GrijF6zjjnuiq7vYm0HjbSJZCo93+/B5K8SD08UNEzx2BzSPgBh1LKQqp
POqU9EhGCeL03sAMJ/jqAb0suxp2cyWzXx4pp9eACW9K0qhNigLamjawxaJYmn1i
6o6EJdtq1qMbfXf9h6W3hp7qR+iyS57Yms2gJFGQRlr9CYakWzfNlF4ckHEIkxFf
H6zCxzpwI7j4TM0BTGX+iCi/nj7iV2n3aigwVJkZAS98FpckzPDKovRXxpJbOBW1
B5k4Wc32L3IkM+c17E7pZzieTm2cKGQo/uC1yY8nnzkE1smbUPUHEByIbWIMxpdv
CpMR3I3s7eH8zA8G91jhSaROoSCU21sLYM8jcLRnnnc0D+bw6bLkPxKXBv9slWjF
/L7yxSovDp1rP+QBw3Pw3BgzgcX9tqAh09LZUNY0MhsUBXVe9b/SCXAb07aMHsKC
I3W3fNmXKh2S/wVHQvSrt/AQTxpdg0dxATCi4ly6P0P01q7CUFKqrFe1MuFHLa4C
2yLWi9N9HVSfNM+kkztwDMgnXDRqBhEcVaox58rrlGayiwW/BpwWW0Vku0N68F8m
9zpgYklff8e2A5ygj/RQUjHx2um2xFJurJTaz0TXpMkvGaynktP8tWzWP3CtdUOp
5MiBFP3n2zAfK+Xwnlt8BaTZrzBp6J2S2Eyqx48bdvr9DHs8p26cnl+gMnxfWu9i
ow6A4f/eQXR5G6CxpFJBUuhA4nmqXy71zpxpsYijsv2DkIJis12+dCBoIQI1VJCH
VqUn9QxFcYzrXKiiBknfZsIWj1Yp8CbdOlnfAUYvk1cHV6JbRYefsFvM7I0JXsbY
SfjQHQDd0J3nXn5xJ6Vi8j3n/5spvam8KnZstoaLd3JayBCX6T1RpwE6ZOUld1oN
so0jgQBNjrV1mRFx+cfK/EayRYErxas5WSaOOMBAmxO+7ohCT6FBEQUwnEuRLUdI
pwrechHlD4dvcxJlFzVCexDTZqn0MufecXzsyxcgwvvGqv5lRotbY1aBoUF8qzkt
FnIf+c6fbEzrQYAvOLn4KX+vPgYJ5+FjG0rQfu04zW7Q3xeRhc+lIZY9kVUrpyJA
OjC527Vn1XUYYJBxtbzJxqRrR4FHeHf3J8kwrfq76hExBM2igIr9RG+5UovXIG4T
V1BHVz6oR5eHd5dScUTvB9ZhRt1ACt5QWlo1L4hN3FN/wQalo49v/q1QbWIViiSH
cG7p4q4y6fcvmSyzX2Vht6WKZuyXVxWRmikKAByObb5NuUaI5h8bwY7GiNDZK0sF
tZZ9HZRrK0FiislnHS/9+HCmt4tnQgZifbs6IhZ9HuryXhSr3hIjngJeLPGhIuCX
nUSw5d+dOylNhId/r/tu+Ryzl2HQiKEAVL/oHgOzLYE0dsf+WTWZVGFMU0oF3RAr
wPhRLqa0P+az/vtTli34bFfp622Fvq80d6ptfcA9s6C5Dlfr9dzmhBOOP6L+qNBC
waocpgWPGkzHElclmPbYGFYZsWBukBf4BFL3nzRiAsbXSR6mUHPWDEiPgOrGSYM1
KIbyrntGgOnBsvRVJ9PXyexU9OZaKezzqmwSD2AjQMgTF/G0I9XSdTRNuewNadbm
2eNiF5JWpaTPg9kqFMoWk0tbHdHpgoeALGja1TUWF2c380e931ZHu2+85RlW/e1/
tF+XEETGtd/BZg6SKsLgSR8vNo4nbL6e9+in8ZIZv2QoMEltYohZtH3PCV67tvB+
POoc8Xr0J/Tl93dLroElI0CMCnAhvbD+scbTlbvGkZ/ICPLm/hjFJ2yCNMb+Lq3/
hugeyb1XEbEqM+qnQsAPXIcNlM3wiJBdAt8FAk1hJtnti7CXzyzy5rqSR3IojaAA
LDmyx08kQSb+6cXhMFUodu2NuaUju1R1syWx8TQULcZtduIcynKGeH1KpdMsv7jE
E5gD/aPNf5WkJ655ZECMFSG4i7uayJsAVU+4VldGFR2+hNT/kYLQZDDmi5H5hYHX
3yW5GNMZ6Mz/ADzhcYMTym/qULpAdnKn+P7FbwLx2qFHU2r3M2tUzh0HPuOzoQ+O
wyV5tgWa8hAWEOKXQsTu4DcDHkoUMoa6ljU2TpORP6C/oGLx7qCx0pc5b3yVRTwU
dMbOYkznSKQmy3tiDo+AwBx+U9P1n6C0+hZ892UX2cJeKV5CpZBYHYKGRTv1SGqQ
G7QVqkkUQS9UMIp5f0XIxjJLZVJrHisI6Xg8xpJnzbh9TQKuVrA4pHBzCWqq1skQ
JDMzZ45+P/TBGZi2t4uBAJTNvjW3TLVqiA7GARZSz78tCyta2ycsJ1GvA0pH9Hza
3Gn6+E48cW+TS6x5H26xiYCzFhIanKufIYCEeDplM9OZ5s+2AJkqG5HRIXP51ilk
p7eSzw25fEEx0YDSiwJLgLp3WA3++D89h7NdlD3M4+BVK0k1Tw6DKf4a4L6/9T/C
2FNWgHnxkouo4oUUqeZDVvfbWDvGT3+Nz/ihR4hRKyoazbkVk0GcwSSblbXGSIdF
plBYV2a9vQoZKw/5GZwrESXzIUrRO3R9kbSrWg+6hVYjjVyNhlsJoeRHeAdav4aB
mEi5sqqSrk2d+KT15FI9EHONIpgdL/yaLgTaU6/o0e/tSRyKohY5+2+xea2258/L
FMkp3cUCWT/argLWRqnmN7gtlO3u+CcUZzU+qUMX3tWV/4jhQmTqmI6j1pPL1eHX
xFQbgSvw46TrNAPzACGeMhy/d3cLhOsN8Kf7DVBkNwOY8d+9K7kZkp6oAAjb38lp
xANwFcxf5FhaEczk7bFAdj33b7oTMwDRXd4QICX3J4ebV2+7zVJ25oeAMrZ7D5GG
n3hehcxwClBSXMN8uhir5UBDV7Ne9oZWgen8Z92gO+QWLzEb0GtDqj6UCCsMvjZr
B4klTAvVbbLbSDUCvDFUZN3gK7LANosXvDgA9OtI+7WmbhT3c6dccPXH1TSK5MWT
QzK/Dcl23UonXFfcEGs8477U/IgtfQoE2msrdw/sSRaldX3gfIgtSjKJqELYWRSP
ldANX58+J5ZYfLjZZDcG41s4Ne0CRKV7hMTa4opwSNjIOYveZ9zyRDiUBbth8K/F
hlOFwWB+Gv/0VOUi/mwNA7EroDdWfxL3xGaxdzWTkCioF+pbKV2noMnaHqmBKl1e
HwjCjv5ssLh+uxIZuLCupGFIeKFRWI20CcvviP8bjRrTK/zhIRL85Ow8utB+d3Rl
WSR4T66HNRT8E1JnTVRqMMRwJNfGuF8k5Fevb0d2utRNYc2toZ/QUEypLGT5sDjh
RxPViGiBBKwaP+jOnBJkOSwOPgaWT1PDV40QVSJ70Nz5TRsHsINzYtTYPMJYyyu0
KCAqk+ytgt3L17//mVscYwLfLJXdlL0oKuv+gXS5aV33cKUbneZmM/ZW2zqKsnvW
wqt1qXhGLWlwjTX34W7KAM8+7PyVmlHqaZO10ugXRGUP4JraMzsiEt2ZA+ZMhc2r
qGp6g/UbSV5C9M7puVrzG8F4Kbh8oKC8VO0VXYaZ0xEeXjlS/oLfzgpoFmfLj04m
xRtQg5tx4HgxsWsuQwMRCgSPy6LR54/6atPXp7Rk0wrFI1rs7KcigpO6ZkWgS8G/
HdybVzRLalIA2VM1KHCQ6fqxZQ/FfUFmJxkg+TEZJ5ZyQaINlCeajU+1CfcmanwM
GYBnl999rWC6pPQUeTVofe+cpUll3qniZnBTPXnHUeq47ZIMO6EGG9ejhMXC4Joe
aKs7sH/iPX/SQ3wXtjR1bWj/boIF7zvrDRDXuLSD5IpdD8L1Bg+IrcMfK8aq06DE
+Kl2SllJJADxBN4SMOWk0yYGCWGTbNILs22DScVu38wSS04QYpskjnkfTARG075U
5pDeUb3THe9uuB3FlITOds724e+fyUc9Nj5aoV8Wk6GgurkQzQAQzcIlgdZvPzU4
EmyAgobQ1wN5bLehpRtAinYJnBfflhHXLTJCk0ztHxlGnW7YLODUTC9Az0I59fUi
N43mELtHMa75qqOoY7xROAxzJLj5worrpTyxW13W7be8+Y9SFdhImf46gMZpdli+
zQyChIpOBQo81hPYhcQOyKkBhsaSuHx7vpg/3ApMMqsErw+LFqqiC8X8GVMs6z5v
CjkKKIQw5GHdAzYeu2uSytf40sdWj/lIMmCL6GRaWlXAfOE0SYeJGO+9xB4F82+a
2reP1MRsSZmerKSaqbrVWEpXoZvQ686ezPTjGnddL5qSsjwUwO8fL56IfH9MpE7g
sUIL9tWUV5TztmJvRp9pA6GdaGwWxrhp9Hr+a3JBtgBw4A8/B6xPatpsC5NrNjvj
8Rclda6F0vkeDS78JiHCJW9CO4rOgZ2xkhqZX0mwNTbApimx84gsBA9Z3/fB9HdE
vV+qXAmDz03W1y7V7aG/zDX/wXDs/a7JtNHCKEENNjMbFdlfJgYXTBmB5klcpcCd
El1ZHaX9rurfe7PaTcQRBnFflvQsaVnw9Bw8M4ydY3e2+4ExjgjbRTEirp57l2DR
uXi2Zn1/lv7ScDJaCzEPX1IDHS8v6HBK/cr2BpjS0ngStPWv1QRPlxhlBOthniTU
o0OK6o4LF4ADVtaKPGV5Qcd9XZZ+MXp4b29Szsl72SkMPCwPi0iotWf75eEHELi3
e9jIL8T3WU4OQENUeu/4mTY42XnB7fRlAy0I/Hbxib+E0qhWSMboymRDglhDAuZ6
zkbbgFO6lfWYyQx6BqR6bEA9gfh3oLHbu6i+J9rWR1p2XZYnODGv+Kumlaonkabt
yrkEF+5XLL6+sXmk6VCAQCE9WMQ0LCV9uSRxR5QgxyJDsooWr8Wuu1O+Gdas4RLl
T3HV/Y8u9Dgq3N/Ewd48Uv8lt6gL4aJzm5axM89V0SGjorExitXvwDDwp8XMEgZz
Lg8WNbzW/NegeuFJDcyC1RwSg1ZoZ5hdp3/1CAYeq7oDBGLick6UbWt7dawMrtOx
MoYR6qbEzlurBCQqOPMkm6KB7so4Xmilm9H1yYc4OjwOIj1OB90Yc6m6+9VZNn0G
09cEPrp11RYE+S7Z9mxqUhSCnMLfVxZI6LwXGrvqksH4XRWfePEWQpfG8Lz2J49x
BGPi/3YrHkgjGNMcy2dsglUJqY0vVs04BO3BVJobowzNYgaiIaBJ611o44DAayYN
Yll0DhkUyE+IXRhGC12Iba/Druj1cEiRcPXjPmunSBxmxKbSTZKM2WwclHBs0wuV
rw/o76YCgZcCzwDpj+B82IMQ01e/pxFIeMUkkLKvZla3jm+Lj2ct3OIyMX5Dd3EQ
7IW/pzQRMyiLc700xo0BDAzx0j6XCZ9ZjrnoY1FevdApBTtu0bcWoSxcbgaN2bXa
nnkbl3au77i+ODU73b6ZVE94mdwhLA0cPf9Tp2mx71fNJa+h+huw3lZNutcO+lzg
FdUgQyuwEYXh7750fY0uHaM4/qUNEIY24nwyqyIT0exSQ2arQXI5X0vPFYK8ZPWx
EHW5vsnZEZKXHuVLujqdoldxJdU+7XnvByil7xdmFAlWP5AiMcFjJbamrfFtSQxI
ik6OmcKJL2w7GWyBzCDFPSX0pgPjfFpC7m3Xaq27UPxHzBi2N9y24KT5JRqlqE/r
z0+3Oy7fGGNkRc7sy82nL3dTK99xHbIwX1aIv1cQJ6tWcMDEB/Xz5DFe4+EoS7aR
og4fIPDPxPgPoSPftji9cFA737A2f4xNBR0tqG8zXr+6KtcFGVtnVw0cc0dv4YM4
yXHqgnuNnnjOjnFcg8Wc4hzHBoF5PB/6lLYjMgjRHs88uEqFpDaqlPxBUEyMPXtY
LYsJfWu4s5RgX/SDbERMJxdfkc0u+t+zjDyKsDup5y2bMXstUFgFIfii5wWB3jqE
ZmNqE6jNoe1sB3VTY8fVwW/JSz565AlrtvwFvfVrZm21U9689tismwgQGWlbKWj3
R8hXEmxjHWb1t9nB//a91ZOqD79QdkP/3DVwVFGajHdeHtIDZ4eWqqNW1DdzBEy3
whTYyvyyi7FlSSh3T86WNN8vWsDzOA0ds4wcfP9iwNb3+LkQYS0Y08xTVOtATDh/
ENl4oVszim32Yt5b/EI6/x8z5iuoYY+N92qMOgUTpCyAGIanx+KhVOVsam5uWyxt
rNmHCS8sYQAJ96zV+9jO2n4XrneBCmX2rVqmUIgx6KnJrj+9hD9ql8kzHU6FhtVL
iscNXikTAaWPPtpAIL1lRs1+0P4e3hcBqbh3Ti1+crdCCMvkZDh0IqBzXPMGozYI
6Ixm2mfNm8Cu0X7FJJdcUsOVYyuJSRc8H8ZEq15T5dymHuinMH3SG8lYhR+jJHno
ild9hKj6abrnj4WXDgRx2cspajM5crhW6YLpKIjYDrzT13dklkEgoLP7WkhmZs8g
WEfuLCB1rbqfe+7k/h4P97Pnws5EqwZvioTGruumqyXoqmtfR/n6xZ5Bu8H5Ji2F
0C+fodqb4Dlil630PBiS/azDqtCK00p3aJXDvdZL54fZrXORo7/o4dLcr43AIFvc
thupM0OvOJJG1/2Y75qhOTP2s4zE0vxMzD12zuq5Vb5sqzyDzsDz373CNlT6xOi0
SGKI2HV0sE0/aRT9Q7h5s0lBHvX1oav52BikYaxhFtYkG+1NxWdvR/OusqHJbIkD
V/jpgespGP6BwWhoJKzFJ+MVaF4sifSvpFo0ZbPmLheV2lP+MDajIcQDK25Ze2hj
7tak5lxCjE3Q092E/dYWrFNjrdfTY9dNNEG2++J3XRX8h17miUVlVtLkosQ0+Fzk
5mwWfVOagAfMTwnVykfZoJWhRwqJTMRbSkreDCu3UzTXR4KgfOlsm6zNMp0wQYYp
Xc5DyZ3FgcTMkIvGYxrdjokTvFjuUIXKyKHhSmG5F4XPIYtnfRQ/WuQGRLq3ogTj
+V93WKc4mArOb4IIvSfpTtlkZtCxqBVFN7wps8ifZOASkVWds+O8IYCzG2XnrWE0
HkOgPcvAYCVKvexfRxGRTD2PLD0SnJO4iOGwZjxgULsL1RgSDJUj5up1Lv7Z0oe8
Gmr5n47ZGR10M6+aCCKhgb/fWttyTGwDj/sYGL/aqYy26jX71ei/I7+Mnns8jWqX
6boiaUFxUY0GT64PCTSl4acYuuuMnWIA1Uc1zrvDt64V+Oq7E+pHO8KCDhiNZfh2
9W3bnFTKrBSfmEJ7ETjYxSTqKCn0mWfgBRcgqstJ5MIwLz1FShc7nhpv0r5ndjwE
XS2DsE+mUCRrCC7J7Nda6O9ZQmohETJo05J/LnJlD5mExhkE0qj9+iDTUmNQCPo0
fa8wTbO5pGKTyMDyyvVaAjgki1eQxSr+bi8hrVKbLctXtBgSadU18nCLkrU4w6Wj
y+/UOmxua7nj1gYHJN8NwFQStOYgYP5IBpdmgzgUh3O01YVTQT0q4/d9r3uivC+d
SsiiLgYUe/r+CzHxZ9tyob7EJpZsF9cB3V+PhIKaTUmW4dBDWOWrA22Z5GAqNYbb
CEj7uZgEcjmIxAUGZzToOfoUmKp/b3/PAA9iTIaim7RrvdLjL1tDkNx06dd2QI1m
DWOJJvkBD6qaheKRQoAOp324tQ2NQTV6vDc6FegCiM58U0//Wb5XPbrL92IVB6aP
0Sxsj53oWWSATHJK2gFS/hEMq5ADnfhQOSvBQ35dmy94MG4y3Nc4Ema2fp3zZxVJ
Xgutrkcd2S7QjjhbfVc2N6ufKTFvUxOa7I0pmTBr1Aw/7/1I2HWlKG8xPRBPMJcg
5NbVqdtYJu0po6Ta13JmcLOHX7stdmFSDWHQaZb3wmV0NVCpHjF92hxIKplUQZH/
9qUeBKBODGXKJO3oEh7pgpgaDzPmT1k4arKCG+1cTeA2YoLfb3WD/NrZenlKFyVT
K6qtVi5G2naf3onbsHFXHsb1kX4/1O1MKJK0Ch2vKUZvaFckb467Lcy3aczssO6o
PfGefsU2Aw4KOye8REllVN1IreNr/UzBOZPAaqmskU8zAfottvvlnbF7PKKBtrhh
Mwr0jhQ7ng8f3fI79oYMK1AdZZT185rxWwmqq1ZumtMnaKQKNHQHXB07GmSYadTy
qxmEicl63kodA5LfGk6gnz8vkBNWwaETjF0DStbr/e6g+q8f2M/EeOpECjaQycnx
sFHqO3HIoxphUTQMFEKaxBJJBnfHiEJ3AFkKzPzK0MydqSpeKGMr5jp0VzLCqfaZ
hWXh22MzVIazPLo0AMKwPrIGeChbRxK9y3aNiyEm55KETP/rlua78YseShYoDFwB
duqZJ2I51MIWkAdwCWcQ6nN4dKKFGxkhsT8MGFqy5FD4SvIoH1E/rm8/nGQNUmxk
2FFcOtLEcX2te35+CNooU543tK3W0lorKXHtqlEJI5w0VH4jToXS7mBbfJZp6zWK
hC3uQlPuOc9kRGEKy6EedL/xfEryZtR9qbgMy8XbfRY8xQG+X1Q18ie0XLSquqim
dA+4vF144aB8bar3EsDJ4AFhL2vbKyFIzDol0wBj91MKjhgFqs9qckOjzTTyafGy
vSUx/v01QnYLZsNmOgXMFu27psR8qQSQy/qajQcI+G8P0G9Pyei0LGyjXJRkMczU
MDJpHzL7x7CIVLvNQamS6RGlN01cmc0bpFZMiZzSGdYV+7E3atrzyZnyZouMPLuO
TFp33uIgjC9m9a6Dc8tt7hsSmky4WwuPisn+UxnJ3USOMf6A1+EDI1/xcB1Jfnj9
vnA8Ra/q9di22RvH57nvR54C+4xE9I43tOXUFucdZc7kcT4PIlS+Z04Vek/bFB/P
vS7gsx28ejZvLJYUCyBW4eei1ppyNkEuDpFqxSM+qG7gRhDZpq5/rvJbrUWof7Zx
D+R/jvGQLTYmwpLv22lOvkY4SACswwd1YKOZ5K1etrdmazY/WHSOb4VDq1+vqjye
Iyo04/D1GVVTht5+coHj5mqMZmBbJ/yQnn5P//gJyDLXRbRl1elMbZt223Kh0uZL
OLekBvgx7jIWjJx4gczxPnQiLvJx1/zs3mqqdDy0BdEPQcg5HpkC1lDjs7Jig9FK
n1h8sUYakbG2/yh+2phu9MrR1yNa2WZbxe7gLZ3kT1dIeqLs4N0uy2c7l9MfFdi5
WeaoSPoMkyTWPmzG6rAVlWWtDEuTTHzI8BUFD0CqX8q/s3qObXiGrFoEmFS4NG7/
ivlaoo4aom5SzDPumdc9xY4nNswiHZh6N587BCfbQnqKeNY+rQzShm8eM1qE0mbL
/34oFa+8dm1iUl/4JeGJ9s2gA1KFVD6IrQjjE6XuZkqg+on7THrqOn9bcF/4ZnBh
KPGR0JPyf4poQ0xKupBM6RFUafR9MoiRH5koZm27oNeq6qzFMQ9yO5sbbC1yHS0X
G7r3/WmcXoljZIRXk0yJip6W2gjSD7VCYWpIHIPPt135x9N6ms1+RJ5ZvKmdl/ZB
G/TKD4SEe0lMC6HvtYenOl2LEAWeoLkRyUzQjynRPG9/QW/8fNxOMT+zPj2/7TgU
RnEBgcXJtP9KWRk8w41ECb0DaF8T7CZPy/fCVPGjMhN4lczbvWUtCaU0c7zYsYYt
FOzT1a0KSjUw545UlfMKbDNmqw25KWjVfHdhMcO5ou/OLWQkp6d2j+Mp1fLLy3jp
zb1gSvmlJdqTblWKtVHdymRrNrNVmUaDE+UggiDLqXb8u5cyTQfEHPnZmAZDbOh6
REv9zvFfGV1AyV4rJZqTpL+kNvaHywf7gDY5F/3gHlsA385UlM6OpQBo4pj7wSJr
/rksvLzsnHYV6kYCVMMK/Ej3fqArQl4tl+BY8mAnYDSRYTiriOceggT5xHAhLyu2
z8LCNl+Fv8ieM20F3Uzxu0pCsvmYKxOBAnV8waqNt9mHc709Pnm/jANWs8CLHMPb
1lToL9V7yYxu/AoB4ysXsq9MSgx/Wv/leYKH/yzZNOoaKO5YuFVqrUhZ3gTcAHc+
f3MnVJKDMIqpKsHKGt3HvdPJBH24ws1P76n5tkPcXIszwWjGQ6DdtY8h14ezxpkC
IAKWZPayajFoLVlKyMBNRRLLL4hNo6w6+cQIYgsYm3FqO0zmrsG5G6dWWFkO5cPN
nj3Y8FPpR/p8a+Z9A6ZOrJgeMNrZphWrvq94rJ/lNE3Kc/LHVEe2DRou6ooch7vo
mhVo0y4xewe427RoDP8G5nBLiUCCvgt98OaUSsDAQ9IvXvxispikjgxcojeKzgtG
btsOONotkhV4o+kIhnqhyJ9DddezKzXaYeSzmMWTaIUOBdIrb31hQCyMC25UXIIk
E8v/dIizkEMMvU0SJWlJDZ+EJJ7hh7kQM0LSZDNAHkRQrsdirNCgPiyk2R3Y1sVi
x1aY+PanW48CsR7BTeHQYuuR8arkrGb+pVt2pHpybuSu0BALkwXGZYjx73ajuKB3
1YqwoHHMKK42sWw4AMoYgkVEnzG5qyIMA5wFm/QwmW9zx+LjEA2vevUhRievUWL7
MpTyY2ZmXWiRQK8YaWLgT1xkAyp2nybj3DMU3V2lJkUjE2/h2Pr/9taqlDKxuDTi
OiIfxiTYyR3LEY3r8GZRwQ8VitFa6msFfskvW6igjrKDjdM6dSun8MWU7+3uKAzf
TEDsiWh+JtgAD+dJqwpcrkF9j+geN7oJARMXOnCJyywVyfx0WWdSZj5rfezDSFGe
619ZjvAX6P2q9vEZeT/KukkBWPiu9TEmfSKEYYM0UYv5/aKLpAJUyYE1rj2SIC9o
5e0IRQrUq1rFTVRYnsMZr6rrCckH1EHkVjfHAcwI3OkY3FKy7fu09Bwvt79SUuV8
yAG/TKRb6MzhRNAUrjRJWelJ+KAWe+JebGJP38/u9tIIx5myibaSfMjzBKrH/XbG
l/qrGtNc22U6SsSHTfRGRH6biw1rbf7a8KUeHpl5HJDy32yVzVKLxa6zwaue6m0c
2Is6LJZw4taZQVngabyqDZZsoL94xYTTVCTWfdlalhPHAWL8MJ/D0kBC5H7S1COJ
zZlQIqiyJ01KRvSbXr+GyULkD3nm5vJ/vp5OWpQnw5/PZd4ipXw7gGXZzrvFRbEH
GhUANdUEFGyKAW9FDAv9rsSDkffdz2KFwb6CX82u6VIPa0U5GXtTidUsYOivjCNh
9ytUER/YQ+8A7K70+tdU4vaButJNAhlQv85FN2xy9OhrdnWQX1RNbvH0r0sgJ5D6
XgG2sqVWqTvqrn0clinn0e0lxgEiFSaLRgB83CC10vkYAxajochMW/kJBa/hwOjH
mGuDEHRFTpszIyysitZD+7ksyQBWCBTsmPz8xBKjbp804lg+upM9MlnmdBJHS2TZ
/4HCU/e2dKvv7m4qy0ZzXsKlVy52Qc3cgPORXSB+pem9/KP/4VSpCyjdXTfUkyal
ZNYu8/mT4HAAdVhyY8E8LRxi03Itj3S57F4b1AdkGG0WNbrz6M+GT62nXUgiXRr4
V34I+dyiibXkyagTG9EOLd41IwlURi+3VixcJ2KU0qa5vTKTGrsi0dXaHV5yGq7a
YOeXER/fxAltd50OlWIGy8wp2SeZEDRlZ+7irPSJgyT1RQrL72gxldMiZYWJ66s8
3nxOKkQAfXQ8Tpaphi//LKUHSTc/hzZ5Z0AnmjMmoE+sIrNSV2yppOEwJsPf576a
5mf9VaQHISzdncRwruKlvLSCb64ADVqhVO0cJet1PEcGhfxJWpCwnV763c9SX6ds
0EajW0Cggs2KWdhciAdaw8w5srfMgAutQTixhJMz2S+rl82twFUp/3yvPmpEwpVm
six1BDPUUL+VvCPa+9RttKoPipPDrOaOBOF7099tqXItSmpsOehIq4gFIx/phDI/
PltrL2Vb9cLYH8E8HVASAtjaLXsYjs09kqIbYWsq/GCKYycKtjjdZzUmE+kvWIga
rA2zFAMa8XaK9DGM66Kaq/oi7tHSYdzGYJgHlK0lZNRwOjncoeZd1unscATzxfuM
CmlftsCqOjWItntf5kkjNnhgKZQBacuyJ6A8HoTNDDAFCF/vMKwnx0brbsr2BAcv
gCz+klL0V/n2twzmc+K/OdNZ7x8xwtyW4Q/BbtB2DtLo0nxfWX75kfkCyOR9A9Qz
GdkdJaLALoX1f8+rTErDaWIBC/bIqdv/t10FaCFMd+mREekXplIdpF6krEtMP3mx
pcMNPy5HFh27IZbOFCcJHdSI/Mt45AdkdRwZqaRdEtrGLFUrPmW/UaJAofDXcfmt
SiNSJY4Kd9p3dsJoF6OZNR6Bi4uiCRTgX3JYVqYRbBynz/WkJ5J1SMu37KX4Yncg
V3jHnFD5dgoJXNzPy3CcbX6Yh3ja+rlBGykzuIkYaM9J/65acj9SfXBy28jcMezA
K3MwBEnsVI4OqdoKVv0R0NQ529oINvPIMQgoPShhX7SQTOuiNlt5EJ4NYmJEQY9i
hmhFHWUxVsgggyu2Njstf92Bc/AFmW6bkpkCMRVNnW+w+YutvaKoDJ5iPve6mmrH
gywtLxS5AvaD8oUxMUDZ1+ugRoU2d7vYJW3UENboxcQuxxvijF631fWKHYtXc3R3
wd3prvbel0Xqlb2kprKucvjhmFcx5g5EQAVQnVAt9dN0F75AFT3LlDmcykPEqBoc
rImcs+/44v0g/xfou5jLqPdOyMJxwSOele+rhJGB6+Z7c8+sIYe9ol+pHL0GE5UP
d6I4TJx4EF583pEXq8mjSR5HzFUeOixvqzfAK3+el+cDm5d71NXrVpJwsF9bMiGI
WHF4c5mUysCY6Jx54fJIVn4Me8gnBC7f0FwwYVZsSlEZspNhbraiFTp1kO8CBwt2
XxcgSdkMgb+bzOHMRJxto6nM6aT+0yFbbBadn3lYGeBWw7zlpUT26mf+WaIUQg+N
PX99ql6FXoXyX6AHW8+2pIe/fHsV8ueJedTy7Orj3ahnHMyFNmLms2vtMoNxzpAP
sqqbSvRVAXnuq675/SlpJ8YJQdUYYb/F976ajMgehbkAImrqnk0OJ3c/SGmZnzJw
lVOMe3q2g1C/5AbHOoYH6/IO0Z/Od5O6NiN1FewJXacJGfSyuMgOLx8CotnpHNB+
0ARCA0LquNscNcUUJmsoYpKc65nsRR4jFliY0oF72wNA4AARuEzuqbLiJvWc/W7+
OEzW12g5e0N7t9wHiT4f6bi0HsXibAMg9gHiUAT7bcSYzI85gNugyCHBCRmkCOkz
NQF+DqejeGdLJOsolBNbbxBZVKD12PFq9znYi5TUid+JwVgS8OvslFkSMO2XyRWW
LG8KnYqFia5YZqDLaKJCBYGP200cynjXhao63u0woqtfvaJhp8PoQpGA1Drb/47n
28UXxQH2WAQHUM/NKX0OJIK38Mr9WCx6voL0KTQLxbs6sq7nm6NoqEMTTBL6qKW6
aXfLZ31CFTpXvwMzt6ju+ig+dziWB78wROKpDnwawmVjSie+b1WtP5a0upJqnhqN
CIASrOtsDpL5STg0hgPrXftUJvdzLd4MkUrc3H9CwaOJ/5fp7/EzBlAP+99Ktcry
SeeKYwmiwrulX7tuC+EqgL2O6gAJLxEpaBrDVZdGWgsfHSX72iVqSFXxvpJwcxFi
X2Gd0cCqYFiyl/9gUgLePLSDrR0BvfyhWE0N/eXBMRcKp4tlpQsfnTlOJpmFFPce
vDcEzed2xXrjKkiXjK3B9yRNhkTNVJO1YV9uSw08dxsfKQ1TMAIGIkKsDbD6+e9v
Z6KUFsZdo6ynKJ+MYv3GQ7CqNe3+KqzxuOvOojRswRee77+3kBc5JOGBdycf8nr+
GY8assQ5s05EjtOkP2qw6mfo+0vl+bWdkgMmfbNU+b7OWUeeQ4lC/50Awxr6Wokm
CqfX0vWBVJsuelEwMIbD/RJBD3mPKIVa86Yi1IxT+COLu2e+C7387ApoLu/aqx7p
dzrrkXrUWxB7C1DI2yMIoeDZ9OU7by614O1jm5lMjCv0fMpVplkTRy3+q1TS3FKj
kWv3qe4nfWQsOwu23OXKUgCiV7TwKJh+CO94QRcgEYGD9nls/vqeI/zZZuhYpcUY
OImsZzSmvu5DrOURXBwKeBLbRrthOeCiEPZoFXtcOJT6/zDRuhj+NlVOoeydv6yZ
zH4pZ+wrIpZGS0evDWdnDlv2lUAIOWRNd9IhmRrYunW8KNgVvlKg7upRLEZzLlr9
M/05M6SQBEdIPD70fs+iWzfrmIB4qVt909W5lnXZyzFUGA/v1yDjah+NU2XsjYo2
K2MptZSMx5ahm5p1oImbO8PQeboJfG7YqxaX3tBZ1tBeV3hi+ZvQSd4EiHbUEKMh
Vnn5tl7tcdmM+oUT/tM81EdStnZVK9Iu06/JDQotssN1GUiHz9EQqFscKm3cKWYS
Yr7PTlheEmAqg++jLmU/FuS4flI6OxUmVvuvgLWvFZ9rf8pXUeSj1FgoeEki0Jg/
EI7u7cLRjLGhYDW7OBb5fygfBvZGwB0FaiF11NeEIOwTmHDLF/lYkGFaKJn8FJoo
hlLDWHhWPmbzDewjm2/bMSJte+IiqvoV5RGT9L35x82prNWrG9Cbc3KXMBX0UQwk
t7hNREfR8AvGeyo1U5OZ8eZCQGBalGdL3Q+oFUJkZ7i39GsByqQ5kwgkHGy8wGqR
nBP83cOwr7uPjYLrcBdrx3pDAFkFzXbvMtC4OdraQxKmMROE8loGTqJyJFqpMSIm
3WujiQaphiZTnY7HP26dNbHomULGVGm/pgkbDXu2CiatGVGzN60jh5v2hKNqO6B8
kVvM+nfOdPFok+P7q2ijb4xiXPNyM5s4hMWNB7NcAmfwrAqunfPENU5glSn3IoHx
dq3K8c4AbtuALlLvanMdh122DyY7ZStMQgVFONpq45DEK7oa2KoGhDorpma/ozIv
BmEhmc0Y33FwIUYGJv9NDPxHuoR5YIg032WurbV5TuFMJT18IDlOPWJyH9wA0jZu
A8DoIHEZmgieFmA63GWR80ps2+fQtkk0p5kfWEswlNJylaBU5NGf75FAEgPrD629
zlskxTSr6KaTxsmrAh+Wmf/V6fDDqzgFi6cSEbMvdAJ/uK9IGCA00elPntA4WgR6
ioa3bDQGKfRfOpjKlfthSpD8b6PFahyy+u2wYDdk81zVSoLbJyHf97GSK8u9oRzq
+KPBdePGQVH4sTj9xeMBdPV0kW/1RCY5FlEdiz5XuiRkqIne7Jzb6VCh2D2hzJ2a
TEPtCHCXiWx3/wthOHXWTgU1bxkfaEWdj4CPkrDLGpCwExkC/D/Q1fSEsq4HuSq7
dHiYphvRe7Q0M61Ug44lmDbSzUeX4nxmcl1a+m7YkwiFM1GLkQvjdXs83+Jd1ITx
qkfl2rHJR519Ti97+Or2UMbGIyJ3gNzhXfh8kxBKmk/9cACQ96ktTEtduWe2zHOT
Qacytym9huZbzjjgRJraOy7IoBnCQ6gH1ANa4f8++Z7jsOcIBhEl2pSgPaofTY/g
TPjWmSRsPgrkm5n00mdi2+ChtkQgwkhyMJBtB3Ic1pp8bPCyO27DvpxLCdwOEKJD
r2DVM0xa83t1Dyg+MAqbYEPus0TC+pBHPwqheHstvG47ApBaVg+Ax1U7HcN19br1
6VEc8Ukag/C14miYEnMVMMNy9/iNJ2k0FSYyYGWf+bmX/6k2GeMhyqxrVL2z10Qb
9lDOX6Mqr7FAr2kxmI9NowL9syLDbKZmPdH8QzlhFpey0VsBq7WQnen+1tPs1a9M
r5hPCWUa40SB1o5n7c7/Z2YZsbINxeM5Z5RhYG2NaIpWUvaGSfKtTjuvkCFEXK08
kZMBkBLl3AJ4J+Po8XHX7n1Dfg8ysQ0GNqXudzgUqnwAOARZ/63YMf+tWFoKXeYI
L1WZZOTdWq/u7SEszHvzJ25kgZTdxFxfrLIieopXdERUNSFqJrzntnrPDF6Esq+Y
Ms2HnGZc8wI9zta2At1g1Ctp3MVeJBYo2aB4vfI6qQzgY5bgS1BcQTTPkcqoHokW
82tX50qY/JDt4hqwCbABrmpGiMrxlZvJYaPArmlwCsJ/0qonlIdhPi3ir9Ocf+3i
wrBH1/sxvdcgPPwZPeozdAQaX/hkzOsqBDyIP/Q5nskmzsr8lZ1HErZkQmr23R2s
oON2ODBDW/2mihLbB8kmFSSbWZ1mytr19B21JHaBsLyIsYFx5AUF+UEoLhtqlp1z
5gzUtEfsqra1TaMvZbv7mFd9BzDJYvprW/M3o3A7s1JbOpnUkaTpeG8AZQWgB/Ct
2Xuo73WAHtM8VomJP4tEfMZVsJWeiEgoeOUGlA9Fiko988YbI62RXCqdFH7BLVVV
WdDripuktaGaPSpLGbsfuC0EtxxdTXfbmelnltEweXHIty9E1E90UNyxFzGvX/FV
xD6coKvY1oKP/8LvRysxrTu4IgK4hnTyq0sSsC3o6I2ArPuFOxs7KJVx/rZOQ0xw
kTq//UtOY259yfLoCw/OfwXTiDc2eNYYEOc27akL9JJoEzZZWlOqJE1cvmwiJDH1
ctNZykwnLi7PkJti8cAl7mqhxYFADGjHUTmFQnYo4eTgRggxnMT8WnQ5alUxij6p
MXw+m1qE2sSPoXq1dwagZHe8kDVwVL+8Ex5I3SpoLWv1+NGM6pTasbGNgcv53dJM
BHfgqDvedphOn+D5KTaLQ7UcAfY6szFXWMDtf+pmTAr38lHvEAvqwhv6h7DCCFsq
3cdeCMyqaoYriyzl1j+0RnTU+RJHQIf6z46eoU8TOHqsC0QZu6mYAbCWS5mRkySg
EIU8XktfVO+xdgxX6ajQ+eqBloCxx0OL13oz6L01p3OelUv1/u0egSA0Co/4cwXB
+bWYhzxhTOL/fm39WrWg1C3HdP2BJlXg3LqohGnNuH8vXCTRu53Ntq+p3WaORG6N
eISchYbVPk12kxsyo5F0XxtBSae7kO3IA3TkZ9uePHFKxR/1ABSCB9+ZQlaVyhsb
d9NBVWaYszFXJfQjAmuVLeuXFQvRINUdwA27kkfx05m76XtiXucYCpZLDf4oEyAK
TYD7hQXHxIVkA4Ir2IDN8W0qh+hnxCEjCZFKM2/hVS2hEDJaHPZdpxfZ4/RnFhs3
2VvqlbyrzGhbAEcqWEhAzuivtAH56X+HsAYldiaIaaBa4xHRn8XDRykeOWm/qjG8
JZKXmbvt4TQcP/gA2AgVW8MvkUyvSUIzXNGuRWmCTyhtI/TuoqfFrDRg9skJsc7X
quFJwYUQtlgeXOL0vKErfaIH1q98BjVY92p6DllgrSQl3LrtGip8R4oqbgEOPblr
jFrs0APvHG0pFhTcijfr4quyORoNmzStmbFJ0L5JHliZboBKOT18AyT+d+i4Tua0
MSPHNkiJ67uim2i7oZifNxDm8qWnrqnBwKeoZafmpuekFPECVNdiBqDEK6iDNtYY
udHpUYRidN6ybZpbBLp8RqXZD9KXVYz8y1WMIO9GnsiW/BecRRzCzhCBP3JTzZ32
FW1MCQ5HSF2HXxmMUriJgVVFbby8db+8OnbC4QBKYREU+eR27BEpCiVqiBBqIV07
7W1EPq8PEgP7RnFy70aSuwHxXxkSH6j9SszavIJwUQjPkX98z6D27wwc1X8kXaFz
d19IOaz2kCGtTF+0WGPDz4AEUIPfDWrJE717w182NGDTEt20158pzEe0yhtXeahy
zeH3CCdle7ppTnBUQB4aA71xOWcXu5eQtYEoE8rqIVY9G1l2GeFr8dE36nICMfai
o9s2qj6pEj3a/MhLXluBwCm1iXvejK0Xs/0sJ05J4V7EMETDl5D+1fYcuNQhJDp0
OadQV+nuU3rzWDKgnm2loDsOCNCpy39VAYG2a3SyTb234zLGmxArqANbVL8dND0b
o490E/KUiU/NWRrx+YLyR/qwrwa2sDlVp/XcNEbO40a1lHlCwFdUc8ur630ikjEb
g0U6zlPLLx4QUIRk2Rdn5sZ/iyvGgaixwI9eSb9p2OsPOChWjFuoCxjWfVEJJzYC
TOCSERhbgOJq2lmV0oyeKx6V8SdcLSiBqXY4cdr6X2QegjorZPB5IW4gD6zH6pZF
fc1kjqlSr4n9tTjZEPlF+Mwmxp3H15BZ/Dz3TKMRBUiALgGveNt5lrd7fGiXsIN/
hVREL+jJUP6HNp2cjMqH/gm8QV4ELy7vg7Hu7kpCo9L4pvAPELdV/GnXVulIzpl7
ZhVAY+btpqYDmFdE3jXURvoATX5nFt9ftFg2EpE/848vph+R8ZMsNuTWvnxhyUDP
CVQRUX3dZ15i+B/ruy2dtVWc9U69Fwe3uxSo1+mNEKlfpCeNh3fgJhZrfBHa9cOn
ZizD9nZZKRSkZYumDM1if3+Al6vlIAQlsTUhO21e/PPvPSElR/CFZlTK5NDGYGNj
oG5j68bbNPpQeVzmzpTJed5u8HdrQNnF10Sg+ZzwuDwh/OzaJRPbqIPCRFkTg5HF
9TUVhkM7HnJdyYLvtsqqa4F8yC/M/pBLC4gp3QsKhA4EVdVdMyd+Lqf80UYwEmwM
Tqz79r09YTXRmYPVmsQc8FpPV9CRJe/PsIRLZI993OCbCFnsaTAZjPAdsEjS3DGd
RIYDPZZhT54wr/ZNOxzGo3EdfO22+Pcg8mf7QzdYjEtlIemteTRMMTlUvTDG1euy
GLujNXRW33Hm4oGDmA3e7Tr3Nt9VT66aXgCNCxGc/B0QqIzSKdA1mG4K2yranr6O
Ef+NatUvSGaiaOgNStbAdeQSLiZEx5a3F1iYQJtIP4l939IkYpA9DuEjCG8qYd78
xff1jneF3RhygdzxpTRU3NxJKzttvbx4LN5krnukXK/78pHfBrgkipmfS6yFUA+S
ACw66yewJMTvZ6mntpsfignYnueT+k6hIJseY8s3cD3v2psEtdqaUs3AgRBgWzGM
55w4BA9BdXii2uG5z1Yy+bSvNnfsuz8GpLbhEk9Oo7HIUtYQidnGpwCFSAAnHHSq
JADxxxhAMbZsP4xvbqlpxurHK1/bvcvT0gFTCjbWt12KdLgFlIHdYGNHVvYKlRdm
QY3gxSvDJBC0QnDNmZlgBWskXTO9KoD77azxzjYGHeWFn50Xj/bqa9g9BDxEEGkD
m8eYiYPqMr6iAt+yiYtfFR5W6x/uiv7arlLld29t1LvAc0ZzPQta4PW+Y0T06SJI
++jBbpog8kD5LKpdDvwb/4uLM0ZJK+YmE8f7tCh6Vem6r4bF/mldtn8HvcI6RMom
F+SKkFCioc4eZk3AuUcJjY4i2UEVkWz3RR7WrP1FZwdPz7f+aURbA+G5Kce25vHr
qlUWED3ydKZpTeUsWaW8vN3MnZJu/1EBU9fxmog4D/xnQpd1vXFVpmP0N7pj4t5c
xE8lykQcU8FbPOR45z4Jbp1eungOnFUpGIJ3Zub0fqxG/1AFMM8ZZoROPC0gEiVR
bVhO4POsqlJT0qG8sr/1yetpl2BJmQEIRGjGHvmqISftjC6L96I6qZxYLYDzF4IE
zxh77QVMVy8lOn6nAT6u5FkRjUo6FzWq2kr7yC4wte1j4xJSkG0H1en0btN7mjHU
QVibafxjQ52jLGIgPF6hIjBGM5fMBSGneDVIKCioi34Fhh/1/la7WVxhcZZ6bvl3
XYTvTbjCDjnc4iraEzjyjecVNnNoo/z7cVk2xOTyY247ycF5YCPcOOf3WGd2Xy6P
1LZpn4cs5BQsx1snwc879OCewfumbbXBFaikjmaTfAC7kMRpUcyvKaP7/XjB2TBE
PjIn8L2RDjW15Ng7ai/J1VZFSgKBNMXXz9rZ/Gv0Ze3OKuTm7F/uYWHR+i0ryx0r
zZkOFzH8lg4lTpsSFk4xrMUagCxCPrchV5H6rElY6HVRDiMXkQwwgjLq4i5XjTmC
tNhW8f7dqr5ALjVc1S6dUm5ZuZveqsV1RMOKVLFbWaWzL7PLbou0Q8vQF9gJN92h
3wACCNJFjYkXLOcIsmZI9YQhbsT24iIxIjOH6aIU5SKAaF4paNHYFt0qMtuz56Jy
u4NY5XWTh8Ibcbx12D2uS6WuBOd+YOFf3mJGfLaN+ZrH6o5hPL0PM/9KAP8eexYo
GtChoDp3/JK+rMKBcqETrxgy2vm1j60BJL2GxIXSAnDx9I+s2h0JFzVsprNI/exx
OJKfjtYrFgDwCFzAwUMpMOjkT2pj46Qr5SwxAIfMH9SCxvIyy67DF90/ft6XzLBL
zyjnnXNy2Mdq9pLGtkAiI+rBzS9odaRKYDfwPEpXXnW5YmyXE4qcpmskDxAwWinG
VT/OIaVd5Rv6HXsgEWQZbzbk2iXcARcnRxpMbWM6IrBwFHgHIDliVAYKqsgwQrwN
DjZ0VYx4rensoHkj+bkRBRcLjuXPA3EdaawL81qZLNTU5Z6jjNQVsuRF47qE/8Vh
4mpUq8icQ19SoiPJa6nsqKi18wQqhLjX1R9ipfkQ7yi/5gqRDwnD5jY2lrRoBn24
JlKLgCb5ux9OCCT3w1VE7eLISoHpt12dvrfOBE1iwdxRD2XznZXL9m0jEpJoXmSY
8dwnTS8qds9X9cs1kPR7zTRrkTw/n6DxQS1ru+oTuR9c0FrwsXJP7sZrZAJRIiwu
LGSDZ38UnmK0ZRGloYpsOCHJXwfULlzTY/DFy6l0GG6hANZwF6U4/WnJX0TTL2iR
h8W44Kq7R4EsKsLka5UmpXrI/vvJmH8h7m2cEQFdkfQPS7v9cuVzScvzlvCXyWAP
FV6FpywSVhUaFBW728MREbAGB37m7xcqM7BEoy+zcN0EYyrZg1PghCsyKsxdmRwV
jM1AJcnec5zhmDUkDu8eIr3nc0vTWFCJbHJ407COaljSjF+38kBVpSXY3xasuV1v
K98crW8TtexCxOg9DqSfobKOa2BgSTzxeHsiF3FO+GX9GIo7xIcyhNF/2spG7v91
fclm0lGb2GoJ5QkLKEpz80TD0Vzz64u7910D9VVgGn9amZ9hkTtNp1oxx/S4mGKy
T2lWGfgmdE4j0hZXv998T35zWisfap5vb5fvFpO8OJj34a8vddI8hBVHEmApb8GB
mfn5XgeQ0iszQ+5pS315lSpTcx9yu7ajDw21SdXixRiCp3LB6dSAn6hNyXJ5YhqX
mMcYTt/alRbnkcn+swbF/D7Pe4wU+IVyF6GwAqHbWZXfMyNf/OJtKzIIyvwhJ4IN
5Ydr87+bsj+Cl31O9yMqwta4n0mHSDcJa0Gisq54oxAK2y7Q3u+cVPb7h+RWeGhy
kpnnxEgQMpD/vqcIlfiHGMm2HcQHWtpZBLZ/EiAROcj710PdR1bY6NCCj8XSNy29
am2Rl01QGSM8tpz7lFe4zdDYqxDP9VdmMGA6WA/RU0qdu4NkLY19BQ1VBfUU+ad3
J0VdJfJJOWP8XlDpn3P1vYj6q0lkAHrt9scGbutSXYcrxHeUf17+moYR9U1iodMp
yghszGRZHcRL4CBY1tiQG2xpFA+d8YbrAGsN8QubL4tdVdvdgFAJFFNH/NIfHBfK
KrEfJE5un3CU7pomCt4EQ68X+51dKhaet0A7VaByjas+7lueAf7Wk8qFf6Zp9eo3
bG4JYvKAo2sEYND0MmSmPKqi+cIsFPsvdE0HDlcWC9bRU/X2imsETwf9sp/tlMJP
O/wKu8WCW1sLOvbmdR0r40ADjHst0OyqJxJ7xBvcQM5rHs2F77Ym2ddr+yjb8NE4
rPTrToEhchBL3E+Ik824hb0/530rBZY9zuElsXHq9lkoq8FXyCO8QOgVGiX7tmfb
4VeYD8fhxoo4yhiNT6be6Xe/B+gEGjdQj2iHPpBdoWUl5m7Ttudjc5BWe41YK4dd
gujV3kQ8S5vTHST6uBpF0wQvxwjzPxIFrhdmJXnEdMg8K33OJfKR+qQF0PS5o0DE
CX3Cx5VHC/OMtcmXDwcyIUv8XPAvtzsiWLNLevCXay0PJYWQrACjmS6N6uUFCdI7
4mjped4o1DHTVcIv/Im95PuYN/r24c+AS4vOCTjbaOgkrGIcydIiDEG1SiKOv8D7
/ggPJ/byQKvWq7rO9tD5LmsTnjkozfDQK1E3+9kaPLTDXOdIwD//DaKMpMOXirPe
I37kKvJJJCmC2npSVVj8kFG+3l9tANOUyBDXiMdEHiQaGs2MWccnFws4APizZe1W
hqXqJaQqW33c285FoBHIRFUGyD/EF3sdky04cL9rEcQabZQi8903FcPR3tdXdU8i
WxIl976ogJrddvpuAsmDQlqa+BO5L9G+lcbpgI+Jm/1xzKDbS9H81IcRraQ+/NK5
S7hTBt5e6e42X86KKE9FQLJRKZN8JLN7+N1dqZKDivQ4xrxTbb5LQkmBzEON2dpM
gra5mRD/bbglhAlWdMC7J6vdg7YLZHJfFF1YvWIQggjJI9U8X0To2bQXHdh5CeXU
CkBAK0T5eq0tmZ62GNFMkIyQZPf2T9p8s97jZWJt+KcdzsJZGPJdTKDgNACb2vvb
a80I/K/p9AnuePEE4jbWo7kn5pVFxFDe/sG4QJL3VuM9yzbBwMhJdkh4D8/eJHpR
rllvnc6yDIwSaGiNV7FZYZ0NuKIuZ+cyYexKA0K3S2wF/DheTnmQ3mgHhqT2+VzW
ObSaEV9DsBqmwlJbDNXvX8XiotmYDIIbhGqtCiEQlw0kvGvBlFWAJIDjURiREp8V
6rukr97SWaNZosW/jojs2Op6jTnhVhkX4Wc83Mu6mOfeLimJoRIOLIfhnMLVbx8a
06FYKTDDG0NRZMvVEuN8jcb5BFClo7vSifYSY3bnTYabca+c7n9RcJDLzYi4R401
SCQ6juXJ9LtLGXajb78vA+L5r2LsOJaaHDec3Mab8H6M8nkcoiIrW0qtl+emHAcw
M9Rw8FLm24L2clA5yCs/WKMzrOOS8B7EzFgrjfhIo6l+SxtUwhw4kWm3Wa0VDNaz
8n+woaBzp8o6cg3L+cADAhHI4j91omUMfbU1jvJuhj50+4puRIhD+HhC0oCwNjpl
wbWOChtdHWal1RbbLOwrV71z5hkK4K573MynZj68EtZzJs17pIgm0CQjGkDBnPMc
VaGrekiv11HkvqPH+5dV65L3eZ7NNDBSzozWSOyjhcNuGZBJNIX01qSyhvOMt6q1
wVUYl7JS2Ql/z2V0KTvGnHKJHvfuCKeG2xPw8y9HNu6DOQQIQ9SM4/EdC+5OLWfh
ElFDTgrb7qDbOnJvBVpiOO4W3hLuHVAb5TwNmZJDW/kvX31pmvXcF9vqUsXifvo9
vOdsNK5bGW14t8H48pVsNHQRfnm5SirDbic0GtGB6iMZ0oNsAdf7VqFhgHBLDgZj
soyKm43Gar/oTw16H93Le0vBteQ7RMjVbL26zQoy1Tx16W2nlHX/9Z/CuTJ4tNA2
QNKQDDDw/FIlVRmHA7EbgLQ50PyAEa8QAXlyoZuhmCvruxQjoG7iey0ZrZABTTQt
pk43SFg9xbyEPiyWz8QNXa2VB/mSpi8ch7ikmYxHbxG8OP7//0zuO0ih7lp0yCHr
djLi+n9PSOfzHY8bZdEujN3p1YLOE042hQ+qW5p6RfcEEZGBQQ1i/UfUQtqjad4l
xQAqpZ7K2DiYbHFHdhu35jlMcBzcXKYK+BZysj/TSD3A2rm8DkfjK6oXa6cMheuu
7PUjShm+FNA0NAZgh3t1MmDEZath/DXBx+zKvAus+q6AtwsK1LUM0JbmNjydV0hr
/uwOZkt2TZs501O8dabuAMe0pyOT0G2Fi9+Mg/nUp2LYJq8YrgXe35wAdxOo+ZhK
HbGkyVu3VIHuCu3W8AMgtTEmZYpWq+HC54hBx0b/8Edc7yoGwF0g23KD6Km7bUFf
mCqL7+L4+cQ9O4uZI4c8Jp4q6xLpbLz9PaAUy8I7eRNOcIL2CLPvVqi7j+PghB8G
oezDuVlfLw8MV5LgtiB7rsBwNcVx33tc+uWibPXa5a0QD8kSF6YtQds2lSvk/+MS
PycDjtf1dZKMKyoKhH8mi4bBZBFMe7qIKMdbAdDInv/xK+xlKYqUT471gWKd18ca
Ul1Tf1nBHqyzyD8oiwhXUsfF6teLgZWUhJCnuVVjXPvSFnccMfqGIIN6YMOQ3WcS
r1/NLCeqGRNjWdJpk31hJfjQa48hkUd15KLZQBbUwqIq2R3IrHCKgTI+6RzfukMV
OPYwjGU+eST1a+KagHP2d1ejmrtHm7iYB6fFHw1RYyha4Mgsem785gM1P0egUT33
1Nizgi/DDxxM1UVYR7+A0y/sR7XJp9kKfCUpRHhx8ypCaTIJccjGeK8AVXvl9819
1nHKqUNqKDKStb/h1ed1MWlob74RrZzGd03ZT2MDrc7XubS0VoTKowN0MP3TmTNU
2iJYK5yR+OJpPmutq5V9lgwCo8dZYMK7Ij0YPt0s+S4ihjhqkpE4YcTcLSUIA3zo
MthwNpqwKhCULN/tkOhjltKHQxb5D1MlufS11GDHY1r2e66fyhYy3PdxR9TdA9nZ
xF5YTp/XX+SdbhYcPMCKRYCBMcvXuMBXGocCRSDizCEm8AH7FmzOD6xECaqfmGg4
keZHB19jMSwormbCCPwyFtKKwODhV5KpgQMh6MZN7wrnsI81MqBOyGE23YjzO7kW
nnQgNOX5IxR7X+S5yfNl6Cmw7chkA4HtpammZ2qTZbcM9HeRPYA5j5sDsSYyecaA
94pKGt0lzy9FGUPm7e7gz6tphrlha4xVWSJdyesDu37HGguZJUBM50UEpg50785h
AWcaNOxhyD4aMv8wPeuQtWDhuSTLRS1I6ijxsLOXohnXAHtmr9KbvvrqL2nVBDLB
3pgCc/YXKb3OOMk1JzUp5lLRIJIJjxRBtqsIvkeSkqGeIrQSajFbKsqi8vGcbhsT
Gg+UM5Rtt+akM0O06JTJxWR3lgVo8XnscULrXBjCJGJFW7WSx1xovUD9B3GG6OoE
kT7QgHdFBSsM0WN6JUL0K5BOsqkPKlS6iUvzaI9Hx162XksmJCAGIEjDOfx0SEmh
NuAM7HbC0fCpFsiaLA2cJ+DaVSHk4O633nqzs2qpApwP9CCZK89hEei5mxtDfnIe
Eb+/ypoIGDaQ9C+FY/HQ0Q1Jav2HrbZizxrnguBSP2aDT8WjjeFygxxTelu0HY5T
PKy3sAePQEaQEpKPJRl3Qd4fVQT741/Kvrz7zybURQXb0eoQ9y7brvJFnVrainTL
/wAEfDYFNJxw1X9UWEbZG15I+tHWE5Ib+aTYhAT1T8lUHUIeYUI5WRPyn1jjnWX/
63vWQ31zVXE5EmIW1wN0IDUlkTKvXWvHfpKygdwktlpaMvvMlHYHaybzIWioVN98
Va/nFQ2DQ5U6gdWUfUCjiHgqxd9YOhsYCX219z4kZ8BzzSBNvvCTn9T+jDLMMwfn
rAG0qYi1FlELtq+9wardNeZuqYZ4+qOO0Q2k8M0YvbaYxiwG6CdwFXCsQPp0Ec+w
JYjmosxn0fB4IwFYLt27+pAqhXeP3JVVPciy/tFg04/eVU66quuHeY/FsKFY7Kii
IE8OQovyV45rF+cdll7uDIq8wEmic5UP0nxfksGC4bebUIMuPhMOi+ZpogNSG9nj
uLXvnqfuq+ocL2ivb9haBfDg/D7Hzs3q1j/+AG1VbcRy6God2ulXnf9644MKHc2A
OxVDtaWx9KEMTWHf6X7hAjZkFyjzt/OZFm8a6R6xcv0VMB2Qll3oPA4rd3aDipPa
8S8ddCKkfNU0xqtZbXPe44ZDFbkSwmUeB+85fbFeqzQifPPFwSUFpTJ1h4J9XmCT
msMA4El3hmGGoZfWiaJHnwU0Kh6VqzZFceT9b/SAEKuKz2kMrRStdfDjvDFfF5bJ
XYOFPyh3gqta/ADEBeoa5IX3HfLptx8dy3aGdFLrVsfOMIDpqHXXdGgMYdKVgwH0
4915VtVxvnFaJ+O6SMstRUE8EcTcykffO0dIlcR1W55pSYQmY06h9VQBDGG+l+Dh
kOVUvPhRbVhC43QjA/qbY+4uJFU8mOiMB61lB+tWKBFEJxrDlokgv2axPxyCuAOx
gdvyRGrmOWfV4u2HrEV2hmGtI4zvP45tnWlyRSv7DMBQhLiyRoyPZoEXdAoBOBx1
MnwhWllPEWYgoLFuqRFKGhWtZcZ0i2s6WtY3S445UAzR5GwbZxEf7s5m+qmU+zoC
2HcxDFbQ9V1vDS3fsj2umKAZNfMwoMTj3cDadgcFv9PQPkjKZDx+5ZQE1BXR31ph
wh02OpSR3c+dlZ+DdQZWYkaZJWb21lltIxeUUd0Qigp5SZ14aRVLRU6YJ28Qy6YF
ztsM1yZDMEtZHyk67yJt1VadrcuSuKMfao9gnFk9qJvDcqMTWgn68UW2cQWpJ4Sv
53kun1iNkO7CknWEkyVq+ItzVAsHS7Ge4Gw6G6YRQW7rWlWXlI7EknJhEkGVNSQp
a7DIXbSpygk4vWZhbgPsXrHAjBL2bwfAXvdYbGdjfeWVn6TQESDG2jUdWeaa2iDz
u5HR2Nca0EZbnY/oR01unuNzMsGogLxU2NbtDf6UKqbcwqvR14+Qz34+JxCPAqPz
k2PSaylHtEKbMCT9V2cBxwSjXMQrLWl3WkggSndG8M4DjqVJSp3tWN5eSlxgpV2R
ZbJ1qLGQP6b3u38LJv+3XCTAIuPOrsgKZupGJRP8qxnRP6EEkcaMfLJsxln+alwr
9reF3ZS6sW/RcHAOFOvWEsWQZRtmQ1eTx5HEkQxHaI2JDHea50nX2nb0Qfe50DQS
hgv5kqzd6HkRFxqs5MuA5eqJJ5i4MMPZ7L8z+moCZa0lLbI1UztvjaDvkg2J0Hk1
s89Xyv2qntkhwN+xfCYunz+RIYqQHOwaAVBZfEmGzJTGEqJbWlaG72fsGmq/Jntf
JUrT+9wYn9iGbd04003B0UbLDqm5hhmEw47AaMTGeV98Kto+PTFnj52mFfZqomMR
8PfwjX/Xkp/Z59NX6iLy3N/aaOlDYYRixkfQ7sRZ+G2dAmBODkUok234oMZd1zDw
bEIrBqlmiiaEDjJHFFUBfUTWKNQ82s1qSDf/ev0GymQDuWNilwbhQfvFbBj4je0p
JgOAiE+4JDE3ztHKJaq2dg1dUAZpXyuUyLXEMTavnLj+HxXIQxC876R1OXKSBWI5
EiDLobur5L/TwkHQkoAluwJIMj8XfKabChPkDipuZzH48wfe6qX8lqnahJByBI0H
L3dK7wajSiwmgfid29PgGVUl4/Sdpq1Rwy7+peVemsRba7Y2gMitUsaXbFSxnb99
f4jnj3/mjQhqbf5aA8x2vt/VpogH6ntv8h16/XmcQfwCtRbajbfoGRyqA7oggMfg
GTmH98uQUQrnL646mTzlxybP2f1mZ2L62QNuLrQaV5wNdxjAWtCpNepnF+BmX0yX
L8a0SSrRi4qhIyp5PPq5Z31hPKasGFQJDZX0fAZMC27eKP4ffPsBCG5ov7Wwy0j+
+GLzGWRWuD4dbnk8Bo1jDXzx+heduT/BI2oiDMU4T0DX7SU3b8Xkb3XecEFpYMLl
26Bf693ODT4NMuE16lSqwZsIeIRGvQCbCMrRYiTpwfbqQFKkU8rZGu28B5YHqQwo
YRu4s2/BeI7w4SveZVNFM8dBEQrlgDSn3NABHaIDAqVf8nUNXRMkyP1+J27d08oL
hl+0jBicScWu9R3Ohush/glosjRpr3feKhWJOR5vcXhifcV795kDuih9VbUCLjUw
Dqm2/5txPgEB+JjcvuirX3yXfVlgtckGHeGSVdKRC7FACuJ+PWfzCxrJKzYdUdO3
jBOyuRnNjGlsNtCWcCTrUWzCHibbjf4RNncr0YtyjoMtGtugjfaf+tdBeUcPsIcb
tiXTX6RY32YTcwcqxiaxTHFzJuT2Up7ITSaEkZ9foNbwCCqpuPydBoYAl3vf43gE
F674ZwKFKbEJE+Pd/C+vCPr6TmlLSPSu/NgRL3GQf10htOitYLla+9OE8B6/lnsw
MjVFJ3jaLLtjBhA9to3cDSwEJwTe3JNswZ0Y/YjCSlB2X5JMxw1jysqFLYEorY+y
RA6v1VCBR+WSDtRWSvsPIoBwA9EJh4hyUNA8LPyCS4iFpckrrj7Z4Coy11BPJ9v8
w4nNlLPUHEWjNwGZ2VBVuavT8F/SEyvxj6RdGMkSk5w7uEdnRATeqcZ4JRds5RB1
Kyy2oDqdKZ4ZD1YGXV/LoGwUTWYn7gHRHsj5RZxBMBvN/qYOndEDakYobCkhxTix
A6M9bIqaXdihTACGZRKUyppeNIZf7SObMezFtK+lwNr15iU4wr7vQyVIo4x3myY2
CsU6OM9wRzWDl/1yTL0Bn8UrgEQX9uz8TqKZmMgyzQmlCj/IJPIHyYQSmBIV58CW
bB0p9pKJhsys+qkQ2u2FPawwl2WQlXhh2Kwr7S7F0VFPCgRA4o2JqTC0DhgvXQ+m
7zmCi8NvJsORiaio8UmKNXMu4CUMUS5d76NLEURmB+nmJHQ1FDClFjNXxbsi9DBt
ZKnB7DBgbdtMLFycTOcapcxKQNQ0T5KW8QBx3APoCpa/SVL09aB7qLNrT5C8Oy5o
IFQOoYhgOptK6h08irNKDdp/uCpnXqHKS3LRgmOjQfxNLoz5w+Yaf2oAmcgH3I+e
6bVYu6F2nPcNsTk9kb5Xdgcw3NXVn2IOpW3UTcHsL6zGuacM9sD0lVu/gNlgM+O4
b62Kw1W2qRLEQy7mkIe8yAv2oFE4QIFtVMC4VTUT+vk29L1U/vuaORkiFaGiyWk2
dB7U/Lv9asRRF46wMt+FXv59W6X595HTiq8CSttqhwChRvrFHBiM/4NLLasSNicm
ScyMhdN/wtVXieBlbebmScInnxv9irhZKG1iD0Axd3mT1Jd7EWN89wi4gYRbhWJ2
3Oj7cg9B8tyq31zVpmu9aUgUAZChMWnhewf1RXblP3f9JaExPfgk6TcSu22I1JZZ
kY+Ox16g9pbWnBC03U25VOqSq4RKZFY7MoVgChhbnKTu509/qNF2yAaxH0PzyngJ
hymxznGesnZUNnYsLNqIFVxjcPXTjWFoQt8MtHjFotv/gWgwk2uL8MLu/epuGGFB
f/RBZ1tJYE/ojR79QLK6Q9T/zTve/3/ma5POaXQ93D+4rRe7hkxcwhpg0thucoxf
PoBQRBb3aTjQvT2JE6Rlio4vmK7OKrYNbn8W5KXlMQLRH6qYPAN2xHYZ8Gxyii+x
8JSxxcaQGoyqY6w2zpEWVVtxSKmuDO7CqUvnePNydShlG4pbC38S+VFLpXDClffn
qhdjVkeycDGUZhv4+p5xmPKD2Q05PiDxSyWPEhczEHUhS1MTwDWM2QTIYt0y4i3Z
Dte7ksEm7no36NXDuApVjZuOdTAt1ZnceSCEA/wD8M93KsrcMUHBgJMKiXuT6rEj
aIKrqhy2YSlJ1x+DlTN/WiRGKG9ma7jOtMQQ2aXMnb5NiKiWd6iM8ki+de0v7vGo
sDqiGUSCBWRxKBp+3vsaaplFOqhcqHoEc09dWcwcI/MDhF4o+bfkubZiv2Jfc/Ms
WzTdb9GnYOI6e2rQUazivmR6XvhW7llBNpwSK5rf9mthS7gZJVnaAekGAqkygFYp
+058QfF3c9OopajDM73y30hlpBhf8JnYDVrp0AsON8bI/uE3GnNxQvLjslAn8h9a
cpYKBqJK9me20G84XWvDCwbne1lhc3OyBogp/FcpfKoeBagWTWe4Fet6aTNR8BcR
6fzeWloYkN9iEWLOsWfDCpGcubw99W7unfCLdFdBBZFGCvxJ3cxcluYkJz58WxGe
l24q/bl/uSpOxhJsDOQtooiUsD69/+XVi7NpCSq3dwrn58bOdsVkETfWOoTzBUHx
2bKgywrzd9/ymTXaekUeUTls3uGLcSSJJhIMeL2ofbsNZ5sCvq039apiwi3QRpfq
Z1goaKbCc0G66FotgJkvhcTDJQ+8mu8IMlExqC9w1+s5gsVgHv3YBsoW+ZjG8Zod
Ow/fdfdffMvDbzspstwQKMmrjaokGSZO19RfflBAqn4yApN/306oT6rYUFlP7z58
BEXs2CqCTgrIV2E08UqDIJCEXXvy7RfH75IR+ZyYmaBxkiKmZCGZ9b3evbRubp6D
jvDpnsJubr+7j58RS4GQCmMRGLHArTIjxI/+nIYCfFWlZVpFE3BH6MKUJtAExMu4
dPfxmWGevT8H6kcEef1SRrUEFbocdAtfizhQX89El62RBsQ63WWvu8tmcITESAEj
S1ak4PPxceXEKG9BAmB3bJ3M/NZ0DhJ/gVQRoXK4ExSnK1MjZPYrChE14uiLcwEU
eCqJpLsg+Et07ayEe+F+08jUNVby0CeT3L2mb8HMfoFYV9jNlE+b/9UNnRSxjGai
p7kWHLd2nJiobj98VPRqc5z+8tL4MTxhDN5J4HS6gJiCXVolR3et6JwkiXJSBrJS
N1xQMDrHSLlRy9TrTPnA97U87fDThNwOgN+oCDdhI1pj/B1jqNuA9UvtDinvgdVi
sDvyIAnNq6PAKIAiEcLGeYYXAHalsP0lmOLQXdDByd/vbiigenUs8K4atSyauAMA
1VKybDNR4OQXN+C7i8/2zE96UdfDtMLB07/+7Nnl0Iyocy3BD2K2/WKlgspczfKX
KOzzGeKasfZy/dLQ4xB7dKPFelkgmECcdo0Yw1PQRjD6QqEEW0rsFYmC4A7lplb/
3gYApGJqB6SsHA8exmRonhoCFbQTy6EprioBdt/+apckhue3rXGljayYpcuDBu0X
fGfxvHfULw69/lNnot/TgmXQfJamiaCeS8WwAyALMjcoG+MEMpmIkvdfARTvVHW2
JsgBgVVSfr8KwukxW5KMbXdbqsjuGgpztsLOhBs0A4a4WcVFUA3z6Td5j0Rhk99L
mdJy6tK04/WGndVujP+JHn8lusMB7NTVUSQeufvNq0bTKLDcif+cGErs3xFBBZ6O
z+VJ/DdUKHm3e/jeQqBJgQcSuHrdpDHMOJUiJact0RhYSBG9oS8rKeuGGSeWHaMZ
oGTqzIFB6YePm074oUbab/DoXpRFzA5e84DWXe49jYm6TYJk42fW6UiZqdRC7HgH
+1FIEOJYJ9xyzxoWWiDFFfbZ5t/FTUEu+LXeArdzSPD0ZYilf7Va3qULTvI7MK0f
8w7OGXplO7bOZ528bbYGjE9YjzRBtpQHG+cY1qKScB/TsFNiZvWZ2OpTXTDcK6uC
Rg9w/rZuv7WUh45bEHk/nJUmaneqEOQSTUil4Nsd6HoCH92U+BiT1HArWu77Kt4B
i+4q9fyJ6dTvRVF8vipMJpJvbONbzEkLs49br3nMl3n+kBJSzIuHysCfX51fyBj1
5hN6CaLbN4by6d1EehZfn6ufI7fy3+DuVHNbEd6gtekwZJFNAPxJIuT7vx2lheq7
JuNOxHMZCpkMkapxBFEP5TuHge0PbEfG1/pmLR6bJOnp0BAcTHAQf5YCiJXJnV01
vAP64/xpWcHMAhaSvibo2EZtbjQq98onUM3YABhE7Flu+TwTT3YnBTL9sLq+IAT3
Ypzk6/++Wl3AvOeaiIuWhpTAo8ZL9qmiJUq6uNcHCQDvMdH0HeWG0oji3kyJGJmr
GR1TX8n7YJUyU4V9HlMlm6o583BHt8f3ogrgjuhFcB29FpaOmb3KYqzK1nOCZFI+
YC/4I3DcCFeP9fzfAIepKCypdfT0LN6uduOhmnfduW6NNr0iExUWo5kS15oFy8qo
NZEX1txtbcn6X3KixirZJ0o0lXsE8FRJE/Rak4a7SYkucq8+4vP3TLIlMFkiyRw+
P5N9pjQEDRBZqJnDmOY03wKS37TmkUg6P5Ul3Z1eS0tYX0FhpX02QTWEZ1Oe0SMS
TK0E6Byd4FMpvROSfSzCWnX8MGpiXTvpJCZCf1AbwKfwS0f4guA1eg0IzunEP+kf
8St4bR8bjr21/u59IG5Pu5X0dwOetThX14NhTEOS9wm5awGT2A4Pc2B1FcSuLyBc
7S+YVSAh9dzPPXTigKH+DMlIuvoHsb2ysMNm3vgEQEAej6ocsS2syuSaa+7t6Ngd
Zl7rWiMQ36AXYX3riRrTkmu6RGNuIOQjC1EFnmlFzOF6fn7u7Qhi6P/FrhCiuih/
0TIPokwN7W5NH+AR9NsxYWL47BwqEW1czaeLhO1LhVMsl5qo1cT+wCa4+twqXCna
zjknSHs4x8Q1eQ7Hi/T3pu6IygCqiEx8E70r3KiMQuR//skdAHBKahDGrpXhY2Tn
nxssMeI7aWpM4KEMsJ3JFgoIk8aWWtLy+UwHJRt4Dr5R8Mu+H/1BO0Bnd+YI684v
DrSLh5PYPwXyeuEaPdkTH2fwNjJ4UDD+1SA6ZuyAw/c17E4bx0epEeQ/UZsAzIk4
QOc2nCmZWu0KdgPqTILPpofNV5I4NpOtIfpc9UYfS4QfS6ijjn2UCKtHOqx1uGab
Ki40JD9kJYkp2QIurc18Oo5u031HdA5moQYY1CdsHWLTGSOVAne7BpXvyD+B6Fr3
0Aq3zeH0ASY3BQqf+h+lctG5jI40v4/my2NS4l1U9s3N0zd+w+LxSu0/RmLqffS+
ZNUABg/hm9TtikMV/4H/bfo3JmXRhn7VupUOq1IHYPa8uJpiDLPQAve6uraZeUGx
dx1gj3nCsGThyQkzfufyGwsooyfBrf7CdRAMrUM7xsBBcRafoSRU+8Tuzqqkoupg
wrAox3qnX8mbE7/8djwhuwHe88TfsQVGGfyeH99ara6F5BQVgb5nQD71evmOYJFE
bPy8rIGXTiRyIz6x4gw9ok8LLbjcaEZsGJYXWuSZqJwFrvQ2v49iFxo6+ZBxBdMv
0dJcOQbDmY5G3Li9PEnPZ0yXos9tbDrwKOwPBHjq44htzNXvXAjPS/2lKg9InPFL
UhCrR66+/w3jQy8U6CTYxe7IJ9qXuhk61GRvHf6BaSf/MqohRN6aCQCe0ytPTOD3
ukVexAgDDuHfr65B7K9t3ULU7pV7XVHr/bZ6u5PUlOlwxRTwkyLjDvJmFy7IgGDm
uPqGdmefCg2LLk+j8VafcBwrZR9eKKPbiHZLBDxfOafvS1Xt0R9PuCoEqSwFCRmM
RCUtzmqm1eiLe/NlS6+fxA8Avr4nq1M0fsPyRurSa9cgXi5pkki9Jak7UegBjFnh
+IPEEwelQIxFe6QfLrocJfGUOHafUlMumEDEPcp8Ycdg3xfpm7ePmsMe7s5YOZ1E
+8rSODCPZ0KJmjGx+exo38aihsYefAIYy4Ixrm19WXdZGT3YdMhF36V6W6kTivKe
hr9qyzzwPKIpaOeYViN7wUyIAX6GqgvpdrBFU5gLaY3I+2Luq3pV0U57wa8XvlfT
TxEAmAWTUbTjU3buHRrKO0VFYKqyl4WWaN007E/xwWq5WBe194eoX69/9+ErpF2v
9+HFll22UE7cksV2+KXqWDInwyms6/alESsSImppaLcVDdpopidHtstjNHCdlVfh
h+WdsFBFo8qgg3JzfquNPGULzVGd5AazFvd1RaoOr1BW9LL3PNi/eGtWlinhnYiw
Mx99kJOE9JKbn1Y9ylRWk5Xp5dWZi+7xTuHkuIT6wXwvxRhBI4bX+UCaCemPf+hk
+6xGAVtkjxM3WTnOreEzASSu92Nhlx6BYKYvQ3O2jozYdB2tLWSG++lN9U61/giK
jaWcm22qosQ7IiWMhsnYOCdggTB6I/9n1xixsk3ntNQ+HfjhWGyHB4VSANXu1f16
nwEBmtM8kfGgr9m3ZCprX6SjQnnb863JDZv0coGXpwShFMAZNYvfXVFJuta+EPbp
S48PA6Cg/uf27uCBjxXbaiZkKpVzbxWtlZJh+E5Yn9a35z4hmX9z+IZ9lR+TSalE
VlMXx5A5D1pH9da9wWlIyWbjYH07S2Y/Q5P0CXrVwh2ZJPhYfdfBbc3sHb7UHA9x
HnsriHUAOlwbwzpksD3gX77Ip83Dv2HsLx2Ne9o26JrI2LjulONWs8MoJ74VDpvF
oIHKD84v5FVBxmy81UYM6plh4k7FPoDL3zvj8B6+dJWfOIavqBmYFlSlyOizCY3v
Yeh4yDMHHh9qft2KCzGNPUkHNBlT9pKLA3K5isciAT1JyQ4IzUhrOHp8xshG//p8
I/ZrfishiBD6bK9CKV3L4elnnaYYF2bixKfHe4xJIclMpDdIztlTWdASi0ivhEuP
RoNKi7K7LrUQNKpRiwnAPpZ0OIO+dy3UZUKQJ3GnQaC1X33sxyk1kg+TWc68EZcG
myCkovh8mcAVui/V1dF6QKzo9Ten0USdzIFK0FgtJsRftxniYBiqfAiRK1dkKoC1
fuIQNqyPMByDealnF/ckzmSoYPZ1grESX1xdBAKn7nnBGLzP4XZbYIU7Ipo+t6jI
KQpqkUssJ0398+Ym4cntOoW6MgIHUNehCGYwBUxwnyxbygJQsrKMG/2CMKDIVoSy
2MoGWbyZUWrV0pflt9mShJ8Ao03aE/648g0il7uoRavtKfoEgUGFEtroeANV8LVv
q2bOhltMDYkXObtyXwKLVkor5goTx/sqJ/VQC/VyJObpOsosbxwTRdDlBynafii3
yPGXgGc0ws6m0XJw83twyNydCSRUyUynjUgfx1FyscJoboOA5qkOHk7WvGx/jasj
Y0ApES8xqQXc6QJOdZI8FA5g2GlCrtn7PNjw6sEr1XgTNOxnVYs1AqF518KMuzsh
8XZby715d9kdF+NvgIc7GsqaGwA2bmRj3qo0zOXDGU4+EOntxOYUAbkn23IsTlxA
6JKh0mpoe9yda3TDnCgm/UK0qHm2zBYqwnHTxoPTZrfLQcmKrHXfSfzGNZbVKpFY
ry68qq09jSuacuqk6OQaMpMe6URM/cjC7vyy/L/1tjTRLy2FTIdtrdDOhAkjjN6h
J2Bybz2qQ8wZ0UjE3TOe+eGrCkNsKfQJabnVuH7w48YH9/MJw9obPa7PW1PHUL8w
j0v8LHTzhe3ILAxQOeWhggmM1JsKrAM6kXp3Ri+dvknd6xmBVgov8046XG2N2FKJ
lo8UMbPwjEzoUNgoT2vDpR90M/aLvvaNScvJuUjfgagKgvzTsu/WkR5g30StE3Is
1Q44eQJLgyz+KwLALFWEsFpmCxMwLDFtuPRyZDlDNIoAtyOXCKJtzB6MAEieREkf
E9NBC9B0zEpJ8fQIoSH/E+73YHksG6B+Fk9FK4wTfPMKnJQ2ww5AWa3Di3SgMlZu
usLz4x5iZfRdgXDGyVNYLzxWGB1fn4xEQIlTyRWPYi96P3aD1sqXDe7V96UQfNfD
32DBjMCjTA+1L3tmitWo+TaYDk3d/VnZyJn53I/2SDc3RlMz/rB2Mja5ClGQFgee
d+P0BHcNIIGQhQdyqxkIM/XKAE/DDf6/4WdWesWcmrF9ayvbIxCzGFhl0XFpS8QV
dLwW3e9exY7nnTePuBkC0tjkhKagdnb2RYsUrSX/3HmrC24LxuFg9D1inDyJth4K
Ka2dISEiUZIJMczt6PSD6mRMyRq23b9qqTu0zKKc3OBrSBK7kBCjm2YZjMPD+sh1
ZIx3WegF8zGm2kDTqvXX4nxFQrjzbT3eXh9IT1hDjEdOeroV0MzAt2WokPxc2NCg
udAmfxD9HwaODIdGlFDZ/4P/kb44ZPAwO/ysrCF6ARTnjLIXYZXUFOuH5HuYt6Ur
f0W9foiA6qR+fdnwIaBcHc/wfX7ob1gUtEk2vK/FX0Hx7iIG5AdU3nrYkMIU5zDJ
YpEQYaQufNsFN3Yz76BWRAGvz6mfQh2Y/0pCt8hNJS2o8a6f3PtlE2jCmXEf3sV5
FaOxrNyfa4IT08NIKYMk+Gjn0yH24/IJrzif4U9HqLN28FIz+ifbMPvnHRcZdeUS
xexClO0YBBDOCs8fpiqZGIc/sNAFbyYR8QV5slhTTDay0RRM5b2a8kiUlC/dtx+t
1Cm5j5b4QAWlMuc5xyOzB5wmVqzJpHc6gYaGZh7xFlAqs8ZumAff2THUYqgbzFYb
NXp4aGlbzWZrZ/qy4GKM6QUvS/r4mVO7xGsDTClm/OTX41+MKiXSYSG5k67L14YE
DXry8aqG3qWqwWJrCv9DYo9dww2uXIbkWNXUs9navFNiHunnz1ta4gIKZn2iYbNH
6HfTFpzBJBRdSNlPUUW5AkhQpCdGwHpt14FT/Un6isNq+94B2JAzvJYereHR77X3
qvwJjTAFcpQq8pRnw1aHK7hSarQRazihMLiQZbV7+GnNN0/+tlsuGDEqEd4RcrrV
Nor6IIy7KE55CVp2rCsR0euUFBEit5k8Xcid2EaZuK/8Ge/bgaIeSCAlN8Yhe2Cu
5cd4du0cfAFIOa6geqdX48ymrYsjyDSAFpUfGuOtl9Jy6r9jwigk0gXFniqTCHxN
fvgEvLzpXkrTxRQ4uIp3E5MmkdCNntbzL3rigOyHaC/WKCNye66sWKRmi6Rv6acN
OEIPK6IMlgThBlsSHEx8hqdrvNMrBa/jUEt8VLNT5pzsqTbdb7OMBsU1rOgBstn3
jbqDqBTyJ9Wo9dW7fbzDWAcya1SM2v7c1ab8O3mK1/92krpuSlXIkrPmAJBuRdQz
B08UfghOeA7cgljx8t1oEii8hpHpTqqOSRcN1PWW/REu/EjRNSapQX/4nkfryK6x
0enAu685UauZFrSD01S2D0G3pvkRhobL6W6YAImjJMfHRLszfuoRMGfMiLXADlUM
dLf0w0s8sBpvepB81tBguTOS/PlrpXi9OH7vesObHm9ZJNJoE29P+CrznZtuofYx
zx56wNnTfKShw4y1HpRnDMQDttQiMqhNoCF+dF+5Ffj1ohPsyZzG+T2WLszIhIEa
S4QTLjh5Cjk+03kveHRqUgasSUqXT2AqQ9wYzy1AeIplX6vzXKdKEyF/OyJReRYr
VJwHBJRtp8X1aLcOlGMHPY+g4OvaL+ZRywJJnVrF0zD5VGhqtR6YhSuncFplnOEI
aa0EjoN+GLbvOV7BDfsYAFo2hk4FZI+XBGTrKyK85pYwNBBDk72PYV/e8AXh5H64
K5lREK11+pgHxID2BhjRIFOFQvirYPYG8xaIkDuAp7O65Xyq6yCPCXoQ4blXi+dl
3PV5gxkA0l/tWSXDGYSvzOAUkNDldNCxyL842HTLqMfkDN3cNjL+SJx/yYA9S/co
h+8QcSi0Po9/RRIzwe/+yNhZRe4arzbIdJRpVbSJceQI9rbd3nID+2b//abVOpU+
WMbd6o+hkhZggzWfdQgwWovNWtq7GQCJ0E0hNvmO3lUEXH33s+iiM/EwKmKVYtFg
lwnj/UGN4/PtP9ARh04L501IOhEShXSjO2YBuN8sZU+B0LcZnwK6sI1OSZZiTpWO
iEu1kK2lt9xmoyfJPL/LTRQDcYnnIDizE185xJIT2NvE4rQZC2UA4uT5HkGhwD73
Mg3O2KEzTqDSj7BXB1pVxq6fNDIDi3JJKkFF6by8uv2e7L3VUpb52IIMIhIsL0w2
DoVpxW2/rZc7kJX+Ms11HM17oebADbAny/wN3+0pBSfjvxa6oi+qrmwQOLZC8mdj
BK2Ar/4KVCnMpWfQEIVWn8JykOJQJZsjun2XejfWnMeCEY+RVqBzwhyL9V++4hTV
14CHfJ8MNhKwDY7jukEvj0+lviUcV9zEfCSR0vosPkV49s2XH5ADY4RzEvML0H1n
35pZaRahgFFLBT668Tp1wDp+gosY9Gehji9lTeh97N/7dWpLkItqO1GapB4Ee4ei
P23QqxksDXxs4E+idt9M7Fa8tgWjvMa5ekR4MrMBkrMDCYQmM2l5rpLY0k+IIiBG
RKnfRtkpuI4dZmM96GjA47yth81K41p/6n6b0otxB4GbZ3BSY0EPYn6oQ4wLSShd
Zpbmw9w8N19BScW1/6Hv3/YCuwP70cIqLntjW9mNSwpyvfbBaR75jcyKa7lYP7oB
moYj6B9V79Q4vnqB7S2CB6KicPCyIrIPE/e5OzWDpfIZCnPzxstr0V1h8KGjT5Yt
U4yk6tuVGCmSGvO4He9OpSk2iqJoiwu9hyQDrwWXV4gvvy/7BG3x+beuznLKdz+m
nnon6fFdWasRMxhOEl8epQUGFeTCP4cPolDykh82zWTNmqTBexeTX1zDaRl04F9y
LpiVjU6sTm8Ga6WZ1yACY4NEenYt+5g9B8BXvKHOuMDRbpjJl5ZdmzKenWLkgVyw
llK1isY9nqr2ye7bGjez1SBQOd/e23/0MXB2peZQ86St0B8TuZ/o19i7Qo97OTya
vMtH/KTqvbWJ+eV+cQJuEONe1uMDk1UQYIt04hVcYkTj5bbXH/MuZEIBMY0zYOaM
hY9VgcY3B8b/ee0r2bcJQwxrw/6gUrk1Yrz2mreOIJ6uRpqC48JBsoLJzzP3+gS/
DlRB1BeNtUbk7/aOSbtFnQezqHYfFoZPCwkt2fOf+vJ+uF/R1i8AxW0ev8qeeuLH
M501jMeJFtaPeOw3nw4rh5/rgk57N9EzzqAlhJYXY8kcOoRMFSvsR48OgeamwlSD
+zGLtIB6NV49o7KpraL9RFsYYMrXYXGugFWfr0NncjlKaOotwybe8QTQLkfc3JQ0
Ht0ECGL8yNJH5FEW9kj1p9MeQNx5GydumJHXeAh3r1ento5wVAxAI1xMIIDewly1
JqP+iPsYUpCgD9pGUPKsMTQELmeeKPu53XkHwYDOZMYGJpnPwiPgoC5Y05ccN9nl
dxp25lnXZGmaxpIyLVAwQ+6eS0kmTZqrxWi6KVTTRu/1B9SEBQoMRtt+skiff7gL
vPkg4scE5khuUdglbQ2fUTZVISsdTrMbGF54mzzSauS5gva5efQLonrY/OD8xOSo
ryLNcXvqUMtj1J8ss4VZ5T8QA+UU2yjyxoFF+3pbNBjTk5PgDmI3FSWaUfjIAWP6
qies9vJo8HLp4cO8CzLKojmOUhx1B/bRFvL+8CGX10Zk4Vwn1qqqoOLVqSUjbRDS
qvMpegB0SZ/RR+5oavRoG7LC2pBl3ZQn12fx66+a70KMEuKx8qU+1VDb9m8L1SfF
9Oo0gGkhw7EtD0bapiZnERCgQ27j8C5IE9gb9yI8vyCUSCaFFWoVQhOn/6D/A6SF
cq7fL+RKMDQRPNOE1cxjZzA+21pavzC34s3BwVfYLbpcuYNFehFcNfmhoqjOKJdW
XlMDcA94RohNRttVu5I3ScOxWQetMbpWIMqNyMC4ooWGQ2SfSthefJSQUWGVrjD/
ISeKPOajXDYv+he2aDXpTcosti+8WUQafk4qfDBxgi41bXC9eJatjKDUeb/H4rvQ
upOBEG1xhrINqlRZeQgS/s0JG14LemnAOavt7GnzLk+5wvfK+5TRtlTDlYUj1sC3
fcZnJVTBMc+SwfkkKIR5dkvtUWjMa5bhx9whnZgzhrlQuSunJ8tD8vV01ZXGQOEV
Cq5FSRVTp3hNqeSrd4zeVk1yM9bQJKEIBKZmX5+qQwt4bsz/QE2KH3RQOA95v3vl
HWpbuVB1qd05hFkJDxA45RcxovKfGu2mJ8rPWW770FOosnPdZWT10l9RAnrnsE2q
lhFz9YfeNFj9qcjv3dKDpTMwEiuCl9MPR9KpwyTYt8VmFo/EsDa6OvLbL/2ZOVvZ
X1QyELMCwWIZE+zDSg4TQ28rGfM5AnVuMCI1vN2+zQkFP3y606Z3h8rjXwDClia0
xxRc62IrCkTsB47R99oYOwcbf5+cf3U7IpbYT5+rn+s5SxE4htNuSkdRGXZqUh1V
jsplZ2Al38BqSjClE4gN3aCk3p+vFM1mBQYV6+s/hFA2Y6a3Bop4v0Ov8Mg2HrPw
OFfvSZSt66VvwsBrAEqkYMq7lW1IYw1WIbL08hhhkpfZ9WctLQmMlsYt68mdeEDl
HBJlo2+/6ssR5L6+1IJvKRmrB0en51AUwi8w6ErB2w6glwPD3uf+cJWwD4YWDfhN
Rl4sVvF+Om9OrSX6Pl8pej5pqS8OEi3o+7t+HM0ky7L4MbpqUzkuApJGDzwpjGoV
aJeWz8Lqo2z9j4qusIEXEKAx/OavKBNiDIq6x3xC7CgwuWja7CXWc0uA2y0YiZbG
fHmxetQAq4vCb8blBgjgi4X83ckA4A9cjnpNPFfjA7/c5aqBrxLHhMakkSH+9z8F
7JPqOP93GaBP4JJsjo05Wwrgs6OIgN4j2iB3OcjKiwdm4f4SLH0e7hOLvTQgdUoY
9FZVcZYh8aBTWMp3tInqRZ/QNn7ZR3VL9pY+x/kkMvLB660ZmXhrlvzpbVdd/LRQ
BmG9qeK1z+JGrMTj2TB0IpN0oWX403U9ofADuiZoh6pvUJHR5ykFn/9TBDd3IHyJ
Viza0C26yg3rQ+cXewfiQ35hoedrBaBMIsmyg2VpsViIwOfzq9m6VswXilNnbzVe
3PwUOmHYV/WCgb92o2lAbCsNLikTkVxiRSh6TvQbHuU5GEVEznog71mmbdcsP1ri
2ywIj5odC+A/awW5WStCc+VpwrZVvJVHnrqLJYSyq8QLcfl50aggEimhkn+uRSep
hiP8BmnKykmg9fbLsG144Jgn44YRis2XHQybSbAfpci072Em3q/0ix0VSh7i6wY+
JL2stHDEbEXzw6dA8ldoSD55rP3e21DwVlq9uikFCMkYrb3GpxKE9xWPhbsWlNr+
iAynS0LlOK7s0DJSuU8HSreKAoB2hNIn8f42yFY2u5qMZVGuiZIJD9xt5I6swGwV
RtzKUy3Lm8dfwI9ckEYhdl/vsg6b4I80Q8f+eym6kk7N4T3rCBPboVStt0bHL7aj
dYEFy92PcEamvIR5b1/qM5ZjG5F7P1ShoTAXSmDo+vMZDo+YsS95oqVuBd+QZtCX
a0BjvimnJaKlF4/70398HQaxOWS+VWtlh+jvTv6d5OEXsPIW+EoAUWdUosjfvh18
2NUdBMigZM2XMf2iQQQlPRv0KGZVxbxViQPn1c8HKqZLA9IkHpiMlTzDPsvOotHP
3H5hrSVAsswrSsazSdWy0T+5qbhLBWx2Ayi1Lm93isobzbHj9U3zdyRathD8qxHU
KXl6Azs4N4kMG4Ike/yESiACOsR/k4eZJzFMh4AvTdKUZMKTBFZI4LsV2Tk9mmaJ
B1P2FwnmxXhEMdYiPLT6u/QYmtfGZHhnSOY7C/UpMHI/E6DxUX+xg+rHLaALb+Z/
O/QbavXp8ViDkfTDEhvBkz47GRj+bfV6vNsWpzshGm+2o+7sS1dGAbs9YIknSTAt
XHJg65DegI5hZ+nTR2erG3vL5t79ABbZSxYHaHophABPCohBs0jESCxFgzEEz/P7
iFtYzngrUyV39zcmm/5e0YpAHnShtsK8n0mR6NEJLKKmKyYQsaLZav2HLoi1sEJ/
yIPPwlPAaoHvyyaC/KOY3uIKIfeplJAbUptSYDvSAlBv7JCN/DpIuiJtPIBHge3m
5iRzEz2paq80Sr8uavJNGAGmnrxmLNPVUBpj0q0YP75GNATJ2jj2/1QPs33i4+Wn
RDDd1O3Ie0+FD8YnLogzi49GBTmMd0qqG+3CB+X6KKqKy8IsueM+jIc6p0Pl7grX
Bfbdq1jWv8Do+rzdSttBfbUYs8GTYb0F/52O/7ncaDqv9NaGrxmDfPE5PFeJmAHe
tp9o/peNO4yGpuRu9A6Mid1+XWczsHlZinj0q1HEnDbFswXWyk3Ep8bundzdO/qV
JVrzPTImmx5XGHXiQ9rac4h0AETvA33tiZ4u/v/JSwIhy54m4Yfy3rXRDhJ4jAzK
ZTwn4Be+6haK5tq21KN8eMO+TaC3mrz3fjaCz+OIBMtFgK+dFI8eTw8AIT1n3jwf
AyGdvIpGBUXfadW2WXzggVJU1dlU9TFUboA1QYHfMSWKpqEt2Cmaqp9eRg/1ifXe
ytQve8/EtnzCMJlJ1CuuwApVyQ4t19XEgQQ5VcFHQ6ZotHoReiO8V3UKX86KG2EF
DRL70oJPXsgBi+ZfMy2o3JfcMMc1ACZHLMV6X3HaSO2NSh1+Vg563aA/jjptILGH
jCVcGSKZu2wrB9IDc231+1F9eKRR2suPc678wcZEK5logmB+gsF/2PnG/11/69S8
DFrWrq+fTkNi0AJl+bwaf5b8TaTtnegUe6I/2BABoa7ytUK7L/Vh6rX1up+2Imyl
xNxq4kZmdH3s1fQy/lPFn2wJTDdM5Oqo83afbQP22MygYSW7eZsRPykV9JXDPI0k
xRRnkQsE05hcK3lKSpYoBrSZCQWGY/w22C9bxeoX2zjbMxYkA/mUeBvMR9iK05+U
d6cEW4vrDC2SyT6MMIwZoGGQypW15q/h1yipI9ZjZCMjhJ/Ce6G/uIywa68FyQpX
wYRsi0hU+k5IdC7aeAmUkm2B+QjnLOXrtw+lgnUhmzR3gCvj3QYNp3KOoct2vXsi
HiwTQCjGLSWZXOWHX6Us8Y/E9bwSnC9se304ecXafDkVmq8ExsK7IP5DdRIrG4fu
3DbGMkeHWaajwqP44A/+vlPHaRgou9ma4MmknCf8MRTNMmjCMkxKqzAoaquvLMNx
9EsavjavVLwjPjgo4KdvuNt391aqKWlQsP1QntFgKVuemsbCbp9ercHbjLcQjq4H
Ben4wDRROR/MYCQjAjDlrO4X+F1ngdYB6OmCFxlbnkOEYSTboFYRDagfrxHqNjxm
JPkFx09DoeZLRMHBB+VJZR/ysUSH8UOQZGqE2VWPp4vMQa385iMMAqixZ3vaQ5VM
yvO3ZynjS4uHIMs+xrEJtaIUqAiQe9K9eFMjcajy9c2R0/Uqx9lSRlRXuJlqxWI4
aWcT/RgUbwf+x4AGjkWATCoPMmSaN10HRHYR8H2ywZ8iOnl52oGit/oXiIWUT+Q2
3egT4iRPwuyN1iXSStAm4kbzUKU0vHRPHz2X3M51MREAj1X6jM75Nw4dwArozmSH
PtW6uqVlMH4rLecNX1LlHDGMJV3g+DYANE1rs6gQRxngewbOBF7do980M7Uu6lgY
2ocUBuEQe9xcuuMtr5ukPZ1JJGf9E+rf2QUkQDB7QMwrts6PK7RRVDOtrykvxHCi
kZretn7re0SfDBGDbYj7/2grC/HV2J5memL9vVA07JewYaOSxVvPzsNg+hhKeQm3
+5IZpCZKGI5+OlRgoTziJvuO9oB479iHEDOFKcLYS80CXMRA4GFT7+ZIdvgQQQ3c
Ooj5IYcqr6jHM08Z8tQqMyI4GZzhRw4XrN1VGfwY+57raUWTmgzGF2uYDA5D7/3v
QKloyi4oi19GzEWopdRchSxx0EN52hgncPoUhChIPIBW9dHALqJaqXZt+ciScZun
yteDbfjAGadE6VbdyP5rucZ8ULIaBIjBY3J2PqtsmNlee2nbNndjxs5uNQSIAL1p
kkoePfLLhW1JpBoRL3DpJchAEvG7rFYhmipC9qcSP/vKf8nkaE2kvj6CWnOo+wwJ
B/D0J68nv1kVWYQD/Wo8eg9jqxdFUcgJ8+R9y34DkRnDJ78ZfKE+zv0gYzFyLjCx
Qv87UkiAu7OqyZRB6s4s607/deKiUBvNc4qWz3NTLycj/jJU2CR6au9BGUejhrPf
XjP3oKdLtBxpj51amXZJvDMzodlgLDioAQ0NO0HebTa39i7pCnrWaGhDDvAZ8h8c
Mw1qvgh4hrLLfvCds+Pby1pAdgJiaHO+q6RI/5VmZskA/SJbvu9cDckN8vOY0BSV
vms0/EBCoxW95I/4vGE+QSu+eqP89XFZ3hQDkHJtMbRvT0794xLAZIBOTpYOzsaN
AOQ25O0dVm6Vhy+Af+3dIk0NalPHSV3qXUy4aWPDWXQi1uYaNuh1Wr7sybXXvgw3
nKi6dycF/NQYL1TSr09ppfTcKF+0UUTf8EAI5BaGPUj54BxxvxRWvw+CzJbsdDfV
4sIwtNL4GjG16trm1/6KzAVLaKNt9zEpRk+8fcfBKfl1jjDG0RNCqrtR13YrTwGP
OJqa2wyGiBYeYGpTJ5WP4usjvVSQ4xs4WRr++d6YD4Phr58vCTtoGQ9LOcLka8Wk
779RFhrI9eaOA4qMd4h2Fx0Sxmtpa7yK33iuspz09Hku1J00DTQ7miqUM2Rh3MRh
g+F8Dm5+dWVzzcHWoPJjLHxk7DCGRSJQrTP9AK2tglBh9HCs/70OrkwB0h5wWkxT
HcGcfsoqIsMVMa04H72CaTdzpS9iKwTcj6iVZng4A6leDpF+12w3MTGp3XveD25G
NOHIQzbppqt8DL9rKK7k7yjgrKWk3b21Zl7Axd+rlRpXFKXlghVO5PV5p72pmKtB
sovqT7iTp2i3OXIV7SEJ+xlHfUj/mZem8Looty2kStqUVC+/Gk9M9ZHWxSlOBTUu
4KsG/Vd+U26yNKnxKj7yioLXLf1+eonx5E2jOsfOht6sT+algTjTrXw3Er1OaQwl
eoXsIahlF7Rnflb9CFbIbjwctX8nVfJzK8jgq0Nrk8jxStLiUwY5s/i4WzNmmYDG
82l4ib4b8R6Qf9F0KHXXpPM/lN6XDOQMA+2RJoSt+1mHScaC379DEOEE0mhQaICX
vE9J2FuGdmQF4XXZrpsepy49/vNwlOcDWWouY/sdvGtvsRZWH421FWhq5pPjz/Cx
e8+ahkvWlFIU5FLAj6w5KVaSYqI25A319bi5WYfp1N11IJnuA127nxfa1OZVmxRf
3hJMHWZKsAa44M2S7jp2rWyz3cptxoIQHNGFhVaE8R+ZYaaEsPJ8OtUT9eFX5JHN
AHgvjCBD4RRoVvRU9fxqRkshjI7fDeB9/ngR/Lawoxe3u80N1nPGfg41KcEvo0ry
BO0oGt8DumFQJWkW//BJxTkNEf/CvuheWAIkA3wThzUXGa4FMkCGFYrF6PnUHJ+E
l+kSeECE2Prgk9nBQW0Tg4R2lpcTa466tH5XfgaFG8e8DavpT6M5jYKMKgOel/HG
JShRfAA0prpASlUb7srYiTMlms6oCTWY1smzpy1uB9e9TVOYcBYsMLA+Q2xOmVEp
bxla9bIlMM4pVDKkF5hRF7U6FBpMF03RfmCkMJ24yAQofvDkGRLw+y+EnY8fWvon
rOlnngWJX/ZH/8fbM4EaJ3NzrarE+zgpaUM4FivsJiwA4xtP8Dxu7XBXNe/+c8el
2rMbNNmvr7Y+JBoP5TMM0SI7u1zTj14IpevKZkn5Ewg86fJAMv1HrGDQ8OQx4wj4
jnLFyK91yFoeb64IAAb+mAd83NwhiHGXkd9eu0QMgXaznrXEAnFO9GFcsiiTyqS8
ZRvc5KQhk4puxpymYVF1ljoTlQjx8+P9zJ7YCRps0xjjKrKOcGVX9/r+mX5t6PRH
UBt5GrHf6bp/uCfYnppRBmrbw63xM9eLfrOSGooB7vgrjeUfSLg6RPyeAyKnc+m+
hPJZAwtO1RnAKg1Iekr4QjohRqHMwDE6OFPgsN/fy+sKND6VkNIP1VK9S+6UJDHQ
9fTuaqh5rTMoB6fN5TrPKRvzQvnxcT+wfSVDquE4fcRpm5iwUpSzCB4ZumPanTVt
yA8B7R6eQ9LdHKQ/UBZq3egwpoPYOGWzVv7FlWyKfsUMHmSp3TaOb48mUv7v1QLo
tMwYsW7bVJwiHHA2OUhKZya/cGfid9IPiL05OG1KxIYHK3wc7BCcn7a4cVpPsXca
i2Bwgtn+f9yubyTBHt6F2ZZsNzepFbnvAx7wOpIoVGrTcGdEvM3d50urZPQ6yO97
ePds+fmBJuhjFzeAi1Ooz0VmnRF+yCEU3SYFJBOZcwO8O/eaBNJKmXVeqAWknHIL
bhThGR3NCc1oMoIOgVjlO6OQ4tJYfj7JWVCxlyEKPvNB0DHAcZJnL4ijVI2Nmaqn
PBFM8i3KoS6D3UjoM6dHfb0bsVSrADTEmolRfDTDst3vjRmErMVivXPq7a8Kh6h2
Nm9LpHmtbJf98vrUBlC5vDxWhCazxEQ1Fznuqvi2nia75b4D5klTcxp2JN1NwFXj
pi4IRV+pZjUXFWIgReYfwtLPGvFJnJjCR6ZmLoPba2difVtV09sCb/SDP3s4rP5n
+lLwVFSCkhhXkR4JArhNPdDMVEsJb0yWvVCosGG//Tl+w8ibhs3JkXbuz6wuGCw6
24H9NFctoPY0XROIZY7eOR8gAyBK9i1jLWURZW2649mOBQAa7Yj4SxxEbKcvdrFB
4DlkCAyRJpIETCuXqfJyRacTH0Q5TRpNoiuwsTzil0nubkNF9eQJ7xxP81O3gL88
P7qugUNT1BNg3SUm3DED50pXdvunX+0Eq0SDUhKDnalZe1j6+ybaDMlyRpBJkPlA
Zz/cMoVmEAXNAkuTIQHcegSM0mhLR15S1mU7PiCypV3rXSq5k8q+K1Zu2F0UkbYi
vjoi8t3OfSD4Dnygu86rswdrEDO/kWs0ABpKDZKXSnKdoXrVYK3DNkvTw7YO9Fr6
MCj2nEEYcTNnKcCXNTLGN9KOxMZkrKXjxh4/sUI88+KAn1jJj09+1a7OykaD1QrZ
ATl2KhnaJca4OotpiLbkQgguZqlCuFHxEHpk0/uVKBioAvIYh2Cx2cyx9aBog/S3
Swef9xW0OIMm495Uajck//xsZZxNbyYhYYS8z5GNpqYGNrkshWgrSm/yrRAyk1wf
RFAPUakiVkIIF8xTdWuWatqoxnI5elZwselJ85gLo9vXzIs+TbdKJGi2DgjYAqls
LEK5y7qYFYLE/ODSBYS+XEMkE+yDIXnIRZGis+T+aCd2ro+ToCCBpTHxU6oqofBW
MIxu7ofR9/pg/pmgo2zWxf9Yw4vhKh8DKW5oPIL3yU3yKzQXYzWSF0zeWdrevUtN
9q6nalYyAkxSxwIil3Nkfnkzpt1EDHYb4lSBcw2nqfwAiyL9Cbhxr+21EEXfh/0L
DKrvuumz1CxUc1rrYYgIHb9lIFWh4EdLtb2QI+gIH9HvuTZdMzgE/K/ALNcz+wUn
7ZSmRuzNmW92qVou5h75m8W21/X43+8hyk/hIlGg/iVxHqfey30e1RAuqT4vz4S8
/9OvX8QE3OFPuvspNdhdCUWlWI0QoIsovdhHCaaz8/KmC1m9KZg2XaoEH8Rcm7je
aonqhwFfSjN1MDrnkELbLDxHba8LCrc3ZlQrY81zZxcjGgI07/ZG4h109oCXvNtp
+3k8BTTAJl3fWU96iZW80T0O4rkM67tWPCctygS/bHnkEX/wsTLfH/21Zwxs8gbA
hphiH6rLAQ2nRZgapUpFkPwjQ6RA2/ko7IFcgIdozRFPqdoo25+LqocyuD+OE4Vv
kGTe+yWb1iXspdHWLzZ04ch9VUlox1IFcNuLosnsRgQcjQoZ8AtP0TJHLOSUVbnx
rwfBbY4ozMD+UUIBX5J4QxJ0Hk75BYJhmqRa8fjUfbeO/4YyL9SK8+ICZB5tafu8
ejMc4nK1D3+DDUkhrs78qZEtza4TeUMGRddHPS85yqnYD6DXwjzXDktO7DUXgY4J
SHy8GlipgJZYgXKDAts/yMLwryO68XWLM10z6s/GnNtZdk85ju5iUPZAZwUhBC/t
wBjAOTzjLY27LEMQ+dPtChRhbYQzJj23b+g32775b8U6CZUScFK5SND62elR/w00
lhNAczDVMLAx0F+qD41BBi9lJI2j4KFpFQ1cHPgPy6LTeFfx0UtkF2okzdQB9CqL
6wKPz9j/PtL2Mpo2EyuTsKsZUCbEqjBOBlG/C6DURWHRQThqHqLmyuxTeuTGNcKh
DEma6cRdWXZTRUgBCRycWhUd1dBpqXa9qZwjsgVVE3z4M6sOAxxUsLG2vakbrJle
MviKrVZmAZRc5QdS+2FIM2L38ybNiaGLK9HJqAbbHXREt5C/qLZjHifcOnkDiCCd
hxuQPW33RrdxGY5zqT8sKm2biN3j+BR/XH0XYUQBDw2XBxm6COgnK+SAeukQxh5M
uXy1f88VJ49C1ttY6kKCCJM8hWpSofFZWKuYfWoAGOD3oPaRYx1fRjJaj7slCrcz
YVf4tlCsZT6xPJU47Dcb/Odkl45uo/mUvsFnipE6xZc7z3QXFb5CYukR6g7KBXHA
mn8NOQhH7MNZFXEtZPOx+jr1SSAN7NY7Imv8hGlmknf59ZAZTnb3kvJu9x15cCO6
52FJ6reV02+3jmZWe8PiaAlEzgZb6EAet17W3LA52NbDgQ31ZNi7WcEqPFtmuWCK
WjL2YiIKOxRHrvCZA4plTO/1a8DKRzJM9MdLIAGS0gAcI9DrK/BDxEMHcwt86Pv9
zhwRH5T7Xu2kYZ/EbEiFUqI4rnp+mHgzF3g36sOsqaZoYfyHq1EDvAAefBCzKa5V
NN2GHNaBiPOm45Cp+fBF++Y0oHmFRcScKPsR94fdL+7nXnTqf2jA/ekVZxk4Loii
si5UIpzwRzYXrrNUuApDXx841SKCUGmD397U/iFTbghmGfhLdam4FW9jpMEJxI6A
fKvKajW18jBd8y9ALXLb0r+tE1Rd2MhlIa7BzI93BhptPC+3VvpRh8gZLalt45Yx
nVVmZinbhDJFCOjn7g8MGNtjbGR6vNVr/CKw2pvQxcw8LOh2uAOgjlKLLcw43uLz
ShYSCsrmZw08LoiNf4aisNluK3U5P8AwRl/URG+WkYvSHuMbYxSngWg/ScjmSbQZ
KtmAEu5fjydNaW0vU9AZYsijWg44TJQnnTp4e8F7KsgP6HHC4EDMCQ3IkxceTtBr
9NbQk4I2gITF0WqjR56tQ3dgkljAI//XURDCIpOZ2v9dGu/b/MPB12Wi2tUOT/Vy
93cv/ME715fQprsKMrjJHHt+QdXHQv5RACePOoG5ILDM16/7QtKp+OuFYAZLhPA7
VzPPXh9DO1gLJEfQF+4SDiSvylM7yA7RGJ4EzVl1PxgjFwXNFGa66BrhNpu2b4V7
1gMtaZEHHqb5wQ+U+v+HMW75Oiw7gXzf7j6QlfOCuMS1yicbTLPtHE++s0+1hLUM
4cI69e5w/QPIegfL9tEhzZ1LcBbLWJWp/cAqx5N9e4PgvsY5E3rnUHTbC6M2yDIr
7IsxTio7wW3vBzhEfL17tARxIHPYVyD1Js0Tz+S8NgFY92MdhbAKj7x4quESDD5c
Z7chygEBV/RdHK+Tlaxbo0F5XE5gfM48qyKp6tr9xxnZIE0ygaylgRzDbAb6QHUi
HkeAJkR2BNapVozNpUnSK/zBkfqV/+7vlYZMgvdPrKHTEmpixulmzJjfZ7orxB+M
yxeOdc4r8pflDRr6TgqomWS8hTt11vLpOz3A0LMdFh1G9NLCxbLGFiLes3mBnInD
T6KrPUw8x7t0aOFjgnwi33lLoCMaUzMD6q/xfdRvG/LIooWwuWeze9aLm/KC+CSI
EyC87Wk2RPBswZ8Eaos5cf6EyU3p0Lcsr4EqaLGouI28jc+DuaI5UlGRW0jRnkkH
sBQzTglK1HllDVnsE+rfwk0ap9T4rUzc8RoWsdgqD6Z7JN8fLPfmzT9VJrFKGOXn
Jz/4VXwNhNA3ZLnNAzg/kAXy8U2BWMoIT+q/f/ofDFoP5/KI5chtq2q+V9lPAMNg
djG0P/J3ri8/bYwRKDdo4rLD8QoJ8+AHkAQhd60aUbzwpcoib7YEjHUMRQlvtsyE
BVlLZPjg3UcO51w2D+g9vffWZKkTgW4w4K+otQpagRh2hd1smx5dTflvoNtoHywt
AWcMRmAHnCHQHdbD2JaGqU+XeLCmeHl01LQIfgUP/L5ImuxBloQJlMS3jo8HvHfo
zoYliCgVwKvpgZ07VUMBbpgJoU/9YX1gz1R13dEVmmSpYxHoZ1SXJoZIzKz6Z+OU
BnGjVh8RcmbG9ds/I8lI+AunYO91CSnoJSo0EdCTqTdQ+txyga5cXMD9SkisyQj8
nxWENGur01wNL5Mnr7w7eI4K5eXP4aonL2mZwrF75HfMVb2ZP9tTl9/zl9fnDJDK
LvssCiN+h9Q0wBUjYBi0u6Ascxqz/pVKjYgUT7OsmTqn9jH9GADBq4N/+MF5PDwX
fk8cjdxCslMtqtCfaBz64IUjg7sNsRar2EIqdKSL1NmbAhZ6DaDCSat5T55Z9ZfS
gYx0n//nzq9NQcFzm2Z1i9Jf9eS4Vc6tkc6ZCVRu9VkY9jOEVP+73JJ4l+y347LX
/MvEKX0lL8Bvm9FPUrqvurPgyy+bDkeHZAR/HnYOBuZ+sVZ0A5FH3TEgMlzzZIRq
AQua9g+m0aFO12Cxrg5yXOUNXHbJCLIfdlLfrB5NpbtxrJ2wPVAnj825L0xJ7V4j
e88Wr6kW/9c5FUOF7us/m8h8laFCquKmwrgcP/TwfRKdcxWh9uRO+C+feQNWrujV
ontvOCMBCjp7M8HL33fK1N/I+KsDXCRCSDwCtEbsDBkS1TOfpIYfsj3U6O1iL9rY
uXX5+xNU9Ju7UENV+3IFt5vztCkzfCNMKDaEXvpF7rGdCQNcQG6Rf7GDWPLgKSLk
NMBit+UFPhqEYWBreMvomq0ForE7xvtTX9pafxVerzjOWjJZw1zmeBVxVfePDrWC
2eaOcNdCBwZxcwuTteSwiBaH579dr0maOtVwLI0fXtTnIUqBX9Mea/vstCzj19S9
npOyZZjE+TRrsLQLr/wKOceNIYloHe1+IzhdQNlSTROhSY1l1E1qWdYBFzctpC9G
H/vNkMHtAPljRe18d2zzCOZkV5AT/DXlxqBiaXmmi6gZLm849ASnerb+YIJBhN4Z
kqGdtd6FvxPAdKKcCA/mp0T43jxqZSCnu0xn7qmhK1yU9Wd0wbYgLSuJYBES8eIW
1ABax5mRoHn7EunqL8xh6EVsINioG6OP5E1sVNfVNE7BQlsR1psYjXYRyJ5gcUwK
QD7mM9BPIUasRqFCOUB6gP5SrbLKADHi6zu/YrBeHgyZ7ahZHt/kjw1FMPvdpPYs
g1Ah8+GqVMj/RSExy0rC84wnCqoBD5Rkwlugw8+3tBHYRyfI1IlZlasTwSs4zDSI
jPh+hfqpTSdNfDzI3ei3w/2qI5b5xmyHhv8vtF4I7mJXTxqkLKM2nuebQZaw0qBN
GrLpNWnxndPEK4AmaQImxzt/5Aud9Ag7gHZIQkm6CQVCl8xP8b3qvsXLRkSsELwK
IK4Sf8Tm1jatp4YnlZs0r0+3dn9sVfQ9AfL+XI2NWfspUOcZcZMhIWNnsFBUe3pM
IunnfLqw0q4OrVAV1Mnt8ZmpkwGjJ30QfJQ8MaZpNqXOCfXB1tzDKka+WAe4Ln1e
IRv/z3QVEvWm5LW2cHbYuFMbn6J8vvSKUIJm4xm8aW2ZD163uK74snZZ9JD332WV
2G2q3elxdt/2DljGrikO12NJgSb/u+Jkzh0yN0RC7HMnS6tMuHVcwdbSr+4E0wF0
DCHUBOfXAWkmp12ScSNX19Yd2UD8mxvtJeT0KBQgiDBVoKEhSNofVhPSrrZYldeo
AQ93vNNTSzpIHWDffAKFDwnSevrUwWhYQMhEtlTIUhTdJmnYleq8UQOAzc8dzaAW
RYmFUlXR3nYi2cds0qzpMHlV2Nlfro+ZGZRhHCxfEOu3Ewrm/iMHYAZZRYOn++bE
nuveK8ChVsUG5RQh6tNlDY3IILyEAH3ox+CxJEJnHSsyt6F/JwkEOoxR7Ab9LwxE
fnQ0V+2yOAKuIxWlWEqdXJpu4lEXRMwEHfKOJfvFDNzStcVpXlVhUgx3RKP5gWzl
3r5rsXmPSUKpM67ZrMNfkSnAmgIhg23l09/2/xjDHNKEcH+pudWFinQU8XEYn1bL
sRJ/BCim9HlD4hZyPMUwCh6uDQTzTSwn2VA0MPSxNOHac/jQp82nTJLziJEEkphR
1JzrkQbidEXKIBSturX0icJZlSfSxAmX7tZBoZUXUL6FXFlUpqQGqeSOLIxdH2hg
FqLgRdGBgg6Ls6sU62oVwNwum+MdixN73o5uHCFJPqLdqMxCpWhGU7kz/dM8uFQT
EzXT+aAZFaz9dvFFi93QVVQTRfHElZg5EVEioQ0/n3DTkCGdFrHFvPUzInDLblZb
A7jTF0PRXCPM/zDEZ9CeDWFG9bvpT4qF1PeDAnIInVrZSivx7r4b9djGArS7D/x0
Rex40RfZ2vN5yqBQ0H1Xh4TZYIK6xgEWuWzcnZGr6VV+53RBpPKl/v7QmaycRkaI
q7sM1zqj+wixQQx+e6EK7wYDpOrhlvBHRrD/iU8Gg6PSRxKqa7lRSomF1fH2Z81B
NBs6b7fSLhqP5BNdQ1whlPMB5jwmI2mXU3NsYFvH9gDMz4qXFP5rh5ZIld3nAa/k
85XWZllaQRpFfFWFgwKVxzMGBPL471pB7UltLZESJ/P6DJi2KXeCiWzL5BPbu73z
rOLiiEomD+7I7kjJH2W7+95+PCGv0saJxDS0nkNu3adjOe66P0WhzAHAH1/+rn9J
hgtX0m7lelQyZ6yj75EJUCengV1llRY7GrSid4RWG9cnOAXCocl5AVbkLDwZNmbe
cnDLjxhPUQf1zvtZthln4Li4Ykd7xXrvGCJdYzWUSg1QPFUK2+RzNVMDOmwMfcfT
3JTeK4qSo3ZgU1bvjQqSLu+tzjeQ7bNC1iBweYDbPOt+cmFZoblkY57Drbe0SmQs
seaYmcnXsD0oyenVVEZBa7X2LkB07jLR63z9kb3fJ6fgNAIivySxy/dlLrt/va35
+5U4YjTCZ8Rj7S1hj/lxTTa8ShQQzR5z9+zy6JKCOJZ7ewVmLqkdkOkg05djbDrH
9I0n7U1pKzAuuIycjgRlbXDIdBSJpZJshncy95xEQJJRzsYRvxLmJvtxlRjx8gjt
SXI6GvUz8+mLZHesLRQl74u/eXBFV2Z6TrG6AvapnMfgjZ4IPGXMUHPZi/bZQOao
tB56BK7cE9K0L3yX5/5mLx5J86dXB3VmhjG2PajAWN/N/Scac14L2Dr7qh63cOUI
3prptkJH756HmmFog7nqLilVUWzzlarxw5M/GEehMsYI782aOxQYtsI5vI5yT5gq
Wu/QlqVSTEBghRjkcaTkeZ+XssNJLpFmGbYhhrfJDGsD5dmNzdbDHaI8NkgPLI9g
OhH/dJ5w4XlKxpfRA38qfR38s8JigZZZbtmRh2YYyPcgqK5IBZ3t1sRlN3kUxDpR
OEO1Gp7V6B+fJ97OA/BeyuVKT/vcPyT5HqaVyBDdqvgg9ap3mM4LXUdLLYc5GSuA
TORVRVZTx2cm5Y2R94azEILqxYbsfNl72jTNa1t5ormLAi0qxrGh18LQO+INL4wt
t2W6Qormq+/pbJLXo83uV0koBaj4m6czMtKjNgNX34TmFCxTheNvllF6g3zqrYBE
FcBgWXouiRCWNArALv11HOolbYOQjcR8/0ZZ881Lc/DyXktP25PAyhQ5khArrfK6
BytgrBt6Iq5k1tRsvJiZaKYmmgM4Xfgd0oFS9dkg+JTJxGF9ESilA1x9i91AWDhe
emI6Mf2QIlTkHUUjrxYYTQJ9g5EbdFF3Od+RCk2nM+QlOji3g3bMbQ/N+XN9XW8K
nED+LmrLf5QjinzneV8HNwDoxmtXkJQXx6FOOAbmnr/901f97gVsaYjnzytXhdfo
E2fzhFDZFshT/aONURcSnXVuBwMyG5koMdxN4srfxYkNW2X26F6zSasOkifmzUfx
p0VgMhxWj8cfTf+n7VF4yS3bPzbqrAmcwiu+jJ3CPmytS1pWVdco8Yd7pl0ayxyo
vAnNyl55I30QUYaaw3irn50bB5xHbNkhKWjGQO+jSlYLFm1km88vhe6V88TaiJ05
k1DcSabCxQSVrsPbxzZ/yoEVakuSvskqaRjfxiv+2lURMEL7UviHj1EN76WUUTlh
7kKx4zUiM2tvyfeo4MX4NG12OyO+hvD1EN17LWEC0t9SsXHjd6BQOERi6/76eZEI
AiitodZqKpI4/b8I5L2s/t5a05I856VYOKgHq5w+2iP7VrxEZpmTrH81TBlW0430
/Yi6CvBmSHWoocWk31kPZruZJ2DoLPUMLWbZykxYlHsa3gDs9gKtx/0wLqgr8smp
J2IB7OloJkZYQV1DT8KjHx4hc69desizCQTMSF04MXjWLPaOQWCogiPGcHPQEnQt
oH2J4gbHuKkr5bmZUYEdBKthHmSNxU5wJc491Dfpfghq4fgHny8wunvLwA+JBxID
cH2rNzSF+SHBq50U+6aZGFAfaI+arbiOujWww7CkgXUmxV4fGTr4qFhJ5VRlIju7
wHDQMRxbP+jL403sZakL7KL6LLI0G9TMwu/yXCYndAMqQPk0L6sDMwrG1oGjdj7F
dDwlI3/W+8SZmvlzt6574t1QIddfL4WoQfeKhtAFNoiHUXOUPBlvjqaescYLGD5E
BLyJ1EIb0Alq9daP79JEEcDEtwJYmRru9uBKEXbO6VCFMZmstNszqMGtq4ZhMYJP
mIgUrjDjvy1f1jjKJpqcmtC7BL1qNuSUHDSJdrKlzoTq6gna3WlD0hoQfx00BDV8
E/FfUd3hURtNAaOWi9CN2PRu3kH1X6AN7ovX78HLF67+E+c8Y5T3/KbKOB8RCn43
BBP9SNVYA0NimTEyICcnfQcYSKsNR2yRVpfkFXQGT1R7/1cngMaqMpZjt03JrYAn
2wYKsWxheCUYgWr3Svoe2HF4/bAMdb3PpP4HHwAfnXrVtalol8e5rNeMRMCrbZwc
jdb8SJsqGYtiN5kw+KcyWDeMNnwWoHc9/gVWhQgXkd8t1X3zD/I9VdFvN9r3sayp
PEvwC9E6fY8M1F3zpR55KA4Kyv/BQsZ092S7B71RBQUlbJ1hGwR1wYY58/BwTTtT
MrLGr2FBtUj8GdCJeYGfBWbvXLCYGXMFIkBkUQIyZoyXtgBX+xEu4awwR5z4cJpw
TNIeTAzxzDoIUI1rVeIQVRD4jocVrH3GOOkbczwEEmNRHXz2Bg5GzNGRa/CfNRMj
0MWwwWzafmYtTs91rswWX789MleVcptCsgj4hjNAsqJEbKlTNfopCbNZuJhWP9tH
kR63p/H9QiI6GIpsq3nwmXGc7NXtrwYf1G3vVWW7ek6KpcOcKaOMGOkZKnnpaQXX
69C/9AWZNjzYjONBVERCS746bzgaOhalLxg/CY0wqEOShNVaGJ6xqbMdy8vHqIBk
c0JkRlyDgNa+YcJ9aIgfFf/QOJWbYlrsbMsXrucfAKKWVDPX2FC7sPYdrJu2BszG
voTuSfCyIrsOK/YAMeL2mEwp4LqlPjL5mRVlCmHcYKq1QH86VMko/ug48gPFe3ny
X3crmFhky+BqLkdAcvOYkyBcG78yqPUHKuCSdQGxl+VVFT6OQyg3VzSo5n7EL8ag
i60wiWVN68XqBZF7WbrWNwKf38e4Rlp8yeF06Bot2yaIOPpLRYeQJWDKp79FgjLE
XwD+rFy+dNq67nljcJMrOK+86tcbCTelishdzTzeuYr81Gle9/hEO8uJAS+SZPw4
EnWdIwLEaz9APVmsV4CmTJTRvLDpQm9s4Vb2CCDBM59gFMkXuSk0dmqbJWWHfG+p
hecX0ABSfPNLj6AzuyeLW2EJn2SuHbcBNAFzqY0ISWplqiubX/uUj/XS2VgKbMgR
oX2dRL0O1fI9To54I8X83frW5qUDnLjf5XjDOby/H4UOWPkZ0E2MlVe5Tihe5QVp
TbQ62cEI+ppAtT7HfeJFsYjscQuDDPZw+xtnqPQiG1C7gKlDlvsQEqGii6U6zvG8
xh8Z0E1UJbbY8Qyzuz8o9usWNN2e2HrDuSfXL8Zc2pS+NDDhDJn2U2gskHlJ46yA
hJwHxhyTjsqQhmo2ZPkIkCjx6ZpHK74ToZu93MmLhc2D+8JBQFx1oomDCDiAnIm/
d+h1vdEAx9IOUAxl/dlzlHWSFnK1btzaIisl/VlAgPaxoIy7FkxQgpZLfCuITU95
6A/PrleUoRWw4AFrY1LgMvAfJPsfLKaPKTtgKbJ23xy1kTDjMeE76cs6Ta1F3n70
qMcYdHQjVJRk/WlpBmrO8AzlQvAtfQQx+vb7ajtJLSloa/e60PgBEHiw6BoSpmVS
UjrEn4L5nmHrE9AcpFthf4aURWXf9i9gYUjYj+W9mkeOkBDnlcXKdjzlVhciNeEo
vwXdxiLDZCJ5VjTwk91KCcxwHWGGCVUjKNldHmNqLlRca9NvYPxOzH7NgT8YZd+q
c2XtvJrLnmQyd17Ff2uEAPqesBLFyfjA1EcFPEYXT7WTO8SV8D9IqEZUlgzRl/E6
OnWN921pllT/N9Qk3P2dp292fmDPEDnzOShzZLI+EQge6OqZ9HfPyloTToYD113M
sMNvLBrPPFD9ACh0IPkpPnLBmtXQtpuhDVcsVIdVxQuG6upl/o+dN8hCXhwPpFf8
ruUuBhaNF3IG46LNuW2k3JmOeFhKdld49QQsapI9d9+uQiyGlDtUD3UK3NwxyM6E
MOHZLdQck1dMDJQzz/WXmvBViQTw5U69/m/Nk+lgmPE6qvLdPhE0uo3M6p/yYn9r
M1rY/rsgWIo+4fSJVki0VuHaBlxmmlwD7T10hxiN4+kmLIBCYntpIEwVSUkuIF6z
RXvUYSk0eA6aYrr0fKStx9h4XSOV8/at7h6tcZqQzCA2rTjOx3XMumnEG2MYOgtd
t3ExVlGwWn2MRyRead81GpGXTMW92TpBVXEM/SqX6nO1ryc4lgLfJ9SPjPypLiDf
IiTIkBl3qQUKk4WJPe3i/BZgg52FGJ6UwsRV86pd+xn/IMgE3RtvzVjoIbeCxRn9
1zHCK8CgJH5ip3vzZ5UnM0Q3capH33S5XLOBOJGAO7bD682I3XZ1Lx4XjSgLNfTa
WAWrolxHt3K81qoZxEEdUaYOQsMCYSU/8CiFF4SL6ahzibvv5OnIhG+YQFDjyd87
4KXNlawy2pNUhhG5HKVe5LGl1w7Sn5j9TjzxUKc0KUSqMK/pIHBg5IVA0mC9X3sc
jGkJBOaqmfJFVS3w/CaCXDwYKR5+Ko4E3T3kkUqIuygoaUjGnDbIseTO3vpnZj8i
0XpA9msjRYLyOWYq9u3TSsnej5j+iUrve6YUjNhG2EpZoYz5Aotg/ANUPxF6W6v9
8GQ2q6BL8KE7IQlg4XtJg3rI8Ywtq6lMj/4QHyuWcdDQJbfc82NlXqCeJF+VN4Il
fhxlxaNnLLGrXwr/+VsEfFnqCq1gahSm3MJlEqkjfbYqNzVFMertvspaGHKx+YzL
didmBS0n5DyzVnTH8C36ARa/T3ku8O+xRhikKvyBXfNCj8MxaCeyh/uzRyBlS6+1
6A47q42KbqKNKRrfOoCdwzOgfCBKIeFduYjTTouSYEehD9Ek7zPb/TPeE+cf6nun
73jC1WraWlvd98CGAz5/VIxvVg7LuE492RySj5C59XnJWk4eL/2IY/aKdvNT1M/m
Mdk/qqt3REvtzxNWKDbTozwXjHxV5hf62/5PNx0DZZnRdqnymckcTRelNSNiFnBK
MSmquKwNbuopuouLQRBU6TZdT65aJM+2NPfxBu6pbp+lgYXgZWRIb5zdoXL8Xtss
hnGm9gN8fa15byh44d0ZQmQErYjLSJFZhKZ3z8JJGQaan/fl4abAe9hw0jEIH0bG
YKFc6P4JU2n1mPnc/vXEf7+/ls+4Pv+xT6K7bDWMxSaygSWRIulZTMu48tmeyowz
J+fsxKoi2zYUIAf4CkvfsEDkOzrEhisxlFjPlE7D0JSq1fLP1r3OZQsyKRlwpwIb
lh/TdybIr87nOXy5+v7YosAa9ILvZRlMQyEKNu1nxIvtHquNZAhh246N5+pD/U+m
dO6z9FwEXkyRD/vnmZU0f8FfQpS3UwOA77YnY25ZjAWqdQGdS6eV90Jjov0NAiRK
nSmrw6vfv18RRWSfldNyrQJvYT/ymafWeg3CxcgWSVo+GqUAw8VyRJTEJvKfmnBM
lz+Cs435jvbjOv0hGGskCuLLRU0uOrs3Bon2L8CCLBMqyDtfOzQ2hxGt3kZTezCb
eeHec/SeKvUbMYe2miaycXm6GCmYM97puvHPRiwX456ra/zIDWLCDQrljmm65Y90
UPSFISpT/AA2JeOEzR+gLeILwoQSay8tJPe+Gf0Wt+y4Hsl0BSaeRvGbW2eS1u4E
2iPVTwkwYPJP2pkzC7BYEpGEjDMKBG7yc5VR6i6qQtB0wMGjY7M5ZaSxYIk1lpfg
/uEDtH+cf2E7u8pS9oj7OnH2l1Tdi1IYhFQpR4/xKlOXdPUEaVsk5Cbw9xSE46pk
am0W1IAWlNIRfWLXcXqHzK3Lu8GjzGO+aEwtZGiuBkQRD4W3poOXhvFbZjTwjABE
m4XVRGPuicDmB8jKhDEaUIGSyLIgzSTV3crPXNNud0tAqnb35zf/ATEc56FKk8jt
ZneL+pKybxprnfy8oqAqXZEuNMsnWB8ETQ8GKCxnbUeMMHgBPOw5S3ZehoLWqKtM
h1IKHvmjp/TUIjS8ApVNXC2UCus/kwLNokq5xJ91OpW5qviMuRUBuHLcq4V0Xu6b
y5pQEJZK5MIqU0UDjtrtPAlgQHSqem/DHJJqy0+AetwW9T/7Wu1QzMBX9X4KD6Mq
83+N9X7rs4kb2Uvl0Ktu/t4dJHNxVWKu8JpD2ZjHOfbWtHi5aM8jjkAvTKfZF0ag
tVDi1Jfn4hxHPC6KtQt6eWtv0lcuqLykIXc8qCeucVrN5exfXcNeu3Bi90zABXNj
42CTW8tPJbnigmmq+l6p4T8O06IrHuR5wNZhIiTF41PHaYqQeIFHDTBSqdcwRF/m
psYbMHbMX853NprG1fFZ5Tq2nyV6QENwCd3xBLkHl4F8rS0C/qbLoeNoUTs7xuz8
hgyDhGO/83ePpxW4PelNW4SdfoJ+dzBRnuOaluhFc/l9zdh4Geo/z8fwwD/NKT8e
1rpWV9tFdi3xIpxk9sCX8DRZ5nFxOsZpQFCpEMJ7bw+4qkoFPPyqlf01V1AzJpAq
T5uk4nmJGBCRLRvtzaXZhBnlHi2dGoJ7nBzm73WPXBpydMFHSgudcvM3s8fliDXm
MxN3Yo+yUs9pto63SFmj/La1DKXLKMJ7FVwXz5MRNXihF1H449d1Ek1ls4r0lmS6
XjLzz9/gsQ2Nh/nSfVkVBubHD8/CxptR2Gw/JY43Sadh3cUMzbd9eyzNBdc0kT2m
5BhESfnoE1TnGpdTTXPPY/OseeJEBUDvhnQEwUa+xOGsVVqHNVf//Ikq0hDetF5W
9lcAlObKe1/PPfxp3gfV1bOSi99is7DWeTb4Svt/W4ykycR46kDI/oa+CoF0xYr9
yUUGaG/wstN1KbIN05fI3YK8sY7S2tnL/SaCrOqK9FdVKECoOvSbA92l+wFcTInC
wwugcFGKEB38XxS+nEpr7hLBZaLlHvMLfkBrmq89H60eKfyYdT2cXLEf+uByd+v1
E1CQixzTnIobzwXxtgSNy/YPA9RHZ2jGDlnjNRFJh0jZgFpDG4Ffd19QLQIujLAC
mJYL7cMP/ufHNkFAN2effTEjxiZvv3vyfB/HwbTYG4VSEYohhCXG3YqSlLc0HYdV
bM1Gd6hvDPKnpoxVjM9ai/CHZawkRjxO8Taj5vxM5V2h69bcR1DR8YyXaI5qknv5
AsQChj4NsKXQeCzPkJDUDhTEY6FHQKZ23kVrUiAYxWOnSvJOKM8V4/clmDivTBEL
9fjmjwIOHMFNE4avkF20TMQwRa08wj85v7tqQKJH9a8Vgx6Cqlw4j9NsojS2UnVP
QsPykBttnhvPtmY5PXlRS/F9yigY6UyKtjBP9JuhD/61qcDiwBLALoXmNAaOJphw
i762xk3MH10pTKGOObHlWXfScw11Rs2teh1LmtoAdZDSn0Dru8M6VMX/0hnYZPSz
jpHOa8PUxt7vk3b1mNh2s1HE5kdRZBivZiHvSFNjzHCi93d0b3XUIozZ7Lc/vbU1
DtYg+Cnu3rSwicWI0fv5o0gUUgDX6tjzQKetVjAoi4SSziv/Oj3Jz4rrxtwM8CB8
V1umZke0oJnpvRBRCNGZsY1Aux7I0NJ2tPwuNtDTTaUscqknV93mONhogEhePDOH
zJG79LOjFHoi2XkVgIUfs6BE4YqullMfbICXAUdkUqfYblsd7t9L6hrvV4T3rOnb
Ss1dnM86ndT8gUUGF512+9jH+7MGnvJE95BcxMybYryMARnDeYIdjfzfXSr0196v
aRNQDRoOyPmfk+EWYdKxLDsYYp4jPNI1kwWrE40eDNpRN8ZFGouQrlozLYy2y13m
L62nsWpkAdXP2FHHyQSGiY8ZFJV3Lr2OUfriw8T7fuu2GyNeE86ALKfEk5h2G41P
32sYttpY5OXj4BXMcy/SB+3cJHywSaZwW+lJMtHVB5/tWmiRX5J9Wz4C/MwQIevK
WTaHZb9eDGf0OVCMfUbGR4+zT5oCSYyRKKfFNFQH4A0raejx4hJQ/bpSGqtUw4OE
UWX3zASrhYW5gP4fRkmlwfnzh3ItYnq7eanD/mhsY1DsJnksDqgG2q6TJ7D3FXWa
RJeec0WnAYvzTEfsA4d2Zy07ob9z7Q4h49yt8MApuMPyliEm8Bh3hZwi4QIAsKuX
m8OSeSY6sOTzlB53o7sFPXI99Er6jHU80h49nNi01BBNAgRKyW9pJWbEnO+m3uHe
Tygb3QevHuv7Rs08qmlZplTLDCNJ5AD6RYC6Vr0cb52Psgbeft8veYTeeMy/dEQ8
D0VvvODwCfKGc6K4uLHg+VM+PFOyu5ho+xvOL2d08nhM1uA5Zh42CUpRdIPonmZu
R8AW5D3fp3AwKXI6sRYTr59WlyHA9qO2sF7bHf39/X/ehSwbbkGIf217dmHlJkhr
uLluUZPUWSk2deMkW3e5nU6IJvkhoqfSW/Je64eml7EhGxBThU5CNrw1UCDegzBB
aC5zCoe7d3OUQ8tsBehHsbaLtywz1zMIETT1u9AP5ksJMGkykm8ceulxzjX7ZmKO
ypY1R6lK68s8ehodjPg83WvgnMLV8QQDLTTIpImBGrzfiVzB2OeUYYfKNjhmWnsp
wYy1ruZOIDP3tB07IPx5+ZCCEQMBdr2eRVcogE9zznFe+/Zx1MMYuPZptISG+OVK
ysuYc1pheZ1vRsAzGOCC4FKAbVEBWmQftOkIOEtReCtH3dj6fHEhwmraP1Y7u0Db
ktcZILql0y9yvBiyRthS2+GvXraFgFxaf7JsDHg+2NnIi2YZeHSSiIzvaoIfqGuW
+8de4n7QQYqKQ276Or/J2OZsNGXZd2VNZhGGy1Om9hLjY0SWRjJB3S6FafSjGqPd
hxNf9wpNxfcm3mQNvrs0+1/FJtV0yhOaYYrS9Jp+ZXiBNTV/UP1aE3yhvnQIsFij
hr3RrCY4IcJZbObHWBVGz/WppS3s7tWD9+cV5VsDcuwejz2h5/AWZSDDMTNKtkmN
kBQjOWZ101FtgkOJn7Z1i5mVo7C7ju3rGubm3bF9IhcfQXZIutQn46Ffxn2yszaw
uMIVFYbLpRXsJCeXDo+Z5KpFO5wCU8Qy6c9rwdQZQ+0aq+Gy34V9DOgJC1j4BgnW
C0DFN3ivyVDZOnWITu3OIh+Ac4h2TTxamtd0FbRKiRvknADP8NgJGdSlZGqkFm/x
CT9na3jz6ULULTvYz1hIKGzqntLQdk7bCyWC1FPcyPzbLfIhIxq+bdryPSucK3IK
1SBObx+KOF08msDhsj1oiPo64NWbbmi39mTJASTG3D9fmS7WioD34ODCXzhMJfEU
wumujNl8R21rLjqzFJulXe2OCvvRiiT/l2/aOiRWyaki7jgWCAqjP+cE8T33aGWG
a9FmoukqJgWwhg5hKvvIJ/q22sGqzEZwGd1CpVnKQpxvXE9FKYj6EdddT4VKV+j8
Erthe3AoQcqF3txNDWu6rSmpAjQGhjbf113KZcCY/mlME/MkrNmQj6y+NloxPW8l
QYRgV9SbbbUKqVZdEQviUzY4hNLjO4JjKrCrOEkQbG/oJH0/hWcjCHVUOky3kSNL
eEGrUS4SSg+BY1u8bBbgSMlxh2KryYNirX7hx1ex7N/oW6tMLK+YELJShiil1h2o
pQzRNwtqfcCxNy5n1TyEJnf9ouyUcuonJrrVox+HC1c8lNNCRtviKUxdmdR6YhvE
jZWQr4chQ9K37GfdgHhW3si2jD26mXpK+KuUeFmfVm6cTlH5IfIeVXQuuPggfAaa
W6MfCbo59Ms+MAUMhI/I6WmobuxVOvTxE2TK7UVZ83jyBLRDiXvBW6USacMDOF+t
rNdHx0fZKZ5UjeJTsydSvKNtvSVCHDi14eH43STe6CGZoMr09WdBpcyC5r5Z09Sg
Mx43bYPLz1XpRmJA3THZi5bgB2zKBOmcu5y4my54eDhg8fJr2aXRsbiPKQkHOA62
eNvwS/ZrtlfdCcv8d7qARfSxBvA3kTrG1V8sHnUjVF7FMMA9r/dls9ZtXxtxYZaE
kR2awwSIcFLEf8tjFIrBNS8lQgF1wVZGvAscLPEZF0xMk+MpEx7TRuTcG+zbr/s9
XgBDHaGl6eBHxMXnBscCtZCe1Ijug+kMQ/SPvUQCsMXKffY9KYH2rYtQeeitgdQQ
WfsjkieKGAcgZQ7tUPK8CziWeb/TtRkoLCKsR54KGe4K2nD2/VzibbTJuyCJasF4
mTYafzkfGgRrXPwdsHer9K6y4MiWEFGSVzNuz+1EAUADQnwx5sjnc+27IxNiE0S8
Epx4L23KU90W4byZekHrs4voc08wNbubmHvvSfdlcZQ7F+7D6GDwd4GaHA6Tq6bn
mt3mg+Bxyhn1AHxNO9sSKVM5R/Oz2kO3DoOXvKPRYVFvjuIZFTJXu/IQI1vyqAy9
judqXk9ei361N+AjBvs0y2fjEsCT4dD6kaJn2NBOwNlOrZKlueM7zDKS4ETDKtOq
U6sI4TxvffmaLWdDgx3I5rTfBn7r/hB//gtFNpgKboBELNhAV6RGWOs1BnPEIrK9
J1Ox/4lKgYxJRL1VI86w63o0B3l3kceGNVl8qBh4e9SRgYNXaE2azgyUoeWmdNz7
dZhWruWcrxPLRoLVG7tFidmL5iCwFiLPq+Ohse1/nrl22dvjUX29gpPJIV6OgTyX
yd3c3HS+1bJ+fQAX07iwBVzMtDgYt79Hn13OSpk5LfvVxEr7Oy79eTbYtOi9yap5
oYxMh0aCxo/Gn9exarOoKd0lE9eoRtivO3Clg54ZS7grBdpgYtldUypSZzjCUwxB
QCLCzt0dPHKPXkQewh7UYVJJTyjZzrNZz4kOSMeAyanRAKZhpM4N+ZbV+bEc3UOl
Y/jZcCduZB4XvKxygee12VYpDFgRwWNI42CtSqsYBw97wpFEtyLx5852iyuxI0cc
cZuQYu7JQu2Em/gvgSLUBsQDwYMRnIkt8L/jdjSzLscCYhpT8zxor65cmagRZqCU
cvt/kUL49c1fUcthkUb4R7RwnxMPhZN7pidwwgZ1XrhN9A9/Ocy3jvtXNPbjzXNF
FddXs00BB4FsqCcr2+dVdccFlyinTxLTVp56XlpLNwQ5mOjR6IZ0ozMeh1EKUz99
mG9TWrlRKTBPbM8IURKDIemyLfwhDYvDE60A6KfJhZc1FSeHcCTZojaELdRaL5ix
b6YBktFAWkMVhLfDiEUUsfg0BAwHJLNeDnhxZmTNG5EH75hndkQd6MkylDucDsZv
YOe2oWrDDGX5xBuFGGlr3Uf5D01TD01yi3OFofrbb6XzXkKHENbsopdpVdQP4gfB
t9N/Qm9MyNBARc7hRwZ84j0Dyjjp7UUUSNKFBcq7BMObbMp0vDnFN7SVxH2Okead
LeDArBQG26pcc/T4X2SVutO+DP/y5pjIJUYS6xj+uQhIG2w4mtZQHWjBD+Pmsx3b
MxgNupaRWK9TzVux4x4SFS/9IxO7KW4Rrgvf9OYf4CnsokDnphMaI7xnDP3IwOq4
TFXmNLVLlqx8gi0f/9dWvSsXe9nmfcSBVkIBU5mCAcDJvf7mcriVnr68HlCM0y/7
2mnL1iKTKe3ESHC3j5oDvshOUgA0vpedfHkCea5tWzs4uZOnkBqegZpbUVDopD3u
ByUS8djQuxrdXqiQOWYLKs5eHAp4+5tCW8V/4JGsYujoYGqqzNstxThZxM3cXb+w
HIC4pOo4cU050ucgDls7Ui2mbGGPh3PN+ONy41uOTuEyt8yG5rDNFoYi/qilLnLK
JhsqjcSsKDQt1DXJ6LcyoHdQsQ5E1M3GepoT1rjtGXbDhlHi5XYH89SXes3H3DvC
F9VgYsxptFWvQozuWYuwKaClHEV0UhtoguF5/v1XBKLouDDQPZv5KviX7wg81Y0j
Z4G1bftgDn5Hb7/GBo+f281mpRx3MEf1wm78ZC8lvZyU7tapFuLVTpEypMlHiLX4
68kwt+utAQ5GOPXJ2hVomROZvUtYLfKzkp+oSW/VerCmPRuYgkEmVSpjGq6eimN9
rMmvYp643fsSK8gKGaygZISWyRsnN1a7j+LFYmw/3P1BQuq4910XMDzFbwB+EjiD
H8r5ltPOiM9X9WZFWgdN4XuKKJQa9uhQND+tM/o8vGnUoXD3Ar1AbiaMbHhP2/XM
i3+dEPLxx6Rw9uikNiBSivpdIH32zuNuDNVHfD5cMBKhbE1YC6iQc+9zkZThqE4+
RKaCrSY8B90gKB8rVLQ44O0OJ8ZHo9ym1XU08zZXO2f8CMG3sVzIgtoKmPBA8gwe
9X+XlY4gVp/snYBf06dlECxJFk4//JZ/vz/BRSylkTI6UiWWMSI3i1ow6N7B5fyq
j0fXJaTMpFDsuECrFkoNziBNgQbR8H/mCxDmZz7fgUTqXBlZpVUHudp0NvGYhZ7l
mx605S9ongApqSh7RHYs4UFaeHxqklId+G72g+wvzTlsQei1AJ0GJXg724JfjnAm
/Ya4uJhLxGm6TGUBuPI9OnZ1XJomQ1fYFKnfQcfCkL9bBLUUoumaYjEDaas9Cjve
ZVWLmlQpN+oQt5bNmwAi4h51T1UpfevZiXCcFoL6qmjK0ZoDhMt73nxdA17Aibv+
+utXYS6bGG8kgWxX8xy4XQ1NpOdiDj4YZCdFIufhcuITh9NML1VskTzuz665WHF4
E4xHN39xjOr3FC8mpKIYsjtnKoKO52r/PH27I35xBZYrw3yN5veQijHmBhu51Lej
1EGtLvIJs2unMjHG5whVasRjvE7rRtQSPuhiE+evw3CekgUU5+95fZUPqwSyB6G2
QDPUpi16uIbciuKKnNWHZcv6tsDadmSr0NvmWgXnTthV4dv9K/ivB8P69A2jz4m5
d7Y3sq4MdUCTfkA2NtMyQGLjeSKXdyDnOOd+B6dDdnhhUsT0X2XhvW9DJeUKwt2p
27vmDavJZk6m94blYlJHf3wNEQIJTdDP0RGhScIX/yrJBsboSeL88T45am9MKWpO
AI4Eg5Dnu6/XqCdfrinOR/25jQFJhKHWu/kPberB69om5IFS1qBKFncXALTbRH2D
4BPmXyE2gHy3RMyfRNdJlSYl5wQns6ApIM3pkYwB+n1ZO1fOByoOaW8HRG5dbpGs
kvBJJigQ9xidpYbYoqYbbLpfgaiK4VeSBT9U3KDkKvX+fZHz/zy7v8JxjjKgtFuH
MZabqPVdk+CI1no7v+b+rerak6u6q9lnELBEdOTHfKiFiiMYgkAggH1E1KnogyC2
KuwyTm2/f4sHLaA8ao8I5Lg73WXeb0KgMbqZSYh3i813LlZEMDGo+49uCZBqS6cs
reJ2/eCIViXtpVZXdZAYa09CALeTJhPZtwhPFpXpemUvODqmNHHYfZbpG2r88enR
j9H3zSXzJv96KuCgEOSrF5w0Q5MWEvdneXNn8mB+g+B6VmoWPe7aAefbmvEYfN2f
aO8ysXLA0E8aqUijIUoQ+JKQRDiN709i1VI5lCcTn4ElVW840QFa2I9eY55gmqdW
njrZB5s18JydpSRJWejrDLX9OG6KDYnI4Fwzv1pWbsL2iB/FXNuAzHM+cUC7vbz/
UvRkANTNhe98xnA/tw15rIFEB2Bn2ldOUt7ovx3HaVndjBTfkUOLPg9b083XwhIK
SqY+I95T23RxoPygeqGRpEEZA27BNbijBvxnbDinTi2uYozAIlLqx6y9fJA2dpHr
UZiOmf6pPNS3fiWq8Cg7tPW6fcw2R6Iy4LRbfuHXoYnCYXghQyzMjg4aM/+J6Hog
ifcpb+hkhYEO8OdldqfXbiyeA4epM1xvX+5jzON3do3SK3H79eg+9Dhba2C4O9U1
024rkAOE8xloidMjrO7QWdTfrTM+eMi1kTyd/IS9Qbs8smlEwGZ50xrZv2krthMZ
Vfuflhpn5zKXe0Qoj8HkaOU/XaIj8+q0avuoqJ6HombrV89Wt4yfPT0W0QR5BZvJ
/0wB9S13QH1X4/nLTH9XEGaAzWlv5EcFzKr+ChzkjNEKY7aZqDa5Rd5RLLNESCDU
07d6/K3jDhKrYVt8NuBeXDR/sXSqqJXaseY/FCQdVgOZ/SsOfce23xcoosN237Mp
Ey87ezPx91zmUHVxeY5uJCEeM/+ZB20cBbrnSEUZrw+i4PDo69LeGEGZAM2fTEQl
xwCZE3SXPsmZ30z3x9Uk2ysl76VDGoDFIWBswA+Kl4CyBFu/Y6S4D/dPKc3hSMY4
9RWgVFXFn10fAkOWop3QZWCGOb2DgzsESA6VhhreT9S6Xp98txpYThpB1WvE047u
9QH8NpBBt11aDrh5t2/k6LCeqUirrvXRLQEPFhFzhTyYnnwPR5pvastmIWEcHDGX
dn1ynRI+KoZFODqnogbiBWZlUYEq9+NkSf9wY6qpU+h+pMtWBf8dRSSp8Rmt67SZ
pY7r+YmZq6YNe34htQmQkbwCww3fxmY4PDXmlk5j4BQTgsZSmEFQZX1LAeHHGesl
xYbjk3+tE3+O9Ms7HdiiJp2obZt9xCL2J2VGBb73Q5kR0LqlBFqvwFxgdOmr1NgA
Utab1DTgb7WOZXrH/XXfH44Sffp24gcmvUF4awNcvv6utW5xuEOEdnaOI0hZptRe
c/7WQPLMkLj+jUYAYNrusmcbock1ctToTvEyB71DRAGAghRhxQ203DdZO7sbeW/W
ywVWtavLbFmBaLlIFStT0ZKBoUuY0/DNtJtR9rkjnWrC3yav11qbdCyrXfqI8uuU
3dOVQa4t5c9Tnex7UJ3UumdySUdvy7gwyL2I/lsW0akxPiTRdHKz5ILb12N3Pacs
Yn4Xay04TQweC2XWtWCsCHhqVQMLbYg85M4HXZfTdpS5xSjS5isQUmhSlZcqyC9L
KryI/iVl/ooAP3g60VWSFV8IY+WUD10R89tXBpn9xiU3kikI5QvWEnYD1G0fPE9I
r62gBDNS/A9IIIZVkisoZCKIRO2NkO3aHEwVHePUx140JciADiZZPN1+PCMD5Rxi
MeBDkhyhG1G8mVo4EIJPGjHDiA8YmUQCaMxbthHlC1b7C+HF+Z57x91LtOPDG3wF
fQViaNbYJ68FlPIsmD+nzfPn8ixw8oCxzCzrX3gybwcEwS7RPvQ1J+poUnOU0ycU
4So6+qg38UK+NltcIIPCsPEPsXkdbb1EjgK2j4Dx6B716sISeLmM6fvSmpB7WQe4
MzEhnG25L6EK7nE4NEsBrbN81aMF2S+t5aIAQbuDDET2A6mxYJpYL36lpXk3mLqz
NIMDBlPB51sBIg6Dhk6mX0WPFLYOcb2zY21Hly1+01AooHHVLG+rnPfVPjmMtKCn
hpUlsHmJMsSxCTIczduDLmtdLnaUketisArekrY2SPGK4+m+5t3b1WAaEZ2UoYar
TFlu94bBxXOegYhtCZ781wlNZosvzhR6tWXdu6ZSZDKwp+gdm5lUeMnEvQMhYcNR
QDQ+EIQerB7WDr01Yjg4iQnTfsT5Zid9dkiL15N5SXpPnl43sGMa7WJ09bc0+OnS
a+FuB20C9BadYPUtEi1exsYSvwoNYi1Mr/Gh3KnRBfwuFmhY6JXbklu7CXmP30hy
lK5bi03UPhZ/ZSe9HNLybnZEgAr9U7v4zvG4L2POGEHwVtTE/fs6ItOThLb6mJHC
N7WhI8K1vXOcQuIokzTlh2LuhA8yl59eBq12TL6ti15DlCCDwyZSoGo+pM/3hiBo
BKuc1tDv+zaNDk2/4Nkoeo1lv3eAlE9MCC4iGjYk7Q3UU+wr8rIkosQ9lPE4b90B
FgtEt3aV0CQ8H4PDyO2beFWpzEXZvMbiliAyfa5CzYmmWRu+xkDK3kR4t2vSM99A
sAVud/y0Y9FbJpNwSpabWLZIO74jRy3TsjxS3NxVnEddbhpzWTH8nr9UEC9ytEH+
KRWCSCZiAoAKh7Yn7zRKe1U877KCU9Y6h2CmHpgEfxv29Bh6hTAYQeu1DHqJyJoF
Su7fEZ3CGTo+qRAhY5XoL4xiN1BtgxuLwJar4MIpM+Hyg3x7liXnaglZ6w8+OgMd
1UILKlv3Dr10riJQRXLjbTSpv+lWSso5EGtm1gRa5Ns2lH0X0SOQJckroWsYjvfg
7KvWc8BSSSOKHtNSiIUVoLLY0FtkigRzburG/iCFWYjW92ryS26dEMWBrcB23Elx
gkwwByYvmR3irdvYCx00eUznqzc2xZqO70GhFabeBON2EuiVjOdresl8fiiq8XOX
sLoA2XT7O4t7HRR5vq7hH1jsD+NM1EshYaDGRaCqcFCACZayaRVc8QvTxqh7HmV3
/dGcXmVevAM7WjzPGhpDzaGfIHCrJNDJKFJfjx29TZhRVOAp3m56MRyKibEx9WOs
sP2J4J+8lbBSOoMsZZX1IXJfaugwt3LCBrHl6VpQ4Rgs4/ocCYdL9vwL35AXfPzp
nx/agFYwLJLK+b/M4QvK4PcIms0xjGnfPrt9/MMx93cSV+zuskL/PaRVXnkvJrXj
n3bbHEht5iikhDeF7YkXCKWob2Um8LyQwf3uy4kCWwBRT2O3wINdZ0rHdSRh7bxM
u45k29yhXI7edO58qv4Wqik2SfjLh4qSpJTZ0MyMovMy97li+os2iK018dWHQyZk
wpRfedydxDslHT3ra7Yo6VnD7Cv4lkX2lYEBnm7V7F0oU9kNPd3iqO+xSVru044C
vN4QcaLJxSel+MeTgf36GJ15oHcWXGthe25cu1yjrzQIAMhL0EI/HNt17vcx3Qug
FpXKTaOkMvXJOirfAVPJY9GrOvnVVJoqfk2gtZGqOCoCS/8pSpJn7D/V5OKUhf5l
9yO/9H+fn8Hc4bsnm22NinoUNdHHKtCDt0IrGs5QmlHG29qC3Pe8O0eW+0J7sZsO
Oq8UCuDn1Wymk5ePrbw8UsHSTw9KwjJBFriNOmWGDzAB5B4KL9PixexQa06GFFK4
td6l24ljrwFm7sc7nbMGnoP/LJDPt5fLOtB7v2JY6cZKwpUKApX2Ys66o8ykBVHs
7byJC9LAsfdgwokFqCf89yKO4tc6g6cy8cjgBfirt0Mpow5HoNgo3u11nuEqJLEV
F6hslcje2kO0k4Ki9Vp6wdNtBh14OV57jR4klscFEgy2Ko3+ave6IGGSsVKZnosv
48pmmivFg5VN3wHaJhl6a7W18pItNy+i7pdvswMEF/Ey0YM2xwtSXhXoNLK1K9L7
DFQF1LPm+aENspDe/Np4k11hkkgZiFbLZ6GNV+kK6/G2+WwxJRzM8OYDLigjXAR5
ZIJwAV7iBuN91Jj6BLoBgi+WgItvjDZlfgXiINuWURDhqhqVEYKGOPk1oavR0F7a
aXEH/g63BXsnKr17EpBoA8OZRP3mf0MSHUVP9qd3K2/bR+x/eSuhFuHo5Hx287WS
gigqLpD3c2jpe7aAFLYiPhJrg6KOknpDDgS8Gxcv9OZhPxD+1Z1E9bb1dgE5OHTs
jWRKAiEuTmn4dfgQ9AQqGB692Vi2muEu3wmhnkjutIDMs7AhCUEJ6OojeNuEKdhl
/lSAoMwVXaNCCcVCw39uWnMhLKQHXzWmLEBIRO/BLjC0XF3pJ7MNCq3EGL3HUMTQ
wCceGRVX1I8P9OchfQMci8L3KoBE2OuzXicsxlMlVJvyr8yKfN8UKmajsT+qCaEs
ii7ItMv7CTUQ5aV77ygSaaH6gsuF3b1ABQMYwUt8tAh6UInJVLw4SmY2Nnt/Ocu4
mm+l+XL2wLXVFTKz5MSA+gA2TSRN/9YmwdBYLu/jSiyzZVCj5C8EyN8W3shgIR9U
ISBIAkJfgXgkruH6pAUITbYnidY3DnlafAOHeYwmourAyLdpYq3fnXoKTYuDsanj
Kw1EFCsymLKWCH+2oR+dfQCPwefahmVKA+1z4KpqtXaGsTOJafNsJMhZE4cpogvk
qNgDOQxo6H1InhglKox+QXbvQ0HG2acLkxryx08STc8r/oN7XaobmUmu9EAeNshX
+Ih/n/utXqewloA3MVBZrxZ+c4pySEnQQ3dDNJt4P5/tOko5AwsNU77NRLvf0+aL
GkVz56T9XbzKezEoGNiFDq/l2O26EnaO67XXyr/HD8GtQx9D5ta30KFFumR97zGn
WNNMhg9mLw4HkjKu7jhPlSnjEXSwktlHXCoOGMPd9J3UwQcG0pN5Xn0cmUpMzBdj
Wk9LWO1Vpe6t4vhQ6qXpb9Y8MYhu+nQlL3ZEb6bK5u2ptDP4ZVln8o1s/TgeHt20
gUCtlavVedULaOreEpGKGURTjeTcCxcuWvj/MJ5F0yp29iWSNQn5+fw5/JOKI8gC
edXkxWKrx7b2vA3HdgLCXb1CLdGyvJe4kcNL4wsMJhm9ORLvHXFPdZj8HKAerhry
DrP7W82fQmut4ld3v6Dd+5+jHhHitE6CGxIwgTe3Af3BiFibOuTlw9w9K2jwyR2d
GmXHzILRYlmodARlrdxR4MYPQLIja+FF5H0DJTu+JJzYlQ0hBGhFsxYflzLEq0JZ
UJAz35DT+NRBjruhRe7qB5y0ETj+7POt2l8Xd97PGcWTTVm8wJUhmNi+UB8AsxYg
T2/HE42pPaF2xipSjFOptMfRXoHO5TqS0Ov7hFitLHB7CD7jlQvt6L43TApTCP8y
NCgjD8KY7ae6HCvCjenREtihp57ZOXZyfiO0j1QL5a8kXgZkLhRQUKIyVqpMi5N7
l9jGBArPQIqkhitENs56UQukTIYtGNuWXAwoS7tVFz1Qrj3x3LpcqKxhEkR4u2y+
pKGFfVveqpiDzuR9fSQhHOVV3ESthnRPZ3/xN6Y/c4V55Prid+Y4+dRgvgmsLjIP
mfWCDiCDWRe9uVXxlNOayzEs2zurv5cmfOrqO4s6qsLua6oEyNueG+njD2Q/yy+j
etzmuMICoW9KI8vnrXn6U8mDMsz65C92C/BQeAl02tC9RdRny2jep3QnbbiI1mf0
bqgspe/uAcKkQK2xSnBOLiNxyn2ZsFS6Bmxh7Z4r1FNYqA/0xmkXgT9U0mDlN+1t
pSeCpzev1I85UkjOvUThK0KLOXMuetpQYn3iv3tUjJo+DF61zGspkVp1Sk/lYMf/
QjOMvVBErIigxXTuwX6xadK85lGq7h5ql47ZBqxIhLrOXtJb4QG+R9KlISpKBCPP
L+KllSBDJOc6ooaxQYlfe6UWOoAf25xChVKo5gT/oagzbDapnWdYidhjC3ShtHPr
2buUdtond0ryfcmguOiliC6pZDUHo9oB1AUqXU1IRbUEDeHIgnGOg/5qAdqWp3H1
wRDyYsNUHHoQPs/eAKUWZ0l+dnqx86by0nXVwbAxDNIqiATTI2a8v8ahRk44vdmI
zN9lTs0e0TTDnVTIPllLnrdQ3W3Y8b+YYumhI9xfk8de4GSPD+cJwYQUj/Sq2x2k
/TVtR6Js/nDAA7febEuDOQv3qu9scMZgiFhCImhcJfxu6mvSZ/iceqXShUdJcOwR
CL/XYxYwgRqzPQcVCear6fkm3rw0RqTnxq4bJBWj41qC6lnjfHUJ0rKX2fTt110T
bp4sHpNe+L0G+TdwGX45xUXbrTPYhbc9jBriNhfmgVjt8ZZkQNzbbCsvi7XhYtc3
4wiQseRgKn9H5XOuM6OHNS5i31bDLPDC5g0++BdPslllQ+yVkKDFjr5IgqnbyWao
etSsOGGssPNeuUByUn/91VOSMkfk8LjD4fAwa4bHEbWlj+7WZVRjW0ylyDk71/Q3
BBphJstzqwTKDUTSpUdpkwU0MRKDAuBdPJqViEMQhiffxvGiARyJPKcDfrmQKpGo
mmtA7GQt6jD4hMy0HuvaQdKTub0A/8FJJF9mttA6qVxBmYARMoJhSTDTUOMVwT7P
gdRPDxEVJALgDC5TDlWxaKx1MUv1Ww/KLHrlhGjQzv3sc0IWACvlyKtVpKHGYj4X
O13z9jBaVYYpHXoQU4b+13IUsLT9Z8QSWSsu/vRvPnMHoJk9EHlgjefz0sAmWWuN
p25qK+67tl647SA1ulOt2r3imhyY22TeUs0YaIN83BE4rAHwjPK/Nfqn2SS5Qf16
qYJzqMncW5x4eogWOwVcTJEWkwTxRkDNH3ezkkls/4NCdxTfINLOaaHPLugJT3nu
mv38Xi+01yKZrSLofPD1yEkmxMcirDpog1PV0/jlDGPZiH7aYh6U0Xo8LeFpZLY5
cs32QHwtgoywHsiE56LIxQeCjDPc6pYc3WN/A2k6VEljdytGkyv2oFM5v1caiT+7
nuDU9GgwdOfHQNHiAOakfRkQGkeTeFMw3MyICqNm9HZiUGi5kJ6dKIxkHtxony67
/2txos+09qkD7ehSoh0zkeXr+34r4eA1p76TkKSk9Jt2mYBbS3ymM3kTD6Gimj4Y
wMKcb/BSOgJh2nluv61MQ0t3PeXaCxxEY5/jOihuj/FgcWP6wsAhlMCrLVtIpZNO
MVoNamadEwAViITRb+exM/f2IhyK0lxx09Gre6o1S8wCJuIYLE2ZZGh/pRiQUGwj
8pkL03x9y3hkm8mcHZVCcaswTNpidSsLudPmnKnFv/EiBJawI3Aw5N1lh4yLVGDi
rwvbBpdEQB8qQ3KZ59HMQrF8go0RCAZIpYgO1yBHvYoqewo6tk8TQ2KMKK3zDgbB
MgKWygZrn8+bpVhP46hR4TtJCl20wHG1zX5aYcIffwGs1z2EV7y5LcCCU3UgMne1
pG7IUQt5tsWtMkkGSJNbd5wM/ndq1JpHYjDuL6JzqZjMEUBSGvE8vw99x3Bo+LMm
//RjY6be4Jkl8Pa5itfWqSsrZPwESO4FlXp7yt+71K+l8UZZpJDYmApWPXlJ7m34
rr1IIM8qReGUu19DCrTuLFXNE/FR3eS6fL79eLlxV15iCpZ5sAHavICcFBOUwwu3
ZVV772ZA0tcPhWb2lMqTMlwLXmAGpRNr0qWMEypBpDol0wobBqG0bT6HGoeP20YI
Ajb7N/wl7/Lr2bhnMp0GJ6SiC2ismpLr39mjTcyMjWOnLNwcMz9G8fb5ZS8i/7AX
wHOeq2nfza2V7Dtne5AudlvMNGdDKn+xNdcSC7zPHmJ3qWkzyqHxHr0AgdaR9fgT
d6/DTd2/StJoSDhieUEfgLvRia3BFZIkCDJwCFvOUxt9K5S73GZRljkmuJQXdLT0
PKHdeZN9SOFIr3rI+bIVsm2SV4htxeV7sggKFy9V/0nhadkowfKjBnFm4Ux6m2Xm
uuhwd3c6kMHe+LqnsIc5pguJfME8R/fIGsVNYy7/cZHuYBat9bYaNNSPygspBosG
MhpF8lQ8o46b6Qt1B2MrMD5++0npceb8JiGer+ZPusFbTR8NhzWCfEMln60dq3US
NnUitjj/S2Hl0GLC6pNd00zOIQwwuGxtfygzaAA/d9oe7+RC1ZPrcnCdD8iWpq1G
XgNsZQYhhW7AQTDenCQcMRRis8QbXhC23lB8Ol2vpKNdJmnoa8Jxnh2kd4pQEAxA
drBagU8m2O6HBDpt4TXL6U02v/hHW+MiSCs3bXJz2kZqXGGJavgPynzDaFvwgGov
CBpTUzDQv8fm+iV1mAC2L+ntQW0X73M8sqmfMFDBeIjvbKrX3I1sJRGUyETfdJLu
TFflbOpZVZ0QmA+Lss9k2YlLwqLJeHvLYmETrqyWrQvJsdZqtC27Uc8bR8LDOWz9
sYAF3r6Gra2eLEtp1eTEPYWRpIQYNCRQWFI40UpWvX9MjOrfDmTSMYtrRGG1OzDS
yrtzNaCbu5LnZ0UhvMYK34ibbGoMxOTltBz9iSJRIGXGBb9DZqj94uRkR9wqVJSi
/Pz9rYxXyR04ld6bpp1XF2JZIo8juq/HfWzJo9hzDAcxnJM763i8MIr8OcGyz5BP
EIqn2Xek4PK5kfkuBGmtuycBA5HsE4ZHlt2n/C62+ANJJtajP6Ie69lC8xIumdeU
kZNfUnc40z/72zqi6MRRmCWpC/bA1Cvm88v5ZtCpbjmjF1X1V9u8WTcN5W39Mq+B
KcyHLQeMA3CVovaI9xGI+dmrXMeaIOce0SdTmEMeSWZKNUa/r3S1B7WKSXq2yn32
BwhhOFxofq6A2zVpcsBQY00NuPs6uZNKhbCj12sHUGXprFlzS4tVi9SGnSmQOd/v
e6zD5xUHepYdxENo+M3EkCWQqmoU4OOwPzzJkJ/6ZfuJS77gUZRFMMxsFEbNhfoG
gY11XSqAur55ygP40OVNwGEQF2EnWeSQs7gQ+khuIycXbtTqjatDfQvV/f+l5Lsb
kpo13h/HPPeQMNnMEvRzngmBgg/ed80qfC/Vg+EnJCPfzOacKNvK4DQDWpfXpn05
QJUCcpjTCTUyL/5z5KGdwFvaZOb/UpPygMQbTiksMCJHo7m5GGtCVmyKGAE7Ggwk
PFN7sUAorUbYzbSe/F+3PnJf9gJQROO/7X3UzJEokd5EEj9DQ8dNApnbomdBxWTK
51DujVUZSM4Zy/N1A+JmyofTNLVmbeeOE0Ah9nux7V014VZzGenNMH39imapUZiZ
5qqA2QtRqWmYZ5LLySzjeYYK4OhJuAkXzXOfMFZcdg+n7PhmyAtxGqPfSSlGJwH0
8pWnchpq0ah4HcoCvnMs0GAD6VuKTz4s3ji8Zwnffy8ohBsRhbwkxCGzf5+s9FO2
OXgJuYmz2IxrNcv8ffYXREuw67ONPR70MQr/fVMX7QM96ZKEyp3i9kuFXf/GJBBa
bdmeBzgvhbRPbd+tosoNqJk9fEVsUK/dyFsPaJO9u06Pc00Y3SC4fcnNVvau2rv+
+blbdt1nDjGHX7BO/vQCiRfNY3Op4LgpT5L0Sclj5t7fpK3MXczYV28KHfpo6qwA
7d8Z/5E0FO0fNPtZ4OdKxHgba9ozSxjVXio1/hIfrR+UZ9VEFxxYmnnYBja1DEn2
NGgD+ROQxORD9shaSC6KI9imTtNfta1s95g3npt8YkubU9a9ZnCAUBWSlSPoI53i
dDhy2xecc3uWbl3O5zjXduCQZ9MrXyGGW7nkQCMhTJZJ9C0axkhGvC9xzrca+tnv
szhiQYKQCbFeQXe03McTPED/V6vKRkdDQq/U/ZK5LobEOq67LymhX0NBNDwoD1nj
XwjdbkyKwYwfJFBpYb0hMcr5GXL3/YVlz8tlenpJV/M/fmzVy4uDJBxMKyGBK2Kz
NV4E4wsR9JSVkrP/+9RMXQHavswLvmuyR/bM9+lgEcJl7n/a1lQ1R9ZwpE78CHaJ
+1AjlzrRQt+kI3kVT/Jv/Bc+k4SekbOzewjnvmhlP9VudKVdD9GusPMASxTtwZ0h
orX5VbdJO52kTvFxYgGX5M0hFdQ4OiU6llZnjfIxv7TxPfy1F8IlpCEL4tXJOnRx
1Q9OpCcjf7o39S5QCbIdP0nyp3LmTlCtd50HL7OVS77jmii+6B3QO6Bi7VKj/bSz
8qb7UCR2TSOFmojSWjFXPD72oN6MGnneAdkdrkqV2QdzhVnnD1rP6+ux3LB5//ur
X1/PfuGKwSvMW0y2IoyG3aW0SzJDXZrPe7fWtaEutkVI3ZRgDND9n0sW4Ct75HVx
xQ0eSbkbDylIQCgr9t1GtmeTmH6oplBdb5V570ZvpRZh1880AaYbyy6hrme7k5RG
t7rYUFCcTTXkbJzPO8OTBH7wbBUedePmC6OQxoZoIWjBLKLBOJUi0d5KC6/f+pPg
TTNwdNm648/EKTUqIjt8If7e5zsdDtJzcfEOuu73cOV0dbqTnLLPuABd90DEkCCY
ekIblB++1bJX5fe+roF56+Q4JZD4mUCPNTzL+GQAVm2Tclx6OlzzCsn8t0U+k56P
Gpmn7I2uVMDExR23lmDnej8sK1NkY173f7FLhgRFjFpUC1B6h+qBGbeYp3DHHH8s
FUhBoeVOnBc2cmIxiSaT0+KsQ6UaQFcKc/XuRrfwnhTuT9UyF1ZkId2MXePaZV7P
wLKvdu1WJwMworXHgKpGp7ofsz/KjYigGbWnl341MyhSjjLFMq9HvRCJK+m4EGhV
3LumOKWLtGhtbJxLMYGWAJCdUtKpoY5vbWmpPshzszS54/+5ATTDPTVrmZSJ35uL
RNwV+EEQPcckTZnzyE6ksbgy1OiDC63BOS3hfscSjxa75RvUT9oJV6A7kFsaW3w4
772BkC8IXjU4TIpnlOqBnuwIS6IWjOF9FqCyuedT37oecq4/1JeFquITISZj9ggO
1xmv5p2CVCbbKiMzyopWl10HYy9QtWS3iQj/oOJ+29LgyyK1jHihDveevAETEi0Y
eXrVZSAMtNKSX57nh24Bqh+XE8LeknfyIcI69EEh7mqNQ1/1R7gTLQ2pyUIDi+cH
d6rR0ZCK6nzb5dtXd7ZCSPqJPZhTnYtM3J2bdkwOI2TtbgdfVSg7uRCIKtOj0Qq5
R0rHOPRSzzNK2sKxwFuR7lbOKWTMBwvXveWKguT1DiKYnRfpg8nLxniL4/8ywKmu
E6YQgLg29lLmtr4B48f4/xWxw9bZkyyRZIqzbuPpXEw7NnZeMBtpOzq3gD0KGyp2
9vXhq/rK69ZERnQoAa0+ufbNlybdZqYIe/A4ogJmc7iaXrxZDC++9Pvot+yz0OMA
haPaYV8IDHPX85MtLjrOWTi7tV51HLkCPiBZE54jsi7/yGshi6I0c5QMJ+9SiOGQ
zAC/j5m0nzlIomNfGeMgH/XqPGitVqPAPqIiAALqZynb5QI5r1z2qr5pacN1qJ6S
kF3MY9gC+bzw4TM9tdmUu3Dh8ZgnvXwJxd1FB+FxUi5NnfFtA/uvVu9AhsJuONgK
W6yiKsFjjVvqHeqIV18BDKoq2Sf4QqRN6ZuZu/vMkVDT8yGGGkjPzkutJrGIZiDq
XvOiIq7hdm6iwcWFJFc6LBHnahMblJuSBREXQCmBZZVt2yOtJqDTGTBKVHhxViZE
ICgMAB/KVKOGuDq9eAE9f+4cP3q27C8momzpVYBlXU9oSzP5+Xzj/auHM9rUW2Db
Nse2O9e0J/HMMb+4r8nrTrCOmr6qGhA9oOxMlbBPQuqrtdKBY5hBDRK0YOrz06cv
Z4/YMhAJOF+FE7pXx9EY0BO9vqdm85I/XugIrfuj0bCsQeceCZNTbNOSTISB0exf
Q8EcaTlSnYTp12+q0e1dtSyWJxd+D0UiM/ntntCKHSPDCEK9BFjgzqCrnX1LBCF/
VN0UlUNvBUIoPvfLIOYVB8R/SBQpkphA1iYoP6hjS/YFxLGk/1hyeWYsScbPgqdO
R/u2GZPfGyd7iTdWvX2fpO0TeUWWfNFyGK0XKYQalqAFIORv0KSod2nHf4jh3U0t
Ej+8t0dNlqGrsO2lkw/rzw3cNDT5aCof4MWcYJXmTtzrCJqytF7mGd3+q7NnkWNC
giDO1luoDqAn6kSVg9sArcRFnymfeNYDnCzTNagzmAFaTXkSAEkg4TrfYvoYc+Nh
FlBLQZHgE9R2taYnV+aBVTqBLWj1to22ZZvvAlsa20WaV4pRrEFtUsX2lBPSGZXB
yABimqzzH6xARgLnKplcISnFJbXFbYdGJXAVn5hpp0LryrPuE6ES9yw+VgNXEE23
N7Qg6fXp1dkujAE2HO341wFIB4jqURdIjG3wokOrvSzPOAZeTKUU4NImPW2CKVRY
0Lz0IowGzIsQWzHuZWc3FEsUZ87od4oMBGkNRt9yJ/sAX5lTESudbYeJM6T+CACf
fSG3TUXI5Tif54YGmtbq3KBNR2hxl+BNmZsEZZysrgvYjeVHe7JnRlgE6WSmNYpF
UB7IdL8FXG+d3ZIEGyb9MFJSyyAQ0P/78FkoaKi79ga7usTHSU/aRUEWVfMKdpYx
C1UrnY+4mAqCsZBf/eNtoc+zdPhZmMBKQYQsI9lG4L6K4GqNFlEfXwD6IZpEpMCH
ZXv2g9lBe1Wx4uKpM+syUc8it7yWzL7R9LezhMabUv6yGIvuzakgS3cf0gzp5QOR
Zyf4cxloupkm5ShDHIbILWiQCtB9XmS00My8FUtHP+bmiQbOIchjfoa8pqZ6swF2
RAnEugzb/U2uRQat+YtwZ85WyY6RnxhGK7c1fQusCHDKhOe+sz0ievuqWVG2WfmT
5hTcQhkweL1HonppCmOCfUllEgXctpb1OfmtXD9snzDVyvDKX0+pw1Rm5pKNKPIf
f7jkKSIS725S6LLoiAj66hyPSDkaj8h61AW6AzvhH0B+lzsmQjqmjPte/gsd7ikx
6BUW5BrqtrZ/HSU89igZVhuZPHy9vXuYDT8DtzQ8npTSAKN7etEu4D0++rs5w8Vc
q0Z9+zbPMhNek4TwsBhxt3LN+/0ObfifQCIMof8Z7gz/mQQl1PUNw1Xrzq5L5X/e
FSs3c8rRs4bWVhfgA6QUGs31xRgRS1cbQxc6UZO1hKmY1ch8ZK4SfstpIStavg+C
lb/7NfQbFdFS1n08wuOmnsJnmWVWg22otyGvkx8N/CWjusfpaDlWJhPruEy8y319
fWHuDC4b/6YwpBVZQ2xorzBmNFtCZ/oRcqLJsPpSvXiek4VzRa1zPrvjFPAX6SRt
R7sEjtDT0f6uobtuMLGUTIWivqEdYxnSm7vTvJ8OhVVBUqQcI/N7j35l2m0jY9lq
f5/fAuJ2O2pQ8yulUfHg5MaOcWQe2g4tAh7mLs1tBy4kqOoGjgpCQf5CzbWBguIN
efdUq7uxHwe8s5dtBmM296exLE8lXmEneZFEkCPJxQZIk8WWrIwCFB0ncuWU2nrX
GjPQGhlwCqc/kXXQmuZG+PBrEH3PCwNU9ofXub4Ta7TcWlItxfRD1Y2KWyTyw2XW
fijyr7IygJVS34Xiqom8ZfUXNC0b44mzab+LvZkgFDPmXw3wh/LTQe+UmEgS7nUQ
YqlWgny8vngZIN80LShdIloYr63Y8BZ9mUQlSSj7+4T3XTwMIjbH1GY94WvQUzWa
pp0RCVOJY5QgFI0PL2HoXZFP/9fmSd8jvkcXXsCT+aK5JiHoDBynBxqo7JPxH+h1
CsK+cTtdIPkuih/qbB2qYeSgYKLfxFSFyPFYIRyJKNg5eBDz5K/vOEw5M3CrSEL3
hjpA6lUJblDf2njmI2X466+RPfFZ1utewtrQoukRXw0MDqt28sulP3KawHY1izPw
wplY0a402c4526Js84IF4k6E8L9fHUYbV9HsAjB7TNNpMvKJPEc/Nj06Hj8YWCtW
VX/XzOIN7U1kswOQu/HcIUFIAcU2JK9cLeFYjXqbYqXIlpCwUdPsNyRP3yknPMbW
z4bRczGXA75jVkVCJjBjpFvoA0l6LsZvuGn99PM6wk8d6NM2r4amLOEn9+UwxB99
wnFV4FtNcVYOz4gYtT9hLKMR5m9DI1B+6mcMIPAQpd9fO93Qf584/S7wZaQv/fWK
Du+QywzU56CJW2tsekYketP9Wq5l0Xgo7Pfx2UCvIo/9FOacKYeRmACned4WE0md
6Bbl5JHmoxVjz0Zps3qNwg/MXuy+KEeYpKqdGa9K79bAbHhGuCX7qsnWWET1weMP
fDsg6qKotQCmqfNgsMV2a57IlO2IYgOO5MBoR7XoX6sdL9Z1Ad1dgLV0vcIps8W3
jAvb84RjtmOFXOv1Ts6bjOszWk8RP39SsJJmgNMcXkLmzA/nWwHtVn55fNAsVqFG
lP3D7KtS7DpmJzJ2jU+BRstG/arjO5FcI4348RKTeSSHhDUEdRq0GarnQgBegG/6
QnwnQeaq5y2p0gZ6XfASdxkzAy64DWARoZwpT7PIiv8TEaseWGVLaUWFEPoYw3t5
VnetTmWY2Jzriya7whKZhXTbjNBywDasx7qV2hF3NNPNHWWoKJzORbFYXZ426N7y
SpS7SSy3/6lc8KCgoOF5FRR3WxzFjyH5pdHLspB/dB7S+uEn7QFIuZGaALYI4ujv
TzuCfj/kKqjgadOjacWI4pBMvpa+nUBZVGwzX/xwfwYxZi697gWAMoCKo7HA9bKO
p58XKHrtaXyC2W5WIUvqXuXS7fFOE2gwdF6f6L6I2yg6c+5UIVEV8Ad/EtOr2Go/
Gl6X1/BzQecaCnJkjsg+2qD2j3C9FzTN/MHA6GhXXecGMO4k9j2ePafCmj9T32jH
HJ/OU/FBdfKfc9t9lOw5NRO5TTLIyZlYSQhtwqaVUd7r4/ndAxSN5eRq1ukeyUcF
Zy8Rz5WJEKLqKJNXwUdmiFBJV2srA/cCuP4onMAyyO6jrgAdACN7yLE2aCg3dd9k
LJgcVMTaINSy/v+/QqihXCk/brjedSQZ2J0So21LNkgKW9jEz7bD+YdpIH9GnLeW
pzwF3NRrk1ZENDZn5tTWErQnfq0eBWGweh68Qf5m/tTEVhTQ0/az+PelFb5Cfr+3
/L6w09QrJXemTB8K/quLd8PLqa0QgYtWf4veRvkcJa3T5P1akMEyXCxgnSvylzhw
OuDcTllZZm//QClZpI+LQP6A493SghNAc4ldqnHh4YsQ8xDjIFOdiLwxA0aJ2Hcf
7ju+kzdTruNCE0kb/HEn7q3VlCSRBNrMhr7ICUAaRn7hG0fmDybCFwqm/uUYCSw7
5qNab2H/DxTomVjchFILgMp4m+2uCKBPbbtQ1bQ10rvYYiuaAK0ihnE+f2aEVhdC
asB/Pnso1y5axwAhBxvIVhOEItIpfXjm8u/zisU/heO9tsUQX3eEbTJDcIoMaChm
+pKHGWKUWKcRouM/1kp4lhMqZpaWP+dM0JmqzpwhUgAQIgFJy7GKtDGw9ctiUAnY
6WSVtwPlF84NRbw+1wY+lZpHukTGHMS2sY54qcH+jMIujDfoaMvt0HdoKd4mXH66
v8iAtMP2VPOmmh8t2CYs943t/vfJHbWFw/PQ+n/LFPPAJdNqLuu2GvDHpTkcJ693
ZEeaK8wbIBk2bepkcPL6rJIkOo9hPVQPrLwpmY3E3Sc5Lo33ekFTVxkd1rH7wO0I
V1WeonNaaHRRcCE7bh5acNyIvwF2YRK09UyUvncAwJuYM9jd0shBBHYjgzfzQwzf
TGSauIXwdZS57F/c9b/QfzZ7ASvtFxMBN8IDvkW9QiKO0l6ldPyRYklJV8b88DO6
mki90TGAcDaB1pr6dZU6mk7U2+VtsSInc7qSqDO3BUtCMVHWofmwZL4IRbFuQjyR
vckyXKVGRfGo/Ep2HCMhHZC5WpmQkxQokpQkwmSyvrbEKgQIan0m58jOq47fhbMV
MKHoWCNCFZH7Rh9cvyoNIZudcy03z4412DGCEHBFsIKUnWkyOlKKVu+Lb2apky6F
zEAY3KREF22XAPdK6BFiyUYJmbZRqi8TZRBP/eWVPTroAPESOB5VT3xLorDo/uHH
aFN84BnplHcNWXwCfFamp2cyCh8P31IF2TdnD2epMaQMtS6mI3AZKB6pMiGVSvmz
CS97rhgIBNGIj62gP4eGC8ZXmBaZ4uQTe5FjbG02wpyJRe359PhblSRuCgbPmIlF
rZf55As6uWlOeax3XNrwLyKfZPDmx3XRKVlxJmnn1LKHZgV4m+K7JH2zwXDyTgoh
JPDOaS7OfXRJGWJaaZSb6zeVgTH1w7m6b1zcwt3bqQ1xWChf2NoKgGC8JaMNYvki
sDr5QkHKFXN7OhFtIg6UrlsHG/Kzvgd0q18wyVxNtNt1hAEhb7pfuOxC7TD5UVbA
GYKx8XF9yRDidrzO5qxKg70cs3vo50yDTsusqs2ST4jRXFzBn+mqtnE6iShMM3N3
+KDgXF9HiXWJ7KXoAdLEE0ieRpL4MZuzEKRpy0skfVdUcK3+9Wv37P262ZFQOr7s
xH3WFDXZySBuxIXdvNRZjuJ1bXTOQXkQgNDYpxRVTiEtsPeCAdl4umhaR+uJDp1C
+obbvQ4iyasIw9lwjsdzlMWy9+L6efMZrXlO3XS88AIe46dQ9xAWRWN3sX3JSQ7S
jwII72bJK0Db89FhGVcSA+J0bINPLRpG+h8DnSrQpu2M1AOKZcejZ2OsvtCvrasX
w69yIlR+4YG5HgVz9991sv5IR3dedx5Wawtoo/X3NLqMsOKrBQ5ngRSJanScKSZ+
3VdbAoZcawF/eFpeUSE7GR/88lYy7nScFw9uQSVtCfpr8eyEgLDhSL/1OgxTUMiJ
Cg+DqPDbtidGWeG5YlSbD/per4Y2kXDJWfB1xlnj+l1EKOAULqxQaon+UK1b85vb
usby1u4dAdsluR7cvWf50lc7W+wbJYkDxt5rT0Ep41+fsAOZNLPJYULlAgLv5Xxu
EKfqYh2Z0RG6k51A+Pk/Od0f6xV9exKvIer/97sem+T9teKk0/OGlBBVPUzLgoZm
ThZghL7SSAOpMSp3vgmYxrhZd63gnKAhdvf3X+a83kobwNbzhEf0Q5Wo1pG9Oxdy
j2Qtu3+aUFEpdHyHraChImlDZotc60uRoKZylNSQXnDn2EwgbfEeKhbSpAZFK9Vk
WV+84ZEgCYG+UEiXbz/lSxTD15R9BAULprVctqvDnaEEmdaO+YVbygT85nS0sPN9
YtvKei+Awx+fnvziDOEom3ZkWTNvw0tRrGSCjUrTnwVMMcGpQ8Zr0acQ/rLU0fXh
tvRSnjXOfv673Xtj5s/kGidZ2PR0umRWpFCOfT+jazhV7lPEmN474GKyoT8JGbPn
3Shbb0cGRryIX2vVadsuUaoDtn3upUxO6wnM98Nsc8mSvdebvU6eB2wUjOjrHxao
2/IjABiia/jpjVAjI0ZANxqY4JeLw/wTc0/a+0NVLDfVmSIoqHN9BVqPgW8r1gmw
TpWU4We6op7cBhuwqJrKCnGNggirSvWndOPryKMI6JHB0Xl3ghPsl9AOC0ZmAcZi
hySkqmYSDdZ+KbTLSORRVGyhjB1H6WegfOQ4NsiFhaD7b1nx05X1UtKDVVqO2z3Q
XOoUQpnVxVtxIcUJZ2AeEPu5kEFWRw3HR2y/E0ga9Q5VWh0vJ8Pl+fTpJPJ0Dfgq
JoduYJuhD+vwqGE+Zzx7uqkLTQGBdNttWOwwrfqhHnHVBBtZWu+B7XzHNVv+Bzcn
gYsU8BoRtVIFtNJG03kfdpUU9S137NzKUUyiDpIShPBdauzgONIJVxZWwttYsHtd
vcqt8573jnSzwpya1i+v7ShAzMwthB4AM3Q6j3NYZKFoKmbRgkpDfM8M5Wm/te0c
ee/YTpbbl4n4pqKpTwE0SRIdPkGmpGWDewV8O60v+jHHWMn9+iko09easObtr+oP
6IipaP6Wfvnkb+qd+xtpGUGOXzbvY5G4AE2m9z463XAbCH2xCSpg3/iGezco9TRR
+iu+afvTzPRupvEwTNzv7ZN3Zkx1BXmI8fJFEDnuWSk6OwvnBRkbfFFKyDyXBHZY
T+d7KzVI1JjbOlLmUWLa07bYAQS3yNBzUY1TztkMmqYmGqMhGV7YmPVEwvZt5CAZ
GpSo5GbHsT85iTsQV2rgXSLd1vY/KRwXSbyicP/fSTFFwbs6UclYQi89KWNeyfN/
5zTMq7AYa+FWrarmmytJY9QJ2dUgREP+CoSKLV+lRkQm2vdVYXDa3p8E6+BbD2eD
2DCUnl1yMZmBcpglhYChnn9ko8SSF6sc+rjvMAPh6cuSVs98ohtwnrYpAL3MP07a
1zfZszhbxK0xNFCu8KuXEa5b3pLEq888TuuqhyUBCpuVUJeHZZaijnMAGKFIhZ1Y
cFuz1Pe6dkS+CquU2MfZB5R327tRbQru+fge4htPJqSSJnqLb0ZBMvhNUmEhQXd+
+medMgnQCC7TexuyE8IWaCJT/ObRy6ME1oJqtgI0GxFkpnfupA5gVB40BfWjJVf3
I4TwiKiHDezs/7ZGYv+mHkkBlQj+aMiDE6RL/jEqmxt87nxk0JTzdQ3KK6sXcQo8
WomsxsATajgLG6dp/IsfTcBrabX4SP69OIwOqn2Pcnl5EHOfV8D1FuOYvCkb7xoH
x5ki69qFQTnPtIkNUsfU0uSDu+Mw8IHSh5GjucImbVhu7QenkK4TuwGewFWUHf17
m9AdP/UsUBnXKAanDy019F0FJAqpxINiJrhzYibGixCoZGxB2HRoa/kV1dJoHM6f
xII3MVI3LvhW71R55XLf/K4KwsEo/bagm/G3kzCUQiK4LaPLzoSQmnd/Ay7hyAIp
f9SD/6h40mlEcx7nk5YRzz+/w478EB0GJuXgxaXcSiRfsvR9/AdOc6sfkbCT5y9L
7LwdkY73EB+xqfptiw4d5XDoJ1t+Jh43PAkx6ltCAVDJpLn6CIcjXtF6LH4W/pzF
HaWmN7AnoHYhkYTSBPwzKukOhCIhuU4Ez5PPxsW1GfZ+EYnOjNJGPWAnPrt5VxmC
/HvOAyEUgMrpJPJftoJpyFzlIluUAaz5LBURnpjQYZaIjXGvQtYeAX9Lprefh1mZ
7VO2+detYH2G/sJG9I4VGw3XksdADjzL48VXcXT6wRS5NtRVIirNA7uhYpoIGJM7
2nFIt3bpTNOEJHiUvoELnSYaCrdNV0WpfPy1AXuoPAHSkvvBiQ3YzIAR1ClDIcl0
1afnnvZA46xTe42eyU5M7bHE0UdI7dLcg1C/14BLCQKJ7Q417g3zilAulJS7mlbK
B1AztJBunpUhrYaUazyvgpqpU1iYXmY2kUE3dLhygi2s2wyw6Fqs6zSxbn0OWqG9
PRb+cJ7l66h7saGVaeb+LuarZYCXSLgaTa0ms0yo8FoX5/upBJVAriwVl7yCg2ph
qHtlwrsmJKbkFlOxzDIkdqfnZI9dDovxNJDnhz62JcO45Bf5WaDymW60OZGXlGbn
LzB0sZYFy4yAGjFhdRB37aXHc2YYVm06f2LW27yqWpR4zftwDidE/txDo18bk0T2
phIluy+9ak7hfu14YU2fdWmCz6AHrythn135VGZaWhlEayQVWxWGiMb/lP0SqhIY
+eCf5Gm2YxMLN2R3VVRQgF39MlH2c1fp2b1rGrLPRpjF0SON8drI7rzk/FK/Dif3
mAI1m1WiwAtZF4PtN6VBBT47cjw9FkjeuPCkfxLCXfjFSuDPkFtmHZ/MJAu3e1wY
hzMKSVe87Igda0P9OZzwxNVouVxTPCmm8ek1h1UtCQJNy8yPQ+wVmC4FSbwPC2OF
/K6U4XtZ7Ij3lIJdC2kVvfFRkT7e3McwrgsANI6LnQaL6bH0bygXgG+RrmFtonIl
RMsh/RNN2NUfRqyk1cl7HcdHJcnsTyCN8k23mgPRiJuzopV0NdpV1iiiJms/6Dw5
OFgoQl9Z65GFY9QLOggyqA3H4qKDa6G/SlZ8z1YCxOF3/JbTrQfxB7sOajotttam
VFR3tzxKY3qs+6q/I0iB/tbvexqccE3Lmxxr4XrFurnQfQB/+hs97etFBJieaZkS
+TQuHGqAElQQNt+5JmzJYQeRHEsJJAdT3USsky6kmyqUgL+zzM26zOI651jm8dfX
+CHZmGeYPMKSKwVkwt/2Y9SuFPBDSdQZ/CoLBWaWmA+iSDVim4SMv5T2xfNjQzn0
R/Zwt3cndyh+HmDJ3e5HHrSZ0rlh2oFuoIyFNJ7k1Q2/LMoJnjXl6ypdOjBwqcn5
3lNWvQ0u3CbkokJRm6wBwfmMEEjk7xTcP4l8Zk5GN5FsFLSILdSCdQDcKxBd4umh
DRtgQ6w2GHrPd4hLC5gkYkcy9h4/te35C09xZEeV/bcSeo9serEbDsIrdc6MFK7C
/sZgHrDjli9UmiH5y01BJEGMnHDUyhB7kOPk1VoCsk5Ewgn6aKGvHMvDCcpVnDiT
XkX9HBiktYTVh3FtSLvVECdBtmyg8jSr3/2FG0K6UFA9+dHm2vSS8YY9G97x6rCe
reEJVTjuBCgJFg5++YbBDpjGyVgSgiPKFQGUf8qwU4rnKhLXTcFhh5nYbkxHvsk3
umCOG9GJhw8H/IAzd0szAu0KabB3LQ1efjSFPIyrZ2f8iEvoBfMdNsEFE0yLVPFX
G9LJc1JttkCaYLn5RTVP0Nk7zfj2xeFGgkMQHa2VFVP+bDYrmZD81yAlSUvEalIn
vS6qqlE4V34JAyMzpvpnxxoZl0CUyKh55ryPuDIdu+VLukfmNN/r8XlasVbMLHhR
i2DxI0P87KFrv1AMmlnuOk6xYai6wB/K+f9C37JzNmJtuHcpQRBpEWv3z4QoWPpa
Kic0VDIt1SSTc3n41+dhSKoHWu+FJDuYqNKMXI7HHhCZScDppmnkJxpf8mV48lfA
SXfZvH4IaBX0zkIp9AuMg0j7GxAWUm//pAWj5kPC/Yozf6WsrO2cWYJzUEacoeX/
/2mibZX6K4CqieE8b3pXMqRzEmwv5oLheBQNwTROFok8E5GWDJErW60icmnPXHbP
wFNXEtEVQHxqXnEXlaUM/4+8Q5OR0E42UdB2V4FJUwxttumE146TPFI6jGG0sZ7w
bAW9RiCdPzCfBR6JRlmshsaPuIz5ex0llO+NSNGGlmL/oIMkOfiPsSCgyPbTitwy
rFgEKkh74wlypGqNUsfBbat6uJhlY4Zt3lYQdkO9Gpu9c5Q2bVMevmbYjKo0cSaW
qbe8z4HHSyoisGjdzx1Z5AkHvDH5D1+HoxhFIi1JGSWWRnFd+5CwxGnnwlgD9Gbd
0Vxo56iTLobz+zuqzoEdNVQ2l/0K0XQkBB0H1Va0i6MrQs8BW+4Av6DeV4LvWqhq
z/YLXPks+mcKQIOxPGha7pFU/apM33mzC62vLTvn86ys+Q2xEt0LdqKPDnX+0hwQ
sPSi44WL8jjcyhfaqEMnjz9LKotJrzGXWlnSZ0QvSmkuLuAtRyocUXOJmnqLxy+g
3GbsIoMl2RSC0D/hUps+wfMVMbtRvlbx9Mu1b+TEhX0pTKDis620gzKl66nVV6qK
MyAvmQS8GNl6Job9YwYz+k+mL0PHHXC3Zwwkd4G4Dm0SsSgUE6AH+5mrGEIe3Dr4
VMB6mgIRGL1L6BAi9gzdUbJ+2M1MuhB6LcXNz2q8m4CRpVoGwPpIwD+1Z8H8bQl7
LRo7js2nSP767DZugJYxsqKTgsi5J67XNsOM7INVQ87Js19+0z1huq4Dn2afMyZv
5co8AkeBWQMd7gC0zsUD4FiUThaNXCCgOlu3oZELCXwrvyc51cNxhp6N01Bfwr2u
Zuz4cT802yRmMJh/Xx4UU5vZFRev2MW/+uTWHlpQw45Y5dFUhKE5mfoV7mnRtA5g
svOn/Gz3olUK/+5XrWpTDOTgEijF4HBlCzKgurI3o5D/z6nsihpsg5DSsOciq6jl
IMBBwZHK74DiCANXtpjJl2XWJdhEoAgEvQ87WzxarfZ4eS9+cedCUA8vvZayAqEJ
XvCHCvKygPdm5TsZ949nc3kFdwvrJlggEdhdt8GVQuz9vGcaye2q8fE+OQwk5WO1
ktgLKotH4vOQZulP5iK+Kxfx6Txd50KIURdDQ+wxK6zDDbKlP3MWpQAdqU7IYVP4
rAIFzHAtsNW89o0euCFpEPC3s6FHlF+s4VTlIXk9121i5/kLVI+JTN7qFFhU8qmb
dVqkTSNMjIod6DNPua7CqpEeCzjBkyTrgoKi0C08TABVVz9pIjb8LVv3KTmNHUv4
VDJgq/vpXbnf8yD2RUX1xg1ms2FB4ec1sRJiIB9MPicRhHr2hHwZmOKce9tZjaSf
f/VTfTKGHFQ31Yb4oTpTgDQrhd77g11y1VlCNCNJ3ZwtE2ReGvRb1Olz2MDfA2OP
/pQ2QobUcoldVqYgQUx8QkTOyuWMX38maZO4j1SVgJFDfusZrsnXxkgG1acfsdZz
yN2dOXsw0WrZJTgTl4z9t0fjTHBSm8ZHl7GEs/PYbbafUUPdy6D2tTu4xPUhmDxm
vuCUyMy9WRtZnJyKfU6pkcArCuDbMRoiNpK7kFS8qWArR3vslqkpuaDsyp/8NRbV
TFseaQJfmA+PcDhfoyiB9+HwBzrDuSMy1qAlZN+CpLL0bYo2k3kXsdvAbQTb3Roh
fneUSYrWtDWccA3JSXJdbNBoEYC4LExwtF+h/Om820lxU88ZsfpnePCyIW5WKcLB
0n/N/nEW+U4fdB1KmMCddHpXpkeR7qM35tU+Oe7TyTWyzsL3ZpshfHXL3yrx1Q4G
iqAHhie4svOnrDOqp75J+rxEr0B4dywIe2RE4uWSgVL8t1Oj7coDJv6QX2t08Fmn
nfxxeFhOijXRW87RB07ZVd0A+aSoGNqqZp0XfA9hPVumbQ/QAGK09J4WWVxQEn35
woMEmrnz8yyiZQisPeJpMf/eAacvNofL4oQXcVmpte1m2F3wk38DHjHHl2B9sUDO
2lamvrRMGhMKGH3W49n/XZaj91fntLWdq9hGtMZbJpkwf9gRPeSiU7ZpIK0zooBe
Gd0vtoSB/ITXXdaIJ+sO0ITAf6eKdliMaWSpQppWsJwENWp2a1zgfTVm092P1hA9
u6180W/jDGA/lKlAtZ3712xsc07EHkfMDbHJNAbhjLMSkyKnoxangkn83RbvX+WW
X8j5Vkh1pEjw4NJ4uiFGd7J+mrXpmkvlAzLOZUUlHO19JX7wm9BkWt1jdUv/bXIz
ulOwIiYIh3mpaV+2bFAgxPDiQmeO5xrgCWktfFP6IxdoBIa7bT+gTyNSRj0ZaCAk
KJ1ppHy0LKwOgWkoTUVrwT3sTnx9FN8fzz5ZehdEGgsLEbvlEbj86UaZhVpnVBEF
NMWwGJF7qzs0mcyJLwmi7Amb5QbyGGLs80jRe9K2Q5tOmGwyOKUY+urg0VuhSxS+
d5Uskp8QU2bWxWDlSZ9gE25fjqAu8SeMQPHvAJizlpaOeKoleehoY7YDRUoZwj2e
XXrbmwOk1twAl1mv6qIbFygGT4JfaMy0KC33Jgm6ccsz1qc4ij3SYXOQKEZzc8oH
d8FoqkQZffnJRhan8d8hfw/EJzh+LwRWFQCtzScCQpA1b/TsO5mM4/VSVwQ2GYGM
GVZ5n+Nxi+y4SCfZkZ58RJagQvDJjqg2mR+F8Vy9xIiQYdY10k4q6QZybiz/IdEo
jCghcsAefNd5LLgPY5TyffMXhFkltYqZeY7uLrHiqOJjs2URA24RvaV2X9Wj/hEt
TQf3bwCuN4zbPbFdzxl9Df6FveM6D1Sf+ODlgbOIGEPYGJ9RPkhybJWfs/AOQk6q
wgwiSqG+FWmgPPAonGUDbBGIC1qm8RlaHV2aYWMyKaCQzYnlQL1/b7pNBDTcIxxe
YOmUOaMURr26MgYM3biq7MgR/cqt0Uz1WmZ//xvl7LwjcBXEgLXG33XEZpiM5o1g
dSDYaSgh9VfnWelH9i+en5QOZX6yU6gf/NfsLDinTrWk4ge6gxkyPv1ZteJOjm1K
lCyg466WvbKLHJkBhQNS0wIcpY9fli8x35MfweILiAassHSUrnmRdiyb4UTx+uA0
78g30PB26kSOJHedMg0Y9nnWQPjjaKJ6PaZ5A6Y8zq9wU4uSW/KC/toDqn5+WTmo
Fy4lbpPVszdQfRF7OhD55JsggpcWe5q3iBm5epHrZe3scnij83MUCqg04j3GJc5W
yoNUFB2qSaAV4vWo8MCiJVrvcWQ9o5Xnbj+3mYGQ++I/73W5bMiJRYIxbG0NeQz4
UpLaN7x3VsoG6vFVcIyLXM1+lqJZBhoC/VzzT9wKk1YEYnzhwcvXyTdnmeEKdIfC
OGd4awheGLCd4H7f+FD8TN0NlOMao57SIgovCPaSLd4H2ONCcc3XjPA5RbWzgRK9
ZOS1SqhNz/hm0npQuKWmCzs4yFsjaLiCpgjARMjg44gKSeaf+Ejl/I/PNp4N6ra0
cgmGGk6cfx8mrZeppx5OJtuvOspKDghrT7qAtAsnjThZsb3T2ZwlFP3hflPEd37D
ZUE/5xPrkf/FvzCDwDRFp9M3GBAiMFn8005GFKOcUxhTKn802R7tqn+igD9stWbR
FiOpqqODM2Qhs7XuB1Gmb57chMgPuznkRGnm+JbG5r3AgryDW0TFbGrOQy0pwwB6
49jTX5ro1WzHkRoumWiKSvV3FlMFMCx/stOUBkwnDP7gZPy9VIlbakpwSyENjL2c
JnTHGcJOHjQl8BD3IlnQfoOn0A5wLZL/ruJZ+GhidPKeD6ZO+WPd70EOw5oaDTox
qdshhZG233liQaUYKp3ge6rk3leYjxRm9obwhkeHjG0Qxit1ipvFAjWlDRpFBeHu
c3y7MfCSUStqIODUdpUQ6kuIyVflFePx2wvDNh4JLUYfEoeKkMe+Ovy5Oe5COljv
2gK/Hl3t5AUNMB0tgAk59KkMocw+k/bcegDNGPN5VumCiUL5NlKB99m9PnHAyEi2
8JQhECi2UmrsvgR5FtKx6ml1aDEPjh9Oig7tjr/T9GTkDpBQ7LulsTRXNd+d3Ifg
tNXrKymDe5oHDBaQ9SWTOkEFjMb5dA52Ndfm53QuV/1uWB0+m7aH1k2UMeim/SCk
BRH+RQxmDZqPlWO/N1ljwKoAC+it7dp/SXlTMm2es4IOGPS/bDmKpfnn1BohE6pg
FCPKNFUK042gbFdsLuhJWNLbfnOMkpkxb5KX36eiKpApYIWisdsFgGuTrpv8Fl31
Kp59ZAkctb4cXY20AukAg5gpFpcxQOHCqH7HYCj8LgQ5zuZdH01qhVNXHu+1K8b0
hvbKcAi+LKsPkilTNsF5H/eJGoPQoYzwPfsNej7LB8+7PMGB9ldrpA36no5ujt+J
n+I2+sieaz0f7UhHLbnGb6jNTHxmIPrXLVuzm2bl2r9FxO4Ft3sFoIAKDyIJmpPm
dyuCrnmtHbdOpV5raaqX3FcfLntTMxtQP6t+E8nMG/uqeHkA6YmyQ0hpFQr4r+O5
EBJwf7qCX38MYCXGLTydRiaFaipa28WGkW3xvHNTmGgY33X32qs2/cvEVvB/tf3o
XVdWyxspO3CsSVVibmRyLQ4QLuyfFn3kvOVFeU84AhVkrAY7nVBt/WgKl+lrcD1o
kObhNlQuypp+XZwuQ2DpETZ/TAfNH2HolShltM3t+nX/t9L11K/exhADBIpyJRLc
fmUSsxACqSwlS1RUryflfj/+vNEtWpUhJ6FrzvFmRG9gl3gmwW9qzJDC3JHXPYDS
GNgA5gUJet89Nd5fbjF+2a+Ht0IV6KxWrq9i+rOORWKNugeq8CCK4BcXUCfV9QdG
1+70aMtWnNZwjbb7dmHFo/ZfZT9ZPzdfTzvJFXxL1aQsmj0FGEIKmKzI8oF6Bg18
kp/ut9t53IpInpYRxTanzoKf3mUfy6DoexHSeWE5gCiQMZsTw49pVVLKCWHnkcf4
sUpeZp+S6+VCyMk3OqUQ+F665TLE162i1H/5XG1vvUH3JRgRDT8WXfspnyMq2OEq
vohtcBLQ3l7oKLmCVGA7yNIz+JrqrwpxBVFwMkDGi2lxBsDXRowqtzBsN1crWx61
QajkgLdTTyuA6EtGCA4DRenVfSxmM6E9Pu4x/lIUl0EgTsW9v5TqsZkVZcE9oWq1
N+4gUZE6s+KxWD4um2e9Uh2nOsbRVpW7VzZha84IJHDxEroXKXA28o+4rr35mz/C
/BdW1F6JoQUzbflOTX5C0z8fsh/jBmOAEzoQ+jce4aFE44CWGpVbM7pZQ+hfjILb
Aunjyw+NYk+LtURfD/wCNIbDXhghQF0C7Gg0cgfyc43rnHUn1C7s24stk8ww61Bc
hZ6uF3IANNXplE21/xdjjn+htYxbcAugHh2rp/u5LVuVPYXJAqz5j+2bRbMm3GZH
mEWEqTSzFoa/zM9AY5WM+BB2b6pF4EdAXDdfNpDdjXlFkoAoncCHfyPbZDQiBiaP
/F0fKKp5pqn8sF36CRHBwEuINBobpx6htyhSuR3qfBcSRVPqB81UpPJsMwJrlcna
SclcZmCysZ8GqUfdmUUVXaQbxZjD7qb6Y1l3P5RyVA84u2k3B91IWM/xuaykSrSx
GhCZtO37DSOjm6zVwFO7jj8f00GZhs15GJG9GcNcRs7wYQk6IHJ+oJdVOdzC3FLO
YEyRpUB1W9FF7sUGuypWkvkOGXH2Vm8CESAnZErKvJh094FAR+V1rPDzjEQTv94R
vy1lCCwQV4Ndx0JiITEjNp9uUg4ATbHlHC8cqaF+o8BZdwweDgSDnVLvOEXz2Q7n
ECu9oC1te9cvSuSm1R+9m4iMMTVedSQEsGlMQ+4Ct0868xeHvIjO0QiDSMRY5kt1
m48g3xt5GViOMJcpro+xuU5sFrFk4pdkC4xTjH1YQ1tcWH9NGVAl5qUbMGA6AGR2
QlVLKLX3SEN11omwtH9YAIYMLUT38b+XtbLBOT6fwcAMc5ZDy6S+RRHoQe7EFy35
Oasj8e3CVW7Fgg1Lkokp352vM4cW0urYk173B99nHc8pZl592HcKTqtPPnjW4vIY
6uflnQKXdpyAEPEYTapiOPfm2gnBjokEB153F///Yq4z8pMGCiVH1IuhlpPV8iNh
BcieGZUXcUNDIY5VJvY7S95+8rSI+Hrscl/vQaxjO0e+W1IpzeBSh8ca1h83loJ8
Z08x9aieLf7wO7JSCu08keiN8G8oownpQfTkL+YmCw3gCgw03JidMnexDE8mdWNH
3brxIiexlthyYZuHEp62b+p0Nh2q3whMufLqC3fekYMehSEZfBQYYYCdsqyp92iy
5CqQOBSUWBvPqUlK020/15BwyFlRUCLdmZiu7ciThfJ7BLgq1h3Vem4HPaOtayQ/
rqYPRN1btdO2t1mc5HKoOi9YLsVXiTdwiLY7/QiMuUWA7pUZOJ4pTz+YwR1Kwfgs
nqYNPvlNSdQqc/ziWwG9DscvFD4QR5gFzNvtFDoW0RK2yokvtNtzGoSMThIOlmLG
ap6blDeG730HV7RokK+7NBmJaKs8OBqFB57ifQkdkfIxd4JgfqAso4j+HFibtxsb
V4acNpgCMdeOKX1mTPaeCOIUEGA5H+nCShjiWIKKHXhsULkVoEPrW/qEUY/kRTzQ
Aj4EpFiPuSwdGEC3DUoKu/6pnucHxWTkIsVuyLnqCpSG+mFtaXso1vJnCPZJlyuZ
YP6HGwsZWcsaTlEIqvBI3Tze/DRGOZhyJGgPJ6/6hRQ5eW0Kgggkn+Hg1n7aakqr
pQe1jK435l5VhzckQBgCHapgOA+3yeaQwdfwl0Mdhl7SvmySmDSSqeqi3zco6MO0
EF/0JUPKkGjjRiMHPQ12bZ7dUwSPDXTKPLUtsIzhjVx7m/IbzizAyjaRFQ67cwRP
wnLm2i9xuSc/dpDNM4sAnBdmBmTLlM8xJPuYKMaMwTderNiKAvt6eEeGa/cECVM0
m/boLgvI5MMeJlnOLQ+AnqsE6ISuusRfwIo6KZVJ1NES2dfiSE/WLx1JmQUPS/bN
udRK9RxCet17vCrsGl7l7rW5v7qhjcTX18vymiUBx9nnzrH9M//hx2mIIzzrPnwU
SpphHTfBGIJ3xaBniOAMullGDlCVqoCJeS+moXx4NNKBh3rysRJDlVm6ef6eIVc3
mO1wePRNK74Z+2v0mUYWOCxdCNDhLsXaQVaiFEa4MUgJZ/ZexnyY8Bryewe2qwHg
XsAicin+WTZdYc12PWG/9AP/wOyOPxpfQrJ+UB9PEgRvsCjmSAs4tFKCi9U1gdxS
qBCm9eOsOCsBgP5rIcKV+EPcCzlko6HXwKgHmIa+6C78vZKa3sBvQ3sEgsTqSLxo
7FCzItwXg1l9yORgku6hwpW+WfXktWXYTboQC2p9e2f0CEjIcgRuFP6awSmdPP9c
fzDbGqbZZubm6INh+zRT2m5NLtGOQqaNeXr/ORIcuARYb285cIWQzVjSgJecDaYy
3DTw7pfMP0P+GMMDzsd07aM2PZvolPR18Eecv7JNq3rT/IxT2+2tNbbipgkAx4UH
ZWu70yZJX+Ov00uZ9N/oZu9EbKioLKWRiJW9UXHTRN+e1kADe+DOTbTbloQxgN6Y
tUHMsICccxwSTW0fHjXRkaLYHtWYxFyX52ypdXPx5qydgy4sDs3T8Mm+I6umo+/B
WcqREK+riHfYyn2f57bUWSeAWfjGhLmz7Z2rUVdnVCRYfknPVrv/BgDvRA5j5/Ed
aD+lmxNTR2wB7KU/N5oG7CgwUWTlSCaZhbO9tGumPC2zOz4n/AxJz8w8e3XAktqc
FjaUDo9gQOYaA88vXHfNSd+WDja6Qs7KgxI9kys8ANyu2oa3xImy59xjTLmuPAFS
soSXm5oU9TayNH5kT5wYW2XfaTnStRnh9W5JBUkKLZd08shpV0w8tV3yk1H3X3DI
xkIeI5mSS38DQhFHdws+WaqtfKb8dewB9OkBSAAjNSGDMa882nDvlvT9tsr0kdE9
hsJZgXeioAf396TkwlIY45uPCzLK4ydnhewqiNyWmemZAIA574j9sGUta58tzIhH
yzfM43E8iXJijY6ew+XSR6iIDb7KtYBsKElHTpcoXOVkgcg+6z1GvCeJ8a2uOEnk
oAB0KAkZbpmOdl+rUh3xUh+BsGQ26qxDzqJZqQRyDtlKGdJHKLRDqoUz66WkogTa
OrBdU7+ruW75xPbG+vYbjA1+wUKu7NKYZcmjyZ9Pucw/iKHAR+ZtR55vL+AaRlpE
5eKWwZzgzsCmN4X+9G82OUrvzeHjbKWU6HrLnPwrRpmbveoYT8V8xCNNgqx9OhOe
akisfrRGxXS2gWy4GjUE4N+G3djntYj5brNhoAnvjKeKnbdy7R00Khbp5rpPPU9t
2+ijT4Awqnlrp9+p4LUJ36POxRKxE9BBPfyfdDVr+LYtiN+9t45eHX9VOvPZv8cY
P8haf7m4kBOofZHGOjyQo99fK5Oujc2TtCRrO7hsX763iCsli4IOmERYVRByev4/
zI9MnLnbtl7PJRrr+HGoR2WUjD+4VHXS3cFxPDvbMgZDJgI7gaMqVme6MaEPblO+
PjoTJh2Hbof7qZEoTTX0y/2TRzheELAKjZ1rGUoh/BJfNbAbfrYkFytszZDav+tG
f786NsaWVNUm4E7OBzWUzNpjbHBiinBH9guGAx+DJUtfBzbczjYMkv3kLhzbA05X
j+9vS2c+4xVMCSBLLQyCiq2TZmt8DmsUwzbAImXRiWyqrsDZdXIS8UBaF6f4sjm5
ic9ajfyLYcakRsFuAw/dBf2BnkaCKkANiHBCavDeBgX5HQTnac2lm+UIh9cqeuBg
p9m3H1qJv1b0K1DTg7LDehkxnftmMgV9P8atYSyJCuq5cHH+X4BsRCjKMsN2G7Yv
QSOYeAsfSw2Dh2kDjCy3Gp5RLNYjt8DSgHPKdOioSZqTQQW2t6TcK979Sf+bar+7
72zcuiA1YRlQ7Q7mB8xJWFPpwCafPVRT9hEP+fBLRHpBm2iseKACS74DklBHUeuj
9H/Xtn3C1a4Jnj58+CwVhfRbQNbP/VqkvrgJycscRtqbs0CZsO5U+K2pJuBxBXry
f7tn/Z5iuQAS7ibyr5pvItIC28ZvtcjZiAaZNWyqpPj3wWNYQvCuJsIbNqhdNiHo
fKVliZrIInwOx7Laz9VsFWaW2/q1gMfNP6D9bMNuueIEs+zg3QaFGXTwCVPWEPiM
1MWUf/f9yqWju/coWAAz6NQ+dOFONiDkTO3FFxlkyEo+6fy2eJyQzu6AWBPCwwoW
go1/9K/NPihExFZNg+5KbzorrpaoS/m+DwAdaNU4U2dNGQMpinfagEaNJtQ9CFLj
RmfZf6yc2MfOHVB4v9eGQ0+Q3fmz9srZcV/NxI3ubV3bloj2nwz/Ip7wRW6j2Hpc
Zbovbn4dk0eFSeGEhLYrPGPFwZfCJTyHZkaEl6wbLkRCLmvD5Axy0TKJI9rCXozx
gd60RlqRpNh5RPf3zl+B/kXRhTveDum8zUZLNLnkLHDfSfjBXrns744EUiPyDKw9
I8ZxFml9DldYLTM7Qh3IemZVElSQwKrVWdHHpzA47LFk5BWXRalp+gz+LGXjr0/J
uI3Hb1nDyJzUZwWIeDXwQNINUq2IpSSANC9MefZO7kUMv7P2GWYTu4yUHCxXFZN9
XnWhigPxLh+DXKIoO+5XkLWtyRUfLIsZ0wWAn6nPqfr/WXu21Q991uAR+kqWadjX
vp4Cnovbby66LNMHyiWbjh78neMKIK7M4dp/860SgGnFaNF6nJQDj43l0if+7JZx
XezH+W3Bp/Z73W8zygww9Hj2Jqo00Qzpp2DjbGSkje7Z4S264pqtYeSt84zCFakg
zuBIq8WPG9QI+tD7yfS5IzKPKlGQnycANsXCxlmJMmHu8nELfjEqtPr7nZFhZpuB
n4DlSL7xg4RRMFNDW29uy5WsX0tI9NxcvzgD3qV4Q4D5JGqG9rwU2U9x8hienmTX
Ef7OaavqEDbUQqOYfMj3SSPGFKxTtmRKKAhjWeb7fr7zLtKNg+VkEgEbNwZzFvul
C+RNWXD2wX0DT2iJfkqsVwApZ+dfvdLdqP2yG1hGUfJGB9K11YuemXMjvyYa6RD/
xHawNFnUxyGPyzIvo0TvYqDLIdBXuHIUn02cNMXz4I/RlPZl8fqqKuYCzv9f86LF
DqD2fdv5eO1AgHOPNc+ENYV7efwp+gb0r1HiatES4/69gSF0ulxiS6Yftt4s4u7G
mpJFLPlKhHz23LwpzGU61nOoHI4gkRhE11x43GCahxtT+w31SOlFZr/jm9dqY0pv
qkOAzwddVIxuuSq6JpAlz58znE2/PIDbqcERp7jy4ltfzTePVAkylLSkle1EGMXl
E84afB+dtda+9Eizj3mhZaig+YiHRm6LVWZKC2VvcigA5Aj8A8AQV+pZD7pIAQSL
EjtJ3xGtFhXYI60ViLBUEUlKsNhtIXvds+6r94oh0IUooCg6+sVxTj6SxdxynKBC
IT063WNtEI39wQqRwnU3v0FtoC/njMm/R1a6br6i+wFiy0BKNkwjRIYOx6MTMBux
zmcGnMQeHnkikaNMtv/CHo60fbDvEwY8iTgG0q9GD1fYf0bBVlvmTCqLHO+ctkZe
f5mWNURJ8HwNKtRvgOh/ksglqNpaJfSWwVNoin1p+vFWbwq1t6BC79vPb/GAuOgN
jJ2YNYocEuC2/TEMlMcvpiz5taGKHWt4mSiipXn+jTAIZ8mqvUoeN4J/fe7Mj6+f
su6+EFweERHXrcTIgP3OeNy5q21zb9NfeKkzEpMT8hXbHBAdBQ+Iw57H2R8prRh1
dbwIuPce+XbO7sih8bZp6rZQhpLwXEMThVEWI1mfNkqd6ZAEEgOv1+UnosMFyjG1
eeRdU6V/3bA6nq7ZvbTIjq6jSx5LRIj7sN5mi6nmYdKMHeD/AC8lK0vB6TgDgSL3
GwhnLlfQuoC2ZiV3UfZ8osn9cUg8oJj5FdA7WHhlccoxBhAjeuAot2GqaW3xZzd/
n5Vo/jBQhbUUvF9p9C0CQu7Ggcal4WXEVE5K+s45IW7rQssjZ8skOx6X13JdnvYX
7ASKvpZd29PzDmgb/b4nYhikssZDokVF4oD+DiJfasyLpJGlqUT31KL7hglBmNJd
6EnyWdZdhexLNHQyEy75bhPLwOj3gRI0e0Dk+WbqeJMjxQlEycBAel8Rj3H0FN1Q
bV571wY5q5fJVpXf9wlC1z0g22D8IFFy/7TL3onoC8KHuNwpEIIHXyvU6MzLcJiO
rlj6lYdDibCrqBYvTEKUy1wpD3VgHShKDpHK7S2dMkTRl11n4d+WUZztzBm8kJ5B
q/ndj6mjtsZ0usdPzSU4VdjYLFKuD7EOTFqA4UTlMBnfGQpDb5L1+3Gqc+sAy6SV
fiIwZFpn7STcj0I8udUsd1KNM9TG9czk+inanrI9ewLeGZ6eSu/5iNydaMqDMHyY
AvGwxLfarmadjLr2QxC8kJy5EiQgN5PhctD3virOD5akhYwxut/2bHOuuE+Srqnp
OiapSKkMDnHrZ+5JaJHk/OqJIsOQCtQiu1UiBGFYg1fW9KKjDuLbA03HDAehZTJx
J5qlomyj5zqSfFZDBhN8FT9NWEo5gQK89NK+jzl/wULoiZTizvtXvAhV3z3L9OrY
QBbfjTuEYPTrjR6BGy0GbeBTrBzvnaboskCo29Wx4bu1nqgqQPjIAJt7orc6Anxk
hdRZjK6ouSRdAxBhWyMGZ02l6k64NsyPU+uWYsbhKIQBUAt7B3UZD8R+FE/nelI9
QB9fyRVq75lXax0gdsgDdA4AtzgUK42RvzaSPbPRqpWAfPPOodf8c/Eht9/tSotN
8SqUA9TW2jA0wQY4KKD2jXMrMhOfRGRRSGRw2WrN12zvdMg77c4rU1UmxyEkeeAv
cbrvhSblUUNJvkptYEKkN6IsgYZDDMtbSlivw3EIOHOE7C3Y5TTvHF+ppIQJKBgt
laLdXDiBr4EYNXCx3o9F2pcaSXOv8ix9L1eBBKOuBC68r/fEZwEtBHASNb/YpHI5
PuUCzBUAmJbkcL5ce3S413WdY2Nv/OSXwrRDeEiv07hIEZLZRSkJl5sQhilGPrcp
LyLbia91DFzCQc3VtmnHoNSsL1y9P2H8kb3gostuQMrWOiQveqsN6gmXDnBvMcbt
oQmmGC6DrJ8Vs7OSAsyU6WTUwBU6jHZDLmpIMgwVH6j+7XY1g+1xrUVPV71BXnXW
S9kWO6dCRie/wvsCj8+vL0nd9JS3SVriegSv9BHqDNelJ7azottKbO2g+1Gz+jz/
zkcDGrLzEaG4kGNp0oFDxQ06oJ8DOOKubn/7bDZLwYIC3Gy5zYsp4nTEZv0uuKqF
O55b2LKrXeJAcjlsVq/7d4LRlOIbThsmfLCYuS4ks7BY42YSRMyHe1TwSkpfvFPb
O38YFXJ+r84RFSIpN1W6Eyx6vkMv8GtvSepkU/HQ7xx51ZjTjngYtVUx09t/HGpk
aythFify0WEgsN3BvFQRl2x5OReYWOhrX6hHZGSRk4wVdOcT5zZbGuS78mAMjawb
amDHYwdnEUobvaAdJk9izUaVlJJURxqr6BCIViq61UJaUH2Vm3urIbVj01xnmzUY
NxmsR0shNGua5IezOUogNA8oCL8ZNvH/dccMu9AeceJ97v1NejiOKiJLOHkwqoiU
E1orL26ekepoeJCEs6fF3JxKtlFxp1Vsd0GeI2okxCvpx0bYxu5WSPfzwLPeiVXs
3wiS9gzN+ONpfWGeh+qrywLwwYceNWG0EBZTGomjefub3/n5+aWblQJYbQlB8LUw
QvPzqSTzBkIMpfrd5iLLHF1d52JKSxZHT/aSNJZjL1+QA6yikEJHGXUrAwdXms+i
XjrkIpshMfYbfaO1tjFjFjAeAopt7WiaikEJmi2xEH7RRM4mZG+dYeX3GXYplHk/
35jiNAHQz4WgCqq67FfCEFRLPcP8Wt/fZCVGs7u7PVaYuXFciS3KuHFH8+knorGa
wKTrOa9bQl6JPoI2ssKjMM1xckAVCUDeNEazFtWuf76BHSzIsUp+gwnZ+oigokj3
LX1UoGgeoCeXIx4kiXGMIc300LSIbqWMCSQVKl0aFelsOXFYdpbsa3aASrgSxRAz
qQzNYdjckIsc34BOUNq1aMhynhuxI6oYhmDsC3/s5qLhjo1rRfdYRSqjsOAqjqgt
lAzsdBL0WR3jzC2kJYY7khCD4EeAZ8vlvHaK9SHisPaluobVv0opDg6IEETlrfZT
SiCVAEmNFGCKbPw7zHxIyCrELuJtwDMfRSAxlAP2GFyJPdVUBWqQP/yaL3nP47m5
VcB43dKOfZycyHpdVsCozFEPynYlosj1Pbt3QhlM6n93Hs9Zu8fZdMDqBN19U9rF
cGV2JkJYJ3B0YOiQPMROzWWdoXqKKOTubKIihsCVb04A9sivTAp9C7YsXpZMs2J9
Gfd1A2EClOXmrMa3FtoP4NBrIk4u16iHEYI3JzWJQq5dnDZhQsFg/KXM+pMttUBU
WKG0xf4FHGwgfNxeX0nYDISBDO9F841yfbWFHIwoVY7O4D8FSR4C7LFH2YmAT3z6
fEgriFlyLkENnilRUUAlG7zBft/iJSd1aUSNGpYUzV//q6FV7Mp202muUuOjZh/h
R0C6/RBQ0mP1yD/CF3kCO/JDR9Y78LqZWmByAShlWR2548GSYZzKqGawv29VG5MA
g8bjsmcfr4R53/7oEk4wyTNACnNTGr4VX9Trbfrus2q09lGiQoC8AGBG24qB89np
rzPkppZws5NRXQr+vc63KbBL4+eev+zUqWVBep/SXEDPW9tLAKYiTsGoXB1ImKgq
uvRzd0LFKlfoR1F1K1Ai6nk3ocAd0YAAhGeuvsehA4gLtvy/aYcGNGv6DeauvF/i
2Dd34Q45lB4bv9DEue9/pBZIQfA6+ty0H+GH0PYtIZ16MJYRGZ7xJe5L/bYELo7x
6dryU5zyQVWKqX2vsAK1DyLsSr0K19JTpri7CMSwDfjvJPKWhjwZeeZ8ZWunblzH
7OdZmmOnE+wvORyZBaduNrKNkzxyH9S23JO3ogpIa8nj5r3aj2OT5OyjlRtJ+VEg
TfqKYoAwW/G9LUPNkga7hxGftqsH0tU8cE69fq2qTMVM/ZPWinqHtuFLDD6z77/g
Yya2GwsNRDugKT5+eKrq80RGauZsPRxs2o7KigPIZT6vm+xAiQJAXJpXdlyzyAMW
vej8HxDBnzyXFYLL6oLECOBtrAcAVm5fB7BLiGpNHCuVuxPGHcAQVE0VLnGgo6tD
iufoxXGqYAZ8kyiaGEc0Ne4HsY9cQpMll6csafg2Ml3Q51wVtlVXQwtD96oK34jF
d7NxaIk3/zLf9g8eRDmugrBcxHSzAG4hguypYmwvm8H1AL6hNmy7jRwM72a2CRBu
FTB4K6hAc7ALyPJ003wcc3v5RMKA7VcHXoOCA5/4IiE0jSPo1Eaxh7hK6yPBh/Lo
KpmM+TDl3s8eyqc4dHa6Jd2WkE43Xp6vcpTuV6EpPoGsKBVR+LRAXn2aUQYojLwk
XAl65vRRI3E+RukrX9w7WZqn2DeH+ZUvuxZX46IJk54rLoEcaao7wdxNO4fsedCq
MHyK1okC0sJILkAzYv3k4OyswSjqNTVt8qG4/725Jn1cs0HcvAM4XadjBA9Cwlue
GHQohSvtJL0rTM/+Ga5ZIc9d+awan3UDTRa9QPsUPsUYN2B/dSXMuN28LQHGLBU1
yFN5sNY6k9nFzgTM1WDWE6JmMHfpNP557SuND7zgW/gwe8g4wm71EGyCsYNvcb+c
YRpbMEQFTaeqO8dceVuiZ2SucxXxPL7xAi6Hu4KCpJ30qB/5Al01NGnS8ja29QuG
+ViA0UHbqsdwD0D3/g6sNhl6Px4wKYz80oblHZd+Ayx94atH9OWzvUY8PzfPvAMq
AQb4OSdxqeww6mHSAEk2Qq4eZxOJN6A/0l/kITYQBLiYgNfVzubN5PcXkWvbk2MN
AuxLzwZzGJiVEs1Kv0VLc5+fJ1lAyYlWsV5v2g2Svw4ykCQB2oCzNKyUaNVH69op
IMNrHwwpHjGa3P9J0beMSQBn/cGHanioxjYne+jJPTzHZbcAZEy2L7cAGwd8UdLo
R290T7PczZXA0n/56pNgTxfPNd9RoiPNrjxlnNV5ilbFx26vnLRIqL4fpPHMek9s
YT2nWWcxHQoKnbEikmvk8SikJ1z1VgwB5F0p+ju2kXmoN7NUlTS7RTj/TprJxJ1K
m19ChlFu+1M8QfGta9xY9cA+Kl2q0Tj3BCnbBGnvusd61hawOYK4FFTrEbZ5bKO3
gwRnZIPQehsqcNJDiJTLpzP6MqBJjg7tiASurbGekD2MH4w+/hs62AJOG/UlHdzM
U1bBEfTnzswyT9bSHbrVgAsPcLzI1INDHrQRkooWfuqeqdsl/z9//be5QKGIWcHL
kp3hUbIEUMUoThi03s7WekiIOUdi5ecg/N2h17thWuoPefDNTRgvGt1zbHjfwe0d
EbvI7SbiuwqVcIrDk9kpwjHKGkf/isutTGQc8y42DTOpyuEK099mCZ6F8KuD9g0i
4hePCRBzXrT7KOBiSvfQ0Z46558Uxz55S2v6c3LjbYMb43so5uXVCOUUzzc9CnLf
FN94LYCUNM+zLYXt5JA1vNp0fIrJV2bQEQdAxS1aT8Hbx8HlEeAA7PGLBOJFAj1s
2Fzy9nSuz+d3olmpILyLNA1Vo5QGVS7y+YTL/Oq/RldL9lSXz5aodCRBHETfowzQ
emoR8jmKj8Ml2Oih9dPskKEKAEp3uvvnXT0PZMnnaXiV9rajgTTBQrB895lwAyKp
7N+G00CC6eH7G2NO9oOAQPsbXHJm9hLPz394UFfkeBwqxohV0twOkO25GIILw1oc
sMkAKu6g6YEk5F0v64+oFcKrgmsWJv3Vvk48+DMgodzZry396s/B1vJnsULEPYVK
GQJH8ncf7dfht6+voABSpuu0A0T7vTNYJnv+LaYwT1wSD8dQsDdk5JHZblZph6nt
f7xrWasurhN/bNzgNKY+rLzfC3xMsMSYHapahrRIrZLA9uGmZsIYk8/vqUBhAeS5
yoK5jNT0LG/IAbPCyOLlCCoDwHdj6FFSqZmA3/tmioOFPDbbuVNUS2yigsltuEbo
1PrrXE66XOd6+m7lhZru+GeLFTOMDF+r2cawMF+r/2ObUG381kixeUyOZTlqvL0n
bFvX7Gdv73xAwVnC2g9GZwPUXV9xoLQhPfDVv/qIKTZ20Vk4KOJ38zj+KcVEvJ7m
EPubW/MUzi3Im3YqeuP9eLLM57fnfld/PEolIVVq5WCeex9J6S0+NzP4Eaezk3G5
XAdV1JfH3uLuZG6wYWe8qCE8ULnRY3jsHO9F41NikjKRQprGwR5l5bKOr6CWYlTO
/W54KMXQ8IhHWfwZppM0aTToHpazzZg6ppbSrPW1SZADeBTvSL/FO8hJYFjkezs7
GAOAJrImSOBjdHc5scOvw6nsa+ab3sW4ofXn7h1tyZ90pcSMGejuf1fJnCivNpa8
7NPqLcqszKPsg/WldA/Zi/HV7pFq/aJlpPc22ThxwQlJNsQ3JqrhORlyaLtf+LHu
Wtyi+wpQTeYo9nk/6HT4umZglSeN4+SK6y9Hde6Oo6mVPe5rTrSBVVtbyS4AzV8b
1kDRMD4u+UV0lrKNVz3fZPCEQ5PesOfx/VuStmzu1tYvTA56ikes8BI+i/V8jQq5
J/BFDEiFY9uIyLj1dIllWan/W+hlKYLGq2tR26csRpiLD7o3HY0vegDS6gXnI7Qi
i+yst4bo9/djVgH1d2DIv1DZ4ZiOw81tflFB1Z/GZlMW1xbyhZUcZRtkb7KVCN7l
fq9Ief7wC9rm9Bv2mR1GNSmd4AIFrzaHYR6gpUC/HHkHQGVFeVMGIh4zQOolb8sZ
rhZiOhTkWO1Dcy107Ri97emuto2AS/7EhcSR/H3l1yTC2Ea41/qzZXKdYbjiJSvG
gPzZigxEni9J5JC6iB4kDynA/D/E7uhz5dALCdzVoJGCy/AfQwKI6v548qk3xunG
IH0mTBI+bieiLJJAMhNx0ILPm/rrr65HeUR6ip9rZ1o/sEiJHbhS7hCOzl37clmT
OpGrU/u7JW6VyF/nKDCF0oRP4JwRAu61fzvLWyw4OlG/dpU85YVS4EWxNVeOugW7
edOcclE+dVnydnDTVUlJkE8KaQrMFtYmcS4n/q+uz2l2SDQmunbBJvgxgiODBNdK
MhCFKVxe0GG/TV3z7T2XISwDsGmvgRs2mSYtt34f15kjwGV43jsMBCStjaG3iaQ+
c76wf4xFy4sB9myrM2QY0szLGJ2bmHhGubTUoF0buuxcPvzHTj3AX4nXc2BRuV2l
2UUMjoV9/iYrxFIz4sTfj/c1t4DXQpuQQ4c9APRiyeDSeNE+ZY6u6MolQRe5MkCW
3fvSqTIf5jAOjyqcSPXpAlI3wVr/By4YPHiO1ogZC5/HqdvcEcCZDnYW4b7vDzu6
z09wUQElzlfoHvWEyrd2PHeTS9Lz5qgCCGNal0oYk2EiEQAJGlU+rKzKuMsahyp9
nzjRxO0P0HK0taeqM7Si/uICC5UPJM5EGJXv4b7q80P7rHl+K5s+e3WNGDKgIIg9
zIWePYUFPn4DWJ9BLAEopfLFWMyv2v6556QWDDP9QvpLSnBelPTebvXIjnCiOPTl
rj3HvIuqFfURUO6fbzhDEtqu9e7ja5RiwPMJSeyOJYw66e5FqbAw6GFSGMKLWGnQ
2ahl8wTKOvrL0U+BvxL34hhxyEYjEMC2pKfIofsVaHgbI/RCqiMPSOiG/+l6nuw9
MLhmTWuWv2j3aXAFQF8bJaRobvWTXVY38BCq2GZK6oJbXtaH/grD/YDt96jvmGq6
naUsYyEc001w1JNWKrvuwmp1aET3Pjkq53fO5lhTX5S2iL6qPXwI5B18s+7XF/kQ
ECMic5DOfhZvorw/ZlAEJYN4403BhrOaQp5NTWLqjklT3ZN4jPzwvo3DM82LkBo2
tFU3IaacEFaDUDh3c7yE0fQz5gT5fS6Td8rPqj3/D2Dbqb9sDlAKvBQbJg/eQ3Sf
Z9yH7DS33gszJ7kSzO8vQ/eMmM/1DVb9sPgpFsn2G8vQ5ImYf4YJSdQIYfzbphn1
mrY3SliW7a94qK45C69AcgL+LZmOuHO7LQwHbj8NMuipnRMbHYjgv3lAMhLMR/20
StCOc7bKPGmdaGw0e22uA/G7Voc1y+7NEP0/8ueDgt/t/RCXRlo++2Q99dH4knX4
0gLyTKwPLOnCGm1AuUZYnZ1KMXUpcaSiap6u/osIfQrJVqGvr0MrZjVlN6vONcis
551dc/5Ng/sPv/sAGlUDBwTO3GoTtcpq1/uQ0ROhPAq6di+Dvd2St3JBnCTjNBji
70qLLDzYtlZzHVdVpycvP5AkJAPfLObmhGCosdJD8d7qhvr5HNjs6qPQMlDBau9a
r/nQa3kGQZVEjVe2wQgGlp/AorqbLr4r+1zlN7vLds8BXFuGSmz7kBpzAZyc5Wr1
FyaYT2N7KZk4fQLTBzhAAaF1O8plmkwmfA86fwDYNvBnhGTdxUS/mxahKCwcXyDh
D9Le8AIVm4oYmV6LAyrBFomlCrHTYGqPZ9qIQbVNNPlsbFzKPsI4A2AwJTm0Jlt+
thoEJMINxprrpavlNPekxk6Gb4PBV1jPQlYvwchSoY4XZGj8vMIrI181o4/B86zm
VFU0j7Lqjluttoh5g41sECe0X7Ivb3m8wdALyEPnusNkiyAl2/MTmNKYS0QufCNQ
edJ02K1JcerErSzCgTg7NFDl2OwkcGQ7AkpO7HIvWrDUMvQNrqwObZHEr0M34xvT
DipIUaTyqICFvvSZyo6aNmffko+kdblKvcRqk7Rdsp4pgiBMzYu207+GByrurA0j
Y8cmQQ30D/Msjzeuh0MhMRc9/EPJgBC4l/SA4qBgpxH/SUuI4qFXF3lw0IwQWLMS
NgfOCE/9DZXMzXr/s6GCWx/PCE4SHIKSETj96pIC4NbITroGpZd5YcEjy2lpTgiH
c2InU23tGrgNiaCGE0YUjJA8nFJXxKB5OZKcTEvID9fUu4fX3CSAMX0TED3dDRfB
G7JK31Y4JjmhAPtKDYp2m+VNKNZdu8AYUs/Bxxfqww6mhbcW9F0958ib0ef34SvG
6qvARUjKYybl7kP9xUpKjdwQzW7rKe21pGM5sEeyAoW+NtfdmF6ptNetT12QPLbn
XohTuM7pi/ooLYmeSdYpy3EXAjgiXB6c5B7xD48IpaQumqTMb6ziF7w0JwbBQ+mz
VYOswpXmVOeCsb6/L2e+Jfuf2Q2UhEqEFsep5hWGn6f2gbz3fzGqMfTHzQtbo6Ns
CSyUyRJZvDd/BiTng8Tz3cuXq7HXYCMWjDVuXYoLRglg6t8poMm1XHa5mYYBghjk
iGb+zEYvyRH3ZcVQj4/IXRSkTHphIXJtErRrd099NuZdqUv4SHagl5uzLUzFOo/E
DopMx5S2xELYtFoZuytCxQ3MCHZtGeIDCayFiX3HqqKq+U9NFJt0HHnk8cKqAdBe
QxewUmbV/UlX8SCr8HDKGLeYUS5DW8PSydTYVIn+0G+zrIgtjdmjk+Lk0ivt08/Y
atE+Z15mkOtnjxkY/vbgl7USsaDM+BSlpn4h+mt7r6fT7XnAfYitr+Puy/u2xW/J
RsNVXXyf61zalVPTu3LaM3qTbDQ+57jzJHe8t22N2hVSc2JpMeAD/blrN2Lx5Ya0
JfVKRDe6gXzOwhRH6gkMquLBgc6HCobOorVsMfVGlFEkT6sDpVIBX927SNdKSRes
3qpL2Hf8Tez0Mbn4WXOOxMOaInTX0f6uVfmypl2yrKRu9SnVPXr21fIThkKwh1aA
FRiOvcqTbhmhr6gXyfJufyqibFNnJgRzUspUjNT2qzvxDkJKiZ81qXf3nV6E4+hD
M9hmYv6B9l36vRUF/1eLCLJKdWoQMPno8lX/VjcLb/dw4Nm6ZnjCKLi2/w6dt1to
YrFawgC+yHfD2KzKwlQWRCwnSiSUBve5Nkm+UU97eWOjxKXUoJcNhsXeqPPJWgOk
aVuaqVYkYZHq9zLJd3zYGpKLBtRq0mDBY4PTYX4uYT0WUoyKOy1BLZHgUdZgDU90
6HJcTwWYc24QAo3S9gW/79ciRDyOQXaEYEEETNNfs4byEP85q5zR3CHr9vT5PG2w
ODkJJL7i+kHkAQRqpZzzuCTPE8NQq9AsqUyeachgb7/lFg8qEvggKN+T/iakrOAH
0jxtxx3xZ/xvWRuDjGMKVifX+EMep8Leqn2efVv1u8V4uGVHOGQy+tdmruQh5F2E
9IA+/aQn726ag3nlEHbsJq4k/6kou+YEYVE1m4g0m0MyvdizeGWZC7KcL4JEhIXe
wUpwun/vXm8BVvmItOlgBuE/AEfx5SPq0skpMEEshqoO+euFV5qn8sydx8laAtix
AT2eKbmvMbzRXPTkNJ4D0YlwjNDkvz8ZmTWkHSTwi5K46OjWBZpL1sw+wBlPKucT
6ajAGAQByfC4RPX93/4msE8VqZsOsDqCRaQEW4ruzf9dy9Q7qDJGu8ua0UySsT47
PklJPFLMeJLa94/GWkSfXbpYuQZiaswoYrn68+cyQ4jMSMO+Bp6Z8F+ZPz85Zs9X
7sbNUejwtdMwACRTPDF9SblN+TpmUZuvmguBgOb6fTx/5qNHoBp5eqQrLTlhTm/E
QtfcaYYo1oH6m6JwCkQGwaRCb22DdBvt2M4H7LXvqF18ttC9I2abF2/71C14OTVy
6ym4z9OhiCTko4ENLg3xVNtZHt/93BVh3WZZwhmT/XtXRdym174OtK0eBf++ydUb
SLad0bXtXQIJ6eH6Gn58BWvToVAx708VCUdH5HHXJezmFACB8wVrbLuSAbcw6ySI
2RI95i9PVOeTNlTU5ZowDkbkrpsU8+w2DiPdQ9je6cMBkosYwaXm2qtFAb1a510M
5l9+UsDS+bjfZQ5S6ISRW1Q/itVToPkASGrLSPG0x9yDYxRN/z7PQhGN6pNcvsQQ
YaPwFdNUxvg5VnizFx1/g3aKdYUEhtTWApKe7rQqdCsXHgR95jeG9uawqb+rhL0+
/TtrZURBmIa5eNfbfjhgFSeRzMAmPaz1x+w0xENNhQQfjvOncMAutAH0hRLHRDwQ
a5HYkFdxKLWT0N4aBYsxcLsfK/SDg/SS+poP62iwChVc71y9OZvaPe+bdSCMYhgu
A2y8v2VBOJ3aihMa/iV8/ob3PsvZGXigU4c3cn5Hlw2i58scJm+3y2fdaCrPhRyy
KpHCc2WjIl1pN0GxuW6L5COyD5TlnCebFQ7NTM/pzAyMNLMQVM4VuLd4+biQr/44
OdM04NPcZ2EqgRXF4TBvvz+4ruyWrkfsUB6oL+ZEoQ6AMF5CWQTAPJaJf1aohbGD
AeAEDX2jCFaJvFf1b2To1KUwvs8gA7zyTeME/UFYudzAjFNc5N2Gl6Tg2J1JgM9R
WNa+K3U4DQvzx0X1j5fHFOcitKKgt17H2Fd5ipkkthLcWpj5isX5QzbUXJIraklF
ecujBJW/i0MiL0tOF6sACO3O1+T4UblcDRNnyZwJoZBAaHfB61RGHOaTI+AbqBKd
P6gPfMblOq9gYg9JUV9jnYVawkM90IZMSvssJ+xOu+LeVUnxSzSCnGMie2t65GjH
OuvtFr5ANxqM6ULesvt6yLhMUjTh0bqULvdH0nnIOMnZ4hEctumqaqwRzX+5RjZA
oySlGkgKO6abQmCffrR8AW6RzhLr/kyaitSUkDU3IH+P0LWAx7AEw3FdUPWwhnAi
hp7bcWaezTAj6ynFtvE5E2prS+LXHlzUqBa+JamGryitDvtu1TW6YYJ2lRcZ+mto
eHaUiJP8KRwbumOyNKSRa1Tg5JhmyA1tkeM5UrBIjbHhe1EMWlneOiW/DKmkvKfi
uBAvG6wa+YlLEuF7BsxGmEixgnt9QsoSon6ORnG9iDTBRaURFfdN49Gai4bKfG4c
Yv4YnhaEedG6Te2DP5HIp2seNcBOXX/TX5jq5f+IW6DpO01RKNYlJEdgg/KWZH/s
rPjfuRLnPkNfjTy66vEQyFjwDf1QURxMfmPqsER63rztX82RNf1Qp5a6ycReBFnN
LVlZQGT/EPJxRGbbhJ7xljr3BW1NAzaQBsB9a3xE+5OxYUVeHs+6jIwOGd8LbN3D
0CBhsDr5hlo1eNMAP4sacWYs8HLaOYbWWDcNqGIr4zmCEHn/Gk1WCtjQl7w3UVJV
/S+dRu4QACdfkkTFi/ZHc0ilxdFDcTHScOOMG2vhMVQuzjZm4P7SFt/lJmCasOwg
XUAb0LskBN3sqYVnEQviOVxfp6c7oJ8YExcAvMZ+qqygyAUnKB5J7+U4YhFQWSEx
0GP79p5ADucA+TNwVp5d9OirPV5zAklDnp3YPt0IdlQ2vCHC4wOU/FRWlOhXpNTo
5SpN7Ibbtj6XToa5wKz+BahvmVyYeYP9Ae+IDLNEZ1nBoNdtewzrwA81BYSyUPUR
opr7b3U8W2SvnwjbJv8Eh67jmBvnqtqN6vfStaMb45+KhM7MZh90xTSZGxrmRz33
YpeV61vJ58O9o8uHPtsrnNO+GvF+LRMhNpAzwPqsnqsPJtTAolc9RJxch8VoKNyQ
/9nuK26ao8hq0HKOLD8+aS+ljNx1UjRxDsMjS1WcUvfR+ZULhaV7ZXGEexZD/909
+2ePuwROrTjlUALV4T6eGdx4h0LVvYlhA4kBv28v0dniTCjLnLpSwNq8MIneqW0a
zXe5R3tMx2adwjK+FZJbaQhtg48QRTz01eeVeF3+hW5g4HCGRkerXzb1nhZI2T+V
eYElkbnt0PYDGf9JQ4EGwzmzmS8gTqBjSuv7QFWZb5J+HEy4kgMYfYjxT0LGPOv4
XA1KmE8E5QsPAm2Mv8TAxd3QxWKgctxhHArELXJMG/yW4m0PVKtvsbORBkUe3xRU
mi/WCMBOvoNaIEP3g6wIvzSW7ugfE0gP05RTvjjJgRa9IkQjAML/sqvt/INmHRHs
MBLJP2ytOlD1tuOdSPAHfMDd/9rmXyfSIa16HcQqhN2pwC1UAqMXhhduLoCRDb7K
zwjFSmLHYqNfBXt/B7+zEyPZStYVcLjtC4YcOKL21cKAGnrkk4iA5cqtSuZBmsok
hzvgINDIL3NjOOWSWTmP2k2IFFX0jRNaFA1cnFFXI26NEqTvLm/uu4Yv6VK4cmJq
PSM6MJugzehl25CUHfJE49QBVWKgyZ8fwmv8gPyNz1ubjWMfkC/4UCMbjU6w8u38
SusmH4GmlJ48b+tZyCnDKAboyRtzBuRAmwR1Q430DzE9iiaR8aIWGRff3Av/j451
XZ40G3evvc2mF1MFdYU2ZRZfLVn5ANuunAx02gcsNX/uIGx74fLY+LNCyCsVkT2U
aFDSxibgZUy2CxpQJNBXAF606IOzw2US+pqR5Dyxc25Uz2lKr9Gs/EymIr0bKkyq
ivF6Cw8oy3tW0I0/v9K8VUTySuE6wWKI2gfFII4Hl9/61ZC5/BOgN99iwZQl3N73
Cu993TQtNxRZcpfmtSKoMmRmIAtWhaY1MwzfhutOO/v+TbNsqDDOA8htnJX16MFU
vmDpFLJvz/FZhTfJ+BgUr6adWjw+qZ5vsMiqNCXkXIiDcF8zG/xdHBsSLFePT6Hh
I80GgcZQknV2VOYtCgeI2KRXbzOM0y28ilRdHcag8CJO7OvuNOLYZhpYwgkNA/9l
xJLrDG8vqdPqLQkyjxEhnsrO2Wb4COjEoFvBxMFCVM7v8yEePSMsP0hae8IplyRM
LhL4jYc1UPHkevu3N0JvoWZ4C9aJ0Y9IdkVB4owti4jLmeaCX/JGJla69wiGzB+4
W6GehnCgCPSQjIT31B8q7deypv49n03cElwAvhJEKByCYWo3BEWVMV8nC9TADjGR
LDRUn4CvWd5EHhf3EFzf9Me1DKOAaROLkplgBJaBF+vPA6rxcQMprmSamaoBxy3x
KKpRJn1r0MBWYwPK7NrvZmaktapRY5NBCtFgsrsvHn+3Yon0FC/6mC/vojoboEY9
pd8fymaf7EQrYiVguL+Sz+YBaWnC/fuqZzAOmVYsTRTYoKK4Z35uRZ5oELuuZi8T
/6YpeTP0ahMYMt3ocPR7ajaWU5TIOEzKXLWGGsRrzZQpCnQTN6vKiMvIHinAGHAH
ckompdfz5rxlXfzzUYlf0T3sKzIszIjl4NE/jgWYFM0TBI+xgStu/ojHrv2jWCeJ
yz7Yi58XTXXqjrqBJCWZrzBb7No/v7bc/qLs/AKSS0iP5nBG7T44JFotBiriRslh
34VWgUJeSmKk+yxv9YLQDm7Ks/4p/5kPQpb/w8qCWPl+6c531wGpc7guP7fYd9a6
LLTV2G/ZTwUjgD2TdUuStXZ6WO2O1+0+vS3dMQNB4yHU+YyMY1HLwBARB+0cwIPW
nXmyV5tT8/F9usW7/j2xpfm3c+ZNqqIajH1b5Pwcva6dc9DRDKTN0Q04X+rm0Hvb
jp270FiezY/vNPoaPQ+RNgzMYBibnXwSdGwjVjmObQyPyznuPpJZPjQ+/LaJ+Vtm
/o4buHVzNIn4mce7NJ5uzIGvTc/4ZM85LBQavoPsZ/oyU+HvWdB48d1PO0GzsTJF
KKEqYPQMUIZJH4SXUEZFbOKr4o7AaHjz+Pd54AO3C/6GuEU9yXh4K36m5I3JUOeF
2nzRSHxaoUNS5TT0QdeRwrR7lTmROaizq+kb5l0Pi2f1NgpYjjiPyJwhzGd1+bqN
NqBjovhoZZ4+IKnHEZmZ5gMFri/lnjDiXUUi4fgZucbXTUsm5Y2gAr4GGWqahu73
PA5/qVmcji9UeVSLfY6IiGMr7kVBRNABpGdxNvzaPmS4mInK24ldZ/ySeGWyJxDG
yb2tGlEHk/JFXEdKohHVSeSWzK8KgwPOKxX9+PhgYgBrkJZ2mzhqRcHWMVUAYL5C
MzElsHpuH2wbMKzNISoTVsEVHOmw1NWJsrGYl7Sjv/PTEsIzSIZgY7kXOWC6Qu5+
RFAH2nttRFgOHCHv4gLqh2dRYqmqlaBpnp8iWks/ar9Ham5OeX8CK9NZySeaCccD
APh66OOoeAE3F5vFzfpyAfIWfkX7BjE0NrNLoAQqMZPMx+LuFOSYWk8ppimuaPlO
36yQuhXT/NQEFkaJ+L5R/qM6LFZjd/e5OkCaEP3aKD+p8ApPjdeULCc5orbZ20zs
uAOxEqEZy8s78cgpbvN1jccE5ex6x4dyaMUB4wnYSUcOhhv0elrSQISAQkvpcZNd
VjBVeNNtBZhR+jj5ud8yy6RPLtNm750CCFqKNthuyl8g514TcVJp6ZwS+2CPdJrJ
hF+eE10zAxB/Z/OJpxfTGMRl6/+6jQeu+kuMOC5znxHTw1qc8r6XsuIGhxuDYFq0
eXkpnDnkS5NtN3y2uB1u2QB5sgQ8P9iDDFqPyEVmF7/PT+L/0x+eQX+KYA753Ibu
HoBxI/wA06BIALf+ZkpkjoVL7DwbdDPDdC9XTkObMGnzwzWpv8S30gKnvrFwwnSu
iysjayK+szVRpNC+aDryFHL/YEhyesjf9KgsjLDonEp6eOI7q5olDjDbDCSfwYu5
ZUeYp+9ik3dKUQZZF4e3t0/u3DTskDZ+CJ3NeSSt+o7c1zb1xWdcS2pj3dwQGImZ
P3wwO45o2MLDQlmnTx/f6/w16yHJbpBb1woEtGZwa/pVK3a4av+p1JjgLrP0AVHv
eN5Pl0HQZWV8xfZXHqanV0KP04y+Zbo0FTWpRHHpYppIhoNCGqWk9eSmlh0mMd6X
cvTOy9cZpKO4Je7KWvyaGOlsfgbvi1fie0IzymtFJCnaf+TYAGg2uTXuyUwABP4C
/fT1eHG37NTztOoht5cfnXyuSbaylISCA6bPDehIWjYK9OnsXkKDKR41Hezxcln3
DYbT74EIyR+3/wUStEg/gvSJ8tQMYWtTDooGqIasOfwkrTAxlGgfSCg9iu00epg6
zcTotQO0r9Z9qWrw2uTc7luWzJKJzU83kQbpbVxe7Jr0RkG7j5Z8O98/uR+7WbFK
LcJyA8EaYSAaI+NbB/efi+iiryIWEq41jiajA29nIE5OfL+UPVmCpJsqKnKyW5Di
GC1ac/lVeAcMJDhxUupOHoXD5bAKpuPt64jIMEozfgIV5+Ij6AGaXB9xBeLCaK5/
/axs1T2uEK2JmOlaKnrQ8gs90s6QdJOJfKJzmw64OLp6B83tDyRGt+CEZu9bGmkL
buP2mFBr/4QCNxzAquhlUiacMV/xID4PwUDGRllT/7T7s9B6xBqW8YpZfkPlX4tq
k1eZ6RYBJa033tR7+bNQj4FmgG2cxyV2+b6RAhQ3QlovRtkj5idXkAgNGOTZep5j
VQWuWrad01fYyIEL4GP4NbA5FAgFS6C6r253uJQwql1kmQPI/DKPO5SeWSZWJ5Vq
swp8czi8EC+XTwM1rofPxhjrQAYpFMc3Q/PS7KlPBY97MTQg11Hm5l0/mRMZ+opj
c0R2AqqEY/fL4M9VsmRyMrdADfnRd5AMofs+oMeGRFKw1rk8pRV9KK+HjZmWdWkc
Yul3roEiSr9/qoC8ZI2o/bTaCnp69VE9WPv9kdTCvGDpg+xqxfKwUXoBzi5ipGaF
jSO3AqnJd/cT1hd/5m3zU4iJnW63QFhkSC4CZOQLVXsATkFzAMO5lK2coX7L6YU7
T4TRplvpAs2XlgJbN+e+7p6402Fr1BEcq+j9DgECj5Kk8v5jj6Z8EkdgsJFIW/jU
duIbX9jmU4tXRw6BdvOhh4Ho4Oa4AWOaFjn+jXuSWcwpV+jvA4mgOyRGvvByITIz
ZcUdD1YpsMdWevaPukf3NEyw2aabpMhxj6YNu7hskQ4pMWu+eQ6b8llHtI9JBW8L
SbW8nJCcuoicNFGgQO1yKxVPIcAqiU1LUJs777JwwqLkuWQTg/OT4rhTgl6DJpzY
37sbd6JVmDcBg2eLhNevx0Nq06eUvTKdIE1qWC4tM0IMWbACZ2gfrmm3EFeBAQ5i
R39ZhOqqLruRbVaeGCVdEmQe2Cj2QNy7VfO4M2Qcw1j6z+SIaIXDdCgtT6SQjYRg
ZBXAkPdkKM0mVKd5Quuae7ajZf4RaYwcS0SrZOsOAjhuHs/JEvuCi1ecKPdVr7dx
a+K8r6Jr3RcYGXXGMcU/FuUbfQlvfPvf5zVJhavFGk/oCRcZ7hj7/iwTbumG90XE
HJ6anpZ6lr+Yi/KQ0QZWk34VVCvkYPvIqRmrP6OoAjgk1d6vDgLQcbYPYxfeF8c4
rKzVoDIB2D2lF6nW54BkmH2MLu19b2ZqVNAIBRXkjz6lYxlSBtRffmUQ46+zc4KT
uP9s2FRjpTJMaoBd9MFMBjAIdg5TS9cXHhjVd4BBEhpWhiz1Myx4qHI/FncwsoHw
fw0UMrwy6FWjph5HZ9hqkj1YW06XA3VBBaeWg2/3ug+TxJo1/lgac3hTkpqbqymt
Fhs9sAuBHHratEsgfRHNqU6rY0RtrgPWxWzGQsfokB0Cb7Hf3ggXzzD1yuqZprrg
/axNNJbng+AoG2UK8dXnyQ8v81QPXL8p5xznJTyEcjsi5GBQnhMyMQVGGQNuP8G5
bP0upwkrkDZtsecZ8t+yWz/gmSkOwe//aY3EAO9T4qNIJ5dcwyuKSMFlT1mMX/3d
hgdxvjiT2ZLT5skgNqU0/p5784ejOzQrVo3bMfQSiZVll8FdBbkj6a5l4SX9y8Yg
jK2paythNtG4FjX4gWWm4oPH8sk6LZfC0UkCKgFWDTHBfGV5BqbBrlPgntU6TRhX
Kc7n0dOorOVXdPfxeVdM4RWILRjRCRbm/ropfN8JTq1k+YVhjKGmty6XWX2j72O9
czX2Jwco/YeglyVy7JepeSJ4jqCysj/XDyghGHilWCh0ZiRAKZXUynsjSML06gSG
NUiybgPFfEURoE91xF/3c/8kU2I7IQFv/uIZE1noKBbG5gVDxptEmxKWXgK5exdB
V8ztnqrSE2guEI9whSV5q8Gv4azg4Ik3epogZ8RWaegtNSg//uxwrpQ+3/Sb0+f9
i2Kw70o+W8ghRw2ZnAQgpewNYW06+1zcoIk4Vr19Lt7Vnf/NgpMjD9vGLbfeyNNo
n374jvWKH1fQy4K//m1izndB5enmDJChaO1HT7XnXdW73kkdDgqGQTN5x5C2GGPc
peX5NJjK28uwDzZbuMwLkUgu8bIeB2CruFWsiiCfPfwm0XAT8khfYLfpoXJCXdcY
D43hXsP2aoAliPJdw2qZu81IxS1kbcYFTKfoxGmLNXrCP6QRrmIZulgAw97O2VYR
a7y+3BnAfzdZszWGFEaOm3mH+fHzjs9bvduqbxSD9/Men/ai9rQvvwE4ykAfrewb
BRo+Y9Zk1VbjKVHuDHUUDl4LOOgirNJSI6pYNq/bIeHFmSNtOcL0wabz/IktG39d
cPCYt2Sz0U2y3i6BlWGbyEpBf4wHSua+G7fezItTaX15taLKqCQZvYE8CM48tRio
E8gFsZWaUY2N4dqXzuDZTZWLHP/muPqPKDLOb1W0l+jnPVnRLaKLcjJedGU/zFpm
qMimLeKT95Zbiu14wSdkKylSNfebs7a7PGmSMEcWRRS/79dqWpHhA14tRfPkb1u6
7ag4mDdmhPxzeLiU+LC6JRfs8j++OrJBUtp/cryttK8W6DL/5d2zim8HCWvZZYe0
np5mBJisAhLuDYCqGDGqNvyr1r4bdoogaOTIla25UDeHxwmhDlwpBEcKRJ8XKnVF
XvcKoQ8DzKeH1bMIjpgcwMLfddU1nluz0BQLBOAsTl7Xiv8cx8Bufh7KvMDAxyiD
4W4D1QJcpaxiMOqHCKnWCKqeDUhSqQYabWFB4ENP/KWvAfzY887HM7TyfSXHErKo
ItL9QqU61WFSbxJpd/R5vj02QO+ok2TwWoPicCv6xZuPOUjU4LMdfkDPgXn7puNq
PwRq4+BhHDWBdU9ViSOtm2JKa6E2+URl0ZY8STQWeSYFbMpjrwfIx80BfL7SPSxq
ii/FbMcbfMhOGHRvknbSdFNVYgMo95JqXkBqqHGWIsGkEzHYALG1cEDpPsyzkHJV
w4xzlBPQ4Px2qwWm+93u4sQUWcvWipMYHxHT7JkyWruyXxftTkL2k99eq9PvAIPg
e80nwQ+qchBwkGg7yNd/qsPFc71OJwCB6hOE5eE8+pSr3+IkN3m+AdccxJtGFniG
qmVqUtAo6jFhLPGovnVopDBdOaaeYtx7w0geM7viIaIVMHFbsMwp7GWDWo2r27Jd
xEad/oyknjiQkN2WZOoS6haYkmkTI80HhRgekUyYs//DgM27vweTQSM+b02unpcM
pqX3R2yCusGN82AlS4S54zMyGgyARpQoYVwvbBnziE3zF/fH+q8ygMkhKvfuDq2k
jMK/vrrQQRHlvvzLRbhq4V16w7mMYJGEneJRHr5yJ+7Z9kNGgpx3ze1KzEkuAZkC
ITGgR49Cb/mhhBzU++Q96YPWLYDFcY1JdG9vfmxSaPGvZ/UJ2X3YTq0r6Po5zyO6
SSvUnw5FrBZ92FYDBmL2eGnRT02r7Ls7K7WBkFhI2pGKHSnwlX7WXpviZ+HTeChM
IzbbSa1fb4S/FXfLZw9ASGVr34RYBQKb/X8DlDnvvM37IUwLSnED0TdJVc98bpih
pkUBBepnJzzHuUgQyRVBGiiJpoOnjgoHVVb9F3PQbNeqD5dSvXV09bzEqkm3wT1J
ghRMmuoqsYXTX/Tvw0lbRgFtU6MTGJeykGYB4s8EMoDytwwAb607RfEaCxFVmWpC
Ibg5O3AHXAscwzFhdvfm49ZLQrub+6Rm6N5UWTCxcRb1PPAOqlS+rAOo473ehAoO
a/GcWEyrf3f8EJBpQY19PRASSQ0DpqW/eaAtaH97fvfqCBQp6Atn3k5q3mcrtrQJ
QY0qCHMbFn5sUOWB5BEi+Pl64g0VHsLPjq2tqU6NMXYCdJCYjUH+hpwbJRjuOoqw
SmstuUaHuigaXkOXnICa8PQhHHbboAVy8UHj3cHRY8ECeE4IbWKInch1Y8LwnZor
/NiA8GhIpUo1SO84IRm8ZWNhpeg4nnWNm82kglozE9HGvRhwENykb+HMcZezVcsn
qXqAzLiuXD3nNiDlB0fCAUvyuevU6EoNGwktE8ZJs+N89vTFv7FBHa+XL3TMc3vD
iznq+EOiWj9BO6GcAZZyXJm3T8mVOJ/wqXitsGiiPMZNU73bT/gSyBn1B2BHdO70
qPkCLilc06ltgJJIdgGKbRAOD0MYU9x2GP7yKQgaRPiTFZpd8TGUF9wisCG2mZDj
PdnuGTMIxemI9qwkaI+GIHC995w9qDAcXlqS8tfv3S3P/37VKLyodVBq01pqU6ae
ltC2AGUL7ka53WoL8Ay0UkKcJwojaQuf1ERHLUj3epqEq05wURaenxzpxUrlDG2z
aWv7ed+Ws8sP1dob7AbazyJeXnJ7DSoXvWR/BgT16W5nOLKxafWRQ0pCgBOd6JkC
EEG0ggBVdOgcYoqVUkNpJcEfvDerNrhZth+NI1D50YUr8JEKLW/A3PryJyFdpIXm
uRUIubECJkBkRlw7PliK/TAYnXCltdOrJRARw8Hf91VBc5ty2lzsW5LAkYp22LV3
OZTUTWL4olAP9Vu6QHo2GzZHkDb0EO1Gx2Hxpfwm5aOetO8vNSTFLZmj19tPRetZ
A3xCrgt8EY3rf8GKbKSy6nzned/bugI/8gUJlFs3nJWwqGEsSj862kgmbsKFRHEm
FFHy4T9lDPfaOlsUukpr1ubEeSNDqhG3M9bjCtbSFwhmZmUSlCcmdHX9aPHNk51n
pAGHOJI5ZHboijWwNv9SxPaZn0cMN7nGHnkQB/9ff/A7fKMl+yljbUA6x7dGnXJp
54hcxCBeaFza5tz6IIjIUtkSS8D88/pAqNjKIkRvOYUMbWFAFViJDdsVI066nsbr
Iu9OUrsE1iB3PJHNoTzjjB5lqB+NSQYhqmmDiRr3fjO6jh2Sn5RID/OPF4//3bCV
tqhyDUB/s8CT1GOZAJnSe7HGhPtl2znv3kNAsopdAcFFoyekvm64AfQxcqT0nURP
dd4hKuhro1Ng6OVaa6IkhclDS0uz44lDBmEkkbIAcJH+8BNewAqJR5QxOh6UONNd
aCtEZXYJnjM1g5dv4c7jCCP4FXR5aqDIYu1lmMZwifTqNvO1FUlHidNE/KOQU/2U
x6hx8egxa+pBMQb1NtFf3j7SyeH4S3Xhn2hdmVAoIuTa6/eXX7sKVJDxYFZCUWmQ
Y+rMywyrsP18O+eP4Lc/PIFcVX7xGwqBaVn3xDQsilI9I9bn/OW8Ss+LsfRrUI8I
XaMTq/m/gQyWCbVYA3Yd6pYxEoeDA0QBpzFtfDZP5HlCS65vZoFULyzVRf0RMjQw
z7RzYJonvbqjK5xcxC09IYd80JkegQC70EiHyfikykkQolzaZ7pifVS86jttjfjk
Younin204leyEBv7oH6Uv15iuFvt0KjGJ9IWfaWqAHIIFPOU2QLGrvBiiuBeNX59
BGtZxdeN0uiWTTbW4Z0bShct6PCPq9hICMKnYIR+tzH4dpC997YcFqYP5DsWdq+M
+dspgaAf+qnPrhxfKDjbJvMIPU071NUwLgmQbV9RTijnEGi6hzw+xwoDjImboyNR
c1hgina112AQHS6cY0meBgFvZocQxEmoCzHPlFqWi565OwaGIJR8OaNpFfXcjjL8
xJrq3O/tZj3L/jxcmBQ7xmda6rv0rLrPmpHhz+Ffzoq8EW1hS/ziZmUEi41I8zxl
Eij66G/Tws588VO39pcPgWFj9suY8UXyeJGyJCMgCRLqSKAQO2DviYewAkn+tbhd
zo8GWhrBoDR+rUuJ2dCozQVm64cfOqdPrypeCMWvGwxv1Of7nnCnMharvFiY4tTo
FeGLa0XaE1SdpPJSGB6Wkbu3nOjEqOaHgx4SknUA+BLtVk0TJr0ZrU2JVg37vfIC
/5clbN+Iu0Px+bs/WFVqadP17VWut0+amyDC/jabKuv1oEkok3gpXLPYG5gMA+jJ
M4cw9qYfAcxW67eAVIJlps95mb8IPQpFngzKZxgHmk/US7PweiCJTD3976H9XH3l
Sd2HI9KUdsYzR7nIIA4J10K/dIUFfdz2F4CdJAUS5y07QAThuPy4AhHslySGzOb8
vwOOeghPEKKxE5rfE/7jLZKY+BIbOBKR9dgbyxb1/ApPFJT7EeImv9E1Q+XeDbK6
OnvtFbgbzOtkPppZF7HuC3coO0ca6HzlOJ1rb2eiBNQKV9ly73ZKtjhHK4MhULkL
4j/ML837NhEKfP7oxWQUbv3OlNJyj7BpxGxSq9nPTSPIxLNgIPBfmBfs74nPFGU0
Gc6L5IFSXqxaaKe1zq5MuYxFQMJs+v8/yrq6LCen/XDgu6+vCC+etF2zor+F9Tm+
09g6ebM6lzp/MvVNobx7t4g+hLFhsmxLrZLYVqK9F/a6G3GV+Xvw5J4ZaURb3ZAJ
9oyJrR+vL5nkSG61lRE84TAoDYd8H13663SjPGSGRr/RUP7JLLeO+brNvsce1qa4
rw1+wzMUlIpHVYDPZD0QvFq4td7Krez172bKebLgdhOoJ3t0j9FfH6n2mLGch6Vf
XS6itettHF8PAdluADeOxHgc9EAYbcUSmnQa9Sa10FE07NkCQNZlvSNq9u6ZE1AR
6rgsFnkyzcEmJenVCHDXVYUSA6h29D51jFD5rOfUq9GsacvB8QymVj3rFEQiYsFn
1a1NrwmBndpd0gV7z9wCFwDk/K4Z8djM7Us8v78u3jgKAOQOAvVjt5UByQ47loKx
eM+BU2O74wWhDNA8pZXUJ5MesXxJMRtZpdh9KtewFVgc+Ae3vJllMEXOCLxVNHyV
CKNluD9OFRfPoFtTYKYWC+6PS3aSFosEAL7gW2ESVY8XYSNLrQ4C+lrPx3kPWAYH
CwE3uFREwj0Lj8SYuWaHamITu3RCufJ3HNTH9nDZugr3PsNVWs8HK6A00QTEXuCD
E4LLYi/Z+jGPSk3SJMptBPDYrxuAuuQu00soP1rcNLJRz9tQI/PwcGC1ZrcKa126
1/Z850n9+Sxtg9zwEiPCAxzFHixrBW8alCD0cD7qZQOrtzraLpJ/S6vPtol8PzOb
bgZ294MSOFsFQgVGc9tiexABDFQGxKZ0i7bOVtArkbRTHZZUnwk3TuwBNZx8NndS
+GLy0KxkmSR/ZZgxQzDNz/TuLb0HeQZwe7OrPntZCf65vS6fCo+tVPdiN/+9duV3
g6awJT4OepK6eemB8c5UfLzjgeo1DoI8F8RZEybSN02baklx8TlWCxdPX74rWjto
m4UTyJf8D1f1xc9YHGpIHj7iB85/PiQN1D9hgOFa/mh45BLTveGlGlavHegTg0+b
PIEjQCdGsBEKMEw/A+3aynH+mhwx3bHrbDT/b9EGGNyuKxpQk1RjLJWqx0+0fU9h
99cO0qGcIRrnUGLgo3OEG8l57ja4Y8k/b9w40IgRAOttKe0D2iFhF5JFBX/Yf89o
RGQsiF8Qt3mfjg1b3O3WH69hjEfKwuXB/MebYZ6ewdfzz5K5uLj3bGCuTRLEHlTP
r9ZS/6688Kz1cvbuM2iEwHav2Ev9OdyDBHh98l6CdmM9+1YnJznbe+DfK5ZIUAax
KtiYBGcwEHLU2lHzWaLdqsMGY1aaYt1tBo7KWDZ/YjD0fbzib4+JQ7nxMQRwaS3i
2S0vrXe5CeXr9lOoqNdbdcL/52WcNcb3NQ5v+8OfpsTK/zxTB2IGT5na5A3kGL+S
sBvTXNW2x64b0xw/4s4D6CqoxCp7tBcSOgtqerThbK3sJsVe0JlMRN5AgHFsJvgj
V1SvGkBNc/fzlEEwdNp2rzFFkt6MWvodWVt487Xwbly7cs9/TQQrsHcUh5Vx+3Ox
el1gpFs98yL2rz/wQdHqqCmIxGG3x3yXozhjXMX90IZNDbmop0zmV5AsHx9DilS0
Waht0ahcRMTSoOsCCoWPxpYDICMKY6DoLUJK8AvLHI0pFjXgZqToSo5j7uYjEn2G
qOdBPQKzsN8itBOFOnZD1La6QH9lSLY/lzyvI7EbSAt7IsJTntWTtDizj0PlYTD6
rDPl/+pRDKEB9MDpy5BUk4Xc5ijJpE3cS+BEoV5g42B6M2qqi23bsKj7mx31QfbG
z5tTbiHdZQuP7+B2p04kMe2G1t8r6BSgtw+apOe8s+8JWQf7tZJCTb7uYk9C37AK
jo1dyozugmDFGuN9PMV11HwKjYCqz1a21F5lzyaDKDsM3nmnWcGa1VHIBhf+dy+u
1h1VQlVEgKADDxDILoa/uDCKr9ikeerHUKsW0dVn8hF8Kqw84QPndZLMCQIoqQ8/
38APk1maOavwgXmWnFT8NQ0sqLoJTleneKs7LAm1UMmvsjrdynoNMy4KGGeG/G0d
Hpn11dULo5TEe8RK7baUCgA/zUXy7zDrLPsXZ4gEfdjox68c2vPzg9mfpuo+pqtP
gLvUcO3SxFkWVgQM1J6lz/Nc6vp8yJ/408/feWkcPDdZDAyO/sgN7bbNyaM1jVhs
d1Ci2BUJWqH1nQvAXL9yUVHnczLgkLaP6byL2UTaF6yr/ubO6B5lsaJqxprNyyUl
Yvm3YL+sAzN20n35gqoEkyjOQzdmaZ+R/JBXWeNwNKXr3Q90ozlcob0Y+IV46qt4
cQBmZp57CgF53vW/egwSaS71HAyCJHedPOJc0K/9QUT0DZDNyPXuOQ+P0ki9tS69
37UYJ0Uo2aBDAo4QzCU3Mt+O4gV1LrqASvjKTEXEmv6MpmPUJNjoQpJucdpcvB0g
i36890THiRdiNjOzlCeSg8okgeAZBCdrf2iuHQzUOw7BCBMm21jm18nLlpeftyjk
gN2xnNPj0Mgs3lZeEG663mdnNtsrE0wNsZOQ9Ca7k1EGgBg1TaHwCouq+ZKzljQ6
sQEmR0HbcG7FVfCdYhUoSfsG7MpP7oGlAek0l5wfcilMDjQ3o5JG9Gf+eUDGexSm
1at6nLLzmJI71ZBB3q7UrokZe9T2sbJFyoXVGUL4LRaw+oJxXnaBU2xA4+W6/2As
c2o+yLM86SflWVCeUgFYr1NeLB3uo8baEca7TTzYkwtgs2IL/nr0YlRsqJ62jdnG
5dZfKewNXblhDtLhobymJreIUNfagOfY4ZdcnM6RBk7myZo3p5TH0M6ZJk8Ld0Zn
pF65f1Uq6xZAKWkMfsHnSrEhw3GcOTvCxfYv8aeKul9hCj530x7Nt7Nv6bpvR96h
RPRfgb+u2n9OZjU6OiE95AqOTPt8o/ra226oPb+uPSZzGtksWNmv3I/oEizR1DQn
WzE+GLZgRs7HAmfEnHoY8zL/v1TtUhfpmZw+8XqxLJbsmm6T5VjUQHDoXNGdFhE4
s+YUBVLCywFYwwHeroP8mArKO7YYnvHS7bUNlsq7k3ZezVmaWw/nnx4TW1AiHzvb
/VjFcVrpQ1qotkklNafTuKTE2pEGHPeheS0IN8f8s7lQrijbICp/I3ehTumfCfF2
6Q799mo0MCBjdU7Cr9blNrOv/DpFWbAy2kOJFHWGIjceX+mPkhd888i8li7EwCmH
kRmtzjF8/+Jus78RvXk4G0eEKEI6EW8Vq5V2Eha+CWOlORiIKoU0dlIwS+Z1Qljc
HG9CIH584XwRilLAjQNuQP69sP5+nhcSwZ3ze/A167GqHDqaxRfjQnw1r2IzYIcM
i+AkGTdTPLduGeaFBARRvyI3GSRJZA88+CPXJSrKo9WAWjfCjLI1SbyctwOo0xrL
QyIpTiRGBQDLLvHgs821vL/v9Gppn58eYWXfyJ3TV9W3d9IAYZV744MnI05FyI2k
jdVdvrTG8y5A+cUqMJQOhe3I+pkLfsjxSudc43CJU3TMiyTk8iLxLXORj4/T8nsT
8e04EE42lTc12xr3wwlauWdUhWJTx287aXKCHTzm31+yxevwtsAm+DkUFcoRkVf9
nnuibBELCIYE7MZly2WS31B4FeWQWQUEih1tR4RbbsIttr6DORxS6PmGOYcd2Fuk
VuwoX2zvdIp+bxGh4nW0hwxHN6KqO/qhf3fH6He5MrUE+WAl3rXwLvYdhesFzb3z
FE7JcwyeA5lnpeQ80iyx7OCA/HoB+eBMz8qIbH/z0e8Pd59OnIdE7WKnnnfkL5NB
Uu8R5JMZKOH3MbvMaR1FkzE9h6iSULh1pZgXUzDH4DJ1V8fVGqN9+q6KRc+uIWu+
E86b0PPeW8/FsUaPiFopCsjsdnG35sGs1Z/LmnitnOu+7w+EAaJlhSjmaBZfRDaI
X/ofE96YKvQF78ATOC3+8E+loa3Gcl84HHnCTGchnEZNRK9RYkNe7mIlqZ24DPti
O5frawa3YAyyVH+62MXoLlkk3L1hmIv2RqPCyNJJ1T38RSK2+6YgDyoidXzu2NNg
ZytqgkGCfPxVzAGhjP7OcQsnB6XepJV+PLuAUZT/BHhBqVz0eYKwnNrTmYATi2hI
tKFhBHHD3HMNTtaY0cI/8e7IFP3O6Y+n6FtoVCj5DxNuOm1V8EASOjxxrRIQgAa3
pZjMnJgYEu0ydsHWHY92dlt/uJMw0juJpbf5+LHCb8Tw3FBcUJIf358dXMZUmuIC
IzUIWRQi4HHpLY6IYThcx/4Wtao6AD1ubosBm89sczJyKcMoWvHgeEMIRB1YdUl2
KYw23FfpnMeWzcP8jlI9s6K9M2bXDRw6+ZTsBIwEUR9Uj3yf3keNJiWYER8elOfp
+ntZHu85mc2ESmPBTF5AGo2HGjSVDGnmWNqKWSevypyp3bltOxuolPMRfcw516BL
nRZBZpCfFznfG6WvJM0tNlx3VXEymZYfNgZWEMP9fkpdPdroUAI9ngxg2sMsmfmJ
Rnzn1Xl288681EgJDJAjpzCE/z0Kbx1COMn3grcv5ODSivQOJOo9NI6BhSewvot7
vK0CeVE9Oa9AWbmWtlWKZtU1xhhilSvYtycB60uyu2No+laicq+MUR19FUB/WTNL
Xx4aMNCA3/LVE25GByqmnb9f0f2uzlidH0Xfv8/jrvwcdy+S8xgQei2EsKboss0Z
C04OekcZdCgjgx/WyX6yy89hZTjxunaT2Sh7MYMXrcMx1CrIJA7T26GHnVNYEmss
30B3CdWzZzVIC8Y1KdRY5+6g4ux6CNXmauPNm5iXuuOGwc6ennESFpkLzzdxc5cG
5SETyYPn9O2lcKB0YK3u4e9Aakb+/1Sgf+0SRnpBQd5gQrPeT9ZB+0i4x5pA1E6I
wojB/6b5tvpI6MUBXW+ud9xSmDR4mlRlsgsF2YznVKEyGbWyR/ATgtTxPfbnJay2
jOhCouQcF2oCb93qqbXv3iEmYIiN8EKpPWUlitjdt/kkmPH9pwRQ0EUXlxFG50rG
kB3i81MolXiLm9kky6frz4kzD1DpA9aV++glI7nUL3SpCrH0yBYGvhcHab9EzSHB
dJZEw0GtRYsOpiIOB1kpFkvCAXixbxdxz1ep9GGFibIj+U26Sv/s/QyxEHQQeeFS
oDgAzN9+IFl6iiGWDAcbc48GfnIy7ow0/hBgFZ9N4zgwT3/yLJzYHmVFIBcmGKPq
T1Re19H4J8PjLJ169z1Tz2fOwTdhNWbt1sSBvQxjUOMPK1hTMWfV8IOpTLG0dUN3
Q9TP1anu3ORxqBkXhPPEarObhF2T8HYxT45MjEBGEIl+THopipIMLyoW/Qijwinl
sNlunzd6jq/03DrB6QCwbiMUE3qFohm6zkwtTQ1Iqi4kFuexraKolXghym4+pddr
7jZwQX/71FfrACSHsB6w+GVeKS3pwdg4DlUGMyrShTd2EmlRuJ+Z6DCNmIPvDr6L
Fjx/GWp7NKu5mKia/5EB5n0JS73KwuTAyMHLTjfxrewWSPOD/bwObF9UB+xOoyTJ
OeAVaMHnnbYoqX/BcKU/SHLbHr1hy8gu1vmoRGgELDaB5TP5HqbDjtSe3Xzr5hup
VfFJWeJAkn9K6rT/mf0PB64VGb1+Cv+GUvRbIUIouQT3YE0D6QrwdQ6Qa5koop/9
zbgDqZRQAzjLSlwPDMaZuatXwlI7nvGb47S5nRmOBfwX5oW71jKY5CavfHCgm+z8
Lmp1ZQkDjp8m+8W2pZhLszKjW9TInOmh1Wi1tNG4rUh705rx2KEM4LG6WzooTKbO
pEkWfIwN2o8HwTeDYIv7s5o/0jwmRjYdweibCDxaap1erJx+ItrbOpV9ja6d7sgp
oqNzZmpxxd0WiDWHE86ci8tuqJQS6LoLvV6WBBAU38vAuPFCqm7J4Jc7wzXHIJ6Z
05zJfQKRmQYtUZcjcAIdkXV5ZksgkckSTvBSSdVrEL1ibjLu5izPNCHT6VgSZ5fK
Kd4Ru8w76WhLavK5qaCMsNLwITIHUY1APGhZFdAOU6t2Cn1ugyqpUDt/Ar6NiP1h
Y2hT2T1jAc7QSaTRqX3Y2j96sY5tyBTSPpxbLYI9TYaV2pdQT0m3uuj4/x6q5kfZ
UBEzHaTNlyiwwsOG6W09rwyDpi3YNCL5P3KGFLJXxacGn/D7mYrEWT1DYJz5yM5J
EK5EmIr8Zs4mxKJDvh87SF9+igC2VvK4Cz6wV3SveEmgeDdod48BQc+J1uLJc0fG
pJiPh1CY0gpaiHvJrf/B+r0+OBBPswDV+WYZemtV26hUtD3zYN8QVdJW3Jgxi2jB
5f2x8OapmPxQPtyqzrL4+D3xS40DxvkNWKVugFQ9BqopnxwGPq6347PYywhVjSFH
LQ5O2FHG4aVIyKCg5tgV5vuu3jJ8qHytYACQYgLSZ88+QhMSpPR1PxpwUyYymUoF
21NlGrsrD/i9tvlNfCm9nyFcqqwoDywnW3Q24cwD5pMCyuNmi+PLs7QfDz9KMysk
iaHezJl6Sa3dDKvo7vdFZZHFs3OcXAfzQgCpMtdH0Ftdmr+ttTbDaR+L0Zf0N5Kx
HahVQK04OLrqjxGwc2GtVAkZqx/DhiswvkguWgt29YOta18Ra41XPjzDxEbDR08C
GeL+LlCo+tgavObwo7WmFhRTbpLZjSYPj9if+OCVhzQyIL2qqFq2wSteQpYrOjle
i1yzL3fxPs9i1EDV9o5uR1pGJvWQjTmnFaCOlbF7y3iO8BryC/1YSb2aCL/ITBwz
p8Csh0wedl8HBDYW4hBQgJeuN4wGsVnRuS8SB1kJwAwSVgsIIG5rUdV+eLmWsKK9
KZ/Puvt3W3gj3qgYTSiWWDFxsXmf49X3J1Et053TlmwqqBjzIrxASKBNVCNTelRf
pKGp53NVFeNQcf9gcBqCjVFSUIgNq5kS5YQ1qB94fq5W8wbJTo+RwAUpEWAExIY5
ZMqI6heMZqCwE/x+gD/i/g0G5ypJhTGZkq17M4KS0CUNS7UROnHp7mvYPLIsZvbF
DaVyhGBypned4H2N8Sgnkc5s/z54fx9t+kNxOWQ9nkUwXRXtpK/L4CuIooK6qOEi
/F03lR6cz4S28NzdEG1ZX892af5PFdn6lQEFiK7RmeKi8raFMz5/CTrrdt7uieTq
4NB1BO09q8MAld9+jWm5vCJp055WukoI1bKViznt9BGC0lR8KBl9bSCXayEN0Xm2
OUpPIwxcCOADzNtudpkUyk34NIW+87S8mb2zDC7+ecBGES/r/MuT2DY2JmAUOFav
J4h0MbNpYZixa1etSdSGEYtj49tI5drduu3yipmJWOGg8R4h97qefChmnguypSBz
RqU6xIKinbnNrTJvzT++w1fK8wehp67Uwrq87t+n1K2alQlENu+swda+0De3WWSo
EflP1G9/pPKFWubBE2U6usAU2rgtR99Sm4nkALIEEi1ZzD8m6ny2WIgLtHDw16y9
qSxi4KxoFDkenAC11fNsQEgx0KTYxYoDPadhQCDetmJXxfGbxYkgyFJwvqTWImqH
5JSyhKen3eYlnFWi7FOpy6sK2fdnACIU1cqGVJKcl8GAjWM7dveNDWu+SWqWT++8
/S0RkYmiuR0/oAs29Pw66YwiKePI4Flk+9w/7PEXvqP2MWCBttg2hixgLfTmbhIE
nOKEos5ySNtDs3DC0NsuijOAPYzuZntg2gMqjNCvEQr8D/6SPEvnhFZLSkLkaqF/
OvyZv4b9v6nsfzNDZx33juIrTuZdSq/pQBWl66flB6iPp7JyAHyKSk/mwD+biTIk
Tu9huSXStZGXa2FcDvVjRwfkXCQAZ5APXhbsZj2IeKCpkrJY/z3XZ62gZ+F1ddyM
/7MeYsCG0hW+JLTLE7fhBTM8d4piE95EATK7jBrTkzriKpep10HVULBvhhj3WBHl
rjP7PF+xUoT4lmK0MTBmXEBHjIdcvPqjmRXb1K5HvtIEZgiGUKXJUuddcrVfvKCi
m5q6JQk/f5I3w6tSEbQJWfX4Wp1tS7soflGhKsL+3W5l0H2HQaVxLSpixeS1A/Sm
wi1ZmQJ5eK2rWtAq1qenNyVt48zbjtvqn9J+W6opE9Ul8MVN0iVQQFoXMvrJyU0u
toRyekE9+hLON8fbv4j2VsregfJRrNYrGNpUeauQZUwUz0IcVE9hYg1Tyuo+Pe79
oIWzPmoA7LNQoPwEDSvB8KLowWpElBWARmzrRQaa/9ExNuRlAYgKIOK+rtVO2e9/
l6cO5FkNfAZVia91MpqFcp3PFGSmabDy+lZhlJ/6yht137YGb/V7Qur3/qRX24WU
s4nnQMV4q1R78DRjSlY4ngyE/czaquvtm8qvBhlF/8Nk5IhEd729rlMym2EI0h20
95vftP7AtIfiLle4FKivW1NqntCqBx2koiK+KeE4Eg6+T/Yp4r/G7dQp22xEF8jr
6PRVe9Kt4OOCDy80M1gxFxxLW520qyxCTOLSSJjrI6hueiRGbQrVV9+FHDyAAK65
w2ify01RLvvMf1z6V0ltY13yrHBychmiUMwuvlSAOF4G3UxI2zznAaf+8106rhS8
lhZJFN/9bhIJwq0zo1QLsVOK/tWwZ71ch8R4koPgMTGOSwtMxF5a+Mp93zGJSAjr
Cg4c4sUvWshI5YNct70QCFGMKuX5dqRCIgWRqx+RPcLZapaCABDgXHfLm3TLeVZ7
8yCAdHVadCiI2ZleE0+xjLO+rYtY9tpyAg3jgIYcTxFLjayPAd/D2DWn163nEnBK
aX12259dzLyczKx6TtFJHwlBc1Efip7tj1vlTza3f0iZACwgyueDhsQaBbzD3yNU
HoqwzyhzfUc6l1/C9x5xEB+JI2C9ndGFUxXBreO2L2Mme+L24bIm6fv283KZyZqv
W1qRexhLkaGGpeMCdvHAehIiOTjZKgurBh+zDZmaEDJOso1cbu2oJPffrJreEftN
J9uKui6w6+XhqLKOrTWtfdkmA+QVqJNqpGgpFY31XxMMBLcrZEU3Knh3QNx1dc57
xaiWuK1Diera2XN8RQTUdDPjSB3gw6JYjUsvyVd3yHvlFtTMEOjg/zrKfWuY2w3E
yd6CcG9Z7xwDkBvEVpxcC4YX5cKO82O2y/0UTP6WvKC+31iaYl2Wl/xPdzez3pev
e7eIm8707fpQo6OJfq7YUNPbqApMsBPYc93MYRG1qfESHucM7/mGByPWLJMb0N3R
1n1XrY/nFExZxTWnDf2+LWGmjpVGPyOfv/fIJmVtnr6PM9bFXWLlCi1Kva1fKevv
B0MLEgG9c7nrtn3NtQQjaXDHYyFg9e27CRIfrNtrannD3WBMq9+Xxtlvx2AKBgbi
DzMpez4SgZoWZiAO6MwsY7BV5JBS2eerFWkmkJQ+rXQhT8+Rh6N65I+RURMmtoFr
nW+nmTW/XXkbLgUpFu5Dok4wjmULOzrGmkvMnDBNb3XQ0EZkL/6R9Si7hSgdrXGQ
37vxPKLN7L5v4V8E7ovh1bJ6Q4vvGAnunxiWG6NjFuocUosk1Td/3EK202ZMEAOW
ijwdB4DOLwX4pNA+KoVjgpR/Hg2QVl426+ABhIPc8n8GI+eM0Lytkv/4A37Ufzjy
+ZqaW2Lw2W4kyDlgo7XQO7c9jqj7+vjc1fXIVGj5t+Bf/V9B5ks3KDokuqez5Zea
iEJxUVfAmjR/CxB20DefL113XThH4uPlq8kccudydFkykmVUgZm7m6wyU1p9nDwl
2EgEnwCvW145YUUV4TsA4VL8EGNn0KfJece3shNGxUg40LWzI5r0EOFxvhd75ao9
A/YCyXdVLdOL8dWixw26tXyxclCs0QpUc6kHDwAjLU2CN5TWH/uoEeWys3QfYZgC
5LdytsRBVp7w4Bgk4rl2/Qdb9Aq3jKGkIaj7se4ol772ahE8NDm56nj2d7DqTeJb
6Bs5yZ1otlnwZ3H/lPN1ZOEW6dcA2OIUijaSYYocVEcYLaiy+MhQyH/z668/etze
od1Wva4jKjj6QLMtxUNLgvEw+GUKHzZ3yX2eNUlqXQQMZgNAAHtNHP8+OJYi+14E
SAuZqPKDIzB/ZIPbR7m3O1gQ2xEEOh6xsQcmxi+jAkFgV2iSzk+RDnb453G8B8o5
Z3T75cKK2dtgQiXTCJAZE+sVWon+nAIoQgZKC8cUmsTdNTQ1PFnzbXx25rQnq0xD
w9RDxApISu14z6H4q8KqHZ2D91EwG3tLatcnzK+VeAsmREGMkEDBdqSto09guimo
gmzb8/yfklFLjGU45U/0fwvlB+Xoo2M5NWOjOYdcTr5TLD8cxRLqZumXotk9BD6O
rdYfYR96zBNRXkfyZO5fy3Hi3w6+R59P6tbSERUgewI+aR4YZIo9iFVyEaAuf0Mh
HCLw5YRpxEuFsVqtccjzeXBXhlGBmiy6Gnnqms1HiS53vMRPKSarkBPrkVF2GBR7
kKaDr6+GZ+P7rOS24V5AXRsln+NkeGo4Hgv/YCcoOyeFunErpuxYkiZ/P4clWFQn
j71wmN+J0B6VrUi55xqLt0X0X/1UQYDZegPoMXDcSrT+MIN2NS/EianTuynFWV6B
2yy7CW4Z3Pe2+4BUH/U/EjmSo6DHptWqoO01gJ1ZCOvzOS0qN4odaa7rVM6ErZL1
ykzzdX4uxTsFKJfKNAKeRWy97f69xepZgK8VOPv0Z+POAPhkFSbk5luoRWr8SXZi
HGh/7o02c9Itw0a4AE7KU5/0txz25KlyIzXjWF/Tta2SaHIZw+rYZddq/+ITqjF0
6ab2E7gbApXi9uD9Z+mg0Xc0YvTxCsGuXB89vlNqyZEnAgbvPMdy78YlvVG95AoX
oy/e8Q6qDmKSEW6LKfMCmQjrr3pAin6cdDb+8F7CQg5uZOx9VhsGnlSCGOUDFMH9
z+HX+gEedYgJRzgll+Lc5yZZayG7656hsmxGR4lDL6DtHIdu/CF9LuaYus/S9OJH
XubsSCsHSqIbRpk094Zbp9YfQtdLNVmNZm4v+kOpNpPGzURvu8pYjwh67EXZDAdj
gB0u7N8Pa0q7bWmA99aJabwTiaOi76QhbovNR9JNJeDDET4eBT1F9fmSzCMjn9Xd
QcIuqFrY4PHgzI2nKVjRx85e6HuSX8AO30PiRBmUO/6HcNiu7zAmeQjKWi//A9Eo
YuzCAZGmms148Kok/Qx7pSCsnFRpmst9T0xaI7M1Jtzd2yoJBqoBySmeAw/ZHDif
GmCIBcH3A5XFZA+beF8gL6B+NTo/Ondh0V5LfR0YB78kbG/6SZ0EibEd4KoX5bcp
4bzoz3sj90+sua1twcouDHfWbEP5kd7292I/xWq7EVNW2zyewmsh+7/1CoJjVjGF
ePW5a8ZBvDxJ4htHtseeCbL4BanlNUA4pFEJpBHvVDwzH2kN2h7PpbJJpIJP84aD
aOCTEDxCdFe7M5Ez6UJTNQnh0TnnziqWQ0Gvk+YacwMbxdhh5F0u3y9NwVrOrWiS
vMiPMRhKRA0OdYXaCjQDt7JGy8hQhbKm6RXKf9GO1VPKB1uc1MDXV9+asSJqukPS
/waVbhScOLc9qv1I0jChibtBmcY6GY9G0+t3WnIUGdt8W6Q0xx92DafqAL4g33Kr
MEa4x7AOr9MtkSYsgn+NBZEk0gMIzClnu0je1mZG3BmOFjeeVcCr//1459vrG1dQ
ujQm6T4wnadjNQUow9NpCfJJubP66cU9p2mmkS7LqfzQFW4ONmLR4gD/p+GEAMDT
d3r7GEiEBmOlVyvw4pAgpPIGDufs3aVu+fPCWglP3Du2xueygUCYnj1Cpe+cf2M2
EGR6hnCyhZJZtVPfMtpkK08UJEWtPVbgN5aUFUHgzMxs7VA9+QAbaaPWlqzF60In
6RPfB8whdJYYza1mCtCwL3s5yssAal38I1kfAH7xgksw2MsydFRczp0hGU5coZS6
tADP/I8WLbznOucU8bydEfxldCOFD5c5qKjCUrFmjvrSvuuHnktFSJXmNX4HdGDL
yoP92TMuCmD8LGf5oO3wpHKMaHcPamlciWCyS7/VtlehV+VWypnpiMFMVwTCg3j5
xaTeVTi0PnpD5LsJAYoIfd601xIN+ce+Af6XhWpN+71Yt5S3rj/fiVCzm3MWqUAR
qTu8Nv+E5AqPA/q8NKRQEAkU8PznZcK7dcY6v7EzNaKcRZS3LrZg4MYHYfQrZNMp
xZOcOV3XsEewJ/vkx/4urjenMUe3ChYi6oOhucDnUwukJvP4sKdO+fZSEkrUNJae
Qw0dahe5+U0HPV6iCul2Hg38lwk1jDgw7R53qJ/qzxcoHX2ALxvdoaQ7Z4LAOeHO
677tKzarxvos/WZUJ/h7+7HlIfeafTRyrSQJG14hUy0fA04s6CI17CJ8eByzS3zs
qoIM9tQ3+Dgy52GTxr/LdJfsJcTJZM3ecwAOeKKk5Sicaceb+4riwjx8QsxDwpBP
1LTYL+PFoGKQuhppX5p0xWeIHMhrKU2bovK21ChvMczrmxOs+4+tnykw+uHWQzWE
Htauoq1S68gJH+IQqNpZvLkBK/uRlilBiknOBR4x/pctlLbkuHR8dObGOfKREoeS
GIr5d2WLHbT9vZQnrfkxmP2cRd8RTx0Xz4VM7ZIpUkYDd9gTyw9bKccI6Nk5pz3F
Mgs8N5xH+rX0s8IaHHW/gRbG8o58+waTwb5lYkg1sUDgARWjKxW2GCCk4ODsypSP
Hqt4uHfF8/giL6DHN9ZESPFnOd27k4EBO3zzwrjLQE3EUoKELi74HabfYetqdxqM
+kf85ztWu7ELbzEpET22MgalqzdiB9p4pIaz2yelYIpuCdN3KcMKMdUYtepDE6Ef
P3h9Uskd5/o9vztzULo4mv0F87SGHWi1Hf3NoAD3Y8d36YDxYqI79bUnqNE31Dt9
6cLS0d7E4FwYEzA3GUo2cnPlfExjL3m3RIXCI1XIZOdEkeSEWtx9Y9ER6t2k4LFs
R2MyYljQdHxgvq7lmxzp7WylELRAo7iDq3Yb1PmpI8ebpIdercZJSrTIkEk83EYP
16on92vcjSZQ8KhGY1c5Lf7snGAursGzQCz8xy4BZY7/52CuPBtkpXO8ofX7B9LB
aDuKqGkDsGKEXRnrH5Ut6OXpp6qGJpP6sqWWbk3nUFC8aRrW3l7GtqjlQKswrhuf
Ys+Ku1TSaHjBQxIs619T993Ukq5KEsGw4Oow72arAE0M4kN79ntTemiB6mXJSiUE
pLm2Mvk4OZ6o6YH2xRn0BXkNWdTPKvTxzG+m+P56sU8C8g9/fnuY5t3qzjxnRXBu
X1sYHidHIaMlbHd7FA6+V4GCwEedDO18qAaL2LlwTKqTHMEhV6UjceYOr5E3cvkw
2PMeHwhtCTaA/snN/wGnhRJiE/3Tgs4tmxEKzeVNDrbvJdRxnKnsYtrhB711P15w
0atDw+WFnr3cKRaB6LQns6/++JL2TWJjPIjZrs05yvxHolba6dCNMzBtB3og1lt/
k5vB61R94IE8uAJ4iAcTm47u/4Iwk+nE5n74XiJzKCwRSu2YN03O/Q2BfdcNjo5i
JfLD7ZtHy234HcdytkFE7pAhSvUd7ldoASD9IzGOyR4PYxaEVPQONzNtqhLbiIM+
IfUmCWWJbBt0l1i36/YDcnGQjx2fYGnDzYEkTqxWSkfeJAzQl6po2f3QEIsYdN60
yJvUfXA1rk7rBY2ovfX+5Ob5r178+m8UrZMvt0CAqJ8qIJhm/p5toQ3Di9IyJiFE
SxULjIAiNt1cpxcskYE4+yu/m8MftAXhZgoAAzX1sKyO1WksRxlCpxaUwAl+AmT/
877H718yCggEhTCTxQTiqJHwq5H08KE/3gFOwpiuXLnXqJWEJGIWgaQfgdXvrGam
FHyYUPxPh8wHJRWt++U7ssp6LPFme5eLZtEf2HDu0hI0Ozu9P4ugTT41mc2XeSMW
IsTRYwlhIO80SH0MsH5IjvJWNVXh9cn1GenhO43WjOkddssHPnIfWhJ+trqs1sWU
JJQ/kkAvYGbZaPyO5N3b1O0cyKtrupNZWDswG2U+vIuf1fhHWZ6OW1Jsc8RFRDff
t7Fr/gBH8JSRXed2BwMK43Pfc8VXXGnDtaV5owD2jbya98vJdgCLlEzeaPOutu4I
vZt+gFRjHOzSFd3kB9C2iFURK/Pn5s9xll2MtjeJVmalUNbLHex65uxfYTBEyiQN
ci2aSCVEFNwN91Xg/rZe3N2h6gbYaPGHzruCuccZizf/mEHEkQ1PH4WlsH/4chIQ
F0HLsm31fjMmHnyg0fUwOdcn5dQKSY2benF3by5T3bx3tDsVrNDBEEu+peleQD7z
2FEcPm1gdEYpZ24VYq2j5iVZtutI62p29p/Ch/hm+vFm4sFZYDQozMlosHkJg/N8
elrNAfjq7KUgr95zgAvv9tC3WOa0Akq8Cq4yRZlVpX6l/0v/xQ4eydOI0loOjWRj
F4Gke+qmC6vTqUkvjvqDK/L/+SrIluWe/FTOf+ledk5Z+it4zQuNvJGPTdcLEjBl
41tH8kdh/OGF6WBfJRe6yraTdZZizmjx3iJMHDw6YWOCp/EbUOpCgAAlS8VoT681
BryvqV90SjK0z8Xd6K+3acK1PinOsq49zEN4+M3yuXZpM4zAJbwWWqDJH3ML7u5s
yu86QEXQYsBvHvuhdotksCD73kjPXMREIRvQwS7qG+o2z9hHe8s3VEathNuBkv0p
QNOJltCEdO3QZzNP532D+05O4JbeL1SHUZCQNjFypYQXtmerP6/S226tc4oimuT9
EOcv9tRIp9XkSmG/TvlxPwyJ0fiLeuAOpirECbBRpHRyzrd3iQYwgA93SiQ+JFAC
DMEhj1wbRliMqGv6rcN9YKZOcTRUtczjhjR6AvKtypiIiywcY3YqMUESScG7Elz1
daXT3jqV7V83CYkAKr/4Sm4BubEI4xlWOOFc5+jwH19Jcq8w2MRkJ2X9Xf3Lsib3
SLpNd9g/MzdprB+R1gh6JFaD1wfJJm/ui6pdxMifrCyBK1xYpgdqu3me0ggGvs4A
wuBQVFC7W9vIzSfNyQbwLJxvJ2UA+orOY+SGXj6G5PYFKRUfJ5HiWHZkuof7sbaj
j32RBomFhyW8AmrXS0KSIIWY3h3iIpssY9Z1gloI/6YxwFAou5AI+qC6AOLIITnC
PKB+TbYZSur/CplwmAEb2B1jVuumFw2vnrf2RI9dxpT9lXfc+rV1nXC5ZVRWQgVX
UmwfVWpzrxyuI4AbsgoR1lNaPU0aG9qf4+Pht32824+YdXP96eiJq++qJ+GRGI1c
AzeHhgRk4OKoTx9FowtJy+aiEOGkTPfHxS/bvBOZ4bKL82TZ5XkvuBaRS2y0IF6c
mrojT3lJsFMRy+f0kB5We6P69jYld2ud1oTngywAi6uUymnBISfX4HaOrcnaqu7P
Zs3NmCPKSn7HoWv/S9X6FTx4hRQ9srKS2JqWFdy1lUPGY6W+ovj6WtXL+TQHiCMr
w6UhUkHFVJWH4WYXvWM6oMx0kI0qDKCtPtSWa/7JoSwqFZhWVnE7tK088AmZFZ/d
44acbYC/hYtwhVuNlC1htVGN0OLl+fseqV4mnyQYZzmnEip9HakHkdSegvpedVdv
6dfU8iBtypbvuKetiME/wonR2X5op5zsmr+oKpniQPalOvxnM0VICj+Gps/7h68u
+HG3zR61pB4oHi0iVH8d4+42kBYFhqAqp0iO/MoWT1QOD8x1ShdComjVavaVwesd
HFM6h8yiehrn2PTENE6J5E2ysqCP0ynAq445SejeXQHHeIhDeHjoMwxmv6UQS/yb
RTsO24NLB4UGrpq/FD6OielInC/2Ujyz7cRP6w8UWDsdebqbwPRDm2Ale4t5FwPj
+kTv1L5BjuZiSG4JvHmjx4I7Awxhm71LYG0CHUMKGYhSpOPl2wCTAMCdnM9LLYj4
AqNJlP4PKGaGDu8+qxn9QHVoId+1yWxanoS76/bAGx31ycI2mTgfNgn6leZ0p2rY
rj841pdA3o3E+RIMzQnvmRrCN01bC7nCDbYwmzi/rN28LIIytaW/sh6wkH7c57iy
17DFv9f52sDRUW0gzqlWDMo6lyC/Hemf/ZyQKwqfzhlyMveqj/nC/yH3u0r+S91K
O52/toiWwCix9rvC60F3pP455mIZj0ecnGAQeV8azPXCx9Hxw0M2lFCP1tRXdQxA
LzUQypAPY0nj9GKI9lOnNf+/dG2vxD4AKBOtzocgNixqrO4cgQlbw8FAcsW088EE
Hd3cniTpZQvcMX37rw0Rmrjmium1ia1aKG6f2PF5CQkYBBm9NVrcp2IaCehGmqtI
9x1vztk6Wzl+cWDKti7UALDYxpRh9kGiS8/qLpYD/hJnzSoiJ0P7a7Q/EAMdFv0K
DCj0Xlg8b/Rfji/+EO2AkUC5kXulw5qAzJH36X5GTlY3fRJp07SLn3d7gkictxO7
dRL3nLibV424ixhWalJ4pCsfHdGPO1iVJtcS0+Zna/NwKoSYbDt6EhAcXhbhf7ni
lg3u54NyW1tssukiGU3ZkeUqDBrMs8TnqIDs6alUVoAdx+qztud63KN6jFoS5aBx
3YWRrVsh3Q/NQjoy8tzU/dLWh+0/Z5Pm1bR8yatY//LSY2cDLrHi+4U4gXpw9ljg
VHAmxBYcwYKt+McdO4qu4bBdK9klj16S3s3Gozdfo3UcD58fF0Wub1ecJlqbmyXs
xMQnb+Yz/C9mtrY9P6mmNglYHnFQNyQh1CEk0eX4dfYa+xA8ecQp65Ed8uvXxam8
S9IwxNR0/Ex/z1/7qqy4E7E9sJR3m/slMPkmxCWmk1haPoXJ5yyH6/ngfu1FD2f9
E9sRk1L4K0MS9/5ONlb8eepUSgRati2LrQRvMmhsBA9Wl3JpFC0n2RBfAxBMu3v2
pjRHToa7ox86H6jbqKUU6GRbwJcRE23l4yJi6emKLKqszg658Q7zx4Hel+kSHxdh
Y6p35UcePlWZxjOS2uroSpR76TLAaV0vLASMOuV+EeSKjkQ9tIQ4vAWumcMewoTr
VTsWeBuSBsRHC8trDFsaNe/6EVMn/gZwbqyW7k5PuLJnm9cRyHDdirh3o5TtEu6B
Pi2fIuaoG4tUeMQi5zAfMxefO7WpeVqaBZaXKcSxW0/HVVBN3RAzgyFPpXPWmoPF
CyumYj1E6h1ChdKGuRNrCbklFV5L+Axs2o6hRrDiUJBx6x+v4euIVlL/WNMKDGYW
CoUH0AdA8LJ4urbFWn7gYV2rrVwCCnBJXvTJLmCXcSFpy6CZ1D9Z8W/tAryIGoRd
Z9KzpxETYwk047D4bRdi+4PIwOJyzLSEUximRjhMU/UeRII2Pk9My543WivwjwvL
MBxLyVPFvfU8iuNtmIVlpapwrLXYAVliBbQVEv2Ti09+8Q1IuFZZ4TaOOmCUIZAI
2ABYu15habKuUx7Ut2vm/gVZm+vVajRzZ86HikatVqCUtQC5a/RCXaF36rG+LPjt
UXgFRVsZPFxW0EnccKkKBwlHJmgzg9h9aHVmNF2k/6buxYP0eXv0ROhKOU0SPeFW
4QFheZ3AW41TGFIY3uNRKO71obLuwIgbq7DRG4mkkkTwaljlT5QiLqDiNxHrpXPF
4kHixI2a2rfSKghY1pURD7L0kEvMOQFphLkFmb66iQIwnzCvStgCcs2My5WFegge
qzSZ0Won1VbjHtSv8c5qjEpXQp3sR9ZWko3OmMHigMDomalobzENNbcc2Phwasam
DHtsdz5/SMrtdAZGhi1U9tnwXknt5Tk+91WM70Fnp69pFw2R7qX3EADgJxOxJ2JA
g7OreChF3nwgWdT6v1TdKlDRfVPNluC2x4Af6fHgdxxAMXUHbp9Wu2Hdjv9lLjx1
q5Bd7U0DjklMayCxVyv5xTHxLNAZIHCYzESah4+Xl8zbRM7L6E2SClAg2RwAbSKg
Dajw0SVF7AWwzwpKGqQ9zoo0SzrxzGx0JFTBQ0iVHrSmmrEEOj6vnjmijfidaExe
4eAhDOuEL+Arc7uV5/p4MzSq80oXS6o5Ul8Mr1XKCSowJxYRcb3A571Hh/Hnap+S
xuBq5qxhqN92CcCXKRMGrovllo4ou46un9FkbrZSXZT0Giz8TUL6913Aj125B1lM
vKOdvOEjeHyy/X8INs3Zmo7UE3ZGbkMoJoIYA3385nK/ww64Uv7Lc/7kAQkJs59T
gf/bXbaWGTi8v6BIXkDhnjcI4xGSxQ+OSVJ9mDDqRMIU/JCrUn6qZS79aB5uj8at
7+EPnL+7/Y40IagHHMK9P3MsD6QOTTb8Dyb30wtSL/ytjEokwoWCBzo9futCCrl3
ai0Q5OQiXuyRs7UEb1dBk0xtyrOC8gr0Z1TAiqBaIAmn7VSSALvIZVdOp4ceEEIw
SU8sc472dPT0nMqOPWISm3KCLibsWfqqXUJ9TS8679rivjBNH/9L9TiI4HMHooU3
UVnNF0r44nMuRySEEJwbc0iTIBEHymRCI+AY8jiQpUqVwU0u7ysU0sa1zeGBAX5R
0hRiPdTtw54mL2723lyqvIDIWG4Vzpsu/0YZbzSRwj2DM3/0ffRzaC7uD2J2lhHb
IyLxJ50OSUwCgbrKYSmJuQK0WgONJ+ik7OX7ty+Yt/5WyaLNIxkQeFwwfgF8GYSe
VmeW3NsD8TmCnZPMF3OFm5nnummOEITv24Y2tHSsIYgd99BeI2rPrV+gYCns0WsU
Z+89XYc8kMpNBISCJDF7tmSxPml/USpI5zSLdkGiqkJSqiBnGanDqgidQsSrQSch
eEWAThSA+wCEZTmkW5bCj7RsU1ZMXFOkymxDr6Vyt7zNWMR3KJZpkbyhKWuD0gZH
kSPjxMpJZ9wnptUTbJpF8XYsGIfVZmrBcjh/V9kXVAazGTjHcfmQZYjWxSiw5Xnu
vFicZYyB5nbIfO9oQY1wjyQeRE0dO/crKVNRd7RhYwL/tZtSi+xmDdlH62Y3h7qO
chDpv8tH47tRbsuERhEP8bWyLdFMdSG61xtguZA5u1dEIOLtxW1YpQUDL0cBeb3h
8gJ+S/Lw9fE+t4+qIOqLXH/Bh549p7dubMTxFhnOOyD+1gN+0R2/u64wsWIY2Jzz
dAFowv6dqPorClyPfFcmzSbh2pbStSXKrF0YlfCdf7ArMo89iNKSMujr+TQEGZ5d
UoCbKy52gcJ35S0VbUaSpKwt3JD0QTAnaU0NlPjbQLcZ+hHE8pWF8j+CEunPGOxa
ddKD3VRQfZGdiKsW+UqNGqpIPr9k7iUfSomSiMZXMbA5bxfnMycEY10/965pg4lU
JlkWD4YalFFFYoen7cmOgwBoZya/feeZBauWWzGRX/rT904DHt7JzosTeWFCAof3
uAGAMqaKzG6EceNJtsybai9nxGlDtbi5Vvw98lpAfLKOF+qQIl9Qv2tGDD7j4UUZ
7iKaOTl/L3XKfslbnkUQ/Zcy1S1dM5geBR+2ewV/0l4RFjP7GydcRe9iLHwTu2R2
yZX0p7Mrd2I7KUmxlQfsGeBJ8j2U3djamTWsZlDGmUn2kJk4eF79W+MS2n62AZaq
KPRPuHYd3fqwAl4f4wT0dJhoAhW0QWUknkQYwFMu0btVC6tPlrBz8gB2S4zkRMgK
+n78ZPZ2KFjiU/qzg75mZjwYgN+YI8gIMMBFD07BgHy9MLn3p9HNUiD9DfjvPr54
pTs+Xhj2u8WaWUtyccFD6QwLSOng0AAXioq0NXpwnB4AS7R4FBbx8dZLyNmoyeFU
gyQAgs5qomaHnVEhXItn0Ag+AQPYbE8bZbs+OAaAqHsvi/As6CXjbd5meKUg+4VU
4ajVKMRheXrYAmRKLS+0TPsP/zF6DgEnDVeT2jHzUZJ4IoS0AOQ72HB0qeH+Y09T
+FQCAOyPjSziMmvFn1SamARD6CKo0A1Va6vEatSTzGPxqfpgMvsTRI+wXi0xHyMP
0CnRoozp+6S6HnCKaBA5BO2Grmz2RbEZUs/VvSxgC63u34cEeVuZsa7ZoPdy69bb
REEyyIpiRFGq4gdsFAK+hjBy6Zo9ruYq8NjhDjGGdfZXdHJCI7uIOWmqriQSSTbR
FiMIQKn776Urx44XK9qSijyxrW8xvpXMEtG+srMgb/nFEpf6JqOlymCfGkh+6LrT
xXvJcf5BoLl3wO5L0dCvYPlfvIu2fmdozqHJuBb++TOIUQQWEt1ZvYCj5640NK0n
JAbDwIBkGWo5KEYAivON9t6qPZFM+61lIwT8ZwikNL6nlNnDurkAPVixkz/fvCER
e6vG8tyyh4LC37Ms5QZCCGEbGmzk+Bmikz3DHdk1R0vYHAjvTWQZ62ujoHo8kiEL
Iuo9gxOWR0C0bbFxE1sgWYfU0JpijjB/t7blpnBSD7EDOhHQxOqkWgg7pstF95TZ
q2kl88bT7aH2Bokbjf8knw8tV5h7Xj4SJ+L6OeTabxgho9sTnVTUo41ZxHwOY5Wh
JUPG/2d+JdNh3u7I3mAVAIuSH63w3AQNC8jOB2OnZpOjd87BKVGhW0KRNNTwkH/t
5PNViZSPjqb1be9rvmUBS4KIvJ/EBWQgkV6cUgzh/DSYmIeWJx/4ldQ9lymi2woY
9IjV2S1XbvAGrr0rGXxnpRxwqnRj7zh2vosECmW8AnlPU7n4CHkd8ktkN3AML4+Q
dwLtOolDGvLNu7AjG8P52KI9AdkNh0MNIx6DE1URULrgJ2XJKaO3DitFLBi6zZat
dH4GLoK1Ftu7HWF2tjDKhOFDiNsNbygkBMj0v0nC3yxzYCTeTL3PJf28GZYot3Xp
nr6NruogtOwjKtCEwim2Xms22zcICr5JRnxaydt82kNv+uuu5YiQMz+fx17kxmc0
PboOKgXaxEvgVuYn+8CI/t3B6Z9l7VYPg3Z9XuUocbpCSVtlS0UEDRnQqZEJ7xdF
YeOwbASf6YClG/kFcjjpatbKw78Karyr784IpMmpyzwUKVIHiaiyqWuAW4aWl0IU
ZxlRj09joR5vkRJmgd0HnSAExyhJpbKs/xemnFrUzMRACPlPBbf0jnxoN0SKNi82
4xC+XVfyCrmRDZw4g4BYShjbeWGr+t0aXAmjXoAoXGePweanaPCUEwE+k5QDcdmx
rQ5QQcU/xXG4idoijnJ7QwrtQox63wBvyhpNdzhzXN6o8o44ZVNLyqa9iDBzbqmk
j7TmX38MOdXmyHXxq97KtwzjTCGsxgXX8zXTwTxGGJFaHqc5RUnt5Wavlhw9vORN
/H0AiHywR/7nySGbZHLZnSTeI3IEcFGTeYkK1uBHZsjkCDgYYFlbDa2WNSwV8kJM
N8cx8ZuKhTwSpfkQcukI9VVdszTpm1TvrkMqf8vM/QKJO1nxUAVBsOyXe+ovRCKT
lXH8Q4RwWl5eFo9M82rnr7mUVM4de9xGz6eDhc8bV+Ihpl3Fnc3Ema2aCHstBj2u
XMO69ac5xwBxrjyy/XV2kQtdjgD8z4czHLak22Rq8VA2+X2wcIhB6Jm3hRR364el
VGQ0C6dRpUuk5uHGEbrzDZI/X5LD1kz6irn8/t/kSE2lIEt2+vnsT5+j0RG0plI+
di+KMqq1hxOdzZLFPuqmiqooQBMoSX2b0HWgygjo7o9AHfGWu6L0b+iA//mvz/ce
jhN3OLmCxSIB2U6ndFtCcpVh54Sk5pCwUXPcMDhwqhVbb46+7OXqBerETjXnLtqS
EUzqSnGZE5GBi+c32SUHI1S2ZVSkcPoqfyTus0up8gUblayCTL37NFYuVtJK0k0g
SWuNjuxOUETCwnlrqqnv/RxtNJhIKMaTIiXBQqQs43cy/UE/jdFJNnTCUrOBaVUb
PxmpoPCh/UGxGYXiqfGlZ8ACs5w7hOHy/YG68QW8+KQPpPRncXtYV9F6Imh6WPEH
HoVz9zucnv5uxwwq0Dn+OLcWALCBimWgkT/d3jiNMJjKiFn4AJegzO4wRPsdYrKY
JarxMT1COeRW4PCe8/tfh8AwV0knKz+slaGYdRyMoBeYrgMT6sDnMERduIFPLuuV
8deu5BzAzRVYtNlxNO2uJIYjXQTAgDUT1Xt7OEva6qGlPU9WODczmMe/xNQ3Ct9M
TMHPiPm6b3wLJk2s+vVsziXq78+5He25nsvGPzwy9tQRHUwC/CGmJgnWUMNrMltS
RTaQ7FHyMpRLi8GkDbRkW/J3wC+9i5GaSxYw0QlqbTf5s8bgkZ1YVQNQ6lBRVCSa
OpRlYEiTSO0Utlh2CwtV93IcUJoLoUXk6a6U4R4SeKPLRREt4cpGtg5Nkj3utnBI
KAoljCLU6AWZrSJ0iIeFvUbXvEd+kitZEjOgVCGHWp5O8XCHyZJ2L9mU4YGjpP5r
SUO9k7LRnzZinoLMVxEDdIkAZrX4PacwP+vMlAzVqPxvnmP3sosZ0QKvzuDFiHMD
Eg5djytolHwDbbhSbhQehIslyhfBACQ/C00iJOrS0OS+YiHfx/CzwGVNYWXUga8r
07izHC6CTSc4bGjC3JwFmRdcJUYEXT5fWvDwli6DnHRpLt6odAyYOPuwFn+7w6hJ
06Gdo0gX99VlDcPXpPkpFDCf6YWs6iECpOLP4M2hmC9nAV+zrJ16rjOg6oStSkf8
adtlDzDCijLAlZdTx8DIzgxHei2HXJdBQSIEr5Y4XeTORPeNospnlaAc+EfQxABr
iZWEG9+hCUDtC/zzgX9ibygPAOw0PALcItZyN9qedt4L1C/uoQC7uJh28vy2Iuwg
Z/E9h6NRYmokeVxGj/0RkED9IwzMbPXnUMuRUKZ15rr6RBYMiCBFD5cCz1keAJBd
P0Vv/WJkfEtANYnLFCDiKufWSJMjKmzq+zSeGA5qHyyAE3g2CVOH3Is+1pMshMHM
0S5SFhIbIV18yksd7xf7/1vOURq7b8g4gEoj0y8tdcdqle8gmeIrkHVW37NCHxE9
Lm/q31WqmxrVuFMNwapevpcOYheZztbPavj4t+LVmx9KnLi0RR6kx4QjS/+U+BgV
G32p9x33Mv8A3y4os/KCtRJDWwjq92bsA6MmhMrrqYuw4X0oFhVE4d4elxJKqsSH
/5FWEHHOrK4CmTcL2QY5RuiUeWsH9bHo8aDuAEd/VFPuAroru4LLArDidCrViwzq
ojRoEfh8NRecXUC8SyIXryTWKmyik688q1ZIVTfeRTFJb9m4YafPWZY+S3U+KF+C
PBbDgVXeOvJzEfuBPQR4kTOw58WyxxDXm69oXDEhfsVyE2jyDPvYn1S6QdjyjEH/
m5/qxbKLnIrPAdkv1jqMwLaeuS5IsmWJxuLSacU0hYq6X/GnB+cABbe2sQwqkhwu
ve9etaEiCk6WDhBWONLv/E59j3XzEQpxjFqgr4+Eenq2DpSKZpLMGzd4tlDDdOn3
A2R5MTuhoefNcQovxsXph3GwjR+VMN6k1kPBi9t/lepmLsj374Ae43NTryU0YS/e
/mam9y3bsfw6bE9LF9DdwQPZdR7RqPChO0clxAWeboc3O0m2BqwhxfFcy4lcIjH0
tWlpgtHloeY//0+4nSZ6a2GFVYrSMgfOkQoQ9GWD7oimFduIMQt7x9kTmbzgduM1
0PP4uwgKUhWO1ysDlggYEEQVerwfHgklwTSwHVl4JJrWdPeInW+hqmPTkoypDZS7
xjc0j91mu/DTIufi3l580YaQGGf7aWoL+ZQpGXcspVDw1W2UHxUJ1+L4YjL6PprB
Snb90XHjTbfnNLxS2JO/nJN/SwUuigStzFyt+BXE2LMCg8J/NHQ7aMYKMd+Pt4g0
eBOZAycvFJg/dMX+zhTxN15fcdgYZ60yQUgrkOdMe+ut1YRd4fC+RKC3EhkCd+Ia
JiW6UOtaJ0BDXLdj9SDtFnlmcVdH1ssu3IHYxlWePS7bHqPE49c3EgftNgCNdIU0
ruqXDLMivkciP/LtFXZQkce0sUG+vtZkyfSbDwVM2QRd3u5pbIzkBHnWWslnlfgu
mMDokzVdtk2wSFIfxlViNxj/1b7gZGyW7hmMJaetixwDsjcYqRIErvBAS1ocWrHE
ywrHpxXbDfaDFuwlyTwienIN6secllq5xC2Xk1Aq91lf6q6cLkGlI2YaTQcWJdCx
hnV60Z0JxDjo9yaHRz0GhHqfcC1MM9ButABVkOtGCYgDShM2BAx0ql85DeNFjCFP
tzo3ssg0dVLxHEPJ/klAZadxsaefz7vAqw5DcjqO6baHM01m4n27KtG0+5anLYB7
QdTT7rMs/JAvVcgRcI6NYMtE+g26CV4PLM8KDvZQETT57fBnaa2xDoBFSyn0SGUO
duFc02e1PI1T2XVgb1inLq4Xm7z3wRdEAXdRAwdCfAB6FK1AK5zjTsY0qq2vYvS+
W51+uDY1achIeJObTAR0v2WL4FrxbHyApGqKEWkVIwv7bJyokd4JoJ1Ll8wBjorl
73UWMpKpj61hrI+o1cQWHdLslM56hf+D2+gHI5T4DSCk6DDid4qFD4kUSBm4aSTv
S9KIFmicCrg0BC5JeiEaxqjUzkJKW8OWc3BIK+c8JAqVIHaxVaGlmpwl2yd8cZ+z
4ZWWjPpAAjxfWzHTzmNOFVgfrpk4X+NqmxkKSagkHXpMyj7FYGLcKaUkJLc7kAwV
yFR7tl5NBU9QtcXhDS59TuhtvN/7JfxPY6V5zCsRSut1uUUv9CTtFZMtmUZX9Az1
DyvLk+O8ODmVawqbisrU4HvTJkhJ2iRQ5TdnQossfFCSquj/4EHUptUJu/EL12h/
rPBYPhXl/M2rms6CmA4XBVKQdryektGTBxkKa/PEYb3QwiRIVqsus3OaLV3E1w8G
9XOfRHJBodAfeSH22qfuM/ZCPm+qEksHprcfzChLRatSy0nkWYSeMtfWVjcsrmDG
AyTu1wKawRxk9H6YyV3jq6Ty1uAQ1ZB1E9adJn9bGCRX1C0fBtUghkKKYEQM8M9S
TmB8UXc0XYydISOs2VQJq6BEUPya0BbT9tXHpWbBCInz5qDSqKBuyfdxZcYs0BDK
lSRGsVNSs9eMKvrKY1RbUaWmuDR8FX+IZXH+0dsRUYs6O4P9FNFS1gJPfHbdWExs
Xt/pIcYyRFR6Rb/JFrwfkS6BeK+Mlej9A/pZkTnSZCjwOu5IfCwNY+FGUFT4svMM
bmAgguNCyVoHFJURZkdH5QSsU3r81MdRcnPTCdk3fFGLhAfsiDN47ZwwFITZHYwY
ttBTj1udG4+/v0PJ48rP5U1VRSS4/qQEZaFCYvCGpPNJRTyCB2DAG2MOS3xSr/s3
jkHUhDJwMf9UxfV3sCaBaimocUIiDzbCmvtxcdpbqS528sibCFOsUDxnp/C84Zft
00qFVH2yyVVlA2sZfNbhBKt+Ft7dYkMt5FwJTYkhljGc5Ss+VM8YcFMdH7U8V/ix
1vrU03TpYOtst38RTeoyzS56OJJzD10BLCxSErOugmaBnFillG1rdGv5bmRzrXXF
rDazboaczlDVZiGPWsjSK5I8g4Fboy8NBrYX2CiDv7Fg0Nuz6RtQbQmTlSENMsly
T+N1cJnzLC/Ahad6s/Yvo852xagwnkDDyTrzkijIQLUVn6Ph2vX7yxewBKTjO5yD
8TEA8sMxAH6eiZ19fkGVdK2V+/x5j5Ymqnwghers+SceT7VzlpqH8rllSVGWF80Z
ARR9jdPYgP/aR3uRtN5TNxUG0pH7Z3udz1Mo0c6RVO7Pu1/wfDZYuT83GD+BYhhL
NGrtlmsfytg3GA56u9PDo1MeMmw43LbloEZg0rRPQ6OJrbInoMtx7kIVm2hC5Hye
DZN2Ijf6TMhUiEHN5CfRvNTAZdJJWJhr2odFcQ2IYMEkQKUktyKrqE/hjb53pbyA
RQAXzpaNNeVgzgxREBi0OU5a7ETQ+y4vqDt4wQPOa0YH3y/bIckhJynbH+J10/nm
0rXsjfm2E/9aW/0kyJ55C+deHlleAW9e4Tf1qvE7V5UtQ6unEwwJw6G0GkaZZjGo
08wlxhvEo7GWnNHdYiXJ3QVOI0CaclclBzuGMXzhePPwSZvXqN70ww6gKWj2CiLt
k7PKDY0nvzMpYqR2RLnukqrsfY+eGrXoNjcxEBdYXzDJiRgKc1BRusYQR278ZW9z
2H6KCPnS5QDuEOSeYyt8U4NTLanjBSNWf5n7MEOAFbm0dhi8CSoQVD7RrCvd23lC
Q5L5TsXKk1zRBgjYgZxpP6RgmVTRSf4m4RdWmGAY3otAovwm+hW3vqwuF2/MFK+G
mTTk2KQecmHoD5P2ntLfUN2HD9v6WBl0Rz8b4/RAhEFr1qSt/vB+mQHQLEHkbiqb
9p8kobSlJjoXofLIBrFV+nXiooMY0bCWRp3aYW7OoSKCRPDfGNXG3npvPWSzLIIe
5CKZtRIiPdmQlFrjrF91fy6yDZbbS9i1Rf7y7tR9RJQgAnBpMqn12MW02G0g5rey
WZmAOiQ0YGtWkxOi4SOCgC1VR/ShgVre/lkAezDWNQHZofMv/j0dUAWEDhB1tfNf
+xKlUzFiw6lQ5Z7dXAvRK78h+bPhIX3+/P7t+swxzDdiN/XFXoG/aeJvFJnSw3qT
R8c+rCclh36R8Yi8+0z9CO14b8oijr0SPe0e6JgUq5WDTwwYV0O9UELx8vH/pshP
5pteAQh2BKyM6LgYuGIWYA5B0HhMBlWTqUuyizhdO/vxPHSjpcv2lVKeqMsFhv1r
n42K5mVvuzHlyruykH2IO74Aw+erjBuSBQalxlMjq5xn+8vLhzZgHnGgNRr38Q6b
yhEKx95yuLXSFdz9ESXnHn2x6licPc/7Pj6aVzrI3zkGevDh9pw/RQXXmHqtDHKC
i6rSb+/UxnYLPwJtHB2mxtOvZL51pFyHoBDcfFxR3PLTZiqOldzXxOdk7zhGZL3Q
rwBQCNfdQKuYaDU/NOxBbQDNxiJucWP/haIfVYTwSVGaIyF3FD5gb5s9aHhBtkTd
efapoxUiSGxYXL8tzfJatydHsbuLzI8QH4XRY4S4+yHJsLILXoPqj5tZXnhvWEX4
dVm/C7QW0luosLiVSYR1H7Wyqnu+69nTxk578jRd6fN3norDbdI5ifLBSOlP6dj4
qxMtFucQlBVOCNmUoiwyj14N8Rcu4SAry5FbrsGE+EBBvB7R7Y9vbiPZwf6NgYlS
3TudBma8Uvv7fvNjvkYSkdzIiQ0Ou7kAPeroxOlLFwKW7jB+2mQSH+dbGhEfRQ/9
QBgnkGBHU5Vb3OUcR3Pm3AlW1wh1OFY+mWCkP/guOaZnpLJDVcp0aDBKcfFgqKoS
sW9oy43AsVHpQMWxEvIXT4IYlmnuAF01Mc+y1GZunFBcYjQc0ekzpUArSe/rgzvF
3/CRVkzSfAb9M0g5wLxTlokwWqyqR2yBMzaSmG6kqolhUGZ1xmtFeN6cTIkEtg97
JRqYPnOWNJOfqUp7Jv5ly68v+bH1XUHTHEgnwh6Kk+N2Z0muE1Bgtyj2Gk7FZeQA
sA/UF9X+C67fbXE/Mo6hrxqeaat4gE2nKlYECx6NMJ1kZuSzplBsiZyX3yTSdUcR
sIlveTvbyQRDkC9aRaGqmSwjr1Kf0pRPq+EOPkDpxVc7h/QNtZu7ay7TXGFuYP74
jktAW/3ynE04Yzssmmr0YldIHdvRlQASxEOCRyxi/o7+5+YZ3YbFmXFw3UdsspAL
q0/I5BKdZb778BjUqKGslrLg1ZcjRNzj+hiLk8d2tQ8SDZnCIoY5Vf7ka/fFzB1P
JwjNrJeycNlnqX0IEBL2cXNiJI929rwsuBmWsb+QsNyxvOjYZIG6y7hMGGZ07PQ1
2ayHj+0eb40K8zsbmB8COur241oKNWxtXsSldCEcz8vJtkC5Znhz455d7J0Qpp7w
ct77Ss4JvhhyRIHMqpSNq8ymPfFIWIbA6KdzdazT5UWTEUnYVO/3SEv9AZdQuV/S
gp3Y7lfylGsnY96YCemLuYwSg5MzNaYUkJm6OULtK3HQVXCh6lT8yxtxgYS9qczU
36NaaqSzCBfpdwbhFg4VAuA7uC9+Y4dQi34FB5ZTkSNi747NsnI+uiEg2wj/Tjcf
tOxpXO6sGPWrlEk3sbERILxvRmGWJhZPjYnxE8Tg3ZjqP+2LPuz8a+qv+YAtzvSI
tvqQEAeGgH3qnyQFUpcbvCq2sD+ns0k5IIkjkBML2uhMcU2wai7EjV2NmZ1x64tf
LdRjDJj9hYgdEH8+KkrMGNG/jIFMzf0gg6fqMQAqUP2dMLNa1OFCmQEPH7g/LuIr
EDJb1prpkDl3zG4HG+yEh9NGit65N3lK/SlqSHNeVVSGJNuZE9LsZd8UeUrpIYc8
4x5Z/ruQocIkGiXVG2N0gH/DSoJ2yUiPFnFsDy2ocgIuy0Pk/LOnGywczLj9Km/7
ieNFD3VKMs4/1TAJ1SB18psuGjLHrxLQ9sDYYoPrfjaser3tcdds8IczhIzK+6SY
00fEKEqDLzAxzo+Qiayu/PlQlgZfaaJ8CvAvKZcmL01jgkIkjWr8Q2dwKqCSi1Q9
KliFwVN4IlGWc5lF7Zm4or41dRhUHEGxmbXNeJWGwahrRvCBOIeyLTRquweMCJVL
C5bo5GNM91bPysmb5O1guoZ+TyPC8JDhTtsTZHDhulWXg8/GkJ5ipiwnDoQmfNi2
lcCMpulkCh0pJVdIg0II11TOdYNqr5npBrr8Rl20glk8es8+N4Is88dWjCjKOZv3
GIxMWikcHxJ4Vt1TN6GwT61U6ZnxkMAq0GnSw1idXgTEoqe44jpwReI2rJbpr02o
ZdRq5quqTX7ykych9i8go+7C9npnL7lhuxcUrQhCcvfx4OxXWT+oUqOB3hPIyonw
HuX7eyH5EtlyIBKnRxrb3Xyz75TuxB01eP6PcUkFZ873y4QxmgEoy1vCRw1jzpPl
GMDdFCQH0COLREI5DdCfhRwrGPNnpnII8qB2hPSYPl5H4xSOA9AWcL5j97M2V8Uf
+QA0ueukLdeD8ncb1tIJY7Aalpn8F9HuDjiqaMiOdtd8ORRVCQn92rm9lcVfL30h
45H15ppEtJvAvn7R0h+fkIjh1o0n/lVeb2OXj3KlzFlkoU0fmNDSFhZyDl0RopUP
fuO7NKoxbz9MqMYz6Rmw69QTFicOP4M+LDMcJ9x/IwQE2AH5xZWGy7bebpjf9p/V
nPVdghr76z9bIAX/CDE3PUyrSvJkqKMRc0b5bG6yGDuTKuFhkh7eFsnA5Ug8mXcm
S2auFlkQ5ofemyKZC5HsHl4Os1/RzPGVNoIeX9sPJgEnKkhQs+Q9GcpysgaxOGgP
yvDZiDTjF0PxewNiD0buUMsCm2RFWesNdHFK7e54kGsZEV/57y4xiTetyqwbWxtB
4ad/09M1/ep2v4WAR1pBwgopOK6qUzO2ri/8pgxZwSHULpWaL78Dn4uNyUNZuRPM
zz4YtCymvs4ucJKC/AK1K2USSuvDBP5qo+uGeJ6lB5/KDvxYsxB+W9mLcBMf//24
8fomoV9LP5bhbuTRt9p/cY2TJSyxgEpwPbwIt8QxMko3AGnQ3dpwLjbt2K2r/N4w
zE1pdCaqQPyxKTlPbHtjRC5jq2OmubIzTNLnzJZTCYCMByrslGptMVrK9aLD3Pk9
5CEYJ7Z8FgCgBLCRjFqEDeX3zNzMt1YNaAqnWJC7KVJ/xymiH49DcL0sZBFeke/I
4oFI1TwWuocPMWp/J7ZS9EU6Kzv4gpl43raU+NodfPyMQCB1T+X06cDWRiXuK3Dw
5EsltHQodqFbBy1sprz16xO4C0jfOHF1TF8qM/90vnJyhf+PKYYd3v5OUcEDCqtC
2UZMUiUmQt2lxzaxWjiJswdq3z+5ljf8qSymcBHBpv66PYZNWMw6c0tw1TF8tvzt
gNZuI3F6bJ4S4MgkaGyXpPNyaSHmbyTaaJcEAz8XlfUyfHv79Usugj5VZ04vJ7Iu
BHTL8brOFIL37NlddKwPaKeAxqqzRYgyJrqKui4FOQrXjXjc+F0F+nOLdH1oiHMp
/SOC9RqFE44JZo6DvhlJV4gj5ZQO0L6Owlp4G4yD3m4BgU+LHXzQhxUc7abQO2op
hp5gLfsbPLL6yN8PyKmdpFV2CZB9NfYU6beLX+QcOL9gdtAMvCSKtjqYsgWyFvPv
W69cJ/Z1u8eJyKk95w9sRc4pGrgzwL0zvQmTe9+xfD3WBw2QR2LM6dz8DleZnO+V
Rx51Y+mmbISWM1Y75CPpZeHGtFF4lMCgIqGJfAaJo40JreEYc5Bj2TjuSgqHcUUK
wlU0RIzZR7RdDMwAsnrCtkY/2zTrlmcehK1899i48mHEYZdsG5daXLzAgYpDHxIT
bSTKqfloI0svEvscSwFrrs+a8cLeHMZIzv1wZHonaplXHUrdWOdx5b2D3s5j1fZ7
VQWed9fqGw+3l/6O3hc7cRb0PT0FQTPZ9PQzmnurN3ls6TgEIVyaCzWvz3geRnLg
whe1o+iQy/cL/B07nta9sQGwOBlkXlwrpQWylnuLwwZzhwVfIbp8JOXcXY5N1SxR
NR+rshWfPxgv48wHpNR7zjDXLKjHV9B5J/ddXJULgrq5zd6MxUBnnt7GEEu7NpZI
1qLddK35naQHD0B+DzkL6DJhXOZmoOPGgcRSEUQxJdjHnxFYEu0Xhv9xaZ22Wzud
6cO4g8KPBayo9QmtyNcg8m5+OXMIvH9xnXcUqHpd3FAyfREBpCMay1LQdAQH0du6
rOG5kk+4SK8Ey1AJvzXRu0wjj91HebYgwTYmpQrAI5HaBkm+qTR5bZ0o3iq/lw5t
1z87QCOTMitRsQR4ZjGoUAnozZJWLoilIZMSa5jXiNfH2KjG0ItaHzPt2berVKRo
I29yWbkhflmgQhxnv27oZoJc6QD/r+snpuVPFBosRgttkSrAdfM5SVPCip+tM04G
Y0hkJDBZI0kUr6c6i+N6HfU/A7O86juRYXqK1SdMQifej1sZde1rddYGwteopgHV
SCAh+EKXy6TkGtLj5Ru9r3Of+KG3mCpEGUYea0Cg48EUPhhKLsdWU/+h7C05N14f
QpN5kyvBesLiobUlY23iJST1IlnVGi5i8X5rnE9c8FFo52NDKi2ooJnWpAc/VVqo
mulqOnj7KokO6nH8D3WNZ3tpWt6u2pG/5XEKXHV9hmy8A9n7mBmlBILlb1iqQ19K
rMH/p0aydTM1WnL0fpnsbGn774zqF5cMXI/ILq/kUr8hxg+Kbh4nXkfILAW9V8/C
dAWz3ikLLx4pvvO6RxhxLzRaud2klOBNnaCkiSbBScmsOL7E8TBxoQU5voGfJsl5
zlQmbOvLpqy3zZUkT4vOJNg/l3AOF/uTIw5By7bUAaY43xwW6bmx1ztLcHdp7ZyN
7YZsrv/9mAXuAx9eXElQ/8cwWjsmt4NrL7UIzPxEXqLSOtpFGGZfdGslnA9xMOpT
G8gXlM1Chtg1QAkpzSrjgzVq9XxDG3AfUSNdlEzwgOBWJrIKIKBWhs4DsCFTOfMq
eC9oKd1Crz2a4NaOtakOcWG51bKWhdT+KoLlHEBOLMERt9IH0SbDpejQ2yd9JMqy
vOmLz2UDmIcLFrQVG6i5IRWhmHgoJMTnO881GTkFF85PKWsXl6MC6nsGAL5fjqbt
+6d/R8vLe9jX8kHHmRiXNa/NIaIRf6frkVln0rjGe8kP4KFm+Wxx+O8XHPKuUHrI
EekswEVKtnQgj8sQr4WEo7ZNqD0ScglF+7nV+Kwtzh8fyPl2I/mIkmVxhU1gBIUm
VcMg2huZKRKQxk1hJG/Nnbk0qPfbh0pLXMX7XW7TSkT5ZXyryzoSlgysHAeP5yO0
mii6IhCZzx/Tm3YciClKwlRXEWBkW/7AQVpscvBLs0WHlW6PicfF9E7x0W29Hb6d
Evlz1TaMQzne4GvXAB2pyQkZdC1splNX4ZLCDrL04OQ4Kbv2fKpqcOk2not0rOtn
QVVtmMJx9X+SRQQUeBE590yHLPW7F2HES+aElJ/FADjG/2hUmPjI+07JRtVSZ1Dr
Sl4Fhqa4HrXv5chQzclCAd/AgCtG8VxbIS/Bwjrc2o6xGZYnUxYhPPvRe4UxQhjJ
ypHGr7letNmK5mq6v9HyyVdqSC5C8jpjo29uYn2VOvlBVD7ye2zg4w1z2PIYNc9L
ySJzhEiDl6i81tjoR5dIvZ/tHMEkYwYGtuS/cRGBOyJgf5C2u3sqIDGeZ1wrJ5Fy
+69il7HC2Bg9YiraTBR9Bkjtz1lUpv0Vop/pvyJ69trg4NfCQek0Hv4plmsz6HuI
oawtGo2jyZysL2hAFn3FNAF6tOaRrbhT8rY8NzeIa81+VCJonmdZZ6JMqzTiYnVe
cMcRuACpCGLlDa4oyWiZUik9T01vejOcMXI+9AXL2MiVmJGtQJqxdruvuS4r2Yhb
zcGbJAY3AhC5K1c0eKBYobJ08Le12aHKvfcIpjR4NeKbuzNqBZeZORJU05FE1B9Z
cNEmbBru/XPtb9SvngpDV/r0eJXUZEyhcdseKF1q5HauA61MdM+WvG6sCjT9f1L2
ZKJ+xH3dzYJSUCUvFg6XOAziSNqg0FO8Y+AQkhaKOpsooOyTcONbdkchZ0z0JwOd
0Trm+JQDe6tH/5Z6cKZOoVlUoJBVtWZb4W3pqDvbDWMZHBjhR5g3wT+gUFEuKK9N
WkOEOtf9S4r7w7X2aNNdpFMO4Y8EJwBv8dBL+ivhI300V08sB6xM+YLzB4RzmbMl
ODr1VISxW0r5l90G6K8lo7sa+/imgGnK/ycrOUD9OIDwlqxBEBsAeqEty0TzlYGq
iQqMFQdSGr5SaPwaSzmx48lDXlWeXlQkzfmrqJ69jPKhbhg9ZyDe2pLo1lWItSpe
Df99Nlytzu1FnEQC0iRCMATWd0mN4GPi8A+GMrJe4qL4RKYm5Egx+uJ+e35CZVRY
bsTDNvXUTQhcqgGwoss71z46rsbftHW/xnZpZfzAwjoOWrZewOwuS2A0+uLBW81i
TaH+2oQsUljbA4DxFfO3EEX/P9pCuLAr/Lci295aDhhJ62olId1HkAdFdBQR+OYL
KkA4Mj05e5YHkDucisZKCgRZ32Xg/lncgL5YkSbOLW0oSLMBqMF20G78/y7Mprvw
IA/4VGAyqCKE3nrWYXFVqL9SL6mZwv4wQ5LyGUU7UT25FnfsR1AnNAcLSVyAKdEI
CvpFcYskyv5eXsioJR5EcbjLYZLSlZohnzrEH30jNp/saG4uaIGmVIh9mOmAFa9l
7MIeUuWDM+dhCqewWffh1f+EuqBPnSoPPAfZmlffkKudqSqCXDq0ovsEm/NPp55n
ZuKcU1ITPA9MwoEHEcAAJayLRKVNZ3e/I3D6fCYpAdxN/hPCI9EiX6GCJ5nJxA8B
dv0LMDperdA6E/zPi6oQ95xh76jF5OiHeZwKVI0LfxYIBAYoJhpoLtwtGoYw7f7k
ZhvgOvU6ZA0ZFQJ/bKHKz1PHeMKzQbOsKujQ046t3FlB64dn5WXS/akvuuJlPf2O
x7xXIHUmCragIcBXD9e9mkNwDIHqdubhs/34sHS5IwMCNRPNckP8f9AXHi6VqbL+
cifgsjhDKgDa+OdMi/ov+oJsiwODqEZS4EGVHXI9uT5ICC/+JKVbnJqqYteBaOP5
I22dxkiTo66nm4jOY52FflSt+KAyit+gqmxLtkh0+cZdheHAbrp9j8v9EPeZthOr
aAKAL54SEkPFTeqRBqea3FALJrX73oJvIa7TFPJe0GdboFff299KoV7uOUGSS06x
fkmNKFOMI/3oUd4HWY+ZRpIw2Wjg/qAaY3gBVDrvHl52d//64/+RgNmqez7Uh3Xj
E8rk518ePncKXgV7weQTbu0vtKSISwlJRw+mewG7L0UZPKms97X2xJ7mEwdxszDN
U4UvbPPUvDCzqAzdfi1kIOVd8ayBVWJvVEmZPMJj8riD0Yb9dbPL/0D447aYIPBE
zjJ2GT9M6Jv7d23UXkUJ5xgXRvukTo0Tn/M9B46CMsq8Zrfy3TQRQZq3idkhvFaJ
YqNqH8Sbx1hSieEsdp9Dy/nuSSX8x/LYB5S9qZx1kdl/+ptvt6uMwv2mhSaj83vZ
MxY+3ge332dZM4WbmuE+DwrwT762Lh0GF6p+rkfXpK6YRJ+gt4rB7IPbhtf52+Zt
K1n61m1AYNYrfblEWnali/HkeIXJ8XLxGwFVlCVMLJU1vDj4wzKRA6pAIdMDa2Mq
qLcCrxs8ixyZQYt+l8VqKUmd+Z01gUsFNBQ56DVesVJ6enJgjF4lukji85ca4v9a
I5Q30MbmWEdju4Xyz9VlqB/VDhaU9VPshIQ4ut1VMIQV21C3ihMkBCIYrGu+ZgOA
ZsDd721S5jBlmMH2rWTOJCC8W67SC7OkyRokmB2IgY5w5+xD6sIBWlzY8gOFpqLr
gZYoqixc+5uFZdy3O5KCN6uube9P8i1EAHz/g7zL5dchmFLOBIs/myZ1k70H56wE
oohzCtEb1cflZ2aVShR0Lhm0h0jnTUX2Lf3qH2mRbGrGRlGOjRUy0yExJcWV/uYZ
v2w0aWqESqP24yItv98JYRjiyGj+LFLIzOzKReI014+Sdjig5uoP4q5MRaTVxvDC
BWn4BM0p+S0WhMTNxoumdF6EJzWNla+pGDJTgOvt+1PHSz8fbUBGM0uyT7QM84EP
V1KtU2Ltlf2F54a37m03DZcKEPc26TaChuSJql8QFUk+p/NlSahpe7TcCQwOwE+Z
CfONvnsERUR/1KIuuidS1DSjz8FtUsKg5LyugoPxPhdxgxH8Vzuts/bEDt30GofV
JJFNDu5+ZSffHFfN2MZYDqyrtqyxnZYwn8XdG3KJotShbBbshGP2w2ovoHluT6lV
uMCsxj6A/rjzUnGd+TV3ezMIthwPRnbcTXhK8DLGFueAGwfwaG7kUOIxboGx9/zT
bSjScZZMVVq4tvn/fRqO/2ieAu7PqOz3LDGii9vEgFK2UX7SAz6Y0cAYGsk8UOE5
yIE327e018TxsBWTAGl1HiMVNTFS2j3HppThQtsuEnCDQfFphrufsEIMHExSrlMV
+aH1pcmWRSy+NB28boIfJah3ufv+rF4XVCeIJQz4AXhsNoFjGuTlkUbJaMgHa4VU
ZnIPg5Ko6tiNS74/AXB4wXzhm1ExJnwC7S6NIOPiNr32TrO6qjw27EDzeSwTT+VZ
6vUer3oDWqnel20x2XqLhj8x0TPhXPZSqmPerYFUU7cLDcH0/WHYPxYTH1jRLE5r
YRbxhnvkAH21NrI/n8hgJ69CMJrPbuL7KMtX4fvzPIM2atuY6FK92XV82CtoPOqq
EJxzmJI4RKnucWjy78HTZ4JVhTSbpBr5gb4mAyevIUqqikaNlv8xQjwXvEm5wryf
wF0EWHegwE/waLrdMA9NMjjiry+Idx+SbkdxQOsvEMRKyo9yTnVpQ1UX2Tut3INm
2L+2xKd3moZaxPRc2UE0j2XC+cdnAcv8Qo6X6jgx30UScw8ls859y2r+0zTqmh8m
0RyBOaviH6wwjhcs/eI10zVjTykvSVLahNZ8Fs9VXbccoQenKn88Q84iHM5gFfQ3
AKeXiZEOdl6lCirNkCz7VHOIF6TGmAW1oLLWkLJQWJdWUyY/W6xBmPmU+9CWaujG
a8BZu74yIm7gxrgY8A7zTGiJEq2eMVDG86rRh3T2+5PJARM9Y2mcwy5KsIrm4gMm
oysdxvDy8puqiDuN8crpenTLdEUQ/m63S2gy8dy8dekc3tWjRxLv3JdNkbm5rjI3
OnaXJQBxJL10kq6kCm4x+cq2h2xtJFsFeHnGEuQaM/LYsTyvpeRhVVale1ZJrWJh
NqD1jtvHE9vhFs2YKF/yjJMmiY9k2N7vX/6Ms8PKvWZ9DAadJoAvuOjkvciA4SQZ
E7ZjEvwj9t3QR2uKZSWThN8ij5PD3FulPXNVb5xVAuurDXaOw5Zt/d4P0BN8AP5M
lYYi49wxizn+fQcS85cb0/vXxoll0kz7X4fi2KBfqcDuOTJbEOIKoyBP/NNi/8fP
J6GgWpfguNtipXICFx+rEsXHnLRqnKdgB23ZYJxAVnEKdiYXEyV+Gsb0XuQBL3Xk
S1QSM2zR66OpkwEu2XqyhWIU1A2sWBCaOlpO1e1BIYV4TYcIJ/fCel4UqUTqvi7I
jc9Be3ZTLmP8phuIla4IrKMWNnnKb3PDM0V1A5dk0fmXNTpsE3v5JAzPZPhPaWoy
oj0kIZ1iqls2xVPQhrCTrLV4lWVscd6jGjP7oqSgh5tvXK8QH/Sx5HAEp3H/BPb5
yaeQClVLu2gpQ5vKFhbHkAwm5VDGsWZu2LvSTAu0egQ/kbymx1O6Lzs6bRE7Y9Jh
a6ed8nurvl10Ki363KX6fEmCpJJOmUnncc4B2uQ6AfYbwouqQqVklzebfb/rYNF0
wotjru0gkC/9Hc1sjjMth7XAaAQsUdDeZc9yc1v0S+9REFud241fNUX/dn0goS74
OBjx/nfi8P4NGu4zV8SS8mVIhKeRxNH1MurZ8opRMJdwacAq7QjNamUmEiDMTT8K
TT0L00qssD9nAgZhQmrX+B0XlFRrco8smMHlvvwxjMZT1msv1wmXYi3G4iTZw1eD
kkaehwROFEY0qTwRO5XrcHGM/RD90IOpt9Q6JZKmt5OoxM+TR+QiTfaeL/8qdWeO
sdrRXcuV2UxwQ2aLDCqx+hf34nWFydmCGTgj8b8Q1zeosbbsPvxUo/KBikKOT0HQ
0pgPPY5vHAjwmGLzt20YwJStbHyuFB8zhqnX5e2JD4pLrFz36MoDDXeeuhjkxCE+
7LxW4Q8qo4RpanZiR1+uAEeshKEVncln8OeDoFmSqsWzINm/11Nha+USCCQF5CEV
TSlp6cLi9hjXSELpaVXw6UA0vnlaj6Mp6guiE/G/qGbv1axHgNk1D8HdYI6Gb1uZ
Tkd2k+V/fBAeXQvarqm5wqwebxiSJobZx18IPGYiiv6BZvTAQYXTlwUIY6F63ZxP
u7Y8H6wBthSL5lmpQwdhot9TnCgBSS0WMz3+1gkX+TjvzKAMcEFZVFYVwodyAiu2
4SoyS7NUvmJ0Xwb5uaDcqjLg5jA1ksQCPObK32JnDawN8/1PnZs5M90DzumpRBpl
1bWYcpR10oppbhXfUzQc6i9uCDUBgcNIKRpnes16a8NEEcp+YCYVZtXEeQC4HwEC
bN799OplQLtzBpVFbKwgUqjRO1MnuOm7EhAvVAEZktcOHMkoYdHrtKENuMnuuiJ0
oU2AslXLAyjkvFQQWECENUjky9fjvbpFl//j1IuBQt7/FC3X0UWuhaALSaLD8XUC
O6Nod/4y/WOeL2sRtiyvmyPC37weigp2/RuR3l7shMQ+WT7sCtqGu/OzfCtqJgKh
kbM8OjneUldESCRu/OwRliH9zC0HET2WjHsWWmX5TTMMNjA7a4ExxvfbE3p/+vnH
XMsc6xjSXmwoP6mdDBBHHsEPjPkAPVQJFLabRiwsmW6qFiuaLehWCQVAK2sqSwZH
UkNPP924JH0DhjhNZo6E/70+64paJ6ZxCCHNFWRBm6+s0KglLaYA9DdPgnFRHP8A
VNyd4noJzDmdmp9g+0rxdCz6MIpjOwNhIZb5fHBdTheyg0UWc4piGF6sCWp5h/C7
mZn5/fapHf3NZu7b5Inyj7iUzFogAin0pGvAvgVP3QGADiNxbZRG23qW7LMdpDOG
iJFDUh1feFxmIxaR2uCuJVsKJH82w93Dx9skWv9VS6PZ1T/0eUx29l0nOvYlvo0E
b4shxAI+z8WFp7TKnhARDbjoNAo+UAZWzGaOGClqMh8uR1ki7rdzrS4rqc0MUjOm
zcnBxuX/xeuIGVp5u9LjC5HMIqYZpuxzcxCeOtelcejXW8+COPCt2kSnKuU87nG8
wDeaRbWCcx8AiPLu4eLktmKKKkQro51n1V08u4+XOI6HSkL1R491fJz0hWgMFvNm
TM6oykbGkaM6SuWhO9N11tg4MxX9tP6lfk5sQYvRmoUlceUPNQj/SATOl4pP8gDG
5ITs4oYnX+9G5yjAO+vN4X02Go8pcZo2qY9RCtwqhFRabrPRbqFz/i/Hm3LCNp/y
j0xNnEw+xOcVO9WZZohlPBZc9nxEFs2p1Sg/Sv7t/hYC8uCk7MZbpVv7nH3bR/Yy
YIcdKN8PPlcRhBweMG7AbWydSyzVHfFW2d7Ni5cWMsVYDechxx9v+rhPuIEtXjON
84bsaq9rUMV3G6q9CJzH1mAmjFW7LWgnmE5SLNDkok33u2Ufdeih4fAmgkztns2T
uPIyFFfZnVi5pHiPyat+heGXpXnFKLf9e2vGeT7puoCEPwPogVkAzU8Gz4viMGfi
cxaZxkgWNGfmGGKceTGHutsNxPchxGBh5knp+dcFy/+w/NtSJ+h4wj8UTLQAQNK+
38PTwggDUezgR/nvyoMxk6HGUOzsVDDWF8C4T+lMgC0afXK6C1XgMNZMyyOP+gnI
2XzTnBX5yzc4N56gjN6nYLk6BJQWo88SZtnTNscfGYDQHEh4GBpdWOxOhO1Xzz/Y
5iSjqvLlGxUdWPmYJqPw0M8x5ciFXZb9pPR7BnsDdp7ScnEA+0H3Aj17S/mVjawZ
cMQ3qPZnIWl6FT3Xu21bLPEX1DdB9T1sAhqyv0UhCzmwcvGY99rZD8eBqUdaHFUe
rTztFb8Y1/Bj23P8IsQ7xBsgK6qtyYsspUKKlPrf3k2Kdw4j2H7VJOIb2gG5NNe/
X/ZHLz/O95GLB6xqy7vdF3dFQr9daNsvcx2PcALx6MOTSQLCNJsm+ghhXuYg5KgY
JLBZ1NZ0/y67r0XNPjz98sDNZwqJ9DwxxkJMMhA6+rH7pQCUn2IU3h5bxLq2RHag
p38Zt6Zk33qf/w1ho1BH1lKrz7OpkgQ3XKbgUm3twtE7IjQ0U43w9zl2p1o64Uxj
L7mBS0ro45xzwoa3LePovlrLmGqmdZ/eoL31S+M+28U+TyTbj3aUfAdlIIirEDyZ
ngatNKcFAgR+TkDogkIzdVMQuXr39SH3BKMt4TfXA8eEIj14HYT9iv7NlpiDlYNZ
20zu/RfzDw5O2cj+t0htEivVjyZr3pLkZrza9y6LO75j1cVUTwZUwC1evPK+MUQZ
WTGfwLG/1Mn9yFkB0EGh9sXwzT6e6GPsdEWjjbwCti7bi1NTYEhnicfumBrEapRq
/dWQe1OP7PoVcdTUr9yu1ZRQ9i4ktnjT5i5gM2I8vGlFf+5fG3lw7zyG9t5jUEwF
FpzhHprqLp7sYCDUgCsBabzB2IUfPXZn7z5w169ZFq5suGPzimJgXihswsYGjdiw
aIWZ7DSu/doJLbUKMZDSYMWFl8vSeUCh1UrC+kPdnXcFofTwaejLvP2rMof3JEsT
ZSCJRqICfKuTq9pMhtjyZ6sycJxFS6hpw+SiVN6zlrSMntLTYZp5tRYs9hYG3oks
q3uloSZIGVg1IZ/0AGAB2ZeAYNKQ0UyxEf0OL4jCIT2oc+mJntDMcj9T4JmzVw0P
WzWTAy1uJk63faoczf5msyMmLHqYd/rUrPWVYuTNLZY9iuhM4gk3Ki0uQ4RI8b27
LysZf/ZzO40obFizO1ShodV+CGqxEGiBJr8Qwpz7uIPW3La62Bn3Q9MTDoO5epW9
PEXdP0p9OrR3X0CxUJ1ujwUBBZ4G+PsGpksrh2Zdb4zOyN15sl/yz7Sb4pJy3B3c
JPa6V1Rj8y1SyCbpun1KTXMSwXCOjPqXjrP6s64f/7QzR5JQlWR0dUXwUwWq96e+
hE7Hirajh1xjQjr1JzW5r1U5Ps6icfwYkswywEV4S/lYhkxs4WxQtXNOVbrsGtI5
+CH73ntHu0OvABsH7c1nA7dZoAB72CVpsiWvd3mYIzLh/x9icnMW1G0SNRTZYdwD
GM/F7zOHXzegx5rCQ4+Z1rdXLpG2ZP2xyX6WtghvAezzckg+otjhUO+3bR72exQT
TpsS4fZ1rq9zSk0FaXHbiQMZ56ICwBINWMiMU3UDczy/2wW459DWlvHweLEib5QS
4ZXN5FxqIqUOJ07ohr/17AM2Dbjko7SGHPLBRJGoaq8tg87Bmu+cv0Y30WUzi+bm
JO/RlYxgc9z5GQ4wGJLM/gjI39dVm4c6LlfLgU25rutXpKUjMIDc/WusS9y00hYm
prw4URJm57HQxgps86D/O3MCKOj8bPNcf2ZZQcxX6pNz1hjgmqtsxiJhL2M3H+Ge
CHlijX+JwY0iQ4n6WOgq/HzZRK9JsE5b9Yvw75lkYg+wja35S/4ONabCpoFQtIC8
9l/mfKw90TrggR3I4R1CZ78y9rgyNjXWIDXCIEuxL2ZHJ3OBtjVIElZWayG5rt0t
fdbZBE1iV0E9USOhM7HdnqUhtTjkI3g3qe/ezcLU4tAPd7XQSO3U+W1mOzSqRSJe
tLhc42ZJlv0vT+aDwPiAVykMeSmdS+gW3py8zXdZRy9D+mb38jh/FLuyfrawFQy1
xG/j+tkxoxKRX2fe0Et+NzNs4K+fxsIu2pZqIHxJSQuw8ThADu5WnfjEp962WZDF
nX7etXULq1GrXVGCNKCn8FewsmayK5x0REAH+qH73p2HEsqMC7hXlYKUqdI6Wzzm
a4bwNmN5adNVU8xHjubtV5Bo9qZMCtvFAXz3dEfFl1Vu90pbek6xymgklSTNFr5E
AAHTkGlJSjjh3dL8cQ5cnX7uPuZQFqPqvPpTIFYmRFvUzhoJoej1ndIWlIkcN1Se
26Z8CrZe++9MLLBrUgwas7WVMr95sgIWw4pNDDkG2TDCh0iAbx5znTlsqcU3kbu3
/1xyArjY68g2grxXYKNHNXl80xOIr1fnmh8Nr9WI+lK8r52TDX+lI1xlJgWMlBeb
2CXzjvFyqsmwJDJJJBjz1yjffgPxKcuUTTn+qPqvDLzupec5zuxL6oJTeiWDSY+1
pm2W59k1PAi/54vfjZ4+7VSFRAE2a3qLHDyKAIk5QPYu+uj1OwVjMjflCx53eS5a
ozBtsnEM5M45ek9HFGfFnFEBkIJfzi93K0IFk8wj3nuYGWRO0Ids/wHTlb2W4iZC
ZtQKOQysoX3DS872QK/eiNhXNJ/oE+Bp5Fq+qCfF6Vb7/r7Mjol/cskG64Fciu+l
1pJ6Ki781jGLUJ++REUWmTIfoBuX75cDWM7gWYwzB7SL0IJxUg+i7EDXUH447AHK
dXU8ShqMLAI1570VS7VpoAJvynJ8EVuKbckXSrPApRaGhAwEqqwcmvu1WigWVDsD
vDHVkPWl6VnBXDlWyMFEIWJEdUUpN2rOF5wZwsl63UGmZP8caQO0/hau4500GchD
Pi/RV8GW1vZ7nTWotkrzbJ8JCMcBomxdKj7GQxO8raEIXFNc/SkbmHuNbZCTya9j
GJSgp6Hz8rkH+2D01M/g/nJIUeYvdCn0V9L6ftKCVhhUhssVeu49pmeKxpm4kR+0
MD2lgJMmSTFsHzmL+FvIpkFHdTCp1Fyvz4t9fUw1i0vjXzinc2Kn7t0rsYNKkErA
bUQx2MMZYZW+DLIiftFWiMdcvEszRlvbXl302rBAdgkss9mIV0QaWzEIpHD/tgSU
lkwag36Xhk8SCIyWrtrCqW+SMfyWX6LwblwrxYhtcfpXM6YAtzbsvOBjrGt65H1H
7//n7oSfoePj57sbKxrdbn5KFeXCCEyF+197OP/Uq3eXZiBPNtppfIk0IBs9RxO/
HAbiqh2S0sFbJ4OL5B51HMD04HmZp0uyEz87++jMPccDd3+KgqHn1jeDglMvvVJ3
vaZqUxR5tfxVQFIYMDRC5b1Am/1cAK4aAstK8NDt6k1oRCtB19seQW+dhpnvCLnR
T/nmnrs9Z1dPHnU4BHd60pdDWj4BsYBqf3Tu0HGJcULzirC70/j/9w6nQB/bfOqf
FxDbGoc/Z3YDh8hKQ2BsQ2xRAGhCXYZ/lVLa02SEoHhjNcYLr/ZB23MvzYx7HHaf
vaiWmfpmpqnLHKm0UwAQkMD/gmEgKfkB2exi/TGhYKV/g8NPRzg30QyZJRoEE3oZ
5SWRKxQcnnUd8+Uvgp7TJJ3LrLhpNG/9bapu/6IE9/q0z+cT8VsQslOzhSVNPSxD
8lkMelU4PoUGxg+q/XbElWdW8Ui9NvY5Z0uP42QsnH7BhuxsWH+qVHmuxQcwCuEy
fnQyty0wiGfWlix++2dvsWNiB5Tuiv2YU1sl/CMmfQP90DwwvMy+2jKM3HmSiIUB
7EFajJAwDq9Sw2usRajJZYVN9tZNOQ8BJ+qvy+02IIEsncJ8Xuagr2Ei4y8/pi76
uOyzCBgDy15eE9sehYhB+RzrN/MDerUa7vrH3Bjy8lAy0d5WdE+Lx7jGOlfJMxRE
FeKlV8QNK3dUPnC7PVGSUYm0P5QUQbvTSAk33CHmCMCa0H+Y/erbYjsbbRsFGReW
ID98L/4R9lm8CVR/TH0jFMRaupb8rk3JKZ+XRn2FoSBIcRB3Tb2q0ylaxmstQnbW
Htop3RwFoip6+H6AGW11eB0IpZBTRso3dxirMD89Np10IZq6i2upDKRBdB8pJB/J
iBYXSzQ9xBKjr0c/3GF2O3Eyx8da3vrNV39ia2FN2spyHSe1bu3DRvM9zy0dbjvw
2GVFEgECZzeXV+GIclXiwJSVESIxMapQjNEdczPbAgwZ4Axxo89V51LETc97YN6I
fDHUryWitfkrZEb4XZRu7696zcs6mBwmG47LxHqV/+Seg/cN5KlYg0VfJhl/fN2i
WIF2+CmI+vG8CZOsXMWfKn7f0UBsdW8DMf2KsVBglF1QrdnJvIbx+KBwEIiVNuc6
BojIIzNtYc5fmLNJIl2Q+sTQ3JBBW+XV4HbOkI3DHLr2fKa8ALWugPyD2/BOLKp2
yyVXmls3upBHKO697cPOih/0Qakoa8KbkzsDtKWiTkjdtuk+eLdqwpdaqgqLcpwS
OP3Xc76Pu1fQ2kzcLyRvaXLBHPwJ/0eazpRak/hdbQZxcUIhUL2vcQ8OWW16nsX6
8MZsUMWgH2Pbjltqk6ikh49MU1qGufaGXrhrEw3Rz3M2OYvgeY6E/yXCHhUw0Oc6
FhCGbRTxpMOkeZfX34ilF4Ai49k+knHCtcC+LAMspJqkhRCDNuhKtqmZ8h74z1Ij
LPA+klzi+CI3SXox8YkopDqR54EOQKCHKE73NtKQd7kTL46dYZ5VK9EMA14kJoZj
p7/9/fLja+An42aO4ympNcxpvpE77/7sAW/DwvNuH5rxetH1LcmBVSziQ73mNQS0
Q4d8klQWCALoN63HMevpqtv5Ge9m3S9MxqkGJ5KkQPFWMQrQILjceKJEnj4iPRL7
9WdFECTMIjad1uZiHxu7XdXTn9pB6MTN17FP0SWDljh6P2MTMCkj92cQpEmA8hzl
PZAJEEVc7TOioW0+MDg7K89AAdIdvT/9HIJLpaWiDuZZe4drSbpF9eW07zynywCB
6PPhgA7rUNVtYXnvf40DywZP1VtsPdK+cFtfRhsDAKJV09kCLPfKkfZGRT37AfhX
d3iWVHMr417YlbZ1wY63cPm1UP6UJShmrEd95C6y3Fy2tALRHhORW3yRCNncBgbl
VV2zFJNOREdzVyGnrtJ5aEK6KBDmSw0/Wcbz985T9iuTv2GjfpGG5A9wKlB6l7P0
0k5xGu+7u4QepuQ7KHZWDk5QdORYemlh3CRRXkrCTmi8h9YTttHC+RYNOm7Dle7G
ha18OBsfCiI5rBVtDkaZxReYqbkSHteLj1JdGJa4euO2+a9SpByj7Qtw4jz2+50i
qHEv9uSzuRCEXGbIeNGW8ogq9ql0nSY9WmTJIgo+NTqK0/ZNuJSbqq9VHmBaBjDO
4WWZzjgdvhqjZ0+C+Sfslu2z1Hfmt52lLHEFyuA7IrDnle5f169YnLvuvMcc4u94
xfTzbHX7VqzzGgJ0ON32xkH/ms2nCYOWxlFkeYSmPiKTkZAeEr+mFLWXIoJmMhSy
SzQOkP23/PysnCo/tGlvwQypTxaZZTQ6dyqRFz1JLhAvKRd8iQT+C7rGniQlWA5c
5YOXS5onQQ3g1B3fKwkupAt5tAaeF89m5fXONMb8/h2kB4deEAiLenpn69rQRvtV
VWjkRq2yl2n2d+6n+ccInyaBm5NN6X/Y0Ku3sAz0DwKKZHzeZynesGlEkqmhfK0P
UukDAYlGz57hOELtYZjZuT+RDpneD33X41wrQbExdKSGGTz7it2k+m3RYbDqZg46
K63Z+LGKqcdZnS7QSVV1vOtDhWKxxIcKjar57/RuqOVVKsEvH4KcQSvR38KVdVGG
8XNP6y7wN2O+NBH51JoMEA+ssiT70i3itlTm0ibgwM2xSb5rfHtn+Cene8q/ZiRS
0TPdvLCxizZSQ2OoTU0pmTpQyxM+1H1/110uV4BHAbyY4vXyOt4m75a/bt5bXklK
U/+5ueHWj/4UpwYOGcMOluMd2CrX0pWwQgtYbddfKrO+ryW8tNkpv8LwSW6WJHbl
YAGxcXvtP0jAe30L9rMHZ4gI6hx8sSYB/gqYpHSqmSAqCKH5lrcIFBjtskNv7kCb
I7XwzoLiCkno5ZJrrLQioDKTox7wVHAw1/pHkRV5P9c78bQRoGx8vqpVJgi+/Nt6
/F81lIi1zRSxK7nLgKn48RYfwGV5L/xmt9cS3FQ2G3/zeocu4FHDiZE8ymis4OS4
uYKYz9yNSiUCb9Q2/fNFSpOxzEHpMIURidU8uX1BMBRjg52+YwnuwMPYW9nTlcCx
zxMYnkF0BlIbWA+hOLWksBHmqyz1XFtGsslp3CGlKvbnVhYcw0KRo8Rmx/u1775h
coSwNrH5m2+fJLUPpT/721N2Obk2/YtcoerSBRqDsqPdwV5Jv3fwNL+TtmAd3Ryf
CRQj2FzVEIohrVkv4GCB8yxqmwgoY+WTdlA/IMLXu4LLzlfU2Dz0RTOO+azJvZLG
hgOLx14+evLtLc0SLksLOz0p+CEV6KKKPC4dmohNxl4G2poz+rtU8zJRIz9h+eQ1
x/YVCDZPhG5lEmW+OY1Ay57a3kxehPAN8cXjJlsE0Jrf3jNPwmDgat1u5+YqoaEn
oT/jKIUmIsA9pnLWAdfNbaRiqJEg8HRDw5beSwz3ZYBz1jQbx3z9OqLQjDKlGsYi
mR90JKhDzzooUsayO8RtDGHVHTLfBZLeyKk7/5vKSLF+oJU+0ayRP2cO0dy5FZPY
r4ibT3nZF6nP9Ba+D+gzoWpOh+gVOpy1vwJZ6Ky41NN3qdeUNFrDcCsbzSLZO67n
RLSV+PUXsqZERf3cs/IV3bzb13htjIYfknxybuIIn2bqP8JIMPjE5vMYE2B4zIuP
UafdCRJbBjYD32sCz7R3pzdD7/ajEaAqFwQZPjuxkEWHWnCf9kfTMsdcFxfTdlhk
kNGhc3qNKF+ufu82H61SkKZZ+u5mFTC5fgwtjt0dj7ogR1k3737gzEnAUWAzSFZP
RXUichJ8t5uJLoC5LiSXbKy3oepwtbY+AZ0E2XA+0/5CM1LuP55PqDu/5P3+Q4qL
M3zX9oSt/oPVQPuX3bF/CwW+EW9xh4KAf4QEcSHUbgX0V16tNU/Pq70WA2ELHsHm
fANh8BTXe9iU5IV6LBYtyZx8rJaMZ798+u2vJ2z47Nyl0/Qj9ism1nsjAgkTHeIj
/K8wnj1+datupAoPVPGddz6WqpcZSAOeJPVen82fw/DDDZz+VD/Grj6Tdzt8pgJK
TBOPZ6Ns/3GqcaRzbZdsRvKpzxynZIgPx/AYKB38Nek3R+RPDJshvSA6MGz+5RS1
TdolooLQKYt/5Q5Gnl+vDPmA/lGGM1fHgmBYkYetmZOg87NVTz/QTUmK9h9Kdqdk
p1V9rOCcUg5e82LACFaj8m2itk5bjJiGkUOI4TNFrXC0EtrmdvXMjrEJ36kBdnwH
Vnj/2g/4K0esL1pBB50fMGfgUwtGvclKi6gyNCx9pnQdz3ool3+9TTtUTlU9SSks
b0xvLtlyEoyzxBzRhiKU85d3wvQd8Ow28b41rqQKlkaMKQKVMAHwbnyoA4efuxbu
XAmjaFm3lIc2iEpbzT7nqdi5B1sXT3agpB2wX2eUDARynk/1vR1Dg0HMVRB4QObw
dBQ4+AATeSFQSMS9AVIs0/OYe4ACrkmGlNvkmK4eioJaShjEn3/hW84iDTPlGV/0
aQuV3mE2Y0b9Kv7AYAQHVV51I8zgFa1mnRSrtldGTSLovcU5Y/0uynwwJWVN8GDG
dS9qZxSCJfKrMTjBOGAHbPgLEeuFRi40LClvzO/fmVk+xyBOUjUJGjFCYaCwxJix
X4+Ai1F03V8sl19Fw9TY8qontWt3Sr70OeBX7hfZ81lxybG4P+vUZ87WDmtnSaJr
nOct7IRqhZyJkHn7E5LskX67aQrbH2xjhyKxqcE7XA6g4ybD7Q2qF7e3p0G8Ex6j
Te47p79c+sX4T6IgTHRghfoC5hPEgIYEBSdJDw2y3I1S3hMrM5hQm2VihJycX095
8wvAAM05+Zi3UnlXlvtN/bfCWy3UDlBZxdnv59MXEvza+GMcwKStnUnSUG+XxGgn
AuCCnteBwKJXzapCg1FZBWt0lLpeusw6w/U0utx+OAkgvIyFweBnN9KkFtJhMo8M
YaA6Y4xbwtgjEMLozItJlivFRpUEK0wbelxQZdvbBZcy9HCmoZ0Ar7AKchpaAKtf
tRaS3rwsU0ehEFE5TTKruoGiTPk7JFpcsJ+jr9tzz1+py/u7iO2BU6pCKLv5THL1
HkU18iagZQtsu4KOdvvim6rHqWSgfnGJLAV0LqsImuWMWPhbnzvTrLtJXM46G4Zi
paENS5rlS1QLTXdOrzlvsJT5VKHJp+EtD8IbhMIragkqUC7A6X/ZrfpfyChoMJPB
1rD2CR9KdEU2sYhk9My3F9G71Mj8pz++GJVXnbZ1N9B6D8+lJp3DYjq3IIRyVYhL
SdIX5fiqzqg7DqrYQKjdYtCqmm+WJbr++leXCdEDcvSdUrjYx9S601ChJ3MQpVFK
Pi20bfR4awO4rgTpevX7cAjI20dzBNppPxZeuaZikCGeyL+YF1ksopvasVTTDj3h
BOLKBH3eHgWIsSGsNLu0oFSKJdwBbyxS+v5d/aDXc7rTWWgweNCY0rPaByyC17Ul
pifX1m7sop+LqbCksTWs/PGD1Jiike4hBAHXlZqv5vZHe0x1MZbnS3D0eO0sHp11
rwOr6aXC8ZwUOX5bGUn/wUy2ffMPefb653lAoCzcBbYNPh7aK6nhiRBnCDSteViu
2Ejglc2QQyOLaaMkzAuIesg/QclE1NvW2wQPYoakQE+6gJUkBT/o6mAIgc+bR+7h
LsnnI8I3r8EsvnO1Vz1G58eVzirqHi5jaO439Q6F/m325VkHygFE63Qvm2Z8xaPf
nzH/kq+nrcThshwTv2A3IJa3vhECXyVofYY4wvPtVbSGgnL4WVezjUdrnqMIjgYN
pKwr7KkfYS0WdxEllYioYx0ROy8G2VFTqldPKdpusMGJ1u+Kg5n/xsN4MSht3ApG
3ttnSWCs6056pBGlhCjAR8Q+V79MNs6TVEqQZbat+kKGpUR4XurnK9qrxcR3/l4y
S+BzoYY+EqPCs1MgpAslTT36T8B7qLxk+VhAdbZtdNw3mhXqtUUV4E1CjpfwgbZr
LrDl5oGU4P5tolvTneSVEjtRmMj7F7grlr1JdiIrLHwoMUPLENS2L+p02sjpBitL
uS6+LF10O0OM9Dyzo5x6p+2khDFP/GPzIkQppc8Gw81tqsd8ItSb549uHPP49Bwh
XQhFXNtcMjHcS+OwaJPfxK45CY8oCTmPQxyODMDlwKmgw43NyA0WceM66p315qyD
Td1EVUdBn4jfAYseO9/jZK5niDLPjrLFkAWB0DNiIpWwmNXKBoBaGxcsaRfowU4o
niXg6vhVjYGjv1rBaPjO3Ppo43MkUxiI6R/Pf71CCTRZYFlTwuCawQRLYjHpk+hW
jGXuZYchksTMiHgvDq+qzrcO7rC8b8m9cuzwQrYZdbVnj2zWetCStjDWQmeA85Bk
FlItJ6KsVNJrMaVwoPxKtA2zLIyZYx/ebfGZGt8Y0p1evDAdYLSVqHPZ/cOAqBkJ
pn+ok3l/5wqHNcIKckWSkpYL3Y7vl+uvBzgybX6wPg+rrkCXA0TbS6IZoqH3NUL+
XUWMVQT5o3b4Cwi9Pn8bc8qgEb3z5puwmI7MyOqqGfLJ2lkwz7taa4Ed3nv5Say1
pkDK3pZTkL6BY0BBEUJpAWutGAK2K0l1wDK+bsKmyg5tfgDZz9xo5kaRsQs15bjK
rmDUC4B/bE+m7uuT2x40O3cZhSk07KxeBsuxABPXllSHw/eAMqODAwXq1mJamlUM
C4UKC/xp6zJlo9A8ruG+bdKlIQc60NafADqIjODVtSbfOUnfZeYV9zpc2nys68Og
lgdMBQ7ffaOciSQFi+B9fYZRg6BKPCwhXARRDz3Sei3RXuNRtApzCtSWto45b2ux
5MQbD4Wo2EuuKvYt+S/PrUeDdKltFO9f9x2Cxp+DH8nLW/sVmOb6z+QzQTi18CZQ
NEhYetRxOmxt4CX8DGZ6rsFiUovyfXpno5+qOk9hmfOU1G8BZaXU3O/iNDo8PBzq
cRD9NRrpvCdugfm3CyjNqP7YivBbTR/u64krNSzeMF0T5WGPAf8gyqzYT9dFeKyW
gPVdx5QNZmzS9yNW0/N/fj6Ln425z/ADwSJ1MRiaWHVNMaspIwBT8yIrAjqIT/qM
Uo7TZZRGRMWDf1l5m18H4TD99DfeOlI049aSUwg4CCWrFjLieZ+KUH0CT0K96qyj
da59gR+iRrxr7b+S7G+mzU5Kwhvb2ER+l8NVfxEL0jhWUvwa/dPfF4RL/YJutYGm
1PjjAasSR6ulbZNxu7NUZLMJdSsPvoCCcf0rl56Fwd75uribL4NxXPRG+LWn4H2f
d6viNPpCdj0dnQvLcsgno+a894dAv4ZbMAk4mykx4UjDiLicv2mLrTqWLWXh2W2l
yVppIzWnHm8BqbaRXYky8psNVtaGP22U5LVMa/N6/jnkp0Wl+OjufZN2L4pNRQMG
hPZMDU2RRZHretFn+IEqiL6TlwX5ZhaVYnG4YRmqsmyK4AkCjhqaN5bqUnlOKfc3
xBqsAIRdVEInqnd6/dYn0taFi4/i8SfVpR3HgiZxmsjd5FFnNHMxgDiZV7T5tAbU
rJqbooOiV8AbzoWVL/JZuMQ+JdElCZkry3a/xAE/kGokNvtrOKbCZ95dwHJDrZuZ
PVqIjps/YtWz/I1SKXNKZhpiit2c2eOSa+iPqwfOmaatChOizYnN03gbXqt4TtaL
MLg6zT+l1jRnu12D3qy7KBiiidpzda8dlm1zQN9K3maPF4S81N2Mtl65Xt8ULDvP
nUdA/Onse/JIzTEtHRlG/K2aSgGpvbuZDcxWI9lz4+wrBF4fnvX1toWd+15bLh3m
CCOuqYut5bu2whZSSjVLXqtU6aa9qYf9vZVTJMwgMDluqU+5iQxqTNTTA96fH6G0
q5n6AfpC4tYM3fZ5JlpPd2Q/kLr2Gla+QZFaIWX1k2+zW0H2j62Q0AGS5vzUZ9Eh
h0SbNWE68DQGKbQeWCEUqq5Z5rIxiJvRr2xdFcEsv7aBVKXkUuHLjUkxigmF6Xul
YF7riNuljZNRkL/uBMvDTqKSC8YxwZ1ZIKR3NltTsFf77hG0Fo9XbsKxat+1oPwp
jkaG4z9MOJxL7P20AeXrrl1ym04pjG0meqzc++VBJWyE7sLaw4bFoQcuj9yl2Dgf
qZyGiycqehoZ32+wuBOS45pRkljM4ypAeveeED7aBlb+JMTFeH767Ijbj3jSnIDt
SyNITmFMiBdMps65euGeakmD2pt35hcZqRVYR32JgwEgCk0pYcpLZLgYrpNoMRD1
fz6cdj5X8iJGrOZ+HIB4XxcaYwRzpwuXrZeMj/xZf5uTBQxM3me16nCzbtf65FpK
20Jx8CK+u6F3MwTFA2nbh0CeXCSTfmAq+iVLuLbWcDmRyVGhS7uF7fu9I8uAEOEp
FOfHM4/bmtLqy2BYN44mvDkxv47jIjqBAM/mtFC0/+27gtQqyapbKF3fnLlQ0EL9
TCK9VmdfUXnWhP9JJ9ey6oja89RptqhwcQRMYctu5WB4vSyeWdnJK5VYXhsqbcfs
HJ1Gg75kJzKX0pfyyFF9J0gSuXbozJ6abJUbV+xuaBbNgaaSV1+IFdt7NFhF6iA2
Dc2aIu6suIeA/LE78WeSM+9M4jyg9vgjcePAnQHvAbOMq6WcxkswYXe3CpsYbjRw
VIVeM3MRiWNnNOmLB1o+pmXHuYivpM5c2SSMIHjmgjPUNcZVuyDTM0wvL0ZPjU4H
IwI8lVvBL0+2Wa0bgJfSoYQxIy+m+uX6J1aS85X3A4KdzKc4NpT3a5SQt1/1eb3a
aE9gzisJolbIxON8hbZ/TaOgm8Vtj9bbj36x3gM6m3RLAdAyBtsLN7H1f3ip/RzS
2/VVe57cdzElZXF1GK52zFxdLFyvpyVfhhcDpXbcmwPGOSsP5Y9Eae0nqbXSbFCh
3vYE+thKNsZj8XhMC7Xb1ASLnt2WLe9La7BF+brGjqNHCyJxNg8J1Q6v58jRJWxS
UCMB62UL2OeJosbNY9kOPZjJOMALvO5VDUcncrUEvZFd8jtKblH4zjp+TZVWyzuT
kXeIaiaUWpaAvc7xjblQ/rHUliniriqvqdrKicQ3+pq7Op/hdkQIr18o+hkrQ7NZ
GHqHd3gALfyMxtPxkX9xIwtM4Qa2EAY99uabyPx6viXFnXBYF0c33yknckKKtGuU
VdK7fD5JS9boCHKbLH8cqKIVuxjeMqgDjcum0+L/iPZFD+OXW0kEHIom7WrZQpQ2
0xj+YQZkYCco0L89VCnuvUl1hoXiNWcZ+dsQO52ytzECAzhrIYnh5OlqrAGhxn9P
TKab9oGxe46qp4XKtR5ghLM9qCQGfcdenPGhkVqUQaJv8NNOf2NyxBRmRtetheqO
RyYhbhan/+9tBbSw1wrWXLRtwbE7YA/4HWdftcNVOwLAr09wFOQsVQhVxatGVNhe
bx4SUaQkp6cJ2DQ8M7gHUPg0E9OAbpeOes5Y6fkKe5Ki6vhG/fjwIFrf82+NcZpQ
Ge+qgXFQoXp/26jeJJBZJ477J3F/iumdMzqEUKPKs8U2i9nvZ/oxyOkmavFHVcD2
4UElVyYEKJjICvevTsS9s5vh1hxpRHDg13vC6unc0GZet3wRThwZmSD0ncNFjCjN
5deEWv4+vEN7sHfjy0ODaqn7m4FhThWYZxiZPxgGF6mJ/bLQR6vvdnNqYaRr1Yz5
bApmyxzhVS9aNU+nBJftP9UiQUkRPTIuK268/aUEWh5a3tS7axxfi4WmUxJKwCDu
tVpC/tzl0YTSY2N40vuScIIcWpcRe3spdSKqgf8bdUfnGeYpEhzj14B0GEhyOpcg
3d7IJaE1HnQO8+zuMUTyjM4+RFJvrg9Ejd6WvK6NmJJihgbU1LxOGYl9ZxpyHKkW
EKX3e6htw7FdUqQ3JVRwA5falfrnZnguNb48b9MqEk9+25LSo6dKoTevSmoOSs30
27uPKihsmc4kQK3UqzcJmRNkhdSL2fdCFquzPFIsLWTKddAj25M1xvy5TPaanvQe
kElvN7qa9rfQj5R/+BKDvY/uNEqbkR9SKir5Qx2KQ0rW24BiC/UkM+7M5g5ppKYQ
SGCvg/S+oXqubvPLcrBgAP66NtDjQJI7oqus8HgN+/RHNe7BW/rtrBAZ9dsv3KRN
twxOm+TOhj/dss/HRSGLYUWV74YBuTXvYUqyQqC5r6EMdYcj/Z/EYHUgu0pL8Xdx
0jLZMQ+dOG0SVRfn0ZS6SYpOM5O+Nhh/943RUgNNHg1kAwlnBGrYgw9AvZOf2CRF
hekvpSXMr12QiLsOnmNMJPqhKUR8q6XwUx0UU51upzdhNfEodmMBvXKVrsvtJk+1
/kc/TJykVW1Z/0hJCIgDsoOXNvpu7dycFe8kLsd0k6TRUJ6Um6s1Dz1d5z3LF42C
5YBiO1r20W+fNhB0SLVh0bMSU/SIfR+pBO7OvEyU1cTZVZNQdYiXHm2In8pEXH5T
qwUKISL/Ust0VdP2Q1fsWRiZdDagyAYRUf9ZXfRj/RJIA1aeXeXqHZSECwKDw13d
QLCg8QG8Fk6f9iF5uuZjIgotb19rsxPHBzpv6/aJSNJ4/4ADpB3IS4wI0V0ZfD7x
FrEY3oaUbIipiZtEBZB37fZ1CfJ0WqsDc6p9X+ydrBpRFBztQzQQC6UARZoBSbwB
ktzaSC02zbEgmAyTURuEdIUM4WNFOuozioaMx6dxXsVUKTLLNvN6XoDhf7hH55pg
dYa/Qff49qRUYWKtyzJ87sbnblkAvJ8AmMI3RPFkqgL/kppaaT6DPcNmK4JMb5yS
Jh43lP/w2LUdY7WeV3LhI5pb/weugBtgPhpQJzEtT2RqPEJcjfPh8VLcWz54xQAj
TOrN41/qp/hU2xy55pYzy+WkA2/CpAHBhEu2QePC4DxCeiHBzwdAZAdNLIePOpWK
XoHvb/EEyG7d/Vgg/zJ3c8v/0Lm1nhAv7SpXeT/IZ6C9i469uOflWxunNlUW35lD
uLavXtBWYsDlEuK4C+4fnYjd8cbY3kPwjzMFdlmPQMHQdmtpUs4Q/KOk8VA5CGpk
hoG5xSbhAR8TbIJzBfUtRbfX4MSlQ2xs7pC7VkHd2Rld/mfxKXkyayZrift+DPeG
0VshiGgJk64w+dVhS9ETSKJOPE2RxShlh8Ut+DMPQFmAVlCzPqjzcwphz/gXfuxC
FefRGD3FE53WO8U6Z8YRyKabhWQJOfnCTvdWww7ZtWtkm46FKONmrlh2ezShfKI1
y3GepRHnp1ZEgHgmR8qIMJq05s2RqBjDZXrt+cBI0hdcHf5n8zB0SFsk9i/dVxhu
baK5FVgyrVlP1lUuE5a0qaxKzTdaQk39okI4yodUIXGoliZNXdHtx0EREFgO9T6c
kqErYTQchYd5g2K4RjQtzW9TaX1JQiz1VcGH4lIN+953EQqygsZMFxnX5Lel0rXE
vrk7y8tNQcIutprJkRxYPrseLu5FGaFFCpcVQGPTiVWlKo1rXBbtkwskw1g5X3pb
S6/IvwTBAANnF5WAepW4MlUMbO+cwjD+7Q/cfs9AElZRYx1kq9Sg9jxRH1H6gUf1
47LhXk37NDxHz1sm+QUmklVk4cpSHErTdpNt3Q1QDWihhglP+WqDdk6dZo5ctD6C
lqy7Z9u0Rnfh4DycCDoeJ4GfUuLxcCEkUNoMS6zhFbmp0C/4GHaPRkTsdKphn7Xw
lEcsejBzd+pQTKCu+x4ztck4rHzi2mVd+kqJYuP+BlFmwRofHdveWSIE8U/jVvzy
UM6F8HpPw0teWbhMK+A+wTbErHWFFNInUrMON4d8nfnLK3mUeo/fLL7zb9w8NMZ1
2NVSR3O/YKDeBFvgJQAq7vccROXDieariafzuaZ/57hVA7vDVay/W/4aWDA1HBOc
0CHZrKr03GhB9kaesO71sw6InVFqwaAjucXouOjmGz3C+JLc012uQOH1RIrPoaC/
ZJ3OIxh1dpQW1lrsq/9x+4S5Tg5OQekbrwoWtVXT72MM9U7Y0X7dUNF0b1hPM9JM
Kg8rwOGn/yFk8lRvBaSgE5mGO3re2F3kf699lwzgmRzf7/Ld3zMXGWxEagEc/Sw/
N1GeytxGxlfY0DLajjXZNe9Q5mn92Bq6ycbQna/AsuccrT2OK2RPb3nJwXf3MBbP
64sdR7edUmkuygAdsurq+kP4LSOhUCQR0eqBxRdY/ruPGWvySLb48BnKRtheuUTv
6TYbZFhc908kgZolZh7XfA8K6yaZC1IVf7O14OtflybUcjCYukg5Mo5jQLz2bobi
cC8iQioxyUi4LoWYhRitVZJh2sacbbTVU58+6Q0s/7pgCNDp1kh8kDtAJ2QUuo+U
Kyq+6caxjnX3oaON1THYTqaL+UcJgbdHs+sWm07sSQaarGJvNpmKC/oZNUOKiS1r
2uyoOzLQtoW8uJEpRvRlu+I2LvvgQCgOJoi2XK9EOhiKggzzDvzyy+L05f0uWRDT
9af11msyxTuUpxMUFyJOhpLSExe8bywmxQSXQlBqbTQqRJ01wIFfnAUw4b8C1wyf
65wpNtG14NMHpdWzoIsx7WlrEqehtWkjBOBqp7MzHJlXlMP0Euk+JaTz3PKaTifi
C93HWZotNgtw7nBi63wMG7hLlfF9JVXb0bhJomUwYPp5vJ3rqBTPAJKpU55VK80X
eCVpimC+k5p1VKJh7sb3OFgd3uu4rqHqQf9lXfUIvng+5EY/nTb2KB4TAtn63PpK
dwbvvmDWnuNvGNFfL4nAF4SvmQKRdG+foAs2w6SO0zLBOQsz9L/t3JnaYPtV5roR
0PrGP+A+iSLCvJw388XedBXRePvWM3wHLva/9A7/431RiZqBhmiVndjZhA8VR8gO
BEmCImXlftRzJmVlOdMaLS5TWlFHzMFi3nVAYgt6NIbvAYyUwPucjVwtU3HX1ms1
eJsmpnYfXs7W6gXyMNvyXE+zft6210cSAW9Jiav9jY9Yuf/aizY/CehALid222Wp
+2xTFdiTYsNyi5mj9QhEENp7xOrPbwzxXn8csxlzwsgHBDIxKMw3WANXwlVQ+Buq
toFD7mOmT0jZtjGBGyCzX0kHh1EXnq3wgeI0BKpQlQqyM1o0bnEfoIMO9xDzRddb
2SonFVmcbyH+TqplUed98osJ7Q97NOep+fZFp0SPX0YlMrvvFL2nCSa6Y0YaOxac
GBWI0QJyopvC4H+VGIO3EyUSCJfFcqD4bSQn5koNUw6Gg9Q7I4MWheBmzC/X2rEw
I6FYXKaM3p7HU0h5F/gvrG6WgxH8UaMAufV/wifBBs/xI9+sx9H1T8IYeZahWbwj
JdyDgy1360VfV9zXVPDIL1J1yFEstTfzGV2935J6GsWM/Hucrtus7Dfxev77Qtkl
kQpXu+AkI7XkAKyMDwp+g3xAOAIVW55gY4n545mE6k46RCet1vyDv5LAk4dLgPRH
TIWWyWJCeShc13cb7XpRrpqkK+4mQOxCPTMQabxjfwQXJAOrc0tQOCPHBY3xgUCY
GfimLAcbrXXrLTZp8VjbmxjvVStMLClWVrH2nvuod5rCF8UVY+zUVmQQX3mWJRHz
r9jatcAE46WR/lFJRSeZAeJCiaxVZ+uA/2pkzAqT49zw3gb7bqUBslbGe4FpvUi2
0R4p3O2EBRmhk9vEmMAvUJwMaVEmc2VtqJXe5mmBFXQ4oENAjmV3Ii6KfsXD5PB/
j5Afh+6qXCTAvxP4V6v2/+dHntZo6Zxl2O/FnL3Ilf4lzXS7kv/4hdd2+bAa6YWu
D235i75oIckbJcfywxm7EX+gldnUHVD9LFgZ1OXLOuKzooXhBKIOp/0gVcUi+Ub9
Z9VnDbK7C0xD8ASTv0BBXnnal2mULgeioe4Z1gHk/Pb/Tlrk0okW+Ol10RsTGN+0
aY3JsDz09rqGw03whSP+Cq+LUZuRpcg5wAIg1ddeUI7Vahpy/O1iQ+GiMLAwXP8B
CBxfjJ6sO2DIEKIh0QYxca8AxNDd/9Mgb/tz2EzXsjAHdm+VYZ4SVCbnQg5ZXGib
LN7hOJzh8vJPXYHxIm6oQ3PNO1V86Zn+iywYdYa/XsWwR0yAkyp9F8ot8IiL9WpU
C4IEzH7vOfX5wVB0NDToDTe53lpQF9IfPx7Djf5aIXbBWsKeXAJZPHuahB5SHKzC
mka03MXjprxcXi+F7pXpx43JWWv2z+B4UXB+pMjSQsmIRcItPYK26iqcd9nWJXBb
Wykte9EJzR82NPaFkvdV4opZnWmz8rjPsOIEpJAXdPqRwPSWP2331k17zlxdR9Aw
2nM8b9g4uj01UCwEjTrOU67koPNhDP5FceX/n/8nrb3AfxpnIExm2GmaS2ExO+5f
gUuyJs4rdKQQn1K8QlvfQENr8cmvh433WWB8viEVhetEluNyXAWDOku4OnwPZfwx
ISEeA4gHkLhYed1QeFs8CnKruTl5ch4dgiFBrLzTojh+QgIBmmDyFy5J/T6gYCk3
aD9gViHNvmZkQkQEyvTbxOJ1V585M7HsQKlwphAAsQ62Xe7WhJwfWaPLzU6sjwak
wrijsEeHg3rhD71BXTDbQa9h3brHyIb4strAsUvko4NRPxihVU0bSEJRLKa4mIaZ
rb7q1KeRJEfOcIgqh74ary8Fkk781UOsT6Ta7br4GTTojas6fKtwC93ZLc6SFjct
K3p+wQDsDdIOoLnC+w46rQrRRQLVHLTqSghJ7pTfk5SL0BREz8Tt/XvcWKwx7v77
bXcR9Cg2jo3vc6mBv5UXCmR+PZs6vzqNMPtaCCzUFZ2O5MPG7VpvJLbz5+XRMDhV
wsapCRUF0q49C+GM9hrujseXOHdypD693hUNOceYenv3HOKUYlDUIh1adBIb9nHY
Phh5jORsNPEDUE/t1CkeLBuFbInNHdYeEMW45dG44vUIjz0BbJ2XN0JkAETvYmH5
sQVMZojN1200i1mSYuox+7KpUFPY8V4BTcZcveNrG9pbXx8MdSRA5QsDz44mEWBk
T0nZ/N9NfTv35OaZADgLvr7pSEEsQU1OBmK+rxcZRywl7arGBlOvvzJAiGuZ47Q5
f2WRjuhRHxxko9zFhc9jeuTtileMaCLuR3bHHYEZMv6aZU1gbgmjRliOVmuRvx8q
lsk3juhv6eK2tbhBIazmO4nfVsSYw4c8dsO3o4Jt31IAcJOx6tp1xqG6lbXlgeKT
mIZHqPoboKxQxkygCMP6dQ43PxambOf1WifnmFvZubZVxhB5MAqKWBHUinYa0O8i
L2Qr8zjjL51ZgqTh2e3iwkvfSj47amoWKQbacXj47pcJndwdVQJQHq26KjJN3WLr
tRBxEhB6QvXe+r98Q6kQGrwXnuSZrxjriReSl3M4poqh+aA3G/P0DJ9fB0EaKdsC
MxEUJc5REbR3VlL2IfG1AsqrApqLDUxz8sXjIu2WOJr5WrdZJpth3FLAhhEkMrv7
QTPCoopbgP7vVsvfRjLG1fomru9gaMDPXx+eTMDAqz3IWyt6rFJbZAFT8nfNFMZG
3LeoiDjZJD0PNxQEFZ4OOvWuGCxVU/u1gU1G48AtRo0riIFW2Q0Ml1RJf3OV3jrH
KaYOLrC/vJzrxlekORurpZ8tqSCjHDmJjJglANwpu8bYnnXKF8nu5LvzTE7hhqje
x5hnnkk7c8MD4IkLCqyDD285BGSLRh6g1ubXTqgGrIrq/RcXvxJY/Yeu9bVwJDKA
92+Vk8BcoHJBw0+TTf3dEwRPRmNaSatj68yBexuSoAxKbSUVlKu6d5jUr70gvQuS
ezbGYAKpxQDpGeovF12066q9JsoimpL1nJwKUxNt4JuGuE0FzsPBDy7H1mu+uz6b
edjglDOH5n94kLnG/Krg0LZQ+PIUn6rfsxREN5kE3FqxpIY3RljylRtp4hClMfEi
CE52nnWTtFGX+QAe1G3vAS6wo3KimnhNCaurA9ymAedNxEU7NpFXqRSgN8Ynq1aL
7uT17687B+dRa1yQTatlNSqVVlRbalSs67HB/1jTUTvrSDhujDAO60Ct7wky73d6
quAS6XPA9t+Cv8yntUuHhjsHsB7Vv38zB2PW7QXjYIpd/HlFkZEChQJClW0Ged6N
exFH/G4Nv3z6Wy12tKX0Yq9z07SYqX/YQT6SIlzk8b42KBWhgpz+517YH7I3bjKo
fW2n1nJEPROj6moIzm/TVJFe0ZR8Z6SIsTfcWbup208XQm04WKvmzz9JdXP1zjDD
JP+A5UGk3Hn3CuZ+LM+UDS5FPaUxy3b6JEnhNjp5YAF8AESCaKFC6zuXt/3mqXEM
lCB6/eyxAoPVYNGStMjArzPOQ+go5po+pr4y3rsMit2ynKZVUmN1Hd98HzHD58vH
VS1XE4yqlk5+lY5rdn870njwEWXyUHnfvJ83tVBSPmkPs34jSseM5dfxvmg63/aT
s3ZbgL8xG6Vi7kwZXYZp8PrbeaSkAFIhMxiARpljlB/5XEca6ECEq+sVLgyTt0l6
sOfw5tW2IcuhKOX0xALTMzAKORd89OYlNtrof4hJhTmZvLaxoLbK7MHB8TVbaD2X
3VwsdK/f0CZqwyTHRTH9g+p+OVBXkKMgbSdfSO3kVBD2M1b0gQViag3pjJpfEEZA
D1HR7sjqr0OrNFNTjK4jjnQLEtXJ5wT1ELcViQhfHCLSkDq+I+QkBIDStmIn/HSM
qKgUFKJ2jYjLp2FoV+JXIpvCv/YDvfjgL+9fYraeM1rUVogDk73LBUipKcTGLpSW
RFLCGs7v1DC5IeWat1Up3gdKAH4CfboEuKwVC2kiWfNNP6FcI8nt9WaDoakZJ8oS
Psvor3bREEX3RKfKiX0NCX3Z5Rh7wGbzJ+NEi6Ccjw8G/DuRGrrOixo0brY4dNo8
mnSkC1nANKKSMkPff4lqaPJnz/ZD8OvLyRRMwOhs71Ii440BOw2CjDusKG0Ch4z/
O/boF8SATa6HLHQMAeiWIAkrwTuFKu0CFj6lJ5/wqjUEAdfL4NxRwEYRnco8QaoS
sfSgjjhpyVxeY7IBhqBB/a8zITxbJ7m1HzPgTvNj7coMMoOlZz0LTBndrxRsWJYw
L4Y9dTj/Zj3MQGJulDjJgrt1BxvLur2NCFBn2PlMtp9jNXJXJ0ZylLlC6RswnODt
ywXzL2GSnPmHvcqw8zhT8z8KTh2iLwicFUOPP2W+dfiHnm6ZzUZwuk/1Qj8UM4Nw
uUppc5JKTfPD0kzFAULxz0UU9OeEC89ZfkpYye229eMCixG3z0oIYWD/4qeq2WU2
CyMPpDqyJcQjDNTKU8CRxnr4oJ/ZV6gSh3UvsF+5F3WHlWho02xT9HVZFk/qPDzr
7drmyw7K+he4/jcuLAzqAsKGO4cxoPNYqnnhmyxPC5XO8yx43zFOdmm1hDxM/ZrL
MZbvuPc50BJFK7QB1N6YhWONnJz4r+DX8zUS70rZ67e9aZUs5BKNGVmLfZXs2aHe
Ce6XUkAZl+a5w9/ta5ihUM9FCQb5Zm+OMGeHxwIErMETYD7513Rk3jE9ZFIoUgBR
U7vy26ciat4aSYlxzCJP5YzQ/JVZ41qxAK/7c1962K7Pmo9yL/9soax6ogqPEb21
Yfrlhp6Dgr9c1yQcplSKKJ4qR6IccG/mqkMTloPlHHrUPUgtQVp1RCr0jhdLZAaK
eJ4XRqpnyewmzag/y/L51sLnpVbNgetmaNinf4D6HMNaJt8AEwQjRVd1T5RA3mmo
tJw5idobKXojtaU7GX8Ex+AzNFoCgxIERRpo0ce6GzPeYKdz8LBP4hwGDt+Wpl8J
MeXvMcm83t6yMR14XzQgR7ON1fFBJzQ9ZhGtHDmWRmYNkJ76EtaJJU0ztvYy/s1o
g/HsgXpcCzH7fRPxwI9AoSAGYfGRW/mC08SV+XyWQy3t3zLGkqzWUq5kS3X9gvb3
VJfSRzBIGiCoqinRp9sGp9rhDSb3qc5anijlqOMjGXkZMGbqaM7MP+98NwV6GG/p
hAF8D3uKrf+vjtnBBCzNWqq3vuJcR6Zp1SKhr+jIV/YnkLeKDW2yet+kd0sW46yY
jZXoNeNa/KDtLjtqtOobQweNeS1Cl+N9UhV5FST5JW0LTGyRKXglefGCQ7SmHT2X
zPUiBz9ZRzMCP1L+7SnOa+sZz++wwn3CSGF+yxb9owmoOiFXe0qTjwNsYprDLmaU
x4t1LgmdTNPT37gM3bK77Z+yUvmh3lP+f8Yc7+WosKBpn2O9NeNtnL90mLkewZ5R
2J/XtGAzfCON92zbS2rUI8YNa1RLNinN9w4tpEsw1KFTWlIwUvxIuIUC5fSD+0zr
eWZ1bG/cDX5DH6AjaenINMY47ZqvhYiCedHcmSsrHyEFMEcexf/ZQ9rXCRNLJE15
ERVAvQ4vgsR4vnxCh09MFdqNPkgI9ueGIP1S/oeolowErZz0zU30cVGxhJ0RmqgC
WgA5CL7KbSmLYUsX6kZPuCwUIhzlf24zlyP7WKzhGQd17ukAeMjXxFNAAXrOW065
P1WoE7fZ/rxmjwmThDTfTFhYCH1qrfpX0yfvpkLTN2qi483OQIzPzB9/iCUdbenO
lt9PhPtYEsPM3PUbhNhHlha3mrvvMVyKquuhZAHg9YTKL3XCn/ee1dXHBuBD77aa
Ccsv94Hjpcx4jxW+2q2zAEFv62/0B32whipe6oX/iEISaBpikqmQekQ3ALAuhQmP
1dLRM6MSW6EqmNyAesNidE+10O/NtiaKSLlFcEjCEzFlq1XbdgvSSsJtiKNuAgtR
2Gf+Q64chVqCfgzXjYNtxi/t6CICJ184E8Vyq1NtfQ+7P5NRG02l4N9Duu3tO8Ln
RauaAm0y56GGtrnodmzKxsx4glXZ8kw4HKlG4CzUe4BgYwMEQ7iWs30wOEZgipMU
yNgVieGLl67bC9iwGmV3l5xr1A5eiAwXJeqTN9QDH7i7imzJGh8dBFjt92woa4uS
NsvJOfJHVpm5dqua43nZI7e8MPlLoyP1EQaLmXSXJ25SXBT+jMs8kqHvhdh9HAGy
C/mkwQ9xLzWZ9mg6aBcKsa/S9OmjfhYgIQRvuBIfLu0RF7cwDZ12U7Qi0op1ZVDS
D2dmtAtt3tXVQjw6HG74DlycB1QJgO7MD5HO09BCwxng87cQXriaAJQ7fmnA8441
ZnanmX6wUSPkELKy3AFWpJ8/MdURh9/74tl4kJ01CZeFnPy9KHYCiMKpWsPJcGlS
pm9TkZNfVtfEixHwcdarJRgzJ0A3aNovqOJMABDGQ1dlRHGEQ0O5ItOMGsX2x4i1
yVzkWAfzzb5qK/OZ/0E+HUMH5NYVs+Pds43jt5+nIRRgMn/U04RSdgZBHAtOE3XT
JCDQkgxfezCl88PCRIrHvAGVCkDMQGFE+8PIchagjNUX+W8gRpIb8nwvzGNye/tG
cfIKJeyqCK3MyjAxCJGRS5a9gS6T37E9XiVkaMbYOiAbWuRXK720g7DRpRxwBvxl
Jzo/P7SHktenR6praC8X+9qlt+2d4Yp875WIsqFuCoXZG1IgJ9JhFGl7J6mxwFSA
b0v/V26iVrAEhMOs6fO6Fi8wNcLkltigMF4X7laHecc7tNSb1eeoqOSqYNBscAQJ
daB4GQL6QybFcJxrndR0gWL1zvoySR/woEdMqURO5hwlhAwnVdb0QJngCe61aJuI
AWj1AEmIkr7zY2mHNwS/m1Tp22ytqXASuM+Cyo/viPlOxrsA5Y1pOerHvQpzBHvi
xHEwVnBr82o1zcmGTZM8yq7xLWFaKLDvFvKq16fbTJCMyVMna6kYi1XyEfX5ncVp
3BbBsFVBrkforsBk4DbZpiaykwMLxKkykWWWzZ33fqf2DtbewECgjIMZQFWjBWlI
nkQPoUYfdvGKWJrlPKNspT5fjySuCwHWYIXqs/Ghy7jfwIwnEnr71xKlyWxuHbtD
HQ9VWqjO7y+wf+n7eN2lxrQtYXWjS1KNhN1i3/cEn6ukahaGznTDGDYeukzZYahl
NAePD1d80lxnfdPkykSeSIIDNlYUQLaLwrVdqiElZHL4DgPDVVtCDt2/7XX/L336
Yh2K5c0bG1jljOkUsc30qJdRvbCwisJKc+MnSd88UiLazO1JrV9G6c0lQgq2ncNE
/EJgfAjTN1Owsab0xd6XKYGH4xyQENIUcU3sCUZNV+9tCPz1PUHg8mdLkhVpr3So
fDSasDwwSQWSYpiwapuQMOP0dnV3rNeglLWxHS6L7T/ps6T04G34qd3BCuVbgiu8
OwcOam7W9QfxVdpzcah1pViEk5r4hY30Lb+MAqZvMECW3dyK9W2pTkRgAZHe4x6J
lk9MS2z+jvFdWU8Hoo5jbyAf64tr4YmJj4lHkQ6I5XS9ZeEaeK6KlGgTfl3bgfgj
t2/r4d929q/uBjy00OTL5mL6XGvLKIWoOXPMBtJbMgsLIz2FnYEy9RQT/oAo291M
g0hulTB82oxwKwtm7SoTg5eJCmDEIlNY6celYKw6nYSqtaVzqNxsVLj/mOmZ46PN
Xq8YfwshsR08SMz+Ot/R2Cv4skzXSykRXLlfVkQWA5raWFQT1kh6OmK1+/Acb4wl
n9TofyMRXf4QwhPLlxQirbCBFA1bn5so4oXrk4ejF2Kr9lIDGAk9j3iwiQ9UTmJT
jKHzbSBhpoGbYIOMovhFLwaB/ixEGXjKMRsTveJI0Jr9wOgSPEaMEEofABnJmU8k
h3E75XoZxobShYqjbof108Ncp+IjHDHydbZBYygqszlm86GgR9mwe9xImkR4nvTu
TyPD94f3z4l60xcspWD5K2PsMBPEUh9XWo+0fIVmJmShNOr8FcpKYh7R1PUUSsed
e2GJK++/gZaDKgy09M3PjWIP/r3Hp483R6157HDfy2PbkK7aiVDvriGCpcBhNyZP
uvA7I0P6oCDhhHxXgRsjIhR+Kc1g9QlsBGu2Lz+dNCKbdowFMQ+a4SS6rUarF6eQ
R0WVHnsy/pYmq5sbeE6dwg/qbiu14GS7SsckVOGgKx9ehJOtX+PY2mbmzBAn0b+2
JpP7cBhXqoq01iv490fLGzGcvMjBE1FVrgJ8EgJaYS2F/rvwkLkeF9GjKlqBCMTW
ylyVYN+XJfKvSEkZokYyZl9xpHg67uYpSs5VeTZzj1Ro6gKW6JjYFw08L9tdP0lZ
jR7toM7cLjAjmY4PfhyBV1VXzyQubcWXq8kGP8v9AH4nGw65+DpuxRSWrLX1lHcM
40u03u0CxmA7k93qfLn0HQFMyHq/0U3H7oDSOuLEnjOAw1PNrDzCoKU/r/L0Hy9g
euMR+bROqqa/TR/ZxrXq93I4sADrIQ0OqNb5ORJ9byb2HV1xiEgOG292G4C+zD04
ObQ0qb4xF2pjIq4sf0apcWJopqByPXlNCxAQFFD9HjlNj7MWrIjz46X4ynN/V/oZ
3gKHu0NWziez0aC6jsoq8LLiXJlf5RYk3PkPYupiB/fSPczay0rfhQoLWm3l/op+
MlmwUkgByhwWK19w6DR5PwSrszQxWVcEQOn0Ej9WRJOUMNWi5UjOCluqViDvI9U3
6kLEfUiyhAqq6cJGD6XxnDIPhQoTvUuSuN3CffmueOxNPtsSP8WbcrKE0B+vqxXC
al3KQS96+tgyH/3Qv4pBQLx1sptJA6IAKvPTImbtRGKwqLGLC7Q5fGFhLkQPPxkv
BgF7eQSwCo+7jWLZ/P1eUs6tjPFuq/4QebDtfWGvorx60W3aaGVR+GynZaxJud4A
CIEITQbf8SGjTCwW/C3haHsKL4Tpye7IyM2AOMb2A5E3keWcYcyINp6DaaUTWziy
Tr3hTQi6f+eMckHq1vSImiGE/KcvmxN2cUtt8POr/bS33pu+9XY/gdki8+kPk/Q+
h0shfKtCylzSlYxCYOwPedap1YHuwglfkv3k0e2ucnJA132X0FSr1r2tiZ7y+7gw
c2iDPgrTHI/o3pufGt/NZMVITD3rSmwG9uaKxGP3q4wTjibhYWC05rBASv/VFI+l
wtMf4C04Rb9vXHnJ45Fg5XwU7Q/7h1FJwdN7QeH3pGX+/D5lhC+OddcYkUKsvvL5
7YhERl54cPmqIGEIMXDoujFhGMHvTuSq6YhoSRveXxEp5GVVw/QF2sWss9Uoq7+7
fiFXY6Z7sWNGfv4uP1fiUyVe20wzSWyM+SaSQZV5rdtm3gKE7TjmbRO1Zc0uPLoV
gDcEYqCGaTz9DazegZfUr08/agzvXFGcITPONuGUjQhTeLzvrwIeM0ShudSkIPCB
0vrZK+lqW8HI3Ih/BMW8n/Mw8ethVM2jxI0ejSY5Z3eavbN4AXTRWwfhqKXaaGC7
h6z9N97w2IMVMDVQyb/sjzZE8+c7qI+H1zvln1b9oq9aHh0lxmynFZtVEI5zYQI4
Eho75F+I933dN7JfNFJRLAP5i10Lzllq4rk+ZCtmX/nKA1nthxQMRsTVWZUNXGCh
Z7t2SABMVFSArhzqSUHaMOLV3nGk41z/GyN/kWQhpWt+J22zjCSg/pCXaH9Uc/1v
JF4TZy7nicyoTFbNJU/DL+/KKCDsA0LTSGm4XqCn8nqpwg/fugZq+4P4ncQFxlrO
9EWLTQ+P+HCFWsi8a0eB2zU96mE03sCIOSXzkYpLxPtpvZchj6ktKF62IKh+F5sk
NrnHvfmHNZbgeXs7r4smYo2lHL4EYfsCFPjlcv/6o8mPkRkxyViQK1vjecESuxdW
xwXOrbFdBVJONWvKbuIfK/fxlWDJZVYsA+Rf+vp2C9Y0xhFrhCA9pc34WeN1c7fx
GuqANZVjxnp082zyJ4wXkUUeDnfSq5j4Odr15CAqxcwvkb8EMrLWkoAgvaKUHE2O
LbZsjejIUGS+IPXTzpuEMR3s9BNOxh9D4Sti3Mn1faSUxfANbWNcaKGP2N/im4iK
314mxBKVFfEi8xJxwWL/vYA6GwoqyrTW+Ux3VAmZO02kQ/dHA0EEb7g2FMeUizdt
r/xCVOfl7UPG1i1WBg185XcQhY/fzKjw0qk2O0zdGZo/Ya/6Ma/cPYzetzPdoOTY
hf+6lczp8wllI2GTZK8cLCUgUxtuBmOtUURO9KdSJFW6l/aLbi9es5F/R9h/Be9O
a/5rBMza/8lka22b7wC0nU+189p1HG+EwoP5b5BMu38xBKLZj/uSl9NtYAbBU+H+
aOY46CrcDBnr0nTfXquNOASLDkaMUpQ38kIfP+uYMNqdesO/DV5ontjbEBEfj2Dc
ASyMAHMlwr26UeHDKBLEOxvsHVYHX/8T4IGogyNh38ETQBq4SzRmQbgef2UDv2tx
7D3Dk/RKf/QUFZF67BTFFk2Yh4UWzqvG2qVEwA8AMGv1HgIgZqI8EDigUa0oFP9T
ZZw5kB+rQb3FRa39XndZjVEeZsDZFoNgfvJ1Dj7NgIddh8rOL48OXu1mh9Rd85V+
oglCvwx0+RrHHbyeNUmyg0GfnUd0MiVflrp8BdAd7rgqYX/13pOFDFiD6mmlXXkE
l374M9uhSOAERdNTE0xJtBerRcg2bDLf/wDpNzHiLjIfTiQVUHpWtEjB8iouAAC7
wk1mg9w2qarbKOYu1gLINoFsVjzzxfHiB+/ylfScpDT3etzqubI0Mw0RdRkNEWZA
o1pKXvnNjg1kW0dZH81bEacJxMJbhfQcuNV6ZUMweQP2osPRX1AOsOi2bzcon42j
9bQOj6RsgpRp+1Ct8fqNHvLQBVNeTcOJdM3ZtLMfnWawJLBVWL6k9s6DIPQpV73M
Oz+rSQVor4paMeanTi9jtr/6/OIMYwMlI8C+VJOhq1zxsGieViF3KCplNI5h4L0E
JdHfx5WD02pFFteNTWQ6KAd+TjunudnrRhO9lvN6btGq+1gu2kfv9+ZHPMLCZYbo
1pvcuV/KSLOflNxIrNRszlvu2xDaNMM8jfxYwrpJmsdxxqnjelibG5LlCI4dvLCi
U+IPx49d/Y8vrd2Q9S9BEoFIwKVBMmqDnB2B8vEQr2z93UKF8vdlohcFAZDvQzRn
Q4PPVHnYOU2K6Sto1/DDpf/vRq6gE1uX0pVnSuP9t0z+F5p8woqjpyjeRe+tdTH2
WeYCnGQCZfBe7QI3Mc3Sg0XPKsEQ3SuuAVydqXHYND+xp3/OjwLNLfgfLS5BcOol
szprN7dc/LojZ+h2F1vjOAJXxyMh0J/Qq/SkdRZhqiIs4+4PX7LhJ2AK1J8ezWC7
6fED1dXCYiH/6Ai6ptaBxywkiwD0oAaFZXG5IisaEZnX9dcFFmQqSYBEgv0spj6R
Lxprtej39zpVdhc3Nsx0pKF5uVjdo6mow/pvSUVNlbmdZab0Bv5vWeewFBzI9NCe
23lh0WMlIAt19Y9hy7UCi3Ky2FX9Sp7hHPvxdklRQmlSL/6FplKzY1cbhIryzQjk
z79DHu1860edXxW0g/TxnULFul7DJvqjqGFL9Iiq8AH6TVa+A5a05Fe+aRGrqDxi
o4CHXjLI4Wx8sE2va+yYpwijQdmTcWSUWfrjsWnxvU7ooddIb7PE6jvC0yigZpdz
+IWUF2FOtAQZw8Nccs73DVau5rMBZbdU8K8fy1oKs9RsppskUWQH8LvX9zTqBFvb
itssCUCYR9bFgPA0l0UK+eYhxzmuani5Q/VmxRf5nmdAqToTmlDeU/1pJx8nQE4l
BTfjIXBR4EWVPG/rI3ArIbBED3MZO2dJocXAJl+FxlIhra0NAsdu8myEgp3Tlhj5
9CpM1zJbbQXGc6V7DMllHgttgvKGU7KNyJv9noGN31LkF9+/Zq4XR2sL1iCtpD15
gRoRJvQyeSfqsegG1vXu/Y875mGli3iBEq2lWFfwVUdhS4FXX5RbTS5H/vXxS/Ch
PBHl6xDA7sMZFKTPOIdUUsUyr0Qma9JAhPx6LLhlUuOD/w5GW2Kjl77RMAj9ePhf
CyZZg12IqBRElMeGRjUY2RFt6Z4so4f9L+E5LhvaKoh5u1D0WPvhml9t5ghfEbMx
S6VMA+dwp46cJb3as5gIidJFpejfYcLo1dJlS29M3G3fVBM67YUAxAvL/35Wybj1
i5IdXUA6bugoEizLpKK535EbBk7Bt8qeq2cYZYiD+cfqO/YXZ8pRSDoBYGXX0fhg
vU6nYgFLiMNd6FHxdkrQWg1bkJpzuC8CF3ST2NTOQxD8q7LDiN3RwEs0GWljqiLF
ulGI60bppDa3+4v1PMe5NALrSl+oaRq8JVGVKP3r5HlSCxXvfBBX2Igvxi4nut/7
KDGuJlxryXq+cwWVsbvgrXPVx7uWYnHVbIoTxLQQuMVqRsWWRHJFNZzoDxdQOA5q
5eFpEHAbsknfvOV03FiInBhpcAYsoUbJjKJPchjnzXxx4HtrvKlfnuJodTKTtzs2
jf0AOXyR33Wc8PpULj47V1OSomncvatEHSFE1z8TVcCSxMzp21QhrThhQSrZ/qPS
xjkQg/ddj3YUkIYRFpzDStL2937wlqgVerTbO3b3q+JQVrYQFACGFQlbqRqWT4UF
X2Op2X/AVrfqWSE9NpNr4s85NjrlpkMrEgw2gtt/4zAqlsFA4aAf7jqgOycJLEua
feRvZLQNfxnnOcwfjlAfO9zsER+6RJ1Lf+tbgav0AhSaUcTUOk65kbrYASYaKdAN
Ww33YtFRW24SLgNdZxE5GlY5Mpqi2E61HtzURKDhYedHQL4phF6CMlS78o1w3Jqv
fpj8nLM4cOyUFwJgpxhXSPZpmRBUlzaqOsZ9FCyxqU62gSbcxY3FdtGgUCgJJDIs
WsilEqQesDYXjE125aN1zu8O96etINGws4E/ykb9YVBMZHVZxcf/KYPgjJkaqfi7
NWtbUwxaD4GN2dB42jSaMkZGOHpFooI1zZU9c0u6K1GRFupOxvLdDmJD+ZMHPgbG
ULpRCFTiEYOxW7wnQ6jcQlaROLlOQx1942MzfA305V9C/a4PQGxoyGCOr178ghj+
OdPt5+N9cAlzSnx9Od8A3M0pcP0jZ8PMxe/662YNjHGHHIS2STNe2jNnaBdu7kHz
vAE+Ztsl3mhu0BuAR650ZNGFFossm5XHDg2kTwUtoH5P4VE6HSHXd+drmODCDYIO
AOGtk/SawyuRbvV22pZ3gZHLwnjvZwh4OwZVWHZwepnkgzstI/+Rd33I2LH/xcqM
qmG2Er0dqiA7KEF8mWlNuRZ4Tm80rDT0WTXuCn3YzV3X9HwGPko2TlJ7G1xbkWWi
Zk7T2Vngs+BkaZ5/VsT7hON8MriuQJDQ31RbgPzGxZLzaelj2F9wy70AwQdVQcjB
HzpgO4nUVLaHy6BXbbBdQYS7WnXQIwClZ2WlwyrFP8r0Z5voR88drylQCdBN7Uqn
bteuk9mZHe/eJa6AEROuNnvHQJ0oxr7ONep+e/6IfS+5h2KT1obk44gPyb3uOK95
gomL386J6qEX/j2Gceek3q8CRdiO7A+sxUysH6QwhRKfDrOxVqbrfzEyJA95KNag
/TtzJKwevn6FRCVo3SUpaycuxRObr2BO28yy11CgzlxuT2+fRlSUTSl2MdszGuYO
5Z36YSODoTwbqsaZqD+OeIp0NMgSK5oU8AZVJYtO/vD3O5GN7yh/lLUuxwenSYR2
t4j3Ldlixei243RmYc+6aiYhPQO0w/Cn/tjwnDY2o5PX+B34ClouBMG9emZV71F0
z1cOntfRL2Qar8AzIGxBqCZScRT4n/k2raXAkllz/6jkf6RmOd/UBFtXbslgNCBg
yKMG9/QodE+N8OmwBBCgGglrrb7UqiZJ042QmL4aH8AmhnX6wYNq1V6aqArtx2xZ
dcXbnCRSJ1Suf+tFZ+Gl6ohSxN9MIj3JmlbLgMOUbJjm6/UnCE+gE9IsbdXn6vM+
lkXzFNVQ/nPLpiIWs9dSEtdxt5S5XahRwjYCtPI/w1Z/XICTjLF77n/oXdRXaZh8
j+ujh0ucl8twoj7Tp9AA7CZQjMttBQd3pxsaDcWZAi+ryTGuzaafiWDoXgX/Absa
0BrSPjeXHuH78vZTVIHEYUS4v7JIq+K4AaI844kxRl9QlfEXRpHASlhO8x1IBG34
88+SyEvyzGCvXehXKsHO2TQa7jMleUyOtNyc3ncwlJShL4dMTdhjaxDHQMKvkou/
z/BD3Q4wnGDI0eSKirT18UKipSq/Zx8mjU5Dutfq8xZRT9yW+RvTBPvCQIa006CD
ni8kSYowCuODZD4yoqKh/zuXFmiV4PvjgqT9fXefwXG5XcAGyN3cMguuq078FzVz
npusyFoC72F8QugnEfTI2Ed2BFzPpR5PI6R/BFLvtTSN7SEcWcTSMyw7bwhqUz0O
UZlmk/S8GUSHro82P8YktYkgTNeTzETVcW3VAYjl+sVowzWMLzeI/5jf5Y+Yd7H8
hU0HIrr3+9mYtmamKWS2BB0QGH1jWM4TuSRkiW7VLgo7CxwwQgsiDvYahzjleVN8
b9nWdluHJ8Yd7TX/d9/7u1cDsG4eMhX+cZEXE1kyM5I7IQHEHggM/950NRJvgX0X
0YrkDKn6JZb/rK+RJUQEmhUinbhPwVQVq85L2kSyLTubZz9jELAssOM6x68rC/8v
EknUNl51YuVvxYdW3/HvPOD+DaDs19U1oWm1L82JZoQDaqrkqQbZoXg+e6k74EKA
cf2LAhtliJ1YnNueJByT+fP2ShhSRujJKFP7m0Xx5nYYGV7qkfgnb27tIWK1XGe9
q7ByohR+IuRkA1BOq143Y/X8UQU0KW52bfuWlrae7aw/jCKasyuavd6PlhxTo8cm
Wb/zYlhNoj2t3+STEKTiVjlqiq9sA2u6YXI8rBGsVDLalSdITu5Qo7Z0c6C2XY3K
RkiuLLdghSCqL41UcKqsqliMsAcHQV32JZ5008e3yDQLxf6qCNWCIT35Apu1Y9PI
JcHeg/ODdFmyMHF8mK3fEZ+B+aF+fjQSSjkkrAgm39w5AlU1dIUxvLDLor8vEgIe
7iFq+PU7Gb49ElwrIQ1RtdBq1X2qjlJm8ruvFxEeGllqaMDtohv5jb7Urv/fGvr4
9KwkXu4FaHNpj9TW9VEOMRkqDI83J6GTIoYCqmZ90LWGS6S9FmkKCPDbvpbSN3NI
C0ep1T+hQATVDdpDWVvIzt+23zaPJFSb21hbE8r80LsisQDuiwnZ+Ogomi2ei41k
6tqMHI/QuZYO6Rs6pknnANElJgd45JHUyVys4FuI0UZ+xiGR2fxNuTN7aaRUeEiY
0ebjWT/e6PAtC7mikGrYf3xsrUivAb47CQc5WXoc5A5fQjHPIO7L3jZdiKhpJx/c
C/XenXBHFcaJWMIV+ejz5uQtuNgDWyZ83Lc56p7EWbN8XDgixH5taVquI46smCkg
f21DaGzcI4kU+xKqQji9ZyplhbuwqlekRQRIHsMg+dnVnSw4Bhl1n6CtWm/k0gCj
nIjewvygZquxLCrs7micBxEmB2ONS9Ke6qFTqueDHV9xjT4Hdp/3wF7RlEIT34Jk
K9j+Bl8JtNlJdsjAHgByulDwNpYHq7TEoKNm+5qgeSqd07hlAJy5rWuorLav/mwD
MPpK9wWiIqXAr0GHyrIB9Skl69UrCpeTv0oJKw9QO5kytkbMn9z/J7bs0bP9fHWx
+jWYWhoxzul5W/UCJJSMk0LAIniLPmbekZZDD/ejKWakQPY8O6eRCA3eUAZ2CvWz
/s1NcAoahKBHO3ypWWCCx0NI8+87frnHgeVvwFAVlq496Jmu8bETal6YRG+6vR1/
irTB9Fop9DFAEYkb5Xs7aaZ7lY6EAzHd08A4er9BcNdY7GHLI7H7DtY8ZmTsfJl8
8ZnQap10y+WBVPhO+l2lsgcMavQeYYBbKsCflW5ClAhRTJitbxm6eA3CktuaJ4xh
r9k1NgoJn3KwGkYSISuuXwFIGQqYWLm/jAZskodNGsFLEUnRH0CVbKhN35uqcy8j
rSkKyVZlckwXgq70k9rc2aEO8+WFRLYarQTfBZ1im9dNUGhN+FAqAcdtdmUccto3
KeOYrKcI+oskKp7sHPDv8+ZEWSHvMsMyuLNxmCh4uM3DC8ST60anLJph8w6seWTa
LgVjeHVUmMFMdArC6w7Pedur7eTHaCMdwnRlYD2BdooCsbpAXui6zYd1oP7WEJ7G
9uDruqnVhI3J4Qt0fYGI29BLrJwPn/oFzNo4K8oIqNHbbFBBfGzwuu3382kCInp4
tnd1mLPmpUa/s/feX0PCfXcANNWSykkRMWQlvSyCYAFSzyXoQYq+jf43BtvouSX6
KsS7iMhQVMEagFEM9XLuWPKUIcattIh9zNLiTWoyNaa81JhFwcFitzPHmgPxs8Rh
/6q3MKYP9iCa3dsDRS+ydU22dlEjRTH45mamarTOOKQfDTujJcTR/gjQq9pj1nBv
LvzTDbmbIw/qOoRwGG08HjU0xDcNDwU8lGmGA1keDqnIe1YyCvgItac/pX/9XFH8
h5yrnnWiFN5Gvk6H/rxmSTdCFtgKzQQ/BhAYaFckxWwcM0F5vC20Aq2F4CNEJgzz
iiqcZyBzYskOlpokZbEHZXFRyBdBgZWv4VWWaYC2ipzqhbJ55jcEGXOEJ0gExIcr
48W1YwTkontu8jJgmD7foJ7O/RdUOjGiqmWhvXtYkvuf5moIuLnHE0WiIj6DhEai
5uLyG9ZfuAnm0QTjatjxuqLE8Xr7kLvthiLQZSqdalrOExgD1Qui57A17edkNgF6
oRhJqlZp5fNsWhUbZuuNb4EliN9H7tJVABocXXVu7QwPhEp9v1KzDyPdPcM4z7L+
tlXOfTyrmKd7qkwU3UpbJ+Fp2YQFB12OEnORZs91J3INCR337CVqY6QDRIjxSR0U
xMGtWqOtdwmTQpJHKkkPcYfWG56shJ69RM9E+s1DAj10W++BgRgysAYV/VDurIi7
TP0N8p9cR2tr30h/wV7+IA6wuXXToSd5/OzHx7iWUzilfn0J64dO/b2QfbX0T21P
fCztrBZBT6l2oBz36zwFArssswAdF8L12I9jt6/VSfsxpquRHY35bczrAnUppADc
8i/8v+hEbEcGRnNJCFq2o4A1R/tbLnmQQvfGThbKDcDZ1zoWhnsoQOa18WxJ0WOJ
/CEtndBDL8RkJRJ19RPNFxnZMjHLEGl87ziRiN62UNSp1TL/nzL+/jV4iVcMNYSp
OuO7Ye7h9AlAzhAM8FRTA6X0VugbOw9qndFIuTtTng8igmzwiw2oxdbwNpHaMDWu
4rwubwOWsL/pbkzzrGQjTal9YSX8cS2QR+N+5Di5VVZsxyqpm6m2pUhxB5bscnTL
yCHyQysM2wnoLbie9RiAs0z1bShzgd7Rua8UOTWhRMNZTOLyDIg1Ti4Q/niQAc6Z
9UL71SzBVRT2wlEOhbcqRMFFbtpHvFgcwgeAAqssHOjoYykW+bkOcbVTNsAkT2Lc
4nUvTdFp1IoYS7OSUMVZzqCJR8FxnQ8ERgg1YZzv9Wsg6pFqluL3ps5xa72P0aQE
VWP2aqJhHnoP/LSb+xaQIJnBcwFzcFLoMgTXeb9ZlH1x1nS7VyXE0IHNEvtEdcZU
7dVazBz7oZBcq75PzbWhz+2fz5+st3JQfHnjGZw5VZJSmtO22iQEDjGZS5huKBs1
/NrR4E++HAduINWp5JIKT/rlRCDH8qQhjhplUQlKN9F3eOn9K60zT2sLL+jlROrS
ZXCb0ncoYZXd7ARPJvREi3ZztSyA56zbQqpcAYNxzSbw55R81sA3Kaasz/Jp5Jvg
Eja6ifuWfEI9EYAjfawjOXexd1LYnffpVztNI3ZNDKnLF1NEkIK1FDCak98bA5/s
ExIdrBgwE+Xq/aeDTW7PcA9QFhEUeq4DBDlu4Ei/JJKJBKC1SZ6K4hdp+Noda3bs
mECcxwKcMTj4d8zWXt2/rYf4XzKrcoP5Jkv+nGpmELJxcUhFKb46NExiIsTD9OYy
p6bxufVmAL0LKrpRsPTd4/CtlJI6VNY02sQz1i+c0UZIObVxB6kMpevFOUh7vZr/
R6DLl1JPjcLnn4RaOM7UPt0kS6Hf/Q1Xq110aPnIXj00EidhONUajQzDueieLNRj
l6Mugh8pB7Kj1RXW39f8jT9JyzV1kgqheTFfbCCIvkf/dAO4t1HGqzU2uBoozyl3
P3JLhzYy33X7lxly/LEIm/xzToXB7mhzyYgpLb4BU8fypkgAhx+Y83oP68fpTcLt
SUCCLUk1NuR+i2rnjcP6T0CdY17X/UnxnfXcBwmwhyrNRCZ2iMNqbD7VVgVw41wH
uYfB8gw5uqPEml5R7SE75NMfSz5kYvHrmfgaowkEAFir1GrXy0Tsnzrbb4Ib0BPV
NddIxYLY+lNx1k3QKNvEEvULW0oYu2zzqYPx/4rckOa4Tc0GB84WhGP8IzXhf8lp
v5guRv1mcqzhv3uJEpSsFCSwX01t76f2xsdDTBz7oSY9+oTF1qcEr+nINnygV4Yq
FxiuEypJNYOzdkITl6T1s2VaHEavfsdt4tyyohI5TCpOdFyXfat92CxYW8zQ/3cs
5nseYGZSx2Q6dL+RnyPTpjK6MZulEDcA6FQH/4nxS1MeAgA3B81UyHzV2B622zs/
P8Zz2x9qucA+sm5un00SHlc0Wgot5PFXwyIwo8C1AKoh5Txs/ROqURmol5gDTiXN
Hn0JzMiQWmz8IGDPFsHemfVNtLBwF9kbqcKyjPs+MF9+GWc+LdiyUDDMw/1Cxbpp
k8BejvozU0Ji+v8XmQYfLw7mh+x2zEWdW6OKDhf5c9Z/T+jjnpt53jlbf+FR6+Ay
wMqUvYrMQHt0qWRqHD8Y7UbM5oaghMi3WwC/twHdPn1/+4EECtP7/9tSb8c5qpG4
b9+UJ2yyGumCQWVqEBj6d/kfbMkgUEJBzc2l/6/I1QuL9nrpnMfchMU4b0ShiDr7
JSaAcS18i/sZ7SdEppTJPtoxcJXBPsJbqVa4H6x7+WqdAAyOuUNy+SrrSe9rFb4M
7GLjJfjbmhJ5KEsvq35wQvjBD7ycHkKfeNDjHHtGS/lYmySLefXO4/FVOrArXdLF
xBN4SYTgR+AP0iYS9+vH/Vi/iO2pZbIxcDZJiR7P7JqZOKmyyHasq8yDHXljKnGl
RZOxUJTTI2zE0MSCDKaap3f+2Cn1PLDDTAcgIOA5p9ByejfJuWgW3AyeyPxv6cAK
Ippj8+DHS1EWQbuhcffJ1SV9gPnJaZ566ZiGYRN7dlYcyvf49sDbpbfGbOrpX5Tl
/+ogTXpKa0koquI21D/FXQXuyIfXWM5UhN/C7PzdnkZfthJHvvu/1AwlREbO3Nkp
Q08w9d9Y1mPTEKIJD5jOYgXmG2tjdfJ7HGUW++eL7HYZvOurGYkkTB3VwptjNigk
HsEOK0m1QICv/7EKJJLrWypnPIIfRftn1vKh4tA4zmhwLa6zmlpnfXQ5qcaHAxhT
2ioztrh1vxWmGr7v6VBJ6ZR3D4ou2ZLbsFAhWx6yji4akSGP2ka6pa6Ost/lK6op
XUwN5F9/pUzNpw4JXQLmCrTyF/dEotCHe0Dr7aZ2NjaZswUpn0UDPtiNTfoEXwcP
RvKJccy7v/WobaRfNerrADQztmTp7121jGEhKptVWYlQKvO1apyt9l1TTOTTr0oj
8kZEExKYuL+g0xgzZTqw1NMkAt6FAMgMVP1GJwbY1/6wYyOc2dA/QqctqPWSSZhy
F9EYo8xAWjrsr21DzeHRSJf3R+Mytz5C3c22TJDuYddQh11gWoa2BKh3aIrRgxJ6
n6xGdXTO5M0P0/shvPYtAwcMr0rzJt5VZYr7aSGv6OeZ6gRUxIO72KJopcpvj/N4
hng4ifSPqXXdVzza7lwJWffHR6OMT4C+Em0hSg7vqkTDx1FO9c2krkw8SAwZ4FHN
M/txRaJw2sJXrjEXCPCCHd7IV7E2gpXCQ4qg079wbPWEGux0jdh0oM0SlAC8MY2+
q4izJ3epgh7t7jtgybX75v/M61jB2wFUrCF/rh5esJ3H2VCSdLuv9Zv7rj3bSpHK
lyEEP4e0P3lMk2YZF9Af6r/mnoueNM1/OkswFpd6XdU8mau7Dcn76zJ5O//phgAX
yDzmqqjMm0RVlbqsf7XHHparDP3nQePHxvsEn6ynwcMe9bb8eyRASqPTZXEI+xlB
/8sbYYrn3zHiDm2HLYQXCWCA7FufnemQtWlFUpOJbmhsZswoNhyy4qfIraWqvJWM
wh42MdFqkHJ88W2e78gSdlttNb5VljwY3BvAdMZX2gmPdayxSFWjQzit07XAePrA
UbD0BUzGD1IXvZKBNVlhooyUuEG8ylb3QPiUPBt0Osvq6VYveI7KWVVoGtcIa5bN
Tz1kllXXlvHNiAbgQ8eONLWI1FYqmcEUNoOP3Ybyz/ceH80JFzJoNPZMvfp9RmJd
4Dk7S0EB8zJC8NR9/r/VSWpYe4st4XLOdJKHbgm1BHmCrnlUlmYA4yOuEoB2LG0D
RQNbVuO1scS6r8eQxrgK9uLDLxXHOBm1HGCHZX23nPNxHXFKVF0CZKp0SUCAuvna
qwb1i+2Pc3tazhIjQR/Z890IVD3AMWrUwaVQ+ZdLRQi3RvPRXnXZZI67EoIlqQfK
4pI7SccQ9snJTItDSY5et342+tlOsTlk/odM5rA0cwm/m+L6veKiAND7L69qK1tJ
5UkgyEdsbEmNjAkDoHzGgSlpHXFlwpp9d8FGZV1Glh81pH2xM00LqnxB2tlouq8T
0OEuA1TCR+bgUdOmRsWA/sSDCvWuxNS7YW3gJURJ526NUl1g6CEyGe4waaADRn6c
ScBKDzsE+NF0AQ0+kiCbKykyjBYLpewTAcnkTwBIHEjUUTEk1mZcnyZGmc6rnIhe
xjkDNNE+rT4T2BVDNsNlYiQqZZ9oFHI9DzjEjC3eQq6bg+NZPtNnttCFt6NQQE+4
ip3pHI5myeQkQQFw9MXyeqo/on6hcC2PUOG9ceY32LSMVRMPVDtFGOLXO5INd8kW
tfF6K2FNQowH36DgfTDBIX5A0vrL3TvbMdFXjlKnv108VZJrKF744qrofJgvJb28
hooOCazaDWNDnEaV/lgwltU88Fcwcxy6o8s20DLKi/zOMxLtK2fWZARNVFsN6IvT
3ChnaSJMDHIdMArG776u43XlUrJxAESU4yASXz1QIDpzIsxDFdB86nTpLT6VOGD9
yPWZ6jq8P20IVDs5nu3stqoXRvU5RqP+2SjO4mqiiG0RUimEzzUhG5ZwVUROAlvu
1Ks2CNhQ4K6+5vLwOOLoanTCovY6ADU6CMMh2+6zn13QDjsIhqeTU8G28JTJmr73
F4Y0rv3yEYguSLU8xTkf8tkBmbpV5UTP+BgQY+Tg9xA2PqtWjyS7R8+9EWVlm9eI
il8pZUXLrmCQHD03Wu94+1OcVPrkKyYh9pdfBBbGrKEKhLFP/1eWDEesSr+5t5TZ
WzLGXdCHqZYzj2EY0UNRihzBXe/cYzqQyVcgFYCHdml1Ea7rxPkXnqw2EHpOl58M
MXKyGIjiI7AJEEDQi0zKhi97FsS4nr4AIW0fwKwOA/rDaGO9Y2q0EZJ4nPoGgn0c
He+vEZSL+qMvbnsW/M3M9GBGmu4NbybzoQK4MMRgcbViYMsy7kHFSLuDu875pxfr
7vgaChobhhP/7HKMxg436kmW7CXubnw7m2GcTtRQ5poLsU+rsXwSMTNU++IBv4vj
7+hucrhlK3X1VE+1RCfsILp7JwZAA52aYIVO8P8MKmvWnabCbVYrBnhgI/gLM3Oq
J/BklTJsGy8j4UCeZfk/7K2NNuWbpz2pc9Z5pLl8KGMJx6uOyvvMadz+n4Ohv836
XT/8yp9r/vW652IQHp22xO59SodLjBvKg8lbOJYZr4rT7oBn7Io19XUxoyK4+l6i
ndHtLIOOHVpAmdx0M+1FA9cnusVT4ZXUjTu6chBpvdvxR+ZeO3gUSgcmkyFHzMJt
qbh7DEUUob04XQ/b2Cyy0kAjWITfFjyWyIZU9E0m5XjX+rkyeObLSYUsl9rdCdsG
zxRKY3W5OeZ4SKLVQJg66bLuf3qtSS/0LCWhKRHCe/2f4G/kY92NaE1JygxCHERw
nw2ELd2oDEqYnvPc5lF5zVAv4MLXN8YQRNTu/T+sT3Er3LJZ3EenLB1Z1rJTWe7r
es8Iquvrp0PV0zZOtGV9oJ7W1fvmT+BlUxZ/7/5P9IjDS0kRepdOmZLDEmnSGJMs
YI6N7TqciwwL8zMk2D1odmBO0hVFxnBZZClWpkTjMaOliap/PbdCpBoO9dY4kYGw
hOoVa0+GplRsmVorr5TNu0uSM88Q23ei2nAw95od1zEgc82IwV2qjSa8JNYgPugv
FHL/9dwWKqGMAt3+/OEcatBNfK6Bc7JCL/9gIvdmUvPh6nHkD63EQK7e64Jq1juv
wp4VSLRCIIhY5/X2bx7crmyOevZO9ZGE3wVWhPPX+fN60WkNJ9h1stmVnefDD5dk
jhMKrQUX2wnE4/vTOFyz44YVqQTq3PBX8fosbjum3Xb+fjPsAFiTMEqFrthKpeJC
chCZ8SwbGUfbjSsKYD/IUyTLBcezumHvN4MevKUaegEH936CMc7ZhKOABZ2oS2aT
lgYq/ZXcs0iLfAl4yWl6I1/WDrMc5jE75qrOcBKZpNQ+KCpzHVv5eS1B0wPElhU+
KMY2aHyr5zsXQIVpi7BLNZBW3SdYx+rnlk02/UueVLrSQfeCpaZAg7fUHQK/ex3I
07DlZU/k4dkIEs7lxN7eZTDFLBX0J3MgGqaBSMXGBPktpLASxwiY4gOMcYEJ9IWD
W7k4FOTVwUNNgthxZ0cntzb7u6a3TxBwHIJZ21tMQLOBO9eR8xAbzZhTo+qkPHyR
+KTFr6TL0Lugs9nFGv4p2QpJNBT5ADExQXh6CFSy19lcM2t9BKgpKPYB8yW+/R2b
fi34pIeQPQeFwdQnXHbAgsql+WvyIyXUlV9by1Nt0o8+thgm2uxq+Jps0BbNGtCy
I7rahg0E5YqNqAdCcCEjUlbDJlhFj8b4D4SiKOtcmbSuvwMX66cPr5f6rFNyN1z5
4KMRKHFfiv3BFTJid12EPairRuyX1K+14PC6itxD7tJ6IchRWfzd8OhtxVj13ENB
UOEyM1oEC3nVaP7MzYAwQ5lCn8y009VSc+uSCYNOG23UlCqHCzh4kZTaQmO+tOsC
vqi/mHiIbcYQjOYJ02LGZICS3+ZfgzleiOH50EraUu9uiQrQ82suIe0yidkvYAry
SAPt/NlUEHOOCehIbJFfx7rdwrCifcH3+nwjO43Xd32iZyJQEYbTo5BX9ulGmSqp
MBvJhUf2jx7ayiW8dS/SnjOa/CmPabSrTaiAM2RAUBCZ4mgFVjuLZnNVpG2XAUNm
wgvFLhpPoA2fUp5fB+J31j3L3EzSG1IDPCrpYOQEOTpyvQbYVvnE5ygvVhzcxGkH
65xWXvYPR6RE8ti4udRU8KYe2na0qNQafUPaAGASpWm6mIasQyVZb2J55xCAo0dm
gdm6hTfGpF7Sn1qLqV2ouBDXt58/zokn0bKd1rtBYARNtHZD/zXZsN2nEzYEUrpZ
ubV7BRVyNd3rW9rs4xFFTLEglHkmNovWjpMQhIu5ykDoKKJ/O6O20YvzMxoUEHkJ
0QhcQt3drjrIwqcwjymvUKL8WO6IkLO4B63aVSi948INs8vkxXISknLfPfs4wQ2l
m0wCvcfNGqJ8vV7qVnDkrAxXPvzmh6aTQ/FKaM7iJmm8JyZxy5ElS17/0NA0rlne
/j7Qmjc32URmAQqrw+SLLrZzvY4MEpwBEzxg3uZoSbbmC8cZSBsptO1gjXwIYX9o
7zHCsfoGze7MSkSGrdscDNjr4mvKsd2o9QLbxv+Q4w+luW4G5WNy/H6xuyTBD9C0
45WEIfSylKdk4FU10MO4ssWHDCb0AvDanccnnnRcosfphwI1jzR4i85igAxFODkQ
islyCBM3B5zh6VRI9/8P1fm2Rz2qFyp7OhMFIfLgG0f1cXCFmLDNQjNEGw32P0Ki
1MOxnLzXfrQPu04C9Q5VicQYeJ4NpjUXavsaMTQ4vww33GkmAWjukG6r7vP/Nzk5
hROXy4nR9QOsPQZ+UqtBWyzrMKeOomTPhYW5c8ARXF2zMvW73jbvswhuRBG70+we
DML9gJWlIQnMXY6GbZp4q6/bPdeRZR6+aF0DrtHSn3guyia3j9WxDJSP7EL9GJqF
QszldRKk/GTU+ZQ68jkRNr1VG74x0c+HJTNctFszaZYsZ8diuyrBgWN46+jCNcn2
KdyRy8bHU9GjYVHrdtpPRVmpZSfNwSZ5TcbtCBpAa6kIEgPynazFXtAoE/a0feVL
ODGfwpPpGCxrNWpQaG7WJQMMMv8OXASoK/yrZ1uA97Ntoj7cxJd7radv9f6VTKfg
0h6iQFJrWAcrcslrybE/bDq4IaPCr+YzSQqROlsV4iTYae8egPKhoUqmmmg1WkRY
9tCUKiMCeGyxbXPViDjHuKeLz4795G62zqDjFhy+sB5UhO5QCDqZ4v30EvFeCxyH
7NYetraY3qlwLWh3DkXg4j6SYxVpoXvYSZ3NvoMsOFeYv4HxkUOBt6R/fxwn0xXa
bzz0w/VoXhdnl0y6ESrBrBvOEt47zGt7dzAEKx9VcmVxfj1bH1Qk/0U7Hic2jw5N
9uYf0+aG+43qrlzdp6sY6qxeTJg0RT+cyNbcJskovZtc6ABEN/vwA+dYe3EQ3FIT
Sax9D96AwK9NasmX0yqzP9mRDcySgp0rjaS/UfXGWcNFc/aE/acB94h9wC/oI06L
agbRCrxqcFnHxzC1/xOZfjJYhvwkQbjpB3iUPj4s56xTZPGEWnJTZGqU2qCRRfDu
ZgZkNGJYXtwrcUwxfQo72i09xpwGWEExTaZ5z5jBiDZt0D8Hjd42P2K4qn6Pi4DQ
Isb6xtt0wi7a+BeNYlZRc1XEY6LJwOQtRvHZ2Tty+NcjyQDiUcTXeYbmK0FRXaJK
PytJPHxLl6OhAlSRxI4uyxQgiKvPUPDwzfEDIbT41p/vhXCocgYtUwPJV1IKLs/W
PWaSsfATd4Zw21ReNorWZidXs6AsjqQbs9xF8C1T4gkd5VPCnzNOz2siGZfJvyVU
8QR7EskVKPpE1ceBSoqElwShX0kklmzKqOGDddkc0mjHDhwn9mXTAKoYDIZ3uOzM
bDmJec6aBQLbCDZjddGRHMjZBxYBS6unhK0Bc/yKBdVvTPA6JF+bd4Alm7kt2Jye
EK56vktma+mSNJJ5e0myGKj5uqJYTDB+kTOAs7av9VN/G/YtFtRtoaB2KGTaTccY
qVlN2zYwQgzdlXjJot0RCR2PC2UQAwH+61SakttcUfVadSvP94PZVl1yNxw/eMUM
Ijlqhnj1ABMQv5hDnKgharebdf6SZ2JIdEtDqIX+yu1rY8MMkyuH9HtqneNLORoW
pSogJ7qzkqxIUJBQOf0BXd3bNIG9sXYmyr5lM3LKYxroQrM34SiKti0ekFFLxbK8
QkpCs93lHCTjnwPF3LkLi9oRoxhzvZSQZv0uwy4njJRDnuVl+lO+whC3imH10aGw
xFc30C5aRyh8Pp8p3004BEKzs53VCwL39Y816SuIkg9EvfnoFmCytzD+qV+mqJHw
X30GHdffamaVZ7de2Ws1CWSmXNuzJ9PZlBMK1q6aLLGc+ctwb5YSNckcnddtTLCB
nXC5R/lYpJ/bRYkPgYFX6CXB4UUZbWXi/TFW7kd9BBVqbt53CwEmqbqekPOHXrFU
9qqmI0R13nURB+bm4UqsZTIlz3KQNaCrUP21EC98JRhVSQUrtBPOSnM8CNOtzngZ
LcPQ7O1WucTqNY9LM3TG5mVf0b9LfafkOoQcCU+L0ugWW4Brj1xvykxCCp7ev3dH
1ZJ9VCtC9XcSJw69oO96FFKsekTQ6SHvyUMA0meaH2k6hUVxRUQCbS62g59P6Qpp
oJf15SeywgCEwgY2S46TFXekRpsEvL4nD0hVppUunK8UsBLNbw5VtIX5RIB0JcDZ
n9rOaCJpS98Y+g+Y8VCrQhFwv6jsjvyX7NRXWv5kQhHNwSEkRX3AnbsewlP0/32X
cYFMMTjP7p8cImS3PD+bqTfolqASpkB2Dgf4Yq1X78tkMUpM/D/E8x/Oh7WEZAMm
NeUUmKYfufLnkX9KzB5y1VfAQvBcGxcEiknTY95ukBdIWZ34upEOYfOZaGEAOYNN
f13zlA7MIasqYF7ObVZ5+WNwjWPdDKWClfvB9CWWpwzX6mXGuPejO9RhUwMkmY8a
haTZ1CJoC4DEJPDNxw2P7KBYS0RZGDMTJupxzMKTxPJJJOhEgUErZCJTTF7rZW5k
LSEkwPKY7nNAND/vNTskg+rL+XPu+g4mJ4oawqtRa92C1QRr5gnSzDtqHelrGvAY
6xapSorAjtfnJ47oeuMmIZP5SGNgs5JPYlqNY2dfJCc6CMJDHRMO45Jsn50cP1jN
pREUpj4Da/vgU6jabX8bqPtCGFgAyxEzWy+t60dlHeE7L/r7USXUA7Zj+p5KMFDG
cQqR+NTzVz9KSCd4lakq07Hmf1WqFCQ8o3L/e+3olptbwK4NNy4TA3hyUoVW7Zt2
pCkAi7Kfxhvdrlb8n1TFIFLqCcfYhM8yrHXK+EafVxewbnyDg3mczJKhf68Nb42G
Iojqiz3aZvj3lWSvNDdLGxEX/XRv9LjQ+jre2IaCte+9DaZiWwfHASLA/01lAFPa
pqoduzoTCT35xuGOxmX3TRgtuL4ykR3ATcMax9W83rgwvQPbIYz95SzErLqepxUy
rstiw/FLUXexL5I7ypsTk94dz1CWBPaX6iVJMQAV1MJFpp6e009W/7fyI9dss+OY
s6U/ExtmN0NV3cLpkdZ3DgBhAsEMKNvyDUIq1dXOV+xxvcFi/NOG6ilcY7fCcVIA
RAzxajvlY0TJHWlFlGNN6ovwPkTrwu4WJaDr+rUetXEQH5PB/s1yXdnBcgtWMdUk
0W0kBiCrTP0QiZZXPKafUE0HB4IMKrlJpNmtAKZC1ECY6DvUiE8xAzkOkLI+m+EJ
y8tJfVn1Ty8JKcSjWmkib6V9Eq4mcIvRxnqpCKCuuM/eQ3ubc6B8yyPCQdX5a80g
G72YnUlFA0u2vXxXsV5Hxi8+8sHPkmrRd+Bzzqmvx5BEdVeWLRa71FoL5I6b6FJc
EaOhnp0tVi8zjSTaA28+NS6i1iTe2GxpN46RyGKZdrp2n2n134fiNvQ/h0cvajz9
6bYrk8jWoIYP0iTgNovlF7nlasqhSiGib3U+1SmoHJkKJAEFJboKDm0oPYeiCIVC
PBd9JRVpWuGEBLAaGUhyzXEx7CGrsNnW9jquA2WQDC+JxK3Ne6gqtY/X6KAMc5NN
I74GuSXi8EXQX/39nmi/JbiGnsLcHl0BIgvqUT4Pkk7pMB7Fb78lGhZTGJv9u8u2
3321Vpdl2g7vnQsd0OXlp8tGDqlHT3ySFLTAGeob5kuRoIMVjQ2Ty1b+gAF1Th4Z
jppqBBnd3Hru4JTeUeq8/6CpcwXb/DECzMiQBbDnU1ii4g51Hw32ZPMTU0R6iCbK
OIy+wGlbHo4XWPvcbMOu5k9Q8hUEQtSsEUFP1XuGKDLD5XCiZWCMwwI3QxLBKmqR
4MWVcKqA3RnB+YdnzZYewCEEo3VqqtUS6qUR7JFTZds+FdTD5nhVNSFSiFnAhWtB
vt//CpBNQ52nJA7O7D71q9VdMawxtRAanFlG6CMi4I1H0Tk8Zzny1wkJCqPmHHNK
wur0WHH582dSAedkadtCM7mV++u9Kl+CDKfPgidjkuRnYoYuWN4jRrT6QluDcfHk
D6z5bl0Ok/ib02VprRa0w4dsDcuuIszdAsIH23Ev6DVrBVE0x0/RXtR+s+Kflocc
NCdU3r5c9gs1/TtS8JCQpGRobcVsyyNm/CoPGVPr/gWFDHMFPvrPrsNX83CVZrcR
yUhgWdvshyPh29MRe0g/2JZTwYfbvKQsf8UqINfhMXVxXyaVlffzuD3mn+KomybT
sTH8esMhhFYfVUAT8KqvX5IFDsGF/+J2wEn97BVu7+ddUiICg9DRzCHM1oyIcckI
uOr4G2tfsVsexXY5blnfnYSyznZ5q8brZnCCcffIFkep+IKA3uSUOKltAGqZgsrn
5cbU0PCV+YJtExjr08CnC9XjaQDtnLjg6MkkKzKONKgpJpYwXmDwwoPhdUYvTWJ9
5RQJOMH+ZyXgvnwm47JpSCLp20+VuIbPHz9qlXU+j2WyCHu514o5Zy5oIr3rCmNn
zlF0hUdP9jE/IRDZkAaKqybGT6AVBhHKSxK1KG4jk7sgq0hfeJsAFV1963IHHKYL
oe35lraMpFBDigAn1CvANBJzXxtn7duRgFi8hLcYBXx7TZ6WqmzYxWj48KWx3dHM
mCv3ISqdhe5y6xormwEZxqmFV2L14n4I20H5wgLhBlNU+D/TXnieIwmXB0QIUex9
7LHY32Uv8k/QUjc5YQzutp3vaMcDww4B4rdS7CCfRMLLuOTNCn+2XIO9asikF60b
a/nL9iS3RDHcHwFA5Pzpt0h/odFq8wCNeQUUXwWPpUJCzQZsmpGWwqMcdMRWZof7
CYwK0ie6pEaIiu5BZ8Jkm//BLayItt+ELT4Lv1VQeoKgayS2TFgfV87Kq5fs6Knl
YkNvF53kNyevIWkwJwGoNy4CWB3dnkWDMcdjJOH6gGm/FjskJAafu171IByeNTFS
ySpcItFyf8ZEDFM70IBPgWJE0SBGxNOEUtt+8Jx8jXV71I1ZdOIcv/cS+iFGLk/D
Nxxy6hJMtk7aUXLP5ih3Za2/edrFuVcbqtJCATvjxhorcWkzwCxx09cyhCrJ//fv
hUQHHZEfdl1py4gxLbPzEawOKGX8qVlbSoeGx5Rwm3BCOwCoG7rlHVfd1Bw+F//l
1SVedIwMYkZ+mQrlvywaXjizpbIPyVg9PJEPVopwlBmmezfr5CYP86BO7wmR1W0D
RJXWIXeW+f9CYYwxn0SdPdUHPspIyX9bLMxh0LToHb9fdrmhxyxBu+WHi/3yM9I5
mxuUTwsLkDjH/5XwkpRsXe6f5oaAD4q+qAJvl0LsS9YQCG8gXOY+nVyc9hiT7ZE/
4vAln0Aml0hvn3UA5A9+iCIaydomGLl/AWy2fH5fNnT7Ui8+j2MYFIS46EyaUTQy
qOi1agmDEIljQhIjG10pP4YqfRPs+msq5oDp41wDH7XNJSep30OesfCndx556beb
r/3oAPHULq1IsXAyHiEJQbgTwA3VRE3/Xxbkw3mga8A+nA3erHqjX5B9+xnAgO/0
k8TjFzoGPMcjnnl9hNVbey11T7kAbWQ1k9kcbqlTkwVfiXZMxHyqKnInnbm8hN4u
QaG8wfQOGecgfuCeQpFt93YET92zJiOQcfXdN5MPankvKyUJSM/FTdj3w9O6NA0U
JQVSnViGR5s6+uOOSb3897+CmAJ0q06yqouk/plk82zjxPRtJgyQ7UkXah9s9Yx5
DDbfbWVQUMn5GyGG1mPcDwh1Rzucr7659PC5UnB0AtA6gsfSjUrlm9MglR1D/uQo
3HtNyn7YQcb2NtDFok7mqpIAUXu6k1T3hfaCwvwbAenc/yfINDJL7xg9UTYp9H8O
lp1bAM55hj4NlTzgPLw9WK5ftgno6OnJPjHMxJ2CEpPrwtWke9I955opXZcplyad
kfCIhe6siGvoZRm+soGyS3MqUNcJG0iosHD27c2dM12ZG6S4AVfVTgpssMRzHBlm
XlgU46D6GXsYJCTZCjVJCOQe/0aiB1gCgHinfX97bKcLvqGoeQLWH+9UcNz3meTu
1dUMoiAdSEvUZLc1NkDVYpkS2KuS5A+umdF0OP1tZBc/PTaxLmobKkdQgWVJ0EfE
o3miMpQuyLJc1AdRc+3WY9Q/sLSdsr1WXhh+/h4ZmPVnG931AL5LLfyv7KXubB29
p2UMD79MSKt1VyetjJHYIvgtNHpvEKeRJFW1Vo7yZzpuBMEPWEusUrTU14c129OE
++s8bcoZERNSEXysUGh08IWtnzHAZFoqpCXHC369Mci4t6aFCwtss3ERsa8O2b16
8j4eaJuCA2l8mq5Wp8otlUTJ13Pj4H5c3PWEg4vu2qC6WZPlPT5SGNFOAQywVkmF
emPegvsxb1SrXpeI+G4IfcQo+OVBXlJdYZhZOuB+TFIdCMQ4nTSlGr09SveIDZcD
tinzxsTDUmMrYp4WDfAdOkEutxHWw4buZ1A2J5GbOee86WakVoeiYZOwBP5IQ+fS
Dihc+FsqtnORmSOvZ39IOaVJIqbgyuyr5ahH3QZMUpxeqqG64a/agCHUMzsa58gy
l/Lkx0ppO0jzOPrBBxMyeV+4mrXCnIUn3eniAN3zLGRQ7l6fCk3ZHlkAftVXxdvA
7Hujou4t0McfODttbhT7DGAjk08PCZFXdzHBL6EdWAVdOga2Bm+0GU2jLjKJESau
/9BAKchkhUDUV4Rc0/85HmChuVhRUzgM6oW6yI+ZV58VZuyNReUNyqSxus55yf0B
Bs+9N0MGMdRdGNHXlvfOlHeh/tk2tqLmFCDDIdapZ518qd3hXX3y/8HBPjYmpUHF
dt59zKRE3O3FJzmuCEqZHljuh/Tr6e6dThpEuYGmuxwkOC5Wg0j5Flr43uApgwhe
HNjbLJrFVznYfT3sJTk0mJLjjmslapSBfKCntU4ebfewG0SA6ajpJ4aPIvvkrYHS
cYrHpuM1miC5hiqfywG9h8SQXhV3Eiv5gx5w6czlohurgfSPOySoKiFNK6fN7v0C
+5CYVmI6lFiEaZG1rocQzoTDqqp0MDvkerdCYFKwkBDp8bLhXPzHEl2pRME9iInH
jqQFVLMuXQthd1fRrZ8rxyScJ9vPebhtxkkH1LQSDxggjNkusFe+fu6C/KgFCRFB
ysh2W0MacJTp67UQ2NGp+FGdF+tqaUyl6uV7ZKoyPI6izy1qBM0E46zQ9CiOdgf5
aHyXj9aawHLFxpuJzbU9lzye93hNoXtukAO6uUHb38wWQVEf+OqhWXIEdSzXRkn6
kDSK1UYXZyO94njzhO/1FC/5/jIGQeODlyZ8hTClw+VA4PaiTavt3qBcVodjq7cf
LjsX1cmb2KdRAi173iZWAIHNYOBeQf4E01V2L6mmQnYoc8J1pS4JrxXSzhTOhApl
1Np7dSGLMVNMkGL7IsfMIXvl2z7Vj9ryNPTWN8dEL1Tt0bJoRn8krlCOjpggIZXR
V21u1x5eIO920m690WmHx3mFGkAlwjQiEQMQrzdnaYgiEdfXXDGMFGXo5eF2VWB5
1WxFVqjFrMGeYVV1XAGhc2xK+ujSpIunIhFyBtqwV6FR5jtvcxJWPjHG0UiamduX
3aRrHHGK/YQmogsGrBm1ifCZRH4aypKxV0cQeAYYv/ejAhRfBTW8gEPruBRn1UlN
bR118hY5W6mYbBhHwjU03Em5jzUQ3lm6mJCf9A8qT4pPFS4wtfQnGEquuT5KbSj4
StfXXh5WL/3H/0nxl77s3ZuaG4vD6WOBF/Qx2eO3IO4qbZsv6io9fhlHyXmkEV9b
jGfsBp8QH/GKM4PMNKtx/aWLFOfTT+sxMJA5gp/NLILWf8pB3OdrQRS44SOoeQM0
orxs0JEqx3VWRVcXBtVY/aHqarl38MA5xyhV0+pKjynhKE9P1N18od+SHdv5Hff5
SeIjvrPMSUHkPDlEMqc5A+Cwsyx9LbYggisaWy5IUM+9QLt0ZrsH6/pseIguCODG
w1p0mCf0sX5CjAzwFiwNmAkJ7fyBdhAc1YEOM1BfU0gfdGLSPXL3x3tA67rucb0N
kVcIpNG8AQOL88hqe+V1kjX/COVg4BsM9egMI452iTsOV5eAIZxqkPqPsCZOOPy7
jrk4ZpMD2BbS9XBgPwhO7Zr9BgkiHnLDj1GyGjNfQRsJeV2uyYO87j1TT6DYSuT3
gN1zCW7lpm8Xb+h+OKHNJkKgos45Zugzn2yBzn0RG0Tjm6wpq3JagfvQeUcWcl7+
roS03FFl0s+tNlLa2fbBpsFP2KaxUEGAc2y+r6Iw9ZALP4pNov+kkSuVxN0YzfG0
P6dTLpLibC4mkm0tXqgehpNDYIiKZvEy3EbCPlmJ2Eu7CUvpnW5D652Yelle38gt
vWmj7RtMJloPACsnr3u0fYxsj9os9aXkQoRuSKZUg0ZHcRJw5lhAv9526UHuoGTA
yZ8OTNqtox+KRVbIE5j2I4kbGhajGggOGyLTvEBXRRYZ6dmqjk58/AFUaeGwrobb
CKlSRWivMDWFGI4EoiJHAUY8tcrGbEAdPZjOqkjK/PjJl67zRCkwWbcWsnjUzBwE
Z95savv9kxPBXY50VoymzZ84g1G9BiVRQt7052ThimgbLcL0n4faqAjkXpa6rEb3
6L5saQgyk6YFxH394JJSUB7Dc7JY8K/Uhj25BJVB+1Zx1U499y6k9lLZZUKUhA1O
r7WDAaa+3ojPrGuS+Iw+tc2m8eBUWEA/A04hNPmakJHLc+YikeIlSHvBXx6daTh1
dYwRUn0Dwbv/uXfrepaYtVd79CP1kSoRPpmCoPmchRZfLghPHtoCu5Xh3EmyGuvW
yW7pIUR4E2/2z6jzGOhlw1rWk8GMA7CHu7poqJhNUq1TvgV7wEF3HG7UKH3x6VEt
0bNZhE4c2JYIigaPZek+cS/DyU5jT12VOvFxOUNwU7rzdzC4Gi2Su+ojLIT0IO9g
i71hVitsyu1BdX84TVP4VFOdfclCIurJmTczprsB4ZuHBynzD9TRcmS6cdY1GZdA
u0vTXOUtfSTymrFqog3QSPL1MU35L+Uwtsmp7KGLjLoUeshS3BIV1bXMANpGMOC4
/uG2Brug7adg0Umt8Png+p78743y13gtSguy7SlT8ERTqd8pcey4otuGHUUyKlVC
eyM9P8tsNWG/Zws0cV4j3fDvFa2hpUUcEPHrT0XRUo0vuaydlHZrbN0IoVd5SIHn
PcF4VxzjPEq9SqblcGF3bIfp2UWXCtFxg+LH60WNJoBs7FsJJBNrMR/3MspAJjfC
WtDtLbfFL1dnjocGjoYlFRrR5fPZCPO7YPW0U1GCbxQBmzeRKBqxqLA26nG8ClV7
s9ztfjmc9et9A0qrQtmOno4TouDXO6sVSeatCeuh/VXgYEzDzUgWx8ICmw9dzden
czku1dFDMBMynrsFBj4SSpPRxv4ZxlmA0K6JPip//KAIZEBcmXsLHUOPRQN37GF8
CFDTqxRJC9d9PnYm5C2Lhj1/AqVy/eaZ9G4dlu0ieo8CNrCdW0jC0EA/4saidx8Q
cZkXoQqaDQlm6JqVC2Hl0Qz94K305eufEAct1Ldsv9rgjcFilQr8EYBjyaRJ+yn7
Q4afrYetrZyIgMSbDPpmQg1rtG25iFdprvSSZmawhd8dsNr5mBrWJSpDz+Cc7mLI
QFoHRXKff1ZSt8kdCp1/g/t/bkKx8URuyDgiaGQ88yKZ1ypAauTe3YCLEVAzW0Xi
O0HMwXNyUkOE71IFAfbaO7dfTNdY2NbVrynB9zilMIVRjUHvEw/SJro3u8yzL22s
x/M0z+AiE5yp/B+9z9/dKScKOE2qQMIUkFAlReMYL40X9HaaIFjsYZDdh9QMYR8z
2dwSI2ZocysfTRTQ4nPZOvU2tIdRzJX13Xuz5XGYJeJBCJ8H6E2ZsU2ceQTaF1qq
EseqC7zsSoDZZZmKGVKqI9l/xK4P6JSdYOivo5SdU8BU9gwvqJb5C2JHD3Mi0cto
g4eYBVO3pyWwhfFQhyg10ez+EEUDGxvoBv9g9JZ+aWR5/sNNn4OefENGqrvXMGUs
GtQjh/Wf1ccV7TTrpVZ1ta6mHKgVZecgyMjAfdJB0b7WwtsvH94k6CqK6mPa+rmb
cdsJQVvzaxBr0/+5+1Pb9HWptgR7+Inxv08OyFSAiSKgz+2B82cRdh3XkwNmJBMX
I3k6HqjIllCE3vC1uwC3Burffvm8oDOpxFGM+HF6pW1tMYXBUGIzkrYHoIsWtilb
/L6fBjeE5Qo9DT99pBHaf3jcAh2k+E79NG6CJLVwN79NmP+VgaSrgzjfKHG6rIpH
LjgOiFg30HR7CKysxN8q1R/0XKYoMihCNYYtD8EXRGL9UdvMJt45tzTgTho/RXx9
1EEtzYkn4ZxEl6VCPXZ6dfa5Jcse+aywvz0tKlSEnk/OXuZuqjEK+zgHspX11+2V
/Iby7rGxvVRzc6kQbCFBCYxU1ShMZJUnIXuOeZevcXrWMBS27bdeMYF42u4YGzoh
R6w4Bas5LxhzsbVrH4CNEV9ePBkZtNiszyYjjitQC8P7CRBaJKynIUmHnFSRwg7K
XC1HjOdLPPcsn07ra+XXa2bJLHTK4uHmI7DySc4i4NGUpIgasK6soBhFwma2ilw0
VZnHY7wDHBtsZnaBSbaqESM7v5RgsUqGESIkG+rkuqDNBevYfM52N/AzP+xtXW8v
fPji4rA08ramRD9SFCKDI5esR8lJ/b8OLp2ls86ZJYqstcSHY+3+5p4/OaqpJ2+B
kzmmhKwH28NEKuMRZI2VJV8kSaxs7+rLvs6sl4wDbKLXFsww4/wCyMNsO9K+x1Fu
9AJMervTrq2K15JlVk2yezdcNQ7HOgW2WVtu8BuQxKZJt1Wb1gLbzdBSRweRNyR3
aLiAMbby/GBDPPIXfEjWGv6oyJQ8pcAmFZj32yRfdTyhj8axzjvSerq/SlESytEO
hvqRpDPf52rJbjBYcvttXkijKvcGE2QkZh33nElPyedTPHCLP8p1BR/L2Uzz6ksg
k0g4FF29ku7ZMUW8wZcIF2SnCJC6jwb5/ko1co5k76sgqXgNR73IAG0jahNjfzoI
ZKWXywGgRPAJ1T2So70c09e0/bMq0xlA4oISvgu7gJbJtRG5N5NBR+2QjqM0b591
FAECcOZuO88VKnGFo+0Tg/k06oKJJKvHKu/qj0ZX+pkuL1GSqzXEqBxc57gyd7cn
wM/RPM/V44jxuSRsY17Yp3vM24F835gidzb8L7HQ7XS8qLHlJJlpqQ6LI1c7zqC5
y/mcWoq8eyEtxT259lsZ20QnfknSaLqiEQNC8Ffg25xjvSZiEAXYrA6HE5Gr60WF
KRuPgRy1vv6nnTXq3Wl2Okef22tdQBkzVs8NgvUNs7ifTX2TTXRi0rhx3DhFYkb5
F/a2+44GKoLuPJjkVdm668ObWBhlZRJmMUbpQBOPkW6Kf9T3TxxqlIpXpEeGQrFl
EkZTq9XwVq6zi/jtv3VMA8l/WOqDScTfZHZHJOFHIj8CYpfRg4Eo8SovsY6QxLMs
kNQdZ2DCZGf6VK4Mr/Ai5I4O9vJXuO2t3fnVmq6D4p3e/S0CedHPKVoPx9zJ6Dl9
OZ4cwkiZ3unvQTNJNtTXBEVL/strFN4eYdM70eByK9yO8pLLm8vQW9SWUGv8FjgN
MxRemrUBd4QGCoBIrh3qdhxtRGDZ+OlyNE9U6+h2m6pD7otwFAC7k+XYeSu+yZNd
nl4GWteCgu7ZFYqln/jP09mLBE7/eP3sUdj4Hg0cFJ9CeWGsM+V/QbM5C2zSjR+I
Ek9xkeybadE2VtJOpchSoJrOMmk9u4LsEy3oJygzznTitZuP+RMVlvAWk+CpQESC
FIpEG5p5sSrduOpi0mR6SPrsQrLT158NtPz7sYD12gz4UbpMVeZltSe7tJomYMr0
/SOMFFurLbhZMp02MlRsw9uBJ7cLo6Vp2tFZmjUAxLNosdew2gDWwbcqSWHPG1IL
oLewTsO7ksROJ7McOqS9xUGOgJXkjFdqv7SgRl5sVMGuM1bOLiwP6NK73tGXhKEv
nFGJqfcs5+Q1OPU32QtDwcqjd8mdTwcoGRJuZ27lUb901Z+329+1tzktz031Z7R5
e8k7uEQ+kQi12y6PidcpHY9g9sZpGSDz/yIdBcbdUWKjImGTd2wiy2LySrUZmigC
Etjs+jG2pNObQu23RzXD6JsdbpQoEOZDiXOtdVOup8VjfaQp8M7qZGitAwFOXOBk
4ZMyKPOdE15joYXIlX+CzbTlavKXhQJ4wCFs2a2bcV2IIl+++3siTkqJp/Fa+5zA
Wev/qnY5qxvOsweCvftgmbFDT5uuOosiKFYwxzxnvvInDrw+VrFc3LLMHxOJp1Gq
IFZdY58NeinO1Qhq/+YZrcy0PsZplKA4vop4NAVwyc5ukIlepxnlAFc5AyYW8Rqh
YJUsBQPbtvg2ol/BMmjaU/WdmNmgP+PQe85moLKS/sEheIUVVH+5/N4xYNbyKnVL
vxvyiV3WozKXw4oRQYt3qdINIGcCtPFq/vb1aRM0LaPteRaXTxUz2feBaZxt6vAz
2lHrw6AGxIEmjOI9tzbAlGMNeDWS2VzQ31JeRiRrNeL9iFbE0NErnPDN6TmJ298+
J7ZnHCGK8iZY1tuRrm3IjRGRqckiF8/fI8cyUeYB96Kq++j1KMLD/mzNqmU1hjEy
sHWLfVjnc7wFzWjn+1Od9Itb0TvDGSmdlTgq7hgsaVHtAaK8Q+64t33VnzVHK3BO
HQQu6nD/FlOmu2m5tvBlVQAztsz5Iq1ncfBqSSY8w7IIKgaZHifGfdvh0h+WIA4+
XB3qmMH/yrXym4F6TIFfT0OmeaPaPAEy0ho3oZV1d1MtBHVdL59SiuXy0L+vkdCm
Rh9lhy6hCzo4lUeLfJDxaKkO7PqqF1w62CHYjsy3IBDp7jb1P5mEr/Bs8ZOjdOHX
s7kyJfF/v+zxBNcJFsQVfcQJKzonNBSjM0b0lg96It+omP/AcNCVZ/Ro32zbVX8G
9vrSKOteTSQsrNDHJZxBSVWU5PftiFjw7NPfo73Zm+1AcB+MakbTEpfR3y/1Nr2B
K4odTE1zkdhDh2Xfd4GG16TLj6T50SurEiR4/yy19tpJ8bv/xmxvSzyP627Selab
mjG1XwNZysE4fURz8l64gezJeZ/dmrZ3Zn2aXAKjlnnRbB4wuH1E2gzns4gcebX1
Z0cPXy5Bu08FTOzkyYGQxOz9PPCKfLZvkjpFVCiENojwHd52dsJ2F9zA6ZMxC4iz
zCqQRbE8E5Y7pBgHprmtfUnxfwVYB9WTwDF7VmqgI9ZVb0MgNHZn10p/hfXsTcQU
wIRiXEvgAKgwhuC/wMH9NvvewZOvrFMLoRxdibW2VGrzRKkUk9ZO2k7wIIjvhzck
XX7DNezDG0L2acB/hJnmdtH0E0dfG3cBxLeD1iR3AqpaFF8+mzR/ViY0dK9terxn
5hsCuBnfUDI6JrTSOEDesJfRmwkViNlU7GSAobOM9jhK6w1cmwYSIE2yV8Ww/XOP
T3DmXG4kM8HrbUCWZhnAOqCY5ZTWgSkQRVAagUierTygabizQyErMOtnmVoVVlve
dwH2bi3Pi4nLjstAVKFORiyi14lcOztM3OcIqvHM5JbSzFGSMProsBupYEpAK7Mu
kGLCudMuYtYK+YHJnyiStYBsP4Cr0RcHUuuGdGn4RkM4G4TuDZ+gX9byFR2ocPRi
EXLf3uEHGnDfGpAkaw1fx8s724vL2HQY0xTdm5TQV5pow4jTf6+EV4nDKSPllIA0
1P2pKovIHuV0wdiK0RcybeNVP+TVp6AndjG9tVjDCIZAX15alzlHcRyjf7wHlP3Z
AUqyX1tyn3DKQVq4Gu8O6EPnlyhGpieIjDsxMknYTsTCXw4+x+woGokn56PeoAKC
l9/yHcJv1A9H3djm6gApG3v5V9yKgPUvZbabMKQFE2dcNACXWhDmX09EMYttHJ3W
5l3P0W5gmeLipdqG0n8naZKxKNbmpjV+KF2GfZ4PO4c12G9/Mf+HCnmGnQiye4Gj
7yhRJmNAOCrpHCjk3wqn7Qrs670VmLtTFnKOrY67TzhKrOy83zZ5r8gT3NiY2on3
HplrX6r5BE+93bFOoqzKY3bmUaJTWe/UXdEmnR2huv6HpUlUMtJ3iAUAkYhVxeh9
/iDd/l6s6yBbRWtCgy7ZI8rYTtrSH75PFssKyJgrLsUrHY3AQrEAC7yus9d2xtJf
irrXpqwfVrGt55qUP0kNMd2VOfSVhQqUy9OOtnwrNh5GCVgvwkqodnJsVNJySQlz
gD6jGOERE6+WKfVBg/0sz8Ir7Jfs/59OXl0cxfZS+WUTFkKfi91/yJ2EtQh/iKur
ZT0KvSu2LH9PBEsPj2yzhTSWq5HqfyK92nO8lgS+cwa+xD7O0zKM2xUN5i4AgpH7
GUKGGwVT3mqb0Bt5y51BJ1WKWswo/mfovZsLHlt5r6iVENjNfoZAfqnSb0RIxk1M
ZcOja3W9HvQlZT2XnBF1B/ESQ7mP0K3osfMybTcCPr+20iqlnROAmEPGS8uxxmtr
100rgzz47Yn5rTU2eWSGSt61sDpxyW9gASybJLsgIJH2eKL4eB5DKgOlX/MTDgry
kUs6i+WAgu1YOIO6lKmjbMFqBoS7MY54xWEt/YnyPhpcrSiQzGWlWrxjdwgl+8Gy
kno2vZLZXscFZjRnYj+DAoRjH9J1/X1u6FZ3qCAmnH4dpP+inJ86wGcFwRmTe4yw
pIUXRPd4YidjVagxgZCkddGJVQdkzyRab5bwiM6MRarUOgXqo1/p05PdbtetDOaI
rtQmX0g2dorEWr3thTmCII1qO2EfFr9osRsqr41/N7gic5Jbzor+2Bjdxvhe0Kw6
zZn+6x48solQMB1rKX0K5jKH1X2LK4WZ8FspiA4WtIq+3gTx2H+P4HAUJ6RaWq2G
vEgPV10qlFRNDs+vkdNotC04kBzLZLMIbqNxRW9/t0Mwp04WUH2ArQimkCNBraII
fTdmOUFaC6Or32f2vtrJLgyK/X4/SD+pelMK5IE46iVUiY6g7TGRcAfpW3R2nnAG
M+GKhfHpLJMhw3o6/x9T9UuCzdlQIKTnH3FuqrRg6EzRSP8gRNqzD86JNkG+2BZ1
HbWnOanbzsP4sfDO7SMMG3FIMRpvQLFqziK9UvVsyX/IsCUD9sOVFA43H8v+Cinz
vHFhiYGKvKq/hXCpgj9my3G3yQigPKqTHbQaZf4x1tD4rCwmP92xKKgzKq3ZqI4A
LypSiygpOoiFzn5s8NI4gm+ejuCeCvon7mPWfCmdeRvN10jbn3y6rB8R13ArIbmb
WcbLNUjx0S8pQKTp+0ZfSgnP/Pntmg6ArePSTXzaNOltvWT1spqL1X/2YrWUgNLI
Du82QpX8ISfRUxzR13UT+9h3mXMMyCcEIwFHreg7BHaXW4i/WkFrj+M/P4lF1I8I
la4gbiq27RfxRzQJHYGwNHcfqCP9a9KHGQAyDLiSQu5V5Fy1NlGCI1iJq51//d4l
+7c8zVZGGyBaYvV8Rbm6GL0W63xQx8MV5eZQ/lxlr+rGv4oQB85c6BBm1RDOyVwp
jaB8bzEj/r+J1jh99FMB2PkIhUudYQkUgwKCHDwQ9MqJQupeUOCD6gVU9RzvX35I
krV1NGIhbGjS4q5oFzXhPkWutCBtBSb4nQXLGE/J1yZ+Jp4hUbTWaJr/UZw0toEs
JOpzw3LogSSfYe20CMXlAdJSWpYL0HOQ4daBLYLy3L8RjFssEBcfRilLmVe2Tf0c
4RFwyquxHibGfrFbdOANuLlC515lQ+XwcHir1DdxHcbqKpjcfDuRi3dZWKb3pr0i
CyRRzk53Pot5v/Yx7NyhFAemNVpz1LlKO4LvZ0PAmvogER+XEKY+LlWFsILVrEjk
YiX+Ghask155imYp1xiI3ahah28FO7VMkQ4ISvLbDDXBYlYhLraNo+SfDGINl3H6
hFP2BzP/Zm6thdUxXNuLUHcQXv39LPIRU1GPObHtZwI2SfYIIyHjSYK9oUPCNkDY
gGyLmD7bnjSXYcsSOwvnxFAuymbfGK05QYS9pkT5JU2f15eES+rSUqaShOfbWqLj
7DBqpjXcvDfnRZnFnjjljN/+TgOWjHbSbtEm3AIjjrA+2Pz/GfIEVw1+xxtwGh6U
cIvVpgDYfBwtHkzmaHVqaY1UfFlaskuC04viwtiSRzS6CelDJUSGTBxHqFx7Ef6j
KviyBV50AMqvWHO34xlRVfSQ5KEwZwrzaCDzzsUFxIn2MZxGCoNLC3Iyq1yyVP2B
aZcwgvCU9UE7vGsx0qO/HWwVGpdv2HuJG+L6Xicqpmp2rj/J1nL08t0tnenZMES5
G6OFPjVif/n/DmYH36m1eywQJ+fPDDnnSXgzO3y+Li6AA00Enl9Uszfqgcr3+3cl
oSXZ6PUQfNIVQvcrtZhVTY2OQNFTzvisOlXxot+bTSygLduMH+7Y2Mvf8ug4MqLD
QSuAN1VNCkkDCB5NIOIZhmh+lMEp7VxUMmg2baJiSgBnDJjBphmeKFrD1qyZAVT7
n8e98n9UoPqLPG4XS5nXRGjRA2SGvmhDscJphAFg7GII0cDLYsj7e1QF/Rw9e3PY
jns9rse9XN8WTilMNf7fKQMrvOOdHQav4bdFgeW2RYLERVc0QJ5+FksQKg+WLMj9
tngohi1QXkvieb76rAptkJ0/unuXTKTjehyCN0YBS4kNxRNmjBg5tkGszhWkSp5G
rMDtUvHXfjHrJsY93NHJA7VNlI1pd/sYI235cSIao4stIcAMTK7Bc+mBmnI5Jk5x
J+nCJZEekeCz0WJVEQ6y9yQsu6QS3HrfFRI3l2SbdVDI9od2leo/23HnIXync3bT
EHqqfp6dc5G6iVYFI8kO5VkVwm7jFWoWkbMWXEPCZkDKhnqTGLscMlu2dqV5aLAC
fI05KajaIFgyheNoJMKkc2qCOGsXUW/vDoRsC0zN2M8isxA9flwVReyIY3DOigRq
Pz/DxyjztBMbE067Sd4eXPzU08/p9isv6131gzjfWf9yqrw8iCwBwXSJLP4plIgD
2200AAxI3lvrZZJH1mRJKwy9vqiN4n5QMfjw4WCyTZ9DlaNM882IAk+JC4gqXeQP
8cCTTr2IdRqbJfhtJNkG9kQl1k/pxB6Okxz0vV80zqdzdS4/hyqfWFmIoVryMHii
LuDcni2QgkrqIsjsbalfPU9Qc2F8R9qX8vPGckBtHGf07REYb2/Uhk5wTcM7jFg+
Fnnhb3UQ5a58uX/k0PpGhYOsRZ3n6oysKozCI+0UqznEds/lZqQMLeRjmNcItK3Q
tV5aSk56TdL09YfUEIP+9ZWdbpsiH2aogQ8jnhoHhysGQcnKgALH6NWtVix0A3xC
Q5nmsaw+FIP7zZUt/WpiPjd4FKNuW7rN2RcMhUjh5BdT9YkSmMTijItsU8XHJTsz
beInGBSRW1bSJ1k+eDDARLk6BeJhz6IWCmHFfnYC0YBMUwSSfVMaQ1IQ49YHs+q9
2SWCTHcEhHKYRpmG723D25JdBm2vB9DVktlM1qz49Q+T1Zy0m3jtwjEVPHOv5d65
5AwFF9JsnVlDvedSFgv6VurHLdHDtRAvL6QcpfV9geirmjighooJN7/AS3vPJRv/
0fxIfH6TR9Hw5PjN5Q0MMKaoDykjVKh+vwbPT2vQxwYSvjaleRjL/YL27j2H808i
G5C+hqEvXAWdC+pt0i57DYMzCMnsdy1ISmGPqE8Z6gAx1jib3k62y+sbFFB8Z54A
5fIfVbITGxCQ2CP7KpspDU2IZ+Dt1iKHWh2aTUstW0skOYdWyWsTLox/mqGY2oq/
kteh/4Ry15oNdkrwc5j5Ja3CtzHmUj1FykNwWcm1brC3gyB6ftpfsbLlvmTGA6en
VEG/tBBX7aA8+3Vx5XskqdGM2rXT/0eoQNafFwj7/G/o9yBFZnDR1aP8I+MBCXIg
b0xSJ6bgtt+2dMVcmo3eZ3IZ1AVcRknlK09ghP/Yp+DODvwuC2iKUwuRfNi7+fKl
MZdu6o4jaGflXQVYDfDfKQZWuLT6SMVdomHGs0sQE9qPjjSK9wKbeXw9NIqo3trl
1f7+GaCwzEo4hua5JKj+GzhkMD37pp007qTy10lPfWS8lzwfFUJbWBYbxDgOxGQI
e/Ss4JBHsSWRFGxWewj9XK1KwZ9TSUeCTsfvWZCxIJeUKg/WslPdPIjH2vh8BkIL
8P0lAD9sgYZtpJoQBlp8g6axdooMGrsp25CpRdPD9gvJXOL0iy4+ALP1J8kuYllP
mXGR6VHMosjlOVkyCYrfI77IT3nwlYromYeFohecPrd3DIfIlNrd0MkQp8/ogxWn
uBm0SuqgLgIGzEaosWECfXdgTtGERebvRgmxp53wyrjH9gGcP6ygOaYust+7uKpi
2hsGniPI4/X4Wz/8OZHWRyhENU1l3Zkpol2R2J2xaWfHzJWMJxK46Y0ANf4Sq89N
zuse9sfylLKU2Ir90oiL/g39sMl+qTd7ntunvRD1xuPAUIGbh+rcQAmawK23Qy0g
N4DauzDjkga875v40K6iEBQLBt94SxNasQmKjnKgnQZOUZhoIBH+Am0kg+gmB9d/
nWf7SgRfAtsLep56W4HKd6S59TmVrSTxIa78Q8EcpSq6N5d3fxotMLPlyz1nJB7f
dWxBuKmL1cggWtB2fqYBIBANFSRBoXGmBFIOz5zWsC8fFn9o4tggPA0VNDEWtrfc
kJytxj49i226wgfXgLPahFBEldkTdh7L8UUyr0BdJbhlOxX/3C/n7e7eTMmRaMm1
CqZA8DFzcVbB3ivZVjVHeKW0BoPutv+9YRTCZ0ZWT2hHUYp0dW/lN4Ecy4uPOq9e
a1M154H0NWzvb4rT/cqUuEi5ioqgEg+KxkWL268TUy3fU/tT4FA50QeXsImBZjrk
NnBHGiz+UmzrfAwfLKapnZatJwyT7ls8gqsCw3xbTkARreJZJdQI7jFl4MKfDyV/
8WWCInDv18CSn8FKHEQ2YpTy62xgKXRRj9M7ZGiiUiILBtIWwljLE2//UoWVqrJB
YhkPOsangRsCPl7QAFlrFQi16IWdLTc7P7V+Wr042lAXxiZq+3VcfzhpuY9i4Gxn
Rc/QGWE/yOzLni1sn3CCOceFdkA7yUix8LZXeanbiuWtvkIjYFeVEluf0CUUjtbt
zrTGrIcYq8L7vRWget9EE3L6DNbXVUUCvitt+K+pCl6gAj2AB2qG/Fi/qxsckA2l
/Dgl7p5JmGWI3LSOhoSSdH5lzPWVBzZ2Xdu017awy5DEl3wJT/dwizz9bG7r0Xsj
qht5CvWOnmLHBofP2hXLWY7jHwMZGYHQNIqnwfjLUTQDmfMih8AxbsMkhKgyi7vx
SusaP4LbzZ3ImpuxwTqxMZajZlu9tABMcjERAO5JH8cPCFr8lRT1dBAx1zHK8za5
LuWYRqTYihc6YRRFFJoCHep/cU9KBMCBPMa/JmLSVbY6Q6yX10cFJkoWoQ/gW00J
dy7/H6tz8opaZxAURF+N0PLmqukqr2S2mcbsHPqZH+uG0o67075CIcigEL1uGMfu
gGGRHkM6MrbqyAKBPU9xNdKbI18bDuW6LnCuiwkRCVLALc+i5oKee5JfZFAOGyEc
u3GFK6IBXhTrghQmLcds/HGJSXpzog6zlPRN/mw2LI/ByhfSg7ASHpnx0wJE5mq/
ImM4QJ+0Vd/rm6KtZFaT27+gDhPMNuSML7WRmV8htUFOuWMIBx5De5HqIxX6q3u7
qOUBTyXlXKPUOri7Ou6dW8z5ULVWOif3/4q1AjTcghCDEWy2a1uuFFxIzQ6O14MF
Gja66nH1MG+hg1YHf+KtqQQ9aRgeDpdDshLOGEsYiIS0bvLdQBgxoivUpKr7NHFo
BeNk38X91Xd7EFrDIfZUaJ7Dj6wazBraifxg3+WZA9Vg8kQ2p/ygNgpoIOOs8Y6S
pF3bRoP2vDSELo7TIx5Z8I3VkYSMaeXo7OiW8TyTxc9ceJsG4Dyw8YyGlpkQjf5g
KUNQQFRtUtUJyzVl98+nXqBTh7s2mWmX13HSW7olaorXG3CCcCxkgBrfwYlG4H01
Zyms+jymNuj2s58JMsOYZ8/8jzz83ABOApWWIGz3/z6CZY3HSLDv5iF6UkAEF7N0
WiCmEIV6FmPh+z3QpvVsfmHKMNRSgwSAo4bqK487ef/CAX8uvSHvaId63KbQ0T+k
7HBdmbH2Y6Sn+kyaOY5TpUgY1kbj1CkSPH76O05nPH8qSYoNj8Yqk5+drqt9H901
XyaaVkhXVWjE3q0M3nFGGkI7FfKCPm2NFSJq5ypgeqmKbCIEHVv4BrJueTcrd0SO
0LIsyU9OtN//P8mdg/ThatBIZhVG7NPJBGd0p3aYYq9213g32FGnCbcq0U4PcoBY
dCOIQEnbxzfyzn/KJNn4dHMoQlRPglT8ldF07AuiRWHet54DsRnq/Cr3AhysVEu5
RZzMP4vE0QnZvtxBTCSaQ5lLiEeQ+8KQfdk68xQw86wdSmnnszCSCFTqwwqwS45I
cpfj3zpctlkzcguZbC02Je0wukGUSwObm+/uaG+KWAFF9y+s11I/L4ck/4j0DBTZ
+k3ref4mAS/flH1nFzOs9ST/yI3Uc0++1EEnXRRE95Nc7sIjVQhbCkUYHL/m5/3H
OrAVS+wiyfkuqeJE2Af7KnznbhVte2+y2h7uo9m/eBk1C8XORsADmu//6DebL3qA
2KnkkXUhBVWjbra4ujRW71kGbF5NGJHUNzk+5Q5TCP/wPKVBBihin7QNT/QSyT6e
Yg6Aa4B7lBYiy2MTEPOnRDBFF3F55tdtMCtJ6+A5sbl6y69U3D0k/vobva9C4H5A
wsEJ0RBILlvwp5wUxusEkgj5AvKSxMG7tRNtKl49Ddu5gj17XwvuiJX+tICMMXAo
+8Flpk7VfdvbfptM3o/mYorUm71PoF0NpZYGwKAsZTDfkGltEgfHsaVb8ttk9bQ7
s6iudzwwhJF15ZE9GNLFVJ2GAQJ+2jY2YuMJkeuH2wNK7d6F7AufsAOShMiu+Kh4
m1VV25an4FYkOtimb+6DDDuBBJXGY3cgafEFdh4/yVVOzHFeg99Ysht/o1AhIDlr
q7g1OSPl+Duva9gSN47fWEcD5zayp2Y4nGzl5rof87QhpkUO1jBC3gSWvC3lLoMf
1ommVh6yA6rAcN5C/qxAyTMBkrNqNsOnnc6vGx1eyE8+pZhM/rLTMboU3Vhlj6o6
QQBCXoA0yjyNll74n7GWQTbcW4vBPRYWaH18rS07rU/a/jn+57NbDrR7nDljzYN8
wpO8qQ+B/xFkOvT+njID3DISFioK+yVH/kJ5ycegVU9Oe+vtMQRKjr5c9ibh1D/R
DLBmeBr6JhIILV0AdgStunGMI3U5WXpO7PqIO4kK91t5eDSYr/cD7hhEx5op6a59
JiuS1oXBt2WwOWuK28WxsYD6f7nXs5AO9ivlokowOeGTjFF89V2pzHsGPpJp9fCc
BXbdapOO73Mj4bf67u8AiURe7uKnNnlNftxe7E1etWiPnFTaNjagec11Fdd5DN1T
U8tHJfA5cc4t/L67B3JWZjGZCvXeqeQPPSI5dQzUiWwcb6GeHk9x/IhFgsNIA2qP
atzNE67QY5GUCFluLcvzSgYQjByZ50ur2rwKji2cCL9r8uEFDFC+cwBIM76xkwVY
99OjUc5LYPqSWRx1vmSS7IZm/7+fkWLoLkl8cZJW9GFo4zpAY8JD/G/SxRxsMNMr
7eirL/kJMzu63QlHqQfb9TT4KS9OcRP1auiOdwpWWtmAvXJK5lWEiPQyimXTvUGu
08rTqOKebWVUD6iVQJJ+hJxjttciHhdJA3HiJkmI4Aw2v3mCYQWfosjfZbldkKbG
kRs2KLFTYmULrEK4VsvYBbdzqksOjQBT2aR5ey6+afOc8evA1cXaHshmH08xrRZv
XEVEqNXRxSdtyW+Mh+voaGgcwW4sncH4O5GNLVomtUS3MLnsxDQWHjwLfGqRzkL4
u7sBKWDgWyzUVWWC33mkNjE1kyYdyXmHXn/XHeL4Ikbvkzc1Vkw2qo3bbGYbZnKY
16/jbLIr1JVcqhhIoFsXKvgu+BFiqMz7JFgQc4t9xZELF+rniK7M3v+9Eijsjxbh
doMQ3IT9f9EuJPre9fu7c8HomgRqaMlZ+liIC2gSCEKmfKc9n6Vd5woRrukHiSX1
rdceCkt9fEHXBQd5sfre47eaUXHREnHewX5fKEVvR5S1YJeuJ5cpwdyQWzBfpzOg
lqFMPbKZKs9GciF413tQgW5ffklvSrfcmDnJ3FRUyznIbptm498z/r4ZnvdSdesn
Xruwlq6J7ae/EhEAHGrxkgHp8ccf6yxFNWyvsQT9VAsOrTY/FEnOyyvVdpkC/MUX
PArZABS12LT2TNBxvZHA77wx/BmuZnIHk7OjaYUVNahwR+6MlynVlfOznZfb0xL9
ztxhBBugA8+22tYz5fYGoltdjVSLg5+E7ZHLLPd9E+/TUIFbYM4T7G6QaGi1zTLN
NSMr7H1o3BTDqnc3y3ndK74eAcuVVKEB/NOf6enM3uhG8IO4s+gxNDPXq4aEnkYN
TPZj1f6TG0QZgg0Rq3xxgxu9SrNwa6MjDLqOqmvv40i7K5D3bbEKqONnn+6EKXhF
BItt6at7KRLlHpRQq9ofanIiI0OF5UAGwS5qo2SOa4I7onF+xEGskTyoEeHVl2UF
PQAUkJ78cqtUkPVK6YVCGnP2fwEZtczE7UnmNj+98C9wSL/9Cs4Ie7glKtUf/j32
vxDuybIyOKEbpF8JoXmvXVV4tOVyR+a31KIMOWsWe28aptG9RSt9VRJXZ57rIlWv
gmxpMZRi/4EQMrjuNoMvCVZcvPJa0Cfv/MMC70Z+MzPSshBCPtBPhM0WN51G6jJK
MNNIbILUWE29DB1o9rECLfKjQtYo9to3EubdLE8F8efP9V74Yfkf//V49i3OWdbD
+IWWakoxLH4ecWzmRxQIkEAWFllHL8A0LRC8+fx8y4k40Gg3eh8xnQV/49owUiN5
i7B8tzoSFqvLh0RJfKzA7C+upsB+1dyjNt8QkGYRMLAeD8Pvb8D/6drBd73BlUhC
h4yf88KokfSVyTeiIzifLRe8gZESbZJW7Ez2V+AxAk0fG9aLKcminvAgJPx2xo5E
CYfdJ6l7NWfK7uLUD4NgcJYI3urIN6tLOenYZiAJYxtMUOR999BC9ShH+7ILrTEs
P148ZAwYtJ5VPpthqUWe81wzwgPq0NLLVzTLgULNcMRVgcesEfhykXhQouIFRDWW
QbQTBCYceZCL5jYNmcH4kE2TmxTDWwkHpbpbCpNlEOUi9+SGPx7uIB/awbMTE6Ou
6jWl2E7k3h5Q5VDx+PAXR1KuoiAod2g42H+4FIvLDIuIBkUnmKJS2oq9r9f1+xpz
M/PwUdpIa2PCOkx9ZRlbzXY+9SVZa8aCfVZAc9IidfSQiqd2QBtApcYVb5wrkibI
Bb5H7iCN/pNMz9ak7+B/fzc69TQVqYdEU27Tw5Tyy3rmeOft8aFczGR3BiWMwCzS
v9hs6/R+6KKE5w2Vj9cpbQS1WedA+7QjYxmoS2TnHpP9ykmY+f01loc8Wsk9oF4D
vUDt0DIgdoNu1nOQzRBG74XqxrvUbipE9wEFx3FT8J+dQmmLKI21FALOYryUoUzP
zUTktxdA56+kB45bSzyfpkpNp7VWP1hwczeCqQI/vGzmsvmPp+i0ogbP6BTMFgFC
EIAtJVXJFCu2zF+A1fljuKxpoISjlYlDN/bvd1Ng5irRuPmoYTtVzSDV4H76qgjn
5CiLTuuUVYZtGtMKDXskz7xouMxJgx85ZsLE1pdvO8TQojfpi7MBW1ONsQAdo6+g
R5O2rBmh+dNN+K6723zoFlbl/G9gEHppKDYvY/ukf2tKnPrbifp6sFnM6pu2IXu3
Ma1Tk60paoX+8VoZ7C6HIss+v3YyV81MlIWoo/Gxi0XUC0u1swLnJksJlhJuTeWQ
/OxWd1F49lBYxbBCQ96OAdYQD7vE2Y2TALvc624Z02J3gGJMmbOiZgFqmayWE5q5
EE1fK2XdEhQWo2W68AxsXIVdYwD6hseNUIJTMblamdKl556pX0dk6Qh/EG261ST5
nG+aDzz7xuA9B4xSczOTYi7C44hzozMlibF/4GFDcREqLvBQ7ZbE9JjXvd2JrNaa
sjmAvuBi/TzeRiXPxgTelsyrjdcjZqDEIKrZmVeffgbjoB9ytN+rRCGE9LxKOYuy
TKi/llb58APR6ImCj+SJyQfYg+9AnFrxS8VJs95wKeoXDfm3uz6qzjK2qeivPjxW
v6I5wfyFb9J1L6SBfnGKLoY00XXSRhNMjbcD5CrOKhNq1G2GvcB13eyQbiK1ek+R
9kenOScs7DRZO9yca/Q1cNrVivk+bUC0NFwdPKOksXW5nMa7xeDpxycHZD0ipEUn
ilaae1QJ2jSorhDuCWPALUS4D++wuH73f3oGDH2JfTuSReNXQ54Gn8ni71Cnno8b
Kms5o8T++lAAHv7Q8L8hzKL61S6HPVTe+RvJWgDWTx9QgHh5WeZ8VR32d8f46uwi
Qd8Y66nb1zmLatFuKOoBDGr6t8Mb7EswQTA/zZ2ngpFpzMN9RxmUhydpVpeLV//x
/85Evvzrwkk0HnXdIaUIa3Nri6WndMUtG7J0mpVqINk1n5kqzf4H5pX6q9+jE4z+
toNlKrbCmAWydlf4aadRyBGlPfTn35pnqCnJjbvbKJK9vN+56fy+2zKv2zM4KZKU
UQYkAqMbhhG9PVAdurXEdU+P3n5XNGB6OPTSJ/LkrKtFILsrkdsEqrl15IsUYzSU
QQwG+NIA9rw8vzzFvnv7mRY/2wux7l5bBN6bp3mIfwsQLR3ijKK+De8qjXy4IBo1
TWffN+Uo1d5gR64H1Rel4GEWo/xnd81nc8+cpsf8Vi8gJIwszzW/1vNekVvmc/OM
3mUc5mgINSYPiAYhFGmjaB41mXieBjZrrhh76n6IkZ6ALyfHsjSUjRMcYfBVQPlB
HM1GH7Zruc19lRmR2kbQdxv/EMNdc0xWDFdx5CXaXnf0M7qmPdaaTcHbLKThK1J7
7b2W+bBXAmIKz2f7y2sTTOwTyBBuZpVyjguRSmhrlHnf9hHUgIvoT32cOD5AppmC
pyjU8mr6hAaF7KlBH8c0xdqZHF8DOonA01CAKLx3C2LlpNtjK0z2zcsi0yqqQqh6
q7PlnFbiiAcX/eDBH0J76EOSVyoinq9CUkLcmW2sJ5j34Y7WRfxFikthJt3raVwv
IXBjH4VX/kDzF6lC9yWQcLVPGLKX7axh1bvO7u/ruIkHKpOLQE4Z8ByGPv9va3vN
6bAD6LSlLkUCZD8VrGDMJ8kVQtd0bjAJTThbcj5h14o84+1V5YmdTwgY2ATh3G+L
b0aQcyevDhVvBiYa4+aBnCLwk+lNTLD5EJiT7phO+KGC+UDJc5yAE4wL10knGmp7
xujt8xn+88NzYN80Yi270ye+SNEbz/4Mookg+T5qQRouVD3mJeOyV6kGuZgiyJeG
7V8VS6dpHmUkYgykfUfSa7D66spuK6nqpP7Xo7dgG07QwKeREXidmgPCCjiOONkl
ww/eQUbgEkkg7KxCJWH8MoyYvtgx1coIK0UNWdDj6RXdcIGU4z27mQOtKNbegLcB
Xrd3Tgncfz4m44HBFvV0mWqfXaj3yuFpZj7bRSs2ABIPGEZ5kBgwlkBfqSW2Cymf
E/W/U4upVx/xhYJ5gSJzl45x5nL2do0h+d8LPspZqVXw5OPmJBiNxI53qMjaD6cQ
C22Vo5SgntOJD2OriHiyHOQQlvsfqxGHUSuCi86d4l69y0p+N1CKhz17riAd7UkS
077wf3djJNxTgynOD0VdCwNOd3tJ9pZ+mHgmtxZBQEiINNfF2ikIWkOuidghbwkh
OkjN6CnLVliMLAec4w/NU4SK8Q+4MlcTiun1PAky6XSYScjpCTCq9c9iaGIa8d3g
RbgUGQ/HO1asqvbfEFi0lC7OtAKm+eLGFi36Fh11djV/yldVe4IUmZumiPz8P2Ae
d5hsg16Eg1sV4424MbOU2hSlGyDhURYAWY87vui8iZgov5704ZvUBIdQb+WQq65y
ApLricpFzAsifckSR6WuVqMUMxzf9PkI1XAABXTUKls+6LX7llGnZOpZqK5ixSH+
t4AoVBzdbfQNCJSpIlqn9YeLMk1zG781DXsArc2l1zcc0MU0fE+rqbHJWdvvjwLF
TpX3V0TPbpsUd+bpvpnfCRFG28B1cBqvbE1/DCIDiL1NeMaS5QJVMwGxmwx1jzfU
snK/Rh4A+/kXoq+uSGF5TXgLIQUdI8TEocYkIVjzs6bxN4l7Rr/uZvwTRXX3HMeb
WoZyzTfdW1R5UjLg/2AfrDjiN03lRdTqyKie312ftBa6mzEDnF2fsyKlPLCWvVd+
z0w+Xl4BIYb7LGH3G8fw9HV3bH83DOQNDxn15StGCicyF8+KxIv6j4wrGtrBl2V6
BqdAiYY3ise06bJC9gBFEWHjdZ7zlHhmjWMfbaUBZ3VRlylCsNPY3MrdyF8KsfJe
cRodprUk5J8PrR3xLhiaSysJ45IgiCLxVxocRWKopJEbXhKK/2zDG7wTqJDFAClw
us5m+ZDfSfMccFGnVJt/+RYfxFy/b+c6VYoomCh+1e73k4YCpNNhznGbhUQxi6OR
UdPtx8KcSbE5bbNELf69t9ELM2irniKM1paClQhvWdKIFNrCWkSLZ14FCqAvfn7U
448NdwO0y9h51FNocpK19rdDcXs1r5ltdTz89tTc4HsFYz6fdo22b43ck68wpiiE
zZSPPIKeBmBTcwXvzf1/tsqCHQE+q0zcCn8z/DIlgcQ++ZLzyOmx3zecHjr6EDWE
rqSNjo4t10iOhuXPsZAfHz56XaxDSs4WGNoVV47aTu304QJrWcPwtg/Q/wmLwJgH
QGIFfBXRlbexpjuLN7nQoN/wCdtH47/5nP+q5BR0F/BvrfDRY5elPa8uT3EEK07S
bYPPM+lBs/X2g/c7f6Mb1qf3HWNvX/oIOgpRZIP21DbYQ9NbpnMnC73SHsdiZ6AW
wp/ZzQa1r4SisZ73r8A21n7tIxDRUNkXc9fWZRZP1maLYsVawvsdx+DpuIkvX763
awoyTtz8kxVWF2oDZSsrnNOpFPphHLCeNxvt5QNUKoWh1PQI8P/HPrqiCSLY5d4y
KxfHi7yXUNkp8iOluNZ/LRUxQ/fzd15t0oduwe5IWzBIWwjiMbZealGHhUzoY6qV
5Gio0LmW/F3B5PdTLMQyhW9quOB76PgbY58VIiFIs9AfSO8pgOay2jFbCJ1Nbpqb
UCSnWK5vp9pb96zRM1ZPwFSoOKa1BD1n3Dwr/GDJt3vggw52eqyhgcn2mnkQGc3i
YItTguMnSmDZ62K1dX+lvsunLeC12JqHBo0bnm0uzYFnGvjXFMKO74bcwIJ91Ebf
NBU6nSPGRmJos/z0Od+vwzn+UhbNyuJvTkne5AJ4REMNQkbNWIk+4sDVBSKIb4TL
XKHH395Gg/6QN0F23YbMHFentUefaaZVQNeFBvvNuH9IFD4DhIngJrOKs48LbHsm
sIxmBBW5zjUY6rl+YMSd31Sqx4wxi+4rO7go8DG62/mV0EEPk8oLAthKiLRZJ7k6
U6nrUzBplzUc8NL9tkXifjmv0R+5EYYkdWeNxwF+W3aoSagpzGjDZ/8MnsmQ4fyM
m0V+o+eagStqFGjPaYYTnq/eOPrAaRFIANdoYYq1wfUV4/0e5+iIzbBSH5qR9ph8
lHVsKpz3iB6D7jZvrtv6LXXj5ilQ8pAoGYBrPYiBvOFyz7ygp6fb/zA2tjjVyuRC
fZE8NLy8fjOjP0Hfn4l/7osnD8e8QWQg8HG8CpgL40kIWgcrDqfet9uJ0lbRKrkF
5KHz+BrJx3HzdwqIC0ZWVumrcHamaMH7O7hqW2WHEs5Dq5KjnjKCG3QqowrLn7eL
3/3/IUIz2cZ8VZ5Z/myRrA2m+SO0S80rc6jPCk8+ggCnn+Vo3i/moRo2f4OB44hA
JAyX75U8xtVojzVjYXetbJsExZptJlY7ZeeCR91AqvlaAVqXQl2fOvHWdB0oXOU9
/Pkl5bXmblHSKO0H5Ywm5c0853nBmx3RWsH8XhzfOZIoNGoFUW2fYc4E59FAD1xQ
8FJw+0BjB5VYrJ8v3aDwvYFWRhkAQHaOaSc24Yr/inKGx47F3JOIFLTds/tNnh72
uK38DaU/vw7FNxG6Tvvv3k7XWZpJMZ3UamHoftOf2QPK9RomDUAirT8L2r30UhPF
9ZcMDO15dTwPUVgKiOza0sJPuX/2OMeHqf5EzC1NcvivvVmfg+0lBMewN3Mxw5TF
yNAj4b7urUeMkN2XEJqLPLuddm3jnhm9RV+YRbT+lQAFiEwDSCzm05J0Jfp/KQkI
+2yOhqCAjaC+xyYR0SPPSb41IYYi/WoblXGdMe4MD8/uN2sWJMWrAMEj/bOvpD27
0n0k17z9ol33XNmomFYYRCV27vFA3ExfeCVpXtGiJ+6k/dmSK7rNdglVRS7LtEuW
uptMKqRlohWWWZ22hCUviH/Jd5/n/sF4mMLolQGB7BPuf5er/V09uRKkMwWmFknI
pVipCEKkz+aLjN/Lf7Tp1uI85y4wIO1LCEAjkbrn3HMoee2c0p0d9eJj5dukD1MR
QOb8Q7zUZTuNaSn+AUO4hXgu16jhZ4BgLJBJNATkKZXMVJQ3FIHq7NegR7jvS53Y
FdEDDcwIqVVKOrqGZDmEsl/8SSvHPUXvafr8uR8/v16ydbvLKTQw/T9rvuYRixFj
p3jzFHoMHrbydgdvx4Kk3OG7OOyODv/C0JZxzVbuMEU5AAakGgqXZejUglzIbJOa
gKezfL4ais3jdr4VChHxr1nrqpjG0qbFN0+RJOk+f4YnppcYzwXZ6DkuXlmvGMh8
pRXe6DEr+i24CUCxo43TVD2ktTovSEN+bsXn3BbQJV9zjf3pukpN3yJ6G9XLo89l
wRpsrsyMkwW+iiafFsxg6eJ51SrwzuLQ9Hq5bKVtt9EKaXxcwgud39WS8kAQlZMh
Va1W4B9qH5l5PSpUHAt3XBZ93/sIl0k54Hs4ddCMPTM6xoRPwNZZHxlUnISkoTUV
O8ssftX5Cz2QEFpALa7c0HyigaTFEAP0Kb1KvzR/b9qEZIqCEOoZJBsOngOZm4kV
NKS94ovagDW6Ia9DvhKL9kiYz3OVDTppny1fUexZK/EYe71sMj20UHq5tRFiPO+x
UVTSRSxHXSFrtMro8rc6kpsIDPpDfUKk8YyRrNqeHLkyYlz7fntQU6J+7HEjiY8E
byX6Bt0w48MYSnbzQky00Cui8H+35b6aUMkxGY5ITrF+usDJqgB7FnzI27XsyY0X
EF6goB4fxuMkyHAXdPNCBjripqKcdQ3alyEPlraTDQ/Bk/8egtKzO7XRnS8y4o/B
GZzBP4SvBt7lb1sZLAWJaKDSCDLXkhUdyAkLEOwnjxO24Di2wwlvz5V8DiHXBW2t
sSq9zSRS+PYBaZ6OpJ5EvxbLn8vAOq9xEI6nV7rTTUGEpWLM7fha+GcGWCNKI/P6
acTnYaf3l+T0OmftjAZ87VpzpsRH8KN/TFiXtGb2e22gD63VExd31QcaCryJAYTq
irAPIaL9+VYto6R9N/j1ZbCNK/OlTSq6ZP3jjU0anqB/LKOw0xAXfDzi0XtHQcm8
irNkfF9f1aCONwPu/QjfY/EUt/BKlXMzZ5vcY3SEWO0ZVO21FP3YG2G8gnBEGwEB
92Wxnb7/pRgq/ZkdrFDFKXDtwsUQEx5LU0/si9NvZXeCxYhqYEs9+yn/nanzNuQA
fhOj1YUL2UxdugpXbaiRWgKNrDwngmEeV22kjhOcMtCiCDmCZ0tHjIpu3g4/wRfn
oEbMtVvLo8QHCBrvgYQnBotFOs23wMFJS5/2MSaR3aBrJ8XcidZeGm/4XeAglOFz
0xSEwGA/UBnx94k5IIkvTaupuKN3EdYne1CLdgJzm4cI9S3380RngXjdffNXy3Rc
quuUCNOgGPrFXaitDbTJmXOSecAyeFIOEo8z8G9rtDA7ipUznhdgGLEzWwrwi/UE
GWi2dZ5w3J/EG308S6xFrMM43e7SjUA+7y4jJPjsj5x+G30LS2FDbBdUjtFyD3xT
nxH6Nn1xtHdI0JrujbICRaFoprxWy17HDb4wDJ64S2j9KAbLRThcZqtB3Au4aP/O
MGI+VlAkNWHujwmyCdYDSQzi+9rLI8u2MlyRZn106dABxclCgHADJZ0L7XbZLytf
DQUgh0D8HuIxOFR5LmxzQ8Frwh8Lc+z2Mx0b1itjT9QZxxXA1hDf/CcPPUSa3dt0
ZwdorijTqFwX5rPXalWbqyUqx4eCNyUnJsZsOHgdZKv367gNMnvFdq0+55IH2krD
ydAkf+FSEcdGze1hy6qzCOt0WaJETzuSe+Pg13e+y8NS5kVCl4qm5SxT7Z9BO/JH
nEoFmbFglMa2SqN8HUgNEBl/z8mLJwF1yWU9/2JNYWrxNtw0wV2b2cM7D4sQN4FG
wOKB0E/2sAGcdMALS7RYirfX4xeSzUE4Bgu3EpNzhL2LtzJSYBL79n/8v2XPzWJS
BzWyXniUfzUlRgThyTOtvMx9sV14Hq8lT9hWCXnd+R8YiuMVqPm2CJveICmdTnQV
qpQKuTu5ZOS6u/c0VeRC93ntLIfek065T95SwV0v7X2hXuqykr9v/016PvvHxJh6
y5Kdgje+PvUIt5ZQU+EaBHwQF1rTmGrUSTRbtfhjJQ+k5t4U9t0sqbxWS3VRdTu9
ZG9P8nr3ng8vj+Dz4sfcre8QHqwfAPnTRSizDu+6arV3YmaTkQsWwO9wZAnm+oXZ
UQnVJulUR46r4rD+afdenzJHVS17jTvj2ic6sNerGgca3vE7wzAx16jzyRd0SAb4
QlO4nL5V4k+22aK1LBKLasoOlOv2g49HLUgBLCgKZtdKDbQX9Cd0i9jPXPHkDgc6
rOPZN1Pgd+6EMgok/gIxxqCumLLmBmOy1Hg7C7F9XSjDXFNod4mvQi5OTPv6Q6ic
yuP2I3qYa5nkPZXpaB99UoyfhijURzMZaGBeWNdEmZhi8tlTEnU5bWcGYmxHCl8k
h8WExvX9MLfAZ+cAzEN/QO6DzxVCq2T3z3zwhsRxgXJe6KPyL3PMQ6LfhXLcHwJ0
8Bknal65SdB5WOOZe/CojN/VKZ6qVGOi61cfiCH4SsOqCV/SoBj1Kv4V299OmlEf
gX4S/Oo0GU9Lruk9PmNqwL54FVze9xhD+LHsbYJEpGRmFbRgF+bYCKsVoKThQIxl
m7yJaw8LCMcuXf/8b/M0EMySX/uB+R5B1QsjYr2jOBBDuhn5eTXR+5s1QNFEqZi0
BDg//y3wmmZRzvPyQbl4FQyZ5JBSXCHyQHxNnYv5LmW7v0wxOXmnhG0xpHmAW3sN
iQHA2xQxpzZMGGutAtU2JP+mGMmRYuv/9Rqr0YYioqfnfASI2AqbQPa2AdZPvckf
hVC1aFk0wQAjn4+qL4S4dZPY6wDC6MKTJ8hd1qD3bFeJJyXzEZGsiSQzhTwIgQnA
78oaYJEiKtdU7hA1oel6oh1RWQGeCK6mzkhajiqvc+W+C/MVAWicaw/7iSATbXQx
AKAvHcNKLhUUxS7TeDnQZCwe7agg7QfI9achBlNZ2/skl8ZpbgJStc694dvXE5YS
LxxNeIfqAG8jkDYAbYuJyylaNrU6NoSGi9Cw6s05X2B/V5WGm8l6u6oDElibeWcH
1OauLkvaM1SMqTmOrFnbkJilqwEB0ql4o2hL7+yj6kvcwWcEpTolV7iYnB0l6FCK
mDWWQw0zJw7+JzfF8NZk/4a6fKlDFDDChHqhLjB96nK4F8b8jHeubILxEY+u4y0o
yxP6+SlpPrjmkoThjLmL5RAijm+iNLJYSvVC3dFmntNjvTg9iftmPkjOTYQuUFYG
V/W8A1QiL8CKZBzASo0zMEWorWxIb6ktljyyfgr/s3rimFEbF1WHTg5vIeNgH1JI
uv8Dl/ihw7OkPScv4yDQ07v3EA/kyoQnwfeJqHe9dUhwAHzBSJxNT/cOP77dTJRm
swNE+T6hDGAJHFVr++hkylTNU57PwLLpWwNdT6ufvgs/GFSLZKE2V9W2uBxPydPU
Y5bkLqv6Oy8a42CJRh2oRUpQ5Mi9zJHQsPfoVOn2wqYZzvkAEjNKWRxPTMarZubU
Uj4xB4sLnnfqlNvxHT6bHlAmsmiALZRy0/MMskQPNEosK/LXmxNAFWS4PBoNj7ZV
bcP5MJJZBFS9aw/5g7K7rAidLrynVNwyqtRkjPetGWycCmhLgowI7vQzcHT5Z3kD
aP0cqBbCNjnYrRqmtGZy07HZXjBdBqtR+QVKtM2La9TXcEKkCvyjjb1rpGnRlK9A
xfCTuQUWgVcc9P6cmoaE/4wpenkZ0Wy+9N3FZtSlWITqj6C/xNlpPDaCcp0wqNV+
/WlNIN3pfq3g+tUMgd6thY5qDjDa6OB3Lt4inwtVfhzz6XWXuTTaxnm6l8st/p67
Wtww99miHUEMTSPLpUODSp9BNnIYxX6tlFpUtogLfcsujWlsqDbs4VpWNKWn4KTh
Rki7zthEcCfLwrMtCZYDnjWDyhcRXZ+E5XTJZmV5Qy2LzAPWnXyRY/jXPK0hwveY
uO7ezyWk3LsTjjtWR4GxEckekjU0znP2ycKLAAkC2F0fuNzTOGs2lL7D7yVK0YMk
PDc293y1qMzZV/zA5juvztyIbGved/piqaaJylH5YUiB7FECvoqei+FGtnMsx5r9
Vf2jV9uk5u5l7RXCVfv7aezCiMs6HEgJJcy8lEl7flRH3C2D66DMj9kKRdLP/weR
VT6uwwdzFNktHL4K/0Ly4kxUHcXyG4v/X/yBQlTl1b501bzpawNqToWu5nCJOdKW
PSh3uxWc8FLITMHe6UgeKEQWNFbwyTPEpp+euxnMRGnNqujcJ03gMfqnIr5fhLUp
Je5XFJv6so4vRQhd9Gy/kpU9woD1lUCZTFssR0W2ihrESyhw8B7J4UUi3zdtSYY/
REWn1j+fFkBDHjoqCNxzY03O/vVWZQbxMpoh6bPKJ+6HlwhUD/whB6CFvCDQYntW
8/fVaZVMsmNS1qK4Dwt+Oo7ZeKF62F8bVKeaQYs/CwRsWexXOexfyT50e5E28STA
C/WtP8zvNVdFIZvy7kYfo6Pppj00ZM+rI/Z4mizzDhgT/j47Zs40EeRpx6KW3Z+6
tBwqevSFxHoNsEzb7f4BWRh+qvdV5ItkVKseS20hDbZYA06DlvRCEHqUjHIqEqpg
PLsyUWAb6QqNEO8YtsI0Vq6x1KYbdz9ODvuHJXXoR5UyL5c9VZ19UMT4a66iL/hg
gP7EmmquyW485ND36SREgb8GNE2fQnLmEX9/rEnso1B4YLk3yXX8bQiSYWPbV4dy
3/mUJaGAHY+g6ehMwyL0EJZw1v1s5BYfC957eX2UTgtvkKcWwKc1ws2wA47nwlKO
XCSivlAYhalAkrLFzCRMh+jbjSfVMymg9Ypd7v4Q82Nd+cwCzTzIf0dHLFxlTpFO
nhYFJ9Jj5gyZyZF4pqIKZaBeX4j3jkLyb9AFbN30kRqfg642L9d7WfmpG/nxFBh3
B+LUIdLHYyzif1pJZsg0A1WnWXxjASeZSTHfuBVLsrBdKLmdRz7l6oB6FQzOyYzs
YWUaYzKMRHAuDmv2O1jV5O4zK/94E/SPz1/6HYjrUu7EuVxIP14+EwGH7Vt/7f3F
M7AypGmBrMT8ghP2KofC9J0psqmci2786aGpAOG/fUu8OB4OLaBcuBZcYLkEbzIh
ajGoYwP0LJR47A9lsx6/BcSJoscpbvttL1HxHJrf7CtiS7AfhWozL2Cs9/9DhZsb
nMa8PwGosP3CSF9lm3m4nTYrsMjxq/nAUeG0whVIktzKWINvoS1IPJCjrMVK/psb
BH/o64B22NjfZ61ATe/MeyyvkQDqCFgSatrc7VO70W73M8Z5f8vs45sjmfoVdWgh
pnbpChH08k5zpOD+uVZRmCq/iKrtGUu7+otuH4R9+eaLj9cYmnFnO1ZvGaOy5NL4
sDaFjy7fNTAc7ZGyhyNAfVo//4i98nAlaRyGV459MeiJUMjsH4BII4WpKGhvUeMy
5NY00aHUt0/JT3aFtUBSCJJbzFmA0EtUUCH5QX6nxvrZy51oW5fPWnoIAMmEHaM0
fgF4o/ix2ov1UxAlpyDs8YWpQZmP6fZnwpoNinUbKqRRQWbHTdfeZm6GSULnz9b+
k+GhFfC2cCFpuOJZf24rDHbY0EoBCgx4sQ+QiM5RkJYeAflsG5RrO6llsfCHsC+I
IByhQ7R+A3iGoVFjgNIM2eRbC7N8KgKtxjRWCq1aSsrXU8E1sVeOEYbJ86YV0UEm
vfCDFUwxV75yZb4OtVlSfSOCvEMUHWkK/CGRPoFmByhLw+DHTDpTFBV96TYs2lSy
o50WLl7GkCMGDrvAuLUWkXOIASgR3eLNQYZqOoiDDRro1qAVJMRHSSEOQa9rxtt3
Tqj+ReePJ8TSPI9GUNiVmzfBqgTKz9ppPG5Mo6M8RpKkhG6skr61/Mf7o1mGlK/r
jWhzz/AWxSxWAkhzTZJMRfZRJlvA9hZmu1rzYYTYp0W9Lyj64DSolW+C8rgArR+r
c4EzxCQJWqE5GQdJL49B6bViJoQKaGEdI4AkYVFQvwPUJyDmjvj5OPCmQg5UltsJ
l5A6mjaLwoVmwcc7l6qqQ8Wr9VfTbVK3nX+IHnSNFhPF+BESqUaY+LKfBUb6WAXY
cTu+si+TsimXZR+iN1QU91pUEZtnM/N1nPO30IZDuNSSp12WJg3OTFQmzqniilNJ
3JFwnCqFfDXNh5t6hz1KlI4Eb1FpMFJPTpGllfGnhI+uyCScTGH6FXV4ITA6/ykn
nam3mtvvt7e68rC4+LXZ3gi26thpPUFuC2C/N72WYRgLnA58qk7JAg+SjjK1M1js
KyQcDzqZSHMujWokEEIF/VIBe6xAb3Kq9GpM5WPgEb2zlykjZ66bSQApwwXY/trr
sqgNWvKojCbcRTtsKVwcdDnw4cs/DC4lgJicb3LVTMG+Np7VVZhLwMnA2i/F9oJf
kzBhwFPRFbs0/uZNX6rWddDdHHIt5L05gOaOyCB8jSCLnFnLaC5v6/dhIOqnLy3j
3SGa7MUfS7Rulrkx+3oaEteewX+qVCSo1I30hImajD4uJ5EHIDc2wTgw/d1TqO8U
NxepW0O2OY8cDugSB6J06bAucbncIExXNihjiTTfs8VmSC+9lV/+lWfS1HIoHgsB
VT8fREii1B1BwkJW53rNjAIsKc9hTFQ+wapMpQ+cM1IbUBcfSb1bHZr0MwOf4o9v
u2WD73pp8xVLz5ukRNLoEKSfDF8mVuhhPFyy1BJaf69aM4Ghir4cFCuK+VRU72g2
hP+RlZcX+VTIKEX2cpun5TNiQgRUo+955pkg059izdg/UBLwhOheDiOVPH1yfUnl
U9vwH7nqgn+spP97ZQeiAHt7D1RraHOuzuEwPQyC3g1Jf/P6fP0E5jRfeiSxB4Q5
9cF1AB4Z/2ZOUmdSASt7yLJZ3C/Ju8syVn9fdxvLmqpXk0xRuz0eRSAAMVguxmPK
pwZHJmt0pZjU+WI9/ROk37wBCJ4WB2cG/+0Fse8BIy2eWcaQuJATlan8IR3sBAn9
8s5fgE1bgt7q0eDarp6dNBRMFd2mqdyuUpYs6dOyxDp/5jPBxVm5gdkAxIPFWPHz
HcSkuzR/F5RyRNomD2jo3tNVrhE3dl9Hg6w/StSZfC5IEFxQ4FyUahwnD9Sq1qA4
hfN11qn9WKTK6OdPEX6m7pcWySjuLjLMB9VNJzQ2NCuVL3vnSxG4MuGdfQKwVpU3
8HlXIRaYJIkj5vXemEl7IoZEwMFoi/tzpGBJmHnvWag7GorpWdHSN1YgweOYaPye
O5jQqmDoxUIotTBJk6lNW5z26uP0s+0OLd9oW7aEOF0zlSmoJJYiQmzYcSr98p1h
ZJA4ysoUv7kg3ax6juS/MWTQNPTMWi+jIiTBxxKgZuqB4cOIDu63Vkcc4fjfnjfn
3iAtWWkiED+Ucdjt98/oz6aPcSmLaf0wv+0fOXNlaox+b2fGx5Zh2yCxkNXkJFbU
kzOEN4J1jlwwE4Qg8Wdhl2mcm/RsQJtKTePDoCacd6GPPWGwKOEYbWRlu+a0k20S
oRXYeboM5DMhsymSqgoWY+vziTSHk0eLsjXJQI2iid9UQhVjIoG7PvNiloz5yM8Z
ja/DN0T4HfcMaizbnHJ2cf671Qev5mp7lm0SlOgAtuMI+tK9Nkvh7R68lHt1O4JJ
UA8PrOOIZ63wHhRzRyx2S6ZKL6XLhDm5J77bWJ+3S5C1ear0gykSyvVdqmhJkNlZ
Az5KGXb3J97qyNT7Dur0+tXlYGk7jO7N/il4kxAcJbozE1UCq/nAAS6TlzggyO4l
zDSRbWGh/k/YexiSibha/hLTkC+fEJ+BjRx400OJUI8F3tZO5qC6MwSoe2xCyvtq
AnJOrkqHlI9cuPO/jxy06JCqOyULKlg2Rpse0bVHT0AenGkiEXCov7s2EtVsgRxO
yT0IhiZs4Jz/YlGSeM0BpQ5RRVrIVtaRPGQwV6ZJCphJK+qLwYMnLLvZtoX/6NgF
tBCKmJwfLnbxpGRoSaPH1j62v2toroJZhQ1ZFnipMyaAMTHNC66tm3+Y7XptBmyu
7ORgdVtiEODkO0BZelPUUPG1oA4+jBIB379zcy16B4W3Ru5ietMFAcsS5CiuiboG
1HgY5VZQfhJpf1ROHS/g04VRDeBraDKKyPCzQ2xrj707qvvM9pH1BjBojPKHP6A+
MsrK7za+vxbAQjSfzyAanNhLME9RpiOuoJnTF5MYmFjlC36NvLtZt0EXYVBWDLyS
wHcze/5VvL8YAqCHE65Pte7tiiynNF0R+fzkEwH5s03X4KPll7uyqOtlIjYXdoKZ
ptxbiG5LICygAio4nWXtcJ2vEPmfljuSXE3oNZYFy1n2B1KryogiM4WFrRB+QeBV
qHHPNLMCpZzCGJPZEld6KCqeVUBd7plmrsjgPT4gVdTFueY5+89oAoC7oIiSyKvz
VjJhcE0h2O/hw9CJrE97w6LnRSvyNQpy3rIgsgMC2D9UP+jeVLgn2GYXOm+/2Kln
D4+ftSqN47TupR2zPV2ILJwo2QgxM6qItKnwRXGTy6YKe0uZWLesmBfue29W/wCg
RIJRr3MIzUDlKMxP3tZQHvAJMBPYqIM41FXRC/ycGTKFmWw/eInqq+odhl4jL1+f
wspmqdGenwPuhWw1QEo+FvGBOlU+gfFyQHxok9BHajytLo73ggsdvZPFSngScqnD
dDH/0+T+3L46L+7ZU1f1YRmSymVCPamHRpGBZrOnaZqrYlWQP2/DsAvd4JcEaHpP
/eb0CBmLVqvChx/Ok8ZtIc3BWQOwGRVWnoWeTjZGu2BAFTP3sPymm6B84qLLUmvb
rCKOjn6wC7/DsRxROXR6r4vqI+UGq7/SFtaHle1dKkKd91fsUZy1hUbXo97B40tW
F1ty0fYDEq3lA1xVs4Tj8PmcIjEnUpQ4Vr6fl/UCdzbh/A2LbKt+lJ0vfwzUYiRX
uIFgEgjLdGQnUzSgRiYVnuXdTCk6t0hMWVGP4wLNG73k+PFTdh4nploEcGUMWDJT
aPNBoREddaqYGcoqxJAF8bGyXZX84lNGa7yIG4PHcPFsTqiLH/v5I5jprjDuc7V5
AWz1e1faTXbu8Uxw3+YrnwvNOUbEQ5NXP67jCgMiRcLonzkkfko3Qrq4zkn4GvYy
ayJnshyt8g0deeHLKrkWx0jNv8TG3oW7B9bLTBfjJJq+eXoMflt23haOfVXwl7ly
LlQLDRchslM450xukeHM04abqjEwy6P1FqMAbqd0A72hdgMxqZtzgFf67u/Rhd18
2KV4Bs8YF+ajMJ4XpRLh+Vh228iSCQGgsIQBqVawlz2/foP8vpepCKLRFDKf7RJu
97m1Iw6JoRip2YFQjug4TlCfIvCMoxkv55AcYRL5kXxJS8gqYTPSWjUlBBkFzoiH
J8op18GxvavTTghXbLrjnM72788V63bbN8bLxExzRglVGSwJkelorq3U0toauQKP
CuLd3GFFry0WN3rBdzplwm30tugL7KfTnKnO7S/gkqo71v9e509U3DlGVDxwjGf4
K4p5OByDGNcbMSUJNGxCSj6Fk5w/kqvYGF9EKGpToBtBAz12UaOVfTn1CwyVDKpN
TRkg2VLVk9m4SUvm36KCmyHChfrMyxF6WNbRx5BlQLHh8Eja28TL8cBM3h6DDrpF
mfgbn7AmVIs/fa5a4WHWbyGdHeMMuX2gUs+Ld37+EhYHjhLmQthvg2r6skUP0dQr
i86yseSMh/kAhSjQzgh6DaOLW0eCiia1PC3rFrDCBEVBJjgLuWXOtAeduYh5SDmU
Y6IUXVl2D5Z9tqljTUL9RDQQH8SkFqbG1Ob/d0iaRZqiI3p2yz/AyrNMUf3nhX48
w1O9wpjdzgd/3TwX4uH6kH/ogF0taU025/P3K7MgJmtfJvNPcRdkjZecHm23FwDt
edJf13YP2PeiYh+nqnkeMKOGwiw3aKrRBtvr7PbmZZ3chbi7PCQbpXe84iG2XnzN
sVqfvx7mw+yfeLAM7V76cklGTvS7m6U2esSij1dUrG+qq1eiqHh2sUH/ywr9r9lg
801Lr5H+OwBKTvFElJf3IoxMRRM5Dsi5VEeRIeqWRxhFv308X45/tI+/JN+jzuAB
gVQ6Av+LGczZvNjPWNWFfBTgeRVTpHItixeKXJQBqYpBVZl51+iKnk3Mg07uSD+P
lF4VFDd9JzptkCK6x2tqaDD/piZmdydD9UPRdAjZGmsNiEJrSHkXjsp/WFEhvabL
m5uBp5KlREQ49fBRyouxqvYQ4BfIhj7ZF+UieVkPJFL/0GlpA2jF9G2Y7MXg1rzv
9ZPx4/eBsMPMa4gyZrEnTpb2IzJ1WkoX+yUfUasEshkiVFgH4qwX0wnb7i0YpfW/
FwsgrCTa3m055jS2aE6XBqVBDqItlfIYV1Z42HdTo9dAEbTQLoIAokLXvUq3M6RR
gfDpguUt2PwbeW3utq/rrLZIUOcuombWudBN+9jZY2I5Xgy+p6Z/Qt9Ubgmp2syh
tQXkvDql42u8y5lZU0tIbubIPVmd+7pRIkDegGtjs5bYBLVF/WZG5oNdrdWZXUc/
fziyQaBuLreHWCb0pa5qf9xuSBOXf86luB992sGe7R3G/AsyxO9hHMDMoWQYnwuw
IVcDCYMuD9ri8avNKXj7dc0nn98sApK+6MuWMORb7QvY9PYcSQ8CF0nkzu7TGI14
3/3J5o8x5nCMgLJEBRiWtjYuKcSUn4X7b2u3jJDIxzA0r+0ypsUa+rAmfmHpiBdK
cjVzGSCyk8JbVCfeGiU1Rd0Nvd+v26kW4YdBU55foagPPzWEsO3QIQAj76uTlu3p
zB3LHGzUPMK5ETRaBOFvZzZaGAw6iB9xVlpSpEHfzacBtU8CBnBeaEOtFXck2cew
W8W7msz579KK2tvZgOWp+VRG3xrX4FEwdd1djJtNV0lL/jbKjJB4AXTQSDKU2Xde
Y8ARZPtFFXtBKqpERerAsyPXqGXptf3Y3nv3I4hAGlvgPRQyEX8hMyvhu/lVpMVA
7VHY57rXtaLPSHgCrlMXUNEDLGqMgLpG9To8aLBXKfWJkpsCIXq1hqbspYOwS+Iy
CrLKy8eBgtCp9q5CuTJR6WdySJBdxbRzxuV/Uwr7pUlIWxE7hjdiy87JdRhwGXCJ
yV1EYhgDHzw2e3mg/b4Tu61HSuoNdJIfO17WNm+/JNrIf54uglNMKtM7dfGy1cHr
TKCAjQuP3IETrtA0jJov9LP9PuDdsWR/sFRtqmXhdNdRzWvf7BPg3GBleaYIOyR+
BiOdRSiKYigzb/ylpgu/NtHCo4Nd/PULHTO7vmnlu8uiZYEvIza51BdOULwvKe4L
mIHzM1eKYVn8vMjpNWGnHKoLO8dBoPapsDo9A1cjPeXbQSBB67LwGR46h2X8BrRn
hoIUnLrdxRW2khzZdsFxr6Je7rbtDfwK1fHmSETBzaX3mNKWe1sE+ZgOU3nOBuxF
O9WuaFAxliJIc9+0MFxkwY1FOhMyI2SdFCYHysjMJomIwGkUe/KC/l+wBU2cJsqL
bmLbYFUuBR+Js2sWV99D6chg6GjM1UDe/NIQL4Zf2PNH2Sk5xvM48VsyCYF1CZ3L
i3Ak9xkSyNASg9rY4ze2v3frmqK0Ws1610U5cdZKzfaTDdeNumILvLl0JlB/ulke
b3rfGsrhpvsi+LLblmN65oiDMFYxkwrKOR0DAyi9v7F5qgITnpAjJIZtjb653MMi
CzB4AE0BIUKb84fZWCkA+OCJqrxP0DtycY+6jB4s2FqJft2IiQxQcwQclIiUH9WJ
PAJ97yd35EAodNlh+f2SVHPNv9G4uDjwU8sV4STvCFuEA7id84/y33fut7pCinS/
KzOrEA4vUFk2fzRNFDffQCwBjcPczTqXZZHmHc8EUT1blHuYXtTMYT10u2cru4R1
eASyHXqwh/jOUHbURlVWUmbpr5gXgoR3+4d93U1Tw9xEo+4TyvBaso7ROSMczB3z
yzwyS0ckv2/L937eVuuuRtJqbyAqVNtnJrKmRQG31ZT+oDUUC8pyd0LRQ3tuEpMS
2RsdF/hRzjoPJbhprxjnbyikRh9nPPMuXqxXksPgd09UQpuSn08uKm/4ALrcMe4U
zyHoOahK2mxKcbpHwdnlqonKEQpjmVwJNAwrBqNNfiPJ1sz2nGkmMPDqQxIGM89c
EDPVOCDipUsU6D1LI36JfrrHald5ITGwJ9q9a8iuq+YA8DFJSyaFcz1HMGV9cyh4
yW+9RjY+E0nxr477/D8vpmlqQVV3gUuUJ8sZxm/9rQOFsMyMuSORtGwMYdRLItz5
6+iEuMBeIWx2hutMU9mwKq60l9+MVXYHzQRnGJ7+K/u+EAvCyGNlm9Ks82CZuwX4
yA2Yq/d7xqRIEUKzIesqeuFYJt3eiPbd1icf/kc5sf3A3rtPKVT8ejqw/mheQ+o/
4l1mhiiD7q76LgmjCISytWs+HyUd49wrMZy7ZMaWKAim+cdpxS2hqAMUHdW7VH4z
3muTtNYd277kfUzyYGPKpNDs7VTmAN4ijf5L8mXx7tNgsGBJsgUDKWEcDGrlW2vq
qj0e+QJ1Dmc1DDqqeMuKiMKO78oKTp7gdEKFNvAqNEOtviz/w7egV3905uKfd2yO
1bd9CqnmwPNZZxPGItJWuvcADcs849sidFgOimwTYDS46rjoRO5lbPxhwIUUsXoZ
4+BF5dFRSL8imlzf+JEAJ/rOHIvtksKIK+PzLZiYXTQZ1F85m8HvnZabsIMxzczw
Mq57zhrxXhkwdWAfm8KCsjFBXaRyKnHh1Uz2YEjsNZzg5Ro1bJoJGV8ghQR1FtOu
YYzRci2HzfAM+XUx5z43lH0EjbjU+4kwPGoGipdZ53a3ib+jnvjYulgLBz3OuxaD
mI6S8DbFwTWM0+QfTyKmtVlFa4zODe72txYE/WGbXEQvyyWSO5VODLpFPglm94Pl
7sG/1hLlXodqxGGWOQ1kI0o0RRwEWeypsSYJSOI/LZDA7fN6lpIuAPUwAA2Q/tCX
qW3r7yqKM6rZmMlMP1rzL8dPYto5NzdwLW4DAIDN+qTrMHtPPDRlN+HqxooMIwqU
vvGnesDfLKyqNLG7cXfYufndGp0TJ3CVDeCB5AiIgVT78K9Devs8hnjkRy24lJAB
/RpwNiI2UXoYMDQftG18n/tvjOeg+P5iEteeKdGoFCDKaAN2AXj9foPtR0xattvy
p5ZkURsl9AR+r+00YkXYsmaiL8aHyv6YS0DIysn7Ax5GBksWLAoqtDm7CCTZpque
h/mkuYTbSp0imw1SpnhHIjcs/Tft2wuaeK5zh0GFKTP+Yj5D4b7BLuNaCwC/6As2
DcWg348TOIaFZFIK/fIXKQfrNybMjkrtnwhQmYF0/B8UDAPKmi2Xsp2aCaXLCHdM
tA0UG1qTXjnGNVus+TE0a1itnKiwR3PSz2qlh/ncdmYeeMAeN7U5ipXZNVt2lOjR
Wa22tQoRFfdYuRqHr9mHzO0vV/HhpL6zv+4bgfmSnBlmj4/pdRyk0SCA018uMegv
rDtEIxd2LmwKRI5LwSEsoUlMxbWR3lVTm9cgtu8t7X39SOUKk730u0hhLeV7l0ca
yF/L/KI/f9JpG7dXXqNV9ZPm4sKCE9XcfSB3Fd0XP+khJ/JfxpEG7IFyrvKQb3ND
PZHvkmTQqgv+a68dDnKlNYUtbydxmESKbncyCyNXjk0Z3ddwIJaocRYNIZsMCafn
zb5CgUWqHeHI4rLg9RpEjDsz8eXXCzxkFCRscUiOZNTuJ+UgcDMzpn2h3H5lHfe4
0rH69ZxLnqE9wrWfeqjNUxQDmIfd5nwPp13N/ySFcMEXDtkHroN40sBrLlwLvxNz
SBJ1vmbk3ClOzOjaLXaVSKUjlsiHzDlJMntn7PtsyV+WnNOvJ5UmjezIzA7q2IOY
c3SGqZbTmJLpo1+pz4VtotUxH2jbit5aeTItvktBtBGV7ZtxCl/y2we9mmvOD3TC
XbouFmNacwKZiL7lb286y9dMesZosLCgmO9ViUytsjkQikzdemVwep5+1l0VOfsm
vYZ8hjRy/fa/Tr/czKzBNPzIODh8qzWRXI7Vcdo2HBAgFzjW18lEf60zutuWnxCN
wPHAwyMxTYmIBtWuqVqjkgVRsWPRN1qLhrq2Z9AaK9PI23rFBja7t43QBNveBizc
2pVXTkFIDI7vajhKeO9aLMxPg6cJbb4OhyZA/1OqbvyoVQXSOwfH3LeLX2/z5gcB
rnUq49JK6HrLDjKc/kN+W0C+wHZByYSUy5MvPX0+wAIBZWFQzQu4gBvYs6GHuQzW
kSHSeXCVIjeiLCujdSVnIUN60vUmle/p2eBygPrCzIyopMp2yIiHAny7LaWyT3Jp
peT0PDOa+3U2sGDd217hmpdJmiaPT0cOhw/bGiMuo7i5Qq96hnNJtY4CerBXfKx6
Mt//B84ywXSfAfHHoC5iKnxpFB2/kCq46ZsFBRieo3MuBKoFuqHJCwp9nJ99RPwU
ypVKgZi5nvMnfhmEJ72d2nPjPRLTGLgX4NPvX0nw1821Spzd/KRz8vx6uCnjDUqw
1AxLvnr1bC/ABpWt003xPxA6oR++zsfCn2BoKQnb0uPeRtYbwSuZMCjN/g7UaRg6
4RHXJBOagaXEKkWNBoqQEjSFgucQJ2GmqZPxLH0H+nWjMDdihD+5HnIFUiI/Ju4l
n0zt0G0PaiPgKwx9iudUMAUefrfXpZ5/amxaJspxBOaTo4kVQ7KyVTEV1nuEGvTJ
MdYCA8Ou9ck2Dnh3bSvUokb+zWApszISEm4IyyyVulG/RhHltBu8en/vR7TpRMK7
BrVLvDQadvZZc2srmptn1RW4ZpteRY5xaZBQ1M4dJmUzGTLZzQPbRwfsovvYLR+2
uhCbwCqk51Hack2fNSlxJygdoB0ewx9on4PVSdCtFRrlvtVLfWtbEIA9jXBB8PJD
r9ZkPBYrT6X/LcfLFOPm6B8QH4asnTHxDofbs+5+TaGvrbjEyhKNXxMCHew9D3Ym
/I/ct4zisvg7boRGLZiXQJ5FmuoZkiRJQEOluiH3jHn4Zx/SYlBFOKxPziPDY/xf
5VoovuZEeQEm13BdnoQXxzZV1I9F5gB6sATbMRJaS+bNfqYNNjdlA1OrM3TDSWGf
pnfRzsmSjklS3G9nc23jxGcO8Fayitczfk0roKGD6/40Be3238l01Bb/XUobEW0r
6fu87whrIDtmdcEynmXszqPnuR/5EqyAe/iN1Clx+lr1oHppI/QXP8mdHL0YlIvK
6b9bb1VGuvUy9+PAyW0Pz8XVVuNVTdxp44BBWxs3Xm3GTZ91HBLheCzc6W4rOHT6
pq6RtVy/ZXZfwOfqDh0ZjfJTQmub/mRemAlwTyJ0/c9wB5Yd7yUk809hOeSE4oOW
A/Fu7a34//qz3/CldFUdM2zwWnQGfn5N8bT7nAwnCQD1QdMiYAjxKIP/MEJgfX2/
PgPa0H5q+Rpc/hPu84BAEhMiVOeBOaKGzM/g5vX3FGlmrZRYU0WU6eoAHop10vkM
r4QssPlV7YXG6l1w0ejoPcsQTAa/Bwm2kDja9xqAg0UTcgccApHnnBf2WZTHaiSW
KbqgWZNKctQbd2Qj2qtub+Oojw72lFdAePQYsLhIuFeRKqyUMNMO3i5p3UfzABNl
bcbeIJeGvOhvdnxb5mjhUaA5sVJIWAjD6cQTsF/VUyGoKu6Khyj6EKxv8EANUO9O
cNYmogkswpJomyL0EOQIYEMSr6hO+7LpMYG97Ih5xPTsapIzv8xtsCr8sa/BztvA
qeIFoWneqoUcZg7lx+CUXfid2TSsyUcvECkxIiNUfUY1B8ePNGZptoT1QMzpek3n
QJuXb4/Q7rAoO2WxTAcqfYDPp+gl/tLB2BVDKdNMHWMrOUGSFjhvV2xHASYE6um/
Q0l27L4vIAV87rsosIjYWfUzYndC6wmOtElJF42lhVS31Lljk8LHWar5gL4iAXhg
gwcsaaxN9rqu54mcchx+DV4P/+ygQKrLIkfZr/EM17A8B5KDeVCVDiakQSkLFP3Z
K8KVUzBOh01asT0fbvPUqK/xWs15jf3w9haAVCSyqeTfJPh2Rgkog49dxjN4ya5m
CF1yQp3nPKHqT1pfCdRogLMqEfEzq+u8H0mczp8eKM2LfDPYjBQoWP6oCaoEEML6
8Ea9twGCA6zNGt7aBUB+Gjg8K/ySpVIUqHkJj7qdwoOX7mIRnucFpyggPccWwQcR
kMnT5y5FIIi3aVengLWZhMrIT56gzLlLs4W4TNduJUiy6Hqsi9sFtLRUzowUmqSA
CQ5LBMuSox4jOfutM1Z7bf8oOKcGnfXdVM2j3q1RmIyFqKRU4Mp2179nzOU1UmN6
eTV7v+OpZqzKO+eMDmjCGwPywmPfP5cdnS/s/BgHRDPNH+am+CERPvkTv+OrGU62
3pUcsytmHtEqOUYlp7xHcuV7XFiTEBEwcJ18LDe+pMGXai6FTSHrlPwqVsK/0qz6
aKusib5KQRx+DWnQmSpet3kcPfE1jnwWOj5jRivMpPpmCX9u0olin1wUdXo79SAw
glbOVbLoefyOOtdEvnRrdQdtCsgvX02dxkR8rxhORlf0BF5nVJ/+9EQ6ZP+Z1v2d
urGsMKECGqetCbtgAl/DRgQsk7jVTfJEEKQP5bxjDli9uzV0q7vZDoZboVQb4HZU
8uj85M0j8KJ4v8pibT9pplccVz46r8qkNdINFaU+BIw5lIvN2SG/RCDnhqNLJaNi
aB3k5KRiyrUMmhwhoZl4lqsv/FyBbe4q/MHcbHoZlVfnhfliU+/VUcJEMZuN7gTo
b/o8m0KFjpwLdccvAky1uMrm2eEbS1jfE/SRInpzcAug+UvkxUzFrlR5QGe6brds
vKh8WJ4rspcZWddnzu57y0EvPUEphexpF5r0BN5nvFblFF3HeXnPwiZY/T0noLnd
yymBrvHvDXVRx73gYmh5cYXkLN3WEBCTlTyy0ZJLI+ldQQj9Ykur5CIpYvTjFUUq
JNCIq7z8zzOcQVyJSMTIDkXRVh7cTHA9UIw8nmi5NuT4MQo1c9R+tVVDtKN0+UoU
Io7mUzCwfs7dokuMggunSAhzGjf42o5YKc7YGMWTBLR4ZOicPe526kaSBaWtD69D
CBPGNKoT987XsIdYE7WI9VFoe/nbhA5VQcd3I9Ryw53kBQwunJYFpBDYYzJQdnZQ
3/eEtLzp0t0WJ56sA+utBPZXvTL1ESGIfGlKWPjT2v2iOmQ7yGT/PObN3MerWiIN
SF3q8bg6dJLjxHzLtaHNqfh7Vn/ipnn7Hc0QqNQ5q963IFDDHCKiaGPmRmDnl0UX
h0n1n/suTIYuZpe+K5X3lBXsqcA668Pli+cdkdb7AvEknQp/yqQLVHJ9A+ievZqS
6XlrtK/rWG2ps/X4tyXGwGtZUWLoj5Q1V1kTifTUztGoZywdirbbdDRxk6DBe5cb
o3F1ESYQ7W8vzUqEK6RKtbbhKouu/MsfWt0sNuwpS+jxQOurf2orn/kvMGA77/O+
T8s1kOK/m4NlArs6lyZqz38FHxVpHWbSDxMqv3B1omj1WgcAwgzbXEfIaUTnXFYU
7/OS0ux2kikOZ51vh8/yh9RqecJDIyyd8nKvhpxmY2VFIh1UoswQovz3nxoPs4fL
vFAwYjq14PX3VFis9zpt7/lWysZ/mES/sPlX/lw7HA144l3LqMmmr2zPTHZOJw+J
9B4vx3Hk3jPlRdwJxXPlN3wMp/eWGocU/wI2XzQeLJ2910CLVFYcHY6IuIIezguT
lvepecN90gdDt9Zb1hgIgouwu3HFfzX3YhM5SbFDXL9SAMtUSS27cRzM0sVUGzYg
3ap/7O6nMXR80B96tr1fzpkEgjy14r5qZiYpUkhyujB8pGIQL5P+mNUvtH5XSVjv
TgqCegYlWruU+MZWA/sogeU/JKpA0hN8+fun317RAAuOZLbWOVm8bO55jcwnrS00
YJPK2+bjF8exHNwFkUywvWzLMLkQ+feWmmtBmx3eMXkzqIAOtbHo31ZFzwfwItXc
dywOn9kVVAHrblb2g15qMbTYPbGuvrkShluiGcyLkPM+IU5B5bNQkij/DQk2aeD4
AYNeeRmahT2g8CkxMioY4JIKBQ1A8hvFCRbme34BvjI3tbpHUOOR7YNd2FEY8YNf
gbrcAwRGYEGGkaZzoaWHxelF8zAQhd6z2qr9ZUryTLEE0lpkfoVolr6+xncQvzAt
QY7pIhB/JQnhhyfF/qMox1S0DfaATeevMer4TlXtBlM7z5TImM0jGnU0rygI8fmr
mRAXaLXZSQk2BCDfTzVdHldOgUNq/megzHAfp+N4PteVI1c0eh4+w0GiFL0rziX0
84LkFkcZ1nqa1iKCxwvLUhSG4FuGsBkNFX5GHSmJlPcYYXNblkNdrEwLcdn0MQJh
uRCy4UBHEAgcCPENVBkWCUVH2xBTeTiR8F6zEJKIVXB7V8ZE68ODZsZhWGmhX7q5
QNV2VleN6PUbuE9XVVTfXAem+Ch5LfWp6L1p6hoRow8Li7hOszWimdQIfP6x95N5
08sT1YStBDYtoiS8fs0FniYOdULW9WOHQ14RlvlhSFKsWqaxcOd/4WYaRrq7pY9k
BDuWPCotDgydPzTP/Z32wlqfleeTSfb5I+kZNsi4jqrKPVCBordWdEaKEJNm70Pn
UftdvyvmE6sIoinezj8C4KGTOJJcX/ry3o5CO6RWI5VVDIYqsTglPtRE/u/8RRc6
Ppf1PkfYzP4sPm3I9H9Rl1nZBdWCwVuam0yYNRUs5BUcQ2uC5Wzy9pBGmHClFWy0
ePVFleKYhX9eZ1lNyvdXqUxfE/jA8fI7237WcmqnewMqMBejh2hZjm9zqdPo0qcR
MxHNU8PUOD4f4tTGJEYymyKxuREjphQxrrAmzzLpypdXca7Epqxbifcz/Posj5YE
+dyU/lScoI3IazOLgfVmMrgvJK7Iwkoe56q2gY5Ne8oDZgbfsMrcz9jeZbX6k/Se
7uwHDD1pA00Nmox8lwT2BFfCz5y/xfXmGuux7ERgHVJNmVvRGAy8//hexYnEsqgn
5RkOhXAHATsp5evPpagDLk7xjUdNFvROy4OdMr2bjvq4HhigzFhKhI1pzpP6rwRQ
XvZnAsHHhLGViBOecnt2cC/8ZPSnvXZJ1OgxjGzHH/oAZGnIO908H1CPN014wFwz
hwtwJCAbE3BeQZvuQr6k9Ta3gBNHwUwxSu4TCdfE23pFIplFxzbBG88irMC8CxJ6
vzTHPjNLBliCM60J3VFflps84koln3o9QnTWRCoC+ZYDZgq9OM/TAO0gJz60k+UO
gv6xhZHgvjAeVK9Fp23Kv6+nxX2zKqFGyxoB8VsBz2KAQX/nuBs5Tsw2M8gQnt8M
uAYTaaZc5KRv89TRbn1MqkyXMwn9wSFHZyekH4DyvyUvzOiX7dukFEZT2tOeoVIu
Eaz7QP5xts8lWqT3hvkrXczID/s1YhXX9L1hK6/4gazIHzwcCqBTSMoGub37YOKw
9Mo5tfCF7K/1mM7tRgB7cBuusIqCU1M2tgSKnv0PzFx8O7Wanuv44l62x87R1JQY
OQdiFIuTfYffAFkZlEPshLepZTN1VTScbcT8SLdXJAUoE4laa9igqjzX0+KtkDNm
ZD8pgwIIJSNxb0/x4IMMSiY+U2XlLc7sc9ZwLmWHdwPtCENXcIOSEeGFaJEnzN8N
HQhe+JkQluvV+MFysbRBYS/9suVi3U3BjzkslT2jUeNYLNaennKDsget1zzdWRXr
/Dzq6FUinq9omsxcfF/DSeqqyMmyAT7GVCn/4BH5DQpd9gHGvD/gxRBP2HbggKwg
yqGXPfBuV84nmGBwYfsG8hLMe7Y5yVrpSIhBkqzAWagJzmqQe4QkTDdePrZap6D0
6H8DsU19SCWkfrSIwuUxbtX1pVPV92lfzdxx+xBANdDJZGzFwmb2NnsgSS1QR19p
EatmOX7zv/6PC61ahokFP2Y8eKlTTrcUIjmQp714jUG1n7Eb4P7zx3sGyDpVs4Sf
KGV5WE6Pv6idkafK9eOln1RSmOUzNjDQXAdRsJuZGScELuLhmcU19AC+Jvg8vXPo
ju3n6T4JfHwfM/TinoeBAbIwzU3NVtKoKv7D8nl2Ttx369OUJfqNSI3jr8tyeotq
ZyPSPLEV/Q+1HaMPlR2zP072CZxJuXBka/V+jkQ5QQXWQ//YH1YX9Ru2yXVb8rPQ
wUA+ctd4DkIrTNmVITGQ1nARhJw0SNX+uKOM/1+t+uzkaFyoyFIOKMnE2v6w8Iry
kceji4NkLVvrAWbCf/XTuOxSpDyhOhlCsGd7FC+Tj3u29I0uRc9bQ5w8+W2/O/Xc
lXkw1aX/70EhaHKECca/vY5YTpjQsqADtwC/qxDn6CYqNuBwqjMDSJeqMoOHXOTA
bIdkhn4lJy0URjMXqk78RHfS0W2fZU+F27pw4gylfWkzOVxtroP3r1PCyuIDFCce
Nl6too3n84qV3DtknvmqwSRoCQGQnpFPd6Gp4AUAG+yEFMtqdhKIto8BvWVInH/r
gBkz3bf5zxZjqOZQi7WQLNoErvrAJh228u8BmMCCfwtwsuaT8FyVydlaGKhMbqFw
b2pvN3iX26YmlyW0H5kqc5s4sxokF07qvHosVe7AHUQrh23NeZzzh1JN3KrL6lLr
zy4fE4r1cZjqMEl18+Cglrl3nT9aWdAwt+FVeuIEQ+sz4ydkzozYq584le53daoj
tgzNq5szUkcNVZb4k5jNk5OgVMwaxGCgeqANxyT6gBtZ9xqcLVEH5gDiqsPMk+TR
2szw/V6xvLYwll0mWJM+SmjMYTDPX2pkwvQA0BUF/BlttHfcZozwSJ90n7tgV0d4
1+O463aIA9sjY4zaFHhCFngRs2kyput1zjqZD5/hgoGNBbRymMm7YVK5Sx4CeNin
tSlroeK66ou9Z3ctdw6IX7RfpYZf0esiNbCHsDe78+PSq1PuVoRIv5PE2wxGPois
QHEaNBxk4LxA3wgFGu6ao5500RuQjovBlGdYR5Fi0KLsux0xDoPFq5VENvFEI6qt
QSoGrtyKRRMzLFgzCOAE54uAL2FadV7o0+yb95Q7BEYkHLcF1JBrvoZyqBYueuL/
Bw1cIg/FWN6r2aIr0D0CahWNpnhFCewDvoA3QsssqC+99yi8buPO+xbiSw07tI3I
NHoFq4vsx5Bv0SWsjDiMKvKJ2bWZXrpJaE7hKZF8ZMSQY9F1pVtU+Hy8QDM32gh5
52QLbma2UUhmE1OkhIB85CdkloxiMYMu8Qrcoub/LL864SogY83GLb9Hp6nRlcgK
IW8rIjA1+XiO5HSi8pOiHKk0io3squEPjcyEX4m7+illnHH1QHvDFI7pTFawrP/9
bSiv0h7rwWf6OvwqlUs7tqeGZNaz1ycZlTOwy59i1PQ7MEYK411Uitg5zsiybklW
apG3HM4KlnKZR+evSniF2iHKdy+Fi5hqAESzVZXXpg2LhDpBqtkVufLEt1srFeo9
nrD9I/jkJwK2YAAPOTuUkoNWWSP52EF5CThvfjQqI2Tvjn0kscar6VeJGbS4rg4y
VeJuVUj2HGMZbfEfaHUGpWVfefXLDfJqD1S4aqFxAVLC1drVTrjpgsKpOjGpUub6
sWHXVSgWyAlmZg7L+DY6potpkVwtOtak8Mk96r2Le8d8D7d0NBJ2QJKz44G8h3qV
b4vtFCevCPvtaDRcJIIO6TeBkT5w2tZ+XSNs4O7HGfD2dMZzdwSchXclqx9ylqlf
I8bVbYc1nXhJUFpjnIOzHq4fMh8xWwPM5IU3whONfvISL2B8UOGKLxMfsS9SG9i/
w/lgQ4cE7CPhH3RGmXJh0WJsLkYB47MUyi/a6b074vjwWzMOa/JztZsgtdgiK8cd
9aENv6g6jOaBjHqhFtkOGe99a5VxtEQ7mJGBQ8aRZavJFDk933nFpruhj6OgJYHA
uuPMKTvfnMU96kPrFRryNwcPKabBNAIefDiLzzcJBfHRV2aL3xVRMvpq2CfJdFMG
H5EcXgr1poBQ9gpHcrHaYberPyCPIOFFZOkAbyA/3j8jHKMUVB4ZO9buTbIlHVn1
MlSB1UOUc/5a2fRi4k6Dw/qUgPrY7+RxtT5ncBP10wwiqlsm2t8u81rQVHRiW9xw
IfDIkGh1/JqkrN31yMPxMquUdkqSI7oa+j3yxyE7m0LhFb7pndJ34MShBtAe2FuU
xuAwhZFgQhASSilKsb4LL9I6Ig+g04dt3gJNnXDnqMfLk+BNJ3d3sMGUnj6AYDne
erp27VeChL5X4BfCwprlBL2mn5DO1A1AC2lpgtZt1tDVxNoQS5msJ7wKc7ofXXu6
UTmf2EZtKW8CNPaOBLW6C6gFYEcBUxToGeIsjvG3PZavaANVPOYJVtqMHbrFXKss
l2rLGylX6k7NcNM6xC4ak/zO++6nOn0nv6QI2hhNjCag8u7H4p9VMzlq3rmcy80X
EzkgtVB/m3C2iC60VFs85F9iNG5qXW9L/jiwUw//FFq6c0rkrIlYt0yRPagnox9+
FJImwoYBz8xEhMHOhQcwkN3qK6hW7jlfF2LUMGMU8rNTMOAv40K5DelTR4bX51j8
QtmUwkTMUR4RKUS5Scbn7DvQ64Qnb5sq2iqMins5k0OJ4FEhYkv392bEu6TKuMGk
WdI7TUz9XCtHLkmGo+q3G5MZSWqJqQ1B5vBw+5j2xa24EvrfbjCwnBw0esEYuGDA
gWBPpps5R4M3qABjkR0TNOW+R3EWjlbawuTflyv0HMyBLN8scn61Gqi+N1gmiCmw
qnQwC01nLuJurw8Pwax6vCY7zR0rrQHzMpaSEhgUmNIqwWyvJOUXqGcG2Fwsa6pH
YGtyaE3t5nIvpO3qm32VpkVBqfyhVpUy92ShSODqMJY+74gHawQ56SMXRkrWoubz
dYibwYd4xSd1RJvBiwTH0Q/cjli1rK4sw6O4+0GeKEom2gIkgyFvIGjTxs9DzzQ/
BCBCd03JA/1zzN77PQyYhWJE8xp/LzyQkNcA1yNA5uWUygZtRSrKMnz7Icpq0ud5
/mt63ffRKyBbWd/Ui2nZl2l/8L00ctuvj753+vT4mfKPe/3AUoVUV+FPVE4/NU1H
DPSLu7/KxiEYNwxdgz8w3ej95z5MUaweZ51XM15w1OsTQQ0iLmzOBJifZbBCoh/z
b1ltRN67kDuuCZIN1IoJPUnk8og+bxURuBQLrHOG3jr24/3+aFSgB8oFDlarcoDk
K8J5prjSE7YxXd9ZnD0lR81VrC+C8LnoSmMy0EeituUbhQ/yEBp+xLJjXIUtzP80
2Ahx60PcsnpFH/quuqmwWYPRbY2JvU576lSBK3Nx/mm3FAEnZh/C5S2MyS0tdyBd
oXrrkF3aQlrrGspk903nFcv6pL8O2C4TTSHrL8A4jyUfIyiUgCvaK0EE/Wu9rJ3P
GM0sMeIjc0Csl36Ebk7myic8eci5sD/v2UBPShZaiSteTwWcoQTVJboZ724cysvk
DNcdZyysWg+tOPtyHxSKroseBRxafxYjcE5YxfLV6vG13KK0u5nn3HY2gLetHxqi
PAkYLe+D+/BW6U5r0tmaZ6hOVX9KbPolPr0SQ/rUnysIX5gZYDp4KcokqidupLJf
Qn0yciFsz9HZglrDEcEs8wjRcG0piRWROjynA3bm7x7z7oGyLRvCjyBDgab6YUD6
1bcdhsVKTpr+kPJl8Br3oDqdKFT1pygQI1X/ni5QDAX7AX1GnCKo7fCYgweetPop
GNStsbaPtADpJrfn/2S/kZF7n46Y+c7er3nxcsUYrfSlcP7q7eEkO/Xno3LWpW/M
/YymE86srylAzQ7eY+OBk4A0sbAlG9kxW1WcIMsuYL0/75UaCBD9VCeECkMNX6D9
DadD470jOal/7VZCQG7VIvnFLbRZ02ZU+dbOPABSp6DQRZWqtOM+lvGQnbN712q3
7uEN9dkjaJbBstB7iZWRo0ZNq17rSh2NUk0S0NqUldByrlSCeto8n7dXW7AwuDaw
jgHlFcpcQ6Bgx/h/XHQTU8WdqMr6LSxFr6GqYFIXvhvdfGUc99l6FmxaduD4ySOy
dowPdjv3nrHtEaCohZtSpw3UCj3poYZ/1uqFet0mJQwDfVXuJ0Ba1GbzbZS3j8uB
mew0MY6Et0aacma3V3IcL4XfdwEiw1JRkuHVUXIPk1cU5KgtvOEjNNJ3/pJ2bTTa
rrpHWMVH4vXO6x7SM/b5XsP0jXgatCtCJGCY30sASDezlZMezSu4WJvJVhf3EG2N
LNqifhaoX9VQfyzsWgpOfYJI/plgWLZYDEwtkA8A+PWwdX52AnTDz0Q+tlK/32US
ZuLw6Z8yL9W6Wj8FSl37v66Nz78ttjGHVK9uni+FJTshn/AeIJNbkHDv+QB/ycXK
24g+UIlFFrXpGGuNr0aUxs8pj+e81INNF0fXj5kCyY4oZnGNViTQ1bTpho63yUlE
BpyY0Eg/XzYiSjl/BcdEcoHmk9aJG9OvKN2mk4KU2eAqaYZu+4qVIvMVbRDXgOyz
c/NzmBqf7uk600t+qZbmAEqarlIghu8f/0ZzX5TWW1cE7JJ6yL48Ml8u3X8UKmnZ
n+yAPcKS0BkUir9+BRp9E7Jvxszi6edijSBy8kj253MwG2AWnb8EM4Lni1sWP/Mc
WywDgqSNbs1ApqcLdxaR59Kcy0UoFdnaUlUuO00pVOn4ndgWfNTRPy6JZ3/VXGMB
gHawlkUT9LELteYEWt5lKeMwJLRsY3azo2l/VGTlQ8yb1CCUjaT1VgnPO7GjYjFu
cKrN4NTaFYhsM66p08Hkeh+wWqoRDpsXiJxQG3OuYB1iIY7qojxDzPydByFFVj7l
DUboNjjcZg9ok5f7S9UdOsVOHuuImmiCd3EIe68We4jgQomkkW7ylsSgTnuQGXaF
jTLTw1/uOKDfS/O+Wu1PL+XA6d25DgGaQJTKgJxwcaVfCqhz+gUEEA8Tz8e6oa08
OyX6rK0DU1OrQF9j7EBOt+EIMj9l+lvP5SfaXYp2CBwuZaK5C2srtnitBXXYGQdx
TfwZoy5Mqp0D4Q/qS9bbqjFXaiPX/ataS+7ywrTmx/d2Arei3q8xwv4RFEoq3wXc
u/Ki1I7dJZmFdJ7O8Dvax7iOEimkKpNiavnGA8J2A2+Ztd4m1KqijSMCxjW65Of1
ES3VxQUzFibBg0JrZXaovWU5CTUEBAlkU5M4EoD2YYepHPXFcWYpdDy22crdhLCd
kHL3oqZgy2Y5J6mSCJSaAqhJIlTPIaDs2a6oFIShShnRilaeqN3iWTZ+g6JFiCcv
vTCzjz7rPDCVIvpkkzjwBXbXIFOiQ306buZZBlQtImKvYj+T3K6NzXU5k25yRfwQ
tBxzdI3EI4IRKn7w2gdmjnzM72h2WfIpOWu8N0YJXIWGii3o4dbaqLrQWJiv27pK
i953PdJPuFq65+ceJ54pQFo4d5tLv+QRCZbtyZVAH8ApU5LHE0wGtNcBrV9ogZ19
fQpGNd1I24WftBFN0td+T7gzWSDk1ZQkqQ8IKUzNGjdmRoIkOQakJ0t+TqOjNw2t
hJ7ifCwPGN26+SRFOytCxMVOi0+mlIDKnjO5WpD8pq1OImT9ZnV7j6QZZO6QJfcx
+dgJ+JSC6UKe/rDR+8aXLMz8Qf4cXznh9PhP5/tszBo++tM0Uvq49LCxakznIvXy
YYfQRmEKVMVnFDGIPADQeNyobfupfYsiZVjoWm2JvFi1MbPJaoa7+Xn9nwvde624
/unfXaAG2hjAw5WgqvhMnUj7KuiJVDUo1uE83OJ0NnmaM0k3xlhyw6KwZh60yYQY
bX1T244rw9YuAY0UVlgpSqNwih3f5S4SKLcq1DJx+NUOQ1XQWKYX4jcciCQTaZ6Z
xfXOs2x0rIY1h/RcCmhw8SPv34FUWXg7hdw4vlxVym745OV6cNuUCnFLcHBsibl4
BF0DKfRSILLWQv3RFz5XrS4+X1n+8dKkhZcSGd4kanZ+LwxAG8F5NytHBDDy1tbL
mukxqDcEW7VLgVe0PuAF3MgBm2QWqS/iekOpF08eLxdxuGDqaYeLpMqXp0WoqsZB
9/uNbuXGMAV0g3dFp/Su+TwfjpwPw75+Njyka4jKFOKTVYlfdnr3bNuYMB4BYmGE
KOwsXe8HkczMs6noxRov/cU69/FgYOglFG33nGY/Sk7QJpYitFegtrIWKTVEk9Rv
Hcxea5HXRT39XZLR9SG1fPjYYC4uSCkJwv7Hdys1dCwbzdsWPLaTPJEsxJd+O1G6
k9sz3MJPGFBrqujeT/jRzO9AyQ1lT13oyfTxKzT4wDXm9zW6+EsRZmqlvFn08kIL
1nsyyPV0prG+IrCPMXgtfKhXrVZ17KGyQlbLSjvU0tpDPs7ONL2R2d22/A9H7j4z
WzzBpOg3zwpBL9Qf7kcYMD1K5xA3TiqKN90jH1gHhb+d3vN4yqqoFJdFKdFNHnm4
a1EfdLeexpeUfrLC2/fkaPUNcJlHZIXDK3eY7NLvMwytOgOUoxpOT1CJe9kWmqte
cxPNoPqQoojGbMgQGzUEu4AVVC2GVVbyeKvJqpdx03x439NuMOztAii2AxNaDSK7
mFtnxr/fh64qxjK7RDUkhYdlzuXR+7nRjdoE4OwEpBrgUmys4lvB6YJ8PxuXTutJ
XUHtT3xYVY0M5N+B2JkpAnOpyKx0PdJgdngKMHVolcZoBspO5dvwpcNoTYtDomkT
SOJ7iWeEImQgC9PwXPCIl8+oxtDTVflaBv/+ivxhnrxR/jCD1Gz9HPuRQBX62Syw
7SiIH8uWvE8MtFie0DfEYG60X+KqyG9/cMPkxqgt3ynQXylBll4P4cGVuybTZUJi
VEFUGWUAMm1GfwBsyYat52dEJRFNzxtVfltfY8W0s5ETDiLBxy0pc5ahlxfG8Apq
3rn7Axe/vGFoxiZDkK9FhM489yUohj5iE7WaFpO0KdwlFTSlWEOuwnjmpM7C6NHn
cLMat3CeBVb2jtgQsaOy3tV1DilJwyhMufrjKUuULS4qC88oUSuvwc+OyrS/VEWg
um1jdG3bNFnqxIV+XeIezxgEDK0iCtDrc1N9veVVskDSRvxtgCS6KfBv38dUgsTd
vTgfxbeTM+b2Ar83Tj/A7uwVbxiN6OzD+cHw9J8nz47JU4vv68GpmCH5sWtwLY4k
+uOFHqfJL8W6S/6uc0o1E+4LF/Ut/nzsGu5pE7P0zFZoJkNpBIcH/4xS3k2st7kf
7xYs1l9s2ZIKSws1E9UyNd+mZ9UcquROrw7ZKQiOJo+x6a8KBl4fpuqRPKB/uL58
gX6Yzk2ykwGM+mWY7rFB/dpKxBqepWQDar/EcznfjozggJpCs74tSOSCYeXrp2/T
O/T2DDIoGwFu7KLi7F95y6e+IPXJdDisPM/blw23hAOvtbRBS5/HBDq6fSXNqERq
vB3aXi5pxIAitRqQv7TUk81obZAu9yBm8O5PziHhviCcAdlR/6t9xZ+WB1GdV0xO
nUCcL7BsZPzHNFgNOLKY7NMWbeCUNWPo85LHuwJmDGT2d5eN4yEnpC4y4Fy/jUr0
vyuYBcXke2VaOrv548eqyVx5Avi8Z+1W9NVcUDc2kjvTgyv5YUD+G1y20YKrMwba
ND+YKbn4OeL5CrXcOPuQORpm94GcZEA/cS7Ju4h6PyGIPoI7FY+5qaujT4QjJpN1
q3XuY8ZYGjev8Sc8rQRJluTBX1NydhIBPGUM8DR2g3a3K4Y+VtjZhBiyiP9Z/pc8
6lOF5UpRVhtta36Z9m3xzMFA1eKZVjyM9NzaIropSL0xiC0SePK4p4MmHATMWa1+
hzxft6K4k+Lnju31XMP7z4pHVQ1gSMhRkjmmANjZ+ugSnoSUVl1NmvmTtDQmqKVv
M/Z1zUoAjer47SehSpYJ9WS0g0d/5/U/fgTEf50ipSC+SsoR9Lt4J4HXb8vMC0do
E4qtRfJGaJe8uL+nvCF/M38jGUNFecUhdz+IHHzlRqNizisRFYqfJWre45vRODkS
SikZwBEq6UQhZ5dcuf1YRUInLG0TGfM1+esYOtvDX4XTYoZuoetI/A8yElRSLyD2
SNKM7lSApLtc+lWd7X+Nkaq83oYNHUpRJkFOSRnX6krBv0Kx4yCf3ZQgnWqzf2i8
c5gYOLzwuX09qm5NTZ9WuELFYCe2SpS7+PYpCNv38BcWlEjXPA7Ta6fUhc/aSX27
tzj7L9YMkA25cnvvsv1UyMwslWxpKvrBmnd7qm5r+c2vByTczBM9//W49EQ/auD9
KmZzEKyAAnpicukjMoa91E5UvOh5ihmsCIFS5GrS7M1nS2H0kozwnu73hDoQKWQ8
Rh+DPrjhwgZMhlN0wV/vjm00bJyeFEHngSxrrhdf9W5PcgJQ9TLstQ4HVs8rUMfJ
KUSm/1G0jAP4EETqAsAa2ORWUeWEo+vZ+USEa+ojRT8WvfVcINqwhLt+Mw45K7DZ
YXD2LvuAlZzV/tpw8tXAgWm6bZL82dx5MHfyg05n+jtAXHx9T4OXWKsKYOFopFpY
3/Y8GCToMpa3LYWTvfHa98CPvrFa2ba7njUYDfpHqrWRpSEcrzoRS3PPGjQl3fZT
ywyBn+zvwdSVHh0Om/pc1pk/x/Ylj0dYWOergr20+kI748WCEYdneKYutgMCBrUr
iaLoAYBCuylswxCcD54tle+xHoacYif74bz+v6qWa0QYJWa3y4dOgL/3ZK1q47Mk
jUF6Nvw67ihoxKwVd+nmQDRuZS1avgXaFVh3PU6gvF7OMS+NdY5cjXdk4RsJ1P5G
JkXaRvGynSfmZkFXzHzSbeRxBzjIVhnN7xDuTbDztRqcH258cbUATvckN87kIavo
JKPZlC5Bv4/g/CWet84kiDo4VOS6aC+yB/RlH9dYjnlarY3RRWrsaCK5bNHhQR3X
90eyZY7WMhrrPKDu0NgDL2aBghV1Aigz/FF+GCXADY4MEl8wyKVOhv/3YnqloeRn
eIxEjpYNZwrU3i7Qi4WWQtajN4dqyjEIRW+w9/L0NuL7mE0cLYcg7UxRRJfb7IAJ
hmL3r0T5qQh+XazQZ1cETXNp71CaY4+dtyq6/scaUD94pjaHQoGufkJ5OLln495K
KgfO8GPEM8zByDBlOC89K5xGYmyfd3wAHNTpYtFVXYo9c//ckubtEP9kF85XojUb
R8BP2/QZVHbznAkd4pZibN/jwjUNfkFk8Kh33kK2vs3/5kg/EMxbyzWVHwrgR99R
fUrgutwrNPKvy4S9gYSO+AWVO9iSL2LZr1Q0bTEcJ5eVpPwduR3mg5O0bBxpfsEP
wTU+1pec1hgZdvsQfKseX8pe4MNRCPSIPTl9J9CTHeFRBj5O6cVTP+boqQkqLptT
n+soSDpqzQmttk6qqP9AAN9nwcPJSBb78t7L65mD7BOH3ZGFsH94PzkfezZVfxfo
SmwhImPtAicc3BG/tMAwlO1E6ely6vssxjnmwj2gvzY44igit5iIyu03YAJgw1ro
u4yz5tihn/LF9Rm0KKRx0dulTCsOvNnhcaJdLvKk0bGSFyktMzSghHbByCdvT5Zj
Q/iLeBRqZRm4lSyum4NB+sRdQgmtEYFSEYll/MLvBuQso4G/piZ4RCpR/+Or2dvT
8q0llkKILjR13Xil/+07Vixy3RMeZrBJxgF8AVZExdd+G2YY2xLPMU7hDXBAtfAx
QZlH8dJ2B8SNkOaCrn9NIAcBEzNTAUqKwox5vpmXF/VdGWFIrwhl8Ft0O8xKVHW8
bjvQ2khKX9g1EaDKoiQBJPtIHEVmWbDzMVDUtrTfaXQLMvZFGZo17Ne7E04gfRub
iqqH0DTIoZ4NIFgDpBtioVEVtoJ0WEw29Z3p7m3DBSv3Zz96g1wYm8P/cg8/Gipb
CJrhL3BBGbKbTGKyM/tmuqq5Me/Xj/o2nxqYguLAdePcZtlMIkbYlsMD5IZW8RqR
YKJSTrPwI4lsDW3LF3zMzQ3dY0TQQbbUNtrk6nWbzkeSsp6PRAvNZYiXqd1H2GyZ
AFrOPrgaXBaupAbgseF1uepwek9LIRbTlHD/ofJQ+IBA6cSIiBYi0xtBjTo0oWVu
ILoYKlQDmKyRriHtNd5ezwb3TmH8JbFpdn9zlDp8k+Rvao+l7GVRTldKXXnf/2xd
GO4K/ozMdotrTn9vyqQOxkoD3tgKS9UvgIopSBSG6TPyi3U9Czf7u70pgKux/OuQ
BC7XD4MN08PRdPphImv5FFkh/WOxbLI5vqj3LoVium4F/nhv6vHod0Fsmb5sM1on
XdsZwSNxGZ9CeLBvRpz1KoyZ9f1iikewwInJYGMLU7qSa3pWQuTILkQiBTgBrSek
JoSR9ksR4bG8qNYz+u5+JFJF5hI3R+8kyUEmOSl7rEVknW1/EiScvpTWUQCDjL+r
mjC1LbeoCkk9zNNVCCsHtteF/SPr2sQptYH5h1mEjKg0NG7njGo79DMSmfSgDdNE
uGOJc4habLSH2tyZdkm19d3tMx+6S/SPX6gf50F+oMBWbe2xRmc+SOJ0qQSVI+JZ
v6t+ySo8N9L33gyXBmLKT5vZXHfS0xQdRGwtd3VBxG5S09hb9NbnlnTYVK+5dsHy
ReUcYZQGpLOFsddNT4NNPpH7rzr7JEsQYMfB4Dghgk6YIFWlxOVF3fDzk8LCVs5e
H4Q4zilzydbJMPAfRYMPuHprBOSwR2OnYZGip0HwOs536KFQIL0xXt7T6FSkfXn1
BhaXsgtSY48rqximXIQZTnaQVNrITrdwVZ5vRRt6CJEVBTjAGcAb8mbAGt0LRtfo
/mAnQblUZ5FJedFYO6MXVvcsD6tb6LYiVuQH7dBge8VXuzhNH4ECOyXrFXadBJG4
Zx386yDe0OW2g0YYZmyV5/+NU3m4BZv7VUMMnq/D1d4D8Eupt3v7P44PfszC7lHh
kzfQuCZYt3kOCzgvF/4gbMSXhhQmeEBmOilQsY2lfWYc56GuAZ+3Rbz+rUmCPdjZ
1qVyTkGhH7tYdWMlPq03E53Nm+RIu29TiU3KChcEY4g0eYqJ623G/jQ/5ZYzLHWL
iBtB4alFzak5vDLuiOlbXDe/6YichYvwqDJThKp+QToEJ8U5OyhVIwwIUIOZBJtN
QieBZtUlM2s7buyymhJ/yY4pek5AKAxA3jdduRbrbaXzTB2ZnapEViUvVupRLWRP
taOubi1+edqdrfFXALUE+ox20oVLUM+9VOY/MqU0faoXgoQ/KKaRcWTfCFabAdrJ
L/zYMI4reUF+FxFx6SIuWEM2kMu6P7063szB5oR2llMEW1m3vtJnH1eSPU9y2L7q
2j0eh5v9dYSTc6/iuKgzhwf/5OaRGCLyFhk9/YN9o0DypPdYaQh8wiklUHRoW0hd
qgZFsYQylZ9pnrTCqVYlIlCVHGYYnDZCNyV3ZfPDbc9+ZiRpiL1EVTKR+UMoHOH4
lGuJ4UQJFXFQ4HSqK+SLTQQZVBNSBkTfmn/csqG5vGmfGo6pIO5qPEd1qN1wJqLE
VHEE/A1WmAiW5Bm1Kt59oJWsbb1E84aYkPEC7T7ppRWYMyEn+kb56u4tMLxmHo8K
Ep05JYJw83tDJ1HWdw6J5gxm5ckx6wypur6dYrvq/z3i+DlrGcRbQx0HIsPT8mnJ
SDu9Nry921BXXLRsfqqV+LRFgZl7eXQX7gs2G7wJ0f3RqYIJ4O3ZS4M+gqL0jtrz
pEyfecPpxmQ2NnZGJEoPIi+gz3gJ6FStoJpK3c1iw6ZlglBzP4ziFt9FU62pug08
EZP1obkM43hpIAUQc0Lpe3Tcy36BMxWAilsMgzqB46xFm6niQhFsrVBBWMdZhp5v
L9VKJoT1NAmSsp6D+iDWi/aVAcBHpKMzOTj2+8Rnh2WmeJBf1KfsUcoR7pQAHNp9
2uOYeuW6QbDhlz49PBPgkBvDnSM2OFWZrWgcQEQQEk/0NJKYCH2giYqw5toTnRKB
ZApeUXYIDU5ZDUN1VLdri/s8+wiUQZQ5QAZG/NDD40qF4RHOod4mWeUzf82qqMJs
llLghmhqYs4YurxFMKJdlPJk0/ro91R0adiTHxt0M3BdYZyWRKEg68MSnGkinQ1V
E0inqtWA7uCazYMgVKGh4K5TuIwcAGr3IEnkjYdy43/e0bJkx53hZYRNcqUqpMzX
TtLsyqRZnYm7iZtpFZI7NWzRgJuEmo7Ylh9+M5LIKD9B1LdfWfxPUKDg+pZqjrPI
dyujYy2bXNEBDrG7AWUf3tfxZIwXNm92idNiDneRbbC53t5hyg9YeKL5bkGp2kyo
Jq9yr5J21Hq8m4Bhe7rAFH/Ghafsd8Fv/0rtdXKCFKzk/REcu9mCX+pCzfd2cuje
W2aowzA99jH27JduMs2uvEj4Yxu26QzZcvkaIqFXyUVw9ty+70Q3CGqagbDxmYU3
s9Xmpgz3Qecd3znZgki4T7ck1KqVWCp7zGMVogbZtkLX86msqn6uMj3QQwGXrIkn
SHayrWtzWgmZ7vSIhA0J/oYNqnKCwMZqJO3bn39ySiyfCDaj8mMbOFUL81K/XsH3
waZ+bb1N+vrs5rohAbAHvhYz6X2rd9oQdfjPlhsczaCfu7359pZMnTKSUJQYes/v
T/8EA+SM2Xr0AgBrNS5t0/pUkIyS86WstXc09v3DsIcolVQbQ0WRv3t2ruBcYRMJ
VzaaRNYrDJGvMHMh8A9E+cdIHV3z3A2NL1F0OFZ5rphaefkg8DUPXzADuNZP+br9
ILPPuIdynemqicxIQFu3CgkxzaiH7pOovnvkygHn+GCYPW9ZhovAI2Lo29xoK2Wg
Wf8QOipg26OsmPg+RKGZxDC6hYIhYyB+ZKosq9Q7EecX+Ue/1bTBXjY+lTx5Fmwi
p+Q5WC1gWmyi19Ftd4SUdZUHp+txZUNr9aitMwgraUYf+/z8tin3/iI9IdLIBJ5Y
sqomYZbBbHnWoyeayt4ATxe8vs+QjiydoDTtT5WTEtVSVjGoY3/FGMcb0kO/3s5D
cHQkdjQEQHYOBEe7GmMl3nHcd/28P1Z3hlMlg+dcusQY4cqI5dyVx5YVZ719+f59
d9e0cXzQGuTCN0LiCZ1n6nadXfblZTCce8vhgMW0G++f6+kHMX44ZpyNI17Id2Sr
4l6lgfEjmHR48ULrmeeDXqxngIM4WA57jCRToSZkwvL4UGuUgAIvBqvhTFgehkl0
GXI6nzxeKJaaVTpbjkSkrr6+swk4EwfpFmRUi9S4pMH5ZdCiCLrwspEZyWSBUROp
1ubZRLWm27zCZY4/+eWD5g1nVHgbSyqxxBLUXfZWmqYSYk9XpwfUhYKpgR1j/5Af
pWGVDPdDEEVxV3uKxM1aYlvFHSmwV+KcyKmwaH4NHyOEmy0Y1Dbzi49YXkvi0oUx
dstXkrzgZJ0JWO3h/c9sAnZHkQ2XvypB/DQXgNFPIDIcbP2nYhaWWzNIMOSaJwcs
jxlvarDiIHR7WRx55Pk5ZPuMjqch4EM9K5w5VNeHH/wm8iwTTy2G5Mne45uzcXe1
kdBvUM3Ltll7uh+8GRXez3S4iQCbK0pxfAO7V3wZNZ0qj3x7WzYY94WScxacVoDD
qG5ylsVhguXCYUzrv1hX8FpYe/5dJirsQ4yUFmBh9eoWRNWli793T64UfpB4itwK
FR/lNxi9dADYSQDvZOIhKwIKllLr7ruZeiysadRhLu8+vf358xXSebX9/zWs7fEg
4cKzT6xSa+k+AF88qomKg8aMzq9NEpQk+g1ZzefBkpTjGk/zUt/SCizYJTIjHHre
x7/QU+Iaeh+iXD7LMwCmfd/uKbyh9w9cHxtIoAGatgMu4FvUNr3jU+rh3JFYrtNV
Ot2y3RvbkfMmVt/7VKUwli4xkOGFEb7U7k1qfdQJfr6eO0+RlXeIv06A0P8iB654
lGBJXc/TuWjOD0gUenQ25gYIXzQ+qUhdRFgNG/3hR7SXr4QYXGiGS2oZugxjpRrf
6p3ZgQnhUbAMfNTCV/TUDN7DLhTwTOIJeIv1gm9OUYTL4jNvI7sG+zJdLem3y2ws
+IilmQAOUw4uzQN7asNBVN+TMNISLIal+QbhqwjqR7odCo8qWBbh5wsRCFZ3GN6A
Fq35mV5calNgj3+gXh7O6W+W61jGxZCofMI3PM9fQXmQKjWLOu24S4WDko+VgSWJ
WuOcAvMKpYHMugfZymyzyFid0/qvZmtNn6lYtEuRzKIQEOB0q8ejwR0CrNMITfaB
02AwkAvUT83Wauoa+3mLryRoy3YaVZgZOQyvq7yDN+fgNt/wHjSXwvAGnHgXpJel
EOvw4FbZZhU3TP9FX2SKSln97G529KqFJpEka5ax60S1HG/xJWxGtJJ73ZXUSvkE
fP23nXT1HRPInZXxoDVPi6Ml1NNY72u5yHKYjQKLaCUjdLamU9dBwqsqvaDATC61
fugWNXBlz4s5Wr6gvmONN/NlufsW7dwaS/lbcuhMAu7vfkxu2P3PRGx8uRS2Es+b
Dbo7P1J9ewMzR+RO6gNSN9HC08r0OykQZASgLtSY1043eIVIv+Su96VAC/LDRh8M
J2zPEPGLJsBEIeRtbBp3mAwqJd4H81F43UKT7TGGrJ+GoJ4E9uwd1YdgPfz2vrbS
ScklJpaRSaomKFsK+yBM3jj6l8FcDWzuvYd3idKqYXyYKav4pvtkZRDZgTiQZ1Pw
piMc+hoRt2d4ZVxrtmQitxAH8NVg0J0WmUxLHoZjxlkYOOJPyE1UjlDhlRBc0/wg
Dg+fUXszjUegdjWvkq8Qca4xkJxGUhuzGksvJQV6ouaDeRcNkgAHL+jHfhNYgDzB
xSJrLAWW2DZW6SBjt6PD5vu8kmoeqQ1F4OMO7ZALN3qrnUri3Hhp/CbIfBG51uw2
ngVvywO+aIULZhZlHhz0bGpnHtcO31IRMSqFJcP71/Qj25UZv6wyzT5dZiJ4HVPS
7ZAjxnnb++C+qroxgS0Ig1NChyxzCf2LZ2+FjssAFOdXdGaENgRtCjrfAEuWWJwA
aH2eUzVXXdhMZX1j3dOGk3Hgu1H6SvjUmB5ecUTgxEd6+k223tUM8MXd30jcOe26
Cr+lUG+D9DOkGR4y83dquKHr3RkH/OHbij90SgHmcuhpAdB+YJL68+fiAxGEuP9x
dFGxyP5yAUqCM0nzbav8QHSKko3SzBPWP0lHa2aZmRXY3joGMCAzFduxIOq4EiYh
yBzr93I6AXd271iVz1HpozmpZwfF0U0xPytQmopNPQbtkfzueTi7Kn6449OCOHJp
NWtOv2Fy+1adH88EE7djnMyWZU6U+LCl/V4NJZqjEz8mHxWboLWTJoCj3O7fu4GC
Sj8rdfMYGBo1xbJ+tYSUL1LlqqKMJH/7GiDOTwHJvDVmUGLcLCpP3hrZ6Lj4OnSA
dweH/ahTHB4l+VNI2M3KgECUlU8LZEEm4J/j6mFd1mvNCxTse7LgKvKp5IXLWf1Q
HpQ8jhnTCma2ro3JtVhqAELw9M9qka7CHCVFu/vXAg0FVFbIfX5bH6Md9DSuOnpt
s94Oz+ENzpqD48qceIXyR9amXlE5BHGelGLZAn5zP+tgTE4wT/NAxEjM4vEmRVIu
bU4gu0XTEB8LbigG8GAxCQRWzbtg+VIWDu8qgW5/vgeugYKtCGmxKz6QAJHGQFt9
1YeVVI0UFxzzxXF4zxUgmatEsa5/4qgrUOvDEH9gBw4auPIWFv1Zv68FrujJBaii
KREIAzuA67ClFMIQdVNjqZ832Kn6zOi7+xBXKzD7nvMFHnyygKMUpI52l5B03y1X
g59aOhoKgAumM3DKD012XJ7b9rmMkoDuGGvuOH3j5kgsWYtPAFkCHGhhuzY6VrcT
Rw22p7i3VlFx8CA5LMkxt9ksQ0pF3vN/l6QaN4iI75NQAUC0W+tKPcfcndzErEsF
y8zHQ4tZctsPufZnD92C7pj/puwS1Tp5yMr3J8fnVx5tWLdFYkOZIJSl5FIv3w77
gDaW12cxpWASN+W9NmYpsVmmk9aDe9ziurvVRQfamSEJAnbLdLQq2l3ln3YNyiII
evfJmcEkCWpozezEXdACG5qphxW4QaB6ExUo/237tl/sGa6SmqbOsGKaPQv7clDY
9lnXPzSSR2TkSVjfTGfK4B8VEr/mG3FAT5QBgyzW8CqGeRvcc/lgBtXC5NqD7D3l
rA4c3gNdhENrotuLJvRbQIva1+HFvex0EPPcQ6RVdgcJEZ13RAf6/oWFgwhtsjVW
QF3GW59Zc6AP4wzb5tlGWofHGp/+y+PQYnKzRsrujzzCSiMFhXeJfPFEGbMgV/Fk
pjpvQ6Vhc2fIEnslk2PmLWf0gpCKmrAOhN+6aBpfMZqonsFJ8Veu6AvaP7QACkJI
ys35fW/bP5uCvCglKkr8ggYS/bAw/3fj//b10COLVYcPOaCbPbe2a2VdwfnKdwmV
OAY3QpEQ0XAGEzUeX4dUH3sKFTN4HxNUmSFfDrYXj5GECsTSc33vskiec1D+Lu3G
Uqnr4CHdo+IQReRCTInsYMwcEUy7IZkHCX8L9OI78C8jgFGuo4xP23d4mlTQPyky
UJlOcRxY1UyB0BryA4u7EHnQL1LOw9bQc9rO+62dnTxkJ3Gkt3WZ88ttnemauNlm
r64lfrvAdvyfKaT0IEOkdqv1wQTm0tAncLXqvv4NmNtfcrJ4yrUf/bhDjpOrEhXy
FGtWQrHeP9UxxQftfTZy+/2EihHWz/Oya/yZAjGGbSXY+cq8TLlzUjN5055epIIw
JjoTQUGWdVNb2PctVYa3fSpIXQ8ZrcSgkywPGH0+9kytgpHnaUPobH/hDhhL5rUV
4fpBShMc4Vh2Ivfeou6bh/hQTZnq43WNKiOQ6RU+Ax6wCr2WUFqyRMqp2gL39kR9
/DbgpIYFMl9PMXVPaI50hPz4LNKVunzAS6CQD7WRMtMPl24D5mUUEhljRetDUmHM
bD3aiHpiFAQZDI2/UbG0ggkUi1qPrsmAIIjtGXFq/eQDqn8wpP7AaWg0oZgXp9oF
I8sqg+9TmUc5r/fyN6t7HBepiJNwBgxhBsV+iPSFAoTC2YQ3vp2jgyiOUl21sdKQ
IfKfw8hw/P0lvIaPqKv4Hz1Tp4R8QpW0WnjCW3SoT+iw+7W2qnna+neA1w7igmmH
VfCVL3mx1Iyb5xECiGCTpP7NktECLNhIPLuxRkAF3dRFXzqQqz2zonTJAwiNuxmn
TgLYySjh1YvN9GpOKpQV2r5S8+0EVlgkwl8e9zYPyKfdUo/FvoBweVYp0vFml1xE
PuJIMDnXj0rRh24yCCyTHdHEJTmoUniAyNT6BbpXlTBnfDobR4xUd0ZTYri0OrNz
eMt/l8tvgCpOdfPNW/YJySosY4GQ7ChTbfBvelWRcqDcDZK1O6+NJugI4AwdVGxu
3QB214+N2WDk9W0RXhDbqtejDtWTOvaviudBlvJXi4wy5iFQBWHPx7qO8UEZSu3P
/aIfX7lQbv5afFvRbKL69mBkZ7uHKOMzrAZTVBAirr6HoaPBMn9mwX8Fg9cqw0AH
RKSUIdnyXIUDzBWj869ef34P3AE60U7gfAunOH8pIqBoXed+VfcQddyKzrPlIyIY
+X55/0SgKjKfXR26X15b6Vz7t8levYlo+K0+YMkbNMr/+TdTqSMd92EHiEcLmvmb
aKUhQPBc3KwH05KgW9JG8C7Av0ddzbGpppyzB7CFb0soiamhmBveVADvORDyP7FO
CEAQH8I+vWsu+iK67WN9bKrCDSpT/BJcyejmZCN4Uv1pBxx3XOh24ttkBBhM50Tt
Zs7CHzZIfjOEEuTCTyd5Boy7ZLxOAuXUP9/QiyJup8vhTRAp4M7hiavE2QKuQMiW
rTo8VVgPlW5Ke8+R0T+7LXITXFNfM88S8ppiQ3sWNXIyjS7JiVvN0rjIT3K4qjHI
z1w/xGKzI3WNxq4BRPsCU9QdLwmDB26+zB+8WN3rYAiTUY8U8xGuiKKc6qS3bH7E
72ZI9Z3EcMk6KBmaucxON0HRFyoQRrKCbfye6JVnUuUsP9prdeV7g52VZO4laaUc
D8HT0zW+2hl4r6VROlD7UAXMDjHQgM7yfnQ55AtfdnqI7qja1UKa/HN/jdPs22n5
rHUINgjoZ5JhAlrZysHVmu0OCF8MvvZNlfdIJYEfLb+37TbvfvXWW1TLsg+xbQWR
WTScp2KXjMdAmRidp4BPznyuGs7cFeIw9P++AZIhKHkUdzE9o6ZTeCRBcXRrnvio
2qc/v7Y1QazcW8hqjE7b/tBOvi6ABEkxREg9byFLYYYUCdqWKeY60NyaZVe/kT01
5LrAABiM0uDHhOhtKOAP5+2vlMPY+mzwQWFfVzL+ZAMeq59f7Ha+ECYDcXsTf0vB
HS7EIrRhVyacIGYTGM2q4TJJTmC8FKmJKTSifHjKruPkowSZPcobuRzXY0hb7PVO
O9OL7sN0VYGtMF68cMSYiW6/fR7PRlzR9IJ9Hh8Y5iNQd1XBI7Q4MQWV5Z0PzSFO
m43u2i/yzyd+iQG54tls9Nd+5VFDzKlhw8/VIiuCqJvseAmep4gCauZO7olY4aqR
zMqp86s+/SdL4wpb97bNn/h9QzxheW9wri55PI5N9C3G3OF+nAXXqRjXMJ84RQ0a
rXgjl3cEwkTNGPZKmzxejGsPWi+96epInavJH0ZmIiLhgYKxQ6yge9bJcZ4iVCkt
45AfZDjcFHGA2qIxRCcnYCh8pbyQqVNlDyGDqbJnrxA6OY3I45ih9pgtyypT47+l
6hlXByGXxpODCKeJJ3L++BEQ66AT76NQ9v91Ob7RBiqfLbGcswR9D8vDiepgUNMp
RXiQqvyZDUhe8t3vCcs1mq2V/B11c52XsSx1+CVpOeWT2DWv/3VbLKAO35qPqQXf
fonQY4sl4YUahRC4uuVcx977G01i0ftao7PI1Opjw3Bbp4a9RVwMOjYTZfm1wNrs
4n+rRmq7VynVfCAk1GCdRv7EyOHJfB2Kb9lnkhzqIkIZ5UhxsUScJFpd0v4U2Rrk
gElgMhFHGSTRASsFDUBM2acKxdDUu66PLcWmuRDFke4ktcQ8kVpO1vv43zONK2rd
mgkw6wp5Wfa+vu6cNtMv7hrCMfrvGE8dPkyBCUw97mQ+ZZeV4u/dNQToTZfwZbLs
7yK1e3EQn2J13wWRhJcHQgOaBJ95V8Nrv68Rt9J4A1uKOqLJkRNBIEF4bCn3tCiK
8keY9Ouof95QAbyfXhjztvCCZMNANTRWbCML7tahXPXXUE45v7rEiYssq9Vt1prV
I603gj8bw0srPygEXwdp35OetvqUquINLEVlw+rAxThlgRW5ks6TZhqFr7gc+i0+
wrz89Z/L2caJBpHgYyLD2JzeJqKgf0Js4sOOQzmBDAXGNrr4lcRfVz4v0Sq9chvg
wW1/DPyj4H5boHjjVTOMLsBmTsvlUBCw96QJXmonXj/ZeiAWiaL1xeWHl6lNwEDG
N0PpPBa35YGCOsQ+ljhKNE4OTDqECDJoyCUw5KRyNvwKKpLHH6ajl4lxr9beF16y
ABDqU/3kHJX0UnpFZRzOshQGBID1yNygiB0Ku4tr/Q/IB+OuUZPbztiVIyOoR+m6
5DhvHBhZZuyFXVJTpG6YIGt13MVa4bV4fFbDAVenLComIRXgPdEL825iQbUsP2iT
mv9S3q7sVwdz7py/kBDRODK/Q94YJrPpO7wJwV6kGcN+IM/JV6cwnBunR/bIGx4f
vNh6MH8IPs3pRWZphpq/XC1uqc8XHgX9NSmbdlP9GM1KCV/tuaxHzQQ31Zt/hf36
ipU0pUYjgmJocNcSEvFNaiTGyiMFXa0yI7loMPXrVzwtcg6a9cmkJSdr7H8RD3gq
SbibEnJ5GR64ZFkhANStcYYiCPO6qzI1A6p9+a74bB62kBXPq/kQ4jPIxld2+5Uk
QNx5sPdks+Bh0naQhfdHYNtaMsSFFI8U7EK2pkfWLiQituUhgSq5Q/g7Rri/R2Vo
EU6FWxnPNFP8tp0Y/LM+ACvlsqgVkUAbSlTrl1rEZKotRH5d2p4gDchR88wcyGgA
bnSbk/RyGHyKE3iAUUPtG9Y/AsUlyCRlnEwrGwCL3hKRZ9UK1YAx3An16kkdHXtf
lzzrQEaXXCvZ2ZV23kn27APTKlELB1mBdA3QpIPtjcD7UHEJNEYYaR7whUdoAjJ7
OQtwOViCsKm84ndY5++aTaeDNZlzuRTwlHElKPKUWFZWDDRshGUoprfpOgKwo/vj
QSQOmM7d5VedSniwqlhqIBQcxAZzlHT/CfOQuCTooO4OyhY0OP+eJqyWYvu+sowo
sSLkpznnT+VHkOCIKIC8zKtEdMz/M0n6+dZHlQuVYp4jXIgnvuEus0U1c+78V5AL
BQojIZ3r2Xk7DdSoTd212/omn5CcSTCMH5F7XsTpz6n3qYBhXW5y4fxxtI5RstQe
01uPeVJQdNk8M+FARXt6Gu3fzmn5fTm8NvbySZHLUJ/8/UyQb+2El+XtFhPDobKH
EV7hSUzrH2IWKkE3FTgY1niYWnGojcyYspy9UMwJor91grbiZGyEVl3ANHGEfssv
Zd75hPZ0dHRHQlgF+TXmAayp+4b9gLUT7DSnkIC3nMxotU++Zr3m1U7B5tDyFhGS
26Gox2HXzLXtWSzeH+F53EiP2E+QE0rd8TD2Z66KCricu3wGfQc7h//XcakQj45X
CKb2NNuytfOXrfZV8xSchoGntILWT5rbgyS7A7dSzNlt7Ud+3q6kOyyjYGmGiSgo
e3xGC4uke8RRr64QREn/W6xcmDTvyjMQhaV4dH53lrXqdsEXGN/n2NllIEfbXOQe
eKy/pCy3YeOtfzPtKApbKRPYG8Q+3QFj8sKN3CU1bNlCZQOMLrDapyXXQk1z6ZOL
uDFevg5L6n1VN9L2rimR8h9KwNvU5jShdgizj/tpIiJMOdHOOCmVDJbf1t83Pc5O
JXq5mcEnU1z5vKcx7OmnecP4lNuTru9uocjOcY8vXpqT551UMBO1ph0/Q4rjEZjl
qyZn+IWK2NZhXHnNkMTj/JtvTT7djpTTDmQUuDcQTwSNLzrr67jJ6AfICYbJA3uP
Dp9QjqWujKswe9/ORtgxkdlZ3Ae62J5wTTdG6K+zg6MifwOUo/X/MT9kTCgcp3yR
8VDkSJcZI4wq7WJLiwHKNtJ6SZPNmQwrVYzLepptGCqzXYT9CiOPYD8H80ALg5nT
u39WuNN3lQL+/5ykhogQEp60l1yfiSTZAcAte2Sz74yuihLdY0kk1mluIqj7pdBM
SCyAClPcIIDCQ1+e06vZaozkVYkAmM3Taio8DzsIA9qsm22Widv8Y3aKKA5pgWqV
JT4pnh5S09Yc/d8uy0vaHPjgP4IBW9FQzXlclZKRG2wHbansjpNDReYFTTEa7bOz
Ek21q2cMn6fsDriWpzRUovlA5Q3mk1FR1slF/Bs88NgJvqFoy2ie6X8sCCByljYI
qArHdGWMu288zjGbit3l0OSlyf13MwNpcq8OcqeiudTmB8f25nkPgVzd/7pvRU5+
zwiZTj6plchr0Fci3RrI1IBdzON50Q85t2Y4ZbxDRWAfOcQhMqjXNzlpdO0vRWEQ
iIK6SVw+EMQjHX90ZH/kL72wBZKfyqjq8T6yyv7kgsSa/ATu6eMBrAZ5pR4ctRYx
+P2JCXcX76MCzDHA77R7zblpHZuyIuuKfPy/XEaP8+Sov6N1gSLSw3NQk+x+UvhA
alNNg73Gtydfw8mrzPvNz+p5pSbK6pa/MuFO0Yt0Fq9BE4pwOz34I29eO2vIPIKu
19yD8KTQ9oOJFX9P9gYKJVGSNmsWmmPE2PYcXz2cmRhvyvo5inTa0AXSl1ZJ2lWa
+YMKQRwyW9Y+lpINmgPL5NB5zU1PGhOP+8l6Kl9VPEqBoPIvzDTvrzyXkZ3txzA+
KGBeUn2iacR1Ro2+Sccew1JsGrssRe9r6IZKdONfJiGJ7iQ3laMHSeWlWKkSQPgV
/IMggA/KoTiTBrq6JRaL82Ya34DKfIqUV5CINIQZg8NdmVNwYjfRFPDorRcsu8QT
jz8jOs4Vl2/ur5W7ivvsq8JZ8UsMeAG/3cdt0BJdrC19N0olYb8snPPJKORVY6Z2
V0Bkt6txYIDy1hn7wtzb8foeyEpIsvtV3ZvZuZDtv2RXkVDWFLextRYESs9WcGdp
0UVz+nfbSXGGjPb79GB4XdiubmtDgU8k+5/MtbWKWUQ8nn4CS40UK3DYRYAYscWR
ja9d6KcKIh0j78sSvLM0dYmLxF0CYABEXXjFMfd60RWAF0GpqP5Bo5Bb8Xn2XxhH
D28qRn4jrwJ2zfUyCfZj9C619zMPV0E4z1rzhJCcoX39dZ7aTkJNYAU8xMVp5A6S
XElVd5j0BeodvdKf7W9DLZEj4CM4Y2fzyKVXSKQOsuCCQDySk21HMBxftYZoKymU
u64D4p/vAYvMSyvyoMTRJ287w7wSahfOY3iZBjYXVGeHe3xuoXz6f7wKi2YsMJxh
T3n+HHUMGCAZEKH04iRLit0IZnC2JhXipH23z+gMaTWT03w/OMoUcuc5DdW3BX64
O+e7IRq2vXzv9HBnqSScow1r5EnEyXwIcUouiGgYBKf4cDpQkQPyjJmqzrQaLEaZ
DMsjZMpLw8cO4EI92lwFd/YggAonyFOcF/2veiTwe7/BVdU+Ncr8dOhm/vf3M4fP
Ook2oBqoTBpJ44lks02axm7jQC7V5WlLWwsFJf9xWOiBi9E7hPneksGR9qbxkREb
NiPF9nl/mm/rrm4SBzY2q5VffjuMNEVf3Nu4S6DypczMAQiXJE/UhIufXOH4Lm+G
AEQ3HifexFy9BY1z440CuLrZLtHBswc4wyCVw/scP09zI2VfGaDRTBXKh8A/Oe8m
e4NxEiRdT+9HmLl0U9Kq85iL3Li6j+bC0/filkwMjbnOW74YSJmxzvWBUDwZHqJP
v8GtWITmIWH/a8DRU+hOjDeTNBYy5hlxsnNpNlBe5Igr0naPcxn9hRyyUr7e0WhJ
esIhM2lhQD4fvkY4Z+Kn2YxiVGsrLdRv0GVYTHlC/0AxGZY51qg3hOiWJpZ/PKI6
SNSFjRedpqkfHg2CfBoRgrVhUpi17y4DUBgDdKyDgN23Qk6vE2f/8wP2qMMfd8/J
YKFR/FcZflO4s6O1CChFBow8qTv16vY0eoNOI6W3Il+v47mrffokisjuUsea196O
N5VXh6kXDGp6RN4uKfcd8aBL6X70vWPLRrC0iH+yHXEH4o0bWXqC5vdckIIv3vyC
8UPkE90dciCIlmTK0NhQ751F6RNr7+EtEXCYXyKmrvWqUEOWBB1pTb7B7/jMbclU
BL7/ShtnSLexpsDIzUwuSsaObKP+lyfsRp2Z+nXV4PA0Kzb96gZm7+cjFsG9IrrZ
B1Aqydg97XFfExTYIboULdoCrQVJNJxc37DbDsnTNYcz5tB/wlxm62ZgmhewYw4b
52Nx911vyyKz6SkkD9xO/o7NP+x4EkOk1utfvIYAw323LaETm2G8DB970dsipSaC
P9ZwBbgGyRvhpc7oEScvAJXNvW0AV2IhBcX/3O/qhDR9BnGVs5KQ8XMDLu1s/HW/
3Hj0cty+valFzjTlYOlsf8/uXgnU4xhWQWSdB/AlBWpkWdYDPbvrC9daKxJcq56e
b5Jk0i7YV3JvZj3fXtVjDd9lc+82GeC2ZrUI9o7lzyXOFgGiuEhLKlbPsPHY2Cpe
+6Qjwt1+/6CUr57nqAVdVBos+d+6VcMXC3TznUHXyeGaORWG6cNwDWaz1wG/Y+a9
H/JOA/mR+M9TwjNUikA5tV5zE4f9Pb0Bh9nUfmbBfM6ZO8SzYh3agsGawYWEp+QX
jlpsuX4jRnAJzBm1DgqbfCwfIntMBxtuFZKl+3hYhhfpxHJMqN2osqVAuGlj4cBG
2kmrIi5fNJ1K5Oa44ZYz5xsMRmilVYVjrnPx98S7M5fbQ5t3kXAnEeImnaBe5pTo
XVQgtaGzKg3mjoP3M+FCe4b2mJ3WJ2YQ+TM7TrmOVh3OQ+7t8tdpnlzrugfd3SVT
YiKR941bnSAkU/YshD2saNy52jbcKEcpokEU5jiu3W05w338WwMVabbSGi3h6kf5
uTkR3gWYF8Un3fCPkbvEy8HKKEWOtnTG+RNCISyR4HbUl4GXmsEVszqVaK5Efw8X
Bzo9vLALvCCZinHNCckylcJtf984v7GsOjXSATZGmaCPuV0lxmzjtTl01E5KAGVW
nNxiTMgwq9dx/natDQyvYp4mr9OG2W0cuMJ6CzrIJccXKAYnSxX0oh+X6igQ8kEf
67OJ5SluZYGG+MZ3aQdnJ69XEunMShzWVL7f/Omh7dbc+wLU/R1IjcGmNV07UVwK
iUzNxlD0pafsL0W15hd5p+z2TUHk3R32fPp8L8iy3wefuy0ls/u7DLVMGWMHIyac
3uksRkpa9p7Ygxf4GvpyEqGeqG9HQguzWC5zv1W5+ifPhGfazB8vXatxkLqXIhOS
PtsOiL3Ln2oeSdW99dda68lgw3cVNw+zuCWdwpVqMwwxrB77SQMhVCZC16KiVSLo
OJlBKHOfRTUgRUd3Ofw0xVcXc954965bi2RvYXIK1B6xXKuDdDGyQWScn9Hsfhrp
TOwObxPJlWnBOfZ2PEQgZPYNEDdPlGADcZncpq4gs0HojC5PzCPr5g/k11mJXyR8
aaTx2jU1Ute48w5KQuCzHfX7eUPEpOqTMTs0Vx1MVHkWTbnfuqA5+kwhRtD87xtV
q8IXcGpYW2uwg4nYuPQwtCkxvi02bXR5k6ssvyL+yvf5UzsViKGz88hsIW2dRgIy
HZzlK8hm/GkEEFtLjQQzCZSEMv3iaFIy32zVNZdNGunxBfv8H9OPDyCAW79ddsvA
8FeTMA+e1uWOhExwZPfpuTTka91qIYh0EyY8PIKKxRiHsykltqFpYrVDIUWnE0x1
SzLPL/3aOpChWdERTJIW5yIPdZZye6y7uRl3lMKZh6XTYd9pWqfLbvrqIbWIun+K
vAvGi/TTamS1+cFQFQQxxf6/WO84zbrPI1m+CqSIKM0wPvlg61ZUnqEdUrNQp5UM
uJ8GjZYTLmnjSke6u62seq9rgryvOEp+oT/djhgSFajbHILxskr8AmnCRv0FWSah
1tTV0n+nwM6qPijyAdzEIeIlAeXOXDzI7ASbo3kwVow1pzxMlzPI+QvJX6tsrCwc
07o1RfSGhOfewf/rRGtk05bFv9OGd2py2rBX8+NHl6qRcAjZqQAwtPnlhWCh2bLb
JZMJ42OxK24K2d5rnYDXDu+dN/4s7MiSTCR+j5O+4VdNpDoRNjAunpU0vc3j2XVX
k24fBScokGOg2Kwq1GmX03h4Jg9eiA3AqduwjNMexPq8nx3QIQnBZvN29LjOAiLT
9Xj/YrduceZnLlXZZAgy49vUdlUqmTsnEkM78mTwoVN+rK3sg9WpEN6jr4FMxIt3
RCnfikO1zR1i3IbaKNUdYj0x5NTElwbGHd5zzw/Tjq7MpcTUX4gm0pXeAxP8slhG
vgS8wnMJxM5t0/JLVhuP6UGBGSo5N6gQcvs8q5FXnTSzb3GLlWCxC0XqsvXfu8lw
525863G5W2m0wNB/pPV3nNKpF3eS+bvtV9HgOD5SU89ylAPZw9tGh57p6RTkAk6P
9YGGtc8PG+QOHzErsm3AsVeo+IdkO7oxBtWGDIO5SO/50Il9Tomsku/J7PmSsXbf
xEdo/+eQntx4pgU3C9YbnP53Ovpa7RoaA4xmdn4zL6/VQPxYWHwbDLhuOh0rucN5
zQ+pyK6R3gd1VOCeTlnq0jAy0KKmQHLbpnlrjCGCW+aEnZdF5Sg3cJELj7RyP8cN
lWOdgHJwwEJWwYEBzJX+kLzPtFpP83M4uxAq9iMZN2Ei2TJzGcJNU1eYR2eTK2te
cRXNxAL6CtXVFBkeWD2LU152UgfvGAy+Kkyj9y0+So/YSmWYg6Ggzy5fwVQiIkQm
NwvKPo0I5RqupB588eQdLa4Ubj+plgddUZ/ct8t40LptQgHY5/AvnaBVcel7mfZa
GCCEhUZiG0t1T6PUYruT/tkvQfaYV5W9ZOwSMD0xUByago6tFL3ssWajp1btgd1y
EfCQUetz1LKbWGfVXm5/WiJGdT4HUYGsYi83Xux3m4AEgyjrkmy2h6kWN+wdjqOC
l/VDuRul9hhGelhvUomX/xf90PKQezV834nPg7G/rnqSex4Ft+lZ5V2M98YF9L4v
f0K5leiOF00fPPvcZD5B+eGKR18Cy0PLb2Ii6/MFL0yos7AQqbvpoOoBaX7NfR/q
R80VMsyIaCbHy+okEw7ucavvAN27LeqY8mzx3b+CsV3t0kvIJqzLdxo7XhNM/Kkz
Kj/EvdEiDR+3ZbJx2rrd0sQ0E3iY4SJLcltNGtOab0E1Vnuj95nVhh3nlk1huj8G
QRSbrKsbAfp/gWygjLMAtzYwOmYMbwW0ljMj14frwWM3D1t8fLvKZomNoBj9M28z
0+l9IFHWqeuwRgMzO1G3NjKc2arNQ9vD5lBt+9lghSE+m/E3WKyG06y9E9cTv0tc
xssjlFkt60eHflIsgSo4FBuVDxeqCJkdOOj0SkDidqJCttkf3/CSwPK48Nsop76V
L9svFpXWTk+OCz50oO7q3fWZlhT6UqTz8bv1SCZEGThFoEcxhhAuk943n88iRTKC
Q8Pcv9eSM6R3u1hOjWZ5uZgOhbrwci7MZdGw8hPJ9dwpeZOtnz2jIQsBHumbbPOV
NNulcx+5bhrV+Tu9jwF4XGUkXCFhbyZZCJHuiD8Pyc58003N71uWUJg9DhkNPlOG
jpfK9ZedP6f61s1dwQa0PLa5jf6+VGJ9UCReV8b5mUC1MWROFvuNjr4xmJWKCiKg
qC7G7sH7Py0ifMXBBXDlJMN7RU8oYsivDIkmlaEkHprN7JMCc930rs35MWDBxG1b
1sJroX1DiB33i5yR+mMA4YLBLTXysSzhfrWJlx6vx1KeKRlu3N4zBvg+DaGCQyU2
Wr+RuPag+rJ6u2f0vv4QjR7DFSRIH3k3U44I4mocEHwEXVcHdsEQOuHf7AwdajBT
I5EY+g9wciCKcyEpcPXtOWgYm3Se7Uq+tIdmnZk7s392+QliUdspnmreJrU83ag1
fKhPWao4Jd6FVqNt9e2gCSy2nXbNHACE5BIFO+feBJNkhXMd5BuqjhSswGmUufv9
1jQZvEg95c8shr/cWhBLldl/gLuYhtyoFOB0CfM5JBccMt4HNa9XFLpMTf7DkWPD
khY7LxwUiQwEmrCd1VA+SDwNNwn5MJbuEU5k3C8SZlBeWHcRqYXfW1Bvl/5XhqCT
FsDXq/ck9FN3K30XoDq5JFlUQfp1rD5rC7Fl5ZS3BEftE75g3V5HFiR2TyEEqnob
EeQUf/PqdmmkhOCcJI0pfodadC3z6RO/j83ynv73xzHeaJkaI5u+6y0BZaCdinXj
ym1bWNf3+6XqZ1313HQbrm2f+odIc9LY9NfEyfGbl/bUzmgYBQ/DcyCWoAw/sup7
HWIDImKcG8AWTNidX1cq6MnXhc22cHKWm2LqZ0ZmVybo3/hctzUFRgvmHgHpjjgj
DAeT0LbBxqEw/Auskr/bFLnuxMLTqwApXiEyFmjUPsHs+411q3ASAJqAL0UMxN6C
dqOvaXnYeWc+8V9wEXbmRUreQF6JLy8J5/KVDKPYgAj1x6SO1SoKkJB7vnf2zCXn
CQeCAPF1PmYP9NcrSh4/J6a2gZABYIMSAWTK2B9hEiX2+440H6vOD+7rPe9pcc8y
bdSSb3TRCsDNN+HplFnHe4erP21tSTG+eeWUtbnCxGU7/EYaiJ+GBeBE+rpLZ7Ac
d/0JjsKsZIgpO/CAqKl1DvaIXRVS8oL+1k9IvX34A3TaTF4lthkOZvi79EPgfxaD
hyj6aX585uVxh5bmycPqy5KwCsHRQmJBkpNb6/qJg5RE0zQ279D2p8XYCRj2MQHn
Kr45GKX3KuafbHSZDiNhzaUYYl/4XkZ2gI1HL4UM7AKQmmrMOr0ccJyFx5E/rz5a
PjnbwiyDs1oywndiPROhOulKB61tgcYRDh91XU16sEh1VWelQbD/r8x9tLM06N+6
4+FkVzZ290PCybqBggf9d7ZJRpHY3iNBfCJ61Q7TSPWRWNBcTrqmgSI8urBdvSgj
WYsoMaB/30KG7cJwJxqY0ZRXfBzm2i/UgPhYSRDgl96qbVN5f9HSWja0nOvAFff2
cFYAfUkgTNles4/gPQ2cFX5L1PbGyi9XGRKy0Ijw9aX1P8pj43fVzNdRNRLgTp37
DBo5NuTAadSIZ4SgekXol9mLvY40c75EU5ol9wWjB51xHdjSgVALbGSs+tsLPTZI
utXhqwERFJ8geujkwvfDwa48CeFu1OVB5o4sHKj4URqcwJuliVdbfqhDP1duD9t4
DaaFWDE3wn6mLfJ/i5OHx4unJ1pGVMmv41Fn8M8h8l9yj7RBKrSIo/49f33kaDJ7
SAHLF2ykXpfVVMav7GFqWF1fRLp68+lLMtC6D/TEjlkmJxf8Ol3RLKaYvUDP54z0
DwPCAXBcEAW845cS+OX/vCNVKmHN/LalKhIHVqRi+a7XE5sPzuW6khz4g749nYJL
YK7V27SA45IpF4hIZ1wxsQqio4bamH/nD6ertOLKu2W7CDanFhjpALhW/QCIwyyk
PR8wBtYSAIEm1xqFjru7bjdQzA2FCFfFXJ62x4IaNjra7KxQrJNZDiCgiJ8128v1
aXaBk0LNpQ+nlSW7wiTgXfmLLKRi0FRfygJb0LdxcIZzo+PRAfCBfhaDej7HUvcg
7pIZC2TF33L8KjvpPAH5FyYfH8Wulj3t4E8QigV9hdFDNitvpC0O6i+tqkjhP3rL
NI7sbaizPh2uqO8pYCQG+v4Vqq2eGHg0pUifn5X2SUBC99Zl88Dbrv2A/Zf3eyet
rkPMDRA8Wur13GF9D4l8Ng3LYFU9Q8h5We/60BI9hWrlNaH89hpsmfr+7g+MrNbB
AIe4OTLCiSyr2fMJnLctpJTX/2npnoNgNEyoQqmLaA38p7criNV1EKVGeibt3zsP
hzsUht1vjTR9DOSNDWM4FKsxShPPRZXUD6Un8bzMpr57B09ywl+/HThgS4HIQpqD
hIkGXE5GaBnY+CZeQQHxdD90oyxSlKv/TzPO9oNPE6WxnxCfZRAIQ0LHfbKFxR3x
t3WOTO5IGZJSsM028AM34jY2OqvmSK8IPiY8gQ2BeNoTwlCSGxyNZWFEnYSYh+AV
axu3EeD9Kl2SmHM8ntxdQB5sJbjvBOogezTLItRudg7MSVg7uyfxJ9ya8filEQTL
QoW4K4YN/4mULy/+W/stNN4aOWfYoYeZlHEPIQX415C3BIk1jUyzkjORFPPCFVwl
gDU86BPub+2iueXFZ1opedCg2xR3bfBTqXTeOsc57FImEAkZNMFwbtCZd9fwPsjN
bYMI2RZUNkFeYZs3rAXIG1J5vsb/lOAwInQKnvCoxFN5wC/+tmRrgavOOiZpH8jV
Lc3MZc16OoG5Vrf+HpZdcDiV7XNU0XmBA8pTyMc5XkLQsW5afJsNADTUn+g5XFar
bcYC3ksYv8D0+JhrdUvfcdRFPTs7Dtlvt6+6qoertL6oBhPEmJ3RZjyEBClEJ3Mt
ilJ117G4zZBlOJBnzC94N9rL/dJqS9lDQIPRKyqySv4sXOupthnZbMROTyWuadlo
NVu68OaNbtMcDp1rg+Lux7BzRpiMpbhUFK5Hw6UgDu3+0eXTd94s7kvg274TI9t+
rvGMbr26aod/SISL+B+A95CyqY7rmqhcuaDzR5udhIOTW5a2nFsXaSIgNg7j2AIi
56GK+1PjDBM8ZOu2FEZg95R2QUpU5iKgJA7G55Q8uRmNKpTfqvDMvyNVI3A/Bvfs
+JuUN3sIfjRp8kYajjp4edVNWra9rwpq0np5KlGnB3jMtssEepqCGLBdHh4H3Pxx
IzD7q9PSRJ+B/djByzrvM5ojbYdaB7KAMR/396YO+GehseM2djDY/yFuED6w8mPF
pEe/uQG7Dl8rxbySnvGm18PLAfBouB9N2i9Fy9/WQYS+9Kpd+YVt+LobVVH5MYCh
62PIyAu5A/nwzKLt+QLgMTj4Mx4z6DLv06xibWLgkt0RfXlNwIgS9Bgtz/9+cUPS
b/JO4MXxpDjLLgqIeE2pINISWhfSWizAltn+CrjuV8PGTdaQyPWoO339nBNb/3rj
iQoa8HnExdWMfMhO0RBjyL21qhMSOrDyf9vC+RBexXhu7vJrsXTR3yP2zucQM86M
q6z3Blvf/padflA7sI+qfvw47ZtRpM+rdlKZCm3M5jlKTdJ/v3NoNgtOSbJ7sBff
v8K7YPIReBlkY1oKqEgitDytPAdNgpzL43km9wHewCvjx8bYmjYLdOPBW6b3hYFf
Y9/2zBPIpwb3EIVzQPwEScxN/csmodQqD1YkedQW2IEHhX2BgXriwxWBakiZsEvO
NnT2rvtRUkn0GegIluFnFX9M6EuIakmWyy//sohzV5jIBrH6NVvGT/40RIcNKp8a
BeH0tk+BS2T7RLMYWPHzFQ1tS+d+m8wFb/Mb23UEFw9wlVkTBanv9gqMYC0Q2ufe
qn0EMErSzrVUCsa2hk5NWyprcBT0yNFV/0GVPnx5GWTXpRqIUgu8+HrlWc1yitg6
6tTPiFEIc8GysXgLCC6a8HZN+gqZMlHinLOBxHB9cfvKxi5HNrgK/JJYnhsajOW7
YKjPIcTHBhfg37xvkY96GkXEGWw9ui6TGRZXmb95zC9KBDn8T5tf734rsGR9TOZH
JjUc5DVUHxFOXApwq6nhM8SytZMqp05ArouezLcAta8NimyaIpic837VW4q+RvV/
lxT7Z0zFuEA5Rqxrtj3Ta/VE0kW/uDncACFKpHyNFF3Jq1S3YO3jgO51T1T4FbC7
gfVdyjIFJ+LQY4b1HTzzH2R3sxKOiUIn7cfT66lrs4lKbjDx4pmKUdD7znK318rj
u33zp8kv2XeT2blXNeE77lIqKgypyHWNigOfwyviFuO02bJ9CPd0kKBJ6OxAE7p2
oR928DNu0rjTz9JWkisNtZzrkDhBbV60nWJ+cOsyJ6oq99Hr/AyhfPbvJyJuGGCe
3gTG2QjQCHymQk7BxIRufitfefiRWHs9foIK75e0dzSO957KLIY7t4h9F5qzbH3/
ViVdRVeg97YUqoIthZL44nSosbnnbVhNUHBLEHHvXmfqWLrYvYJ2p8nPtte6DbgP
Xo/CDGA/E4tYPoRsMkmNrRMEG9Bjo352fgfXnzQ703sAUKo+En8Fp3jaAYW9ctV7
SHCQjUniEZ//Gwljt2nKwEJtVa4/oAW2FAL3kIcTY6x4m5+7tsvwsyy8rudFx7TX
zS/0Oc+oXE6jwaxjtzjC7AC3wR1OGeTCjMzxp+w0AI9vfx7Fa4gYcSnmLnRZNA8P
xOrZ1x/iTzVpbB1QfEk2H0gQGrhtbaHYbxEZf3d7y+p1mfe5klAegoY3z92VrpbU
abGCQMexAJuYqQktDNkpwGHzCV4HrMjxmdSzgy9fpABiXbmLs2LSPsT2yPErVSNQ
GcxjDsiPDboNpwVtw0RTobKPn/NozR+G9hAeuRD1Yep5LyXZIUE44cpQSwOftk9G
F03102LnB+2s5HUy1a7qoZVTj3o5hRghfBc19LjxCMAT2k3yg4YTlsexdIge0b8O
BXLzwKfGdGKbMeDGCTddj70VH6PgUEwf0rsdy8LMjJs7K0n8BldXRm/veStcMYSx
FhvAagVYYYDo35nth4bPX53g3o5b9+7haw5fWWhYIcZYlm60s8WzXJmuPR3ofky2
tOsSqrCaAcoogHj6Ghr9aPgctbp3gCTnUZb79YAwLSErdzuwwblOzHoIi1Ew2ZIa
9DGBFpx5IE5m9pybXUuhxU0ryEtuzJCmY9/RJYttPDxgyCtty/LPXZhd3IvXeuE6
J1R+PwUAnti8jZ65ivNb+RwqkslvuIn0M4cOsOBJke4Sk3hBedv9YNtENCkk0wBq
ezWheSCiY059ZjxAaSnOrKn2XZ67qvUcH869GTjZqWjd8ADMk9KTc+WLUOTygam4
DgdFVNdiwTKnEezA3nrFTi+Lvj80apwaupiDIMuBXmlkZgh9q4P2NOP76hvnae3P
AcHnBEIz2ZKpj3HMK8u/pCVh4uHfg1P4NmncOsbNBHJtFZjS4uKo7YrTP6A/6ukA
AVa7s8+/OXKlpFFAvZXBrGFfPMQ6wdp8upqaZAu+Q4S7A5IdweHtpDXG4c04rgFK
p8QxS4r0QFsjj3gZAy8LV5+VNcJ3qHFLGWko0wA800/S9etdun+4S+YfazZmV45r
PJxkjXA+BeuqJd+RgZMxi/FAihRfqSZ2UJcDyX6Gd8s3MML4kYxgd7QN3pwrb+tC
e0z4c5/mv3ydoDQnj4L9CJmKsumDkaBETRYuy+oodJQxtzhLmQbMdV4Ii4n45KzF
Pv0rkngG6JxJZuj9AJ88N20LODrnWYk9QJ51w1ab3SIXiIn7z9pEYUsVbThE7IvG
wULKoJv2SDGHla5EDb5DKjVABAlOHeMPrmuQSHDuqlGkELlp54mQWPRRqddvQhlz
P2atwHykcLZ1pex5Z5mW7eaueNZVcynCDYZs2XBGzViU9sJh3mrL2sUygCZv3d2e
cgOy9H+RK5k9dKZftualoJWmnrI4w0go3Oc4OtKNeeTmzcE81UwtMTgLxVlYyuqV
KnO2Owh7YDWbOiq8LRk7dDu3qV1aCdk4dk8gzXTRXG+TsGc4hodJNcSG1ZfQAd4E
JASSDZHE8Zhv8VjyQjxeIlO9fKP4aobCLkPYKxx/xLc5l599zqAsSODdd4NIOiKh
8Xpxq+ewzHfee1Lq6H75c395D1zylxuzjvxdz/bXMIIzS08akN3Y4gfBjvjRDrsO
Qe46LoS1rKl1qoBwdlGOTeq/87EEA2nCit865609Mc74kw/4C22gDePtb6LzSuCN
ELVdSbSzBOMBfOePi39UlDeI+77ChVQQ0unyUEQXhTkUJFvgOaoTCPqa7+ejhmdv
GnZa9J/3H3Dg+gPwqoX11MFh9N31QB6I8bVtjfce1aFYEEWGDLSvWR5c+9mMbHmm
nf428udxKXZixiWPbSgL5rMnK/jsSd4KnxUgvBrlLomWMRNeKmde2SEANB3Y20xx
BmovqWgN/2i4SmhU1mM4WCl+vnTnEUaL0IxD+oz6LZyl1w+gReNIfjsClq8h4vIl
iA2f8c5ADmQWzK/p1cmsjlpQEhwb2cc+JYHmtKeONH/NI9UKogJpusmTbVM3kdkB
8KYKaYpSOTpStcc2XElzFT/GzYKA69MTR9BOwhn6u33XMYJE0EexGZ62fK7ljSWt
Vb3l/U0fV7ruQjqY/e9FUrV2DMFe5/va4U6X0ASinhB4yNEZKfvHW3Ac78T2DHCJ
R5h58g7nYjUlS3VRCNfE76RGda4hKjFlkQTHc9ilo54kMgUFx2ti2rF2lPEXmNAg
QxL32/5znnzDAIFvRZJBRxcmQUwECmoTPROBQC8j54JekRQsIQaUDdHd6xGs2HpJ
dYuK2TDdKSUKxZBKF+YXWBNO2qwQB6ibb+HXo8JNe1RoSBG2qA6VdNSSU4nDyhyE
GPgg4eUVEuT54dZwcXl5WdLtjIJ9PZTx0LyJ7mjHEQswOD3bG2FEukYPheCreG7w
BhNvgAH5YIHJX1q98cm87xsOWozIPbmMm02k16YDdgS4YZJRxXlAUeryZhN2qApK
Q5N0IH7kBHj39rklOE3OQ5hH0bZA/g6nhtkBSFw1fuvxfZO5gthJ1ftreu8I4GmI
ILz2o7n00DU5Q7sDRK7o2YyfZJoQ9q6Z8Dg78HpfMJRCMf37PSLIM90mRnMxRiAe
UigVA7upyRoS9yhGJ+VPVxP4TDdABp3VImiPveTTDurJA1FPmiWzENUIxPrhoECA
vHkIuSrqlSB2PyVzY4b3fG0MzPIeVJoc6P/C1sXH2Fw31Y+IlcwXgi80UhKv1pZT
fcpMQIkTHfPsq4xZPh/2838+sHe5kfoZycCgGrmLJWVnYN6SgclTrmjYLt9EJBKq
9obOubTIlkctBXktpQDy7qnkody4xjfpfqdEVpqR+jkv1L1SnHXncZTLOiDNAX7A
22KT3/pG2OzezHdjNwwyW/IUMq6y/Y0+SCw56BWfx+hUTMcnpO1zZbfO8WNyvsOF
fv0LBmbaoXLnEa8Y7mjAT16zN6LS9+/siW93BNHtFNJ/HODhud8MPqvCEyHNRKIw
w3WPvTq4gO+iKbTlqq2W0N7C78XMxegttMHvTL30hEs84iKO+PLm8TghVfhNX1bV
N0e4xt9NqIBE1eyj1Xq8hP15NBf9GQhjMDB7ovskmXpGqWFiu2d54BWMjKNKAuiP
qM/DWg2aGP2pOxIubCvIuuoNVTgAZ5AXUrhYa2C2ybahlHU4s8H8CaWWGZxADPl6
TlE5M/rzo3395MRmLYl2zCPyTdDbizu+dksV2xoFBrpNRtirqiQ3xMYRTw8i69uh
4VkcCaey/NAv5z5MpjccYcvt9jHWRPUp8VCVxZUzBLR1S4BoN+CQNeUgWwM2qa0F
5P44+RwoSHRWmBFSBXK8FS0NEFWSG4BmesmFubttH5P0Kzk7Ip8mQUHJNSF24DSo
nTJ6qt4cDRYgWOqYGbix1Msw8eWS66vwmWeGJ1hO7rOM8Uix4lFFu2KJgzcBBFYz
/tV3464pydLj5E+oWiJuGbo9Pp0vaNaGrOT9Sc2kY6Q4OU1pBM+JFfqr+CZaO9cp
ypEK1X9YfIIff9TrLKBUXHQ9zGD0asI3qccgtlN7IQ0EtUX3f/W/vMMdc9DgDYs0
7z2lyYN8K5CQB5EfUMkGnZVX8cPN3AReJrDhGMeTCZ++LxWLuPjh53Qt0TOpI6eu
bxnfYNLqhQlOjoHVOm1NApZvFE6fV5ne8KV8PVpsD65ivbMLrJ9aUpXH+E1r7rtJ
4sxVqJLGFaF50BJR2QzVZHedVpX/IYkaYng3z70PPrD+vsh0bgljUY7fm7dw7Bjt
FCJqP6y7TfPiBdapRgKqf3VqoJnPieQYVD1riSXbLmCaZtY2wG1tz8c7eyifjKUl
I9oXv+iKsVV+bQHZp/+lkv9wAZR+mfsibeNhR/A1Cg644kX3ZoIVjySUkEMAmAeG
ffH5u8srwyOL0roqLrneC45lsW2gpKKUrnMOjShOsQkoJcpGZMdUecMOVWmANLxo
uf96WPZkawqnWTNhsCdCygp7Bd1MDdjcFKKLagYQPeRcljcBh0qIu+ITSrihvWBj
dvlL4h+9kO7mq+4mbW6A9JGydZSrIdaO7R/WDRgSWeA1IAxlXeLrenJ/DY7BDj46
5rvhCbeXamixsHJ8wDCI5V3rUzlnA8WG4MhWMQw+YENCSeqYGRoNBzH09+CQ3A5T
tAWoQrggnQVrTvC6z4Kk4unY7P3MpcqP/GF9L5sOeryuHYmJfL2ji7vdHKed++ri
bCSBXcc4Zc36+3LBV1g73clR18azML1AoVvY/guQIWhP5Rn3Vt8nTWq5cWxTvhHA
HQl79vMxKBlSJjc4NxSbbDfHkD1ck40C0VRUoBKSsJDoM58or7a2BgpspH1EFWOI
qo1Ef1iaO2BxlU422EcuDuAZQVpVRX40N7xVXhEHXc39Uu/qXUcYqF18QXg3hrXr
0In8ahNvvI6QeSLym3fPdb0Gd5mhYAuUBqXaywMth12XregeKozZI3gUkHL3DZ4Q
SWHU36HSkC4rsnYZ2Lb0MYeBzCJrTL4Nl/l981osbFfuLvDFcxJONDluq+3vmQLU
arr1uYQI+5s+adH8vGc9cl/uanZieWCp8iee0Fhb5Z8n1ahRgHadr1Kj4pBVmaip
ivArMyvcMXHBq11DSU2/tCtJH2QcHTz49QOq6SpTY4qPQiaxvXBB66bBa6WdYH5g
oIzgiz/WUGQD5svxMuvWFAuYbfq71mSQ8o7A+uKCX78sCeW0fsg6h9EtL5fW/SEZ
F3Aku9F40pXxUy7WTzWJiXIls6DKs5pZZBxg3WdpQGaKYb/Bys6ya7R/m09t35dC
XXmJzsKyrJSQZnpXmHPEQn9YqD10G1i/jsdtuXfw7IT02Hlir+5hEZkPObmyXoeV
ul4bOX6BjA5l5msHXMB0HA786xT3YIEfE4yD3tsIFlf5OckG3x3pIQZLYjsJHhe9
csGb0tWEnUaXbiIunh9tQzlIqu8mVyt2QyfCt93+Ne8GVeliX3LZN1KTBgpGiAxq
D8OcgbIGFccAPOhzd9fEu6C4eMrd4pcIEcyWiC0mjypUzq6ny/QMTcu5ro3V0aG+
Y3pZ69Uqn9BKM3k6UdUxhy1GUuXWkmb2GzNaahf2zqqgK1gfv61jFWmr/f81ctLS
2JfLLLUBfHzsWct527XXhHZs73vNt4shr7IqGijzRnsJerKPL4rgW4nRynoFR0nc
OAAhqEEK50GE0JfWP608aXqZ+p8YgLJuT8vIWDDmbQYna1xC1OQxUwP5GNMJ2kjE
a3MKH8/yT90TPBvwm1paeSNZbOMmz6am23fUSRNtRTQ2Ra+Qiq2AI8UGaTxv/41m
yrIXffZVlHRE4NiE4bUcVL7+pfI2FXqAClRIwrgc6MqBvPD3bMCAIQ9YE6wtCMs3
+qgCT/ag14Hozx8LP9B/y7wKVSGO18FnG2ooJ41a5BLxJWGsfx+dHoJ2F8o5vAr+
/bj7XdRTQgZVlxf28ixaup9Dj3jltnPcvTOCkU5Ib9CLeCZw1ZbrirIGJ9H5UJGQ
jYb3PqbgiaBUWcoGX8/ZOPn23+27NkneogMZGKEJMMvY/Zz4Iaw6wxNR6QcDwqIe
AyFctCJCe0SK+pgTlGJx+BA3VQuOWI+nEEIeHpiyVWsDNpdd17m02EwsnRZANnGG
nxOgRFH4IxvHVia9qcfScP6AKSTl2MjjGf8eFHT3DfNyCHvkxcZ+dJvPW0MH+N4j
RN+C26hXm4pXI6fBLDdPmGvQSuyLzYeTyThoLVdyhkm1shqJnDQrJShwP3NZh21r
SVKg68YQIILeQiDzmOLrNATvrWPWRlljNc5jMSUQbGl0XOWRRjdToGaXW9Amlwx5
auUrwkVTDbqAVqTyTYB+V+f9+YRllwNPA7+o+EzvKUyBMWgrsCIOdsfq8hqQzgo+
+XOFPE/tEZsPWqhhrI2cl4ODcuBRYIEyJ/dX5UO4WdyZOZm4zG3xt0DKbB4pqdu4
Tf4KQqBkZM1tBHJq3E6EA0ZpgTR5CTpUUqPnAFrAX4k7dxsBlFMDI5cJ1Dl29K2t
i2DVWeSmSpwrH3nTD8UFmhg45RpEYx639t0+sLTn35o6lKQrrejyeudx8RvtR+zW
W+NefzM8tdB14c3KvSFy3upFyYB9rVPIvPgJHRFgDjkhJblp6FYtHFP+39qNrTKP
RCM4UDCY1x3F79xGkyKFN6yqj0GgUls6Pz7HZPmOtDfj/4RMyhbXgKCo0MA8cJvB
nEn6nE/L1MlfEE4/P+v6oaVwAaDvJYb2J38F99rdiXlEpztJbwjgEFCXKQFYiWVI
vnaGUvk7c1v3ykeraBcf8pN51IuaPu2mV+f9VsUxay81b/Ite/+wmpDtsZG/6Lzi
mZcCYjyBc5FaWLpCBqvnMtsoyKCzB9zNTLGdAja23+v7+9ZyJc9tduKFnGKefSS7
wTUOmgDTaJIEFzu1xvUZ6PC2mZFlkpjlPg60/F4Jqzz8UeAMF+DtkHzFbwfjak5P
+sF/9yFbNLZ90gv4tCftNQ3EhDrD69jGKpUhH/FcFIXg6uAGmfH03rBLGlMf+gIB
TF2PzqwhqbN0C0PFTRdeYw67MWDkv3qPnTeCPQ4bnMJyWMkAHJT7j3T8uEOqHnOC
qS16fqYTZ2pXV7rVFPwvuere0iqO5B+JhlWBo82faQLnf21NLzafXoUKN/k2UfFN
8szcz7lVUN9AbArGFCjOSpBAjggxBoDRkCv0J9dNZ3NWawtn+p8OSbgs29ZPH9j9
AvUrGbDD4UrmrjcuOmMLi0/fYzcWB2NcFPdV4MJBO41rHKQk7fKoU9Z2XYv6Hp3Z
Evf3173pzBlsmZOmvgoEikcliOC8nbxRtZczxIFkk85UcQf9xxQEugR6MG/Lztnc
PwqZmXSL7BjnEKJBpRJ04OPjnVK2vdpIbX0BCdcvN0GZOW6++oj+v671/d8mltlf
kopbnnkEhAqZdJcK2epOuYBoZlZoePFuBcyTkHm2qNgRJc4AFW28NwOidSG0PkA5
VHi0CtQoQ2gTOgOSxJiYd1GOb7DNc2vXCVqOE6yC6h8Vy0xxaOEH2LTqZgW/k+Rv
ksG1u1lgaMGLM14nRjPAGCioJCo7SM/EJ85ZN1YOFENyp2HIbJT1fNGNRTA2rfkt
0hCPEhDmzlKkiKDb5FF9aCIUiKbWwIJ4UA2f1YVNN8lnn/niFFQo6nsXCoo6hagY
80FlYGR3AfPE4jWSDeDQCJgizPikkv0GplV0HsNK78DtB11sCGlhAtiCY7Xt9Lhh
vUcUs6MP/vomJpPNizIp5nLFhZqbSpc0Gh45aqfwy6b7YKus0adS3yC1cwp7FIMK
U+z9keN/uJ2tBRSll5eu6q9w/y+ZDVVdDPmaw0tHXHh+75VIL/U1hgU/jdglNbbs
BY8F5qO3l9Dp2gmdgjySwmZkVrDiDx4L+sJkpX1zx/LL3mb/lObFhQKCQIbOfbbe
Q3bzzph5aIs8VP842b1Pa79AEFG7ig7BfAERbcjsA/ylZCxegjuOxWfYMMShPMVL
E5cV4XzS3yI7KsQbFgj4D4kp5MQkoePaaZmm0U1Q4QlExEmkX+O7TF2dWjQ8j0yU
pjJrueIy09uwUXUuXWO461GBc9gJtWJsx92vcTx2emuz4mivHFp9jqIOqDmsSUUm
tv4atPbuTf70LlEAKTLdmIayOzPAY9bSDWtZahOKsqFuXwz4TFKovBT9um4vBQqE
3CV5b1VTzayWiWfIefOTGBieR4AWYAhqJecfR5BH8PSWX//sGeaSeAzUFVtSaONJ
wBjXthDtor0p9SVGqPPEIvilvzEuAf1gt+cQ7Eq4zPro7wkMGCbz/8Xctjr1JuFl
oeusZrkLRbpw28FsKNnr0qXsxRX44kgtQyobFJe9XKZWcKizXIIjntmiLTBvFoUx
eAmqOA9oFJNgSiiz1of4cXIn7ExYTGGHD+Vv0u9v47wrcpLZtksZySsGJH+CRQDd
al3LP+7v+J0enFJsca5qq2gCsDmzq+KIYGEsNSPeEYeKt3CtZ2+XHRSAf0lBMYWl
czlWMrSfTBMOafCEdVswPOSAD/1SvqsvAx3zN2dni5WC2m7JxHeM4aY4c9gXf0PU
4ivco+Oppwurm1kOidqYFReuD5dK7flr0qejIFWPiWHxFFlXC68yHDlcOx1ka6gE
7Syeb1GGsB51ohBGMrLlzTJidQYfe50+kug/OAAr38pBSpQkgjY04LZACUHENM29
DWomWOVcN6v5mGD44B+JTpTyDp6/ASJ0mAk4tSVD+asIl8WuB8QAdYguAmKgHwcN
XGqeyXo9OUIR+xvOz/vrcewaGEvfKM/2YFcE8H685JCS38tWcjlOl5klb1UCJa0K
f9DSgC/ZJvnJEkoXpY+ak/amynGOudeUlWv2gB3rm7DEf7esdVGqo6RpExtEJfNP
q4TeUrikvVl5W9PkGqUZjeKEWQLrc1+siRSEi7snOZHRtmHj7ghV7FlINhzSAkRK
ASNi3mKGYHqW7aFLLYCcoNHY+6dn4U9s+nf98GtUH6VsL3OW3r20W4q0n48OvH26
OQwnxZbFeKGNg8lrPWN/NSy04RNIrFV0WXS+7Q3ckZ+naha4aF7/szp3s0zeAswW
70Ruoq8kBcKYLoU8YqeVYvi1NSUYTK1AZmR1oJHdLwuqhN3lDyNw2mus/ClgzeQa
r/BsG79y1M3RcP3sl3oLzLu3XOzHlrrwN8Ky8JC73msXXNkSF9yp9whBOfx5E3++
DQhPX7LaEFhdUS8/P+zItUS8W9FhqTKNzCkf7aWV2eo2fqEn26n0D3e80w6J2PSP
GDa/BPnI10xPKZ0qkKW+c0TuUrMHaNM/9B0/ibZUXUYNJlofDbX0R099O9CSSy1f
pXU0TGhW6jomR2ptnKYLlCG22YNvTBSyBkGjEsCyNKkBVev+DcRcSFC8k1m300nZ
pJE814JhkCanLRsiPndMg/agfEi+R5aGusGt4cIu7pPY68jRWbM8+ksPi1mLQN5c
wHWRyiVOvj/MB2lULc9/SwgkPWI/Wm+kKLbdPZmm751uYK+7CTXBLIHoc6fxw+aJ
yBN9j1YrTt/vTPvasc6LQ/a9a3JllvR3nwKIDvG5V1xuPmyuadmQcdluWudOaznD
7pm4iNXDUaMH6hASkuTPApZMOJ3rPXkNU+h/v93OMGv7wv/VJHOJTEM0BCPefOKo
HJUKC9AiDgXi7CCciyBFCU0dzxigXgO/aeVuJ/BexUIsBv2CEmyvsEZsrVKEngsY
thnT+X8iGoKet3Vdh0Xh1Q/s1s764nF5iqZ+8P1w+1T0PyIHDr5lG2HEGT2EuByN
rGHkK9H0GWIUGBVewGQBPpgXZYNDKwD0SztzlVZZ6lD6NdFF88V6il8zwiW0GsxE
e9HliU1kpg47+uMJ7bC9e8o+jffa8PPdtoZr1X2jyC9cBgA8s7TqDav/E8IrYN51
/XEoFX9SjRNf079E1dEknOHsC+mE7Iu9YtA7VeQ0J/iTEwCc2JsgnZAHbisRxw0D
LPol8qcck0is7DW/0ArZPjIva0zPLYq1sOYUDn/702+YLnuk6m5SEkPxwFaIbOVa
MsO6L7gZeLux5S0ETdk/Skx4dHzUrGhcAcO4tXzr/8FXPLxvwG4dwDw7bukCrzAk
Nsq4obOdyAgT27GCINEMD/oVQG1i7vfAAMd99Rnuvi3uKd85GinRlvxl9Ttzik98
RK17/Tv7woSgiCXX121msT26CRc456k6iWuwNbjKl07tK+w1LDFQbSTvo8xsSFfA
iCTB/LGnY4eau0ZP15bNe6dIRRCIvLaUEhYTSbGZuApb2MCLQjSuzU2XdHlcqdf7
Ky7TeJc8RRe7dtOYVw+MXzzBlo5NFKm8EfycK1EoWKVK2rJiSr8+lyrk4Qp9iS/O
y8NpAOrPEGaXD/4AEfE0UUSx2B1vRo6GUyioAk8AOh/0bI4+vTHGo/loqSv7M3zJ
hUTsf+Fs8IyTerGtFX+nKEeEpBqFjhGfMU0/FOpuDv2RmdGnYU9JF7O3aDgLXq3c
w6Ov075rshUuGgB+X/KjCYD2UKbDyjLsKQ+/T9CLf1OWtAtkJ0mHAqKxgspQDU16
vEyvo2EfE0hcL1szAijgCYLYMKkTyz2/IzVdmx4IQ+t9OZanjWz4LOTAK6f13Pu1
FeGMDtnBSx9ogN1QaN3WZcSYmiRxwQjb3bTkpSBI72rBSxRxXL+fvMRNBdjUfucg
8qcX0SUf30r52pEhavOow7TbVnoH5pjHOogTW/H7RgPgHi6I34WxV9Bi0DbG+3pS
30cwyNLObVt2lq/b7k3FkFdO6Wc8sxAzdJoknwRfpiJq6TFWOYDPDo+0S/bN9oh8
pnxvpLnQvaIzDLi2CoSCC3nSFu7y5u2WxtACKVpI6w2mQCLQ2UMCAYpVeaxWhs8L
Ard+dk3icDLD3lWjtuWUrylyktl0q/H3IGSS2TYUXpPocaodDMF7+dHcE/R1Xytr
RfkcTphnnnj/CPTJiy/Nw4zfAoIlObGOLJ8Chp0xBocd3QGlvX3B06jVDV57j5VQ
gF2zuuhrtJOHQ3jKZYMMZjFh5P0JOd6qXUCiGe5fgGLEsPbaXFvh16pZXda0L4xm
t7n4sMs5B4nCouJpDR8/mhR6WxYJukvyuqUgJMagFJRLqGIP8m1CQXd9Aivlrb4n
/eZUfYP3DbyI0crluYadTcR6is8qBuO9KS3nicVpQ7CDCsH4al0x65Ea6XUDH0iq
EUaYJP2h5ZxHbOoFm9qtW5VBEyMP4snm0ISGlWDf3CyyXPxc2CmnHk4TAthI+CGk
OFf/GDGOKK/RQfL/LVrEB6sWT9f4tWlOZxcTyHwGJPNt9yeacCEQoZW2iZOzatCa
EBoDySUyciszCPohB5yb6nL6E5RoCE8BUrxxx5R0je3e+I/w3I+v3eT1gvQdEPDA
jwdtBIGFtoIVIL8DK9Jchs4bfrdeI907lpuPKmA2FcGciB4PbT3r51B7lGleNUKw
whOfDucCDgrEJ0bpucQfu5es9q7ok/B0nMboaCHhVn7wX3p+uew6fmZIOiQtFXKJ
RfnV4VCZCKpTiCyeBrRGfmQix5hpwkl3zH8etlA5yWE8s6feqp7TvUa8O4Kk8lbF
eRBLwyfWqQDZ7MRwyHtqmETA4m0foA0wEw0qJxadQPeWVelQ/40DB8mVhZswM5Eo
Txv5Nl/ica8M6hE1oNNHQpqz1Lj5IkbFnwT353lGnziGoA6b6mN9zHJLuedlWgxx
rSSMuSsbzvJPyDi3nv2Mz1ODGLKvQuNG1UEak6cwH6T5K6mKpfHuAOQI5oci7t6c
lsUp++3k3FSfIDDJh7JBVISyANoqXxCOi/AHj04UbUL+FBp3IrkhDvRE1s99wbB8
IUaz2ImRSJYEtLbNWbQqYIl4UNjp1aXgRkb70vqWaXnRf6RuEiGlAonGYXlairfZ
WhZk7Ak/r0N9ByQpWxNsezQyspoE2svvtNZKG1tiuw27+q3pVu5NWTzVFdP0+zKo
KjgJ0ZLkF6/uLT4SqAFVEKeT1MjaLZcf5rfsDR33U23xhHhuJjAfsfRt2HP+7cZK
Mep5KmuBGs58+kzuw8GXTVX7ijkM0dDmpVOQtkp6K9wwMzk8ecBYIyy/mCpe/yAI
aImF65pza8ItvIORT0qDDFkbaF75frFaFrthU5uo3AkUxeGRx1aNwagSoTOU/rFf
pb/yDBi5G3P7tOFojeEavYj5/uhcSUvb478cg69sw+7thE96JokeR+9gr6bqV1fb
5wgTuNCi9rOzvtZT/MlxVdIPOCtAy0F/AsK2rqZBfeF3sQRh3Q3xlHIZHpQtgaCh
a8CvCq1tevoLEinfMCjtWOBBic9576JlkyzYf24GgH84jkc2Oask6scWmQ2f0QxD
GPUCpsTsb8XA9L32/W5ZfRy1scAYlx8zL3ZGckdB6dY/wP96NEjDCKpGVQL4QVWR
kbj0g+Hc+zHhW///v03EnJOMOaZSrYl3+rge4HtLPb/SbP+p1bpA/bM9+2n+6RHn
biO8srzZEXpjhTDXh/XI9ePtVRYwkdqZMyLO0e9ZgO2EwSdksDcHBavotk1QtIlg
lZTTttptrspXsqVNmSSSITEYRv+65iUfXHXN/Qtiv3n6r2KfFecAv77fTQFP4HKp
m4OhNBaTHU9FRrKlojGB3FbTq03pxwreMVjL9ZWJ2mfX4CJ+kJse8pAZnJIaldaD
OFy2nCtw635scip7aGC7eAbA2OzihEve3C9Xq0/7tDhETv2T2jx93bTYdH56+cLj
IKi2ls5yAaVRaVEUWulGfhevBShvP6HrWyNJuSbeEkEde2H7dUgwZnAcIyQogMzi
OU3IIPyeV6ypqaicOmzcMP2c3Um28EZWQoASGxwMNZp2LGEOldHJrllXogRxNvoW
gT9Ah4roIIaNhZO7m/Irb06QeeYn9XSG52z++rOOCmotK3OpV/ttMynUC7+cAHH7
NyyUB1R5MNeMJF10SgbOzGd5M7kDn5Z0Gy1kAmpvJPXI2EW4EjGLrqZA9+X7COPH
LtSq17T1594nFGTix0fkQxCaZwXyUNHRtV5pc3Y8CFk9Zi2LKO+YzMEmOfGEpxdT
lKtYzBdVNYJzv5bFO3mAd1JeBMcBmudon+AjKx4pZ+QZ8dFo7BAfMeF7sD1My+EK
EWzDb91AkjlIUv9p65pEsoJMKAoMBXzoEOd2AiUhBh/xY+mxmlyfydwEzTw8/oda
lH1rmPt4rBwja85OJw6WExQ47+ItSiFSlsItYsRqWWaQTahWzUNM3mgPFLKWTfWU
Y5bfrvlePeFDdoMy50jRxHda0A5X16UwYQnmYcJbP8NHb+RM+6uYmEEJidB/+XW4
ZeCxWTI6Xi7rAmmzLQPINH3XL/25nkJ6ei1xDfmiEA8qlRzH3cv/uE8nm+M/5v9C
CGeZ5axIAG3icVaoTc6u38DRTIahLxy4XCRsK+a/7jcVT67RyR4llOOU8C/caOLI
EpsqqSvMNRqCMeQsSPP8KVLI/g1W8qK10Ij7iytTNm6noCJjfCQsbAcNW4aLR51h
M3a7vqK4h6xdgw7nXkXsOFWEU4bLcIG4I/PY3R4whfWIzGqQzx7Yo+F8clFL4CL7
BpilQVMQmCyeBYDo0qNlSHUCQBJlly+omU5sRgUlQF8awiFRvaINo2vUjrBRmmus
KbVDBb4og9I/fWAaDnB+60KqviSUVT5rrCim7eOpI8jOTHpf64kn0Fj31TmIO40M
9ImiER7BY0kTn1M+kgfuCBPPQhrOJ65Lk4bPgAm1qjfynbLWmFTYyGKmNQIgWdXv
G2ItqtZV1MLkhTmMn9wMTwhuaoFGu2HGpglVuTOqmbX11yTTacSHAIWhC2nI6S8B
xKiF3YXneXSz9zfxOD3RX1pKe/+xpTtDF27Ywvp4YWngembDDHhU/i/s5Eut7ao+
ynbNbQOUx3+mmDToOq2kL6vArhqOGdGKt6CKl1AfNS0L92VC5zLodugIApcbqj7d
OutrT66YhH9L2GBwzTaLPx3oaaQIZlPuTx3n1SA3pL8/mnn4RipDo+rTPdjdRF7R
phBw3jD+QQ3UugYoGjQDUzHlJ1vynY7OGvyCE17ds9Dx5CyMfGznDlQnMVFwhPZ7
zf0WlB+zxYGx3XRA0RH9KmdpxghnBVRkp+SV8gZ/elDeYWA0NVLTDJJFbvk2MSnw
I+vYqtcY8Ia3HUvaOkxcGYnVTjBlibVVut2SOxEt050mFAz54xoqxYyEFBX1cSN2
yYo5wvR9f4dgqxAvg9rb54Wot9R2s3Il0m1sMRbwObKfYDE6Ywzw76AYw9fT7BUE
6fCxAl1x5Ik8ThKdDx1mN6ODIOU7vpL5c9MZ+coPxL5zaMTubGFQUHJe1drf4ZtT
bYUmW3OfMDhjMt8WxaGuUTynDasgPLo3j7akV0H6/y5SaPt6QpvU9k7v6QHNS0p3
4Y8BBw6vluhi3Hd4iaY0Z+gg4m2g//dJdFQSo7DpsgbhHOb8aBM3Lgil+iJ7NIlA
mXK4DWvenaFX6Z19//ZqkcBZ8HG/RAcEjIXu+gw76vh3GY/1yEqkqt+f3EVECU+u
A3e9ZFMlJaRAHT627Ef58bq2ZcrEI6qtL7/sBV04FiYV7QFu75ePK+fMi7IVpyoV
gFigpNCV8miRf82IPZrOmY4USLRbxD27shTCRA+qwYE97SDlmZiBJ1oEmXAANcAF
n+0MdzdL6dn59uvg0NiBaTAtE/S9B0R3O9rK14boc7X/6jtITPUGO/9vycUwlOsR
3l3d7TK+EWEHGlbZP81s0diK4V643DDMX8HwJjOLVQu3L3Vwz7xKullMnGYvPynD
O6Hg2vnO+/W/9imZS+tu0Y+VD5KjfqdsNz19nV7Dwfgi2MBVpvju8bppwAS3wWNe
q+OWxMO4fopxJ8YhFtsYhygQjJRGFv3M3tMY5QyhmK2ODbx66UdJQX88QungP6z6
6izGpWyUnlbbWXIub6U0Dc3DW1O0gnb7VAMgxRwRyzDoDl222+4Y/n80TBqFV5UZ
QSh/B7WteUgBo3QildEZyp62JL+2J4z8MblImHtSehL8ue/GTnH1ZSQyEAqNLTX8
A8EVFohtO9C89l86/xDZBqGaW6HPULFD7IjMlqAIYfrQG3nS8M6XKih60JQpi3w2
ITNcs2CzUD0OCz4n8+55E92qpe4rma1ugQ9OObgWdfCa3BdQdP5nlIjdUsIQ6MsC
FOyp03PyZi8RcJxmrMBpBq+7ZfP1KYvpmFhdtzCLCMpuGtSPwRkTwmUtTibXXH2b
aqy+Z1vUsBoSltViiYDWscbAEofNhIIftB7t1rKQ+J3IaOJTueP5SjNt6B7Rpzcs
AyN+TaCXigiqqIrW7iIzODNJ+K+c6/Nt5pcZAhbkCecyDNXU3nn6klVLKuumnD0E
upy3r+1xZiBjCDYVUeXds6zk1qCGgqGvbJexXPpMZ6yJ5gD1K4qkJAHDfYKjKUqm
sIXF8yCuOCKzhbXw4ZSyKGaBajmbFc/68D8NZLrQBRBP0kXx/x1nueuGvDEpkou7
iSAh/bSzrBHuoMnt5EpTF7UqHGL3et9LD3YHXGEgSw3EyZkq1JiELFswU6H5xIeO
x/FHLmqXZYnU1qFQD14jOZeny27Dy57D3tSCROFDmu+WPTRF/UH+/cICPhd2wbTY
UBKXDsmdzc2eiIz0qJU+HUgdLz6T6VcjWYutnfy9sW1UtoT9WiCzKiY7Midue4j9
O9gUCOHcpCaN6bT0Gn5QTBKmYiBfOxQIG7wXmT+ChtUybP5zXAVdG/5i+oQkXlQq
Nuh/83BRr02fIX/gFsxBMmX/CksqrIbgLy8bEkAr88lYcRGK+VTdS/dmfUQ4QFpP
slMt8pCB50sc0Dtzjj98vdT2Yf0AqdUi1S/gBv878VwBtIoZSP6cel/2Awllsihi
u5qoM8BpSzBcj3GfpQ7rMZNIJIG8eRle2jMTNjjQJtsz0wVgrm2vybaRaJQdnueO
9Oo0tmwVIgPI5lNipizrfsjSoUU12NBgRMGZoNuFgq+3TsuXaBSdbmRvPBaFlNmS
6DrPsW/C/rNDNiu6T3fXkgcZu+jq9rxYl7JwSmnJDfSkUbPOX+h3oOOVzx3CWDkr
bEKaPXe8pMpCd01DzYDtPu/FNIyN/MvIO9ltX5ECSl1C1O7WP96YoDww4RKDOwcB
4RA+aQVMNtt7y8zkzCnDhnP7Kp8nVUgvfpCZYKCF3v364czJDEimfOPebgDi/1XR
UQlI4d+37bkqlp2A4/Y0uCkhpNBpTISZMvWsq3NJfnEh9WrE8JQwQtiKfZN9hRY/
H4GwcWwI+sdStFnqPlxsHWOy7dsr9bCh9j9OpRhPwo/8CnQBVtfzRGezW6S6q61o
Wj5BeU/LTcVwpp8eEcOjGHKnAT6nZcVGTMNtb2h2+Jim5z3lsKq/yts3cpdiT/gL
6S/F5mfZjAEkuPZfcfDe5vxhLWxperP2azWJ234iVrMjqXJWIUPqXyK/qnrN8yqJ
1hQyPt+6m8o49pb58t2pGC2ZwUYrmzuxkz6Jg2BQ1wOPV7JcnzbwVH0R9IVQgCyC
tSjAW48GWfSyr/Fer+zJAfZk0TFM8lfElgddU2rK256oBcUeHDJsdlcRB7P+49Ue
OGYAgz9ttU0lHbRf+qTR6BmgiTkiqvmJ1gLy2SI3p9EJMYMaWoy/hbJTNgWG7Yv7
RhRB40hlRg4ld7SyEdL3LVJZgHqI/7xNPwlB4fXKZ02ILdInWQ5UUZuLAkvVxKX9
8/mF5AsVE/zBpSuF6T8JnjzL5VYLleXLoSM0BIQscyOO5CU9Yztqq4g6C6r1+8of
Q83MNmZYFgu0/L8WlsDr+o7I6cjCX3I0n0hCjpUnhn5CHpqfN9JcXeXmo2v8aFQA
rjyIT2lrpETdNe8TAQZA3SVMyPb3YfACt0czdf4ty/uGY87uG3P3I0H48aohB5cc
BNSPvBiuxixmFkPZg9rHyL5YMvZsv233qrmAOqcyxutZIc2RIyGWoA7XpuhhyZoJ
FL1Na9B0UvQHqMgQll574BiGfpap7i3gCbk/RcyyqEBZQhnTdAgh/UfqJ6+n2eZD
DwlljfAkgIYiFEnOZZHlTv/xInzG9cWzUYxPmX+/LfTobBa7Wov/ICzhWUo1iF+r
82vNoFfbpmcnDvOshNw4S3vrnq6MnMFn1cBuS7gEoBX0x4cRLNFHKhBCEv0hmVYG
eIeU0eKcUeav8NZYcl+4W04xIlGeYq1xPtKQfTdim1Wy3z8WLr5kh1mxsw9YzcjO
9EpL5hZz/DZRSgrCvkwxqPCtj2dVN9gt08Ep7pbfCj3MmkYiPzo5IcUaaEjm2y33
M6If74kHICadiG1m7szkCQj7fb1nwA9xTeiYyfWW6Z1h79zuBtal/RWvJDQUWdDw
O6PKMYCQqcFTEsAMFIOC5RZafZZYBwG3keLfTwME8jWgwtyRLpy/Hlm696DFqSmR
bJx400wF9M9M4J7ZsnEZzkjf3uRDBFb18RwWaTk+oElw2XEBa8bD87+dLJVcaLEs
Z4+VWG204MUGdwLG5nIonkqQe9YKJnDWdeHf8qEmtxKnC/tmmzNPVScYk9A14Bab
hKg/iSMceHcIK5Bc3Rm0HE5O6kY+7Z374doNvPawdn+S3uRy5ijnY2yYI8g7rVXd
rA/E+Iho/++fwWgdY9B6ZGhJaToSBD551KQN+KwzDNFdpw0mGjBWfdUV8kclNWNy
z6d757HNpl8SCZ/YyAzra+MroeMPdulfRUyg2e3FcGFtq8TulbK83wOktEHvI3Ew
2kq5I4JedF+E5mlJvfY6BowtT1a6t5wRniGu2Bdfo8iMNp2F6HvV4mpDjPv40aCN
qCpWxY+/6vtXF5oQ4nxtyILATGqgbnz8HTeSvBVJoaYCEHzXhaEBdwlmveKA2Vx0
N0oAl9FVSHr0Sjf7poeCcqkuCJli6bERRE2wVQRuV6FciTG+ATcurokXzOFr1dn8
MKzsXOY6/lly71aUisX+2UfiNvkXpcI3tkQOnyVrkNUeFY+HO7ueblKigopclaXv
UAYo9n6kLW05Lrh+H08lzeQP3p/fpmX8j/vbL5jjzt78AJg+kt/z4mNxrL77NvBC
7h0rLeu721Fpdp6KF6u73R5/UIsiyimdExstale0kcO2kyxvbAKewd/owKGOzGeg
VJl0PMt2ii7gUJ7/e2nnNWDKBpUb//vvFOI7QruN6HHAgALTt/o1JbzCjCtreYwa
Ct/9xSz+y8iGthQxn7jBlDp7EMcSF0iLhzadThpPRuRRBmN7IKAWDUHws/2SpngV
nTW8Of6/9rG1sZZRYw38bItAbogmoOjlNnVVA2XszTNIQnAzYs1FnrBTtCMYwUiw
WuHtfayGn/6A/bucaCXvv0qD1/QUUOlQWayyGYvM/KY3poMi4H13hoHiiAfB54Jh
dvlvmJPG52LnAI7j91WPyD8nK6idKuA+kVd/J17/pKjGyVnp+yfkblvRkAfuXEN9
yDuNVmgXKnHORa0ylcS3a7uYhaYpac2A190p4BwdMOkVV7+kchKYZ7LuwZ5nk1/6
X/ei8Y7wyKoOFaHaQqcN/iQDOzpNYTWuG7X1vhY14Q8UBGSegRChJhJRgyB6vFyB
6DECSWa4QPfhKbKoclnJ+8hztcDTXWu+EIzcIRx8eCxmPPAiszHQobM5L1eGvaAz
HwBn9DAL9FDRIkb6ojIekDdhmmu9dIgbzm6zBD7sXJh0u+3qIOky9ZtTRAfXh+Vs
0bI72XDEE15LhR2JUc/hTKC8hEYbJ1/n0PiW9kgoL2fZoXD+hhzSC0GprwbZu0Lj
5YXYzNog2+qJeZPfCOL9fHES41e7mHKjNmnbnnWOHrVUm3XjUCVdqsYsXm4135Z8
eDxhhx3g+tTJXjNmmHFgw6o116iToeo3EEQXbKT/v4PGGMqaT9PYpAQUI/c9xmER
uY50GWH/D37h8b8/pya0jEHge68zQr+LfxpTFZ+uCihnwYLZlMQHyR4XeScIafgm
yulyly06DRdZ4DX48NOe49qIb5XjDxaxqq25mmfZoEjQdRv/EWgiHc7ATTBytwSa
UkZ/E+ZBh0YtR5Lit+hTm4WLH3+S/UCFOtACGKvfmDh3ul/xESp1s90EWaxdA3cy
//DX41lCi3l8sjfaSMJzAqOnxnUP0TmVCD6zPDm0o5G7JydVl5W1HYc2MscWlCNb
7LWKOgwwCAkvXxvTVF/m5gS9n7Q79ECejJTbHOMXMqFdXHiuWKjVOlnpBOBzw19P
WoB3jlD4VLqTB4QoyZ5MS4ZQLf8aRt2ff7z/pkGPwINmQMhM6r1SUgPEbsHo19q0
YquMYJ+UITKCIwyPG11dwBB6N5n4tAkV/Xgr5OSafc0uztolhBT35JcfYO7Uj7lt
jqVBHRyc5sZrTSbCJtugLoCpoj3qHp34xFNNJK4dq+CSqihJDajIjh0jz3D5J0D0
9Ko5nRg991bapR1f8Z3SMFBd41OfSM+eDkEKt0eLe0oq5AlTxvGweBRVi8HQqIzu
7ioCrK7lKAoyaqqR2ozTzkwlfq4yp5nwKqwPOI9/kP8nm4J3i59RLvNSdI+NCVLR
yWMOPqlTRfncBzHQQdG73gUJxU84rXEbC6J+u546BWi3CdhwtzKkwOOyTtcTsCyG
edpY0fSihDJUg4avqpJKZRyPprIK10fuHzP+Uib3oDvw6IPxtlT88lahSxURzRM1
ycX8qJjUlP8MJ1TCOGMeNzOmrvYVOb4J976+AVxzFAFJbANHT5vRXERHXwdAB+I9
DM/3MeCHEu1DfI0/pr5RaB52Ss1NTp884oGPUTYm2cutuwMJUYPyDJFFFC4z4oAL
YzRqdFCAKvT43SdsZ7s1Z/tf7NgtQazbzhsUWXknP+t2K5ovIqSQ2tl5ss5FefaY
JTIaPzMgN6WWIKpGTNfxXBLw5W6gkg60/2W1xc8ih8qsAA4j4Ys8alBSrn/F/CCe
8QOkIQ7vcfMfTkMT9V7yx/srKudikbMDyptc6etFaxs9JE0/6PNUNvcyIHQwd472
d4UOpoRvl+X9uMJ1Y74QD4JJacv9w/iDCYhtCLyswD/kHiimxx/TlvBBJu+3LFI0
4ALhW2Tq8t/2S1ZCi91+p8TLqS9YickijfTyBWrFU2AF0MBwJz7Rnh7nH/aAT0ew
WrQhngE02rJfAeAvHljP3XNaOrH3N+x1IUWHXBZx77DTB45nM7xeW1m3XSN3HPcU
om4YDm+Jw3HgqedFXulRvv8mEKU4jltPvnKlylbHsmHWry5IQwGOUOehKIEOYtVi
BHgF6erzsflIdN4p27SihNg0BshFbHs2BDIm89M1C7g4NWES3PdszcBAcnImqXdW
f0dYGUFGCCGHKs1+SqyGJ0/nRTmXUakXpVXQyWB4yifrEhdeIl3XMIsIZeeuRIBR
gXKuuLxD7eizEZc8OX69sMS6tjcZY/VxXWJneuBDTgw8p0ASLKmJk76cUZscWqX9
zP7stQAcov+KEJqjQQQFs5L/CysPQag9VMbao1G3T52yD2X/iEy/4FXeoSoZtKfs
26PDGhg5Ingzgc/Z5HB+X17M3VThIfRNk1Ot+ITa/USWsIdw90yxO6sGGkFmbqND
GY5ca6ZKG7z/XDeX0obqRjCQOIr9PBoQoW3I5nrm9pH9od0RkSKzZds3tI8UEkLt
4i6E8MFSTN+5S5ewsW5g+1J+rZGatUkvyqKEnDnBV1awQug9n3/oqS9whzcUOIXQ
mcaFfYJLWFjsRmoAjAHhvqJne8FJOCZXXp+12bhVKo4iSJzb1U7U3ObH51ykOYz+
EqI+wi5J+rGwM1AE6GgrrFHNbedYFClpInejJOc7yzQEPFvD/UHyWp5BLFLaC6zQ
ZRJaNDHVdvIuAE0XMRM5vSJNB8bL5yyJzf1MFwC07qCI3N5c6ZgVoemN1HW24vMF
/CxU4fIGeA9KeTtrDAr8dOGS2BysnZ4nHgtjUjjYGwoxigHytBrMOZG7iA+zkTMq
5Q/QgC+ZLUqjBCEv1KUNqAyEvZjlJkos1uAgwUVj8NuUoNOyAw/pfuyEFtumGG16
elYS/GCv+aXb/DgiHYYaYwZ+PxeOScBREgmmL1LUFy3BsStj6sqE5aOjrqm6V4pl
ojHuyXYH3PYNF1Yvfdkwwwu2vQYPB1oquxY7T6hFc5IKIPdqTvxIjg5UUn3z85Do
ZvTGz6FuQSx6c/W5orbpJvyaDMlIXJrQE39RA/QXCNIfT2Z0k7PbLWPFOitSWgCP
gx2pnFRwq0geU2dB+PfxF6mPbnzd03yARch/XQB5xgB5o5HkFOGyMgHdF9ReMw7A
JrTYmCeITPtLQUoaARhPKcjzR9kY3xZEr8vvs6kRUpococw0A18R6Z7Fl3RZ6EHx
zyNdYq+dIK76yisgkVnM7zMjbEyYUAR2pkQoY4XIOjH15ygR+TK+jkt0n2IUrp/U
9hFFr11rW4uRVyRFzNsaGnJjKkuK077HQDdAObMfsyP/B3VGwyFjlNmqzz0gm+kX
2ZV0N8rRvn7O8FnL55+YilRTWC0cDRDo/sK9YwTRjSVJxIB4gnQg3d/eczY1HeDP
oZKBflvQwGhPfhRofDgCOs2TfhDRwvicvRyQP367yAdYbQH7Nwl/1V65fawGeiPr
A14FiR+EsN+Yr6SarKHyMfnE1agH6NB941eUyXFTsqZDTGD4sciEWJKjVc2/yzjX
HDgFH/KS9fXygcJOb6vHiRhmA9ZCEljgyd6+syNvN5hxetHaUOUkUgQmTa/vKjr4
eQ7GpPdAht+BQn8CxvX6hgq7yzm8KROVTpVf4V0pUhaIn4Zx5/opfV6+nn3HvCXI
d3Of5pbt6aisgB73x3jfjEuX4syMY7dB9RPNN982S0Euf7tjcNqlKOyO185TrOyg
jUf4hW+o3erx4nDzKwsJaIUDRPcMneu7MS1ara9FrQ3bEqtkMZIw0xIfrbLeJ7Un
KhJ4Na0qmV6M9ZGYbiZERpwHJ9B8EkcGmXnPa9MkJw3f77IbCZMZgOCurYJSd572
qpUmSwBofNvS03udOZ5G9LkL9R6l6r6Mm9HAZqo5g+OhKW5VVm4TE6F/NgCxFzVU
Ml9okf0FQaGTdkYblEMFzEY3g483MrJd5t5SvzJteHWugjTQDH/0LjFAJByyWUCX
4oOElzwuSppJgiOY81ALDBluEDllcQLjY6hDDY5ZKITVNwcSP3TjILuyeqEryG16
SIrGS9fch3Myi7tDlc0Ab8icNQb/UnciR9XJn3LO7nJdVuqnRgA8s3dgdGNdNVgJ
6QzCwcB6uGFnI5QNbc3O2kpK1Gdf3aAD//oh9EVL57b527U1+5hvqwqvURpaQm2n
OmDdvu7VV53ZcHhz8VMXqLB5w9I+Q7kHpKWNShgMCatwCl6GPpwRIUigsn7IGKGW
S09V716i430Ie6PyKBj2stfCiGYH5bp/8VqvLmO0JdfT/Ar7ich/dHtEgg5g43QY
DSmZhYeztq/ypv6V9SL5IoKJ7LdkINd5bVHPSCZvMWuQbAj7xVEMAVBooRKs2K5I
pCaVxY7l7/8hgITJ9WoD2OgKzU4grYMmYrXaVIty9b7ezEoO5zjSA4CY0JhuHHkA
PjtxAqqrFqyq35wxbsvZwnqCQqIKyRpEVRmxbM4QBu5WGE2LCiYDnYEmCLco2thN
UaWDZsYH+gxstJdOjf71H01WXoxorpVvNzfCq2fnVFZgI6lCrEUyxJODwPu+eY7/
ixfksnHXh9U+ClG39Ijf9AYqpP+EwY4/FRyT6XBTjJGp7SWa/5xQdBuI6URbfAsk
hxKhBu5SywMG/57XQQ+wgplJXvr80L1cG3J8I1ySxuIh+2oXTElcCG868Xg5yxcW
pdu6ZkrNwHQ84rkOPOKZfq4ueZ/EOwC3zdxquEzCnNKVvL38FMCRGRB8Kk77fxeP
KGhJ0thCLiF50ok0w25JccAbBXrWzok2A4GQ6U2Jxw3SzCsBLSHm8UiTuFtCi2Hn
nDYYKVRcnzg5y2SmEqmkMw4XnQtOqR37VoDLPqaTYRAkMkVOV/vZ8DrSPEEeERpk
v6KzREoGZMjnoAouhmPnyLFutPuklOJ5mug6W9p5nXb7dXDALqELe7ub4tZvqKFo
L/FhNJ0IfWchJYgYqQMQ9dCTGtVIwHUvJbAXSQPXXf0Z0TQrhxfotFOdHZctCZyX
injSJiq27uZbJPYWE9t9z4ArYMZAvPRvtA6rBtZv8xwwq7p9sQhB2247AIXtlLkZ
TAT8M1CEH4Umv7cn5bkjGNT91Br/idhEiO6qWluxBySpecqWyR8mHFJxqg8XPwjp
HcUZBZDitTZgX/es+vmu4uoszznWO+MTAS4Q0kkKBrMZsoJIF/wwcQbjLVv7pX9m
Q52cIxBP2OuRLlHKZgLdzc3l/9ccot+zhwargQObYLPh/dzl7xB/dFs3Z5yDqvx4
B4bZln74psGwHzuPcSZWaFAT4e2MUJVEtWlzqSUVKyWRqEuzING0+Do9Tis8fTEm
GGIqSmuLfynjkMHPC3U3uy9g20UFlHnKZM4EwL2jmNwfM7+OgK6lqmR/E35UcTFt
JVeQl7dzjW/6DI6ek6ASymz/CyJWlqroNFZN6j7BMY84e0ZqU7VvYUhWnwsBczqw
/+m3w/yBYo/S5n05AXvlaIo041rOHS5s007YlaO8diGU4ZYvbHEoO3+me+dDuIdC
vCXLk0cEiwxDE6mBsCIL/yBok8XbXRVZZVEL3QvoU5dFW0+qHa7NkwYd3eDoSkbc
jP9TbWQOOHMZbkQ5CRaDky1WmrqJycI7G+Mx7u65821daHsvSyONZsH695j9iQ9g
nlOykHuPpxJJgipqsFZrl0flbiH0FuFbJOpBNrRluLkDnIT0jJSlKVyf7RJ7+eKd
Hr5YwNin9+3fTmFAz7bvG7gf8rJ5IOm10MtDvPTJgaTsNypbLn41UXlOFv9L7XGc
4m2tC+WLZu4buqvHOIVMbJTMWgJXA4wa1IKgZa9OjA3rtEaCzcf13vr3Ii58HeWn
0a9MAHr5eah5g9vVa/ncSXAdSaZn/MIurMyIQxaUfjg08AA/HnAndseZ964fxrlq
K+DfQsszhlO9g32oOGRIKdoc9r52JB+z2BD365s0xjI+MbxvM5hPpH123cxkLaHh
FfMQ1BzleQKmCdLLPT8TiWbS29DBknO5z038mXIzbJmFPwy7NsOaVG0uJKevtr4c
P1zrBjEnQ8WM1WwleQ+A8cFqTDZTxbcrPZtaeRzkL+KptcfjkI5Ni9O9tmbP18kG
S81qiqQvOjtIKSXQY2t0NKLf1wD1ZO8JVPTyr48faDHVWjXF60ajtn+U0+Pe+Z6m
9uX1aRVHwfFYNPjpdkfIGQ7LVLsm2YgS7i8nu4u9mrxzOXoaFA9aEOZGDX7SYXu8
lqdyg9k3GgqpiUE4sgU5RDriFrss8edG9wEWlFq7VWacfvF/4NPocdKG72hG1Lg5
pLZOCAfNJEvZLGFwsBplI1lpOLGTrFthZAF9HH+BlestfjPl1HpO677nma8gdL5m
yfpZifXN8uGWCjAC85NDHM42GODap7LTALAUvJHfFb4YtelNAHGNik4TbU4T1rw7
uUlsrUeCe3BTVrJwoEvUXpmK6B65QAoBuvS4XftQAzalCMWWcDFxMkn9gtU/e1Uz
MRJdrIZc5uQvwoefNY3uIQTKhGlqRUZjMVCD2M2RrnThYN+4op/kX/Q2lyHteBVH
NlO+jxmYFP/xtildlUPp5YfDRZ3QWpvt4DM6j2uJIhjQDHHLq1Ul6sLERi4RqSwb
rTVW9kqUeQ34KTVeew6eRjvZYzZs+Ojs2SUsIFGK4nGsb9YW43CILmf6kIP3XB/f
HmJtk4SYPd5gIja94Qy2K/V0cgVc5+IGVpv1ikvaRDItqgZ0REKPHeEIVS5p+hgm
6HDTK7XRXsVrGrB9xc7A0kOOPjOHgxeT1RyZ506WyKbp8x2K1z6QtUy8SkczcIzx
bdk3DLCTsPmLaf6jVDIeyopkhWEt8CZdvEO5DEzizCW+Ld0Xncck8FySLXknGoB5
hN7LTFtsMosRhzyrEqJ/0RU7DCzT7dRZ9xxw904ekkxizxy0wkrDT/C6s5dF7A5B
xVXd3U1R/UP0NFMITnUEOSdPjpzhS8ao0uYQlZhXyAwwKKT/96H07iCauvnqnZq2
0B6MXysqh/DQHmlkLUW0OWMoOuZECHxujyEkFdXWX3cnUdwaOjhw2rmwAw4iX5o1
r1YK7n1A5juHAvP3vDp5YMIdmC7I44ewbC0NL84COxVlfHqvL7dTfZRhzFiKdMmr
X9G9bv8aUI7jAb9p9rI/L8AQwb8MkYmH5AcqyT4OUydBajGtFd95Y868pF1F0CAL
qty9ofrlv5tk1yd/lXlkRSNL5KBL4K6D30HcwMMdiC4lEY6Wxs9n3KqIAseicvgw
SgBD+u9/FzbZIJXSEzPgxR51NzvMvxpqjBoiqAJ+xpxM67niaueH2IOqZ8swHCbi
Q9SQ4DTIwdXMQ0eDNzjxvKtDQp9ZSeIhBxfBhCQapjrVHevWxNwdouoOjklx6rAT
3k571gcGLM/dn/RI0SJhCHtAEn6lSQ8XD+neskn5bQA4+ESy2xpQR4/nO6k+LUyS
gcjf7XuOy1TB45OM/5RDT2yCXgY3+tngFu9I7eMnpth5YoW2cNTAALfh/Y1MAdsb
QR18A0idMeixzzysAc1EMqZtVhCchzQof+6Oayxo2DJqHCs16QbcHbxeW8BBX5TH
0N+o5FfcKcx7gdC/jCyzfvhWEjlv1l2diUvD4VDuleIEdmO3z4ZQMYCZvYw1MlRC
Sz98NkDl9y/KQ77qgZsMLqwZlw5FUetCRzQzj0Z7cBt3XhqlEyrHrjgXWH8nnoMO
qE1RvpIk9rOBpcWysgRojzkOrl5Wi9ez6dnmJAuQ/QAjwxx9XeuZbdJ8ANktQ/Xr
ayINiZgalm4z8yf/ptWco2QHGIo2X2c7Mxzg7Xst0eqG85hDDiq2kj3uk6o5QNpe
KOkaWUTMluVuTebK/0OYcfWXrs7oBVPeiZwDZDP8j7+IwccBsyfuCYhIdODkQ+rA
xzZF2TrRtbA9xA0i9dghRUwoLjGwIN3l//Vu3sjnz09p2uiqwF5visIdeO9nxZrm
R9SnTcC/1R66fAhwS3pQOraN6SUg8kZJjuwjmS58WJwydHTQr2HGaMmnAo+l4w7a
f5IDVe9dSZ6btkNHlrSNfmcUdnNPWSEEgKHB6vNRWjz4o8GkeBuK1mdRlQnD3PTR
udxqV6HKG/TexRuR7xsnBNstW45ml7M1Wh4ElSsDb6BCICNS9KSVBtJIFsU0rZuw
f6c7eRNXTKoVjeizgHfyw0Lw6NJ1zvV3qW4782cfQqe847bzUqmC8u6Z4S5KA1g2
Cow4EtGLJRtcy3zTM6hY2+tPcwcRK4VAsMep7WTVIO9UM8oNLwes55pjAe4BuvfE
3i93QH5PbTs3cjUEZDqkAC8MoClnuB0rbI6W8rbwrx39vg5yu4X9UDNutLnxORI7
fzCift6RFDFiAb6vi76mPNwQez7zI04J/sS87x3l3xv1SK9EnMJm0MI3W8hpy4CO
Tu87cN869edStrMu9eV9emcRk7I5LXRWmqjAC0Z9kCiKDfaUr6TDgGTzTW0zlCnX
dtGDrePke6+XJTtlNM/u9GKm8Aczol0dEXhwurCNTSBOGZAFHaeysOY8e6HolEFB
mnUs8BUNsupzmlJ9yTL16ktBKmESuGCMOo8ZWgIgslvrPclV6cfBt5INCEKwJm/4
8SBcf1LCbOazzoEJVfiAySR2YhXoZbshHl8kXJ9sdaLJ6+DTgw+jSHn0nHt5XiPf
zKFjry4NzsFzHGmx7WWTkskaMSJnNEnWAx6eh/qFbPlIftlZNiT3acEOyy25S+LA
+wY045yDe92gB9N4AjMdvPQetz61/746aM8IZyC0k3HfQ7JUaDnUkk5TE6neB1Wx
7q00UfbzW4NaC5lo298En4KdcNR3If6y2Nk7BKEMMsYihMWO/WTRaUA5y1C3/8fT
nEUBLM+yTxIIFPd0pUiEwVcTRvaQIuXJPgf34x4Fahcg384HBa1uS6UvcuIn/Fd0
4felTZ3D3JL3ytZvAWhbDua3I7mvFKa6xE6LnqBBueZvX0II8gOGxixdT7rWVwGo
pXRoCWp/eJ41+st00x2yQRjXEnDVWqj9+XwVfCDlIIEsQQE2x6djLcsWqxF4dYpy
m9t8D2D4tKo5mpIL+Azj4D8qe1HeBpnyxIH5KDDAQTLXU8sOK9x4KQQEGR7PXA5p
zBcsS0UZpCNlFLEsTU/IvYfcNm4+3G3ailvRcMBGNV+ZvcsKgugXjcxih4Oh3Bzb
3CULE7UnYeoHd4wFmLK2IrFpwiRaAkCNgYDkRDfn3dTht9g+H4a4EydMRgKUbV0i
uYDzYQVfehYZx12LnZ8Pw6fKG/VPrifR5pkYzr6f3MF23g58ghLUTmxj8gKZPE9b
qhuaLWDHmEwvSuX72NeNnyNSjE2ygqWLGmm1lR1Z1ImAN/xJVHNalMVKyXHki846
Zz64UZJ1ll4BBpK1Zelhn3PgL/niw65QkOYM8VsBX1JfJYVEDxkODKfNZhudgPkG
aFJ6WvCoKlJzAJqr2oAA6P4IFebOBju8LezxS0TLCtG/AUf0AHYeYkutUCbqD+hN
lZf6NcAI6fWnTR7dRtIgpD0fRkqOhbGhbJn89uaMqqM60UZWRjEVr93DBhtyJDlf
vj/+vLjN1YQgqg08k40AlKqopf235mBYY8f5tVFKZlTOawzi3Yp97Qnmmk5Pj5u8
91Asmcomj2kdAfpCe4d9cWCAae6Ek6+SCoOjJssLDpVpGh8jeou062eb+HebFav8
B0QRwFWrej+tmhmjU6af21VSXhF/zuLadDn8315DxvyF/18FVHFD6LlaK9ZKbFcG
ZvwKklLqq6iJ52yQfCehLxNyndRCuSsXxvfoeiBJ78Zo/PNKeue+F0pCim+d4kMU
ikwT/lGzsY0CQ66ArqTohDHJnUgV4Tbthr0kJJ0C5pF/ExDw9tdStyd4yKgslfqm
T9qS48mX/n5t4QTHrMCNI9rSb3rFzWb1LeKlkuCtOiI/SQygurluXGXZ8VkkxCfq
oFAQJne6lel2dX9+XHQUR5rSpSp4oTcA3ZaG7+a3ZKEkQlFtXMp6QoRPX+dpLe3m
xm4LLmnRRqY2PhWowWl9docrR/IzfdtwEV0IU8MDV3TqS5peKrRJLH5259a+byE1
cmwPdAwGEprLuHG//Z0pPp2oxjIZ4ysNPGOQCcVdzMetLeDt1rsfgGrldlcxJhvS
fyxzPxcxLTUonY0nypQGBm+v+Q2WgaFotdl20erjrOW98f4hhpEazWpvh9LH9bU/
iqFNkiJ3ubBz3vZMdIGWQDewy0fzqObFRM2q+tBCWf5jdyomw6CetQ6cNdm+lFMH
6SZzlHHTX1NCR2ODY/p0UM8q3MTIbmwSceTU7Fr7e5LwkjPACRu505gQQJoASlIg
6Q/QTcNNGzMhz6+mURsxwE86LXIstTda7rXSKuw+v2uqA1FGUexPbtRYBZ145RKu
u3pRO6ZzeynS0MrvgMxbQOxOQRqqKxl/9wnxJYa3fS5ipAO6hi/6yMSFe0Ke8R5Q
0m9Z1Z8J8DilMs5A2uEpPZT5ddkrqaq/+C6hr9z8Iri6K/EF4mDa6XOZbQvb0Mze
ab1egxH7k/lHV6RtHMRiePC8n4ng1Yb+pU0rhqRG2KYrEypl6iBHE/3F5LnBlBuS
QHR88qMHCHXSqA2/yaiYLtrI55etS6Le3g+b2ESw1Z5LcyK9XkqTOyV3g+ucARSw
oEF7BwhgUqZ3Dnqy/13Lf1XUJPTJkLKtPFtXmR5PQNEY18ZCN68UHE5oES/FhC3/
kuejqVV9HXayWYaIWBhrmu0a9Zisg2cLehHEa5FbIVXgF1z/piBhGIiK/Uch6kuj
NVHUifxtLp0uZ3jBAAOoLZgtpS3NXjkezxifgOPwaBwsyEmu6PL5PdyT5tJNyZUz
8nniJpPJPJD7CPTnuJ9LLr+F4A5wS49+bplqQZNuInMlgPd5ioy+S+r+f7Wi+t+F
61FyiWiODJ5wxvB7500c0EJ/XcF/p9xEsdU4fnM2Z3WmKR2mTAlbthDCYii4kgZy
vjYo0W2gaWCfMmyyc4d4cSrPnntldIJQp1O3FHPnGAM0wI+tgaPTq6fHYVbg1X6R
2lgMUqkJ0jhnsJmiO/W2l6SfyFKnURMozRVIxf4a6n7/p843fsAPQDymbUyRr5x2
wH/c5mZlHwi3n1BaWyuFlbT5IkWxm1cre3yquPoDLTrTrn5paCIPiikENdvp420w
Y/UfJVTJk9BcfH2RJF7Jzr4ei7tSwPW3tHPONwEMAtsNz1Ar/9H9ebitEDlI/h8W
AA3sF7rBwWG1UqL/gdkG0uavsfzfLKRaOzKGmUmi/N/nGmgPSXNotKB6RSUvj179
uXXBJUJMIA4UhoWpEWyPOj/ZGLkPzkaaUHtLGfAmwPV1zFd3vxbWJlQqMs3oYQTc
3445isL85LCOH8yamW89zFRbprOGb2Z4Wy+SDg0PmTG07vhSWEyt4TG/FBImgAaL
45VxDWzSLbwyFze7Bgq5XSAp0ObT8/X3rV11B08kXYZa8vHg0P8tacfKPU3AyAh3
PvJ/kSj9Vhu3JI98UqzkNBzdHbsDFW1HuIqr8FVqcn7QRIai/eI0+aXOzdLDL89H
iRuXySdH+rxrOSDkkj9U37FkIjzlY2lIOsYtNO6GR0digGw4w8Vd+7hzBLYM9CMQ
B65TPBWC0/nxRfsuwYwa31zJjcV3fVsDWvHXx98PKgAmALqlLt3dZDAlcAFtS9JE
JNFhIi1wMGiLmYkXGnQb7DUcJiwcEySxJDhkspCd0TT6wpDgu3mcZKEbRA8RAyy7
F36zk8UvCtmSprwxlvT4S1jktbgQjNhGL0kBnZ5QC0IWpIaE+zX3Xbg9EUAzc9Oc
vml2R6YZwiwKe7DEZiJQAP+NqdJB7TMm06BaRdQ76NON1wOIbLmoiXoBWKaGV7Sc
2jYr03kly7wCcByQt17DdZWboHa3KqsZlxYej2RH0ti7Fpne2P+MzwXsFBLDpsnz
nVzlQDdqctWI6iUnvZGSFd/eNxK76A3vgK2cbtRIF+1QCCYGyUblkSIerh0pXZ2W
jr5irt+Yt6Qbj+413mKEtpwLfgec+2BeWeUuWQKC0Lb410bCxjUBLsUwCQZenI9E
OtimJXVMgZsq4OuKhMW0fbE+c53iDyoAXf2/M2z6ERAyZVu4R3DhFN9h0sHwUZ+D
bXFwYYW7IetULq+CQ8tKUEsIb8zOyq5BRAuPYzAQYJM+JqD9Afq1jbbgbf2/Q6Yr
seQ7e2DQXXcgapaVyl66s2MwtIDe09oc1A83pvs8joNwwRU692lLbQGdXjxEuZ5x
Ib4bUx+V9aoSqYaofNmXvQ++j0X5gHDfiBXz2zq2XvDE9ObC3R/CFef/7e0nR1SM
FK/8IHpOEM6E657CP94TqkhWWQdin7gRO06fi7bNb7+D5SRn/DYiRYRPlswQRaMM
j/wlEOY/39MuoaA5Kb36GQHaXGtFS3qDrKk/GZ0/SlpW9jpq04DyJdcChkmUiZ9i
MN+J5U9GxmLVC14EkycMbujM5cuKbU39C5MfGe4PYSz7SCFTAshHf6qbSvJttkfU
wSpRGb+v7A4kctzdJ7b74gYffQz7/GoiWreO257afD90+66STeEDNHEAzd+cmOPb
7x3w3tEmcIJM+UspPxLJNN2CwHxhuEAoMdklxiUPu5AN+8afQqHdtVeAE9fuo4XC
W2BGQsEsDsHoIW8jL/picY2kslc8Jaif1CM7waU71uWm1lQxbXhrIGCSDc4gkAW2
GBN4+xVaOxHtNwYhat2LT8hNMBrrmk78AmP9QPiJZUfaknfEFNpM4mFwj7lm3hMZ
RWPm7M9uUFt+Ooa5ZlCrDDy13o4jt+tO3y2/ebKaM1mze/FVupujdWbaZNqNgUyR
OlFSJt8p0VIrH1Xtu4DuJeQuVw3c41NA/Z+cxM5rJLeYwPkxqozBn7rG/r0lLPZy
97s6LquUyUjv4gWt4MhywnQgE9m5disG1iwPwtocs+5G/7eKgk1Wse9aWKfYx5he
R0EW2y1Ze+rdcioiNTb6A6Y+hqBEV/pJj9SRLXwrT+dW2YpVZ5VX3pTHctLxTvkx
wq+OlfPwoxsn9jJ1a2M/IUIAA/SbCqxr3t4t7/5+iehNOV38G1ZDsKMnHAydD24P
wfcV3UBUdqH/bMMZJfQ3LDHoy836KO1RO1eLjRGeKXVUSFevBvFldKoldIUoAJC2
Q3s0CcEgPwu2KAO0PtdnUcOGAEGXW15NsXDCcdqQ9+9tnqtB6qJm6zGYl2edfm6j
8euF0YdVNDLQbQGdRkIyj5XGU/50/tAOsWVPnpEkzlaY5I4tTeTntE9t5kPMjrfL
EnFcse1Bjx+jNdijEJ7cTKTP2tj8bwHxv+C6g+KKnZ1lfU32qYIRTtkOMRDDine7
t0/OA7RPySN6QNlYRuke5nsL7BUKbo1hiwLPDl1/yJPIy5Ddp0E2WM6lbhZohEms
GLj3+x3IrqUOIEAGhP45MJ3UWjhL9fwWz5u97JhzD8Yh5C17sH/Zjba/udKgFCCA
e3G+uApRnGfHwcACMX6+T06lAIwF0EkOEO6jP78aDB1TN4U/UWa1FKRdwiEye01J
ngZqnSSF8P0jy/DPNubtNdgZpMzS9Ooxe1IaPDRj9LGBXJE9qynQsHc3BRCPXZYd
cHM7cNA9nQP/uVJlhcdMueoC8mXPzfgSX2KnqYPCGXWndbv+qqZWxQA03T01WWOu
LSHnT7IDuj4l7SKgEn5qD4uIInEGXX1inVSA9w7pPaOxVuEKIEdfC+5FeJ1D7Wdi
ilFURIHhdKzBsJl8OKAqIYQo0SdZ4n7lUX86n+YJHihlqFAdr2FgInB0OYshfDGq
hTB+OWC518MV6Cobt4qUSHmYbg2onY3wVDNkRo/JH78DAXtyVZUfO6TYPlH8Q5MQ
rqQLIJTUL2/Fk3i59tVO0NH3r/PZKyG9YDtFCk7udrubjpalfA5PVUqg2/ssO9IU
fEUJdCms3Y8V4BDXHlf3hCNnpVZ468ifFizKj3hzrtmnVMeRcJ+9GLtd3Rnwu7/w
uEY/9973ZLyFEOD/8HNRTDlFeMA5o8VfZg5scWspZsCShWfVS/++2bASmAOM7vgo
QJIQtHvOEKtI6RDZMhVI4I46uDPup1AS86PmzvDmFcaSNJwoedYS/xui3/cZ/3wP
JiMuPeA4jHe1BXqP6942nxIzw+aonxX1o41Mhxmw7K9/zQF+1UaXVbS6kpz5I+VI
g8mPmCRa0JUYJxSe/R1H6N9Bcsk19YF6q1CmzBYYeAXlkcRtcrnoZd6YKSBskvtE
gvx5Y7rrENjgyRGf7UZRh8W3314/8Wt4PR//DNhOPhSL5t2TMaMabYyuoJF34kSM
qyfUHK6Jm49qi+VB1YNPN8ZgQIaOoLH93IY5FrbuzzilHQTrxayib0mwbSAc7OGG
UYskYCbDnHP9ZbON5YLHwtk0YbUmkkxxGF0Uo2VEqB/bRK1Hkzm1FlNre9LvgEQy
wkGEbcA8VuTy5SVnSlP6NTfQq0UzRp0+vE2Mi+XTvEMRblxNAJTTLH3gaovwaUzc
4tsVYcb+h2+Da/O4MBAehKQps1GWrUn3V/qfPEC+yly6BEaEgTpLrLc3Em2SXO1F
f/XyGr8ytOnWkMGQe06YhBZrdkhoylH8DWLsVKFzuqGVXn+7BQ+NeqmOLZtwIOA8
nh/Wk9aCmKojuJosLtOwz20nQlOpP2i5vPWlRZL13G2Zxb3TtPA96P0UPX8oWXqa
REplo5Ax3kOdC0FjhFYKXci+KisXdD9LmaeR/tPP2FZBJqM4KiS2qZVhKERzZf1x
4/YgS6jlEjVO/+snvJ2xXE5R48hvJcySXbbKIZ1D8vo1/JY6byXLagEQELbIxX/t
oBVNfnVFZL/qPa/XpEbdAtUlc1tlh4qCycWlJoFW2ooLcTtmsxlSLE8N/TKudtnt
t6earBvXrsCf0rqru0NaebXHsNAKfG4g7ozIa/eKvPLvbRd7EuCl1wx3gy2cXmSE
pq56KJghG53rtEmjBb6k0XA++mgiNGy3ELpQV8oTvPXegsYoj1oKzEMQPI7jJJ/q
rbFOgaX1H8zrYkBXI1f79t4ohGfCvybF+I1JWo2I3Q6VLtLtTgrwjbWyp2U+7HUN
AnxFWHDCIy2SacH2tmH+3MdeiYmF9J40TBpoRAN369wuWAd6UwSPY/PyyHDghw8j
wwcJysoRs+nPPZMLyqqK8/GwO+PnC+9Ock81FGlpQFq83z+4+9XhGE0NslDS1Tsv
BW/r0uSrm1+OtTNOm1rt7TX6Q5t2mIUX/qUEeMnxILwH7SaM3HbQH5DMQHfULRQ8
jhW/cPyRv1HptUpnLiWQdY7aamVkYqQWQ4XRQmy3oNfQXDYS8y3nli+LEF/QdQut
m20KxgNVqX5//0u+NDHHFyAnd9fhbTyzK2GXhQvSufigULZ0H3oqag3jgEWcg/jo
7onDpf0RW1BcXWqz4xwq5/goaj5gnCtSA20nTDMA0/os2G/lq+eIqKEmfgVAj964
oFpjAV2EceSy8qfX1zVPkEBSX1Hrf9gCJ0tLefyygqK3JRl5niGSspBdrF9vvsk+
2JaPJX87DBGnLl2xvc8q5VC55oHWwJvRapcQc+tTK0mXfc7pShQ29+LZTZiKJhth
nH98Enf0U2V2I8d+XqI/KNOEHyRtodxB/xzOS/iAYGzJCtbdasWJCIYIjZeUEArE
taogvTPEQyzy8VPWVp8sDB8GOXSH6CnqTk+47MHUgYBhCzbsPeEVzw9qtNwzcO6j
YhuJiMjxKfcqjWZjN23Ms1viWNYS6TzFRitFyZiWc64sznCkvfupb+u6/D+4etLq
uMPE4coaTwaqLKoMYC+mMPp5kfN/NIBgdZlF9Fos3PThdVPMqFggJ0QzhlPsQ78J
7RLNRfX3xkB3dotw6nsjy4i8fJBOyJrQ1FkL7Q/lAxcjWkCl7nZquLhzYiiCWKo/
EW9HViU9HRaFs0sZlj8iWmsj1/wILPdGDFnTfINuLpry9cYPDJxAdlxZSu562v2P
Y3w/IHLeOPStPXwPBW6lRqZ/rEDD/OnvDfRaEBNmpEujIqJIn5Ck28GaJAuBPZAe
DFTyL4/KX3OSCM1gur8u4s5jlTS6qL+GwCoLZo0shyUftDqLzXSH8fMwrNywtV5y
K5L6YQVMAZ/24wQSHznFGimlXLw9BeFuMp5PDA99FskDm5q6cL86oW6NRNEQQ6G6
EtTVAV4P3YVEC40XV8AU5l5cp7HXedESAgKtz2nQLaeoK5KdsODKUEHNuPX7z20j
tJTAwdHxdIKOg4L52o2QjxDYu4dBrdVwvehgmdbqrunVRUNbKcGkIde/jlXyM/iy
4rfirMWgzUqIC/ZAZawv4BdeYznfWqTfM2x4YdWGyzOcqrY6TwznXD+otoa6Q02R
Lr8jB9O3p5fEc3mJeZANrPch2+4h4ivaTVZBeI5xpq2BRwUbECZqMh3rUknr0t8W
TZXhVEriBUx295Et2Sw4a6kte5lqgsmm+D0t+B7g5mJd64tc4djrrD+8EtaloX77
oILnyIAd23XJyAnUhP6N6Ke77iCOhTwsBLGFx4knxTRKaL5u1Fg4uUFuLfWogxJ8
Aa0QZMkAOJbXx1gAHFvgVc+bYcoYsleTATDMSnDnaXkbggMoVwGTtdPMAvyZPCwg
+L0o9ePufSSHcopw5/4iFAn8kV+hhsxnXk7RVAhhThwYV5Q1MRGWUIs6h9F4IAhr
s4pQ19/uepuxjMFkc4OHhDPlfoK+/5HLuPAHQmw4zcViJnydvVDHZMuTdf+bejj9
7CkDGsIOdZAaFzSX8xBN15q5brOasgVjAp4ZfKdIJUI70gBPVyxxCjKoujSoHveT
tXUs5vWZBIU1NGUvzp5YK3mjZxy0p+rXT0oqW5iZoTGmNFaarcxRHDOkjq62D9PF
eESypWj/Y0x3pj8L2VFApEIyfFP7eWEBbwaAdCr1WvUTEi96k+3yzAV9ZYqaRTgl
91MrAVo1aMxLnA3/5AIBdZwU6Q+Jhz1d4SCUFYxYGT8qqtvicPZRg5aAlA6vSDWl
de56gBvAL/GNT6dzbYk08WWJZ1j1eLUUEOrnDhuUeH/OJStElVsuFUC1nCRL2FS0
9D4d7VDlwSNhF9wCVJylsCTXDIllHqu1fvgxT40ikr1ZOgfXj4369fi1QBgYz4In
8VmYYV9sFGo06aVbaTOrJi1+QPdtq1giVCtawSqFBL0N7xfEHSFkgNjCgCasIVyI
vN2pHDNQXj8i0lUsRGvshA9RLlX3+XdpSDQylQEmxSi3NB99uCzPYGShq3MFO7KQ
/1ps9tqt7/ZdpdEBIAV8dUsrJ/xvGWOf1Q/gW7h2/YFyACFlBnD3hOUBh7/Oz9Yc
JlpOvo7Hl6Xv5ugstFAsLRmqOb3tQkSNP9cpuJ1Ng8Dainat23eimHX/IJ/XDEJs
OBryJpY2y3AU16QGBDUyZ3141OOnGROj3tpA1scKKDKGWXFXS9w3LPpMWAhDA9BA
Y7+Sble/IiFa9ftGhARqAPBIrKwZYrrULs3MXSXXSpVVCMww+4ak0T8kho+sJh9g
bACQo/0gwIF7wOltY34/SWjjMexRM7c9zi5dk//Asm46NYVXWerZnsNDntM4UsSD
uvxa3SLvxoCVA41lEErdXK0dwV1F/qMYucV0bZPvJHRPJMcKwbfUqXgwD51sS2UW
4me9O7Jou+Y4DfN8UpkplGgrXpj6TDmtXsCUhtZxLRk1AB7HrixzzI9bS6wl9IA+
Y6x8VhqQJp5HB1UeD4O828bkemYb12qedSVvc8vK3E1goIbMPuHFzwhIBkF5fbo7
roj7BqL9NtCEVdCv08S/IqDE+pyqvCs8XRNAVKv/FnJ3AJFkqSuGE+SE+MFHPnog
1L4VdFmNQ/ZYg7kEs3HzMv0AoBBe5t6k3cga4BrZ9fN0PbPkzrL7Wii1RugyW52D
aLscYse/YbgWQhdEh56xP7uS+aXdZ1vE4BTjZSG1LfHDiHDBiVUaQSxGPhoPE9wE
I7FI8yw4ixzmzEXyPgkdFVR96jiTHWmRJk8mmIQfI8ZVtkMcykNWHWabQcnc8/RV
wD7n1RrXbLt0rXkPhIYQhkgTgghoBEqWeXDvCsR9UrzQam9/TLwvOAgBMbfDdfzt
9wwagrdB4Mhy5iFBTEGu0ZEvGnlbid7EemweO14GUgW/l3CMjZAR4V+nVUbfStk8
DkhzOiespTAezKjLCU1fk3cLYKdxG+Ulh7Ap/YkG/Nx08BVTSp+0kggrJwj4uMFS
dISBOJTR25LZ/KKrTm+LwLVfqUwDnYtcKh+PYomi6REWqUAifFWhDbt2hZEILWdY
z57QuiiCX5bLe2zXN53ni+189tFtX4B0WccBOIspDCUhGkeHTzdqKgAEeCHjUTiF
QOqCfrTBp5aijhGgugJE9caIx3m6VVQDjP48deurZMnh4e9xldXqkFKVGGrQWuZE
35D8b6MErpa6NCntjoHDdz0JzutEwFzJyUTOE6ls75wi2YI2eQ/OK3Q7JRJ8lTCU
d1woOvU3zh/f2wohsd7Kx9kXuuP5QgcoksAn5+hSixsnu+eVSlBdj2Q40SepaaaS
K3VA7g27bVvScXTTZr6J1nm8VfKN2sPGsnijwtkTwnKgL8ovE0sjzWce8lh3YaNi
nAbPASjcM3nd2WekxbrimvDlL5vF7ZGMnzD43Si/qj7/+Br9aadOblVln714pAqe
s8QB0OouEhUbH3i9inmI2sPJ3nDRGUUo/YPtSA6NRj6u9Ng1wnh4LhwyGLOne9xG
Im8+0KqvqMhmZJZCSZI1C7+7TPz0M71RrWe+3X0N3tIjdPufA3sijlv0RqUfXVh2
icfBRm4w1x3ofjFvnaFqQNw364KOLMP49qPIgn0YkvaHNcpq4qWfSe8w7kaSoJvb
W9IRJeI1QZ2+SKsyhAdoaDoFc8cNxBPDoiPhoTZ6q8Kq8pDXqsluhzeAWfn3wpZ2
sMyubJ1tADZkCaC8y/r6JmyPF2kIALobS1bJQoR4Ao6uLr0VQQmIY2i5kzIzEWMx
8Yt9ryCIcv5lyvxXyH1Jt4JPiiUhfQmSvuw+g6hVOJ7O325wvtRWeg2qflcA8CSi
SvwxwKg7l5CEk2Awyw1FzvlDqJupZRXrA7KEYJnwsVyBXprFkyYS4vnKKbZOljRe
mh0yXzFpRdGdZoeJtOEfGJgilgJRTH8Qjzni5JZP8ZmtK7uv4Dp3VVGSV05H3/J4
1vYOp2heTDsAc0QGHhEL/ldBxsfy1URsZdVi2EDX+bA06Gt6iQY/mgdwQp+RCU8G
mYQkFIZVL0w28YVve4HeMKTqRfBiEY260H+uWgqVNpeihMppMPaHgqa2toGLFRFn
T8flb+fjr007hl81cS+JSXuY9WifhQtEApgfK8fjHeE2w3Jhctbx20WYgqbrlekG
KT0tEcoEUJsNxwzi8uhHbcymDpUjk2sbhijnN0K+wyNmh8v24aW3aTSOrOJwbmqt
XWm8ehqbM/ip91D198149IlZHu/BGe0HJj7r7IlXMvg85JQYlN5/dPlIUvplBl+Z
mH5FGY0rgHLceLwgbs1PQWxowvW3ZRLnROE2TFuDwgNdt1b7ZuY56KDvmX+DogtV
zG/lLUh1XnDSmpY8fTSWcx2KzRLByfF2XSUocIoSrcXp5GcIkjuUPxeSDpffm/Ta
IE22mqwx068YzRySom1WoQr6bbUGZlHGUFwEOnyBy1P2y/nc10RiMXKmTIGj47Fu
tVipBtkW11tqorkNLpzbYDxS1khm2f2Bps5RsPa6+doqzFx3ihJRnf5KbqpHurB+
1HMt/Wr7rWSgUGFH3skRCn+2LhtTduOEXJyJMLS+d11/Hrv9YJavUf4Ah55I6n9A
M5iBuH6ewk33ZoLp9VdT4sH/Bnd74Pdeos1nElVtW2KvcE6ATOdewiWgMIVEQDxy
3uIwjpIoeMJdfZarfLcApVohBduTmQsKbPoxAcx2CwHHJLwaeRmgG0UBO4XZHwnJ
D8p7WZKgPApYYALsUFHSeVrqdOVPfbuXZUl1gSC+vLCD6uSmLAAsWRn9k6bOPE7A
nvGdcw5Dwa8huLhSz0oLyk/qL8mz1ru+iHCAkNGMRE9xEBUO/JWWoJq28es0yBzU
oInWrElOe3gBxc6At6qF5VWKf2WoTpGxwSfgL0iXtzSaLc01ed+mw7mvFQSUjuA5
hRcdSeq2WeJrTAQz/H3P8xbCPjAfGvkcPm+vunmjCGcleXtnsgzw+rLRjSjB9y0B
rZxDHn6UIebr2oSV4+vOszq66hUCc26xGzQZ7+1noiI8194QrofZGisponkK6CxP
TZqk+X1QtygZyuxFjM875N6XBcWSJNv9rAk2/pElDkCSLkwwmdm5FVehHqNzIOVj
UWiq+4e4weL6qHcmjYBw04FvETXrKe5HFGCsXH8RHj5Yq3wvvFQS+jMxXxy9lMdU
cAEoS5XIS92fUlMODcuE9AS7vrKav5nRCamlDLNvRyDKsG1V6uij1fcsuPDRqfPQ
Hfsf7dbffcEJDqheCaK3xxBI9uHDSxW0gqqPw1sROgziIca8A0K0unQz5LloCxNf
mT6UDcHQDJ8LYi1ojDklFBLbXPze4F9RIMNmIpGIa/1Yzw9eGPHQcvoeJuyMHEgv
+mKWWnDgeilTY9+V0QpDct46xFGr87M07fRjNdvPIbtfEbNIASnbZvpesdEsJGZP
vjiJ7b5vv125/GQnXRMcf0DVcUY+98K8q+eqW1b6WHQ46QyvhmTRW/nECxPN0BxI
RERhVIQb8JzlTcIPLu6BvPKOkWigrfz6/964r3e1iao7dLxW6jczmJrS5O7EwaXw
ikyQ06k9sxhMGn1NBjFmB+6ktStoxzKj78xcaCkhRA1S1tlP9WjDAWZW6OdXQ6RV
A1wzeF6hTNwTr3cOsnIyt7XAYsGnkVkLEZekUvFZ0tiAFSymALc4WWAyhoATRYJf
lRZWOKDHaIZRCLuwtakohC8YXaRgK+VmhslRrUElrfYQZpaLRZgVea4ab010YqhH
2ikzgn2x2aW/KSLOtw/w5CVd82KAtLbg+hVAqO1cFIov/qeWxdxZsmPJHVsOjRON
8olPzRCHX+4ram4zXbS1e3qUFnqLRgxlDHLRvqWkFZXVeevznblksQItbAKt/oCu
TXAcNjXJ9FOhEoCMEUkolURvaR87F3sWlWmDaU0hEN3hGkYNGUE7tddu8jnGv56B
60ZVp1tNDZp4ewPp60PlRE5xtwXirR11dUAKn08DvuZ07tscunM6MxjixGokdLev
jkIH8Dm10OgBnmKZnTHNazomIsgorUZiKd4rq6yk2XD8ZJOpIPs3dtM6FXSIg9cF
BnvigVzMWSPzLnhikapen0cZNIzdUWQVvUKp/gTmCjOdYXDig16HV/bNUpmLxiCl
QM5TWPl+yb1vyh/AbmpO7NMnU7uzOpdw3WZVoMGszLqr78Qw9Sej7zHHBxkCYJot
XYCWmERFKNmPPA+pqlkueUSsexhPbEoogPARHzsqMsjmA6EY/RS44h7nxnpPcKr5
3x5YZLooPVwFVDzu9Z635vy74cABABB5n5MGHuscozzAGgKBarSydUKVpdTx1t0/
YCFmSo8WVYxlSDjr1ODyMQhONSsQiOP6SdwGVBtaP9Fo58zsuIhBze/I/Ou8kDWo
EqER+I0gkMs1P9k+UvBndP82tcO7HwRLBsvacx1zbrnGfCMFoxSIGCgI4vlVwbjv
R/5/0zutPVbof/Lmy3rMNTWQAMC970l7br6wLwfW/J03A72gz9ZJjZvnAkP4sl1N
WDTq8Yk8QBg6aaN65tvHb0IWqGJmMMI/9WWVexZ873IiytP0Exg9ruRerdFaHgXc
VOC6vh8nTmhkeedEHEJHe3Bb9j0x31ps5ea+hjeudCKnoQHpMRIiZvtdhnBSIGl3
m4uTIu7qDw/GYs3cxMD2fjfLpU2z+c9OGtI0JRwCP2K4YRjvy9QVZVXAyWi8kaGZ
G5R7ZRw5Iq42iTwXxMVbpypY6piWL4PWPd5EZfCa74mExufnGFYsebyGDEaoP8LJ
5FP6CD+jR1ltY+eGpYnV4TBvyoAxAcEqSBkHjKFK55lZWxT04Y9S5NEZhkJZwdR3
BoU2igM+xBie2wlSEuazag/JZIjy3QOdPm+H2rhZV/91lKOapz8fPiBawzr2Buze
db4FXMCX1OT+8FWfdk9ga6BWuRBWQGZDAEtPVRVI+9J2Xhro/Xj3nzF3H15mIlsb
ACGalyrJNp4PiyXDPBEGO3QWlxylBX/zyDkkZc010sm+XedJmYHPc1F9lJYnTOPH
rBzwEDjpnhFc5FTdD3Zi/GrgOPjS7Fibi2N/bj9hLmdYscMrXnJWgVCTtYcciEro
zWZJuzcmIOHugDilJ6HVwBL1dyrgbuBhZRZsH/5W1RuofKA+fhKuE6y1hfonfKdv
f0nrMf5AhnXQecLoe8/VrBouL9FqREc/jD3aJjMh17GZ62b1NQSSXmksocu72vGC
N7b+3ZTAL5ZuzTCA/C80XopIt9uxmMJ2ISH+Yjwk0L9andGhCLVGIOfIGu2TlmFe
3lpGLlRUXPHaJv8x6Vm60RBV+JA8gjuo+FsS6k7DujpJZQaMj0j0r9KEGT6VBJje
OYkSyiQIIrVNNM38lpdIhZbt9CapgMmkwPOXIpt26ShC2O2k6jL9tByqszph9N3m
VVJMjC2P0GBkj9KX/pyA40hT0wGtKnqe23nQvTAg/59fQUA1frYSdnQw8RDGHsr5
WgKMr63p6cgRSYiWVyNZjl/ZGKNZmF/W8WgXgqAgJp2NHQtWu5lycszpfcYLX1KF
878000s4y9x50+j3tyzI1M7k2Gq11e2kh5Mb+XmD2g2zFtnc7GwlLgxD/MIlCVga
eDE9UicoKppKP+hzgmcPK61j1RwwYfvkxySthgsYXqHWGO11fbkguwc5+2PkHrFW
iYUyNeGNT9pUNqKEACQdsKL7Dscyt9MUOVA8pfPKHyCX/szzwfYa2XwYLjj/rZsK
yB3siWzSTI990dC08TYaa88sji59OT05bHJZ67LicDxBa2mdta3Sc4GecyfKcW8p
VtfTIIrDK9MhjAmrCLwBFopZP/vmGytt48w8zr0AA/WnxwiKniYsqZoqrCAwFTfB
2mr7fOpvX3kIOvAnQXpy0imOqNp4DrA+g284/XX3tOqFGKyAkNP6IEiK8t4VIzyG
HHTtw3qz5H+AlC0i81ChZgPCw4f9WTrQNUWHDOT9Dlir7poRd5iC9ZcpsR9wdsU+
GpL3katEnY6PFlDmixyb428DI796ZjypFtFb7EDjghmFKEI4gA8ZGBv1n6Q+sIMj
VhaLd26DDEnUPvw3UNPTj3cnzsm8HHrx0BOfJLPZ2OVQrQ+M3S7ac9WC94hRhioB
i0X6JmracU94DObrowQS0vx2SguUBYIy/HQEuJpgy6yyue8Yjg5/9B8vXlF5Jh/m
Ivxyt3tU5yCsh319q4AzTHqcu2Te0/b3UETQIFelWhtw2AWv4M168nDmCBUjbvww
0Xg3lX2o4kSS9OI64milanJxboukQy39r1pOs8YMvff/XGuLGgvptmfyefXAmtQ0
gqyd9YfPCUxR1PQWQSI7VCTyodQHLpoMVBteq3YYW3UPbsW4D67SkRXzkOcKhGyP
2i2kSDFcuKocP83JcfIyz+0XT3ihN2oPI7Eec5EM0HdSRW5KwT6+iNqDNcwsoQ+u
WDDw2R8eEL7bQH7kcYk6nZpp6HfLhsaEbG3eF5rYltv1HCh7/CKanEhUP7ddAI8r
wcwt0u9ZXmYq8PfVrVDGydtOymzgE3Atbiw9UXux3y9RDmENHi9eCaq/C3IFYVPa
PPgSqLMB06IugD5gAlEJPE9cuMDAIB1ou5Q1G/Xu3qbSE63wVDx0ZGmWHlBLD6lU
k6DaAktuTCzLjewILcbURiZCOOnluyGUMISB4+8QWGRhqJZLpVfgoc0BsHf847mF
NSnbm4yT95Im+j2vk1PsInms5204XwqegX7ECC9Od5Gqg1dc2w3zNb4/XmJediNI
rgufbQPAGLoYh4FdXYpRpac5vuEsOFPRfpp9J9uLl1rt3Wbk7DM1abJSSecIm6No
Duc9wz+2k18aJJptAFpdCkm9RojkE0WBPQXo98g7Ubyzxu097BJ33w7mWLKi5dTF
pEvEoCdzbBOlMFfJU+bH2XP8f1/3DbAZ8KhXteukA0zJIjRGuUfEiOWAUArcFo5U
IufxLqXJdfAmNNCfY762wWw88Tl7maEluSBKvlbKWgbRBgLH0nDD2Rpw3qmViF7l
Woy6EGgdUMNvRjCl8jkEbNsWq1ogzyhVAKx09ugZZtbDIBg+zUl5F7ZyXmtD9GjS
ekCL1thzKCWstRQGXcHREkL13HwOiOc3H6NEQYJSjcQx+BYxLYJNExfOi/NvMZsF
UYaetrDEJPjv0tTbXLCBZMwP6S9sn64yANPlaA3rYM7hZ0bzbgdqZyNrZgdIyDbQ
BhrbqpyR00xN/KKSMQzKzqfqGtQ4J784+/JjvBtLw5JmA41j9q+sabtEWt1bzihS
HCqQHp1EQSr2uyY6MeC6cQbRfgBIP4wAKTN6kZ/QQTFC0YAED//ViG9MzLncD/Kq
lo6SUtTH5jhNJE9sQpazYLPWrk9J+z149DLQE6cstKa1xJIvcK3hf4Mab8vR8opf
oANOHatB9U+WFZctuMbfb8xKdrdATDKv0TWvXZgJG7qUdnzsUPr63/06bUCt7rMc
o00l/L8pmc4Bjoe/EtPlAd0soahNlCho0gxZHrX3bk913HlaDvEijjKJT4cblT54
gBUEaILVgQ8ukOq23qSt5HVZ2zMJz1AbP8peM3AizglM2VWjvcREcfj3xRVyLoz1
0mD+FxXi8mF6LpH1lJDQ1Np6qhnY+QvnxQt7NJE/HsYVwWhBlsNO4ZlQH1YySA+w
uLwuAttSxrHy2fpAspZ1gVfFgYONXkgcsd11ZJgzEf/cpevWMxsLbmgoDmz76Jdr
HT5JVvU4woLvp6SiqAnseSenjxYztWvptXy+6MxAtLxzKfF9WfSExTau93WihzhV
ajCIJHk0YKhLeKVjJLsV1RGCCjBZqQpHL7uyA/j4hadwQ7qeWFGiuCP4NiHm0hFz
wGHf1J8IlKrDaoQcwkw0wvRNwZUGpzhDg/nWu35aKteTsOlwEf6zuNdLEdMJOkM/
lh6S53oDAZkZX0WYv0ONdl3VLWmj/UUwHeG68EPO9gJtJeb2Zl96QynY84k7hn0Y
Jd/VW3I1RvcFpVpqexhcMqbsV2k1mqGbDISJqZwMg568Rd7rLX+cP7cSgzt4nRVg
7eoW8pRyW6YZkptOz6DKONSSNjzDjRgvHECIjiijUmlhu2eTXv2LHw1GFLFQ5kSm
qt66VmLEAISLW6aFP5suNjpeppL5iPkjpgaMl01dbHTpE/HrFZG5XLZ+IZtPwPIc
qpCgMbBVrblDjA63BkD26heg5iRU0M4br/r4Ys+90k3gz3a54nxhGoehKnyFEReX
EXklpOarJ2FrGbTOuugOjUABwl93Fel3Xk4Xr/O6/7HkzR7Kq5m6VMug1XufCtmN
3b6YMXAGSQbxfqTd2DRkKs76uYyvtwlVd9w4/NUYHMbOpRgGFb2ss4A0iTiV1FPR
IScWzhruqy1cQjPFfVe7jun/IPKKNqYzz0PQJ04bWx5bB0q0cTsbIBtgVF9jZHj8
Pp10C9GhQ1IhO+B3iYx9rrTmRl5WIu2LSBrKBafjc0urKR4w8ShsU4BKpPr++mSr
Y4HMJUNJu9py9nb8W5ES7ZMHERO7ollwQpaGiorAchCN+jloDlLt0G/lBvdhiNmz
MtnyDm5TG1iEoNMt4xwoKWIEuuo4ds8zBhqHyYvw6x1urx7pr9PffNrsVb5kxvwR
Gs1kg2N0CtAIMsdR42trqDJhWGLg3kP8DN5dMiXUwVmvpXzOyyIhCpamMFoBU/jA
zhkoY0x/J1gFJTFjul1AHktWqzI42fk/EfuPJuLMEoKECTQ0GmAddSpim0uBbLd4
g1v3oIbhrNVNaT/VR0yOfcVbJ2MwusTKfR0T7eYmc0H2zV4WCs1eJ0jgRIFD0RFR
LHBkn+rBtMaX9Ph/BmS2dFVOm3PkjI1zzDgmZ7KJGDD//drZK57yG1DSMT7FKS55
5+surhIB8scTSugWOu7evdACrT63uU8uwCSFJ020NDz/yO3LFh9SjZYZBHdzTRdE
+lSNf+2CZAVnLs7GuM70xV+4/WZcG3A0YBaD5VQyxUjYygJDYToIcoqycc9FMHTy
Ss2vFwf8SrPdAaqt5RVdYOVtHIJDrKw3XgtVZiSGFzXPwZFsVm5Mi2LWW26YRaoB
d/3/rKeeAcjbor+3u+sVeA57Tt4eqZfG0tfXNEAWmNQxhyr8YJZDWp4T81j96mbm
tbZG89vLrolMVRbSOd8e7ryUs5KA3TA454ptUQW6JlMnlPjRbtMWcIx5uRbFa7py
LDC4imSaBM6zBUXO7KvGr/K5gV64/RPDpwARDHZgl2B3oi9ELlTMnSA9CrP6CehZ
AiDhyNZGEgFVPfw4x21w9ft2MgNm5qP7C+CAY59o1H9TsVEQNPAYZLyi3YM+ZLS7
FDp0y0np6Nc8Q7GxZkromgTIPjSEKTHDBa038O1HNDTCD3L/BnxwukeH4XJSw4Mt
I8Cla9B2QTTjXjia47DbtQ0Jp6VJbdpb3bJ95tslf58yWEDcqoWh/w1h0SdBgoGs
iZHVHMPW8kifln9gml77qzfmVa6FfrXzVMFH0LUZusyjsLl2ADxV3xXDQqeQLMnT
so3G6bNUyLQ5g0CpFPeuutWw3Inw7+KbgQlIc8NdlN0hVncg5Z1bvJD5fBAcc/WP
ixb/Pwm3W5XqquXJ3xFK5rAI15THD6OT1La+la9DtU5nKI7oZ9oU3I5u39kTlKXx
5UP9H5nerZEdNe8pN09m5bQkna6pztwSpqoXbhFEKvxqozeJMyJb8u25yTNwbgm1
q42YjcHig6U1bkQy6186aR+jygLBKC8HAr1/Lb2xWrQ+/r4AlGdhhvU0R3qq4Axl
NRcmBuZ2tjJtDQKFX/keVvxkwhJU+l7hEe8ni9ztfvLxCE4zs2Yf5DXdRolVBeVD
AsaXM0uNzsDF9VNBQRP80s+F8OvMO23K9+1ZbCl5NE5VQk7kEXbu8htWswVZk0zk
ywZjw1UxdcRBA64TFvdpJqv+l0e05lOJD9WFOpDRfWL0Eb4eLOHJbjz6BnC1YmyY
miC01uNqJoUOjh4SMD32ERsSUyZ4sdnQgqtVaVGPRDfD9/wJBFHreTtUOiU2ioMh
w86WdMTDx5COYdi3Bjh0IV9safM02JPLmYIR0pl14jcvFxBgVCr1vEKFuHT1bYNg
Bn8Aq1Ehdu4z3dfdlUXNNKXl94dhXyVD/eKEIZfjVvs2vT7IGs1iOdHhm//04uVb
osuF5niQSt1IlwATb2kJF2CRMAEqZWbXnDRymCCjEK00RJ/8+VnTnvaV4JGOIr3M
XeGnFKvKg5p/QHb/XPHrs4HHXFUDEYWSSHA6z4Q7LdR8hehmrVeaKnSgowzl8Fzi
gbV1hXQ8X6lfHswKtbfzMTax90SyldtrYRTsTsvosLlNQiCDdxmzWeNltoU4hgAn
zPHyuWrEJxRpDwBU/WnERbzfbEnH1ltR7wyIxUJFbQdwUSmVj/dR5HNHV+gi4sK4
M3sa38A7Nuy9el+Oqc3RfZifZ1DGeGJ734PN+qGRfWpxXphHRClXxY+ET8ywehuR
nQPfgmDDUZc8tK19f/T2yFhqwgHzq4uWooSdawQdgRB0bt5gcB+0oOHbstC7+Yq+
i/ESJqomBDhSGtEffIDK3+wpe88Jj+qKc6+I4gNyIvS5q+QUTtWjUr0N60803aLd
2AueD9oTSQ5aRhOle3nJo19QjLSS1GikuPQEiorylTOzICVl/YZ8C/UzP+0QKt22
Ct31Cpo5K+la4CZEUWhgMK0MW02hjE2SPS/WNU9PnXMP91H9Mjs3osAZDRWn0IHX
LvjNzHAqX1mFgw6wYAQ/28Z7F+0iD/YnPQieqbgyJxrNRF1HqIWfiXczudH9bI/T
/vBr6r6qNzfrRz5HQF4xoBVjp8Hioy1Q3JT+FxABa2RRt1s47gjTF9wlzG4Zc7KV
dY8KfeRRyL0Qw4vt7I5otTFM3OTSFJ9Ds9HHNB4QSJWBlo1aEHUlsoWgwEn3wwoY
qsM1aYHmRuy1qkVjwQ8+uxIuhHvarhQkcn+nuXf400dR9Jq9a/lOp8B08NtZYXvs
/FyNSnkqlL7pBsqtucOwxaJNXs/vzgQ/kzpwINKjF0tEKUxsxo/dnfDhTp/t59Es
j2gaPrszUwWRu0e78rOxsT/QsgI/hCxLFZPzpGVoA30HK79uihII/LNvSV3vs7XB
qeAjVZ784gw14lWL0wXtANltaJWA6+wG0TO6hA+G6xVnB3UOjRTDWwh/f6xjiEiF
5P8AmHleJQp1x8Pwg24eR3sbdBGl7x3NCu3CTKbXl26Co+IKhlvNyuoL3EX0lF18
FbKnzMV7r5OLcfjDESINx2BWkDxezJIqXePlsNyY3CM+TpvH/89RriUDcLElIjZB
NkRMdmZTdLUd+E9roIt6Lh4nYxSgw7rUywJAeXqFOeXf3+UUQkWKsmsPy5H31b40
nPht5a8fFbjZqzQBx5y9eswt8qqK7DH357b1M+gnC5E2RLekX5/mu+ofNZ5wA/D/
8prBkI1DeIWCK138wkvZsq9ovt+vkOHoMR92yQOGnyIKCdUuTkZmKllKoA0GFBzF
ajp4wugsxkjNghXWX1LsK/Du9nj/bKH9kkzeQ46yobFnzahvoYiHsMuFi8p6Hm7V
aHjM0OzOWy6+70u2IgSRPiQKtm9hJv+Ph4YNEl+m31DXoYI1WXNmV7yUlAhEwYDX
evp301KqV6Kk8wuOhUgI/GLIlNWockJnqx68XfHKfPQaIDO2UwPz9C+b/Umx1Y3b
FeqkiP7D1HCcqstFOLiFrZdG+iYNB5aW8VHv+FZLv9hVdnjeiw85na9eNpr2FXOP
b1G6wE7hsyxVG29zJl9A2Ogb97vz6FU93kxFIhb6w/P82c1vOCocceKguyBELmeU
icx1++ZAwfiuU7mP/g7cWSMvtsULb3Ji3uhe7dmj23xsUOTxfl1Tp/JO0gScYuO7
amyU6mZ4tpWwwf75IGJbglYHYWJ50YiW9ZbS0FYIkZ/AEqVhayKcn6IZU2T3Q805
lTRQSU2xprQl7VBLpnTGzb4udjwzluRNVz7j+ENai16tlN5r4sPA0XIYeoRbyUwV
MbLvcO+DtqDjWGgRn5KEFiHq9heZLkN7yixleA+UOWX44aOvqsWubLVkanyitfay
zVUdrL1CxFwPbLSsqTtw6ADcC/H46PSraLafSeKMgj8nzX5JprAcqMPl967PlJvD
OaAGTe2xMr7REqu8XjQav7azuohY2gKJd8rbSH3gL9G36uw62OjTlRqqxe4DvTl0
kkVzmF5mzwGCfFYUsP4FjRoGhtE+ZepneaNY1Eb9CARZKhHHee/uRTfWW8b1VYu+
CTJUQEgPV6sCmwlOnBZuXzLBw9TQS7nEZA33+KZAhuT7aVS02Sv2xM7p1lMNPt9k
vNwkX2hKYazCI5C5blih8Z9C2nexnis8aPGRocOeOkWbRL2vgULXeL97n3RLhRR2
ek/ctoxBBnGhGWMCnFU64tnv35mlsvdl3PfAeYajjqccEjI+th52eJS7S+y3BjkI
L3N8tzSP+XrzbjdVelVoDRwteUCfMFMWcZyXpkUTlliMDyaofR887h4WGWnA9jYq
bf76Yi8TAD994Gjw9ChAwTRXLXvmwPm81yJYDVm4rbfEIowwhv5fTXflTR48bVBt
C3sD4gv8ZFteTttqbFGxmjc3up6YqYg5OQRBBwIfi4ooyRvsVdWcXekwGKH3ZJ4w
gMwALm9hAb5lTKE8U/KcdsPgaIA7pFmfyJup5ZEqNBiASRUuDWaMbAg8IGnnopKw
tmG2kqB4s2G3iYvPRZV06Ok6yxhpe2xGMgGiYllfpy8XUjRJoNGELE454HregPiu
BtGByDsXV+vNkAAyVug/IJwOrZDB7KI7ZU4Sm2FRZeeO0L6mrF6C3kL/RL4NHq+u
d0Bhwnm13EnGBQsPrmsCqJXSDDF5DnVBYltzICuGTQSvkpG9BX461Wbw8X/qH/g7
EMB3G43MbR2GVwDKSBKjdA9KTmURUHxJd8ijUT/aek3SVYOG/3covtxBu5SXA6ak
NtkJuHO1hhW1o64CxjsP9OBE5P0kmowHk8rrxZAfJyHAn94u7KvLtMTHjm/clgmn
zVPd1D4pOqCMHVpEgtKRH8emtwyAsXFym2yd7klLHsl3NLn6+1Sk5U0wL1sAJB9Z
zck161sGLkux39W0iW2Z3+ofLivV/h7URv2JUYLzAWGB9GQjQjw5bJVgA8oDvpmP
kgUEfEb/o6gzjb1HVFxx9VLqsbFmFCJwSPwECI/bgDXXu7x1qPG38+SePzWV/DVz
pWTtWnGYTMHlV/W0cX6YIl2N6DEv1+9Cn0nB57A8N9pky0JFBa5IBNFbhjFu+xXw
8XXBWBeFVHN5ws/NI4uwzaPRH/UnNihLkmEQedRq3fDRokdjo9/UY/dneoWJpEWf
JOi4Pz+81b+HDM83wBwhgLTvd/aIACz3K6IGzbxWrpyB+RcMfPY3WMV9KRd1UVc+
BbtNwQToV6rKlAqbQMNLDjtfW0/XZtR5uKKXTpU8Kiaq+i7dV3JVyM82aXgTVaNq
QVHp8y4jft5OcsqZ9hLpQNd0ncohbVO7peEg1NTZijkaN0fkomO29Pa8PbD/hRF4
SarIAkXcY685gtqXsEtl2XzgFE5e82nDVz4ksZtqhKCUH7whxjKGE6PAX5jRZjB1
3HXOQiwgxPSMjFa3S+HsRq0/44BnBp0zuTYD6gaV5EpMzukAQfxkX2qdstEwZkiU
DAry3tf+VvISwmginTyeaF63srerPklgIzsmDXuS94bxN4cfxeCaK4L9nTcTRLRI
DBwR0UCpWsgXYSJ+Mn7YJ9q6O6F/MO4Raeg7dZnzNCgPePJQ/Q71ceWJBtvSlEPC
fTXRFBiOOpXxnzT+cgdJdSjQh5LvGyLFr7uU3b43cszfMM38AIWrKxl5669FFu58
j08NnRFbe3EyPjqn5n0CGuyKdxyMTiLIuasU6FWqGN76wdaiQttj5x4oez5hxi63
zCKh5cc24jBkLuBhxvcwTrqLHyp9+uyyf3a9tS842o2EIEjNzhh+apArHknEnfu1
JDJdCv2pO/7ejN5UUqT/ToGUyLwoXXb8/mz2PVFEUEcSPzNo1LC/vXbhAXjW+b4Q
j9Q20Xesazz7Vv+4Eeu6Iedxc15S8NsLdGrbQCBnp9lzgUteOGKhlScq48udwlY2
Ii1DbkjyMBGM2Fwyn4yE2+8X9cfee3L42zus6kBH789RCvYtoZqFj/fR64We++ca
XURm8U4E7oRfJgueTtb1p+ycOdXKYiZq+psA8z3QWdM1A4bACT07EsHzDttyPHz2
fet+On6J3aI0qdbbPMdEAIHeOzDs3UcQ+wtqsgSoWSnMrveaimjSNQ8Dutc+YqAK
9qKIslo/DB++fHO+ZYht76aPuitLglnLtC9RlVLt1it/fDP0zEb1K3IhR+yLD6SK
JwNPiOnJsQmu8ndSORWvBpOHxLRB76hWggJ5HBpCqaOS3hOqEd5GUcgGpdydGylt
0heq6n5p1UlZKVU/mXg7/IXCavJ5xEsXmi8MmMvJp93wHoDPao1jiDmPVNDin/ya
+qkZiflzIcjpl8Yd8d3KdImBbwlZrxvVZcoqRvypyLT3/yvSDX9EOVaHnkMLTs6O
2QjYHLQJqajl0+OkprzWHyvSfDXnUfpN0v17JfgvC1Do63a1UbgunVkZeBHL02nQ
LM1909t3wV7sCVdsAjV/gnxTB/KBhQl5gU69KSBNDeO75qLzjtweqKr26LwQYdKm
ULrXgiAkP4IZJmoq2EuDFF+ONyFVmP0U3SzHAQCq4eoYGTGL+2yz9YMEw1uMbGJY
6WiL3B5W9AgqOn28pIVOBTPGZbRKJAQVUBOg2XA6H9PtoVpC7vE49JU4+OIP9Na+
BVEAmHQ5MFLR+B1mbijK3l9BK1m64mEeSFPRgiU7cXNL7IXGGqnO0Bc/3NchBJ0L
k7uUtTuWauxURW20peMcDrTs+m+nYbuZjl7wiSfSE4sqC7SB1Wi7u71p0msHXolV
RChqTTSBtTHt+IPxLzic7sT2U7REjSJvvJa+v4IbVhAVYFxrx9leKW5I82fmT7p1
mDp9zB6JFsgVBqzJbNryi0gGMq7v1hSgsXaZxC3i4hsnUnkbyuX5+FOU8wlyjowU
JrekuxjX5ggd6s82D+jExoRuV4zEAYchBHk94U49eMW/ES44dCwfo7j+4dumZLyA
ceN8hchWciMRJSTFe5bM0ExhsX/O0hPKz/6OBrJL/Sf4tSdBrmgKUcchytRUJgqh
+0UlS0Wr1Ys5W0v8OKsDYzxDPSlSg1qhWWPUqS6XpBnBRtpr66kAZr/nIojeDIMt
2ftKtJ4t0BNcNwjuGkEXTucrxFLjjM8l0jnmdPnSr2icVHRo/gG4EiERnKL1etxT
RI4/HMyUcI+/u7rnWsnUCotH0mAHG1ixgfZX08JKKS8KgvS1YAJn+qnoZRuW+RXA
56iIS1s9gYemTCZVyQYfX2qeyfBz4uNNv34vExTAHoAbsCFEYprHFTWZOs0S7JCE
qij5OPnNcknD/lgehyZfugE1SjpHk/TSUXmCJENlNet/G2UdT2ZQZrjR/poRUovd
AEitoeRyuFDv+G3aaZ6RTzhfnDltPG6adTiO6uFGLj5wum2nz13MLcRoKd/1115S
1Xpo61UNxF47C/y45oAp2FvYLJ/R7X+W18DgZ78X6ugLka+uS7sUayX8xC68Aob+
W9SbI++ZOhU6JpLtNpyy0J61oCQCC9oYKyJTrt6v0CO8SoxWywMk4kVoa7M2CmmM
gBIj1iGDNwpBqaoIQ5VdMV+VNwU9RaifJcJzvtFQYtPoxhV3p/9x/STYO8wBstrZ
5/UkM6AqVhNzP+LXFdZ3z0MHT10Z9NXfWJoCiEqPx3MDQUlhoS3qfzZm77XO2XJH
WU5KSo7yB5CbJDDqnJb/tP1mN6iv4gdmBk2QQmKQ/OtuakCoUCE0mLPxB5MZo0W0
YHTPObhxVC2fAziDfk0/53vzbBQ1s2i30VxPUrV56tw+/yHthfRWozY7G5G1YQDs
+gDw0lP1NhBJ3sxs0BIvS78MZlRhmCsirEEKlGQqd0lac8wMHMWoSXPhMjIIMW0/
fTtpYjjeMX5kxXv8C40GbRZGlBqJU/GdyH4vue0W4oGghG3AziOq6th/qzyetuoC
JgDD0KSVso+VvJINnbl1A7qjFqdXjtGT5LYDKjCnAiZxmavq3gfvnrjHRBQAWkKq
pCmP41rKOtN2lKLFV56iB2ZpagMgVnbjKAs8MYw5bAugcR1UTC1lKrEa4+s+mB17
i67rtcDDlwbh82fOBvZeJLY3/1tnfTYxZId5vLU68dmkcBcl9rA4h6eLmcdoPjI+
Oxv+whlBBZ2MHNmMoPUHKanzQpi8w4spc4VSIA8J1t1Pq7Yr755kAyu3Qcfj2xT5
Lgc3OrPuzRmNUQQozLJiDlvFbDwB65L0vttUAyBYHZQYRou/WireauUkxFpdC4nX
xQ/maBS3yCA+GuajGDjIG+Ngo47RlL+606u4LzJCyHIcQGZ1Pb7+6Y5N78zugwQ9
G9zQw7Ti/c/aqrHBBE4XeVBPln1DDxh2mgEhUdhrSgngieQUD+PEBDiLKjleBp+c
IL6jeB4647kE2jdvhnBImeDtuvEJgTH5QKmBHLJcuLzOlnaCapv7MIiSUo/VvNyD
buxGhUVm+AE5g9mYYHPYPmlPCVLtMUsbPWRal3IIE4mG3tXkZ9nMIfONr6FES+hT
yjG+c5Mk0YOL7OHAVmvXfuffiKODgDj2iYzmvgezbGK6a/hTSQPLY1dKjYp3ME/n
hdK1tqGRDkXK+F/XCsSBlb1jKOUhCokLbs47EmRRIr9Ow2JLOOFlsaEx5GZTXcKU
gFc4A6IeBnYjA3AMjg8orksmWEAdT3hXupu+kWX2p8PK5CEJIHbj/r4d0jCPlY5R
mhX3SmhdVy/y0rI7/+zvO0B6ZHkyXpwJc6od365ECZGx4qyjm+k3ryb86OTDUsSt
tITUct/sjH3JnvRaNRb/AMEnvvD6hn+qB3PGTCSlOgvoAspwIIjJ95jbOH2FsRre
dhGh8yhmCml6kf4C8EpPpGAlMI+Jhk6HY1dyUH+XyBBLb4mVVcO6UuzLtDvxHluW
UYu7adytMzpDY1kARTvcFwJpvAb3JU722EkfMo152ODrcMZwwua5zB7AeGeaJggI
ZeVQUBDN13p0PA/zbFN6IaB2cbvYJbU/WxybPQslZH1dDK+ixaQe61f9aqFpp8vW
nnS2/7Rjix8YRQeW/fYizKlPc5/0vs0zq0l2qlXAN3mjhE/3KqpL9uODLP/5j8qU
mPSqoRyRfHA4YgGbacpYMguBxpazKHkcTpove29VNZNAdk4WW8UaaiZi045OP3Kg
qc//lizxL5EsMYe9/ypTm3XxkAaQDHV38lexDF3JUKNEUhrF9SzgYxNDRSltLtcW
Q332e8ZxoN+ujJXlW4/MxwGlL7OcbtlP5sa+Ew0rQlaAYesWKY5CZ8wf4lko9u93
YEnts2xHem/9WpXXVOpYHBQYygEZyr2l14Lq77QkgqioIClPy5WByYqGuvjjj+xz
TMtB0PcvDUlA7/hcKqJsJdR6zGmT3ADb5Sr/BHL7Ors8BK1VFBro6Nff1u++nb2F
8lO33/Xxe31mhaO9UZgUPiKEgy3lPzEf2dzpwUfgh9yoR66WwCQ9TOhRCory95b5
OuSLCrqjzQR0W+QZll25LJX/hdbAMpnmgnfH94Jc/Tqzls3nt3ed2wxs8adzoVgz
HADs7DZPP7kCaxshp/GwjHvlvutUgNMOXqOvSAHL0Aa7U2SwZM5LxwQnH+OpEAvS
5YLvgz4kR8pX9WFe0bB/TEw2MjYAMboawQbuwksuhq1kmXr2Q+V4MCTh1Vyw6s+y
JIGdtyz51swa5e2eGXlftCobu3pgD97W60+mPSscpWcp4waHkoLmM/msi4lHlCfL
ds4qBNZAbX8Y9FH8KwVYfRDx4kBJvPARLpKMZAnpG4/h6VbKPMJKs/7hjfPL5Ti/
ZIgCA9Q/XV1fvo3rvT7AivK84NmlPW01efX9RLSpKLpewudwKCTwf+nP6Ms7iTJr
JpJE2SysqNHY6VVninVlB2BHHLxB4UDyGZ68UkcbRkoZMM9tldtaUAYZq8AOwdH0
DUTgz4lmwZRCk16Z2WqFmWN4n9LtvdE5Nkd7WGCf1uphHSZgDFtgKPRO+zwQ9gZn
DMigy/r1XsyYoGLlw0cv91IPcsTF8wCYU2mjjH7+pgX6/jDYejZoZakKV2oJ8P47
MRZTw8tx93JPHbxHuJOPBmk4sc35dV1cbq0byCuZTtQ9rLjbeg30D4XF9q83UFjG
iu15h8sTdWBdo3LSbgRP33GNc/J5gO99Hwdy6Tg0ZGngypbPgB3tLxXKNltwMTVN
jIriy2LpppkdGDF+VFpF7OR2EEX5uNTHc7ednMWK4JBZ7ZH7L/lBt3Raw1XlUpxD
sZUahAvb9LlIZDVIf7qOgY+tBjwBo8S8Mi41OwY5AojNg1kJ7VsU1W5KeskKGt3K
48XrJHS8uNZe57cJmbxZDtBL0NLkXtnP/d+zl+b5VsoQkk07Gt4j0T+o7tgmuTyS
cT04of9fTnVECQwEQG3kwcY6wPOpyyu/Vluxa/L/LBjCD/mkkMU47+6v71WpzIgl
yQzKLyVLHsenz20mz8plKF+QcpyaOHzmoKeB9BX7VqOyYQJ6xS88R5TW97q6uZiC
jZBkk6fX5iQwKC1OLIRnL505YZM5VMVuxqE5eQPbcdcnogFjEVTxQ2s+h04l53Iq
ojNkq5hkJLqRbnguEvRXNKJ6NuhLKdFOCBA95B3epNXUtIsVN+lZlI047jvyPbnv
WBOjrYhXHvrcrOvlFPHcdmjjJtib179WKbbT8Az51+nO/WoePUO6olEYF3sUV45L
sIj8dKerDBlKzyfx7ACfZbOQcfa9Oi9sWr0PSBud+TX74fr4a17pGZMGY77NqRRr
cs7vQQg+XuT4uvZiHUpCra61/+EIujppUM65F3qXgY8Z58Ygx0jsDkP8xPMjipKa
tNwPNMqEp2l6B0kzTfGbqcj9ovIGkFMoFhqpCn/06tziSQVsX2B4JFQF4gI/jXMy
2Qc6JMp/oAgGs63f/e62dkrRg6hfj+5i4vx4IEtpE9Inb1IRNnpR174Qr9LYmCF/
skUTjPUQzjSL//MRiMLdrksJi+/BQ+yf/egWn0XCCuqYmkkxLY1tkNUK0FP+2IN8
7lgUpf9F63lUy4rX+QOWmU3u+pQl3UOX7J7igcYfMs5nmch6VDZUw+KQI04+7WjD
7mvnTKFBabUGFDh42bA+KbHDNscVSvfxgavMAAo4/5cVhxbzmq7mKE6ePHAD7RY1
YeWTuuc8/eiVIOq1AOD7wLfRykE6mR6GYiG6cJzszjr0WtLN65Mi6OnasxGkotIX
XRlLd62lpR01TPhu9kAYcH8XiIUYnXXy0adWTuySpkxuhCjcxh9gKN2CY2beEhNs
zZd/0tcGKAOjLkVX6fqelMl1A4rzDO7pb4gh6H2ZDAxDVWpNbqzTAuJqAgxrzflp
AOXquqdVt8RiA118JGpnhGXev4r6hKr2I/JeGYnNFlwr62bWQOviYQB0zCHdxOIk
rvhNyux5EeRSf5LENSC+HPryxQwbNnoPMZXx/yh+wfrEFg3O3EV2Cavi5ZOcTdGG
QDK2zphhiAb4e18Z9dLDqkVmLP5qQCQswzv3h9CxaA+9em6xv5WwHLM15/Acfyh1
QlnDUp8T8QjHO0gvWfnN9m1fgXk/txPYLQux5icrczzlYtnFdeTV83iGMzoDo6aK
UQyXnCjxHIRcCEM9bJ9E9w+VuUQVvX3oTLMQK27DzVR+jVwpbUpT0yOWiLjyAgJm
Y9V6wcqeXWx18vqhFUI8/iwUp7MrE1JummWmNPRUlrrJq7UA72ea5q5C2aZxE/rS
ccmGgrxhj0eRl1TdpdE9ChvdK+nMdPUyTwvSFKQeJ2DHRhZB4XIP/jzBe13lfRVA
W5jX6DmAlGH5QPdCQTOM0Spk87IhxcNefBE7kZN9rSzOMo+Ry5DWRnv83IaN5jNW
4IfUZbFA50DWEepycVnAY/GeTLrN/8DD1HnoTsE8HE+AatSUcJsOebMqLazgRcOC
Twek4dlNtuxUOgLXWiyjBkpl6T2SyGLkUv5MMGMl2oxpuqj28yScxzqeneGbUCq4
AmJn0cZWaSvMC1ygP5Ja5tJ1SLK+K6gmCHvYtorDh8Dv7/4QxSx6uFqP9TfpG6A/
DTX0VhXu2VVKpezN+UVULcHZOBr4S3yek1kOdPvC9N+KYTxTgtLvO5+9L97+lSST
cdLm0m8zCnimWGIRb0wCbEcuAV3o5OWr701V1gi0/k1HcYVb+KQ897TcHRjYSXGn
Jwb/46LBksLJSCZa5zqmOlJX8JmPdXSUSlpLLlGiv9/RTpejvwmeSuw94miP65dM
MiBxL5ASTLrh+S4wWppDhccbXw1GpH2tE8Y4DA8A010VU1cdVItzFWQq+aEY1YKs
uI5dc9sXohtRJDwuSJWpOCgRBXMb9yEV3ICUELcrNz0YW1MUE1k4GiwuPsqtvbfb
OOug0rxARv8CJxVpx0Ugz2uWpH4zhEmeLTYNcWogV+GXkAPUXs5KXrUUHJoqVjfL
jLzhe6pw0fipJtzvbNBolNQqmowqVEzh9j14uzlshLK9mVTeRmGGeYB6oK0WEH2P
+Sif7D9QuR1sBfbUuiAXrlPMGUcSuwjhrouW/VOedJvqQvNaxHuBlufINcNTD1Cj
dhnDhyEPyET3aC9HiqtCNSbzixqDqChj9XOWILbncp9otISPQxMraR6WLk+kvg0J
H5E/eCcSYo5MRyA/cmgGNRXt3Frt3L80w4Nv6ysuqhRny8YkK/42mji7hpzGbqDk
dNkLHs8d9tPJN2EKPorff9qr/QTDTcgG8GSAF1iT9ZoG8wZL2KOTOAY7X0oGlAK0
urF+ZNkVUCgt2OqOemAb9QE/WX1x2XXrsxyrnIcoCqOopXjuhlfdv+ozXJUVh1Fn
dCIpT8x4clp+DgBujAb6MpEl8FBonLl7JJFB5VfO3rZsTNyZMaPkm6d6jpHatDu9
zbohgXJOG9+YC6Ll7g2eOM0hpIy6hil2CpL8BYajrblaeKjjqcQEUYBWrGcllK+w
X7NmGEu8qtHzUqCmhLHEnG23Vs+XWeYgatbwEgE3UQSdgQ9NHgV47XomBMLg7d+f
RZU225yHAxIvd63iMs5appSKqqiOrU8i+cdUz8fpc+v2Ob85HCksbAQL+Ms/tHzJ
SWs4JqDKJGglpje6nYXmG468EpDWP4X0Iw/7IB9xqalJhFOTe/YBsvR3qZOO5NsM
sbAyxvuUGQDVnEsLEPy+JkOG1A5qX23PCA4LuWJKWb9JjGUM2QbHlANKlmY9epUZ
KFBbP3kNNwCFHMrWQL+AIkoIsQMgusVUsRGJMfavwHlw363Ji0BuI8HySbw9KRoR
w7ju0a9GGZ/udZVz4erm5f30RiWyeViKKnvLldZAqQ5Gx1/lvIFf7xxr3ehsgn22
8Of38WwJ40sGwxRP74SpkMt91t1BOuTVzL5z6yhQtjIQXIxo4FSPX0NWsdzG/74U
B64JZroza14kNKHpdE9VfPDQmfa0X7n440WwD2j2uZTdonxqfMDOmH0P1x0Z0e3c
6qR5vVIgT08Q53t5kBvsfGBxmr3Hg2rTLn1tN7CrPCEdkQyWXueqFACBlolZpuW+
vtRnuo0ZZZzXNfi6LXDdPSdhkKjslSb6wpUE+IFNj0PVjOR2UTd9IAFdoeNMnG/Y
TqjRyfndAwMbCj2IN7FtHwRaAp0G7fX8UkDjZfIo/NloCQcnjKj7peJYbS8mKxbM
Tr8PL25uQW+bFNfLzQImzQmyyu9YjaMzjeZoToSE3lbveaq1JagmaG9uWDUk1dWA
VHn4nMz2OSRqo46RGOo0gBpMQrnzQBfjK/1veNa0eQo+EQID4bTX0z7gr6f0vyCg
It2HNyw8HLk+pxP3Z3NiUqFpspMcQhJsicTR2K30qiezGOuh9yuNl0heJHr/r/ZE
fRfJAVlKiP8FB8JhYa3ataQ/EmCaVdpYa/pUI71M8jIIMk7UUq2HUzWpeQ1kzeWm
3QZ6wo8aNIVie7YGOBO2z1Owu0iZ5UFTx/Acr8MKrYiSrcFRQPWyI7VrGA3/pyQ0
q68tzknVNECfGvZFHv4gjMZFBlYIb83HNlLK0NK53DcG+v+pEoz7lvdnocmFhKKP
6h7nDEB4rOaUB7cCJ5aYeUN89d/SI3L7BflnGnYd55HaXqVf4abHaSNeXvDLpYga
eKvVn3gRJOQMpTpeV7r3gfoCVEIujoJ6AtLQmcycYc9uZi6AuKU2ZD4LxWp41EuQ
YZP9yDXNLqrhXQEh20C4Gq+916wlp7j70DhQGy+Re3cOzhgaOXYGfHaExtYv8GOU
dCHPh2Nit3xd8DrmqYHGdk876xZjoQZov9BwoIRuVRTVNVCXNu6D2DjxpgR33Gbw
SZFp8aWcgf6EwWAcHbhEoosCuxSSARRKPQWuHTQKL1FRzTfdHQaC2/B0RTaKFyz+
61fGdFu27boDiH5t8VBEaavWZpxfjI45wjYNoYWyqeL2Hlep7O08lnTtqxArLeuU
tP14AGTZjkvgtqbXqaxKxSm8Fq6oyqXs6vZWLzWxoHWvDm2S5b3rNDZaM7cvPP1A
dmtR13Y7yf7XuC/yAxMzeAbltRdfs2BjaGwvHEZuIENBd1qt2yAby6fwh77TKIic
2RDv09wg6gAoNvHvrK7J6zmgdeQEDSTvq+A9pBU3nyOpJwSl734BD2xtYqNm+DHL
X4OR0le9Onmop7IDesqUfxHl9OJUX453prsP5p3+k6VUh3mdp7Lq0W+MzrY+0MeP
iRZFtmc/KvKriXMZhPg6qpRsM3C2pPaBVRGWtOBgCiF91BsAsRAQZ7+8gIMEm6xC
jd75W/1RMOSFERJxCypq57RBE4s6d1aB5wrlLuGFAqU50IwM89kkDa9HAmWvj3fS
Ge/QH1mUAblg6zMWbRkUh7TUYslSzg0sbJ+jL8ss4QOhZRaa9CT4yFNwqhFTO0hk
YUkycGwWIa1kSwhjhX2z5QxMr7RslvHxk7iM/QHdCTrBwQAQF15Lh3DkePOw8UAu
CpLHaAFo2AITAlfvBkaNDdWv28QvOZKxgIRbeWRqTouBe5T4Kpcgr1XkmC2R36CH
Ut+lGxJVQrZJfrW9W5yWxmeoBhStKY6d8QrMR2FLdpOpS1Bx6rMAO4wvL7ONINDG
HWhDbSTC4bm8Ra4Egs1snseNVS1UnFmf9Mhc/ZjtfapHO3gqWuMVjlRikG+aJwak
dph5AABHQ1QxRN0cNs3GG2AStHH0sRwEucGmB0QJe4NwwD7SRx8o1n37IW3IHdDy
CRMlLGvBlHu1Np11BDx5wXApblZ2dS+Yhdx3MI6AR0fsbl/Tt3pEKn/bmx4KvsOX
wpMi7AvXvot+rBMZY1z+J6BDKO7XaiZYr34Ah2JhvkEA4fNzDAJjBtoVue7E0/fD
JsRdJEonPgz6FAsNFJKLWilDIsaM2R2XbMc2Jt+AwAKviNIX+Z2rGKdj5isicmX6
iQb7kEkNNR3gAkiK7TtssLq/OtPWI/g8mx6X8SaNRSfV3iByfdKLY2zFpFpzQAdZ
HRekb9sXQDOk3SLX4DRFhPEXuWuqvOIpXratupeHvYN2Iq6Fv5RFnKWj/XQWD7BO
caikLm0vVB/0srQk2tu125td70JJHBaM0ckZYK+1UGvgoq2OWPKXW/h3Ks649aJU
HoS08qrs7DgE7NA+rOQnC+fGK/jiUyi5c2jJyNC0XxQf3xkVcwi8qTlFpz6r65iK
a5dBKjo6AKeX8Z90V0gC2PqmzhINTYvBxNmRR76JWfKBYW7xhzCHJujSZPO4a18G
GFcQ6d6QlNLRWyU/Ya6vgVuvktPN/wyjsm75tasBwCl814tKndytYl3M7ZzrEfVS
L7BsD9Y7zKxLfzUuhT2W24Gm8XKhziCVis6tDZoUXoHHdPiRU44OknCFoZocqfxR
U+zo6Y408Y7igUJ/zdMSCx5d4fdrYGB76xVz9HoivgR7jz0Xg4jQlF+tZhWpsiCR
okxKOtrNk9q780f/UrH7mcg9LVpV4W4OQGUWKH63ImhTPLMiW7nmSNr29SxEruu1
rVAA1RDlw0/S5lEmSChu/6Ia0SXGOw9sTpuVoACG6KjLq7l0+98UPFpUgO6Ghe+x
ctJGDfxhyWmIIhogZWIvwZXHLxZ8xrJ6ZnLKuMjeGJD9zOChHy6o/JuSTkObrO/1
00CmMYHIHBHSBFWLTEszm4xx9FFZ9Yh3ShOI39Iog+N3CxcDtNTwLMFyBGVIn/RQ
aTCPPLxz51TSLbykNPV73rUvRXeiNLKdr/i/yJloEdj1JWjZNGFvtfvjWEKz3noB
S3vXZtmwNN5N1ypk0iq0DiGsVZ0ivy5TbizGUNJlfQIScXhoYy1io1SzDXGAqv+i
A8MZpOJvPLiaCnE8d5Gvy8xrcH9ukwGIkeQblR1USCbuBKdDpnvNT2X7K3BnRLO1
mmeaWcU5lgzM9p2KIK51WzuqWP+M0RYkuIFX1V9K9WizrZkdAj8ENWZRAkArO3UI
24Q8eZvj8RQav0SXRRRaj/zTjudMAxdz3pJLWYWmCZDeBYzolmyEs5469LvC9lmN
6mCZ7ANuLqSxQHja+1ajy5PsrGrveXvf9KCQUdrY2/OCTD1UqbaTDFQkxb3+GU44
B8O4SXs9rSGi44+Sqkbbr4zwZ3+CxbcngtvtDr73juz9zXmQca7WxC4uwgmqcJ4V
ZCKx7lnVXWL6wOeIB5ZBrwQWBhwGKr0gI2YEos7Jp4DFta2aTa0+MsLeqstgpTTZ
4fLI9BF7tX4ZXcL5eFZn/44Y5WkcpWMLG2VzVL93YILyjIC+VlQXgHyhlARM5EqS
FNRsjT35UC63A9dTcfb5eERJqSlOuettVZapOYzfxNUPqUaYu9tHeWqye8uIw5rr
cg/eC/Os7JedUZKnLPpF1watUO5RWp6JZz1c3xBUg7O/llDB8UCXckBXCrCadEx2
QnYLC9ZwJEX93EfVE2epV9+pWcAVNYWZpYnwz95SGpRuqRhbTpwJUdsPFjKcJirS
BiSDTR47ceUINHWxuYQ+1GjHqu1wvaqJi5RjzACdhEGU1ekqyJlywIkg8tBCTDJY
YBwLzF/LLaQOeQW8dei5mjkf0M5vFkARaYyMi+V1WZLtr16BZ5a0WKNQAYl/Kni2
ZElCKtYdCeE2E9Gcr0hY7wOQ8ILW2tUfu7vh2CBZX9wEIbvnUsijz8Sw6AK5j0en
uw3054ZYVAo2mFaSZRQhzeuxv3S770lXEdr4sKtOhD1xVF/r74R8nRMWSKOch7DC
XoCBJdgKe4hlNlp0UJ6F+QcDE+N57vu+mxu4biELhafEEy1gWf8ZuMdg2vbPprhP
viBpwUpFU12D6fK9WaQkYtUwLJZ6sIEYqBWOhLfwQbHftYFaoTjx7ay3jd8ELL5r
UTOgfgRRUGBXiQHSKdgfsIBMcGPwbsCAKGn7w23+P5CJDY2TWTPUXuybo39q0ZzV
g64WfLobOQktnl0hRu36SwtEhHf3aCevlpln2N0Z3rUMXqw44I2yzEZTRPosN61a
oU1uSOBZ4iWd0Dxv1+LKdcXT4ZWSHf92gsHukb5gtnutxx6rTuLTi7bphOhQPHV6
sQNzU0cO1ezxt3VuJN1MkafxvRYP0/XSyPcTzPJgkbg2tM1BI5q4TcOlhlfSHutf
lyKFJTymC2L07bz9vHYKAzklm5Xf850s4T/+ZSGFCeEVquBamkLuv0TGw/NMtVnm
FRbifVSmIug+x682SZuS9PboIIbzDGNQganbI4ACq6/JIO5mvgcIiqjpvp3omI5m
myk1CxSIrDFqnTwbotguCZAgdHrnmMwk1tkz4qCwSTEvvM2QWjeygk6Ki3NW1CWG
0259fwpfsOyLdWhUlrmuEBWxJi+3Bnq6AZpqwsgmnQJmHElXZMl4hfBg5M0SvSmQ
o/o2JCnCRJwIRFXFsxReVud+Xno/ow9cByyUBhC35iuoF8fFoAEpuk+yDVPqbMSF
DmgMtppr31IMm9ep+ELm34w5t6h+IXdATyyRhPyai/fK6P93SXzBPyJ7SpQJpfSQ
9BdnuH5H+NZi/gfFUBJAmpU2HzZsKHPa6ZCb/eTy0DRt4/F7X8AtxAdUiKzAlde3
38RV7WXMMoltUwfH4C4JbDO830LgESzZWoht8Soe+fa5fc+HSaYHJY9OYAkzWVLm
lt5Hbt6KXB3n8/64iXY6LDes+YO5vGvxjNiof7k2qxPBVVE2dqs1ICTteTgJSsaM
zXa20s72VvB8W/nx0WEIbWK+T4eLPTLzmR4ho1xVTu1jrtuP+SpA3Z4Y44s+6Bcx
QVIBsv/HRdUrZ/G1Rhf6Bq8sKEGBhFHp/SC8ahd88tYCqhwpobzcFsKgnQ8+vrVj
BdiFxFJN/ZvjZXI2/FCzdGQRhz6Jx+xJeYtPOSxzVZk/NmReYTbTAAW1JuHSgYYk
X6oX+Go0pshSci0vop/lTnsFG+USlLGZ4afLuZLAJ1bw2PmdZtEwnGoT3TCGznS7
S5rNudywsK+xuDJEVstv2A+qN40OkyFau02I2jul7TUtTd031ivdkpb5kxovM1YE
oB6rU97EAohCFe8xMHMQ1IfYh3Bj8xM84G/oBNAWBGpYciDH2wSiXpnd1xNFUocx
7v+1Vd576R0zR8WEp60lMLwd8ZEUEA9L+Eq75bmTez8p71zsefSOuzY08tHC2zd6
s0euFEx/xcBdh0CM9MdFzYb96vog8ouMbWTUyLplm5JXmCmvcky4JqMWmJIyJwK7
WbW/qBlZ4/T8POrdLf9/QrEHXEaoDgcVvrRg+dv3vonrx4xtTzANuZHdPq5RXo5H
R1J6CWQkYqyXeT6Ulrj7h3pD4oe6icPvpXnNdOP8l4K1t23lXomMDxQBBBrRjSsi
l0xpRpyXK/Sg1EuQFuWGcouJhgdTJkQUoIFYHiI+q/yEOO45NiotlVIFgZQXuGr3
NEh1KK0caNhSkhNd0/t/hjvKHes41EO7kmlb3vlPBTqKAy/kqYwrbTr1mBOKcg8p
6ze0VdAOf1YBYPD2Tz+0lZ1dy85BKzVrAQWb5ysXEUWj+SAXeGtjpRyIAt9e8e0L
4h3TwcamwD2t7NYVSsXj7OYEM+XD6C5/+HQrsKw+QjhidS7kVgkJxR/tzKdzrPzv
XELpfusrxY/hAeWaPfvdv5ZyZvsh4yV5AnuIu2Lp8J+L9HSE4kjt06IZc0t3LmB9
Z2TUxxDR+mWwX1O62Q4LuW0RMtI0w5rxPzFs4mMRYGgWVx8bsB9EGm5q6dQNN5Bj
kziGJN5KZVqLp6mgCc131b3jhkD6Ct/KjQ38raH+cJI8gYfrs4FIyIdtPwn6tLcQ
979syzVKsX5CkachYHFHyh0iG0DstQ2zfiKDr/CEBsmUQa6dNrcYvT4z4xj6jvL2
gXqyo4HRYSlgvKIDc+B76DP0CJWgdAsQ3OP9MYgMW3IqDUInq80zg4BLBgH+0RRq
Fj4p8nXnYQZcVAyfJ6KQbo0TkNh1xNCiIDY1Ey19a6J4IbwJ9kx6Q1YVWJflO17h
gKDdjpMp2Tcm+VA/ouDCh+zGLoSvr4ClU72y1M/3ozw5LtZWcCtulmazOpFanzfk
oRLWBZQ6w9Yd5yX3yW75F8kPib4ut3vyGmHJZzh4N1CuBSr3mLcVGqBzsX6S4Hi8
jHd/sXMLh7Kqnr5vT+DDip0UkekvAF5cUU2sL4EbEGHvURx21Xbgwbx3Ygt4Jadp
jatZBOiYrCMY6S1bkmDqHMKvwMkELda+BTCFnR/QL+oA2vnoNz8oglyRWzwSKZU+
Ug6uJteh0vQjsVBSvK552H710Ir27r8q4CwpA1FRDpmWhb9LthA2sigUKBCmJoAk
GPuJUfK2QT/mgnepylsnDZ4z9WhHTLjKMySw4uBQEi69G6wFxwxaN8zeEyl9Le70
aYRjdY6cs9wWZ4eZpqhvXPZK4zreeXV5P8Lr1G65Pd0Di6h4S4NbjGCd2Kys505i
6sjxCsc/AQ+DMccdn/aZPBAON6VKz3QWY8IpmwlL5CgZ7HeLH06j7mVnAms1tC/u
AubOjJ8rAnodGtfigVOfVJzED0N4ARx4dfrNTlncir7EsEgQjs6giw7OTS+BfuG2
Cjo2Jd0hGBHgoo/gI9XRULuavIo5frKV7llhiOeZBp6J72D2rf43n7hP4ROY4nQv
bEeQKEJZb9U+f+QiY4E4UmFnPI33yBuVCury+QWlDCfkVNAzreJIIm0VNcAL2hF8
OcZWhtSBhXSmTnQN/HF6oLiKoJ8euLXnAS0xEQP0+536hvpg4xSVwbFcdxElLWvz
1mwLusCQRu30678TrYwoW+ycgA70XNpDOvqSXedu2AxUO+Fv+jdM8Zg9D1HRHALw
mNCg6xi/8mzf1ZYk/BUGAwjA9zTs0c3xacWXOn8YiNv+HTUnKoILkBf5qoGu1/yQ
BgCOVSmOu1/EJmRxnNDzziOTUXQeNAXlLKDzLSvp+M9IX/ejay/cxPc/BAShRxfw
jvjsZP1dkObVFDozzkN5c5p2nlRt6SksAmZywr/g6s69jfFvn4LqX18HrQpB1Vmc
YfApt0P5rAEx+g7MZdFjWtW/dnjsd58RvRaVKOeaYbnzcJiHgoqaHepz+ADQk6b4
RJc2yEN3Lgqd6MNhZerL66yfA+b6yK+0xuXXg37ad7zhtKhMjh5ud2HddYr19GVg
rIMwS1Q97FRffAqTIpJbgT137bFUmdKu01sKPh7mgAQDjgzwNIZRIEonkcgSg6GN
MuYMPHpMt+i8MsdBAbqwAKR/kxFhpubywgkP4reFPwsyY+aqkn1GOWK50cSSVkiU
oe4l4X28z+uKfYxIqLeWJJrq0CbXQdJJ4/fdcHG5gUIpQFj0hTz3gRy4ZLVMMSxe
+bp6tYHO5bBz3TLKGu1QBaXpr5l27Htd3cOs3YVaqn4aa3ApgUw+rhqpUrPQMEOY
MRYp5CA2hPB+kQsIsotKEaJYMTkOkqe1EubkUznXdz6T7Qvdd9DA0zicxLAIr1pD
/YTDtSCs+tJNVn4XTXou1F6PzFzT/8bH0nks7VluCOcOA8YZ41HKrnuSgVhCVjhc
4ySXEykILeAiwhhc229XnpSmvhpLn710aR3gL8CvRmPYlqt+xrSZzY8iU7amh/OS
B1oa6VyBu4LnHOQKYvu03oEj41k3Fv9u7Q2ZCjHKZn5+uo/ySRtLuuUT3kI6INPK
8MG9fCCmeN/kqX17ljIyN/IvLx4yk25kBD4XbveF7UydHbumDNXNOAq6TE+zsbaY
uVaYm1cpDwXoc+pYc6au63CxJkCB9QqNzTr7DY1MRmoLsybK2NloONtVS6sN28uO
UUCrV/V+FSf+h4l5Q1tai9ayBoUPTB82TaCA208BDNSEGQYB9QrQnvYuTtS9axwH
lPRnT+0dISrDaYEcy7rM52Tm3AKUFzvXGkJ2BGQsB38Q7wvW2qV+YRfIdmdogIRZ
dmZAZDtY+5K2/6sj0lmQCSL1t0pVNBlppDLBeHrqcr0oxLE5HZsZt6YER1OKId8S
EIAB1EWD4t9f4DnzV7O40jjgDUBlRz23OaGDwThXRHilcJb1Sbi2BMAvuoz60zmW
AZxJ+VVsOca8Z/In0hNgLrWaSicBzkum47yiqRZImgixii5/s/xIEOQWpISsj88l
pmygMLGq28NsApwzE5j81BwhtP+KR0YXg4+aat1sQuOmaL2XIT+K8soekts4Z0+8
MAK3JHszBVThmpaENT+dMfSNlbP/HDehYXfHp6CzjofWITGikQAMpd3LG+E9MSqH
AY3AlkkotfHttY0qkDuK1b2JkNEqdgvX2fNCT+0+8o/bQhfi+I6VduxuSxEs/JW1
quAvhhrj+iAuo+lPjJ2+sqoSiGgi/jEamQuHVLezwcOqpsj4u5n5useFEllQ9f2E
bYelfUCLe6vAA+/jOMVC3xjTds8VyxpXVEQLe5FX4arSairthafsA/HbuNx6L/X4
IqlZuQSe+cygjw3aVdyFx5a6G5lvcfBdazHjExAhjBk/JA/xcG06R6mUkrihPW6A
Im3ZK1HekzZ+pxrFxSFTALq7A+cpKOCgmCOkmSrs7geNs0VSSBflqEdmXnXgJN3S
3DdSMSpq4Tp/wfefzpObZvRs+HdZH75nIl3w0+l3Zg8UXbUt8SyXZK2DBj6fwu0n
jMX3kLaS7pnFxjLiY0bqzCYKzguFoH6tzkiETeMwDvLDNnvAMwB9FOFQF8nKCkS3
4lalziwHmQjH3Lct9yTTNju9ngidAHvDABbh6nCn7njsVR+xpTkh2TBgDmFHYI7K
iWXhP9cLG3HFOt2L6NbIrTZsXZLo6pinB2YaKTBo7u9HIJ8wtPnLHebzXwC38OyU
C05Pk6lDa895CJHPVv/0os0c+mJSCmu5wpZAZpAbqsPiRuZXGqYd94OUmucqtpEx
y5zHr7Xhr3/jpG42dZSSKEB6wrkDJOGrwg60wkpjBK1ve6uNSUlayhqusalyL8Pr
JtCX7vjyOGzKyrRmw9pyT1LPVGgySo3MR029qN28yhZvJAWcFmp9MjLex3+T7QJI
MS2WbuIlN/rrad/dsfwkjs4rlgipknGRndLO6AQ7SnA7EfdiPw7sAtzeAq5iBo0g
RC4BlTsGO1Ebg6smP6TcsrXyj0YI/g+27CBQYIRuLa0TNQ8PRWHWzz935ijc83Wj
MJxrYAXSEHv7SvG9uLnHond5mFfJ33dxezVwbtenAZCp5taejzjkbo5OSiR6z/rX
o7sslb1xNXKbq9Ki71B4jArnJthxf9ow3jMHhve8HG7zq9bID7JpCFyFzNW+hQUc
mSFTM7RGaZPzop2MTDUSyDx8OTdW7g4RbIiskV+kuDETKBMkyG/KZjh+az7022tX
Vl3TURgFHuv7gbtBMBMSeIx/cvTKyBdpotFHpU0W31MBmREpcuLh/ATpbYVQWS9D
EpHeeZLE2fr7MFn0Oh6Hf8tYSJhHS/Ut99cG/wNZFYWxyH8d19hTaJx6jKIRSSWL
Cs69K7OJVyObXsTuFQQriwpaOjkuLhX6Whpo5YYWdCKcUCPb7+SjgaYmQUJkRME3
7lNz8FmytrBn11ropeWHmAYLd6EuAyer/XkD1T4TLiSVLbu1CYKtIZnZ4opPR2pS
TryK27oBrZKCLVFDJ6/3lhRkP81FGZFxYuTcFYlsMj2D4zKwpmBBrFL2FMxDi7Nh
5/WRg8jKIhjjZ+HgIVcMBLcTXU0FLPYqY5XOE+/Igma2sE1PZtQ6QGK0W9GEuqys
NdjbYIkpJP+h+TwT7sFBxkKSMsPtSA7Yq3mx6jEuPbohVGP6oqb5pNs0/Kj9Zai3
HF2AG9QfxqI8orqWEGulFdg1Vh3zEic75mgzGVG70kQddvikpHI3YF14RkizobY0
9lkSDY8kbE1q3BeVVUrUgkqPXmm0cfKSHNstkLWAtwNqYZzmhC0fGxoh/LC3wXYF
hEvWhjtBqkYMTznmAcrCZHXlfUmqI2FLUNhe4aQcd5zaSeEfPXlw6BMM3f6Ncja7
Ypg2cQnZG4ktF6Kv0cX8/1U7OT69IVAGisKKt8fTUhg4M5O4ohfqz7xE5gVzAnOI
yqEaKWo+EXz44ueH2ywc4F3MSlLCMLqwCDgofRSkw6RI9eXrvBkogik4/9WODkI3
X3x9rY6aBAqIw+Gk669o9xqqKiuhrG1uOzJrAMBlgENUKzcDFA0/APN4zmiMJKzP
yG5eaIlBfSvihZ7UxkRjyFnIGxvPvDzJd11AHOK+PHzwWoIhV2ALRZ4bDwIlAYme
PimFOld59dVvv9oC914EZrGU0DHBrsjgQkCvGKzSNO4VFXHt4XCr9wcTrgC5EmwP
zia9FalLYy3aK+z6BxwFJDkV5tRqNReHFTzhJhOfOYXRZXMxoX6o1A4QQhqL7Gke
4MTJxqm4gH5+JSuUuvYKmTxVTQEStRew53x3C5nO0XcJVS7YVoVYYtoF1OQUVGno
ANqQewhlXJNDmunEheVoV3Wh7kW3zXxNQUDlx7DnkEHL9iM2i6bmazNO0dSeIHiF
CWKLqAc8u5WRif7UA4RoPPUXEd4Cw3FEn6Bwjk/3ERrf1H1sz1vYla6LUApG0mel
+D3QhsYLB6D2CAvGdys4fM99HD1eoe5mWyR/InXSELkYnddHkCjJ3tbFAStp+kDZ
fxMxRq0iKsVDRSeVm9EBw0N2l4894JRsoT4+8isqecLd9+D6EtZUffiHNA0Kkw5G
IMCt0j7/VV4+w8sQimfIxd5uQEe3jXGLAhxJKkvf0Q/x68o8PgCAwZPNd6drNBx1
zbbJhszqUYcQLFZZ/RvxuEgbYL/gxpdYC+931mLTYxRj3Q06EzzNZe+ZB5ltXiEG
vzBeTgg11mF9yqDCST/LtKsNfQUWU3fpSp7JWZdI9WtxJEMhj82if9+BSRcO8QSN
UFqWM+oE0MDphJiunaVDlIMU+N1rP/h99iFV9vFLfoVIJpzcd5j98EdywODiOIZY
hZJ1dv00oRLwFF65gX9PlBmocIMBv06AvXUPGBz/49XfNZkSoXZXS0qp8SlQTNnh
uDO1Dl70IcGELVLOcmpsiewMZe5cJTz+EpHxnE1UEA2d1vz/Z+ks4QEw7iXbBlr2
/Fpj6YJwq8uKOPArJio/vCkWOyRqUGD9hSPzLTsADKtLEm1OsFi0IBeGiLib3Qo5
YHHZMv7RePInJgATrovTtz+vsJvfBVnkCFZXKKTUDwEhhWHa3NSqHxJSCnkQF0E0
w8iZaZpJgmN4NmaQQt+BUkSssr6kpF4q69Ar82/pfTeYzpyIx81y5g4mdqBkfWu/
wgDNAZ+9daUsix1HjrIU/W8Wti8ZWVWNqikUezvlgjHKFgkuUDFWEQuxx88bzYKx
PrCfI2WG3xpStSoQ0ipp5v7TANj666f3PBb/zKhYSCGo6rM9wzr7RSWoDOqkmnNi
XDk5QgIOo1fO8AXNNgxYCNWHhf3R4wfEXhr1Rg93lAOaMlhdzXMTGksxg1VDvTNs
VvONz4QbkisXFX8dYyjyF8GzcGfYTohrR3JBYikOLGjFNdwuwmpaJ9CXLEG4L525
GfN1oYfE5O+FAa++0k4Mc4j1l26Z/8Fm1AfDQc3QhS3qkvwo7co1VURgL2szOi3a
Xiq8vgfqJ2i29XeK0z3+qBRbAc/oLHSczoUYY7WmvwmLX90ehlzcRKATkBcfOSXw
vJAc+WxW7vfzwtb0rGZTOv9NnpX9xDTl3QgCTeVOMKzgTJ/iYxO2u7SoJYdzjaLt
z1XeGAPjWx/arQ0WQ/KMhET17YYZPVsvZymZTbcFmxRbkBuz0detFL/1XBxerKSX
lVsiLjsUXt33B/0YszQ3SR+f/pHYx5lHIA3HWkw+uv94nDLG1XG2LYVFkm3y7eUO
7Se/QN0pAz8fOdo32YZFYCWHoXkaHOmp0vnmPp9MfRO/7UiROLI2oEpJJPPBThOk
F5utqKPTGvcqGA7Z2+YLzHOOhvuKNT4E2Ax0jq2K5Yqyr5I5W2VG5dwP71H2nll2
hiX1XlOMeX+bpByQq0XriZpVA2JmplBQj0e/hRVOx2tqamofAZT2jlxclSYd5JQ2
+hQBct4Mbc9tzguoeqP6nOdGpTN1FVkjoESg6GY3N85iQH4/MU0maHRKy6GXWJre
A3O8ne86Sphk7pgcjXDehcVgLKd+mjeHTKhEq3WrKrCnEGfHAPoq8CfWPmQNBXxh
86toTXJW9GG2GGixPCFx5MQZ5rvrpWV+acDMRJPEtTDIURHBo1I4gZtQngDz9Gu2
bfhkRb04+LGbTmxFs+iGwwbgZYKFod/5pF5GPQjrL9gUL81+4FSs4JhAqsxPur3Q
uZdJWaqL4B/6uyfu1tEwPs3PPSg+vjopzDF4YPgCrOhlKrj4OrtNvg0pFMhYPepk
ctmpOnXg2tBGUuHGqz1fxIFEiDKtqZwPlxV+xUpsg9zDtvExHcyid8ubtWkijCXC
9A4xtBFmPseQZCELh2DcWT1RyZ0drf4hP312EvoJV9FWQQPYeSCHwsezYfjMWj23
RH6qLmO+FW6n/5wBNUp5AxjwN4bp4rJFg0egwyCP1+ZrB1QJnUEjCYwMu/6xUGEF
pXykaJ7d0giSM2mzUyIFPDf3YrrC0Cfm/j8Ykl1VcHrvFkGg5sOYOcf2exVbBjeH
iNH+gwLYAYBo/RkKBJ11fCWA/V6buZzEsyBwG0gAJ/enSXpl0byrMbxuKE5iNPAp
kG7FsAOLNUNpq8/nw3bGrCnr1OaDKSOu1KtQjjtYzrxCiSoEdGO9l3Qwmwt7V0ps
On3foTov9jHLKIFVdfhg2uP1R9XHLILq5JERjF7GPClX0mg3bXRO7NjIqO6jwUlg
hA3aT3uB2gKLo/dtYuuDkm77+ZLhF8H7FBrnbO5/Epvh+uzk66jSmjuW+ZcHetvo
AuI2Q+RLEpBB7tnYxw+ecvDemYaYfeciNzOpoS8uo3j/QweLMY9+ZBQcg3Knwns8
rUGozfzZi+qMPyiRGhsu73zMDWOKBv1cP/zsrSbAGyHRwaSN8zSwCbuCC6N957vh
5HY9I9eD6DfYuJPf730NHFFOqO3QhxpSu1XkLCq0+fwqELwsXz4/ZnNK2D7ZunlX
bS7JGsXGiysS/AqbYYn1ZY3xBnymNelatZQ+civcDxwZWxR3NH99NYEIbTn1CW0K
D4sbBZ7Q3LTWt36lttHzHkjsRQxMRDHRO1f7uj7AGsSSjMSHDa4TTzijI6b73v2I
wYGJ8kGhK7jSSnQqIu08giSQdkgKNGqCCbtVW64py+xAuuVPcu1WL9HozVsB4EpS
q4Jg2T0NGNvQlmz8IGBVXhTSEdBNB1LZZZD1L8j+kIdQ1I3rFdcRnGmkwMt29Fsy
YATZeaBnHL/vrf2SvitU31aSG1rZo0b07fPYwEudWu82Zr6+HNz9qu6U3/51Vd/J
7vG+IgfTRSAZ0gy/1vBFnMHq6Dm1xm5I7Qj2Y2aAdpIKllFktzDztg8oLHfF1j/x
X5cgfKG7LIMi2HfOm5I91/8GKdl1dvjfCwjTlDVEcL8tuA/OZUKSnqrhlwDbqw6a
U8N0Wl68fjYn5kAHC09cJMzjTsDW8dM9b5I+f6CUnmHyhyDRqBbv/nUNgNKp1y99
hPuDJrggC9UikEelu5/chftQU/+j4wl8xtncWHwzzyiLz5g//MdYsIN59pTAu2ol
WyFpTgwwFCFOnGe3ZMRa+oKGaazMdovMJ7DgEizcVW2QK8ROCWDC6QoBV/RjnID1
tvJMfQJHzQnEvlfV/1tTY6hTl3aFfxJbOJBJiq1GFjqWp9cW5GZy+JEmb9YzXOmm
zDzQTwzsot68kDChfxbFfFwAeIcTfV3REvXmPIScrrjJCum9d/AIPUV/5vUTO+4L
HxYCjnrrJt8diD7KU5/DfzFvJ/nAcX1ZGkkPt1K9+zebMyYLfQrg3UPdzBVtfO0P
XlgpbOdc6x1YyRrfTOeHGRan46L5rfZv/DQqXNHYlhC/dRboZUyxazt8C2Ib58M8
HUvEMe7gfyXugqWkPeesY2rZGZY6hJ7BPB+vFuozEM0WxLZB9siLAz/foVZLq81G
1i9qi1WZXcZIPGVpIDmGdBIpTkAwpUD3vZpfpSgHotZ2pHAudfmqD7k+fLH7q/XC
qG9KS1D+d9FSW0TBjRKCLz1xZ+H49ZqnLWJp14kMj4or6HNUvbvvB3dZGsdiCx9M
f724cdjZgOxcLKzTPxhVPYdB8TmuzqoyaKXzEOxXpOpOQz+R6t8IG30hsp9vUycs
/V4ImelarKixe9yk1up+Gnv4vlT/8gkWInra1P+tMHV260Y9munkgM2JIzRNGr6Z
SFOxovVYc3d22xmEeMGobbiRHFT6WYLqNvKGNmMJScS8NfQ0vGoL1rntFv1xDg8z
iNMidoBFS1buN9foRGqTHIhALRju1xp/4MdGEpGfQZbIfRK88gozHiL8ahLbvYgk
+Tr9ZQjG0ApsYBuWwtEjywmkMo8qjY4HCfEHv7VqDfEWzCpTmv8LTG90Yh3+l3M8
mWgFu6ItFa38RMwG5pzVE6DOelUHePMmPMuR3xe8cH+MqypTaOGO1bguh2JMjiYD
qNBzgJ2srxe9JY82vI3HzCFIxLb2FkFpF+GjCvD3rLdwcRncPxRdj+CXLv6Qvbv8
b2kEToIpGHdmH07Vx04Acf2q9yE4VKG0cYWGP0ToKCcxgNrqobeRg7OhRQyUnp/O
6NhCDBHJSYP16De2jfnCk7bMC2C+zEVDcagL+dzdgQXtWaCaISqhM5hd4XMdcJA9
eWnkwgSM6o8rtScDIx5is8NaaIu3wE4ELj0a0LRuZi0AY7jyCHR4UkL2sHjQRO2T
i95dAIaoj0HDD9UqvW+QPfOPks9tfFTftqfd9g0JX7GM65c3PxbzTHURcP3jqy6D
sIfSm45XFS30JRyG+XZ8WuDBdWxxbaE3qG2oBIvlvpX2a05ar89m1wS7lCb4jp0E
FUKFHJta8ZyXkhU2LA+0GXGtF9VzSMvPfxZAKYLzIfmqT3LskgCHoM2YUgMWo8Yp
OUPOnFJyet6aZn1O0aXCqZIh+DA2hDUuiSxD1owjZfQEntBNUofqxR0R292P0eyf
PWTsGXMf8qSkEjOcL+YfTqyYaBJf8iE1d6X1dbAFg1FzMaAS7AM1mKepIX23hBNI
3h2F6jR0Oa7A2BHJ+0qun63biMbT50UcmETIZMGOE3OvvtqItRDsFxC9wHcf+2Ot
rotOqrqN46ORHeGYha8ahPlJmhfc9kZNBtAyJqTfP5pms4W1orf7NEq42XrkgoKw
ohr4gmxGfqFf19lIgRkLQpNKGmLaZLt7JAhIK233McFobv20dExqYF3XpcO3HoV/
yTfejNbSbWVjNJ2BKT/ZarSmP/uEZoIw/v0yVRDgLAQHbbR1Jxyn/myfIPU0w4I3
Y65/eh1Wq7Qh2I8L4+cwB46902/nCEwFas95FQemVPPKEGRVtaZWRII62auaUp2I
wLFPm0IDVXOwHIPSSLCEjBvhvkRwnYPvjp5vOzRiH9e1aCVbUUeZeyA5H3pWz4MN
yT9OFy88yU09o6EkkI46xbJDQ3tJ/nwjYSFYzCi9thCER2GoHMs5Yc+SjOuZ87xB
uo1OY4OkVZfcvo9E1DNM7Pw9q/Mg39WjfKp7bi3nNxStul++OKiyewXRQbeZJa+U
ajKFsS+gGx8YLnTRKKcX6lLDlT8Rg4vgnyjrpi8sCO8Min8XE4fNKhdaXLDUJYhV
OCyYXq7fwsYrzs11hVSHAU8YX0kflDFYIUEfFQQXH00Zo2tx7wL8nPmS5xJwy6e3
10DGpdK5u2Fc8C6h+d+e2vXH3skPLDNgEbFis4SmD1MPD2y5i4Us8O2aZgfXi62g
ggOn8Ay163U3N1qJAtzxcXTj3Qq9ixU0ubBAVItFv6v6RF6yrGRHiJySvOXC/7ug
uNt7Kqte+cPmJiY5vFSFTeUN1bUhLl9iIdqD3QwNxqDnDtzZdShQqcr/SC8q7Ihf
GKKGVPut53592ToJTUT+9yRzDCyRw1tz5yUFXy84d21lmsEbe/s0debXbw5gwjlT
MtL1tMIvsyfSL1qPlJj4oPIMy4ET71u6qRP1E283VlnNAvb54Ca+ooAiLOadLeA5
27lSh3LIwdnhScSYk60rvJMCimCQrFYPzs2OF5r2y3KXestYq12Aft1otaU26tS1
+EW3/gqqXusTRHH71YGqpFBnMO7ru24tpprDdlrNhBX5c6uwC50RqdfTMohzzWsV
RDEP80OPor/znteqpHoHAEZR/GzbaRN7eL/3oqx+9pQQazATdpxbUFYquyYVTonE
8vEktYWyN1m5kobrLUM+PPx6OxzGAy6/J5HvSpgegS1PHcDEmvHn0mvuO3GZpU2m
beTgyWMj6pyLo5bMXB8+hlTVetaV8kM0eZB1a+4KvT1U5l6AfIck+diKoRO6rP2J
t995a6b8/DnQzItuen7RqpxfrSZaOLf2tTNsqdSqtFyD9X+v2xlREv+vAjXj2IA4
PFJgx+PyS9imFU/MFifucK/7ErInJVL0RO0gdXBx7S48PLGX0QKs+aawrk6rqfWw
o1jUKskT1mtlKLmf6OkIQNaqCNhspB8II5k6VHqJaPZVUIWCO1p9vu/whD3ZV9q6
Yk5M6H9xbX/iS1x2aWZPRvwLUkxZnSfsoACLz62LFCNVwgiAjl/4z4gKtgaUD0u8
uz9KuYecgEn0KHXEy7fm3tOLVNyB6BkzAD9VsGws3gz1h3+w9fbPtlZNQXry94SF
RFOUlRE5IW5Zp39nAN9XSfF4emYJdm0eHBApKy7se7iBJReWqrhMDTCVgzo965Sa
CGcHFTbuyfXS1eUzCxpAXYsL6g8+pVHrwwgBvqZMVrDhCBMcfFdUWLwJv0kgFPWt
sKdaGhGL6FPf+y5mNk9NQiIITgYTB0/NVcMPyVI4+/3OGL92J/xnP4VeAmNILjR/
MoxxggD7/QI2UgGc/oQxAIibctDfelT7Os8l6cypIaVKalD/3QKFpbZTroqGG4yT
Z65IkHKfheofXc39/dRRaGANNeWrGF7K1Kk87fNGgJinY/HC6wFRcP7ZnzG+n3yh
wyHXyk5Rd5J8db0K1mVa9c7uOLjaMauZ/PNnHnPhblku9RSpEDCABcp2xPXbOR0S
xHzB6JLIbFVVYHKMz/uYePSiSIG4A8Mii02S6B5ocb1A+Gaaa9/HLutdG/KOi2q2
b7BhCtMRpL2jReRkcI4gJGL1O3iRnPaMnf74x8EtR5rQQNfC7aaCWxD3BNgRmUq5
qsqEXYf0eyQoEGXkyl0LCvvpyVRYN0FyXUOfa5cb4PwEaINI/d45HDAkcuA4dWYE
4+w/ogvoynnbKnZ658thvOQbWhjOTAnzBANgdxVo8PrvaDiVP+lx7u13Lz3Ek96F
wFwURnUV1dfaSr8OhwjYB4PH0IBhPWCod3W7wkQhYpmL0oMfB0ZoS+3x8dR7XwML
WkyrA3YGW4nJutzwvL6/4qmUDzbTmdUEhbqvr2rROad2J+gkF+lLru2PSf0FrzSD
SMc/sRE0yP9ItSw2LKY2o3HSgryLMzla6NA5zmBLIL2ToX3mNM1Q7uAfACyxki/2
kEv5sOHb4l6SqhaD101v4+ch0DQoeyq8l2IjZ3ElSp6A5T9/Dg+t4idT3o8R8d0N
M9wi/cIAlq+D6LoGUAlog2Uu5k8/3mzaskcaZfQ6SznyxItRKIHKeMiXf+Kg19q2
iN9VjGze7JpcmYl6DL2frNuZvljnTH4LdF07zxEumeQQPF7r48H5VzH1s06ARGqG
a2t9um683PU+wGPVJHlIPck/F2+XFbHXwWj227q9N559XI0sM+gSjnc6uyqBdfoE
w1pguBktzTERuy8kBdCXI1JkjQG9yDtNOfjp5Yb2jYcMgn+Nm/DGF/K33xJ6cupG
G4iQyXU6KaxAf1Yw/c7AIwURaC4aEnRtWX18CmXfyW9pHkf1wqbWUpR7BEhr0tJu
2K3pntjP7WVQVuiSYuWSFpNWX1NWmrQR9WHkm/o5xjHkaWUL9doaRfXmRp9S038T
RbVKwGBvP5DSmRq8AqvV/uuqbHZWAshLNvO9EBOWaRNw8M4bO1FXbbXtM4k3eFAi
ZXsvQ+UGmBE+sT+d8jXSYYJ1NUe0XmJtI1+GmByCHdwz78HD3Mlhx5AALs9XCSQj
tOhKo+5nk07apjvr7KjDR97yj7dbDw+OW4TcGrd0j/AVo4qjNb/jBUDIXVIaMXqL
C89OD8woiszWgcnGEOgIUZGb9lkkN73nZ2PQ37HW4YOuvaRVFJ3PFfeiIBK2k3XE
nAmxrv+0nObWJCK7ITjtm2iQJ/obSKiSQGXpQ4/7sKihBrUtBW+N6842GMsHQiPi
hp5lhE3dIIFAMrZVfA0wDIdBGIFkjgJIRbt5AOUL+0w/M6ZSLrl+YAH2HYrq5fyo
KqUSIlGkNhfYwWZv4n3HzkNK2uFj3bS87rMbcWBrLouzx2sLZSMqWZPjU3l2YD9R
zWLOHyhNR2eTE/hJ1D2wWjPkSOTSsX6nomjDrHywEFFm25Zgcm9SnSXmQoDDQ5Q/
qPbEfaSmDxM0H7TQ+zAix+QC3j2AAwWfxK+Tk1EyWYCdOCgP4t7JA0LAeWVu9HPD
Ul50lnP49RZtfMVmyfb9pR2KPfeO5aKK0P0VCFNUWkBQrwVQD+Qea9cpGSfSrPUD
3IdushJgQQQ0oQw0olR6PMa/HWLa6ed+uceIHwSY5iThBMX3KSwzt+p0LzYi54ye
S4/Rl1jZ0QpLPinStouY8hA9BO61fj98B8AigE/ahfmhX7Z6gf/66l41ppRj5yWi
CtryvbPEkICah8RAxSU7PtcsEL7Y3DtsVs/5+/uYqBPdhEDSGVsfqxflqEdXNqnw
BC6s4sqFYrAIhuFCHse2Dk5KoJ550FdV9D9jvemaG6ELTzh1vkkdIfCk3IYKgF+W
7JMu1XUGlmJunuRzWq5I7qwek3OypQng1/NWMuwoh3s2jtdeHMyo8Lb7OFGTpXex
judKU5tCdl8OS1+aVIS+LbZbz2J+ou+ZcVgTOtgT2Yto8Mp8U43KpwW9ONCLlMQX
WvR3jXSl7SXgqbJtOuHKf4aLVsXKjjBKgEvrPO9HABTH6CDTk99MFAdjw6K5bBWm
c8tNtRRJGQEysBg2gunbGtidvM7fMyituSvC/ZaJuhcemOtzcgNZ528ebSgrgh1m
jbGkwXmauL+lQkALIsn39AbuQeO2nK9ggh1RuwDbsOMmWhPzjyRDGf61mHA+mM3o
TX5ReAPWOq8jzKmecVBm+KOvpEEl4bbakNqsCWncVTMUoO4atjTByQcDVCXpzCBc
bLm5ZqlidrsxwB/lQc9QIad3ixUIYQye7CHxV0G2+FD29lhus50LcLK9M3GuU7gh
7p9GgZHzApCy38+Y5tDPdZsj0tY/Ke8YRGNK6TBA/8g5Pb0a6u60ufU8HUlXTo8n
nrNLpR2BYR6fjoJzDdRnEOPTmjigDt9U937ggin4sqHtHsjcHc7vMpintfx2Q+V7
m9f9CDNmXhYTedzdTub6RBlraC1Ju467LVNXH2Fz9HVcmN3/tUthNV/1adawAO2i
m26baFNNuHYJ/8B7QxTLx5EefzzV6dclT1Bz7xCcBiXCck4rZ/+95VO9/l/wNFFw
ZESh7qcQGbr1b4QsDh9F/EPVUARAYwY+LI8fG/GiiFSP7rKwdhZ9sF4u699//UVI
arj75pQkfyUGg3C59LxvT/MoQH8Wd5OlHBjAZ9wJH9c/38je+092oiBHZMNjVNsD
9iVOxU6kUZtT1NJj4qIMm+chM6QL8SK2Xz89jnhf3COy0nXY4dO7lGhvFA0SmGko
UD48mGUKe1/1hiQiP4iVd1uRNLPlMCN0AroYPas8G7f6CXSKjhb9uJSRIG3U+IUy
JP+yil/bPw21CkH9P7ftjcHhLKyGNL5CR0jcgxxcFxrptMme4pWIBalpz2dgeFfX
B45NRFYbyIN+S3abDUwLN205rbyt87OjfYcF7XUBQxyS21EpMM+OKodCTDyPndcC
hmhLpPhVPMae0cOF9M6TSBwMtiQpPGZ+Ldmo0aVgaM79H9Ub9yCgP9BuWDa0mwsN
aJPIpExvXo9NsMtdVEgD801xnTDfn99Qq8I8H2xdVuJYQRQqt6M1EwYnPThPzSK9
zDV9gFwmhevyaDpxfytixfIH+baS9DihwcbVsa8JY4PBW2dFWcKAIydReOxHs8YT
IWa+/99eZA4KDtlnEgwG6Dyf0Ryr5xT+7/xv8lx/BqjQM4EeOs7iV4eR8eSBFv7l
mBUWZfULJqqz8Eq+RcYbEfGa3XNyaQwlxUSSv87cOn9Ly/kGe1vtnEOMGdNYH+P7
Ypd+cw+CtjpO8FwUJ8DBmFGdNRKhzQYDUY3+vrgF7v8l52dsDXscYUuke7Rnxuok
oPPp7wnAC/qKv2KIO1NVMt+dUEWnaSzag2/aar0Nf+cq8oMZTuqHPGgwbkAnLhny
MG7eobEK2SkBsnyx2bDU9IW4VyuGTXTx/5IeNSdta10bHQv5QKD/tsQ3nUK6bMwD
yTiLRG55mBl84tcmqOEFS2q7zxOfpF5cD6EBUm9IK9HM18OuGdS4BJOq3dutRmhp
9/VGP/HI3+sV2niOzz5cdJNhFxMchbfHKBbxRU1rgqpGFQSweR/25EOZ9Vqu3ddQ
uiCduHAvsAu/xowrge3ItvlgXmyCo9PvtallP7koSur9MieOBqPHrwj1V0aWxEuL
FBVQet/zXMeK3H7Ck/QGEymrpJxNjuDvr4Bp+s3H2wXmxLtrxSGtcPI4J0a9OJHq
PWVytTXMrdrD/O4e3tm0ytrjuPZyAH80AnJ1QDlMcFxU580VTYUojdCif+kVJO1Z
UBcgNKWjUqKMtlrfmnTCmEvezrtDlw7FoaPATcNVn5y3/3UE8EYssKc4I6k1R0E9
tZE3BE1TYbM/96HDj/hZ7QG9qQLi1H3E3hUiS8ycgmp/RLp/Ult+Xjo1zw2KG70E
NFrRUnI5C4hiQOwESwWo7wnv9bX/0EkGxiqJWkOraWJACoV+hcy4454gg7boUU2A
beq/zN1UfjJztsS7BI9JxD5EWvm9z5w5RyBWxv1Liv6FVyNioLUHuxdVcWzmsZjr
flHeqGDezG7e5APjd2rtMZwFdSj38mzEdFPxJcUDiix4tKAqVbsWW+xnS7dH1LXF
xoEL42r1mkmiIDqnz1NsEZ9Cjk230XxsKRuxs25YAdQBfb2XMR7E1SYThL43rolW
9c8WPrZ+S1amqTixNiSYzljT+ycWjnspLF7Y+oAMieTIkGsVAKcvNeDaSAFYF0Wb
qwp4oXZ64LZ/LtL/Kuc177etG+/2ymkvhSF3L59PSGKKelNOrXZAEZK5LyDOCheh
5bsC1tD+Zqlk3sjcxGBF+RcdbzfWfASRLAIv75KCb3HNQtsMGizgpN5ZXXIkhx3Y
F84zaO2t+laBNf5VIJfc6VfM4qEDabCgaDUOcOCSYkUbUscw9MsZIyCGM57qK8Of
orSpLdy6LfAjXyFc5NTDqAORzoSDmcUkt/OeOvnxWMypp4wyuW5WI5/lnZyOFFze
06WPVzOLyIA87j4Yr63Oyyw9CimtZ+k07D8QKgcIvzvNhsa2qbNwdhL0uES3HZgz
zJmXE/VciyiPr3Be6Bm77cRjFhr6ibntipOntAK30HkRUVSeq6a+qk13BlLshEaL
YjTAJ/k0S847/tvhgksEobKuuxd+37fDr/meNJIpLmT2Uk7/PsyWkVAqi4MOd9eM
KuDX4VtD9f+M8109D1kYa8qd3cC3mpV5mJLdaoe6gC4wpHwcOyFAAwSWAGtJmALZ
BSLbvtddceK7kX5yig36vF+jH+skRR9S4BdgK537BwKgo7dHbh49MbDGAE4CRnBx
YL7U4YhcIE3UbtSCMlJNSmE74RJMVUClKz8wpK/Gi4VVw5hMjqOWpwZ0QhTGl/OC
pDl/5A87dSA0vM1K91wlfgYMFOLFgRSIcG2UnBTuIgva/L/N6BUiU5ZOeg9gzHkq
8bA6HE6LFBsKLiGMBAzDjKYr1ux+A2YgpBC5GJp8ZiZkrHzL++8DhxMVpbrKfsDy
IGX+FA5pYcbmx616XtNTPcPk/RRD2nOpG4/joD8zSxlBYgbcNLG2nExc5Mz01eOc
+nWhia41kdDqZD9ZZs9eKByzEvqUakq6lRM5Bs25an97k5LnbdnesSMqrDp/R+4e
7WDQHbussaKzqlltghgmlSIEqenCgS1MV6JnxXFm0oXevyexIlOGxMUcGHqMSThF
Lis4JDnDfGwmkXAJUEnvnGoKBvmzgaBLJMbh1ep4ojd3naxtQx2RI9hswDFsEcco
ajlX1UCnaTbMkSzuJ1ptYKlKzUvHdMWNay/f4uCLTaYCnDgfmCJOlWuB0gf3p52P
LRa09aT/XmkPSbbZGODNAHy33InzPVyPw4i9/E5R2LfB0OOWRF/LCay54j7A+1Xx
TT/CBitWpMGSveY7FXiHkPJaXRilBpJejm4rtcRPFs2NpGFaR1Ja+15EvBRwHu7A
B6NZKwCD3L24Hi74A1OWMnicUSIIXqGHCgm4kAtfDEWygGU3L8xd2TOdYvDKfL8O
LTQy2H/h1gMf1yewyQ2ig5At+DfeRUxznbY39I2W/Q+/r/f9cBRlhz4vGsRaNv+E
wUqZqB1VSfGMy0TqP9/I5bYiGybqGrMGPPv4vPMlz+fW6qjWYroQA8O7iMMjvvve
U9oWNEuZMG96N+InicaiKCiBnNAVHteegeKE8S+Fz+YZpsnQYrzeWi2bV+U3MaJR
8zEUrXdCuB3+f8NXMjs48HTJfzHXRaoOMaSgDxYPaCIbCwJIOv4rz2EiR/0TEFsJ
J194V6JNCclO0qk3RhQsYQ8WNJ6JdON/jJalqKtgHFGpWvIDax7VrWX8FDQ3dRLU
1PMoogL9Ej5IcMAmM9pkY0jTGeTl9g3r1H5KliEzb16/qgzga7kQCtvTmgLdlDfb
3+0mBvY5JLygyYWd6k618dw6WwDJ9bE4zjhFCDJQ+OOR7xweiwyuTib0m2wj6NkL
w53Hqr/tr/qvTCbmds8ZKYwv6QF91N+kXvDJUHpdpeOzsM531P+zv68M/rtJDV+d
uuL9q6IFtYyBSa8X0heZnOCihBYyoegkIYyOzDQhAuWFj2yK5N6I+co2YVqr3YVA
ULdCf0D6NYNOe5BiCfv1szvlmNxlG/tAbOGCFm9ViP0nc2LusavY1erlDETGK/AJ
e8ezxx8Q2jfRVWq127UFYkzLIpGWB3eP/59lMgZWQy6tOVT1SjyXOE9kBEutQQUx
BY+LL21nkQXrhd/4192JnNwBCj6BPJqSNWT+J1bZdN91oPjisl5oXcHv4J1TsHtO
LSoa8nV4hBFPt4sbYGrUmdbVnb0JESY43qMmDL7X0bWma+vCuhSvmDg2zVpgRD62
3JcYz7SuugUVerrxrke2uHiyTK980iT1Lu1qL/nUBBdtZ7nRNPTDxLt4ga2c7V/g
EsNWI9gEwj6fR0VFHRaqyaubu9TFRVu9Hq0vkozUHp0OUIf16NcqyhX22ewaD6qO
PSKJI9d4yH4v1gcvOwz5p4oKcUAt7PfkPG3utlWR/afpqyvms/FHXRmtqgotzWfo
ipWowpak1NIqr7a9kiVmOmCgE1o3vFPJzPPjqyFCEe32PQBNkssW/MwtRgTGiPPs
2CZrQkh26zTLA1wnf1CW41lgarVHllVsgEVNlFCCdxrIHx/sYdFJfwj9l1E12ASl
EcDK9n+beFQIIIsln4Myf2uYZmcuD1flJ0Ovn3uUfTk+m2Rb6OJQnEA74s3uX28W
vuig871+7RfTpHuujzhrnSyrY8uIAjAwYrUNujH71Uye05ku5tS+iXtP0LEl2dTO
YplLfs6s5H85qyfid6AEqD1PmyzgV/qxX8riyqesyCDPtu4ftCqVcTCeiJt9hVXh
b7scfFXwQmCKBir2Vbdo+0fVn9g1o58SvC4AiMbdBlSCBObRom98ZxjSPgV6vMZ7
nRwu0STQ3FBXaWAVHtVZC9pMpELgyzrjeFgPlAV9IKPKTtjoVGfGtDZ+oAS6Ji1w
aBUvlNBKTSgeUBCYDEurapziddwl0nn+8uiasjqF2PhX8DZMbStjb6ekIDnals+X
emKy2KXknojNtvCOyuL7QSuui3DTcyo2FR0vueQFf9Gn6dDKFgImxKoAK+Nxgezs
BQ/qjXjR3FOSUQ77ygZGhTHdUxre0AhNfUTN4j3sNERxtmLJBGlJtM2MMFhN1mpZ
hn28dtmTnC9Fovs/hlJByWs/QqKKh5fVp046gT/Ff5LeENiuljQx0iLD8TxwXh37
B41bwpZquYwic4ACi2yS1KKA4gVUzzj+/OQ8IL1NiOK8HKA4gJ0+LacCy9Qczfa/
VQny5d4/rVb1jXUKBEk8lkyHlKsKhkw1EtXYdmELJVDqwMgwFCUVrM3sakXCq/cZ
jr9ZS8i8Wuz+dvyaDjxSGKRXFxcgh2pnv5lmx4BBLKh/SWV1Tm/M8Uqajs7h6tC3
g5UNSuhXpeTncNfSQQiJAUAp5Lxlvlpd2kfg7fNNoFnlKJsitbyj9lh/ajgqj/4g
4KA5V5vHwkzF85NRLH1cF/bneuTUsJ4yoiRGZSfw978nkPc0siS69NIEBRlgkKgi
erub+Urz+OGYa0wXeaoxEntE38t5BQ7VCBIK6a7Qmecan+MH5P5Jxm2bpV/9fxYB
XqMPgnKjYeRn8WCUiBwd93XSP5GdLfuUEzOyEUplM25JeEmcSvHdgOWHRvOKBtpm
hZHYIZBferfqyFioR7OHlWqiKCtIlFFegH4TdbxqU0wRv0EeNjFraaAtvd+1w3Bx
eByI9QGXYD+pa4mM40ajT3MOWSsZT7rqE2bfpKzI+Zr5H4rTw4diMY/GZukg+nGp
18jAFKQIZVc2010XGvrY0T0uoyowoZ7T8EYCsCzH0DaG32+cs2xz3fnM90i+vOCg
/3APcvLsgC98PctsNQ3XLQohTzaRdvCM1wNls9WgCS7nsxoG5a/ZQAsKs4vLMn+p
KwfsKepsM8vNk9f1qu5WV4segw6tzTcOMqiLEtVyAqG6mWJpU3+tnZ2aTpuoPdPp
fV8k1+kchbvVU8QEwQgrM86wfitRiGdGviQe4dNnqbbNhi7HK5NjEW9CbUhvlQ2+
NzmaKiHXj9c3LQko0M2T5lwqL9EM9mihNVjWb+r7XCy9ap1+qegmqWgy0muXoPZH
9b7qcsbk2wuYC6dUSLj4oQshmqhPw91EUSKhXLNHem5zc+oaKPxjzzw7DGScTLjl
3uJ52wGPG/ROjqjBmuow5Nd24unxET/v7YTyC9y4fSdaXxvSN1/c02acTvDmsvWx
Or4G7YOxC8Py5mOd/LHoMQcmrM1lyQYJIqT/teakQDVRpy+rv+qKaLb+FIePAXTy
HPhbR6ml/JfUiqAx8UaOVuqwjoemTr5XAtbWWa/WC+Q5Z3wVGiPwWo6siu5ZBF9P
/092ekjOJHhNNBrbc85UaQJrvr8jBcn8eO3aMLt/g/0F4Kg1u+yFt0iOk10reeMx
0c+fNtk+58ZrSTc6+nhsX7cmmkRUoXbCxDiZpFkbd3KmsTUKz06cy8yRXTr97IG3
69ZsoW17G9edx7WR412x+dqj03QIdVbAgCuVN5asZN4HNXFDlzwjd82tFZkev1WJ
DHHoyyeJJegRvgAEUb4QXuuSUImKf7AhRLU7YpMW0SEFLdo9Aw42inxurQmzR3x9
Zsp5rMUcsSBao8n3cDoCjafhlGt4VBRpDklbwHM7ajcZFIaLw+zKNcIVRcLfuLFS
3Vp6p0q1dSROSIo3k7i2NhMRFXcCsVjUD83k0lFC+znKGWLVvsWCWONQbsT2iG+A
LaazpaHzmE6AXx9uNqqNGlR6q8Ki2CAHsjY0nMIFfOmsKfqKQgkFCbo/LjQhVAyM
PceM5b7ljZX0H5mvUfrIhl3K4da1TbX7ZluA0TyfUylFMHFy1dOZ4zKyU4jCmc/b
lhDl7HcPRcirtMMlCnnB70Qw9uYb+t1sY6ZffDOSzWbdiFOK1C9VoY89KsOUMrDS
fFw09CgkMtxyrLcldt4MqKo5qpg0nmkLpi4M7bNsUSLkLIQuzHAbYKdif097U8Nq
s6FDHFxyzszlvWfWNxOTQGpL5RloywQpQqyiKUgAsc+/e7Gd+8BVfTp2mbwIcpC0
CYT7GVHh+eV8+qyekGy/fq8mk8bVEMV1ZJXph44pmR71ZkWskVDEGjfUlHTq/fsm
MzPnE7kBQ0Eih4kT7PQKf/aAPFYy98HdvqwnXl5ADn/e5TAp512ETO1S4F+UISVL
Rwd5phYcwDy9Ry6lPge0nrbd6tqEBjjEiGwBr3e9ZkhGXNCZbh9uoUP9yGM/fybQ
6YVLWgFM6JqjCxTvZd7mI7XP8xMcY2yPQ2lWRtlbvW+AjaLge5X4Ux/F7WMYmUup
ZQ9sdsqxVwvRkFMba0XbSGKUV3GWTnX1dg4I/09YZd7qWd3wP6ykZE7FQfq23kGg
iFJmPiMLSX3l1kLlHCRCiq6dKkI+uDkla+M/DSKgprNbVaicCMhpWnZIBSqGyRHr
ykBTDFeper/fL2thUoL4Xe9LBfkah25GS65WaWEIhaLBUdzgnMekR32Om6knvEiE
U3eGEFUYXdivLahG+89sW7QNNB6QambC4QNWWtGfKEdDdkQYtxk3riyPpD+7KSxi
n7LFINwdDIFwwg0dzyPRuanva845nQdCvSkGx6AbxAq90QW5IcUb2jzJge2j/N0v
l1Dcyv/QI0fbwg0577PLtL2JOb7rOr3nRw5e5EhBMY6Yhtwhm2zixTeRkfXzb/Ow
LSmSSnaJtSPs6Fhi3NS2u5i0tKewFwZ4gw2GDn04mBeedTOWSZSiAkHdaoebaB64
kjRKuw/fDVaOlCL1x4UVtBWlCUYf82ir0yc77E9c9MVfcAU/IfUoxR3yffrClbE0
laX+VabM/8V64vVGeXg6RVm5+QhLVIM/TTZ4yZwjP3H8I+mOx1hsjEXTChYhCa+x
NLoLlFvs6THWyd2RU8UKNTqq19Whq8ppIUbQ15fPPNS6QCs/M1fmEeSzyi0KdjhN
1+7w2SzPCqcydWW1nYm9m+wTt+EjxnJfWKXtUNRMlvAYI3+n8IygoimWnkvRole3
aebuNQQuwP9m75CzBLjsx5X6xCiT2VIfMp3eIN2/6DAQ8dpq+KyBRIPtjeEcIM7m
GoZ3V+N/KjSp+upb8ybTDeDk9kJMsaW0hsRvpXDFhIy4GJTi/jOngy5+gD+iqm1o
yr1k+W2PbsHn5iUnS9ixZw0v3UcnAl3g/sBscOUkoiP0PnTHJ0LEqN0w1DRLGQoI
PsVGxX5eOLuVZXexiFUt3OqI3Iv7KJutKUfpFerzHdMkpc7tEY6twXpFbdPCq2Jz
IJUD8n+ogPCYGOpN1b09qNJt3ABfPpzCJgxOV6LdnkrUuhunOCTIRAPeI/AUiO58
BY8WJdq/OOwBNzX/NBv4ncN6quWHjBJ1xRSw3sxS0+5/r8cH66lYMg1VcA17113v
IzWWX9clY34G6s9072olcUoDcbG7ZiEiD/Bt0+LxmowiFLs8p0HIma8P8aaKyUYO
t6EYYZSvwHjfOxosqYp+ADsosjhSIrCdfhg5jl8ENVJ+nNHwZxKLlrMQQnW98dp9
897JfEu41czuhwPcgJKV+n42tEzMbFp+rbpppVRcDwdo00Gb8qj+F6OdrPDdp2yA
1QCJMaxe0sWXMePJcoIUBvf1Nz06tyrtsZYbZs5LPWFiIxwuuWJStuLBQcxeIfzJ
Ni7MW3KYdekLmCb3CJS840hu2vIEZ/PCUd39Y6iEqN4LcGBxEyQ1aHsCKX5aHIgp
KHOgKkD2GpwwivifP+3zh7VrYg9j7ySAzMkVxiqQnpgi1wvP+fCUp/d7t7H0EunX
H9FbmwdlKJHMy3U9RFUFkY+/6Lvba6pI45PnBG1wQby1PDmRRzbXVyMXmyJqbezx
2SfOmBjF1AILjCQ3lBjJXZ6iggmNCnc5MUHYSSgjSUt+llQdjyrMLGHvAZtK1soR
HqUcHIRs6p7a/JTnPRQ4GKkNAhTMm0CK426ZmGL7/58zHTIynuPKKWNa1zzFpcka
29in2um8fZDJ/81S+nJrsvXZUet6S2N5uPy+9hdfhbM/8Y/r//YVKZmWYr8uU0B+
JRUhos9K4I4gXvVx6U+ByZ8nUfk9FGore9GR6jHuDskAHji2Ig/Dl8FesjB+JOh7
g8evQfWLGbhAj8OGnJ1j+9mXTDqcRoQCkbRbpArgxY5geGrlM91luU/vBXDgz6zV
NJ/4b/RmHM7HRyz04a1nthII1CG5HB8AEr3F+2rxpQN7SX/n9G2R2P3eeB4I5LW3
iMU189uCIY4AX71XcrfvGDiLU1hgNgD7VPCpaph+6cGjrVRvLi48J3id9DV6HcE8
hjUv8ahCkZzC9rywRCNE341EWsOvZstTo7eD2Q5Bhl1bELfvHbzjOar/aH3SD4Gv
1gw7MQk6jhsYKvly8inDyRnlWLx/30gXAL0T2wAp8OmMkznCP7KzpgzcECBeJLRU
9llx47eFdhZrinhIvHnpKHXDO3LesrqnahwviFwaOZ2kGN9WY12W1IZVvZL3UC6E
0UsT5Wrn3pe3F9XghdYGRU9oJitQUzhMymwyLYzKZIJSbu3lqIhd34XzLkvZDdlG
HxY4L/fyNx+qiwY7IUGqaKORVzosTCeOZslWQ155HWew2riPwT9YDPMwmfE/b1Oo
209Qa4TazroMA5rBSIvFxyXTcc/cuF7DEhXukVdMS6zCXDcW+p18/r5HR1VGE2C4
GjAZ8whWMtDqMfpeLexoNyesKlQviSThA/y3znrrllQovlLz0Zj3cgcGb/jIF2nc
/4ZXeBbn58LAxma/eZkZ3EPh3pSvfaS7+o8XX4VjgVEPeQYwmW/b7j+CQGzPZJZP
2syEt8BG30i+MtrmAGuV8Rk8fXiF3etk6DrRSc0jHYLUaXpk40P8TKoJsBB6weFo
kFbS66ptQ0B7tjX+Lu67NY13EnvEDggddfd5i6LFST/f7cBtEqFLZOUtAoKztrqH
bbgFNkWjQGinZ+1iTYw0vLB8p0Q919Hu6ui/JC+Uliw+Shg4PCy8pgEis1TAHTbJ
TlnTdUIbeKHrVT8krdCJETBpNj0bkIfaeDY0sRkKoMjW/w1udaJN/70Iwyzk4x/c
n6loHW7BJk1RBpuSALdEcg6rD1e8UsbK1prkutB77aOg1UlsA5JnHOzU/wugYJvU
xswCEm1ATeQEn0An3b8lAyH6bJ8icy+ADRef9UcK1urjurGzPhWY8hrk1hxYqr6p
wP08D6kcwneOQ9AqGdeURqbo45N8cMh759cN0euNbI4g/NF/uu5Vcqp1HlBLCamw
puCJs40YduPoQNZvIHGZ+yceaaWjz/lzlWGOpHRD7Ftus8C3qW/mnSK2VguJKqlf
L5CpCm2/XWc0WRLWJVoMxnGxKrUFgkMp2HWgmvAJkDimlMwP2q+YfCj7Dfe/ipdn
KwcjeR2AOuNdMnCTYqSqaNTGz4xdVrBOFd5RH7fgUu9PlRw0pSkDzUpfihT2Nakb
wbIDH7cUF2XtIoOLizSDTJ6Nj9xPW2moTScHmVilb5GDnYvcFg9TJ8Pz2HSCkRhd
W6U8hqx6D3Y1VsL/wLoYul0pf/BISPIGIKYCH9DDU4xMN9dogWlRClXfcJuvFcYa
GCc5c0DsfY393pSga4WIAMCTSDMn6rgNZ4UrBuqjb7ftxokpzVY9sxojciZrnj2F
qGr+C9jZ7yzrVioX59bn8lch6+Dgy3+tZfqmK9dDp9hFShHBHJbqpg9MX1qJDYjC
IXR/EydpKAqPz6jUwZ/7Aw0WSP6VcIxwGZZQGoNBUD/sajN6zgPN4/DZveyhPyDX
ugTfqdc3/42aqHuFeAnzUurgJqZr3qgB3893miL1A86KtQydY0PEMDuOR/+YP9zB
MLzL+9FGfcLrwcn0BOlsrYgAnEwe0iT2dMLL+b7ToK6L13Guyx3kwgPLXDBWXV2k
jbh9yYiNYOs1O18DtKlBW+GmDfYN1QLL8XKaJrV7ndzkT6zQMlubXxkiw90WdNrt
5laxx+1ZYak3Kps0aZ8J0scRJVmHKWiasraSUqKvVIaTjEDBUR1CukytmtKl8I3O
lEExpUPhrL2rLhUUtIy0yLhDYmUsp1pMWRceIDy3t+Eo2ghHV0HWzu3jc3UHRHRc
SjGwcc9u4JKFvyshFy5cJQiur29pOG8SarXUwG4ROc/M5aEoh7CPD0BMFMS3u73b
CiYehbPSPuy+3MMoSPU1iUEPztQa9Ow1YscGmlJlsekrbl6yWM6lk5eyMq2KDPBt
GwrFXX/q0d9S3Ddvs6QoHnoCjW5GrXgkWn9mHBEj+bdAOPZwD66cqgHa6tN/Rqn7
S2OpXYfh2c1cL+xdxJEMxU4uYEKiyvRcbsaxs/fSAPomIOWLEvAIb/mCnYaJ/zAh
E5hMN1IxYK/H9IuQI3PZkQeqOQKRA6Wh7GU7rppAJiH8hrYA6vgbyJl+Qo+th7G1
XZQvItF8E9onimMy7gKo8pkE+1jbgKP5cYf4+1m1HrPzfvikIJE46mByH8U1v9rq
1pL7Zvol5TD9GMadvcwZfDQoMHogf3m5Tqr12qSmGwNjazBm5fgWR6cJqpcCsq4k
87n2XTu2u0lO/HAzs7bZIDRPnZ3pWWK1C9r7rMB+0wg94EJLMYgsobxI959JbNE/
pkOB5LWS1eyP7jlQPC2InMBb0fdbLUDIfs17fOhU2+v7tivZA7oYWtXTjZKyiZth
xCEcxmhXIjPxmowcIvh0QN0JwXZQbc3UAHbTALe7LjGE8XZ6RKlP1mKbbrruhivT
NH4UDyJB3R/pYkL+Hg/KflumeMIRP/rgOnBuAhceHeqGKhHxZFpzAeg/3e0YsmDq
TdZSP2jdSpy4rlctciMTnWo6tHbo7Iw8F6KmmByX+X0bndEj5AgHHeaSgdIYkgK1
FnM5hyMx753khp7DI2jE9uQ18a5zXF0sRV8vllRSkhpbRshayIcgfhQk0scI3r2R
bq8PzFkIHBYjur5GeNQ/tDFpDh1VVoD35z8N5xGZlCzNMVHCC+qmg4iMWA23kkj2
OgHXPOII7u+4iOFAiMXjVOd8oH/05qwSD474cBE4xnZEGumSK/XWYPYHHY3kvxG2
OyjZC1W2mLOX1zKBJ4jM9PEduWQq5K1MwCYManoYq2v4kGneunlCsqVUSChESKmp
o4FIowWRoh3DWMnfrZ/cCvqPa6i1ODI+iF7ond7xXFQKr/RBdAwQ3uJCFVjQv6tx
p3mJwVI5hd16JlvaRzKjPGuI7PeEV3DHE8HkCktd6JW8RwwndcDseDqjFkLU0J0x
hxMwRqgHi8Q0WonDZ0cl6CdbXqHNejZeWMgw1ajkemFLpMDMajzA+SVwGLDUPOdK
bk+ZzaSaCvFT4G4MFN7HYK3Ty2/llPEaUDzbFiTpoHFq4uGq4C+1kioF/Xg7OMGw
LcnHxBfMdCeFJfZrlTU5E0/5vwz6vn3UQrB3XhRKVveFX7mX1ciGLjwaP2eYB6EW
+L1kCBLUXdJV7OzoXSfHXd9hf3YszeEGzZ5LmB5mZchjEg4WfbQE79kTg3CYB0dQ
iEiVx73pgcpyAJ30nE2JpHbCSXukwNkPsQIe9Ul9lW30P168PlPqWB+NBebjNDIv
9SpmQ+hyd875ygt8JAUnBX7Gpx9cQIifHj69Q+C+tG2rFj5H4I6S4zWkwmjK1+Ah
JCGW6xu7mMlz568TzpddDeGmJD+yrAY4UySA5uT1ybmb1zN4l0emAw/a6ZPu5Rr6
djwcyYlE3zVv1flTtVOUxmm03Ky4KiP/dD7JJHQNYbckD6nBIk6jsVnoDN6FdwlT
o0Q0eIZxpbmcrUJjrHMrLPB0hiydJzL0ltWO13vQM3kcuBRVJb+OXU7zPPo6YVSR
A4d1dhQwn8iAMaERp0mPVFOo0Z0FRFPqXd4gMrcmFLJdBNxNNTR7f+YLm7ebYgDv
hTkHROrliOsTIJsqjxOn/pPRiLOIGvHFN95lXCU2vwqxOexjkDCU8jCU9nTKF0Vf
7W2DPlqrRCXpZtdJSNc5V09OKSB7uScoDBe9qD7o3HoCizHzym6MYkP/S3IJaUPy
1ccv9RAEvPOPJDz34VEz21TduxuYEm5ge/GlDzCK5uPS4u1wulbSVSQ7oTJkX2Q4
SAgPRSXY2MgNoCkNvc6rZXmb+SZhVr4yFte+mTTbTyeh39V6YfXfr5ugCz7L+sOm
WSEN+yfDoK0DeY3LveC/EAVRP0X6OW7UujIm313O654oGxoMc5iKiPnh72vNEEtk
cMYeQwbKlnY3ic2QMxGDOBIZL491z0dPg9N6x8dZKPrBYK9v389r8dSqjJ5GAFSI
MBklTbUaSQupfw4IMo8LEZFbntDYFIA7JodrYpAbHmwzjNyI6nBOCycVgq0nQSCL
fbhJlufwMm1GRizfuSgFSVVy1Mn9lqSpj1nFZQ8dUQwEoOzmmdNOCLpMf05DTEpA
WWUn7TUjovN2AacQWgF/6pUM5Tez/uusMgm+ZfHwkJ3latFdkYpZZS4x05l6MHDQ
rItikVmTUsaBrMoLF7L7/cXEPkKkxzVc9x/6JiYtkbWnsC7+ReVhMu4d+IT5dKac
PIFTDPbO6CxehDT9/br+UFmiE14QMG/JIcG2PgPes8u1E1BlY4Zh2LoU3nNDPn/A
0G3v5f1I920Aao3jpOZJXFYuHViI/iEQDdcAgvM1Y9Z+23prptBCiGYe+xZIna/D
nIsVE2Eq9mzyB98wE4rfHBk+GIaMN+6JcJIC0y8bP/iEodMDeUHrHZg9Bm+B1Rfw
VCZJBIPJdEald4twbkLngVP3QZ9tRovAB7m4G4dGXJxltMti7av0UbxVDEo9ZEIV
YkLT+7u+SixkSCJe6DdH8O7vfdaBJ5WHoCX9+Wmzw9LcHoiw//wyRD0r6+wa2MkK
IJnQ1G8q7I7pvwot7xuOcMCPETm3sLBA2dt6BzTuZll2LkluO3tbN0oHHxpM0jRx
Ch9DD367IbA42jEJ4j0jZny2a+XEf4t7sITEQQR63OFsUrL/D+GV0xvJnTJwSgtv
4a4Xu1o1/YEZWcnS42N6Hb/Muh+kGDQRnIC6JuOGgVt2X87aC5ngJbCsc1TbKeLt
vteT7EsXUV9WXo+xfB5ZYoYxdcXmy9sG3QrMgzBkZM9T48byQhgHd76W8kfa+VIZ
L7WC4WKaYxuRT7OgoclwxNIa0oIRf8yKyoDf5gId8WcxGBcB/u1rlW0ueBIr+Jsx
tTyn6wW1f5YqHtjYGy85wyxpXNts4RgWPjCfZyJ0StHmXEEXXuXW1VFJNKVCOEbZ
8ZYTh7XHy1K2OZ2VXNzo0up3jfnjvicohuycvSVGe+0cmw1E6GK1QjC+w+5ONHdV
gl8QuF/v/8Fb/ioEYoMCH3S9WPLKuQYufbRraV7KcANG/+syw0OvTBQCZfzI/QB2
cN4/WQAv3Gk7Y+423eLhlR6Oke33LzK9t8h1+oa40/1bmqI7ssZ7fv2CZ+9VcSFP
4CJbNnI0LJkVB/eLvXKZl4YAadDxRr2vH9ZvOXSV1CAnoNUJuO+zmQHNeS3eavu0
2wHIazbVuYUTP7IHJMeOa+MOtjgPJvfKpudWzp41LU5vOrKeVrzn5BYptFp7kl1H
vyk3nvVCNSU4q4m3tWVnHUDqZfdpJvaqSXFcJH1isfmyiS5URruDYeF68uTlNXVX
/5o6dh9cPQnnftbVaRa3FJSmYFzcS30ofE2ZLKVK82IoGsZXzHSnwz1LWTSuwCJ0
Fj/be3f1LZI8PiJTXpq2dd5e2/EMd+/CeivP4LBlllJzXmdCul2Yx/PeyAQdV7EQ
Pbd1jMux66pxynCVixTY8OZico5UqpzCJ1sJ6mBFHaAQtw8ERKUUMW73BFeDRvTf
ThdqZc5OR94KXFKnnDs+bfA29gDKhgnzflbfI7dLCpZWTrOY2P4JH78XVCLrC6PY
+FwmVyuIaNcCN/g489XJwIndgfAYf5RpudWnCOiV0AI1ErnKoUTVxfP7rn6vmk9j
y5EQfb7L3lKdJe+eifn4n3wr1eDat2vyW9SIdjQ6YVtuWuK1MNAJomNNhyRJUFZw
OMnBpv8+JKUDPX1nYxoJI0HuVlJlBymVmGeZhnQLoo0Juy/F56puTemUJwL8Sa4K
vEAS8/U7EuHiYhqftRj5k9831SnEA+J3RLadkkL+Q/HKbQLuuw1Pc5szSJsAUBMz
Hb6WLETk3VPrmK/yznFwVpIUzGsg4oB7E0AgwFBOwFxDGcyPCoMvj5hGR4tQ6YOP
fxr+tYLBJ5bl31QKvz3OU5UDJV+29TtuM4pREz5Q8RH+oUm9rqkJNZSavPLppMpc
/avD3/j/OHvCKTkVAjBQlDk+V0qFRe0AOVFAOdXZTvardhAJMmOadUaPfply8buv
Tgb59UCzGBYo0yhT3uB9T9SVqCqizKMrMUj1WspEsiL84Mi3nRbv9L9ANHb6cjJ8
F1tmHQpaCWGVNBlwBnFtISCQbC73zi4MWkxZo2KQ7E5nMlp7PCysCzE355qtP5Kr
mYhGAPMgIt3dmnwrADShqagekgkFwjjyk97HtpYc+Iw6NolyP/I7TzQp9G3fT5hq
3Z4LZcY9mvEM6dmEl0neNIEECNOW2sBmrxec8DkfiSCEFjcRRhCGcj8Hn/yCUGVY
OUw3wbkIfjEUU3EDY1zlnJrr1RXaEKvfcwktmErAGSr70R3sMnd2Ae7W5rzI5ASa
hNBXU7Jt6pROKb1235CBQvjwp0ZKbRciEkF3qT8nUCx+b6Hqf9Twpt/BSMNAVT6t
Vu0/CzWtrLkqk10Z0OD4iRCGlJo/vwVwGY6fl8jNdGuIhwABWkp11PIH84qE+w95
6TkXKd4QJjuUGpVkBTBm7s1q7xaw20lVTuwgIdk0C9SApmeG7b4NPYTcV22VJnN6
SY1y2lVtN+AhDhWfVLh+aENDQeJWrF1X/WXKolptWlHfoom2QppBv160eCWa4QGA
LkvdwsMQDHRp+SAnJZ/mXNuUWH6jk01hnr9EH8Zt8tLZngFNYSk+48jMky7dn5HU
o57p11PdXn0fqF8FYDrs5wdNvXhtjgNPs8LyuQgTCDPIbZCowfhuVGqcbBmS0dt1
3I5nLnIShXS/XbRGHdOoxACufobg8Tjb9bFOhoB1E8dDC3PlltNC36MhlDVbm/tb
eHqITRE/NDfLsIz6liqfhBWTNKDNNnuX9vSMajkMx+K7S9zxdXGVKiKILqsSUTuz
ks51ysV3G7DqqdlHF1j+EJS0ebEkHwqCMDtpvbO48A1owik2rzlqvNoFbxwZscrN
UPdgzPP6AY4ivddw3x6VCDQiIP6lYVmUyRqL9NraGfEnZWnu0FIrGWg4OfPRA+FQ
8pQsKGZlyeobVBluXh61Dh3IKxGlSrIurpqdq9jL7NQFlHV8qzPh4+XhCkTtq0ed
FGR8bBA0AIeQoJKvWPvsIR74BpQiyuUjD0LytUlvuSA49G8qANK4KEnkWVlW5fcy
yJPUBUdbz4+t1bHhc20IHhDCouO+eVfO+X3XPJ1WHxkELXUAfKGFuQoQ12BorZj3
IqXef/7Hiyl36IzlaApVbgTKAslRW80ZkR45TB7Xb/dwGboqeWyyKlTU7161Qc5E
uEerZuI/R3SZSx6PbomL3DwRSbP7J+4RLOj657org3mIG09H3u6m/VAugKTMlZMO
fcxW6AuWA0/80VvAH1iM2kWtuKWwNRnSzyCAelHWZnadcpsfHAirnHVXcBwKcCkp
Rlj9/9RZPHQybFPupFI9XiB2xwMBs6iISHM2wXDSD3MpvU45KSBZVCk+oRDknbHv
8596KrArcqjHuyc2uZuBz55oJyxrXJ8UtSM3FAOdM2a2qJGoE+b1nkz5r2NAcV9H
MrNYJQQpkjOfDTjWgAj4FRHTLfxXx7B34HbbxuiB7L7wTfKVzuBtGQjVmzLdSVub
OBM3cksvq9YPKHFCtVORyzm2zWLCAt/1Eot0Q5jmylJreE1LtIa8fsfayzfo0Mao
WKmSLb8HktyUTxCJACeMm7ztbprG5/dXy+ndRpTV4eHoR0bx9H6CNuliZTRj71YR
nTSO6xKzW8pMUXDh6OmzmM+/o3aA1YmXzmdxhjxR1WxSxMxLI0mOjMI70SWAQ6+e
Cw7FDnC30waM3hhcfTcP1hjw7IsZrfXbJTP4Fybi9JNp7pwm1m4m82jPOY2zeEYo
cgioohuQbaXLXdDjyoPim8hqsAkPO4ccWgX5l3F8KMJy8O5qb4ArhRlpT34MfQjs
O9Hp29F8xlC97WDONY43r0WsygESZAI/pt/ZsN8/yzy4AHFFsG7/UaHaeVEN0g4h
Ij8z9zkZ0FJKK472KavvVmeOl4Lszf3bNqy9VQ8FI1mzYWZwxk9nGrMff6hlOobc
46GMIGS5dmajos8jF8XSAMmreBJVJ/xMvZNQvrRyLVTJV+9DxSMahwaIHuKS/N36
H4PiML4/oNYBJFZzuIUyXwJGB210UOqtEfqis25K0N2/aRg6fbbfve0/LMxJmEwJ
Wj2Ld5ZRM4aC1rvHkO05kLrhR5TlVDGFI+X8SB5WpWfUlw81xL/LIl4+ihwdvjlX
Ub9XOb6aQaHhpZ0HFOITIkiXlASdSt1T9N6q0CHZXfdzAj+bBUz2KbnIl1pN7yqn
2CQBzHx3MyGjig0Vopa9NWQCm/eD1suCPWQ4Kau2qSS74OmlBuzhOwS/AfNeWrk7
kHhEqYBffSbuuUOrccCv5gAiZ1RSrk3BhO0aP2y6P27MQ1/CYKEQ4+hbZLC9vJVT
7LTR5D/LVodAlt2OQPs55qPyb1tton/SpLY4J361iU9WMcB2W9OCVPDjJM//mLEC
K/mpcW+GfYU8cdP544nt6MweA5HzzmkJTnQX1OX1Q+y0wLzrPrfvz8EmaD06VrKt
alOyyx0V31VgQ1TUy2phZnYlGVJZWynQKHDOUsf9rmHHXzcXNK/w4XswELBZKbEq
2oGShCSQKWKvdcApxlp0RF2KzPnpYp2kyCSwvNJXea5x9Mmi9N2VdT3JRAFsN4M5
WbrwPSwFgjRrf2x2hhhWxMty/V9QUUOlrca+0cKbHv5KbIiz4ptO1qKNu6VSZDom
6Q+m3/KpZRjzFId6QhpU5ssGT+9AQiiJ92TaVfoavvZS2rdYBTP+tpTeZZT6Njm9
+HpU4bNKZwajxE2gNtZ5EHPe8qYDBsFb+jTDS0m1X8A6Vk1W+Uj/DhNxll3vrPxt
z5Jvybl7mRe411qgDBngP3kBKKPDR4J7bKoDru9jH1evKzmrVEPAkPWlPDNUWJD/
ocd23eRhtSEOUtn7PmAypuFYXLNM4t125+BvCXVW6rIJ02H7EpN7rRxIzvzTzQ3a
8+KAuhvloM6GJ5fQOPcJyNs0j6MOvH+ow8cS8oY1qSLxgIpjp9Dhkh25t75vvmhm
J6CooiQ/0RqK/NgyHmEYVRokmAH9YXRE9ewDtZ2ElAQ+7A7A9eH0ZyUnNlccYU9t
7VkggV3NUDkGwmxsOnmIIsPhjIOaj7jGwCST/TFTJhlg9LSinoPGEarX6RuUqNgk
8Y4wdFwo4EPM/mI40gjfcDfhcVi6RIzEx6e7TOIwM13Ja07eKr2pWjyU47cZ3u0/
tgTXkhSDsajtm6oiLYO5rQ8TEyHwHpB8k+VTm0smHZHPqmLuAPBZKAFlAXkGcRgs
0J/Q/9UaAAsgzeo+2Q5N5/gCbHIxZOT8bEnB7Pm6s1LUiGgykbC8CPsM5w52VgQk
i0wSSnwxp0FOgD0cyInllu0cJH+rNV4GpIH8Dx4ZmJkwJaULXz4ToNf7UWh8UGxN
Au9zV6yRMKWggi6t2Ys8sPwF6snzBVdE2O00l+B2ZsNMr/Td5GMFOwu9uTrFYhv2
1rt086m1qGj0V8AsJjP+VRfGM7Y1oz9lPbuJu+I5lLc/L5dVA4hpD7B5NIx2tu7f
IFYMzWIzZIy1RvACXaJj3SlLNyW6O76VE0F0d9o/EamYPt2BzMQ3I6fXw4jhMbKd
AgOrrXszvMJNd/BwX30dz5+wnyfJZbHc/c+R2KP/cfny5ybpot22btn3vCGv4Oso
OT24MkMziBYieeIM7NbEtk2uB6flEfItffuQmJvSTExzr1Y4SJLDyxX4C9YeTm8V
SjRznYeKdMPSXDNSS4SdtnI0/BN0oDMKRm7vwxDHPhCUDlGGJzvBdj2bsohF2s+C
XLdTQk8tcNKoYAqcDDtrdtxNufZ2t7uUA6KyKR/I+pYh9l/Iyvk4ym5yk/73Uphp
TC+QOru+TDbYKTgNXKshydLtTBJfBSgHz5Z9e9LUcxubxdhx7SxLp2sk/b5hnu56
+0Oamo9WZ05LGuhkjZSd75UznagiY+UhV24DhhpaJNxEIjqG4WGWcfyRvJcSOUgs
2mWGXcQ84uAyN+H/zZHCY+Me+Wz1eroTrASC3QPCghHGuCaEicYzPuokStTrsYAN
lJ/U8E+Js8u7LQ2pIWtPbXU92bg57be/r9G9DTenmmnaYGMBkQJhkM4TX4fGRjj9
as6eT/rlvMTn99xisSFBLcoYEIJWhazHeB+9pttn9Zyw59NSPZfs0VIaUL7PFZck
3mhOirdnFEf8S9aui0RPL26AKNc7PqpiQfAPSIqO0KflxUjMaoXbthGI/06VdgD4
Z/SuBJ2drQGC0TIRLx70Y6YIg4Mcem/tTUqkyqDKFMmXa08vYW3MilcYzkLtLnO7
wBLUXIxTIqOjiKXBEYfoDjxE9gdMqKk3k7iaN1zhIpgkkpWgWCh5vFWuYS/oO4vL
NZK8IjpK0xZRxsTgGRGN1SCZBxPoC5QuUOfMTJOkitdl9IzbmkBG9faf9WB+F4+1
gEWDWe/O7bGXGDVG++Zp9fAZV3YHffuM84UDCJpqzhTcHjHMfwdD5jTE5SEPmWps
W2//yy77MtUYkzI8HzYtYcncp88HzNavIN2C6XY7+JVlXFHMu/hbFlOixcEh23Rb
+Es0HBJGvjzzt7CjUIGkvGZNCRGweHGl6U6QB0u/8e2BAG83FBCSuTUJ6K5ejuW0
kKRgSFZccYydj7zOeNtAtV8/kyQv6WFtBdnqckGF3QI25dDYBC9ZxDpaCKqft53E
GWQsv7skd8yGkUdmjvGSJRNmkJbHmql4pBEVC/qaT3c6Dp4Yn9yE4Ttx3GdmW31l
iLMNj2fvx1EVRhpYqNUg3BV7abhtcBjAt/5xNGodHpi8Cs+mXeCh4xy8vI4xnXXc
+MPD3ggn72azjs4gUG3FOPb5M5QnHM2Isr9Zx2euca5aM5DdProJQtTxsJ3l8WMN
nfsBg7+gHPeh1la+sWjyz1kccSCcEodCT9kHSE2aVCRwtWt+fSc+LFD6SK3e0MQh
N9JpK6sWC9O3lCaLVqYCAnoC3AJc/pDfu06twvg5cXvRTEPGNN5zF5igqNlUgfC3
gqUA51KWGa6PQYEbsF7+3/ImhPvIgZCQx72twxLggx7mGhMRMGY8PKTiZGD5LvW9
Aeek7LAr1WUfvdJ9ZRJ6bFLy30dmJeqTFAU2qlncbol7GGWahuSkDgu9UT85HDDd
cT4J47l8jQcvVcReEJn0DaGyh1flheJex/RaDp0C3Nz/89hbjUr5r7i3mTmJ0+QZ
c+2++DbYpGNLJvx7K70cLTvzTzV8NBqQBGbZ9cNglsBg4uhtKHJhbfjql38o9JwZ
bzRztQBS+7W178AwPZ+91FN3G5XYPnCyjo/RR1eHj6ux73Pg1jw7vJhusCvCdQSg
MyrhHOw9b2m4Tn/xuUh87ZI0AXT74+IsQaEeJkOEL46XEMjLPTZieIxjmfrbiG1y
+blF/7zbUlBxtA2AjFTAi7ymHP8WKvrZsf1MV2EtlD4N1lN8rcLcT8Par6kxpwlA
LfK464Bvr5kFKZ62Gpto+6uM8U37p5pRvT8oWikEpglNj/W4EJ30Xd8+MLUfiDME
y575dXVRc+Q41xvZKUU9WWSVJBHdfQ5NKkoAKh7thQoqnUS6qkcsIr0/G1rW6rqc
smsgQKUT+W6drJ1i2SQHD55aXETJK8fpyDEKqFdBjEUbPXjb1MrfyZWdpN9VgPrh
mDY01WMIrDP6pZdRPT0jc2Iz7HW3cMg8+Oo9ZOPndesJRVVFssYUGitnAs+EtZXu
mbpPntispGtP6NQZRglf1XShl17c8NDFo99yhukHAtoUYW1iGk/7B8vQ/ATmQOZK
UnoFlVS+bD6/ervU3GY1z04TEHEVEosXyeqUZEG1lkPEWNGY7Gi5K4WaYAnzcJnJ
Ecey1lUqWF81t23UqmYl6gt6ktDyQ3JqVtdQknezZmvDKUQHWC2jt+ufK3MPIPuK
gHQHyVvXWQRRc/nOZUAW2ceimATKGEK2FE/L72rHdT8kljqfvDBvnZpv7UHImKKY
BQeTuY3TWagZq8yRKC5QTIgjnpMHGeAcX/LELshdqWSBkpwg9bobd5Lp/3WTj9Ci
zVaztdBlG5soakTLf4FBkQKvnDzTA7xSzZcOelbbdJsPo4y424dtNq+8UFONuuLG
SwIyoenZCX98sB+ULXKDV9qcFulKvfqwP3Jklb9xa1DbgaxnfNc/jtER8XrtHOWQ
iHE5wMc6msxHOpG3bQtZUj6OfsGiXFBoGgvn6tvZrYdqE6xekERrxPlj0b+SPqqt
wQC5QluqdwbFHw99+rGCYFwpck4Y2hJXJ0GIFnpDdXkQPUkTRjn1Z/viyJN83LE3
T43iFjIZyUhG7Kl5y7qwB7ZsAziUSup65vVkiKzNXpM3v6WKwFg4cI2dp3rO2jeD
oepQ9BPSvLOKLivdCdq4FcEZpY/rhmyZLXsay8kUlxgXjuX1FccBlQ3gS7iEaWOZ
xsWWUpA+tfRKq2W/JMz+rR2uYPojiogZlAcs72qjemGP7Dqyu914SwgPhINQBZEv
53Fcn0EO3CWSkKCdowcsVjXHVdRpi4EoSv1bECa5hA79KKQtMmGiU9VqLh3EeLcF
ij1EwF2e/WVhzRHffGYyPvpJY42QyFMpQwPMGF4QJn/ib2sXV6R7i9DBKV+FX7XV
ZXbSwoyxA5yYJYuN7oJ09wmyTpuJQ+4yKkOtiGdwAD1vo3nAZEb68awXKzUSs6ai
2rIcq5QBM9G1xNDZrB9B7fbW+kdiDTDlR+0QF9mKqdiVSfY3/GDRyoyBPww7iNno
OpjD1jW1k5iMiOwHxh/BW2ASaXCU0hn4XW5wXvZtpIilhu40ptXu0bYQeN57rsCf
z/X7isqtl/6ULZexl9K125UNrl/S+yCwcIJyRdAA/tHL8qIByoXTXYw8Gd88tfAS
61zNhYoq2/j6iOdK3zWY1JHq5deonnR5/dactN8D2sxVnXjTldB3ukgNascaOv+E
42RYdc7bn2O/gMCnfKws6ve9hSBzeDquF0AYA7YiKe7hAiUoVTBlujY+dEJ0jSKl
E1S3Ez46s/GUkty2r57V8gDw8WI1Kj7Jt0uhhYvGAzKsJw5I/+O6FhtI2z7seoIN
8JxkrDEOYN6licmDE51SscQO/GAKWkYXfRPTEVMkoWSDQiZ8dxttDbYOz0l0aMG1
iTRO1QRlaRgbQCZgj/u43y/0xMnGHlKFp3ZF9O3qwUeHJcKHYtNEkBLzN5bKuRLJ
LkVu9qZts2czxePr/ueDbkDMpMuitR01TtKKn7B+D7zxoM2Vuz69DI1QsT+02JNZ
zuJRi9r1VXAG9562MUd31QZJ3qSP+kHlf4zGDxjCXay2l9BeRkkbTIfSYxG0qqlu
CNvcTNQ7bYUxvGKT6PfBnXeJM1sSoSHnFdKUxyq+2M6Cyh88NmWElZ2QYvjN2xas
srVNEwM7c6d0NKr+3W5k+2L6SICAemG6v2DaB+F1An6S+oDZX9lAf5Yhg04Gt7QR
JW0SSzn2iKIKvS+r0Bah6dybDn6w/TRLOhyV5T8OdZd+KGGmzaWUFWYeZPpcPXU5
wzndww0Yu/PnmGV6CkJR4yIHNawXm2JBhuH9WIxmo9Dv4llVYIENFjnCD72O+Opk
1kZjfq2k3KPONqvZ674eDCOIaT8X9CqFPqhDwzMK8AW4yNVmbNfn8ZLvTpereYjI
6JOspQHgiRQiBc1cyByUPNYTe70WyjGmcfGP3vxaqvWrbu/GNREVLjAArXp+1LRp
om2XGgxJ7NpwAj6JkCfCQwAOivlAr3FhLvbFi90HRS0sxePQLBxgHEKO9CY8mK5q
7lMILBlIQZvYDb3Pcy4VY1YDUkh23y4gO6F5o5YbX7Lg7gc79ZtB+IvXRpdMdiry
LdRn2NwDFu9/hxppETuXIx7E6LL74HdCS9LKg2y57EWxZHo5AtmkCV9ixYSURqvF
uH1aW3Kp6hpUVBhwKI7XCIVt6THoSOwuypO2CR1jUVbIGEqQ4cux+Oy4I4CD2bdP
2ywF487sBHscflRsLCviIqOCdIxGo9JTriEJv2NjhQNITPRIxrKx9iPOdo260zP7
Ls6l015E5NVOAmhOkYfp5ZaV6Bbt7mivvPGkTWiTUxVrsYAv6vMKC/PXn8zte2+J
jwZ9LOG4rp58oFH5HR4ZVZXfZOYGSswEC0Pl5Xy/hHlq5zX08XBeWpVxpoUSBjJH
AkIehUbkPIW0RoZBKs7eog6HXiZeeVmfOTbB4QcUzMyWJ8SNQS6QKSgnb2Lp5qdC
EComFf1vQPGSwHs4Vr/eztySSczCigag8NjkbV2If/5dzyZkwN4xiqzDi/F0R0+7
ShtShwgPgpEJGv4bHkFe8iKvJpy4DV2IEeRLt2rqf1skgcdBAvmm1+yNJTgqxX1b
Ps/4g8fSVv705r1fZrxZpyKm5wySEIZJleCS0RbaULwtllh3HqqfLSmU3i+2mB0m
dEhezkfP0w63+B/e9Df/sG92334E2uQSnd98lRtgdDAHzZLo6BwA+s9BlCISyOJW
pz1NVQQ15oB7ijDcVM5nu8r4td7/dvweturqlED3IxCSCKymMdwbQK2sIrO4GdIK
68eJsR/TW+HT7ixvoSe7zBHJSMywfzuLhclqq4ilShU0SI8E7dbar8S+eP5jSG0G
29Yr0OvCxHXUf5HiSRSWxnn+ExnLSVyAXJ1wpZX1GHlllBgJsC47gxClR/8cCzHy
gdDl8m83qa//VwqQ1w1xMUcbb5kkyUt2+ZjncAQBzGUtpyYzwsH1eHAEobDvHqZW
v4u9nNQ2m63zcK3pSFR5S+8OCCzjEWyID7i4TlajhLCSeUMFXpaR6TCWmhJpoB+6
WWq8rq3dHOrC6xt5/clWv9ZvoyBLadRkgaFSN0AR1JqI01dRWhyo9oejOqeLmPT3
DhXKVe+toduvFJB+Zq6u1lHCP4tZ2Q8VjwM61FgEOxbrV1+CMOdBjuRqMIddC96w
aY9RBZHPGFaCAX8nzxIZeR4yftIGPhQtZoVWflCD1JMq82C2rGsmqJgd5PHnvWeV
TZ+KEa2S7+ciXAg14R6Yet3pYyCejg7GQLdAlzrsCcdVHNPlWJ59uVSUKrxN0hMM
HiS4dKrJIiC/dCWR29xCq5hBkePPPSKylXw/aATTFaVH+WQvUZxvuroTvMM9x4/D
Kt5X0R2txYVxQ0RZcKag/ZRZvg8C7oGMBGAnUVXS/zfD5HIC0VIGCE3AnI9Oay8L
kBwyR+xHyceV/pD7nSpBGEPOhiHMhRGbd8C4m+iCJdMZ/l4xv5OFv2D+mF2b/GFU
WbzRX9hKLEIuuufCOIGG+AOFHikEA2vAyiXpsU0YdyeUOR3tOSHpwAOlPVM7g5Bf
ne5f1r7EceIhNjun6dr6hdbS+ETzh8477915zH/ODtnk2hUXB251FKjk25vUuwIc
M8Ke/4ySRLX8DfrdCDnVgTW6HF5ztwlj+39fB5acmhJi5u9RMb63/ukmpYuyt66G
MylkzVwXL8SpoiswQstEl8BS9xHu5tUCI3+6GrSbvqreawYL/PAWDepNqRAu/EzL
+4eiEK0dJgnCi4I5d1uJNoFisoZT1SSDVfabEcv61X4Wzu3QU0kGFDnQtSFSIJku
MFGosUIMEW2Ctf6fSec4xgFPwCeT0xRBbnp8K1mm3TQpX7WC6/KZhd299EH5YSQP
aOLwBfhQWCujZIE57yeXoxFqN/3TALQdE60twv8aBNxkubph2TH9CEnt7XJUluH4
cJ7Y5/o5ApecnSKAjF21EQ0NZeXOocMRPAxC8U+E409XN422a4Ab4AU2vC5gUNgT
+1O6Xp1lxz72U6j8CIMhL1+4Ro5uYfOdd9sodkTf/iyCioSxtRtj6xilUaRDiMJ+
/mZp9oUkGOo+mEcYQwmBTO9cUo1kGQF1Deim8i5vb8/ZGrYCagv5QYXUNTaDjBzL
hSwli6mziNj5/6wIiGmfo0EWGpnGPesy4Te+/V0G8wQB5u1OQvZI+PhlME2isVvy
EOYdW55/0v4uyE/w1W8ohxYKWuw0OhsFkwTUWIlszNejaW8poHu2eG7Ll/3SMKDP
0mE6MXtVyJlx3fOr43aZWd2FV3AOoLh8mUJQR0ZvzFHEzoS6Jgpmlg6fWIxQkEQ4
lQygYb262KdN6srxzZjioR+T23nmXsWG6siE5a//rB1u5N/Eq1SdfjDpw3cERM1u
FvWTi+RiSIdeAHMzlh2zBYcY9pxco9pwnLLpcojMom5a/2xnxb5cUDII34qJOW/B
U4Fk7tysvcB4wHzgrq47W/xhX7dwRSWkIw7GT8k4DbxpiLp1uhJa81QfitVclkMr
smyxB7QaUNHJEgKLXYy+XRziideG3O2ThQZCteOGA2Wmk0dfkDktSdoLqheBnhZg
sILqlaBO/Fl+lMJHVSOaN6oVaiIU8JW3S5AQ5MvtfSHzER6eWjsdZKiqi6J7BBs7
o4SEr0L1Ngss2YpCMVXjgPWS9R0yGre2VytJodjQvzISFchStX7x8Y7UV7Cbw9qr
/cUcpDSz5ZzOky6ufWeORchXEmZZeBlgCYtsVPlykogfEgOodfuLEMnUW/LcqCXp
rN4A1bEw4sByNAJHgTUMlVBEYslMm22P6wbgFxphMLxcUBMcDsd71FfzEe6y0mJq
wn02TkcBEeVtICU+jTIFihEdR34b7dGZZcFGhafC3vXMgv1NgDVBDOffETET6chJ
UqOwCQ7I2OHBHx2w2zOHw/3FdrkzDb5oz+nA08/mhVyLE+xPN2UmgC+5U8JkhvC1
DdE+HEYq0NDrMMMp9Tg2QO4F56vL/wU0RGEtLkLb9IQNSAuzxhRKVMOiIMrVPd6j
d7WOM7c5ycVCJSc5+OOm4WnIRnZFWEjX8GVzDe2EG24a5HGR0n8uIWVqK+sm8i/H
rhbQEKdWVceT/oji7AjWSSGP3jzNfvRTt2/4InRpCl78m1DEjMoclB3bpfNklW38
7qtdOHMAGjB6E/F9fclGV9x42C9xMEfugHE7BJjDKw1DelI2fjvIT0wFHSEKTOUQ
jdWaATk6j13jBtJgas+MtC1eIXND0lxObAwrN+QROqlpOTYiXufbkX5uTYtI46FL
eSXGdXhjhJstGllyftovSl6jxT/cKq+Y43kb+NNXJjMFMg5shKSIHCEA2XcGqTiA
S4s/k0k5+J6FnT1ea+CeK1MFjB7KWE/Qc4FWAbz36VFaPIv6tUjZOKoV9koNE41r
zUMUTMD2qq86+IF5kXZ4gx7aWU4KS0s94nfifon6qs7BBMog/dr0OOi4WMs1fLFe
6Q7eBkRvrYLI6PoMVdH+d1IJbTf6N4hhwtUanHkzfgVF1Eq3ysH7B7++4ml3L4aM
n0k8KKddfCdLFJZREsm0xRfT6qJ+fZoNLd+d4itIX92TBqisavRfE+VYydk09pHj
pJ/WeAAsJhxMietovXBm/Jz7PqFJeM7Zm2cAXTqJ4xz7+3SoaUUjTfchwRGAQk3L
Meunn5Xru98MZ+oUF2UTu3087ELbA114UxUpboC1h3La9PCMfjBlWOy4SgQrgJve
4bjymBPiZeyQvCqnscl+Iex16VQdEy/GT8OaNHQiGej1cMtgOVKb99F6gnZm6DD4
3PKx1mqIi6grwm4iPfFLBJsDvNxhfrS3umdoKZayqIPOmXQb4TIxZB7hsqhDCG/N
PylPjfS67hTYJF2uWBBax8plqwEuUn4wMzjOBKdvLHN83IaOATbWAE/vUdr8tGRv
W3I3ufA38LotHqt6VC10yFjD2CSuv0MAWq7JSuWtFKrlTrb5n4oI2DHc968ViLW0
znfR9CZTD0uhZwvF2o8uSjz0+5Q9wgZLyju2V3qZrdsBidV9OltKLCOZVajavkYK
hYO5gZA4SZmyc//2IsITM22sM01aNtvl85Rqg3XrcGlO8T4EuTRni9E8I9LaNFtE
qEdWTXjR90EOycAE1DktjwwVZwWjKju4C1GpiXLVBlrWdv0/P8WUccW9sTNLUgnG
jbI3SygzgeoEDyXhjyrzKOmSVdx9AASoio7t9SRkCVo7diuFS6T82UDf5rSdRRFk
EQJ3nIddlbibIDx3EjoJttZZvHbsML4CuDb/6l1WPuRJpzLRuiSr0jtRdHMcjts8
BXPIWH6TmZJtR0MNnuKwmLm5U5ttcm4v1Le6SGO2yfPLfCR91Oljf5eZhHPIJMYj
FBbMlofOSh7LWDi6qVHia7z/jasw+hlddkb1ML5IoZ+Mdf6Q3CJT+27CSZtzL7jT
20K3hmzIQDM67DUUavUdtKX8x0S+xNBaLdmlN8z4+RfXorscuCrGqp7J+0KnjLhl
8RjibPVXNUD58vvb64uwu2ZIbTvnkt6FarfkB5BgqEDsAGOjXzivCocViVFWYVAt
w0mjF469qZyGIT9a7z/KbSVg0t2ZZUV06h/7MGfIFRcEoAHXHHsB+b/Ms6URz2n5
0Jv1lXNasam+9HkGqumjy8SpENWwjUMlNOlsrxJ1TH52k/YycoaUlMp5lUB9S/mm
LhpY9CyvOXUpf6FJyJai82c/Br+vKMajx9K2HNZBoRKHNGklUd991soUDAK96IA6
fU+NBnKuZK9u6MUaKMDhPYuMybrKu9ibcYcQuQhhDt4cxxO68dyfrPvn5B/AAecn
1DG7Dt83Ip1fNe1/CpNv5GaBqarRNHoiWnRM7V2Np/dfKlfzeYDJF4dG6ZuaV47w
vqiG+yZ3aDXoEGa1MHWrJ9RULVhor4OOs07DrHUU402E1mfkiNuWY+vmyi8HTxVS
6FVaNwGms/QrOTXIyFxm10uscryPdc1f38T5Y5JoP+slo2lWgZpxq9ShH3j2hgBL
5vXFLAGk8JMI/uXrDClkuA01fZcraGuOX2KyjFaONS5NlY8izxShqxzFABxOjzaE
2u3G4RFLc9I6TwYRToa/5mAryE3s+HmlE+uahXP+8HPbS1fzV4UBWYgQJFIoyo1n
qMYdf2idDPDkWwRkBwVKjt+x3QxqwTFv3lYtqT3/l/Boj2Fc+i9nWAFOHNQVTlHv
WNZ9Lb3FyOV2kI0F3S/UEcmdWo9gnzYjrs/u4NWcvg9d+t+PtFfoedZyWv2WKHIU
A+uYof3w4V9F/efa+3XL9haDM1Jt84MgY724gc6Wk8DzxlJgpoP0h538lalRDC/D
KpxgpXHe3zCR5jij5Wa/0lNmvEvu2vmDzQKvPD7KN+gER20ig1ZShy3nyIEHmEr0
N7nHsHeyeKc0r24tk9UiMQL7bbQ6XKHp/Jwi3QvZ8fg1SMNyKJeFAnyaR2cVIr5l
XqIMP8MKCNzJ6BPPVYsEYVH+ENrFxvLVN+vTdFDPP9io5/cpYqrJZ9eyXWNzL/Lp
UhN54nJDicTZff6o42ZNNKYEozPqoTY23fHqLjp+QiuNT8L9jnJcoGZ35WEiJLZI
A8IH8Lwpn+PNP8gNovtAT74/La0KbrYOnEjnaEuBbNBqyoUn77MLhSLc79I4Knoe
2XALqoy7cazF1/FmwK16hp3B8puoEu2KLMDn7sNu1JVa8qUZ0yWETgcR8wGKpP1i
KKSRI/13EAei04oG3zbnHW94DcHC0poQe29LyOkaJBW9jWVC7b1Dq3wUxma9Ho3o
mQy+F78DZE5cSu27qyG1pdixUg0rGKJt6MXQCbHKgMAgBXDP28sutnIq4eLkbhu1
77nfUa4Z4UPQTLtOebFlxnQ8Xg+I/s25DXWllr2q5r0iZj+ICUfsBVFAHHf+24QW
Xe6M88PONzniRRhNIHIjqsAn3XmNgVUw4lGaa/uLJnsL4OcunesGhbDGNXuNzFXM
h+k1TsQY8RmrcxICYihFoHUy40sOW5Bmn3RfCC2Mmrmd6SZvsUY7c3LRmwCX/eUC
tQmcSB/zie/UIaW+QuguMykk1r8t4rLRCoMKui98D4amjj25DuFSe3ivV+pdek5C
ACHt9zXWB1ZdmU6HzJRKchWySRUynfMziZQi4XwEqux3cd2N2gbMZ1NCxl8gVddt
/X3aVvDgPFqtLedkxgL3Xm75ysqVis8rspwIqSUjH7hOc9Oxw7mtF3nHNaBaRDlq
MGDA12fNekHacsN0f+SjO+nYQAnhhETWq5JuEjkSkKwaOWRrrkixAN9+RqgccPdW
5B2CoqkNcvedQJWFIbF4yMYlJiZhGSHlD3moine7TpppjlHM93HkHo651upQjVnl
1La6pf/XqAlAE8PBtOx0/EutHS35MOo7pcX6zPxY0JNJJjHUZARq40Oc5zLqF/lr
rLZkVQp9WPKHFWAW9tl6Ic+L4NRO1VCQ+Y9GXI3Gvv74MKkom+sUxen/7hz218Pb
laqxu32df/TpKoLWajF6DtScpXAMM9Cj9vIbCLr8UC3fsDiBwE2Ype0h2E/sAtuj
0yIPF4sYSMVBosXicUA1lmQo9F8gGxDN8t4nLWrvOHAS88r9Ns97WG7GVj8zg79t
Vky3ilgiC8VYeN/NKf6HDyPcuWCVA/srjxtSI85gkfk09HzYGsnb/bsDPsyCeKGk
siVRghssNO0mGDQupp5cDD/mf4qTItd0Xbar1BJEkjZKDWpBy0vnZlk2+LKl22F1
47Z6ouR3ooaD+GDWGh2y2uPCC+UIyjKbf/R7aSgHBVjKxi8PB0pSjpzjsQnTwu3l
hV+0HcGjD/x/vddr/HQYAp0lRiliMy2UwPAeYemMKj4jcHpCFTvijqwrdDcPUXAF
XBWbBHtecnHCOqXVnMEMQzHU0U+qi0rwh/03Y01K8dWRp9fonnkmGz8pET/9BXg3
KPZQgFhez3B13X+MyWqAATTRQNFnp456YdsBtSTkF+yRMhBawPME0Y+m2tspT7EK
cCZe+wiG0NaYxWhiWfyZEd1j5KlsuuJroCoDJxOMESD4lnzLZdy0VpF68SCrrhL5
inwUDD/ezu5/vvy4THZph5Oh18X7JuZmpS/ESbGNWfWjOHmgmioe4b9+I4UlgQ/Y
gTwQRnpMmyEYm2DjYJz1lLef7FDaRDGQTW8JbAMYRPIBO+0ZaDhCQOiAbZ8dZiL5
wzf2nSfwHJFmpXiWdz2njwHYNPm8sXgymWsGPwxyoi4D96wJeDgoYdsDQnaogrYu
rNiDnBmqbWoTrE0SF+Cugq+dfGHNlk237ACPHq1+gyGLVpQWGSSAHh0UobFblmOV
fOy7dh3kwNdyY2pldDPgM3qBT+642fuowDt2wTDveGhwqE76Ul/5lApxCV+9E9zg
qjiPmdp79CHMEROIjHPY2UKoELrxG/J/N5FpolpuOglBwkbRVl5bGo20qevCkNXz
9w/m1gqiRGmTul7cuI2/IqIjuWmmx5LXmwXHcrlwOSujip+cPg4iRmpmt2lbVvF5
S2Ef3g69rDa0dmYa8vOSqaiUfBw4lzEHWVg9qjABDruf3nmlU4tKceUgY/ybPEz/
W4T40xUSxqcmLE/Wtkdy7Dp5tBh6LlpuBJrMRwnSOFUDMoLi9TCROyp54epJCYqx
mzM0NR1ypkyesH7PUwhvrJuleg7CyjVDsvN7VTWLndM/H2I62KmG+rSRGydFWzBh
RmRbmh9U6A+lcJgetC5iWnbdt125sVLJoXft7K89R12tFbKm098KNucNBlkFjTQ4
GF4ZtG0x3k6OFhqNJDlA8dEq38KQVcLPOILFpuMBwRWFeFaFMHjA+JnjQ0hL2Zxx
4A6gM7bgoEYJpdZm+2Cjx9mRhyv1xiuM2bbjTlrIP7dTufHea4aNzWM/gBKYo4tO
EODa0zOs6Kv3yJrVxRtVd8s+irNnRagLoPCBdhYfx3NfWvHZTjHBbhn0nvdGDyeF
JNryuWQu2meUHWSZ0+8HLg5g5fLO9jB6kp4HSR/xFw2NVHx7JUlHTWQ1lqQSBC0b
fwaUdbkALseX+Ce0LDPc8E0l74OW6WSdpUQo8XZc8oSsgOlSFno0UP9A5HzqsZIo
TqH7GjlWdF9t418BCX117B0naoTIeSU+7dmp77+auUcANdkVN9zBCeeD8Ijb3isl
ayj5Z+d89BNQgujkkT3N6szwW4zwgG8oQHmPn0QUZF/Cdr42TVMiwxSYklUm46PH
3WPDLDBWJxDJXl1lpTVFCwbG4YYEaDBizc7P9SwckOdryKDlwRP802H96s37wXNZ
vIPzU3K12gDIUQzgcQbmLg49ESwuF83jY+4nfKNQillw769Ev4xjVbp+kFJ+N08d
cSBVwaqwLa6qV23SlEpXHX+cQFTQazyKS+uExkCAHNpgRu2VmDG8iimybWQ74Q2y
9ktQEoUnfFBVZW4joOIFL/mNpkhttmePBx0Zq6jrw9Qh/uF18rC948P96eKdyuLi
tWPZDGAF4EwL+GMBS0xGLZhsBhFPkO8g5nbqKxPOQpDn4Ef9fsoGWt7d3EgWkxxk
ZHtuzxW6Cuaptenrfbc7S3Zq5qdDUh8xooVT+ZwHSIWekWNCu05j6EFEwmZqEsBV
6sO5o4CmHLJKBXjDDVveD1SL7EERIVwgZsTZ8fWci2h9oZihld7HfE+vD3bA6UMA
Jwf18KMxBtOyqPFgcJ2YI6ayd99Zunu0YZx6/7QMP0h/TMQZHXuNkWA5XBUy2ktS
NSLplG4XcmlvG3xy6L8tBxvJe40YcGMbZxlp0PKEhqJWf1pEwPfljRgHJXL45rJA
JEsagFTpcdaTaHsmMgW8idsOYggffJmvK6kX8roeIxhuKUdl9SoT2A0IYP6VquTn
7cPIpvRGWWD4Bkv3MfW8TL3n2qMypWza8EqioNnqGvKNIDF5YGf4NoTRUQr1E7aq
Y/1EKCLEPrcgdWrdPLZwmOVCDKWdwsaeRiUh/RGmN5K3N1lOxQZQ9fM3gfbYJCbH
IvsTNfoCbHuCEU8qwJQjXr91Bl/Hc6kGb8A2vA1hNonGwYDGBD3HQlOG41uvhCBt
8KRnLUEzsSkOw1kknO36aiq5yJRUa9Rsql/wmvw2Rz9a54jAncz6JYxvgaLrRrys
5kax2bw2vKMCmShddHrAlxTHWxrvFwLu344MTCkIOjcZfXYLoj+lP8A5ZyEmMHbQ
5/SCf1ntMPZpBNJNzhaYbfFQMr4LqhIgkEUTC8hboNYbQoiNCYN1p5uq4sWdMy54
kkkSvp1+KnW+guUB+ytxiWlDt23iLfDptzAXwbi3vL3nPDwgrb+5FterCCIZ0EDX
mRS8rOjxjbk/3EZyO+uqipiTfXEekt7/098GU5kHNz+Ium07S3G2aGU9r4bBYhdl
lvSMf7qo5B8DDHRtKZ9e4uGkN9JObMAl2BONaVBZoK8sKE8xCSHpiXF9F4tZuJFc
p3y9/Q1zOHT/eTqv9PeWnaBqiztDwcOq19upYyufGJO5qw4KE3P0HCT9nhk6XE9J
iVjhCXI4Ra31Oyt2UHdqDge4GHaLOy4D1K+O6afRUy3FyRvIGzkJ6FVVKVy1EE2T
hLezoE6dqte895vTG8T36ENHID/DBpQISjHRxaVJhIIAIqs4m2YGb1QYk8/1GXPg
aEGCJnEJk9AJIXwhHqqTQoOMwGnQ+9OzKBxKO+T4dq0r21DH7oh8GT6aRo3Fx/AY
mCRjPBSAOqVTv3JOvDN2ZM0bB7w59b6kdaBq3DAQNstCNuIy19I6+XfRaRHnyABj
zKWNElD/9M1HN7tpo8Ioloh3Vs8njCVtczHzZeFcsGjG9sT+GLoW44k2cVVnJ6vp
etkQjBjiGUyOwcxuEBTMUzJsrCDWUjkgMzRmZa86Xhpu97/GGMoj3uiubXVQ9J3r
RrQmzpOlZot1pLyTXcJaftjGeAhVR+9hzSEQHIp98JaOWaTQnAvCWhdpFjgjUfvF
PaerECNP4Qk8aGfrvRLCYg5ce8Ft0K6Zy8+mVkQC0x7Xw/rESjXGqWXl2FDiSkPw
3kT6OA8P3DIfzK7HoNV8TCyjRus8dN6Oqio/UzdPv+/r/SPc7KddhZP7MQ1AJJW1
OnAsIJQW27sjFFV7KmT6cORe0aDUqDsUjr/ywvsRAzySXeKBQYgUF+JQLxym6/H6
WgL6yHDYq1zYPVX8K8hTLFGNrxVll0rzwZj4eVWqh1SRUhe2KX3K0/zccide6G/Q
URYDVodyD+QzH9IIUh/CYliDgiJG3gWBusoGBUXMceC7jLg0imOzDDETGHIamtK5
/S96TpaeXcjhF7mGNzxUd3H/H5VpxTgqlVvsH+nFKItUEGAmfsycAKuetJMkFwMm
P2qa/iwIDHBebF44MKnxePr/P6rShXsc1qEfeOdtxt+d0SdMsJa+kuld3DOa5jv1
5rEjDHz/IprROHHGASruuxozxDLbxpU9H12dXXAQh7bKp65lomtUwerh5K4p3n9O
zTFXlX8NmcjKdZxTsUZK1hRoEenb1us/lmUJMd/68uaSoptJw6q16P3oaRj0AL0B
n25cveS6Hj8UwiwIz+tl+u+R31URv8MEGzFGc/F3YcRGMCw3h+u8GUdrYaLFd1Rv
uXKxXvw9q6ZkFF9xmOlo+wStZOFrr9hVmfp1xad4xWf+dIisHCz8JTE4KkUz+xdF
ixMqc8Dr6H8hqYfPNQXzXGAx9tZkoMrUa6Fde+N3oTXAq3qewb70Puk//uYYCfkX
aRW+5jOBcdEuJ66oGIh4RgD7U3reTEGSugd7c1jCmw7h0mYyAH9A2/lZlckryCmx
O351gyAyIHZzWIOUG2DkI6hjZCipousT8H9s3J09ZaYleoasp4pS/C3eEsG8OlZ0
b01zHXdWEeZBrkjFXLGfGL9dNiBiasOJHTqRNpamLLS0a6SN6c0nHxeWn/ztWfAE
MIX3MknvlIQlqYKTM2k4Cy11BpKXsOhNMmiPlkN2tLWWrhpT+xXD9M8RmMn+guGw
tzUgGaja3Ef8B893je8Mk9N87AZVK+EHIlExQ7H0+tnYP9tc2ck4btB8oHLQX938
8avSkknto3mRXZHTaSdTxr1F4qKxIaUKqS72jfD4IlxizKm0xCpUm9u6xQOLdgVr
pvbgXpI5CUip4VorzljipEmGyeCu0SrRrCV7YNoar26mt5pZXwyNx9cGwex7w5Q+
Z2WEa7OgbG5YSjyItFFw4pLkRsL0Q8leePk5ElfYQpyjuMSeD1SB3Gwi7Ssdq/0o
o15nahHcDRMC/vlneeMwtgfL2HFk4lTU9fiu/qJJT82RxT+RJIMDCwuwsdmZh0gu
jdVE6J2z9p9tNhPaG0ZvJxECVq1nx15fEdMs/TZM9/M5+34/6ub2xvWlNVFD9NcE
8syV3vR4rR9BhSKivua5ByneW5ngW2dH9+FngkclN9uNdXqKPeF1oKBCOxO21Nx9
86XI9i4G0Mj1zkYM7RX1cyykaoh5zQv7GArSEP1Yj1pwoitBWwpptb5cTTZmljmq
aRmxOauBZ5oyQ4yr5b2qx3Ry8uFPi3OSCkt5WfpLJJvllNlosUKoqgcFr/rphGo0
mG8S8ccnUK7AL8Ah2hKraVg4O+6ayCkt+5mopIStBvoZZ6qfMc94CkNhfKs3pL3D
tpjIVV1cQ00MepxOdU5mevyc/Fse6XGsKeLbYQfDLT5zogYjE95rdj3hGaNoG2QL
fRd7SfXv85hoh29yd+ftKAqq5m0X+cGStx3ntl/00Xgo4gdSynysjy5fEFL1tjuI
2RdTaDJhVOQMLD00ErEIxCvBQfdyCi0Zf71LpjrFp1jaawrEris1nK+/DK7PzrFU
igDlRjqEGNbqAUtfF2mpccgijOy+btK5meOnVWjN2NZvs3Gs3lM06FBehZ8GjH6E
ojCHE/jCk3ApxjOFzcrC94ZZXEZCTz/80ywayiHNpPhUluWg8sW5zNQg3TN6xw3q
Pjx97huF9Kz4lCl0aj08+rOPswjBiwakannl+aLkz6TXHOjp6a2f03vn9DKQMuas
kqRZe+gwilQE9ucjkxrA0gmT6h90cO7YN7R6cFaRG4dlkSSgI3IYQ91I4Oj7oiCe
NSZYliuxA8gH5XCzisZwCsnoy4MRKBT22qnam3hoRQzJWEtYPl/j7AVaJgMs8Urh
FDXrPcadaQTZtQGPXtIzGa0AUwG44ib3BR9N9LtrRayks/E26DgonxBsKDd+Ij5C
A4j0DFRtCnZnVzBI8HVytPi2NUYipAk1dmpAXqeqjTw0fJzVrgyDvCBX/eSY0jCH
7oVHyHXb9GCEU1L/3XhHmOFJ3M3Bj98R7Z8nI3ij6mL9aGJS0Qm+jmFT4shLjKly
lO4aw9X09/VYYmvjsRi2mLcNZ814Zqf3V9oplatT+oLwv9hf/vFed0bgKxmAKJhl
Ix5ujvJulCL50eYVoiT0k4soN821+877DKP3hrHLKWRyxfz7vQcg8FwEUAUs7IiQ
xVI3h13d5Oebi0KvRRVpfVZA8DDpwuGp5J+qOgg2exKjRmDSr8+m8Vg0Ad8X25UZ
zCkHEVtQCz1bRKrPZn8aFnHrH+eWsNdMPeqFILPE/LRslk7eaz+EnBmX8vF05QjS
UF7ybEqX43uzy6skSdSR+hrUBy4M3PzFti6p4GT6U/GJWZUjS9BG6H+3QTRiAD0y
mqyH0tP6uo+bcPfcKkvOAGWC3YPN5MqyCbQn33YQmFIdMyx+2Mwjh56n5HGdF3ak
t7XJyETd5C/0w1o9AHqo+NM76SzkbVhAzqSBBynyg7kiJ6MTKWxRRvjSF7+OtCf5
6/M5lBAsGX0uGF3P5SlORB3MaPYxdgDhiBNA7XU1BJUapW7uZApbsyrgsfaRzay8
a4EIM3ix/PyugocFbRIflR4wF9pOVHKWmSct5N08R2u797cPhXQi9+Iwcq+jXBCr
81WVbEtfbZZQSB9wKw9UhgtecgIuTn/KR3/o4MxlhEJ/UjjiU8v1GhOfm1Enfge/
iLBeNpqIlZKFDobHUhxgYstJ0armnS9BJrTkx7xvUp30hlP94kLKLaO6RNnHO3Fs
yVkZ1iT3L+TzvGc/arcJ4zbshKlmh7R/zqfUVhqLTMmCw3Y+YA2kaEYiXuOHZvq/
zfL5cMNK/Clu8/gg37MchB34ppEOgGOTOXPmaohussm/3lEhzuRwWgpqLqlqFXaD
GrP82JMMxte+ufYbALWP88EBb0cyB4yMBJtjBIGzDfQciL/52SDPTHll14QDGvxN
FuV8LPtFGUybwLIr3SZO9c5NR3ZPd3STnQyDpJ/q8JQ0uKymWDgZob/4qzWeEexe
PnCDLYQNc4GnsN2RHBbg+wH+LFUtbevig/rF+UsWLUby0+O2RErZQQ+pnz9D+kG3
UCx4yJPaT6v+9jg5JMwC0xAHCfSD0FvBBQB4aHSPxisjYrrDDvcq+s3T44T7piNW
xk89x4UfInmEHeeXWCGto2UwmREihyYroTYLywlo3ogseyP1uDRkNlta/q9QRD2T
P+dK5brRNTSOOhQI1VKXPlYkyo9uD3Wg+LzuBvCHmioGjPlJvt9Ozr1+FFbog83+
KkSsXtJVs+663tE0hXMpa59oNewzS4mG8AwDPUkrAOhZHq09S0PM+otDq9KP3jKu
Yf0dHliM2K2uYmQH56EhhOI3IqoyUgNubj6avhnECOsmsEC+7LvDVZfoOnZvwKwo
1wIwItB4kWgJil4Zv9KGyRVOcbRLyihk2TUMsuJ/zSMTNsGkAV5iaP8YF+AJH/tq
zRWDberG8eyBRorVjU7XDmzE79jb2NCL0eEOjMLEZm8+4gB9Cjc9wk4SIO5njyrz
O3gCkSjvWUOnB3NQVSlQ+POQaHpx95FBC7mamVy/xRVTw5zMXfUso0eo1gvKFXSE
v9ufGwmlc71ys52ipNYyfK2DQ7AXSG4Buj78g+DVn3hjEzclWtpOds7qd1c7aasC
03fpLvz3D+he40MId+I0ekCJZZ3h1ZDnAzAEvHPYAkraebx6jQpiVoq8VIcOU0l0
dVZwFQW+vE0EgesWxhIEM2miJLa+mVi52yGis7CNoSaAzGnR1kVbeeIx4AXS5zog
DicEqT8AwF8rMdlxLYq1k4BN/sqSo+I3GdRX8PRuLg2g3GeBUsPu/misKsE0Gio7
5aVx48+865oTPSY+edmoHB7iy1GBwPSztHRgmkqIKJGRVH/OTEWFXkGMDq+aNvlb
yC3cJFquwWMJyoWEZ8jMe+bQVTLjBb882aKKKcaLdMlITQKn7K8J4ADX8JI8fSfi
F01mmCFFZVu6R1cY9VLgQ2QzoswiIyby6kUjOxHhbVbjZwsv8nalVzYAX5xAPOSI
xHIUQ/LRV5oC2nDbkCq0yRcgINobT8Zx5aJLkkonv/afjEbMlY0o43cC0Nr6bxCJ
JKWJvFMNT+EDHWUVlt9Z6hGrd88rtL2lmnTvgHEqrrWOpoL24xXnmDxMFg40NHgN
q3s3egUYTmUPIW7F7hev0JeIEWRPZOIRLyges4wR7pvFBfF6a7NLFdHXbr6qP/+O
yJkhqd/mV1oh39Sc226t6VpB5iurnUteT3c76VciMW1SVLgmCRhq27VfxrU0K63v
oBpcBJZ6Nv+HzOV4FhT4nzXEHEa2d09Y7UBGjeXw5nGy+GC7xviWhKbWB3kNIaY+
pOSrepXX7aeWjxiJQFm/392Maylirmq28hIQzdHamCnY+MuZbwNQ9gEp81qs7vKc
Uh/7xTs1eJ8UvcaHcFizCNo3319MxiaVbxMAljTu/W83K10dKQzarxiuNdb3hpxz
PMFuPMRdlL+QCEHQ9kxPIXOZV3wQIbHg/BrVZPzyohOp5+elvEqKcf9bbPJ5ix6b
7ZWCfahZVwcZTNmZjQ0058Q8tX3Jg2N3qNDDlJ98Zayo+E5cusVqQN+XviefH8SZ
ZG/CN+fPOUQnU78OWLz4agzIekIclZKDGMSExi0K3FO89JJSsOQfISi1kU15zENH
wP3FBdyBVZMXxOM/5uiy+1w7/Tlkdjv5WbPXmYtKs6H06qDFfyzCT5K5O7oJyY+n
fa4z8kOs5BWIn106PtsE5/+c3h2Jgkh9ZWoeoY7R0mR8v+ETewsvnl/+WYRcH63S
WCjsrFIRyVTKcw1LSewCSqzvvG/crR8A4ga4e9q1VqqQsR4VBkXZMTGwvwm3sV96
Sxzf+EqAOEjABbz42YbIB8K7TVi869XrVf0oJ0NYIy/uQMQ/VPy57ga9fZYf7pjX
ZC9xI8wTEqbl2VAxJwpMRQHH8z3YJXaibyZzmcN7Vwe1mVBNilj4PzYQymomPz2E
Es7KallphxMJwfAxVbkQU3Q4j+QRqxB6Le04k0k8UAzuHhgCiDTq30uiiFvX+6Bo
tif+B3W+c+andD1iIp11RHtP55jiwNorNPqa/p19BA16F9HYn8Xi0nF1ka3kTTAV
Gm7Aas1m2MUqBXj2+mq6MhQv9/2l/jtA43QT1Ia7pxVHI+I99SY5ZZVFQXD09wk9
B3SgB1TcEsmBwK8e7+EFAx4hRwKBmitR751xNkCqQUKEB3ane2JKIq6TznlMP+wF
fDSz4onfjSxbQM3HB7OV9lS2bJhTQwmneYCH09dZGZn50f6jZeiWggTzFCcFrbTj
snlhXBjLj10k9n7WtkZZqdl57fox7HgwXNJrTOWqy0PddAJtLWAwrGI0RXpe1bfc
KFnHOlQJNNOuMhrFnx++df43y4J8yp+mqdju6QYqnEEe2F3FNkbjZBKpVBvU+9VH
RUUtHqE3whqRcuhke8ki6tqjNk5DJ7k/lN68u+17qgK4AyIwwZ5Gr17aHoCx53hM
Jk4+cnSjNsE6STt56sLSBKwtQ2FrmVXQO0al//FnnI7tiiZfpYjR+A3Eyv2x9tA4
jlQF7duqfLpBe7Q9F2RvvX0/Rk5oRc9i1RqmF7tsvrpfJlAgl9arl20Hw0f2Ses0
KKCBm+Ya45JFSdsfoEaeqVefJaoetAjyqzqUbCGQLNzewtADAfvLffodwxWhqyOE
X9Z+9CmksFMfnxukfSP4dDpKynFrcpmWvFAxgQOZ13ZJVDvvUE+DkJ8cTwHFlTBU
XEJ/RiKb+0gHcuoqsHjlx/sdMVM4Crs90eFaTCZWl0mussaxInwoEU+JllAXSlSf
a/NxF2Kicw4lOkN5TDSxysls5nzJOwGijMiXJZfm+7L6dbO1FI/RRI0Hte+Q+Zld
gJpQkCisRwBw/iQRQEhSRrH/3aWn749t3Chbb+lpUwWE8soyiGO5GxqPGuqmysEs
RqreVKmi1pHs1oIYE0mY5hnuydeIqWP2eKSFXN5UyO02QEQNoBuRWN376Tey6suV
A4RP1zBSWvb8YZRHuc0gfFrX+5V6Dqj2mLfri6SGqMjhKIKy+XIYdoSrQ+GuM0mM
2gA4JozUG93jClqIStayq/z33ae861Qomls52laDyRxxP/hubpx0d4bzP+nPT51n
S7jBGy4c9YocHsvInW3vURT1BqJXXvv9vC4uBq4FNZtku+xR5sCLYFT6JyLq6500
589vvgDqN4/vBaMUmgoljLOMnjwAC4udM5hCErBF1t7nBQ2SqPnp7i7AhxG5YEjs
Rs7/jDbfm+EKH5E3HnIAJseHHontnGxL77G2/AojpqerGGa585wV+Yg+2fjpni1n
eNxPP4Mxef09GN3S3AYzQh63ERi/1g++Idlwa4EMxUxhpY6zVnq0kuZpewSbX3jc
xN6PrX9wm8U8hNof1Oh5aHrekMoisGQ5ZzJSmez0RmEZ/U4zdhpQ4bKACeOmBDYu
QmsxYYUwfJXu2OxOD2HsWRGQvRVVvfy6ozjYiWQdHtjGw5Rc2GiAm5Z2rmvfTpg8
ZVDTPex+Jf3Up86/om1Mg3U4ZoekDIteBCtMXpka97HpKXPg1a8DmWQ/XVDftKr5
Bt/v6NEquhKpJdF2THVCqtdjP2lvuujbK7d6LTFz6o9wnrjFGXZkGdAaFMcxJxZK
Sd77DjcaWKlsDBGtxyTeFYxOTebXJMI0KG+GXscpuf9jVp1r6Y6lWsJqKnqE9AWt
4yBVblVmmmALNHjJwKF++duyVnr8pP6pEo37JCHU+/q860NnGe1e7fM7Vc2a/NEu
xXrmw8IMWBtfOWMvjqYUPBJuiuzF6GuvaSiItmMRC7LgLeBJLXAN7OYiwlBiPC+6
bqx/qFuSP8b9cE4etvVMUp7KB6Dzs1mv7PoFSPV7BaW5bqpx7Nw+nmsP+ww23/Gk
OJTfeCoPRyEOhOxDxaAO+D0FQKcJLhsqjMyziETSyuEXPQZUT9WN2DH0ltlppJUA
2EBKOHbTvtClhDaxfyGtKXtr0eTw22Deo/LrR8yUCE1y+H3juNpNc/Qm+NM1V9WA
Se4CJ5qH7RhZlu3V1Xha2+kkmRiAy7VIuGTgVEnsn0klGuf7QdWAoZcZj/hq+8q1
PCKekkJ3ii7PPNxyzRZDYVIhqcFa1Jo+xhF43Se+HmWbIc7D53KLK5f1th3k5Mwg
VbV89IeIocE5uMH54H1mxwrdTEIImDwSMDrivQR6TiY3JOjEsm0Ue/Rf0C3fXN+d
OgvRxlxRSp9VK93qHSr64p5BPuNEtKw/F0Dz+oO0t6Hbx6Tu5UReHJd7J8e8CipW
/NPN+/BqdSi8lMmncAkbKqCExrq0hhB4Awq4BxFUD5wKPB3pbC0kpxIZWEiVJx9q
kmpT1FJXHYfE8pyB2CG4Ob7hV0AxlmnVd/LAzATDCJpzPeD24kDXqvv1L9T4UBUU
iiTVj5iH/0gOM4jScdeKxB3jlBCAwW0LS2DcSVXFOqdBZLGOy8eF6Iw3cduFV6V7
Ky2E6uYmWPHhhmr1EUTbY4IxDr8NgIahqv3U6MwTArJj3MzgA4oIyHH0tbmhuQHL
ILA2XYyrTYVkHWOC1+97EvcMA0vp2OuUdHM7noRZD+EASrGp9jz3Ulcdjzi1dGuF
h5vQHqGqUw7wkDAC9b+c5LdX5/plFXUxg8NcROp/UF9XRH4EYYEAgzUzYwtd1mom
7Dhco1aepytsHCJRnr3UUcqc8DiKBVapHg+khak6gRhw6K2J+5kKUhtg3KygBGdG
eiWzB7MLfIhWFyZckqsD5shETEDgiIwmKwYoLbsL/iONKzlVQarky+osgVKP0OCD
UWa8E/7X9LcxDjg1oCFkZz3N6J3B7UPv6hqvJItoiKzQAiauSK5ikYLbYNTIBSL1
L1kiJyxXz7df3s7i4ewqORLgt9duTSI0EYTT/CPsz+qurnEpbyV2CXOuus23g7+S
6sB0c/Y1MdeSez8hgZjOYP8SsCftpY+eD2Yu5HFNBmX2bHrcBBKxjxX1EDEugpR+
PtM55DJCHDbJfkb1lVD9l6vLRiBtD5RkeL6wt8fjYcFQoiBekRFNOGV77PX+LNQ8
Ad6l/+8jj346Q0KAd3/7kb2u82ovHIOmkKs1PZbuiHy2voO1bYpcnWGdOLzAiclV
VpVPMRFrOnEusd2YJ+/ePqnC2UPqI+35M8dDF576qM30fSjiRk/VsO82DHfZTP3b
Sve7sOW9owBXnd7vCOJ1GlRn9ReAZHDJPw/onM3J55Yfbm8ikBFAmDnHIphJskfV
yP7GYKUS05AiM84NcyDb6wZbemYpUJi5yswhaHh5KnYbOVFNAGZpApN4+r6ilLkl
d51aBVGrGG5NJUQtYbssB/xYZ4TevnpAbcz06tSFXU/a4Xy0eAdOlIE1ZtHcmLuF
gVElODa+XK7Pdh8AoHgUm6Xar8EA5JsFi0fq2mPgZVW4JaxpsDVMKZRIbD1/dVxX
0t+2qJ0gf3idKhrD2xVbxmrlDGwWWe7jEc+aywf27+cfhlWlitUMxki2g9FgsM+C
FVL93+TKHQfjcQ3a6BhYplvK+BJ+hGBg2F6DgA0m2e0SSVxYNUD5afwKhxZIi0Kb
rtwrK2XfLGNB/7YsEqaF1LjrJubTCeek6fMqKiY5RqZHyPDeylU319bWUm5Rxaga
DQPeRwDX6mF2dUVLsP1oHkk3RjIgQL4XFTTTG8CfcKBFidwQrPwB+HEFu+3K3siR
RN24zqR7PCOUskvRPgxCYn51vhXKL6r2ho39ypRgAksrqKNLF/pZfhfucM5ZQcpP
FeVWNYMBakuP8IPi72P6Awn+1NYrXRCtuNI+ssBMa/xud9/ixPxfke8MGOZvGh3p
CCJWWvlF0SepWuVEVQBPiNjwh98eHGsRjiUf18ngs0HcU872W0cRS5p/sFZsMUIn
mC+PtGo2QG5NSs7tYQHqw7YXCKEosLbRQHLhTTq+QstuOcA3kdinwOFgvzADk0Jl
oiXj5ebwoacS0fwY3BUnCagMC3YmjrrqfE95Jep//B65w2nFSD6t+A+HgMzkbZL5
Qe7xDxPLsBadvz2xt2FcGb+ziTxxytXHRR2qpGgg0rHKomKl9Ll3p9lrKH/E7bvA
SPQtKiFuiCW/AW/mqA2E2pAVz46zawCQPBvzZiIxmuE84JBpXyIIy49CPRchKAf9
71xmlAPLvGeuxEq8M55Rc02jbdU9QtTcFuupJuBDQ/uvDgNotNJCMEHMKYFC5T3W
YK/Eiz2vB4FcwJjwroLULX7wuFjYI8YtRWzVXrxSVaPiRlC8+BDtBXZyd5OMWeet
pCPtRwH9pYiZ40C3GOnznj53PbGoTxA3BOOpZmW7LFrJ7xsVBF9+DPnEhajJxAp0
EEGQcgMIfzueCEu+C3NYfQxi67ftel5tBhAlS4+DM1KbKrpFEhvmFllBxBJKNwhd
Lztx2+V85ay6lqD3NwM8QifNNHa4XNj7EUu3u+xo0jofOq6Q5RzRjjF/xeYndyqh
vyUHLqjV1L4ByY/YG/Nnqtv0YkWBmRHq0ItaWfJDWcsqcFTTaFHSoTdmDjkImNNo
htS7O0p0i3w80Yqb8BH2VxsfmrDgP2W8StX25elIlUNG1CgEInJepndBtS7JMzJT
hWwJdiNINONFceBvuIAYRnx95RCFqzYBewwy5xq3qbZ4i7JtsTxZPFTm7XxV94/l
GP8mNpQ0SVzZEMk20WDVk/0VmjZ1+x1ddtj+FTypZwg9GKBZS1lNTQoKTYpDfSPk
X0n1TAiacs4I0Ifz7g+BB0TRg16you7Qls5LFkH1Rhd9ISvpesV50aIlh8evYOC4
Bc9E2RtnSVHPn5Ny1lGeyeSyhkbbu1xsgrEQXgwZrOLrnowXda5ldvOj8djhl46m
+qEaWT65OvEw+cO15xlkjmmh/oRBINqStA+AFZpxwp1afFmKHqUwJxNynSjTbBfc
ZjnFjqabeIAnIEFb/y/R3XtFP+y38N91Xzl/f9FhAoToVkuiCygFSORdXdUybSzP
Et8CLwmexjwcbdCPNw3ka1vTrtMTHNC6+0pJmP7gyy+DU9okyJPMou1rKpZHX9lc
AXGdPdW6QXABBctW5x+iQtMZqy9xrYfIcd6N92PzoAJu+8q7fmhnAbXb8LrieJes
2sQmggdU+2LPMMYr+FlqzpFr6Q1xl0yqK2eKZDpZaXQYd/RY/KCs20yIvy7NIkHr
8iFoqjkRRvBkvptUkdKOIxDiuXWmbIq1p72fDUhroB7Vn2F4GwGNb9qDv6bZOs1e
/g/IYLaRIZ+ZD4jOvapYiEOSSc+krJE9SNy212xUnhCf6ejSwq8O+jG6U4Eg2lZH
/oZDcb57bzNXjL1cdwiQkhNLSiP+g3eDElnkfTqDTNqXOs2Okd7VUBqJkkNr6lb8
yDjfzv7DgR/Qw60FyFPn/nI0bdpA3tVf9IcmSrc/aISM2ZgLgO1imtb1n0TwERN3
o7CrWzrhW9rBP0S67LksPKranj7hVpJm3aG6qb8VnR+Ja0CwlIEtkChANFh5fb56
7RIdVAJofSfcBzT+ifn7I8SqTMApf4M4oL5NDdyFzYRFcj4qgT5VY77skigeB4uq
wxL4d3XZzXkE+M3pCyrUUrtLi+Upydeol/RU9l5a8Oo5nBdteXee8drcAOIeGDmU
7Qe65rPR/egDyZB+khCJ5CV9uwza5+nMZXyQn8X4YORWQk4VahF+I1hgWra5tEQl
KFkta+ZDxQhSJW+56JXDFLXyTUcRmBEuQG0GdTT395yLWMvE8+iKPBGzcRovZl/Q
vOzmQxMIdfSpjklryyse7iPCLX+XKQM75MQnQRzj5Gs6vixjQznS4KsvfJgeseR7
YdqzlKnxG9TovVIkfR1YwMVtSVysXd/N1tybcQIZPUATSdgv9JdDmTR7wZl0WBSs
y0/OjCw8JUR7pvfDn3GEPIi5OlJ6X0oSjFxBPNeaxH5JFzuerIzI2q6wgZxzMefQ
ZMqf+V1pSRcKzwjT4spjiWbxv5/rc2PMh7jfGBClay07ZzEor48XkIrxUwzOdrHP
JPuleHlnXOZkeT4NDSZ+iqpt5vfXUbFHGP2VXLFf0+gi1r8Gb6VI1+ZtThlCLwgq
VV8gNc0si6qnCCwgAdTr6WzU+qXfKS9G2mRHw5yRgDbIZnUVasFnoiqMbynJUd1b
H+uZw+4VhzOFNvnp7Oh8YALmA4m7VqFKd/4sX/LnJbIIWNO6LQz3Boj+/siEuUjv
GqTg7tRJ1ePBCL2n9m1w2Ynyv7c+EXG3kG031cQ1eQo6RMe9KUYthBDHhWgoJH3H
I3t7khvw/onNHWJbXajbci3DtpijT2Ww4dgr55amniouUlJe+8gqVQZ+3DdLNG/8
+UxUyTQRsY44haddwgvk9hdPwvFWjGnWdXMwCt7tmMlJOfB+S5FuPqA+he690xsD
qE9kWlx8cpUzXDLCalPiDwCFyG9doWg5VMIAGhuJzi9KQVstJKiyihulbsLd0LrZ
8VRY+tQ4fTvwhec0ajyJ1p4rCaT/9CrXOOzAXh4dwrY/eFXlXcTma4RwscMPAjEm
XhNfvJ8LvZLhoJC3MCJT9K8vQo6LRElvv2fWzbRrGJ2s7YDmoCkEGbZfbx9J3g/b
OC2mW9U/YCio0rWKM24IZpfoJZsAZn06LBwq24HUJ0XZ0Fk3NS9TQlrB366SAxi1
fCZZLOEHQAnseT9vW3+ylrGZokT8LJMOPXJUha1IoIRmqEG5+iB+6huQASNKeJgK
4Ba0Xh09oARYMzTmAx4htLUKc6lvFY2MtLT8MljHOZ1swjRZ9WkZ550+CQQHGCKN
TlZjVNzwp+c8SxGl3MD8jix8R9rAqHksymqldHYJyPrwfuZJaf/dBj67kZEd9AWU
ABDmy0M26wHtarq5CLyZYy61BPqmTGoYNXr9qTM05+omp6ETlqG1bMzs0lVm/i3B
/ayhoDNR3Qzw5p4gTzNrkhV1j2dTt6xSe47+veqlwUsHQcxa5gc3FppFok6/srCg
6Ax9siurCQur0UBAOAs2NmygldBYGmoy9wJnxjZp85RJJ+jgcnTQzFLHj99amAzs
eyL5xtUUIWphRmdQKzykspfwLcHAvRr4PyBT7ngdAhmttaSs1ZPTl393ZpGXrQPA
K/ynTPuy/VPsCcAuXLbh8rByU3r1Rp0b87OKKuF+MmcLgSx0ZP0XfcCQsm+Ux+fX
zelZ2ArSCu+2Uy8cUtMAVjAJpVq5XTvTq+VF2vnOMbfHD+boA8V1JDipSoaS39i/
bzYtFFaXb2/luN3J47x+GDc0nD2TW8no/UWjc/zfFrN8vj/x5hBLLw86cuQI6eLS
Q8bd5eG7UJcYVh71CZ/DOZijSV22pw2jEYL/kUF7Hgmrkwq+wUVi2JCZc1j0v28l
G6wyYd+JU0th1uP1CEyaEQaU9sd1zOGazaYg1Xd4lEhv9jfqo2nptnACtqPlGleL
RMwpl/Asp2YDwHbvt3MDfqBn29hC9qiXGp+DrZiwywd725RjC49V+e5fXR3eGMIB
eja14RYtGblgGeaO96ysksV38VYJWaiODkSCipWZAEyHLf5EoukS5FbD5g1v5nC8
OTan6JYmIWP2w8/CBjiyz/55tsfR1KWegzQVSNwQP5BucBEgUkaHIvcmtkRNDjwU
eyNqiKfeT2EpasiF4d6Y1QnZSPoxl73FiWaO9JhFnwUdSllBuOcUX2O2Ceig0D4f
l0c4cBn3pFh7NkpIOhH3Zpjz9DnSnT58t7lme7khXH/g3rSYT7QlJ6xfIwP4Mmph
EQze5uV+Tw38XmHYrMAcZR+5PSFEITORW2DWlqnIDQd0A57G+e8HwtsHtzZqa7d5
qH0y57wrGQW+1d6jKusNpVXezRTKmBNycEzdGsu4G3U1l9Bl3yHt+cfcNL5wABiJ
WVGIX6U+AJ+RfLrP2DxgKFMI79VUMzdL8jq2g0LOdOX/YuLfuJyKm+l4QK0B625H
I74LJh4P9TAgl5k/Dna9gLOZC7RtFHnWqQqjsLliLHvOnv9RP4C9RsKMMjW7dcvK
aODmWwsHmX6qOd7xFze2pFkv4EtaVk3mwSAmDzBoavMX91Mri5fDa90IcYnCKdzO
kQ1dNYJ64EHvwYYjuv9XkPNvuqB6u03hTCfkmoa8N45Z0bC66cnFkcxGi3uxoAHv
frcfwI6SoKKHTno4a81eQw29FmDlJNM5XNBm3EArlAAQIH15C6cOH5UbCW3c47Et
daQffom/DeHt7IAArbWf802xTumJh767QqvhZKK72OsITC7OifJ+Xg/Xnf/ZZ4+n
WE1lEdG7PszP/MPZqe+IEWUffTy96fZerRnqleTROsOl/hCxDFWz3cOgkdwNKYLs
eFvt3sRhbIP4tPuz0izGHycsp7fHXJ21B5iwlLVY5zC+GGn1XrJkVrXJ4Ti/poKf
Lpa5glAcol5xdytikCeL1qtHVt5SCZcffnLgEdRtfceWFLyIjgNzzgim6vFwOsD9
wDa2c/gUUrL6gUjMjCixXmW+8AWLQU8C9uKvFUmOIDPKkNeAAyHh6zaYYKzRFr/p
w3tKfOHsUR6Ye4b0R2XTZWcme1yBlKNyFYO2Nm7eDKevo2TdpYa+0hJhXGlo2lW1
k3V31z6P2kE2O5IFQuijxfADhGHjk9qnmII+smdIOwvTj0VsuygyaSdz4RPAZH3h
c3X6ZCZ2fian3xnZ6YRRpuzpGLE2lIxf0NssM6BD8PBR1AdEMN7OI7HwtYjUsTCC
Xq4yAi4DpSjEY/+4GpkS7ABU6X0Hu7nwiiF41EUoz4Ui1h1kOuaXFZ3IQ0LR8PeX
1X69K+2Ve4HnmwjE71BlPcDzgXcXbUJG01rqKOD017G62aePymK9ejPWR1agY76I
HJKue2ZJr7GmlO5vtYDVx1HfRTT9V/wxaymChFqv2vpviRer+pmJufXDpucyeX/j
DvbiWX1HFbw/ZYEGB8yGXe4baoyXThfWYws//J7qWSteCNNDt0iSEuF4lMjxQS4g
BfwbFFRsXhF9yd5MKX0AJXyUFFsVmr6pNM2rYwPgmVlv0RyZY6f4S1GEiD5aBpQ9
3jfmx7h8LH4Cop0EqATbpg2iNc8P9pHG+Lzwr1HIAWrf9N9TcBUXqTfN6Tr4+apy
qWRhd90RMBQxlhX20kqrqqQxRQMd46eSxT8kbDQgUTf+PBGtKnh2WnAihVYG7aQP
9v5esvTYerTe7u++E+nd6PFHJb2k3eRG68JRa07LxREFY11Av9qVm+tfX9TRVeDL
uiSsIjeOUEOGWs5/kg2y6q/wjb79FANzc+Yk+52lidkjYWEisVsCx2pHQkEbzXkL
8tobnxJay1m5JKi1ykRSUX/avKfqOYYyRMbnRb9S2VVYVT6xuCo7AzsX5Xp0kf9M
teK9lov853OtntLnPCCKcvOYaG0947a97HTb1+QBtYlaTFhXy0V+fAjaqcTqlW+1
pjqWcl4GZTC5l39BJifgJnjz9bMAfUYfz3XLiiivtCVy3c92VJ9Xm3n+F9yqGNMV
T00tfwAE+gS4+5hJgYIN5yfS9x40WzNGcEesTTqrlXyuKGWeiwj1ISwd1l/l44Dt
wxsKAQD+jxZn9Nx4QFcBNWh1a0LoXkI2yWIhoaqhPmtN27DOWTVSLKfzOguIuwD+
46y7b9WeU908VUhRDS596wGHLtSIhutTUxWnAFMTnwvdMj6B1H1ZfwRayb583Zen
L6HXdKScVRSeLD+oOx9XSEI2S/sm0cAx3bIxokUp0WOU+aB2eYPmSBo9IL0fm7QH
3ALoR4nRSmbjwmDR29aAMQ2bvp3CMIXcJ8Kk8IkYnvbOadr4HSm+A4+fsfngKsjc
z5kyedYQimx1zy2sV6++PExf1g+wAu2Mu4XKNKJX5sLnywuPlKv0bZKloUH2kQcn
WLegijVOghTbYMt2TsuZpxqhOgOWhkZiA/kAkjCGbOwFExOH3k+mXrQQypm463UU
lFNgBnO0Pcl+rpeMjltAKZLd74GvYwx3xpJZFfyQS/ciEdZQ5rkG+yPbpOzVVV9c
yjO0o/mNw7iFNKnNoRzRN1dVMZs9STAT8z77y6ju5vYp2/8tvhnMluUmSD8z3GwM
yTMdBjVEeOALxShSS8+74xu9nHsPf+7gXCXCnT7i8fKv3d7hQBRDZdJqykUY7y/X
z8+5d38uHj4UXZ9guFExVcCqVWWRxA/4jj1Ln88i0kyaeAeq3JuLdYsEksWzworC
OuLp/YsdXE+2RpsFngbXPGAA1BFfbtvRjYS7hnclxZE70ySRKMfhoYpRN3xisIMw
nIrNJaUlaWg9C0ZazEbG6/zDDbDYT6DohIYErUd2VV/nTQiqdiXPgCC90EVHqiFl
pNgZRsqrIsxhSO7uHn+lRN+LMXd8cmj8w56OE/PAKaotlPYsCTi0RfwIdenewbN/
SXfeESYIObFNrcCFdLqyp0hO3p+42S68uLQIQg7Vm7DyHvG+yCKC5BwqvOgHNtDH
wJ+8Pkt5HwNF4VXgu+tnO+cmK524Pmg6sePwBj0hV1AeySKHPPdwtIJ64AQow475
7GijIvWpOokjkDXbtbuapS0kkBS0osX/2SdJ76uyu7DFgXTnP6mFI4Y47FmjyD7r
T0J6MQZvkN8upmPtAJYoyfrNoy0JwlLeLoyDlEYezBE/QS6/5aMeyZI5yUFGh+MW
9kSHsxVo9gQ/cTx5WthDfe4otzX4zx3KOEzc5EOInN28A+yZi+tE4A1ZgkvQk2vz
ClHh0ZGGJWVdzZtn5BC19OqmV9KJN8oO81nvsDjqzKYW7jutteVlAKEy/Lp1s/A+
1KsWqBMhXOLt4yr+13GiF+fqj45srJ2XpdsHDXRtZdODdEHuggLisjidlH+6Kbuw
2nlGp3QWJ8phiUq7wpVOS61v6chlucdRh9hzd/4Cn9WxUE4YhM2WEdvPSED1N35K
g4Ad0uIkUx76rkgD70CbAv7sJxbhDdib+gIKqB3IcpqyRhx6ROUBKqyGcTSe/YpZ
4B/88bFs3pK8dMCsLlfNd7QRZ67cnqvfiHLiuhaw0g6nT7iEatGlbPvUXVaCGrOl
0xVmux/3kiDbgpOHReIF3nTV2P2DzkjkDL5bjySRITwMkwHed8h9jie5jfysFE+V
cCK4qjXIDErhJYpGKOpbomwMR4C+Aew/v8LYPuOESUluiHDWNsFLQqBiceDBhVxR
/kUXcxZOpjhYKfeC6V+PeVoZV1V1BDxQerhbV+KNKxYNG/Ijzaz+G7/BgTsP3A1w
kbba44KqGJSPA9G01Pw5Dsyf3PvscSrMbPYaxnfGrngEPWY5eq9Nc9aJrnWVmWfn
90AvWck37WlOpR31M913w5wqcMR5nUEUSZgzUurdTMmeV5g9N20wl86SFA6lh3bJ
ymXU+vrUJl9aukbMngPMoi6cL203c5wL0arQx8Pbym36zMJKezcvHbSA9/AEHM4K
35MI/V+YRJLktdTqhx9UBd2q/CHX5qZTL+ZNkQcpbjUpQ5cqBMYNE0YtDb2Kre2K
/sPes7LnlbGHxRjzcK5DEfFBdWJbqYo86oPyaUktPztCo+hPv8u9yhtRQb4r7JOu
8WOur0dg0Wr1UrTsiW6QdAbE7xsQVnKRamiMRrwp/eYsRFCRz5g+Z5/j/Tkgc635
/Dy2MyZmlj2JnqDdzwy46BXvB5t4pcMJfZo8OmESlvbGgqpcQwVPPJD9//oWUQ8n
ObYLkurkaaBdW3sxlcJd5aYA6MKPsP3eeuf/mImLZPlHDMjzBlYY5+fsh2+lbnfn
CKO+UKgh2US8MTYxqgfaypF9ICZc+3nsYoSLSnVKXqJaNZkIwzaFQNxcQWbRVq6/
+SKZ4Q6EvDWgQhnDwq9uPVzz/p29ejf5R4J56SKOBqaJ7IsbqmCeU/m3nTzHdhJ9
vARDINr0RG4xMB6lLb604o+53L88Z6flKDrvGn15RMhkw6mek3WFbqhIXKn60J9B
+9yqcMPIAPeoty7DHOInkLPIQVSc2nAjVaqZprd5h4z/0wtMu/va4ricoLWEiXGp
csKDUBtIiKTL/h31wlsvt3wMAEbcxQoMc7J7wxKFsf0rAIsp0qpQH+RRki2ZSUrS
Coetonnpp1SlApICuezqs9TLVs034nHfEoWnnMiV96+8rhTY+PVP9vWQ4uFafNOZ
lbI9u/0cu9e/eoJzBapZ/OH3ySp+1/MqAKCluhOkiGA9Yam5Eak+2qVXCdfWNYK3
tc6uL9zjn2BeEF33N1E45PF/qCTEuWjUDwjfpleJ5LIbLlQCWE8mGr5XckmtZ0Ml
28SA1W4n0ezy4WU6CGGOtQHbNAsNTjN5O924e7AFTZB/IWVRFoiNjQUn9JYUByQe
pR+/oGDK08yHXl3HtgZyM5L+WsvIHSxazzj/tCu6v/e8ETkQiXFlM+ld1UgOhWIy
/tsM8GWV8eaeLVAezDiCQ2KIvXcAtZ9WqOSrrLTkMa7hhUp7LOn3/E23C8TDYhrw
ugzzuIsbo1rUXJeqBctQHFHIrls5MDrVaGIV3TtDdjB7wuOjoB2iOgU1P7m1Cdv7
BG9mbsy0cTAn9Sgz3jVkALs13shT9ZUk0HuXcUnIDxrQJzGbdo3crjG0v5dWPpIa
d6Aiql4wKSLhTJj8EQI9mhZ+Ks1Tt5YLnxJiHwgIs9OeRI5EOBgv9tCGv9ds3J9S
JGFkYz6nguOCxWI1bWSfNWMdQ3hedFG+sAcDgKf7N90PWmnF0UX5GqgWlN49tSOM
JXLcBR6hOEzXtqjGKVYgBpWzSkoTw/a5BaVd0zeo5TWi4AvAQB+4nkQlYLv0QMhH
6XTQJwEI7TIZla/jZfflceke1LFKQKe6u1MIy+3BwHp8K91ZtHQmgPPkrKnFiJeY
ASR7iJiyDIpzQxsmZ3l+x7gaZi4rzcmrFgJV64kQHyxVQUgsSQ+hrX2BTt1d4aMN
ZD2RFXPRvVvkbzbzQiT73+EBjZvBf+InL7TCWGqXeI4v2oz7gp5KUvIj4kZ4jDkA
hdPjDWq97ivklWTESS3zGffKYe5Bju17scCqn/6v5vvvjyQp3NErVeLxNZR1rm1K
Zr3tNZPaigqI1k/Et3o0l4vcK73G13BRr4f1AfK+5Az2uBbX4QOpBtwlKvXfmbL1
/eXMcFlc0/e2bIUp3qJWjFKxVei5zysKsjtFKThrvUx1rBQ1P9X8dWrEMXMOtHA+
VzJQLxAVRxD2UmxxlHZK40GqRmBo5LPHgdsdUgsxxylWdb7KfYmO8nQaa57L3s5r
VQveBlRK5xnsMCdfUEc8Fq36oT+Z2QClapTlgVXfnM2nf9xAYqXrtjqJjsSpxujm
UCpOHqveyS2zlNFp3Th2UDDuFS92NKv80Rs4HRQCWcq7tBOfQKYRSMWEjIo6HTaQ
vPArXZi/nyGdxHWbKmMYeIdbnwB3xPh3YE3GUZqG/k1cgiAAVG/tZHI8f1S1KeZU
Vepep5offJ2t/sE/UK99ld05wzxSMttyAa27MyZUx7lU5+5TgKvTDNigAEPYw+RZ
DjliqRrtTKz6q4yN+xV0OOyzl8aQQDchRQ8VJGwqynU5eNxLH0NGdJ7H8Zc6xp2v
NgJqLRxtBq2tydE2pYT3HvCAx+JBr2L0Fv+Klx51LuHogji1v3mli9xwSjm9Lnm+
H1NdhooNBICuXP+uxkezQ5Amhdm31Ih6oauW9SAW9MIRFoAxV8H3AWfCm/Vi9KJG
2s9t+jtmiMxSDxKyZxyY9o5EuqnIE+XTiuVkmp/yir+HRw8DrVbkIOo1uBdeZOrR
Z8C3/iyBxx41ee/BVIySMYtMp1oa3WUS/qGnJB2w98dTyuwjkj0YgDemEkkgvH9y
cKEePT83aYSNFQzECJsqMbJQXEbgTBmGeqye0Ln8+lr7TwDl3mEvxdsxLHNMMGFH
HdngGe1sAGyFUgw3wBvhU8I/HOSMVUWfoGpqcaHVsj09dpdLWASyjCjXkDdhh4A5
+UDxWCZdOMG7jG/LToweH5HSFxJmMfMVyJFcraHC1cDjs9FfVDMAB7Zkz7qXqGie
C660b9m9oVuTgmlU0N+nEgh8OdPjG7qPT5OKK5qIDY+kLUjiHBnl/JGLjQj+5Mrq
P0MfPbf2bRYtEnAqpO24BSzIXBKfQm0u2eQbf+rinlGIuKbkHDSgOW1h8Rrc2kmM
HVQnTK8EuQsk0hlDWXSOgtxMCQoMlfsBBdvJtIQ9con0GGIFfbSQdsDhI1+NiIC8
Itwq+IZoyeaefHX0HIWGKoHG/KsG3rlDK+jKmJpx3GoPNKMC1OkL8FUIxUZFTjo/
mRT9+73eiUvBLiR01AGzn3z1JVa1hhp/2cxSt5g+bEwnFjCcA44/C4PGybkx6mAr
ncTDSubrkvOUHPDQhgc5IjGu7kRj37I9djAXzIiGc6dpfwU73j8Oa6yQiV/q8jeH
hxSXpQDZClQ7RX3+eFEE3HPNEpNNAVeFuS/olUMrDh1hGxEZB+u26ksbtykLcG5E
/BgLI7xEbqQE0+A55/IwCiI63w4xMihq48pYKiVE3RuDKfoXp1jiZHfJtgI9HBfE
GwG7k0b5yjYVGQlyJwuo50Q8WcpVBb0iDeSQHNiQVtlsqp3KbqKKFn0eqb5HnfKn
bIXooxThrawQbElbfj+lXAbxuzErUlYfXA6SMB4alcO38JiG7q7RKA/PhUcHc2aD
t36EapQbP5bP3qowloV5H3rfIgTReCS0DRI9vjtYk+OHw3zHUorWIJJsvxzCC3wC
2xcIScW0UQi0JjDTmxku2Co899TN1gi7Zz6OTh/P4wwAhOi4OKOKVrTibkAW29ls
um7x00vX0Y9LPnw8LYOFiMwgWXK7DlmwDOfBnC58YfB6QwDjIx5t8ssQWfP50cQC
w02gabIduLHMVxD9nbLsoqqhF56ufPjQnP/a5cYiftX6Jm0J8lR2YzxS5NsAKWyh
6uQru0gamSWt+WX/DgdZcCL4q2FYg3oq4afNB997CLYhx6Z2uUr+j13YYNVdsohK
W7efi3LUNZdlG5E4CY3c1LRaSTsM8P9R4XqeDleF3x6X7Rs0ICthQglOPT3vmHJ9
Q/rkoJo07F591VONTSleYKdNe3DAM074Es6Mz8+/0exY8lYUTcgMG/wfQKe6QdbQ
AVnbDznJIDMV0mqm2IS6hwr8s1vQGhQ1dQpo7rvZPmP507DMRB2ttjLvKyPY3Utt
Szyx9pOpWxvHuGjuKDu+rqLYkhBZb3BJBRIZz2EARDmy9SzHDU5X687fg9dsW1Na
kSgG3/5cgaSZswm3MnIZqS8OrmCfQGLaVVmCvVghVtODinchAYr/En0nmqm692wG
Ick+n1t6mSZTZ5J5JLVcTIhCWrreqlM4/1PoOSG8zkXXmBy3XPfEhirAc4xptqME
Chg4EMHrzAS6oSo+fyimGz/xbNfvXmM6UMZh5kkeK9Zqn5iGmhS57zsPG/xOra/p
fjlKMLquOiyAUIq2V0Y6euswQBTZecPKL/HOxzB3BFBw9igH//4245zQ540eX5u4
bscQdP3PLH55exjFEK+L2mznl5A7XdcND0dKhnGO7j5OOO9tjjdZJIT6uS8EPRia
9Rbt3HQI95ozqMacApTd8Pfhm5uS++k4w5oy5Unfo0rWmgnZ0Cq1I/hPJJ8HCaPR
IGViC8QJGBr4cNCQUYy9wYKdZxx77g4WiouJrR4Z1sGp/wzy0WX52OKl4I3MAThY
gK0F/2rUMnB2aEdXLcZnYWI7oX06u6Le2Z9wZLSH+cvjkY1CvZdycFkk4iA5x+Ri
YHD3Wf6Q2co11aGay1wM6EtfuGxTZgFmFU7qpz3aJRAIJaSCFyXfOpwN21zRbI41
oLS+Zf//dMwPKt4STKU4XKzGwnDxMcHIzHdue5WNxhTwNlz+ZBJR9kshslTALza3
5BaRq5T2irDBO09UBVUgqUinAiWzrsuLwc4dWi7tr+acsSguyzvzi0b9quq0Kw/e
GNhLKxBV2XGC9iArMRYxK2R2yuo31DhNrme9K/8Y6+Slb4IThicaTepuCG4JTLg1
4BAbo7YDsU+myloVjK49DKz/kaNDHE5cnOHFXPH1bjnukPygI4i9A3T/osW63NI8
3iholgSQB1iY2pFgKQDRmAVH0nJ4jR6LRivtWmf8ERLyISZO8ICT/6HGzDvC9iRi
Hj6Yto/RwY2iLs7oNeDYZ3Pq6UBaIIE2oWL+fusv+eQrpTNa8EcH/0bJcw2YxAom
OcmCp8r5lIwc/kjs+NJCHkRH0TVwC4Q6S7Iv/ijct5QccwQIv9tByIkLqCypL87E
pVPWTVk9cdrfd4AeUK2Enkkmd650wK57W4tS4O0Bs4Ugmyp48zF5MDJR2Ly2rkY9
xexP0lzU4D/PUcxGTyhYWdQxuIIrW0go9iw0aMU899WcrQYq7ZD4t0E4GvGhn82S
rvPRqLGhCJh3wTyEMUxFaMA7FQ5MssIY2LedJmfRzPn6Qo4lPFhZ0YknnAs0ghZa
FCPhyAJIcoQXf+U3mYfttfRIKnTfiARqrJE+0sK52ZuKYiDKZvYkdBn6J/ct/b37
V43T2OheOlowER62psNiEtbvF+v/sSBL8QiQH+3Zz1Eh73p7MBaULp/RAcRGCix2
AO5fh/7iTL/7QQrKV8V51MKZCeFQIPrh1lSUAz1DpQrqYpktbP1rwEOidhmzALXT
EYmXDNiE22UOyd+WfwX3lmlinKd2ipBCryAB3lE3MLP5AAPPsvmGEO5B+BrtkMQp
dD4y3oPxwpEvyP7szoSZAGjoTCv2mYA572HHGyhJ8nn/vjyY1DHuWyAxPZRGdcmx
hrLAztbDxqP3X6UVIgM8sLCLHPvhEfB7IHS6FIxegUb+I5T1J3q+Rcbj8csb2jMh
P9lNvtoB6jRT7UF9Ye2phRPDVuN/fk5Bmo+lLJF0idN3HKBeZ/QDD7ls+SIiQx9Y
feu6y5mdSZglCor7Sn11DdrgRYt7qo7jfe3mg+fcODvL4gO9XHOr1H8cTu62011v
4v2CpYl22DgFhLVi96dMy1O+/cfzb23PENlgNJPY08e27ortbahrcoLLfVBCq52I
tdl0qijz77g8HsjgVJEvZInOn0gCSK1lwNIN2KxTHownlurgyA6wj8Mo//bAFmMO
3Ep5xKnA175MrqxU/IqcuIeYGYVEyj+dLvyEpmhJRN+15jnYgwgzViNWZc/0p3XE
TcNe/43HmPF9jqLCouHdh1qrVsHvm9Lit7FJjVUXTA2+HqxpyO6lFotJy7Broql4
d7AgW8PUGHypL5TE7Bh0FVrG9yDrr3pluv80uonuzJDhEvbNmh/kyOb7VMvFmoeU
nAt2wmjJTymraJcaZVJAXBhho4B3oreXiVLtB/TpVSs7Z5pr0MslgosAOr+UgbLD
ka9CQFyzBqzZ9LCcFkmCgqSJJLq/NnKw6QB/vnYkzzlir82+v6iephNBD8zVsccZ
Go8yF2xeG5VMMdQ0GLV8AMZWzEObSMPdZsglL+uTJvnh+6ujVw5HHVzEgma+1c+Q
yboHD1jAnMS629Slgly78v1srBlHxzqMGvqHfrf+aCrYkKFNwFeNcF1NoXODcp1Z
p/rwzkc7hv+tywGqsDQZYPcFq2YXN8Cbvg2ufq8bpU+APXEGDHZY4cj+vsLrbJnj
ppTvuNERMu/ldin2J/Ie9AViH/91GZ/1h3LLti62tG3lhQtAdd2PJnINjn0rAcGx
cOVMUdHANvk08tO6XID0f+bslU5UVy5Ml2QMwgv4sPQ48U0uXIKenIaWxxIYIhv9
CRttwNv+QDrcCNxbYdxOzlW/fe2F3JVAWWo15GdQfGjNbeTbYK9XWDYtaEdIsLQ8
155fQgkZG51Zt2Mo5r4KDyl+XzeNQBECsm4g0GdaKyu1sHaUep4cSZ8oIUfLN/3v
As2cLnreKCjMH+MczIZPuPzAeyJUpb043cD7NcPvAtr+VwKUVCEhspyChR/sE+UT
/yaxfbcEp6AqtdhH4umKyZLxk1pH5yu4s+jNrWdKYPlthFkNPtQ2FY3u9R8LGHNz
h7oeJXJaZDnO0NnEFInDTnsE1LhJgT6MRFPR7DZC+XHQUTBGSSwfb7nn8IQprWbX
0KBFQiY3AD31uD5KD6zot2mZyVEyGUXmnr9go8i7CEVCSJCRz6VwH2a8S5o/nloq
4Iu9ifmW2nKCEDTFCcPqGrKNBagWyp+mqC18z3gTQi6TrD9eElUaYvZhO4esfikx
Bz3zJLPspWVgVAnMGVx5XAEosuqbRgPr9dhbQutRMniQcBaXXlmV9rMGGMBnuBkU
nsB+hJpGGNNb7xqS7vN/Q5fd39zcZpu8ECLzKJDOWXhkf9ya/vkbFuhnCxWHBVVp
FGLYpK4ZPuokGpsVqSAzKyhjqFFu5Xl6FtC5NdUoSfBpQ77H0tERiYnvSphESuD/
U6N/3R4cRmc4B50Vd7Q6Ge+kSNDawkMdE42hEIZ/KrqlISimoAfFf+nnTt+IHbSg
kb+HhkKc7mYAiUpgCwoP4p8ng683vWqUUUiewY/53KL/shujs2sPzhyG3Z5kkKJW
NaftQWUFqkcti1e873kk7RaIiqbXvmriFQkTmzq//kt/jjMPLEczMspukhWRqIrH
8Gzjy+fKuPd8P1gDPyO67oGmMVjKL1fJOjcfcXcfsDtfvUciec+hsfXPoce7b8Qj
vVn+ziYWo2cWVGdLGbdDrvnb0Ofk81X/QoDffzYBVia/PTQy7E4mVi9QfgOymQBy
qnlGxrVruDUb44qdwZXt5Mmpb94C0memwikBbs2o5wPUnhIFNzP/BnuSWFnocKuG
sZu/QHQR60eGr2IRw3s4z6g6ugWXoi/cX5Yvoiei/XmWcrwzZ9eYtj7U7QSSmMpi
mjhtZsMdri6iJC0unsIEZ7zaLdCWNOeD5bZjV+mxzIRMukelqdHyV6DOUkm1KCux
Sokdrjxwcn/lNJzMhrX/f1BmXUNzHIeI/iTVO6ccoD6zRomWc9cs03m1T93f5agm
rurHJZNKiiXFoWTKzt8Kh3QtFJB5OMQiCJ78bcgsp07lqLYJhTKx/Qua85NYfQZi
XtsTQ/SFObE1cJOAOu1M/8Sb5wrWsd5VsCKApZJUa3BfUTowuDznab90bJYllmdb
kK07qGSJJSiyFjb8r9hZbxe38hz2JCSfw9+2LbPDvKolh+WAvL0WSeWJ1cciXrng
OcyNVPYVHx1KWh2MQBWajQbtvcR0+lt0WzMwlbntw293G6QG0iaJBpu3IgPjZERB
dVwn1M0y3hiz0tmZF4AhTT0g9PkJeJdWdl811OuHzOBM32NfJCMD+3kcQ6HVG7tJ
oHMUqVDLlzHVAs0lTmqk1XrEUnGtgm3i2fR+aHlAahcuvK0jSBx6bngeFQyENdQe
os4ndEZ1TJ60bRq4H/HrwgGuBN+a02lZEi0ALwLcHsq3fuOxYvb4oKzaCB1pq4es
wDt3pcDeOyLRO6K8E6mHzaj6Z9qdQIWRAcN2JiHGbP+zHGo66fyRCILEKg6luaNO
J0jIfvNBFSWu72u/xzrycWBeRU+fTWfaewmPVm70dE+K9JLcBxhYw2VVnP9cSy5F
JVuT72te17y6/47C3dyZMXorAT+IBntXDDKptHzWfY96DNdfwMNLvdcca5MM49t/
fdSyRGrh//ksP1tuie040b22JHi3SgiIRZxOw2z1WoCP/Co8s+/dt5lsoT33NXuy
xTnQafisiyxfER46DRSce8UhKYpfX+rinymxsOyc2Ew/2D9g6YoSjeIqvi/QwD5A
Dm1jDBwuvPx2M33RdLulWbq/Gx2OMLP3USRgemQE3ntgiftc/6UckZqF6h4r8mzA
na0v8tG8RCeLTY0MSS+UmRjJBwk19UFxYVTYYMfGlmsAJ6nwbmUYzGpcC+SudgyB
FWN3xneP+P86lqK0J3qDZzipil3YHBFiCjORzEG4yPwXXHFSuMSRV7AOwl2YGsJn
zuKOrLT4h8xsuWXTHUgjdV7oh1a5rBQrHhHxgVELK78qbzmYg55VKgtppRNq9n//
nSHNXcOii9VuMCrwbK+xGmCFqcqMSztFMKJq28BKgzmxMxaDwix6RI1TT68zEgcV
E0daYlQd2Llj4gN5QRYFuVSqig9mHyXRj2q6AzP2prR4HzQNyHJ+MlecblU7eYdr
ToIFdTq2+8weN9lXGWc38585tIbFQfQ82Dge6f061RbCl7LUwEXPGJXY3ia6QwTj
6jJe+5pztS9aIP+qExcNbSfWF+rOGGht/zxvETMwXox1MZjJgl24SjQjWHvSfVNi
PPaj2JHmRw69rYjBl88JIOi0CJFuIEEA4aclCww7L4AKCO4YJTrZYcc31DUA1I4Z
7ZoJWaH70AE4vvYjsAeJJSZn5+morOvQAhWzgZzrmVUNBYMfn3f8mZNnqr8ochpf
bHFM7R16hGOBA9HMBiUayyhZ8TWIQu+4KrR8ewynO2sIvaBs0+/90sCmoEPyFGz8
T40o04uge5rTmpjLWiRtSaFqDlHVz5+RKwoU+DE8Z3FQo3A+WQxBc2sYB8EqeygS
ay15zTxBzq/NDMizvWM56Xx946Y/33UE2W+zE7VlewVZzdl7yD+0XOZ/CQ2TMgAe
u5FGf5q65hOFKOV3s+gGNN2xXUnTLxZk159X0IHmgBhdqnI1dO7iwUQL5nCZLqO8
gVS6o2CrHaiJr8o3NraGzWMFl162LaNcMFB+OJJr5Mwo624cc6H/RgFOmBc880Vd
RG/Q5YQ3Li4eZvwAbJKKN4VyNVGijgeNkyw7GASYM8X1HU9dHIofIYyhR3Y3tEmV
qV4GBPv5J8H1PIofCawNg2vEDRonIRHvIXNMBbx1EH0cAp3X1KuwHB3VrjtmjY6B
iNMw9YpeRhS8Zmzilmlep4Mabb8v6aH0cpdEEgVMIzjVqB8HIdfy6T1LA+zyJ1p7
JNEMIO+tNw8iovRAvtFtvZxSOo/uxV6igNv+ZGSYxlt9NK/AcPFyxUgUQXbEx+4K
EDlwciQOpLaWuHpPRuF/XCKPKNZME1BjYajkJN5DJMHt5iOMb8gtP6pII21O7O1D
sxePEezs4GVqc+rzw8a8g7sunDRUplR4U2oYf7PeTD85hLSMqhQNAwt664mnygCI
qVzknEj6uyjXwCEbo8yhIRISV1sb1hHcKhzNHW7qPEQQvqVNFZbVFolxkB12Ee3d
A2pAJ9G7vz3LSl7wRJ51OlVfdfMKTNrn8e7rB1RWEwGyTb7uu4cmooWjjV6WRFHi
S33mCK0CHudDNn17sauouKHOeeqJ68FsrwCBi/F6hISDGb192ttiqRlZDAX39N3V
ng8cCgoi616P+ieoDPcQyLcPWy9k3edKKyRMhQ/v9qJ5iv1OzhIZt56YBRkzwVOX
RhPueCsHzwU7gIUdTeNQXe0RA2xitOiQcGv9KFUCehSXCZIeH0ISic4/I8p3OlVZ
LRe+TLi1cu2gNibb6PfDDg2GXxxUxUoCu9DFZQJAbPWUlL0KIT+PQ2Oay283HqyZ
WSo+uv0va5I/gWqnfHjQl9xlQk9+IUi2wPxtZW0aiBW8yi547zCLf3DL4DB1x0ep
4Y8dS9jPmSUnrPkGL3yEZz8ZwFq+5uy9Qjcbj9OuXH3gNCUsithG6OCseEQ5Y+CS
u9qdgZ0s7ntGl2Jm9N/YdVFVO5sZwNpzF3K+4X5FTpGf5LWlOKuRpYlB+eTM77rK
VFYefVuUCMYyVKCHSHlnLlLMs6FoKOUPkly/PnxAciDZ9gXhvw9//iYixbNGVoHZ
eXPAE/K4v6SlTHZFFpHyyC7LjmT3+lOxGvsPuq6cey0C408KsWG37fn7bgrnV4LW
SpUBnCeRpm/E9XX6xCDXm0FStBhUiw3M3M+fMlLNCxdZx8PfcdJeFQwylc+DKMgH
cRbUiKPZ+3TqqQhiXUn1DpcaQ8OzpZRY4t1yE1oJSUZc+KNmibK7d4e+S96yKkZT
S62X2gHYrK8ubRYejTxIZd4j031A0m0eQZ4kuLzcxdPtfkketgxPU4LWaKfkW7TW
6YPHW42DA+/VEHPMh2z+O28O/RGgosnJ8T2PD+IfsFG4UfJFQB+8WcH2AtmZ/lOa
22MW+RCBZNif14rqqwx3s2DlGLtkZWaoTTGoU0f+H2Y8GXZ4THfc0gixoD0eMhuP
9No9thrhpE9Pggm/qe5akUl/Eun+Tg3gWuGUEVZcaYD2Xtc5srS0vRwlk/a0Lj/0
XQOz+DQ2G3nEyFehRfIZ1MGpBcb+oXatzpGzHTV0w2B1nArZ//qMnSvLzduzqK/W
/cpb8r/p76n9vC7q7aubZE2xhfJ132BpVeb/a3oLrh0I3g4N4hPcwBQTVlvYKydV
m+QldXyUfuXLUd/fSTfKl5jXPC2D9HulDJLdXSfR8TfNCIQKVWLRanoALiSeHUK4
GDx+cJf8AdO0eg/NxoQyABRKvZs+iu3dhGNwEa0r943yfAChJHl4/rdZH+i2iPVf
Y/NguUETlwxDFso0fRWO+CjTNGXLLQnL5xpUu9lAeXyzQy/GSIJlu9/Gyrqfuiqb
CCjFLNofsW9aqj4kHeavvz4CzB+TFbTksyqSzGhdT8jURlF2V9HAR+KmR69ccG9m
mIlH+SjvbUW+4NlJTx1DMqQcFWYyhTy6ysrD80hpSrrA65OjoLkxD+LI3LWS2Kjg
R+QpQAKWTju6uHsywovBB6GV1+pFrsLmufad52kj+NSQNiTMoMcpykxJgDSAr0WL
joX1kOz8JtPg3huB2UMsCTXqlICL0McKOtFWvy+gIY2QebGq9kOIJhh+EF6MYHyY
JmF/cwx0S/KcWhNDhdPgycB5CKAM8RWey8wyU7DZMGc2Jhl3fmrP6VIUKCa9KA9O
mmyv8TjHPhdFgEFo7VZ+o+VbXujmOxK2wm/n3Z+InnyEGd0c8VAdNJ2lKz0TMB7n
HgbKMLFsukX8azhua2xpN6ivu38hOJG0P0KBDJbVTj6wzHkH7PpWjh1z5LNOTsm9
6cy6nr2CW2zqUuuWbZnaS/XV3mbc152dqYtnU7qkrmQIFODKdrDwHJRFVX7iGlYV
7+/lMU177IO6aZebucUVXTwDvMMladrvRr7+3Ef05bWLTptpSLEdProa+U6EODhd
OD8UkAilkmDV3sVqqtqCKs5F33BtMCALpwhQ5ju+NMyGlj2JGkP6adCy8vHR2rH3
ggdHaFUl4WqfEtziMXvN4FPjW5hQ5nCHcRlPjTVLo4ZlDTNRzGf2d7ZzmXwOTzjN
07bhUeBzJGO/E+OaLp9B7DFvXl3eAHTBT5ZaxJV1369fpNtxkPDZsEwvvtRBK8W1
7LtrUKcyvSMYKETSFcO0RPiBx0Q1UPJQCXCKKGuQQlWuWgN+7SGPvzRmCGGnoM+B
7wpTyVdcwO5hEsBONkDR4qhrp7pJ/zibN655iEXoRH9jAG/v/hRxBJlRod6iDIgX
W/9Md4GPbRFk42a2uGrIqk10okJikUNyrWa8tTLp3PNypAeizJpwK10ujOeQqOGI
PzHfx/IdVZZdyfO4a58XqsqE/eA3hAK131ZIVg3w0nzfFG+EcIbold8jINamgkKI
h5e5Cii/T5dHTFTvFAaTBjSGA76n+2/8upI9P/rHN4Ifz93wyE+dgtstxixJAPJ6
3x0o/jtglarOyzm08g+mq96zjgIKoiMfJKpvgmxf7vGmLfYf787TBHGF5xV2eF/e
7fsNhZ/JLX6DnV8LG5e1JDTelHGmDhUdV3y2N5eUK46EewBQbaHCQqD/TV1QgYD5
wKxNyE6YJw8RObfcm4G8dkacGIeyfbI/Xiethc+X4m+/fsTnfZC0HOQiD3Wc5fr/
tNSt0isDhjcaunJ8s4lYFeBW1N0Mka8YdE84ckYWNOD0uIf3XkaV9prKKM+5KE/d
ZEJb94P+avegzZ63+bk+wb725BCiksfCrgyOGVLR4CUsdbN+lXy0xSJfO5Hnlsfj
dygbwLQ9/xWwfxOefFmSIjJifL+q9cXPwP3/jJs5/oTOSNy+UNCKMUVT4kMTRAul
5j7a6FWLy1W25e1ZGMo5A/DXpjbFukaxTjAaQzBmZaYElEhOX9x3D/fpZDG/QrZj
hMMa9tK4ngxDmUkirQx+mV39qMb2MDbavaZqrc3NxDjeug16nJHnQOLgX+HLDrZK
GVX8wwPz/TZQ6MadP9tKuOqI76m5sbvdylGtzUQCWuj6OU9bsvxIeg+A1+FKCC0j
tEGNXReH0mDRRez3yNoYPM2i6vzcuKFN1Dntdl8owCrYyM0nfOw7j9WbW73Sin8L
L/f7+2dQxPl0jSAJDe8IBnW+jgCMgKe5OtlH6yZp+k3i8420H4oqYqcz/KEkSPPW
lj9vGhoNtW0e2mZdNGhWbrvCczVoYkwo9vHPUj/jxdjKyQSgsYv5nEO2zg7h9eeT
XuHP23HYrcsZW4RhOAQpHIXnPJgLLr8qDANc7OWecCB+zH3Ogf7929mTUWj0VrXd
h/NiGh5Gy2p/H309oAcgVono0dHiXA4hGl1J0BKd3q00AVCnY2g9mS4fPBdJY1wt
aI8wCo8AfIihMRWT0+86lj42h0ngE47QpkjQ2/fIN/BagVDlo65WxCBja9YuOxNq
w3MG3G4q0+K8Zdu8dBxW8CiXKsWJRjTNyXPu9X/wipVRWi+ki+RACfXDx2pXRFVY
4vm6RYdqMAN2wlqum9Oo0nluEWbAK0AXb2fdGLfXc0f9/QExX9jUIePXoK6JcJ9m
Qkqgyzfo/yJi8IACWMUD6eRHmi7lLhFq+zsCRXR1e3RCFCFPyX7bgKY7jK3i4UWN
RwQxNBoNlM0SFyWrUC3Z2T3fs06wMXWKvcIpIJm0mgiC87eqr6ePTPDoeSmX3u4/
bEiry1DTjUeiTXxdxj5zQ6KzmwLO905Vyhb2CjlpXSjo6K0O0I2dl9KH4sZUvVoK
9wjK5LZU7Hux3Z2RmGG/Bb60dQkuz8vZq0BS9NSNlrHT1c8Ay5UoIB/olt3NZN2r
x1wrLdYjdHY7HGfNZ0BHF/qrMJjEQfU0LP3eKy6KPrLW8WdvPcItYfcsIyU0nJUS
hOolG1m2L8bkJboUyFg/MTZjqsoLOa9XtWBPsSt3N9GB+/TRzJYC5hfII9QAXMQx
jH5nszBuBCS1WFc+nZrU4miNaPpk1C7ovxf4ophTOZXpAnyMBJrEEOJIMVuS+rB8
JTGr/k6jYxW28Au/SUlpBxU51LZj1zibeb3WXRTMj5evOx/xz5hw5/tdgZdG+JTj
5zPik1IdcKNbCz2Xa52wQX8PLI/2eZKT60piiowP1qY3+3soAtmCUjlcf508z6Op
MGclaI/KSXbQSg+aMSt/WZcI7TTfHksjjXaelIOV/GRuBjsv/2BtNYdkqklQfKI/
WvhEPUbdQxegjqNMzuyKIYRfjEPQ+ruG37hQhZQKkkZiXsNiNldVGmeKx3P/dbPM
Y0gt5C4JKgF99Rw1prJMi2CmAQ0ZbwyDKh5llIwYBmVzfepsT1lVTJdFdgN8m+YD
oM8clVv4+i/FghNNOgHrw4RLJajA2FLdpM4JwUbwZkb5Blco+L722DkuNk7nxdCS
sPabXsAIz+0dD9aeXR/elUqTY5+sjE28f0XH6BZquHuuQEgdOD2oQotj+XBAfsy5
MF2TeP7E6RmwHDxt5qyqKfwVp+vYN2U6fwag+721mOUvLgrHpHFa7oZ/maHSYBK8
ZIsvfsfQtvGG5/MALZ+jiaAj1nbUMt9dlawGjuU6I3E2KAZiKz4al7mowyv6Fivs
woQvJ65BzLvDfgAQHYwu8tb4ZGYp6XPon3xVMxPDBTfVZ72kQnZG08CkeMlyaA/0
m6FnvMKswUhwQZ3zGW/3xoOiKXvYXAHANUGyC+laVktfnzRB0yqna9E6iAb44h/S
opaNOM7MHokfRh8/A8y1T7X3VrcJYIPco6BLAooQW/xiIAAZh9bnmEqdhKR98ANB
Nh0RjVe//xU2hmxgD879c3R4aZFkagzCBbiWzZqFwoF2Lf6GOI4J0s5/ufASFYjt
jsJNJiTzF3GS1QTlsKXTnM2pXy01muy1z8ZbvBj8u9VFxkbGgjiVXukRePe9ipUr
wD8Cq1zFwqPvDkz119ucB5nun75775vBSWahzKoS/NhsVPbtgly+wSF+OlrNZb96
3HZgDNRuv2QpuekIoyEPdWHEs2Q+fVodjM0RbLd8Y6Rd9NdwRin8H/hE+SxbY9WX
agIzZXkMb83zqEcMNbUwK9AWscDAAcNZMYng2wBVmNJRFL0IuM7rlAWHtLgpp5kz
papgjBil3sRX9sDBC7peYKKXh62sdAUyzDrCpepexJizaskDhIyeE8zV5igZm/5e
Z9gOp53XXDmdyB57PJSLTqVfZvwFy8JVCqhGDgghNfiEr5zBIolQQUc+UX8yUwJi
KjvOVbDVjL10xRoKgh1T5aZXz3hyUlGaQXFkfgFIWC+jmVjzt6RNyVIqnEJyuLay
TCHEobkpUDjJBGFmrCsuw41aRZxEXdaYr41PHhlDJVfr+J6COFeqxX6z7YWoOtxc
apTE+5UF/fJXjaP6rPudMrGG9/aBaPhVf/VzZTdTK8djS/TLfpKaLDrb6XjD1k/4
oBC8ucxDiMK4eyZWsnUXkGKlntQUtWoZgsmlD1WWuJqOpv8DWaUbsXDpu2fIpEud
XGFxDTzG6+e3zJ4dFYqhsbRxNRX1CJgQxuSOFMNcIN6wXC6QjtK8OZo5tkVCt+h6
JcF8wFGGle4hyYef23dkECwFT4kBaKozfXeDlj1P6trakqD3JpH335raNF0nmv3/
guCTy248+YeCIsXOvCaAN16hP6iVtT27m69aQTlglqQbcxeSPCPaKZdghiWnJrZ3
pTdQTFphZcr/kDi+QiZYDQrDYzfRqP1hCPCqUv8VQcmFubi0SwaOFSWLIg0JeKn2
Aa2SP3at7gdzYR+oAr0CpzrH8akQzc88cCVBxNciAjuL302yIiFVy7MX3aHejtfE
R+cyaF28nz/3e6N3W8+w28OX0oW6Fjo6PY2sQAbYTvUFtk9q9dEuUnHZWmUDQmKJ
In7zeAz0o0HeMtNESwSomwQsneutrNZ1rUHyO6/FhCza805Cb2UYSlTV8FDW0HjH
DrbfB/jU5IiNwwod/IlTt67vIRRbX6qJZojrI2RXEEnjYsQDh1sAJvP/zYkSX3go
RregypLE0nv0EDfPgJBkgwhrSjcYJANvDnRwEkgR4xcEjGtTph+GIOWtN8NYTsHx
vATkDGqajzeFsvgEOA5q4PoiD1pROvqE9EbgkMVJ6ECnb/tCGYOh3CUN7WhzUC+X
9D9M4pfS2nuukdQ9Gjb/+dyhx5XH3vVf+vtfaHERECNQK0Z1mlLV7mbJB2LjIJl6
osdgwlGEfwRJZlnA7pNW7NZ+kBBuiVKFLcWvbRj764hymXzdNLzQf8N21hFYAd6p
m1ngdptaI+wYluC6Sv5SynQqJLMabJzFpG4MPfLethIopw1K+vVYg1TDRNRy+b+X
MHHSyrp7wr8tR/MrAZsw2rSAVIB1S3SVgvv5O8Xmj95kRu2Y5+DpcPakbCbL0MfK
028IOAhFSBaZWOmJkLwMh0jhsT9FPksTZqZyyTJTmZVDuS8y6AOBgZQaa6pnOB3q
TFBNBaenunH0qlswHPAZH8u7BzrT6cdKHTGQA2v2wsPVr+wG4t1J4PtsMWwApDQC
g4UVks/LWo47I9Bk+n3LR4VvojzY8vCN0nmAWw+zT5lvmhd6uSzqu6zZPOPW9VR7
sSLLy2ARfpk3+zpb1LzBqnE7KNcy/reK6L8St2h9JJ1Xzw/19Kx+dus4cEhSsC19
8OHmfPCnSfev18m7GtrbbQVBPUaJOiQjx8dTJqKdx1aD9Yk+KhXVnKTfei7/YAMS
7TXyc+hppv3wSaIKl3szYNQRbR9pYu7Pcm6ABRL15jyrDTcHDrS7MtgzLhv7T9RC
4KyCRLYgD4xEA8sbBJIjknCXwDyO1xxPWAC62WHMZwSeGhz/8RdYyEiM8J/syGhc
Ow+k7CEMsU3/rgw+Hjym4HpIkXIAQ1Y8JCKWllNzXLNYkDnkZ0yoJYcY/rdwX57r
qOcChpIW1Xry1Lz90yZ3nqSsYCNbmhE0Y8kH2zU9+T851D2Yjx5x0JTPtlBkjkQ1
1g8sOpMa1zHOhS4bviTuk+LKVK46HCh2Poy2Xf5V5QjOXP/TXRcA49T939FjSHo0
UZI0iwRAU1IsyLC6m1CUp1oZSIvbWUebIGJaYCFqC+PzkbfA8N8IynJ9gXY0k4u5
jnL6l85OO52yxQqE1Ou/6Z74++AOEWsz5GNtK5spHZrMPP2ZClVswEEUvIF1yYB7
wIA2NcKRfBC+C07Ft/BlgOeZlW2A5aBIz0O61ZbRvD/ckDW62C/qkhuSVTZhVR2R
1rU2qhjvEocb2CTPexqaFsXIGOMInW9OD6PdUVpib7+kbCu3/ixnzd3QSWZ83AEo
7ea3J6gKLx/x46aS/vap97iSF6BCj0d6/SI32qhjPTQzmwOmVM20LwABPj1EWyy/
t0XzWWJqxuxWUHBRHgAdRyh7luDTFZ/svygk3s9UlEFNGQf0XpUf3XQFefYV+02n
YLoihRc195qw5VwekdZQS/dkf5BaMMPR1ir/ga3gBUGLg7fziJFRYeRSjNIGr0Dd
Z8U2avb3F0nLo/zbskTZJmtBWQpj3y06ofU4asdP6IqO7Dy431yvATDDd8e6t2gm
3DPa/7hPd5iE55wbkGvQtR7JoZy242k750mGSYFAWsq6i2hZtcml3+TxNr3AS4P8
8ST7JhK+OMx9AEr1Ja0KnHdvJsCEwTm5zof3Rn6fBijJmq3JodtlNxm3M+NEqa/8
V6oH7xDhf1P8vgf8cpiA62xvb8NrP+g1aW6mR2eCPj6uqIXMalokqVenpGQ7C9zx
mi/N2z7hw/Iqa9Rr4pyWILLIz/jfM4y5H45mO6VjkJK+kg98qkxk/zgSpNqhP+ui
Ov2qn/npwkGYsgL9hgV5vlmTI6rRsyLhFDErRpBmsB8HUx9W9iNTPsAfIiuMI8NM
YsYp2dQeihmsPg6Wk6u5ggs+0ddOGhWE52ET/a5B0JN7SrzDksneLVp7Xuaa0uts
cTQlYTeLlYdE2dZKUTG1KFRm34//WqtUtEti5QvJS/8P1os8J75GhyQW1BkEEPKm
tBC3sSUtNcaCpqVDcbctmv07sBOtKmUlEqN2dSV0zBptbP4cyzzefJHoKC5zg44l
VjXusXVjAF0wN9OCs5C55q9Z2QLJIy4CbsDWWcXfOzpBl5x6+hB4CzJbbkhVaxsU
NjHCOVwFZT+w8D0FHbbhQqtdtv1yIP6ad7v3A1+0akXBRAgmjavBshfNuIdxI3cZ
3qBaWCrg/FWZvnraei2SMKTMWDRLEGhhAJ/2Qg6D80wXjM8NaWVV35bLVrc+IBOw
D8qsZpb9Ja6YpFUpP3wqJELmKnYyxZda8yN8oo0na2eDRHLOnYlU10xzyAuDYNIX
Du3K/YtOZpl2GBmNbLUohfX9w5Gb1ZsZ1yZupY5mV1z5PV5ccX4WqYW0bYUWifnV
DKgeYy7TYJz1QTv9qXeeGdHyTxzJOhDvtIW0o8wLMcAwd4yhRxcv46Bt24ULH8Hi
rMZI+T37Q3GdFfryqDqh6xDBZhwfvfV7qivmLjutFeJa8alJJC/qQSoJl8XDrkAt
6aLpcQBIo83N/tQYqL8OaoMs9fytkhfosvq4ZGeH2YNaZ68OOBG+RCvkT7D++dbx
X5JASQo18r5QsWz15gP4eu/1BpZos25KjtZxWACYXJkXQ5ypZVn+Jf/WVTxEThTP
Lo5fCXPFAAZcQY6J06kUHvTd24Owc6cZcR99H/dlhXUefx6bKMF6pRokZ9riLrp1
WafgNo/eHK9khn42pB10d/dkRREI24AUNxwfv3Ef8R+a35/HdWhkGRQ5CmRccWEp
RilVcylf4Tk9t/S5zIFaWbAeGMZ6x4vjbxFBRhHA0h5KG2BriAl/HuOfexJMT3IS
c3SPPcc2xNqV3GqN1Q2u6Efc3TlTY7RmIXuxaUj/lSgmGz4H4kj/4786wpFMUOcM
UoTaVT6DXgCkYhwjpXoOO/E2q3Fydq9zx6a263Ph11iw9PcYhM4qeHTuPCVfQY5D
oYU6otVh+V/FjCcAwpFkZGXO8+MSKy1HRxHphyD0GTUzAMcVBrZ9tu8oTl/seYQl
Bwi9AYrE7aQQoKxyP6trxQq+xiNAOWqHs6ZCt9X3QqVMaG95sJWZqWgbCDzLjmsM
ra9xQa1bpF7aur+NTshYhie0nUodoqLzw4v1aCU+0ONwjPO+0QPb0qPUx7yQT+fL
gB3psPgnbbKFv3AewRqmvTahrKmSilX9L/r86z7Fb0p3UqY5pi60gsz/pbQH8CbW
3F9pCz4E5kwJIF2NJTxWFAMRp4wWAES0JPF9+iqB5r8hXHBGSDgmKvp4NY+Ocm4P
ar16wQG2+44pnDN/xAWMXA+Alt0O7/vqJt/oJK/ReSGw7HpvhYs9ibnzZlYY0Y9R
tb3tu+D8RdvZLNJpDcVbTtiGYTrLDkq70MvFhBX4yINfx4BIR/wDGOPnscZOE57M
NZ0rJjWAPU3p92MlBeSZEOOjq6Zg682N3N95oS2olubHRm/vTFlNvmFDmaRiHOK7
a4bJBZHVIittv1HPZ8FYIRBF9bLUOdc8MYGOdyAAv+WRP4yh+ZLi/S6AF4Ma6o8B
5YUjO+bL3EoC8L9cwG7W3NJmPPadlgswVRtwnd9UdiILK7rAxSj5pQMxkOv/wFya
Hy9lDHMeUEhdBBfxvhHOLVbKAJ8XKGdZoeziLiQGy/IhAuuYcdw3t1TTyDvaQ5v9
2rD8h5WFp3pVsX8AKDbwel0YkrJWdN+eRW8OfoQV5bkhk/0/cpFLaFTkG9+iZfqW
axlo/Rmkk5kfG4Df0zka4fLlxsEdBZnj6DNqrk1NavZTGjxqqM/yjz7QsCuS2cZY
dct6tXunYsMAIupdElZv9eSde2tGJ6C2JSp2UkHeNFDxoNx6BnwDwMkqkd/+lQY1
g4HMvvpjVum49Z1xYNsF701xlFCHriwyz+0nXTxJ1hybMYLcCeQ7HVp4VG7DCya/
YDL380s7CVcL5ozQtWx+itKqTvdv89H/di6I9h+H3XGTXMVr8/97WtqCwxqryuP3
ZJN5tXaSaKLU3lcrWz6/thcJx79VSafquPfN7iMgJhLrjeSaNVrJsr2nculeU7+e
I/N99X3S/IjqQtTGck6UcKZUhH7XaxOVFCt2AdJ3EsrWkZNLBpyP+L102+vX+9/D
7CosUnXZd0sT5FaX0qO8JJOo2FfTQL/yndnMkceHNjRjiQtBSyYsWCf0pA7YRvpi
fLI8+cxl5gsG1/ew8eztKSruMwE2iJnEf27u8ugKRM3/ifnCxVyQmCwDmsggvGYX
0tfPj+1Gfwr0mDgV5kztGFRaVUAW3x+ITn7u7N6gOg4d/8+R85mGdnpZy+U9kDFe
tpZfsuVgP/oj1a7owur+Eee4HCKUr2+nA6YA2ymQGYbx95onYbhQVGW7FQjrA/AJ
EbCKJG9+1jR+kOUjw/u6fK2ki6IJ1asQL7mZ/2GeV17FpKAFQ/sP/lKd8uH/qpjI
ZmTXRfSsj12Nqayawmvx3PtMuKLICPAajro9/1JfOuk8HpLlD7GGymIDOmaOa/LB
oUuaH5DKdqVU3AMdHmnG2b0LnhXSFHw+k4HLURP+rF/PjLzF2TYqVbFD+AEhHu15
Qm00tycOPoWSalN8FZFO6i7nQoVElIZZ9IPKRvXHYeclwdcGiBxs/9WNPywzwthH
e5C8puz85Pe8ejxsFFQDfSc52iPZQDiEm9BsM23uAZ8GKl26MfScJPpEyZrmOhUh
eyv1BC+aYaZ/JAaO5CFNrqBlJyKAWHu55P6iA4qQB6Q5fapg3Z55etvz+ZCOzi3v
PZAUgxtw7Q5OlK3/QuiNpYfCJTNflLAncadPPWDQIFKyAKJv82fGNbifGLMCIZH+
eiE19mh9FezUlCCXFHqsEWGtpOP3lp26rsIS3I+MAkLDo0erkUbLpUTymiDI7XWE
CBhnIsdE8GgWMG0D/VRgi3v20fUqfUpos6m+VgSul2q+r1l5V4BVkr6p1DeIgNWc
ciFQFhxyNf4levRNPB55K//INXPcTb6nvzBahedmt4JFar+ZF2cQ8KZJnjZICqBZ
XYFNgIRtEL3mKx0je993+2zXiGfOTPEjMvY+42gXex6H6qf9HtYiVVTlKlRpeKX+
B2Kp5i8NT/9DveSbp8b0V2BOB167GU4CfEMD6sj1niyXumIqJ/nvu6O7QfPY8tLU
Wx27IyItHMw050bzx+SVF75nZAGeB0a/YmRhP55f3OxVN1GOcSfGvjyIeWijGNep
ghE9G3A9bZvZ4uVIyrTspJjKxCTwOqXrL7lpNAAcc3WRZo2NtVTInAOHHRujV9e+
lD0FA+ZFE3gltUHan4C4JHtWHuEXflarvO9g3e2P00e8hKP6X0k6oDxSqrckxWht
fT5Wm/kPe7VEAZjclasKOZNovf1u+5IjHfS/57hWIXrS3T1EOO4xjMCrZfNo8bx3
ch7FdO7EfF0qs8TXygY6j6wN/bwPd5sNAxQP4wv1QJzpPt6LNi+qYueE6mfRSCBc
Gyea5atUR81PM7DsaHdw4zyseF9xk3zsxzgI9cFPna4Yz2GUXH+SfvHLFFvuAcsU
Q4QIWULiAvx/dyj70OA2EFELFaoEyd/J7yTolW/wz9ChXUR/N8H8CF+t4vpcLevD
sJsNV36d3lrbL46BHhnoObArc2iIv8ibgVxSmD3Y+lmRLEbefooAWOpZbFWqEVkT
L51L+1x5DnJVp38C71bWms2XQ3VkQ86o6TAyEMXBBPVYSVEzD9eDdBmBEilXudEQ
lZ8uqdOyjUvVOZ/AH+1pRcJMYN9gFbPo29H+eJsNhQ0kprtHAe1kW2YEdKUfxG89
nyAkIZ5fce5tIzi15DJbtexybVcvQTU5P+BN8iexPykMcZIQiVZ1rFQjstBjcEf7
CcJ4eA7oYsXGJcyM6VGnnw2R15Pm6PeA0T6INxeq6LKgOw2Y5xwOo0OON7ldhdVr
Fjh/BS8/Sn814ezqDaFHwyOipxQUGykX89YIap8TsDSFQu3qlDgLxe6uXNtdh8/1
uuiij3QZL4rq4ppq/heuAUnFIqdkJ7kHvtLLuIjH4IPxH00gwinQBP0404VNgwKX
l+D7MvIyGSzLo7FxMq+QSyQR8DaxGmqNCpwy7bS9HtET14OyFp/VYH0bawj3MPxU
siY+eP92aoaREwQKYVLPBz6fSX5JN6q7GCIascjglbeYIphR8aN7LHinulyNUPjM
epJOfT1RF2q54F7Jg14Q3GU9AfZE1axi7tfF5lIj3oAJ6Dc3Y/h9qQaedgrtUq0f
95uulEqK8lUwyARIZZfr6fxAxS30PMQXKxlzogPxNTt9ala5CUZHuJP6FDEcwAac
BQ3DIDqqFAG1137CoM+u/YM5juJ4N75HNViWO/sV37269zz3AO8N0bO74XSZFE2a
Lpz0EejOAZX+rL9d1RuKTobUl5nIc93J/UBHfajWIZozhXwxg9z06eW4m10ewXMi
z6l2y+hgENtOz+0BuMA0SGB4daaGWnm4SUmwoE/gA42kQquON4yqPDKuPQ5/QvZu
zEoDfSukZdDepWrMTB3J9kEIZf8ph0yITvBRfdrcjwc+SY8Nl+qrP0+yel8rqLrg
C6PPKoxTfdOGJRimbTBvIn0y5r9ZddVfj/bBEmxEeLFDP7DEXQiH3aL8uHfQdxWP
hLVhmxqkAXPOOSYA+DAp0kMwcM64gHEkRZ6l+jCUr4sqLLfAesWXtKcfb9Myh+EY
OWTqoU9GyqsMInirYGNyI3nqZpBwI/qKEBdLsmgz8Y0FyMiyAXYHLGZ43ry4yxq0
ASy2sHX1cK3q4eHVORmzbhac4d2Q8QzhvN07NRIaAZ2H7J+mqrpz9oQgvSmkipx+
+lCdYQnuMOH/eTp4A6KSIpDN7Y9XwKuIECwa5xxzTrx2LG1LiinTSRtwPEtQJM1P
lJoRsMgOFuC5IlGKKplqsCmpP1dQ3PCnzJe8Ehq/AWnNaQwQcrIu6K827klQ25TR
dVOkyCURf73gqs3yGIP9MM7U3szPrgm8gTafMe6a61Evfu1MBKc56lxkB6sYHt/Z
TUQ5AsHyCRZMDGn7saj5UmWtG5aDChA0udopFW40GMrmCND8tNa1oJvZgU5SNuYm
P+CZYoJW1MkfPMHsQvvn+LhIEHf61QssExBjRZl87mecJQ/8YiGzuOEcz0NasvVR
+P+6AT81r0TRYouUX1DQF51C47DDG+tIs/o2AAuvpRBNXm2FeWz30e8YlKecF7Ft
QPhLzlt7R3wlo0RBDl2Z5IYVxHHWS0hu/ILYWJBWj/zU4TzVTve24hX4dQsMGmlX
Iwy4eereqyhQSjuRQa+K51O9JCfT1Cl0z0DMnVUbM9Fz9qFBw61XebJS+4WBBTFZ
RH8adak6CMVPKw5ji8eTDfJorWeP6g1Rjqura25Mci10bCqmeOgiuvNHIDoEKcqL
GOXHj9jg9PD4O00xO5IlRm9KNRDeWd5wdqh4Xvvteu9z6jJFpRkp98oAAiVw4n4Z
YagPaE3v+RuF7ZRpXJX/xzC1uEBztHuTtFvn1h9yglfSYF4fop8/wEpH0g2MpjuY
Tfa2iSd+u0W48Rbzcr+kXSr81LlTRk2eITFA7GS5rreDLwLxVng1BcYnvhXoxZq5
uux0sae4/YaT6yeUBUh6eIXJbK0RtEU3RpHJxwawh06C77K6Bt2/xLM7oOj33JhP
XyXFc/Ema0cijU+F0ZA0HiiK4yqIA+Sr0v3cfXcfKN5b7fAijr+t5LixH+AS+LEp
DDSkQL74Mwjj664k6LFMK8U6Dl2ZSD0LzOVu9+0QK7+PvraAd4wjQ9Ii8gLN+wRV
MSpZmCTgvtQT5IqIVMY4Ma8XZ1mXNcI3VJmA8mbmup/PSNwSi9XU2qwtltKjrLub
XeY2PzxtVuwUb57ZCxjN7j5B3MAexugOCYtMw39erhC/6pxNUD3y1IZJnmQcmhcR
pn6cB2sqEfovjnm2jDQ8MGjo0SCue+gnHcwYBG3Ar3DBi6pyaOdNqheMvMcf+IHy
t0/QwPvaDdY4iX89yfwiq2wyQjImW33GvAXqyAwwtKGhk37ykszQ9jh63wydn0Xq
iRcp14e44/0wh4Rp8EBjyKX2B8gKB1lISgvDKbtLoy9MBjBTp/MPo4aMwe/loFYy
KzbUno3SB65XbF6Nu3ZjfWquke2avWA68F/AVBThx7tgyUjyMw1PSWQNsGYCTzZm
DZOWfEyMrQWcJcjgDo9PsvBhtPOKL8Zlpk0cVXUabtpWFFC4oQ60oKWGRFcmQOUz
V8kN3XBTYEeSvWuWxbdm5gtAOFgsgPx9ov4WhvuBm8anOAsP+NbpMLanib8NlbkF
TcCwn7fP34aldhdG8n2E1g5LQuMvqe66ZjjyH3ln7mhO6TDuJ6GIkVjG5epP62b0
YP6DEG3a60pPK+yo77IOAEj3S1F9R3i+mwkFX59tXJNNV2eoQXDb/RmGICwZRvE6
3GOnASNxkPXsOmpIrbs6/NgKbcKDOm/JFIQLLS0nJDyYZqTsPLpxhNScTFQhAfCE
PWbden5QrBtu2Zp1l2lz8sulstVp4i0RQ3y/VIbVVcQX6+3UnRuPGnAH2kW+ID6U
86js1qBCWTzENaR8zEPoHqwJHERB1Z5au9hj8R4RYUMSami9ZPb/jMn6BZ6jn4la
tVly29518YKiILoW1zKGYC+PyHnbtw1K+bp2zBOOkMQD7JOEchCw/3eH9BAEUqHF
P/myNktUhRifWH/ipai1Z2CzR7Ha5Bi79jfmmfM4hjvj6ICU1E0IxTlT2dGaUS7g
uUwMYF33SWUaN4S45DwkLjM/IfgVsHaRB6Q7GgroX3xI+sraRdAmOXUWIkrTScFp
N0qkxK5Fpbcph6LROwaX3McRfHn5CrqXiY4nMshAQjHGFrCb/qIhfod74SVEKJJb
bKmEb0guCzCk2PBviguGUUWtD1cl0fL4xBrNCFRiPswkL0BkD5p96mdh3QJS/2Sp
yzrLS0/3i9FFUhSfZWaW8xT5zy4mwP/Z4pwBQTrEDTATwC/6q0nJBpiVhcBl8uGV
uyRxqXDYlaoyYjJ8m+VkvP/iq8id6oCYk2/bUhbZVEdHjbFLrOYRcHzQzWpGTCGg
GhEl710f/wulNYDRR02nhbUfhf11N9M7x97Z6C0E9AhAU4ltPLM3Tkg7zwMaeyb0
NYVivbnj/VQQH334tAAXLDtW2pwgj4cEiO5Tyx3BCnQYtnBL0hxlkYwOfI3HSMVn
xsJ2EgjDeuTAASy0ANoDyGtBjM/lfSVYW4JthWKA+Nl+DgWpyvKDMWL5py/tBFbB
21Fq2Xt/jvqYnkE3Gc9tOrLFgoNiBT4PcK0bPiADxpth6yMy+CskBmpCN7lZCTXc
FhCuOFLz/HCYWW65pA3dXjvII/ce19T/w9dn+WbcCVCopGAFTfpcQpzu9kNMHaQE
YZDcl62lOp1Gw+JreqgcrroGeRJMKq9VDSLnsGd4M8mgzbCQ9dS0hwIaNuwxKViM
l4hdZdCBFREGOGrcKrWQO6hMAmoq/saTwe17X41IdGh0/RgVXGyToAKUHiWn+4eY
JTewFcrA4XeBBf/SWV2ZUVHWJmge1LAlIHSeU6OxEA1SI7S65s7Tu49rjiSFs7Z1
f9NNU/JZ6VIXMjjxxqH8bFGURtnB/0m46Ju7x7ftlb1iHmgso5q2GXXh5Ytv9LcM
PdKYzi3x08TcGsPkr0EqiPdd6YGq7uoxeXh1F41fZhUBwtY/XMQKAgZWaeCOYfAp
1VbWo2c080Agmk/cFedbgy9uNoKh/ThFYeUOQjzQnD1SOjZF2gyazy7XFtx9Dgkm
mtvAMvQBLRSg9ikn7K7fboEq7bQWCWhLw+ubK9/Urwkg1ZEaVU/++7WpveilC5zN
2WSfmdsK2UI+9zJ9ddd4O2n9APPTE2rJq6P9zQXee9Tum9BI0QV8ECUsYdEGm7BX
JH0/4Y3YWtGIECTzC2uKhEDMBNLfKNWNgwoHOWGf1mXgR/fT6nAIkBvVhA8wfN9I
XTE4WyYA9ciqoR0I+jP6zMAsxvMDPxTVKvK9EGTwBPbNcjU0A4n5YDWrCbn9evc9
mZc7ZGuE8Uc/ec52gmw2cGgirTY1sBabcjZHRAqKe5jJ9UuBrZnu4z5Nd+XhZHna
sUmTJ5D9vu7f53LOI/OMnKaSMEq6YGOmM3axy5QWUzigFbaoeMph3J2wTPmAeGpB
LroPS9vM1cGC6HRPvpucpxJIPSniDcuNETg9PkUdpTLV480NNb2l9Vu1wHJjgMwu
jqIrCT/MhxUenDJE5AdH04Mp3VniQSH9eI7iC2I4LTJub3xo/7SKCnKZPb5rxYZX
RsrPJnJ3M7L1RIj8rElPo4/1DpWe+GvQgEePqU5X0rxRZC/wQ0k+pwg5+juwSnRj
0oD8crZSsxHcd/dz2vRqLK8yDJ/jJxn8is9sIEaFUPOO6GOm3LQiidBQTiPHLsW5
1eNPR2EcmA04WrqqPI/DB5uqEf5UTzoI2hq9u3j5UO/wFQ9f/uPD6qLHZBTpQDeN
wIWpGsiygYHbtJ6/lnfoycsOAWzlYUggV70hGreos+m776iVg1Xx5924HWOcw16H
VdoCCURTHMY8CbGF4zWixkLqwjaUaUL8jCCuO/HM+2cyorCTkDOfIKvXYlmHlwrt
P9pUB9oY87CkCqTKeFJIB8EMBTZpEyaPkkK8DkKD3WABRpbPlseKSYpxnM6MCBl/
IUfrb55o7OZwrDRhh7tJXSUYwbaxXvoEAha86k0DqKv7BDjUEvfKf3cQJmVdZ9Um
NrJGldpTIPx6IB34yOSta345FB6vPAyCTR/D4VBYjFBh1MFwsUDL3W3T15IXR7jN
1NBR8DfH+EZJ5TE5QYiu1+IQQ9WNk4CqkLt01h0hBBhRGfmlbY02u9E4P6fcxwaY
1OYVVQfxQ5JDaouj/Pn2zXPkqEyrIebeBkERqwHACGGsbfcaucmubZPnZb5dJ0hL
VdbWpUFUtfvjJU4BTts2zSxBmx+SZ4THyrlivqjmYjWiaLZ1J5kNRGxGwb2SeRah
zA/xGgLBeMm/P415ZiI+8OV5SCA2jGU+KAGJrF97WlmTZ3C5znNxNQXb6am7FqqJ
5HOz7Foz8eBFYn5bpHDcZr31PIvXWtMeMiqilC1uPDyzsW4FaQA2MYq80K0KEqVr
n5MHeftr7mdXLRsdz3TfOSsNsuYCCi3EMe5vi20f4h8q/tQJuovUbUUfChiPvXLz
rfv2N0bhAXU3q2sqq+JNsAzMZsYFWH2zSpf3TjtvHK5YfKGZQjm2GDp8nvlSZ147
qxEGOGsuz1YPo/aqPqWsLzwNEH+tiurIhk7UAuPG03fhDcouvBurJF8jEOdCI6/S
OTs6H4WziwB4a1y0In+LnqGuTByfwNKgPv/XXGbCViRfxXQR6uq/mpUzkGobnXu6
lJE5Fh1o9Y1av4ogurA67nSJeW66MUoZqTibL80n6d5IlHd4nyyyHlpdDpcfJBn4
vrGJ14ph8/9XdMrMojB0DtKdDfcTmugcc86NzGFdC/gUnsK2ywQbrAw6K+QP2MPd
BANwavA769exybLMiv0KGCIX+vmwkLxNofP9k7O9uB2P0rWhuxc6VNEcPgfK6xsD
K+PnqNLIhquoiBDAdsf+p1nfwtpJxukgB3+ON92PNh4HMlKCaT4HckCDkCtsncd1
E9vecQCaJAXw3l8Yse0WeM8VkHwMYAA0ImN4YguBH7ISEPUF8/BiRAKZmnp6jCWV
lhQ2/jKfQPJQHQ5zvcgCqDzIbAa4Fve+aRA/pguNpbSfhWYGcnd1wx/ZHdgOE3YV
TCyBmg1u9gq9ZoLuyUaVG0H+FRPIb6lAxtU60LcLb9TP4FP4fODn5HquMIuedUG1
UfQ27TrzN8BimxShbGWvuyiTh7C1Zenxfc4XHifD+M4TZIiRW+rk+KNUb0C9u950
i2ZBkuq+WTWGf+QsGPcBcEz0e0bPYcZml1K61I6XULbc2lZNjBFDhr4mmMmffP6Z
gcb6UELQbxcjow/MC1RDm5gKhvxI5Z9zqBfQiH3Hgqin1yOIMxOjfJdWCWvaqud7
Ku0qxuCxhhjuq0G7u+FMVDNjVMTmBXalwQDMJUkBbAF0Su91hslTWFIdY8ZN9sNy
P4IoE3MMlpUxUZSrR8icMP6pFfffsY90BBNGq+ISXqETx4JQnRVkAkNGhlco7miP
Dnja4P/u4FYTBeYtT0mNPg1tegDOo77omJo4085GhVwV47rJNrx1cZHZUDtwneJb
RlyM4gamSQL95qEm6E40hK7NN0ygYObQzJciM4xs3UOxEmPU9pithKyEdM43bC1x
C1IJ4kVqqHXItCw1P7B3DxeoyclO9Li2tEsMYlcerlY7IKI4KCQzbWjQl0pTLQCQ
5Z3oQBp6ofLVit3a2mBXcaOFhQVGzOtEbkvL05FCcrn2dUk46uFN7cpBwJFQi0Tc
NvU1cC1LJy3WEURl+xZ3cjRHzlRKRFwf5BMb5G8P59txlwFbVMgMSCgfQULFMjws
MNBg7hGAg9bqYIAiSgV414+kdQTznt4GlfDFSrTIFl1RDNM93KPwjiUkL//RKISN
kfTx0sd1qM1agdbOUp9XkJH8LQ2mU7u+FzADNEFL6NDh/snw6ctPqHaHa4ZSKk0s
IK02ALGMn6dwoCrPJZku0xSU6/7cgLLuOL5DqO+aPaNvvYGvEUORrL0H5VTkFrFP
Okh/ZVwoqqhrr4j3vjwDOPWYXv0NjK9gc00K6GdDBsflOR7FWHxuPrPYkswF6rvf
qVxeVDi92Y6aKcLgnNnW8oUaurEQw7TQ/ITtCTLLwy8JpuIHxRybJXa6WlGqRcat
RSlVi78MW/2x2DjX3eF/F1FiTjSqFokV1CDzs3AOJsdyICHBloDeqbZqnwujrIdK
jQV/kqE2HShBDELtsODEr+tKArB++NQVaF32TlAhLbbZ4z6FcBCH3FE2Cx34hyiK
140vyUXwWhLq40SbhFJobY1tj+6z7hDwJk7A213/HqGkF9v8rsTF715WlHlnZMrb
jI2AFTbU+4PKKtDt0XIITwGFhwMSG45yokNQpSqUTc1Xcr41GiwDCwUr1wd4T0w4
7PnduOEF1xuZGo5ZbObEYGBfkDHjRMWvVSljSYWYRy5+b0vHgFo53lYMCKFkidMi
E5Krg28L5+t9snv9NKBJQeTEICCRbCwu9a35yMRkYDfgVISLTZDrm/XwgP0Gkush
uC8jOlUwsIuhgbukez39k7PbSJImhix5g+3MGXhngPEjscK6cccjaSDijL2BQrEn
/jio4mVcjZdS5zwyGhKYKuY06qtAutQAk5DRQZksO2dQukQzzvi+o4Roka5NrPIu
sny+Q0lqjIVvEpENTaAlScEgPhYHBDJEJTQ0XcmYLEpYyy/kMvaTbM4SbFhIHt6S
SXiM/uLLrQY2QRcOqMa2lKCOKFmSUFN8/ARyes1D2DNrAsBGWYp5isl8SvB96fzw
HNl8D8yUpJjbPkU3B0KVvHcj8XItRtPWbr+Tydsf092i0pCYMfbRQz5DdUT62DbS
4U0ZGRbzCkSpYzOLwRfNTSHYLQVe9iKvZAxHfU/NKicHlOf35QY3cSoZCNKtU1b6
46X71CbMnR8nutJUQTEGE8HlG/op9r6xsYeEXzdtQY+WSdKSb0SgjhuRZQHnYt8e
FR7OlXvXieV5ZWdsaXNZ+zEg9Bmmf1LMoFI5aBkOnk3ekjywnBA656rsXvqpLM7v
TWEQiyYfZobe5j8NdyNfr95tr1XNxHvFYV21j4pCqQJWF6orZhu0ob2WTXu2RH8S
z+lHI4OGdDGiUIuvUZkjWfM105T33oCOqIFt6QAGkIZYsFM6qOfy4xInRvAL05RU
D/Mh8iIctu1vyCe9zzx/unE4SgClShiuq6YiS6U9vkE+AIdDcVF7spFaM2+eiIm2
5ksZ5oPv2jG+lFMEQO7C/taZSL+vsjESxj4SfcKWbnxjz+WWljPdYfMO7FzWBbsA
EFz7GaoYbG0YeQR4yVbQYfSKvJPQiRsZGfBiDnHQuDdzgSDfCHA3QtYg0JCCyc8l
Nm/dy7U8TZMFWDwjNusHEsl1s/EV+OCqi8K5lMFidGxP4jq65BpA1mBkmPqQsHxa
r6aCNI+NmU6A6TkbuJqUR+ybdcUxIsI6Lcdxpc8WY0Ohloh0ztT/S1jx0UIFfVj/
CRFjyk4fPAP9FwMph0/+G20gKO2nZx4KatSvtCpO3VbMKf+ibtpH62YR3m8wc6ri
KXZuEYUaibHiP0rlBXXGYryFT1gA4ma9xYRtInb8aIiuJrA6ECJkNwlq16CnLCz5
m7aU0/FZSFAuD2PUvMOQk2gcQuIp1Q/9POyQw8deMaiZ6vwYsGCcnudAPxDxtg0z
Tg500Qd7DvK5aYUbAKjEl9ZMxWWJRfQHlth5KEWO8qoKidXOL3xPR9a587rd7k95
6aKnqTZoVwTQcO1hIMiH/8BhHUHPwC4YcWNp3IqIFWNY9pFGcqeH4dtaMAfGmrmh
uSb0HMGik9Ee5j2iclFqPCz12s8OOo+eupjD7B7oG84zOpZLFyL24MP4u4Xq3uLP
lFqkk3fSf68ll1lpG7xL/Rkrz+aTmJXxwF3bTSlJ8B1QuPtt9+Hz4X596tH6Ec7T
k9sTJPVKJiiHnQ3LgnSQzxxn47MSEykTV6hMlZLY6ugYBjQtGVPGNsUTiZ9Ox6mI
V1FeNw4yS0CmjXjBQOGb8fK+mlgvCXchz07Xrs1SWhELB20j3xB//WUXPRQMcFje
H5UqJnjw1G0jZvwRmiT0kYu78xGHozRAtCiqX7SgfAQFFLp3UFAoM4uIyGzd7HLH
sL9IvYkwhFVnYGHNYJhvriAZX1MMI+hFOcAXgTa08RuRshAGlF/4/eoEoqqP/WZe
56Pz5Z28ZQTPJymPWytLyVZSvCo3pXriPv+MnMkiD+gjU2l6XO/5248jcgYyL1eu
pIgBzWU+0qPyBsfOmwm34xw9zacHgIHEwmn43o1HwFsO3xAlBCOw8DxiQNg/HFOr
zs25IUntXcjsNk7zrW6u4KcsqjfaMLNDjKjpiNhhIIYw8dd+YjklLTOw8s74s9ii
1TEhCT9guH8EAu7YT/W1Gpm3JkKDJT5VlMWZX29SzD/wz1u5dcEzTQzfhypWd1Y6
r6ACYeR2UZ826I/5r9A19jATczrJepOdRHd9dNxlju0p76YKdAVuKQRqI8DGqgj8
jlMMoLz3YZ0sIXrUcSQfIApY7cvXMU+B2j3IwHJ4vip+uJL2j6tNpvGce8guPsp6
M1jAKRpuC8uusA7QMH2rzwaOw96yQy6DmEGzxXvxJOPG90/APv+w+62DhVLMMYk0
ceDoCBwRWWHP/0KXQH2TcTbzgywHIyObkWCf4oJeIS+Ltf9qEiTrPT6VlujYh3Vt
B61yO2iug6PUw+zRWhG3IHv9YucuMlVPINqFleOYRDSAHi/vWV76F5OdtZurUXrL
MxCkvKiYlQTK/f3ba+mh5oyvXaMrWX8cSeytAK++djTwxC03UlH7TLbC3WiZhyE1
eoPNq9aMBIJ+2Jc9kTyBoSDd/2AHVRYQW1PLAxYick1zipJpFg+tj0ruqoZN6O5P
7yCdtKcEQWSb43QPfJvE9wibGjD9IRCOTs+CwN37QwdlpZ1RCFXdo5dcKqHy8X6f
CHVn/gEfHIjAlV/CE1U0Ewvq5uyW3HJCtjAhKNXvpwTpbKxdWYRiimiRnAKY2NL9
qYslh1sJNqakB4j22TpVnMNlh34c+ExPk56htLNBJT0CtbBnJrsUUWtAld3YTkLQ
ZRgtWMjRAnzdw3mIEC3dYSuq34PipHYIXAI1BVtQAo+GEUDNnF20RyBlhhmGowrk
fv7YitePdYWkTV+uSjv/ctUFDZovuF9jWDEXyA454Z+uM8r38DAAH9Jo05iicRsB
Hi68WZG9UDA/bNBA25hWoLZlwLvZTXx+O3UzMgaK2vn0hNYk0cmPfv1f2sffq8Xo
Do+VJ8piC9qPL9AxHYd+oQH8LAHjXSZV+sPSi8OwrdtCScHSBlA1tQpSU6+8izIQ
JG2vPOPORlPs+8mEkcn9jGAqvpI1ijm17qxbbXqiK5zPjb+GwrUaHKK2nB0YMqXj
TIgABEg7Hyl0W/6ERz6cpyB0PBjKuomXTNWtJiVjAAsy27BmO0GQELsrG4DOkkgA
Yr5j32KW6JSGxvgeHly1gH8o5IApfr5nR1mjfFnL88vH+dlYWE2Zn99qcn7wduMt
sY6KEFlmjmnsii1J7UVdTMBq8aTZUP1wRl9id08z9bGRPec4DiMZ2bHHk/sIdA73
xKFe6uT2ivPfR+5iysHUurSDWixeND86MgoJEyXgjC0VGXz86pr5Xc2XG9CVDgLb
SzkWgmNtZK9NqAmYKg+PGDk3uoOj1bLO7+S/BpagkxDXI6boABqD3EOs2ngJrfQ8
l2Fv/Jco5q2H6QvLykpA7Z1RWg1zimdBRvx5f2kAUvLaBP2MPx7OgFazLNyEOLch
EiTRWLNhPZEUmiX7EkVswQemakCw/0MBx7oQ/5bv4aS6auQxToT4UYyencl6qw+U
oxGa6cWosJTyPhGZxrHAzdAQa+qrqWfDYKb1swLwKLwiVzZDsZjUBxsqgShWQfT5
vp4fn/Vynr6UkyQtA0sTYh5If6IPx6fo3QV6wBZIPzDwDfL7nK9g9onOKXaryDEs
HItEowqzEMurbJLJI3DVHbdafUe/khu+y3Dd1vwFsxsYuxM1kQmJc6xPuPDRn+g4
FdWAeN1v2cFjQNnB4yvLgzmC+WloLxkQc0WzYvmc4DAw9yG8pnAtmf/HH5xrUssO
pmbqtwIo30/F1k4s7M+BphAUrfTo4ZlqrZno7WdUI1QmoJxCRvvFyH1idXLjaNe0
WlL5znN1pNy+f3Ql5GiFwujax9pG1CeeJwjFjMzNd/kEFuwnLMQm7M6Ci4LwJBSg
/5b8Mq7AVEXMWibgNmt5SMxiB/6v90V7Cmg0RVKPl47//Zg6eiJVfdBRHo/1hkgD
YVppCtjnPntkjjOPnnHCIxlZbT/zBNJhwtGWhmYVHDGeR3c+GR+tHz3xhCvmyaB4
s7IZAqqGBOad1B3IA4xEVhkQuGbOsIcH5y1zzYHhwOSOCbEH6Hlb93cgaKB/JrPu
3Vhp4hlTINNduzleloiRzb2xxx9OWBwMerrhOXOyO0iQ2hUibsAXtlVBr22uOLge
64Rv/M7qu4iPXPAAqEb8B7JWei0L2q9ORDJXUwZRyYj0aPDwTAtHXxVDgBEABGm7
/uLtR3zSv4maDqQPjmZklkeyZ7/75045lszQTGMB6N+9Ku2LUhEefIpPBgkxqE/3
mvLawW1NJMKL5Xu1f1ra14QKOHnYZuYCKB4Oik116IrPgGVyU9lcxMIURLsdumLx
zuyoeV0CnPYvuoJILy62N4Npn36DmbHE3vq9QEZFOjnvPBozA1io9c+dSBVkszsc
8VltX07hd7nxL1MC34n0F+PzHolE6VMv/aHIyQWCwISk1r8gho8mzBii7v0YI4f7
uLKDLmEWZ3kPLHeAQzz5/fFbR1IHZIEHoXXliCW6pg7J9nw/owSP3ZN1FHyss2Rt
8dym3NlvKyGpxX8wwaQYSUT2scYOmzY1e0ERfLYNt+lemQy/SlWRTD0nrkXqQU9a
4ce+wlusAryllYNEFVXbdqIMmytNBRYrkpe00otjKggA27l78zwTJVBsxk+9Vg4v
lcwH0MOOTU0msL39m0ma9moWzD8j1A3cNyciR79Vvq7prAWLdQ7wqS50RC0ijJhz
NHwlV4HxZtFyUUIZI5PmluoZmkKyN6aqy3diXNdn0sjw8JARoxzz2KpVOq/fqJ3L
ReOCv9FmpJ8gH/IxypJT1tFlJt+DbteLL8RW4p5BZYG+eAE8oXYgm+r7P+WWUBTg
tHH8+x2Ic96XnifKOFqijYuD0D/A/JUragO6VlkMMFdZWsqIPYSyDggVZPzSZ+Ds
E5BMkD1Rctkkb/7zaf5JmaZ6teSHH4NS2Ay7swmB2UeqKNycRTKH5Hz/OfVUxpao
+GGvTvY0OR7amdD3xra2gTc4gYes2jVD9OTAHzGICn+WZT1ldPQzOkCjpI29lEjT
Ypdfa3jEWmYhH3B8c4I940wPsLzyslOevzVv0inowygiu/14nqwNigki3DRyxhO+
wud8ksBeiIh1UlBrOm8h4SeqGcRmpOg3ZuGOtKfktq9nnrSjAelQvBgYXWTjk/Up
TUfZljZtd6j6BycG47l0G291OYMav6p7LwQ3zG/1aPY01g/WlTGFtOUY5VP7XYHk
/tUtyCnQo0HzDoFmvAzkX5xee3k5LoTYglxmH5MVKiLkQm3AFuK1lP6NboBWJdig
nRuPs1OPhAbVmOnCgh7B+7I/zZKDJ55hqA/7sSJmvNqsFvObtuAON2Ru1TX8gdnz
5hTK0/azxXq8XDOa1gag7qC0HMLz/g4cjo2KtH4rSV+wDR53+jf9KZ8iw6HYjf/g
oPgkYMn5j5BiUZAmCAY5OukC7QVhQuclb8x/VWr6GSejbqq6EVxz6B9Z9r0y+W/C
qOQuPqsO1T9TAjTKj/xh7KNIH3r98t+vAke/PGRn+YhjCme7OPHEJdDXHH33G/1t
815M92rAizEBCYCufgNeJJaRK7RPJs3NEZlQIpAQ5/uLIvtqMeVhLHBCkp1d0N+H
tBBaerbIVJqC59T6Iz2y31ckJyG4+S0g9RpEGrD3PM5uWngoejkl5/esl33XmtxE
OCvXg+WGNZYch21ldyCjLdZfuwUMgt3NWd3CefxhbYBhN7BjVTkzXiJoTFsbF5uX
EYJDYHXSXg/XpqJDOTwGz1bu87bGncBqzj64R3l5ltDL6iH6nBVacFSFVY9ke994
0I/Kj703m4Rmhd4awXqSdQ1BLx3grWCXPZ7r/77a1186d/PEPs0XV+0SqrnjE4U8
3vkeOXDkEwNKpGRZzjHC0/5sD8ynvl1x7jdLePYo6RuatI1KTO4TJpRXOJt8rE0b
ZtCupmvor/EgAJCXc3jx3GGUmIysTGQStUuzQccgh4pGj3tN1pfpu9kHw7mbnNmT
FtqShRRl3Y0qLURNapduenGuNGRuklUrYGS6iH89tDOLRURTRnBb73g1a8nKOkt1
IKsIFDRi6RfCWh5rH+7RUvY0gjVzWVkgxxNxoquUm4FgXJdDxxjL0eoI7YodGX0l
Yw+84tOTciVvWP+FAUbpe8eVENcLfPNNrjS0TWC+2yVwQlhKxXgLtbFncro9gFKk
wxiQ7IvvcOW3q2i74Wf1iltZv1pQdWKN/PblkujMujnsNK0vzKWgCX0ctPTt/DdW
ckR11f4i2fi478sTizThC2pMv4BZr5Vbt8nZDvdyPOMMzEsToawNGLoD11+m/tQC
ZdTahWANXCvThIKkiPU3Kv2RBqTyJjHX4/jTavKzT99lNIuG5EEIuHux4f+Ah6Ze
X+YJE4gjc1BK3tyZCFfttJVbGMGH5JvAhmYO8PzH0svgsgaR/wt8AzusGfmbNmDv
9nllEedqjhvLDo6JyhEKqzn/tQ8bqKNrjSribkjOa+ozVisfC749V5Qh6UCI+dKf
j12TVC1jBKMb2N9tFV9p96Tcri4/mxbQCfnutSx7ahtdvZInsOGkKGmXHb4uXqhW
FGSKJv/JsuEKBV4dWaan4s403NCyOOn84iHaU8wbFhtSJaHd0ouJjomAhlHyTAJY
W2NBHzexGIaclCOLPlOtGPSrxw4j9kq4XQRhK5Y0vBbUilpoGNdl+aTyLo/3Tsb7
cQJesfs/1L72i6ND4H4kpd60neCGo64rAG2plRK/TeVgzaLVDXq8XiC+ki+4cCp9
G2K+WpkTf9+JMrz/6NruGqyjgC10r7rfOOQMjAw6y/KcAtJ/kR3arkF5NpqMATAQ
1rdEIdIW9NGRHs7v0wIXNnZ5oCVwvR+thc4tOm9wLyN9NrU28eZZ5yuu1/yJMook
oIHSPhcuEp+kntPnO2XRRBdFh1Lvs+23sPY1BJcZNPDJe/7ZyLcJiSfrtg6gzYoe
7+B41ZhVr2YWJE0n4Mjb9NOjCz/st0APA4MI7myafkRR3ybpXfRf6VEmUNfrfJW6
SpuJxTpJ/A4J9dF5V/CRb89cMHz3pb88x6zed96czGUI++kP2xHWrKOi/hX/G2jf
hUDDPcOsjVEjM73fZiPYMVygZPtIWc6YdaxlaRJCKHvZil5M7ZdsBGH95tw6hfOF
nnZu3a0+HvHP9YMo/Mobbd/+5VkTSAu9oIqaH3BwB+VPOB6bAaz00nW8PBXrB+AW
IF8Buf23oAEVe8pTQS/t73e+7G/Np13JRNNfba8BGLbZJEUGCk5e8OPNC01UxrcO
QRtZm/CiPAQjbxs3711Yr69mDOBTSOUe3h+o66fOxF5HADtQyHPKiEE67td5IR/m
9Odke1/XGFdFKdgRza8MMEuP6B+AGR7OZ++sKInkiKJ942YoJeDa8GCNwRK+6hsN
bK8wa9Pto//VTpwcuiwYb3oMAWcOPy5dz3JA+imEz9HMxmvSqfyNNDbxOHgvPVk0
bpeLfdzFOzs5LBZ84bwLIXBnvUNlqsm9Jt6xi3UTWnSxGSKH6CTjwdMDxxwM1egT
WGz/qoMtSq9ytFOCHKRY4B/qFPq2WwAG0foOn8wzDWYJNkeLlzEAs0mhtfKLZoUJ
uzY/r5xLVzHsyntA9xYGLBXiA40yse5WTtZxYBOb3zJjFXcXkDCzyq1lq0FinOMx
mNyMF5LTOcN4W22ecWF/pJfzJzTc46UZCWtqY1nuh8ybdtLXP41oj/nM0sbOE+qb
plqeASZ5AtANqMlAxmNYRwsvi1miMWKWC4nflxw9Rm3Ev2tJu27PUwFqdddYS9nI
SzxYUMXHoZpUsmRlYGCCNe983f7D22cfrF1RVb1tTJQELPwdPNgBiVy3IVk39yte
XMDHYLDXzdrTk1JU0DVVo01SV+8YGGfwGOhDQULfIiqM2Vgd3qzFnQ2PBY2wodKe
7IlwaW/B4oLMaNrFRrQE7Z2E+/lzdSJkolJhKWyjwD+O24vMKGu+XXWOmYQGdLJn
bKKwICHD/HrDoiTfH7iZbE4HzAAdUCWIp5/BOm9sotTDT3bfxt2naZ9b+sSB+R51
ZhpG6h0VLOcO4ogywGRrvQOlwdzthZZg7HqR/1nHBDghTFKYiUw505Q4j2gVnGUz
a4qL2os/0iCiWB2jzUNoH7l8L0CbSZ8C9cfQU/HjzZTau0APaXhiecetIY6PXO01
x7mVZzDfn3tVIT5qkKheOXhNb6W4G9YKN9TG+5Gq5Bapfp7TIDlgDw3TyMGyt+wC
Njgm7m3FADFyWZ3jXxQcI1cTi23aQMT4ee+fXrWH7hXcu9bHgUx25LKlEPTs38qA
9teKW6/fnmpHdo7qV1AStVL2SMm6UFeY/VkEj5MQ/jZ01CYHRvFXWdbjmF3ANjpF
M3nUxwKcggncR/O6NsWOIMyO0CgDJ/LaW5Jsawlp73zbcMToDMS3XNmtBfKA+B5c
e8QXoHs5A/DY4VQIaGEnfKY+x3551JFB7/0NGtiosHw7IizFyhUoYN3UpaYNuUZJ
UAOJnu6WMAkNRKOthMnbobtSCasxfkKi19mJKY45Gm2dkeHuhtwjJNGIZOS78HNw
Uj5148sG+TsaLKwiDH1uwQ5e7vNrp8e05YW8qwxlAaEVp7Q7ZZiq0MwfYIlsO9CS
MqhMd7z57G6k5YCiGSFPYJ4WBie8kGSql5K2EjmnCoAR+J7mpsQwK0u3JL20ab17
9HennzRd6fTPUhoF8vZzAN1N+BQMEi4HTcXCbWj75vV628KaVb0LETDhLhIDSArO
miRIXHeymAy51FLzdE+rEACns/c7GMo1sJ+5DhG/GikZuLlnHGYwHm6PUcHF+fIU
n5NcE+tEX36+h8FkX3vy5cgIbSx/cRaEypOQ7s/WjmpeEK/awq9bmKhG/pNamaSf
+pzGOHsigqPGhl7SDhXEWPTR8VuC7xLhAlr41ZQMc7/8biY2ghHS1sVVF0C5CcS8
d/gXZkYXCXZiOZNQiHpjpTR3Y4JuEORiVfuqeW9ff8epIBfHbTkHH2NJtcQF5Sq4
DFzk19jb4YcFYSzs8IC3lsTMvSVjZKHl4dWb7GT42JXceK9Ixfrh47faJv8Hlgb1
1ypYofgwzO4RuFUqjp37anL6V9S22HZC4gEmq8lcqOAeuvWYVCWs0fX/mSDpoL/k
4ffJwv9Y3YIRlEGBuytJGVOp2J6J6EXAjBuZvs7JcUPikugGHUYAtqHZNHGhkKiw
OetDlaSbNrjHOotLNEqJmr0w1W/+GEk9UhlA/UmzXh+PjSsTTG+9PuVU94ahTuTy
dzVMoLIicWo7UpGBSyVvYk9b24KXXMF8THsYSd5x2hBXo9mUk6tbll/gIHJeiBbH
suL4KEiutC52Yidwkh91xItC5fEdvBynoVeV41HzETeu75PWXjHuSkSUc1Qq22cS
Quh1VunmgUj48fibEPrVA5ddYY2j4XdFCpu62HdRuxiJcoo6EANeGiOm/GIuRRW0
V1CGXcYEKwfZZPwwYzVJmqjxZU6FRyoeyqVwCXnf4K3KXB4LuouHBIuQ4eUPY8x3
52E3ebJQZNOYgMQCPEe5uU1hiDo/t0KC8vsK73udWxh6LQ3akBdJZAiWr+DA5puW
1sK7No343RxIq4zX9/t2xcTOnaB9tJtd8DcvQih94BRO4astxRKt6fSZpvGcp/5r
mt39pKVwqPl3OoS1DkI4DevXFE+iTWLxdsA92+S49TDdfd2ygVSqArjLAv/6paYz
tiX+QNnLPhPxUoo1XIA1oDbjhMA5Rwilc5JJogr6l5KEOo6B6oxioVAA9iziwmD0
Y4sNlfPFxVprMh31czkbh0lnnRAItuuBfHGc3+nJ8khNvL3yDSI0n3/jmhTjIb7Q
utBcYmAqye1XaWEByCpJLCIm6xfxNQL0BjGseFL3jCAfIVTZiamfIaAsO/Duil4l
NsqeASFa8OA7j93fr+AxWv0w877D9ryqjt4g2V8/RMWjtV3hpyRV9pss6RWcUVgo
2aobhH9JTYPva2/EA2M6WuIBJ/qe6jQdPwudiLNZqS3JQR1PkbNKFGcJTWRQ+kVJ
vbFJycMLShL97I3jHUc13zrYIEpY2MubPEMdVz69Pj5blNdPvVOUJ2sgwDbxRqKb
V+AhYLI/Q9nb7ncxMnf7bnIOxuQfVRgO+dlIxkNz8BojFz1hsA39o/98EN6qySnC
qYD+MGOKTiZB8l2qvX4HjBXzD7+grPG5YPpHNVtjSWDwxnwuyhRBGYTAHG4zeNsd
B80pJthju4NCnj/I+ghpRSmFoSlWWSjopWpUFg8pAimmjWOw2udlxonnxVp1oWwz
NRNv8qDALzqd6ddjBqZdoGSPtM0aMSWeE9bNW1Xj4XUY3YNsyd7t21dgPLfsNe3G
AzvIhUHFO8uqls2xEKqgKBodujN8H+XbkF5CJrQDJw7QGwBQWUmxslP3v5RltPPf
zTEJn97yM0uQl+1Xh/OsOacR8cke1FIQo7JA9jdrIzNwULJx0hjOdZEZQ/mxgpAe
WXg59wjxfWMnwp1c8ra0gTxdYvtoLKuz8FpXBnODhKsdiKybHzW8qTONYig0MQxY
rrX08Z1QoGx0jxzc81Y3zs7SYwqjjo8sWpLLXYsT7+Tp9I+AaEQasgCr3QT7c7EC
TyVeIKxM6cs2lV/3PpOp745F49n7FdZ8A86hajxvpqNYhEjOhN9/ADnjCQ5bxZUP
g8glMZ5gNFDwbK1wdaYQMjA/qzRoOxDMLKDYc9jXO8U9afMQvJmA25cMi0BeOA0F
FVzEw90fygjwHOvDtJkSQVYf5D1evMmS0VnMj/ro+AqZ+uVZCsZ0Lxq82UCaCvp3
RLZsUxLBdjBxU+OYm8nBV+5qUUGeWweeTF2gg1LRgBUNq1wTk5dyVvLQNGGDnOrO
RPiIILyYdKQ6qop7J5xtz6+1gFwUQ/YOY2PDYUI3x1UxO/wlSUeH8JjrC+NUZSqc
oDKcGYtBl0aMKPTKF+MxQZBkU8uCKMuzytOvNiKky+xNnidIb14XmDtMP4hPrcYs
eZD0Kb6nPgUw0qNdQ6zj87oDSDiXmuG9X0akYil7hLEXKCeC0LQ/lIW7wbyVAVgB
cdLwJqVjox6nn0PoIIlCCMt/WtHPTzowJ1VsBnqyG8Fd/3+Ab41+aM3ccHAgKgEi
pKLvJR+kotCMCHGDDmOW6EWVcVlUG748iOKva6iirYuF/RLWXcstyEDEcfmjKgSz
kBvF7IE4X+7+zJ0ySKkoDCfL+fns8LFFumoqx+zc9VLkwDi8nNQdUyPuywG6I3vz
pI62DJdlC+K6g5R4K+bWXr5nZBG3ZITTK7NQoQd4tODEqGn40I7Z4m+d57i0FhPA
NOOTGeAcPoBmO+tMcz3KTRn/rfNFAHtJGVWgiy29zIKCp1HX41CCxOd4i/Qo6Bpc
xCcuYKdcPDvleThwj9cs94wiEP+KpxvIEXsxcAUgD8S6ItILRLKIkm+0nd5+bI/P
MZzNiB43WXUiAkZBVkLC2vJMNpr2F3ycSpV7t8ojHn27JeNPHmA3XHTXAbyORc9D
pLZgIUnE4R+oYNfrS0Fk8+AlINkmckrTLmLdP6QQAOyMVws0iVa1d0LFiN2NCW7n
if+eq58y+QddII1mwkSmLyPdwNdqircuBpdXChQHNGVhh8pQnqlJNUNrOmJTr0oR
ecO9wdBqq4YbVKfhN6ChTZaMHpFyC7gj13i9AxQ9RImNO5SYKBirW2OUw/ZLIwuH
rTeq7jjuXR/M7yZDKoKQwY8fyjFH/P7ACq0vExMAHMTNpQS2bP6JxeXsKEO1bkHL
ENDik8QJv0lFidEKb83skJQ/DwT5LzskWZlM6dZ79xb3CZ109Y3C26HwAj7lsRsz
cKgimNK832er0xFCnu4QgfhUMCubcJBH+3rIH6Iv349m5NHmgeLBYD1DpjInBSYk
PdPL2KNmUrUbTFfj/g8A/1myLDoFRAGFUQF7pDRiW8lMRCklWpefXEsaPZMGAaUR
Pk5oPHJJpI6tR0bhy8yzIPgb0fZP1yET+iSxpQHoOaE632wdE8+MOOPNm+MPq2QR
MEfD7bE7bAuXWiUypOGNE82DtLuoMcN8KbUj8A3gprszrvdZ2hkmDaxSlyguKFbz
3aB2bxrKTBMPuy0pJBVpW+s/y0VmfFWwhAq8wOCe3YO4ZVjv96hKQHcGiizRm7xy
4yQSAs3LR3PiWm5kfaxDLEdsdZBmIVuMZMykX11podtMabhLX9umGYB9CbZ7kVca
YtNq1l4DQcN7I0Rjs+xna85GOyat5SovLgZTXdFwM9h1D7OCbliQayl18eD4+Vdo
f0YNfYrQhLepeZQg8zraUkAqOKBViswTu0ChbjlhYSwg0TlJgoQ1dJe4ImadZKls
Fhq7TnF1tHPWiQaFn5Y7ElAi1lm+jez8CAyUMdm9WS0GWvuCnH+Qg9/IogzIGw1l
JSNwtgMpJLCm4xi2FNqVVwMQC93DC1eGmSGBJadicDFxtLGjSVJ/qk+lT9lgT9Ke
RHCapCVA6jAVOwCdwEOhpAK7LvT6xgC3KZ9WWRKRuQVlhXEMh5WncHEU95wCTZn6
l4cZ+wwQW5jnKZy6mb/Z4OOFyneNAKWzP08afr+BUVbBORTnMWCsby0ij/uH/qDf
zR0ao1sFS6SRwYzxHjpJSTzS7QTPUVEHTQjvYyzYspoaKLIXyLtSJ4xCQvkLeenK
8k43RlK3pVbuMLfHmYmm75FmWjrRIKAJS+7HTHjxedPqRzmY2KQREfljPSiNG0oD
XuFolra/J8KSSwHtoLNf0LYXOWJ448keRXX2td6MbAthy9WB2WRwvfsDJh+Hm84w
V0wW+ObB+kQ7dlpSQpCriZfKrUD6SBBUlGbL5mvqga7QtYI/qA0xOZvaX9KL6weA
2gfxEavmIio9tJ2lcBte8Ve1xPqPAweQw/hROUDCty+IfLQQ8EVk20ZiI0lPt3yK
MRUGYcsdeIa508Llyp+2zwsCTcS1+E3EgXuY319g8x9eZB7CPlQcTPhVd0dpwrtf
CPxi7P+cUcEeVMfI7e1+HYNSCRE8g8WI8wt+SE/cNYNqeAip9QovbLWEhpTj5csh
sXnij7KjdMvMYgIjxv0dYNrldXvoUoJBKM5IHeAuI0rGWnGskTzRYYo2UDy+8bvh
fpB+s5rVlwWbLdBz5sL/AeaL+9285wkZPn6tTiXjOFW1sLmhoDDI0qSnRgTsWXDl
4h4WkO41JWHNm74Trcv+fhWh+68j8Gzp+T832VzF788XWkFIqnHPSD+VYpvSC8K0
2pBEWu64CN3Zl+2UuffvK46WHX7aXOxaPMUyPy3x9UYtgdQw6epfiuwLcSkaN7zu
hu2OAVm895ai4MZnWKt908MPsWUv21TdsSIVX1eswE2W+P9LzlR4NT12D2UcpRhQ
z4LxfvmGyYIihVHuLnIkMCvZ0okn4Kv5VsHHBxoBFWD+cnD+AhmzFBNQgEbqsM2o
ZNuyiJKBwtklJrpL+sSeI3IaNT0CFFDyj76o2u59NJCerr6BgiZ3m5c1h8BJN59P
iHmdd8y4GybA38uyVV02tRswHf0nhcB6m/8G37jJ5rzliyOeKceCj5dIPt94pib4
sBYQP3XYTe7+Yqs2z9o7LMmwV3h6tjy21tq9aoP6mldFNmBlGWrcRRFdXqLqwLUq
iAiCUXkvmL6edcXsLh6CJSCHuWmjUhCtu20osbWrKo707KEMhrsiRcnT3iAYLPrx
1SOiJs9+p+XYFTDziVmAoWrAhszM5lNaJBQzr/5jh/VF2pF/AXXcXnqvQCk3/9aH
VJ954ajBeMwvTTDSr/N+blGnw3sbLKOiR0k3U1Hw/KIbhK5cBZfPeUQ8slelGjca
7LQ7tlnQJHGvukSn7wIFwXYZblI3EXCFGO0gUgznn9RWyKvFrxOiUxNyseUD/bZB
/Uwur0m3Fqoi1sjKgPyDiiM3EBbPhnuOIwyC2azee6V+dG5dmj61eWEPJ4lWI6sB
bs9lJ4Ykws8TAONbzv5TLWXaCeHbAlFFMgOxVI12u3Qqu24neBwXA1Kgkns/q8kg
ENyq4wYWnXbZBpukhaQ+h7GMOnoGpplMVpyhWsQ4IDSf+vbdPDYNH1FgePbdif5T
ffE0ls8oNT2V3WLAaG8v/3CniOZsh7tNyFZEpUC1b+hfHxwuXhbf24Aerazha5Wr
9M6qhVqmaWVOECAYDmoeC1f3VCLMwFYN9TGm+A/2X8d4Cy5r1vz2fIYdu3PbIt6W
KDPef+XMo6Xd4ZFFxW6reuESEJFajHda7rrRcN7G3+aS1oiG5UTVb9lo4CuewM4J
5fz6ctKSnZs0FdYbvHUaWC5XVddtRqZjnUD3gpOR5nzIUXh96J2Dw08zPlvpXtcM
yqnFNyR/82YJFyyZOCFkRA+Dg/9IXjLTiwFH0pNXWTZbcEv8vj4Vk6FKONBT04eJ
dfQP9hqIzm7oAVTxSt0fJwLSZ2eotVNOvo5GQ8frg9yFuuNlL343bErvHzYa8+Zb
wdg+Ntyov3Ys5W2/G+49vZY0AC6EOYyUVZMQun8z1uslLpT2mOhLGGEp+0KYjxHV
wwG371vwxG64epfyLYfGRnb745YUYy6BBJA0JPdxjDPBgv4Djk4mYnuFIxVdCrzf
Fn/lpzdnTOC6kPuGFovZtmDayWCZvK5RC4+be0jB0YEDlSL+p9ZEb3FQEwJnZm7K
fodXKrg/CxC2GLBDW8aTEQk6j6wO38qz9kxFihxRhITYA3vbLtj+QcWVwL2prlbL
MiVYH4PuJs7TtlANlKJWqLXNvk4mHzBexEj1/0uH7GLjLmbl/+WFVXMCJYWlP2Qi
68wroTJwtAw6JR6yK8oAsA/+5gc73mrPONuxA/aAwJR5oPaty6TI4NTRh7kIN+14
hZg/jTYoLC5oytg+pa9uiVYqQqK2MoG5G30DLSfnxJUEdGvcqQc6jpfiQnbAwTWq
6WWLwvJejImeGH3EM+T18/AkMsVm+zztFcYPPlIMYaL1sEg2G/b7y7KvfpNdpp/J
mGo8r+zTl8UAMi6AQ/6onseUD93DjxfEQw4ewzd6IkbEkoSyNeqQ3kbobW2/pbLc
pG1HqbrufJH/tiXCSnpUsDRYP23MPYbub4KrcvUvAkW8izU3ANJ6qqFV0C/HR7AN
Z8F7KxHF8T9h/EGGqJmWLhjVbTjYpfendPp+qhTEEmh55A13hExwv68/8ejUbiRH
qf0x2xrwvdufmnY8OSXEirIMNOe/k1lnqnh568fKN1k0obkiSjGCGT9/ov++ihXV
SnTqZNyYgjlRRi7X//ILLk4R4VBVyVmQ24vf7AhgmoHClcqjhKEnNtar3LPaecgm
S3HXcFmHb9dSv1TKEXV229bOaxIRaMgFsIPLwijOEc5earMtQkW2Qbq+/CYBzuey
zpQ/hUUHVNSorb20D5JA600tHsy4GmMfu7fZcnV7czD2Sn2m0HuIJIRupcU5UazQ
yB3FrGPX2BhMwKXeQ74xjCQ2i/8GViT2Bv4Rutejfs/mH+mr5jf+isoWsCFBOXjW
uAUPCr4XtZL241PdnSi+KRo5GByjw9zr9j5BJN60cCEeieit/6YnT7ouMxBB8rrs
c9sq4/1U/GlWE4ek7TicHwO0FB4kSS4eyCgLs1e+k2P/TiaasRKbQbu/DGfvvS24
a5StxecfCW5Ox6ws6O1sa2nU81v2ovJBVWpgUYKJlCqzIgJTzDjTbcvLkUMs5apa
NnLO9Ts2V74Tsvo02cCIZMHl+68TTOer7CFy6lE3uky8CS2r3DJiSSCjb/pB89+y
SiCLmukVSRbrvMbN//L37rTzyOiGQ15/tWMQ+scvn5/yfOAiuQ5Q1mghIcmaMubG
xjdjZsSA+7Do72PWj7EKFhBGVje1QfVpekga1BdHtpssrhSXNVUpaOH1hwJCrrtl
jMQBDcns1JP8GUHSX5Jp4GXviqXpkq18UgmqY2xvp6NS6iWENTy/rbhheqd+PHa5
G3H7y40sTR1HltH7DgVpW9cif0AvQdd1u83jC39SefVpBA4FcSd4tC2Y7smbkA8v
t34KN8ojna+OC5a+C8znOilYyO1O7n2BWtvfvMxSQLxg9NhR24GEJifkBjUP51b4
96dyR0coZQT9F6ZDDOx6jVqW3jOyQVHSfQdOyamdPsrDauVQkDltMUstdc6/kW1b
/fnGmnsDZNCZrL87aArQx1fr05ZVQYVAgxpJ+UKt2GdoMS4SMAu0ZYbPpdomKmb9
ZK0x+u962BjEmQe4DknysABWVSRu7hukOB0rcQNEb9BxlzYE0JLxRKDAd6Mplhbg
8wUqWz/dzVSVJ/nnVQPotjFl9+mUTNQaGDsSzsex/xgCkv5rQLcZ5BDObZ7gk0IJ
NoAz0SymoeDvmf+ZzMQV3V0abjIqu1Prn0AO5buFR0vaM+1v9ajd8N75ftjCevDM
k26n52J+JZI2uB1qOqhfswQvOANXz8hqull9tgFNBnencadK/oOc5kQT40z+4Zp8
vMHzRXsPhwdg30WaegQMc9YtLjRVUux46nBf5Va9gaek0Y39Ay0mYso3wAEkNeYY
VxoKDBcDobO83M0L8zC24Nqs8t25jcmUeTUVWjpW4NwTdD5HOQzFnDfn8YqfHkjy
7ZwSk0QrlXn0ZR5dkSdW873buWxnS20yhsoQvjxlS9vqWY6pQ8NuFUkfFwkQCgfm
JFR4epDI6//SQV2RCAbG7uygWFifxE0VxuwJ9dpMSAE+dVewQub3lJYHLlQSFusP
w59oO9DrArOJGiIAB7psZjEl7sEbSNV9DYW5COcJNtSDR1MjxrSwAcrOEItBpt0w
1CuxZ5fAWnK7HKgpfr1FyNTbRtXBWU0Loa6hjc/k1YGPKgJgtFrrM3c7KhDP19I0
T3Cs2huPjJ1DnRo0zjqEpCRQA0nEQC6I/6qe+n41AO63xN77bbc6TjW/IYj2iKDF
caSQNNpqTmfFbNE+6VoBRTu22BcGuRVEtxibvXMrbAzqqZfpT1sBk+3q7zPxnIXz
MjQ1hv0ep7yLt6gzB9OcXw6VFkyY4e6vTTyfI2ccu1bqRJygDcLiUzmTFdH6k1/S
5EPSrR2sflLpk6ISpu0nxJ9cTG+962hEPG6Gfm17FS3Bic72DUgtGxMPJiR710QU
HhHn9z3wpTYYYk22kVoKjbN5dgn1c2u2jlmRF7MSFlauCDl17q8JMOgNMWrvCGsn
CkkwkKOVChn/FQ7Nk9iGIl/oYiE47x+LO+iQmGkAMoJvcMse1GUARAtLQdDu38ot
e6c8Ci7JSpkR6yz1o/XVVIL7IGXuHdRT1Mmt+HFegZ91cIQF85m+9Wqt2qq8680F
NF9HbnGODPSp+OoRL5LfQgnqWqIJSo4huHuK+m5DYuQvIIEMnUkt2gM1L6Qf4DS1
Q4Uzw1bUu0r4D4TpJRjMvYvR8F1q+vcW/HANEgmhZuI8sQHG5nzJzY9t6usPpjms
6ZpP60d6yQtLa5t2hQUMNUR+xLrRMxrKnDxRzc2Fg1dEPV6RW9FjqYqYumY1enP3
cxNoKvf8u/TA8axjQEJUBWKqmGAooLMIdoQWuuAtU5slVo0fAZ1WOsc9/DT9OWGE
QyCFn62Rx4jD25h6pCzlel+kEvbYeFN+8nfDK7z4m7AIrb3QENLk/UHX/3tioe4i
PkkWX/8wr+rSRa2re/OMTC5mFg7VSUBQUspmRjJ5A/8BWyHObabRuyCCRgOmqN/3
sDr+xzH2hEqI1osqIXHbV8bKU1k4iVcSG6RWtZ6Q9Gb0mtUmp1ALoq1jPVqiuXjH
0ZJZpLrKOLUSICn7nBu5nbvI7krVuHflVc3IQgfLOb2w1BCAV6l5OHG4xZ9bMjZ2
D81DkhwSGgShtgdpn5SsdwcZ5EPqVMD7RLl5YTvgH+Vb2VAaKE2MBrhX1SqShn9G
B2x2gekbUkP7tFAv20cj9FKgPOga2t3cXVOfNtr7X/pgZij6C4kFx2H+l83bGk13
jKgS8P+xxTfvt6actNb3OVDpPMRMOqfqaErqlnCvYhTkSffm4Vun97CWuncHnHjQ
U49A6dOTWmJwWVXi2hmUiBRs3qpKLokjIVXbJ6A7d5/pw1TXXrJK2v8Q6wmxhG6D
yS0AAH3kxTXMQ/QgwJ1O55+CorDsqQ2v7h3NYE+lYe4Oxi5Dqp4WD3Eege7rTd8j
X44JV7r2NJJts2m+8XSMiooWeHuxqQUUKSopLyi8fCu77X88eWZ4ZTjjsZ/l61qJ
+EbjLFBjluXg9e59Xkp2FP1lIFV3kxJGREczJ5sBSpqIuBmmuuW+REapW0U5Nlt9
dgjPTtLqltP66+avlaps9gA5D6zlWHASj6xfa8V1QeFVZPqUS6W4yoQyTik9VXUB
RDw5hS0Y10b129lPu8f2iwIt3Twk7cVdqRwEiT8FjTq+T6oUlmj13s6GSom8VQPP
6XpKHE7PW0TQQv+0poo6KDCpTrZtj1DtDGnDVMxTSJfFTRt8+9bdzJNbqSu8rzEY
C0TA5uLLJLtr/vodYNsnr1tEgVfYjsDJqO6yldkyYwzbkfdc1ZsXTfiWUR0+xkCK
q1FYS8lVInjHxeM1/i0tVBBA1ZmnM4levdIp5xXOPyk77imbyjEseDF1/Obiabeb
ZOfFt2Vv5yJ0eHhwEyJ8r6HuafNB5DqbCdHJ0kDKrmV1ZuAQnOj3XQLpOBdOCyyC
9ijaHnQN0A1FTCa/S2e+o9UhXLEGjLok+KsUYAcTVXh7nX9sEV8f17w/9/Uu8hNT
e4QDMuoSQvsgdd1WhjqCBOu7KYcgqt8HYWPQeMdxzBNREoy7x8k/fv/aLLR3IG0f
cFhFKlcTYWESVALkfbTIVh3BibthK1+uLGUmGhx1nKAt5bcZ5xr88eIugKVAYde4
sWziDAQKdeuTvgWVI3YZPSaY5IHWrWpdi04NPfLhsLtRaT2yLr0CdFsjnmgan2iK
hvFkJv8ovPJewasF9zmNNwDkengTM3KxTMIDnM5aPYgk4Sc3HeFgP3t0iA03pU2B
ytNJk9tUCQNnX0X51qX/g7t7V3nwuGCsCBzgQLRBHRVTdWol1glsJ4L4tZfQ0+aw
RCChD0kTwzXRQeulGnc8WssMB5DeeMtxDmmoemKv/2eDnb0UzhidWjM7rRPEpmUi
EMbOKiQyq5XtPX+dQAXih1H6+MdoxKOQhcqFAW3c2A0gih2BKbhJCdiTM8GXdpxe
TklJNNE3w6Gngka8vJrwvRdLpVbaPXZ2cem34CG+w+fmgq8T9fJlYAMwtFZcWqPp
/53Y9Q1CvPnnkprHgBurCoMhNY7YtJocUtlUaq/G2ZcI+YHXPh+iEL0mGNWUOcVJ
IcSkNkuIpSe/rtJHtyCBoPHwM2iObQf7iHxmkUN+Evk+/CU0HnfZVyoy2gix2fYD
+jW0LCtGpsoQhp4Xs1GlipfQD9jd2WUeOzsyBIpEXqsr1bHidRGYYB6nvLxZVkp1
NJVdqTlvT3y8h6zEkFANJM9knLmCl8T7EdBTgt7VTMYdPoy3KwwJ2/sc5kqXd7E5
zB8cMr79JCLagJumbPL0eVA6pWWKRQ25PzjhnkYwLlQZG7j0LrS+KuEajn9S8gPt
Uxr/1smnrwfDtsoJ9ZmJ4rTOA+Stajgb+OJlqClJE8yhr+3VJhHe+aqa1G9+V7IT
fEetIneGCnervHvv0PJKVrCmdKBrkPAxmi5w8d2O6sST5M18wfznjFLhzAm7hPpM
S2HMmTBDiBX6XBvSRQDDLx55KLLSrY1X5DqNWx8C2ynY+ZzKa3JnaF5RXWfTIK5I
MO/Xz58pxgopf+FDkc8zleoXNL4SIFRJg+3FctSixCINbH4shpANaUax5XyeqjJP
A7hNDRZYGnyGLIG1dSHncMSDql2JSzu6NDkb/P+e2DoXqbEAFVIUoWJyjexuvbjC
NJpnfabAFh28CwiIREwxDo9qzQofyLImU1ZcPk0IZTrnNsnTtyrYWPqpjlmGgD3g
DceN9fvgVheDBlRDYW2Wn+p9TOKf1N5X+JrI5KO1CMl06sX1xKoHfK2bHKERFg1y
W1S1bb0oRWEdjlrx/NLL5QwFxx+SgMTpK8vITmmOS16BkB1hoMSfSJO16SWm4Lyj
mjviknQyl23VU2ohd3nxRzXXjM+EfaO4s/yHCuSfCm/wk9MnM4wZ2KJzZ40UtkSi
71cvPoQS9AOppeDvJyScLNp4bAORCFw89nuwHn4jK77vLjD7m/foFaQGTx5sFHK3
HjQFer/K9ptCPY4J5FYdtYGerp1K6n5tvfdUWPCPwIxGkbOiYGnhpaTq3nPezUET
6it2y4s7nTd1cbMAXIdaafVCP8oQKOHBKUVn3lkUJAXQpCLsGjVJ9JB9pSI+JumZ
HqjDQh1xETpSnXd7Cff5JpV0grNJiFQVeVkzNf8S/W5Jf69wzhwRZLo9T58XXefp
1Q85GRyKJVtUmnVOTYHl3WAd3lXtzjYKh6Zi3qiszAXuLCyp93bef/m5nkFFG/UU
Af12vcYE9QQZoqd65CB2iN+oDRMwLzQLOAsV4U7iidn7R+OPg8Hg4EIyOBEYq0MG
6tiZUlhSEvUxCO/Hvwg9HDlMXPXeKssaYhBSNz8xVlZcTEbIZBSpXNAunvaatpt3
ThymVkbnjmGOPycjNF2yV1nNvzxqoMPqnJgePF+ay/I97j5bL4D7fcTN1mZNKtPJ
v9Gna4a0hxcR/pA1te2Vz0hziqemd/i8vqBq/EDXzOdTejewvBnQtHJnYK8q8DhB
4+0RflQESiCK48LsQHjqRCFtdyWhZIg1XgFqn3TFEm7B5ITKN2FC2UpCVBdfCiWQ
eeu7yJ8GNzo9yfoO4plrcsevFoNe9UN41m3xYSir/HKiY2+D0dE+x00irZnNikLa
nmE42G7MidpPzeTfMHi5ilpQyXedl4hXZhFrSB09W+3LHALwJP8vMKddEzGEw6+I
l6H4UwwJ02APWMupk/DSMyMFZZhP1iB/xxs3JS1scCcD5gRSnBFGMFlEfOM0+EQM
YzotWhcFOzWqz7OtmrBm2N/YlU1tQsX3gZg92P6Vr2l7hBY8NPC4jEhiAtEBhtV2
uJGmO7aJH7eG0b6v/tiKCHRphMAxqMrBZmuyPG2SdHZQOEI4UPWoFWAmGTG2nYtx
qk5H9Q7a3AhwRAqy/bdB9wYnJU46I2ZfcYYVv/wVi8aNAFykiX589sonqlGdeHFO
hEQKxxgmabPSSuYXk+xXPTf0FCgY7QMzIMREnq2fci3YVt+q2qbhlUC7STAlLoqd
GkDY7BnSqweN8I50QniOxk3JWfduCMLp7Dc93Bl1zF/QdSEk2qPZtfmwKR0clGCo
asTJBq8JF2r1OPCSrLK8OL+0mmEZ5LFydH7gS068O4fsPd5Xtk+NelmWHmaKQkji
iU8DSA6rAmisgFyHUWBtBvO6r8r0vp3wKirz1vZ5UXyKRsExPFpAVVBUTpd6zas1
VFURhpxVgCHVP59uksXvcxYoAatr0drNJ6UkingstmhwhwYTcm2xv/uOj6XNj+IJ
CMp0lkp4E/tKy/czv63ukQ7/imMq3s5VgPVDKUCu3E9z6cX7RdbCnLPiQUZ7noMt
OSXDcH6MiDGJugbkJnytBz6yh1ZdMuB3hwOrt+zV2zLkFr94STqkWGg6ufEBHsp5
ReIXB0EJHwj2ZipLcrar2bVQFVJadsm8n/zzdHX+9iZ3SIxyW7h/YF1zC1tY9KJT
CYss2cysXGUm14imbadt3SbdA2cYGXRETa538zWcI1SGm5Vpda6Vzr0niLAYw6eX
TUYmZEQVxoFf2VSU7sWRilmpNjlphuU+h2y547AI2P6l7wBFj49MxN3f03BO5guD
FJFZxwK4L4LcGDCGNNhEgxl7IEaHx3sPx4uQwVzGN5vD+5/e7l/FAtXIFUQsFzvF
EZ9atAchuj5/gvA+gwHPqROkCDsUpEn4AjP90cPGMxTnPz8NVlbanKZliA82oxoq
EFWGTFzUejxzO2Y2aCmTGUTETQICWJfpC4xHbUXnghrD6devDnuI4RodNRxymCAa
TDIVR15kFbH0Cp4AN9zq2mRCQd4JWC1GmsXXtEsXUA1RavcLHE4jv22SOU/Uekv4
yMzHsenkil3oWxbbRYlFEdq138ItMnedP/y+QFB2rugRTEFvau+BhxcftxVdnoxn
+IHKUfSkoAGdRNTTdBnXIY8wmfUmDFO9hxuy8y5hoK/0arAohGzi66r1HDpLdc9v
eb0YhT8fldopa5snCbr5InhxM1FR1z+G/Aih0WwMPcQPyPUIfELCTs/6CPZgSuFu
Mfkd8eW6+wY4XQ7VLYleYJebJmmy8A3XsKavU412/H++1cG74KrA5h5NVA3uakkn
eLPH2214CYIsn51bvO3ljYfGwZtSx7U5r9aNyamCECLm5lbC9Ie0hZAOWfsIISIo
6+N5Iok8BTcqaXvMwBXocDuIfxPwukIY6GmFJnv344fLemZehC35zOd214x2l/Gz
IW+SZr38tHhCsFdveWKDCSalWEOAwYphpU0V97IxRdf2ChOaiZxpDgau2Mb3x0U2
No0T2ZqaJfo0HzhrpXFPAgUdW0R8O+QYNBig3ZR30cYsMl8QCXb+zTUyI4DTWlyv
eB2FkYOoXWqkFfSiin1Y9ApjWHhGpCLVI+MaOiiN5WfTC2Jw1rNOZmfR+9CpLOM6
3MdOqGNeJ+mhmEVN7yP0MUjtCkcqOnvZXODe3y8x530F4hoH2BhEqUu2g8DjX2cc
L9uKlKdbXea1v8LweGDPStRxV9sKWBuhmn5rHyoUzwRR8GrFXXdoFLPXrNQ03qfs
F7UlIOlKFoe4XFocZjkRswkf6Bw5nG31nw8y/N0ORVwb7GQVJEeHAfFca0xC6bC4
6pqPKvkl5FbZbDbEkk0RnNJFw8VZ5cDP+eNekpTTBVVoIxBJnoE18bGe6uDX/tsU
/n7o3CywfaIUakm4bU55HUCp3HkEn4pYBgbYls3k1mJTsvV1m1OONZCeESmtjgeM
ejZdAkvy+3eiT+P2C/JQLTOtdOX7UNbO265Xm39r2ABfHY9FDBsqCGIxgw/mPBD3
pBvBlcO7tZCYKlZZoWpXoiT7N8lxCMdLCcFqwSvczrloy6aWNzZCo0VGT/SEvO+k
gxs+xSssi7+6HPze9za3dvTxnLKVXU2mkxXJh1VOHHB4qb8ODl9kkD4zWUJ0Porr
BVnBOmYw13djzABPa4/9PUZ+E6cJHE1+TiBUtXZTwD/efIEXhjIhkP0Om6S4A9UN
fp4Mkjh5LgZ4fdddpdAIOfdEgv6aESqAQE9BvYFotG3HHwjmtNX9DZkYUgKFCt2z
/oZP2+tBxU2mNBlH28KYjPrYESyc/A7eS7Ia5aSf97iizTF0ZcByIkexBVNL/is/
gZxOC83QYzMjoNSiZbIFd0jPAQPCTyOnAFaeLqEupWDg4vFISw7JBkVsLludw41X
Hg5XVO/pw1oqtg9wJ//RHtoHqxGI51uo+JGznnWTH03g0HaQ5/yIg2C8o4YBXuy2
RdUaYmnPAtu+dxFIAD9c1VvFairAiuIJiD99PY3FQqzmboiuxjyh+pHr7ZfNMyUG
Q2bQuvw400S9E4cTq7nozslMaAhO4IBqY7Qk+5zOYSI90oBdydv5xcxaiEHA2Zas
w1S6XCyAVr0TQgiGev5GpaTbDlYdey7/0oQO6LyZGDmPAqjRTLWw3kWuBFWqNd2U
bx+1ZHgoBG0lX9mCSKN0Pzre8W8T3prAvzyKbkksuNB0uFMNvQT196N6JoliUYOM
/DIoMfKrwjYxXVVCugLHZ+Sc2dMuScSX0bgG0fcr1nclWY1AUiZx4oOlI8+t1TuJ
WnqyricUufykEen+o+hfyjqta7B+k3qdUR9jXYqhtT9oO+BfV/oVSzxioO+eP9bN
liBodP0Tp7wOKOIkCt/5XEKgGSFmI3ZK/x1XSkBwo5cy00qAPU2Vz5Y8F0f4jOfy
WUC76crIPamhLaVwwJGS46xflfY8P8x0i4Np5n4t4qNVpq+UjEEM+H3Z4cORVgTt
g9blGwu4g65c4ZDNHUnq+jkQLhwyn8jn4t37TQxfv9vKCRb8pngjHiK6VgH7Jmps
umZUQ0dZKYqv1G6Qxo3Xqun5P2Mi9XEeC6RXZSEe6QQIi2nY4Bq0KM5nzSoWzbdE
h7BF5Np7+f0/ZnEGQq/jRUAewMLDEjHa9T/1gln8fZm/H6MjvumowaLd5m3Cv/As
qy9OfoExaHTBGawj/g6eD2YjZ0zMEu/djJofITXLEWCPK8H48vm9KSlDAVoI4sOh
g2zaVPwTGpsbt+uYMUwY+wGhSr6acZ6GaBGaCjqgQn+WnoX2EMzvPOlZAZz0uiYV
G7MpRdu23NsaoEZWdRDKqqb3O6bBJz90+DO7wxzMt4dhOxAHH4T1viPvW3xliHJI
icUYj5m0fP0ZXyjiBLQtXmbWqqOweMqtDy+K9PwrAesT803Kk/lacgXLxjTYrBuK
fz5FyxPVggQcG08bMUdFKkEs7itGmNhjbf3mF90E8rOQsBSAXPNzoUkbiaTls0L2
5GDQRhG1NYnKJbBI7XqltoSUd0Cct3c0cdR1Jhz7Uk4ruoRTfR8BZGX21vqHm4QJ
02wlsgkuW2q8aLS6b7T6vhZlpNiDM4UVQIdPm0JEDIp4BDyfbEzQjH/Qn04nQaWO
h99uuBzTdM+/1TYcSbcSSORmHaur6fbHLVjpLPbHVl/9R2J0PreIXa5rH87V34uL
Tjl2/hJb3LZvHZTl/NyACmMNi36MVK4bTqcdRE4AsehbDPgKQHUedYAPW2N7mMYg
ZOi7Rzv+qQTBapwAi4VhxQTZ2PQGEjW0FVfAGRCXei0NAb+0j0kcXW+BubUPKFdT
oMWzkMvbeDIzKyn1FvEtD4yxv9oAZfyImmIbxP0lhFuRxnxf6/MNtcuig+LOM7u4
6NLqpdiT18/xkoixdU417WBaMoiznapbSf8tBaLqV6fhfMvqrIWbpIPfDGCuKtPo
L12IQvLGnxIqmYjf4kBo/2tEpY20ilF3mSGmJtTZ6adXwnn8YwAHqaVFnXn7uSFC
WfZKijPj16aDaAbnu7cNUdFOXrQhG3ZsyTy9nvAjGfb+KFZ20urigzygQoOvwymt
kfA8C9kUJssvwV0bvNJS7lh6lGixdpHo03xX5elDCYsitIbdE9OBVxBKOnGuzE9i
qaQeAsXBKnLdcqXBsBkHlsHmU0ELJMBXGjakiGmLaCpOC7cRIw9/PWRQF91K1ANb
R+kjZrYhT7SwG63uOQHV/59J/z63czrJttVrOWxsUD3lB8pW9GyHPkRbpogsL4l4
I8Xdpm7AJ+ULpYGw0BOq4QAzBLVq7XL8IWiUI+jzOwxs8SzHa4Kdk9Y0bL/r3HyK
iv9SPMuzMmKuj99CBOhXxuAmQ4U0SLRLOoboONbhV4rr3syaOKf2D7SwJLFoKmdq
dx/HmqQkczzjTaNcoBvc8VATzRqQS2PvBSMJau+ncUHQ1V3qWZMtReBXHNXizsom
iinXQTHektKnIICDSSEkLf+wdHcxyx83P8j3Y/2jSkG+Z2mSH65wc4RJFKxacKT1
1Q2covF9krLfodYZHO1WWFMxi4kRVaWMmyHRAJoYo1Gg82lO4isbi3ZM301LI6/g
tOA8YRUKHu33WZ9Z42SAJXawnkogJomgwkiIQr28QnHMME8Nf02rlw+bmgzlsrDe
GDUA+XhZ6gh6HvTAGVc+UJBnSGFAwDzfL321LXvh5Y7UvtcLjEqKt/TiWYC4RMNd
EY5VjJJi9FFdG07lhn/OR752InnH9X1T69Ogma0vHMKLyaXO2cOh4J2m8xxsZ+/G
ed0BDCu9Z85hDEqgQBOMJDIQhlQZ/qTDNF9xNPrxBfDHVmXqmyH5yxW3TJ4LZkG9
ATpJyMpgwx4iKkQDrN2CDTlpwIbmoajXxDUS/bR8/U3f/qtmEG4RxZObmxNT6oMi
wFHVV48TZnIZfoiIs4JOSFosKOIZzjE1/98ClDgILSj/jgdrkalf0BRdP62yA64J
wp26pS1M5f1zY8OKjgkFJ6pLujzMIF/0Og4taddGd4jLNkkRJqq+YdmhIbJ0nYgs
+GDqfwdoxOZjehNQgKyggRWGebS5IbO4hEIEUzeI+QMmEtZpap0Pe7zg1aYkx4vr
E59v3ThfXqSNwtZe6eU4WKCLPCowoiEiCj9nEfaYSHY3iCvXFyAfTtLZooJNn04w
w4lnw6ieJIDOwfHCJcMO8zpdGDtgSCPLbKFlXOawyN2GKZT1YqkkeGvrAgUBQLcO
FSpCGPddsBHyRsnBk/43tTCmTA76uhLIJnVH90Z9bPBqThB6Y1JoUyVXn03ERS4S
I/HAyOxb3bhG1FwbMwglGjozY6mAauHVbzI3xPG90EZlXzA37V1vy+rMwP9MVzby
Ec6KAojH2Reb3HAOTKPzv+TN/uoNe7oksyI94khwtdkuIHiqOSziG0iNjhVwj8RV
CKZ3anVx0ip6HOf9K/ceFMEVEGdO9bbZySO6K4CeaiGTacyOWyG6DaKIxQAmbQAL
c8mRY9/s+EcC8nW+cZ+uk6qNav90ySAR88YvJBEDYl9C510j7n5RYrFojDnqCVYF
niREXivkqH5wIr+HIZKo/b5NrlX244N2FA5YIVMnWwY5O7JO43w7ivHxXazMa3U9
ajLg8T+MTWr2f6hwJSzmc3FaoLZ5C4VPVl5wrDyFEJa2qeIul/LWi4b2YO89Sder
7M9BsKI3ylsctfki+epjsz/U+CSlcsfS5YCcBxza+/k26FJfb3hcHKTuOxS6tWmH
IUzXWZESBfkm5r7CEw+720YZCI0vn31ozy8Xa2PTyLwE+Qq/x/qpIobEq2PDgi8I
o7IgvJcFu+SmbRnKXjmUpkwWN8HNhqnS7cjThGffg4l7UUwIrar4ORshG0NzdTog
wijn5luwlII2Qj4UalVuCLtTJsO7j/P6x5PL/FqFIK659UNKu0PzefSt1B7iaeVe
VZMgdXowiCMcYjQ7gGU0AEf1bh3szAOwAjbcjf6WaCZQiJGjEm/TSC0LVBVhGepH
M7HI8/ID9VSBg34lVAa5W/3J0osWq+2nrNFSaDMIMg8qzn8a7dsR7ELajgPS40J0
xoPzMURQW7CjDHtD8gIitrD69VWOCyxJ8KvkdbZhV6yncJ1SllPoX3sqZGUVAhHj
BEyiHPch3U38wHSIPeHBHh2o0tnRCty+7X+/M+MApKHZ19td+neNbDgRWkFBmPm9
sXFxlZTvU+DuycKXlrZNuLL+8mtyRN0iYfwLu/r8wzcdaC3Mi8pWkr3hRTX53Rwk
1jx9P5mgcvuP8wYRj51Tp9/IpwyYHHA4P3c9DKKvMmeqEDmluAHmjqBcgQSPbTsg
GOevy46jvonAXBL7BaU7+nbBc/HvV/65F4j8uCvIeHKLyKAZvsj4u5yqHUXJV9SF
7UystUtIWyFEbhqRXVFGQXPvfbd90kRxEsE88WAE6EuJD46SwmuLhvVr/SmYwPyD
vkp84ltRQW1fTzprwawbSkrvWhpKqd9NLNxOnpvdllXwswOnayLosFzCABAcmNUr
7y3lGYYAWVqGtmJ+db8w+UpIVw+osOII9+TN6y0GBihKD2OMdNeaNSU/sF2ODVHD
ZQDejjgSZIRHeiXA3BH7L01r6ketCBaromE5LtAxly7uCA4Whdu/joFHTIzOXfQJ
rxtlpMYeMGEHdDlV/DulGpplMgtAMcIv1OhP7H6yEVEEtm91dhRpBP4bjOQHQYQ4
BpYJV69Jl0rtNVs/b8XZBQPxH7xRlnvFvfAr1bYU371qlq/3TjPTYn7JhWQhQjrf
DnOuPz5jCsBCoATt/qZSnyznutMFG1LUofNb8NLZG27UGM2IjZiOquS5/113EWST
Oqwhz0c/2EhXh/JaowbMuOHY9AjnKhknsgnRZx8ffGtyrUcRCUWvgsKBEcs8Bzr+
hg1y28mSJu8lqeITGQGHOZyCv/HNBYIUyKtSwR7sSegtEia4UcGpkKsFA2ZeS/fe
8TeQb++N3M2f9dXomAHrAVGKBiROtW2fDA9zSPh4RLkc40EedYS+2tRdJeDGYrWi
h1d+ee+iPdzbI2MUrtF/r35E8TANwEEQNoYSvtBOxjF4/IQWqXaomhR1JYDMZ9KH
HyMQZ5a5e8S2zW9DObMUPINaCugLni1vcm2MDRY0TiSUqDCAHpIWE7DAO2fXc+1+
/yQEC1n31dIHZuEVp8uNGSTmtSdLPwDeqOW/zUNu5jsJd0CDbJecovKGnPfNWLC3
5n4WGhEDdqvoHUU4/V337+OFmWioYruWPt6cYpdq5j1rJgQsHpPYgOP7j04yRBo9
1AUX515TjuYVoRISZ+NLlofGgczXeqanTIVgfpojFWdyfXTvGTvVUQJGTO1yksBm
l5kxYLJmZ8rY+piEPioW+Wgm/svPgk7MEeodDEQAo3K+hOM2znEvLhe9dmGKqiTW
MDH9JYPmx4jDNnBePWBfsom9jNsttZgNi5TpsY4Z8leowoRqRBrqPq8U8iPbX9rT
iVH5yJ4CUkYxhH475IZypJQW0OisgLdlDg9AFFmYkT2eT1xMjPOBhpCFMwAX5iYi
3OYQFUaQKr7JOR/wUXVIUe8NahvP6AWE/NeWfSbp8o2csKf6yiPnz525TWLwQv3W
iViuAEsid04QMGFmp4dwVlK0SjLBVPJ6YZZE09Hlo79Xl824SFj8Bofri+JFqPyd
mOxNXHYgqoHgTJNHth5RhEmaMxsHkPmg0F87Gq5biMD2BPkLijTeJUvfThTrrbU7
kp9E3shzDn6LzsYMyfydh72Df1cTUAGPfzRwAUamijgPaTpCcHNfFt6+hPAH0khO
euC0k7AoZxcDsYepTrALdsAVLuU1Mgyz7wqP9KbL+D3GWqOkAunJMDg1VkbVBS2l
zv2aa6+EpNcQZFlKRneQmOOuD6A7u7kacLIASDebBYTGH5jzab8Hn4HDBATaGAbE
bWtzAlCl617XGfnBreTs316oMdT6ivuRfMtSkJbpAzD1M2Tr9XhhUj5DTYbt5bVA
/CM1f8TUQTmEZY0BnVzInejLkzfCzK9My2IZn8STc4PVAQi38EfQQwoV3ciPflox
D1JKLUcVuwAJD24G0Qw51jqaMmxEgebXsi4TJejS/PS0NadhCOCqq/wpsc+ue17s
Or36rqzZEqjprqbUWmjkbGLjX9fUhPQP3c10T5SBDxxt1NtXOEWH46gT8xjjPZyL
+pNZFH01DcTp3Y+o+Il7UQbJKq4jtJ5aQ2RVAJwY4WleTri7kEYl2P0kwETtCZdt
3b3z+iO94XlrrBAUhxqi2Cd49y4tGsAPOA4wU7WrlK6qCO9fD+72VKY3/rqQcAiP
NnkU4UAg9OIIcEgVtOjz7BDyHCHqth3/JshBmbI9P/kBh0xe15nXn75cmOgPovN0
U+cR97aCL+zStGD5v31O3+/NE14k+EOMt5fa+HfXjfK6Rbd2KsR71v71Qj6MIf7E
axcG7NciisFiNgeYtNY6SlXf0FDh/x+8s9xe9Oe8gK2osG3r2fI3Gu67OHMCM0WQ
VRkWTGs3ZeZ3yln4nWehZZ9rrWG0f41r4hMicuen4oeEdk2s5vjUF9xTPxImN0d2
jHvXZ4+zsuWLsIyIxHbJ9KYS/XUZLqZR5GXosv/e/sPjUf+cRME8/6/bzTiN+zLW
tiQcj4idJRRMSvVtAE/Wq2tFKculpS+XdVck3PDkkAAdE4GWlcK+n75RLrl5N2sJ
5K1ObYq2fnYOcjliHjtMB7q0cDyUgnXmkcE5wyOPtcfwTNf9BPVQ9rUFIfsM70Uc
qx2sOoNbzRt8i8PvdXo+BYz9ly7K+c+b78ge2L9Q7wnlbE26X6opGKIxmuWmekMW
hdi+lkcnuGbIVriUknVVEmriTXwB7Js/K2OdNgN/kTT3jyS7xBclL/1iFI9RRAZQ
fS5ShKcwmrHeITphtfCtmSfukJqR1jBlZgGWVchW0lAQ1ILET7mqdEgEaVItgMyz
BiPtRp86TmxsJ0wuGBX7/G+qDmz4tAQ0x3R+DB0sbULEiVSSl+JHgJMqoekO998P
SRzDmSLV1KCPIrcIuvb/IwhtUwSDWvgHMj2nOm3FnX6l+x+Dmxs0Jje8NYsPEM4I
NIsDB+BlextEYU2BEBg0aGEjZMJ6cQSE5aYWDzReROOQeKgw7vXefWkQtKV/HBp2
cw3OnTOyIFHv+zS7f0mW7otJVdddJCf5tWGQMH6Gw4hyDcCZbZKCgUJsL0SL9A9O
NnOBWrII4tmlvulAhGDOiLURlLTNzMOgwGAf9rqluyNW1rwPVi50av4fD0uHz+74
xx76PNjXOf1768JBt44wQD8BLFNzGxpvFYzqFOTanNlTIYtPCnDcHLC9Za3hnBC3
5ehOX3ta8Y8NKjUw9+zJRyUNZ5I3ST+JoSUBrUoh34j8Is2KLUAQEKk/k/1dGbAW
EODz/kIZg1hnx6ymBpLip23wvtftyB1CjXB8kKwkPfO3KWK158YURgSJL0/A0Qb6
Fvl/trLdvhC1aCGvIiZus+uOZQIlhrwVlcT6CD3wNl0D8z1W1GLALqsdgnGybyNQ
o1WC+zvSawrIMxGDnAbuEAMMLvKahU2a//qvLggYk5c6GbGwKqiXrWRK4FKkZiqw
ULrW2rMCEqC6RHuv8yW+w/r1Sh1937mezAZZ4m5tHewMfJOnGyz1seoex9ZHUE/8
RwXQd+jjdNFpuS0rpDL0X+ob8Vw2SsT1QF/pZi3OCz9G/U2frzpJX+8RdK0O5KB+
q5jXwAg06RlBREopd4dZCMhrcd5JMXrfxG/spKclYYx3HVmPVOJ9mKJrX8IzyGdY
FphHkQDXpQYOdCCRz3heJ9EUG/IYpGjF7oz1ELf8WYAU0p0Jjn0BqhIS98L2qwu4
xKyarBklQGlWLR5m9ey2HE1//eN/hjX/XtYd3iXSVQqhVAXdQtafPJXszHuWIre4
p5G5nJ+1Ch+0ve5jh3dN/rvRmvErfIKphSND/XcoU7gpAT9RaMJ+ycBzrba/vEZ7
IfTYuZA4pAdAEtO7+bby8SYZmzqu9LFrndob8yrqHSsMCc2ie3bAO70K3THCPHdj
ObtJuGAsa9k/eJXRrZsZeKAc13tE/fSIZARWxF5D54MlbIJZkMdnklxuS37BWgzW
PCm7EgaV0ul4bWedBcAY5EgXZojqFrVdAMzJJxelmDWBwIVlPxvssMW0o+2EuqUk
9WrQxpahxKkrkTxBRipouYBfCxmRIWxIsE0HIC7l5ykQN58bbNMj41zJH4YMRiNu
JHV5rK77PRs8fSJCZK46Yu4M+hMwFrbSeA9n8vSXd+NeWVuvTSeDc9DeB7sRA7Ob
144IBGx0HKgMJhHW2fNqS0jPzzG3DnkQFKx0twLfuo55ovelVJzh5fIY0bbTmEbB
OiWISBgc/1zmSGqDMn/FC91dTXMS3Ge9jcRrSrLEYODYUThja5Db92kjDIWu8Y52
+F1zehuH+ZeL2ZwfupHjctgrlVMasGz1ljMdIGgxKVGk6PJ3XidQxhAO6npQu6P4
GW01Cvpg5O4YLnVt27xKRe5r/FguDEN6aQRRGo2Wq2mBYW84bAqQCp/uCTHqsqIJ
w4WXXs+cBj+Jv2H9i5yn02OQzQMLSPAOh+CCyOvOvEJCeYz4AEt8IYoJgq09e6Pa
Z1ThHQcuBHQZZKXqLVrBhcjkTH+iz6tu69oyaib3C7FDW+pKYQcYRNBaNggBRwHn
0uZiFpmzt2nejiSIV1dZTQQyznZX+PzGAnaP0lXglEmANRsozTc+PULsiSqwkEcL
lPtoS7ZPfevT+HR5mL0R9/LiA2JygxHeAL8g0eJjhiZkBW5Afoi86bpL76a+DsQU
AQlWbVPSc1tcPu22s5yyvTX5XiPg+UEhCjedOBboPSZsbLOBsY85t3OWdLSWuG3I
Fjhhr9B9CSZxq+5BfeQ4G08FMyyhsLZH4aQJC9h2+28+epH15F2X2xaAktcpYAaG
QFFVeQs0sk71T4N6zovALgoDr3ZeyWzHYdTqiadr1AjbCLhbfSGh7y7p1QUeZOiZ
gIGGHCcaGF5gRHwZnYwUBCEjB14UQM58brfQu22R3TJpmIoadceC2T74iUte5wMz
dqmSfEcve+C5Onz8vAE1SEHHtEWhxY7lESZLI65vOeHW98omwnF/2sKQhn4dVX3/
vYC7HDUBhZ66Sbn0YFXBjNn11dq9BCaK+kn3zjQ6XPUvu+xXGccbLp1HJq+zZvsg
Egt41H3ZGUGWhNlw3L00NlEikJhuNiHX9HO0r77atBOM5wbr4dOEC+KsVEQWd85q
r9gQ59XU8lZW/uw2C7rZbC2WGD4jN5MOXty2TJksN2bw1CN6S0boUh4yNkCsSGyr
GW7/bcihC4tR/p2c3ZX2h4blQqxm+xp+d4h+9LgR4jQAIBERdqQz/WJ5ogCdEXSu
JlUu0Ihz2+Hy8/KOtkb5XL8MRgnsq/YHopfX97c48c2jDTMjgCQ78mp9SYMQ5M5b
HO7D0XTaA8mlgYqfmL3tCnLhmE2PEhZyboLeNjfBPkIFbjAYSa47dFdDQDzHnInw
Mx+L09uGfZTga1jAF8N2TgmnQi5ObRLQV8XI2LD6Ly7UCGM0nRk0kiYtJ8wZzBdL
VVzXYwHv8la1A9EcYCWIbWl+C+bv+26ivefDBC5fSSYgWuqUGraQvDk6Qzp1x4sA
XBwiOlgmLlRAJpy0iHLDn/NU1KAdy+Qnccd0uOq31HAUyQwk4hDZN5wdbvOau2oy
nRi0e7Ort+cBT9n1TUAYbbBwMppK3jD38g7yf7RZSGNSu+rI9/drv6ujx7AuAAin
T0hhEajHLyWvNNsGpM0/mmnUwS222GmMwUOmn8X3nVxJ3BizXhdKOWAmvWWkGygW
tIeJ4PGcgy8gOr/WEI0hIySNM6uuWvEmMj1ojnNHv7bQBUTstV1Eni48kms9wlqj
MOHVMsYHZ1xQjIOW02b77mqPA1W6ephslmoes1riuS5UV+gzL1GGlEG1vfRqExk4
x4smCoA/xRJNjundj2YbWHEibp7P80dZSFUQVkLy31qndHRU/IoSx+yEauBZsP/Z
8MOuvPKWa0vZ8OLkKQBSFzSlKru5j0SxL6OCAnqzaoobC++RoSPt+kZ3RiXQu/JC
zKp1xJzDFJf2OK27r+u/EqTM8/cZACckd0Xdrlvm1d434dDHZ1vAWn1+7q+/G9XZ
g3Hpm4ViKYHW3IQAhLicwah84iFsRWPPlnAhbtm1l5ERlEZjzd0u42TFaJoba9V6
4MHeX+PHSe/K9lr91qfSFvCX82TXsr/mL7uOif/ZopwchSsU5UbPcRMmJjeyCnHY
ZJXXNFpMkDAkQIyFn1DHyAcdoOLeJJ5sbbPDt+3BoKobZGl93BCLuMfIp+cJ33te
p48SjrkfMvUV3QyHREpI3Upr+So8V0jMrFCOidK9MA30mdwFZhscoIubI1orOnw2
//GxoskNC57ylt/dHj52yuuGHBp0L8nUVePClrQHBxcMRRWcQ2wU/uZia0hi2mE+
Hqa3swIj0aU7GJUHMriDCUbSzThCEF2wkhenHRx2SWiQkDcL/JyCt8aJAo0ewtsy
pO0cOYxVR8de38GU9GdhriLdyj+VGfFVdfoz2/g7XcHbGab7t3SuFm1yCcTR0xdX
+LbEoJgbq3GuYUm9FPppW6xeqRS3HgcT+SayR7r6frkNeba4e93v0XOfs9EiQ2zz
lJ8pgRpi2eAWhe51sFCINhwdTxfoJC23dUNPypnzQtWegkssf6FUj7ocBKL2mwOW
jMsQhOqc6zdmQaFbqS31U6BZGPdTlVrxfW7DfbKT0uLwzqt5Mkd17T1+3mK/s8Ae
ySqdDJBzMuNIaan2e4vITkhYU3sdy5DXrSokQayEY0HvTv+a4z5oTKGxX8hmdJ+P
+FXW44+LL+whw8zdMPhWRgbtUUFdQpW6IzZ8putzdNTg440pZy/boFK3cjofEWhJ
BeXJLPgNP7R9XDYhmw7Dtyo3st7eOEzzhCVdD/rO/hOThI14NY70RUrTG6wM69k7
1Pzkab13ZPSBUwg+QJsCI90tEdfbNVJDZBqc8m3n0d72WMaVQl9UDGvDXewEetdx
ajJ8bScVGVeWa87UeJLXf54CRoGQD4bK4zQC7pgCPrDaZAfdTDlQoHKzw/ggMbvs
xe9sP03aqeMu7xrLzdPYvQIJz44xpbdAksrdPodOgwfq4k5Ulcz5S6msu4WUP+jQ
4k8HvLiqfCWb3VhRJQrplrCWHG4qLhUXwShf3zNLCOjzGvF2CIPnTt4UWx9rHY2B
+T1WT8PQVmksEs92cG1xFmuvhi/Hha/hhuLhvY5jrYURy2KyQpMlUGMPeiZdedyJ
FfKXpgeqQPu2pwMWPqyoymYYHIPq3i/UizbumHmJHJ7xHYjsb0vJQOrS37MNE5Mq
QfGQQ+KfoQSSoJ/B8PnUqOVsv8UqaibZU1pEKVB0udabWg2OQfad3EpbG968Oms3
uRwqx8mJtqplgrQza+DHUFdNU+yIQqcaak4/8on/hes/v086jVnQC1AfaiQKjSVS
OgRYEKyxUm2yUjrcke9c3rVBn4nUtuMubHWJHin9cfFBBAbDQzn0AjA1/hD9oF0l
eX1FXKGNzeomVhevDjJMUvFjZNWkJGodjSe4aHa3GGekWSMr+/FTAzO6AoQE+kFQ
jztG8ojqmMLCYmMtxbq/Wc67eSccFpHoZiAdQZaJQ+MWNuGWlKOdD3mZpM/+MUD+
3vgSqP/P2QBKfX0pl2OsXqpK+CEa/vKjnu+ST2WzZTi8WHIUIXQ4l5rdeovSS1c5
lQptMEPD4ltQ/6ivTqJmUAVD+9dzRx7rQ7xAkXljdEboievZCDZtUQBGs1e6zXCC
PJaMHVXgMZrsHEPujj+zdWYwd8ZgndVfPvyRBzZ2Jg4KQDjvUEYQ34Xtq81m0Ip7
UexjIR/TVyvJiBD3qP7MWqFJyoFORfXdYTWs/pYunmmIStFAlj2Z73sV8UqgmF+J
9WLjlUqgX+ULvOX4cLafoMlh4rh+Fw5DZJj2Fhbofp0N5xx02t4s5tCC4KVgzYSw
JFmqfglSjsFqkH1j3LfCFtCMiTOAJ7Vj4DQCsg/h0FHQqH/ljdUVpx89P9IRkLKg
pY4cXj+oVC6MKmGRZTD1X58PPuH/Smep1WXB6aoyqiYdK/x8jE6ZRKSelOl62HPG
3JA+mJuXrSpvq6PE8VWzCyYoyEKHHFEEs+t/nUs6Rmw0gcdh+vJxCd32tVEwhac1
nS/v0/gZ6PHUzQjIP5eROggsScy3Lqr2EdWeSu4Z59l95nLKGeDAAtcbAw/1pgQn
d3hRlryXm9NJD/HltQGKWtADtQgBD7mUV2PML/CzTFB0mp9JoE8+YbO9Ow5rECPy
yMhBx9S9toClUDeoMudrznjDms5kZXAWpwIteT4Yo7fKkFfoJpOL7WU/9HMgDw9L
HR48nwivozHnBKxEmr/wXloyiK3vVsAHBoyZEUE7JW1YkhhoYRyyw3V1YoBZhnvm
V5Xg5B6qQm63tb+HXURJjr8X/4h3jYKQXmD4yMg7oo/UVwI0IViCBL4f3VxuCufJ
pESoEzScDMWGUGmsoyxWr31B28JdUw03ABYIz7CHObMgNdeCzNOhaWU6rW+AdJJg
ZkzBsq+u5eF77r5jkP8IQb1mMmzMH47E53zBCAny17YfqxMlVFKU25D1D4jjHbbr
AX/3bpCkN0Emoi7mBbSq1cbHNQacaHR9KLXeeXm1nTJo92jA2K6LZKLQNlfy+sMi
BB/iyr+RJpDNGbP5QTm0B6snrO6/zyh4ZQpSU+0khWa5ijAfp34yuozOqPXr6OyB
mdIqIV6kT0wYq6aauew3AkuXRmv6YIImlVx8W/EK9ip7A6ctbVPqxS6n4aqMyeTp
+/kJUxoL8ClpKJ61P45T1SeH44asPLzM5D29srp1z6hCNcWUnu5pC2oRlxfj19x3
8dVi9WPMqzB7nD41ObJZ6ilp89HEOzFjex2ztZ4jYM2Dg0P4z+DcBJ7D9vEWacbo
gSCqSs5rxTlxka0aUoCoSpgemsdukOynwDmoSfFjkkioQktCMnv3NCQiFFhsMDLb
AQjkpP6HoNQYowsbPD/j4IjAcuOE24meUWhGtTnla0JFoPYy1jFYk1WgybMCpgP9
fiJKFCyUP9e4i8qouzahT7pZdcfEyZYolLvF2mwtJQkMCGVyp/KKSRg0zZeaH1UH
6n6iyp88eUq/kGCmA6g7gpWgB9mC7Ju519NxuBS1gGHsn91mYsqkOZriRp1E7CXh
VzCTofvww1vXIZxtKDOmH+WvJH3VZnFVXTMo+Kd/8n9vBicSL7wmZuykHWI4hyfL
iJX1TXZk41oE+a0GNG2ZbVhLQ3Pp0b7qBhUmmme0oUi58PxK2xmGQXMKitYD9PLJ
lk7gaVk+beEyZDrbsUX935T8zAfHi8bFkNax+/MphdcVE1/VPY5ketK9sYMI2IM5
hvNgzFDHWSyliIVAIVzyNSShO1RFhpoFrt62KO5K1lj2QAJG0Yn5Z5mutzDTvbPk
vm0uSEt5ybpcLCctnN8kEbovAvRbNX2CuAwLhNbYArj7/9TrVAmgUf6VggWtvn/c
NPXYSoquavubaoaJ/tlgrN1s9wUWj069z2Itk+8g8BVXapgbVBNXTlNSOGCh0eHI
OpEN6Yikoolw+rmTplmYj5A+1t8E2+AKL8ZK1m1aUJbIzWsm0hEK9zzmIJD+iBwt
a63WDnIC956rQYJJZpZ0XdkWKEit2Q+teZj7D3TZwcdl8O4uqY7DlZgjSX7ZtDkB
rBDYrg7XuY2w+Pu+VojmhoI67I6RJey++6qJjXv/l7W8a0cJUop5Amh9ehKMLAve
k4CoBrI95FUKGOGzPvi3exbiqk16cbsmrJ+5FQgyWdtpN3s0S2rUP9SSnrLSGo2D
sqBAG5Vfkhizfd94T0ZCl+STrsbKhn47/ESLId7PNUyV3dh2DVux3u9O6vkRKal1
EKBYLu+0MIz3Cvrq+qHnC1+hdlsvCeMIvKq7TM3KF8eojgfYvqTI3eeZcMtF4/i2
hfw0yHXLLPQ2YNcc/wj3UzOUAOJf4XQHbkG94H52KljrahAnJ542FDjFzg8jSdBm
GcsN+5www5ek8WzOOO8+GtEKmgGSLojztC2UJLDQuLOvkD6Ty/E6/ilHrSsCtKRt
/aCow/J+mVE0zzMqFZSG7RFzHjhnIhq9ZJLlWPVpvX0xxubgUanejx+wSVJ497IW
IPl0MtV8wK4tkJEJAdzSRp92A9L7H1dA5qMR8VjfkM6kPPUEnCTiElXeOzybVN9r
9fnC0j5g9yk4xWKjM2IojNivqQ3ovQKjtI0arXmaMyVLjNBxOkcMbgtq4ZHyeHfh
RGpa/wno8lTZ2Au5QYRJC0CWmm7jkbeTD1UYXa1zOpiv4BfCE+7gXDnawR2oEcLD
K5eqk7ysAnyjtDfzytCU1le60Zm/bkclSgOHWJqSKBIFhiNtzgFBmUCID/HEQv+W
EzIRmqAbiOkRQDXUzeE2+9CQm/TWP14C5pX0R5r5EXZxND9ExBurC0ph7Fu77th4
Sxp+J0SnDp57Kqgk2Pt4kHrRdcRShZ7cOIKW0ilhkT++Kf8TPXtWtFw75bIknWJj
FithDmGDbc1PHz4g2F1rHiKNIOCnGPor+orNjSrzR3JlKaQejIHUY37LNMKvtmyC
fpmLlpgvM+N2FqR5+mTLan4dGac/b+MLdAK0qeYGKe8Sn/eWUgvnaetUD7e+3S9B
gDyyu4VtswGdrn593m8HOPpRx22q83mkxxUW7A7yk8HZ0owu9FlrnpMNVxB+RTaf
O1ytYDWLgXEj35r6NNM9K+TMpWw4zeaR5u7LG5O1gMMyRaSxDCi5yBy0TtMOrpQ/
hRhMRgtqJnB4lY1hrJq6NCLqh4qi0VGKXOxQ24dGo6O9WPDeRvv3JbQAz88YyFKx
qCAsD9zK9qOXjhA/gJX6+eX52hv06FJwA+YVRCvob3DkNywPD7nAE5MIYQaQQh0K
dZSM2YA/3fnfWPBMCd5qD0ZKUfovRnzQm1ZZFW8cueQe6vjTdkLcO9P8ivj4x5BA
waImb0mWDrsKx6/CoQAfgJ70jQy1cPYhuS1Y7GepeqdSPGYjdry0iGBQlWdtMrTk
kfcrvdrNROX3UrMOFK5/OB7dDJ0Q9I11WTK+qcNJJrUazCAs9RiHV2pdNgdtwSgM
ECSaCREnkWMWqV5xNbWzm43eTy0Wg6L/O4zs9aXtFTaiZYeRXOJ3rm0VZ7rwcxh5
O9p0fYFBpAfp2ieQioiHpdolMbevHqA9Bl+gpj/sofk3jfw9V5naWMSJwDQgIMSN
3nvaqqCtIxQ9Jzgdrhl/eWBgR9NlpoSEFcPsrobkLb4l3+qBHPjkV/iABrx2BBRH
17IE7c7gpJOO/xO1KqPirNrbp56bdExxj7BsRidEGAFNV5qbAx2voWzZ2bWu3fBg
p584SQraWOoWGp+YlDTKMBKKNpZo7gLbudUzZ4/QIzZSEw6Z/ZTBitrTF1kL6D7B
YlQ1W8mhoJ5tZu2pD09RwLWBlOgpi/jOt/39TOPHkcwtj91muhRsWpNe3AHMysDa
liUwMHMyWFG06nsR8E3xeyD1NcS31LO0GePbMpj0+XFG2nvaOem7bCXqpbYJ+F4P
rVRG02+61LdMviEymgAIN3TtOsfX+QCxrWpMDNsRroCX+QGsUWgw+oxaNucvjQHv
An1BAzuoe4T7Rbmfpx/dny23eu8RekD4235cEDU8LMymGVQEjG5swYFmGdI9F++j
JEOCmsAk3TjJpx0kExJkZbNuCA3e93Ucg1cwhUuXojZhOFtL2M8Lc7VpsRox2gpm
BHq+/Lo1N+svynK6En5DOy+kU0txIV2z+MawHUIbJm5N1UEQ1O+4rW2XZE0SaRyT
EiSoM5sDEOgtLCsOuNYAqOw+dSs40tzjNFx0eDjDeIITpJMHnCdKLYsySMZP8aEP
6F8r2bt+ueIdC01AisFuV9bD4iKF/s6wtKsCTQcttzKdoRKU7JA53gD+5VF2HoA4
w8B9RcxgUxDW5X5e0uknz+JRKQMA0FTq188HL7KRRdIO9R8XgbQ1mJU+48iIw9N0
23koQWJ1PZb4j3DDtoKHiurKbkAqpH6L4lxFFVB4s1TL4YDRCOpcsQI7EjL+2wZT
AnStfhYebJ9Nx7DhoZmO4jVnrEmYaDzmGhXxIimQbrYgAml10YjpW/SaAxGqC6ht
YVQqUIbKLPTsmeqkrmC1XRE1k7mNwp4/rXjA7adYDG446mspvD6NcXve1ltt7Hp6
RghCJlX0+tPXXQ6qG6VciqTEN82B2t8ApDu+Y0DWtvSY/qXOkuHigQ9+jOoW1AnY
VV1LEI7n65pm/GCnKpuKdRi50K2yiH3K19VPnLoKnLCk2WK1gcrb9qgUxR7uSDP8
Yx1i1DTPNlPHyCTq/Yyt4L6uxpzROpsSQrtj1D/unVgu8MhYvcIk1Q8By2m4pGNw
czpBDTQB0Jefd72U33QkRRduW8F+8EDzOw3PqcH0iPZElGrKU5hUVK/tAHmTaOAM
5zTKycvzyNjDkxpm3SLDFhNJt1PR8b4C8cLAr8U6yBoImHEKCzqM+WaIa4aZPtn3
tNy286BuUpR9+K9RTcSyrV33ogL4maq+2jTWDvHigmjsgvX4y7XtfhKWoQFYuTRq
X/06NJ5gM0jy90KVMxzornsTPgFul6C+ue+nBosiu6wfo6ZD6bYzap9agcXYFH2V
iYzcwP5MwHxwLRzfQz+nBMOIP6RrzOlRF3J8jLwZlI19kca9wTjt0r3gNVPplnW2
fZHN9dyE89TUVRMFmbd6XWqaGeyCR16kLe8aMA9USuDE7AoMYqwfT/2i3sovmCfM
3EMHkufrtzRS6X9tIZ+Hi96A/slRN9U8a4NnrJLw3sZi7Oh1KpIrpcMN21+3Xepz
aw46++za1o32bxh0zObeiaikExVFzZ/+ZZXj7zenwHrgExtwKRk9Jf5Zl8NugqeM
GQ1pXHnE3o9qPif221p0uG0eW0Mar7wLFrzLq7lE7b6RwabfZ/GTSFwPhNs2vYAA
eruLnt8ZoyaVC1JFmhK4Oh+8X7VC1q6D3ZZkH5UyVR1UJ7Sr/bqBfuTiBVLmA5WA
3TQ68SLpHqg60N8bNv0pvqdrp627D0rOp8nn/U0srdPyOzIoFrkWHPdPS2Sjnpl5
uVSqmfB2PP/DdlBQvrdRuvGUhw0Ikoua5pSEJpP4a3J5EdBEW1CYcumU6pfyady3
9LCIfdUEFVXMlhmfZ1Yc7iiojtaOicBpSaruqSqVxbQdzJFH4itljYTiAabTdJkh
uZO5znyONLXg0UD1z221kCUs4CQOyAQzzULwms7BSAmqnA6AFl++uJpuBKolIvIj
flC9rkxTtF9wXkO7mijXuK3CRy84seVoEfrFfCE5UVIhcb3ozaaxic+bdpv6JWJn
LnZ+8H1Dn+qrHYwmWggVCedpsFPCl3W/rUBWP84g9uhKmeUHKg4r2wNWByxE3WYV
MAdByx+v9PA1ONtnO10B1F3EdOrztHQFMyGsKyiMYF6VOxCS5q0hNs18N21PdS4X
MNdt7TcJN08CGcbYUBPexoYPYUg/ixfuFa8qtFryoNYLYdtB3EbuK1/UO9pkMgAx
PKXtkMSXlwXtOWhSdXpihAB0tZdq/ILBCp6fB94ipihJjEYKW1CYhUPRiRPuzkmp
LoY9PHENiJ4tl8La7s3I3YtrktVD4eTCP0Q+Y7IbgG+Kaog5t/3vpJ+3VzboJoMs
c9Vr50sJ2zhAQR2lPsCI0YE4yZtAfcVF/ouAviXOlj12JgMOb+3rnVGOZ7WL/p76
P59YDxtWd7g1xmvnN0IVf25GBcd1cwsHjyPegvjVJ1Xi+pvFQZRPw4EEcp/TLJMa
jVdU1hWQ4Xr5FTeRCB5f+KAsPWXP80F+96X5t37GrEeedeMF1lKb0RC6+IOqgcAK
HQbwqv1n1Nnehf4PWMAyu0CwQTRuCy0HmBrlj+BFA+OCUs6SbHbjyakpALY3Ox4k
QL8cjYip+tXYZqzISDlQrSCR2XeGyfKEgHiQaJs9x1M7+wvrHqUz3C9tTQyfmiaI
/LdigltOMDjeUXbntZP52KGvsQYgGE1x+XjuPNoprN0gOktz51HoxiFIaEtFIu0x
wbiQ6Ht/J4DvUZr4PVV3VDGY1W4v1wzoKD3JFl9ud3/nqSIGzZ1eKWtQhexLYN3w
OgZmRT4Te2ritOKT3ZtBDh/LnuKDk9NRgrZ/MpW+IX7Y/4KmbhRDNP5j+juPZgpF
4FjfnkOujb1YxsiRcyaenxzRhAJ2rAfX1/D3upYDZ1wqxSmFxT/uvRMs7GpDp6AA
Fhu0r4e1z3MWPqD1kUqgRtJ5XjG9QyaGWCfZjfeFb+/ZpjKftVu7g3Xi4sVYvedt
GnUViC+v9IDi+wTIzyJjqpB81C0mL78ylTTgUYFSMghfpbuhWk/K8PswnZZkrPa7
kJVVr3RBQsWcp8PFEjNf65iBVUAEQL5L3BbmbS8js0J6dVZHi/UV+7ESR7rDIGGS
HQTYZGvzKSq8et5JZ/zL/1Sf859Tiod/WMSzP89I52SSGWzFCUWvzZKEo3NolJ8K
23NQboSjcC83+YFJkXkyLK44FY5xgJmfNeg/Oj9jfxbOBE6AO5FZBzMmaRP4JX8n
03kfeLYW5jmKsOGddRy5aN8j1N9ygqN1PmBoK9R6JzY+0l9GiNuG5ule7uhKBgsp
wnixkG2eb9CIaNVuZRS4PQXRduaQGHO5A4iGev4PgAqKWaE9/9GD3DFSNnDqP4KH
ZHXCwYJ2FG4VxLITqvyPN7VmACeop3MCDrmL9/jw5Frcfo7M/uKxQaOmkS5R6cVa
B4JYTBe+FZnfY1BR7v1hRt+pqkTsurHDCrUUAL2ABOQ6lbvyKrElY1bZvfZ7fBSU
NNgjmP7uxp6yaSjI96yen2TurzWN7HQIBSL9Y+YOGS2HpmrkUdnh+S4/6uk2ld7V
k4SZyDgi9mfqYrD8RaMLYnI5DsxKLb6kWRpFZ5XLjUEcr92RJcC4aD1SNqZYeVc1
LYgJtVFr7C4piggZLkkujOsePh/P5McnOjay6uz3rsOxRKyKSXtRPTFdu7TCAYe7
KfwuE4ttJrxQ3YjbPIJutqJiMFcpFz0P+YlkwKeA+/n4z2Wzm+DF9cG6WJrsk7Pj
/PLfh6I1Cz3LmbWiF47tRFzm4Gw/BYP679IN+uq2k6bowBIVdkT+L6uXl27IarzX
QpwAJiydEtHyYHweMc1KE+KjLl/Vreo9hY00MxyphYRIHWvgwnzIo8cFxSeGOR1J
bCWFJPvFLdwbwUMCXdu9elMSfW5APcye/d+UWWX/qWbqCOxAmVkhUSGs12OJXzV9
VSWRGY0Ze+bHObmnD6qEsr7i5AT9o4ZAGWFL0y6caF+K1UO66ATZjWEB5vcOlGo5
68snZcdnwckVWe+vEFMHfQH0s5z7LPtw8ogkj1p1DTU8xwr5/o98JTW9vv5x6jxQ
CejCUjhT9yFzCa2JUvxKrWJjeEpm8TFGqrOawYM2wYq0QXznmX3+fTE+KBKpn1h5
3BxRk9IuHdkCuXRgLY47ub9A9jwwlq6OpxpqEMNLdc+xiGkfRlfpdaTkkfxfOv6K
xH3PBetMdM9l5EnrirMd3ZagoqS8tj7uCRV1KQT7DHXU7iKeMzDNKlKq66WsgXF0
C9T6ehqfvmgEWP5arfI5slIT84tDTnbjIEtQBmoiJNZJUUkcGKVFlw7v2w52Mte4
Lyi/2gjQ7FOIk1bSJg+LH9WpYoJpMejgL9Hb2SVE5Ot+pUqfIufB3Vj+D4dgAf5C
BKYBo7VAeGQ8FyAkefQpbnsiBojd1BAUp6Y2wHAMCjL1De4UBySTIJgOlr1fL+xJ
XFBlkIXisbq/W/Rv9b1C3FpiNgLFMNjdotdeaSZ6R8Ztfci9ddVvnyzwh/yPwTyr
A7qR1XrhhY+jCyWfM17z5AzHVrspA33E4d7BwsH7jPcAtspRK5w77iLh92pzz9yQ
msMTSCImUrxXvWZm8hcOgTM+E27OWEtVMF4JUaWMZS8Xr7YQqiGPNLkocjHIxm5d
x3gEsiwYeBo9sa8Pg077GTOHBPSiD0grn/3+YgTMADgh9hdHm5+KB1Imgp1Dd1ZT
h3Zu1GBjn5WsW6x0NBht8IqsyawGkvZrvvfLbuP3ff+oI5uNIkA79jThdYPtPqip
i9g4AMc7vIzj7/VA3VR2T+8WoVvdb8HUEHtROv4/Qaz0RxzMpvr/MRlFeVzW0a0t
zfbKeRQAeIDXrdU6PnIgtGyKH0VvnWKkorunjH9lIH4aPiaCMW7tF5u+UJo69rbV
jcQCTd7rpM08Z5BCE+5vYg1D1NXD0kDLg0UHJ7qgv/2mQGXuL4RkeLin7XesoCDX
SS2YtFn4vGM7fW6aPvv2w7JkZjWrLZ7cUzJ9QShm1KjQ5rX3gM7WONYsHizti3Un
g9AjW47PnG5GFNRZXahoUtDxCpkHgUSMkc+Rz0mmTOupEss8HiJTHfctpcMozQyH
q8lSGR25QGt8Gxz68YugGr6FZzL6sk6sDKo0PJ9PBV31ONPA8RLERxtcsAZhINIw
kPK1DavCjAMKazy4+O2ARNodrLK4y0ADgKiL8URVvSy/G3SUjlKM57YpTg2jlyCk
eLudD/4t4Z/11HYa30xeRxQngWqy4mL9JkvUbUN9ggd95+mausyxQWq+uzQyghhh
ruSIgkd6hk8ylf3jUGYV78DlYYk64t8FA2eb0UbFYN0gHLHY15zldTx9T6OhGvB/
cOJen0TfoD9wdsLFEmgiQIshYEUavCsi2rNxQcxoWZTCXOzj9bW1sImE5s2pjri0
RYSkI0fJlIbjqIJi8ljq9Pc870Um42pXqHFEI7jGfzagYsc1Sd4EANrZMXjivL/q
DLs0BogNenj1MXuElyZqpqmjhblixpMSQH7H3i/OP/A6Bf1+E5EIlnXa2+6NTuIO
hcqDSJOIPjISZXels6x4YQd0kfVfyqcogS1JXkPSxsvWz+QqvImy8rLbFxEDBG/U
ovlloadgqYUare+hRWWM6M7kaoKpigGfRknuXA4OxSQEAWB+CPfjxJ/fsUAJnR/C
RaNuON2qbQEalUkOSIrr8ZtxqBDHuyuKou3oVEF8xF6mOEeIYT6/rAYfrjRoM/Vi
zDRNSjYr+D4vi+qm/Tk5N5HVJolWD3YaCZqyKaQYc8wu63mCg+KpoaavMppRe9bU
lW+cg4sATL2mK9m41PhP25OLLGNDyXYKH/ZKOXKASLf2ZPot3yV/N2pj8V/kgO/J
SJdh5FHoBXPJLaqjmkSIjvGZJOjt0HIdV+BmeZfhywAc+c/bRdhGhBUAFvA5DlLm
qByIwp8rcCtBBoUWQ9uGcdoH6wxa36yPzTWYBLBdVbvd1WsOqv7Cf0K1mTwSyPDV
TSBXui68Zg8ZtQrVxrHGAqppS5AfV+g+NU6dEnujRF5T8bxi//Z2Co85Lm77yzSO
fTlOhekILIvo4DuRow4oZjmFYqFlLYzH1THOn8+6Gldfgy5IeUINJmDkFReduMs8
Ywv92zC2HeV9ySpgOBHV4aeVaHhBROwQTU3yVjdu6AqjzNFZ/uH5kM6DO1p78V2E
fHXg7SGj7s4YKBdVgyIOuZIkejNp3uLBaElMGapyAREfCQUPs6wEDrUJnqFLdkCG
lUv1e8occMehR0ok0JjZBfT2VQoD1eUjkNfxuX7lVTbUfOWwSPuC6DB87JrnJtXR
ZvY6/XmiPvxylQsZ+EmWSIaTtres17+1NUqEn9tau4RBNoXvyS3qBBCMi3H8/O3Y
cPijX0l9vbCAYg61NXcegPXiWUdMONb9NhRp6s7pXXqF+SzMEDlvs2Wuy7zwlpK5
V51euj4W6sYt8Y3B6mus53W/UOlhKDlyc1+VDdtelDTto2qD8SoPJ2pKgprFrGJ1
NJqB/jcAeVL+n3n16FkYuOlb0o5DOyId7DVb0vaIMkLv0sHTeHQ+1jBXKAbLNYWx
UgvIbtdsDSKQwlXBbIPnPkluc63KPSvuEfH/KEpqHyQ6jLogkTKBmEOBFdTQHyzi
GIGBC0I7QI/gNGaV5z2inEX/a1DJx2D9sK/ZGnyFRA+Q3VX91dkXf1EZKdfoxnof
SBZmG97Hg1hyiO3IvdqEYORYDSyy9cStPxf8XNI0fHGvRJ0U/Y0ewununWy+kDpW
WPTAfMbgFVdcyo0CQScS1MzsF/kMPKhxyiFTcYlhq0crO4aUWRMlbFIWfq922X6s
44Q1yhKjV+TfRIvKKeVLl2btX9VRz7jt8XX7FtgsNvca6QZhQ5s5GcJSstvgaW5Z
07Yv9Si6UMzcw6fltZe32Mo5NfZ+d6bax4bCnVC6ORbtAJuUOCGzo6knlnweA64B
g6sXQUlb+nnBd5LEwW2zBFTaBDOKJ6s6TGGmL/myV5IWeRZ2sLKYzCof1H6EB2qI
KHWfT7/zQrA+7iog/4NygkMR5TbBDQsKZsd5IgRjULOP2WmkqEChNTYRU+oBDHN8
Rr0rMMD9TxUslEpSLjZwN0y5V0yWTMfmXBRfLERp1IGJRKlcgz1kxg6ssMCxEz8j
6rGHCiTMMO32tk0ltznamhAXK6FZwwkS36lsynjiGCUmoAB89vtdD6mfvRF8a4fV
C/YaBTR/Gxc4mbOcM62lQmTvcrs2W9V8tnHkQ9ybjwMHsjfVV+/8M9kKiTTEcBfE
X5NKmJl5PtMV0MaRMmPrxiRonvirCXzQDF1iFZ4AGiSiwbmEYukEBa6kOT2xCSte
3NveGLfw9b92ZjQV7K5GCwyH1rZjcXtHg+6Q1ecq9sk1jyOjCU9W8f4bT/ROgvpU
OcfV6dUPOOKYcCS8IweIWtZuEKcpOZGDSg4VbGqOWNlfg3602C7tQEPmvU7+rE4n
hyXSE127ACsdi/5HW1YCoq/tWOkzFPCOgsE8ss1WqV3F5Ygrz/VBM4ahzIjU+U6+
DxpZdUHm9W3yVi76WzEPR1OkZsAJh2n7vgDFkyRD/XZzz1/WV5Pb5FllTEqMceWA
27gl7k70n8f+CX8wgtr8cVoTepl+G8ORjN2SZBV+zROqxWa+c8AeCntSVIrcke1f
aAemTK6qZqr+Izuk5ks4LcIE3xpXGcrr4p4OEKLippzLfOfInT5tZwzBmbQn7nGB
MmjcPE6ltfjYUWY3apAeh/OnIE8EZWv4g4MUtg+z8RyF+FetwuLWW3oCo2YXvulx
66/+yGiR8ya/fxTSv6BI9quI1YcLwbFul9VoUr6WDk3FSZ8QkB+aSoiLl/DQ5n1+
9K+p+9X/jJY+/Fonk45+a9NYUlqUDlfzdYRTZhX4GXMajmTvCnYv9T3miQGew3YT
Nnsf7RhhCxkUahcwTpY8+8kX8epiK2FXQgRdC2cJ8iRon/N7cmHlTWiPQcXZRmEL
M39Ve2Eu2pgPMavW6kSrl5ZBvat0HuYkE6uCsQ1a0IgP04zyzs37VHYKHDlcvYLQ
OjpLUuzh99tLGLxTGy+obja00wC3LFcdgPy0SntfXFn/iIhG0L6Eb/faENzx2tK3
IAZVgHkI/1PgD6GXkUieMvt7L06Pj78gu+lqM5jzUXZF6gnw9ZpNJdmkJ3UaTeOs
49YrRAzDIlyDLBu0j+Qd9ErDwgDUMCzU5OGQxt7x5UkEVeaZixYBDIxrspDED1Yo
IZTkBt1W+Gg3kUUEuYMLEdWLs2wRPfu/Xeq3i0NuNopd2mPvEslkRYH9Eys5YZld
oT9kEOEscwNMPfapGcB32UK8q1ahSmsjT2/w5vdmr/2rTTPkweiVCQtb3ESVewE/
/fJBBGJYVJi7bEuoiTDURs/APi7wvDq3o9aTRhpvg/tUiIKToqFeKC13YGqsa/yg
soW1PcXkZbx6WPxL8HXkSwZrX8R9hXJi0C83sNeLgdEM6KKvFrvgu10fRCGq005Q
9vHiTsD7tAlR6926wSXunxg0u2K+ASrWi2jh3hCwHi90GoKNcH6ONhsZhBLRVi9J
pZYzs+ntoM1F7fvNLWApoqya2giSBgC50uIrKH3WnfiFBi82ESGYu4G8WuG+t2F6
SBCegbeGJRVr6GORoRiJIcwMWrEk2FUbllJSLVKlyN/quacQAR/+LQYInNnILLHX
7v2BPMq4FHDs1MiDxZBtJ5fnvOTjN1MeJ1CLCbtkDUfMPI7QCVViBWYhkRqObVns
5FQzc9iXvCfhl+v3ijR4eK76af5b24MaaeTKcCPjuZBqX+LRCO/paDwJ6puPuX/u
DH0OCB07GVY60Pg9VFbofoOW3hQMjtfya/WydEpoKuKnBxBNxAV84mv81WO3QvXf
C1lfC1fzsSeflBg3E4rvT+EJ6ondXAfCGQon6p0jO+4tBTJ9R6X2+ZzgC0wjClhp
o4zOsvKtZlKFrveZ/9sycmjecrFjbwL4EguAhJvu42PNpd9YX2yHdGrfmiZjtq+x
tqzEAZdeFNiWstDmwQJhXs1Wpj/8cpsIEx53rlkd7xRGurWru8927LSpJqazPYQl
xEdhhkpD2rogvtzZXSpvDB2f5ep22KlqqJayaOXvGenyf3j4LM7DMpbkB8wrZscO
BHZjf55u7JLXNZvvxwi4gsVvX31614MBQfO/hIrIU96pLPvO9Ap/71HDHeVi032K
JCpUDZEGA0cgrhcM9NqhYN9Kzj400Naljzvu/FpVi74zq4x0akYL9Z1XOciDj2bj
GmAjAYKLebVYOu+RhGCcQqtjccHKWmv+OWLdC4nKTdNsYFywvjwyNkDY+EwltB2A
PX5C1U+VQZhSx5OrenuW1sm98tN+JFMOjqGju6elS0H18M+N4WPXdvkp+KKJDNSD
PxAjWSRhhIJdK9/Oi8Lo0/63BjMqfqtKySLMHrBWjKCC8kQnmzCrixw2U794aiNg
V7qmq0Q/uekunTEjdok3hOzVWWedRwLEH2DoPldrcUapkmQzHlt4+NIg1NyzeXzy
5/EFf+WLHxV49WFzjZSaXw7iVnwaeYKmht+owjAUgovrkFdQSndQBbBdP1b7IvLT
LBKuipjaPOj2ilrdUrx8FilzsJOEzd8R67GDMxVfDfmgag1MiOuDS3rGZJHMXOuP
SjLWmhMNdwAmf1C5Svt3yHxpUCvtjCgouwYsaYv3ILXWgerltj2EZl4uL9bTPOIy
KACpLhPp9a4EMtNIjeyJQaj6lDGgb+wOd3dpd1VG6ccRBe7eqQKflXfL4EKxpz2P
FUcDoKcV4jTaT/pIzmuuG7AEBylKguWGj/BdMGibPjjiW+lX8iR0Iukt3p/czG17
WvqcCz/hjXuzuCudblzsN6MOVr1n7Lu2rI85dI84C+6JUwFoUquNXFIebg6Z9m9N
b0BxjXrt7RkggwKP6yr+7+7f5z+TqdT0swc6COq5a9qKt/DkdJPxZXroe/PqWu+s
qLwQueS/L3zV6LNEJU6VBAO0xTBjkcmpDchnxxrPKJAECa/EcRUU1Ig1naAEDozb
pnrDT8o1bsf1VLFqYKVtvGvSjlcj4SbnNRnvAwAlSz44/DuoV1ldy1O7Y7hNCRsU
v1m3EvNATuI3Yx/pm3ekssqrdD33jpRt9iEge+Wl4M2KMs/sPtnd9FN9hV5BWjM4
xRl5qKinefkZ2LokUPLq646Jte73dNDvlLvZchMtsJa6tYTi7QszbLiGI82AYLSA
1Wss9b0QA3tYC8NfkwWjuwuAN51yRc6K0uL8Di33uej7bIjpoj6eIDIOvQQ66rHx
HyrSNdnJoF1se8kf/WnjvrhX15ZrjGE9Rwvn92gwuA7YlmPPvatxUhKCxD0fLCFv
atceOLpt/apiEZodrL69Jbt5+gu3350ocM7kA3im6cyCV9+0H9vWoHb5yyrw39z8
Chwf2FvoV1BhTw0j4JXK7Qbl1j5uvHKSwIOXta6Z41yVXsMcuFF+c3mhU2CzXEK9
D521i70lRYxDNaKdr0rMsfp331/XFaCcBvbjZfky9S3dcdxbRHYwOrT2Ucj8dNCZ
TwptgR8+jx3r8lIqnJ9HnuAP70ijdzSH/lSGNgRkudwsGueD0AetttuGHQ96emMi
gdRxaQ+9N9x2KakSXcSYygM0l+J2Vl6b0d5/XqpmY/kIcU/55ig1D0tKcT83PI1W
/rox41wtwQokEF48lgg0+F5N+67wFHlA3EwpZRp7PZrtcGxtCW+CfQhQZEV65kTW
XkPUiTO51c0b76Wyjjq87al00Mb5dn5mhVctnxaBbnAs2fLKRbmVWqMLqprspt/m
6/beOsCTPCn5NzqtsJr1VVxeT3CZdsL2FHKDCBVxMSAzzar228cVb8vkQRJEMFoc
BFRlTWixf0tjTOFR1H6VKBgTTMyEUaimvo/I7GDjXJxKWv3Ss38OgasHrNJGxLjy
Rri/nlCWiX4X/dbiOWEJ2orpV4r65KXukpBCv1xYM43sjv4k4CnJvCozanw7VanU
No5FJOS1Q7e+IwXfluAnkzEYbXII9vi0dx7pMKrBBBE46PBd/cKMoyZYfVb/XcF5
Qwk8bJZjMQBdwTkW/xywptAzwRMNq45VCDmanIJ05psL7B1ZjFkWHtYQD7gxIASN
3xbMbiQ6qgxwJnj1PH4Lcbz6KvnBZ7bT55mTsPkmFNolaU0I29PkF8XZdZXC1a4L
sJZF2MihH6w47xE6z/mvVzU4ftoH10HgatBFNNanWgSx0EJY/iqf0SCOKnSz0MIx
fdwnAS2GTVlCWfujvKfUHjYuJdekXx0Pl66lnKuOCIoDSIDn0A7/wBi05lCxglOy
bVlA234i94iHIn76sYyp1W4hxeBAGDvU9S17GU6ZagkfD50eLkLqycThLLvosk4l
WMdZL+AvLOy88DtIJL4w68HztP1r4mW+AFZ9DQF6+9J5JHMV79kYfBwnBYVtgfDb
9+Z6C3fVRhE5qFudLfaQSUQ0v6Mz2TmR+CRchPrO5aU+QrX46Qw8VH6kBQN/IYXG
U0RsAgXwxemYuEZBzARtVE6SO9ZRpy6ezPXdIQj5hELEnoeVvvEN+jQ96I0nuupQ
OEUEsqMfHcn1yuD8DuI1aPojdMtisCynGv0EWeIq5loiSyBQWFAdcGjnfZUbCEr9
g9+jxeiAb67yQK7BDS3V2aUj9s89fdZT6NqLPXFTb6GUKWZ8jazNzg6wO8EtpdLs
P7gqhY+gyuq30NQUHpHo1fTg4M0iAQg561yq5ZhY5Tn2FNXb3+Fko+mN212TYgM7
wm99tt/i583BVQfWWtA6l2AwU2mJP785+HMkjJKAq7/mkpf3PmahXGNa36LNJtsR
NCMlDuYvhOquO6C8rIW8+f6A5PSF5tq0MQ/WtXu3f++xJopksuPiVfqKD8keOI0v
Y5iCowiMx1ExhcvYAvAGtz9l9HH6lEDqKKebfN/zipG5ETWnaXF710LwRfO+EzeY
lW35sVTX0IrVP5yq8t1gJCjXem5mwd63cz04vsaqcF378w22bBCtBqNpd30htn+O
rZpcWyM/1qNT3MqVazb8MDe8fJqTQPjvY+wsE+ZpuDVPp8Ye5ScMLkHe9lUNkiAI
AG+v9O828I5LRJcOaBhDXm8Q5SVlxQS1JPK3gRjLKKbNZrJbBvqJNrX43sotzNOT
EPlpuoJP7uUq5gF6v6bVCYjl19S1EKIRfoPUDKm0+aHlX1Sma2yWcYSz0G4ORgd9
mtcjLgqfupOTJYc9hPkaqwUmUYsbTeneJKPayxIB9HKXVpcP82Jwv38CiCeY6G+x
RoORdSt1MF7Wf9P1S3jdU3tds4aHVWjw3RFN6UuekQ02zXvklSKfWlJq1kBDMK2B
iJvvxwgzIS4vof5RNMOWdCL43IqK2iEArsnj7wWB7zgkC6b729NAVwFhefBrD7YY
cq8ZqhR2BgHnO0IegJQFVIMc4g8nzcSkGOjO1o1U2QJAkfh0FLUk8oi9lC0Qx76N
f4iND63czyLuH9Ci7PR4fM1tUM+XPuSTsz9qmHXqtxbPzJt38M7TmbiHYGUHMG2j
d6GcQam0HYQ2F4zZcMF+B1MyuXRw02cwDZSz6KS8+tCtyTQ2XBWDyg/TQMsgfNK2
59Zo4wjLMJocgMOGoDKFAgqwh+W+F53mXv9FxR+J+VU1vSOZl2nYBFTUfSju5HbT
z47FnVdz4yiOgU/EFqBfkVaXWBrp7MDrAlypKxn750igXxYB6yh1+yWrJ3HM/oqo
odm/FDwZgF0Qq7v+znbX9PQqi8RYHbtGtQ/1VJGA3fA/aMIicfWKTftvGe4v/3yA
L/X7O1OTrSWwLAAHjD4D7ez5rmUxzo73hipkasw2M0+3OFweL5zsH0obyNZtPCpW
+3W737nbWe39U3YhT5YZLPPP7s6+VlyOjFv6Jqw1BvS9Z8jnUKWZZdpR6VfgZr/J
eqQsSs71sJk8sd2YDUpNgbMD0xUROvH/Vc324PHSiKkr47UCMNR93Yzc7hTEQOBX
AM3dM8CWb6W4uqV9UINEDrqcfVDqPcpVO0q4XgaxKsCWpaETrR/Ex5gXLaGInjiV
WK3qZo3OxXIp+CXN4thfefucRL0K7N/AyrzcNZVkOMhBGBq3+rJlxxFR/eFlcIS7
Dqr/D1t1q1/SqyAEroRr74y3zefDlpnqnO/SOhOjLF7FuD+NsQOJIbB1us3ENzvg
vjZunS5ho36xVl6Owtmc6MpSi+9k5LwyR+rSLkk275uI1151S74GVVC+++L7smww
Ji9G+31oSZhLOz3ET/589MR3hnX39GiWdQvJec5A2uXm92AtEj5upxMSmqTSPYF4
H+b2/0AWLXJ3hKVoNKeIZmzT/YD3gRFsBjrwW+ZhUvvhD+rcFxZ3X/wxWh+rV0JE
alU6f4euXWYh2dYLdNhGkJybVaC4QtYges+VOp4MZINN+n+6PlYopjHjU1a28Jh0
WTck+tP1ZyZ5DhYPINOcgtajmdXRihI7gTncoJGo4UfC/SSliH/n0asO+FQHhrrz
Rtmp0+gMvBE+CulwaqbhJIImu4OKdFiSOF7TO3v8tLq9il5NUEdX+thl323DkFcm
uEFZ5HtdVcUmgpupUlZ9/lSOcaWq3ck6naHLCtGUsKCyQbiFsj1TbyZ/OnESYZbd
pfRi9MgbVYCRvxVVOUFSfTSwn12+2zFYT9rfc8h+KzFYdnyhfK1NDUQfwQmLnzrZ
0Y4j7YLlbpXyzmJFaKxXr3bZ2wm5xUEIj4dOt9fQV+A0yHddZIUOHlHnYgKXtTsc
Ep6rVjrpc2D2mAD0tdilrsP2g0IFUkRlk5bu7/cqr/VnqUBNSuJ2At4ci82N0InB
rbOxKJKTA8r8Rp9MY+Idokjl4gVwVWiKH9zxcJxPsspIwJSf5fcz+GnhVe2Ko3R2
3+hjpMb/zgzUjMbRHrlN/yj+dLIvMgBHAy1OmEZEICLHB1VkO06lc7HpFrumF1kW
bfjgz4P5WzuhKwob240BJZ767NWUN2F8NYGru8Aj2rd62FVw/+ohI+beYxzLyHoq
oCrXklz8DwuYEZUXt8VpVKJvItAUSPuOLEncoIa2qSk0M2vcruqBeZy7hDsBFJ99
0j1jMSNWsUaTBLWQamrfczmN5uc0qKStqkwZrVWedO//2sHY6KytoBopGSCNBgRv
76Q0y/gQWL/PFPzLCwFpgNPLadQdH1e6EaSUHeJ3g7nitNgnSoTVZ96+FTlTQTZl
XaiqJcjBK6n0YRAj4WEDdeRiuuse9JOmTHmOuab0XYbFC4VUYw2UyNy6mY1cApZF
oY9L277kh48KCmbxISG4Ln9SFt8AdEDCEE+25sNjCxLAYa4fCTSke8J0ce2dzYUp
rw5Y3RAJ+3NeHAKp6ra3H5M/6x9U4liTeZn57DccWa+3FWeDgftZXK8sXMFbQSce
SP8eT29jZVXNHZT3Q69f4QWViFRFMGjueEVEM8DmZjPW1TtAjzo7PMnqOyjcW2T+
ddgR9jzCJcec+p3KUfHYCPOCq9DF2ctBIqrjfbdeeVyfpTX9WuZXXaGyRD/6sq9F
VIsbkaVc9C9hewO2ox8ltkesvHb9VKqqJHwIYzO5nh/CQFeIprSByR0PQOMZy+aF
TMdaalROmt42y1n+oBt7FjgDJ1MNWYTEpEIBEG4pz+7itElKeqEfo5x6f2tuRD1O
OnRqk7hhnxRDLWWEiW3v2U3K/ex96fmlVUdWfZXw1HEGrwOedB0fyZrOhwy2QyB5
7Rp6VGpCl9XXXEaRTM0VagudXwMLEKzD/ttRDH3fJt4WvA/MOrlcmAbqOxWmz55V
9KB+0JKvITPbMZ9XQgXhJ3Az+W25SdU4nHkUWD3T/YHsbph89cQ0LT+YlDk2jJxD
xQpNBcfYeEl/NnrkgIK+VVDM5UeHsKMZzsoykJD2KjeHsX2rLPXrF+otwCX353q0
1siauJNHHhYcc36/FABv6G1D/ya8f5WiN+Aa+rZfx29W+1c7ZTHTnMCggSxzILki
rzNpNIkKDXE13leLQoFQ8tCEE0e7Q6bqM6QGdKyrnNcs6kQnmitbV8qukfod8KIx
k4qLkKtF7dWt1872xZM0uE6KXc7eqc4uo1yoTuMX9yFzB0k2Fbv4rShc53NcNK1E
ZMqkrPVavxQ7dpUReWT4zCll+t4nuydImnyN4HpGvH22Zj5wukokF+YqOjfahZq1
IaZZsCG0/XAd+yf5tlbhgUeG7L42W4M16fUMEnxXxKjyA0JtBH2N2rCjrfnw4DZV
78TySU1Hii9xdIjD+hrPOc21KRykgWmW0svgrVk46LJFSRZdttH8DNaRWIRWg1no
Ic9Pex8ToXAUwKWflEiskfoqiPC73f49x+tTqfGR8rDHAPcg/eYQVdLD7MPLTweF
RfTZVL8pSV8mGGrHnOAVeAABmzQcvUyxUspii/iidpvTCyADSHTZjrDv+vaP/PmU
Rk9bR6wPLniEyHXwnqSelr8Gtj8GtelLzy6ZGbLP+7V0F2jdM2FhEtcRG7A9Om/Z
LV2xTaJoFqcqDzBv+UPRYbW6gIZigoeoty0ZNCUG0wRBUjid6jsYnsJg7WVWNIge
WR7xvLvlrRjU5on9u9qw3askKElGuswRazXpvIjafmhBCteIRVFbV72kdo0AyEB8
4u24XpFRyQGepnBVWsmAFpDZ0ZXlI4iOq+fW0Bdfl58Nbw12kGjg6sdNjPiFvdat
65197HDHTMDNgi8F02BXPz88iAUO4EqGqrHdJH0kDUCU3zL+xiZ1Gx82/fMVXxbw
C0RtIwLAVYfm1Eq+oIC56Rpf6Q5BvSpscJGWyEd8HaVCCHAGbrNW/nGhlyzELhXA
gBDnFVuny38Vim2J2BVOkMTYvMoI5hogN+YPlDRFyRrp9+s09t+wap8YgG7qdTsA
7wAkiRE6qsu4HWLFwc+iJxaJg3Ey4jqMhBsTeEXm9LPPhGRfKBVAMiNgM60dCylX
8S9V6fzyCXBXXwtg/QX11Tk/pR7qUwoXGlTLQwdvzdRfaTMfcVRvPZubt4UfxO3P
FCcsexRF9U9Dq2Hlg5n5HIQCj68cUJP1r893MV1OHfVIe8ocI6+HlZM/PsZhAC3Q
0BQHg7VyBORkpZ8tX729Xu9JFW/2jHSDQ0S0lcHFTUSgzOHzLm+PLOKyKLIcIgf8
qYRwhQh0mFQ5ustgYjf/BeZhy34Tui/DJqgFoYenNseTR2Ca+1NU+VjSrbergbqw
IGZRvvl+ABPDoKabHBvuQT3ULytUBa2t9ym+uPxDg/CvBog2QImQC0lCi4eXhOL+
/oJ89Q9B0BvK9jqyDUIVoXvk5mCE4YXyprqhXdZUeGPO6XoiBgJCQ7RnnnEQYUQN
+A6PWFOYAVWfKYoqMqAKelLd3LDs1afCmvLXttETXeS8v+hqgUAK9qY7GbD7fJuO
uNHyNR63vOE2a+tnrJTosBpl/FHCIUMmPy+DVyl8ZS41qZhb7hy3GK2YT0htxP8o
VM/uw+4pFBAmu4EUpVQCocEbjhMejAkpSTyu4lqoi+VTAmN9N8ywltwBpYPUszuz
mL5Lk6eYG+sKut52ME7oktHRVYkjNWyIwHHqs8mThYu+vrhPpAaNU1yYXSQPVp6Q
U8ZPNvJXis18fI3aXrPV8iqY4PYHC8af/DqxJrAdQ1G+kpZoEZwAN54zb0FXiVFQ
+m4CPRHeoWlyJR99Qld3BlT/8/2FGgmwVhghkPRBlhcRHgg9Qw6BkW7kSayBUXXm
rIz6RIs4LGKfb18wc4JGjcHR2s/421zf4II7W7C73wKgtHkO+xP/JfD6cRulKrQS
915/B/3Zospyeln3/vFt9X3QkOYc8v7mgR8iiLfS8VkRzTZ9esKFZFa4VKwRnb+7
S/yPy2nkSMASfsZfIKddNhXWYt1bHUglVWcU/99j/lM8BSoewB2jq7rrzhWCn5xJ
+JXVEVxemS0uldQW8dFz24BTni/7o73bohTlgT14ZTpJPUW3llvF0thsAyyo84Ls
OvRET3CggrWwEB7KvjXqPnwzLyRmWDjS5qvc91zTFe0Z0o0lHYTgumTeE+Pa1/Nc
bFZFaIUkLydSyMzXtp2jIJTmFj7MaO5L8W7QWaf9bw3oskkdz+71A495w+3M0baJ
76DU7nrn0mWKpOVUWhdg8p7eehBEeghuUT0U15PQM1uwVU2dLh3BoBldI0zkAlux
TmYcfiNh7YnccGFee3ZHpsPoWVhZXDgfeNhnsAFMq++ct7E/4VblT8bloCztm19P
4YWNffC2qEFBIUb+XMgC6m0MO2N+MVOjfTXbpuyTtNzF2Haajlj6Too3Vpd1xfhj
TMjXbyTtNHYF0AcSkIhQ/cZihbN1U86/Yn74UzFMBAlsmAcEFvfTLUTBreCLC3Lc
aAZiNHqQ5FJ06rgJ1qpFeXA5gwAsXnR8fw3Kk+7mcEhFkBX3VGwQjjhtjopqOPp7
KMJnji+S1gIYPpOL4Ob9teYJ+o+YulRhm08GDFupRxrfwozjH3Gbif6YkI0DFBjU
cExtpn3x97+R+BKaJ+t6GbJyFLmRLgMSgLHPLwKd2u4rLlKfspXmGkqwSQTCYJzY
STUaUrIb186jPGmA+wl06w3YP98txwlRU2t16tCpMQfwOEnDjma5xWYSp2T4uYHL
ox60Vyq7lGIyjvbUNUeWzYQVcTnZ15krQY3oh/wuciEnn/ZP4t8bRsCcMA5W5pCN
MkTM6x5vcfOJzFUyJhJvH/IXMfMV3nv4s4VyoepaeRrWdypSyaI5aRHPWPCWVYjF
u3HMu8VEbWVgnqGdXkxe/jOlnxldkMWrR2bK3GmpmLFWtSyJrkFHM/55j/iYFP/T
D7FfEpD7a6dxnF8QOSau0le6Yd6GB01CVNMm91ym4WYQajfLFXAnqhABwIFR8VQq
kG0BR3vlg9Ncl72z/cHhngkvIK93Bo8U7EX2FFOw4rnfgj1ilYAkqzJbOfd0EKLZ
0i+oDk4N/8CfvNQEUPokuZ+mJYhy+YbEXePFgFr356oRuNsxvZQXDWw+bJ2uG0Ej
YJU3Xl5VDIl1IGZZKxxdLAHk/F9298VTEaioIIpnZKECdljsGD7JpQ+sTDv2JBgN
/aXRul8GgqJiYtiEreUo2obQ7aWCm72G5BgryQyP3LGNSsB91246y7wS42L1DKTS
v4Flf9K3RZqcP37TewcxYmT7chFLcGqmj5X3oUT8BdAybQmio20bXFuSu+WzWW11
3IewqFSEXhL/r6aZlSp+Y+xO8Z6+/hp//bKwOMZqzHdKkV3qIUYAHC6WDVX86Dxx
s5G5v8zl3kXXH+K8gFm1CJ5j9jHo5j4FUoZ/tc/js9MjHkC1PqDjlwPcXBSI6bjs
5NPlRo2ADckKbv23Lw5+FE2DUPptunuvR0phE0PNziZj91YSO7qajHCzh04G46jq
G66vdDvsfDfmYcMgoLvtW//GpFVE8tl7myxlgN711neF1gWr5T/YV/feBkleQmVj
KSPi+KmiPUCJiy2nWtsJEGlbwcnalqjhwG4T6ji2Qdl27UdNeTp5kNGo0ZbYM2qw
MSNHmfZuwBgO/r+yg8XridIh8Z71ZNW36VD93ksvhJ5BdKsHJdH1U8kXR2dSuP60
VHU5Dmpvp7g0q/Qqx5dGDfFcZL7zlpEcPhAeuDIcG09FQpO7Dz54lwk1NUrCo/HY
cpXVPQj2uf5TCP+/vUzGf8O+gkw3FHwXHnycU8yTXyEfA0EQW7bttJZXM6K+oFis
+OheMXG9wU1OkmONgNSOLz/AO3ItV28NZYeJ2UufDlw2Vv0dyRHyv8jQffWyBpe2
Z3lJvtvlIWPpBFvgAkfJsUmGVmRkGG/IjYvCpCOxHXCIrXtEXBCg4sHgq9lQnJIy
57W8U7vyATQtjYd8eoZ/sgjVN0eG3skH5qxwpqJK/yYXKX9OSVLE/K8tl7jcS2eb
f7C25DijYcu1rTYb2L7eATEXZz5jA5tLW5jQHMOYjfapypP1HlpFBbg7Q2HnuSzJ
gkU5Gcx6yjx/xExVSf4JGSTjJ0DMgApGKcXb9BK5JHuLmwCuqhra8pKMAYcK9/F8
2XwKpwKNNftstM3Xk07i3TutPWC8NDWdVWuurzIKmLH8B8/eso5xFgtPZgqBsZnr
etCFFD6Rr5QNm4ix8r3FeBmutJjBNJgYFf/Ox5e4uXJatbr/eyep5wY4NShCvrtN
HLt9N/k9XsyjV1KCzabGZR4CMj9UEHUlzxqPPKFxUxp4wTOY8BUQptdhyEKTQM6q
eEjHXPJUxl5pTFo/P2PA+38fTQYa6rjdRNucHT2Ga7H+RKh8BNWVXuR82y3Kcul8
8S58tM4wVIFddH8slGwOb2jDQxo0qHqLi9NQSuMIX/cBnMcv1sihtLO/qhU1wXQ5
rOl7D7HjKUYn8tGj+too8to+LOlkaS3s6vZGn0T/Zt7ZzfxoyrAT+2gDaiDXusvU
SKcPm7Qw+t70s8qVdyS798L5kv9FVtMBWB8MEFE2IbH4MVkcCycCcwHiJXV3Bnnv
oUUDvL8Me4G3OG7WYZODjwMc9PAbu6i/ADHjzsFC+CpPZuAdR0tB4MKXoTowfsjY
wGd9mVyEIy3R7Fw9NoYDy4OKkbvWgSSDLXXD1Bf6cV1cH9zcVsigcMiLdWaNgiCk
QeJjXFQ17YF3uI9TIz6gv4mYVU0/9vcwu49wIAH04Xi1vLsltVLPm16ArCVQIwih
2CyVRelnedQNmq0xTTE9Wft12clt7Fnm0RqNWgxHGRKTmC6FhfScmD8uNiD2n7yj
1r92H9TYQsu0ehFNls8nPrEtEhHAP6PD+zg4zHSCASBqq0qmMofxRcDS6f3m3tXK
mDYjy0HB6b3TohKVObfDBIvxerH6etkSO70eoQLow5drOHh1clKR2/pvIkfCzihA
+CmyaFM52smEBdoIpFESZlKUgXAhU4Ar6Vio2iJN4TGapWctS7nmAmeKRP68Hkqh
nus50HB8ZyPPIuDI2F7a9zEmAu94d3SH7Nf/MKFf2dCsEGvTDL6SXJL51s+nLCH8
rHBW9fOckAxtpzvrSzJBcNQDKLc+IUSf5DWsGYMDqTuYBL/pnT90Qvq/NjaJZ5r9
ICCQWGM46Ua4D3an+dYruWU9+akeKonBmhOasrOBNG9++MO/6ReuhksmoScT5PNQ
j8lGUidGNASrEFG47tD3/Y+6jcrZT0speoCG7j5L4AKpbhs/U1ckFJMCRZs1GPNy
B1qKEvW48J3sxsi62UsbElVQhN62BSMz6CeH9R7YQ7e7GVtyAoRFyW8MpMItWOAi
crmmFJJe8mcuLeX4T+fU3gh9BhMYEWY+hhAbotFcB0Cj3cdpk+wxddMYil2yjvwQ
FCLwLQiMzm8i+GGMeBqqHk906sDRKJ8UkYwg3l5xzivNJrDSx2ucK28EGBWn6LrU
/Bv9zd/0LyBDWPX2EEVYaGHJTiBn2JgE9ek0dFQiWZpXkUHxVEg5KdaKBnhmtaLq
J0ZfGISl9vfwIBZw0JdD74aXMn8XXP7g5eCMR1vO//jK+OLDLoVoUR6kDLyipgnp
YJd4/pbQK498iDoDdd0T8ejxcC2Z+StLxrAjx+ckIhcWw7pqAm5u2HAEiekZJxn5
ILPSphCF6JW6dvryfb2EonxZ7dVMvf1w7baAeJikm5gl42Y6BnFObQjohSRDDNy2
S0F4j/XRB+dWK/14ZGQ42G1ch6Tvs+ut5NcUBP5nbCwl0s/U4CnRloVm2ctMz8aw
tgfmLOoDi43Cmk6hk7PbNXhWDnZLtjMDACLddwKgOqyGdrVopflwlZJbvMR943tn
NZ9asFMNNfrToaj9nMGrF2EVNgnPl0bpsQD8VMd25veaoeqQFJ9fPl/lpu3OE6xr
gECOlmquMREAaESu/af2+SNhjpqy7srPY8mtyEzXv+NeNdXrRzYCT8ttR5k7s4C4
ImzFxezrULotDT13olm//UcVq6+IQnVpF47vaSdSL3S7kzucfjieaT92QCTx0UIe
p0cCvesoM40Lqd1BjxB7pKPIeWrUu7d/zjFKUnyd7znCZOxGpum31XHnfYSewRmw
W7t4JR/Wuyzz8x7/UhQRPgH69gZx5oOH+2BMICoVN3vbx2j3SSjXoFdz1YH+NhUy
TWGNt0No9EyAeO5HKHVztpYiCUeo+dOrTLMx8PsL5Ifn5vPCfPhz6eSABOzoRxt1
fKudNrsbTcd3Hp8bph0BoRtMX0bhRFMcGuBUilBYOg9m+VzAaAO0bEbRdBnt+EB0
VZFyp26Srak7QxF0sWVKpdLa32Mb0/8BW8f2e3IpwQAt1BzMR2FyeaXY/OW/sQIr
ssAU+INFzamaiWvsuVd2MSoDFXjtyISwDwkiE8+W5oygx3UjdVuNGXXyrOAstp83
ZuhM1kR55foG7tThQTCrg17vaM8cziOU4WiT5tIlob3YtprLBo+iIX8UEU+tOjAl
Wr4h6PyDu8vQ8QFuQzeCTrlCMK9QWU5+zw68cunMU5n4gftjDA8D/7FHHw5+HIFZ
GibVHfbtsrtS7dCw3WqI7BslBy8RA8XYl6JBp6rtv4vJv4iGlIYMnRxlnJURcuNn
+2QKpOka6XtNuTscIqSLoaMEUYFpnBgp3HyBOgda6XV92sdf8UZRcCPjI1U+shcw
+Nyn8CR0R0LhNTEUFhxLhPTnFiIfF0vRR0KCvlMTBPnm11EFEprGrYodFoF8wZ5k
U1HoamM3+A9CqoIEAGDXWqozks/IZaxboL5tfS2iBLjuduJMxuU+JgadbL4tIvnZ
LkLufSKCoALZqrjG03beRov7UPQDW+08z/ozdi6SJCm5YcxKkCrIp54YlyBhSdL3
QzJ9vdoBe7JZCfve0xq5EllnrxMHldA/XvLk7WeJy/NWgqBp6QG40Abvfqfn39wv
Vlii2e7zBVeyrGdKlKCl7BrZogm1LBw64HD/5FeB/i7yGldk4Bz4jYXuU5+dQKHJ
LlXEqUxTyxpuMsFdKAO/y085no9B55439nNm2qxdBrdFVasIXeVqpFOzcwG4bS2q
/gG05xDzIk2xVGq1OkJk6K8v8PSvCs1xOT379wQMpv9yKthYCt796pyP2hGwDW2/
WU8qQImA0QQvsEJwbgep8fPnEs0swKLRcL7vr5jOVgF5xb8ljSV2OFmMowB9JJaJ
i1+FMzyF5MHGxmbujJbSdfsNTPlJZwhbaEtwyPX/hM3laD7vryVElmISHu4hHXg2
xrCUoY5zJRuthG3ZhnlMxCoWn4KZvxOWm7/MPzuTJ3eEjyZaSxtHo0S2us8qZyjh
IyzXk62M/db69p0999/+jtGinn6wMyLRPlq2o9Jm4NUI3W9pROzMFR8bhHxe3P+e
m6ePgk4p1xcNihKdBQBrCdEeoVGGg5SzObeyG2XAAkRVjGdWumh4HnfHPAGNwmO7
DFpm7F9NXMS4aJ9ZY0gFyYAogLUUVEE69YNaXjx4p/wGsPzR13To7ZSwDYhJqKcQ
xM05xGIsCi4UI/oD9KxuL1+UN7fkq7/Hk/n2qGPD4dyzj30VzvAiJgtkqC0i8qAR
R0H976aG8LxVtn6DGeZEOpq0HZ1qSvyn71G+nWbono2JRJBveQHWTRwYIbl9nO17
J1VTUwlyZ3LhVF4J3H2QaveMfXSdt6zZFTlVXTA6eMNercdMwA3CM2sgHuhUdAEz
hfatT0g6v5h6k+MGZdqlJ6occhb6Usk9kX7sVGtpmQUroW+MixR48c7q8Cp2U/3u
fm9Su15FBVyAA2tCYDeypuvPl3PMOmfOH0N+cRtCIpmXCSMnrzHGvhDNTKfcIj+s
H4Meg3+ut3ZNtrKK943jTToxrDQKapAgS6R5i4epujVQLT5DhUDIzxOj2mcMmRJY
2bSzlHLeZdg68FwvNbGmxghd5e+qmxndrc+FpwtvWk6jC1lr8NccivvXnGOCEk8D
MevVX3WHrFoPb/2KuRqGFls/3QavpYiQIwd/iVE+dLKQVu7lOVrBwoajGO4mW00Y
SfEwMF1kEf1F3yH1mo7xmQc9Gh628wYZSzVm68hcRF8xwMA9MMLJel2f6I2yb7oe
Bdzex12VDzQTbjazsNaTR3Wm0EVWnabTMWa8SoAyMVZ7PDLEEH1YDWK0chz2zkPU
+sGEPZPPX5o1hu4JUjXQwIfUdRfYRlT7HTJ2b0X9+P9lwhugHCv8OGGi7zSMq3/O
LucwqeQPTXHH0/ITWnyMrH680sYQ5iudRW6PtvKFVhpkVYMx/hiGOngyeCmFFnfq
8kOdzOVwNkR5s7NqNpxIJgUv/Zes5mHItuHbQGNySgOpY7rbQTUHDZ6mykkHphAT
bCKhw5ATldFDw+oKnKI7+6UDSbIRpnUPVme2+Jn1PtJwkSs+mW2Y/ojXI7oToozi
3vTGOI9+jiZKBEoDCaJkOByV8TBvrwBDQqwMOHyGOLE2+I+Dvry2GcRrb6jk8aU/
HzWSAzyPs31hlmmd5/1BwS+hXtjTB70BzuU7KRrsSTKzWFyUTZD63OMyoicm3jMd
5s4Z6Rh6EtSJAI5v7fly7cp5jFrGZ6jmylYAme6F9uv0+tujSJ9sApm4Uy/sqPr1
xA/FzKHdTXQRQ07hJnQ+j8U1hAiBNm89Rvy6GKEXaIg6p+RWqsODcoqtm2V3Kypx
DkTQYLADNel5pHMh4rXsPTIP4GnX3ShpBjcZYJoKjXstm+nqhH0Dl8hO+TUvAtzr
jmxkSq3aBa142SmgTK5zpncdeiorxu0f42KsWRV/Y1Z+c3tSqBrIh/8gslWiXFdZ
RHLldZL7jD1QSm2rSurwD4LwYaOeNSYY4kVgMsfGVLri9i8xWKE9OwMQsO4ioFrF
uecxIeOc/tMflqkABffD6bPeELF1KsHoJEZlml1qDWj1zqNttw1VN4BGVPAZDBck
/0fAwtgJAgGa3VNHkqv8SjrpV6FSXgUEb3Kj4OGboKFX+pxPK5kYO+awRRRFzGOg
VUFuCdbnebiPaZBXWiLpCSZRSO3VDc/tKuvNWMLi4mfZoWu8I8CCDn/kXfswF88u
a55SFbUm4mb/KuiyijOudouDQaqVM3x621SFMnRkKlRSOptQFGmn9lJMgdBkOzen
lt5DUpBBIAO0lP7oIIW9zF/LKwElN1hWvc3nqwPcQCq/A378RdMOg/qnczmq/Gap
F4G4rAVnjRqz1NE0FYS6PIkaQLvmHbPUBTMrNEcQpus+EKJD1YpOi5DHHEb14Fri
P7Hn3ws+K961qstf+A5RspYRCDcEzokMaU2Y4E1SaagEHu5t3t6+hDadgddNsWrR
ZqTT+/WkEoLc/BBUIn3cR6ICUKVCDv3eCI4WeKXlec4I+CZQLoCj6s5UZU0/tBHO
Orsuvu9GHLouSFnctmNKvxpe9vf67EDILtq+hciN+wiXMR+Umiy6zPRx4OMuyll7
oIIGnIu7zJXbRPYzOClCzIIx9qJRDArM75JysQaLuc2takP7cfL4cuUIyKVm7r3a
H8aVJiPEQ3L6rlW9MS67m7i1MQ1IX9CL5jJ7UXcMsgd7uzi3ePPZvbOWvTVOhzMX
aE9xqLLd0ZchVPNRhUOR6tqOZirEcDhno1TAVorE7lO+4N/us30+7caLeWnrBa0y
dUgfjqepPkSiq0vOkXNd2tHIlhczC/DnqMRJ/TyQkCt9rammLk7YyYnHpxHJVvQY
NJTS6edN+4O19UrKfQcS0NxZwHZB5AubjFeJWIGzjL4fAk0nwUlNqjZ+jBH/YFH/
va3x73elRWccvK3ausH+xRR2GsKt654AtQUQ2pbkIefXHS50109ZZC0M9Cnm7uVd
rRq73aOYp2CT33kwyxhb6OU/uUMRipSp7uSxzOU5uj/XJGuH+N/N7yz547he2yUq
HuMPgO+LsTvhOMKbuUDkHf4G2+ANsMonyRYlTv+/i0fomeY2ceIwbhsNw/K1l4DI
k10onFUImmcpzfQ44dllRoiHr1URGY6JHWQa7XcQyZrpmY6Z4goQq2CXwu8XXhVY
HcBWcaKoJVi0vgH/m1FFx3qUC/6UOzLhjhz1XDDiUQLkdxW6gnycZGrsAY78W5FG
v3g8XYLHxwL83v+1Q6rEmO9pQKezvaeDERMVccofQYGsSFPiBuOnc30jPnCC4Pg8
uDBBB91wYFk12cWre+U4axDLUkwZ93uFvNAuD0pW19ZpU4pIu0XfLyP1eaO6Ma5l
EJJduCYvQMELudgVyy0QZpNt4v8e26PLHiUZLppe+Vv6kSEEhPmc0lvoa84rw1sW
iUcEzat3sytScYJH9B8k7rzdgYzEorkYKq4D4w4pM80wc8M+/YZz+OWZhyfGeLw6
yhYmfYTfJ8WpiynZnnMGfXB7+0jLVC1J7z4mnAJ3qDj+C+qp+3Z5j/J3QyLD1DKV
FM9+huvzz2uQRnp27QMJy/I2vPnITLkTswt3IUUy1VmedGjY2uzm1b5axKT2KjOQ
bFFct8mCvwXAAh8y1meuIpiLAr7llmC8VfcYeRGIJUSIklhubjXqtyeH/IBwxDCg
G7b7r9NcnTyGxB0TTlMDOBYEKgk8Xz4zdS396u8niPEdfO4c+WdwHHX9j0eXm0g5
3c9MQeb2jzcjjMEAASZtVDlDNu9aSAYWCCLQJMMNnoIuzm5bNHS8761BdMG0/9Re
xEq4mubJYIZ0xOAgpi161EJ3UsMafn7Q6Ef3MZlUTy46ShSzqdHZU5QPkaXnTJWU
oO2p0EbFrK/ny3KD5lAep97TA8IY/dE+heOHcyWbvkpSQhvOR2zmwGI/Wwny1Ro5
E+rYLdza36uurAu+NDmdx2Cg3MxIY2CPOdLw4IQQDySRcRpoGTLg+BkzqMpUZHP8
cAy2OgoJCrR37aZS0Kss1ktCQPBiIwEY3KySch6ez9i5QqG7Gcl0A04OkzTrmqPl
t8KA/I1hShQ7aZ1OBUnAkLIeYz/WIOjk2gyjXWIDxbZWExE+04R+IA5wn0y3lL0j
hYbJpR786QMM9R3PjrLp+HRNg5ltmm8daofu0KpNR2tDRbdT+k4OnEd83ZjHy6Qi
/edBWbsrYR+x46ML+3tolEYHoNfq30RzfkxYjr+O7xlcZadbGW9INmR+xy1Ga05l
iABb7YMJh+bg4qs87hrad4T4IQtrhhJgYj6i4iL44ohjJGNGOasH7V6i6fcBgFI/
zZlw62lhh3ovtJi0YVo8nt6EhkWDWVdSWWen2Boiaf93/pxnyJTb00oFooeKYRAt
ez54hSeaSQCJ5xyD+BNwwQCsFO6JmPVdOcjh9eoA3mHcG8EB8mPJ/Lt5RDMBzhf6
KYRUW+I7aimU2PWQHwDr9JKtA23O0V3c75t4O7VC+h+xDbTyPP3nPhtHrJZhKTT7
cECZY9OIuz5Aajwt+shNdnc6ucwC0Xn37rFwg+Bv6oXVC9u1tH8ev6cVWETL6QIq
F19EislUjNKc8VM9P/uaFK2jn2Lg6SOMJImmwYfgZ+/7m71VWtbS/S+Z8RTbWZVv
KTGYTq382cpzNaJtXBGGbyptZHhTMaN6kfYCdOBNWQlDQBMkXKsufvxxTq93C0S3
xOuVs1fKgnczxZMlgc44cUSVHuh/q09oGgmPzQO00Dn9wFyVKZTLnpcGw0g+Dx4J
tDXaXceH3PGa9qx+g93QskVTg+m24TycgPo0YcFASNLpJEtPKY5+DEM12/NAdS6Q
WQg3hktrBotEzzpqAPtjWe42l+JNfWixFY8nzQg8DQwL9rwIira+cMHi0DJIqQEl
HrmVkGH7qyokVq3u3g0/wmpbqKP4bmpbsL3SvDluYbbwyIMH4LGxitQCcjYvqGS6
YSakRZ26C1SJxNuk2mPD/WKXLiJ4Sg0rzmfShBGW7svvSOCtEcHfwZxAWwJxKSI+
4gUQJtrpaHtlJoD7oKdQGc0Pbd79AK8wllrQ3QhcSVYLPVdq/ACMH1wvKy5ay0hc
5RMhl4/RFQp8Zsvn3Ra4rgc7L9y8agDYfF8e52RjMj4f/wR/gWGi+EbirmftK/bv
lIoXcNPNPxloCzN1qodo7ldWTAAlGGpegTW/BLVIPaQ3BsV3OvX/oYS0a6svv8+y
FRq8KpB9uI7OU6amo7I2dKR+WyIdY0mq8WNiLtIQ4ZrUyrVV1Y+04eU9NDXiiobQ
5A5bDUNhmBBa2X9pENw60ZmgjEnp/k5IlxsUCORgICRZZW2aH5A16PO0x/cYxc8V
zGR/s23Dxx9J/R9jufc0yHBDoYOegUfYXOH7NdEX8NPLy3f4B0wOoIILBGDsJRxN
3s/UYDwsKUfANRuPwFIQkyRz4Up4ho6Phd83yk5Adgv77yZOMmK5zojd0aFjXkXF
i68YpCQOFmeYNdg44uDKy8cpjfJgzkhs/4qYava1taQLQYou1Ngg9zLoAcgDzA8I
0bdiXzEdDFDz48v/y5GMgR4MFTvdBFsPQA4K0vtxh+4PaiCYGJaKwwe133aU/c+I
vKfLKXUFCSa5mk4QbM3j50SqJiHsgQ5eCnkoAcB5PZse8K0vxJzO/5NbLDZ772zY
9OZlHrbe7U1vY+DZa9brUj30xndREmyFgQj9EHEgmQrvEfV8mKF639A+e7+Dv/8Q
7DTIznSFlcdlozfYwZm9qi6N/xHvDtXKZNSKl3ZiyXDS70pMwaAOsCGrgJuzp/yg
28twb5zsdjKGtobsJVTQTjw5yiqWJGu2Y63hpHxmWUTi1g++PDPE2Soxm7tabYkM
3YIExln9SJ0upEZPyCFZEzdZRh+ad22/21s8zJJM1NjLbWTFCREg+73T6yKWyrMt
AW9LY+mVDQg3k5YTkuSznhAbiX/JvDcjBgqTn4S2HtVUOrpl5wXflhgXkNZcbuyl
ZG7Cgwyc7fDSgQ1CTVeyD1DpqLKeANuLsFozk+qA1QtTW0gzqgF8d1rMpBeav67B
HAk9eOGJctMgWd/QMzAatzKnpNJn1I6vD7/q3oYYZxeasYjEMGyj0wk2Wy/Tn6Vp
wil+BJ5/uyj5R2GCyF/Xipkbx/HdW4pmhviWEtoOE62DPCp6V87Wvi8AmLKa9Q9I
DbgkUEQsZOfwDnkmcSbuIz4a9+CbW6Ba/mNuS+rFj5o8w1TA6n6DBIQlsrc2yNDX
mXP5sZc55/guTcMRbNNuOt9J7QHEoE5aJUKw8Tx79vD+X8rf8T/Peb7orjlmHfRW
RtdqLjY92T5QrJQ8lhlmsl2Wa8lXpvbQ6wmF6bqIROtwmyt3AXlr7saOZxOU8Rf+
Rl5zQgXDV/4vc/Di2bArgcjbfadmGbHLK68d+eTidNbWyunPJ5Vn7Hq6PtWXskGy
Nqr7okPjnCwOdJDQ5urIp/pZZCcUfLoKL0mQg0N3YJjtkCBwLCte7evwHm/gnsb0
PWfk8+tPabppCxCjANxFLTcKTm/orAei+BR4lS/wbf+lUL3gUdYiRWXwCVHeYfhu
MZcad6kj3/cCzpvfowMQYVhFgRJNEgqj4lnOm9xeIhhxJ0kBeBTTK0JeeIeIYlFp
nX2+AJgaO84je24T/6uL6VxYbu/w3c1cZQw7mj4eMiFzNKyX1MpKABAnd2m4lfUX
9DnCeDTpKM4518m2XtqprCFGlOh8XRAIFzSDqZHJbOzvnAfpC22YzyUf3n7KA1iG
+3QAzy9dGGoFdaM6B7LCgVl8jYXI78Kyz3ST880AOmU6wBUHBjTkQJfOcKA9H0ky
zM0LsKGxMI38B+WjgBY7VgjD0Z4tuH9V/kGJmqwuim8aKwDd0pkNyyr41Jlhvms8
UPB/g1hTXXd0mcZPjepU3Nem8GBpBE7ltPrjkC3iAe5YLswqqJS1dPMykaL9/AyS
9jJNz4xIJjVznct67tXV2BvIVdeJkSYRwM9JKwwl07kN3FruTK9ySgH6tJqBoobv
ksRJc1+g0PQ/U4OoqC8Ta4vbLhRA+f3SroJWz1fAwQjPCmQ54Vd06zvUOaWhuJrM
3gg3uB5HVqL59y2n3GR2x3xJMzTi5mfN8oy7eOIvAhMPzNrZajEhpj5LvEyf3kwO
Xm6Y2EMrKI7Q5YSs7jfgAHlO7Cy36cmaMO7EAysE9dkP0CdzeYzW8PWQ7SgNcmzE
XJo/b/saVY9bZDPmog3yNEUoqMfMy8/fo6jV5k0G9u0ID9Ghh3lwMPn5MEcjX38S
ikjpydA/HhUN9TshUVMs79JzcuEFjvvmSRl/LXfq5G3Pf7kxvabM1Z//xCwVNOY7
P2KfB/ywvB/YxC2PCaCwMrHfciz65EcVcmF8WJWEIG3hXYBFTEWwDOlqHGPSK8Jb
/+dyvL2S3Df+wlhpdaQ+C8VVZcK7vUhATaOeQgfc+qVNcjV3sTeUCkdkR3+sPWpp
vzFQhZknDf4fKZMckSnXcv6wN3aE1hLm84z0qGj7cjdCoD4FfL8zqktxhgeC1+w5
zr1uR/IG9PiYc6qz3s1KnO2re5iGag4B8EATY6eRIXtDpKIxS9WnQMukLCQcldRI
1cSR2UjL3bm/QxT9Zov7q3NkN7LOj+CnEwwgovanGa9UpftvOy0P9RxzLzMzClKV
0K5FK0a6J7VvjQ8opiAQoLrIVIUQFsB77KKbnkxwKITGH6bck1GoD8jFDqJH5pD3
wieXaUSMxYvLfVCcqjvYvVybdBIjZGiMHqaqAr2v2Un9Mn+xtL66JWJuPV8qVCEi
3SejCa1wea9mD59RWYNFG0K6yuFK4u1Z2NrbiLPO/dzmiOz16iuq98WzCJn7NHjh
dDybE49RnNDTWOOlvgpYSxDEerrPq5r2efkbqJlx0d7xy8QXL6gaIewkmq+Sx9YB
QeNWGR/ULwUMI4fAELs8nPZf4r4qELDZmwHcx5pZaUbRxBAWN2q/tFAkbLdURuyi
rD7kvAqxRRBngk/LgecsoNnfk9700tYsBcoKEEpKLKrRihoGkjO0jwygkEU0YbG6
O3mWB9vEgBbSyqBQD4uaVWElr3/6GOY6rapWtySF75y2+Fm2qlWd4P01xlwrHigw
0rGzth2DGbr3libfvZwBRssudr6lulRWh9Gk3In7IBs0XaMS2/uehn7vmcCy3kdw
GHI9hdh3jrJlLtQaIMa1qTOEkorhs+MsJjGgq8/iZDqY46fiDEoJ4L9LGqbbDQ3e
mRaWTZQTpw1cdVBOorCuUTMBwEeb3ZW+Y29YLjTWR0I4Isqh6/DQmeQ/53Qp9V9J
1PZXKKdRTHXGTXAtC3F0gC7kYdRgCoAh5sHkVUv4KIXE+mnfNfDVUUFcZXO+DIVo
E0GxTIOgTFLmgApyVl7VhLCzBqMQ3mSJTp9EV7B5iINtSK1pWqQQ6Gdy4kLrCKq2
cDPF5Xge8ww43CVfCnvJ6EjXBxzFz9yc2kgDOjstoB4ZohtmFGhY0Tx8fTtSQLJG
bXTp8NDe/JDOSmBrj2EwQS3MSYthttf0PJCtZ4crcM1BDped6zFgNXrBlvmKOM75
FCWPQKPcfP9FvJgqGnKsWoxNlRnjXjl/JH+UThWXCxdMHzMZLcl43Ylt0ub0IsrC
0Eb/8vcOqB+IuycNEd9qWUkZGNeBNJlDInY2yrbRRBEPAnsEfDKEivTvoQBQFShP
72vyZ/XuseJP3SWVVaE+H2DMgACUPhX+5Y7aD/FUmGw6poRfQun761xAlfb+O2BZ
zazyKsc2leadAZUnkZJeZhaMwZakkzs+kaN5jR+fUT+iBsAWsP6in4vLf3o3wEpg
93GzKR8MQCeOW0VfTl6r80oUQ2QHuND8XzGWo14Nr9GIASmAPIgVHXnmW4XxLu9Z
p6Qio+h0skBGhAZyF5HscD9E1BrCkfDrcpFpskPcG8QaZic4vBc/A4jc/ehDSYVe
blRXZnry6bSIwM2ftpNtk7yBtlnatpmYOLyNeI2gmP2p2VasZX2hUlBO4ZSv9CyD
LcUFNbMIXz4nCpNQ9utnJ6dnAwmWnhbys9He0u6v5HbD2NAqEBHDnPbDGrNNU/HC
HTJ15JDtOzDgUrTcSkuCSCSp25C0YgsmdlwCwADUU+qoK/kJBq67XECvYWDIgpSN
wUSMNI/DLI8slcQKDh9aZDzFNtlApgBlQ18XC6132r4dxqibwSfuiMNQuJ9MPbfK
j9HyHLQZvYEUQ1OKqLV5rb8/TQoc6JndaNcR6E2yfCCL/YHNR26Ggei7tOKXCJ95
GcbP7b+Bj5NunFyFMKjSLoZcTaOQJhk/rCUDCbdeacLZysX7PyVd/Ywk55mriSKM
evGOp35rMaxcZ31ireeyBzIRgnULx8IJiGtRCTJAq4ZNmpi5b1TAqFrUQJOgjPQ9
yNvKztERemRua7jU6zQAeE0Umk7Sb/CU5lUQ3Au4irGQUw+JA/BmMW+Lz7dJTZg6
s8Tzp+NIiiPV3yQtd+JM31K3BIwNLb4Tool5Uaele6vSsivjAwRRyHPk4ANTSCau
BNo7K6BcSMTP7zj4wJ/0QPzTJqCUtOw8E6jKZnRYUHsQZtgpdTo4WVJzCfjAPT8y
mhqxy3xiWIYgNTO8sHZBEdgj7HOuF/j4rHeaasCEvArqUaOZS08wYxJi4uCbW0s0
BChRDf0OX0gG9L7zGl1XvEXNYPX6fJukhuJ3SKlpqDGh5+2095hc6sZ9h+S0Duui
qmdjkXiQ8C13Tr+cEVps6RHO9/59KTNfLLEp033b4IqIZCG1PoZsY72TLgbNE1K/
K5VgjQzcO3tz8mfeDLwl2TLC7CJD3cAHVahaH96v6JdlaVSk+hw/HhsEp8X1BPtr
bzdncRTrds1l/5uuH21/Y0BrXPtPRi3i72WpqlLMBSnAGYB9cktEW5uOi4vD4bLh
0G6z2lE2+zz4ZQ7c/ZqTqkEO0uNGA1/BSPYK8Uq7l5krZM70hznVvkpP9RuouDku
MoD7zdSh6rjfj95QDfnMhBRRcmtacq4lJDvgidffpWt5EUFbQqzufyFQGKjS4OB9
ESzqc1oXSNTuCoFQfdCwrC/5rVU9goOx7htnecDUDfTN+nT42nmtdATSgSymEXID
lDrVvzqFcQQK0JW/2vepS8Tkf8wIk2I4QNB9uUmSSvmeFGF9EPpKqIYIy7ISrDfL
cO51ZkWsmbP7RHjK5urINKmhV/xl57t9xuGmHwr8riZ9HKYaKRegv1HjBzUJyEoF
XbN+9QQQJQ6Y/afOaGx0W1wufUl8kbgBNaFTMhDn7jU31HeB33pxE3VxkyWQ5wAo
vqObg+mnKoiHNBr6dB2fS1Rm+qCUdA/8g5HIa+DNzKiaCZRHD/y8VQ9nsYyuGeqR
3IqtS1m5SwaahhBT5ljKHrQ6RCgdQTDIMgcFIE0DBGTl89qTppc8bUVhczZMuT9w
5NhWMkm2Srr/tqJHVJ85n+A7x2Kss3WBoWJpRqERElgZaxOx2/aJ+ibdYEO1Fxzz
vgQ7fcHCV07BliaKzxvYNQ7u4CNzB8J417MtkjeoiGTIT4O2jJysFVJK9F8d+A3W
/U0y/7gAMsVNFgeJ5mkrASdnBrs5VGWCiwFVVfUMIc9V9yh3D0OBWDPwAYa7WuAP
nzXatQjin4JX1I4Y7w3mTaDhR7QDv20cBXPnYgEa5Qk3zixxjPtEImiHSrq7TYUq
MzKiEEKJ2p1lEb131z4na/zDp0yY9LOieRDhVbNt9A5UFUhmYAoogsV7jEMDOkB1
WCP4jC9fFNgP6FWWzipIymx98p08xxYCCSL2hszAIzWUqRsUJZl0mIC1a1ArZHE6
lU5iv6ljeWeldZyTShF3Q8ewHblOz7wWzVkJJVGDidxsh/owU/kCPD+OUTRUyVyf
YDnK/SSL3Tc8W3GxEMF8Lccb5dlxXYnY8sf39VdpWH0KkTTlz4FAUac8FDfc7FqX
EMvBXc/DbbtaS/kLhVWiIrOcumBm1VQqFQlCZCP+OKqLBwoHags95OjlH5i5Ixre
K1uxb3uO+3POFBZ4dURaypdN/CudPHRLF1Ak+9RecB++/q2EcH6gJBv1lwaG05P+
Yb8gMVv9DPE+y5talZIhjBZOq/Gqm3RQ4Mdst3k6sxBEDZrdMB+ARSisbpuEywQ2
KAFY2s+ko5UdtazH4j5l+dolz0iy9vCY59NWyMw1sJpJtfv4GYVfRBD4M5uXgKs9
8kP4EmADk2p+UlpHrnpHqTium+/ZOLnZmlsMgDLZwDbxF84/clE+9Kn0bMtKi3YB
7DFx5LLe5X5AHeIYfMlfEg6qcdw51Y91g9/IZfSzUEf9OHWOJ1UFZ1LaKL3szj9Q
XiC/GlHg8jYdKbPKUudIEswGwZIH6KM45LrQwLLpvUphXwtxVtZNYQrAumAsgMZN
nYkVZlYC7wsstn0DQ2d9laD3A+HybolHCuHjZpA5iZkL9BUAiotBa4vgOccre3pJ
7tG1NQHywUw0ee8pTZmozBnPs/c+uZX1yY0pbP1WVLixRc/rS6qpEmsDbm15bgxW
hinx4V0k8ZOqdCRs9z3pT0tg/Xj0ya4Fx3OcaqTi23ag5RCOAr7tXgGh1FBKkFXl
CuobOrMLAr2fhc2vZZA1GsAkFw99QfzxjU5H6/ryR7Nhi5vtacRtrd/Tn8uq5/cd
mD0LpbR4mYECg6fbtjxiJg2u3Hjt5zoDJgtW1SV6DbOJVgjQ6kKXEEBlwHSSSMzZ
l9gZ0SxHt80aKYE8SiTIE/za1qjyyf2FKpAhTDyZEX/UJnCeWOLA13POjwJ+UK/q
yNoEiwpmZlipbfWvq0xbQLbIzLWqyHvVRgziZmZnSD0U+ZxUFVCHuGkbSjL449PH
ixOLGexHl1pMyE5emJb2+3y60fobH4hq35EZCk3/Ood7YM4vaWODhgLfYqSQQimM
371fQZ1l+Ai6BNIrHmjs1rHOP88kn9nH6x1reiJHS8XoJwm+vKkbfUJyj06wlgUY
e2Ojar4E5IHz4BmuSMA5+2y44s3Q6CD056CTmy2sd0dpWWUamC4uAEjw0er88MuI
fB+ZyLUFBVE0uBfthwE3bXQK4FUjNWU1GsobsJ6dPO+wKq4LuDnqJXfV6ICnxDVT
sKk4CZFIt0qK46C2U4HVCYUBlF2ra01Fi23mpLb5lTpnCsmXddAaqmzB8Ai9Fv3g
h9QEUgGeFTZuu7psK5k9pS9T2FV2nMyDMappmxHO4mr9HIqfzWTUSXc8ZtsqvS/F
1dW8q4h2QnxkL2Byx0ORWeCibuO+RqAlMWvzYn1aFkgiL2UMB6TRK2/xNrp54QiP
uLU66KN1qUNJpk9AliMNyWjfg55or0MCkNSKyOLtTnqmzGpMKihl4+OafQ63Xz4p
4QJyhswbRlMLyf5c6INvCCBS9FNUun2JbRWlsjLFzWTE/0hTCg9erL7C7kN/2/S2
L4hxCOz0WjW427lVj3uXM8IvBwO+2DVWcUGAe3uzg4pftGHuPdJWr3NKbCEsVPid
gKFKALIsKmM+/3Cnt7OyPqkpiJuORkJhjCoKjW0Go/xjtXwuWvBDOoijdfyJ1cay
bAtEO5ubp0Hpi/rFCyl5BTmQzpWo3L+P1j44odPi/nLaW7JQx2vlrItSfMKtesAk
HE+vl86R5dnZyUrwOqDTHooG62IxTn/09pUcp9TS4p7lU4UdgGYSf78LjZ1R+R/S
LnsWZDboCtLPhtOIOqlL9v/BUKaaS3HAybv6R48OipTyhh5vUw/CmYqbIKdm3HXc
vrvJdMCONqrQHLKOMCKGzfeiOjnBmOTngXWVrodFgLM//dmtvsGNzDdWj6kioGSA
1R69w2g8yar3TthTPNQdsVw1rOE/K61FfhOACVGViw+LNVJrR7BphVnP/0tGYr23
3xd3vDbjbKQHblWz2B/mzwvGf52uWgWnzyGMPhl64Gf6Vx0+YxaVs8LdaIzlxBRD
W7CGFPbJoycLfAZwfo/FvLkMJHJOujvUmejX6JSnyPgrD0b+HMmPE0YIqoZRMVpZ
Ht+iKBQyFV0uhprd9t5TB6hTRiCzlMEYF89PAjIs8muqt9VrPh6Ek7dTGLsfMjdw
cUbhqft8WBhvlT7bsAr9sQraby1826eCUdjPOYXMIiZyCLC2JXXBGL6TennTPqZw
Qv6eBpyPWCkwlWUZ/5T1tbQQ7PLUE/U21k5qSCWxsiP/hqe3gEUSXINCvE0KbCJM
ENHPVszS4qFO1DwEzo5c/DiM7CxvIKxKRbpHmk+PMofHVCvrNatBI99xEO9j1WJq
dRWs1yPn9wXPWoGeZF+7K+dcDar7tVOzkqfQpgWn8WVtorU/RRVimLkZw2F19pyt
ZKBWo3WoccgWJMbGnmiBs4mOnqopAFtaltKILr5q/La/4LCV0i+MsuCbYQ9dPY1H
64lSEykntDbedbqWWg/prfPMubR6tcjZty6LK4Nly44oBV3XHEVTr+RVqVQL1ziB
+B7eIQ09mWxhdVT85WwJrcsLmvWeYfx422x9tiSImZztOWBqeeXrPYGThJ85tU80
hKkf3a2Ci49H//323CXM45XzZ9O9I4HuZCezneYTU18zTLuRiDMirgAbAc2QWMAC
CRhk7eRMCAzghV/11bTLqDaaAA/JUjHHRrt0KYLfrajgwSLDCYD1HbSmoDqy100w
ZKJt5PEVJ6LYKmNf3xTcJUxLY06GLvwsyonrhPUPgFeoULvb7Fqr95Jqnr6dAYNk
bVif/cgJzMOfBUsZTXTiYLep6JQkspfu0NphNzvV2r1rXcDwOG/yLN7RghaAvUrA
AIjjdKrrFFuajHIo5EdZg6BRZ0FotCPyqlWpvRuXjoA5ag0XNCYwiU8Arm6KS+Fn
p9BA+RFfEx5W0wIrS1WWB0lSjxn/mlDVXjCa+g+TJE83+YMUcMPlKzVoB2mnpUoD
7VnqXiqbmIG+LhuRq+8t44pekRGMGgYo9COX0EcXKUSyENYuyrJOv8553HE/gCD8
2YFfpuMrOiFUElSaeY7D7bnnoSS/AkbGj+6GiWG4Dgi7hwY/p8WCF6VPweifXEH5
PEV9zOWHphuRvZQWDKah9iqUkZg4kAlpRtbB/376ooayMKDVxR8IVP69LT5unc96
syoojBBAgbPcqCEUglOfrzn1Jp3etnhRGtRHCPKX4r7UtxXDjX1yQBZRir1yL2Cq
Gmw+OalFa+LawuKN726ABtLMC/68Q4VpUHv3par3BqUzBef9syOM5ubdXONH7yU0
4GEEEpp8e6za/UtH5wH2m7+hxMUoZMz7FCHyIh4474OvpagTQeli4gLmoGB7Ernx
XTHxu3OJqC7341bj1hHOApwXZpeBE95Z5fTN16eLxQKpVx8SvcQ1TD+wHvsvHxat
hYOf2knf4kvi6BVZSWlLHsUxz046Ge4VxLvzokx7G/sZyzsjB6v689XOf0aqtyJT
8BFiOaxKlBPSDiNwLDOuaKEGXMEkXTL1uwGPNUFw3hFBbKOcN5fksII+9xwe+qOA
0o7CKme/+p69vczaQ5IcAP1jL3uyb3an31R9Tawq2FLhizGYFWzE9EvHDAGfZvy2
Bej5j1INYVvK94dbG4VbWCpmB4izCeqrMJlDSIKRuZwwhXyYO5lWb5Sgxs3FZb9h
WmoVoFg/a4WP6nc8esuuqZsdTJYvribZq5GokMf1bG7SeuLrewIzG71ifnS2zT8m
0h0IP90ccDz8SN83HFBAaPU8YfYitSZ04u/yyJEXtSIH72wFUNoVWnIh884A4PqV
Wuvp7Ce3VOdrqcpq0g+u3LW3VZP0Xj/PpXlEnEQ8zr4ma9jMkPVPZVaiieOBY2VV
TVzcHwB2UN4cI0akTWgA+eUOfU7m9poYTmqnpAnAUvW2QOTiMIhFLdJJrYVfCL78
y8eOTOrYgHvPVaolIgqpdeqGq9WgCF6Kw2MZ4SiWv9apL4rX/SYJkPl71bp0i4hZ
01rvorLe2Yl8aXl/Uq2mlQ8MpJVufp8dwtB1NgtJGFmGmuJVDCV6W1todEnhk9+I
A+wZCkxkxA8FlqKOzW2AsLbY9lykKft8AzIcPTjKSktpplbmbfBDEBHHIneh+VRv
82Z01t2j/+vP3u0CP8BVqgmI9kdsjv0C4i6f1Y7GSifACPY4WNSm5QRmjQe26eWw
lEjnE4RNBFGm7EY9cFRDzd5aQ+9ms+eb5hHkdnbYjfo0+4UXamiaYK8YOO2eu5Vt
TVhKGo8YrAesHb1kjBpThrlLkM37Jc3wyljEpq3/0KnLr0pkp+tbEQg5O91dRc9b
cdutv7WAyyCwktk5XtSwJMIaycfhvHfbYeXp3udZfH9rpIonE/fOnc1ciHkSYqzE
oC4ssvLREcjjaidRnBkCyIuSV1PkB3JOUQW4B+AuJTVN9kCMGOTvzKeuIvtpjO+I
UGNVFo3/JlyWrGXW2Ys3Y8zYPkCZrDHZRrMcdsTm3ZCG61u15JelJZv2mDSTSsiX
5siEW3R0eM6upyy3zufVv+wO+buf6U6UPE2q6tpSI9lDkNnTt16ztBrN2pTkmDD4
hmcigEiq1Vp7E1w8Qn4gwGqINe5TAMX5QxOCRZbug3I/eZTm8NV269FX5BJ+oNj8
LgAhyTYfrCB1aP8q7BMHc4cQdEmg+Wq1dOobjPBhZOuaXBt/iNgr8uxLvoHz2b8z
aDoHshmr1pkeJKq/YbSvPgc0R2ek/TxSls13fiBdhYLeodpRJJc1R206JaNzO22b
tbxx7jXt5S8wko0m5EirM25FK8LCj4jYL53oQJFrQ8EKxi9KdyDOk90J9NC2Uq6D
OpCmtLPtsGgfUPIXxRcBZD6aFQw0Nt0pRwQXNimd+PbLjt70ZCjnTeJfgTy3QGxS
2e8APA6CynYGy25XZ5tR7JXfSjrl6vIKZPbS5sSIWSm75xuzsNY4WNr039MgCWKn
SRy8BDX8smzxIYYiTSuuQKqBw2roaArMAo/jDpgBg3MgQ4YLo3ZScYmM32ZglwYz
/HPz8ZSzvo/1tQwaGVXSFgBkPiKsn1N5u25ix+tnJpZ4XgqPuGL9BX+HitfBZ2tS
EzscBX5aP1lET9arSlVPMZHjYe6ae5vDK46EVpOQAuw3afoKTTeMK4OqcorfEPBM
BrRgShkOtGe4R6kHTwW6FhlHXxsL/al27b8h1wvcaK0qWqzljzawTyYCcJgf4FZ/
ZchWpubiPbglvbhYlbbsmUA4Q4xsEOxpekARu8WmwbfysIr/d3eDtzKs8cX4C9OY
ftkGjY7pW32plU0miNVL2iUVpVOpZMmHU052i0hpChxUxR2+ki2Nw4E90Y1fNMeF
bs6ZjRhzAwzt395Jz0cnYDGPc7N3Khfhz2VVayEZjy7LgA3NybWSuQuFgm7h2Pw+
dWBAMGtbSJ12i5W03zfAtQqvMKd0zjnAZFO1E4dIy3NfNcaGkO+5l1oUQinwwUMr
G3YPcppMV5l3IKiQu6RCW9K4ijkFEz/h7SW159q1dMF1W5pgyAFsJY23WG0suE7f
KSka+oYcTxH8U7yACzMUFO+IlZdmIMZjNPJAe+NbuXcX+u48nLY1XLfaz9kPn4l1
QZOgvEC3gGx9WsAs+gLXcCQM9eMqnRQWmdfkDPhQFwXLgttIu0tBCARDV1HKd46K
NlKWD0b0vccOb2vdbOh9DWPMhuApXbUKJD4ZCgmNRk0AtBvpPksXNtyfg63eXLVO
QRBnD6Xpkc7sKZrymNLRfgjpOSta4Ij65Wmpa8wl3z87UXx8YYtwcIF62SAtzOdQ
XXw94pSC6m1tGiqptT9wG6x9ERmT0CltfhfE06oMd3Ru4aEAyNwadFEAHYm22sCP
FZhIVJkjRsHjpPRyqopqRtx3rpuAn7U+bcrPYbjN3ZbyJ5m3zIpIPrLCF1UAMXs9
JfTOp5OfJ9HQN43FO9899GCEqWqyfsXvCz5A05iQaB22UYT/PLNty/bT22J4WFH2
4pcjsbZhCqTcsKvy4SGhSKLmUeI9ZZixMbdGI9/YxLlcL+b9EvkJZqK/gF2dJw4b
9gJfplCREQuLpL2gkcIcFFfSNOw3Vhw6fj/wcqXadKaxVqHly0OgoswyPC5C6BsJ
eL0FLhWIpk1bmZjxrT7NexTzBV8Frxyis4oHkAwoL4Gg0nBoZruZvNOV1Bs3yRql
N+ySdMxuhVLfMAjnxgMz1cp35Mcb2KOg+ZkeKs8bp+pSA0DpVGxQxUmRf4XrToG5
U8yg5r01StIo8BAf0r6BBP71APt9qQajrjaHolv3RY+grpIR/lzvH58olQk+VZWf
bSxlTfoCExXvEgmzGvbPI6fGX7LQZbvuEHsvVh6rnaGPB1VVhT1Vl96zyGRkjKKo
8MnZ72/iEx++FeNwk0MJlE+KxLpY1xgt3TIQUaFZL5e/qQRTITIjyXpa7jt0NOwN
2lSVPs0e/FGtggTR44uYRlIjOjkYbAdg2waYMMjTPZTSoA1keltQMpKMKrfol3e8
ZXbu89safyKMRfeewg3xVzcoqlXRhws/OolRK0cJWu2bNT0I3fHmLzSBwuP+11gu
rxvGPvPdmui/Q4YZGzOFvcRzzTK8K024jAgddagyBpRmQ8Z6Iv0E102+xktxmA72
zr11MRueniVPTjPKs1IVZLOAG4+LGu4MKqw2ewamJgmmRlOg+PVhqGQLRV72NqDs
R0N1bWlqG6npgTiOL1tlqdW/7ma3ncWuUfKqsXvWRiKFXbLADP2xXlFj5H9m6jsk
FeeM817Zk+0Axok17adbpZdMWCPLmpIFMN0HWmgH3WSYIvAdZNlL6Cbpkr9R0ooJ
SD0enOEp7J9MgrQ5iFrA7c9mFSQ/y5EBDe1PqRTf55EBQlRi63wK/Cl9PhzGCHeK
HyfZrjbZctRoNEQDgb3n0CwLLV9HDif0eh0Lg1wlIRLT7o178alGfMFK4ZEKwwCv
YnFQcCVt8Gmvseyx3z4t6FTjWaDmzhaf95jHB82RNdVZLBYEgFWSJxNDIdWejYKx
vMlo+lXim8Tp4q5GXD8KuXnpp92mxCBoREn8rm2GpR3Qp3EjBbQlO9LOrRgusMPX
BhNi6azXK4R3P+mm95MTUu64zQAsT4MAqWoc4lU+Asz1orxEIws7r3OAgmmDpMad
H6CihWTc3LNG2ghe39FYkfl4TCyOW+/z07Jghl73aMD+eKiCfLaBcSPlG7jb2FnT
l79G8u3Nrr18SMg6dlcDfz30MFOGf7WAiJ4UFYIMKnp5KIe+wgB/s0RKkYmDLwDN
H1SW6TzOUCa3C7gBaqFJwD0Ipt1LZvpAD4GIVvFDVTnrIdvRwF0+Naw4NNiL/yWQ
6PJs3VtkM7an/gZrT0tEcgQYh3Q7SSRuxsDEeWN66fY9YwVrZVHCV5xb5KJ/IC+d
hkipISRnkoUObLjV07GdLUC/x0jKUXG73qhjeleea+jmZWFQBn7O0mA4NlLIWRzY
i69rFV9OMUZfcxoj6BklCb1skNHR43iGeHElZyS2yG/JdORkMh3LtGblCyxOzQ2v
I9b4frTRXx/pNuuJeBxOr/RYJMKaCS9MKkwCnejbcwON8/0Shar1xyqgpBU3Em3V
9yXHFVVZfeHJg1ruTckjHlnLHZCQ0RVjQgUEWouoxERkC8G4ogOzqPQd+G1ugcfK
hd/ZP/bS6y16AxwKlGgQ8dKMtGblmg+unMXCfQhqiZmvnf8r+8VuKM2CVBzGtBEo
Gep88a7mcF1X1GsKLSz4Av8Kx/O/PxbFpJ+avNYYuEFCMrDObro85evmatsOjpmA
Bl/dSVLYDpBEhhW8wcB+cmtWrEUNJv9ACkAIQdcSFLTMJDt0GXKMjEWJTD3Hut6w
7NcW3lT5FHhLw3AzfdKEHIz0nr3+yk0Dafc4bAJhRwRoBsxnCX2EqhNARyG9AsqL
AjZP+zU6GCAj6bxbuxiAeWKLmJ/SOAIJN/P9YtpzNOXXPJdg+KlwFLjFhws/KzIg
y9VToOM0gNcvGRZ2AzXJ5M69RFJ7JpzG5Blh0VCVL9MsRJZN/k2tk1cG8F7CR5jH
dwv4Di0ui0g5nq3mwFpoo2j7wwJein1DLtI07q7MeMkgag4ViLIt8HAiFIzgUu8m
CL2ehMOjTt539sUFjpCFCek0HUk061H2xCXR3tGPuzDKobtCDYb99QCkH2vWuYwq
MqCyrliGo3gxuISLc3P77tydmVRK6eVoK6k1G6fHTvdsNDoum56gt0mLQJyROPR9
PabchbFOMJ3tOUmIBQC48gXAo7y/FhUzqut2nEzsZOnedNpIZK1znqN3hyw8LIvL
C5SNOqPWaj61bXYsso/+U7Te6iwbXSMAUN5Z+cGaFiX65zIOptDOyCRvu2yV20EW
fE6/dop26dzbr0La+Li/wcq70/w0Pzyat+1qdBB9J3/cTkBSzUQ9qBxOgn6s2pG8
fE1wmtGqG4+LWUaQNRAJu7qTsuqxNUd1YFU3RObZ1gtDTrSyAsOAEHYEQfoXj+bR
PWf6KwiiPGXW/k9KM00IpH3WfjVp7srLbff87ZotpvjLT2gWAXgwjMY5zrJ7r7Kw
8sQoJUH9Dd5+spdHTE4/JGIPUXL+K5oj9eewONETq9z1+flPArcRt036Txi4KYNw
Lv+UkNibBckMCwzMV/8lZkA5JDqm4/8yE4qZ4geZWABXypGh9eyfK2dp6azy9520
gD5BPSCJIHANFNZZs/WCiXKuTkjc32Yohtqv17SH5TEy+TcpQ9Crxfo8oFjAw4Z4
ILgLx+gjQeGSiKHEjcI/rOcYppCqQnj+hWBFx5AAA4puMqTzQxnq9JjvrdIgDDzu
EAU4H/9XmHKaS0oZNVSOmcUXME3Z05/F3f4B1ihLUuDsGWYBFGQWcmMPUwldvdn9
AcdPsd1rprDhSbcJD+aCzyic8lEx05OY34WvPvUnYZ9ojNJXTltqKWvF/t8mt4QC
cxCvEcBGu2IQmuNeFAqYSJiuV5zaO1bmt8OK7m/OJFRChWqBtu1pwc57zyBtstKt
FLoGoimbYwxzaJrI0GoD8s8uF6Dlupprr6LK+CCW1mxCVkl88LCi3RTCoyApjSwh
XyXZT6aozT6KbpUqHtJn7rvN8OBTh9mZsnuaZGHITkSXRq6ITaiFWFy8NnD1kvB/
7sa7RlF4IOEb+aG51qqNGbpIg8BW3/vC8Wpimsn5bnykue3b3tOqv1R9kzAWz4fR
+YTRTLYSLvVmw9YVdKfT4tppb9rMKHC6rZkqXw6Gx94acYrXXSBc7kK6wynvldKP
HHpJn6KvC5JZRzrFSymXYr/8tLC1TZpmrSUpw4v98yjpYf+KyqRlp/0RFiqXdXZd
aXYeYKSb4R9ztLUX3ewZcVzlUiWhwzMhhnaPElZ91NuEYJn/Oum+NNhDl+1qm4P1
mKupWXVVAfYXyQXDDtarKZS1enuXOyzfGJzKpM7Rp9t14LlOGVXmiulUGEgasawe
btwSsxOUgMlG1mh2FmopcMPMvYWliwwN7UF8Oz0bErLw+I/xsvS81z9eUOgvgxPC
Sds5ZIu90gSXvFbdunFkR15yxwP+Ig8vpilzSLKoSxbHmTXi+zruOyB2HkcORSWo
imeV0AUjPtV0UDZ/rVvUysrAqsj1IA9/F7jquZwhjMtlGl1u6kntKLaTuCXcFHVQ
Oplesk1z3nQl7sP+0xwQMrsmhLnlRG9N+uDMPt/dAoTxnC9WvghaljurnFVyJyzl
2MB5S0K2inNrlO1aoB8d0wtgaz129nb2xi/X3bUlYd6UnKn8z4MyOt73Hn82fFQA
UPRjqV+H7yd2pb43rziB2+j0RjnzlABz5V8Qp6mFZAo7ZBH4hAqZXeqU/FS+nkWO
qkM9BOh/qUeacwGmnNYC0UiYfLdfxVS1OKmB+i9ZZ7A90Dz3HWKFBvaXfAcPc9pP
GeATI0kbXzyF/u5Xgi2bHRbo4xZGAbv2Vuvl1maPLIy+pRylqStdfOFWR1USB+RI
n4MGXXtmxIEmw32AMkFKAsDYu7S7gFcipas3pwVzGPb3OYcveszzDb6ce1lI40kE
DDDS4dBI2A3deP/Qp0VgSTjdglSGHB1gJIXYqRjDhk+i+ehUobmvc/fV3XiW89fp
fztyCSKq+CKYduseT/HVuOvGwtwNCOj/BIF7BRK4FhJ7zGt6tq7cT4Bim1lLELfz
qI4NAQM103pu+UsvaUKuwwmSwdE2OOK9mPsckhi+ZT3yWGJDgsjOjBoPwnwFjyUu
jgm7O5iwVhexL7P1dUYQtvRxaLR2xdunEvAAHT20UufalChjNzep6S2l6TZXFRLk
sGBk9/RKIdgaa2TRx3R5EBP8WyZd4mcoZEXw8J43LrZXK8bt3ZoQdIT/0cOmpOks
lIN9TYPQ1vAhIPRkP7tMHBVA7ounCW2IDNwYki8BQ7+QWErLcLaxieghsCiLdBoE
ahy2OUR07hW3LlNIetekA79P8iZ7tlKaTPP0cXd3TcbsBrgsYsj1v4hqsouh9+jV
gdbU1Ep5q6S/tOw+02NpBXR7b7DT2X0Ho5VoqjZ004/NNrM2j01GOgq8GwXwuYhU
7TJZdsm0PYtE5sRuWC7nqE87RJYNmXPHE8KXvNoMPd7IVu39khN2bpRv8ZcN84ko
itYXZd8rMJGOUEJDGfVdhvjBPMWmsGGnsOSbOLvfaIV1yygtTBCl818Bg/RN7kM9
CR2VPXy4t2Yo+f0WHMDlRCRnMVgvLcQbOstRybdpgsbWFH1sB4rd+nLvRm67/o2x
s/a6dGapEeWdJYwNYOqOR2WiyDPUInV+HXVBX93GBBryqs+VY6zv7XoXfcNKgeua
+bLxQgWqTBDtSwSycfAwawq+Vrxm3dntebPjTtLFSi2/AT0W6mTBvyyG7wph9icT
2MQnoIDMEvBlwTMhw14Xu95SCBRlZ/Nj5YG6Mqje6AxOzTbZOFUkaiU0hUP/DCkR
bb5YfR06mdn3RVyEc2SYdYyHGzTkoRxSUIkEuUkjgdGvpJYslDwTZKQJwqmQ/izx
e8vfxJAMrU9n14ZzpljrimLe6K+c2bAK+2q0JTyKdVbNBL4JMogwpX73I4+BHlTU
F0jLkAb5o4M/XEWag1FT8qj0nFB+BqOP5gf4AA+Bwy04htSVYZCgeIHgo885dzqJ
mJGhQNPcH6Zco9DsTnueti3u+D/lpeRCJ6r7lqxstit3d7REkLm6Yn1fcO0QtiZf
GhVyv8XPiHrjSVyIqNHP9TdG5fvJBYSaM7dZrG5WU0P/rJearujgT5n2Z6vzanq6
UjV4p4OsytYEho0QpkuyyXPO7TPQVSUCMaNL9VpShIr/GcFQfgvEYfnhCiPtCSIT
YQuB85qjZR2ppIKQu3bD52ZUdMcspkG8SUe12j688iHQPHMmcHn18SgQ8baST0Ku
+apM0OzO1WMTILxApyyBU5NoDvrwJodYURtFITV2ocTppUYRzD5F3hB7+IyiZqNZ
H/2r/YAzMiae2kTOwEInonwep4M+7RwxLv/WxfSIJzEH0D/vjZdsNkYrK7YQ04YM
mgOPFshwsg6aqkyDt/f6RPBFD+67xXraTPTb15xVmi1212bDwJdYM6rt7Ns3vVBX
BN0OvRYFULDJRhSyfAw06KEOc5k7M1KpAve1dVZxNxqG6/B+acw5VPk6RTlTYfbn
tJbPrYNLvT7+gDBjvrl3C7tvlZkyAr9NCe+ysFbP4UOIsmycdGZFeMsdSEdAisbR
OdjeC5paXvznZA9AqhnqqxfpkX6V4wp/toQEzrposZ6vdX4PnbHGdvIhYNwxfaAz
xSzaRkRdNMv5riA2g3uN1XzgEQ9LdtJErflh0LJ1pX4dZhmlJkCgLwISFExLAkUb
AC8Hi0isdO39xXB2O2R1KhwtXsR0ypNSfePuEa6GowGSz3RcoElVnTVbSc8YkiGr
AfJZVbMKr3V8BXGmiUMil2jj8f2YmquDl75i4vIJ1NU84ZfJgaIqBR5IolrGy1v7
ZPyt1v4GOoOBfHndjSP5/68j0qDOJuimiUVYjoZ/KqbvhdKKubZFCh5pW+C92sTp
IxBoQrVoyLLCdfBBJrKq8GZ42uLvL927D0eC1lm7YWgYfg/n78C5+vwTb3SCwoEO
YGh0koBsRGN/voNCn+FHHqhQNV+2Rys9H8+ApNqwp6nyRwzyhKMlNgavr4qrmUCp
zBSXx26vVw2+bWNPFqhfp3A/U9O2aHkbFWfLAK1qMlRabL+Ad7A0d07uRODI1rLm
xZzrN7KmzyDt+5YEP+dg6+lcKtYShiypjkYcXEnzbrlGMnOezZX+j+KODH3otaaW
k6h/aflfCWnMFbDRdop3Q8JWmsXFoqzgsVIXVDd5JFW77c618OMNhZ0bWFKvF46C
TpJx+68P4PuU2LKawV70qygNv+J2jlz1L7K/6jXWR8uNoKgK1Qv9752X1bH+xSCJ
B4eeg62BOd/IU+sX4YQfAfouq1/nvhmrVgQESIRglOzozI4M9FgTp79H5UixglPk
u8H+XT9WpyjY2mIZGcSzU4FSliy7nbpNKMYoom+lYu+e4YKvoRtCDZ1e+vYPrdi9
myProAZPX2iUKSMXqCGnSZHItVd4RXcY4VjJSt8U9av7cDGk80stdXYrmS5uAStu
3QuYK/SwaN6SqriGxdUgTZZx17itioVuw3ckcuqUbETbbFbf4TrTflcvVj+0FoCX
k4vmVrBCVRa4wp1WXbToiNJW7qS5hSKr0HZSywS0RweyV9JhQnGRsGp8EMbMnG11
6NBqbS35R9GXOVNOzDvzTOwdMbyZ5NGOGUYdNGwDXklI3jUauDMY7sqZwvq/6SOO
dl1RQlhl0cxbebW5eUe0L5Ft0ibMdhbAwa3KmgjV/13cvPvS7ccDvordEkBBDMdF
1eO/snE71xSDfoPYCQYxA5s1q0AIJceN/5L23nPEi7A1X/uNIb9xZANbyyPQ8hpY
865njbyC9kHsK+Ail2ov9PYQayTT3vbrbuegj4YUhOxGGJlRmU8rm6v55PUWhRbl
HtgGhug6HXVmR1HsswD7RN5A1KzfAf3bHU8qApUVkigdptvlEY5WY1Esi1w7p0ZN
3yvqwTQ3l34nmn784FKw5e6ISMxkTYZfjl1YZ5B1MwMrbLpmpDPGpBRYiiODgBT7
Q+8Mf8+oG+hvFHJbLSs6XgUB+y7K3b1b4J8roaXMunwGN4ctXMhFAND/PRBQCUqc
yiTKpvHX5TjOGj/L9VZgeFWW1gW5v6K/ZQb5STZoNqXm3GGgdjh2ssonduaKvnu7
8umjn38IOIV9uZZs7FleT5VYoG6qkgCXc0ibdy8jebvGuR0f0JBK72eEQVPhJbNl
w7JNJtSjVBkD8H5eAM5Iakv7UYHwmwFil4IMCWj8a6ZcZqDItgTRC/6UpzQSrPvZ
WttxIfOPVxQQEl+C68IVNlhH6SMKbGN1cMgPKGpTl8kn+4g8vUP4uCQZt2k+XvKO
qVFSBdlkyD36FJc6yl1EsJ4Wz7/rHHu/xHeZXytNFOHRAHdDyKnNbXTMxlKK9d8f
Al1EtWtKM39CbOp6qUsY3NhLTgCrCSmNgRiLjUs5iL9VJ3YYXEcbj29vuwFuspEv
qhNLAfiK9Cyb4L8XoERawkq6208ufVQVYubiGfX/x6dta1A/GaWpEIi42ZoV1yJ3
6wWRnKYd5gCvt0xWZsGaydWunjUua9jTc+lk7JmY8j6lR20e5YWPXDUsnEPs9k5E
oWlkQ+4ld+ebXDRbeo+0ilRHK2gOQIdtweOTVKoirW8s6+Z00oR1oSHoHpOSw8CD
cAOAWLUMdhtYO6f2XczmWYS/k0885I1LMTmQD8frrTEuzi514fLLyKN9fw/PfSsW
9eTD9fqTVtSQIg2ycCFguH3g5zw4VRHuMvwa8lz+tfaKdxbHMPD6dIzA/3GhCYM3
0tKhUM9EN1t7bowoO1PSHfBeHSbg9EK9S1TJKMg8uPsTq2i9dqJF4o2TDjn52HuT
2J1V12oYVF1TjbZoze9vl7nrjm40uNYWCOj8Jpz9yIn9vtCIOxTOfuk8D0iOfz5u
E3wmolmjDcwc2uehpHt7H+8sQcVF+Cttdpeg/oTny/xvCGy53zCbmas3XVutSKYQ
Zg2g3uhXvTSp4BvSu/Ph4NTnLvTFogD0ZhSL5SvmBmRTZGoEVAxu/PZWED+EqrYl
6m/n3CP3ThIWTPwerz24L0aSNGeLiUBkbMTwY8EngBWchF8uTtM+GXaqMcr0Bd2p
NN+cKpe2I9W4F9X94vJaGjK1k//qNC9gQBiFxkUV+osWWKIwZRUqmH54cUUR9/af
vjY/Ewb+dS2bG/aY5YPT5Wl3b4/sp0ZtedIPWuuL8r1as2NFkab/3R7Vr7/1DYmi
WBQ0QAuWsKrFR+MgR0zMq4kP3ZhNYzrTJBM67DL1/wvzxdJriwysGpLY12I4GhvR
fbPtJRg0xGjWGhuPDS2kfTFkjiYdz/rzfGG91HQZdLb/NQ5jI7W4aT1wqiYkRUrv
ycmjMlJzebyBYsWTUDiTcBbQYjqTTLjbabVj0ZJ44nJF23/4Epdda9SKcy2W6DPa
9w8TUK4+OtykP+oucBuu2B0K1p7oL0bGdAqYU+YBNdNkzrLsv5p9iDM3B9En6Dtp
Bmeg2KHJ99IsN6UqoRvsY+UvjXbfBQUMYozRcMbi57zyTbJDJIP2exRL5OqdpaId
3ttab2UmvESXe6Kebfr+lYdIlNS/rEo4WDTR6jfbiiCMEUxWGXCHw/gKDvlAw9X6
lPlF8lY0iPQrSV6r4hVQG8mYkQTHmoSHLxjUObfWQmBMksiQrl9UIUeF3MKXb2ML
FmWRaZThzTQw8/38MwJkv0OcZ0J1mliCMaNvV49tJgG4x/kJDrceF4+taiMCZ9HA
NYju60YzbS4fMrYRCvU1BxKr0kWIbP6CRs7JXutNrnwlFGXWioNFjc8VWf3eZVCM
aEsEgMCoysR9/FCl2uctwLQfZWiLbeT+FOQlwQEx9lZaV5U0hRlTIP7Oa/SWgUvW
dj5uPtcASG1c3XrRh5j9IOQBy8y9npNqyBDS11w7VT6EWRWT9hZJ7aOLRXT9m/W7
MhCMqTTXvFEaln2YSWLVYj4MaRRh97VjW8XOoajJpSg4udVwZY0ragCwV43Z1z8o
jJFiDgD/ppzNqQsgLYRdFcvwc0uDr5cIdvmQsqw73QArB7+Z7ePQUuOWwCh40L13
F7Xq1XpmGXvAcmfkgV0eoqHV42D2PeiWt/yNRc2ZN2mTZSnauzj4IWkMNilgX8Le
darXvfCurFnRnk4yf6bmFugkjh330EQ11WZyhgvDG+B9MD4MBxNGigthbuhlvrdB
GPAx6K+99Q8vGFztVBA/DoN3H2ahSHbAwXRoydZLzOV0bHM7NTy8f5euoSjPDA3b
M1ayTkkCJuwDz+8o0GgYfaNn7SS+DFGt3iKxIJYOyF2OA7T+FXOPS66fzRqUzWHV
7rpBgV//NYnqTmsKIElntw6aQs7Et9xKaIezOuiBpRP1nVUjkVkjMIT/QRYNP9Gf
+t0KRIv3tKx+keZWA3L0Ex4mo1ZVqFu6pdn8FmV9cVwuONPGqWr2tA+h9bIzeVFj
EtQcbJSjYSbHsogbEck5Ny9N9Z58BvcaggJWsNoXYly/JhN2xt4UUfqFZ3RIO2x5
biOX+QveZ9daazbLsrE9TlI9tD5gZk1/a8l6HGb472F+anZrAtbuZIQsu4NBtabs
3JOHja+NDHKkTA5Sy/JwntVGmhylF0NtI6iYOCqAAGvRKrSh9AJa22suelxAX9+H
D0zrrZgR0WVttJlk4olAKR8u5KC/PipwwMkV1QB+YAsxff5vQWO/obw1B4iaL558
e8ibG6jSUagF4OvBxfbFuEpsv8sUE4gqByM/JdXkVhKMk0iiz3z1okIj2b5jzesr
+Oj8bcHzVGcoYfkFxQld9r5lHuZvLSsfeoDI2zri/vK/hfNsNLuhA7ktQ0N8tZhJ
uh3IjDvQC6vgH9cQPS9cpy7wpvASC2LnLyhIbvuTbnrKT6oZY5tyX3hThO+tqQGM
Y/chOFbvg4m08Sqyl5u2UV2kJwwTnSk8j8pl3v3cuq1fvBlBNUOuZEsRImG+G3Zz
nTyl8cyFcW55jn3zi+8NIzGiUUGvz2ZJOrkBOBOKDZv0z1GBQv4Pmlib5ITyHMbf
e/LB59zSyqSNM3q+2ghKoljK4/Jvy5Gp9ayofmQ1DQezzOOz8qovkHjcy6LXo8G4
Me6vxtQfDamBGt0TrmjL3YQgRdinx6tPT2xmpZom0RsIN405Wh8RqdnYaYS0k53T
ox8TLmrgKTkI/a63I5jQDEov3cV2gVwkZ2i1LxPjnWZaHKEDm8UGhAH+QZdyNbco
PK13weQRkubgtJn51rT49jEn3NSp4xXgHy2yt9SwjOEmo5y4jg4nPpSewVQw16Ey
C5MBsQEABvDLONmDOWYus3wtnd460oAN89aQRUmW71WXD/KHbDrsIv4Vv8PRH66S
ebFyjiE2/3nXDqEHUo5uE78DIDxhOVeuQNBa7x5vgOIHBAZcDP85a3B0Qojl/A9v
DKy6N36lwvMpDk7YkDdqfjpl6VLSxdNwcmtMmHULxDcQd7/VWquctvTVR8HnLJQn
rRhd0Ak1ZhMYxHrNHSm6cggBrROVZjNgJDzlw7m4JkznG+2NP/f7oHNvcZOfV429
WXZrXbLnca1JTtnjCp4rLDknWC5EspjCG46v7Ev8cLzU/GuiJ//kipzIpZY2zziz
1sMWtj4ObcCTgSAMMgaslLHmuQVA6mYFpvEfI2ikrx4l0NYBcbhxKjS0wV1QUV7I
rqmzqBlB3zFn6tGf/EUO1TaRs88l/V6gmvjJuA63EXt9E/7c4XQqxTgLEVkYAfi/
rvu/vCK7saRX11VWGWfcdWGkwcdAfvEtVskAcCmOJNme430KY4WEesSZ5tzWMRZL
b5V8rHsy9bsol1racVjF95ZTIVoJB6IGtGJ9zWmCsPPuHYo1blDQQc+qs/IK9hoT
p/AG/lsGu0nYE94DgE+caATiVj/Yszu4kCxjazK+iFAtrrRHRpoeIqHaCIv+r5XU
z14jpuTHtWmjzfGBa1sZ/C9Cpj7WWVq4KWBD1uCE3McauRjMW0WhtbCgV9mv4ktb
UP0+y9jmIjZDWenjxHCWRoHgz3SCCB9CEiWL6YlKT0afSFekTypynFhtbI/BA9K+
/qfpkWiY7ppTNY8lYO6uUw7WwqZnJkGs3u3uXFXlXXeUZInXqWRqlR4SeIYQELn1
25W8VeZGtK3rJlYKbpp6bG+VIcRIfni1c/77mQl/gBxtQ6x/1rAyBmJfVKyEnRzN
4wndvceTvBcarijEwsSYaADhmBXC/oRPjxnJGqz0HKDZaelHZp0dsHJzF+uYvMW/
CSaVALX8GbfiAkje+zSP2bjAqsCyCEFuoHesMtg/CrxR9hywK+qCyAI9uPtpf1/e
M0TbAsz+GqZU3PlB3na8W0giyTFqHCnvrw0dGT1wR50G3kUEt2AULJmBWACwPqyb
us2JdL5a88Y9bx62FmY3c4JHOkst5uFFLQcmreba56HBcrkLJSOqsJvPed00gNmy
eRPAI5kHnKD+XwTER0w64qfACI7a7DkFboS7lr48FCLYidlA2f4jh+7eZvBT+1dh
yhOZhuFibaMs/OPvm+TsAU7sjugyxhCrOxgxvdRWyOMhDz7QG819d1qqt+iHt81q
nWiM7ehr9bLOTsOPUM1Bi3Sv3ifH181i0HaPBg2MG5CYqKdBRfrHLmNSVRz6MTu0
SX7X7p73xkJJCS9EBOCV4nAxKS5+LfLDTZbFvRJarmS4HqfisjETNDCg+M4IUlAa
2kJehXYyvhWeEyZheNZ0Tf54CM6wRj/dMvuq9A386E98zwij0go1euB0uCJe3y//
RcRYlQv+tZk7ngdAzyJ6PW2IxY/yg7Qvu0x24oKVPsoI4bs5QOFv7ataVXPQmvUv
wqyEr2qjnjeiA+tC5C7HjTAN1HyBiOXoZKqMOnQr3bXSz9iFsHo+PCguLS1FWU5f
5CyRAV1MH/GOuUPHM3+vxbpeqyC90YSQgIUCmXeGODA8xLhQkVoktEhW3h5rGtj+
ZVFQcpub5GEu4sAiM1ANb2qotM0Jk1ATwWMNGIcokBUu2ZaWlSqmAsfIdZFHcKU1
IYicF7aVC6aGoAdCTwwOBPLLNxm5Qis+LNpMNsowofGSeh1GUUpLViJQYvLyTXSQ
/UInfvWJ2TcVvluqQR0IJbDwDofpPJCABfErFSyO4+M2PD5jMT7+2k1Php2l+bKG
ZFpgyIzAb017mmS/yfVzLXJwD/SXpAAgZWO6qktEyb6VmeoRmn0XZFchgqSaKmnK
+sU30wo2JYCSMnK04SIMsja6aEMu4TQLbIWImcIJUc0jdqLTtDSGPiP+P40PQUqv
y/krnGREhbjCXQMTico/9QOtV0jvctU+AJbo+pAuZZHMXeqSYBijQN2tLScLWhvl
SADpxoqkibWkStLCc7GwXmPVr5/nec5mvemqbqaImS31tXPYQyypmORnLcMjhMvw
F0OPUqyMKVqMTrr55SHs7GvAPQWBB5q8+JIGt1n0udumFFGwknUGCwk73gnZaY08
XTUbgmbdMCAx8zvqGE84NpbwszptUgQyAq66egD39Fzvxe818PH4IE8fAbsjmNi1
hSI7cyLvKzaV9NOcfcK14wbTonB+17ryLxSkoxYPYRkIuSm0mOVJQX9HVH5oFYf2
tVW73dlYb94dXF//WRG1WPWAQ3RBg9HYQ5Z89olSbjlKBCSl5TbOsu2MzjSUWohu
TRudFMdj9TT37+WyjL67lhB7i6Wrcm4f0OHkLEC9LY1VsO0YwC3IeENYuzEBmVlS
y6e+izrcxTQkeV7BpRVQ6M5n71UxchuSTNxm1fNB0Z4nyAhRCR0GRZMLUnyIVlRt
pNwxGNSLGTHeToLPG0gnZJBYTUpG16FPU0pNdPAdnDnUOjEbRSm89GQ+DkgRCLu6
BWFvYcuZfAbQAr64qIIyG6Rl5nbHlP9H6uFlrwzfGnbdnzhY/aC+eNaUQS5pBnzo
KZ+ZXhaSbcZ/xUtzSp12YSfpMJTamO1QEUyEykwDy20jGkcYrK2uzjKhiBXNksTy
Wel5WDm4igfahSEulKuzsCyaqCZ41s2j2dUoFhvTIW+tF+DiMGMRAuPMH1Ao0bMI
mv1g1/LA+ON8e/FUNQr5ACUCQW8/HiD076Ju1ZsskyUi9vsGpuCYpMJRZTJxfJoP
JWqJJZklNtPYeNXpbecvEQ9Ws1RfPFCjlRF2BgOUUFVXdnygz15xQ5PfZyJqs06T
kJxrkMtegwPod5S5xPoZboRLkpSvLgaTXL7OgHEAtDu6xQWz6ubKdaaFUN6SL0ue
FKNLHhNGwDDauK9I20lUlw7F9sz3HuomDuAIXOFJzTgBj87lloDedISIw/qfA1K3
H5FCF8yR61IIAJT4jvuZApA54chyYJVUWYbBGcoLQhD6Hl6WnOVAuPbeODKwyEr0
eekhagguozJiiwp6or84CqSYgUY5EJLK7CiSXjDhqOm0CassMDhAk/R3XVbeHKx5
ApU93znRSYwTFQQE4wHK25bekZHaR5hP6Veqfw1/MBQ5pTohEtX5Ym/0UMhZ8oGM
F7/4Ug7ILk2CFkpVRsayCadCXXU2rZKvDL24kDdXXqKozrBv6Bs1+5bG7eNArO/C
xdN14nZDdx0Q60orxAmVkiFCDRF3TlMubjy8gbgYVrvVj4wfSxdNKJXmLDhIqd1P
Dhras+M0tJt4M39NWfne4+QiY3Bk7WJ7HecFIqaqsh/6wYufwWXqboFbEFF0HVjE
o1vg+Yk/Vl/QkbM829OEqNDpFR1jqpneDm7wePgrWZJ3gJ/duZkD3R+6ON8/x4d2
BMcbYJ+bst7Yy91YRTwvQPIJqNmxTIRnydfwywcG1ub7dIG3LydVf+T6AuVQc/Fd
zMwHJhh1hGcd770ZkfjLBRLuf6Ae1+unTE84ISc6zf1HtYsHSRAYZ+kZKld/FqG1
l87KDuHyLcoUgVs0L0azLw/vmub7SV4H0DTIXHFj7S+ugRgdnoap5AD/x1QBWtQ9
T04abBMBSRm0Ab95MZxUni/7reZI04ON8AlfGXL7ILbatFhKSFIfMUVOJEY1xeuw
1Eb/zzJ1lj6HWu9mZfhv7jHe9yckYCkAyKsJ35EQ8FwFMxgTn8y3Av4cvyHakvtF
3NBioqZizGPzDIClxND7ugmEH6vVeOw1OfOBa2XGBi8mV7yctrvuZXNpwP7iv8Kq
mMzm0PN38UTBm8+2dsfINfEOyI+WwgNhJQ4lrzXbjd2PfHPpbgfkmzOnVEdJODch
aw6YoyJUav2ZIvz69DbQzeeGnwV78/mMcfyf1qVVcgJrTgD1428pt2rrEfpw/QQE
1YeTrk82zuPCKdLjZUguM0XUVHK2FOtlTBc5Tu+nulL0KRN5pJSgkxdlBQRuy4l1
6RkIwAdt2RQqShrvDs8xfxcGYdsBXJgPyJSy9Rhb7HGYVutiUfJf+qmpQJwX/xXv
K6K/t3QYR9FRFNyuPmCQz2aun1OqUCxEPOGvJHhlvBKLYemm0HdAmTd59fZBcz5n
x2f5oAFmPEVr0bzShAMH8poz3tBYNHcYk1iyZ1H8nXGW2F/nv0mjSpEiTANpNe12
edsXQmmihabWjU7mVhhHkvD4VNSzyujOQ98LzfQ/eURIX+lazbEK4ZwNfWbuGYH/
WLr1dcgFNNbysNodK9HGKeVNHSp+W+YmWgbtutEsjL7PX4jw9G4Vp6mN6eKS69yx
HKFMVfDMTlhj1hyBdARhCZcLlhJ+lXlYJ5EENeZxKUancBaWk2tvXrX1ZxD8+iut
P7zz9NmzW7+z7VU3oHDsMQfPwNmB/k9bmyTg9WM7Faf8hFQV+PA0VOrQRL1+bv6v
ELYoHKlqTqqqMnMU+gvl7Aj/0mC1NYcLD+Bm4VKmz7KCOXjfLk34uWj1y0pIEiZN
zOBlTjJI9qCKj89ofVG4iFLUnrCywUzUZfWkbGbN6KsV+tLsdrHoJtq+LLX8tmki
dHH66zH3zip5A1Df0cvxoGewwCJ/+2d8JqkS9owEj4E01r1Fvoacleb3uDU/vGeV
uWsLawDBnyGzYxfX/xj9CFTKG0LuxXLJ++RQyRYA6ydDCoZf2Cf13HyDrUANO024
/9e6kJeSAcS4+brPm6D0q8kpjL3a+91jh0KvI7mm43Y/bT04Us3RvBZcGwqqDhJM
8aOGKy/vQSzism6EMkqpr5xXGFzBIx68VE+uURIXbkx4oT/lqW9LZGBqIWcDQQ8o
mAe7nRFqYSSgHFTNS0f+XOhOQba/F2P7I2hDWjhG4qM6b5d8BwzeXU24n+oNZIdh
t+YdCvx8r9rJ8bG1/2ssCKc6mmw1hqA4ssVftyZXPs1mZGD91z665n7ZqIgKI/Uj
g3FmbA+bFqEqfwG70F5hQb8azr625BWumpU9xS8SpZE8pUZvcFaSBBgtAJ/15rAq
AD0yRg0rGBSv7IKnH+zbB8lWhOJIpSQQpPubC/xGnkhzyeVGs6MgwdITE8fdnqef
JVI503+wDUukV2XECOd/HFx0nVO91NAqFqNGWD7fqOpo4I3ekk8ODBWHKRf77OvZ
9MfWRWEXHhiP3+Bb9IUAY8mVwpEqjrGXJku20d5lfi1xL8lZnw+tzVA+ZxIr6yzw
VB2+C2edRE5qTH5bEV4iP24vjl3YVYeRebkopQodFkaGCeOXYErlp8Hj2N0UMlHZ
MRZVZi/HP4rAA29mSHJEluXTpQ7WRT0Ti8G78BXB5qRhqZo3819Z61wpcNqaTdAG
tD3jFub3C7EYeiUfY3n+tPo5QlvFG1GEr10iSe9GBwAOIKhoAy2A/OSZjqLRCCxS
XhROtC/QKclb1IDIcS/0GGk+cXRFm6WiDuemRXE2GQYpHkdYM4Uxr+Az+qbqVxBz
wRHC0lCgCvpvkfMbOSLzDDTI0ZLGpTzDwDCdem2nQ1dwEUk40p4a/dV8Uk5UFyLU
EQDtObsA7fkrmtiO+M8qRIcmNwSIieTiQ41fGv9l96YSTspx8IKhJfRrxvw4jQ7R
58A32l0GUc/1EBXINi2yAG+dgqurdIkSx7p7FmT073lahh7MDK+pPjV/aypRBTZ9
pSedFWleoPxVLnPvX7LjMBB6UpwdX9EC5hk73320f7rRXeunZm+LDMd9YSDZ/jgT
4UN0yhPpgI9n95vNiSXuR1ZG9/q/x4ZxU0isoYuvrZkLvyS5TFpMsyex/t7rItBU
dC8LgZPg/+s7egKiP1aEtsyBh+jiwWAJ80acHIzpyuO/z/mhVFzmAlswzygT+Drv
ieCZ8gXbivbVlPF7hYjszwDXQrEyDhojRdZAMVqIf3B7yTfA27jaepOqBq5Y/Hqr
1bYKLMTiJN93tcdVJijMsNlim1qOjrP7ibf6tOtuzpn87RZXBxLdiAYKcp49xpU7
O/8ZGixSm/BlNFqbh3iikSFOs8TJvaT9xyFag8NXJFS1L85Xgk0SzOpc2mHsG57v
9OfWCQqyWE6yOt8quMlxU+4N93JvBfhmKeQvgIukkyX4YTiEprP6swvlY1mrIoPE
JIRE5KXDpADGGR9+jYS3db198PT7kxDi45EY7an2QjzjLD1v3AsZB1/9np+hi4DE
oFbUQxvLZZWFZDZ1K919z3ex7x0QP9ChAj5wMme0WtAQA5KHXhWNGT8rIYdtFqdZ
S9quGqsnp4RPyL1HUfjSK4W22zpTd9vI8XbWULJ1/3N78/oSuKGj2O1ynaFOyRez
c9s64JsPO2lSh43AE3xmclVIIw5SQIKcCKO7C2ylGrnExI4py7LEl9xcetjg4pLm
rv+ZTeXCpk+XPgG7uscT2KSSn3pe252BrH/hFap8dE22iF+7UMLqeQkE6fQ4aPnQ
8fb7wy5DtP9a8bvjkzDxd+ZFlzuoMo0XR1P5qMnYTynshj8iEAXkGbehLEgjDtoP
6nEQv2p/YGGVBqbeCdFtwdk+U8t46L8wBB7UMkFf7xxDd0oqTci4HaH5TOS8n2fG
kzNy+38cSNBUFFs7PMqwzzm1nOD4fpu/Wzvm6d5AqZw0BW3Une0C63ia1vUCmqJX
u4hV4V5QX524wbY/aXNeGZUNVQ5jo3PVuvXttLqiiRIdy/UPEGlXj4WsS78u32o8
oDp/Iap9wXdzUx034t0deRMuCLCt+hiF3biR9Jp4dTMFr0YNbuZflXWKgYdmLvCd
EXl0tMxqKzeNrM15h6OUfHAr5374OjKmVVg5KAK2K3WxeSaZJwQH1mAHtSQ4YTpJ
yu/fSANLmSexLTeUmWB3xmImxipVkAgoA/Z4O7qYGnaoqzfMLLkLJokzQR1PyihH
uFQh95sfIE1JFkU7f4n7kqHSscbt70/ovWqooqLY4SV3yWmjp2cGVIxWRJ/ahR+e
FKTbkFNnp64UZVxmM6z5MgoruIkOQdaTc2P+sBHRR8UJbYvqz+mgk77YBSEO1Ean
tRHQgNdWdg08Zliz1/MvAy7SWg/yJNOA1c0dwJxptPSaoLfT0WGk7mz14K4PYQHy
VQ2U8cFCaWO4dcXhkFU+Et0Gf8ODgp1A0vv7/pgufsJoXyd4tyCYH/gbCQkcqfwH
f0RF+MGS4BjcOGYRK2Awo2pyC2Bb8XOGBL0eNiHKMv3kES1mS1K/WBiAw71CgcMV
MeJy1ywPvE+EQMUHVdDpgUwdDPp0+mYTDlSym0OwDiBoLz9yjkQdAHUnxrbz+oFu
+4YAqe90e4V7mLJ3OduZn+Sb4Unuqsokt2opeY7AM+u8zSfbWFHp7WstTQnf/fNm
e8dlf46jR7qn34WyCD42YQopYmaLmPlYuESP98MMXEXrZoph1IiMtK0fME0SV7Z4
CR3PibrcnNvmD0sRblXz9L90nM+lK325xkLxSRASZ9movKne9zHZYeIfoT13qGd4
/iNg9jm+UlCTC1O8QP2aFsjClkLxxmI1dLA4fVDjWjuqgeWDMF11W1gxWhrhBbg2
fvrE5VqB+osL78OeYJECcvEjQxU7+LblUvv2/1nSaYGIvCRRVm/THmTe9gWAVOBS
LUCLWAQHY7aWMdYCcwQAdPakLu1CiD3pWtOnf+gB67gUmwzygzwIx2Bj6yAZghyw
CM6tFjbC4PM/BEHQbRc8DYmQN0Chn+7FkdKgxcJhCgP0WMMYynIfpB7tJ1UbtQ+U
KTHemV29AzlT+Z7IaNLeRKVIe/Velf9ebeseO2xs60aa1b7LsMkoDVBI7CowXK9I
ZLO+wBiC8j2aV6zW7hor+C8IrMlZzOI7KM2uJmCFpmopuZx0it5rQfYu6YPd6ujO
Bty3tQIf+4WTuuh5dBOoipou1CGt0K5NbrSXeUhR3oh93yBXOQI8R2atqeeoNGSE
mBKOGKxwJfrzHLPZbpTJlxBnNyw6w1GNhFzAwTLAckMpfRdNhtouHKBPGtO2TX3J
RI0WBysM+ySRd7awoTJShLwS7LXZZ4aD6KpLfG2T5Sd0HnD0sLnc0Q+dK3cBvkXS
2GrGA2uzYzCAIl77cJyL/S7DxWp9EP4tGo5+nfRZx0aemH5K2HqMQO4LdT99X1wR
eTM4sw81P0IcRiyCymS+Jy0YdCCn7Zn8mlwQMtnAKajn/2Gqi93vvHI0hooXs9Ew
B0ElY8huAvkLvxPi5wcbJwiS5wk6IB0cfKkzzhZh6+oO0Gh/cD+DlzDItWw4X097
5SIvRW+JR5yVz9W4xkO16jpGSYJsSMxYA0vgHzTPjqZLnzLjTmuR/soC/jwmdHyM
kPIEFFSt3r23eyvLTaiBAmj1KXcbsEvFbyVhby9pnlwY5qWCXVrLJu9qh3+xbtfG
8E7poDd9JwmY4RwHtmQfnbaprlFycWW/X2XUubmlnPdOyW/nreJ6msxmPgc3chvw
40hSuS7pqfz1E2MOJHEQ7tjNA+UpJrpynzOwQ5ne7M6NONA+1tz+JCT3J/0vOCLA
OgEYXpECsUcAwJ7UPSyXiUVQzpomNqMsgu3H8NEgZoewDetQdUPZU/ATzyb+TZjR
dIk9ecs38Fmyy96SLbkKaJFe87U9ymOQte+fqAT1ylJX4FLqvapmrTOaf9LPLkJ+
986VrQU6Xo3e717CWCGRr3TqU0y8qmPdM9RhpD6qfLEhk6EP6FklL0VsjICnqjJB
hz8Jhq22wSYE9tB4s6gkeMmAlOyNyJXtPxInuQWudfl4NmcQxBchK1QT9zjBNRer
o8uk0JD0mk4WqCNnHoxAKCR3X42ygH0I8SM1HsZDFGRmtmBYalFJKz5yLLqWw2ck
3iXlbdYdcOqoWo5tEc3OUIFVS4Zixk7EvhBiEn0UfUVhvPL7SEb8rUdaTpp1PYR2
POwVv6NizJ2OOdFnUvlI8L0Hk0CWZIIm93kZGW1OPDvejcHrEfMuXoOgjRrltVLg
1fIpQkKmgo7urBHtyQA0GlRrvw8E21+jLZmHV9EfpJvTc5s4CkO2vl+ILIFUcAbF
vMv9BzW66yqcCBaC+Hhngzd03iJ3BG60cGMeFNvUf11ygYiEZXuN596rcDafquVj
7hSOSNL90O8x2YfHN4AbglkY84ySo7X13rWNxFUtLFJkAujyG2tyHEeoulf6T1I6
PjR+yRRuxbZF9HWTmnWjBXXFRDwtpOYxscvAR8PXIznxHMxo7wdyAXiXSt5/d//o
sSKoSQvFE74hp6cMcD6F3GCI/i8Ahkdbq0szy2GosCgsWlL5Q9YG+8EHk+Zgtdfz
5EanPwsmUfx4SG7GGzUyLRxcvUSNpEo8GX8GwQWR0WZH+H/SbrJI9S9Zib34E52v
JNZlntvZc252GHWmHZXWNnyccfVneSW61mG//T9oQT7b+FVg/2XwUw/cpBD5gnii
lbglS4c7dp8lB78SwdzHcrp2nZJIELDm661ywhELw0C5ZHyL6SnvYA711rQd0YzV
sdY2jeXfN93+9EFfi8eE+hJtvTzBnEHtgsGS7jQemG9Y56iGTfr6AuJHf0HuX4Qz
iWryA2i72vixILJG67pG9osRQqlDmH9/uIUd5h/vrabQ7i8+9NwvjDUbecYeyN3p
oL+hkUtXNfRXFIcmYQQUR+QD36B5B38RcFmk7L6caq5d5EVlUm+8pKNKlRNew92h
XNCsn+lrz27sTFY3PrzcBXvw0N2E5kdBRGqIyBaxmHns+0x3tfMtSvxebDe1cfum
HnpyklpQywP9pZvuVVUoWaaI/QLhsVTlEbM+uK6XRLiMVx4J2paqtMaUDLkS5x3D
e3ZUWl5kPo47A1Neve3MilqFGwtksiDJbOztpLYP2Ed9q1DFEZk4AHzyJyMAhR+H
t1sXkJI756AeyMaJFG/2Cb9XEDupmPtPuFQJ41nO/pOI9yUTZ0Rlyg+gluZ/cyjR
F3NZOdnC5MQKsO+sOw6EwmD/L463aNeT6n+2OVCQICXTNAh5+6gfJWw/LADbJK2a
FsolnxEkpxBItF6+EHwkG/c9SxhYjeyfTQGHZZtwE4x5XCw0IHC7N/qNTdg6RI+n
D8qQmyZMZu+YjQay6XpW6OsQpfHmPA0e+vGhonLUNe78VrBBgEOdTHtmpCLnk+5K
r9q9fRbQ788sj83tQ2cthmm9K+pUhvPfHVISgKcfhbqBkZ3lpjsQpsCgstosYqLo
lePyKiWOPMaoZaZGnP0eZROQFHz3xi7pnTQxJJdhbPlNj2ZlUtwp8DKtNiQAkTBy
s2NA1/HbfHkCv4uW54PSMqJzdc2PAmyftIjRJYwdy7OFddFFuxDW+pDer4hT1oMn
0pjqOClmk4+nC43GzFJMDqZWuOzJtSKCRX13J9/MnTB+5MNF9OWmy0guYmfgx9Ew
MbobtyWO2HHkEIy2zb9vpsz84XcoRJ8rjHVQANuptMUFcR6GZCiYDhxi17Muw1S7
ij3AdaJIS6c7+RLy6BVV458+z42bi05vbYdFlQXpxYxEFU/4yMdLnRgGQ1N4H91w
u75wLvg9uB6DMm+ucwYuqDomKEQfviMROsUicUFalfCT8+jvDHn7SFpUfVi2eRRa
G/yEDRNxOUp4/Aeq6WBDsmsSBd9rHEwJ1XkJkKFMmYF8oMU5XKejp/HWnSTCTMCV
UK6nJ6LvEEdDYNOjbhiBj6duBWR6ePyjBUxan2pgBxKuErCF8TURXWok17UTwlFL
gueWGoSheYVLYPYlpzOfWTr39uWpbFi7sKRKo7Dnw60Bx7lZlAIBUDL8WauJR3xP
ODWL57k2tMW5UmyWg/YMJ31l5llvksNnRCHg8wNdDmXSbJAEz+BYLjNgQijP6Lg9
jUqAxiER9Ciss/NzseToZ7SA0qiNCh/lmMtvZmIsaSc7r9ivP+PiMMMy+gzOYmzs
fX2castLDFvlbHjueSxQVTuPJnptLw/IuvkBzkp1cbEcE0uFFz3dpqcLgqJam1A9
gZTV3YYYSde6go9GBywroGRHwBF7fzTxF1cuWgHf5I7aG9mtmYmBsSkMgwivHVZI
xypp90PWMfZZ/mD2UhjcyWyWgHq28EmcScVzSnHYcLbjI1mjDReuCXc6QucdamPg
3N97cbFHCSnb7fhjyCHO1hHYJiYS2tThIbNaUIVadvVvR6uGCo3C0Y2w2qqXz8/8
NaMryk7sePNtQuXnlSt1SgFALggOmLVZOI/PjB1YFyldtnJfRySTXQK9owfGZPt1
x6sc3yuUAI9OCbJnjj0DGI9g1/2aQ4aaPLrE7VxlNmHPLvL/xfIN3cVzAwEl56rN
2KuUZw9zZBwuW5d/dRgODCigOiiSMXTRwx2VzwS15EIiKudCpWl6K9rivdul96AT
zMZlubJYNdZ2Gx0ET6pE7P/TrBrx+zW1o21jwaKQx0rNwcYo4aGGCUjfTye256G8
qvYN62ns/Cfihl/d6E+xSK9J98/EjhNKDngB+q8Qx3yvagxvr1RC3V2QGyfNOAYb
Q3Vn9gvIqRrMHDis0EDtfxPvg1VeIi/HiFnxkH2v7yJpp+NxIKPfsfnGrAfyhipX
67hMkHX1NGauB95CLdtRMKrdDOfN32qBTLuJK4glPrJp40I2MPBUXSE8+oRd3O6K
FysYg98WF1mXt0UPuZR+qGsqMFn4W8VBIeX3oDsaRAlzX66GvbZABos4CGSD/3S+
y5PmyTB+XGZcUf57qTuUwteAIiX3c3iAmmq+p2Xa7ZASPQTDmmIBYxUaZhTTCCcT
VUeNUoKFLhsmXCOpPJPmJ5CM6IYwUiXO0RNEdXWjUwC+jJkaYgQErVJTdefIF6AM
H4OHkaHO2UOQ1HaiQuyJo4PgqZLDR5sx6/xjQRMUenr/FRpbpdwQTZMptWvMkgGt
N+bJAdY4Bi1MdTiLiKgi6khuQXmZQ0REy9XXmCWPVlC8FMM2UYMESEcAoyHfZznL
BmYmSPDfeE26oyYiUrS2eoQGH1RJQo00Aqha6H83zKWQUjWfjjUpvjxhf4DhK4jF
tbfUG+E6+6flxsf2gRGIvFtuhhb3ZMjDIrqWF1Cw1/DQE07yFId229Wtjwh9FdLx
GZLxxf4IJY7k7yaGWXDwkNevqXpMmBc1xSTNlElVyjg68vsPCxfDE6zISHSxixlB
uv4ql+LfRkag6XHX2Z/NNprRvhxW6srcosuGXo6kZ4KhSdoqglBA5koFZxfokrdR
9JCU2EavYxarZnAOZvcKGFkwWIvH2nH/GoTcKtUNbpEouXGtsJqW2L79yiqpBdDO
RRaXhzG5t0ULaUU5jOuylwJYqVaovgYFOWirLK2KRzT3ORjXhafvZV8j6LerEECQ
9mDeXGFT/sYJgJsQ4lLUs+WlhaPPUXNSTYzJZdeEp0F74Lhe5nYnsC0lhVVo0zFh
cSTT9271PZU7LGzQAkcX3ZmENwcOsyeDGHWgU89aEJ7CiZRWewzaPc5fXdFiKgJZ
TkZEtBSuFxsu5L37BJWXH2s/s9OZ9+BRLC128YotlZyEU0FQg2amoibaBYyRSjR/
Tzk4Gc99NkiNH6wIvLP4FxdHeqS5A+aqEEtGaRiE4LHlVfPzBsO2NBoVwaV0HBd/
dAdGblzyin0XC9tVlHtU2kM0om4vcktbEJiw74Cix2x+6imtt8Rb+8epnjcbnyvq
+6pN8f42+pGazqwHxlM/TiT7DmI2VAq8nAoKiWDCWB9Dd9zFgBNTxdTos63iwYgl
+o2Bf92XvqCJWutKwYwO3wsDvkZ1ET02vpKGQH3GDdXwsvsnF7rx9QEsPiU2VtsD
Qmb+6wLW1tvSYJvY2TCsScqbo2g72jGe77yRB13fuZ+igaG3b0+h6lqKHfC/qtBk
/eTKzgYaz0Sokx3DiOhnjjV0FAtoZ69vi7qlVNP01U+3SNIwxDXPUuCC7Eoo3l/x
clnzGLzeQUpz0/oDzogixgh7/MuTBUrFt/1RU/3H/YN4lrRsJO4haphoXCMuHhjR
KGoYTGY0oWnoylP3oRy12fpgN0qT+++BxTd8Lc0qmkeVaXgQuaIydMbgaRMt08Rn
wTtJP9XOIk1v33INXL7bcF9Ta+KG6cTTdUW+iWcNYGpomq/M11T86ZWN5rSPXOJx
7XMnniCLdqaUBTQ6MBqRxF+iV4HQwS7LqlvAonUMzHS/qydriaKPvvN4AmI8LMAl
me0zF0Fv++JH5E0dMdhX/9B0TAzwukESqms73POkuMB0RakLdXmgvJDSPj319xDn
uxIu+BXxD2gxE1NC7Nb2zfeKe0z97nXpyfkw/ne+mdVuWPYBj0JhfFJFdMg6H2U7
vGyCqPZprtHsjyxpr+eIsOzB3PIHA4/mrkSRA5SvFYcGmmJS+ZOTz/aRasqW4N6V
Iw82QnLpj/mwqLm3YZxYTJYClQsY8VnGCxajPWokU/vv5HHci3pOG5rmtfbMhis8
E9Uoe3ik7Qzhh6H+m0jATIB1faG6z8v0oS3JRvvsps7VM3eMVO9LImrBkvNXcMhJ
kDTQ3Cq2kH8Iog7Xk/kocNfTNh1n1VFlJstQPOF1gWlo2U5EufMbxKN74Hxd45os
xZSHsIJC18oDUS3Zc1ciDPj90LsG681r/4GbBCoO3J+vg4WgnkvFv3TN2kfvMJBk
BslA1oQXYrLDcrv4TdW0uRWXShOvOOMm6Q7AI9mo8iNVBP/Y/7v3LGNrZ9Si/775
TnKo05CNzs4jJn85c/5zb5PoqRu4+mx4vSk6VtNJlNfyFFv0VnAkTyVS1dNSY47h
AeXvqEnSp23C1RSos6SMNZJHQf7/Ii38uIggg6T+0tAH9d0pvQ7MV9Bpc6NrfuVz
4rFpHw1493FVq9mQXc+W4DLd0N+MO+bQXoqHqDIUGPw+gB7MI5kWk8U6ErdCTwZ5
v/8Rt6YyAE14xT7MsqCjwepseb9qovhuHc8DX4U+Jucyw+u1rloESOhjquIJ0nIA
mozYoQdXNiHrNA5tW8teSvLhc8G5vFzm8B7H6SeQ7BH6cGXiWf68BvlpNI3aWqmn
L7O+TF/7kQg6jqZ1LVGvfUvq1ViYBu5HMcHTv3ILRgMW2bCKwmPg++IQoCH+pFc9
Q+JEBetYHAcR25m5zAkGjictFmq74z0qWImnI9CtgIbfZDWSjPbX7zuk6Of8D7MH
PndcCdt/QNVsCiYOhIo3JbVy8Yq+vSMjC67giPQlpkcQ0kMKF2iGLFgmxNYxi+Xf
B3+oKbC0NaA7hD9T2YPc2fC+ywdJxZGNW6T0BCZlMu+HlnCKF5VynTwMi1IAChFo
1nidUgCX7n61suWO3yrZHruMvSEM8RJQLWP0fHAjtxiCrEgeMuOOJ+NBjP9THx2J
aJYwEv+smEzYRS9AlLNulcx2lnNKW3A/WrNJPj9yXouVn2Kq/OvyewnP1yiuvE/0
mZiGKnn1hk0QbAd/eJp8/SeN1x3V8eaOq+3V5hAbwC8rkY0iVF586shuYHXulzIE
XUAFTqMYFjs6QtS9Rz5QW0brRMx0nB9HZfBxWVauGFRYYXDBGrMBAq4PY+1VxxdZ
ZBRwC3IvjXVzSOH9AGoY3RpLLgExFAvCbrdG7sxJcjPWyskOSVZYusQhZXqYohrn
cJMKyYeTKpulJBdk6AbM52TRZPrZKQcCFB219PPz/cKYtzqr1QYP1h0XAI6nrXey
TPEbumllL75KiUn5AiEgYjpcnNPLXSfQCGV1MhSlsMtrClI1khBY1WhQou/5pX7A
d/wKkrXkZTy+EPSWBwkcRcil/LAbFPWeTjOVuaryHMyafKvCLchoQ0+rntqX5ZCY
w7RwxjtlD/qKxNZzF3YOp3T4txnBAUXI9yO4eLfMVIK6LQr3YSm35oIIeK2h68lm
RF+3aWKOvuELmgOKx3h+MSjOFQYYJcD53IJa7AMEfecuWq/+FOqgSmnsBzBe413B
HBVrChw+jH7eihiiY2Kia8/1Eyxgb5/GBCF4mUNVw7Muy41tcLXeT7E5RG28mxsY
MCj6FnBpW95hWDYelVgDbVHG1e/8nqQWY9AwEqTGP+YvH/l6wfUxYJQYuBMC3DT4
SYOn1a/3ozFJAUNWdgKbo88yaKXUSLY/8pbVbkgWVi61ftc6vwJpbMf6cTSaocDJ
06rB/wiqyPY2t/ND11M6D03+4sfMpdkFlDjBKz4A+SUb477xVLYpMay/jlC/4ADI
56i5ope5OTZKEtvyllseHmPrkSsLDYJILiiTZyOEqTGMlAqVXKEwkBJiFKgW4xX+
7VKN7ASosCxWfQ+mz+5WiFmZ4VbyyAgReUIL1/htjC+ttL0ILXPF2eqdwVgtR4QX
LiRM+Ctc/8fI7PhWjtIxqd5NkNo0lUpeQf7tV6489GcIcAddizAMYAR2dA+bnw8o
pNKvIdeVGNIhnCLEXkrjkvAHFhlR6NDAdDFYgYxAdq/P4PFuXNdDriLRLoVerku3
V7SWKsAb/Uq/0zlRDnvTsRE/NoNxSoOmpjJkho0fLrEedmPrND412JUuifh64guS
/hEswUg5Jq0D5n6ImFTcqfOv8f4Q2vkgDdg5bmXW6oCde9TPItwX+Xe79vfbvpzt
Ca00+u+RATYFe8AKW+lZ/OupDecZt5vvDM4En4udG+t+j+KPAKQXGUYcw2tx5Ql6
16InJp7i1SxkjT0JOPAZcRjBUNi/B3CKI9eURhH5LezYwK8v1wRdQpYvqdC36bfs
oV4dwEJIMyvUIy5UCJVDzm+0SU6cTZX3wqTcKziWodYDY/3e5/RZbvJfLWEIFoNJ
JUJbdq6xQcomok9q1+XML5QL7HeqXV5TP/TJ8cpcWgqbqx9XIBZzAWFImN+jpESi
L3U/3P99fRLTKRI8Wxkeg7fTc+wCAzPXH370ZeYVy7tLTcHTzgFJ87k/ed8CEpbN
yiY3gcg/K/6YTTcHSOIuTqWmeuLcWuIq9GKz7cAbeA6jxfOFZzQ7YhqFFkefa8Ni
6kOhbD42FZjBWxXCWEYNsjDUXLAc4qMk/oJqBcvWQmg/zcXRAHoHhNViiOjigFPV
YYamLa4ssnZAEks7Kp+N/LAz55LORsX+b3dSb0FsNb9+NLThijHWkdFMVV2i1E8z
LLFwHPYMbSmBzt3AmFzzvvpUtScgUOgqm4J/+X4oVkm0daHXIw9fa4II1BxEUtqL
DHsUgrhyFJP6V+w0kmjGRRsjjYAK36Oc91rP/NKXJ7PREmKDAQuU7+4XTQI0ls1B
jCKRbUzXc//Fc6ddw+aelM1YYU59jWaSxJP6st8VFK/hMzXeX8zgwVjYSpBIIZmY
oXqJRS7/k15+kir6ypsXEwa4G8SqaXLpgXtq5BbS8edhlMSOPS0slUlCakenNSqn
7e32r7XOmm1262lavECH0o1StWQE4LVTKqsyoLAMcZGdA00GPD40qqpD5nmbSK54
8BzmIfnE/nWuZDHsdLzdecIokvWYwmQlNIiUI3nYBkqvf+3wSJ8lx5b32TxEsA3P
dWCnikk+T2QkJzgYjqJ1fHN6bFOJMtgs20phirsCailC28gV805UbXHxJxa231tg
F+8wNus6jlSMtU3f9AgtBkYcgRSWvpSFsY1aC6tatfU1cKR4U9qwopLbnV/mE3YW
IqoYWwCJ1x1MvXzTrpOGbqN5tUBzktqVoPaLyY3Z9PNuu+YUvbjPNmc7kmYtMFl9
nfSzxCGgWXIvGoTQf7VeDmJiIUWovR5MLG6/PEF7VnU8jz2AtZU2s5KFcUTif70m
knEOoFuEALkFOl6N9Kb8KH3nuj604owzcI9WXqOoAz6J5exrShM/iuvmRXrNmcFP
+l5QPcUCd+y3XgA5zck5txvlPmQNJ90Wisgzqs7FwwUfTbyvdoiehdX4bpfo5OWB
rWFbHfd/BlBPPhkWGxIjoPd6/tAv2QmKtZRLdIu5xnAvsRjbXSfTo6SPTj5w95hl
4/5R1skKY9B9C7w2dcSrda9LMhSVAa8dS5tDmxeXQz7cieJsxX1gSUEnCS7SqYjk
f8jb4kzGVR6uroaU6fM3lkNYD+VP/KEOkoM6AeHiqU/ZPdMMtJrf3WFReidmHM7G
wK3Qk6IztWpt6MiCw0C2geGjqFjwiVL2c4foAJjvfyjRXR12OyveL/AtKaN3+ixL
2uUPbfLrWxfncLVFI+21WzvHcWU6fRyJLGeR5HiXueMQepX0OOW/6XHmPh2AUPcB
wE8RSYNOEsOpzG4DYORUEmtEbzbON/pcwXwdVjQIJBa0KbnH8Y287SeD5UnvIJl4
ggUCo+gJt9G4v4lJ3wep0l2nI2g/Z/DEERZd+OTqNbK+4hIFDcN6JWWY1Am8c9Y2
mMbcEIZA+h/18FIeATy4nl187kZEaSTZCLRKnv9Gmo/QzP9AkBbxc7L38jPOzfKm
qHVYBcRV/+4Iv4Ampv24q5hV/B9IysERZ/Xb4ApE17JoDW1iuV8vlx5ZElbVJaDS
RG4wUt1y+AjYYc+zXIvfriqJ4tMcFvNOJgGW1p6K79nBOiRbIhRm4bNJ9+dIuvh8
fTTIenyNZkMi7z3HUq8tq0cL/443qHzCHiz07F3eUmOaB9sa49lV9UU6i6N0vNg2
enF3zp7tZM2D4Fvo6ZauEr7aV1+l782180IXUQsZaX8d9KKXWMEOryNsKuMznD9N
aTyNUbwQRe0i211EC4nimKe03Eh1wIfBfKKUnAN2IKxKuBZ+H6cRwobWYLfZ2gT5
4p/D7mbuq+6Sr9qT5MZjWogns2CBsWyJESsKR/ziKrjXFM69wO5YKDKxWBlKo0Uy
x2BxRB76HCxVmAuaNbVBtKU24e2IoQxgKHLAaKLQN6Pf/PsgTBgfEiw6uyMCbeMT
4WU94vBfRGi2l84o3YKfGfL2x6OcVZV2Jm/Y5AmRFoUC+hUHj/mWLZlM4epsw9O6
02Ilm1Aq2HmQmUDP+bP6/U5nZkIq2dTeKF3Jt7YBkN9/HMAFa6RdzzZLe1dN1S9w
zzu+oBW76cdQTV7/UQZyncyHuwfCKcdlktH2a/KDAZb6Zl7fvg3KgDfXK23nyBfE
uzgMmrJMjaMJqDStHry6XbGxJmNn1YdyZEOJ0/XN6PbRoVrR245IDHO6qjqM0Zpb
uixisyYY7b9G3CvgYrMxs8wI0rUo/xAB2ZcY0sWPe73DoMPUCiu94tqcVsDAEIZa
VGY2cR38j0NHbbiBjIFKfDkJ2BhdQ1WcDzw+1FmcqfSSgq0SxAHg80RXuat2XlMz
pZyDxVMkfYdsnvfNuE3evcvUFEjrYMKAMOewfjVKH4QzFMlFgiFziIrji58WweCU
Uwd8wY+2NxP8T8VtCkv0Oh1CSku2+khtzpuoHlRv7ck/sZQ2cPyfTjaBfQhURN/j
QoV1pYlKeoBC3Gftvkf1AdN1qM1CQciaA6D1R+P/1HV9etJeGGMEWTGz69ZUZUV/
T9a6BTANutVYvD57i7qS4gnCT5sp79iCrwxp6nAYz8AZVEbG91NKDTNibnLOeNql
TlaAVm+HRFN+0EMqpTRNK/YdgSy1fHLXqMalQOImJC28kaIhD6cJtCJhLH+D7JLg
pz2cjCTk0W5a5QW2b08tZACrbtUPMM0+rRLJuqVPwNkholbmo6VQhgXnFTEVml7V
tcL6brVdw8xToRTxmuH9I/g6MXmgl+ArChwgaPDIz9iQ4b+I2+QqUW1GTSTK5aTP
wOyO4NPK3jW3whHsF4GmEp3yBLSbRm/BTgj4jZTFSP3FgqdOIwDN6pNLGV8oMQKx
s9YnLA0zfKQrmusFdf+bHFSUX5Unig7A9YP1Z8nF8v9yFdcSTljORpKRvSPbipn9
G5NZ9jeXNssBnGhOLLsEbnyaKjq9ouYOS6pMNaP6b/HtXCpB4BKDgv3jjiYNZOQy
s+pNPKvRmnXe6FuTql7Vtj5SEdGVAFTNFruPlN8E8oIvK3dSLUW960vtqUOD4W5+
4hP88CcIUqX3bDKeygpYrzsJmLdwSsJee7GQCvaEW6u3bg6PBEM559y+3piEborV
3W8QpffCICoKDczDmCrOBnXgHWu4PuLDhl14xU47XIJC5SMonT/Xvy8kpk0/S5DF
ZeqB1mQPNYppA8XiuLdVtGrZa+Cr87s4/qvE4+8TaFLheeeoNk2O+upTD83nUTsX
w8GYfZ9ld6OY+WQI/BPiloRhU4SVoDACOZgKceVz8Jy8SBrr+u6Iw3dg4XWPpYJf
l84imPcIgJv6a5IphXQkYLal2BT2rm2iy/Njd41cyFIymXtGqvDPtRWGW1euCcsW
h4PSrWnwawjyg1AG749CxxM4ftNgjXoHsl7+dgvr+i0aQ7kmohZeCI7wHehGupfH
RBIiN0+vBYiKiuGb8TZAz0wTvG1ySX61kbhqEKAaaHCdXh50EooeVLfQg3n4VC/S
POt1us0OnPfXjB7Sl1SGIPvtY+lKGKvVMqgfw98KovZgWrLZd/xj6mkrLvmqebY7
GB390DhlAGisj7rto1e/ys/bqBOMBSd9yrBG5m7G8a0IYWUGtdfSkmZRRoQGOl2v
epUM/D2bVQ5Hjel1CzaIHfij+v//NthoyFWnPdMASHneEa+Pm5CIB2P2rH897iGx
K3bRVZV6xSf0+tQJhdhPaIP+A1MmgGqB+cd6ecGP2G5OICxkjnqXpal5977Z5WBY
98vyB1jbSM4kElXvbyl4yF4BQAJ38pAD/Nd0b1XE4Lu9lVQZDva+1zH4srSK3LiH
Z0q4Jg24xVCWXHm0xaxYsleLyzfRJdd1vU6taOStGzkNhWGJ13guqO3n82uuXnqI
swlORpz6PQfA3ADjSoZj2CyjbQ95CC1/zwgremYR73w4KypJWDKUzLQEJAcJE2jH
jZSPtutMc19ZTwmgPqGdR6n2Sm6s7LE5lXxWvBCrAJi1UeWrsShh5KH+hRIERjxH
mObc1Qf0S5BLEoy/A4cNqHNQ1vM+y3Wt3gOV3qXCCaL7I9JfuewETKJbxgk8tiWe
B+v+ETLzTkGj3bPas+/T/XHj9dnckmuVV1bc2HHdSJbM4Q6QGFZwhxsGOemnzoLR
sMfxQIM1+bEUhfcdljmA9N/Dc+Ic3zSbWE0uOSjpOo5zhmSI1HzRQf4x/lgi4FDs
oeceGXrQBIMsL88xthq8fSrD6GB8a0hobtpXjq7km50lRaeBimRoZozDXjjWIbMq
cZJYNJW4TLjqQi1Li+X+PA8PQ2eADC8pPnUUirS3eH8P+iiWta+o95F9d1kVhIxe
PAhXbwgskPcKNeBIfaklOPUrx8g5jAz7MqKetzxkpR9t2yeAvhIzS1Q8dE1Cp8vn
JQyb3JUbRc5nZNR9z5iZayRpNum+/Wo3hYSEVkjd/n41lDMLPvy//3eG5oMXrNyt
TEW5ha5lAsIU0XGt54UCObqfsc8qaDyVvdAc+q0EESpkjmuctvdaah3pCs0HPnQO
NXp9uCp1xktqvcbbzlf6ihVGiTcitEPQEP0MKCLcFU3JkytZ3BxlA8zelSoZF6VC
J0a1fE5MVPnoKHAx+dIAMB8KMHzNd7EaWol9foZ515sj/1EwgRbUDytgKmB+Pxyx
c2hLHoe6jOxbp1m97R/bnGgVPZ6NE2ZsCimu6MoG1clK/m2xLQoG520dHjQvLccB
4oYSYQqVfUXgdS6sqZkSXw5AbWWdehf0ixmhTN/XA2TT2h04WWyAtWh4nh5FiITj
fsLhJz6Htm5aaXYaQdhIBDPCeiIhJwTdB7eOgVwTsWktcn+Iw6hSeoUypRkMBbrN
lglr2nVpxzX5inWC6GhVapp08EBZIF7Mc/qT8qNXWY8W1nK0Sw6enfHpT+H775vk
btAifVHqC7fp4T4+RVa6TX7wo3po1NViqGOjoTbywAlxmtW7MnZudKfhmJQd70nv
3w8C7c+151yQ5xFbD2/dYsXDf+JTU9bpy+vqXeNj7yPcX32KiapgJyEHkeDK0wm8
BDro4mHcSpeHoAFjzx2CHWmesKp3Vl93HsmgWNux3ze1on49vYiXaIjO5iBfAK22
t4LoCdu2ll2cXpc1Gp7J7bmeblJcNVU6TaWuut8Z451Hng5EnC7/oLI5TjuHZbT6
6E7MXAg5w0du+BGal9t5EQS5tAPwp/YRBI3suEM7PkNXw1Z5AK/886uEj9O54FeV
nkbTDj8GUmeslLLp87fH276xYazQ2PznGzNNa22Gf02tspml6CnCckkkGdFezb9O
yg+m2ISmG/uCrYs4QXPf5lCdBP7TUbj/7zJ+A/ZavgGxTD5Nl1hasaxAk+wlg0X/
YW2FS3o9RHBAXZOL0jlIUzqFOXKtgrU0CCrexKyfMpQ3O+Q+5F0+nXzOPrG+yhcW
aIOH3d9W3+wn77TAlMEu+LYKObOsgM9DQMev6ftj0Q4EE0DpSlRhJPzyaZERpwFN
rUfswQkd+5HmkgInB+3RTgHECOgSF4/mlIP899S59f+vEtQRGlp09Bqh8hO26ZfD
vS6ty5FwbctxL3Q6BoFD9icQMPEyLJn/0XGh9HqhL8zYFTFB9O9UNJVpPsBsCURa
EzUkSYTtuBgm3R3JNvgEgEIyikAfn4loi+JZQ+PzdbkGFxii/ZcUzEQioDkxr/eq
YAMybAGR8SL10qcfLi8xeNWGv/HCo/1LctMpNAwhTUBzXIG8qnwNnERroyg8TybC
/Lx9JVQYbrP1hFALed7v4QcE5wM1ks/GoFjWFGAUDUum7PnwILKlm1uLfiK+839N
qSuV0+YKkdKGUnqYva5VW+bRemAJ38QnoI1sZ+L6o82AJMz+5YWLdWSwH5JrqdMK
sivXLrupXT94ek1hPLn5k3NjHbABTKgYqJ5HJ3k7c2DXd8RERwISSeChbRtMFxvv
kUdgRxzxg0quMGuzFbSnvdHW5LNqMUe/ltSiS7kX8f12IXt4Cie24frYrQMPqJJm
lxzsugDaWIfG5M5xpsrBog7sdZ1tFRkZQwn9CNQ4egsFQWppazICHSBVHUbI0b14
wK3Bjkz6LNicngR3gCXSQztjVGxO9bFqr4nK8D6B49ZZJYFveo2apMmu08Zo/jjX
vzLBx77Qt/Z6jOw3ToEL6PZPofZT/9WB43M9crexOKmU2LEdy/hNUla4yUZV5i9p
Ds3GgnRbc4mfCL3ZbZ02CeJDqxsCMboTRDY3pvE+ynf1Uz2iq/wKn9yeMtZvrTeT
pX8eieo46dJHRSIy7QiLuwQUKv6gdJdquBRQJdu1Y49DS/CrFoM6ZVHRKNUyZMhY
bmFm9UM26sAKluQggf90Ap2pMbc3MimU7X1BS220iNet3jCZVUQrWILGVzbLPSEd
tn+vZdXiRSQIn0bg5AGOsuyCkG8TY2wwXqpxq4p42I+tvtFHJoNTjIutIz6J/HaK
4gNC+1GO5yzx/RE4KX3nWdjSr5D6K5mZ1eILp7mwrnWkrNf/pzhLWGBVQWucYMqL
OuHepffJoF1MYdWW/1DYAYMhCy8FZsTs6XfRHo9ypDPh260KHJAzaMZf1ox2S7M+
72RWRsA6cUOhdRitVae9eYQDJNfHcUo4cE6N6cHhzlpiXoSUZr2640st8jH4U1KJ
TgfpPCr5s+jB3cd0dj/yRdmJ9RGeVXSFhX5B7nm/bvakgP4Q4eyEKKgC6TgolEQA
vnYZdeqUsD+S3kT5Pkf2rYv2zO/ykQNNP79wZSAr7ySldYEnO9jNxNF2SaGl4sE1
FDYk6jQzjw64055SCFqxbO8VwmPcNnJLFNJdHnOhicCXvvYdFuWYcr8EHuPy5cZD
WVo/OyemL4DHcPsnKB/c5Vn3qvf92mHM/4lmTtUHSTGZScFPyUixCppHIK42qT/Q
QjGKC743V+XJoti0DVcazSM6J+LO63+qqenwZHucb9Bhknqwi1G2vDryBdJfrnEM
+nkuyRbW48QTHq9A+0yFWHIgY3HrWNgYt1EpkSgu8DZEv/sLdSoypePLYEC6T3t5
3fIhB4Q4FKf+/ZIgcAZIFomU5Ij4L1dubxIpaRxp/ySA8y6RrAUAVyeVxGHFv416
+8vXoXJtbKnEPbnjl81GSozfiJi9rd1iPm0VWlM5pabKTIPgZNjPz1SyMqAl3+i0
a5+KG5FT0EXWlXcoIajy10OWSR2yScXDT+8B1V4PGcczMb/wSuS+L/MAKYlGnPqV
cQTPbOvh3LcPGl0vWAeGc+Va66fUiUJrgYFsm19FR43m3xzBGZ7LgXBoAdZzgXkP
rUTjHkU/in+gGGPGD1e4gB1rGAW+KNcr9vzAHn/DzRrDFlG66WNa4Z0xQGMgIUOY
cbASr1hvDhgjoDRCVFX1ncPR660L4CrCIJu48B9O6CHnKDo6mSvdW+VQU3SwLQuW
MQ4hgGg7tGhtvEzLyCTSKhu1yXkjc0IeQA7PMy0/eNzUh+GNvKPBrJarx8C7VT1q
Lc/NF/lAepP8Psv0NEXu6a127fn4oe0/vwwA1mChuob4EAqLTHC6oTgJVKTrxbmC
Jz8Y1aULnK59/YWDqQqW+RUCEGoneFCTGmHKGdLXSs6Ew4A97FRt2XG8ahWpZk8s
BZX9pPd0xAFLovvKBJvs7QkkLc4dY5eMtflahUoHRxsUy+WnNSBpN+chsjUtiVe+
jqYgZHiC0DJlcHBRJbPPXGroxNjRwanaOZ4PC5GB761MRXYwfL78JvX8XkGsXxNt
pECHk8xZIu2h8EEeZGgS/+hfsyoLzDZAUT/ZfIrbK8G1OqdfwuyFIMBJqLf0Immm
GNI2oI2iioTCaW648U+aUHKpLZfdpiFjwik6ghnZ8dOdKthaG8BiDwgmPLeSNyu8
HWdBUrxgUexoCh/LIVr+qSjv4QMLlP8uS6EIzN0TLeQ9XRcwB8L0qfRvpmGdRYz1
kuL6Qq6SPxRQKPxVrun9w98Xc4xWZ83bZRjnf+dwctz+rWZT1dpu/gMGQiyUu/cb
my3LsHiXso8keGChRo5y5jF5a/G/U1KC4KCAx0NxGa7rBUdkMCvD5nmbLeuZY1Bs
krTaOuDvQXS8VUO8SxJnPXSwNDaFbnPM0e4YIrC1jMaj7UDG71EOhu/PhQnlQcr8
VIUqERrl+aRdIBZxkNmHXvfWlF8xSPfyGLxUoBBgsEqwPzOC3/eKkWG5nlIhJyeP
8ziIU40bneYq7ljZ4yOvSEqU3sdguePSMiuebney69SvQ1MYdn4aJKx+i1V35s/G
iDJhyGxs+henUcleeWQrqDnWWG8lW5nODhl37zDzsAx9iIHPNGU5Y1RZq3pHNPA6
AilRQ1GAyzRfTVymiv60oJ3hX91AdnUFxpr03NSqkLsukhDrREwcIVAqy2oHviWB
0CrrPZ6MpUn0a3al5r31fV4kISGQeueUc5DG/nLgPp/EzMsUmHl9cNnLknkhxcf8
hsZPoyGm51A7mdXPJDmlIIjgmlJcn46Su8p/rX6aBZwrC+wMKcEUG4B2AQaHsmeh
py3jqMCAIHvGSvt00h9R1S7oeDfQt07g8UCrTJDZWh0epAdi8UV9GuYOmJPgf2pl
0X9YEgOn0GrlhpJgcMLw4Xo3qXNDKR2KbJdE/oJQmH16quilonQeqJbe4EI1huFP
MGZzy+OP82dj5m/WubdrKQU6Kf67EOFqfDQj/LMRVqwt44Xgt6wIEUYqhRNfCLuY
4JOBuMZJefhbgFT/8xHcmVS3jd7XJJ86hrYHzX1eLWLY9Hdfw/4IGeSxFJdwDVqF
oQNn9zv4YmWHMNGMYOQpxs5HuytRzO4Tk6HdUmZXskMbQfFL6r5a0b01p4eVBCFy
QPHADtLfZa7X1c4BHxLMYGD22iSBZW6h57vVEcxtGJ9ybP+qH/OSzbBq+XyAqxsP
2uAJspoyJ9p4pnVJTxDQGUr1NVW+eH8N4/jgjghL2SDVVq/CiR8nNM3BvKohzTuO
u7nxEbct4uQZRVlaIWNw3rIA/ryZKAOM369hO2UYcrkm5p2+P6QMpTUVQw8+a42S
FFtqdnILIvQYVdUg/QHhWrALndP+z2j13KsanvmacvH7gg4ZzK+/roqF3vcCW2iF
jCjdsJsyWpo8aeomboWoShocPOCl0dmD4Ap0SHsx/yTxJaGK7H1A4pSwtbDxqYqb
xWHXMG+1NxKY29Guxsrwkh2q3Ge7CgMsc7iqs3kK+6OFWgsy11zheB4r9Z32OIEp
ab9n6FyXneFMyrRYQ0C84bOc3b18ZnnPAK7bBymP7yLDZwrSz2wl9yImZwSQTjpc
cXsH8yoySnEmZw6nxd+sR1srvoMR9FWsWb8oeZn1h6p2ZlOgsyh01jW7W8KgyUFA
D2SAEN/pYplwSVoM/WEP/CuYKjDPB/EB1Dcfm3OXpaLlQgJUheFAkn19vaRbY/I1
4DIQQSlyDmfNI90NchuwLYT8pZsi+ZuF6RleqydRisEcb3+s+FIoSg19wOghiY4v
a73dR+jcUC5v2uoZUr32Aiv0y7v/IMXIGYUVDMaE66lulDShw4m2v/aFMCeD1Sk3
Dx/k28YujxK9Dfl+hDkCzj0xjlY3uxHRKH/+U4bKQBGMG2Td8bdYan/aiyKgUOKv
u6YA0UH+Uc9EQ44b5UXMIq/z4DhO9Iw+Bv5IOPxIszD0PXBxzGwQxnlRrp10+lqT
aA4GKtop5AlJhcrSaHn3YaWQ861ZgR9hVyXN9A0tFNKijpm/GP30jxw+CiCpDiYe
FXTUOn5jW2ubPF25fSq56WzvHR3x/5UBFsHvVVDDZt/uSblzuluhvLywKK7k5FTu
K94oBwC7VFf2jhj2NPlRixyhRP36rfIhLg3aXovZq+mm7sEaf5JmyzsWw2uvCl+x
Ytne0drkvQbxo1yX7Vb4qnmCdL+sIjrScif1A5/YJIPg8KWD5wPc4GXdBC3YBOVm
PrMvCShf2rnhftZ87itPZRzcV/u+5WMo6ayzVySZpniaJaQ2K20gAwo4wNmkd9Zr
rp2120QA/hVQvbyLOEs5J8C63vkOL/xvjPNF+hOSj6uU7mIZYn0KQGWSsGAvrjc8
pi+O2RLQpfTCju72bolfGdhEevp+FyWk0TpMjwNpB2IdQ11dZzOc/hBENgeAj1fd
SUeTfYnF8tm2YHM78l3NfitW/Pa4H8Ku5C41nm2cydrofC49dAtZ3UOMmemucy/O
ptv4EJaQmwVEFXqvNH5W9f3fmgv4rkpsBDm9ih7dqBDJHePV6/rce5vCKt4Urx4j
YeAAyoNBLO45QS1Ez8HIW6j98QKq7zGVcgkAn83q/oRYoeihCqq3u3+pTVHi4yHJ
M1DNw98kZFOAGLVrC19hBkmIMi8haymxV0CUovOFo1O9Xq4ztFCnZppaEw0Ruzfm
WqN/UBVlIE0DPYO9+RIT3YyUeeNgX2moAelHlwdoYiHUAt5teQVOcUaQgB6K4xUe
rLLX+i77+4utXNUQwJot3LSGU+gBOu3YcHlO3yJ4Oyi8oaCOhqyORyoEW1CWMvgT
WyncNNHrM3qnfG5wvt86CIuA9KP3UBFQv5pVGRc+fFkkqcN36wX/rNfskR0O37mA
yhTzFCMir1QB7/pgt1lLMaqhSqpj+IhYCAyYKJLpCoYcsPfhrYui7TwX2P4eHdrT
ynntO5fJ0ZfN8HLg1RVLWPCWCTBGUl6pwDgmtYdlLX9m+pLpViAUymNYFgue/7G8
mEfIaBIUDUx7D0JDkbZ2TXPUkKvU/bBxMRai5mxjJIR4pQReh5HQNFKUwthlQkBZ
C+yEi1Nyee2KUkLMFB65xT6vINGy7cyPqvCO2Em9byIs/heLeG3YX4HYpKj99ZRR
2QUzK4WxK7evZ7jv+ylTYLh0YiKPrLpP/tnPxKDmbBh1D2GFYpEo+MkDpGEGZW5D
U8Br3MkN3E+EgqaAfmM24fTZuqgwLOiGt7Hox9SlTBi4T/FCs/HsWhFO7FQQO58V
4pqsZaEXwQbyJioB6m42sjp3q/aa3UEA7I20chR4mqsb6vdPiX9Qyk49wjdx93x5
BHANSvvpSC9P42w2AZHq525stYts2+MH23j32EXjR7MXAtqk/I/htBF7CXKWtWFM
6FFPiJmnQfzLGqPWdYox8KQgHrBLbJXVKz8oIhyVO96F539LceWdz40+db9S/0N+
0OqT5C+G9R1hV+XvBqID0Xi76p1mY7EQfYY+mgKkqjTp1M7cP/BEo0+Cosh+6jpD
PpqAeTIDDObEN8Qt2K2W/kLDppRicx46zszFANnp6cSVEvKEfcdhH2Gkne7eO6y1
IYQhi+CRPgumb0o0S/k2EjIZWOT+HZFqk907tMCCGUHKDeNQhcwTog6ejh6zZPFQ
MJB++W5zGgka3+80XOVed7wn7lNKy31zbul5XW5h0l8/xvfxXaybZtQDFMJe2NCF
Na3i8t4Kg0K0P7TwpCESOgK7RAIB7+4f2pWBkBXLEYboaVk/rcHS1fabQO0nWYyX
04RrEEAFxT9vSuwMrTsn1DaSrMIUoVbp5vfD1C5hK9fhsBHxVG3ti7ax5zmyCgV5
rsvDQN5Np+u7NtO4PXeqoN9Iud6wkEUQT2eGWFELXRhpoHAp5tGH3nG7uOgQZlGH
vu9b7yB2zoyd7LwMlG11rg3IkoGyeZJWLLjucg7JbK97ExKjzdaIWShFctQMlBIA
hK7iu3GYftXuj6/TbJ0Ow7gqETDeQhxVIxHts9kMz5mBCVef71CsmAOTaSuR7TuI
P9b+cLfGxH2LQOYlPwEKHsUZ+c+prq/eKDIxt26sFaJY40WI/sVkk3kgEeXH3odm
V/Yk1NFf7WzYf4WhiVjGSTbMB2RSWRkVHRfa/2MKbWah8jsROWQiIDxqVtZCafhg
5ivWJL0QJvpd2OFaaeEciGmgJDKiLrvq36b12LohlrmurRIh/P39TT3eI72OYypx
KgstLfv0xrAKk2NsqLgesDvTjMiw8BuW/b/kGWu/sVNGV/kZdnPQTEpg9Swa/2qz
faoTHEyuOc9m8a8klefYHD0JSx1/iP7+DeWQNwf1DbiokDjb14ZriLqiKqbyEKgj
u1OOWepusGKdIAHqH2AxlefkpcHnVVZTzeEuO20ZyDxln6F9ieFpFVZ0+b2J5AW+
UvJybMVITy7jAgrMh6YvWdcvUHxoDO/ioCRMMj72rzCE0JmWkS1YRINKDbPyn+zm
bLE22hIbr0p2bb2tZyDgBQE0jTUFKhCupVzFK2yTkmeA7iOS0/qAm1kxFdtyUTD1
ekL/9VHgAMGoH2X5Q8kUbMVmMxbgI7ObkBVUjXBbVh1hGsNDa5MQozkzSTa/1ZXe
gIm1qf/r1uD2Eb6ZmMk6Ye9mYwiKf1L923QUIyGk6v1X33hCD82LQ2ec6ESOGzdT
J1lEKbfDyXQomfGgQhwSmEhKVJFcuYLNxuqobRs7wTX0nLCMf77OEEnVEFON5o2t
eFkGwbHnbH9KPEu4hKJg5/TFxDtnZV66ZDEjIND1bOtGOA2GHCuGbCAbze2bzq86
Nu9eVHVwtw7hj7H5XXkJFR7O+tiV5F78a2SbyejMw6Bdh5OUoJin7sPCJJNupqG0
S25Pke0/nFXoZJBnZP8L8q09Iyv/xwtyxfQTyz6DofiCqKEQgKS6/WrDZzJIrwMh
3UmYklEKu/eGsxNzdoXxcoMqGCDXh1xffHbpUA+16UqsORP1CPbpYDX7uN37Fvn9
PoXQoo6ZwbIhZZ9YdkULV6hAMt9tt3yNVTkCsa/cztYXTO5FNQ7qt5DS+d2Y4Hwq
WazM4yk2DGF67mbrLuQFH7W2rTWQ7LsDBwstcl0j9kZgyxwyY+m3sPW/8exYvGOa
Cgi9HmnzzDmZ57AwCSb71rsZY1RFvoxI7BRcPUw2odkb4ufj3TsUZ+wJjf+JGuwX
96zuIKBWMkwy/HeXIIMp5HP3YfyXzdTxgwla7G0eJ5/WIUOd0n7TyEf4GztOyuq6
POdAIu9vIu9zZ38/G/k/ScEMATjiJ18t/GMhHtxZDDUCC0wXzOlD8wmLBDvVU5DU
JwJYSCbNFkBTYgXBu/y71uaE9cdo1ob/YYIhIIOsprTjMu7yf8wjkKNFLSPJy9Pf
HGU491DgxTjOFr0TC1I0dOU06JXcQQfgWClaB2ydII7aEEtclrPaptxoonmB7FUE
788PGH9xecRoZht3oMjA8jSP70S7Z5dMSN76bp/s6wCl8X7UMPIfjT2CvNGC6sQ2
tgn2W10AUOjYQuSVApa/jg8fJi0C6zAGqf07eVZWYZwV0HIbpDSCwMZpMb3uvG4W
KoWBq95ILWQ5V5ap4GL9ONq5NinR+stQvqxxDquFAEqcskxJCB1X+QlLBjyjoyb1
sZLqYYHze+lGp9DKiKA4iFGlWtej7QJxooHTiLF7EdmW3P6ylYHTBQd4fuN9BiJg
rKJ2VOWM4LuxQ424TKCTupwuMmaHyslErFEhEh3wzQt68VKH6oGQ0qVGbekwgShm
OmT7sASlQM43kMkjq5OXtX/GK7EPU/W68RDjqPL/KYAbE3Sh7ALnKOdmGb+7rnwI
NjvSYv4esAhJaXAbw0P5fKF7EDPVcVuVOepicRy7dw4Tw6pDvaI3Kg/xCyoAr7en
ELpFFmL3xDge220eTLJYKlaHztisUe6Zgc/1ppXp6IjUPI+5CGvb1VII8iSboIfO
lfgM9fNSQ+AmOg54CjWDDIcFLuxdcCoqEjkT8IeNuGLxlE/rI6zcoVlyzBoRYC4h
nKxgxEJPKp3BBcxscTSKLbB5utETtU2iOATBIhIBPKUtOUdWTZEn9WwX3mr8K+jX
GJWxL2ir7OTg3z1w7X7AWzUA0Mtept5sDRkIR72h3dRXlRl2DmOWPyJv82yA0xa/
vcLcW6qS/njmTkvIx/wCu8JanaQuRToos9UM+9jCm9p3VzQVqyDeG5fyV2z5bf47
Mc6Fcm0h89+CddZGO3SzniFLpcs6f3+VEPGWuIU5U4xonCMjkRlw+gnK6tZk94NV
D3ZV14dBJ0ZbIl+DfjMxhLG53mzk7qaA7eMJ39dnqNPaPiv/fdlHY2w1raAx1uni
DkXb88sjLpD+cL80SJ0b6uZbQkCapt9XxYQXKVc9jzbwqtiX8RNt+4ffKjrJbOBn
f/FTZX2fe05zjoXxHFWeCC+n6OJWgWJh7SrZDpv+Qf39oGWd9kmaCYabVPTFv0Ua
5T/YaCVU8bZVeZWf6q4CxFL9LkQhQt69cR6pV+p10C8uRpdyAsFmzW8d0+PRa+hr
mg+ad8FR8sxRp4eV7mybJ7NYNfEMlwQa8qDNYPEoe/HtQLXuZpTuFO5xc15wauNK
8PefG+tow8yoegucWPaIjpIsKKI0xRJDlOMgQ45mmuerw5G1ZaWmTdN7E2jgPnQd
JbDaBeoVRnYYz40KOOxzbPwNCCjWH+uRPOrPzc6sJfrf7TgFXC81Xd+dJT7A3WAY
o6wuVeSLkOcVTKGxBTlLOWJZEd99zhQ3aQ7JRNLe8vElS3Hig8n/UitVDuD0252g
Rsj60FBhiJ5OUEAE+fQngLms3tNfQv9o/5o1h0G+j/MVNTG6ZvfNq5RPKzZaDeY/
QeoCeuqS8ofNR/AO3eH/ti2gu1HtO0i4u/oVchNE4CEZ/fJ68g5MxhOcPAkiVXIE
AZre/tF288cvrJZ3JQFKVYDUnNSHdEd1uMXzmVQRlRJAT46fzO24aSV16QWe3tNq
lOfIugQV7Hk1aIaogcm7bv9ow29fjza/Ip4kO8xHC6OO+BwuPWUcESPxvCns8OeC
Nk3A8pZObnwRbeO/6AHtEmJrayj7Ht2ohKemoAWXuQbhNqTcH+5LLzMyw6ZiyfUx
2TXo6MSljgkcSn9qX5IULOSztDsHzsLcqCGa9ZDHkIuDTSy0O2eQocWkR9NHVC/X
cYtCjjkl7cL4n1xW8WSE809XU1XiMrtUGo+PIxP8/o55Fsycpul4jxbpNznNXkEN
WRI3J5AswwHLQORysj0auz1OI0Zc/JWiv9qAGvTSvlhBSydjlAR4ZIqvc66tFdIs
87uJhC3FT0dA3hzPjoSiaPfanaG6nAF6eLD2lpTkR2IF/9IAlamepQVitsexNaXD
el1Yhz3EYWi38AqqeQgajp5sAuSl+EtIIXvPWqP3bQOjqqQaqtdHVZlgKW4SDNfc
7/64j6Ys2D1KW8qpvF3I2frhvt+64WpJ4SIJ41cVs0QM2kZ3Dn76y81I6/KCMFdg
/Y+5QBX9+23gtrkl95Jpi15y/tJuEGRLHXcgPFl8VYplefi90QS7krwoopBRBfRv
Ek7dLel4WyDuNA7yYMyR9+G/r14fFm3APGAeOK+U3RCdZv6i8D5tMNvAKKie+Z9l
zM4XkuvK9Cjl3XlKK+VNmNJrw9+McxENaBQooH1Tvb6C3gUjf/tWJgYrHwB4MD+v
spdKqrOCqO61XEiAXVCTejEMz9jN7Y4jBclyT7HdPlaLrAzGJfecm9OJzYNP3M08
yQwRMzhhjQn/Liri0W07NUanz+LpMsXCQmi6AxQGci7pDGVRA5eMQiHoX7Lv1aNx
rcaTZAW0KgEP+t0zzyswAlycxljAnfp736/FyEInAuARNtvyfkn8kVfiZOZ+pHqH
uWCf1kzaB/7st7lmwovXUhP5mp12M6DP/YKsojnMHPKAsU9bgJ+w47+4GKtcA9wy
viy4MeAqidJCalLqhO/Pph1m7oc8XLbolt/EG+bWYjcQjQjbAx4VihDow8YF1lYN
i0+DbSDwGaZ8yGqfoGp0DGI86Cgt+x1UCC2LbysMHDIzcUf4WMNoyU8p1bsIZ6ti
MAh2Z/nEoShS3tgzTk8opME1GOrgPiVZApO0oxkGIV05VG4gQql5/Jya1hPMaFQb
g1X9Vlq7B8tKVgHz+yb58nXdQI37Mr2k+RRSOjxU+VWnSiQikdfmIrLrDLBHD/I2
gTOLgr52bOFztJuQsCymK48uMH/IIVCpHBpwD/BY0bV69HFmDkv8QXzW3xUTeqKv
wGpumeHuM7AA9C/GuLlke7qxH3DQ45Dr/7/9z/4Wv+Xd3WMYXXY+bkMmeDO8/ZOM
R75eHT+wn94SxNTfmq6VgxF54sEe5ksTBZdxslJhKPtFfbmD8DN/Bj7T3e6ci4NN
EUMEg/HAp05zz/kvjyXm6GtqDDKUKJTduHQ06PHeMisaeQJIRZ1A8f3hf0TgCUw7
PP3NSSR1ztT59bLhSdhKzKnH8zaM20L9w/Zloukapg+tAkSh//IaF1GQ4JbfYw4a
R8GgBCyvJSkH+UG2CIWroIJQ2rW3C3Bw46KH9s9ZSgPPIcXqYFVIWRYoEC0jUT+f
5QOxT5pU1PFB28iFCnefdPfobFpHvUM7tSGgRKEUMuRfDo8cB+EaQk6BbsOBjzX0
Q92aywJqXeRWxsn1za4esrTBu6BuhPzuvRzQRVBzmwYWZ+PQ5KXDCHbabysK5S7m
jZ9EJNMz3eicfZSeyilLMOrDn+VPdok5z42FxgG2KXPJopCqVQUpS+e2pFTUd94Y
wLhTrMqM0TOUP8bUm8DdEuf2Rr3ngQlq6RO/POH6Ome5fvh/RfHDbDqzcaJcjWSz
+nPC9Z3anOWF7DYTqm0ChWsvIaVWvSuWku+elebrB+XWdWjeT+XB7BErakTrT9gn
mwcC8G2VO2o3iG+KZodAJw6XNO+Lo+zACmZGEmLLtWq3JPH86AspPQ/tXJgJo4T2
kWWRH0XvWJzjCkGYVmw2BxKq7I23p7YLxNi61jv89aZ2lKMoU0WiVoYnyFl7Hj+X
eRG+/n7jyhOIaLaWQXhIBUWvBhtqih+z21s3bZmU1H96dL2QJfuh7RtUTrd0STI1
jgg0K5yruYIIfZPZKjW38t0vK3VDMlPLNpRFgXiIIU6/AtsE/VDy0SxDxfXWGypB
/zvvbWkbGHPW4+npotuwEx5HMnU7qqIFuO7gy+dOWBEy8zRuVWolMhckbQfnKUVg
nLcBYpLQHu9Q12PBkd4l2u7gp9jsykFHbt29r30jy/4EjptGZxL/gkPd9QXCLWbb
4fTdMr3gLamDwgDMARnY4qiW9GCM/28emz4yJaOvP5K1/Aqi1ke74nF/nci5hf1G
793us/XwElmUMP3S7i9ZXjG2sMI+k7nDS4UqwLB2pwpVyyGH96kVxgwMHx0R6Rd5
1qSZO7aSoPj938YqbpmeUvVo2us7lXg6032e+tEnaLreKTQnOeXHPuCmC0KZFCUq
9zL5dEKOKwo1pdGo8qQ/hK9Lt9FlCb8MerFLe3se9U8tDzMYEztI/Nqyzqoul3Wx
VpRDhCNoyKnQQ0HfOfp27Qy9tl6mcsRDCpsUTIrGQR2E7dFySJ7n4SzBeeVLWyzH
R0PmnFFcjWmR3NXTxI9LWT4bEsQhJqNtBP1Y8HyRy5PnkEjBOz2QxeSlc5Q6Ws+3
A3dr6X8dPKyLXLocMCHCiLenl1Z7zFV6yh0qG6kQUWRJSnG2IDKy5nrRiKPAhJsu
05NpfNrS3Begf+BLX8ZHgmVqgEXxkOY0Sx2E4/4MqC60uY5H1OiyYz36Yjhgyjnn
7eJCZNR5APB43XhQI+mhe0jeMZPkqdowLvrdeV6QwCh/pq6W+f+cRoSWWDpMOm8p
NOcCkZYvcR1hJ6NavoHhvUOWvNA3lfhjA7mPzq1qyMEPKnZwxR+PL+umaFhrbYv8
XduhZ1x0w1yUbbuOMOiZzmv7tM+S666KMKRcDSRI64Efdr7xBh6JurXTowxVJPxk
eWKeouLFO3k4RfFGuBH2z17jZVcgv3NgP+KkIHPEHVqsKwLQqfe5shy0mgcRGa6D
cGQktfEY2FC73q1KOOg0Aj9I+jEpFvWhmQpLww5VR18qdFfuzmugaOm4tb106+Au
NzzKiknG/72xUEjc+zlPUTm8U5kyRp1IL9WvgdaYiqoy+oCMCci1G5RlwYws+JS9
gpCbA+IUZqkKJgytMCXmIQVfdW23FqnZmmdwgh3y4PMpBffpK/IoTm9H59Sgtord
a9Bzuo8mcsJ8Ke7lULHSgIFeEAhzCgtGMZJNBu5B8NIZoEmuEr9lv/nhoTk4oHQh
f3JxG1UH1RAXq8oe8F77sCYSoc/kN5ZWZO8zteNrOt66nVvdHo/1GuRRVIjnkddp
85ESha+G587PKW0j0MfLzKHt8aB51pmi7SfuXZvOLhSyx7JLfoHHqTT1S30Muukf
d6Cf0ww/G2bu2IAkjVBq0FYV/ZZofvHFIgpwZ6XJg6fRcmPmrOWTztsdIees8KjC
9ooT7QuO2xOjtetJsRclUDlJkfhDWSZGzC7j6j+yUpOsSfdGWJm8/cGtYUzPvLi2
0Jr5LIH96WduAqNQ7FUxB/KUn9rLn061RI8oBNi4GV6g3aulnk3SjR4beSeYIgFr
YCjfV8b5XOqlJFIYjCS4eDtOeK4nrEqrMb6p19zs2HASy9NTZbOq86msLYk2Js+d
05fmUp+Ex+xcMvVfou/m01G6G2+DvhfmAbcUbcDVoLzICqY8BbEZEDO5p1L/k8kV
/oMP4wOIqP+HceZMFXV7A9PR/tp6H2Cd5psgdioYcVIST+Nfcq/LfUmHvPgImfx5
wjzQKJX2gBhpxVZlNTtpTu3ff3dK3dK9NUkJdl3ihsRUTzh+EtPlpl5U02CVBUEQ
1cDGTwvfhbPgL3KLE3H6AMQBh+5G+maN5OyzDlQLMnuf8mbevIWl0rawL7Gf5zAs
usrs7DRBo6RMpP7GviPCFL9bOkqSPxiy5VjFu1Pb2PanKBMkb0bNaHJQhzi79UQ9
E8+nsLrifiwGUWP1RKInAcNwBGdoHNw2EVXjfsH1jxZowg+TOak8v8VVAYRNvXvh
s4nQ4paZ3L/zJeIlabq2bZ4QOx0/mRpnqYy9Bp1thDZge6zms066PXD/bkb+5yzq
g0LuUexy+09+5ENksi5a/TShL9x7x+a4ULsVbCK2CTYRiR7ey3T5K5g37SlIadrL
wKujALdjFaxq442teoJrMtzXfNCWX5+3Fe89e/n8aLcMGIujYqNaQ9DhhMqyYsUw
a45kQSkI6GCo7RLi4K70SkX35ANKnz6H+wBM0qpfzHE94c4EOxT+TKrZa7yjAlkf
cgKCN6Dyfa670EdOLUNmTMLlcvP7r2WJuD1rceHA0PcQ1LKdkP6N2+fLhhUZokm0
0JtWIIKM/KWgJE1peSBB+HFfvx9m1Q9mxJ65CfjTkj3VUpzqF9rmL25r6Iuc0Gub
IXFPd9/dVJJaDQejek14jS2TzUcf+ZYPNi0l0iUrFEAAutAl8Q2alt+ReuOE1RgK
hIzRqnxQNGk+st44YbZtqYR4HB0espNFjb9jJxXBpOQeuK44fkevVETOKGA/XtyB
5BUkV5snt28teR5u0aa8yd9ZoOEKQeuZmjwGvrOL3OXqkTUaYQhfYwhbD+jlU4JD
Dob7H2aLD9wpsP2F0GWhcUKyi5wa5GunR7VqOQSLzaV+7TSbDXudcvlq4KrtxZa9
HchBGVSElAeqKN0TXvTNe4uf7g73FmmGGzKoVj60K3bxcenvDe0Pdc58puelOJ+i
t4oXvQjCprre5hVBRNxf9ynFk4WAy/+Mkdz4TMz9B9/xml8hsC28HRlo8lWyd3YU
2HSkP2fpqWkFBOOEy7bf7zvhwlO5blP9g9Dg5/gE9LAQ7az56asefTsegX9R3TrM
ACsIXG4BKBxJ0qbGNbtxKTF/Prp1hG2l0ykZpoxfv8hM7wrbGxRNpRUWng7sm/QV
WBeIZWLW0yl8NPp2V3erpYzRDBJVCXqffZjO4CDyS4UILx75+MloqJLa7ZTEfyVS
bG0afOqyU2n7JI5Y790s5PBwzWxszoPQAgZmqW3SHz/A/wUFEFeM4D2Gv20+kmU9
JUGaslvh4A0QOAJO7c19tLn2RYF3szRr6f4yFU5R3rN/86YId09jq/VPvSv6qpyO
Jh65zkRBKTu2MpcFVx9i9QSlJXT5R7gdK94ILtFUeca4zCNB/4Q4k84VU8g5IUqJ
cwQOFaaoh9RoR1fkufEs6yD293DLqIkDqKaPsq7II/D/Wdm0v3O/OvC0qJhouRm5
+DoaibHB2RC3vuRCOeFRZIvu6Ti2Vf2KlXyN9ZUvvMbWLpzoEY8hR/u0F4xfoC6L
zTo77nEK/dphnrSUqVd1z871k1L7EAiT2GNe8+vlo0oqK5IKSLm78SHoKY8oqXA8
npMsdDPlg1LQ6Kosvma581rF3TdKS2mtxXVfgkTZa+Ip1YcITTbbS8eY2z4O/C+m
yCrdkAsRKn7cJnrXmCInoDMKNh8qblFXSO6NRM8iE1VP4WIpTxZcBl5B4puCgckc
dyvJ28dv9+zSUcir1WPi7MF5S5f8ZPhzE/mIQ8MJgFvg8ndcJNXMEfinnUzqiSWN
YNAFZSOG04p5hbptt3KcLRkHqN6NQ8qfQOneD5RYpwBzLcXvUNoXEk2o5XznfvVu
0VN3YAALtX4FX1NUBYSbkH2uRVKFEGYIM7IhY0yPF7azpUv4glbJdo3te0+/eZX6
tyGTmUESte2itqwHgTCSpFFhH1n6EWefVqO1Z8AGOxXngLPBSnLgR8YMgPBLZmrd
H5AUpY4hVR26wwI/w25SZkfnboKu+tCAkyWFwZ9DLMql7nc3s2OdT79aWidgrX39
1vXaJ0NrZ/EOL+YLjwvMuvRSFkhZ2ecfK3dwjSqU1yzjuuJI8QAMd3NMIYsjm7KF
FHHBuz684tlDUPqQBad6lXxkKKoJTgSp3bGthsFExqcIkiA9H+gjsSv3nvlI4Q60
R1T7Bex1+pvx901TEJctR2S8qn3/M2oFl8FZbUQa6tjEXy+n3YZ5+HmGDZ85blrY
MAJB2k1/revezzz66+HijCdyfd+d+q2UxOEHZz+iuCwQhgqrCR5e/VGBq4P4LaYO
CN/uk1+HsaJfJvfwb6j57z4LqYyvxjA0iqZJHv33kiK+4u7YaZv3jzNi8sFF8i/u
P3EhGk2+FEUIbSpRBGfRQvukqUclsqsccjnIH4FE/sNDTRaQZzP10xl6xkJSY1BV
jRRsPCGpu2JgoFs/oR4KvScF1AsRKMhHz9Poe+R43V5JaZzICd0Bk/bel69Tomgo
1V281d3koUU7HArF8sZwjD5Fqyk6csS/CSE2J/fYmYAViS0dgdvV1JftfwXEtg8f
rIV6pKTU5pnXK/GMOjNYcAxbvcviIFmCqkGhETaAESMKyZwt7MJFm3/EG7kb/C6U
CaSbN9DqVXNFMiQ5v16N1GEwnxsiIuuFVYjbnvhtED+/YPfxDr1JUJeSniGzNyIq
Yf58Ya0XFTDAMrUYBn67sT78I0GMXtveHJdm36FLnDg4nbWjLMjmktjp2RhricBF
ERPdmDG0HUIxa7S+bNfu7MpU4eEwivenh5bp0ZP5FCW3kAbErsC+5Mx7nLjIRc/n
XwZcSth75aYGLYIHkARTm1+aWgzDmmtO6919U3rUp518XYmH+2jF01P9D46d/0N2
RCHU7314WyltPCbYQRG2cbu1HFZpQ5Xgv4ruJ4tHX9DPpIhYVDCF+Yb4Ifi+vzgv
VS5AMu44ZwPOR1T7h84vJeEjkialkKz/dGFxz5a+d+0DerzrUJ/aiEYi4U9sLYtc
XBk5YwWXH36di7BiIOTfwWCtIRDzFp7IoEFRFn7pJ3rzXn5hjmu5MxqnStUzPlL5
kRzkisXAVxtOQS7Qc1cGFzzt0NxFW47+bsZwpV5XwYRslkef+p7IfXTFSmQVHH41
43EW7zpfTYz6k5txvEaTe3AVDo+OWU/Nbj1N87BgkjpTz86HK05Adz2k+z03pZO+
DXd0Ut0w545x66OXnjQUlYoFPaxFWKDFseaCeapG9Meb6ZXqqSJthQUTR53KGKVD
NHupo+mTfA9cH9FzK8Hr5B+mynAfyipD433TeuM/3HX0zO/9KL0AbFuGf/yhgsT5
kvQL8YniHJe1ceqIY+sim7pJB0O2D2pjnnUb3S2tYC7t21P3X5dQLQYrtQsKFuPN
MUaVae6vTWXBE+rKOPZbpcjCN+T6Q3IYe+LV28/s3Dxqs4Kwrrq6kcRqJ7gBZ1kp
JiY9jwPJg32ULyLJLiki5JNmTA9PTVCuCwfAEJeqkQDI1jIB2QKa3u5CeLUSsDoO
scW/PzlixVqP3t6MwRX+V23PYNLLifp6T1UN2/ZzCHVvzJnhc4W1Sj13EdU6fC8Y
XaM4SqUynuGerXCtrsPqF37wk0jPUhIoBUNxUs3SkB6/DLJ+OF9MCf36BN85hKEJ
QWDBg6VYmbIxoz/j5miSSxLFpwIVqHOmxCHNjpNK5Q33VfU2eUVFZ6WNO5Gq61iV
H+qiHOLnO+PjUyZdA79YFwI0hun88DMEeQ2OaLkwk+MaO2zy1avvnK2gp2C/mm//
lh/q+5Jq4VDBCdChRYdvpVipBRr150g57zUHt1+8XwhbVUkswsU2mA7yOUeLvGTQ
6vgpN5Q4rR/35jS66EQUTVaIfE5sqfIkmtnl5zSOc7sWfdJkb5FVtg6lRQdvWOlc
MtvZtZoeQa/MeDxDoxYSVyogKfbNTRU2Wh7ZOIoA+GLter0MClQH9BIYFWiwLlFn
v1LTfuCkTT2X78jgfwTI2ZM0KO2+0YHLBTJi+IulhPv98IDVth5r35L3aKm6xIWP
gwbZJzviUAI77+ZCYA+APRY9JuRRYec2pI0sggF96MlB9zr4y9/HJN1hNPXj6K6j
3HcIBh57fGf2/4S37aDfw5tPgRShzpVEHrCh+/tYYffQpHzO+UyaehXN4wIWq/Yx
pqkER0LsY57Fz8SLVu4gr8Gky671D91GMG9adFKk9ROTRV6g77FPwbXUrJhOPdi3
YONaWfoI9Sq8OErP5MKTQ3gy4MgzBPNEKUZtN2jQLdRKlTwkVjIMSVwqLiL+z1mr
BqsCzqTmdwDYXGpHMtfBZ/SQ6bqwR6fZQW03Lq+0SM2r9gm/LPI/D7ylgTzlCvBP
54LRDu1jAbXr4jm6sNRs17vjo5eDlBjGoiY9nP3l7LsWzC2kEek9skUvV2EsHp+1
hs0Fd4sifKeVAi8NCtSmFRy0tkpOmWHCRgL+4S9ZD1EdUc+jV1uAqwnCvszwjwW7
jwMvQTrPZcNuAli7mRE33TsiPUHD58UVmdhYeVfKVYHTi8mYxWfZo83bBp4vzVXx
BfIlVjucleY2/NNgrMY5IUuqZEL8rbvSCAnVrXYpciIS2TPBS6sc7xY5y0TCKtem
tqlv64h1VtHIZXHYCixxSv2dSLKmUX9xfY4L15PkpkmU8wAcOFmBwgKSxZB8C/0R
P2tFpWLV8EcDYO4OAo1i1hBFDAL+rvqFhHQ2qf1iJqrc8Q4yfZpB9sg4M2kVZA+H
+6Y9Z9gYq5U4manqhvuaSbwRx5jf/JqW01ZP3fJoSLfBAfsa9s6mGidvmDKw47Dd
KFbsz8Oifse6hKsOYUTgeg8EtgrXy4MHGt3FDmH1hBqzrWWfUE3RpUGG2yG+yNn3
bii8PD69iueNKaqewVc+WO+oRsUhJryiI4uYqi4qXfXge8Nt32TXzLNv9HljdOju
XQfUZ1FicVQFEUKOiC2llivXKwPqeIbuZ3hnTNKSYsKzkbLPGnS3n035fnnQFPl+
gd04jXEVjWzsF+lwkhc93WqKQPehTPgLJIsQGMp3RAcnS+WFZe0ArTJynZkVVK2m
czNQ8Zh29Ubm6N278Gmrv10zew+HPjFhyXifsVQjunDqM7kco1J8+fgfl9XzlNAe
aXCHsmHcwkTSzZkPNKzr2W90pMr9O+qKPhFJwmLRMmoECAsmc19eX3mgVKd0GgjM
gd2VgoTcBHyfEBx+h4gFzyXirrNmfcMbph+h5kOksQsRzSRU2fiCakxy6gHuNJMU
KuW/WQhSSTSCO2NHnlV10KyzlI5IxKqfuqqKDeKDNpEI9pd0lhdeVWFjVJM9IvSU
8E/o86AQjZwJPEfsECiNxFkyrNaPMi4uJKtzqJs0llgLgVPf7y2je0n05eYztRIw
4OrJ+q9uFYcDjVwPNkbeNOZmEA290oBkKV0iAVenMa6p+JbXx0aZw3MfLLcjWohS
QA04IKiq+HdhjJcNpJt33fINqr0dzJWYdCcQH6Qdj+dC4nDu/Hmq6SVxlrr8zcf8
cj7Xq0qLI4+he7YTw8TaicAqAGXEMOVsUqW9cIvSVzpptcLghVDUwExJfrOvGK3t
6QLMiHvI9eLzmAULiiW9fnxhjLFpnLbhmZONVV3lEEOTrXzO8Ydr7Mn/KWyDByGq
GXbmPNrvVEiS0k+Kwf0I9CcEM88rHeEyxpgA6HafK+dEdphWl6Mm2CGGU37DUeo4
jqIJ32/3W4w8FetMdJW29szrJ6Hu8Qg8gtEMuGMGfd2iiQzF6IbHPS071Z2JHczC
j+AtQr9dkk/GN5x6F414nETAbk910pml7DmrDswJBiqnezs6o9c4npHnfQyV1ZBH
OLt7CeGt6mOF95uDZ7dRS9PfuhUl7doNsVOlZdzbKqRXU+4nYIqhjJ0ddDjNGjAU
vLSdHsXPUWWtapKBWFskoexnrEXHFZCIMBBQW0PYd703Zkh3VpjA+fZ/6ZwTUO7s
UJYLWTVz0xvU8kxDdAbBUGVbHH/bg9Rubjdp8sAYsxqwnfhR5xILGqE6XGz5X/kI
3rWgZKpZ5w8ygKXi0q1uUiEOtxviarsaNfXdW2LWOSTo9Bo75yNZ8IaVGXL3njwl
cs0uXStlR2oguoEn5Gh0b5YHDFTPfLOTW6bY/doivgGzY60P9DicQw1Q2FfPAWD5
GrUAmDRFWyID1gqiVuTHz+TnrlSVbjRe3BKjcTiniJVXlbky6sLb7qbKv/8743Iy
3QVkkOPQ8nFqFmZWjArHg7X2OsOZXprp7nSBYCJSZklcL+yj/zMLvz9K0zmU7YLO
543BPhBsHB2laNxXQ2KrxQTa4wsIw4ZRXG0WPF3LqouRAu2oaMcQbLwW3J/Vx1Do
BFgYrNvyh/56PsjywD/DsgEw+Y6MnICcxzCnIDa6gqHl1PCEbkS/3VERndB+yaKD
TiHTTHIvs1oPxbaVuiJzgc/THmdualUO0rxmoFNjwS4g+uNTzEPRc2fkw7tzHZAi
Z4IpqkamGkRWR+Xlx59ojORmjUIqvGEQMYWQ1bRt/r2gLm3AaVtKJWiHBJaI5GoJ
UE7zrDwKASU9qODHkuSvVMEbXErKMRvhmHw5w6IltwZ+t3okjnEQHVgnVNEUHKs+
lO2fhIcfHZFe7PGgz4wMvlP+9l+EXn5iwG+g7h72rh57N9wz3LimVtDZCUSuaq21
vA/XxUJQDdVhsyQvpQMnYKvka4UvyvR+4Yl6JLcBLLB55PlZUCox6DenrrTzIVyF
8CPyvhjeQGRDhhddRFWp5D1nijj6n0z7PbXc5Vn43oGo280A9B2MbOGbqFphjBhM
jkVtYDmQo6iP8f6UKq1p5R0SbFLFYHRpvFl0SbmHegeycpYZbCmSti3G1OISHfsK
lImq98hnUho9o1RYolQZMvuXyiyw1IRLztMtPuXllSXLqgHUxDx80ChUDYzuwAed
sgCvhl2sJwsUuhppDVwjakYlVYCu1Cb47VBk7eTEBSnzpyVYeqAZVjWBUSBTWNOr
Q7xMEBsV/98EbzEnAqbsBqpmb+nMti4dcnION4YKcj86QkzkmY536g3lP+75VLeU
SqzPpZZYzpwITE5ae/dBiYewngiw/+gevTIeviNU8dbWdevxuFXk/1UV6aRsjP6B
yl4A87hP46/dSUiXEL7tR/CbtS9Old0WQyPlaE2m3ktC+XGls5oom0TcL0/Qw2Yt
ajQBX5c+MMnsWleJtpvMazpT5UD6SHWwaOBFRGiPaJz8XAfKyPf8Oy7eNFTIQJtS
NdNIBo1UySbSkE8og3TCdGyt0qCZ97E9F5QOw4GjOlD9EeAtfzsswBesfW2inikN
VsG1/qPAo/QLaYH7pUtyonsec6Z3g5Qo5EqxdozUFHs5k4afYEkc1N06MBszTBPO
+FccsLRTEH13ul7FCjCXGKrbPYp6WwemLt+PSYTf2qQUHJe6hVhfoeBpUzXDKzZN
WnxZnN55RtX7czAjQdK60qXS7AxQ4LxDdJ2wCQSXmeWdDrwO002rBIoVxwdU6jQf
hoOxyYWtrwntucGi7ULxJG/sKXTirU6YjtSfgdKayyYp5Sb85g6xIlQmHw11/W09
MS/UdYrquLl39T88i7u6qe1G06aZnerCmSpITTmtpxjExqG5ZKQ5SzmbeZBDBjhw
dgf41MfRjXtilJCNG+3a1HbOmVgdp+RguIIaYCQJcWD86l3+oa3VNkG0JSHbp15P
Jjnw6OM9c6+H76YViQm9l5ATl7WEN93ovGrvm25ddZuvAQEfc/RNOIg45vEduuBU
0hwcRGwj1Yn9JHPSi0xcpjmDQjinKyOBO8z9en0gBZszRii1cTbdmWGbeP/8EDoO
L8XfuVXvFXxZzLY0KKFqNgULq+WEv4FNFm3/GGoQ0tU1PYlNSHs4x7KQC+zPb6ez
zyI9T4zoI6uGeic34yLkhmdGgHVdvJ84CsZnviPZS4juNSYbQ4oxbuX0Y+ejxlFz
CeiCo6QOmv3iSVQTOaDVG9VRpeUSG2IP2XfUblFB1j13VfvEW4sQtfIoiGBjm3xX
V+Kf1x2DYk4wtFkknTQrwtamw6e4k7MreJU6B4wqf8Cw9/2mq7/d4/6Ud40NArdA
yt9gDKKOhEE6oahCLqnlh6IiWYOQmbOevKEQliVUP3pku3tbgfuRzyt7Ewz3Zrlu
lLAe0YmLwJOYU5Ovgp8NORJxdR54ql+RP0XfFas3DEbnnQf/skERPz+kz564Ulmx
GtNKkWqgnZiXrajAC3qCiJz+CxRHGlm0oZzvBJpGd3fINnWGAkWaS1Bp/CrHAzFj
M3O3YACVWPORI0RVEkjBEuFnYD/cC4KzM91Dq7wPuUcewCxIOVQQxh5rTW57FXsn
IVveqQhEfZf96DDV7QfG2KOAMSXn194xkapDVeLwlMblKbnlLrj154DISFHs6tj+
Q+qMjkVibhg5oG93aKwdrhMMGHbOcFJNfdzem1T8aY6lo+CIO2SbbvsQJf/x3jfN
tYpkptKqekbv0ZeXIVIISf12486h+cgPKAS1dWdycjGQ130TORhS0wa7o+pgJTXg
Vl1bzfdIKkz791r5uEOXE9h3vs5nXV601pMa8DUNqbIizfK7yQ75M9JceiV+hE+F
gz4cUvGSKv5BDepAe69lVr7loJAQSbIrjedK2bTqUDikdqe7tJPdd2ccHTCk/Hdi
S9DUCUlbkO05JtP+mh7cLV8M3ArgvuCITyxftRNC4ein7bQ7BZsrj8pNgOBrX2Xd
CUWyTbMLpu/sENcKhM0oxqlzh/vW9c2QRvMk6WHGrqbAvgXjP/hUS6+FexWcHiNB
+QWrutAXg7AhR142cFGd7QUGcXKdQ/SMHZZvsRkUkhP09b5RbS/AM4RyOQe0LdiT
DnW19UFDNPO3d73Pit+4NNsuAkI/UppIQrSDuj7mC8DtXmGRftF0VnUmFbR2dOoe
kwosfRMjKTQBFFwrYJOQA5fjE5hB1F/37ja08aK7odCupXM+XEWdTo9Ggf9q0Rrg
JNoXwIouoV+aWcSv5LceYWmGl+2ju7iVdLhfLg6p0REJ0L/QTGe8OaVNSMSKm8a6
dRhSowVct5NSseESlTr9IVU4Y/LvsP3QYWM9gFix+Ncy4dnOUSFsq+ysJStF4vXn
HNtFbgXhD2m8sl884kSTcj0yD4Pfpooz5PHWOGD0pQZFnyYmMhGnuAxWvUVjuGbA
rfoFmpJ3ynaThie2GBOmeE6o/ewCJaT7XvbVQuXT3KAK+rDeSWzhpMMGGn/xihkw
TVpNgGFFq1Zqg5WrTHVOZHotMnw3xIIL6WCqY2L5vIQvzNICWRhV5XSriKlUibLd
8gP1qiZr7Ky40Cup0xqH67R3/tB76TwVmTCIFXpxpwGMukzMvHb8OB5pDN92AKjZ
vPmPvWksy44c0tO2d03M5t1hgxggoHMrOspnFUwt8oCF1a226scJuvRrITL7LuqB
99ua6ybjPvWTGrTftEmZDp8BiFkbfTQtGB9bXBwVIy2F2QYojRl4hYjg7haAMChE
QR5LL4lXUfNy7o9Ggigf9G25j9bH9tsGjMLY2yyXpYzpsPliWQmK/TlZeCVshcI1
bdv2b9sLjLsxFOkJvsAr4YY69jS4fF16rffIW9Q1s+Qg762axegT8v1XoI2h23jv
+Xl4OtRmKHyV+Z9eMqGS9mW4oMh868F0a99sn4pOSPEGvM2MAuAd9thCHlCIhmkb
kcUjjDqt90Qs1F1H1LpEMdXt9lY4dYohHoex6k46w0/wT8+lN/MPJU82gljG3i1B
pk3J3RQG/HOuf0HXszSN3csFxsBS5bBoYn8J5i9KTToXZeFNfS7KGNum7SxkTEKH
z51NQIlECBd2vFnX6nc6IDXOcv4JRfbd+Ajv+ZfTWFflh3kXfZCE2O8F+m6dhrPw
3y1hgBZHiOYNRt/3dITCtFmIZxZlUKzMlxcLZYV3/XZMEzCqZxCcDMW30Zx5U2R4
jd+G5WlOXtxKxKKrc+DPofdq3lweAkxR2T3e3o5afWYGjhXPYuuiGj7Py98QaYE+
AsN0ZZOOAezkMndsy3oCculbPqloMSxdv6+2ojTN4ow3TNj0e7Aw9Jdh7qsU+Wzm
IoXeTWjqsH0kdA347okgHj/+0Vzo2jXx98CdOQRenbHB95/9qZhKdTZgT7uAydo3
/XlytsWR3CvpEtiniGQG/V4iU2CSaNxM5Aso8GGCwF/s8Lla7ifxLpkSG50xo4fo
XYPh6rje9gRRLu+Sbs1UJTPf6BXJyLT0EMCc5kKpsiyTXytf31oBjXShAC1UcXD/
UOKlMJDr2+vS37Pyb7X0dvbF+P0q9aaxeG744A4olbfA+RqvPFDNwnSZoTfXXoss
GaExgd0n4b/mEu8HcSybb1FnBgzSTVGgaR9SaJed1NUevNBHrL/wLb6TiEn4DNxv
/TuMBUMwjqxgWl9s9N58W6B+Jot7329PxS8cjM7NS6PMxwp3mUOozd0HJl6me8Cc
qwQTKAyw3ZZW9h0GOrYQ3jIn4M7gwh6p9RlXEsykW40CixMWlols9nI1Yyew5lJ0
OsA6xdSN6y0atIzDVKIJKc6WgeXnJFg6mBAKKRo7xAhy+mqxfmafPGV0FrM9eCnW
3Cpa9wmba8HIPVyLHti4qO3ImVn3qwLuCbvcCYu5sBWlTMPZTmaN2qrSan2oNKUM
nY24QJd5lef756WKmnQEnZyRzT9p7rAD0Tn28am7kVw5s/L8f8Chykvxq3MJKlMT
xO5tv+nsgLGmcHiEsZl8ebBRaREgiHoksw9k4H3IkZPBdi5yKcgOLAwpmvL1Yrgc
lfgXGm386QapcTZw8JaFpaHV48VEV/RQYLULumjVeiudtVSZYdlILtdKnSVf+hck
PSdCiY19bNfGcMLCu80E5Mi4jZook34YdbJBaV5R6WKZGZtgjopcmyzYD4gTjdAQ
AAYK2FUZDMQMYOY7WcHpnLv0jg5iWtoP4+1lrgH84FGAUt56zygNEkRbVLA8Pmt5
YAIc84Gz0s5b1S6vyJvnkWzsVP/bz8xLKUlPMMNxkNLLRqHwwm4W0LJNBkidx0sV
xPiRAuaNuuMuG1Qq2f32umtmr/dBdzoXdF0m5m8wDErzG3gfVhKUFLka93wsm5FT
IR/ZzLtYE4Z4MJGy1MYvQkgU6uqg01HYpBH2SRwvO3BxRs+Tr9Id9PEdmIO/Na9B
zjM7Bec4HTo6lnWINsVNdDuutiCbjQZP4gqWANrlxlG09P+lxEKch41Qxb3w96GZ
Hl3AtztG7rS6XP2Ny4qjQO2P04osNEOl8wJejicelzJODS8+IbCTj4aksyUAOibI
M3Utv7aziZlt5IARen+iUpSOU2YhcFQvbRb59lGCyi1RVIPay84bcwLiMmn2rBc1
Hug9qtUfwzTse2yJlEUhX9NFWV6+R/SwmTE69Uh8qf4fCb8TAXpghmIA7CpZIw7/
TlspJMn3lDThXsbcAQSvbh8s3cfVVk82wYr2yAixkJZXOLH5yhzCCb9qFWPRyIUS
jicetEe9wfWbPB9kgoR4RQ+KNy3kjkmR9L3+MKpdvSEd347QCfEFWavDkEl0TzII
0dWAz+RDRdP6p+2BTpJj/C2yRawqq5BheIUJqUPCOjGbMdLiNRaFsWK807wIDU2o
5zACXeW1f2TTCeqD5y7bPUNS5h/7N9DmMIhhSM/L+g3LcJXiYMQwDiMYAWckV6LS
qhSHv/UqR8r+EmAzFYRaw3fRte2FzRWZxksMOyFK1wOrJyMKtEi9DD0FnaCGUyQA
kCfbbzOHk/WaVOuOICpxLPEkd7/qSwvhiLMnTw1/QD7QTso3w3aEisVe7ycasmlF
Nzwd6k1Nm22K4/jI28GXO/joPGy9ZovKGCnVrX9w2Ih3dLqxaObcmUivXcn42Uf4
koh/Wwnx6sHHh/Jr5DGLCxpdSstAsSbgF4m3sJxtFpqvvJBu6RI4VB4mEWrf1Yyj
BDmhKAKIWb37ulFd0TipVoajvMABz6zLxe0Yk+/2jIv+uSMwpakfy9YQ9eLWh3h3
nAUF3jcj9woMdI9zXXoLjcquS8XYytc/pssk4LlIIclqOP6D63HgCdNL/CHgnuAx
jhUXRdfb1hoDpP1cgaWCBSBoteZ8b9Mm2Tw1zWZvc53UiFMNzKTzjJhtb+buayPO
pHzwSdrKr3BK1FuFtPXOfoa3hFoR/9PK0ksipUz8r04TIEM73Y80UgkWvvRfMJPw
MuHxlZuojFfo4n+Zi0jXxy3ZyxRw9Qoy2NFklmI9PVZDVq4VBziMzS73V2Af55Zx
HDIsitTqMGkLQKw7Qj6NTnGuJ1iYKXE+vb3BCY215buiZai4Ih+lnCOOY2IVxfYv
+tvYrTI0P5cc8dxEbnnOjM7dgaEJn8JzV4zF5U+GFW1x1OBcjQ4FC7RUWps/xPlO
DPv1cQ1DMVO5p1jBzaxrYXg95Kn7BcsOc7BBH+u2gP1c0lhC+lRnE9hwKaIl4Q0J
94OhCS5VmJnvorbDzHkTGqgIg6IVI3zVkJJgw0UdcSN1gVGWZQVEzfSJ+55OMFH4
9YxPw+yi30bgVyAuSPJX+evC4tBO2bfsF1plJugGgVyajOaAHr+VjqnajHxW3X2Q
VZIfzWiPpIGB3lgWnofOXlPSNdrs8N48ArFadR7rF3uEyH4XdpO8I4M4TVhnYh9c
1in5XB3K9oyNLIqo1T0jlViOZIJ7pvzUaey7Vt9doBhyiXW0WdhK4jusaSVYqLZC
R39TLgeI+EICaDu1uZcoEZF98UOWOJg+PfYI4B/HMtx/45EAkjWgvZTOMPODL36c
E40vUDaS5E/XIkavwjlUPsFksoYgRUkFLe48HrwpdibB5WIEYEaDn2cxVOcTSiG9
yTJS1/FRMlCg4Mk4+NrJtK8iLuva91CEcNt6yhqpdRNFFvZC9xRZTHCSIyImoxEt
AgYPD89r6qL+3ExbJI6qwwKRC3odN4Jp2tW5Jd0EG7DZofMyv+/UmDB3AqMNR2fD
n3dwsrBmw84b/BHMt0kWkRxI/m82tmZsQEFXgopoqBDivmGg1hzZXY+1nVi/rjsz
zLdCpefxCYqwphvASOnWaFr5T0bclcDOzOoywzzDv2r1khXWcqFpT8/kMDBUO41w
A/GY1mwKvC+Ym58kdwEnsznlwXD0yKtfV5nOcK8zgQukBtA7NnlJb5hgA7eA6893
S8K0tx/3m+IXYRAgOfLiuBNQgiwjGrxwSKBbX14q72AtitRm1tpaojRMu9hl27s8
l3FYRbTDHeh1krArjKi7e2TaW0iNy9en0q3Kk1tfV4cAGaFeon6Zv3YU5YFG9b4P
Ka3fUBlbmLIZkvv0aibk5I3FnBn6aOhfpk/1rn4qUKIrZfYN2KiOtLbfpInaOkCX
SGERVop2UdrXHXl7kwZKU0g09hxFRsdH+zoSfULn48Ae+9DEykuluBngSD27Qb8p
S9r+O20vGLi2rHUwFbmflXHtrB811pZb4mwtEj55lAU+lec5C0YFleBWIFSS8kSi
x/sJtLehEiodtBiLdYLMA0k4it3UrHXCsnx2HmSs6IlezeQ1Ytj1zbl+nUmSbgjY
BTVPWcYa8FbI94rf6jSh4500yUxpd4YDC5UzP5jncH+sCmtbCsoVOEzjRHADsytc
dbpsT3UkOW0uX3nnLv+yjQNSRxP/cMrseI2CWU7TrVDwRBWjHr6dskkAzrv+W79J
vl8VEBsf458y1OgPLvxFFiKOCZhaE50rTutiBMzKJU/BaN4H0qHtHvLkEfLVA+Ge
1eKIQuP+lG4GyUczseJuPApdxP0N7t6TFtjzQsd8d0VRhloC22qqY0BmoSlgZ9hj
YABlp0j0WxgTQOWXNwsp6SsYoa9R8/lf7eCEIAs+ZYGSLjaGFxeQvioT0g75oiw9
OOXV+h+REIf1NggOHDa5J2C3BeWUbcv+1xgll8GcQk4rJHLpbCgk9Btp+feEZiRj
3IJfQCPkAjvb68qf4IniqIXKNF47lz8KiVEnzGWzSeocSS1B+Qw+I634afhO95lg
b/VGflscduCgCWqRGBGiIqYz3DzBNBp/d7WhdZTDorGbUZeK+pfzqB56VP4WRrL8
Gs8T8UJYhl6g2CHT2kiHdpuAoWt8J3nmxzhI+NFK2doYXG6tUheMbTuq997NWBIH
lpNtZS336W+0tncfBTQErh1om9dRtirfRggrtY+YePPHAh/RRoeIsacx08uhgnI9
R0Xj4h0eRPLZIz7/gxzubKjIlmxKdeh8TaJANoRQYFYxN9yOKyiwEHX/Q2zKFYuf
dKuwJGtdVvB68ck+RRYuVj0H9hWcUFZ2LuGrwDWirZvicwrj5spbob/gX0eFCEXY
KAOF7CcSl3eDEiApJlKax3D8h+aZT9Kw9aCwut/dUHnNCrItAUvZCRwgAvWcCzYd
DTze527QI5111w/uBCN0upvElnIRGnCDz1Ik4Pblt5qk8aEGEMmKzenYLPQHFSr9
mrB+HE4AIQZu6/FOlOgLAGbpOUwBibTJwYFKn7s6R3stIqTLlUnxdF5MVfz+PSBe
mWI9Ow2jEt3tniKKdPzFOFILnYWU7h0qw0Pd1SDbumz+PeC8wxgABlRTqfuEWvUt
/DC05vi/NmLJWM5QAb4T0qeNF/o2NkHNZUEB8jnAkv+p/M2cHPobxEh/sL3vrFrS
WCOers+G/ba3z/tbz+n0ButrzBebAzB5kIeZSSJ6OvRIu8FKGSdssMHV5O9kcM8f
LvKdB5DlzZ+WB+k8fUqnqPZmeOrn0LqqoRjZDovy/21Br7rueOqvoZJ2+sR5Raf/
kgEou6liTJOlY8k4+GgIqwNoGaojx7BCnyfVn5+Jv1sZXL9wFxXRtM2rBAgvSeo3
fn1lk+6olGKX91287foi4MnsAEjVVVNNZ5Jceb/gQcRcvjN9r3bM6//TvCBwB4mu
8OKzlRpLs7KsAXuQZLuh0ftDIw5RXxgeCk+MOOUj57XtbmLvyjSVEBzVBjbgTfsz
KMx9A1F8e8jVxaFfCk+vmDR5IOTLdYP0m5NRCqpE4liL0obARYJmCvWJs0fs5tej
b6vWKZ2OZAGG4gLYHqpx5wey93JgCzkjf4BWn49F9kB9i1VlAw76wIh/Qkpyi7an
TlJJuZJ1FgUN7LGiqyDJifSMP/oFU1mVvpeEedpyZnx1iH7glLyrG1hlTbQsyKU3
kyY5phs2zVHgGc2cjRLV+N2/WPF0T/Rbn64BJ6Q4op8LCVXtBL1jMFHg39ROW2O2
by62kec3mTTJkdsXDk6jnqHQ9hMEh+7MyLU2holkwrsyhLh8x7p5k7HQsHYugpg5
ivjGYrHAdViMlgG9Utis4XoVEdk2sXtSCzb7G/bvg1otnWQ+d/J+GijTXBh9+SQL
y6tu+7RJJFT3QDjABgS0+Gw05hiBv3gjBiZc4aJrlc0rbQoL4l9SE+1pLYEshV24
yryQvK9rQz8sSYnVKSRFPDqJtYylT0DevjBs8yoewD1K56RPflIIfC5HUl0q8bgX
Jgcb72FaPKl2S8cas5MyE76wdmFmv8obYZOkLM78kF6AGh5qw7xvHKUg3RRuH3y4
6SMnEQUoanYFyekRaBIor++1b/imFx0bLT2qiOntXns86DrPaqR7ThizXPazai4T
r9O04hCf0a39QsaxMAPPW3Ck8fwr9+OnGiCTBs/iCWQA8s6VAa8fRE9aLvPBbXqY
/AGdrcV+12jtyh4GxAn3CrqzWzGmjpEFzO+ntxg1ipvhwTW3SMHQqHxZQIe2/k2i
tK87Jnz3aYJdbwl7DLDLOWQYbFNZlHRZ2gzlQbPakyGFsLHlSTn7cLPH5sjeFncb
WA58e2vt1VepYeafnwZOSGTipqpnGdNo7M6woNTBXymHxDeCYRzR+ufDDmeG6F9g
CVnS5rdGnwYWS9pjvQhidkfm9Z6rgByGvwfHvOXWRFq1Nxuh5N0+HqLAjqTOzjUl
dqDjWxnfhpiZ+NW4rUEMXEslTyudCTxOLObrnbpBnLh01NQYKfRGkZhAiIq5Wj3L
J7ceyjxhINCl5KZHZA9lno5pXPz85VK/zCGI0ZfjKCO0fxRbvbE3jEJz8OV9uNyw
DKh5c8YiaFS3yTSI5f8fVQLdAXXXKJ/9q/zMnsEYk4uvASs3aohDvraS3uVrXtRo
spdmkhKjv4V8fjT13p44ebBmSmmfASHp1dzR4lHMkhl77NobEW+Uv3rAnI5qaxnm
oiqHFkAeTKhuyETzGSMvs/rNGwNLD2fYeoN7+FQFt0T3ThjQi/BQmipp/KCab8wP
pp6gXurhB4fvLMqUorng0mG77oo7j4yoHVi4YHjcS3LxPnlAXZ3uZ1lxAGzq8tVR
Nig0y6ZTtaClW1vsBgWvzzFer2PRQQ3vk0tjEUzuYF2BLibx//ED//hU30CYE9Re
X0EjgUfI5PChi6yH1ABVw0IAR1pYFa+cpm7QRgSxbyqs5Eih4Fw7kZJZeqURswAr
ymKYvfRlph8rBHVAbNClPJwgqQHCA8QN0uf/cyVyAFodB78WVgAhSnBJg2enYvOa
HqJj2eZRTt6gmKj8c1pdTob7iB2ZE3zI5HLKRRvS6VJJcHV7BGj6dkEEZ7TCTsDV
EmCSq1qdHLvLhgkzZYabQjnkjPRhM0b/ER6vT1ycr/hdRoWsXS87hVbJ4QgVcMfw
tldlR6fiLcRNydbVB8FkZzEsa98cHM1jCf3YFKO43Xb8ai2l5tOzWnCofNvsV8F0
WPM0zFcIlTKdjX/rwCovmv336K9jVK2q9uIHvAkVrNwmCfNEVDlPA7sbaOLwugZt
qvlUU9qc85mNv2IufO+lFftcm4+xCJEPdkRqB/9UMduq8AqxjQqylR9jGp7EZmVf
BI7HdpYr+3s0i3yTBy1x141BVIXs9DsVOztj9VqAy3dDQYAzwy8PEnWWCsxSe143
ZMg25BljBzA02H4C8kqPeo3qleE1HOUtXc6SdNOeT7JgRzhLdduXYTynr2hBn4m3
E+jj3LESyeQiM+WBesUwnjV4FHjutOnKwqLKddypsbbfL90dCdtcASitSt2dTtqz
26fofXW2Lltr/BCqAaZbWGSujr/rFlofvYguAjtxd/P97CH2kPcpK+/8LuN8T+3Q
9gX61fyTHGNP+IIivsXharDUXtPH9tgfdRcNkdUCxKytlYySWPM0swt7XPRFrsUX
da5Q3OSXsYqo65KsaFHCcJIYK13bCQjuELW0ubhcfUjK5IXm9HOfq1GgIP8OPPM/
7jHYpr85ma4JMjEvxrXa7SLooTsx1WHmAnDLYJ6H2yuIvnLw9OPHX2a++7oWgUNc
OfxUgocYOlhYHFktl5KypK+GRNudjr97GE7B3vR5biHeT0BrsV2TTZKguZvB3WoI
BRn9VmtyIkmxTKmRB+RY8bCuPM0BnL0ua9AVBafAiFih5b7JowmA9TqizohfQHST
olqrIgeg2I/B4PQtyNZlsF6g5dYfpw5YRkowCL6j+Xhk8wZraMyx6uNUJVEUamPv
hSAsK/YF9eV5qxRMg85J7+zyOkflXxgWojlIZEGzON5Az5rNRO5jp8d2uOJRPIHn
rhZ55G/HOOc9nLBJdyTwjUx9MsmPEZCehCvxbqeglITUeesWn/P4qERHgN55on9F
PiIEX+E71sJ5nFtND06ZEa60g4D4jJfpup1/Bk6f9LRqZ8DE7a8wIaO431IY8d6Z
w1wGEnW8V6pwhSgscvhr87oHNEPm0ZUnhK7zABsAcCiC4kVR1q1xMqTIHX5y/nE5
9mfgnU6fDD5GWObBS3mD4OJ11EQK/m6KyyvIUP82WmP5ETXjOSvSpCKN0YDmpXiT
62eLstsdE+fnvvnP5HlZthQJi0Empstfr9wQxxVof4Mrewtq5VSO7ZzHHfRv/YJy
T5EIKEw6vM6+xsRCySpsPjtMLVOdWEY4/07mCEs/e0ajvcFIlE33r4HPsKQ12jGx
K/r8ANKnhai/agNS0krsnwfVKngMNhc8pyIYd4WsY5qS6K1Pg63pNIxGjfhBksAM
nBEsTJiX1cKv6JcFbw48fOIAkVa8mnse6njshZ+JrLeIXXboVOloovDN4hfAvEDn
Xm7zOW6xpXoecCAcHg1UyQIsRgdBLCzJjMVHDVKyXlmdGqb78LfgY5m7YG/DHcGE
7ldg8lUAQZQ51gyUv0tifkbcXrIipOp76+R16v+dzQ/Rkki6VanT5rm8ebmppHBd
9KjAVVNXgSvxsCkUgCUtfXhQgkujpniUgrcvzGSXLV7KkUgRHCI7yYBBxLm4mTfb
3PFdiqvl3RJmyvR3icMl0tGjnPm5aCx6YV3UJj8DoXWrihjrNR+JUqoHCXKbTqch
Gz7l4J3uxTcx/hO04JHoePTYFlgwTjGx+vi0e/OlhyMu/x+xJnxVgd5qA0dBaikX
Qzui23cr4ZKTjhCrXG141CX+58o3sxe2t6jlVNPAkgADWntQO8vPE3ibM2CaoTRD
OdoLSxgAOqn1BBDxBggIpOcZ4LUqF0lQcX+CqerobpijDK6auk/EzDgRLUGbDSqD
F7ibsGwSe+LVLftz+jVCQ3C+u8QutG9N+PHYX7/y//juoGZ7D5njaBt+nMdY47hA
O1wuCPqdRp3+mcYJ8gP15jSVkODEN7ToQZrILHbAilmICTZs+lJg5a+A6HfYCXKY
KyWR0yP+Mw02JT9Wd0TgldwbDXRu3Wq6BrXYAiL42NIndyVYEwFhWz/lLd59TtbQ
yd2ihgLTXwJayCbYh/yGA6uNAzEtW9QbK1TjKfYl0wrylL2qflSJjcjT0PHyJzrh
Ufg9DVqruyb7u+vmjKp+EREXhZwDhMKbfHPqomaNq10WKBJ/q5YvGzfS4nMGFyze
yh29iVSVZi14EcIv1ELxO1GnBE0hwpU0CHEtoO4/n+E7nQdgTSZRxqfSAmyWqqUf
7RiaITR9kBB/Iko40b7Qv1j2aF3593KzBKnLxEYdnXRkzSeF4gsu75Gf43T22deC
WgxCK5OgninkTX1QS17zc4fm6MM9/MjQ642YdbGjAdmXoc/e3wcaNrZIwBi/ejp/
x026OyQaVFECrjU55gHCrJY/AKxVyaKnmcuSyYR7Cim0Or8BTAHa0Vu6QX12QemF
fbbmAGqdhsaahghnVJMWMxg7qxCRSXUbFstISDnFffwiFMYw2N3+XaonFTpzpYRH
9ygot84MtN+beq8TzvCSyolPgj1NLxvQBpWz/pIXEkp+apvDQm48mu7LZG10B5ex
gVN0J4YcapqEBiss+bvzjud1ICOXVQeCNC43BhaLIlm2uNRsnQnD98t5pJHG0fXx
pU7Z+0S7SbC3CLbFM/c/gZTOKi8htkG7JKWfDe10flw5bgBVYYeUyhF5x7kCB2CC
JkPxscf6ryEm6L4j648+O9MWygI/s6SAx7jN5Dd+V5efd4/GNEidYoD5ynBArmCu
Gc4FDu2I/43oMk1Ctca72zjI7k23UPWIBUpERBfG2GfDp6aZhSMrDhplkVUUwT0m
KXCfTIEMb28biU9rNHr9DWnU1C78VU8zw8qCruMfECqr3sB2ek7soFkT8La7RAk7
RoRjUj9oGYU5tWyLAJ9TKDlOhmwYtAgK1pVTvf801e8og2W/azUxGMPd2/UF3ajH
rMk8wKZWTAYQjlSSBCBxcfpuTYGNxWpqLJouSW33DtXj8WIrRqo6EnCtYhKYUsPU
61ECT2ve4NfWz91An8CCDLNGUi/OWMUovgutskxaWF0xF584PNZ0t9LyulB4di8/
hYKhU7NDCweyoNeoc9vUdYNe2VP8K1+l/en42yOK82B4udsudrFD8Ouq9Srtyaww
ERr09uuzIAINy98+K42UBedxB4OzGjULobsyDfwOmege0jnyDTkJTyBXiz4fujhG
9aWxAS/o87nTCWTRyf+bjE+y2GzhMRDQrDqQWKqeygemxpzzjWLEYEsR3cuKGNr9
rira1eZbv7PDp5bSiiW0bC+tvBDIggRPi0d/Q0F0cyL1RNANGG5ZoSB5e6Qcdobp
CHoZ9GfX4l+o6hu1zxsB6uwgzS/Wpq+rDrZP/5SwznZ6wkvaCcvqxEEjXMuEzsmV
ur3ssBl2ImhSTiSoIGkTSSlbVv+gi7XEjGp63Z2zgiukHFW6SMY0+E8ltacBuU3p
0qrc+HmL8XLOACY105fxiZXUDBJm+1JnVMjRNVYyi+o0v7V+voIH/a0YTNlzlR8v
vCsKd7y4sOP5GQ6BGZEoFfGk+/UgYOk7I3UvvvHK2q6A+a3qrj4etRbDTNF7/B7c
BWpA6XdWx9Th1V/ywpjUwPZre8uwgX3uswjbwYFRKXIv+PkQiwCt9kwIyqLRhkTs
WrxZ3tzQGCp8CuWv/cSUBk8bNHpGykNp+Gr/JCioQOv+YyqttpiGOBP2GJTF03H6
OgEiQh0jRoXKzeHo+yai+BsdQdn90spqPCbpVBDYZMzo8Ad4TRQO9w9rdaB5rOS5
tF6ZE/kX1zPggyjemxpsor5s9DUGo+o7jXjpHIc/ZtLA2dLFotkvLJhian/EJSrl
qpZCSN7pIiKCJ3xbpub3sE2g+WEuttP6Rw8LJkEWExtt7xp61VI6AQtfV5Bw8gHc
Ertv10wKMuu/xRU+Z62qUTyQVItudith+6tY94bBjybNuac5c/nwXVukYCJu2Wpv
PLC9sIHUS8nw04LQu17Ols8Q/bR41csq6wSrKihCCNqz1LC/qFXNcgbNLBK6qjwV
ZqbZMcT1tmFT9jxJB8SVvDGVjKlO5kfjitVOreU4NL6g/ORB3bgYwgLPqQ5E73c0
4qdShkKVj7eMdNRXwjutydRSajuxqp8Sj6iKUV7bwnxavXdzYWud51xFvE0cz7Zl
LCOBwgQmGvtCcsVKdIxaIPxigCnJRJKYtaNdwvJYft47VtpYEZlEKvMQB+bLBsST
/vOOSk4/pjHSecxjcgZ1Te1ILvYJoh14V9TYnrBR4IeL7pErkcvLoH7ZvweIWMcG
Lst+KUjU+vy23mVmSx63egSe02l0+eeym6uzTHZjHoJarMYjVEyaX0X4k8SlWNwo
o2ERE11luUFoBlpzeJYI2LOB8E46x0k628n5RZf9q5rJUS0yW9er6oTlfZY/jxx5
hjuwQzcwQkDENx2bsQ2upnrASzq/qrABGWJZmVp7ksCuBST7lSFvIagz1qb+2G71
ZG4bBA8KbBLf3XxjF33ymslFX0cvFLZFxmF7TvbEsiHFC7UKy50QULPiYCZG5bMM
O8x4DLBsUDkaCwMW1k88hIgVdG+mmYjTkCvbjFLxHBFi0AMtbRHL/OWLO0lYW2/v
ksJBQlkY0J+8DwxBrmX97ONFg2LlJFZYJK3OEcDeFZXzZMVqV/jVECgG2rkvPWtl
ncYT+fjzzATdr0wuBSczidLPxfosPD4jSDlgHdgBSE/XwMV5c0dmzrQbrmGONz0Y
+0ObR0ioJ+iAPS0Oht0u2lWuVdH78ZdIPN71eKVp9Fk8ZSVBTam+edCy3uaRVmPs
YAQ7HMyIgvHF6vWOYwhbXAzmHiA+lfvAkLprdvQBFyed2h33gq4PFpM8PHluAuO5
ooNHZRPS10UnXR1tkpLZy0UeMdPNrDdKufeVr8xIHU7ZfMsHP/bRCM+hozMX8oP2
0xgMGPWUVeb6SwVn86/DAARronEito7/FB2yLirTUbpNterdARLuyn51U4YnpyHX
H5VnkAghgaNkzpohKlHb3eXyJXuoDu4BUDmEy/tc23EKdqW997xSRafJ7dwt+CCg
Qb1BJuYd7mKlGyA35lqIbpBIvAryJkQvjRko6tZIMRhhgW6WjiCseakYRZSNYElN
RLqQCyrXV1etuW948l6NofRfB5FzROJJgYwyMeq7hMqdMP2GqEAa+RGRUjYXPvo3
LW4KznFAvYf38aZiQmylJbMaRIE8FNHlwY23B/Jpd2aXUF5XT3/qdDyZvOrhZA/5
gJoLLQLI7TCm/RfQlcXMTLFQd88y9j+hkBVfhcemxB2YvdIkmVHg0FYWWEAbjv0e
tjOgrwgZL9xDvU6QL/EsEG6XXicHqggtuZlVOUmoNn83xED2JsznAshLuKLuMdw3
wWFlGs7hwLiP+7JzAafzR6Hoa78dw1iHpH97pYg6MgUdcmAVtOsgE2OpziXdAP+f
mITBJtbLEGxXlyU58vth/qiycDhhh0hVEWRYreI/FIDq9l9JE9SvVlFJdeLxq/C0
jjMGh+W801WSP2fZzrT5rAwNkVk9PAmwqSF+UjIhK4bwrH93b14k3Muo8jy5POBI
VupF9ZDuIMS293mFIZS9ivjsZlPvt/d5C9XOw8fpWPEIJQMam7wzYR8lyp98iNHU
ZzUasNqYNCGVwEvzEvLd2CrXCqZ8Zl05VZFAxjUAWfHO91SnuBoUE+dWe53vV+IT
5MGscXWhNYc61dzZXXMpqYHT6xtlk8KPVoNbpdhHw4dSYHFPWUoLy5Xt80OK/EOO
m4EL5lK2x99t1LK7Zqymp957bjSY+B1EpZmDsAVt66NhMVYDREj2b5/WdPK/qBDE
BMWcJApklXSgjIif+Ib+tLM9ThAk3Fx1PO3WeWkUArTbngZstwpYP/hs7Sw5isDT
qmydOFhfAjLSlgBd/Kr3Y0tt3P7acR/+rl7Cqki5Qk2pj1ej+PuqDaMnk89RuHRR
SVjxpzUV9FJyuO0HlHnn+OByttt17O4gN/X+gYLI4Sdhe9PFT2kljG/kP7yt9NbY
+EtsxlF/o/JeABh9A5+AqCnp2mr6Un3zD5Fz9MEOB0I2LpYJD2apMY0o5gQ3xRBF
fjfbb7+Gzux6miU/jNug5Lgg2ek3gxk8FaM8EvblYVdwo+vLf+HSMnLzzqACbJii
15kz/GPNYA7+Gtm1RF++ON8U+dLP6IVT/abOsTOTPVvBXEXXaQ4niyupPgVktHbK
5gczqscgZ22HAyMe6rJGv3qDacPw+Fk+EoJ0VJZ7NZK86UhyBanpmpDdCtykUwzx
HkjdR18SvzPPi3DkpG/VHB6RxJRoWUUYhaoJoELTEMs9QjXmUbpYFpwf2m0VMXcD
pyGG7CLu5TG2tWubHNjmtdihYZgyknv6Z1CUWXCjZGv4jz9i4rQpbpfCLR5liPxs
WkbZQZfqE7WyzlrEpnsTJ48pX9Ko8jUjmqeqAfj0WVJeeuDn6zA8zRb2bvylUUMT
qOEUecReWiha8Zrt7a1lpglInfFrbNT4Oor5UDhcrhCpco254ismfr5gZQz9XP/8
CeeCFoBFlV5QgaN3SYGUVUVV2ytcXjMKdBMlb44vXMS8nL9umBEwAHqCdHVvWkcb
cayCrJgCjozYFhlnYj3z41dxsVKi9cS0bFRt7WrAy6h0HX4NqePXb384C8Gv6x3k
0aY/bfLRwuFfbgISfk+kfYmBHJkHl2XHElcclgooeWNECmQouvuZfP4Sc6Wr47j4
2Kr1CD3iC3zq+W9hpryfkAjevHrUuvNI2AcizqjTjNiTiO7Qhrr+QbvT1FWy4Qy2
iuBaspthrN6NwcD252ZYlSEJaJ53rm6S4vq3+t4FvbjOLCjCfsMwjXLKdQgq1OAc
zXzA3Hk6TtD6bHX8c5Xfxuav79K/Y5bqjNC64qrb2CX/N2qqBBqWAEWqD4B7Re90
QITh/iRw+vhyUvDAmeajny4BuhXn7sNwy5KWLCrUsheFuUBaJhrlKVyIT41PCI31
EMk0vj1hKe01ERLG0/5cLvB4I9qZ40HrUtC6X3s5L0ikmF1kTJuAVEa3qGVZ2hnM
1O3WhdzecC7TX3ryaM+r8AAwTTgr1HOX+H20FrZwFpMEW8tB8d5sSJoqmUPs4cIl
+URo9QEZzbGz7anHJH6qwwI70Bh9ja0dK8To6jcGVDEjMALAqREu7IGhVWV24Jif
Sk7/ugSe2QmmntjyXOKnw25RVJBFmXJSkENv1XYyc2EVB4hXxUFyGYCHC3kmncRL
4zPuTATcANVLRiDkoWGYHTAwUkxqYq5OazmZkOAyjAPcr06K40tGgkvHNVlAEDzj
h3M/MkQ4rN/9wQWcJ7TQlvSH0w14iJW1KjD/lbE1xjE1maH7O1gssSTfyS30sE6T
QJibg/S4GTUnPsgF8RptDNYsiJvkll/n2f99HTsdfsLgRnzcUl4lTd98n8CyNLOt
29mK/AKH1GCfVIV+JH+zh/anfcJx8rajPqzeUGmaZrTUaaD3RE91Vdt9MrMWMuyM
cDRiZH/S50bAdIKbancq6/j0LQ2F03Hi+d+MVOKWuY/2JMEhC9piuhU2Yk/vt5lU
lJsUpAkqzObVQNC03/m81EzXfdJg1YpCwqSGO0NsOMdUWqUO4nODzpkhLaCNGIuX
m6DmgOB8j9HLeX175bl+q8jhe4TcqrYJptpLQD8wKZheJkEY1fk7xaC3GP4nckRL
vBWId6aOWBx/6h22Nu/VAXEwVgotD/cVr8B0YHmzeiwCXaYqOVCUBbY/jomGM7/+
mbwaeSFKDHkOO12DoORSn/lZQenNhmfOHtggZXyCtsMlrMlAC8wDdYHCGRAz9/+n
9T57CsGelSPpXjkS+Bq4ZxcVyB6suMSrrXPeVwSnUUCNqGiHYKpQ/0OZvr/uVM83
aj0N2hXyqOKwsXLEYrTIMOi+YTbkTYk9V6rEjmnIOI1cem37VXHRqg4BLWeIeac3
UotsbLhpkw9oKtzen4kztsB2n2bYp5x3/IaiArJ3saG/nAc3ETunLPNBcMGBSf/q
7ezPWTd9EQAO8hzqp7weswDibeCOS4znPqf1cigK7BhpiYot8/JC0sbpWPLo5NVL
jkFGuguYnI1mCM2ZihUfuJpI28YTYeksaZwzxRoQtWzEgznm7CgavDVlkY5xBZhu
YwJsTUCQvSdbMP+2ETCFZ/mjJvSMCOBnzXfATmW2vM6JbCrUGk5C3Pk2yFW3lZUS
ghO2S6yANhdX4OQZdhdnZFB4O71btpfoeTJSRkZxYk2R9zlc6Z+YNZXI/0zArafo
yk4EuprCQRs0HcUqRjkHEyRksBlr/V3hVxqjO54K4VAtLKrDk4hTKrg8lfOpvwG+
v9NplHx4Bcc1k0nIsczVZrZdZn6CyDT+M4gco6ZSQZ6x6eC9kBtwN/fyyMeKUDMS
0YF1x9BU1Dv85KAd02Fa3Nl7eg8NdjPYxVl3ZumYQBoQ+xChY6aGPQxL0ibcUku+
x3ynNUkv+VV8twQw+5iN7RlfzRREzCogZf7E7OfIhng3FlUXmXxv0X/qAF0Nc2U9
9TJdVloFAb9u6aBT1FxvzEL72hJ0p0MKj+ZWOxWgVSIylEDi80la8tqxQQMHOlr4
Ucesk2cV/G5AEufkK7Ocy2WvVxGZwOlJAY2BHqA6LAQcy42eLv8REntct0ZkjKQx
wHiMQrd2yFIzpnV/6ZEV8ma7RcEpiP5/fUArPpAvCn7MTo4bqBxU/7+hA28PmL8v
xjoIQStEMkH31LvyNBv7wSCaZW+Ftl6/C287fBAcpYYNaQ5VekYgbtInJE40tA6f
3pT0yl0vPnWRmeqF574EUeaVd2VWQ+xf9SdwpCK8W4WDLjVtmH1WooxiBcaXuzHT
zdMU5uMMM6JGLsEHGQ9RDzZXwHXoU4yIE7+jORPDflB0Q+w6qagdG5bnqDbN5bsv
HOlMtBO6LZs8HM6ZiPopS2atMEBuykUmqHZXYCEZIdoKWEmdIxNvENHv1H2EXlG3
VmGo7tuFXnZJ2zBW+9V92SNvl2ZNIi3AWAi2ScwKf8XYQsb4zpFH+g70oXcihrfg
apQIN8/y3Rukn5C11/HwI+DkyKlpTQwU0H7KUUObxuKIIi2M1jeYUwlZjL+i3+bv
A3slnczOdf5T5UFqYTC3VApSp0psLbaS+I/uQ+Ws+I9M6giOH0YSujGVWMbLxYEd
hlpTBK6jrCpmQXMMnncjFjLe0aBkAVKxPviKGhYCNFVG0BFlfsrqQuT6VZHExTfQ
nrAZEdGQ5kVW104k2mdIPfUfoJHMbEOwmlmeJoVgjERTAtEClsY62SvP5gQCsjPr
CC0WN0roh5kbtJU4fRw7TKrql2v/uDq2FgslbtfeTUdjlZlskKUdMA5UUz0iOflA
OhaVfW3MFbaYU2VviAGNlMy3rL3yBuvTrbE/HG3jYCILwBSpkM47yMBS5PnmclLR
p169xQ3qySxdrJOe3Rwu2Z+IaBqzayOwVtegk5Qbcm7eyRi1rJZfGbdO1/1VCJeq
m3fOxWpKoMpQ/oLk0rK/vqdfxTWJ6FCpwmGNIHPNh0ks2yVE07rg9i7hjmq6b/XQ
VhakZqMmAWIMWFNT5f7O2NchI+DKqZFQpPaxETFDkc4qa/TP3+LJbfi/jQgCEl1F
T1dbP2JN+yOM2aErjRhy4Yp0ERlg04atojJjUybQoPuBPXQ7TVTqxc2lZKCbGxJ/
0IFZNNPsCCXWYbEhsZe7xB8+/aL0Cx/18WIjvOOebVNi/+ooenXvw0VGjCnR6k6e
WeCBmQCybXrsbiaZ5GtN9OB7Wy3NVZ0TlHWkwraJaL2vwsjCHvp9DEP4ulxfAIdt
IcG19i0y0nkPeVbZJ6jeZfh57SyfsN2gW+FUGfv4uNZogV8j3tV5tZ46ucWVT/qD
Cg+1xZy4OAsLpfOC+bB/LEiXJy5SGwR4GrfoRVJPD/EN1n3ZPBXzHgHVk/irsyWB
s5Z+JiynwqxHxmeMlGSLFo0TaAsN561IvKkQuYBgKcja/0EE+fpcIEZXGAYeATxt
Gzj6GlG4BPObJCKdOx6rlnKlyPripQwt2ZxY5p77IpXkMPtOdhl6pPW0lO/BSrdo
rItc+6g8I5BKNQgQF4FMli5dZK33JmcmBKoDJYGBztB6X2RKfLR05o0Fd3sMrOEa
oyB9jKp4NRGFcEGkRo/+quUK/dEU39XIHOsL8+cVFWTn917urVHRmZEzxM6vjUZQ
QfweBCE0iTb3Bi1jbz+Nb1IARhwnIGtdHZLzs9Zp21lnAQcT6zXNqDrUSxdtRdoM
QIJi39cZkhVGyiRj0ekAuksa9AUKvBFFVVdj/6tNKLqG5Eo0Az9IopoNc5sPgi0i
luQ6Fqv2uhqvk5xI4BmQmH266MTXCrflZqFSDPwNJsQfgLYob21DAkD47o9sF06W
p3JFdaKqNCb6ntydMIaOorQxrMLLj0JGBcsV+hMn/USaLFZrGgP3O6Ns64zqDhA6
8RU4DsQwlDQVExsPaF7IECnM9sBVpy8gr/9qG7H7wig+Gzjd2DLp3Oh9BMmUG5cI
PC/onn5lxJs5AZMOT/hUx6GZulRhmPlzHFmRTKtCadSEEbfa5+Iaalcq9B7FTq3s
PVndfo5re34mmK/ZorQ8gbs/mzuN2zQDMyHhL7zyqaCXMA150YDkyl4rYPfw8tyd
PkAvVvqlNGu5rzu9qtBOpdA/uptlgcLxIBhOy0WyZTv3xn7nFvK5ykSuXu2vGl4a
PsfE7ZSZSnH7VlPAy224snmVsknIpJ6qU5pgqqRLa7+QYbLrruoIbZwbn3eg3mjX
1+D+j2IKBado58L8JW+ZsiNaA6rZmMJF3rFowJRBfVUnnKQ+iNtGrV0afZ3h0iOw
ImGeln7puvReguYBNJbV+fS3Bh1vJGQyi0tLhGAIAbT29gydbfsObdhRFih8mdhr
tfwB1a36foEyEbs1hcSCn9IHYpj0MyfEENBM8/dkFvA4uhZ+e8nW83tQ6JZwHFPw
UE9izb3r1PE2aR+3MIzMGdQl2jLTLpzWZXS5mDa0LHfo1wy7fJIu/Vr95pGjxyQU
7LM/Q8JO4P6oAhtUHoMi5Sgsnz1zzqZoTCknCDsfUm3qN0SvxBR/LeaNJ47lKnma
LNnWSQu06hU3N96XycmrTsoeQhomXBtYTlPMc9W7oO/0NinSghs14GrPdBQGrMC0
LvOIheNf2pAQj6xUwkGplYRx0p9pSdtI9WV8lGHAjvidSYyVxu0SrS9/sdqKfr/i
mDtAWnIpvORh93MP/hRgnNvhTT/P7sfhE7yh5ox1SNyeXoHu6+0WVSYpYha1gNOt
qDCIiT9cCKxxpr1WK6hOKmztfT9UxQ5AUCd4r0x9OKDMObRIQgrx53JPiP2pIqZg
kYUuw+eGy7XDRkWoDJMU43gqCvtY/Ct8yTHDeCKUsjIVc9pfsk4rmMCrFGgCOPV9
yqmrmUUeQcQpLfOLJHC+iFv5Ld2ctLUf0w8ZUc9ulDoqYjJlWokmWGdeCjp5yAvd
j5Kz6OO1hfAaHPo0TWfRG4EvtbFch866/q04IKqcKT7ftQIckyNLndTsIW16MBI9
L6jynKO9mM05X/THW6Ga55cvBaQgBadHwWFSDeiddZiEYqzuhahM6dSYlX4qR+dJ
CgSp3KDN85nd55NLV4epiXQEn6bL7hG5f92kjvcZa+sQrhqO0WZWsa41YWsCgyeq
h4R6zz8pS9K7zfVZQJUKjaOYW6JH3Y9K0QwEicZk9GGPLewkmQKLXa8fYn3rHVDd
qPHyaBNH6ORF5uNoXPr3M3QhAiniRarAHgfXA53wf7bIWbk/grzDrJy6KSDYRcAZ
IXW3AQ2z49+7m2gqzmUlBWZ4aH/TQMac2pPWjcDmON3P/GcpogA5OJMHLEgNVSnf
16IgAIpew3tdcVh9lsPgv3ZjIaxr32gT1YguwmuG9HRXAJwCzYeKcA4OsP2/FZoZ
VqmGRiOlgnoIvHYDs9GuaEiJoEvB0/2pIcbjEJUApppan5VEI8cNp7uVEQFzrJLs
Ri3uzQwmjzkD+ml/HGaoisyBFQp8AKdwLr/vIG9uq3tgW3OHsRNgVe5zP4FCPIeq
ykakKeDxrRXUejs8xFXHkdy3qNqm756RUWvybd7otUrIb0aX5VXPKWqqYlj5AbrI
1591q5WVwcXZKZUzgMunc2UGis+8ERb9fQgBzZOJanZCJv4tD+PU30uvZETujRIh
7I7u5Sr+/rQJjtisqpFi5G1dfgqHVh8zaDHBs+XgDCHNtVOSN3cx6zoOiHIvvc4Y
uDkuDUoiKNSghnUlSPTaWFI2db8wN+5GYNJqd5crr3nDs/EeSVKLxdm45DoWRoue
Sm2R1UtP8WQHUmocpgCm9lsJPwCA3pVH2849LaY6ccx+6Ddg4wCqXMPYOds+oDNc
MgfAZAFmYQwMGyksvYPBL7sI1z3QwMSbULAkI9bSgZK0MKz3JrgLKGK7KwHMgJcV
G0bloL7We+yTHdj2YL1+sf5q2MPJMyoNlRtCsjUnsFvmIeXyKXCBzZQZI89SsRB/
6Omewtx21yRmfLQKBghQCJfdyxOTY7CAXYmrd1rpxqDhoG9+p3VNn6kru/q0K5fP
rsMHjvFbVWhZm0LBbX8BbIPYQwplxZVNrMucEtCX1/PrIy+fCEPf6J6VqEdHwcjx
TPx3q2mV9SkYQkkXxgCBDuBt0Cl3tbboaIgeOPlODNeXUT6tzTgsfKgezV0JEh3w
uYvLZprG9ENxh+1NpRHn1p3znRWvmkU5JPl1aUK/7jbwFjweNoIR+IjPhwL3At3K
YblpbpDp8KiK1IVO3umZk4wu1lOAKvgKoLvYqLzucZ8DUbAgTa2XLnLdoQBs88jy
xljT/ndh4ALUtNiolPcPcNqkGdeBZE7qhUPyGr4Zo/IGQOeVXAMBJVbVrRgTPK6V
bUzoBBoCu58kmIMsUBo3yHqirKIQRJPlX9OBQX0bZmQM7yE0+PSZnfx+vYIR9knA
zh57CTM8SwNKJKZmQxAqgNM7Gq6/muiUAQAE7y2i65XjN+BnJBfyy3n/EqUfR+Kj
KvTVjXJHZnf+4KSi94Dmt/aGgQRsa0XZjqkytaBwE08lFHOwnLfGNrsM1gTIgMYn
2SQS01oHIBRe8zTgBvb3SA5fvGFxc0g7/WKjTWUEPZikwvCWhxNVROpBkBUaTAXp
EL1ui/iWkNc/Tmanlx3nNTHjiGcVzeVAN3tsKAcNu6ay9ISFPZsg4Nsk20YSDXLo
iLqUEPhFwxDQ6eHtit97rfOj/mWn/dUdhyG+tZXcp29DSs36Dhp3nh/AmNfWm2FS
3doobyGjLWaq1Yn05VnBkFDogMUbMUuvRVtr9PvFCZTAGHKO7Sn4SgrdBrf46mSi
DwhBSlYr2WOt5Fz0mcxUxKYXSsyoKK3PCzo3smvpHptd9Uynl4yYpyueXdM+7/Lu
/Y+eywA1LtvvwiigzDd0A/EHh4nEAJVkrNMatn8KhX+wl7HuJZX6kA5ukMH0sBhN
itfniVmJutmTbdC0T2eB1iIzZkugGo+WNya3LnzMBFwpOH92EsjxaeA4kjLtm1Mc
OwzLHvxYQlJA9S4AQrKSEXnhNuSfbiwB+Ah2KB6P34IRCbdSNS8YXXwJsAO6o26k
pXjnoFncixJARg364zwT1KzwJ66Uv318V4bi5yKmCByjXYBkGPjALsnF8052tjkl
7YKkiD7r0mvzohift0Cpyc4sU8NgfSaJSiTnblGOSlOWXqdsOahWVzgVCDMRo3eJ
xZedxdupAVf12PGlx6jkn0J5g3lJ4cnxz/+6l95bCnsHYIuu21vtLB2pMwY3wCJT
hTNeeVQSq7R/j5mo9vcnSSNWRlgleDbBRVQ6vzqxFGj4c/zwlbKQLWqQrnfD8yU6
zqRViKY0mUgxgewRcMqFslRWSUKbzfcBiWosERJlqEvN7JuEA1fqa8RxRW1GSi6Y
1yP32qQXj3orR4Dr8kdiLY5bVcC35itdFnZbdbDpR2l+nTC3rNR3tV16KZICByDw
H6ogS7JkSPzW7PEcgYYlI1rLDve4zPU15A2FEMx/KKFR+B2VUExx9Gl7UIQiLd2Z
x/LMEndfa6ShEOeLxEM7VNEM/qgyzUPZMZb26qsV00R2YnBNrqQlixFiK3oOe96s
GOOAxLJ7UbWed9MWA/doVn6Ud0DLGMJdx0lg06SxGAdLl+KFbFKgCQbG/vWc2mtz
NXj1fiHw3sKY0uTq/kohDi77W5wbCIjmHBYiwyGPWSlBhdrXryR9dyzyMj78t0Cl
cjjoih2nYQrg76Z/QzIMCDf3HwD5bMeVZvyuwTa6zdkmWaiNFwsnABkKh+4g1R+c
EBVL8/QZrL2Z6YdLu99y/lk+if1WIVVIjgmeIUo58Rs6oJwhVfM1pNz/SQzhdxnZ
6uFx75En/Hox8VAfG6S2teSq5hHcCusJeE+v46WJtEEVugb9jFdaK60132NYnfNx
6PMOs6AvkG30y/Pd9HZb4dfyumoePMTfiEB1SFkQrUE4tPDsg2ree2afeMVH1Jod
oCKWaqlOswF0l9kKlMbQRLTx0be6EsB7hsHhGStpchs2iY5mKIlhBKa3yWvz0XNB
E2SMfuvSlDdSOp9KYWk8hab1tEPso+H2sz74YytxANjyu0/NHXwLM8UPvOYRsvK/
GrtfT/z6tbHXR7BLV5vktSb1tGgt5fKrZGrQo7sG7p+y68F0wRfcV7GAluGPvKTY
clf9c7wbJfsLllZk4GpTZ32kIag4/tnkEHY6e6BwEgCaNmNtpjoq3fS6Pijuh5Pp
U6cLJG2cnJgLIZ+pU5ujxDsFREiAdu3ftY+qlHfTnz92UJgsARriotFeIM5mJ5TE
ZhEPAVMhUaPQDzLCdPX6p5iXDzIgIk8IVr5AF3IoxU6pH6CucQZYH/ZwpQbYow2P
X1kCbw9ZBlJZKqRwhGiwUB9xMMapMlBCkDVPBB8JgNHGJ/UGHshR+hMKQF5Pj0+Y
roiGcDxQLPPkiQ6JL9ncxTsXStOWIbXNfH9m10s7SumczB2THbRcmWZWXkk5CWE3
Bqgc5+i8GHV3/TA2bz3IOLxQjbtUKGzfGj/xZ+v9lB6W/ZRhQe5/2AbtTI5dlAWm
CL9x/dHIinrLEKSGxXcJDQwDNpRK6qjKNRAZLi1xE0J/d5reLFIIvV1ZfqSFTMcs
uVbddghwczKQsbf5VYffYC7xnkTEoui24wz9ytKovAvLyHCLS8rFT9If7nRuTb04
Wxrp9JX5peRcYwvHckMXwxj3wJTdrkiR0nQVXbm/i8VjiLGTl3RVgCO1dWcJmp3G
s9PyWMgoYA11uIUfp5XxEf9KvYSr8nkwO2U54UuPtJ4FmaKQETcK+v2aRjxcg45J
fG+5ySIknhR33pHaAXfvEkF7hMCwaYz+KZt9r+QmIJICj9/K/QGqO1OSghts32US
X5U1z+TA/j6mIb4wlp+guXKjLB1whLoI1pfm8uUbq2B5giMDAfs8RleMyhjUkL/j
UeJRM0RuqyrIAViPGknna9eYpFKvmahXc0h6wn6DJY0xA3vC+YYSugxRK4gFp5ax
cB7N9EzXNTGA/GsFaAln9llIcQnRzrkviaNjykixGYUQXOV/zY7Jcs+PgMKI21Q0
OEABGVxuL72Xas+HEOZyCysYuuP1y7k6hveO8hpuUGrTVxpt8UYrYx7WT7qX91/o
Er6+XEvbjGy9eHFat5WR7wMYYmImsWoXhvataO5sESSMpchohbhfBbPwV2v3zbGu
mZLyyP89yegbzkpB0XsZSqAaEY27zvXGM9Ib/2AdWqK05o+o8w7dCsORGfV5C3of
Kw4e5taAPWAoPq2IiZOaSdey64/JV0qGjB1xFI7nfADglf0v3I6uYyntnCY9hCsC
7uO50bHqPlBabxjOX3919TrDyXsUevkrfikffE6J7GkllROv3TowTZ8YFT1cE8RS
T8DHJVA6EB9UWox9ZzYj7d1a/a5ax97hH47ge8i4n2Xp5c2j2Evhm5j0okt+YzjY
PzVIY7rO6lLM5ayWS0LNMyvD0cKS2EoFEMMFTr5Y+cRTnHAafeT10iGJdduIEfYz
zREGCemOcm9MCFRJAywbtpafn2EeO9GHDBYqNbbT/5UEK1KNgcjbtw+3oGFHEGB9
qUhvPnObq3+4phrto1rnwa5gdJBxGv31AtiIbsyLfYjEKfsBKEjNWJSHqBA/pB9t
PCr1H/RNYPmAcF36slSazKi4sGewHdER2ZDkACbZcsNwL7IUAudzUEQI6gUSEinZ
+xSr/WjUPnVDjSTET5B7SKDuPoHJYs9LsFQAJ8LlQ8M01+bA5tY+TtlHGRDvgoVF
llxo5B3WmYCE0Le8wUUgmrs2CCdYURezXWPKceIvBocnMwZOmB9I88EDzBtFp2U3
MDMwtSgFxK00tSmOJCVG2G9HcwWbzl04DWKXP+uFLahyshEfpLLf9yh0c4PmPzGF
10QiR9ixsFEvW5Xb+BJyjSDir13LjO1nnNouTzX6NrTsi6K+qmcQEf+WJP2w7Lg3
ho0DzALuQqqgqsiNyDPsB73nsXsLXnjzmx3DbLj3VwohkUygm2ZzEsWeMWEcE+uF
ViZWJGLZFRPHJjCK1a0dVyhXu8Blk0a6YTNSVQmVEmbdZGpQn1ZZyUt+9nsaHx/D
uovS7lXFF/6zyzmzH/qzz32uwTrRpL+Ze90VNQdMUysdmZMeefGFnoP0ZFAkyhP9
9xdZZEEvgUkMV8sNGCp+EoFx5h/IRx8m0h21gn+ysiwn9wKBO2JXPC+Y3wrhMCsx
Guep+uVHjnk0zasi3eLU3OfHWCMf1wpNVtvHZPAPYd5A22FFOuyoKFv9rQzlBioX
zokcui4dZJhxAHLI6KgmnovsG8QnQYvwtRmGcwqpX1u2/QUgQG+w487IkQ3T282F
jomLhQTg40SCe2H2UH3N9m8jdF9qekGnejRofaFCQ1HZ53EkCeTHfF+ahPojZa+S
K4/ghJaolYHRCIsA0+BoSs1o6D3/p26ogUza3vNru+9dQnO8hvgBK2kcZ9A5Bke/
Bu5Mu6gZr6mYb1WSD31Kz8LL5qVDlZKC2aHGi+AbPARKmUTeD9qEXBX7xMrGpSOh
lR+clGasx6B1tln7P3XsGQLrwT6VzBNmwlRXj6g5bhrp9c81MjklvjWvzR6lsF53
11eFPUCf5QNdxa5Npxfq3pbEvYPTj0rjJL80brUTRHoe5KskhMP0YMyKc4AfkEgZ
MmI3vSLuzcOLpm6xbJNPSa3q2PdcUr6bju5Sr1TagvekLH8/JZdDsiiRJjBKmtvb
x7LdJibZSk9yBuHh13RsgVE2X0jHixfh9TO+wZBHkzUlKMvSD5B56j6C+GwpWsCh
99sXVRQpk+KxJz26xKlft9TEsYxZ9ww4oBETyT4hjSSC3UY5R6/AvWVRjIUNQrWW
21cDijTP6CHJ7sNv7QosYmhry0YqqmfpEDvxawJ6Xw6f9Cb1KiFJBl6E8NUl6kct
BaUTQXA/2kfzaJ6uFj+fXZ+PKMoJR2uD40LHPJ8MvkYi+oDm5H1FooqAtFv3MlBg
AV+474Jp/q7zebotQV5TAeIDlLed9Fm5V75Q3EzoOeivnWCqMDaixtlWdRIVHyNt
v5B1GcpRI93FOfaSsdrBHhC0ilzzr3ExMS4RUDZ1TDkjB8ot+0pKWXpI8ZY2Sm72
LV1MM21iA78VIKBtZmwM8VVSDPmdMtQGuGEKKeE/pRRy37KDwgB8QnYWpuYxpSGn
tiPINVpiE/CK2C1Aqnqucncg+eGmahIs07fqY9MC4vI7IUBDRvSbHLy6/9Md8QqL
OCsZs1rCTvRa+zTguT7o2gz2t5WgQOvk0dOUbFly8L1pNtq+MDSeCWj73fbOK7G7
yNdGIWf+whkpqJ5aVbTtuMobWxuUfgRsNImbXZ0pRKpqJK13gmZca4aGW5xKcE+o
TDkXXxTYEiMPh28TBv931Z0s2Ubrp19ghW4fwmipldLs2olca//r5Z/c4k5JkOef
OKlzc+Vqk83WVWS/9So+VJ8XhQHv8bQa6DbbVitCEYUgok25gu16Th7FBL+aHEgs
d3W07AxWS75gTlF0ribzGOudfKQ8e9x/xyiqjmqoQke78tEGXoa5KWkJmiokyZ4E
Usn8b+zV8g64PdpwOW/ONC3uIPutEOzieZnDqfhyL4/vtOxwcSp8w6isktCm/EpR
g63os7loCQZKa/ilOB+QEFridqxymQR7D/Wtl1ZUmLctWdkvQKSP6j4aKu055f7O
AzizRL5Pxrh8fZ8Y/WHcoImPvUkA1w/Dy1FiOB33vEXtrTwdyCM9BXyErZPznBlx
8Y4ykFwUGjf2Ga2BzggMxtSqD9txk7d75YQWi2Cze5O7JjXngc2SkjjqTYACnra4
2B8+YM0tkZcvOARxDbiKYScvoIXmpN80/EfiiMkgA0+DbTR8AJCe9f7FIgZbE5PM
6pUKjQm1XMaVZ45gEpQZhXx0o+7SRtNlSDXWUkPIkE8QGaT7FrbsICLWV15ggD/V
EIf+DtVDJ6GTzQklQLfbiiDom8Bwg6aaLixpE+iQ0ByI3iXD5y6gCq9+JASqHE4G
zWAaF9GJyl3Jja3iuk7uGJNR/ceeA8j8Hk4L33vBMtHGJzVMLh5XDpjwpsyc1N5j
+iwtJaE4NjoThFptB6vEt557Pfy3aRujpi4AgZf49ggZlatMKRroosww0vVPKLgA
+dh4t6xk+6RcSXgUKoxIUxXVUJ5GqrBluj2FZCd03ji/yA7/LmrC2gecDd1MwGzs
KSiv+4NiRv/vx6nVMp5WMu9kqf1HhzUwfnnaKGTUScVITaXYlS3i71ELcBQR/ysT
8r40sjnOWmlrmJIp/3SLKfUrzymYY+IN4LtFfW+2h/J0lSrscgoqQcoKXWesa6H5
4VB19rtXVksX77mcnXCoFM0La6Yw6CsxAenj1o1tYJgao1AUldlTDmTnXUVmnDvb
I0rwxLoOKl+EfP4CbHoPuYPY37TBCA3Lcfqk0MX0okByUOkC5GaGdCBemTKLCDqi
k3mhTqrIkaPdkLCD6dPo/u3n2yRgdEu/FCDFggLZwpt4jKEnDKGwHu6CuItNocSg
PiL/eEoKJiyVCAhKGFif8VgibsJwcG9XQqS7DO4rNzhIZlmz2dRFtgamLD3LHL3R
+/pXPy8HOlLGf5PcDzoxKM46ZPyuqAaS2hmNZd25mtsVsUsBfhZFNL4amZ9DMHJZ
gBXtrOrJl9Bf1Q1v6okXSnwq7QQycbcYrNEeOlz9lcJeHed76YDFvqYsK9bCF3PL
upzoUliI74AsLNytu7q5oGcqeU6GU62oB/2+YQvB+hpNe05Cg0Emdqho6TlMMbIC
lhn0lNaNF69xjrz2HuU3vHO1h6wwQ+O9Rk0Lyy+oMyTpDesrT1kpvqEUcoO0vGA9
C144X0zRmX5OZdc3+mPJ04RhMDv8TD9TJdmYT8uPuZNaQ+kjXkjdpGnxTH+eokY/
wVQ5m3TV0H+7lzgmtk0BYQ8iQ3x/Z7xB9ZdHvsGb45nJS6n3ymfGBBjPbwaF0hM2
OIhqUYR8vQoRgd4pSV8Vmwd5YW5DJC8qfIrQg1ymBxNF/VWLU/e/q7ZNXB1Q7nEZ
RwRuSBnROevmhj38gmtK99OmqUcEIkw1P4cPkEFvYHasmttvLM+OPZOXamF5Rvqr
DbOgXJRSxhpKnQ8h9qpf06gWM5KaBNXyv0E60D8AOIYDNX+DIvBPwF5dhOaDhEYS
+fPtVjVvcZEOkFlq1J5fT+sirOlXRjgQtRiBtYm0zQIeM8Ddh2MzG5kW1Jx+0q3o
ktarGFJ29CG+MFaz+FqA0Pj2o0srfi+Pr0DYNkZvUXSBQa9djqkv/zfhT2DX2ELR
e4QEoUMAZsSvS7cXY+wTeGp3ZBZrO4RxQcNLDtsI5y/WKVAaFsMDqFVamdFZ+iYm
z3/wY6JM+i+RxNDhmIjsyXIuEwObgTra6EUOd1XMB7BIan/Yza0yMIIn/txh4v1L
c5l25vBpEJ8KsswvRYY0or2kZCEea/36RaMB31pYICGzY5IeSGARjF10+yA11l+F
TQvHorKpTiqhoXteMCRKYH5pX2G7S9ulj/lbjvnpJ3BoppByVFYPENMQnnJzN12Y
GVBUlyOGRQ9U2lyegvlE2MwGJI4/Cs41aiSbovyL9AsfEJitrg2V7s9mNGx4iSWo
1P/Fx51NphtuQtwaFrIjmoNm+OExO0EyIsOkiA+rRVtPS8xTzp1mo1jYIfTulWqR
7bqqaTf1pvSQk8zQKnnlwHwpx/05Bnc/p5kgNpvqoWWC8PrdBhloS36ch6Qt6qWT
aRnKNFiOARkdXhj4kHJG3kQIX1UAz7OLoPD9nIQB/MPpBQ8L+5Pnq9jeDYsAADT2
ZaKeK/BHti7+27khmTz3W7ItB3691pRij/bnIG6OpewUblOUMHYUr/wWqalxHPNn
UNzqIsIi3/T10sJMspCTt5sIyX2ODMxFWCeewtw59uuwmyL1ApG/Vi7dQAp1bTid
pKh5/4u77bJAaVpTme6J0nEwQY3HwBNfNWXsWc31RxcSwWenJI1OnYU2iKIND3o+
aZ3esOG+/V97csWNNNvlcs37eorzkyBMkFKF3ql541xlMZQoZqIBC9dbkYTetQNl
H5ULxZjqa4pbm+C1xz8zuoapbYPUE9NHwvvKrCTTvNmgdbVWlpBOW2hKb/tgVOOH
/q7GLpj3z2ArGCU4IdT6+/OETCpMHFfmMOAe5zcrUQhgntLN2jcDaEAFQ8YVS2Nn
S01y15E2YZUlh2EOgh+/lNEj2sjyL5M2OqTzKJ7yj+qdGsvSL8kCb+And+j+ONTP
ZOemf4ax7DHPiv8grS+ljTFRF6VPdb4QijUBwgxZtOlBH2rLtnRHSsK+hhhmalU4
PL+ESGyCXdjlFtXYQJ0YulF6irm3BAzRSHEJGMPrDuh/KYW0Iyn6DH4xnk9FaJY4
vIPA9J17ra3ZZCj3efPPLHTdTFOQC0zI30zO2y3Q1QlKkaE4YTxlkyZyRFJQzWmU
4uGCzORIRwEfUb3FBp1Gd9zHf/CczbRWAamtUpO+C1Ztt/5iU52Yy+MBo6oivNYT
nLq04OIsTmnc66afhik8wSVMld9KGRiKBIDxk/FCLEnNwTrmkV8aP7owKMg8pNzj
Mt1k7ky810znSawqL2Mh2VZ/T/16DUlIj5c6NuMKSz96biZHHTzqOvLj3MEM7HC0
szlAZ+rzpprf3qnaMU+I6G1vYFz4P67vH9vy4okFoAyF/1X9CUcZlJDD0/zc/TSA
YzgsN9+qYCwlwIJh9STfSI8OmgEgmEf/PdxIkAyZThvlseScXlWoh/COI88W/auS
V956mvt4Gfk6AZwf7C/4TJbqTFIREjS4X5v9wEwBScsAca9ub5NpL3NB//xGT3dp
YlGUSyPWOfnTw7pwfD7iv/ec2Wv8DiqPjq/myFR0YlUfHP3YcgOxpJuQQEAqCdJt
eyNa9SxQmkUspjskTeJZVK8YOe5iyKVIchaBGYpwN/b863/7kB2u5EqN/TfRM7dF
yeM6LrmaQjkIz2yMnV9KYO0eCWNdTEKmWFCJa8AdwNKxc81keEX/6Q5Swk2cR9VU
ePUu712FarpWBZgvxtGFoGEixyTpLrTnsDZT3g1Qwn4i5V+JR/3tW0OKlNiaVJok
nO+sd8Dk9EAYrkkM8Gw4t9b+nOzUYNNDd2xo9O1yqplSvwmEA9qDSumko0zKkZQb
RL1VBUTcdJehSUxkR1tiBZAtY+wjHWAEtj6FnIotIZIa7obub5k4iyUp5WGiBGNI
iO8QxJuwnoKpfUrMrPZVkJLtwfqvFnpEcVu4Eb2LoE9v8u1vvDAychA0dv5ezRKs
CzrPKbNOM/OCWhKFdVqEEE1GonvgKgeJmSkHp1m2b7DyFWireFlG+cYUrDuVi0Zw
ViMdTx/Yyx2VBRintEPX1a2Zwp4pGrK94vaDOWUz6bHLYtfJRQGIAGnjdJzK2gUe
cA6ZMqoHb/6h0wODVAJ0SYSIh/5PWuycq8jcJoxcbSqGVxLdS6t8niyl6/IqFwq+
mTRCZLUvg7cU7XBLYgvOPr1LrOEMQ2f8xOrtjRYOpV18FvtJrtUxwEfeVYrFusyz
b9EU4LVV+GpryiSKcvMVKaaTNHiZ3Bj2EnQ5ZcLoTyLFhV6xZg/zHELBHjrESKpG
PNTseMyekzM0KY6oxPyIaUF+nnv9xJ166AkHxZCbBbgtxJu2sGGo/g9wWO42WUay
RkVNUNJ6obHKXAp7/LCFKSku+bC9xoaQDgk92+FSyhXsThFu9fqPQur+Ix5UXtkF
IBxag/C1D3osAFbpvM5dLwtR2Vb8APT0Bx/1RtI0nsz8jyW163zheXUDCVJ3l2sk
sCJsuTjHXlXc8dsFykB6810Ew2WII6NeiY+XyIMHZOCOpbJ7jHbb4FV5vzZ0cDTI
gB41Am6npyQO1XrHREaspqKvY6Kx15fnVVBefMg7NnL8yXbSGr84m9geYZf4gIO+
hD8mMvP2DJYokMzjuJvljoNbP+/ER/ksQcUhIr2HEY6QRBa8QnLmrAFLHS+N3eis
CRfJzdCQPtPByIITKnnBwroQrdO64/yL3io7AXWn5PIxMwjcxE9b8oaUIsFe5QQf
4S/7kVHi3rgLziTH67uaE8yPNMkB9HQ1OpTMDwGUdHlW3oM4QmV+evrvSiprLAdE
NOYVNe2iPGh32wESOJjurVJyluk8rLjugqt5ZYtsFWMZeeprmf+OcQ+BcHVnDor4
PyW/NdQXfIwdsRjIU3HUYnS+XEhKcpDOX7tDs/t+ZJjVTpekqYDjXiuuIrGC8eeI
JG0v7B7VqGINtHaQhYHxNQkYgAmNBIBzWPRCbSxR3wx4OwIaXOw40xr4Xc1SUNtc
udZPSqDHkZIc58e/v2DPIaloKRB2WSqYS63hBt5xn453lTKSTKLbhWpmS94iUYfq
FvT1i55Vd6sMuK5BcDPu+UBI/Wt8fmHa66wMo5XxieYXWSnqvEMqr6/F5fOpBXme
wZUCdAuKIgm2BMnwbuGk/bFkNTfF7H2N1OOnOYRJpecv4rqnf+3uMsHAKPZuOtQ0
e6MWs6zHQzdRfSP6dvc81/Sif9L+QA9IjWAQ57q8KhctOo1K2D+Q90gCB30Pt8px
8h8kwJZjf6Cx0IJ9JptJdGNfn1QQa7myOr6StGICA0Z1nm43gMcOCenHt3MhxeFq
Mf9fhGNLkhQiAWvqnWIMb88u6Rh9amLrr2JfhevKcSBbcArTEPn2XGYpn5/lbwAd
3SvW5cev/1Cvup1Co5fkmnLFxCY6a0xY/XmVFGTKUKnQPFKykGontF9sHW+vFDLy
0F513dRaJRiKrGRrirMg6/+MEGORgUGb8EYDyHcXKLXPNJ4bQduvQCQSYnqR2rH9
ogku8nH7JfqUyYR+KnXu0jfmeNMXk+J5OnZAtnjiUx3pzjjYJjuxfPI97vuz9P3d
SYMsZs30x92s8Q/dN8uZgyYZ1YEWP+aUqiHMjvvxCR2E9YICYr0UVhB1KY2jxRdF
XFVsMhdAy2qqEE4q5cfDGUCAx3hE3Ym8QiZUALD91Hu+MRbCziordnbWW6xsWwu5
anbI0iBwfr3ZHZGUKbkolhgl87my1QaOqZx66CrnIXKhXLiv4YRHNVT+1wEL6UOw
+pVwr7ZAOeItPC0ZJLIUZXN3ixSQdHyHT9co3F3J1cUq4yhwTFtpPejMmsCGGzHT
He7XSrrugsZjzLtZW9wNve6dE2OjDNyoLtvKDcFbh5PEmbO6OFeF3WZO61Sx+n7T
yEZFIm+eArRBVy/Kia4jKBNGZMmoI93JjLfLOHNlmSRL9UvijZUtCZtqQRRd/AZV
omXdzbGYERTCcasoIaPIUymZgbp7c8RmVEe9bnabeaBwZ1gXbQKmrcXKH1fmdpaH
+pGhHMgJrildJ1X9o1WjvMHhuUxrWMcaIfNYlPoqR6ALuMB0REegxixuo4Hbp/C7
4yVU8TZepGRnuHJx5RGdrDobpznRHhXTEDiRxsP29CC7GQpBBdg13+NhsoYDy7YV
+rfcLLDzprlo5+ZHZ0kgf7VPfCewPlGOc5Pf1AcVDaJJTVjq5eM22zzb+fkiyh2N
N5LXHt0LIr7LdK3cfIt1is07EVaOkRBTRHVKJlUBWnKOAxn86omVliCrtxcLedDy
Fw7kFtox3kPpmgn0rnc3karorAKdwYQgR6GSF1IWCoDYm1wp87FsrWg4wC3BdMNI
DZbiJ6STc64ln+Pdit03c48o4mhi2dvDnFtE6WDwVdsOMgmmzexyHN9OEOZjfbJY
IkkIyHtJwawTVUn58UeBnP7xbntApNelSCRVKnccosWC62OH27LqUoB5jELFMYzE
Cxm6QC92+jXvJcqEYiSKBJC263SvFf2ZoY0bOJ8NRjHFuJaTw0b4yIii0H7o1giV
e4YeiM9GBny2FHTqG0+Fq37N4+Ijj0EE7Q5hodt6ePxlonUXcR9jZ7Fw7Clg9K9z
vD/nPZ8yNfrt4LW7Kf9nFFznM9ZSqR0K91d+zT2+qc/vxyPJh68SIawLR4D568Gt
57IYj2Or0EsTCxVjd7dKAugQEU/zRzW2YV9nLLZZJl+pTk7rMpE+/yzcWGs49GqC
rUauF7fuS/owr+xCIBvB5RMQu3/OI4gnWwmdTj1e7T/u+5ab1Ar+dlCINr0k/yF1
QmvgvXMIymjdvFaXdJ8iJQR1pIl2RZoDSDmwa8ia1YNOxvjycI7RmGPsnmCi4yR7
JWvwqD10+cPYVY8KgMAL3bp7elohWEmojX2fc74+FI4qYXf/0pZ3Euab46opgsaM
hX3EbFHK1IbddTxMs0/L5jPeZcbLwZv1x7bav1zUVva33De8fTIsAZDbLFcUc4Mk
PBzzIZHwSOskd3MDr6uLlxHgdmTKOYwHQGOQ3PiyDKv+5LxqyTrKkeBcBQ+S0nB6
VKHwMmmTHG8wlSQKl6UX+d/Ygflw3LZbgYNZlyq2S5EYk2+PXwyADm2eVIeQ7Mas
VL24zDDBu5av7mqxRQcTYEKuk69hgGUgpI/BBoW2hNKvTPKiLBqU1M+jj15h0lVb
gcbiwqTnkIZ3B92xQKnyDYU20BZ1SbSbjnYdzYvVVNwEE0sLMnE//10n8MjYhzG2
SSSbUgiliqCNAI7/zGFVlJDT54V4DWUBHVV3fWZQ2N8wdYtUxzmKNg/uXvkixeMY
M8WiYUKEA5U3D5O0P3LA1KdnFELu6ZsV+L4tSjN8eFF3jyY0Xzv5DWQ9b2tYDQkK
uwxlYM2vsgLfpcM2+Higdt0wQ7ZESLlHbraw5t8wwB2obeczAcmG05p40iZn6M76
MRmgPdiODASXhoJCxZdRPWRKgsv31FEtYny3tCNPh/CVS1fKLgbqbtx4lrJU7/0e
OiJMpNS+S/yeXqOz5/IIds2WcU4Awenl2eSFA6Aw3dcKzeiPC/KUW3PAXwvvr0B6
fmTL8Qz2MmteqsHFbEIHjwqZDtge3b+L9NEWRkSIyheq9G0pqlctEp+Th1lQnmIr
mpeimtN/a7+AolyRP9xOJ8ypNaN3Ek1qQqmfy6rXDtlhRxJg0MRCzmvEfFpkPdUJ
axirijbgo3SioZaErMP1h8vDlH6YH6dxhvlFbV/qnyE1SzlzMqp+2R9sUMgjt1Qi
meeXZsA+IvwYXsnLW4X07g5pJIFmN8KRXq5GWr18VcEGqPWJwS4X25WUslLcTzLB
Vx2eACxShX03BpSiLU5k/ArtewFsCVXuvBHqnzTFNehwuM0FHy6ptTzn11BoTODC
tZXEm64OR1BqSwkP0b1flbnm44knXmVDFgFq2xuEu78NjGM4I/PXaxdxz6WDeqFH
WZjbYO81t+jz96aXDXADGuTm04TxhrpygXvplw+taxlrf/1mwHFbuW/ALhSO7Id0
u/QhFVK0H80oKMCFqf0D6i2nwYm2pDiuEF7KSUcxW234bY4iWs9p1zxoxy34H59Y
e8ghIthBkNCNQVeK6xL5VtWGAnKIt2Zw0iJs3WlYEKXMLq6nxKCfnjjaBpZRE4c0
AGCakc2SEff7pesFQXt4Nmj7dG5XQyuoTb1ZFgjRy1ycqK2z6TC+EhQmi8hJhknf
FoffLOr9x4RvSq/H02/xa6z3iEFjW6SS0p5gVzMAopieIDQ5vegsbaTwBlhcSmJk
Dw19nPn36mD8XnItrBt1Y2eJBRm2bAmmN4XWtyyr6cTrz2SMqLZ5o68jMwqcXcX5
KO5Hy26FWlBDILuBD67ys5GTOK3h/wr4ZUVCzT0PZaXN+ph5y9Q12HCsAHUs1jKT
F5dF34ydy4IrPVBaCuoickAcb3bIKSoI/65STDdAKYr6pLN4bqg3lMHhvnlV7nMd
Z1twqaiOa974NxYgmQGl+IkwYbFacG7jjEUTyv9nCD/LIPCO5OjC0cgP9A+KPd3U
uCP83ZB8Mn5McfXkTBVkhuvxALAIGxBRoOGpdEJ5UR7WQfjq+VkvNKSAGIPOMlZD
nEpKkM4cDsWa4UHs4XnhFEVkAIseHPgQnnapYBO6x9ZRN5js8I+nZFPo055xcmsu
L9bSB83qkUdq5dn6ApgooLB8X6vEK4jNLV4dZuB6ryXCC1wHgCSEK32W6wKTBie/
Qzpffnfb7nFTIaYDSED1XCMz4pjSHi89+FAGcgq4/h2uIB1WuzFJ4KIpy8Tb5VaO
G9BQrEGP5czM54wibCFq/jwIjl5nWlQFY0b5A48AkmvYR8XdTm8DCTCoa82ss256
SBcIqv5RFxpbG9dClfzz9Yr1gJcze2yzRuRa0ufW5fTVlNdGSRrA0YAwAhw7hiif
O75IigUx6wPS3Ous/9IEAoaiN8VPSyPlyRxWgCUQZbcgqtIeULOx+6kXi5nsg5Nc
+Zx0p36L1uuoYxLreXMju+D2287H95sdhnuBrVrtWIA4VsNBY7kW2EbLRdCu5jFr
O3/EelJxOMe2H2R+NXp+WwF8AQCRM7ph7wbGZ8daJ3xNDkn9lkVLuW0PL0TwpBZX
Ttx0ocem06RnjNJiXKqMy4c0NpyYDN7N2IOq3G00y2g99sdjcKHrhh4QrMyq+48R
4yNPdUhtXJs6Gp19SjHVfQJzMuDMSldBbURENN+nzwW2FML6YEzZ3oDjrdmnQf+M
Nj6mUopKJyQyRZJzDv2nKbW6i9v6WONAuJm7u3oY5yQJtkMySlhGF4qcxIIpyXSg
3y/uBXAYVuNO4TWwtd6tqJ160iq+317d5BGsdiTLy/qTb2w3p3D48uneWaxvJlM1
vez082EFkpQiJzQL7RYA/eJN8JGNrTNSrZw+6TUQ+/y25LioX/fH7v8ASLoM8FYI
wruSiEiuT4UgOUbAHeZIDwuTpKqv7WAcDyswZZv7awR30+9VFpewiRbaiA7E99Ar
VeMXpxVD+WUn9gVLeZ6Uusc+RQH0GwDYnlVu95uSdEmqYS83lc6aOQl16QHMwuId
3NQ4o+xDjDT68vk7duzZaRQAMqmqnv4J1pLtbTAaJphNGrdcWcGTn4l45IkOAoGp
eO3+tmBqQmnYAy91unoaZl5I9dTTO2pVfOCJUimckSGK+P7hV6yru+25p8yp0fH0
ZnpXdBwt8yllBvpXjzTEEzmr8iYAo6v8AJxzgbkKI/PBtynmPdqEtKBrHQq4hX25
RBdbuqaWcdvvgPJXg1he8J1p8g/TlOmhUncXBfebmRMchlBhnTxN+0/4x4mffFL9
tXnFZztNO8hzxmrGhE9m8jyXHBVPbhvOH7gYgCXmXNoCk+68aS5UTEpbjCU+RhlQ
h+PpWv5pp0f8d6AFDGqbNc25+5GOfW/eazy8yUbX2/8elZGGavNpETBslE9Kw75D
ejFOFwprS6I+YZTaRwze+1gYJAIv2CeKa+/MLKSxJViP2uVCEwdY3fwTvQQ7EKrA
6crQ5C6OHNqAjpT802Ok1NTEYCCyWlE/lW5zVM1pYH2rpAur7zXLcF9AS2x2N9mY
SEA2+tnESnpi7YbpYiJi7uDMOtnCtCudWxTpndoeLTNvvR/x0Rx2P7tblAmr4SM1
Dy/XRIk4nYoO17PCcg5zsqhW0YctdygQE1QKHanWnKC2/bdk//TGq+Vhv0L/RtQg
6ZjXWn8313yETUF4LffesRT8Ww5aZq9BlPwVI/6+T3aeDrmpGy4vC6G9z4I9iPr9
SOz56FfNbPuARG5tl0UEt3qxeND57FWSXdRGu3pPDRDrFHK1HWpCgz7yjWWLWtGo
ytOzKGTi7IX3hnA+nzA4hOCl8MqDeDUksYNTLHL2jhpESZVOCE+qNLJu2Wt2zheF
Kbz4Zxqek4BrDrz5i/wcPiV9nT1Z9jwwNf7IL6i9/db9tReZL5QeVz57OFkUjdl7
KHttr6nR63D3EMDIQmRKM1g5JfEClE7hMRB5uv+3fuoDnMQ6BSR4ld00BSjjq8pM
6vT5a8BQ4nAGxR9tHsa1af84ZNXtBKIuVnJzR5RuanQExf4jcpLShY0EAJVw2FW/
m8vYl/po2y87DNyTgGHSvou0R4y6R+epo5hAuPQ7lrrxFZ0AHRTBLp6w71Wusjfd
danDs7MXGfkBcPPPt9QmkXrtf/jlX0qyKkg7rjC9RGnBXY+HzmRcwAksaGBttiqN
l2Yu54/5LO5bCBkA8otdRWIZzkRPWU9xa/2g6fBvI11fTUHbwfxvoZMah7XvLmIH
C18HqMH/cIj7mzR2dUJmHunO9LS71FxAWxfdrf8CgbiteB2bcxHdEBmWyWB4BV24
9OUw43SLCpLKMverqArK/5oVdTW25MyrUhy+0CR5H0nyk6G1mK5BaReiNCm693T0
HxGnxmTAAlEId2aDWNeP+pWbZoTrXpQvS/lw8UdV9WKHkVXvM8SUaNGqIHtOp1pO
J6qlwRwR5yAm/ycwiQvZiAhNegBognk9PxfkTxdVhaIcAK3nPmvDTT8IRLL2K8BZ
SHL+/I0U8LEUYarkSKzJW0WE1dMMg/KjKo2JeUnhPqnUdu8w6zOFerq4XL3OI52C
4cMf+P5ouE4lyFIHvKyIEq4LF4PjmW4E8MTuhSTtQrbsVMpYql4ndYncDyStmF+Z
SjfptVNMCzsQ6TdI4QveOCCN1ByegTxafBtDxSy1tjPRknoD9OItdMzPXv1j9BEn
jrblZ+IxvEJ/YswI1KZOn/AYEdlhtLGYulMZVBhyZ+NmBfSBIE23f4QZ/CrjqugD
QTqenT/8IocXyBZvTjOadhHQ7Lqwwck2gy7PVE+YEZO6ZPslU2icm0QfSUFToFOo
bLps0/mNZOQNSfny2kAGkYMLxwAvAXE6hZD4lcEMj8JZ/i3Rtn86ipvPzUuj1uH9
0tXemF4f8CchDJNuXOX2ar1wAovudUmqLVk63K0b9oFjLP2ps4amDSV4U57Jyizl
VOy7op7P+8RDpgw84/2jb0rgejAu8VYt6PVI0p/0P4rjuAic7eBAbGEJDTFb5FTt
EeqOjllkz+GHZRP9A8ay6cZdPQeVGbjOPjFoRu835akLjAEtRTqQqJVWPDNEKcPg
hiMXtXPJbfYGlcumEayMk5WpsUxBg3+mqXgJL+TXJ2V2kV8L8TGUGYYwon+r9Pah
bt1Bdza/QQkAWHCzpG3Umws6fK+wbSW1sYRNVa2Q/1OjKipTiExWC7dV2eZF/bcV
Wbm/JeTFmYTzhK11JKEUmmNugDVOQoJumI0ro60eKne/wl2F+QlXbS4oCwiyDni+
/XUjL2VTqoI+m66750wVNcEuEbMxfaI1uRUeOKt5yWKlZ1l3yTA5Ze67D2WttauK
R0REWEGMoGIIJfnfhfM2p0+y1nRT1iq6G1ycgOMwoiwgzVgEKrrZ9T4fQ4/CG5AB
GYDvk8OfgmkV35hFazptGArRO3BeJ5limeuUsDxjmexFNIsrwrvMeg1M4Daxn+/b
0knYbyw5KzxBOVWJmkC9rUW6aR3/sxY22W1JPkP0zkO+zeqgC5B69GY2tdjK3eGU
IvLs97HrnTUdGfBFzfTaHI6uXrFme1M8j3GBY3YLPil0mf0a0VHPyL34IqQEm5nu
og3RndgWS8uT1IPAUVwlbq3+7LJpWQNkuYAsidKDKAlZkul3PsZQGUNGG3CoTJeV
8BhvKBMhn++Q0y3imyrE7hxwRAh6ysySToQb8oo+A5BJneZJJoG5DsvaLE67kYuw
NUSEgDHesDAl1/EBzVluIZvhVtFg/lRCwtQGMM2tcSsQGog5m1mWXomSChgWZS+H
91i1J3A9yTcbnuOfp+C1bfNQ8YMX3zG5dPqaPEV9RnrE61lZQjyH54LLTjQe8B+x
qzFTLe/1EOVNMoAnB1j5JddRO49R83QOTHGyGmuuxhduoInVbtYDGdqZ7su66KIb
woRTtlSbX7OKVCjiKLerigqHFxf69/WpDzNp+6TDOw1z8WeqjzdflA+6yiXm28y0
xNMpd+TmPHacE7ZX+80kfeJIjK/xd6vyqCS0lKa+fbfDPFUj08Ftv7KE15mBSx7u
Yaq3caL3SxWNIleEowxP3b9ad6j6Z/Ivvd6sYOxIRt0L+RFFaLI8d4ljGEvQNlKu
Kn4bc7/1P/6M/SOOuoTK/MitjEjVt3qrZweJMkfOe9BakA+G1i3vdCu1auiRcwoq
XanHxcpfBX2dSqPcD0A0TPq8/lSeE0RMwx+krd61qDgTzgMhRoM6UWRNyJXdz6Ek
sAHDruXENAKDTm5E6CXd3B1H5jCP6iJT17iJV3Ez+erQ3wjYxq7K5XabdiSH9e4j
sheF0z/A4BqDXGopeneMi9fUQGuKn+UyAHmE70YR7q0BeOfRY+pBPfXY/G7KP7+t
fdL5BQD6sxJM0IFL1GUZG6zDYA/VwOVyh1GjBdA3wBNBv3kXG9zIH9qpGVqTBPVv
xs8QS1osaHQqZK6pAUFlA8ZzvsaRhKCX3maPa1TIuL3ymNG5mUcEUoEjUDEYHnKR
PExkOwjYyP38LsQQ25TxhRG4ThggBX+RoKlCoGNXqVj5NTMiZXeRdWPDChfOLj2A
rmKdD0frJzm7HeaJ5It2Qk3GldiW7hErMOyAzVpTDULMg6aWSW0lZgAbDufxlu9l
++OmoxYTNgK+Ov9Ksfg/+tBvDufiEe4eDh4dj7Trv8EyejMdfHn68jz6BcIwTWhd
iTob7GkmH1WaQRnvOt+qw067fqQx9ovG39MYdN8lzQz0BykvQBLd0xmmUb3U0v++
vGXPVhWeoG7fPDns/crEulqfADU3UTzr9B3sXZhQC1+37MMYQ8PtBzzWOvIgtFmJ
vnMuyLeOjTaHqc3rESr0CpURFd9pI2ov6jxqwKfFIsKbyOkrCYr4p46DfGFuFjWE
69iqW/ZRNUiWoFJJ6ZRPsb0N2AcXW0WTzdWBDMx398DVpzBb4cO4tF/RZYGQWJWL
2NI1bvsqIDpkH/nLiDBOLmgrx2/zg7Up9Y1Xu/Etrvv/T2ezFOY2DMqo0qZ/fuGl
e64GxWhCUdlXoAkKyKtWNtOhO3dCQqjDgkVSObc+4ieWK4b1BCrGQ85V2WN96/ko
/ONCXN926ZGoDo3js4w1gizZywDFNDL2a61uzMkafH9dCAnHC0vj3VqGYcvTz6WB
xo8Rjw9th977h/2bu/qB/qS/0uijMr3gpjeqX3xYo9Z9hSTllnuJEtUEDAR8B7Yb
2Egsw6BfrJ75J4KthystdV2yEU5rDki8rggKaYciS9lALKfCqkIQBChYVRniIB0F
CEBNpEflX7iteqCGky74bnhyMKLlCNCP/uliktHeUmpA6VBFaI7Rc4Uj2PXL4O/Q
yov8e3Afz8aCEkYeBT4/G570aKU8Dfbqv69Xswt0cwK6XflIwmDJgvCvdYwNsFDY
rStAKQtN1aM6/ZqqzvZMsp3EADQlSCoG4A1rPX/s1LS7S6SbzFgrKe7yKHK0OE+s
/0xKEUpaNLJ61vGR4q87E6KerotBhKUIbaamDAy8icXpd3hy7NQdYnxPQHxOPo9c
+Dpmhd8opxi972YgN+U/oU5SoMMmpLgJ3YzSxGGIfLpYr4qTftJI8opyMvGRThzk
CSUgB55Pq6jO2BAp7KzpEwzV7gD9qdVi9bNKGgqTOT020C9H0IBiR/kBwGr+1sXU
hNCMkQmh+MjGPG7FuoLtQsSiGwqm/TcMD51r9Jc96eE75DDFXiIQsoxShXfM56Zk
k6/O9It8vGKUQ9iBW6mEWG76R06xzonlh8iqe+0JPyzD4aGOXZCaIOV86D8BIXnh
1cJaHALTITPiQZjpWKTQvnYxegAq2MzGnb5pPp+TJfPUIF8Gcn9r5um5J1eltYSB
JYbB5WgTprY7vTJyXYLjmD//eiZuSpWYTc9u79fD8QDfigUkJ310nv0EVpYJc44j
Ii9S6JNU+9DV5Sv5l2qJyI71vGeVGG2uvpFOR5IoOgSIpP6a68U2kb9W8yK1cTo/
nbpUNKkuMdGTo+oYxYpwr7SEU6dhR/tyqbGaFrNw18sEFrPQQNJBNptnBbU4gM1/
7RDyzbHdw1Lu6M3aBxk2oFO/svOMisMc9Yuth5Qxsum3zkFsLmHTE6LzQDWnfyVZ
XJuuKwtmeyqUTdSs0jMY1EdZZmC2giGU+8TU0VW8J7tk0a98Sxkdea5G8SdutXCv
tjSZRhPg6WfTtietmU+78MGokZb0NX/mEm72vuRtC7kpkbv8D10iopkm2TkxfB60
qUIQH53y0wt2ll7MIotYXCjSPQTPT3wQHw9RRYhuXYJKjgD7f5eT3dzVBA3fnqxj
X5kg1z79+3GhkM0oKTgH3ZzaDcER49DQab08k4lT12a3HwKn8N6dk7ptLlowTrq5
bXL3ScX7QEFNhOGnvRqenrPQP37Q/BH59mKxsKbMRv502W8GN1u4yfyotQlGOCIn
/cOd1o7ES/SnMslJ+A2LLSExquPFTQFbme04gm35RE6fWOKXnEtA0WvfzPfXLJs1
GFN8hmZVQVnz3bR/MQuOBeum+c0zpz1vD5+rdtTWw1tsJ3s90Re9WW9EI4Sh9Nc7
lV998qy6h7nRjU8oxv7J6IAp7JA5Gwwq9JptMkhhnv34ns2tuJFzX/7TlcMmmeaK
GD0ze/zocSMzvNfM90TfAg/ci18lvN4rTAcKW6R+inYH4fZhZhUOa9IiMHT1qKYw
T05QnpkBVOdHZXC5n3/5xzAi8qGDAMn+netOUp2QHXbXgsrjWrC9uV0gNrBl5lKJ
P5nAe1ZZ6BRXKz5HBaHzBXvoz7tMCf6kf4YAWPZ+Cc8v5h7/mPRxyy8MYk17l4Ea
6z95+rAZb+bjkJRLwkvO3aeG8IV4RLk4F7fZ8fTe4VsyVuOENMwvhHprl6UVqWjX
hH91WC2j86SFxCX+KDytOe+VvPZWdFdpI9dOpU056wTSWvtwfWVghdTqle0SsUso
cw8FPb+2BpSKEwUN9QBSZQ82bPqj+U5UTyBVUJ9fIsgJ1Y+VFqoQBesDZP7kc/bb
yBtSbxT+4nKtWJErheYKCEukDXbpSDHa52naNt4sSyhr/eB19XrJf1FVToB3Fkg8
zhvF+UJwckeBc339jQwtwsf8mwWf9WgZZWrDbziTSvwnUcJAsVdbOgNxMswDlWP5
osMxIarE1hiIbhYvtGkSg/sG1ofsO3zRstdbow8QZdC3dDCbHsuuEuBG18J/+WoN
5wpheqc7IjpxUCnCYXqcxLRNOP4xKRhFUaLZiDIHdRkPYS6qUL1TAZtlDaNg2y1c
UmTPGsaFCDTqTh+XmjmsnWOoWRtm+xoBHJS+JZTXZ3lko0duu9A5fYtGtWRmwMTL
RQA0AwhAEkPc6oOjeOcjjOQd64PIeF4kiK3yN9t2FtJqLiijADOG9mVPbcdnDZzr
b0oNqL0mkHdn46X3NuMLdsnKSNH8fwVOUbWhWMZjHBE2/63FdUY7NjLERmgi8cd1
nHdjwoh/NIBWGSNru/5/2/J1kEvJzICxDaWdYzGMUi6BCor4/0z7Dx9+0xpQklb1
SbmJ72ANTd8/W1+pVhjaMbOfMytSc9SbpDlb8hTu4SEbmjwaaYfbB3JMaoWKVlN1
Y+vY+TBy+CBXkpV7uackVUtkc7TAh1PPrmUzPe5SSOsQdZhYtRIvS58KBi8nB67H
Yp8nUUEGDG/LCfUPU17T2wnATHfU0jEjElhCbk0o80N7C3w0ZG11Jay75qpv+NVK
clBfPMYbjuy/gjqZDQWxOJ62BSn1RF0uApDdPd+LyezjEjcwyvX96j43YWBqW+CS
3RayD2h2CbkoJwlepWkKTw+2Ue38VajLQ5ycUoiMEIgIdvWm4ACIyjGAb7dhMd4v
4K1ihIMoFAb+/+vakQ7n5qQgFQxv/ZFRBiV8R1EeG5JQf0cLVwmMrNERFBapybqG
pntp26j28+GUAYvawyns1A3XhYxdvlFiNWmgJ2DXZlqArqpAx+n92YCs+lsIzpV+
gmYlN89Hm8EFQX4p7xYN/MKK5zolS66lAh24ld2LdKsup/pM2NC6s70tBDSnyxcl
kyEI87V1IJkzx7wIGfU1aoGO8rjv+htagi3NvfXrtPqskOg/DBBy9GrOCCqeAh3D
NPquZKaFjFrL/rApMmcJ2V9QShqIjSduCNcG175hrSIsf7j34Px5NnldDxZvktbg
68CW7BrwFqr+bHrMaaLtwgu7Ju0bLZ9K4AWvpo8jbaf4hraXmqe0qmK3q0TaU9pK
k7YzAnVw1eQLxOar3Z/Z46Ga0E1loIzEahvjpnDd4vDMomOKr7QR1jqcrwtFVujU
X05dLX29SVF6ZQ+yOLOyN0QT3PhaWiMhm2XB1604uObc7k22mHr9aCbKpmI50x1o
FZj1pv/pY3uSeZNQJL0Z4kRvX7fgg3w7A3B+4d9D7Mxoewx5I3qHHywnH8Owpc9D
gc0okyOn8U5ctV0zslkt3b+TWMMt1+1chrVMRge29UXdbm5rfIw79j7hxr1X8mB6
k8kBg8hFVxjh+lFHpYoVJvLMUMpc9IavPQRt0FtOjucf2NN9DpsZGyv8qZDSRL/V
a03XprDjZbKpTj1iEByCzq9lVlCRX2fZhENP99ogFwNr8sw/mW9q/12pTjrACb0y
ke7JNv5gtllFlotIZ+z+z4pLGHz1KCdJuv9ftIWzwBEh49BAxnpNSVqP52oEHHcq
ijCZBDTbPsja7McScSOPIF68Z3jfvML/RUxlqjOdUT5AsLDXGZV7ykh6RD+0vDwl
ocI+dbzqCmb3Na+VNg5n1Opdm2IGUrbkfluSzI/wfhgCdUZKF8KH3VY1W1P5c/Mx
IFSktTruM+Dr6+OoHpJdMEV1O1h0mru+I5HoI1iVkNDhtOdV7tCW6c3PnFbEE8C7
EQdd+HYfl6HALBWyQUeb9zHrXaDlxO9b7rJaqWRBVqBq+1QCQFt+xWwIOTX3mDiA
xBfVreJjWSpPNtNrpdcuVcESslgFoBWqrKMdypxhAUzYPCei4YRJL5t7TYLhOTl1
ihjMvIfF/1Sy8hwpbEtqWX9YQkw98kx7GLsG5XYdDDrx1oCYFopH9KFG/8Su29cY
tq8yEEE91hOSL/NPow7cyuKB0mgZncmLB/nVVyeAmtRvVCMUkeixF1ThOFOtRV4b
kHdgMJt5ZHjg5d8aA+XEMZPfxrafsVd03rbrYaJLoaVnvPUVj1BjOg93P2/OogIg
Bk5VvsiqiwiRFDsNB2nGMOzLv8wrpFEHO4zit/c6abaLVzV7q2wu7W+K5S7AIPIM
DrJLSpY9ziQ914Lu0Hu3W/mDIjH05UO19JBXDfKBE3fER43o9bLs5HjLcQB7Gb6Q
7Vndn0Ynxfvl4bslmiJLo7oljjza8JAVqLRHHnq3Wa7f8ecdWodcQANnmuyk+NJA
SunxHisFuIz9GAN4yWM58GghlFwrXlG/bhDPQGoZhMmEHQprwS8lrBy3PfOEl0g/
mPrr4M+CXrZkvZZNjOe+5V8BYRoR3Nf0v9ZMCNC/u0wBxzhyVUzjoOsCwMsh4HJz
iONrOqxZKCfWX0Ierx5jaI3dwZibsPDBhmXTSZqz4e19G+bmLH5CNnkgzc9D182N
AGMR522geb5uI1UISYR83vMYxf7ZGTuVrvvj/S+U15Bn4UM1rm63qdxGYsvyvnby
EJpAxlPol4WRKEKVMF6ATXYHzVs0n6lHgKw4Vo31cfkLoyQJitCd/NDIRUNU7LqC
jB/e5dBh9P1+cgeAVaUpXBTFxTS0WU+9aqEOc3hOp9bD7sBMEhuijc3BTb0k9GO2
b18EVRyd5ndt2xDpmG04Wohe84ye/a1KD+xpSK6WT6EqgycpnvyfP4VjZkGMBLOj
k5k2Xa9UPUtxXiSt3LHXBdtjFFjwCm7brNYHFnjsp1PM8aRElgYAbvIUD6osn7mc
OpYCC2xUDNPWFeho6M41r/JQC70RBjTdth/+DVnWrQz2kk/Oo1g0vJuk4mGxfdgz
waF9oVKWa6StGQ9zUZBK4ExtaA0V/JWM430sk+zY0NrwjfcMdehrv6nvEcc/9HPs
viTdFN16YX27VrSDPv75y3sjpQAkeHLP5l4g0X1riA7DjsmT6AdiCmSKV/GsqWpU
6mzvS8Tw/jsida9eJkRT/w3c05U/GXSr63aDX0C8morki6Y9EpIcA7KYE9BMoq7t
X8S2IM5/l2kkXrsnu5UF/YcONV8vmHIw2RIikI0AihdwPw54dfGD71t0Nu3aY9sr
NblR/d0fvbMpd3biFagAzcV3NiPyirpP2uUV1jYRne+cxrYTznzdep1mShuXzGf+
HPQNCP8Y7wQ3q+0MSGH9+kYZcy1NqJ+IdV3DX+7kL3r+CWSQCBjeF85shhGc01oz
NMXGWP19T9jId2u+gYvoHPf/lHS9jdsCFkcwgtE3dlpkOm0aHnByB8X8AwOAaiwP
BSvsCS/ZnU0TtRKTdHjUxXZflReTfvkeUmcziIo4G0z5Q2VRHmvZtAJcuCPXHCFn
X/arH4C2zJNT8AMWEs2C1PCp3GN8vFEmr6kBt0x0IG9uGcfn21jWLU6ECzrdSTi4
kKrT8xcPqNCWUEUI5o+n+Zh2cALL+b5VJD6smu/cqQkPM0+Q2gky37Im0WlSuQK4
CkqfKmTJwmTUXvckq5zxtzHCi3DOqFLk0y2TB3mLUAA24ZFvhAWZbIAzrZe8Cyb7
wbKw/ODEWKuZj6ftxGB4i2JA2PEYdabtI1c/mvEr18i9+6EheShoYq8ag7HX4ClU
cpWtF5I2MuieKCkvPjLdDEbteML1oOE7auxgNYmwz9ehQcgwEqbUQQwZMPauOjl/
GPnou6opSe4tqnTXUbm2KXFeXJBHIkpRCGQbda6A0ly+KYD/SCaSsi+aKiVYCsgD
OYhoyOwuGbMgb0aAIrHlNXt0422phtHWiCq1waAv+dgyqCybKHkQESWaOgC8FZQh
4LQoWYVspY5Q02r5sZu9/6q1aFoCO1ktjXQNUQsftwbD7pOasDci3nxbDT43nRv+
s/WvcwSzmSz6X5VowKexzXRHx6XIDcFkevpk1b95PbrJpHxahAqFW6VZWK/vwVcx
yqDFUvC5y3vi6dhANqtC7n3h3AVHqdJ+9PZXjbX8GAPh1xbh5MbU86oOhs+j4RuT
qYLUE5UVr4k16UKUq2qNCZmpZOO+Kkrc5u5gg6Sb5JH9i8I3VT3EdJ5KtkeBGNxg
Rb5WRMEngpl0EWeNt2fGqFucC2JtQAAvcUcy71fADEOS7jTQCF7WCbvE7zfPt/qY
ck2vXM7zgOKBpL0sJ5egEgDej0jxkuBTGTwzUz2GNVYXedNSeunPC3Uy+1MRzBFJ
rZUOQAyaVl0ZEsx3bu9cedp1px5VUwN6Ez35TzlkMxQLo2/VyBw6WMno6rP4OQZr
d3rgc7mSh9sPy/ulC1sWwW6Y3rf4kF3qhsqn5JdesAIGgfxotuCbbqIaY6xS3jZ5
jcUB/hUEFbDMj1ylhjnQtafPB+ohRZepVJncsHGeeu9h9k9jYk6aD/1THQ3epjeQ
6/roQDJxeX5OfPjBagKJi4kGNOIrp1NIuctTcj6DLmPtpgAzT3ZoMGTq10r3vm5N
a9z9DoQbRHZo1ImYlzES5BMXuLuc892Nkrg6Oyt6Rd5T/aGApAl8381iPE1Wqz9O
38TuUU9S+QPn5CbymWV2H1MC0rEdCL5GaGSni3VHUJOfxCts0njYxpglSafYTrXA
GBbyfq4xAmxIyoZGrkzca9cMnAE8HP+MHQALUXiVdL4lGTG4TUHCHSt11ExUdjbT
TK1mKKar9KR3t3EWy7Wthzm98h1TUUPgjeoEpukyf0VWb6Oa7NoXWRmQi2IRTgXc
2WD4DDq/vo1ZCrdbRb8ApkQhWzyXjmWuJSxNf7kaBiL9HAy04H1Lwr/BH76bBGQo
CvFgVyjCDbOKqJLEpEVVWj3h4LhldYCnZHkqd8wiJjMUwL9c2LH0+47YmVAweXpD
TWfuewHHLtldBpthCggZRWYcPi0TPxyLvh40LcVMUOmTyEJZCp6iUwVZso1zUEIf
Avv0I4vDF6iYfdohoRcynXG+FGG9+gxJC18bJb218hJBTSX7l86C4HjO2lr7DFFz
ViJaly9SaLD2aHTCSJ2Z8QXOovcL90/9P6y1gSjlGNEAZfqoy1eqjKwWHUizMA8U
a5yP8FWC1NB35At6T0ah1wfKZ83am8ll89vHQD0vKtrDLxO7Uek+DJMTz08AsBQf
DYk5+a8OftRlvRYnUzIGfmhDY9LVt6o2ZNg5aLGbUrLSG6S7vfTZ+ZInQiV2rsGy
x2qB/TfkWv73ibW2jfhIA4H6/QEj+5YRzaddRfZQSoKeuK9jn9se2SgePv5uJF9E
be0NKRfAUQ5vnzS9porhSGML6C3VbDxRB2IXzIVKk/VbNFQEQTdRRwkqrqCCCpPR
y3XGQzarh8354cqbHvkE+V6fHmB4nCgMD6+6XhRVQ/M54S74jReO8M1Pe8ZNXGBJ
/AOlX1oezXUNDrmlyJKTFIss4MdeZ9RLzQRa8rusm1iLBd4sOqriTRWAXxOzj1Q+
pYfTtwW7WAhv9y7Y144tuKAKNjKT+6IRLS03Hf+hM2oetY2LECPGiZ4tQurFsR+a
jmASnO9++LVo+XvNXQR4Rxd3IMJEW7B5oPRXXEQx0CAvEzb7FeQcJNsYqE9WYt2O
PW08E2o9uh6yv4Wr00m73ACa9Ns7JyNC4Xatk1ovVwzSJ15qc5fklen6S9PwvDHJ
Iqin8PddDjT935zYPLV/P/oKJVjsdJ3jwNU07ILqVAAdqiSvklX5FDJ7iFbsv8eh
WfppLtS/mk9mjguhKVffWuoDG9gvuiGNki3Pz4msWHx2hzyL2ufu7w6hiEjsa2N3
Mj3lQ71Qx6a1HsaoXUdaunXUUoRK0yVa1VnDFQFvBifHrnHrLz4uOzATGJJ+B0nM
nRJy2YkKBX5rPYAAlMQmz/ah9Uj6z8/DVr+DaHBSP1jOkshtcMczLdlmxlkN2Zlz
9HhEpTV2o/5C/XSkrdk3s+bvgMT0YY81XgDpbtw/AgJUpq+H1XA+y65W/WZ5UCD9
ItY0Yq6EtiDhc02NWgbH5mBFe1jwyIzLVSPZOmSAWexlMjup7XbKfGf3h4tR2P/q
vc3I8AUGFO8o2uPImZhsrNzk/yYKSnSzhLxd6BT4aHxiS71KcCwW3mxJsQSkusll
0nSloXWSROE0Uazh7hnpm9ZK5UCblIwOsQXaeBn8FZdZ1EBkY4R4bLw3Q0NVs2sI
N7r7gSzGYmCI+ObQkGdBjxKqrp6BbHl8goA7eOPI3lsMV+Ng6rdFaYHEUL/Z2As+
0ZYy209EcbOw8SQQfA3avPFioVg7iHj6lYCKOnyc7qsc8cRrt+aOl2III73uV+QX
pWeI0SPk+8ndvdjiLyUMl8e1rei8BtHlhYrQ5nOvZE9c/1k6FKANrWC4qQPEj6DB
vuQnucFKFKfZq1ndUHOUOF81ahAuyNjYroPylYETy4Pl+SE0Sq7JyPWBpki09DCP
06Rh081EjJYFsTwQ+3t/qN3SwgvifDpBgbp+FMIzmXBpCEitZkub6HtVupFSvsIU
fzeQ/Rz+8TXCjZT9ENDPabb94VJI9gVRz9gTrwFn09AOzlJx52/ljdzxz8uiGR+f
gEWUFeG1cwpy4PkMtnKCfFMiH9mo8BI2HnSwkL8S78uy07y/P8ly6+WjxCqmA1IQ
otcqGb25ksbnGCls7y0PwxC2G37w1CnfiFXxF6SyG+QyIrNL4nhuGaEj6jGOW1jk
Rl3Ps2X2md4L+HFr38t22EtlHxseCFESDE0hD0wHr70MyHNPh3EGOlj+F9Gku1zZ
OWPuDUePnkT/Kbq17uBb2VTQHBPwTqnlizmsr2TkW1sIDqV/US9hjJLuZ+xQk9yZ
QGBXKspF6xFYhB9uLZf5dMRtOm7Wb0eLfFDeCQhsp/smikJmfvPCPLwNyQx3SMuW
uF1vOcddBdhh1Aa4sVvkhDvoo6a4hnLZ40x0q1tqSE6dbuTyystAbMcjoEYpJOWZ
D11ZnnwT0Bok948+d9xSr45WjETx6rMDfD/jf1qYAswBfTA758j3Sea1gRmGEY+A
74+YjMpE0+nVRYDodXv0eaepCIO1aJoyTTC40fKztzgTcJtu1XKgclRo6tChSAQ0
ydHI9fDI9yEdKZbUFIxmOD365bzW84uITROM3vwyqJ0zI+ob0mK3GMPj43bCS/MI
ud+997h0X7gpraKNzLPZV6lML30NcqH/inTu7Tepl9gLM7snQLG0PMvm2MHUv0nw
weutp14MGs7rUj65WocbEL93Ho8AqsBGzmY4yAk/HEOXgD4k9OFAsGZLWb0UPx9W
niR6LKb7fW39OfPpUDIS9K2S6VRD6MySewdWX6+FxFWVKZGAu5GYGSuP3Ims2bw6
oVbUd2F26HXWNRHbN03OqiZ/NM2d4mupIwHctmIQt6WuI9Izvdwkniq53aJSkMEV
67EbyRcHH31XnhhaISy+GgYfw/di+CD/DgqidjXdUyvV2P9c0EadxCOUPujVi1uJ
+U2rie+JvaIVVlPfZyxUsl2NLJ4OkKltjGlUhmglpAM/UqSA+H/mmD2XZ9iQ9ELC
HkDgj4xQrl+JquG/S5ggzLPP9+G/ClDfjgdzK3XCYbD3/ny1gowIBbSSniZvfNSV
ONnt9Tle0Fg/xAodvO99Pc+ek2DSxadGNqHHNob8xSTwmQ+puyOLWghYSuU6jW8H
6OBqsF51YY5Ke9EG35WdNXlrs4y41NI+rkd24TwJpmoD0aifyWp+ppTXP0p8D2dX
wbuf3fRYbCk4c5Bt0grDB4gplQLFn6DIZr5RUHV5ebb+/0liEqN2x8su49HtYDzs
mmRoaygu5ZZRc6V0N/ytmbvEBiW9PU+25LnNCd8A5SLJJJVImsXGiorJ2mTJ8jAv
QfXHFsVER791Bk9iMCvgKvqUkm2KymOwE3EiFkoCYNoSwgObHpxhfm9coMSlUBEE
fL/Krx2q3FnhseI8rZyYAB8Vkz7Mz8se9RCTeYNZLnP+vmoIXQitBBGO3nUNvWF9
cdpxuhgnpPdVoa1aIQ+pb3X/YzeYF1kl8wi2zyEHiT4zuIGTMeYygC3g8LvHiNnY
YdWN8B9r5HnvDNmZpIblknDxF9YNH/U0ql1iQZNkHhhYXFEavixiR7GzouMFCXAl
SldyadWOPAbDQSnRtMHu0CrmNga2vsXL5u5zdVRx0PX3/TecGrbVnjYYaieOL6uO
9N5MmPPVyOJpo+HuAs5Y65TOwIkkzGOyKQStCL/ci6Gw3eBbaSbyVYnHmrqZVhDm
ALpxdKgK2ReMx/6dfU4Yf7FuLLiMeuLbNqx4t4mDok+2K0+xEfnDhfP1mtNhX+Cn
zIK5BKP1NFTdtNp5voXDG73e0eKYhQr8S8Hdv5cduPaXzKwc0isynZKP9T5L5duL
y/78MfYQxCSAWfu9rUC34a6oXe42HVzalmniB2+PXRrjxmjX/ydteR5f7JcHsGZw
JSv7uCTWJ2Jy+ZDbUSTl1iiJjmsc4QlJrwx7aI23SwfNsgNJvb/CWlHtUQaskdsB
HVIneSImWqjBquDg1eNB1arPIT4822HYijpK0R4OCI/2GmDAxO0MR2R1oeTsI0yL
x5uy1t6VUavf9w3PQeXA2bbYda1U9PR6rZUNGGe2eBj28SfahV6nGZ2PYylXg4vM
ipmLcjru4o9tPCbMdOiOTli1l80lOa79cc6F12Pirbi37JEzed2h+cNbJWBobqNI
l5SHigNxFYox/UsZGEpvBiL33sp+7p0ukVRN7QhCmDI5MnhjsNuZLf15b/p0kskF
F829QwlXspVVogZamLcXg5aBT/gOd0g94bvAqdIRAQvvQWcg+O9hjyM6Pdj/PSjL
/KmCVAq7nLPIdkT4Dr4uE0IdjNGj0LiPqguFf2ZdfS/w5+8ucH82jgssseN8Th70
hTgmnTnMgz7KTP3qPsR5NQnhCMOGbIAGtih5NVzXrs2WxfWNhWz8KtmiOGImLTnN
+E6L+lhBqDYmh+7tcHtVeIJhS74072iVvwu5r3n4CyGNE5xVeDdBriYvUAqpKXVK
M4g6aoAZI1V82kDECBs20iq6jIdIwcrcpCbq6/+0UET2759e1d9jdofcD80A35VR
DTEkwS2Ms1SSplaRV65CT3P6p7Ktqeo1HEG289hDGIupkyCHqkAGoWUPMaYPCp53
HrxjDCZnceLgsYLicyeRclyHNl1yN+/NtCSjdlRHb578isxFV3xjRMI1IJ/WkAgd
Js4f9q8r1VUVaXuO+M54LS6IpqnrZwlOsIB1oTxWa2CJqOYOgoxiLS/BMxKNcLra
92/v0Dh7LIa3z5+dsdpEVtkKBRxrGGpC5hn9RpQgVXqS5+D71HhU2pbxDXlS7jLW
dQgak4kK3gU4H2t/K8dH3FbYKHiz3CHg2hgrytpqLpimuFTQZoxlBAatufpQVT3D
S5kLGxAq2rDaESGIWk83PRdDRfR/mRgULuqNaMlpxjYr7bgsJSXa6tXsLVIecr51
UFgZld7JNBTCMjoOr9gnQm7ClD8IvXba7ikiLlCkgNr06joU3HGN6im/Ykj69qh/
fyPWI8VJtpGwyA1Wm8j3OXBm9tL4qcYue81nKx7T0xFxN/FOZPTcMSOJEI4VB2RU
wn455W+yKj8up4u94txeTA6fVsjoSjxD9+ophVFhJtVS2tNbgr8yGr0OY9YjEv/0
F0taKHyp6j0Fg6+2bpvl5VyiuEg1fOdBxymKZnhf0DFCFy2huJhIckJKYxdjBJfF
gkAjAbot5Sjk4rsotyRaeTF5/+M+gtboBi7B/VJlrBGPFs5irYCsjq2rBck9qkO+
3Vbu5PkUnzS5bk7q+1v7c9cr7e5YywkikE3T/RCkUgU+esJFDSiqawKCKqvipln/
x2tNQtX30c9FKKWu5uw+9ZZorlSKSXmeD1nLPQp1hr5PpyhSX3dsFuTkJ1NgJy7B
Do6GAfKRMd/I1c1zO6nVksfT065AOo/0t0LJhpU1GpDVoYk1C+rbxJVWlAf4Ytyy
+RiPN7uBZ5tHNCFc/jUrMKCNv63F16U2oSDs8aq+1fOssGgIziXfEv4MCnlMkK+B
QklfHWNpjRIEc8B1yyb/dr4oGRKCW8fmaJ+vkeBRLUUbX8KTtiCujT8dV+uMrgjT
x2pv8SsF4bbuVqWACq9NSao0TOj6XVf132/yk6RRAGN7BG3C7qvH1xc98XhPngP5
qTbOVDiyT9lEzLSKhmbSD3yyt7MtAkPj61fVHg+SOHIpCSCGMEvhxIkNSuCvXWkU
tzlSS/wuRt1xp86Thyqvw/gzTHgXC9WKJwoPu/qFOqbzw1fcBjTfJND2opJ7wSdM
lyBS8FCV1+C0frpSlIwn5MbiioCLOu52egiMIhd8F/YfUs+jbc4a0lKVWIcX7jVg
yXNv3pwL79ePOWJ3u2qzgdpsWBRu6fqdSSwAbCfueKKzYgiKza2w+jucDOagyjo3
cN0sI4k/SYKOvgEZCNhNs2qqU2ol4S8pJFhkqmOeTxffvGI6eLU9o9aah2BkEkVA
z5MX71HJcq675PVu9hoEGwB1e6Oy0afXqLesEDl+DNzMOnO8YVJQbPdc++/iBeeN
nixCFhhZHTUuTQ8fyrG3Ibm+aLyhkZJCKGqcELIMLCTud3Zt4f7ZiIZeNkvBRqgF
5YhOd0Hef4VZCUU6i53r9F5QjWt3u5ZaoWOPf2GlzTFTXbwiWLWeJq27oQab1PjU
LJlfFMEdy48g9t6V8m+X60ECdLwyUL4iNIKteh0w9hy/I1E+U9HDn74EvpEQbFfN
mC4Oz6ErZzhptMJoJL9WLEHRshi1zbHgIvoA+yc2jhAfrpkh0/wwpgf2ktJicOSz
WGYwXfr7e/0I9XPw1/4eU9obNF4ayKqQ874EpvFJDvtqypSVt7CaNhSqmtNbF6z9
XPUF2CPRohwkNWc0wYxFNccPaS6tsIMTQowjMR2l+8SOADZcZX/qMHalLmsC7oIh
bZiqxZkijycWRgGDxuA3TF8uKcMThNa37tLK0gboaIbYjeAE996yGaVyDGCjXHac
aLyvRuZQVIls3C3TVMvJUFatpY4UWCOdDgjVHe1ps9PcNxb+aCUvRiXXJJhHzIMt
OQ/qVIKg6ysKfqt8klBVny5ytv3l7TxAMCnzVXajNiBgrvAGDCkOvQ3/eKhYly1y
S+G6JK8VjTogRq/Pt7S7UnZ2ZiYOKBVdTkK6RF8QLSu5KG4LuiWv+Z2aMl1Qp5I5
xN2sqL6cIRHEiz1iboyt/vZuM8GUq+CjdESMg0Rfn6W+dQML0UA9WyPRtB3rc3Rp
DI4blwhAT7C29IAg4hinYZ4njvfLre2NqSV49lMu6ij6pZqTVLmxVcHd4yE7PZWV
y4YEY3G6YPxN77WzLzzoLclCchp0yCtQIPHp8bk5F0SOXJRxcFB4H11B3ZDA06Cs
oEXboVJS7M+Kif8iaQjiVJmAzprOZwqgxzmvX0OdIC29HGhJgY5kMXgeI/au7KK2
qnlciagFNJiZjnU0Y/zlm7i9LrDhWeOLSDGggqqUw2mJqMAQle2jOH2FBJ7CPl3U
0+QBwUb9h6R66xaY35o18Q1ZLBlOSDGVmCzbfs6LrVf1WhrUbPJXtKH6pbZZvYOo
DeCrSoza41z8HKz+JpBCeyKQBDmLfW+bmz13iT+n8Gf3r4KdmsunwTPPYuvAD+Q2
vn/YKsUz+QYmEZ0tGRFds7ubHoblEUshjVi1u5N4L9nlGt2LfhFkrkCvbQZ2bhHv
Jw6UZlZ3xdecXvnv8d+dVwAk2N8GETBwcSOXEw0UetXF8XbDyqpK1Euwkt2eokA/
IfRE/XL0MDxJWGl5ZlZzcDAwX+FvITxEaGXthixHKe3yUayR1yuNOxyifbW+o+pk
AVMXJ8kM7zjCk+TXpfXnsBDp/YBZs2JnDeywClGO2lp4BLlLt2lLQ4WNy9zIxIWb
it6/wJZjShuJrxu3/0dVXTdw7AAMbZSb3+TJ/t7LKouAdjjDy7cWCLRWDSzog5od
l9o0PW9E7kGczzvjlTx50+8hF8zop4YxoPfq3fYAMPn3Vz16Szj9+CIUxlU/yRQC
Tlr9uJWI2n9kg5qm/rvzsb9jsaw1LOXkcNDsXMheyHi4HvGDC/X/ltKBMkF4moYO
vKdDX9CtJUYmriV0ktznWawlejRPv5d/ohPlW9qkfTmpGFX7Exhwv1HZpQLZ9w0X
5WXUZhvifb41JtZW21PbkozB2fbNKrA2VpW0utNZ20OfhphH+eUBEnAr10SCn6wA
k6puXF5fBgsHNK7kBRfMsZQJ+8T9+UQhoxDXX9rX7fQWEihSZrGV4GQ+Kk4WCFhD
B64v1REVVS3dMQx4Zmo7QXXstQCSxLCxOZM6qDTF1jcQ0Ek/MF/OUFvTSiLgRGUi
m9rtNujhKJXlKA9Srw6HixhDXrhuPRE1W/1tXox+z8Fe1QDfwS0oxS7ZqKa45Map
ghLB4WE2gkEk6i9QDYzUbMgBF/t6nDJ2p5O2VOTt6vfx62c+EJUJgcD5dstwTN1r
dFFpC2J7KeeULa95gfOAAueAyfdPDUJ1E9TWdzDXS3uHrWfpUQSSoF2+CrWj480B
O0fFTZa51+kdAS1oCyJF0TDkwi2I1zUx5qmNmx9PK60101FebUIc0U1rGYFQPqD0
6mxLJnt8NYBM1ZMSGw6cvAnwWCoH1hIa6ybP6ErSf8EHLFobQ2QYcJte/jA0OXJl
HvMVYgRL3y074M7VV+d399ZZ+wS0pyzY1yZQrG5zNx4Qb7qcywZ9pEQ9vF1r4Q7v
5Y9Gz4mI8e9SfdlaA6jr3jkJCyKq5r//uN33i82UYnhFcQ/WHlkCGXx+U9FYGRPU
I7HLV9tzj8u+QV3+azYmlDjTY6nCvcKCP6VJidE+n26ZgKFEx7MnUnEEUjJR8XoE
LlCZXKNAoXW0aaOeC7WJqIudbY6Bed+9PbfXwsmv0s/t4t2qDVI07v2ZfQsCE+RG
jUY/Q/1eH9HDr7TDbmQxZeZjwTWkuF6KU2F50H9ZMzYoVp85LGIRvod8szSsfMYv
9KrL+MOVxnBxPhBI/xGG61RFoMMyPdWP580+gI6QWub+Zbuu2C2JVdfXCsHJQYTq
OhulDu1wLbtqh2pFBICANoEsGYPZuEk9rBFrrmCqYD+832XPVvc2CNNLnkfa6HqD
Jin8o1z6Bh7xzU1bFCMxjrJkTMs1eaWFUE+5yLwyO2MjZo+TGjC0AqfWGMyt0jBp
B3OF9U65GP9E5x8xnoYCEVAdR3daVHHpRFugT0RaSlUQUmykSDG4WzK39rlm+KcD
3AqFtv5UmnWpGg9nN1iZir+AKmJhsuf502VYok/Ch9/ef08SDfQQs2BZB0CR+cSh
YuxvJw/8bJdilebKTl2Xw/1Rv7vCIkAZFA5RZTlYNiiAqUIyb1sKQv2iRF6oo+da
uzc8+QGC6wtDqpcOqwGpdC0viWnVDWvZYySx06XGX9W38PLotTNmuhMv/mw3hVaa
FJqLdcL3z4BSpWGM/+TU7kf/kmS7uP25y2VtOC2JECJUcBl/OtlkEJBlF7oVyNbt
q10rfGW3dtm2FhqVzH7SpT760178ci6bLwMZU7O3+cgLgSp9Sqds1Vw5AeWqSVyH
qj7+np8uWPxz7WqROpx8t63Sa/LVcXLYOA1BoiEeCrh5PCTo1hE2f3yagP4DMfeD
5kFA7aJQMKBCGDbNLNm1LDBLnE9odLiTyDjmoEUXf6cGzY8OBjl8XAPpZ1jT0Z+o
sf6eArRZKMKwQP5tJOxCopGfoStJ+94baxSmvaBCrtie69YfmdMg9/5Or+KuOAF/
Hu/UoZ24empRRa0H9z+ponFDBcRY3PGn0T7tXcWvOFbgQvjnvYbDv4mb7gM6aNk0
mNX7cR0vCA4OE6O9Dn8Lso7nEFunTLRrabfZg0TvQklv4Fp53BWIUsgAv/l5s2D7
NU8yda7ALRJyRmlVT2FnEkLqySR6xndi1ageZj2KJ9Yk/TZcSzU4j5YmU5BqhDxr
BOMd1Inqlz8tDsGuJigw3heHYfV1IrbZokotmYsYMt7yNeKK+fGLtypJZ1cAwfVw
4Qpz00pn+tPhsFv4k3/0aA0LHfqjyVvcgGfpSUddh+f2kAniCrqRHqek78nZujNK
SeIz3bVom5wJm02ybfLUejne1BSY/3QlnCIkcdmeETcRs/PChCMjlBM3eqK/IFMN
c0FBTRyzXQgYpcCDfrKIyW5O5MobuFryIT22jMmGIOPl+9nJxlOzfmxGK5Tc1dVU
4j+QcU2IWkmXPotSZANo6U0BWNagfO9cvEZXuLFW/5WWkv6fc/cuHpWdlh7qj2CF
0A5ODeQ+ysHX7987CTlFxP5Hqc7FxLCwVoLxVLibh/l2mIqf1INdZm7bZgUhfs+u
r+SzgK7vKaOtJ3TNzpHbV0SmyTVcFTGsv6dVeRkezIWdUBbGMfIetygRm3BcCBS5
R75RjqZbMNmvo+c34zb907enZ474/XdopW9X2X1n59m9tELPgNVz5N7bCjDH5NA6
5G1cF//P+sgQnYPyl+JM1w8uqdNl/OYHDHizaYdEyNDjRvTYpgMLtfLYKuoW6SGD
m4wECGspSORSUeLolCmAcD9BCNr9J5RgX8RgsvoZhJl/VEoUdZNEEL+IkxLepCNX
upJ1vxRQf3iIgjaR9jZigAYiS9+jYCRJDn5478No2/Z4/LHW7J59GUeMtvnFzeIj
UwvPdqs+/dACxZ5lrWgrJYwS3sUd/qSepubmGrNhgckkxi5jMtzw8r2sOQ1YRoZg
gsbISsbAIPhrEqede234A5R5BcKEaKKP8S0aGeYhKPStWVnx9TfqeInyXlA7FpJD
2SATUs6OTIe9HUgZXT0UtuFBgdqvrZutTzhkIACjiit0NZtfA0ofqVSVaS0VY9ba
r69wcghImqJVkOVvFUY/PpDDl0JelbG47VsPLhu/3VSclHlWcG4gAwqwZKAM6gCQ
9XWnxmqZDk8wWXtmDaWzOlEEPSfqZXX4K2eMlPop/puDEcWK0XOgDUD4RSQeBBno
R569huUzK8Ui7qCLXNvMv+4dZG/pdlhzVExy4aaixxUy8vPuQcG9suGtpJMHmUrL
D3WeenBw0J2PVbdWyT4Xm68Fnez2ikLZKeeQWqHFpa9RAoIGKPS47anv2dANDGYs
2lrwPqWyVWVw4Y8RDfYMsDF6YsZCqYnR+sJGH/vUR1iHR51wNftWB9PJWhKKqafV
BN5GhBIzgxeyZTEVMMA1sZKHKOIwUGmioleRpUJG60XURCnWrB/MZAvY5oJn9wza
QqiU4fjzJLqU0hW4Qd19imNzC1WqmoF7cyvNu5idIQiB3vn7aRMVy0j69SoZbbWR
fzu1jmxN6AcZLXYPtM7lwklKDgqAhU4yUGuYjKupGjGFvg5st1VYIXuzdt/UBp8n
USeX7PDDxWojTaC8FfNL0PCwvs1UwitVYfeIxeMqagRpjdqJ+39Y95Ir/Q1MSXiL
HRU3aVYS4gjdGx0AKPJ0cDM1gX2QizBOvliXNdp7CLLCc4xBKKs7EWP46+TDUZyT
n33ig4fN62lpUb84PmvtrmqLS0p1+yR3bWXIKk8/Ac/xgZ+/wNAkdCYwG+A7jft4
t/Um9IiU2INg02AxqfuZqA9CY2v0+bjtmA5PI3R+stjJSwacL0iVuUadTkfQDvO0
E4bjEDjfXkmKycb2Qs+ePNssdt7dXvD0dLqlKDZLYlWt8punUxNccTaNAlwyf1bF
4qjzdtIr28J8vyw2NXMVY2oe9eeb4++a7LrcgNnN5MezhR0aFF38bPZvpSsur9Xo
NgWEHlGxfOC06rl2jOjekN7pVKqWB27fgxjI4PW1gqUxxMEMkRpnqqq0Kps7OTi5
WdHgASs/rDy4XuW5tvPa5bkLF+e2umYxj+B772zDS270idXKWI65gjhU7EB/wFSw
7IZvRVlQisjcDU057dfsiXTsuI8Q83UOU7PUxulVQvwQAnd7eM11iXGpA+s8e2f9
dk7Sn7aCXgG5gd34QN9tdqXmMdt3NUa4eaqTsRtsVfO5sQhPX2JBVikZpC9+du/S
CkChvrJqyp5vhxh1IWlDuHdaeXqiUCwaid1KMtK2s59cQ/zd3MlsDZF3ZequzjDY
sz5I7qzxxub4mXgQ7c+0+BbZP/ZG1aXNB4OhIbGMnfa+wEGIRnGwmJjZhXBzKkpp
f7hgVNA3r9AJqSanwenwkTg2Ux/8eGWFlWoG5VnE28DnTTidXv3OnKK61ORl/EbP
cbaFbDxQe3cZZMR7Mj/DQCopzO48jM3aMoorf7kK9y47gAUfoPHlUDI/bl+DYG3X
n0CvB703v8BBeIMT5m8jMji2lyKxGfgAc3nVlHp6TXsnwcTPREKzTJKzoVPeSUt8
/wqBzHGbWR0k1HS+4Y8jRi7kGvfVlgxVN+lNL3R8zE41rwYtAnm6x1rur2/slgTi
vzerUrd1w6M9nyprAacOr4I4gbLDin2FSqM4fw62IE9KDgqS7gwG2dOTIq1m8nUB
R8a+QZCtnonDSxc9mbVNDuztHdGVtCXoHTqIMeHAHP2b1is93Uz9teAIGtTNI1ze
RvigvR4ivXrXbdtd7rvTBBP/Nijb4SCwCb/8tJj6FXSx+jxYN1t8N2XKD+gPec5S
kCOXY1lhGBnVya7D6f/gfEP1gREronBZamYT9VxnvNa7YDnWVl+iQ2WEHJQNCg/B
93u9gkoV9BlTTvdVlLvxfylwqFeMElf/7NLO6ZFlRhHYPFAIt9mboE/medRt0laL
5CqPGKx/bPpvfNSgq3lbc7EImTRfbrbXAJ/cEMWHlnMkEKOmeh7oN3THzee9TtPQ
4Gz3Y+iq4dkzb9kqppRgjgaoK7f5qISZMG0BCrA00Snc9APetmdIUdBevrkf5Vh9
tTnVpIQ/xBmrlYUB++IRg8aErJLgvaiQWGZ/qy5vhM74FVYUgETrxco59yAxVEPO
JuNx587eMZ0tjcgLgUg5Y3j+qG9NzcUy3DjU+wbsx52agIe011ICP/MgZSSA1fmv
cdyC77ZfrU7+FUlOuu3xi9pfkhmIKMwQxqP2QHPgFTgIxMn3Ox0O9ivUWE4vlknz
77vh5VeoPHKb+Wxn5I7S2Z1QnSgBU6qP776NoOk1sutjAZI5A8J+N67H8kWLd+i9
mev6Jn12qzpbfz41LSZyNM3qxZWzyLpZlPv8oNtvIKGx4/0DXSjcQhg4dn6YiaxD
yj4vpVwN39NFDTVzOAHW5+2SF5L0zp+8at7jRdTDQdG6UKjFqget04riB8m7/QUp
+Bdho4NPg3SGNQ+37kB89vmiEH+xW78BYq1WN7VaYPVq1kGBfAI7iLUH89Lg9z5b
j+pEhZymY3leATBQkOLxEprCFXuHmAAlplADWMK83iQAcLR0Qn0bP+ZNql+xITqo
DCm6BcnCiDQY8hlbkWaNf/q4zs6TpP68r71ufAHuUw+RK2DaBNbMp2uRoljQNNaa
uP5q21cP3byCW+LuLvixLed6954vsJUlOLMbeBEuJm/U6NMiMCWfKRtViOXQgGbc
V2KjGE0vm1Qnk97MqoljBiLk2V0nQc3PD9Ip4f0EymzB4KxqwXlS11QlH9zu8vJx
y9l741yPKGCEa2muWR7ST/2+jeoIh4yhTzBLGIRYB7WMZ2Sn2IXiT/BiyvJMqwFF
4wvxGl/dQ1tV0MMIULKdLPUUuvkKZ8MlOTTH62oBkby07g4py7TrmyHbNycDqU1k
Yy2JaqWXCkMdZRCVq2azPYgJNdq+Vnj3vYMmkmnlNirtN051AvUeFhqWEvT/apV8
ocqgLIjlLuLK1Z8VhBKOhucAMVin0+o8fvu4SlQ/xL39lHsSi/4YJK/u4YmpTeCs
wREYZPANfjyvwdUUYuPbDxrAF6F/qief9uKR7tk0tk1vsZmNECqP3jDOU/ue8+tG
G0LhHhT8CR8t2CpmgWDI2gOmLe6zggWHH+9SNWEhVHEglwaV7ROw/kzvJ+NlPH6+
EGR0eH/fzLYSsid0k/at2IwRsxYgQluc0NuKZ9fIwyfsviAe5JTa1evqE5o9Ap5x
233b/WaCKqk4bYckh/APtiohEgqwe3rOVSsg1eUeLVVGgJuQRuzcQ1+gd/Q+ueX8
1viEFmksNh1hy4OquawdnPf0zVqZED2YEFet6r5dFxWIkNGZ67UmWJ1uMCUIipcV
dqUaKQrFimZAvV/ZS8LBd1nIwr5v+adPvcfuFkaLoKecfeQFRD1w6l34TGBuC66g
TG8MtHzSA9GQ9YFrBOf70AYwxyasYvp7t/MbYlJKZL2CjxB9K/oEwZHux2zf2BO3
+2wdj5o8xOPnCmHKCfpcnpNYApgOfJx33I7HfAOGTCxUMF1h4gZH3ZUU6dA759Nw
/RC83gizcSQVJuDR3Hp/Lv5UhinUBvdc8HI5JtFq3tUZ0fMBCEL4A0ZDSC04dwhb
W7ARGmrdK+5ylSgeQ97GuKSOP0he07a9ANNZL/3L0iv70fy1UKKE+WV8OxlSDILl
tcpiHhHNG+2ilVIVaDqZr1tk5BNrpnO14kdcFXWVP/qkBKHSaSYICHejAylsn3XH
9hA4i14yxFxDp4H0To91QfTVUkWoQsusdE/G0Vu+kaXzvpHUTdFVez6t8g/ZFVEb
NZXfK48mumcCRe4btl1CkcvGF/g85q/l53Nok3/dY0rP1e6kFABrmKkVPlSU0t0e
gKDwAW1fb8Art/f3T4/D3ZGakJ6zbyAKNIdMb7q/vvrKhzMOato9Sjv9rZ0fIZ2i
idm/Yo0ZVwf4wFgSqBC/OeNEqSAnH6xfOFUcCf0I0iPkbGWuH4Kh23BiqJEoy8+P
+biimgZinWDoyPCOj/f6k2+Be1kKE0eh/6l1oQpDHMuYKghKqG/2igck0XE//RKg
wdTubpfskPPTvjMeuR28iyJ0CatbwJkiWEPeqxeZL4D4sPLh+ZEXcEgt2n1KYuRE
NDN6+nXqYB9G//lIgONHTuUSqoGn6Gr0zrnu5SUHUb9N0X+osTL/8wlRlGwgp2VF
wwF56PUan+dLwyYcFcWg60WYGsMX2ygkQ7lPP+BnlObJNUY+Ay5F0Mm1XAFhNX2s
FqaoAV73uz2S73yXI2vXHjirFXwNCG57vIuY1daFLlAUJ83uhrIksxlA3HA1P7XF
+SE1FNeZAL8uIWyBI40J4faLLH9qJmjptXzqmZjFXASb/pFzaN0rCx63iE8kwKiQ
M3MlyZ8I1WVBP1cMiM/17zsOtMgewIpiHhvcCv7KQQpgrvJKwcqZ6aqF1v7DArVz
Rb4wZnfV5q+8Xj1+XSdbLHKRdDQeEbbhh8kVBzM4524H4n9J3rufztT8JBpPD5Lu
7W2Z1sH8O6hv5GxONpKvYsZZw3Fy8ckBpmEORUEyQ3dCD09NU3zS5av2QHSu4yhm
Yiuz81dlROifw/vH/T1l9U1ptalbubn9I3aFLGdsNwa4nuD92wmer55+rXaTDvCB
f0ttelSXkAUtANlW7CPHqUVAbUVZwqm7iPUpsunP788olpo+WQwGGvASOQ2Ytkp9
mWnKzLs+hWcGj1UYB246HtO13jyzY80z64U2aHFSBKTPjW4Ld6JQDbIW8OQi3Olp
ubk6rHRVM7eI6/H1anZgco/orMjoTAivjNlwcoNjDw0mlQlZIIuczRF/jwGAutMW
1XpccSTPTG4qpCDPzPiBmt3sucDL8FIYxkLJxIl19xIOT5jkzMaENvKn1pmpEB6P
Mr9fzizQ7TDDxh2jCUDFY16u4JtdPlozvdJ/lbNgfFj+UEo0fqGklLY3SAYRRW5y
+wMAWWVnZ4NuSvKCzn738o+4GyZdN3RGFZj46UXFyFTaqUyUi9bTYOGgk+y2AixF
Qf16Tsfw2YHYPQKy4oHbciReXNgXKBKgRuG1kfrjk0+x3iwkd1pqdQsl/RmlgHLO
SpJEkpuhBIZXhkl/xVU9BxOJdWe6E5rNczXgy2G+9XxKUswupVkzkMMdQI6N6oGn
75QQ04bISohbm1qZcyY7DT2rBOAVGdDuSrXs5cRX6B2p+siTQi/wGZdECuoGFZPH
QBRrErpciFJv+J8I8Ijfmsc5gaOY+qVk/RCqFhHMEgtoOHc6vpbk7+1mRXomDymy
mZ/n6R28E81Bk220Uus3JQaE5qED9ggCIN80WaWh483WqKcD6Y3WQhzGfX/zeHyz
CWLmv6csNHUrr2zqBf7btmKALTnaiLqysTyKQz56LVfBp8MPQfCX7PDitvV9E+4+
ae1LlY3r6Ou8MIz7gdvTIdTsEuLt/8dKIh3x/n8U1p2FHRlkqVWWRSzJI0mCyRfw
6hbpDIActYdBJKxW5U29L4zYf0acjZiNcy7qej3oCRC7a+GNMuRmBrbvmsyHDX8w
WEvTHXVX6GQvJs0xmmWzMZDCrAh6e0Q01+0dxVoMwc7Fp/wy0O3ucTZXh2JKIdm3
5I0eqfE7rpW/F4FBnnrnDvvmpTBjadJt9rMmDPsLgMCHR7urq5se8U+SAJBpzI/5
f1nEJKMCFVcqKBrQ3Wlmc3b6kQw+sc6gfRGZnstzY9R1B/oDb9ECcqVZyr9U4ctz
OLyAuOoMgrmC+J/RQlUY432duRk8gWCyBegGe2SEvxPZjQ3xCeNDt6zP5gEETRTJ
am8gkTzgayAo7poLVbO0Tf0jLJ9kEGdgNSOZkdagXak165+2C1XvoHfOjLX/c3a0
4ax1NRH2iTXu/it+9FrzgqIX7TViE4UzYjPoY0+fP4d1G+BmShWodlvzh0Ft4rO3
GV6C3K4SbKtiXE788L56/8TI5hU9Xno+F4PAEeXjzMqz52QaVKk/3/L2ZLCxP440
evoQeGYHQnYR7lDjo3XSdbuGGw6/inFRIYP0Jw9LSALjOWOWlh2KrIj2OPDxGq4L
KN3hY6LcT90OSk5M9iBHpNoguKlA4nWkg4EsmRyOS2fH6lAByeMQl9xd3xqJo1L/
29779TllnDm7Nv9VFn93dt8b/7tJbuxhz+g8nTeRdIOvmRvc8/0RZ4HBIX3b9Ipg
Pc8zLxG+ZsVlPo6MlcGlPTRiXZwucCJlv0CH4T3STMUg76oo4HnWHSxuDtAVkrcY
VASc5sYCt2n2WMTZWnPkDAWFra2Dpgiz8898TIDcUiZwpi/ufj+IoOtabLY+7zGT
AdqUKL5GDClP4ZVGZt8AS1KQkGmjRWZoIz6Wqw8+B5UR6eFbpm1ID8hZSFxdfs3Q
zDVZITTcPYk3uUFk1tecMvD701b3DpNTlz87qEvTvBM8b6E7p/X8n9peTs5vFxyw
eEM3MQAE4iB4aYjKrFNKXzMMlsJnOONU4MA+vu8Gd2Jnc7ay7urlIcXhItZiW/v5
twpseicEedVSpjsRE7jDa1NLXzk0+PuRDYvxiBRGSlMESn/2ESmvjpiXCEzbDtua
ZMgz8kCOW7GBpTPlb8uW/tKqVyjjMqVp/7E5vmp9GvPzpUVSfIyPPN1Cve9qASPZ
Y5xie+Hk0WQ0RzrMR0urkfVIf61P+ZBuvoHkD2E0iMp4GhgCftGF/8DgtA45z8Sl
9pXfAcOXRQOfFd5jFvL6CHXFN9Ui0XsuB0/jp5TE1sLpf7of86g59bjGKmJp+D3m
tmqUJwU74ZchmfMItNUqSQFObkz6vJbtAOVcbUdpDvpMh0I1/v+7kmASYaCzH4z0
+Lmxu0lybWyTdyjHNKwCNeEJGXrkT5BinwpDA6SldYBr+Lpe6RtJaanCuNboOqIj
jkSlGAoHWLC+63/cZIqYoWj1jzebEI/BVu/Kjng+VjttCfbbwOC2i+LJEslJklcN
gARRnp2NKxFdqv7oiclPEllKqpJWfakBKC6pxRfeXm1qMcozTPj2pw3+X5rRis1R
aVZVFl3UL44n7+6xinySVDj+XkQ9aS72NP3JRiZxugeYCDWuYRb+HukBr6o57MMY
00OJlGr0vdhqoLuXVvSmVKwN5x2F8nrWzSxNKlIp52c9mJZ76QQvZeC6KTWOp1st
H1nl+49w/VDxnvzx0YZtstwVS7PYOJMBvvvuwTG143GxzdJ+lWzSKMEFmPNp7HZ6
/kIu59j+g8j6zf6OPGcXjZfP6viQ77fTf3KyGRnMKOSL0LadNwqXxHq66p/BSY2g
/AIpk3iD1GfTOMbVKy4AR3RdmTWH+CDmcFgkBdZgl84IZQ+gYHFYqnyi+mdlLq+i
buWC1mLKmd8Lmx5TiKzSHeFw4m0swHdpnPlClmWK2lrxcpkwTkAylaUxu2LrGBR0
YUUe60O63lZqyNxbivhCiqGl668P9z7Rw14jSqfeMfn9i3AyRvjQkWFJdtgZhVE1
TEOA3ZUoGrSXgJNrwmrGlCKfYfMEeoo5b0Ndu3tyyi7fNCfkYz+0k+QSa/uFZeaj
jgjwXAwTNaHQwsMrknejvdRbRRiB6MoXGYRg348G4ePwPu08E4GlMkiWUegj6xuk
eGaRwmETqzNE7aBzr49Uw9zhcZO+/mUwWHsrpoCjyRveN+CdK3vkDkWpytnD/xbw
jM4lSfreptHMYUx0VRlcz7FWJ5YJNOyUxyZ8qRoek9mFXeV56Y0FfRNc8qkYLMnJ
qEgYu3T5QFrBLezv38Mc4MtDtRC1oBCIvTnnxoAEgI03TxTcEWUNFA/VzmQWIV5w
BFbOqzloDdRWdCDFq0ygag57UdiW10DUIpc9XsGJ9NjcwzNR8kAsMbOkVb8ZeD9G
5Sh+hgOTt+gWSVRU8J0hT40XCfyFxdSYOR8Clt3q8bLRbtqejUpeEPCImbzUhRaQ
LR4zvVL3Gy6kBQnieoKDH5pEEAf4R8HYzD2a0L6rwSZK7pYatZ0cDd0/tlI8EoUJ
+58clsKv7XCeebhcHSQ0EOGmqEuQPmljD5KAUHuE7zgBO9C0FA1f69UBLri6mLHR
YQo3azp9dHmptrxBBN/9u7g7QmUNPxwpk3vNK++NH97O6lsS2FWUfzy20Oj9MzYc
dxHe4ZvfyFLPqTaU7d4h44hZRB9MlM1g2GqlPw8Q6VtB6m6PN4PfjyIwRL3FRf44
6dPOmgvrsVTVnB384QIfALJ4q4pHTTL/11xYy4Hp2lsNNL5NZC2jr3i+Dnj6acwO
YOBMvqwpfnsz8djQ0VafuK+39aJDOt4nL6nSkk+8pro4B6LMf9BLQodBmXZH0jHH
BV7+uHNqQK5Z96HJj22RTbnTB+nilLelBo8XM/TM38rjgrVudJ7EbbVCjIqZZzCO
NNXurmJZ61Ocl/ycZFReEQQu/bLwai71uKHgCbOJ6ZmYOa9jT4MaXkj2H+45FL8Y
EiVW/s+ei4L3AlpPOhdtgk1CQ0aBJVfzWQT8S2drsE0wWuCXi1jGZ4SYMPGGR7Xh
9AaXwW1/c2yVn/xRNEvBDs1J24USD4s9QU6KcW86cnWL2vIXz3NCDlwgyrBp+wOD
yKkFmCEYKTz5THSD40LBzvL9FAjmrxGFVs9FCAkAQiu+HBcL9CtjxZ7VQa95gIDa
sddNkTp0kHfphEWavTLx19CdRVBCXAgkuyjEtW8rhS0DaV1rse9CWo6krqFam9iW
oLPVlWk1rEqvXU4GDys04VQgPeOcksl+Pn2cl+L5xK3RSyHURfHCUYjZ8yQsloWN
uh0hOKjYQpSS/WKlLhbsCfjenDYJxqX5TZOJJdKkBK/g/GmCUHCA//+oI9uKCrHR
O7B5QasVNqymgVyHG0l1qpWIgCaCbNLBKAywJwDmXlwPmx0z1FDAFqxbaLroWiXv
PBT72wPIAPrALdadCMwWm+9fKI+p/MlfOQYYrbiAb4gvqkCt8zKQ3hJysFnE4pyZ
62sMhUWBA4mN/OevUrthoBd+Zsa0gt2nbHEwrIDDUP3kDoYB1dYp2N2mDlPjhD9l
nDo1LVqNlC09BKTxxO0y+BcRu50uSC5TvNaby9pgrfQyybIbcquih+tiE9q5tdNz
psA2WHFE4k6kI6Lpmn3RpCa+ci/qPiXBzHTRF85FKrXB4dWRnh6L2C8xp3Tc1KmH
opTUdXo/QuklMtXqVElZRZ+oEFYGrTz22aLaX+ZwWvdvifW5akDVWYX2D+gvRtsx
nofP7ggT7YHvl8tZXSzWrIXO8a9tRShjctKyVytLvpYj2YRRZJcMikhZIrF3TPxk
rvltR8ZdCqVtR8lgwg/g2OHu4n/8R2GsRGMwSiYtnX6YbpDiPZCp16ZVBKyxutav
LKH3/g0EbAExjvOYm3Lm1jop345AYXkc74dzhFH9scy3tILNWZowRWW89hYsWgk7
FUopnY5LBs3NRyHe2afXmaFjQ2VxAR/m69GCbWuIY4iSrku7XBWAi8UUOka6IW2F
LzJrkjFgIRWATHlKsnz1Z7lJ8B8HNUWrsPkfG8i6mjhyXlbALRjxd6XYuz1/JAJn
Rh/J5pmhdZEKC0c0k/Y16oFSJ/ATlW1es29oqYGNq+xcAUPxUKKoY7xjuhC7Ylws
xzETUMvl4jlaVrJUAYbbw5sEVYvnRMrCQYZYYVDQe7zeICSB3emZpAm7T5WckHee
khIWcjHXB1CWnlnydF8JhyfaYtbCX33JKhAF9H0rfNzF9G8R2DeqYIJK9dIT45ur
c3NmiBun8/rqGkyNKFXrbBrFRS2CGMu3NK/ffqnW92fTWHJ/tvdhVuNRmZUJGihQ
1ouraydCSQpQWkQuFdplArI586Qy4fxxwFAhy6lA/OByGRLPGNnTjuFEqVGcjPWz
eN9zJLL6Pq6Qp4IeSSgG3vXFtruliXrGqBMerW6w+i8objmr2ArMC++U0PUjyvKX
/S1ZsmrAAXDazqVFNTvgtU2f0+n38YsemgP4Xw518i4KlmLegXmm/DXGZoHQo5SY
p7x5mkI0OEGzxmigbidDwEMvBG/3RVT3YZrwo7ACU32KSkKvrX48/0vsjU24ekvT
z4mbe4KmKq7DWeMWgwG2AR9glTOM8b9uwgVLWGnCsZD2IH0iG77NWeklJYXQgUGO
8GGqePceLqmSA5t7261K9Q6xdxFm4uC34nqEyblgekKB4/6dbd217rGgD1kzs3W4
XZTFnnrB6ZhCVxax3Qg/xs+jTO517WUkbbw7CW8Wto6rbeNznEqmHqWr+7NdZl32
uoyTFlegEx/BclKCkXprvXq8mtL6cwqVJE6CL6sFm9j60yFZlN9OV4xwrsv0sVO3
9RKqbAw7+iqCeGH5KdBhVYQn135rxgBDPKWitxnMA/5zLEXoX3/tgjElomuNT17p
plJ/t111J9ykw7lkO0Lf8SQMCeORwKrgU1MwHITDl3zpoXlB7dFA82s71j+gHnTx
yTzRTK73KOuBk+cG+gJQ18csW+39E4kzQjEh2aulzzP8YopmddZlZ5S7VqIkFmM4
sa3x/dO8qpLAYaRk2ddri95jp0E4nJ1Sxv90JPOvPAN6mHqVljWUkkvx3YbOOnR7
ANachPhP9m15Ce5xS8b+v/c/bjtWM0OEoGaJsk2ilKwZUAJqwgd7QgtOZF2tkbte
PLI/C05zatYx8ULesZkNN/6rGrLo8M0ZxaxMYrzAkE4AU7xOXThM6up6oCJYaMzh
diq6Itqz9gnfJ5CXN78zyh9IkY/Df4FFqhT/LsjdhGm+zlmjriMYh7Ep3Uh6AGae
5mPpjf8IagjXwmNFqKVxNiiIjrqS7VlyyCCnSWKq5SOG/TxKGiSAmPlA5n8OGw9f
SE1QFaqYohcr2vhoDiBOjDoPljU3LhM7uKrSn3Ddn84h7H9zhyRYDDkbX5yIqsLF
m/rRoxFkcqtoBMffhRpz58XEjumTjhmVsj2mYKKc35dch1n0KQtNtMFFLY+Ki/Em
Vx/3/okzAz7VF80toQq/rXadnxTD+px98iSo5PAA2ZrMeg+1HbKb70oTmSsEQvxK
KQlfb9TmKCF51qwCMN58Ft7TFbkJu/fI6FvPBW4J54t/hiwQBQ39MDvSHf1O7s4A
x9Id38Bv+i+YrHgfQQXXnm3XEiiwR+xm8uWtsKBiSNjNk+nAFDbgZHMxqgW8Co8v
pOld2tO/rIuT2x3VcSGYFa41S41y1q7LXaz5FXw0CS1oxf/C+wCTakIjfIEiVJvX
l20MJ6Pol406x+V6x6r11f/Ki22Rp1tIzeqI2l5qBN1uAxiOT/DUK+gGkqxZLOYt
CyYT9vTIndObOfLA/AKAz5uG+YYI9/7ybdjvhREa5vj74QTMeWFYs4jRMDANw3VS
lmIrIY5Y0IU2yjQPH08OQjUhuEPxf45mkfAibiOyRcaw/zfWKdGvxEIkunX/4iMP
RaCmg51o/kboiO09ZEhMzoEIBotLF+ey4RXQC0jyObEY8oEB37S5x6GUt3HkDVKH
9h/MPSu41QE9/UB85btjnlFGJP6XplAo6g1iHGZrpAc3AgFB3PaUVGl+T5+Zp1JU
Ja2Unfe463vgubS+DaeaoocLiClqryjrJQvei3oaRvenYObpZ0xp1LuDQ9pfemGq
SVkyn7FF65ZQAWOVyt8aWgkmjy+TCwFjsxemlYrSZ2X7HxnMV4EP9BpwK+qoN3u3
I7Tze2L6NJzJAOrdLV8PTKVHf8HV1ZV3YG/tVDgBWBTInqFYcseJkQzHeOH4+MCF
UzHYPP8TUb2QBhFpHSn1/NTeRuDqE6+hl+qfgTqxkm6qOkaTSxdR7EGE2Eo9ML+e
SWwpgITyfxWtJ7xzJccVj7gb2saHhygdR4POPqkuAoFW2K1hnzCwUhGJj+rmwRAh
rFfISBP8wt6+J4v9Dt6PAGM+YB2SPNu88fQsglu5X7BK19cv/HOfAK+8Q9sVp6UW
DVz8yiUb5yasICQ7gwRkzBO6/9ER0xFcTLfUuuD/gWcWCEGepGh0NfHHRotiW6oi
y233FBIbPXwDmQJOfQIHM+mBVm2zbe86gYsxs7+oEh+iVT4q4bS/MWW2jZp6HRD9
Wfk7vG7iKZah9vWcjl3B0wdaJ8UT8IukWk1ZlPMDwDlDB8SDMrq4LuQH8gJmNNL9
e5opTgKFcwfpm49QQvCIjqPGmDqQ1Z3viI5rm7Xkxo4LpjXyh3gVX3Add03ZUCCu
ZutLkS0gStIGkAKGOlTGBRWl+4Eoxk2PL/sLfwVacS8YwM6wo8C9vek7g3Cox+xn
ho/w7i7pTHJ5gFxqS1maNKOdzBaas/fXO7BQTZGpw0oj7NXZiIat05L3pZG4E+GC
q2kau013PHJ5ShQyDhmpqZblyewq0zMUyifnp6Ae5LGP+Ou0sZipimjgGoaYluS9
dMxlAtaEoYPriFj5DgGFt3yJw61x+AIUmRLRCxfd2y3Wwc4Iu3n4B4u4XhcaRPS3
cxEb+yu98lX/YPasSWyGWfIFJrlJNRjztWqnR5Wz6Iw5X+axkXQDfywnfCVTs5LV
hfMB3zGBU8WdbHXggEjD0WTVazVpI0OBF14qwcKWmCintJFzAiZXgYNo19sRCOin
JctYwvslCib4KxF/lydGdLaAxeqf4X3rFFb8m3rVHIum1EcvDr4c2WWG5VKldVts
FP30LWtbOIvWA0kIRO5cfWjPOM3APUVFKDWCNs0AWQ3WKXcnuPUs6idBRWQ/7hxH
Ehw89+cQ/AoK1bwgEKyi+X3mcI+R6skmAkAlwcvpHPePUwDXJ+szZMqWUacB8evh
G4lfWgJdnTyjSUrsTHCzfSwtuzO2kPmcg2Z3jefCNYraJRSCBKkcWDIVAP6UqdJu
AF5YtMSjudShGgswPx+z2QaGXOUFAggLMcU0LDJM6Rm++eS6wLMYfAwolweRtfdi
nve7POcoMA7eQW1Z97Ns3HYwHFKfIZ8eJ8G99+xWXJzkiCHSOIObZl7x4nex0hjp
j4XPnbjhPSbvOzYvXlD4apX/Qn45ftjCk3SxRVQrSUbMStZaBGbAB0FVsVVGRmhf
X04C5LJkvebLhVmh4SeUf+xJeB4Zfxgwl4VpKVPj/z0SMhI7GJVje9I82eGeV0mi
YECbPTCT6Fvru4Efk/S8zD0KURxDvzCm4v2FCNB7u62iuB2OC/72v0sDGpVItzJ7
aI7dp8Spq1dXfLWSLaELdNE1jq5Q7vWK/X9fltWT8kA2rs9w4dLajUv7XHvg2KOx
zWeRMyEaQmhDVzvKWo7v8lREx5sY0/t73bYcmiTUt762dmVufDLB3My6GbJ05P5j
vItDZ9708hrUcTkyZPFYK0NFeCFa22JJdubVNGvlxYv/vg+vVjpQClhLUriwt3Qe
b5Yi9iAfpNDE6IbPznaNIrzhZNstjNNXtlniM02/igPk7FzsS5Yxlum6LkvUFSqP
6/uN5imIcjVe3+T2rr9Sj0zNyW398KpS4LH2ob9o2ODN3KnQ/RrcXugrKLx0mzNO
Ve95aJtwYDyQnGU4vpWDNr2ghqXMBK0c8Y4DmO6pUkGisaVDxa485LVjEoMx1Au1
tgZntGc6xwoOuxUpAnq1RZ4fPSakStGQYE2XXGlNR6lOAAaJ6Q6ysLsihKwdy7sa
T1pIyrT8wad+bvE8MnflkQVtDWFMYutE9ilWZaWg6sjWfoKkEhzRv5YDLlZS4Cp4
ubdlkzapQDxcw2VRbovGZcba9OVRnFu/cDTNKBiH8ZnKrZB7aT/0p6eckguPuYFh
z+64Aincmr7+WsAJn8dZ4oTIwlWJJRXDEPv/hrNIM9BimFl3M99vHxzfOsqiDjc9
YdtCwnTaFtEPFA54ldf7BrvT05Lds0QZajPlC3XjIVUq1SCjr7Kp65a+WopTzged
kelBpddNaYuZi5m9FMxPKQHDDNLYKDpC+JPQPsZniqeYuUUtDTbmFQVehCP12AH4
PE1OKRu3g/kLX7FCHrBo/DmELBe/WaPQX4zXcy9NQdWUHfaKwLuY+FR2sify+Msb
yQmJV4IUWNfVrMpN3NIijknSVPvieh4U/GoVsSnOdAEbWr3IPlZ0JioYyuL+8K9d
9ROJhsf1kjaUSptngj6Tw56icW8NfztVG88n09EitMV/m9c+0bhJAkxRYZn0CvLt
sHoUgmXT8l5g8qWz7wxOhZiZyEC/+0+Im1I6etpnlmoEKCEBRJxUr+9JOOkXXYi9
0150tx1Ff0xBI8eF+3mJ2VimQSerlUfAReXkHIhpohXsIDhZ4i4GU+MyjcDl7pS6
nuF+rvUxrEFsov/HfiFqrsEWN6HPxo0IACyI3rKo0JJxFzbHuePSBYhxPRnhrZSx
+3QKmynd2iATCpzJhq9c88kkyXTYHxgKPTYWDgLzXagqleA4F5qLPowazRLaYpoI
0lXZO/sDhjuKiWPWppfzG06HS/aM2uPLDEXWJH07BK45wmBopFoc/qoOTxvKIHND
JYat6d8WBjgnlXOSAhdFbWsmeYAyPgG8SJrSxUM7z05yTvYu9fuUJURSwOUQT4eO
MmZsvdkhHza/9wduCU5UABaXMZuHNks6Ujq/yinV5QFUPN4mVvAgPUOExIG4z9XV
jxWB/MWMj/qrPJhJqUxg9PInVokrE5rqOzzbORt0rIALEMSKhJ7sTN7kdEe/b5a7
x8KtqqUB9GeNSCWkvn7fGLLgNLQB8TOXWeODjK43aDJnEY4IXCCncXMHpNIPK7EI
X3xKXSnHpLaCiKFeUtfj3JQeP4vtNx7h6t+DfrFB4iHsl0OGxmPuremoHY9Q+/2I
AuGuu9/Op5fXYQpXj6q7JWPu+K558UehtGAgemjKkSqvOhIJIFoBHeni4iZuq/Ne
t3qs9i6FCVGikyZL/cerHGiG6P82jNO8ozMGRHivuvLRtWrgXz/VsNz3FdY8g1UJ
ZmwsA3/a0Ez+QR5yuaQfaAICvGYjFnWY/3yFE2QgIDFW2+HCUZUKcRHs9/Nw9syo
rAZ0OqfBNA6atPf860o4+SxRt2G6aoAySbFHqlbUn57nkSEqA6tQ19dBkYq82p/c
2s0QAAJxLwwNbbjPSe6s89qd6Qo7T9b3FWrAF+sONf3AyFYR4VcSo7mMi+JRxivE
6M7T9BG6SRYSzhChi0PXUMNPKXRtRP6+WrwfB7v2+CpeS0OYwfrDYnTzoBUbPiPu
rJctsvTxyzjGun076MDfg1GpgZCCMehkUNCbWt/SKxbxa29zCeKj9G2HKzbbBK4j
ghrJcSnGnqSbRURVYfXsafJ7BLfiy2kTn5Etpq39EM+PPEL9FHraVSyriaOYfmh1
DlxBhu4hm/XjXs7IkkoAM0Pjml2J0xbVOfEiVCQRBgKpoyL7ABPC6gt9tKwWU7Y3
oH5YULhlRu+QNHX7gqaW+J6yhGrViXrf5KaAOnN2dSryETbykGkM/R1IhfAs9Jbu
e6vho2x+xJG40lkNhSgLChFk6r1wV9Gcf6hGkgLmw7W8trxB18D+m1cZP4zEUEFN
c1WPaELV3gCidmFoZsTRSYI6JIuIc8YKD0r8sQ3Pag2tNdSOKrhxvoMgHX+9AotY
8kIUdVFu2ekCxOwMS6WETqGs//KBAZCxYxspIBIiLwgyv+jl1snVwzjbBjoNRKBe
HzB+bckiTaERn9IRqA77PP4l+DXsm8wIS80CkH1YZNV87RZqkFycwl3SzbKpnYKA
4gIImGn4DwEORPKe2lACXP8zTpYpDQoxpS7ugMjiLIDQWwyDbzwtZWZTVlubTbH4
Y56WHjYOWpO0qFarxDKRGH/Z5ddap0XkFnzrFdO8ET7CCX2yFSV90EjsnvvUQlQT
lshbs6RMw79jMBvPn4SFO1zEcnpp/4zEPDNVMVNJNiNjrb0KlNQlPye1hpPziRi6
qFT091HtLEQVwTsk9STJclorhDfh60M1ss2ninm0sJYXe38TrqFl1z8qf7WLl1NT
o72OKjx78krODdZSyAB1PcXftNuqyCOtmCn3ml3p2a2N5Aw0zjQGrstitvZXZ8Vy
TcCC2SQzTd0mlCSMbZtyMYTt1v5c38CXn+V7i4eu7VyaGN9lkwQ7eG+2dgZUi9Fk
oFysRDcODrncMK8LsPZVNpawtVDzrTUWiQMJuQcyzRT13Fg+zKwSNq4VmJQ3tfX6
PpIygW5zo5hQg6KQpXpIvZhEItli4a61O/IDetLjs8oLjF4Lt9MMxbVn3qA7ScVF
NZVmK0vP3T5WksCxs3pccCXl1FnBND2cU1IKQXrZ8jmeuphtK6S/47d0VjMDWQC7
IJPQ+z9EUAfgo0DuxCt4v/C6fcgJAd3+xRBIY0jHB+SHPbr4LUHOFcSEsW2FiMIc
s4iNc/H3mq0+JWEHxVNlmvz4wEP4uC39xGbdNgu47YE1r4g/SMSQDyByynNjamaq
XUWvsPRiczISDBSFUWP5QccBnuMhYhwUEIc29pTwTDHQWSA+mc2SiKWruvip5cjR
0vePsDOob1Is53fWRDZzq92wmz1H+jEnw32eLRzSd9+jMm5fmjhvk3iCHRShu14I
NK5stYNJ3CF4Do8hh77XY2gJq9BlKkmbfYJD3Tvs7x19ob3jVrE/As3PRKAXGDOe
LlknaNT0YTsafAof8yJjOzR4TgNokJGZvsMW2efevmJK0W2t/IhzGsw4jUD26xos
QSPQ8Ob1R4VXjXB+GmtBNQk18wQ5IyBy8WSASd1S+lcAR4P0BL+LaSW/si4coIJs
G9AX4zo/xxDN0UJTqdn1ig5KR+IRWcwB231w8f2E5rXHjUvnEvy85JkaTBpd6Hm/
EGQpv4mPwRv81t5MXNgWyWN/y4oBnRtU/a6ehP6qNW2T66cyHvNaHYuvkO9ZQMhF
9MONQIMRKWN6PemH/beXT3DNQ/QpLXs4d2/c45jM6xHiD+SQBv8psw+gqg3sd7ho
2QJAk2kyV1zNMYRAQI6TmV6cFhkV9XLF9QLPNdFNpZcnDqur+B80nvMbPoCL9VzX
aVw2iHYY+ydJ3r5hHpUNqsyKfoUDVJRjSOAYJ1TsFLZ8n+RSbSJufGlysmyhVQoi
amtQR+fb2hAJFqxjlulJT6lxhBaLQsShZ+TgzWjzZGwbe0WhUzZ8JPI/naNXEStA
+lX012KmT2ALJ91bF/1zRyTIL2XK7VPVSkpiB5GD8oe9hWPeiDmCb5EbK0xaNtRH
y0w5YTlcrmnvzolLY7IZRDwHX9l92Y54U7JBr0bMPrBl5zBRxdlU4PUNngH4opmY
iNG10NElsVLuA91oPKIzq7bJiFMDImfHEvECk7TmhsSu5CVliREFiFEgvyQs7TFI
lBEVCC+giFo08lkJZkyyTbsBMYJ2Y+CYCD6ZuwKgD5L7tHfsH5Cpfh2bDHQQtXWU
uMHUpCdKn1Zz4XLTVzG36X7BEuc3KQNn/BiczgmcTcewpHBKrpW976wYZNsROL2i
LdRxX5BLQS5xWQD8euW67e4BSYUWeodYQlg3I1Mwx14CN1o7sTlOFXmGRtPT/M2t
+Pc3Hj5/RsgDpo8CBo1WRD19672alVL9K5V6G8m4hfHK1ytiMX8Jn/x+AE51cmqx
f0uX7eBexh6MZghv8Gd1pfovA2ngNMmUwUA6TdVRAZIogSxehJzIqTJy8aCFcgG4
c2F6qQiCk/P/fZnQc4ufXE66o5HogqWwOTLXUE6RkOvcCpfCAiSBXtdwwPh07yXc
8QkM1KJLme8lplse/eKAOxAE9DzrP+2FgkcEQ1kTNh3IIHjOiQsZJ/FDdGGWJwQm
HRXMvtXBOz8Bd9f53ehxPS2yl00YSqSghbFOkE1iVq9uO/X0T6zQSjcfUeeqkvSv
CdxN22jA+SGURJA4nCOHaFeRsaahvIujKMFAMAA8FNo5HtiW1hTkJi0e419exuV3
4/95htmO5/Pkb25NQx9oJ3QosH7tDviyXHG8NdrWNjz9stj67fgbmcSWmisRbC+x
lduDllIVec38otXoKJDlBkgjy9J25vmcHIXn1aQ1f9U2hUdzqJj3R/vXb8192Bn4
CKP9NhA8ugUdS7fxjdtBTrhRwMqsfn6C+sIHFDYlNuv48o0rowiV7vz5a8jJ4n9V
T+8rHHKF7fw9utvqdV8S5Xba9Me2We5xx6zvd2mdKHuK1S5UMMi/KC5DPeKCv5MS
/OqH6kyfhuHTSdwtWMdgnn591p3FSZXpYhHcwiV/yTk0xd66qlKntaR67bpwtRO3
pwgsp7fBEGsyQ7B9xY7kd3o4DljuvctGlB8TqM9nEN5WEuFCexG/ccv2zJaMvKow
nJNAQXdkYnqKDsRrsRNykE/lJD4BH8SgDCoftgkKLWUvprk2iOyf8rZ3TYLP4VKD
vM7nQUKoayNQ9CDU+0HyRRYCIRypLHYDqp/IKmEwGRhFy4I9trM1TGVSWXXJIcx9
bKWbYd2nJJ+EYWTPD1twHI/BlhFjLiHOjDf/JoaOQF2ISq6cHsbTjrFjJLKFgKlz
rxgdQ1iKpGrFINlAD8QvSgOR4pshxMQTCYoOKSt4nUMvP0EKgH9eXdSUBFwsxxFn
bJRJ5y6ArBZGtpXtkIYWD7Km4eU/nkHR1AuFzCAzIx651kv8n+tunTzpHTIqjGvY
G2U27Zvc9uGJQrjhFzRHzzaNvT5nC+Q4yhmcqjBsarioslOTfU7pvz6KZF4JGiU5
ekzOe8ynSRl6SQaXvgg0U24CWlo9MswfPKG1fXuZj+T+oHavuZtDX9Eupkr70j2+
XjfiWVbseePgqmhd1z0wn1qQxbXeamJhLkExu6fllOQ2GwvjRanlvr+ZJ+E9G68D
OFipaKq0ihUMTorUvj5rt8yVtVXuTVJDk+8DdtHqa6rn6Su/g9nCWImG8+/lPZcE
4ugMyMUcZKMDGyLhXQ6VxxWq10W3M73YAjFH+a78SGof7jzImkbX04+G3GHuZ//3
QavucNjZ40PLbV8QypnZDddqrCBhwr5YD3gXhuh4yfzufqsfE6eR37eIcALsabaJ
uQEFdjSi2t893L7mbwgpZOgwwD/f5pFe3yrIBbaI4LWRgcU70OYuq9InletpbScC
wzsxL5A1NaQTfZb6fA/N1Bz/ztQsujbjWI/bqOP+55EV3SpkJEOx8GmMN7eVgB+t
WTwclKwUH7SFWVYplO03XpymBG7nUGAgdvRW/4HAu+vqDLVL3l4E8qalSY5b5GZW
1QUBcPut+kBQ5wYpj/IZ4F19RNhVdWGRR7++Gjs0BGpUZy/2qhiAbOIHPpChJ68i
zX5jNjPSbL1XyS2/MuFw3qQlntxIC80MgnyvkWSbN4qHuZZjS1sE/3YIcCcYUJCC
ZIYSMDVRduiMNcHMCjkHYR4cmoLefbKlsE+6izZWQJ8Pv/XYxE8pQzzXxWgty88w
D0GsONpMzlHaGjTZLWTpKyG3IGd94APSTKH+3zCl+HJ1+bTwXLXXOiuLGeZfrVuP
AyGkBZoeR7T/W5Ts4qsPauYZRtR4UF/DknkHgMEJ1N0m12JKPLcGCs5Ipp0CTY0p
jHjVpphskOeAHE3nBKDgjVptnrHxqCcI914378AjaTKepSYsiMe06mvtT4j0M5K7
vIx+OhG17+YvqsI6IOUfpNpSMS3iJ0f7Sm3Fxk3gCqloPzzlhgvpx8WMPc9R2yLY
TNQpleIjViDXBXn3GC9Mo3VQ15C0nsojsTlpMZ69v/kK+jkjNCnGYLigt6P4/fCH
3j0uWTWx85RVDuBgKgdHRS6No+PGClzSTwm6NhuWWZPe8eOVTRdH0GjTVKjHKL6D
eAUEKRoTEvNhPRykXEs5FIKgbq5GI6k7GMMZm/JiF2EnDD1NHQPtzMPh0rhSPsvI
2fhuXxHm1PB5WvIsClgBu/uKluu3IyIM7dSt2uce8RtclY4ZLd3B0jQHTWx2iaw4
Fs0XtUH5cyM84rOY1+HwgdTgOUftZWwIufRMkRSUnvdNRU0kiLWfno1ONoMLkHnm
xwcnm8W2hQxRgP3yK/iKLhjaCQ3t183cIxMSHsvmroGf4rR/fyJflBXAQE7y1GVZ
ob5iDmI4QtNVclZVTJJ1HEOIdt2UwlaJyw34P6HjXuFu7byOoOce/aV4teZq+Fso
j2wO28eoPGFb2Q5d+NSA1w0EVzM4u5fptJyuops+4F6IRS3GleouExjfCEuQhsLM
JLjr/Ji/eqEfpNkiNye7hjePiBqyBhYK+bBeqKF35HL5l3vehXpcqQa+H359KXwz
fPGabHskjwxSmOt3D1AjI3nqwcAVvbJrSwYFzfl9mJsEu8Dd74GindgsggqJBKfS
6PGmF4bPu0E1FY+KBnqAZdMN01UJ3gKARVMwPJVdPfgaRgKQ29e3GkgGykG72/eW
8zsoeLBohSWzOM0KJM6DgGG1bri0JGJ+/iiagxY7Ye87n+dr4eSlSsVGYXHFzCpX
GGLbdQ6gm7VEz1Ko/VsxGFx9sJJr3PWQJ0zkVGJBs9pD1R2K1shE8tnB0cYo9jLG
zqyvpQZ5tpIvnACd2Plea2rz5lgkPQSR8TQuVU/qn0Dmlrmiq5ePSbRHe7Ir+DK5
2K6uyLXCN43sdcUiLUdq2mlIf07ZdYvqfpuhC8SJqAdDaw5+4NA0HVfjLBE7dW37
89LQa4DcRYMvHAdzm6bBLeH9qAF+zLmpNRaDlgLyT/JUjf1mSX15AipK7veOOa/D
z3yM7aWw8lLSb0XJJO3LAuNOrrdAkXEdIhuW97czb4cpqRy/MizOXMwYWC4eEUpU
y40l/4K+CUWlSyCtW1LtmAEud9BivS4g/p6zsQTvxipfz3t8kJBJonuYUchXynQJ
Z4oThg4BHsJQpcrFSMT/c4iT2CARwIGXLW1aPGu8fiTT+uYzbojLwfZNaPD4zjlx
1JRIOsiPxm2Ym1KeiYNJkt0gl/jCN9YIq8WSfpjBKGZrmeL5hZFOsvCk8SzmEr8i
KnUkXe/ZVXE/jq+nheV2+xEmc8EVRs8Gii2nT+Oj91IW6YBSJinxl7li/K9FseEn
rJS6/xSfE6m9Cf2FuDF1aUir8aQNnQTtbk6Q988sdBvpqeRorJyvYqtXEPeut0IS
8IMeJiwGqqBakCkViudzl2hNXv6RHvxj5GdHsfXeN4tqm/KQcv/yq7UhpQUeqLij
IHQUIziy5Hq4sdZF+55nQPyJz1RxgvqlLliOHo4INQvF/+L/f7jONpt4c7CCg4XW
fVDQa/qLS39g4P3H9GGsPcRwbmGsUonI3trWL5ip55GqIOETs9IcUZQrNZZwoCBW
hUoVhUHGTLWkE2lO+St9zWX8Ooyb2IFzdayNJ2b8L2dqa2LqYikH7uYlN7thkuJs
pjKAjvMtFITVhhhiEK/hB1XjP6yGTHWXDSw2rli4VdogyFnFvIUZAzyuulBhcvpM
3U3qTuV63bRLvhHwgxV9SlEC9fWqc+x9fTsP2XPk07a9XA2KKOY/AEyBrl1JUnGc
4NqaSZd6mrXKe4nx9Uod5VTDRpmCYgldHkZtDXf2ArGOv2hkzIs21os1X7hOAC+I
U3SWx88fSa/muU1Tw4hsllTZxvlt5hsc66VEr7aJiDeivA72c6QpRicKZHjo6cOC
drhniMdJLl044+C/c5kxotC8uVAOseB3LeoYaUibdM4iRvFX5m1vetqU+tpQXD2t
7xxyWOkoOWSW0A2gsPXArPia01aPySGIdOrO+EMXOgBCZRj5leykWQDP6CLx8eTb
W11Alpu1nblzBqo89FCSc/K9WSLD21EG0BwP4KCDGPDQ2Qe9HbQTfeQ/T3ggDkes
3+xKmbMownOccNK3zqE4tIzetxGRdGNR6G0ZzqUB4FhD5JA6t8UfNMRDOI1hakzf
V37zX322xOSmwGMvxXOLdj8qUY4bw1w+wo5X/A5XadGuYDmwfVRShCJvrxHS6f9L
U5Y61vrbzy6bw33nhnifPR3R7Cno8J/a353PDjKc0DSp1GNIzMAGiRQhax+TcVZQ
0FZ3vx0S1VwwadeXAGwoAb1M7YVRkwNyKATIrQiXvn9Myk/PpLE7eXTvxqUFCSsJ
axG6SlQXT7Mt/Ooznt5ymggmpfUWT2p8ebblWqJcXxxXA/XJLRw/UQyxyDQsgcyf
GqCwJvLmGCSoPvXzAJhWH+dGVqyXnEskUeLMOSWBXOU2EJj4h0mQGEffrgKQgfaS
4lE3AtT5WJklfG/KgFO1ZZqz5ak1hCf/7eIhkzcyl4y6424Y5ga96iF28iVo1qRW
StYcFo8fHHRudfwwOmKYTi+PnKZZe6zOpR6E5NQm4WFd1qFyaA0wndayW3sF07xn
kPEO2sHnRlStc3XqMnipZYePWLjgMdCN3vZwhR/Tp2gCUIP5+7tGqt3/afhk0k5w
PpRDmLENVeCST4/tfPOhwKV3vVQZD2nJutBWExU3OTh+0uq0qJW8VVdK2xYs6Krk
Zv4ZiGR4KIdXtmgSGaoN31HuiYMSqWLuP4HL4i5lq7VB14s6QsaMRTaVAx1+4pfO
VOwzkd6+zo9BFE6JQQu6qctEVlAN7hi/Uvzaoav6dSt8BuF189kjN33m+RVcq08r
FuopcGLrDmDSt/S9ACxnMh4YtHVSDoIhAbje8r+7dTtfcg+OGBAh+3nw/ZxCuhjt
qGk9ykUXxhqxU1/E1Nnk4jXDaLFIZViHbhsILn4m7zUMoqQMRCopnvgY6lExmWtz
miOFIIpeKURP9imeGXLjf6Qj793rjW1gLoMMucEf4zY0VhQL/CMASgB9wDKAaA8f
MmP2aEF2pgtrKDjddqTTHzaNFef82Zi/C+ZVM9EVJY3k9QJq1I4TbjlRsRgRedL6
UJhfat13jeyNJ13gl2dRzwyKV1BPeqtg34K98k7pMctgeJjtASGiyxdJNA3Y27ak
vnsav7Tc1Nc/5i0nhcORu9BuZDviXqHEykv5IHcp6MvOH/tFL/5KSRM8x8hh05AK
/gI0hfm0eBgNXwQKITYFPOZIXDksbfGMbVehw53I/hRdynk6x55wSjJqCKEqhHc4
17YlEatTTNXdegXn0x8jlwKbRb+u0mZRfpGt1mi+fkp4FPrq+vI5hcaRE6UgFZ2z
92M4QlanShqy6i2vW5DyP+8GgR3gMS7cMFSW9+lj9usT/go2hxKeSSNhkporurrJ
hbAl8LUqP4a5nNReefEEcwDfHvpiekbalKt49BdCL4rSHUK0v614BQtb9rG4+ITe
BW43hP7dHahGZuW2lb8qVSvZfuKJUhZIS2rQI5ly0lFWSHBMa+lAFEW+m8ZxyAsG
L4iYdH03pHtojMiL6Ww2b0QYUQryYTm+PHBzBYG/9cdvOx3jEjbsc14ccROtLfcx
V0OLEdq0ZJhRnpJUcnD0lFwJ10XgYKHu3Fj8qMbdHQYqNjyMFUZafC7AxzTUpWm7
/4NSpHM1PD41NEEubiDT7wrwlSsBj2ezOjZVL6naeKYgihHCKAT5Yz6S1AFOVCgV
5skyQhu0BU8oGs+jbEg9IlDYU7MSFb3IUzNkSzWnIHR0ysIm6qf0fsCIv7xHjP3P
uLMjB+M45U6eVGz3ELTTG2CMa3SeMFBtWFfK2VS5OLafQPFqjMy5I3KaE7Qh2Sf3
0nkXm8cEzemKHGcb76CofklraOPJFqTykoV2D/v7c5oiPeHa0+zbqwVi8+MZSTt2
FqeeghDspbaZAONgNiqBxe7C+WmpHgjq+4PDhbEEc7g60n1WJwDpUCg1I2amlSZ1
izVBGxcFDPVsyLyaN1+KOYNBwb5dtrJAOyo+Vn/0OAwdMh0KqbKEtbo8RxVXtgF2
C4j/TF+9Vpsp1g6aQBWBC9sXhQ4iJ7YdjzTR9e2hCiWj+BoLJvhUNEIRjLq9yFtr
WETdAvll8yPK0EnTOJS+qWZ1y+FrEkmjmxdhiyKfydVkbIo+KDgvQLxGodxWNAD3
6l5vvpXFNxU6ANYVHt+Tq0vLDdArLNmOSzuPGUq9YzqZdxNi3IJW+isGHKU9ntcJ
v9cJmXL+XFuPMSGHv+3N2gDO9Oe4U7VPgPsYSlkgP00jzRiWjT7BNwbUxQCD8u7S
pdNNCjb71ethlTZdXhhz4GU645lY/J6DnkiW51MtJ+q+jcJFOZ4707PQ4JXV7nc3
KJGTCDuWbuD9mnC0qvrMZzp0uFI6J47pqwzdnStYaHJyssAQ/zkJg3k0nZaR3xAb
o5ATw7b7SGWA30sIO92lbNwCxfw1GNJqrBBwcpZ+pE+S5gzX5+XYfFpG+9rbTkR6
iAl2PLxYA++RIdAiz54zXSLIBXBKjLYSWkPiXY9lOOvHMjdCEyRFMnhc7pH3/vuJ
lU23WdsSrfxV3B5e7488+M7ebyDncoaWDCpMV0H4t0jE7vJHNb5g0a5R5AEakbt1
D4v0PR39HMxtPdp75ZlD5vKTkcZT5UnVF0eI2Du/Vpav94KxZyzmepqtYHEI8oX6
h6scP8JFaXC5YfrtdtLMsfcO4XZfCve0TNuMf8OWZ4S054ovF+gCkTvTU0iTtNM8
Cai73JshrnrcZWM/KVhoiZ6MAP+WR1PIXAqxcOSdm6CuhNRy82mY062xxgXIrrc4
e/fczDQmYpTvuZHB41fkqMvjVa36G2lihGckcdiQShTI89DDfOJNh1wwf6NrhIIC
no0LT/N5A1FdYBSiAd9M2ktBQx6N9/ff8cByMcENwqsKITrql94CMGSc/cGq/Dhi
iTvhVdCjX+IibCnX8b+bk5s0whJCQBYqP/Mf9doGBGZ1IQ6HyXTXATUHdpg/V+kl
B9Xhh5j/9Va8WyGZTuHurarBcrJfMQ2hMbWxIOEzGCJwHmG+K91tin1MJEb4tfRb
8JHG4xs0BRfRCColDtLyL0H82h2S1d/SCTr13bpHYzmZePunw2b95Ph3inRqExL/
KXEmj3sFmbjUsoilDtOCQxtqWyHScQhcZftBhB+cAHL3y0wA4duINedhkbBugVQ4
ShHzI6e+4iiFn5JyiuSDQ4Ncjz8YL4gLOFekJb557lLNOhKZhNLtV3kOnapa/9rb
UUSbBXln7iMWmQWIYrs4NVbOlYBCnHItA6gcerFvqexGUA+YM6AgKk51GnkNzqKh
kXevMNLrIcR8DyQpyWiKMMQpBlE+zlsnlLF+Iam8Y//jzTIE+g9flc7AZtBpedJA
ZXxXbgdcPbUmMxEQL42gdEdgfPlzwYD1RdGovHS7+wm1hpXXVOjyECgebfjQAyjY
Vaf9zRxQnHo0HwUd4x/YcoUd/7Wplv9lN3f7j61jUD9BWetNWlu4pvM8FAJaUMKG
NmfD7eSy/GORSrctwP6e3SwGJDtVdlE5vimmN+DJbgn+gYJY9sTBFrWX6RZcS4Ul
TzVe8NC3GfkyAZESeiTfrcxeSofq9rnX4WReylOleCFCFF5aPIxX1sW6LKavIi/4
RdE+1FO+0vBD7p8wuQqdVAHZj3RtJpuIgrJe/ZcwN70NEsrsFm3n7XbeUS2lF7W0
ToUiyqgBEcpepTlfRtG7LaBZKpldVS3+OCxPpQqmioz1oX1CV1BZd7lwttppT2DY
PPQEGBQv48CuMxbxhrfu34G6t4ctwbNsReqj4NHfOK5WHbed9sb5kG+2paVo3iyZ
5FAA3Kr0Lb/f4DdUYMoog76ZSCKaOa1qqsGA/qpwEdC08OylDkEEfvwJsWJ1S2ur
6oBN1GOJ1XkW+EnEbVr0xJa17aEoMrytmeM8DXLamWDp5KrCrFK/zW1CHQvHKEuO
xvp/smmuAa0fF2AA8ocmHuyk/1bdMpNIFJ0TBRAELuHJ0JwAtSlFYy75ecckQCL9
q4RQMQ38sy3HNCMK7M30hFeZ5Uj28FTtVqs4cqmM3mnoSNPrZRSlo+kPg+YPRN7O
Ex9ZaEy1W3plfiU7ZX5hieDm/fnhvfo+K6zxBlH+/aAjjoi/mWNIROv3eod+e7NA
BvMh830vvyB+bPxjVRJQk2Mjk4nb4kwuVXZzGawiVFeNnHHyGNGBkL7T/06afsYT
0lDSdhpvbt9FkMECRBXW//WLtnlmItxzYGElSwgyA9w2hXMFNUOv8UvF3SVEJ7Ax
khzt1GlqY8Z0XYvOQdU1GK1E+fAAWB905EekcFGfjBVUXT9kM+XrqTg2CUVIBpwc
lhqVG2+vdju22R2ovwd2BmjietflwAX+E16bcI+fhcaTpkuuUmzTWzOpAy3RCWzO
iqEq4D1uclQbZIiJ5x+Ibj+gCt/g+ZLL/KrHAU1QuFB/z1d1NHrS3oaGmZjV7R1G
ReXNhW7ngq7ZWVKNE6Nn6+vCeu7tDnUFS3fWlRD01q695ZouBtYMn3czSHDSXVR1
r4creK0lAqMAvWFaRBPI4wI/L/RxfUtmvtpUFRsNInn+HQCYq+vFE7p3AN4jyXzM
yc4cWxmfjeglSU92aEoyl3oUYKNZSaKshwK9pz/r6+VvhFBBnrgkkAM+0k/bTDIV
5MAOUiLffdXj4YVvbVRKPjOAnMaYVlruBR0Mc/ffrcgxY92E9Go92NViQ6Q+RCZY
xZyZJphbYJ2M4McIItJaPioq36rHFfCLzi1qVt0jH58fciDYR7h8wG0FjL5X1q8u
yF6UGMrK6iHp9tTXD27TWfibz5HLiI7n0lADx3jh6Xj/YabZctpWcRcJgrVbZPTZ
djIJajyrrvnRv+l7gqXUPYOlB9r1Jm/MKJzl0tmh1P/P9O18KU+3ZwOUHfq/25VN
26yDRCSNpO9SZnoKd/LLR9YglwG5ukNkC9DQRILollyf5LE0+p65ohl1XoViv4fg
0jiircMyylwXYu5P9GucMaT5CSrUt5CjDdC1Mk7nQpRcJSvY8bR5rMAh17kIdi6T
OUOmQk0TyC3ML2fOsHtARBT9QRiDIiENhnnlbZr8lzlNteEND78obda6NPJmeOdX
/v7NqtVFeF0rX+ZhoCiyDcRBg+6fNDtmyCIzaGmOp8Xq3qW0imqR2lhsa8iCQmL0
INmpiU9iW0Eu1PEJQUW+VL+vQDY84cAKfO6PhE9LAEFHCihbJvRhzxVhhBiwJrua
xlwvwXQK9y6b6OKFdsH24GSGBXE4UbLWcjEkA8kYExRI8DWDdTpZmdIxzg33uBAY
nrBOkBe9tegkCOGeX5vyYxDsfkWmUICAGVCfjOVKdKdM9V4oJJPQuQpVgrNNQLnG
LxiGcgfd6qcnVGbdoVIhQgbJqucGWnxOFFzue1hqNW2MIWv7iaBYlg6z2cnG9l9z
OdysmWrmrezQvN03xVIQFbHd0+zZGsBinAFtDgzf7OtMeHX16Am0uTZAWtSS+8Xa
99BiV4sZVwTDSs7ofNKMpvVmLa4pUIi6qoJX7rCm298FVFqqOGVKYKwV78nuyGB3
uWjxMSSFE+RW98yoGZyo4ybBhERt5pRSeSMX/zfQsWjovJn3XOMjiDZkdM+ARXsf
XKYsDVt2UTS3LgJDnvcAjwl2pA1ca5eQH/wsXXS/PMetFy65xkEufegdnmkScBue
UwCaDfgT8zJKf2brRTGxbUksVB/mWtPb7hT6uOYbjCvvD6xuTkioyH5DtPSPOJo2
SMfAl3EkxYgQHaUatNFIF8V833ZEGTRav8o2PTSqLG2FRmbjtFvM63Whl7s2Ylh+
yNgCrCqaW4XGvLqbmSYcfxZN0m0mmoTljDuqI5FhKXdbyHiumMcAsuWLrDzh0q26
/+mLKTfVmm3j9Vff8pCvJ+Evdifkose1YfkLW1GTysvqyEzeLl9J0+ZHlMByJJ0q
OWBR6r+5xlXdKZWNWwW8Q+9x0JuX3pSaV5KmH7UlvZgwlxfC9nUy037nemWErbb3
da83eZ4D65kEQB76msXxM51ppOwpJcSNn/jTaxNyspXFjXg1u1z12RSOITYhhOVQ
wa+YTffYmYMdrfXgXJANUa95uy4sJVznTJNmW0j6kVvgraZ3qP/b4n7KuED3v1sQ
a/4Z2sGRIkmt6V8UiXK4ufO3RO4n5SBDdCSIcqiSReuwDUZ05Fuk8ELf28sC6V3J
Zga7ipAvDP76IgdOWJwiXpKuog6GLCN3/Hf5T5af6BbFE98vzcJfVZVjy43M9KkP
1FZlRCfH+UhbY8suAMxDynPuxnPw76Efc7YFu4CZPL3wtEv5t3jVxMDp1PrFaJI3
rCQOuuzBCf1a4XgVB6XLrxFm9iB8nA3trQiGLxfDhRwOWL//cGGYF5S60p22AJgG
MCIRIYJf/XLZKycpwkX7YrxM/jLfmOZ3LImr20ZA5UHB0RkKItxPy7uZrmyuwFg4
o/PslFWseqLZ9XcfdQinSFVQ/GK4/OUSr81nmyx/CIHGG6qVKh32tYx/pPYuFDaH
HXnDnwWq1UVuoFkV1hxzIxCYc7WSwJ+mGojRTvQMLajMVCAQh3GxOIFN5PiasM/F
ZSyoAYLEL3z7rCTXN90Dejy1NtgQXfM/7zv+AQcVNAuGKnwHk+Qmqi/tD4rz21JX
3V0iRIqbmEuWUny1TvIrF7gBjxyc2HnzxlcWRq+fYPF3GcpAG1s4sXZBuI5rW9pm
CHkVNZK+2KwJBJWwwIjwrRJmhobNbzZPMCaHK+OKAzrck5PVmy7Sqx2TLeRXLADu
o92dqAPLREQRay0Hfuvma9+Nd0Tbs6wuH3O0d2k8I9RysYYDgqKKdQTd4/7EZfZV
u3cNc/cGnFzHtwU0Uh9RyvrJj0WDeCEzYMuaHxnhm1hQfnLDrfpvp/8jKUNkU9EJ
DVem86ic6gpRvqDcQRbs4+1neGtsFj5sJBgqsGCkKAUL5w49uqHl3PPleol1NEBa
P9WMRACKEXRvvQ9IoQiWCcRavz6JIFOsgMJ7+B4fu80gvVhzK19whJ8sFfdVPDwl
cozKjaaZD/6u6HmERSySzVDE9v3l5R0UMw6PBpOpAsvTw0qh674/NIB1eGxWEEQw
OsQ4NDIw6rR72ZYTDdCBYW+9EOh4zR+YNkhE9xsCmZfYkK9NXgg6lAbotiufUl+h
V9Q7LoSd5rbM8PFVeCA3CQErmVh4+FmrCPQjF5Rd5zWePebCz1iio7VRo+voxM+u
LdZ2OVjg2Ko7L01BVC4qiHYeoVffI6sLd2b6dcGL38yIyzjum/6HpFOpW9gEEjS9
MzIt1XbytmYRvPIP40Ez2hGHoWG6fbSnHAkjumjpGNlncZrgFXa9BKgZCk5BfGTJ
fGg++ylUBP8ddURKeCYhYrB9YRtv3OLXZbkymxzOWIt1wCbhB03qsS1yif1NjGXL
Ipxvsz1HkWOVeT95ztAgxzYY17fFZURHFAalHs/KlVGKxE6u47dW1uSd/gPNTDAm
Xi7cs7g491TpxRxcdORoVuhg7X1l7uSr8Zfiw89b8/xEn7wrcbZ6ANRgI8/LgNQO
AEt304ydp8xG0StQEzpf/tMqbB+nCYqBkc98vkJGbQzKl6rwbJmprQS9D9RZ8S8V
ReKXqmwxIvInQzNc+AgsX4ZB9zD2a11un+WIfoSiJd7Vsi5wm1GMVa+NuKR8Nb3b
lgRYB9mPFwLwtMMdbeCx7IGLZz0agy6hQ9jgeVrdgcz67ymFPakqAtjU5D4oSLjp
oqBDu6n+C3n/BuLrGq4jjqlXjh+ZA6QLIyh+g7MzviIuQCPO3CsbJ/m7JOcJ2Diu
TqZZP9THrYK7roM/87w3ToHiw0nHZsT0A76kjEDVMjUuiNp1pfIn9MYkkiUWkn2A
+ieccf+kRGIi26DxUrUagvet6k3fBiJWdYQNz5g/WTSBCkeDqwyfw43Oly/MUETL
5xxMXslW9GEmPQSWLOkoTjzrchyJLFBDa55V0aykXTx6Vny22szfpme4pF5BVzZu
alxpQyK9hBdrp8UJMXeWOGdWo00xYitIXlnryzbLwOeZLE+XSGs2p6PCr5wwAsOe
ehg1n90XmVVjLrquAR3CymPzR/Q1i3XaBa09qjCRmhYrh/3jvEPS1NTB0ywVhWzk
EO5KRdh8GJMWSpSWW6a5GUc2QwFD9qmpyWnkolrbP/WA34yzlizQ+j/0cw6tr8k/
9bQ4IDTGcPQdDrpqDXL9YAz3xs4acATFRGHUG0Putkke53wKSBoUJsNCe2/YkMP+
eqCAVjxfQjlKGsdVmaVu0Jlo6iAzsmSOY5zT2UAjO0jzBUAy1WanFau4ojxFps30
P8a/OQMA/y9yutmi1pV9K8baWJeO1Cg2irNWK7CjieSzcFg9o8OQ4TB3Xv05+F0O
ltRRK9sIU1HcVdQIy9ntSshu0ZvgjonmOHu0vBaSC/J1oIdpLIY2aQ7I4DOSlg3Z
GcWea2MGTJp0T/Ld1gD4QqLa+aU/MhMtG585DhU8/esZ2QCRyFnAxhEnMrz22KjE
lpaFCRdxLD+Uhia9vs/RQOq9StkWNe6AEPKPHMXJt1VS2zmM/XEiEqUNdvu/vYG0
klSZHS7+8LeAXKNVvEhVoNZRrcohRT4rdXsNG4mWtA4ndb6qpyIm0BzpOqYdWAqq
b2568Jeaga1sEikjkAQ39XRLCG13VH4bdi6JUdqTeab8W0aJ4MKiquiCTZprq/2g
Vp5z3ocB7tS9R2posi4jTqNfZBnFgCcNiCG987mtMZ20PA9lOD3qWMfp22krVUNu
GhHi3m5MmPT1US2SvSTL1vP7SW1vVu/3LLkQXSh51jt92klLf04na/piBXykZ/Ml
F9QW3EzsQY17xq+Aed7BdCYbUs+HkL12CklQy3M+eS4etjrsENLtbL62ar/2adhg
3Dg0+ZqNJR2tCQ2kj29RKChOJ+W/MCZLfHuFXl4MyyNo6SoBIbGnfKcUka9s1yZa
Qv79ILC4KB7fRmMkbqWLYeBc6qZV25OlWSK4jyZXpgUDEKWCQqfWzC4iAsXpJ6dF
gQ7WXaIooJwwu1+6B+JDEtN64KWXX++VCD7gLktJgTRcT0S8f+7Wgllfs3EYyMcB
qsUwK+/ku7BuK4dtlaUgUPczbKhmtN8Gf8nl0q9ykmwNR64f0Xs4X+qIpKsaZRrr
eD/Reg9fxQHWI4v3LIoO6HOJF84SfLNi6YqXUcYGwx6xUmV0Q22T92n2HnL8PUE5
0eceq+L2QSbfDkYIMkdA7XK8Zzcm2iSM1ICwl/Surri/czJ6cFjNcxYBWPVoHlDO
Y3xsm/cFPWW/f/r2LAPOU7lUuwv6oUmVkd6BDVwicjgowiTGOFWv7mwyM581kzsC
4N8vjPP8DrmHprTWuzO/fxQPHvgOr+GOjBHUjoXrzfYFQ0AAtxzmjuHGkAAGwcoB
4+k893yoK3coB/UoXX/6qnKK4LPTkcjWW28fhz8HizTU8vSpj3KGNlI9p7SRzMuL
6NxvqDf8HJnXuYiJAh3nDJU+P3GHdgGCquutCOHvt2BpO5B0dRuSLZmES5IIc/N/
fWoPivQMN/oI+l4yV0MZ0emmQciUV+Q5WsoAaYcnF2cPZtksbP9w+GYIYxsgadDu
hHAi0CMPoS5TAJc809/3r1vCLWcu460vlMI5Z5Lza4WZQQyxh1KyoXuYFjbjvccM
J+mPr9NhppgM5pfdrMiNhDJTrIl/9hwIjN0lumGQks8RTNJu4YAFjI02nnHx39C8
OUoC8gaJ0ChlOXa1Vrud6m00FoOzo5g++Yh9CQD6MiS/JXNKTjHFqioEE38YtW5k
uJZWho/DY3MPJlb8Ve48dX9V6DXVCWugOYjiEwrbD+CJIoplYyQgkuYERaaCVXEP
B319UMNvU0Wk/Z7yMfZZp9/D0Os9mPdT1ByRVEiyxvHq/Mk5sL5i2ofsyWTUs3q1
Z9Jsq7OPauhCG6ALGRL0rey720FGhknCxmYWbsDhGdG2rzYH6GvHLcQoWodsG7Tu
n3bT3kmsUl3Apnyy1ioSRWjHlUdsofTUZm6JEEkZPWk9PcCyFIi1vGZnXS0+TOOt
m8/SYxOylqji7segvtB6lz3yEaAnO7pnHyFn9iqEToqyhMhmWl0kadKdlWRpgr9c
7j/Aqmk6ytzsvA5vcdOM3WaSKHPNQXrTg7H/EiC1Ijk1rGYZgFATZs7LknSunc8E
NdqaiWAsV3Kvbv/Is259shx8n6G03j7nWGC1Fi0wFGIBfhIrfIB2eqGiqnihcoUd
PUlkbXMHCo+tPrJ7qPIjiDAMvy97KjcrUyvnAqgGbXvKS0hi4QnQfZNCMpbjGaX5
cyr9KJVShRBbXqahHlMRuqmRxZbr1tiR9PGxgOaLkOgYnE3POnPGEaswot8v2Bt0
IIfPLPb+ImmJ4voFT/OmAOzaiL6t5l3c3mHLIlxq7lKhRJusqcKs+z7v/R1RamvW
tA/2gof/sa2Uy1zy9ZznHIWvcRIVwno42ojVFyRCSI82VXT+twskeg5cy8PRiAk1
785qt7MUs3qlxTnmDESdoBeDYzY3in5ZJGKGgU4L6vvnDEHo3ui75MLjwLKlzC2F
uFwoWCuotiq5qUeDQvf3IlwqGBq023Es2b9OS3z5hPKy3VR8KibeZVQwPJYvWRIH
OotHxM2ibz/hmRqSnxI/p2V4o5TEfxZz8sTRUHWPY7/D0A2BRC34Np0t7QT6pKcP
AwqOiKQarsLqYX+FWPSa36W5mK/Bb6KkgcBiE0LhOpBHb/uZeuxJ7mP5s+grTwTx
5n+DernOLPPpx21Lv4xb4YKBXMZJMIsHRhYPqiidgpYRwtI0DBsg1fqHbBPnm5EH
321vCbMLoRkcWIriyuGTEPQOEJve0lc9Ot4wLeI453lD1e2lDKFoXMAR1FAE4T20
TN9a+/KJMryClKh4aeKEFtOcHarHWhEeAIfApOcQq4IY82tnxK9CmmJJiEjVwS2j
arNrL46AlwdZfoku02bZp3O3xCsbN8dqCi45dneXs5Mh+WJU4lWR5tdmmJihIpjo
hNuK21DPdzEdYm/08oEnDoEmEzdOPZop0xOA+D+Ha9JXx3RodZYtDLJ9xuWao1y3
ehqTTSLa7ehfQw3IvzwdG//AQEgbiZKbdGWg1pE8GU0VKb2I67JYY0cwQVlCnSZa
tK9m+rEo64/zo9E06dQdsSPiL0pt34Ll0bXggGyIx0S3StHw5/ii6dvY1imCYArF
SA9TeuZFe1sGCR1PvlEd6b4X0AYQKgqOp+s46EshjOLCx6Ie8L3+GViXKTJ1ZC7i
2MJB/69vtMXZ085Nmhskjy8C5prRKmBozlLsxt2IhQKl3/6vQ9NhIbTg8imFLZif
DEuM1ufGb10pOrYF85GTzBd2GRhBAuXx4xTcN2+tbEDSPhAZIitussmPDVAcgLwT
v/CtDxsAGeXzKGNMFtuQB26VcHnK/Hyz0J1bOkRhA1ueDj+EtNRJkKilXJwpZTIP
WaEVWMvdWlMzo299n22pBm/wUSYOOJzFFFM8fw2jQELoHuQ6LvJowzMlXscqiPPe
tCQ58Wgth8ispOZpQZxQ8eEccxCAJNESnGj+xWp1lUWVjWiaZHRsEIsjGMM0AeNJ
uPH7ojtgHLzj3nt9b413Xoo8fKCUQ7GYE1KkD1+vq/yw3uXgxs4aBLtKzV9K4bBF
8Ry3I5/J/5BcRbZxjeo6fLcm92WcyxFeSzq8IW4fbq8Vb/JJ6VXQ5sOUe8dbJm9a
oPnL/HR4iI+3swteQ8vrdzuSyT/WgxjLlbKTC1D8h+qfJZMHn63pJj6KUjRFs8ei
MrFNa1XLoN+gOdG9WauFedXEcSMqPIyPBuuQKWIltBTEjr9sSoanLv2rpCKw16iL
gLUUFRV3q2XOWpcWzANtq7oU6/WSvSeaWh/EL/pGKbh3v/WfTaikpc2OttIpFSOC
TYpEqaRtKGU/cWNvyY2QjjKFcjJ142oBuNAXT6ncfYoUVsadZiWgGzpbOeLLbSaL
ZcWG3jDjZnM/Is0Ql167aP/+HJ4b5SV1SCXjPFE7/LlfeOvAthJtdDWeK3DbrIbD
ezoz3taaFSuF8EveT6/gD4B0DOz6Usj5bGOn9W/IwLCYVo/JfzhpLGmrXauhqlUj
16RrXidKIQJni9GEZGFxL1I6HJytxcayJy3vXWb/Pz0iLA3Ej3H0Wc8VXXytSAGw
DGGoXBb+Z2Xj5pNxCq1LGPQM1NeceuxkHIqPXCa6PiG8LQx2LQK37UyLtoFgp8Ji
3z7QfP8XvOJL6L3gtFaJqjJuKcg4oLTRLXAIPJ7uPnwALCx0zvuLjgYqxYEPWQIm
6rKZFUdIuusIpMg7hdK4+yKIwxlsKFet15056gJK41mL9KN+Pq39NvbIUgArVs6M
TnPIo8OSXCMi9eYeq4Hp1/0AVXfleVomuKYU/g9SXl28MzQkzDSUv6dfFEW/CDnM
RKFB+A9jDGafEG+PJ0KQYykI6N0Mri/3I0H1TmkPUWdopbhJIygn0v9Gsw9zwDdX
Zr9xOJQ4yQ6WtKqqbXES3K2m2inlZR9KD+1QAVFjkD6HZgWVPZxBezY5FyenvlRu
DyL3iN2IiHH8h4lg95q/IkFIw/I3gVOc5HMKhxg/9LgW2r+/EnyO68H/+prri5uT
1pW5unxn6BnYMKXPffh6esZeIfQRz5Bxft0haabRbC4IKfbmM2r1zbIs8ILK02n6
Zacn5mfV+i1xTRMTSoAu0CM8fPAX9rPsm86SPvdTkfwWlWMC0GnrRH8IAMJxf4xu
7rv1DCHGGDnc85b47obqViPRfxCN5AStScc+POLpxzLJ5+iyoPZ4mmd9yQ2nP1PU
kRKyEIOdwGkHaftzl9axpDSOaH2wztr57E+n7iV2D5Iz9EXfNYa+r+6/RP/icNGh
BLVFGir8vnqbF2dOOp4EhKnLwPRcRdCzVZuUFkzDxEqCrH5gcHC8QjSszeCY5JkA
+qBZqF4LfUlBUB9UOD+ltFyu6w0y2hLFSC7dXdSS8/UtocXSYJ0daGn56Pw0xX2X
LjctbHPYomCJcZKI/50hiTSzxSg3B8MuJUj2vr1q6Cfx5e4W0XoWFC1bkI5T203v
jkjbXgJJphg4OUStPARWOjaF/qvE6RfL50Urx4wyVcX0y1NFCBbeCpS9Ax5ic52T
bsZM54SnO0n/mv2RjYJRGgyhBNG/+90XZ6Wyl+6X/VfPvz/f2RI/pG6fz5mkGaHt
HcKnnmQq5rMwi4boC+WIs7OO5iuZGwkNArQYIy0LSJzUYeqRzEBLDyi0U0NGvBvM
FAXLr4r4kMqALbj+dRPp0zi9n5TeRZwTU4bCaCk998zZa/xcwbTYCMqfHgYpa6d5
PPJSYBptNIiCW3BLBgEr1mDA78703toq4u6RikCkoHrZFiwiFZZ55MhEoZO4TTZ8
8Xeej8NXXwoqrXAnNH5eHhg5muRCl+o6mdKnlhjAaaNIECQu10Gh/5ztklEAffco
VC5HSIE+qiONnYWk9GAtJUrA6OG1tjorGBYaZ4nt9RRVdeetdF6mQIXlEsENR5BX
lYyMpCd2E/RjXwpENJC6B1JVNWEzwz/6uFsPYFQiPBhwhMHVy+4hp1Vq0tJMp1lO
8FldY4ea2H7l9kNf0xGByEL+GT0mDOWKtJ9XJOXrB+b2tGEXhNwHiqee2XuPkelP
TzJjUld+kWU5ytHe+T5o+q8b2nYc6F0WSACyxBc/7omJxn+0Wz+rE3YbzRKmY6AB
kY0pD7gmBIiCiiFO2bWrypIm/uT22hU7fE0HL48SVgMb8KcncitnjC4F2M/coWHW
+7UA/f2RaD/BIDv2maXlFJBeVllXuDoJQnEZ0owCXGlYua48XFx21BAGTDOk6QvC
MEYPe9oSHnf6TYLXY9HPWswcHPhvF+RDvGDNo6VgoOrqtaQUtjJjYzR8/bmyvf4l
3Wo+SU7QTg+tcxGMjxT+RlBWP+8lBFUDqV5Ru2UX4fRaUwaoURzLyykosIRsXSLZ
MV+pOzGue04C+SIPL7gUxOFbqhUVhUquSLXmNk+0hzlMgda7SLyr1q86XQ881GTh
pYRngPQ4B5AQyOYo/JW4xPjrP7RfK0ZgOqKmmwOvJLunnrj+vjMROzH3bbAX0RwQ
0rRL0iTRSoJ1WbOrHrfNPjmFJ+WrTHniZEFqwkUc70INbj3ZN5AH8UJVK7XhxGW4
GTq4HopaKZYwC5CdwexdurBw45oV+eD7q9DSdIGoyf+Xv58Wls+Rq1Mj04cOgamn
5I14CWjG8UoZS/F7OwlwbywN57SU22pC+lJCr2PYMa8fr7BVoEDom1WEYK5i1/SM
ZN9AHrbTxLubnZcVufRR00XJOdOssA9BUC4mCO+g+eWkMw5abmuxEjrP4X3CSFOR
NcH1wQneIJmw3RcbWOAlKs+B/1XuuENU+sJxdLXtJOv4tG+nBe428pzotqX+9Mni
te/uuNjD/RPBjFuPnjyundL6khIfGaiC+ODqL4o/4k4Hekwi1lSZV1f/maHb531c
D3m/HUz3ZqD1c35KmeE0UUJk+sTv9BVh6JFUoH+rWf59Dynz9Q4lZn95b+gjY+v9
JtJQpXHLM14kRmeITfZB6/4Ya3aphEDy6Eeyv+OscRTvHBjYZCH1+9r4ktVwCpde
FnwaZV5GH2pwdaFvhzKz83CR0E5ax9K6jr1yvfnWhYidLyLSi6EIiF+tMJXnhN0M
pPhNxNOCHHg7mpkCsnp5wkA34/5EKBdTdl5WM9Xawz9Etz6rNcd6vU+6k0m0I5k8
A1LmKVty8ak+xJTd4I0e61vk+KOcY9GAbJqo5hHisbqcLgPtmkL7wLrZQpwZdY7U
i4bk4Kvscoz8wxBi1goirGd6+hR1VvZMXTxgqv3HCqVDv+f0pbj3SVD9YitgBFd1
iMiJPHoa+ujmIU9gnZoKY21bpiMmCIpybwIqT6pQTGkQo5TMQRiEfW7FGukDUYXq
oxHRJxolz0Gkffessty+lhch6h79vNNdCuIi/qkEYDe1Vlkma68GVG2kakAvYPXs
heEYTgHQfkn9Jrm2mRY2zvmcsRj1+F9K+wrkU1z06+uGEQr4yAnmESoEWYNU+f+B
WE3di7paLieXM/2Tp2LFG0r3qmAgSDPIboEtdlNspOrakjDfSBVmaDkDuOZZACZM
xw25g7lnVzmCHtMdP548avea0pWCyLePb8W1RGlTLjkw/0rlAUzkmFfj2+X8QGZD
o6QdG8ZBLtqCefw+U2z/lE3T5ANv3a4NVshqVGEE+/W8OgEus2ir9X87qAk/4suP
+160nkvSb/GYebX5ngf+s5IufV8aMLITOcuJs6i4GystaDv05zOCb4kmgnCaA97b
Kc5jCYq8W6FILDcbebXOfjL9lz3oIqhxwF7bm+ziK/rMbvhwYrBn4irWjkz5Q/FA
lWPBYfl+i2meurOdwKgsF4390fSE9UMO0uMFxkIeg5/F66n7WpDEqextCS632PXu
1t5512LKQO4iMgmS1zv64LgRR03+99+9yvmXNMeBpZTb3PXnlSzslDRsJ33cJYXk
j5rxZBCoGCgmiHEjklvScGQgG1M/c2RO4gVZTkZHsRJORZsmyoJk7kL/rC2b0mJW
neytAjxO8vH3uEFUUC+x17+KCrNq9QeZs3tSOXiErWd3tFBXito52hGrBmTBhc2a
0svDAc3Fb6vETwRMbl0AMG3v0FUGyoer+ZuyN/W09zCno1FNm5fUA8Sv4PEfgeqV
8o5hDvCpTQo8JynfWrlldDdwk+AmHVEWS9lkXZkmmn5e14hwDnTRyWTs25j1trYF
EUfWVliwKaA06YOeDX6NGIkOySFBT/b6lPajXVWwf53AZ9bR5Gz8XI7PuqSxjBBT
zpJPmiAYi2pzelmLEM0ESOTUC8vuXibg5qmJtZUaSPGomK5XKzFQb7w0UkiS9BJv
nlJ490iuRNedPiZTpgEJhxoA4ZDmKmzKuBm5yv9iY7W6NTdHHPg4zM69x+2dIEUo
uRcsp44U+t5yfNylOCONVefdTlmBpHbBD+dYnhi3ddmhCIu2n1fYpsPln4aC+Dgb
9w899GDCAspTx6ofC+Jmmi2A8m9EFkEcFSDUzqWM4LMQRgStxTKLPuVy8reh8pt1
izxLhp5pFV20RftFRxyocCEj/uEzeqN94a6A6VFHeHO0JgE+3e6xmVMC8wQP7EAl
FpRnX6nJWRXIUfgtMjXrAhJ8tKBqVk7OkytrN1FhsgEFuQ4gNxbg6L+1uFwbboMw
T032StY1sO4f0KJBzaCEpQ9xGTXwgJ++ij8FsOROm7p9s4vT1/Cqya9cEVMUvx97
4GZzcaprT/wTmMvTQtJyJ10egQ3xzHHUe2La2SveptvVRdppjoAAmsKx7tgCLNIU
wiO2UNtJZVj3BxlTclmv/Z5jrTxyfKLgZQneIRjfD+NyG3yb/KJ+VkfsgaEuYGpW
QxDITzcnuOZ2Bi90QwYfalEoZ02s+OjOMUD/4iBc+QZFwVrSHXRdk7itwOWsnoV8
q7++XO5F9keobEQV4eDWVeBaJbtpxND2w6GaOzaTWaJXgi9gNUfxnFSikwcgeYhp
nvL17CBUjt1tLCSF5ZqGQR7kST/t289Y9veuIHK13tMmA98LGBS6WJuDq1AHPuzl
mxyn5QRYbrIQrGPInwNlDB/0VyMbNwvn4BmD242qQOkji++lmbj+1ZPUJhsO11Bk
GyReiGIHaYXneVExF0wP0WYe+bAHy5sDCsnkXB+UFgkzmVNjC4lb2bSsEXE2M7Pq
6GPVUp0NnaD4JTHu4q8Qz+W9CYcc3TRRdqthYoFraiUrqbgDozTH29ID4oLELIKw
uFvswWTguEUTsLF74xczzo3N251EDOL+EBDfMFCQW2u0gkIG8FOvN7uui5boAv9j
yFG8JO2PYkBVNRwmEKsIuYXcYhjKGS6J5tAOxEKZgL+eMpYRlBVwrQMi7pjbaSHJ
0BOzMM+G8tO/S6vYvaLHp7si0C/b3QBhOHz8/wKZKcS+GA2c74DGdI6OvMcQVOvQ
jHA4i+5e9G3TUsRR9Xpfn8CkzfzAJAQ3WJ+6us1HTL7h6nyWjuM59K5U63C9df0G
+Dvw2/l3Mn+I733W7H6aus5CMEzXkCckgfYcMNcKLFd4Znx5sV/Y4Ic/0MjyPV/j
J8ihYQVjvoTohHNlop99yijjvb1wbNxTNXYOBW8yhKGxoI8wUHQyKmx5iQZ4tV0K
5ItgnhuNqWjYy3MEX8x1TwiKfadKs53ku1z/lWB2h569JIm2TCCB0jqtWFBd9vb0
S1Eaw6XMm6JeBl7HTSGqpxE7aFTCftK6DYKFc3PGmDxCSVF1hBRFn0GshOuWOuXO
wuFKmzLw0bo2M5Ga7hRCYOU9rmnpcyNBg8X7J0ZC6/aOGVhsBQXQ9O3TqX+MQaUy
mJCmYOW0IZdWTOaB092bZihNCOP76kEHPQm9Zv72O/kPRF9eljw267zsVsRWCp4v
04iaAxrjhKdo/R2XGdUDd2/8WIaQGag66UaI7s4VuF9BxsLmAhlfTXUaEoemQZDe
WF62DFE1+8TsApw3Da5U/qnH31BJfq/VWjSOvPLLUh5pthxhFvP5A4Vzl6bxjT6w
Alp6JNjA00AGB/aYa5qeUrC+5N97pMQItQjWSyaUYKiImWHSCZcWV9bKXWOaE6va
TJl2KYGe7ap6AQOie9BcM1xYolxYr8f6C5U7bFQXBcfidVLn60ukxL+tgv+XzWRI
oEPs8evN71cSbokbzqPKRHKEwrvpYqewTzfShVhxwVkCexSPIzV97YDZnpjPWreZ
wLZAqxisR162WRqyeQTmfFccfkKRQH/YJs1bliqeaACgo+oilY/OQKzUrbZl0c5z
8fTk58F366I5edjNAn/jwNC6oySezUUBFPkPky93qnoS43HhgYOCxeg6F30eIU7x
R2+2dXxx+m4zbf7pVOty1A/PVX/O46Kq5tnR6PIS3vgwTHtoiEo6u9mK+TqjdpCJ
djyUogNjYAMYHdEZbPE92dfTE3l/mlIAeh8lmwJ9Y1ePoVH+plj6Oug/I9cI1iwT
A0GYb34FT6By1pipjVTp882dHlmZ9kK+tt8RQmd+K4S4QUKxEZuhJTYv6Q1G3VLQ
oVK2Dd4VSEsbfliUGi8Uosc3XTfHgfoFMvM57VCXlbt0ZVZkCgrEIzHPNB/YvGcQ
vP0wni1XQf3pFlY/8HqFyBbfFKwU3WJmKopVrIoIxV7vucjpGd7fUQWOaHJVXnsy
SMjI/qR09exgFsFqTceYQiEluP8LoBLxb5Dz9kf82qv4/6b64Hxc4yYJYBtYc0td
OCp1x2z3cdWXSh/DYV4olZfGW31OQL23CGhiogKfTEcFlL7kr21d/t/P2wzeJ8Zn
ZNXDW5fM91Ie6GL+oemcE7M8OVD9KGdaU6fPJZuDiKSMFAvUghBIyfPu+orRTHeR
bamgdbo9YqIZmSV4z4vXlZADE/HYOty3ZLKfokQ1bOXajRh7dyP89boAn4JGQ5FZ
gMU1OsgFK3xHLVw5Hur6DEJncHMh6LQbpUOuShoREUJuLSGD6+DahH2MTejLyBzT
JOeCvLGADWSXTIMYM/51fpnoMk4BnixvHQLhRZBHeF1pDhPaectKmBpV8WuIQjUq
584oUxUAnnjMoLHD2Ne258mEBGr7SBwPe5pTtcdl658u9E8gM050URqqztzIUhV9
iEykNm5FVALwKkM6btLnscaWQLRZtN7uXNOAOtesuwWyErYDiISenr7YF8sOQiH5
nn1vDXqNXx9sJ16jDUNt1GI/aUDmIFqeN8GS2CbxzdmL+Gnb1BfaqVWg7BNHtUeJ
Rv4lPmbkAeP8cgca0gRoRdgmJeoAXW9PoYFYeHB1/BGSQcAKe5GJZisky+Tl+Mal
Cy6fExQvxANYhCxmHtnrcdYYmS/WbW50v0Cn4VirldiYu/7+WcUyy043cPhTRArE
QD9wm7MBAIh9juFct4SlummVOQIJ3M9XgqWD/0/nUzBrUQx99Dh+TdpmVY9lvn6O
9jWvraUwFMz1YetYL+6V/NyJVZQNADzsc+qTifqXqEVmoDyy91mzv6oYshdT/ai2
706/qt7u2BNAJsWDJ2EUQbDOVmeXdxJjnXamoZ1GJA2lAce7w+Qzw1M84u2EiS1q
A2QONU6HcYZxddserlk2d0wm2Rzhk0HyV8gtokTQeznVpqiavRpte4r5kS3Lmd5U
RKdCBj1h0k45dmT9uaz4YLnNvD19PntbTygFLgeY5FsobGPVCRFSKSCqhfX3iIOL
oNA5N1GYfPkf1lhRiS5TS72WHUZShDL/6pSibeiKxLb96vHFDQE8nI3k61go48RQ
qn3uCVkajHXx/CzBnu+omkPp/1HkskFwY++RK/XKjtHMwk+6N8R3chuO3tPYhgpb
U3VB+gKjja5BgPgJcOQw9uaPJSFxZ2iMlFzRhcHKEQnbnN87g4B4e2iFFsVHI5L1
4FaSVv/wh6YQsjt2+dLB7xXcdkX8Sldi6UBq7SPXnqNzrBl1EaLdyfMFuBwuJnpE
fSjAah8+jWqboNOdMucYxzIYichOlflAXsDxcD2aMyGtFSs5QBLDx1sW+FUBvY1L
BSmPOnrm9QRt7KU6LImJhcFRKe2FF9y+r3XCXbsQMoRiuBGRL5u46bFXfddQhpaZ
EgMpaSxVcVm4AXrBdd7f763Pwj5HR+Mgw8fX/PDXrapTFoLst1KkvnVV3FDcJ8az
B8X6BSpb0jbbjjrEJhdoQ1HqHG20AVkgMbXqhyFjl32jiafQK8xQb7tq+PCyziqm
jK6LGwZAGzVJ0oAOgUDshzsOBCgSw/0aQSnm4N2A2sEvkJXUfituSTv76JoakXSe
Ap09lOsZ492KddE6gaiwL3c3cg7dPqQuXoq32WNTVD10qduGCY06FmXNvbfqfPyz
TJpGx5psNs6G7EMz+fU+nXAVVIcS/cqpR7lwziH7eSqmmsFeJNO1uB3K+IbJhi8B
XrnzzwCYghJSgbnUA7pq9NXQWTBKdjnBesm15bPPYJ/N95NkYFEpYIq4zk0lBqPD
VLhHdX8/7rquEoSXCyd3a27IVzi1McQfeSxQ/wd80Ij2zt4cYnys16GZyFZ52E7v
uoHs85GlgEqw00OL+RlapGq4iRj4zQn32mwwuQysW2FgukIfx5iX63TLnDarFqgY
F0fL84DfSgoh/eZzZgyQxEInUIIad79Q4O/AaD/gwgHt7oZT8+a9bTzqfFlSM4eq
f1guNv/8l4WdRum+x47BxNN4u5n9YAH7Pq/fZIOcOOPJ1fMHPUsyRMgdEcpnT8fa
NQQfGfjn7+vUWgqD96QvGG4HLPUGyOilGVTaaeqhbVaRrSWuGLxB1PfORMcbzoQV
a7peH6YvJ34F42lLnvLf2HiV+K+nI17qOiMAEGD7C+heSdpxfD7oB8Mc8G6LdWeP
FTJhnbiYW96MTmENsKK+zthur/yWH3p8vavYN8vbcxPwCnJpVsdz3Gcc2+bh/s0G
M2L2dKHIPzhpSClRQj6oQ9fYGG9xkLGdyp5EpN/aT5wqcbgK/+pgh2WzJICxoP1B
sWiR9+MrvnI+RO5YfDck8iFahCb2AsD5Kv8i7Kk8qDvGcQ/heaAqSEtrYEpJF8BV
7Bi1OelTJpNA0BZudNd+4csoLR9f9YxQC1DtbqfL6a0/OWW9KNVBWgdTDgh2wo9R
mwjBvzP3fvNPJYTwBWWim32wmPe6NKSfJO/Xq8lwPOiCtfQkI1+/oiLYSVM1RhRW
O8Ru4pmHSLkmY+kEWOfDFiL+O8E1pGkTUT4luwRnyxkWUrZA8sBYmecKWE2nEAqw
yBkdTl9nNTRtSUBRIyYUzqUc4wm7PzDJEDjFOwZ/QsS25stygeGDIRQql3hqllCW
dCb82lXkUtYAeJLNbNGlVyylsiIcQ0NEbhCerT9WCDQvhSKhbxCMY7OEwx3oTcHn
qrs3xg8sZ6O4bitfCkK64H2pxd+OEDNgWwoc3iBq7vWiMEsHb0OOm0oBoxaKyFJn
mEQuQTVkiYbJlG4mluTTRIWd97REFV12ItBRw5zNhkMyz7uggIBAuxz/jfJWnB3G
Rk+ffSAB2AEfR8sD80IUZlI3vFGb8gvDV6inGhhO/wqP4E12NljTBVQ9mxCQHjNS
8KnrPSQOUksv9tDnsCpCqo120qj2piKfMgBGIKOjpqRlOGnbGwk5NmcSTh5z8cse
/a3xGC8rApRDILpGwbMhOILJgWsFsf5f07BdU7eLVu7x3OIS3vySKfOJn66uVI+n
/ZLiiWKAARZC/nvY2wI8x1w+nGmDBNRkG//V7vVLvEWZDCSLopVtMaMQHIEo2iZV
8BsZ4NUAIBKDL50V+9a/mw6C7zeA8VBHlDi1vS/xm/1L9NU2qSlgZUK5SIJ06Zrq
pYUeT0X3AqdAav7lec+mZH5s81YRvXVRt5J9aBVHjXZRXKZVK1zWPNIfZOZiyWN3
tmRcWDhvko+QDV8HRQzruO0sHmsbMtYc0NQdQCwB7ErBaiMs3YPjDOso6lzRCzmU
+s/CX498WHuOphjdNSTSzBHgfJqR7dqlfsGoFi+dSa+2g83s14/PBufRig5QhOJR
/aNccAq/OzFxppIf95N/vBJ7EExchOkZFatLLGkp9oPBH0+7ziYNwcIz8iEEES0Y
txTT5qkR5n1CNlU6NsrILFa8q2CkvRfeGldCIpsMbVGGM/xmuKR24vEu1jIF2OfW
542sJDhku6DFIJmsgIxUaXdmL2wi+x1Id4lbbbgpnDPJhslxpjH2ry69/+0rwcfc
R+6TtB+MQgqhL2VQmBfI/CWP9Um5Ifp0UxR/j+CPrE6vqbe9kGzMPk3FlaWkLkJb
ITSLHbmHQZZ0vNmprq69e1r4HxE+RtVmnCcp5Y9OX4v4oq0/7Pj1CQdLNLcv/5QM
Nkoj7bXuZ+bSU2CfEo3aup4MLak/LsurfiuT4hTiQgrvpo+l/uEmjc079Oy5A457
827q5vG9e1d/dEGriSB7mPx2mBMrlnnUGKEvR2ktDguwBCBEghq6+N6M8++0d/I7
vHuknB5ItYWttR5rxkOi+yD09AUcia/PKCLPvRg8WmoTqIG56y0VnmwbybTblXgK
M+d8dEz/HWHZyfWA6sYdylRBA8/JuKcEEOr0R/7WnkMQvVm7G+dedjWLw98F6mz0
SrPjWwxpba9zeoFeLxG88I6t3vfn7fSxmTK2E8SWqXFUysicevG4BdyLsE0BFsWL
xfGKQ34OebIt/sFDsSfYznnb4hPcyBBLOP91eWDosZR9xgbIhNy6HCrGlRKuEDHt
+yMQhYn/L202kObx1hi4Wbfgih5icQhcATCavWvrXtFWhNmy/WiBgmQ0d35dOIhL
0AUep2GWdbTZIlYzWoLsfNhvE0myv0OtJ0aGmvdGovScMHDRzR1VBvqMHyA2L2vy
24OZIi1uFZcI8Gw0aBZl0DxhSdhBIFobUuAsLCcplbdEZwk6ZyXnQTAb8NREekiB
DVRwEbrbjTPyE2O4ampWxvolJtjG+Ku2rolEJZVqIm+eHgTv+N52z4sHR255ZcQ/
tiGz0+7F/dWORbzyHAo4QQLvJVqEOAoqkF3HlMs4Jl03ylDHuscXxgtvnCok6yiG
+OSp7FS8KicZyQ8XaGRIZAY3G//VHnGR7QwRa14RiYVdnLVMJ7anRybkzEksBvlV
D7/bgKsBJZMAEpyP2M37GGnAPoQ42xsCRB8mEl1WkQk2Ns295MiZOpkmyUOihNkD
CJwdSuaIyuxQPHqlYGPw31ZUta8INrbjQYqP9DITuz388oQqVIFKW7G3MydVeW0X
GVmFa0x54Xu+FowFGIRfWf2k2LjE69RqmCiFy3TAuhyIOsVNxPXOMEwW0CZlculk
YexJkcP06hY3k1ecu319BKiKw93AEUeaGasVJz/UDyIUR7Jk+ot3xpIzv1aNTz8o
vwZ3usVmgmR1/M25qFnKr8uWxR/veUzh97U+yCSm7NP/I+TExIO+tjChsQMO67EV
mGZ52JdUBfAUgfAZmYxqjeh9Xj96gPROTqI26HsPE6Hj79e6+9hgn5dorgfcxp5S
3gVebcPq0A3dqMV5GksC1++hJ7oG1/7BAVMK7nLU2zs7LoG5kfb8Ab+8ccTkUczB
5NTMCV8tcpF7YXeaH+cJe50iwWJGAZ63yvUkRve/1a7bYZILCz8GBD/BzIWMo1cE
wCh05NNuqWEyHr8gibcR+pgrLeXrmHN5M5E8p4o080OrUDiCSlieBsT/FVBG3RKe
c2+cXqZtkYDIzFM7Abe5N5EnEVavm3bV0esNIFa+QQV1b4IEh4r25gr6R/jzzpeM
ppAyBifBLRGyi/lkcWGQyCLnpNrrW0WB4EJZVZrrw8JCpf/pryAdCRbyb6hXFCP3
E3/7iMAIjVICgavM8yfZ/7O6RGzX9xzyI1SJiuTxsHljN0K0Czmf72IuP4oPMi2L
AXgBeiidq8zb9ZncTZ3K5sGDuoibtBNlRqseGeq3npvEkJd1Z1+IUub0Ux2OpADa
XYbpU3Ux7XSk2I0cm80sejmSk30s9tscq7htk3Ix5GbEHtjLHdel+ndebpQ1346t
y6myUHnO2x1xFyz1ExZ4jXZmWWNx30GLal0lKFb0Da0l5yUY6/7ItF2uCjP8xk/5
dwQA5gl4VEdPv2FJ7AY8zTmSqRLVTeav6qRiLYhSMzh9vuW52KuuB6TqWL2PqM1l
z+CkHWZMN3skyewXjWkMD9Q7S5w49gPVA634v8QhUg2C18RSQjsKN4gje9sqFHwE
vg34S6ee6rNlpZi+5o2IANcs4M9GxI5whk554WZS5/6ybg9NgctJWCvQvoMFSJIm
HjeKpXDY8WrFqkmu/wVS2RaKFH9uO8yALeWZUq0oaudFqieawqi3GelCeOwJrb4e
WYxCObkpRTpFgU38nX9eputWDgsSOLiQ9F2L94FzKWQqy0QPOn4g1dAa09Pl67aA
ngYRJaa4uUBEaVUyKHiV6y3MaFyeIriq04XLKlPv596FBlA2Dvzgoz+0/KJxoCfK
P0HQtgHW8fuZ81E0e4lLh2zdPjVOk2AQ+UlN+nrca58xk5QN0u8eJZDZ91uPpYKx
9rjItsrIaXjFciflh9KDDa26r9EJ/MjbYhhdyyA5bOm07/6U7jx96mWKXubHhj87
/7153Pdnpz39eOntl9qOCb5jqrvOlwoKZ7Jkeu64n04bNNBB6aeBe82RshL+2HUD
ge75LytfIxd9P8UplFAwStWs1Vb6HnC6jTxAI9Hb+o/XqYF1QOJymQgReBH09STX
R6xh1g5BR+C2eBGUXnLhiaK0tN2ckWh8hsA+rv0l+FpvDnBb/7A93cWdjUnzO+U/
Oc5HGSNmq+spXcVX+iDFkrq5haFH32zK0ou+oL6ujp6UPbQuDnkuPzwMmXoxbnMT
MTZunIMEp7kCYdTj0VIvoNn44IoVOdtCqEYqV1zwLxCMJH5CKCNSwQ+lACmNjeuJ
v7g3/LLd4+XLSyNPsPFugIezr8UsOzLUrGfFDGYfKB6x96i8ZQPwE6eOxPEGElCE
T8xKB0BEm0Hu1XXSxQsidO+Ai7Rnvp2dUna56qycvBX2NL0BF+x7lrDUASRGMFZg
4zeLC9/6w5dDuVVExVrfdWgI841ynkvlyNmkFXDSiw086lGTflCov+K5tnPDk+gN
dCXFJVY6P9Eqt/0kM/Np5f9kv/ZO4fiom7XEOgh335qEhkAZWqIU/SZb/uUl22u9
LZDRyZRTKVfFGy16+4I9R63/iAZjngijEKmmLOk+BQWLdSLsp0Zu+3xin+yCOR7u
fd1xz5se7t40kC6jVD+WKf2/B6d5HaWxhVhcOblEf5yg3yjMIRvWWNaOOG86InI0
xW3nOzfl+c8zM94usIUtC50nx58nCK13QOhsIKagZ62ItbdJSJ2OgiaqGNvdkRVR
AUUYZeosV5B1i7ANeJMBEZ25y+Loceb3xTI8omFTXlWl0M+qGC57z+Elgukuon+y
PdOjOLHyZ9Vx9SiZ7eTRRPwt1T1Cxmy/KAdinFNZxDz9n9vr5KH90UutGtC+6etV
9pJfsIEcP919eok16WyVvam41kzxflaBfRptPZU2DmssHOvcttNAWmpQ61kxFVX+
J7SUOLvDYqbHO6J8hwsLzrCKmm+IK+rFMhh9QTj4Mlfu1VaDhBsFdTXdhQrIq88h
uqOlcmDZvaIH5tddOVIgxEssCY7owLUBSIAwO/rlmRUp7jNMyXRrsAECA2knels4
JxRYO/sh7Y+jp7/xlx8xgwwFOuPY/K7QnLU22ACue8h2cT5jRurYS2pXPKY0msFp
Q1+FATwbFUN/TY3798IqpksLsmLlus2dxZffbwnPnG1DCJRErRtIn3+gwTYvgtZe
7omTkFiyUthgy/cxTxCkLVDZMqLXv6OXXaw5vNsxHoGljajM8ApCbIM7qgv2I/TP
xwpYtmbEKe5y3SGabaqWa9Q+iRI1DkN8mr1ZyQhCbIUvhJIIVPiEMEriSjdsu0T2
ZUhVVHR5iFvWwzQkRuXku534mOeb3wPzj2JRzKm4mxddlLZJH9vNROsG8W/obC3K
Fv/gV1rERUFJY22GpDrZCTQwTDEbu5kBQTRI1FwiNO1pVI+RgAriVR7DPGI+mCbv
t83mu4xcz74x017PDxYuHw4l+Iz8RyfyORmCMe6pq9j2xfKg/qPayXjUY1/bnoz5
PD0jSxx9sUROjhB+764XrJBtY2DvskdvPAZzyWV7g+KGiAIdH6DTfmMkTh4gnKqe
m/0tTJb/tHmR/unnfXdjPkwyi9LofLV/Dpq07Y7ypxjF+dh1b5/jhinCcu/I2P3t
4Xi6D4MtUSRcmlCNsweLw7n13hP3yM5UIOZ8o8CIdi++Rzu8oIyeo64OhK2OSsEO
aJPwuOFEL8fqR3DCa12MsBHMcNHgD0GPQm/H1bF/D1Zlwgf60ct4QqOfXzd6/HHN
2VtLZV9O7bzocdBKgqC22FASjlz0gxZvWoltzrLyQxlKaWgi3ohoF4+hAltE7JVt
yDip4jdtrDpyF/NKm4LdmpK+XHkHSGXiv/+yv0zHG9URQukCWNr8whB/7TlgzPbz
xCrRtePhWnga0vgsIAzKtsOyPzt9UNyX0yAkzJrW0IWSy1lWRhCfa8Bq9Pv9BzoV
cO7GcDBvpHLYCgl3Al388upK7/3uvLaQXlQ70FLrgjHwryYX2GzHwmd0qzTNjPVx
pmVOjTiLURUCY99aWFj3+XxcuaHkKRF3w81XgXzi6peT48vIJB/DyXfh4HID4OdT
FY6EAf8KxKyrYyYEmBHOggNFdrOSuBQFZ5EBf/nfuZraikUQQVe6jopjCCJhwPTa
Ui0Q1ZljjVQLR9tKIFQzzn33ZRO+OaorfeFcbvjzvYYq9QV8dv/EKgQ5IpjxjUNR
CaQjKE9VBWI4qvp5IvX8KaRPo4ovExnnfMlXA3VAgVQiGUxUvyD3727VVvVaBs3H
F0IMXxd/ZEDKOGfRQ66MtaKygri9gbJhg0mQH30Huvmix58+uxRjo9WYUoNTC4Vb
H7Pik/2CYJ3U/FBbatb12/4DHHI2iltmDFK4/ebMNSbXid/rimKyrgC+vWf11DWf
kzGjOXKY+CpsQPVgQ8V2toZfmpUnfCyiQek8XxMHYAI4hZyXVcu2tR5ROo2iD7xo
7cTubnbI3X4sf+2Rs1xodzkcKJn/GBGKX0WX2lsqK8cdRm+SS1mhNPibE3GV8M5B
t47g0NcnzPPYLm1yhS+vEIrgyX5WagKeVksmWlsp8Owa+zOa6RxSXIyPj2JHjO7V
aAGu7eJGHgwDGx5p0wvk0xUv+3J2UbPf4FhUo6OHYOq2nE3aSUw+wVBxXbayWmHE
kSrJ1eesNSYC6AZsHABSFkS4V1HBK6MByKPdTj4lo/XwhFD5kr2rQa+c+JowBZN1
vsqMIUlhjuOSn22UBKA8OjKUqNbJqmoBKTw0RGSmhC3E+zZwlrTpa7iKyBh52T+R
tekc+HL5eLcgvwnuB6ia6BbD0P8QqyvFPkSOm7hWMIgafUXpq60cvEYfLxcsQv9A
FyjUx+qGNs0hjGIa6bYQfbaXvmcoY0p7Cx7r5XeYmM+2pSI4/ax1pcyx5VOLQ7lo
U2ldipkQXAQJDiVEkzxzW1FCrpkrHNukLTmnK1CeyJutE0rzxDnRRkXtcDkzIfNg
IBtKpgVnJq+3CquH+sIvD6674Zj9H9eMVtLAL/uAEsuSqZ7CvqPG0nfV8zVfeWcE
e6ZdIImARS6XvjjERwjhr33JWsBAxKk3dBAWAM/lABXQJfHZiw7aVEkI9WEbxTGO
7jVbkFgu7DpHoG2appAHDcA4Xn/xVaQfZJJr8CkPF9rNIIPNkXzsee7lIN7Es47c
o8K/yIaoGBEzlUELJMb7AOpHX+8V8V2o6cirXE0uEhgSN0Xc3XEN2Zbk+C7A8LWQ
FdsMfL1R/nTaWtmEwNdUG8DbR6BsxQCbq8yM4VsnKM0ekNavPWWAwKbJrWmMTLaM
j7vDnxi/lOeyBQqxE/zPaHs2JB/HUmE8wUCKIT5Ifao2e1fSYlTjDGPt+UQJoV8p
jGocAaZHM/g7rhykaGbJCicsRik7nyfyxFr/S8x75+kquh44e/TMZbZaOI5E9rlk
+m6GBZfzkhG8UAAm8wOGDaRAg/9B1H7ZAr4qbdXRx4C8eHI5Pi0D0dwX7jfVpOj2
T9agGaLJE2F1IyWrGtlvUE0nHzcgBXGqNcQ1mFk2JEJH3UvONw6hfACikEO0JR+C
LkJ7QT5HyZOIlUyX9XaxP7fBZ8ll/SHauawf2RHl1786zZUphM1vv/sO/xWOsPSI
ogso5SK0PLFt7BVb8nj72QJClGmtmOe9UHGTnvYNNGTlTQnLAl5FmVOzKp0drXth
7jL7EXDnZzK02obkVzqsNQ24YLdoKWQGIqxCpdSfYVGe5Uzixxf4ygXsj8hVYjZN
OWoN1F+foFP6KueqsaGF0CCvXHEUXnx4O+ZdG0QCjXvxbBDJuqG+kf5nkQIaE0Q2
xOZ6FJCC/uSQZoVpgoijtfHGSBjXT28VsYZCl6lS2Dafq0kwSxZ2G+YN4/3kJQa9
+XkJsrx6XVTPEIixpf0b64h+HGVlzJQbXs/BnqEoPKTHqJcebZIGZ2skiSr9d3/6
035BmAlzN5SgS4wSA7fbm5GxdOdBPLCnBFbRvS6A2tqH3S+8KoJvpKnZ+xFkhDtd
HeRZAQRC8kYPJkCDzh5ZqgQWB/SDLu2zLfjj/SFOYJIGhGkIt+31rJKb0L0DlQyV
9AijP2NOQ+t/QEOSuXfU6ypxEHGiWQinHoCZ46sXJyUp/In7nrsmvm2LorylSk1Y
qhYOrJmWmt3T5puqqJk+mzoub7iBjzr5EilgcaQWkvQ2IACr281SRqQ8nhdRCuXo
6+zlaG6WqoM/494/s0MH+7dAVAiJ4Z6Yp/CwnW709VnH2Jmrxiq+h2WkP3WlNirw
zvP0yT0ySz54BavgdNkplSZjGEudTba8UYVrW0uamDpBPp1EUu9GYGOLzots7YmU
S6iM23EXdlwK6lmmelpDmc7tqXUOw2WAewTT/SuOaFH7bTmyEt4BTTo5UiqEF9fl
QujcUEMzFM0lK4Vu6SbLsmaM5oM65Zqz+fCcnSUo48FkCDT5eUAiXJbtNw70Ubm8
pcbDL6Ll5VDjAvcztnpoIvCE9+eMNKoKWyrhyIG8badIqjW3q6q8MHBErpac8WfW
iMZ1pjP9cuwAagxB2bGTNOb5JmmEiNBUje8C9L2mWkDpKltnJoAayQjdApY8iWq/
QKdvBOyd1eZnV4DWk16Ax2iv3TiVi044Z9vYgiNhK9cJWfbOiN3LlpxULt8+chKO
r9w9W4a66sfWB1zV4WVGrDoxnKtoK/mnO4pOd8tsxiHZnSjlTLT6n7ptNDyRlvLY
5/VpHFqYKu0pJMOMXVWP3z40bliwioweCBqEYBjR6f1WQiliaYhogJ3L9rxU9uYL
0hmM32U+ZNG8nOm/bURIIa1HSkcjxOuqk0wV9qzoGoWnWqk5QXnqFTm5GOv380xy
JDSptm02ikkJIGII5AQAprJJX64tASH6UwXTJc92hq/CFqyf1G2wxpEE95WL7Pgp
8phgKBKZ/tkI+/IXeXRwRGvJfdWTmW2ynYy7/Oy3lhUpFNndn7YqCN56DROnSPho
3R7AAqA/Ua42MgfNhJbZIUuBqbPhmefKFGgx/gEInlU91eARu5p3gN5enznulYKM
AVfNCKXiCE3d0AXMYOfUQoqBYysbjKEaBFF/K9OHEIkUH+6/JNqB79WE4Inqh3xG
5U96pCk6gH9igvXjluJYakuXWy+3nu87RxIZINKUJi0qIj3Txl7Ep+fen0d/jeZV
vVInOsVprFL+yEnfX/USJFf+6IY0waRNXCa1fMunADIMc3+uZsvD7/AB6/Yi6sBE
p9onc5v2/Ua0VxhBppwBS3R/eDs9CmBLE0Kw/igwDw1FXVOVDxxgvppEvXtO3TCv
HjVKLNb6clrNw/xS3CRgFwWxWobgcNOtxyGFettvnEvf4FoZDIbFGilCMABu3gtQ
BSCeuQl6JXh16wU524Gki7A73cyKUtpCBRZtb+e0AZWfM61rkk6ns221lNSxXg7f
Vtjl0xV7Q9PmO6qqYBasz0fr5LdpvqYhMI47H2Pq2j2HyL4jRHI7fex5ffEhgRUs
Q5h3eapENfM5Zb9VSTn8h03Gq2OUMmm8XapWSLz2cktbpkDE0Z1+dqL0V7oj5oYp
zAPRteU+A/NvHHux4YncsVmLkQAQ2p5UyyOCc2lGFG8oGux4h1REcWhjitPllq5m
a3jYRd4vcajt5tyj+BGz5YxuXOY1jObQWHFJPgiPbszSrDvJ49bcUWPq+S4Apnoj
1beUniNkawfM1ni4VZFCuchlhfw58GlysPX6wc4crbIyxt0BqkH2IlnqOqocBCra
DAC3Kd/EVGw2db8Kmf/ut2yiyk7e2Ph6ei31ryeeCYllHf1SyF622px6/d4Cvqw3
3V3VExVSY8whLOwUvBQTKhENIcgEUJXgbL+3r2lI4PodsrJS8/7I2P2QKyl7GJpZ
WRtCcFDpo8/zEh+Zi9EhGNnD4U8r80NF4D/oNudzEQG4d+5Cea5rpDpH/wk/rDXn
H/RhXDpyf+3hpR5o/MpllCKyUTYTAs+WvlnsgJ1Z/3k3LK0CJ7qTwyDJ9JdjuoJT
Yhu1NCAUkYQotWgbAmlrCZwdP97Ka7TubwImyx6TTFiEr44QEPoEZaYjSXjgnmOH
Udi/0BQ95v5qdjshQwTXq4zCNOAq/OzuXJoyHuS5HPE9HWVBkYaktclImUNfziaF
WgNLQcwFvUbEx5CXINRlh6u3b27XFoU68ChNBJANcznnGkgwcm+m13qC+KL3TOal
hz733zyUA+Ygdau6b2dwxkbLejwbirml1cHwNv39Y1J6o96kcNx/zuLesCyaJ15r
qttPlPivxgaXWiSlYgfVoMcr4WY8vAMLOFUPT+5seSejP3wXOAJT5xYC0w3m/6bK
oWcobigBN/JMUV1g8SMwqlgyCP5UYJNlOoCf07kFNdb1A+D38rRt7HiCAgVro0Eg
VNmZIbVHnN3QHxTy2UZcG0YPk9RnuPiObmcmj6CnQ75EAMxtAmQON3Z2qd3/gaJx
V7L2sVqykzDBUzWwxSnV/R6urDS32BzFQrtNKgACELiIGZXb65iFymh6UVlSMTRB
rlCVQ1uXIlU71E/J8RwGzyMqekkxB8Pbn1biV1NbF3OZsQGnGNVpNPcnqaRjBGnj
KvbK2n3C65YKC38kMKf0PtCyiylLyCQV0ZBw7t8ssrF3zmLJJ58UI9kxHOzzMSe5
lnI2wc0l1OjKuHrxoBcBGSEUAJKia0SdbivQScdz4kkhMXzcY+ZakRLjv7qx3A9r
hSnBM/ywApAfK4ZcSEOsj1KfPohhYTUeVTf1+uN2AbOwiWYZxU/wAYaYWFVHhRd6
xYTWPceko7ti/AeZ7aSmiSB9DqXM4NS/2BdnYKZKZ14iE7Z7zWU0W5cIe5iJHWZc
1t7K8EAWbDnVbUojDwy8NymSkG9ugoPrt1OTsMv+2sdx1p8u9xwzS0rxV55EJ2VD
GJWbMQHXV1mhdtePvhh8hlEwhi+FrTcT44XL+VLWPHP6VXNJC0wuKomI46nEUEpM
JmsOvFYoHzBuKkbbdJvG6Mo2sXj6sXFDoyDyhOFwDoKCSREcp8Bbvo4w9MWp7bI3
1Rc0gOsU+2MFWA/MFPCWfSwOoRgtR20+mwOV6o6W89s9CNIINSbeuUH1sN/F/oUV
sMpX/BntdpPSKNZZMlcMoeLtA28tWSzZQqUfqQZ6iXWMnPIUZAeAnv2rlyINwVcG
4UQW0CwQTbzCBuyPCjvZcjUuvteVn13RTw+m/DnJkDPNX9TNZTVLgzx0Jl/eEjY5
L3x5ve0GUMDmKl/A6B9y1HXEa6iIuiyO8a7pnWQ6EymphU9KoVLI45zCXe5as+OJ
tvKc3QWLr4ZpizYKv3uD6b2Ln3zvW09MlOjaLRUZTmV8QnXe1R8P46PnXaW8zQ69
do1Db1e7hkEw0vptNjIJD+hPkoPrya+ZYtkTSciz9iLXVpaCQPyAuSvF+7Rs+Ggw
pASgSVboWyY83S8L+kM6dkDNAzPNujZhNUJJezNbGbrv+guU6qyMdUTd2yJdBeHb
Mh9ghKI19gJyk3jj3yZZ8KM5ZvkFo+caOxumxkwku23fAQju28SMv6n1kFudEZcn
e9CdtOArcT0CZQ7gtCrsXgnJNLOtLViKpsAbC50fjGaBSMb+7Piq46vIsLNpAL/6
1Qv/RE/nv9ck3e2kcMKh6ATbrPa4os9Nq6Am8Gv5YsLWW4iryVCuRxg3gyFgYw5R
DYz/7aONlt7ADdfKPmItqUktrERSjVjeNe7CjYiFudsGWzFYj5qSFObCXa2OUMjh
MHYMQHUZKsKRT7z9/Dp3Oh2JnO1vXQApFapbg9uvMyMs8B9BFZ6RP3oqjU0hWdTq
6FZau72uWBGeUKiWJorvrK8RZDBmnTaoUjuMe1F8Q5TMHkZEvxltrmjBxMyv7XwV
ffr6I7Hzw7rBtRpWDflcsqJAaFzMOo/vM/ss8fIDHTdJtRLoOYVmxt18u/lsTMrP
mz7HOBy1iRfyP7cUz7GKUIY8aV6YUmbP3ICQmEBQtAJVRhTo7IGj43BCT3gxAq0i
E0wd7dJc7ErX/jwG4K2wNChocRje2ZlcYeavCw4neTPpl2lK6po/Phj/+ARzSTI/
P9ixBd0q26mjf2gW6PtCt/t5l/q7PCyho/Gao8CpsLcQ7h6MNhV6lEdiSbmf988N
rssmR4ootCstvsta6Rx1eR3DvxpxfPLj3LL3ua2qb0UE4hodKx7xdejhSfrrXMSt
i+fxu6k6T7wX+7pqFiR3X8aDPo6LKNNPJMEi6BIhgdrWC4kh3/QXrtrWgEfBrzKv
gX1ECya5sh3o82bXuDXDN2ZbgmCJWUzvuzfeB4pWOX1utTN9qUUOjL82Y8XubOca
K34fK5DhFvf7QEinoUdPtxkPjHaaBW5QBnM1nk+/6BNGn5VcKFljJeEApMM9p2WO
DqBTdEHcsZGq4CUnghVRYo8In/6ZM+LcE9MoM720OaxmySd1HrOPnXAV88lAtNad
ERxECuwBa0z4Iqhmc0OO/9uIiOnIRY7ACG6WgogjG5mR05PPMHIebMQ3Ax6QVT55
C2ST0nGAj73Z9NlQC+y7a8aBJFRuHf1G09IF/vhWkCUeXJUEaYZUxU2VFilXyIQ6
HV7B8U9+wXyYznK98nKzm3YSJtkBwpuKZ1vmTk1+4EEPUgwj3y+s/RAxxOPaq8ah
VQvMgHvUsg9rsWLS2Lrru0yCH+LfRRp4hUiUKW43zaVhxofBwCwm5rsXft8u1eM6
tkBdU0mZBdCZtSdJR/8PPA3E+NLSstVYrxNKcF938Cvu652kLDVoek9Vv46RmyrF
cHFrl/QCR17gNTi7D/zOS1G6Mz7MExQNJeeKQloeXuKO6z1QyTeNM3vU2/515E6F
KUl2DLSkiWXGHqeLevgRbOWKFw1UVYG+jOvRWOfS+aNBwVZVPC+XhZ1dF2OFipmO
I0+i9urYkJ38PvMEkCNClaSBXSXLFeyXuN6aAIdmkjM5Qr+63X6zaAJiuUZvIrm3
lGrUsWKs/TUaLK7RluVh7px5Fzd8LGxiCjL+goQ28J8N+jD4nb/sDjLRhSmI20wI
hRX6nNKaHhoqtzH3Ute++lFcnyL/14onDUP+k79h6lQGmARdQ/5osZkVS0kLeQ7Z
ce1li8YxqA1KP4TQE89mS9rwskjck6Gaj5jfodMHetKotpNLW6ga54oXtGj784n5
0/GenUYgvnqK6yH8QLCKnSrBeC+5GY46wiRelBInCo8Sy+7yDl0QSgu94zhmgiua
KJlYJhhri5yZ/UYfMtubbDOEwpzmiSDgiG3sWjScXZwvwouk0HHwOhYGwoDsSeDh
ru+7chwAmryCxg+PqwhJ+FecXLTGwficxJKAvQJOYdoH8owJjnGcjIR314+pt6nE
GdJDqp7xVUrjo8FDwiEOeDpYABoGOxhe1LOPBoOObIMqlONiukH0YoTu2xS/PWE2
mw4ofyd5zKZ7mxsUHqJI/ojexxz1R2+Zpe7Ul7lYf6Ia69tHSK82Pm6FFh9ugHcX
qXy/0fkjP1pVmS2pR9D+lA/mdNSYsDJaF0xYXo4ALqGTTxKSPNE03GbR4jCvf9vP
tJb+FijGLho+dhOBHTwfF/5Ohn2sKePQ3DYe6SmfGyBRrkDKP549H9Hml49f3rgO
sWenFPiIhT4RmQnZNQuNnGRJzl9O3BPoWfR6zpA533B1flxA8Ca+EocV2dwWw+XH
/GrbQlKfuSYMRcRF+Gz+7E/6iTYJTIhhaxOg+AEAVMqqW3Em5f4YIe73HgOymno2
PBbnLFM6AW7B2G4LUx/oT9LORxhvegpuHJvXSN3g41rcocqyBQnpRDa2zdhFUWRK
e5dXBqUBU7yl/7nK4NYNZDwVA/SAc+gtQgQRsBmmAnamJ0kAbCjf5wZ7i94eja7s
RENFh5eyz8hvSmC1aaBP8OrpDgyGs5X19W4gsvtDrtxbv5nz/yJXLdJHI20tGKmp
a4N8fYxCT+YjUgGVPfqwhTxjzxBrel51GM/OjEW4yLVhDWDIRwV5qQlZIrA1wI/Y
6MBuSnddr5kZ8DMGPeJj3DMKhHoRrWXMJFWx8deC1aUMWGpD9uRwa5/Wffm9zSlv
CUsKLnPLZDHZRPJwc52Ld37rEtMmWD87s6yUa4QW/XGbm1STKirirI+Narwx3f55
35m0M7aD+FrdkB0zDYkKGfkU2im7TLqkXjjwA7RNV731vo7kO6ieQraYX3b+K4EY
xihGzisYUl0LGrcpjQ7iR9sU2xdTkyBa3scrXNMsPSL83puBW7N0Buhkr/NZft/E
hq/6TEHQPqJZkt9JQ7DrRRbXOkxQtVP4BIMbMTT1W+/k6AYxjbXrpk5BPGp/8cdp
4EVBYbg5mZDUTM1usZgDA+BfRjcLT1YQkfxJrjd06zygV4d5ImFHzjpxx3g/WnHU
7mh6+dR10ovjnNo+2wV+JVf4qxhw/4zWp0xs0EHNsAxbd0e6DmaOIgX8JjE4X4NJ
cV09+C3XYsoTkEtJQk6/gHwyzk5qbo++51Qxt2gXEfU121B+yRP5VZeYlA0vwE4u
z+9c7n2JIpsKkj7njzUEDb+/p+gKqpJyjdPL1Gn60jLv60d8TJLu8hTiggy2Ix/U
Bt8d3rbTQqaKsJLFmI6hi/93FvLAS0NEyEMww69OxqCl5nRuSNZ3BHFNiAGCt8vJ
UsAltrrZydpiZzIBPiBwivnlqwurNW8Lm11j/AYY3hTuA5SauWTKz1SMXzrDxB/V
AhCaVvGMeg/iGO4HGE4Zx1Gr6gfkyzL2OPLXrw8isYKlUAyxJuS1rhz0hNv0cCGe
YoCtWQTiEer+Q3wUYuEQDCanGqm35LMtAJqTjLaR30uB9LsMBSAGxmqAk4O9kU7y
JPkipzzd2LE7DoMeDBph7y6RqVvUWFqFuzEmGzxmVegpDn7cnUIaFJnlJvyYlzay
ijuokdvk5SpYw4eQzuAeo9soZ5G1i0Cd4zsbvv1GpmP/nIi6IyUgP4KV1KTkI796
fTzE6faq/0VKTMGn58Q6MLJ+k8IEUvQ6yAlYL43wZUO8vWXM1C49Jz1kXdu00Mb4
n4PzdpxIx7BN0/UDikSRs3/k+gx3kpotSyVTHxDtr7S9rTjJQp/YYAOhTAykywAE
YDmLUUvD+dtVmxexERtrKgrO0w26yL5o8m3i+mmEmAZBLQeeidFQ/P4Lfn6f/TVj
5j5zmIX1Hymo+gNH0dEwm0G1/BD+fqNEoWXrA4t9iGcORXoEar6oaX/fl+zU9qFf
k/p13wkjIJJhcTIihWwtKvikmnAEqB87flDrVV1orMV2/QJtW6SEtAOE3TqzFB8R
b/GvVF9xuquIR7jXSkzmpN99zjLvFKXsIax7JzWSg983oPQtgf52llNBel11vIlt
/+m7aD4BW+IUVLJMoDWQsy1eb8PWyCO8VC5cRSmdjwqcHRoXr9At4VuMJQ8TziWz
A/uQEmSkAtsbss6FtBjJpqZwnr6JMTN65GaaCpza76uUwf9/IOrF40LumaOOzeE4
namffwMjxPvgHtnjm3ac0hA4oCIPancjUWCz9Aho/lqu1yHfLw18b3cJ1hPnhB43
6plINH1OFFY4kbJ2dBAReBz7f0qMfEZUUVYr987asMP638Ygbq48J4lFTAjWMr32
83B1AdnX4VLLN2kXvR6ecdcY3cpbrdhk2JQ0uzlW9m6ytUIVLf5U+bUWDANGv2ri
HbzAUxiZI7zq7h/mPCDCmINKDXFinp2m/y9Sco5AhQf78HlkvzyTxVSAcGcuVaCu
OjqyAH8w9EMV0fbOl82XA28RHluMUhOVNhWBQ74OneQWo3ev0QdfY1q0QaVGJqnE
z95t+Zp5p3drIbZdh/f0Mo1mAeRQDk30uIc1ggRwqdIrvpI/APzpbOCVsjw8M1sA
gytofuax1n6LzBrFlFerpDDQkxktchwq1Y7PnSpcz+uFK2/rHfxoPniWDhMRmHT2
9HyUwYfUDKv1NPwre9sJ9YcoDkU3gLM0uz8nEfjCHx13YlqN7h0RQumHzrz8hT+Q
71ZxukBtK1RZD4E0Xi473qFwEaoCnK7Pv6ba6VVsRKCbSrDzNzDaTF1rWGepbbFw
anN99GILDdI0RArlyS+q51UmCaJ3A+MtVFgWPU0pDi8cw7dUXnWu/nIO5/NeKj8u
Hy3YiI2dHfkMfJVFfUGbsmJm7iNxUWQtZghtjLvi+olUSxZt+lmfvFL9SkjhU5Lm
DXbo6i3YADjDYJj9XHb3kYXwbyBcuSIppG6f5SjKI/QthsYSANE15BmvFg7zWwd5
m+f5pos4SHpKzGr6b0nd/1t4IjVgjabnFEihBFIxuDghbNMK+D84TiEkAAncd661
zmJlG9cDH5QAxaBJsdvItj3kLk3poijHTu46NXnGAxcTEsXM5NtwRD8qA5puKj80
JIZtEcFC93ovoxNItz9Wf5dAtPXslZKB44fAhdcObILk5eLinlkIij9JCcd5Vhji
tTemqIoYy3xPJg72oy4+Rgq+m7TSzTnB6Jmffdkk1FmGToI9cxSJHN2+w8plVLJq
GtcWxaI8Trx4MotLAg6qkUaI2gVRZ8aFMBA8J2+0q8MAtKpywE/R0DqSYG5V5gcP
lqGQ8PykfJCfsBeJUZ3+0IUORHIQKJRGamGaIvv5Gr/fpSNfGUYEPdhub57WdRcv
JWepstJbX6QC8WQnmnctDE9c7xew9dD+zEyv4vJhBqeHE+JYZFo3uuPvIVSq2y5O
tdrRSFPHoBr8pDAH0Z/BWqzhvli+GDGHryesYc0g9nqZvC18Yg4wg+FMUm5T8XDK
vx+z4b5wryPMUtfMTpWEmqqC6xup7eEobK2SDedmuk/e/3CzlZ0IpjEUvy/fiPV+
Lbe1RdUe/OWGBVigwBGNJwRLsxCoZfBO3tb9C+N15ZGQ8P6C+iqQBG900H38QtO2
1c9FW8RqQyPmm+/EYQE8JcM8tbVsLuVcLvlcF/EF2h6BkSdJZsohvK7Dxn+ho3k/
OAbhpnFrPZmY8KulrTQtrQo8c9OMEcc6BDGaxTb106OLEcxwOZHzQDcPMgeaze4T
H+HxqjV2PdtBz7j5Q+xDgIpRfi5nLMCBE11ex72DAvB1czBgISAgK0WCe0TFxIkY
3s5LWIVRWeKtYbEshzofzJegGq1qeMI1szowk2jDSq8Bt6bhpYjW3lp77B9E+TRi
vnlQ3CC9ARYuUKcJnG+m1RMRXMz53fY8mbhRaW/yiESPXT3j2BDWpo9ox9Uwyo0g
R7cvJACbxTWmSTVACLKRqEBU48WtBAgyXNwuBdSFUB47xhBjkpGHo74Ic4FvdI0d
bC2hgkFdmLen2WEqIvbjCU3vJU25c01D3AI80r5HK+NgJQlbStM+sqH/f1a5LAPp
hg9TlBAt3i9yiUCvYJ7L6AQFNgxrp9t1eFB0nBR7sLpuHS8s+U8m6/fMrZH3C8R2
zRgl1Gi3tIK7HHNyMFpfV1YBlkg07sb0z37DZVO1GoE7cI5xWRUzhrGHtjCm7UKy
A5GMp0Gz5uyzcD+AJI/0wNshLZGe8H37kz7HXZ+h44Dy/nqboRVQ0foU031b5Ird
z4TrAR5ui9BLNRNx2iQhzUPfKgMzKGL8PgtqPZYRCP2NShvmhLI8pQQXKY+qmWjd
A8mkawuQ/gSBG0hwiGnaC7doQzqYL2hoFjrriYuWT1HfpPf+BM05DL/sawfvFLUl
AAotWWbqM6LXarTG1qZW457SIcA3IZEOnLPWmmAG8lEo6yR9Y4ZNtZvJh1YNzarS
W+j3SS87FCvk1e5wf9V9x0VWmcZIHX/z1RWMPDmh3kBMrwPPLNnHcAtq7+p4a7H4
5DF3DirFY4vCptI6ucgcSrCHHKL6AXYtoTiWhKTNRyYvy7v1fKnmLV6FaraU0xoe
J/k5GE7g0/jdGMcPoJtMlyzZ2RH3J6VVcKILNJW9/WrDjxzMr7LsvhOOdLgfAncl
EcsLxGWoceZo+nY6hnqGvR7wUlwwSeqZu+XGxIKtULyJLq4FRqWw8NcnvzNXnfz8
P1DqNYDwlXuInn25s7gF+xHOAkUkZ2AEjXwmuJjGr26eyi4VYEDw0wntidGWzor1
Cg+NBY9rcsrLm44K6hx1rDgqyfkqDEMT1qO4GJXXjTOA2pWIE3YshU4gM+/oBHbd
XOzPhhZJ08QLILXvQL5Z0gnF/0j/jZObOjs2m5eSs4yleqh3s6Ok9fUMeaEFEdag
pSPwSb9qQjovTXC4HWiPlPoqBN4U++uWGPUPK6CWhAmfxh1t619/kBsKF4KYY4T8
21QjRHtj5PFql5KEXGG/TT3kw++spgcD8jaHh8atFlL/BDx2/EpvYROS2TbIzRwn
hsGgfYgK+V9p+nx4dFpPi3Xu5dg8d5wEiWNUuih5rldK3uXn+ALTHflHT+Nm/Bac
Yyybwbx6v6m+U323wHmtdGPQlIb0AaHQUgFcF8Ct1akr0XmU4Pzy61XM2tM2zHYx
PenPYVqAq0RBwQBgtCXz+x8vIhYTi4CpYeMj+B1xbyZYlGo8DD4Fy05WKtyCdEy+
0goWuXSqBl5g6syHU8yLv81pQ4vqvSQa+D4UStBNOM9YJ1X25/0Q7YkiDrcFhFZn
xPLQ1Sy50WJNFyr1VZ/9gWi/Jo/Bq7VfY4V7W8WlbGUmHzcxUSTOkhKzQC1BUTg8
dIxIK/dGRiH2RHHN0SkYQuGlomp6n+l+FtnfKGmC9wJcIdAoyvNX2qcKLZNmhA2C
SgHfU8tpvNfpD/pntci8zXD1N7D9I+DPzER79jeJ0AMg2rYFlPx9ui+/0mRU0esa
LcaC7O6E1y9leRKQkfQtDX6XU3yxvvnuuM4EfI/+Thkp9ShTRU8jNcUq5vImnwcm
IzFvXA3Z5jI2nb/R6oHuKB+7NJlOxq+fObt3A2yGhvgWie35bML7NjoQRUgNZqTr
ObWYVryTQUSCf7K28z1yc8hb6KG958i8yYlq0PRzWzAODFi4nNL8p9L7enpdPOY7
jS+3JIFWKDKgfUeL6u13GfODy6buKc/MiGgX/r1kGUmPrfhu519lQTDq4ze+lxtL
ALqSEBopDhHX/K3M0Epv9RFamqJs0IPfkb2QTuGcIjAl4UjT98Jm8pB71vn26SpG
e5t8cPQZkEB/ugZwtS45DRc6Fqfj9wvyFjXLPHWgETpoKdl35EZvktmWQFoFmxA9
GCRYbQpj/0hTeuoB86irYS6KuzCbsDd9BfX2rrf5Ksj3d1Y6wQeSDSHnXvH43P4u
dsbjMIK9iu8xqtwshHYbwk7xoSl6BUFwYS5BcWuX9MyLoue1E95JxZIJBwn7rHce
DVcDKWTSgUoQMLA8TO2olqkP5w6WLPO8zHo2wqd6KeAKuXOXUr2RZcWpnE0aMlP3
k/0i+52pqxe8+R09Yg3CVONsGtWQWlAkTV0Y1dFAaqU/3jPoZeqvSnn/bVIVdrqc
yd/ybU8Qs97NejbRfG7gxbkx2LQEHCTSbvXg/Ojqkxbh0hBiZa1szMI6mQ98XUDF
RExCLHEEFtGa66Qzjyp3a1KnSXXcoeXyCEApUBzvwpb1kX8MBvZQaZPlE2hN3Fbq
Y5UOKlkWm61gelwENy2/1zBA+5Vfrv1wlCiasJkzGK4ydJHUO7TRDotlgG7fAhNM
lyZciwRTjjaG6gBBvLhQC323O8GaI4SxaSWkTsrGT4/WlkkLGmE/3cFyuHeeikcU
BUlgUVGM/VDwIAMMV132Lgkl53dlfaqsXoAgz1fBozTHuSjS4psaZ3T7jxZ9aOT1
4gNZwHxZbPFfyT7UDn/IGVz2cKp7gnhwRCndsyRd9a4q7LW5nz3bJMHzB02khPNE
CrFg87n6KOuI0iZ3vHmb81P5SNoLKuBaRJBCXTzFymxEv/QunQrfFguJ9pphmppO
JRmeR5ASeL2Mp4914e/8HEJa2cZBH5C/n9aoK11njQ2+O/4ScvjlsjkJjlM5U0mk
sqX1VdXVcnGHOxlYk781/2h00BUFomfhtaVfUAn5V4DtZc04EqH08RPfgZETWUry
emksVnbYlG0RDOHY7c4CJ0eQvL22KYwyVO8+y6OOVhQCP9ddecnhSc7J+hqtCSfn
eFQenmgOZFmr7z75iVWhjRpJCPDAC61sT720srcZZE8FVYBW5P0nxC1RePEusIEM
fh03tDJEFLoqidpf/jVtQAyboYfUjUbV4nL1TY06ljk4Z7l/RyNdwo8qjIcr+SPR
5kkRzNgUOFcQVDJpSl8lIEa+Ka2kurEIajd6icfkTUHDwvcCs/403CQ1AnB9ZEiF
I2+qKmSZwvX8bUpdo/QZsEFDZiBpEh3ZFtFVhRO8Vi1hDeBWm326ciDcFoXAGtRQ
3+lF171i5nzgNYbkJEOTXhOLjLNvkCBRIjWp/dXoAsrYdrbq1hXka2SyFWZ2cEbF
YIMp9AhP4QpemsVzVdqM9ZTpeAkq9oltAI80TVWkuUNOXE6ZWHOKqP6oxcPR9Kbu
pm0ItmBXOsJb13RdryYER+D8O1xXPQ7+SIq0ejRRT49JsFhwvO+W9jBPjaZdZIl7
DUyDSOeHoM6OXBNPcB8+8fZN12Dh2MzSnWdMWYBlscHzYaYyH46PYoGb/8q2Jo1g
3y8Xsn8j9PGY5RYbdZjkb8mYVDNpqD+7WtA4Mij0VqyXcMe2qinQ30v2iZPzqxgR
R9kiM7IDhSyejeTdcUpyDfNn9vlsWbJzoeuRNarWRkyA1J8EEonSzjamqVS7B9x7
ZvLT4Ao5vjtMgumahWWy6wJtNnk8n2VCfYfHVZQqVh2cTNEbXN6a5oRB3BWOTOok
UuO6P+y7ue9c5oL/lanzUkGxfpBcqLdxbT74KsY7fQ4LtkLLE2VvubQS0b+F8Y8H
guK1KDhpnZDFke4eosVm8n38buIaG+ARlxJeXeha0XWMH0ard5z96fB3G6973dp5
9EmyCDA/0903YUrDtR2A/mzNraBCg4TtI4vMQyXNCU8JJ0kO0X6Z+offnkqAYppM
webVk7XVmD0XYyDlpP+PuvwfDNoq98t8/xyG7dT1GuRRa9sKfEqfH7IBCx57UNBF
DcM4yn0h2shB1Z/hpKQqo646/l35S6T500CFkVprZF/X/LevLRMhM5CS1Zh89Yqo
0e9ORUD6/HaTNXSqNiEkCzeqKqAfkl51dP5obCnXIV6uLL8zd3789YVeDAg55sQx
JHsgiv6pEIoTUUql6h+HId4x9D6LHTAqV0Cz6/hJdCOxNvpBDofnbKHE47WCMy8b
N9kPCd4SlUuCPGNF2HDwuUgT9kq/UaRVSg8sWpRrA1iRr4skZxhgzQMmo8/WDcIV
qdM6rWHB5gE+QlQr7BkjjCxKh5VaVw+Eh5lf+vr0cckFjn4YkotNTDlf2HjL/5JN
FaFsWowEwVr1aUto+ZuFyZ1VxpM+19w5TcEhRs6mJ3KC/aylG+I+TVFSw0qtI9XL
IXTx6ltQBsZdmUu1m4oSLvMf2/cwiZQu74gMKmTOJ/6OZR4NxiOnQRVgHXtYeI1t
T4p4yFjwdVr5x9dkI2i8dFbHj1kWkncvv7oEvaEHIi3end3Ew/MQHGfs94uJ12mo
FWp/hWAhHBmv1W2RNWmuzfpTjl6xXL5cX1doAWzZNJoZxldR/8osWiBNGQs2lpXo
eMS7i2eQRAiJhHgfOOhInmXNxemuNK+o7m0m5PfDszDV3kKtwnMTZpfqPsES43Ts
xmtm0hn9OjqJvCtC3Z25snUd2oegErMa55+V/wmtzHfm9Nop9lLmf5Itpi7CpS99
oPg4WuscdhQVbt75gZ51jcdKJHhBIj62ucimRbF9ohwwzK4cOwkRPvzTlSR2AaLr
nB0PSf3R/Bn60O7BMiPnGxfFanA/5HE2tva+EtxzuEYfKD6qlATaT1gKh1tOzYX8
KkyHhDHuLkqU/Yh3M000lO+xynPSrk2hWR98cQ0b4hAVBuYmFzrArXtT+GPRFbp1
XL51/smVvvQwioz72F1gs3sCcuM2Uz9x+bszQCi4tzcreTQhrq6p71/azA0sEpnE
c4Eeohhg39hfwRah4YEfwN6v8TmYXZ89henOfqNkZlGD/h7aw/p3hPz/X1B0zYz6
nX299TiZb7LDx6iLOfqnkTUKuIHTOjJcmjSgVPirgB2oZFMKh5xZthVxn8NjfhdK
oOyruz+56m36jZgMV7WYKFaio04jXTpBLh7T1N3164DaXS0cifhey8sGlZUJsKXq
PcYmyCSIFya3A85hTSjichKQ/BCJDP6Xxbqj/vCyaf+fvGiKUMdqywHwza740A3a
yJUOTfig0UvRtZfrX2flBVO5YhdbnQiU4BVDLXgMI6vUpHNtEv4Di8Xwtu44g5tQ
xDKLiJYC5sMfXZMMXUe6qsjq0343N8zeKLo79Wq7mDJXN8839SggKiX6oZLOgeRc
kUGQbUCXfsPwn0Ye2FU47nC28/6Ew2z1n3nkrJFW31yVblkV2J64VXmoqyrQMzlA
l6qU7U5V5nQWqmUrj2YEv2Eq/NLkAaMx70YaBdM+BLWySzIErfSVhrg4FXSaFT6a
e+BMaZPdC33mRYvIGwwwBL8uJd1uVCRBG7w0fqk8PJOZOtX229aVNYQVxJ592csD
yAumEdro3zsrj68Mw3GxQhgpqNoZD/eppzSpWFeYFGEbghmdTlEHmE8D4J95NE+w
DMe5ApsbWiJRGZjbUoQlvvXVM07wrzDbW74OoIxCgGOJjtHV3tjLWzW0eE3gwLHY
1oZLL2NfSppo2vVDMtNo9Ij60i2Ihok9ynt5cJFOdTj94hK46HXpL/0TlixVLqec
kKzgqVaKrtMH865rkmbz5XuFSe8wnfCjhvVlKAByMyLrZtUkCroZaNrhpDYtsguy
n8nATQrGGsD9hnY/gpSe+w7b+Jlv8Gm+ZyO05MSzQ+oPvPZQ2ShQS27cgP27qfLI
1edHTGBQagAi4kBypLXqnm0RTJGxtLqd5uTCENc8wruZhNePakDUbpOWXgGfu0Cb
d9iHeGBMqyzK0PSBgoH5GDbYhetMzpih9F8R1WWGT1L8lB3HDcTP6S4wW95cX2ff
R3Qv3JQMnf1TU33a1aVxYmat0ma7isIEYf15S5HrzTQ0mOpYMaaml7urWoRF7L1L
YIyfRDNUItJvJvj2Oxlg8ljxRMd9deb6gobxmZX9/YP3GdljgHD68cIqZmTXdHl1
Zchk/DDfFrF835KmL34VWxMcBxmWx2VgleZChxnyWKppZggQk164jLVqNupCId47
3WaQ8WVc6Ya9XzB5dmIWthcK8He1DoQE1lhN8+QVNsDkml/4sPvfv28bRJSSGb+3
/CR9LcZAc9wDQMY8poTQtxFoM77YjIgv5Dzkl4Km6fduBIP5m0yqKWd1QuRl1dpx
NoGpa5icF6gL4RsBUpf7f4TAfLPW2DPuWB+W3NQOxUBrPpmbkBk9cKuFobX9bEQy
FMH7alSdjRg77mXtRG9r7iXIVpXsX3GURb5YKNHabK0rsVjqCcbrzJzeSrNyRu7W
F1pyfBTjy7omPm9roMSluAbh/hkZRH4FKfSL/dgslQsuiTluHhdItr8UGF5CG5/2
W7cza0yDfEkTHHaIxcdgq4kKJLGDp3xgE+x7oEpmQxu9H7ySVJiIZW4uREnIzQQ1
6CvbhZf0rSyKD1ywAuukv7Wfg0KTm3dmCO8eJbI6DrgYbbSHHftTak+R4Zv7uQp3
IlkN+ycxkonBMDnQdIzA/Nrv403RNOgfHUuTL1haEBT1glEWD+fW4HBrACzOH1/2
D2KFGQrfBBFO94/fLowdYa27vUGNUgBGiNLW1O5JESdrVv6MPWySkFNQoGY4gUoI
PZkwCdVfXgIuWX+rql4w1bgvUBE8A+yHGlYGZ15vWSWjHo0Q0n5aeuXOKOUFP1+g
G+DSJAUSQpN26q8tnehmmqdhA4ng81PHegKJdOhB4uL3tE27sMhsmdOKiW9WYaou
PlHeZEKZZcDJKgsLzDFDUyY1mga2eNxpBRx08v8NQFBLQ2gtNTRGQYFGLF/l8EZn
GrocshhZVy360go7O5UQFbTJnjK9S6PBSFVJK0+GhowC9i+sCok0+ED1RtrEiEUI
BLgCtiJ4uUP5+j/W9lNJ2FadaNkxk1MSbSt7P2IWZXA2AXtl2pJDPhf+vvWsA5HT
qXCYvAGaHWa3xdubZsapzhr2wkRHvJZUiJdEkzBK8OkjSzx2uSLDkhN5yHJLbGgq
MUlfjTYmM8FUMeTmZKiN2jgyTX4S6rYfhdd9JCkwX14q+WiE7iWXBmJKlqhABoCj
uIO/EbgZD41iKVxPiy326G1CTI7T0vJtgzuyhwkwxcVvD7azVfY0z91VfqJowGrh
unCzehFgVTidlMS7qUDzbGOMZDQg+LbgTh/FsrT9eiDj7ggw7g7sHe0/W6lnzPdr
K775LGTv0k8SrUvLH/1xEyLd2LU4ydWZ8UQ42r+xefOj9L20SCEIWWujsQN8SUyu
VYZxAHxBZBqiZp/8YQaKknL9TByXNiI0nmyKU6CnTmNBM2jNwojNJI61RnjKGh6X
s5n/A7wRciE3Y1hLAjCj6vCPOqByc+6e5+ciGsV+0BIOpo3vHvYP3pb9EEsv4Tnl
fmJVTNQQyEFsoW1uDGGf1u6XA+qRddewWrQM3jxViwYr4a6pcoa0r0MwWtlkeCSg
ae7y+hzV3/84ErprBou7QjNx4IozhPGlPvn4xdPI7vJD5yIDTVWIiQZTSp8zFyq6
QK+XId6oNeXe3g2qmqv0+ZruQFtSJZZGaOrMZVEDdPnPSkGdAXiJ5kpTBEN6DN2e
X/TIQrhGMeWGgQUMhzUJxWnwVy0yEDft8VLROTsOl35D0FG4nzYQihe+FEYmZIQ2
cv+KFpBSYRv6fgs8rnJW/EhMOqrdC+O9SFL2jnZb5k8tGDjh6EtGD6Em6FqM5Pgb
sdbndToWReJiUmF3vpJofT7dYqU4zmEw44HCz7kFEEXcZNcfKIAo3WOZuiFreVB9
+eV8U0G1vCsiG7GbbHBf+fJJ5lspiKZGg2tRz1Bj9HOYiiuk4UWlEUm2BfqyknKR
zmL6NVheO48y7U3asRBZwDedrdOEuATF+76LpEyjOFQITpwqzJUzSt7g2gSXiDqe
wpwxbNAOo6n2aYYupxIfnr2vqQVA5aeAGdfK8VwIyD4dNHsCnyEommTW1C5u2+dp
MEijWRmrVyOPgerxk1XsLhCwsdwBxzp2/2hwrmGGHrtMSNzUdkZNyPDFFw+We+ML
ROe1/4fi6hsyyIr3QJqmth347CegoZ0VTYzv1iTrMc5ZrthNS7Ollf+kGbDkbBEr
vnOr6KDo8KGJLAH9WJoTK9FrSNF7fJiDt+GWqz3cf9Y22jOCFnats4P2mib0+ggg
99qJAtqyle1hd40MV2z2YCGTCsNNCcvUz6MnABKOtaayBRmohmOBwiMyTEQVAdfG
u0zvtxkMBTxZu4icrHmk/SNQHNuBR1s8dGaFf+/IE91GeAc00D61lfd++18vRj1M
+oX6ElOkYM18je2LqJrF4X91SjErTOvJwPJ9PV/Qu6qxdRYyGyVTu1xoJ9Pene1O
vWlr3ob7gfTGjqUvTq2x4UvDSIOQyyPGCdUKdTTQgfNQOh+sWu0KYmRKAu9c/qZn
6hm6+mSZDcRw4LeWlU7ZpxlFlQXmu6QY9TGY2ORl23PBOUofNw/5cYGfYTUArScw
3cWTpON0gFea8TpuI88nSNtJUe684QLJGueOcVqiz2MZo2lIrvgi4jO5FJiG4mBe
N+vZiedWbHf8/x3CPFRMVzjel3kP6B7GJIzIoMBxw9SvI52pCB+wAjbBgyw2kzxd
9/QXccMVvrF5LDyUY3ER7o/hqaqsQ7oQNA5CFsFj4YcZhnYUqLQnsRwv2AGBn23L
jtm3ilC0LAGajI3TKzMLv+bUj2GwjrWHF9JWGC5L/Rz8bC9MgZHP7Y7QIurcpDV8
lUUIhmQMDsgdFIVAoag4ujE09CWtWpdg5jL6X6/hxHvGkJee1JV7itcqwmHM5jq4
wOmaGsreqB4jkrQrq9ii3GC+88XcaZ/0QTuT0vs8zVbp6IlFEo8oFRY5C4XUqOu3
CFQldZv5R/AnOtQVBKAHVY5ULse8pU/NJPmpftGp8NZazqf6hesTdyqCXFkWi7EJ
GbPObybmB4Hpa9uWAMuR399LY2VSKXPPIWZF/AE1ez6U79ySfgOQhouC3wNj21m3
gW2SJ+pPrFnuCJo1hUbgeNvDg3s2Z1rPuophydfs2MOzLYuXytdBSQ+4ROszpRgR
S7dzU9a3iEiOYmmSMeboJ5L1TDQLjAsygwgNEfFvgCofYHow4n+3hfn+nQyxaGEM
X/pf35dQtw00JsrhPQEtcmu4N/mKrWuoFpZiFgDxiP1q68GdIU1LT4ys5ESM5Wd4
o64ZcjEi6JF5IYZXBJm0f+aAux7FCde42hZZ4oNvYB2FOg3jWGjUnMtT9xflnc+g
Cy4Y8I8GaiZQo9IJshM121Q8TDNwhhWDzgNHNVtIB0qDfIZ9ABWKkLQ+HToq5tHu
T+lS1mbV2c+z0nlKkqoe3e48QpSgf/W1lnFKQE6YF9bgl4i1YUPx2rRbI6vlD/KH
cuFOlQ/f2Agyrn3dS4Aa3WwFKsFFOl6WplmOQIIqoWjIauFYHPLBpGBR6pFTv4C1
Mkm1cQbPxjPuGj7KUEmpIng9h7L5LnwG9whhcQeFZUmAXyKJm3z2K/a6Ih55fEmX
xrwjUY7WW+dwfqp6FU/i4GzN/ledbOzKHzXEypyu4WFJ2I+ddtweuLuBRfH0GJIF
du5tMO6OSREZ/7ZA6LA+8wdOIm/mcn1lP/iPfRM6wVgTLKhR9GwBsBCe2WElHtBf
PYdsGbc4vV5SV4NaYlF2kDWjkWwM5CVS1tweR2axQCMYwhmojQ1lwBIGslvA/6XC
NgMoV4uOxYiy89LCvlXBR/BBwk/RSTFrDjhejD4YsObJaiiIU0rOVQ2M1H9vbGe6
ieJawZ6SzlEr6Jp1Xi5f4N71RwczAu3Hia+rxKu2+l1kTeexus8g7tOiTxDx4t3V
dWUIpXMhdmq+B8CZqgNK1cganaWoNWVnRoGTcb1HsIwpNuvH+wgdwf4qxtwrQZy9
ayq3J1mB1zMRKnlqWk92ytq6DMvWoBBXjcEZE5IfKSoPFRouT5I51K5yj7eC9/DC
ZmWc2D3Ae4O5VVfz2FiD/r6pkW7nb/PAxP4AKWyGUO72ScSApPHuaC0jlGJC6ecy
tjNtYhvgFvLwjVsFmUKYbHANtiPt2Eb/Owlh0Pnf0bAs3nRaOoqj1OVhZx9lMg39
wW6fWdC0DZEmuNxcY6ddzzFTcQ0yDybfXPh/PHS+cjTq+tKLnosgbK/Up07qlf6d
9LL8jtV4k+EwSmGgI0rktvXtZ69zBaHqmHCK/nsuaoXvaqO4isZq/LqJs6nHULSe
hpk0IDJFTZaqEIAS24zqvGpLPwO39cxVViPOBc/GBvcRisUtzuelj4U3DV0FH526
OqpXNmMXOfHKD5l64BcMnsn6tj05epKgCJKCHAT+kQ4qobbe3DRtSox+zZVo1Mfl
Ghgz3kQxxcshK+V26LXMXNGj0LscZPb6myOrRXWVMjFSKYCobR30vvlTBqLDuRQp
kqw9Gj3HOyLVjS/soH7c6IAqtI411T/9Ghu5SxGdfkkeAlX+J2uhcjJveLw90/QJ
Zg2ZesK4xsF7lhrVNCt8yA3NeuxPuzjfv4MeIp4czaRpOjwTvdPoHyRbylySRKMv
wif5Gch4BvWQtroIp0qQoxfn51s2JIMuYQhVkL4ad3f17m3yys1fxVsNisW2bL9e
W+z5bSz3WHcoDvCV9F+V1anraa7/XIeBblYbZPSKEA3ZyXQVI3aqaZVwf6zJTqUJ
plXKFaJiMW1FZYVpAnXkIm/+r91JDFRFN5TdBY/VqmvQRTq+Br4hS2kjEBrWn0Ew
x+EAFN+fSqa+nS6GkrCL9y2xBBwb9cibv7HWMc2n4YF9ABGsZQR+tErKQ5w2BRHK
LGEdhoM9JBx0WgMUhV9capYSuMAeSra/ImTibD/zCLqtLuyg08D2boMifIrWmLQk
/q1QuLjyAV9YANxy10J8FV04jzxOZnNSaVGiH7jXP5B3Gtzw8Zys9O3t7lYQP/K0
rzAmNG0Q8YjDczg9TM7O10lAOnQ+rAFmwaC+PkDY0GXYDdFX6injeAat7MXtGdmk
+Zb6VVGtmiGYBJuMc/yUpx0bQNZ1S+1BJW2ck6Wsg6+dfV2HuupcAnsEd6J3wuLc
f7pReEJbMvAKb4Rkb9IeUUBRMElpXlT9Iz8sFHTsvBVyPEKpKD9YRtR4mPBFlU3E
A8ky2TyU4VzKSwMen48zE8lFEO6Of24oouUc02SYMXkMBCi1Gl2nFMFtG+oMyS+p
luR9PAcQ5WmijaXEIcVr4ZORlpq65RgAt/qObVZ5bF9peHPfNIp+P8i5QZ9vGGcB
/JP360bqLoRJLFj7PfG8G2K3X8yDtRAQXQYSLoGGFjML/0se4PCf8RRXJOGAj6pS
on2c7HJU3tUblj5kJCoC1pt+b81pm7RtSaI4BL2HwaPDwqhTfjUe6xTRG7JYjAi5
d2bmfhd3jlrLs1jUxfKOJzQMCIGBCUDJjjQEfqcCa0f3KA8g9XsgeJvs4ioy8iZD
BdrouZdCcsDffvFEIxNWh+3lGz268BvUN/Sc9wFwHgMyLgpyXr2N4XaOLH4uFyXm
5UrIIv/4vHJHLJ+byrKJSOlqQyfsnOaVFLDGTB6ARXLWAKqGyq8s9jPohuFFjxA7
NjMDNh11X5YxdRuB0S3mXk8TVgnYnCoYtEKICBbIMxcDWUvP4kyZgHk2+sWMSfPt
ofCg36Trp/BS/P7mT5CjP1jv93vPFpdabVAkiLbtmaNjqnSN6t8YNs4IiYzMX+fj
jZw9a/6uTybFKC7IPSBsPpyJVhO9QC6EJtB+FXUetHPyDHyMN21ZafpvkskJvfzS
KJmuscWH8smnqLzJ6efuQGShEKBM0zQJRzuU8t9gr5k3j4N7/8aPlJ6m4Yc6zj+m
PDJjIaIfB9nyiwiQAGmIj43MKY148Wl3GZ78Q50f0kdQH8tGV0OgPDYAANCplPTP
x/YGU+Onx42V4Js1mY2YHS6xKr0krj+/48d5qfoShjlU0zfnoGMEq6Xb1P/DFP//
qFj1TMcqtodhHc9XvMG1ZSgbpzIHzL+TW0RJ/NKR/uy95dx3+AHvtWcUnoh4JQgj
05lt82hkgln6isPLUH4PyT8WCeaF5bZZnDaVd4CSxJWZ8egOW5Oz2HgiAQn0KB8b
omOQd/Mdk2At0oVeRXsGBTX104LA6+jXnKdrVO1XtsN/84E2wsxuRRKFtvc+fu/E
Ib5E8/DP0x88BMuBmh/XQEnMiTCqa2hMD1O2Xqi4KghExs5pw6QPPzbfZPVtVsCX
w1bMCPXD6PBWdKeIsrugh5qT6B6N2XMe2IXnU5aIFa7vDkX1+W+5+/OrX230E7Vv
F1FUKKelUynz+qyAxiUhXVQtTF64qA+TAWHLPBSKx6u5nG3W+Gm8zq9YEZFCE2IQ
EWM/zpL3rdkHmNy1WFsjB8qC7fWISNAuhsWQTKdtq2TXrozSj28Yb/oK/492Dz6W
iH9bQ68yTp6ERH5e4A/RCeLjDaegZTwbRls30rUnevP7SHDjuEu8V+6xT0dTC+I7
T2o044/sgiD48txy0iTNnRyL+GohAkJbhPGHTAdHc+xSjeq2e/cbtdJlZZzWJ0rC
zy0vyJQvPXJ14ZsKl1pAq1DsYzLvGHQE+6Hfqx26OWrrRGuW0ji2aE80n7Pcf0id
YrOOFA7j2kE9YZPAGXzb0kn8x7T92QWT081yR6ssLy7En4aiEZKi1ZZjyX84nUdH
42Ug2p/+ZoDS+hxGRoDXjQfzD54hTJKYlXyWA6ldorfS3UMSVfV+Cht2Qrc/4HMX
bE3xyzRRBHUylp7WZWJTrGLaN7dnTVEQX2Q/Jm9z6m5s1vfKZM+0W3BmRnBDHvDD
QNTRDuGKVXAPd0Xtzctz2jlx8tw3W5LYiwjBciU9i7JlrY0l7as/VW7H+4+ekTz6
FLMO1hiEdNdTYHaDL4neUxqSQxsXs8fGZSj2+j2u4dtobFOfL20WguGFZK/4DS30
AosAafqMmJVJd5HoDdV46v7PounQTkx35HpFjLvlvixylEjBoPtfXibifk3ykawu
NHkYEpHfjS9QKSclKYOsZ1ReYWqPL7Y69Jh4LUTOZs3/4p4TTweKxt46TbefA2+1
436JM47gkzSx7SoKApRNGoRCcj+BYxUucnob8dsjNg/2dSGR+6N3zLK+3Wsdm8CI
PuWYpMHa4oBBb92HtcAH3rwQKoKAUKIyQt8bBMPRJ2CG5gDw1dcHvVRwQZT7xCyz
8yqLsvXW6aXJ90DGTQNIx2cnnsm8LJmpprQFVuPNhU051DKjSCeFaRgPN3pVJHwz
LD+Ifdfen2xDAYGKfr6u2xIXvB5Kxzzk87zqf8gP6SjWGNDHv9k77a2IKN4h12lq
HcsXu/B7uGLcLwjGPuds25dJODqf+FFwx8GmgazD19vQVQUJ0Z8Lz1pM7F8xbTpL
ozsEFMJ9zYlF3iG2NsYv+UDtQ70WGUsLy08otVwjUVbjKPagHoFBL4199m8C6z5w
XEAYrl463gYj9gFXoCxX6shy+JFIt/4QH1B1Bt+PEAFcjajfZ7bA8KEP80wlf9Hb
yzwvv6N0IJ1jzSkVHHEyyeFLXREsdwpf9Vn7nRZ88IDc3rdj8/92pIIELlY8bFF6
olYszndb4DWUUuc1zj2zbd1kCbTbWD2dROIb1y2ne7eUk1rMn0WWDa3FSRUAr2sO
tMyaXxrGPqCVtu7nAz+2VxZrMq0iUMFIZ/WlVEhFzJ3iD1LrayWV4sGXiU1TkC+M
oKsBxZtPRrN4xWODneTMkY9O1oi6BW8oY5PvzZS3wzMdurAf74pAR2UGHLr9oJr/
79zYYq7PKvhNUolkqNC4p5ftuy8BdgxJXLKzLpukVuvns9wQoLbvLGez4Edrzb5d
auOmsvAVX3k6tPMDoftHIx3hupCrqPP032CFZKs1cZzCsRWgpjkQ+lUUAdpOGPrN
BgCp5PdAbx726c5/gK2LXqtkMXm3jy+OJ+2fijCtynAHyp8RDaL3xdCv+hzo0FYU
4a3H1jxwS8COkzYk1wECwjKR7CqZB3+8dJX8uF2hJdy1eayeEJKoN4/RgN1rQBPG
bZh2rRoez3aqdV/1kevcb8ER6nQNwTbR8vkR4c19BbsaTElK6ZJAKHG3+vYBPcUn
YhZrzQ69DWXcE82f5Ay/rlKAjPYQ6I5+6D6Kh/s0YbAvnL8Hh1CJwy1X4aaKypiC
REFLrCUqVgiQuIByNzrlA7OEZiOHsFXQkP2EhVL6CxB98+pIyRB921SQFO0H4Uft
KDsKqU7Z4QeDG6aaxf2aqrWAGK9Qk7I/Agoyam6d2Da5X5wcmpKHE17BiuMK34CR
RdQZHhBesMKowg1pI1lElxM4BTk+30Fn9JdCser79lvUNYTmhYqp0cvSA7Ljae/f
V5H6Ps45FlJSrvxsfCuznlpBElNcKnhA7hcev+Yn4Jnte8UFfp4maBdG2obSleTj
Cmt5SoN2lXaBy4bB+Z43n2NbChmL8LvVm1lJwmvGDjHWglw4w46dtIi1AEL0r2kW
O08K9X+3NaL5GKmSv1hY3OKa7V3VW+FG5tXc+Jp7lT2L6uGY+wgJ2gxnCGhYSUjp
NENlEF22evGUXaDb84OtLPjpvyD63fLAhlQ6Z0tlgCzPLoD2QhvNvdasbe58EbaU
JgF9SPNxq/yj/Q2SXFlNTRaP3Q5xQhaOoQIDiO1VMsXo2LHc6x0VCqIZM92oZ5KD
DnjiWKVnyX80+QGJoDAOX9nim8I9tCaGMDQVstqx/KZTnYbl5FFSsj4R3fOr5eBM
jgYcM/lCwkc10msivtRYi7gfjVBBiOt41h5DGg4wZsd659nm6LXXWN65ZjZ2BDrS
3CP8DquTcw5g9ZXbRkY/2A47CdJAQQBDPEbINd/2eIf3gTSt04SQ6i61geR7Wk8/
2qkjLDqvvf3a35EaS8Rv18Km4j8r85ZiMtXsP2aNHty0KVl/uosJZDEcwPOMiXoq
vCou6QWopku7lVN2hyJ3r3i5ywI8XAIcMfI/P6Yb4jU51E5XDW5i1cB9VzbuBPSu
UVowdq8tdjY9LPtEcrDjv4I4zpREI89GJgLM4FdJKR1+UHWo33SXEpSPTM59iy3v
vt/sKIPMd3nBIZp/emntW66+bd9hmkc/uDVt0/0RPUVpZ2gFvyvPTfcULsXKqt49
cix5OfP5qxW5Z7CWeRtF/WYA0OJn4vIZVOjL93x5hjzi3rc4N7uWqHFrgLlyNerU
bZ3hlvtaCx113KWQMfz0Zy2OolF7ksrUhS//SM8FtV7o+mHE/eLIC9WRVDL7SjZP
J7VyG3C4FEY+TyP7UWJH8nVwSDJCkwZ9CxEit+pXOZKnHMUDg6gwC/EPCT2f5ocx
L70EuUBn7cc2IMWs3yR0ciKCVE3H2Nh9W3V1PS8WTLFMr6XckmZ/I8evB7jLv+me
GkuiBDh1H7N1CNdm6TSEa39LR9rnyEgWpg8QaKC/nU2pxKDlxsJ3mWP7IfamEpWq
SknF6gpQeVVQBiv/ZLR/k9MY74bY+KY8hBhyaEAb9/nQ8bj2l6iLDxis/NPV9Tc+
t+hS5FAW6zqvlKScndcWDPX5rJiQmDldiDsRx+N6NVot6BQJIzEtQgMK5z6JIkCC
539L8Us8TED+Dn7GaEz1jZl17104+t+0hPX8WnQfO1OSjc4YEVlQW6uS6PanUwNu
97T9fNevLYvOc5FRUX8L2rMncLvxI5fA5A6m3IQ3k7diXdnDOtZPd84A490kmPzI
M0zW+S2iJWKCb/Ux+W5TF8HNJ49qwaNZOs//Zp+Xaq2gEEKjOIthOdnYARGmJD10
gNJq/nea+ezRegxQCfCSO0xGCqq0ch1tc0pEDE0qM2Yf7KRQWdO3/TpOxVpdiYty
YydMkSMKBAm1QHyeTLOwqyZNo8CX7S3LX+zDN5thQoN2aiLOklMtWuNwBPErq+uw
LVnP8cK/TygiZZhlOuTTKznaV8ykOTi3lKS74IDQe3d3zbnAo84oAgQ3/+fW8p7q
pPxT3U3jTVNYGqirXrLyh9u5sc9OuIb7XV0hL8fyiLhgbUVO4ZqNt6rbCIYVcjnT
plO7syM0thNglT+piuufH/D0uRP9VUU7zLoMqr4Qa1QDDpj4xG2VtTgj0dveR9Uo
zsNpLP6UdOKfCoYRIVi0Q37+axclBhmi9T+68dVRuBeczvEb8SiU3mUF5R0Qcq+m
JuMqEL1MUnRI0cF4fZ1dF6RnVUZUQP0w/itFBU26x26tvQS/2X35dVDfWHohZ2xt
9uV0hgsuyt+rQ5HJX5Qtu0SkrEQ05gePb12kE7bU9vcBa56Udf6QJzTnpFAFxYVI
AJb8MsyScoCTT0JqzMsgAPenUNAjnkt1Emi53KluNwN6JEw1gloN82DAoF8KBUur
dSVBs2VvKowUogBmjjt19sOMJYqm/L2X50VYLARs+pEAD5BSD7g9qfxqA3ImQXb5
YNOWnbYzrmooGj6lYnH1q3wK5ozC8eC/Enxuf0WuB+mglnpsxdlB/J1qdBP19MD4
iLNm7M1qT0QD56XHK228O8RDUX1ngrinM39lacYDJKwWjnUUEFxosx9tAI3SMvUd
CWHtHUBnIIO7WOKCYhotGvfMR1clmUuX4wnmblReS1tfjsziSHvFJVaPKcPS0QY2
2rIz5L4RvsHifQ2EO64CuT+ClBpd9YCuKHj+U5kRLMq/AcZy/7YBC+BAlcK+/e+9
xGUfGPagOrbLIIBUGyIBg60MBkElrOYbfGpgxWFNWbD4vMJS4AzHB/h7Cm/V+dyT
gozLdSSL6TauNCIBNNAAMqNj/ftinrMqLcaYaiJrobqD2w4q1jIWJmQ+BeUXm3hO
GxS//j+nOy7XHhBMQ9ZgdmPawkgrtBUhByEZZqrYL7xRsWb3IsgvOiuzUtxt46Gh
4KLGr/oP9oCq4RqlBaOTfpAC6sXoyVvI64+hfIxW3Wko+VVK0YyQk1eTdZ5oJSbw
PPtAoRSx7gVZEsJMQerd0/5GVMqMnvv+tWRnDZmHWDf04e1RlURTFz/0bONgrkiR
EkcAM7m5zrpHETNG/tbe7xWQoG8fy4OMwKQjI3GC9zgikjgKlmvPgY+IIS5BFcuo
2yQvHB2auksevDObBnSMr04N+YvzTj4L1h4roiiTZB9rdnGFZpkrhN7JVGkus5Bj
GvecU8cQibs1AZgCrr0MlatG9m2iF74tJqPd5lMEeKJ7yNDFhUyih59BEhlFsoQc
+jHgC/6kT4U0TOU3OphVCQGbQHyUAN3DBRMpJhBES9q33I6Bw22RoRDFFoOWZUc8
+pn3xCg81MGMtdo8mwIuYi0PUlFlAWV1O8bykCLZkq5m9jCP0XA3AcVmEIkNjKMX
i7CR0XGMOi9hDoczaU58kS8tpIMm0muHUM+m96G8TjSlOJpgPM/RY4rXEMuM60bh
1XAXPPRyhE8ckp9tOBnyt96TiZJp5PVV4xtOIQhcKWF2+cUERicBr4x61dx0AkSQ
tbcB4f0yIoqTgY3d7O7DP5+H6DUC0Wf03hU7TYJT1eSHyrBq5ktGmNajoaNceLQF
OynTUyRac7j/1+RVSJxptxRN0Nm5QIoGvCn37MjhLH5eFr9Y2EOxY1lGque8S58i
lPQgcg4shau30uQ9+XVn/IrCev3GNO0AQc70j/KS3YaebRjh3TLxWR/rC6veHWtn
ECXQghatI6QORVqxTfttHl5KmX5lATG0heLMnw7jKk4sg9LvS3Kfr5Wi9HbeQ9RK
Mm8bcAY9UrTET3H1lez+uc8YW0mJotJJGkt7d1Pctr2+7KLIcYcWW6KmjmC+AKq1
LimTBNdBX+yUDYmvqk4sxnnXG3XMs41jrmiEChrYsAiAqC1nqveRRE4z/YwpjyQA
7eyhbmdQKlmoYBDoSsXIFtqg9hiKWO5KohSc9V+fa7FL27FztgYTm8KGe5OBCUR6
MccI7UcGEbCvVFQRi/9Ol7sGOBIQdSPHnd/mQWMjqfZg3rjGs+EEVXY5wYl2fVX3
3i8v5ayJ5ZJ/K9UxjMmx91PRm9j12/3ihbisSWThTgyqz6RtW7Wxqif787Q+CSui
is3eIGArUo+z4TjvQDbLdnv2bLof6ddbGODOsLzaVL7v+rX3YZD3tL3r/N528sKB
XDpaH+MRUmyE/qEM0xg1yCVzd24V7dOD0Makc7emJwdyF+uSkS8acjfJ7FAhAuJm
Gxw58zcNusdqwRRSGbHKM6x5EqYADxC+AGZhFJBsy7A0aWCV+M+ZRwAJLGkoI/Jn
OOdUav9r00TzSyxpwQX/nxcMrPuAzMq1omT2PcEVmfJRJIQCO3Qudd1jMq2TyTJx
QQsKlNx38T5ED65zRzfklZrWQuYzRNEJpYylS33pgayqslU+yU7XeyFvr2+3Qx+P
C0tYfdr0/EPXbNX0Tlnmq2uGZ2lHaIE6wbzi3slv9n2Vde5UWq1nV6XBlyF+a0lG
U8SYlruzheG+/XwFKGR6xAec383Zwo4ZMklfrgN1u7OLKsZlZpJ1Arw6J4/jFlG0
XMcVUavZAsXfLZtZGHYqLYQ+0pfbyaStD+cCYfXLMbE8B2lHhNNhGJSy4hjRjnIL
MzXAsO0d5VOX6XlvadwNCqUXECWWmv70maU35Jbf2uhKgSv7nYJTDYI9IB+rh2tc
f9Wrl9For5gZ//ljQ9EO71SqXqgfn/GuCrRhjpeLripnCY9rLxicnua+Cvbv9llA
lwtBzh6lq6bvdIwjIW21OCnze1JtdiC1gCNBDfcaEUYGoi7U6ZGs13COXxCCXjdE
ulqtuYgRxLhQgy9j6rbIlikbTQrxSq7AklEH/aNBQDnGHh2d5Vt65xFzv+J5joES
Q/+RT4PFQa9oe+sSgulnebN501VK/WpL0EM2M+q6Qc/P9IaIYVODs7eK5yjsL7FC
43ds/wVcEiGRXKfQl4lyAVqSdioFVSAemRB3R/+NBZCVJ8nqNofSAlDK/EglHH8W
LZtTdjqe1+q7Tg9+10pCIgg4G8e1XoRheaVTK3muJczEzgQ/kdAslQG5SlOW6n+U
34HzoHp0tIIp2/1nj3Nqf0Npv83/W+SFMLw9E+j3+jMLs27VpOVyf9Sj5AxU/uYj
tGIhfZCR4l5uZXL07MmzwVVcqS2I+MQZOGS1uetLfE4oNT5CplROChd+0MJLVNCQ
AaXtgvnWMCjxCvs5qVlICXv2I0cY6NtpdBSv1hambhblJyGTK+Mt9JPX3WwvYowD
b7I8hrCS35OkkyR5yQDBe+QrxDDlH20iLtv5wP7lfttZORyVp6vgVYaXmt1D4oQl
FhWe9O8f5Gk3FFlE1hEaYr0WLLiXP9Nuf3/OQIwHIqi1BMPH+BFmDiK92uvYA8eb
QOh2LmSkb2xafz5uCEwhj+YgMG+nL6pRO9oa2uxxjX3JgMei21OFkBiDV6lrD8cH
A84zt8S6XBEhPaj2YWSX5ORSmkXi2YJWtd7qGucAV+ZGMmtZAdepYtm5uc2Y7Ou8
wChmNE5iaRG5vwOrszOXXYYIkx8m/5ThwZEHUm4q2E+PI6nrybtUj4DEUwJNdb+n
8QufGrOHnMQ2QH6kncQsscC+EEvzw7kcPvTH5fNtUnq+QLfvjbDcASCIFlxDY/eH
0rArD+qeMxNgYKX2t4dOYkLg8KmxIF9gyP+50d/wUypfZS+OP1BZkL5kLS3cbMnZ
J19e6W9d1WqGHGaR7EPHqP3OUYAuc1gLTH6b1x2qKe9lTKT0G9oDotzJafqvg4A5
YV9pQZ0+/ZHL0R/ZyIHqvgC/cDeQXpakCQ6sQmISWls6U/dKwml8tmD2vFbeY8n1
QtV+bEX9tsYzMPXar+F3bl68b/BUAcH29G+TcV2VRNucb4DlLcfgq48GG1i3vgO1
7yxu12loETfvdkoKvNJ+wIl+B0qHk1nRS6fZBRebQy6QZkVEP53riY7Lw+33QUgz
WWXImRBY4T8TI7oExzUV4ornqHZ+8+10Qi+arBnku8yKcAeYeLWsGwfWQyUXngyw
QyzptLct5k0vUF0KCxWVp9O1E6WKSa4TyZLmJcnssN04DxvJD8GpyEhhtyxp+zb6
G//6q5Yhh8Tvl2V/ncMFAT0ADHkFi4tq8iMM9EQEwU5TrHWUsLXqmWaYsNoO8Gj3
b/3W4S0483ExsEPtq9NZ8oXfxTY4CkOQnW3MFsLCHZF7JXVgTI5Y67OUMxp+76c5
sjYgyufHntA1RPlE39sOJSOaFtXMLLHxIvBP9sToJ60LisQk9WYgfKOAF0j6fiGB
QEoVun9EZoOEuCkjdC5Z5ntz/tPZe4DeT/YQGmR/LV/NacNTc0+TPRam56l4qAiI
HX5KkViC/2rp1ZiBCCVAgNzwcDGGUou0RKRXoBVbnaRFRudBnD2Z+/YegZsqpw+P
u4xR9qeqyZxpAjlGO+C61m44fd0MWpyBCW/LYB/EwxAlEw2AVPTK7nmA2aq9JsFA
pHsajl/gU8fbvsrWy7d/w4VD5sCO6BhEzW71lhmtgkvV3zejE5mgmhIvXxWaNTn/
hP70JxvHjWwCXbza8kXKHtYOgZuE7iVw2syVnJe0/1p9FV5YA1qb4+0dyxi66xpz
2PQyEDm1nNXy8CKq4FNa6HYFCj15Voq5RJn5zKYnQp63lSg8/DOklh2RFXRdHvvs
HiqdTDLXF07QMlpYjM/YXng6maieEW16+7tXXZufxWSzK9YDmJmmONcHsMCl0rG3
pUp6okahHGo71i48p5ZhfaY8RYjK4SeuwPW0rlV9Duat0U1iMQuhtAzIqao4tkao
37/Z/+2rGaba8pxEhJh5wjYl+yoQ8C9OltGVBd/4pA3LMVNsLR0z/hG7KV9GSVgo
Z48LI8jlpEfK+8GY+oIPkOTw7hB8Jh9B8yItWM9lVkrJyU/IPTpsz0KYpdsNZ3vn
F/WfjlvJKQHCRNf6zZbh8KBG78HRg+qvejTD6BQTNgcdUEJz0V9FSJpCH4j2PB4v
oRzvHpUXCQaAcayrQvqBZ3P8qNfiUBDLekrSfaTREWJLF0KLCBnt3Fk24FSbQ96g
/vwxtf+qPaTlUR9jCImcAFUirYVrJTgQ+WIAUBXSaINJ0b7f5i525OqogNikVpr+
ZXhNi1s5Vqh0CfUtxruYTKObLDpTL/k3XtJl7nlpcy2o18yN3Wd9dyLYTV8K4QGb
sNtvAXpnOq2zGtneqYmpDlaKMUunwhiKcBACY1NGTB7mzB3q08HAGPKGsqCfAV9Y
awr7X5tuAf7tMbnYfyBdHO9CRfZwlmr6w2YNgRzMUAdQoBwFx+BoNpUkqFmOHQs8
2uQpr9L2vnFlr/0W3nv9Tv54PYHvjfW5aed5lBJ9NJW56RxZWExcinyN2IyhDoSB
L7La0M0p6D+sL9nXtOKWI7rjbjYI4rFIVq0lCGEucTb7xnfcr+WE+FERoqlbPaGZ
lex8VXOEX27M9EWPQcSuNQ3f/aisr6Yl820LrvuTcvKqvi7IS61SnIPvORjq4rWT
a9wYVejLSzsn1MzH51L/E7ODbJh0ghjp3nUr7QWWIFx14rodp42Sljx3VESYBeV8
7O88KBTRW5Kz8ssV8UX1AaBND+qA8cCfJDMEM/bif0H7ZRoZ6kpjiMi3WpdIHTrN
s7XLrX5sVu1cMQ4KdlHTefopUKZvjwW74maNx0WXBAE0pK6+mUzlrJLzEjq7JfH9
5IoTaaBa+HA6G+qlwot8xb0OElhv1l/f/F2XlrOQjCRh+jzBFWz6m+VxCXxnwOl+
IbpaqobldX26561geVa5fAFkqIYuiOouMbJJQr4gi9NQRF8UBMvsmVuSGACtdN1k
Ms3weO9UHHSIj7MLhT3BUUDg3Z1F6ReEMdL166fth0CcniOv1e17lG2H+jBJAWcL
Ea7kvwrDLvXddS7kL9v5tsnU/amP9nE/yK86PLEiQDL0TLuJ9yYbQTbHC2o/Oabo
GQzs1CpIVeGRbBnwFWStTt2ckjap1WoDI6WZhg7QgzIHrdeMIqBaR2Hq1WB7mwEO
1hWB9cje1pShmf0DCUtn5N2KmfShfJadrPEVlNLAHZUuOcQMwschKQ1vNcJqCQRX
eRqSSpdpa6F7ciKjacf5AYacqsBVBShCeG05xZLle0polxkgqglvmfv8Z91go+Xw
Ou/gOTh/04YqIYn5qUN//pABhArYAb2VMSaYUzoNrUaBMyuEfpC8rsS124Hk4yGz
qCbTG1KPSk6VJlTmO7s0PuMIFKfxsrGDHYK9PBVbovAjdQr1ZuSwD16Eg9penxXe
dkAfkhhjW+w5kTnKf31/FgYPqYPTX062R0w8p2kkuwG8m9P+vcyel4uHzWHCaPPf
TB637f/rbpogPc+/8IZS64eWRfQqYytfL7mpeNMmOjhsD+lLqs6mQeivsOX3P3Oy
4mD13v/lGe1R/lQ/xzBP4G2EvdYoJiNfVdYOSMTzmroqCLQMECdwtaws3pFUZnXx
HuvjfuLKWdRNmjADaaHgajxDbXGZ2r4nZ0hX5uHptHIUEeSdLwzvqH/WMeVHWAHF
edrqwBA0SHY47G05CQHGwedY4GVdvw4AvXf3clwqUFkjdMJGpUH1IKTjyPZONslC
Zno1MzDO/1XppASyZMXtDO2XPxaDQzl0JrPVu+OGU+7HrqpPyD7k412HpiMxFZnt
rP+uEoMh5zkeOOL5J0+h/btqTkJp+t2DTyXVFxCzIdLssQHIrN2/F8loT31hdlaY
vJFYmYH6NYBY6s66sd124g3uBpb5HGnlSBjEBVkEn2/zVJIvwsaRl34U5FHMHy3Z
UfDqLzaPl0Tt0b6VhWdTkSTJt+wUIy+3zNmOTFFnIF8wTI95g0nMS1xYo1khwbJi
NDclH4+2UJngUH8O8NyYmdyeVuKqPhdSVhaiVBgHKJ+lTMRcLCP7ltzwfpj7V79v
A5oCyizAzOfTOF24xIikslfDvWSOf5dcAmCfs/D7ptclVOw0C7IY43Ov/3BZIAB4
UrI8RyjbLVtP+kfSDnodNnGny2VH/tkc/M5+ffaLEjbcOnzCEFKZCOJvbEq+36hV
rSAYKrgq2HYzOyQDXgqaIL0aWKYJsE5PLuo4dVr1wBGZRq6ZgAucWBWF/h/p0Et8
ug3DVZEqXv2VxUtmNT9ZqBAa/sZRBDcj/wy40XX28Ucrhy22qTUuSBUKhNHd2Cjy
AR7XWsmdT5wUpzQsTvzYu7moMM5G9588P3VHLNmxriS4p0ERqNAYun/yTx+It03b
H3TKcNN+eKj8xRDl+Z1gw2RHBrulLa+bIzZunjSe0s4V7H5bRzpt0O5Pnp8Zf2OT
R52Oau48SBD52viqnhBGntUDEy3oIoRYEE9yfbYhJVvP5zpHIeFBRfhZeE0hoPLA
y/0+GYlBzgbhZaGrW7RiKJ2G0LkVOtdHN5Dc3eQ+Xw8tjHFhqPx66Bzx6tmRJxGv
zq3KigvrrW+m3kFcPXOs90B/Yywg5gPADhRREWN55+xNY+JASDLksE3y1I3Wn8yN
TpZQu2xn01mSuPdQV1kgvhFvH4YYKxG5xn2pMZCJpWi9yiHuVHjzczWh8Ft50RWk
5/5N06Vay/hh8eWYLOPild1sSQUSKrfA5JAH8gQZ3IOMNB1pPzVuRuTAxhFVD+tQ
fyblPRWi4zMs0gKc62gAVAHAZfQ4LJ2/uTRzHOzQq8hhi42JfgFMpBS2HQYI6xck
oXzQuyWoW4X79mUEJQaMTEtS1egMKweBxxn5UxHaxzNq8VabE6DuuxkeZVsYJ1RF
O4pjb0EgCVdnHsBDk6G3cbCjFkgSeqMHmedUZkLf5s6xYpyk8v9EPizDi4Ga/tJB
Cxy9PsQKDUJaiwMkBbN5sUJ5T0UV7Nsmu/uOrR/StwmyrtW6nV+iPoANFZRRRIr7
fb+sfpbGRMApHweLL8u+IIi7xWG8eotgRmcmmaJgrZoVb75xLH2ji5Qj4ozIKzGc
tca2qXKHZzRkY9RFCWmL1VcHIAM5967vgoEeYDH/tM/BC68gSRux4p38piL+e7eI
lbIOkPUTdsfr8kc4pmfz8SzXVgZhJJocwZXKOJY3I8bKD+/6LMCF13mMPI3bIHai
jjGb3ouQ5L+dGTM8HN7wKf+QBQgSOyUbGRsfZfDAwjVnQ8ZdICwZzBQp9qx7+ROq
7InFPoBT1Dxld3WvHEEzUDMhRXFEtUY1UT6er/5UH+4prybBcACwgFkEi91qnLLq
BQ36t4pZbiB95PSbVc+K3ACDSv+fWjJ/8a1rcp+F5KNyLsdXj3y9JQmFeMa1mj4M
fzg344FT8qgEgfNG+MvL6Wlr90QfG+1nkHV4rkNKhAqxTnOd5d+vGqY5C2TQ0v0y
Sy6BQQb1azZyN4+IV46DBzCoOaKR257jmhhal2vYd6GA8PSC3QrUv3bInFOKgsb7
IrH4xkvpKD0m3MNHNLy3aXiQ++m60Hp05zbqJQ+LudPhohOwrhdYPiBjtxUOs2AP
EqhJv1diszb4NefgB85HVSc4VLOkc73Q9iUTk1jh8nffOvBkb9EA44YHwxs8ZciF
2+VGAXj7LIab8TRX1wITQ4PC7fohMjMqUMW83y1XN+vTArvf3iAJCO5EwgVxyIGo
sMcFWelFGZMBHBxjLrEojQbNkxlBIvB+HcQ8dCFaFAnsfNeZxSoHrM6g1zXrVQo6
A/1YFRgQfb/RfGQqGOPGg5RAaUoK+ZDa6NugtWUimCR9EWpl8dGgYDO7Shw/Qf9K
vnzy5fbpJrOp96QqIi88bREYeWYDXObGu+813EWH4o7dtlV7i73jGENkzYXswymj
JJzuD8gJ02AwNTI3yaxenWh6HsozbVfY8FY6OdUOczeMKdx6f19jL3W4FMp+FaJZ
WayIQ+dOq1QrdLCc8qrLGa1B1L3SE4nxAm6OB/Nap++z2vd84sH/mbXR5EvgIZMV
DdD5V7jKuCB0fK4Af31uyd4JGt69lSPQWm7pcqRUEzDMpY6iXzraJ/gkGcOP96IQ
0cF/HpHg947ydI0J+payoQbGLKmpio63tkqPx0huay3SRxn3gjAs/mqihfjYC7Gr
u+6VJHmXC1AMUsMU8XJkFLR/SVua9jANe3FeepJpRvMVqGIKpdmBJb/0eOFQmS3V
fXrRoUmiafuO+WjZNxYpsgdFq0qZXDk5ztVAe9l4iYPvGP7dvQfPLKujM9WJ9tSj
dkll3pPlSPWYwO2LdXJbGKcw30eL8029SJMaPmJk21vK0ztcCyOxs9bsQ3dzU9fz
wvr43vj8lZfFL7GAjv1aZWYmOfX4Ox8uyfSBw0168Bx+h3jwNvYVtpBiffrLYLQG
losths300bnm7CllTSHdoAtCgf5Zk0Y86zrYa1+adL8066wt82UesrkJxi5mYdMu
lQsuig/HjMWAexdsOvKYt/9uCn9TT6UfCTsniSoC37UcmJqVT3wofKw6Z0tUXTmA
swMuvDStP57Mttj7NCfKoB49uccboRifZsai+SUJR+sB6Vk6tvRM0WJWciIFUYHu
ME9ztKsxvFNtHjBFgk2rHN/hfKXqbnsm0JeUnP3N5gR6M/jcJWtrIvas+XcKIsGm
Uu4Jmxn8noHzknjBKhdFTThg+FNfSMM9gYVenhYidc5CuSECYljvYPzT0FuU70Kb
KtdmytuLAhEuKV5bMOm6fSB+0ibF6Ht1xXnePIWOtVV0fZi0nvwQ35J2xZZ0IGsY
yGQweOrmZH3EHi7EObFqSb+fvfUqnoHBYehUOxgVObYmlKtEKkdDaDqp/mozuLDP
YJsZhpvuGuyamPFUE+9Xzlh1YH5Eov6eo9hk8iZkHLUpPDyIRSWPHvFtVXC/t1ms
ce7p8V/7VroZMTT0/xGimpX+/WyLn0/0A2G+Ib+iG2wRHR6XxBTGIgDlfHiAHKeR
DAMKE0qLzU1eKsnoLfqqjs4fXOMa6YYAPCt0599KZJpeYJwSWy/cOXow+NVNDEQ2
Dg/aF+87J9lD5/Qk+1jhM0DqfXE4sYUbMRA8nPnTHLEGGKHNwlqMQV5m2wgg29Vy
RcM0xuxF+Uo7W587j94qD1dMx2x6y9kZh+N4bGmGyGCZoKiIcXK+RmZIyzGtt6NV
YqIVexVG18CZw2tZvXseKeT9cfRrjA2WHnkdYcu6YPByf+l2cFnhFFhht2RdCGtA
J6N9zMvH5yyybI0T23nWqMW5nVsLdU/TjEWF/aWS4drPmKvrlgXl0X1orM3NrgJ9
ll+gkB2jtlMz9NpzJHhefvldDVNgHZV+vCfJ29DcwKLKv9JJi7Z1KTGUu2H+m9f6
7Kq8NiL1QTRv9d6Cjai6vEl7FGKbB5PqNlFZ6pBmpTeJLw/cvRaFzR5iEIPYmu0w
xMdVQWYIyHhStv+yfVxkJ6vCvvXl9Tf6XzsK87xbPYEFJ27ZYWlUmuAdJsfZiZTD
i95swJQMsxmEe3lg+ZaNFCs4IEuzP7GBWLQEn1k+/4w2pbzttbs7+xLUj6RZZ5bp
AGnApsP67oFUz+iynDsnxW0+0iqfnpzgmsSQQjJj+1Xja9bcdBzCo+yLvhz/MsA6
h6VuTtWVk8DqTe6V0idxFJUc18UH+/cKIwDffuOnlARWUMMGgcap0R1Z5wy8FDyE
R9MicWpMAiW/1KSsD+UN/+mRDfTSSl0h+Nu+KP782ssGnIQtHA3ZeAxZkCtZIcH7
viDbA1rti/q7ln/hZlHH6MDl7AenmGAxdERUAP75NeJM2sFpmTd5N+RInmzpnuEN
WoO9VQJsDoOCGeED+EtOodTzIXPHzTNtxWyvjk6ku3zZSlurvvQWKgTfGjQpwd59
8Q+Jm4RopzAeV55Lq7qjeN4HOl4HyKV3/p9xGsoAzn0I6Ihn+HtKcicG0rByXqOW
2WzYPMWllQv+JFQdXv8gEYapPRP51jgeUgJtEJ8XGEbUB6icGxMWQYChe4Ns7E3N
+oLa3cUTJ2PUPceAqfdGofAWUyfj1EfJlnVlNF91Ao6la1oM5bGApzIcgMaJK5xu
zwsHKgWNHblhH18CXXx+UskumrWfn0gGGuVRqRZjBshff654ZEkgUDToqN9IxhSA
TP5FfvBg0auIoLQnn0T6EP6XTHKcmOjB2nuyA/WOydZTtGDnpeHGXyIhTT2ngIyP
bj1oO8d6kvQIpsCWkk9Ew1u7XlhPY5KqFHSSFfbcU0a7ECbahHnGVmerZ6/bHDk1
OOhhxEk6sMk9+YPAnbnlVtJ0wSvJEVwaEkHApVuOlkLJTdTh1vMX9qqG1CHF1xrG
o1jP0qh5NxTAioJHc8mz+0YHvQq+bC3XmKih0/zQVlHXK+jQZzqZlCzEx3BMm7TS
yn4lFn1msTeJqy9JYAhQlXVR+SCuLf/01mbi5lJfMmNJgodyWCL2E7Xdu/Hq+9UQ
L1jMsK36RHAp2OPucLa/dg57ptdkGybftco7HbLI9FpvNC5RQqtX/3/H2Sw3FpUa
zXkwo0w43p3THey3LLAsxMYaCSwsHJplr71uvIb5kvOKRoIiZkmZZJJ4drQBdfG+
dFp5S9DjQ2ABGwV4Auyl36bYNJrPXdm0Jw0mRo9yV8VfltQ7RJ74shrtzHQQEbzs
WEDMB01kb0PixMTHckmrX4Q3BEGcR4d4y8ruTdo9MbQipDe59K0o3AEVqitkBJDT
GNbgcogPUDz9zm2RAC0BKxYmHP8mqBt1p0/TPcvUbhVviIzynpuXsQcxfPZd2PND
rFQVeogJGl7DyhibNWqVg/w5e4O1AHAOE9hkfDulM4ipdDeOPSJSnryotLBaGAzU
yo3jbLp06i+6Vv1SKEIoIHPh//BSQovSyROpKRVdb3eFAsLzutFxoB+QOR2QpAG9
04AYre6WBezPvuEDZhZSsxKyVQUg1RJ0l+ZuIna84sQq+MCzEcl9+GkUAwFWXsRu
BgUlpjVUSR/8/cPtY/AE3Y03BUgfgaDbigc/b8V96OTo4L0jwPu0RRKgNPuHcas+
GYYJnE/vDPWRXqsrkFouvx6eTHM57+0ofg2TAqnr9FQBhHXkb0sW1BVtlaZk8wSe
CjH+0VXmxMn1AzH4Vjx1iemKS2Wkf4l6x4SwjOvkb0G+/1hHbv/Q4m5nh4nuE0Ym
cbw6IKMrTazzZRUaA1IOWU60ES9cs7Nj3D8F1M8Et8MV/vbJl4hspjdWK+Sz4IBu
6Nt9EuJ4Fl7pGH6H+OvZuTB2HT2uXoskNyHYJCdiyL0Zyb7HorkcZFbMiehrTpEJ
4RQ0/dFRNgAjRABDbZ7z6crr2roMQwG7dQ4KHFHSBlReaJBZLRWdEXkNA+WOkFj9
u7YAcafBlA70PR9XHxqllFh7RaF3mrFMU2Ke6d0hfNnl3x2ygoGH0XBROYKWLnI6
PUGr1Tr9E5QMXo8HU+qErIP86M6OQs5vcK5eMOviZsiRZRlD2EOmGK3jfwt/m0P0
crJBTqVwf/BaR/u0mY29MuZK3v/wEngo0K53AnzVJpvWIy0bicWX8Xpikw3L5nTh
73vgyZ4NTEzdKU5KlK5jQSJDBADskFcQ3cSIglLukaONgExIj0tDm4zZtBo4BXGp
cY1T7n3ZoZnLQ+BlkcyKET4GTVXqod17s7/LUwsbI6fkGICD0fPsO5YQGXEcOFJ7
WFQ+XelWg3VyXjv9IjIHicxl1oarhEa8SJioz2AjqiHFO9mQEeiUchqdOMXclDcZ
MzzdMYFs/8HpZiiQ2eNjrxqAnhxZY9zEe8N7U7qMk/9dAaNLvP4Tz47iHkFnp9RL
Q9ApNATdDaLnv2nM6vrDnrSTj4kpQCg+yZ4NDcNqSiuAuwiZpzDYPuZ0TQ1dGw4W
1wOduFX1wFe8XZhIUjzM+us5iqPs74AKb6h6ftLiqZJpd2LL1p2b0olaD0/uESn5
bwmUB43Xlv7LcZmMXyO9TS+xLoF8EyN0vXL/AJFTkPEEkQmqdtNSdwFKUqwP9BVO
wsWkNrw9EeBw937zi6k/r5eBGTMYNZDqf9VcWs7V1iZ33bSiwLrEBZGm38NddBzM
cnmhXYwFz4nYa934y/A195/Gi+BJsVNj9fdwnAXA2zOTR4XAON2AqItGIdbcQzUA
0+4jpS2V0CAZ77aSb/S9eX8N9WbbWVLF80fJsucl18Mjt3O122HERT3LykWISTTa
nDSpygMftjbQT2g+yWtBGFAjfMW+bBBAGGRKGKOrCKebSwDZlqImiMGH94umWi83
ELzr4EjDpiEUsTopN3TAYi+2hl62eZmwyXsZg4vdv+/08zzdAQM01jB/2BVxsRug
H3UUpZMEc0wFuWXavPI8LI7DlLEUpwoluf2C5O4aHrjFkWtyaiZ45PJhU7E6MeWD
rZqDdTU4ItpJTILWg+jOSfIKO0Eum7T/T9FxBaOr9sQvaUTsOU/fHT/Hq0bWBUkd
lOwtEYrj4wbjg5GSNqqI6P2M4Us+BvyCjlKYwJn8yX0Awn4BJbBazI5pTRCph2d1
1I268JxEcRB07D1TfnnOJwghf1mfIdId7boifsXkpzW3zHKca+wxud0hToN6aHDZ
r6wwZ8xwMy7A8RV6MZ7sVPMAou0LVM2h9iFSI3C7LzOTT2GG8dNLFERPgyyks0EP
q3rNbJ8CRJ2RyViNoCWfMG2zIZFCDfh8TPqPrpISJrNk5dGyDuNaUOuOjMx4hx7Q
/MZgFM83HzEUxe4St6PtXWv+4ZGECUHU0aCo/o7xqGYg8JleVtlcWDuSwo6JEBWI
7rMFVZFYtzFL6iB5/nsKqJO29HXCmHk0rcYHrUJs2EjK6mLUpFdz+f0y+rcUBPo+
LGFLBP8BQFlhKsUmBTILCIO654EQVCuBEZwpGhpuxQMEnXTFrD5aFcrCrFuf1/jD
jH4pD02FVkZ2IVsbk/IasZsfX8hiBoLwRwBVrJUgfDA32t7gCi76IjhaZaOt9jZt
vg2sRy0aEJ07nnrZa7gnOUGCwcMrlN3WCtoK25EH0o8V0eVs4YLs+E/KGGCLqI4A
e6X2DmyNdaLck6CLxuzC3nWNt+2Crl6cNQVE/oWVthTYyp66K/FhRs2jLCBOIrf2
F86lyiym8BjNnUmhc1atxwGmkD2GkmhuRzN0dvzNVd0pQFxpGSqf+mWwUrkoUs4z
yEZ8/7vMw305WnltMpXCbSy3eGyiqW02tbENqhIjemqMgPGfUzl0NzQZNId53KKY
Y0BkKir8sEp/p13L/YZsi7LUWondWicRCiMHpr1SQTgQ+n8mbySz9cvCuae5sdSh
2rN5EhnzA8qMJps3QWJaY45h+KDwdAVmhDdIj7G5MIt4/rRODnQoNAoixVNjhaCc
o1+9FjscB2zyPvZT1DhdtvKNybRjSBOZGcc4loclE6ixYgEjy9dwigM5JbbWf51G
PCNB1E5riVeNFTXQUQxQq33pHuhiPkonf0cIRrWJymBicBqnWcuowTMg4CsTObbo
wgnf23e0JyuU6KHHB+bSpdCbl4DVDThPPVTGU3QFfxFGKAqQOppYHVpk6by00ExN
2coY/mARlRXpwqv75tr0dtTAO3evaQfjkadPAyan3YkDb+Vw4lu5AJMRwUoFlhAd
7xEvo1PjVowg/0OVrth+PwEx/dpdIrWS1LtOXVk1Vwp+00iZOPeGs67epsdj1puo
910nvEiaG2whA1yp0PyjVKijgZA+lqRQYegrYfIfU3YIjE3H31U+Z8QobT7cFfKI
ZUw2fJ/1+29tAd6s7MM82/PFjNQiOtLJReNv9cB4/Rb1/xDdPjXWBNnupaRv4f4w
SpeFC4HfFCKUyuM63gMlXdXUoQvD6Pg+O06t6mRpvP94tnrbf1tHHwKPA6l7r0kz
gPavTvs/TB0WJrUGVUmBIWRlsk15EZrwHAipD6TYJMD5IP7e+GyC33khTXVUZn0p
Qwdy3Z2uxDH/o97CUrkJVzOrOPKkKj6KnpYu5UJSmVuK13htx8ptopkUnxOApbZs
0sQeZh85ZHEOypN9HdMRVT/uxtCSHxy8oIoF2Ohk6VfcvnWbePvyDuCgF+/OL/wY
ecXZRmqLiOJJT8NGSVO4vqCpg1CWjjL/4M42jsCtbkj5QzoKrLJIb11nR/1QqS0X
A2UGLaN1fLi2aVz4neeC/g3CAZpm6PriHSVD88n2SlzGKSR10GhsjyBB9YE86U0g
4C+1b0vC41DLG96gyineoXmGaudCqKL98kr1BTZUSNWUSojuXdW+77ywvqO/nCDj
f/LguxY4HIaqTW/992EoFqR1lSzo5NvarMJQreEgiBXr5O49dqfwTcZXW06gTzfA
poirKkAxJowPqOS/M1S8f8f8SepUZ1q2rx3cIpirzLiaIosHVXC8r+NLmMIbKj4T
mocSl0ESP1PFsS5UHs1srq3w954sF8rnSn5WLHYJJNDVl1EiJDzfuHBxJg5fgzm9
qT3W9jTOVQMvPVRT9XfOl6FZ1x4b1Lh0ECwFAANgePlWNMSxad+1P2pDxUYNl+nV
85W2yZI0gM0QQ/gKugo0o5lZrqLJC7UreXcLJyyKEzSKof4uXRcq3SJNPRApcYqR
et0+7sdRwFJhd6ZUTGQQKxjsP2td4/BWwCOcRhIauE0Hx+Gqxaz33V2gzYYvOCOs
zBOz3tQDlf1eKncFwFxpjkhDdvjZGpk3LTjFVmpI1JVI9fYaoyRxwTdNzZTaZ88t
kWxZz881e+nF4NINuHUezVFnWu8ojkl2u6cdNGa5p28dsy2cdc+aFcY/OGpub5Ns
/MO9F5fCUQl97dcgOz9fh+nMIjSVK1Z1+9FubZDMQ1JaqTmyJWTPV7XDLhF1IJ0h
5Ra1rVgp6nOE00N1AZZtPYNEcD6CN2rvgtqP7z7ZjpupO3mx4AUtGOYS7VkM5+BU
90CFMULgud1TkVRkHYvSaq15pGvbO27rt74Vb1udteM+GBez4heRJ3nMT5v1Zif2
jHqjN58d50Xx9rFpPVnwhh2RfEDHsewtqaGzpDrarYsqNlX5FulWdxGEn8u8CsqQ
6cWu8s5laHi5M2Hkbn6FiVdAVK5qjdpLA2muUXdpqWBiJvPfCBXcGBunDbMqVWiG
Ftl1HqzO6WlI/CLJH03Xx8z5GYJm2OM3sB1gEcqrY95Y7F+Uu2APDPvjUxJDuA4q
O3u6PJ9QCvpKabAh4oKjFbBKSOvwp+e6O8noV2Jm6HBIgd2zJpuxFQosY6L7cEIA
EXMxxgxg5M12B1S63K6KF60U3+MLvsu1wv0uNIZemZSerQJKewd0Mqy413bSyuiU
o6xAB6/96YLZQ8sESUwBs176+K0+0iAHltvii5WBFkZaIvrI5kUFvVlXS/viBLQw
fCwAaCZIJJT/fWJoqGEn28SYGD0YZrBH8gp1SfywIQdylwo+lrN8ixnn2zMXUCFu
MYFweiCXm76W6KnoyjxgiFU7Y6qXg9cZO9QkMC7KLyWIfYrHrd31f4mca553FOwD
yEHiSdLDkGTPjwiTz4pN+OEhALO+Gsedy6uM4LED5sKSwMh2OZ5XQj4qexDYlyhr
AGoiTBECjjnvK6vnuy8qeNNxmA1ZGsmCU5pFfU6f1vbybJolPRWGi1SW0HkZJKih
kEhwMyh9K3s+P5zDDdk+/7Ljcn6rTHN6v15+h839pT6a7TUeoq4ydswAwf/5b46i
T8xHb4SsIRnyX0tVht4d+orJ51FSRSfA2KRNgKiMWWFKDfR4WA+6TuxegCL/MRg/
1bvZJcOzjBCy49loRNvK2/+KVErhK3ZVTlhkke4YOCumSfcDpFjku5jL0v2kQH9G
HtLGvDF3VLg7ZTz7TjO0SmnV/iGDHFX8lydPNtyR3BYJrJVpyYZNYIW/fvQbbxUt
3XcxpeY554Ztw0TWJoFAfe8utJ625T8uCglvYGGd/CE//OnQD+qzuxJj0ZGO8TxI
HM+ZA6YH2RQu7HVgxZjaqFL/AXFZ23Ws5HB7AoWACobdC/okoqaSji9/FZRnsCI1
CQ9rD1dYeZn7edEdnF1lOPPSSgA4qtiFzzq82CRXWmPxrc4eAzjIAwITtnPTuRHM
WYTAcbaiEfMxotmNu1GvUCfLQkZQTBpT7GZ3+MgyB+XlPMA0SVxgDG1afnhbSbkA
yJhpB2jICCLd2fOSTVYVXt5sP31Ir75KflQOdtNAz5t+AJUc7ikI8GYpPatkaSxO
AdyBgJaTHMdYfTXAne+GR4cUSVbJCRETfQCwl0oQ1zz2NqbvHPCWvdUG14NCz+MC
CMXkiI2i61ntO4+6nPk4UOdmxb3xoVhaFlcSeYm/lvkNTgzEHp4QMoFfaHsP+M7R
imveaIj12o7/o8w0GOlJbRd0rAVvbxWtnodqiyncoBhprO6dHi5K54t/mRp1ksR7
Hoc8XdFP/8zynmNVnzJ8bQM7IKrSCS0h7iUpwOAaqpyOCtyJUOMsOKaKCDoD08Ui
V6TYvr4CytZM6Wa2/NQPz3v6JJrbwEKXIorEotIH8Ahxhv4bSYekLc/bJHcnYCA7
cFGMjkJLZ3dKfy5Hah0ZNJvOJwnRrhlw1fBspRYTZ71OlLEPPfRDCBHPq4kfUEng
IIVI9TEfUxtFzWRIXxnSvt1mZ+ePEe3OkyCdcP5cqVbv0VPRFu0V+y0nDebjiFNw
jF7Gq2/05BpvOljvJv0NYHl8mS7TxJKjIaTgNDmz7yjbQHgER37dwENa+M93nxtV
CYP/H0vTqcIKyIW2mVwtNIGh+d9VK6Pw4KNsGDHZK+4X5vJt/0GVoShB50ZEZO2A
OtoQR76j5O6ctY7z13W8rmU15RaWVxGAlwBa6jtiySoL4Nc/8V0DpthO9l2n7q2g
Fx+l31Fuk+SIVWmvgOAo9K1W11FmHgGzxjogIPehpTWwXQP7xf0kqMn+h5IiFAis
zuixt9v2hAs4CEmNRxvDPBiUJ0ecIDyJI6MnNn1edzXCunjDcoG6zGGPvLVQhBjx
RcuMm6ZKZoUeTX/h0S1OoU8eiCpSVe05kFEFWEMf1r4dYHQAORyAR7fIoDxCS73b
Y03FBAkMPU1S3eLSbkdg9ld9au/tVEJwUTz07CUREtD0rqRzBfeQr36eAqPFhHd+
a7WtBkcILvwbEXHetqfYJMaGE2o6+QjV8hcc6L7zNxeUmlE+hFEA0wI8Fc56UO5p
kC+29UuJLSdisuxo0189XQQMhFANdqt8mA74jSldttmISyZxhJeLGK8lJjKWUUb3
wC6R3DfruA7iiSrrv1K7f3ZtDT+Uv2e2HBqhpytJqbcTLRttt5pzkCXZfoncXYC1
Dkamj8hyqRo8EuaTo/rIt92nhxm2OkHvzKlke7v9epdDUHRlbAx4vzOfZ5dIODwD
QMEqylem8Iop6nNAKbfkrRm0/o6x65fkQyZwKdl3+uH8A6JJ61fBy5M2/2nm2npi
GFD9PacUoWrMBVkgqjoxF9IrLUQbFm817DgylHt9jAuzbYEmMZB7j2g5ycdqqT8m
uamZtPzOEqcPa9dKXF7NCvbS2yuUvvz7ipQcGrrZ3QBEhtnV2o5ZuBQbixaEXKNH
saKNSaS0G3n7z5+Q4zQyZZtrY+VF4UP8yxffFgdhiBnvCYW7U2+ej0sml7yUbHo+
nyyn5qUzxa+oT02EiyXTNaH+MpGWFgj+mxlvMKKnR3OwclF80iy4VwGrqF/7iVct
A4R3uf8QZdCBRc9VBCqL5hoLhSqOpuReocVjB4QCR4//FgkWictCmL/i5Z5Fzzqn
HnU8YmAnnhaJL3BFZbFioLK/WHAG/dw158jLyEhyy1YbE6x+IrfJICU14z8ihnKn
Ej6nh+hETopWuDdC4qEJt30rETWAQ3ANnxmwOlq1w1mZ6HmGj7UFkEesBqYuuhTI
sCwnvw78iRAmeFU/WSdUW9OItBcld0Uq8LN/xhQM1EM3hRUjKPHtRFlHpjgeqX93
jgd873j6qC4QKLl/IIBh/MowARXn7ttLWosMsJZCuc3A3sj8Kj4Fe8NSKFKv46Xw
SUv3HvHa7j/hHQ1u0dZQYmyX0qO1fuYB+5QDwBr7h0iDHJkaE4DkNp1wmrdSKzEa
OeXgRM8mU6Bpr9y/l5BiFXtuFask7FCQwdoImMjvO5GgN+RlBBS/eICQXLQDDAue
WbTlGD1RmTqb6zfbtj+UTwK0sSyzaOGdcNTzqXH4OdcqYZd3/IqKInsYzbQNdsSI
XLhsaMPxnRDOM4IXy6j1+saC7Dp2EC9bpYycNXqC+3a6KFfYuX6AjcH8OZjHINSW
mThl4Rrjv2hBIhoOOZujYkCo7AFfV/8PSBSd3Y4PvDCZ4wQwyaGwys5iDKE4kMs/
LCZeMiMH3EnHnow+YhjbK6LnZQQZTUjNrZufOV58afk/G0kz0SkaVB7lPzleVQjv
cTMRXeN08ft5T0QboEZA1p9lmyXOizmn0t/L5dakcHHxmERFZ44BJhbr8pUQuTMm
EZm9r44/x/+0Jw9Ithn6hW9lU45udAuh/lapCU3fgUNn8svz3eEEd0Zvzb+G/fdp
Sqwxm21M18+8AUPNG/vFSyZJyZ1AW4S31Yw2V/GZVOJypWI/NJUjx8eyCYLC71X4
DrTBpuBfiJCWWM+zMe0ihS7crKSrMPkmo6sxoFelGtJs3Vl/hbY3DMet0+P2fUvH
g20pRQFkdCpztfsOlHc2AncuN7zpxbH6aRTDnruEUgW7APgVsEvx1sjrfGH5tuz4
++57Pe5unHTCUAU9wU0+gvplv+9RC6TUiUN1Vh8VS35pAVMG98SXvy4Zat4Rjk1k
u//Asrr7eSeuzI1Koue/90j+eDSQnN5Lcexi7nfNAnma2xzoVe5j6YO8y7WLVv6J
3vDa37FtZp8XOuIcKmNzx793yTLWVWr847USImT6y3V7tMqZADqmrBQRv1RMKubJ
RzYst3B13NzN0ct0ZBJe+LDWAbaSO25qC4X5hY1kXV/MOeLl1hjqemdegQ+WwKC8
acA57kpOG44kpEKKGKHtihB0ZCvtYns1+GlwhIjViP65UxZjZ/ezYGjG/cWcBxn5
Op8Lr2RS7dCdtKmQgglZmKwt6cUcpz+/o4YkC404MeutV5OjLXn4Q4yKpFadu47G
2prZHCxOBrMid7G48cDhQSQ+2SNRzj2By8zR/5o72Lgw3d+5n4Uf4GC3W8j5DRBm
oL3CR/NAaxvGN52q2ioFZIRIdeH3qIzI8wgfRFyxs7WrZv/FOrWQoOtzYkRGoLF8
aSnkuiXpBiNXoemqhSu84HV6QbWImIkUhb9GYsT+iRyymB4NlTWSrfAQyopIvphu
O0Jy0P6iQny5KGecp9+1T4pAiT2xhD8uSVquIwoTO3KUpkzqX1WisfIREUDxTGUq
cuNt1piMuc02M7XS5E53OqWrTIiy8PvZGuWodeV1cIVAktFlR/1y4tvN+qeNqh70
s3GhrMTk3dqKfWmlVS5KJ4SOz8HWY0uS7yvjJTApIImRCz6QnHLJSekowPLfnnEy
QLT8/K3WUal5dl8Ej/BXx0c06NbYtNDwCH6/qWC8NrJLwL58LdxwCMbJtnMGiG1g
mAVbGUbi3V9MaiIjMJQxMMTeUAX9KwE930WeG6mw1k37FCF5SigoZdTann2QdXu6
LwLWTr7e/K51Qnb+KDrZpoMQoTkJPQOm/kL5vYJkm+jnCaH5jd4gCwlOHDLiKBji
eiKYzZhS7AiOp5OtWArz+at3xmmkZDtaWy2NvQbfakfqBxIE6JoES7u+j6I22kMS
vSDrQzYQ3pJi/h6dcFg8dJ3y/2h/pK758KY4oEnRTn2o4n3+vDgpzM4hR25AK2Am
TS/1vbIXL09XR5ZyTyzdXJARLDxSuT4/c9C77ApkoDOh9eGcoyLc+ICkBnHg4DE0
2SC7sf6esEK2SQVGfvWKCBgxcrYXyA7rlFfL9zHXTBEzb2gAEaSaQ/kxiKu/5J8O
Go9acjQq3f2REhlzswkrTy496mETzHdPa1MTZyOtHFywVbwQ5hxD8CSu2GMcHbGT
RYXOIq9Z8ZKRHbKrLEPUsT7RRocz3fnEPok/MiRbKvQp3wdkdspQCYFaKNNzxVfO
4FngZA4O9SYzqJ4HW5dPbfd0HQJamwIjUruP23A0Z+mKJiuelfXcGaUi/dsQ2Lm3
ZPn3jZnALfoNbc3YPKT97qj4YdaFf0MCjtkHAMOWrsZ56cW+E0AiYmjRuO181SyD
T/kKV5Puljo+P4+6+yd657DKS3GdJTW+rvjbe4a3gidwCyJM+9hgjOPD4jBS9rsy
dKv7MaKHu9wN4uyUoxyhm18zgEaYSp73x95fH3AJUBWcHXXJx2STg/+kaZ0nQ3RU
1cldECsLlYlUu92/q8CxqA1d1POw44rnkayRWLAK11CXi1845mJ2ND3yNDvGGavq
F0uexmFDAaFRhNdr0U0sCzBXlGl1Vy4lwPNBOi/P+bA52VWmobE5yuUbydsMqb7b
cGT9HOf6OmiOpN6DWGgAs7xobTIwvCP05kheg9WaMtl0pXYRdHVYxAojXP4WwP1d
Q+Th89h/TLERPFAsuXghEst2DGLiKs4LBywzlCPfBGJMPABHPQyxEkv6I5YIyu+b
pzj0ZpFYnVdMtQOnrE/ez+gyb/qGuk9TJj0zqIKjD9hiTy8BuKzYWKeVVm0k6J78
HCrZQC47hG8Yus50szDBXxOTwXpQfzJah9IrB7oCTre9BoGMd7WNXo4h2CWbSD4x
HD0qf7K/NR4f5IKllw/HjfqAIg9QRpMcSgjk1wlE7GKlOwdx+kpEp1z166Lj+trD
EhRbNdpkSH7wY5GJAZktidr/RHjYIpaa5V+La8WmDfiUkN9eGJKoTKHUIZKscbIi
sfna54Sz39poXQbL0vUDLxWd6zgQa9gDPtCNPGZWBgBN3xGhDTPFUMA9w7Oh/1Qc
2Ucknwi9g4NICP6Vucs0XQrGQW//7hCN2x2BvYJUpCDZijejKuXZNlIl9sYY7Ery
3WXgKEHVV91BX80G12Y7nUaDsjOc1Jdv5Mt/c5zh54gm4sOV1vv1CY0yUotUzCFe
87SiEFVJcIn5RsEz0cfKnA7Xajb8wcz0XB1p1Z9DkLI/G8FYTSZ5I6srbErZRggd
/KTOy46tP1wvj6OGfv/3mOK1QiQQXDN/ApbhH1qc72EKf6fI5lN3wuscE3mc9ADQ
kyWYrAKedNKwdvpv4/bm27dK45ix2W4z1jMmfpzSFRq8p8O/im1GMbjsxK/afF9E
25pz5ybxHf2eglwifGcX03ZkiXtqf0jZ5kIM6vekd4nu31WqO8pLUXyH7vrcwZGE
2i8YAu4cHvdK9dfRn9e86tdmeOg1agMXO32vdo3EORrygVHVhyO4d5gZ/YcCouUJ
l7+67HfcLNosv0DbJWLs0k4eXnzNClUYCS25x+TbHpTYWT6aF2vAvn4212FtLM1p
rvDeiYHkhjc99A2rW+mmhr6RfmK7nXu1uVXEAXAN1wmvYW/cercecbS91/ZwfV84
ZYolfmgwYCY9I0exfv99+o7836XU1Ilek76r9QMeBwAUG5xZ1GCf0YOmNZY/Bap7
KeL/5O7MBTqbm3lrmHJouJllJ5CPS2wEnDOgXa6z5EGfOvayjC2Lzoyj2fL719Pl
RHim3MToCP0X3wjPC96tRhGN6hDpe4B3NMOlwZ7fQMN6CSUCFfkaBIibm0BtatAb
v6iOQ8BUSn+VRmjQtQk1kI59IuWRXi7oQdnd7DAurRQ0qcnViqcGI+4uT9y0g4pC
6K2PfU80aeM8yCzMewtr/U6MGnJUvaMZNJEZp+lk80PgHk92ugKKcGiw0Z2F5nTp
7mzI+ucPpLNncq1dGRC30UBeKpCxi60+y8OA5LrKWPz9tVR7++GSBEnrIHatDweK
VW9JcGdKVqlk+49w4j156YgDvitYu/luC1S2GwL+GHELcbk++FYuond7Y0yl+aWi
X34SWjjZZkJSHbbUTbozQy9OuMc/xPDHGdnF1uTrpk8PJ7VBsdK3xC22YntLpZg0
Y2OdDkbP9Rly1BYx7TAsJLhmTbyRju5hkbIA2+t0V6mfF7elvOYi0z9wwxt61wvT
6ENMqGgN0dChLxtaJjkWhQ5VykurR/iTaavOQYb2QbZDEQISEOFvudfH9vJJXoC7
Z/wEE22H189w8uexZhZNg+iBk1bfNFPC+Ci6CqzBL3cLVPcRLqit6+iESWpLfExb
x2TnA/zu/HC0hFEuF+J9npwWDs08ubjzW8phIQC0wAJCBmgJWnJRE5r+HPYhCK2B
WYUlG42Vb2YtRtHW4gbjcGtT+0veRxCXYx/gq0mnnHm4VAPwnqCfKLQeXCFPSfBS
GrOs9GR8YtP18rMPabr82XUZKpp0bYhycoik06vrkQNqiuRuhDbZVii38Jnn/DmB
MXA8Y4bC6V7x2+aItXKavrHV4Fr8fFLg+YpyC7eLNFD/IIDcIAvMA5F1/1bhgeJU
7IY2fRGxVGJgmPEYknenB7uXiAX5AX1ZZHhkqqPwOZmScZGTO+gwa4aNLkmCE/LD
qa2KRUZGppjQIGQde8R2SJSK7FuHLftw0hHqJncPnxeiose6iKrjlgLUGSqbZeZd
DoUk2kc87p6J5KV12z/96MfmruUlaCdrttFq7dxI4odwi6nhjr9BJUGjcAcQJR6v
ELcUzHPaVrkbT5i1UUU9eKr5vZTEI034vBvW9s8y3fe5ie8NZgrC1NTpImnVTYLf
dVI9EvHPiUqq/VDrDYaZzOBZylE0oLRc5/LcIFN2xvA65D2+CfI59O4nGIP5nzTb
wxuDu+yuRXryCsQGA8P/xV3jHapqYE7jE8ES4rrULZbzA5r1K/9hYjBW73Fy+TQq
1WgSQ6N7r7LlXU6eeyLchh+LO/Oy9c/H5hJZPAILFJJeEhMeVMwVGelQMY3kWobk
QrxfinOOguuyd1Zrms9Bftp0Df2eEy+mubx2K4zUMUmUBdN1Fm4TAzGc4bH2SXtL
bv0tHkXWiA1vMEEJ9TUxVkjpi0oXLLcNRq4xOF6lRPZrxbPa0kavOlVRmHguw9Dc
Ebmu2+ItEM0ArlUW/Oh+Bngw6lwO5dycWMGT7ykf4AVPKr4Wr2jnGl5RwSYGicw9
hXysE3NyO1aniMZX+nSluiGTttRD1BGyUHyRSzatMJ4S/8KA8X20ddw+sgTxAI+K
S6rCO7GcoF+97+Gu2DiHeeuLVlNQDfGN3B9STuuxyommc1/5RkDFVXQuSw1sldpl
ApqRrkKYgMJhda6oy6dKyemsVEi92abf9YCFkxo+NiYw263spfYg4xkH0huhgsjw
m0nsS34dPX+E9SpCdL8f8w/mizVTg5fxqWHFWa+ZX8bBPjixPCQqgIM4knriS3ut
cW4PANcLvYVXlnCBqXp6zKCy1h3BXQDn+NEAiBHenRAoT6NiKD1qBjJGXmxSPekb
yWH2rorKbmRko5g7KpFZjfbjfM6KZOPnvDk3R6b26Ugn3mKekxywbi6f2KF2kWfZ
P1R3SWg6afh3H0xsuocCBtLPgWxE7CllT7JELn8xVpTzTfdYaPJb6vFApkLMEaW3
ArOjg06P/Sbpirb9MJnYZLpgDib1GzqzKjDQzWpdIFCI9Ve8UbVEZ1rR4c7DQ+PQ
SRJfEwwRx8HmGAinbTEPmj3lce4wysoyrKW8MpVj+hhVdBb0rHViVb4J71uYsUpj
J7xrHHVb/UftaN1CB90lr1URqch+qctWL30tLWDqPj0IG60XB/xck8oBy0INfSgd
ZziDUjyXQjvMI3ejaoG8gsKDkNUhy++jMc1kUj6EJdcBoXIXe+bJx3Z+qamK9bgV
ScotHpUjdDGbQ4YS6OJQMjnr4qAdmc29er+OmhwzfouQAQ4v7vnT1Ipjbr14LYv2
xeLr8/iyrRqWgMxIa6XUkykFcEwpQ9KPHfW+tPIpKZx6uMmo2Tjp5zl4jeFQRvc4
OvV1sYXtFgCqlTfDoP5BDPtLsHFDf948MF/Hws0giY9UKyEnZPZjqtd/+8BX6Ga3
FPL2W1Qz7S1RAPvJUZYrhwUYh1fPePEC3Sfy4ooswkbNF5JQTlR4XeJfW+5Lqq0S
m8GubFmDpDnTdO97GTWsaJPmV+smqyJjM0ZK5AuHhPWFWryd+rN4IIjiskTJOmTr
mtkiEnYkwB0L8stGdReQTNMw/njHb2qdFx5KwPTgpzD1EAwXyJtq3H/Agd/FPO1J
B1xuV1Aq57/pBaw8qjbRvEHjVus913qV0mO99XHECMMj9B1BzePwkCWdkQDeadmj
OfXHZItLWLBh6fFErqOArE7httPVU+EpLm2a4R+QYd6K/jGjb8IHI8msWV4PIL4W
ODK3z+em1HNhPPkp/AIbs4JnvyUItDTo3x39s16+j718+UfDign2K7/IDDkmTZa0
1d1mfLTaDUsc7hfZY+EVx+Nll7WUNDKdaNnxWC0SY4Crwdz3HlZj1jfEB86KA3Zf
kJ1tgEHcdZeR7zApHP9zjkwCjOEBvf8DDS7wJRil4+K3x2zOBqjtVgcro3RxxEHe
4MkZhPPpJdjjQlVvTc6OGh9YBxf8HI43hUwcr9/PDLC/odAzu9QOlGc+acUQag+r
Il7bTxJP/tQEmsVaWDC69l8aeFc/AUYKfxq/c8scpaGn+L9qSk9+QNoq1LZRVpBd
KLI31K/axmf+yjeVs6tp2YQJ2NIRbAPmJvMGM/N5733NeiP9ZtApnnDydfPVnH5M
u4ZRUufk8/vgjlFZMGK3ZiYUKCdopx5RvFPYPivaznHLj6+GekA1mSPwpCzzCqij
3/6WeyPPlVoT7fQ5wCDK52ACPPQeBiDZDr278o8asv1IXtU/CzrRnFawx2xUUrC3
+W9mrdZZfwiO2lHjhRzfAUHL0oMtm7bi7zYQwdwe4iWMA0bioa3Y2/FW7DhL29Vb
9/IAOOziOzgEJnNIK5uto9neDrmfEfBsM+Xsh0idFw863q5ca+aIPfBuY/HAtBhF
luCuRh/u5l1hQMTzcq6FSQWLky8jB47YV0wNmfqoME/KFL/Apa9TGYZ/HSkYc5oe
HKXYKMVF31UTIPf5HB7+YcGNGOhMUT5Wu8BSL7NGj4Bc8qSB9htYMJiNEdiE1Hy1
YPBZBu7MiHlfHpvtJxwj5I8R/6QF5XK3FGzu+rfReo+0mgQugCfmwc4C8AVLipxs
WUX2zBQKhlMQ7JZ7CzXvkr7RaEJTTNSGEcbMT9KIcnO4dGUHNsnWyk0UCc0+bti1
quZJ+ifEfVOCluCbQrv/98NFQFFJLmJVZkMR4p+qgEWmb0zo7zj1763DEEV/aotx
e9Z5ENf5rQxqbNWjlLQErdMWlmI7UHgS6gAO31rbbJRlBAMhLLoAnBdBWFy4fmFW
cYvpBaUTFGm2vYQsa+LmZMzlrJCGk81Xbo9V7+TVPt4+v4pbfg40qTDSvFrpF7bp
vZXeYcoxknOT34OgQYLKZQoZf2GqeMyUUkc5FS3yF+hIasBL3Bmy9/Gd7P/Q68n/
e+Bz6+kl45VgP68/QW1Zdo0C/sMb8V29CZMGeT3MRYye0Ixf1GU0VoGnBukWT+Lz
qngW16Azx/tZN3ET+hDUkxoUTMJq6BqzoJ/+hMQERkmIWPh4kdOQHDsM5nkh9BIB
30N9y6idhPab/as0I94DGjYoJGi/zHbVWUB/Fx6+hYg8NnmxuhopjnMwi7mbNBe/
xmSjvCPARCiUW1P1teP8r8MnXq0EBAty5TzTZK7f5wzamkjWeZieb6spEGthrGR8
/JpfuSEyQP1/zgQi8tMHxWmGjojwlzsBgyaz5sapiS5SNLhNhvECemez1dVRLuq1
bOWQ7E3+5YnRKKTESB0B3cLdf+DN/l8ysXUvOy9jOddWHrA5Co2ArudXzPxLkGVK
JIhFNFk1d5qYKvD7EWe9To7x/CDceucUFM69XFOL0re/TcCbgZDOrZ7cqHesZHc3
Zk5RyjyJsm/TBk6Hu2VDDxznxoYU+h68jBX0MBo8a5nH1/6shzab5/RONuFExS+A
UK1nzSfCGtsdqsFL0OAZkyNqiuEB00ID+BdbPaf2eqXDBDxgn3Fsq1e/F3tqkZem
uR8ECWUMMXl/yB2Lo4ZznO5I0JL3v6+rc35KO9P4IiXIYqdQF4YllnoixGBuZTuc
bqoP1hRf/oTe+Qtuq+8m0obeC8w2SW5Oa4KxHlj1gSfjSsiNpXkHELgDV8CEWwyY
NV+9D0cITLtFPmV5mPovHBq7mHt6d61OfvSajcgdZymR10KtSKagtSDZ8ULYdUH3
+OXrk51YGtRO+dq7a86GxZIvWctPHYxvhO6EMxfuJJ4rRj68v2AY8+6sxp0SiUbZ
hx8NVXupZUXEIZ0Bgd7M94bT54Stslo5olBKfzaGkPpFTE4fz3Nhv7LGwRhfgJfV
3KGE3zLmrp4uB/KamyC97mkRUdPkCARCN2swcPGLvb0LxAKFWF79f8lzsK0+klSY
HWBnRgHP+B+T+kf0DJFVcqtuykEtFHI8lTCZ8F8glA7+4hSai+CgbiORNSOaZL1c
QqkpIThzYkWAWbVnKCLE6pQ2tttmS8ynw6QTNDx+cxzBOEUGCs0582UcvF1pkx99
rChOVXxr/xxhA0s/dhXjrT80WPc83xs+DlBO2jfyrY25Na3BOlkAHfTmXOe8wgf9
bhertGYfj5ow9UE3OuJEJB7nov8hJau0z+PM5MOAV0A3xCENKpVksgpwX7IRcWx+
S+pgKiVOL4Z7Vb0rhrTdgBjgEolyx++h/fXbc8aBEcICDdgD6cCca5Ng7OxbEjMM
sQZJAdmS6UML+9YkgVR3NaM7DyK4vDgUUG6aReLM8t2XWUEpNzm3+w471tZEl4pd
flEo+TuLSMLhiTa4+IMt3Uqp0hy6G+9qhDKiQgqzoUsHBukv9xKicfgG0FwLz6aJ
mSLhEMVTBXJMmOcz6FemLjAcWYPBQZhJD7R89NaL6ahdX+wALDZFxF2KU0+m+1dp
elprJQwN+94EtsOmfgwCvS9d6Cn8dr54M7yI3+yYBb7u1zyeIEp1Jc2FhuMfg8Ue
uGdQAaXPImIkaF6WBHSE+XrI2cufEmrz0Hg6hNXA0Ov7i/PV8Y7GjF7+nsdmaaKb
DB+mBuScjWEJYljmLXI12l7sFElMOJC123fHCpKK8HJDcD6hWsPNC9zLfn0uU1uA
hbUhUxCDxalZtidL7iuxabJDwAYyDl+qpc3IAnBsLjeepW+H0yvGKrhS5yYVUFe+
rb9ePJvy9BA/dh5pkDEgVy52PRJh/a01z9lJ2E1wZYRLiPZxRuygYfcO4VOs/oKE
84ozkEeaaWVmn1S4TtXSNOwDVVnDk1yaPg2XLcmTzgeNmJBykNrfnuoBtzL6lvjN
JW6twoWF9xnk8UGUgCE63LFfyWJCOkXcrCpPgtnP6d1CsOJ8fUTO2silq0Ivabpv
sEzyubibNCFha07cX1UfCtGo1TArglmFyUZMctRSQ3N1eZ5Oiz7Jh8c+XeUn+bes
SVPaA/jbiwvemlyOpnEDY/7kSdsb/47e8ciOz5pFMc3o34VEim+h1iHQjjl+BaMT
g0CaxgUm3Yv/09c81pTD/qOGuO9rcSckNHp4j3xuGuU94wY4d9bdYHNgPtMrrg5P
n4nkhU7FTGYwakhREHsXlKxc7SGpD+Uwd/+/ApxolOY9xaOWInUyg2XI/pl/Xa/p
9wgDxaai2vhBi7+z+YlBdSx/FX1tPwe/dSeJS88v5meR7pAzQXHLLxHH8mpXNP/9
A8iDjvR07+4qgtsWANfGLl87X7BXJJEL8lKHBcUW/h3TZswwwniM0EApZw80P0XM
5lMDYmd9pW9WbeQ+ClgmMiK6oVzUrVEnCgoCwUr0qTt/071W1+NJlTo0prRXNzJ4
X7aJgb12qJ3bE+sniFhZ+I/FielX7UqU11HVtYYf1dAm71q9g3XcMgJPsyOx8do9
GYV4wurWdO63Sl3Ji0GOPpUqyjCMOsA4jVq82faViO/tXoSrZUunORK6nzRhp9OM
JDiNJUx0K62ZHVPrQ+JJUZDNZykEBNsKLSf1yHNGi1K9bi/iL5mgASaH5XyQzstW
Cjtl9W+muwFEAqmqoM2aTOx+5qwFgeL2i/9n/0dEgjm9i40f0vzTXuStFtEGG9HH
LJboWe5ogyKzaTayJWi2//lbv+ykgwRD08QITbfPjSOXJp6x8mGIobl9X+djzwZT
+EMg2ar3/YzxefdMa6TfBfUVlKJqxUR60xUkREcvhpXqT3Eegd8uM6PLoOdMfSJR
3KGIB+oKI1RJxFPGPZttq1A6Xf3I4MLOgqw1KBJ7HNycOB1/x7gyn2DsPImmFPqj
u2YZeAwzcDoR3eNnAke6PXcf3sN5Xxkk44x0NxihWPsJLAbTgOuaKc467Wt5txxK
R2l/9oHhQNP3pEhFXxCYbPT2iX6ySp8CHUw9EA3ZRSObX88Kfs7n5OviNXE/M8T5
A9wIXyePdJTaggwA2U1pNIW6pDN+twlMnc8N+yPieHN7N3u3Ff3q6ETJHDr9wo5r
gOTbqrwJ1ZM+knNZryfThbHLiWqceNc72qPZd1tVhv2BITWEgsyY44HdtU6WMJP0
XWOtJtVk8od6ZgaqOi5MBufDuGLk2WwIWp1LfYiStEE0FDM7sUMHbkeozDhEh0j3
nmUQm2BoyMhDB0SdojahgeeOBhvXFdZwmEFMnILda1syeZe5yGg13gQrekv769Zg
7X9rLnbpjJ3t3JDeKv0ehAJeh2V7/IlIIMlja6SMTXyotPSe6w+mdby3og6xkFLo
ATksZ8T+WJ87oyy6kjo7pqPI2LnC5Nko2rYCwWysDkgf1Y+U8Baoi6T6Ryw3RxXc
CXAvQZOgpqjGSXW3FzVHpLfjHATiMUHA2m/L/14UXS1rPQQQT0FiIrChr5TSWY1J
NZ3uMfZtAt8NnqS7g4O8kOtIo2SNRvwae15GJAuPM2YPG/viM9+zMaZaFhn9wQos
ovqQqI6AIOzAJ6/Kk4FHpbHzAt/XTXb1bKeGNOV+RHDU46OSPMG72e88ACkzNFHv
+GFeqsVBxc6PkTAiLHfvZKaFjZLrjOKqjUrdRKGz0tqN06Lufo/W+HHdyxrd1Qgz
qEmwT3NqjKGSpDQ8hQrClKwSIumHhxg3dU3PLlvyIixfY893gqAYTs6fDWQPkkdm
piG2lMOR1IQKcAMVjZJ7wBjXOmbgvd6HPYT8MduC42oKY1i4Yq2i4sCIUa7ZbDgd
Qws5VyiweyAVnS28kxm1dc4R6SbojRe8EkCSoqefcjMLGhVWUvpcRI0Qc6UjJ3DP
5eZW4iBVAvhZh7gUqomxApuLawQKdKiYImxGrqk3bbWxfYXi06ZItGb3blIrkvev
nWbv19OK5wGmp/GyHREVK9Bq4reyXEXKVXDaJQDSdCt7dW526XyX5/y/nFT0dJNc
1xDLNzObBTcCyyCbTSlvgSpDD3JtaQaajsBF2+bl6jNF4hkZVIbYPdRARgY+nQ8X
aWYMO2b6W344c3HjseWseKfqjTv7YXzQKRSh2OjWbiSO9xUa+xdkL0wLYg7N1GNn
FJ2USjb+AdjXa+dTfO3lIClKNP+YvIkobVksQKHlt2Ri16WSOXZFh2RQ0lr2Ov7H
OAWvPcfhmoEj3NA2oFeektjQy4xvW9ZBOfMsZh+2fasKi9ap3AGSImV5KtyNGhvn
UDHoXv20gUT+vti2hDDe4qUwxmQmh/19sGeLZnzQuPoyFiffug9mEHKIL9OOZPNW
R2lFhgPZHpIiGy5p2dO9+88WOxJV2vn3WClhoQopAofyTHd2dFE6bor+3mKVmx84
/Bl+k4GatW2U6vPskxl0Y9i0Q+vkoAMvbgfbEIMUOi5CoIgUwNNnJQGEC5uxnER9
d4QpC5H9GPg+zzQxVVx9GQ9GjzknhhFkje5qMco++v1aW1ySCie7ot/H8U+CHSc3
tpVXBtf4tO+Gaalf4N3LM+JKq/APgwNrFSFTioFjAgVLziZBTABVW9OcNiPMONfJ
Aokg6rNp3kHYcxAMRGvIrfcRwr75JZBDOUiugMWmu4ub9UUGlWZwBGxVB+eG5MRx
5vDfLPNC8EjX9NHO4R6pzjmC1WHS9VV0eaitqLc8Rz7K3mVYQ2v9ZSkYMrZTAHrY
n0R4/ObDwjWM2KxBXsbC9xUmyjCOrhQiIc9duU6xSlk+iPQ7vm0W6oVOvTj60f27
FdVVfN6JzJMR1eaqLfXeSub0ynIKOlVal50ojyZt5+4qBNyM68sZH5mId60FfTfh
48V6yuMRTEO9gpFiZTsbWIYCv1neqxtEAXAfAazKJWnSZH6YlEliFDXKmMocGRFx
kFFdm//tAOA8AzAh01VSSVCuupaBI5E5iPDv5eX6kvB9PCI5pc8SPnsQJQ5644SZ
HuEUUiGuEa534h+NLEGwuJvlhjmnS5IHCFV1XrNmTFrKG7lmgmUYGBieAFz4EBRg
fAHmd1cG8cVxJfi8z47HKhmsSIirMVffiQZ77PYmXXmrNSFQsaUwLVI9GVCUucni
7NLe56/8Vh6Rm1TgsJ+a5+pXESu9tDkgQ9YEHFKiTz9AwOTgG9PjwmdPvJgnM9qz
hkFI7UiVOCVBE8LRjhrQfWd1qSXjTh2AAUPFfoLGPfwxTKNJ+7/ONqwIPXAzt1N2
qNLPA71KJuSFxIqDw7tgMGCG9rH+YbDeHabc95ZiugMuiDLUmKa0iNwhrxGmZvTE
uiVnZA3/DyZzOW+sidPnwXksk7HJmiLfCPrLJnJ3j3HhQh91MI2j4HI0/fFEWULo
u87uQuRFHkYGvX0wYeVdYzAe76m++5cN2i7w3TK4iYSlnOfOfxJSiNAwdFoNvs2F
3iQIqo2Mw7FSMk0MyqRqiNLsyssLXQR6DhTo89kGMhJAgRrLOY5uBj8ZtpT/wu+L
H6TBiUOZV9oytTKYc/NelvrHDw6iOjfiT5BkT4rsnw6WpC0GJ0v3p4k8oYf2ostE
QBp6uV3+d6UbLfuo0PX9G6LTtNo7IyDgFdM1sLtl/5x+YARjZP20C6CM+5X2IziJ
tCTSQ9vjDNSoTZkIAtqXsgGwIlvPSvFfz7VW0nrhuMi49nISLL6cO34rbs5+wu37
dDmhG32cgSqCpjKOzYQKSLqP4ZD184xGXN0y42dmu7N+awu/ZkK8W9cL54fb9acZ
b87IiIsj39DGi661yzJbjP+Lr8nFOwbCXDD0ZrSgHGKHklsv5K91JbELZJ9PwT22
ABAOSZPCeD+ivoDjpvrS9mNTvsFr8VrY1qAzEnjWBt1IaVkIF6HQsUfevEV+WRVJ
oZfio5TTVGdrb7qp4Rwje9FHOX2irheKZ72x2mAvfpyWxVkVYIJeW8Wz80JumWUE
vaLqW/emnt8KBfB3u5xU4FKU2Ak9l7gauXS/bRwA+NlVn++PoXEHUZB67KtzKsLW
q26PP7Y6jXzLHl83r3Q7EwWLgLPrM9Cy8I9BsWMMgbcOwUU5Ov+dw/GUT29oAumZ
hfG/I8/zGITJoBGRkbytNX8ulm47WxRBk3MGN0oeM+kSMvR5K4okNZpDzYTOGW2x
n4b1FmAQS4+SFdPZO7SzV2sYq9M1ZClw4ieBqYhmk9EJ8YKG9s/IfO14b3Mjm+2H
KZb02ikB9BaK0CLajC9b1Yj7Lobe3PG+R74FzpwFtF0qqwvJ+aVQLqKD948gbeZ4
6+zjS0vKBJ8EmfanFFl8C9usl7A11kfT5sfNBmlqkmTM6xV/jb8NfSy4sGx9OVfE
MnmsGjemM1cwwPkjE2scndJx6nmaT+2F3V+ik33iZ3MQboqsH5dFWFw2UzINx6tL
EWlm84+oYZDRnFRxeMVWApL49qhLIgc0piPwtRBK/agqRccc1lzwUBYoJbrLndua
0Tw+hBDQXSP0baiC539dS6gCwRcPz/t6AdzIORdfau/6v51jGQzSFJCHpzD2pIqH
2KSKPYFs0Yh9zeWFgWhKy32XDCjN6GK6DcQMFWMk6Wl7DQf5r8a0wdCcTx1aVdyh
0qjPWIFmn12FAzcTYplZ2tp3CEPdypu1ve5RNo5GPZ3zMrX2QiaahzhGVjEKnWD1
LYeRYSp/n6wJdW3D78Fx3L5m5oYwcr8Db4Dvg2B/sVVOlJnC7hC70/8mcxqDqUjS
TdICpdBocnTYIV1r7nPdIulkE14LVKNWb8+IXU4tB7HDCWz682FmKHwmwbGsnoy3
df6B6lLhD9s0pSa6IOxk+V2xKqN9UA0X63on1+qZhpmyfJ5gvjbW/yf/K6nguoug
n7AUgs2QKfVkmuXyNAg23DxudqXKEjyYzQw2zyV7A3++4w4KiToEXHXQOG9SsiX1
uqlbh/HuelACldZm3ziZDHF1g/L/52lF9DWXWHUzJraZadq8A2aGqlOeVnvY6wt8
Vwhjz8/yldl2vficODGVFajUuXOKKWNnLwzcOqkfkwccRB5ftjUlGwFBEMqDIbVM
I1r1WOF6Mi4RnQ0iYZ9PJPwNv5/PWYTOD19NImAQS9BybXBrcS6BrBwABKs2WfDZ
aXVh8R2FmlWN5ligu+v6vOjuLe1ZhFZ5f+fXCZSuNo6pPEqa+bY9kSHtTQVD0DCS
qrhilavPfIVnvJVkIigj2L8+E6FapwU42HP98gxq491kECNJmj7i8O1dSxuOKYfS
3LuAZ0tRdfRWkw+BGDlCng3PZmBr3RltQw2I/UVsBA0ncgg0PBcVan/QUjt+7H4T
2IFPkZibTyfWLyvUriVO/T30MRkPS05Cl+lFF4zw3R0BM40hUbPQxUwS23D+tqNh
QzqcZgp2DudibdAjQdMZtIopbyElDOrhOQceNHYMG2yR1SeUB9oR7EmxirHm50ow
dL6XiXo6rYoMUdQC6u8diNjJxCXOZI6/aZUNWDz8YU152XsXzG02jNAMCuRuNIyF
p7CQi7Q7NUWYxIYrAtiSDQuJYpLJ26m2uzR4vhUm94tLoLOrq9VnDUtun1XZ+Q3b
W7Oph6RWG8IyDrRS7aoXPDJ29y+38DXjDZTIbBBdu0WHW9Xl/cUZ6wDWVrJxlHUf
KisHWx6URTg4JRQPmUstnoxMHjfv9V6rPz2Y1JEhSu3deVwv9TTTFRxDzbRSjE6O
OehtpcRBzdpsBBWV2JEE2staLhUSbLRhe5f0Yl06VK0nEuAly9WB7km2E54yQ46e
fz4MOAGV9Wbw2pE+2S2htXy7Mb7Erp617m8m8lHMitQz4DTqDdz6gI7dYiBTH7Hb
HB6I8Rs/9ffr6Ud8NOxiQLF5+gQm5Dsze3hTob9Q/piROU6YTCVjBObA0s70Lfxx
x5w6/vvHn55EoQosk9lD2uZ7gwm7BLmakdqDCKUcLATgx7q0hyD6F1AASG3mx95Q
09fg6WNxC1Jhwah8JEAbmnuY5pYwC6Jl6rrEvTQu3AqVejJua6ntBO4wg5jFlW84
9u6IM5VevFtUzFy8Q2xJzmKiArBXT6Z1xkGdc5ZETBrfZyEEma5WwbP0MRoTw85X
p1VzHqZ9ZkTYmsvIOGBAiHbmXnUtpsPVXZKwnRzzvYMx/XnCkr0pLCqDeu3bvAPj
DoY554T01r1hprUOcZnuL+KTFt17K+PQtzp6vV/9L8VgZtcgEzw7p7mwSn0k6ShE
31ICAvfz06gnP7kHfPVpKgbVHrpIqzZAiSCGS9NJXtptMMax7M+38+Lc4PHkvFiy
yjiFvHLpIld+RQuOpOw0CYGQkwYHYvAUFlnqeGPWLYynBRNl/NmC1/sXSR40pwaJ
q6yZITnFLcLcGI45+PLwqOlrzwcOiZeurbCRteGpf2IGfLcje60YoGfTBI7fYSwr
HhQ799loYTxVhzAS0wt8b2yb6JIiZcnlBMb2NojQpBHPXuDM1teAL3KQhFSzbYtE
YALS9zeLBAGl3vy3O2T95E7LRW+qSeWGghTSRpG6k0BkpnpLPZm+z2lcg6s6pEnm
EVhG8meIZboeBnJP3uJSmKXyKQqTLxD2IBSUntjVkMAMJxuUJcb5KwhxpGneajf6
sVHRUST+6fu0WbJ2sowZr0oHCeHtiOTqShA/zB7J45VRMeULkHlNJuN2CVG2J0Xj
t9/hV1pJO6v9L1U+2X39m8qQBw9s1z8Kjs3v4E3t8b96qTg7Qs0kdYLpcWqThZAe
OqH6LlYtv454B8vpSK4YZSoO7fqflRq3EIJsOnST4Rz7w5XR0Y9SO6dgFRdTzLKe
hQq+CEYlPb8AI88HIJxIdGMDTBhMYk14GXs+BkY4yY/q735cSzq7EDvxwk88n4cJ
bGBwXhBt1xeGyTKRsEF4Bp7iPPqCRm+WiYMEswwAigfiqxvQHXW1bqNyafpo25Wx
S9NervsmY+hU5FgpOiW8EkbBgcEvPE73oUpgCIqo/NfakY3NN9kmWQsQl5GYA+rd
YS3SQIahiXyn2pYFub+E2tzKEoWCjtRkN6Od46/HguZcNmR752ht2ETf9y6jJI4f
Mz8O5GdUD8+wnaGF+VAyLw9R9E+wXoipFS1PMNeedPFxOVOnX5SCAOb0LH+u2uyI
fKqjNAwNST9FcPXMDVrIn+WktJVsKqriAyjsO3csQ3/IoDp3FXZeax5M7+tY92c0
QF15WYGdoZtRad1H6d43FE2z+n93kYoqtlpwnAxqR/l563ASpJVYFLtFOBNJM5x9
LKLesbv/4pOJ5LIG7IoSIR4VtPflnrgxBnCj1gk/y3OI9DarcKGSuTp+j0DHagVA
dOjmo45hk1cpczAwmLgJM/m+o8NiZKPefPf3VyMiPxhUljXBWNlASunLDRO+cqfC
dZYQ+em2ZrbMb1I27uqbai4sw9zLUIFCMmEXEe3dAzoxKpCa6JSU9qVth3cKsQi7
+qCzFTb6xrweBgs6Ksm8G5eYPGo65eWuVGW/rqC27TREcXjKfIG/x/+Ed3JmHg8K
tEcP4pxLHIvWXg4bb7BtkOq6I2tTzEvI7JGLjtHAZHn5sIcfhovjohXyjGUSLURv
VO66yRfTMLZvC3O7h4O1AHOlp8NpukQQJMaH0/mQm8sXUaZWZujVYKCzZLJN9HTC
8rmTUiTHysUY+ca8Q89jdPKZqj4IxPWGqsvikb0qvnGkORPDAPX4HeIVnL2/xkqN
uXoNc6i6Qp2Thtx6a0BbfWMOXbegS3QmvmdPoxP73DUjp0Dsh0IxNhZT0ot5inVq
lZlQU52mTf27WJNxEuzT4ph3Y1oCPOhiLYgHTKj1etS6DNk/yCebOZ8Dcld5VMTX
A7JoTyJcfF99C07V1gZSD1o2071ItoAofFI1MUwAnlWhsor7Ojt5INhEtGECxTzg
TVw+7Kao3bHzGU0s+K5jlG/8hghZG49XaQdiQI+rgRAibcN0nT+jUNhJUJZQyKSN
JMXK14O7chWvXdN6REmZ26w6M/lrOvfDY0dFAYC7MDpm5zBxnwkrFKjfZRZh0+yY
VY2pX3x94FTPwDHbLar3KBd8k4f5+Mun+VNmARYNxPLtfmuxnlh4s+UQQOe/619b
J4aLgo91u0s/X/+OjfhxVK6okBWu8v4yGH9uKyGU4mtEaz/E+mvhGK/U6B39YUdJ
DkBwY4Ow3i6oWIVxqNcS6TU51CEiV9JnMXetYLhd1uLBfPuFaSpQl93djEyVMKxm
lKbZbtHYayU3ERXwkFwY0RyfhKn2ekYwsSheEHrb5IbP7MSylj3WVfkAobPZF7+b
tYFFop3ui+y2sxNQAb9zCogynFwlpE1XULcRM/rnHvwCtjAUSdXHRYdumUjYPFPA
ooDsR6neB9pSw/GYNMj/krAmpJE9NM96rl6tQQfavD+Y231azStktVq7niYRz1Q0
cFKtk86YiZ6KVlKX5cb5o554FivNcRJy//S9XBZMydRPkdGOXDWwDFV0GKONFrq4
BuI4lK7fABncfxtuDwIzebsjZ4MuJSMndymnPLoqo6nZsyo2S4Eek7vXgWd57Koj
yngmL4RMliRQ0FmfeHZsznPI5v3tIyLfuenNTrOPojXOwwX/Pw64MeCGPh2L1XEZ
DWPX2y9pEWFDyaSEGzBFFdo5fwy68P07ZnG3RibbTcawDJbQACVIznn7cGfj0Bcq
tGT+TuV43vtcWX7oyn/GQvoXJdAAk+VW1xD5YiUWmv0bRiUXUHGz3A5QP4Xbe0oF
gXGEazor14RqQliAmiGxFAu+dbECjzOmcKl9AuKSUqVYcJV2/ZPtXVz3ERdkpEOV
PtKgi7z8ZwFlfs1yvNZjqiqSdl6i/NQC1B5EsIY3lmEUyba70MpecxY73c/rLds2
Q+L36iN/hvgTG/1FGC7nkXx56WjWDXgLw8UPf3DGpx51+Pu4uwnravss2VPgL7B9
L/m5ygTeivpT2BWE+dw/GojwFztPJrQulEwmPJaoECKcEnPcLIJ8+aZ3yMXH9toy
MwTMjFNO67mvLcECLLpI8cWAGGwtARHGt5n7iAK8r8EH8pa20HX2qljNHgNIZ1UL
7NAbYB6hQ5zCbELjQKHoZS1hMiPL+8+Fe5HYQfou2O9ckk9VqqNxOWICmqH08wfR
5YzdrJb38pqZyqErM9uDxFeWdp3TlMf3G9xgOoRJThfWCYK4vvjvPxi0ztC/4sXh
Xrg0+mkfv886knEoeqD0K7IyvVcFFurd6kLGZX0kj03ERN/QYtV9ph9HTRTO9FMD
Ef3PuYX4HZHhVvCV0Z7PBLi97GWsZ/vkneN3zIXrBap48UZ3lucXgO2Sb7wviisH
wWR9ztYzIdxikVggs3tgARLRUndpS/xVeKV5mXfMECru+jG2pvguf+oDgBlbYGBo
szZXBYTZiazC9Dk8bKJPoCW30nvwLOo9mM4aFD9SJiOW0SoQiPswYyYNnuX8KZmp
sCAq/Hpt7VUeJM1OZrW1LYPTY/sS9nkxUujQVkWWnCavMHkUEMkuCezAJ7r8gKtE
e4eWzXm6d0H/NpIXugp+BgqT/z/Xdk2w8jNLlIVghaIFWjuSnom9OHyX4g/EP/cQ
pV4zPV7SmlJV8vsKe7571x5PVF7uWHt2Pjd4cxDc0pgBRhBXYzbJ4QRMumjHRqbA
wy8Dnl5ojIdJBMHaVkTri0jthBO1Q3ei+UF8gtnM4EHt0SiEmkgLdqiCmTncEqOM
f/SBjOiu914+xmCyyq/PteZiBv8k/Uq0hAPT92y7fJoRs2F9uGwW3iFE2U2mlrxS
MwPOmz+ME2aQEGGCA26UtEDgRZie21vULfOE9yY9wQYweCfd5pxsmXHEyArycFDb
YnM3zNLglCHPpteV0EYyHNcbhUwSyqYN+XJYFIFJ4q1Nv9+jj4GgdgtD3IfVfV1X
Gi6hlKR9m8H2f2y6XrHTZZEq079Uv3MPVUzXyRDmQ8yGVvTtCQmmZmPgF0IS2gD/
DRJAFuo0VOXDfQHf/8ls2fF8HI/ptywChJn3IsBqPEBJrbxE96WEi6/yZOxqwziB
j3uNiS07YFci0mtMmBh3xQbZK6EUDryq33RNRZ1nSNzVGrmlhiANyVtXHuvK7nEy
7yVtxM7h17Wv/e2xKg26ZlJP/DP0GOrsWIf6BVS1hKRreoUfyHz2rzTqfr6128T4
PKhuJCzC0xnJZVoCDWDgHvvgQv1+60/jvwBgwiF4ZFfrSRnUWjbkocC9jkS7btKz
SJuVNQhcrB/IQXd6QDw/q9WgMwZsVGomfpDekM1ysgmGKPkVF97RqxkCaJTgxxti
/GaMxZ0GPSON2sn85ryoWYrraPiWFvgRg5ttrTa2C7KhTUEaYtDIATq8aBRTv5MN
gllwAStENw1mUmN6fz8L1MuQB96F6m5mv6F5VNN7nD88PgWzfGnX0dlOvYdIub12
LQ0YXX5faW3MFHRE8JpVv2Yx0lj6AgVbElwXCBGMNJDFGXawyf52DrGkGEULUdFC
xQN1CjLFq69JUoHQZvxpRvsL8q2eGQZbLZU79uIhlCdVfs9w1dGaDqRwK0uwnt3t
PV2UgkbcogCVmQqilsis40zHr7407E/WeloXdRgo/Eb954pM37xcOL/skVHKkdog
03w/ZLcRW0tAxjNxVZuGoX+nBf3yTSRf1kp9G60I3Ge5nT+qg33tDX5bBh85+6p1
QERW728uTQhSr161DckXhKD1dqV3hL+ZUrgnPDhjfhjNfPOuwOWy4QwQF2LUtB+m
ApDlIx3qY0fDlREkXgXhtRtJGM402mX6gPuu5Xm3o1Uqu7OiHAgjFaTdY9t5A6Ma
JXrsinVuGHaFmMwsXp9N9DDMyY+HBovX4PsV6byoYoSxBT5/pDYXEQy/50JePKUt
ZXl2mrSQRVBZ0DxW3OWbjAF3EE8RAfIMq56ffwZGZgyacBB/uDOrk7UWvv4q8Cvj
pjWQb5Jwu8jGMc0DsQ8wUrtefz2MlqOBrY1aWcmR0+UNGRR+YqSe3Gq6w4HJNNQ+
2fW+S8zB27PAFD0cXr6OI/zTlnWaUg7Dj82Vod9+KtGkfCGWmx8k5297E6rGuufj
C6Db7zu5FBHO08pXe4s++V9pMChn6huEWXeUjy/oJj4P+XkGqZ92IjHfK79hPzq/
wYsNgR/eeQs+7ZpdCK/wbI8bWWf0kJ5mmo7oQO+OvMqHWbhSf8sNPpMGOTT2pe83
m06ChVYqgaMTlnPI4sdvxbobOQDWF0p6t7Ao5MwJqZq5ine6YLKeBJyg9Yn9NrD5
7uSpWkoe82bQhF1fuwCfYBr3qW8lZaeB/vqILIWArpZxoUkOyO7ucwJY29DhFuxj
1Bbgy9iupffaURdiPmW1fF8lXCMT8NoFOe090u0Kf/0F6LNtlYhDDGjQ4qxAOhqU
G7al7/FfqHKLGdiwCxpLeSo1mr2QH8nvNd+8gYEDkqtMCAhX9pJjlAzdvbvZMsg5
tU+JLNmK7LQRQMK5SdCuIat31zctWLFpC2utDGSLRiwgA7BHtQlQWwVwI9mlK0rA
1ld9XqSFI5gMIcI0xbs9UkeoIER6gSVnHzk21nJm0F2fTBb2gcTFEndveyBiAs3D
nETsTdkOFAcxDcZLLu89wq6pOM8M3BIoqaHF1RMA/IZNdxWvL6rJyv3zPi+ZdyvQ
gTzWqrlFMtxncHkjDWdHeO9A50uher3+XPpLwyMuJ4QhSQwUfkbWiqfS6Hxc0gmR
0/+LN2x+20yMQA8iGlLPBGctBwtSeed6vouuwbK+FVamEDe5hqE1tICQnEvTmCEw
PXp8/Nrm5lOpw+wXCRuQRxwdQL40auoZN0WO21h5fN2We6iPG5DsotfvA2dNn63n
8PY+RgQDCXokRcd5+yfVcYObYEw2P303sg4yRPs4+Mjzq+E3Q/ncmzekiF+kz70J
MAwT6vBJ0lnFuolh4pRiIYAxpNvWLzjgvZgYSL5dvP0BztXQswbquvtvAqwDQ411
UdVyBDrkeygsPjTSqgUAOEhvrNB4xo6+x9yUEoDjVpRlMCygNi65ZPwwujLHQHa5
d7hsQGz2DduowZrF921+LCbJeRXPsrJpTYnUwqtT4J4+xwbKN+fZXtKFGAvilXQt
uCtpqtUwexzmzLVr/2NDNiyojc9myiTWjEDdQ07pUbwyTonmasxghCMJLvWAig+d
rxQj2KsQ4DUewoJynPZsiQqwDj+ppHi760WcNxGy/Q5UBJ/Cn6NZvF02YkUwxIa6
fzIw1sYJePK+mwgKcs4+PQaWY0nQ/sKJY5w0AE+BSHjJ1sgTQY01HpudE6gFBCvB
n/JarDTnEF4d7vg0MSi5k5lxY7Wq5MzN3LrhFNR2th8KAAM+xkW0NzmS1AKLjvhd
FXZgxH/74CWrVadYDWTbn6YY8y/t8LxoU9Dnz8PDGAzYwNEt0b83Vb/onh2Z/Ksc
uH+7n2sZk9GCeNzmiKh5ODFzAsLrEe8zt51sJI34ita95q98PWkUsQp4Lpddk815
HjiXG2AVvTsloxWDFh0niOjiyGIAN7sUd13vALuRydWizF0lvpIlusCD8S/9UxzN
/A/FLXPNmlbUJdDl7uNWTRl+uhPGIMBjb7/mHxkyOPZ4NHEWpd5KnKrLzNmr8+t7
D4d/bIyN5a85eaz0VUWWCYjTjNoWSCOiwc/iZ+X/MJzllqCSROGbmbVdYfEx4VLl
1mm9r1/TLR7M34Ven6nUpZFi8deBOe/juVgHtTwTz6qIZ5EjOZ0/jREu77SOCQyC
vo66yO3mYkeuNQkUypgr9BdQKrf9EVOZIsjL8nBPg3CurIALJ/bjnNAXMcdq90oG
giVkd06y8syjIRXH8pd4YEbelC12vSVXF9SJhuFCfx1GcKFSjfFCTLd4IzEns2KL
akev7fTKgTGncTGPcW1cqsyN/z3zhT0ryYCaTK2/vPgo4RGqBkHzxGs1oAJRT9kR
bcIlzZWrsU3EhRigawKimWvT83Q6fcOYztVZjvcJrJnXE8i5QXuMXigbRtBGisIy
HiNwpr7iZOBToMfV5IvKl64EI1eAmHMsW5ZjJaHtS0/wBe3Qsr2YGPgTtCybsN5R
5OI6Au423cNpSKsk6uLrXqDGqVIocm312PTT91Akg+ymhlGfd/7pUidVknXihCUq
kM1YlmwrWG/CW9vAY86PaAfcGPuUHVhsmtMfGeH1305HCauNMuW/BX/xxpte/ghR
EVE3xnJ+urdQ2YXpcsI8AjwIVHNn+owdVRq2UNfIeq2Q5BBju8UuN8DtyvhT0Suw
w8CKd2t4XZdaSEklDnMmvvafu5GUvbb7nx1DvL6kRl13zU7AuG8koxwxCNRELshz
R0OoWtGmUyWXFkS+6vfsPLUx5fz4174ADoTf5aLHuYUNznPksbySCv3ToDHfmPQ+
EL5H+MX7o6SBqzrO7UIjypBk3mMSn76c260cpUbCCWSsa8QOHEgEJ/gV67p/6iDk
rTRQcEO53zqWUiOElpwA87EMw2J/p9A1QnNLA97hR8yBe3MLrTs+M21d784ZvjsP
1FLg7J6172/xsSpzw2emO3CH9tzQSS2JSEp/FcEgt3b2DbyKsuJknyW5oFu8VyzJ
+G9ryuC6WdZRO4nfxvfnlCPBvYC3vfA4T96QetDnzz9RFhX5ytSXUGS9Z2P6krlL
hsSrVKIvFU2q7/1YBa0YtHtadoWmIm0J6PDOHqy8BfvyEOKCMq4bCvwXDpGoC3W6
2Sl9B6Jvf7ICJwflVOIB1GlThdzYFnK+kFQUVfszlI+kkA8S5gDU3YLBAz4VJwuR
EOwKIpB2GEwHEGJSZDtQgxlr/gYqiVXQbLWrT+9+ibJeAjE+lTXTcbEMom4CoKsO
+dwl3N7s2s1sLxfuCv0nMlgoWHTIeX7qrXWkBGZY/30FDkjDHqroRninPcUKAH30
JvfwoMmnwRKL54PyFLAmRZUubWQ3edJuUFGkC4onPzaKTBVhFSai57WcKXbs/+PP
BfIY5t2/01LG04dN65G/Ds8TUa4i1kpZUXilxdopIXTQ9n3jzj86mVi/Zsyr0sbX
J3dNEJ/qw1GOc3nBsWXrraPPzZQIDbb4x7g/Xs28et0xqtGASr48WM0zu2nd5M66
3bgmrHyOcerSr7Nd+WdiXS7BX7q2OqVfWKNpf8Tpnw5zOW9x76117U16kHD20/wr
kPgJZDz7PRMa5VdrqNL7qQgFvlaDVA+VtzUX2Gg6uHwd9j+o0dJoDtYcNtKeRhgg
UI5prVj10wS7zdFZ7hP/xVP9YpLO7bIY4475t4vl8LMaLjQ3MUKb7CuVBoQJAHZj
l8OtGuPPtntjKTCEuwN0ZcTIgYB79W9I38eXf+OYyOU2JlTpolKfEB3ujSp+T2TY
ee1Fq0dVTCGyE4a/9XcgRtNN2TmeqdYzCDsivm0Oxp7QglUb+oAWQr7S1DPGJVTd
ZLij5tJdAIjPkJEDJ8p/dPAl/JHOTjEcYxRNg/g8BTZGuxSo+o2R2yYXp4U6h5q8
Iawf1+oqdGqc1Y0c5ViFpRMkGqSzVEgjzUgVMR/+S0/Gsxp8Tgv0vhrFAERPgPCJ
U9pTM1zWlvBX0JfqcNqXCyAhBItt9XfkCaf+xBbg80wAYLKP+uxTE+xAC+yH/qik
0OgcOCgxl/aa8pMv6ZumlYO3/6ETuBT4CdKKs9MxIr8R1R5TGvgfF1CKYwVc6tlW
cjIemOMNc/cAr/Ad5WeBbgtQ+JsncswPG4EA2sOyzmBu/M8BkoZif8Dn39YUS9Qp
FYBUhb7JoUAcghwpJzVB3vFQx7l1rdExfiRk9q+wzzzFW2LsxM68bEo6D9B7lmSB
C5HcgwKHdvZqwS8LY1uIR0+Xnq8X9KyBJNxFevPpER+cqHvwJCoEag4vJ3Pohipz
rFxR+nzZkzXMkwJQtGjy0UGt9e5ZZYLad2VjW6BAzLyHVS44np6HLvQokDAjYZX8
9GcPz2+otk+nlD6pQX9t/PxBiBEftCce7C6yRlpljTstX9jdAX1/Ej6VtQnsHJjw
rsICApH9QDaT5MNRvqmCD7+ek3iNW+CsEhLQbsfWskeg/MFvF00HfuVTqZ3gZCoB
MGv9Wzf37vLYMO3eh9NMprOvEV90br/pyEpGaUMA8xdXZQyWKiCl7u4bGulTqAkn
WzWiQpFkky13eT/wIv8zSxzWQgcdDybj0QnVOyHlVlLtquQrrOOZKiD5l8sWA02A
rtT2Mr7DjN8lf5rfpmW3W/pBIXYNy+lvnrUR4ULpXTwm4XbviegUJdqfJl67xuqa
yyhzJUqPe5P8tZZuICRZJorLGEaYqv1mWj7oaFUFIUALX7erCFSf6s8S1oYkyJMk
V+XO50onnRHxIgE/3PoFtjJSpNi5JRR00/sq9XbdYYNov7ai24XS5JEt2Y7XCBEf
xHInJYIEdgTGaIIivEe/kfmuGCC8Q9Rqe2oBntL3/GWozzScP51c69I5eno5TsU6
MIdMuYpNe3XtYT1J0YbrW9Gw+kwE7BExOGL6SMglo8ZRvyvibcpd7u2ngb7nI7bK
9VMK4eD7aFlT9w3nDNsYlIlqvf6w9y7D3aT7vyiAJnVYnEFihnZbgtbksyn7igSr
83XoXuoerVn7AycJ4uLnjf+CMWbl40z/Owipf/f4qmO0ma/Ucxx6XxVpA9NivARU
GAgZwQufxdhFOjnHRZa2kE0mCGuLGoquaLM5CMLRdFfQfxLGmhpeIOoNgFcsAJhz
tlCOXi17iLSRnii99kklOuG0TZ62QRFcQxAHGy/UtMY5UAC4HakcI8tTWRrfGFiY
552lXPI/DZQwe08yCCLd2T3oIvXadpi+iK85mX9lvNzU0q7SoW+Q/tjC0W4n9NtS
s5fDlBFkJ7l+7LcgcnFSfilJJm/sYSo4zer60PEHMYDkRsab9dV6rLqxYEDEzrEh
RZblNqNLN2FUbYrSfNkRDt+oWmlSV6tcqjjVSyXkL9mbPQ6hcfEpcNixZ4dXrdv+
zIQ/HwlrTFqL8lRsZeD5bvkvxiWsq41Gosda8dyZdVqVW1hyUTLtOW4FBRuOhFMP
RIfyIEwATZMNNB5IqbA/UIDnszaeaZyBEWENTs2iWeLSCEYoOmfDg1vujLanWguM
V+qKfVBm5NQE1w84FrlDFuaf+27bUZP2TdQCXcyAigRgXdjB482sU++Dgbu4MEts
FGarKhdUSfqu1UPGT1sCzhpQDGTwFeg0WdRtyQ38UBYwWYrFgzzApNetQs99pLS/
JLEumhyg8QVK8JCP79hubED4+4O4CsM3qg3C09IVrgY6LNn5sfKeeKQIlbGfXnZF
Td97vwqKCCOAO7YkEAdRQoaCL3XKNCAKyVGHP2l5UawqmQI0+LmD+LHvo2Cwy1To
hdunK+Y+5k5Cbu0+ZlgPnssuknAhKzrnlLJMtMvoGxU/CXS9sdB8ssexndZKp3zB
C8b9yAmAnxHtOXo8p+ZOc8X28F5wWCzU0CuSAHPY/utJwGdfASSxG2r75Mw9qcn3
LGX0m9HGhRnhG6pq5eNeR2g87H0Wx2T/ai1H9E4qoZ/+CS9ezb2jC7AGPTNlIyPO
0HCqP5dhO5aedjCVIo0yKWe5oNpGf/ckHKCQbalcvFmXNAxGJvRr5Zrto7lWliTw
TxYEk1hGtt1QrcH5YLcdWUWbnSyROKnIjhsJoDJA3FhgGKoPVPbld+RKxrbxb6qJ
gh2EKBc0Rx0+7cg3nc/vxXQI3JhFTP5JsLudRHN5Wc4/0Ez4cmgIT+aqjXiSnZCL
dD9rb4ZT6/Yo/wCpru3/AC1HTK3OsMMvZgGCNYDRQihhGBxNRYvwk7PE8XkQf/iq
NDLIFYBEavGqEnXbWVpYki12sfkQ02pzXKsv+qJI5C+Fba9DR/IXEOOW4aJ3+SW8
qKr8vRKWVmDjIiKRobnRGw8/oFy0sg+yKooDXsHtSsyEcQkLFr4lfPYzMNF/oEdg
XJ5GG2g+IccucrdecOTM6Ggz0Aoycb7ssbJulynLbQGefWC6Z0pcQ2ewKWHGKeMG
QxIP2VixXe738STzzy2Hiy3cOFWHDyZlqnrg3n/5+qsllMFxM9LOPRpIyyMZlGTP
cozjAMz0K9SK4gjRxYCRA8x46xRObtGHdQUB/QqqthVXSs7Cqr5B7NnQclAo1STA
GXMwiveieBQwevH3A65MX8MOyKNX6NIOOuZHiW7+K6VVnF3auxiXMKs2etLj8T+h
hvUOvdZ88KbdaXHKCqQ5c/uu+/MnMLC5YLoXBE6Nd2ahDsgOe0DjhH4af/P+5k1c
E9H0E1geSA9jYjoX3skOSFbqdETgRJMz50a3R+YyJSp/vb0DkUxPiN4yuim9Rnza
8sAe2JHuFwGZlxyT8rV3ru5x4z1Y04kBZfvq65rqgrmXh6KGfbMXQn4EFY08FJBi
qV/Av2+nVFOuKWiYdcFvAQ2KGl7jzrE3A700Uvxoda/+e9QVZVjD7IzsfWGXvnYo
FkcmUxECKQPenqnE/bcJ9NSmSaEn8Undnio9v+d54KEkEWsvOveVAePTP/wXAC9E
Cw1vMztiM14lU50e59V1cEEYShyeTIJdVEufNNBkggfDsJQm306FCSLhEM5sDBig
5u5i68h5KV6btS71wUi0/QlFAkolSHOh8q8Vs5XKvw6p6FjFoxqrc0BIB0V9x30R
BGT6fqe7Ajzg8gQd2ISVszXU7Qujz2CbtZZEWLzHm/VRRdug/+WBOS109bbZOgSm
K/yRYA6Xi3FHMiyBhxD2xaof7gs6yYDA8e/l2/N7CTriEGHhwx5hGDy9obzMQanM
J1h/bDjAGE7QncFEzG6PIFE/UWzmmOqfSVoO3bFXS+oKlmad/pAst0dB6sENYRoA
iM1V6TD6pmfwfW3BpqIDZU4rRLGnr2386qjhP0h2eO/u0fyqOHTivTkC4pnl7afw
auolJe9XX0ESjlMK1g4lObo0BFZtX/Cc1Nha0K2T1ElEO6lwmycEIROa2Z7q/hRw
iNjrd4Hkg1/Ji8Ol0Z5ufUS58uscmPZboo2BZLZzhPZK47k4QAhb9NI1G73w7yp5
OmU6F2hmry7gOS5dmMMilHc2wcovyw4ZdYZsXagUb65ZpBrQbx1uyMuSBac0dIqd
cXx6v/iXmR24sPeg3/hfTvz/HA7jTfhJq+GRhvD547SXjZ/AjazbxHdxPVyrqrem
4LdAUfm6N3vg37c95DQnJ0Ibowwmx9a6mAHtoZ1bSDqIn2MUTmrcjWm2/1zt/KmF
FTV0PC1BkAlf6DeiwzD2hqti2mC8VF5iWk65q2f9ZfChGE7gRsghtGFQQeaFiCjg
xgJBffoDTjJ9C7Lr6MRi5y96riWvO7RjwreWKWRyxuycf1vPek+EG9CtzASP9NBq
l2UFweq8J+Wb/gT8C/2nFXAWkSbrQ86tGnDxaPh43/DUMvQ6UN3xMaKQ9q0EivH5
/CENnQ2X+AsAoj76O7ELw6xsciO7l3arfhU73SmPPnNNDEIu5vJt6T04zT2lwkCq
Pnl1j1HeJej0L6WULVuRyL5kCLkpn/3/ohTYt94JpHNUoyswauox2Y46tSlUsIuU
8mQ4Coxpx8+TmJpEUmVyTi04LnwfFunUfUYVhLfGSRAYUIv6kD0iZs3bkAdaqczq
QMjy0zRYNy5SwgXSEFOzFaiYnf2YOBhtTOUNWqZpDdBD3TSrGGD4iq6lilDNdYn4
f9YhKYgqCwmtlmw1dtmd3mfKRmJb0ysDSE+2iwDCCqy/VGJ/x4PgkrReud+Z9Epj
VzIjAxQyZJ2e7FtFgYlOkyNfAV1PEax8d4zWy0cMqI+bo0tonxL7CFUgdqikIAoz
kPeHIKyATJfnwerupd5qADYpazGnqAr27/w9YIH7+mTsDDwCQ3C1rQijMrScsUbb
cu+h0yjXy0VW/SvwHTtnovmqXvU0PfJKpTyhoFk88UbsaMB+h987BbOwDgJWtRim
EsLsatSwoMYYOqAF7X7/GNcgOwdS6+8LKjl9bEP9ILNR6SC2E9tUtYhAegjqEXKs
eJJm5ERfOOtqfCxbs64UEOcdtI84bGx/tDRfczVMw3Mw1Wo/9Y1Kzr0ZTPbOy6tw
AN/i4iFDuiufUwvVx4jWc8DUnJ5mC6vXSqodWy4pLfhj1Omh42BYCQyjFnb1mAWA
5YSPItjP7CcUtHL/cMKz4W3B3SEEo6buMLA5jUJ4cO/HeylEFBlNnkh17nKJSP50
fH2coLC9MXQ4ikA/RnEtVHkkYBxdu/wGGdUwA3O9RonwZxebxsufKmmqdlKrsQuk
EobrUrsrLTl3uDEaMvKTozzqqhqIq0Ss+msNwE5bzTdH/o3JCrWbVUIkogpsyyfx
CGJKjvroQfRAp0AcwzHHl8lsrBmkpT7el3rCVNFF8hjfcCx75/lwZ/it3beVxfsW
OcIJox4+oJOAt3xXNeS/KxAwh5lyKt/uEUtH/n8F0Z7YGSXaRA8lamh+AnbsdwVb
bGcxBr+13c0JZ+1eHO0dTd6saHJkhvokwwePHFKV1WCGHDUWwJ2rBBEW0RWjS02q
XvMm+jMr4qYzHkQpakch4g459RATc+hi0636wZchHc+F8T6q3r9gdkw3dlz7lNC8
NXLvOnqcyOdcVbOHmb2VZA37Yymz59YOOAEYTFeKsEb+/TiagZdBavNcsLjDHXtK
wlzyogBlzA6voPMHSDtSGiEdOuhKcbJ7dFs2tDdL3Cim8fmxBTkp6ym1ZS3DZ6FZ
Dc1OD40Cgze8Dr7IwE/Qg943MtoSIqBwaj1DKUhqctekrmtKzkP740TowWzgpzDM
rg8GNcJIkOmyl6CebmuP7az4etdtA0nP1sfLaSIKudzrobpJB4+3W2JYknq2zNL5
GgS/uedDo7lTejuvioniWzJSH/9n+NJlPAPYXMPe33IXocmu3ntX62NGAt68TeU4
BdM0pA0O+Ly1fmoj+KBU8FuZBLDwbMaLCmvc0BVXrGNnE76t4Byi4SL1EMtjTI8g
JBkvwV1cO7XE0ovd5w3rk3vcv+Z23r+ksDXWy1PqrW15FBtr1V9XjD9zWXcKglyQ
2H1+DmOgrF2nsQR2EeQCej22T9BXTroTROU/+BknU2c4/55OOKmaoN24Fj3l9/Pa
RREHRy/SgqLxt5ItBqJxwfGvAcWqCQ5hDCZg7eplRlyXQ54vee7rvGttWv1gj8S3
zQvd9oMHPaPstB15oh8bat9zwJJPX1d3BaOvsqglp5K4m8THWnF73kNxwlUK66I+
/tNxvxbFoVej3Gx5UrC6LbZvPbMZyDufsfIZxHSABOQqMILBnqtpwR3N6quwpYGS
Ezg8HF8pCSHHKTdI9xx1Ls0omfZQtOKQc9lnNrJIFm6IA0W0lwTrlahty3josoF5
LRpJ3dB3k/yCnVsUVJ06BpxQvlKAriFxyvmVHs1Zv73RvZVY4lsP9+xIIDzmu1Rs
fTtH9pdjPOZQv8iM3CcfRuhfUmKrWbrJjXOyUcQ8clOXvvqdxqxqM2OF/Mb7/WtS
yrzwC3cS0n7mCOukqXj65wlBIDtRRo9fkQrZQo7S7lR+YQCW3trs/W6KSL7WYK8Z
wZkm737a2V5miMV6KuPatGZUnQvZpgC8cUd4d81qG9lLkXwONMoGSfkkRUsGJKoW
zwftRgcC9XlIu2KnL1Rr5LPCwgy6+K+ww5jLLtJosjS2Y9IvD4pIKyoi9IRC6qdk
OTQVuXzlSwAzdwCVMr3KLQ/ZP7virsdLGRjy/el3CT8aW6OAMrSGdLpugtEhSOY3
ny+ayU7yEPx0FT2kmaqcs71gXhnDxX4MFsx3WWj/zB2quvI7XKnLQwKhdoC8zIIJ
g/jSo0WpfXL5EQ/dCmqgOalBIuTcr3gyKmsLbcPop8gPdt4y5y5x7JjZzTcwYdaI
fPR7hftVsm0Yqf0bHljfuGRpwEVnKyC9kYHbPaeQsDSGbRmph3DPQTrgM5A0VDLk
8ixn0cZLW4oRhtvuI8mBLz/fzRhWujf8LydwHlkRJb8rDzJ3YOjkm3QtV7K17qjv
dmS0ZujkG10OlC7/BrtgyMeo3F45zCH0iiw1fqJgFyZpzOpmCQA/W+eG3LJyns0H
d0OvT88JJjc3sPP4ZKX5iJI+Bi/gSaMQHm7xfXw4+DboP2P8gPxwv12ERYzJ6Q36
DqBSZ92bCVzKp+29Ehh3Gso4TJE3fvNELkJIXZpDoOkdAAPiCNvmMSGrhdLsCkk3
/UgYInhi6Kd4eshNSl9fk8G+tOGolcFnROGLgXNsWFlS/cO23sjUEy0JEDHiF5y2
rl4jeiC8FeG1nVih372sfKueku5qBdNHc6G1J6lDlBSzFbnLJkE/z1i0ARzKkvdo
L9a+13GYCj2mXTaCyfhe2CmL+jvEK57OiRVBDUbY9zy9ceo0ap8GHLYgza8WjUen
z1d2O+sznUO1yK2OGVPsc6ZWsgOVaBIDRN5YiVPVgoZe6S4PfY1iLZ8Fq3PsXMKM
swdR0AFiwb0dInZw9RMLdYq0HPe3hjexPY//10GOkTSDxEX+wjMd2fYLdHyU5abg
s3z3NxxwGegrqzcUzuaYAWfP8Kvselu33TdtKsSLM36/Kfn3p3hci6Q4FzbhIZGe
v8FTMn2zgDCu1OLWxg9woMPqHdi/xbe4s46tjKbrTa5ZVI9kbwOlHUzLeHT41VIc
Qs3p3H+yhgCEg/SqCTd3f8y5qKf7ZDl0lEfXHqzLc4bwasgx+Fn+J41U+RqZXdNB
v8mQIKVZKIl8ZLvJ+Cm5RxryPtsbWs/r77LYLkr87tPaH7eU1sWeC6vgw0PcsxP3
4wi4xpnMDA0kUpc00+fPDMhdTncjuR1vtn8zauGsEbkiJJeuKCW9pe0zXinFtuaW
vgD4GXuSBzwK76K4CL+Wk8N+Oc+HXiEOwh0xUyHd/4WaY+19GL31cApa04rMI0Bx
+QkrzKIakbKNnPoAOf4jhYKM3HZXAs2xKC0tylLyuK4oWYy86agXxJw9rI0zH0Yy
5vkNorIv0jwMvgFbQxZwNoj4ZCA6XQkN0SIpQiMUG1vHMX7E+FlaE95YPSdz7mzL
KYQ1yyh3I4iw1O7zAyqKgKpS4H9Lb/ggAdFFsXvEiAMbDVp7y3Nk6F8TNQC1THVw
LATqHeDUANFvM4jawBFFcJy8vu5p1K3hyvdI2WvwWizmuuP2qQUYEcpmGZvvuOvG
81DmDn4MLh+3Xv8d37UhVRhcykRnLEDUy0RU21vY1Ctzgg9ZEwyNxmnx8m75Np6E
YoxPm/mw7gZSDpgqkLYPv1hgVTYA6OW2GEeHsPD5MhiIYdFP29hNRseiqCo4GGzr
+bfRFvIKpNfQ9LZ0hhHXDnLvc2FsHx3WAeMkG5xNt5y5QNM84iS3l3XaT7br8X54
vN149hA+Qzb2VcR2sVDoq0PRo3SU7xkdG2SAAcrchglYHyP11POgDbU3tCArhjQ1
cQf9FaRznhpqiQatbJU8S0fVr4tt44Z+p8nl1gNeWn/903eIQm4Yz601hvdbix4s
KC/CJ8YpB2jnIeqpEIKFY8PwaUcqqBfHIYNnlY1010TLHpHK4doog3NNsmjAiW3s
aUIUIGwCcFl4cg5JfXpgW+zuq7YKgRFMaJkmZ0JB8Ag349Cp7uSjmVJVIPfQXGEP
uDJb3GcJC64p/ggC5nGmidZcJ6qoAbKTRo/IzN/SBTDsxe9EA9l6fRLmwLzadHCN
w5Cn8T3NbAjXwuHpGfqLkyTicIQlBnUnD5H5ukeFRGl5xfq4PvOwCGsZMd480mPR
6l4cZFnJ87mNhthDizna7gv9Xykf2tQjyFxFRay0LNYXulMXnh12jA53nwV0GKe5
wbVa/FiIj3qp2F6W/9O0JniWKcEtBbskpdxHEn7/KZnt3hmt/Uenm4egKLmwxg0V
m0VDHrSlXjIwhY8q36oRR9rQEvsfDVpvQjt416hki+PBKVsO6/DAYHOTowC7TVw9
BPJavZ9TTEA6e6qwKa8/GunTTxhxhCa9tgPxcU19SiUiJtjcs32cZxYgW2Vjx+Xc
sh3UOOT0Qy6YvixyN1iIh6pyvQnkFFXFX2tDWGGRGbny1SrVddQscSxYFca16436
n2QFzt4aQmEh7ddsnJXYzq0FLsvWRTCELnCY2uEHjmIPKw00ujqRSUjP9iLs8zAm
NbfYUwhInoOwJBAlCU+sKgAIHie5rXN3Q1zPS2S8Ojme3jXcMl+X2aopHJ1g9TyX
4jxGHFUEiutSkiCrMfwu+Gb5O4UqTcwlo6Np/YrpXnmzpwv5IMEwUFzYBeOI1xCA
RSaBesvA/ho7jCDVFgZQbT/ovGi4dCH97e9b6MKATT49KoZfrTx9X9kiY83hGvMk
A3nszPCQ0c1Pb+h1R23O9pQpRFywAB6eO2PMoQRkCpodpbjog9UsqAjYGhBiI2dg
OmMrXn9oiFUNiTsHY2EArVQvXwQyEaxc1cEWW936mvezkpt1TgL9ElC7cjDpTsL0
3dkSzN9EecWNBG42FziKDr+fdNvgaroOpQOGCVUoHwG2JeC06BJAHb+tk/9jM3uP
6GwoIvp+YdClB7P1LlrO9jkJKZTjguBH3lCnJJ4FlW+aFKNtVba22CfTtExLI91C
V7NB/aGlNLI/jmrV4iZ8Usk/ytJuIaLqFWyIbYqECN+o7Nk/3daM7UoCaIz6/I0K
ZPS2reNnyBNYWcUb8BGm10usAp7PMc9n0g09MaIgPHOgg1oRgLTykkJNhvdL59Ui
nECBxE9KSLtWa/PwamyE8yv0v62Vl49sUtZjVZP/1ULms6/PaJbfvLUu/bErcp95
GqnTEMbwA9qSmxodbat3rCpR1kfANGL2ZZqhoNilpjZvFbK3v/PrF9ycLLLfS/ji
3MRG8e5YaeQfnvioDjLdcooDJIDGGp8V+eHfT4sx/nroQBkHRoSu10NRZPxRUdBu
NSwpCDsQ4seYQp4wAjiUORC7MP2IQuR874PJHV9SGqcSJUBpAhQPflRlZ4RQ5Gis
HnfJGTwvS1ZqEWMDwDVw+/UDU3/ncd3Kpvcfd4aBP3m/I41yLsD/z7hVRUfyMM6Q
TMfa323/6PdpqCJvTd+kpGLrwIqa6eMeasZRWc2gIB8urnG52m+i9PmNGeJkBcWq
hNm0oM+TocrmBGz35mAiuoNHDQdIiPcoUtdCgq6sJIV16dca+FmD07WbYCCluUku
LPVu6Alg9PX77agpBimw3N42Ug1G69pPj78HanXiGjP8dYsWL/Y6700vBCAGGc8J
rQs4cT0/gJcCq4iZU6xSHFjjjaLe0Cbr741ib+ZbINw7KdH1npztBeNs82VlzDzN
YkXHjFdQGjR19XhC4sp/RaSDGAMf31lUFjtcDY0uH4u/lYTMVm+m+U52Z1rLeDFr
mjm4Quhf03oWjtOE2oTD5W3hW1vFfTEtO4tsVLrwLsHeRdQ4p6wAd6G5zZGXs8I9
D1UfyA13j9mV6kZFndzoukQhOBSfuaH3RsnC1nB6XeD9l8zrrU4ReskLIDVVTHHj
RjcYE8l0jz6BYnFwIaW5xAhx77/Ykets0WTdkoTkuu0XUvLRmNYs9b6Nw1bG+d9M
cJ3tH8b2GePSHWzkEJyFCwVzzAddyT1U80HV75a3FcC6kThBiT3FjKZin2MgDsT1
E10SyVMugPmQn1UH6Ybwgjt0PeHEWtvTvja3l475N9BfxB+vVwxNqJfo9aUV314J
02gGsNuJL8IYBfU/Ym3AxFf1KVP2gPeGmjhywfAWut3H4fVJSeeBCQRsn3v9FYhU
UlEwszbstn5SXutyc6It285p2bmKFEMXUAILWDai8I5y1mGG7jzapLc9YYDyrGbj
uH+BSS3qXzqZEyHcf8kCvzY+JY/tLWGlB1trtIZ+zANS1Ji3/xaDbkAPNt6OiF/3
RHf61GrTJT8CljrfLQ439diKmyQVjFiZygg2kzrkw/5ViYhFO79mbsEjAoMKAP/q
GI2gm3JQf2bsoH5JX4H3qqxjM1dlBZ1n93wkpK8s5sSEBxUr3nOet1xKLzRQ8bSr
uVNi4Gq29RuczS/L2DqjPuLeQTpHfWWeQAyw7UYcPVoM+4g2siURp/JmbRdVl+sV
hV3cDmp9Es81Y17uoGwusDxHeT8PaWaumH4GPSMlUNeBEa3tjKsSOZ5PcAaV8OMV
6OrVJN6knK6AhXSc2/ZArM/I0EvOP9CZ110Vz25hgDwaQ/bxd9ApG7wFKEBpFzci
4tcYGpchM0n8alMV917iTseXf8z6SbIILlhUDXNDrBCJ7Bt+kx4ReL5ZFhtzlhJc
KUTUlWGW4JXSU6dIW+Ovj75x04Yg3F7i20iVgobHnCsEjioAqjkFArzM39k4vvOC
Vk/bVcMo46NgIlJTbsrqHgcGIgjW+PwMCnXm0vn6f7I9mfFZTIYhRvSs/ipeT31i
ePVa0iAo6CGtTg0UlcwIzzb4K/WVIMzwKUYB844o2r4Z2MyPBI+Lnyvl5aJOuQgw
WndMpQS8vvW+nJ6XkrIHmieMUtby721qheJGulfmn2vuBzXmxuj5T9xi8ki1EH3E
yPx0RAd5Dae3HvLhuoU/b4JKVtdRO2iNsvKxPnb8MGXMs/WFLpnpHtCVyqcpg1Dl
tGFovoulXk70NIlWV4xjpLkpfPn/X16NKS8x7wQWAHY2mGZ2MEHQ56rSaMvdSE2x
H7Q9e99zN7/CaO+uj/rTMFs3onfMWnb7ghmHV6P9N0EmW8QDBOylkp2so17KHIDR
NO4gEG6Hf4fBINL4HUsar6pPp9R0qEYQ+8IDltEp88XgJqD7RuDbsuPeZ5m4LfRT
Vyq8Atah3gYikC3dF8DoWqDygzdW659J037rF8JLg340HlvFe42ty4IMiBk3hXp+
F2wx8vUo6n/KOpnInXjRNP2wJBSQzjp3UzzoRjCDcyN2PuBsL7l0Zr5FqN5eDSXS
6v4XkKxRlRnFOP0rS1Q8aWNSqqNtOVqX07ykS0rBi30vFWOWrsd5zqPTBel2B4gK
YwQAnv7coJCQlkMgbPYDQ76x13DH0sMip2I9cx8EKLUvw7JXdqEsYZmD6wthqkvV
n2JASXznxoC78YpcZCTM69Z6Q+fI9J85m8yhq5Vrte1H1/XoZVYYTQMiAk/1HGVk
d9ZH3WO7YyOB2dWElZM7EHyjET63QIrDg/iGrXJyx6P+N2reUEUN4Unak9R+vGmb
4dk2uT1N8f0I5eIieRQJsPg1oR/hzvEP4lZK0a4XyCqcwpDE3nCRtO1PoYQ4w6EG
tr+mOl0XV/RHEfIW3aU23SgOTaMgjtI/InQRVY6cagzz5KM5hdp+haUx/FcaTkM0
CPKU4CrIkGgvPNVpJ0dsJ9AuKTU8TgqxlCP4bndN31uujvELTjGUSchl4Mq1X0p6
gDaHOIo7PuceYd43KTbd1qWmzQ0Z8hRHHZhPOAlJneRjtQ/gcbtVmTkKI9LGWGa9
erFeceGcEbGW+W2a+pJgTkFVD9jz4pBnZQTnrzvYOrdzTgjaclp9IbrnaSMPgv/a
/5xpL0GyNuZx79WCnv7Qu8mf87lYh37PQ9k9Qen6mqeIj/xKF7/ymMfp5jSlw1E5
QfpZAAXr+k/Btlqo8zdB9SFgVwkXIIgVj371u0VCdrWKy0nGCG19e5F1G4QNMX0I
MAGksYVVSm8TJXXzjHnwGt4EuMET7/EfpvgCTowkyZtXNOjGNl8CDcHsTNFXdqKS
SAhs1gx9JZ4B7KcMno4QQrk4TKVSpsrHkzivm/0E1EyQy6+QAudEU8OmurjZA+T6
GY4bDs0eF3vD2VmwJG3de+culp/NNi1sLBHz8xbCg/H1A2Ni30Od70wvHEf3AIld
M3I7UfkSOMQDSayt/tDGD3WCCWZpOoYSvsneiVINvNFifB6ELkWeY+pQGkZH+TzR
3YoBoS+UoaZYYs1KKJqa18KJGRAm+poL0qvNcchTZzDBuOv2sxyjeE4pCf31zI2s
RGP4igPLy5XcI7uGL3newW5Qy10tB8BH8i2Id05nfFA6pi77XT/FU+fDFCp47k3T
Py14BZ3gtG6ykSY/BqT6u99mxkCR0mlqzCTQhov/BX+7uK3jieseK/EG3XqGqkJD
8kkKsFbrRXcwo69WbdC21GUQHgXO38irLkHwC98mDhd380EqB75D4MSrWKM1o2iO
cSmDnrUCVBsgq4lrZr/0aVs/HTmO7InZKuH5BOvYpBXXMwUdFCH4crPO5PxQy+tp
xrS2EAPVkoS6fasV/ZfGt6gaBJDahxQYpjg1PMGOMUQk/OXWUKe2F+HCDi/okiIU
+9hZzcZPY03wtg97fuLDlckg6BwYXNE8ZqzfvSd+WxlYvY0l5r+OEC5o5NLoQ5fA
1zIeGZyzIyBmd+6s0hjq1dm8GWyioWipFpIB979yUULoIW0TB7WMn1Y1JzZL6R1B
Altx7XCWH+AeYVmDxogqLAZod5rDe2qnXp49UoffVlrx3zEcZUvpAatQ2QUe9WOI
P7WgHiFJDJv8ZecU2f+6jOpV6oHdzStlacNljKQPtwHnw9Xv9ITv7KNyIk2GYSME
mPNE+lemff4LCE1KyMgJob+vI2xvS2utTtrJqw4MdkDk0A82LBbQ3P7Vr+9+2His
Njl15AgFbaSXgnVb+4IUA71cqnp+L/qss68Zd2JesJH/r1aBItPBilC0r9Dvvigy
rg7novIdfm/k19QujjEFmGIzLHHzVUEMeP3/epn2BuAyRSLUDmiJcfHcNB5XzQ/A
pjCfZLXVRNET4NsimxvAoJFE4MdvDGG279bpWYcup4i4nAJBLL19f5U7Pwg/cgIg
8+IdzyITETRcK44aGh+6DB9LeAB+ipBS9Ecrj5QVGROX37sww3WOvashZOa4PE8E
+OKjJVIY52+oUAP10xw3GVt1BMNf4ePsrWXwNWB/EoUYsXqyQrMw+69O2APxEH6L
YM70eg6ugdHncxjoAmBqs4RsNQxaOo6Fv6G9baOUaZRocvS0NGNNVB0C5xXrG29Q
vLzMneNoynfzaG1Y+KsTRJ9CNv2+OkhbCHRclRBUaZsKbFHLQmfpAFGbqWXPYTtf
bCkUHzX0FT4GOYctWjUDq0r2uLBGuXL85GjogU6i1PJDJfIhFkf6c1X7hmGFofN7
F0FtZ7akNXYgS3M1YR+sn5FtPRB+QMHVQZOk3DwXs5TVoBZotbH/IsiMzlZ2XoGH
OiR5IXDMucswRXUyl4HxIFv+NVx/B1AjJTMnPg4OluC0J4Jl3QzDq3b4gRPG8nOE
EL4jXsWhfC/zjfbxrd5iVPukr8Zm7krlINWKap37S54+3Pa1SIQDoVMpI96m0DQI
2xCusR+8oxTG9+IB/Jr9aKndNFQLWzYUSghj0FE+z7fBumiM6IRoItD+xEX9PXkc
fkKjnM7BQvYeSLHv1m+Wg6UlEjOpXuL8i/OqHa+kR8VxxW+lDeZLvYwvDmv3p8bn
FhoVI+qZRaxboYLY14QAld+pDvRjwgVeeujNxXRC36MhFE9mT6XvkUyIQ+ws07fx
kyUgkufR3PdEbERext/V6vUPJcsmmyhtM3fM1jXjoF1JsOZqhQsUm2NPxHzkp7ek
FUiL0hgNVGvWU3WGbJRySl/X+087Ttd5ATAWNks4VOsEjisN6WHj6wn+ABWV9HXy
XG+oDfnFCjKdc0W9LAoNfEB40imgoWfaJpMFkwJmFk5PSvKAqo0h8DC4oV8DYuYd
C6LxD4ZtrzQSSgF2KSxqG5nQOlPG4VCi2XuHOPTwGkaaJxtRSG4SaXnpuEmpsTp5
UYvzTZ/A6Mv9z90U4DjVfmq6VF7zzJKrYZ4pfPdz14R0rT69yqkHlH+qTXTN/c7Y
SARAAsRM7VoOLJoTzmi9zwFTi46wm0O1OiXz4jy5Mave1HazYCV3IRuenlcOXrJE
3aGBKZFutKCgPMTUVH3lre7mQyVitpVty4wmxiaH4IF2LVw7Fxz28rnuZ+9BLjCJ
wr2lRnzI94G0yifwhVNaolY4O1m52BW2tvBHyTarU1bM4Aew9bVZIOcAPGvYgZrU
7xzU2I4khGfEBr0kA9yvyG2u5cWiRZhcjzzjTjPYA2Z3XB48cJBUiu+0LZLqkNnO
GtCpsozaK2neEaJFmJrugvClcMzq5Bi1l+H/pW8ilgloF7hxS9MMGnipJSVHjhI3
KC/NSKvruzFGPHDmQYL4q3b2B3Uyf8ew0hH+D+qucJHsNU2X/Yuzn9t8s9YiDMD2
lyVhkNthVJqRA9IWweDkOCYITS5hixA07MyyVHF1neZNym3PHSWqFRysvJCe/Yk9
r7JKwePj2fosuKEw9VK0ncZSz7kxrjjAaHTZYbmEB3oIF3XpbGHzkHiTAVATQSoK
x9kMTHx2pU1sAmD6hew+UYR2NLUnfBvg54d7TCNiC/rerjGUQC9rKSAYTJ61FgxU
uh62SKW6dGeGBkSkS02JZ/kWAIGOr3SMGJ0E+scQWxxUf2JYXSFHxYA+NTCYIhTe
WH4oTIwDI6hw7v/6XuU4J/PcX/9ecK9WnhEZ5xaakfb2uGUbh0VndBxhaALsy5Jh
lFhoW5TWEQsJUpwfadaPGGYsF5vkXYAuoPzay4uIuxyG2ElFq5z1JaMKF68SP4vM
JYuRM13uJLvBMXZxjovQEnwBETOV5foDK66vPoiopE/oFD+tIS/OYOK3CTUJXiLZ
CRI8jnv5q3xzKgRNMUyrPChruN2Vmai1Nryk/GT2ErbBhiQ/vwL1aiaqat3xxnBz
SWpg5ap3JCOHMGBChJ+BrExET2k89thX+AprcwWrWqYg/EbpcBIUYXAQv01PMsgE
gOYZnBI4PtQ2NQWk6Ax1G51KLq+AbzMML18enjylykvk/Zwyz1uW7cXS2RyoJoSq
AId4xj+R4HZDN8IA9Hnwe/0Thj/7nMIn0dqqXU1alkQZTRDh/dOFXaOVaBPRF6JL
JaO6mw8vKUEt6AhN17CbI+r8OgLyyr5kzNiPDPJBQV94eKcLAYaPmtVDclr9jeB9
WtAcX9v+w7kyHa88HxOOJdagPymTnlTpomjjkePw7bcaWzr6Bcwavqci5Nm9rmI/
gtLGvK7dPzAAktBKMxrE4H2XTEdJDkPlClfE3/3pAUvVBHtt5zOhcvi6IfjpoWnL
CCRgFHIS0b7QRNXxOA2aGOdGYlk0IXxhKbKop8ya59Zb4AFATvcSYFUhJPX7BAY+
m9zMSuz+IxBThdTz8VItw2mvdEgXNG34QW0pGADQTNpFsUXEOqlQxD2chwrR/4eh
IUQrQ5T6m4U6CUSnmYWSsh3pnsTbKNO5RAmErkzGT9rpQM7MRvt2693y9g1W2yL6
wmBCzUAgJmy/7mFSuczGfxpcWBL1vI7WKnM4wsymswQRH7e6QeJ5vR6iaTYxW/2+
5S7iyJ3ahcvdombiMnyEjvVnRUwm7tM/uDlJi83LimB0fTjZlJ3IFt0Pa3RgR9Va
cNfW5i/xRpBgQl2E4p+0Frr2oTxRIjYzo3IKFZI3urLR7k2qIFvvvEUpLIcP2B1N
gH7FA5OH9uI6uO1N06q69ySVB4nGpPw3/kLEmqoOdtL1NyZ/BROqmHvL0Gs+fxoT
wtPr/0NAQQOtA3FQ0ULbTOc4NbC1cMQ+X91clEhpRqOfN3SPPJZzL86iIevJJada
qEURpaBwe1Fs0Bu8lBKetUXeA+/gao2/XtFMC1uXwnDe/OIC0MX92qZKeHPXqDlW
5ElmHjPzZQ62nxCeLo99GCQIXr24yXU4qp7ONxvH1XQPFK9k12Hco1iRNI6rJ8Vd
e82fdy0clPZ8UMA0koFcYj26QloCcjodVww4/QyUFfR5XFmRQhQ8UvceCLgUmYmw
p0zwZ66HpVnBEBRk9tJBTAJHSHXyhXXLUHaMY2A9i7d5vLF62ZekDB7XZK2szgj1
Q+CbferD24OYrLtzcDsyzTe/8OwvRRpCRnVN3Zwh/vaWc+TlBWX9qXKdxk5Z5VwG
MTv6Mk4cM3OX1tLmEgdNfPbinKkUxJ5sPYiVSxpOeG7QKuNpJ34rVrdWUouPEUM2
Et2XS8wL97HZ0szhITwcJMRzUkacKx/Irkn+a5c4Ffo7+FpbC54jksV2gPo3kf3/
lcaXJM7+6uH9w1vN2tTLImEHK3zbQ/hbVxomNJWQbe89iylAv7VFegrhvEwtpk1b
4KH5USF/yl3e3aCK3CT7BgVtbsdQfXkMkJm6329yrpjj0iYOew/jJNz4a+Pb2TI1
GrEkf3/oyJ0Dcrt/e8MEvQ15dN1g2a70OYACmiwX1dlQqPN1zcHARr3nDeJxmqcc
3yhSzn+t3rFhao+nXJSTjSgU3uIDtXqxfrUoXxs5Nt8HY+v4fKzgCWJ+5j2VW0+G
Xnnm07G79Rny6QVm6gDDfRZ7z/Y6CS+h70yHvd8/zeIBqT7CV6a38LgnAOWFcCg2
HIZBTGHASJmplmBT4xinKoJvEQ2E0cGHK/XSa06IQ0Ttbt1eOpr6FAiph+Bjv8el
1tA1eFazaMaprmXxFsx9v5XkJxL7xK8lJyq7XeSIACLt9BzomypUlbs+SyPEFrjF
q5lAhGR2rkttJ4/U5FngKPIMPeZe+szjD1FIZEUBrupCP2BzhpRRZp7k2/LdaWcc
14aWqfVaz8ubYmxMZIWushPw5nNikb8n87jU7ofzCpIuX2brcghlHgkyIP7vgQuJ
XOgL204a7fakmHbDHaz80cwTZbhtf4PaOJy6o+RclMjfJMeBhD0ajx6xLeQ2qaU5
9Mio3VLeDe51ZhOmsPAV5iOThBYIb1npjj/FkCP5OH/qkcvxj4EH5Vy0aafPdq6H
2yblOVL5WBSj6cHV5UNYL98RsF5sj80WEPmGB1UdoeIWnbaaJ/CGdcLSxuAuHWkw
mqmOrIlgh9WmJYwf24JrUhixci0X+90WT5UwGDgjrc8Nt6rhymk3XGtNVn0TIkLt
WVtIzfwv1W9IgFbKtGxHRyanONaRQN2vqXRjhm5o/S36l7dhKBx/2JJpd+DkIKJH
STeN4yITf1f4wANrYbpYwwBERtIVOoi6xBBGHYmrcfpq+spwsqdSmhsNNrFx2v2q
cEr94cQfuTXREU2eZCmKUQs6wG7vC717O/xJDSLCuglmlRAgh65zft45j3OcWjx8
Btaoy6VEVzfZcx+rxNVJubkDtFM3Wl9rqtBE7YNvwjdFEW+hEtG7gnpsCp39yyyT
TswR/NNF3qUsZwPdIQ43YdSsT8HXgie7uhSEl2dDmvwd3E5RfBnlbTfonxt8Gi3x
w4mmBOMbP8ygBl2Jv/jqPjcSGYN7rIaUW6Zub4wvzkCL7si3FhvXTwNWxzhy+slo
Bwjm0T1VyxMTwP2ZLE/BDmzaK/6INYGYFzs1Dg74qtEG0M2O80cBinQ4Ev105bX9
sERr/S8LnRaeedExxHOH/cVGCB+d1NcM4eaQLBlzHXs+yY1mTm/2ypcvmwJhjJAg
0OH8cqdN8CDmch5yYMhxN0YHpzIQE3158GN08fFD2WI1Rjp8ii3VGGJNdhaTy4S4
9c5pk6ww9ey7wuEbgZX09VLIGhn/QBD2tV5lUNnHe/lS8lUY3+8laDKyuN8dUxEm
4Pfdcfl0UAqx4jpi505iPwH9YsbIRR/9TgXO7u7aHX3nCcENd6kDaWJu93kPfku7
yEDAY563JU4n6Oi8eF8IAFqC5BdvGjVqgklEKkZ8EeVH9CKVLmUXKkoN7QjkcXK9
+Hw78Hwn33Q01R4SZro8x6jHA2TRMJmSz713EFuI5GgNXH+pqAVBPlCRHjnWGkw5
ezrPWJXFsn0UBMRi3BS2RS0nEZ15x3au0N9sJCvact0kGvg5xrAMpgnvYbfTBKH/
s3M8P7tP2hE4oztLGmGvPEBGOiinb99FbH6phySrKuRRDMIKQIy9busslQzZFuxK
CiQsKPsoiNirTHWdSRil3otOMf+X/BhD4ZY/+vvtKuchO14SdcDpNE1ih5ZNH2mz
rNHPeENZR6qe5hBXoTieDvT/4kuMrmeHTZpWXDft9D8KN01otsWQIq3XnpjNCkit
zW41j+iXEH6wS8Z2+Ovkt+oSr2M+c5v5KdQBClozDuvXXqFDvztNC663XrNmxEb4
GNLbv4apErOFCURfzXloJ8A3RVm95dG5k7TPY+krpMpXciHVl2gGgLc6VO05l9jS
FuxXWX2Y/9o44EnI8ILsL6RPoFgSwpqqMFa40iVgZQJYnEct2GtvfQ3xW9JHU+QZ
y78q4GO+sEAPDMVROcScbRlZsjCnohDFRZlxyAioCNLIOyKtzAVVV24QAPH7OJXQ
V4PtFxangROChp3gWVfgnC5fmLm/EzKJItvcvUSYbD6RRWBRtXtCU7MyoGDGDzYh
w+E5H2wEfAOCwfd5zTufU31MTTYdJFE+qu1kxkitjSIoUZ4c0k8Id0fItWpuuHUe
LNdahfGZWo4w5UKlNGnN9L/EuLyzol1gg8ibImINO8yVNKomOearnqIKQGXX4jax
5nfi5pmjR1cbLyAHWesdXY6wV68rRQpbOywLQXGQX29azhX40jFZSXUfa9MFyUxN
T2n1CF/3o6sSLmoGbktSMxDxKA6ZNWXtULcT5+LIih3MnXRHvF8hvyBiiJ2h+olP
sUlPjAdWUKqj5DlUJgYtm939czOC6gpLP7o1aGtg9xCRU4Wqnk+4rXnYrHLDB1fi
BHmtStZgdl5awBAYaNSB+rv6sQqypKFsTFrlVDQm21LSDYWlL6VTyjiqUyp/g/9h
a8v6ERBnvSMDwdnuiGyGkjQ2plAdgN9LhGpykvFlKCJ8Qtbl4iZgkHsaYCa1N0NV
NWUmMzpsVUQ98PHxAqJZLC3RP9GZobnyv5ZehTmNyHL/JMWdi3U5KEYtkFNGp/Ss
+AG4NJwu4vTT/oZNeVSOPK1Sx0L+hIUvOjrV33wAvKPSjp8NpaCPvSwM+I53y5VO
TVb2mxIMEgcZGl3CJQD4GJKZzDiioWo1rBHRUlKL+CBOAcmeRcmpV6P6uIK284bm
DYI5/S8o7XPwyPmVZ88lZcCQ+uSVfvPTsStpUmRjzM+3Dzw4vK4I0OoS4txDLnQs
dm1ZabV1+iK14mW5FSMUYaZsVAtQZYUWNpqVs8agPqev9P9tq09mpVTEtD64LT8n
Km6v+GxeND2cKetfPDY6u2eS0MafFgkSetMEdopENTR8OB4a1U5EeqToon/tK1zJ
xtAzf1vZ1693yHkNQuIAjJER0PBcGYgYhFkFYGjLG2PgPwFq8yBqhcg4hIgunzqQ
mE5T31IeY3AOdB+Tp/4h6k2hVu35CTrm7qpKtwkXNOzqMTKGUxt/+C5cJEaKBa7L
0oWKGj4sIGn+fPBn4yaBef+zXIqBEaeWlsWn6Uq0q3AQulpLPpqOru6nVg7ZlBih
f0xNAVzn5e0b+AOlRGembu+QwYinMQTrUCJzXN+jBYrEb1aldQPDuSC6YE/diqpx
F7kZ/UGe71Wp15KaE4ypzMZZ7B8CsYu0NT5ew2gNMcB+JhbCk7iQAx5qe0v5tLkV
FahYNd5Y8+3yCdDqGhFIiikSfk/7UtTtbDiizTwMON+ijEa88ar7tHcMJNcUX49W
NVJiyZlABdew58vFNkTM9y78JXkA6SaSMoKP0XizCa/ANYWgsHfKlDZi4W3XB9Nl
DZhXfxQhMh/8uqlBhEIC07YDrUmp+YMbFYFfVlPkmYpcKjV9qIExZjMm5FKYoz41
PUweyG3dmxz2cXarHezVFL4wsl8IDqhDxOa7zf41aSjVguO3dGpieB5fHRLgNtXg
ox7ovUCAmF5ADER+Lq6/Kbh8hBTAHoi1n9pe+6UmCh1czNBiWijO3ndd5UX8D+Id
KBhqzkFjLNEy6A7ru75YOkiAaKOXrSn+AsthXa93YlFNpONI1NCONX+qV+axYtQW
O93O9JsnJVegqCbpv5qjfyZ3Erg+T9BzI4GF5Q69wrtpuQRY7bp9LpHZSM5sGjBX
I8KESFitGgRxEovU0RQWbTXSOyDy+70dcEEnqq5gfLxzlSKWW5byc6WTa+0hFeVJ
GypeKWtqfpP0NY9gU2LOmGZ5UzecycD6Uo9nBI9QHfsw5s281ghe1tGOv7hucRuo
XHtIYawgXbgwJZ5eFe1btv9+UaF/inlsLm8q9XmIpRUPOqjTfwRfTPBrC3Trc0TC
ymhHXUGfEZeE0JNaoM0xUMsF4A1fjT3x8XHFO4Wgni1mX1amrme7CUwKBJk/LbCI
n4FvZwMo2C/Sy1B+bzERs1ugPhG+YjxYb3YcXLuuN9EKTCwbw6klpc+1p4f0N//j
o5UmVK7JrkE4MTcvgYYmIgCdkE7uTU4/XSpE6GDz0ZYH7voQB2U6BVXi9re3wi06
7TIx+f2b7JTf/v3M4nTnc970IlNSH62rm8g9qpycgpgTAykMzKLkTTTtx+lT7ylW
qcHhnbrNZNGAkDjXyie7lrvxXcy5uy+oW6dri0ogSuMAiEYfe9RrMbyj1FlXhM0S
auoRajLsGHqk9It5qw34PiUJ+QaMolnX2ac1VnuINGxVuD10r09nST+Z4L2WCOh+
CTpY2TLofnHEG/gAsdvecm0KvsfQ+T7wu0Uv9nqJMu9yWuXIC3/TwJbLhTGnGadZ
JrRUMAgMvalNP7HEqbcuXpyY95Gk9or+vGwOpMXULzk1atzCezO8rSoMcey5dpQV
SjuFKLp2gjLrQBJDgroz95P109sdvIBBfqKwiniTNRtX3KiT15HkffJPiPPeScHQ
0llqC19z+ARsH7R40t0XBDItvEH37RiEhh0eO1gMUSufsPHR0qhXILFyH0eAsQ2T
egp5rBH02siBV/f4/5mpGUe+YdQ/6CFbTZUqcMckNwtna72r/UTEoHfvjkIQGQIH
+aWQDrCPQ5A17Uq9lT+ftMG/+Dsxzt7cqBAF1FlUdB0QhudlRu9s80CxibYg900z
NSDy6OBsKaeQcY5LUshKxJ5xgREeeYpl3BQlPpW+hJV36FieX3aw1puq2FUnc6WU
Hxuxe4uPSaaZxKBftrl0JnlRuOBuJxBB1xhK56qmeJCE9UxtCav5QOjkUKhNaW+e
TfT4s4e/7XDtbAvQs6iqrkFCOhbbGgYPBaerBTvTFGs1bsyhW5JRQt/NmphDz3LL
YF6WR7q5CkaUfDZrXtgWWytFYcxKcbLmNo7y0Pt/2CUYDX6m/MiM/jD4ELV9OJxT
uvNfwJBEg8bHog8fGpSyNqAduul9lbokJFs6iK+Gz/nMUj9hDEjQWNZqzTiD7kuv
7Tkrk7C/fF821RkpmqUh6Hi5x+kQ7ernBy2dIUrTTyd8FMzfRTrwhNxgZWgT4rhc
AWee6ypmQ2Vu0vqFvQGCw5zmAKYp6hm9aGAot44M2nYtIClMVITbYdoz8uYq9T3X
D1MXEzAFbW+ofuluXQ9+8l/LKR/c5GZbB1HDQa5s4wIyFe806qQXsRWxkuZI+ZlT
gvCIK/Iz4qTR/dy8KqT+S4I3fPAl3zZoRoy3H5MuVjk0RPoiAVqVbmh1ORvwAHjp
j9nUx0EIrLbJhDI9pDBbyCwl+hFWd/5ylrVv1m89lU6DRWH09CF3YJzlr7YT9eYz
PdFkbtFc1ZNB1QZC0lOvbD/R/BxOrf99EZ2VYm8x6O6p2MT/lLche4kZhiRAR5fw
gdUUmdpFZUEyCB7dLqKhPau8uKZRbLCmGo78PfNa6UZMVp5mlhdK55UknZhKZ8xA
YjRV/FoFjMyvFVGTi7vwb4VvZbcpYBAvXBPXsFj5voApWN3vQc1IAMQb6MznDfpR
ax40zETnTRZmTzgFWZVXkaZiWAaA7Zezc9NzVzKBRmXmaQNAZ58pFfxSLNE5MTkj
E53KnvzdEpKxC4fdufj/dRkFDCnzOArFxtE14cEkMQwXe3PZ3oIWG/7vAREH1uvm
5RxXs16hUxdhbeYDouRQoKfzUjU8gwrnAH1Wx4fQRWxc41P7Ma91VQsJzAJUjpkj
QcdK8qmAF/JW6nidDqj5q2P8+2JQ5dMd0FQAex/SIE5rkHsORkAIilQw7SQTuyoF
XWiJgTwOqO1UHz00BgY2aSW3UtoElyjwhJhdbb4+Ej6uyxz+gTWqvDRR66xjJjbF
64sehI8H5M70bw3AMBNIPFLlm/wHKCmQgqDgoFZBZwFcvs9ybWQvKRDzepIkLqsA
roCMIi/G+AXJ8SQfps8uU8IzF9vNcw03H7Jz6bQaJsLffGa4rsRlDsSD5KTigNxS
IWmUg58qW1/AmXTCXbNitHwu5LztDpg5MSVxxNEatNt03HhH+VCMNlzaIjPTgEHf
7lxIxCa6irtUZoknGAMJ5GrvfF1e2k5IQ34KUY/M46KesqhyIAWhRjNlax0PI9/s
1OlRUA9Fb1zOI2vixg6piIKowkB1DQ6Edc4/mUGh3otK9WVkcIZELlM0Txkta1OV
BgKr9fT9Ef1OzrggZeoqnKs31aO0DdHfT4B+B6UdASfGtLMuBLWGyCVA/4gPjym2
QKAQ0DZwq6doDU78U4aSHT9sQhHzUgoajF7X0UlSdIFsZWnFAOjoK+l8B1kZIRyz
GySM6Nkq+zws0oezQDKPU4dmj+3BYuxHaeqnC6NBXgUN0WlBc3uD/e1f7kfngw/5
1HuBSUju7JT71OIOfZrgbH12wl+1GjCo4KImkNBvQzpz6QiUCBbonquDojlMRmul
OFDOVTBSwVCYkRqHsCj9yMkPdQ1af1bLgHSCcdBE3Rvx8nnxTM8GTKS3yX6At4ga
4RQicJu0AqGMAzWdlXplQhkMF8wpl3zo/rdmmOOOSEPHXld7H6KVuEJOPGHHTAbh
ok7R1IHKRGvMp6LbFeHPbLEOphXGZ2OIGzDPRbiDKOmgyueZ4sRajG1tc137n0Cb
c/LVQD+D8aMg3mbcFzZC6RaMPkQEYoo6OB81KpBNOaa4WQmrFhGG/3nhrUWDs70W
xX4jn87t5gmdKx/vaq/71OWxy7lUj9P39n5Xs7F27oGvHIJvdvFDOD96VNlsFbDf
9ZTU10YREpoVPVI3FhApMbri1aQf6odyd/LUWRSGDUIs7MOYHrdZekMaYh5SaHMH
pJGaJ/NoLtaAjReqnyahWMIpWFWvexYondT3n3MGAy4+M3FL33C6ZyYzGHEOegPL
NOVBD2KJEUiBETvMfym4gEhQ+yKMs5FKKeS0vpgfmXKR6cLTC+LFUaxKgS6Srjux
ocSKepQdu9XYk/DZ+GOzJfls2oPKrcZmeKgPIYNkAmrkTPaYF3np6CsyNNsizWmi
tA38eycG9cAMK5jiWdXkS3x0uqspoWVlZ6K1RXPfpTEf718FFamYt26fft8+9d/X
SMoxmx+PB8EcOCE2lywuxyH9bqr1lX6z3CZjxNUiofWHuU5Xv9VHwR97eszQFdse
aUMcGwDB6b2lS33S/nz4S3NJNBvZTsPu5txkhgdP0dthVW7KD43wqqF7JDItLg7I
qn8GWmQbOqD62O57aFu29feYmYT+K1HGSldly/STksGz4rD8Bdjabwpp17Rx5tFB
5k9MjI1o41M4BbW3X+Y1wOUKuZv4T6wBLLhifTBljTzuSqDmABkXEfqism9kcRdz
DC9k71BOpalKB5b/o1q66VS6MiPwkpEQJDNgn7excMiLOgmizoH0RppTdAVNqhhu
F2HelgWTTkmkEq4aCNscRfmPBcsQPuxmOlzU2k/77UyOXEzF4mJHwuRrlC4tG/ki
2zFTI0RCKTR9zODXKU0cSQfbnGw04qKGOU2UzM0ObbhWxk4iKHAiKKeYGMH9CFXi
9NgXfjlxIGmp0L7uibGIsB1FKW3uFC3HE95HdbIboZpX/tN0ZEt9pNTkqSlaM4u/
I9KdMOM+WbmybY+hZAKNbpvGCIiD7pGTJr6RGbmH83kQ77czptCbNKDNbIXZRVjV
wY23Q2MwPTSen0PX72KeLJRc2sL/FxEGF6tbzYjv2F9B/7ZtVXhqjIDfsXlQ/i+D
o/Z2U/135uOBGsUEJqzxnP37Z0kD39T0uW5aIla/fTFtJt064h1fOMcnOqpeDKCO
3IEchM/+z8MYgwmkiVXACN91gcGCCkIGgjSsIma5A8qMsWaMBQ6xteJU/g1jIJcx
W7uotmSWCbxFNQQOHzq14K6Gx91jZgEK3+CpNWGh3RXGnNW69tiRwlN6kp+bmG3x
FA7/4NZdA+V1walnFzHp+d74x/e55aZDj3y0/OB1NovAvMoP6/b4ArscMTrt+NcF
Wan42lniQnHXxR+iFPx2BTBnxCZKw2jlA9XG7xvnE5oXnJO5VtamNvrL5EQr+3Ia
EzyWyXZznglU4yhcR8aCo8a0+TSX308PskjbrcZbacR/PfExGSkRYjL8XgfHfZQp
ZPI1NQwUUbNEJM15YMC8IMgpP74J31XyYECP5Ki0pSQ63Fg/xPBsjzlGzaisTJbc
gTT1PEdGjzCJF4pf7C/soP8H7gE/Ur6qs48gCXAUrNd/nK1XvFH5zi67QGzDyV22
2o16zK0ly9/MKZ30Hj9l+luPKamJvXDvLtHqJDGeLMaoXGMF1xtdOd0jh/Bxig5j
wphyGtQBlI4jJ51zuFKHDpfKrA3tGz29UZ1VQEsenqE1ykOzrAmdspRnroRVThyJ
X5Li28ZNMWmBmA5BgS7N6qWzm9/z0lk0a8JMqVFE2uMqxC0SawYEsn8Q0ypiDCKg
suC1+zmP+WAHOoEPLvixn5R48Ny4HtnKG6UyPQgMX36dh7P59icrFy5XeTiI2ARD
Bm6k4jPpV+vFS6FRKdtL5Rz1TtM5ORPJUFktbZAVRymNgnPALN8ESR13raUJQu29
zcBwiekjyqgKLPcf0iwqY1kWCce8KZCG/yVVDRK9kIkuY4uwklNPGmZDNH6zMSsM
/kzTKpNlsnHZFkOHc+rA5e9rUpAOq+jC3LZvWNhfbIdewDIRRl+okPtytTOF3UUp
GbOXdJobBgF8ffUc7WjFs25anik20jLtnWKwhJcPd8FpInBhUJzb4qt4F+MDwPPe
fDmJypdZN0N0YiC8n0RNVdWZzjZp28x8bD9/wJOVvisDdO10DUKEeOrdtkx3aCkG
SwB28mC7AmVOzAt03wIVuv3UbbuZ+4f7EVZXKnmWKwKUsIIx1Xysv96BLrCR8qFn
CZNs/mhAs7vvNimEo9YHA4ISZZ8hwXQzCAEHw8ZKizJt51Dou6Zf57Fzaqjs2KtB
7NTKXL2VCblv15fslegSYF/czQPGoswgBM4lHH6SMw0xnf6boon6RPvbt626lzib
69Mo7bYxXzZz0vAl6ZMCooi/5EuNahuJRZxtbXLrgKK0lQok7rXa+uM9VWUC25xK
rgvfnrOGck5V+yN6ygS96pbtpRJCcTF0xmuKSY3Xhgf1+wzrQ/OECBhNnXg8CVam
E2QkKHcZDYtzZvhEwtR302uXprxmjLMa0jQbEfWqUBdhHfgBGAEE8vbeRzC6tUhJ
Bzii5X4qh+xNM1raKJu4YTIAATXDZaaANrZrftl2hteIs3mvGZyoVab+rA4wTt+K
gNFjAPtNa9QZzACbNSR6ifUL6SkoOlzKRAR2r4H0V6etJvtsh49jzJiIOoGs9GqP
OtG2TLk+CNdGy7wmSLI1Yq1wmugRmr1rtKpe0SbIoM6/mV7yTmmr8F/+ttQDHJFq
PZJJGM6AeDeafXsqRkLVg8rIGOStehp4EBD+oo0RGfFqlCWFMm37zGM+zdFGcDcM
bXhRJ7miSykh7FEytYd0iwgI16rJf7EglIPwCSLAaGkKAtsAGDqybdanPfn/31S+
VLJ4zbSFAj68atdiD4sNnblwiZKK62BA1tQ+YAGrveJ2EVEBJp1ETDfqSPnF7o3y
EZmUBY3+RUhNsWzzevbZf7qw//prqTCUlq2vlHoBGEEcvLezkCksc3314LyG0VKf
MYc87AQzMqpaIDCw5148+1Cjcy0bo2GEzYqh9NgHfBXu8bAzQebSP5rF+qrunx9g
ZFf2nqQYUs4u4IQTIRb4TBPVhSmA1hKuffAF1o/prkmkeECn1QCFPdLQu3froH4T
5sEZeTmHOhGTEDTDmKa5wlT0nWCqRQiRlzful+w4qJoZTL8H6TA3An6Ln8e/aXh2
AnbXEzfYDNudYMSvZlG31VwX+mFwS1NB6v682n0aTrEYyvf1y21PeV6ZgccbavYd
LQM1qGaRJqWVpMu0qFe4rlHNUo80/vt21O/TwbSEhwzSgL3UaS38G0A5yawUPkaL
gY9PrIznUaUiMfIlDhfuTLRbpoPd7CENyqKj9FQzNaHF7BTNnhNM0Hsx9Rk5hw1v
N7qrg9RKFD3x1nld+Q4dn6VCLPa1iV03OmTODDnzNQV+IkU8TxMx/7kfIA7tYJtz
T6j3ZewZx4uzQEX1fXECoUvYDyotjaIu4F7HLgqbQQExIIctsN9XE6q1i7LW/qgF
YV7dzBS1HttyDKqI23s+vRnXXTu/ZBNb9VbbUGBufvMJkB0KMND4EvHIsgiuPYFL
3/dbgsDUtKyxJ7h5mFjFzRW09s/mufwdzjedctHM9gdj4HCd7BUASU+KvyLwUXHa
0rN0DhSFNL3YqPFcoS2Y1RD9RSpqMRoYAu6E9s/NUYS2bAMhvfFzNqXBwnwOSlNh
3oXMqRzS7FkjqJe1KKldl1ggd7nYvtX/x4sdapN4vepD2Nrt3Gf1Qd4KU5mLC3id
6Q0rVgI4d+2o/+LKASvtyVa2JtfR9eSHXqoJBFtir3OVIiqAAaZCAW245DeUpxuL
kg7ZrPLfsa+oaMGNUkjm43oYaB1/VLTcCUEX6/jmXS3gwEEjrFTFIdRhMqtDT0Sx
KdlkRrbg+9BnTVg4Px7hwgNARD2KxskKLm7g0c6/hRN05///PBu56e18XxFkG7U0
pW90E0E/dRYuF7W6qEGMJXALIcTsjf+LErtlO3gxaUevrzqCev8G8tWzJubrlng5
lOkmSjrEUXPYM9F82KcBuNluZOS0OuIpCauwpP9boBMz/em0plThQcnu+NhUL2Ez
3pY2cdTJvPlWvaOwv4cUemsA5RYEb1FjzRhAzncESSuuqFZG/jppqQX8FZ+zuTOE
fTeWHxP/KCiPKCsEleMOB2nPalZGWzpy4kY3frdYQ7b9EsrwLYqWPI0xIS56hwVj
JzLSCH3ig2ZBZiz5JpznQkKKNAKodpUo/TOcluSvmbBlg9egv4ZYjdP3krprdOuL
w7wdrAXAIXYDsHWZZqGTR7wJ7jR5HPp/ymd4YtypspsOzcQrSWab5hxf/psOVCqM
QA9pN+1HLzUwNDD/bY1/AlMpZHPU8hfrnlpbDDO5mZhf8Ww1eYu4RCmkZ4Hd9kHN
ETqHQw34U71wcgPufgaw2AvO/Q2XQECeTdhSrPbDww985k7OyYg8Ic4+QDHIhYnP
6S6dGFXNH6E+dB5zvNqU14EwKWiw/ARaP+t1Zz9H0HTIZMYwUOysnfGvMbBHrAXl
b5PuYxdAjbduLxlMiVA4EfL+A7CuomjbFHg5AsKpTDjh5qj8lKUehNWfcLeSMqXW
yJh4kpZ+qXkLK4lF0TOLpoJPXo9B42uuIiJ641enOjqBzSzplpcwQASygM//JaeU
nSNW3BDZTJOGfsg0qk78UNGelO891bWEufk5M/7YMcxUKb2DEntosrOr2pBjFoaz
xU+obtHVLuFrYaPoXjsyPb3eBrJuPhFucIHjMNA0qHx38zyWCkO8olES253fgthO
CiStmiEjxxFjbxLwNjxdjs/hMHghjx4vK9X3zC/gybd/YkpOcJo03VX3v4Suf+Ez
6GjhcdRYNpWPOAAsQdBk08x2s5Lpt8o+7/MWN9P1UTJbzFlSEsO/MYft/EZTaPC5
j5PY6tlkw0+cLvE/RfULx2Vau+0FBLaFcyrpBkCd8HPXoSpP+jHsithjDaHhfQxN
mJEddSHe5uTqQycUZ2N0fdY8XNa529UQy7/gdPYbIDYGRurBDdPvwmB4YJ59wnix
DpOWFgXszRCSviU/ExOG+bejhMmoVbEyRWbEXJbEHlbYQiYR2GkVf0+liD9FUdEV
r9A/XfbmOMoQApt+03nWRR6Vhvi5IEQMIj++/drf1x7lvB8+zbLYB3ZxLByrOmyN
fAYZn+WqrcNshZYAZx9iCDrUBhYnwYSPAKRZd5JSpA9ZroJmibMM7vUaR7A8x01A
+SfreFXIcN3zeTLmXG+QlMr1k/yIzWJc+ZSrjYGa/6HMSD1484axf4KO1lhYqKdF
/r66ykWF9VwEiGcliEoEk23DfbEID506BroVdN3EfaRR+p+Pr8/k4xo/fWMe9zrW
59ilD6682lRDK24SL3mlIaed0OMz1SLW4Sil5MVsD/ya8+kWi3Zd0AUFW+662IeZ
xnk9fMre0aeiMeU4CHGDAkf4skMRpmpmcqYYXb5RQNFlWhBdb2IeKHX3iD4uBWjr
c0lKzDwyhmD0HmAFa/MfOvHyDymK0PUur6k+3NlsSYdlTySLwdJ97TxkoAmZ4o6F
9SRISEFjVmH0OuvOpxqHkcUVanTKCK1pKkoXmtEwuaerzzq3i01jdE7siowaAewG
yVXR6q+FQQFleO9vAJvzUyzCoFQmU7lQk6DjHr25ez6TK5De5T5uCqkb4WUaBazF
vRtsmYQsKXlDy9N2y5gqp3O/Q6IDXUA1BiXugjHnDybCMnwZhfg5HzwNjpH93ykG
Oz8T9p9X2tcOfcl6mrKzqAWCGKDceWqLJ5mNLQ6dVJeagWNSvr3VlB1McrocQoww
+H9vjgz6D6gj4S3P6ku4Mx9jVrlNS7tuooOzzrXgUDGTVSLGFmkbi5MfhWGJx/DM
/oYeOcfaLCNlX8ca/dm0+B56D/OOOu4VTuTfC8gdDzRTUFMEDrqOD+NAr26CItie
//K17J/Qorze7ZHpzkkCxBfUxGArpv9yBQmyDOtxhA7u/6n5y99u8qfsx1n69Nuu
1Z58zfkqDyqDanMmIeJj+OFFQkJpO0Q5tztnELnB9VEDFbKLPZpcJVPIaYT3o6bM
mbh9tFl4MYGZj/X7sCWcYBJzMGNyue3YXGEcjWWPsFXyLUo+nwICmqkSvRTs5YBR
VMPEZEHsyRiQHoQtvjkmZbA2tH1HXTslgxvHB796wWmEB1nVJhMgueATrW67YbZu
l1mxU8wWwbtNioZwOLoBL/nV4PfwtDKZ9EcD9ByzPPySkYWnoTLwbqF4L4bwarNx
7w2MZzKqcI2F4CiqL5ezP0q7q4YhOmmeTOb/nbK4EOrLdImMpHMiwvY16UWchTfn
N4DY/szt2tfIt0ewc6RV7a1sooR/i732nwGGzkjK85fSHiJ+YjEryGcTLPQL5KYh
bEzvENtIfXUpH8257l3rleZjPE5+uTQHgXc+D5nsAb2r81PY5NMkWKp6/iMaUphM
J1FDCDs50XfUPseHOPOhM+Z6GgKdWM6rJtuaU3WMo9djfh/4rh9/8PniWtkkKErb
g0zBKtNCi18gAwLLLTolhSYtlFnSyP+ugpffAKct8H2cFKlokVPpnQl8PQeJkPeT
MHeYKtFyDg0A24/MOhkO3Bghrm+CgvVxLXjc8OMAMIOUr62hqRfLSZ+8dpFb4R9g
8oYoobuTyegAxpYidiyVZK63OAcQvlTNUpw1tBsRwo6PVS9H0kXrqfnhxnj1wncq
xk/vReUzzyLWG9bizm4menmmfNozKnwUpbK0QP/EV6aoYa9wxXr6y+d6518x5vsM
hG/0vIMuVTV047eKh/dJ2GV/SneujJpCW+0icM34lsWOa/GaMABDiSqRYcRpQGXZ
WQPr4uFUs/CbVpzwlHAYVd1vx49YxphPzsRFMe9CNhNVwjMU/AlfyI+H+J8+RQZa
BYvu36bLJiQnmaYzxOz0Ma4pTq3txjH23C2Rj2wmpodgOUOrRVabM91e5i0cMSST
QrIi4/kEzNHpiHJD81+jSdTlRk7pL33TA5AwgrhlxwubkY3XmqXE30cFo1HY1rKj
0tJRM4xjk9Au00f0TVUNcv+7fKDWwGsMP2uVC5opBBNBtDrjHkFUGyOcNJCDVrRn
mUztJSjsmRbAhwZ5ErHX48/JWkXHS681nb7cmcXq46Ef+DurI0pg7CchaxKjSCij
whI6cVT6aj8sc4+HthoV1fPcJf7xiyIodmYoIch5Ed16OJ7Pv2aFRwVCs0zqNm5T
KYigd9jZoZnACvIJ7Cv/EBDg4ThJGG7yz6PLTMrlR9To/FafDC5ur7PlvF8L/ynf
uBwxcCYMASnKzliSRaC/uOMKWVwDn3Fk+LtCeUsstFWCQzbflz5dp4+Nfpws8hQ7
7sq0toG++5W8TWGsuVfxZpaA+Q0hdayqqh41t8fBeqTgySRA1ReT1XRSYtH/Vhyx
8/UA3i4d5l+2Zaa3WW0MI+Plq2FXf0kEXm9eOaHlGso+X4fed5rI050ugXG0N6MG
mrZU3/WTwzqtYrVOVbaLm+sBkgHxIeJK4vjs+gRufhJ7UaPDf92npvyiNa4NXNTZ
QKzHD+MwNmP9iZoaNXQAg0SyjZek05BWx41ONmrRkUEO6nKbxFLyvWXqz+cTSa3U
lZ3kKQB7D5GBaYpb8H2amKPc6j5biN4yx7gCfhw305WSsDHCR1m5whl8uAVCETP7
SiGgp6qaUCAyrQuvAttPvBR1lghaxHyIRQedjkr9bIb9T9SeRdEMKAqo4/AzoYTd
1vymsel4+yfo5uqBxpbBC9a54Stml1JPU0UTA/jh20Fl6gD/cuAb8eDqnUyBojKa
51BfLs90ERu7K9GL7EYYCEcqVGWgH0O7fkOZ3wDShuWDZk1W9vjtr+DgaxPFV5UJ
JkOLskPu5rD3Pmo/W0jExGA7pA6/RTML5DAZBJtFxHppapbT7IYblbCNiYIQLwF7
iGw6OuaaoCqTyp7jrjRdwEIKAvixuijLPi9mBMpkij1zmYuCvP4xoF3ojNQuurXG
BNLQDz05TLT3srooY2FgiRkKk6/kWaTqGg2j3J20Nq8rd5mTgamZOEfRnM37yFK0
M6nZT0kDK3tCb80fsUWEM3IYDxYrrE2F2MT/KvxBNYYpxrEpQkxVImrx8JrTC1KX
MmGZbWR+ZD/Z7gkOug5zLiUHFSKqRq0u2DbO/b+fdkh1ZUdMvsNCsZ90XYOWBYFc
oRo0ZrizFyZzUGd2gi4ELMqp7eliNIIqKo3h7AnqyYfCSXXeh7nNQuj9PNhHzIqk
C/TlskIzxXd9ZpCm+LhkRXhIlmX8IaEEDvwyZ+xd9Jg03GCCGocC51zsPZKluNOu
rVRFatoK8a8kbfY5W40WW1yOPI/z+k2keE3Y5O8h77dmB7DO6DcmmBHim9uN0Jr2
rJXkU7Ug6D9rX+SfGchn3OA9eSSEeIpRWLpqBtUlyJPNpGZVNKJGWIDNLJiS/5Dg
1kwWzrUdSJPsTK0BjhzJ2LG3vbvZYjPud0aRxsfEwb5HB/LAD0VmHWE3Qwlwo7ZW
Q6sQzE2kNqAtbV6Gj3+C49uwieu4UCtv491LR8XX3RDquARdY+2amf863b14GSUD
CwTr7aZCLngjpIquc0P3rKE0IYPIO1SyPSwIBgunkBtXDHQ6n6UcjPzaECsOVRBo
EyN1eqlwdvFNM8/AT1yi32Y0DBguXI8f/DNjwolfn01OEAjn6GaStp7nA/Zc0pON
pbLU0NGNTey76nKyWIH0OGvdbHSU91hdcei1YjifyW9iQJWO+HGVg3T6qomaGBii
2sNH9LZn/OonZijC9POeTTas3jGPt+oGSPyrl6IWCyOZVzVf7Jzd7CZ9//HxT8do
JRli3+sU+XSvPM8TwON3EN+p5HJpywRHQPiz59wgf71ezbkrFtKilzgqfFM/XCgi
1CzqPBnEr6fwrMzNIa8h/D6VrCRxzOjiWdBDtUWwPicrwJyYHyXVxw2yhvOJ+UJt
oCctx6DUhuo8FmuqexdS9OlZ37ECgSplzUaL/Bq5qcGVQ5vcU6QsvQBVn2FIRecJ
u/hxrIv61/6kS0DIifh5/DQluZw5Q5UTruSy8tyYWKZ0uqP96g0qUPFUrsDcxrA3
xqg6yVo6NS3tg1T6GTNIV7wTak3B8eFGBmRsiV1bONiH/omvLwaGzpfwrv5bfcGz
IiQ9tD5QoqHyXzSvxngFwxexQ0QqKh68QIuTmefvZP0cJunaaIM7XFayFWN6bqNy
poYoy7M+C6DNPaU5HZUeW2s9kptexS4IeTVSodY1K8e7bPM9Ho0jFF5G50aDpjyc
YUrni3IlxcuYoEYe763juDPxRV1TrUG6hxQMbesBK78VyugXcImhXS3BkMne+9ni
yEk7MZuyEFgwWjQJn2mzOOMQ2eid9vZx2e87/0428L85WsJ6J4NEbMH8FGACl1XS
V+fmMfAEawlyLgKUMB3G5sm2fiooC6K8eLYNmnl0rDLc3XMbB3dI2cbDEFobXHJq
S3pUj/KYX2uiHx3QaUD0uAV459Ie94BXZNvaYdDtVP0ooi4UeIyq+t5LSD7+MOQr
RLSPWXEJgwU36EqXcauNYrYzNmSgS1Om92T0QZb8ijiM2YBb9bgdExZa3DFEByK2
TCSiUGk+6z0R4ozu2MeZh8/4VoqGEUTsBOIGKKTK7AYs42jtSEKeytZusxUYF3dT
iAcO5o8L8Y01LrPqV0EH5f68foEg5bCoQBCSsdbxwDwQj9vgJ2W/qM+ERNB9VLa9
mDxdipRB+9SnzMoRiDvih4X40HA0j+HsRu89FimvbSiNnepcDEyqMZyDerIOzGQt
yO8wKVm1hAQ3qFTwhH1m+qLQRww0LyFB0coceZbjukFQg/JhG1jfT5BAxZmJ5WyM
s3Bm9aLmYqrW0SdR06xubZb8SxAm3iFJEUGaaV4P4cbGY01mu1xOpxYJml3Pqgre
PtQRp2F53gcYANqvL/WgPtL7gYXNBSeoBhOuHeHu0P1LwcfUXvUThY7SMuvRkLT2
HEfmQSFzcsroh/EjAbq30Dqx4QSXE3ck8S+AkZ0dDZ/6O0BBnFIO3XB0SZLwN6IH
7DgV6j/LqvHpz7B6L4wOUZJ60Ool494HxjUB/9ELHUzIJFmZgB4+iB9uerr9PrLf
UYdXt5/APv5c+lru6I2xQn1l1CNqfMafmjKFJgCFL9KtGWT/w7gtKJ6+o6nw3u7r
XiHTpmLPPmaTpeGVCQB8PEu4SYLdr7D0HupfFzIcF6XchDhM84dUbaodPKIjncgx
cfhBKYb/joa6Cns4XsbZiI2icxdtR9zAGD1aX4Moe8u+Vn51JmBE3SuS4a9Uly5m
i36XO4ZbIry91DPdBlx8ijBHkQqj3fpnv+zFO5BMzwwA+SrLqWIU//xdtxw4Q7aK
WxV65rca09eXHCQk7x9F8iskmUn+ObyTszbbDhu1MZAJC38hu6AsYzrE3lSWNsYR
U/GtwPw2b//RnoiJxJ8eLqyHg3g18KfpO+REL3sCUA49Ymlur6qdSKFeKez2qwRy
XMGqSil2UaSUdgSvEVNsQH+uwcDod37/H7ZsVX6kMquoF+AuWS9ZpSvcUDQfI9gA
2IVN09pPihlqpIJTLFqjE3wu4UNJXETAwRxXIDPr4K8cqeLant5RDaTWxbyDpg6z
uu4hLsJydKpJvJfpWe0GyRW29D6LHe77VvwUU+EtEsQXxh/sJL7VJdMK8QxI4cse
vKaQg8dV2Q1Ic/TIsDw9cX0Zew0Cc5QY+VDvWt0CenRfL60c+6pJtmaVE9vf3u7R
06eWv7xzxAa8aohv7J8YqMKUQE2FjkaBNtbFQo0JrYbZwBNRq1xSZyB452BmPOd5
wwbU5FIgFRSwJQ1DLGQeSL+LLAWD5ips4gJK743HrYn7QTgNeo64g9PsWC5/lZnc
SLtJJNtG3Ud+o0aH+x8bYDMKDf8rDimvrKohEGGvU6HGQDhQRC6QviJqNxDUk79R
qcxzkQPCyXUL9wnNJ8hgdZ6pb38ktBuVPLldniPYlJf3v8Jv3QmTs2jBM8nrmYf7
Nh9Gf3SWNp6dNtG77c/YN0F4ANMIKY4zMQ1Z+xFdXV53oud9tzI09uG+Z9b632xd
5aqA1aB5FT9lC9eIW1mVjdOjY5RdNnNUmSxs8jWDIiqGP8oPx+96LIlpOJ5Q2DZi
EyLOWfWKNvLKzyGs5/Vvf2PsajdLzoN1SVaxdzLERrUGAeLQ4SszgGOLn6qa/rKt
eMLFFFoyKjqyJM0GrDhGwBkcv0SxrFflzv087TL0I7UGkuyG4rpZvQkuK5S0ecsx
q63xVGCIpXWyD2pc5Sz5ZypLYaEGxbx2EQ6aOt8vjgSeef2CPSiWXO7Nb6Ogs9pB
tgYlW/GRUcmf+z5P7qrIgg5pCydOQsDzFzYtDAgpZpGgORZMszu/CAcCYffu3HRB
IZmirsvwf3J3zM98lLrM/o3QAZNLHzSzlhpgi6tiIMjS2RNfSc3tooIun2MUoGhz
5olEnrk6C8OTNOU0Ii6s9rOOOtZwyys30aRDBreLeKZHn2lYccxxkI0J+VUlO7c5
ZSPtyx7v+nMkzRKllMkG1W71j9mG3y+s8Muq8cv+m4XsIdP/hsRpIJlLcDXyfnaJ
Low3iSQ4hFN8bWVozwt/I859WICRSpENn0RumKjENJO3T/0+Ymf4/L1mk6/E9TNW
NB3tcdYnJbD87Ckh4H48UIXVRG+Z/7Ji/8XxCcbrJfgELg2hJLenixZBlMfI2c86
XCu2rjyx8yWOM0dzVETOsk4P8Ys4pLDHcVdZ9yWtRWiukMPjh++RT0juhIuLo5uj
h1ZzuiPllaljBrZfDPDaCmne9+3UuyMMnU3PPTwY+r34FAUXAqR4fM1FOnNRnA3G
Xg6J9DUjMVXEQmZzoq/FrZwHFafbT7C2FD0DON+XloYlcnDJPymlytsE7aOPLuEC
eynF764pzjDg9vJpQA4m71WeYoK5hXLBZGWKw5Up49Su3LjYICRXUEFZhSOtuK22
RJkyrrsZLvdTKZ0RmTLcNj0KvyE5kkS9RAkSdOQL5uuCFCRMDFk7qVgBBygBlAvg
TFkb612+yT2nfD8hnTzNR0poHqBe748GrpIO0fDSmzhXvnfWtPuKi1HIRU+ErkZf
wQDs8ScoNZXlX/c9SNJ8XVlbNQAT93fjKwvZ0m4kTw5ZQ2Gr9Rv8xgGd8uWMl2b+
ClTssLEAViqe+qqte4mjXWkuPbQ8jSYLt7tyUcyqfnw2TS/POUeegT7n8N6/bCR0
hVXHk6vofFdXU50Cl0AqQWLPDeMWOA34LhEcT5KCz8Oh6+9ZlWG1KWLmOnuOhVtC
y5ypplaP8PUHUp/ZR0spHanmh2qRk9iwb2pSqRcnDn5nmx1Ty77MVmmHkYULiI1n
i7gOLrYwyHNpTA8zZGgb9GsGylGeBvbblUFUS6d+AIQyS28iolXas3VSpPxg8Rvd
jJ+RLn57ZIHC+ug991+JRqx9Zb9bUeX0Yf1kOeB6k65T1AOkFF8zJHOwDeybIrYH
Oj2unuw9H7fHHdlNh8eRmuMLM5s260YUCF6Ib3vHDNp3WXuJerg6shKdW/Vmw3Qj
H2JsvKIPT5syhf1GfEVP+2PUBIR84oGysVLygPwG3OXCmAwlTm9Ph7un7BG1wDeS
yEmTU2V88ebnS4ksbKGsAaFc/Uz4ZKeFhYMA5FzNb1JI66v880OuJIbj+hj5TjM4
FxclgOWU/kEGQHJUPCgHtnB/xU/0Kg6+qAlq3dMsLlDefzwkpcC9qzIoR5bOiI6S
bqWQ54uAFuRnXCHdF58ywvzY4tZCkHF79St1TRno/G74lQ2j1X7+fR2bigFv98Vz
ryro9DH5q68aSIUJ3jJChz6Ov/9d6E12tfX2SWO3CRSHu4MWNBYIvDyvrBcXJmfw
/pxaVFKwIL7xtFzEep2fLqmg38+yU30wXfWtugU2qT8zQttYuynSUzcYC9kNEkol
6qaimPaEBJcXisTpRJGDKoz+/S6KwVPV21BkfkYLMjzB1eBd9kIdQs3Ue8BrLS9c
E/RdE+lze6qCyNwpek4wWBqycfmqUZOJuhk0kWDRscA6aMKTPL8NUsH7WqA0pNNF
Mxq2cphGgqpgCUAQ99fBU236s1l+vh9kOHGezuf7E0p70QoiiQmE0VgXT6nUaDkP
lno/PmTQ8+tbq/rkJlsOYBzRi/nBXPnrOLoaW3zkn2x7RlttjqepbjfLZ5+zmHbj
+1xrRftPceRxPFxNrjiuv4XGs+XlQ/raAwuEjTQj3e0qkypvfVnRPPKCSLK7ELt5
gzVdvpG8lnS9seB8BFRSqGyFCROqnNDxLBjTE/74aUHs06cpJJpZYOlI4heVaBuv
vzdN1XRGXMV+jjHC1MvRxdrJawwL3ywz8NX3Iq2kmApK9LVUoofJ5iizcd5Jhplw
gpUUojCsfswSJ+RnAj0LmOi1KBuoC1CGKwjHE5rVIHqqZW3BRHEAZfOx8Pzk9jr1
3DZ6t2/yfQ7wx1AaxcMeq4u/qBK84YBqH4ZIcuFGngu+G/z2OYNleWng0ywmm729
0lT3JErD8ZL8XMo87x4QPwKtuB67GTidw/cZfyd5xBZ2GuBFpLQ1RnfghejFWKZU
vyWpwZ7auJiauQJAmdpOKbCSZ3m04ks59zcg9nUN22IqWfzKXF/zkoHYC3AsAUv1
YbZLDLBqXC2lXauBiEAzLZZCA7sgUJybRKZ3t3hFu00cey5DffrSbNRHQCUzb4EM
zc9ZjMha3LJiO4J0rB0yOXPPQZGqYnbpdQYV9elbRj2i6T6he/k8163GmUf344Xg
b2lowVTLE6rUucILDHZzti9b8lhyqctgcY9kUthq8GspBzML9W8//q2ZPmubLZMh
V9wkHw/n9L2Tc/nj3GZkhca2IfLYe0LGuNf/jMiseaPRVogeLf1gE6UVl7WXzd31
wcKzRO3NEpQZIzrr3II9aKT+zGqDQt/jjOyrGd8snOuzaxQTsnBFguiV1UuWEqKP
GNy11lCYMHlL3TkoUaxwXS02ZijtVzQLqmutQ6qJnCdqtfd6XKqnH8T30GyppQcC
rmhPdaMqw0E+WzJlFth+KTKVeOvuRvYHfwewAj0tS820WTXMi+aHzLCi/icBWDXM
DLGo19nIiCXoB3vi1/sFNXp9uQ9z24zI4Nerqz5uHElpzdLbF+FAiRTIae0/E3ZQ
6I2b+G0OXAYmLYcbO0ZWg0d1eFh59x3TYZyfchs+DyzQBQ4T56YXpNz1m1+i/8uN
ksp3ZMW0XNHaaFaiZINi4XTBjMwB+sPKvfdI9RjqASADmuXfwTiaGy2wTcMflZgy
amxlIdiXfFG0TMiSoHMzShFc5Rq3aByZVPEMxYspLEVs6uP87zUwiE3hQfBwZ4Hg
z6b6atLJRV14NE6OUCPf09aDngIeAw6kkBE0Opas0Vcigf/8sZrcg4YbpI+Tx5Zs
DlDQHJHHlZIdc42dHZurblM+qSbwlgcz4qAxE+5gMAyUfWGIXXLfy9rKWo+5ZsL/
bNBrtsQil6E2rVrbxlINiseTu67YJrriwAQ++Mx4WzBv4ehUYb4gmDt2+Ts+VLcP
wSIIUaS7h/+qJJzFbve1Z8zbMCFIqYu1yP5nZQIo6noL7Genwbm0GmEoUA1UniR3
FZCgm5Vo0y1jHzRbZ0RkiraQZQ1CLMKRBhI9r5nN0eo7074YwW3ETKDN1Ale3Q2z
S5GKusDBKFsSETxMixhPB4HiDFV9b8GjiJdWff7NvATmA6PxQOGT5tgsEGc3c3BU
LKIV8Sw3mgS5AkUw6wTQyBrhxfv/QfqSCVRQG9lgYqip/30lxbt865s+JmEAGgaD
dpTls4YU5PoL9EEtsV7P9THGmj9QclD2/xzl2EaNOYeD5Itqj0dyl4AF8EACrxNk
jbAgLltx3q4PANfjpZcYbT4Lm8jZmc0joqh0pTkZ6cUPoj1dHOnq9R6o8XLgoh+F
W2QeDbNdrr0VrmytIg6iJ2Me6uzQ+mMxN1AgtzFZ6ZO7VxNvt+08jYn+HkhV5oUD
tvtdl2/PdIoB4y1zTfKG6U8HL4vrAEvkilrUSlYkHuvtalCRz8JOcTaucECcK9mn
FuPUPnuYZHeBL6jOHVrh/7zHcSD/TVWKMjEu9BQ6VtrtOY91pxJZG+HhiA7795yz
QQ9eaP2T8WXuZxSUF3OuthLzUH/8jESj2mtGh063ICLnrAlAj/yJId3BGghS+B1M
xgmxFSEJKqc30KhhyX6MMy5B0jVDB1voOPdvTJiMnXKZNz4+BS7TpzgxS63xrNWu
ezPbnmR+PHKalH5+sSu0jcnOSExBUBVFPxbFgm8MT2dHUiWfGm69KYKFHYpcfY7z
eRb1sD1JYmijxNAifxlZiZFfwkw9lYSWCbQ2SoO9sL5X9JyYJGewldC4mVP8hUCZ
ezpV1IOxDhCnp9AlYtZ6EljAhM/CcjrfQ0zoxlTnKXlOB7izsFO4ltSk1DwRl1qO
Yn3i/Xz3LCiZerzRptWu8LcwQoxOh29sFw4FnBxtZLm3SCfxqjQuxF5zOGhTApVE
lLw6HJgRfkuSoxOvwa7tcatpqnGt5IKMa/HT2vLlcp5IS1HkE0jvvD5BfKY7DSwF
KOe7mMG1cY/TRgKhssufdk7R0cSpmKcYdCiIie1hd+CTjGBSd5JIOkce9pdD5SLX
B6fOApqAzIMVad+9nbzMLvDMLCV8c2Vsz+y8m7NgkfJZwlk26pi3DfI6xD+njPwM
kLS7SPEOFgswEz7AAGZLYRgKaluh0PKXXchcQ/7OgXhB8BLoF7rh3MW5lgVPcRmZ
IVAlFtP1TmDzpxSftEbCyBQmXWx+7R7A3/QK4c2uH8gk/WHz3utOxfX8cLZobW8E
IT/QrK+IBNU102I7bPlqZrZOulZiajA35HbV+GOAOayB+t3uM9XoRWyxQQ9wwNxM
bNxxk/6fXj0GDr9CXApqX+N5WMWjsC+rwfDJijx4wqSIUmLhX/lqVCIck2tAjhLH
re6Y84lzuYQBFO0Rku1yJa5tpfmKiDrFtLE7+EZl3KKJMnCedq9WpYwSVPWHqUEP
dUZVGULfDckSICHi5FR7Hsu05XsvzGZb35OEQmT/iD5WAEuD/Q9GYxvJ2lUnREz2
NoErewmNLoIXPAM+D9JepyGxcSaNxEfFxdbgVmc4tF+6uW0kw8OwHaYwfBnhYf5n
FUdZKYeZNaKORR4o4YFywSwsT1FGMtH0wKwtwTy2pUtXx3l14zX9N2/O4MpwIpTh
0SBWJkBGfZi6jKssyj6sRxFzA3SjsLICainESmVZ6XnmEvcG/o0VjJEGE0fxWxCY
nnbL+SpwGfNdTvea1LP+aOOZ7U63o4QuF9GxaESspRSK3gN1YS9W7MLtJ/q1+Ia7
VNca9JVFgBWy/LOhbc4cUL0Zqy9gVwhGtLZtX1JEATcodjP3d9RMG/yGhBRElOAf
LBY6GX8TvR+YxHYyDsmgcil3nr/bFmtMSB0J0C5+gn9NKWy/87WwSD6RwIs2u04G
5p9ouHmaPhUaDelmku0qzU9WHQ2yw4IJO0Xtn10FjtqLwDZW5K2obQhKJqBrkymY
Wae+s6nYZ3B/4TISf4NRMCqYe0Rz0PwealUxH5Rv81isKVjdo7JJTu4boAB/YrUo
GlRzNvmTyuebZoTuf5YEtGeLAdhEACyoI0AGqvNxFfs+6B8OW9BYScHi0Rxgp4wK
MEjrTB3alTUuYBvtyOo3qkmDcHuUmq+l29YtPGUHEMDMjS/FFUa6H9yoEhEAyje6
+ElfWSrV3Mb2hiymODf6T9OmWNjZSrweOQ2VqkG0R1Lhjq31dBIxgz2uJqyvAyeZ
y6lIMzupmYXKyaOWiIx4uzvTc1iK8JKJ8KNygM7PPNAuuFhUYVhSaX/DiUy2GDR1
njzWmwRAt3P5s3Bej0YEhqyfUOE0fsztM6y3ZpNnWIN/uXJ4Nf0aFy/5olKMJAeA
+DiqOt3ocMBNQsmQ/BUXXDAeteVVpHgmZ8H27Q/97OvemOI2IvTy0Yc1aTRjBCta
z9pruKlvkSdXIOQbyzgn3eYmDPzE8L5D4kHvOU3UFuWcDMY/p0atjAD/8eObKoAn
RdyrlyPGRRjFNFKUw3it2oPjDZls7ZZIBLsud/eXZrDPyyLql4RwEUj43004psJN
IqrjYsZXYjhzDuo5068jATJv6SjE3MOy8V0p23QrYyIbCpjCIbIMGexiB52OxBH+
WuMivUqdXjRvHBmiqhFFbrIF8hyGCK4NflW4veZ0tJQDHnoBnH1AZH+cuoQUMLRI
WypM4y3+1YsatQfLKQsWSTSyZ3Hq6kQ6oO6rJKHcHQuHqTkxxgPwk/zrWuiqyuI2
F1r0m3YyAFhFIRPnWAQu9xRhNl/B9pmhgmllVj6E/NZzZ6PGiVYtW7Lu22pJ/1dH
OGJ1JoKltmacerbm8Jb4Yr4oFUmB+OCiP/BC1Kua6t9BkccrEqNsBWzTCRw1Eup6
zjPTB7s/Qs9gfxPxXaISbHX0xUMBcGs6N+xMRGoM7znSZQ0beC/VVtJmwtd0ORkG
05iMTAqOs9LYE//NH88gd5TjajjrgErk5TVNBh2MTuzlc7w8oumGE5eJR29okAN3
swpccSEV+F+KfsFtQ9x6DtTo66I//lHA9xRwcjbOOpjHantmk48B1VhuZJTZsUer
u7Q6lTkJCmxgOE7ZWm254EgTz71RdB+EfbCzKQjq4Qew5OpbL44iSFpHwOy6uxKT
sWbxYJkqZZVv6ogeuePcp5SbJEE5sP9EdSo/Cz9XdKItNJ6CHQjsZKBCE/GBNiE/
b8KAQ+pkUGiVaASMdoz4rqZrSRKyUEEPIKWe+OPIb1pRPDeNMsIKZhdJdLlbwBSt
c8HZlOXkQkJmJkIK2vcdGMTd0/jCkBOBAOTDqsXxcnue9jj2lQXAmBrMmkjIb37J
XIzysgWAqYgrYRYpDu4kzbO0J9Txa6gxqqZgyJQc7PPAmesGlGeMMn096dN9BBFs
GWUGGxdyzypJTsehO2ElftsxdfllKozDerD0GwVCj+S2dhIZ7dpSCIA05taEFplQ
DvR4JiVCuY5VsVli76VPTkMRdfCJa4OOyEfnEYxM3gjjIMeAIDuqVCZR6Ss6I0Pj
qurWFCxNGiYyRdOCkW0axAaqcZ3Fd2xg3OFnPwyeGdFRrvqW8AG5Xq85r7gIFFMg
m3K2b1I4vGm9Z+4mZ4F0HE6VfEhZGfxfiPL/0nyzu6YCm5ohAbcT1UrGmR9qcZlI
EuQMBfQktVqfjIeY25Fip8ld3YSU4lb1Bi3Bq5J8dI93Q7PsHDltvw3FFUeJg52f
ymdpVtdHU67Lv9CM2PuikIqa9eUL0WQlBrfZ26yJhIMdZac0aNKpYiD/rIM1sziG
jqLY+aBxThQX2naf57uamBNqEUIlZWfX7EEFpnKR5UAovyMobtCwCriwkFXynqsO
2ZVpmyKD2Kz2JkSwLg6CuCm9XGMvJ2sU2RSfcOXAnDf/ZWJzCp07vgLTXVRKIvAg
NEcJNExeKIrySqg2Y+ymqxoT+EjzO4x0qDzhC1lVgHoWGnEDYlDoDhL8O2wVN6Jv
k6K2n00PCMgSLIH6HjTxtZWtH2r2+pgphkhlXAqmQrfrg5VDVo294kjBYe4Bm4Xs
ez1XOsXMKRUcOaV/YbnSiAWXOuyBSPWnxg0jxrC7zbW0o+KDWYgH9A0X4K6tjxU3
xLfiEavIy2YoePZ3Hg9QKzWHMYtLtyQIVs2PZwWjdLSwfJ1pd81pIe5bWf2FilK8
+1KrScWMAIEMUpobS+u6gpPSrkSFL7sMunCid9SEK6UFaT9+XOmphq5vjYPfSsgX
2RmYPbV6wnZz02gjOpgV7xKukMInV6xJVJwYr4h27jhRPtKNeRJrRb1MJzgqM53E
AqHH7kGeIkhSs7DfHB6p4wzARdTxFSdWcCb6DNu16v42/etTqlwhtswQasQD2YzI
RJvOiJhwOd51GTZZ7Y/22Doswa70ZX3UNs8fQaMCtT+54n9ySquAMvWvnWBLpmiX
WrikwP8Tv8aTPTAIyiVQpWqH0BVy82DU1GC2mBO/KhD2bYF4avgHd/0WmmyYAC1l
nXBNbVId8gzkIweEFNtbS/tbQwYDS7HHx2+rY6chdphM55PJbmWDzPQn/DplWxyu
APIeH3J2JkPXQK1tlROs4JwHW0go5BAGBWUtMRZxbah2wzAGvaKL0gXrgPW2QcLc
/7gOsezx73uVfLcePGCqFCmbFdOKHKvqYeSON3C6Oq95aAw+eoF0fEeQROoGq2aY
Z1QPbb6Rk2xWNjaAguhnkk0Cq8az/mFgRjmYCaDsSZH1bJh3vc8odBK6wyl3/21W
hz5zjsp9Kqj0Bs9+wKSXo+IhOBxX5UzbmjmDPciFI4+FQWtmX5/36JUql+eUxO7i
j7uZN+381NlBsQ9yZZ3xCgj7kWgX8jxW+YiFidEyh9MBi/h4JMF1wgp+Mqa7o9ht
t9VDKOhUBsm2UDJEPk5tgUg3fmPL3HxIvkH1mkgV+lmtDA50VRQVJ2+j9pe2uB8B
LOeFmDymLbz66InYviczmU+qILrCihb0c+XNZoAkQt9QdbeVImmSJ0GAlw2Ui1dr
Nf5DpnwI3/FpDKIM1WQkkWeI9ZWY6xJN4qotk6N3M0GY4XJ9Q6Mi6MQxGwxVjrOs
X+oXEwqkJdJtqLIDvCd7Aqlx4DnLg5kJTfyo0z1a2/kpedgw+gv4PGhjsUUSqUju
lKQAj9v5c/dvR4/P2XmW+XZ6EmEjHfERtD18S6dPjOOtJ7dG8GZRP0AlBOoRpN98
/NuOBi6bPqx7wfOcbYHhsmqXQ3gtwXX08+W+Tqv54vvfjRLf6EiSQDwiCKiNvpWV
mCWo3mFXNPwGEvGQOrFbbB1heMgT5+cU6NafnET5+mhUuJYv5gTo3HSfbX78X7d+
/kpsMVsH+ZSjsHvgTVr6Na9DC1cEJmjao2hTe68CilrnsX4XcdlfePCfdKWvWX4R
Pois51hY1L4BL/W/xUXZZK4HvpMavGprRMJtreHYXi1ox8ICMY7BuAtBQLlnD7wT
5uP2GRKx+M1sCIcaDcpzqRDillJQE57AwTvNUIqgcpEr3gO5b+QPaH7zO0aHm580
RUToqxQ9lTqyw7ahWa052n3GLS8sLMv+hindtF0mlkNPpTa5jqh8DvnZX0ZYzoYt
YuM1ytGv079uQ9JqIP6k0ahmbAm1E9CDA/nbSh08dT4s96S5gxGb4NbSKPAO4+lO
BCMJUicWOduxa+bYbIfiB0XoE0noKnkMP2+CO0nhV2xxad1C9wzJshEnZLyOnZYX
BtZpbZYnTPL7y6M8ZvFCZumPiE/wXX90L1PjqrHp/E7YOFL1jUCHTYHOK9xlxyYZ
WqRo9RLBDPKrUrG21G93e25P1jVdva1rhP5CrwdxA8Lr1E1LpmGAKGLmH89YVWKb
lXKTMvZZZIWI/ohz76cRyP8fml/nDfVi+RDPGL7wbXViRBj1wisvmmIHPlrVCPoT
KuIwE20XJEZ9TaQZwPsUomC7BF2UCCZOiA5KFIKmBwSzQGj6xBmND//rgls4XqfL
Cn+Zv6Cf2eR9HOceQxzIH6JqiFFeVS+heRBGWVJuHeX5MVl/Q3lyVBVn731tUzrR
GoYZEnYpK0sjHlHJXOIF/5UipuSbajqmhTzaKQBZQOXFWDEE7ojRJUHIUNUXEoJp
IICxcQxLFysBM4uDkt8azyCI+Oi2seDExPdL+U5B2dsYEJj+KglCQXwd7GhK+gb9
94jBWFRaagfYxpR654JeDyPuvWfzs0BMxk2NWix5cc5MrBCy4jrA6jhsuI2l9rt0
ywB08Roz+Dza5dflFNVUWPd0mxMzF86lOGsEfcOPD+3/qOAFYC8L2v+l4OLEfrTT
CLfFPjQTjRHI17QyPMKMsD3GpSCcAUQexExZUqvMRcWJjQuw93aKrkZoN71WA0oj
RsKn0K+TkUFoQhhXUT4ZDunjfH9AdM3+poW7wD5g1QUvpzRN2qfRkkAhnLl+yese
TlvpS8oXewzuIr+Jl2kEkSZw9fz1SaFIVc/BX5doCWQQ+z5MEkIOMvrqcOeP2QHT
tNTmT1rUdNhfrXbGRRmATmEyowBd+SrP+laU2G0gsWJ3VufrwPqX9wruhnFMzcVR
tHz6EnplkDhPI4gRhAr8oKQbfVkwibPbL4WmAkpxoaNF43qYxsoQG0NAvlIswaMn
UnZ+WZNlE178b4cf+ofMSxnzY2d6E9JBb+VKmGSENuFutoq+iUfhxwgqu4U+0vlJ
jTbOm4Pbf7Uz3nQxR1cACZPjVRc7+6aTkvy3RavM4VcI8J1a8SBdPlLexHAIa9k+
M2rDgEnnB7y39CWaomzt/QkSjJWnCo059N/pLl3UmIwxYf0FQOTYIXYUp5H8BElo
/ovMujaULuIc88A7pKhJawCm+0GI+EhyZ1i3gRc1yr1QjBIkK5ntXgf/qy8ff44D
Iw3M8ccTBh3FjS2JherhWs1hi5QHAFebMykkokwkGxUMTdP2U5VFKBVw6k9nP6Bn
vySK2B2OR2d34PvkcSpXuNy3c2adnj9vlVOe4vlLEj2RFz2QwdoAf7E7BtQ/c7b/
lN0D1MWE5rpw8kMUDVUBI0dz08tp5XNpkbNIQAWzTWzzBBrggnSBoquVW00KM5bZ
3uvdcHfiQsjUzdn8cl/p97SSIJxEK2EeaY5ebymxZeeN1dRc138UJDeHqnYwMR1J
d+3IwqABdBx8zOP4h0D4adBc9/ya8nWGObbD2mLwU58X2QpiGSVqJYQZ/gB1ljju
9CiIMoed1IcaAHzdtzSLuqsjq1xHGbqTQxlK8Cfn1ZC31y+x7PG+CkSrtITAmMoU
S/O6g/M0epvCqND440sFBYmb8JYQI5vk8HlSU3a/Pzp/yDs+0BqxWQZWkfOiAFlv
3woL/J5N0R79GgpfyO5AZz5lPyVKGHziUAnChnMf4pkgiIN9s8pCB9aHC1wMfeF/
y2vXPujMJ1f4ELHPlzlqyxbbFImGXRO3d1kWYHOeNcobpYMH4PMz3EkEKGxKqAzW
pwJV50z3zzH7TOMXqSt3VF5T1k11e/5gNd8Hi2eYETeEJMmII+k9IjuDyEtr41TI
7YZEUJkhkeZBB9nk8g5kjoVciKGAPHNjX6f3OD8zGmzmynW6P+ncRCwnNk9ZKKxL
CqzLMtalmDzyxTBwAGQfAt0hHOunyOLlB6fDnOr56N/L5z4EelxGF/gZRUIQXp6i
JCOBsFxmCH13vNVBKbOsYUUfz/UXUrXc/CQfB6TrOTF3D7VnQltOx5B3QL4hJVLi
aQN9qmHS55sPmoHKF6wyaZzrfJ3T08nGKWtQ/iiK+H3jpfyABo7eJ8aHzyXZY3q7
Sr3LC4VEfj2IdtI6ipNBATkaY3Pdes6o8YNjVJMDQqU7Cq7WtktS6jG+2M4i+5cZ
oCPU3AlqyNyHMpB/SBlJuFe3he2J6qSyhdUGjTbX7iYd3WfbUHMUSyehB1x0J+M1
GtY9iVxyUaHMhP8e7TK0wN42iMC7v8wPaNLgFqM67I+UKS1yV60exjcPk62uFCeQ
PhnFJbdFhK27WM7Yxgka4UI/RmE29gnsR30B/1yzAkYKxsnYvMUJJkrt8/o7Fch7
8zAeutvQmz9MwIO3lc/Rd/ULzBkf+uDWecfB5lULdEqU2HkFiAPD8kEmJkyb0xjv
i8XzOuAFTbDthCNCcKHIymtYAqGzTff40z3aQdya3eAXuvs3PgGORI705KI63jVR
TGPOoKrnTWRwStxJCfUBq5aH9/vA+iTmBw6yWiCoEN6TxKa6ykUOkDn3HcG7VWcY
TfQm3mw9MB42AWQOR0cIYaYoevasEXtaNkb2xalHVqWX2keKYKF18Rtn6y72WH29
vVaEtx/ssK0Phan9LtUL/cUF3Lxb0CiwJXmP7iG1g+6qwtWN2LioyO8urTpt8HUQ
Cghmu0Zk4NtiqxWenVHYhmFYA28GfOmI0h5uwFbRS2aqJSMbUJACAkTFK3ilA0Mk
yP249yiso+rdl1EQ8C1cZI03YU6llxVt2iDm5i7rkcyPTFLY/evdwRlNw9lljAKA
ETm9nEA+DcfVQOdMIIALamebbOI86B+w50y0gj2JLp9/7Oc59MB/KoxTHk4phPyy
pmEt5zcPruVdgPBR9yiD+KjXjF2GuGY2u3FqmYQwj1OyJMsQbWCQo0vKMOGmYZtD
TNbKDnj4KyY/yZpbaACUWo27mrxpGGy2qOD3gZY4F/0kModK7cDVE38QCl9hlOFM
dKFOUjIjZt7t1EgzGcsKtdn/dKaJlZT02dfQlPz5YliYG3dN1RAjMe78tQOIRGPz
UNeppVT+DgZELlNyx68GBv05sJSbtZyguf7MWNQwteaeka8sEH/aBj+m1TNEfqWX
C/lIiBZjF2/H5hipOE+RBqSSRB6tHKXGBBhdY7GRQAfCfG5RcyP75U2tMkIC6ux4
63a7/JsQ+A09+SsxJbfweemj/5zGPemSfmwvIHeQtzPynH/w7kN08IKZtGDD2WlY
6rgzioLckLEWY18TA94mdmMuB+jN47TUUao3zh06os5YPwEpK2ixVcpatOuaNfuA
hrzkcgubndUCTHpFDRm3ZOi5hT3x1pfFDeeyusloxE9Tx6nu9XZOMx935554Tta1
3+oiS6G+WRQD2SI5wYnh41+ih2Pn/Qa+evBJ/OgmAVShkSKV63BGnXTIr+eIjE2f
phU6TwQqixnXNWJXagYtHq5pTAHSU0DbQpyrFMA77Vic6V4AZizCve+xiM8mlPjE
lJUs+RzB6uw8Jf7hPqb6ifmxKkihb4FLJEHJW+lyz7RkEEhikmQ6QZWV3Ao+leGg
JqhIgRR5lyvVLT9NVC9gvO0BtJr/XEgFIgG3M/LWUM8EXTZqZjMDmtQ/krEfmUBX
PMLgoNBDhhUDtG87O4xoouOT9+JmDPYbagsJOhmMxXeqY+sIuF9iDuHdZAlxODEE
0dGPPC++NHrhr7S/bA2ORLpitSKvOuGkptd+58p722v/QajlWhU+X8aoprXO4bAe
/afhMFDi+nFUKKLk4bnx73nSHCAB/Tv14FDrmwRQIp3UOETLY/GrWGSUtjxOyg7d
O2J/M5TeUilwgUEIKRmL7aN5D++gGnfDnl7ReRBhn0bbXMKMBEOX0biJpphrV6ev
JouWja/ElWgIU+atr/eoBFlBcnDlWC+1WmZOg8P8wFpakrfYSFrG+SfOXhkumXbf
qPad/WtqnJJIn1f7ktx0Y+eN6yh9v/db5sSGTSPjyspkKKDKUW8Y1ydKQjpW6Av6
utulz1Rbapk4OAJh5/s6xrRhXfu/QVty9fEX6PubTr8h6tLLAwXaHMJctcyupofD
TvrgET1o9W8TCKz8DZY79c9YIIYSTtPCk86ZVyH2kZ2Lw/EMsmL0NPc5OgbSVwRv
TJUC4AzaJLeAPWH7XMWSDsJ2oVK7cK18YQIiV62cqpDxeecuPfq4k7GBnRdfpG5V
dM50ODjNB5ZWEqZ4bUFsn2dlJUyViRiYZ05sT8kcVz9q3B8i95pyqDC8w4OwVKik
IfLGFvZosk0b0D59vneE0+bD5jUtipXJjnsylMcrWtJk1xb3pgRAwGSFOOQQJcgH
cxVpZmLgmY42Qd6KgUfpqYitOwqQlp6O+k7SzGt48ja7TzE4PoluFzXeJlB5XVUD
8Y7/qHRplZJqhlNrB2qWrPV8SWGFff9GI9yyS8DPadJoDeTGCjoOdVzOL63BP4rN
ZjOcOOTjfAZ9bGb9iSX0+B5rpoUt4tK7P3+5NTaGVphHxLBuNLWg9S/ALd88n+Cc
IqcFM/fDI1he7L8jMibF9gkgWa1DXng9AHmZX+hlvZm9gjAhZpxWEbzV8DG7SCH0
S+7J6HSqTzc2k87Yh6ehf3YtXRj/fGlyoQ7MKo8ghZSXyOKtFxsqg719dUAcSs0p
96dpeYXsWJClQncv/kottksXv8RQEBtkWz6z5vWZjIyXRun4Msu7kUx/yKlUB9P5
yZIBUIdgzNMTiUZ9NjrdWUaSGsmewJIioRjOfJ2yf9GeLTPfPFHpICAVDDXKSB3I
VoInb20QnD2RZg+s6ud33Vdl/RwbcoT76VXFewfDmnqqfXDfU5SflEYnivAK5NJj
WYID0t/gPBQfKhv7MgydIvJVOcJfq4BavzlC0G4Rxg3VuseGYiq7nYSXq9UHOHlz
3BT+AfFflg9e693OJuhPyjcioezX1qIf0qOWNpkFc7S9DuPBLebtfisL8q+vDfZf
AZE4KUQPS+FERNLbskKQv6HzTWF/Q0TN4g46jmq1Mus3yRx+dWB1dn+rdHSESh0m
XpfkIZ1ecx8KY3875dWVtoguxS3U8yxx3QKKxuThBVdZC7QOaMTqC8U/fyddKwhP
vcdf0m2GcHCeBd8bGQnkKY6hgQwP4SSLMnzn/mrr5wUdFmGILhFvC8oN9fXB4OVZ
Nm9xytAyd69W9i2DexwDt4+ktfmciT1gb5LBogHdb5h0vt1YR1yNrWjfKj8oECqL
a2/Utpip+wdK3RKw9q5kaGEbo+kMnLDfpgQtX973bjRVsCzoU7reu8kRcZnQNJlP
NcLVYApABE+tQoUHQIU86VeagA555CBROvliGro8Gl2GXtAZyf3KS4+ye2Km/LeS
2dW8OSzzlY7TDKJEGCi2U0sBVrjPdM5OVQU9PRW1AnGf/jWe7iogNQGFQMcWhl08
73thvwFB6diZtG8+kK3k3GsAcq7Xs/Ia2R1owu2cSiaNMpV1osbRGHRkRLecxnew
pXDDz83lyGG/jBSKHEgbzQU66rnws5+Bzv0Akn4p2nLmo/7WdHiQlPw0ACjf+Fc4
3I24IqUXpV8A7pUr16Nh5QTYlneU1sY+3MzOPqyhMWROOUJL0MSNpso0W6d6TlgF
hyuqrumWMsDLk95LpGYyJrosXgCEM7d3y6iVD08k398h8s1OevQYeRsID/y0pwIR
anrgCSHnCZqxWXoIJ/nlza2CpjhIuq7E44FAzqd3DGv60YF1kADkbWRW952rxnlQ
venT6ltAoCI/tU7t1rJv89VXgvTAWU4v748vghnBOUny8DtQo7ycxlaFfUF1UKGo
5wQwGd3kxld8NmAc7tq0pKrw4xOlEjQEow9J2k84SfYpZNFHZU6Psj1h0GSEl39q
2xSInnuP5Xbp47Q+enoQZJkYiNDTAgAzP2stCDGFS95DOgAWA1hdPU/pDbwMZAhq
28cmNEiF9Y4Zzactz/niiuL4UYsNjC54vOCSh4aXwL+IVxgWyJsvbCBKFXC5Ke5f
ZF823iZ+ZqQSXCAeKLWPSbIx9hh+WESxbKtuw0nBD0txhlw8R6AopAZfmG0MiwTP
a5EV6OTQCqEjX+tAu/MfwKwgQcJ0ura/QSY1X4rMeU/GV/Un7ksk2HhAhGwscqC9
NX3EAR53ldkRKd76x9TZzp2FMOye2cF1jxqDkNDTwgemBVeMLY3QPW1AzugjA0sG
gZa5K5Z4aoA8nw15FegoC4n+BpECgrL6CsPPuFb68MbM3TflGq/bX+at/7YaWzhd
RdH3VIOGM+aR3oUwXKM3q2RrQuBQD169o/i0AqkRToTpY+TNvs1ZOjoufZQRn/gk
agJcmbe6R86puRu/rnks9ejLKVPKmkLSWkaTSlPsaKEVYFns6O2G2/ZUDsTYLLh9
0D5BTsvOJYMYSsUtIWGD0XUdCrfBstMrwev3aXgy5pue7WmxK2pLgS93FAltGd9e
+IozbFn1cDyRjcLAov3QOOo8GUkJPxom43vT+jD7VQFuo3JxNKMERMGJl5EhXkIU
bwKt38i+7sH0ogbPcUx2FB4B0UZicbLjsC1tEpcx1cy2psZDc4jlvImTDJTd/BVc
gH6zpdpInJKpn15j8IVzbPjxWuuCKjn7zLUsiY3afRVVBnJNBFtw7jabFF0YLyBu
dN1v01daKXi5Z7jbxdWuTOD66S7IUNobEAsLsyF+aFO93yPF3lziHiKeFdiZtAj8
Vxxpyv9TmCz9Ik0sLnZdLwG08g6A+CK5ueGY/vYjLqsK8Hb3cKAdHeC/1wqu21Xs
NJNr0LQ0OY3ZaK2GSqHnL3C2PYiV7zsHVcgEc5e2/2ICpIc5sbaYc0eNyyjc34Bt
Cgh2EHtohKRU51NMFiW6QPbRr5nMfnPk0LkqA9R1rVhJ1y3y7glCmern5YPJt0bQ
liMX0/zpdgQNnuFXOpSdpKX/ls1Z8hdRLq2Z3AGHZC/OK+55eFuFm0Bh4RI541+n
B+D4JQQp8FWGtYq4ZOpqZ0z8TnzafUXMOrkCJ2QM0TukhOhrxXXaQ5YyRUCbt6Dt
4TwQcG8xhKwcRx+t5I7bt0qmr9kDlNswGVUQyeexItVFUN8/v/xvQEF5tJCKqlEU
cmeo7Gjy+UnVJzA8/sqf30yAlvYD6pyQnv74nlqcU4f+M+yqunOFnQTa7wCmplF/
G6n/ZbNRQJCqzVw3Tgn9Ci27GIM9sdlYXfsbpEwFUOKymRGDGQ7vobqa1NpD2dj+
gWVEqb4CapNWIBoavEE/CT5X1NIX8LE9RRtODpO4maPTqRBuYnOilHu5XFnNi9YK
CPaAwTmPgoHOfooz/wBp8oqTL1Osnt173UQy1geRnJj4in/d6MMY+5buVNOfoXNf
B85jBxjSUp2hw/YFq6JYvWuKn15WTe3RiZDExkxoqzv6nI0lpIKyqKmZtdRbKmoM
oIwfXnOVOzl7WNt3fY7H1zvniUZHqAw7KGDpWWIIjtWjruF6mGDTLFDBSbg8kYKS
dKY2i6z7zCQiJDM6/IMiGvBWuHzRLUYOTDjnTEE1xHSuBi20+moG+P9+8qtEEuGh
uHZfW4MAec1HgoK1GImx3QrfTs8IbHB9COPIpKwYqMOs2uKvRjqNxejKCEDb06f1
8IHPQU85RGQyBnfo4ojvfbFwODGfvy8OKfFIur/6YOWKj6OaQWxqYRltGdWDc/AV
XkFaqvrI14tSoitGjwH7ZGxygTxV0d+5FWcv4xplR9TxohUpS2zxghaGDkibcsgD
wWpSt+DU9TgsGaoMUUtgiCIFL7tc73hicTeHK6dITCWZiEFxzv3IAUZILhRuwkaV
g8stbk0D4aHG/9QbxWvFuyP8yb5/pWhrsRKHUZKQqpw9T3e9yMBphBLxZuo3akcu
snUbZBthuMYu8vViaVRGWoFHvcI5z/hL2uSFm357virIp7T0Ktpj+e1XLZ/KzF9g
KbEZyt2FZmOkioRdfQn0fr8j9Ufhbi/PpdeV4hMkfJfL/KclW57sRlw18UWyXRxN
3oXMcXeu69J47LsLeQ+Bkx68HBydhHxC8rpm63W/zRlZq3AC7mXbbzqD61Nk7P1z
SHvwjtQ0qmaE/lQFUlauGFAhJHWnEuqklcu8XtaIH+865yBicrTz2Te2n96fd0Z3
xU6qixh7p+cEvYURjs1Mcyk5y3fwLOXVhnIBHQF48srsfEvcGcTeiWdWM7QL8doz
ZRMTLCleIqJe8M1cmLos/sLgl6Ss/+TnMGLCLXDfuJQk59Am9ehftHHEttf7CTGN
C1H2V28ZkY3fOiHWGNWcYpzjgZ34MmW5Z/3r6T3S7OTsSHY+YD2TVdR4Kfx5PAYa
8+L8DHFVNSjURNL39d7Uss6fwAAkUQGa6IAQA2el0Se3FUfwV8LvmdLw/yS56T8j
PT4mXcCEGJJUWhJ2SBYKrow9M0U2MjuDD7ADxY1kD/3qppWpzNPBe1PBMYswC8pX
v1mCkI/YebI4FyQMLhx1t+GlWxN/tr2zJ7v5g6PfdOCWcDpBzubS82huFE26x15U
eGUZRfw/+x+TXVcS9GOYQDXlLvlscd9HEFkxczDfheJ8S1lbcG+t19eNGG8Rmi6M
kQgBMcH2fk5s9QdJN0dHVmmv00EPetEc2xwUgR+1o2uCixTeRkMdwjdswsuGin0W
SgPS0IiJ9vfXCNeuhxSsYPI0d0RT2dNRr6Q4L0eMcIrjSzfVqboXPFt2YNu/qPpl
GtTOUHruP/wUCBCG0W24fBROzgNIsVRVknZFXruSitVClg0Tm2kDbQ+vYC1AUTdc
Q8gXEGi0kCRpGFgmkirNDvo/xXADzxev8Zvmnxv0y1ODXrWdU38NzTISyrQKaWWF
5YsWEO64+hvr8B1z4N2o9sZnZFiaCp61ujuW4Nr4mObhmRP9DkPD2iPnJ5BjBZcR
gQPR00of+jNBhqUPCoFAXADfl8tfLQ+9nlhADVCD1uA5ViLOLM+m33vjAPNo5jKQ
/rf2Db1d1iIzOkesivjM/KHglkK9xzA9d0dc7/x2zfwLBF1c7yAh+QLqethGS7FF
fnavQUV/q74WqaGXyO/lXkYyqTjptL64AXGoKFjZx0ojFIqMTwlAVIitkf6Su46O
JrNFbLC6rNPfeidVtzUEwD1Z7bxJ6ahUJ2LkL1rzHc0KsLEa9vTgnBqW8yeTa4qr
bZUBLTq8KS2S3otXX2nfxHhci/9FrfCsn/F6CKDadqBQoaYGO9p6JqbnxBTOdi3E
R9hhbOUaw8qGCHvHSCKTpvNmImzL8WnFPSQNEMXyrdp/I45+QYrEnUGRs0+VSR+F
Ad48xnUy+/IqDhkLQI8XnigNpC4dBsRhm5egJHfxltDvLrqD/OLfmj/QQQ+hsNTR
Fh+/lnG77ZiLocgw/OeAwIxZda4YSZ2UuIrZP48RwOCp33MB1gQsdjVjhnR24160
/apdwgM37vBCpsHb2Gbxc/JNKDzfQd9yegQkIJ10wnEprb91kvbIycw0ibrJqCAP
OSHRJsQ+nnO8EaI8tLjCF6P8/X22xX/pKvbImF0Isa/ZP+jiU/NuPr2raa0O+RSk
8V64CJvPiNukWOl2JGM0VAcGK+Xn192SeFMSplINd5GhpBRr4ECRLXb3D5WtnDG3
+mqoxwSHSk9wcg9HfTYWasg11Em3wNCw5AH+dhyW0zVccxJSlin3sLriK7tmOSFC
82oDb4SSfEdGVhq3Eyc/jI9qwguHyLSnHwdE4elTk9RtouAyc+CmJOnIKKDkDQN1
7JmWX7ssCvkgvccKwnfZTkDjPG3wok21VSKkwp83/CE3wdTut7QtxEr/B5xz0vhq
x1aubBY9ui1vL7g4nObxjV/p0VqqCazvzvjyXAsBh3IHK00Fiyf+5TElHOpvWQTW
Paq9nGOx1UJwAQPjybkxiaCg/+OWKg2BJCzMhIsq8kWR7n85kQQZHfooNBrINRj8
oN3ahyDpPrq154Tfcp2U9dux7VycG2CCpuGp3UWEVcCZnUWSlI6nos7yttnnqSjB
cG+YaiR4Hvutgb9KIuVHiGh0ozZCSAiJ6dNG3vBR+5o4MWCSUqyWXRpvP/nbeOPp
HFoWedOKorAwyGM1enDtCJIosrDyxMoQ2PQKxhlIa/ogPNJ6BEYsyO8UqDyUYYxt
CfI48K8+cbobRjza3oULJgShV4eWPJMXE8KfhkOI7UrA/B90Yt7+YPZoXVt3hsY2
OoWV7dKlcWzZ0Xk3GiLSwDAN7lR7ZEQlvOPDqnolcwKZNTCGI+C2KrDya4cB9/2v
LVT65EuUqfDemIg+Zww8modfDX1BX4S1LdrsDmwhVI7iNQxROGZSRJxkuf/G2t1l
DmJzi2PeDia7BUKt2L1lwseyf0twcyAFAh6GgUSiWbwEJiJoS+Uq7dcKYp0+nyW8
OGs6BP3/HVy61qa6V3HyuJydQhGyeFwiVthwVjUMgb4yjztBu0G2dZCeiBjFgqLw
lEvnABtnbs54bxB46sPr/8X+bIlRb4CU6To6eonG03xXY3/0mVqxrGYjILkpPl9i
zdvb7lHcbxnQxEREnOjVw0L7x2FM4CzdaOQLioWbWTjZKCLyENW297AtOlPer8D+
driLQG2ZoXtUSAeCTYsV4f5BCQbBRqlC4ODVV54H8noyz5eRFyynL5Po3i3s17yG
kFkdkHnV/0JVAFH+9NAbPs9JTncywHRyJ6HY44K6mqsgx0OVCdNJJ1Mv+3ZhfyPa
6ScaJJAIoRE/xWPVw8elrB3gyzOPyYLvuRSEH/Z526mTTkbzVqnsZTnfRYgtOq2J
tS3zC+UBq5DK/ntQujbVXmQhYRxWwTVo7ZSN1OxWJ3H1KWWpVi9TC1PTKlZR+sx1
eJfXQ5qEwnK3wngAo1SNhyeYSdzl1Eqa2uuthnsPSrNu6oY0jwwXQdDtfYYwfKO7
7JQYbI0r0Vr5/Y+vkLNuvuPrwpfZniFfamiqBe0FqzWiQg9WUV9W5DWAwyL4S0aH
8ioFLZKlZ8vCq7RlANPieBVpE+0wvSEgshwJKYTZyhraetP9uzswTeVzuOYLxSUZ
x9lweYeF0u/opr3EFayIycG8J5c7Kd5rQ3mfZUecilZ1GPMmfFbaLnX4JyqrYeoj
y94syCx/ccqcQ98Bh4pzzdWLkYVuTL57AYki8mnnZW4H0Z5vIHY4ewfSNyfJBFYn
Sg+/ZyYeb9/SBvM0uDWE/CzkVgPBVVqoLimILGgc61AF0ANxVmZagZ8Eoq5j0FvB
vKOZkJWe6diK9qT4u4+e3uVQLbzbz6E/LDy9Q93zb6xMNhJDhN//Y8fDL37keRFV
OfTpAiVHJMfjYJmUxaRV7uD3xxSkUZJO7Fwfr1sJ4+qmyISHoqlDAeTQLKuM0Hdb
XXgqyLPmZDTAAMbvjZb/xzpPzLgMd+9MMFVVFZ94OPm9J8DMtlLH4QusDxKZme2O
ok1QqlwDFgnF3DKdoxG8rVoEIa04TOj4RIPZGxLjfn24ylmgkl3IpKhpC7p9S/0K
AJqTfhGZa7Nz62y3I+0Q4koh20GRaVSwNTKB95iPk9zijvUgfTDFtumfww7GNeWs
0ekbM8NygbwmrDgg4nVlY1J1ppOwQZlPn9OkmYEtkSxUWisn/NmkN27+pUbcw2ar
3BzNxyJuBYOjtBvDA7cTS44G58095XF14aj/TBTbZ5uEeCJigim5mc80WuXSCjyP
A7LH+cu8w3FJjtVSYqh4zLDXl9jmso5kt1UhsfktczOewqd9cnrwr5VO7HjLEcSH
y2mr4HNzDI0mKrVaT7tgSfWoUXl8kWScQZYhJCXe5sLjBiuxptPeBaVdcJsD2Jva
A4+uJy1CmE5H8V7oXGC9h0XFRsMzI0LOjQQb7oBPzXsMrZ13f8Mp+JmTGB0Y6Ctb
dgsh1CUMlXrFDIeulCDCwOq1Mc5MQJwuWjxY7xHbszzHegt9P/JFH2JKEm245l0p
w3oqlHd7PjR7ZD3G4/9UvvQzeFS5CD3nzrl26PUUSoJEx5EtMo5iv6O+a4QOgv+t
dMVC1MqqnTUkGLxvEnduzFlTSTl1ERRVG9x4bExBwfmkRJarsebHNQhhglGNSpXw
5nmw+1KYDg8WK/7BtEVNMVruHYxB6XrGh2FBMP8nZFU2lDqCNMFwhAizci/sn8Rt
5jd/HaKw0SvqhujQc0kdpJtYzVWwwWb5ExT3BXHXsEE3qb+4GpqSTFUNIAs/LCr+
yv1R0Oxb44yiVmI9jCG1KuxA/cALzPh7qV5iF9uIY9IxIMwtQXET54O/LAbmpvCh
4jRWUU7aWMoIO8GSACeKPbSFPPYeuEIFl5kaLY7rW5vLdVLarmvWIaZck7G1MKuF
wOVcafLueclWdfTR5dtyCvtgew/o0iKGwtAJHeAdltNlzMVFJqAhx9DjbwTBZeoo
LRSK4s9VP2V+/j0c/+/2eHGIr/g7qwUrHRCiQ4ROatMBpQhLPlzWh+3wsY5HFs+N
knzjmqqfovyR3bq6NUyTIfxNzGp8dY88g2hdFzCmfFzsB2VREXs7LfakTei2L30W
82cXGV4fuAfLirR1TJ5yK/w5Y+fW3deMGVyb3CY7c6oNk5n1o7q3+RNVAVkE/Lra
qeoQDnwe4d8rnhETzH+stwFqRNyci1EkIdstX3MTWAYhp/ij0Ztvupwqjp8gfPYr
V2KL6pXilGLE87AsI/RW26of7ZqRyb9os3yeGLedwmMDKK9N5+woIpuCo9+4u+eq
/jw3ELYBIyBfa056Yf/kTn6OWP73GqOBHmbx98ZmdKSaOBT6AkqBMxNc5poQX2HD
GDG0deeJ+zDyL7xTtLgfBdkn17D5I0NbgauaN8SCXh8OjFDNfo2n0sQcsTeNj+uD
LjlF7U8xHe+AgDz8IG35uR6CkUBsmT5rs5K/xvtPFA+NKKXpUy6kSH99S2o4f+hQ
gOS41P2xPq8VtokGQ9SHHgw4MiJy+pVtlP+/GpSWH/vt/FQQZVetTmUW8vIrQwYV
/k4fgbczWChQd1hWtfH5jw8tEjvtpcVVAVHwykNNw9J6eF46rw1QsNC8OJt2V6wl
3xygTYHUWIVVc7zDlcK/GwhM3y4uKzxjt0d69bzPhypYQqcfA9WgC7my21q2khtV
oyUz9mheDBB+yrEOp8qnNGkn0rzbYyCuubNYz4eNcPALgEj5hzT6lQk6dXf4coP6
HW/XGfRhXhD2AseCoQAVXiGfmrU95TFI73VN9Ae9loWrcdHxaq0IsRFUdpcUix9G
HvwzeoVhT3XAnHzwvIY0R3btuvoYCLT0DiKpxwIyPIIm/B4YEFMNWb7SDOXqLF5e
ZmIhZJ/4KhzktRDBoJ3dBlbhSVXBFqLh3tdd0EbdVuSzsifn+33DQlDkaSSSLgmR
XO78QTJRN6UiHf1ocu/Psq+VIFnasrK+sWSHHKmQawDOpzk7Lxectl0DSSZP5kJq
F8nx/t7pf+Bk7d7WCkr7kRfQMM98FkrBftrVpIXbeu5BgNlj8quecrChTEEyIm13
W1Abo6YE4OZNISDeLQ8vkl0k/sY5RUumedDE5WA4aVqf/7BxWpV1/OCDE9xiVgZ+
sjfJSx2qcfIVJYVX3sImrXJALgQtHw8BO9vJcLDQdpYfv7Kgi67IQnz5ce1Cbzj3
EL1uUZyyn+oVPL2T5lgrOGJqTr8k6hmE3IpJi0OOvPHNXto0eYQhuT9yKfONXtIc
o4ZUBfiuEoUwH/AKiC3tPaIrvPP1KNrGdlAVKrL5fpYoqPB0fXp1fatNYAK2KWs8
C4ZtOY963D1RYqVqvYGmS8BcQ1JU7H9QM/687Lba6qOASx8iuDHi3ArmVjMybhq5
EZhNcNXkrzIbTSPtqEH+4PmK+Q3ttETivjUjiYSGh1pRF2KodMRqXmz1u27CWrnC
iQChOjYrur2OswSsQBWmBK3pBJdToV+BuXxbwnsg8lajCaXhEzgtYRtbpCqDEqWz
4WXxrvEPXIWlcpFT1f+eT/wl8shZTOYwdFPsfnkhkdeunrEAei2Xh6OZNWZ/TAE8
GOkGfbfmqOfySCXUMkzYj75a44s7XiRzpn77vpQGsNnf0JmQ17RJfnIAWeImJYjx
PN92bXpdZL926z7lc/b3x9IltFY/5CnyGfg4X11T7UWW58QQDBEN3iX3BweKUoBL
piFuofeB/UIJP97tsMmLVmfincFVjpzvaOq0Qt7vJmgp4zkKime24Z0nXGcm60WF
WCrfU6eaX2I7CCCQ/sa/3ubbGxOQTavdMYZFaeoBI1/DUz8BrqKkUlWWlyyJHpOD
5nGYgq+Qim0WGahfRswOb0YVYgRzH/gDYxjLO0j7t1Yxp6X0TR8eZG0KMaeua3NQ
S13k1HfhvZhg/VIVP70tmGRq0tkJE79r3C45jZnPxKR8UU5ubqebSgd4nu7g/sth
eUH59QlmF3S76LSHEHQIPLIMFnn0htwPEsMYYgVrWUIbcsG/qP1qGYBEicKOiUta
/qU+d/qf9M5Uujmjj0a212oCQ56Io0zFAIQWuE6pZLEWZNag08ooPRD+MswE9uh3
nr3TA6EfZkG68EHRzn8TqXbeB3g/1k/Zmj2pzAN6k+PNH/UIzGKggd1lIA6PG32M
YrD7DODGpqbkDKMxRBfuR8g/73UhJHYaq9Y4yoeNxHhpVhlg9N32JA41i2R6+byu
VJPEgs8KCe1u2HllNcD8Xi+FONQqVC+Sa8vAaEOVgmhsC8k/AAFPReiPDCGl6igA
KNiAaYf/rFD9mLLw207Cj5eZuBttsZ6RppNekstGFOUywowbLKWLsXOENBVn2Xpl
YfeCF95nH/MvTAdEAQFYcrfoamHQh1eDDmre0IbJExWybyJNWHSNLT1kw4hN0Ezt
KXbvAFriokNaKDUbT4F4Z4yUyboVlWYMHALZd/0zCib1jMVIESLSb8PvpvRzfVNu
c6/i4WjRzs2VvrH+xEXqu3XiOPY9GJGxI2pKSuzciNki5h1LB/FVRq7aloXNF3xp
l6n60qlHOJWNMry5SRnXosZKDxfVu9oy3BPnGHw24nGQ7BuVucubjSgaiSEThTkZ
2Erj5UE2M436Vji75/JkMxxpEFlvDqOKLP7bsRbemSPY+zBDrkOt3xsu7yCG499n
0pSOdSTMKprN0RLniB13uyUQHNokwAwaZgbAEnJOGSBiMenjcIHvMKROLbUj1tkG
sPQqfNrNOkX041/WsXCrk/awqGnmFcQRogXEgMlRH5fSDpsmm4APDbPudVhEJALd
+gDwhXpYWJVIu1yh7Ymx1hgGekE5V0A8cQnm7fcswLIue271oWfgU08QhI0B6rqJ
Hp2CtphEZoszz+bjo2dbFV5NesQd8DeXbWURfZfmVEZEQe0j7D43BaPEjKTFULZp
0wg/wOqb/DGbHWceid68KQxynelQUTE1pUenIHRgMxah5SJKTmdzRYVSSSvhp3Ji
ebWlCwXIJQzAm75Y2Gp4gT7V6YG+xH8VaVyJgtrB5TyEhZB5FBu7u6Vw+5hzQOBB
HUXb693HsLWrzEPW/wRmP2pAtV34WYY09VaqtFXEJyvGjV1IHvCSw9to88k509/G
ZmESHPO80tG4WxlW3DWDXo5WITCuXqMvTbViTOvsOAiLC2uHlf38lnlIgISt2ZCl
0/1ZTbbI4WcbT0jwHmmy1M2KAfj4tI6uMrOHvpta7BQ/GW942HLyxKUiJLbbBE16
R+/HBf1VdcXHE8nZTWIZaf8jSsa9N4APN1iXn+dsbO1IQCZdXEx9zWiSWDyBiig4
Al+c7D+JJEDjJe0tzuG415grIj9NGFbjrabm8qFAPZkftD4NORS6cbCL1l9+dCuN
TEV9vosg0+3e8dB/2rnJUOu2mrpsluwtFDwG2BIt7Qhy1+hgKZ2ol9bjOZnkZV1A
E8CZqG4Eql/P0YVAXoHd67zYtiOPI3HuI8JdJzDdncLEBqDX0CNC2okGyQX2Hb92
/ouGZHwuRIsTGxiVy6NtYuJ9CrShlKFY3BTJ5cnJN9f6cc5clV238WE+v+WYdnZm
VwXtqlVnoswazdx3SiPcNV81+Bhu9U4+C6Xj8O+4xJRkHOm/ERRpLbjzMd4sxJcc
0XJ6HQuBn0sos/kKeUQsEQzCHgFlxEp/hHBiApH3o/zDvse1rNBLblZs+zspr/oQ
M1l1eNyp+hsSwsmvb2j3Qs2hwlCVQ67Txy4WT7QPtqGDCBqbAZQpnQR/Rs3o+Dtu
8c7CCF2F4kvP4k5hpt9Rz3rDkWL4wZebasgBubrSvsu0XckguVOCcYzxf+iVtaTR
pdpk6m9hQexsMwEZnQMsMNeeUgxk7cmInuzGol1J2IyqBRZkJwnEdsDGPlZQfYXa
FPfQJqtv3a7x9K9TkSk82xinSSOFWk+CEd0MpJGcCO/fVHmbpMZsF1LCE3ZnRJ8v
NENYfgqLe+BEsZkVJCeNdAvdRpFA9XrqG6txZmi0MJMIh22wLS7ccBdVcZ36+hQL
E7OaJHXjEXfxQFyWkNH0R/4RdMgqLds7Y3gMupAbnIRzMKWiSgPv6fcIJA6u0Id4
g67M2mQSRpwgxcy8YYo0sxmAGhGKsxHhy5DITSc7Zda1guCv46o2guNU2punlckK
D2YTrqsAox7taarLkrKyyWGk7ezK2Lrh06E5PXeQMaEIGq86k3Zv0QUXvUYGJ/Qz
ZJPETBDLjxP5rawdy6/dFIbLv/IadN6sggc+iiBQv7I0sstrJvAvlPBJtWmo5HQS
qin/UcLf06iea32CLTKxRd1bxxQqgsTmnU0tTPp8najegsVXQNU4/FRGtuIzdLRs
1rmnO+sAjLoQghr887TAXWCmOfRkdrCegzLwIZNSfeEB47pywkAGDY9GpVk2Rrvd
rruYN744BkWxr53R8WxPq4YlKa6NHj6OoIzau8xXhTx7xDZ6mcG5w5eOZXQTfHiJ
Hn9N7gwLYM11qj/NmpGaEGKYVVcHE0Ok/BTIsun5Jzg5JdF6n/6NQDN5NTMRv762
zsCVgEIc/LLhl03izEGhXnt1Mf9mDPBW6F0B4vgeGXxB6mZkTcfah0NLo6qiC6si
S/tKeoKc4C1fVNlOrQjuXWzxAJ4fX9iJBILm3d5tspASymHxHCx/RNZqYsGGdtfg
fMVIYOHMpMKVn/rTLO3eM/DxPIoFTPwqFpbT7WKq8pNpaVzH/wH7dokEomw3eO+T
Xx9vd/cEec1kVc9poGgcTd3N/r051YnGjSzzdsoelhf1fwls8D3f6qU5zmW2mXyS
gsnXiHW/wmneQQTHMzHmgZ3botr02w6yjmT6xMYnWRek7+UTEMvoM1AVrj5mBcE6
APVT8SMOQlKoKvDB3BU7jzYzNeopBX5yBkHU0RMRK62SBgk0fvf/8HETGzcQ4pNG
H9IBX9rZtCHytKoyU6NBnwzcSxmq0Qk1qxwCu6qTvC84AJal8Ymf+qKaD4VOUXkQ
7hYNVdv8UZtDI58R/hCzEEGcp592U8AUg9foRfaTMuVRegHYX9npv7TXejiDdfXH
jB77d+0jCuxQsHxCG39AGTLGams5l3ZSHAkquUYuLbiz/GiYTxv0GY1UDk7S/SEK
z2dDfPbZpA4WqhpWDcJVfoM/WWEVJKwzfq7MiRL+8SB7uw0UMDJ/nTHzCXukwG27
al32j6xxn7WNaejMMYpuZ1xscYD5OGWNSXtXp/FuaEuUR/F9fYfQIOhPiOBCwTw1
TQiETWhc2Ux4o8H0Lg79UNkr6gq4obr0HjFsj4sKmp0sz2/2YSS208fp6ko2OfDu
dH+p66Yhx2KFZwCpczxXsMmLHcfsZnse0ovTD15+causquFsuxZ8mYNEPyKw3CMB
pemjgj7mAFqoInkBDC+L9DSov8tBPT5t51sL19RxSaeKuD7vQEzNNlRwCPXiNZl9
R7EJWZIGgCV2e9fvOSqzP+PH6XmzmqvggGUjo5+eOux/VE7XPUW3L5o5AwC2+TKo
eIH2/cXd8kOLrAKBBlZUqAs/4OKKfsatN2s0+Ep1/KwXM12J5BC1jQ4SzSDJm0wm
PL63IWxGCbVzRSJrdfWxp498LYAdoI7SwhOtOg4cpRivyX2OibKYmWOxZjEj2Mdm
978mIvy7ySCcXhEhTLWRsbEucd6I8KgikZnnYmzeAyNHEw8aeWHnV1/B93ws/F+Z
NRxmrDpvF4Ns7vUaPcBWM2dWAnybV63goSFC3VgUzPDdbts/GgTO6O9c1BkHxXnU
nl2MNdX21JxafIpA490ENe/Sn/CZ24aLKuGRMUqxTSnSWcTmp7pIKQcMFwQt4tgX
LAcMD9Cn8SmcL4YiejuveFNqBHXpy73hUt7sgYJ6z9rkL6368T6PgURdWPcZMfDG
DYWNep3YxEA/mPdCkhypRIARI7iB8A6OOQ6ASH6rXChH6yTqK4Bg3PskMO04/3Ih
XD37FOJ4lOi8ye0Csiz9ymOhjAU+IBKi8AM0QGV248KMde042xUVuqRby/w0mzuQ
VZqB1pSpoztl9j1WH2/VIBnv9G/tjtP3dMTVTyu9ELXokqCFwir826zwuO5LJ4FG
kOgkP1uExkRSeVlMEClILCQ/Y/X3qeQKQhwc0S9a07xlq+MlNajDrWHjbGXzBJ6e
YmaI+94umEE7xe+dx4K1g8y5E0lflMNGIsYON2+GIQ4U0RuyajlBvHKMzX91K7oI
ayL/xKY7SS5tcIRubjDAz03hxSpuXNRv7t/bSMTKyWFs6VFgPgofkpvLTp8F747K
MECae79Z+YJ0wR1VbuKnrGWKVgWWJoCrUMWhvKcrz5QHRC4iYXJiI1wE1a9FH5VH
1STT3QHrDi9fn5Jlpk9zTDIvh2bCmg0Z2WH4INGxPpsqRtzGeiTCEFzHvtWhMOoB
CQRuqNc/Pv6k3cToCR0Xy9ABO0cGYBvNbJF1DnPeDTDh7SarELpM8xSdVnI+c/b0
mCe8A5CngOoLXviSlPciY+qC6l92u4gPFRExWTqn3zRJKoKHjTFTx3pt9KuwUPZ5
S6EeZtbHAbLSiFQCa9Ya9sVT7FKZNYq+hGLTtG00WQXP4nF57bvZaG4JHV5k5zj/
pp5n0X20j7yiwCsxf6CNYD78i6AWul5cRToILmO53WqHS6gxigAWUAH0DkAQOoef
O/2ejCYCBwWG1IBSZpOiWk6zESOxh6cyBsbHspsUYNGgZ0SXM7RVRcbyHD/Za/Oa
FYZuL2yqxhP2mzQY6m1N/2bHver8YezsgFgojFeQS4u9f5qUxXIAco5NFQN6Zsi3
i3xbMzmZJSHCMHuAtf11UV6B+/wj1AiBZeqME5lcEG88sE1eULcq7lNPpf1r7g+w
tLvTlBpnTTOhXnxf/G6ubXp9iWFRFgi5rAWIPrEKeTXIvD8ty4KgLLlIqHplqlte
48+Bu2gq79QOB5Y9tIWDC8068oQkzJ+ECMSSgWnvhZvN/iPOHphR8cB5ycY85Td+
N9sHAUlA1B0idLJLCcDiH4R4v6x99BRmmHDf9awUf2wXx6H5ETYw1gQT7o8K2Jgw
mGsv+3ERpYn2dODEcOUZIGTeWFQ2RuuGCyCuoeuoIvY2UPCnG604OxvcghdXHCtD
e9GvIZqYG9yEPmcNMCj8BiU1wefDteAewwOITLo6GEv0RCw1u10HjF8UAbSD3BGO
TjRY88rjlTiGt04EGSAP7/3kkIUGTWtl0kAbku5PGhDjuWdw09a53nESufqTzxBX
6jUHItxdXpFpaeUlRJOZp2ZVKa9CWdVJ7rFl2UcxEn5c09EY8v9jElBcs+hylHuO
N+iCS63Zb5+x22LhVMjsFMXKaknavxNRjQ6ZUa9Wp805gYWHOGYTQtOuH3p6PJMw
T8dj4dZHSsIQJ5ltezjkLSaIgmL9qAV4Jk5Eb9NETzSty9658sSMrUCa8yiYOtfh
U2dl3fctPcwLpGEV0qPgYOR8zY3/QL4Ppu5Gd74iRl2NWx4tzIfR5IJQ2zqc9u5K
3JAOZO7s/UmR8r9eAG8/WFdMorqAzw72KxoaSPxXzXRrpJyvAZ24cD88VxmnML5+
kXWK2+qXoJ7+UIxZ4Z7x7VSVplCVujoq3I5o2lb47HoUEc+KwZLEjOyp7aWL5ouA
1vjT8eBL1+D5PMOy9CLmOGVmQ9L9M74hDmuF4u5FwBZCdD58srfXV9vLcu4n8WcP
tROJk0oVCdj3F02/A/2YoDuTn8WXU5nWhDn/e6GTpsubjZlvzIufP/1j6Qw8iUWL
be2B37YOy0bb/2iXs+Xz+9uFSzMo2ZlNhZyGujLJcL7Mhn6vWM8VnaeDNM7D4fYb
6PmSS/BRgtK4/TkReuBqZsibLm+rNfTHoJMxk69VpKq0+Opdg9EyhdfM6R2Tmkc6
8OiRmjhZauMnqDF1GCVtkUzXm2Ur7SHdY09i0uBsGCPQ+NW5mwovns78dxb/rWxI
Fewn3SAyitZGW7MCSvFBaGL6480nUET1Xu56B/0SL4GScVcl8y/Ek/HXydSFwPoO
di7t1CGV2sKcBbBI3G25ewytCERUgTNKxKIVRzdp5itPbzs0l9m4fqTrhmkgIazz
lzyAB8caofW8rtelj4qT83ucRdvS5ZjlbNSBL6z1AjdUG0WlyxDs01sZsCIwXouv
bo1xE2ufg9vNTg3JhIFPUJMn5BqS99DhlpSmYGS8I+zN7r8fuXuvG/WmEzluddw+
a+Tjj6Fk2w1gzgtrK1wTR9NBKAsuVX1b14P/WHYrAUtlDf672Qxgasc1+rhJgBoP
jf5MoDQcLJpAylEVEI5rjBBsMcld9sdYqvD7qbA3auaVvGmBfj6S/sxSwNp5BTqS
fBOv/ebcQhUTesRyxpDZjtXNtlPOsVybVy8YrCcYq6w7xP+JTFxVQ/LxGAciaw7x
yR5Y/CoV6HbusWYjp5WOXnGBV+56TuUWlWn/1N/O/mgEEPG1si0j300guWjM0+dX
T9UQ2U3dvS6jAiBFJ9epKxRwAWs7C6E6skcqwQTALQBoQ/+CBnLhEyqx5yXCqu/d
jRr61KJpLDSGxNaRR6HtNOLUm2eKwZyp/dEmr+Y+oixD/1dkAKzjP10PpWe9T6WG
RDV3Jko8kvIV3t7o3OqQrvKYtBElCiA87aPHiM+BKNllKnGIbGHu/0KziBs7zMLk
dTiXukI5RnQeRqtbRSPMyGkMZJ5Kzp30rjXaJKWGYQPoAteni8h9/l/OwVg2F+WS
bu5QyT5RP1UkfST8akzbXSRjwAyklY654cjlziz7Nl5o+C4ugFF6oo5wC0ZIQk3O
t0Xtll7EfHp8Z022xZPgp7/nsOhdXQIY565zEL9jcugoxVEmRHpHP7ZhPGC4/jnb
nZG3OgiVBGh2WZJBwep47Rpet6ijoJZhCC7BOSkr8Qa+x2Gt8KctVgLOT0S6lqhF
9VG3mNuut6SjcM53NQb9uqMPzhbRV3TUfuDM4s6ijHaEZCOqUBJ7/dRdZaJFoj6C
6u1RdiIuLNNscz6YgevyqlyVygZ1BXpbfbZzhg/PpujRGJhBmf6GY3j9SH+u6cvU
vGLDucoAafwgDHNPhsZ2fTTd6w4a0/dgukdhHZ6yIUnUOEZDuKGjGoqgigrFcQVo
4bpskd3yMKYXyAgcGTKoDF2hfD88KjjHcS7fI4wOj7ez/DuykXhmkgoZ6FJ8nuPM
8u1+58qOdA6E6DxE6EGq4ts7Q/eQTmsCi0qekYNq1peyZ5aJMzoEHNhjp7hj5rax
CTC324FLNpgNjMb1y9ikDNICWKA2ZtTT1n/7ulF/0ZWd4YjWCSJkP6V3MkZuLsdk
LVKx41aKDTfFBIGRJ1kA3scW5f6xJie6g+Kw4vtIw3bUCrEtlAwyFLPZhF+A2B4R
VmAXDkYU545OCtl9lce9vpw78zv/EjuEEXAxQdpq1NkmKuuwzMzQHujbLum6Bn2L
OJgRbv765L4qYrEH7lHr+iO/woh7wYoNgf6w2CGx367Z6g9BtYxZ6MzGE16xr/kF
uM2b2J/QFB715PJPGNfBsVApIDQtuCj3EQSvYvTZsZ1ZAUI6uw1D+BZSF3mUpx5T
1ICzk6wrKYpuvqwify+2MZ12n/4QxgNw38tayS1aj9IpMW4WSwEv7mvqyRL8MGye
+7o+c/B/fgx0e3DMXS0mkUkg5XU2zLECO2xvxMyaY5k1XzZ/RF19srRlghiMsM+o
Om2Vvtmp0O3keJLdn5K2RW/cc43e8iaDKg6of33uv5AHim1jYE4szyMiQta0Reoc
xfQ+coOVMa7RSOp6goSq/Q4BRzze5TLwY0IE6B5XVH3GYR6hCZY/GmZ4CORL+QB4
NJMrCVc1pTGDkEB7o/cpxrzbGTIurK9mJ6GCmSUxsqSf18jDBZArKmDEPWXHd6SV
vJcDjTdjeCkR0jAVgsscjbp69DXE0pkHEAB6Xpo1NUJlpCc78ilHwmOUJ4qjY6nM
QZe0kHEZE8QnisUMMha7NXhWvfr+2x1jhxsXXpIfpJo/tN3RuF8PuyrhCjI88ZdI
pFhJ2S4OWgOXNyDHAuRr7upKCWtV0dtnebH6ep3XY2e+OcPI2SLcnHR8hNYCYrHC
M5h3kQENa1hqAaU9wLY0q5XG7908W1pY/ugTXjGBuhVr2e6wbmYt2IR5zMCCkVri
Phd7fGXHP6wLXkV8UQ6GvLHOF4BxC6jh97LYpJzrzcvCFyHT/bhVueJydQBSdISN
LzC10+homd2gkcgJzNaiaWxjhu/Z3X4qwQ4Dl2aiIf/gQ6dRGBQjxmL3Mtb48OwB
0XKRq55/t4AMH1sOsfbzb14zd0RCA33fjz+U2CmS5jTmoUJINmZTXJnmQ5zU0xkd
L4drgYqK4ghZjOmIJ+YJM8atr2BllZAKMuDm2wKvVfnECfRzgMS4lvBs0u3N76yD
nqetKMqeo03bETSUp4m0ivW93Hh2vtzWSqDH16sG/QhiUJ5HYnVGHKhK2jXQ3itm
7x68QNWeNBXlczA6XIAisDG7w5BZVKxL3EknBkaiFlLv3r3zuoaBW/hLzVcTHUwt
zrfdpGrqpKbnIon1TKTp90DKNBF1kCimHWF73fiHzDdg4HvhS6BnMUtURW3swrzD
T3dhU3fHyV/PI/hZ3kid039MzzTmcV36s18aplmoI6wL7COiJQoKrpv2AmV46sCz
C0/fFUJCElsu8UtY/IwRkRwK53PEjO0FiwOy6UG9+23UwXdd0tizi9ns4kB+E2fZ
WH+/N38UJM/opNeIx3v1qofnhC1765NLBaX9dyt6Pb/L9GLDcZmTW8LdphTKGy8d
7jyYf7xFXto2Umkuf3kqBWHZbfL0sIiSTbu3lytrqfvxqu69DtU9tKF0rGCmNx0C
fb23gQ+np5Oh/bmGMrbVm88V96JPF8zpDJLDpp3dvOXzUiV7aSg1qaE+RUQdBu6f
ODP2dIZzs+dppjFHvHSunRdp4j5Oea9xwlzWJoZtnWK/H4Z6UnTmtKNZbGIhwft4
zVQd6BEsnzTKAQ4dD10wCI5r45ztbiHFRiF6/OzwzHIGiAjU/9UF85b0Isgsjts7
ZheHg1wSwoVlOuyuJB3+Lxbl3m9QNkJ5ko3AB6UKtrWE6W8Skw2F9ZwYTKLnS/rW
xkvpzUqAluP6dODBb3uLAAjsxavZm7cyOOFQQedhJ04fBqkR9x8zaN8QuqiBnuTo
hxUwIXbqQMNd90mgWl2/XF1EEqJRvks8GIiH1xD2WRIGDpgRZ0IWn0E+a7KyKfna
U+ikZ3NiV+xPjNSwkSN3ewdDFwaZSmw+0TxLRuUfj1eHDa9knbdb8qlDaE91xNaI
EhjMhGg6HcTuBcql8YBAF4XL6+IRrphj0LMQwm4S9hxI8EsrbN7MkWC8hXOUb4hM
Kf/CcaByQg+gWaiK+2kt+DfH0AxL4ctiayNgK8OqiPwkOND3nghnqiegu3MYzSWx
NI6OFLjtSIagPK9Bp/7GEoo7PUQ3Z/QHPpj/9VS/qUEbrkKBfpXSSPcnt5mmKILD
uzOeS1KC8AGv5+GPsjC4aw2j+ZyQzwQj+6KHCaVW7R8TnKLasRQKlW6gHopV2IFB
x2a+VmGr11dDo/JjuLWc0aHmGyObCreoTe2BB8iQfMgwo83WIdM5y2V9XnuBiOtZ
WevchmI/QHMegKDo2se0264LJcCMOuamcMIKpamr4bs/uUeUH7puVHF427rE2Kbw
rBkIHLC6K5JQS0lK8PqrkwKt+CHfSzv5Iv3jOz6xuQXKSqlUg6wBMUten/OihVO7
7JxkszicBSslaBgfpXNKCAwlKrmaos7SW5kohgzwobboZ57bgtCiNsanFT/ZMBRr
cKPEB4FRmBROxWGgerx0Lw+BHLymlc+RrL7azgnf5lumJA0/4mcYIwRRH+oqFhIh
Q3Pv7VgSUuEAjZZexrH80penqbADX27fUWZ7lTmgwa/rTFdeOSiN7jVF6/OUQsjX
4EYtNJMM+u16jX5Wvm1Lbi/dAnSNONyVExsVczgMyxhYeMfgXFdxalyehmAdcle1
QytF5CvNPzibDOU2x914BuN4Mjj4YsvJ6gSyU+Em0as2yBQDGIyh9F+pNNq6wQ2w
6oClMJovXctjz205W9oTyb8Nxkba0u87gp6v4sgZcUkE1fV8dKMJ4MeWzf1HNSVs
42wq5C5gnAaQgbrPbJVZtM4L1vYeO+oedv59hC6UWMNzlDP2Fm8bWYmYR5tlTON0
lklSUofdBlXN8o+TDJnhhoKJ/8km0DUOI+yC28IvZjSjwp4pLzmrD51aayW1kH7F
CYmciV7iU6enlJTFB2E/Q/zHQS2M2H70boysQNfoDWplCXpIaHoO3ZIYZEEUH64T
4NT+ZzOlrdq1V832KrrJA4+RifmZyM8Nsb8mQAFurDSuQ51llyGO8ZjTYHPgmD7U
NDjTDjzmzFec1Pp5Fz1as5JgSOd72iqc+8pmXKuRrbV9a3vNII9N7hFMyCNWyhaB
x0KjK8o9ye5L94ERdQ0/u6qM8dI3t/xzgjr17rOtaO2t+5/NtuahoRJ8y3W6MlTL
VidVuuKgochzXXj8qLzbe8nDAJUFmdNz85qlKN0pc15tvhJwqU7ZMtGJKBtIdsgW
BA6LEyE05q5SJpxZG+9b/dYGzGvRxM+HCPrNXGq/DqXuqgvgy5PCPR7vNciqnmku
IDjvTze9t4B93l5gHf3Rzvn4BQdUz09YUQ/V9TeyBVjJqo3UFTr/AHjz9qaOAKrE
XiQnpcIFkMvLTo8rvOZzLhHsSk2iiDVdZ0J8g0H8EUkLOoIf00v7RNrSLwFU4fde
gso0fD8rOYMgtadhe07AFq5hiGXyVsFNhiujEYXt13HXXspKQGLWQ81+gXS0p60j
VxdNRgUN2w+Md73wfz5c+ES9q06NOo18j1yQuY6OvO6xyGzzpdSmU5l1xEa6bT8E
Q9koTlZ6v78qeEuFG3L/oBOf/et1UW2jF39sb20DVdVbEVJZYp9T94+ooVosmA10
zGATix/UGnw3jmEBoY9q9S3zQd7QgnEgbWAiwI4YUSnyhdZ9s/MSNjCClbpXNUWy
UvMOzTIuA1qrJdvU4V/vpSDxAzraU2ssPXC0Cb/sk31iGcqbVKdZ/rKNtKqjk2wp
f7TJfHUXwxQPWd39lh3tCF8JsJY57Bq3EEDBHvM8NbK+h0+ayoIeVVl9I4dObAPz
AKOBRNsz+RIUvuOB0jD5lC7c3Ic3y1fKA1diRlt5IzryxTutRdRZAgbmZ+b8N9CK
VY8Yp2fYXwy/KXb/RrH3WBA+G7QsYaUfr+1t9urFgjrA8cNNtWZI0ZOb/sppl8jP
zzilK0A++gj77v7EF7eZ9zTY/xa47HVtkbeinrpjcCyYL89M5DR0bBOLVBVHDWLg
9mxs4cWrDA+iunsH4/qu9DtqGafeAjqyA1cmNsQ7FpSRx8e52/sYGoRCu6gU2WJO
qcBrPUp38h4LRHItAL8j6KgidJ5sM1iDRlvoQIFmZnVFIX9fFw5SjcwRgcRngVS3
nnTQprymu2sh8j/f1jp3P02WBx32FwC5wiGF6vjfjHn+eIWaCiLADVMxHByc1z9M
UCXSMaao3J6wXkBu5/IkpI4ilBatRJq/rAnFqUhThfNxT1hVjrGrqa1oJoBy9q0p
DeyJspDzvAumbrUPeCxLDt1NwrUpqvJFF94k7Ywi42npgx82WebryXVFdHmZA7Qi
YSrl59cJGeuRVwix2ZCsocHh5AaQ0ShmB3WRTRzx/1PU49NQT1PqgfajAZrtOoBs
Xwf7pjeElT8eblynkTluvSgP0bCSvddGG+3tm/bbN3AuihpQN7jUqrI2kwu7UMSQ
W2bx/RODObUa/fZWoGOneuF2w5YrQn2/l5hWApOuN2CXllq6T6CSfTQsE/b61TSm
YnlYjUGE5U/+g13lYCMC5IspIPYoJ4CBd5EBICGOND32jmxt6IwhFPih52orAyFR
GrKlL6pKYPiKDkyZu/iB9z+YEikQMhzMoLC59QtJddQqInw2XQINygyhyGI/MdRa
A+SYCFUAJwYFdh3GNge6AfVAQ9erL32Batfw8iaU2Km6FQvEHW6d08fO8udP/Q/W
eY06BDyjYJDkZZ5xrWMEhYFZW8kALVRHhj7B+ERiQNzxeidWu1NEs3E3cKDsEu3O
QedMzvExP6QDOji4zJAb7Dua17TmXcyWYiafS9Ai9wdZZ+w4tsnO/RkJyuN2wsTu
HDVifjK78tkNgyBi45db3uvS0Zd9QFYbyEjPNK8HICBXymJI1IbpBJlZ8GQCCDdv
xD31QO9JxidYjw8VpVW+3veGv5I303yGew167JIlS9SFGmeGOmm2sbG+5VYh9oQJ
UAt6a41OJTLO7q1b12/0OF2AdEWdKw9G63jpTz4kvUn10T9o+1S6/QXMyxUlj0cn
5uZhuPAhC/3zG/trh2QRcnqRn/CMSYv614A9a78lI42I54AzUPPiNDQSXmTirhgT
YTlqTyUksjkYdNezUynD6C7eKnH5aNy+6vhoa4PGVPJxo1+8an8ihqypCx6T8Rlx
zXLupJS1JA4JnamTmtZEAUzVSZRM+eZrfg5JIn+55oQqZDt6S9txHc29vC71CBHj
/vFXsahrQM/zE9PnezGBC+FA+ALCUKcjptG7RCf2jU94O6klAVnzLiylzMU6F5Dw
nZ8JVOQBLq/XLLqSu6mU2BHzwNd6TR0LXGXTTC4gsGwH2I9LZF7SvjmwCp9LqnJM
izGqFG/jtCnrnD0aRel/C1oJ5u2JqSSQF2UOZrnaDoZ5CrTIrjT5/xUn110Rt7Fm
nB9CVrV+dzhuy8XEymBfVleGY2vUamumApyaDgTJtB0O7iezmv83RDSe4qzXvhgK
5OHnRiPzijzEAhNnhKWyzw9DRylQNc6qz8cbyX5OBHMO19JCiiKjTbvvatKnD/g0
fnxXfgLlo4l2WmkTgrw9app9AJ62Vm1XJVxy9Buj5PgVI9sN8qSkDA1Soq9ZJ/qb
DmlJat4R6m9fWur7EiWahwNHfCkZKmNmvGoeVCZWdtiRMm8WyoEwsJviUW0jjYoO
0d1xYz6T8DT83xs5YAsm3JdpHuM83m23wcSbQTjMEjBFvmKiQBULq0FNW96Wc/sx
wc0puV/Um7NW4miDzRk6DY0KqtEI9OX83T4dn9ux6WpqPvtFpe1XqfgcdYcRBVFe
uujO2+uA0Vw4iF/Gt6+LrixalLtGeU5owTzpQ8wWxuV9a4GRtapIQpYEgkpwWKBH
d0VNlUHA5ghrGdYCqAWpv/cgh2KRs8haYFowf9yL91NklCGkTD6r9AXnp+G+sXit
qvRJXKFbeliwGEMDKKf5ecQle6noXD9quYEdUkaPZ6gaaJ0gA90xs1J8/5eHftjf
WkCqEBV6UPEMw3f9ZDsCUega3PrqQyAe3fWNi3oHVYQKnJujKaQf+wubGKZKQPda
2OhOPDiFmJBevVd/cOL87ztUdeCHaRUzsMzXU5hhAwSerLrGQ+OtMdO/bVAb+UEA
6FicgmZjiBh7fLpyyxMZIh6qm5DpdA0ICH7cX4QiADtYvstOCOCiiZZ9bOP1PCyi
HiG2epI5BYnOvKV3MyDsoly/xD8+d1jThGg+KIe46CGeZjysKkkt7lrmR+GVsQbu
6Hn2r/OwvR6R9Iq9GgIlr+xZXDF+ZVsl2NyEM8E6HpbSHTsRL0zyWpQMeVRlZg2k
MPRX/7KGKeZhfYvLgka5psfwQvXloyp1H116C5K/X+IoGF344w8hoXnO4K7xHZnn
WpLHJnKYuJhVGAYZ6o4UbmE1MkxTFQu7EdTd41NHzBqQqJiVpDgFAIXBNLVgsRM7
kGPjd9umN1K1B+DMeC3E5cOLr2Of+Ru+RSWHXHVC0TwrY9NbbdFeB1bNpezAskZR
3r0Ksm0OGh4eNpuf4iC+4hMiMPyv2m7o8qJFtb9d6/+2zPtj3CUjS09rNIkUNTox
H1GC49eveEq4eXRCicGdICkB22/7dt+p8ftt2rnXBX/ZGgrqBXkleyqQ/e4Rzdi+
P18iku7VINYzcBm/xpiMo1Q2u67942sQtG4XCv2bm7Jqa44ZuMVBEgdQWrEEIhDy
RPK16/E2iufkqs4waWwog7VxrVlzJUjXcqzhrhMVSW2KJtzbPx5tY8FOBbeHO1h9
EAW50UNT3vtmzVOJoxKSNO49rWteoH1vWoS03u3p6NPwPqxf6c/e1i5O0wtqb0uE
9ID1vU714i1s5SYEv8M4+2xzE4/ruSI50ffTt32UXDkOR0lUXEteizI5FW9LXvA6
Y1OqPa9h2vtv5VANRBBwJgJzyIZSQRiVifokjctpfQEZKI1riuhKGX6qz46MffoH
J8sTO5L1gHI6BPwHgXi3Zkj4VRsdp83zV6RFnuFTwyJOe+f7+RRr12jrT2EPJwNb
DbdRdaQo1GfSPUouRjfI1SXi7UupAfFYfmtV7TUucyGG7gPreBdUB0TUemI7CzJL
anKeknhiKsbu2PjVw4kZ2Pcm9+L6DLWMRg26+nNpbjSxr/P4gR0+Kfe4rSVystav
CJXqxOnrCxBCOVPhX6fXdD/SLsKDMwWMD/1eCCOrcWKdFekQI5RlCkvd67UKcKGy
VMQjW5vj0PlaTTMnQI/VtKWmu742SeACcHkbWNvhqPpGSNKXoFUraJjDZBRciaw+
E0cyYurGR0SziN30dj4s/akzNtoVSiu2ivCCul9GDv7xVUaCvlZJZx4z86L8KjEj
DL1clRJvSJP/ccydkxAe1kfzHJby00Ta59WDTt1RwiglSXbmCE7gKOZrTL/KV2S9
WRPDvfucrkwVLXMsqG1ySYwKJuOixqjR3JAga5rtYRGu/X7fvRNf3dynjCN1xmSO
J/kSEyi2PzjYrWidUim1WUc8XeUsBlknMnGiIZdxM4yCuGkzo/DZ+N6jI2g957Qt
NWKBeOMyVM21BKIBC6R1C3uJCmB1hDcxBRPgl686vdqWYeGfpMa0hBrOKk+bVWDd
DHRQtiR435DY1gnvApiWwdhucU4c1ZFLhjJA0cQy8S9gtY3KSsRcbkYxFhGZfeqv
4/eUsm90DDafhEHbUzLZBPResF9ZDWVx4S2+BfpZu4tbpYDT6TeAyioztMP4+VYw
FYfoJ2GaqGfB3HNwElbAlM0hOvoyGbfllNYNxnBnXRc7j6lU16SKRSiEvsJkCfm0
SKUfZ67a/EC23X/W2R9fDd7b5BKapTiHV8DUECCQ6QIrklzMizmqg4YTndl+cvgy
Wsw94jWS+GznVelptH+xEioBk0ORpKopcXUO4O/M0/JwbFdY2/8yyHmGHRCaQEv5
cKTjeHBBKy7hRQZ8QHGah6HLgeaYgKBvsjQJFz3arp5mQTLMs/UkSViZws0NadpP
YUdGBQJj1DEZZDXArAmGDKA1JpRmJCOCf3+IR70FGPSFTzseiY2MeWxX0TTp+71r
fW2pjqB4IYRWXEO4wogpzAPhv3hFMC1WsldYFVE/DbBKIcoIZtp2QtWN3XYj6Irr
+tbmAUC9pRRH7hyvKkTy8IqgjdYkHGgIuinoLX/NF2eMn88DsaLj/hpoJJBafYPw
KKYZ9SxaucT/W462SuIUh7983HYjMdxXEd6TCQmVSGAqbYK+Ha+cAYYpsISYaFgm
uoDvDJvLQlMEktHJxe1Y49BU/ydjnkDgftqZHe2rU55JJVLdGI/7NGltvCN/F60A
sd1a0d9FgnCm/MCv6om251Mel+cSTWsfFvd4fLLh5PE/BMFzwqpN722cGCtFT4KG
PhSiAK1FaURAMt6lZ9CrdmWJRqjDVAihMjTKaI+si7y7JF257B2fmR71sJ8JLu8W
zf9r5x4usfYzoh8sIJPgVj7aJBKrlM4ArX++WvZFYeuuFOCzbwwODnrVwPh8x5Xu
N0DeuWgW/SzGrt6oGwnMe/lDr/W0Mm2ZsT2XZl5iH2CW1Y1HQ4hZZyPjr3+5Cfv+
WrwKLOaVX2heE67J8AS7XaljB0qsP8YTGUKY1a1o/yow9K7XG8IrNQ3jK3av7g6G
F0QgQV8g0FyBKVyIdezHw06gNc9tHH1vBRZL55J7JGn1G0JieQrGoebpaoN7XrSq
KXCl7u5KZEDXb2fxAuTH73kKkdNpfKoBiXp00hXb+fuKcDF4neqgdhSpx0uMDtIG
Xidev8LSCVSPzHB/N533kfe1ct3VyMGQRH5RdVQLMaBea3jPgRfFDV8Ppzz7vu0U
Mj3C5CJovWRosstho778R7ikc2sRxfWpqJEboJPQ2EDXNh/ilHeNbbjxgWIpot09
IkXux0Mls4Dr/63PRXoZoxgXFlp4kZuQr7ac3ozL4scRxk92MSUgIFRUriIYAnD6
uWJ6S6tnRNXDSZnUxMfKDPXBceBGEZ8CbqYXHQM+ak4hZCulbkMW0jpUFJCUAra9
FajvAPn2lrmTYYOzmtiMkEHOIOPoj7Vq5KVvTx8Cul3L50CwZLRoSOkf/m17LMe4
qGjlk9ICB0Lf1ViHPSqLf8ERkf1+3raLI8tiXSAHE6wi/X4zRSwykIN1weyUrAyg
8u6QhKQTciZG/5EOKq1W+BwmKvHDpbZzlTqRMMxMhvaOkfYoiif5o/lBY7mmUcGV
Kradk5TD4PpkQSsIBhOKgRhygKB/35TMc2g443QYqnOxDxHxv2loBuXMv9fBfPm2
FpdVB8FihrLE0fTuVjoj+nzdx2hJ4+j/KE2lS9NhUrFs4zDfA7VhZtCPp0y8H0d+
6xYEsqTn9EPk60egxTKXc0Zb1lRhsukWqt5GSAINavxCEThJ0BAmm7dhKCpgBHt1
ULq8iJ3VneLo0KIDyMA0oh60TICCVTYcrvfklaTzk3KfLgCf/QKwhG5uBglu3RVe
6g9HYmoF22YRfOG9rrxMvQU/8014dId3C0AehZI/2l8CUkW9iEpCyhBED9bWTndi
+0gkfovw5T2iB+ObRBJjS3HYPip26TZ0oC7/fx/GwISIjLQD0bweE2Ack/Znh5o/
ozL8frDOxMUkUEQ71DnHvqaIjabOBHH4o8UVe2gxW+hTNMiu/KzIF3EArMu9chRm
47Z2qGAH9feSPpCFvuNLpJWUY6wTofl5aYQbiQIk4i4pN3rJjpNu0RXbXOsY9q1i
ahgIprE0UrrkEj8vTph7FgXmH0QFIX7BkOhPfofWnSa4wlEJuO85N+75FQDFUI82
+laqupSX0qip4cCmbh76xdZ+lblZSF1VQPh4b9IrRNJl5WchvgRL74bFiQYjTw2P
bXH5FKzCo6f65mfqhr8LihYJu68dXSkS0zqOpZ2LgVlsdodPR67H5gn1SsaJzJbO
jWmoHq1ViGFBlmvO3kuFIl5tzpFmMVidnvWF+oTQNJHZZowI/6/S7JbyP8GhhRH5
hOC0l0jUNpY9/C1Fac9uqgpRHehKIEx6Uxfes0ovewDZWkdU7R9NTtaQNV51gsFo
V+y2eKmLM0zAKeimmP+ZOrykkTTnHKfqOOBcDnAgYr3gTyReYRQvSqQLcxIh8mOf
3abXe7wg8lJ6MiMmo9ckwp84T3DXb9Y1hnNcO3hGYGEJyGo7BCZZ+LNELEEhcoeF
nouZBPjpgbw0YtGNanjMG015ewkoZT9il+7KGvvuYH4my1VYYK/Cr0yNy274s5D0
b/RcfA8OzmCYNsp5u/dzJsVzreIXFEL7SCKdlv/RhzEiyPD1CJgMIoc5+mU5jnrE
7glEGDpqNQ+XjEU7Hyuf36OgLkLlkFaj42RGgv+NAvhz1NqbEMv0M9xNCmxtwb39
TEmv/DswHNseCFR3thk1hOYZCnh9DYiHINoBB23xdUTeygZPHwMTY5sj6AsSQNuj
2/aKtzqj+IAMeeQjKDmNvBNmJ/c3Ww+75Bu6iK3R42gZHa9omaDuCj5vvxEKVQZJ
VIK8qJBkQyJ/nGtqBq8yzMRCKIHl8ZFlWdhBNHoxZSCs3IJwYV+Z5raXx8TzBq9D
TRYCzsIMUv5AFCp4mR1ni5Vqkh1dAIzdlPqc58VVAEPGhvbRgVxhvwfI34G5dE35
4WGqQMaCqDDVJ8fxybfLql2xiLvPYI0EW7wp3KgoIDsz5T9aARPSAsEwajz50Wgl
Eu6257St5SJZOOlxtM5tlaisBP7pEd0xKDufZr7WRBnDwbywJKoNJ8qx4Bwn5XNS
LYqoPPOIu+c4rcQ02N1cWAoLu1PsnMzh/CEj5dhwOjE1C6FVrVKfDi7xORLlUOAt
leON5HGHQ1AvYLiPyXgXRZevTYRTgiVJaFLSsP9pTHeN5izvXWT+gJ1yNe08lwfP
cZJZHPJ1Vu1Y4fxgjkaOAZLXXanWGy3GbCiO+lgjE7psSAjEL3Z7r+ZlJnXZ2JnF
Nw0RVmTrVjfqhD4K+pkVMWfysYoWjQyTO/eLQlOCKmR/B1f+4HmMaPXowDP5k0zU
f7zHCH+ZEt0eqRukspk1R07+/Ke6X2JQWceFeVHWV6Z1qegg75aVYJIM4nCjC3GF
/yeVJZBz6Ku03v20mZ//XEVmnLnAAyK+U0MOZhh74kkAWo6lIciA9GSTPu6FycFn
XJht1d+wHjutzFNMBqgJUgSxLlMgVHl18hC1qWFYkGnLlKfrym7ceRE+MlO5/ujt
rczFtmg/TzK/V8OMmKUNLm11I/oWSaecv4gVwhu4ce8h7dewwdBfcIjwykC6NrpC
2EznLmzkgUdtNEU85gxIrMaaLGWvtF4zWaNCplZAiB1W+vyvge0lTb1zh5F7TmXI
/hKs81ourRTH8axMlLm3X4cy4KC14CJj1H/dbmf5LdWiGkJLV7BYQm2fUg8EhjRk
ywUMl5Ls9RitzIP7BIwsLilVOpQf8BJjYRx9lPARHHyTDCjxdMF2LFfbvqVuF8lJ
ZZLj6W+6sEajwyVtfYlhk/ehFvbBv9T5x2WdOJpv/F6A127FWgH7PbAYmnGLutqd
tm7yqELeTkSYSGtxb1ZXe2ZfRH058YQ0Optrq96onEGPI7W4Rb5RpavYCY0v3QK8
MQ5aD2nqCzxQ1TsEozP8ARHPZWoTJAiZB4aI02VTM/NE3SDkpZ32ZiWUjnlqjoM4
HWLSegxRlRnOxiXNd63wiybyxIxEVN6gqNTUnVRIX8zGknojrX08E0yQTF6LP9CF
PGhx98Gdr2LxuVuhRsnjRIjhVOYcxmncMOCLoUjcYpv+k97GQyy2JlaF1u9jy2Zc
HGxmIfZGdu/RK5UByyiY5fwuphMer511WkJyfDMGCiTYUpl6e2IcMSVbgl+4svS0
3P5M4bE3RaduX+FUDGqO3zvNkXOmcGkqS/M7Zs/3zQG7CBBzVo1YHZX9+VNE2upE
rHg960yV8oq4EdwasKmcXw8XouuSAGGlXbhmMB3AHH0gfa+4YMKiuPfF7/x9oiFg
xdbICW8RJx2qm6Y7snxNHYc5uYWZZwV7J6HtIGlgneYxeI98Az03zh4TfxfzV8Te
7cxIboFNlmW6cukNycHDFsi3x7MhlITJ4bI7uIj1yjJtn4scfoQQwibEsn/z5xKV
bvNGaPx1NY7yO+YQ2OKdm7/YaJ94p5VRB3CLL2tRctA32bCUHbkWUDLSnRSrXcvq
Ql6jllvKVoiNROnPjsOmFVF8EG0hDEqJx6fmCYr1uRjgIaXx7VsdRF5O40I5O3JG
r7WLEz5tS8xb873KsxO7gTxBKK0MVoyns7JHUUPoSLhqCROcuZYH8YuagQRYwCLM
WQHwxtjYIRmOZnIQQXAQZXVxvQujNKpNXfVO1oULgszzxtOxf1FYyjO33LT+ZDrF
IZZvlz4oDaUl2qa0lOlQXetUfScNWY4iPHOqwPe7IbmCkEvhARzdrqYrjPu0vK5Y
1Zs7sCyDArnW+yTHN7kFDIVJTpDTQUuRAil9i1WioOaVVQo4WmaLG8CrpSfO+2Pi
YPDjLeRxVtJy1pNNq15UltwpIiiZdVSiF1pSLMs1xUtXt7xrF1crYSQYIOeGJ/vU
aJE+RylQCVWAAY62eIiHvcr8L6bRfyX/d3ueViTDTkskzP6/QFJ9eTFRQj+e5pCx
s03tUvcSjQ77FYavtdkmxxPhaoRQy/WE0mnv11WBIsD1fUp9RcH3pwbvXItx5sjc
ySYqoQ4yYJ2ndAhXI7q3jOvgoRGhKoYcPJ+5bPjtxkMCcMhr0uUSJFiRq/or4llB
JZ4uAWz7TNfQdwW2/wuRkdjk1WANSBPo6oCGle9DaVh4drmqJZGY2g1WH/cd1SA9
EK3IlRniRaLNFqetmE7lNddURlIIOYfob1KRVe9MuNEwQ/tCxLIsYyqvhMcqBOO2
2jVpKLKe72MHTbkd7zcacIjqoPe8IdBnZdZ+H/lzVbHEvx5Tbz7//bny1XaD6W/l
5SYdaUfJClB5+Etvt7fBd8f/pKqvJY25+2FkcM1ZDy/K031wChQG8tN3iLBkpces
gvgP+vBm42fFzNsyUZe3SltTmGAa5Etf9RgyGn2MUt30DZUubTxXtF2K0cH0K6vz
DabiJtTLGfu2VXNFNpxtLspj+Ti5JidTzJi/br+VZihmP0c1C+5ZtEmnq+RvNzHy
k8sfnu2wPlFQcaUgD+SgN9YmPfcLQUGm9gDCuLXIzzHcCk5zmGVxXVBFrbdNfVfR
MTQF28YMmKBuMoQfv7kfCulCuyMw7Oz0HMwEgUM5cgshrQf7ESOiCtDiXyIYHWJZ
dQC5hkszne76CWNlHdJ7c/9nBsRuAzEgAm0nJELLiC2aSZzvIVWoIwOPctktlpEr
Won0mvCwl1PmT/ANgeOmx25Sf9jjc1RoHwlt40rOyp4amgjPwNNNI+Vs0THR4NKv
bkXF5g0OqLvx7tShfZDyu8F/PBF4Bpv2lVRYdAuKMv2FwgqDcqbjO6trpLeCnvY1
/aaEMKjI9ivd70CN+gVz1ybUtJsOBVCpHukRSLB055IBv+hbHbBF08KO5xtWGF92
rtLkLCjE+gGVcfLjXYMOlU9R3zvjXMAo5OxT1Pu+0GYdBkBfF87xnY19KLlisf4l
I9jpTOT/YcbX/xMH3JhH8mX4uodoCH4LYa3SVlsJLQ2YSXmeLHKCnc8pYzhQ1peE
n+baE8RHkxWXlI8RG1JuOvkEuoTYgCwHxM5UxrI9wQP1OfU1Uxm4b+q9SMkBjgnN
c0SR43hbb34nYIQLoGoAebehDVPObsa3Svq1qKSPR/MJzvue92yzCdCBgiWq4fp3
V4y1VCTidXPS7gfS9GW955dHJuEJL+k0vEp+tFlfmOwT73a83q3nNiACeQe+XU5R
4qrhthQLEZYYmR3Lsx/e+i3yyBZaxkZVDLhJ9fSJoIZGb9vIM9YqO5a7W4gaLiT/
gb05G5S7uu7O7NU3D6T7+N4CHFgFJVinnZjpKiAXrvCVpVyDGnL2FpEXGrSyvH3M
x9TeoWQj+y9gNYw8eEgWNStfDGq4oIn67oVDN+7SG5/aB4ELzubHFEV29kaSyb1F
T0Hz0N1/YvGoujmceJHbz4mAGwN/kVH+zJgrj20zCRj7WnpVT6+4pqiMG9ZVhScr
UTv8dfCX+Iyxtcu60OBcklnyQzbdfBKENfcRxScq5X7Et3c25dtFm3Sz+2+LGb6h
GpBGDi2iiDwlmYn2UXZlG1KY5Eg/GUjdlblIzUhdGdLRRojI4MKjjnG9UHvj6UTn
0JYvEjTTd5cR9SP0ddN/u7Vm1gyHGVOlYsUBoBEDiWBqUwInZA/ZK1th+St4D4je
cKXV1jQjWOo/aoSzK041xGEjwp8o3NGm5GuNdmjUJwsNHGrzYjQOXwiMd0cQ3jjr
YrBslgV6rJulgzYdiK/8sC48erz+7d8eqwWQlf1kya8/KQ7/E8e6vT8DSsXA6h4u
jyH5NLW8wH2WS7GZQzIidRo5gLRA08wha4WsgEfpm7AUR5CrvALN6/Ldf5mEx3hk
hWQuKlYFMvetwigMwjywDrV38Q+83aq2nt6nDsLv7gD4aEM38ij36lGZ3R0Ce2Wm
Vqb/yWUr1EiOVJtVGQAkz2N5EcdQLPNX2bTThLmLCfbSIkiiyl+tZdwYyaUrp9g8
KG8yWPpUgjPf6KhoGNFxMs4YE+kP1nvvYOERHlQ8wa/X8MqamAKZCEfb+yPMPSbo
3tpwV375s6YSgpgOOwJMqkcUgkbwHw6R3peTRt/g/22gZR7LQ/zIVJsvZM+lXkLl
ApKtvhamki0j3tvfFnXpNtyRIPiDGEGE72ScaAkk2CT+k9JXvp1q1DMY7xSzDCtk
ynGfQZ1SjbaK9fqNMkFIIbNpdkPk5BRoiBogGs/GDHEGcaNhrFoE+HfAOC6wzewU
bmj1q7iusky2PBgO7VixyySzV4Otwgl58Xxsw/PzTM+z1F69Bec+ECWpjAhnwvYe
H87gGKDCBg03f89FD+9WBwrSNY3kxsSA8/PCxqucNoo+ViOcT08AGrrsUBj/iask
NOkkv+vl+7blpKMPjIkLpsK+L+yKAOa2WK3nKI94hAKQMVbIhjKH0n30xB9iA+n9
DT80femO5wyyjXYLtfYzTU2BUxmX8K9Ie9u1gMoMTmzICEdWORjiRhv0nveIb9bM
Ss8eCS2qLjbnu4Q+LN49a2mR/NunU3LjvgB/n3zDoFxOvMTTjVeP7RaMxAkOK7wZ
PJYo906R6gRhb7cKCMU+028Fa80/0IVD3n3mzBKqY7ZEsLAW6vKe9nNDPhK3rf8D
3a3SkDmyl3XlMR0dKpNygnxy1US70U/cC08r9uG3WsV6kjUq6c3ssUxLJXhm9PxK
4weQUMbln0H6CApSnlpv8vsdrBMypn6nDwXm+KfOOe/e7Z4602ZZMbQheDltFYIU
ZkIsJPFxtpjac0P/iNM9tWpRoKlpk/4k6BJGbTgc8yRRP/OsE9Bl6Cvjfm1QfgRh
d7+j9B+H4SDq/DsRB4m266M/lD7LoVhyIceLyxVDXKpIU979N2mB12q2x2km7unp
cG7mWzKp7uXIJTopgkEJciDghOIho1W20fXOgbgxnZW3nDm948XcvNjgYAZ0k9zs
WlMcY5Cs10mSC8HNRDZYTvLjJZD5lDluoMO5AqOM9hohbKdGOZxswzAn8RNA3FEg
CHmxwGl7O1VwSZkBQh7dY2uz9Gx1J+32TTFDoZIkUF0p7WDphv6cBu+tz2XVMF6C
QePaJ9rSW1qqZ7PoO+/wSjV2WvUCpp5hBJI6Db4p4lI4qKlXl2ovFCUPdDt8rvGw
sa3eDDv0gkaTZfmCpoLi9na3lZMIW90i52S7D2w6JDl5n+zevTfLwU8plWjucbKx
H4eqGiB0vMKVOcACZ++0DKU/j6ME2WBpZaksLI7gSwo6v2NEnydFnP8fRZ4xk1jy
gvEq/zIN6w5883DK71junZM/C+PO4Fa9XzYJZJXz/PnqZ16TaJ4kAmxHwt3SdL6G
4OrMVcfzoD2WpntyuO50/M8dPeXk2b3Gi9maeVuPOLWoV9VC3GmcISDhfuJf1rj4
M2u8LQF4YUQgpRu04aPxTuEqXUokK5jtdEwxzgz/gHqqT4UGm7vWsxbxjcRmeKqD
3r1Gi5Dbza/PLdYEGqjZLL4WsAKWfyvZeJ9J3a6Y6rhY7PJi3PjBBaJhymwM9qDT
SA6zet1Qm+kv5DAS4DlkwtUaU80VPp3Q2Ye+A2p84KcitjGWhdd1BZ/DrKKH0rcF
11vNyrVBx+e1fWcOIuIX/8fzjdlxG828SCWMuZcP9G7DY9c28fpcfmazGbKNgxIK
QDONHpd3GCHPrfvkMbeQfDil7jWwLyApf6VNVFQfFH40CIYivVlJYeqCap3d4Y39
YA9a8Kh8ndMxc6Sixy3Cv2mKpjH44RzFQ47zbYHt21b1zhaug81aYOF6kpBU6+O/
EcAu4W+BT5RPPseJKmNZmvaFc+dSpLdireNwu65dJbH2Nr/NaEHeFs2g8uEBh2Lw
LnjJFmjoJ6q7HGYsYdg/VuMmJcKUD/chkkAG5+nNJrYlS7dHuw2cpuias2APTOHp
WQL3YMm/5vJowA84hI6s/fjEHVH5rjn5pfBJ7QCseCSu6/ZMsDUbVDUc5kfwD9Nm
tKqMGhP57wetMxIR8KnDmKtme4HHybeJAkSrfcyd2WBX1EtnqN/4Yj6PATWiPbC4
Mlkj60OwbhvDx0cEZv8PNI133WeVLVHV4xJBaiyIPJlBOivEInFfqXDaPhKE6JC2
m4Dy2g1pGFGPJRb5pgsKrQAymSU3paTU4ABjyBH6G2buGqdJbpze1hdKDEHECRTP
6TlryZPp/Jr1t08kSUWk95SNCwllhu1UIYvTSAX0O1YUpaKFKc8AOo84pYzmNgKh
6lgMcPOtDOUX+F2p7Wbdvzh4xkJTYeYVh5w93VYKHxFWZCR9klS+LhSTWuMmALSs
58tVlFrPSUASlqB8DirMJb7uI0eHb642/QofqGhPUU6aPCgFcurnJBtCFE4lwcCL
Dwp+u61PByTebiKck3byrq30fW1gv3ilrQ5ahyotnwWGPguUiWC2Xdo8HNkC2YwG
+G7fCZqEZW6XprhBzka8pjI7EoAKu7SaD587Zo8VPnWF2zI5yVhP2Uaro0PSByHP
kFivhJGLYsiN6mShBRnY4TXtkfQYnktoJAENxIx4vr//H6swf4cY9ZVEsWh+N8xL
/avYD6fED5qpHi2sxxwtRjTFaKkm2HFM99O8lXQUv+vHlqvlzpy20x2cMJ8skUfM
+iMy0GaMVJKRFg5pRW44Fk3XJk6DDVJWmOtSSVinANSq/j7sGPjkOEymPV0JKDMq
ndLXj+zaucnrh37Ix3bztrZMJDSIdW8w05YwZqIpGkYImZ5F6xQpTckYDOTpF5a2
eXvbbERvgXpsY1c4hiqK7q2qQ9luebstvrb3aG+MTaPgSzmLsp66Ub1Exkp5qF+a
E1cCuEnC/Ag7dojrb9p7Bf7NUTrpJkbOp3tVbkOBbhkfAc9xqBzB11T/DDWaVeYF
u7Xz0i+5sPAisFoYAqbv1gTUtCosfCHshCQOwQvUGLBgP0+gHIrP+f0rmd/K/4Xi
oitS/ofByp1ubHe2gnhtJep3LjT+Dl1qNEcDc/Gzux8oliXjThGCUBbawyglR5TB
7S5qXRgR9j8Ns71xkFAbUE6MshIhGxDdgTm1rvS6S7EANR52uZB6jKlZZG/Wl+Pw
Miynz3cUN00Vx0PAxgs1ayZtbjN11e4SnsIYnoz9esMZAYHm/xpAd7V93EQbPsE+
z62J4vQgR20VisLIA4o0KGP9btSFU/csgtar4xj9l/eypHxOWZWmFqJknXeN1Ko/
r/CLuN97ypGYU/3BVY4bae6t5lThMqfx/Ra59+h4EbsplZNw+toq0y+cEeOTjO9J
25Vbk97GBy2iO+PIEWoO78erGm5HZMzaaPtawOcD+7LFzeiOrYtw+AJP+/8aODrX
nwdRL6+yv3cIlNypdsZjDUqqb2yb7wIf/B71N2tw4hU3KCf2g8L3qfOf3e5LZV02
sVhCebgSvi5j55syL9+FzzXtuI74mRgtIaHBHpsqxAbY2pWXGx4lDeXq/zWhGLMa
xCk43+QAi8BpLrR3C7QGsnqGV7E44YnMfBGxYVnNBeo23v1d0TnuoYAJy+Y5FhVb
JjnQsg3U07W7oe+uKUNJG3qZv5bJb/D2GdDEn1BqF5w4hNp1QUuYkEpjqegjsSnd
wqFsuUV4NTSYPuKlGBVLxPpXmsPYhG+hb111mg2bzZWJnj9tpIkTIuqtVDVDUjju
WzkUU+qL3+G+p2dinp6YB4k3yijgrby208R65yuzVhEzIQ8v8rvZetZyzJYOfh/y
nuHFI7S9Nq1PnuKEPCOGT1I9HrjUnpjwsSewv/k8bjvZUveCsc77mlCgQX7tBaCa
fH0eSVCDM1VIKxtdk9zkfC+1w9mp5uNEQhMYjv25R/Yst51F6Jnm8bUp/O1lQXz0
7KZbIh9l+7z/jwsSnMtzV42CYX89mfdkvcc5YtaaPV2n8pOPwm3PfHMuoJ9XfYSu
vby+6rMPCEiN/+of7OMLVD7dkuKnM+2SCYu6Dc93ZUiDLwhaDdUx4D67vA/pzTIS
CMRzNhjxjXu0Iqkj1cDkQa+x0Ru3wAjD6GZvIv4GHxUPW8q4DDHGLSK0rH5FAWfj
9pr7aZhF1VdUEArWgHmFbQ2SyLzZx7SWkn6BMfCxmFboE3ANB3a+3od7m4ZEJXx8
+pnb2pWC7/vZO7Y2f2h9DuKUNPSYgMZBvC3d2n0gcOJt6/nbSNXwYPTomIAn0c3p
O1w38T0LLTUrHg4IsUlJ3l5sCoCesm7lv8fAph2GHCVomi/SxaTm0aEmzax9IGyh
e9lii816/pTKiGFdZPpKCNAw1hdt/sSHU/0I3o0i5Gc//MxhEsFUnUfgIet3jKMs
OQkt90FhltL7KxsnUVlKv5x1TULhlA02S8jQtTuoKrIk9mjuXCfK6rDCilxAovYs
LNKRaimPe7exjgxrT2slCtlO57qvAZqgoiiRZ3Rd/D2WidDDEMZ3Ou662bMp6ZQ3
iN7O8qYB36JyhkQvAXq834v6IcBagqgOxkxmFgsPsbCeLjMwB25NlF4CiIAhVXkA
XBnFY4tbcYFWLDWb806Sg+jaRDEu2KAZVaLJVVxUceqUJmPAvBYHboJN6Q12kDa2
+FbEtLiA6wwZN/GWOvIi/jXwtrPYhZ+EjyiV9fgPHXZaT98OlWHMxZUwqeJw9kha
QXKnloxzRlZ0hDZ66X4zxgV5TvVShPxqW6BAC3nKsPE9NyXxUDPOeyJoOdYcnM3D
OMY7pPzRqIbazGElYE2/I2t01K/545HAlNuP+d5TI4IBKxXxH7kUm4iVlWcIrpxv
VxVnnGFoTDFhtJUYDdMglQhtXl8mhzZyTB3RVKicAceY2EvmJgogM7KY7dImAwnK
bgv2nAnRJkxyWNHOHpCLXK03Qh9KgvPsSLm1ZJC55xRy7fZXxu7aGPxTUrvdQb1c
Y/tVuQuTaFzTJHOE8qPUaq4/0XIYSGGN6Lqv1RZNOdIyldqy3sXaYr+H8jAJePsP
Ub5izJ7nvyvEX4rNVQedN07kV3VaxmsRiG7xbil7nDW6mx/0eCEINfHsX0M/q5dM
FewEC22XnFrS3hG5dfI8+OvfVnsRKabXE5zNi25Ij1yT3reYHR8spGbm2ZmHxRoO
8EYHJUIXdgvAWGmriY+KYQ0K6zjKwWEpXJXvAL7AOKGW3ucbwRlc3LcLgWWlTPwj
3su6oC4urbiEYl6oTBT1c+M9sIB+MPUJof3xq8yAVD/5e6QHvqI9YCWZ+YaNq+Cp
NhZ30oW6oPiQnlu4qdJsUF9uwZyLmYoihYITVqRKTWJKOzCHpgg6sKQVMrmH8agt
VDhrP5qQuXBbssP+jdOlG5cNwmWlzegc3sxRAlVIpDm2fG0IButPpCo5w/lI43O3
cEHA0zUwNFQx/bXgenVDhM28MRlk2hYIzvZFGPKeWTPR9F3rkQ6lDI794RfB2kMo
fgQOnnVbPHl71aUAR9/oBLcH3Xc0B6I6EtPirKeAClUiALCo8pmS+ba3+R/Q/1G/
O+3g5TAOMXtPE/5CI4qu4Lq2b27rWG2ea0wTZq5bmZ9hOUF3VNxjL+h6jf2puTEa
kmCF8ScCFXL1zLaK4hm186AdoxUg0CEC2ICEdc/kycAiD2gNdV2ZqDf1zmwN2pz3
0o36NdlcO/VDd5Xbd1ZSz0asynhAwVYffcIRibOI5/MKXTx13OBCsoFfs9ztaLlj
Wap+b2KgHpmjmWJoE1OPoh+4jMD5whDk9l4t4f3IzUQfzww4GS2LD6fufZtMcv59
dmu/yiaMDtMpZZ4vLCgpJO4FjkYJc+rqnsS/Ywkg8lYyyEE9rD268vJt+RqfnvyX
iU7dEcSYs9+rZsR9jTY2PeFSUiWApj0I6EU/MplpHQzBokrz+gp0y4A2rotNIVb2
KMHfyLDRoPa2/8HNEH3RQFMrjBi5gt5CCMkTJOzXPrPgw3e6GUAaLN1o6SuPE/h2
pJ25hEo9mSrUv5xeUDJWFBg1HlBGRfuvsP6jBtR/hUz1iaF2ZKjqxsspBGjCIyYH
2g/BX+bOCPjYsPqtscoK9HTKYcBkf7woaEUtuNaP5bGuSA7gQNLmLalf9lCeDXay
uZz4YR0vY2rCTK3Vr7A1FUHqkk8rZWcIRanfTIFKVG1Rid/tywKggDQrRkOiicxR
bMkuCkzI2EEK2Ja3F7QxS+k4WWAgnxpsOY3d/mwryBptSrC1Ot4va4XUCvM98EMR
PFVMLcUn7PR593XJYdUNGQRWDXCgfyFnzGPExfgHQpFbRQvNVftNiWalXqFYlpFd
3/i05oB6G2aaf9H3FWK2eenSyd8W0ZX5SOZuyKc35OInQrn4ieJEbGOJhfuSTOiC
hzwbXV6ZopwuWkCWpSAcTZapIy7UwYC5U5Ih4R1CFt+bLBpttOaKDH8zOmEDccd6
gedJshGM3uzi81GQ2XqDCd3jgjOw7fS4W1nrpTmu0RusCIE7/J6rMR0+I6tAjvby
W09v/Zjg7CjDAA/HHaiktgvjD1gJlqvFRBK6b1jb0nPkfnqQRXaFNNNYe3zAMMiR
q4Jeo04AgHwY6Ux0cU6m6kljMLEIWL/qST87GC7F0xQQ4ire+bSGhXbaV5tT/ocy
1GTvnM0PQcohs8d5HDI5vLnXXqguzqB2ba9ZT6EzfTGEaR6bZseOpO6IBptGm+o8
zfYcx2UUu9fa/e1iL2t3MYM8rzwH6gf0VRok1mV3pHeDWprznpoD9mxW1AoBHyh9
qJPTfzgQbMYQEoAe73cdKoSZ3EH8zNLhgNHNXyxvaa6j3MzDXiXoEp2w/b/TkUSP
71dU8qc0KiEcnQz0qlXI8adNn10682VfcvJR9xr1unCwbHvkEEvsQVBC6XxzGlC5
OPnWCKQDSBD1PClkxRbLA4flik0GpFeuAN6fPJdpHupXvizxwj3fxlYwWlN/tizX
AFEg1FLkqEuQYlm5l6dyIXOp9J97uiMAujAKVt05BHg27WlUPFRVlIZh9hOVxy/M
AOkoNHlGrWOIxTg3gm5qGHhl4iZ8v6YqZ8gi2PNLjQFOzdxJJBIITEpJ/nVAnT1u
NkFzJc/l69mzyI08xQ2xMCpqM5C7WTx3eCJX/TSdwbGUiiw9HZYrSTjhkF7G0PRT
zW5SfE6bHtSqR4V9a3Ar7ly+aZSuZfCvaJPy9CGuikLFgBxZ/+6ejVkN8L7zuDkE
ZXe6oPH7DApFxkQTR+GxgXef5uNO/HLnZfO2spGbw2S/8IQ55PPAaT3yYilosHFl
+Gm4g6dkSZH3c5F7mCIouvAw50GyPyauFdfzYdo489j65yDF7PmAP2PTOaf/svl3
CiXEWSkwO6O/2z6IsTyrN+VUG9aY5AwoAh+fqbIkqSQWCkqOT298oBcREttRCHNm
ztjhP8SmOYpEHWuU9rMY/0uDv0+ZEkmAFHI1upyUpRx8BNPXI+5ajGG2m/t4qFjE
TcmnzObFupJ88xc1NaSOUDiHDGdjfPdtSll4gfDSYM+i3zg6LTzZhalag2YisyAg
QH1TIGCs2FqH/zX/WKzAG7HXM4iTd5pJHLHVqmO5qoML78KtkCLHuUiitL0MtYti
7BP1kQeft8tm4jvNc1Kut3N5Cu/WJ+cTSJ5bJMIgc23zTrymcQr6iREbvAowiTci
HlNpzylcfxcnZkAEPJK1D2ZEpK7dFJhK7h+m+4ie7L1p6tNEjmXwstrDw4FpKVP9
p3p9oaTpqw7rVIqV2dDGN7Z0rbBjWidAKB0O/3qMz7CgvSuUGMoABGhsv0JrWIe3
cSUndyHG8Vq8fMhHNOfnjN1IpehRdtvtW4wPnIvLizRoi1O59P2aeI6PoEXOeCl1
wCG2Asqt28qQR7DljFALN3ZImKFzwbmAJ7wvSTqZsZ4jPLLbXGhH3MkgoqvKTsL4
auGnhxPvH96y/DvP9U/gJfKcBNOdsvmP2Cs2nsOsahJgBvouHtPUWxq14tHNCie3
AZ9n6l8MUW4stCIpPPj1ukq06qc9nhkB6/TzfGzXVYroNvVKE1W7pzPsJjdrKLJ8
mRTxNpupm8aVq85W54nSRfeBFvqa17XMleSwoez2wOTyr4vLoEqjVHa+tYLYJJOR
AtNWETvhFenK9MzNVw+PXyoZZ1ggE6Q/gcozvdCzbVf4IlPaPm6NC9S6cv9Cj/IL
plmEIKadG2DD+/XbiMNGjKDwXxm99ymJH1a2EbRUU49rPYdx6W9ju1ntQ9Xpv6e3
AJ54pWUYzwFOekb5nvWMODbNFZ5G/2qP1RzPiUC8hsO8SxUkfdhsFZY4x5D+AUsP
5w2S3Gnmc/rMPCl37JiG3mJmnuulIASKHM6gWk/xhNV4FEwgOCEKjzHiw7fusksd
DXtm0DHaLYxVQyYL8RWUBMgvVlo4CU7JGHGq25TGmrbWkxhYRc1cmWDBxtNRPiNZ
E6jSmBXI984p7Gl19xgqpHpTVFZTUMphQS3ORJAVAqjFZjm1XSNY5ZuBWFpspm/e
XnEqEgBhfocowSl99yrdkU7QZ+gWeMl2rIG3E/MO9Yf5eT6ewskKp0+TRjMqTASI
zrtf+nyVQqm1ltbnksNQVlclzJ7NC8vyO986NWMtfiiPhQwFssQj7rEvmDdzoxVV
5JO287/tM+8Dphw5gpiAy4Hg18OJYCsKwu7bd8i00B5aMNGT7rm3bpllIHt3DQ/P
/BV9AXinO6H5TN5I/LPGocyTmxnIjg7l5lo3WkzU5FGCw8hvnJVwfWDiKvDBVONS
sPrH19RFmn7mKsf6ZJCbRbwGOQKTpDy8gohbCItP7uOj6MyGdISDT4Jd4o2kKHs3
7ZKJmU7DBDzcZULc3Rb1gwhfcE1RTGm1osuQad3tcTMrGVscuEFP4lv65Vezuatj
RVLLGrX+P8dvCXmyyQ7RUTKtPTnfyoMagPJzmbVHfDFd3+GNfNzxP3KGwr73wAJ0
Z3vrQYehs0uI7QuL+YhsKJ3EpFOOMDLXu0AfFlHHITVZmwnPVNVzKsm8ZxAeBlf3
oE9B8lbQouLImIGWSdyb66OtS99nuG9eQDamWwPtsNRB0b+8UyYy3QZnsccR44uT
U7QlO2VadifasV5wyRRLV2ncke2KDdDH2qJDS24VDiGnLeJfKoiHRA/iK/ZdWbXR
ctsgEjKCfUHAJDIpMKYY+Eew4VViiglVx55MpZTi9amrilIi03zPXsE1FTxtGLBk
EOmanUzi94qeAgLbHvagQt4KAKrh30vn7D72Bs536xGnETRSiSBkzwptCby3Qw1T
YNMrYCyuGQU8ZMawpUMG/jN0vx2fAJtKS7D3hxZQu2oGPB8MllF3cCLqnSguf7Kj
AXo63FJxTyB/FJbsgQVdWDZfx5v2njyQ82uGqd6y8Q5eQEv227L9QkMPlS2q/wJ6
v0JWvuy0MU0+QlU2xnKht2+jISqSVXOahE8nsADWBSeRm8iJEJCltPN5Eb524K92
D6vBg6ROVaNNcolMlwkiHeaFA9+6P6RLKYfLLxcUqdzMgSeDl/jRN8qyNilW4LlL
lCjh/+GQ5bvoq7laielnLDugpJziWqWAmH73LcMCj+3oZCjCtwP8nlKnwPTdL5zu
D3FxJbAOFXbhxa2wIGKtqQ9zoLk2qRz6QwXpQ58RbMJpW0Z14YuOg1K0JODvJ1Z9
I9Uax26zQ/lCU5UtgRbqdFWcEd2neOiw38R+Y2/4wqSbEyuZJB9J8fMSbXBP7htr
BPZXKnClUkXTyZpOuXNsb7GWvyXT9O0+ucL6YVXmLithKJWl4ZJoYAJ/YIEeuEir
0G133Vg+XdpwCRklik9vBIiYXzed20664eXP5Xx9Ve6y0Vo9Jzcj8DxfeMOKmDYK
2BPhbOH7kEn5OKhlh1fIExWVT5F1qeUz8jXHIrlykzLbPk7I4XlFIN9uA19sW68M
1m2osQefs9VWKqYeRQH5eR3mNHKszdU+HbY2L5CDimnoy75oBrIq0W7idSE8ifBs
NWMKgxhqSoPfDWaTY/cpxrXXbiIa7maMGJsFgMMGivHQyHsFO2Prnnl8vKKJoHB5
R0tPpDEIBO3G2Fh34bTwOWgXDCwI7tldvYFGK81NSVnXYbzFG7XVAPn/hq4uBXsJ
x51TAfYK0cV2BSHc/93ELkaG/XiomGWVhG9CHxJ1OkB6eOIX9jYjzIIaDRfNNIhk
1OsczYzcQLFrCixrgb5CM0zkkgJZehSx5MyafVx7uoP22NSTgGAavxHMg/LihhX7
+Wk2A4H6L/H/sgow20f9BDCCMpsgBYsVKOFxAgYR6ekxhejkBWCB1OyyUOSqWDAb
mkem4qTb0cslLyLcw7WnojEJmwd/JkV7riAhv83g+njydKyPVTjkvsWLPaiywQsh
NNH9sirNa67WhS6vN/iTHOYAi5N6sK8DS6vlnIscQp53u24OWM1z+aHu6VSiu333
ilAltN45GDk72+saDdQpEYpMMFLgvtSTuGofvnSvpTZkWfeNs1d/zsOIZzIv2qGm
7Y7L4nd+tYmN+e7LoDIdg5TkrQEgFrr9gvnib0YMuI62ELTEZxn9gUUf9hI7HALz
J2y3NX0iWL7vLazr5NIMvZ7IX2ePwtB9mmz+nX8ARpE8dy0HBqX5OEvLxJIho0Kq
+5TSpOilFZJjPxBjFJgoNGNN/4Ob0d9qVPF2UXcMBzjNdQsDuehZVtD51PNfBqzj
wUhdlh63E+a1XmrMhqrcKU0/e0WYaI50DXaJ2Dji2C0HZci4gnsPCLC72wLFiHn4
oIl2vYRJB7Cbh/KjOoLeGvtCddx4J8wRMslITKCPqNJV3jEyLA9x+QwhvT4gs960
XQEV+DCgfh5YSTRDrizmarkNtisguF/bPs6opDDVx5HFepnCr2r5zIecqox1O9qv
ojVM9xLNLTNdrTVcYiX3a7P+ufu3PxpHtWMT4rrj21IE58EH0tsvpgEm4ukjrFay
qklTQR2isU1Kz53z1EmrUNaPc70f1a3S4S/XMjIfYY3/1U3JTAxOwLRR1w1+ok+C
IgX8q0IUEZEVWswL4k6g6uIsOCC4QZhMWI2HqDW5vfGHYcVZkaOBi68BvFppqMea
Ol4C8XGLfENZkIaPcW3IYZ7/QlbemXiJfCyzNiCC7ptd9hE8i+lL7ZF7uxCzMH7M
ARd0ZsK7LM7SKVP4F6YiL80GyFCYu4dTZCkV4M43xyqia0gs2ef/JpTMNDhWWqjL
6SiNJQ7z3glJ8F1MG5rQOYmHs89W8e/wq9M7+uaj7UHK/HpaajUyTq85K68VnPqd
pnAck6SlhdvuqBqvAuzciqEhSk+fQNyMJKpERCCQsH44RarUbCib93BMQo65dQ6m
hJDTk/LQyG1YG89Mrwg8pX9id+D6zhhfHfy8IFEsCFoK3rJy7ZklWfJqzoGhymlp
xQ0SvwaFP4w49TIgB688I5H9JtqhhXd1AbNpyMXdWonpShGWl7z7z9cwlbKKuV83
2pHikhYukAdclzbJgDAXVX+ZOmsoT9zaE/iflH99IMdK3IQQKvpIpDPyWqdZxwGO
BSqcOF1ZEte7BfQsR9KY+7mx2cNAvxK3/Tn+fv4UqCEzWLm/QY11tflu4vM/ipgL
z7vzQ7xxF5qnoKgEAl5tcAc5HzddU+zpGIlTwr+QVMeVSiWwOGw73FAccOAiX7LV
UvNMZzrONjsCfDW5UYPM+ldlnW+NI6I30mquE+kl/a1ZsKXAh4Y43fm7fWZ/K2b7
NkYt3JCeqboFKrc+pW1w6pOylGD7hnfPZp6KVaxYsdymWPpYzTaVu+1ly9n1nhz5
keHMT2zwrbKVfgUX3ECYUMGClqn+taXLwCvg7+MGmyyKtZ7RbeG787rMvYtzPYp4
aIrt6iEDDZeVUM5yQYTpzC9oGLqnFvhLftlXXz54wHaEpQSrj3cfWU0MxLMDHLVT
KKEc6KhvBBJLgV445hBL+FEVDjl0PQifPb2mjun82N0ZyAEJE1OCSxwooonlF5i4
U0o1u0J8ufW2GA+jCxGtttkgtDhTgOeYs2fi1cKDBKkTOxDQl3ueapWxJhmnxwES
8+lnDTtdwsTIYtqO1/x3hdl3Q6hBEanCnHXNxaOjYIJ0RStJpObd2bL/MukqsYMK
GGGCJ7EVVhmO8uEpyECUchskrlxos785cUfxCOff+D1jcOEfSS275+977YyRqFLU
6lR0qLZhGvByu2GRvwD/W/ojcpqFVSXtf8ZbWNiQUSxjXQtFr8qyOduLde0soDNQ
cjFmiLP34kqawgoDWuQq7yBay/GJMv9jMfqcUTYP6VD+ztD3Mip4xQXqDRkPAwTT
xNVb87TMf6Ggpqn1geTVF3jlhcyPibg4qQp/PdV/mfBQLYe/uty0BcsxypBVyBRR
Ye9wKMVcwxaLrbiwICMLqYxGTufAzfZVWcWVrWehb2U44tip9DOG94xNt7QF5biH
GnqOKKw/5fMJIQ0OSaTV4A9UQNwdOalfG0QKVlrq77w9fM5dmpknOYbKoc2fHoii
cP4yLel2v08gjreaeibLbQvmmqdf1do1bbhblQQDDM93cXc0gGQuCQgEwHlrUyFR
2aXMuF0T7ZuzF0/wcw4zrqBNfTxt2dtf16HII2vArU1NhKFf2ADyFSTNSBInMrLg
CEVdT6etX8KICOxtXCitqw2n0l9cG59QwiPGUAktcWcuaj1xx1UfEmZ6+ldD7fM2
JrXj76bqpwyYCCHFfOARRY4W/81ynMMdWiLW0DXT0egz/2DZAZIUL3tcrvgpILgN
vj7xgP4hlaQ51b59JDdDIQaqTCO8sbKTzvv8r3Iu1D9is8IW1o3501kVdKoMIyf2
9rl1Kpb63ZoKcyTpa3L2IcvWdYJxgQqcAeTAa6MwqCzpbIJEgCyhQ11KRfnDCAz6
djgGUhT2ZnU7MBYHAy7OXe/v7Dm7JtCieMIZ4vGXeLtruCryjPKPDjv1p0+b6kR4
Hc0ELJkgGvaG7XWm+RU9np58g3C1v+H9eJQIp1qYi9i9KBzE2HWlhdmbz9ZS67Vj
0vcs2C4mVtDD1XhjBlJfMkbkOqiVKwNq/MrjIsq9h8cwIyrW2m5qduDDALf4/dC+
K7soqUijyKBKWYh6wI3Ot17y82FFtkbQyGtafd7IL0bP8jNBHaIFT/70KMt+WAXU
j3OswVMireBnWQCsMxxNQlTyfMbkzRSIAT/NQXqTyIEwNDmaKqBKvbOwJdFBLU10
YoOpI8HiQfiaKs5IaX5VbsDK4xjUSdTtENb3aYhAwjU1QjQv/h2HMCZ5XKVHAObb
XdXLTvPuUNFCINdW76monLwUA4ZzCyKLJqzAqCVULSkkdIYSs2QlSZ9t2uZEIFtH
+SyDN7zNG0K0Udz3BF8+XjSUt/L7440XhHt4WbvJENr4ybyLhKHm4E/mBQ9OpKfY
bfWStF3t5b53eq8uZzzKySJQqkwC/6Vl/FVTV34hHYclsLaDVI8hDvDntKm5Y3zl
siRCjHb/31zioYF4EHo/pVJmpeokl+h4ZhqakICJ8ex2Dxi6pabZ/JYWWhENBGMO
3ce8vQn29ITc9XKvWIKfZTzPChf93xJmhcr2GY3vUYftijIBlzZ2MvYqGCG/Gm0r
YEMadznpvcqge97FprvafhRKeYWcRY0IrQ4fba22F8QuQ8hUi/hFZa23V2PCY2ej
tnQu/T7bfRzhblvxwsyS94Vf+PW/T5XIlp155vGjyq60etgk5vJDkXNlWd0cwz6N
BB+G2sbySZF2hAdOkXFgLJk/UDQQxbgTErzJXAeNYS7+QczGTBbJC1q33+IPa6ox
Yza+M/bpGdWuyPXwaiNQNL7t3kdtZqeiA9hbV5/DEGYZSu4pdXlDY4IWFn41/Rgn
4mFyFZAD4shajIdeFd09eHg07S6dqt2z/I3BvLyBjqWPh0f+nE/19e4JOPSSdMP4
pAanZeBgzHgAiOiK/TUeWOSGHd8s2OFttb0zFDJbQLrNvaqWHzydvkjRWwPXnFwT
j5aCCZMe6jXMlpACYj0VcNNR1Sycxi7r7f/z4V4YZWdzv5v94y/Hey+12JYyIMpr
MgUxXVyMbCFDtcwFkvK9h2neUgNy6jMI0eV5tuJa253XBUNLT9uinY6z9SlYxG9w
Gvw0pGPVinZGS3Kvacb/IVQK/NfHgr+647vbsjT8ufGRbBtwJStQsK2oSuGR0Jdz
LHTa5mQ7xRcgoRvh0y39bH/2dQHgzUFcjQw1bz8x0U7GROMTJjdCnyARMlQv6Ov8
dFcbN/ucJBO9Ib8wtNtSPbN5RgDfO1OwCNLU2zPsvP3ate+tFB8nH3XCCuepA+fE
qKBly5lAidut0EdNkM7KZaGQUQlt4EHzxan3rNlCM5O7oKMJEvknGJHV+xT22xon
dXtcjwVEHq7mt+1jHSRY+wsReRriZX/t78iT9GFe2TiH40EDES7DyvfhjENtB/NG
ozOZWxrGx6uV36kDzAqhi3H6AIUtIX9omW0HAg/hVuFNFPZpLGqZ5/SDLJabTwJx
as/CHQm3w/YW2FOIyCeYiB2/Pzj+14IXgU7JbcyraXixibsb42dhKvbhVPn/Zvtm
SeEEYOdfsA93dbLr7k9MhepmcVh8E7z0ZeDbC8BImnO8/Kx9Wq5qhc9IcuXmR9e0
ZXCm6U1Lx7kXIpA2NPOhCYmr1x6lEeifOolTtKhCnYF4N7t26ga3V0NpQQrTl6KC
n0GMeK64A13W+Mw4Qiw7yBWwq0t/W2pLujt078Bfd8PsdHUu7Q8SXOQqiEgfvqkD
fTLL89QfhxarzgoqULBqKD9DQh5pUNyOC/MniGU85H1Vj5y+1yMvIifUWNR9+bJc
WpEIQQIKPdvC8fK0yWC4VbE5RT4fKnHiCU4ro57upGFauZLrEfg4GrhEXXh4m1Id
84zfeu/+FWjGYGyTqNwd0CLzs/oRNqms+OuY2vyfLpWWJjvUpxZsNxeukQGnMJTA
wCjpEjHKs35qETDRzuyiS/kaO4pqa6/K1hq0KHHLXro981kvLL8mcssYV2Nj4jcZ
UcsQ4kS+1w8tikJABmrBbKcXJUrZm0LkvTe8JGW/Emq0FoQNsn4HyLmpNNPtuWZu
caqs2oFp6rG6qhNNqW3u/gaEQ5/jEyinIyK8P8IA1rxlM/eVo/2U7Wejtgj9txMX
rY0Zh+lxAbEsHXO5UmSZj8DDhGBNTOBiOJ1mHiTFZyaHgFA1VQ59qEU1/VBdVWoh
uOXeYV7vbemXeYrtz7mloK5F6VvOkHLjz5T9odkrDvYwJFHWWdEhH2AO1owZNqhT
kW0MBgCYQRNB6eIgU7SMMAWshBVn/qlPNNUcDF2DenL52pUvkdRgoPsxgCw12QSj
04cDh7Lh6mxUDS2iLYIrAD3dGTNYEjey+T3syGq7v9tne+CGKSNsNosQT4H9a5Jz
/e816g4V9fk/DWm+RdfTV/d5nQKv1LFm0DtK+83UZyTIl2Uo69YFbUEXOaW3PQdk
AVRVxxpmHDfSfTNEPB7rr8SsXcfsJwmRfbKpfltA2LKbX3HPgmHRwPiLem9/jNGs
rlQgke5BuBPXqaYKIxlYK8EY5Cbcsip8QV+xakmrHCmS21+auuzbIDJFAQafWAf2
aBVv3HXB6RJXW8FcEDp7hw+kt9E1g5xMdxMD1P/snQWY8mcwECWS6/78qke7RCjD
QZv+nHFSyM99tzfdg9L+41rw31aqx9a3n0TU0V3RlT8dJOV/IdHX0GvPYKDwDgL9
YWFQqoo+PBYG89BQL2ey3MCT70wdueX7hRxEE4fM+YYkEwb4qJWtf2F+PnjdmM8q
B7A+6iXaXvKWqQyU7+MLCm2TnizrFYBjEQfVGmxt4FT/+YA13PN5Ytw8M8LI0gu9
8CxXEG5Mw9ZkKDZrmH66vfaX92O0q/ZhTxX+Ssc16/madj99uec+iQpqEPIz4OL8
CvPkP6Rcs7QVMVeQiWobUPdOgQbMlm4y5IYTQ29t/OQp3/9uzFEF05rTRxa5r0j5
xRniW9ciLmrjDH/cR5aohcmV27Ij9sUSNI8HWThKWgNwdrANnmeVaRBxW7EMkhtt
uQ1DZlKZa3iokfWX0KjIBNeC1HcU8DJXSETTmMhvoUfceM7h4qruS9OWUVy6cjk+
j5HzlAtCv5EfywggLw3GwHImQFD8Lzf3gToEVMKuzzu6pRAtgGxFc0EQWn22gl6t
3BQFT79IA+zGPGgi+gU8Wlz7j0dqduZtjXiHCg7pNgJZG2n9dwe/cBsJpZ2MbKBh
1I8VXrbZp8uJz20GhjriZP28ZD4X5JifmEfq2ZXkMiQFTh8keE3Mxlf9yUt7d1jI
yjFMV2tIE6z/EN5yxeQOhRPZJg/JOsdNvo1jdBtQZyAtn9HeM7osZwj97w1PAmLe
lG8i2Ik/DPXT0LkKuG81QBrtHuSuV5lxn63g//7K3rxLd7y63rbJEuE6OdGVM61L
AJ5UU4wxA7Zn1ZOzvSZMFykxfV+SODA098mQEeEhZ0DoMkGhxb+GpE1M4P8As9ed
0Htcv5wk+mIuDbemyakCZmuM0FF1Pj9jwoqDmUJD6fYET1B7ZhA78OMD4ZNTM4nP
bThUCuYrKlGoc6mwkCuc2Zs/nlZKuHwt6ZQ5xjE1cfY/+Uh75xycANAvpBbPniJo
N/m1vhWLK0/o6+0OqEHY+ca6qwFzjAoCkbVCEF9YPOu/ZHnGYQMC8FsGMFCJ+cRL
5pgHIw/Cj3jkyfTtNf0jGLNXFz/jdLcj97UTJJ4GuiwniyezZ8na7uahXwEWudho
jj3S5YLjS89fFWAHJvbJqcjJAVEJTFRzAgNfRroE1jAdIyDK0MHAFZzExOuseisO
qqVHl5jgd/X+bcS/VyN8p4mDqblgqmsMiksGaI93vBVOS48xi1/tjq3z3rNtnZ+b
7Yg/itOQKtuHilJZA9QtFUr9nKZKT4hu+YyKyheqdTV2F6+A9gZ7P4gSWUyf0qnD
T9TA6haWp/2iknJ59hKglJaLaDAEBPE7i0Ywiv5AnpBHGWeOaqQjn5BRCiqv+vs1
NWhL2k++lMgSGufdrz7DAhn0tlmEYaJT73xmb1DB5W6OWqRgLNGcdVJfgV9iYNwd
h9iGAowrU+mhXdGX0tghsyWnjlAtyNEYJtLKnafU1TiOAD4liygeT7W3hs8lNWr3
Nh/yMUsnazo27DqFIa++Df2jUBCYXJ4MFKTCO6/DclZTNRicATvHqZd3p26WYitR
mo6VNdO18xtDipYScMi/seI27MZPbAShTaE6KSwwu3SVK7WP7fVDOySD+cGf3g8V
o6fi8bGHzJTk4AVitlV8NRtYqgfFszYHCpeFFN/Q70DJKi/mDtn9d5QSS5UHpFfI
i6+ici4GjPSM+B88ADKLgcbb7Jhk0gDfi1rg+8dKbfcZh/GFM2QKjj60g9UkCowZ
22MpUlahL4lrgA49VBurlR2yEL6TcCwNeunGFLvS6Z1kqswb1wSYXCS4pREzA29g
vKQIUD8AIpx7qbAY/dcy2TfAFmdPFndZA3vctkLOshghFocVAe5zxHccPJ1fz7Xi
s9vCxzJpY0XwT2dslyZIVvYM7UzrF75+5FldBK6OsHttMby4pZT+XZhWLA/Pwt6G
qIsiEGnI1W90FmRRdYNMoBWMKkGbS94wT9FjM4aGIRr/r6J+VFVSwhzM9I5H9BhB
aC33pEfZw2CGQEInJdN3CGYnd/4Dk/Gtk9rXEm7Y4Io4iUkrGlSvqngz6mvJZl6y
2GhQh5lwdcGgxh/JYtkRG3EkVdqwIxv3trPgs9jlo9by00DhjSQHuF/sdije+3W7
ZKxN/pDSLx1+bfXJYUun/fUSM9dgGda+MEyJVZZruZK68L4PBsyUPxNYuaUmU1Vq
NVpXW+pNXqaUctY/DixVtKEVuynhsdnridemRJ2/ro5tl2sZ+KzCOrGZiiRSfSdk
xQMMRzte9P0ovRakgbIDhS3lIs9w05F08p4v9eZhiWVvi9At3alsIXKsIy55GfYA
9xu5XuSFKEkxuVIDPhjowZerSpaMqUNM8U1BRImtGg20qcD+F0D3Kqp7xCGWLkql
Xla3DVtzjFhys9HVGBAQCkxpym2ft0G0OGUKxbPc3fnXr1dkvJtKiAnuYuCSXhk+
nbQVtKwJlQIWiLFMe51TOd4uvYTp5gxE13gljrSE0HAPf/hX+iJzrcuCHMWGeoQp
rNa80n+5o5asATJWjDtkHfvgScCR51C24q/ZnjSyHbPlhNEeFMZ4pBos71/YHqIi
XFtjpyZJOEVIF5opMr6hyzZ1cZv7OhsW/FX1xQLgL6ifYO4ZXJauOJcDtaePgFKT
7ZvW71pxX1iEamsl/DecMUAQuxbrsT0o84FgNnXUljZ0ZvzUiUef4BPZLRp8mVL7
q4gER0fxyciulGhqplKEmHUpWORuhPTdEad9OoHuDubErl56eMJqU6vBz2KeWPV7
mRZ9OVg0/mCE63/nZELQ5Go5Ml3w4oJFfbQnEmzk61LPIBsCzEYvM6YbY6H7iy2C
AcVgYC9GnxGOFL8yKnU831oZLePZR/QPwzUM3KFAI5M44Mp6uX8iGx1UBYYKWfxT
DxzIRHie5Hp6W4fWIfhLANgvnN9TYnBRqtyR+FXcQChQNsmtHK2ZPpIELR9HDOSW
0G8nm/KNpDlXx+qHp2uAL6caryMSUkeT72y/yQpdKubFSZm0TWoQYFLnj+P9FQLt
VuvkRC4e95jkDxDaftmXuA+L62t+Cja/a7Dt7JQ0ylqiWr/yGhGOBD4BodtGHEHY
CbBiPnWHvTIpsBDTzz7F7r3szf9m2FKRYgCtUreUyDihuVgE11nRYcxsF3ZL0Svf
PlIufQNxp2CjYkbHJ1r5VTQ2y9pEDz2cWkQsGKyQ5yGnRmKn/mWWBHerHxIXSloi
2lj+t/HU3YYhIYlwjI6RNh+Oh8E6vZ/lPMpbrB27xqgVPuEiJl1Mhc0rF/RBi1Sa
dHRMijhkuPPcb/plSiyYVCxIKbmn+ymUe3D23xafQ5y+CkP8P2xgLs/0o6Wa/mlG
MSSy8yLUxKjptx9gO8XiahpBWYl+J4/uUb617yJPseI4w8Q/f9JDEYCSL0IiJ1s1
VBEwOJIwCrd5ech6LToh0/1QSYez0j/fd7E832LKXdVTAQ03sS7IX/6lxoh0AS+n
YPEhrDnrXsImebTFvscOTYJhncwKJ+p6ZjSQBWLiVNTOHEu1F+IPUj6yr6LITA6E
lUUjfPJEklJ6M2OhFzKLeo10SL780q15CU6u8yjdyZ+5cMJz+FEAafg9Uojw44yW
q5me1cVLDwzALnusdY29NTZsHTHByTbcGJe4mwQ57V5/yvjUaYZbOOoFJuF5NwiG
eTdHXe+fkYnuKeF3SIjpw47Abjd1s3nbZ4AEqsrQPvUJ0zt+MU4n6Vv0CimDqAGj
Th8gUPfalEyFzEbENWNgIsbZM/JvXOfGhz5CxGrOiNNBR8AHUurxHTsr9BFQg6p3
NwLqdRPNKEQ7JEwdxVtxL0DMXba6qWRSn0W2N3EBcwvYvRn0t3GGyZ+tdiyw+mO5
8z4NL7vyBh8PV3yX39phEgPnOyu34aAtpBAuATv8E+KONbyB25SeDme/ETNLJ1uJ
/wKDkhz2JJY+y/aTJgjvuM2bzVjPM0K7uj8apxQV3+18vUVLieG4/XuJF/5mo67A
mkY02MKJuWLU5CfzfHIL9iu3V3wP7Cne5fEoSZTwF6c+J34KG5+zApXyATm3Y7ZN
wh7oxmrG/Mq30AQbOUxcoFkSqGLrPkcDQ6r35DKGUxDv/2eeIjWO3aMOKTwpm2a+
G+t0zFq79SwGbfcsB+hIwEhbmXnCIrB6IB5dce1iG5W+7SigLlelFkTYla4PS8nn
ZmnG96sYPvYc5uTxwRQQM4XFHzmge9l/PiFqExVrGWAPtQAbgnBoTkdnD9+65q9s
7kyjBgKw0DBQArQm/MrJbDGbW4Y+9/5nzxVmSJRfM6tyGWpyOA/UAbLMhQ2WEqK3
iooz6jaXuHhRSfO6BCP+0iOE9xZtPc0TNW++wgRWTxbIJy+B8NEF2ZzwCRG6udsd
IlnstC7Dx13Mj1wTNvujh1/19/Qk+wlSoR5chntYtv0XMXsjOjAeVq99X2OsBLJ4
79hEn2N1sgwva5UQLRpc0MG6K2c5LotJCJ+DZE5LsBlwLKPr+1dP2OZOoZsJhNoU
YLorAJ4iO4ngd2NfBYCphFIEU2V8z87/+cZ7ZO0NOy13igD/r2ES2WfTqacVM79Q
7Uw5C+A2OVx/fgvl2z9GBgp5soFzJti8ON5Rmc9hg1pLivYWm5g34xcfnUyLUNzu
6GPK6H9WD7fKcs84TtDQK7NOYF0TKJJHejgSogvye9gsM5o+3tfISVi/nDybpb9G
cbgy5mSCAZ2LizbjiPghoirHJvBRF/jl2pSuPnyK1AywInhQogUJM4z4yXqhtC3L
togaPhzQcmS8K5eiXnb4ioz/CP/EbiBnra9tx3I1qjJWyF2II7iPglonAX4j7GOH
BrP6iyVRTcrm+EHh6bkWcaUlVWwTLKuSiEcnI0Vms9+2imf6SWHXdk9NSxv7vv6h
Kv07RzNjGP6VJpLKpS4KoZqvyZOydjWGkYP7cOrSuH950vlK65/2vtDpzhrU/mOZ
Dlvj2vqzHQKu29SSWRblJu+BWfQvV5+k2zYONAE+Pq7kLXcPdGGsbQptaTpAcsfz
AhbsPYjfV6DPxqGG1y1fq4SgR+u7uKwpAWoIjBvjM/yfBHz9lXsArSJruYFMPt99
vAsey+DZodAR36c4VVRtfWqZ8Nl7kBLK4/xnfKU3q0PAh/N9zpvPHSnc0svtKI8G
uRsJpQJIw+5cFVisCTpWwA+FOWfuGWkoabm8dN7r13O4aENpeZrmcRNCFwCN0Tnu
uY0VO4Xb44tREou9YUnrn0IpNf6FiIYvvZQLxXSVikSxU5aaeoD1sngMUVCC/hb1
cbINcDcInRrcaYCUofiAeawXV7jMUQEI80ROnebqgFzY/j8RimPjgpb6hkhR+DwG
MVZYV/sJOLuzD8r1tDedUlsuf7ItjbhzLIikquGSXWGe8R7K5eQFYd83mBGGFiRQ
mmAF/LvSmJ9UAKjXXWThGqpnpwvjdXxs7OvlQMRcmIPkn7uxUxjiXaLDhbXrvgmD
KWfhUFjAfSzBf407o1274tpqdtZCOcqb6FcbIY26dTBEoku1bFlhBsGz/jQXDGBR
Dbdek6lENSa1dsNIeHAuukA+PkLFWTgeajLuGXt7QE9US62jy5DNe7MDW7XSpGzZ
SWRRkAq5cvvVTEUUNkUqCKvV8JBzZxUMSDXhJ3+ZHhrjh3SIddMCoZ/LPuuO067Q
cAr9K/bnKXzg3OuXfi9uGe44rS5247oPLgMvujNFGXrV4ygR9cg2UaR3OSJvuStR
hwT7p15bOZAdOpdUQCx51oYhjPCr8ZyUSOw1GEUv+iQH3vuAbOWielG37AYILcSP
ly2ecTZl6jqPANS14VxPxKBoWue5u+WBGdx3+R79fkP8+9tBXGJeJvToFmc7ubk+
sLqOOMSJFTZKiIybKqmwjIAp81j7HFJCH5WJaYs/WZbkFlvKmS5WB6zzW6eKO/Hq
2hZLRCuEWa0lj4paB5G0s+VeEf70Egmm2qDeObHLk2uW878K8u+Dt91rkceG4se8
3eOy9lij6NJvTSMXT3FRK1NU4U9zH2cV/G12vt/uJ3wZP3BI7vZY5BesGeX3FVEg
lZ1lq4XnEgvlEnBY1VQh0b1kC1I528R/q7KwesdtT3ZUguvCYY/GImNGNwWDkrB0
y+Qn/cLfDj4cWclHDgrSzrSqtu9uFzvE38zHZcmbRdyFa9NCJoZNwR2z+185/KxG
fww2m2Ldu03N9BETgnVdsGjzsz/FrlqklcRJLWp+fRQPIs0qLXSg0Lv8pZLsR0xK
QejeeEp1iZBs1sUqBe1VNvN+B4barB9+PQnGbmXpvcbuHdMAaqw5hmpQC9921Hhb
Ypnv8SiRFONc458D1gYgMG116vhXdG/hSORqOjwT3bltgrThBnmOsell3ALZv0wu
07Sv9yYJcLSHYC5qQkR+Q2lQmL1lhog+SNnYq76orRPhdwbl58/+uLfG8R+4+6Qe
pHHOzMsHX22IQ19keefh6pyjPcrL5qvA1AiyERe5zPnaCsrJ09p0XinMD38e8K+D
IxJCMBNdVh89Kf9LC8x1NS2fDbY6sG6nAcuONipJX7LJ8zWeEMb59A3RFPhDDAvM
nUW3A0VCtJUrsEEr71E75IbOW8ti49wHq58CIAko41nfQHZH5uINYEM4oh+5cR25
v+u+LZOgihsESmJAdjBn/sNwWIScXDhSsDuSDT0rDMU2R1fSidACqE2sMqlbad0a
FXG4GTkJufVGCzjX1ijO6wQPUOyDlMCK3Ai+bAt85lf6fkM6rgTH+3tXsew9cD7R
2WiBkDT0Slvp25jlIC/du7LwNC+owNMAYERNJvmMqRmvAxS/tVQGSU190POPwh50
iDlxg+lpjhhEobxKVSPZLC3eNrClukTqFqbe8VOycfXztIYEyen1W6ysTZPb3PJu
+TrpBs5Ra4eV1EXuPEZDa6esxcMSjdjRS3oPUK9M+lTs0lgFcmVzVdQjYdkdvNcG
jX1ak+Aebpw8WX2elpxv8Zcr6qqxGWiBxkbtggpS1b+ikHQ0l0j4VDfG/WWb7+St
4HxOKr6LXmJaIUnx4LckNz6pO+av1a7AFcztWAQwtdOi2dXNAuk/7BdT+gbOWTYe
AC2iIhyb/J6P7/N3/hzhbiOaP94jA47ITroWHAmvsHzqmgwzVyy+s1ECnWP76oUz
Qsc1V8tuGdIYG3srM1GFn+Yu7ZXwRaC0VDBuJmbplTvVkHKj3OEf4eZTiom16A6w
Ut7aVvgTdBPZKW6mA60xuzGzB5YKwbVDQ5aFwx5+3o3zieMcEI6TqFwuW6SGcKNs
o8u4h1pNtEiqCs1ZUUMtI0dzhfO5E/SCKvCkDGWZ6M8k8XqGpSLXLgxoCxxHmJuR
o5q+eVHqfYe28o8YVuZAXPZ+oOPrHzJ7XstoltbmRAYtHRnffcn9jHeOIRwG3nfu
usQeNVEReDp38RcBUAm1DM0sDZGQiivxxtKz/TZVUnu0lbPxwBOg5N6/6way20o/
4bOQhREl8RNYsDZcyIOuylAN5HTicU9XoE3JwK85WIe6PiW8Bf3iTPCPniVwQBJx
ScbRULPJPGre+cL8itrtIvNTcr1I2pwQkRbrQau3RFuGy9bKs4GAKQF1muRjLD4R
eHy1D3UPjtoXHXBzxgZesaAaNSzOQHRmH+GVfXIRMWdOmsQAsgGKCkj1YmGJ0G1P
7iW3B2HahFDemhV8uTQEp1Hx73XDs8/R2HjRLrl2rIklbyjc/K3hi2F4a1vbAkpQ
y+WK46wqrbIiHMgVl4zW5igRKUJywEaDj/p7z++fmYpeY31/PthuWOc37QCYbgUw
y9KxoSom3E/Xi9mUDTZx1WAqMPgrC9t2oPQcXrzedi2TWBuZFV+5u/YNt7bSbuab
logjMwBnURm04phhgXf5yzU9ELNbnKstCRl4AZ7s7mG5LsegAMpiQfO2bqWktHx+
TSkXyZ+koeD3lhMNQTAmH6xzWCLiu40fHw+9LfGRrF1w7e+/vmbamxzP9VvAFIOF
dOizaUGskwLncxfGUuy/cM0X/ARAgE3rMs7sQqvA+KMfc9pRvSrwiFvJ1hfjAquC
2Djw3h3f3xyS8pZtVz57Xet59zMZT7GvLdOyN84LCiYXiSN5Cb3Unh/mV623vwhi
XkXAzZt1pck/vDXQ0Idyau+s6fI+6Tpe0FKfVnHBfIr5nwHrdJkgZmf4TgNNu90y
DgKaTQKlH5gRfTiEM28uIhXX/WgmXU8e2EZQdYZcA1QnR7p7toEV7jAchqnPVNcQ
TB4cZgMTBzZUE4qn+gwFSD11/+cIphXtd6ayIOLXhG28r79mKny0vNaIquMU6+r5
jwqe2QG7+GO7HTC7s1UUaZkWJhv8ZGSg4ekxBmH73nhZW1cbW0vg5kfLq7LHAuz5
RpTWgMQGIyb33cHDoIdpT1G3/F9ADglIVd4eDq29oqyVEyGGzshK24H854PoDIQ0
Hd3R7kxK4VaFw4g6iakL2Y62qLWPGcWts1MXjZD0leVpT52Ux+g6P5YyxkwQ0GdY
NwrQh0o0hv6YD/gNtS/yfeo+lQRa8PWatSRmRWvZ0Qbi9JuJoNbCRw7eaWOmNkk8
mknFRxqvfeLVjpw1aguj6DvmkeXbpHQ6GfLkdeMmb2aagw9YgLcppGql7QuCjArC
C5dJkpDtwRHv9XiGbWIiMVLoGTcyJJdRlChu5k8zrLOoOKkf+zalj0uce//A5G34
jf/RAQXsRRRmiaruO07LN72PY31lTPHKSkIKaiKmJrjnz6Jydui92xJawhm6UOnV
wnbQdmPhw4eTjheMqA5gkbxwqx0+o58C0XHDJV5EgJkOUm69fg1e0rtPvky3QEbE
ChlaklxJD1Jx7lS2mtI/1Pl3dyvdtZ6H85YgUkU4S9EQORi8bLAxFZYQIGFzxm8+
8DAk05CRqmMRXYb6zHdlIZPwzIIN+VhS0kajWRyoiwRCNtYb3rzatr9BxdW3XnEv
ObnJutPS2IqO5SowAqSglUbWLewRINT7hZRXLl7x+OzQuX2fgUCEmlY4/rr+9EHP
2JzXgK6fYh4RpV3m4APVcaZAM28yS81jA+dX358C1Cg0TnuOQuEG+fNZvD0AAPpJ
DbgBswkz5tzDT4cQnN2lWyi8pdI5KzAxNGfo/QpOyWQOzN1tyXlp+OsjRslyb+5o
bVLWw6BRV64mwMtEXg2El5fBRV8MbaFhu+CfsxMX65Gl90KZ4sgtjWyRUliVEPdw
DQEwEFPfeL2H6CivLU0iyep2FRdkiI5R6Wb15KxB4/C2m38aMWfqUdfSpy/4t1Sd
jXwj8jrwXOtZ3q7aBgwtUt+i1H0848hQq0kYJLba2qgRYE6WRrglnOso80K6nwWe
3Xr2rXNyhzcohi/zvtFMA6wtgCX65NsnZhiiU4JOra3R1T/CIzH9G17/K0U8DIRX
6kDwrE/w4vvuIDXBeB/T8jTvFZf6sLQdz4Z7u/t7jNZVTTQ15Z7cp3uvZSujHXZ9
xAPe9fa6cOlxv92r+Obm/ULUKWOAMjwVkjy81kNRuKDK8QQbKfmbaqrWTxOH4fGA
gPbE+2n3f/+dOOD+/HRAP9xJVeqWdCddhLsFdVKS2c9Wed5qWHymcfP7QxXRSfEq
azxDfFzdZcbbF+cgFRnJ/Zi/akC6XIbv8CrHCfXLdDJCTzkGgOd0PTRev/Najg2S
QNHhin421T+SscOeAzyLkK6CRsNXl4mPeh6GANmWimjLAPcn6sURf0KMs0jEiB0h
DfzRUrkKkl3Pna+pCNKo4zBKxjGyQ42Pjd6gMQUi8Qh8pfibjuEL4iG9ad9wT6HG
Qnbb/Tdk7/6w/sUauqb8fgYHQckLpD8n7R4oa8QzJ7kkP7DLcfjBRKrmKegfMWZN
XGYv35g0pRg7GIkhKy0sYoCi4KVI0ko8e6Yl/LIJivENju9SQE3nOc/NVilslr6p
ZNB/53v7ml93qVEIkCkuznxWImra8Pq+R4PhVVsZavC+w9HwlQKasefQHMzDiyxu
iu3JIB+VuSq955x6nmJjJJ3ooyMxcsYlHk8RZ4Z9LaYB1wDqOocNa3V8S0bkwCpy
6ZzM7REL9r+VWnFq/fFK5BFjlsqhu67VciOUfW30Jdkoa6Y05NjIC7RAQ1E37ZcA
j5nwO721Mt7aTKBR6JUNjUKovKuYB8iRIHqZsyy1qAKjwPpAcJ73ElYckMcKrZiR
U9kOQYFvXmFWP7rDPIIOEkp0oEe3DvUl5hoJbsqmpsl76ReEfOdgreCRVfDblYUi
iB1/QGG8awTgJGUurirGsWvubt9EGB4dVsyFpdjyKL/e/og6Z//Ti3dXTLCb3DR1
v1cSZVetML8enBpneMKqhohL5C5HCYlvtr1Ravc5W8yiDVxzv8tKuwQAs0IbS6oc
/cBwylmVns0CIoIVoV/XEbaHdIzVD38WhKpzQ3OO31rRn0pyyGXpMqh4ZhTPNMvD
wAduuBmJT7g3kVA6P/ZrmWmXczpktulH+IT6w0ToAr9VwK8eVPRzB99SK8ljgV6A
Eo0Hx9ps9mO17VXx/aMZX+xiD9bg8SSa7B2FWcc8N5hw8jn9gH/I2Q/JYtjNFmcW
zS0YAj82GowXK775h31ShDOnXetXq8BSTgdzZIMMJkCBfstksVZBV3r0IfTZU1GH
YdI5RGGprJ0PpcGG41QR4EaxsS0EASKCReWKy/yC83IZC6GmVHpqHXA7bQigoixs
m6xL0ckDZuwOOQIu+A6rve35uJayBMT7u4luGsSeI3H7g7dYa9ZReobwO4aFKbfM
gPTor9o5ecubHS//wHm82qoK7w9PWrmVyOmTO/VcPXyywAaZg/CIkWPZVi8iNCUX
HlDQaVJpIRMxHuOVzQ6lBE12ldrtiT00oNBhI4XehF4906ff5S7XEvg26mHGuz9F
ptGs8F9beiWfIRMICchNxpc4aGQU2ja6jcD6CLCPBwJesd/GNNCw4umcELYm/Lhg
0OTG1+dLstzH3SmuyC9BMeXmFUHV2/9iZkjye+nW96tYG7ttQ346QSYLQ7w8CclY
8c1ART4wrmrImOclUa72lYa1y4HXhM9yuoDd1drtqTbiIwmwlMSULOl9ijq6So06
mOHcjxO1h17GE6usX15MjaNALtGGkZg5D2yTwxJaEE+PQvMsYNwaoAPQwrbDJNUM
y77M9x+GNDc2bZXdL+1YID6jO66J/8F4/QkjzQiA3DJo+JXnpucVU2PAzpgPTHcn
ODIHbGvg1Z35gcitwruyaoR2T7dgx3Wma0wGQLvT+oE5uIT5DUZDkM1Ea6mf8Js3
DtdM7s8DAowoiOrnO4g12aYRonF4K/woOk5IDFacaAZeceB05AoOVXDESdrVlt9x
ccTIbkd5MEPVVnUmU7UU5fqfUdvwJs/iaUkqDmu+sMjRwZC78JRs2n5LIVczJEAt
Gn6BTF3yVyuT4W24M2weTT/cpfRBc7RQ4dsCLxqUDXura5mezvyFQlQNot6YyZrY
9SAb91PN3gLoxxR1W7lhksf6mFrRRhDfwAyGQCAZIWypWO8Dloz2K4+UP5Eh2UWS
J08qh4eHZswQSntMNAKuQwjkdWVqVfJ2NpddAMA+k6wslQRIaPakTLAXuJNQTsS8
64Gsiy0aNr3ONNQFuH4+UCoISrC1BYymOy2I/CLd6iCvti2Vb+jLyvAfZVDQo1NB
GwZ7xYpjsYSV0LKJpmixbLVsHx3DmlofYgHLkxNuwj/PbCnpOZqDWpBNAfuH6OS0
hbOhQafhXNqfHu1alZTfBV/NgnKW744Yn7Jm3+xhepyaYTMNliooP/SL3tq10dOn
lPC0Z/tGMDhhbRoudK8Ipb2aw7fTk4rE58/r/L/VpPopyLPMoiNpxAAscVZRuIV4
1b2GYAQc2mo38hPeFOOC7pql1w/+fhZ3INm7LBv2itIFzfHpRYa7tYPm5K5bnPKe
NO68pX+uIY4BYPbPWRCDnatNXPwrL6xF7seB9pnDBseFg2KbgglGxbo0qbk94GIa
PGMWxHM8t4G5w9TT346iKB86LA/voV6mS8lc3G36bZmVAdqffVl+nuCtEHk2q7Z2
72Rhr2rg+HYxnPwIEwpFYnzqx4Nac9D/vm5HslY1b4/ThJ1sH1ZPu4a12JhSDhtl
4cUZpHW1UzsqYnxypazH6uoqgxs59N1IGuI9JoVghZ9sk2wRt0TTdMxCi1m+IgsG
JC36YWMl3EA+aPCjsOpVXduZxL8XfkJG7sPWMj87jhhD6tivFsBPai6n74CIFs3Q
rlsoYxB3xwCfGfARH1zxmtzZ2USGrqJaoqou4mpWIZTB41Dz/dUeJfOi0+7WwVLP
bpvgkl4JbwEs1ApY/55sIlzva1mbzWlRSKVmKFs36oHRTt4TSA/V2lmSydPLhXYd
Lb8KntrkHXNV7vpTHy5OWRkAJkxSKSSIwOCh24KrACiP1sv26Fg/JHmxmUzbYFWY
0MM8WBZhn1Py11VfYqebGb+ltHJNYDNOO7teLWq5+ISteR02vvfXiOuI4toS6w2P
29gXF/Woqw5l8UpY1HdrtWCuNxMCSHc2cEs4afHI4gelPPE/ixQbjhjbyg/mdDjZ
e3ou4IpseJKfOqdh3yY/jKF6ixUbuttVAsPH682yDjKUQSRY+djbfEB/5GHw48d4
3YkN2kaKsKAzCwePsHDMsiKapyJFng7/z3RdR0etPKjXRyNfhU8udUysYbDN7PB9
HenJ2MPPwzsfpmXvhm04vJjWuh1mMaSBQzQYOL7QmKebRPdbQijK+22/q1d3Fpfp
cgSgqtbZFuGZWnbhnnwTLHiLEUVI335pE0ht5Y5p7F2P7nSjfBb1C5hCuNmTvh8/
MWkd3YBIVZK65AL7Ci5Yl+DSmcSg6ev+4b94shMyFacLQhzVDwFzvm4dVw+1K5Et
FQmXXQ9qeU/4W789TelnZUpTbFe0znfUOamksOLptVCQJA4xIQbi/pvk07Eh2cnF
WifuQzuwliZaLaAtZE3sq4Wt6Zu+hpXB/IZ/iBELG7BwowD+ZfHodL6dgszTMr7M
2GPDvSuZeamC92GGvgEbb8dpAs7Cfl1zzsjADoQZ3Xqa4CqXUD/TDN6adaRO5dXd
bcLu9otr005xmbP8eUMJvXcid/FizY13Kb5B/8k46ow6EF+OdOvHaPL5KsI1GNCw
P0ypXqq1fdLVCCAIzEzSxxTlsB/rRcZCU/Rg6HrkTZ5Ff+EIyoqQMosh+LKTPk5n
Y4/e1G01m4XIIbpzNEfo/WIjYBpmY47n7ghfaFeacffa9faxv7ouj52lgSezKeLQ
pZvts6UiQhAYHLxBpYmjRDhJunJSLA+/tx/tC/9JjLDR+4VQPoFo+gO1Wtx+AQ65
ZoqnFOFkmytuxZ9m+edXrFu9Wma9CesvnjBNDR33PgaCwMyVDhcNC8q+gmFjuydN
NACRWpCXLjHPI17TmeFqy5ybK9SCXIjecCshqu2LEcHZOC557vLe1U/7Bug2ULpa
fY2qzXBkuFhUiHwMAg3p8AhmRkhAfTnZ/c3vX4t59JjV7WiW4AS8XIMnNsEGElsj
gmjKH3gD51rVRvbZ1hF9MPPT89n8jat9LwgBggUjqfja3ifjYZe6Gl1EOxWhnFK+
XPFvUbmYY73EnFUeJiaQ5kazpEZhPE7eTI1zDZkiM6ZvOa1d0OGsgebz9vT1J20D
M34K/fEG4pUWLTXefAgHfKMOUf6tLo1Q5hlgj95UkiIC2sKE2/CQKeXVW2/99UlL
ateVgXxsv9yWlmzdIADsgfFq+lcIQvrDS0f19J9DCmv2wt/T36sxany0D2hZ09S4
fYJGPNgvCBM+s+3JvA6XRGmEptWAgdy/vreUxqzHxKZ1VaX9JkLD6Slyw1d7wHoK
acyMjRgBLoJsgWr7elVJv7lEAyobELp0ZnfNBrffWm8hUfdDdSvIAAMx/o8Z/cDD
vdNBKM5rJjUKuUFoLQyWFdTAjGqPrNWRZ3cDm5LAKA1Mc51OHoMRKGZma9aELk5y
pw586QX+quXAAUGemCrn2Gaw+YDPpATGLjvLyQc5Xrt2kwGGskfDRLzQ0qWc1CjQ
JaxvSQWX0JaNK/WwQgycyxheBXRhPrrdHz0lUofs4Bb80q6DrY21sCRamoq8ab4z
QpGxl9M2nnKWoOOM5Gq4u0m2k3n0FksD1nFOnA1ZVqHMcjMGg12YilM7feiYxoHJ
jmnh6sQVMLtZOCQhiVdwwuiG9DZ7ya+te84yQtaptFaRvmCfetFuoxEQKzKdIS1A
Gi96voaDmsEqE5+goi3Lr7AF0gwsRasJ1rDayoPNy/u9CdQz0sIzslcZt5R/xsYt
u/J+gyp/Stek5m2E/f6a4AfqeByzLcfawPINFzclsTmtQ8AsC9OKKeWUCIA4EhPI
0CQ9cF45lP3HYLzAxRzLCe1u4h2Fw8iu5G+4+JANLn/OqbyGa/XzdF1XyHbiYUIE
XHb5XNmHwENl2hfRIMvcAJNHYzDTamwGC99dbnhfWoyTjwvchoDpmCBhMLw3VZly
8hjoq7/H5rLg/bm+Jmi0iwVM8JfAk2xsNOOIXLgmwQJLyARyf8Oc4cZm+64zPy17
Z63ts/kHr1Vizf85cHuHzw/8HFwWZGOKgwgKo3gBSE4UNEdoCg2h6+dke6aR3WGQ
sxvH+ZBrK/3CiD5FyqteEfiiJcI2Hvi8/NMQG7v9cAlDJlhjx2xXxKD35DwUpQuo
nTdLY5vD0S24E44dtZZ0OgXBH37oohhPZ5ucz3KLn+kb9EsTcuMq6+7cN5M/t/wh
QzCjag38IdjE7B7oKb0HjzrOFmGmbQ3ofndhSrzKmqXxHVyzckizNNjtxGTPOGe4
a6cesfVazXwGyzHufxtqz5BY1OWDU0+6YlkhvPfTX924+4MVBO3i22HhnhiWDe6k
yL6wD6rxg9z8qvCBYzAeFwW2WeEU7i3VurCgY+4LV0zQin/zbsMVnj8nK25d7uRJ
f2nG2mrnp1VHjVAvJ7JGcMWPRb2VTN+NXTEJ5wED9mcZVvBYNJup+qSl+QwP8cqr
Hcmob/sRqxWroxp/a4+qPruq4dEjmeUuiXIEfTB6DJthq9edUIJR3k8L4GsMh/Ib
umM8xVxPUJIFcHAQ0SpLRQBRyny1gMsdyMMMI3qHGfibsuZSC1GmoAGML7wc6G/A
a4zLA47VNk26SZn6RK/zibw/4Bx+wgwcO6ZPZEZMsjLfHo4VGZ/lMeyC2R+Y/t5I
5sNg7V2l3b4PyS8ur26A38Z9nWIOtStp5xX7bZmvegHosdIuhq/oSvurRlZMFBzJ
886d0TkS9I+VxsKLzvWCGz+GPSgh77/aKqFgNb5jMyPsDtNOgy6PCUnHUj6nNpvm
OtyMeMonRvI/Htly6Mj1Qpxg4UxM70EsysNReNNO/rW45l5UcV3HvVjBuKp4mvxg
ff0IglMQIxLW3o11LsYwhQNw2M8NtTJx3dKXtdiyjZGkZTYRio73u+ORsuCY/M05
pZ4FWToKknn14E1GXuzMryTrGxFy/2aHYhTA7EDPoTslPn/iOQOobigqLxeasgSo
LGiOp4i2ZrfEVA0FP9wxSJFFe7lA9nPxeVoIWCbFAxr5bOVVw0MfeMsXiLglCiEs
TOQUDZei5YxurS6iQw2KJdXTx6zEstZkZOPTEaZ50mXN/cN6n2pRf+VAW4OvRY/T
phK5hhSww6SA8dtw1DkjUbBkuQ0uJ21f8Vzow2DwczXOQ6X7E8I77V7DQBCqS+Lb
dHFbaPOx84aiaqI7Q7xIMofPjDq3Oo/3YuKIJPlXWn42o2zpA+zySh9RdjEMyvEr
v3OuPsnKAw/8Jt/YFzSafS8CT4RmOrsqzn1qEiPyg5IePNpMeoZl36cOumopAEeC
tpN6/av6Zj1Ly7yqD/jqNx556o6v5lWCDLso5yZ3/HBgIOevng+uuATRn6TRHdVt
ogQLX4P/Jj0UF0XEEnPLWl0vbR0yMmQaJj1gsnUHEcXZuE2y2VvzvICOKo4DJM/M
d8BgGGTOXInn77fXHk2ePLxS0VRtojV0nkrkVk5+F2sUF+AosgNHNjSdP0dBNZ2i
OJCbGWwlvqsYTv75NYhnsepBuawa41df8LEsTL68ePTuYVhO+t43Nvc9E2DQPlWV
7nN5xChSIFzaMOwsvXYUEgHx5D25t4B2qygpUT5U8mREQcDgsdfOIhrbmCC3rBYK
wkdy3OQWqS5bRJBe0lwHWf6C22dTHjswNo1dOKFGVbB7Z0yl/X+S82u6B7nNDa96
q40uSjDEQjIjYNdNIWxbF1sMHl++BhBwVkGtuoSg3uClzs0Xr49RVEi1HXzgb2n2
zPMGTYz3xRW+h/9hXvyl9y3Ie3k4aR7V9PdOvAWdBWwKXCWYvTdCSfdCb30QqIlk
CeuClyfxQmymVgpC7ia/bdTcSjL1Mr2q/7C/vM6tczf+yZl/vwBrRTB9/ckuQW0Y
V+JRLJ3bCqdVZGwe77ui7/ieKQahtdqWrdfdM97tOkupcT/tVdiJ0XekxtT67f/w
Tk2nez2JNO4rSgCGQ/tLn2UmOTJIn819zyfw1Sg0sZsnfvre8+9IJq1pye/nN+Ya
bLrM5Tk9CaePpJoikfpRZSTtoca9X8G3Ua8N3NQRuU1NaVKiIzGYLS3YiYcR0gg3
P2PDxxX3S5Z/48v8K+v56d9aA7jpsSHt0IuuAro+XSa6O6gye2SLH6/lmnOJG6oz
qTls+VqA6B+0S8hIkomUMf7DCZR+hoQ1q+wlri3LWY/qoIH+fJN6doWABafec1vr
FXNv7qjs2Pfz+VVxxhkpdbVPvIVRvQwLMZFBqzO6VndtILkD20+vmsIkZu4aCky9
p8qNaiSZJPJqzhnRMy1UdeSR6CscUsT1YxNCP1jOrOxzyk7xsPJYLjAQ0+ajTg0J
9s74GFN6dSjuEscED02OCiO/BDQUaSbt5m6odG8GV9A3yUWjE6ZvdzY67CsHe8yw
xG9PQ68TMnpCa3NKxspUkL89a+QLaDn1P28DC7zqcy2OvgjRPeYGJDklVBS9s++/
07xmRAVApgKm6XzXteIpXlfRxUW/Otv6TPznJ8cjnGYMyKYxHioIcatbGsOUQfHw
YW5jBV62t9SVHl1cgewwLa7zhtraMoY0r9agPkHIAhuJQEBL9Ys0SQKqlHy8+02J
b05Har9iS7cVRjfqKpSpUvbQFimFAQTHCof0AMKkkUYe5TXnbN5rm2AEFb4UZZHG
8r1PxbeVQw9VsPh/BIN7hq9yUNsRG2NPmEqWY/VQJOWHrR1U7/3TUmkc75KRxo6D
3SYUVGvBLRRc2JPDp0yEz+7TR86EJ73m7fMU53aUxFOpwnrnBBL/PXDnU91D48iR
kmfYEagnl+2HsGqyw/clK0cvfd8WGIWv2x8g0nGejXL2IgLJkW6Ju2l8sQJtdEfk
5U8olpH3/zEKMk5QhEQvi6bUVUeZ0v6pBrlAQsABTYYY5XD2OEgjkUmcGqIAviGz
krWadaWGb7AU/YQuupt01nVT5M3cu2Jh3IAxCMEoLd12yBWz1dExZxAqSajbj6dd
Ud/Bug5pwKkCw39hdIGj5+9+N379EYLfxXO9+qVzvNBTNgGttqDcGOMMe3y6XiLN
BUZznT5tCR5Q7PcM6ehsB5nT1YYlavZ6+KZsfMYvjlYSOtnPb6uC0t3FH4V5qPDL
IL83x9lDONKUSbQipaGghCYX1sOc8EbCQRI1ehIfwLFI0COO/mEPUiKoLEDrRP56
9aEpK18987b8PVi2tZBui1hITifh7tgH/79V/z25uEm70I0rQRuZe7Idk9swdiRo
72NYqpq4nZmQkFRyi5xyAM5Mse7TxlB1/Kw18oSyqhxFZDfcM8hQdmmukhlIOcyQ
B8WsmSEUKe6v+QZCmcD59C8J9grCxoUXfVH9CuQMFaTw2njJ7j9Mm5aXPbwgb2kE
/x1DfLboi3I0829ovoVIKgP9uagNC+SXrwrnPn+Y1/ePubhDaRl+NTvHcSKxPyLY
exk98n/VsRLJPeOcrz+RxPxtJ8T+9n7AIpOW1Tx/6/xi5OJSFffGwB/5LCO0033x
ju2qLhcYeGOnNqH8MV4QI3JfKFS70lz2v/SJ0UV6o1enWNdsOCt+ii/W7WFt2OBA
WRD9T4xt2ULkZjLncz40rF1airvPK/K69fJYluAQLqdeE77YndrKsW8MjBtNLJlO
OnslvSlgSegYAka4gS6ZMK1SCPr55Z9Yf6dvL7aPDMz6VCrCXH3ah3HmSgwfO81j
+B4Ef4m0DS8P6AazPFp8/kdYN8PcQkE2/OrS9t19VF0Q55npGs17NhTkdUeTls96
vg0YS3h9eXZQypOAHX9w3dwyJUjX7xNqACn4GGmo/pg/bUy0HhNvxAG4xB5axrQ9
/NfDxqlukkPqO5ytZ+UV0byn2ma0beZqHeF8wSxF7EDx1rkxj3vRr1GuNgdnppoF
EQpqaqixyPymxMh4q+U+yPBokEgO6yRwNLJ6ddMGtXmQEtHf3CAja5twnIxQ9IqF
foaHhaxW0nBju71HtrEz1lsRc4PHM/JfPvo6SHMWrXL5+jrJN52njky3sKkVWSbq
kz0ocVYQjbtLDRf0A+lcHKZ9BbYdOFBnw4ql87fFA46MSBZjbYVYLdIlNxF5S7uq
6ZhwzEsTBAtelO8MfhyB0CLRULN57bklNTPDTbxVo8fN52iJS3LtMBnua4uJbjaJ
s5a+8E9pzWOYk5S9v+ZKdSWCD3S20ERy+OykxE4TQvqs8I2wDvp49D1iJaQdVcn0
a8rwrxAt1tSWZhemCbkKvjhziWuS/dq6Fgb2eddGekJHoEze8lbHC5jD8QqTMWWV
qIxyoKYOMcCKoPCG/7/RKe9qq7+OYr2WcSQybaePVw/URl6AKY/4aFjUJ+BK1AFh
QPVt65A9oX26pkje8LsgtSVX39OHctnCAoGCWksghGr0b8JIpRzjqkfeCHVSfjh0
Mo+Z8+x8RVShzcLMcoCAx6NPFNE8Yf7x5ayJqVvh0mPwEs6w8+aZgvk6JyiyFg+W
wGHt/nHTYPAXbtoulO60wS/Nj+a3R6MZauM6j9zD+8zA1kFhBwwUKoH0PdgaGEJF
6yqF4rZEr0wCticoN8QaMcpDbJglGA0DRsRTcBSPmhkrgRYVk1e/oTzJN+ABvbjz
p39rRt0vM7ZjGpeSuHtgLJM3vIFwJvpQ/BY26S9wAMNWPBOJDLyHCc46CsAbkVOG
+HldXcWCx6qEvxYoQINDl1riO7gs+7Y4UfwamS1nWj/rJbrEonSL35XLfPWExr1g
MvCbOLLi3no9Jes193XG1q1hnRosdaOM9KOMqxCnEvhE4C3rORLYvttcVDwoApYj
kg1qwhBkym0BIDgwOp8jjyaF90iKu75MIiuu03nvl3IZCJtAq5kS8oxERMxksrJY
pSFZVT1hJ6f9wBSrbD/CKMh3xACIMBLAdLKQf6AvkcI60l3xPHRWAYe3P4ZGSLui
YkKYVAYnpptPGVw1kG9dcTK81t/OVBnUfzEf5fGTH5a/oB3QTazjs+vlgQ/WJeMH
6Nto3AZVA3SGMPqutZpWUYwEQLSNT0iW2NMmE1VZlqsHnTom9aSZHvefpw9XnIzp
v4+VAxFz+2T6qaYURTOiDEFgfv5BYKHgC135zqKbStrFlM1sP6ol8Anq4wNF5VaO
NyiFK2uH5iEwcjPQ8oo+R/1gsyRSltlUwz74rkZg/Wvv33pA1IF400I8jYQeBKsU
wfQPyyk3juGZndYibtyOT8QStdt3RpLYWGAnG+OOe/SwJyAYMPjHJ9W+7FUALeze
6owmLFtnDZHMHxQX/6fR/DW9H12+xeAdqwRoXMitTioDnk5J+KXI069NVFL9b5NC
49WS7pAEMeH8v+AmPqEgsk88jVMpIUdzh8y3dMhPgcLJqAIEVg+0NQSg5qlOS7kA
HGKc4ENVfn35KW6iNogVLVuo35AtYIdUBtTfpxieVC3jHpZkTECV7JHLnVL8Xbim
aU94k8vw3Pg2rOtVGTbFTOHVuQvp+wj2PpEwrUtsPliULBS22aPiCgboF1nNX+7Y
RId1uH5CP8OsHycJunV/I5XgvFKdvSTox7beSx+07Iu/j4c3ZyZ2HqQgX5E4hw5b
Vj6qRTZRBJej3F9wsgZFWyBjNAMhmmRHRq2pOukQ7/NDWKB8ztMIAKWpzpOa0Wnf
i68P8EihNZwGuTMWGTWVCGiA3KM9uWus/49nVYsMbX3c3q01jRP9pkjY0BRd1bGh
tB+J8Us66feTrXOVlDwFg8fCGe3bcOT1LHIA3wGO0TkNr2tyNiqwtjTxM8Vmpu5V
dp968Zx+LakaYUu8hAuRU6mT0Q1mybQ4jKigpysshb/2dPiDtJZ8y53o9fia/AjK
KxtRIWWn1wjTh8Rpt7UgTpGszLx5Qexwob8KbUa5f7vIQZgqT3bxFJv8i/sCVybs
pGoe+ZDSLjTrpT+4/7gYMBZ9wr8C98BiwRhEhyVu+GbzwMZpr4CE7+t4hPtY8yBu
/onNI9x3dImJhMBqF4Dykw7+rqerzGjKoxbmqtPw1q45JYMcxhS0V2Gj/sIcwKK5
soHAArjyiyXf9U+3Hblo0ZPDHUqqwndZ98o/8IHbqIpL2m+TGMvTw6eScXa0Smq9
ECRCbq6U/1HMn4w/cnOTluTMPNuJ/uV9c+fpQH2Mjd3hjNWqB1QbhfutJzJxFYix
JFLT56pJYVbBEdSAWp/lvLdeijNR4XMsBqX0L2pgz7b7/uXLsBtd7IX2uQyzWrYp
D9LkDpaJEaOFy5/JG/hR13e2il298L+KPHAXaYm1Yp78GPFip+t5vQTy5CUAl4XD
tj73b62kIYgux/SoYguk/5VhLFYsFuQ0qHSvimMEczi/XupAnbmB6GPEprmYi9JB
Ul7XaAp8t+9E5D/N2BZdKy+fF+3mwPBJscCtDJi8tOTEf6V6S+D0R+/3ajTU7ceS
MMJrkPY2fnLf/r5lgN02KEfaf3m/YZV46Yp5djnJKbCttgz6FF3gaPHiYdastnJk
6xhto3QjaXw6klirqZ5HFFHP4+mQrcSmOYVZ6I2mVoQMKaaAAzMpaT9w9aYHtkxt
ffMqAYOBRmVm2Zhk76qNlm6VBspaDDyJE4GSF5L0vGuvPFGIEGIyCYmBGUEzZiAJ
gSKWAiGn/nnyAfsMyCZTh3NFacVS5xsMjgEEal7EiDQMYUFTfeC4rKfo+GnYa6oh
qJ3UltoKjeypzG+J38Sv8PVyGbAUMuSMKIuy5od+Zm6PTQvVtZ++8+HGzTmVfN49
S5eZTJziqQdlNU6xkKz0kdHqwfM1wlJyQIqoz76X8o5VHeNok+qFbqYOXTAJ8xUG
aCrGB8LzF6LseHg0q2AKoQ7RbD4uc2XQh3jyx3TFpFSSQvtJJ+RQpBUgeD8BAk1n
iSqXDrhCUhILEVIxg4Sc260IpysexHA5wiWT9RJf7nocfl7uhIwMi2kXBe6h3n2s
cIsqI5c27ZWlVEBLgsLuIYzFnuLgKkbyl5o/XJh/vBilbgAbbPpJ/8s6ckzXDkZ6
8ebAQphKTfUEMUFGSK46ljYuSdIyMBf1Pz9tUITsIkCDOZjKFKIRLst8s57COhZq
Zg6d4imn0RlKINOjWOwJJApPPRa5wSET2GVFE8XK3BizEbIqWnGqD4hCYxDR9hsI
KjdaNCHLWm+EwYh/0vFLrkcTQFTL8e3gbizn+1ndRVobQsXj4juUNAMQFixw0Oxw
ZU4C55pcCjbFS5J55+ITBdHv+/nihW8/ojOKjhqroTh1T2YpWDGTW6TCJtw0CYOf
hnVGsdxCP0k4Ec9VEZsP2u8KMeEQZ0MQ1dcswsz0PhC0ByCr+yCsL603sb06XApR
UykdnTvLg4otyUBNNyAYH6SlSvhvgqxA4H6kqhSk79k8fbNxlHrPfGIKLrDDiZHv
HD3UFZw3f4fbns0YqBm4ZSNC5o3HtU73GoODvAk6Nk61LXxx5IcMIgI31oHJF0k4
/qPVeM9z6JLah4zx89JfFL3FcmaIYOSN7zHW4w9VLmg6QhUopO3b9F05qk+W3Q0n
LfStvmQM58kKce20z24VhSatHuPcQj9NbaVrcxv61c4Ar5x8kymbcZNGK2Yfw5wa
RlKPNxMMkW5qhyRV5/04D4+RUL3TsRLfB1qKKTMoUQQHQ7nX/5bun/Hv6xADT1vn
IXJwoWkG1zZvJrTrlGQcO8lMlKTbbIzua/VUhtYq7ZxwmKOV0Fro9zm4/ULaE8GR
OnZifzjF2A5ROqa+cMpASlM57zFK6X2/WwqVO3Yi33I2y30FfGXv7er/5b/H42Hr
1XlKp0i6SdCFiajBh5JRUhYFgKJiBXzt4o0FCgaIGkPsLCRN9q4eOz/Q6ckxz4H2
T8uDed+9YK0Hxi1paEK04apb910iRBVqa3FJZzjb+U/2+fd/mde3uzd2gGoVei/U
kDmszYt1GRYS3AV66yCFr9M/MZjm0C9mi1modkeozw114s9/xBeSWHhE0LozD0Ln
QOSmfgV3hsxQplCt3x3VcXwr5PCEzQD+bM+1FIFO9CIVAI5GWXMOTL/p/H3i2EAj
rtBqk/8L52oewdFURRQsLzqqrXARj6WRGLFoqpiEIn9cns2vlfwuKNzVfI4mNHpI
F3bKHRFs/0EecO54Vs3AuwZ22t5UC0q/w4MKEnRgZmH7bDxqbgi/YvGsRudi5Hfx
VEqpEJUqmAS2ySTpAqNXNDt0ZmryoaSbTBbc0f1RjNU6sLF8WV8n+V2NXyj7KwAd
nhnE9LXUcX39U8t8IrySqGeIN/Yi2CvkUkDkQ6V6rdGH63oACawgM6rukzmPr4Am
UO4cTIHjo7QayCUQ0/SL4o8adp7Not/m+CPSo7o86+kmh91l1NNSTbnoN9ACpiSS
s/2KhNkwa+V6y99lUPiGEMkY3LkAeO7Ve5Gukj/woM8C6CjnUr3Fm1ukAQDL7jrP
dQBox7hlez4YJey1YNy8lkVqie/8SOBQWVonGRomVL2GNDeqKKkBenVIs7t57p3m
1zwQeVknRRixmKs4B63lM4m7CNgVfdCILX3rWGCIjUazMdyHhz/nIVXg+Tv5lV/R
cETKfFn5TeO/wMT1+QgSK4QhNJYuU7cppR68uunytWMSZlazU1e8cFIY48X3l+Ui
zCpg7PSLz/9RltYwbFG8cfKKO4nqLvlkWSjRya5XO339V7KXcFYs6gviG84ZtseB
GLuBYnJaqHBPKGQnDkk9/zabhKmfe+JP4Q0BH2AmAojam+0t6WJ1QrC8AXfpBBRL
FY2tnCH5fKrKEBnNpBFhmzzpVJgtY94WHOSeEuUWQpR/2jAHPF2nyQ+LLwV2ck22
qBI2aAT7bNKJjQdqx/T9CJJSsSsN/P2lMvjHaZy6JUrhz4MKdubEAyVpp32vxKrL
inknkA4zXAFpIG3vhqc6qIqRI+OK0An/6KjTXbxN6EHAOAzrUCVdqvRTnxbKAjab
JJ4AKI6LUdve06SvJd+YYeP57mSNUy83GV0xtly6qreqF4dCHbOyODcLsYur4kHf
NO/4TCDj/fi04bDOs7mWynemvlh5KpkgES+lIqEtPoE4Rup5Z6z7KBnW/oYGiSqr
5xOx3Yh248Ij9p6iGITcF1uWVe+9C8ydm4/0q2HNKBvR35ewG+fciUKXvA2rya/F
SSEjtLN/awJ/sO8AJ50/+0DclZxxm16dOpmCY5JWM9tlHl6ScgGswbWs8dxQQIdb
0lxfSFUbhRCXU578x5Ff6twG94iey0P+yorCYhDPykeaJh3R0ppDs8h+7eI2abj3
c8h/wS+oCjBq1Hlwfw2bw6cOTdOoqER8isneNNv1MMK9iOYimRMzH9YgRtte0CAb
xpkLMd6/OKHMT/wmP9BZUWUkV0ct9TXdGzKTT82iM9QuuNHVMIDcLw8Zvjk4KUdk
B8/WPiBMhug253xrHC3H2db8027DqnhR7j8ONriSw7BjDnf8HV47g7kAY5JiVWE/
GpdBbmVdBTKdzEqjh90nFMs3DlaTWaKHh+1L+blKJlp64e+CNTsrRjpD6vrYYnp8
LOvsUFh7yvcqhz66vcygaoehkRS9S70C9Fz42mYDmNC6axR7RFyQHr4ONx2Iumoj
xcHWDcf+tvunBbU8LKeOlTPl/+zAxxCtV5A/SL6nosj1pMGc25txkJDbS5A9oMoR
KpE4a86dCrXmgDeeqbOIkSjlOFW+/p2jMLlK4XtQHXjaZ7hd2A/BpYuTRVMEZ8Wo
vO4tUntfoKeq1wQy2b2ej8sFHh7GaDbQqboRgYTcpds/mVUbv5+fmBg2D+hQKry0
VUUBAWYfXDemA+2xYlxxaL7WiV7o9MV51PUzfirACAPm1tyKvqmrLRju//BGBVzJ
MZA9CwkYo/S46gY201POe70HsKwHY609Re7Rs2zTtH24nDlykCv5xTCruZ6Vxfnr
UFmwM3AqWwEN0Cbqdm69/SzYuZyXjHTaQXcsYHcsUSr6r8Z0IazlGYY6qOUgd4e+
5OJ2im3NjnEYfDyIriz4/5YUbfAFJLIuvTPDx4nD6xsAoaFPqsQu40jMUbflehIl
NyZbr/hxXK2atxX0dzet+AFyrjv3U8V9i9b7Givwum7vLC3I113jYOkjMSAoh+PI
JN83ghyGjqvk90n5BKD+3tD9E/neZWkDi/4LBT5bgDmiBU4fFtBCABp5WPoZLqwR
JGKnd5HqBdvoh5eU5IhpVmd/GEhCNukZDUUYQVTtf5pRhzDD2YRYaa2No5iD6nLA
KRDyB2XlxM0X/8pZre1DdgVjvZgtYDGi5FH/9HBm+rp9HadhTokJ+3nol8koylHI
bksQ+r7cbnqWNDtfcsu8H2LesqqWItz2IxsaPe+aZD/J5tWkQxAmVC70ytTaAzYp
2emaaIds8tUN/nyj9LbpXtH1PImji4cqWcLD0MjliRwTxkDOWtj+patObROOVzjw
RviO+3QSd77jPhc1gUz4nun76Fn7MYz+6aLhRoF9AhJL/MIpx2jCPnvpFHII3gbO
6Qqtcmg1swJ+B7vJu7I+RG5g/gU5chd1T1BWbPHhb0yF574PHnQB6Iz5YvuTIq8S
9HrEzpK/8vbWdBZhBhdMp7ZzZTLZGLScpg5zsQcbu0b0KXE5jpJdzBUy/gOSeLIm
CTtcO6I7qDR+oMV9wJma8QmoUPsJCeAetij6wwJQX0TVlC1ElWwA3TFs/yy3rxcl
z7u67F2kB87jzHCnYnm0mwX9d7Yfbv+g20Faow9Fk1le69XMw0c/XFOqc0oAnFje
Fjr8uD3wOyWkoZe4vezLO8zIbSUPawmYjvyfQ4OkBFCGQkKlxRTD5DCv6AOTkqSH
0nD9CTUXI4PukeObE3719JfzLK39xqSY4l2a6czAePtLCy6/EJJKeWFOUJV9KVA5
j8YOBUaD26HRmopV09t8cPavKEo8u/QVgX8I3QrbfDqnhXtKau/YXvH5ad6L49G/
pbfTyqmKLYpZeU/gtT0e/AVnbQ/7G+iw/Lz88449QyzPl5q6Q2wNd5nNNxIvkGX9
9Fq1+P0PvaI0FGjp8Yawu2XlQn58bx14YInobrkv7Z6BiVE3dDJd6xP+ETLtImKi
GM5hruS9rJprxmxUjPDJ7KHBimFcqm8W8NWLyP76hNcKscAkgIt11Usdch9I2J5r
FgTrDaFFFqhx0TDwnDQz50JEQ/H9m/ijjfJY7nEms6U2B+U/jMXz1JBFZEfNfQDv
f5Fpdq9Yaxm6ACEPQYd9JVbkIp3/9RaOJ88r823sPSbQmnPSAVJC9mae39DmADEv
069xBFI+XTXKmNDvvJAinBCtYEKzkyiwXvRz0BCVhG7/UAYQAUu9raXlRyDCmjAm
VEJUd9sRvdL4/2DkJflJMKzd/HjMCcI2/HoRkHOlORF5pb4TG/6hUzDNudHEohFE
VeveKWfUnX4O3KLa3cChLjVHjhr3jPgPt2rP/kA/WrQOnmnFXI60Yg+HZ1CYyAgQ
wlA96aByY/h8DcYi9sNDPCG2WAaIN7+jM2f2sc/hrRJxM2IizV7S0na+Fc1Gqwm9
3CPR8+MnhYJPDighhK3YLbfoqPW40iVLoCu62nrh4Dazr/hHetuEfO49JkI6JEti
x3at8Mwovr81MnUug4P0K6PcWI4/w1mTzd1Lry9AYmy2/19C9wVAxBIZB0iHc7PQ
gmNWTNGY+j/Z9ADWw3/sUkp7ZkO8NAhD7oz9NZvNWBWOVHDwsui94px9RpoJzwwf
ByhsETtVpaugYUKPSSYqpJFE5agwWN6TBHWIawEy8ppwjqCIXiit4tZNWsPj72Qx
Ts/4Nyku+q3MZw3DV3d7K5xOJhcGlkNB5JSZ5SyfenLAw2qvnombbZisP79UY61W
fnfHer9vA7gU8YMnZV5P6WZp6H6xwRGNm4MqlpT4iRGIpMgm+odYWX4V7r+hx5zN
SO6MeSozK0b9M0hlh1TokHN8q2aBADDshKgcw0swmV8LRASAYjNVVKctYSlOI354
GfsjrrQE0qsTfYVDVc08IU5ktP7PcWiHOahEYcsHJ3Fwsk4NwAbyqOOB9Y1bTEoJ
qCX0CiszWzDa/xoEAOprxUmeLJ3e+kmwWUzW6CbF5hJ/NhWFbXUyzqFqJ6kaBRLp
JDFTF5KRBI/20UEax00d9W93dypf9aAFaWMSyCeDp+XW1LSpONcySXBpmXTIcsCo
nUorwALHPvCjR8L1G2W+Agk5RnuqFauu5HZAI0tCl2sf+hV+pSMWP82Uj/gLHUY6
z21DpaaDnzTT8001vTJ1uzz4B9Y1iqlruebneVlVPn36M8z2K2PuNcwAS7kAeZbA
SOUVKaZIp1TDiDq17gEZiIKFfhjIbQj9rXVFEV3NRnFLRgTMzaVLqkQusKmuGcWS
iZ6/Icu1qqDVXUZkwNMy9jceIXZbio4ZXEpQ00ViF6/FwxBFM6jLdWKGLc1odYwo
HLozxqIPAAjXotD9uF0Pq3eBqUNdctUlcIsCheRX4NQYCO5wKqZDa3adDzWIW8Ru
nNFS1KLemCSbtajBdZP4j32g4MZl4mu4u6Xwv7XqUoUzb6r4QPOPnf8Uz+sRukOY
xxT9d39L61ArDiDDUY9tBKgP1RwzezivcAI716zZPxAAaJqukytB1mXq4SbaYPgE
eQWt6hMF4FXsAU6fYAOgLrp8NYVXRmvnM/B1fo1OhJYlw1o0iKdbRHfCIr83Xlxx
y1j00iZ04ItXaKyCMZlBU5keRUjP2LbZMe3pNCrsa6XxTY2mxhxLDd5ymuPjCkCV
+FQRYUOV3iVZbzwbpG0b1W7f3MWJOCzPYMQ2aTzMrAyUeTIPq/rEkNq+bC1beiDV
QSJ9mA6FVLaHvibCmesrmXBxbWcOj43zHbAexVqHgDuUGX1JwbpyCp1ZPx2HNYwQ
032MiiNBfDvOmQ4Brw80EoXYCeMXHCnX6T9ILw+OdBX3inRlWFwxsJLeb0c5Ist0
bb26MHtJQIK10MhmGtm8WhfiXMDVlHCqX4O2ZEL9/ZrC02Umrrdgjc3hs+FSVrkv
/I/LaXCCd9bmO7+hBlKsfxAtz+826iyuOVhKbIX4nPW70YMHshJ2M5wkgI//rtZL
KDkbtWW36SpunFzCFxNkXwRxs6ogv//26HvP2M++vSkW4rvWLqAUND26FKXRKLTM
rFt7R5oikx7lgvMRUXlvO8MvkC8OhugXYLawknt50oWt7HVqI3e+WYN49XaTbuGA
kvatMmJ4yu6EQu9FTCFkBJmolXAjZre2rglEr/wvLNfwxBkUf3oapDzEMvECWHXD
VD43PisBY7MnkuSX5ftKn526WhBPPYHdLgUVL4Lswoi0Jn83O8RfPqYKR8R1lvIR
iU9VT6Wd5zhrAROeQwcd4KHelBT9409ZyizTsv9PAbwFC1Zy5g2r4BEe9XfCwtux
/hdxLP3nxeYOtsEaHJFOyiAfziuczfEHwmeCfaH3HN74ptCbm3yRSAxkWEbixDik
tdemPJC010F/94tIrpk7YHgtT0dxwXE2w4hEkj2TAo+af3CuurLeEm0XMhqk6yTY
ze4y9idY1n92WTAXz7Tf1goZgjgUMD3fb5yPFlPbVoJKsN4zh6tv/QaQplqpF/9K
c3wg0NWDIG7loH0gbvK0klcqhKdQTW/qMrLYIPXq9a+AXw424VuhrNoqDcMqDjVk
I/D8WonB7Mi5P29vgMAmnLVmp5HGM80nw6jYFMOalMpF2u5xdNAmzLep4WOsBHIk
6Y22+YGbJ9WURlHlWC+0u7GqPSg826NMncNhtSBIMfgAD3/S0phcWSz8cYO8gQYy
b6/FRbdav7N6RQrNECxQUKBwDWriNqLEMTN99NNVvtfpxbKBoYPatidh+OSv3Aaf
/GnDXHH0NczdhxgUwoelElz+HpYrPGtQzvtTdbBB1Zqye5WNyb5bOpEIrA+o6C4I
tDNBMlG51QTAs/dylwpU8t13GQeBZPnPZP6nTov8n2yOyDC9VRcz9YxM948J88zM
oZR6cZBzvKec5xJiCF8aEp2kB87zSI23gc8FfAc5p55cksbByLCwZAtIRAMcn1Zv
DOI8dHQo6lZNLPUiz9/aOSXqEeDDQ39gN+njUNxnxTpSdwFJpDiNI+dcvhx4Wc65
qYXL0NHJWlSmmA2Clf+SuPOe6PGfdUAIlyEkXlXrJqWCFpMqmZNl19W6I0yNgsfV
D6OpGF0S8JmTzaQ969alwrihOd+HdEtKv2Fk1QIK9spbVvIsQur1PMbv018CbTlM
MyZ6RhKb+djyBYauN7lOyRyOMAovCOvpinSz6wb/3EuJWtUtsQoLl7gR0w/Ikk/G
bnIkZplI//oPmUSMpOV2Rq7uFL5SXvPfdTuhqZVVS7fHqIZao4YuSFRhzTU55hnC
xteSjsOSY2dw9pD0RR77tR/BBhBrAGd3w+T0LcXIzD6X9MMRBlkUkKsPxkEd46JA
dgUGPUfS1uJbNQjbZoQZacTK+/2mYkPuATS+Oafazwlc5aTYE9KfAzJAEyw5v59Q
P7REfQDMutQlecUYz1MBqVhIvDANaZ7rdrJ1vcWWbBXi0ef3HDfzDZBmgtXY3KAp
x1UMZzpypOhyMjcvpvyH9kAsjCNyshEMwOJbVBcv8E0LZgUJ0gDOJpRKHsNDKALa
sB+d5Y5M9UY+M3RAzW+glFcKRgUXKTaM/feB1j9ADsdYGvftrRGS633DyYRykiMn
bB/2eXotJrCBWy1Fc1AmHyGnWkiYxbOyBeKUHsi/eU/MN8kjdeoa5nUy/bwXTWKx
wtH8ziXRfaQ1WtcjBRSC5EA63zNcq0RSKKFHlFabJVuns2kcrATTZL4mRaEYfwbd
hRXCAFFIfzkfmmno5d4tjaUFh31fCDaNxkB4jjxW89qcwoQICEMV5qelDakLCKdo
gRZ00d2MmkddoNvrlLb9YzzjO1o1SiWg60l8LQ8U1Oo2ZwcxelZtSpg6jEiwaMJX
ymB972ycaDfcyM6vrSYAHy8pj4A2Rg0pzMY3Sv6SUQaLrW4/zhVOMDPX2+tldbwg
i/tkZL/Qsdaqyjl4RGPuOniPXXdtpORzyE65dj2cQFEEC6vroMokViscgWSVRhRN
KQX5B5VhJF6nl6Ef3ldptQ0ZbsJfElWFyk2dJeQEKP4E6yuBAsQDW2eho33X8rrn
2muUrRrTKBZFzh6b5kYepbb37rzZJC9QwWqkjg1YDR3JSkde99cVlUcU/1/xLU9w
s6L91Opl0byHDPzgOqHn8KT33//rJzHtkOLtx0/6k++q3wt67w36pkei+Rbk22GD
ljyqiTqIOc7Y4wmG6IYwurf3rHqjmOaKeSDjCkm0cfxHo8g92Sh0Ci0Ei/gXYh5x
nw/uLt4+zyY9d6tOm95cvkVqsi8AW2Sp/7tp2AZi4T9W95HLTT12TIpVxsa6v5bS
iGON2L79BKXCORSP0WKz2BdqhZy83oIodA/sj4T7MqFET0cqgO2kQMo4OMHNtvDE
8YdYIyopxdsn5S4XWxVuLItbmghPTkznddHbUyhJt3Wycj076wJZidDbvYG+0usR
yB/zNw/IFdkO5fs2nX0K/i4sxzYZ3I+4kZwM6JbI/wS6jztiDnvPwg7flDDZ+dUW
6u1YuE6zkmRjv/b/bXwNOTyY2hcYunlAZqGLAIPkL6y0nIzd4HoK5QnX45QBQw+1
WcKYt6mLUWyQU5lLdIQUPbq3vDaynN/NPj1SohQulzgxM090PItSWWOIGzXcYKgf
DHJFMxdT2HQn9DUBz2ADAAKyOGacUNDijtWT6TDwrfo7csDisACSOE+NJvo7kf/d
jrzg2XJ6a5gkDNUkyJCSqw+FPih31hyn2uOW02hOF2qcBSZcyYfOPjv/7W2UMlB/
TbCHXqr1lmL78onUuGWGeSzSpSL2kuCA7qfRVjp18S5uMHZnvx387U32pAZsm2xG
VghEL+WYvJsxR+bU2LkW2/F4Q83L+RCUxV64yuqouHK6BWGFKzyJAag2A9hfpHGL
REFXFzP6etWJbKsMFfKgdZjSH4ZNdb8aPWxu4z6s4/9qZuP3DEXv1lmGm778TlOI
l6rd+yGcKN/rspQJemScl4cxXmPQq6fA8qacBYdG/hBcGGgf0JZ1ekcGPR33sskO
UcAP1WUWJ0utsLcPv0hgYTYSRK4hyY5y8X95df7U5ybAqEJ+1+/ubbFVqZQoZAE9
FtT7iAuiwaZYWmJa0uFRM47ch0uk0rglONW3OH4YEn5CI/wZ4/+N0ussJsFWRLyw
ier4/IYs5FqaMkJtfjNIgTq1Wx2L3TsBlivsp6P6htpuIT8b1fWCf5txxzFKlyYo
FGdicKgVPgcZ0bC+xa5Dh9iLD33fN26ceZLDbSE6y5jMDad68Yrc1FwvYghkAKk3
uuvg8mfVZr8HqkvYfOV0OG1cTJpZkwCvDLV5yvOTJhL2P/5CcUX8wr7BqPiTGJyc
qSiSqlxtv0DOeTyeVMV7BixbcluVPbXU5FC6ji7UlZ0S2o5gfDfTL01LlEwiifZi
N6lwnBVTpHgkAM9uxn3yeNE5FrtrqlOWWTbdFkY5xbz1yfcuDbLhxLfuAHE19kM+
4I3ewzMXoA+wnhVmQ+eC2aCxttT94fuuMdh/Hlj/Gm0ABvUPl+y4Koycbv2qROmB
G0lCByrUVh82+JrBaG9twRkPvksqcX6eWiygMpCOI8zsjHPYpkfxf5O6xdKuNOLz
GIFHRkHD/evVOql0JW2gBpk2FeVPYhj5qtKTEnm5iLl7ORvAssStUfCuAb9I7yTJ
i/M7RL+mtmT8iZEjGeN6rSNF/1gM4oL8qd7XVKCQbRg0W9BfwRPwkXV+aQZiuIgh
t4xsR4Pu8hhbkTyGtXMbFFt/HBIypNyFr56GM2IYfLomfsscHnvy0mroUZlNZooZ
qWVC0gFI0ZQ4RGJQ5bECe8osAVKSxzpMIil3V/3ndCuwLUQXYjjL74cZM9jC4eDD
+er+oLW5GC/qFClYTaqY1tc+nriwcNo3TehJ3mripnwI3cGpAMMx8uNvEJmIzltr
xKt/5ceaMe2305AQ1BTlxs3bnqYDP1BMWqMeH0UK7fz2AcMkJxzvzzJKSb9Ii0Ee
yZONlDraIaoatUoXDt0zweXGmPS28akCvZqMPG1z9YTnj01JOlonTOfhdVdNiCdY
1FfPIOaYf4jOYW/F9R6chX1FxPp0EBzlw4gfJXMvsE700wl/TxclBI5lWhTJfZQZ
oaSq/622IP8djAGpSqRwRjB+MUvQvnMk37Hi8849HSVKbV6VR7L9asT/dTcvDZ8o
u6mc1J98qT/MWnqu/4oxtPfe2Lr3twLZU3H2vyF7rr+FitjwmYLd4EBBN1panwff
JwIVPgs86acHa1RqtGnoVCgWQXeDnke46dZKLlR0em3Y94hsdk4gQZn3TBdlv9Te
PgfNd82J1EirvmIltdJBsgdK+b87gD9Bdjzvkul8RUDQzS2D2XFXsEX2I1D07Xt8
0YJ6mdlrXO0Tl5/qQ5VlK/q8+f6jma7B6yyvVFwpUA7h5xRpxo6GYJrLZaB3/gdu
OjGb5S47wNFGFNtlBV6rP1N2hptwJf9W4cdlNANyVnRirxPJIdWgHVgb7UYvclHO
fn1vchH1K1Z+yIs7Al3d1VlJ4K6RIi5CZ7i9QC+EQ1vXkTppOTHNfdaVh6lBpijt
Vol5iV5TRMAIPVYfxt6Nme1sUuMk3Nnb7ZTNQO40wC1AYYNl4o186blxD1ub5Cju
B7y0+Ct/bBCtXlopuAgZhlnYScIRMm3KmeYK3jPANsgDHD5fF9xRcb9bZQT3PLmf
pSllLHhvttw+E11ApOPG/s4M7wl4ianWone4si9FYGdy38C+tjhpKNJO1HBp3JGJ
GhZGoIDFuvMIrIuCNuU6us38rwBzNofkrls2eeo9Udvts66bnqifpdjqkguN56tg
I0lDKlTmz9nfQ+QQ1OzAl9KCk7mpqoSsL/qo8mijUOGtrhx8SKzb4FQQpArV00OS
282rue1+Qj72wepJCflSd0cmbwVncK/nPNYtpnvB2MCGeEjkPXIPabD8o4RpmOm2
5lxS6Awd+UHsfnULeq+duUifYK6dGgqRvFCImOdIrnWTQRvm7yajz6uHeo7AmNfQ
ehUGWdJZv+pa3bniYhYalEGkVtrD9dDGIVavrv5YMWfPVU1GaK9a3MkKum18B3V3
FxDHI7FvPm/xzucdlpjZ/BPnohm1DoTxCgm3jQOxMuH1tO3BPvMKLFxoXSmBasrR
5NLwF++dJzJZvrWV9xvaFqhl4uU8wsSCkpY9QvXT+zynxprQeTT3TVqsE/5hr2Kq
7XU8hbD8jL6KV+UHC8Y5El+QnRd5P3Z5c4g10vKWZufe/GPtZfSKwRyGvVYLgCcO
aI7t8MYT0pkN5F912agc0UHXI7ZZL/hQCqX9/Jn50WfX2PJqToC4BF9A/lVHaCF2
Z1jrgrv7KyRWFUp3v3wG92uD0pF8YDiWXUbW8vt05bRuCHFDicgz3JaLnf1UC2vL
YhF8IqIQWqJWQNlsNLXyIZlvGG1pElIhEosGAly2y6LZE/lwEOhiBHZrDiEbLlo7
ab6odmiYvJGPti7RWT8lJ81kUdpWTS1hdmWRSppDG8/KDKzKs/BOCno2LZnP7V27
XJ6XdlmeVIoCcCqDXxFPwcw2ClCHYOUpVno8ZFoKf9sdI5fPpyXPMWo09Ibq7as6
3hDZGOiFcdOdf4ZwZFEnZaD9MHLvsEJwohHaUBilOX31SWjfHEE+PJp/jIjGTSbo
RUrsinYAjhjFYuCI2x1F34cAQUU4LSgODS2K2RLOjhCZbb+hK0/JZ7S8YkSki8GG
Km4j8s4KRXFp75ey9XYbu9C1w91E2iRXSm3OXahl8KrYROERu39SZQQkNm7cUta+
AhM3Xt+V4il/KaS4JMScr//vdNu2+tHjsmqDM0AaTzqR5ZUwZb6QFR1G1OOItYLr
2hYN91aod/TqSHJTkrTRmlWncohgPH5J4FqpLf4mljiNalx8KBBe5exEHFe95bvf
u0hhBzk/NgJ4MM708GQqKJYkyOlFBLekOxi9CfK5RPBxNQUYAJ7MPqxk5TasLndU
xCNTO6v1WF0o5Wyev6v0jOr/7zWkyccyyNlNfXv/4hWKqWN/APafjycVeunRmjMh
4LhdVaTqb2rR2Rg1KbggoBfY3pR2wjpCnrswMvP/+RfHwzdrkgMYQL+aDwgmpDCc
L5tRVDMylRqABLJn7m51EN1/gG03T0vq6Wgx8rUavxv94xzPcwkBfenH9nDnkdGw
oGOpRCV+nqsl3cXVSFkP6iMjzSnQXKuAoXoBBqn6YQWBiRHfGQNkoSmvI+jVszJm
ZR04iEGNMip0Wrxno2u8EynvLuqS59iGAeVs6ABpewamwzSQyjUI7aEETJOHzcI6
jFuaRUmcx7gNWmuUtcbJt8ZOv/bQaccjYzdytwbf4CU35sh+8XEiTMc8rV3Ni/7f
htTvP8cvospUAyrKtDpyXXAe2qug1jXZdrFZnpaHx43D4CAjYrWXPUoIbc1Tfzaq
qmMOhimQefXa0ohGrYkcLAu1QWYVOpRITuyL+MkVBNhdBFQq4ZtH/pXP791Mpu3Q
R0YGLgSmEvSaiZiu+Iyg7khFNQYv5kLii7gpSe2r7vau3uKjEN7N/pB5drhy4pzi
nh/MV6ewxeFOqdDaItJGQgcMYiJe497tjCRrun+s1ibjE82U3mhkT+ga/vli6ASo
pcAmUBnd1V4de3tucQqQXIPFFXZx9XWxwevUQmlRQuzRMKr7x2+UbwT3rz+SJrE1
8Lobbo5GLoWCSMFomZBCMFtEhmPtjoDozW70iVQQzkedKNqXpe+xQGHidpy1lmqx
MxU5Bq34gtuVoViLoZdLIdZt32NZCqLRCXvoIYG8Qw0K2YJOYzwA0tLG8J91YZ4z
WUR/RttWpApOARdWGz7FlS+82Ai8WXBI/r4eOci00fyU6bt7ZzvfhEpxvMgO/Js6
RsbxENH2fcS13jII7wz/19huz+cQ2BSbzSoAE5iPaKQWj3XOYJ0KU2xGPxji+mys
2mYrllSrEtncgPvEfT+ga79JI6x4GitzozkkUVQoensex05dPtZRiVytORqk9Ftq
TqRf1ZsrNN6bbXCpbtmtUPljW7iHbAtQbVa42Bx0X49JUJBmdydAYz5/38OugERG
Bczu7F0QM+2OivJ2LLme1OOAv17Gu0NmKo2AhFQjj7ImWgs796qU0uRCgutHer6w
v+U3cY8MGMPJ2tTfhqSJQ2kRo+UFqifgtJIY6Oz5S9KGpuhtS3KxgTmB1y0hNl2i
xp/Q0MkNDRFApHc8jc82a5pVRz9I4uIAp68rxmWPgxgI2fXSNNkCeuJRqJx0zcUB
Qi6G0rh8QoIE3rUjC7Y5CgvsvkU9iaJO0xqaLYgXdwAmdxFqUTBQzCzDVmLH/vKu
oTfeuNrqwLy3D+ItUDZw8w+e5VH/CGK53se+1Ck/0QwSxiyfxBZq7xGMBWTpQ+xe
mjEW08De+94nWNedovsOY3YaGbmvJrP+LkAFr4ighXad90IBipjfvUTSI2uWSYRh
ogBq864xOYNceByxcK6bTUZLaDhCyXT/sNvGUHep0OSKLwgiQPlu4FrrE/PMi8z8
dTA/FZRY+vxJ7CjLKwpKecPNBWNq8OLecq/39yJJJCf8Jyuk9LZGNaEV+JOWMxk5
T217qrVTgpqn0PcTH7najdcgC/xz68kX4oKP0nIpVpb9O02f5tVT+4ZSIvypTIWi
pIpKDFI5u4ylhSN5+Q1NaMFMczDQq4XNZT44V8cPpcg9Z2+NzQlG9dBw77wxu9pa
AgMsLO/eLn9QzN4qwzpBNxvmI9j9PjwEvPoaNkvnOMl1Kugj2ukMALlI9njI577k
HjmqnpXR32EWFiTJ4RKbe2swyc1CNiJYXulNsbMT2O46kf4hg78s30mYDxgjDMFu
pEJ58tw2a9zH4mIMFqTAeGQRmuLKapwTyd3MuDwb0mZVD2+mRZSua8baBZxLV0Bx
YS+bte8JCSe9XO77EyCyG+JkrEsARfeOsjIvwkSUeGcAObsC6Jvpf0MC1GnflCmP
uzR+08Gd8Pssp80m+kzGAPtc2iH3ON1WYt+tJlq0Hk+w6I67FpDbPmza7ftn1vcK
6fIdeckzKcvIS/XGjZaetpGPMbyrdTQ6F3+tQZmBh9DW7gKUQeEznakYcAHm2EkV
clJVjMhKcWTH5ZoQhsfA9RnbvfPSNcQlgLFVhIFRNzDPwKSr5mELN4SmJANjbVZw
adlQc/b36Zea0YTz1ZYPMWOZnRE+Zv3VqVVEIcSXd4+xQyLQwy9vRu6ZakHJTBhQ
SsGwYzwI6h8rXKk/Oni5ReGuNTZ+9FfIeq0oNyvHOGOZsfJj1+22pxdeY1fAf6aC
ecwVdPNi+orSkpTMsPmZ7VqhrtWOBQYC7iCIv9r/HwtkgKwkzCYTJx0QVfYaNycd
ErAGbgl0trQmYEDcp/pL6GZkdsRRXPwjCykYQACb8SorpILoiCnAR87S6Jo7/Z44
WjV26ifWFJTsz+UGIg1vXqs3yGMkUbGLjGqh9vua0vpaKLJyMLNH+e9vWcG6qhTJ
TXHChdXQbXTltGltXr4ZmVUW8wBo35qpJcLQYBkNBJ8bCpfVf3dznnQgANBtLaQ8
TM+KrZ1my/x+7Aqf89tZNSH7P6g40C+Z+Ebwjf0so09oFkVFfCsSdg7BSrnVDO+q
tgXOyD1cqu0Dx9/QrZuF+NkS2W/ApsV8OPgP62iVA5nch09x0d0CwLFheIHnizn5
LhUQv3Jm3eGqo3YbngjdCKsCmFSlcbmwPwKlLG+IWdPUqSPpDEC0KweP/DchvNCj
aRYB3eFqF8nwzta+nuKfpePGyQlSKsWBkH/TrJfytbyFJJdVwvCiL0snzJq3IZ/o
Ktzpz7zMGxxUXTSOvl4DcKN55QEU3ZSJe96pvyn2pWarDqacQOs5oV/jbjnjT+Me
yl8U4UTQ9Sm6u+piNVMmOIid7e4lHj+XNQbq46Vs8tWWzzutNJGIKooCrFE9ZQ4i
oIH1UZUrWC7n/0seI2+ThAf1Rnlew0uvc/8DFWEnLdtUSRixCSiUhPv5L6m/T2eS
OE2qiX0oKmDCeU6ElzjsBmchX6cia+9u3WNAljI8eJAf/MXO5MySr2VetGOp81av
q8SHbhnTgtkUgduX9nv1whna1QSZEHTifdZ6bv2oCpBBjDPHTRYqtbTwpUFQLVzq
YSRZm/mu+3z5MC/jzwd/Iyp4aAKLkAqMigXc47YprGfQadvLzCMdqOeN9wkQ5eQ4
3yFrKhMYLQoCnYqEhy8hsiNn6DggZK8qpLTTgV7lMnsZ1r9ydqJ2rK6hzqca9h17
1u78Otttl4XXLaFuMVuuXbJOI+RzVaI8ZU0ugUujDvw/HBwtOAEJUcb5BY12cXA4
XiN0v6Z2cWNi/cf9iazm3DpUVC1MgrwgDWqP+pSD0/Ge2+6aNZ6fAEHqGUywe4J3
dC5gTU1xsGU4KtE2IkjHPNNlgWZtO84wSlet3Mqwxc0izCyDVrWREz+1pJL82+nC
i/N5YuQkwMbjNW9jS5Ry5OHIFTWKn4weQ3qBTAZYTiYql0N3UwFwoecW0Gjh6Uls
DGYQu7AKJ1Z+FuSsT4ylex2Eb4r9lsvSzESztZ6R+h78gnit8q62ZtcSkovbynCL
VJvW/ThZcVMgflJSOKyVj+ptGQUpN6dkrgQbsKMysP7CcKh0KxPL8R0AGRt8uTix
JNbzrWDdESfqeKKxMPEzaow+S9wPo8f75e3upv2Q09bpIHf7kSr+XZ4T73VcGw70
U/PshiOIWjqj8vESo4JI7tHBxUwjPbgfEUnh+42kAS9uTYP3PKRdlB52KPkIqt+3
Di3yRyIaYiAtat/IFe/U8rnmLYY9gjE6v23kuAl+7PCCygbN+joLX/ioHPWeyawk
YtRktc2AAZ1DBOEO8guTvFYxiYRPI4HJ9VGhyYS8tffvyOfqoqTz0W0tDBBMwUsv
GDKHLyNoOcKFvUZC0nKfXtM4zzaD8T2U40tE6XHhOsN7BXU2KOhdQzBCmM0/lpUR
upzYK0Lu84Bw6Iu7kyDR6YxW44Ti4uMPeBnRoDsikXKY5SuAmdlRCfK8bn5PWAZm
05uC/4Car9lprNN+UYNS6eLTI+DiMvbzkJkRP26LcjM5NkVX4EkLI07Y7shQ2mQ1
fq4pvcy/UeEb4pstwCyNTOSpQTO8mXVwJvJe0T0sVsZPTjxOH/2lg4MOBPrvgXU6
+MZL4TrgwEhSe2DA2pVmG/nygiVrVFSqLjzj3hPTjczIFV+p+xmu12ze7MpoTfkv
WMTl4pvHaTr5mPI5Wf5YdlOX0gGu3ZhIAeooMom0d501IwTGVAb09naiek0Sz0MJ
vI07p9avwIHqHNZQA9Afnfed7k55RGUFkeusXg6b1U+uBXuBAXQVQcXPjb4pg/Sy
BaX1ggKmsmIF3XegBmL8vHyd+NEUyHv7fd33NHkoy+03CpFWUGodDm7TVVXUeBvN
8n669Gcpno3+I60kzK/sWxkMYdpUdkA03k92qte26f1kf3pMoE5PrLn23wL4TkVl
LJ6SBK6mxmsBgQp+/6579qgQBLZOLtmojO2FqfD7/dXixhP6iGC1h+gzbKISSwuO
CbQUQ3vuLZEmgrAqm2wGzxXfS0qUYOopc8XEvya0Cop3a2skhVGCDFnYPAQKl7CV
c+iV0rNQk0jf+n7p9f1s7EOeF8KBza+0YuYzgAN7sMI2XT+EJ2AfNdwlGO0c7sQU
GohZLk2MIFeSyl72tX6eBpCKyiiLBS0+gVxDPeOLDM5BWFjFU+Bpj5L8vVppgqdd
jYq21GlWoHmE3moZb9ViiMHzNxcY6g7rLjYMBgIf29+VrGlLPqEFMOUOhgv0mx/6
X4LPuM4YSWFD8emR2++fvc6tG94FNoxSxOmsfeYCIQJwLhlc6TynKFufd0cnHQAF
1x3FSLKpa5xvIri6YM+dtG1kIDL6bzG0xtwf9zLyaDptoamZJv+Yf2FKm4/0HQg4
VHX1OCOPcgucb/QeFnMKY1DL0aUroqFcH8s/CV8NcVr14uhT0lHz3vSVR5Zix+Rl
ZlUh2q4g7LC3yhpzQtq69e1vfPkdFbWlTuLPnskQ+RvZ2+IIkZYdRlnwKhgKivJE
itNwiqPO01XwxV4d9lT1jrJHOZUtuauB0n9nQa2H1Scg+csUbjjPUCZ8cr0Dc+RU
QWYfvUqloGnPcCSIqyayMGGhBxMjRLeSl9ki8Ph8OkPqCI95uy6Ki8OTz9tKUAZr
BVKowKIRcdGwSeB+CnkdRM78lwngWBRMOeclnq6XRhtevOCbalrY1U4uOjcBIXd2
fC3KSze1poVoB3oSiR//+pmIXKnHdG3Ca0y1UPknep3FgoffostMZ+iYewvbgGSm
4+gwugBuZ2qOsNQxpR7HRBJ/8u1R0SB4tf+D3BtuPc/6pdZluAzDyGOYYzGcDoxx
WwiCI/GT3Gj6167y0ETxcmV7OhKywmGjUNP8zCdEVGsDonmnE0agQwzkrK2ZA5D/
n4EuTQAR3EDlKnpAR7IcyazRS3YDx8EJvuqIrW5pFZQbQGrhKiZlrg98nyYJqrQK
ZXOYAnzMk7vGlzfB/X1J1+h3vQExNil6h+yG05sQ3lkA92iZFIwEnqYB6do9YpK/
XSgPuDAV/X8qq7SLg58+A+bw+kZTdFb8GN2kwz512cSQjS7iEEJF0Vj6c12qcHC3
p8ru3bOCJmztvsNYZyg/fWReYN9YeESJAayjzT66oxnCbr1rOfKuQIcwvrknygej
OfI1POoSvWZc8+7mmdhyhfWBDJb9LBBgNSDK74nJ7uoIm0+VsNxrOtK0YQ6DS2/F
dNxF/+TCttQ0qFNP9YZYU6Siu/MTpkYtuOjpxlMZZ0WXQDYLl6L4dkexe+AnEGWS
uwpDv+A8wvhg+GmzrmX7MZtpVmNbPWKvY4RmXuFmwthQ3mRCA7rCKaFH9XIv5Zt3
aEw1t8qaFk4e1/kxY1tZjOdIl8v1ZlQuh+bCM8Oe0WTBOTwAi0YliKRMaMb+VPji
zRg91awcbrKf9KTIvRfaTrv75nlEQyISZ4lI/gVmnjZj/wuyZxPSykbWK8BvK/GM
r+gvkU3yVgL3vy5UxfvPUiV53V3JkK6QGj35jR/vY8KH+3ErdW++fUIBVA2Xxw1/
Jhdx5tavdXBjrkhru9utSkzY60dLA87Yp0dJ4e5wrvrv9rk0Wo4J8iK3eUPqBuRm
4ewnSvV51RknKs/MSu/MLhY4yaIljYXBH1N6QLLXUeZEDzhYZTfGpFt/lqiZAmm1
qW6MkoZ/8PGLwxBNZYY+nt/T19HzZdsjSZjtMGlyI31l1d9RhTCIsDQH6BBo1QJR
ZIe/jV6B4YfVIgbaKAnXvTF04UpWswvbZYSmEPfTSVQmCTclvKQ4EWOUGRze/OU6
6kAqE3iAnYAOnIZi1vq88N23ZwGHKOuKyDf3rgJq+tft42weTaUTOgvlEk044sGL
nLP3mm2Vl94+QwOmtI0rjjOPi6AC/Yw8PVOJru3f7LBLfWa72KWwx9k2Bt68PUz8
r+p9IxqvERfB/v0i8URLPhm14/jbIAsuTHpptLn3s9HnUeJ5AQE1a+qyH1PfkTqs
g3bliITuZchJE6+6nv4jxPc/FiWaRuGsQywA9z8fsOJ+6AqGjk2ddCWahW6vrYXY
V6Atg5AJQtXCh1uMUoZrgaylu+9SbTcOfnhN56ran6H9Mwq/IlITovwH+ragOP+d
YK+RUqQZ8ng0JKSbko+zFCYsjo6Wkxbn6G/hnyuZQnw1rAJh/LlPYu8pqPn3OBBC
gH8/WC1rjLNXUt9Hir5mV1SA99dg4+Ic0c6M9wToYNqu9burEZOfVXDOFEsuB0Ss
AG7HvmGe6GCrSy8e3liXEy2+aHRN0FormnUV5E4JEuGnlipq7CtPNpZSpzbx2TnQ
VIXVlSBN6430CGrEGqRsPARiUfXqgkn5qZd6Y6G/3Xk25ufW6tl8+jst7TK9diT0
YHKYtTHlNdExGxyIFIBoNI2cxXhPlfMNUY/DN2pIUA/gYZws9LuV1TJom+i8WBvt
/CY/mtwEvFVt+vMdbbmCiavkP8SzTdOe8/UrlT1+DACJdhWl0pI1fkDDFovsk/Em
h3giISF5cKQRVW5Rc/XcxVHvTgmBX84m3cYmI6h8YTlZDvJ3NwUoz/b4/KPlXG/z
6EhmaOAZbbcu9izO9unuEAAAjOP5hOtNrLznnAwGZdLVHIFr07VFwVsQxAqEH83s
2MCfrulY4eono0VyGA8Dkh4EsPL/EPKpNvbTQjpiFYg6e7iRRNphP0XuJcUoO1oG
ZmGsP0InyQLFizSFS9jVL/ZT7KXJCuTokeUEVodd5O6vIcI6Zehf88fg5ORHJ5ZE
7rIoVYhly0uqWNMyQzCbihr670nw4pnFEUm7odrIwjEEFAX1ai3eHOywSLS54oOb
hgVvYMJR3oZzyGRuXE7XsJXFTctewoY9nIpsoIvtzrMUm9I3tkrPgFV+PdmSbptA
P4Y7nnXN2IuGgvCQO2KFIsOoQHmD6wAB0KAA+1KIN80T6rnnd4CNsAkhunEW3u1F
1+F/9NFnCPds+cmWCg8dznYpYvbZfuJJ7SR4RNWXm4VQqZwZdgz+/ReTh1gBKtJM
ovkXdG3h0S5lN3qHKD2cjyAitK6XOMs+5lZ/rV3GM7/CjUzVSdEs34oK7wamvv3I
JXJ5VgzVmCkv8lj6zVWTJL1femwZyBpjJF0cqmGFQ5KIe2ZXu5JZuQTr6ukMi3gz
ymwMhmCXW+DShGCbXloIpDt+FhPuU5SvZAkoL2713WsRrJKLAlQjarXDkHDQBQIW
Y7j9Yg+gLuDYi9LSW7DqWxJdnyxQC0cGjulPmLd15MaR0wlcFghPD1uEAeJm4335
5mS+jBXe+b9KpMlVC9mUCPSvxbOubnuRHt6DIwK2r3J248w9uq8V+n+CM6C9rRt/
RxRR3n2FwnyqWUCKpg7z2QjyvjMjVHtIjLgTIN4fy9HmV7Vebhr4ZHJ4Gwk/ijcI
r1f422QhaheuyraxIPHNHRN2vfIGMzSkMIWe48DNv0eVi65yp/SNXgNwxPG5Z4ad
WB2zHQve2GpH5nKN/S2NiNyW2YvmxlXdr+G+Dl2/6hFt9XjUoXhZOytkzTaDKwfE
9XBOVtKfcdra6JyD9Bt5+dcMK5ItKm83a+pp4McH+IjBJXlng/MOzKHnnHFB/luG
0LIzoRVq1/YnAx1Z5BhnXAf768c6QIxhAVp8KAAkxag0JMaVSJolRd1HnL1Z45X/
IAFfRBw4q3F6Ss5aVOujpI+lvrvxV70EV3rGPN6J43imSYYqBAD4nbXlkiwb+wgI
IUMz3A2OlOQ8pRmWrbsRLgUo6SaMMCLXcB20OVA0SkGMUCNkjHXk5wWjZDTG5ogJ
06BQhtInGCupiQ/GNHGOSV8XrVqFIBhu4xezy0gLo5MZgrykWPSe5DpEyjbXxpkm
5EWN/jA+hi5+n2J5p4ryeTsMEbqH5MxR5amP8FSFZlQtFMOIJJcHNEbuQQl8aUq+
XjUjBzU6UoKLvQkwnVCA59KJR3V62irX0X/xT56VNPidd/sz0p61QRIxJSCNg0IT
vmiQTcog8F5CksZ/HXzmnwMn4rFzgzmXwXOLy0vxCRJPr0kuFYJTNcKO79PnMMox
UfhuoHQqS1To5PIh+/mnS/ggYnEFHrYg5Qj+Vmb9JksK9eJOwMvt/hdB5auvaid8
Kj+PpJcmTBUF6exlGkKtAQ/XwJIoHd68F7cXcnI5tetA503r64lbRimFyuwRuAw0
U4eUd2Py8moGSQVWrJPYFKk3+c+WMkbL8EXayjim5ShzSF5XChixNLWhUHPm4l7o
vvn/hGUdhbQoCiHz9h6Z5vx6x2WPNfyG+/xLPCfE3NfcMWFW9XS75dA62Ub8Gnue
T+N+0Rs60VMomrskvsL5UT8+LH5igj68qxojDG6Qdc/69ygFnDWwEqGr1lhWb8Mx
qgeQCqNPPjjV/dEjxDbFWuc78yg3mJMioYIRd+sZGlKcpZnAVek34/paYciAdBoA
EZR3ObLJD3Ik6oM4rju/8cAxNkQPmjfQ6vQrOpqiA2Rggvl1ZwXA6/urk76V6Iv6
/Zb802Z17zUE/XZYtTKKunHxnFoXgXVJRT0g6ADTpgNig0OUmnGtKDdr0Q+teIZV
1hIrZycbxjIsOs7cEgPoaqW0LRZx3tgaHBd9pFAp/Hzrw0PYO3NakPFwkSFdVlDh
R0SwmMMU6vvx5pxV++5J41Jo2PoRiUkTePO+cZeVgB1kUEhY75fWK2mVq9sLJueq
XJ/wGgnp3hzO3N5BDYgMH0zOmFxppuFxyPKZHY32udWnZmmTZiRmKWZPxz6g1eeX
90WyV0NB/UHaCO1HrdykLqJcleCY1GNcw2bBQT0Y6gKn/Xp0fJ19j+BP11vpqA+1
W0eGKEisE/sMNLsanxK7t3APiWkv5HDQ+hVHy9hDMtxBAWwrAtJFjseBSvFRA7rO
PNg/puDLUDZZRLg1YM7TUNT7vidqYdOdI2Jhk/3QcoFsyxA2vOeB8d016Qxxaxse
i3YSveT/jy6vv4fhrRpaWBasXQ54O0lpnTOz8n1mUD9k0qAODMREfoME31j+kHEW
dkAg3aR2+y3t1P1ubZV9V13A4CH44EF/l6Zpj1VXQZBBxgO+VU7qTTeqH7lRhRTX
UX38GI4HJO4IVfkHyBGlT560vHzQ8QzMiomh9Ry4kD18KHV+UoySJRvRwMni+5Qd
Ud0DN6khySAIx+Agnz57d/HgXJ+Ug9ACgcmuZasRBRfnLVVrHngpN80hcSpikw9c
OzZF4tB680vsIAlMZzDpGHaudbCrcq9gCr9n1KwhREC8T0Df/ZzRFEuRCPqMppBq
9Y5/YloMpLzABkPI8VJN3720ecrMyg39wbXPD+pgH5lUsqmdU8dTH/iHZtTNHIOR
gmKmrtwGDu4BLtMqBlR3YPMHOWR/Anh+VHje53bAh4D7vbabfDkS6Lq06BZKz2ct
ZEfZfoVqqXdpm3Bb3GqxIeS2qkJAIvLc+wq0HPmz7JJ7WIPNjIVDDm3rlyzCGhbH
TLsx7fkKI7XmbRFEYzM3iUXuJ4Xj+qE+pKhuGdl+sOpA8Jo7Nl9fu/aUyYBbARDp
fP+TxD94k9U8FfmkLzn8kSo+Vfa30flFnFdI4B2/68TmK8l0DZNtTv1oLT/LIFOX
GPlyJ51T2x/1len8CjzukyjX6lhO6BPNNTLIBjl+ydOPb8odMzixVZE8Y19rN2Tv
f7bng/hN9HjnkSFt5ZXuNDz3W5+r1/mMamTHCG3BBILNwFYVQvkPMh7yn+NTJVxR
vwPfowtO+gjnOw3ysQ+EmX+Iqtcm5TuJP2NRmQA4+iwSJ0NlyNQdzoyLfWmZIrcd
fn2rs6eWAMVUyy/AnqIw4KHDhwmGmfKQG4TcV9CYBwJb9JENAW3r6co8H/bnFDPZ
b9mAWyPEgfflOxniB6jAwBYVJYSgwLDSJGma5gRB5tQdgr5dAuOCmzJnbgDbZ11i
+Nb1PV2OhhSh+J22QuaNeavb5bUsbWRbaVBdp/zshGKSoeSGxz61ad4/AFO0SfZW
Ow3fwMCVmFYsJHnizf3GqASDIwzopAcNbYQej+BwSX6owbQrdsuRnKepmIzzoOW+
T/IuHuarFfzBdNY9Ta09lmh6zht681eLiJy/sBbSgS9GDXjiP7kL3fGxfXoliSYV
R9dySOH24MWOrPoryPclAAb2nOA9QXzSaIczl3YWuVQs0soVOnl0KY6LR0tY1YqR
CHX7yr0WWPFJcOR+WoQg4C0WNNpbpwftUyWOVFASQlvLpYRyiyLiLRZyE4XwDSW3
vubXAUXigxLadFotbi0hT9uYbcj6anheczw1SzOkCGLVR8hXi28G6Pzwok5wGbi4
hhcBjpCVlR8RiQ3d88txCJzK/sgyqEnVX276cTW/ygLAh/UgfiFLJs7XXcviMKUM
V1MjPDZAJIMov/xlHkiXvqeRx88bSKJj8UFgX+juwW8KnqhR8zN0Yu/yY3Zk74yZ
eMHclxw8lvdEsFBivbm8zd6+ROF8t8HbBZWcbItIKzUTSY68dGoVisH6c1ooSrrG
jzTL87Il2XBGGi+lOCijcxrkvWVrwcCR5f0Z2pJpfprdyLQPgGYoK4/J5HAu+hZ1
JtZoPQadRgUTwSdMVfsH9ZMHjKCaeF5krQi61H6GmLqpMDHGQQKpj30j4PY0GLBn
u1Oxe9vDVNYjYJusF+CzUFVRGAASwaHb7LtHgluKR3NP9llDcskJn7JDS9x/RhzD
PTWQy5aAjhTcq0NLb3d5MQ39CnX4Ne7vGtlx72FqxLzAgl/4Riibm7eCMd7YGXbJ
PzIJ41vDDRrwTKJhaxfVBfOYrGvsNyeX1Va6D2L82jyMdQvypzxu4I+eotvxlRxG
WAGFXNiR3+0MkILpdEYTSAFF/D+Q3dsrjp9Z6BonG4VaGd/fAj5k5k2siuTh3EBq
TAOqYRTXhiZttzAejgBmQ4AV6nZzFmU+s6eNKw88Xvjna1SSPRJLjXT8nnAAIwkG
Lgeq9v0opGXIOjD+Hzs28ctcEXbO3ObRMK3OV0UL1IRn5crYLv9BOM1pqSPA1lBh
cinG2o0UC0t6M8LJAOlzWpYNRehLjY/Q7DYd8B6wOHeA9uuwsBm3YdCvqRCNqUo8
qGhti9HiYhjwk2FUpWt1PteY8bnzj0rl+8cRJoZS1zD+FqYDYx93OSIgV1KtaRpt
Jc8u8+9/yq5oPjoz7DGkqbgd5sVSV88rdsqba3qTWbMOd8PNuUSKKkVCtgOm0njT
3h0bCepWtZPRV1o+OQdCwy3A3peCqtQC/OmcJDAMyN11KLG4JqC+rM0VPTZ2LucC
xHMypRVhT4PsDL5fSc07D1QVYVG7Tjv+9HgbJT/0KO3TI7Cdb2c/agl9aufiYOM0
9N51mkLHlVNhbcIkIHY2sC2ubeJ+yL5wNBPZTNe0ZWZpf6yElcuD31m6eRaIaje7
ui1CKAS/IZgrKsE1Pn6LjHHWtU25ZzvhW4wbhfO2QC5ZD6TC7QqpMZv2I5rDuBki
n1/lTcTEMhVYCWvWxgJ79lZcX5f9j9kjgR99V6PSjRE0u+3syffkG4Wsn/lMUBW9
UGJEcsdVYqcAnn5IkPZ5Mxj1G04fWitVzMFdb69lCUA4W/v8M1YeHuhC0r5Pxd5q
OAZ5GYER+yvmVvUWARhtFd0WhMzIbc6mRKwtREcp46BK9x3zORAPacXI472F6B1x
2t18AX/l/WX1BXWtzKzvA9zfQ0+mfPtZr/a/1A88+eS67kyfPRhkYKbvEQ00Kn2Y
maytMaAInK8Ae6jZ3+VbxzUC0HEmVvCp6BcZB8i1ERjV43lTBZ2dPUFSzA9/FX86
pdfT/+KDebEhxvPYTqBAO+6fVKgsogjFemJpBf4UX48Hd3F5r5sDUOPzL9raymz7
wUBK+oKec82JtE4b32nmSgQ6ovD7aMQ48WdM7w139UMjDlHXIzQAgusGcogyO0XX
I139S1xZ+WKSH0SE4sx4oKuoZjg03UfxO4rP0zTXuAsiSuKyRaoz/t5BQ7F3js2v
W4jHG9dpDYpZ/8XuKlFuMn7ds1+83FVnqxA0LXigmgwNGc0XD8oGhjsWHphPT8wN
1z1O09EvufU1p1shHwR++sfBn8fn0Fhxw99W9mmteQubiAi+IiCVrSwUprVH9coz
JY9t778UXl0Evrul0gHW02zIJxQNpr0xG+mcC3BmVS9+DkPZ3bW0U9wWOS3PiQOJ
O1Brq9Z5mGUJw4JKZ5SK7VoqgS1XqSn9DvrqxjwG1moZ5CXdKkxv3l/1bJmHqSB+
DvUMEquPe1tysohK7MFYb1oqvG+Z0IHyvCeINzK5rKYn45zRgGCHwVkOF8EKosg2
v/xgbYZKfS89KNcoUzAU3MR0IlBeLGiYw6vMf07SpsfJe9WWv5KboOA0cwSpoh84
avFAmp3sTNqv6ELm9ArPCc8I4obxNEPXn7h9CExOFSvVG/vHtNPbrMqdofHyXrHm
OC6kWQkaAoa+ScLOBA/4sQMhqgi2M6NMUtH0YqkC9T85l4/+lVm1l1oupriPxgDv
8F5iPg49asAvBzzOpsjyHoP3smQHPFwNQK4nn7Q1rNHuNw2OCdW6RkemSQKw+FvU
zEY3vumxJjcApf47jpia6l3l8ZvzFBhXpHTX7emj389HQgV4xWyv6djfShYAwDEq
/xoLSwcGG8mvvichsmMJLeq2GY7ghsfXyTUG8FtdCro1T5Q6DFmzNibYQ8hId923
zF6DOBGzrSb1/5nBsnVZeli8nVtAd/ngjmeguS/LrLpQTFmQaPWz2fHKpsxMc+/K
EHoyoQD/HslHiyPlmJojyJUXgA+HkLYJnIvSvHo5DvNIDv83qYKs+qVv7ts85kdp
MEu5eek1xDm+KZnGHKa8mf+2ylhcSuYBlDfc6atW2YbXyxOHjUKrKNfE5yJJT/78
5UHcY8dznnR9s65Qh8pMWT39YhdEStkgNOt+ztEM39g/7uL+LFxk1/BwnPI+ek/U
4s1unydvkLO9bukeTOiJuIF0TlAfLteXt7xhE/F5wg5Il/yo0+/0G0CFLUYJemZI
yNy0K3fHbe8e4x//izUV+jmofv5hOUnHjmp9A5Ao/wEhBCc0AcUFwryHJXuuGT7V
nQD7RLq2SsnRTtF7zegTuoFFKAxQXsGbgIMg2s4J2EfWniw+e5nHfMlgl3WVvMDZ
7bzL+sz9AuWEMmYequRFgmgvs/q4u3L6js04zkQPJrL7Y2smZnEGV1i8ZJIJHSUB
FsAPf7Vp0zNuZcZNJUz3vAehIpXmQeF8HaAeyHVdjlqGzqLGZltNweliT0Negg43
uZvmoLyLzdGpLgtJmeA/ObRC4mZdsGEjPUOmf0HozOsPWGplwyMtD1+A3CzUr302
1Sa1TyEE5erdmwavTUsTjGlHBPtK13++JlZoNvoDoBmc3AZIY9Dwp9de5DANG9FZ
vg81liSDsRMW32O2F71BvdaY8HYn49H9pQ2AJ/cPU3kb+vnlTY559z7RahJKwWKV
HyDkrIVepQrI2v9qMDoPhw2PxYU0lR6LzAtHJOVINqdA20+vf42+cUCAr4knTB/K
f3nWJyBw4nq16YoNZjtRh5+d8D894zviYkxoiQrN5y5OOaKbR9rIYWTe49dIy+XT
qmmZwqQ+rrBdM6Jp/G9YwN9Hq2uoL5ytgeKiW3+kNcKvqHd6yUBLJintXCByE+yo
TiglBVPhJ0W1Yf5DIKG98VKarmoPi1iLrcL71+aHumx7j5WhWgVEly5DMgHEA4P+
qg9djH2PuiZrs6xxXECCp6LT/L7nQtOtAMzJqQer1faYl6qWV8Dv1tcNweyfSFgO
FNxIXmdKA9qDHu0tgalBYW+VN7axK1D8mT4nYPytgN2Z24jXDWNS4a0E/WoPMhtr
h+QDinPsmnXiX9BT+rcn4AHl0z6SNqlPoQkYZUMTbCJwZqOHW42MurXDsFLa8sek
Bbh6V1N8986MDC61s4g720S3aWY0Kn7UAKUiFQRNzs5hql5Lb9OByD1uIcpZC4JC
8PGJHYTsr/DYp1FKTj2be12Was3nx/4TfKJjUuKV7H9EpVYS7MSflgzqiyGDcrGS
Lb8lv9z3rzgw3DBcI6eD5RsQHrKwVgfYL7Dbniwyyf75wSpp5KeZxNtqcg37djY9
/JpC4He3dpQDVnukViEW3tZt3dR62WxiPEvrWPSjfyOY5MAW952cPUij7gUph172
CqX61ha2dviLvvQCiVy6K2oonFK3r1ZVDbqNovfnLre1B3grj24D7Dx0jYdygMEL
1pOdbej/RNsKWIrI/W6cMEj6R67bnchPhiA7Tk/LIW1R+QzQAeBhgdm6BtpxVqo8
PpYUzkoxrLm9hpkXZVnPvboL+vi4YN0HVoBVDF8BpB8pAs5/R+q9173lLub4fLHJ
CL1Q3w3nTz2bySmBe6MW5fFKUglkmpIJsCc/eXZUqePJgnuBkMIh2Pt3uAGB395/
2lIw5HtedKwhJKtxHQwn3qEo2dVe2c3vrZEZ8szAZoBlt3BHGPlvCO3IL96qxzQF
mocbNVpDOoI8N0+WUuOkTDTGYqkIdtOrJidgF4PBio0D9GD+5BjHtdPbsMZg1m55
WisY16G5zoRd1gtdqy49Q6EZII+LQjuC52Iok4kQk65vuXVaeprnyLZe3E/YJumT
ezkSAvuG2WrTJcOPkZkawPZEy2+NAgji62P0Quz7Lnjab8fY+PTRMds4RkgE3KfB
hqyqY725FvYXbUw3NQNP/K32DtjGbynxjgUwOwiPi2vLAI+stM3UKz0eVCtN57Sv
sC0uSgb/qnfGGQgrdO2RUdJjg0AScPVrakAq3Vlx7fJh1u8JAHp4b8wuI5IqoddK
bGQzjQT17+WAtDMpRiVCM5TUWPtmDj4X/h5mGhPSxi18zxc9Ygzv40rkpGSuyQDy
NJ1x1K2BAVKDA/TC70VmdzBBeld2Zl1ZMVa4NvQCg9UQ65ZGKwIrdLu8JwhBy7t+
02d6qEOIQpRLDJ7nHR048Yld7Td36VWq38WCeQhkXB93p/hLrmpZtdQH3eicKmXU
dysMcq7EfAH25yujh+hYrk/GPjWd/9ROaJxcbXTjO+2N091spf5imYMoLFjO8cBX
UmWzCTqSrUCgh+483JkGjs/EUdtKwIltZvVQrlbiUDLNNw7m+OyyGv6F+8uh9uwU
vRv0Y3rbtU4QT+T0DFdI/v3nwy2hJ3m+MCajhPuCxKthU2sTwWdWFExga6Qd/WeY
TY9BwE+MrdlGrsyGPVlB3MZeSWDwk3LjZe67uAFULRCiuoE8pYx2efKIu7JZSWsM
4gApbUeUeV0/q2rX3smgDu82pcjvpywIZ+EMXd6I/AZedjnWHsCV3vH6QalAR1WL
L7DCm1GSXhK0osbWQQRNLPvf1Ea3zzsnkRFTCCLR1uWFfb+x/H5oIskAgUmgHRxj
uXfLwvsfbrQ+5lu/YJJ427qhJH+iGseE54RaomYwDsi4f4B4uWPg77JrQyn5W4O1
f8Mhc6Ds/K8jni8tlbV1FaYIzZOyxVC0wv7zwd2dXIFv8hRp3ZWwHdjaBvDEBQMB
2edBsKqunhrtxTWCxvXSPEkwg+jumww2TUzQMsiGOVQkxxrJ2Gq4BRkRtK0MtYyg
xMxcY1l+OOXpAV1MBFuap3cFp5v3Wi1uePQYGkfQ/3OdCEvruB5IBbuiV1SzhPvT
aX0Azl7iqwocOw0yLdnMG8e+TSS3SPdhyAlmfYB6ZuRrRNB+VzdsQ83DH/zxVjcD
eY8Q314sItQ1EqxaYjJAFyJnsOYYdsT0wjT60Cuxt6qi6gyx6gfE6wHlv8ceb03V
m9+vzx7cwdbe1gu3gQKgVt2ulbjl0rvMFBH5vhXzwj5j5gPbdE5+XCuRg8PyVcBa
GHBJcBWYYCpX0swcr56cDim8Tq3uyUeKWU/VGPlo+IpXjmUDmj8UdDcF5uZLvPG6
Q5cVCQfGccqrNKdqJgnd4gpjQ7ASjxyQ3bSDruyGtH+og3TLZ6SigTa6kIDhHyxn
a9TDogj4CndUGM8gtJ8lWAimahtzRmMDsaQBGM9aqu7CZ2UwERSZHx9mWIqVmYOb
dfDTvSAM2A9YGp8AnduOgjY0FhKJJnEJ//ZpjJcA1SlImi8nZB/ZpV9dUFIBjDDN
rA/XTPqAcqQGZsDSDh4Lcynho7bgD+BjWKdOMZiA2US3o5EeeeKFZh0C/sMWIH3x
5liID+ykPoGbXKtsvwVOBwJQHFwMWa/8vKFnS33gRpE0lnC4ppQhlb7BasQtAiMy
c8ePArViMpH+Zx9mDcagADVatJvy66oZr08u/z+7LVcFZwXIb9fMkfYg4GVUwdo1
hywFBFHx6aZ2wamcTSGP93oPAazVzRlTB0Q3GReHYmE989ltLeBDuMKEY0PrCIuT
Y1X1nIiWTq4/zboayaNJITSnURkye4QkiSkKJ35r9Xiso1sgIVZBqpQcPlLCbYcx
67WOECrJvCSzjaPHSeWgTFguhyQ5kOpjj0Mc33poMp26MtCaxvilHk7Ap+lXexnZ
jZsI6H6kJ9oJZNzd9SDwI4AN79i8TkP1mFUYqibmsMmbwM5ZVa13C6eGNKo9YWYb
KTwlUR5KeNNdVT40NcdVzz3KpXxwbEXvAg/jLc1nxFIBCV3LOUgnIFYZYJDKV/gQ
S35UvTgghy/l32ycXFd/M11DILh1AYGizwx+ICMbp4qvt4FGVlqnPrU1GbkrwC+k
glD/fyiYkUVL5kP8jZldsdrWT7EOBt3YSh5MryUlLCo8yZ9ADd59dRz98j19tjJf
+wxFDJovM5/vs/50A0WKj0Autf59RXkd3ioMgTZ3RK+7Cwu/3Izg17dNvokmQA0y
jGKno4VDXqS8iLQDjKQOzxcE31yXkAGlOOduoCTZVKUBmTJ4aq5QZB8UHD4DxmMb
kXttdyOgQqKKTRdgJIhnuhMsb/zAQGYMrw+HTTgzvYh3VljDToxIBsCWKwT6cukr
YigFHokytscBQfzP3cmajldvijU6OI2pIhMk+BEPWe4nTNnn6C3/4zsPXRSNQNqL
wJ2dIgp6PBlXyCkJHrvMW9zT/fsVpCVQO4ivo4U45bchBU05Ux5SKCF7owPJomHT
4o1It3cRDcVAXJwQR3wUmjGhcVqNUxH/Gw+VK4L+HGUg0y8cb4pDf/Y2w/CIZBXY
g9YKCdZVkAFrUiSf8KgGyxBA2WIoqbjraL4qcdX8WnuE2AqjbdiBPZwUzHyI/YK9
bRNae19PhG+XL/odtN+mSI3G1m8U5Sv0rzi+rJ1lFzsCW5L0bMLtvB2E/uc3Bd2o
WRBGgL6duM9GeEdlcVDQ/Ro3XPLe3HlOuFXrrkJLlzVriKOYx366tBUEJsj2zznz
k/fIM/9tenV3LZH6AIAvBkYGRPXtEGus33Kh7q7UhIUSKcO8CLnKSFuLoHcy8WJz
ydenC7IJpGYrr4pzU8Fl2nN/EAYz+eOCgLP23dizpVOg6bvKLB5aFMTZSfK19GDh
euzUDcf1BP5lbNgLk6X9AZaW/zaDJIfvqZCry27FS3NH5wX9V+U09cpAmvr10zG1
Hl9PvUGUMPY2iod1BAfyr6hQBQLtOy9v3GJJAWqDzlFZzAQ4D9v4ljyhL68/b69g
5k0VGrv4fkLY6TI/tLujadl8psMMciqG8YJyKe3fMpIapRWJSG1s1qzRiKlFPVDc
1i8UgKEUwIemXmwMhpPs8hhgOlupwvy2L3U95i9AU7t+JaogGN4Wgu2pE1rgmvVA
U8OlRxOd9ZEtbPWCvqCvhiI6JhOEu2xvfZrVXoSk0pwaDTHZRBr+ObgkBZSqDiuL
kt08WXaM5QQyJmga9HiXmohMEPfFpzzGu5mP4vqFz2vhXKOuE8nohcC9pSic7fPp
aY99YAfJfwVnPzS0+EV8yWE/p2o6JRTOdck7KkjE34xwixMpluU5sPQNuDHZMgNC
s3f4jROXAtjCeYZghP0fbbVluh+G3hZVuhojsdTnkxHrY3SlNgWWkvqM4DKadZ4y
zotU+YS1MaKvcGY8lQkmuQE3LkXq223zJy/0ALGdNGPWNC1IX+uLL84jTL8yEZGE
Juqe4ooqbF9/oycB/T1j9pKjjHjCSLFmrfdZ/hcyyFsDNJ1ejPtiG1paCTnWyGni
0+IRtLsil4YbjxJqA2GibkLSNJMsxywcKqQ09bBZQJ9ay2EblVR1pJWBGW2XEcTk
KnyI9IUBgCgxOgu/Z2+Oh2LUYHK+LaLTdpDCNoFtzUDnXXjubSxQXrXUupnkSz8v
luUuEB2oVCdvUv+26di5H048iZia+cBgr/ctFEUg4/kVWlpCmWoT9VpMjMhVNvA1
vSaRrs1EFPzRSDMRFchwW1zXUSqyb2u/HIWzutLhOf3LUBZONEjYconaR5BO7Lkl
lKjZBEKNQo/nZW7jsZTfNQln3J4Tvw7R35hXYrn4/Vd82hr4n9t+xnHGTPg8Lywm
VwODLwtAyCz8SYk4JtorFmDZ7Z2r51NULltvEsiYe6KTSY1gDlpJ1OvjAwtDnIn6
ZMm+VhlQhnKZz/OvNBjdimifoeYyFcBvzYB3EMIFuMz0DUiJth3kHDufMSLu9Pia
i9GqlNFAsf0dvDCL4QqN82Rhs2sMNPniMkKfNHC4jmUjMD5uE2LGZ9rcjhreHRzw
LVeT8qk0ADDRrDxF8hdG5LDCgDVNW68qmJUsrLFFNDkiKz3DAqP+TZ1MipMccwmJ
NbLEVQxjwbXE/ZJUMRAwte/iNOmfsjZrx380fj5dBf6inb7BXINlcBUWTA/PJAN/
CSQ4YxzbWusZEuiD4blhTXvNElzrqJs68aUZDcAXNs3S7LVVlyraAGC4SSIuItRO
aJ8Gh38qxkETiInLfeQsd8ZOzgVSKLGgt2IvTjnqvLNjHfORpUnPQt9llt8DuNuI
O26XvvPOxAYIgtC9uqFuVFDKHF1gmpttLlxa/Flsg++KDPuwhI1H6R+vYEOfKAsS
jWPmeYmysWi4YZWs2cmjBkIv71gKN++bFmfkRwbI6UHQP11Ugo+0agm5O5KKl/n/
PiZVSm1tC+wNA9lA4Ie/TPB/1uJld65AQYd2M4MMoADTEIMupmBvsN17cO9PAHSQ
yrUe/kEji5k9Kts4Eht09l3Ok1h4sRdyi1c5B+UV46x9snIwWaJ1uy6XFHsbT8Fj
W97XEq+O0tYvAd79DQA4uGu5dn3LkWj3FSao1tsLV62KjWmseeXamF+yymfZzsbC
osfQ7hL28SwlheAupZoVorkq3aJpLIYfJ/gPaVoLXGuf2JBMFxcBdj7PRSqMrur9
nv8j/aRCA2uhlD2EARtBuGugszZGxzhZFc52WEA1pVHukGSLz7ttHzfwkWSwkpY1
h6/P34/saDoG0/LPYsYvvBmJc2NSaMh0qHdyr6nxfQMKBjVfdFeYD3JTexR63Uwb
W9TjI5vfDP3du3epcYdtfJQvNM8b3avbFEXu7evHDA2tfluRVs2K8Jci7EIa/RZI
gndbivMAfgp5Wl4A2eexJN87QX0+9F3bE2XLqqAtLWqWhVTX71Y9qn9DkWOoZGT/
6Q/D3KaomXNi2nu54qtPWzip8hFsJ9SV3Sq/DbfoXEhE1e/eY8v7Ghceavc/wqLr
kaGuUuwYouYEE2ra8PlIwXiz+GB/HQ4K9JoBWygmM/S71u/J+iXhW3aCDKQl4ytG
d0CWeHcI58qU1N28dwuLnqhw1mqFA37VYRYwP0MgV1vSqQD4B7YvFdYGRIBRQS6m
hu+AWoJOKjYCr6XtDI5/UlWZqI1N+/2bEmzBs57s5aAZWwSyIAstyuKJQFBhNSYS
Ot9pWApD/pipwkX/sOj955VmzrRHv1glum18I6dfRQuFbv/otRBAQLJWOu+cQs+H
IBhAYJ1FbYxBlrUQneV0HlmJ3gvqVB58cCDDPHGIR9Fe1immWiGdKf5hIDYLtwTX
TXpkn4uVHzI8Y4NA9EKIuDOozMNll9AahoQJPh8gT8IZTPA0bdRMXeBG0jKPp+aO
3xWPfUJx7kJ8h+ZmfAIKxhzBz0d/XaAH9FYtCFAB5p1S4+Wso6Bem2yuDxmqRU7G
dFs4vWhtVEhRMPwnlIfHeu+bztn54PWvxKFlCaOO66UpzuWk8p30DuLxgd1uHKk2
vJq7J59UeiRQAskeBgf5cJR/GulLSUiSwaHg7+oOIplYc0TirKIsuPd9q7iKEEZA
vrzzsBEFsk0MHOa7zB6obX8OTyP6VM55txTIA8fa5KDHjq6541UqUZbBAYZHg+ZY
BlA+EwBaSabUpOUGm3DWhPaTS4ZBIk0xJ4uT4heXA1o+q5F/cEsKV+BOxsG2tJoA
aWoOq2x8XeA8TtW2U+AeuBhJHjyV81rwvY07IokUiTv1zKsrMl/cue94xWRsxjcc
ZMKmmWhfVDAySvPVa/pYDMmpZgBfg9mDfy96ka+fW5Jj1a3FBW/5K2zDxe8z7wjL
UFIIok8qGa9V7Dg9x8+mRugpLl9IZOIKDeiNWlUxOX2aRmsH4p6k0EoUv2QDq6J3
2FtLeCfqs+TZj3avj+eoKs/NYEtT5M+Sq507hvEyxUIaZTz7uLRWhf7uf5OjngS/
8wPJxISSsZpNlEjE5QEsFZrBfItE7MjSd9uH2QuGtq6CI0uEWpobDrCo5bhf23Nr
pLqHmTnMVwl6DIRZuGDD1koG2VaS5HkTDoOdNn+nGlEiFcpy+tW5f8hv1QVE53ri
zp/oNLa/OyD+TSFJQdMtFlAejD2pGJxtMrLZSXsKv5JbBji8WB1fYFmhQmNZ/SiF
yijV68AHIZfJJ5n7PIUX6cZfU7iQDjh3dE1hiqToH6eAUy/fDPySNVTxHGqnZNpY
A2HCKrtzEn1DJp8rLTAjLxUlTvoTwET//WoukZvILCumQ61zHXH5U7H/stdCgAyI
6398/ZzonDmVffYU/AS3+YmTgvQoEENHw8xiIqVYbTQ5z+3/6809kW3y5KNhlwVT
rAhwhel0H1LsA7H8PAVSp+eX9LFGbwilIlOJWcdkQxepGKuKGQaR2py+JwLjqsFR
xcV/zkb6YFe7Fgm30Ne+FhIUwgNbibn8XDEG73OCzsOo7a5E7tp9HmTDUTyQkwKQ
16X1BkFEgeaMGQfvGp0ZF7xXT3pf3zhlzE22VynUXVj9tOLW8bN+AenJXUmUceZX
rR+zvHFoaZECyokIsmLip4R95MCVXtP3p8ui4XpIat+MVe2r62abCqsbC9W7g2QB
mRG4V2NvHhibak6CyqF88YXi0MxCB/he1GUSbVYaBh4cu/LX7pX4MJVfPp1Azx6p
J6gswgYqzGFVXsAnX0rb5fxc7qCzaTIEkr1lc0jZYiKsv9u7sPRJubkghZgklO/u
f/07/V2shDE8lfG/i4zD240wr59ra1bQyuzIg95LKJ7tQf+MVd5k1foh4FWdzI9d
TP8084UxpWXlqbhK2u2AH5tTkjZDSMLycUpgkKDRO9l+1TPsPIpjJXdtmOzKe8ng
6J8FH5fWok1u7f3G0wKSdKPEFC4DdcczYDqj2zd8ewVFbjh8yd122p6p+XDQuqYm
eq1lYbUCSoAEvv+RmP0tSMrrawv58M4OGw9qGKCjpA0K+SxCUrqR3RkFV71V9/+Y
GHqSPN8yZdshmnTGwvpkXmivupAHeVbJqzcKDXx+sIr6rxZUQdOQNwc6p/4pQRgg
UOnH/zhnSxX4vaEE0RvzKDXvzU33aNzmTHZVba91+nAqiJXOVycorS85EkJL2CMt
k9RxBJMU3FCOKu6VnS5pdR54DK4VCCe+H5yzeaFtQN0XJwuhDykmyf7yisFMUKyK
rch+IfBsb/r62QwrT0roKh5jheSDYN5+RFlluwsdkcTADtyjfHDiUELQNbolXoq6
GyyiTpcZ/Z+A/Nqdm7ayHb3d6a55wK/+ANfQAbmKdAVllsktUmfSYyfzlEYESduu
qmyktlSs/evUGALWnU2q6QSeXF1mwy4YWYZimX6YR+lw0mM1WTp6z9GEvaE+3875
hTU/eEOcXtPVDxBShjo2k6/BtHcijCGm5AOLKkUB5qN9xahWWJ7pQ/+4DS/uPWb3
M5J6UpNXJlSmZIzUWktvru1fINmWQAhxsnhW5YRh4QfalFLSroKSzkDqih3kkCUi
eAQMHhWPAgFm1hhY0CtXmu9Axv4JYyo4vbdGPK0OqVgdCgIUd4810pLvZzh8CYT0
Y1JzLYn8TGzWh4fy+L39u2MF7x4J1kDc+oloWJIFylDu9Ww+WWw/1lh2f+qKT5dC
FxkzgnzFxDa+0nzID/DYp8iILLn7e1cY/2TUmA7DydNG7MUM1Sq2W//58MbAvazp
qF+YkyRHczhkYOMnHX11WAnfzp47CFXbjHavcmSyGfbvca9EByiQONX7lVsDODOj
hZp+6Ux27xYoespfSIKEsfmW7YCDejoqXgFPlesJaY1nP4zz2W7p6Tvuw8p1Honc
VxIvo80C4r9qM1SV29GT8mZQ7YlaSHdpN2tCUlZ1Kj1sJQV/W9fvUpOQj4fkFjiV
K1wOYP79vcsBhF/trnTq3wseEPQFI7a0w0/AHine28oT25Z8W5adzNDCWausks8e
jklcmov7cWAphKarBnVVFeM/Sw4+1MjicwnBQDkW6RXnY6nSHaY+6uY0mLupJh6U
QRpqGjxtfxw+M3chWzlExdGBWvIM4w2PrxBNBJn1DPeSy0cUeiN+6VQ+44KjYOeC
1zEPAPypeQeoNF8CYcDqZJiKjdEqeeqXSiBsa5CAIH+j9gG+bJoTv2+FQPz1NsA4
sUu/BKNfYhDoI2R7UCGDaRe0s6m77l6YNyz5iHPrgxcFGSWHhl4csct+HT9+vjhj
uXoqj97M6hkqkl3Ju8p6H/bJH++rP4RFmJ5YY8mONjiRM3VfsgHzUb8wNMHU2SSx
j0NxFCtDkq9WHqbLy2YKUaw8OB9Hwele0q5se/kuPISUJ+Y+XJgBWEtfWiU/dlR6
QAKAWhApFek7PjSERwwdCJJ5QuiUd2uePrYlgLuZYhMtHJ1B13C7P3QoBPQRfyAY
uUVQCGOI40Q702i7I85Aq952cYU7aX5awlmun7lq4mU+Eztb72y+gWWcAqHPT20N
YxSDz/1ln3IUYnBW9eLjeN0ZVtrBbnmZM/z/X1lAFmp+j7W9QFoOXqzTyNAdsrRp
vRwSkoyAfs82Sb4q36Nn7LjPuvlKB0aBQkiYPXNEaZ33bPB3MS1TrkIZp62+kl58
qJpjNSZpliFoZmuoER9gegumhG65sNhLMuyE+DiUkU36JJ6TM8HYfgHMybD0jiN6
HZnFyccJgRYxvnHk3aDHgxpmB5u+dQMo08q1CnUMeSgQkuZkJo/ynsSHig9m82G5
G6MKm1HTxyn+/qSAOA9iRcJ456NOR68WDiTrdhnSbtumHlzM0rCHUlRD/am7IDJp
Pnb9pOit2eBfn+yLijWiRnqbJ7q2QlJt3pCGtoLjpwnSKN6qVehNipAUoYappzW6
BLvYl71ci6QrDnGMApju0QyylDtaD4l/uGzpSbKpGIpM+fGJ2m1nNrFDAlkxiMLn
Xs9xVEjkKgbQ0eJEi3HUGcB0zt8tKuz6QnbvL5fR0txcYddHOXU7yyJi52yQbtIm
yjMOOcyqh1ZNmtX+uzIstUEiRo+Nc8DabSfJA6RffhfTaXa8RKsUVT49OA8QyY1P
Vnr5kx5KQeH7W02HQXzIz60EtMI+GF11GSPFN411fDZ2vSeh4iL/9uv21W31mSHc
6sMFDk6TeERZjiICdS2ePzni2YuJS+T7RAFkl6kb3vnjpJH2rnSQHcIk14EbVn3z
csKikahg8s4/cm38IJSeqZ7XFNDdXiANVq+SSV42DC6jUHDKZ/KyoENvWPjWDcFK
WYwiyeyNhEk9mZHHTwAzt/6zP9izALfNnq+bfCIEMOPLpprb3eFEwFDemAEjucXL
6F6FcGOjXlRyt1l7m8yDE5Bl/BlwVWkn5tYOgj/orx4VXjwX74NNzN86rOp2uHqk
j9KZO5L/tPPMl9Zym5JZhSpDAEIp9PqNxi1MG9Jjt3ZHUsEdDAzk6KB56GttAp57
RO3ZjrUJUEp05Y7fJgBadV0PB6t9Xe+57S5HtNGodoKuWlwgcI7ZAdAQfghboSNi
XMYQM4v/LxtNLRtxlwqYRRgUAcuiXr5YvRZ73WoVbICPXswWPVnmUJDouba9oaF4
ORE+fS05dGLHlTRey1ZQOjEC6bMYHHPgmTFwrTv+n+f1kkKgr2HLjQdrexRAf5SC
UzwqsaBzOT+JWfKcRtlfhg6lnndnmm7vwOVqaaijcui2hXn/XtKbd1JEKEW2NYnH
WYI8JfU5KDZdGKK9juRIS1g/p98B9eHNjcr3VPWSqqUnfa2AAhfRkfgiseb1mOVR
tuQWkU1mC1GkzfFIGUPSxtK3R/ox6HQCPRrvtJEqb2/hudA7Esw/rzEG7M3ek3vc
ckwtAA4DBbw63ClScxX1vFNt9Ql4PCt842ewhx9dCnUhXDuZxSzLZ2jW2HswFbw1
8EPIjttfne3CodmJF/w0chjGgEgEsg/u8TzDCf7zmo/zek0jlhxYEUgDopZqKHpo
ydqDX8dcy2LiqsqorpxPrlGUiN60y/72bi+/gS3VQYIsjP15qxv098Wr0UMG+l7d
2Ls3588XYeP9fb/Rvg/4qEJq2LhYJFkWDWpGgDx0Njcfvx+9rL5lGIcwGJfgm8xW
v7rKrh+v4LEK91wNeBF+JqGQN/d/bt4hZcK+ZSK81uIspzHeuVy551PfImQaMOC6
Lc/7TkfR05P8oZxHSdXngQwls3H4/EM3Ul5UPOFOnyIRx9oKPA6pH1pudbsxbnyZ
ZxlSTqtrg1tIRchY/bT46n09pPHvrsMfjM50QrwaU6uaujDZDfuw+16Rav1vf72U
R8NZaxSVx6Xj2QbSQNDvjMjUUFv25NjQyqQRSZgvAA2ohPBJ+ROmnPnVRQOkMJAq
uMuMmNnizisoXCpcFJT0o2S8k4/BPauqXXJne2XsYCJc8n6IN+W0M8uymhuUWzIC
oMjlK8rX+4/2essB+7vPVccCG8OlNHJocXAS4I2qCPB9ObYArmeIAvo3iDiKq9HG
TTrr2LuOLaXVzQ3YuKdaWQl5w7dOjakCESz08f1IVdV6iYP47gp6Rbsu1M8lHwKI
cGojbpDMjHkHo7s8TQ8sI4d+sOkWCmKR+q+QbOzvtCn5147fIkTsGe/rW5EgaOHg
cS9PDZw3UnqvZ9KLA4aHUAHDaUXqhWojguQrvpw98WkEOS/S6VjYvhkNSPrvUyd/
VVnLFY58zBk3H+sfXoQaxWfQ5Q/nFelnPPLRpMwGDKOvqZr4S7vbjXtJSJdmShlC
i4+XSw3BfPveT9KAHDvGnTAqhk+5V/CqmsddAowWgfbw+ybYGBfs/8gnNmrvoqhv
YOZz3bMqZtvOND0YEGAQL0pgGT8/I4LKs2KdjlWxHgcRjLJh7ArvrQE97gU894H4
ovbILy4kxldCKaSTcEbo2rUhs49ppwzbysWaPdC4CIKdY7l4hW+rSnN0ltWhhaLM
I9Zx829mjhgGS0yJjwZHLkRefxsZscK66+6uCrTwjaXoAbhlbcwlbaCVszLdKURj
2u5ydKtU+kt0HIlVGX5ZUpj3kJe1pVYnWBtWV3q/L8MVCgG0ADKt8sGfcH472byG
Fua7VKBKj6TpEVpOfB6kaq3B2/2RpkmLBuW1Bns2RKwCqHXs2pNyw7JHA8g72U9h
hOKpUNplnZGzLciiRibHSZg8oLKL3xllkIXScEVdgTIrIzbotS40/AhwdhN8oAck
3pxavcJ+AtR42MjXmLhUarDtm1XUQ75r100vCxIvIYn+hRd/wmlmtS6A3j6VIc/4
guJD0lAHhDN8kxEfa/Uwlb6yxe19orN0rW8dCmiQnE0np66AFUdDKA5vWHoCIYti
Iy1xueTRoAno2hyGUdhxVOnrEzvFgUVKPQQjSqoiVEJXBuJedxbRO4LuubSyNgsp
+qGw+opUgGJaIXRn9gZB5aRAd1mnAIug4308QqW4YxdvBYqn/H7SdR517ldxaLmD
f3PMiEAYuBb7HSDB1sNAN53on8p5rf/OQmHeV/3VsWz57gMaEX78vthkNIm5LoPF
rbyn+QIbT6h2Ka/PiD7SIdJktVTMNMKxaG0La0hLjqmLRn1LX0lra1+W6rONRX1C
eVPiTlRlAPLTKxBbXFkl+O1dpPqc3lae/etv47uLMHeOYRw5f3ag4TOy7gahUbti
ZogiIxGfWNanKT0jgcZlK7f9vMmMQsQaFWM1csbvU3mZ89hr10crFtqJ+KvCzZAU
9t/zOcsWWdTzR+JuqApSrvSe+f7MHzwO8ZEM9YotTb10dHysuAXY/7sYCo9S/iKK
9ptBaazQz83uOMowKyVFG/vgsRphYeTPD+OqLb0W5an6bF+ZLbSy1zxln8ZBzVjx
60b3fiErleeMgwJrT7q5oxCOIYFg6gLJvmeURzXZFmeOCfV50cw8aWMoeiC6rSFN
ngY5cm/PmVu8DVleniiK0jvETAFmxcELy7qxpmtP+QV1CsfcAU/OVCrBdzGwSnRp
TiGK3WxijQ4p2kylOFx/0uyJZUAbHamMJWN2KZB+cfbPntAqGNvPagvwjzuBL9Oz
qFfUN7aIUHK0lJwxuNQqoVbmMm5mSXbR2HqTbqPRlcUF2VuMycTmdRjAxHTwQXHF
aQhSYlVloxTqZ+vdEfYCXq+/+7uRO7yLBSnnq7l28UdV0gum3DtCDcL7squVRWBs
Fa5kJI0jtltswa7YvwyfCwwLvVW6j4Ut0xKy7GwrpXBc2bWFbfUVAASfY8pcaChO
IjSrH0dmv7+T5zAd2zdEuvkRIXuYfnY8Z3x8HpzJrqWDT346UKUGjIjD2q532Qi9
MwFH7k9s2Bpr+ktqHPeUXC9FdavPZvY5Pgohr+RGShZ/jG7fL2nYHg3qIbgb9Rfp
9RTzo/DRt2/MEXIj430utWKpQAFDislcPRv4/oaWY8Krq5NKHWk20rYY9kYe+r9i
h9M6mny55qrD+nZu5b2mPb1fsPHLGBOwwry7V6aFx4kZBY3gidbnEJ3e+iT63lSt
zjPtrfJRN5Zwq2GrZitWwXrD7C96HYhCjJeqGPOytcA/WyXPDqeEQhkwJ21pP//N
SiQEWQ4X/kXwnh3zzDKj7Et+uZbUWqgF9HKbg9iwnfUrkxQrRY1nomzuItQJDIfs
4Tudwd2WM+8n8Emhn0sK+mEG9EhxcYJJcYiy0/Jrg3i1xNDORr5cpWFkCfXgxILw
xPpetLUsZ9vMwaFYbMdKB+wOcA8CW0ppsWRNG3i6bUvRB9fx6iNU43OEXPKNRXR4
E6sShKTVJtw6u5TWXEtNWMEuLIcbQzTtk6813AebRI4qzS7K2YJRLTixSzmpfYAG
jC2ZcRm9e6H83t4YaUeNEjLeNQZ6dMM4BiohY0XOiomi7SXFl6EsPFYLz7sxm+U9
OS4r3a6LIqSx/KBeMWeYC/D8nHc29F/3WbTfgMH+zGFxX68HIvPtSDaD5lnbaPIV
tYaByU0MTIURztwm0nBYuygUW6ZEPY2ZgkL1GZsVHOKQcX8DutwdgAVGJMjZGAqh
1BmI8CYto5OQu12CIrg5S6P2OmgbUgVzEohALzduIncbljX93wQ0F4P2csaLGxQe
mdWJ6ZgVmYboKCiGbD6M/C5t/G1hiJ4PhfRzMtJ98AHe6nLllaiF6bk5GxVPo3RN
CM+jpH07zFqTlZvnp2IWRF4dwNV3l9pV8hKjDPfc9bMWi5HZmYa2j39l5g0/o963
f7saqmibowrNeJwCv94ndHw+My5XYGeETDBBBFdtl75FD5GuXI6zsOFJNbpN/Daj
vOHuVqfcw+XYIMDJnRu2axD+OByi4MqScqC1sOiIZKIhDplFbwLb8hpwbExCYbe1
rdWOSW3qPwIe8BSUiO6LutL+hnztUTgEgCNfU1dnFzsGtYRwa7Pz/rdnJ8w5xBog
CHzoS7RrOYb+13rsvTOLtWJCRFUTW/qLbc4FlXm2XBYe1KR9pH+Qm/P4Xqb7nl9a
fuawPxYK11hyUWc0T/Acve/RAllKkTHt5eUQuRj4sNnaIIXi4jacWcK7ZO1PbXDn
+CFoMSAjdPBLMN4ziMq6YcNjCJVxabCpa9TZCHOdgLtQp8tToh8+cIS7H7DEyZnA
GCIyrW1iLGp0fav++htyuYNpJVQdR4jHqjTLIAiisv5pH3iSM3HIqUE+kFOeQ5IX
P2CpIEOoCPGfT90ZbGdHSET/k6GU6AoR59EdWxN2xAC5+lTILagEWQMJNPeo5TOV
zP1RrLzGJogIp19S1SzX2h/uEKwpBYkkY9875wjPFWH4g7jLIMc5UGF+6QQ+6Zv+
CJX81YxHVBm+prxXAnc+m1/FVW40P0PRDU0ZfOTV/uDVfg0aaFJjilavT5HuYOlV
7Ngkk7wXdwscGBdseN9DprQYAf4qVAljYstf3D4SK/Q7RsjEkDGpMeRrZJxMeUzV
2FyOokw7a8yeYolQ/g3EEKidYjsRpMquEvMSQTUCo7I7OE5f96dv/QuReVYMZvGc
rFFXnfOtyQ6mnA0BY4mr6xKKMi49KTc8eFZjluRHsX0edkS3uu2SQYcsiHmQRMtT
DnV4m0zsxciRwpiVeMQCZBdwvag0pptfhRSy1HLViwEw1DZ6PhFnyl3CATYW5Ab8
ZSQ0nS8dBvLFGAkxl3xXdvk2kJaGcfY6AgJ6o1r0H59RD0HUycXqoeqeIssX300Y
52AATrBJiPxXGGkU/iKNhgUeDkQWeoaQNU02R34swzLo/seTlLB/URNUAbk9RiH9
VQuLFF8b44WzIcjT2xEv5QOOLvSQyybwtN38AZ5OSEg6Gry0lXNhLwVCSJ7H5AQn
Or0wthf0H05BLmUHSCqE1jWFZEEGLjNx2extW6JdtY4xfSW7nXnspKJimIgnwbnL
yLpUHEt7RKNa9CTorP0JNm+g6GAPosEOrhWbt7R5QfzDqhHfuIp6wI4a6PUsk/2V
TggmebQrT5VoXjgzGUVMSifiyPL6kxW4hbg9vSzkbDMoTf7n/mGJp666YAL9rmLm
3uXJPm5Qm2LBhCTX9mNZov35WXUkL43FomWB8QwhMAU9x8pVU0RBcu5M3IAfb+vw
RmyuFGiamu36ZRn52a8sSQzBBwaEaeIDItvz1MztZeTYgIdGhFMtHEwo6E0+HZ+9
Umc8t+s9gTERq2guah0IMvviIN4rhKRsEOaPFnhsgDTzRaqxSJQhWFl/9fuPMjfx
CQm3BRzzxGXn51DreZwmMA6cZ3nwn00nwQYR88h4e/HZAhszFnzMleeD9UJmTLoi
CSXkIRa/IvpCy70AGCIJjJ9hbEWrXfg2Chg3jHneIdfBtlLkahctfWngxgfAqLsM
vvho924S0RuPLTPoivW+H37N+y7NYMb2bJsUMsE44YRNMMkkhqrV0neWDHj7e7PP
woCIAX7agSRGfk7uwliBk9F/mDwfC64EuMVU+IorTedzPJMP1GOYzjhqImFki5Je
f1MspQCOHkqLc20hpv/GNnSrEL/gYdpnkD5prbtnYIT6vcA0lrvXL3CjsjjW0pkp
n2NEOV1ov1WMMz2+A6gdladNqOqfchExgtxwYyLw3bg9HEHWhBz+/t6wno6F12u1
51xNwcGlJTqfs93xvK5nM11bqr6k5h/h8x1b/i+1Q/qUUDDc/wu4ykT6L5U683k2
iK5BCX0lKf6UXFMaGVTlsx9fNOj41CkAGsxGCb/Q8IK7DMlnNROSzPfRR8SYnDT5
5bP7GZy7jB2L8/dVE55U32BvtMRcRktgQGa2cloD3KxXZtzYzOpR7oejtLpzTlsq
/Yy1WnGcZspXzcXBH/IvNOEGzWjjOp439629Gi4F/4TqAB79ASNQXlHi0om69WY8
Vlt6olk4/7UgB3Vo84ddGxiX1Ca9IQp4qsWVGwtRBzX3T/wFUU9iyZXfMnWe5Y23
jPmQCEk+qmY61RwyHotVGIo0B1gkOXyWCD6fe5d/Wpat4zRXhY4XJ8aHHaGNyJ7A
aRkXxaEivRUY0Se08xsKLUqbpjzuvvWSKRXN9HH0kyPv/jou/e5Djdff9xGyh6u7
mul+u+JbduzF4GOrT1z0R7xBZsOx2L/aRmQpfe2SqasMnq/a/uJjKh5pjioeknVX
2LU30vGy5x4XKVashHqsSp0S6Dto+3XULQsfAg+7Ca+NPCCn/9kU//qqmcKXEQEO
dNMXP4VKd9sLHNZGbuJzffz54FFLL0muGpCGZyAHkx9pM6xjPlQjG7YPneGfGCfe
zYDnBWImCvqTUMgCZmbV3qVNrT4evjY58VdEpU1vaczBlxURf9vRmTVDaeTaKapN
WnaB9WljPZNqBwum6/tdocrM09mmpruit67DIuEcf8WeAI/detGGHy+EYSyKluNl
3FuPDPLmttgySs/xWDUC4iutHo+t45xnmkrdHnCEiu4QAujBhCHCn+5f1fMpR6FH
41IM4Yyo0SeVNacB3ZQ2Uc/X386Lgixb/X77A4iLekUQX34BREW/Nz2Pd4T60zXY
+/5N03onp7NOLMwm2dmTRqu/XklxmFADdqcAcJddkEfMGXngRr/rl5SGu9ukmFwO
AOx8gwkfJjKCVPbstwKT/me/ISjuCVO3Nu9/0SkM7DLLw70mRGSQ+9xnL+pfCsJ9
A3QKzfqUOTGVWA2XnclH2uKswUq/HS3wl59W5sKcfTOlkDJi3YbP0pH/1i9HM2sI
SV3nCG/WwVXV/G3B91BYSJeZiOWHgvmeNZDp8BTQX5UpWu8fz+w1IjrwFZfqcrfu
gn0VF80VSjT3OWOza1DOjovQ3Y4Pzjze5P9BVHdY0uwcWlhNUayW8eFchvnHS5Er
wpqZOWFcqwftVdx4fJfHIZJvZYfSz0K/Za0MFedfRqELLTgXLy5JKyVYqtQoh09T
2nyNkLMCn8e0/pmX7YzNBfoyx8GbQj3ULdQ6p8nUaSFlBrgh5XfmxfLRB27F8tcG
TEsUiPcACZtwSxXocq+XukO8xyRc2VljJ2vEubG4qYB4mJw/Jq/WOa3rcghdDxq7
3LILDUYHNCj0jYp3BPy9zmh6mosIBjlmh6uZdZMsBEfyfVL+0ghR1LPpiPeixzmu
89np6C/YXUfxtI2m/8okPurVMe7oI3Cj6raU0IIoqbUZl3ynbg5N6f8iKqVKe7LA
L1mkfrxlp21kK/HNuqe4tWcHREp6SKIalO+uyoNq8c7btXqJ6phnXQ8LKePZxT0A
W6MvcvsCtlO1kNqWSQ/7znEJxF/BzRiFexTx+IZLYEZGWpB6rZv7XnUdhMe7Ry2S
JlwREOZMVSb7le2s7QXTivqphEt9QypcykVLz5Iga2FxAJ4G+FAbtRLph1BKMfVU
nSszujxKiX0XsMlfo9AvveQD9INGIPiWNr+K5qh9o0AGaT9Dzf9VFdtA/qHRi5BX
xHa/nDfJ5lhHGHku/ra91B0W4fkjjZgt4NvE8E4oYeNK9AQCzaOYxQ+ixzNXoMFy
BqaFa919XDiiMiTNvGYi/RvKDxDD95raxH3bvgUQWLeqHVNdvMQo0ml6hlKlx0EV
s67AdEYSMu+JWpa9LGbWMUTTBo75ehixRdMl/mfbzFlooASd21BAd0Ac35fhq0l6
APwrq5jl9fD7NcmIDwrIImmQUGBvJd7c8IgEDYUfpTV6LMgvOWi8D6BA9On7LXC7
d4DNopGiUTWCx8Rp4G9CxhhWAfntX0rQBhUXFlWRBQ/rj/UXKET2xS06uPApcusY
FQMDA0iSEFR1S2W+cF6EuTcDvv0czlhrRMpdRg5w/7gg6tEztCv9X55vb60tjcPI
pe6b1xGoPZoZdVFxMnk0mvSsoAo9Ty6Ztvn6qODvXtesoRUQ1i3feOyrT/9MomVV
Bbia7LKsVCtuYPlrtcjRCoWoXLLRxIIIoDX0/0u4Oe2g2l2bo1QHLiZ8MxU6yc4C
XNF0dOcWVmngW6nYNqhCheo7doNV5yKD2SqEKPc53litUP4P6CvyUWS3EYbf6+RS
VBLpXmGMB5KlMppnb6eqjHcGIy9pFLVLfWWTeewaKs29qdWQtgfqGCkttpGvrrR1
U86JAxjqYqTBsAha7hJxHkEP9jSbEyAIO01EkkWPOBFdsVhNUG4KH9xNNQORXdNe
zFpu9x6P78gZ1O90YTPUm6Coj3semcvuwhgTWm5feyrPsy2Sx2RiYOANYGOVF8Di
/Rq4nIf9wNYzdbNWZt5nK9P2zNnGTa/VBN5zdAtGEXCnyUVp0jkF0bhjq7hsq8AY
7bLqZ+3AkIoZC4wQw/WoE9WW2GYiDqBKh7VmaosjprV4MdjpDIMW1h9GdWtqxVPv
Im0cLzPsuBukVn3pCc5UAlwObgdu4bYSDrebUq4uviFVYb+VXRt/yKttNBnQimQv
NYgO4BaBIX6UX6N1YKRoEutMo4ioovGO19nlGhoUVBqw05kKk/Cx4CZB2uHKgRYO
29m9k/n0w0BAhxDs/ECxxrcpTffHPL6KUffywfnb/Dl2dIp70D15UvfaJnfps4jw
+lqgjvwbHT7/73F2HPIO42xHEe6j95N9PS8AWxRWM6d2IKf+Kn5gUGhW3VM8ll1t
A7MgcBaGkG1CSRC49LCsa43EiVDiTZ0L7BrsrXiwjyqxz5Vcc+zvSp551OPgr854
mX+fO7/fQQsefBAobeLtzhk0j75KEmFzElt0D4+RoGwehgeFJ6XlauQYel08xGW6
sw91gXxnoFuGEpqwYU+1aoPqyBHVOfu+L83/+zcbIgMn86sDiUjmja2O++zWwEO0
aqu+YccexkMLYpZohsZWBqrPIsMLxcXzy/oKsZfbbM/CP1LIZdsqonmr3GQXLbSd
glFkwkYYXv5KzSEaugvxqxa6sY6N6cPJWycPqgklz9Pw67I8iR672zDqF7B7c5xm
R2Wm4lYxkWNiaUgezWftmyopKMYVjsBVRYO61q8mcU1Xx/+9c0h15KzUMF/auZ/f
oRuFZdEHbdUS7v7LGBZj9Wjbz+Haw6Mhqg1XiBKvtNj216hU6kxtuOXibm1bnqTC
PojqezGNGmeZWQh6uO03MZg8J6Z7RP0uURgvgDKX7T56eeh2fnEGNJRMBNhu28e4
H1sa3UtPY1VeG7YM1zrrhtZojA/aeZiIhdmu3TCU2O3doAjzwLnLyc+ZBjjYpRNQ
BQ5XvObrDG8mdCwmUWu4NBeQn1CzKKBJdZByCp2giriKjz+b2jyCJ7vdW5HDxA3L
vX60ukz2R1yYQ6+LXZOkWVpL8HYcZkZvVgr/owVMnvxY1dTU4tB4v0odPoCpcbsB
/+bKVFwtWMy7dc7LlA2A366szD0548IEE0UksRVnBj1WAXbJRLgOVJCjaAX74U6d
BqILqczSvS3IfH0dEh32o1VGQIoEQPHTHmfJ1gIgTqs//1rliPZs4RmueIa1JrtY
T8p8lNz8JpXH7YAyiGZG6kyfljN/jTbVtKMgXFPUjudkSnX5V6UhyI7yymwcuUiq
+20NKYdXkVhFQk86C0spP0HtBcH5fniYawvyWGY6FHhpXWYTEkkhar9i92kt9wnV
ciVXnB9ut2yr3jHNyteHJQpZWBE9gf1a7U7uUyfn5jrf2FePDYG7nqHYctU2THfK
8Z08ZfvaRZ/bUp07thKeif3Ez5E0tSkxWEaHntrrxfLdSxUniq0A505E2iLz+K0p
KLBDLzLTKbyVjcpWH9oMwYiKcmsGL5hAYv37Fxb6MrkS4OSynEsYU4qL/Mwubcut
mrtPpB3ylQnGtVP1ud2O7MUPdBYtax43LnEXYOVvSBX8MTQ0DSV1TkdMyuhKinZo
ibZSB6hR84j9chpjns0J4ewowE4QZ20pduimzM2AERKMCCQg6CdbEDwDzI/+uv1I
410KWFIQm5sr/f+H1bXLFMzqzBFrsTubnkMo4ha4nmMzRyce3i2uSkc+Gq49gJ96
lhbpqd/eXtHx9qpAX7aU6V0BNLtTjAfWyTp4JR/XQhKa4vyK4cGUOAuSnsDo+Vc1
XQa2IIlmRHQPKa6maGoIwP/nD2r+HtRAKp04Gpp1QQFNezCVMjhjEnps5RTxEiPn
Q30D9/Z8uYW2ZYNq6e8unwtWUiEkt3Tzpb1EY2+6Lx6fjbp0X4ueC5jSJgvxms0g
GxAJcUozrCKv2RB7Nm/M/uiVV32DwBfD81J0IEX/Yh5CpdfVzDEnjdZdIDVahzl7
1+vK8I2s1z36Kzcve91phlitAQWknL/qIOYBR4Ht/GRYSpKC9yjRjEQHYyCIvx1B
s2E1iQYo0aQSMfXjkg9p2pTmjO1659WKHMcPwr+6k7IHeO9Ns48GOs6RQWWxRVDb
c9w2osG2E856UPKnKizDfhuwogxIsIuRrMdCtwoFyRsDcZ6tpUiVP5uqfAInbXO+
BCknx4z0AGpE4U6z91/THkPPedh0S07Jg+/rye8os8xulYxIHAI091+a/kNL1yYn
dcLTrMzA5WqhpHxXsVUql/20x6O/CM19jv/LJRW010CysbUKm9FmKy0+FOvZsPeT
/Mbb+7FnLNsfF2+jVmgKydH2jWcPKpKnyqY9/H8v6TfTou2S2wO+fAskylC6vTNB
XJfA/TjdsPtF88y9wl/dZNJeAlMTpg6rk1MPgORvFPuRUpKKswv9/vZv7IFJbWbF
L4AfdrVt3KuImEIqo1lcgFAc3IyciIVIf79EIoXa62v+ug03mInD8ykdrcu/FdYW
lZFYCk2NBzwHI/vROvgp1EWHkB/K0vTAg/Ri6Sx7mgofPI4uQdu6vSPH28/hWGQK
4saFE47vl+JsPce8YtPuJuNRfEgExImYXe8pu9l/O9GPxO8VgeCQ+61KUL5vrM+Y
DmS8M5+4Kk4RD2+gDIQLMjUnb0PNnZl/mXyWz3SSqJO5kT8msDk4L6kYBL3DPG4D
T2aUiUXFQ/sbuaTSYB03Pr8GQeP9qDo4RabpDt+a486tuk2eg0E0iNoaxWOzB8rn
jvfO85/zaC36nES9TxIZY4OIzj+E33D+bAE2ZnxXMQv0f5Dux8/4ElT6yVoAaqHx
kRtlJRefw6Bnr6nZce5bWrHfuHKXrhoheuGJAqVWhfanIO7Fk2t0Yaz9ZLK/KPze
ZA05hYjvhlAZti2cGGcaHrLKgMQNaxNKkSJKtuYDRHN+gNeIIN7dnZtvFwPtBUDZ
NC2PHawPb/XAPWZuuDSYZlyfn6rBvgilI8FcOJJxeevwhlrqO4MD+8N7LSf0Ji2l
/TbXfi/qUEsMKvJZYq8XmkF6RbwnARXn/sYAHIP1xfbaDm4O0WSVMxNsNXtIT4JR
zjBfF46MTgeDfAt0JiUwyyeE+r4WWTFOG0oCDKxXSfmcWnhU8zMGSTqOojUagu6V
w7OMLrfA3HdO6/NfHy8dRO6X+zDe4OItpjSPZOHS+6Tj95rcpAR34+c5Kbcrm87a
7bx/Dd61L+hI5PaJzXxx/crbyGL8QScjFaLWnMK8Shwyc9tMb/2++CaCA3WHd0bN
pxDm7gLNur/MlYJO7pCWD0TZ8ugR4bCWDPXIKhjHAJpBl3DX3N+Jhq8nsROkFzn0
SPrUh4GImZbIG7gXflsHAdDooDIAA4K+NHloaOmqgHEU+3FFhy5G16uQfz0Ss9tq
XhV8M0CxOoPn7lAJZGQhw0hJmruSYNBFI6a3xj7Xo+SApDc4CR5AfIrC+kl1fVdl
cM/isR0PHwd2/HygU1hGCzJ4Npc9uLity+rczw/HxWLd3PVQ0p3p7Qy98QUzXbU8
JbeEHViHT/WcviC3tTOCsofFhMfqXpbv8uhT8VMqToTnJFfwwccdOMcjCoyx7esu
GszFqvcg2yuCFDABhLbwAUHh1Qj05kAuCULkKFZ9P9/TiaUxj3J0L1N7y8pjKxWO
9x4KPrmK2A2LBuHYdZfiVSuGvdekMzrQgJ5ctjiQMIEXCuB8vDvx7IY404ooImKC
tg9LnUy5sV6goEYy85qH0o05TJgVHDMv/d9mSkvOO2lyH46iu6IB8zzcASxUAlob
TER+YHHZ65xokxnpxbNoZTAmbNgcoNhUiwfvKpe3xKIOaBOiNR8hlr1jrcy8V0p+
d38qFnETB206ZdDAK1X9xCRyaO83Z0rkaSAG4++vQzDTs6mHjWwuqVHY+/LowbUt
ns84iW4ZRXdznC46kBHRIOkdtTsqbxn/HyAr4ipvRbO1AYoU2Fnj4FoH4w47VlEB
H4+okRVPvnq9K30ZsI2WbS9pr5TzP8Rn0H0xehExNFM5208Gz5fWY68ofBgI2k0S
b1qtce2j9+YoGyG3TBnQ/nNr8EykyiEOuvPNdT/nEP2OM74iAJ+ItAEeL8aBF6pd
HavQrRvmZr/tQiXVvatOqDfdCeaj7+wFMc2JkUF/rBqxTlj64NKICv75IC7Aeyk1
wwLItep41sToTJXo89eNpKV+9D+PyeqwqljK9dNRgGxdVkCng+XIcmzlvf8Ees37
YJXbDkXvXu7NXZ7vL11wNUcFJxkvfid2Sbl6AyKf3VJYpw/Ah/JnBd/58aKrwBFv
gsFkNvTHDpdeNP9XxoAj6Vcmavr35/0eLidS7XmW8mZJy2ykRN5Qk8MeCZ9P/zjs
fUWmJDcPa8A5pFMt65d2U5M04dRXz3zn6fN0gJUKdMvyN77bv4mL+a1QV5+wrdCq
KmHKda7dLVQ7op8MIt0NwVcbxYNFag3HZ6pB1gUcDDUVZZ7DgpGRp/oIkmbZ/L9X
l1ZU771ZZm4fanhYxxR6u+4uoqDBEx5VsJ8cZbpGm00BxauoymUZr9yjVxf/ftLB
Wd41WnJVDEO8UZrVXT7K05rV50fnRUD13gXn0q+QfK8DUajXJaUfzyyJBYxQG15P
mlmV38O3XgGaGuEy+nFadwzMJCGYiyDh8GnUETN+oXWVoSU7NGReHQ1LmZno2/et
K03Cy6wKU1V8jTxUG4synKQZP3llXmV8Krk6nl0yLsE5kReNUA26TSrHFC6HvQkA
s6+bGBLybDIMFJSAwbp0NwpG0EBeZROUSKuEl3jsulR3nCvNLeCDCLcRjabELtmT
isFi0B/QwqrsSDWsKHxAJVustzR7/s5Sagh3K6ehx/KtrZvdLQg+NjfkOkudte49
zYgsUfVFEZxK7PwUj3CZNp8QEjzhmomMQmPkQSJJ1d4+bQ3xgFlGORCgMAKgeV0M
YBKLNf4tr0jld6CqgJ4ROkda4KnLK8l+EkSIORL46+6Rc58cDCpDXT7uWUWgPvGf
8f+xeLHJDfD3WXMpnKI4te8eEljq2WvmHyHKz7U0W85cmKMCft+VzFn3kX0H1+IQ
PAq3K72JqywIZ2F0+uJLv4ddKqyvdXCq3UNZBRAg6KYb5ypWUOfD+hmdyZHmkSZt
KT9jmE5DqcWwGUfQJJDZeDkm/MHZjEw8mkl0T6SpSyO0kp65X9Z5mBFTRa0hFX6D
ZdXxUeGd1Wpe/AiqkOrDlXR3AdMEK0wl3slvGHlFLsA8boUNcNFnQEuDABfbfF4U
SQFI+Z7KICZ76rSj/4r6wyY9TYxMg1Djv2vUYDVYTC3QVEK/Gcdg1L0VAMml67sU
QTUCVUX7BfmHYcIzCpFYy94RF1nYq03dQqqvFBGaFAB2BPUzQ3GFB5vL0uUKYuiD
6zj7/u7tkyF5fToFz4mb6SFWiO9PuJ6P0RIz0hV/JVy1l4Ft4K3O/y8dLsk5GrIq
ZMMF7zb3L5xcMxu+SrAh7bxTsSO6A9LQ58/RIWxx2J3UVDPiP51D+soyYuBjQDyX
dGHIKyYE0qPpVzriKajaf0e2wHMl0IdmEyGSMowmpqJLS0E1sg3A9fEF0/Xawgn7
5wTe98NzdkMlP6YnD0E03RYDc0FfUPTIQ8z1d12e6XpoZ8B+82xZiggx8JgfzvFW
/EdQMWiPf6DLr3BgAap6Pf9DD4FAVMfn48IfFyvjo6qERnoFyRVp4jf4zFK+uRyQ
1iEeyUFCc8uWXkuIANwufXcedHZJrzStJT082YTRaLEZXTzugzRiWHbJgJyK+x1k
cq0D1vP459qrwZNM5jT3/RkG4wOxHqv9QkN8LSMNDdTMVT/19tiLJ0shFbVcVSYH
r8+8mxrhdZE9LWaraDvFXJL/cGHo3zbFZWuJt55w0ljYcX6O688u1Cc5pzwrpYSd
ILauT2PpwsY6G263Hy5xr0VxGaEGffb6fvLi8/rKPtZ6JY85azZd/bk8RXOio47i
72nRWyjbynR65mYrLW6e/yJlJZXH11O8VdNDahWIsiq8/Qa7NhZ324pWnbdMB4Ua
2tZhqde+wWfAR5Xelj6+7pL3iNn1N7aVe4VHu2x7PVR9iDX7dWoW6foLSGdZB3NV
oPw0zkJ4L1ToDUXAvWUx+9rb77IEqljmk82CGNOf+ZacmGHC/KegkpRZALm01HUn
hfq3+wGxKuXjRhSfYXvVwhCZbU/lsRD6juu1E+Vo5FZm+PpluGHYfn0RIxen4V8V
fcouH4oJ1+0GpyWlsHMAsWebxXvVL3zleWiLVqNS1yPRwPCjE+9JwcO+oZsCgRUw
4CqBh5AVG5TxCDpHS7Go2lRYZn/J6sXwmaqugSUkpjDqP8RRqwXvK/RQc2k7W5bP
Tth+LCxtzJMa21zEYVofqmASZH+a/C02pTAOYml2WtkGRwHr5AQgC65A4GH1nf22
s+kuXY+ewzVjiREMXjCeeeHn1IoETL35UPqVq4400OCt/gYRucH/e8ZTFm4Ob3s3
UNWO8u+3GGx1ThwShj8AaAfEMpS7PqZCSRs4lWBWvUVMbUo+MVtwGa4SVntv+tJw
5cwc6GANX828RHrAmqnL9nlZQMrkyCPvjg7xH0rZ6vnbaCEfbh0F1PdmpLvvcuQM
WsIxIuMVMt8Mn8nORhgMoPFmlRG8XMWtQLxbs9J2d7a4POqq7xWS+Umw9c2l8jim
PH5XbCtfnDYuynIR0gRK9WTjuppGaiZM+kVf81ZrqUnkkDMhteGF47G73/ij16nK
WgMqcOBzH6p5cC07xMLaKOgVIgjtkFd+j/R/+K2u3mjPpaPewWQiI99i6jcbLquk
WUgcTyf27G084Fvi+OMpcgPz8psCPuYyYDHQRs5RBaSwcGt7DytevWQLDOTlgg/o
xNfsOMjDEmw6qK8nRoPRrHqVsyxOG2cG0x9oOHsRFj9yHnBLyqC5TmPICc3jpQ9e
7uBsUQh9zGpofc8UuxTiLTcK7Ygp72ox61r4k1vx+TTfvZ98bWL7Y+0H58UV6sof
VBAqW+1h/pE+3aZrZAkqtJZVfgZ9S3gQAW3z5+KHiBr7lmaETw+tfXI4EYqYkhjl
snPkoAEE3wpycVbzpDMpmYOODWGUvyk5ebRuQpp0YPuB0RVyWELwFaq7IuDDVrg6
j9BhoNCivYS0lDlbiCJ/K8ul/gUTrBj0EahgZtB4PEIv/7q/ZrEOYutGmC+CNJaG
cWI6wK2XOi8L2eSP5CnBAhXD1YAIpOj0RFCgy3GlQpi6Q4rPD1Ba4PTLHEXKiOIh
xTXqwT6JjZJ1l0EXNTixR/CXsj4DaQv0dN8jZUKbhBIXECAN3KL7ltW5oEI5UTZN
h7jQwcrtNyKSs2DrMN36ya/NMFortsrEOue1YQulGwkMq9/i6tqwqY6rPb94mGpY
m/K/cHyXjcCVtIPYzm2l862n47HG5LRDx6dHGuLpBOzTD6K1Ez/lTQvVEbnfmjbv
I3wDgK9wu80wjoNglQqs8/IuLYhVGvo0/y1H2GXDjiz5kIRYFXQci+kp43mgIbCE
uZHR5J7XPwP759yFxNtcwaozN68Vq/sxTdKxub5Rf0n+zK4phv0J3uEKQaknFk/+
nQoYpHCCMHtQSz6joBNspuNrDLEyKjR2pbNX9otP03hj/Fa6FSE/o23bcLnVFhv/
OyExkVXjSit0Udzqy84Oahwc7XryM+m8VXZBpFeQ2noJCYnniU+UPUsDoabnL94s
NrwF38VN6YNUXRnb/TnA04nXmqqEgALJGmFmQ/myE6RyTnet5gpp+w3jdVFuOvC8
BCEeUVkncDu/vtLD5RoqatC1saC2ZeP+vigq8CsvuLlQIKmoxkYRgFajfRnYtL2R
qrL/zoPrLaloTWHm5QcBZI6Z8hRTcy1kW3NNzn8d4dhJMpFQ3ST8tD26zaNRPH+P
BIp9/1WSvaVL0R+yGWUhaVD81my56+B+ObvCA31fyClK/UkiWPwuwiKle8+lmuRZ
1XiARurLJtVaMH2auszY46WDb5SqfrZ28hI/jjsPUMbxzNNWLB+nNF4bFSmfaoQx
rtNU6S91Kv26l1Nmvlm7cfcEUfAyE1MbdHjXdWsPEW9mwcirvYvjAiUHEQWwu4YF
VbWtHgL6wH1jkwoRrn9nWnEZtlU5OLLmUdHgxVmzDL/gyhKcAfhn+O6PevCafH2Q
G2wWmJWvGJR6Woqt93/hg3WNh91cAlzqJJlJeDn8YUIA8S962kEFH7qNmI3Fsmp6
4FtxYRwO3FFSGwHbXthigAuNMQzGDwumpjcGAugq6eIqK07Jxd4/thm8OMPthEcX
nKVueDW/jsKlNH+2UjXbg+vEfAVP3QgjcuGx0B8IET2rsWvOq+rwGDv+DXQ/W0qk
0xRPdHo+k9zdG16DQiRnNAJaekVyGfvduRip5EVKqYycnAuq0rVHnPwG+Yw18fmI
/7o77A70BSlXd7YUaebLStGIiaBVB3F3FKRNn8dZ2FXj+ypQbuU6Pick9G18hJe3
c9zUNs34cQrXf0zcm0o9mdhybLU27GrIOxVJvnzHUc8K1Idr2jfe8QCtf1XCDwtx
h8aY/lnhqJOn9o/h61DRlBAiKoA6+WoSk3uhW2V9zSli2no8r36cCXYfbNBro/yO
XQKzMAhC6Ud0i596vipN4tROhcMmfVJQDMOoXrsA++VZ5K08537xhAoeY8WxYl43
oX0WlrfNbCTlq06n9mf0Zlg3tePqfTWBCx+XbPAu6pN45ND5J0dzis7KEvIMUtUL
a+s1pQxMdgKJvSLHf43mt7Uw4lRX75xZ2uVn5U8I+5Ect3Y+Gk6Q2brSSwXmTbUJ
lgrNrtcNDAsT1XbP8tZUFvnh2UO4DlRjAMKsNags2duvw43PGQ8IBTFZomSjCTvA
4U3+EfQJR1R9F2/QuDoARGyB7ge4HUJwtl5FslYoOOmb1GLVPPlfcKBUu2Nn6fjS
zpRiXApW3d3mjnbNeTglI3YHMYoBO0JKDgPITUO8UjdNDrFVpr0OQ62Z4gQNS6SD
XlZ8/IU8czWIV9IFJ4aUcunB0SM1DbGwuxnS4IGTSabTJXbPjSiXj9n0lvRUFE+G
Kh5ReWdiC+UOTNRFWsVBYeh+klSxWkuYHFW1Hukm2zoXkg6DVjLsCWBd+L47hgBp
I3frpfnAWaI7W1bQe21WJmGE28MSoiOBRogEcVHfDwq4kLGm1EXTCHMoAOOZ9xXQ
jxlBgeYpq6XnVjOWrzphlTN7K5GoWt7mgDGrQdjAuxF4SEPF5gI/MG5XvPPt/Gtx
EK3mhgg+s5LZ4g+LPJAzjudHcIzIKVMWmEYVyyMxY54sOe4oiAdLxZPAzc83J114
EEO2MROmTI0Vnf9EPeVUpMavIgZM11xbQ38KKe5tNXluhgM1fuQMrjjCNYALUTJ5
pIoYTyJsAmkLOHLKRU0keyWgvQYBZzy259OuM42TDVxL8IzV/dFyTnztn/9DUEAE
mca1Zw9p4ZXkzbv6RCr5s4fNvT4yKsexRB1xI6APn3YYqZc3hoAtTn0mWCIaqqx/
PmKmdm0zx1DDKt6J8jrDRSpBsR30qE0paO8quT8iqTa1q/+jRiWbk/Mo4kyMGUXT
uRwaGurpU0zpFbsIYrZcbgpk4rBGC2gtwzV4bQdozMF4AZ5Ga7QcmnYKftwejDnN
xMIyXinf/KO/7gCN1IDq3iBXbFfm6p7PskD1qH1wW9FjofCh0qKUcz8cJcVDJIKU
dD6swjqqn09cXhX0lCq+rm4VbX6qYbddCWMiEvFN7WIwW4hvf9domvMRM9khHBSS
jQX+RzGjskORGw2Zhdf0xnWPnqxSyF7mxhbEM9VnhUd6qpn7YVL/pt5AGAZVlmS9
AuCA6HjSTzDBpx1OtbSUybBO5tFHrDS1y6esE3WjKTdDJdyu4tIcHRn12Ckarf70
V2P2NwN3b1PyQieY3w+enZFd1Bl/jJ1HkEwxih+rL6bGxnNcOsKT6SX/aBqitefu
muR+BzOu1jaLAnp3kPlzAAXCfqkJ8EwgnBD3lkJQLErIJAeFA4v0w7vQ0ZCvm0Ru
PpXDnfdf+9ahNQljVFoJtJo+KfFAUghxySFBbiwrjfkHDGU3qsmO/zOkj7Or4MBU
Co++MY5fOaeeSHBhRR/CujmE+CbIlOA2L2f9HxCoKZpkMAnbZu/XLs0D2ujvBecf
5/Ijn3w+WRTCsCA7Dv4+eLX5dyLHOzuirCmYx/cg+JsvLttlbhwRFZ6zC5LIl5xr
YFGk7JsfF+Cf2yahh3rz3ouCI6SLxEjqN+IRUVPmKWGIwYVlNiM0/5oYpOWDvLYK
VY4a4qooQOuHmnWP5n8M4ez6Oi6s3RL3x/5KtV3YE+w3rrk9HilPJHUHOLzuzR4Q
VfzVMatSyOIqWQ2/RA3AQiuxr6lrNKbQnj/KLbAtcXiMKF8YDzcnQzhqtNUQC3VE
xcJ9UHQBu327CbIj1PQXu3aZWitFABZ8UHOwqBqGCNrVKBpwOV8vMb62II5eihel
wTLek6wWQTfmAN53ZxZcAxJexOJevibrPpKKwhtgZ2i5IDF9i4IB9eG3QTJoMO3F
6Bz6oUTQbkUTVvzF03YsUimqCGujLSPy1+kh2ThaiLlvDcIvc1azcCqG3MQBKKId
bDurgFOx7Bl4uPiniX9u9QZ0xg08ORUEfyIOyuTw0L6mLtXJGx55dbP5N1uGoMyW
ZYUQIYPL3K3P2jew3N9Eid1OdmkEwCf/esHmMx2n/gHFChIafiVucq5XK64tEsbA
OOHd+ghcdYrZitirYRhvpXJBl79V/b8ebOCed0zdsRyzKNiT08slwZPG9p/81OlQ
lZ9MKXcLYrTlconAq4u5ROS1kRh4pyQ9sRIDrR3q4or0j2tToKfbIcwlKkRZjq9t
HmE9F8omHYEzheqaStYq4tLqlQLvCWdl1RJqHhg58+S0zTphJNRKdgE62HWrfSqd
VfAZX9UokDjgSzhJQh52k06LVoHdCEI+b2N6O9BYGdwOgGhPW/YXPJf2gqois+Gy
lws9vmqu5BOucXVDHtPp9NfxY9fXDz6udbcvvRhIJKFPRg07Un1KoK2vSzTEt+7K
jn+9ESSW39N/G3WZeF31ZQNZ4xqPEF0cF+BTxqdneWfDnFflpX2CoK0SFD1DNx5f
YbPvP1PQwz6gCFJq7pgLA7CRYIa4afAVUy9Xnf9TjKQzJMCoc1+cBGmPqM3R20mG
eLU21lqgBfkmuKPivVom2e+7gIQHeoNMTE55/LMtFQy/mPbXImZgpwYFKooDJucS
IB2knLIGW53k6eWdOWHhEiagmzlG/HDHFnP8vc2Ll8w+nk2zqgH5DXbFq1BIf39l
P/6KEKWv2cPvFtovkJLvUx/htQJjnLX3a2l14TxrMYo7q3qQFH+vbeRnxmVzUdwt
Dvhs+nKLtpjvdw2xP9TFwCJgUrx3JM1I0+tXWXvkQt+nhR+Vf5bvckOJb3eCQsLa
n7lICMu+NAzb84B2+rRUgEz0GbqurHstZE16Tww64YWQM6iSL1polynJfI43IV1H
BCFWedX9ThMdOsTMpo1r9JaLUl6AaLLqmuSXyCjxvphmm8TWDcHxmH2yLHwlwFjH
JNyJu05D7wMkvgFhcoSehCRvHMtwxF5srLqtZhQmKOVE5iHVjXDRmn9RzdDGvUfZ
bzmDZrOk/xvTYSVBdA9DC/pGR7DHWiLKZ5CasMzb1+kc53Ayv0F8cRBUwXnnObx4
rH1M1cRnmkYOsA1hojByZ3pLDHUWBLiD/7MCvbmF7ZU0spTSfXQ1lQQWAyo8YP50
CMqgtessXk0dNDTrGJymd26Dr56J7N5hpe1OscYbtDZ8AA2RMb5wPHkwiflt54o1
tsq+86I+0wUS3HKteP1nPjkjZdU3mDebPMwH4kWzbBOCEefO4X9sYFwPaUcsnlOb
+gZERDStVSTulmeD006LF7BqkPZ1eZpAEE/3IWe44Qb5bCOtPpoJB/ngRbrXUEKd
R9HYcghaLtoeIjTheuxEQ2SwBqo/z/POYXHG1t1huUZacLycgsmbWMpvdt6HkCqB
8Cq2grjw+KA9qnUrJO8OOFA/VNjgWYMy/ghRGPHtf9HSyrwweTj/76l/8AX4Hnfr
eL44LAOccdeaqjelDZkLaQMxWyaT455c4WyIcQ2xo46HXBSyvU78pVA1tp25MRjT
oaoi7DeQ/l+Dcd5GfwWG7HAY3+6yfGEu7zSm2z4dWHClID+dGcZI+g0Mvx07yG+p
3BSC1yvNWMtigkyxrLapd+ZyuSweiroQRQmhsPEQzJPYBBWiA3KBbpJ1UMALUNXo
pDzCmODhC6HdSUkMt4MX+A7CnPV2Yhwrj7bPYf8vVtiC9TzL8pssx0CS4RLoV6bf
qms8qqlVE/9Bxy49alzqYhDjjsBd856tMLxHYg/tFXr1w00I0nIWNs7o4Qr/dNJJ
1tbjlUo10nkhVVntf2uRcnalGtfPb3F+ZzV50Cw4vi2mDq2yAvGa50cDKuFDMLeY
mSiyldeSWpc3ri+lwc1PIHFW5AT2a1ok4GlYuZmlrJ022APiUyVmKPeEAIIWDA0W
it3LtiM2KtqNaVzVYjo13TPgn0i5xOjK7N8Twc0Q6MfP2GAMlX7yNjjBoLDyC1P+
5zb67cKiRK0nDe9w5PL00z4amzYIr0ZnW8l8D2i7bJXCulquviOxeRTTdLnblGVQ
kFaBeqD9URKzslv5ss/f/dn+ghri0WHYi2k5VhklO+MT6EGAnPYbaxM+pfKQnXir
qv2xC/POpmo4F79fBUcATytlo7NtXTPVVfOpULAAr5jUa+ztEM1oHoAhQTDbsmQE
ohFR3BJLmEOdYLmB3603sEwhw9jTivSRBFlSFoJ/ol7y0OKuIdhnPGT+W5PJdXY3
OB8HBuNfdXiGPPv4ueakbNsJu9lO/qP1n64zneEcRfGf39aZAydDunv0hTX2X4uW
Fe7Z5vJVbJAex+cTqGQCdfKueXEfgYb/WUOZfN3MX0bhXSyCvdlSuBuvjTdw3ATz
9MGoCR0T6azfdYitwro0QglqTgVfZaTnz7vSlKMJNeqENw0MZtCXCXU/YOy9Z8C6
xDAR2Uj2ZyBIDE37u2ngzJ4cZ39Z3LUxCA7JfXgkDoi5EAflfNdkubhATWraLqa2
yRuWJfcPWHoTCTMfW4VH/tPhSBrs4T4zwKUQox3HjK2CtkERJQnsbH0FbJkRhoal
9eYrUt1QCEb6Wdmwkc8Wu8zB9LFCtY5VJ3wSjwxRAi7/c9iS/fdkNjs09ukZ6TNr
JM/clS7vJl1PiBT7ogtG8M/GdiN1qv6JKo082dAEPQ0BG1G682SL/g+ffasyWp1J
Q2eI4MrcNGnrYQFPyoBC/VATCTUKukMoY+h0llw/HuNXv495HR1JhssbQB7QAyX3
MMN1KRXhuHDrn/D2dGKh11BKLL+ng0v6vtKYB3MCqbJpvdUA9iBU82jg8Thhl120
WVMrmXG/KMRpEwXHK6/xxlZtj2j7pG2Vvr3OHrZ/+TNJj1ypH+d+Xt3jtlhez315
t6q+dhpXWGoqu6oDigCAXXz6k4aqGW0BxnUq+8KMYll68Ie0VVwGPm3MXw/833zR
i1xOHpxlYJbdrwACDHlt6Ux/a3PUj41dMfGsWBql8M1XLL0c1aU44f8zTyoyNv0O
0B/BFeUtrcB1hOGStiCsCv+Qk8r8zAFeBcy+/cPZLrCngQRV6/0Q6Xdwny/Vd4VF
9IQDHStCg1ihxAqcxs+rsONcltmwbUAUL3s0d3Ua0TDktW8lfyOnaruz572RkKcL
iLO9neSjnCIQE2oK2DRCi/Uw9LdcH1OCkQ50ZnmCxGbGkAY+n4mbpotw8Lbb12IM
GGGTbQudnwpdjamp3p/PbS86eYMNRs1W08yjTtmwTvH6i1cVBBEiVFkz1PWKtsGs
v2FAH9MLVuTy5+JyxveqtnDD7bjbTOMJelcQNpSVpuELII9ZeevFqLLBF1IP4qC+
XvcSc0L+r+GylYjaCD/pu+N5q1DjqzwVFgeS9/YuEqd50p7sksY6yRtyaJCYGV5G
L5QV5eGj/2JGemfvyMmaDLc7aLXVLSWrsQnbykvnaDcai/fGDQ7Y3KV7EP65E7f0
r4XImcF/PCzOddEV9BFO5Bf2RmZEkIJQRCCVph+hqDfR2FOPCO7pXlKqlWBeUGq0
72+8sCFlem+TOM5JlLRvX0K827CD6N5aLm46+SIQOeI8UoV3jjDbyhN70++iANgl
QAhMcbSTJioN8zBBgG+8KNcPGExXjnt4bWg3XDVGjH2ZDxHv+JStZIjG7ycAJRvv
T7f2jGUs9FNZy6iPmNJKJkzXgofBie81QSnxJwkLqzokHevnY7tuZkTqDlz0TZkO
KYi+Rac4kfKxeiHCfXQWjPRc6J3mAIDGF9W1KslsUfadFG7VLnYINF6PKBk6haZv
FPcUXA6ueZeXXsowY4N814/adfrdxVn2ySZYH3KYMKfUY/lwI7soS4D9gxHziOyl
+1GOw54oJuGQ8IIunoq2FwH+jBEqh6EcqRnxuNgus8a3qBUEJuX85YoQXNAL3SFH
9kN1JUClq2veJHio2Hj2/wK+hzWKL3zb773dIjNXgd4HJO7BDgRVroJakIhR2C9V
5piRZmvA4V572hv8qucX0tMTj4typNaa6tVtPbLbUZb1yEvXIrCj4H7HsvsOmwaY
qlkA8DL+eF7c9gRYDtpVAdlyRf5Zgm3iLZXfCznh5Fduy4MIaNA7LoCFlh3NtMtL
P4SAz8Gu7EspKS//RhIImOv2m4clYQAO5rRaIGfXjTEJ+umnO0v+LjcVUAEsYiPn
a2OE/o8I2hcwpIgM/7zOYt/5ZLCGptBy7oYfgbFAVoqbAexz3qKhUbBYgUdtm1g5
QTjzNWfhWIAg4wgr83JK8xlAkFj0FKb6YCeLbPTMei6XZ81lKaQpM1b6vMfNjnVx
f2Xz0QxfPTVXbv1gSxknB+KBy/7tAhH+/XPVIpt3OqZR3tO0oQFusQYqmE9ueETL
/BaxPwCUliVcN1/cKFu4ZN997q1BBEZ53Dfd3R6EiDBUIhkIRP42TyrL8y5thcSo
26WtWvUEUTcPglS154/mxmLrcbr+29NOjlDurWIgRtjghRsYV2DFrtIqHQZ0MqTj
Hbni04YNnC1QOpwKHpxbgeBWMCu8VKXGmei4b/tKHhgU1EWW37+6SqHCiQq4Dji+
i35N6rdLuBuJu6t0w/M5fvEACE2vO/fgGvpudy+8NmEPq//MPM0KBsVXbr738fRn
vnNeGusQfh8KgQ1gG7VC8JNWQSXsBW5Ry3llg08UOWFI+gZxxu1jw8LjNmdfYpAf
fyVawqWO16kc00W/Z+VJsum6eTBHssgHNVC6BOq4M1dKjRUafX9C0sm04d/l235e
578ZddK0L+wCeRqBOhoXrYa8p0d71MJKWTbpvLGP/uV/wO/erA9nq0V5kHU30tJj
TYEiH48QFHDHTvhuCV8zkH2rm9i4Y7JuwQyeZrG3Ei0v4vLh9imi2KPntoJ9mlT6
CFxNJUnlDxbnvUjHRjXtGUoanGH05KQRiupc6xISd9IwaqOWKePNtJOGPyA1wOBA
v6qGer1tRxYUqfx83cgIW35AJdXOGXmlAKqe6PDEUAq/EpOwX5Ojw5gy5ATSI9jO
8uVtbV/FBUxB+gyvsEtPkLLZwspDcw0glQ7V5WyRsSEFCe9ImC0jLu6YmN3T+F29
gN92ejGz0J2y33cS9FCNHXdYS60+dORlHB5dMpS7noI8iTk+eKuxKMBbsPiEEw5e
Gd/+hR+Nv6vbgIDCPhCRGNenXRgj1REuMrJtc8S8MDJx6KJ0XceY9fThPqLAazf2
HGzERZOVDdNvf1yv5a1D020gLJ2BC4nIZvs40xPuKprhLAdXS/o6+TBtl1ATn/UO
s1/uuwO+3wE1E0FhWJI0SkPKP6Wk+o5TzKs1oACvIxx8K/v8EW+9wiBpn+koy4Nq
newCPJc9YmxTMQEqlVHLpUg+GL4Um3SV0PFdG/5vXC8ye+kArxWAfQJuY3Ie72D3
zGRHpDCv+AVv/FujMCIgY0JQI4R54oI3nmO7nlf1afzClhC6qVWcJnDhStwrWYy1
d0DiLIwffYEqyqOQXu9NNEWfg0NOAiwycP8e9uNTWzgLHj6U2NR8grGKU3Q32NuL
w488sjvkar+GHWG4cd0XnspIvRk2YqdCVpyOKAgrPsdhcNrQndYme+ZkTAfaoZwb
idOGTres99RHJe2NBTKtDWHcEuoGRnxtwwLF1WSi3x6y6k/sCIwvOQufxDmjjtrh
rIkxqblVmi1m5rAuYwQSaQ7kf0SP2j4tUyeX7imsiXaFoQ0PXDyBK1aTiiXvp/Ip
y4KxOrOcGe3tts8oMRTRuLYxKSISpEoixQmI0CJL8Qvn4JrrYp3WfljL7xg8BX+L
GfRcVfiduX0DXg7owabv9dt+ujLSUzfpd16eXQ8vk5i7FMmRNT8UIaCvAQdEZe0k
9a8E0ZkxYoNAioaRoVr/oochTo9ygPk5n4BOLwGu/yliGVmR5+UZc22NlAdGyfxM
hsC2BhWNoG8rxY/Mm4Hl8eSI02rvm7L9EN+GcwDEqwOfCzAm0ER5nio2NCgpzuPM
vDFrKodm4QhDTj6SjNDTifVQYB23sctJt7xgxFhkhXuoQ6lcv1iquYQAzSYKZxcH
lXM5rVTghslewabeZ+MDKnP+Gl/qBODx/Ww1QL7GcH9U9zIr6vUM0EoFuJXh3IJf
M2mIfh0fJkntuEU5XL4CH7GyZAcDmsgMhhVY9dwiDcXyYJckAHARPR4jdGumdV4U
sX6lEQn5TZDYu7t6JhtQJkUXvhBkJS5HWruA01SdZLBkN8flP7nVgHcp7LHGEN1N
SQgUCEb/cPgy3HDP4BrHGmQeJWfTnmy31A3wDDp/D3VFWj3Qw4buHx9UfoQ170N6
TG/HjPQCFJWplhsCxAPpiLVGxhPVrtiMI/5hWnp0Kw5Dnze7Z7fz4ju3OlQ7+fPr
M7TMtg0AvcYzdKnmeOU5+fX3+m8dBVWFgSM35rLEnxUESqXAKXruI10AN2n5hcm+
NOMzz6frx6QwTZgeYwI66t/iOHUs87MBdCrC3wWz9ssZaLSOiEpwIVwfuX4FD3YM
cs2e86DmwuEbTrkJ5/+QNUoser31qBBbEn05CivbA2wWHk+JANbeewMIK32wIDJ7
gR7qoa1nDia7Tjv/xOyEZk/SyG2bBB7u/f2DcUgXms+So1wZKS2go4eEkOu2wRtD
XGiOYhjtVFwOV7suRd7SJwgMOOIREuHAbiwPBk6wyehMoTot+pFAZvA+dpJuH8e6
hv/UtLTMSpZFD4mA3Zz1tL1/58QU4inVMAHbfzY9GEJw+PrIV9VO5qXi4GT1NCB9
dWEB461hH3RwZtr0u+KZ1blLdvJiNpBKzRumuwSG043TVS1IO7uiFeI6fAPbzVRd
1U+W5E2LAY20kPWNDRB9NvXIoIYtqtQYJ30Ohf5gaza3XyqblYTm0ShoBDXNB9AY
sqQTNNfDUmulNkx+60oA+LhF8RG/+Yu6eqFZ6SdfomcySxNDJHcrrk4Yh3DS6UuI
CTRXqKK71ykCpK8FiF124LbhqJepP3fLsov/WS0OcVGyBvonJx7PKrXNmPWoPC0m
yxArWUSBsEZurP0rp64TLSYumoaEmHIlCGx5uN/MtpYwcQftbEzF3Y79/3vs2t8T
J/P+rfMGivSjeTQJfldM8SxvhRe0ogszuCSvlCTXPrT1YdtnERLRf7cF7a3tfC1k
A6dnjjZnhNv7mGGeWbeHyMVFmIMNFdHaC2ou84oUaQ/vieYJbof6g5ilgt57Da3e
+mersUqJxAhQdoeV0U7Q3wiuIS+BiFOMAzH0M1x3OD87gIvQ2XMjJX7o+n/7IoHv
Gx4q7DOlzRNcguF0SGfffzoR7f93YywEAnZkOZEHuFpFPpkOPAR6xUKuKloXXDHS
rb3bzFP9IF/P+zJIyLPUZ+Yvk0SFSFIz212Cv0sFTVixDerbbGbO+D58hU1byims
Fc8/IfGFyV1frVIIYdNSQsyDQ/S7TTkfe5sFIxJgWOVZJYTqJGcTNIPuq6iigM3o
J3Feq7Wl2aoiK96JDRN7gHyQ/KT5AuSylBbfo3pJnHmrLzkVnSyF9WGny5jDPJ6N
Phu2774PS0p8Z1qmUrKUIhMwDP1p28LAM+/Y225WLlzQtmZiduBgTbxlWG7rN6GS
SJXjq0i68E6cUpmsBujtXZgWmR3mPLRNcDRJU4JgRDrnVQ5BGmOOz/xd1HfHH2O9
WP0Db3W7ddzc04IaJpwMhutpxDsl284v+TvSMxjoJhOis35XCvFgcu6OIejUhXMd
BfePcI2sJLS8gSb09M/Kl+wO/8APReUfdcYrZOdN4IWhEQu3tu2l3b/3B91hV1R0
ndC9OX5Sx5sR0PvUKuV3Htm4vhXFUVCv/hMhj2PIsHZ2pvm0yB0yhnHgR21mQdAd
ukEr+ySPHNinCxV6VfU19+HMYCVx+CA/0sKyqk4MN26fJ+Th67C2Eo04WdL1m14z
EbGQJx5KTEMmsFSP3iCOcOzOTHEHjvnbTMXo3mc46Zq5id/NDO64FYbLQFA3/Le3
TB+Oezs9YnW69bf4+0iChJIaqw5lQwC2X9SS2RN8jgHTY3V10qimglJnjPjSv6Aw
fLHsTAc08Cy/uJYq2P0l2vbJ/eTrRXjomYuzgb4OTDvShjDYPX2SJJxShHEg6QiS
ng9B5dr0k69h/+JveE4AzmtyOFLFd1H6tu5dyoo2BXAPUbJvvdYIrLy8DMCPQdc7
ZeS7IFG7G2MbaWpfynjDmGgnVB0aAcF456HVM9hcn61EsBhqhb+X3O51SdAtSU5L
0IpQSTDDAKS53t2fnTLix0eUBrMJo7ZsKuX0fFVwbWNeebeECa7T6cOfio7+e3vb
3xTTd0uDNY0eX/VgABjHItDX3vJy+ur71BQt/fIVrO38udBAHEUKXsr79xF9eZgO
ECtYThILTrP7LDi8GwfSZnbWWy35mEtgfq76W/wheeOPbcBEFlmLklsmhyJzgz17
H6is2VOSB/VCDFPJrtmLiU1zCtABKeFRpHjkYqAvd13brCYE3OWyf2M4uWlgsYKi
/uQCPXUIQlgcwT0Z2krur4qfx9g8XhdZpE4QzRdvZ9WDD3UZP313Q/0U5qp77MQd
x5ZBcHzE8+b+YG4VE5zw2qPa4rQEWuoiOSCkZTbDG45Xulje2f+YLICsdqo/7xni
km704lBcuTGkshUn0Y3j1BjXuydmUngH23oq+64hSjEOy/98MX05W0YlJkfiH7Og
zXysvlgnbC8PyLtaxaeFREiM2fTrBaspkLhyUAfc911NHiSzbfroR7Wj2oSWuNq5
b6yqE4DQCF9ySMhWvYYSsvmTDt8xWXAJs0iI81KmfpvXTm8ziSbyt20HUaCCTpJO
8Xu/SspVLLKKGZfo/iKLPnersuABSXijccM4y0zIshMmff+c1i2tXu+9u4xb3n+z
4EH1f2JJvfrPdXFFW/TYIVyJ3liyDsYEZ8yEHKtfFKZBQDHl4WgU8Dpn+kVD2rvf
ogEFV8T8PC26uBVvmQFwPXG1xfg1pLe90p6JZP8m0c04pvYSomcwEEde4Rza0CG/
k2/uBuiUWYa10HjtXdwyZxkLlDaCbPFml0bzv2z/z2RSYCs8dY4+j4VMjZrg+R+N
m9Ts6NdCqcjU+2L5ST/QjhpUOIIUATygsNrMj+qBgZFBwB6IxJGqKDBFNri8Zb80
eg+L3LpuliJDuK3R+2EuiIdjxNTfyTjA/H2xyN6ih0BoryP3ViVwal8FMCP0/Vz0
AYBAcPyPvYO9j1BbFWCYfbw5eBq0ycqfRBUxvpAD74mT4gEoyVRjBHM0qAnmHLoJ
opFhkH+kprovLmgT7q8z6FgnT0ADwprjq80mH3nuMZn4yv23pY24MQ7VAFq/Q+tU
Z1rgJeIp35NosotNUkM+2LG64USrIi0/EytWYLYdmtWdWfrMBPHOS/RFwHFmyBT+
kp3UsPeg3P5v4hjWo9iwZM7fbGI/MB/0rYlKCT3cMj1LvaKF4FcKahDk7C945zDH
P4hdd/AGg7zuVZ0xeJXGQ3fc9IDxuU1734FAGSz1o6j0fLO3BXiVa/jVLJQPPPHU
sR7kG9cqDYFVhC1D4x0YB9P++UMN30OS8qwnqeij2Wtxbg0hmI1sCG05y9ae0Nng
7uqMfWkhGBWKEBgSExQFGNedVRZ+XLmwTpKZG/AXsw6C91mQSK38ketyx9buQ1dR
TUqsu5y9RQ8z/8UcRc3gMIa+btVOTD0FUY0sxzw96QY83EfX6dMXn+d53ySPN5Mw
N4RQZRPRYK+na9STPl5J8uEn756L2ZsLJ5V2bNq8l8E8UNBknesBiHrH6DKp/zLq
O4qPvYAdT4C672M/zfbmY6vZOsn4J+3v8QZ0QO//pgC5gEV2DUBKTYhRzyAcD9WW
IovTb6RF3Mf2AGljL4wo5nmZTOjpulpFST2faehdZ+DW85unxhIsAJuy6J724ykQ
0YrWaghdahG3ITKmvjWib2dx0DcAdxOT3SRCG9xMc9MVuwPvZmxINlyxEKER6CTV
+zeEDZCqRdMQpRCTmeRAXHyqMZPTWHirIm0zRaOtGjrTe398kVDuOYwikl/ekjTz
D9FxHOHBByfKrBu8VYYTml2/1pybsssY/oLi413aeJrmBnJTsF8HwyZAEFmuNHNN
yrjktbnODlEqq3UEYD8ZHiFBO7qx8hijgIr+FbwyRawm0EqoV57ghiLcNWG85ZaP
fZGY5QxABJVrb7X0FK1zexAfYEKQ42Qa7TKMNu7oHecr5BuFQFdmaTplFcIgdQZj
Wd669xl+FnKQKwWqDAsKOlp2rcGteRJFEGpQgYcqJDkxgxp5h5id9GA/97pqhWC2
nwH/aQoLDY2uOj5BqNdur8IPNgNIBu9oTiJZF0DKyqApXq83yBj50W5BWIh6kbx1
tmMDhMaIk0ICuf8uXgwJWUffqVAvMmFaqClMBlR7L8ZwrH2SmLKxDzKQU7v7fxRz
pBe/v5/1YyET05efy7UFue0o23IoWcO5v0Zoy9RE0qzmJMxS2aNFC+RdqwRTHWOg
PHDZN+cHIN9YkSdPBnUaoffKcnFJ5OWXchV0yhQmGtN2UC86Z/Vf/RH0wUrwd/Ea
bcX1rDxanh2vEcUEMBoY3elycnbKKALZrkwsCHwyI3AP7aY6CnIx0ZbjaLE5EZnn
f9Kzt/3C8fcpSk5E5hneLZm8CREZXLEevccLmKjI5lF199+a/cbfc2mIWFIIOKBQ
V9sFd1rUaO5TIoXVR/G1moGyD1B+Kym2g0+vpaInBYojvCAI0yNyNMUfDSv0BJyK
13+9oSEOYKD2wGcPzsjM/uFLnFtZ4c/+DQmO7+9c4B3ZBpX9jSE4/P9H8cE14oMb
OuuFsyXITjxD7BNzP7aEej/gEiU0UL3G2BjaJUmgtP4z7p2ENCgFWznJwLBDFy4n
sAQhzpQI2lDN8K4YFQCPgoyjeWCZS4oGwC/O4kOIjd4jxwIIcLnxnr+FUg0Q24mB
YLDjfopB79ZyX8kgCLf18A+PmLZQs1JUKKEGbJqrL6b76MUqQuwzx5Z+ypSoQhHZ
USBu45X/GKgRNLfOPTUq+crcLCsqvaF3PU12cKOfKccIpxVIsyRz8hTLBoLrDGM9
PynnAYwJLkhIa7uPN+70ZRjvr15/FYddrjWY55V04+hqLXwFd4Sn/69Pq40LnJMh
rLqZwdfI4eQY540xY9nqvQUfEz1HaFmeuaHnk/6fBkgY79FWBVdjpmmzrDXmkGwE
FPx/JjoeiBzeHepTmBqsfV88UziDBDJj3mdvBmRhDSkpttVGJJVJYZsWz+maCQjR
j2ezzGzRcXkgL2NS0R8Vs73Qkq/hmgN++xO4eSHWZwU+LHQn04wv5waYiphbWJMX
zUQHcJXNqvIurizdiHozbvdD4tCFJ3a7edfEDstlx+8waV5quFQtvMx8MO6wsr+s
+GUGQVhMf9aBoTfIHGoDsxMHLmYVOM+PaIZudp9D8LvqGfLa7EXnd5v29Lo87dn2
93MhaxUUmIoh3xuGkZMAIeClW6iCFhsv9baFT1jdVki4O5JEIpEQViJcdr/MImOv
Ygvnv7Z5bUd3o8mWt1q0QAwW2RDjNdjP4aah/yTX0FXdBkyT7gO/uDwsCvAMCp5r
c3/MZElzsiQCvyaHJrJcp1RrTVVDPCSxH04tul5P0CTYu3xbp/ZL9DlCJl1XjOGk
TsFjeqZzrgqFsLAfvGcr6CEfVtSlpc0K6cED/KT1zFc8GGwUUBN2SlkkRbzeg8hH
MvSaC1xcOf2CJfBeJEnKjq0UU+qNlbozOmVj61pVuV1qqQBbxHYRXAd32PZjOEPf
nok4ZySYxMKSuO58pnkHi+N7JMUIRIbnyXE3cnBd8+47XmceF65uowMvb/e6EWIM
qkFdtOZtnfwFG0BTa9uTQjhLsaDOosiOgb2KMPKzo11ae6QUsQm7ZJNtMfNy2123
WEKIAGKSP5P2ugb+iuVtIq9h5dQ+BhjbeMQm50+LtBxkgy3oU49jlmus8tvX4j4R
25TwLydDKjgCVRTQbJ4V7NgThysg1sp1syVJ+jQ/c11wIfyesAM9chJSktla8dlA
UqnbvmDGb7l9uQoDsMXwO4hHcmUFPuYlRHRkj85Rq4mb7gYYfnSYm3Z+5nfhXlBJ
sanp/gMv21q1r8GX7E7TAgEgtuKMd9NFu6zKI/mCng5t4q/sPIi+8jrnQlWKtlmy
2x/8IiEzQAmiGfK6FnZVluozcMq4JnB/ey+UGTfBzeEpeFwt2obtJkYNX+OMbclV
BytiQzmZHAUnTWr8DczBDIkEEmFXBycw+I20W7EPERlqSbeSGmsQsON+XGZ96U63
lLQJplxsDhSsKW1EPoUi/kht7Z+HCEJZ9p+gXavQ6hZBnEON3+xJhVIScHZuCKqe
phAClRqeKWyAp6h9ZnqTq4a7ivDZPrlAOnvjWVpjUi7ffTHXXe9+MjTGJszZZ5R9
XBaM9useRqnFgIkLkvjs9yk6go1YLd7UmQP6xfamBdx7RnH1kvx76atkxK3KI0dN
mo7pM2y6nolKOEeCxj3HvQffAPMCai2fKx48tsIZiG09RuBzaHrcHegHLkFcxfCG
CfHSAaDDzxh5hRkoU0+mKKBKYoYjV0QivvPRYlftQJ3pUlWJ0g4qd2098INaTemD
flf7z9RoGAcZAT60PbmJQIoJoDztaywQpvwMgVdMIjxdD28LUcXmAZf0BDKzgPsF
s1o/zN7B6OwfqIJXtC4+krmcYKtIR/0XiXCKLSWsKmfEHWuJCsa1pnx29moCgFKn
VOHjWpm2EtDB32HRVpS4nN9KJ/JmYkeimgjY0QBhNIWnKbqTfdrIS8jxSgcPxv+U
OVcruJc4V0SWOni6YQU0zbWS/cNxHWR6NCP8S2qAggLvVwQnw2/Loga8JAIN8FxN
VbhlmjBOjZ89XZ4d+INh9MdUjyj/znJDcITuZ9vh23BWJ2BL22seSm/fGbhjuxru
IHN3Bcs6pguWorWu1x0hO3bEVbSSjusvzdRfryowki1VFLf92/RZbws02xZ/P48c
6uLuBkjjUH946M3Bibvn5bwIDUtW2qYHFe4iAIySrqCsaigGGo/dMV2/dwSPTZ05
jiHh5moB9tZ0JHY0CCCoJJVNEnYy20DlN1Iul7HfRdbdSTARn5DaD/n/0Ar2KGXq
7SYoayvRtDv5Dc7wrMT8rx71qXAchFRqHKjzI59lFStYEVJg9idwlpK9xM5e7yda
vhiqx6kX4p0JLYMz9dipz3HP6rQ8MggPxOIo7VCgZReYFCdhe5eFAsaoLPjHhx+B
Rn5Q/5GyG2uzbnAQYU8fTHQn9kkfTRwggNOf6qQZ4qKpBsdzcUafzycPxgj9KZ0C
6IBoi27A6aZ3FgKIydJes779VX7yJ7xk/2GM0bDK6eGw8oN5CsblFquIzs1uO2OS
YCEXVCtSNDPbfxyc6MlZUatgenVVGWdNs6hqzFifeLm0dopJlBOCedqaH966Mfcn
huejKkM8Xb6S/tf03eLMOcu4Y6+CfZIkxs3loH7oXsgvBA60EKFoIqYApWc9VqDG
Dyk60Lb/Bni0k9eOLU2a2Y6ipK31wASq/d51xk9j5wOUdrxZzGjxZr7MOveHz1mF
3H7a26N6LDtWmgxEByad5YVGxnNGUEty1W8jGtvYvRUF7+o0soBSeEFh4EZnUR9H
ZQHLz/X/uAAT8HIqJWebl6WATssVhkpgqqPiOyThxnNpQWGL7eQ4qqs97c/g8y1l
w0uUzd1IJZp0eIyvJtGc2z3mEdh/fTK5bUP7wHxgONoCJ2dcwZGsjIIkalntNpNY
DouXl41HU4j3AivPUHhHzWGH7lruKJOLtdnARFzhpy5snrDCvvxm2ihq4XkeXIFY
ArN+0iLUklM311b1VxSHD+VDJYwvHbKxF8YBNrXnFfvJneGPHywZXgHuyg+Soma9
vDU3KJKWEfgiXsgNB5daeNFwY1PIKhnA0/NenQcNvzyrUhYzIB3vk7gaeR7rWxGE
3TOVOQtX37dx/1z5mGr0bkWUBpvBfE2xc6q521aEw6W1taq0EQ7Zi8CD7j7ZBZbW
b+Urx7L/xpo30W85vb75saZPs3MNufi5xwIs8vILyeXYTe6OgyZ6oLfEGghxeey9
H2OHrnwMcuVvwc2BWP5mzBDvWJLi1AMyFmqH1OL9endW0GTTwbhvICSikAhRc99l
ybPzv2SJs8FZzkX1jXE9pdC4uDlpkbvqhGYkyqa/zoJdh/CPfXO4K/W01BvIG/bS
BDXMceaFPkTyCR8MNeSI5LkEpw9gU5MR7Ny9tZw8irlWLzIsnAIzwCW3fqwAGeKN
LLrfuVXws8mcqc3L5rKA0WKcruLO+6CT0zQpqkSjxHxSzR05n0R9k05b12H6sq66
3jQo6nexvvzIqBZAWxiZuPtVBlG7cXjfWDIB3pjMFCt1dKxheXR6ipEFBCVWExaE
rjIW7QoXKKpZCtkSDoIfLBKN3BxeKuigoekTWJqGjLrzVC11K9MYdOM5C/+0pDcE
KNs1TOUnHSsMVCrmKQVZwueWg+YGyuhQfxTKRTsvFKGJAF/v488k+i27gGy6I2Pm
UIhCAWlkFKa5x1aZ5FGaYZz9zhFY8Bm8d1Rm2P7oCpvGDBGXs8ad9VT+30MclmA9
tT/646VtinNCopj0xK3fufpHlKUK0EzYa0S8J77VnEraZiGmOVKdqvUATVAn5FI3
uejZbRfr0UHcYGvxuXHoGgZ64yfX84h0/JMEyLSjEm0kd8LlhaGne9QFnf2TW0pK
tAqRfRh2Dyg4WmpB6HC29rIfTbvh3SGjoQwD5aLfh3zEVnQGoGHsIcn6bwuTKfOL
ZScOX8hDLAAmX7DbQQyD3T0nj/QDd81oAuNMoUM+iwTttKf6eaNiDPPywlGwsfvc
wP5t5t44Y7x/3zhi0mKt3rJPhBjnl7MAv/HXu/dpn5BNKLtZYfTa8gPnmYm5w5E7
dIYA/l1yGfl30Lw+KKqNNYzkNErAGxHEEztC6qUGeP/2psfWvfWLqto/4zvkHRUU
7Yfc5ylpTe/5QF0YO4wa5IVNLcXiYZjvkM7aRYjOcc3GRhdOF25O6OvW00qeD9QO
uHWNTnwkUbgXF/to/JpE+kg9anBFdiYNxy+QT9McEV3V5ZzUsotnuh/zKtrJUfnM
A/tGNpK77xokA7qqHEq+9CiCNk7519erIgQVJIdY9YQV1UGdztAww4ufM6BslUAN
BLSB1HejMSCFMYRKxnZv/QURm6tpPI1rbZR4VION6qYUBl7W9GxvficPVHWc9WKl
t6gfEBmxtApXc5AaXbRxVbkWRsCQ4wbrq+OmXNLUGht/gYfrQ6zZutmRE6FJkQvL
8hmqhIP8YSvxprRMsDvWToxhveqAeVgUFS5HKqsSegkc2WAcFb3/DkQcCk7e0xCa
9SEbxtK88Aj6pyzNEuw/bA0wqWbKlCA0HWCYRSRL8wlRxWEBJ2S6ZfzaVrQ0B7nx
uF/8hs5rnpG5wa74mjUNdzFEufX/zphMmVsLrNVRIFESsIzqrXxpUO01wtkJvARR
g+QmiKja69KjebPkR3c2liDOyaHU5+VCqlg6iE0noCxiO/JAd7STHrgiIP7VBhip
Lb91kVJHHAzqo7hZaxVEctJ2iKk3WawclT2Uy3veHGtQQeHu4L80c2DV1mRwQjIb
MQC7QyOSq9LEVjHbJBaIo8bOupQ1/SmmSpsOJRNSzD9q5hG9Br33D75MCr9mimBn
81QfTUlUVpik1CXq5iB1UmbrDB9WDUf5nku8LslpP2DzkWzsqDlGOIMXF5oNjqUA
TEnKJdOWddXI9yGBJkbIdfaEizBjH1KnkAJl8LYv9VfWNKcEA6j0gpno4PSKR/B5
xotIbZIG0LwpSzk3AWQKTKwWlu9vCC1xdQ88WzPtcEtEceOfjlpwUxS9vw3uwpi/
wm8PAqE8lPRqbsKR35NnNIwRqKXRoKGB+u8zvZQaVn4k2ffgLrE32BAdu6/xvb1I
kU89ZfzSjVA4RLe1+JemGZJVw/INckq8juB5t+bS43CrDDZM40eNpGEQwfkGc0nd
w5prVZuK/VjBbP015hMqATbvv/H5YyRvhgmXzvoRfrE71UT0Dg/8kIrZtYe+AYcS
go/1LSza2kepbBHEW0btMPmk5UW87PzXou/ejp/nHK7lykCePGV4475r0eagklRb
kly2gkT1spZ2KNtHwc8t4tjYH7OMLEDOzsJc0Hecg6R/SEJ+OCTTUtWKLK+X0WOa
pMKGSGt5Bbce4WkDmkZV3xp4irIopAJuDDjaqShixTXn+MIGH9S7ci7dfGzjRvtm
7j2pe/qi0277sPSyIOEZi/5d0M1t1QkMCgrMEqfHSKmD9bsGLS5mX3ySqNW1KYcN
0kx0rkzrmUnikxgaKSvOsfxu4ZgGWHp6B31gvVSFFP7RtAx2Z/fIfCNyF/Z0sqtk
EZDP3jEs3vch9RRglzYTrsfdfkx7LyV+aEoC91uMdRM9JKHKxJiF2oorSQz01uqJ
FZjkX9W4HxL/ODp3OoSYz3cbVv17yRowusXDBGWx8trPwjLQ1kxLqqvSxrKP1txE
53cS53FNYvLTj8MvCJTrCFHKExnAGz5Ii7LVn1ljLXdUbBHWjvaKOi0GjHwlOFjC
eqAsvWlQvcz9cwvmP1pIbLOykfHIKjb49HGTXctfFvTt7vZTsPIk296noh2v4THu
/uDJwrFV9ebzrqjKMRXpEzGCXe/RaWt0gSw5F13QozJfbEZ1EUpxXWbv+1/8YAzN
RmFyiDiSfWXfaeU8+Or8HYSrGmrrgB+lcEiX2JLV1fUx8Qb3UHp16sR3Rff/VxgT
0JcFEc2znXpV9bXHoEN5Igzv2kabh6AaAoYcVYX1LPGI7RTrDclNzazFQwEe14/M
6bNpifPobiR+I32xZwRgZGYPqrsfwL2Z6+DpoQEDXw+XQb1tSzTJTJCknO94eiDu
y8svksu3ixxlhyQzDTbVki0IU+36Djl1pdr/xRxGaDNrpvIcyazcKI/keeoE1FXz
XO/ZSM0aS6A7yhYaLBXo4PSbC9xwLUeADML44QichZ7DGLV1bIhrkAcAdZBTkhJo
Zl90x3ZOfIhzB9f++RmR5h81PnPoR4GKG3RWCbM4ihPOdTir9jfW6Rg8EicYaKFF
kE7WbaTZUQttzZF98rTaCwSmfObTWse/B74jhwHxi1CcFa14PH3IJoN0EbSoGEQg
h37jfT89FxysLQTccG0C7BK64jVwUdPlvlPp0wF43MXnNgDiRD4lk6/2FIyzfmwV
xVONu+EglVD7tQ1Vr6RjN7/7Ez0v8UXoBh9NOnFgdTOv4pEDAvhDtCORKU3MGzK4
MTe8aLjM1GGiFIHDRBroS0aCKxLCBUCzwILAo1ulLydGonX3jcg5AfbOPhNd/r2I
U+PM0zZBJ0cCYHD8g6Be7OdgCRU6uaDvCJYa4k9xlPzeOPmIkT4SynA7gsMlun/2
fkFX48b51tF+w/HACH85Xph+lQwbwGB6SVWWil0qk/GkJT8c2FiVEmtwlSZ0pNNs
BeKSxeP26BNa5PGosF2GbEUoWrNOlGDxjLkv3pRUqroNgOI1h887YFbv7vNxaFXw
QwcqcSACQ168MeV8Ya6ia9ZHLn2AV4vyOhqM8+++MUavWgwGv5cHk/zT+uKjG15F
O3UH1YdltHoIlK5I3Qi+uhHm7A1Y+roiijKR84VhAunXfrTkRyF6YFTQQ/7NZnVC
KL3ixikcSpb/CFEbuLwyIIS3DrIVTu6J7AEjx0G4qeY5XjKAmGGNktz5hShxbb/v
p60h9itQihGncysIr9SzNblVCaHfyZrgVpf9uQcJaVT+FhhM9NZytkt621Dm+H/2
3igZnkAt8YVgmMEVsSUcWrDlsRK4EbyFXN8gSeZd4Wot/j1v0pDbPGnP2NcFoiW0
KDH1Uc2uUEa1YULicCAZjceW0r9B9sowOwL6JW/hktiYWhoEGsGBfhaVHcdmvGfV
HnWJm28Gy3FACeLFB6Ffc9H3DHAzyuOqndiA23p3LM6tnIYUiLjvvyS7o1TevNV/
3oOlj9elHkWUDghrNUmPrtX64uuSpCEyCDShjKYtwsEh+jL6eqd6CbEGE6LSV+UX
dXUiiumO+BV/ETXmyazmyIRnBa3IXxE3JOfCa4RvtO+VxmHip+A1TADYp5DQiGcH
iXLRmcR9+MFs7Tl6vqWuaTgcZ+NO2QoNdQUZuylI84Hn2Q/f+W2Fyq6bN72m0adm
wzUicqC8ESTYUriRveR0P7/vKI95V4guB48s54W1A2Wao919geigOcfTi5zhFr2R
l9ObQZlngF0Hd/xMVtu882NZ8YYfCH/VpPiVQo75qVxrugZerGMKIH6Cagcseb5s
KDRlhj/zRjHM7gXZU7RiMK0FgDXxoyq8CzwfHKS7d8jUqEow+YXFg65aiPKMKaUl
YM7lcOPnbyXGke+ZyiY5l7pj4nqwyVfP2tnPlcUHa+qugicBUU6v1iaKHlR7mb10
gLG8ae5do+NWEIJfMbcaSt0W66ScSS6wzebv7msYnOaoXSTCstupmr9ufgClUQ8D
rnoDA/hI5l3Wj9Chjx4se4H9YjQknOP81yLgYm9VeJVTxYwOaHby6Mec32ehelG4
etDLHuOlHStB732gunrhDN1i91ZPIAKMcPtHGAisCj7qLRlLlJVdFHA5SyQHrlYg
Egsh5pPVYpsS94SlvlWNbdDXs7zcH2aZ6Q0SDrS9Cjl3E23Sbdn+y2s1Xgzrg04Z
bujPMQjBb6TT4y+kOylx5KhJ+Whf2lTTJLfON4+s1/aaQMbg7MPMKT0LHRJCDaoQ
JdRzXgP4VRno2PLparCxLkC9bRHlFrJ06gsBpd3US7ctsUaD7th/MtA6VNXBuIAd
xO5eiex1NmndlSMQs30V+1Zz3r7pFc6DTKQNvyvxXbi/E7Jo2r4Oq6A7PeZDzTx7
Uk9OWYPWkZr9uPc5rGedsBbfWz+iHS2qxDop9lF/lXd9wfp17Ed7YqOzBoYvkcxb
1pQbId5OByJRMhBEiw+ULDMXvtlpxSwq3FpDSQR3QQhuTKm9zCrULEs5ETC4mOT2
/nH41ohVXwUm0rgu/hf1qJxgP6DGt2LDqE3pJwXKCZsy10GCLCnqIxB08GwZ+oHS
3jL7zYI8kMjGDb1LIUXkAuEXOkRm+bHtaRdgWMG3lG0I6ipneIx0zUaIPlFtOK4x
3RmGDrCwdXzdzPnaqr6Ug5Bqt6x3f5qqdI+B3cGcunLxbOpS/HSwC6VcDmnqlDdG
dK3NBJjKUmE6uN4s911EoNmlgGxu1kiOjs6784zQGTinWkC3sV7sbGGDG2M8OWte
GHfWP4LULBEGuthdpsRjBKPogR+gqDkkQqnP5A08oBRSBYi8YkikRah8exU0/0fl
G6fMvf2XyrVkpOhiOHxSvxEc7mjd77fudIDM7AoqiUennAGiPAdoK9FwDwtzW2j4
TKX+ky2FCRCK857ILm3BKa82lUj1Q/9IahObNfH+QcJmptGdRYUwQ7UrPj1SXcLP
3jg1LqDcfdWGilc+P6iFAIlLi63VOEK7jzVPGMBSt7N1x4azRhLRF7dd0J9DoThp
VL+qUjifSIUUDxFXgNvboemIVWUsIFTsiobgJaOyZ5dk0MxVtqYEzyeavuMe9xua
bXMJ3DiyqGzE1/HJR8Zep57km8bdcxcDEh+fkHPqKNzmrpMkfkdl8dD7tvlWQZHL
udO9VruQG4OyTJN6OvWIBBS3QkVNNYWUQvyRZ/vyQG7hc9AbTNYEbGH5hQdWx5+r
WgPIsz0J5933//9I5/mbmqJxvOaRQyUbFbLTJvDMfS2XFtBTYHaUws5th9uxnpTI
xtqkCCP2h0GzIdtdsPXiUqxtyaf8o6a68xLOnucG6xbXJqceQ7CHuMm084eNpRPz
pOZy4q56cPApSeUIOHnAGgasUwvlS21HgLMQuHmQqAnr3ViLs/6OpTsCJcZ+Qphf
8cFxi+/90/EQ4q8m5ecFsJsTmZGobZVpnoOEkWWs1UuPi9uUgJnNw0FLAXLeiMO4
uFAV3irS/bIfc34rSTPXRAxw0jlNzgFY48ZiZ6f6Qtq0AKHfqJczd6cMsjim88J3
YuLidsPuEKnjPPCe+RIzZF0RbblbKx+HNlqcdnxys0EE0OIciEwzk/LT+BWPJwf0
AQAllNPAoi68/tMshtc5tqGvoK1pF2dAYer3YvzxpZVD4JUpSGn0iTRDwbp5XWoo
pWYJNNB5KRI/68EApR5773Nq9bng5MBZcHkNN8K4klOpAcego+gPDT10/09yCVWf
LrKFKSjO6gD2undybfQkXB00drojGPojAIxCpwJUVfHnsjE+4ye71BBuehpaYZ/D
hoQBByhiub05P0Sm33zcLXnc00XwpFOm6qjADhm+9sMIVW60krpHbXuXs6nrxCey
w9tuytY9KwHpj74pq1664epAnRrWbPT58NFNEdzFUWvU1oK2Tp0vuCx5y+IjFlfh
lbClVogMZe6vMljSvx1Bh0+4JJxNlSC8EifJSmYQbUnuXJVBFL41H56lZq+hBlxS
M188jwvkkHVOpk5vbQhvXLH3u2PEEt68ysAUr5a4Lu5P143OR59egjjhfSGCVOpV
lbrm0YfB4krzayQbJ16rB2844sWJtINTkGGrlsJda72cqEKbHFw1RFuoZ9KTIJT/
XTnB1YkHgTpAvv5CV/wS7HZ8X6ljdES0YHF5lRcQIv58RsbWrmUMtjvzlK8OWALX
sfQ4fsGNLBD4lgGuRaB/uCF9Pc9ix7x1mrVpKGg3aPCiCjWQEoZ56bL2yslpC4iB
sFYoOOyYoik+f//+MlF7KlNrmn61G2vYKPsm4adBCS4S0xetF4j9fZuOxgutzM6S
SiTgGuY8+FvvURJVR0Ir2Kirzqb35sjjZkc+jzgTdvYXT9US2SVv/oaF6xrgOz8x
V9h/yNvEsfXBLLHMe54UQ7sq8y269oKRfFd8SDpxOAZN1XsRR6/yjAL74Y3GqGF7
KSnAL1mgjyTPFsvRT8VjyX1brqzGTAtizDlWAP87Bfcn1ZW1TqoTEzfyLAp6H0dj
W7fUZTFw3WZMNZS7iNs4k0HQWnGtOySinmJQyG7BGb+XFZAmmctWmhzzX7iQZLLB
lEcnggyD6W1C3JYPfeqBxCCzWbjnT40e8+x/DSby1hWnCoIw4Z745+eeyVdCOrZO
9z+wHcv2Lr9RHVlOVhRk795+iS0hvCFzXqMTix0C3Gefx1BmXKnz3MbRRB1+obmV
yH5KeDGD7VhmlzXUednwILMEx3lM1VJu4v92GTkcI0Um1rF4p+KPpe3SclYBdNJm
HGAdJhxVZSjiR7xRYUDwr1fvr/vMxZMei8tAnZSkoiEiaKJq2oNEWxI1jXSNyH+w
ziZ95lUZOlBgxfScQCutxgwvG8xpjHEr5YXhDKgESd25y6pKBTrFoRSPrkbnxHLB
PruocfiYz0E0Q3TRLhzG1fMY89gCXmdCU1JmGYa3JTCQBr7n3DaoevZC59Hx/DsG
EUTm4qlYTYhroaXVovcQeOidP1+MBrT+MPvvcT+ak050Ftznz7vnV18H90YjRZpY
m6Rm9N6PUzZLa1iElWjQRuLbymNBBJE9gtXgvSxrOVeFGIZiE2zo9RPebGdSLUlb
gC+vvt7nnUfayeO6gmdIoGsCyN29pWxY0rxSppyzgzYnsPC7VPjulozOZtwDRRDv
EZ55vfInN6eOD+pJQHJb5j7he/gqmKQx1GfD7q1b8bK5WBLi1AtLqN2HSYTA4qCw
zBB2CXK+A9LSWUAiCMT1xmH+xdUezZj56Nkq6u1bo/OJPNHRkqwA4H5KSy3qUPAl
8npNjW8AB2i8eFA7F2an6rKKrBe02JL0lskM4GKrQ/l7Y+OY9356noiYlgSWbwD8
ngpvuYprq8v53xUpercll5QRimF2OoWnqbrwE3DYMHyt4Jr5ebHMZos7NURXWeoE
/dUwRF4Mf84l4ovXoCvt+JmGL0VijT7IDfjQ8320vgGusQ5BlGa3Sc2oW4YlUM8B
iFJS1NvvB74nN78oKewrvH40cIwV8HqEcwVGXpSc7jhIOZ6yki9KKY07EF/2ewxA
JMywFivplEGjhB4/Ux4/qDNl2wN/86qlLzFxzVIqPB+cHozJjIp9HJVJd/jLMCmc
kDDX5Sv9hqhfIPR6Oze9MfudQVFH09cDjPG+kmJ7Xoq7/AF2uSIO1y0HTJ6VqAWK
R8zTzWCq2GyZX0nZJQb/ctQxxtQtNjjOlKa/gGHp8Iv3i/Bt81Wrq1320o7mDkzW
VdYe4P1mufIggi5/TDf36eqXLcKJDrcTkVJRzckagBJBw4MJxJhe3a6erOzQ3nYp
U+ZmdvRfAsrC+H/KEuwpiQnmMw0k+htDzUTSKU7EzwrPCzHyB/sajpox7dTjfr+v
FhgvZTOsMhUf4Wh1GjwXJ93oCfO+u97P/RC8OG+Vz6ogn4kYF4NSGLrgUmtjKh2E
vcKGE6O/J8vQO5RlaxHvOwb988EYOhZoeWFmWKegMcipwdj3ctW2btEGu0iZN4MM
r/k1iFwW8ocVBPnTensqOtaTTqRXsiCx/86inu0qVbzfnq+xROqT5DfqJ5Id5hfv
I4MFobwSSp1TPgb54v3weWFmT4AOk8LQzNYW5OxP+yKaybefbaDDe90BRcc4HgeO
Xg89hOrAzqfRu8wYdoLLqBBdNGl9BpuXMLyLutrqQh5NqH+tH/wsUHqK0W4VGJ+k
/4IQXZHJJZuPqvKFsqAX5cjAA2lS4709oHC3a2LeeqA8vThsDRVSj2N0X7pSB6mn
fF1ECuN7lvCv4Qvs8CHsuMZnx7TOhcmzRg0bz0qxVvXE8O/cteeSSZnTaXEvnqLp
NUOnD+LLz1WZOjRp52nQr5pm4dvWogA9edSeHfwwjF/wZO9AQvF27O6C5Ps+tY3c
rBhwhNyJPyNz9ibU9gkyKCUaOsaIm/+WcJmER0PA8C23KSx/AeB2rN5H1Fa45LmI
msQ0PAC+bY0UvSaDc41yscyo6NFRGVT8raO4B7gDcABY+TF1WWds2m1MswT/0j+1
hau0kGW5s4qfOhiTDDKUeytfk8opPPxRbsG+SqvXLKppZIAZggueN+BSsuhUYb2d
U2ictz3PeIL/HjnTInWO99yvxQd61VJDCai+CrvtzP+64bzKdES3P5OyfCAfbP5c
pJRxDOC2ppGKxuTijO+oJO7YoQzXoqstLolkSvIBgPdaXKJcvGpVPmCBtYHtJjIz
lp4NB/PNYD9Bl7lcwcf3P8gPy/xc1rG12gJCGmffa0OUFjINrgiGiPrnkv5M0KN2
yrz87nqxaNZrcBfZI5q114Cqe7e1hpF5DYo2zCgMppVDg+lq+2UilXrkH7CSIv1h
fEa48+iMGVEp1jbgg8GoRwsv/a9vauOb5WX9rWptfJZfq/0TZ99v5hewjBnbqSNh
tUJL+jlgNBXZFUMlrO4ti/4hre2TF4usF3rQG8OUuzD0y6STWRG2+VD7y1ncDpmu
hn80HqTWcMYxDB/+JKGsWHKFwPqphwQEY4zc7qYwWFovgdnCSiX8WzE6V5dcE19P
JlrR22nlxBG1zSE+apPJM6KO2j05Vh/Vva/QjC4jekgpjBRaKiU6Fp7JFhFUOBCj
OWadKAyWS6GDA9sxgdi341PX9iFcF8sYQyYK35ZhfmyY4h8QlipFK8mTUonG47fq
u6AVszL42XdZQhO4NDnCKL7IfBYBqM7d/rL5IhE+XyL7eWP3naSthRg6sMFZN/Ex
kWPjC3Js2TEk9xLjyrBu/9S+gMTZmXErJyeCmwtZKlYgC+/2cBrjlFPNIykKZ6B7
oMNDS3GryoQIOFDqKxMqRJEwhrbUGaLtzu6v/4gVi3SgUKNJ14KAieFkc66uK4jD
6baxfD1vqhVFM7GJpXHmkAiUc4GnyB+g9Ii11URmO4ojnCDsvCSb0lKQNPjc/uqH
XBcksIyCswZ3Gh1HyvR08UD7shIhSh+34HAYbPE5Ph2O7YP02hVcQNWiQR5eW02B
0YoCPuNt2Sn9IZVYcfrmCCZ3ejv73J721OGoYACfMaTeDtSRNoCYwmbj0gOQtsXb
ARuAa3s2jbSGZCt5C5Bbc/tQgmRn0r16d6oQLEaP5vMP+qPtwvXmSSenyNvx/wF5
Hg5gkpRJTJ8kUZxsSv/8Y6xsR8ti/onG3sbb7C9043cfXSTfCwXKvKWM4tWK+Yq1
yxiv8F/JRsq3yyG0uAuSb688qOpHL77wY3eZ0xCbIOGMJuUO26k/o0Ard5CtBb57
+gAC6W5EP2WlFEZ+SQMmU9te1IUqNcWjj+8CIGC8CVGa3tIdc1FWPvRWRv2fbHxo
gT598gOYsYhj8uZ34DJVf9ba6VTrrzNPIoUs7x8tFn0DrZ8cos8u4FlbU684XwdS
UtYFEryJdkMuhC9KZXgP5xEwb91y53ijWdV6pA9JlAjnADTk3vPZQYHh38MfWMRZ
iZhNHEvzXPYZLcD6M6pBU86poVTbo3Iez/tVz4aiQ9HZC23zEl8Rq/rw/9ibG3Bc
m2fohL6LLLJBbJHWgv/1zjfuZ923WW33h1982uydaXPTGE/Eq0uKBA6s8hRJAuSS
jMQsZhGH/0uQRXxiPnpHnJ1APvOI2kCZzHVOSB7VBO1zveb6goc1G/G+6lUbRWcR
9qL4STwW/efPKEo3igoI7iRxdyhw0zapavZxTQV+wqB53GWER6hRxkFiLPmuszDu
NmwZFb3RsdlDf6Njzq8CdJ7EnKxXmyPQLRVdc3ofJATmjzz4tzB4HQ7jli1WAFZs
3MsoyiVQH1w2nBrIt1PGUlfrwPJ9C5Le36UW9MDv0pGp9JxQE3UhxaoYeBVYpTdz
A30BhGkASriMhTsDexu3PoWBqZ99VPbS6pfF7ivEr+ib8c1aJhAkFWWQJoIbuGs4
RA0wj/uLCCXyGkC9fixLrh7jiFcxR3nacHntYnEkcyn/7B0HSKGK4EShOjJ9/LHj
nnbJyH5RJ7sOtvr0mjq4rk7ty3eqwi74qY6ZnuI40Jjgq+COZRS3DKFd8ljaPfng
J01EI1KOlTOlOz9QhE+DAK56gqksC5BhrqLOdjwBvnAMO+26eDiOvALoEU2XP7l3
84QCHmoXAv1nat6M1ITPQTWiCTKISOdKv7rLiAWx8uh194BPJ526f92YflD9LY0Z
N3x/C7usidviTh7iUqDZi0xTbl/ga5ALHcyKYO3b0+KXZkiassJ7aIxAU1da3bW/
G6FZO6DjZbO/KCohgnySO6gXf0fxZlMqYpGiKhCdE02MOLziOeIjbFBQPfe39Bie
P2fz2ih6JZ1P2o3sgBXNKTdsFxXQLHXhH2BL5/m9kCE/teweAeYm3GyJBruwjsAP
DYACyEB5ZlvyxNWvZooPrEiJOXcqJlOBI+CaC9+diBTMceZLYyM0YAVfO5tE1sSH
9zCbBlbsf6SXX5AonuIwFaQJFUrraLzdRM6yDGhjl8I4AGSeFrzw4pm+t44j6ADQ
hGe8DFILIo8nhk8nLNs4oNj3fZKSL6FZyDem4XVNOFsVSPs0EE+Ke/1bnKhGObUv
v0Wnz6VuhEiLJ+gLTsgYnc9GRWTzS6NSsxephvYxsUh/GjLVjg884qMCNaCzEcC5
mghaJUkbPLOHYz+BZa8BI8jqyMSuKbZNWqaNQw1b6BMTJd2TcXj2s6R3Of599zlx
l6vdHvqyq74DDQKPA5d6ZIzvVnkYrSdUPs+bXPfyZ9HoscIGcjboVgjq4PUiyMYn
+pQs5siLcV2NjhQ3nRxfT2UNGS6IF6GaYQE/B0Pp6rExUYsAvuoHx1iwtyLcVo/i
n1Tp7lCd3EeOmhzHfIkYupYu8AzzfDIvGAnvMOgsvriYbYq9TYucJddIDMV5TJYV
mp1YuWCnjdBZsLBgi5oUzUe7Ykgo5Pp1fax4HQtAkFRc4g43KfwVJinvHsFrNb1Z
Jeym6M2MV4Ec7ArJ7Zxit+4iuBfe1x0sWAEK9SeezSfydUOzT3zEqUgWzeag8FBF
QdDRDlvRDjrJ0xYKqFk85IijdssospJRa3SHZtUYQ24KHO2F7WzYom2lzn+EMx4Q
yIR2JAoopBjoxGbLMDcIWwBcE5rEvckfdnovamqPOQ5ffcImGpRaBBEf7xBl/VlX
C8X1Mffp3Jvs/S39S2H9AbNEgBiSK2pudcE114Y8eM4MFWZZwTjn3EEnMc5TJQVk
kakgvOExDiTBtOHk1y4C42o2bmuQS9XOhcf9CuuI+UzN3o6PVWOij/QjP3jw/SeR
UL40oT7e01vYhbUERldfDUTBpHM6wOp8zZhG5nP1tUHQ3cskuyKXdcJo+fTfRGnm
aURR66oVRowWAHmFDx4XbwhuzrTxS//6qLaFDtm+GY+f0EdQIGDY9e0DbD/6Z8pu
Y/PDIsbF/frctNK23d5eqeyifMu4bWO55HHlipjNB0XIsxBTFsse4yoeQiQhGuAn
XHrfXOhQcOz0Z4bgnpqggK/nSeIxpV9kZ0eIdj40pV3RMSUFE6SRwtOSw9h40Bid
5+HMM4pj8apdt5wpRtJR26gP+bozeaP5m6E8AwM0ZPYUkTbl1lfKcosSrR6mQyI7
J2Xk0S9BAWySPqnXDbxKykBhOaEaZukdWYFXoyFiXnG02Dp17qze301SQF9bhYqk
wMjeQ/eHsIMqEqCsSki1hC/H9ITBw2cECuB36eXgkwnQmNO63zzha0XcUJtbP/ND
DZq6Vn5M62zP+6ipwUdc0nIILBVObB8XWWQHgR4oWm8GMBvgc9IT/0bydeIMN+Mr
MyulnWRFPiUsqMvHCgAiBBp5yJCSxzPiR7o7FJ083as06aKBQmTFCjleHFn7hTcF
RQXsh9mlSgrx1MxAy2gb/YfK3z+SKz6eyMXgVjvyJLhNac3xIVZLLV6/soxzIOog
7+AIRUSDkXrYI6eDFu9+lbRPafLIgvVs4w93Dazl0WdN1i0F0Ow4AW/8fy4HJ1RM
1wzpniGAn7opsR04sMCWgL6Gt8VhcFUhQw38hsEn4/MAh6JboNaxAZE33+4BhPDd
1G4wzf5ztXZf2tg9hhfEltacL0gJh3IK0ihJwUtSWQsQ3iwjNHzQvOHB9Jws3LyO
mPRkULpyeEHDKCB03+EZRLBEFwzqorM+F2mxwVtsEPT6Z/P7j7hDKKoyCPNQynri
EKklpSCHc7rrZg3pfTzOBLpPG8afX2ZLprc2tHCFkINeLqW3CQBaPOSKSahRYCSY
54TkOLD4CXrLywXrhi0axCysQCINe4MfZ4YjTgmJHEpx7hF3OoegGGO9RKLAyTBG
IHfuK+wM1VglOtOQi+C2X6dxHaqEL+ekkqtOjcDhTJcwu+8VVLAF0y0FS3lhfDnl
V8GkgnNql6CitfBzOEbkX9Gw49QEnwnTZUpXBfWNMz9Rna2DJ6kI0+MeL+zKSWoW
5nY1zTWtJqHl9PHupha08o4H+CWxT0GBXjtSJoK+Uo9EoBzMtmMDqNDGWbwTjkUI
tW7Gu7b6fqd4nkFrBu5/k36/nFemwRLkhrkWXLDGIbaJOdzvfRODcbye5tuy+byU
WOaOVo5rVs8bdf52Cji2wdiF75BSKFvncfWd8KPEl+in3N6PjZKV4sXlWAzrCmVP
IXO0UzgIj3XbZX51Yfp9SMrZ6EMCu0iy+GqPdscGfZnOqTBSvwehwie605rD0uky
D2z9Ed4+TAQk+FqREXeBQo/yIUd/p+jBQrezGroI3IT0aWh2xZKXOfOdFRr6h6gB
rgGHyd3Qff2e8tsjBMVAJdfPvlJfY19+kyAs4TwJPnM0/Uov8G5j+os57s/+apBJ
79m05TcPduU5x2NrNRrJBN5fmLUisJFSOYMLZHrnslQMqkPqKc05rBDWWWH6FjBy
vaxaF/VkGDPwWIZgl2IvmFMCZcPMErV+k/ASsi2ZPUgTv6lRC0eLw+F4GkvjzJO8
Ya+nideslVvi5EDaJHo4ST9kKECzzJbRJcmiCF/KXYiIGvCrGR+Qp/XOcdZgkEyb
s2FdPQMsh2sv03+NNRg6VcOvGUtI1iCIbr3g2Il87Op4sPjeITwKCb/+HpYzhdD/
xF9yjylH9O/oepNuGsOD4xhQ8VSnAP0VubEK6OJ8R7b7nYSqG3TBdJfMd52CnXA8
IAlJIEuktZMXK9mp7nPqpYfOf+QAoPYjV8JUKU5z6BN4P2Tyy4nl5htvgeuvs5r1
1+qzzu6Rl2T5P0eUqrMMxEBlWllp2IHiQrSsbvFCigDrzdLo648L6a27drb1M+f8
Pwa9QhWaauq9yUkgFDvogOvbKstNm6He2Ghkn2eqDu+fhM76z56LAhQgNUU/wZBi
3ZNPIuwnftBsv2NihEx73nuo64tg1gIFhmnJjwTbaT0rcZbS51xBRlNNBTQbdvTW
t+aAC8FAuDPij1r5H/oFDHxL4Q9YZ6DRsqVeIbUYklgwHPQpkcFz2xrPwxEcjN8x
rPhpuws9mRiMekIBTl1OWSK62BZcmczOxkleA2xvgl+ISB3uex29Rgd3LCtViHxx
OfNdgn542qyqaHWprMGR6R8z880+OsEj/u1EL1QqCtb4XSjuf+BaRAbBddVUSpSY
bJsji1/N1RMi5E4xWhRTI3BCW+fAxnxUZ9bfLrh25ji3U4wVgoVPV+tn4vMVnUTh
YPfswHRpFgEb7ojqbAxG2nq9ScU9dwu/YUD81TX1VHlEC0FCuiPbr1YxkSecXjnl
EFHulvQoSiMwOHPpfFvYvw6chxgWK9oJie6Jmda13p5gAYchqFKSU1cOMKklIVv4
lYiidZI2pHY2IE46B0N/rmiI0vIILW7HEPnqvIyGg1560SPEfIvSYm1PX2l0IKxs
2PIakgiahoSxWQkcJA3AaFshVwDBwO5mWKItEjV5dj1mWTB3D/i4pbPmHDmFc/80
zAWPK6+Tv9++Co30wTjohrlQkaKjRLAMN37osB98O/GeQ1opCqFNfWhk/6tlWmqr
76NiYdZpo09qH53rDVTpsL+2WbFiHDTT2xtoWbuw10bgXGBgYSpMn4arFsebdr9/
FPDKJYAyzColT06H2FOTYozFkEpE7HUwBfS2B9z0dOn0YivIVIY0MjPqSaYTC2YT
2D1am2nUFvJoJmXXDjCs3gbzzqW+pqbk+02UyqeZDn6r2q6eKMQOlhbzUkICUBqN
LAaLeV4qOZOWR1HnBm03/RZpe92D0sTXuZ/btaIL3i7EK+w9nTwTMcp31UvODySf
wIQBb5vKbIp9CVWx6djs6kraIDN5nQoEQVt107sgX57w5xaLeHP/nKhMZN5kq9kK
3cn8MW/o+o3o4AiykvRaBAnNRwUxiI7Epg1jdC8Sk2AsG209TKKHSqGWlYFBvRKc
BzUIzuXSCCxF7aAwNESxD4sKIOeRmTXy2yWAtLbPbI0Z/WdsSHDmWCeQxZFx++hn
NehLoeaX4d6Nhq1JLaL8VJW3OTzXd05ghpf1D/Zo81Vpb2HT3Wuc69rfVAAKIqXy
Z86E9kkSudHi29JHDKD7HZ76IYiO3lg9A0l4X3VbuuWuFTy007ymmtWfdiUoCaIs
aqqv+Jrgwa7JRSDkpnHYVBpDLqLjWEPD0AwIi9TnffXSSFadHx1f+yMPCB4bpC5N
uQWmXzorGdBKGM84LqsTxXebXuce9ZE9MQ6vmEDrjJom5yppjG1hEG9SwmonCAFW
6WY8HENvt/pGsqzeiIeMczdMizazKXS1CuDveX4OT0KIVBQ/a84apS4IWvUiCRSx
JFnwy0HSkFZQEhdcFT/+I3nisl2yn8ZeTm+kUzd3dPGEZ+fBzd3veUTSh+hSbuIz
vni630D2wrK9iYwdq6+BrCCt3G3FAOqY+6DB67FcZVblsnbnjywYOLGGxrJErfKK
ffoaOn+YGz9X2Zk99Rlj8ge6/E4n5H3XklXeCQZ/hZtuT1awTFY/altsHiZOMpco
xjW2IfsvIHTzwtrlU4/PfBqbq3tBeNsAKFkazWb26APY2jKIrHeP2LdTNlwpLMIM
TaNLinEFY45DzXJEsMpUo5E70R0SfdSWDbryfirE8nxoolFxCmcXC2QnPFDcBoHw
HLvemKcen7JqQxGyaYTGcm7oPv4erixaDGdZlpYbkd9wXuTF8pKiIvQXuGGHWr6v
r0rdWFcIh91SMBt8B2GlhWllXTscxc/oC9Qoq6DlQkAQn5A/llL0Gp/f12vpjYd3
q8wrJmP2cplY5Qcr0fc2C9C/EPRkKECCi8GAAKqsjM/fr2aeZQMJUXmB4Qbhpl9T
k2UT5dHUmP0HqTBT3kq9cGLut8uiJMKVeG1anLO5duz6ULVQIfj6y42UW0TF4V/R
DW7EvqUJadcOicYiGyZmMIIC09/Le+XIf0bDgUgEPtEoUmOLE8kcFN63y/Fl8dUR
N1Al9Fc/8vIxZyyxGndVk/+j3Q6yG0MiuqVXRkooHXw0YY4iDLP90Vl+P7sAkPYt
nTSOg2RF5ixY3OQwK7VHgp8ILlLSDESU3h57zWwZZcdtrCeJwDumRf5kCZ+lagbH
6qWrh+S33UaR4QJJZnJa+jhRRSpozD8wJ2suF7NY9P2zKA/LJ6b+MaDbJWsntGt8
uHpGnxpsiamKeBqmUQx4L8SSx8kXdA7Chv18H8HEmlmE24OQERM9iyBBqzDRdnVF
XEeZQVSD95EdIpWAEj4hcURC2EFE+OT8+vMxBtDB74wN5m9wQd4FwwoELMpZ+tYd
Sd1D7tNC/knGvSfDsk4sOyySjAoQ6pQzSCm+WzIbj0oAdjQ/tmERjd0+Eb7RZYzQ
eqyaV2sXXDoXa0bck++tEEwPBv5Dvq0vjrrpgecf/kfrXPZTMZUpQJQUD5Bcx10w
IUtDRZII0maXYjhe/UGs5VKLHaks/Ys9rYuSNYzAl+oe83ZET1EjcDckFl5HoSYd
oVkRrf3wh1A0q1bp9lfGZ+jgGs7itohN9YMl8sgXdOGTP0t1nUxoCDLLV8dzutPp
jpD4OjuveYntFjJmSSIJMNONOs6vku2Gm5N+vD/znpFVtsqUcVZ/xps2Z4Ye9J3M
UMmx8qJSEiQVRQGhYhpcUcBNE5YKa9AUDzpnUyG3sht9QiKU2F/mCpU/ZaLTbrhy
2KTSj8JQe/Zxqx4xCYmYr3xC5KeTPl4KFqGV42ojkxYMOq48s31HaJwxK4l/Eca1
lKKJI9VCduPvXv6EQ5A7OKF/VPNlyUqi96W2e3IlSciVisiGmlr1FKJ7/DZqcJDS
01JhmxCCCHQjVjMGA039JUTh3yt0dHBjxXouUpKO/lXQqlUUJ3xEsOpY/1rQL6Oc
7hRbDR664eZfIy7WNlU7WXy6+DKc+CvZe69jrSAPQOdmkp5lqj0nB786lNWke2MD
LkT/a5CMkNx4gwm7fKUt90J4HhsOm5sMMQ5FJWKqaY5CU+zhq+ZlzMAEzkNs+phW
BIo9ZOREvtdLvkSkMM2fQiErMQKl6r/6d2zQQjVNr5F2QeXxv6Bzt8MtIyUCH1dW
769G2r/gDA44YbH57hPXMP+XVUwRJC+K8y1C8wCkSh43BmGmCorhn48SCLars9yF
GUXUOz0xE312j/gXU6744AJx7uMVUmM/6M9CaNkYzObkLvi173u3cjQVirLYo6bE
io+wmLwgJ6tfgm4A5RdHjkhTv5H/kdAc4MagrJOYD+0+RLekcqU9BXHxqX01NOzY
0caruqaUIFnhXwk4Tq4Xjmx1Gf4lD2YyEfgNW+BFBCKYMhfDmTLwWvDEBR9vFLpd
ikj54J+tIRBGyKoRG7yj1mswZLLEw8GJZD/4lrI0a6itsMEQhC4LnfC7DZmc/bvb
gX/ylb93zkWY362JSHmurxmb/TwAs3mm1egdYfdTikQqcJfHNIMp+l86PrXOBfin
DjzBEOdg/rI8cKXPZhwg+rTynEhaiS1DezAekJGcaZZYwJO+1YYjoBCrd3nxFmqO
Ysejm3GBPUr1zZ0sHq+ASjld66wyWY/qdZw9q8GNJUi4epdS1q2Pz9Z6AxW9oCtA
E2Zu6VaaY/0Ws8nsF9KQa74gieyMdooAiXAbNce054TyOup8E2R1EKKf6982IsqY
xw16//cEsr99CaIidgFsgq1FXBTyMESq6R3awmynho3wKv55Cupp4IuVXAV4YgHa
Tf9XkjpJkr28rjERToJKwPMm1FTOLdMtuWu8kL09D2C9/cZkaHZN7i//figrNaSZ
Rw4p3aV4Zclrj/l6QJWk6CYgyaAC5+bovD6M1FTUrk53DZ9i+vUDX2hSUJu8mmmg
SFawAzXvbevLJrjEeP8YEV+7SELTD0aw93QMGWm4NeJDzF9E1I2RoY8lyCbRCTfe
YLHxRBF2c4+T+mnNlRyO2/MlP3G1I9bTQpH+vO+nuurx5E818WgqnG9Wn6ZCb09E
/b4kzLfAfMbhJefTWx/fgTpFKLezzeNOGB5FgKBm0DQHKlwXXqiYLK8GrqATKR42
H/YbBVO6M+4PjFKG1Zb0BfVOpDoY8J85V8HsRpqiiyq0HzMe86Lsixjbks0cCDa3
N3S9ZwbzzBKbKyWXBdVwlMK9q3TXlNG06y/kjbCd0pScfFM3vsr2pb80r5aAOWuu
YBulNIy/QsYeCtDm0Lfmos8RU/FWWEh928Cd2jbUCeDAAIt7h3QQw56DZhrI3+kW
6a+7QBOMy3arVaYAmjlxhaFht9dEUCX20cUEZqX5Fvb5L7NwR0dIyoIs9ltZ60BN
Sh+FMKA2x7GNOA340Q869uPj4xtD7htvb3HZDiWDJD+g5S+eoniowU3ItUiRAXHO
Qx6EQx64+3fSvJuL5YIlyKWSDszPsqdwA/hy73IZP/4e4/qJ7Vkxcl0V3bwiJUW4
cWj/inMk4Ow8L5CG/ZJwJIN/uBApXjxIS+9fpd6NTvrnnYYGoq9zQwZab/ja6LQk
9Loq6ZmZVucgmANgsyJcQ6vzBwDrwBvW/C8ZWDT5ZnBmHv7AcjH/KwWl62c8nsrk
AQmsNNX+lwAIKYmx0SaRsrkqumOcsbTNBNtsvDqTV2ZzKTEs4v7Mju1wSPaTeDFH
XUsu8xk1857wCY3RzUFMtBq2LVndDqfoXKXMMYxxYIbf0At3HJW/gwNh+SQcCX8w
kfuETmOEHvIZ97PekaL/wpPUSk4NCE73NQJ3KBQr4CzXCW2Xb1CqvZn/svb6sn77
Od7HEwUAEnFvOqooR3roBpVM6LvW7K0rqYp0Xj5UYlnX1IrNC26JSZhuyKOg8CR5
SsT7YWuShLGg7og4m0WfftFccoY71+jcmz4SGWyc3NyDtFR/jucO3KqlZDXR8Owb
tfYArGfmG0RyKrawSSSztM3v7XzD0eqUoFy4u/Y00b0et3v48MzgVRkYqmTri2rW
XoTZxAvzn3a+xqK5C4F3WTxc7JPdfammU0YVlhCFYbEBzswEYQD/Y6KZtZ4qfX55
np9QjqrTolZ9QE1w7P3or5miV/vCutLjbRd+c2VVp+s2g7d4/N11GydsYT+9Nxda
jnmwUBVhxPVuBuSyrAf6+c7hfAKTtCsjUsfrytkTvvrUw1kJD4HYJ6W1NabKtrSi
GKFt2JxQuoGFYK45uU9wqKRC1056BKZlwte8cqZxDQQDkSRzGw8gf07Y3JoTvr6r
blWTbPRInzzWgC3ijX47zMYIZNU1INf1oM22wzTDGNGFYwSmCpUDRMGjhUCudx0C
QVY7JXoADxdOSoarAY2nc4g6EOU49HB9bNLhWVfqcwloNeBIKbI9FH3KkYwnCXgB
0XWrzyLYV3RpfkfEAxGWK2CBQ+bCNgu6SvT+HohTaLUkh6wrsansvcwnvwZ/MHCC
syhvwc2nM8jsbA1RsaHUjsqlcNDvIsJskQPoYcWmDlwdFrJo1ZY5leAikr35OjuV
2kmwKB/vsmK5bP+Ryhy+2GzlA8TuJmJ2IvivFAaJGNw+HYI9H+QMKlr2pStt222Y
PT3rjCQ7XK8yDbqZmgbDTRMgmBWg4s1fjd1s2zSOXO2U7n1OW3oEfKVIc5AFLTwo
Lgq2xH8TkEpeJRc/Vkv6h+oSaJfMxFgXDl57oUex7fV3yZNhWR8Op/wg8qlhuBn2
KNt+eaez6m6h8cikk4cfEfES/seq8TzZzq3W9mjK3y6yliZIgeAa1+ovGlC6MtTU
9kBXI6ubmmZtrbgjUVusIzGqCZA2dFuPCyZUs5ay02vH0SLJlzciao0kZwN2Tur+
DghQoCPRahl+RvOxtkFhloyANcmXdriqTzkBcOZTOl1JiiGT26U6HQ9bAastcsU6
+lwvHEyH1ExX8M4vuoqpD3YA2MHoZ7gPWkjrFwhTgggy41itD3934ooXApFUyfSe
/fSXj6Dx8Ccb6V4DrVAUspDV1E8iemb/Im17DaP4s02NgsUfd2FDMoXQ/NGP4hyG
40OMrQoCAwdbPPOegQLXh5jsSYuQucxIlKr/Pt1lY1VfaC2B+PRvhtrLGSxjE1lP
PCMk5WNF58RyxToerYNrKbKl+oolIqvzwc8JQKjc6SmebMz8CPxbIAPXMWAkMSq9
kk7A1SWMKiut2GaCCa79nEcG+CZ3ASZ2Kmg76mBz+ii0zgj5132ODdxOtVfMYSfx
rKzKRL/fdfh9GfaT9oH+qJQ2ujUcGCWL8VJB34Fu0mKdDU4KbUA2qtbUUCbJIe/W
DPco5+eW7qDzDyko+8dPwlPXIdVEpO6R6FvLJt/y5ojtWvdLKqhEE7Iv5X/aGi1D
5/SGZkoR0BMQJQdcXet4+uR2QRxr6KdmcMtjTbYc/l0so8m9pgypDFQYsayIvqTr
620Dox/Kw3uxT86RQbOHk2DPSQ7E13yhHI/QDctnQJwnlZ3zmwSN7sb8FTJT9qM/
buNm0Vyuz2CrOA6U/B6Tr1Yt5JDjFYdbna0YG+AsLo1y1YOhHdnyaDyZFhz5s/HY
5nWnvzycHT3n4nQkJdC9p+Ju5M/WZ/ZGSDw0vPn3pRdb6+iKZRJLcLyt0f7CGDf7
x9cc5rcxHM5vykdp6zCQtD4BJCwxclRm5BigmbP0BtvLtNAdvvLB+bg88Y0rm9AW
YxoIlk2B9+CcjxKY/YwvC3GjXIEsLiujUJpgVeS/T1RpwL6ofa5dLMbrttrE0w6w
xpS/qmQwocHqTlh+oPsVyKmy+cQDgaXAvvShu4vpLTD0RAvjpQoDzWAu0oxflzAh
j5urGB3n609UvJ3T+oWdRCGYiHUUJYG7NT/XMhYKDYVq2slJpcPpPBel9HztXjE2
uRsE24T80YmHQVkvdDLua7kGIesXniiv0ePi8kNwUzDGwn5bIelbwm3WFMI/BKqV
bNjkJFB/otlZZzJPwnjpwO1clpbK9+H+kqA8UP3C4GmgL9tQDThIS4sWKPIp3y6w
EVfdOZ+sC5S2IpAWULWcmGuqsB/E0b4hGcZ9x4DMGoZd7RZl0+EUrmNeFwvEI9yG
+rM0kQr+s7FT0d+o08deqxfJtplaDPWBtuAg1VthX5u6Ue1aaVDv80+LOL31urfl
xppjHxCtgPKtSWQb8+5IVeewx6umTGNSaof0ETyRlqAKxnCpvJZAhDpZ6TFKXV5Q
Rd/lmzfZQeLIOykOo06aGI9sdZ6bHHxnSgYGnYjK9EfPwMXVRl3ViuWobHpQb+Og
cnZiopcdHZvJEnIM+vvYMg991GFr0THjSEOX6+9IrKhJ90qXv+261Lx3x8RyHRWJ
UfCkeHSjxGlwNQie9mJcplUS8qsFNqF9vaZyochlj5NgbvtPMrILoI2izcbLYcIc
pDTqQ1qkxCHYA50YitmXlA1O0RAUmQZmGL/P5wsizKwc2tUgrCrrfGiKH6bEbEbH
hs6sIpMxECfnBFoP5eAONm4yUwLWL9Te3BoOVuUQ48AO7HRmKq2IAyNmkf64UkAh
OIQssjzrTgizJz4ElxUE+FCJVgk41RK6tC5PgJ67RzFNP245dSxy06OPq+/jRiPF
MZL/qbWLz6xaAfyXA8jtaqfuIDqgonzlvpyctrLbbu/Z2VclOOIj4N7pOFJD1teU
/NvOZKM3fIXc9UDacIFbmhhwPWtbzUc/tlxV3Uh17EghsZewUCJiPccuhWSx8xDD
MvR+LMG8jBGsZTw9zRA858Pm5AX8+vjhq0GsZhpIzmcFDTYxOKg38Y6NgomUk/lf
aeWXQ8ALCcQp2Y5WYPPEDGHJCd5hyJconr5QwYt21axU3aW9EOBgGzequ0+EKqCD
Ilkpp52E6CP4N9o/0boa8SaNPKew9wLqTS6K+/HEUwcQyq0LDoak3QSTy6sCFmL1
BRe8q3t0cw/wCbm0tw/NuLO2VSXu62PY17xU+WseSoE2pUeIm3k5pLELOGaCQ1nX
MCAfWw8qeytB3nXaEKGoh1zp1lG7Nv2ZtBVqAf1lZ8n8epqqr5Vb5oP41AgHtkei
vrcijQX860Q+Wuw/Ee80vGzXYi2DAhBZLemYc1FDh8eM8Xs2EKGBkPZ5pf4XSJux
+eUxrJus6UFHpr02rgmpQOI4IlKxl0cMoWss4Wc5f7l58QUTKstvyIIRzWe+fOv+
rCF58VuQdkNk+t/lCr4pTcrdsC4NDDZw1Tcdeax8n1I+yK1OG1pBCF1sU0Si8g0S
PWqM7qbtncoyjMhinp/AmO12xmLrRaLzPlpCFHruXEEFBf7x297GXLrb8znwj+8A
vL+DN3J2B6g1q5W0cWwZQMUYuS8mcVxDYd5AooWb06XpWe1DcC5BmzamsCeuagBl
kF7rYsaTK13bD/RE7jd68tNNGbP6V4+qs4NLvQlduPgQ+OAfOhCYKk+6/qVyA84R
Ao7Q8on3tOfzj2BMa66O7Mq69sFGqB4OtSm3jEkm3LtTO5/ZVOv+Zp9mkfOWWxJm
cIkNt48CSPaN2DHeAiipbJRXjtresC+3oeahr4/nk+ISKmsOzuIurrHYhe1MCsaF
wMNzoArEu5jQN6kdTZsN+8329/z+/fPYKDM4arvFJYFUbBTBJnUAeuwj71hPWbpZ
vR/YARo50TzHCXW9L8JYAHkJ341JEQS6/Vb1TbDeS/FwyZzTn3SRoM4sBBWNHnqj
i3AIGXFlhobh/tpxcH6SuKabGBPtWmU76jHRH5ha4jS8hdfXaDAOeZSt/OjEBLf4
5HEFErP5qOGHp81kB2QGk5gs1/9B3pVYClDWefBYXJMM+4vM2PwypI8qFJvR/TyG
53KGWLnmxF2DiPXQ8zkqTwfd3DdaPf6oO0Wg/7H9X7qJWpfvySPvjMakN4I65tg0
UOa5E2DBhRSLROKeg6fI1Ws3EP4oucvP9okZuF+xYhC0Muwbd0g0kAzodbss/NZl
omuS6DwRBdJtidzyMO5haU1j3VLdiAzZGjQCYP6mKGpF9JRPRYPIP3GjOXzibsRX
mcMbQNCna7pdMVHYsy59eGR2ywbMGeBuuohkSNSqct/IGdk0dYtUt1sjFJiuT9eu
MV2lch3HtZ7C4N2G2X2bvJKZdBw506ad6VbxpppLcjyjrWwWkSHTRux+/T6+Jet/
m8wkjV6yBzghIv9MWGawRW/UEQ0/ognxbyYjPL7v1kMlwB495on/y0SR5ki+q6hy
QKVVDDNwkvB9gfgOQ5QwMJse19wPsS2dLhAHiG+xc7Sjqkw/zJ7VJpN2OhQaWj6S
ur8N/T4H2PMqni6KfIE+uTg+uiKa+I3PxlkCDc1GrXJCfl9quK0wTSzZCmRWEiPg
G9dEnv9L1Rl4OnPEIPxsIN76CtNGJdZTSZMvlxhAMryFgegTaBj3PlLIOSFordmW
fHHKqRFg9khtSFhWPjEZ7hbZH7vZr5MUT5TLOSP/dIr+AchMAzk4HGbjbeo1yXB2
/qMfJIbI1BICnZZ05tn569DRicGYY6I7+czs3GF0GJ1Z3GAXUMhaWnAa185K9IOL
mJvVU6mNPjV2EUIH2GKJYs1+7341pmF8ZYJ19eJsc2xwqsuy2TqaU9IfC4lMTZQC
75K9Hnz9ITZquaJhCg9m29ZXYZ8WoM2Imr9zA3Y+um2HxnyQwOIq7g32cMecOanT
LVCf0hTXkVS+qna/iSPESld3eifg/rF3XZRd5BaWEp18Zq8FUcT1XdCav96CpLS5
wls3hPQYOGnLaUE5YplO9M7xY34/5gsGtVPMwEYGe7SXmanNwgwyIlHEiQLSwIqQ
FOdwWxj8dSIBzJqrq3dydn4vsNClg4YHinfY7DTx9bFalbkW0DqM/2hQX4BY/dLD
EzMWWz/Sd/zxl0Es6KLkVhqQSLVXiAlhxhAHogC0d8K4dtZ8jSos9ZQCt8/oc+Ze
LL005fevp5Tx04yyBcUJEA3BAoB4Z3SZvAFrOafNnDTr4qPm8u10/J1fdCE+Jc3G
pgjQ7VDLgcBvo5qR7pk5ejXenFhdvCTKYa3QKqAYZd+H0t5W4xcLDPzg9hhvJX8H
assjfcZI3zEnAaMIstX+9ivfzlgQixZLc1pJ0neZx9HeUcvRXZPpUZ8OFe3jAE1Y
18V902fjaPXtB9ebiARRt/r5UliRMKlOR30rm+46mXiTmwkNG1MCk9hpAXp+qofY
VKp4ovKzgt8VI1zeoVxz9Y0naxw9DC7gTdQ0m3ecEJYiwOn0TzkgzFX77UEYBIB3
fFtqW9eB+8GRq8dub3+VFubEQdcj/q+fIzNiBQeNJenRB95EKkUPJNWgmXj87Khf
NNK1lhvHh7wswVWyPdaCv9K72dXCLm7EnipxLw6tLDavhFK47qCTCliyGGrTMi6+
yNsQJvTcKkY0gfSigWb8u5n1mco0zR+GrBLL0nU5InZXRA0h4OJfEqkOwbH1hjtP
VKuyYALcFajCmqIIBdp6zwI7gohUaOzJKl1wD3j5z37bdp2em0hCuR6oC75KUhAK
SG3zi/Hd5cj3OLEV64D2T1CK3CBEZgSve1eeKHSJnSzUPeG7cpywmz3AWEOLhzdL
ceEigjuchhEplj04Hkx7/58Xyx74/XAiitaohMJ3dsl4391an4+QEX5ML7a0JIyh
r/dFHi6xPgq6/0J7jB9564q36sptT7s6Zw6jxCDeH5olbHPGHpvjRs2vAHH0R+Ah
MQd23iaMPPdEnO+X/TZA1y4Gal2vhIT/daU8+wsU4frKYAWOT/NvdWXGSlFcoaxf
UOSgU0+WRQuCtt30Wi9KViPuUy/z/LrTGA7DCG9ynjAuIu8bratzcbt4thpcz1JC
CBbZz4XAGabjGZBnSKsLTe5j1698d4cqQX0jARTxIvjJJ0rleV+N/wT0VXIXDNnE
JLcLtx+dbG+IMtG+vnkh/mSsWlOtNnid7QRABN1jzt5AJJepiFuIWpS4iUQpyd95
t0OU1l0EOkoAObAJIobyQsxmnX+0Xp2omkhMDwzxVuiPRvpPp/dh+L+ktknpiKAc
uS6v/dqpa9OAPloPTFvIAiSdizcRVB16b/RX+ThRzf1dd17mlU9rWbNsxrc/S+S2
8spPHTuvdJrpm8rdvtF2DbtRX5ceKe1jL6GSrv7LMoEofIapniP78k8w13qfdcnY
gOrxwa3WOsd06MS3+YD+yVemwVtNzzQ+/QMtkkPNY15gqf/eKaAKbO+T+0Yjt/5W
X/c+RkXmp55fZvNaXLlGYSggQJXJu9r/uxqTkAW9VAlTsykOIn6Q2mWGP5yMgcct
1VUx6JJ0ktcCe1GF0gzoOxmznub0sPPuFskS/8+Qy3EbrePjtraD7/+EvM7O4r3r
ewM7aQgSeJjTuyRpSXb1H7KzNhElqcDOubtWwxL4Pw+bmZatS9ssNEF2PRY12YO7
k1vfaH4TqPMuH0LvlejmTfr/QMNSzEJEY9bUxznO+93WEXYsJGZJFQO1RRlouYrG
KmBEK93bd4CvYTtV0aMKu8gylZaWyLenFrhyHEyANjmE8MKTGLbwxicVvMa6DkAu
LXWY7PfDHbHu1sYCjIvJIZgUta0iqgxjV/V51T0NR+2rh7cDNIqmwKWtQ3ANJDFK
dpx+6w4ZLrQ5mhE/X0eXYT2cJkotgvHJWT34PSq8erji39RZ640huuaYYbzmbivP
coGlouanGKkvl7xJJNfO18fpqwZVLasi4lSGohmpJKqnaD7xO/6bwjSIjjphzcxb
ESIGM5ZVqEwM443Vpx4H5NhRJKhtG+r66RYF0ehJa9Zhddkagq4rsLFB79i9WxVK
xVbzwL66P/HiOCRqNdJbcK+FeZJ5SD2vIpWCjvNbufBTR6sK63O+mcanXnz1gn5N
oX40pdfdUxQhsKxL4o9xwg4eTqq7q3ZUCVl32sGEKybq84XYVD2Wi37Sux7q2T+k
TRZgzbML3l6HLWf3WVfmx/6IBw0O/qEA25Ko01T39mSmcKxZHl9dKyRCHrVbwbt7
nJ0lWJaBqTJOi/b5O7O0b+RbErij71TUa3QnZCGQf9/EzMKBatBKR98yD0VOKv7H
y8DFyrCYVKGZT5AkwhYIyuWrSGeeA5Rn6xCp0XDPhtpZIssvR/2shhGsg24mYRGS
lRp8uZwh4ZXCxR04O2VsUheCF9BBoaaBnBzuaj5PVwNXi5vGUjPd9zzMFhsDYpNN
WMl4oARyT67bz1OOId6Nt/1qHXgv/lggx9s6LmsbsIxhfEtq8ACyKPiECvPdhFCO
QShxM2ZqdjHjT1kfq6uxYxGmoFXSUSZwns/sr1Hj9A5XOnsX57exKxJaajovHFfw
xLiqQUmlxYhULtEo+GsNGDG5v3ywytndPTtDHfWhp+ajGbUYOuVnG4gKtRjzcGdv
3xNDlLPAgLx3e5ZTGi96JEix1HgWYpz6ahXxOLr9ts19DdCm3x83pgwY+SyvazCf
sfmpY4hjwt4rJ+ttbpqAgbDmzh+u/mqkBEkxBKTuTTsAnlTKhAJuWkpifVK+KCuG
TJf6ewJAAx1gbQPB8ndHlp3b6YEEesnIXHVxztC/hvh+qfNdsfyX8Ptosx8d0vB/
X0/+C+dVotAB33kLP7IlqvWDUo7ye3GK/hOfu+5g5Ig3Vr/wVbOVBWeD4EJQbwcQ
eX3r9Z5Rl8wMQOMEtDRh4vF7QoNyiZZ+wvqPLYgQJhMCQCeqMTqqvTfSo7dYqOsv
Rbxx+bYGEwOv3BA7Go+Cmg3VvitehY4z80+YabgoZ0OGsS23PhQ690YKw2HM82Py
hMeY1xIIVHwI/N2T2EQ1PZ0QHhQwwK69SqZIHLf3GnjsRzeUIBQgcO3IsbZodZ7+
Pty4+bRpjGODQB4JOci1n7BKIEv0JvlKc3Hi+606YFWPepICtHMxVi0BFAX7T3FH
4SvwKJULyBmZIFQ11GioqBwAMfG9yS1rluB1cIMveY7T+PPyE2eSQ2uASqlaxBZQ
TTsqji0q09XHCYPNh70mifDHa5DcRipnlRNJV5/JWh63q8VmpkgQWSrShQzuRP5n
sBdRmFAhsQ5NQqsdYyx591EEeAPCyYeRFseQ4icpahySb4t5sX6mQCjrciM8WlyC
Gn0A+YxdgBip598KTvbRK8Yju63k1cwSsXiJ6VQiFgTfm4Vl8WjcWCV5CqbPdN40
sJVcJDdSiPSwwBvulxQ0L3RqvYCVZYqQCqbiyGxuL55YW9duHMU6sYoPeqr33Lyg
EjWa3hbgilgHKDgkApzpPoBcDUO23cCBi5Y3HnNKKZPnCYuk0RCZhibhyGld3dAW
/C0Kz5a4nMdATnBcbnuzcxRu3+eCAkox5EepuzuFFqM0q740Bv0VZhqtQRZsaS68
dkJPQp7Bidwy0Ma36ku7haB49yHAZGz51qp9H9nnGYV7X2tjKzuJJwNFradqtfsm
u4Xvdy7Ep+xs5PTwjZIERvcZWGIPfhPpP75STv3cS6/jTqBQFm9GzQVF6E3B7mbP
6zwn2gMmhQGwP8RtbZzvwbs34SzZd8EFHQADJ+0ZBk3ReRSr2S3Ebr9xh7kiujhV
v3S6BubmSdqPpbYF2UunHSyClBM47Y5Xu+QZr3ybfAVBaksdiBUqtOlknCTWcslk
QTcxBN7xL2yecGZoShh/nPOQ8cGtRcL6Mgis9I7QCg7lSNeZ0kstTAHHe7M6kf89
YKAnt6OcZnfiqCWxaIoBsvKu5f8SoTLZTOr0rqJQxdS3fYOYRJpJ1RS4zlUIQvkZ
z014zxVPZeHGbURtTyGPEczrbLbdilb7sfyI42Wz4AGGCF1FjwP5otho74KV85CW
f0Ep2TfkU4mIxx2PN/xQn5pl17PC3EpXVw3OVpcmcqk/n+onsQc2Z5PwK5qJfRjn
bZovT3l/B7dJ6/H9DPADorjPiq8gLuq4i57VRCFpKU01g/tYw5xp6Nh6TZCB8UGU
otZLlHZ6Jx0gbpmRSHyirfjsMSHKNVbrspfI4pa7wkbFfwHqL+PXCbSqqT7wV/w9
Dl+bqNoaGmG4HDFw/nKD/VOoI3kMzh8B/ToI4o+1Dm6STcAu0rre7lpLt99CElIG
OcnN66voP/kVKfb4zYL87lSe21J/M3t5NYZxD4zh+bcdyYroO0lnoz2vVlLr16cC
29lo/VHgP6YccikpEMbGn0BAN1gSj4VOgVQZmhtYbOOrw9E7py2FFso73LVDGgNH
d0myYyYOR1MrUxtKl72nM/izYp/7BFwynC1day1WjjyKv5m8bQNBcII4M3cHCnys
JUieXzkuZ6K4LRUe0tdcFHftruV5z9jIAQ6SLZegQWuAgVF3OobRD+ITSPBooVwK
//hSkFGjIUzVu91nakNZOoopySyH5yC8rj8wgi4ty0kIUwjGu8co4/zWu1aOR+by
CecHaN4mwCBUIqTcScgFU/hA+AcHnOhCzyOMB5SvyZUHbTVaijvWATNBXwsGkF+S
bbO+tGaqT9n5PpjZvX+y7N5CVsnS7yj608MiYksbah+67ZgC4wJ9xan97EU1TfYr
F3p0dwDjxiEzJvaWtadB431Pls8EMKpt08br/EyZMgyw9ej5zBXuWtqAq9hnyhbm
PoQSYxXUVJ+9sKNdvMpA//AbHBfo9M2m5eKs6ZM+uSQzxFwh4+HbbJYzfFjLRlnU
+GUemHUPGQw9cPFbEJHxl0T4cYPr+YcF5XB3SY7GANlag00jdaChadCCO/WiKZgD
rPSbvIOP1fdaOTp/5bqYgtQjv/f8+QMqmcGnyQoyJClNbeG/sixs1iH/1sZ4pSa3
yWf6lP5GhbGor7S72aiZzBiwJTD0+Pwnf+b2HtNy0Jxg0hiwokr1jLsU2nHYX32m
fxj0sfqw4rUxqG9APzWu0swp9UuWWxYjGge0mqg3jhtLdqyyrMPcCjzhGpx8SKB0
lmrfho2uq37h7x52gllnBVuZD+qK21eVharqzC7vipOb6ffnlMpcoobpZzO40wfb
s4+PTBwuDewtxTt6dl89K/yzwrS14s/WydtUrxgkxytAk5/qlKRRTnL6yZSHEFpk
tXyaPlSJpx4sekUXNUIYkjyHKi43CIMFWiR6Sxot0Rx2X0jj5Fu80GPihcC8jyY+
qpHUZ39Qfb5sA1k5QdMa0eLD/TJr9ualEws8JX0//kU9TDsAz/XphUEn7ZBK3NyL
JJWNancAom45pIXsDubHujzROUwco9+wPYe82SWFsqq7/CFZdJDdjxgqxq+YmHk2
I+qOySa5XrAcuQwUXlHSJxCpImuX4z1ciyqtgjKZUF9JvuoAUMrmlnFqM1VeHBCc
9WiyNxgeK/WqHz2pmjf8Gmoty5occuhoRz1QGe8BV9nNpSDrfuW1ZJ2vPjNLGy/F
Qd73RrmRXHMVUT0wfcRjG1GSjSFeEoIyqku7RwH1FaTB05cn//B/w599ksPKFg2K
u5EbYob1/bsdnjpT01lGeobw9XymkP4TD3N/M57HlCZQOkpeXb7vxv1eNtxXLmVD
xfvIa03vC+GK606pL1Ct9jz0fs9cIUd0f1pOxRoZdW/XhThEWEg4Df4Hv2BKyBBM
thuUqxpZHWB5n9ygXa/SLXn4ocfvEhh/QWEOCA+Oa0NLoCYOHpDeXmn9x8Px73cA
pzX6EGKZk9HElDBNUQLZ2fqTnVQpxBGvcPJFyHiKdfHVBH1u6MypCcPDXaNQGNp0
qYFbw1pMDtI2dUboDm6EMsTqI35JVRE2sTwd3x2a/W6YPgJeMWXoYJvI5T0Yev50
eR+/cGw6ia+xWyma6kWzCpYNAV8b+CLRJwUrvSyboUFRdIPpcWmKfsy+8+4jdu3a
gTzwsaxjdYR4ukzFMK6ZNl1L6nTmPSXfzipb8QW55z9jvOWewCFS2ulFkuAPlliV
nL4mxYz0Uv0BcIkw904oc/04eEwatSuX6bdpBsrGd2OtRC9emC0tiyHSA93kWdUY
LYgQ/u9/2BK0UX4MmuyTM4TbT/CpM81SeerV3EKlICZZI/x62ReN97FhLLPTM1Gc
7gD3xUnWA8nHBnOaD5lHgGpilVS/pihsd2g4/E4qUP0R8iVhIiDLcvC+IhSqFQPr
EW+73bNWcfEMg5zF+hVjGUUht4tw6qOD9YQxU/otX1vpuKFxw3c+wx/NDhwtyIZM
K0PAMORhuODs0vH0lcnn8WhQOHlubJvueauHdLjCCGhGO+2YNlZ0E3SZcdoqJCmR
N9H2Q9m7mQxxg9WwXRoOjQpZFIoWP0t1vVMJo8GJrarhftk3N9RGl9HkXY3AMfRI
agM2yZCX4F+pYR+sntpvCm3lftVnK+CJtsv0wKF7o2uxyhzZa1IODODYKDpuLesZ
YG4v8NlKXClJhEjkQjzA91tYpqok5vbB3jpOfBplcqn6g8flo4T2V2J7D4ysPeJ+
P5WM3ZbG8eqRCUDHwLwkbVcW2vdW0h1v+oLtEtU4IgtADo3G4t8tBolY5B7j50Bb
HN2zRCIXvYqrIC7qf/qMNRJdVJl9xNr7JwrNrlWl3fvy76ARFF4XVaIq8vF+ahin
K+P0wabLbMSNx+EcIdYtXfiOXi6iYyBXmGMqjeCN5A52KBkvrhxh6DgdLuOtcav1
p0bxyEAIirosdWsvcWO9dtueXbRUxtaAyQGzAqoWCNV3t3GqRQlUwWyzmHAqm91t
fRhcotqq6/zudve7zCBz5SIXE08716hD0B8yY4bKrAgBhU1LgYaHg2zsF4l3iAAj
/pGmYfxuQfajpQvdsoQiJMxj1ZXw75Dwrc3MlAYiktTVibiziaKcRPE88h9ha3T6
mdBayg5U+NPQPigRhdBlCow+35nddjNv6nk6IXrVXzZw+QFx/cwsiX2e3OWREp3e
IEGa+37+A6qmjs8uc3f6OswjgnibWRqFTqt++WPepW3iJ30d+OMreN+9TeGZNYIt
FLPHw37JTOKTbjrOvtsUHYsku4eDq/5Tu5U833jtuDq+gm2s8n3b0vwyZ3VXpPqv
+xW24GM+f3aqGkEHS4ula39zWngG3ECFSJ35bm8mhyV57Z4ggnCk8ZXPOZcNq9bE
HfZl6kyylzF4DHGPqROxUuSA7SVTAhbTaW/rqQyd2mi3N5LL1N1qTrRv9Bq+oaS1
iHDWHCTUhCwSiUNySwKCdNRDYKw4MCxmuqoTizw7J9k39RcO078kN9cYylOQzK4u
jiGpWtwBuSsEuys+amC0YWEdMmHqjb2/M5ToxtSIRm6D7yov69Pnhk4iUF0w0SWA
7xXTIv/6wYulPvk8Tw2OAXUE9OYZmWxfw/0WNaylya/yDoONB9Bya57pVGOMSMmR
TWGghO8SR/N5DAcJi17kYbQFzjoca9w1O2dnnDWqcNPDF2C0Ed3tVlfHkb1mwnB6
51K5dk1jG8Fy1ElTNkNuXbLZq1ZJVmYqgsRPvV6Yr4vfR8WpUwYFFa3FlacYIHfl
EeiFwTtzgilKZwI7oFOSSYRPe70KoNIXcxC3xRkAibt6CqIVWso/wlvMJiDBpp1s
D2JzR4lj8MiicXkytPW9TunpaAalFf2a1N0V4AkZNKqQqRojmyXfOpZoweNz7JIS
DP0xH81l5fFGSRhEac2cu72Dnn8HtPsOyL1StVXX57TZ/KNBsSOrAynlBxWOeuVG
OVMczxUg52eTvUcQGGyhdhDab6ceYhH52KuhvLWqLaJ6GMjisPIzsOB/EJyUWzVL
FDhelxHcBwMAhnwq/I8XBhh9swu3jzaZu3/Gr+2UFMKkJsVj3uzAS0xRnib/Teyy
oGWogvVoEEh6ZwwRGbZKKdA4oHqf+8WzOa9aQ72NJQR9+U+sj8QGRAESDLCu2eQI
esK1L+7sJwLK1c1D86BL9picHbcSGV9k9me61JzEPdbZPaR0aDu8Sn2pS4vARI34
Wcr4t9YPt28KPt9syAhTRqclAhERmrGpxwn8ujlaW55LQhpqTtdem10u8MEbTuuI
pzSinIEJbikpLBca67PxD2yv3mh7jkUgar0OnwZqAK8naAJArZgqoDrqEVtgnJqx
+jKLfwBa/IJMCc35CmfAYpUErk9lz/g73cmd2eCZ8e8SxlH6iOujGT9whn5JwQi5
XXGMH2njb07kAlAaoBoKMsUymPLxB2G2kxLgX9MteDrJdUVMf60oxMZjo18z09Av
cszpHm8NNOi5tBh90mC0qw6d/XNEmNGxVpMLXgQOAsR5CzZjQc7jS7W4NQH004LU
BzS8MgLSvbTGUrBkQ25SeNhPUrQeMws78HW3USyACptrg7zxuWKYYma79O0gkVNR
tqdp6LQsEEwL+wXhnoVMxK4wqNKa95wFSgey6hh41btz+Fxlfy89B/BsUlzYA+wc
zcXTsY8U1hp1oSpV/REXLHIG+1ZBaj2I+xY8d16tw4Zvc3uaHlgf36jG0WSPxw1F
pPcHKel8ybVsvmIrPusFH5HQb9onxdp4IZaAupr1RxhQukRpj5t2eAwiM62jF+8W
0d1TNNyHlbBrEOzXAc90biMHgc/i/DAX9eDgLZ7aFBChFZ+XiaMUQelKQSs2coc5
78hJva0svOv2qsbixps+B0T2TqwNgZToYsx+5zA7IhwfnpJRGsK24e6ehINsDQWy
BZ/bPXstVvXW/vRlpCkPMLstvKoJ2QInG+7eJwalkjTFnO/apWQ0xrA6CVB7zZ2u
Hd4PAv7+3Ua59UxOsorYZ1ZJaxJninSW1i+14R9xsOl3PvNl3ejOt6KUci1ftVKa
fBWF05GNKPfuRDusqhA/t4g2ByApvZHEq3UZ47FtGOxGHFx8e4R0IIwNwGX7P9dH
9bb8dBmowhkQAerRt1KmtR3IIwVD1faIKRBWN2LzfldahTLbZWWWX1eVa0zE3S/d
1zmX7axFf6LxfRuxkJwBwRni4IF8Q2Jl8RsRB+iyguUsLOv/QzFF3H49xoEzdw9a
N8j9ehIjlGb0k81nK5TXaO2NwhpiYRBzJZ/A8u3lN4BEPLL8Y1EK9ggElYgSjAjO
mIQAKlM9H56xNNdQL6ZOg1pcsquKM06oSQk2WfaGT7yj6z5ce1XWxlol5cz6umF7
n1P7x6eusU7TZN555IL9ql3xqoukA9HWiMA/ddJdSq/ixPBB2bZu4R00BNT9SMAo
x7vmWXmy8r3VZcIYeaWaTRD5UEkew9KXqRrIGz4UGc/2zZCNF7Kw1WRn2L89Td8c
+0k621piSxpxLpk3jSYybBFp3/rndNqgrV4PrVXJugLxBTfS3rRJD9ToYsReiHgM
+tNzjRcmmlcF3fIn+qpNyqaT/NLWtjV4kYEjpXjBtejoGUcQ3PVleqhtd2h+d/QH
JXYa2xbTFYtShDnhzErDIKZiqpL5pqsQx+ZVuMuI2pBJ1ydbIhy4FE5GgDdJGEbg
0X/E+XDwgqF5TsnYJJCvZG7zP9EJw2SGBPzNbfCNqUO/n7Gy4xaxhJHA1CMgsnJh
ZW0r9VKgkLzyKA2qgpXNes4zI/ddUEVcAwq+UKa7jB62a6+By4xRczGL143/4QbX
MLWPQeZ+2fo2yJeupTRZx+HNgjU1E7W29UrSGNfMfTvxzdcihUBfs9xNbrdPVQwt
dIPEIlqsHXDjBtkSaAR8ZOSbYStBaRVj5Z10h7w029OFN3ijXCvTnQwzczIB6YoY
CmfTkx8vkolgbtmvVT+sJE/trqOLpe2GMJCvt0qtZd6vvF0hXiSoIsSI23aQJMha
uGcaGQV6mrOY/gedQMMxJdiP+LHsyrRQIUzoAb55lSQW+d3PMVzzlyXv3VzNp4VZ
VJjOI6NzAIZJJpAfuxOwtqVQtqI1NGans9nLIV9Qf53/a0PhFDTmwW9U/GXogtGo
ShZ8LMqKalbj9JL9JiuFbVwoHHAJQEMcdRnMcvJ2OGzIBF2RjRKzjdGwQklegchp
gF6Y4RZo1+3Ru+W1QTCik5qXEV7lLXbCM8UnXbHpD9vHckCAPntTTsa/iBwXGnoS
FRObDZIkW1FOg2FLe2cgDZKGfd0UKaRHX5PoTE0kYDNRE5VtL0zTypdeRUYYLqEt
CXHptAE6MztdDGnlA5gaYNZBcu1FMYH/wn1FMHEdeSkkWcty8ODwQDyFyxbPpqsk
pt3K7EMKGfM8nsV70hk50ccigFfMdPJJ6qPhPp0JqAVXj0sxrYSQ+gvzanfMdjz/
Fqoad5GrYo52dTg0QbnWY6sHIO3vXCCSzcpAwNXgKO08gMJss1arxtl1TSEv6kgJ
80pWpqg/zBsXyz995BtLdyATkz194PrIOIXtf1wBmkEQPFb3JvX94vgEUf19eSC3
JiiuwJOTWvfzRDcb00ZGUT5Kwm9Q2gmhCFFTLbSgJRZqS7xRXpVf7OXTmBQyPPVE
bFOLMOlxJUCtTJpwR0yQH8ARMEV7g9O0ZDeCMWwlJic6+4hMY0cccH/XF1GuHRwB
iKh/H0I5tQN1ZXa2uVqh/sGoHvOHn4Xut2MZwDsPcTWZlzuN5yFWnTKp8h1nGYgs
2WxYARv0w+iXXypigE7/MBrELcdaHTyXVkr1PdwG91fy+p/jfFvbfJIAxgM5wIkC
YvCf8ykOeABEcrJphx7aMN8i+2iq8fwLgznscfHLFrhG17iK9UxwFa1EGzQG4xcG
bPBkOKsmMrllAWLQ/TpEcPhKblTOiSmP8Q3Zfz6PYQvo6WgZlRkbhj8yaJfEZvNM
zUGm0wIdUkEp+JV0HNGXBeYgiiGd9EAZ0aLGYHfRlADrdKvfYX/1ur4VBwA0sZGN
ULpCOPQKF0CgeHZxyCfhMRIlBB8DylyPaWfXLX4as8uSmuG2Eanc+uyLBYGcUeyr
0WDrbYKAwxPQUtWggvDcZp7e/HRfjUc4ZdJeQYxVPzZyd955fXiB1b6eD2/GDqgl
o5XeEc8H63TBmIXvt3px1B525NkN8f/2Lb7YxCVZFzUc1q5Ef6qnLJkpjiU+RCZq
kffKf5puqXUyvJy8RaBv1jSVeEyUta49GKi8vdqFKjliNNZOVNYq4prN/OXdBXXX
UC7/jrY0RyOUa13bpojNM2BjKeMcz5r3E6Fbf/rhYmn5mOf58m0PXmtoOxh+kfi0
FXHn7tcH9XcG8vq2yuB7i8MlmPIIGDbS74e/I5qbpoT0OFp/jbEOVVG7e9zHWb6z
AB7FxZn/NRaNXETxUcoNB+MS7WGL7vku2pEgubRbrNd07a/t+QLQlojgi+DyHf81
0NTRO1ga9yEquywAtpqp+hITozjoapwUd9dHNo6H5LphfWoReQD+Brxmm5cWLonQ
tLpl6fFPuSvdyJKxg5BeuVcQl8NjtG6WWcHb7xWsU3V/0r/FZdDTbtP+ATc2npqZ
CXz191hNzQNK8fcOJWxzb6jGN4S3JZZ41FjcCNZHvZCx07SWb+IrJpUMnFG4e3az
OB8esl0whSu7oSC2R/vdxAYns0sVH9yV7pJxM8ck0gPEK7if8DbUHSBnUlSLkufd
bhJlAzposQTeJJ6E3Zyc9nr86a+xmZGe+Hq5gr9x1KAhrc2r3ehmO+kkJX0dnxvU
0uoruU/bJbSGtHAv6RKYTz7vs/AHNIXFkpJEV1mV2+8mIct6MYtyU/TZx7tsdjMF
F4pLJjqPqT8g2LjLFBFyysPiuC94yHfbdGh41T4vTm7asGpYX+JPgOFPuQ+zFl4D
HVFbemSvFqkn9bh1fu3iRP0dVF8zs0H8BhajCzC5otessmvmt8+rkCWjzHDHuKe1
7Y7NoCPEWYaPa6JKNHW4XR1ii8Qogu4MFaSKw9fXcbJOPJ9OP2TbcuZWrwTT1Gxh
asX3+jsR5KRVn7uQ6i8KhMEvKZHcks6t0QmKYntrOkWmbScO8LwjeTCrisX9IcHI
lR3NDvZ6/M/TVV+ZgCW2MJNJ3GDgUgXpTh0z7zwlU5t12wa2WR5K4Wtm7d8rDnkS
6tYkU8H8OpLeY03XNc0fcclwGfTxSiY98l6cHSMZRP31nKnS3Tn2g3n18YrLdXyd
gdmr+3PmefosDcPO7qtIeaJ63HC1Q/o7VMqtAvqK5gUiX8RUxnnHlEzQp9sp7y+C
8TGrD0+VPhnedwh9086hGbRnjAPMLIYEyR1G/wNQ+q99Atq1oy46Tl1GlFvYPIwa
erMRRcXjGa9BqQqOqu4V3RQJhBRe6ZqZtHyvTpQeuKh3W8wqMFt1F4hHPuVpAHdb
NM9XkyKDp6Pw+i47hS/TvibUB/2ICqN/6xFecKmNALdV+nxnHoYEsIPId9fItYa9
b7F6U6IQVoBPHQdgqGJEtCJZO3ENpcjwNy064VOYeSvWlpltT+LyJiGU4juzcM5w
uRhHfoX82bfnFaFNQNvMHebV77dsCqDd0ymLqCNySPoLIrmp+gygKRtxL+jTGiE5
7dHanKwpxk1uMiVy56Q5cr28jdPTQL0bvA2AUc+uM5f+pQ+xEu4yvdb8flo+vT73
JCLW4Vd7zMHuLkAzERG0LhFnXR08tByPTylm6D+TtAH4fASIo9uF4Pq2szOU/WFU
ZuGsXEdl1Zxn8yLyiFPI8ismZV6U6vUUKga/W85Gd2lIYKTnktT4Ilyf1Eewev3a
0c/VOxa5S5Z916P7I/TZWWmIP6NrwSWwfZMOtjdVB6oBnpBJxWulWlPlikWDayEc
1mMhOUw/mn1PUJ0eEIMGycDWSSf0tIelpe8IMlRaSpho/6+zMexKtvm7/Zxw489L
fXskTnbjhcXxFtoOEw/jiDUHMPbRovTOoLHzi6olbJ+W+UeX+o/UmzrckjYIAi8h
Rz0bJ8aa2fgbfyppO2cdgYExtWixZ5Zpq/vZp8dE/I8rUykiC82SUFxWkMqWqcPt
aOjQ1c9pLGdKoIkcOeknICfH4bSwkkfAoRu070Dvqz0Hz25tUtaVAFVmRP+ddieJ
JVdSD5asjirmdl/y4P26zg6dZYBnFHMf6RavC8HV8gTRRu+l0GabURnUaBSnfdk3
2ot3A1AcOxcJW/wcMgKXg0dR7R/YYD33qzosQrq+LEFQ3y7zCDW08dK9MQkCpMyI
QewzjYLk3rA5rWLMyuJonUV1RnieOK0GMCpjDdjzaxlhxWpSJEzR13daRylgCz7q
gdUYVb8h0RK2hCQe0C4UTSLTDIFc57ReyZ5EY/vgnsgJgUS3tqbqEdmJ2EUMfHXz
d0drK97S0hqeFcYW4vRbrbP33CqjvnceSb2dyTSj3B7o1zKFVN/PVJIvTnsa5T+Q
6wdp4Y5Pacl0i7YlxtOFT5mDdVtFx90rRYLGHfxCxfgSH8a4rVF8269OhWPTRPH+
M6fsiYqi5F4bkoFjA+TuiggazY6r8WCnoPSwYpCKy60u22NbZCMxmXQS7vLd7KnI
K/56qFVGJVs4ho+gX80bUat5nmtl8g1hlIiQLl9w2iEcEWrmsIV7GEQjkKbzzJui
NgchrSGL2P9OGQAFcIKE6CYz1+jrkBmUEKdpIltbmtO+TVf/260mxIVCu14rhKcY
japKLHLgaQqpeb+P4Qv4k09b/ukVJ6b+efOelqZfOmx6rj/XtcTTyB8gUZyoDOHr
XrI41LGoW0+AOiA8ao2So8kC9un0ebim4Cbmhg3rK44BDKetqzETW71zg5GzKb33
2zxvS1YpmstREDl32ivuMZ36dq3Q6O4HI3DT/iXgYwzWJ7ti5V8TUptwMT4AecwT
MzzHAvxW/PXTAPU6Z1ySwcBdbPVUM5F7trczNzdjle+0d417lxJ8N5BK8/AG+nYY
XGLC8tHtQ7sRYMSRqBzv+RYTSyU1x/OldXLk49pl9Dsv4IADE4R2/hjKAmTxo4GA
JAJSi+POa3MHHaifruVvu4WeqG4rmATAxm6HNs+n1LZOoqE/McRX2wo2zVBWUItL
edN11cclK6IZobTl1kkhLJ7AmPdXpu6UrRWaUDlyO1Pghw2N20Wt/JjAfJjt67ai
8wqzrYlLamuJ35O07tih/fif9vAH3UsxBvpAxvpErYlr68mmmf93V6/uZiUX3pMU
wpQAljr/OYvkkNqtzN74/U7rlRBauk/d3t9Bv/Yv9IwcEp9TL/A7I5t/PJvdoEk+
GLnenj80zIXXcZXYqG0vI2qVdxzb/jwe/wuKI8NyqWlcAzC4DUnXje7OQoFROjF+
4wAt4JMtrnbbRu6sgNbqYbq6gDJW6jWl2J43y9tE9Yxk1xHxHof6BgN/VjUgLN48
z2xBsMOZh6dyZm3k83jTSLNTdjKl/FVsVkRRGWsirNOmcjTB6Z+fWNTPgDlUhxpt
Br7UayCfJoV11xcNzjpo8dsp7I5y+zPXVwgrMv+acmSomRD1VzDWmRIPBVe1Hs8q
mWbBeB4u4Zc+1dF7fJM4427DRU+WclIxwZYyR4ou2wcJeFxBCNgHa9sOTcTG9TnE
XLJ0RjXVe8uDEZ6N4fDeZS7WNkND6dyHNe1mwi7mkz71QQ6rFfu/yRZpu0LCz/xJ
lXYGAn2C/RAwUaySSixOWva2nhXrcNyxOhY8l+xCYF9k/i5+rc88G+KtnIOSvgdp
eTxz0eKT4Mnye7QSEQ4Tif0lnXYHf+i5cF/C04PG8zVDubnWEhrMyjjXGjxtqkz3
e2tmXIQ5VDbAO055t0uxtcMm/GK8XHgR2++XNuXTQWG7zfzwcpCAp8TZhfVdQqVc
jFHbzyyg4M3kB5gULtH91k54kFq/bRRw4OhxrwRfci8mFMZT4Dj0xmzPJstvckFK
wrZl3HM33mfWOkXofLJV5T2sngxMaGJZfam1FoHa8aBrtsy6h8lh5Ec7rvLeO87j
GyZmSr4lDl6HrxMGzTc2ZnDCeD72GoBZfxBOJ0taX12qWy2Y8zG7DfxXgmq7q05t
I/x84rCvmiUbGdTZEOr//fDvvURaeKJQZJTNbxZaMcaqKTCDrCOhgH+Igpas+Str
BrhZ7B6tOGhvpbyWiT3flK2Fhesa38ToggDKx9No7ettyZXsaQBjjEqHwl0ARvL6
H6/4evR/VE/ZEt8guFk3n+NhF+C5eMluUacN/4UsDfNSc6axUGSgw351W1qqmOJq
SWbZMLprAwkVNcdHRRN3Tdlc2g5Rcer6s3fqGTxIaDvwxqPmiCosIAIshi/9D2r5
nwjbrmXUKRGk8HQeyeJE7oHRKjgLT+S34etQPwkHTD1ES97BD7R2dzQfLCSIYZSK
l9mm9aEg+RrWxMj1a/rViUiPGhCiCQjg+ZBsnB5pF3NQqL2KEPbmCyBNp4OiQ4Iv
rIbDMAFEWOsRtHxN4mpSQwdLK+v/d0shK/8Qy8p+ooAt3FKW9b1zorApiMZlGVp8
eMbcFzVi/YKkzAGXxY9CX2O4kE6yPxYl0xTd5WEUiO6D1TEWoOHEEEa7wRjVnykS
MOrDbzVI2Xwx+G8vkj+iBiqpRIA87uOn8ZJ/OZgPjEa54WxRkYmMZCUwgC80fQDK
lrXU9hTteEAhJzadzvdk31xoyanL9d5k7GrZQNGDuNOUw5+M75EJZeZfiA24CCzG
QSAltHGrJVMIsx+AO5Sz8pPzx0Z2PRZHJmmunzDDZgilhrYd9Y7ePJUKwpoM+tq4
gUC5R3aqEreeIqyM/1mBlvsr5+V5va3oiiaXrTsJcnQecI7R/MTOAjz4Awiu+FRL
CYzVVeoYMFwO/kGRJlFO+vByyJvb2FDHJbQX4D0EIBf/FGlgvgRqRZA7jGbdXO+2
jWCCf/UPJ5QKzdJsk++648927EiBB6vcHh843K7i1ecGFoKTDDC8rQ5a0648lsdD
1bDTdjINS79PcXStvIhFVuO20OpvPQzqhQOfWLSIQUUSROBYhnoJWB1yuKvRTeHp
HqcgrPsPa+7dBm9xem5AXibf3UgTiHmjG/Z5EQborgLisOv4elTCw/2i+nxsmJFR
p6Jdt7Fa6sigksoxqZHCRwlBttBxgURiMBjJAixPKAf5xqtm5/3rd19Pxa1T6nrr
DjU8vhvN6INWrREl5+gxF0sF7JMYLfEUbZA7OzVMa3xgjL2axkh9nr036w+ywUOe
DjLAWinaZB9/VDGBUxH+0VRsRXJkCzNCQvAeIvhsBiR1+C8/KBBGFOj363ea0PLv
eXmGT0kU+FPwSHdL76MKq1H5yCIekASqJWeSxIh3tL3P/01vHM8OJJRW27IHGDdQ
ZePqX8v33XVjYh6dQM2bm/BfWLSAKyBgcOFk5KF188x4UyQuptHkVjGBDNcklPcD
gmRzx9eayIWd7ODNzphG68RIC+OqM59m+G8Q/xOJHHaubdmGLS4bKb5lw9fTjYT8
TD5LSvgd+C0YRFFAd0lN8KKmA7VE5djqtmQmYU63BjFG1cwSqLwMQa5gtPMe+uqk
4Ttl/N3fI38vTC2aZSUP2pOKe82rstOWuOqMkE3S94F798UY+SXQ65fIxaFLdKZl
WQ3CnAaV3sqyhMvAx8afOnN4NI5Hq8SqINcBjAtT9qrFRikukZhaEPZznHi4fRCK
bLQ7UbwzlOniAcgVEqRSPGChPOnIQgfJQbzXlXqILlAJi946xPjvXY+Bmkdt4mnB
Vq0Nz23secc6N8EruXNyc/g+F3OXwkzMAez95+wRfo5SwbI74UHBTfLb71XWe90V
22Hx3+csuMcyInIx/az6xIJCS1W/U/6hQ3ArD1xqpJOXJ6ZOKMFR6tXSdx7QmgCi
IpfGOWnCRuWzshdWDrNu/9iwS7yGTp6tW9Y84Iq5M4deC0eKZdRDSjdKCJx0fUwv
NgrBwFAAACLaJBguV1BdBGGg3YtF1/APB27orYp36fc+dh1Lh6gdfiD5GAF8itUy
nPM6zfgr0vgPKQhZ2qP0VY+uhEYcU2CnuuXQPAiE9Xwu/ky4dTgrFe/bPRtnccv0
w8ZxqtQ6SwcVVER41Ae1Y4S+8oqDcr4DxwQ8V9z68x56smqm0EdmSG+2QBU/4LLj
mSNyRrQmhfPJNkm2GMEkJGXqEbzrHPW7986mugvVaraI3FcXZd6LkMHlNWsmQHz6
c09lTgRZT8Ow9jk9hCNzWNdYxwayCEjDFXshoEMk22pyf4tGDOp15OsSslHRrBtD
1JFAUBQW1pfnxhO54xCizvH5AawIH7GEIeYQ0dJNbnq2EG8PGzEz3pYQnx6KgtUZ
CqihykXmldeRMKX+q0BGMmVS6E/rB6V2nbhQ8N2awwJZUysLVUtAhfcpL7x3Mm0v
8KSw+rdXaYut9nBN1Yj7XptQB8OA7INAghjXYE4AMsWxaReiIVlvDZgY0mSfmHeg
fIb/BKYxdF5appPkhumgHHndcpDyDWAYDEB9zQA1Zchh68gBGqj4Enm/T9ZXXWAh
QhNq3Xlu6ck11zzDHYiR58atT2V9O0T+u7Ib+welsZSXQl9PhV+w4rJaabcfS51+
LTaS0K8NfEtMDmB2KWxwQmefdfX435QmLoTe5wrQ/bpmdo7R8C/dyeJ9LO04ZpFY
GTawHTpunl+4dalHhMfKo4HRbOkvh3pbNjaqqXSZJYeIWeuvsV20xWlTWtOY9PRf
BoBlZpFqCjeQzkY6CLiciHLRFjjciCjkoxCBlTbj2CshD0wwKDRGaJdOGTdqkIMv
gAZSS3ohcE3fljwpG3ysp1wp4Ry4Ujm77WIQ2VDP3OYCuXScGjZ/fPa42CI7Cx5/
IxMiQuACgM6IN6bxooi4SiEw5EU41DOKvJ5eMrEKgpt3mMOEBPvxF1nFjH/HdiPs
jaye+f367wEFC+8HbcWUkkdamJvFWDDgMp5t1NmqsclxE9MnNlTU1AUSRzksgVn7
fF4IIj1mFnO4nocWf6bxNzkBMXldnwoyS061hPMU65KzbcFy4s4qWxK07It7FcUY
wIZzvAhhlv9bHSSdn1pdL9sclYxe4NaLkAt7him0fLmaFeO5Q8OkUahEzuRWYqCd
g0PokJwWs5VoH8B8O5CQqZAhVsTvSQ0hnhTTOHWzjsL+Jk8pj7FBGvEv5ZIEN2db
wjRfyl8t2NoaSNlJbzaVnMX/eBQbNhG2Kt+COyf6C6qio6VZwzaHTVsjDSJmbg2N
NzGtzcEStA8qLQF8BnT/L4DMjmCpN+fUA171/UX0KfE0+5noG8rLahZG4dLPfsPB
Zt4Lsm9B8qo/Nj8uTN+0sD0ALzGT+QlqqWC8Ns26ZOESipkFG4WDpqGprbxGi7ng
7h524WGSLi6rXyoBoi341HT4egwS6342cWJKqkkD5DAwCXwLD0/jdA2J+9jZu/H9
ehXslPoXJsAFyc+n/EUuTPBCLhSV0wHZUPN++n1A6DYd8/hG/DoxbgqPleXCebOT
jHTLB78yZ8Gllq5reCcFv0Ibh5kuMM7bSdAzm8YoG77KZqw0kkKJVX6WIIy/2z2W
jI2Fed/nurj9tF9jQ9lpVi4UDFXJ3RJWVKkcx2/BVJvMsFI1C0EopewyWCR9Y3C0
VkkN2hOZze2rvwv3cbxj1XrVgKrsLV6br02Yv5EnFx5d7tyRVbS4DKpffc8hiqcG
JRk6NJ0VcGLLLpGfX9jusMG9mBrnRMpZUX4jNiUunlmKWEuFx+8RoYHyUc+muhNN
na3xO+bAVCOv3rzw7/1jCSH9gRfl98xvCFcQmE//BHaBEyf0f/bVWIZbMOkM289H
L2dwix0ahCJuW3npnVxV0u9m5ZVfqtEsxf0uunJmAFo13cXVKfsJ1WXYNrLlQiho
uxCCiotnRdo7/7CfpF3y3hWZfXjmcX6OUdfRmnKDEC9JyOTwZYm2s+79pCP8F+G9
WQrB/RMOz9SJk8ffyVaZpEJF9zYMroxtw5J7MeR+A/fg3HiO40RDgLLUgbaDWwP5
HETzkZMhhPqB/GthGw5ksKTRxLHcY+9f13plgnIPzU6HqTIhpi66La71+TbujqoB
6l6zeBo0S+nEyCjzcm2AKZMRiRkIa4OEAZqhbdL1Ikc7Lb9X9uKq3FuiPDY3xcA6
mzWIKCK79btdJ934n58beCAlnswBOZaLsYcSMo53Mpu0ixAiItNtmpdeuEho9TSd
D0A33Sy9qVZns87zqU765bi3Xy8abGhKDKsaKu/qprd0463ch3EopzPoEEp82KRk
tD3Cf1Vdbh8832ovDPOUrOdesD//Ud4xGJEjheBUlIUq2SHItReLRE01DYaxB8uA
txoAVu+8CEpnX/eGiq8QSAnrzM3M3QXCrR1c5/o936DwGFum92yZbmiafpN8Jlr+
9XdP+Z8K1zeSbsitOj3HmK76vCaJV0pKsreP3YrbpOBVUcbY/sBv+sER8d3/ogwg
d1EgHcDlHxvqRZnBpSPufiAOl4q5cEglqSrTH4dwXWQKW+Zak5hnU4KhFQQz/yaN
GLvBh5xNBBLOdmw/fWoq8RowQTqCvxBTUl5tqpuuzY8Bqcjnzr7eB4ikSlBvExLm
lDiaAV23jnCxGZhHXL6mNuGmLBX6VIyjy+Z3S1bhA/K7FibYfaa/02vJqb2zt3I7
Gi0+SIhUJDduQydi5c+/JKcXkfg3aoFUGo9CJyNVULM4XGQFDj/UC93ZJvkH/7Ue
CE5eZLWTdZnTMOd1l0UbmF7eQG4s4z/ew5a8381/X10Pt0HBUx80szVFJjPy0CJA
WeUtcVqzqkza5PhOnboIQ9DH/dboXGPvFV7EeJfaaMIqMY0/7wQ9oXPgvglJNcy2
P/v9Rt0nfJRh0IqOP3wWL3kkEiD8fMA03iZGeJozX+EnlcZLCyUz6rMF2li4pzJf
AZiBgamQ6GgN+zceBpxaIKeYLuk4JcvLT6FEk4ByRyjdu/bRYcquTS9ZGfQE+hJ2
BOv76ZfB9Ywl2vJQhiI4EPJD67VyXcsKOJBUleCeAXZYuy7QL0L8PFi8E2ic8J3y
AGKgfKcAf/y566X7JMNYTNyhcO4avyO7ievbgMtZTCQ/PRJcisQQKtqp5jspIB7s
cB/nGiOYKaMw/sypznbpkJ9B01JechOcXHdAgANtqAf273tqgx0TKnpdSfPH8AkF
Joq8bLm2b31dV0mJdenrziOZ+G+b82UO8asPPZDtC66eEc7Wa8GIqT7OB2jEYXiV
6jHRMcJ+qKK5LXstUkgNxnLUMOvL6Jf0FWKkEco00MO7IS19SZPcsOcWqcWqImyv
RR5bVGO1YIaGeFQvEG0k2eUxxlgD62GEeNHgmk1wT22zMxkUPBueldewI5zJEqPS
YO9lzyqMXD2owwLjvZ4USsv1k4X5DwlBU1kMSDiKKbljwLxej9Du18NCZpu4cQ7O
v2ZR7JE3Kdyqe/XuD6OhhYJ82gkx6Qph14MF9sfrTJFqe3Ry9HmlTIKHDehZqXF4
d0crLp9gZKyOfmvDovfrarPncSdbsq75dgMh1vXMDBfMqslbEm8yqTFXzd6uInYK
sCKWd7KSt8fclmc2fhMNp1JaiLPBCDLkiRVAYGUghHtxzC7ZZqh0pgdP218ap/3q
O8MqeRntEHmS8o25dp/1y4GqiREYMXNHDS4CEMr/UpPa4Z0YSoSNUyBGL3s2gVAE
hffRJeMrcMHKuAf134j+2VgrpS5nYWLdOBzlgOBL2GbhFEHr6vUWdxWC0+yWInjQ
visU9lLgGBxEsXdTyJYoIdbxBHXniLp7PLVDFzDJOjsyh0caYGN+m5SsGmcBmqB7
x2+CN/t274bre8ubedPzK+naIgjVtLguDQ+aSFkHHe3v6geh6FRvetxE1wLJKxuF
Ol5jdskjqHOQs3hWjswa7RuM3BEfEcLAbKKT/HPx79TkFFknTr3yORGgxj6ev69o
pp2MzhrNndwL31gr8o+XPZej2i98tYDxdf/YS10abBkvrwhmJxqAtRDiTnk1g8ZK
jY6PGhIpSD7OFQLpf0SJwZ8W7hlNMXvUrWtsgO+vMh450TB009Dyk3mTuAIhL6hg
vxqn0VYANIsLeWxZ6wmXuwhaf7nQfytS694LtpPc7rAznFsi93dT19hH48So0vRn
fitkQ5TyMjj1SRkYOUnM0l/wV+dQRHOhtawoAW+o/4hdMRAd6lSqDYdjVHskCo1a
thvPx0Qx7mE2PcQ/6mMXSKaura6eYswhcWTdDsJxUWhZfNhK1f+JVmHQW3yOtuRW
CalgdJd1Aelf4rwGr9zxjnOYL9reZPAt+P9wfX2dpCbQJvkMBvLVeGYNrdeM4mlz
LZ5XtceLKIweaVX1LFgHky/n1d/EihEIRg/YQS5KS9Fa7FTz2jwNwcywBxdLoox/
802tMdi+9cVGV8p9+ElKD2Mny0iZ2c75lHwqTZWmeTJRbLQClNOUEuPOufxW7G/z
KE7d1oTsEnigQBKm6gP+GvdlHcDF9WP90AxzJbGnKXwy9YiXEKV7uMJW2dOwBueS
Z9zkmBf9Y2DMl15sW8prXGtorV8zCirDPZYgexXvzWFGA4e/8styyc/UdGrEViXW
aXbpDSP44rTnqTA310EQ0WOVac9bRgLIIiQG7gfhsYyHZcYTVGPRmSheJRDfpO4w
1Gm9neIjvfjJaZmIrBluNngqHxuxoKndsbFZKG0iwMS5+3B2crH3MWWZNSBej9XY
rAEFHUALA09FldNgpdvTzOIB1RCvanRb2KbWLbQiXqgcPM85F5w7jMtxeY62cfUz
OljgB/65nMiyQrkIaVKJbWGyjidnuOcuL/GkfVH1J8SP++yMu2baMd7q6yAAdmeT
oP3INFCONcNoaRoCM0//t0a04faw1k0NUdlpL8V/Gk1Udi2T6DZa9UWRCqT1TgoV
OZ3dMiLIlhpnnv/ns7yOdfZAWjqBgrumxxbodQHz2TTMhVZEhyy9kGwNk1mniZKe
5Y+7F99qR+prGBawXYQlKH3ArjzG6rwtmKnlnESb5zxXrQElTl7P8ZlwpKDVLosr
aFZWWryaQZqftQ1wjUy5+pwB1OsoXkSX+H4DDoXK2O020HSfTJRziLOzD46FWMm9
EZ9XOF4nhI+7ugn5kY6dnHVDwXzoQjsGad/xmGfQFHFrR/lch9QLAlgpPW0lkHfp
oa+WOlAl5xKS3Ym1DP38a09o2jjUv4tU3y/uq876g20hoM4vfQ9ptS8WqF9MVSnP
bpgn9ZBZrlzfTKItJGOmZIECUx6ESzidgeHrqQFYwZLjMtvSXdYZN1+q/C/HSTWE
HTXnEZl7mcvO/+22YhDOiWz+ETblASDFe2ZXWtHnSAb53UH+fPK9wQlE9ozamABm
LUnZJfzuC4oZr19TlMZEiMS0MfEDlYpKQqvKZO0lgr96CKWv+t+Gm5yv+s4lqivJ
lBNSkp0HENTW8TtFbEaqr9or3i0Dj2cXhFN+RRgmD2+7xx5UjULpLgr+yAO1OZ7H
S4K6HG7p5CpV6YZNTpTIj2/Gv4HBlguV+HLsOucMap67kV7z/ivjUnyrioSVd3qZ
AhocZMX4NoJyJMSoFDrL0cbopQlthzpqb1z+8VdomkqHFY7r8Hh5NZmJ5VoxTnzd
EPLEvkZp/RMZ2r4wOiD1jYry7rU8OZW/bsvESE93hMiQyFIzyBdb8m3au25aiyTN
lGmxqUFln5PdBSl7yDzPSIkO6SulTCVsUWU957Lx2iV98FJYYmLECthUykAJezMX
RkXtZeGKlAANW/bTQ92HWVr3BkCkr0rmXawFHYdSooutF5hmKZCmWbScruJxWXah
2Q1moCM/qrD60EOdDjqGNLOpJwo8wdyj4FrZ+ttx0WO4QS039yBWXaAWYCHA7iJD
MYGf5lPOstol7+4ZEiKGi3AMzdRhjgxat5Nve9dkuFmaccTYqItr9F7bvjjYZ4aR
WmAhJubPFCmDApjvWAGozKjfakscYczHYn5YsMay4KHbd4eSy1DlutDx6/VwEbyn
zNBcUBXZ+yUt8PMIDkZeMIh+8KGQFLkWy02yHof1O8FuMwO6rP8lD2d0/xgCstq/
72O8u9HQXAjE92mwKdBUMZqFTPqblMlHzgcOAY+hkx0OXp8RfnsgW37JDeGR0gwt
UVTup9U5cvoA+RNOrmWTkG/PnuXsGDKnFGonfjLzZIod417dY4H6KB7RpxrCQbDt
aqnTe8JfYDEJIJV1wHHKZGQvsVQGPEkA81YhAgJm8MR/iND00JcIoGl+lr0RNnLP
mKDM+vaoxm3phmLE41FENR1MpmaB3j0rwti3Myj3BCLdp9NcRsRU8axHABWyeHiX
7v9sI/55mm1j43NFkzL2f8EubRMUpD973Q4wFJ+bHXgkgKqnZWm6xb42P25Op8Rl
e+OIpnrvCXPjwiaTMJVmD9+u0w3Af2wj8UrbP7QswDHF6buchuKOhax7vYH/AYrc
DWwkOAyudEBlX7CPeiwxbZmGfBmpP3JoFaUBAuvYPxkiRng7SO5Kk2rg6Vo9nY17
Mu4C33vzg4TstgkW/xdZgQz+Df7zw7sxp0JNIwb6Yp5VNa3oggCCJIXjvXBXgAry
u9nBrZiKowZVALyothOaog7syZ4kPiDoPxV2pwsxr/SbWOu1YIwSI0HyR9Rs/Rip
mbL5QcaDKh45ZsWulpK9Caj2FMjgNfmFRdbUlYIYK/Q5WmpzBU8YK36cNfxkXJzz
m2Z5NiAE8aRy367bNYtQNaaaOCsULvcpZ0DM1VcOCb7fKRyswe4tT6C7mTxGZhbO
9kRPyi6IDrM4uPpJ8GMcHVsTISW2Hap9TmzQ1GJLEbKvpV4+2DCInn/98rTkCiZt
J8qnlU7PA4ZDNzZDTqhEoqNhQblmn4WJUcfjENyET1Vym1TqjCBONbWmOdgmrch+
XEmkRDLFPgd0qKWUC++z/YuInwnZ6x6UQAk+RXILz+2j+9Y5lOJl070KA2KivHqf
A2OPCeMbmUcrSHBNRwDfuyUuvyvCsanOFdB0GLJz+zbMCEVOVMesOkAYLRqQiVis
ZyxAUW/2a/l9V+MfR0hzdBCXZKIZehIbIRZMeSUvkQZIp8cEyvupIi6Q6KEYeQu7
qbPhH1ykM3MMBGLRkuci/Dz5W5MP+HowoBmGPwdFFCYefvDmViYyFOIwvZpqm6v3
S16BPDFdWRb0b5JSH96ZHQX5UMKd9LvG4qyMJWSINtKPuZ8uW5xwMk1SltnoKOag
Ugxh1b3wTx4v+J3XFuk8+CdSWSlFedrDW4dfOrkoBhYXG1OCBQsg+btcRqZBPBQT
2yliSbJcm8E49NQA8KvSKJT80323N3pibGAn/Z1Xw1UP/tSNjtGc5cC+6/UczYsH
ei3rcdqyK2V/pQWkuMw6tWmEYJyHZ3Dce3AId8bJovICzeQK93atI6d7YIfQw/qJ
G/jrkAf8+N5uvU26evaBQmlKOa3t6d8D03T5pEOtVeGK8jXJMKrVid4eAyamAuct
2PofxYtSmzwLINQJoAjnTNQZxXhbwTsQajZ9XX6MoWt6f05xUmo2Uq8J9qKXbeTN
ORgkxJMUVgNgnaju5YCPgdr6mdXNfAx9eyanj2ZgLoBRBgeYmqfGn+2q2u5847g/
HhpbEyPjiOk7t6VGw0C00qktVwHp+lf+6ZS0ICLZ3k8JnkAiKrJhutK+Qc3RkU0g
YOmTpVu4qSPOwduWzxhZiOlDykhhDCz+pmeLAtRYE6YZBc+NzZana8HwI+sZDyIW
vdwsnaoNEAdJB0hQoivZB9eCwZXWXfeQwZ+x7/qZZOpNP4QvvypF2TPnjxGh6Myi
ZOnRWRRCjTJ9iVI/Adz5tdx4W89+u6CPlIAMKui/q7+2jCY2QBiG1tQHVSrO8tfb
bRKTzguICvAd+g/jBHPsJrMGXWcyVPT3Rq9Vpo7zLJLzZ54Wb3la06lhFc9UxvDb
jABex+gDFsWWCLvxALmtIdvWAz0llIH5lYeIVAeZ0Ug1225Tk5GZkJmPusKENChp
/XPAFrilnaqQKG00oB5P6l0tf4h7s0N0TSSZ7pf1btJevqEQrAnW1t26gWe3d7au
tbd80A+P/G0iOKPD/HyXeFrYPy1BEe0aF15QvqXMaKzn5N8j1EvQS+tMAy4dm5QR
5xjcBIrhGdP6fIdKHejBLD7M5SAdHLSQF2iZPXdMc+qWmrTJA8yblKdEl+HNap8F
n5SgvhGSgesgffq2dbPsxcjtEHVb+rCcGV66eMjg9S9+vwH8Ugz1CDtWkl3yKfsy
RucyM0cAr4QeY0JJvHJb+W7PA/jB585UYUDZK6Aj39wX3QILpAkehDY9OHlTBMuA
PpXr4YNsn6zZcwGgDyqKgl7cv72C+yzIaynD1eIDzeMG9Zk1r/uZQzbsZTkMfp0F
iucmO/ldm1zLoHHUj/I+djBjEWnKuGkd4BYjO89TdueHxT9h3y+VBudKedf2HLx5
23hYP8L6yDZw7A1MAKp1hZulsF/+73pm4l6XF7OEOc5CGlKDvop0PmcttWdMbo7i
7BgKhgiuXgrtkIGSAmgAuguQSBLXW3K/0vnaD49+5JrHIp8cvILDrBqtQlGxJVBp
vV9NjIiL31kQUQQhVQHI3SQ3GXLMNN5OLry6l0zwAW21XK6w+lGDDz5PYliNhmJU
q1i328hvolQiz1kJ7yyEdFNI74bxl0cmq7tA59mV70S3HcYF583NacQ0VC3TOy5S
ggsAyGj8qfaDKi0a+5GA3JmzGOy+z5Drcv8shUzSjjL0a/avYzUhm8pf0tVc2UXq
khpk7w9Nc+yqEKnXEVJIcAK5YkHozdQZ/PCVyyOcvvlfKCpi8HG2A4c/K4hO2kyk
0SzCjDOBIrsq86ap0zcr2ZIS7FQEKjdNA2wgH49/d2eiiyBGzkyDLUCobCvgecEv
zRhEGsF5wmcU5mvppg/2zQy7zNfmHRzxfn84IqLMWRS/werXEwnqUwzBL1NVSwg2
xfweSt8YGVxudAOmS9+5LgaIihsZMYWWeWEL8tApt5rjTY3j4P9ojc0RCbJOs/21
xtlcAR1l4CEGAsHhDlB4KJq/m6mirAgUR1+R9ieN8RpQ1a/8NmoWp0ePJGJLWG0K
pNqFksmySFfUFiV8ab3HuoIVMinnDjP0AcsITGJBbZgMpfthJGUYLrWyOfHxSDB4
nwk1rejpfXvUs+UMXtFf6xUA9KMhexzxDXIOCB6lSrk2QWMytjQevilr+mCYGBlk
/hcv159X5GO7JW+Oz1J1O26ICJpMRSW6oWJSVILjTfcwpYHYN6ptDbMvFFJ0drbZ
8QdfMz/V7yLeSQZrJRrVts1CRckwnlNetjXNgS2XrBkzbFAQMbV4FsO+uX9pfUd2
m8ZRB7qNfETTaWF2kgTe7e6jnWZUJ15k0yXqHRBDwlSbI2Inh8aGt2aHccjIHpND
7DKU8ZKUn1PyJeY3ZEvSosQJ/aWjpypc3+d3VPP0iGZozaR1or57pbW3Swl08+FI
e3/4/P/NTHMTvhGMRdQhSAhipP3EyQBA56VQ78XawRdRLXAqGT3pN6b/cFmBoz7s
6kSc1UMr0Dfw6LxRdaEVL4UTGOjvuhdbQCSmZCzC1p6DO5qTknhDgy6nf7vV8ubk
PEdiUV6Tr9uFhH6evZu8onqYhLXmqN6GiyuZEYb+t7P6u4q682h0p26pruQHIvfA
pmAkz6gTv4Gj+YBKPVCZWc3uQeKGRwPvxYgeIcugJsQJPWjuVFRQ5D8XcULHgZu2
zzCvhnz3NcdyzPwPkTJ7pLPZL/oqiXVCquc0WdEwPC67BjOcM+WPBv5c99dXf9pD
w28SrFOwnLx6IClM3zSbaJOcvEjVk/IkQ6D9SVAoGijjphHLTsb+R3+WVEOt8bUl
O7+5/p5F8IbQiC4ZV39jd6Koje3fZO6NlnMkHft4ERyFyNI5PAqD28KdG2hvyFjW
aEmppsfzYDnbdZBcZE3/CxHXnHAXjY+NJyeaf9MRd27HgIWP2VpKZZmYCV0J/U9E
yOcb486/tO0LWyg3b4yt7/6eWlGzlwegP6/qfzle+vyMfGnKUfD4iBsWVDa2zjyU
Sd4oM2JLzmG0bDWVTxSwcFQ+NHuan/l7KcJAijkxX+8OsFsNCiTsvmDObCAJ9pqX
w6Gv9ppXofdDdBrguevMch1SSWwWpFnpcNP44P89yfITID1amsDQ7TjSaOLaALYs
owJcTPUU6LrTSeCXtPiCvEqfdnZRUpYSdNSj0vTgipt0Z4qYXwz5WiRXfpRj+NcL
6WEEAJbYEUTyQTlev/mmBLtYv9xPGOwElkiJPXjSG+qhTG4bDEKjVv/itmaY9te/
ON4NSP/FipKIYpCm27eOGpjCqQGmQWqWODHv3DdJ2/2EviTVIwRU9CMxgdDJ2/eb
JzEXtxb/z/w4R9zF49lOdcJNNpDl7JH0fCUP1DZYRpZyV7f3cv9hr7Kkx/ZfT6jU
PL1HhmFMkgxneo3YFEv18Rj6yLnV3C3q7Q2htP/mwxNmMJLOjLVHXoIj2GDzRcn4
7VKBiULvIy43fPa4PcU3+gdWfP6xhdgJK5CMY4ga8uh8H14S1rY2RLMF3PqpzvJJ
lsbz8O6awr/xp5cLuKXIf7V3POFnOEzDCfRNqJEHL2xkY6IS5kq+2HMqIjPp4p1G
858OI/PfcKYlK9LEGpZEH5Y9FqtAjE1cSf9/x0JPVfY3ANticIbf26zbhujoxagL
msl/Qqk4zmr7J4IDr+w9yGMaWQnfnXLAeeyrpygYdijmen+J5f5uuwOy5l6unByY
kdB33ut/pSCrBQmiVA7Ap8ghsg5CwfaMFwKeQaXu/ZtOKQcQDjADO3KnpjXc2u4b
GJGRHqADJWR48n7z07pUkHlg+29EPFRd708kco6ZIYFNfntxNfx+kRP1uU2G2Vgf
Qr5xs3Q5itHqKoPIAKcxop+MVhv9F1AWBej/p9ESbhcaikPYYY1ZrfXflUlLK/W4
p0PTGtKXC9/34PvBLg8V5YL5UXwSD3WejV95JBRTKSKyOQpiKxCVtnonVA5lNkNV
bDtHXTgaLnaXbD1ekiTWG7Pwe2hQCz1kkZRaKzeloM3sYQIhoQzYBC7ozQ0lXeV7
jzhIeKJgB87B4Q8z/lQM4xTL0yRdIP4j8eIGQZlb4HSmsLn1qa6UD1HtiYbv2ctK
PGtVLBeMSoCBXcykwb73bo4lZuZ5+3Z2m+PpVdWDCEVu3rQiXW7axt/P3VuOtWyu
Hfruf9UvQbGGphfzv2G+RkswfzxLTjyHGWNu/c93WjRQpiCEjXgGZ0sTIuQtjHqp
deX0/ypshk0Mo6GvCurXI+lkWIGhPhwH5wHPukJKGJbz7UzyqnnriBCQDvL6BMQU
G9rIrGUpcvLAB+a2w/20z7sPp981Dy5i4qTKXLF+n+UTnJ+PelTkMT044Y0YH+hu
tjarPvQPt2wkHysy+R3R0qTE/o6vlgnBBnhssJydwoYLYPRnQ/3u+1qrXMNfVHbS
CvvZQV5FOosVtjC5wSY3STTsaQRgMLkm82eKGRC9GsKX8L5BZMontdvrD5hGYNe9
JX9yxrbyL3okWwKjq3G/jTl/6S3zTFGQ/hr2qi3mOnL9B9zYAzYe2kRlswd0aFvs
Cn9Y8IjgGE1RKiVdoBO3WVAFlfgotV64rfMjlF1EK1y+WeKIO2DB79Emd0iecPZv
SvYUnGDhdAWlPoQexNTscp2BpsEBziynPWl7ExwxqAaQ/SwFL6zM22KGqtUuAwkG
0g6mE9XwqApSCb+4HHFauDDwfQZApfU30EiUq27Gp+TpRBb6n+gf+DuIad/nX1xr
9amHmRI3Wd3Y6uPx94aVKXu/VIhRGgkxyRBTKB7H4UoAwPBVGl45HJw11yLz9jzZ
ne+rVCFzW+XbyTj5XPGYdxWDZ3H2fAkziR0fSOwT2oJAOzr2hMHn8zKAXmGWwVJv
I+PmPJTGjFfmyZSlV35udC0Lw9hP45E0EN4RLMadf/R6LxlCsukxd3YLqPRXsL9v
EzImwr+2u8LMuhDU4L9ZEVxMErbpZW33O+uRqK2z/2d0GaCpgMqnzXXd6TKyim7T
9RPrfrxSsBDVHZL18U91ToAABJTwIlGrMfB4X4Mp2bVYUjE+bQPWC5coT4mY2fnK
Yk5uWbg7kmJbOSF9sajBwqPWfIREF4K50m0lUK5h9/9NMYU6CyqtsOVzfWsLfeyK
2zRgDS7zF/x/h6reCo8AYQzHSATGXrI3GfyELmJ3uxHY3ASK84fddtSQAcjThWDB
yoHoXQ3lWqfa+OZxANsZSB1iKSKkVB51VY8JL5obbYajnwrp6NyvwxHLzkaCjQEQ
wq8T0awdeDdSF9owklH74yl/QVj063Z045zsQyPir8ZRnY77gFezYpfUZD1L0uhw
4TxrpRb4VD5chUaPMuEqTFFsdcbY5AEG3uC3p+/6uqYrE0+ZLnul5fgeSotLLsBS
/wCL4c9O5X7k1XjbLjYz98E4SEQF6nFf4EZyTnBKBql6JLBrH98STu15+Es56Ilw
+ow7AWpB4twEyNHYHnt7pFbyXtlRNXAcS5vZuq1xlJyTpgOfYqAZOTnP2GjOQYJQ
cmzpPFj1Cdtot79B7T+RhnGK9m/9QJfkl3bYRDnIt6ebtvMVdlzNewRhwe2jx6d4
0b6R5x+szemdXGOkWoamWHYT9ZL/tJ3Rl9QMMbz8/BHqhJB2RJkvdNYGANRRQ6/h
qLNLxRp14hN7MaT2pxxMQ+YCsiGch9TrPuNiX+SBymbJ+oUIN0jKnGYFQxufU/Le
J4XPBE1bEQgDZcPeG4qlthv2gn1DX03vnW0/ybd0c8B8vXGEQqcd/EAPn2NLKO1p
qP+D5bwCNroz3zkd3ti4qNtmS0MI4wz+9y1P+8ODNsi8sKX3n3/ObCoJ5v/VFEji
tVSzFVolz/hiujGOK+Si6qKLlBbe6I9DJIv6DHyzmnMZT8s69JO0tiVsBm2Brpho
59SFXfwWQeXl/sRkZoqVf1kW/IokWGKj3FvF8qzL7RZrWM6/zgMgMt9IMQyK7TD8
BMB6P9dvITj+CkQz5MP7SxDNCkVDkjYYsV4Qxl9OBCQA8aRlRWjwWjH6fL5lzW47
vhZXS2z311r7ZkHIY0q6+mVaNrsZCPnSwEiDD2Q4SCu9NZZ+5+MSgB8/5cGT3rcJ
xHNTF8wuSDYqAUSShHdadMa9qmmTV4MgYAy/SmxD8YXJLOtCuqbIRLa76dZY/pjG
W+xuYuAzV6WXVh3cM/uLjWsz/N9uziRNp/CmfHCom3/1pho3pfel/c22QUdJxmBs
rn1R0EtEmhlBJD26JD2qiOyH6QdutgMHk4wrUx/qFVtfISYO8y4Mz4rL9gleLxeh
yaaJ/FGML45EJ/ZPDp9CLIFQusP6d6kBuPzStxsvA72s9dWf9fhvs6FyBlryKa78
j9J8YDaLE5/anyBPkSFvdWPzaAljKe9p/bAle7JiCgBu1x4ldT/CEK2N3N0Rp19A
v17PvOOyA1NPIv1MCmJfR63QdMu0uu5WOIrYCOngr1pM+QDVaKjxI/nfKuURuWlz
I3GLDIRU/uNryx/WzFGMK4Hx9NSAZkhajZ/9EubO40UxVd2NbfZv260mYpmbpmZa
GepNF/asFiRcADVYUjAGQQvP+o+bEzwMrLCo3ol8Au0JZYwR0ZsUOnmvcE4vRC19
D3NhXKqiQ3FUpfGMSutn4fE49BhNGxVHAEYdi8U8kq15RxrCxzDbu+4275fY/kKN
oX/xu16F65x7XYeHgGaq9QFLb730rYNndfSHStEj9PP8qrrwkFg5XjgrUrgDExYr
+/ZY8KUxAnQrOlljyUnLJz4CBG1nybbYO+IRO/hhZSkYpYBpvGsiOrAl9iJ5PuVj
7z7TuHwvRPU96QGUjN0+9PCWAXsiinu1A3jm9ykykeiqoYI8BOilFUdLvOoqoWOQ
p7pqt7AI7RhtCslXuTuxAffLCjt698UjkmSio+w4jm9nHfnSWguYzIfczwodARyQ
8ihaDBw3en1FZMs4Lw7t4hZpgcisRgACFGuDTjP63P3+l+ZWkYyskHpq535EAmrr
LYBrubSW8tzNVkOMNZwl8g/gMu4LCj3yxa+2fzw4epZcVzH26l9OzCDl10oQakNa
a25ZI5yBWnSBwnnDo92WFh6hOIGaouvCDl26LqDzRw9kNFDSPchCHow9nec8867c
V/GWZBpIiBQn9w4NAMet0+Pt9H485AGO3oHr1dAinb6OfBNZvHJ27o9fL9CspSgw
ODusIuTRCZ5rU1nwSifwCLP2oeEewgfLXbyTbIA0YIkvXDBIAzTjczHrv6/bB9Hr
mV6+fM4DSmLY/2NnUrKlJwuKR2nvghlEYEHqR5eRol/ntd+HSo5eNdEhXJps+7Av
DWjNfn/4HxBydgLfGo5YTalGOm9zYwB1Fz4u6zq96ePeVpIcULN4ccxLAJqVkIUh
M1s2sahI0sVShlWadHQJquTueyDkYK9FrbNNIVpy9zB3yAwtsrSCpSIEG45w4uhJ
TIUEMCFHorjvHUkK+xGS6tKqQImNBgeCUrbDHYW6eZ6+jUHMA4vtaacLfJdR/c+h
rhBsCNOzC4g5XSeEuDkAA0RV87y1VhlhPQFNYbjJfG3O8QQn9H9zfoJ2kuS6MstF
IApRMBtf+ki6HuNtk5u9RkAgBNzTJnzvzkGZy/rbMcGfBVDMOAJ5WcXjbvy6BUgL
IJbqqygS5xJLgre3kyufWFpCFhUfaIgv6d/3MJB9pb0RFjjGzHQdl5Pi8ka2NEX0
t2g9FaLpHGizpc4BHH0rhxHU9BYxyF3NKfkxHyswkCOG8jUTSmteiHHlN3iBxdtP
rzVp4UMwPHD2L/JugCq887WjCsEotCCIfLmlzNwsS+c72hNHBRmKydZ0eNubThDO
War30fqtFXp4IT6HKidx+NvJUti2h6ah3A1GXV7DIFsqqVPNVgHnRnl5HpWEnfGA
ZZqkUr5dHM0BVidDwwlzawGKJsP1OYVDzY3FdxZ2RRY7qQuS+fEVgggepz0eHgnF
Txa14Kvw1npVyLYVkfNJEkov+j4hGzbG0Hoqu3rjB2Sy2VNjZopu3EwV53CHZXec
Vh0RLrppcPnS83+BkIKJfsHVru0FENG4l+EFbxKz/sYdIfP5957uhq8xsnnbAyip
Q42FpbK/dPMtspjPo97rks8Cy0+Lu2+qsvW3AgYUE0boKoCZfYv4gLvnZHcIRPlG
IroVzbdHkzCw7/vxuETf0Szffrgu6DlgWZthf5V2DWXVavceUXLFo0b104Xx3AqU
fpuP36F8lo8r6X1I/kzyKdnI8OrchsT0XXLkk62uaHU8vmWJTItDYVz/YFMKJswf
NcRazab4ur1YW4Imb/a39+fERuFPbGtPxKoAQuPCrHY+zOyBoOm4cDYQo6pYY/pO
yUVYsMdaxqZM4ZStrw2Dm1yrH0mM+nYJOdmbXG4qNUV9EWigGHMeQE7HxDym4yE3
+CVkZl3jXuOeTYe2uY7bugt6kC8/h5rDg8O6NbSIaYAT+PNiALK08t6mkSoZRFgT
MDxMPangAYKmZqMUz1ZUs2JjkitLIySyLpqiln8nnUHuwV/0B+aC4UY71st3IvRp
kmUS0qKrvasxLn1ZOCMv0aIXP1CfyTKaSOTh0smj6ZmR6V6UatouI5s0hNv9fUIZ
R48rAZFm7KKImiBXmwnZBDKHdPfs3DPIPk8WPGIDjlIkHxu9o+TmrvZrEKANfih+
LGSBifZRG+gIWQbLLvsH2qPjOTmuv7xh4YR/I3snPzvA4lzZxFnLXaGbQierT1VU
cgp622xdX/c1xcVjtARGoRnWD7hkvQlqul12FKsmjlNXPTlRLaXKrtRoQBULKTaL
8fK6SxLxxr1oU8e5RDnKiRqdWSLzgKe+XzZ1553xceSreV2zFv6/C7vUJe4HPgNy
tMaVO+uF68shA61wSJ3oot9kxBlgw3eZ+3vfFhx0iHh4t1smCY7t98dt3r3O0Bbc
2JF2sRTGnLSpIxOVFCJV2YyF7Jr8Y4WSDaevNZeLs3O1JUn3NiEapXTi9ztRA7uH
1svcKfAKPLJkTwFRu7FJMyZPLGP0492hZhwb/zt+mA2urY99RRJx/JzHyc+LTqBb
weviwenYG3TnbpOrV/2vgd1IAB1BNeRjFskqDxgaFQLbg5GYowAKeRzu5hG/HZJi
cx0LMGZkY8QZWBwraeqnw/jMmPQwVig8SmiJFGj6Bq7EHbl3rLpBw3ibvatfnxNa
CZ1zfckQzVNocrW8dgzm5YmL0ZW0xqbcwWzyDqfOF0LOs/PUGek2PomVVTH30MFP
8IHk7zdYrPiFWfTF/4NHOdFNyW8dJDtqv+IlJ91EIuWh9x7Un8yoFC+yCW+hIKOt
qYFaAWI+UtzD281hZIoZ9IEuDYbC0CSTkwGUUcOyPumClBsSxFQB4t0oDcnIb5+y
qgjVHomsLYPuI13iBE/ZZ2GX2fa+ORNlccqaneWpK8XO4JQf+GgFTdlCvFK4dvw5
qgmqCYOW/KibD//0QQQYaNVrbkuia1kGiktec0yz/ZDCLJbmCdHOOtP3ol2gTXxo
l4XZGlbTIFPvIvXyA1+b/ORtiIjwLTStmpq2VcKvoO66+d1ew0524fgsfxhYEtCC
GlZh/344PivOz0/MkeWg/b5QmlrLqkvQI50Uxfuaroc8KMGD/sUbVBvwtPk+8cwx
MU8EMvgHIfw4efOIiIAVo79NZuAPMEcJZFoOuZgGq4kyloRgKrDbalLEqNWJHSQu
BIZRe1dnf+xaeMbHnJIjdmlfr6GCRAKuzqAh+iFpYT6NPrWw8cuJKLyrDmdVuiQd
Mf02qdc1X5NngyZUhWFf0ToZbDAbR4vq6BJBLA2STfTt5T8fFctF8y7/OzRDW8cT
sHTr9Xh1iq0JW83OOls8uqr0UXysraz5WidenRU511+UjqqHPg+HsT9s9DB2ckfS
2lN7cYW18UjLZGe+kl14bt+JJpe6cszdW61KHSqdY4fhus1bR5aHeGv76hqtCO4G
VFV6e8q9GtTpqTSyH5m4gvW2mwYNVDzixpqplC1L1r44/If1sAEp1I7zPcdprDgC
AACzHqvm99nbvQp6z/6KTSC7TGVgBGq30z3yxrZahs/2e8Tn8IiN5VCJsk1nmajs
wnHwYfk3cvpcjYpXe7BnykRxsPVsKrfhW5Aw7FasmY/Zo9jRBW4Jh17P3U6ICTTL
32j0EOibYgOxwgVV7BRxa8pGrJpDjBL5hhilPrzo/CBtzrIzwrKJETwZ/un4D50X
kP3TMkMBXIrufLjS7c/3IyVNyERfAWzDDwQ1HwEDSYqcsnyM6x86Sw5OXd9MrjXV
aEjxuOyBCb1I4m8x+OCEe4IQsSY7K4Z3zhhaSE4IcB3FRCJi8KpUW7vV0qrt1bi7
03+o47NhKmHZqUbmqzv2NyHiezHSPZ++01fja7pcEB8bn1xdIfhk4rLLZRe5IqxY
nZ1uzQrmpEYS44K+EmhithrYZ9ppZnh6qMHpzGoufyAqauS2kvZUGLXykKFBToXt
T8yn3PU3AW48K+BuXCA96DnrF3gNEnVkRH3VJITpo6+fL4cNA0He1fXosMPq1AEi
1nFrgye4ulXZcBfTpKDtUzyhgqIwRTUZyArGtwPvi3EGInOC3qi9DdrxfZN7Fx64
rgOfPYRHLpn+b/G1GX9gdC9pboo7z/iSUWoy9DcmREgl+Oq41z0XmGtP6JKWLf3t
32RKCuD0F8Q3zgxSReDiX3xFhu4tRU+kfgdCjyclFRMoIEdwscONwT8YmJQwmgbV
oUTuH2ywFyWpAH+8kohYBevIkrpt+gPJ4OswNdJxgCGXog5yCQZii3pHn8LLMSZC
FJBNPjmaFpK3kEumR2jAoSu8RSidikL1lSsyr58qpVjMyuGNFm/0QoDzy+gY7CAw
xJ/BMxXRWtmClNM4xUebTLDzqmgkFQV4nAiEIkGB3kD6MYlNubJTwxerMjHU4Tei
6fIN3hwZr5PDbWq5KF/x78IcZuBPei7rU02wRgNryV6forDFUT84olVTKfGyoft8
uKgyYo2Evr90nZ7uW50Y6PKb4dVyCZR91k0WvExgBPLPt3mKiXj9UXiKsxKtw/Jj
S30Nh8mNeh3ZImtHxUARQBcsuPuMNEDnnrr9AG4dvEx2AOlINvrFQOerRbipoYdS
YgsfbQ7nHOk4ywWasYH7bgMPOsXGkBcH3+3M/3Ag43oPJmhkv4+3Vq40jrmer++l
ZZpnoTyczt2+GruD+JB5CyT1n04l43ynKJkhz9OqXMrti6Kqpu+x0CIHgXD8ctV7
dSryi4LMaIPhw5+J1gUOBG8g+ezb07KTiWltZI8yyjAMXSu9HBHkUscsBu7fsA6w
E1ickMJGKDPrp3IKgneSeJForuA0KPJ3DPnffWXku085U1IrUEh1FF32oRTKYyGb
0PU9kD2HvwhcQafyYgojfGGYNlOck18ZDJOcXMb+cdLnfzFdTSr41uWDPREISFVM
0G/28EwAPPpj6H9ZcKwYJbahECsctTOh0LW6EbOjtXXQB5MtQgj8W9bsJKtl40/1
KLl8UwDx2uPVzxjJCQuKGamTE18Dun2vaGi482/FJ871+oLX217G8XcibO3NqYZm
mUtQrjn/ulDKLZkZRQ8ZdrJLJ3cMtpti5APgsn/Rhq7YmaeYaclJJFDBEnL+6vSJ
VVhFi9o2mbPgIQSh9dGRr5J3nbbtby4YEi5JuV/acRqSBHy50D4NMigz7mRQ4K0g
WMMyg4VbpXGTcanH25vjY6W7kE4RPimxBVmECU2iOaS/y1xykgHWmkBWZVrKOYpF
RUVFy96y+4irK9ecRJO3uNKEvBS0/RUpZk1HqJDGnNGgMVsgxOdN1zcmRqRWK/mo
Gta3pMBhP6cS7SM3XEd+NgPa7P3dcASsg/6i5/AL4VOUZHwc+shDmR/F4K8li7wv
hihKb7FDANzuqla91zS196nU5qm2/NwdhnyX84VzXUVuyLZCYTwk6dEn4fxSvF1N
lxngub7fe8T2CP6QpUE5mxgMP3TuiAsLsWgERcouWP+E2GVbknLNqUS3i9u61CBd
PRGWkjnvhFk1EvcUug71wFIlNxzSXAfnspH6oAQtCbmlIax0XLwzZGekm+TqSZpM
9/D8ypEnPtRQS2UHhP7uYLLqwilrPUh2NAl/3kUTM7rS99gmul2ZynnPyjsU+RfY
+c4SDE41fs9bJSn07pMd7Sfd4fKnzYmJyFi0w2BUf3rnzkvF62p7TshzgesmBxkX
bGUqnI5wABdiZ+JoAN/m2adOtP1OBxXTtaMWqwEvkjiwTlCDYcLcpXbzRI//B0nT
pGA0CMYA2kjoZA/HvMvcPtIPygVJPoDwrOTdbtXBXoS0v2kzf0ZJrlp9NO8SldYA
Q5vqdAtKaWy86mDS1DOvrrHtGtI/xmu2SRGg0jhBNO6HC0CkBJQSECZ2JT3Lv3u9
7py0rQoz4MNVrMlksDzH59bi9xKaUcpEBoqmZgE0891Gh9WXXGVJm5Ggis/YwKZn
XHrvKYj9d33dh3FMuvYn9nj1b8GjXSbSaYO8h8yNHI/2Zn/FxUNysnPR0aWkc8E+
kz7fQ9J8tIDEMxb79o7eYFce3cKpWTe5170paj4PWoUKFXbcZHI68HYv0hLCQYkJ
71n+CGAv3Iyv9VTG/0q3JXXsSrtwGzQ85Agm5qWfzQaAIlHDD3cU24Vnj7xDN9p+
buReYWTAPw7devZ4E/diCW9PV7mvKcgwPvVqhxmVBp8dy+tps4Hs1l6f0eKzdRfg
bDGHJrURc7p7wzmJSnf5nzj3VsS4C3rfSBZ9UDHBzm5FiMtxsPFvlA+YMWtrOQPQ
k7m7rqO1xBfIXml9+GKsptaB4J4DZuBYJT5ASCoUak2IHo3z+BKuaL+fN7WAaOj0
NncHVLEkCtdve9+FcWh+OYZStI4zznJUtKwUyencv2/2Xf+omKY9ZsuMtWBdywmC
lM48LiQcpMz2KBs5PdqtmZzPODc6WUvo45okMur4j/u6CuUrIP2bdVMK2RE3SYxm
bLIl+19dAFsuwKo8nIndWjkdxd43cP0pt9e3dQVnBKaE1Hy/CBmV81nXp2g32Jip
MTgbbPyvo2vqkr5nYI7taS2434Vmt2TZUZ6Y86vX7Vb5CW0NWQbEQqIPAlQUBMgP
XT33GExNMR5dsMvJS/Go5VzEikkyVDjw6D40Ber9tZoDvW7PVdWjB65lEgBqRxxb
sNJy0wWX9rIko/JVTjnkQ80OG4j3/eRNT6IxA8hHul9uYI33jdGU6IxQR0ZPfCIh
8Ne7E89Jna/N2RuaUak4FGG/Euz7VTv2WlTRS2VX//UzHDFcXCEG01e2eosrHN05
WixBG0AYvACE0LDNiGCeVz6lbX4De0F+TsdXEecQpiD+WGBPfqjh5NJrlQHgMqzB
fs5PDC4vovBcI8d1lW7cOYNAIh+AhHMzr4kMuNL7sfiop49xUf4uKNPgzp3I0XrZ
Cfco9WomIILDI1Tza+QnN52edxCFKD66xQiv5m5T7KsRAQm/RU7iK+ung7cXp+w5
Pcpgliq1YB/Fl8KUwCgU4+7lBM3MZZBqicrsPki77YmsjBiEFPTSnmI0/QMym+ei
SLt2yMbIGVrryV7ZZtrdHx/9AVe9Fmla24jqh2RTl3bysCbV1DB2d75gpjbSITlL
lYi7BzgdFuK3ARsRnLJsLmxuWPiqwVaOoLvOaKmK5XqwbYNWR9LZCzeIpYZXQBB9
k+9u/I//9ovPVA95Pr8QbAhpvGTyCKZQXOA/1rgGjUR1Sh1Luiw+UBa4PaFv1jM9
xm+RwQ59YzQWgxQZaIHd8pUuNidJFOGzvxvwWacRzdcZDCoyQiT0Bzya16BMvukx
iMRNiVxL3VVZLfoVl7UB0ceGdjU9UavskIicl+AvYr/QCs2i0ySqLAowiCzmdays
A86iV4Pine852rABPezQkc15Bv6/kfxofU9gPDVOzXbcZQSR5Vc7UHETYeHFPobj
3UXxtTbvERajbZ9tR5NgA+FX3hxXag/6kXUnvtA1INUqGO3xPbA4SdjDJXTBLWHy
R7rM9ISesSnyeyvBIfkzWkvsHGJ+55SNqJF9k5LqhYkUG1CPSQ2BngdWlbYlrnIh
hWk22dMH1nuM5Jv8Lb8G6QnNxuZJgin5nGXixx8mhsixK/rQHkndaKIB5PC0cWRI
af3YT0lubu/BO9i6mKAjevjvXwxbiC1f8YDVOf5khW4rGupWN3ZunbwoHLHpS1UU
bv+oy0SZGV8cIBnKOIwq8KZTjwMFy80aEZQwvQJuVFSqkBkzTLy05hD+ewHCTGot
wPnq4BWV+dXkeCC9BoZSLl6Jmnbj1sSBPZnwiHqeONMC6LLekQfo1FssB6F69cJy
PeoITekWR/C1UK/5T/0loutEIv8QpBPc7stXKxgGiimgj9h/4dS/Gdyf083v5fnV
jbjVssUMHD44cdB/1u+azWldrDQP0zdoPCd6pB6rViSt4SKkUyDLaFozSILnvsy7
TXFWt9JuTqz3rXu+lyzzM0fLElCSnG23vrK6RB7bRsLPKIK0BLiivGtoYAp+LLpM
hZBSLjOafXk79bWAPoZzksC98VDVATdBsF9zTwhbs2HQa8eofsnbuPzfRLU7zADX
yoesFGD7W3XZWpYjQ5eZ/N9r8lA19VuUxHMVDWX0/xyvoAljXnlYbaaM25xw51Pl
4SYEyfARooeGvySKm6qrftoflwZbx4S77piekSni7muJ94esbkvJeB/ZH3R/7//L
J30et+Gb1wh/Ngyzt05eF4YwqpMFsIptKbVrJNfd7qS3cLvsKmOSyrHZ8+N+DdGi
MKWPJsv8USplMPBZpqIkz9JhlvBj/wMM/T696J1R7QNYZlTl4ggdC/zXfXtL15Uf
ncShmhMzH+4lFcT5WCCH+KyqzJ6tPazUnR1/OqI58eK+ZhPEKLhlb9KiUzmWt/Td
rf7H231fCQMmNtQyMb0Zdl/wHWRUy+PDXhnNtWGjln+Z5qbZ2ehGgKUiujafi88F
yNhKgXO6eypxKsxuHN+Th0cLwHvfvZlWXh11DC2Jros2OmMZruH1Y1g5JEOSp5Yw
dN9RxWO/2mXm15z98twj//i9A4vS4cWFsjsxSnM/LsplNLJzhgnAkZmc5r/53Z/2
pyL0viRxfZSGYLMhcTmS03XHOWR/SdLjbvcEfygrakx1b5esa4G4xYH7NwaQv/4b
qYn+N1HemFBG0XlSYSu2/ih0KzSZD1WsPUn3wC9d+npjdE/6mf+L/q9JJ8YO3phP
eRKR2RqP7enqMdHEGXZcfBJsxnqkC3v95b3SgJtJaqiL7hMy9FhHNkwmZipdtjMi
GBxY3Fs58aFYZvZzze+lx89VfMEVRPwRFxaamE3XUkuJAikJGIqLfnZy2jL4lwsY
n0aaB0l62NekczojcTYwM5JiYB43/rB7qdPyxH1LTaKq+55ueQdxGbSRsXA0xqHZ
Qh8uyTxNYLyWi5p1XaOBsqrizhaJUxqYRwDcn34hrLlHvl8DQEoB6JAiuFVzsf2C
XblcqMvAZT87RhkFw8TOlZj2DOt0+rsVi0fLUaqyyoIAorwX8nHCu88jVqrtK9ko
auOkQYgHlgnH5xbEYwzzVDYY5idi82UbrA+ped2lZ/Cs2w0x2Zy9cq4BJ0IFYovC
AuzN7zI+tGb8q8/apvAaC39R0H3DNbaP5BLrsTcogmLAUYs4CFQLifaRpYcBv+Yb
EBVoMgibGDY1jVTng9QFYX/tmPk1636U3k0MQFCLn+jVGG2ya0D6Z7Fl1XGQ838J
Cs//J5F2LFYdvXGbQKYrZKOOKN/6lPJc9YRe1Z0RcianP1r+qrZws0hcOiptGHlP
6MfnE/Trp1AL3lsLvJwuTPjn0VgE2EgK3syD46awMSfkEq4wsoqCmqxqvGiDw4Cs
Q8bX22VxjURc/03ry/Mp0+7LlQU00PoQ3DuR1XxsLtAbgZgCfMLAcFWuMmWRIseU
hD2c1FUF2NIV4pZxNDubc8t0QT35j3x2DpoCGcUkhMirF7vTac1CViZoVmhTOjMG
1wqen5OddU5U7R9nih7M2WS4HUDeHEuY2fuhyyTfPrB4RIbLBqCkiRLX/djQ2top
zFxNHnr/43wtk32/x5eebv5c7XKa1i7B6VQLC5uFcBU0MM31d1KHYLK0DWdRIP2Q
APxBP6QFpK8arPIRuy3dSJS/wHJrBUG5buZUf80e759EOJUotDgFd14+p+VHxt1B
gX8mL44Wi25ThVyT0762HVm/1uR4dXv1oUJOrTv6mIyfxWl223N6c4ADL2QQDKOX
o1YM1WeIsB9K2/wBSkl6h0htGKaRBmYkru5P5JjDaLaBINdCYd8f3pMil7c3B9qN
pvjCzoKBjlTVrPmqt5qah7B2a1TQR3kxY1phalRLb4Z9KTWm8FB1r7rJX85sz08z
t9dMsFr8Jl+0WrEDHQmdm4KIIPv6+OqlZXmKqlFGKi836666tf4SLnoN/KemSg5W
Je8S3zRCqmOKDyG06lPKM2RPGnZ3fskBEQK1/vU8+EDVF024Xe6ugib1JkC7oR2l
P7Ai9OQO4vrF0Th8U0iovw9HPRKV01pNjbwT7naTSzTlwgr19EofLQ1b7elpYkgI
JZByo4tOPrsGNYYUzTaj6mPu0/VNLAADZZ6h8L9tp6j58plsqVhiMDXzLxZ8CuyK
LCHhk0xhuEsF3XNaENk3rTf1aWXUAY3fic/sn+Nn1U+Y2RLyOx3eVc3rEUk7RoUy
94ulENhUVkZVBdc7AXb6Z5LFQ0gpMmA3kPvYqKuew+F6IBRzsdK3ILFJq3YUlGhZ
pUBB6xV86oNY0djNNJ/iyGYTcE0yrpZhy3l09leQnnd5e6sYOcbfFx0ug0VXyXjY
ngRoLHp7pOyKfRZN99jChEl/5HBFpMvSUgCu66TYrxadfM97DvSZ+zAeEH7vmWIP
Xj53DCyvlnFJOPRE2zDV5WrJhU1mVVaiLsv5EgLAwJv88X5KcinbXPe1dXG5uoh3
MXC2N70FYqC05IreEDearrFCyVK60Aoe2yWqA4DnHF+HeyWI6XhWVWA0KKTYx8jD
SHwZMayGpWn8dUPuoRo1vQquHvQbVQ2bWFhWCM5QFycTxyUpqLQTiiDiOthif6Wr
Z8nYVdEarcgpOMrW3JFKKMud6YF3EcZMXaswZg3yZ/fbqtU5KJsRFB68i+M+jiEH
VEbcArmBXfcuIe/Ig5Rxsefr7/U9rzyYozLAsnhsNy5eJiVdLjCjJQEgH4ABpqMH
fVCPJWZsfMLphF+taT15N4Vp36B62OReshZ7vrIi0DC87GfeK+zXbUA89gdtdsas
X+UIbMpfCbIU/eAAGzxYZ87pDeWzz82oJiCwV4RL8Sf40rzy0TkqCOaL4Bv87SQU
0QAYdtGvPWNJ3HcK7iy/WeMPZ9ztIMpFLCZmZm2NnaGqK4qfCq0Cr6kt1ZOTH0Ay
3xG4iPMcCvLSusZIJwHOqabJnQYGroJBYNbbNajGbkW4cQo5MmFWZzHnEzEIV6v9
rHQmpwecx/xJvuN6Dh/9VSRVuh80TGDwzKJP9Kc2pU4Jyvc1xGT9LVwQua2p/5g8
506r7YaCKKmurYGyNQNhLDhr6/aqpgYmi/rz8JIBWlvt9zo8q8M5g+GfsgW/NJvy
8mKUYW0UmcPJcr1RYJAlvEVfZ/isgR0YVnhqZKG/tDNKGtuwFhwGFJyFZuWUJLnm
pDLpktJ+IR/kMNdsShtrTdurL4c4kmbinYfeN5J6shOWuqjORbnO256q7YFBaTLp
7k7zoRvLroxh9QgDv9hAu9BdAm0ujwFylAyyYIe6EmweAmT7yBLlPUagj2ph/Afx
wGxUfsdQO/miiwgd098r92AgciEMOLwV+J9EJsCsfz+m5rX1sUYneGmjfSP7Q0Cd
UcAsSn2ZYrNTlzDpHtMDqv94pkFYvNDdtXBQCoufqfdo3wAU7wsb6UYHwJzZtuEJ
nn8nVWHQcrLt3YjrLc7M8yrPehJPNoWMu3tAMc1vR67cyzYv+otfE69Kems6ikDo
iJEYXAyoOkqW9ZvynZsLAVXo9dIotjv5x70lRa9foIWh361XEYadLkihlgXX751Z
W3XMLhNCrHigWe29iX2ckl/5ked6fOVe3AYS6I8m4RkgHMya7x/ccg5V1xLbHedu
QPH1xIikyxUKAzC5+ST1PFHbq1+SeHmuozKw+2PA9SrclTOPtIJQLx7lSoanqkud
HRj0BIDuPWKEEE25XZNspjSM6te/ZX+SvxF3n6kWF3aj2t07QQLNvYwFvsZPSNrN
mP30i/axVJvtL7zquueEunG3tZ/auBpz7OEcgvNgUymvUASVMhdhKoTU86tIs9pI
pDq9pK12mjQNsC84eD0MpqGrJE0jP70gpbCXcnbMmgRZBuM8VVSRcWWoB6x/1YtI
XyeQmMFrbeqiQHu4Ch+18k0tRMa62MmmquIaP82d7iBnjdfxfb1eYZhK2VqZ2yah
wA8ZubDzPW5FHV44Awwhz7KtNtYpAstG83ALFpddekhhXuvPPBkIea1JIwk/XLSj
/JL1j75hiwzVXvYCgGvqtVaT2tgrwfOFESU5RSC8FBGo2dpPXAcCbJrVO7r6B+dV
Uvd0IGCc1ltVnBM3USGBnCN3PoUsUgsB5UrGapDzdRMxSF6GpOtDwEwg9WvEQtGZ
R3iCuT7a0QvMgqUVMa96RCAX/EF46hYvGBuNQlRMynpUA9l9GMzGpleHLCaB8q3Z
Xs6qWjdJ3JUceAWTswQnYCf2iNtBQMeRzuAwYE4ow/gOC6bdKbp6M973hOXK2GD0
sxeUhB5E7ZsFVALGJ2Gon5MR3LS9JVIC12/AmIakg5nkZKMIJGmMmrdi5DynAtSK
DHafp4LUzcW83NKphBcUPlVCWfcWvnMbSf7QMHQBR8Z6sUf/NoLX3Q+IEqj37C8j
IWEmrqsEf6Lo9Z5C9NUAEMB8la0xKQTPk6CDTHFKtuCDqlHXGkHmKUTUC+ixNetD
9hCzceeQEF1L0onE4p/iW+7g/j6POeKjzzeAt2CKSuVqQLPpUP86SGfH/522OP9e
WVDcwtwpx72tUn12nLAtu6LIA9fnulD6cnxD0Qu3nQnAdh2AdbcC6dGBSj9eR2iU
yDHlnldeH1Iyd8vT6rpH+PNBTmjRm2v33f1WvQccC3QnAIJ/CC4THppVUNO6eCuk
1JlsU3yaq4nh3KlTPVSdCsCRPSzL89IL9F0SseFP/+27NqOCdDdn8AOuKBADx7VU
cgvQxnE/zkEIKhNRZmC6c1qhR3FB7lq8gxmZrRrfwj5MF4cAKlL7v6H75+OueUk2
9UBNhAq/YVbFr+wpzJkeDbvIMGvxoCPhqco7AoZDgxKKMAh6ldUYxcvmsFOpgSvW
jbGUlmuXVq0agOi7O+bMPOeMpwSRvFlHD/PPEWdOMLfXFK1UZd5XJJD3cS26idN0
mn09rb8nSUr6ofPzO460fMPlyIldcW9YkNiQuPPhiGKV5zR1HXoxDfXqvOGF2/lG
5fiQ4U0wRmJLVSuHdW5FxuqMg8+ymCJAR+bOVpARDXzm72ValtEieZ0qWdom+c0V
0d5+89bK76n1yBQjfDCBU49qcBaXB0ulXUAt3lGNANFI6TjZfutY7qyCEYOxGc1E
9Wtb2IMZj+Efjo/yMq1iQ7ZEI5OlVhAXLBQQfewx/VXVXubvvNZJ+kl41yU+up8s
t07qy8UkFexPn0V+r6b2tnYjvcc+RvGYKQzYb1Ip86JZVUK/0DVnXR/VWlNj41Br
HyLfk34Mir1a38VYuNwBh695roK/XpPHOIpfRRHp2u2Z79/0zKO05Clml5vDfxd1
xmljtjO/xsFdbklZ/A/i0EqSWPbrA7MVlT8l1c5O8K+ZLfFGrSXkAp6oB3EKs9wh
tMMbYvadCMSWqMrRq+2cBf94gfg7PPm2jCV7wyyrQuC9Ci8J0Aj2OLRHDWTmjRem
1shHvolgntmsDJ6NX910t1osj2pmcHk1cOURQeLWZUnETbj0bQHaUsB+8VFkzQqO
QBqBzYnjWLpVV+zqgwmWUhzmBlbHFg9lmGYNXWOCsZnAnw91eAjSU7go98mdEZnK
cprORuyOYvgQu5/EudayllhDgl7IkCDMLo4ebLVkeJEzBzQByopG2woKPMS31cP4
xKocJFmswnbUL0oaf2NtwOKgP02n6zgZCDwfJlz6H+Zi/HliWqE/7yHP/BRjGA/9
xnDhuk0VqY+qFPcJ3gKNi98Jp0gj4X+uxNb/58URK079vS1xYD5vvuzK25pyHFg6
XBx4wB2QpTlukfAOXKKmzUshWCFQ9ZK2p0ZSIvDZm8AAww7XrsTPGJVa0uuR7u77
Ok7Dm4dmYTw+B/Ul0um4wKnXds3roTlEu+j80ovJ9Z68Zdq/naTlFM6a3epzoX2n
mgYbHAxdftSK8GHzeIL3sjRY86eWKzdm8YctlOz7C4/J6ZsLOVeFWfarMwsZhKD6
k8nLiEVJWvfpPDM4a5sKquhUBrq/ygmLGba4Ud9KBdXlifVsg0MqrXIyN4/HAtVJ
aq83g3UfVcsJbxGBSFhwGd2FmnJWQscEN0RbywXGi2aHyACkauBSVPp90N9h/3Ix
+tKwPw25cYRR02460sQsWINWkAHvnybspIPrPbShLsbn29H//0onu3MeijF2JxFI
0G+uxyqpMHtpPrx8sX1Z5vFGSfTCppxQoK7tpHBSd50ml2oFK0l5ETTWPE+8f/2P
sH/H0088OMcHIy+o8GnQ2vH4Z/VUvVLGANyIGmchPczX9INw9vkeQCH0owKQnjg/
t1xlDnYCEuJPr+9rOQAz7SzGvOMNUYU/PkVyvMufO4ETmlpZeKrb4xbpZi6pahbN
PRGx/3XQjMglKEcavQuLOPI1YdHHPvX7bkK3cDFqIbJ5jLM3Yz9ADjxxtHr/ie6J
K20d0eRrLFncdei7CAQFM5tzwjvo84s3eSl7loF94R7k6OfFGG9M0nL1sWxJh8f8
Kz9zB7yFf35mHSp6qQd0L49Ymex0no06ZfQXh+kqiu9RYs6VCxav5a9QotfdVojU
EjaOyBvTFOL7zUL8PrAzm/phUe18KlS0eVjNtZ0ASerEPntiehozThd8D2AFUstj
dk6ar6MwF0yB5Qcu2GNpsFWvaTDSIMzemVedxug5o2bEpc3a+k8eS1JlSgykmw2V
fbKLzld+hJL+C8Se/adS0w+MQzNuYmuefRC8QAfxpldHT2ypKDkFw6ZCpc4tRa0N
E6Xlau7E9jXZNW1+0pjM4YnMHPq7gByG2CVJdN/5HGjthh74fUhDxVFnFG8hpsYw
gu8l7S1UYlVQ+4v1LB5E3UxOULQtQjZd+QK3O3Z7sQOhij0u5Ei+diZ9Baz89RR3
3X2GyrwouOOzfoW+mzkHEgildGtT5fvheyJ+pRWZlMyjUNJ3WRyLRFgzJnLxNjbz
zEAVNYpzn0GaaTGFSHF4cRISKn3Ssgxl/DPGGdQfxHky/fecJu1wImXo7CL0tGlI
n9RtN3a+UV5vEmJ5CyCJuWUtmeTWvu0ARXm9ZYoT6L0RQrvbUm+LgDXTPUtK9Ocl
ElCKglOeAInYJ/5mMJHDK2MWYSBYI2fgfFuPdXrzm33pdW5rH2s8cjm3htSDFjxI
3imOkyS1a+tNmvu/XKRj3sj7YTMtF9TE2H61f/bi2CIIkwSDxF+54HoOy+zUB8l0
u5ueCnmkNR0XLQSKTnPSqn1NIETQ0hKGGEEd/gyzPr/re+G++oCYpM/1kuoZ81Oj
CwFwEXZY93Z/0+z+ex/pPSGv76F/bzZYjtOgjMAuvEHZV4up+6SL5frl2hQxI7QW
o+6AAdycYKvCrD9WpsTlXXK124litp8Le1nMhxviJKrDCb9ISwDp9bBoDzq/0rJ9
LlC/oA3oOmuxC8B/il/LXS7Tl0MFb1DGlY4cesh7knY9yHwgws4QnhT+8dsk317W
o3dt//qL9DmqtaLZL9nFW03oatt/kTZ48QYtGe0reJHIkk35u3Ho4ToO6OR31XJL
K3fleupVsSOT//0gm3nnfBLdwG3qX+DrepG71ZhtEkZ4GAnPEvsPag2t0eUtzpLC
oadwM6MUfn547XooJxMUecjI7j+vEK+nVKkgxe/HnTb3byok+rNXjpZKr/SXNZBj
ZgD2VIlO8KpTUW17sWOn/+EWLYyklv9yrgYjEGl2Q/008FOagIEj2j3nQOR0ouuA
uGlODsINQwXu1aCTjnj+76rXaxvfGdW4cGUQkuGuV3qvIXyu1jQDF5iUsUCoL45V
Rpj6T7OKjZCzXogx9Wa6V+SNdSH9hIjqjSi0S2e1xnP41k58xhTcaSg9iuuX6MgF
xfPMz1rJ/8lWPJgDE559yRRTvvUjYCwdKVSbyZIRIJEhkKuiSfuULiveKWgVSq/n
5EsLtE9+/nw0iq6m9Z91KwwDa4HgOmLIezRA6DgIBJKDrURRr0464+pB64RvhiKJ
wMKChKoODW9wFW2JVzAVhn4XrAa0yEIS4mdx1gX9uIdokRi6dZduzulXq36yv3yt
B670NKvQUXio1n+w/JwxEHLWyvEUonLOSKuTSm7BeRd+sWzp+JbEVKZjE48mgNQI
xlqgYgf8S24EUhM9g99waOiqtbZHlzHjFdqgnqYDoqU0rW7OB6CHNZge6CgUQGWc
dJk0ycjxtTe+ZvW7CoBVeEKBayYU2y61760qYAt/bwmTLICANZ4p9EWI5dBEDlWo
3aXY0fmzCli/QC2bds1k0gUR4mcimZiFPyBHOnt8Ey+ywp340TtL4gdkAvXXBNlY
ZmpuCXdXP+BsmJwuv6A/ggZ8SQztMmIZTsvVQOAHzo2e/xVqyzyJ4aTLkLHTdfpB
WgdvXGbN6t3VIce1eKc+p4j9c8O+anpUuKG7/oVfUNftpiV72iIzeZEgY47L4ZNa
0fomJdnrCd71ThTJsecqM0TMom3J48Q6YQ8ETpvjSgifcxNb3j7oOTbgcR+X5GZQ
8laDmNHKAN29M1Vv1x/4Gt9fAKlW2bzJzbacOyKX4kDuE4S0CyppDcN7X4WMHIjk
n5caA1LqnAMLsD3tLEN2XWReUY/q/Vb1JeURgNx9KU8V12IZ40RPZBQiyV88sHR6
mMQQ64V/wYoEi96In7/YuxAZxFcVFpNRCEslOKW2/Eg3eR5cYAmHKhQ3FCGaHT2J
nO8z9c2cFOWg/keSL34Zv3bBZCD8j5mXqSZDx1mc/fFUEr4rGjq2iUIH7U11LzCN
JH6uwyeljwyx8mgYk1thHBWE8Tl97duCQQKGhvuChvQdvCgzJ9NhhisMAQa53WIS
gGW5+EucRJghVJjxhfsb86GQPDogUrrFc//fmfwh98GvUpFmSqdk4Ixca2VRBaX7
YoG1LgqmLaaD1+Z3t2bjmXci6PlTl3GCCKr1R2O7hxWvPT1vV2VTEzGvq9phyGw/
d5600K8PV8ctsfAl3hq5P6vUw+ESLU27wcDmITPu3rwz36Dg/ajOZAok+ujZFME+
qQDX49OBN+3Ik+sv6h8OkUAhgCkIKJHAkNMdBISiHLF+rPGanh/WMej1+QcaZrcg
q+X8iH4YAGUU/GBY5zQgsfGA/UexU+r3D/1sSAPfGvnbCFN+CQSK1LhSEqJ4H+1u
QmjB59pOqKXx7dgAzH5SpYlFCex1aFIWlj0kyFO4bYlfEikbT0QzvmeURhNm6piT
Jlxc4ND30rdJZ/RzFxzLGdhR3LGprOFNa+9qltn9+vHIF8zAvwNUFvfYe0uVwzY9
wAwSTKoixjvW2zy8YIDWB6IhRtF0T87IojmVjLd3HNqc/8saQZVAI3ZWtBN0eEoD
g/e7LPvWp8ONozQfgB+/kB6W2SRdY8JgRbgSRCr+T1PWix7nn7N/h39G5tKhxM/q
Z8SLvDkKCmpo9GyMzAKircKjQv4Dt99F1RwCTVbcVhYonYf9H/Xdbor5eWUPUtCB
QW9H3oNM8PGN/nrofV5rzZIrTREZm35lqBQzj7H93pW54QTBrPB3bUEugVQW/fwz
Rxy6iXDk91+w/4yCBGfhb0ve8NLV7OkV4FaObhS14+2U5Tqs6Q3hWgCemHQ0Z6ND
WvCFEjjdaOYVYqGGkXhswiTdR0P+wz4uIpZlmNo90TJiqfG5DtwFBGSoqv154D9Z
I7Wvq+BtOvwSJPRXgtMQpxnFHwGSSRJStt9Srqp+6Qdq2/mj9ODmgo669BBg6DxN
tyhYSQnQAshhe3MUIvRX8GQqt2OcJKpumjmUtpkNCehLtoywtNEMBKaXgULYSacJ
/eBJO9hWt3LX5JJBQ+xBk7cI0SHur0Z5sBR6Yr5UbVefKrc4ZTEdorhM3WQcPheE
EHe2QJt5O5p+IZCLFfY+kCJvbZ4Khj5Mg5T6FdntQK20SEI9FIVe2gZwA03Kfdc4
QxUi6BzWjJP3c6zk8xEkYuCurvBIib0xGOjOzFFrLRPOv3rYSe5RieLnamAp70Fp
SCRj2NEX6ASpifJMHk6Gta9ya1nAUVZpzS6EwLmnA8DcUW8yLZo9EWhpPRhBFXFr
HmiUOauB+SDR6rGiXgbqb3qCG9IV0RBL3K5+KpUKiVjabZGbkHjaq1lJGTlCbVsX
r6x54LvKJnwNrZ5drL9YrzBuxSyk/S1SFiCnWjTVcSZJWvTZxhrLbkH9t5gwlwlN
3O2LGbnAGqGcZv0Q0p+hJk4QnXxwDrUcqEdWxhTKYXWRfNp/Hz3O5GPfrTBTInPj
KpSYPcEMYsvfFzrc5Y5jnQJeDWPwU9983PiaUYC0JR80Jd8VRJa9FVn6A4QDRM7k
6PIarf6IBLEGz2zSNtMTYV+x9VjFIH672TlmRIeCDQYV1xDOnk3QivJmlIm8ey5D
WFr/SxLzol8EEWydXccDSfXx7+vestBuBPcjWbnvgQQ5T/r+GjoJZcfCeFf5DLFM
sdHhMGPzp/feYBBBbYk+4HcDXai4/qGQdXUeVcWOMKy5gbIt/qJiWtas+JZdFe/E
wEI07VBCTvC/Rd+FKICMYLLlzxDCvwMOkFt/gQHsepgcB7rkTyZgNpyVRcAXPUsr
69VgYN+Jz8BaaHr61cpzcO67BY3NuTvaKQn+cxI5W/hzcVOQLICvO50Bsv7TcooE
EW8BKdzT/2Q5ZINz6aJ2cXXS3mdg5WI989BjV38+jbO8yqdFpzXWKrlsqcar4g7k
6XUgxJcxvwt/7mygDz6yNwt0YPUKzrAkqC+9aDV7Est8cFPaYM+rI6ku0Hd/KYGv
GMAEUu+QGzXDRbtal/SC4vFIWcqs3uLjenOeXhkibt2pmwZFdatEAzua5i5s6G/0
3oCRZT/YYG8W/asKlrWkV+1zGiQuAjw33Mj40J/0ds0dy7V7hZBsTKctTWo4U2oG
rMlKCxyIbs/BMlQgrls2RE1hTa9uwpWYGARnRLWv7t+4yv9tFOQ8/7UV0l9nCg5u
7HDAqQZnWpuVTm+GoRy8fQu8Vr6AyvN5NKtFx8srxikynr78KW3xaf6s87xfnZTL
FlstldCmTNGDcpRGYRJQXCksBkAtMwxUrh9LPvAz8yPXMJa0pEf2hQxgLDx1I4Eu
nQEpzgftvsUlawWNoKtfsq4o1ojpCUsTNS+r//nrlwXvMW08/v0cUbWvExITT2Pu
rYRVbzzKQowEzvPy9sif9qd7gKui3C0450R8dXEZvG06237T1z/4cS1g9smQmMIM
O0cJ4pCcliCNYQhjoxnMx5q6m4I0+ypRP+3GLRP/sAJ5oRiXjTqjZGvQJ9CcStDB
N+CtIAl9vbYwLeSZQbGHJGIVgNhbi1nl7GF4GCfjUWJNowGj1uBBLY0rE57B+SyM
5sP6+3wvDpXoQU48phCknetzG0ssbcBfK+DDySCZ4FaGwKEa9JqFEj1OVW0NzMIy
/bDSWyJ0oklFCLFVf5NlEr5rinZu422U7DZIzMKEv9DzRAYwtTGBNNyg+K2D2OXC
JWO9Z2MCgSa+DIwNZNEwxXcErcVkAjioFDWOQEzbShq9jMRX2yRqKrkb+5/bF07u
j5sEogZ3Xuns0aqYLj46d0IQdTs6u++IouViD/XSc3S3cqosBaD120gMlUq8uKjq
5IN9NPNPb1UHVO1sJqJoSF+elLuIUVGAfG65wQkUT3Yb0DOLYSKfq6rwo7rm70FV
gf23vqqFwCF6nUG+9KG2L9AiZ9QehC8py1S25aDWZxSKibImjmseZ6Mpqf7M9pdT
WTdk+3slRnViaWyBtBPItaKQkeOUuqZ+/K8bybf83bsZe0pY6LxlI2Stg2thlADp
6nu91I5d5W5T+6K2g3pcNgz8zyVxWqBV21BOgh1EPBYgTvvBQhg6ToT9pZKRQoG5
gkE2Da5mXdUeFrQpmVT4h4/NGNVTdPQCQ7QI8bvA+4exY5dJJ9h5tfv0UoLnpSdE
hDDzh1vw/srXZ7SuJlfnGKuuqO8174Fxpr4XafGFcJhGd3SUYtGZAQVHmhqEfZOs
mFOhksClIycsB081eSw2CfYXe8My95XjrnR6bLUDHmAI3fGpKmmggezkYEm4FMwR
GYZM5b8LWjhV63OEsrlzudeyO379zJf608ZEEYko+9I2UNiCc2vmQ+pKUQ7fyMdB
IaK81FEj7oUI3z4e1TQnKoXDdLDOOpHuxt+8RmyhjhrUBDwbdSjfcLzXI+/I8yKU
tWx69gS32PBz2aM9mN7ZsCcZFkLwfHREdbKbABqF6Vge1V+1hBf4xPrgvkS7Vcla
6VQ/7w7RLK/RY/DuyIjq7flGa7RE5dniuH1SdDHzBDKTa0/nhM7t4HYW5z6kIxqy
orT/Ncm73+0P/ATQQ0/NEVaivMvxKFcBQW18jl9Z3/MtdPXaefIb03R6JHyfmxrt
Je5Ca0+ZTkpgqh/M07XY2P+Haybi3e2VuXz0aCM9b5Yo3oi+njpitq7o/Arjw8X9
Zoy84zvYhRVSF5HXQirOFiBBlW5KMX9JQjLGiMdNyo84UDQpqggbDyW/u1DeT4dT
+fmmb/zQ2PcxjzBjSriqov3qBgvGKYK1YkbhYLIUtRBQph00/8evF+WMnrNB2jr3
DA5oSbQ4e8C9Lj5nyhWuYXnnA3hJSFywwmXWBIpmIHZ7k30ZAuNpxp8+K3/Y7y6a
8KK0JYkq61pOeooQty+vjIytM48dgd+P2Fh/1cuDmK5yc/+AbGuFTeWQCCEhfvcX
CnRHKd3WzTPr9/JDWyKUuHlZLp3PYxTNazvZixaDOIjsbwmYBDnMwiMxjyOd788v
mJlMCTmKJ+dsuL2K/h0yQoeRkjsjZWr3c5h2YtGevK0dXsRVxB3onHZE3OVZ7sbM
FPLOC91vwkqjhpudYaI6PLq610anpUmjcis7AuDnF66p/5WkXsE50Szkg5lA7V9n
TsXJFoNfSaVa4UdP9W60hWeU/wRAtQigLbDAANa83uKppdgvO6T7QRevmmsjIR9Z
CfvDrumECpmineDjjMS98hTXiGe6k1f7+opG9oHQTnAJP0M0qJM+Wz6GMZDn0qxV
uxfAz1xavhrCHd9FV4tlYkef7Li3CM1+iXs/LK+/twHAtcSoVpnudbjCSYMAO4Su
jcAnEf27jMSsyU3ae8boPCa1n4MqsLkTZvpEmY4AzdGzobH2lx+4M0a/rSY+hLq6
O9NwhEBut9RnKhScxUucAmpHorLhVMnlJq3GDmDUz5o7Z13ctFhFNKnoM6qlge0K
JHB5Rmu+pfyF2Z9h2ydJKxanYpZCpQRjHNp2VkWMF6VApfZARRg7ydlUw7CIS061
uiP9D1pGiepz9pvbGlQ2ndbDKWAl+GhQ5iMv2S5JjHhPwM+pdwXBko2xncmDfEKd
8M47ujMwC6UfxXjzL+vCjQRN7Girpfb/ya3vXFJ4emlOScC6HlgAXUd2GbL+cdvx
k+w7XtxeSlYVZNiMSkHOwpSGgrLVK5rvKX2dfX5nbTevfRTh7OqflDjPnQKNbi0z
xMA4Or2rDVu64uXLEvt12f/EeoCih5sFWF1kN/mAjLjC8SZjr8+D1q/c7pth2Atd
hvMdtP3irdlIFBHeO+HP50qjBdmSyrdnMoMOyTXV+bon8BTmg0/etbijeuggG0xO
wDHK/1DJ9iKY1KVgGkWOQCB2N2snMAHdboMTzDwETOFNZUggw95F0ZUfp+kwUyKo
zelSnpH6U3UCaxtlr7ANbtitiBz8jd2ZJGFx2VRqLPh0KwlZx0Er7ckdvsx5pOm8
6odx7gq67Gnj/ZzzEtwGl02Nk3qgipjc+Zx93rdKe4H23uGW7ZSQS3ZqZYA9wipB
hV6cu7ipRUpatznlmqA525mzIG6D+VF1E4uveshxIOEABVkewormlX7uQEsS15NF
6JwFXknvIxcJ7lYe0Igx5JXsTFek2/esG/vH2eAghgI5z9JJZSqMN4eaPOy3PLom
W6usP3VNXSi7+6/xyImk/+8G41MWSMw2pvcVxqF86D3ODKFxgVSUaII/s1pD/78a
S7nJTRDI7ol1JVxP+eBHTkiKHeHPG0JYOQkHf3RJA9pw4C7n5nPMUYXNz5YBFDD2
YwbjM8J34yugeuKnvSlO8rsjdEL7JU4Do2TLIMaH/etd1ursrCosREM6hn+Smj9r
NmqDONfjxB89VOvw+SWAdB4UE1iLzfRrFbWbujlNNBr0tAPS1veFEOagNMvXnVX1
U+CwR9tFLFelVqz2rkOyqhYdkE4d+RTQvLbDY1zUmcp058WOlwCqvIDlNQzxhEfp
tFx7JfXeB47Ds/4SBOeDhpDT3cWJi+3gJlWrAuKCWCoTQ4UTEzH4vPhk0BM0dCmS
krp0/gIliDXrJnmWJGZ+CBYuLlvsJQibIqwj4OK5KfVJzPm+SeVzDhrYrwteu/l2
AYQ14JPrbz/osgh+mtu73VC3dym1cp9i7CyZ95HEPy8cA3p3y2+w8JbSl5uXG6iI
r4MvBgvBRWaOYA8Uz9ajkULdVgbYQcdJxHb+hX8S1Oo+Mn00pa8bYnOOUe6/WVjG
xHMtasIo2bgy40bREP8W1dh4SGKGYGKpyRiJpdjs5oCL9PkdZqhmtd05c4xkQEbJ
uK8sTFBA9NixbhfM2+xeTwJ6syPjAfJnIoa+Vdl3Cu13B5gXV+Wu8gavyV6UAQRn
ywlocVmpfWMHx5KQ9AYknMoTU+hLpq8/vdpqogc0wAjSSAZETOZDdNGFRaUbOPJN
4m6H2aFuJkR8FfMQyeDpVD6NM4y16aclUF6uWGz8QV6d8EiImITG/zbUSiFcVtvZ
TyGq97vM7XAmXBd9YWz/0jKaa5a3x0FFeZxaie7adKuvlkU2sUKmWjXv0p/9FXVd
jxseyWHWBb96dldhH1VB+LSFulcvPR0sn3z9F+FvypNHNdd4QhPLJRrc06DvTOCY
tJATdCkSmQN1NlH6Qo4a5Oux0HMYkqSAgmtejSs40OAdoNoM1PhpVMH/ZoxIZJJm
Pt2nlKWeLcNnhrmj3b+Is79AwEO7ib99ALRw3kUONzqUh3yHIhveJoc6qSO9OOpN
fu0DGbZ1PqGbek663Bd/BAurZIrWz4X8qnoZMxFW1cJke4eQ1wpb8nyzB5Fu/SpD
DbpsAbisaYqpPK8bfO71mYW9kjBkTQcpnAtMrShH/tRhezK2xGLIzXffUFtO6Z7m
iSZcRc6uQw1zRNIEyNFcA61Gh/b+muCH4Tdy+8vO6tv9+IVeYPtQG4lKRMddIv2d
+rxKUdFLMmXWndAi4bpGBjlSi6cZYz26QKSuZGnCXdDkXhvk5lM/LghJq26UPMqG
i/ko6uhcweXMQeyuJbzunICUEamtNCsQjPAB6+t6/QoWgJbcjouAUx9Ua6EYtmHw
HIkBlTKyBKkpUnS+Yf8EsrLKOSud0N3gJTnZkRSRKZZwzU8bcHaeb6oa+lz1jiw5
HMrvfSCZl3MWYCcRGUe4OLC/nzJPR6xeNFWq2B6J3eRY9u6/tjoEQVh157+W2BEz
88srqH1tMz6WaHKxB3i/5OCdc613bT/NL8H2r0B983QXXZFExiFhYQh/yodnVzbS
6FuZqiulG9uz+DnRd2otqLgI+brwBAOfmtTb59DRuOOgapXwj1HwPhs2DAnnuBm0
hzTic878n7PgoRpxxi4wShg0oTBcwN0vPQQjNjoktAEbUp8UZzshGoiBuFU0UfRf
bNc8uXoQnobWS8GhxYMVARqcF3Av6+qNZkLAPrIpzjaTvbs8LJ4IKYJz8DJ4QWbz
I4UaIt5Axd9oLvD9m92Yw/XvHbju+emRRcTzRYDYV6ttKFWqVqj9Ec0IwA/IGyKO
+Nkeo4wx/kJ58J3+jGCzwd1QHLZhxGCMzBT05IChFcEhqR2BZjg7X3wpQnos+8FQ
oIxK2WwENbiOZuMZpJi1zi8xx5bXgMd8BEq6PwcrgxD3PLB3GSCToU6ZTjWmfa5v
Dt8WvrGTfWG+eBiNyyNnDesk91s/xMrm33O72zGTHHC9a71ckzABofRF+SbmKRVA
WR0b2R5ysIyN9CG7BCb+6kwbuKBAV4BNKRcrZCXGiMxTIEtNxCX4COTW9wXAF+wu
ItH+1W/SMEf1F9iIm1Yc5JRyh5HVbVvSNc6AdMhiYzdXQrxfy1UmfhInFLtykEZ0
/2CjFNTHGHvjxu9M19jqjsqfXD0+OyLvzR/FkQxi2MxZC5W0PTIS1aZD0PSXj+ZM
Xl5SawCttSaaW4+fO3/FZ/U4W3wDNCl4Qs7z0nPCrfVSbLFVnC4meunE6Ub3wRj1
h59gTJrVZn92glrXMXpcGlqUs4tGtVXePNJVGH7HOncH+rbihxrTA9XYNbJQQCom
xtlT4ngDFkTfUqEcaktNOMBRqbDPlthvRph1XZTpaytCYHQN7vLl9cUygO22amHQ
6Hc7WhLEwbxPLdOAsxbPWb0Bam1GcuBUhMgy33SZgd9OXgwzr+0GOgGtigNNcSJ8
E+rt3vHGOrBFYGYPuWFr0yEYojNBUCM1nAhPsgpsUYZ3ooPrNg71ZIPyYds0SYUH
J2tdjuQXvvXdFmDENJ567bYr/OeXqM3yuOaR3JPlBj2ETXJE4F+vk43vQcczoPQn
GwejkidhccCWe/QNeH5b5g371UgWQQLp3cCb28Voe7c5mSmamSuq1nizlKU3OEF3
c7O7PZvb+WiOgDUaiNmH6FJsknt1qgCR8LbbDdQYxXpn8ynqV1uEj80Ahk7sfvDt
ue9bqyXET2hnLWmgQ4ek1z6boNfUcUk4DuXesJavKNWRNGCrFLQWF8ksb0Q7cS4M
KtdGa2tYEEbF/gte+h3+S/OfoAlHiobSiKdviRmu7u0NpqaPuOcIZYscAyg6pYNh
TbC7+1UzO6guiOZmLGrL7EcBYN7opTJkMV16EkzSx67nRQHSUGcVsAojBNXuoWDE
32i7o82a1KhgfJZFLCRpEmKX+JsJVCWaQckYKn5/Bh6SeEAAL3OYnnWaUUx4gu9i
o9QF7mLgfVyurv8YWJTxvIguqI1LYkDF5Rui+v4XVVIJKjHnU0qm8Nk0hoBD2BcV
MqoZZClXrWGuhDuca+YSoB2A50UmwiEPrK6ocbcMC1BeR8FxZfP99w4a2H0a5bzL
Am74p6DWzwzcxs6WBHHHvfAVZRb2koa++SDrVXSThlAEtHVfjOczaDBTJvuKOqM9
MFzZnbppfirUdCdd9biWGftTXsSEIASsChWROps775Fpq2kGpuyRKjl02bfR6MKY
5mZ1lqlOiGd7FK3GGot9/qmVyqNrE6XFRdKWjEMwwFH2ahCnDjbsc/npWXAwgbD0
TVDe15gVVLUnWpVdJSjLObtfHAsHFawnhpIwtI3KPOnhVj7PKUFFEZLotSxPeAQA
Un8yYf0h9x1ryTM5emj+ewqfefdfpJUclVeg3V9QculnEegwFR2diVah5z7O+dO3
8JEjxyOloy3BR49i9IEIxJZIReTRHFjSFHf8+NmmbTmL+jrsgShzs9klS7chnHkp
fo0FbYJdBWFTqO5MnPJaRljcn8S8SlqaJWHePvjt37mod9ZWyYYD6trvE5Y5sTaR
RAqFZLpKZZCyF5pRH7JhXZXSv9wLTllruu5AI73yYouHVcXHx1oZockW0m1v6bDi
lTVqBCSTIo+YuDq4U8eviMU0tbgBwAEN+qvENnq6nx0k3UG6DYtuIBQmua+THCtU
SapUJOQwoSGK6UKxkSBLVNco/ae7gbIGMhuQZuov6XVa9gcrt1e1gGZmFmUAlFjU
modoXHCZqSSEAjmZ/Tg3Fmr30q89bA0haFusdKTIUDf9uaEz71YmTnYESTLGAy3c
qkSQiOGoNxZcWtW8lXQ1IOIFobCCKIFRgTQLssJorHXGXwIhybld4kkcuR9vsNzs
Rol3awaX5O2uNfTzltmFJ6ClylrQ/eNF8ZMEPZflXA36MC0sNQQZGFVawLzhdgA1
gY80bbfEuPgkE+Qms/pOtbgJbJNvGV25fyEEh86VQEFLuCDrxI03Z3mUEwsc3Q/P
Ofk7cnRVp7dAY+hVI38t3BncFg+9IGFk2mG0m/ZuwpdCoG/nztv9zil6z4vLlhHp
MXbSSBRtPKDsqcwH+gIGo2X6FMuT9RKaiEvKP7eWqCLU0spyZ8yQBA2byOok6GP5
bWXo8jv7EyD//MViWrtKVqP/QFD9X5KPUEzwpOVH5Uq1NVqKuDNrQ+5myaD/cgCB
VYHvWbUKxuf1+UPhsdw6tSMEnG7y78Guic3YYNwTUgLwpXOQPRGV9ptbeAfgtkaU
LG7Z2qqlX5hVMViTKi3Ie65qVax5APTsYjFDaL8tC3d2yf/zF8NKlRAaubaRfPIZ
hubSqU2Yibh5VwPJwMp3+jrtACzU+ceg4Q3RLZ5yXx6nS1JFo501CrC475X0JrWZ
WvCFmd+22fQvO+eXVb6nyPL5xIl4LrTblZF/Pe2I6XBcJ0htA8sIZBWUaWhfXiZZ
0epw1kzXTrjDR6j1ggjF0TtKhRJjkJ49QOajmG8RwuJfU8/12esUxs0qRku8W+hf
FtdYhWRbldw4gCt1VBUC86UnwHDQcsXJBhQdy7NUNzckwMi/JUV2F+i2kIlTPRH1
6baubeYccq+SB68VG6gW8SrtWYJEd7LUVn0TJfsruBnATbogbWHDGL8LYtlA0WYK
qmaS+43YIpM0ldcBQincViRB1gnusrHQeKsjOyNTd1f2T9SoKzHWErVzidqBVp0Q
Ywpn/7I/RhK6ZFoY+Fk70iDNEwlTfMiNYSWmqQ7n0GqTKigQCRzWLW/TNOnfR/uk
Hs1hvXLUAAvwPelI4QywZ76KBcRKUvhnG3saRL6TBzg03ZXg6b5b8Y+RDvatQqAl
aY00/WkF3bkGQC/2E59HR2OqdsTPGoPWl9Im5bNQ4wRPyfnEYmVtdZyZSGwXP9D6
SjOP4tfFAFX5ntYj88YWYJtk8ORyDIMQFSGkUFaxzdPIx7Splvl/IIKgMrMC6+mA
b5eZbf+nXNeMAIwDrjaNaYPIzls0QCl8h4PvWSOLRy3gzwDvo4lnjdKOoVmGrBrN
lnj6bKZ7rPGIzUIUcm198BnPPXJRneBVtWj8NPla7q6Zf8AGhqKzvQy2yjbBDNsC
P7Ty+VVITG5nGP05GkJuFtJprrfqi5/tV6wM6ePYtSTfOdfJSQxV+ULD1/fxY4Vt
+caRcqEyMKactl7JccCqM+og5jIN9Y6bEuECQBuLmjwChE0XeWo3/y95SuhI7JRf
BUdSteJkvFe2kZVlVCz6KIDumF+wLbkGZHYRyVosvuIC/AOnjkJonEztvfFFJq3p
+yBQWgkkVqXIc0+TiSW0/Q/o8z2vUfAIFBchoBZdaGrbh93ky5Co4iYoNWw+M2xx
pekqy80vPLVaWKZP1kJd0SOAwQZgqehVshQjMeP37gufGQYX440U2RQJbw20BRxf
U8TAi8E13g/8BRYcihH/s32uJCyoyFGdXUhKTqB1DV6N/uzHYFpnouXG0RiBJryL
PF/uWYvKnlLNiYY4ELWaEqSA8l7Fnb5jDC9mfK5pBIL9qja1ywIwGZEV3Te07IDL
JDyzAengPDpqYT5+jYs86aiwl9HVLZluBzV42T3jG3fV0E/gY3TOkzWWpEBk6Uuq
13QZpzv+wsEvE6fiTSPfy74qDk0+iJhiArmWlzoe7I+E4hzoEb/Ry8jRCtyxc/9L
E6k8wkEZ10h5AZB/PS1I8EiLmK2aZRnSZMw6PxBgxsG6IgpCnft9tSFLVXwPANTg
kiSNgIh16KTLzAS/DM5j354kEPfUN24rRpckyctF4IB0P3MXwVXelLOMtaVbkE+T
UoTZNh1yK448gxFconcbjfQwv4E6lQm3Z8cCtQSyqTJaNNdYIMUjvZyUFcXaWYaF
Tnl7tQnG0xR2CblnFRq9vNYjfL4LSz0Spju9i4rI5Tpx6GVAjJCChVt7EJENtFXt
HGpSl4fgToIIGLkkA5TERLwD9msWr6i40RYjt9Onm3Ej5Rd/ozRb7zEIqJEojvcO
crn+ZJkR1PKhhoLnvJ67WC+VbfMKK0eO9c40KK36ly14hNXBRxigp8JPEyNQA5eU
4qvGJtGsyZGVO2AyUzAFBrdXsh0+U8CymGf8QHE7WuevKQLna1VhzLX+T0cd9HLI
I4pPaujW8in3tqnB459mETUPqqikducpWC8wljEieneKwV8kffjtxvr6x+QrrOEL
eYKE5bisRrlGaHQk/mEWB5U5gpm/AMpWOyYwKgeHMPbxo0s7Qp57gGakBYVwKSQy
zdshO5MNGVDjt0XABrpey85paLhftzq0CP5CEVUEhJAl416KkeFArVv/Mf/XtL4D
XjkCNbAXHYtPT/uIzPodEIRdDX+PwpzaQ/8kfNKqoTah/9xkDMF5begKeJUvmkmw
Qljl8iLlaW+rMZUQ9aaJukVqrc6YbzLICWf8mueDp885SU4EAB3JKveMJDbbVGx4
FaZyykAGpnKcsBa2G3f2dnAiKfgh6n3kBvyTSIE9EbbydWRyQB4FKNwud0rrF0Vz
vzAwp5bs6sCtvMiGcrOA3RGIoJRukehiyal/zyz0OK8+ECHzVz2l+IejFj5Kq5r+
45isjb2fuKBTD9UscJLW1QXGUpqrZpPIjuUXJ60QrPqRTj5hOtAZCLTMfzK81Oat
Y6feOr/o9bHvrDTF8XX9XoYThjKfysuspJ5Z0pAB/tJoQHbsKt7z/X2LZvQrlO9o
6QHo8t8vkcTsm/ECfHq+Yp5F5B9kHLqNpkpW+i1e0tncQxHgpdIHdEsW9+HXc9T9
lKIcIktdvJCQo44zlyCKEbiLm3pfGqqupsTzOPJKCw9a6w595dBuHdV48RIo2I6j
DjrZomcSx9Z4jK/fwwGEKWpg8/r7Q3AojdrkF76KZ8Z7z+/Ek3t6BlupQzpCq8TG
QNUKsNiEIBpUltPGUnktv/LAY6USiUIusWDC/Vhnt6D/tVhW6XNCbKt1ZI8TEcjd
ZFtrzDyO1VSuVGDHxPMr+JiXu6tJp20baBXXG3K4J9YyaN3Kxv+YheIRGSaBT7bN
X8LWUxRGEMp/hsh5avV16GUixvZiGfgN64rwApPbPtfIeuoHNs7LyA6EhvEur7SJ
NDEQDu7H4gjw66BQNoPeNMyzabyAIIevlFJ2V3XnnS6xvzWje0uCssnKi/gAjoLF
KR9ShYkquO1Dbu075vxpKuPHRUX1P7OqvPg3TNLkU8Q/1k/zSEZN4hwgShxrl+Nn
iZEazTk95nIQWZjLaeFVltt9SQx05h4DhFsItBOnPbEMJzanp2H8yUVdIxZZ+tCk
Ge4E10jh8y21k7JsTcnyD6a0Dgpl6CKJqPMtbD2g51RMTCLcFJ5GXfSO1yqlIrCe
d3+5SRdYb1+1gDcZkq93KinanINDIgnDE4kDi4zWaVWTn9RzToghphYrwZ9guLkp
FuTqMaV+rwZw3OuPV+/3LIsexGcN0w+H8B8BGiWiDDUmjskmDeXNBIgwLM4T0VIv
1KXhbfNq/zlCQar5TWAfds39+22m+qLjQhKOOa7KlscMgFm2SSX2mUbbmoZQHdtq
AXrqIT+Sej3mkT/yEa9Klrv0krsQp8bM9uhASl9J0OWngP96HTww0OCDsnaY3Sll
JCTbbxrFQOBSj8Z2e956AL1hiA0e0N7WWGr3XEvaPumo5itOMcABP/wMNE2L47nt
H69jUL0YYNJ0eai9t54lAdNPzbv8QQwr4grXkytHvUh/FWhjHy3IIi73a60CtQh3
1ZcjkwiN1Hql7Oam1Hes7YejRZfBsjnPg8XnOPm08E8Dw49HFxrhzS32XL7O2uUr
8WQ0iNoY2mZOKujg2fbDuhexPt5rPPF01yzxAmGKhTsalp5SVpxA1dXJ1YjgWmzB
LQWiM7ABur4vpJtB6pIRBCEg5nWQh08KDBXdbrQuxrlsvuc+oPJV0c/RTPMRGzf0
GfPj0W3zYP8Hsf4VCgemV06AYTp/0UySnFhU6pU5CWebuxx37atK8ijcLb7DRx6w
UJC6QLSXifW4sc7SFQzUXlSyaZ/IX2fR3tm8YlKITxFPs0a3HJnUADH0GoQAYICF
SiRcyrqQ/TzsM83hgX+iwaR3c0aJ2v4GevhHBPwGueypah1sa/pylhJrygMx4ibz
5G7Gs3gTZ+nIAPvagojTm2ZuPZwjbbKICSCihP9mA0f6scMcjreCUdNkhHvzs3my
h7msQ4DnWcavA8BGoZY6cI0uUL7Jdii2AOGv9SPT+ipjtjnonE9VfYZ4nUkLQMIJ
rj+hRnKrmidohAi0U7rZEP8qNwZh34V0WZHybW8jvrYSwjrlwg+DCplKTtvSIE4p
CjTgGRvPkQ+j13kjB3vX5XLSyvQjnJbXIQzIxVU6ryTwyJJ0P5qMcDVfKLM4xki3
NxKdoN+/952iUt1jLCUcNsawbZGozuj429aniMF6kQ67o+yCw0FwBEUZIR8KHI61
wHtqlbtxtEUVT0HJhT92TIkj87pb31VS29K41XN5xmtG3fEXbtysRFXyZK1ugmZB
O6YoQD7VFGZjkPANw7HHW9jWtWtLhi8RarSf/ec3Mrk4ovk+6LUF//fN57zWHagU
0Xg0AfNmfR6QF+p47KhrZstsOaxfY1pKxrJ4QO3obQJW7CjHSvpts6ajjwiO9o3S
GIsK30Jgmx9kWWBIJubcjRUPSBrEePbU0/g4RiP74CbwgMY2ZCyt5rssE3E0oYFZ
XJn2Yr6Jl2vf51RAM463mJQoIdYE4ur8Yiiy9KwMa3O4qOPl8zoFaNtROFpn3NCB
+fWgFs2MiUg7coItyS9KHP7Y+egfr53aBH4x8jmivMbmLth8AvZm/WKrjVPHH2FR
NkQOaZkietnDzWLbBrlj6h5RuzTjChR81+imje6VO5tfqZS2q2lIA5xtivVzPHeA
p197aqAXxoLzx/DF/QsobEFFmefnrl+NzErnY9BdjpqX10WkAJ0m1NwKEJbTMqfz
8VhqWy0hGqdBs5m2fgyT09lnTg6jOH70ORKpBCLtjHW9QlSXEtx0g+hi9P0q09tl
FoMpxpkJ5lIrljGeYk+2P6tWXo+FZGKtH7PsG4JPX/O9WWNeMvXO4McJo70I/JNN
n2L1wBKKgW38h+qu/ohLJv3xhJtrKjS5Cb5zsObMeBeX2fZOMErNmsJlh4uGLbYR
4Uv3oUk1FtwLT/8gSU+LHxiRdA/h1vhftQpqXuJdsqpvCHZmYa6E40d6pmOrivmB
K2d/rSpiVXS28twCAI3yGcFdvZgdYzEsAxpd0kO0lk74bHe7orbrGmzVoQxcqsgP
Epidi1xLfmaNRzpHu2II4kGCzwxq1Pssx3UvSVVJFNaGHciimfRuiP+vplYQOFzG
mLBGGh/rOnKh5yfLikk0SRW8cAl2pAJtaZc51chkTRmpjhwHieHGrgQZnFlIcf3F
QsPI8A6Zt5oZaUu8a/KGMF1kKWNWuaOqyCnj13l+uIWursxSs5/qpHc8wEsXfnm3
PJ7dEck7Rof1lKdnKIfdy9ZqL3IQIH15TRId5gYcCxAxxkj5SgNrU88GGpzD6CgP
D/7Y+MG6lvIWU9LitF1qDL8S0G7PxtTSOWOmdlcxv4qIDwfqgxEozkZ2ZqTcjLNS
CnAWkE0SGe0rcJ0km8Uo3sEoD/vfypcfebfxJqtNG7TerbXzWcev5Ajun8uGBkVl
Q3dUDaCJeltQmZ4O9mG2DLaARUiBiheIratZufM4+Q8vaO1HDkwsFwVX2Mf4LeCP
nZa02FgXD0NwW9ZqzNHxuZtMfKgTql5hOvcNkyE4+IHY2XVsg2HBRVvs+iL9EDAC
n6pzI5PekDoYG69TFi9sVAriLclo0PrQanLUjSD4YHPKCyj4MfpUp8YgnzpDWok5
GhsN9Q8AJ7Y+TxUEuKeVMLzJzWtuGkv5YDY9fsx4VsSFSd6pvbwKkdBE/xFuTAe1
9ylWWPwZ2m5yxx5udFKDS6TE/26n7dtW+b9KuH/CcSVcUxhQqrtLXTf2G2vaeuva
SPddjKEmS91fn78xtIbP4ryo36y4YvLTApfwudBH6keM3/u85VHRpJXHnrdFdezy
Ps8LREPfPoaWdlHqZDoqAKhYxBfHjSCpYoTs9+mTQcoWpVbp2CEVP8OIjmatdkNW
h3QSVb/K88kCOeDnhSUNNaqe4SmclkfvDmvAKqlNauYFYK0h7zbSKQU/Bigt7xL/
8mVtUpPe7aNuBM8E0nuCTPHNUhzPELx+lzGJYe0+fdPJn/6xB67vtyB11E5Xm4KJ
K0HyT6tLhfYXdkuvg09N+ElqTlTnJzYEYvORHrpZAnypkfYzVq2iT30kE20w30HW
PEV8jJSOe3LOQFFuFslCAMGVIT6LTl3OLIasLSa287dgpSD62TmToS9ze0C7/HwM
pMwVbWHYWrdhL7kZV5hF3tnCHvUwVUon2luOq6w4za+pL1AKvNcGB+B1ptmIVxKb
lr8qAsySI05rXZAJZkawlGjHrJYZjX2T/pOzxB7w172jmGVO9A2aCK9sqsG+YUs1
WkSGAOUm8iiNNNhngc7VgNCoUmVpwUNgxRKy6Zi209cb/wgBmOK940WzAQQaWnyz
G2inpmVm0oZ1fFinL8xXd5Nz2SFSI6tgWx6IfZcvBsj6bCewVJm21uXAZ7oSK1ao
dyIdenh8bYxP0MCLxFirHHCZqppEND5WNvxAct2Anc8pqI0U4KnSyYN2Hv1bC3wE
htXVr12rlekTgl+IutHAUzjlY0ay/SwIx9r/umwyvBVmVQplcRYEJB1ftwd5pzO9
Yz/p3xv4e0gU4PhDf1p2RMiv/JsI82veeng2hNzx21yP6uhYvv5C4JUGGD7CJJr5
pXRGiABxOd3HK49nOi4PsR/tE9rrC0ZZMbEImVnCIS+xeTGd4HMeDXr/Rxog0e/7
n7v+xq7TPh+AdgDXM3vARanI4Lhvux5YmePoKyEfurMC3xUFW4nRZCZAuPcwADQ0
nE1bc0TnkNdoALwrhf/bCrGBw9tCHQOC9Dw825tXBqbnBI3dYA4eW+pqbWz22wQX
jbtsFHG2fXxYurh9vH/VK61MHsjlXgiybge00cjKAhM8JhK7+cxIGuK9wzJwyZjy
bR3cBzwKvi8OU/u6IU3MW4mqPSNoucTYPvCcHpxdUrOl0NCxK7r7AZqUxroYSzVK
i9LTbYJ+W1JdWbWVL1WirzgFQFw04Wfc9l7htdBSXOsB8QMpjP5uX/Yzz6VTr1vJ
cvO89JaG0LXM4+hPjgnJ1+8hiYoKfn+NzgjN1YRxTjIWsh2B8GY/F/+cOxluopyO
KPMwOx9Bq8BvpvTS87nAqwtP4+kJgNeK9tUx1t+0tmn3panJyeoroGBnSRD6RRkb
dymj+nAjGjf3AS3KzoRmA2GpNmUaX4fQjpv11jJ1RSnwVxAzb06roak71AicL7X4
sk4yNmA22FmsAORTTNlfHdw+yzU6nUQVlY0Hr8+k0vqOlgwvI1kHHE3Pqznk0Uas
ll3mx0Z1b1V/UkoYoB9jkr3l1i1ipwfgXIBr9F0tBsx5H1hl7oZYxIuEK92XyP86
4JpDOBa2CPlCdqJVmQdTGVN+BCgRa1Y6ZmjwSjJ8Sxm4/bhdoX1Zbkv31pWPof1d
3SAi09nmcwmwc/cIBvLPVYmCjlicKKEbHuqpKO8mw9NwceXhV8f1YLpvaYHxIeU4
y3t9z9Q6/vZ6M/EyD9AJou/RZxuPV4c8A46ohAv0ipWOUIbDMbV+cAlFwvWL7UhY
KRu/hKSkO/BLIT+GsCh7Ilbdv756f/pCgldOcT7mrjyzpIQJUo3hWfd4vWk04Co8
GrlVNZWzKxXbGUW/NI9pv3EN7eA+KfCe9ZWcGYFanA7KyQiYz7IJIR1PTv1TlNVP
zjWe3sEagbK5c67FmWqT8R9mXTveQEjYdljOYJ0nXAPTO8iN3uCiprt+VMki8eFb
D5L3LRnl9DSdpGSPw89nk7Sl5JYEYrTfy6/wFuuVD0mmbkJ6p5o0Wy6Njd1SFojn
RMAp3PuEsI44GQbIrw/K+NffWP1q38EQiKbZKzyDJSQAR4Es+S8jn9ZXP9XTfdCl
IcGMaz3Za0JgiAFLC3qiHQIJicCJNdDAgPWqLXuV5D9rIrz5b6KOlTkw5cfMYPsx
moh1YYBhmXU34MIjwasCMa/4rhLbOvFnsw7ByO8Qm2S0P5Rl90wykiSS7X7DHozj
qqF6jDhGR6zldSuxcHHejI8Vql/kaJArDhbdbCiqkCp+lav2T1GCSv2ccbk/D2nu
vDwm/D6MsI/sOrBzdk9PVR8gbw3a46EoSJMEEvCFfZhHGuSTpGYAchJHCoXCvsIO
tQfveJ4z6CoNJWuPod31+/qa5q21w/+kM/kuktYSMr8DPbR94Ik0R/LTe5pqgnA0
kmj50AT3A4zIzqq8PB2T9MZuP0bsFg4rBOUuxr22iK8kqxN1cSAjdRmCkdu3docI
2S35pvaBHNFfYCfjWR8IQvLwanxn6MsHpWIzbjLmwySmLC17N3ciLwyw56aUjnag
TXGEqq7satDZTrcxr8WTFAJoU3ncoKQzDCW8du3U+4WMbLwCPBxPLgWS6VN8nsGN
3Q/MarF2nMRz+RXSScA41DjIY33JEuAoV/Ra00nrOcYZ0Jl7jeCiFsc3V8T2WFhF
P7LS30IuXeiO+oS2kh0vdgRm0WIlDdZWU3ZYEQBmRqs1gnhKFwbjRmBiTCB8gF/4
WYKd2OAgmA0oLy9+nwie+wpCJKClDyIG7hYFEPyLMkOjQATH29IMi/zXXRDpjI/M
C95NRpjM1F3mtNbV12vog4Uq7evGxcr5W0i2SatCSe8yAl+WtwXsGZJ6eugpRpcc
3SThsroGy8JxTGOfWUeXok7byd2tSqdQtu0YUV/mNGyuggRMGnM7fHVrVw7Gbe+f
3XghLNVjez6YqfZBFcsg4UtRrSGGA+k8+IFbBq8Uf+g7xAsgGrelrA7cZS/cAQF6
A/dHfcLlpyH8WViSbE86A6MSVSUULSgigilH59LfhMd/qeHJvDSfIUAjUNsufcP3
YXMfF9poltVaW2lTpEhcGBPMIErTxwH+c3Re9Bx1y3UtRDvASpPWlqKvv3soezaF
0rkymFjLL6PsCFrPyw+cElG3qjwAvwocwuOoCO98duUPLld2litoCe9cQRZexvax
Hb9BfxDBzgeO7ZTQwHFbs1CLo/eDAt8Ju4puCJmbJ2jnnrwbEIAIHzTRsc/sb8Td
9U1Xq7I3ZWdc+cvHQRbQcos3plQNsdPbz/Ab7wVAwDd2S3U6S2sV2X07LmLoqiu4
MGcvTQoq0X62s273++6YOrEnwMLvIVIVjXwcsp/JQfV6teXEXKt250HbPSC4zPL0
Ca7iRuAZ93HXIMOQNZnmxx3Bx74QLPJ+5WKbwbCN1X+mJnemlWfOGkwZ6XwR9eVo
4zaIbb8EwxdVz9WgXhfpapcbJZG2qb9GpCUu1Tvh6nDWqH9XJnmzkumSDisraz45
QfrYVLcf5t01iiysrWNtOlbrc/3pLa1BMhe9ZI8ZwqnXNwm5AXGFhthiXww/Drst
aD4AvtNkQJE1l7pScZf59jHGnnp0NBysouOdGzVyYURpXJvJUF0B02C3Z73AkFVE
9kJ7xaiRPw0ViL1iBbnn8SfSEhEaEimArcuRXcd4FzUtbzA9oQDE0Jq7BzE3VQq/
ataAP6LIWLc7pOCaVy+UVZJlLDbka+kKstUT0s+xSGtOfu30W4a9Wo17jXtn0ESg
5HKtXPEDwm8FhfenpQ4TJbanYyw2Z1MwAxR/YmnSWdzP5PTX5LdtxWae5hOIO3Ba
W0a2bgldUFs3Q8tfS9jLc+DRIouSQqgvOl3oC2m47aljjzLhAVx7VDFK0uwA7hNi
Zvi5tqFinxbjXmQ4+mXTouuDVJfqeOFgNdpITmSy2bvGoZ2dTP41L/b+wEtc8Q6n
4MA7srVARKNJcCss1lHIjM7NGnFjyTLNX5B9gCcEf3GtUltCM2l0cvSO3q9prpqS
WXNGzaHehD58XBAkeLRF4Lw1hB1F5NtNBD6fOAgLSCXejb2Lu07vx6sD8cmHzi8W
01T+YdT0TJXq3qRbd79m+/zCkafDkv3K1IqavT3g8Bq0ESFCyxnNijFX/6zBz2Zw
RH781JEswQvZTYRRWfxIpZZCO1PH3rtqWRTZ3Muuo0Om5m3AwW/MIgOJ1MkRi6D9
pqr53exr2Ve+EXGxxbobyZaL/wpQc9/GsduYSI2/zpaWFvBJogrtAi0vkJjX1mJH
ogiMrnwUMZlu90FD1z/5JyKRj0tpQ9dz70FkadEIACh8sQLnpHfxqG0LwRMbEyfu
GoK9WcEeX+4vkZ2tow0jgeWpB31U/MDz5imoSexY5HNBAPCxzx0NOJIsD6tzolu0
XpMx77qAHZAQ5W5IWy5MiYId1kuRaiq95Yh0O7vO4eWT2wM7xOv+OrfyXQPYqtF+
jnt018jG4ozKLvJ904m8eMfkgSbhA0aydRIJ8QirCVQMLJTMhgh7Qktj1RwaI7xd
eMwKc2zFgEGKwIEIP0bEgeRXQ7MFTW1bwOur32LRFWCI4npytF7D0SU2baBpqfIH
/YMa4FfoQy5oTk4RHzFN1QOpfHlUqOdlugZte+6XVtqym+n1mirs9VTsk+baRi7L
HV7qka+oArfM4tkjiwSvM6SD+RA9/61SaXa+/SF6kza3ch/DXaOkueqFgqGBbTWG
OwELd6RdVwDU7ddOX+I9zHLQdN8PcptYYjrM/3Zvy2pV+kSgUXpjaKJVsLjz0LFk
cCav6pf4ZK7ipUzAqERfMQ2e80I0ncpjaumGhlgKEr2US8IIVxf11F8vOkHmJU+K
3o68PRz5tHOCVaRKbEaiNO/RIwAnYdi2iQhn1buIZg+GGOPHSvCbmYRKUtK3Pu3m
vL/gpHiEu1PpXdXNgx1A4rmcUeBDiFR8CQgEHZ/dJ4ts2oH4Cl2Ttm9wOOqr/F18
d7x+55UCRzLvWmm5FdToQwOZzNXpICJfGIBfPODIZl9WgjfB3xTy3Q20IXsIntJ4
XQVNDI73LS5z7+xTJt0tDmkjyk+T6hpRh75VC3rtxr9MZuyGqmSxs6pLsSoetT8V
09E+uRRm2DZEJwAuUcnkm0KypKScSErlW5lhkmWAQ8CKkIcs2lCrd4uX467GmYjW
72dund/wzmvELDbV8hUMBXiiOhrA8O+wzY+w4WuqmPC/EZzLb8Bobtn5NfvvX6n2
Ldk94FsJS6u9Q1tZ9hNIaNTQMkKPiTGA8w7HjQs1zasxU4rCkz10Eeio3psjUIPb
yFIBblxHEjMzn63YNoK8vBPDaeocmnD6BLGakMj995HJvGRvrEO4VhNPbrTWjGhv
2hGJj0FsRIQdSaGM+awia3UakrEG18EhA5EXxkA254oR/yxGjxE1lxxD5PScfxv+
OmttWOp6742R+sMMtCzoh/Byfv81NH1rRL/zPGUXU1cQTBm6x/D/1GNnJ7GDQ/8G
lM6JZqFXFq/G9xRSOKzva0HBEHeDubeVXt6Mu/mExl4wBdvogmUl4s0RwgakuOLH
11RL5PEqUhkNoQuOui4dNiDHAq29rRKOxvhMkK3HIoO6AlI0px87ata4Gq5d0jpK
5dagbGk476t3jQc+FdtF8Mg4HnxbFFb4XwaNatKKGHDTlh2AqcsUtcMLM3HBlCp0
hBrLZgDeTT89yYn8+A7Qn95KctN2BRK2BTqgmIKiUAr18kOYl5nqH+phpYuEEksO
k/74Q2r/8YFM/FHc2hrUV8k66iqx243Y6f15xtLXMJD7BRlQGydvYa4caZP++M+U
RkoVIEpyZ0eJkldKJ/y4tE9Qt9RFYQ4G+1WrfQtbO45WWnQeU9EeTB6u5nMqakSD
KeFLkwqU2gdIvpNxWBjRhpVcSz/WjklfQ2wwXScpHiBBOrudp5WtWY2+CT6eOHv2
btvRDBuvaHR0UxDuucueQgFP/3E4lk44mwJWwOZMKblmSgO2zT2FAMb4MiixOH9y
uzf8Iatheu7DxAVvpb7pGoOvx/27TZyfhJhj3910Phq5Z7CoF5eOAjIshq7tnvZg
Bxhe3K5FQmGeegoB4dClmQuzVVs+nla+rQ9Kdq5KMASo6qxWxPkLgekDJt2ueWvK
4dWcfhd7Lj2V1I2OmyjaTrePR3LyHf6oAprthc+enHSLpPzs1ctHERcd69/lo90U
QZDiXmp6hLZeOfKSgCFyZ1tMNIhIbqi0+Ejny/je0FT+5hNBBNk3ugXsrsaQF+Hw
eB1hmCC15KrhwJgkwCkak9SC0W2EkqwK7pwHVyl3aIO6M2pZw1jOaoU22cpnyQf9
wVkgkp6f8LyFeHkZaSm6vBT97yFxzXepI+o8HVt6bzMvG/M25bn0uVKab/hrBXwX
38z9hMWd5xSJOtmGHKkrXR8h6H0MtgpJdAjLfmwTuN2L0/DrgWkV9WpV1d33J7E0
mRIewJr7huOs0EFyFiZRSBP7Qu43wFm6A2nyyjnv3Y0GSVWLhvSOLnJBNz7CrApX
gJDN1ZRB7cTn1fIFKkTZFOGkELi6E8sDgchE5uV/nEaE7xP8AjnJfy/nYnitT27Z
jf5LruBxbq4iO12+QjTInO2ackPPXHT1xoPvDPFdGI1nn1JCXtQljgrzZxAmsKlp
6dQ85yAkUEZK2xcdEGYeQwemUneDD/MMBIRVUBCyL9zBlig1Z18LAA9LKi0ScrkT
Uk9m8Ys3q1Z5Rim7myFShHFjxEX9npcMmt0ZWfb7kaTpGTINyJqfWRquZzdnHp2c
QpkIVDc+T3MfW2/UnZBAKFXr+RQ0rpOrPb8wSH00jblWclP4/kAkvLD1CvBrL3Wl
CQRpd/nOUKnQawQrLKzK8RT4xrJB9eYmcaJTckTJ8kuUaSJIdmkLHWsMTubjJN2O
BriTC4cuxPZELGkmxMHW3WwWM06RHOpvomz3I2K0qJp1V3byIsJ7ql20RKjqvSul
6bViuz/fSHex8hXZ1mPcL67+b/0ymfVMJFyqNCNn4Pte6nPoG8XqmllqQzh9K2d4
FjHiNQBh/qgLehCtqugZYEPaVg61apWYcEFpHAEiowp7pCOQI0HxM6peRTG2f5nc
GsOJc08JW/d6oMRHRPhK50gaD0yY3v7tkoj0MUfz9kofNWlO7O2xUUorXtLXHzeC
B9x2CXppV/NsOCz6Q3jL/sV2S0dzzpWiFMe6Oo0QjaL0okLn005JLw5ZnjmouX9Z
C3D2Cx9zAayy8MevVVj06fbIOD+FR+uilgggT8P3LN1TbKSXqKttmydujwZ/V4RI
EhXd+2J8TADodkXs6hSC3QogpJ5zcx6LL75cdyDFknYs4OEwLJDhb7xPATt53x6b
sKPp1zYbHFKYw2fGfgzCUqYDlT3bRCfMHkM7PfMZnd2dbf/xbHoe2KYtYbkdEhj6
4ysdIxa3MgIvUlAkrhJE91hbANIaocH1wveOyz6uNTrDjIRJYWUu5r12ogeyJ1XF
JujqZPT+6ccklEC0RjjTT7TIEplJ1bHw4XD7nYD61wz1Ml6f/rw/XrL8HrdKM0mR
CKYCRzssurSxe26P6ORDicxth8khiW5aPJinhekAQQxcqFmIpKEMyjsFmJHsXk15
1Dz96ruuASLnFbjRRgI8SoG6+FXMk6eXI6UhZEg2HlP7CPGN99+ZeWKgMatrx/yQ
rPIfuVbYtcAcZNBWfmoEdxlmFVPdc46YzcxUXFruhp7omfzWZq4C8w7XbrigIRcj
cDsOHleecgJBSTvrpkpCwqrFRNbKIYi+tEEJSD680ao09RT/o0UJCrfIMckHJh+z
mCob+vIGhKG1FBjzCn7m64+IDbDOsECNEXnJXezpHoDTKgBZv/Ni+m1hy70n2k5Z
J3y1aPqP8xxtToQLnfZr8kbo6UOyVefM3bQOSyzo5YJiF2D1VUkT5yn2DufJJqDe
K9fWjE3ytAMCXZ3y0khhhTckT+zIXQTOLwgQrZ5+tK/TnNq/Emqs9WQdM35y+6mr
CnTjQIgdo/5OtPUY0pkvxqbshOtkQA1CnTn668GS9SJPah4rY/PoIv0yke+7T2lZ
IDZT2TuOYe1qFt2Bqi/HWr6mY1LiJT6SF9NJo0M9mcKanKdvTNlcIxiJChdd5SCX
rwZz5dxM2gkixjTqjm6M1J79eYYlUFtcm5M9aUt3e2pD0C6oFSYxO0J///E7VO3l
xavQe3ABlihrSvsMtALb8mhHll/4jNU3T/ho/CG8PMXKf0eQav9/ELepr/04+aIV
hSfdaFA1WUmrrMK2eKGwrz+tiu3UqOl0WNMeL2JUwBqVqMtaLlP9+EYQ/hrBdu16
E0KNLcdN6ECV46L3X8zNIJlpmWrZ3K1qLUJPzjYYt1FecUQMN/lfCOTZBgkzzuBv
pRvn+bgphnlybSy3XxJJ+bvIAyMXqm2qr+F13mrKeYwGJCthRYKW8RBiBU6+/hK8
W7HrsvCmRKywdKhjCnnE9QymyaBo7h0/tUlRBvjPfbJnUa0p8kl4LzgHUEEwHoLq
zvAKqnl9n1PG7I1di/zRVfhVzjy9GI6L7hOUC/A+pr83W1Oelp/6bALhhrIDMEgg
e/w4YR9CbSCwgKQjLxVLv8I5HUJ1m1DVMF75ixez+1UMpfqiUtiM2ycFBYtGdXzC
v1lJ/650eoDbEcGrvIHdQbr6oHHN3qFkS/MEmyf9twV8/bkRzCnlIzf9sS2R/B3X
wN5cOVwzIXHQu3RSNEX/cvxI6xu7nWXMS96zRZ5q9+8pXFDGeJ16z3RpbonzjeHy
h6Ztuv8NpXgaobCYKKMS/G892SjPrFrY6skSdTtLq1kZxAcVfx79aOHWQWbZ4ujR
0mz0+Tfudzht7F07CSwOXMQxQBov/vFJoi3eJESKZ/slgi/+PP0l3Ab23+F9gtog
QJ0HOxwg9dS7492PbV5U+AZwCR7xVSrjrGRv2CliXPeowBQgeJhQXLrRUERimfr1
8azKxU7HD04XowulMLsSJeP0O5QAUy+lK0wHjHdgq23ZGMg1Pefz2ngynBa8XaUi
nNXnhDocp2Aqlm7qQE8Bb1tE0W66J7JuwfaGZj5mvYhiDcGG7KHqf9sGwRVXjqM5
yNzIJwLfB1UKo0K4A8y4aDesMR4fUf5Ix0AjVjqFE49zHI3BCLhX/2g6a0PGcOXX
HYE1CC78ysTAFLQLTyvr7OGa8yWk6hIBng7qjBikhR9oS1cgv3mSVrjPWegTqw0Q
xrRew7r0pBsnoK50ZiCEdMP+hTkyjdtDayT9C/6M71ea1WvOTkLzZkq3B8D9KyZY
Y8eU5sdRq6QXh+KO/8yKuSIeNQYJmTsTiykWZXSNGbz/q4Bh8TbZgehqeUBzEOBy
P7Ov3nrBKfo/3xKOJ1m0a6J8Qr4RsGQQmuGbF4E2+tyJSyesHbe8RrtqLNd0aiqY
Xe6mtSXkKM2w/+iVV5f0p/X5qxim408LiogT9+ABH8faPK6yVCUD0/juoioAn41Q
kcS2Hr10z9Ats1pruCOIzXxsyCe4eVHzqe8KNWNREpbiXUs5W504xWl4aPJ8iobT
XXZw6Mh0bicoRIlaUg6O8D+S05TnDAF/UOKiGRSEiM3kPxV5mupsYVrhS/wpGAno
jtCzfYYQNHcOwuMgFTFn5I0GKC0TSGlvJkWC6dNvEjORF0cBzE+QIUS4ZsCcHJns
gLBTFJ1R4GTueBZuUJddCFaUdQ7LObKfJ+v2Pyj30Ba7xLYIm/iy9GqB28kVxOAx
KVcBAGxqf/2KOWCZmQazrgLrsOhNwm/wuW7CsyS+hgSwmuPGDVoDGbr5frjlRJ6Y
KCksA5cPH6MYT9UXChV/J9ZnWgKStBnFlDRBuFAXHcu2CEL4gdaUNPQFr5WU6ATJ
mCGoWFRKUo+xePHHI88N4XHe+JK0aJdv2fAv/2Du7HlBPRfL4LtIpDBiquoYH8wc
ZaP4iY5T3YOo2R0OkeRHZJnFdKr+cXY3x9pnbrNvgVrfvfMeg8kBaHQUq/zfUXsA
LMgZ/QHcfCCxS56x6IFAionV7GXyWMAumw6xItp3P6PNwP3B1LC2tVeh7w1VgR/E
CxW7lIQc2IqN7jBd1I/k4pzaZYPosNQHq6NOkHcUHrmwLXS2YmPPOGxC9YoLD6Ts
Z06nc08aQoYdls7Q7hOcjAza2C9bV6ekXwNopICd6em6WUmMK4gMK44ih3zX4yE7
2SWGTb8WWHQCQxGAIsNx1CrvBbQV+iipIEwC+lhMxIORs/UqzgidGUS8fLa3CElk
FnfXPpbpZfG8KJKLPKsz8JYigoPMJpWpPTxfWBpvSCxd/CvkKCpkb3DWh+bbHnLA
iBC4Zz51bOWbV/rXjineTeZbindwmaN6XowDI3RYciQ0iw5uTikDiileXTfUKUox
NF0JD7iEqjJSljw7xRCUOfRGdqeMNX29fLCSwaijidfj79JQo0jS1P+F8qucUmyu
angjX5c8CQm+G2Mfmu1jsA/Q2fb9OCQCPkoDaTIxT6J9xoMOSdEo9pDLH/FtbM2t
tmFa/K4uO6T96Ab8RoY+Q30F2Rih+ItR3WgZ0n1bqZz5o7308uGXgxY3iw6nZeit
lTSD65KWJY/zezjxkACJom0bmAXp81nL09i6CKGkxTdoICsmNgzL62Kv0QyPEPNl
q2LhpHsNoIWEWnKOgMf0Ru0s80IAYZMv67rAkM0XYJaguRiozQmukO55hvLNHCEn
4wcJGFq0xdzSpOvADqMthKYBInpHRF9iNCguOVwc/bCtr81Ai/06R4hWu2eZs5dW
iYg800CG3fDQb0MdVLVoDq8qPqcShYyBo1XTxLjl6ulmx6HVew4n3EmhfOguof/B
P8VLqMVSZwVDBJOV3aaEkxJrC49hn1We8aK0CkjUyESJlW07lzpOm4etu1akN4Pb
VQzYndJiPcqAOIK/ouyDzqTL+7eRqyiiKt5+czILwHVewE2bx2FJIV5OmRtMN4Tj
Q9s+7v/kt1nKWwe3IUtiUSzDc0FLgHLgZcYTtV8v2zXST63g2SPkSaGzHEo5Hwwe
4cvHY+Cchs5rEQoND3PDQBYvZCLIoHphqrnDAIsCQmiAISzThJcXMi8CFsgS37Bd
YQfKmTKCRyJ7x69+Go7Cr8RsiHW5wvEDXuk2z9WUj3cXaESPh0kFdrnIF+XjStWG
yce1vDshZAy723tVuH+WLnI6n0RZK0Ve15B6QqmwD0Bn/A2kWYzOcEQoL8t+3q1e
u2eFWv6z5ELy+U9CwzhNDIyIImvgePb1u54CLsct5mzAca2rSXFrDLqiLY/uZfu0
gBut5OqITImMhlghQTKpomtUI5XyLFIRqeMK8CEmRzGOE9dAY9dJlE2Ku5hwQMa1
2eCe0Qrw5l7kfVHFPfqNXUyxoCeVDMrbf0J5wcQA/k3xg37sNGpeEPL4/Pw7cYgJ
9FSCUuIU/e7p21a72uBhgwrhS2ayPK1EkNXbC4862gWQ1i3mPwoxCcVcKAiN2gRy
safpHYwFTx9ghzFU8PpA7oTtKfN7GDU2+pMJvsfLVz/UuCRM9MkvNyU7bKT+SPxl
PjqQiIaapCLVZkpoKpdliAlwpsciawVGDztN174WCIu9pQ/EuO242vRwf8dxCFtn
FpRa13lv0gbuAurrPUVFvkOFBlahaPZOs487b8FSl3qSQ4bZltMd8xnbAZ43oDUF
DPPSQLZg9UqfoRlK+ux00oXGs0pea6bXgh8HM2/yY6QiulsuXDFXh8jq3tu/eRbP
gAKzhjbUe6iVqb6nlSeFcBOZqKRG46ZDcd9MFK5b2/IjAtwwDNL+ZE/i5B0PUPD0
2SjAGh1Wz2HUInaCz1slOqPqYSK/Sr29QIrr/KV6cbvInXoN3NXoqMSOdp8dNWgy
99qiH8rJiHLBzcnFYDyrw4K/3g65RgXengDqCr3mXtfotELpSEAqNnEyeXUGQRpe
+bYDbfeV1YaVvw9zWLLUph7zdGunF3TovrGN/eUu4WWkeqMvF47nUSolTK2jmLR7
KwkXqvvmKiJItEr4zBEiGgNv3YrePfzA1ByDRSN9bu57ZZtyVbTFn0dtSkVEAWw9
ipGuo+wIqEhG/15HtQy8fUdb5h/SNVffXmEfT00J00xKpQstyZV3pygiLloYfk1F
SPS92XvICY5cIKOwQwt8tYGATqrLLwpj4JASqjAH9ZHadBKKl/BpW3SN5QwE1u3O
AUboJBdM5AEfazRsIQXcBsY6eoapIlpZCkD3SOFxF6n/VW7F4YXeEU1A2EQMQ3eQ
C5JFe1p8NHN7NbputlE3O5m5QOTT8Wg/uH3Hl4G9Kj8XGClZ/nHB1idJWLyLIv1c
lD2Wda4h1apmUvRO3hNSTRN9m+EzSZEeVbJavlyN9MsPx48BOYOA0ObzLhnXnnwM
G72oeKq7MOhkUsAiV9U6wMC/pNNtdPW8uZ81XMP/LB4vCURL/lhVaHeXR2IdxpMW
Pu63mzG8aUUOifLTLsPnOm/szQRPtjuq7Fb4h1XcfhmFaaczCa5fIsnqvZTallgQ
6OzP8tOXwVzSiKTJd6zI6Izh3ECQ+CR4kf9mpaxh8OTYdR6hllfS69hgoEmqasOp
kbST0vC9cJR+mompnZuRZGHKYpy6u5i4zSDT5Pgk/AdWssr11EUH8Ma4+UNHB+tl
G4DsIV2No9PBZfEG382v7A6Ju2uMMd98PoMOv8VZHjiEDnsxCKas/+KcNnFKmOGw
cPf7egzrL6lF9gWV9uQLX2MgUuSJdx7rDpw9kmbuZ7OvhJy7h7fsim04MOnnsXSX
CmgardUZB22GVPp241DTCTOLX7Q557azFl3cyQzu82ld0A2zB9O/PzEMSsjGaATY
8oaYnvXVkSu2Vptffdl3APCb+7dUB8eAKhlWNx8PArF+dS4aq+JLwTDAm++SuGN3
K/sdL++UqUSiNX6S899fCN3GczxrLU6NiuIXsyYrEZ6OLaIcrGNgHmRlPJ/MSBKE
keG7HWFgNiXspxnYe8viFzgZoDtDbfwnUxhj1CIqL3B3Xy+PRBSPDsmXBuyJk+ri
+ncBLlf7kbUDAeyW/r5gm7C/BpcuFPytuB2lZRNztTc3U/GOnQ8bPNrzU5NTVckH
0CN3o2HvvodJ13E0ppyf402QI9O8CdvGfSh9fb2/2qYGeeE72eLKHDdK3A6jhgeO
URcskyp72yR/Jjx3+o4otMxXowDVPQv8tio0hecW8KZpwa+raA0wt2ungGGkXMvZ
sMK4O7uoxtsrDtdxCsQob0FmmIc5ozcOm2/W4GoRz8YC01u1xNh//rdQ/4Cy/yQu
YbcIT9vpEhXnF2SrPW0637tZVphaFU2WUixI70aLPK0XeOG2zIQR5kJHd2kXQyBq
u0boMudurEeeUjwAWZHfSzvOelvPKNhjUJ5DNFjGuSw8NgPcU5DB50i6ubbaJATz
6lLIdjiOpRGxD4sH2KZ5hIX5zKiGmsH+Wq93olvTzIW1JVRFAUOtDA9yr3aPw/WS
4+vOchP6zseozUvoUuoQTwF/BiaYSsUVJxrEU5uoBKG+oIHDgdgH8JViVpSB+UBU
0zXpSo+64VFU/x/7L6OJzIpI9PFGGmmo0ppBN0hb8EdB758S2uECIct8qzoWUREm
smAEqRYNg85jTlSVADY7niE8duYuR3sQJnStV6qTc1HALXZC6FIHKU+xlSR2MGg8
8gmlG3LUedKqi45mfn+3nEyHR8LOBZ5NbLzst/hnzWfNzEiRSCgt8bz1slyWuOl/
gH+c7bnXsEFppM7QJJBEWW/ZSzmItexvyN23LwEISIu+DrtQ1m3Od0PoB8RmTCCG
yEC3qraSwBSw+xGKbLZeg5jop7hVox4Tg35By+rqMYkewqUGRWH+W7O18S+67ZTh
8tLe0Oqq7JoxLKMNFWaQhVZl/sMW9e5hK56wOlIjNPKHJ/stP9yln+kVp3zweGMk
SLAPHzH+LoSo8Dz5PSTIN051S7cw9IB54VG2m7Wxqp76FoLtWw0cWFWXk0MDiQHo
hymTFoyLajpcnWhDkjSanGLsMklAT62gu1BuWgJMV6m38YMACllHhhdgBT7mWjIU
xHJadfGY0ihgE/KTG/pofyfF2g/Ynl6Yy/vw+baxXCv+XZhRsGidfRWIs6od/p2w
BveanunSOg2OZ533V5LbqKqICycLxHGR9l0D71musHk/sAOkywEwP7HyiYsm9MRW
q83BQ55rH8Ij9G9vdla+Qume6KTm357Tc0U9IdK1spdPgcM+08S7r927NFUZbKql
eaGxqu3CNW3d6inmrWU4Eu/dm7pkwZ0VexBEPZcQktDb4b+jFNDSsmZ7t48L2OTm
kKgOlCvA2TlJUvimbebr+oengO3slrJGZcP3BpsKMN0F5PFvbbH0ur54q3W/gmX6
M8sQi1hwEgdeGcFQV923x6cZ32EMgiQLUga+k3XC/cotZGKww/yPZwUkBEyOl72j
/h7J+UExdnaKfbTSlXEIxg0APeTX5UkSRx378EsapbE25oG7JAkYw1KIHbiven0s
/jci7otp1AwBqdcdjtSoZI1w4r+WVZRymeul907HGuemh3gEfj9GRb1otosCwhA0
7f75VnHnhFKoK/1n5ALKgGG42FXFlgYYmRkjYTKnMVKF0bXZNZfa3Q1E3XtniKFj
bbdPbTm5jLtpPCcXdv37AujuwHMJu4PVg4pr3JHzifEumTbxA+asKU4ilEt7lWUn
oCVGvbo5hHhoI81z+650eiDRSB7o3cvOFF26ETaWkQurGjAXp3RXcPCimHfDMJMv
cVaJIegeixFitv6V2zbVjTOY50XVbPe/S52/HgeVyhXLYwx8VpN3wzgmsUVaMj5k
nqHCRV71jWr+lJfhdpDeRrg3aS0IQoIfK8Q0qXy2RPN4W36gND8WAk15bdYo5FmK
I5UB9MDNTSPBD8Z4OgY+UF5P8CDwZi5oA9UVVnm5pnh1P2fb8ybc6T4JIWM3fqXe
a3+O7yS7Zmi1i1KKNKvXLpcczHq/VXhdd+Ukk1UsizSKmUMOw3NBPeueRV3hV0j7
gpjDvjV6TwJmNlecXJoir1wYGB7LhsNIWZERZ6FkuURPOiUQURabaDSfg+1p+rQa
E/AJ+kCY1LJ8VQ0GUiP3xvIuCfYfwKHfJ15pXu0Tmycy1cnhSblhWChgYNM6qzw2
xmn4BCMV6+PhAdYVtxJ/1NgknMnZ+lY1p+lF112gh84qFTyer3k74EBw9+I/wJkF
ol2EABgglrHNGD5OkfpvG3GSguc1laZgLbpa+pTPn29Zx+pPnVn3G4krvbzU0vuY
p+HFUlhQdo3M6ff5kDq5Gq1pZAGaD0gFSrEK09IiNwwzi1Xe0JsqHeT8Fuwmger8
OGls0XPi/qAdtxS4unF1XyVx4Rh9xDAaGk8y2/5vxd8h7qIjIX0MhcokqZwCAC4F
Ulz3/KTGee+Z37jP2gMfAyM0cCINdRqUtpfe68Eg8jHQ1jm37HTQWwi6Kg1VX37H
Vgb8nd73LQGdMBSkS+S17OcQWE594Xet5HhEd9Fz/bUKLUCBZpreD0fVWlTgNQGS
jgaknjqDAqV3yhqYbbgbwtQGT+edJ9iu/EK+tVLiqXGhNn4PkPuQwnGLO/gcFxrp
sOiJ1CK9ULmbmVVKvn/Hqi/rrqVuHoDx5Gq1RSqPPTW3MY5rG7EWuMq3p+Evp3GW
eHtED31L5ro9er6HHtUmjsSg3ZzyCKYF0pCmwvfGvuLpO1eHA0fL6hq4GsChNPpY
Rk8dbfzWMa8P1Nw8FJ8tm+TuPA2rAL8MJ2DQciH6A6xXVuIcj811X6xVg/GfRaRz
kv2f6HsfaOQYJWmzDEG/jsBKDPrjT2cAatB7jz7ETC9CfS666MFWrqSMBLdhWlwo
JuyIMI0+HU02+2kJktX246GarOhxILdYVdywe+Z8qepWIyqxmAaT3/lAFB9N9vFD
Ju/9I91tPP/4IV8KDPTdyGks5bWC+Y0ZJl+TyQy5/KUiLEEaQXKV8hqm5WtY5bKV
S2NGFreHeDDpv+JTzFADVQGH3OjfBougss1Hb16vEw+XO54wWL+pqsBIZ6LZqtpS
AHlASNbp1P/h2HxssoT+1qVEK7H5uZ4Dg8zaJFk9l5eiLawWbzK4hnG+HHsTjUzd
4tOziAtqtuKyQb1mZ5S6gDySFY9njPUzEUHZznsR+sFEBumzI6Wxyh9fmsx5KGf+
unIkO9U47WpLUMEqxTH/Sja4DxGSdn/svyneKPnh9yiGZ+41nzs2TNCzsysL2ofk
6Yg/HWMCQhmiM35daLdk+FRHnEytVMtnedugmAXWmFGhGl1zKK750j31yTvyMTXO
S2IRFvv2eRze+KkU8B4ixB6naufZBYsk55bIiVvflFOcanHSJ/rU5KLFSTPB3Rw9
jTuI7J/FT7ZPvwfdFghbGMyY1wJpN8/0c3L5lCrcSSlZiPQ7ihcV58m/ODoCqfI3
BMQzDIsOM5ndIkf9F5pYyTpwCPSxbb5gDtRQjEA2q65mCu/pZScE7SpPInvu4V4I
iL4DCiIugA7D4X9WJ1h1mlK3jGehtk+HxPuO8kKRxBDDWbxnvWRROzpiiUCl5fh1
rt3TRS49LBvXpr1ZiBW6u4GzGB9MLbcxaB65KY9xqtbMQ1GiyD1XoDhtGxaV7rsD
uN1LLF6xrhSFxJ7EpSEtrstdVuudU362WnjdschvalvYmgoKwUN0WFb5M2hjaWqB
1720jQlYRfjGwnl4DyQvRLnGLmxsUsut9lr1DI09RmP0GAOG4piwWaxBnugSaqvt
Ey12UpoxNLFWWx60tS9wh26WCDZVDAEX6KctJ7yRoqZU34hOmiIJuv9gkgH7w6Ul
jEcWegU65w9pJ3HgD53J5vDR9vi8qW8nbZePtphmxWFmcvmnOuLKCpMto8JWFToZ
7sm2uwz1RRlwrkcJ/gM6SuyLhPyjcnLjxNQTluUfOha/GrnFwEumBceC234K+to4
6U5KrzboVUpgqRNjEikNRzL+EPBV9JiI+wXf7dpyi5nMNOe69/FgEyH00+u11Qyh
CwJn4SqTbtamFaIlmcUGNkkyghYi7flzdTw5pZuJ1Kcs6GPmsFkmkNzT+4JO9OIw
YSJKfGot7cz25pVCEJZ3JnOCHIcih3RUuRBLCGobmdQsRlRaOBEr3Gqb0rsotzPI
zZ1AoF42Ej6cB36Uld3+ALqzlmzUXz2JJ1pBh4R8G0TJ/BGus2lKMzTsxTHtIj+B
zfGkdNS+1b7KST6Up8roJaqvcfVjy8PqKeFCZcgEGP0fRAe1tP1571n3L0Z/QRAV
5PmKGX+/J75OO4exMqqrcNL5WgoV6OoJq7VvFI2+n3BUNVVzdmSb2R6M+Gp2Rm93
fdvf1YlIs2zvDjCgViTmM9F4i76DGi1bC2v0Y2iANWJC09iuC1GTpiV6lBpiYtXj
uvjFkFRpn76ABzAwMjM9V2UIeSnDixfOVLBsCSZoLSi6AIqGVdCBvlgfdGKcqaaK
RBiD8Ja2gmRWOEZx5bNYKApqNtkDmhkSu7itb28AkWlrpdd2JIETCxeBTW+bOOjJ
UsXN16MDiF0eg+qyCdSi4vFKaVF1pT2pQH3u6NReAGi9uNpxdnf+W/mdl9vM5aii
tQKCeAg/vJ2uakjTt7JWsYFEmMOwITwtTeRsMte7jJERGfW2cVeZ2lmvWLISO28U
v+FRYJepo8+VH0N4qZLFNS5P/RM5oTFFdk1TNoqLnMV+XF6bPwoln5BmulHAF3Sf
hdoZOJK41rqQZlf64zRL5K19oUAzTvLM0KNxRmW9SOpaDZ7jlZlXWvsHhB7TjVnf
AP/fi/YZZMwGidlPqtk2YzcP+/2I+4iViR3VnQJKaNlu8b4TvtTBZrqcYOkBX/9q
mN1jsQtaDApM2zOVCFIHl/tdwjPhvdjUk8oZ2pbyQ3Jg9qHy/F1SGmV4WL2hN8aF
N9YYsBfrfgPBMnaUsEdI3FYb2HWi4g8s8PhiZiLR4vVnYZD3ucdYdqjtIxdAZB0D
x8IhwAsclAe0D9i8n89doyBqvaUOPDjtO/I0IkIy62SHSR0LLU/UKtzWHdmzukgY
NDtt0DMZD9Z+GEmypuchgz3tMHVNVq67hSYZFOCFgmzb9oAZbdT91e3U7YTn5alh
4kMDMJCbG4P70gwpa7sGQanl/rGBLJ1FcGPfD2yiimnLEd14NELjn1guPnKkONBC
TWShnpY7JzBD4E+zGikfJrewCjjMz31rBh6ICdvVpeff8INEzIomH4bNE1LWy1iP
QXgEeRai2VTMQsm/sNPKiT/ZtlhyTc8Pf7NK+7UhoWBVsusBR085H5sFgaVY8uQv
Ja9AXgzis4EYGaND5DBKIXAVtWZZmtQw9NIhbFZFsuN2MaL5iPMUK9H5oGbfEx3F
KTzKCYJx6AYkydxRcNg1Qmr+pVqG2E9MlunwSBc3iQHbfvw5CakFaZ81g7BiscHQ
gviYo/DUO3/XIzzwWcoHA3NGpV5foHAFr5C3TiVFApprouC/zXvdLp9ToFTeIVJ4
o++qjURwFqooijOpjTRpHtkArz1WTyn8o7UQSqqx/jkUDww5uyxDfeoF6ioQ1LoO
HwBkmrB123a6/XIIajtVqqQ3sF9FwfKyiTSGfWwrfkJnT8SISr42yQJ4RYVIbp+G
BSNi128PMg0Kdr9wv4K6TecDvgBID1HBJbZiWNFxbdK3q99qLIFthtS5aaeshVhu
ADYcIUpRwXcdJWGbKjRBfn5N+rMmO9onGlRZZ7aJjB/YivsadE7X2GvmGEl/w+0v
w6MnrDW66JAaRxKjXRh/uZbwiJvmsDJ4eMnjlT+gb3ru/WYwOLn4Ijz6y4A6Evht
iI26jdOPNkXNPLZn/QbEDwaWfwvqxxXswcQFs0Itv3uPZYO8tCO1SFdN8pJq1Jdh
ce1RFrK/WOKIDOe77GX25zJL9u4My55YPnQcGeo8Gjy31POxv/xoyOz2CIAFqny8
imcVDOhUW5Y/pqtwjKKHRcpdWDIL5A2SaK/JANwE6gNFO74TUHxKF3LwnMCp67i3
NhjT3zZz7yQk9sbMfbH7EQA9g55DKYEisLEsjmjvaasmgcx7WEIvOG2UGQezgtoK
IfyiEVbIJ9mKY4uapi3TKw+4muT3SwSurOUWk67vFy5+jfocBlnASg4MXnH1htRl
HqIlqajCb9kMPYqXEOZbb56ECBMc9V3oq1Cz1V83XFWFfKgDov8jbjb+vU2aF10V
fUo3DFqnKIO8SunXtBo8Nk9CiAuivPeQYVLw9WygcmG0zW/wqaz1bj9hTdDVDdZ7
IdzPSiyaqT/fYvKjbWxNvSAZy1tJNgpQyH41gvh1Cl2lfj+IFeypJk6oYOjbi1mc
wZTqL7v2vSVukPkKNHt9XrNfN9CUKxb7x/FRHuW+/Z8PRA6/v2zFA7EFhC6/rSon
dZP1yqLLYEdVs5ehec7IjOzbzj4tduOPxWWZg4QWeAluugdqp9dTrhPA/57Yd3VY
ZMIuzRRxh1gX6HSSRbHAyySCJiaMRG/G4Cu3h6PJFqy+92smj0n1kUGVamUrLqE1
Xpw6RSn2HVNDyWycJlKtEwWgE6rCT9i0EGFF9wLYxP6vY0zPUF7k0Ymo+EQW/+9B
MzmRKvHZK53kSkkTi3xDfgSSeNND7/TtdaC7UCIsSc/1Ueegx1XgxPLXQ900jzVj
RprYfNyZ+4aSIDEdnTulQ/yFIxeh78ekg8Civ1S+4AExoLnN00AIIqz9CO0kv1y4
EjqRFJNA6pSiNFi81JZEgfY5Sfjf+WuRIwTPfY+fDy2e22GYmy4hlch3lh0ougR6
4bJEJK5IUTG6Ut/vqII9gsccBiV2APdCkOCw3XMUvVFtYwgpHuEmLVYF5iWeTVDp
cLWkxY6JGrdSgyEcU93HGWHdlem3toH7SUTEa0gNuL61EW4fxcaZV6C7+v+gYXJ7
77NKeYitMKZ1cFPWJ2c1E6BZUwlzCI/ndnkOZBpTHBYZwQCUNE2DsrNSEx62ulSt
Moeo7IH0sGoWP5SrzkZ33FbLcv4CFuzHkmxC0j5OV8ibGc7Fu6XL/SEbXm4tPsTR
E/t5N5CR8hEeZr7XBq4EQUl0JdbzNIbHrrIFmaTslGMUPEeGixHdQUWNOvmYeE02
1qHo8J5GX54FwXCZGlVY1DYqJD6dY1Jq3SrGkkfzpKLwdZyoodellLOWYsw4Fv1t
hHT0bfVjOMwd+qcrI0MeABKjC83b/UUECxxlPjXthWbf29CCBuXr0gJQ8MpVuGPH
Zuok8dWCLsVB2wnbfn2M6pFop8ceIp7IDTCfPsG3nA82x9MF94SpUXN+d5xAC4Ih
ana4T8Tz8j7gagqvj2MCuoJkLqFkdRcjdIylyTiO/xdpn0FdxmUcFdZYqF9AgzVb
DjknX0rB6t52FW2Tpf5XlsjNnopRSNxb5XpaNMXLTgKce6m8Sp6Pu0tZfN2knrHx
X9d9hIfmV6RIyW6sLYekUThkwG7kUI/lSDGQBLliGZCL9hWdU7MRG5p1MubB1Zwt
H4soZRkTA/l9d95mw92HsK/VGdJzq4y3ORfk9XOEmd3+yHAwKnXpN8p09nf6Cc5T
g96bR/HENNezmW5WUTCayD/PzY+HTmC+zHZfkrmwD1olZgmoF539HdFYU75p+ixA
TxHDGJhx+0jtsje09OhFukjEIUtxjBg83pRNOHPD+C4laIaW3nmbNhd8bUHqNh8h
J0C+8FChZK35Du7tAkt6S3vc636IzZPIw4SEHKdQtYFs96BGn/7EI68H32VLHKVH
FmnLrZJqrFCCvojFsQ/tkudkZW3PNc2PPxjBRcT9FNyDk7zO01UQEKrCu0eUJkRj
b8wHsLdsf+Bi5ZLVN9dPQ/1lIXQzTq4UrrsP0fjHite281tlTFfn6w2RfSvH8eBE
32udYNO/y1irOZM6HrAyMJAwuDRqnv6JHdaL/DC3e+TkTDUo8ywYSEku6mgup8vj
5i7B8TJeZw94X+R8gzNcpq4EcRb/8HlbOP4w9XnJmNkOaz3xJSpAfouxosEAPEJW
kkkNEofV2fI6guMOQSvFCOO2GkxxQXgnOtJdnSYLDATY3wB1yLXGb40RkEPhEnvV
VL6hGBAw6ZdvZf9x7/KtAaK87V2bOjjomgO+adhY85weKgFShilqYayBt1SmLspo
fxJBbwYsyqTUQOARE3gajOE+nHCvM3XMgSKfPzV3zXD/qxh+gF+ASJ06fpp2DLiQ
KB8nG9RNhX2eOctWJ8uRuZazoZZiro+ILxdTlWGWuXOYDzaZDszbktdR0TFqg74d
SmD7CoO3Iqs+x51TfuOr1Sc5//GRc050MfEeJPVxlzs/Q3PV2UcPZSdxmESBldaH
bCWgjyOzJqom5STj4Dij6UZ6XC1uFmB6hcxerA5+hhpDYX32BDcaVHPJY7IrCZQx
ncyu4nBcZrUpVRxyNlOIly8UGduYBubQ2Jit/dMXNthomQM/W6oLimP0UhdgcedK
DeQ+poOKOffbjeo5qeOc/VHVCNjAJ7fxrFwgdyu+tlPpdAEVGWHgHyO58ukw3CUL
9lymHYMkbBLAbXC/q6WnKj4b5H63kMjADIhQLy0Gjo7uIcMBVw/N/Rs7T2FMOb8U
4ACwZRQTjMyFnXB2Atv21dy89G4LZNl3iB+TZzBx5YTxOAnGvNqNaHh/3xUIgs33
xEk3alYzcy48b5S3+XMejir6/WnInV7LP27/MQeO5h3G5x+Db+7rniNm7OWowT3Y
XQWTPqLx6CX/MuE963Hey8e0BOQeA3kYFOUusi4kFnqcEQlFeFeCfmm6LLeUCGia
QBWAsbLUa2NWXugSB/hTgVTZK29vnR0JtSY7Tn94Wa1cGeRJ/XuKiQGQ6k58YYgZ
J9ciNcJ6zLRgIJehgxT6faPGOdlR6z75f7yJgo7/KI1bHMMKRGw1CYTk1Au2B1vH
U+r9+fKRRhj/mEfDnTSHN/CeeGPvM4itYBf2xc3C2zNu9i9yS43Os5dj36wFs0QD
dKp6OeCMakYW1H2faw0CHu1cwKpgJYrmKQt0z6umui6QbECCTDk12q2gKmdHDzfG
fxYN7k99SX3Hq6nE48/qsDV9FYrfz1af6z9gw1WBEOP7sRQSHZo3t473fJuqyceA
795D1oWtCggJ7mCs36Ji3aHDaCfxdyAT3uu2gQRcmds5YcBpnNwqFLuM2gXwnkAS
YXd7zLG5J+rCHzBodoLS5u4RZr+Nn2ODDP8NlThN1GOZYIdYXqPLNEjLNceHeANj
wsGCH3ildTzeLAFVIV7Ou22Hn6NhvF2ca2zbj5Fye6lapL4dcWEJQScN7XR38jci
kIy+VNRT8dqkxUUjib68rNryyY8yw9vYCH22hLiuPqnliZtcBujCUSu1mTIAjldV
p43iMvTpHpj4gSGBZk0Xan8g9jlg3BKQuK9hM5RR2RrRq8sIZeNfx/lvJ+1NOfrh
Wiapdt6tFyKyzt64iLamASPkTN6WCtm7nEd5LmNh2tyMKXWWjiZKcbMJBmqSGZAw
Wf8+hHSVA/ypz4ajcSSLW5lWfDHj3PN83x9HwHT2mpoai9fTOdAxYYOufLiJYF3U
PmLIfv9iDwkDPbqwB4tFFMSM+eZBhJNc4NUDfUgYO/r3ZJI1RcFsD1p1Pu3ltTkN
fyjdf8vMzCmODZNMWfmNLP/kyZ/9rDXbhwHziGvhbehyELCxuAufn0CEN6hVPliO
kVgY62aKFGf7fI0q1pAyKNuJeNv8jDbSvvplZSwVpW5y3KxmKB63daHsbDmvlU9P
difRw71dHYtrglZjonZ7zljGkmrPSDUDPK5PNxADx/ozVdBXih3ic0paAOU9jHxl
I9HHu507FF+PHROP5XFo7fOI8a5LZiXRvAqQPCQ6XXCQayIux/WK1WDzzPFHkUu/
FB/AHea0Cf47V+1vzNYLPUoCzUpwF7buRlf99IS4Q1MpvKpqlGeSEQoPRMyA+Itx
ZKTOPGEjLFIAXvATfIbePRgTZu0DuLLU//jvYs0qDbtDKwt24rz/xVeQlpreP9Ix
NaioXN2pt1z2/AikfmctTzC8nPVk2yJKCeRNhwwrYsgPdWrirQWwkioJiy44sajN
cHZP7P/RJrgDk5VGfZERUHGuYpKP+rTIXnlgMrXWlBCsRnBZrxU4vyKHkQTk9oW5
lO5p+zrgKCGVhMjiewHz4PVkX7u6bnmZvOedyee7lWXAXQN0CyQzMF0xE2tdlHEU
N5BMAhkqqRTlwaPfa3Oh0YnRm6yE5lgCmB+zalSYHDQsRB44c4325n/cxWd4n26E
x4xHlZZqaMTLcZgYcIH0dfvIVW32tIMW5Y2J07itp8VeWkuNf4IJvqPAMF1fpwRq
TI8H1P1Si1iEHPmPy1bK7ghLr9pAWhk7iT/lBYdAiHUZHv/kpUQ7nmblQfuPnM/9
m2iasL4OnkbWu4iTPkMnvt9xMfubg4fyose2kmhc2xYThV1oaggLrdrTJm7hsuUf
wVPkRwzf/rbPI0olk1AwaX2Z6QNogeoVMRQeCbCQpIhChEFhPIHDICRt7COxwD6i
dCTYAYXCn+zcIbbnENfzUOl8gogpwHNpmEeGz1vPWakHOrl8oBRs3jepgd0miAPA
1rl+/xvgvIU4bb+/CilTMNePz/lKD2iAJdJeUElQc7s5ByBU0rcqyYn8Tyw9TutY
m31b2t3TcMg8aseQVY/N4X65OyAHUP59txcZtSJBHJ19Bbh2WPMQzmUJG3XwIq+a
/1XmX9zxFwTJknIUFMKjPNL7qnwrcvGmOdG/nmbnwAtiGYgb3tNnubKdxhH1hGZp
ySy2TS4FIafN4pFInlw+x3dKamdmZWJEk+UYmNflY8kIVDE+xuR2gSQUu+VtOnTu
gbgJDkuHpwAJjDUab08LJZ5LgB5/jNmCkgh030FiB22Yk7n85uNA8JBFN/+YSOV/
YW0vMyE6NT25obfzKwDKAoRMceAh4hLwYgcL04z05rkOikQDBx6vu/9Nk5EGs/Uk
V8/fPGL4zC3nUTUKn2hlVPu3XwI6Mtk8b4n1YJwCwC2+0uzoGkpwahN8G1tgtsjh
B/3dR7N2AMINzglTdmIytONPne6xQqP1TBWFBSiTCkTbFRkBdkLXq+fFEKT7d9gA
E04VgAscxr3VgmMIVVsXEFtrlWqLoZau03tk+ffF+kEGPFvAmRf48XpZTc/IzmZo
nqccadUaa/gYVPYgMRohUfItLgg5tQ3+ym/IgAhZqZcm/20iizvDGFjkOKrEHYiD
O+WdV2mfP6Hc6GSXW80BMR4nCQGzQUQBhh7p2uIPQx+QhdsKWilGG41Z5Mu6skb2
oAZcJmH+Ebz3PkwMx4TEZqyWWvKa8HZwtJp1hZyjvOngv4BtldzWtWwARiVRD6JN
dXIt08Fgc+kewlT0pjy4Y0AshT06bz1D3JFTM2u9V4VEs9veqO6B3sIGHOpgh3uq
NGTf1VgRlVmBzz4QjO5dy7v4A9I0NjhmIBvu1/ksFof8nkD/P/URDe64vpVcDNtr
QFidZgSauBdHg4nJ9sXiSzCrptmPL2VgaEPMrM3A4b5pLa3wlou//qXjR5B5unhh
8dmlQFLSufW1f85xGGvwJc1Qo4S8n8bLSxsaE/HqCslQBoh+Opi+3A8bLBsYvKjy
WoY/ZGTCnH+JgSd0E3NmWlwYVPmU1uNlpnAHZ3hfgEMEZKiBadX6bZlQHKJP8F/r
4OXKupFotHyUWFsxXigkHqv6vKIXiKUUQd0QUI0MF4QJ0bSacg++/QJV+xa4Hkjt
5szfux+pehMtAt9xJLDS1o7QqLXQ+T4BvQca+3cYih6HkQ86voLtubYUCtbjaEM9
IFfo3RSN0YLj+2Z1gjbfX0QDICR7ZcBBwrP0/S8il9Pvfwq5Be6lN9hHlmjZnQaB
dySjzgCnnNKIBieageXO9gaNSC2NVgkcnM3FMMntiKlkBVEv4Vnk1a/7KwRKSkxR
wLZRrtaqjzoRCwHLsrJm1M+iVvb1KG4OvzKzHOygAJEdIZbDXf8hMKds/OoZkgCT
gQBTiEtziDWRg1ItYMUdSZiIEyDpjiMHsGzmJDD568K1bJ3aKGNHHa69zMx4WREA
Lst2w512ClVt/iCN7Tk+dO4mh/NscqFBeWZ5A+cncoQftMPKWSaHtd55Woqc85lr
XnA0J1rbwIl4QgozL328TgOArWWrzHRjmiNfcLvK+dn3so7aTfHRiccE6rwQIbyS
OuxVdOw3C/Acqp3l4d+IhU3UGWMFdn6x4SRhRJfTrKLKTs7QO6/rE4uWXlGF9FpZ
YnVy0lne02LtiT9j+kCEEMlcU0bJczjCdBu+7MmmqqLQBMB6ZPkfaitWuchid1nO
/rtb2UQJ7QmR4bpS2KhZN2OGAbAhPpdlkmJJagUGYTb3mg2FGAtGH16ixpYRmpgm
1pdbuH00mOwvBLXLnvc5nayP4cbeM/Go9p1SNJR0UI7pAtGxX11YGdIlUJNCIGLx
lEvJ4nT5iXPrE2QpsRVPlEA6kkwGXHGLyl0gJwljA3JRIqnX0dRJxyGoTwG1YB0h
Jk0I3mITGcBDmrb+WfArQlhSK+PND099OTDOFg2quXRD91qP7SIYYuVdD+pV+53s
WlWWYYix5roLYwXbQ2lr91w8I6hQnM70E2jiUes1F/Cw0g00hVrM5BgO9teqJDP7
GGv8wxfw8M65Y86TdKDr06vkd2tQeZz6+alDYcrJmfSn7s4oZBmJUpKaea2dBbNA
eELY+VB/gg/WYDnBmM1Zy3k+l1iodw3vLzpPDV7TV1UcNDsyN409qQU8K83onvrT
EZ0NB6DOJkrtF8W5OjpdjJm9dXsfPCpyDi0M/EhyP91c2Zk1lxPVYIrJl0a20TFM
ozkkhRaD1XnjWiWEtfTf5GvXd/fyGD0AENG9JFtnghQNAEJyaLxzwcPu2RYvGZ1c
KyVAz0T6TR2fCYsH2itGrZsiQY4Ud6C0qJVurkbCNC1FsVNSEVn7t3Y1BNHxVvmi
PBGzKo9eRnbH8xOw3scFpWHaVulVfu0Zgg8A7ED26Sg+H0KLbBLRrTYWkCAfqQaU
v36Ger+zIymwU242w6eHIV6Blv36ygV3msAr6LvaOCYdPYwFA9GNvR7w1GIlBs75
M59Ry7VixndkgKesJzvc4k1g/kW5RXIGP77QKu1jqBqlo5Gem/eKsIZCCePGfqw9
tYaE+1x7VRbuFtzQcGkTN4wD8NaVE+CGQgIsjaDrLuRGxtmcTrzSyJWjOVvv75/W
YIrVoeMXKE9RyOsngMzEtg45cMNGC21wLkl8NePD8bBBwt/1OLBHCUlrnHA2WaPa
IOj66/LRlo3Apvzvfj41QvU+J45yl6qArEr8mc//I8/BllRCekJxFPtf6LlEMyhU
gPIYJBZZ7KDNbn7qLTUEBlm+ieVtPV24/H8r1xiMgJNg8IwfW0b8/2mS/WhBn44O
m3Vezk/dKj/aimpOyp5rRu3oPDvJ7LbxzAL/GIGRTu06qQjBdeOWJNe+EGgUXaGw
XrXdEfchwAm3Eb5Eb9hABye1I6KIyBT5BMVN4O79eea9Pi6zFqFlmC9UedszuaZT
iN94krAZVupa4Dj4cyEcHCqOI/HVgXmrUHtE6mHcFELl9AiPRErDY3tAItVaH3Xm
VawCXiiLpiAQeqaHYkiRpo7o9uoc+ktW0A1/YN6uDV58ZpJeAF+h9oJ8jELnvvy6
gjt/TyVhAfENcRvGwmsN9gp/Na3tufM4xqCRstaGEVLN/Rm4Y/4YusxhCNKeW25U
ULDR2VZKkZnxERwr3E1RIh4LGnRwIhad5MyujF0wObpb1PuSrfxEVe+oF3Jk6jmv
70Zckd1urtgxQt4OCoAAFS6rNQTvXNsCWKV2/123szwYhTRFeFWoXBpzBZPAQnab
/6MllfQibh3SkzyGeSGkU45pgJxgFu4LhsjzWfFHQqmA/e+90x8NWn8TVCcwpciA
g5D6xEf2r1rQtueJ+8JWMLqfBfj03m7S/EaSi7gtQ1+25L/P8+WGpPUL1U6pjW9U
1k7OYrKQ/gkIx79oE9WjsddDA0ed2JYo12mjqlT+6GHgU+X093kyjmPaGV88a0hc
56FLsw8JRNqWytbFx9fTM/jYFAiEP0K0boWzmeHhdm2DQdzLO6g/MKOI2MYjdqjb
2GyCT/LPB7Jap00ade16LJN7vwT2fknFtesOY00ZaQUBY1ZVLUeO/sW8aKS7IOFR
yjSobsYRvIx4FguzwkQpwa4WX8/8/8P8+r1L0aiyEXT1JZVlJL0ZidSilZBzqtrY
gobZMZMTOMjOkkO884ewbA4rEmvL0LgF0Wi/+cmbLajQ9fmFBNGo50v4YDLblTMy
98uu7R7bovnk2/jDMA04L+WWxPBf+/widiTLobPcJamZD3l4eA3XBqfmFY/rvyrP
wysW2V209WVWUBh8eeGxxqstnHCxiU/xY356MN99Gid36rB3fSQ+AAdvHLDJkX8C
qauvlyW3K9sxKZiPPdV2Q7hpjwaNKjVdyaLM66uHhgOrOTExnpqje7csfYUogHTE
oh5Ax60VXjFg4IkwZkgq99it3/3jfdRWJ9fp/W0q5fhfzy6IW3BnqHxWK+u33pTg
U8D7HoAR9Fw7AyVAhQCcKytml+XZhQ38AlHGpyDKFfxFJFq+zVBdusXsReDJSkiA
D6hzV81KFowEHG6YdtlOGD09AA9yOqd96CARUm2Nm+kV1jRdV1p8BGerp+Y4yYvf
JNFEBvCTGrND76tgx8cVv4XwSX9vUS5na0BD6UAkGji9iemRb8iASk7n35mJWesG
Jw2nhvloxI2S2ABXfCGEnqAWR2E2+CB3azI90dRTrZAp+FPmBB1xNl19VpmZsUe5
tXSX0l6cmhBK6ztuVLWMbPdYR0mDYZ7kRKtBCJ72pTP5ZPMcgbEvNBkcirX9aw4x
IoZqAntRDx+36RHpAgiuJB/6nmlOaLfbE8h9783+B2/UCjKw9Ctbdr5nleXQwlOK
rg8CRkymT4kbusIw/EVcQzGbkLLtII2kLE4IjqwGUG5glun6PUY4PoqWBhSqeSaB
LF5LHzKgTU/lx3tjQKkfAODW5xwmqeAisTs85Cpuj4kWGJORiCHIenZ3kk8TTsJY
bNZXlbz+GBm0auG/1Nw1tOWZmkuUCAh6IzOm5nf/0Ew/MOHe4LNu5nSJ4K9r/G+B
KK+clNBuAYzFXw68W4FeJ2HmHxoUfLUeXb5b+2RWhFVpaKZxm0G8cnstGy9P/BpN
4oUll6CcfkITDiEBS9G2K3nmZOAlCnAZqBHcdjpu9ETAn+VoVrl2P8dqByilQ1fN
r+FbBcA9Wa/x0sJWGRoLv28/4dEBfAdXslNcT6uprcCNMuW7gB+oU3d+Q7Uqvk9l
+ka5YrypJ94jRnLX0+UQ9hHsqBXE/tCnHEo1EpYno1TyGUDOl6zPCBgRZ6Yg8p7D
Hw6p8hUeLH5xXiSqzIDLRy0Y67TIEjkKmZYlk2Ej/ub5oXp2Ui7eJLg+WIPqXoYU
E6MkBcao7r8m8SRc6vkcFBOu3yLnhrXhXsG+pyPvhO4u8MfLEspeqbmuRKK3Yt89
4Ufj/CjeBsCg8qF62XtNdCC6EwewlrJRE5MiXnHjiJBU9PMjmeVSj9jBHW+1AK1X
rlkT0BbDknHaD9ZHQPKKdY6I7yE7FHNOZyLCtqlR6V7penImO9eGU8P/lVp29zT5
6PLpTcpi3aIGAQZQqEJtE6Z/GJjyBgS+GNX/FximKDrJ/cjvyzn8A13atZkAU9Ww
KROATvK1bD3T3X8vRS2fAYhg/7/0D+70s+D2rO94H7B47mXot8ep71Cm9pj5CMS8
iyA7rrtw88Nv/f4zzH83e8jPKXO/YE86oI1cRGh4D5oWODuCatBTp6HEkw+19AmH
uC8UHuu38y9rPessNGNpyMPT8VTplZkPEFdGSX0eJ4MTa8SVUgdB9iBErIeFdqXL
1yPvnRWIvbSCBIQUnSWB4Fzj7IGjOHZJniK4DrSWhawTT4mlJE7UC13SAeOfqoz0
On36bzSP7X62VSmqkPtaqQ0bQXKBIWCDrsGUusBKmPFEZDZZHlcZhawBAvhSvCo/
StqgZdHD9q7XyhHd1Z16sm2Gnkgo+zsmqlayJAqzJ8pgq6R4L6D80wIBp/kePg5K
mi2OZhRPDv+Y5PXbyv0KrnaJV2kgea+p2WjKjik/r0HDD+lsgrHsjPBduXbx1ElS
eAgrs1yHlDGh9E9Zu+l2qfHKe2WlNAm0UairBUOsD18cfP8Yaw+PaaCUiadmvcZV
J79adykW/9crrXHg2MCuZBSrDKlGmYQU/wO6/NhE4Ktzr68dqEUyN8LePHwtDs1Y
wkJdX0Srvy0tmP/xRIxOaMUfe3SFpPyQ2/2ZTKXvI3n+T/gHe2UZtyKsDuf+Wl+S
zZBRK2IeyRzhfoR0V6f1aocP2ZlSuqvlFtL4Jb0x8RISXA0gkiz1BQ4p24A713Gy
rXDqP5ui6MCKszuBF6k0ekr2XZVRYhnjDurELXuxTRxOtL3dkSeG8M9Ia7wTycty
lmyh3xUjpZqAc3H1Xnj2l3vORjasDkDf5WoPoh6CBEuJEz1DeJnDG41ziFQQOqlx
RzMuiD7gksOoD5yxnrFNFfr01UzwnPgt83zODHUYXnxxd/a9pbePQRgfyoxAtRXn
8nuiJMQgwVzIalOa/mMuGO/td22iCqiDh44p86Pw+MSy1Rl7KYZcG0owN81N/CPW
rNYuYdBN2pn4CjVXzlZhevb7ybAlEVJuKZJ0aAkxNEJfDjWq3tJj+pQj4Tn/pfjQ
0g4Wcza8+UPtLdSM5jxrUZySMRO9QhyjaDbHnaPHDLtci7VUYrWWmCR7Uyt4MMhc
MqBRPzbF/HoquETyWNw8R6LtZZu4d34vbeAkehpIQVMK1G9omQSXgnsImegBStu2
xfDXKCpNInfRxDHKLGk5fl1oLp0x4XOmelouVjwMz9pV8nH0elYsUaBoW5+cFD0c
cUAnLLyWriphyLHtOUgA02HUsw7BNZ5gzlL5kFH30LLaJUT+XZClTc/0ePrU26h7
ubc6kjlROzxqVlfNBHYar8uOYM7WFX99tpf4oAfpUF0xycmBQBGta1AqsWzIsYIF
dp2kLNiVWOoLvwn2+upihHGjPD4LfAwqnOrqoEk1KqI16jwGjQio1OaUi43KGqZJ
De24rEp6d4XExm+ud06CxmtNU9E0N4KSEE5Pt8Cn4/vAP6u/PSOuLz2PhKN9rX/A
FxUmzpK+kh/URrFQHgrzUIZDf5R88yM4jlLEUIRunT2nETh3uZVDdRUNf8s0/sCP
rHX9dXC0a+3QVnPlIejFQt4jD+lJLtvFiWj7+V5Mzy8s9qT050jdbb+g+blpn3d0
rwAYFvEBom/qQzOjB482VMbiPY+bwi15QnlxmhcUuXv0x3FnpV6c9rkrNTpMD8bq
bOEVxEhhyCvcguR39BhAylaISm4vP2GBwnawoMWfcVJhCiuxycgnKhQ+cMClbXaW
/YwLGgGcrz6OwZOzI3U0Tlu5beUKnF3b6zCk+xU6IeYcxmqVT/5h7m7yljahy0+J
FuFfa0hkpjfNCB512jNutNLAYsNqbDJIR2wULYPWqkgRAPfQoYB8wi9wOAa2ppIi
fAvVTmixdABAmEB01xNsN7gVXVudjKrnjYrK8DJNrZUlXvVg4Qumj3cL8+qRAU9a
q2Wt5FyiK+2nGsD6xZuVBRdNO5CTNYkMby1NOSBRn4V/nmaXXKm0XX5adJSX1duQ
9u6uzYZPmcmT8DeVlRcN/pEmb1ioN2TlZu/upLUf0JrGfkrxfChFxh7wHY8ht3ef
yRzgYw4i1rtQfE+rL3SgZK7vzQLEMtwKg5hCug5xSoch180Kc8pvH8MZc/1UchII
VNVJcxkWGwD3jHWE++00macT7ee6HN/XgDKOkq0DlgRE8vLNo0f+yYoon+pMRcVr
6G6QJEE9Mobi37gRkDe8gHUAdDYnOdCmC7EQ/D1EYVacb029Of4+n6oTnUrrxA1h
Zmzd3RXSRcaFWfomF8ZG13pE06TklUn6UMUvfmodeN+31h3O96LKZ90oVPdZzC0Y
0WOe2ZhbrldBOM1FRjKnjRgP3IXzLebDJONj707mNtVIpPvx50dRrszwFuCvOdum
+B40YtRUUWjfp/VJCI7PsTEecV7fPbrtg9AtVr0uuq1sXtntIJtviQvJoImqlNha
YnAUmkTamcoLw6ork4zOedgmrQyjvV37scwThN0396RUmdxLwlNNMTMMoaq+ss6C
Ktelzh8Bd3isrgqeaw2pP+6F35Al4YxAN3HdgdqYIlwKgGYMLmJnSdkP2JGHV0jm
rp7BXN/8De3IUIu71Nf7MSW5W/HhThsHVFv8e0Bb1Y6OaXnH3ion08C7Y2MlXMCK
9iuosvHZqoi5MPLE7hXqqUTrR0Ncq1NgeQMjAIC0uGyX+kEc3qmUeFTpv4Vsxudp
Eir9aSFNYtRWagCqzVmp1nrXXio1nxkV6Xd+b7cDy6l0eq1PxzMTy6y/7vpqOMu2
oAftXqAoTAaUAyNJDK7MfdDg4tWCitxz93Q0oa17ij9+yaHiL4wgadUz8YDmbGP5
iwzLB+8L+t2lSbxp3lzJEsZ59WfYDleK2Km9IE4Cn8DrjU2+kFd01+vvtaMyLrRs
xCCu+bkI3UmuGd06DxxRwtFc1plVR4xBERDak5T+g36J8NG3P05ssUxX2Xss1jWL
U4bAOsJdmTTYMR8TM2ULfbm2A2rDcTCFm03QFcT5r3msoKDNBo+KrxbQqi00ZiXf
EvAcE2QZhd8meNgjW4849w56vOqwZjCbigcsz/TkAElZI3VObr7NSTIDob4niLAz
Ob+S6CTViaMK+I0l+C+wReqPnSjOYQ+ebvYKZ55mBnw8UkyaxhnOC80hajtCGWAa
hEIeJpOnGWrICnY4S3kDPwzZog3OIUsFXw7Ozy11RoF748nT7RAltJLHWkSa8l02
AkWboga/PnJ6oAPWr0oop67PA4SSJC9BhRiBQRac9lLhqKV0oxa54bv+En4LjPMW
TA75+7xQM2gExFsFM9NHVgrTOvJyMhoEHLNwS9gF/uG0QN7E1SbtdMN5X75hjKfD
Gf8bLakhxnPAiciOzlWbO4wA92qu/ZjtQUgHUEU42UVk+WeDXnBAir2lFUKqTidP
aMNpG+1sVjeaPuH6ckkIAmXHE4wdK/UHkvWRZ+xwdMP686wu2lCghqo9nm325F6u
FdhZvWy8vbvOQ/xvrQujIpGcaxdualRO6J39W/kPmCXWKSq0G2vm3S0684zFCV/X
BOt95MhycYsQ+ChL1ZbNDYR7GdziaCrDK9k2w2i56iFU8AGp7T4MFoueyNWA3t0h
64oXrg+fWqCbUQJeDYRZUeQoPiNynuuzvGlWM8ugesRunL92QKknF9PLvwq6Js/v
Mcb3c6UKPxCAAy/3Pw32GjpEkjPwLFw0M6byuB20qBcDLsOzy/tQ5BuZo7oGbxmh
ut+PxYdZaIU4BF+JrGcK+t/0drWVWdhg+zsOLCCDBx1K2Xuh/r5K8wNcg0rjEZYR
3ZlMJEaSZrOkDHmks5zQOCgel0LWYbdFELNh5z5FqIoXcTddRrDn0lm1aFDyRVAA
rsG9G/JUnG+EfCOM7O6NkbvfHAqgH64az05iu4SDV1PxEei79L9ETJWwrnej36Di
4oPzVkYj2DhpbrSwkYeI9ZQnmlgsFoBdkAGSoNaUV8vyfjGLYxCYWYJx1YjrTeYP
8k4STLz7ntNNVNq96SgT83ZLcuU6tBLYV6kuxSEfFLFCohyNHfG5vJ3pTziwGiYb
fPUB3SCFy6fgEe4ggP5/3VXRYWtkRtSXwvDK6gehD78WSrzjMLltOoO/waFsFcoZ
Kgy/Jes/fLIF39BfVDe6VVpia0fYlcpedwUInAocTN7YXw2z43k4vx6SPxDMtt5F
rip2gm+I6NlxyuWemOeqJrABn5jvUdyBm/xKAevQu2XcqmVKBEf7EviRpVjv4FAx
fkPRu2r8bn4OeMd0hzCO/9ZQ7Fnhqw/x7wYXOZWX/Tp4W9XxtJ24YYvqpjbYinPF
jlw69JzyhqFwPGq7wxp3ObyFEQMH6PjKek0RMbd1uzXpJah2yHwDuvckUF2RzLeM
IkNZheD2sSJ1B38nuEQUorzJIuej/Hl8p1f13vGJDkUfsqkggG9HRnFU94yOqtxn
PwnDQ0mTKQkoasStXYwnZzPauo76tTw9ng178WPtUplrhsOEg75NcoqDxCk+z8mZ
xAJWIzGJykJXyZCMRGP+jTuqsy14VUwdzONVmc+jyqhHPGRwKk1BPpRcbTsoonkW
bMfSbBpaDDQ0Szq4JNWbTf6CEoybMNj5J/y9YvpJJrUrEx2x3sbYirAskaGxS984
e83wnXSDZOEx6BiNJG6KAytBa+E0T0Q5yPP+HArWqE+opDPODRMnbzV0sLXx9xpL
XnUKF7chP49+ow/b17Ua2/z+wMUistddXfNi1CzB7Dwq7bm9arRS0/pZIYD8HTK8
jrzEUL4olzQzifjzMcDLNsd3JLyUEGBFrCaJo909idjfFit0dCnuw8FYgSgPvCih
7iaOx4w/9fJXl5C6osUsHEQ4andgkC88w9dNFJEO95sFhVpWYKFH5uV+jy5PNOwz
/QFyJxzFZt5URiee0NPBo6nY2A/mU+gh2C+w1qZdVgeHA59OcPOqq1SbRE16Rj8G
7WUxAZETJzk84sWMzOmmgrFCG+qpAcItVzqSQgk90N2cv3T0I4XHzFhYEN3hng0s
R+Enmgc+9bbPM+sUyb3WK5ecWx4i1t99c9eEZs8QtbM3ceVy8ebdWcqkxOBXyil4
yd8raSxAz8emn5u76/vvLXULYnWi22HTfe8Bj8CnJY0lRAKlJVbIKspoWHUz6pTk
xDgYSv1mqkGTmLUuF2MEEoD5qFRUStklgPIvwSHKeCzfStufy1NOcCw9SSX9MJIP
DdSRoA8tsNUABrdriNnGDKCLxsd7cnAtV/t2qH5wrlm9/9/JfLOjYysxnnYc8S9v
0PVXtJg6wp8gbKp5DhajmQg8y+s1YEeHxpkz9cl9IdxbvrccP+TlX+YuNIyKdLCj
rnZYoP6PxpNB2O1v0gxxIxBoNCIDsBces8ZoHWc5l3uWXyZw5L95imBQ0eFIbQwU
HZA8Oe5IR5nE2YS0XMkT2/Z7vqTc2Pk6loYraLpwVOAiZaCtQDjbxfL7MBlvLt0x
S3nZ7zL3W4VlvX6tk5FRTwXFQTK9ejTOr/liqyaIGzMwzmkacVZ+2egouY/nU59f
kQuJ0oAs3o4OjcGeiZzOAWKUuN/HXOUbkE7nSXcsnrrIQqL0jz2m8iV3g8JNC4pk
jF17+IieSe71jyY9juM2jpek/0wSg50GSKYTDytahJiD86YOy80JkhNbFEhJSswf
7ohEKVERDrTRj6PJ82GucLoe7xVsfDnoQH81ToSh4u3R2yriRN1DMDMDCzWRwXbm
heqBHbeBmGg7fl/RKCUscvY2lsz9Y9hsTaH1QkH3hVo2ygLY6Pcy2c+RcXZCegOc
NVeNYwYTcj7nPeIv31pQwOQaHvTzqslCMvu90olAhAJwNG+GDdaZrzA3BJKCs9WC
lrxAkq/u7rRhtTYUaI8X3tujUgs4wh1MrgGQgOpr6JfXAaw7+TW8rAnelRXe/Hzd
SeHBPC83PhubbBeWzJ6dGSalyPP7r/sS+Eer9mvrjo65l1sceSC42I39OEdxD+fi
JEzqloZm5Rkx5mIcR/7lxHNjIAC1Tb1DLp+MmLHPcsCzUFHMYBcWk/D9M9H5SMFH
5KGcr3f0cLzbJz+xDAogsKF/PeNymwnEIThzSkGA8di0ymx8Gz1hSAF/vd6uNKrR
LOPSG17krRx55uee89C0fk7FJxDcXfZnL3hlZefwaVvuxu2r0AyokmDrqzZHoWOi
T+D/zsJhncIb4Me8n0bUDyH+iTJ0irta5jDvpZw0RIYItdOtcX1nifxFyb+yOahu
Z55uoisAwpFx6Bn1U/TOx0HgPjLVkJBdL+RwQK4fqrULDWVKAqRZf/z6Mh5ePjpc
253huKu13oKhtgcoh3BdFwteIMrDUz6gxhR4Ii+0UQOPW4KwVckWU+mtpHF6ZDFI
NswzOtRq38/HRIyvULmjFiK5PV8BTIpv20ZnG7GMD3+vsdzhvN5T5WBQwRZz4vcS
wb3BgMd0HIM193bRazvpAzhe1m6l8W5GltxvJAfDRSKObNShny+LQcReLTD/NSr9
+BwqFvy45/h8F0Xch0CwDwAv75Z6P/qDKFBRJVryA7Kj+aa7hvrUZuHMgVr9ikzV
4xAz64fPEzQzmtm6s2Y51FjhxJvoe0ZPde1oDR0aZUQ96mzj3GsyFRjvokP652Kl
GZmNhgTOmYGSh/rqMeyyTiwR2xzIbU9Fm/+OeQoy4h8ugWsYtzKqlFcKNcjbFbYG
u54QWTDZiUvFkLmwWiesisRYADlOPEKd6rQ2K/4iwusMEOAfW2khVHh3VxhvXbDN
CglzOLV+EzsDgGkD8wLNiHxH+XeFZObp8ZwO0L2CD+CLxVEYOuJOtZVRuA0bDs/r
SDGUeGVy+7gxEhRimf5YfkveCaV2wmqjqAT7wXpOKi5+ykol2+ToqQIUIhuNjJ2t
c3MFfmpohieogp7idObt39NgRzJ6kExkCKJHYWb2VVCgrD2f3yny/6MzHmaP70K9
alsHy/Z6v3qetEGDK85cscNQswe+xpnifiQyTzDwfDt3Bx+F9gpZTJFjvTBIngHg
Vx2pL8sFSsSHH4U+FnDhuGCfr6T9vAS0DkvL0uXbGF8ScPeZrYzO4MHtXZHKHs4l
OFxiQjz9EXTb4a/beuhwEJxTWTzhNNo8OazG7HgHYh67eCJHO5HzmN4K7K/iWu6n
81kSRAAgfsXJpPpTHG/rv7lz5vGD0ciK+zJ8ADN35+boKuj+pWV1ulRiqVJ2wCV1
rqPA2HMrSj8s4CylZuIaByk18t4NWpJvjCWeeJGnfVj582+qVdKKH0hQ2ll3n3Jj
Ui7EKsiOuCxR8Pv+dx3j1P5LlOreq/D7AsU+96DvwwZ1KRF1GUdq1WBILHghGnuw
22y+Vf+v49GVlspN0ouKa6t8j5LqUJ1MWlC0NWfVTGIipSbw0e1zld1jZiFLxqfy
vBAIpUrb1xeeZM0FrKbZd767HFU0Oz1HTkWAjAafJ3ws5H/W48Nl2c5yscvfn/bN
Kw2jebRKf4mhG68kHCz0+/vaMhvxhxSQVTSfHeQl5qpUJKCsYz8y/o9e/wDE9Ljt
ezjybKtkUvVnryGqsnjcHzeKz/LtU0ghQ2l4h4IJCagTCZqP7J31JD7AqW1gan2a
UNu32gfhu6zVc5y22bNCiydTq2IwRhqALlI3QqzODoQMmFagih7oRrC2E0ZPUgcK
mGZbmwGGfMuK+/JbM2dem8YShlAafu9l/2gB/KtnZvLB459XK0i9NNkFtcImKspO
RUMNNcPJ7p+vnf42gWmcThgCk7uiIzOX37+H0eCCEG1+pQfLcu4O+R6cOZvwU1wd
iEZozKQxVAf8tao18ICiAJLz3vXr/OcfxvHHE2g1hKM9UDSYO/jkialjhmwWP4S7
NU3aLkZYSf0ZsppTX+we0Vf1NUs7jIWRuSpinm1dNiIuju82oPjiOVgruvmpUsFp
N7sNr/GzDTzP3pGQhpJpPDYY+iSGGa22tF/jW1sx0f1C/SatnW2al8GRgBESHADi
sYVY8BxjUVF0OJmojK1IYGIyq/yxdCNsuoPWReUan1T+GxBtryLKu2dvqZYfy2W2
cj1z6dvJYc4SwYIBV8Euu6+Syz31SXSU8ExeN9LC38Iti7Pr8m1uOZ2YREi1pgfc
RDoGpjjTg0t+P/Q9k5SWWTwvlWHaMXwIZOCKS4x/L1lEf4ZN2Mik5s2cIr7MF0kg
FhBUTS7HRy4Jy5Z7jZxkUzItPhbxpH9NuB7kCdP5f53RhLEHZ4aJAPPYWYjTMxFK
QCimKyC2C+bYMYElexZcEEvCgr4aoP3KFtY/1FVX0PoNVPwEZhfrT7b09nmXMRMM
9MkdwHETuidU1oGSLD5syKNwwxwEw71GhHe529UyN+N60vfBIiMZlj66X4mSFLlo
o4n4k8XXDuD8ub3V6n/EdUwwa3EVdiKS579DDTYflZtQg8kx4X27Q1zzn71iU1Hf
KALx+LYgybOSsyJNpVCuVPHn2d4L34Pi9q+/0GIN98W3VebexdvOsJWmrZtL3T6y
0RQJiHFEHnCiJzOI03YIrhq9vnQrTyWKGfCL6B9aTeh8+QCVuhtSHm2p5S2E39EW
2w447XTgCbc9njElZ40AcAwKoeK+X1ji+/Gp64XwSWeaBzdg5/u54PEjfL6OYwKr
OkrCcTZgxXxj1JNdfHQAC5h1LQqFMvfRQLk1ew31gKrGGREsebBrEH+eSGzZMVA2
L9+pSM9IByRc7Heob042a3FRuhVBUIAh6IsLO9wCgGHhNbKj5iXHfD1veyVfYvnt
3bvQre0rr2UU9sMJ+jkkHaHlRBLMvF2FY52jhjsLrvyJpu+9lp7dRrnZCNOI+inS
V35lregx+vK66iT9jc53cBP5AOhnFaVHjWc0vGmKoMnig4kW18ZoQGUOvZX0SpcL
fXae8p3uOHWAWDuwJpLcSTh4aIRGc4chBEHzCkfzSiIWM3JU+1HBqZeuwNstJ+GJ
wwRNzy5pDUS/zdcaHEeuf0GrOmhexXI5ZQdWH3tTTXmENtN5XTpLOzA0boc4ZiRZ
kx+WmyD6TJnKPi9/xV+l72Aj77PMMSfl9T45ib95WRjUzOxKwsQcS1MrN4neR8EZ
HxLcslM7FxXorfwa0FS9XZmbfLLk/KTzAFYS08RydFmSzjTd3wBbepmc5z1qp4ss
bEgT3cVw0jssYHTvM7RpTwCvhBAn9y7XMM6StCPkkoLQpejJk3NcCdBhw89HdXyE
Eu3WryiQ9ObqLvWZwCm4CuDIWt9zxoOgx1otOJnOCTNxST+FXL54SqJsxm/+Shi0
ZJ+X5ZujwD8FlyDNaO1r9cnCmdj1/FKg+aezvhDngDN/ABGpT0gqCLBPDm6+sEFU
st67CG7zqBYbPt8/NPVgOEyXo9i9r0Fd6KH57Smyt/Cx/W4/GWmdpWuJKdeiIUer
PezVErES5/1Y6AsCD1S07bSL4JjxT/pyjjLR5miTRk2e8kMcmWSU7LWQdVmQGWqf
ex9NIctSdft8wKskGbmv7y73OtAyA0704wfKvDJZ4AspNdKoX/M58NL505+pFDLi
D9NxKqoeqwrl528W0ADZWcC/0MUHxFrG9q2E0RcfkH1t/QRfpcGvh4cDWjK0CDNb
x4ChamKd6uSgyog0Q1/k7Y22wlIRWo7aWn2PhHp40zFNUW1YCXLtNfAYpmpetKjf
DAnnUIpmHY2waNBo2iFGxVl62U99ajN6K1lg/AYaAUjiQUoEoQGlDcztFWLwKOvJ
xNDHnH11X8d0pHgb0KcXqOPlivwAbU5D/PMk7GVKK4i6h3ohVUVMVp3mn+8koDGf
+388NIf+FPEFDrg9F/lRtZiXIElNn/Tkj06pU1RifmEjcklnJAjDRj31RfP0uGyd
ZBmhiNI5HM7NSwDlk8pyuy2qzuVVQ6v8Q5DggW4pnkt3AkekRMweUF2b3FQ3SSNs
HHdaIKkayb/IaZxHMhtEwdk3jAjNRWEDRaOFp7SwYWSrV9aLasRpyFxWFUIx/UQx
KyeMi4X+iDsvD/wSgsqkRgYAnBZWeObaRU9KUxutIOXL4uslvcvLWSbbrl8C5den
97b4YeR7BxiJ/I+a+6dsN96kIXxgbsN2ZsGIg4A6miLuNrZURTH/GqyvDzREHWrK
jOZOAvs9F+EBqchPxWvfXu7wPX8fNhUkhZxylZqGCZKnBXGa6ZnY/q+0uo1OgNZ9
AcVGnKiGSIwpzH/pfaC4GWcPGaFrlknCWbUeTJcoL1Ru+dvvIoUa9NbPQlYLctXD
0OzOYDnuv82pdvZNImh1GGx5yygQ5LUpwx6VLVFQifUJmTAPQwlfXPkP/0648cel
Plx86dcdp6Eyjl9uMiLYboU9ldzMMKfoHokU5eIHxcsiB7l33ulFeAHU0z/JlJz/
EmDghx2Fn/ptV8B8hsobOCou2Lyw7tds/n7+Qz/w05V7wtTuV+vj1CdJPWW3Dm1J
pUytTJ5kR/FEm3DOpQ6FketCc+NlX68xaVmCLwJneoi68+wMfKEl2Qtm0WKpQh0G
tVT6ih2VeZOeDIjEfGGhND3CWEvAZf9KKLrS9IaBoLdmKe67SRxsTA8/VdcWsVIx
oCSvAURLBi694AkkAbT4idVx6XEsMw71jTgWHn7Vpab6beN2Bot62tNwLIwQotAl
6vay0QoHviOrTBksVovuQdNyjx+YHZCF4Rphm3B3dexa4FYQxSlLCLuoN8cJxbWl
ulTLGoOJL2wq1QTtA97r/R5LP6ThHeSKvUU3Ql2BJH8k0NtsPR1KRVyoiN4oTr8B
X4z/ogUP9DSeNDrnZzEnjxcX2XD2+LGU0L8vnQBbZQ7lw1lyVfBEkADKLKerUPUS
BNhMnU4J80zZrXx9RgVLcB0d6w8CQgAZq2KvMUPcOqd7KC4xFwpzjL1g7xWb6hkB
Q81j94EXx6aMWW5AK0j0E9JLJYygtaUGJ/+B6mM0DwaWkIzCsL+gf4bkx9eVve5p
Cg7axZTMaxhPnTB1BdefUZnlelaz6azJy4IxhpW7plR/LyLOBgbYCS25dWoivuMj
ViVuyxXTbCCc2yqys84vUdZ9PIiM6QE+FeLLuIn1EoYOJ+cbHZ4jaO9rd4dtE0dZ
h+IwfVcSFx6Ij/qIXc1onCXMM1hW62YS/QKtbuLcSIZcQ5S9WzhOMgeifSqwQmDJ
BECXFdID/2bJ6FgidMkON4/VfLicxevhQXxDVAru70jCJmKRDKZh06xp27CmCv6h
SKIqiS5yefu0WUziT22tecyfjUG99Zbp2x+gRNr/SJ7e5YpBWYlUpFL+f0dryKB7
05Qd3artf/gD516YW+E11R7t/uuce89HSmASd9j5KQHsIZnqTz/nh9BM1ZgIN3BP
/4zALdnf7NhVGhBitER53tXwUkRqQ6JgjSX3uefPwNbeWyr1xi3MoYbw3Ao8vHzw
3cyXl2X9bIe/LhAtVDxrARNIb0i2fUr572q1hQmPjRDkP4ZFszANKp8I9liOM3kk
Mdbz3xc1sv6XcOFwkNJQYgbqeWKMCBTgdZfRBa21DWxapQEqDrUJfdcJ0JOCNXAh
G131p1CoUgCLubC5ewM27Vpna9go/Lb95Pt++OjEfEEVfrkpmyUsjXCSU4BT2r6n
2sCgBfbkct4b8UqzpkLvlFagMepv08XYa13oALUf9m5Gw25CR4vGE37TI1iOyo47
kXETC8JTbwoSGn68dc2AFM4rRyC+f4JRde2lmfpJuZ+zTb6UYPjWYJkPX9o/lyuv
6fx1k0CcgxJvERkpTPduO+I7KwJiBtd+Qf2/2wy9GpafWvRM7OBY3CG76Z+phxbD
RsjkaFWintOV5ZI7zB7sNZ1tD1pNHEviMKd/DdwoPz5bvb9zl/ubXYW5mp9kxMD/
GL2x/bJTkHrwzX+covfUZCllZZraWYquEK85r4/VMKrWu113OAE0AvlZeBLc/YQw
q67VHq8BIQeZFUB1KauMQ9cPxnxXtfEjiOWjDEkaZZFjp/WLXwbmAmD8oBxWipsc
c1iO37ghR9s6JNosglVWJkNsu/UnMtyhX2YwsFJMAgy4LFUdm5yeSwDBd3YwLXpw
f1HE7u7aMJIqRo1xKW9co09JQqgfMslOrnLbTcBPhlh4roggHBKiMuk8eadb+Q2t
Sxim8ut8vRfb+/W6Vetd84DnbcWfxIXdtrRrM9IoEyXuYweZVRSd28Ju0EXE3O7j
gIQAbsvD646FITnbA825LsgRa/cJIaQVrx044K9RebTO4JfBT/mmnGZoBsS4Dl8z
KSHMBvrjCm7ao80FM9cS4+bfLcK++NImb0067kcIHKDhLNvuH5XSu2K3KoAU6e6s
Q/z+K4Zer3xpDBqfafY+detb33pBvPxUWXCAUuR+Z9O07VfvzQHIRa1y273zbg9O
78q8dnw863LzO0UUObnX0vvIv8QAb7fppN9/AxbWJoUBbF54sgNZa7m7A9+M+Ojs
1YgzBBV2yG+C1Y5bbUUeFxKc1k9/DSsv4EUPQZ/5gef4t06582ZtMiR+qUWrvUUP
YP8aWhiTfOsOa+C+uBDDIxkESrnkuJO79BHymQ0lFvw+jrzDdgoChCv//sloLNNI
00mhMYRXzvQkwhFEdBfF/Lo3zyIa86+ic8QgWg0uNp5jZhqEW7og9WZRt0NeN8HY
3t6WX6MTs6Q5pJrTmCcej0YIo8GOPqJPa7dYVXvhggRlV4rFr0BILHm/WMaVnaeD
Jc6FLE9ppG+pJoety1kE2QEVVoy0NzfnrsvTm/N0IhE6BpRjePHDgwZTFvSnJxFj
kOC13nA37r435Kzyz0UKgJfIQKHXQm1bZO4hOQeG0Kv6utKfDBP2pHYxtC0pT8Df
oc/KgrWPiLYUwjALl0W1iYCXF4vL2UyC/lTLvSQjN6oS8AzCtSUzzHm9uV4VeBZx
RNEdYoGJ0CfcHeRtfDmUDajanAvSLvJQYkpXT4rDb/AbNMOuG3Dhtx8N0nrSCX4+
wJ9YJNpMzx8wnGqO4sT/fBWr6XYZlMzCmHsd5vR+MFN33LQMqD6njeQK7DGFHhVL
sSKVbSVDyM8h/4dsSDjDPgxO7ODg54ccRWb9cB4loAvjp3+DF+lqqm7ptEuD5v8a
+0p7hxwSnWMtasvX2CDE8CCdkAGy4e0ojCJGlrmMmUY5zh37ozFI8LuHnHWCqxD/
ySerBVHgMxH1rvfC97mTZt3wu5GVBe6wVJLs5uZebzsDfsXTaXQFPXV66gxLop1l
8MWZ/BL9sqCsUJt+We5RCdDgUp0zli3jswD5h+bUXLFF5vIrwz0MpqVghC+7aT8E
nUB2CWPYRykZVtihE8AP49PIi9BdwEAA8SKon1C1UIJWxRKjBClSAZsn9FYx47ig
iXrDRhmcc790Ms8vWCZiuevHZg2MWlqRIFf8f1ePhSQq8PWbyakxsmtUEPspiFdF
cbo1W6bR3KAyUz88W09EZ63Iu/C5BxvfjWwNYRSrmuNjWTCmJs0RmpUoKsoF/SfH
V07xo+Ot+BhQK4vr80HzbQGgmpLrwBlrfY1OZfsygTfM61if4mx9F8EJUzubeZLS
X7bgKdEUmmUQ0oWo3zbau9q+fkQvJNn50ast6/fiZmhvKfxloMFJQJtLlo4olki3
dQtUxNJztStQgG83e4A8eu4eCL6tHXiN/TGltGajXXME5zxJo+XThQu8PX1J6INm
xCgMeXlOTqFGVjOduXtxwIdFS6KFlJskOUoNfrOTcM0oGPTl1tZIlbvFd6PjIwhV
kUAK7PdP0k7LStUoeC6sEYdmX0aSMpup66Sov5HvBZhypMGo2iqGM4x1qqwhCAFR
6U8AR8/UdBdqgQhf46fFMZ13ckHcSKdKT5Cx9XAP0MSH9xveQS9YmzpfHL5n3Fd6
oW2e68tm40W/rG/MC45WlFKlV/iQUPx7arz5Hr7FGRLkvF5pyh5yv0Fe7KGJ/eQL
5xMTjc4VVVvoyldjiR+p6X4tpRhU9RxKTypcgpwTjVpbNjS/CW7XmScpjOfGEXRM
0dm9gVMJbW9i7bQ7pQIqGruniajFCOSIikmRKpBOx8m2ZcGCoYpQJy5bDFLU6pWv
N8N5vC40wrZS/CfmmFMtrwAIXGZa/3irygf9YI4R4sBXbHomuiJtnO2A5QVV+r4h
r9z9wu3d5dn6xumAbKFtBMenK1dSdF/V2jPgoVWjYETXUX3p8yStVKLeDt6mgaV1
Wtju6Py1ZoaMIwGqabDV8Dsexg7DRUj2fpSGDAu3a6A9VIAnwL5/BhR32erBssrG
PUxYlNyaFURNrYy9RZ3M5Ve6fKfIq1EMefBNx/tbtnD3x0vzwlGOk9nLoDA7Wywm
tl0eDmHAKbSqg9HoSRfIAa24jgn/s2s9eq7hcbwtI4M68vi/Ii7lkzQ0Nmm+1LOO
5HPq4uk/685xjpHbpEQTzua+u1vByUmDD35FdY6iDci+/e4lEr14MTzAY797IFRj
1CeL0Tqn7DpyS3FyiEd9Tf3tkP5VNOOpJ3ZyEdPOVsx/fjzKGvpf8YA8W3RH3/f5
fv7n/8hNYStBOtkux6SaE5/qf1JfnTkfDBKBGEJzjR1Qw2bwecdNVo/jfA3Q2wat
DfHfXCM57heWCQVhwu8VJWJcvHq5cwKwbdaKDDrBznfjOoxFjDE9zgMkygZNHsU1
LsOErSDVxKTRx2akSuF8I9vQ2kVp+uws4RIIQR7iF5enQ16lUy4qUO1ApEMk90nU
MxI4b9I1xSNkzbyufwBmPu40yeDmTk3JnO14AZAHbqFv8wlXnOHBAPCja1Bno/1D
roRfuWXSDbT9j8bWVEFef1TC6ZZzsWSYafDD2bgWMvu7k+TZnBS2sspp/J9IMugb
uQv5TAQvtMY72gq1KgpTKdR+3ZUXoPZErfyM+MF/bc8KLDdM4MP2oAVxWJeWjCK9
VRjAUMt7WQqg8AYc+G2eCNyN0We5hv/jEafYR9XJze6/bm2hBhBUGvHEDxdBC/wI
5Ffhd6rdD7/ejtjF5rtYshNluGfTKqi5aq2ho9MGUhCYN/s/cgVvy1GAN8HMnri6
ouXhqa4BGaolfkP71Ojm8aLbB7pQUr+8AvFhZm/at288RiTVAeqSdN72ZuWxBUEj
lWsoz6gicpimMh7wZOk9K8k1wvObE8vDgF5NeiVv8/9nbUckDksKbD26F3SYOJUZ
SdFhMrJCh2Eb8y3tJ9I74kaKOGmf9YRBbC1+yq7X2mQV2A2o2VJw9X42K/srWxs3
pUVvVWLZ0MRLpVSpIOjp8Ytn9tHjnC7UzNyWqlk8uBIOAUwUlBvK8d2izemL9Y1O
c9rQTyxaOBVAjmLOnMKBxau3PZqWyGoLOVDih8wu9bUY84AfBPiyfhl1npxhy+tr
iaEyNsLYG/v2w/r+3t8QOCJobXTFlOgKFRkPVY4FO6vmL8qNCuCUd8OmZ5J4Zj0c
Oej/ZSFoOQoHLgmZxIx1pZbuJVTO7u8F9ChmbjQXEh/or0j7Rf6eSQhtVbA8tYsA
0AznU++jEd30BoMnArYexWC8Ytlqo2AzZCnBLQou8VWd8DfAWKDzeo8U8JNjuNOk
I9r3IkAKKmymZnWUHafh0zfxlQMxk+u74CsYEP4s33nd9PamolHlbJa78989FuGE
2ThZwRUYzhVGnX0RzupsdKNdILqsSaM+zMNCq4Bc2o2fcRA+rsKhISpYJALRMYEc
o2WiZBX9n/tb3O+A8csjE1tzwcYOC9TM3Bbl+AJ6y+snr/3DIJ/Mj0BmahzFJTlV
KI2NmynatWFC3qTsIz2z23Md1cvnm+2ni4/+3uAlgfTjhNN9UHyGSBfGXUjN67bL
1ewEzi/ywC2A1NGEWQk3Nn/PS9JHUOKKNYRihjMUXZhz1rbsMiQPNKJKvB0lQYje
ApxbiwzwjG4HyjEkNhi4ypQoFr/fh4RT1SRHWHznqh+p6eThnnQ9KWIqgNxSt69/
5w+DITUd7KhYnWrFU/YJa16/P2DR4AsOcmmLPSmsIi0dFkjlmlqzqHYqrUk+bOv+
l0oNOjaFMqqJhUZc1kSFPdWDcQbynlSo6hmg2FAD31DhzXtd78MupssN12SBEgmA
jaOgkg0l5RqQ5fWYwLP/jhbOaRR/xZ0i1xL3aIKGzg9DZwFnGHyxa3ianQzhVtA7
lC2zbOv/osIXqj8HYuzXLVpLA9KCrvfOlCEYFdzhHcOhS2bJXm5Qkwvcxl3Q/Wty
N+252LZ8QeZ9a03V+se85Eo9jgsf519BXD5V1p9hodWgFHKoLf9filux6ca0GWTZ
JRBCR5xNKxhJROrCJAb9CxA+P86PLQNKqRt98x2tkRl61zIx86SfjafBprF5GfQx
LAR8zXjuUa8sE1GeGXVt26otDdI1ciGAcIFk7uVRDotv6q14/B6vk/upFFBYUWFZ
/DC1B21FhDZihmWMpxXcIw8d+adVNVZnfNeTCPklZrSljefsAaODg040FfvN1FkW
Z0/VWA91ga/xBrr7a8xHlthhNHsdgFshCj6i8zyZXEh45oUb6k0TUIImJiJ6nLqn
LrmfSQv75CkfcbIMw0A0QtfTlbPzA/cfwAsLbiBLSaCyRc1OOfQLotka3aaBkqSz
AqwO+DAyja5T+NcT/nvIWCY9oCt1VjvEEpjyJSYlqf4kvRmJidcv9Hz+Yih3COK7
aLdsexeqU28DHks5xvnTL+SbRdPmw65+2pokPo+4fTfammUsp96tCfEAccR2cENT
5xwFYPMT/gDcizxRPqkMYCEEjKWvMr/4xsGTUq4VCeen67ue9T1XeVJy2gGCv/Kg
7N2kSYbATmkqbLdXtqHLmLsOWqKC9yozHT5MEUEJO+3x8FDjBMDUfN7hFvN/wHzj
VVbHLL4gSz1bGzCoZNBnRpP9gTTbDmqIYsfGMZqtEa/wX9/go/D5drNXY9uO/x+8
OuaFMJZdXWmw/Y0QlEdi+UZrZxHds2BOOY1jghOccFEV9Z2lG7AFO795usNz/Oyx
aF470G+Ymm2UtjrRqrDlah+a6rqwKYnc6iUC7HFDAPkL9klTezCH/zZw7SnBagiP
HaBKslYcT/KEVfyDs/lbozlXMz1h4HiTQIp2ADaiZTAQ5RIonP/As3O2EtogRNdZ
r6EY5JMtS5yRMNzK6rnvZahq5Q9eX5YMmhPz5Zs1OYxQAr7D2TLuHku2R4sK3mJ8
kgMSdM7ZRRHijWxxTsVy2jI2IZREydxIaD5/DciKn45yw2pltKvazLw33Mib9EtR
+WJINtJMOxRg41eH1Bj/JLXcg6KAPT3VO/ylyYhOSxQBYV0tsc6IEcXQf9Hj0gXZ
WCkDbRVjYUf8Vr9+F6AZ6CRjr7uRCV+/yabMwtienfcR7jZu1OqYsKBaHmb0FrLk
H+jGuKyzaml1LbAr0Miu+nl/3a/GbWmXJPVcTtmZp9Hrt39nOXGjXO5Jxp2e0qOi
TIvgS+dv28I4QYT75k1KgCiDVFiadH4wrTIpTa/Sl3KbZBBga4n5nkY/4H59pH1t
3d0dwsYk9Pqx4/jQwaalsxZdF2+Lj2b/p+RAg8SlgWAfam72a185vPRuhzZwBcfO
meDQntv5BNSf29Yi7PAwZr0q113K9CJ2E6zSTA8BVCU0E7pkxmmPbkG2m0LTGI9v
PqPS/6NmzjZtJcOr8zc/ytg7jpRM9QJmFNbgMVpLwAC+fLuQleSinL2F6jfs/dvx
pFp3UvOi/VeeunEXrPhxe8XK91P9YyJXd5zdesWwBlaZYWg9WBP7vyDqXoJAMhnM
5wuXKfDZdaQYuLYfhT621Cv/fA82Qx7Li6yg/G7XV195yLTIPdh2v+Lwb7Kosus1
hXOlKRF+fCipAgoyQ83ESFsrdRoT1jTgYaA4zTTnAfC1gbXVYJmFaXDelD8/LHHM
nFtECxk/gpklYQjiJ1xLlDT8FVehDNv05G3Mw/kHWlh97ZyB2dgyzD1xp/bC3dq2
2Ke1LQqb4RXBqaD8tIIW/3arbwRxmkkHizFeFnXUzWLGE1m6KXnxH9/nQ3TDw7aZ
dNIzVsyuMOXVGRLr10lkj64s090hD9Y9vKTfS9O0he4YrkNPzwCv4cizbU5+5p1l
CBVJhjqRw4Gnt//STQ2ekbba97nr1fozFMjqFmFCvZ17cdNuxjpVEe+YqGByOlPD
HC/3uZqkrMnfPxxI/1uR9dANLywM5KBfKqy3TS6cz6CDlshicr7M4A/XA7MjndZa
0JxsuGsV0CZjhrrBoT/lbOuxV3WvoGRHIaJqSG3TCIvqFYLWtOJbtkTXhbB+/nRH
HIrFwheRg1TI5UsmGtwA7XEH6vAAVVODMhT/5+Ut+nhtcVvgtyzUfRc/wvwnHCeD
6u7OGBLSPlBK4QCbVADRSmQiBnNVD+lZbGe/c8AVETp7xqGOtMmEVg8rX10WNxS7
dzw3Z0RtGWZzYx/4UXNVTSLeWVMG4CGR8G+M5sz9YzFpoGufPaw+2oP2aolFIT0d
2uXmAyd1uSxXF1Bs1Z6gxJEDUvc9pH2MPPi44RwPoh2EhY41MQoAyH5DbNXDNj6k
Ui870Fo8ReBZ65haKojAZeLRbkGv8UW0Ua+mSjp7LEdEhka54w7tGimvLDOC2dQv
Xo1KSIVrL/S9X2luIyHRtmdiHt71k8tw7M4+IOHLCDHe8pJcSz0rjXQkk8SyT9ta
WM1LlXouAV5IaF7bNeW98x4gNeQMmnkX95vCmEIBi6UJSN0JqE3Rf4Pzv35I6hQp
q3F/2UrnYG7SBHbPVsqmEQcQGL+tPwEgOwWLK0DoyxTxs/McRXKFehcurW8pi7rv
UqSJpxtF7KYWo9zb+UmIMClCZ8hP5Xx6Q9x2I22GyWumPE8ZWTuGGbRXAOW5SYkq
r8WHnx1jL8N1+61sjRxPdxsWcUOq0OOvUBw2Qq1hd0yWRrHeP3oJlJHqOFSaHGzd
nP8Bh6aH76ckyAr535ckNPHkpN/gj6zUP828Zd9SQe1tsUb47LBXIDGuXLd5oaO4
8XeZ0Ze/ZvaziwdF8DzQD8K4E+40trfbYhWLx8ASJpbcbkOcjN/pds1WWdKOFhZb
0SfgKohBAvmuQZ7b9LqRkySyFnZbsgAzJiTpAU6XVynYDR/WNOvKHs/jnhjI27Ut
aELc0NiZln9Rpq33cTYpWR1MqfAOlvxkWMGKO349V01YHUwQR8c1c/LFNeZO96z8
51Qi3f82q94TZ4SQg/rXi44E7/XeTKMpN5ypgxifsUsWHGpeR6Vtu/z1o2yOqLe4
jMKZpu7Im+O9W+dynx9f+7DEjgujSSSqqQA61yCxak0GdmRfpHAaHABs1vyTaLoj
jYF7SvdTvA8C78md8aexMqHFSeULwitmy7diMXeZdfQ2LWkRqMpaJIRU0C7gBfac
E5UcJQAxOJBZJv4EXHgJuvoXYNnaT6ZZ3trbt7pURhdu3DBxLWfB+qz6M6y1QdIj
Uh8t4mMnfSV52q+qbaAjMiqT7cJh+7ulaJIfvsWdRl+uWiZew+jzZcSavMhhIH2e
aFE9T7Giw32m+9Yvpkdn3oMyNOiSkxqWBQTJ2F5ZuD0DMEfEujehRwhbSHUO/JSm
JZ/Jf90+kSqSas/y1GsFxQ4y9al9n0YO8wWPid3OPICv0vWmpscXm9Hpyu4GZFgo
sixvp06nlXJvWjwsc1rm8mqzMd/BwGecSwgtOZWhgo5d6FE8ua6Fpk0dur814XKG
ZeXvLhdto1n75/ApJR92TynhV+epJvDC8qs5kygF45fK24goreS9qScVGKG19pSQ
DGDvTrdLz/16lsoZpBX8nBPXkuNi1T95tDWSK8m2pWdZ6sfJXmbmG3UY2pOs51bL
o9lniTQnHUlc/lApmhsrMbtyomYkFFAhTYq3JEbU/IfIfkIpWUeyNCkeq6MRh8Ac
1uWuYpjHXVrk8SVRKRrnA1qPjzQSuMVjTNHOe6Io1jU8qQisqeq40NOAgjsZG/zb
PIdXrvHFJ8E/IYJydKmD/J7F1ps3BR8dC/e8cnUfCHUMJvNVI+g10fZCL3uCE/I1
ACuflV8Uqrv6D+UL0B0nugSli8+5FrpNKSMy2LUXhw//+A6qXyBfgh9mUrFUHiLU
ym1msTFz0J/26+0I0K29ig1YZRog/Ul8KjyUPB6x6BCgZHiw0D/BYiXUjtPzxeGQ
3ZoaE5AevpQ5QdhSwsw9ktyZ7uRE53xB3qjQjaprCeYCsGLO9z8nd/sUE4dq3QyG
9bNdgHmWrkY0KAc1Y7Ta+i+BFGV/P2FytFiUiLfibxj7T8SGV8K0z9OI00QtJZKb
7VoChnFkQAK8Q74tfQCMBjabVYEsaFG8RJAa3kFg5oqBHxWCXIHNea7NYKDoqp0b
TnZMwJU5cQAwORqPKdR/NyKs8Cl2kTYknhE8kbvo+t+XHcmqRQNlb/Vcam8/hanx
GLqEanJJJXI2gR8vsgsCJ9gsS5GpAKOsxPFT0wb7Q9qWzsTXsOHTB6w5cunj7zTZ
00ql3XpKTR93kJcwcVtbvX7W8VkYKt6oLPYR8Sy91eOkR2uU+peLFCS1ZbEzl6XT
ycWr+NNEm25Z3C1dh4b5okaLIS3YezNer9mjaNaRyRrpR7wYm5YWZraD/EnKPHpI
wPEHkhsYIQJeCdcloACQI5hOMgN69O+wlfaE/cfuqUIGdxHXrhkk4IzJJZLOTFXQ
zynhadS6odlGLrZ0h9GyA/dF21GnQi3bUChk7nPXc1g+IqqrAtm7flkDos0DmJyD
mALEoM2LKHtTsVNcTyzX37g8pmAiNIG7ci47YItRQfDsGxxQutAacHM6iPmKv3Q2
YFYXEQJkTQ1KmPRqtjQSKI038j9kg0252B2K5ccoOd1ggrKo3kuYqqejWIz9jvm5
OmC+9ugkaQdWSVjU2iI8ZgBxPiMwyjSPSwHrHxHFIZjoxNoEJGRiH/BVLEeBh4PM
62FGi0vOlrH5V2VbEG5pkeWPwdoNgCtki2nUPCVdyViWZq49A/s0IEZX3Pa3ovw8
r3NujzjQhb2gCVaxSffM56iVhqNZkuriNurXMAwoau5JRJezMJnS9mVb6vKd0KWS
2+ku95SDdfShjbCqsJznyEvC0u11toinWFURFRZZ6iYtVzFvjtTLZxs+ee9Eb3Dg
Td5RT7/N4+sOvNwIZl6W79w3u7QXLec+YjpZDH2Jc7mUazl0Qxk6h2GusL5u5YB2
o4EvDdSgVbSSDmdtHL8U432rnhrt9Oqc+QhbluD4jACyiO4SH87T5C6525ftU7bZ
WLBsB6bwbRsGcWt1ZKYVnAT0xTdZ+BilWY50k2O3KG6+EKNT11njHzaFniHcfpQH
iz+3u3tfWQRjqt5Hum6nyjxeBDASCCUIqIA0S138TemrdKuW/h8m0GwQXMAmdk12
yQF48BMhKAIiEmpGIdNKnfFgcLixBM/DKs0E6LHwNMXhF/6CAqZW39tDPcUMIg5X
xiLvVf6EmggV9dHrEQ0SxuGWugLxaruTurCqfU49G4lADpYUUiPregZH8PAbnpu0
viy9I8uz7T4X9E7N0v9kPJV3X+dIlZYGuzeWHkBIluH+PeoJ2Rtyim0/LM5ZZbIO
GAKK71abxnIFMx7k6PlEtqgFelvyxZlwhJkLX1++cbVSelE743MoU6xuy1qQxX75
7Vl3gKi60Dpz/YBPvcSXSd0xTXnxQ6MFwt8GP1xJARNqHnC7RDOorX+PsAqDH2Cx
fwMbkMfG1d5dmobeGMU1q86IwAl6+aEbR8WXn/D0RQH3NGLKMPYkeZAxym1nO5Dc
yknZYCjPDK8Qin7lGvbzhMRli4vu3CFOIgRjkyHGteH/ymJtr6iSdF/8+QDOd482
7JMQIwFZBUN2H1u/7Hs1o4qzILv3HGe6MRDMOdWHbNSyn6w/Gs0PeWzPN4Kz42km
4W/We+RSbAR4JKY9qJyOFMZQe+NAFdPg+AScME6LeHshmO6JMI4PK4ap+dfdXVA8
/d3K0fgbpg0j7l5tnjyGB5zU6gUbB4wCUCCtXXKEuJW+vJRvy4d6vzGLgqLNEwLE
RUcIAKr5zPyyvxWi0RfHAHP32BXpxvV7v41OU4WlBxYb9/Op6B/S5uh3H5eiJDqb
BhdtOa2WviU0MGErCtK1tSAFGdbDbNZwAH5O3Iy7USLPiFVfuUUT5lCqJKet3cHL
cQ9tikxPQgagoKUXQGYvC9JfyfGv39vMrozf3dDywJowa7uHu2drtlECKbw3Q8u+
bfFURP7mBB4yJw+z8kvKuK/4jj4QglJi7is1QdUZxBJLFnp9qrtzvDR1nrVUvo4K
jRqhGzmYr0B3d8ou3CPS/QWx9SOuWDZMkFfFfTLedvPYwQ3nc9CVFZHkfyciqFHC
x7PQOqCgNx4qa8Tbh/BmOaCnQUZL1o0rbWDMSmjCzGhJxvFP0QK5c0tnBzdTnAyz
YDqkW3dCSNVMmzUm0j4y78lupi2KpK4mfcZionOfZv7qb2jBet/ohxCCzFPsCxeC
U3HPE0l6H8MASja4PVhC74wyL4xDzFvJwMYSWxNw9cclzw/te5Z8j9yZrEigY7Ej
6qCTxOOP3gNgbxdUx5ZTCxrvEfgu67eeduxVAGQE+7LQs69jf8xSUZyLWQhBAdYn
Y3p3DajY8U6DKdnfVoyA4NBQNhB8velCK8lyFfJCiAMq4Ok8SuXMsUNkZbAhxvwt
V6+s8fys69ChJY7fIczC8s/8js+k5pyul0DLPMVeZPlfVZX6r5EYHqsZLeDCHnAw
/eijm+7CZwWc1fB5C3Q3Yb8nGN9SZQg/WE3IkMsqvVy/cNZWnxodLif1Z6YTJT0o
JUPSLeBqu5gs1m0igxlrBCtIDd0fporoX4xKq9Fe9/Axm3NmyfB0Bd5PC4yLeHwv
lOd4g+gEFiWO4w3Jzl+/Sglgo8mChVAHppoW0rjRC1cmpLFfDLQU+bQ5+iUSBJqz
U4AIZ7mKiB++fYlDd+Os+G2KqisrcSfIYhLOwPe7iNdmk0C/rgC5s+SsLJL7/8Oc
JPELn6ozzlzv50rWW/QhK8SDNCoqV8cqVvO8L3S7eyf31cng3E8b5bSdPpAt+1+Y
gEuYGEz+aeVROfHy5GobUTtLc+RxALOeczyZwUDQtrgIQp/mC0n0r/kR5HeUQfM+
vB/5UgxvVlmCDv2EjTQGbzKQw6UOCFjWKe1MCNnUliY+l5/jGE4x4rsE9RflxzvY
YycrQqG0gwzF5L8D09iq6heFItvZeKc+oRDV2vQbSV4uZjhp1+Iw6rAqHJU9/ngC
WIJaOOwOtsNulpPwLgl7EPE1Fv0SRudjMpLEdzCSEYm4R0DYdz0RuaCBBTn8/2sN
vcvv/+lIH9Utb0zKdA4B1Ej7utH+I3NGg05m5L2ytZ8scuwfTl59TfIpvH5CVtOy
sqJ+kDcUSmGYzsRT/VeYkoLKcSAFnpfaSAF9C7hDCTC7Btezx/vOuG9kGy143qyW
Un711O48PA+KzkIgsVH3+WpU+PdRyMHf6mrioCsUmhwPcDWZtpa7JbhYk3PS73hg
lpa2mLQyKpgPnLIou7UDhrL6i8kzFwPvq2+kUZZR28VlzZwqK7CB2MqhBFU//vvT
LEdY9wN3GjUjmPP6PMXYEAvWbnxc/PoBoYDsbXSKibNIDZv804++j31V/5sVumbh
FVh7x8gY6aPBjyaIkETtWqR6wDS8jj1/dR69+TO8DEokno9Nj8FY/XcH1teca1cL
ulIOs8Anido638ZsGn0PB1+ABsU3kEKSXP+4t4sFMtYGOx95KKftWIkqoekDWN2q
stmXOKYTg+gagVNzaRNkgNFXg/A/fyb3C9GLT/azszzleyPi6xTBJi51sX48suO/
HJO/A3gx26Fy2qCci5cSAK7Si+gYCBAz64SEGbna9abQGmVGgXBJlU/fmU5BENPH
P88UjD/e0hTc3boTbYpP2tgueg+9Wb+8g3ZAMISuUWewKStk+kog7fGHTP0faySx
S4KeROs3tkXHZWYdwrSMcXTB6u+1SJRptpM5ZTa3SWvZ+3vBKu1hAKyUi1sZ5Wws
sbP3aiA5eXYIx80cI1y8R+dX8X7O2KDTYdaxZfQC7p0kzWlspe51yS8yQ562/M10
Vj7pjuPiF10sPign+iQsIVcx4FNWLz5Uwg1Ol6ENl9IVCVnhR/DMh+IXXwq4YtLb
+FQCC2kC/9cLmkVogmmR725nxbqvEsSQLOTQJ07r1uZXeIV6SO266w3hIaPRQdij
KfgXJdupKFlMX9wND13kxM6XQf6SEd63LilEN+onWRVIOkt3+116iMAV1ctBNDHF
y8kr5T4aId2S8sO799JGa915w4OE9v54m/Z3FYOvgqiHOkQcyLLb8JMUW4CmDiuM
+nrGIv+LNb3v9sL4vY6itNEF5RgsNuB3eNh9d/EgqlFFeO32vcJIBwMOo2CbrDwc
NaruDGOVYypQxy7OOjOKnvPVjnuIwh3vfKauX4e/xO9KK37vhx3CDNaKTKSfE1jr
rlYQfjsrwBV2dFKucXtvGGIgXFz3p0rEB4w0dy3d9vKiL3LJu1A2cMNOI1n0jOPJ
D8R3r5e5e8OZRWXl1JDm0fvAvYmIJzcW+C96SQF8KRR4rpteVUKUMBvfR83Xd/4e
emqXbysrtU/fHHnsM3HHIBMFNGO6OwgQI4SCh4SgiW6KodtahzAO2+X3xBe7TsxZ
sfo/Jyvb1Y/0Sy8WWLFCOSKW5PPQYQQUS6WITHHdTDk4+6VwK3pRwCn/Lp+dFRAm
80L+m4qPqY2MKZypp1h0SxeY1ESE+p6DRQ40Bx9yem993nLwRjA7B+5jUoUG+WJu
BSbHqVtBAVC2y+h6c2BkFW7H9VPZi/kLLSkQyw/WGP5bDLGONGfF+McBPU1AAKTn
XoU23svo4d6Sa7UuaWsVem8zRzJr00vyZ/jMlIGaONr/w3UeVtGGKKnCv4KTF2Ke
BmyJ+h/cylw1Yt51b2vwAwigcB5ZbxLP8FabaHyRfRmzaODD7IsUedoplNtBfqu0
zqVG+l9TjTXtuyJIXkhngg7eXYT1w2SCznvXryQFn0uQUEEEoMLqRjgGldk1r7/g
WOEYesPVOJblnKK9OrnFU0gO0VZwgNRZPstqPXUMbvRInWup9XI+xP/WcJCSk8t2
Qrao74G2fdXMKN9XqA6or0W8bAlUNFz344GSbQ/W4fGfplyZm0NJfM33EyVIzWOU
vDaLSdQMD9az4p+HLbyEAde9KaotAWfduCd7Oy77U6PW9FOm+UBbv+zHn2x2Ptiw
op/9HnsipqCsiJoz+UB1YYn15Kgipm3zaGFTzOcReWW10HAyDe0D3c43hNO/Hlzx
k8N2r5i+od3NlBqyvKJPUV+Lh1AtTK+cZTxxRrMccoyImc0KvIgwq6pFDMrfR06g
sa60y41CmTDH2QdPxmytGblkKosdqIjz7+m6jIbJ9nAJmkCbfEWKuAvp2CxTU6o+
+OcujX1Sp4dkIcqtCHDXZvyUsPBTFX6Sgo7a3vnhhWSIKU9dGknDoSB2kvOo6Kt8
koO58FwWl8XLtOzOnqpt3yHWbBdVxCawSDJm81cH/YdS/ZILsqOiYyxIvQ5f8Caf
Qg/9KOLtC/CqBmmDxDog4AWWghaQ6nvaTgY72JKUFEYgq1Zj6++w/q5Zs02X78ed
oTdY89idHWiwB0smaJePLqvKiy0gPH9mGuu8nqXlETsE52NkUDgLM5sY+r5LBHuz
h8NmXq0x/24K/iRid33w/PSq3w9qIvs0FaphzDvn9hOa8pLK9Nw1CKe/OxxBFoA4
WW6BKNKXQ64seneBgUy77A9NT7J6slD3Vl9v2OS0GAxgCTxwitBl8s8VphLOHG8i
A0C05A9eOPZfHJaqkcFGBvtZ+cXmZoKS6wgOP+wx6uav5pAAlX5EEADOIsC509HM
Z8ILYp4Za0/llfoXmA7OMEtKtP5B0Kncc/YxEjACmPcllJTgZJDsfWKpiFPz3o7Z
qzlST1e5f9dwOEItwnslhWoeuE2pBBBK4PuznkzbOlfL73AmO3X9FQgwdltCtQ1r
A/5RzxmkHW12xegzN7H/e9T3e2cFrtQVDV//rhDzaGYtW48p7HsBK7EbUP++a+EX
fb4RKlrng834xmgfwfCzlIGpoLElsejbsAyI4/GOjJSH3meEg7lhywsMQKmMQWl2
pZ8ElqrtDM1QEDaocc9xZAtsHNBVgWckECU+V9i3przFD6kMB4tMCzlNYy7BTxUI
BRIh4SXnb+fT0jWT/zdo/rRj6HqmEhMuo8SRLaNFfptl/VxlwQn9NNfwYhK76hWf
KdaDpFapc8ZMGwIICSQoDLugJQMvbPesTMEU0G1JkaVs8v01SgT8b1ltq1Ci0R8f
1augY+VS56pXnV5Bt0Vr38ko89UNNmK8mT6QMx93qaDhJRCrPTLBb0L/tLbRZmV0
inlfuaVVqPVYkJ6uD7ZilUJSzBeAN2BaVtxGbvWbUAZIG4iheh4YbJr9ROpqgqfR
edKhAvehcTLUZCEB7oc8kY3v9ft+c+alrFQS1xPeS1Ep5su4cqyao+Fjt6Sh1s1X
aagpBailNeUtbQwi5JQuQi94WzFIXYepUyffBHus/82Bc9yJdyZaIhkDJAagfQBb
C2E9wHULO2IqbStslBb6ccocF9488QAC5GzRKgfcLOjb072TGG6IiKDERiGrrR1V
ReA1qJlpWusCHefP4KcjCNe2mVcUXHokmhGPNc7z84bqzQQUkUZrtUUGYYmDJPpD
maQQCge5M0uofGVKvkRAoqbL7XEYtq778pXMJgKZhsZ4lS/G1przf0/oOISNnPnI
chEkUPkSt+akJTa4G+A9DN1WQbudq/ekK15Bl3rqYdH/D9h44jojB+92azXzRhAl
v3s33ObWPX19FeMtmBpoixutCHz+khEXA0+9dhn0RgwKk1fPOx/fGP1oXX0Odq/6
274BeHtYX2K9DPPkgK6397Ajcd7c5arwVNdxdBwqWRDom0qKnZSnC4jtV5mGMmEq
q6tRtvR1R1abBrIM3XtRFlkcvrlTkE5PUFE8xxktzZkF3+6JRRMEbv21Gekbe5aK
S5p3dsszAktVyw47/Wb4nUw6Qw8mdmaH/OafeBm63ZoUOhjonVLl1GIMVtqNXGkL
sNtiJdO0ngPpJRmvrrL07ejmeiRUftFne2+8u1DfZAgPr32onMpYcQvs6eW4VvcK
wwdpzkh8L11OJzlvjCGHY/LwlUWmTqRUvW3n/gXEh4nkpQTXljypis1k2ouC1AZ6
X+bRorWkPMJcPz5F8nLFHQ4nXiz0gBwixaAIihFbwO8TlP/1GQ9Ps3U5QnUX8HrD
ORynLcPd9NZQAOhcEDk6r4P99y0zD+wpcl1h8XnD+PPJ7kQRYaDrtTYPa2T/Dj2s
eLHWy9GHKAmGqpqnP1+Onc9wSDuXzM6jsl1/im2UiY0/HoQFR+MxB5ZYVole34dj
UKc/DkEVsG7DkdDCVfzCwwhms3tgKQ4NbA5COboeTqaGl8vavKtE6pXdeoqsoCXS
uWHLtcq9E67MhjqxacO6O2eM67hsc0lLNp0sIqwKCJRnwpRtGysrRNDGzKxbBXAg
XrTbAHx5aHeU6NF4Noom7wGZeRaXx0/NEFiau8zKeFGekon2m/kJrg9LDfZMGZ0M
m5wqMV5HNwHP7H4rdxJRml5eHELjTkO3ToSnrhdJOWEcfa944+ZII3Mh5b+nttwe
yvfW5CPLtqIOYJmwwGK0EItHr7HAbrDC7VrRCEb1ucz9kIwGXcm2OWmDOQkd1v9J
y1bB9UGZV09Sz90xrJNvx1AL/fBDYiBT5OXBtKv6IPeHTleu7pzCuC5gH7ppi0nU
a2pihkcI41gmkNAq7aQERFpZ7vnY+GswQATaIopL8kLApfycuE01QX216FpKfvJ5
OgrLmuf5mXjjD4CRH/4gUsgXyzB/oFZ7yHPy5mDzI/DP9V6S5kmeQAwV0euQIlGN
wBYeRM41yKkbqYIxJQNHiOJ4lPTCG5PnEH+0m+evJPalkOfVcQicoD6daMoIqyQT
Z+MIZ0EdAM+bN65L5bHap3kDYdcrKaVU3/MDaO+kUeQVapmbirNP+3fXOt/qFkqF
AAdc8j4O6a/IR/7Sf0onL9t8rXN9uFEaWykJizmAacSpRmr9cXHdD1n5uZ0/bmcK
ESkii0fqtcTbMIauTcNPEc6LtHaly6ViL3ElU5qcuf80+MsH1Ciu55x+3jnLqIW+
lnzXKOI97dgNCVAwisHVsUsokStBhAhh/+47xYNjb9++NTKoYmLOglN4UCLNURJJ
vqPTzOEQzAq/FmR6vaHvNlXqbOLMhwWHa6h/rckslN8dVPg3NpAJIAzJ2YHc6f28
kOkCYF44xKyKYbeEzK5/eujwd0oQ7gs76nAoHwHDi1+fzCYV69UX/UFPkMpYoX5t
4xjPHUhFdW/249fIDq6UmPZoK+B7/MDKp8uP1RElIE9RIjJwrMFrLaa9DgdbFdWp
crbmd0HLtzGGY3Q5xeGBQrxqNj2ut7II1rVwcABI+5547L86p9ncvrp45dsv09Pe
IS/FLmnfb4j8iZZWKBiQlgMfAyhI78pfoc7UNLf09jA1oZXVewOcOTuTnVEAil7Z
VPBsIs2ZUnzLEV+Q1MxW1R55/6oGok98hxBwrbNvwTIUBmGsz2gle5KREgB/86po
Z6vxXrCfeMmvq2kSRaueHBLELEMc6EjHKofdeHCrr2yr/g1xlwVhMpa0mQtm5C7s
Ei4jnu941HTv4Vdgjy7REZ+73s/E2D/phUzF7KwNryIOe14wvyo1fR26MOqr+wSy
FhNIurOD7iFnKW8ehI+QNqHQ8YZ45eaTSHqZBGSuifolsnknQGiFb7b7nvVvOU6I
b6aFSIOivb62SAl/4tQYTycuA23v7RLTvcR0e61qF8vBhbhGbvfj3eNgKQ08ekNE
JFpt+1KF4FwDSMuUlbwgIt6tWQpEACJE3DREFEBNden3+3r/agGZPPmAPZ7LVJdc
510xV7mmIVvjq/8wOKDQY12Sdd5Mj40joMc+IFPPCgARxnJNi/qopEWNP+EAKEnk
imiDvJSUhMnA4xri3WxGEZHTfGs55rPykR/ymKWYisG7z5BEAsa50gy3lJTdmcjQ
z3kKoRGwAIO4pXzTD2EwQ7Id4Wi2p8rr13Ejhc2FFGAH+76BOopd86tVDmXbz3LV
QQCOE6ychiHR7Odvxx7TY2YJHVMTdAlmjRt1EoLLupcoIBm0Q8fx2plS4ZFNsPEc
GxjP+qg+qAp31ilXhRsBfBabX0Ctto/cqFlwAHg5DBSUyzxU7tKsof+xN2+/LhSa
Shu7blOEzfbfsgtEroqW+1ap/ds3MoaB9bx041yn7BZ3w0OB2p/qwBG6arTum6Cs
ALCPSjRsBi4dAdQwP9qzzNJbxZ58jCWJ0sbNq8+jegfAAFQOkw9DmB0gRr1XzCcL
HTS279hHLM+iZH/IDhAQNpcIkaZTpRZwXHALh3mmTrPmxROjZoCk9SvfDLzBmCwB
vlvtgZDqrOmvz8tgjjla0zMUG/pi557/Qc2AYblleIL3pT4W1TMYO5xxFu6Nyev0
/OSXbzuWClww4UHnku7J7gT+CTWZy3v/IwSfQ4bf43q9+D1X/wCQ8p2Zz0gtWR9P
GJYBw7EIie9jpcg0JeZRRmip7XJnfPXgtXBsJRf60XBGKZMgucO/hXpJfI/J43af
AUgxWbnbDH6kWGeCRoe03P9qtV33Jyf8TrqDDyfjSe5EYfChRAgkUoj6yOrKWqK8
wSv4X+/Hlpe+wHFpoSkJtvUJ4NPYltWJ7fkNXpzpD+iYDvqIkUZ/lNXWkAwphk+P
pkY85DpzKEfIAVY35PhMoQDnOPfvT6DcCtjiDN4LH1sMookx4fpJqvEFVBmptSFp
azzK2SMSrPuGqVfMoJK5m+ElzWD4E6wxEKbXS6l4yoVP9KwxWebazBsHCAvSC881
LnAKULTt7Q5irv0K5peqNpWnbku5rzOBD3e6SasK2RbW1hXRK6HZiD1NqFfvByaw
43qpqNjCX+mcB0YJ3Mc3d98MbVvKLijmUzv14yJv8Gtas1RVS3Gw3tloLsTOV3ZR
zkdGk86mLyKreUsAJ+7FiYC71TENnXfYZBqNFcVynlGdF95Tzy6zqsBsViabYmAX
29FEnlLquT9raGooPw8oHiJGh51JTm0LhrUyz0mU/1oO39P4QvHIfR1nRANtLIu9
LwiYXDmonNeT8hzoVwkEBqouqHO1/IP5iDiqUV8HkgZSZcCq8SvKSWown49M6z2q
mze7/o8cRnRZDpFi4nwKBaCP5nE5dIGxB4wO+8cr7TqgQIPrUQJ831o3/PVDJ353
VgwRRhCDrxNfkyMTU5aTzvu7jsljhiGkDwEJdD2NEg7jfJnfPoFQFtVpsPeAz7Gb
qeU/o+PWP8TejET7ZsDfDTA2ic27G007GrB4qkv6KlzKP1gwtLeqruwu1E/53viU
n+w6yZKICj5KWNf8qZs3fIEWD0UqslMBk5kP817kjcT4QBSCGbOSC9a9efRvm5gO
Gq8oVu+QadhE2Akp3EJMPlUTEflaL0tihwOMHyle8TmZxT3S/rRRuoDXDUIAb2AC
HRjRdqEm6cAWUgfMIX0HU4HtyADOWC41JtRKZyPjORr9ZO7ZNC7a46KUGY6Khvip
awPHJ9gSgUY6tECQD2jWoR54ibkwY8nQ5k5pmeauzb/FkOxTgoIJM6k4TZxa5+Za
fIAJ9ORbnX7wNVWko2yqBGlI7olhFLaToD3wpe2XTl6w3jQA4vk0x5mo4b0RQrDM
FKjcx3PNBDTwfg4nRJMnPnaDletyYGnaOSEnjxX061Q4kzPvIJ/AFJdvq8kexKsr
UzyGGYT+aJYuUsMLCL3/CYYPr+vAVtP77ZwELvDYivqO/+zInb+xd0PqM1dsb2h1
bxIoIzDRzMDeETLsMk1ix+ODPe1srTWTCCmz+Wc88fUFUMJvz8r0nLiu4um6hePM
ZQxa16KGGFFA9NsGij6JKGtqBx9a+TPUMCSXYiKXVh2VyPUMkBDrR1ytXZOsn5z0
ak8+qoZf7H/wrMIUQlFQ68PBME7sQVHYRS9O6/PGouQHbdtTbf0uAH2SEnPwA8za
J61QHsilre8Xp37MnpigBSfq4P5CSzKuinRo8pJ5yb7H597EybfPmdmVE3SXffHY
UA983n0zfg7VyEv2or4HwFG4frhp4bNYSBX6DMn3JDGoIurp/akOQbeOeJqP3MNX
ja4lUUvoJrOyM4j/lg6kVJwsPzdzy8NcqX86MuH1DQYH2BD6cJ31tJblZnJCFSpR
JNTMCvx+3OD475Ol3wXG57CUQ1Z8gNjYhorrMfQKXnxkElYXUOP2WkDf/8ExtGhR
hAyPZ0dQLjBJrMJNJoxtRLNyQD1jNdQbEzmgPKj6ZhFfBQsJbrSbSvK2lKcNtASt
o5YxEB5OJA0lAnjowswga6/x47Km/tJF21GyQIelDYcNwvDRmsy3imnAd1VNC+0b
yWReS52mb5aqoeTO1Uv6Kap8PkUYBaKDt+zCswxsKiZEhv1qNilFrxeLYvSBfE2Z
lsizA6Ss9Cb7n8qifS/k6l/++XxVOdnl73FPOGn4ln16VVvwEoMuDTLPL/Ly0tto
tUnMAVYOYexuNJyLWjRogq4I2bxhJzqDIcyKppq2MUhyfVJOY5C0fUdlOTrjaGUV
gdvWtYkjeNNGquOxsWE1oelktwGDobmHQfSrLzQHwqpJK0HqlO7wYWvlbtOyXcna
ECS1gJHec/AJMife4KuAKkwsd2YxQlOd5ubYXy+dhJ7+F7Y11Wwdj7o+bU1MgtNw
WStH4fiW3TgXNBrGjEeyjReh2qysf08Bb/MO1A6JtSgYiqYB+ZUowvjF60PCqmz8
RlMITLxNu/n170+ZAYyfr4N6M4NtbtXIKLFN60kmRFzwjq/HlXI90cFBd1+CgGY7
TMk1KyYjT2/4hrayEZfpUgabZzGDOOxJ1QpGXLT7A1i6I4Ej669WzylabNpVZtfJ
MtLLmkSuOSZgJuMl57cv8YsbzfO0s5xI7u75eHzWXSMnqLqsTVGfMY8bonOt08C5
J5xD1PZz9OQVQb1F3AcqLxvpggHKHmLMykjG8AvtaCuNMAoPXos3xFXHmL7C0LR7
56/4fW4+yJUS8px1zIfz4zWBN0IMt2xggrJgfet9qldQpUdMdAzi2RMBB7gvkB7I
Hi1p9byxFUgpH/oiUSx8rbhuWy4NFPuqMTf/6QSMO5aLIqipA07yozN0iqX1mTcx
h9a/2cPAKU7XGirJd841KaF3eSWexvTQek44/2AQctV2EQX9nFZf7Lcw0nAzpayK
DDKic0SpsKMBtajFw9I375Xv3+bOMePgzzlAeouiqL40ltepIy1u6zMDxi5wRub+
+XzQdMsdSUXCMq8FMBWvy1xkHdRF3d3v5p04Xa2F7//Nvre//XZOtDFlBTZCjAYZ
MJ3QjJvQVe1eAFGW9gKtUM7iXCt2I0+C338iM1TC4DpIpdvEQ2SCsNj3Go131ytd
eYWIkZ2m0bm10s0EJi0Kcc39o0N/KTlcEjMjU11ETPYknhgtXGAsgcUE1nq/yyjh
3WjYzPOwHlTTtc4KeRmcxhwaqkWZ+tNKzMsi7Osne2z37tpuFmf8ECXPqskhBqvS
/yrBulPW2bExGVw9u1p1qLKO6vbp+3aPNyXuK5mwwaCJyb6LFV20GhSS12gD5Pf9
7o33ez5kbhz9Nf4k1CIFvhjANOtexMoccGih00+/tsmwuE5HyXjOOVkBkybV8m2H
SCa9hWaWeNlWriezUPVPPo0TjAsucFsAfUonxHe431bWL5hBIbuKbpv6ob4yUa6Q
Ad7iXvUs9wVgCIrQgz1Bn568Gi9CFCIYGIZZcZHTRMecYxrylZOMovQD+bYEUCA4
24kBAhjjpc3RtyUhG/A3x+9xl8oyVerm1SfwsgrIBELC9kbZY9lSdo3MDSZHGBj2
3j8yWIE3aBXRriQE7CuV4tvNesw6BYXFj54m11+epkuvghIcGbIWzqOvQPBGgA6z
g1eyJeZyBVakmH4qBGThnMZSVjYNj0DzRMGcQUfsrXffq2JJz3w3q+EooAjlghBI
ud48uHc3EPo+S+7EHtI9kDR1SbifY9dN/LF3sYDIvYDXO/6h//qHjxmqsapdG4KV
b3BtjySnW7TcIkaNtpWCC4SuYVxSwcLIhqQ1P0g7mB0HWFN4bPVMs64Q5kwkY9yC
jOUwaCNsg3yN6zwoOjhvMGbvbuDEUfNvzQim5GWYnEwprgowi6K8Bkbnv4nO0GZu
k7+VBlRfigFEMgzocPUNvNzW0N78rfDto40HUiLph5QAqiYhnRcXNnCiLDXVriyG
mjgL4S+N+JHcU3AD38Wras8e6Fl6FeyZVCr0vSL3iW0/uMK7D74ZKocJxRK6W1k0
+4wBiuTvRLXu5+2FMAsZolpbfX0iBKCsMjM7rEqoeebhOv88kZrGggXOisHyRY4k
OmtMBJE6pIui9BwOND2O+aQwi7WZTypl0rqrRMfbZPDd5MTw6th186s/Icxh63Is
33fc/HEkzXou1Ub6IZsqXN9r2JgM0mByeQYq7ZU5k91QHTGQUihcXcqSnlUN7zmy
O+0qaHfI379kIvj3TbSGVq+DUFm8h0ZCavh4Lu+t4XctkxCLZdAregT9sswzIYu9
o895JUonal1R6Sgv19qGfcgbb4ck1JkOWz6PHJiZn1MPjk0juZ+yTkGOs4DysR8s
7IelWaRxasf9qV1iRMHzKc10a1aZyu5bKGkj6jtFgYCPbQ/4blzhHUOnubuMOrVJ
h0X5H47kVrxNA4gLmGpDwvJBCNPlwTeZYoFgJCWF/209Czo7nhJ7TcPqElL3B12a
+6jbdcsKDe54SwR7BK/NmhlK2ujqAZlcFVT6KbKfI80riTqg+tZJZpJZoiLyz7Qg
8fL62ABkuYsWp5GR/D4Wj2dLxioqZ2B2Noj9QPbG1Q+jVDzgE2vPiBACce0qUMJ1
0sD/e8jlvenGQjdiiaexNMI1wHaygOgfxAorP1Y6ERPeG3z/iyL20MII5utna78Q
+CBXJ80QPD6XdNvAqlaSgu+6hiMbb2nk8iFv/PiegfuHZ8dxSjt4E1VNY83sYHRs
nlzdXR9XN9qUnD48suD2x8dANWt6x0ZlbGdXdnjjeKtv+dGaEK8+5f2l31oI3xSq
7KUcSpngDT6J2xBf/iBLri8ySHA++amOda5MOOnmk0lYRXJEWRKJ4utyIctRtK8/
Il33UKQSrSpvFe2AVdH6fObxqXsbGqFiCGCX2a/+jSF84LGuoL0em5M1bGdkel1/
QifvoxNS1iYWwV734GuYIchspJa/fhoHi3AbO1evmeTnhdk+jzyHCM3D98pGcSmO
FEfcKKDH0xWd6IHuBlCxOv5qFSffE9rezkbAQ/7Ise3Ke5mHfimn5gwitlIUJLQN
WCnUZUQzkYJKNnExvHOCrc3NuD7pr7Wc0RybHUqUDIIjErdbZG+cyuvi170j0cmW
qUf3x938DeNF4dMt7htk0vV3ap4GWPTi9t9KfW3DYB7zXEtm6J7vWARcqrb2sFTD
0v6Exrrgcfidou4vcQFH84GJUn1PAkACI35hJsaf6CJmKG9uH8eI1SDRtam09avI
XMDN7KNb5NlQITAIGqgBsTefopjP+rKA62t2mR1x9SkupDlzmm+AvQkm/caCC7oU
qbyX23bnjjP8suBjFWOQR/cQgHM1SOAkJKlICLWJRgyc4ZfHwpuglT1oMCP1NzVf
o+/TQScltsf6QXNqSHI/NaZa9wNGHtwydQno1CEl4wqkQ1Pt6YofArM9KVwnJpqX
i2/EP8pUmmdv8brhtGBtwoJbI/0XhvqwOEiBeJio0wKNOGeN7X3reWOwSOddY7Tb
8ztcP1QtosjydABcu9wnPed6MagnY9dj6BqDlOC4oKQpgyInaNpRegbh/+gJs/Vi
oSf6pxzDjooNwborwwaSz3o34UiokTRGE6Jr+sLrgpjRrivLPSzVexvDEVVcyfz4
+MjFIVjI8x0H25TEDFsolnopyloPhwAeNplBkJcviqjfb8QLBgPrpX/P6IejGBCn
PsgwQKRDoCRoCfgO5ykE+fSmWvv86cGHhpOhgbUsxwzeZsZDhx1tfrtXaaJ1INrO
BzV8rkZE9XcqKQhWDy7SYtol0DpuFCXuXkPLl96K/sUIP2k7qbv95We7RfwYiX+l
LUZgyoLljJYWhe0zg3MxirkZWotQJfu52U+X4ZM9Mc9T0PxYS5IroJpI32yh52FC
mF7MzWajVYdYLAAUXnHJ/HJN2/o5gVVn5ABuSdDzLssjz2r/PXHZ4xyyCLfuy1kR
sNoGSFZa8XSxEwHoBmAvCn7T5XFWjGDavtbkXGH0wI5UQawnbLYl2FNjgjKhaR5O
PzvuyX3pKcfISVq5uM03N/c/9pN2gHT4E8NdoI3aNy1VXwgpHHbIV4RFX4Vkouug
VHDeZWhmmTIlCRo8SahnAkxzx3HXTkl0Hz6M3Q7EcS1mxxE04sKiFTdjJDu081oI
VNduJ/yEPfmsB9OExCbKwj2D9bVZV9lsy23OgImQTEQAyM9QiZ//4d0WZr5wADHL
gKJT4AXcKgvANx8f2ARK+1npdX+2Nr9wATPxDvhQjgrS0e7cUq9xxrBPeTJWYl6N
08FwQO+4m9cTHoaLNcRciLczAGE5WBqdWOt1gSs5NlNh09/CbyE4id2NbwQYEDKt
Fx57lOze1Xt2HCfuXjV9lDducv3j9eXagyGvvKlzUSQXQd6R61C5Emxy8YxFQTgx
BEviJdtP4esm5P6ZffAiU4xqGpuhgT2pY2J5Wib7Xr/Uv9GG/vA/3nY4dREX8XLS
Qut49Ov6RD5eyxamAPNGIL/0RoBPhoGsN6ZvNLYVmPh9gRxexcq50Q8zPVDLwEkc
qCRq0ZZ++OK5+WNOmM1GaUGfRYcUU0sDtpaP1FKQPonTMfDKHM1UpoBLxtLqWTK8
smKQbfOEMrtebBjSloyDiBkWUdGE4vcgud3sXdSSShBEsLXXiVvahlYm4EMXjt2+
t4svFi2bE24DQvUGouhlIWm3eEiDlijjYPu5uMVEg76rKtbSDCExFEkjlge7ae3h
H/0ugN0qRde7cZOS1Q9OYcGWKfbYZ5nqQOo0S1THj6mSFfkPbpCwQ7dNjgNhIwrW
HllU6nVqI30UzoPnGLbGUu2U7FvQqbZeO/9e+2j4tqggYp4qpy3o43bihXKngo6f
gd9WKdxZc32lJm6gZizRu+0gf75NCIvSgc/qGZV06z+ucqkQVPOvevsEohvAGBiK
msrxbUyJ+nqVtvXqoVkeFItYKAF9n6PEBk32K9YhQi0FNHg5SQ9JumuM7p94hYoh
qOUibu8+rU9MwgZaDurNdvQHaKW7ATC9lA6nn8C8JNlXjegQPQUykOet08kAOJCB
ps4wQ8LeQ/k3Xknp3Pb9oHLVWcusmu5RNfKo5J5L9aiRqjvqi5eaInlC2n41cd+X
YJ5ju76btzyckRsStvV5+cl4xXx6+eWNtGS2Ic1MypaftVC84H92+pcjpmK24fu0
Ja45He4zCd1CO7pvviWF64MhwoRAWqwM65t4wQeHkn+IdPiM0MvC6bcEBUGrG5Hg
EO0qINNROc7bwCdl2GQlWLXY1oAFRlQUgCTw4XIeIxUPpW4Qo21UoLqAzZguX49a
Dfus7vPbEj/RuUgVYa9GkbACMHQtTCXJIdz8XPe8Q7GCI+MKCcGUKj7DrB4/8+YV
2dsFGIoM22bS9VO9anSViwgUONaR3+5Yb1XzJyrPIQk3YrOkToUdXa4bF0WOQ28f
pJCf4xIFUMeS2300IrsqLGY/Q4XgovUfIx5KqtkqH2edJlAg2dK7zNIEyymA9CHR
Aro3FUSudvXDl3GGHvWEvZCx8fhUN2jHRCDEKtZUaF0TxD239fOcennGRU7kQxxd
je57wHfQt839rG2kT71+7A2E6daVNSDfUvDyNBXnbpWsQQQmOvOtfUXrkrpHe8MC
IafMF7kpZjW83g2kMAnFZ0me3PyVI2oT6S5pD/b4XYvy4b62gccc1rsmhktn26ON
bk8UT2pteXs+mB86+Tx/YfaK1LvItcUnhn28apvo5Of+NakCNK543nIq2cu3rynp
lBJcTafNPoPMQOxDKeLOLLCeVil9TKqk5fVTVzA0t6Z0eJLxdaYjhA2KkyOjrq2s
w367es/CxJ4x1TVVjkDRhm8WtpqsWBXw/wU/fbqsjPwjNhSKr2VNA8zyeS1/ehM/
NHgW+YHbqd/0++970SDObY5f7Wmo5lEZjhSyU7nzROEEV5ngzx+xO048G9Wn1A90
vtvIPVrScSv0Ca4dIrHaZ0N2wHnEkbW5FxWnL1V/HDHxu+8JtM6TkNsmxAEzfohD
GygJxPxXYq+sd2F7i2a3m54e9i4kQMEiYLXb1Q2aajWusIw7i+q66c4QJI6RW4J9
wPT50SMlNKvnWS0neoK0u1Bj+QZtFc6x2PXF3sNB8W3hEWDM26s0hecRKV/+rprV
MCwgMC+VAeHNn1qe2O+tHOX4n5lWsimqlz5G/tJXWrlt9/KEzqmfAhR86+xLalSo
6tSx6XeMyOXVi+65+UpGITtnvXQKdyjFaSc7QpII54cVO7bR7BtMuozRw3vbwg9D
KWmJUkoKsBy3ZqPuMH5nugCel05nlmz3q75gfdrg6AR7Lod3rK2kIqmmd8CLk19o
aJlEc/TtujrelqYpUdyV6HPHu+QJ7KhNQwDAtIX0kVxAs2qovOB71UsSXYl4yPDb
XfWze0DSa55otlRy0TatgWWbxNNA3kcHjVO8PUYuPyPyJdJUSsRIfJTmEX+YiGBh
ijy5JB7fW7CWLfV1TjYs9yJ83afZBQOuZuZGvqOZVLSN0IhFXP4etSHqZk74gFVu
j9FVxjS3K5V4XvPQQ2Yk2XuZ2J3xJPyayx6ZRCz5kZsqt5isMla0ypIn36v0hiue
tCyF2nye47q/mL8Fj7u73TEcZHdf+oLlONuudq5Y1HftREIkoKVMkZ42FC/KnMW8
LtT4/U0+hIwsGA9CupYr4SFEC6GcaWIZd3ITu+ZPydL6aL08kpg+IQndcmjgSWfB
ms/9DIE2QYsmyRunF9BXrTEcWKexE4EVvE4yRW3mgkvIWMyXbHpDXZZV5U20mYUY
10xz3F86Fee101qacSMiXhW3dlJ7UfrzexcNNAuOC6F6VmuDVSWiQcLmU4qsldGU
45PbXq/tV2Oy0d+nVtEEhW19gbT9/+TNdN9W9ceELXtoVrru4oe9I6WsIGnGnUM0
aHUVxEuOHn/ZzEmAh/tu+tJj9smKQrFHR1h+TPTXWZObTRvBOETKnfTJJn10mmcl
NEQXzgInoKl7DWQ1zNBCArBb1JXHG131wlcHmo2MZj92qDRcCeNSY/Rpwa5bcoLz
0FKOjRjdFnECePoZ50d9VlMimRkFx2JQyQs34Tf6IGmo2wvivy7GTZDBVLFOWjOz
DpuLcMFFPOrC0nb48htNiix60IQvH6l+z0wERlY81s4MSXiBpboGu+2DP/wDSvQr
WtHtQ2x1dWahsTLLT6umb1dkTS5+xU4f1hEvNznrJLMTvima8ok3ycQvmpHzIk9c
tLquwqRjeRQ7oSg83KKOpclgEa5FhJtyFK6HZNRnVDSKuDbTVX8Ip1NZDSPEJ3NR
BgufyOTjC4wpzLQZdr2uzAEslhM+XKIsaqY+Kr9BqDA+M8JGXtvPpSBNy3eRlKkc
SpRlcBxzveTmvcegtHIQS60INeTV0UWhzvofTlVF5NYrXAVMnvt4ZPgohgBxR+gX
iZLMFLxAlmSgF796YjPS195ARmmmsKGTb8gICkG2SQt7FZiz6GSo6mR2ikUURgrw
nm2C44jw5NXHk2ETQrJuKE7c9uqEAuNEcLVcs8/kPL8FlHoiNHzBb2xMrGUg4gwS
0uk0ghNmvzlwQpkMWk958TO4F21b+p1cVLXuM8NjjRVnL5zbtbri704qZBIh33ab
nw72MM4Hx0LnYJrkk6ajG7gzYaIg7Wxk0GNZ8C0j2Qyw/cSMJmgiDTf2BYiFgLqN
bGOjwDX+wZP0hdFfT8Y6/l/lFjP1of4iLp/WD3aR//X3y3V0zExMpxqObf1W8j17
0mSAY18GsIsHo4wl3ogiJiGw9YMuC+daNV5XmqbRFR6AncTRfnCK6AXJ7PaXn/n0
1O7E0OD3gz0DLfRjWOfex+rodkudOBzI4xAmPNb0TtOfcSlvGNxU+DEA94HH5nV8
RzHjcgmWYlmwAc0Ela88K/BEpqSvmAKMLsxdfiuluDKJ4Epg0GOJaY7HYCCesEzy
5ksZnUQTyO9lKfyNg5Bezp2jGnf33csI1+qmziPfjTVOCQ7olGCIv/IXMgT1vx1e
Sgzv70PVlcmfFBE9UH/I2CN6tErBkEBiAYmYTsy+kyilGeY3MJ5by4yBmrJGzXOS
SebITfGKELGBWm+1tyxMx6xDNmxIWewW2DqJMz70SgQ8mEDTGUSATWhUBN2ZzRmN
DwNXJXXovUGsv9KdZ8tsikRnvoM7I7tC8jkzfCQvaHVtdpzJkT5ZOIW5K2g/Pazm
pow0+mJtSqLd89CviDzJlLvFtIfL5BU8QpMxIzWpI1VBKmr2E8IYjMvGSzfDjQwc
O7NbqWZGl54NhFMyDLBKxq2XFDV5b0XyNePA30QxUd939SJM0lWJxg82KIy2z1Pv
BJAFWL7bx07IM1Q4J+vogizzBUF6orJfXfyT/a5yZYBT/+Dl5Kk9z2lfHysJB7Ik
pYaK3huK+hGO2t9uCWd0iB9VIYZudIUhSwRNvkLbmv24O049pAlitzJPR8VJkaKg
ec8I9FuKIzpFXcLbxnUryQgOxxdO2Aeg/KFL59w0D/67vAwOSAGtkGOvAJfQPnQV
lbFwEQjx0MQHXAke5BsWtUmYeBvkOzRyBVPl7x5VY5VrAFOkCOkcYVvMQjZe12R/
cNwezc7vRdCD3pQu5oGOBgsSZal4a/+fK1/Zhd/he9oKUX4p6OY/lmtuT71X8629
xYX5gjUvxndzcbU29ZSpB1taHuhdmChKiURlRP+/V8VZQz9PssgL0rq9w8vK67M3
5ZBZ+ruqq/TZUZniu9m3TlGQysK5EHn5ClrRq8YTmpTxt8riSCHWb3+mMKHf/JJ9
bLMdb2sYsnQJfvEr1XcgYe6yDva6akPGKfS3BArFYLxjClbDnfTzAyYjP31J0TrU
Z2gmHL2TFDIlWxt9xWpdN+c7m9NyEzbNF9EwCP4pWJs9bM9SZ99UvOFjcWHafewC
slvIFNQJ4gja+LOfr1bhGxV0H3kxCKzLGNKMMhB8pks2FaAV2GlmHNxTCFsojenY
ih3XRkvfWkoyKSSUxfzzyPcb/pvaV35EjwpZUyncqdTOo9NsRiI4oupXz4IdBe2v
8Fl1piySn+eWY9BMG+GJh8iFYMktH8woEpZMKm3ut27+utbwYhAd3BA7txrKGU4x
7K2BUV+VZuTp0sr/qYl6WdoGuxeMw+LV7tGaAX2aiLb7UV3nmgUNKRSaFg+YaSBE
oGmMFKIkcGi4Vb1eEpUU4uZBlQ9IfyHj+0ou8ZzpwfANyzxrStAoQYxKiVMUDTDG
Ft+djQIA/i6724l6QZFMpR8UahJ7kt9DOXNwhEg2ncSg3dkWc0hWurF/fniw0wD3
ZFJd9FWMw7+sNn+4auXIOF98leo4he54y7gRhjksl4dBldAWLtfY3UI+vK5RymKm
KWiN2b6rRsn2YYbcyU8+bYEfMa8p+OUtd3T48hOnoaQyzhfHTissqUvh6mmbLwpS
m8eOC7LsrFU0N7tJ54QzjKcT6VfZssDlh9sncVvgGvMP4vzyg9el2A7wUswHfUF3
zavtxWL9MsdBHA9JoNb2QEOP93qS5o5DUo756qUr0nbM1byHsuQiHbbxQ2/Cyjv6
vudo5HrqGRtHLsqXUaH/x+Ju0TuJg6105L7aCIcP8lmZV6A8BgwsmGpWHhmNtu2p
Kp6VnD0De1oyYosWCdcS/en1OvsUSwUQvrhW7YRcrf2PnGgpWaGdrzPoROlftGQ5
1WmFt2RYsYhDtpCsRDnUK3Eup6sUUH3Z9xx3eJTSZCqYMd7SGB8Fa00kWNVkhwlJ
oVrefe5zh0UnU2G6r7VSUASFPwJ/4fQYlWuQApYAAcRwTImk9fFTIwuJLlt/FBTc
dzfQT8W5n51XBex/8jUm+kJ+mnT9wZfW7LpxOD2Jq9wSvaT+Z++asC4NVkPb3scx
gksvcIqqg9lLEmc1Gu3UtjBdo9F76+MxQRm3q+NCwOl7knAFo1D0K/473Bh3aXzg
DX8F4vUEp2BOoVg455Rz5P9oDjFuPF/mqBLHQJDQLBgP70dlsqFWScu4anIpIlY3
i0Xz8XZBLEAys3qqROFzTssFc6UvgAdhKHkZR3MhMYSwAYPsmdwZ3PqjMT6FSPnd
BPCDmDRMwgiIzyOzf6BygYpaUrXma+maZPsdr+ysV0ff9ysdtyxMlAWZhIbrwatS
3OiUGYzIcGyC84pXXQtBHH5jeOauY5jYWXPoHAOWUn+lrxVXqp52EKAmDehzO0tm
QSbUJ9Q1FeLR1ihmwzfDDvgPy7zCo3ZX9LC55223gA+qQMcst3AYnAxABxOEQPlF
cliz5grWvbdql1v0Na+G8k0B3SOVSXE+dQz91EUjatOTI3cFExl+y7AhJWOxTITC
Y8zldSIKvQ0yeZi7p3uvXpoSCPzFgTRugqMpx3bYjWXSs3BMqHHVIpP8jOHgxdB+
mvZFQVOaVe8sOAogXfbAHs3hz7V/DKtScAQsvLFAhS9Ss43bVUR6KlelhNBR3UR0
HI/bDLHqalO/y23ZholKN7t4uwjk/XMjU58uTBPan6XxZB9g5+HYDbM+x6Wsix4k
HPCyuLd6+ZcV/e3OV92jpcTId2BiTzJGXrSEb+zyPOqk1H7gfvqjtropZw/YxtID
bEmaoqOGrlk2pC73RaGyYd9KQ/1hq+QQTNGpGq/uujUov97bfMYMRBD7u3QQcrDM
R7J6450cr6qm3V9MRLQUSo7IHyQqdvQ9tfGezjgTHiI4zGm43VkMf+o7IRt+0IkX
qCZWmUl6Sjrw0e7adHc5I8n5z5OMFwqaAJGbGHusB+/Lb/CdZJrRlcWgbs3LE6KE
sy4BVEjE0+AG04sMjP32Ue19F8kRSBhnSElfQuw9H4mC5vlmNEf80oIjVnzEI4jK
6rfAOUdvnbRd68uNbMnZziYJyXlSmV2S6BJeRiNvZtZE7uam/koj6A41b46ly4A6
EIbujJyqIs49LfGbM3piK5Fv32tt/yiX+oin/vU6cZVHkvpe0IYcLVAUK16smvWE
Dqsvim4Mz6Yqf0dvSGIe/PIekFxdnzAsyw9kz5GZ30Lip7afokmCuDc6Dyh5JllQ
tEpFxFdrx/51J9P/qlkLhonfZ9Yrzwy+VtuGVStt4m4ypr6XAmi22rzoI/tTPmYX
DP5Wz1qR3shCZjBD3mS/vAyWtXmLXSv0J7jXtkMwWWuyedcopbfZMSIeVJ48p4mD
oSaV+vOFovpK2//wPL3+KrWXRTESgCqkAdPGvbQvMGBoQN9ECq11qpqrg9uq/xe2
4b1xKCNsMbem+K+0wVVEEgW0i/qQAlZZis2r/RAOEEVZ0X51aDaNm+5HquXfj2bC
sgI19bh55bust2T2Jj839odLZlE+BgpY/6ner9MWwhzcPFGITY2Z+4mVUMqkSoB4
wTae/NZuqnPj2gh+nvREju1gzI/qifmh0GBLexJnGRe4XkgfGcKeN3CltVp7C24O
8Iq5cFgha8xDPjhqg2oQuBi2vGOlj8sNo1l+NJyX2xly57bw4BtjjQkYfnDAHasn
/9HnerkHlBcWJsUZK5oxNUJ/czUg8RtTukqnofXmffepiWmIw9+sBwGZzOoxze2b
Cahm6FkHC1p1pM6u9uioeDL7/oihqH7hTTlCxE2RBAZsDxV+rUEapgBPDzo6XBIk
q8VbqbTAc3kNNuf7qmS2h01m6zMtVnfN0kA3Ijr7v7WAUEzhh6lfBmC9t1D24Jxm
sH8Y/WrDk5wwJ4cHXqW5VzWwwjS/Ji09HVCFxpEOMFllRzmJ/l8mhiBM84gJ8T3/
tda4f9Yan5gQ13Am0wkJwBEsF8XmISSVyq1NJ9mWtQTWzzmNsdux75FPyNDdCG1F
Atjajmz0eYGI6qcBzmD3qGhwIvXRxJs7sNKIayF/kDZr/WcOozQtHqIPJ6De09K2
2jCr6vy+vWMpmrLQlVwpj31FvnEuOGe7j5cTAE8xp31V/VcfByFRae8jRlY3xNF2
phhZDgeEfcIPUH+Oqj56ymytuBKX4q+7z9CzOrHArQUt+FMM4ZBtq6CXE6wlTqzY
PtX2TNF1nKluHCEEBuOZp6pTzqDB486n6DNnUq+wIHmSQ0A4+CBFDKYqhoRhb/ia
Ed2JXZeTKAMHP0EkcQMHfcwFNXxZko5mPA3dws6ZrTKB1OIbp8TtERKLGG3HfUqy
7POaDyI7soFNRoszY/DGPQLgize1zLrlRnFZM4/bLn1mkya2pJ0IJi7LZHn0Fppu
dqXkPkMSvwmVaisTLKJRrDlOyJN3mVG4jznFzELs2qeLVrEItTLmOPomKB/tG9CG
GI6E4IRlK4kJ4tA2Oe+pTOp1K1DLP8WIGuMzdgdNLzeBL/NX6fQ1mujGYmNF5jU+
dSbzZ5DOZujOihWrue9jGhNF/goIn0U0W9JF1bMTnJN5eyzcV8YTxDP7qsnzanbH
PQN/CQjbqSg/gT2w5qjdl7L9aTxcAEWULC1WMEk2mvPw1pH6inENVnZvaWgd7p/Z
I9uoCa2Oi6ZznN59P8geUYbIhRsnpn5HxRjdo3f9o0mjai0mvS7BpP/2CvlL3D7G
uqISaqVNDwQ+L7OJSUT6EbZTnQS5FE15GI1mmZ8F6fjf27v7Bc0o8UGcmdUx1+dS
1vV6Op02kMWzC/jfxWaJxoU11NAfTjRdBa230tHG4zdstPArqgkxGgSXqvP36ui7
aTxdehl4K+koNd8y64cF0AQNB9FhNFgScQV6OQmdi478d08Rfvp4uqztACELqYfr
IbMYjikvpQYC4+ny5Sf6/TnP0IXikOJhEeIhedx14bdVCVHpSOGodMbdgNiSN1V7
NUAlCeedp7wOP/0BXdo0TBpF3jwjZlM63zvbaeTMDfUlyMmX3T5NA0jZriplPuFT
9+6auDHhQujrWLUQXYqUNDksiX87i/0pwj+kk6AZCP7YUus0scEOuf2G2IUlg+Ji
S7TSwcwafGotilBmhdL9puQ59vmHm6e86+8YyeSUtyzP6M1DjkWk09UrRZmWMwFD
AZea0s9/yxbP/jg0jkJSX+HH5eD+zNAlSb7T63tFe0z3im7fA9M8a8J4OW8/kp8q
WjTP3RRtw/OcrXV6bcvzl17v2orY+byPdS7qEQd6HG9ZUfq6ME40g6QXBXBYH6KD
DC0kZb8O8gUR1mcvHgP9xWx53zRlPmdztPLix7AELDAmes0f9PFH/KvVTFduWLqC
WWCWMsdx1JNq56FQgQ/R9VGV6ukWbBlDmaUF+aye9C5lNN2JtbFDdBKR45DtQ5KQ
RcKE1yAkNROKaeQXlt3BLzjNhfjZMgPrIE7T803oX5R6ORZaay5h8eeKT42hy1CQ
oqHwxO4lViBJuH/My9yxFEyC/EJOWYSVnwe8kHLAnU+L3p+6Su9Eqxt2nRMLrl79
a/u8ZatiuFC7bZ6d0g1ySVMtiLq/nzBuL9whSOatlUMkHRPUHV5pgYqRPbkIYktM
4Wd9V17IoBqujKMw/KaXP/J0kyi9VFks973/AvVtY28f53BLRe29eY8KU8IanQXc
M0EJU/JmRHoAfIahSXKHc2SYfTAuTvf6XDhrNr0CiCmNwYh136IpdUJ9PYckYSiv
aDOBEVUskyiGGoRQ/Y6rTccEl/oxoCjXT9pPUi2X8SklrTthopKP4Kw1H5unnwtt
873mEHLO2Fkov9FTxBzZmOGbzh0TZ402B636BbtHLJWmqN88Fx2fk0PGfgMp+Gqd
+b4XoqjSqcoby/oJXvFJl2L26cBYsK3t2+m+/w2uKx371pIZVGsTEeiO8U53jImt
RXEjClWR8jTlNRXlVn/IvmWM86igIpEIrZw99R+C+fasfQ3HZa46pBW0daarRshv
fqc6DyBCJdGoetFWo+D12sSoP6TUsU4ArRICbjqQ43tBMp7XSA6vcj8p57Dlo88G
RfoKvKooag8IxNJkyfR04dxGezW/0QRAogrkw16/HF7hjyKKFF+kOBJ/iqXMhb0m
IQqzKAjYgMLU72T6fkntvqwd2/fYqH8nGpsWu6TndxqYUU8PNAd7K5ueq+PoqcyB
Ji4fY8ri0YIHaiHBik7gXZINF+db3tL43bYrPrhR9xpLqCbyyUbifRQffSdoXWHr
kBhrSl/c0pg6dFxZwdae+m2MFx/7B86v4oxuy6RkaQ9RMyXc3TzIs8gixk8TcarC
FUylmcukY1QMShDbkm3+W1dzBudbiEfwEBaxNf9u+atoHqty4oNT+RXNWamy1z1+
V/H4rPXfBZVJ4VSkhGU/LF9hpF+eKmINF6EikhbVEo8cmhVDGJ6BJHabdx98Cuxt
YXPSeZiWLwgoa8eJlvRGU18+It90IxDFBvkzdFmg5mDKUfSEKSCcGLy0oY3c2zrC
nFVFEzqZrjq3NhC+bRHRA0INcE4BTbkmHveGDCXEHzbrEvzMDD5hGJHS18LwDjZD
H7cNqDjCOAZot7GMUNtVZy/oBMyc/ToDgmIJaqFwYgYV9w76XL6x3QFWpFWKRFK8
UP4+QW++dK9Y1F/gd2tHab9oc0G0QbWSgXsLZnFPpptA3i7UaUqHbogKIsoYIREb
BnwpRCufzldH73MkHJUEASKgqEeW6ZNR8VNoCkSaBGy7Qs9ALhDCyhEob0+izjlW
ZPHYx3ezO4LXpZD4XN1aJDGzIgcqfC/9h9Ibrnl4HgDZUixEnUURJnA9fw1UwKki
ecJIj05eUYTESU1WHF7O3r45grElIFxjchmyFlaoKZcXKXJ5NDzLBrUUVF+mV5XO
Pg7s+YHQN/ovTTzDVkzy1FTEkN+0EBds7vgAykCcqeNO8Ca1/U4ysWreaGRjJnpH
vcsCYXcsH2dODZpdmmy8Phuy4wjWQt5uUcTcHUHjvDB4GNMKaGH/nGK9gJ4zJ4jj
V1GZjCJlmdCR7QdnwgR32KXvTjUBVgemZmA0Ffv2pmeXU34vccY6TKi/xn3STo1I
991FhlW2OoIrzh0IXzSlSfdU6hF7pi2+g4MEk2xuU+uOJ0jW3+Dheu9oDx8IwAVl
aZBE4Y0CE/Fe8P8Gbh0yfLz68P1VphmVZjsKOtwbtIn3WtkgMt7aaAp/fWqDcV2v
R0LsPXAHoMPGQkNyfRXyJHoMBRFFJUctNmbJo1wQQKcy/UanzNE36BkypB6bh6+s
ppImk6dd8c2UU/1AolVH9mvCe3rvblRAzMRLxx8Xsxu/jsFQW8cjfa7/pDk4Smqv
N/jl5POKS9aX+1C9NOwu+PckOMIuoNdXWf1UhXAFpC1RwTuUnW+UTCBfuih9BnPZ
qaGrF2mv+f+MUMqrzmRVGwNysd26RX6aKWiXgG7gAnN9NU+cTe+axrFObGGIlw9y
OfWL7LrXBHwJ2SBiXhfUhCL5ka9vU+faYEsTeumXfZq5124ewaaBSiEFQ7kRHD5K
07xEZgGQHrRnzCOSzlyku30nx6/EjN0wmbARpxjKNl2oG6R62LRzB5mDldcdb1Vl
4gczaSohqhofChSMW5N1x31mz67UKwNrC9INlChcb8iCrnfmrP/fZ5RrC+QonoTY
pjM/sBwG1r8snAUYSFNnMR6XOm7jGeMLN99qdGmOi1ZiAtR43HezPrh1Ba68PdUa
lVFq9YWRQHvsrHNPiP7+mtPG+6xj0uNYVFR0bw1ZrFKiQPK0wkhiYAfptX06p4kk
yiVMB4TL9IJ8XT0r9pzFQeQzSepFpexks2NhuZE67swqb1npLDznOAW6hZq9/8GG
kQ7qypgmRAOlLJWGaOpv9Hd5QCyTJueCWJd84zFTOPkcHpp81fJRkDH+HKIpMyjE
s8m2fr26CItwkmvOjwZ9ok2UqMVXYgAYfsurqUyPKHTlPGtBARUOyMMbWKjwN+ks
Cej2dlKJ05AkPUNcDrWBOmAMI69mAqYTw3MlYDGy387vMmdpe4GPYx3p3XLo8tls
EJ7gzI8qiaPi8RQ8T86QNoAa6LoYLHh4+5R9UatdhQBFWO6/Yc2cDGzW79DaNqCY
NHaBB2fQjA0DzFHSJDv9fUSM9i40RLloxLK+jORyr6YtD5cG0Ki5eJxbJsAMDiAp
n0GSvjjCOWJKDhfN6z8OjkdW+no6X/kfTt69BhAJhFqNWSfmM4/iBhPlLzYHf55W
80wHR0Gxre6UfrLFg/SbHuYrdIuDi/d+le9CFr5U1SrZeqQzHTtPJwujERSznen4
YkS85a/NtmJlJfw8Tz7CRmJgr2NfDB6nsZ8DGFEocbAOVT5uBKhCTidCb0D6z2RZ
2o+Dh5e77k7EMtv465oXxDwQcxXHt55EuSi77E/onm8+aNWUM3Wu3oLECAiZ0Oey
ksLdzdRRXT5ZJdrOP/WkV1E1at70qhbbrPKFEDjpJvwlviHIdO9d74+2OEj98BzF
0xzqjcn9iP4hsW/j/SbWXNEwyJLKTRyyxLiFlekje3LudFvOQFz9ldPnn30da2mh
qduLnQG30sXmN6FPRXHPbUMaU8ZtdgvW42eCCDtlxkvHK7OlY7ltzos5IUa+SbL5
3J9lThcyL6HfEGEgy34fcAWJvqOHaFzYqKl5h8O7g36bD/oTn1Aa8z+Ig38o+7+n
2MEkaAocDSlewRVhi4zYPEzyM4T2u9cHdnMZenE9UtFNkCZ3QjULhiLJ10OdgEnn
Vcfu+lanIKD0/7w7yfv6m7Z0tIGChY+bdKj4oHTychtcaCQol5bfgD18577dqsa3
3uGF4NIhYs0ylClk0BddGcpSdwWOXJAGUP5EhP+KA5fn4R8VVfaofsMGGjTdT1ay
5EBx4x8iILhfOs0YtXlsuIXeKFr/mPx7gZ5CWuSsRSd/gjFnQ8R1HUSzHsy4VQJP
STzQEiU3d2+XN4xwVGZwx1VZsa0NMjAB+2TrRvaggGgSt3qQ7n3cTsM1UDF21aUT
27RAP+z8TVd18iM2RcNkxlE19wnwrBWZwnLDP0YOckXRiwdmuZKhJ6Mea50x3iE8
7bjbG83mpk8l0Yufl0wU8IokLu/xBIl5324P3a8en/jC8jXgbmEAPjO7TYydZ6xX
5cyzh5IbrIwbzsp6dy8c1x/E5gOwfYN/u5N9o4Wf0TlHF44q4BOx9KmDFJPFOK58
gXFMRXsItgiUdgEGVTXJTlPXKGyi2ZyxAIc6RZGHhdmLMpzoFANyFFbaUujfQaph
AB/OI8syMgEzL5T+pllS8x2oSpZnqzHsMYOPhECPN1NRncjeqv9WJ223mAQElqJb
z01XT72XKQXb8ZZDa6cnEafWBqH0aCAHqSkkPrvg4X1AL8ulsXACzzbVwrCvtKi9
A4P5lFlDoN5joJU3UXqpwzRmflNA9Fwlipg5VH70eSfT5ZGU8zLiKha125F9bJ4a
us8PahF7eO8nk93Qv0EAzh2xmOzPjz226t4/do65M9D62Gg9zU/Vhz7FvIT81gWt
ZIzckqU090iQIa7/n+ZyvSCER9kfCZ0Qa63x7RREUCkTEmIZFmuiho12iW9r6Ux1
OxW5Q+N8bZNsfZBGCgl7tSho43AAGAX+7rk4c60to6uCbT5/Ngy6GuheEfozDe3b
0B9+NpDyXI0wTYceKc3dhHiNo8pfpK6FS/1CQCbiRyhwb48IJdvqtyxXCweYcQMi
1Rs+jAAeu4bjAhYqNE8v+BCe///EIcDsxD0r6OC4fYvG1Kbhsc9h8DJm/DAR0bm0
p9VgRZOiXLGO9J+NBO5U6c1S2p6xxMbu/sLABfBKD5WITkohtU7Ia4yS9ykXeoap
krJsqTi1pL/jxovmhH74WpelPD8k71uSgQ2VLpYIUqf8Z4XDcDNjTYPcHNaYi2RK
pB8h0Xu3PrvtZuZI7fsgLQhu3RM20MYyxEmLe9q1Qk3997/VpOQbLgqEFk0fk/9L
I8+dMpvIwEzmxV5KH5AnIBoZ+ppaTyE6XnKAyedQZcHlX5JPgFT4tT4hufBMPCG4
oaZf61o4lZTMBv7fxmilhgfxeFobXkCndmZ2HvChn6pENGHYn1EdBrhEsLi/Jxwe
WzwmWqC5o/UgjCRM0ySHpeFR0zQORDAo7BmScd3H2wq3THMiZKeVJrL++ljEWnxT
NfoOy5GAuLdk7ji9u+1tihK8ZEAc7JA7mOQhMW6nDUAg33TapGRx6V1A0dfJWlUS
wnRa6O2V3pMAim+B+BU6oKsZyq6n2fgXTpGnSErXCHuTgihuWF+vHtsQL1hCI/bc
dvfGyoJrnn5ruUzHX12uyBZdQJfN4rZKyjq/+FL0asd4geod1LSLnF2amN2W0LvZ
1F9cEJZlqXQdRD0z+8zTrrSXSaK+8usvAZf2hDp5nx5+vG4tgukLsw1FEOyBaMO6
IHN2PgDZ6hdaZNBV8jfZN1Mw7wmfGEj3tWDTNm82E+QMcf+jPJlzZ9MHREU5Vlq3
kBhkq6qX6fSw4fxryJHeETLg2EyKJ8hgnGHyZ9lLrfYUdGa9RfDXCXVGV2kKthaJ
v5d+Vs1WFTRhxW05JqfHsWHrXnGP7bCUNXtAxRj3o/teS5x0L+5VFkoY85WmDvu0
kCjt/CvyyM8lryn2Qfd8UmYe43N0dwBjcnXGWZs6auSR5g1TJqMHjyiyKEuMWTQj
dpdz+ygx4LJKQn4XzszUvcBA+v+eLOqa9FtA8Ypau4/8bgd7eUnAzqvgT8fiu7ap
NvUZX34ESkgs6JS9/Rqxp8SbZ4+5s/9f8XMuPSw3gAki0NxA4TML2VR+YmKVVrhb
yLEyKYJy/FOMGmBUz9r1JdTnLx17ANlqefCiAoMgUB0BnWAJwkCKFxD55AJisV90
63Ubbd3tDt1ObsdZJwPTFo3Ym4hIfMOniOTeaZo7gjHgIpmejDqn9xrbwtpjIdM4
lTc5LNfOogRj+j3OJjyksviDUaoNMiZqtlXRN63UEvG9VYJsrtL2PsXs7oOuw5iB
mkTfLk8P9oYqXkwQudsdjJnxlX34AqjLj6JVByIxXqECpx0qHeMpK/83ch1Zo3ik
kL+iL+BCwx6p74g+TZcligoRd0E73gtszdKqR+WQRxeRLLQC0Mb8WFsORsc3NDgV
OU5TfB1dDwM9AC/PBvVa3N++CHfaIIN/+asU1HCo/0Wvv0FhEL74pdWLHLHm56li
eOnRGIkZN1S6SVYW9IJX5BKJPu1WJpWteLTxfjD3EdUZeK75twRz20pF+AklSADd
RnX6yeP/Ou+0JQ5MvqnqTUME2mlgi/I5GHXugvbfb+slczqOdB/C1jYQ5If1bdc2
J33R94jzWc5ZAJl2RIqyCbj5Y4EYngZT2g2fLzETbWZd6Qvf8ah9siM34pSM9tBO
NWaC5Cg1PD5H9KFiIWxvgcFHvdGMi3lQIT7imKJeluvwFolrKzIwvBDRRlFGsY1Y
dOtqoPMjydpHa9EVpgh/NxY0hvcTQ624V9CQuzlgGsK1CUHcDF6Y2u8bq4Y2GShx
hSPmjWMzYQAP6nce0aZXE2dun5PwoNyBenPis6RKbX3iOsiHxPaCLms7EGP0NCho
YVHIjypnyPQoANiaQ+2mO0FlzW4fO8bJrIAe52U3Z3Ir60JCc3pgro5Ndtr8qpZo
BJso2M8/PsWUjTy42lM+WklVyzr/sopEC1sX/8i3OWDJaXMuPd9tvEEi/GjNx3Wa
g3pkEUb4Un1WVaL7cXQPjDoeyP4R5v7lLraeScJMw1E4yHMkxbdjEUfuHAMYkt0F
zKD99EEvGL4NeEWXnwzUoCGiwBW96QSZNExrGeHVkGh6fqfdAfamaJuWMkw5Gj43
OkKpCFfhblfJ8g4JbwySLemUDfxUulgb2dQ7Ay8W3gzcuy6WmUjz/BmOKfmQIm6A
Fk/QivjocPv97wiz3eT1Sw9ykEIFRXgqLFPomakSe2nuha9Ispzf4YVfCI+h7TBP
riC0HDwj3rC7MUbccxVyVBwbF+MdNUpt6lCYQj3XQuJqFKf5NXfVNdKD49EyohlG
8ekL3QzvmjoVKVAcSABCu53oI1tyqfC2X7RE/LGNNxeYDDpzpW90A6K3MnW4CpRC
I63LaGSWS0lwHKQtRY6Mp6LLw/JNUs8+xvie9EEd5jsMJduZsL2hiZAiEF7+H5Bq
9SrVuq+tL9+kNO7ezLDDYqWNoOC3ZhzwZ6BipFliIo7adE7AvGUhmxkv7XsW4yAf
0kGxY4kaSnnjlR+A9Y+ojSlgV55VyLrnAiYt8nXzDN9VexUeT5RRp0ieKObgymuO
vDRI4qfpUO0N7hbRKFs1EKiM6R/j46SfjffyRZ4tRyg9pxoXw7wCPLx/cPpcebOe
4vkfpmqcw/3EONKOH2u/Wy0ENfi6nu5GZYEZEER2WdmukKzVLiWzBuL0jgaUPvEm
8NHGMsWsrf6pGEVN8/BZyDJk8idtQQfs5IgzamWFA2ZCVJhaYa25v6wzFmLun5w0
ODlCPOCQsmVQ0ncQ/dKjpLe3xkQlHwaf6LBwL6YxXJHc+Ap+vNl2owj7esJJ8FkV
tGWdyDq0imc1qqRN5KB50r+iK9DKcBz0JNYHq/ffuowY+WTotvVD1RGR/EP8o2Ax
WjkWQBqov7etc82Tt9fEMqXvhLsQiq6wZ3aidRHWs16J2Cok0m121YODThou06u6
FTg41gV83byxxYDK0VeZ6GwtDXbWVLhIlCzvSfOnSP+BmnMHW7B4XpO8YIfL8UdU
CnQ6qw2gn3/T4vySvTEOQVUi4/Ymc37UZUZpF3ENiNgCp+uHx9x78UmnOSPkRZM+
JmxA1XzitssQhtdjUQyMzc4ZkRrWmGHAgrdSkIAx6UdlIYn9JMNwtQdh9glnkFhX
q2Q0m6q7V+txtTfjMEuSE9twq/uW7DNONBHDMLlVkDbM6Bm063jUNNyEwh5YpceO
VFtJevZ/M84j6XRAAaAKAfqV9b5oILp1PFkSYR414GryRFoLo1oRQVqw9gaTLsZV
r4FGmSSb7dxATwJh0vZOh+dfXH+nqwiESE5KwIAVMCWaxUFzJRyf4FmFB6EuL+kN
Ork4KnPCqYvI7IiTy2hTu9fKlZXPA+ZWV9/HmSEleIL8k45ExGi1zDlL1p5AcrfA
Xm+jtZqygsBsLrPXmgtLBJ1qz15L6qiz/hgNtG8w4sK/M5GQg3ePekoDv9p+YvE9
qtfFpkLU38w61G6VBe4oWqwOXhjvIHioxNHFdLW61PMzlT2dM0/pleuFVTXJpMDl
qieIwdGAs8eAvwDFYuXgXhJOKl9D4xzx1tXIabSYx2Ur60ty0P+YVEXpj++pxuKh
HkyhgoGrHmB9gCVRbuj5AwfckF1/F/vCMq9Wm4gA6Q/Gj4fgyvWBskLHcvpU6oI2
F6SqqpEx0AKI0wMu2yjI6/Br0gc0C30N4q+qPWI2NliMYRZxgsiGgIZ5ymqhZvga
eT4QPmniPIfWiS+GLbxwCtir1xXebSchmGutYNPDTDA8Vhq+VsyrX8sTF9+BThHH
13Ai/XojfkAmQ8MyvXbk+buA2clmi3bNqyHiVOyO8HKh/tigdgwLgRQVNs2H5itr
dVo0M4r0U9mF4soJDcrENYcZVpOSPNlpRyGZGJb62uvlSWJV+YW/o2HQlApNigoF
SwIwT1IG3Hp/uIt4Fs6V5yHOy6o7Rg4zlDtQpaEOTcLlSjjv71of6v2rhs0Jpai1
u/iMllg17ywkzA2OAh+PPOmbmQOqzpBh3yYneMbBBMVG3p3be7cbjngCsqZ0O9kL
AyW5s2V7PqBwuMdsNdxMeXHszkNE+bdfREAzxc2E+eJMhGq4DBDUeHP9lOxAC/9k
D0Kz5IFg1YM1rMXln+ntbkKpuqpaMuikftQUr1SqXKCx/fET/JBjPNhxvRjTuzfV
0qdCsbJT6SQX9NQWZ1eL6uv4SkRiwm4HU+YGP/NtkknG5cskuHzYUp+wW9Ha5jem
VlBkM6a1Q+UWJSPEY/ClwavKDtq1zj9xfMlAw11/mejACCjYAjNiXc/S/RYe6c2J
PUF2Bl8t/popfmrt3TGpSuqQcYHAkp4WWBmPy51YCB52sygKd4II9wgGxIZXZuqD
6Ja9EuQYTWOBfp+E/y9DQ6ju7eWa5qORe1/WYtf0EO7/+7/n8LrLc8LV3vIg9Lyp
N/16S8oVy1r/feT+n/WgdNbrrKISFa2GRzdipKQn4CQhvyosfFDOkwjqgzUN87t1
6db0M4h6qkv07SiXq0o+YPImJ8Cju2Gce7FPROmLzsIqCccuDFriUXzm68FSP5us
kv6V52VmKVOumB/dxmmq8WM7wJBoqb9Wr22/gIp8Sln0+X+zPjic1Xcfj/ePb+J1
S1FUvt1gBZj7Vc4LMYTwzqr+ohyIuRWyIF1vJlx9j37PwVWIX2lAbZwRzfuWEpI9
8cL9VIEs2f4q/lqS2H+SJ3QD8Zrd98+2QaylU2Yj1+g7j5N6LsOcZEnqzKbQK0jI
2fmsEm05jaB4E3Fk6PN5vi5rNwNmx8+/9fmJaWwkncD/RMO6QH5ZbF65Sz7nR3ly
WEd5ANUsZy2S3pMQT6LLMTVx2CB3lay+F2uUsC7bfD+fd9gN1sqs2zuy96aresna
5jXN6AA0PoOxG9DaT7T8aLKu4u+lPqUmzcCIw9P9FnAzESlFgGIR9z/TcnvL8GTM
xQ2jdP5qdgmVY7L7P2qHYdrpzBgFKKKG8wzZIENY9F3ex9mBslvry8xBzYLSYNQ9
EOn/f/oVoIbGCSZtqbUCFByH0RTJ3d1wEpseCuaqUTZnHQTNfZsC7WdRc0Y3t7/F
rYte00E17Ev+2xVp/mQV8pbFE+e6Fm+rB0Ak2tnqCPwRabtIA+tL1YAGTIG2YGBA
U9O9tzjnu+hiLOC0lB5w4CMTak2IiYJXixElKHFIfcS50KRc6DC4avdQVm4xSnb/
XLlou7MRSfMTJB8DBnCEXN9LT9Ig1huZrKFoJBFsJzs3igodbo4yrkdezuduoSZC
KwzLcYowkJDOWreGkmTHat2oBvyyqCJn1cxLte6W4ULoIYLv6bxqCusrBIPRk/Kl
LCtsm/jJB5njROEJ8Ys5MZm1V51rI0Ph3ysy+Jc1bs1FuzzZ6l7zx235sxEzRX3q
RJ0G0LR5Gb7xvQr0GFZ9qXVVRqlSLIIRi+GAdtZhleOXrctl3fuwq+AU+gCEyLqS
Rau1+OZwIE2mcaX9gqyKABNC33hvZxp20ZA21ml6pN9QhUQPbhG1t+CCmb3R7n1o
ADRpfXmfzfsoko3507ibXEfFEMwYwktwDVaBotIjcSiTLG5YZBTuG3NF+sQ2BUc1
HClG0cKK1hzOhb3seiHOU6LffL/YpniTxlZ8uvRU/e9LznWs9xERd5j7XnPBBq8x
Q3Q7l2Wa8TxIpAXGbCA69bCYt+o8EmAQ2lXaB6V2tae7vQ6nKMa8jeSUwZuHl0KM
zXxC3l03MIgkZPdmTsd0s13XqKAgz0vQpiXlVFjKfLJxJn8KcNibnAZavbxsU7xe
Cyonc/jxokEqyooW1VSOLJxqnK7/Kh9vxRqRntgF0VFNgAraoIRagfJ8uKtgwqOr
d7JhpPyObq5iZM3b02AcVIFDQFT3F2+BtzC2pWY91UwGWSasQU0qdEhq+UJFAASP
b5e/sekW6+kzI9dT5Qvhqrng5atoaMLIxi9dF4W/GAMMkCET+SmCDvJqdx+rHfRY
9Wy5cGOoEEuUl7rXDb9AcGpO5MySClYedIG3GTprMKgOIEDRtBMVRMxaFaJ7PSWW
qJrWB8JkuNOHi74J2lTv89sL9tdTfNFFYM8HeIIRN6UxmGfovLFAuKlj219AquG8
X5DbYWLPjU0ipfw1rCpCYRmdqqB6/2xnBKyMpz0y9ucoYB7l0j4AUSKMLEvi+W+f
N7VCZh8H9cP2WZSOKH0t/77fdkAaKIK1qYC8O7SNimU76SVJgNrSzprMXsehWq0H
f/H71r+vKt9+cz+xwA50rrxYlkNPtTKCZtIo0SMdpSkdJ+mF9WxxQV1Qyo7P9tgz
F6QoEeDlviujr8aHwher8RSIwtMSQyx1IUdqeY8AvqMfTbdg8GP3++yeLqMslYIN
O2j3fNJMYINEd4OGm/bks5CE9ym1HsOlnpE17HkoKbezHbExIvBMcpAVlNHAXV5o
QpwV/cxoiOUS3dturBoS8ll1c/aJ4m52VABwfYCiSRI23xo5KmIaCFTEaTgI/FA9
lppIB86RvuAiauCt3v/jQnVhCT6WuA+rJG12v5avimzr7VxvYpMzCFkU64o0VOZs
uTQ7qEaTLY8Y7fR1GMeHL6ivgksdZX2ihS4P0IRUmV5Q0QC27NF5cy65Bl9WKUeA
1ImS3kYGI92KlzmzuHk0MgJeadhI42OhOovkCu7SEAzT6cFbC/JFYFCqxG26x4yJ
eYw1SnzolBlNF0UDhGn0IU7hxUAEXSXjjqHBKnfGUGy8GdJoJMz9CLXFCAeg7YiC
kNUWnjV0DQDU7epXKbJBel777alsjhXgUznZhIp9/Ndqf359PaEk10WK2GzbOgX6
FQi5eGQ6QPd9QIU/k0ErKrhk31vic9yPNvbbYOKwk2LzA9o/1qvulLbBkRsKk/FJ
yT/76/AvOD9igkSvHCWCYclYCsKDN3H7g8xWuf/guKHRHkErUVC8MGhvs4YilHpW
eY59xUVSk7MGwCKQyovvv9u24s4yXsaBk0ZdswqKZ9E9lgHJ1gAzGzf7QLoiRDgS
nFqR+ZZbJGKL+HgkTxL8w8Sa7mZUjesuFR0Siqs4juTojzmSR45GThPyf5QIyNMJ
PSv9lgU1wJ77ABYPZhvYXCYfqDpjAfBW+pgUWKyCJ4INikpAwuKlZkAiDW8+3CQ0
jMrIg1t66hnrsHjU+7wIWGCVXQUKL1rdLUY0ExRu696dq3jAHPaD8Fe4vBVJY15+
aGT2+bq4xxD4/SIz3OBg2kxr1BxCTI6zg9GALBge/+j6a3k7KhJYkFLa96gYvCow
1zVmkR3jJgYI13c9NzOTL/kHUmZ0ZcVuR50YTz54uBkQVJo674wkxRh8rhcWA1tY
HYeL+7SnJAn6j1xrQdjTssMctdx5lUkF4e+KoP5ZVnLy3QlgQeoI+Dk1Y5lquMB9
7F90pkaWFUBbEud3l3Yyre6YyoKSzf5vy/IaB0qyJnAG+T3yvNVxB4MdMWuCcyVh
oYOqeN2ZpUcrCEt1vMVdnqryQ665VmCEB+N9iMCbdHmZOo2JvqXZ8eEaw50FxY9i
bMYQFEF01ere8Ub1S5xe9m3M8iYZ0Plyr4+HH5m9lE8Ex0fYKK7h7+306ZdwBV1x
STFEUekzqYej4+QX5s1QIEHurf855JZafDIco4T15W2KJ4VIetomiMQhZOXNDG0n
jV3PWIM8m3DvNnrjGxafAl2n5SlFFG5TtYwSLHqTL0ef/q4NUKiN3kxe1eRDRyt4
SQCGsiu8KDW03Ed+5d1fQwZLYzKt2021n7YcVRZA+GtwHZ5MEMgVrUkAiAI1axID
9e6x/iG130fY17gF/cky75iYRKow6MZxS6FNPJ0wqznoxjmS8zHxRqLKUbyaRTcr
VxHilYgxDjAlsLLKFFag4qszB6gfWKn7xpk3M4xGOF47ZeBkIpIuO7wYkIJXQqrg
ik8j50a6VwDUZsOePYj8pT6Bm1ZgrW5cYtMdR6ipa/lkq5H0sR4uAxnJdTyO0+9t
KjP9xHUNIwcc3BDaTXhuMX7bTHWj3oB3NH+iXfBY1Fgk3b0gpflMgojqorJ4RJ8C
fu58nGmjOdnCnA+PMxEc43OWLCP66btwQFNZHHC7isL47JzUSTxhxxUDROAbRFvg
S3Jfb8eZG/MvfV5m1TiLx0awYuZoepYHtEbyY+Jy1qkuMYqRydccXydW1L4GSLAi
1vDCrQWKQu3oMeYs4odwRdbQlMXjvD366foImT4TXh8Gi20w4ZsjmftWMT1zWjtx
UG+bD2BWbZ7TkiGsbQ2870RvBTPjlvINIqQKljebIHJwJP2HFaun+vmsLfiX5CQq
bEmqvFsSa+6Y/eH74928Lu3fjm5TkrI96WDhRQF3uXAmLWVk0NfTj4jc8ANp17eq
nSc7VZe0mAY9JOnKRKY6l/FNydNBqZH2Mut6QEUWQKFkN89gXKun1gFBZeoxY5zZ
OKd5sx0ahRECCcvYdAPokw6E8Yxv616fp3iDX6NnlWat2yqdeMyEe8ZFKYwCp+dW
Px0PSv1tUeP9qrGgN+ry9SQhGyKVTR8VpxGpxXv09xN5Ep3KmAtVvNLqGPoyaAuR
O2M7n4UQGzjQpXKKx8mz8EsTHl3qaXYTVKByPKGUG7RQY3RmSe+f+F/h7OTACCcx
7FYPG1+7qMZhr2+khZrPzk4Ly1iWUPM80XzgzgfDIw8Vo4J9VHfByKAqalb5Dj2C
5z0b3kIM6HaPB+P2j+NRCs/1lsynDl++doPWOEWR2sg2M81EhmBDSihd9CntS1v9
VOQnIlOrHwOyLz5pd4Mzb6Bt/00gtq74QlZ8oQflYWjCB4FwWiUP4Q+cgLpBOJiL
XtsXHmJGyNk/kfPZlx5JWwMYWlbVp3/HHDlswfLTuOSJcUiyWdeKu+11DL+yiNzb
dlXdjHAc0BUb0GxyXWDAbPiZ9EWvxPuUzMiNXpX5+Hc7hQZEFcvN+n4hHk0Ybdsq
GUwL/VBdYgk2OOGeauCnxlfrldLHab2Fl0mB0xAXt5yAPSM7c+J9BIUqgnNgRcPk
Rsh1EUHT2TcQGGqacNd+/fLsw97lz6xGvA6en2TCbLQR5UtGzIaY0mX0UK3rbOy3
AKHJLLnN3vcUf2p0u6cEbVdQOe/9wNNkCcdJ6P3M6i/s0ifJwSVlbAsd09rSqFJm
EVxRSir0wwXbSCe95S0lD5Cu7thaHWxFKUgpyo/ClAnmp7R6hQkpm9+/G4rvEymd
KerFTNRFlWAqRQkDs7thgHNMoVIALn6olmYSDDY23kOhxvClroiPXfOk9LmUcyNU
wwxaUYCOmYBCgAEGgJ7hh29IvZo3mlSSuXjfX/EUh+V2xtjoilwfEt4IMlH1Y7P2
gkZqoIXkntk7iyrijuBiOzVTGzR2E4xBAnQMrrzXWI4YRaa2NX03gwQANc8ZY9lK
VNwFYyjskYFvcf/2PF6eRtIAbvYh2ae1TlIWk2Dzii3kg5fUx9ho09GTzcmM+htc
eljFSm1ULtgARiJpXiz31b4zcyUQ21e4BfaEe0hbMBcZzBui2CnBtGfExm6C3wsR
EmDzNcYFxo8WylX6phvSQDWSOQqrLmNAVbcDii4Y+LuHGiyyiK/BI83xbH4jPG2j
sluQ94AiUUQpnoCTzo1uQjsjt7pLZY9ePL+h1xtao9973nxiuX/UIz2qwHGx6Tj0
jNZKrUoMb2Lnedm3Vt6LNqpYJVakVTSyyYs22OfMxR3baWfYo0fF8Ny48BzBDfte
R2PN70vZTJU0HTUpWY5YzG1rHovU74Tq9Q3RxFqJDcHYC2lUY0d62qzZACUdChnJ
JHAjBFIuSkxuZo7ETu7QBrfgosSVh58ZemTieE36xnw9BjZLnOX7tpZcKi1YEIF7
17i6EC010h1IUwN0xEsZR2oqWSvG6IOCXn9F2CdTvokwf1Fkf04GZMjmDXOIbrkm
0jwtcJUuFyjAyI+1QcGOiyYjMrBwyIVLkSqTDR9e2I76x5ytEM171oFKFnsqsgVK
JpBRNVCVk620ZxLRDQkOp2snk7icF9n6TbjIv4Uxd5Cw5X4JLBgmSVkW6I7c6jz5
8uLpuqsMBzpG8aE1PwJvru9L1GTN+Gzs5zMBlug5LswbnLywkl7e00BcF3s1w0gx
dIIkMSXX9S/30u7U0Cb8ni+RKvX9tUwBtfwwnhyJeVseNQo3l7PIfQuZKm/+BAjU
Uw2/rWys+SQGzqWdi9M/t03RVsn/AymSuasB1cyGJbLwQ8x4CWDscY+FTiKdEnsF
hxge30x78BNewAqXtVjmuftO4792QUBfv+y6Co0AtLeOk9Z3cB7L6vRRAFFeZ3qc
xJfATFV+kdlLg65kozHWj27+fyCw+7S6Ydp9uzuXps/hmmcj/uYnSUw4bWMhRrtE
mSNFH8CZ9y/96m4wInJvVJ5DvdFwvrYoOg1PgES7ipH1/P6vcpxQI+3FzWWFsGW0
Rb3LiFVMelJYRYDZAfTnWD5K3FEPaIND8BAnSIGFl4Snu+4TW6qZqvS7esnQ/A+P
WQKR9IFW9+ZQkddBBb88el3+TrqjXUiJe4WgMFnuAOTRtaFcaLeR6keal129hY1U
XEuVYUhM/PIUEXqfKqAVfw3ZCOIQvROT/OY+E1y4J/TDCAidieJfuMnxkm4wDR/Z
cEbkaz4x+IY3wpcJ5ldwkZBuXYEabcdqyAHYWQhWFYeixB3kQUA3u0c0Ce+wbDMv
+IDJwwdkwOwAe4odslRYoI2w781ccwFMOZe7rOKezjrTWSDXTQbn0nNrpjPkfyv0
sN5sEAjLJzneIuqVJPBJw1tGxwlASVe1r8piq3ccJlhh1k5mWKQmfLYj7ZDVk+8X
ntHNW0mdbQgjOHVsdUlJtUHqmeMZzqFStxXpsbHH1kfAxaft90XSkpui1Pq4vd7G
EV7nl/Lvgzg+V7RqfxFlfSKIKIADHJoahK3jG/3nj4AjAiEDCsjDEWwe07wA2SRF
q4pFVHsoWHRy/kY7T6zUfznr09Yw9Jx/VRGV58Uj6HW+fxqxKo3rJJqMPGy4e67S
jPBeRjwyUfJu7MxYDf9oC/5pgIpCa4JLI344pnQuncXYihUZVBm59WdiRX/AvIgM
MEtvwER/3OSXvnbhmolivLYkJPInI/CMDyloYXStdWNn7TQjNzYsGPRCpksZS6JA
m2/DYptgzaF8dgg1kexbduDMkIBIG2kklHVhf/w+ao5SsqXJTZjkgEl+O8xkXnex
3RhT4pnYOoodPTe2gFbKnU+P+1EGBYRHmE84JilY6HQomvanPT9cw3Qg/3+gvOJH
Bmt7F0gBpCeGs7IQ9vGJeqr0VxHasnnc1qpcNt7nKA1fy64LP6fF3OmnlHrkK4TE
sK8TIdn31jcdBBXN46VlcObrxQjn9O2wwMgXdyVk4jUVGosuSmU8b/upnhoahMop
9bXqxCxOKC4fGcz9ujZ52TVZWWWHbjVefpHbEUnPfauR1CRzJcIkj4XmuLeJqVcr
Zh7pngEOoNwDb+lLFCcess8gHwXeFNn0uar59IulmVfX9hlGWyNxvrd2+M4DdLXr
fvaGqn7dNEnXhaQyYSb5xszMwN5oMsuf5fleSTSc6mGTMH4TLat9hr0uTRusE4PM
IW3TFwtjSAhFtCxjPdvG2QnXp4fNREs8Kpm2hhixyE/POyUKta18adDOWmXqJ/Dg
z4M9pN8Z/inMCoXbLIeAbJhjYyGHe4OfyZgv/GBIYf1BmR9BhY7h66BQFVdD1uWY
9Z9wbyPaeMjuu4HLgkVCdjYmRgWyNPVmFyGwDiLR0QrmQbm6zwnXSIT/u8hlOLuf
hnldf2qPAx60G1Fxnu4CASyLNaJk0y0jVqeecHvOZyBWThlj4rPryvT+bhc6sBVs
O4IM2BGJffXwFc9i8KYPONyct2iLFPVJv+m4oeUjUxZFs8g6QC1Fhp08YoWN6Lje
bdB+bOnXD+EAmoK6dNH+ViXARu+/J3Ph2bHGCauHJ4vEMhylODn3bNi4yPypFeEN
6tb6h5efEZyJp44kgBB+mg6PoFo8IJdlENdS3ZVWP7ZPWUDepnMC7GF7hxJVMNwG
uEgSeNHtzBvrbJCej4sDZS4obr+Sik3rmPT8D1Z4DxpExXivp7bVvRKiYp2x9ZC9
iZosS3USBDw0ykjuWmAoMWfAo9heq9N1tYqW481oJl356H3dApD4GZuzWnQvfPsM
yfvOSJ9e0gX2bK8BVoPccafJW7mdd2BhCnHxK3B9UwdPw1E3J2UrpVGNxEVhM0UP
0mzytOirM3s0sMY8UThkvGlx/5pTMK+3vxBocPSz29rs60JYqvr5ty/m74OpiWE3
lPUo+AAI6mbOiT1/Y+4U6MhXlbrqPk0sRWwkOlRhsJSm3Xf+rCaREPhpyNwZffG5
SMjE0bAV/RBxS+kTIEPQSpSFjBAX7sv03kXtKkTH0Xpoicrq1V37h7vBw1YCXe5J
xA4GldVhMmoauGT4NeT5XXVZVVyvieru8kC5YfDd7q8q0Xky1T15AV5+noYZt5py
Dlb0Ghcc4B8RUlFzWEp2wMYbeg3uNuUsG4yed/zt8I9HX2MHmt7fQRMXfkSA8pNj
sGz3Bhn5MS8XeRxDx9d7G4XtPK69r6KQ37wA+RvCWeoMlz7q7XtEA8saD7DO+yem
EG4lteDn8do6PHNVZNdCARul153DHCYypv8SfhtJ1yXv15A3D7bHh1Z4iphyGshf
FaVKnUqBSxsGSPTU+i5+cTmF2nSA/8HPQTlX9lSEvUL1Q+Ry6MCs181MGfExIf42
Jsmyfig13k1CX6bHIxS/bDXdPieR4CsXz302axP+kpee8iQqqCijznWvTV37susc
v+ZPj3RSlBxVVlW/GD9BU1FEn3wfmjIw2qKtUqoUaAFQRr/+C0anN0DOPGEC7Ma+
unjp8Mb61kDuA2HldbHqT03a0jp2F+67vEcH2O75FmhylXXLQX7iX+M2dWp8Pc9D
nUsXUF6Pmt0BsEMbWBSC9AFrwQT8b7+czePeHAYRFP2n6jsfI2hkxziKoMgoHHgf
gxa3xGetruq+/xUosVyUNrLKFfUw9VwCdg1+IjykhzDUSjJj68Vl/Ib/LCk7I+Uy
4HZrt1r1ps+7WLuZ9Lv39+kMdhX8VVU79CgH+KxrikBWFYCQYP+pBjNQdD14jVet
WOA1QCYZacmEkl4NLy404ZsMLLnScEaN8OOo1MS9RIDBo7/6GCwXdgLlIkOHssQ9
UXoc9T3dmc+PXbngCFo+HTVpqPr0RUSvCX9uIEvmpq1GykuZ3yGCHsPIuEMTuRkK
nmcYEE4RjQwmF38TOJf8Rr3dv6IFHKIQQXxGYpGWwp6HnzhD9B7JDs6hkk+qCwj9
pPl7cDiVoDC8+OYLGSJtlDkXiJsw5YilJGyvpe++FLQUapDfevjMUga+qRMmWGgK
V+VZ0bWTtn9MjKItZy9Q7xFVIey8tmx5tCO55O7VF/dgVE0UuAz0BIP6FoH9PLkW
VwCCFLaq6CSeUfJrYNpRvFL2TS44q/xBVHW1aglSxSvA0OtTq8/Gx8rfzTixBdNp
AFGIIjAmQpZw6VtfB7O+aZk1cfhaSlIRF/2t+q/coT0QYw9IqgdqRkn/aiVogw2R
u+Xj5dG96E1fK9w5JyORIYzVZlXymzKXNp2gL+Yfb7xMgj8SkvdLKlrru+/50TXW
tmSWAoYCk7PDpVbMrAJA0Djitxx02d2cY232vox8gO49fY4dLlyMSW9NYuFpzRlN
psW4QHNFV0mHSgKdY2QxTWsXmocpYsTbs7v9yGjbYSkgJGoz/TViDXJboBBT0rTG
sYmV45W3nxYyFC8sHExdYNM43YRD8Df4EYWC6QNRqO/dLmhHe0ubGNRdAIL5++1z
UaZ26A6AKq7bAE6Tga5S0z66SGnrGb8gVvZooKT38jd/48A1lI6ohGluqGTGe6iu
zy9T6T7wWQdHTlZziJhzCpKOwhuqZWc6trp+kSVXB334mDYFRB/Z5H8wk+qKsg51
dVJKXMOOfoeefILys4+ZCwN3Rk2vppuOQngDl/NqYaV/OMB47h3cF5HGry966t2h
XTVv1hIq9JEY0m12F6EsaeoGb8hT3kNhdPkRLg6zYUshXTXE5A+HJKYnkcKam59T
guprXFiVI7/foCmyFolOweZyCo5or9MgVIIjAAjUq4iNktdSTzmHjt2QZabV5wXJ
FjILWdxeSEzdpS8QmrH/y73oCpcgisPMmYC7flo7FhE2pJSdwbIW1ahSaUO5xpP2
/fzPfmoWwFR3nka8UWQVCT4xXavPG+aXBaGvMxR/RApC9AQ7v8DpnNfG1eqmAPwh
hq6VOJsNjVnC/DOmqyJaJlASWnngPpev2tkUF56ZSqwQmDPst4NhnUBti8p7WYdy
8OT5H/QSWgv/6QoF9uNV144br9T08VN1UcOJg+ngVkt679RcQWRvrClNH7gzs1yk
fuiTLrsetvuDAvAaRaaO+cfRsnIkcfSX9YXnAP7BHsfJjK6IneOe50xeS0DlTFLE
kKc1GLNrJli/pesD54UhhkN8MSZwuGWHCEpdj9ASxO1qQnBpDUyajPk6L82J4P6W
XJePwHBNbovpSK2CkM5bGcEDnRfuK2SuJX7ER4NiVT9mcqbtSl4l6w2NkJ6A5peB
4l5I9AN9Zwq44LEI68WZp+TLreIfGMYYW537ck67h5QKTXamUNAwqg+THSqX/22e
PyqBhJzs3VoqU3E/0HBnFguZ5GL4ZX/O66aI5OFiamyM0b3zyI8hJEDsjUiGnh1R
usNaYpov95d1crkE2/rFrUp52nsty4as0egFXBVGSb1vNGDvFyUBRwSq3nX27gO9
nJiZvlYsbSegOilqvoGbhiVUsfy+oFuY5KKWbxP+ih5X7+9AJPQvEzl8BrX3kjDn
OeS0dm5xTBIa2DcX/FVxjqA2V0d/xcXDtrGNE0+fAvYuGBc+rOUK7t5nFjK4SGAR
4seg4BsJY61OKI638GCs6y2KT+wS4tV2nV/hhAjnrdPjnpqDheQ69pOqEd11+yau
9psesKE69vezuSzj0gPjij6RtZ9RsCNV6KKYnsxjb10KmU4vlf1GXT5IWG5/iIRv
+UpmRtfn8gh69DnaIQTg7DeMu9bZGig/urLAJu8MpAu3K7J362ELG9zKhPfJr/ym
TKtQsqH7UsF8yPHIbA+XL4BLRvYNba3OhouU2ndKNIY5ibbwy164O/la7n1GF8kB
Pmh0v0SVMjtaOpwEAWna0TOkPyeaA1HHO3hftw6VRKdqE9znSE83rKkf440EbLJN
75aJJnYVUx67yG+Cu0wVga7I7p3sAoEqLHKMpvPq8/wtsa3+TBfx0Xfi01R2vNFV
TBxrNlvlQanKxDakBoWT4IyM407tEeJTBxVGOMrW/YgLJPGxkcb5dlR4Ru2wUQqq
jA53IG1rKosyiizPQC1e5ogsGu/RBjLrGa9aTgP/JvGmVYD4SZWeNRdlqYlI4geu
X5LZcKikcLbKKx47GWrQ8I2RFOV53kofIK5OTdECG2RIedgieVHfV+G5XT1/kX/W
Akw4fTBGM+XU7Jj0q+FPHJ4iwpVB9J4dfs/QbkkBDUffx7gATTRZGDJHCzPCoG2j
r//MONRs06c+dcGsAhRb+lekFbjPvDFkeLAsre33GIiMlUJH/a3Z9m1XGMXpPRDu
F/odyKv8r7helIHkpaIj4Ov92dBolvTWtITI7oWtHH/tIvtj9gh3qRNu8S1XRRcB
cH312ivArsl42UMJyVgy5g5WRPhfT29ITdRplbmq3z+Bxm4MzYlEM3mzyPE8DjRv
mmdo3/BIHM0OWTcCeEcklUWRBuy7QuA1pXX/N4ADE9x7Q7uSsqws8ng/wOkndxx9
D3ZoXqFEGy1A1bbjh0MjfIU26ZfldSDefwXLYuKC7A0quIw1leyPtNCUzhMxvOQv
1VXN+m/LlU23LGPR+SAtjaP+LMlhUggOSOu4sMxrKAlkMfrBXkasjVKBBhQkoKrQ
PcBohgyQKAFM6gr3jjKAodfXfyc4SMJcMAvVhl9FcFuijqfUqKoqeZQHnV+47HHh
4XnZyczBH/0Fkmm4/WERQjMWmSyVCI555oxN0fwuinLQbouh4hdmuT5JeaHvsEhz
7zaEw/9p0QULDzSOE8a5xF8Kx0zqPp+HGG3E9huw9cT2zD6O9VRgjCs1CdLGUe4P
JKdTtF/oMgJlnRkIf3AqpRvEJ6XadFlQuQxv9d+CJQbXv4i0aIDsP+z0sQgW2vIe
vOcY2c2zrFsHltRh+zlrgjMHxzFBqvhhcvGx/RfAuYFIjAZBQUavBRwyR3pCakvN
S1fo/yGaVgwuvodp1MxgLRhN8dfKjCo1I5spot3men42eyLHzdAPy0aRP2DCsBrL
YAAlsrJOMwTnRSvxjNUaFcF62tK/hr8XQ6EDretLPqMa2FHQFLnNn1biNE9q0UcZ
sgnc9Y9O8q9fexXeI6svfmgWlNTj6Gy4xhmD5pjfPRevUbW0H4ZNapP7R2LUOTmI
m9+WNlsaez7Kw3otiyA5L8CrT3hjQbVMscui7Q4sp31TRAV6qWjnFTuESUECkuGY
+Et+4F/02G71wJgH0D6EYaOFySQTMv19A1iuvm74kIT1lD/O1FV8Uc7ZKuFuQyYG
PNye6rh4KFAY8wNC8u8x+7YVT+IP3+t5vb8PU/nniAgIFIL8nYimAV0BWQ8g+gXq
Yu9tGqrOsCTqz/FgMTgOEYuBkReqPWJ0hvfhkIzWukWDr/pUaClaxWQ6IkNI6B1E
vUEH8z6hMGU2iajFAhYAR0/UZqwzYVW5AiPYmTNd+DhAnzFStBIlANYYtomP9wHR
70W1UY+owE+g47aDz+Jy1J7nYLr/sFK2GeZp6P+6iGWWOIf9RrAmgI4byndJqHqF
HfU6uyoyj2iIf1jR1mqwnUdxnzESq8BkQlJYAY3uW6X4q8LIbCZ0LfXq7jyPlqjr
gQwXuwXUnsiTnpiRY6djRSO3Wgb1qQdp+DMzVo7aZ0vgNcnh5Vwdd9ucFhngIzbp
/DmjKFVwVal848kpOKISkdYOunjlDQsSfqRBpy8Vs+dUIOhmQoSpRnGwlZFhWq+f
nizU69O0qetYDmK2Sslij1a2Fa6IDeIaZweiP04YnELHhOHsuAEqgvu9gmQUwszN
R/A1wPc6Yn5t4jZDzxanc/lxUkqCa6ONy7U5AVB5Its1q0syFPyCVqUBemDS394P
EJb61AAJZqtY5HcAsD1t5fGjE6tlHzXkXHXFXjQZ60kqWnRqloi0JVbuAZpC9GQW
MNaqZ17zTVIwYruEA1SBlWV28a+GfqgJVEO3+1/oqRdHzZkFvL0uC6KEKQ5kixzn
KQ0ecsKUV5w0m8pOwALDPOiVQPgMSpWUlUtalFY0/mp4Tb3TYrhtKpNFrAaYME/G
u44SjScEQl/1ldLsG5iPy+kJdz7NsXtGwRi2CPv8AbSiRvmd4rMKXp5Wmdsqgs/p
lxbO4euGEKgqhV9KRhF1VbVr4Ctp28WHdtKsM3fMFdJNkCDzYt3bOPPCJqRSyw9I
fJaArL+AiMT3dcb1Ifu5xERdYTyW+lIMbPUcaTGCJINZULr8N7TqRIQYRgBHw8mn
aJuihIzDO7FF73bTpEhcCzayHpQtd8wIsMDBtk10QqXyhQzk4cEkObxNry4M3Roa
QN+WyMsNLBuCi4uNteUSsfRRSynlv5h1grwH6CizNoR4Q8tSwNlYCbs1OhZzFHHf
Q0cbQQt9ido3rD9cUO52O86BkUKTO+LoxKEaxZfm6A0f29Y1YCE+g1lMzLe2Drv3
gqEZwWVSYOpLg5uGLoAZ8evafvhf9oTMppVEs6ZbdwiGqu2L3btW4rzthx/Qdrwp
mJOOudFJ9ltEsFH+uMgQzhLT2Fs3vny1ojbYD03b4/YgXJWcNeMVvGbjpIHonzrG
p1tjLJugE8xQ9lHFF/4iu/cee2rSLg5/CEagSQ4An0FU1+0nwd4iGIbnBNjilNRT
KCE8chk9oF80sO+CDq0eYjFesXHBaKhJEi+rOSrx3gECvllzWMhi5ncjQ7+dO/1X
uEQ49FKaOtr0ZA8053HPzVyTX+ebgNyuX5dFjLS0Cl2W3EMKkZCL/xqddKETNBKH
qYgbQBJz2Ohev5D7INsGT9RqRXFXxETEHYkvrghAJBJ74obVN0Ru7wra4zmkpksg
P62RfYcPpqk9bXRC+l4a0qSVLfFmA8vNWpyYTwUGeVmIO0h9kWULuTvpza4MvdAx
sYHrBEvm3ZyXWseNtr4Vi02Hz44BFk1hF+PSo+xhnPqfys2kvftWhs1cDxtvIYa3
DkGKa3F6tTfeVlX3EtZw0fww4abMvnCS9nMQj39x/UmSxeUrMAAbAeucsSaGfZzp
aUruPYZu7j1zCgOK7V9QMtoB6U6tqEaDexrzgHx35/pE+mji9Z5CZsS/fwU+NfZv
6FJpqgk7XbQ3bCY7lZr9qHg1gFjdyM5bxSwY9EHX2iln4vuy9ZBFMkzQVc3LooT5
LWBJSVANEtK10qP8gLIMqp5R7e4jniwRZyo7cMvgX/2mxlZCBUKoD+6fRYqWHWrJ
gAalb/hChxvzfhtuY2O36Q2XhCAV9JGA8NOj6UAW9O45IEd2KJCd7lde2JA+GJ4F
nb0M+yoZ0Dg9BI9k4mkCl+SIRbH4SGM4rErsnNHVfVxsbWiejZh9+5b8zqiEicbK
j9nISritxVHJx10qTDm9243xKQB7JtONtXj88Sd874PRMvifWzJwzcpLZpKDxjw8
V9Bmt8nsPbFytfS0/Tfn4tsxlYhR3eF6lYE095mCUJDowSqg+8SWNgGkz/1CS95Y
IEE4J9yx9qHYVXQ9e33imYWB0peupdZ6Yad0SyeOFoNeGifaangPNMwcL+b8FKND
muT1k5+mKhda6fuY1BE6BjL76+sJLnnYk9Ynq+vULddJ04EX1MKIm4P4f6g8Q91Y
hWdXoRkuzfKpBVjR3cOiZ8uvK+rCfPiIJ7f7Dst4NEihnIyikQJnCqUb9PDP3HdJ
1wNT+I77H9dAYWV79TTiRLnJpqFsSsBrqqV/2903qXmPvc3MuajgnSFWAlklLJwa
mgNIfftYaiK9zxBpJdmtXXxMPNWNnOXdjptt75ijeWdZq6OOWbcDA7rxHMPowram
QHMiijoFaooZlc6fScrLTNK2UntGaRsfyRFyy3s1EBd1mjQnfNEtDOCEDTL/KkEv
Vy6fmY9PEu4YjVkJxRHGruXCqpxSd7NdmxeLu7n7sRiqRQNzNsguh16glfudF705
q9GI0P4oVcUvxGmfWRAWb8ra2ru076yRTDqQHs+VHTEzatM9WOTDaA5qD9VsLe0O
g9wbt27BFlKqjVJGE0Cdfy/aKwPck7MamQhoBfLZSUTj9gnN8hLZyXk2sP5iQghA
6EgJIYdXe7bTJM9mLph1CfhBF6XYUcumuoX69YcLTUP1vU+RyEEyQaWzO2eP3eu0
SiX1TNz/1HyJHt4gEO76+cGy3/89jtB+Xn7VgvRCCAM+r4jwP2e0/ohNsoP6aoCQ
NFUz7xSk5OamI04TXQyWw86KmIboyBstMU9ns2tgGb9TbOybiXwpzHAY4+QxIb8X
RCFSZN4XI2UGhFXKqPFhZPewxikFAzdWvNzhe0lrGhTlyAPYPgsvLtwQe3ucefkT
azNRqKYC+PMu+BWIcrY0GKPyr/bypezr+QRwoC0jJ2VSbsWyulPWpVcO02L5TfZe
PSdPWCtiGz4PXnlBuX+B/A4RLPkQDDEJeJqfjW/0f31AvprJovNCvMm4WTtv1RIf
crWSzhmp6GkebMhEOzy0cGs85YR/B9G0tC4uAv/+/KAvm5MDYf04l3gNxbsOLCuW
DGh299OCZP4i3p5kHB2tyOlNluF4+yB8tfNXGVASCdRjhnuhjOuCjhN/ld4/U9G7
OUQJiGwg79zt3nmXemoH0OlxXzPcKe3W799DgNBuC0yFaMlDgyeMcU6QOwpWtZmk
AlMmmlEzUq2wBbzEtUOpVWl7eMeLe8L8V0XkodXbLRcGFLLXjUol9PtMNbeqQihN
5p7hr0caGS5PRtjNuqvY+0bQL3eaCp8ngz7XMtccDMGmqg1s5OIWFA0rKT+ab3wi
ZwUAY3vDf2YzdcumyIZb4gywpvVmI/8wEx8eIRFJ+vLbJbTphBMjXUFYfQYBU+yr
rdc/amnHEnuv2v6GkQBWAwpi8qNet73ECQcZQDLIXrtlGwThCR+Uz3QMLdttP5+k
4rfyfdbsA04ZVr/88Y0eFOl4XG/1z3wqt0rrMolwAPwtIqazLQ86bD2uTpVTozmh
A44V8oMTSUpk27UADV0I5m3+qBOJ5pmkvLsYcSLURCEz6okxyp6MVO3XFdS4wnTA
+FRNQQOcnERmS0F9P+CJVmL1xVhPPtLyn0uFgfO595drsOo70Rdo5VA81rVTt7ra
qBndrRVsR8vkW/S/jeEAUGOKCCnYUrCF7z3sNOI641zsPJRst9Wl431gRtVGqyzI
YfRqRqaZpyzzJjzRNm6FTkl0/3+A4FHaHWEf9iGMwA5nExlgvlRJzxfIJA3T3yrk
7ZUkhSgOVzg2bgzWXVF83uU5LmjNp2hEIKw7YKhoQ5j9RXmC6QGlMuyEynB2nQze
T+Nz5vXqznFFAS6kUf337BO3BWQTkwwKVtkljFTOTNOvSclWvj6UNxbnbkVsxoFa
o0Bwyp2MVzTcLFGNBvV0HXqZIIAcUXv4mrFfcRF6/qka3MW2DmoxInGhcqEYT1DV
dnsP8jTYxJp0j5GQ8SmcqT99nD4Me/K2N+p9pNudwrERKSBkch0lxx7LEr7IwTiS
J+jg/gTy09k5qgV2/iE27A07VJifhJq6NC6c6Qk15rnKCtxr/SI6wD7LLW9AUuD9
cmg5UscBcyugaoqyXlyjFLrxsz8jMDbNSC1HHli41ikTsajEwzzGab8fYI2arj+S
B00b+Jo2uYMARCWzsoaWgiekxWcaOOkMG+YUmS5KH/dh16dtiMXYwbMD+FPEG424
fhKRL/uWimuCGZ0ggaffIDIm2GEvkVdhZaGlETgtMDV8FHO5B7nDcmRojmbieWfV
ZtEAWIpuEYkrOMz/kscFmJw8CT1HzdnidDXOBRi8zUY+ijAl738SjtPxgiksSk1M
fh3X/Vj0ZsNCH3zFiYuzaQRBGk/cqcVePLb67pfSZ/Dm4jZ1dZYc6GMNpwjnNIMy
UBvfpgeCjRDgCNEmIengdJZXxxYuGtuZzsXi1joZ09G3FRfDDxSLRGVI34iFQHTM
rAbYdPd6+qN3DZm/kUZOkLpt3i7a73uKD2E2ZrJs3fgcev/BE7lC1tADYqh7zuIp
tpjpF/FySt9LZQ4OE4xUsC8wmehSbCRxkacjNSAo/pbrx4IG5butnvMvAa0TNZlR
GmPOpa/p6dDuM/jP/ZVYmawmtDaGLpWWi/OYX6rZMoHLq6NnEcQMFWFGFVpVdzX+
P3RTCdkDPT+2JtbXvd/pQsL7u8kiq3XJzh/W4+zdpBgqD9P+VUch2FEuoKUKI6LW
H0+vKBXhnw07lp84F1dmmUXzw5H0SEzRy7dB7Zeh0q5Xhq+4mUb99/EedblmGAwg
rqAWNmpewWziyQrvaTnCDJvKrFtiSsf+DyfhuP6XQccy697inVuYjH7TSAF/uoYh
1ZdCb1yD50fyRnRvMxf1HJUVs1rGmQ75aAtCtPYPzLgvsqUpoNCFNYV2jusO7ttJ
JQZsxoqWqoRik1F3ANNgykXxgw42SGkMkcXOtQQevV1SGwbAbT3i7cKz6KB8ZBHC
AJiOwqtVdbQ2ilRRx822P55mmd66NTayuqr/Ff6uZlGq4wT2RatMiOHCeTxhW04J
aAfyvcvsP2MuHxFRRtFFq8QG3bZip7yWUT3O9vgrk7S/8RlrwfpFRkphIIJNR+9M
NMAIHybUvsw45RAwZ2x6egogpHZEjmOQeDqCrTREBhu+vgnXUXMozZT84B2L/kvq
dD1WWKJWT3Y/TxXhIGJ/EWwR4P7WsWHeVZ+l+k/2g19CdDgDQNI8RquOPUDLwayM
2Gd9BR3zhRuZ7ooV4a8XI8Y3pAVfkRcNVuIK0yZZtOUU+WaJasWhdB+6iTpGPscQ
T7GNRC11yFkZA1Y2IjPalrAK7RF4SYAmPPOHNicdyDbejWSXQOwfPC7vaNcRE2aS
5rnNGVTU7Arry+fC6TS3BhocMuJbzESc8qm3LXT9veQ4nBvaOds1/JZZuE2Skl8z
4JK2StoOHK7JB7ROReVIVT9tPUyntg4UV1Nui4NkmfhdLXl2+pu35Schqia85QSG
/lXH/zuMUzZ1KcOyM+jihKX3bUbRFIbtKNgX+5gJvYu42Ig604Ei0fECaog7BPf4
Nr5WQotd+91FYoAqMqFqNtvS8d0qROeYevQ8OX+p7ivplLfVGT9fSGf5pax1i/C0
7cL2G13Vt3SsZcz44XEmrmI2sVlOm2lTOdORtFd3ewTVw7SlcHqkthEGqgtGuwSF
9DQa0sqOMt6elcE+lRhZbt15/kgm9oYOsM8sysw9j735lmHfbVJmcAdys5FKKIhz
8fhnNL53o+kcPoP2G0I4AIEApru0HF2Kg1+9dkEBT7pcn/63mUCE8BmCZLmDcy3X
fa2hHXwERtWK+/12uxBNlqcr+70rq8Kcr3+ggY0f0hxQua6qSMmiFjFOK6GP4dSP
n4de/c9tHvK6bOs7orPg5FwuQoepGjXcM4NsyA/L+Gr7H2bL1GQ27uWyh1iK5ZjB
+bu0WUoojxo1jf7rEXQZIPhCqR0JLykqjpLZvRPuG/tYX156PcMGxjDqmc5Yg2gg
XCdW7PIafc83W1vUSsKIB7oPN3YyiWhd4VwU7VL4RCLWlzeXlIM7esg4K3ZmEeTZ
jjhSvKCv5VO3VQVJdpuTjydYY8IOwhjLrZnAs5iVGmjeWGH2JDyVVeOlIBEqiRb0
o6Js0Vf/aTSre0cAuILuR6uQxEJZpbjko3H5DXBDyvQhw7/cz9x47UbH3jHM5S9T
OSqFdRdqVzGlU5IEvkjmkwt7le7PrjcTjMPalQMqzEeVnT6oHMCdlMnCEgmOQeBj
Crh207AuDHeouy7yareK6RiRqhHt8KoD8IXufBkMXKKT8NPKm9wP8zC+vMMzb/3D
IWtmzzj5QjC30k8X6E2IA1fkgZNImq6c10rJI+LbdesgI5f2vHI6BLRLH1+9AQtQ
Fp0BoGijLHK+otyY6Ii3rHXdtxRCPpk1OGTsg+k4BzN8h4iSZorLCY6kt5HTKa9E
zn4VGDg96HsQdq3Z1X5vQtOykRw2Qtnkh84HvVw81oIH47KAcANDO8XclL5J1oYB
UcJv5xlQTz61u5PiVYG1qaxds9eHufLwiNapDquJuHHa9LHOmx9/shb1ZC10uUKH
PDipj80aXzObeUMuk55p2QzBUFWi1dG6dbBEMF8vqlOS3h8YkCDJc+WuhT5ppyvI
eVwpMlAdTfx41KB2I57tW0GlT2jQ61MTEN50OrWZgxvilueZ5M4U5Q/D7zHtKC4s
cwNbP/dVY7lTzRv7L2ikoXnFD3ygO66mrwR3JeM3OrUN24GOw0ngWI0XvJUC0fvw
t6DmKfCXkJRqK3lySMPYh8BD4spZsLhnN6fDqqq/GJ0APKCiRbhdsnKVonD3Wq8y
hfEjuRWQchNtXgXWEQRIut1AdcH6ahxJOmQG1O/XBDGNngR0UUmxUxXZEctDf9Zt
w1xEaJvtY0X5XIrheWozbG+4qHNGVgOWuWCOaChGghMkoLET8jRi6DxWVz03JwWx
WrE00lbfyUw76QVxbbRRTQo9UfRSLOLLeKlXAQEaKAKJQd2nCVjMlPzeKQH1tPaW
EJ0K2FeEKow1GFyq08DtPUYIFXv4CmQqdoM+J8M4zU4ZmHGL4k/iNubDKk8dFt7y
EBc9IbK+ctOQYcUgWMxx2xAMopBMNQOmrSOVjToqujE+tRjluWjg6k5s7PihwVAs
rUFwkSxmQiXMHPUL3S4RZbaKvcoi9i4qIDBoVZDEloPNcUYyu1Qf1xsBDbLpc0vz
Nc8n5xs1cypwAG+IVOvVXQi/25VJPSR95wbhk3GEP0/GwaAFUd7hCObxkdYmKlGx
z4DJtpxd+afLzQ4PpcU/W58G3GJdkuvvysKs9JtTL375Nr1IfAblKQxqrj6+Fn4F
Izk+1IQG9+66nXpQ7fODFzZ3pmiNVNnCpM6AFw2Mq7YpC+PfoFCCzDW+B82b7aWB
DZvtgAGnvIebIK4BecrvJiTi8FrVj86zAvL5jN2qa1MwEsSTnXkUN4DXfA0X9ocS
VKIjJ2Evcool4qm5cj5kh7DiucW7FrVqM+Rl7qY0fMEdxWsZj+FwNHKvM3r0TbsS
zB7uKxI1t1Zb6kr/MGkhNjxd1E1/aoivhuVAqhlLbvW++JzcpxhCSgpnct2ICSBi
2+qt1+tkTRZKjZnAMRgyv03bTU7aRUi+U//mujD6pINzGiDsahbyYezRazNO4wKp
rumVN/snTknglbI1vwicYi601XetZ6QXE1taIWJbnePw9yyqduxLj/f/ZsvbThMp
f6HsQlUyXnPvVywcOTJXvqtc8XR85KII5zpl2Fc8Zy4X1a08eidn8k1V99lVmA26
ODw7QnPcCdHQZyUV8IFRhagrLi9GCV91CDAq//7UfJCZYd95m7fZqHZW9f/Xi5ui
cqXWdckIhHSvO0upR7B3bJEMsQVnB4yegTVSiIi0mtM9bSjlXodXFb7JVWaquLht
qHJAdut+IlmkkvSNccVLlp/3zdMygMoaVAfZ7VUIxID9XYN8bcaVPYaGn7xX+dAE
CAco2R3tov1htuoxp1CCicARaY9GAfoZFVY/PVFSpf9bFPfY5NlLq4CAgQFATkAq
eo099U8OkcZ7hasQ9n5ewlHLaQOZrR7MOSiQD3juWNMPvIEz3sBKDv3hIjgBlCM7
vBgahHclgs7hxGcdFBjnfDZolij9aaeSKEoprbMQJgDZ9ztPMBV2oA+lrW8cqr/s
K0fbjk9VXkhaUg8jFLCu5HQHtFxAh+hXV3nLx8l+ELiYmtZwY6N9TOpUuq4SUtFF
T+VsG21DTVW3m14UFw02QD/iCZOQ23tf4a4xS9+dWCbhajkmKtiWXaLqKH3KEtJs
W6/8M2ph7E9KwZyklUpkfKzfOCkFKJnPfWBVAdvnSYCyQuaIRGmgT8mDh6QCLRbI
AzPk+6/YhZhcmthGgyZy3i6cGJ4bSn42qeCA03gSnvpZqnglih9A9VsEvev7b+gY
MDjf3VdVVtiA2GpM+zKGe5Z6/fYTzNLIa1iLqsOa3aawWFoDAyl0ys1fAtLRupu8
rgWP7AOOonCabRZH8XnbcLbFDuTxan82SSc9Nisao2FO53jKFrCngJmOqb7U7rnE
KYqwWl18eowt/Jcsu+4VeDZcA1Bng89Nmca1XEGTNe59/kisDojxVpb+s7noADPO
oIloJaIZUAb+7fk2AVG28igE6vKBZpnJVi3O/hD7qdWHGnR1oCYWuTh9U3IFFlMs
KbHYy0NoR9D73mu/d5l8XopZ5jM6u+qVgWtogjHseBQe7BEgzoTMcgiUBvEqO0/Y
TAquPwW/l/8qMb4ZLI6xXe5RWcwR3raavPCFp0gL3pxdoZNhocV6CEp4VDgIxEIz
VdCOlPYaimH/r3EB1xY7TsM3UD/BIbHJG837ZvHEKv2lwde2eFDocpeY7hQX57pq
MK5aN5vMQ99gdpjbuvGW8sG/P4dmIXm4XuGki04kVPNHR1daCO4rDYDz82EGHcUq
+gi0PjdvSyhypmqF/sxSLuvgtYJvBROsYMbiTiDDo4MV/apvwzTnF3Qv0/rrvBiT
T7mqdYBGbIstsJTIzqceVaPdMrh+Sa5GWZrULJpWCFeDksOCILcV9drF7n77evM+
sUSdfeh0ICQrYM8JN6QTgFcxUcBimZuCJmAalXA0UYU4GyF1mhWqa//HWDRo2exB
71CmqasS2u8NzeeBBqqfHYgmrnqATl4427IoxKEkCbAnIZLQyEufGWdL41nb7hno
H39fdzMtMrX1QOC62zHWz6oet7E7VaZhYSijEfHiWsldij04JrUpyVq3o8EhH9eA
XSFojA/uyZhk/48lLPdPzDPv9Cbum1jalq4kIy0DZnEzViOOHxYyNv9ttEHhHwPh
DZiEuFxqh7Oy2Ptgsv+t4btB+lthIg05x4ULkpMAYotn5DySwJuDRBnOsQzZtIgN
hLMjE4hawqepxTAztaqYq4I8faZd3+X13KLls/J8kmGZT8NKeIR/ZKoFt8KBZUPD
7Uh20QSV6MfHA2YNHPPV/sSt5lXani/usU+/dY9NDlfkYLPMLIlqH2Xe3Vr9HnRn
1lovpZdffepH0ge0BumORw7VnGtcE2OKia+TRRlrENTkwFp0mPBAwhZE9dR+U2pU
osEqSsHiZ9lIjQkG7AM732nCRGmYekKG+Ipn2dZ6AY9MtGTWtHdUQ6R6ze6X+5Wl
xD5xOsA+xLibz5vg08iXfyyl4GPlwqwCekKgKWgysjTq8KiL4ac03B+SCdERP7il
3rJJ47v5RH6XLxWJw0sxedqh3rtejB2fKjXDBdGhPHvMX5kocMh/P3Nq7Am4AkvY
xYbizrVCJ8QvObqLxxQ3koOw9rqyeJowo04qFOMn4j+89TNZYqa/MV3LJw9UCkjJ
ubRLs0UMnaya8m4ra/9OnnEev+uCSlxTpeGIAPAPO9iLZYRvtwS1qijeU4upkge6
4b8Xw0VdbHaH1BJdeYMpLwygS6iAfAWCiBBaCpwcJ7NAebv/aup6vykVhcVbm/Yw
Ma1J7v8YJeozh22GcCZPnZzTiGRgGHyorhtCIBJ1Utso3TKeK6hBzZN3jPKNVHWo
YhHkVTbkWVKrwHyKL0jKmGcaR6tllvnQy1CJrK+cvO1SlIwUpPTolo2cI8x/6w1C
lrQTzYGkkHrik0ND/X5tUb+vYQyt8YHCRvnlrqhaakzBXebcRRnUAs2p50XPcyso
3p4S5fRJ2V+vaXJtdYaaWbt/KZvHs5NNvzVwNHl8ba0D0K62dsTLxXX8El/cnp+Z
A/iJWagU+wZCORTCVCaYOxJE+SVjNN654pkh3RMULK2HAA9ptb+5c9r90vbjgi25
Nnl/DQB/bqG3OBILSt/By10Tc0G027x2yNKhKjhXbavjXFSk8sQWGE4ZzHvvnPMX
MLzxPlK8uIndG854iyZtFeyStdk59pLBzHDgCMTuSp7eBX2MiKErwvdPFib1FlQV
8ZZqHWd3UNPuN1Axv7BKYy8wG9MzgrqroxgmJNsOqVAuephodLIyFEyHXqj0f950
1I2SUoJTTHwmMTYIMyyahb7cmKfXb9Iq+SX5gAL/iEuTcSG6JfjGkCYJL0tJJ5l/
C+BVAMRNvP2RUeI2YGrFBP2Nd1zN5MOGHR9M/8hhvwyFNxBFOxXiBuolRtjJVrCn
V9qMxLsdKR9t4VCcwR0n2OzMMWesbAy0vA/U2FR8J3ijr0CRV+0vAC0X7AZ2o5zM
ZPiABIaJ6JlDcmfoyc0EB8i3n9M2OcPRJj6jfnZxBohCMGV1CU9Gf9L1m+B/SHVI
vsHpgUD3AcEKT+JGWhMnjDwyS9efBEnRsVBm3yZ/YkJk9gQN0c9PDKaNpnSM5cXh
f6yuQhhwcypaVx4SvOUJVQ/y7iZ8O72tIwhbg8c5QtQN4RLvxja3I2oi5g00zHs4
kp4UQISlk3BBJRoCYbVdnkY5EjHNNoBBU+Y2WJsLyoQuD8uM1UB7WTqk1ggZnFt5
rG5q9lrxOo1LSK2wxD7vKPBMlcNVT0Vz3poRltk2/+fHNuEa5hv9dWQ0/oRzURBY
u7Dsa192Lpt3wkCGU3oJZJMP1Xy81FkW7SdqSAlTs6Z0TioFDvayRZ/q60HT9zXd
LUotx1aNOfCaEp/pCiXsNiCv7+/6O3WEH3N9TBloRQ0IEwDT0pYMQ7SivScG5HP/
A3leydc99j0e4wMojcWDGf5ZgYfUQ9SB0pQGIWirp3upE3Qzlfwxw69acgdp1h+O
brsGd2WLaCnTXv+GykQNg+Hqf0CDOi+27ZtgsjewjxGUdnvK6nDIINn+c7Ps5Bwi
lWyjTtT/i9/DJ8LhmcuqPzDdEmxxAbj4OXGy2S1JssXPDNPRDQSDj/xhW8T6C2No
58K6RO0/X0yhP5kHtKZ/iK1XLm8Ny69w2j05AbNfev1gBq3+Q785/WKaPwX36kAS
DZjs6j3jgH6O9UE7MxH1mbA5xRtsiPyS/1sauzb9H0i0Eb14rtLaVq1zrY2OtoZE
kbLySEpv+tJjHR43MmvN526a9/p7bPX1Sdubr+PBPb7+uGuyiLkBZKZ+RZvWpBcq
o91vslg2hqSXdNbqVfGYzTZLfjOQFfkqbB7YCQJ2NgEFM917rbaaF7oio5kvXBfc
97YzdBoVbPP3k1CCjxTKxN3LQ7hevNEUzNYz3UoqixsZRCcE5dxvz2vHMdlDCMO4
l43SGvJC8cPOWDMRAXZ4zB9/GdDTWtLUBfzNTm2Y2aYRT3nB8Lgk6kKL1qHdNVlM
O+jf/UIGcXysD7wj1NWoDbyrLIy9QnLCMocCjsYtGAk7gJUdm1RFOSvHWrPcbIIa
wIdUVhN0Rg5XQ+gsSHtkebBhHwvhykbz+4fy8aGFThu4iRVmRotIOfhxKCROP879
Mg0nN5A8Vu+7Zwe1z09WI3cBCS4ra1QHwqoHDT5E/oztoo+mN7mRlCVXiKlQpI4j
KlesJF7YOZXdqj04ewfDXGX8wmZgu/NRNpKYIx5Yb47nb/pW5ev3hiXpBVzY7AEL
8S1xNla4hPPezQJQySZlOVRVJVGHt2+BigQcYddw/5Z9l24LEAMxbaXbtvLUqKZr
syvwOPi1YuvmYJzQmts0kbEw3p3MBsyOH/ORQ6FyxRKzTyXBgbkaAPQCbGhsdbtw
btBc77jz1OTxMpXJB2i9KkQlBsVSD+wkR4iX/nlfKxMmasELGbjmBLdyszxJGAIP
xIDLHnZnLUW5tTtJkBcvSgfenUGJGrTdh4XkEDADUDToD8ATfkd6WhbbwnJ6p53t
Ie6LbCOaT5i5N3iqzngeQA6Nd8gfMze1/h7LbWeUeHR31H/Ufox8ymqch8l9cbky
T1F0E8abgK/KzquREMGztRKDEq42m9MBPk1O2t65HNuA4OldAMd40+rkk1fqAbEy
52p6+9PMKNQsxfsXVxmbjukaTsisC1hFcf+HOGsDZoyYfE5nq3DjLjzsYQdU8e3F
jSe4TXV3fccQR0qAi+aC+80xewECIbPcn+JK0POMhEcoJHRi3BwbBJm8l2bjGQMA
WjngmCIbGg+HAlSAzdf8Eauw5JFa3bM5b23mgwxWISfCqAp8Vuv3NFpimk301klC
w6GCpM3d52y5FstA2CRINrLftj3r7v2W+tkQx/+KPBdUZoMDlBKlo2wLmmH7tLYK
/7VtXZU7SLi1ajTkqZwxTe0ksQe63s3JlUUJ2BitgeEZ5lPQHKH6P/O345gwToZ1
1oc/IM+xBlt7Z1iEHJvBmRW0ONeqYtQUd1SQjErUuSsxQJB8TKYWjs4YeR/8G6dH
MjljQuxP8cXMcV8bGDi9lI3b8I/6AhvH2dmDMOPfo3HOprYiATdHqdXFeuHYBZB7
0dUwQHkVIjl37VpAtp8ZQZYVWs8FdjEqwhh+iER6OUP8sV6XMg3C0c2Z3XOT8Ykf
xIjCxuzjpbFgdLw3y7hGyVdEziGi8DZFwxjWJz/KxW7UohSbshINO0mJNX8/0Fn+
GGqs1cmAaxrtMqXeC7MYjc7mk5FoYDUF0BuKFgspHyQvibiWAlHcaiLCuW6wdyV7
bG4cvz4xp3BaC3v/cVrLQRha9uI+r2/MfN5CvkfQq7vpp9616Min8U65hmUHq8Ee
UcU+EVc/sBQgqCxKepb/n0MDPBbLu2qcue/OP1nANe8ecFOiQczmNrmDe/0CFfvg
3r2i4nKekiEHEjhF7aK/RL91YYJUrQaZLhPuMFsk0QO+MrZyyAJChykYnuNY33+U
/JloPjdImzf3KtqRMCDGaT+itsxvzk9XmnYV/5etYVnTZM+ImzO0i3oDjP/QvE20
F7RgJAVLxQDoUCSa8m7Y9pbm5WSYMX3zN4H4SkNn6anc2US6R8II1ISwjTVILeAb
H21bQi52bNNAWwWSdBVFA0/fXDjPJlvFhoYkzggUOXyeIrgH9UQaMZ+1OBwTLYx8
XG41Jz0cQGqT6MpLPq+VVb8XZsiTQlrZJ/zDoXVTGqrdxs85n5OxmFYD4qtGPALJ
9Kgsx0APtWr+y+/IiL/5KpdjvwE+309Zfo9iHh9D+3DG0j0tJVmUxyE+zPxbs+Rx
kjCqIXju8UTVVSl0YxowwB0uUkUIHQwdtOnz0bggtPcYnjCGsWJ7RU+DTr15Cag7
ZpDSwylMUYz/WdIC+MX3rNfUPFb1/tHpSH+zdTjZGYJOfKoJsolgK3Lk/S/SnxlB
bEBvwxWg5DKJGqIlvanHBMOZY3QUQHtsZreFCPXKuyJpJU4ojsRtbhMahy5OpvuA
AiNUARWatTITDkpokqR/P97Qf/Fkf4ccoLVWdbPoCdIwBirne+jA/AVXkUcDsL7r
WYs+w8rZCRQOoJO+S7t6kA/LNXc0ZeGMOFY3/N94bm8vryyBNVo/fMKoaQR9IvLc
KX4/nC9EOsJrA7LSWspHQ1JUOJNJAiPgzVb8X29NwvHsKcQJYJEareNZwahs73Qe
T/d5+G0Rmznx4bA2gtsaMyNdLgRJNBrUnSfzml1KjxAUnjw4jysDCRHULBxWLcOZ
3vuPA4Aqj8yOHlN90Sj3//y7cHln48TejVNojgUryM+trvzfsKCsJyVYCyy5Rqso
rosqLx2oKX2WBTVdfAKssgmC/Qk9tSESm0rXK4dPkQQIVpwxUZoRkGoO7zj/oFGU
zw+Sg3oXoPz5etnxwea0KObyeeh250uc122OA8AgLamj0FasgqUYitlucdT4wVkZ
6IrxVrSC6GU3xVWU70x/6jSZNrGRIW/oQWoRKgEgBwgs5TWg6eYhh28WLQ8la6qf
LtYLJCXt6aC5fUVf8iDMAx8rLBpk332YorOyiHxUReZjg0vUJai5q6X9B8SoGiXG
yV49QCptJbU34BIhV3R5ZWQu075IqS/6SZ9QNLm0SHUbWZakXE55dpob+7cxRYy9
ZZ8nSNdYdQTUtfzV/+S8PqbuaI4K2TfjQL0CzP9l8dwxRZQzvVRxw8YiaV9kk3h6
tI8pZmM+0X1QPBs9T7+x0vzjlO90S9ieoPeC7Qlyn6KZ4KI/bJly386pJycpg8SA
8+smtujvIm2CxwPM49Tn01IL6Dwq7ttFjIzgDWgxXE5ZvmBYc6MtqxkOlyRmKr8T
bZudHS1lJBfCKoIB7BP+vVb/G80RVATPc04LC+tQuHNiZygdHJSlzGiAmlLhwoFn
lN+NRYWbqnIR0/2itnw7fBpxZBnIY8KoTicEvAHq0Bp3LHXMbsXOc+t1PJ1MkX4W
FK5tfWvnQCXdhI1t8F48GgVGUQUNUDylTqVy6g7xgFpwXeUuZEdWQUbYNpqx3RFO
M3wF/g30vaHjZctlsT3sKtxt1kk+ZGYTbAfVY8sFQq9fAu+QkIKjjkEgmPi0Faxv
Wy7gJt5AYpy10HUxzp4tPag8E/7JL8ojc0qHyCdRGpUs2DlzefTzyKd1BiAm9Ngy
yBKpmGXJcURYfVizzdU7Xju9tYljWr6DLmjO4tUvnB4mO1CvZfZfzJBwj4j8OziL
WL03ER6GWg2a5HeL9k/3A4PDzDm94X6tUfdncgeH/r+hHsb6Zga5/xQRN8kZlUVz
kesw037piIOH1E5imLKE4MUfAe4Pn4KgBMHO/KLTbxEGtMdL0ELHcEYR5tUXPnFo
JgAqtPbAXG7YVzuT6DtUJnHRcpkXows3QzBQU3AeM1UdMvPancBawaIgyWubW0n0
jjSgShVfuJWGtsX+c7JZcU6zW1NDRcIuf+MUJdXMqsmwUDFC3w4SNSTgtKF/n0uN
fg/Ozm+rsd2SkSjeCcmThyXud5WLGZUjfXod2Ijc6rTR/zdeH/hOAaZWX+9rFtLA
TcFqrkpJ3t/AU/7Uu0ANZZhD5DARKNPpAtszsbvIfGxJeMlauDVamDCJYWf0ZPJI
G2tNViZC59Vd/+Rcw5RLCdByqXm/dQ/0DqoAIRJaWWHrJ4QqFfBbEvrgt7TtP7Uk
8ws/Tk5e3iWkb613dWP2yjcI2myqFnHUvIrfL+QNYNBHfwk40xIQ8lzInEr4eZ+B
U4Y9dbh6eY8wSnxuKFg1RtigZlNjmCeBy9bc4qk6uRz7IXdMBbWrJFuUG2Hy2Pik
5OFMH2Z7fwKoQFXsK1NZOgrOchAQEQdwgJIq3h3JFOsy7/r7jriSGbYVoALOJ9J0
WwEL0GVN6ERgiIrLcDsdqMJBRgW2nhmQQF6Dxi6J1YKsXkWZyaRdKcIG27l+4UIw
pyCejZMR7ZlJ8EbkEpcjO5dMiH1c8dY3jCS60auDqIDlJXbMtTD4cXJcNTgNrSuV
hYLfOMZN53QQfeNBeglr3jre2T8P//Jq6/bp321PIXzhczJ8LEAJU1rKKazNWk2X
II3qo59ltWdJRVB109MVy0R9ZX97N9dqyk530m+1tzZAkjjT6M4s/dHRxdCsPa6a
ctXBIEpyL8EDJHGRBSd0uIX5ujqtJmHeV1lwvvad96wJbq7s0H7ZX+rnaUM04Hvo
9vxWeLlUaPQxfhwvEl8RL+MVH8bskpLlc4XxPu3jtcblLiIWxx0/SpdX9fo7qh3Y
3KT4DU9agtDJKSRzoMtFaMhzAEa72R+ADugkWT1bZHfwRW++4sg0HorXVlj+dSjQ
QB23IEAc7IppUwaKWW7Jm9kwzikvm2H3XjXXB8WVq4wNHg92NBcWV61JtDeMJD7l
yx9T0PwT+wATlbNl94r1W3kk/7bG4luDZ9DoibmlDSbMyQrTKeNu9le34Bw/OKGc
CSpwbzsZqhKZZ7BscJ3gbPDFnrjZOtA2o/2GwmKGlbCwDKLPhmu+HUSR3RkLTGz7
hpMCG8tskG0cTX5p61bup0a4VR6VaZn9GySfM+eldkS7rEyG4XEWYWlFVLvHa2Bc
dw4Tb/KYWg4EUP90PQx/nGkt94dr0mByH9nWNHP/irTDYNG1X6hkh6BlfgVauSTp
CxsqP3PQRiq1od5HNEMib6OwxxHLKUhx7tUgXuq4/5+HYDfGC/OX8CnfyDSoGZJm
ois62FLg1iOMsv5WlRvoWYCyT9rXP82q26gr/N25/ayKbzHcO2vmFPdqjze/F9NR
3MpmSEqih4vLY8jzku1frWz3h5NadihjuoRqYuWZNpMYNIi34lajsylxebLUM6WY
wU7X/5pGKU8mYM26y/jZf1O85BnDfLd8nG++BG7x02fiG5POzY4yQJgpGfXBVIgx
zHvWxLUY7Em8V5qcRIft2YDOfgBq4XtgdgDTvF64pZDTdSK9hhdzjHFowCXK36nN
TaWeCSx3wIIWK8mR8m21nbnPTD9fq0+osTbcBmL2vQ6qcEvgd2UF0bQaPVJC2aAQ
ZtrE1EumWhvkvzRK1GDCd7CJ8HRXUUCUZKKH4fxEUjbJFaw0klFiB+E0oDKDEdtd
elgpIeDmTA9t8TZnj3j03+tRj6LGDLrruUJHJDEul3bnPoKDFQxe7pwmnQkZiHw6
20k+6mTfADMeUEVUiK97oVF/QMjSv4gCrxYsY8YlbuHwk41rxsJ2Dp3UZuwvB+dI
kH38Zggx1jhsmGLJ3ErF7OSgRlyHBZBa58Gep5AT5aEo0BxIS5YyFQNNdBWgVI/B
tW6GQS9lzy4ZwHLNwota3IRHqfP9HrQQ/sAE+xMJde7JsMC+AlddopTmM/C5FW9g
0Eys0TyGV3XlGgqdNypw/PO9K+oUiG3E1Mpls0tJm+kVsGxj/I56JLpGMw+wQy8X
onNQUPoQsAZYWipmv+GzHwQycOAn76TaxSfTp1yKhkX7Zx9KMdy9HuQIhRe7F5l8
ngVWLoi1Wf2wY+sXeXENA6Vcn2eNXUDth2AN9gBouY3HE9ayO17P/D3LnNbR5RXs
407iWmOTdp8I28ke1kTwp0Pf3qgiSlL3IErLc7Tj/5SrvWUtJavmB8ByatXV76JX
Livkrhu8Sk1xuOfSykB5264wwHPaAdF+rGez1zVq5M50p6EEEo2/yuh+KZHDzj/D
dqIR54POEqkZc8oVvYMcUXjgzzFiVftaogwH28TnlVk5pMMVVwksXFpPi0HhmkoM
FK0FjkwOoq/NliM8eZvtT29/BDIC3ZMG2/4h4VdS8afvCEK5wcCB8m8ENvMId0d7
Bl9sZdBXMEmMKsmQ6nVLRUTcbnmQanRVNMmyk16RmHuhB73AyfhlVp6nsbEDPOvN
IDNgE7aScu9P2XkEqFXWQG1r0OssmilQaH0hNbOv/2RWi+qMGa7qu93SvcxTXxU4
IF7RlEi0kbIanT6S2uujvNbC2jPr9dxBjvDgc1S7sHaa26Vm0TZWrkNF3pZ0L3c1
1TahV5PZLliahk9kx82sr+/Hosb8MpZOeq9WofCIwBum63Cqe5T6xCD6r9ZvW8+G
kSYOLuMpcIn2e7Iaj7miUtQMgMqlbtzp7sCE4SHi0kRclq0BULTsrzPMPF9Bav/4
UiMiTB9NQsKaW6DBJe68dxMFDVn3a6kOpDAOG/TncMrUjoC9ErLi+2o38qMblfjT
mmKZJCc95G3DviNzOhhRqBwyvG3Gu0di+k65OpI7RIw4htcONMnuECcbTV/RBE+Q
5zMOEp8CA6SGgAnkOgnsRttb47XV9wF8fFZtszPeiJYDKsM0QyDlR2ODo6ABZdFk
5RWmDT1HIFnyCYrOE49IaHoEUTlCw7sHbA6bsmOB0I5jSSOzX4K/xtwYBW+YrJxs
990A221PZpsfSaDdtdIboXXwr05fkS/0nIPqmppD6lVng2TkFOHS0Mxf8gZB/DUg
cegxkvsyzDrNcUAEYIvOuvbNpDp9RtCy6qwDXzTFwEi9NfI6Aie/AM2NI7GTVveI
snEFpigQDXWCLx3UgSDHh05VwVNh1W9AlK8ZvITSTaoSAltkuk7HF+Xzxl+R4jPo
9tO/jKk+w2vZyEvhlC6qhjebnGNiu12JjjjqKmXTttgFBrLE/Ju1ylrKSGCWlNmc
J0fiB/HOXp+4kF1AbDW7eh7GkY8IfoQ4MpWsP3FWEi0WRQgBSMfWX91HDzple7ac
c4dFu6ApI8VRxZv9BJIh3SfNCWWEzlfqbY3GZkkGOYUw2WgzWqbrTVLD5MM9vFAu
iVsEknCcA/kIXMwRbKosV8h5EVMxoyk64dSUtNxmkDQjwBNp8p301gJ0faOFhZxM
GxINejMuAJih73+itXPJANKUxpgVX4tnoOdCwNmfmgljfHpdjtCuWlo7+0X0AB2I
Q3XUmBAKZVH7gFKU9l+MVKH19B6vVRcHFFzRTViaOaXMnlrtNQnBTGXJUu84GhHm
vYejs1RN6dOnG1ZAJhESezHYk2rPBNC55nDD+IbciO2Zci/2jAHQIi/y5gww29/l
ZekJHHfcQ9Em89yurPuXAkvtcO0CpGgimtasuEfOgtrRX/oTNbtYwvGoX8ACpnE+
NwsiJvJFdlxhnLYwvwkibAlXAVpE0W2g82j/o0CCQARiKE+AU3lA4hi21Z7qmhUa
/pdjTc/2UPDbGp3MOFiCZ09LvGiTo7fXHdTeCwj1y0Mh6rv6+83/tmJ8RT9eCCud
dZxEn9aUzBVuqT/tqaoE0yi+cWzQMOQVqUqVgHKbMcFz2MA9/AbLVjyzhwYxvDCA
UUc8UNcmQTgQoHAhen2Ggx2nOIzqn7lpNaSRUoG13UlfpmO32YfDdyZw6BGOMP9U
1CCtAjvO1X6dDS0RMbn0KAFdonWBCazlkq199oXMRjX0o3EOCbdlDh8LPgEp/oxx
uKIKFi+d+KZu3dtJHfLSvSrNPkGP9pTTtBEM1p4zHd6xo1PQ0HBXAGhKliTF7Wxo
xaxlnb4Li6eWi9mqMmU/zFudnRWyUL61ZFyYbghH1xkGMgMD2cD5YQFbaTrggfap
EwwIrl4p5Hlf2yjH2cyBpbHW/LrZ0k3L92+g5iSPbXM7iTDsjv4TwMHBxhoxdGxQ
SfR/nKrhZtbzYe7T7clug8GnIMSj1tDoOs2PsjDafy0iZbsSi/Vt3hDXfwV6DebN
PW5zw6XBqRg7mPzciL/nSjBotPTWCt9+6Yw7N4a0dGHZ/7XFFFlA3lpIEJb3+tuA
C2HuAGHrwL3pogNg5+4qlyIjH1MNV+yFe6lPzUR4QJaEbxnRYhbioOEfqbCkN5oZ
XXkAl3TQeC4URfApLqckl8Ki47snx8vIkxV2igsf7BBrqTe4rVgt535boSYRx3kj
9QUlsF/vzOkAztW25uaFL5Hci35VLVmE+BMNb0RfUwzdQoHAI0G/L+CYrGc+2lMX
VCLB1s8I7nEpXK4xmjszfSvYlZlviynfEEidfPdPcVltL54dG9msbe6u3SuwvBqH
2/y22QmKOuqzNwKS5vDEEQiGqvkMZ6gvW50/jVNv2gFJWbyFvcAfx7dZG96ILMjV
UNM7cDQWyCQsckEzn5Ad2et9+fV2/fDS4D7EriUfNjZ9Gp9EUJQnGMlpBDaXzkEl
2InZwng/41Um1z/x8b97Ts6ZFZ4SvwMQDPYjn4Ft1aHlx4LZSNhhbC9ki+Hl0p40
+YUuV31lKuFUkWCnH4KLhQRkNGVTO/z5bbVehNdgzHXInvbKm3iLiNudyn9O8XrF
ZcBqjsDN9FandFNv1eesfWUkzu4UA6I+38rFKSoMli/7rv2o4QzLMPJET3SG4lUZ
ralT/L0Lu47TdYEafK8wn1Q63TtV+gm/ARmvT08GOnf9kikuwDfy9MgbOyp1aEYJ
L62RPflbE5i/kXgCtyBbrWQbD4ok7z3L5bR4/4w4cSQ+wpzKgFqP5R2Xk6zYDJBs
gAx+mSaTD0QkzWNnIHYU5++GZwQuY8OiHdEpM2qzzBwhYvhvC4qef4UEX9u5FgmG
MWaULOn7sQLRp61JamSGFEAwB24T832GtsMKqyc9RJMUPLormI2B+biwSnkOai7O
DGYDoax4eFORu4c18qrWh8V5PvtkGUQLCgVB2EYx/vRuBv6imIFW/2yEMni9ECu6
2OhgrHvX1bzzAEdfcAIE9eJl+IjwBXr4F4MZ6x92qarnDj9KhCvQ8DVW8OrSDIOl
BBCtfJfeE9eDiCxvxgW7/ymvCxf9OzY2ZVOIm4yQDWEGpeKFvefCfQNZUWU7fGeW
/75iuBCcm+5+zdmix3ulVI6Im/ZpgfE8Q9zzNz6QIMPEdGp7pchthA0RJcDqoD83
7i7D+fuHrQpK5+dB4nPzbPND7ONvgZ8xK5rnxK/695pfgY+hfDEfQ4SM4wB/boOa
ahHz37oyS//rMW3WjC9Se0qL66fCSIz4+t+FRJtBMyLi0wLo0ajlTYVNMGuJdJKk
EF5SBOFPzKYZXsBVcT2TKI3xzodPceiMBcm3AJwRXQo1vl8YuKdlrs6ztWC/A8e7
vXUSEmZCqLfXqmOIUSsApEFPV1dtLEEnZFCz2hbskROIu1fF0F4+t+zkrdh9bAtk
qffl0lRGjBjly0+VZuvbh7/nu/sGh0RWkk4Fv/5GHS7AfEC28DaCJkYUSeDTmG5N
Fe36kltznLHKkNWBhL9kJkturYswX5bOPNQY2j9KlbXV6d5y5ZngrOgPSPNxoWS7
SbC8zktJhG2S9Jv87Vd3HnGqo5++mjZSJ0flBwVBDKPpHh2Z+kafCvgzBfdDfc4W
eNwJjiVZ9p9iyT2plgTz+EOgRmI36K6WDrX2th1hyQMhlcV5ZaStUw2gl+f+vt5d
FzmITgsmorL0AGOWQwrH22DlDJe83bcl7lVD+M9sKKPQJYeSITe2mqMWb69DM4XR
KWgZvvT8nSBPpPlEyAorVS5v/bkHpYp18LvvGdP9FfALGxLfUU3jgPBWlJOjPxH0
BqkSjTRFTrcu16V2wEOnDgCINPx43pjEL/k12cKJ3Vwfn2QiSaJ4BlOCN26owe87
caLfh+91P5o6Hl4VrRFUgbO+Wpr985r4B98fwAEnAibmu23KkixXEJ8jv/1A8xNP
D7Ji37nWbFUzgmOLsAetDX5YUJoOTjLHOPYMUvi95yt5dRd6lLejQAHQvvoUy2Vv
xN2tElvStavONneZNq64UsW7h6dOUTVbqeMEfh+xIxDBQyu2dpZk7jxEiUbrMrXN
R1KdCrQnBFnj3ZT489bqowT/HjB6pDlkP+Ix40QZeK9Fvr2ozEnuCajwGcr/hYzz
AonmSaAIa4T3s5y7AIePUR4zkRCibt8cfn9vYfZBI+Y6vDj+b9P08kHbRfuHLRIs
7NiJU3CDV9yKFD8XmXCRIfJS8Og0qSdV3AjtIq3PkhTvukX5IC1qnd93M0ATmVhs
5n7vi/Ph02uDwAj8CL/hKVxXwn1T3lzk4sWWUM5xz4yD1xc2qSCt2iM2aIwk0l6C
dqu39L/anAYNpklp+yS0B5mpqTzA5PpvzoGkAf/LBmFnM5Pek+QcptaQ15QV/RL6
d7Nr5vq+Yu+ol2wXAtHaVD8pKDYnYr8p4fbjFZxR1AVjBKL0ouxBxVqaXb6GcFQV
h1kug7zZ+F0jqYFcK0hnF4F9TvNNY07pYYw63hyyrieVxcTuwHbfBfcyLGCVL1ru
NF9PpymOm0Fe7vHzU9WCkILFHBDdgqFzJQNRnkKdsQ6D7KFA5PqqWP+ezecz8fNw
F0Y5OeDM0C7oK54I18beAMLClF1pUX3YY55CDqSR/OheqzuuzucK5ZNkXP+Tnooy
IZ7aXzO4BnIbLd0Fm4TzJEWAry2lE0XAwLHLtgfTPQ1jt/kwsM2Uez9yArl4HCcg
EbkDJlWdtQ7GglCimhKke08bm83lMsduwlOsJG1S51mQ0k9Oyiymv0m6+X644CLH
SqbhN4a7HC8YvCNgzpVm0JC/pJL27Ensv+zX5fxv92SqfuZr2cHm9DV8gPiaBUTY
X4QKpBxYbNbf3A7nfCtvRiI+OL2EXXQjGtf9FNh7PMpv5YExPK7gzpenNitDh1T0
hyq+BXZK53vXd7SDn/uqAROJZKpRL5jjDrGJpCZroeQPHlKLEsdxCT3M0snHrHNG
drPTXAZSTdt03UJqfMR9dxoGljypdh+UAhsXG/NJLf81wBFfRaLX4ee2rlWOijhr
80fFRVYFuLnQahBLUleI+jfgLPVUuCQj4cs6iKP0CPcdsOQXvVkIWI511Fjf3tWC
qOVWGgxmHyS7f+eFuSkiFM5tRwpfepjc4dbl1fOhZ37/RSQFFwpf1/DUrvObbaji
MRGuBqvcjtSm9ukX557sHX3GhCbMIsVScQsA4r+OSJYD6G+8GRWNFZeozLKON2D+
xABK5nZ6AeHG8nT6hGEPMBDTUnTFyt4D75KQplVOXMM2Xu3Ns9/REG0uQh6ePFMN
qqNNB/XbYBrOpudZenX6QLhgp8CyayH0ghN+T8bUGjQmExKG5AXxQs18/1hKftfz
rMcBvyIxWQkIFUExeTUkG1PPUgUQiK5xHNs9aIICr4OCY0fI6NFk4Xlf0bcSa+U1
YcItG0xpH96uAwkyLi6MQTmaiW8mX4aKZzZqgiOt2dg5uTryWQ1Yyz+ygA0fJ+m+
e/vj6p48FhoJPyRaKXZmJj6/BrYN1QoLTxHKYH/Kv0FaLNh/NiGiHUtw1GJecMUH
n3CZjqKLD0/Whu6qTvhmSro7tGMkOGp4ealQ38w6E/lapK69z7jGBtPsaTf8wR8J
PD28wqDEQ4gB7x48pN7yWUGxKzF+izAm3fSNEIy0iTs6HQZ2yXF0y4aaIajbV141
x7ruL3oLSOVs2d02apRrIz6t7JGzQ2Q+N+xjxpHh1zKWhy/J53DOd/VJa4ZD2JHi
/s281gO4jy2vk6IVYXzqp7QiwghINHkchy5j3c4HQfJmfVTisGp5mowWaekVKh/k
5zkTefOn+cHwtm32KhzeB+EGTTkLfVVn/XEMiwe2di5OgYM72E2+kMCQjO9B30b7
EuMfaXseOg4O6rKjTj+QAsSzcOhtt17NEDfLzGq/xZ6YCzXskEF8CO34i/XGsQKr
wJYMUmiFFzwokhqBioG/BeVi38gkaaTHvwCVnVU0qaUDgvg17EMbA6cWi3emQ+wm
Zvls6mr4ZUSBqVAcpHZNMMBcviKsIsp1sJSe6RVYNcufjKiGo5YyNLQUEG5gQQ8l
YC46brbRMGbqhx+3wPlkwHIZBTWIgq4Dz5JKsYvtL3etrdOcbAzE/slicuv25N95
2l/WUZnPhrTMjCBXfsRlKBcJEEExKMphrCaDS/A41w8b7ChJzSJHmAOAmxTpBthi
yNoXKF67hZzjW7F22+kYnOo28vVLeh/uzZ7xhqfF9LZObNhzoBVbYNNR9rZ/rxSP
MmDCMIMWOzFJa7oRd9nF6ci+n5AAsc7AgMsb9S3HNgwwS3X0CHjLFw0wIykNxRwQ
hkR4XHnHoeW3nBHA6KjlDHTtMDvoJaKvc/3zKLHsOKfi4T+Bc2KSYORl/JYxnbBV
Abv5bzKCBaYIi+V70u8T3Y3NrkOaxQNt1VrOzuTXJK8my9WBgOPmuPxAv5fDcMJD
uBrt4SgBWXv4dLP5SdebOm3RWn9uQqI0wkD1bXe7QD0tVlR5/IDBwq/k/Jnezqbl
xob1zKYRb1OwGIAkF6HTelfObNJ6kUE/FbWp0qB5RcTq6dDPke94lR7/Vh4KdFL2
qyqGjSBx+x1jZfzagKrGbatGrR2I05KZMu42zn3YpOWlfTN3TWvMkrgC/82lwaqC
6N0r9JrUl4jl/ibPq4GCBS8RIhn2wjXHyQd6ZuYVUoUvbt78C6CKw38y3u7c54a8
/Q/h+GKmoOyVJoCwjftE6jUi9gbdokXAy5YxvHuP94zL1U4XFab1h0w7iCBzMWVm
8vssrOnkXkROtatSPWVE8CLFcqYoPBtaCYRAoidJu67xdwt+SUjUmGWSO3gZ92//
AWVaLSfoiB3YYYyD41QuL/WGobwI5P7NLfoDEPAmw/jtMPhDM7wAE5/knrX3YHpv
8Yf0oxXezWgkhcHxvWDXvCg6x0UH2g+1Meka72wE+jTcJqEhox3ITJ8umWDK/IPL
f5G0S05iroYPqZLDWX8KFDS56NDFYNqAz5exP4+W5qQ9cfUynxXdJxkLBWUMa1Iz
1paYGK5iJOobZszF7jCxgzSoI4POaEfwzvvRfov075OZHlp/cJMonbx9s/adMpRA
FYT6bPnrRuxkcXxASDTztiTb5MQYuLbj3nApW803mUQtxfsoAoXss6vdFUadS12g
j6YguSnF4t9Sv36VxQvra0BrSEQ5kx7sEHZGaYVYb0+5PSOesvq+6CL1LnRVJX2v
jG4amdmhJFUYf7dnNsPz5bfDEaT3+gWMH5EazXTI2lygd5ms8HVJIWnj+gWJSuOT
kN66VJXioj0wkL4DKOu76N1obpE8l1Es71usZCLPZeO7ot8KiLP3bFq1XsrF7uNH
ih1iBbwWkWiQBBIfYG8U8LJAr4onLKlQxO8TZ7fRNcEdwWHgmvPSb8J6lUGOz4r3
8BK6c6p7p3vSeH9MhiGNcyKi8c3ORVeyuFZvt10K5V+p1glZPr9ovI1mcRPwFSjA
KShBSRw0b903d7maKUU7YOtW222bse2jUOpI2zzpJYSjLjayuucjsi31Gtjpjqfc
cto5iAvhOh+iMIDsyHpuPt7j1z3uqGuhcq47pLN+PnEi+HLTjfnah4qzozX376zJ
yY2DwxRg4BansWpfk2q2yAT5wH8fISzoCRi6bnQhQIZQLxDfhY7SBwfd9JneA5vW
//v8fGVo6vgDACC6y47ba+ywymeYgAX9fTNT8s4o2me6s//+N5+1QmpS7n2e2dRj
RdEulVUr+R+2iyQAu5XoeSPD0ERFLkC2jExY9pTyXAsX4pr55LBKscOyOLMdG3yY
MXBSUl054/8Da1Qg108IBTtJO++gpyy6kayQtnwmZs9bT48wFfUFNbkklKuwBUCB
bEnPNj0Td51qQTXG0MIE/Af0c5UTK/XEi6gpQXvDGo58cF9wj6kBihOABlz6cBRH
MQr/rysgs4XcqVUg0Lb5j1NYVV85dSKjByBLc0RF4kL0nfGvkyNSrveMl6uTfAM6
Mb/krj4n1zz8Bmq2SHjAqWOktm7M5J/wvdHM6o7Yio7RkU7vcccEK6Oe668OFyFX
+hPJHQblMJRWHpjg2xRSE7n4TTYJ52ayqZwDLN37Bn8iqwNBzMelrE1iR0LzfOol
c9d7Gow8CBfAZegUBiQlRdImWNwhfPidNQrzAVb4JoHP5/rOqy4606y6KlwtkAfj
MO2px/2zgfSo7AMk0BwsxAtSiw1F9xIJ6N3en27ADbiHSsJmFWVaCyjy2M6xWJjs
HvbXYRTU670+YV4rzBwRImZCtGYdDk+p29Ar6UOhM0cPHvui4D9br7TYsTDGccgz
dxFscNRcdXi+ZlvWrddgrE8clAi7yOEBpoA1yu8STq/7bB3ZyOflf18SFmEJPfYt
hv4nHHzRr7wW4LijbiZmpU67Or3+er7GCmxA8I6VlOo0MC7tCukJ/NUcH0n8UcDh
+0TTiNqJiOliY3O0cM+CPVDxGdOzPRXhEbU9Mhbwzl+m9yDhLci5QjesHYcHHA68
/qTSzEgG5rDCxHSuzqyixW599FGEfqHPtpF5Wr9Wj8B+cJjcmQxeUTZ896snaO4a
y86b32g5qSRzIlFY2fgMJ7xvjoz0TPI8hvKlf5x6f+iGE4TfY6w7Tnwo1XVsfdQZ
kTBL56e9vGgk/3VP4lOHI4Y/ywGghPtpicCSAcXFIqDPmmkGOMQ6mxwIxR39FXRn
EpiSk2szWjBisO3mXhNowt8yjh3jr4XmallBtMD5Na65TUV3SeqgXYCRpqFWU1hX
s46plUwNWH3KKZGGkvX0yALsnyO0eaPzh2NKFZJ64MQ2TX9QP2mCiZZdhOD7tpE1
A3rc4rutpqB3H8xowKrAHnDGQW5H5aZ4watRxm9aglQk6Y5IUa0kvL6y2SydDyn7
0QinO3TNd/XXDkB4fHMQIeu4T8RnpqLfag7EKd9K7Du8n6yYUoE0tiokS3Qa3nTX
AzuzmKxf7Ren1sV8dH8qE2yBp7qPZXXOEl54n+tXDZ0rjsy6Xl0NWjtXQ4R1EFKQ
gj16W69zeFPA15RbdT0qaH74StVAnOzeml2mzmyZiQ5HlXrnWipfyM0j0MVfbRZZ
ttaba5Muu1yTPoX+nch5ngM6rYxVLmCL13YnOHEScmFSS8oPEgzr237raRvvSGWq
pQimZ+35o0tq4+a1VsBAd+ysBQqwU2QkrIX1QgM64ksMHOGlWw+21Wto0AOJxA2Z
uxZak9nWVvFY9nXT0PU2fWaEnS7YkrMmX/mtS3gxZsRPxiBh8s/savzA0j7858JK
dEbHLDRfe6n7oDegM9FKNSe1w6pX9wgeqYDe0nMPpAaUBO1lp/ZBfe3ZQJbAz6mo
S+OtX3S3P8ME46G4UwxvJ0f5VDBFak/4V9pub0+v8j86FKhj83g++iIzoe5s/2WR
YluaiXkQCU/uO1ouJ3pppTyYLjQD52+gzSZgMK5r2C8x2sxMsUGoYcYgj53LICyA
2r97caPYod0TwPL4to8iukPlcJj8S7OO4IhPcDTnzgejNiv7Dt6wTq03oUyTTi5R
d78Hf7fhdW5WRdE6LKzCqVY0viBkkuzdbrducrsCit8K4IhMg4oZ8zFLAUcNcfs2
7m1A3nRTH3/8bR41mpFxxbZqV71BGxJBhoGl2M7fsNq7V4Y+ImEHp2JjKN7a5kmk
hYQqmxTMLg1YBoujpCP3bPL7M06dP31S/ysdlklusbf3rzUuC+1rO0glWAAaKO0O
MlCz5gI068P3k1plHe5WC9AoOlTQpf2sISMrva7f2rXdcmfCG7qk1K5ub9t2J+2V
SXxt88HsKrQk84mkueZwFFh63GYwid2gGTSbhIUprOXYXI4L3v7qRjlf7FXarXaE
NQm4gyJeqtLcqwQLZIdaGsec9iZ9Q4eSxk/TlBQ6IHzXjoCxfD+7cEuNvVMfSSbc
7mmNmhbamqhwN3ZCFIEOMyuqmMiAGbt65L8ZEvn03Q7Hy80BGUh1jNPfiq+AzjOW
HhvWbcgdUUap10Jd58SRjTqgb3k6LDLFekKfOyNvSZj3pn6bj7b2e0NJcygqoUpA
cVCcblNCA1pzP8++4XpU9ufqeAu/Oxf+2Qf1EzQO/TgdnWoznGpoKqGIfGiyWHyc
fcSiWtvnne/qXzc4gZ7lm6EKCj7pqzKca1g8tpgOe2ehjIqiIy1dEy8ELmr8YZzM
UyXl1X9qYVyAeufdSMd0R6/TQUcf77p3Ih3dxsqvZ8Kjp/sOwTNGfoEmhsrg1aZA
vAa/QpUHG6svERVMmB9KV+QuiRCgdf4b3DeGijzd/7lZr01ab7aYRquGRBlLAyW5
4nTfaxXoPxPgJ/FBLPcf88UBP9NJFBs9Q7NjVcx3A1HBFed7nT5OpY3wntC0SjYs
l8YQGHUTdfuI6zQ7Z3vbxH8EfPSnHsoySi6YR4Go2q/rZLV5jThULiBAfoF4nXhv
Bq5nn44w/kDOMx1EJm7ALIP63OmsfjhR5zMV4Enf+1fmubv5RstuqsHccc1G+o+e
lNA93Ik+WWji/y1aQnXUbBMXlCj/UPUL+d5a5mInwaHyEU4T+4lPIqlpwuZLzPkN
L0jDcVbqM1R1F7lHbyObVnycCbFhX6sgLwIqg358gWwfmKhyRGG+FSHsFueNAdLd
q1/crwZse69XbdDM5jw1TmPWekwi+RuihjMQHLy/04VPGOpbdpKpIQXPA9d3fLft
nmvdrzdrdh4xJ5VqCXiNYCnNuerUHSss9Vha67cZY+pdI4Z+F0wx0uoCa0Cg1hJx
LIoTv2z39JQHDHpn562MOGFWhoDyMtA2HzjUO3yEDJiB6skAUHAcc7kTR7O0YdVB
sW65oYdk1ZBTNSOJ+8BO/w8ngWUo1TWIq56r6KvoIiiFfi70SBiL6TismSoVAuim
bhUkB1m51yl7UBHLVkeegBbCmWMXZ4GAFa7Q+40Mef9ncmPJDyqrD02qqZZTcFGX
p3Gn9Zv8w8u2Kufb22saq7rhbGJpDaxnPx/VL0KAuXV/KjqPSXFuoUShWGqbWqTn
JPkg5wNHwKZwxONrqIqVbcIGbufxAGf0V6wfYRsU1H3HwYq+HB0JpMgsbVBRnTdx
PHEjzb6Ufb+CBogbnykm7mx5i44nbU0UWrkrV/SxG63xPGQt229ZJp3em6MIw0sW
GAX3K+VSmoCfwYBaoiKzu/5rJgIiDuKwj1aTzIYbibWSzcdRpuXECSKiFBhHl7/x
d4242pBhlF+6BnvF3hUnxByly2NQPR9neF+JP8Bl5hxODKbG7KPM7xyOvynM6UTl
VSTXbf72wYThOGQAbAQVl2To34RORXZJnuD+aKfbH3VIeVr6TKCRL6yskvtn9BgO
mgzsIboUSIXrZOx8dDAZd8ayEitWLT8ZXiUjChu8g5h7fs4cFGn2VjetZkoiqZyR
gr7B27jnYRyPLW/4YKfIyPTUDiCoDSCylHzhf7kE2Jq3Am6YmyfkAFNty8oxivAp
ll+b8dfcFo2HwI2Z5ZRrRWK31Go/tU3pewdoGr4qKFn2FANyVlS5ixCa3azqJER9
WY/IgPhYABiSAsmy78e+EOTsx/EuOVfr4kooxov6YnVVsQxPvv0oeHkcIJQst93s
TTlfBFvQR5CEtno/SZ6ajT7vXFgs5tRbPnLA2Jjye0Y31eXOMcyQfP7/VliRZ7jn
km6UzVarL87wh0Hp7nwlCvkDtJWFOQJj3Up11uE8l3CzWsmIZh0htDOxyCHottQu
X3Rl9YQDv35gm/mzAp0NFbztesjDyXucp8nNAFeoQlCCwy0giJz/eTJNiTXwu31W
9V1niLc/LMDOOjTcwZhLOk+PV6PLj9qsc1Y0wUb1dv+xVjqQ9wwhWQ97gfv9b5ko
Z9AnGfhL4yKneDqUAZdxGKqUdXdft5SnrITqU1T8SvKFc+uoLNLlHK49mA/vi+oD
aWannJlXJXG8g/ZxHFfZ0CkY7pOBz7wv3Tt+kB/rnhPPIW3KIuFVdygks0/en0+6
iYOBObSgGR5yGiRPMNlRp2/k4bQfKY1i5IqQafNNat4TQQbMjdppwhatIMSgXSHW
u7ta9TCn3VXj372PuSoGv4PVi6HGK37wWvA2fXVHlGvdzbDQtBRz5mi3dQvwx/It
FTkn37wLaBC66UlGWaxPa7mHU6qkY8+SdaE1Awvcn+kUrzGfAsOHnMZZkFuA6/xV
Ck+D+m5D8VOrLhVqKFQLOvk6AvZrQgsh/CwBE7JsHo4D+7bVoNL1xwQNHrkhJbFN
Dhxu5RwuMN6FMU+SzDvxYaxnxFibO9+GtSpGU8+WfODLRuWJy7kzkJBf8XziF/dP
sfsTPG36iTk1U6oM69gG5CqeL8vDG/DKm+NPamRvGoKI+hkCqaRkVNuSy9IQrblw
3crtxOVdD2COr3xxl4zglUyTJz+9vc0Y+suLuExOWw4xceTV/GnwmjjVOjPU+W6n
/EJUKOQtW93/lvZAiowlG5KXOgyqTauNpOqpnx/UzzPDwcWwS1SW4H6tBBZmDxWK
QUTpR0+0Tnn3Dezq1AyTTwIkx6GbujOl6/q/esj32+qvkpInRhHfYJaZciOyCpVz
O7msmSzTEJI+NH5J4VVKC0HDPl05Du+RbOXEtnz73jMjH4m04oGjqGhEpkmC9jQ4
cZHlJ1nYEvxw0WWhPAwVbCL+9sl9J3+AHRyyKaL3dccQxLvzSSvqh/2yzigOkro9
ct8+xifbkWxAgK7qh5ZKZr+MJ1hvKv7XvfX6Bl+RxDQZalctIky91SRQOZ4GaNF+
qkObrU1xnLAiGstnpV7SovdSY1q9hU0yG1kR3NPimoXX/Ibg/WgOoa91Fu2oU0Xv
UxaTqOV9wsLoM4Z3WMvxXzi5T6ikbH6hmtxmn9alOPrhS41i94YIHzLTZ5um77A+
HvAm8zEuH7cXevOIftLe9qmZlaOM+cnRDIB7HoNpArnaGHU4Cd+7YmfCj2cH0nTZ
Dc5YiBoOskTpVrzm73A2gA7Yzbb2vaIb2kkwRRCMQo5Hyf5+QbLwBI9B0vFmXm62
AT4zKJ7a8yFcASy9hekv1Elva23Q31MLkvFrkiUBl5obphE0ZG0GFRa1ml4NUWim
q9l1KaIOQifZALZ2PzyuMIC9Ci1ZsDMw8DZFYRtly0zULeBLZpcfa84hmxx0PQP4
7RGYMNG5kjrZV93q6YC3xCCBjoI/OXtf1pzUazTFCPMTCqcBSpzXUmAd1E1nauR/
io1pqyW21mV7nZ/fkKaDqAdTOfbbi5gHERMc9pLSOXU9a+b8WY31WT4O8dYC/+5S
ukshgZ5thh83Y3vqtx+xMQeNj2w01hMbF2DwlZUR68SltuWYQzGfixCLALueaLtW
pginFpboFb8P4AVCasEO+6daFuW40oXXKA1rAy+I+8OF7Oknv4AhA68UM/KNqFna
iCZ3O0AOhB3f+VcphsfGEJjwVbC042aKYj17EfYlpBNZWReIY/jC/yxtTayLlhQD
fS7YNsAliaB5r8dSgSjTT48Nd644/MmORC7WVELaKvfcDlkwpiKY8ZYQzTz9gTzd
+3a+xnC21z1w1x4KFct8eZOiMsbtOX+Ft7XHslnCDbKrU3LzQzTabak4OTRmHvZd
WaZryJzwlZOKwr4bQ4odwGrvurxkdb21f3rpPwMBAnkX16Do5WSskRkCC228eG+d
B2wgj57Gbogz34gmrYGOrlpFY3tZl48JcyM4Pd/UlND4pxnMBnwZL8Yeu6wz7JQy
7eBixHtygovWuRCI7FEJ48d5fN9zF1byJViispyn4zkw9llphJbJPdZ+Wuaao6oK
9jg1/y9Mu6U0us0nz7t7MDJ42okYhVVahE0x732VuZpas1nWPhG8bttvjF2iUBcH
y8eWN3seCEsZBAzlQYYkCCHop3OYOYMY/UMGdESp8yB123uY5957RHCM6LKrRARc
cKCKNrnuDnQgVqSqJ6F6A98lWGOn6Q1sg4lfsWIXmfu6afb/L2BBZCFDLvg5AgW2
t110FpWxjAADYe34U+d3hs1SwqbdvxnKXkOaoqOH6X4JUlQ0e86mf4vYfiJOiN5B
OSU+EWeHJl2dTv1IxqAokai7VQRggKvonaRQubwEND/7CnUctmcx6s4RCZQS+pTg
yHtNa0R6+u54tUD+/eE4pYyAE5s+rdoIOEMvuJmsfMuEzq7o6nkm3QXa04ClLqN/
kCc2GNonflc3DWhAnnFafYEZKkuKlNSk8YiGY7b7AZMAu3mCt0imuDCq6Jby8Dxz
6/TMBAIvD/z7S1p17Rg5johwJN1XIpX3RYcOTfpeXA6hNxoFdY7cUQq3o8w4ZWPp
1eFB+iNgl/izq0H1gZfT+pYGA0e6APpGhtcjzA6b96jS2Tae0cVk3vQQ7PJ0yVIu
sdxEo+waRGPPIPlA/rMLd6vZKcg1xzAVATO/lXOrM9nwFzfvIuXgDyJ6KrfjZSbT
jdQ6AWcbbarWALf5nXn3yCOL1vKQxjY/dS1rih0G3Iq7QtVBbxJhjC4I37l0WGB5
Zkcz5XOiv62m35ZLMsCV0d3ONUPec7d6X8MKTIszKRx7Zt+9G+f+IpL8CqUEHApY
U8NmTncrYLs2WAgIHBKeTvMM5aypRKXRal/ecGzoM390/cN4xGGdFfIwev+OIkKT
XHp1ZRyqBhNxtZqV0E6SCeMzL2kZr63QZbYvB6ifvt0AUdFkjmYMYvVWTRP5qDsb
7ZkMeoN3dvoKYHfFODsO4mTIBYcEW0r7rM7faCyqncKU3pHoFgsFGmXZ1GtZHqj8
TzTQIk5WBoc3/WBefSO2CkO18vhHUl/wAkb7v31Nj11HwcPoflkCG+1xZKVvlcRL
MuuYSov5HPtS95/8e8lF+fF+cUdJiHIPVoDzTgF3OyyF/4AmrmM3XddOgJNl0PHz
mOkBY98w7mjFI6g/i6pqUi152a2/9WtCuql5BROmJd/7mZqncINqfCptsq9ol5Z7
HX5k01nseuR7lt9iUg3ZPyUPayRCz+o7cyCViAYT7MVnakBtoyqF41dlPbqQ9/jZ
5zXOpctwWW3UdGnXQrBA3tG1Q0zEjYh9QtjZRKnVDZcKQfWLprNLS4EOkpCViO7l
rfo1gitHIsFC1qD9QJj31c4tcV7Sfn/Q+WDiySIJIr4VESCnBzDq95S3xs07jRdL
9+e0vP8y1RtjBGd+4LsN1e162JKb+A4WI68lmz5a1V2T7DgYjY0J6bTiNpTHJomB
zOqdfplV5KrsMYxkkkTV/ixJ6KH/S8q86/hIcSjCGnlbePmsQwvP+G+kbYMS6MQ4
yTYsYb5zHp3pbtI3OVVNXCELeAxPUsw70A+98b316wdlBPKYVVqRkyqhEunjXmY/
aQ6vgrVmBIx5L8NvA7qDxjeeFJGznu13oq4Yen0hz8w2AfIiEjw+h4QVpLj8LMth
w5rFcSjNyT3lBwEb3/ETRDZaHzTbiwU4zwkdLOx0jqXAAuaZifsioVD0kkoNJvdb
o34j422lf9FcbT6cof3ddB5pIF+0Lgxu0ZkDWQMSIjjsiz1++6UEvb5r7Xo5boPe
JhK+wcddw7E2Sf1rvNEBohhIFW7LSq5sdDsmdKhlPXDrN0e5a4XxaXAg9rfHW+rQ
pbXB6RBhnBVk2I08WszcuNpiA8hr3TnPRRrd15C80oJ45me0vbKvANVTTvueyTP2
z0e6wN154UXnOPdH3CXQr6M0GB37XxWU58CjAAFFXpf0WNUkQ5+1+tHfAGw6bmN7
B1rTUiY1UuQn3vQiQXvH251VLIfNbtwTfGEp3+MF+vY/vleAp5I/ISfq9wJIu41F
bHSHHejX6NlXonEdFAxd4ffChJJ6HipT8xOVwhUDXcZVolwj3IlAT6O6d0HXOR9E
bfnnCAA5ChHrusbm2vEjHO2XlgbyM14Ps454Iy6lPZdeMcdMpR1cUMDAzABRnxHO
zviDr+xxXxLSirrHhBqM7iPw7MXBlFR2yiyHU/cJyCkLl0T6UW5d+tMWJy931yEO
syxZs72byRXqpO98fCBjrlh5Pc6IR6yGRiZUgcKNjtQCZC2iKIuIvFat2zxpUtgg
ns3aRxTn4ayjWpKb4ju7QiYJj5HiR1+dAIwG+8AahUGwWBY3jLmodK3dsVLi4RNh
iaiFHHHGrZXrE0bVdA2nr+hx4EeoUFvAsMjgNB4E5EvcgDrN6etNZC0ocnrIHEas
In4u8y9sOr3ewBKstRjUvUVopVE2OGye3pqpyrczhY9raHPHJZR7I0wwmw63LDbH
HyBIXvSXkD8XJJ7Jy1sftc1WUrGYuWjKn5h0AG9ET8F2Y2ySbhdsGKlw05AvNdlL
q6tqDDfzwLLyymdVoYso3BN1FsM3iORVbQhIPC8Wq/328NS+rHEBnNor8picNmtH
zu7eaBmJWgOh84lyZBRA8g6maG4EZqowmgmqY4Ikuok9WKeMndC25RGWqJFvaprp
JVnEvMesOwBOtP3xmV/PLBa+PdeaaidOauq+1x3Cx7mprt/pmTtxvTHUf8C8r2EV
krKkYxMwhpARe4JxwEZDiHUFPqUaP1K5+4yRJdWXjRkyzXODJm906+x8e+SAqKr0
8RBWKP3buxe+VqGch/eTOM/k9TFw62RZ7zP1VHMfZQQv2m/jl50hho8SWcCN6lJd
0SnYypt89zePeoTurCnL2OcNa+wGOx+EcJ9SHmRw7bE8ikU2FLGzypG+Wpq88KIq
khj3PqIiA95amY/I25pFb+f10htTUVx0MajBGbOzN76P2fbcH+ACSKed3fxqMpFe
LO0Wyfg469rfD6nt99m1PqNtlLHI/Rf0O+xFP06NZ56hgTbJpP5fQf+cfT1G69zS
yvSesQ3Vfvior69+R0X/VJHAddCnsyioR5wUuXRDdMn6u/VfUDG89TiT2bVvYFOO
wCd6i4aUusz4mBd4zYlJ1Lv0q964cqQUDZQmBSSHNbz87WoOeBApCx13jlB2GQE4
Gq22AWWKF6t78a1grLB9JsZdtgAXB5bap9eag9kVN0eSEBH+Xrqqtcrkg23Yik+y
eWL74zoKs2+CSiEujDdWQTe9CcWdB+epTmj5pIFqb54vX/wnA8L0+ICwJnLvL4Ew
/Q2JRYshCACvKdEhB5EuiTnNfEnySyUZSPct06W8bxDEajH6D5gwqIhkRv93fTId
XnGd4W0f9qSSEEOCZLao2yuaEywyMf5l2b7hZGAdxk6iiLythULtupA0nqy9N8Mt
2aBxTIRDdm1aB4j4tHIlq7/l5YUJSdENmkU3i12CzeKY59YV8dXYlcWxGjKzO4JK
fGSHk2Oc7IuaGm6zsvplFonocADoz8SNL7PgFuWYD/l5/bpkVwfyf8wqcUD8mjpz
AglTdGhE2/r8YiLYP2rJIVPJkr+tWsSFm0qz8aEq7KWVMY+/ohjuGc0Mg1tbIgK9
WcHxRfWfM+EsZKiIP6w0LutCNfPdSnyZSFj9OL6g7br5Eb5l8GbUNn+OqgBxbPYl
HeLTYkGQN+nHeBcSE8KBGgGApY1MHM0T8sGRBx1QM9wnUcXPhW7cCDD3Tvmjr+Iv
rEC6yekQkW6MJwHnQ9f60mb/6B675qe1EOzsWE5/87dWw09wMGOnDnSqL86kPNRa
SnYnt4rqQg+e9dCuUCr7ROTtBy16FB8+mamZdjlzQboEJwjqrmY0plh5wXcPTgW9
mP7IijJfvY8ocVh29CFzcEafDeY57ID0T7OMpnmobIa8mBgxW0NffTF8FWzZp684
0Fh6JmUoNpOsn8T9a+rouuWeTVpoK2/jKzEURRnTs/8339hkl2KyeNlGCX5cBwLh
813NWONOsITc2DnVg8JK0VMa6Yuh55sZM5qgFqSSePsdkRbA8RnNK6lISNFTiJPa
TqnfVlx2mYOnTgdocoRzvkQqVW/ooFZ+GIQF0C23cBHMvqjhZr5svSvoada3dXAJ
FaUl5WqBAeu6+xTP4a8WM/kw7AkcQWL5X1kFGoxHo0j1ysDXEELGOQW/HgYEBsVv
nlWONSmll9AkoUf/re4vCFFRBQOmQQBpLkw8tRyzngZvP0A5RAAPIkWhQjhX8/NA
09Po9TGCF54aN4LWV0EFGXj9PdhNDObLzKmVm9bjfKkZd16kUcGf9O/tCozIZx1r
7ET6w1vFRlt7JUQKD3YjWyt+kg8S/7p4yGFso3fD9D0z1LcsIYDrCjRFoDaG6RNh
NAU4sXo9WRapmTJch7Scf+Ubv90dsSUIyYdYvgUw3DR6N5Mry888lZy0BhiFJrUt
yW5MNMQ9ePtwIwogrTPLUVAlhqIyTg4kDnf4ejn1j7Sdpf02IKnW0tlU0r5Nxpc2
EDD82TTHjgX7fN7/ckv0vxpO22kkOyjBzeqFBQNJq5QCSIiZuSkW8WbiY26GvXH+
WdOGawR+sAxjlBb+lP43OrihzedatT8LS55OAa8mm6+blzMai/DSXYxnY68CnMjB
pMI+hGbzboRcqT/gpyaM22GpdPXiB58LcAjvqqZSHVjb/GMzZNrk21LxkegncmGB
9feOtw1q/fPa/Q8wuUBKy3eLLcPf77h4z7OQsIxDtwjQMuPVAGGK7XOiuDQzfdmD
irUwPKqyUEZjclFMcYKHY1LY3IGwbgr/M0/vV8IeYCglHKOK2g2a8jNumpxJwHbO
nq6a/0wEWPSSio4SE8dQlCnC51Mf8XVf7xjEbHcunQn87pLASca+ycvSHNd+amD0
zuH4+PKzFEnBSdA+tz1fzGA4QEHTe0ytP9iggi89803sWZBk5zOwpNnbwX/ZelwR
X2gacjjfPapaVw+LyM+rw+YaXKVVQS5Vk2+4CuQsEDkGzJwrVr7FsyZVjEEaIYP0
AZNCTt4LiZGW2zzMGDUA5InXQvPuaNbFy4QNKLp70r81aW+wjQIqjq59yMqiyegX
WZiqOAaOOPWsUx6uNwxqSEmIv26U0ZPdAE71kujkUHnjXw+PH0o6xbUvCmhuxR4K
zBreKhiEswe3abNrpqa67dp0tXOzpblzYbCSkbjqj82nRp773FD5nuEutSDGTvil
Q0lie5OzVlKquJkLAxsGRNSj8PgZN4OzHVlw3De0rKKxrzVpxU45gR4EA6th50vg
t+hb5MKzj/nlgc5ZMz3hmrcqC8HNHCnbwgOA0NyI8icIEGxtwE/etuHtq53YRpJy
MldaKYlMJDSyMOaKUL6H9UNybhDpMXhRYEBggTC+3p5UtdUgcw3WQv75sD0AXdAr
UEgrNOAu31JdSueA6/rMCV4cHIT7i8EF413arIj6ztv9smh6etegv+TGxrJcIIJH
Kd4x3foiyn7z6kDuKUqe1zwvcpyJeSvXznr2Q0RU+0b71f2pb/x4e98E+1DBqAq/
g2n7tFRlTYVrmzgxw+DjZhFknjVvKVPaZORCt/0mDIc0sT17kFQw65WDLAd8K685
cSnxTWf2zJfmUXfMoh50Z2NwgzOo5/EV7oKQfwVG1e3QXez9cWorpD3CPd+drb+b
zDPBy0ovSiBEnWlnLrLhOBdvtEF3nZbQN349hcXbNhJ7RQKazCGNFj9aMKkAyzR3
4ptEqhMFT0TcJLcnq7PBFXLv3Q9UXNvJOhTM27jKqjwD7Bqrz/LZy60Z8xIyUH58
VTN9M6Mix42+OKeb7OjT9U0ppY/G8dBJMY5kx3aR8UM5kV3DDavDwvgozrsB9lq4
UuPXJ8umS60zfG1PxCkj1sKnj+LXWcBRITyR9i6JGTFpNDf5EzLRE5tThIIYsffd
GiWizgvZ9TzwruvIDEKNt554UkeqDC/zElXLshTN/GQW7+KQGcrzNXPF/DbbbXIO
80jq3s812bF1qeFTAy7rSa5Lr6Rw8uRQ7bDLQB+n3ZYphC8qzPJb4pZfozNZueOP
PUkaCtwLAeWdPcRM1IlgU0o73HsDqlVeEUSdJ4gXg7FGoh+SM0p2Bq7wLlIS0IFG
4UHAX9KU4v5iDsN+VthDWBhvKF4YEObAnziK//uSfHHj2SkS+5g4uZtENZMvF2uW
MjuxmkzGu1NVZg42RLcnG7036bCvxcrCtz2zbkx3urjTKdtslPPvjo7un3C6wL9V
wXEmAMurmFRDLcTIjCy3eA4CdJolwfpAhKFTBKmYuseZ7Xpz5CzrRh8oxVJW3ZJk
xlXnoJHjRgsx0jybkuRPnzXbTT9uecgG0HRjuyRaBhAhBnssT1kaF/piu4wSgAcE
8ZBzOsiwTr9dgUz6Ou7/RL97kVtBLc7yoqCS06j+m7yDIRwBUh89+BFs047CzMlT
Zsvq137kbzlSnNPIMqlLlxSVO7ohVOd4ouHsvN7Y+J4mHRJzWzGj5StjwR2duGNQ
b1XfIq41DgmO99puEDccC8cstrCDHyhkQ2HVk8VFw3gFrQGampVqJwbOHmuQ/R2E
J3Bib/8UIF+SgWVR2otVFEL9J+/as2s2JEDVFPd1H2bIBafKOTogS/RUicZ5s3VX
O9f9o/V3H9xyQXWNmMK6RDlatcFSgXZcXXuZQtEqIyASCErOJFf2llj7clnEG0BW
EmKwvLayE9apa9KAXFMfSFryUB3R00jAw24Z0nfTS6YafEuoLqnVf63p35l1i76Y
1nE8LqKfZlQ59upC2xWqmT34vrFnCOeBRLfiUvAKWQpp+bA2/p6zKR8e9wxQCOrj
INHIhhUsxTX5JVgKnbxND2iFJaWl9LdoZY1sboD3kBJqC4YIA+RzTrFyugGaPuPV
OxCi/9x7pmf237Ox5YoT3FNyrbdY9ucPtBrorsFJTEI2HjOajdysCN0LWe5ntvjm
wZbRAC81HjX/bHAOE3savvaACTgaMAZhYU+k8slXtTTDCwVbSRd0bd4Afvq+Ur3s
hOaP5p0pKfLNtMKZfqAg0X/kCl9DWv+icB2vtuOTxPYAGDm7Q6GrLFuhzC1jERbm
xlhIadinE84W8YN+fEG4nB1ZMIg09ylr1zuYGocCG9pCUSUCJ1d8Gqic6x53dt4o
G4uGPWAZ240VrP3O80lhsTCwsUIrQ8WHL21CHUISui0ZNDetuVGXouuq0/1NAUAA
ZuAr/2RlODs6NZ9F7rQSLHv+hVNQWi3b8NSYjwvYln3JwOyxUh3X/c79dMEIA55I
x81qQd2J1V2Db/CHw2vS7iSSeGzuD/YV7Weypx6UzDP0SP1a+mdH7bSJ334Z1FZW
0FzP4KBgsneuD5lIi6bDkHim+fCGViOcH5juEqU1Snj6wMauuxt8wbyN0+cETlgz
qU/6lrDnWrHt9YPwW4UGHj/zUGtjBt4955xerhZc2CWzG8Na4NBUjWlz8EvwfV+G
AJC+ehnNOVyfcV6TXrQfMEsKu6TyyEwaF2bs9QRG2ZArRzMOsDL4trQ3VnsLabpz
WqDIMnDLrKsqOUuS3i/U3XS0UWVnJ7WroPY7wFOAAZGjtNOF0jRj+VvYhZpa68Z3
kiQ8ZSM+WEQslzAd0h6HM0T8g0flMyiqQM9/uEXDyEGE6vD2BTyhSQ/t58zM5gFm
Yc9NuPpxp9BtCf6lsXQTGiDYRXHk1V7+sOKmfcx8OUNew6I03GwAyjpp1+8W/30Z
nAqOkQDYUYQH1RFEkoFbeHuWoW+dHiIdgJSHwv0WIuRhw4QrzrMqlYLrbwN/0CeA
8f0gj9VcEpepl3RLNvzOZTF8sx0liTLCWekdrdImnq8rTCy9pD3GOZOMVFq7s6Rq
TwSOIklqIVZvyiL2F1ttEdkeVKs2wM0qy8yc/jiEptbXWd2cZIk/AE3l+L6on/fy
A6Mt0poE2nUltZGLaPVbOS9BCduqoOjub8PvBvSv/HuvKPkUgsVVd1dg/Y6aBMVF
GkVh67mUQwFH+r1RoiM8FpZXTn4vEeWqoNw52a47hfP9bOKtxFFE52CLDJtEn60j
jPPjrtFU4ylDDBdZoEqS+TUgamAx3SwqpSiFd2V6cFriksYZGkE8Jalz4CP1aTs4
XXsDbHG8p9Je8k+aBTb86W812Mn97c//eZb62CxcjxfskIbQTtZYWOvFN40jv1/b
j/UuzM47uKD41k1TnHHDzosj4lvKKV7G3S2cidYPEuoHqbHHBQEBp6x11+3LzjDL
fPGRaVR/Bvkvz3bFQG75c/q94fifr1QjKslL/Q2aZN+6DFKvhSkIKOC+p76wtWR0
NxUBGjn8SbIQWiQhInNBtKq/xUn4y+u+WWB3/s0uXEPWnmtZGRFGp45PunSWFKN4
BfgW04b4jfKY4uZdlV7xlmsBIuzFv4aGcxwM3bDOsvf4EckgcJTq81J8U4PcBo40
BO5e3882QKo4Q+aBt1oQZ+GCdmBsIdswSyd8VzyCFDKXq1TX1UHA2A7fjt2f2tPL
HtC/xdaZJxIOU2NSqnFm2U3PUUN+bdxPk10bG1Jx1gWoXBeHdrMwaw07ZPtxuIMn
RY2eRWbxlFJR6DKfh56JD9NylGI36tLjOn3Sg0yXl5Zb6zvv0aZFrT/QgPvLkwB1
S79+1ZWd3gmSGSeRWLxk0CJ4sRFyl8Gzse86MRffhsciBYNdjemHkXX9EEDcgf0T
+pWQM/kCpyqQxPznnxf1xvtCq3xR2WAHOWHevsKrd1vYakAYF6rXQ9qhKUS5TBQq
LdSk5AbfpfjgE1WbUoNaKnZaVBRELtzuXFGDFtsRcc5MIhnBUYFbnrULJyZgjapC
qP9yGtt1u4EhSyVo3Kr4dt7RqGAjAZZ22+Ho03XbuQTwGGSSE5BooQWHLVKuUERO
NB8lKPd9ftssAN3DV7ktkDmVJOhK5j05SvwpnwnUBOauB6N7hBDalE5xzxjrk6O6
L1ahDSOluGI8szVRRiSIXo0yV3F60iX4ew/iL7SzaXY8iqWmIHkptbGgPse5VjgK
Lh+EZ/kbxYDjfXvsd6KkRcJttlNIM5XJAViBIu6mrjfsKfsb6T3rXI+/8QOneqnD
BrvkV93jfmmxiyv9fnmWw7xfLBcM0jiMOsVqjzyXCo4OmIOTfqWjq0s68HNgj+DQ
hzdnpkrY/XHFZ4B/9eQYvzUtwDJsoNXtYe771sHv8SCamLjFZ4/oM1pq/t3JwWh4
u0kYFORtbv6s3/QP5uNmq3O7nZUwJnDjacR6Bca4Uy2I3+0MyVwRcW4NdofL0yXb
KAwP9kI/SfFcU3UQ9d1RbI1sxVAT03XY+615+W80p5Bq5eVjh13tAgHMzaJhtY1u
Fs6708E2zzuQFGITW56dXyfrvYA9a+ddkMTDXPLDy/Etd254gcCyujGcspXJAESM
Kv5MWhGP9XFeC9cat1G2ScH25LRPp5CjiysDJ4gYN/jhjBqCK+pJDqyTZeNt/+kR
VmIhxTQkKm3S1IdI+2xE9DZ/LhSAtDiYoWjn+8dBaJ6CQ4gSia1d9qcLIupJrlco
Dm+6TAIo1515aWTEW5lU5hjgS6+OJBXKvB7ZB7b9i5cL+g8aeqv6O6k8QnmMz2lM
1ROYlpFPi2UqtRCVdCPJHJ6y51LhR99COnDbJUojuieqfEH9PXh4HBnQ20hvGz+U
XrNK5MfHPez9+qtIK+QW6H/sgUyrZj2NQWGoriMvrWHBdC46p1yFyHMTQqfgUw1y
pHf3X1exAsF4nkzERUqCswAtcsvtljnzGPyi8roCYv5BuOXq17dbzAht/1uTpTrR
GGDs3wWW4ICgrDt8jb2rRhsEsEHQmWvH3alokw4pKtcL2yebLYRwwqIgN4JAw9EH
Rcfx6sWTG3tIQUH0A/oxGzUJNPq2aVHd5y7dKB/pYv7dQGPzNGNw6JxnuHt+Q6vO
6G5m90+xlD9YMpODKSxb2aLQhvnJ6+BCdcZVK7LdTi/oPm0NnRBFriOdMD4Zi4vD
NK1Lti1yDFqvK+8Gsm/dEjN4NywWX/23xbnpgtrqdSLj9kMSSW7N7EjoOA22Gn/W
S0hvXrpBQ+r66ZoKGtKQnXI9VVasXGBwKilyCYt9OtBucJVBJpZUtBeG2cBHzhXs
X6j8lLG+NV7xrzSY9U8eGYTmFUddKE0aog62l/Dee07d4KhVlvhveqFexMqBZjvd
hOBlXIWzVql1zmqyzfLM5GAWkI4lJJmcaSzZZ0Yj1INqQkrgpG4rEagYzcwiSGRW
ANaVFEy3wjFsg0AFVKXZ+L9LmjoSR4ONNpBXuYN67PMhlmOUT20ZfI/Es8INE/z9
bB79OxKttQgLSMMEPEGu0M6DrIAsFEgGWUCwjRA2/Oo4M1CZExMN7ibhrkty+Wh0
F9XQqbQSenDx7SJX1RrmVRNPVD1pmE9U1e5rntjG0bivJRefyO3denmfA7nacyg4
hvZ6QSN7UhR33bTkClEsKJZhPeVFmU3CXYZchZDyuKPW5uW6Beve+yQGDChvnqOT
X/QpkJ0c/Hu9EZZ9Nrdbdhh5UMtwxtc9G0j3GX0n0HAmb9arB60rbh4m6bdTiPPl
fNwXCbIYVFJmhvfqB0Wl3Hd9sYB/C/7SPWwMlJdtMzw9Q5aWu5qhEFVKxVNY0lqO
Tvkdq2MPpN8XkUkmpT0CEyjLIGRHqlyHk/Uz7ujjx0tnLYnXo423wUakNh4D5haU
V8M7rNTPqvktRRH6R3RsTrj8WjPZEIB1ldhqQzYZqjqejEnlhSp96P876retI/bM
2kX8TRlXJrq7iN7tUVxoiAyA4Idy65i2d+7BDiTlwN+0QtQgC/W1OYX6TGXrtUyN
UsBx+wu9j6pazjwSuGZhuwNTGLr1BQklT0M4nd5Euj2UJNDQlcgsy6pMJAIHZoKs
g9mTjMnZFv7Z7UWIUdtZ9wTLX+bAbkZYafLkzzTxyP68Uls0Ode74tzj7pVWZysk
tvSV/8mPOXl8Dzj69GRQbnTwGxjavbbc3x63UW9lKJWdOhmM11m2pa8FFYb17z3M
BArFDVaHj0N07qFtq+u+buRQOcrGL/4PNYLkd3a4O9h1Cps55hN8C/xo1DBsiHF6
OwD3pFhnHQqovlVMHuExZ7WDFVY4D9U2BVdAFjmFraCfA+GgM52F5ceHeFRWzHEe
rkoDczomzfzsOQu0HsUNHmIUt0dkHhI9IjD2eV+pvUT5xub042ETI/xoNwWfsssB
ryikADUtVuMAzTAyJQMUfpzSEBqFyNS1J/ftn9/mczGMIjoYmwGeqGLYVi3BLDPv
GKwcM644xMRCPw7Us67fn0zivPHkNsYUVHsuP/HJy8fn70DJHtSTwNnXvvsITJRO
oSrx7dNWPvwHtZN+Uki0Zz4vxM/RPQwaBo/w20oTOxxMQtIQYprUeiJ2hzmLx6ww
8Pwr1YLB/E+h1oayUtAJs4VR6JX4o5EK8JZIY+c32Mqw/68vP2VHKijJVcD7s7D7
oF9vAidDb2xMCTFnL14tgPG78dSs1VVw994SGYHF1erbn6uyKMHbBWwUpFpOtDmF
eLoy4SiLGPfRVnNvUhr8ZWynUmRNhoc7pF/+f43rFznUKraou0KLS/50nw4KNfTH
zdw6qWBAnaY51faJQsChXVgJA2GOdqOehqLJbMt6DTaMKR0Mhg9jQKn49I50lD5h
W2fZUXhgshykpyXCfS6aMVHODBQ16PTE3Z3iLCpfrQrVKo+7sTY0rz/ZaxASYtcB
u5jYars/pK7QoBwbm1xWES8IMiuAJJL4ZBQspY5fQCGz6lyASRdq0dCl4am0NZHX
4RHBBbeHI/R3HQzJd0knnk+w8RJdmuHVPd2b2hW2weWN1XcmUh4s1aAv4r0bdGP3
/49X1MKuJVVFqKQVzkDafVmv8SqRuoLC9YJvolGK4ecK+n6tjDjLGciUr7MIlNtE
Xu4ZRDuRflZPwmuNOSjrwNOxPWzRfuV+8PU9DTLqk56xo8oMTO5k2KGhnPowtCc7
8NqAD/1Bm1bqtsPK7P1yCzfurzpKbWqqwJGlp6zwiFxhMMFDfj8negOCqHF5Xw5M
1/a2iVEOTjLJWUHzBVzVHf/SolSKukIQDxDcPYkRYnr8W69IYp53fqFr1daeW7M8
Ol11OmXGpSPH/c4BUqUgp9VDBzdqYh4pJbeefc0OIcnWYMXW/fIKHb/vdgjc966R
WruAleJ+HRCg2ZWKxXwKG9lqgO9qHeKN4s0+1xr1cZ4di6doH2lz+ADHGOAdAdFW
24KY7GoBgi/75cNTdPR79RgU2c6zDXrZ2stKxLEZ+DwapnsMidDY9yDqzLmP40po
L0+VlTrrIWXvidU8CbAKcmTjdYvQQq/ZQRfy6SCjGAihkhOdLOpFblx81zQqP6oz
caEyRdu3se2JLmBUP1c4QdrAJn1B3ab4wHQQahrSOCQqbg0e1h6gR4KrTaRazNtH
4B/UV2yD4h+Rii1081AFrlYmYMIj/W5wWSJ/9TdD4YMHtpsy0r1p4M2StnU3g0SC
1fO2Mp55c61bkP6IIt9n/2ymM3fPWfaNAt1dXl5taqye7I2LvMl5PAPW4IE6u7R4
SK1HVyUqbuackJno25AG2VFKN5B0KQr+gi9JGsVClttu0CmO9s2gtbKYnCedJPjh
Ku+fHHIORCHuFHPCZBapS9Bal18SPfS2sFAduhDMSX/UlQRlhPLszBvARXBTlDL/
wR3DN0Bt3xpCVO6qjRNACtfJ+JINrSHB8jolMA+JVwG8nIcIaQmiZvVbemERKEVF
inSkwflfzAz2tdxK0jVwZKBhPGoHDd18wGQ0A6r3BKonLryCdjJgj0zhufeLRtqd
GYfvtGmpAEnqdRHjVf8o36x/ErdA3UeY2xARzn//AkAeN5tqtlFD3W0FMibRgtPC
nQl9ouAHtiCqdYHFogX0LfWCY8keJnNdpSj7Mh9eBIQJkm3i1gmNQOcBoR+P1Etf
m8QMP9kY18egkIAqK8kcNsp55WEAfeZVuP+/Vz/6FN2z4QUnfzkmvwPzkY57ic/v
3z5R1Rc7ToX9iLA31Y1PuuLbnlvztkiP8wNVhIyqvkUWfsoWSPPWXzHAuJqlIDtB
T7HMTM0WozqsypupBcbHmJ8z7PDnstSRtK+VJ0jkxNImgtF847Zmr2WbjgHR9Nn0
P7aMhkZ1hgjhZURldl5fS8qGcpxzioRiSEmOlp1Wc1j88tmssigOC2DBS9lukjL/
Fw78TTW9mX7AeZW6SbUVFn5uKRO38084Mras+mwS7qwNzN+3w/CIPdJeS1L/0RnA
yD4GOKBRbM4l0HuRKTNgRwxjeKuGQuKy+XVMCCT2zebFnyubeYM3NDw70dhOQVwI
GL8MyhiddtHBHGjicAvLktsKs42UZN94pi1OHLNrITH39+p6LKQvQTnON/n+aPOf
MJoSYBZC/7Es7MlZYohKIf73kVMeYJuQ5ur0926tO+pKBP0YLneYkPs+tm5KmijP
9OYQDPoWknCibmsZA/lWojfgZWnR5S8Fjc/cAeU4a43xS0sfvxVjtsqXeDksomHP
LcfmhyqGdEfpMFO2CcNmxwUOLUz1UvIz31LMThqV97oGYU/FJ0IeHjD4/VpCGis9
aC/llZEF335WHRq2c7f1OQjL2lWXEIz7RebxGGHQDMbghLbxfpjjJE+Yt8ZV8xSs
0+5qwRo5+Mocf7fOopaDBEkZV66kd/H0Zv6SqO3vcvQnu58q34Uw0sdEcinQBVxJ
u5yUhxpE+0vHYBNSeLokjMC5uPHCeEFerfyKA+L8ZBGtjOdVyfd+pNisPd1DlhoI
NPPQgoC1Zuhdx/J5PhEacpR2rte7INplcQHLz2oIPhbpd6B7XpFRCqsKKRUUN9C9
Em3Zw0dAjdkObvmDKplTzH12UWTlC0g4RXR850ypHD/iZ1KlQkiySRjHutkyH8rc
NzhSZygEIhNpPm0m6RBUHiQTlN6d33LFU76MKevccTk6B4oLkPGSdE0gPi87xToW
i4JbfoJQcjPujHFIOBAbTNMwDFuMxnY0ZLLudiwddKddMDqLjMp+AYYun9sO5Lk+
UacAm7xbdzOGYi5wNNoiKGkXhAuDe6CEZpZObkBxagxcMB+5saJfWofPgQz6BHre
pxE4S259yHsUBJHv03Tg64kH5deUwz9qR2O3wM9i6Utny0hKuHo5WAQD+Htmm1HZ
eeGbJebZfyz3ObJBDZnAg0uIX/UWXcL5Ghr+U8HA2QwCADnzUsqU7xQx/MEp+xQp
YvhnO+8Umufdf92X4xrrA9VCsrRhLbOM3Z59+SqW4JeFWPxmN1u4K3hVRClPJaBu
RqkqEcAK57CcL1PiFJ6HXHb7buqqBZA1VfX+g8lLH2IggxoMOWRgDk3rkFh9Sqai
fYB1PsIZqk7IQ2NJdJ14GMQqKYJ8W7zvu7wRLm0UJwT7A3eHyNpkjfcxV/uv/JEE
wErUY9y/BqCbTm56pcAAJxsU0iLZF07XGBVPIByiq7h15IMQaaQAXbgYoGRnlWlE
8x1bZqmYL5HyxBlHA5xNcEVZwmt/h4iyknU6bv2bcFojp4RsOEFVyOADqmJzqwUf
GfHMjrfHeNrnt/c0ysYwUHgMV9vwmXviwdZe5yGXgsugzJRGWPDjCS4LHTUOHIpg
stbcaC4sHap+jKGXCnk/DXpPSwIE3ybG8XUSRRygVUlChYy2G+RCaTU8sJGZlrcn
1UscpFsCb235ITHWRQy/99B0lPx0vSY19+4yipjj+jXW11G/+ZCiFbvTBQ0ojkTH
7vIyY/SNWS0Cfrh0VE2qLprT+bD6IOaMRT30mJxCRRxVopuPuInbUV+DCeU9V4/f
foCZGBNlVKWO3YREXipL4WzZ3+tIvljAazTacBdyuDu9SeBE/or/P2c6OYPoM3g9
sRPWQDY7j+f199V17vX2tBspq4MLVDjYzXZVqj6LsjC5cn0x8uXhUJKx8B/TxPtr
yAIoz91ydOzT7HUEzN472LylrE+rZc1b2BBVX6yZOlQH7GCOL/Mr70eUNfOQFqLj
nvF/ERwKA2idEh+TAiVs7DziaYVHtbtfwwuKyAfzCr01iw01FiKiUjNJ6muJ0ql/
/Q18dizSExJ2bCbNrWKjUhoCgkJc3ZcVF5tGeL/CXLqljy2sMvJtwjO+ypwrwYfM
RzX70vmxttAVVZgYpUoFXREqYxwjYFS0r0I98xGoALrgaokmH1+iiTdKmXr5qBjx
Jy3zH8IeTZQQJ0L0TsBYinZRd/zecDtdi+K7o+Dj10y6LJEr4Zzui8Mydh+w6W4B
EIe3Q1so5KkMxU4SEoKbpNZKpVaBiV2j4RVoE7onvZXbahMh/2NpogE+f8tWiH6z
kMrlJAIZLvKcoi349Po7aOfwoWBdse5AWx6RbtOmB98BP/unOmokg660VjlJwM9V
HrTu8DPlHwYVwOfGwuCId/Z2E3q3ZVUF6LLCW5wEOZOdRqqk7QSmv1cmDuLHZXNm
YVfEIb/aPvibvdKFcMyHxXFunt2FXkc824HNExdZ4mPHAFgc/OvTKMkHEIrNQ/am
X2iALXmb19MfDhlZ6Y5o6c8HTCSLirXILtlHm3QVQne9s/mJLvfmAIFVFKygVEeX
e8yP3U+qDVplwwSzNwOKIrYXmuVHBQyU7QdqE/0BqqQ0Kt2Fgir4E2+XyC0CpoTj
4ELiSWgdj+r/wYr+8g9J6jrPIc9TnzlIk14ix1GjacJpuBJVZjQb2tBieR9a/THf
hu6SBpp0jo75bloXWNG8nGn4ASfq8NTlOUgYCAoA8RAnLxLKqjkp2n8awcjjehdq
cPTwEqxosskYnpgVFri82DiccZLATVAEu5eZDaZbHG7RSReeTQPZqTb1h6EO2k7W
yonFs4GJeCd+hsGOX+nnoRyQ5sqE1E/tClxFzsCp6KLq6hTm8B4KiJg/8kUCz1Sv
gz3CNaeZIf/WWSA3v1jSePBadj/HpnA8VP9u6T2euhB518V8/tsYsMahzFJdQBDr
0+D6VI+ghmJej/SUrvW43sYGh0DjYBDEBAXbNOhcaxRv+a4a0SRrtrC3dbMZXoR4
NUCZT31sGltnXmgjaQZJmrBv5dwLSWtP7A5Rp6c+G34+ov7RFM1rWSK3vs3vbtMP
w53talFlo/3jvk4WjacV9Vl4SFlTcG2KS4U6aIou3ohna1dNcxXgO+u3786+PN4o
4mwfyRgBpk93VzlFUMyoYkZy1ktAdHegBpADo+P6Ey4uHoJCmUH+IbKRCA0euMa8
+1/MVAproreX8Uu4TOZW45v0wyIgToTuhHKrSH8HSDsUmRTUTYF989R8b2DY/Oh5
dntSiNHLDmSdsj2U5ZEqyaRuPzqYWETY80gdLssFTRoMDaMKudoR1zel/wDo49v1
xmtPK1b3Om32FzGih0pLzSVMvjh4wHMygBsKN3JLMP0NK+63rv/N0ZH6kR9ab4sg
fg7PsF42GOCspHykzEMjnw4UT/qa6pytrf0ZaMJL7j2eesS6HupPPXQHZ0BvEwEX
lSkrNvr/CpqDVivacCRcwB4LS7iefju2eNHQa25JxkhvcH/i9fzrEZ1cjBY73rHO
J34vYqOLZKmjDMCJLjY5+gGVg6yyduasCL4AnxWVXVCywklWhM3nOEqma3IooL1J
TA4XcsPcjInJNELqQyN3TvK524GgqbFG1RqQVA1h8dC1YpqOeO1lWUbZ5YUAoab9
wLPISUp4USjDsNkHEO0kzdENLmWP54Dw2r5hyrKDh4tDlBlXFiH+GtVG6Blscnak
OfCa3Kk2E2ce3KX8fAKBZnSq4Ame8OEnIB71GpZPFXhIeJyKMfrL6vqOgxYvRzQk
JhA/ctJe6Qggy5GOUlMDN8IzQoDDoPxl0xNF5tLFKBxtIYNhaPkCL6Up6i57GQVA
VM/TBx2z2SfmAa0ispUQZzVO7U5ygenxaGnvZLfcD4xEAlbprwcfZBOe5Gu2MIat
7tvhZXVNFPRuQgfE/alZks/fOag4GjBVM2p926mIIe/AcqlmVs6d4kLM/zo8wVyz
nXDFd46ZMllokVhLdH/dRmviNuF3p/KSj+VEmzNJ9eywpQE+pX8MTsCkX7cL5p6E
yaDxHle1nVcX/AN9c/UKKLxbcy2v2rVEXNeqjFVW6uaC1KE+IErUYBXusDf5sryV
LZCLptZh3Hs4xDkL7gexGUqDBED7RsErDtSi2t4rnxTArRLw5d7QAECAGwEkXTbY
Jvn/cxXyHge2NIShORKxdi1OttCJJFfJa9UxrWBkfM1yDZlonXrLymAweNVT5wjN
xht5nFRBqXNO6AdCtt/f3Wvp0AyLDbOKO6FigEphGBnnyh6X70eKv2iF62RKa8qH
ofl7E3nawU769FOlj3pCTQmHfdux0qYQlLpUz79Kcp3u0IaO8rKJ5HTERBAoNEqV
OyMX33GM4VJ9EnStNI00ORsU0x+3tD0VSkWD7JTeXx9TWqy/lAiRJp8/+Zj3Rewp
LtZD6ZelToMFVPIXx1dKqwdI0IRrYEk2jCaiIKUnu+5UGygP6pfJ9qEa65UKIugQ
3bMtaVnCc5FVdwwdKFaz96QzhfjWuxi4POhIs8UxwDMPO2R6BU7OZVjE/KmBjUER
qD3ytxakYOg1tDaDC0o3gTjr6lDnmLLWLdihx96yV73gfUQBmF5WvkuFWq1Tul3z
GE3ceRnKU9etehPOl9Kj3g7WWMp46zOpUJHJyeWT0+//FtffS0JQ+SP9+omDpif3
GyXdODVzBGHxyAr4eNVoeNoqpjhmI3tcYVzYDg7fbVAdD4qXc1tv/Y78xbk/xv09
VGcZfxMUguyHUVZcSYS+J5ifYMirrQbnCPzeiYfHCKz3nxdkext6npepynnP8hXC
RzAMFh871RdR2SMQIYflqbqARtsvT3mdJHtDk2s0jHwVxBFifS7DO8yC1e+ryNB9
VNV/p2hzbzAsSL4mIdrF50/9jdU4hKs8VG/GyRzFxVoCNc15asa7RNrDIcbxP1Ul
/luUw1mZsvZGWtU9qSdmN1OEciC6HrI97i/ipO0itFHaeCGHg+oTDdPieGsFKSjx
bXZaVmxbtI3FrPjNxTWZZRMZcnufM+iEgRa+J/q1pyl9fwj4i5BIKlIWqJZoggRz
yqEQjqtnqyMttYa5vb5obMlo+dfzR1zLDeNS+7N7SmP4XnSuflW8mf2XmyfZBXAt
24S3Si1l7ryH33mcOa7Nknt+f08GCmqsmWClT6etStfx9H3H/Bkso0+wibxUvQvg
+N5Si9vAS0AAhnGfAcx1Cog2YekJXH5OF2gU3krgUuv2AZYdVFNnPKOPG/AlXk1u
fj6F8lmTjy7lrTf2POcDXKcHCDyL46kWY3fPAU0EvvEhvnCzayod5tMmHe1IVauY
Nx699KrhsK6bXPL6tyM07IeWtsAifQR9ibkHSWaOZBauYr6gRK2LWlxE2tC4N5Y6
3BosA6z1eny0oSJbDL9soj2HKiqEid2AvsocAkY8pYTvCYMwaohYOLmlnwfwLiie
27TtdC7hbZQZMK22IiSSknro8A/tlaU4VicNC3cNRzZfHFh7yfdr+wTxP89ZNDDV
MrzSk80Imlb3bzpwH+96Y1AhINTkgtWozl2E6dLV0RPPDDXRRhJtq9zSZDFwjPBB
T6EP69w0FoEAgcw9cSlrmnJrQNXTOekpCA6adukbcogFWvXD+dFmZ/gOgxoMVAzE
X6vhzofyiBwqpdEgod2GSlUi6dFJbhM4ibdyV2Z5a9jufja/+R8KbmWVPjcy6SCS
ubf2PIx24ywFWpt5kFo/hSg7yLIyKzXhJ6VQ9nv/mu8T89RPrlyAg8tLP7Teo4ey
za7JdxCS5PmEAo2ah6koxqp+WFcSbWMHZyV3n3RA8bxjbjYjf80Hdu29lLwsmWJa
CzOiisEkt8lYPytRsftZCJEzy3ZHUi+8uLjedXO27VbyqtOCe4GGaL4uRUHU7h1e
1V2Zps1eD1tMPvLjpjrb94D7UsW1ft5EBuzflr3owJR0+LQ7kSawh9EV5p66C9Kb
WNhzMNuOCMqTRI9A6JasSrXfAgJ1lIC6H2OitoB/QsZ9q9Tpp1nHLHN30gcbhMGZ
duwkDZTIGgkxdBmFXIy/emvEXg2m1aY9g0n1clhgVb0Aa8s8c8T4RulQiPUjuSro
ePHn6lQJ+lKUOqXcImM7dMsONWodKEy877lm2Jx7yP59uazDeXlp2L7C4CdhIfm+
+TMM/eCBWPJXSwqY3h1I830sadn2Kqeyg9XjMgw1wjcWtnEOLWWJ/gqFgA8dSHyw
6s/g6D6LIDghIpE7CIz1EsrIm/s300tYGfQk0dvvTBviUF6O6FiXNf1v7DxY/dhP
KBMjvH4EjRv/Ab/nQKTeZE4zodOsCs7vcr69DGFEj69DqUA2GBv/PatUDc2xmrRe
pZ/hDJaWGqcNBpyREm1C6ruy97Tv9ifrSfLyi4x/5WECdPhplxPaBSCMJoOOXISi
PggnvhP9HYsnyBztd/7tihby2EbeiLmCszVqpYie4BQirvy1i3gwvlf2xhncTsVS
VueI5y8hqWUoICrDKB2SH6bLycMUTgDV5BHlhyxhKcdyFfSQ8mZSs96oHlYGE1Wk
rHQb8G/KD4SAlwMwEWHVvWaquIXr/7hIUSXd4CvVhdsHWivIPy9OP1edERp3IVnn
+B7GKWV/FaujLEziScZbC4+Bzg3ofTR0G4kxjsEoGKvS9xmaHfdGa2N6AXIedkoa
R/0F2RRqD4VeKrnpDUrvkeeeyL2oJi4S0NvPMfaIvWrwaZi1vUTaM5FirlgTOt/Y
DPRQMzwy/Vpier9NHkY+wGXNeAaXrOs7pUeRKTx3bjDpRWSJQMfajIQeQRzJBSjg
MfmHlX18j2ikDDxYFli8RVOzd5Lnlnuku4XUigp1xLbTYm/3z0ET1D+a7d7D1AHt
cR3Ha7Yhs8Fas0fJDobO2xjvMOLqO1EcISPw424rf+s5Pu5tha8HoLyWEJsvOdjA
OZn2JObOgooz7q4+nTAbDJPcxltn8349UGPC1Q6XQ0hHhvgJTlFA4KRfoCp1nLEi
Hn9j7Jh3zmC5BKRSWqABKgPrhrs8VbtqBb17SRdbu7LnscUqHa/Qr6WzgJ3s6ZHW
4qFqyHHH5mlglySv4ImWlaJVqgSvaHGLIlZKcjteAD3bQMaFta3XNzrY0X3+0CEd
jnoLfodytNEgGCi/1Fn48mfuv3sm1AKCr9RhBhr6l57h2ycjcCPdQr0rgJEAYAD+
L1JlcolN7Xs331UR9GWdbTArbY4gXJqSzYtrssQeyBpy7rMfKwcuZzXojnNZM0d4
Z3lKTCjbShzcl1ZyFrQgXoLbOpca3fF1aDzKEdX+UBotkJ4NrOoPSJL3WC4b+VfQ
7ivaT31QUDV9hGegBH7gXsrr6aRgBQZt10ZUEBbYD6YnEDoxgOxg+NxfxtDy9ylW
tqK+78ZuTyC7LudLUrsyNueKEyNtNIb/YEorJBhyh/yugxCCWp7oWoDFDy1M7SXr
KBAG/qJh6b6Ur3b/jZDGwS0JxctfsAJcR3NLMzLGHWqcw2wSdHxrTPdQ9oQDzBTf
H3s+KLLetKXpIWwscPVFe5RSviazrsyPYaasPzZ4l4M/1PyGVjuwdU/QGUj6n16e
W8Fz2e8mEIcfMoSXfdMulN88mH6b2EFSp+vWJDxGt6W7CS5iP14VrVus54a2XWiW
phtCGPFmy+7FcYtAZvRaxBsORTUEErUDn+nWsDYk9aCB33AJ03vvhTzhaNZBWlJg
iJ5dXYIKLOEnjaH7rUMUA5/i1QXAm+cabNMKiUK70QMtTBg/iYX0NEJ5UsEuL8xA
9k/6WfVByeKDoqTnFqroqQwSodkyGQAaQW9qwgd6xax6I7WNjhS0932gW7KVAj5j
0zRfs9ILXrNkXdNX26M+4kyF1lZAjILSpYYbamKVc50geGX6JpXk0OSYZbCN5o2m
Bl3rEDSlHgkeXzgR4BfUJGUSD18aF1/vzj/fuiiliMvL0h6dv7iL9cLROMq0faTV
PXO8iOCobUtzn+RmZQYrzFJDZ8GyIOg6dfV1fPAWzwEuhiW1HwZRF4Yw4i67aLsD
fnaQVp92rBbFG5WPgJ9HR7geJAGWfkJW6VO5OMXzH85shNTK4Bpa7VE6aRhQmMgV
TIpu88ijcUeYAJz1w2TwsG85AlaSunEX/LpKhBdf+sXRN/jfnrp2IFpM5mDbyQYI
Jn4zL57vg15JE3KxBi/86BGkdDpWdpAqs5stZpNdRMfE/t8K/i+lpKarGPSdaze+
uUxG+0wqmqlxFaPxCOaQc56dAp6yPM2OPCj2062dF5Ub5bABdbQWQ9apL47cwftU
6j0qLnyuUD1faXHxbeqsAfb7x/71d+UOFRu/QbmtEWYwru6OLc7dUOqy3tnnLThF
T3/5TWDhsILX5wdbphaz1YhN+Y+rwZfvhYlZJPb1Sd4n/OACyQk5GjzWtZeiaRDT
ektOe4drb2SL6v01PpUfqzS3YFkLnrquFNkQ8x34WGLxyYbBM4S84CkBERFw9Zul
Izj1aLnk0RTxqDA+eeLxGLrcWC6iJU3lMyg7OD9/5tZYhhgXlt5+auLBEhY/CqW4
Ih1k2NSbXLW/j4N7qlDGPKaR8dFua99S97dnkuY5FzYpENbZldblpt7wL/ci8Lj4
WCNIF0t/zA+JCaGahcgan3gEc1WAP+ObPyOB17D4LyKrvDS2/W4NGMH2NfsbAMex
VAzva+wn9r5K6zYRqgc4SXnJrrKF89SKSOKdM8QgK7i9UK5PqWpsBXBHCbKvAfBo
Um7+ImedC5Z0jub/tP+5nMicZuxzKOCrt7aE0hC7E+pLUpOHZcAhjQTzh/Ciz8fX
eJitn9qfPpHk8H7eCGL0nwvg+2hNASiHt2FKlJBRGtmXiO271cIl90rGYKMMNLhX
kj1lOOvZLsO5+ltm6HvJWQ59yxOdq+jqZ1D3OFAlLpxhYXy3Q6Zse3Qsz01sMTJ3
xuDLQf+/0sUkJRBdQ3A14sPntTPpHqJlsp8r6SS41+lz122I3WOiwlsDFrw2tBPU
NKnFmf+dud6yUIMjeLICA7plgF7j6p/ASn4cTisu/sZ1i3JA76i0in62f3WaevVD
nSlCoJicCCOg5WF7bqNQaEqHtKtSEuzzxHC2Bq3f/LUZeN/xChM8qQvilhJtSkCW
CB+OOq9qqpxpZr49cWC5Ap1y2/r2OZ4eEMkGu1fKaOEGyoeRSkpx3+w6bh+49Oi4
Y36DuyXMhyNUGJHs+IS7NN3yLwxm3ZF8lHmVWWdXURNe3K1GQ2GH5ooNF/fAjezF
MVMbv3FZ6qKm3zWeRT7fQ5tuOKWYZUz+kfht+hAEkW+KLv77ymx7d93lCvWKBvCX
1WYW4T06xTGmprRij4w5/6XDgH5F6RIEKcyWpJo9DyjUaKvRST9RcOuJBiK6Qxqr
A37iYRDGGGJOOwQCSFZl6uPNhjqCBn0otQPdQDw0PPjOy1lUHCW8CPWvdMB810vu
KOj7DN/K2H357PSPIK51x8++h3KR7SdqAjHsSOsjqgSxYO4ZlV785VHy4+UbSJso
IN87F/qTOumNS17uQcoS4pJpqJLbKZZpUfIJpDUnHAVBfAVrvqJdj2BqYJjL5yJM
/NRgovjoVdZ5oupkajCm4ci0aHHB910uEhpjmZfH1ae3Qa/PyF7eg6Z/awPRdrBc
rkoRHfxw08x4sIp7GGEvNbD+T+RsOWtLJKMgn1TV9EhukcjXY1Q8TUXVsciT9FCy
nyeeFmk840ymcr02K1TrvcZXZ5UFgcsCemr4AmTa1PvZlMn9kN1ZhIcf3fIFb8Tl
/C/PCshfYZYBL7OQlGk4n8SXm60a70vLwyzmqdwd9NqDG2mONM2MKxsfd+xgiJQA
UXJSBtptF8kRMbjOYbDdt3JXWaj2sjYWol3bChU2RKF9KJYJsFIYMB+Y1+QHjjyh
i3iHAmBTOjNE0UCeVcGZ/lGz1M3zIa7LISsjSCV0UVOLnvZEfQsEHlh6sLLVuS/J
9cXqb31XkjxeTWqjZB7sEvAubGth+DsJk1kcCiqiZa/dG/A7rgd3cC6kcFxmV9rE
WKrw+N9OOm7GHZSWRjo4V9XUuU9G80rO4oHP0QERr13OVOtZ7OjOouKBUJoZZWq4
fHw0AGfjOkibTWberF8QoycILL0kpsOmnDHjYqpGvRT3QMmHqQkfnNgPuRonntvv
xa0uZdPtwCx5abcOq/zpzIx38F5Wi1X7bV2vsemg5r/6/Qr2O8/gSUOVqafggT4A
GE4gKOHZu8E6zkKmUYT7NITrcyRsHyy3liObD/aEbaMIg5NtH2OZvrJ5HH//5TTh
nYWV4YD5cXp4WKik9SekrDOee7fz48v5MTPP07H2w7uj38tchFEUPK8cY7wFXl+P
7lJWiR6DLo8C8OVQWdbrOfheHHYvDt8yVWX397k/qoqVcRTg8neOBq+7sl/aHmdQ
BhLDky7gpGtypxS/SE19zx/nMXLOe+eN3FyYT6IA4nHZuqCBRGZrN5O8RfX1n+1r
iyeYcirflFllTepi5RgWGH8VfvSos1hDCK8+uzmSW8r4RoffvvCAF+hrklR5gvP2
ZowigWcCYibb7B7ZGAtWv157OWPASzVc2jAOgkEx8gFYGX5MMFaf9rHMmpTlow9e
zKtWaDiXaRxSXjZ38F4z/SPhQ3Byohf2zUbXcBxi0SW66G6GsFjKIVUFt21X01DS
HDW2QnnVMqIvB/Ca0f1tU/zinOkpDzjzkHLLARRybZrYZ+nBZfB3eqGZ2UE6BsOf
8zT44RWVNqjFMLlnRVwrbc8u/Z4kCunMZMF0aosXNdQ8eUf7UThHpoAI5JZzea7R
IgzdfiRejUAtxzEZrxr+a8Or8wrt0/oBRjfOawLCAImrxdXoyGqcMKkNKGorKNEz
/IYQ2FndTZ0+JXp1SD5m7Y7KqWvA6DezCeSdbGgQb1jIYJdGOXk/Bigx/jjXacUp
l9wTW5/zi7jxcCe4o8uoqacaoq62mYKSgj9Za1rzgihrE3IRRhtzNS7xsVPKFBlT
/KlB9T495l4FVdYZOkpMzWlO1VuLtzDPtWlH6BvTLCALLlGpkTucJa/A+BKOjwIa
a09xhe3nuRriNk9HTgpeLnglpG+1JoxYcyiyPxCqY9cnVeEyoJtwVERatS51+hJm
xemVeThygvb+0ddXjQ7N2C1wiJ/ahFDu1iBpbnGmoxmZXDKw123kSuWPLMBbpR2y
wu7y77C0197ulIvB+wYUOxNsEU2G9jUDkGbQ+BU/j5I/8Rkp9ZxS0ieXwRHfoPUe
DjlXwx4R/Pp011KS3SQLMlA0Q6TF8uSjPxiGlgnV+iIZrZayLuc9UQSEi86P9lWx
Edltxsp40jhx92PKSXvh0KEIBrfBnUvBHLB6UZADD7aZWQFRawRhAdkGTSOptivL
Q9vxko2GIxcg8aqPPtabYVI7pVKnEX6ZYxnmyGV4qwMs1NkzStnQmA9o6j+lUafH
p81YAmZMxqcRNZLz5KQ+9ZfzDKLMtUKM/Aro/OggxqWZLczwrmCYRLPAPiHiihP0
u7yHB43IEn1+buUaiMrKziahMq6m8ofbq8+t2Nx4xVod9J6uAiOLdxwoiG6ETgR4
RFARfNDv57zpA/U/5mxZws4hpoghby6FTNwOyZNCfI/dvJ7BckaTxrSHeWNC//6N
OwFLy5A0GX4pE4f/7XiK26peiwBMD6CwnaXua4yFjB3oOxs+h47g/9mHVG3vrMaP
S8cgIiyQqjm4YV5eNf8T5LgdWjubjXAjPrdNlSlFK4eLTfAnZb4Ba9Bu76YXaDmA
cJsS2Llkplp68pt8pOxTevXIv598KxAtcLuwW2QSuUS4ayvxRZLO/l4YtUcVOvZ1
FD9aW7BGtJoa7Gzt0x97n1o+ddXK3nBMmwuADL5OwyeTre7/P8nSXngsxxd2Bxy6
OPqTVsLNXwZxnR7IE0dIyiUcK8bTwkBLs8W7ICx6ONeWMXUAooGqI9NTTzUB/+b9
7lbxvZxyRO2NSazZD0MLH8HfgD73UDv2pvIBtMrG79QKDbdFnnO34Zx751WaUB6i
MKg0dJvNN9ItG0it1M/Q6Mkthgja9A2G0qwWC+ntKPGpi9d0DouE4CSC1Ca+em7l
7KR4fuCsitqIF4N0B/HxMzFq+lmB8K8fXhHlYPynSL45vR74BhoFHX/1FSpAX8Mt
KwA7DVF5cEPBVzmt+49ZPcw7XUQ8hnxXFoQbxyspt9K54rcJQKFthXPtm3FjvZ3o
anDPEmuo+XCekM+JtYbOqb5EgvcPBmVzwlwEa+ikI5xAu3uKT9KnN2p613CxFb5+
0TCIrJ48VjhqwduUcDgqct8A8oyWCh0+J7Pxq0Z4DgRBKHS3svG0S/hv3WU9PSSy
pLpjobnXzz96JhFrHoVKks5/yvfv7JTzHn3t5bT5O5b1JQPYGnub3zbUaoB1ajRn
KpFtFEQuTace9q646RY6dC1XCyjbU4te4LWAHdqcHchOYy8bOg32Y7AI4wJPBnnb
834bMKPbr46vT5wul1AdCOIqfAc5P/8r9xzLWRI4dzoCHcmqz52WTIJE63loh18y
ZFo6QttJpRcalEsLneYUK7RKFcMoVinEdvmbtBamdWK7/POXeVDvpqq73mMETaKO
VRsEdFPPWrAvVZlqDk9Wu4RFP2+frDom06yf9QKU/faGakdotXioVxbUNF+fpqOi
/MpTBPASu3fUCYFOrEGYg2zCpf2UAWTyhU0c5wVUW5chDXRjDnZIntNIUkTxVzaS
6pqChuoszeK1YkCiYwCCh73NsfeMYeiTpKKeTfu8Iu0AmK5eM00mi+o/4p9+d6UP
dPkZNAjHoXlEbf1hA/Gm0RB3IBEoUILVQCx5T9R6UPgCpcbOX3cXWwVWoTvOjxlj
Rus8pqKnTb2Lj9wtUr/V8ygbie5Dt3K1p5djMy944WiK/Jfx69FHelOB2ZLVpCdm
DI3A3ToVsOwjZUkJOf7GEyfLD9pG3Iz5GAsCSMl242XeX9gbC6P/x3O4OJPBBVRm
bQqpaO/V8U1Pusro5AEbgL1wmB+z+vwDMoXmI1metjgCGabUe92us9GGuCALAvX2
zfUYXT2EYaQog2zBPbs7bYIibZd2bbHKBjjj71U1Ek2AuGvFY7o+8QTU7BIDo/Bj
I00OIQd43Ui3DO/OkKBfHtXpAytyWgkAkK6Jne0qrKfwS1MpdiWVAMd2rlQeG9d5
wZ7rIzjux++IwDmPy++n5cXGInO6ZVEtkfvWumqV23kuC4vQO1jUBHuHr+8IjNW8
ufdYCMfRQDP7/4nvKITEXRdTUstNrPJTURGUHqz9tB02t4eMzq3XDH0Jf/+gyzpc
iWk+LKUcx3JS6S6f9Njcn1u5AGBSBYEadgxaZrxuBOQAU8j0kXkKQFupTiPVBX1Y
5Z5O1PgWYaf1XVbH+cofPYpuCWl0uxFGC4yMzqmKwKNldray2KdAFNXPjNkGBiKW
Y+vv/jgnjlAIpVnAKEPQ3wn49gxBzpwXMchtQ8dFIljBq5PDeKbvvYy3ApzdLgb0
/7Wa4eTsYCf/Fwj7FJmf+MOsEXCxD8Iw8Q3ZC4PLeVq3erIbsToZTHtAXzlhtPPt
EszT0czvHZPK/OdrFIZUh/klBBbXbk6MctBzB1sqAi4mAQO7ic0D9wIwzDi6oZ7c
AhVdekK/MpTfij66xqGTd+ks7Ww26iVQhTtJ856lVF5Bh6etYuTj3lch44CgzEBB
pc7sIjyG0vhRdBti8d+Ivd+c2Sm6HqSvn9shEFyN5CsuJlp71JalqRednfezpBym
Y4Jb/+o5tWmoHhb+CBhsMBAT/NglEaYr7A2Di6S9bVjNnbto8/O0dNQn1Q1LMdWO
W82XmEu3qwWf7UxWpgQfPMcgq8JqWFaTwVZZAMvO+BASeBNsTHSczySAr5iyDtrZ
7ic7e++Yp+Xh7YVD8mHRPnfhQUPVwgpel8xmA2SpRe2J0zhCVK+E8EtY5B97fwUv
4X9AOTW2lrBxAluES+DeK0IogkYA2Mm+boaOxhuvkNSfRMfQZF7T6tLZ1gwZfgLh
u0r/g3DpQOFMKf1nGVCnOPhJGNpP1HEN0P+XbekZKAQvcO8o11VZ6q45/Wi8zFET
aKqvvj7SmnsuVqLz7bYtXxmDAxx35mDuShk0OoJv7mHgIAFwkn6BiIzrcClhBKWn
SRQb7HH+8ykjsju8opTxG52eESLz4c4Jm4Gf3SL37eZKQAzqtc9DEb4Q8mv5PsX1
IR8Ll+rarpNFwEwDqFxLid5YQyqHixKoogjBMxLcrXnyTBS2D+bmdGTWrtsiJJIB
fUQ/g4CIUyVzIlPS6c6PhDLsnUP/vQ8LB0xERHJMQjjYwM5EIqo2MLWFPyFfO8PG
5xiFb/u6op1OvORFR1fFOFpingfX7v4iYVsWJdB63aBU4LXW1an5rmpDmNGFNVXZ
ZQqZWv8x1r1Rr/w3y86li5KhlXEQ11TZPR/c04jP+jr7W40GdVkfGHRoA43xLPSP
Zgubc445LvJjxh/gV8kFwrxNey8hVoiKaFtwlgrmsIwk0DLNkreK3UfGbX/sRz5n
GSkMgutMwvXEJybNxyFkWhbgEyEe7IpDUkwjdDkCiXDkmLeVIsCFfqSfINmn/tJX
2a1SFmxG0eh04705hMLDcyTjXsWsStW9WL60nq99QUMYv6ei57klfQAgC/dV/t5+
4OQzeWFcYaQ/xB+xmdhDwKpCGX16e4qHWUNvLJjMA0nh5U3Buz6Y5UAZ4z+2h/QH
ERYlH6oi0bXDkT9rq5pWFZ6iz1VDXhfatd+JoQoWMtQDaC34xeXeuCqCt2RG81l4
XO+UYokzSwaSr7rachkqPaWtNCPXvfUhgDEvAWOtJ9k+8kzR3K2ia/d95lfNU9A6
wHNiGmIjeUiRgR/tQ1Jur1ZzGLZ1KzeXSBMCFlTJ+Q2znOA9mOqrM6cUewXpbE8o
r7p+KF2cPi3vIJM1Jcoscl3oXUri+0qu55XKTUyLfKOXXxeN07tO7CBYKDA9eKF5
7+3WCYOC/tdn9VhStjGg7J2KHc3kuv4ahvRpFtlnRFr2aUfkU/n2UlWeu11u/KEq
nxEYP9DxRyCYAzf6W4EOZJ4Sw3MsMkk/gi4Bwis0Y2NziEe/II+nZWXuIcqu0Mir
T3SlJ97E2RqNDze+Yg6ysznu0ocEQFTYeczIxpSFuzxBQFMTBS6EOG2LEYkeWddO
yc5sCvlhKbJJMJXeqmkizGTEXxlLPoCWu1F3F7d60JDLFUGzxLaEsIRk4/6CNKgY
X8nDgCbCpgMkPRdid6yUMCh6XougnkogAfbhdIMvMAFpClqyQXXPwdbDFg0MUEK4
XOFxUZmz1bzDoU4MWN2sXEKO/Kx7t8QV4VlfUlOnhhVXzwSnsapR0OMkFAVyUYyN
6RiiXAhNv/4pSOfeVwcjVHnUuVKPzYvlW7vtI74XgS7iiqvc7YzrPOzYrX17mIZ5
574NcIWO16JVFEa1Q4nqWm1Vj7zmGlOetQoSSo5Y5hx+PzBx5SdLiYKRRijEDvk8
+ZefkRBquGvkkCZ14EQrDleppurlosgskLlM+hozOxR/ZwURWpGzFbkx9sJ0oERT
GKp5hJU6EWF68Itw/uGQa9JVBaXB2I07fttjZUKzRi5PEuD3I+l3LPh9HkDiFDbJ
Nd/Vt74eQdyfEd++GZ2biG8zNsoONLIQCNqovKUOql5ilU2ofOil1506nvZAAYsz
Ck4Uyn8sjcv2PETHCeUSdJZwL7WOw/aIaCd8Op0p+jHz1kvfiBSnFrrz1T1Iqx2j
d/os6tBtsmm/3RNcONVIo4M8wuakGjyQGM2qzT0C8sH3tgChSaSeRiur+2DBv7dW
rq2l8HIZzMPJ/5tMwrCmt45Rv6Tl+l4y9o++neeqEPk7/fWDLHdmHkmYSscSyHDI
UV/RPKYLcMz/0SIzUYZLgrsvLKaQD2Ghd1Fw50TatsP9A1YbmexnYykv4i/FF3TZ
sYdq66dFzVkQUVv4GCJR4Jg2UjYeBPYE/dJcvZIo9OTAI0H6QoUqHz/MM5+tjSTx
3LRXjUxFPpDSIP5dbjBbrKpIgJMki3N+6bU143EQQ8YDapq/aUYl4qNPBAtWPywj
3IVrqVJQKE87wgcl7CXfmlcPmtkfFgDuNxI9PIY2LV6GtJD30MG6Q04kvn2ZFsBp
5tjFNKEMWN6Ow26SP+ow4Etuf6rQeCfFs2qlSTsEa6SvvK1ZBcqUALMFqsptYuCJ
q+5XRnyYfgmVTLb6of7HlHxrs1pGKnvBxBefBZyMPDngU0yinViLn7aHLKBSUtlm
dItnYkEIeCMHULaM/N9DbUCt/x9aoMm2t01nZbbFB5VLgv+8B2JMU8K66nTaSQsG
se2Wyl7IU2QO4+MN1eyoDBzNXupf1DZ5EltpHMR5oWS4Xsc69rneyRLj6UaNQqdf
UCxO6vgZJU2RAN/peJ+xS5Balv5xTZsgn53tP2y1qeN02cc63eiq/JhzXK6Qp/Fo
7tKpxXeB3/UOk+b7j/AbS9GUZSi1Sowx6PcVQ45K8Gam+wYU02zRAA7/ba1Fu1DR
MRAJk9dScm/Qnizt4753CdokCWPLcjUUJfqpKM+hqYX+YRTUnPtmtP5l5+wtnVkr
7s4yBaIQeDl9EnO4LtN/xWaK5rDW0WCybwoh2m3YCWJ/cnBQAbmhiLp/0yzEmSyl
EPFOxb47iVoKCY8cLPdkkUeKXxKKphHGIt4RtECsG08p6B2MumhINnwj3Y58CU2q
Pt8Z9XIf5HK//LCg4uZzy/70v1pEqsPmfB4DxGSvN5o6c1dPwJKsIg6O0vXa8vCY
UV2xA8WJ61A/+gCROW1uHtYCNROn/258I+5z1nOEn/UYDUZBVYpkboNpVHu+BtD9
y8jqPiuwB/0La6D9i3tuyxDC+RGa6hJuj1E+aYp2yEcUt2gs8w2msw1yyybs3k0U
tOUxGgh5fPaHRi0NLdv2U+/2bpoMFNKzBSGuS2Zehj6wJC47CzpmUxTLK/U3HzS2
zctLoAg+C3W84r9C7dvPF+rJoKmjHX4D3Wsx4Ce/bKb2u+dl+Z2LMiJYN6xrz5Ap
4V4ghO6HSar5Dqil9AyhX9/KA8N9t8BEmekdxlfdlGt6daaZxjkUyEPUPQZaGo6F
fPsjVpLMEt3ze+5VISgd8drxKkVBdOwjsy9dI9uDykbM0hU3gy4vsi0YUxGbNZE9
frHwjg51tMYNz4gqS7W+zHUbgoYjQHgXK+X00WVRn4ORTjJOW7XiekmgEGcNKjv2
V/7kuecOW7D3XI+58mPqJ1G8gFXwDXNhGHeQExLotf13ivwrp/2hWaMtlc0Fas8G
YH4Klkaug4MNgzTwzpeNmIAlJX5jxk4TDV4QAuliktOpLP5cKcb9bVGqWf3r9iiB
D1+EhrD/trWH+STwxv9y0yKGCAAjw96fd/ju++Jq6o7qYHADVbZTxBrWjoPDqEiX
mzSFYBB6NlO0t4lFKwovQ4/z3qrNY40G4pPw0nhV/OewitqoowL5ZtjqzxRJJpuy
hSe3X8Ss98VF6LCjp9HmEJFrfSWBt5uKod/uNBEsvsuO5EvD6OEQkbJ1UX7Kz3Os
sgJqPZANf190o6i3mKfzjc8VJ20xLxp+aaUTpyHQTZeiqiEoqhYOvclm6TM7FbSt
t9516nFmXjDGsD8VYO9IkMnmVgE4k8WeqH2S6f5NYnK3maamfs8JJRbW84pdyI8T
dyvWYJKHIX6yt31v3xJe6bU569K7bNFp9XqSXu12oK48GWjQuj3D99uUGn+gblwT
4TP6iZHdHBBZJpd69dtGWcYqJon8+2yb0BkEpDrQNcVLwNSJOk1vJSKKkXVXwtLb
C8uU4/N66ifpMgDLtsPf+eGo7SqdoDn96DorJWJnhbG9NRZMKiQHxPAaX9l3TgWH
9YInixuHht8B6wmxi1CSBGFCtvk8uY/ccjhU7Or1Z1ftEMDm9YUx5WcVWt4YUrbi
KyBpzLHaa0RTD0hQ6kpJqkttN4Jvi4IYIhfMD0PDLTTT8JuWYkEXU86zEXOqLJz4
PORAEgGdn1YBXXQCALApqHdwNj7MeMbbjitBp/bFDSXYgHjb/5Nrt1s+ocSDyIBE
c2CpY5CMhyLYR67pJQXHeJicj0Au4UIuflP+p4EBdoYwTyIBpitX1FvF0MRo/NcZ
XvsK5qZ3Ba333hKayjE6sF/BQ2R8ySMGZyk9BqxreugRJgG31wSMOnEYJ5+cPcQZ
yaA69xVimSXekC/FrbXzJz27+GiPsRHQF6i2TyuS7RmUZKR2fBBdEOPhCzQvWWfR
jeoR3ihGyBg3XSzCqtyxrAOZvMgDASJaeZHdzlaj8CUFA/NKXeEwUPpCdZktv1D8
+QKYtLOndMIORtyzRDQx7DZQjaM39fcJ5C08uSbUiF3Rb8XYNL8PzM9vu89H3vXM
cAitCN79XOIrcRl6BbP0trF2SUEmVtDLFzs3pT4L58+0UbCEC3ij1N42/rYjkgDO
9hqj1kOjRpd+WLB9XlX2xenZABUHbqSFRtqhSrjaazO803jD1MzcY/XmgIC1B91k
cA3IS4S5hf2axOQIVaK1KgnZ2jYGFn/9ng2ImuFBq49bNGVsabB5rXMLkeOrvfg1
ZmLVPnTEAtafohqLTAJQE+ZWXOt7IzYsVtzzxfFRbohNNnYQZAPfLa8YIlDWA8X0
fZ76bOeSmj3wYNHNgxdaYxBuntif35Bq3AdYFLYDnmsdU9gFtrMHVdNCA2HcyyIM
gCI6aswcS7/d1epbln08jw2krv64kJ3Tpeym6oBj45if9w9f+3iCh/B9/tLnBD9V
CnRKw7ab+i3MYXaFJoV0BurmeLvAeFry9vSX26nXeD7s15DIOQJiywLAVPNhXVY/
33rBESNNj2rBvylaY0H2GSXkvDqWW4SefTCpjnjZfMhEHR2oIopUjz6kGSVAuePp
VxtrkxuuOf30eq/zUal6XPYKhp/5ONN/HGJNHYxsGOAlzyNkOrD3OWW1mqK5b5fs
jQUA1k6ziUZUhuLS4cLQxUq0W02sufUJ+dg6NOh9Fg2GMnOLuPkxLSYdIoyYXs9l
R1Y3hOMMB6kqiCNblWl3f/dvzWzZFt/BIN1MBd6ma4mCWJvt30dCv7R+Kpsvj4BL
eMlGfIjCLfLpWt608EzDuc9mwCf8jwk3ItWwZcN9S/VDKyALnh7HAF/ylxJIVRyK
jbDuspsWxTUdotB5J0gXEijUh/BJFdPJR7Mfux4Tof7ysVDGPx4KSc6pIWEmyqbi
8Lxa3kZAGGMpUX/qW4/ffXgz+A/7tfWWgu4ffadEGjHPDmE62lovR+NnoePu+G4j
GmCOhmN9x8jqiXlDsDwSRanNDxInx23xsXf9cfrOv0bMXdjByRemJG+j9EdgGa8m
KkgFI5xqNyW+rSI4GJR66YV06Vp2/szxBen9x1yQk0IPxnttygUe0cP952PoJvlR
Of39jAho9GZdr8EybehRuLvBjYRmVY3LQ+00kz3I9lL+Iaoj6lmAbI5h4A9qw/xp
EJBynWWYz5bqka22BXFYF7/WVpCT3CfX7RVpM44AsE99IR2Iy+WFE04mTdNI44d7
PCuCP+bo6rc7JZxXNs7V34ziPMPRZYPE2U3JQ86knDxb4no849PUloxZ/RYIlIs0
2AdjBUALBDp/ZLwvtu4Gy6Fp6JsIkY56pNiVmR+xknmMuVoLDslN+19qkGEkppLr
YJd4vulP/VIjkKEP2Qwwz8PZAbfyhWIudemvAzDCP97yQiSHcu8GVnZ1CwcJFzLr
IoqDeu6yQJj6KC8ULtQSr7mV5fF1YwnSXFYQsV7Cr2OR0Tb0tDmgtPMiXZDACrlU
KN9M4hqqGK9Y5bOd6F6FcfP5Efcndzl1Qg2L/ddpayFEjA8IYpMbD+YYQTYbJcL4
DOmGF+PzBfz/EGqdxAgJUE4umtdkg03ZJhjc4p3nKIR6PE7qGG4GFXyCptK9eDmF
onLD0kQIB2jadS75DdTs0zq4+bRoIvAeGJYzc+7TJ9UY9iOu1tk8aj/Yq5TEbZ3S
rPDyBF/BDfmZCzy08IM8/kqvA4H20FDbu+mafYYiluFCoZlNxL0MtErkypLlTubP
5SaIdVWj5UZIaMCNHKJVG81ayKWMM0cXTSI1FdC0wg94DTdtf8BHRW8Zerr44iQw
qETT8BB52drXqeH9j4bX7Rnf+60mvr4A+92HCoomi2xRVnKYRx3X6umdHWpxEKsc
upAE8XznTDmAIRkq3yMnJ7c8IKuO01rttw593MlCoN3SZE3/6eDOij4qwpqyUzBW
ToH1dCppdnkUM4kFD+/hEzAQmOTwhBZoZdHA6ES/s7UZJkJpUbsl1aC8afguyvNO
YblI7+CrWh1HfBCpExBjloS/RTBZg2Ou13BzFW689RJgd8G/0yoNr1FCXX/21r92
Yawqi+igi6WER8hPlqD0GODEeCMDl+4sQNLq1EWoC2WCdz3sAmpmJdHnDfemtP99
UQSRAU9LLLvS8GPP9dc/TqNWlVayesd4zcMEZJdVcJHXUH+fnT/x+2f9/tiLFPbD
1a9TvPQQjx3yDllEGhwlAywUt+4Okjc+t3wQvwWPNaHnn56sait0UzmtSIwCORBP
2cMuAIjvtfifYlJrNHUXN0YxLW3zbnK+edZaLUVkw73nyaO3+ld/AdLmhpXHxgrW
WGaFowdyAzMSB3h5Fw90O9AJSWyNQKRdAiTiRwXf4x51kcMD7nJwdOR4oyHnZjoT
lalH5o8NwByoHDNmsIafZtaaybW1+tG/ag8Gf1etv/rwh9pPuD87Y5n/mtfntoIk
gEphhPwoga9yBSh2CK8G//DHQmY1VQgFZKZI7IzWv03KscpcGyQWETV6VIVVEit8
Dw+77xAXGMMC6OGPxb78rvUkhu3tqbRINxjIXXIsdy/l8xHOdxoe1MUjNsuL4x+q
ihT0axNGoLUgH/4M8yx0J7VAkvh9Yttezy2jXHPLMFa9Wwey/Wkt4yKDqq2LXwjh
D3PrHrigeNGhygS/zvZ/6E9vyX0nggW2xQ20i/v+eeoJNj3feqz+XuZa6mGytmZq
O9yjKEa34+pBP2IimA3NbEsvsc6cxLjkZ34ga0SjTFrP1KS1me8vtfD5AeZII7BA
45tjk/dt2QQzxU8ERZvyWefq3FJ6VvBkEjYShdxqfYHXUcyECOV4jCRW8y5Eqah0
sEYXTp29DUsEejxYc1cY/SWrpt5Circ3XP3QzXs3IVyN5Q/jF7l1tsrzPwbRTT12
57RQ4SPjNYvdTE7lQrO4qhd0bXYza1nwGAZ+wtiwHvOnS7DtoRZTIjZRPhwBcrd5
ZL77DYBqTQfDT5LZcIQrN4qvVfyWEvk2ev/2jGkdXmibhvZS3zIOkn9Yp+Xn9UwG
MCcm+8u3Z/Aj49+ONjLkAnEKPJWXyCA2MNaAAPUKiOXLnvhJmO/pDGjNakRW0maJ
UP239RrLSeVWrexBUfCRuxv8uuD8xhZm9Pgoii+zWnVQbl/GT+5urLmwzbF/RXpq
hzFTmtuXuPtA9u7DpOB1dVSfH+3B1sVf38q0dABuALA/v0V61+rpSJ7SVvcT7j6I
JkHerq9MJqLUdLGHenc4oXltPBWGD4a+OV08i+cbRfHw7kRccrqqyJL4n8aaJwNX
1j/LHAjFm0A7PSpxnH0jWDtgQVdQw5IEKr8q2srQFcIpCp6N6K3Ybv5jSZymkmJO
8ivrYCKrQHohuSyY2BsWroP05u5KgJWa41xlAVDvc9WPD5+YJv7pwibI++V9sg0p
QDGpOjnJKo68f8xwKLQ+Y0a1K55INZiiPjyacbcY+pPTUaXtJK7oPtsnBzdkJcM4
sGtXhzMPw7zTe/pMrP7GDpxdmd6BEkM/VmKhWYpxXL30OragKyvuypOFC1zueV2b
hTR5alBWyADS3wgptGYo2YIYWUpuT8vUubdeSJfUaKBgMJ5cqUB8BxPsIj2ek2NF
YJt95D32Y/Sf09JVIhIY45/+z7y0PB5ndxt7DKgKbFIfYuxHniePT9B6EbjNEIi+
uw2uCxsVHI64Y98X2KT7ep/gY08U+YtvlNUN0n1X2bzjXTHNlIlraNBmN1z0BOhq
vYOyxtuJnE8xmQdq+Ro5EOJg2HAhM2GniqRQEVGhJsxqb1EXwSpSWQ80VnOI55An
qT/MFeYb1SS7VafQZxXzO53B1oq+7E8ED0dBXwyR6r6cvSfDBbVzK27PXXjvDqG3
in2x0KzRtQoInjRbeah49YsSgJaI6vUmFWe3OC1ZjVlWdZ74mrdFFDM/RvIwp0J9
q5Av+qDlCoeP2cWlGDdd6nGFHrVRMrJxg+2dMVhuXVyii6Pn87wjBPXQ3g8UpWuO
XOde/CMZl2eZ7zPNpy4Gy248Y7cHOT4z3cEJ2EKQgSVgVwYIsKvBbmH3VEWA31BU
yHiRko9kl9ZSR9TgyK+hJsR8xACt1dzJAVmW5cmbJFpwP1dV8nyMKYzmuDgEIZ8j
KtsgEXO87v09yZfLQz5jkbZAZ5cHafA52VDgWwGvQJ4yecacunIjMDQoTs0f/NU7
QU8eMitmmEwd7BJa++3gbhmeYMT8d2FA4vMamZ9t4LtS9osdHoInsZr3ME7CaBvB
jH5+Ovbxr5E4u+CEX/OlOcxQjAMFoD8OTCwDwMF1qjwo929DpdVXsF6RDR4GPkY/
L1kbbCy0Z/HzoDfy1kNVIIdcT2F6BTzy4gGg7F/AxaJx/bEOTawlrkgYv2WUrP4m
NbK79vMBApMMVfdaaUzMFDrUYW6VG9h1vLcQmQNfZOyp/lwS3MRDUnsRtgbYjoWP
E7iZtE/5UX2Rpp6Kxf4AQkKiF9olB4jCXpruX14Z34pzv8hi84AwL/K+WQySBct2
AT+DRdAnG2/rrAc6v7+Wrqqhu+KrTZ4NWb6V8n6I4HBf6JSdcbeE6sPQ68LQ1F0O
NajO2hK0uQKolo5Xe2VsGKajioLQuxYBPyxEjQ+Bu6MIUdZuKRH1qg1IWzG0WA3u
ullsWlvyy7DWrf5kv0vJxM2W4T+lx2ndMIHYp7SX+QmNkl1vTSjROSmyeaZtf5m2
+7fCDswGfBZLhSkb93bYxRlIdX+wrUu8UDdXooiTELpXKyUeXu+5RjYpkwK3uCw/
V4iBV1F4YVyd18DJOkzNBfebj7ljtTfV+fgD7g8CS6xmQf7bjW6p9xxHSu+Pf+dr
2T5Im8D2za+dAiX9g5P34qcd2eCmNl3Yyj97G5SU1f7nUg3vy3HAaQYOsA2lipBV
IRPcRh8pX3V+agPMdmXAI4uPg/4FuXGAHUOCefsWbObpYULX0zI64jSsGroj+fOp
5SFp+htviKAwir7M95CWxrgbjskP34zxq8+7/csvElRjRmxib/1UmRe6s6363R8m
/BaUzgGrtT9eipOC/0bh50UqZN4GhuLehrmEGhaeC0KT8R1bxn+7urmfeHOpAhpS
N4ZO4WJV+8Phl79ZhAJ61OdgLhxq2iHDs+LvVAUEh8d8cbS/BHkavatvP0HxASQk
WL7jDtq+p/Hskmhsl/ga2uBmwBl0nkppJFIz4QJPRadxZvjN+5E/tdt7Ml8wT63V
yYAYV+Fyk3Wk2QXBOIVPykfW/OhBDyddWrVyoFZ9N1lkR1iAKtv8cOm2TdDHXoy5
sLuqJWYrnPIx9MhNQNwVnGO0T8z2f3YdKxDXbbQFf4Q76uqEYtzGPyCLMovzBQxC
9XtX3vbVDKyhNF5dibdvZgRW3T8iPhSX+hwS6XZ0X5MH5kGUeopCky5D2x/Invkk
UC+rG29RBFuwlMv+XV5/l74o1qoDlUwWuycydLnr43ahxQOTr5LljqyH58Td4XYG
7aAMwiWbosMPiv5oye5W7GWInZ6kY/1lDl3F3LOLWhSDWn+9WkWQ/GaBsvB+HnZS
i0M6WNbZpMjiTWghbEBfgUkFPLpfcWqCZUVsOy5DYwVEnoW29P4NaWaHygDucJfC
mfv6Cs9OhD39Mu4YnMitJYNWNMrEObqrv5/wCQ8AVu/qX/z0wmH3avWrXwwAuhJJ
9Dfh7Es5hb4sGlYTpDpFGtsAcqyck1HbhhIW3Zz4Y+QuK7wd8Ju1EPwodujnBsc1
jLnctV88hmtmCIpF7IkE7DokOBc5xN6iR+ZkB3xkMuCZ+rzJjbtaiV6vyPBjmr/o
JXPIHA736uJOQE9dYehVetBFIyaLCqSbhLo2qi6IJ4SRdR6v8M7ufoHaqDRzzT+q
qTSzZllhkW0rC68x36un0ijKok/DxD6uNM4uuSlgGf7BUVWJVOeKm2BJn/29uxEW
wn1/MEeU7XlU2pKpnVq7NnVVUbjbYuWUGJ/wkA4mOC1ta/KHabrfMbBzFZEyML6r
POwiwL1f1aken/xlycCt/lUbAEdvsTncOZJ6JZbl4q+AKJSlu4iieiqOInohtWqV
M0ngdpdEzDh5jGqLpZEfGpiwFPi3Ry6gxXFPyb7tbaKGUz3NkDye5pu6qBf3fP0I
uNRYpTa9PG5E8o5SLRMeVU7w8HYELcAIRu+KypW+o6OSx97gbBvDnDbIEHJEyyPh
KsJuhVCVwxQP8kTdFAzXUbmyWkOAqzpzVoE1jGeQCMLoFDtCw3wQO2PtbPntvPSh
XE5iPSe6tAZpy6y3sFrcGdIUSwdEysLz/6q++Y+IW0g+GW8Hs9U4JoPYD1x0Z1xH
jPijMRaI8Cx8MhrqQ7uuf+iHq2maTS7e6uSJwITKcbvzK2v/8nWoUWXKRn7NHRw0
0qs8J7Yv6CI2Fb6kuknL1PQGl1bd8gjLhJZsqBQR2nc9Pz3Gkspz2qK5ytba2yo+
dVlIPUsTo0F7bBGI4KOQum6jraHAlWMagtqxJrkFKc4heAzAb+PLugAZXSHZNHrL
5VgQrUp7yKb0dDakxXuav+SfEvFptpzAlFb2DaSlW+rzOz5sV7vWSNLLv1lyf547
TLp8Vu4EDtr1/2L7/7S7AYW0bav0gS6bVp2yqYsgmVHulJ/++F0V1mqr1C3YNypF
wHgNRN/fRZjsrLrqBpGmStOr2PQjFKOreGiJC9tXIZIfuChYXyBnsp5lszoUBDq3
jGssSrYNLa/TuZ0dv/cHLLE2k9d7JykwfnUq0zSnM/+DXAgoayFUbCSAUrS2cMR3
y8SlaVuYTVuwEvf8rVofD5aZvz5h+3uWL70eaSicd+tOj0bUjH/oLdMuDQRdJGiJ
+oFANAvnhbgKBbYBXOt/pUNlwNnPt/8En1mkwYwQX9Pkg1riv/E6qW9DuQ3eXrgV
O8ZspJXU17ItTMcvps42+ws7DcNoxDTzHamHJXos22R9E3BOAy/W5sy+bIMNucFa
0AFLwKDOHwDnUSYY1OhNn6M1JLho3gEafoIqv8qUIXPs35U3twd+BEdnOM39Y5p4
LfyrNvdErG1I35BHSnpa2KnlfDeLhyjUZAF984srO5lesmwjyoyuf5cusqdk4uzB
X2HxoFA5NXu9d7eywpfdvR+5LQdLkXyE+cM5qL4I81HRpPZYkJlZ6GKLWejdXHLZ
IkkZ/weKOJ6epupwqjhkiEU77gshrWoaco6tZACQpbiZI9fAhOe6evuaVn9e3Hne
x2Kly6wk00b+iBU0ZEKE+qzxvNIaVO5HDxZ1atvmzMqEJinvYRfGOV9c74V5L80X
GgOYidtx4TelA/DLQ3LAw7QvY+5OoHCMl6cB4sxDitMMXgsKWnUqLo0YuSjWM5yT
bP9I3jYR/b5xZFbP+YzN7gHRwrDXvp3iHWM1PP/ytYnbvuACBGrX8ZbxSVSiLiLq
oo9XjXwTldlCSskAmC7QFuVt3Q349PIAhsXVJit2bINeQwD05MOWsoYab1GCjFGU
jwIp8132y5EjJyYHwggRCXlNKA3y+W2oZzhZ85L/YsEX/L7UuVB+JG0GXfZJEis5
Qz6Sm7jGfqq60XFyq/RPcWS4tTpanmWAbdI9myyiJo46Ar7HTGmgDStJBmoO53a4
AY7R/IVyIfw2W1wMFX3NW1mZ8H5UtoHlewHnNAa29Q3REmaMxpS3YjO7HAZc2F82
CaTXKvaYYGE7zhjmrUjTPW0zyolA3HyXXKsC5+jsgagc/KDo50270LD6aU0lMv91
v7zjWCTcQhgVJj0ojNWveFb9DY7nPFI62wqOcdNVj16mya/7QqlfMzV0pr/l9dfZ
CWgA8ObbPlLnD4yX6mteHCRdPxF5nW8Oo7+bv+hWiMUi5uQON3lcrxzpiJ/jaEXT
AfpWvkdFMBfQi1L0bOj0OhgIuAHAbMTFeRuf4m31fyvE2XAWd8YPK37joGHrQPMI
ES7AvedVUi96iEXhyG0zZB07OsHEPK7uAe2BJgdjq27WAnoaGMRUQGGkhXPL6GPq
obCj895KXwKGB0pYBOSJJJmoHtkmtVhI8xlzEOl+3mKdBpcbY3otA+Ww8I6SEXfH
darxuhCkPCAJVuaUqMfPboZjr0Jhttpe4t5Jo9kVcZQNK+AJM+7M9edsjQwi2ZYk
zx3CKej9pe9oOUJtaecl0PF786J1uCpJpgkkNYvLGvF+mKtQz+xT1x29VHSoOMpa
vikztG5eFAZXs9LgZwNbpp0N82gx5yoagf32qheCtgogoYJByM2yC+WEp5AmzmZm
63Ya0Ek2cb72WinY3CRjeAK6sOmUyzqgetm2BIcjQFZP74p7cf1cTVo9o/i8pnI3
/+g8EFJnNXlToRi1voDTVx/CbMZRfhuak0BDd2UtDil//c4eq/L3hU6mI/psNn/g
kwGT7V0nsKHJryp8+ug94p9ajOX/hY++aYJqsW0b6wlkpLYRwR4HoUfns/szDWQa
ccAIPYT0aZHPXtnb/c1L2LQlFZXR5S+sJ12Mzy3nr3dCS8BwWCWZeHpMWtIl29Ra
GLFg1BWtPwSPsfTYlxWqL3Py7z5vKbEo77qberEJ1Ce1LA4wm3d7zD/EC6SvGBeu
5dEM2xZmKB1HKjuoKZcLYwT7tC0LZe79UO/XtH4+LnRdFUrHsM5iDS9RsMeA9Qii
VYLFm/jm9ZrTVFp1l3nPw2BM9zVp+0VPMa/BN0YRZypAXQ4vTeonETOKpTyusJKr
wG2IU/EGSd01mrWi6Ev9lcZ35Y0xkSPU/xg6XpDbdOQzjeiFS0EVEZvXbhTHunwX
x5o+s2o4/dI1m7uQ9++ks5oNgSqlNhPep8z2XCaQcScDCCx4WvxNvnCh/S9zJLs1
nvIehIPJENbcQOA1RADZ23eTrXkCYu/wFChFuEd/IUxR6PH+G49Kon0aWqg+OGwn
AB5cJ6m7BHbLJBc1Qos7A8VdjDnmioLfL7mMosnPv9bQSbO4fhSb6gNXZbDjz5Bg
tJmWXfbUs0Cu2jTGPorb26ChDgSTdyKjjK8MYP75B3sWLfOGd+RxbG0b5hAbKH7N
2uWkX/anBWXpeLb/SFzN0/3yq1rLIpOWakojwFBqrmefQeOoUrND84GrwyhMvwI9
3SFX5kkBDTPJzl3379sx4DQpmde6R/gfQ40WnTOPCp4c7QMsvMzCW220omU2DDsG
eQXikb3VDm8A5vi3gixvX5za1s9eNJrUaiUptEIo28huJ/xwtYrFyu27UKkiTIcd
w5/p7m0uaF7XbcWdFZjBX/N72cSL3yaCAc1WdKmt/cWXsN+OMuneQrQYjPibp+62
xQkyiOlBAcsulCzJNQkG4dZOD+wxAAfda34YNlOvVscw4h0H9L/oSTFo5G9hCElG
Mjweldpvc1fCkqP1uKw6bWmDo1OSsj4PoLZSevGf0Xjc0GWQ6CXcsxfMQihg5MvP
/41TUgk5FesFD5T0es5QZ+K8Unm2GvqCAlmvRoIQaIDg4eISOzFXWJL1sir3f8b/
vEs9DwZdnJ4SbH12DbaOVBpb1sE0L+nYRoK2SlO8q8eW9HzJfYD8tzFKJkwijeUF
sQ+YwA4/1vGqXwzU7p0eIPhEBIKK6wiewstLavUmDRkIxMhSbJGHZyE24kd4zQGq
uwCUOpYI6+Yt65DRPVxsd9s/RW8ylwgcLG+dM3SzGambaH2ol3I/SCa1lPZWlwpD
TDdbSprA1f0z1quZ3rfVEBFlKIBh967+1Jxt/aidGLtGnoTpsXMNoJSIxs/vtyuM
BPvM55ZbpVc3h5bPfp5+vzIMpIeeE1ZjlOK9s0/gEwhN0/We28GYILMPS2MlsJzK
5x8ge9IQ9yd5T2BY6fwYBOhtoZ71OgjsbVezm1a04hpjmgKlhFVD6FA1Vf+J2aCs
Pvb7FEJ0Y773Ucw48MVc/RUN5KV1a4noAR2+7xFZKzjhsXm0A23xjO+TmIEWtWsp
jcx4DjQNtYCbYfCvV03PA/uRlmr1kGyab/rrqNy8ypvqw54VTVQYjvMPVIpezqAX
dGFFFkQX/ItIpHxBqIqFok1G27NXZHkrE9Cp+CcDgPuXmgWKWFBmOY1l54dRLbcq
aEfNFPiBjRH4zwKwq5/QDginsm7Ylc3zjq0cXRmXQNlOJwDAjbFy5DMPH/uxCV7v
SobtTUq2PAU5y1etfkLNrzd9Xa/tOF+RMvyDs9pVMfOQmY/tLoOCXD8DDjg5vyTB
qDVshMCrKCbNw4wOdMiWkh9XYxAOj/q2okEZDureGiRR7myaboys/ZaduLaBZDNT
XwVqZ6gVPWRLb2PBK+Z/qjWOs5Fu55yYnskFpnemWP+/QJrNzlSkeHpzyPlmulHX
E3cRGQ1nkJshSQw5eKzqkief+cZYqEa6fgZ6Y47+xZkkNN0eGcm8x1sqBMuK4XOw
iA3BlC23t40Gxn66yq2+qKBtzr7EVMhqkL7Hqhw/aOiPVt8Fxo5qJa9Zz/iU7/JF
X1lh0SRf7ukX7I3AiVUEZ9bTO24/L6Fu8zCuNiFngPfTK9bc+tG2Y/3o173aaUs3
CPAZPLXCTi/anVau9LW5d9hmEnUzl2sxqlBK6zjeTS9AlDNEKcKYXFKuXxHRhWvv
XXr2pmz+ldbdFJ8UGpOdQ0l+aL/rb6MV5O379TiSBDDYLuronZaSyUlg4uetP8FI
3UTdGOQ11cQhJP3E/bWTgjTReFXDdMA8vkUjxvxxDrA/Lxxfvu0RGLqtqtpVFNLD
ZTakqnZ0JyRh54Sfz5XrKpzbCShKZvhLEL37c0afQQOE0xBskfZOVwCxmTLmZ2HB
fQEm+dNISckYaQ1Tf/GPDg4brhpfOjvOeA8HwPhfIJa/lw4/Mi9XjKlUMWR5QyWN
afcf7Bb8c810iPStvBpmtvfcwz3LDuMBrmF2h0NHwBj2kszLhhPmwdD5Mrewi6GN
4SrDjpubNI/AAFrTgde9KIap8y4l54UcPaXmzSbHWoysliumkrKquzNbixIu9XqQ
2J06A9FdWOnslbi+CGejYmi1g36V9WIsg2eH5hMFohW3GlWtkAylBEV5/qlIROQS
1FbNI5XlCFdkKRElzCWPogUXsW3diRSHau4Cd00L68ycED1e5ySzqt/sYJE7f4jb
5Fb72Rw/gJICutOnutVNPB3btp10ugC6HCTQECcAGTFT4NETSKBk6y9VDhfWuxt9
0LOk77UIbUPMbbCf4bpYvsoOlkjpBZm45hRWYGMyzX9d5gIbgTbeqfOj/Kg3mZyI
CSZgSzSfBSuAHrl8Hd/Q/LDntG5g466YmPobfifY1+jf5ngaEP2HkU+1RUBI3E1T
dYRAy4nij0U0fwr+PmCTqoIkvRaWEayp3Wa1nO9k6fOk005debildmtWb3sETvSH
2Py9OQq9gT7blA+DgnVWUP3nKi3VTQZJgSkePcDOUFIOypBzQ4KFGTg+oUeAo5o/
KotqyZORK86ylR5wmS+7yAZC7vCK7C+hs5eLROu4Zkr++g9lMw1hvTDvXFdFkIfR
wakhjMhZEF3ian8WrGdwO7OybRFlnEQZ/ikWZ2oed3inv9iz6otYD6VgxchB1KPr
yFtAKdwEgG10gekDOaJBkeRyUeEmLoZGQ3c0Q0YtOAtzLN6VoI31JXtLehirnlHT
1oXg4fmZoHaUsPzS594ntifVQ0Yj6vWEg2weMywu9mSWMQyckB59RYqg5K0d+JEm
keOjJdT0bSqj6pM4FNsTGcmUHSw5HZVMADqQh2Pg2Jxc+jk/oVtwECJ4G1x8j7nm
jqbU9tA6xHTDFFlo0OTR7SCmdOcb3hLOrMpa+LsTEkvs6ll5DX23SJcrCNoMQeTu
HNQvTH1VFEuoS6NdeA41yzPYMYYt/E6WmU9mApVS+NWC2PIdA+pj9DrjdlCU+VHm
QDGAwnR7YjWvFLt8PqDz36JU/Z4qxz3Y88F4Zlk19Xo1LkEimRCG0+S6l4olAB7d
aulo2q85ePuIaaKeVMnbYYroyyQxVt5s/RO1tsuZbohsG2h2xu9lsH4CTo7/XaBN
7mv1s2/5x1zCFckkrfl4TYOhIuoaZrOcE2q5Va1k8qmzDdY9TYXdKTjDPo45gTMY
+hMTp8mkA7yFHBKNrjV71zRI1M9SuDNZU6TGwRLQ5PJI04044N+xujZ53DX+FOG0
KvCKDds0pg1t5A7+iAryMCInZe2tWcfbBIhjqKtBJOYRj+LY2q6O1/NuPPnhOV1i
oMR9/+Vz+94QmlqS7nIENUlYA/a4D5K4Ypg0QHhDQHj5N2zVA13ykR+w1mLf6Ic4
n7u+Yb6O5qeJ1J+CfkcL+B0blp2ELJBN6wFSzS33iyELEe0YEaZ1/ZzQiNC5ouU1
8OxGxNY1MXfjp78kxZf5YlnxBLXfHZbMjYB/Ig2AktbWiSPRIMkw7b+96/JWBPd5
bS2J/eJwcOCiMPx0FCZ8piXkdl8f9APDjTdCyBfbDxWZ7+olnwUSKvg9PjJCjLae
HN5gc6M15v8yg8bDIzxwh1cf1Zd8Qq/TZCwnoH5nhJa3Qb/NCMwUoCbqupj0HOz3
py1F3S2SdUi0mi+G5B36JDypWD3UUCSu/+RKc/hkBiN7jJxLvw5nYizakkD6aWQq
KLDu4lbnLJX5xDL3ShYqKu9UwQ/3gmCl+M+NdqnZ25hLcKBAg5YoMy8ZrXG5SGqG
ouSQVsQsr8cUKL2NLq9YTWw9J1kN14gkRSaAF5VrIxkgaCaXzMfIIb1HZLvnZja/
QVexm1PaZnDXUHxqCuDIuBvolsfb1mhqEFAo/rqUu3ezxeD/9qXJIAaWbrII6Iis
NVE/FU+HHIsXEoZ6MvRp4KdnnREANykDvndJUXmolqL3Fbj5tUIyzilYiYzXCd/G
v8CANFjASVSFQXe25SngHpvEuZVo+ORuTJzpKsiuTBwwBXepNrGnKoZeVLPkTMOl
IV6GIJXnuxr5WiJICYEKSbheRileCSXN14RO/AlF00RWMtL3YQiMAr6yna2LVjfX
0jncGeend1JPvcrVDGGGJj5HY224TW46xdjIqxU8OoVw2dklw+lFsetO1rw3sZbZ
YWWyr0hiGTLA2jYwFL+qHF+kAX4+1Td0ZVEuT4JoOG3NTXQXOGC7ojBBh1xlUB2C
QfS58kOyLIkwn7jqtZ5wcL8O4BDl8SDyHTgGgNz2tJstmYvPFXBb2Dip2FTj0cn4
GKKmvNQ4sO0wGX6odJ0LRnHOJ1l+i9ai0VN6Dd0kGRIQv8epve8XZDx6kUps81GS
2kh7gGXgl0tQ/V89uH0B1kEGHh7NV5lh9ys0NgEizkDfLC6DoheDkFWf7FuZdWNf
li007QDKITfGiabXa4SzV3T2iNHQiqvd+RHbX3E+DXSQABdbnJnsGBl8I5eLJ0Kq
CDhojX8eCR4xOtOc8YqiUmbDA0ZcATN1t8sg/Y82RfZ9DrWy4eZQgeAt+EQ+qBcL
UKG4sUID2nelOu44+v2UfE+WpC3IFZjA2EGCVdRMUa8+G9+KMIhveX9JH31jXQql
uburUJ1Bvya+rwTYstZ/MVofPm0cDQiGljeBXJbm9shaTUawrSbMKY9TE639TlZ3
qBCBswOZWNGjjn5KuxYN162QuzutXhyOGGFFBvCBBbLfjyeeOklTJOkb8q+PBZj4
Ujxf231AL9sy2/mLYf0qKKaWnx8VsLb96p3LhoRfttG6JsleCRBlwQr2LvASMdV7
NHcH0LIMwYM5ZR/Oxi1uuqHiaDfiiPThULbBP3g21Ym40/VIlb1BlmGoC2DXTIGf
uQmFelRYbXeSxVov8zBI7odZGMOHw5rNslrcv0xdh7sQTryeUZ/pK5hFfJ3SF1H9
6TKCqQdYOhxwf3Gd6sE8STMGcSuXTDPAGs5xoL3Fd3ybkm1knQO43pGjC3lvnmGD
dDH1RsxWtCf5Fq4B08JsxigmKgDdsiYdDnMopctIK0XPLefZzBXyYV5FuLHM5kEX
q50SxUsAVp4KFuNDsePe8kTTXPeLAqxcm9kdRWCVcztnNXgTNwisxhIxMj3qc9H4
e8zGFVIUZVqsVwevMysl0khI/MHwg8AJKawaDv9302Q6wEgtX76qwrrdi7R+MNSf
IiMN9yLVKYOiWJCEJePGq/NGfaTMpNuJ6C4hfUMm1PheIqvEU04XeaweqTOg0yEA
bTjCQ5h3tYu4NjTpPXqPTA4gfOXeUWGwwk68JyViRtRzF2dT90FyV+T3fbJ1bSMD
8HucTK6l2SKyrOArQZpOMpkrQi/fM8IGRjFkV45c8slA6DKxkEGE+jso4tR0l1tf
gt3Wrkz0HS6RuRFeWecpavq+HEG1SXlJqRTx+IuZ1mOEIu9petbtw5h5LSfqmJcl
lpvLU8hbHU9ZJ+vej7tAZnK0sc2CRAnS2AuatSN8SmlNZNTZ9J+yycAQ/sCe3NBz
nj0pzfsc2GOiYV2DKOi+OCfrBAh6M0mVRazT6uz9wZXztC9AVFNjvb0oPmA5D9iT
DRZhQqaYCW6+e3bXXdz2sF73AJejf2to0eglboHMHml6Nk1n7ZCxbmtAhEODWYjs
2PDtNngHLcZeFB0UWQnLs9+IsKQnQ6GjIQrvxmC1mEXQcoubNCMcakSe5N2LVux5
+Nk5Cq4/H4t5G5Bzwr9Eem66fDLLvLOsEGceQhwMUb4zuSo5bYn4G54dMqkVoJTS
vq4+rAv/agqvGWmxe+F820db398xFWnqulcrCOenVO9l78VbJwGnB8F2DM6obh4p
jun5E4OjwxZUUEdkbIy/6KQ3P6PDhi4I2F1xML5Y2CYR7cQy6I2LgWpDsDyjTd4c
gn2q2Yqv7UjGI+wJnTZHKa57W+Rgv/ofi087q8UixXEFr028nq9XTy3aMApULAGy
U7BXj0aFgPI1+URkQMo3csSOIgFGKF2X8ijIzBgu3Jl3TLN806pQ1+Y+jLGP6fXQ
CsNSOdJF5NfuIxFv2LVGY5o+7ysDfE6jAt3jkj9Coo/rLKOvXZfbmo+5WD3GyCGx
BwDae8xrDL0T/IpQ2mi9xNmBjXkZrbqUTepdoyV9P2Q/hvwX4/7micRcQIv7Y6I7
WyZfqr7ASWglXOs3UERXocyOgt4tPPkc/lXd7cWrMmlnsdU4/7O0/Cb0gIc2YE8g
dPBV3zXm4gyOje5kCQlxtRPj8BaPT3Qn2VIixCqdl4h1aZXDfgmVCDxhfxUxew2+
drrwigmK7KAoof+lrq/cAATUV18BsX9kwFQ0l5NNXwYx5EKCBYX8Nd+O+jEd3fMu
bTwf5NXy3ypD7RNFd3RTIc63XllKShfE0cJ1H0GTltPmigaGyB/XMoog9KFPtIVL
4QUBGq9+bB4Ip7fI2O0cazQ/uLRVcdnuMREmyV15mx/p2ZlVifYk+Pbwtg3ePn8b
WnmaaRl1mwRIsMjGtu6Z2gjECCoZmBJTXS/mUzav9ItjwrsduHWFsu+FbTCdXiq6
SRbGHtE0X2Q/WszhETCjIqPdAIyoUpKWTdFSgFyQ1aMkub/W5jT733GOQq09Y5e9
0lNsvor6hLLB/jpvI+chWq4F1IFwwmJxVvOa4osdiibCCwL1fOe3jt6SSUWTGcBo
+9oZmWrzi/wrMz9AEBR+ZQ8VZvaM/Hnyv/SPqczS7GOSemvk1kNcPe84DaJrqp3D
GomiWL6ZJAe7JZuDiBQQ/kE/7qm4hMPsol7oYC8gSzAmj0BXWw/xafUMhWTCEep3
qVsS2HMmjV32Lt5v+0/SyN2md1FYfqdYEkDFauc3KgSeALCL/7rkzvgPgCtYxJne
PlymjBWLS+C4aPozHvB/znNkNSh21EdFO0cNCbHxljFjBq4nczIGEG2WK/CRkqkC
7KnB/c5IBg3gpBCUEz7Jsnm0kSrxZZfye7Uhv0iBUf5dYcKjCOV90YcgIG6O5ghA
1OOx3HUv2rApET+uPx30kjNXRTWpfkOpG1uYBWDISsPcfzs5K+w1zD33Hls0L2nm
5g4x4+F4kwou1ZBLHHBjwaXNLzTO6+UnHnXUDhGE//jdDi83GmQrwBBRgRRPSujV
umUnh3MCE1Z0YUEIeu8QxIDyNYncX7h25apvHknFRCBi6PwxOsPjhUmaBIgmlEWV
UnM8QPZ1MpklqMFOhn32LeWjDBPE7XNcfeQz948kNHqHgUAHQnc7+WsCGKaYwSC1
jn8q14XyL+M5qghtJhW86Ai5ziLAWuHNG2qthWQH66M77wwx9KWml1/hwyu+A0Pk
xwG129WhKKa1cVYoB9IIFMrY0SNnDamy2vp4TeXW89PkZGh6/G7St+K2mmf5j/ma
RzXn9Gg/68yUGM3TnQn7ZW3o69vf/A/S3Mw/xESYhu1N1LwMitbIP/91ZxkKbGwS
bNjxxMjyKV12rX6O90tvtm+PLu9LJLNQA+vYMOHq602DiKGMQLN1HGIY15u0OkaV
0N3dUaI/KbGQqlAfJkxNHlg5pLNtb2Nv79SbjNl7O4lAymc/jEMCMScR2GFZxxjH
d4JSeIk6G09Is84sLTMtVYJbi4fy8s8KNQzLnN1qQ6oO3537f5rBccsrqS2RplG6
UtaDRM1I6Z533XCCtWv0PtSpke2W2+oTSPBli4bhDZJ/vxhXu2HemPsJutqkheTq
7uhSb3EMWpto1+5+m2HSvyS/tK9dJjPW0PezRJEpeC7jRAtj9IEdJ8pWcrm/zgXs
P5VojaVb4ZgvccZASmuJOUI9KTavZqW0j2eU+Yd/BzyISRwrOUxIFzSMS89E/CWQ
bvG8c/bnaLJqp/ccNrOZIti17LZNtSV1bKb10KrCbJRU04t2ek1leUvHlvXM0Cea
BKCWHBJg4/tBxR0lQDzG5ZJCcnf52hqnK8QutKFQzC70nY5Hl18hmz/0pCsC974r
2UYCdnkhayFMrHLkMewtWDfuhgL98SSs4AgdK1jDSEQqRXCsCgSQ5pUs5YYF0jRp
OmmJeQlUNtAZLxrWLF2qvUESuaFsa4xfc0RF6khvc1djxwsfN6hvf737z4rNTeOG
Fw+rwjWTs27o4cQinqARQ/yxA/tvC4z/d8IdR6Xpz/GE/c8AWyHxvijEG7s3CCcY
gHRpk7zotOm7ebogGXI3U9AeEfYPegbe/wvlfBCrtfs23rSMhh1E/eAHn8sbHBU/
7FMNSczS9yinyrPN/dNJ/QkhOWblQIR9IgY0U5DHCG3uZ6qF+/3U8aqc+F5cV+0T
BOmr+FDor+7w9dVHha3OhFPd2pfxnWvBSpXRUCIrfO82f8K90bqBKC0LyboX2/tt
GJRo7WZO2mzajG/cITABh/G27rbKaAy1SyNshbSOKZyfbpvCK26rGEkabetwKmp2
EzDVyiIQjUFSLLNw2s6Nmdpd6n6cO+uoUFhpQxFI8jnXhz+XQqoB6co2O0ezuIpN
+1UTXLZ3KYZYgLwYJCACip8Hv2hjRYHyhdpv7XTq2XzWLBo9lR8p31RZ9E/X/H/1
9qAFGz6Xl+ew4TvwsKcl7QzAfRPQbQTwnqM9GS6B0Foo5ocnzpVsvEGMcq6aKJ6H
19RXbDVjYKZ1Jsoh8uH2HnzVXzd5N/Qa3tPiFLvRo+APSFv//KDhYu2zT+cP6YXY
XAMB1EVcznl70T/T5+ZRUSTSvzAP+Q3T8hyLCR1NNsftd/DNqoM2m1jg7ZINRZ17
QN0qWVVWT+jOh4AYMoohsYb1uc9bLFPAEPO0uDx1GDgFw1DkJ2CsYTLos5dcHIBz
nhODfVUjhOAPGj3p5L6xlWRFbWQq0gtvogVS1K6R6d/3vE7nAwLa2NzQ6RTM7svv
AHflxVvYOCGF7PaF/D1/GO52/oVoxBRUIiJigA7OX3eIZ/tpdH0dPB8fQnDzHyEw
xOEiNc88x6uhWio3yFa1zJVtapziti5qLFIDZU9xaGcRVV6SnwIX4wJ3Q8gsTPFw
NETSrWONP3jga7h1FchR8ydTeTIYpFTlLYMLofsdV8qGZoi8WOoFkDMmKf4aTPHi
b/DdjudiakGPWvpAn4HR0KtiLj3wYWBpnkLMj7HD5yvjuEvzxU1vBJwSd5PnQGWH
nsWwTmDP87uR9AB41XbhcjmxT+XyXHaI8fkpelWR7d0S3SCtcVkugnrUwhU+YBDi
RCURt12gYZAz0Ernmh6oRlIX1zSO8JxtTKZJnTXppk0JPYY71NJ9R5UmyueC1xTt
SBTJ+rRKNIz6Dr/ylJ5Gtl9yO6TaN2RPtBDafAuCjUXuO4SzPc+qXGxtLwr3ZaAb
6xUlsT1Fw3p4/dp31PMk920DMt2SFBxZV36EbuLEx8ipi6ej2jRJXszs8Iyt71eG
VR6XViS3JD+uFNgqQyehGTnUowxhjLOtlSxttUrFXdAZAFnme+3nqZeYGL8R3WSs
J5hXeH3s0qwe3zvuyvcqKvK3w1Yee6/8Hct0AHfQzEvxCM1lUPaozeouL6y1HmZG
ZPX2NY6/rk1s3nclXebktInV/NFcyiYjSbbja/5cHZKA2O98y7ZwPiIlJBBRYxT8
3lJeMqQEw1ZE0KUs1SinUbgUNZoawKe9TzaufVZJoJRZCqQi+tl4LWMAcX+Z/LRW
hzdxUbktPoAvr5CJvzF7RTscHbNzTCgfrWV8Ltjy9+i2MgeGNTKR8rBAvI8Rlkya
ugWy7yFkhkFw28ZKAraJg2ba5XG2RyMWBYZPQJgh/hoV9uN5ZjYN7IB5+q2JLMDL
NyYDQaBZfeSqovOImoPBCy0uefbpi7fBSCRTRClmI6m408AXCmUoOlRkeyYdJCPN
Z4WBBGNVkOOGtskQ15A7B51gMkUZFNAveHIiXE3Fn4BYoTQO3lvqd0mPJbHvRmdg
qggGWJAd93hlnI2+s3jBj7Tj7uQBlPKBe352L9JmO6ufR1TPV2JBooB3Rpqdms3J
SrjJdBMv855KbYMJuaUMI+XhGqc/XTIZeYgw020ySJ5lJ1YrhEKmAovcr7zhMeEv
OAkvG5bjwM+WVE2OLvp42ATnsZunxiDHvywyVRtKjM3i+iwPlesmFHR0+cpKAm1s
oWD8kdA9RKkmopkRPHm7xj9lY6xvUFP9y9HkGGiI3vGk3nFe4hjIUc806o75N39h
Yts77uqW7N5Unj9OykWKTVXO04hpg4KGZORaML0/Rm0GMRuuBcjuuStKYDJXRmVl
oeekdH7oVQ6Ri/PfrbcgvUM4UyXgf8A0EQKuZu3PCX86v01jt9V+QgVJSQjYKIGh
5miXh2SHFeW5eZfuTBpwwGeo+q6nu7yjQ0EwYUsQczovNv9948QbkTse8PkI0MSC
EDfS8mlfDz5FhYRAkmIYn8Jf+S4gQjYPHWCyWVwEBeV6yfjQpLXZG1Dlrbr1+Irf
/EITj2vmDZ/XKKt9chTHkSeHUd109rCdc82QKQwtXIgux/0oCjhxOXX5OwRwHPxA
JkyEYhdjj1uEt8CIwjUomHjQWWu/tOHJK7W6l/xS+JeKu0YL7mjm9YJ+ktcx4uPP
FdXUhEPkiqxEbW5ifiXfSK4oKCZm6AGAfB/qUKLkj2CchU/SBKHGHSmq82summ7q
PQiUYZUGtR6wquC55qg7xZ2QVLkfG0sc/Q5jFMWh25dJuq9OWGuT+sw8B0dPZ8wy
dNw6UJNfgqtuhTaKPf6cfwq8B32KajFe8BO/eADLwNvhxV8+WSaw9f88N+446nds
nuw+NCzn/5mkzDF2edj8o/NhGt0B5niXOEPmHu28Glbj8WLMBHbOvbq+ua5F1OJL
qtJ6ZQMhJDr5SlQdAqqLZrYP6+WiITkT7Jzvig6YMfDveNj4Uj3Q6lgaz9OWBDnO
F9/48QMSiUgULKOrjXZZgNuuny3GoSFYIR8vuQ5U/LTGSDc07k9+pc0pRIrUcOIO
ZHRz8vtGqgcCJQ6A+PV79T8Sfzk+SPIHuFjD8yyoWITuSwyYBKtneMKokFilt0NR
/46k9B0mIeMzE7RnrwZN5OGDpOaDCE1xueRo50hSSyOx+6PhCInzN9l0bVFdwnns
jtz6GsmZbfFPdx/L5vKbbBu3reNMcXrvh1UBo8QNwwcSi3g792Z++feURYWi4OXD
XvXqAR5/YIiVUAenYqV5yoO2ZShJCZLNzJFR2s2rQTQfd+Kvf5/+TmaT3XeJ6n8H
v/gu6z0QyByBp7GYdw1YJnv/f8qcMuSxnxJ+BMsIKG5LeE3iq+zFN1qi/GTgQNdL
muROpOg9iwLnMAArtbNiOjtaN+LFonZ+6QIlP4pehxap2CXCFOrWt7+1XEVMVzLB
/ii52Mhy2JqxJqbaS+i8mdZwzD0U88NZ/MK0F6KVAKpWAo9QAOJSx2vW4yF7aeY2
bdkzsDz1NNAhyZ5VBf8IQakwtgJZve2eaR38JB0i60l0cz4uyod0xsjR3GZzzhRN
OiqFSF0ErVGHy5bSyYy983Hlod0gpaeXfN3HFjvnugG7U4WT5N2snxLXtbhaGukY
bckkx9WjOsOMIvK7usHV2dxbqouAxMvAYBbAFVI8Sb6GItvI3Zj3jVB90zjk2kUu
ZOSOU7/aedt3OTd88anOrpznUs/Dh4EPvEwaJmZC9072n8mhO2GfcldzZP75eiSm
+xRLTI+sgz8EttRIUsi6TbvY8MPMX5ddCsf986YTWhPreZXcwqpQvX7auRN/sftR
t3FYAwCOHQN2OR23/4YWPi5NzJM9+qdveDHAM/jyT+dVjD4WkTW6IWHYae5sD/EY
Jw3RNmfY40KEnz8BP5x0we2ZkOaXUsUaipGSQTnEXQggT36HJ6hcQ0eVgvuBjVsu
HgQ0i9mq2EI3PbwpJeNKWr0Z8M9gIcYRt/hbzr4W3Jt1F0SXXYvGxXzmZsd7eoMg
ftn5ndV7NVQ4vG7pCz5XdTJgo5xIUVgwRDrxZyqu5jRzJISmP8Uh6emFAMqXtHQ6
7jRdIRA7Tg3KCoj+Sz5qTPl4d3DsgScef8GZDFPRnNa3GAzULT+pyA8ZuLcxWrDi
qSwVWsiGlzj6qqQIvO19rwAnuRGQfUsuyFE3FvM1kBk0aM+fpgBDnATJMV+Bj/qU
lgDYywtJXpNiHjM3A309fWVThp4ZkU5QCXHTZLqFrDI9yyUSwEOKcvkrlrn9qyUQ
bXVOFUb7F1+lbyH11skQOA8BsoZIZJPVibWRoXchdQmUjebMGxssrxpkcOaSk6oA
8trFPUh1DGNdUvhU1P+envlTo4NG20TZuP+kc71Fxg6WBGHjoMI7DACljOoBvpuq
k6AQoZ9UZfvZLtUNI/jxzPtvIp5ds2R7BVfd97Vkl6IrmGH+2JsToave6KKYyCSL
Y83Kcrsr3GyX+8lKzQ7Nqa27yYTy7CACGm+o89QE5shnFTjGpAZfVKj+O7I/Eva5
cuV1lSHH1Qjpa2JVAZ1rrSQ2JOdnOFuKhWpuAwnas1wRmu7sr2+BiF2YeApUphv7
nT+MNLnp16Y74oK6B+jfH2bvqNl2ApB1Ti7YZfrfNbSZgJc+oO/umVhTN6oqJgCf
dvfQxoYehT+7N2JniizqA1XDRy4BzvDB9rVtmHT3+QoWmPeqsTiMCjNXGXNocaJ/
c6WpHACbDGXN+OdMQMx40dIibnb2YW2kqJB254oYhTyD5TRUOMFpinm9frA/3ISv
UnR6EYRwcorEYAIyYcdhPJaBbHnYN2lvyyXAsqcnEfnmkkroJ/sxyfBalDRODwT9
Iuw4H8BdZ3tW21cwoMZzzUxDabZfkpW8EndAhyKFIhZo1CO5rh1R/VDu+5KD38SI
SroRkUQOCLjJvOF89NOW9NSlcTqgP/1E4fsVBZvDRTe6QsdNv/ac6GB1jGN2qelh
bDk5wE88pZu5qiEplg6ZRUaYke7rzi21oH7Q8VuN4UPeGH6bot16oE6ToxnNiz0A
CQxHE3TXqhI5hoditbYsRm7tym04tWSP3vYdtpNGa9srgqvsYRYrA+irHartKTUF
toRv+RsecybPT/74srWO/iZQ2Mwo0A+Ehy8O47tKRmRqCZRinayXwLDFKDgqEc5D
yd+MqQxUQvrbacpDkVdvjcFLI76GtFnN0K40S5l9q1pCa7wvTNe9jrjpPr1Gdo+C
jRGc/QFAWAd0PDSND5kM1rkKQAgFZCbcqN7Kedb1UcZy2j3bSYW2rH8n57/lkoEw
C/BxAanNDb9aLUu070PCKjhu88u9v9RhakMsRiZAMkO+734tld2cDEowP8j6qaM6
z1y/wRy0LM9a7XJiQpD36m4NxSBIEzBOMTtgbLd7LDmCSvuL/VFWUBnD13Hrm11T
sprVhHCClLfGkRT0rcH18iw8Rs0vGWpFbXhYWE2lXUSaOvg0AUc2V0AUffEIrc83
6X6cuPpx7FspQC6Ev+8GYnFOf4pjMFQGBeny+GBkN/9vSMa4KB2Y+aqfO1uIMKeV
zvRC9AmOWSwoOCfEGL7MIJrq69DgZGIrH4bso/dyuLv8StYKVPRga+sUwCFjm01m
YwFz4LHZ8aFN9ybx86o1yDosh2LPq7Nxr+GCByhvX28cZFCgSDpdVyZS8NNtuLi7
TZ6koCe+PhC87Mcv6b9kYdp9fSWrtO75fhh5gS7oV8tfbTPW9pCzM643aoldI67U
xJQ/ysGh8BFCStUSmk4phKn+73F9qnBqVe/5p8eyBGp2hRwXh+d+Maf3MmbAGjys
83rxPGu98HcmL+c3YP36PPwYOOKZd5wQ64A7xdSXWlIOlrprYUMtCxNtUsCIIWax
epw7sRIOAk21iGgVcPoiGBVyGKk6IAZWVSPoxgVqBmsJrE80XX84w88U9O4nIc17
iudJQK5zVb/G8HMNsJHMpV1O1rqOBFg0Sq9YZvmzKplGBnb30yZ6UZMguvwStUpQ
GJwgOAX+8stmNGHHsVCv+XvRJgVkcBGGvy2tT2vmtGfCZkgeRfsPbU4NMfmIdbW6
ikw91F7hs9FUHYOZawEyvCYUXKSo+otqxwuB2++pcPnvAlp3jhE8ClwfJCB2QgxL
VcFo1k71MnuVDIzOWXDzo/MIiAivN8+bXL50QBNrJwUp9ls79uw2wafR+4uGEu4u
rHBpelZga3MTVCjheyiJHIyh9yIYbcWeTfxEJXP478+h6OQTjWRz4iU3taqQvewL
TCIJcm6EEJirpn5F2QiIKC1JwPnqeE237cVdV5DXNw1M6xlaSMJk23HkgavyH+Ce
p01a6MXFgSRxLrBY4nh1U+GMM0vnKckbsoiRO91ZNkOgOwGuL2b5Ww4sxJLk/YOe
FcHBPPs2usZhEKBWlSeR5cWAaiwJ4qPvtAbdKxvYMQsWJvxV2Bc6gR//qY2PXwl7
BDSX0zEtdGFcmcpoSxScwyQAkVHgIWxEe46N9/+TTumOxnMS7W1CANcy8Qg0gS2E
4/XH2pyN9uv9zua9Wzqo08HOhI0Not0R57v+6xneeGX6grJr6yXu+/ML4qAh3Qf1
nDGWg2YVHCgTDYZp/FqJ0Xl8PwS+BqAvB4dOQAMjiuTToknkIzOXaYwkomRfKYvC
eYP//mXLSe43SrXQJfaKDXTRzB3EZrv33FhoNEGbiNePNXPwuv75pChWnZ4c5e6Z
NLVQ2q0bEMqoyXD4qeDmLAov1Zd46+C32kPTqx+gOucedRyxrT8h0YqMpJR+/2Vo
/EdEFyemH6Mgyum2dEQYMS+pNr5bWKPoy7GAX82jZRFKKtkSp48wGB05omjlzhS3
sNZzUcNR6ajcMXj3ZY7OfRwuJqwNRvodJHSWTtcPk493t+mJtuKOhB6n0VzLeMJa
cZs2nScjD6PV/KQM0o3iSBZaoO2/+XABlmvZko2DNr4doEqSrtu5fZ0p2DkvCDov
wAD7D0ZamyRREeQ6MFb2RPrUJgdjQ3kGS5YENFEWudFTbQtF96c2ercBUWNTLsKG
aojMPNFgjuV8DHtes4U1D65KjhRy5avPicrR7lzwGqjaCSmNt86voUtiXnD3yE/8
UDY5BcQa5c5dyI1/82HbJcfnHZCb8dlf+wrXviybCrv5DfRk9JIGaW4+sN63umJg
hXnwOzha15MktrnSEo3n5TnRGkubGItDc16B0jDD1EAWPv6jQUZTDax1M4H0KRj9
nVrLMkSgbDi8HLtL08JhMgaZ0i76GJ67VBKPCeAl4LPWbLKBRBj/kUogQkaYOkBq
cIr4mLeEr9RngoMM3+XQ7NB+CizRrdjzJcqaz/TwUjpqbYwyOVLQ/y+wYSKrNuLQ
PKXgX6LhwTpXTCh0K00P7g9pRya7CcbJgEWa0DHPHFMfe+wHVeKEiFAULNjxKoCC
7GCG71itYCs4tit8zprjb3s+21WiNuRpvgMpbKmlYdijtBLUoMwsVjrrrewECtH6
nNBHXY3ZNP8gDc3Pr79SPVxXGuLuEfEdBakbUJPOTx8WPRrSN2dCMaiEvWPF3Ys/
2gmCIOjo/VaJd8HZLgjVn0wKzYSNzByruquevPynMals1Sc7Kkn1P9/MR5m1XApO
hg0sjgIvVNWABQxxtAfNwyk70LQKSezj0clMiAZ/Asamkj0C47HAEWDc/dOC6/C+
hceGmmuJkes83zkczqLgRobSyoRNP1jLs62oLvQu7zBXPgK8o4/dY9CaODEYu0MP
4HMdKdIdbAC8z9oqIs+Hve7S3+OUjmjOHnPojwcUE37GxD0xVMARi+6SzpdF/4+b
ZaOvJc24k2xNkE6JyyObVO7fG6TfWwZusfAEzYJkJoT2J6MD2d01kgUHfxWLYF3j
30tMKwSfrXxou/oRIjiCxHlmK+B23jKodW5HLKJWbVfGt8Ficdhm/pN+6swufIJJ
UKJyOBgGp7Ep8aHRLdendpmVTOpPwRbbjb9+6b4rQEcppFZkQ9n9EiketYiyUIfC
GodrfWfedH//HgP6QCwEv1TTigSLOKF47GIW3lbkFjQIlX1fe2mTfi3q1JGh2YmX
ZEMPvQhwJFisNzk3Iusyy4Fa+7EpqzglIZnAovUnueU1K6x5gBFy2jXjqlswiiai
ILq+0QYCYrdfLapiJcxPuTARXVTjG3uqIp8RRhK4UD3MnqN4PPxkLEucPGYzYWaf
/IOsrM8LxHUhu7t3XLEgksxhMT2V2JfFDw7Oza8dXfq1f17SF9cF5ndle51zyTZZ
wdOWrKUfPdCfFjldFHgSzuBG7zJBTjcyOFWpljiNj5Hgv+i0SWN2fSyj1T79j3Jm
d8QLBq5jZuEhIGJtZ8TJysR/OOwPNqpvxoc6X1CzYfdnJKNDurqCTL6vPaUWasCZ
Eznq4cNNS2NaLOtfqFKtLBPlg7pnkoKdNGCuvu95y3xvGshp/VpUyHUB6QQo1GmO
PgoI2Q4BtOmjfldIkcfqFxq3fhDWrV1ivsS504vJkEenhiV+ZPK/qiZqDrwB4zZf
LbcjNPjholrf0zQeDxBHfZaWhF0mXCEVLxs0CWXu+HZvVI5vRItvApGbfRRUYLgw
Wb4eIwOG5arw2JsTIpABoHXIqFUJX58bTfjjg+kySWOO7vUlm9w2aIwm+MGV9hAM
bkNSTnmvnojOGJNgmPnKJIax0N7yDzT87+DzWJ+YPZQzUnv+wLledrsJx4KVKx8p
5wk+6aHdn6+S1KWV/Mg6oOtON7NF/8piUIqZqiL+w6ixr13F3J5MaO/InAWrIngi
T264Sj+tGAZrZwdIO6jWVGnBW4GvXrXF3qIbzPOb2pMh2ZqAH/QpIClJSHa+Srgn
AhCvzwVPj18JHeyrYhMR490y4UxUuKRYlTHR7MRk7rb6tOBsU1s047MmvKVjffKJ
Nnty+amGgy/oRpE6hM5soi0Okz8Uo/vjwqCoSIP8fKoNHzs8cCM8B1+km+LMhXJK
JZ43hRCgdJyEqbQQwIJkQuj7cXgLCWxFO4HwgNr3jjQ1ONnvl7gyHcCzkqwI/J4X
HQt1hgeiUg7imYRKOnbsxGxsBcq12m4c4ZZsOS5C8fmbG0Z8enMBKwvZjPFCaLk3
kz//pbe1ZH4zAUnMgUG5n9ukyQrNf4M+AWPjCZMKCTOqK1u7G9zTfQ9t0MPxdoUZ
gI112I5ZhtWOMOg7P0q6kx82KunZ3nUo2nmQQdHYbBjA+RoOV8K60NDWAFcga0KG
YZ692yG7pGdBpd5tpzCBTO+FpxyHoqlQWyBKRwDoojTXhbab9bjK94VBSRQs+10o
/lOumrL4pxKypTS1b0uxQfMx5rJhNKMYQOhocsuzmYmYSKDzwKD2c2KWHTEapA1n
52Hmn7MAOivGRrxs8YdAAKjUKKy+UiztXOUeVxLZ9ww0bFrA3INhFiQmNcykzhd+
/onop41Yz9irLHQhABYdgKktc+nHX3uKE0+sbqrgeWhtHDTWmWgVuLaFwNY31yiO
DdQJxG1LMi4k0RbdZIxlgTQzAS+6A5HAAzUIZAozC5V/2QXLsH3ltgvUFEqc3Xvm
R2qHvFnLs/++hn0SYfeTArTIdvgyjU/sK1LkLJxslOinifABvRhNfqtgN694YN7P
JgOjFzkinApLaEyLa05c2Uunn8XrgZqJAI4btBiIF887GarDgBL6m9sEyEhSDHNF
oabJedhyZVKwWhWl/eFcZnSLBemnCoyDC/M+HrMwm5dswBeCt/LrRLZ+/R2bQ9nh
iuAAcfBX/AbUI1cRRWBpLdaodrfqCG+9OvyWAXLYk10h5ffybHef/RI03ejeQ39u
i9r6t+sDH0X+FtGptBrKlQ6W6f50NdAeURP+0Rg3aHSp+tw2sVLzhivgA6jkcN5L
prS51sAfvlNrMh2IsjM66SROpvzekfp0FS3z2Qx4Z3SMftcruk7rittYJ0v/m3F2
qHHHIg19tYgufR/fLNnEjGuvoN6bYOSvmQ3aMTZddcLM8up7k8c6unh1zpoLMJqF
HPyuRiE3LtaPknvth2qk75WO4KhCnl8zTLn/KMBo4VMhcKCqKq+VNS9OOLo/mtya
jO46I2eCTsPzGIcYNUL41Cr+LlBTNQxIlDuaoNlyko3/8WSkS3wq+WzW3YxISR+g
TThazVnQaldQ7OzusNg5xtWK0KJaHEMqrB/AjlxE74easy9X5TI+OhswlAu1Sawu
sInA4kqJTxFFHjpremzjcSMmh++o/cUwkR/tCl/yhTkOVGtsL2b9sHdPE0JfJ6t/
nLEMaJT+Pt/P5lIhyzX/9L5MNzAHT0SgoXvva/JGzaStVwp30f7zeQNk6mxXUU/9
xcrOxyoB3Ry2VmUtfOFAxohb+r2gcriJ22DkFGRuS2WxZ0a/fl7IZxGfigN9SLKf
+l4iefZGNUhxZs6t72BaHI7WHxXZnaRfdeJ2XJlidpJ71KzHJ8Cfjf836ILTrBIt
PoFSLYQrS1WQbG6RVAxT/SVDqgTPN7guzGDTT6jnSSRlMlcdCT3hp4K6mP7XvvG5
XQ0lZWk1agqfq+Nq1A2tFAKLwH9b1Jq6EOcJ1xEmuzU8ZmMUtpnC05kbIM6ou1Tm
XvzX0kkotAbhjt7+HManYpAnGTgXsW5RfSBMuOClH9SJRT35/SFWscu0/7fo19Z+
fzfaHrKAI1eIhvDWkW/3INj7oqrJWXAy23SJJXbsbmNbmoIZ4wj26fag/BWkJaS0
U9XspUMqLtpxKfBH2cWVuu2c0T+EQXVG+O/n8ho2yexPMV+cU1KLu46HohQs5YMs
O/pLcOjzn1rfynkcqlSoKbyfUIOYafaQHiFqmJzvJeLfpJCoDYOP7sqsNJBxmxdW
5+YB6vX/3jCEl3Y4mI/tRTmJHTL5J5zXCO94f9agp9DLkdoumlpCdWubfYjE8L/F
nwfwzAb8E3xo1lsLRdajpGU00yiIMQ+DSk+Ad6Y8VKA4tnrN9HvpUmDTDqUbUNeR
h526RF9uDSLqIIanoUOGmnVDY5+QdFULASAqFE1lo6ZMdAgpRmfTWX0S+fhghfUO
06WDP+z89fizv34OgnzJKDTDDQlHJ++cgkVPXknu1D9zxORVriUpg/+21SKuh0fy
C99lqu81QvbuLlberYh5gYz7yExoeTiG/v+5VXHpHTLdweniPnq36YzAGxzb/V2B
aBSXJcQrGPSFjHw1yUfR6xdKebsp6qXG0U+lGDfh44jBkRoeVYhG35IOqykyRd+z
R+wKspT62B2rTav4ZySknD36EEUOEDx2Lyx4PUHGlZs9g3EN1IJ1hBmBCYECx8FU
in8eq/GiObmEilbZtG6FjfHxT7W2p+n/MORDC7bbJJvOQINcG8rUZn8jcNKT7iGk
4MWR98ahMRorvCYtHZJ0T3m/Q5IFnMUwHo1zHM2Ev0aPQc9ZJYUAl9FbOSobkGl4
xyonq2/SYls/Nt52kLaCs/wuGEHcum8Yd9VGhlRPo7AzmDqm82AW8R6zfWg0i7OZ
4mPZ6MQeh5ubTMpxBJkteAc7IZFyoT5lVH6IgDhgQcYW38CGvfTGqUcQ0hagD5/r
D1hVaUIfwnAFHUcX0Ze1boo9w/e0fF9IrPyN+IqmqkYL4RBWeTRIZ1VGfc8mg/UZ
S6yVgS/CPJrXiPutB8nMIEAuqpzUNx3/TesJEbmG0FcgJyKqGLFoNQYdkNqV/PU7
D9BnX/t2U4ZfUSp5RogWgQW2lRfRGoU6Cfd1MD4j/Tig0FaJLppSpXOPeGbASS5s
r/dwg6fqDeKHUuQlaSGdqmcgH0lx9Gtfr4jCpnZ78rDOoKJjpIdpA1OY22//OAiv
uVsm7vIQzOL+pUIku0hs7/GjC3FHiyW1LJ9dtD+iSQgFH5DhVVrs6uFcPI+1Zgfu
iu7KpeGlucEOodDy7wBcdtQq0nrgJ4W+c9xvW4fTCkV/zIA32Z8pr9ORPmu4Ct2I
QFUFEzmh3m1vN+jOmw+v+S00hECjy6CC5pvbyD4gA03Ka2lwwahDVTU8Gd7Wa61A
5xaqqmXDHKYFd+ot66DSQFzKO7PzjIJATJe3R9wRZDACHmyL3WEk+9ol4qjBm00G
NjHmmQsjKonIH0Y/3Xbh+nYwzKpNP3MjQ7+kZUaE/ZzAvVQF2ylepyNPBAsSOy6u
tL4tO6P+GzI9iVMs1F8DjBBNXOywSc4UwwLwndr6cFUcvLAXJ3cjpJkEFpkIXpZF
6FYv0LE/K/LkEwkx05siTAQFjvcyU6lDme8GPAd1RjOi4X+bkLjn4tN3oPjDcY9k
NyPXRvmYAMH5aqtXRjWM0J9cQnud9ZOtgoIqWBwVt86IQTtXP/n54aLhWWP5DMjW
+SyCTuAkPeCHgTaviJcT7+omt2ND7tm3Ov7ETOQCrC4kfV4U9aks6Z2x81ab1Hp0
//5w0+jsPyTzDQ+6YMbMM9ag6xvsTAsJX+xPXp4qluqAy8kFgOymioUrL3FGoQc4
kzjqzYZIJuPj+BarLbRCxe0noui5AtE9R+Is3sG423+mAncrCx1ywL6cRCzfKS5Z
kw60l3NA1Pvrb2WTRrvB1/Re4kYWl05ocIWUUBKkOA953jmiC84U3V2p+zeRqlEs
cXzaKqtjE2QBa6mv8Ys8tiNV/500dRAflmHMgTNUk/zg+++A8oCejnrbMxBSXVWM
3R51G6BWhCyi5kFOosINpI2/Hz8aTWdAF8awLbrTddCs62NoKIeLULwaOT4tutyS
IXuXnhZ2SwQq18uZCxC1HGWFpzj9Y9EZkTnEVmp59Hy9WSgAvR3JF1CGGvxODMO2
hqKBgJXxWLwo9Bhh9vs8kwBoP54m0DY8Dq0aPhJH0To5G1yY8aaKCFiI4g7RaCql
BFI72GRoWb7cjW5BWAncz8L/jAINhwgEZWXD9gMivLdgDbZpA6ChAV486f27YsdR
xtxBx5iiDJhVLdpMRSs9rxdG3jJObkQ+NOOlaHElGKMDUs/yNKLr5tgfDC4F50Q3
9utjce1y3nclmohrdMVOfC2T59Lc/aOHHsHMbWn7q3cAa8rohIeIHlP34CUNecmT
/x9UjhQ61vk3lUyAuGThfmlQaBI/nmZj9BMSpi1yPK6oN1N4+sHEXHM+P8NOVCvE
VGkAWF1BZKcLZBsbRsJh38L2YSVHuWNkyXY5ZoPhL3+sJF+sdFX4E6/t/0jKmCIA
2altk/9cvycALlyq6ruS3gQG+O+qe3IqwnZlBpNuQMVibNQnlnd7ZKDb3JboNuGt
HlY5risA/q1jqaHgM3LZTDXxlv3GHy6852umeF/DKgRjM8E228s7RXfTUYr+dTWs
Pa2q4pFDJzxKZ9Fbve1mEKsAJNptnbNpiYeFBxVDDh+KKavF670EypW45Kkj0gg5
Cxx4pw7qdIk9/OeHbGRSwFt+QSyQSZet+7aPXEzK928qSekgLEq3I2kfZwxPGXb9
JdUjClQvsrvyeYdpS1c91jBQTPvqLcyhTvNR6AJ6eFux8el+TrN0cqvoUuw0Yuha
BQO38XwhAnyqIPWwHWzr9ZA4zLdoA5ENfWFcFSNZaLwjhFXmh5isHllgFyU3YhaM
xF6JA+fWzjdzVxb29PR7MJNAXgkoDwMKltZZ7CwhzYmUTVQMO5WCpAuZS5nJRM/d
3XhrElOgeJUA7ztiz+SMxJztgbWzJPSBHi4E5niqNeuvMZMc+OPnMzuFgB6zByRg
j3WrbJ6GvWU2nVqUwSsaNKi7ojHEkQNV3NyG/AUAIJlD6vT1X5Aps3YaFbimDZlf
kHvB8aNAFNyVJOP46nDOTdTNgUaGrKDbsxULE5H6CS4fKcOSGKAJFe03OLGRshNV
UFkU0OE6R5ehNinMhUgicGmbyAO3ggFKqj+yjdSOdYHLMdIdhd6gCk9X6IuhfYTN
YxvAZ5s4b9gcJKTIB4rsemBlJUGXNcS6VzLj0WrL6U6uAPrVFHsCyBUNEwc6DmcJ
mQaJ/UiTIOVU9EpqBoOnMRVhiYdEj4o+T/b2e79UYp72sxXqo+ENBgeTgaIsJkB7
5ZH0GCcJCtZI7Cax5PSeksM7M2xIyY2rp45MVl+iLC9UMyZtiqxaY4uSOdC6oEvP
CxNJcBy+WW6tT1ZKZJMsooaS6EoTpjcUvcQjz1BA4mBVO/SeTYhKGh5USoLKlFyM
sJ1nDkCP0jsrWl3sVmCPbwt6wL3YFFY/Nnt5Ulb/unO996VMZjrusOyKYES41Nb8
TA70WKYUYz0GVmpbbK/X+s4xauyXJs/2gQrC2mjhjgJ1ZImkFfDbplBFdBm2BN0L
FipvixMVwLYVBNoOtujs/q8jEnxJRHgA/TLXibY4LE36yF2jxk7OXmvhzBZoPZOY
hgvDiLwXK6xGaS/D4Ohd7YafiN1eU/xkxK4vZwLiKxgbC8J8vh0e5PvZWAskBIO5
akmVWGSV2TfdoH4AvxSjkAHc2Inp6vL0XwWgkIPLAk6qOWmy4mRB7AsjmFurSl8d
rT9Y/YBIr2buac59ubDcbhLg0qQGtnfToIDk91q/hbEb4RK5vet+TXb0RH95PFcE
6KWon24CL+CdLDWekv/eB9utuMfYuPCKdyA8sh131v+2dQKEDBJ4z4F1mMgY1/rE
tFQhzXKWGoLdiVjQf9WLHFTgMvxDnP/hY1d4nFGUDKyaCFJWRfSD1r3Tn/uPyoQC
tZ4xLq6xAhm5d54qhXGJ+ecyt/Op+6IWOM1qbDoQUmdCtyNw5cSSca3rt9TJhZTj
s+qePFB3dOgBFUsHCz0Jf5qlCXUkNn4vGxygOp1KoTVZHHbR2bCxU3cb7XP5eyia
crL+437Pa1myp5BpBjHmVQyh5Lz0c49ZCdHxwkW6yMw73aOSgy52vSQcuFnSCMkK
kAE1fbUiaTOYp5z3sfnr7t/jKz6rhraZKBAMK57u4sulczEVCpwiVzngsYX2rSUO
tj4NEQ3g+oPCq5TXUf4Bn+fgUZavjuqBx+y/kt1FR5+2hWOYjFMCO1wUu5F5ZZnG
GEbuuwuOI2YcjIY4wicf+g7gSOJPBvYTNONVbF7bSAKCjWaJ+6Uvqzwx7fr8gtan
SA8cEIXR7niUoMsMIzxJ7zI2rK7DaKqhRf0ipdS5x7DHD1jHPVlN/pRenMZLwj0/
Z6eItEPYMEr+3JvoZYDpDr2hIjD38Fzg13UqqidkFnTHZtoOLlz1pohptgJlXjCM
ZUIAvbqyFAAUxVUF6Iv53jSvqTQxfVhZPyKKPtbkCJ3uuB+tC2y1Z1X34fq++t7X
jpnfhqJcCgTWIF40tB1K0Z0fhW/OqFWZklNcF0vgQbJfRxHJKosAH8x0OZAL57Mw
2zVfwT5VAxl50jwMzuIm9ySYVOm1vVqEn4QPxYTH1n6ydMx/rxYgvHfMHjD5P8pb
V09k7bJVshpt6pqAKnrpYOF7MBm7vOvvXIoFm6r/1eB/kAQ4KK6ENHm7IcFaQq18
GjHv2puqXUbbm4fw/QijyIrVaI+Bt9Fqh0jdSST4uh/pAaNT0U/Xgx4lvNuSXpVP
JH2t25ocfh0Q/i2TbvhZ+1CmQrXS4G6pFo2tdwYXrldA8aTaYLUsQkD2mLEZBRUn
tGCqx03bQhKdlXn+WNCZIAczixUuu2bBvyWadokEGY7uZ6UKs0N+iKtyNPf7UbLu
xxFNS+wtwEnanhTZVI1Q/N6rJnYjQbi6gjziyuB4tk1V6y1jwMhHpUMa4Ge8SRco
Uebx7LM1e7Qjfwn4feSa75dOJQt/xuyICXJursp2ubuD1Ze50KVvkFAJ/rvohA2t
qi/KlZaFjxZ6uXExfLF4O90AybYMiNiGq/NqF0V5YBvZYz1jh/VdSVX3s/P4BT5T
xw1XInzrfq0hU9r3NidEn5MJabluVht8FRbZUGYFdeb/aTLDNhkJD/jsO/Stdlmq
w+g24jzLj2Q7zC8KSJBceGPLNGpWIt1y6Lvmb8R+zHadBflrDTbUH2QRU7GvJwaN
3gFNKAJW850sXfJ+m13prYB5S1bbruYDNLBuUcQkcjsOK7uM1wo1AKLwWEjPOLuU
gzVMum9lGJp/sUysFckYEXoCugYTiG2LCigXOIgtjfKQadVCtz7BligGtS5qYVfc
i2qERoWfnJ7AbjS56T3gjB2Rk+9piKk+ZP8C16b+12n7GnRWYjHuSdN+eIy0D+B6
cmh/ZMDLtENozMz+1x4KFWOZTMGAEs0QxW6+sD+1c0fULqHTUXmsHjeqbnlNKPiH
8e0/WziMpc/LdCHm41PqNuSaDqGm/s1FKOtTSM6ulBzMRQe9y1Nmi8I2Wmw9ySjU
Pg/WcTfDZh+ZaQ8Z0nixUFDuMHS4TOF7o7SeqiDKNBBM9KHd0OzkfqGK0Jy0kQFY
nRpCCUKoaxUfOL6tqOqjDFI8oHKzzu505nw7n3ynO502Joyt4/jH7R9ybuUrdqex
UBpmrOHtJzF01nheRbDV/Je98Ffd1jOlWVsuEq05u4fdnV9oWUUGY5Dca6Xw0s5A
nF6S8aW/ftgNxlM4GcD8KN3is/6M7pxEJFsKwVaF7e8Ohi9+kcDHtdP7rh/VNmn1
nZyaIT91jAHYixVZbbsrsdqvhppblohyS/LOptWqMZ06NmK1PfrJu/7MdlRBbdYE
70UfKvDuyqVdUfNb0Ba/WYmW0icXsrS81R+MrDVFCkeyfY+rAijmsUeB9cEjaPvF
NGqCIge3Dg4FNR2gsw2zsoErmBblotlsPnMwvPq0YpzXFYOdzqCrl6/qCY9zbh9S
VcX3d3Dlipys3IxHT04Lqb265vA1MJ6tyL88fWmOKwrokJEiAeKyZcJd1xtMNMQc
Wxs0Qnh7nTD2K3w1ZHHa2z/cjN4GpAb74mdVLQcmnYtPz0zis1f4cGq0R4qG89lV
Gg4meymXxY61FoiqaDQ+s5LX/GxuHLNRodFwEouody+jGhJYwW5hE68MDbz/u4aI
iGzmRXLjUNQTD4hxmsSXUsb44ZK8g+4gHnrVd4wfWWS0zVo7J8hXyI/GcbRtVFEL
Zdy12iU/2zChxHFy7sPx8NPG0uPSy1JDaZRWE2NCXUxWOw6bzpms3d8/2aHE7nAg
L7D0cSAVLROvG2n4yNa8Woy9ZvDFeaORbzda1X5sw1pMwuxIQC7V6whrflRLE1WM
IpMtgOmxXUkgUAnbSgP/W2tC17snXyEKdoGBdOb9Cf9s4aV53L68Mog1tF9YBLos
+kxguEE3zsINevDD/4NIYHdv/bnudvpbGMhc9sDIH6wAydmuH0S9+QieztrlAC7V
3YZlYrt3/v/SSSVXHhewDiSVwkVFQukWYZBBmchIhHnCAmaq9Fj1ze72Cc5Yn9j9
4V619xWk9oVDGlpslPNtRXOmAinpZthTQJm0V8WzFjiWDnw6fz2TwdUArCursD99
1L4K5jz/+LasnFI8MKdzXdeIxgyuMmyhM/ASXe9qsDtotcFOdm5u+yB00Ts61uVb
mEkQuOvhOmAWR3z7N5v+/vEnb++wi5JlR90cYjNx/7H8PU6T9WEYiLXaCPJh855E
MSbSHpz1+zComF0SqERtdIBqSquMPcGQMAPnKti/lpMLVdwxDaagAYq8GEBRTr4e
ZaKkD2M9M0VjRymlkwTTK2J9ubekss0u2l8TR3/jQNuNfPKJ1bUn49SxEUyEtJQr
Or0DTII0gAQ8zTh1Gcq7rg3i03RWEN4/LyStdU/f65ozT19w0dEQU8hKDnyKPesM
v1TJ9cuWhKaj00tUI6TQYi8FBz+2XC1h63Ot4uA0EghPV1FfZmOfDf1YOZ+vUiAt
nQm1/UjVjD7ZN0QY5Gd5hQ/eFjl5DbqACwvvn+B9ukqUq7MXVFZisMLUo2YMIMQ5
1lglOyiM4UH1fsaBmVsqUY8Z734J68V3scSsNGp6kPK8+xRWeOPWF43LsoBD7tEw
IGz4B3bYAn2U3skm6e6mq9GliHhD7+gXfDose8PL1W+3wW7Gyebkuky2uOdebmmA
Ip9782ikIP+W0ekUbOmOi/KwIShuJllRZIBMCFCUBwGNvHlsp0zWTm8MOec6/TYf
0pJSckapBDvhgqE+eQ1od0cuM+ukYcilBQBuQS51A+88VPGMkvtLgEydneRWc4rn
BdmDGGkriMwVWJmoBZ5TC0Wi+37DYA+UvvW1ayQfpM4Dro1ze0rJCUaBA6Lo1U6p
xHT2JqMlYtVjQHq9aad0xDcLq4YKMMX6ewxV8g9AQbtUtqhHV20w/vMLDfVm3hYg
TBXZ61jJyniCa3boNKgmhKMVDI2c9eKlHokeDvnaNDsf4zgOXj1SsZZR+Y/gQ6Ol
V/0q02m2uCrVVWASYXLhqbaQCMvHP+t5y3TPA2j/2tNZQkgf3xf7+/92MfAJHnoS
bpqWOge83j3QhK/qmDsX30UdIXc+tICD9p08M4qJyh2C2WxUMS/Uyajus5O2TuXt
dvqh2JQQZCOKclBG8PYojSRM7EYKP27TvRPHBkrZ1b5LYhuChwac/hclCD9IizcB
l7lxVqIRfxgTl6nWzIgbc0qiRmdofSb2aU5RtiExDCte5Xav3T1pgIeyVl3OCZuL
ZAtZVzdja31y7ynPZgv8TLXnEGWTUhw9BHhdRXnMB0WwikD25PXdJEx7jBZu2rxi
tWSyCluwyVpXw7EbkwKqmA01xfCTb0amfHx8MaWvOqM4OiCz3QvVQEKIK6f8kVLf
KHyEQbkXUItVfpe+4hDQTdfINEa4M5lmEuZKmTF+HSXx/GLRgM0L5bIIl0ca0NVr
NDn/5yZ9t3v9DKuqn983aouSnGVZ4k78VT0jrY33WQfi/wHZUTsRZHrDCoQ0zECe
rOsbG6jzT26kKLu0K9k5k54yKTUXsWyJpf4BZnWEpj5tOPa3fkihDqEH9Dm3AGMO
/IVnYQanXJvZ7DURR8Fdzm+fBFwV9LlHkRf3dxIgXlSN/6c5KkeuTBvz+EjOtsS9
aPlCV+WZ9dGi6rsYVEzg90p6wjgethWQE4NM1jMf6A5/3Jm5q4UJNURXBxekkbc3
5b4OARXqUsv3uKoGVy+P/gkU+EfWQPHMbSphy1yEJ9SPw9e3SBXb88beIiJk2hqC
JuQ3sm0WTQVwHEpUrlK95TIOkca/dahsjcD8mlWf1D4JV1Se6VEft0iW58qih8Xg
NvbLtlS7K3Ueo7qV/kkGPlokti/EVCPakH1jdggmThif3wui/VHSBcLpSH+xabZk
ZeSUZGzcFgXE1KTxLNKV0b1r+uayaGuaO9ZUGhwHWogc9HQDVBZuIabaFd4WeHen
UwoxpUB6jRNO2LnJfh3W0TYMKl6bBIsi83pMUSI9GazhJjhEQVAcH2YEpQ3BNEMH
h+NZY1bbiknWFRP31PMnWN32H8TZ9QxgvVY1QNmJ4fswtYQsMdkLr22Nj0VFPOcB
BH+1L04xnZRYTsS6bbMcDZQaN2PSLXvHEr7oeTmBhedlbsJ7UG3f0TUjrxUffcCd
35Ow0/wr6yEgwBxUfjzood/oAp0w414ae3QWN1wd4HgkumhjXP0n9uyFebZjrvi+
4jTCoWGO+9gAhT33JcfXAOFHaUVnkpf6O8cw6H63q4GJYPgCcWgahXlvUUcKcbDU
6xk9CYP7TYs5Kihudj0Oc2dhWbN7WyZ2Ykg2RdSnxptK9zozl/smZO6lo6XnhtcW
OqMEn5Xn8UcVRUin9W2eZpc3S7cAx6+Z8MvEQ79L4xZic6hjCDqdA79D5K8/9eVx
BqMogKgr9Mytm1gEAbnk4SUB1nWTX/goxYWQ0Hl0pxuwTkscqkF8BVZl3IIoUeKt
imvWwlVpZjtaSOaVYeQcHIXkbMFzg5WHuoUaJ6nRfcj3mS1T5NmhngmS82ScWZ4d
euwfQgI3MJMnuaKTYv22vNEgDz2eBDkvwD2Na8qtT/y3PooX1GIeAlki4W1gHfoS
9Y5g6pCGGxb0+/BudQFAkiBtDE1o3hBspG13CFAyIxbZG3bZTzCGrV/ha8gmCXPa
KNw5FRbFGah8sH7Pl5Izkg4QubMG67Cmyw8jcUo1ogB/GPIDFBbdPHpgEkFrmecC
cPXKF7bFYx3E7tDFaDcWCSTl33EXYISXs5Fa2zpuEoGGrAXp7erHPLGaOveuHc2n
mXa3UDysXF2BwoG1Yd6ECa5LLnR9BfJorjlcnn8DLsnsmKY6nV2m2UBEk+cIJT3K
yk4uurRtesNO2BRCVYElg+tpoaTGAKFgxXpmn0JY03urxfq0UXUrZYESNf5l8uay
G1yNVChg2w56s4BEG4hPRTR8lwmgltwbwcZ/Hz0Y3RVClGZ6fJWWmw3K7atkZ4o6
EWEo3ZW3FlEoVtPhwjp0sMzgPow7id5YJAiFAJx2VS0RlSi5EYD+2iSxkh86Zlur
uHtTdBrq29YasNsggR8pDDreCJaI0KM/dLhu05PEB7TxHthMs7h3QrGB8eAqszH0
AaHae84ncDDHTL/hLznb5T3rA65QH/CgB88vKM/6ZETNvxFWRqn23AQFZqEicwp/
ZGNlio1tnsC0GhgUilb9njJP8CBf3XUp3CXP/bQYgzsfzsZOj4nZXktcOoeX48ZG
A0Tv0fvd+pMHdwIDppQ48HS5My1umWeqBGAtEV/cjEl14q4e0GICZOrH6fLzIt6S
mVgLfWY+A/Lp6i7R47q/mEeR0df80gDUco9kRTQHP/loBA1xv108hJhHm0Uus/Kw
W5tFBCVJ0eFuCme2aeYJkzjff/EWjvAHMKyX4LgqFrlC0Wu6vatBcOFjoS8T0pEh
aWkecnYUDemPo/J7oXyiXWGinEmLHzwDmoKKvE1nT9F6Lk0CPv29HAdcA+STkRDu
1GBtWkd+r9CsuGgbWgiSjz/2flFXIhxzuv00UKYMKgLPUkD/HSqOXTLmxxuOylvm
zM/NxGvgYUBObgPvSADChr8TE2kIturXL3Vbqalj4fhrrUGbl5M9GyOBj5M8asPt
DQImpS+faTxwWQ0Mu8Gy8/tzNTnZ9WfbQNRYKVTCHbHfCuajUNB9B6+ffGiwIxqv
dFy4eMrdmOinaXBvmgaOBxHEC2M87Xu8KVLYLTg5+pOjqDI2H+bs7OQG00FKfrTh
kVqczy21m2O9vzr6pIpDWrXv+bhRoqAN9DhXzfUgqm3aRSwUdY+9CEpv52jHsuXt
tpk3slJz8RU8kLG18KGgT+xSt4WhupvDvVsgPqGbAy8EM6iV9k50CQAyk4xJiLar
29ucqFNNvHzuRYRoR0b035eu7RKCDKoXCYtTPBY3EPZWlsCRT00eEUHP+HdznRtg
bm+sEaqDiEeLd1ga7DutGpu+4YxgnF4jI5Lmg2vrcwwmuskQI651BrN+1W7XFh0x
9MlcOVVGpQVz6CpI2KxUDH3iuYapg7fin6GyLpPDqe/OLTel9tOQ6y5k32hVbnVp
VuywLuNaFiDS4N26rvRKB+A/bGXeMo1kvEzn/lEpuRlFZz4OyQbstG599u4epPC7
K6qoD8J9pkaQMCSdSNF37femBGvOwX6n7mSMr4LbFJWNkp5Z83xyrCw0M4Y3iovz
VxruEiHKQfBS2V4e6uoH8l0MlNam8/c81vstOY2tFLHPy0xZevk40ZDEFX1nAaeY
tcLd2/Nw43WAExT8whfc1+p3jAqmz+FKCC3l72kwVa5Jgs8cDhzINahLZjtx88ns
b+VzZaWsOrDZMLNHGJlogJmizazzp+p90ZbXWqK3UFp1cilvchB52YWzjTC9d7yW
ilwPfahv/fdGKt/FoP0HgZ/dMlAaoQSTgxAKCfT+rNXI+sifD/pTlA/WalCOiwaD
k9gd3YyCwwPIpzQZJUjMVAr6tjD1Alw+iLjdEz+ZDAjpHtHPGi5lxbIgylG3CcFp
O0gLuZDB6WhTJ4DwGqQNGcaY7uf1B4++dfCLMQ4huSrReADdOEyuL1BYmmbTt31E
uIwkgUYwwFj2ZMLuHVKl+pensVlfP9cI/d7hOypiPpIPMWlM5Gi47l9kvv0Xm1vy
+CyGW3157mzA76/SYRR0UHlhgr9Yie9vbLyKZ3lsmEm/b3qnKmgQQCH25pqIPKZ5
Vo0LqUoYNA0CrDofnX0auQV9mvjPmxF05JFoucVmBCmFGwRl3GLgJouwUGlVUYYa
YeUy5+L59nXk+tWjv+aWn9tk04fuvGLV8FuU0cCLo5dAEfpINM+CNCN7pTNbmKzN
7W3+UHL4SRlDPzLKaSv0NkB2+0oldGXRkcng0J6ZBSNyAklHsLSqT9kzx9d58PNt
KbCEZaJ79QS1+a1zUzj2H2l3w+2cfCm60iquSQNl5OTOOywwMtqgdUmZImO5r6OE
L+Qc3XzLr4RG4QtEkvm2Cxxdx5rMepfyBoc6aJc2+M5r41NRJpoDvieVYQMDJOjH
9sg/DXi1bc9tqlmOEJkyck4qgizNInXE9k+OgoYiXQWpPhm6kKW5MgBANc3dufNk
ci7m3yKZsQXdB28I7UED8DEI8JfooXxDwkIYMb2XT+YT+B/BdlrC6lKUsaCMNSDA
mFknaUDAUbRqHlM5JMbxSLvGBj3j+28UQYBv7e9NuJVGtwF1T6/SdrSWnhRqCJ0l
6sKcVuuRW0epjzY8+ujFPca+RYBVFPIYv380V+dBhmsnW9Cb4ET/WMsV3C8W+UcD
jN2Y5K9OO3of4zFtb1b5R7RHO4k1VDwmumwTGO75ps+XNlF4rgpnHX7c/T3Jpj4m
Q+I5I+0/9ge0NYUisfUtNRF3m/RrRnkDutPe7ioC3sX7zEeJWiVE27xrARf84rPD
fMmEinESh5FgvNwEkdmImh4rrIVldQ+vfRU8wuPVyWjzwWIE/0KRAOSuc0ueYH4/
ZhtHjP20s/rN1katk5CYvhhVAocBM9zK6b9sE+KnSIGCODcn3+g25D4Eprhxn6hA
inrAn8FFh66tkXVJ8U5PsagCcGOVAH5gca4di9UxhzymmDgwjftfkb4pkVGDhE/R
PlbWTlH9yN2oG6OfcgHgONwHrVpG+vnEa+Rxy8029frXEv3KwK/zCF0skZ9tnyry
ZlW3U11BTy8KEc7jjzrt3loeDQd26A6gBl48yfxJp5+/LA0vFOfuJpK3w+X9+aPj
nVVI3yw6qAILHEBaGSaeJ7dUUTyxRlDhGcbpIoB+a7iyysUL6+u17Hwf+5ihHPvk
Y67CDe5jrbZ+Y3z97FzQ5PVVKRoDLSce0xYt6d0ccsHcBpIcGXjlSfXbRM9haHGq
WuaHVjIxHXwyp3xhiAVlISMA9Foz24zIOhKHtraDIBG25MAleep3JrmUCbqUvycC
AIkaNoa/EAfSsW3Rj7+82tnTO+QvDmTahIK6aWpfzs8/s37HPuOFd3CxfzLvyUEa
7TAIT7KbV+rqRpafZR5JadEC2qfIohSyXnYG3iQd60mPUwBL13gNrgWDH3m9koZ/
1Ityve0uU+pIIqIB/78463Mgmn9YRxOMxCl+6BgbVEQ/JMwyI/FLPVuRQBptnm/f
Nm4qjatArUI/ibhfTeSb/yGUAYxy7zMCaF8rjXz2t/fJl2dxS9XOrf8VvI800G6N
xarkyG8kDNpkc2IX2kAVFiWSUu+rMmnZgnsEVQKwE372IIHp1NTL3u6eNZ4mJXz3
6UdVPWHwn3YfBocgVH5fpSgBXijNRVZYZIsfcJIm+5y67PJ/q18KDFXlD6S0Owf4
jSIirGHSiN7N2D2Q/byKMt4QGp8PiNDa9nbir3XNN6IdYDpEMDOU6hhYVEXoS4gM
zh031Ql0hGBlaGId/Y4E1R9/owMJq8bMpJgJV4Fksk+gnzf06O94fo9r9GmWP+Pp
KC+Aggm8796RPpy8M+UPEbFZjsytXap7QCSPmv9TaKw3ppEN7A907LD8fC05UQAs
hTm+3GDtfcHvsUFFo3nH2SLfF0hATTogQoL/vvUrDzmOx17zHIfuIUt/9ppdhUzz
WCG5R79vXOTmwB/cwAj2BnssMGMNdnRxcyqtxv+WEvdOnEKcrtav3AKj1eX4zJrV
leEoUgtUAzL/1vt5qs0iS8w8li0W2TJM3unQ9Uhn7/eCkJZBb4kQSpsuM/rqeuc/
NRQxsuYAjxbV1GgJgeyClkJ0qCSRaGI+x8i9SLyuPgUUY260I+DY3Dan1PjQLRBS
xV4YjseEBObXxLmurR9EJCGd6SpGdorLR99z+F2DP9NJsGIapHKmD+nIBdZ/Uiz5
WrfNWcjLWQ6sB51TOsD55l1lWXPjAJtq4L8VnjeL1agNtKcKkviKFgkUarBRhfYV
wpl5RC86zzXc7JxJQj0dyWPWFQkXw7Kr2rwQ09w1bCtc45Yq5JKXm4ErND3ZemHs
zWPfZXSKwIH26DdXiGJNKqvkCGZDI6vivBqB+Qeb9FQN299Uu4SQQ9QZFcWNVe77
4+OmVV+vuVlEUanFCtdpnNhhsRsxrcsbrR3c14WYSH9sxKPzC93fI6mM9q8io4C6
3+soR7ngGdXDYW08sO8/A/k2+KxZaQ0UZWuMfhWHuKZmKqcOscvpluY0Uq+lWYEj
6PNBK7kQUypO19d6n7tka7XsU8cHRQyKvEubZcgZRDj9sJbOm9464i6yCP9zI6Ge
eqBCyy2rCwkkI8YeW1BCIv7YJjUNkxPN7XkjgQUJIY+kO79Ir0WVIZsl4pjyw4Pg
46r/xkpZvfNLKf4HoLxzRMjS1KmxhfnZ/IIakYJ91FEPhsqUK/e3tAVUWKZgMISl
/uvLA9Mz6XR5i+nQldmj+xQ4vmcHCvgNmkAHwGOmqapx+qxLWGohvXNxAZJHsPvT
KE4aJlJ6q3Ou6iJj+Q5BxUIJ5Jiv6iXpwdNNI9fxzqgp4gUlGv2hZrpsmxiE4QHV
cxv3j8O11zfdTmOdUQi6XTfiMltK0VDAIbHOkbQEMorxAF6I+P2g140FIUum87GU
cRcuFS4n837Bb4r9cfXOPqN4xHIfMISWVRyT7PymGOLErTb5scgMlvjPYKIkyS0s
dviTnsY2AUBStCCEO3a8NHAhIvaEvKTkPnoiMqScm6jWjT4nK44G+ehsLx6B9YX/
PqzwJYMvT+Z5VVGAahYfvtGtoShKHc5KUyjFK+rGwjqWkFACrQbj8doPqh0j/LeY
Ih5TirgAKnqnLdKOU5ZPE/83ySm+OtOx6lfWBDRCLUZ/kNaboRZrJUcH3McmFVH2
Q1ChFmsTHWUzN5SI7UrkPNk/iOZpQH8zDTIWlqeEx6wYx6YepaIx2Q8122E3XCdA
RLBSnSKgT7OdDSf34Ifq1M+B59FzBj1XPwt0A8yrerzZ4PtQn4EHYiJ5RAFsG/Cj
3lNt7vJuZ27zQFB7d5kKd40+zLsrWmaa3vIxEuoniHy3X77DBAVCYBCpaYeckbX3
AKQ725rB8VT/i5SFOpdigEeKMOrZY3DFz8f9sM/b2S0ErP+V1QZ5l0VavUN8Tlq8
gfH4xL3aQtsVlFaZxBe4Lyvpc7/CA1N8qdCtMs/EvasQF8Ceor6nv8ozb/bA443/
HQFGqcS9BTPXlvIbaTczskeMVsDYW6qhHZh7AcL/4rYWshZ/xi5jU2my/uQ1U3KW
T4qprmhZ9ka5Dq7HdwwU+3nJHRVpPxZcJ4JTaBR1iOIaJqiUZzwxfVvV6AU2c4AQ
112DD5OQWVyuXcWwW3Qaz4vHIa39laYtv/qmgAr0UmDx18jRF7OJSm+5txu+xN1N
TcFezM2wHjntpUdxNG34sOIqWgsTNk6ag3v3elAuAJxPlhcmKGk5dIg/2Eai8kUD
soDKTId1nJEb1iPfwZvcpNbG3vWjGOJZvbUOS32wLAacKPUk7hR3+tDRrCFwijOx
uKEiKnPExEoK0ufkLC3uQX2FrIjrwKqKWmZslrsOF+YnsK8nqHKJpnMqjM3m8VZ5
LF+4+rVQqQSlhVYRWovReLzMYQZX2KJamtr8k86bu9jd3IvcGx6+xxkYUPMuFiT6
7Mu5feQgpTRDonF7WcY4bLSgH6NP6WX0dBI4SPM4LFLADqxLwpA2s49sY9t7RNxC
QTgL1xEaT9dhnFcQ656vwHzZDm6txvpOaUyvUrUKv3KtzzHWnnF+1glaZV077PTo
9eGBIJ2gI308v6I/ZbBzmlN7+YwFmbQP0bWAxJJPHs68syUOhFxmu8Uf+xlXodXb
ctQGrsmje2Xb73m46dR3upT9Xq5rB+cfnVERXD+FXfb2bELI+m/1jdyKJv3cMuww
ArOU20Sdh/gylhfjApDxV3eiz9A5Kjpr1KctMBUEELIRPs7eMivwGTLpP9DhWY4r
ZhbgYHVuhPXAUylgYTTUQk2M5LZBm0Uy42nojcTz9NlEdOuEOBqxhQUNKYB/Y677
KTksIlb/ib5TgrwilunABzfw5UzykhmPT7KZDo4zMY8SYMhFUt5ugPajksXy3k4O
XEmGiU4l03g1F9kzja/DK//tHnyw6kxplNpUS/fUoapOU2MK8bYSj7REy6680bCc
tpBTRwLGDKKHGqcFrPC3EhRyFhCMH9WjpsBBBtJ7Jgbs4gTTpjzjZ2EA+D3RkeyO
gYrF6sFG880Gi/EJNH5K8SQfuHW+Bqemt36KBZz8eSpAof5g3E5H3sbINTZakRby
8df6RkL459D3pIwrWvzkYvGmAv2niu8alc4aRzxleAzhukTDrUNJkTnF4L2ogMg7
+7u77+hzFmls9lLP+NyhtVcY8xbsAQtXcj/2eDKI8qQXoJ3BMTo85kUC/FYl8YkT
YJ2B1I2NHO5KthiszZXazZUMcHuxEthYRP2wzelcgpKQ95TQywzfSE2j2KZuXZ1V
gzqBZJPe1i7MUq8mnDchHzLIc66tQ3lnkrx1UrOoEosb53CU4WI45JB5sA9m/uwA
nTYTCA5LycPT+B4ogWuSCfFTnIklTsfMynpj2EK5YKanFbrdBKGUOYnqy6E/wAnI
PqKpv5E7QhOV9DDToLqslmLfKcYxvdmT07YYMA+B4CJLO688H0ISmsRGdlrSjpv3
PhWFHf/zUzpSdX55ASg7DVAyRTgD7SOys+fm8JLFsd/Cihk+CX/oOWYnkgLzNRIa
QzZ7HpBP0LIh4xIrEh+fa/H3YQg1RVcaXnWhaxldsOlUR8ko3h8FbR1EwlyhF1Ra
gu55xQMkkEo3rEzwWCl8dUgMhOl8z+Tzu/10ROemzUh86MPIcl7qUuNvTtQ+mv+J
+rdWVaZ7/iJ9FZZm++uxHk8QMVm/hUvDAjTlidCM/rt/KH5ieHwCuzw0BuzAZKnG
Xbh3GWeguWOSFrDulvBAYHfVXJaYZS/80OMwTcNKhudbUe2GTEx0h2/XHtHBzT87
EdPNGRWX1n5cijC2KBK1N32qlHyF8OcL8VSNxWNuG8e1FbOVl6H8MeNFPk7W65GP
d0DXyFreRqiHySSGGk/oQ+XNZOuJF0NI3OFHW9eqxNkuRFvQevEyn5wwjkxZzkPv
euIxmWKLNltDbqJ2ZMimJWp/BXTa+1MSsKQyikE7fO2mY0ah0f5jFGxuAxyEmMzY
5bmLTA33FE9VUOexihHVs972bX3A+wpuZv9MDMFxlcx6LqaZRuZYn4F6AHCyr4fN
+DQfIGHZyr91JhKcAQI7hxWzFDvyTX/3BCHOGilPmKpAB27VInwJkY0PrChhMw6j
7aWMSHx3zI/yCeZWSnFjzZoyzkZAE1Aat7wRaEvq03FoLq50UuSbLpohxHCzL5tH
iegkdbcdwmR+z1c9pXpQeQA0KgaCgZi0XZee/6c/x+JBivgsTB6Dwal7vVDzED63
zUaOa44zlGR0izg/fqPzrdOqeUMYs1rgqNXrFkTKKYhxZBnqSNanJB4YYOQfQlRg
XBp+MxaVKQc3hgpmhD92hAJbrhx9g1x2y+BNrYVS54G5spGR5bJ2DHPgleNIfxr8
72+s3zUu0GaLTzNvZcuzGqWiIUyNPwv9ie7B6EbpCbUIDSSuxpTG5sVVsB2xIbMt
OqM1XXeKHNB1uBqNaV5+X9CPScSXofehdcI7l6GXM3x9eD2JrUvDs2qWc3BepUUG
o1Pw0DfS4D34KUk6Z9Mr0+I33p7hw9L0xaolmX56mngCPKdcN8l3FGQe3TlJ5fjn
uuaWcwx61k6WX8B77X7WvA3pCxda0ZgqyO7VRg2BoN1B9VNy9OM9SP+qBsNkWFee
AZl5y8bK31oa5yx6fsIxZWi/sWjYZH3Rg8kWRoKmaHL0+ue3jWiWpLToIx3epMvA
Os3ZH8yhYm6xxkliKhPRJ13HZ+JfWxLtt1v+MmCz8nIkXsMG6VTiEqgONdW/PpW7
RPoKvRM3pfPN2BHBLZYF6IXybI964sFCpdv826Qf+LdAS3JPKfwXo1+HTiTyntY2
3dlcKmxRZa80CegdhqnibEaAFrKtpwUS6HYx6pL9g6zRDJ4EKK1fXVVLtQlHyAN0
NxEnQTiivs6SOEr36nwtQK5p7ka38JGWF17zT2SAxVdfW457o/qLAuzdp/wgyAdD
46rTlERC3imZ+KY3sjOQo4PQVCYhyjfQLUkdQ8Cpy/dV2X+pxvXZsiXox/xwFvUS
pS98cXH0yNeGWM7bUoqQUqe1TJfG0nmGz43cjV07yLvFHjWK9dLP3tJvSZbu00yQ
1T/4WTfTaslosyZKMCQwOilq/osVwMaTZRewHQIDDXZ6MLsiF/mFvIsryNjFzt2C
Y3SqQczm/QUI8tmLt2YPaTmvD9Co0l7+KQ1oFAZih9xeHb9VFPfue52+PP1oycUY
H6CLngS8yLrLAbHP48vCEIw+/iZfP3LtQWkwfTwSr80ELfsozE6x3FOUzO5+pm8q
X1M1Id0LaM0Jue6p0amspOfnpgyVXJDZdhaB1Ou7E8g0zBVl0OsW5PYowDFZwcad
kKfsvV8w5tLvk0mc5X0hjBXBLPfNKIaAmwwvI6P/LBzBRXWOBu/3gntOstRY7Sam
KSTWOgokvhejxR/Bd4Ua92GrJ7jaYNYtVLMpJyEBycSKmvgGgi4YF/51zFHa91b+
XXCykkpMaTjj5+HdqhijQfNvTdiVp9Q7tRmC1L5dF5kj6Sz4ZMB2mZ6srvYdCGIA
RxiBVlntClb6Mg7pc8BruzFj7GOZGMbwgtqWAzjZF0XydZ7G2vvJR0EnCcVE27xV
l6lggM5hk+mGXI8O3d91WaTVfUvXAZy9yo7X1ok3cyIY+aPkBP6C4Hqeqg6iSlZJ
F6OHa3W4LmCXzAfDRGdH6k71WFve9xVzIp0DwZyESCEfVCtMM6sobIlVuTvo/zjh
mWuJrDUuwGi4R4zq1gBBytrZHrRTLeKb/cd1+QrYyafqqJtOnh7k09h0VZ8mV1k1
NeMWfw3jnXLJwqq1m4K4hpzx7YeHFwJdkrIsYvzx492DnH76VjX5IAOe0R3iQrAW
f9MmBFcf8Sa6a+bBAsrmzbSeQPKr36iHT4vAWGC6U311n2YH/+l3z7gYqhwKivWw
d2wQUI+MlpFMxu/mmNZuw9wAcs7sjgUgiM1m22a05ay0nGrMMSNHfCCQM9N1CeTg
DbwfdxUYLp65M70TV7BGS73mjdVnJ/bIAA6DpcXJcCFXYyyXqPdJ48j6+DhUnnZG
v4pqCnvosqewg2ncT6ySHrnTkczzuvoW6ZdWL4RdE4sAaMku0gia14atXbD/a8bS
LzN2Mv6oSN2Ao5nlrDLnzkq8mrdj0U3pG369jHxLuQ1EAny1lOprl+3XDgN7/zeV
8U7W7qu381KlUoKZ0A9XAU8nZ7jTI6cCVlXo26Of3h/G8LS5RAQl1quWPA6VjLBF
rNY66bc7pMe8ZS+wWCi0I4KUzv/sNmkLmZdsrYD6BbkxwVDjTG8ijUhyTPewChgw
wuQmHEa+qqW6Fo8wJDLo+aIW6Uz5Drw5Uz2cLiR36eUcteb0ynnSbKYr3K3LS2r9
EXSxWfefTxR1IAqkYou4S7E5aTtNAB13bsHM1I5qjCVncdQHM21cD5E9JpxUC5nh
RuxdL9wC6zg5AQVqwwvanXd1KbD5JfKgpLUNkKeckxq7gdEfg6vftUjw9o/b7JK2
h4nnVuUlNxuuiPtQ1wAzV3u1l6hc0vXpeIKefkDvxoF/NDLKV4scCNmnk59kuCG7
uMX/g+0r4oPbogJe1+MlWWPjxbEsep4c6OpJ2Yz2y2Uta+JnscsC/CpxJi/z7S37
IrUItvH6lZejDu3lTSwaX7SlSojecldkvOOAAjNA8wJnmCnf5O+Yd+k8Y6dBi3EA
YXnSyVpMB7bNKNuJadaw/9S4x5Rk5q/F7pO6wO3iuM0z63BMQAzhnlxG9skVl6yE
c49MKvfsaA8DAu9sERnyIp7Z5FR+A7YIc+kqYR5IMoFbyhlPDoSrBu7iSCIJcDc3
zDcF19R7TPaOTJKMap3t2/TGLby8XXUeXpY80wPXkWM3xxMgRmtoC3nYTYe/jki0
VvCbqrY6N/HHkc4nr1O2cEfWeJnnRoJuzcKTX+mH8qyShqBsTwOoVGdiShra5o+J
bebX7MpFRWjM8EVIssMwEvCJZMYofe+NfnU+JVdsAA3NJtm/S44zvyUpIYWXPRxV
5D5nxA/w1t0kbeZ1iBEmEnm+c3Tkgfctz+E7RM2sbgTJ/4Krmuve2HUPXal5prck
bUUx3wRObvnctWfLImPHtKcgvIX8IM6ouhoN4mMThhFYPYA6xlLRfSE5uE60KGN3
bcCmtKzFOOeBPFL7gRgzMZdetCZFGmav9MuK+6/uyI2nQAvh/8AIvow8SL1Rg3Um
J+gl6FFWJs2h8WzkQ7cKq82Hg6ZE0/CbhHqMq4GpF30UjVeXfUqhHkT19Dqj5H5r
XFcss0nJp5SG2rmMN4IZGOosI4OYzIMOBt8kENj8XJPc1NdVylfC/qFP3hxaoDEi
nQxDsmJFfvEtsBvw+IwlpIHZpWMw4k7iFoc5+6ufs3kv/EKpV43uMIyKFHEHnHwI
dZFLCcSu25NnjJPt+bADQnPAE1BmOAJ/DGCCtOY40Na01mhDZ0eweGFI5pVuFxpc
F14eamGpkAuOpHQwjnOLF3AMoszl9NuzZjl70eGR7hmuZ9H6Nz2MgzKOamG2SjIg
kmoYy7sZBygeNF0qDiL0X9+qIHJQdAOahREgJj+cpA9HomVFwEIg2uQ1vAhRA+Qc
FZmNeO166Jgrd1t6nLUTe7ieUNC4DLoa4GnE4R1VMK2kuhpLxf6k+XOEs2hpubEO
4VOiL+OGgFhooqQBlkm1/jSd/WPxC6EHkGznycZ/riol1bwMAgIq3V9q5Dp3RhSy
OB/bxVB9ViJbfc2oSFUmAVQDzwALBtE16DJzKnqgOp1CDTIZWScpU3dk23ha9fQT
CUNOaJ9Mz9DaME3nPkK2/NK8wphMI6cCG3E2hD3eoJX7mQ/w/sWwepTx3aK1FRNa
+GgIKahfDDJC2WKxtF4Ehp3/bl6oCY60PNrp+DxLU19paJp56NrPgep0zJeHzoWX
osp3Wcd3eqcyjpoN2Jh5gmVLKd5MaRdaIHRwvtJCcutC3hR/TEqojyPlG5LGIadw
Fpf6j87OWyviR7qFPYMbkLlah9l1IzEsxqSMVsB9h6Nxk76sgHK3QTzUQ2RpuQRG
BJ40QpwTwRWoT0OsKnPNwiFZJJWStZUYAUjkqSv0jOmd4lWPapYWuOuUb3ocr/qw
D63NpT02U879ICh8ZqODg6T8nKKghbqWUnVaE+doMJwcqi4yvALOfe2f9uv9Ckvv
i5naR5eaFFyQN2NBsOmf3qVpUE0FJpiKMuQOR0no6cxSshAavV//JTG3YISlGM3V
V4cXTcE5NHkUlNIg/jU8hg4cKS1H0HE0UI2WkqSwXToj4DQDoySEeSuA68pzgh3+
1Th5qLQkdrfzPXDzSVeBczzCWxLMIJhrsBbH3D8xgFN0KIrEZ57AQfHDdleonMwW
U0PwnX+AffVBpAF/YhD2Hrl5kn6CVUz1AX8bTgmtvZMoFBs+CmsN0rjk11koqSSH
gNxtztra3GKBhPIzE/wR0uHkYln7XjQp8CUeFhDEr9RVcxn0mCJH924sMcx76jt+
x6Q4PL/ht+/nXMLuWouZ50UlGs9T4IuUe6S1T0cgdWW4DV7ZXZZi49ZStaJO5yAJ
bjAQzniFDrkvLuYBp0r22IUys4OE6YY/n6Y4qThUWSbK22lUELX8t577IyGKhqk+
YenzP42ax2o27i+iVfpQUdaerH16NeEQxMP3BGOh4nAKLD0z/M4kHYYBkWWZyU5K
c8A99Q8H7Np7ahopGmdCxN5uzgPc6/GkKTxSWoAHdyECJr/SbF+RzR95Vs5Pmo8+
zdbHqzw+UP6NYXZu0ggDQJRTSB0u2Vilm3uypLSAnRWdJUu1SmTDcVEmElkBzu1l
alk2y4+dMkjIUn0IzUD+GgtfAvVYzVzQBIVTsP8xNl2PjjDX93g8YqTGgG7g2wQM
Op4hZC9/tpK+ydXxqyqXiLBOHtmVnrKUzXrSFojgvj0S7Udz/KhdyLOdi8mhaosc
ixvhVlOAPDhKitb7P8Anx5Y1XoF6JAq3Ly2aTZBm5CHtxrQkYFSXLcpO4lnZfT8S
Yl/WivrP8pnJtNWltCY1D1HrXFetQJWunYgS0j6zVdtmFSaBmpdJJNZxYDbxwvSA
lp9HyVi4bwnPDm2Y40JhDEN4vcddBx9L+KxR3qb2s2uXBYWID6Kzp+lnbA9PJtQ2
EeVMBbBkW4aV6h2ChONKvFfGyd691c2Zn346LHXGvw0P68Z/lIrRpJnhGqFqnFjR
Ryly/1X7PrQCzAEqaTbGkwc8Dz5Su2Tbw+MHUb+AyhTMfEXIRAV6JrAAWdi9Td39
zUjO3MHKnw8pEZmOb4N74gft0GbtzKOiQcIIP/SbT6F4axnpovb4J9+WVkij+E5m
zJECJ7cR510I49h/WvrndoIpz62QS1EMUXW7JP2In9wrRmsJy91hM1y3rnXIy4Ho
+NOj8tscmRiFuOIwbp5Fg0kQW8/S/UWwzm1RnYP6DsgppG+TTvMMO1Pdau0e+a8a
e/Z3Pdj2c5W9nz3PfssxMdBrAbrhxwlKPoI0ZekznGG5b66nxjmWevG9ZtKqWOwv
grv94dZKkGtU6J0/a3A3zx5dlt4sFt+TUsBEKCd6j0skdErF5h1Dp0oufExZzi5n
xRkUXfH6VMhDWuBelLYca3zx0eB/nbAYhBXW597QmCRhFgbQrJiLbK3ZUfQ1oB9p
qCJYo3faIAd6m31XNQS+t07vc4bWyKx7MghmmevSeCG7F6BHsoTLdMTC+OjXm76Y
9nDY82ItNKA8n84uyH5NYuvOJivOxAVR3oR9TlrXlwI/dJcfYJPh4K1p8nEJFMM/
gtCcuofxyNAVCKF9AqLpXcU8WBzzE9AI5M8QpUdmWfgrr7e9Kvk/RW9KzupCUO3a
PT+b5ea+07VfVjTm/+amJzS9Ov9QYXR9G/kw+Pg6FON9lXSpaTieMqGoztsvwoJl
C9jUyZaP6KJNv8ZA/2mlH8tLdcYII1kAFPg/ipcNNi0U6aH1BunCy0u9OZZJYlqm
FR8WHuYGYg2h8FwegVfDSJloEwThoQV50/nOWac4zfCztBl0YTXUOGT5s9tDNoIp
Jfz47NLhyvRUy3LGJpb9niktTDbbzqLQm5z6PtOiKuSBUiknj0ANOX9jUPW8Y8NK
TROfHSDi57NVFdTXKQR3fqfjKvfw3gJxHSbM0lrpHw4shEnCLToUTnTsrQAvIbp9
kzZiXwJL/BxqlikxSa8xU3w494pcT1yC8Hf1H/SHx+opC+SFN25IenFukpQ/vvj5
x7RB+HqzZPz7hSmSRndzIHyGUszAitWx/1WA0YZHuw9MUOYN3I5Y4ebgJoZcH22g
sGFbWFfoBeC99sRR7eDWTAnrQM+6g6heNicCGS5mP19OxN5tgFf2hTNPuRafMJoY
Spnpmvfnf0aofNfJIylvePhXzUTtQ3QvEcNKH3ymj/ZTN+fuV8qAwAVCRuCP4laI
WjS9c6MzLEKegUSjA/y3aokH2VglDbqyxsLwj0/QUmgjMTr8TPO6djONAZXMoLnW
bSWDKUVGYCAZSKru+hQNzb3JoCUU5a2jG44I1E3k/TMcZ5KkR8KXGFLh+Mo1ssgz
DqBb4XYuCbZovsGFJ0ufF7sYVtUEw7pXh+/tWg/85kuRMtha2yRYsSeAF0jr/Ur2
AlRn4LeEjE8DMfS3cbF1vF+RGRpO+tBv9E/xTb5ZQ64Si49wx82Lp9OVhm0PqIOu
8v5DXFd9heNMH/zRlkdaBLpFvik+KScD2KPgl48XJwiOWGwS1o5AM1x35rIzWfaS
HNdAwZsHer9JKHtL/JbXBmWujZPhRtlO+Krht4sWK5CqwvyYhdQqKhl6hvXrJ3aw
7qzXjGNMyYkznxxD3v3PkVhMSSHHlrdfYx316nGB6Tb8GkTB4SCy9Ib6C1ObXkTk
AwOsGyyIUZUPPA5YqNT1SPBZyeEbCiDt6PRdpOVGz3Syw49VUBK8EeOoCX1NikMk
LS9AVw0oEcTv0TLLrZ1fBc+Qgg2fmH47daZB8tpVaN1bHjG/nVxKK9OkJR9e3575
rhaM4XzmI/VCaztTt105NZOb+zNleWU3dyvqUmyuIhHvoWVHk3D9LZNJA+MMRbcV
zsvweCkhefuEIeUlO+Azv7+9lsYnlU03v4wW3Jw/9sSzmGMwPI1snbpW1Kbop/6b
B/97MUZUI2H6L12A6fi21A2j6JNQfoE2jrh70U5dMuPiErJ9c2jj0qJC/LztOpYq
2RSwu7Ro4XQgbwlh6EbKfdOCmCX1lR30/4bVp8ZValTYKwoWFy83LKk93CxWtC3x
4q4dccVWFaSblWZPQK7vkM/8M0fOz9roHpExZRYhtVtMuwqPxJttLy3AipYTBUDr
nbzlIdIxEhWT+W5lI8zJeK0tCor6ch+Mty4xNkBI98F9vXADt23oHMU1YHrvYAr4
1iji4wcEkbWyYz8UY9kd7c9X9PfEr3PRfzNELfL0f7FquiL7T6u5niReYsDc0UF7
PfDv13LemXw9mhLyt9Afx1vmiWu4SVeUhjRiwMgcJRrrYun4z8sD6jA0NNAJc7L5
9p1jl/bWUT/Q+53evz9Fcq3Qu5euIOWLKJFfbVqEkR6jMF3BAvJS9W3pzWfFYOtX
kVf/2hWCCPtwYNWrKnL13mJ5iIuXTjz8faDNuqq28zvMMmORuB5b/XxX+Tv9ioLV
ZUKD/rI/oWU2zd3Q9YI/R3S5743WebBp2q89SPO9MY851vCrmZsLKOvz4ZlaPt7o
NPWT2Z3Skb8pwvWWmQ+q6FECSixfXvg31IrM45PDr2e+lsO60ErZjqeaq6Gp2fE2
9YxWuoegoSuhy9SnzGW1N8xtKbBdSbeLztjiBUBiRL1PR/8x77V+VhRlUN4IaduF
KyCB+RLuS7nNDzc+9AqkoLMiEmbOBDtl3REBHBd9ISysH7GbGblodLVTbuf9Fhhk
CbM3cdwcZQsCJ5tO4OJspLFnPDvAc57tjgtY7+RaeEGOMmTUGnSOv6RosmlLin81
mSHei3584uW+kUOPhtBHkA9XpBYewsNNqJsfDvHxxTiTw9GHItVIcMTVRkcAhqBg
on95ltv0WT2C+yDTkiT5voiFxFRKsdWO326hHYFjtk3dSlUyiwJphhQEWeV5mVlX
nAIuJ1MjeSyR0sH4HOffhSf3MtpZl29vRhDvhbKptnXVEf1rgWRTahfvdBAxr8XH
WuIcJ3fPvlE4f/i6/syMums3tOCrsc9Fc+HkCGDvdnNAzGytfQ0hS5W2/5bVe4tP
pjHY0VP94EZk2hXcT3qExMsOL44w43LbsOSq61qWEVJ5f5OtAnSkPhG+tELzz+8p
0EqtvrebYuE7Eu7cQUiSpJZTozqQgmldUjkOUHOQN1ViTexPUEaVBhSrWUr2awev
GPrlfFl2iTrVT4ye20FFyAkWr2EngL4MebaNlgv2wOvSa6UX6csOCYtLVyRt8XVZ
qYo3witmlQYnIEFHg7UE0xk32ns5ZajJCU4wv8KjJ+WtDI3TcTq1IzgNSsXAdRb0
c5xOZlCC8fDKolFSzQ2Jd4JFx0fAEK5cveTrJRl019TBM7/iaJuEmQXADcIhfD0I
79Xko1qnkn4OZrk15/ddG3BvfZ27etbKVqZeq2WomANZb2SO9zkpdyu9KeLeJ2zc
lblSv2IwRpohoIoWOj8ydjiq/P5sX8psboZZCDW3dhYG1d9qApoxA2hwXtHaYK5r
WoQPEpowgbZG+cFACmJkOWYEV/Tdxg8L0bRwit0kfGOfXMXkng6QRhFKDWPKOn5R
Rzv5bkrVSvvdeLZ4iN6Pbk373N8KmyVtZ75sUGRpPXigdPQ1UpU3IcrDHcf2Zv2C
JvmI2/FN/CfrzRNHoCsCvhFVMwpQ9+UecwrmFos9T4TGzG0HmyfMoMgGbEXow6cA
TaCohyO6x6rwKvr8ot/8ax9HEud+MPWnQISozP8WwM/vVZ2XkkiFyvfhxQ2iwXmL
pLrWMiuZpmMbUwoPgKjRZ4Roa8eul5ke9wQiGIBVt2oQ4S3DB7GI/mRKcLx0pI0V
MqTQ1o1Sjt6HqBpJT8r67sDYDf1Jk0z1Gatxkm1ek0WfkoQ00nf1d8xtKsueJS84
W37H8IXQ/ImLLvxDw7P2v3log5SL75v5wyWTkob01LiTNBQ9KyefW+qZrHWzVvYE
2dCRRH7RUy70J1nGzsBrr+QA6d8FWNp6QFJqA9rC+iLFXN+qmcWS/6j2ljhjgz82
KrQ/k8oLTR0lOs32Fbxbx1EWezRR/CimuUO5ohga6LWxNtP6qUm3FRvSha22Q9TY
A2wPvRZBxXvlf8FQYQXs7O4F1Qun3oJf9DIOGpFkDE2ZYHl29Wcx1UhsmnJEaDuw
g06qJPNNnHVims+kwuksQdVYqaOlt2TMW3A4+5r0oyIGkZnq+RGXm5C483EuSEf3
vp+vMseLjrYpSnUe6OMxYOUDttMhwUH0KvEHe08QaS+0gzUW/V2uXZclMe8T6lx0
xMUnbWDvSpA/cAts8lm/x5TiVN6+9Kv5TjcKuoYCj8o4D2DXSPYH+QJelcaypZkt
lbXlOTYV2l1e+6eaJLo4c46CW+1jZDKxKTMZptVmLN8NCG9W55qyKvnJcTuquaVD
tUnIR4opiumgpC8vnCie7QknzgpvbA+0B6Nt/2hmr9i5Q7EyvoFFgI858VzeiaHM
cjTIClP/5qJ+jGv4B89kDNyQV43txui/2IK9N77mDzF6XZTatFA0YH6zbUWZF+kb
hDG4Nd7meK5P4zzVdD2YlkbDZpRDK6KIoZD1q0/B1ncHn1Ca8zHzWE7xYhgV2SCO
zqvi+6XldPhan6e9azBbi/TLvrWbTNkuOSzGNyeiVWsydOO5pnIU7HnjnZnqqv5V
9RF5dJxKTkrUWoKJjLNywb+WfqId2oK+GDnMQ7XamA6sZAcYS8HCsar6122CMF4I
/9q9m2ZvZOFl3oocTD8sQaa1+vlOzRA8WGkzWrKHogl8+a8uRs8OweIckMKv8Skw
U8CwdHywY7t1ogJcNgyEY17b0JkTOWHyhIVh/TxtF2AxK2FnAQ5jmUsw138Xp7nK
cDap/KlsZYVmJU3+BZNpzL598igSWzW9+Vw/16xW2YtBL+FGF2j9/+gqJH7e4rqC
xka4roy/knwDjcbI28iilSitNXSIxGGBVcjqjmPsXe1OGxDS1Lyy6xY/r4sY2Z1q
XYbkgugjtU9ktAXshK7GaWOsV9LL7Nv8yYj4F1eFOofIIETtYe8zq1wpQVzLDpwp
nQxwTja0XBXQwjMwSqz4I9/agQH2R1kbo1/yISZ6YezkSbah1OXRL/7HJMBC35vF
X5N7IW3ZNQbQKHB5Dm0NgS+bC19wuZfgabOS9wf+lUwIIaW2Tipy9hFxy5wXGufi
eAuJD5VEJ1aWRYSSxEuZKOsj0pGzfNbkhgPL6P/ZT4S8EdZ9K1AZ6JakBWjIYnea
nBQu9rQNpu9dzPrIClAb3wS9y39oQwmjPjV0VYCcb1H1De8DPZ1uCJFV8Z57T/1B
DR2Gk89t5xk9x3Fbh+nQVVcQ5sVTbp5EOvD4Zo+1k0XqE56ORTCWvOzCe3uKRlV6
VUQSDeGjSOdfQcZL5zS/OkOjOf5JyVBdl1fo3BpPIopfX9Rn4U0ARk2lyQ8wlybr
iFLxGMhsZTWsiSOyJlHMvTXgUfUl4333UKwb/r5Bk13dij5msTq5YcVljK9RxYJy
LEFB3R0nIXdRg8ngovOCk6okEnIF/W8k0PEtUSLHtRo0K/XfTDWSMSzaXUaJqOwH
jE6lD20mPu3EB8sPL1j5ouYk74H4RcJFN5raspDLZqTE/vwVE2Xi5hktwXekxXW7
VCtiSGvZN638EHY2SJ6bgcWSKiz5ejXoPMoEELAIzljb3+Hb2RItuScdsLAGQxwd
c4+j60UW7mlWR1t/12b084Jzdiyu9OCYUIN3TOtPGTQ3AAb5btdDkZ1YI44VzNE8
PM887D4089gxrWlh2cKsC9nI686V1r8Vofi37Sp1ArSTTLmnJxq1599Wb6fFtRxO
IYsV2fuAxGGjAArlmoR6spY7AS5Tzv9OgsTB1XdJqXw3N6tLyjefAWoNel4HKAOy
oZ6GLxFx5MIztO3GIIPi4/MqZq1p989m9WRJS2ubU6H5dSpEZOk1zWucDqoCw1ST
A9Zyyjqtm9JmHRtTMXZAoPvAknjkJJpBJc5nyXv61L1bDkzD0jGVYYerLjr2hrkj
Qtk3/qhu//1XgCK3FUUnqWOMTxWsHqareJhl25c/DeFJufOlgLjY24Xs6OaEenkq
9bmNAjn8agm2htN8WP5LmX/WtoHumRVUgjNreIZU+TO/mjDt0Q/9xWYN24rZnhEW
D/ImmIR5CJ+eVPjlVgEA2iM8zcb7QMAw9lp8bPdILwpfMisrd5ueGySFZMvKMqN3
B8irBD/2/w7mvQVA69rXVj5+uobtHfCmXYdNgRfeDEhHo8wBMTiPk/y3nxoK6XCq
mWS9n8rybcPAL7noSOhmTx1vWEU4bjylh2l0rzqyThch6KyJADutrp3taS1F94ZC
3zgbJJOHxLw+cowMLDLOvN7wigkPQJpaHKFWPpky3/DAouz45kF7JokgYccraBhd
/D47bl1NgFb5MR73Wc7A7I4wh6qD9BT3yXNAbPo0e2txnMtV4Yy11aCHNCtRB5br
88PBNT2XVMxEYZT5uI4sV5kYosH1dcI146WrnLCDNbI3bWxtkj1Obz5D8f0aT2Gd
s83+3i0jL32V+TzvLh6dHBr1AMgAo1lsCg6x0Xi4CvQ2YDXjG5yiMiVf+O9ZyowY
Ku7HHS++Dhlv8ct0wdJ0pqXSQsnJjPkDDhG7isSkUg9gWfcf9qcEtThMs3nBND2S
bfScpCFPfpkJQ0CJzs779N/PJctpPt48GQKGKRGNjDnNdUW2jyhGp5E2M2f3mgKe
2nJX9G7os7A6fgC+2G/7+oTcZTtYUrB9igAVvrprvhbwEA8Sc9HF6CJrK+9yh0bW
9skcgsDP0RMCrUfh7WoNGoaw8VYHwnqar2eOI4Bkj0PNHcFoCcyb3APHMMdE2pmW
VLqkL+TbILLQnbD0Xl++Un0NzV0CDB8MpZOtAvVAoTlEiEMNzOZR+cyozVBsDw5q
r2mHVWVVc6b0qK5yOrlM4y5MFGjJVTHmtmO99zJJQcx90FuCuA3aXonpj4YtVIQh
sVV+qsGgGLN8Y4tEP3CUxR0qAiOhYKqUcH+Je2Zx4y/8Q9s4CK3PDyMQp7m5JXeY
5jrbEBzI+XIJA3IGLakLWo3ppLm+DoWUSaPJbdDliInIhzhfHfDm9DlaD7J2CGI+
aSisITNhZIHM/SPbcnWiRSz/iW3LX8FOFe4UJaEZtv3faphKrwrxZ50Enrz373RP
5548PnfgXCDydYu8pYctMRu+4u4D0PDjmiSQ6HOOcECRUIpTpA1s0899dmsLHpUP
1t5igr24XEJN+QrEr3t1nMTUEX8dEqNj1GWm1xZDu45WTmTAKbSh3GWnG0QkBXO8
dBgUUOKAlJePOjTmUxwIakDI59fm9kIfHt6fzCMKrnU5AYRzm/CQgXonisW0nwLB
Ff0zL06HNuQ+9O7ze626Tvw80zIXtVh6XNMOsXSzNqUvJd9axGxLD6yA/wz/ktnF
kEULQMxWw8bppTwuqy5DvEEWjuNLxx9YbnpHI/CHCPpKKp/YTkGgJA4u4OH9kEWH
XQSn1OhUj8BUA6fHBgY5qeGXKwsiK6wVKyLF8dJWD2EBKwuFYrnJ56Fr8bgNOgSQ
CmKrbORBkR2NsDNO7l0otXyudg7r2ef43okMD9CJMkgfTk7SRgIzTGMLlZNQ0Glr
SwhB78rqJD1b606yQj1mgMjy6zG+JMhhH0saYjfV3N2alOqt2mJghPDogSjq1ug1
x+dmYrldGjKVTJZ1rqVMz14uRF78cCO5g+UC1ceOKqwW+TAG1HwYuXTdNI2lNO/M
sN9ghUGwaHBuuS7F+JNTw+o8MMGhRoraleFelG5msUQ+eXfhNrSoMVESPGqHYeJa
XGvX4qyeFwR6JQa9cOzERPWW+FJd8B1+8lUZguYSf5/M9xiqGtUN/xv0ElDd/K8K
KWPdKGzqwmqGL9x6o0amJz2Z8t3YI9BTvDs4fXXdqq0UvjU9H1RG5SPb18NMy94j
H7Z/DvSTc6+s9Xi5nMEvJFZKwAm1qXa0G0eGU5WiJBMRquASPg8pb+of2F4755OD
Jb+o0Zpkifyj4ssQ8vOwGE9EMkaCbT40ahVmby8UAZ0OHZ6Y+RtlWosEUI7jbiZ7
qi/GhW235AXOr6/jruSapSGCnE4Q1QCaNH4hn+5WW9EjuOrBeC7Aul5k7eWSwRw7
8xd0FM6PfsaXo2Tho3G+pIy9801WZIZHeN44ts3llW5KapEDHqQXuqjfpejm6qBP
Z658gvPnqbPBniB7S8bTmN9zKUvuobXlYTyEU2NAXNp2G+PChEqDpA845W52JLVt
85TAoQ1KKFuLVzjXAsLaFHqJN8xz2qWc/ILOdNvoU8uILYKQIriqG2APlkA3UXOo
kMpMHeEuKdju14NcED7hiK3kyl9yXwWZI/4WwKbkna2cG5fjsJ2fvTOzf3F2WsH8
fidPtaPT2QU4f4ognTIFIzcq95x/F+PsSXMWu5cGsRWWRgMpIKM7eRctOty/nCey
PRs/XPyIG7o2A+q5DrozRw3LDZO1O45p1Won7jubtS7/WD8wPC3/VbbRgNA04KU6
qVIrw9bgiyuf2xSXC08bamfGoDKJ+HVP0dJ0PaalHmLVIQhQRMMl0IpZKnw2ghNO
WPiZDxEAGsPHmuHC88d1fjRlRJA8pu9kzH+djw8+9bF523tzf7TyWs/q2LXhbg84
gkYGjQKxOrC57FIrPcOFyIFcshkOGH592TtVzTVKIjoW2joqjQiYuSiQS7H+Maig
CNnzjxZu+TsEUEouujG7rnbi7qBtG1uVBlz+LF63j7CEimjUcoAMla7xCMOwIq2w
NjvxJA6h8ivB+wVZ1lVDCgfGv5v4DEBVxG5CW0MSqp9AGI3IzlDG8dwwk2vtUaVx
2ZC0osccET4NXz9i7y2cGuqDBqF2GOtSp9AHHf4xvVxReM27GqKF85LtR9L5lpDl
M7VaseTqnDYOGzGx0TUz0VdwTmiW/ExNQ8B6+24y8QPHyezSqfUzp9JK2cZItB9e
Z+Cp5bIEULfWHEBhVJhO6BgrIrLFJhNfhnRV8sUAwk0kHlIlthsTBoyg6N2DL2Al
frHpekeA30HsmV0LA5khJUav5ZlR/1yZmI7YHngn+X6E+uQ/cV4gxTL8z7R4SvAn
RrqvOjdkC/eZEhXtlyxheNd+ELQhoHcAz5nvEDdWkKGlPCg9jHPIZJYesyp+60In
iEeNnRtxmT0IW3TdW4xSJy99CfnSRE+FBEtoCSrSp16gK8fUJB2mgoAaJQYYxGtg
RMzO1t8PavpKFN43e8IUNPjWcO+EckJ2OGtStySo712cXgsY5ut6AWvWFvPdRlQq
6ydYHG7s4Ou5lJbUZCEWEnpU9WEHb//u8bz0AFbOtTSafZSAoOey7BBYBp/wGWtS
Ljb5i5G4EIa9jnr0SlPRPz1zS5QzePNp4UY8mq9sK6pNCjrza2MG0oAu+/fYUtbx
kmHJzMQdXcR3qFp9gDi0qq2zuCqG2r0rpeNRDKuEo/Na4oc5qeY0IgPyktB3je/B
17JnH7fVrUvn4lZljuWdG0xV/deDWNhQkqF2JyKbvGs6AvHzJsHJ0P2S+lp6Fvy4
CGv/t12JpxjJlpJr1GkIrHT5S0Xuqum9afO5Ary1KxOfuXYHkPVKFCTn7s4aZif0
WvYiAR81IB/7vxDHfRRP92Yb+e0/Yh20Ex9lErmiOpS1Fbv4JiLDp3A4gSVQDXzu
QbDKBtMujsXjPQc0padeCJBGKeatdWDEnBGs658K8ol+RcWZH45xVFGYyavubUwU
wnKux7reUDpJTlykeGJ+XnI6ZPcUCNAhPiIsqhUvhBiv36rFcEkBQnhx3VRh+Q0c
FfEAqHkJmMuCvKQM5lXOyAv2Ype3JGopcsc9MSW7WHnD6brBpSDMgkQ4YBXqEISx
h4CVrFIxeDnBhJvoL5BGyIaqjeETLD5qt3Hl9WiM/SGL+wOBZJnvBK3e9Orcg8Sz
7bvqZdclFKlGdq9/qpT0yUiYX1itS6FszrNUy0TCr1shuLtzHSTn04TMgM/KPiQI
M+tkvgaZrIU5dBmvcI23aZuR/fKmsqiDD5QnoZCLidnOjaaX6pYFI5VxO8fNXhpD
bBbr6+aUtIFgKwifReq1Tzpx/4yIq43LhgPAwu2xyOvJuHKigT8M+SF4iqKgT0Qh
pmzy9vpmNVDGy086jGZczayRBsLaXgoUtSiWoiAzMvSKsFwSBD1u5NIdTI3RAe2w
U4cCg0b+fAqVlhFLBUkWLzUYFQbOKbmOmeVX6wzjzFZbROyW3uEPdYtGqMbx2Pld
Mc9tm9MrpSAMqtngtEUGQuRgAOffkUDUZH01Mnwl17h/9HHxdEecYtcs76luEQmI
1Rbd6bASi73o4YQZ+xi/YYmEM5sib3437/kg+ntPId0SrykLgGEI1A5pAZ8/eED2
16qAY+EBz8/Lkrb024FO4W7n+B44EB7CYnfE/74rTD5hoaTfy5Bqi6nDos89gw5A
3ItIw5hUBEvo8/9K2/TTpyIu9he+NA8AZ+NdmQgZeHoDBSkQ7zFZdVlIMRhcFiR7
eo/fsViLALS+WALq0itbDVwMiqzkFTGykhQ/BLRHOjKxJHmzdZkuGLi2wp6fwqj7
sQ6YPX3ZFh+BvJgiiYTaN6secPqUDg3DI8OBFyXIJZg/4Rsfzq4/zPwesoadbSS8
n0q9yWBJpURd34ARSSvENjJ7iI6+SZF12OtlE0FLrlS2yoM4Evm43H6S2faA8WRB
kCNbA8++CURaruD9CJJ1siquN7pU3qc6TAZ457UKFL92L6ZTvz4H8XyQVyUMn1cl
U8w2lXzznjdJiYOoJcKL7Een/GRnnWbFqidU4brrDycQnNyqJDMZNl2LyxEwTqrI
UjqVj9zSlnOFAE/pZiS/QT4wmvkxki9o2QX4LdcQOuWd8PsADoR/k5X0KyoVk9yI
Tddw6vvZpaoBEaz9tEC/wYEwL2gQyCl9BFDEL8qjVmNX5li6GYWRPv+KblLKRuES
lFyzqVs2TB32iD10ea99qRuOaNbDz0CtjZUBb5GOrypU0gR+g8n3XHeJ8lmSsyYb
LdaGUwEPpJy1cDS0eFxF7VRJCaHFX4dBUY3utZO++iE3auVOBu59QPIx8N7N4SyU
KJLiz/FaJUFl9ZqZBFcQUmIBUrAFbu2300gnMehdEAo4eovUs1SFjwe4qWP+hw55
9BnR9jnVsWMKi+64MgCUcIw9uUzXwkBJMTaBXMCScSotpNGblkNGZ2nyUEegSvwJ
WIdyRH3B+qJcD+zEBQ4fn5im7hr8yu6/ZFc6/m00B50WEACU7Xru95BaPWgHEEhU
94SVtHlPYdb+6pTQCn+RBsatYTQIglA0cwZoCucDjAOlluWkq8GviAxMR5pTbkSV
qxSA5KOvxA//MCBpU+AgKusbbRh7CAAXhEobtuOULV4RgRjkPqzax9cGnZPBhOYO
Spv+oosgsQ3/1P3YAo5n3Pr9Wf2w7OnYFzh8UDZBRQkOw61vyXqsUiTTvv9CQofq
nNC4YvS/r0BE4ec684kUhuOXdRF08os5X7Q/bV2kpivUdgpvsrSU45LJw3yb2OM3
48l+e1miuGf27i0kaGSRspLttodPgyLuHJ/w2zD+jzkbXyvONgch2Riq3eRkKWt4
fWKAIR7mKC+T51UfvF/FeFQYVuOEXBud1S2JBZ+Xaf8Hdn41mdP1Ks/uiuXj87p7
53NYDwtTmcJU4XIi81oTn4wPLWvsF8Kuk8SSPKx5Fb4opEmVggiHq6UqntwZ5YCG
eVBflUdiOY0TTCH2qxclaWGLNe7r/DtX3WX1PG/gohZp72V3XmParJs+ttDdgNso
xPXSbUX6n+EyfHrRX3WThSBJTcoY9PjyKOzmxMObOMSHSlDm5muE/BXyUZWlVAbZ
NvZ6ETRXTmqWM28LALa3i3oQ3sXt3Cins5MMM5a58T+8KL7okksWABAFpZYvVO7L
fFEy2I0+9EROSknn+IwXRLScDWtuH9wvsO350DouudbkGUFgUODszSw9dCkzk5bG
XrR1dScKI+UDONajd0sEXJK56nfDTsWeTPrwf31FW+gTnoWhKwcPDG97Ks2TC/O+
m3qSCPkcwZz7R+giahkK79G2NOY3FarkpEIRU18rObAsjEmRGXObtaWDWTexkVR0
CcNx3JrpqEWOjAXDLXqM2QoSVX3FDhL3fleZ6ZXv+HEATyguH7PIDH0j1XW9+HLd
uVFcUDm7NCbX4zM/Fo39HTblT+AC9MX6DxUxUm6J4HPB43Gi1JJhDWf4xiOdvX+h
TObaNfJIiQvNuqpcF5LlTbifhxmlA928tVn+OZv1AQnNtk4VnlVu7+HIr40RlNSx
sc/krHyMZqZZW4K9KWbQpXg6Mp6ctOCx4DNQlmN/obzumUhxXvCqPGt63mjxSQ0D
ykQ6Uh9bEjltn5aH2AWoq8cPXSmy9ruZ+QTIAbaqZoS2LuY5p+AinB8DrIyX4TG/
QG+c5VSzeNOwEkb6A/+JRXgDYHzyRyGZkSYZJOaRsvo236PDsW5bXkDT+ZQjFMxJ
poH548h0CbNci+RVD4vtp3hae20bzHXdT10wTCZflIHtJaVwLu8qlRDMCiMhSjT3
kmA7jmLiM10tW0xjYHXH2gJew8r1C11UPzOC038EDhAy5SFcVVrQLicCdYmLyV0J
VKIy/jhZbJMaH8iU5MD0gAG/OU+R44tab61sycq5g69z5pBY1VdFpBaiFZlk/PVg
QBrYFsf8HoxTymcDkwcmxx6snkcfp5mbslnbNOXw03VHcjlONxh50vBlJCtBC3bL
Snrr8Je7/+dLLiB7BwClm265X7hc/nzYzbU9zPIMMRvt1gDVT8UhvO254jNSKkKX
NoYGj4g62nTCMZVnmFvjtkWKaypGV0VApVWO4iMpcoVgs/IlTgGE1V4Hq2deh88h
iCzkYjzTE0hGiaJY+Ru/LSBJvqBfuhQuLlcUvVTRzUz9hMX+iKnlhiR2pWU0J47f
iHxwSYdUKMxOcZm/fyEokWjBcPOR9UOTyuZbMAw32u9ovkf9PA/VeVpzgxcnIN9s
ISqKXpcjoFUgnL9kzXS/YD1E/OGxxCZgYpuQke242OLzAi0vhO4nfNuxU7RpBP+T
ovHBjua8KFufjAOk0p7ZL+R2nJI3uQJYPPKzkcAvl4Rc0KjEThZPslOjlghP00Cx
aAi0U2p+yprJjOu8KMt46H7USVib+tGJMFi5RfbNOLgyVgIgw089OhXPFfimIZXx
9+iElDEKrWyrrzQHbjPsaoyVmf80TNIH05LiZtTTJ231Pub9EZLxdYhzovXjv7hy
m+d1nH54MWeMoN6TY7mg6HwYanBn+jYRfLiLpbCVrZgO1IzUTa4RsvlUykH+h0So
KgBui6D0W/1M71aNVRAbD6VkAKWfbCRBAXIpjhvL5/zFDmR6zhprXzIDJLVrKXgt
UgkBIRwnyAeVz9/XUb1gKzEJJMa7I3YYcG53lO6iJb1bHemtuBt9HAW/omXv9Sru
aB1Zor5J7DgVcv5MZwD9HlHW97+LRczhptEmZ0mqENH8ZUQV45duoO/X+QacqiKY
6vnUh/iqyJzrpHrmQknklRsqcy8rgwzfNdZGycPSs7gnFrPL3y6rfFuIE1C+G4q1
tXGzeT1nGBjIN1ocF0kYp6S7cweIO08R7No3mB9vrPBxTJioG/gJJzhKX/hK3lHl
oq2H17mYfAH8fc1ERePI+/gD2KOABPriw6uEMkFJ11yHKKvnweuB6N3UVpgVZV47
TW0dmb9IyGHEIaufAB9y/W4pE2dG7FVYprE/J78y6wFn7Pc0IQBAb8lbPmwhdkKf
EKN3nmNitxbK5LJ7G3bJuZhd8Jbcbt6X2xQ2+qpc4AwOPbTJbw1XHangHK4F4pna
0qJOT/tKp6wMdghSpiDk1dBdyu7APhFdd9kzVxA1I3UkaIlG3+/zroL/pGwRN/xc
Ft3Kw2fHAaD8hv+GipPD/Hkm4d5VdFFH//9sOn5MNTosKUOIM1KVt6DwKNSqBSCu
FZNy8dmlnonLcGO4U48G5rw9dfge+pHxQw8IHaksQdW6G1nvdYwVjXW0fbSYYoRO
CCZ7Rt2qbGZnF2gReQ/83+MJgKHG2aVs8YQVGR7EMUGzpgoXmTty+500MQFLPssY
yqrPsqJpRmoffp1DLbQ6aYNtxWICTaFsU6T1OaHNrR9twLUh6P7rxNMosvXy5D4k
9pyqmm3G9xlA1LPkrXVo0aQjE0zHGKrOJaFgqrHcdt2/fTn5XOSjCnvo2cR8wCXi
u+YNnnCf6j66vgKO2zzKsHJp6QVZke0uS1mp4NatVilPSfTtpde90ZQWN+p8c0cD
HbgLE0+QQZsWPweVoOwpGQHuK1sNLl4XHQXztC3ToVCfU71R9aTOQmr052zXApma
jJ1cAiNYUe/ifDDLap5gM2gMdkrTe5e9XopOLZbMRiKdgg5Kvzt6LW3lmKf7KBO6
PMuYtoj2E8h21PrlUQ9CJI5EfIyIYKp5LlauInOY8HfCLFgprfaDsv16ze+kGcki
WVdZiqh3qAyvYW4QzbBxrCdHssujuyM337Ls4B6mQTK7fKEwvK7x/je8igoS/VsR
0rtmj5UIU1djdIeEkUw3lN8NwSBuLSbWkhmedLXl77nz9S5QzgPFd+kUVbz8EMFR
cR8VVJXohp/pW7FOcGPKYzkIGbVZiOrxF8lOMyhFWscghYNgk8jMwZFEEtimDKD6
yuUIFhwkdaQcGq7Q8iSpqliXAu9vMwMYdSlgnzGvq4Lbc0tYCon6YGczribU6/rk
xsqBDj9k5fZUP0MRMi3l/8BgxHr/UCwU58zZi/li5EE42OG4BwoUv2iXtL3wOhVy
HdlfC6YiOI6Bxg10HlVOjXhZOmHtPFPwZrhD2ihCfIZMSFEezSNdJhuXXAGcxePq
DipQRp5z1UqoMWUWKVzWU00U7UzP/SQjPBlVT8EFytRhxTtPUTF9KBD7a8W+a6bT
vvvj9MDW6NOT++GLYmcmG523l41o1xZuutazDGyjhNa9h4hCqSwtiNC5zIuAZskC
yGFzgDSqOOgIVfI0ixYx3fUEFxnpZfwaHnEr26+uIAf1vD5/b2isPfxJZwlyLs01
frpMJc7Na4iPuKxDFPos4MNh0Wtp0TNUwXStm/r+l2QfaUSoxdfqZ/J/WYYRru8f
dsK1GtjtolZv5lOevXAmVg7EYlZgwOOkK6q8laYscQbpH3Ap2otxEJQdTzdHkUxF
+3YK5IMWocrNkok5ytpeczClVs4+QBx+9afHo8/6PAZ3kfFeN5CxOdXdTPnHvR7X
lnXTerTiLCwiSnFBFmnpj2sDXDqg1YFxqtSbX3oQnnVfj6hrWu2ZlQdxjx7RueKw
acZ0tUhEqLHqye6quYWX3UdbLR6BQyEkIrTjRshCPHZZH7rhVfto0pVezefKWpDH
jUj8ARd+N0Pjt4veeKx2BcDxKQUVsw24j/M4rNQXlEKfo3gRHxdX1S+vLcgorTsS
Mo1nkNeOjMISNieeIX7jXnkA1lyWyzP43xCIPuaTmDDdhCSrZ3tQwwX1FLBer2ql
rG0foZovUxDPOKLd7JpxBIqLSWdVgjM03kLpvrPcf+jTBRT4rFYpmNMxqudEaJ6h
o/IBNXgs7oBNafxyFc4LOqYMzK2Z6ACLTzHYkBxPzyEegDQKl71hNnmqbUV/pfKE
5bvtDDDoVtHX6BBwrBv3mRSrO8arxTHQPVBQLQ2d1mEQPj9NtjddyJq2vX/fK9jo
FtJ/CgGZjT+w2Ba7R/chS5M4bQmUOq+enM9o7bb1yWI/JfqLl5hZcd+SpExzBpmM
ZobWDd+zybTKh/7Q49QJjCthljV2ZbFE70w5DVYoKrvFTGsX2vtVbMmEEJk7v/Qe
qjxe6hjFqGqhh7qm7oyrTJVE50T0XrHRNtlBU7KZFbCOdqT6SgbwuzcGFAcyOxBX
cyx8lNI0AdoCYMAjJf5xtwhdfnK3tJTdmO2zs7zeu4diBt0YpUAhAGmiueadpmi/
+La9lBzGMYXLOtPTYY9n/5hypzH2z2ZtpvUQ0yVBhQEltdiK6wWjctsLv/IIa7QB
ief8606M7F4SVG4Q/X8URnyOxDnALIQkK4IUvVBTi+0tBYABoT+lnjdRJMx8njX/
Cluk2qsexk2JwPKe9+JDybRN34CfG1JAKWicMsuYURT3PAAVlRVarVKKlAtZMeOy
wlnkcLtoEoqWDEYTiE9hpCv97fI4+Zu9TiYIQL1leAxjz/R1v7Kjrm4ZdbmO9zUm
MRkLC5IYxa2qaagC5PU8eUX6RAr+J+j8JtThy6ECWD/lpcL1TEm355UqoP5u2/9J
/1O0wSmikjDB+REERXMgiPt9pin0C25s0OHy4LFJScV6u1N87NM0Y15RLW6hp19W
1mLLAn7760SSGlMsWry1jbM+ZrCwdeLQq2xOqUHgCFnKO+1uqhnogrbC2WdlLLOK
NVRe7Px0sieF/57Bm9Grj7gJDy7DjkJu2Y4ETVQjIq9JTe+Jo81fr9rGlX/WBOAy
Aba0b6tuwoTF5DlON1EiJIHZq1NBYLA31r0VSk0KPtXfrWAbujTncw5tqDYbOHpu
HPGWS/YWDcY9AXyndMxVmbmEc4zyn+hxqj/mnlh1DYPlsIi/ABoSFkcRn+UV5rbE
D+DdrZkLsJkjAshw6Y822p3+bwiNh/SeINdbdY4tfUSWB/iwMWM4SJlAdFkyNjjA
KPCa45eGzdhkHU86KiVECKhLTG3AG+4H6hZf7VJf3IVlb3YWy5FxFPpL0NAafjxS
g0/o6LTYkYOi3uMvxG/Wnv3slVnP1o9z4cf8FW0ZnnxnODmpPFX8sPBP65Shob7X
M5VQqj3BBCaOFCrVOE6m4lUT8FiVb2cxvy+dx3G2HL/2TvD1OGmpTDGLNubeRSBV
iXRpft8QdRqksBr916X5wjkj1dIsxsnl8GtUmeHtaaNnyOOdJNooV+FHND45uvcj
t4YHw69T7lfwsxR1xw7HdIXMkmZ6F2qcLeaJKDyxqi/teDvmduY+R43OqWmwnbdQ
jEzDcLzRWS9EU0VhDo4oZb5UsgdDUcBQFobhda4QCk9tsE6fGgsrOvm+cG+aNsvf
ZlzVgg37/GQ1CIxLOIu/r+0PiPJwOK00f0K2C8T08YJqwHIKDlkq2U2HG0EI7tvp
2B2H0fgHr1nv9l0ULJh1hNma1sobYu9GxFfAcwHC0psfpI6ccLOlYzS0Z4jqH095
6zAWuW4+8FyZR6C76C8Ir2+0MXaCfNEzb4i471APi5arH1Cu+XVoArUHkYfMNLwz
fISld4Fkn2L43qSJ70t3/6f/SYYCO7CoCXi0Afv0V6lLKsqsh8QIQnr9uYxGhqzY
MY5/yzwv89TxIHdF0LXss9OoRn7j7KHrNlrAfSqJxlxrMjZJxA+sYK6OyFY+232y
v0YyDl/YLT7j8tMtlZkgO9bCAq1MR1d1jZ6mAzPLmpvtpKE2XvaMDYYeGeX/Cpwr
G1KpoRbNJtQA52hf5Z8Qe+DrYDhZW/kxxA5pE1XZ4t27lnnHPygpQ87I/lAbFI+G
6x21KQ3NYzJSBQm2u+5uP3MrjdlBf8QPKsKGFtNI2dByA1+jwM6jRMnQe3+1GcKL
OyBfjNRt2wWD20t3xRU1hpMC9fjJe/+wncvD3IfnxFGXHMwajUj1f0K3+BLXWBcW
FliiqfP0ZHtPy3mIF1spXQlVUMxi0f/9eiS9EkWVnI9TyRqIoz8zSpmwUzcys9ab
RWTXnxw2mcGun/bxUTygplDu9sL2uGWC/d44DGL3/QFayxLwXPDCVGsXdWP+9+/p
4C/lkHff/5XJAbolgK+jjik5IZZurDbIRVRQYDAd4HrvLW8C8gXdSWdfdVXPLXk1
P1xs/sZi2izKbppacIRC17vVjGssgXD+sMTk7J7FgOrLC7EOagO8uq4qMr02ZblV
GJh4qOQpK8G5qS/REJjB8Z/Y17s2tg54xpc4hERgVoSeCf1DkPfTNV69GEAKYA2z
FOdRr50Ce0GVjx4Cb1nsgkx7w1qFt+WBdk7tNrl0zFtMexItnIYLzzn2EiFPFl5K
Fg6bVJy1QKf7Odun88OqWG5XZ/RJFxlbBugUEHfEvgIv/MJrgu3jnbzVbyLM9M6s
oPYHi5e93Z3sNU+nExQFv5Sn800rP+crJlH/XJK+HyogyTXUM3tJ3weFm7VeZHYW
jjBtQlb7hD/o2GZtJ6yXkB7j9VlBW/5WCN/PUi5NX4GPyWclmC+qeMzt49dAuPzZ
MPKnDjsilQaRJi7rlHybel/x25HK0m5nvT39XTowGBU+JgSw1Odzp0vgrpMxR8Kt
WG5tm7swDuCFfL6DIj9GgiwlOMpbohUcVLBrbsBYwyKPFjZCU9PBqfbVhxXG4F/B
uwTxeJSD90ZBWjkq41IpAE7rFP1BH7nUmcXNA0FWI5mOjX/U3LgjDr04ilxPByUF
1fxZa2rP0RZc80nT23fYIoC3cGaENtAPn0McNGC7x/Mycj4epbXOjCcS2Kb8zQLd
v8LMAqcw49tIYyYPs8dytBSI/tzRalHqsGxpbfiUiOpUN6Ozxb1jrefPAlspSX9X
4cGuSesjAC6H4MnDqcDvkulAVF4mX/cnkABtZNiZ2Xfh1EFBEpDWlL5V5RhGimt2
OP7lZLhi7N/dMW+UdOzvP+cMKI/QKSH7qtnRpml8po3LVltH6r9CH59j293iaZG1
PE3FUdsyHDdUvbRDYSJ6g8WXzkLmi2tJvL7c3MD62BtQszuJXhMI/i9ShXHZ/nE4
kmMQOTBRv3ChFp31RwhDaXuG/CrwKDRykTdJ3P89+gJeI9G2WzFhL3wCmR3GQmbZ
Ldq+crlwz5IRNbt/1wKgwKtY5d92LnQHBsZkQLzszg5xFytQbQtRhAcXsG1qLL2v
4OnmtKciESb/xOD/0Y4ww2MrJiInR0QxgZnNab1jj0Wu9Ltml/X2oyK030Fx2r/P
rtt0ewJATSXcd/GPs4r38rWunians1/F7Bm+4kTcQIgzPzJhnp6Pdxu5hc2gZqTc
rxhW2R6uhSgzYHkNATJewSWz0shpoHpYuCXorBQ9th3UJA1xaV+pb7BvRWKQMHOc
D0LfQalZMqkxnOngiLEvkitKUgK/jvVKqvLKOGlv+IjdzSzPgaEuqsevACJGoeBu
tu4HeefxHQPEhwYKYoF4H0S3V1zp0mx/JLYdu9BiqpZZllmygb+eX+BNEawVltLq
Ct7uIObDuom9P3iO9s528aj+jWjeZ4IAORzZCPaHY3PJj+8H5+4NmrZ0CGEX/jcS
89Lrt1R0i0xnl0i+wF4kWTEN5nH8sCIdaeZ53v5b+QegqYQVUeF9o3D+3X00Pvsp
RUTdRx2OPhlVd+sQoeCf1ZRKjY7pYM2ReTmDPb+vBRQ0J5xTQDiVIHLzccPMcDTi
0vMQXaRkBWrUjhVoE8Eos0WI7MzO67S0718hYuy4LncI0hvhsoVXZNarkhseCksp
tQM+wkXGmWkQ8rk1oe+UxB0o21FG3Xman3RTBY1g3R4oEsNpKXhKO+ybZsDth2uQ
Gnh3i8lZuxgP8QXSIiWEhsQC6ET927w3rz5bSHC2TZrCfz4ZTUxuUj4awkoa59AV
FOvzs8fXF39tHOcRVKjndj2Ru2gGjOVt7zcMSBQ20at+hDMVQe9GW1Yy3dzdfCaA
QoSnzUMot22LOsS5upxuF1WCdeLytsYtC2BxXz/AhVKPiUL6VBr+cnnXqaDCt7KK
yQ/Rbgoc3QQGieBCe60+LBTUE5o7+nfPcTy7+91RkIsdNMhKa3tuPRjqpciXodhQ
83MmqoiTc3mv77CYs554FdoKBiN/4HjhrlWCBT//VHQxtRJSi9b4GKpDEA3VmOgY
oltPMtxUDBOQC0G00SJqdQzdjNJzzKF70RJRulBXBV5PvwnthjOhcEUInlrauGbB
Y32CJPOaPQSNzEYD5G4F5s5Y+bePayeOlAalDKV7UAMdvM4SiXMT1oyWpdxFYa1z
vgAT02TYjtr/ynlaTDwyGr4EG+PuQy61P+vxM9Tl9DDPfVd0CxdXd+NNhlKNHNlR
Aki8Vu3wQSjt1IuE1DGWyPud4gnnTxcaEI5rTPckDDXoY5Megeva3Tn+7+6fkuYc
C8ll2t5r05+TUQOHCF6PjijNXSnSpswOgQIN9tyUgEMlJ1h3+gC3VYdLM+nqUbld
3DYQFDD3zdaKcJT1w2ZEBfH3+l7Ix6y9UEhBX/WP372FH+i3VB+d5gU/JkOOkmgD
CL6FhHVGQFNg25ezH/XAv/GTIsnmw8O7jetBRNTBRPQvb+G3qX9K5E+YGXX/BSP1
A3/Qg9rry5PEzgoGY8dOplN+cM2/LQaM49SFA9coiI2Hh5bgzY9ePnyaQCIUrgSp
6HNs1w8qhtCku1ikJ+R4n6sF4iKY1uh/7oVUETKBmjV15twbf2Ej/XT+TDpWvHUs
LHVTELl6iUqHeot7heR4A76jIoOIVDwQk+evy4Wf4eTY3AnsU+Vc3duPZg3QGJ2c
BlUNOYx1OxhyUM49bKUoMZv36gIhoddDL70m28xQVviO2ond6erMNnp07pXPX028
n+E238s/lqnXadDkhJSG1gzEMkEh4Bcb433WuWlOw7jHUwheNaT/wWGR8wjXMFBy
kliGXq+DhliIcb+51eMCU/MwnSAwn0nUEwgw4zzCGc2pL5vHaF+azr0M77gBLUgj
zxqb2rK3UZ0zJoldIwnfJseKnN6gKeqFMkidcjhjkr2qkNatZJ3sawKFHFQgEkw1
XJva05/dY9WEUb5pK4miEzOzihozcb+Alwsxh39nPttI+FQ3cpsv2iZV4Wz35P1n
J8emO9Wl715dAqMqY0k8wgF5V8BVKlOgf/gwkybiAZJdeUfdNBg8QiHtrh4Ivnyz
DD2OHlBfVsamqm8DsacrC+aQ/5cpKoR5nNxhMGJ8NRtDG/slIBJH9hIWlrEI58OY
zn0OGjqykWH7kha0CURHsr1QmmDRVnRpSZJiww4epBgGLovC8OBTGvSJIGpxH2Fg
PXXj1TZ7iKHt+ScSFUuuqIaSbSSoI6aX0QO5aKbJmEWeZx6Hfj3t4+1vPIjOljpB
gsO61J9iSBYNGlOO99EyrISnEGfXmJGnAnuOTwFj7wXtxc+6UwDV8oXXUG3udNvo
oa8iNA/fWgKlvHjjUYYwZPJzfi1c+rEJUox1Qr38hH8BtdV4/0WRyn3HkgyF/exX
iY5VxqTajzTqce7cp2QCKt9pWhPG6zkWf9dXTIXSEU8UlUla6gDa7Soab0AEr9KQ
LqH6loxVwLOWLiIFs6RWUaypJtqmk+JMz0aIVbaggJJBPHvgwVRTbGsA5GRYvI07
8s7Zn5QhC5wKsEE//3YZWe/u6EOIiPGPZCqja6sFQDS0eyUF0M7sI/oQIOx2Xt3d
/Z2ZJ7unC18dQA+Hh0TWa8xfrevyVgDxyiSM2Ok4tqSvj261cM8ydJ4q0/Co0LVi
s6NJ4jfYV+K0QTqF6wkvEUcrBo0q/BYtHQD1SsP9bWKpC0JOWXIfIeVEfLPZHeSz
bY+diEV2Z28+Kcze9MeeSjbUrjCbpzcviO24rv/4RzkNm53Cdu1I2afUZzxFoCHr
eVLQBIicgf1CiqlJSYn8VwlfOv2WbgRM2a9kYVAVbyWVWK/+LqGmDDLHo0I0IYs/
Fp+AqCb1vxixRZyMMYpkcjL3d/NnwFTkrb7JYk+Cv0mljYVJINFy+2kKGLUaZaF7
e8yZ0ZGjrcqMplYCqXANzHKBG7Vo6odfOI8mg5oSdI3Z7EXh/aUOePQJprnxmMU1
2Lo6eLwulk99zGzZxplDi9o8iGJQ398pVGeytsA7g7WhRH6hHa3P2mSF6swsMK8J
JxPZb8wuVC4RydM1TPwKhshu4ai2rbvUQE1uTlipk1PfY5pAzZ50Cvhv8aE2nuez
X+Fa6cdvpUTL+scqin4INdJCg5EgYeCoD8HCrmc8lD54AIhJirlsb3Vql6ItScxN
ARp5om6V4ob9vGpBfj5iNNwIKQ35lDiwbWjfhFatzAmw37Qx9rHkV1nLMN7bjYDb
8WsI8ir6dJ33yAd70s5Y6to54Mgg/zDgHh35mLvzrt1bCse/bW/8qfqOYwsxiQQ1
t5/QXwQd6PiLaSukwUuolZtyBqKzr9gQ2TWMpfjwSMNafZMS4gd/WizuKwdvIKJE
m09gjXX/N+R3h/B5bvtpSDi/HZZs2o0qAlbyVjzbKemAJROTf/Rap66ld4Wprqqh
O/CAEZViGpaHIG8Oss5pbOwcQ+sYcKAwMIBZT8EU4w1+WjChDTXUcpZ0MpPe5JDM
vZQsT57VdO+YhQFKP316YdGOdVgmBWxHneQ2jf/SMySWDMIyF3zh/BT5+JtM9gTO
TdRq7GpYWeFu9pENcMYCvKHMgIt2zFul2PqxqCQm3v5biJkKrLkJOleW7yrs7MLA
RX9e1SNDWxDxHQXmd3O+7tm0Nbr/jwunlGzr4GgR57eqH6sUPJrPwdiZv3ibORfI
2nWXYlkZ81cSvgIcI/4IobLs0b8Q2CjBVn7tkcaVqPXhWE2wGHPFECXlDX2obazz
sNb1SAzlHgLOFoS/73PyIxxQk9q6HJhgmBnBFCEGMhRRHML+fZesMNaQ5VEs+lIA
5kLiSZSTPl0qY9nztqftSp6fRu/KyZ7JsUDr1XZQawhTUrZOIhyd5kPsaxGJHmBk
tge5sQfnTznbQW1OOrQrWSuedb6n9BRSgVHgTprjtC/0s4pvNNrDWjF70Cl4CZdt
zeowaBBlEEBl2y84DwdoIdlUmWouoLhV+BIOO27QX+OPMYlO8AL4xRmp7RzpLQKu
aM+xP+Z54GfyorIkhi9ziJXM1OK6VO2QrcVR1gAfpBnZwVtWMCk/H4ht7Yb6UTnS
t80eBrudHG9meCOMHBsQf0+CLHXMM4lwaY5y38R9dRjljW1ghXbFeD//8fpnZu0A
p+yW1VqxsVdhZapMZ+/RjO12pQqEuqCt6aOWMBJYU+eT+9QmWy/NucuOP15qwYyW
A1SfJ4m59MZVxR06GJzNLVPnL8KYeuk3z2AyO+rexdAagWHX9FnAqYVJyKJEFgRE
+EmpXupBudPufr+/hGXu+XsGYNbaEAxpHZBTROGGpumlStlmxNwTLZ1zsaj6HZ+k
eWHMstm42lns/S6rfF4OBX5tXv2nhYVigLRShVFfK7iW3Ha89oB+PJ7DPVXSfqIl
nLtQb4CN5HnKVDW3K7M/eZVImMjO1wQaDyBB48rJrL1knZKTpbWwFGfnCf/RfD6a
eTjCfQZZUeoTRQzl5UpmoPplv11kaE1soNSDe6OWxalwA6lPeFHzJ5FCmKFbgMSD
qM2o+9e4nDm/alqBsxE9kRQoIljOE7Pmh6dgzxmPqE4vetQLf2hAy9KxKj/Cjuuw
wjjKCeq65eDDb3GfNkt+1S9MHh5IvJFleQUVV6ODjG4WnXKcGbs7s0Z7ARZfkIJu
dZWjpmeFvKrT5EWnubfl7NMPw56xMpWvcLL5cYkC8/BC8i+vul5l18HxrNmjwKeI
P2evmrOzUi1DmriAJ6Wh6fLKlDIDQxFpfJ65xnSFzkECko6YQ00T94QfcVDaRYwj
0M13bV80BGeYldIdZQSeYcTAQaEF25MDpiz9HSLvpP5bHB4pz/PDPALCXVH3Xth7
Kk0qy9Rrkq/wFOpmMjXAqqB9SAXxCMWVKTVcMUUFqx8gSIwoXF4JTZ7eLn/8XqFl
dxTan/x9CobZ1T/ENJN17erOF14/Yzw64i2ykg/ZfP+M5FtE/7AcfQgLMTlNYXNL
U4/osvnfGEzrwGl9jEbrPamVtwzataPVxgKENWVIk82n5nlZUwyPV0oBg1SFk17B
TtPyi0sgupovsVcsFiNsnnmFawiyWrlyJ+CSzKhPZ/Yc/7FrfwD0npLMuon/Ex3u
5ql0pQERmEX9lVWtPFbD84qE62MaIcgyzKOEQll+TQYCj+wRcogG1PWeIlc3+Gg4
VjWM4EmQs3gEVVTpBuMtu/1oZOICsZ9306/wG48XcqnaUDVzMnjBVv2vKQmmJaMC
+MSqdEXxQ/0NNJLN0b/TboBAR785OJCYXXR33Fu5jmFzvXb8O4cn50QY1kYqlexZ
Htyr8AI07Eu3wyYOfO7gey3VN8M9QGzj1n7FY5Ag1/qngbt7H0td5qcq/c4/D5KL
C1CYACZH1eGpmDaEsw4XMztFrF+B9Vl8Lf7QgH8ES8XJa1sC8yhAN3w8UaJC4Mo1
1t4csE8N4xPsIaz9AjkrOa+UwtNYNfS7AZxJ+M4vyTOi6c6vBX8+G5IsmR92WBM2
//9NBOhUG/LI/jBggtu8Gz7jDvl2w2tZX025cslh7Pd0ideifSRRadjglrpZMd8m
QPFcy5+wG+88s4XnDKqRalGQKMrKhfrIo6z7p1HAWiMSX/j0rmKJ0eN6XxubVsQx
mX0lCJxMrRe3l9bMyoed3fmTlvTFSK5UEWUc0//X1xxlrNfpDgesO63ZvCB5xEgB
3NpospX7ihSFzqHAaaE/lm9wq8HH5uPvp78pmFj+mlxxexpTC1J37WxOxVufnP9y
a5Qf4Uek3NItUvQ21PdRg0sAjeA4HVdRBnBRy15TST7aQBzvvI+nyPGoyDS96uae
9+9A29avOsVU5LidinaiIayYDskTwZ4fsRU/HpdWaIZ33qzAeOp4G8c3kKiE/hd0
2hDLAkMI1RDqIYnIfWubcJEiVGxJcGv5DNupK4c88lMEkehS4yV19+ffpwxG/Hxt
iSbUXodkiFC5BC7ReQ3o2tqCDMeN8qKWE2C3zkZmICqksFawNtM0uJh+oSXmI7Ez
H4NocTOokWudVLRTLMT3eJBUJByT90G0+TSDxaQdJ59mZscAB3fQMyJXRUAoAY/f
8SXyfWJk4lV1iwe1QcJ4MqYRRawP0HI9maNoyh7vh//0je0n8GlmAu+NXM0cUZqN
aMaQdOqlGUSGFYod1XPM6P1V1gVW52lZuaQoljVe/lM9fFiwQQsEOhlnRrwF5i5Y
X3uq5lMbmWcBqfavjkZNuAupJEELCSdUF4hIIQjlo8iFxpw0Gswq/tIJWssvlnIm
AJ1KpsFfxhNwxQL8rMz+do9Ub7H66pLm6Y50Nfb7qeOww4dQHbIFZTgrRwvp9O0R
wwP20+hzLy9aSeoTAoBG1N9Zmaf9oqe5CIgO+4BdJTPKIuN4T9NKKbq/Kh+64ELU
xgF82cbzvGQwU1arGgP50UTyTZf3A0EFfpKnEemLs5Guz0hdHfB6EtBeJo4kzon9
ah76BKvuIHMvYZtqEGB3xgVINB8yOQtVEVavCjQV/gDsyx1E6GU1Sy1qmaMRyDNa
I4iOFZ7U5fQapIdCR/26l+QZr1Ktv+0CWveEQ7X0UZ84Bq/4LnsrP2+WwYmSJAEr
egrsjjPWkgkIiBdTBCEHVYKbF14XBXDTNb85uIODtOwW+L1xX7zbquWB/cGK8B7Y
Q6NiBDy18X7muBkfcWoExXWdmu+yXG4Qw9xx1pzjem8QoUfYRDBlwbU/VeRepQl2
94cTaZF9w7DhGbgHfpPk9FdeDMMYfU0DnG0qyJP+bLlJJRNpvL6Gw5Vl36KZ88d2
f77EFpvzXNnxAnAkRUVUjtRs+9Nb00tdXpvd8tv9RtNDt4oFIOse7JCQalY1GK4u
tE77rjscTxbfbmCIDc5k+WZLu+fDSilc0gW7QEd0nIX+1Q/z8YtMDo6Yh3Y5bqaD
sMMX9irpRYkak9+NuN1gkqG2lpr6bG3KPPLwVFvWgVwb4Z1TLzbQJ1S0+ePz1xw6
QMwxttnn0V6a2SR5rgl//d0XWV2XBwzWG/sC0lZP7K6Rke+MoBKhQ9RddkN0Nrzu
/FmU8Ray5EBP8gOrqohd63CSPX06eS3sLAzdGgyNzV8Aawe2hCssv1EORPUQINX8
cuDdbR4logL3i+GMa3floATUoBZqoUKJs7fPUy6vPp8QIDpFi+sVJWAkEP0aOveO
VQkq5aZx8YBADbLYscJLAZV7dtoa4gRpSKYDQVPtypufgckULEpUV213J4kWRwC1
LisrNVPky3gbqmOdC7F8VoA0btEJ+6yonbDvffbSfbVlY0hXq4pQIODduagi+u+q
skuf659MNKhd2qLStJGOcEkDxCU4LgN/4blOgIfC+OlsUTHMf1SYJEP8AgWB1Kvh
O/pM8wjxQ/Fk2LLhvXKEQH9mwYH/a40IKd39nxCki/nO33aQWFhCSlgudwL88q77
gi9gGOagtEA01WNfyYZ1FahYbX8wKqmqtRM0XhuY7xxVAqbi2SXK3pRoJYOmd6Ju
HyLu0OH/+wIAik2M1Wqo0yqN3OFsNjW1wXttC0Kl5L5IRkRbaEqcdGQtrfy0Dbct
KT0i5ysBjadFdZPrpINlErzylOtZOZk9Ri7ZI6b8jnGDfbRbFLWPvfVqyl/XGN3+
/s/qTfxcIvHJ6rssMrUPVoYARPzYXoJiD4cFF1EX0/yC4WLvxIf8FfXPPKc5PWF5
mJoKFWy4uO4hPWMxFmkcDkvXmqCpcRiNotqemRuslcgRelgA9UZ/DT0xEXqyMk2x
8FOVQHOGfjfeRBaIuX0Aps3RKdFDXw1uCvTjBo51hIDM+pvGCbbG/VZukaWQrtOX
OYLMLbKnUD3eYfiu1VvoDm3tPJHu07SPKAVpA3fvPxjmDxFzDBAKtLS5fjWroEBZ
9c583dyx2oIkkhopo+28ApVI3nVfZg8HnzTVEIVFe+7MVDnp0KxZxGoBD1SkTyMq
5QPxac6SOc9I8cNFwIXF7ZkH8GMtCLftKn6b4+89hMcAqSuc+8HE4UTrgV/CqjCM
nnJqVMaasuRL4Q6ifeyNrX5pksMvtw3dqiPmN+1qEReRngLsXg0MJwLDyYQJciPN
V1yAGgr8a9UgAP/Qoyss+roAMGonItCYFbXo4Mg3VbNBe3kg5KUf7/dIIXa2fc4c
xAxaN63/zveIZI0pljbcJgdpAjA0afa3YnkG4ldBcxCgRb2Hc5Nlc7R09OQwipCn
mmOC66W/5IyA0uLV0scFXYxBr2nSk8hh6YE1eLyuMtdy8xjj29GDAaBrCIFreJOF
kqC/65ra+z15p8Nd9R6vogQkTfIEBhOpp1c3XNdjUXZ1BmxNx7MTkSyM4cEjkVcZ
NP3i/co5SO8h3/WHNjfau96bCsQfnAPCCJkfiQ/S41UiLCVAaLTh9hutopH8sXex
2GxUi/S1oonN78YhWsSgfC3x6+J8VwPeHbS59MDGxK4R4io8lHf7m5D861LTgW5p
Xsw9p5jqt+9CVFgRKyWUFGB4qgx5o/TSKnL+fXjaxqk9CQCCaAulURimtGuEagtK
OBzhn3wSHUKSAlnS6QUxGM23liHV2jRdNbWPRnh/GU0Jd262EG97GjFSdB9GP9hO
2dw/zKd6q9vMyiVBVvorCKVMRoKYt2+QnTiPFMU/1zeWEQruX5K37PIz6ZZwP9xJ
b/r2uieLXX015kVQPm7/P4biNwmDT7xx1BMGAEB5318/74YhyOKdi4xqfjwvZqbz
yoOZoGnGt0bZ76rTBV+cWZUhfwkeC7yWHer6eOrbeTOfcT5+AVRYe1DmAH85hRZY
8XWcVPxXbKEaYj2jFcnRp2SD3zr+mxp3ugGfLkpW3jebGjToXgevcAexnm5dIwkT
ESxj/7NST5MW3CHrHEPjzUSU7VYaT0wkiARz04/ngOMWWiVpHpKpkTI40NwaWEll
js3ZiWlgcdVYtA+TQpsteUZtoSEHxZKZl4qc/j8X6jiey6mrRP41dYT1qjS92ne0
csSi9n9yyat86zAgZehRzPYRHn7iR1fd49U2fHsOB4e9BWNxV0GncQLxcd2Ar921
YfxPejkmzf8Uc+ITM6H/uJuT0ozo0v0s0bJuYj4Ypb5mAyPIuSt+hZ62m+K4WHjl
vmRvKcdpwgsb5WQBE+eVcqg6gH6oaZ6E4z7mw4MHmCHZwAgNKUNTnJMxieM9P20C
wof57LZp++X6ROXjgd9MHJrrW4UWAx2hMMLdGkSqmSgJqj9TJiab3tlFQ7g9T2Ye
rYn/R2nCBq+qq4OfcXYK933qygp5bko3cU4mkt3BeIvvaHfcMxW4JDSlYWpFFb25
PbCL9dgnljw4KjMyhaqVGLTQ9rBDYE3a9c1LwVqnQ8tk71KB34NWJ5S54BChgKVg
/pcQMoiKVFqpyswHiIxbUj/Pf1sKNoa8ZKCBCfZXMTo6UkBd9VR3ZbXaI4i83Vzb
6TRbu3+SRrVOwZ1O93gNguQJnUZiUimy9WU4AaQX8uWqZHHKyfeyaOVifraXUG7u
3rKUAXRYR8L+cUL9TzwPVtMeAUMpPzgDoFvAzwpW6Osq+KHs4xG9OPUg1RH9NMtq
lopEsIJPj1GyI7rPiaYLbZU7hWnonbj15Se8S1ZvK2LQwO9IDf/QQ3DJ/7NSpz2x
Pjs139kmOiAOTP7rrhNaYr0EA0c1eF3DnF6XZ7g/QGe6sJWAOWgSRVtHkDqWIJXc
EZYhIluKtuUQ/QSjpQNULfookcNcX8RAZa1HEeHutXjpeOM+PKwboOjDBdLV9BPG
stb7i24vcBGbjaqaJbzHDx5DY0vO7pv2aVbw+n20Nz61hCwW/B4Dj5d6qYhbkypz
eJeN0LZ0irT6unrBUTSODbMVxB8L3ulxDBhbYJ1dGBd06U4Wgfq6i1ut9Uez0wAA
dPjwcCGrAIV04iGyp1xM/fEjxD9P1r3CgbYMqXKh3kf6wiO6gfL66Z0d8Ony3wJZ
ELmQJCJyeIAR/aE/xSRzSjDCPIpse3ET8eG86dnEehp+o3IgW6ePLLrAXgQrc5qU
ssgTOXV4UOddSVvCKzTLlW247YJMIUlOChrZVGRYwZGUwxLbI6KfPt9RdgUiBCIK
mLUUdcGsGL+H7bvDSmoP8J4CrnWew8omB+Nds/wSpK3u3K5VQD6IONdOtwsZ+Xwu
idHbrnmZhJSQe9HtSeaAEHQV3EmFwdDAVDj0shrmStgDBz0IOWZxXOO25QxyfFNO
u2/6fDZJDriqCkYgkLkDEyrvQKhDcQ/I0A0s1pV75/e9+Nt9TyoQuRiVERyxd4uL
0gNs6fwie/XhDtaqPx4dIueIOFjPPZSsO//6PE3YMQ5LKtztUztZyMXzWv+lZ21p
TT8cwlr0VFYnaqdNlNhS6qT2AEV/6C7mgUOlYpTkOK1IlosCBYqKdCb5tGafGhcn
vrmLpzAZ4Um6xgH8FMOxxlS0G40jlzsmVtzNNsJfDYGKjgAbGaVgG3phgZ6hw3TF
ktw/H5e+2XHoFLZL8Ib+gWkAXu1YEJxn5TxSf54zJONs/wl+2kvECEB5PJvzAPfp
xcr5uGVUKf8RLx7Xw4ezWxcSk0j8JidwblYyZhpMkHBrW2zCAzi0NVBTvzd8o1kI
tls1yIp30AnjAZZejYqVZffrmHPWw9TLmtbmMHuWLA3jMRnkz70rLo9zP5UcMjLX
wzqZGQTeJIun9XcB+fhrpe1Fd/lxlqswyAsbrhyrLLoS0SKUZHbxcZX26tB+U4D0
lncDzBxeqExF8bI+oTx71/LXOzZhky68vD7rb1wMmjbbJUqes2/sHmSoeAIZToge
Grvmvu9QmGLswG4fAy4a+RQV7eZbOuuZLSifinlQ99oweViBIZTj0ddUIiIdrDF1
6Lvi4ZXHN4TWCK3ibvkzJNmNQOSiqTNAS5EodqiKhrWlqa/hmPC2oHua4MOhXoeK
QgiFn338g0B0B7iyuk+5uREcIKHHS+jYrwJ1IqH9YcEp0Nnr/3a6sqh+/yDStFGO
51ylNzo85gzt70lxeAZh9HOD2J7Zbb5zRuwd2sQnqwH/4H3n6n5VfUdDZMpdYZxT
GKDCxtPBA4ieIVx1Un7T/7gCqrK8xW/UPfSJFBK558sM59Q/USS5uWYHXTnbJLTU
DPafwrFE1sH3W68yevsYm2NC8haJlcwXewb2QzIOP3oJ39gLNZVsNhv55IMskYFl
5EXEpVCwKY1QFkWy6c4m87z92UbZ29BifYmyvV6yZn+Lwb7c3hAnSVsRQY21yMRH
s77U7oKpw2eKtYkQuDUW35AAh5Fl3N7+UlpkpvFxrwQvhYXmDmFSqSe+vk5lGyRD
FYTT+xf+RZX2bkSb+ZVJ910KGLO5M/ynrzvwG0pi8aftVQ8Qz2RYaMMBqhUNjTQ0
qW84VU7qnvAVSpgq4zBBaw/9/can9zAswW6IgekSrRtdeteX6OKjB8Zu8gTUQj/2
Vxp5n7tF5xtrv0v/Ec2CpKxzAqHoqSn9sUijPGVEijWBom8K0L2n3sTXabr/c6yR
g9y6MJ60kyRiiNs0k4W9H0tzqfo1L9UVBvy68o8qqXqfPkShREf2WLFk8qSC2wsU
O+zGd1k+S5wFVfsHstYB6Izt3ebqj49klCG0ZUyGtRJLcZ7UFRVn04lMPyaCbjS8
Pc653g/umjUWAJRfLGa4lRpwnIupB2btffyRCS3RnO1Tk8t3Pdz1tv3qLeRi/VQr
iJUcsw+kWq3NxyUbsRspnXngUGZaRF/PFDR7FAQl/E32RnPWV97FtscE48PCZ3KC
zCF1nA805i9D2zKCoHs70aIc/k4L+3Ge/YDBHY4gopI71brZcf9RrVLdHq4/lj67
Phua/JOS32g4rkTkrPuVG4fboOwtkf5yoRTqjcfyRjbR5EBo+bfq+Y6WUZ7Z4axh
rLIb6iI9lO9NL7PQ9u7bfgmeR+vMXBus6IiVEUKLJrp2GeHWQv8DoN2LwBhBVHIo
tII+KH0CCI7ijJ6i9Mv8Hz+JVQgHVVDpuscRTfJeichu4gRIrnceY/5kG4z6Ba+N
QZVfAGsJCs6gpcgS+iHd8+6KdFtO44WnEuCFA/DBQq0LA22kkEa/m6RKduSCKZnT
1mnqqDfbuUnkQrBMa/qBbjzdgKp8dXHCmQGoaShFRGj1R0jm+BzB7kUh/kukvpDn
BPip9ulOGxrK8e0njHwpRUhYnrNVoqzsWtCM+YRcGHY5J0wfiicI9QF8Oyp20MQJ
vUh0fMgjv6Jy6wxtRJ0IxuLuIDCfUi4dOnVsxrHyItrFlXhtM1JnNfN1k6uxPTzT
69Z5JxQc0Kww+Tk809TeEC5W65tQKM01YNdojkTh+vhb4qVY0c0bxwtFJuwxztYC
qxpQqVw4Q9n8nZRkQzSK7vztPcHWkBq2Hs0/mcNCsrTqFgvgZawjNcdfPd+CA+ck
Wxogq/gmFcwt8knKgy9nZNIWmG5IfMSIc472ubbROh5miQsO6zXi23ggEb62DoKH
tZKneTcL6zCa8rtJSLCmd9T9UbtPVGudEc1BlP9xIb0JG+0RCFxIr5vb6Gs+BHDt
nrvRE5MeXc4a5h8sbDe5WnHv0ywkDJwn0TxuvGhwH+C9P97X3xc26fzDEWuruDIU
xF1pHGFkACTtwctX9xHUROqSwBFYvnxEWOrgtv6s01vq8E2pGWiJdC6CaYqvYUgG
sQ/F45o1ot8ZeeDIj4+JzxDJ7wYwUDPC56G6dpLXr8tBQr5OvEsOEOQvG5fhSx1u
My66uFMkqTQiKAJ4J0Y+um5pi9+N/UivcCI9oKPZPTNXeAPkw2psUg0Xl4hd+z1w
uGRjMm2XslwbkosRMorCQPTQTgjYmo+yy4QGJua49yp5LTvMmvlPIV5SJHToQnve
z8fCPiQQj856s8tUNfywDUaxPYnfcr7QZ027e4eigzaQOLgqrj9MLWo4LJbbqNDX
zblzpKLDeKkoIBhvB8H+UwgEy3reqGXOrXsXJVvnz9j+lNLz2JqP3RGiJcg+1RHG
YkpqiSG3Oy8QnoYOpapFydlz/VDHVr3TyWI+/vx9v0qXbRWlQ4TPIGTjY5fPFxt1
QixMtX5b/Rh+Y/pf825Z6BOFwk8L2B+b0lhMpaJnO9bmmFDinCi2y4xycWPfsl3s
Rjbssvk0uybdPQORes0liyKAZLR8FBr/FPQr1HUu8+4m8z5omC25PCtc+Qkjko4l
HR6d5KNxD5qzN0dGx9yzClZOBOmbiOYlw0WoVwsQ1L3gqgaqVJHRD7xzkDXeRyFl
En5CKK12pLDLDyH6OOybz39UT/Nlppujjs7lhrXgdKGsHaLgybAfQEkiJ4SQS8Lp
QoxND+S57tSCWKhc2YpEgYuXqTuVad3DBNBkUAyZG4lQaf8+s6OU5pJyakp8JXTq
Tg+ZDtIaW5qfJLSonIr+sDEb+W6O5lScmrfZ5Q7emHORtnz8P8bW9dkcLf9Aq8Cf
e2PdZ61EerpSEYbXyrCx2dUOsjhgUAD6rOmHPYltE5OFSB+rx7kyRqzfVsi0QBcq
jMSpqyPrgO19yMdxikvzJU7kxdkhC1Pmtybfoc1SBB36wMjcFmkhNRSBaFMCcMAu
MvbuFXnbY3XHJBDZvxH2nqh2SqzugZPd/BxuWg4picc5dl8bSzxf8d3jOKTfZlNP
XwJ0XcWJ+Genu4SKa12tfi1TgBCuotJbgtmN1hmuln0DVbdcPcQpNt+rf+RQAeI2
YDeZ90anBh/clhOOAu1mLI+CbsK+SVA0ebCoYenncbTiDd4AUhvrrGniLlJB0LtH
Xmk9184+TSd7GLv+TFHg/97rkAv87PNFFEWKaZ6+T5qYTjbpgR/UnPQl9R4KENeA
y2sTzKisrAKhINAebBG7m1RAc5XLr+jCdy8nHi2hNoJqFHMtIf8JKzO3DdXl9QNb
xd4FhRaX7TvQOIbd+8hBYuT8dwh1HdGtzodP0h1F6wVfYSZmPqYVvISQAh0HNX8Z
kVlcJp0fWv3ZMNbqCZg4XO/u8Y7t3QBd83hkuqKUl3sa8e3hm5xbJzbaslofm5El
TnpWGjHC+8rBiYEBbExZvLod9apOqiWZir2RMhw5rSTL44hkE2NnVCOxECUHwggK
hrBNkAFavfGFIx3aq73baXwISYfTyMJeYL/4+ImZkVxddYV9hQuIhpgemOz6RAxJ
kDqWK3sDV6KET8QEJ7ycOW8HLYrDQ9RKx6IP7Y1q8qmHwC0Jka83JB0zZzH8ZFf3
U2aT/oA9Nh7AxvzkiCWz980yGHFzgnT4fPbUMpOKHV80CCME/LjBrO+rBlZSVwBf
of7cb1YUXoeBrfVZWedHct85IAdAeczO+eltRGdzAhVKImnBD/wghCdToMECMkLG
gXSLH815VWrRCQf4UQgaKrd48QzoS+ByFcRgFW5jkykO9hoCoWcCScrDyeJadDer
Nx968ud4K8e7FOBGYf/Qa0GvPysSSh72nttVi3LydUJiOQp6RERSk/jz5iHSHrSP
1DJ2FkDgFz507ciUz1N9NqUibOfNtXmqBq0Cx1sMvFJTfMaiSNrsMyu8N2EuSM1x
Dwh3tk8e5TSGnRlIjos40OiJ8unIo2Qogj5Ny2PYfg3OVlGW4s1EKPJSjzCx/Kf6
r8kl5Zplk689Z4hvlRzgZcEzjgoxahtMl9S08WAEhQqSGg4PfjOt/jdbCQF7URac
57r128oxp5zDM5QECgRXk6Z2GcSvnB3Tyqx5hZabnKTBMsqj5RojwNIDy40+zapj
QnJL7hOmI33KnUkgxtLrOJX4SvJtomM6ctzrT4kSEvm/YmYTgEI9Ep5SP284J8f7
FPzBpj9yL5eTDhxvu5++xdN0uOY/bdsIleN+VkoAt5l2OVJdijb7aLSYotny4P16
c5RPFWO3+QCEMaXg9i3XZlIZt5C5xeXnKpRYM61lUQNRBBvyzOqusfoOLDLxaNgR
0dhM/EsTJbFIqh1xqmVOKX8L4C+j6ufimxbHB0dy9Ok3ya1elqkHxd4FSimw8/rY
z2nJ3sXAKkcJ7QRH9PiV8j39bIYltgHJsbSWVW3JpALadxKN8oZh8V688knUoBSr
zhGz7aZaenMWDRufGfWD2iXeq0XzYc3ABMcaJLE2J40Nm+y+4ox0Ode2I7nUC2CA
xTFCyqE2cwY3wwEWc7YMV2Cj1nUKvmiJQvqFvxnWsS55MJwTsXyM6sGBx+kAExtW
/Vg2uE80ZGMRGxwZxCV8NgUCWouiLu2hFYJxjRJOoUaXU7E01sjAKs9O6l7XGCaj
zSzNXBj68KyW/YY5D3TvqXtQch69h7aNhJuwAf5oodW/02o9le9Mmli+xYiAWdTN
N2/3NSqeSBQtxvcFZmUm4C8o4Zyh7lOig3+22pMIa4Fl4z4BMdVKAPR9SbCfcaGI
pbxWTZzLlMyHN0N5MTAyc30xSibl+5Agw+dlaDLZKW0HvWNtD4j0rGF9DcK1ImVo
MWIg/aEGd7lKXuoJzL/Q8m7nd2c44F0go2zAOI0y5IEZD0kL4GTSKkexLEoRfdxp
XAAiDclAc7wlOM/1yZAFmEcfOODPlN30ukdEkxoojbbRdVPKDd3Hm5fB+/ux/RMZ
CZeq9WlnnoQ7BqXUaOwTct1Mfs8wLQESi7i+6NPVJlFR7357TXrUr4IlbkKMUo+D
dz+cecLbNMa2CFMw3ZNB+h7LDsdsD6J5ZlLbXoT8UT9KAQcQdLNaodGvhV3Ji198
gXfH1U4JcaN2TuTKbpmTYR0DFyVTVd+xOJfAfoUhGCf0LPM7IEJVJI/b7VzKB4rl
N69VOiFHEV6U3f0rwLA6MZ5Uj+VhL3xyQANMWq+oIa3GZflSavz4lo/gj0RX1ooO
EEuAz3DoHpPXlOvLqT/VTSIPGMH/lCEGGqhMDylYzRWVkTKcsH29fsmv2UidLSi+
IIpwHln5XzXwoVKDVZPhAjVfPh3hDyrJTw/WTJBY4PlilSow8BTjsJRBgI4T2tKk
Mz67rv33LEG+El1Hqqz1cf7btahOhfnTsC646BhOvD5IK00x/55U6nOyzS8bU7YE
f0uhDEtEuGH77ykcC/T2UmB+hLU5TmPAsuj3X7WUqTiWxvy86CJbaxkuleWWOdm1
obJhCkQnjJVSZEoik3KzICdRqJAtMw015/H/yy8HD2QMEAt37tiAr2QhG6vngYWn
TxvqsPJvQVANjGQNW7fz2NglNhNlrl/uwoN9uuWZsKddGwsf+qj+3U0EYtocrL47
npf6hs9SjcxqNhdBO0LeyLM/2HTtIGCnhQz1+b81g7efvY75rF74jdja10J9rJK6
mCfSm25ezOxVZ74IXbVwtrfCYygnSpYRLfyYT3BvE02vh0/zORCQJjF346F8fRdW
rYx1haPOFOvZ5c8Cz4fBtd22H9arhg8lpzBN/eN/CNP6kyAancBAARayEmKu1ilb
1U4P2omPbT+q1ZyUwoBbrydStHd/uf2HPAjhczG2I6QLZpOks9kgqlkbGyTBF5fA
xslL2X0vqSwEUI1EaUjaJ9JNoOl16wT52bWsXFqVxbwAI5ylYYVyw7K/jsu7c2lc
YPogf+i5eJNbqqfW7fyXN64za01PENcANFHXYoXQROWskwNxtZLBqyE4h0ytW6s4
nIA3niquFmEoKqHTuCLWX/fhrRBl3YNWmayQHRv64d/2izWoH+15wc0zsV1FOPfc
KUgyicAcspHYgx6yYXV/U4qEjz65xK0ymNLlcmVt50Ly562vBniDtYIvmdlSnhKp
d1Xh0iDNDbruOUFLG1lQt747iCLxm6oBR4PY2co9HwCnVg6Unt7jrkd415f8ivG9
tgl+TkacM8hG9iM0d1t0VgPuYxPk/HCi4h5UUu3M+boD4UMQ2HgU95jEKM+myTDv
AgHbh7C8UQIGXZqaNg+G+yD2JtaGXE5bTCsI1BIdr/Ov9ZjuOb68RPgf9yrQfI6H
Hhc4lE3uS+M7ccv2pfH0+peB/0niwG9wOS6fzsRJQsxKwokK17AXU3LhWXYHTe/Y
NUxg0qw1+u2VC0Q+s0zD2360qJNjNhVXTAtDM1yqcsA3sdewzJFROUC2NZuIGvLM
EKXKIatmlLYlsYQO6wMjX4AZaK/EHy6L8YR3h4umHDp4xEgjGLJT5RySupWMUjNa
PQt7FFsb4gbNmBw9CPeLPlDQ6zJ8DKG00nmDnEAFITncvfT+V5RDkrJ7NIR+JfCd
OM3FmjbkE9gD0le4IeUXZO+nm/cYK+SZ3Q6Gyl715dm9bEuKfGq2k6v/zyk1kN+I
Czpn/5TZ3PvNHwBXdXpbvRAs8ktxxySyvKIEYI2QYstPSeCsECipkggOuDeo8eJr
k4UD3QF3tczU00xJs4mYofG0Lt0OUs2z84/RmhD+vrrPZtnW0893T1ZxWugbMOYf
R6cJJGchiUkFuUEiyBROklk7bBD6iGkgFcsMNIYrBqoT1XL9aZ5B8zJW0Cqs439h
icS6Vezq+E12hNK/8826b+fQ7ojC2BpaV7BrqJsm4LEVWd6cBfcHUVoO7RcYaVxN
IdcJtIaGw+PR9GKRshYVK3NAKxhTvLZQbtiwcV//AjsOut/b0ixUYzTOjihIxC+u
0Ey4B3PDn0LZLN7pvOAtLtDLsRuINW1sudZK0UVdWS/Sj4jPXWiELyWkqppF89Ms
FB8GqfgeUl+mC6Q/A2Zxogju90kEf21t5sCTmRiYnJ/2W6igKn9aN0fLDgGMx1an
ms0/I+wXdUzpMTR1UHgkJJ1po87A5ms0VsuugarmJa9ITpAALwtdItNJu1ghQc7y
tCPpa/mNdm4MB+ltXrdYsNlkqszelEpYWRWuvsJcOLujYyjPAmtUi1NvwQxhneSW
Qm9bNWvB56Twsr6/5FmE7QURVasGd4HBTRNajCZ36LdmucdP0vbzHdggoNbZtSip
aMFlaokQU7m0SX/PMxUb+P4ajRBi65QpFbuHHeaMWZ7mjRJV2x7ZT9cmpWzYvq1b
/WoNJzdDO0EPsuTOnQmVAzbSHdpb59oPsxbtChynQ8Q2vZaLi+n1S/nxwJMn3630
jYigBtvXjsUAuwzsBr/EdDFotECkcWo1G5EpMPHw+ARiJkr+D6xIGUxcc2qHK5vN
BI6v3AKUSMezxKuAnelur3KEN1l4Ugs6A51DiMZXlkA5n3s3+Tt9v+469//3ozRg
BubjfdkvnjB46liG78uqtJQQ/oLOQcQq6uIuns0e5SPlwYp69svg8ZCURJqJxId3
l6IL9MrvpOOZYTehlPSWXMmbT3nD1abrcSINeHnuYVCR6go9oUEMY+L8KWXUGR9v
k+TzXRy20govpnv3Jg8fTArls3RcUhRpdfBKbwrdkQBSPX2ONkTj3TrjsclDUrKT
IFpWgkaEOSD//u1SQrY6y+ZztJh2a9k74leIFPkEd9zr0hv4asjyztbx5On3Jyrz
uVQ8oqeYNUDRvaZ07p7UxBwPLcGcw4Luy1K9d1ds1Ek6Mw/qrTFwsg8OXxJ5gU1n
4Ba5KWwa7Lnvj8wPcqJov6fsWh7xsoJb20yC41YHQ8NMH1+6wMFUD+NE3SxHpKNT
ZYRIN3rNEl1q55xeyldjgB2vL5KskSkrrxYG1mvsvw/1iIH4iwg4d994jDedfDef
ZXZGrlfTR+SyA4nCHBAewNSVOPDWf5+30t1UBFmYkCXrke4Zxi/jC75iUEwCEX1+
eH7g5ZK6TnTTBqmfHBfrFYFxHsE1tjAqRC6DFo/Fl4YcGSVLK2I0vsQhX/w0DR0H
BbCgrZDD3poEZCe7nMFP8BlvgQkkybgbvTu3sa1YuKWUjnIwPO6tF+vCvxqPznuD
+98/RYvbFtxGEfpcvPVvpwL/0qkseLmtRbv4xbAdOjrL/azXTrqzt4qPlGmxKIYb
nbIqAgJQlqjVl66BYPkrdcGv1qfmz19A1naKChkjfNISZmJv8CwqYIDwPnhgRHMj
AcnQFMkAAbHuafGBmvn40gV8jntI5MV0/L7r0eDZsglIY9ocl+ZCwgmfPqSkWnys
Bx9Ukh5lbJBftTZh7aYRUVI8tC1dpqkdRYgnXuWgF1QPRuh8xFnApbi+G+54eGf7
3Rptg6g/sGI5kTIQXjKg1lRZOpEXAGDueMMqL/fqmdzMe4m9jKp7SAR1/HIAXkTd
N1dwLu840j2ITTDFK3gngf1PgtPcdc/IVDYWzhYG784hPDH/3PAWqqaHAV3Dp66y
IN03d6qvvPS8yzZES+s3i5jXcKWQ9wAut9mvLxZrcBDZi2hMQFbC9sXJKfVkc1iM
1Z/2xASp/71tc8FcHBgRSZYnhKSLkaw/h7uBuN3qBDihJSWukyhvom/qmTqwF8Ks
hC4QZ+xh1k1U06OwTQjzAGqrtNZqFM+pqqnGgYjUNu+TlS2M66dt9zzrMWuTQuDA
+CV29cnIuKVPLEGnH4eY8wVyHjUC4UlOXKyXJ4v+7m+YlxDh+NDxobo/eVWGoy8/
jl0DWyehEKDV7TRR/k5iCoEeUwUUCQ3//Uk+1pa960bLe5q2BC0dyLloc1NDp+Y3
VmJv5vQDyhjhc+a6oVG5EpoivQeBxTEkGR1Dv/fBP8bku+t4VDvSQMnobQbDRZPI
2U7lpS44SjfHqUQTuHIiq+32VOhJPeN/MTleMfjNV0BcEjrswLntisAdF0JqQTKZ
W/iRjj1Fw2aT3Unpgw9Gj5QpkYiQY7e/7Q4zKZY+9VSz1CmwDlcB/lN1f9BWCoNN
boaDuRAoPtKpqAdbYH59x52AipSSzqEo0xXpwPk3pBTimr7wyiaIUD71jFmNIYD7
V0Nh8uQEYPMXHduoc8oS82QYtDJlzqFOtxp5P/1OHnftVBIrbHMONUvgAnUIg/qx
ArqYvAjH/WFA7FWGHdIV2nS6Kl4LhuNimMPiiYB7DbqXvFcSa28uPpQfFqSGjqHl
zHdmPY1hF93qTbl+4xNJKcbdnNPH9RqkNFLpiXz8wg7bvkaaP/z796AUMZeUW7v/
xvYC82+bF13HDbLA048jQkiCv4rqarPWOj0jmzss5s3tPSMMrVffbOJGkYxqcvn6
SxWu1ksqrLSFrvI2GTcuRjAQ3/ohGmrA7OcmeBDpCCJPX/dMCf5PBzmMroLy7U3u
suJWA8Wn4H06o00JKF3ySzaB6HlnIy3TTT/zM8pBq9v+6iNxgbSS5/rKiJrTCexy
dd/k8JF9TzQOXs412HZVVDBSiw3f4mJaHscvn40+mrMZ5uX84wUuWdfQbXsCF71A
HwrPuiGeRpZcuHmeeuRK3490yfNqhAmHfF/eIQSxUZJ5BqbMiEWyR7nv2AFOlIRs
Cm06V4LkMXSMYRFAjDY+Oj1l2knjwseqiiffhfTQPx166u/i3qhY5d6jAqEM/zw9
PJihV2nuw1E31QzUjeay9Xeb+Xx0b5uUXWwX1qsCgs2H/ILlBP4NmWamXi/2WW5+
sgQq27ciDUSGiB/XqtG9h+wogGq/L0tQg9HVDIefh6wu9FvZ3wHv37z8ChMpHq0c
e2JpPU7E0pHgfqwOva27Pe0r/m7W/TA3OBhsriVSSfTcV/wcD5SVWX4qCXxzoUSO
v/WuK1dkO9Aoyq+6sLb8ioR+xTweCXj1cwwiNXMAoRXA/jSVusEZ5H/xxrPfy1bg
9SrGiVbZgf/nNVeIlE3kNkW0I4ZRkqG5GrD04JC9pC7rigroiDt3rAr6D05fLU3b
MX7k0z191RljtKzn4fe6vMOS5agoAe2uTk4Z4MOME668aGeFsP2txx7eHKDk2BXW
QwT4PsJ7LRgg4ZY0KjoJOAK+/mIheJgPQDlndx+XWjNNpF8n3Cy/Zg5L0LeH84WQ
5QAxXTP3N5NoUmgY0TqscrvdZjigwxIMu0R/zzq+vFWKZWem7BX/AdvwSIFqZJpq
ltGt68VhaR5vwbFT3k9llr130mdkevZwxntwIMGLaB8aRIJTyZZOzFQbUOyJmQ70
6EfPYPDsBV04eN0cSwbkFO4eCc1iKyL6GpAh/Lmujuq8i/WhU6KINUfYoqDcXlnF
ZwW/FJJDeElH/tPROw8M/7c338oVkcz5HkHOYm3qWzTfNt9CRCP16Vmx8z0D7GfO
fRreVjGf5+Gm7NXG836kReniVsTvWhotOYTNAOkovs6L3CEw9/Bp1r7vIADQVP7S
NnNgvJ5+dNU0/eyTr04EqsJWuMpSw/S405tPVuz6tMYkYg2f93gX/noiyYimc/iu
874K4MDAHS7jO7Yn1dlyUcvNt/JX1yb/0PEQp2AcQ380meGeFcs5pjHSPszqid7L
sPnoK97hxQVTBXbvINgGWI2ncYyRGDkCFl1dSexBoh+2FC/vgreCDiP/kCOMq15H
GKGQL6Y6DZAM6FK9qlZB6dIXwhcSM5PcF9POP5yd4wcN8dPlFyjg4aosXbvKnUQh
15miwHhhnVbsDh88yoW4U8svD0SdBYUG/4wpZ5aRnl7nPQDqQuE0cXQoAGGvX0VN
P69+fbnrulK9E9K0Hm0/qAiC4/EYxjf1vmmuX6ygx72E8vtwx4/068xnVFYq37h+
aHNWfX1Mp8ocIoO8OQ42heGffuGbfjetdrbJL4q/UDB9/CLLKD4aOkwrfvWVBQh2
rlPdNKAq82NlD1pYgpN+Dz9AWcZ+PQMCmquRIz/FBvgJeQmwV2T+uq6wt3NrvMqs
yRbhbVGhyr039MmIeqxXWo8efHPqamPBT2cIjeT0Ft11qVnP+qfnf6/Af/X2Xuxb
YVNYTZyIxxkBwZ4+rHZBoyswwDfiuCr1vZ32rZyMqmVY4Qw/jwK1FkiSBEPsK4PW
TAqzByQjtFLSmmadpXTCOz3JgoRl1fRBGj+0faJGKsJuJYX7TkJOlLmuRDZbB675
plQuJYMwMd82BEZ++awmO96f0yzDeVAZ1Hk48ychazw5sCorcyDMKQs5QDaYx68J
U4vDHgP2S1KAmVkIds6YOOCscSEwm6VBDbj40yf89+rcaghzszvQ69peVsOvnl1O
CqdciXWqIdoVklK614cQgL8sjfVGYLHOjb7/b8gOikvhr2RulVL0ZClfxHYZWo8Q
Bsoav8IrZKGwvfyDPdaY2e7EXejX90VtHq9WcBKn6vs7KZOlQ/8OLcYBkkTfOna0
Q17PbRcZvnw0VB9vVB3DW+LSUPEEgdXGSiOMj42fytpdd0cqmNNwZgt5i3pZ1LHQ
V8IYbRJKWQLgoqSM7+6nbs0bSwYcObcyqfJ8WeBjMiOeMDpTpl+ENlNwCtYkGoQE
Mk17yG9ZRCOpr/f9njac9j13D1rxTePoRG+Fw76zFj0MnAuuSXcIcHEPMiXYbs2u
aEXFOl+DHo7k/VSjLUDR7X9ckYph6ixY6g5mjX975yjf3q0WZub4V4Br4jXivGHc
9oKJoO5VkASRXHoYVJWUzO2jZExFjCDRJFlGjQI/v5QBucpEx7xb3L25iiY1xghi
XgIoATxSuVHswNkGvg1MBUp2tMVzI7byJt7CwRyV92xRgM/aTe7ZWGJefVU4FFdR
t/5Oa00JW6jbQ7c59qwLROdRkq693+lsLjWBrS1LaP8yTID9UpnH3Y+GlJ4fKliz
1CIQMB/+zE2pyWm/VS3ZRaH31Vlahkhn8zdeQrwG1oPaQIo3u40TpYFJovHhpKA6
H1EgjaqKYqSBvaE6YaMUWW1r4xV4uZZTPeug2qMtk8FYM7RrUBhuihVa7YOYvDNU
Uav5SH1YcJphooIrvCV83paejdufJp5FozuLHV2QQIboLfyUhTbzU85f1AZuZ3M3
aiQIsRychm+qLV6yKSYkHDif6CmhJW70fJGPtROvi3rsV5PWH5DUUaPa9gob6c+m
AgYCY1sJMr5YcPHOhr4E9vMI8nuFkliRiEXh8Wt4flBfD3C+muNTov5KnCxJmZwe
mlF9njZdqQsAe7B+78rUdM6BTj+YMoR5+llP3BSUnML5WXJH4DdDkbqBewCGvCC0
68rKTX8ViysDHV2FoNSsw2c+9IwDSMS0JrZZImAqG1K8vPjRynD+55F97jiEQHBB
d7XKLkqV9oth5XlNEV0KXMsg4h1T0ODoKoDv9hbziOHNyY2Cv+SkAIUnzuVN1HEa
2x47ccfpo1HNU3qcJrtll7wJoXTgciljlRjNAgNbGDxjhgFcYsl5HM3JLW7XTtFH
dSR822D3F9zKy0HCeNz5nYtRj+668LaHezh8qVgEd5FUrZZWfQKT+TQcojisFPNo
pDt7l9p4LznaAwdeTm904vQXfSnEKEEbC3FO5INAzMm08w+DfezUbLljRe558HRj
ORo2ysDWCA87DNA5wS8EKOSogCsj/fjCnLsRoQMm5hvm68luhopzsKcGBjNenEdf
vWcJX0TkUR+AKI4fUa33SzeNJFi0yGIs131MQg1IKpheoHapwZdRsU3fZ30bdfgk
utqghgyTvju9Bg6UlO9gxiA0QlCTsA8+aiOrNTKF8qsplPcIDafus+6NvdqXPJX9
ywslkxT4nMEALEREi997su8A7i/6tOYA2XxRHtX/2+xrESS6hgWvH7yTshAaXdkl
dEhPqtmVqoW/syUaBhX6e0XP9RPhtsTZ8Imi7T3iRaB5kSLfhPccAJokE75t/Rpe
UxZaGU9ir6ts3lNzngWixufbbcdISfqRDeJg1y0kX7vQf+U+SEQpr/003f+GvuUB
b+GlxyGxW1U8Ylcnn5EcefxFGNI+ZaspyAPRGsyHFL0iqTO8B5gVnUseauw2pApz
I4Y65b2JXyRxQVbN5Artu5SI5j4kYl1t41x/UtBRH3SjXmFduhI2+sysDZq6E9ct
+5oBRPZifagsbaO93yc8v03pCtu8l0XF298gpHGgqJBr7Y7qt68+TZPS+hCypVqd
3yMIWmEad1nPO1WEAMiib0Nm+U4oc7rdhvmLsNOfqigwlOoeTVT3ZSiPWZaumvWB
2qB1Df8mcbCreZ3hKv/EHPVdJ5KitojQFdryARtqRHn1Hwg3UeyZcNmoOl51WzhK
aXfvT92LL/meL668gNzPXsT2DjbZSMU4NPoFZDx8GfyWYR4nzNA7rPLTbsTeUrQ0
AuKScNsZ9zXkJdYL5zciqXeEi91EcQoUEJFGOuI7htjEBuxKs8V8KzglbHvujrQ8
FSkZJoIDEGNpA7xLecE/HIsEtuwsxYr9PgIvqmVUMqrg6KEjif9KGEWpTwv50PSb
HNP9k+NK9hAuJdlro93sF+jGyocAMS8lsegxksbwgS6ZNVD/Mw75lsQV5fvCaSEH
HN2yphQ8BJVrcFCpnymq5XiTlrBb+cLsbZkC8jXfS9tJPaKaOwTittTaEw0OmKeq
iAsOOWhuvA6beY2nfu27QJCvr6WCd5z1nIbHT6fAbjYo8Yjdbg16D7hg4lxyB4uL
7tqUPcRDoX28nf9vMKzMAZhF9p0F5duHc60WsM3IUscMSgX46xxPAYB56BsaWaPv
WtK/7FHGigwBCZ1NsFVZfFi3MdjFw6lcl47QAhfXNNJjdVhPkT5XpYH97M5UNOiy
jjcuNMBwic+/twjQ9akpf1m8qBC9yA/Dk2Jy4edb1Tgpn3iLi8V+YmoeFbcOqVCb
CeksimT7QaGJ+AYmntz275ZrHJOX1DCyA48V5B2oVZ0HCJ/pQMsy4Xtfi/cx7TA+
tlMYjtxZg2zOAoPZXcuFXC9V259VUrxaifD7UaIcZqp6reZNB9Y9y/Fh4HSDYmOW
+3gdlitr8P7ICtC3DA8V+bO9l24aeWeGmj4VyrqrkWwP/gP8iOFV4uQxjNszNEjB
+iWhKJ0osjtQnjNM2S7WO64m7O4wvqpIFWaelvbvyl5m93nvmNbh3npuql3U7ohO
nE843p7z7kyKMVRAygs2jIBmIuOsIx2gUM+eLK3jL3f08dsZ1YlG93PWkPcli1Tn
JW1viI1OjeHAeg9PofcIT9OHpJHjTlhUoGo1UfAxiFqkPfD3vVw+oiozPo+l2o5l
df1FlE7etQ8C5bGoi4+gIzdZj5eC2hlPTMtBx7WKIEJUK9j/zcKOrrn701YfEl7z
jCyDASF0EbrH5rcDVP6JSZydbmxSEG6Od+KxAXhQ+DTQ2RKOBLwaRKaXeW4xfZus
txt/byNNCTb7Op2vt9937T86H4pxuMnfj07PtAKCzCY7pDxcI9vKCImpVS8UOdU+
PW/THFkyYAs0uBFIseZfDHxVE22JyGFQZkyamWqq5PvSnI9NDyMVTKWbF+RgMdYm
ptZfUiIs12l02AaDFB6e6dc1AvNPdIsx+kf6or3GpSSOYw5rV8qkf0XYCg3Loz2F
lNE1VadyPGm28G1Ixtb3otVzXytp8oLWqVjA4+Cw1/hQtz46/VKZ36ikRAIF9qKS
En82jKm6VF34xNKWr0mkX822YGd4eILzu3QiRQ4LYVcWpXo0TLsShwmhqyDllt4K
NIFxlDib2GKtTZhjlp17VDiu7gkBGDlSlfnMFdvfz55O9Itu2oR/LdA39hiCGNga
GsmnE+ltJNNjrn3RfUok7ukkM1oMet/Woc/nzfY3NgnAs6zwsPhwhgKeMrgxrefm
+gIqCGALrFCr6DVnnp/EvBjH6xvSXrHEDuqy9s7gKgBLJicKXDGeUbfuJvSDqkTd
wn8hQpgsbYP+9Kb3sBRY+vck6DzsiphRFn1MLJajbOl3w9bkHViSOUDe0mCcEjsV
dZXx2yH61E/lxzmiBnW+dUEdJ+A5mBdyzAdc4tVxWtJrgIriljya/WDpS5Mtx0r9
WccjGoEb+Gi8YI8Qe3C6DVrBQJ37ELlv+nAbFmSuEzXqHmYfGyVRYSiE0YXKAnm9
tkMK8qN6tjAhXsbXjWZ5tKBl+ZXSkXjcWcDXCkymzsslMSEvmjpOGz54b3Hrk0tz
OWBJYXr9cxF7XyS44BxQida3wuZ6SLPw6jwpe+77l8Uenu9vqc8vM+oJkZr8Tgly
5j7MeVMckb5bhgd4f4qdr2f/296S+g+RIV5sB9Wd9QOXxJvhG2e5MoFyPCifY6ng
gFE+pL3JZzwutAqw0/qmtJPqMlZ13QAKEpXnKjEGRxbIvI55jSNMFMCx8LPDFupM
j054MiMmtjO1VGs4RZVZFubrGmlJ+vu/3dretJH2nuAYhPCuaXVsJplsZ/AFXZk9
kqgrBwFgrCAbiQl4s6RrLNDFhVOjzYjfVTlBpBhXeNfumuYjD5HKFAkV0AB5uJ+Y
OOOtXKjvpFAI1pyvkPrYjjgnMWYZw1jFUJ0fXZAy9msYDtxx5fhzsIIy0fVw61EU
lZ2NWmIomRixYeotaz1izpzCKhu8nw/SHkTSG5YQsA99BYm+OOQEsrpo/KI1wA6z
mHzbsuneB09GmvTRYwfK8mKG55lWs09yfFfAWgUniHcHhzR66l8mxVzSFuUmfApq
6+RfOKVUT+6Kvj0PBkB1ZMIl9UZ7O2mhSZP/Lymm/EI5jsFCuUmxZUbD2hVRG2zj
Cl5YBDs4EzDT7CE0WBWVlJYFbNSQGDFIg0QIbiBI0MZXT1NhwXFMxyv0dXadx2BO
oqmFqkbJ6SgEbCRthED0aONOJ1WyNYutlja1u1UeMqGZt4xK+CZ4sO4/x27q+r4a
gp3TQ4OFVxGdSr0SpPE4ss8jNYS6OZDV2+tpbAoRESnndla/jh1sJmxT1iHNe0wp
NgK6ayCkjzVhI78Yp62KE8sosY9ynyM5m+0YRHnmm1jWjpnBpXMrlxEQzfufi1PF
s1EaXmxzxpKYf7TzjryzIIcNYxsjeZs1IifmhaBjsO41U6q3MqeV/cEh+ttNzCJ0
e96JRJ5dLhdNkDRpO9VOOouQxvvRHtLf508Ex2O4om+2qTBvgW+lIAf44qLcAcxn
MFaz09C91Fly0f/bp8LY84c8cG6OkdjdB9Priwl4H/LxVEBszX/8rTtOtM8Ne/pG
4KE0x7GIIL2wflyjZNDmZjzOwBqlYu/MjCZTRvpWY179sMUsrO1/PBcy0towPrqf
D6Nw07i3QNtzJU0DxszCCgQpI782z1/nsobE1KR4HP076nN8sbsoXxn54ggHw8UQ
/trDOVak1tL+IZoZsiqHXMjf6tUSFUO6k4cBrao0ySb5wT2IewTuQNSzj4qz/MPv
F8qrf1GTXpm5i+m4GalEagHqRqSejYqvT+TQ3NL/UEEDeJOebe00FRRAZHIQ2fGx
i6ImkYLHyhZWu9rfUzYPyaC/QZXS7MErcR6kW8J8lqPI/bjatu5ZbEuSo2zk8LOR
r+PoTevmb/cG2YeJS2VvOVPVCvRtxGv3xDuKXkYuQFrZnZqcliPFlY24GS01bXgb
SppWhP6Z/iakNt81XXrzBPpVsT3aLOsiv7/4rOrLN1UyP/U0WGVOgBmzRSGhaYGZ
Qou9VXXA1v8dGuW8XQbTB0fb2wRzYoV3yQZKXd3mBCjYKSZjcCDX49P65nZKlDLy
mA/6diYZ33BxgA02UhiCAkeMubLv3Z2Yr57zfLxY06eoKfqeXn0kixs6oXFbnbrG
Vjsek9n14C2b+uONiD1OmM4coQ5+nhAdR6FWMhJcgxJh3eu9mkKuvzpsH3VBMU0Q
+Tu3jymoIbn0XHMGJX0jQndUVWe0g1NhT3bEi9ng7EFtrR3cDb++d8mSPo9LsPxJ
EO5+JV9/Y7P3SsNam3qUIIbcO2Y+qO5SSxzoNFBoNJ8eMLudKweviQInlWqg+NGO
NUNsOM3IcIb7omtK0MOkAiZ72sffxpu4IpB0qeb2BSspMTLmmsrNeYWd5G0E2e47
OL0sFUJd+nGDOEZ5pyCa6jr7NXOIEG5Lt0z60evKEleLbb7vFo2DGJelpdVF27sa
HHnmg2Jj8zKhvRH01ReDP0QBADYV0PZDIvoWlETH3Bp5JlMLv6Ulq6VflJXMbRAh
/wr7Ibpz1EbCObY+pJDYD5WZaZcXq3cOcVqk+8Utwuaty8dBnXmQlkSb5XW46iHK
oK5xaZ/rR+SRZhuqKwKh3RvdmG6FNHaEEOom4pSMczzskUTXS3s8W+LgmcsYqDPN
tN8PtOj9eT6L+IniuieiWjLyk7vsbYZgG8clo6HUOL2L9+NM0/8uWXeTtj4xzzij
ppcQ9wKZRH3gNVns4TG4/OGfrk4AUj2huu2ewMETQbr3zjQ2+DG9tVqNuKmuclrl
k5ODauVbzmqbJ75rSJ/dkvToLxLJ1jaqQySZues40YMrSheMrRunxefb5NXhD3qQ
WBLUN3LVNmEitanQreWpXENX/aPeocVnATWTZ2nOYM77nwj3qnkVVmvwGaFeD4Nm
aQCrtwdEXJzFnibFYmvrkBHzQEodCHC6G8pc8QJxXwpUte//eRc3NAlCSlIyzf+5
f7xHz/hLS0AVFfi3R1ybtkocB5PHUzVuRxW8dlB+6thxbDbPgD2RiXsKXq32e7rm
82urz6pgF3/1eZanKDz/RIlQNP+lHHDPi9ZlhDOzl4487NSAN2GO7X9SM/g9yjyy
FxUkrE9A90s6hgHybFIMmUJ9FeiReKcU7zm9LpBR18egHDW0RnJOPWELTl3wVkcM
0XptCBwKP5nC7DgaQRy9p4VOjqjObv9/D8WcoctRVN/I4f44LWt+n9RGHTB2xLvJ
Q5B6G1NeOEHMPkgZ4nv9GB9npKLa/I3oI+u4UhtM2y9tfiZ8xpD6glk7htBIfSA6
3BBGtU/qvQIm8lVtslFIuXiUONCBcUXiQ60skL6I+w1eYtzzSNyX7h9WzHlg3sKp
WVQB2VDOqYqr1OuYahiU1toyDWHDSlcxbZOAoNfxKw2xzKe01tonTQG4mWurUFEF
XMQyiCtOlhE5HCjVYV+sjIXHYpm+uokuTtpoS/MDXifeO9cWWuBdOYmTqd7MBmeB
nBkyLoWC3eLT15mIEUyx9YCO40zWvubN5CD44vvp4H62WwPdD58bFfrkcGW4ZCcP
x21lelMcxM5rEfnAx4pQtJMFO4kZXWlAm+Aoi6mDps5PFive2RXXlJB+UQuqhte3
fhhZfaolcRwh86xvgEP+a+nRg9rCPJzbzlhQu9hkZUlNpAjGUlYx0sJlLJlzKCsy
ozhWHS1WqItB79DT8xvsMibFJ1Q0jEp09VmqGHeu3ne43dSVCRX5MRBvHBQ6iPzK
3VKZTg+ZNfW4L27pLGNfG1F7lmx6xKdADHTuD6CBBuYlP7k8v98BATuEObxaD+DG
CwXOjy1ml9YOv1pYzfxAghikq62kDYwECdXT3i29OG7zrdMbZnzWvlb6iyqGcuZJ
WV6M1RmcfBAEpIzT/3XqNxqaldaaa/sM8oJt7FLfvHviPF30u2DT2GF3I//fFhWA
3Z2pkX+43qbC7/i5RGhc4sKnKf0YpSv+YAUwoowl4wBL450KYM9lV6toLwvV9s1e
JHKO34VVYmHw25+Q4Xcl0QJuIx5R7ZPMH4hZCfH4BJa3mxPQ3soBOOt4QhrO+aa0
6J4QWn1VpR0KH0GW034j7Tc8+GIsKM4M9JhxzwY5tJSP1xmMgVkuNNjn8RlEejxE
eOiCIjMp+SP4ljBgNRT7Obc14kEoJVpoP4WKHgS94UlkEp8bUcH36YhM2VC5Q3xR
X66WSouzky6sZ1GXDnm+4r6n6dPsx1vB5WhBUeZY4W91Ldp37g1d3r6oJ7utxDVO
i0W9wCqmOH1UktW0nkOvi0FGpKjHfmDX0Op/P3GPvBpCZAIT04CopwGjkhy4D+r0
I7mgRSgk2Dh4m2wTqkzwxePxcvy8t2uMUkrHyUtq+O86hhYJjsYBTFD3GNmOn2Lf
EUkAmBSo6F8FeZuR6xQaj6DCOrT21BsLd4ispHlXR6/W1WNktBVtJlCzLmCbEo0H
0D+X6Xaot4odmk9uTNTsE3g4juv6BjQN5gibA+8OHD2yIpbBAyjzwDSnzRKypAr6
l8DXP1rcGp7N+jgIAGN4Ig4a71Tw1+WQ1oC6g+6wGrefLpPJ/4U13umDUqpHzJuI
jE2AInj1INCi2SDCaZICuCXvDzGo3MMmaep1tIeWP+lm0TvRh3n2BW8LAusZkw8t
2yfc8Tif7mTwY7pB3BnOcQ+6AUn5T66xmYT8mRofsbsb+a/kUrZd3N5BjAgq/Sou
W4GeCqTTKrSjmUOhHCYLUigAFzeTVYfqG5mARJUOP8tYsNy0M+nmXaVUUkuOBDRV
b8NiFrIAWgE+R1Kog/70NS65VSvok0jZm2coQx+SU0q6xEopMYum0aQa1jKP4eRV
IxGK7Fc4D+rjxoLICWfU4oeNixWknlJu6ybzSKBLnO46kDzSVapdPoiof+Sge0Y7
n7rmOe1vqStqoBkBvUlaYmGBmyxmdlAT1tAWmGbyleHCIww+gpSprSyG9T9OYg9a
dbv9A6l476unf1prsfTnzXIkfr5kmkgvs0OzMH3I6fbw6X5tvhdFDNJcvxu2fzwo
ALFlnK9dpzV4CIMWzEj6mlPxVwMOIk6Ithzke4bs78KwH/RGx7dza6EP/zm6XSjU
vRPdUOvv0YFT9wczUi0SjaYkeSKic9Vjr1vJkvKZxhXu0So8weCf7CUULH9QUOmQ
hTjJdMDucQtaI0/JOipaK2YM+n7+2p8QZYriLR+0kvtWV27bx8P/1jCRD4kldcC8
q0adY5DRFA1aac4R0ngUNDPh6lhwnrBupQhielpjmE+aqjtOB3flaJeFafwWm4PN
wGQenJW+W4Dq/6pV7pHS8L4FtfvWb5URbaM19cvsM94GO5YaXvR6t8odJqbUIRSW
ABKxi3+LlIDiFamdXBGBycNS4P6ec9golTdde+MsQyJMSTBUqk3RgK3/6QoeAfNa
P6UlIfT1AN+txIvG8oL3MDYwh1K0Ju2iqbcKP1z2r1x8ccD9w21d51X/UvTaOIPc
g6I/mhofwdjWBEL6uLF78ZOA70ocVB4mcS9DG9zFkCo/dVWp6exPfjsQthdkYs9/
lIvGOhtJst8Qz4oKYRyngAO6kO34M7Oqr6bcbNKodaUZUaKmuz+oYlvrvKuqFFFk
f6Bv9RtDbCUthOMst76jq4infQDFk8cYdxUuy189/IRmHYzoli80Poweh8LIn1qg
HOt967o0b+Hmtr0bxvY/kDxoTdgithPA4vhe+kTrikvi3hP6ZTYD6zq0cLfrmX2O
cX0uxEftnJ8ynKEcQAFVn8FU6SndCqlxBUHOf+SfBmWGz/vbugQ+733qHOlWd9Q9
xUK2XOPWjSsZY3BzHs+9yciq+Fqm+/FWNafIXYUsf+CATrYkoHyR22X2EugPq0Bk
9avLDiwU7JnjWsh7CqDx3Ka6MdZmljhHgmbwKHiJIXcTxsZ49JB2Z2y4Q3vCh/4k
sG9hB7Y4FJlO2rna/SGKZQYTrxb5EEzOCU3RTKv/11oa8dY3Yao3YAkNVCo4/VwF
PewXcR6f1ysfzQsbrGt5YQodF6wSsPT3pQxgRm5b0oHOkqc43a6rz8qgs1X7J1Qk
8PDVEtQZV7EqWpqXx1AlToEhdd+JLEcSLhIFbACxoymQTr0psElkxrR3DnAjzMFh
6XZOexfM++BUadxGNUaJS6IbFgtQlDddBQRxD+qB1A5oBp0uTuxCQigBfbyYNBK6
ggNzqjCHMmrk3Ppjrh3w/JkwOz2xMgTFBoEiSTg4zOg1c689kvmRPyg/wxo39qNx
dhKqtKreDag6j6idEWw1w6sDXaqWX9xzKPsbDQZmDoRpCGHVOY5SRECkEYIidEHu
XyDtBOIsN+8l4GCEI0hxB2fwy5NpymIo9iiH31hX4xkz1OgIINxCzboyE91oiMVT
wle09zjUEAmfPo9Dx6B8rPxtvYje6eoVhFm8g0+xZjer89wHLKS/i8Ph4NJEhnsE
xQv9puP2rtezpotoUu86ZERwFdMxRVRkiDpiW2CxlEFXp5xZ50ElQGpstpNmtYYB
MNGIqnUWgQ2SNZK/RVtzTch5P4EtJyP/IVoASWgqNZJxBWuQWYnXukGdYCQA6lgi
EdkFCv+s8GPlxp6CTCwG2BAlscouLIk9xdHSg6qAzN7gN6eTu4QIV3iz7qfqLK9R
70lfubjU5+KWVKpE4WVSSFUURAROYNpeJi/qESQLX37FlcC1mydSkh73xfTG+aXf
cNTD/XyG+kqeHdrKJbOrTCid8kRpkHZGJUvF+t6TrfZAQ+Ebu3AhoxKzoEdDdgCI
xoK2kFhmvSYI4Yjc29O7Lgtzn9FO/cUWIlwKfyDe27vxJ20IQrhakcAQr81KgXrn
eSGaUbUBBKZ0zh8Ts1FCLdXDZcCttMIbyTb0SeVQdYkUc02jLdMCzqhTL26LFIu+
DPba/xooh/RdP2UKBpJh0JLCf6Axs6Ho17+e7a1Qkeyq8o8M7XS3OHLZ2GqnpdhY
V/JSLoLglC8eCOJvN+puAO2b1JU4XrPkee5K4idIclTYDP6BN031Ul3+A4E4YFDi
ybCHclDRn8XIKFWsX0bhJ8wsQMO4UW9FWj82mDQwHl/6AcIL5qnNMKjY8D0mrL9S
itSF/1/BhAFXWf2xax7RFFABuKAWCLrgR9E/zzaHGsVNaNtubRmAHDd6QT1sNyN/
PGswtAptqyJt1YlmDDkcfylzqaLqlBs3IaXdjcqU9+Y9kAe1raAoY+8nsMnb0UMw
A18c3McednuATHiyNkUDUYNcQT6+pbgQaYbLj+gkkfYL6beVYE4E9X+RLb6sDab0
6DU3PNzkHfo7QMLw92DyZE/vi1dp9XHRLI63WsM3ZrO92PNiySHQksNvyyhUt60F
xPFduw9jenWMOoc6Z6nr6o3PJ2hJ5NgF6sWBqS9vgz2ziwPY4D44DZ54kXWon4OM
F1JLRo/xojLFLBgaAEL+5g8IaFv/qGKnurHUcdPAgEeKKrf4klj7FwNuvnopaLau
jUuy8uOZAHgmWwQTzZLJa+JOaZBN6FnByACG+k/JTYBZDT7AlyzpSgf/qHoyuLrD
rNlw9q1x6IglVRyexuduX++eXjv9gktUGbb6pFiw3rDHlgRkAleIkR1lHtWP3Rf2
HIEXnBJXppdTy5QAQrd5RCJiwS5G+Ch8TfopXAeAfryAW2irkq1dRocCXczqaCGe
IKGo1a+Dlo1JLZR+2qPpl8s4ehJTUFwVdwi24O1xmiP8LfCq5wKQ87PFSG+KMSfw
MlJrtjXhQqHf3JAaSja6sTYIoYzLc7z1PtaQ9nHaIfaxeDiR1dO8KCfqak4cP6g6
YE2ZMJua8Z+1G0PQWaaG+VUwGINCXu5jZNjsmAptyzaoOoj7AAQ9dqn7DNDxTJP+
GH02yx1K4axhcDijZ6fyowgHTjjGfzBBlxD3yh1DL7nqhT37qUrunwpLZlMgalOO
234xvLd9Ml+vN5aMPMU1/3tVKsmYFYipOkl5IvMIv2fY/ypSOiWh8iczJwLwn67n
OO83TeJkqOjnZj05akvzmw2TVKbYD1r3XEvbwhlByWhhofdnjNTduFIy//UWIx8F
StabUSWWLkJkzCjYhA4g+qTnYzHCSbQqdbjlcSXdttQviHcWBUd1iDUNmkJJVOoB
4UMuRLGlSz7hXagSDi/MUHaOfWRfKkQpM4ppvHJhIX2T7DmWC4U8R+Rp4dPUB/DD
zLmsGcOHqnMv5y0MDcNIM8LdyLpw5GORvJIe+yjL4ADWKlkTlZ6xxKvqcOGDK6df
hILSyLCDz1NJWhjEpa1FYWVFy6cnfL3J8yzxOXroMBueT5QSNRimyNGnpO7LOpkA
agN82XBYGExLA9YzV4KhNdeUiihXitAWzW3ljiAVderWXOhFi3VEDYfpz8m2D/nR
AzT5HX2UIN9h575w3axxPSUDbawlsTNrFuRIJn1a5Oo6jdBFLwqzRCZ0B4HJIeDY
3hf9zGLWa3q7ZFsDFI1IYXfpPbfZlLyJWUUW3KNz+f+W1koDzoq0x8cGrow5Do14
NSC3PMCFPRn8UiJwdkyyVT9cxBmeqT22nwzUalNCpRk+zTjsnjujq8BeSy7X9cKO
6e3rD0Is6LmiN/N9qbbmK5y0hKGCRJYfO15LxNelXI1yGP9ZPHJSwrW2Fmp0HzDG
YXx0/N5I3fZx3Z460zCGvZuQrDwpEsWFxUE64eX71dW7NKs+dr4Q2DvVJ8VtoTLH
A3rrkj8rL4CoK3vMk45VOjZlU9brds/2yslAUA0nsWLuCNC1Irnwo3Gxt9Uqp/js
IEG0j69EvTgTX50Ke8qR3KqVWFqRtn11MWjLn812APbtXbCOSHKht9uB++UUDL1v
RnSOmsNWXKmRwiDcOK+WivlMDB01DgFkWkckB4/uZGVk264QRfAfQ6aSTF9HOi7d
u+bCqzRj3PCuNLbh75aB6Pqwwbgqh/+DYKcHTKCtSiwyZIZv5dmdxqZDflRdzcZO
rCM+P97b2D+3PusppL/GHVjUMr23qizW/JWjkfSjgj0RVDxtAEUvEjH1zEjovSmw
aAfNWY+P9YM5/+Vg72AbmyB3HBiZqDxuoQbPcPIkXEalMg0/pL1Ym+noHmvf6NQT
/rRF5BISgaK1F8ApYuw+bMUs0TbruZ40Y5flbm3NWhjsT7rKp2eYlDFaIlhrexnJ
ICYUjH72UFFmbd+D9awocFtw9D80IY1rcoU6fCVMQ6WjuvZR+89LmXDU0Wjsf1tb
9UVICfhm1Vgtoy/2SYGTVx896SDVDYkrIPyi5v0yv6lGi0sefSxuKC9uXdb76mTw
F1ocNUlgLnbBafLOSDv32BDJSnfKhaO0Klm6Cdl5yYwvTs5WW3O0BZnWdUeOYPL7
KMSe2sCintgTi0CnVZ1gox5PBDo3mTCmQNQwj1sUwv6Encc/d6giAQvxRluAm983
52GHrf7Ab3P2g7va1e27Gw409Cfocl9RVhETW6Sqw/locotZ7GQ5KuNE1501hzFx
mdViIqBqKHT/uzIwD+l7SNDui83aB0vsHduJLQIqss1JQeET5kDQbgYgDHL396Q2
WydOcaijaOCT5Fw53tu/nNqy3C3FUoIlFx/zV+nF/d0P0PhRsCK4BVMLcWn+Zp5T
nB7cHwNSMEfqyv3kSMj8QeX2NsmmMTwpca4zbgyRM89IJdaPxjoUVMkkosxnOpVl
2Q82H3CFNhkR3TWeHmKKAtEUWHqO3YFTAZVsDnlPVla+Hdh9u5JsxGi3qQGbpbOC
t+1FRt9ME+Qnky2/MRjv+dEzpniBIu64rv7ZrhfyiK0abzGVgX9fJ64BeQDsgkde
iaVwHAqkgjXDNZ/iQe9EVX4sxga64VDYafzKbw0owPqEkGVZsxeEruzLKcAH80rt
nY+6paWo684v9gCRTT6jVXKqPNuJ6yFbASZ/qQRw38eV5O97DcNhqxk/V6IA/ODF
VXka2o+vor60K17jkL77X15ZKgiPP57AB34y42+tu/boaLbHNdapi27rMiu1hK+M
vcuUuzMh56xiseStlj5Cs5O6rVVGyRqJ1UzRJvjBRhvetuUoM/hsyG11nSWdVAOE
hVdYqyeYWCdk8L+UxUyVp4b4BkN+32tV35bDBBkba5jtILZE1A6yAF3pB+nlBO87
kYZJU270i/sEPVf+QaWI+vC/wmDikmEisV+Yke/lPoxYdM/UMC78Y74pDuCt9u3H
ycHZEe0bOpumfAGiiN6GgvZjA2rk6FJ2t4/dhSSGrOsyVh8MVk5XghR1cjHyLM3x
zMHhDGsKAZ6E1BDWpjG5EDBWFoJOMovKNnYOIgPAyphNCEeelF6+enQmkPZsRyi0
0IAmNgpQWX9KnrY+ccfPy2SZNcKyiMqaOxZPMSBhB4Aen9hlL9a3uuEttteS+v7g
/FsPPcSXXlkQKFJhCyN6jCTGyBfux69Bb+DM+cvHYHlfz2pNPGJgj9pFtmZekYIA
Cq1CfDgP3jZ/Nq/oxu2WjnYthoGFrnqVpZrL9yfCFNf6MXgPa8jc7AzWPBflXblU
TXTyjyatZuAl2/IEgFXRMGr66gwAYt4fDADctxdNwXoiZOfiUzIquw3Sw3raQ/MJ
OZ/qgtEEwaaVjLpVyMyEnL5LyZRekIPKL+DqEyVtqR32avOgvWHT5+bMHpp1o4iX
btnD3tCY9+lrXMglinR+ywn/WYJ5n2G2Wlu/IzItrSlcd/HskacbnREg32w0cpYg
KGMYYVwjYXq4X8if4Ya0ZXoah7djHCB9B1A11j0Mvh9tXBaE2vtFUhnM0KZWehEq
5h+doobAwibJ1sgZMmrPzbMZuzdnZe2yDWoNt62k2SLkpZESpLDCquvRe4Zh1LZi
RUeSWtyOMS9oNFHwtRkZ4MYwpny/tSLhLSsSeIQXR22WZjGsB28YzuUBbbIzTIAq
1UyS9OmSFhu+pWT+7ThGt3NW7+uKll07IQ8peJ5kIW+KkaWeUYA6URyZTg7K2Qf8
SwpcqX5LJOa82Ar5z+I8uN5jJqZdKpL/AazThr3hoOlunftoMkbF7W/sHkFR0UPm
Nz3rKiQdBb2Bt82E5Bujs6BU8rmYl7PNE6e1uV4fhBC6em0moexBbLoR90V3KWKr
3AJ+8WMlQpx2T3MXVAyO3/juoosSbVYuyXZiMqY4GoDUATSpQn4xUZIKODuVaFjK
B6jyXKJbivf0Yt+Nd5EkKUm2UKwGkc1Ga9jm8V8PnO64899Y5NLkD2g1f+jxyVVI
S7CUCLl99NY0FYOpyQWRNHOidUGSGn77pS447KjA6EM7UzFY7cOxELNDEGJo+rHc
zF9+rRia0HHKFp/JVekpLmi7CvO3Ma+pWsWtnQYSG40YW2VSXzDZjDVUwt7IgY/j
5HAYzMB0H9Kc3FS+EEGqWU/Q/8uKx9MZsvLPKQipq1muJDEi2PSluYBNXh8zRJ/s
uGxIj9Wpm11Dp4d8bLOzqZ3C6fbEKIEdV6v8vRUnpPFNZxMLKvMveNJELFR2v2HP
ePtaODvZS3LEiTznyEPtZFIkX/rCZg6u4EP7qmiPkU39jvEHm+zSzy0R6tIXcZ0x
VlpR3gOnRthkjPDlQSI7iGjPZrtEBnmJeT4lHWvkwegYZ9i1NqWOZ+0w7tCMDHBO
u2v622omp4YfvoSDFhG29LeKwRJP+pBih8mgq5rQHDnmi0IoWpZdyNiM+qibQest
r9c1nPkQ2zcNPIk0ldukAZVYNN9N0VOT6WZG+PvvVkBJ1QwSe3EA0rU/ZHDt4CMN
lZPo9/NEijSXa1uHMyez8V6wM6SJACFvfkZSZA4R3/UdquNx8TlSd6gGjgRQvpPn
Vv1gssuzaudhF6Bqqm0Q1m0OxnsPNWGQNfMMnYO3u9Gb8YK7w3HcIO4VheZq0C0F
VIiaziul3fzN0pBVRXbzNQ5jsaNz7Kh61sXQLZyqpI2k27v2NMdiIUTrrzvlTpRj
lLium1XKzATFx/e/ProaC4ybps67AgF0s6uL/9oS5aGUDdqNyIdUepXLcqm2rOdC
AxlRmuNKTxGfgZqlP9T/IcQyW6uk9js4vDKQmr3F3sl8Ld7avrsFb0JqvE5b5h4z
jf10X/7wwdTaSP3lACOgbyp5RRBjB11dtMHHX1Nur+lMZhDnlnHuyuUw1S3xKsCN
Pd3FyRvbQDcI3j8zz2lszAwYZWr7z+MyqD1FHaKAeVDFOurgyOXdcmzDmCZsLnfi
8GHk9G3JODb1TELmIFdsgr6q3axUHePWi/NZDtJS0SieNglkQf2RqwCi2xbPho7g
wKd44aXt1DJ/SN+ogenyrDjXJngCbJTxgAOErklc4y1E3OjjaA3QblcllBLyzVKd
Z0GusfgDELWq2ih3919k/uRFGlPVMFaI1sf/08KxSE+c/VJr/KbNhuF9+0XsviHU
LyOZ0QlETDuiFVcr+0UGayy6mSrUX6D/MWe5b1DTy5NG+TnfXp7hNcVy0gL5YwsK
EA9ti+5bJ6fVuF/5GtC0VgVxvcFvAqmKsqNLCSr+doHjfC29SCB/n3W0Qc3CTJph
rdakbNRZ+nd0F+s7IhGg0qjx+3iLkg9M36zlMxPZIqXavWcfshPPfgNotYg+fha0
iMu6/yYG+Qe2X9BjGlcXcHGzcjgE5dZdLCfhOhPOjzWZDpOy78iovtaPxZUujUgu
aBOBbFnZeKcEedxVBjZrr2WmQFknfVvafW5TRS0WevMUTq3Rh4NuMAqqn5/iO5oi
gFb0X/sYHx19aY0Ry0qG9yo90t91HA/29EEJLIwKuGbFL6/uASJ4QTJHQ1n6GlYt
ijg62StkZ46npK3qJvtKY9yYNiBZf3SIWnI06wDM3hH1zxOlEde6FfhVFBjKMKYU
Gk+G3d4NOslVN6wtaeQNCxHKJwrJz467uMiwHPxeVPIfLVylh8f40mcUNRePSbxn
L/qEAKg9pRORQJ9hXDdvXXuTAiWZYCEgani1FEzZYRP0q5W0IDaytuDDWpZ/jScK
lm4VizjUuCl7MGFXCAP7KxQdZjn+lwSkNOlrcLOLvlGjpLbqR9qnIPkpfwBUKRvv
wBRJcwILpH/Qc30YcfZ5aC7eWOAX4WNnAMSd0TileXVPOpLJoZwUsYrWo9JWA/r1
UZidqaPu4TSsUi8e/Vjsni7PljITSHPW6aqDc8uz1upfb4eCiYefadQdBWcm/1Kr
SkyjaQbgW/OzluaTNGrqRWsBOj4ZzstMwpP38BEQH6H0C/dXU5Y3/RHhJCmRE2Vm
zYG2X+NipSfURDD8bUM3zJJnMWwrBWSKCt4rz5rtzg4gaQo74EqwVZLS2LKRCnCf
F5V15J9ym/ECXU+MtoGShjw/NZnkEgzRzRUlxyP9YnLBnb79sZrSi+870vM4T6Gd
6Yl/Uo5ASpR1Q9kFHib5EbKLkMcbkvgXTAUHP0Siy2GJMmrS4cMwZ8Ygx46+wd6b
MDHZIXbA99pGOxfSs2bXW8pxRlYforxg1Me8jpzVYkD36kXwI/WpWQeJdWC/vtdM
2aLUOkB40wWhXXNmu+HYeIOKgIiOK7V1xMWmItaFO5UPXfqPd98WuVKXvevCD4ly
H73+gMY930V93l3eTH3bDH/uVfIvj68ZgnWFN9ND7APUfgavDIXvY0RoVbBbLI95
UvPLwWtTF1cZvFFGgbWbcFiFISPsNcyhlFcH2TktMMK+5yN+PkCROau0axIm2qat
Y1fmV7gG04fe+T/mJBs+Li4fmKF703Z7NROGm8RS9AyABf3UIyVvVWNuLjmeoZrq
L/ypTpaV1jV3hJreZ91/3GaHbb48cdpuiOloLjmkfL5GSw2FLyuIGRxn/famAmCO
k1DyvbCmZD9+UtIsEbOkx4xMUhPS+Ok3Kj77BNUx69NGOz3VFvhJsS3FmqF0tAEn
fd2i/nllqKEk28BOG03J3M7K7AOAt2igkT+9xnLbWeN6VBvOimgD3CHvyUL8sP2W
L2D2m2MIPPw+7WmRwr5l1Lw8/0BVv60LVUg+K9g9jgGMheNvsqBue4lBPgnvNYqw
Vou691LaBCMzTd03SCuCiOqBJcOduN7UgydcFn3qG5HCVxjQMHWVPLJFldIL/3PQ
UgnxTFq/UzMRhWKTwgkWTGnsc3+JFWPeIrMiDvHbdCW1poBSGxvo1x/revByGs2d
D0f9JT20zkjIjBaUB9tPEzRL1lN4KPMvxooFrl3CIb5BlKpPgSRO+kUqZxZXJ1Tf
hysZ4a72wxqG71eRYAXYIUS7XduSVvgi86oZ/k6ZEHxb7jE5PfhOX9Dw93gXtAK/
8jxkzNHwtBgMZGnGvV236CAY4zU2B49SnCXPTo9Isbvn0YcKwirXSpTk8EHnwSSf
5cwjXgQidmp1haTg6Neus5LOLby1dlo62pohqMMrMSPz7lAl3iPx1bniHkIrvz8D
TSj2zcK4cfIXITVqOb2lGyE60h/yhQcAhpA0QB02nQzF5EnsfQVTfkDCFsjx9UD9
Mq5NZup1eB476uEZDe3Kkcc+5xlhQNCzzONia21v+fSEISyr+SUgzz6PhCT+pwmR
okgDsYNBPGC/CR+lm16jMevbrqxUwgUr3vs1WhH7H2HoNCphWYJPvOUy8H/n9UWC
ifbAC9yTuLSeF70BWYzcxifLyTYZ4s6AnPVwQ6ppx7JjVDUSdGx+MBINNjwjBANg
rwehQPUngRNA1xpnLziBG17MIyZ3JBAHemCOIb5ipiDVsHZCDS/Di4ul/EMqoRhk
BLhNde5PuHET4924kGmS/x+qXYORoG3oX320Gh9JbAO8c/WJ8CA+vjOtlyX5yhR9
clw7ccK1GNqsIgFqnol+8OOBp812MsR6rEbmGVetBfBREnYqqiklU0N3RSJzVKuv
h1qGFpytUyRa71KPWsjrmAnAFoS7XjC/GnabJn+yX/C/JUNEyDE6QG2aLd+xuiEd
HET4NZUdfN5aTI8E736+/l/zMWtTZ5/65FFIRM5vWAUQXEf6IRKVUEn3heHL0QTG
XbXgIERpgZH6UqoBBt4woB26luy6Qi3IwyJ6KV3LPfeOSCwYfwlhQCgX5Ns7I8yN
0VaLwXcGe3cdsyGmYX3v5ABfSYeMSv/1wXm/VvfOjzVl1ZGWML+2Mh+jZi/ND2E+
Qbc8ayOwY5LFdSheyTKGqRbzAJgkCnCEdT3cUj2tpGZtpppWXhN0Pdn3H2IRtywZ
PNyNQTRrMUVlQi8PCeYEayB282G18+o/nmi+ESVxnBmYGVrc/E8MqjH2+AQTO6cm
JY5CfuX9oIUvzyMAkoo7sHpdgGWWDrm6OeEX97FplnZAgDw3QjbB6LdE3Y6jVhEj
4ZESrYKWxGJbnfTQUplirJkh78ztjCFmEBHhnaUziH0dZ13F8Xxy8bha5AYbxvnE
QDBHpv4jn8qJhjm/8o+fKcoTjGhcjzVsM7hac4LXJvEuEh3FLiEntJSam9F//NEm
xGazsfLSUNpM1YuwT2OCPO5OnjfaeaYDiqWZpP/tNEnrLOPGIrLBAacjv6/718Zl
k+rv01hT6jgP2umWvLT2r6W7kabZllm5/o4IkF32t15pdp+gCy5zwr/YJBA1mn5Z
fL3BZp2/hi+Z4O81l2DfZxr12+np9kNA0u0tMwqJyG+Gi0OkR/sahKHxaR52Jv4n
77ktZ20c3CPne3MqyLXJ3EMZ1K64muXA3j2VcVXjnlEObVFkKRRBCbzmphU3PlwE
FhcGxGlqW306elgXfu447q890oSiZG+ICVQ1hRO/XAIxzkc1kwaOXPyEwLpWPDv8
OFuKaSe4YTvBTGFBYFCL05eZ2sp6F+sX3vhk5vM770tyyJ+/Scc71vQN61LYt5S1
hYWZ+s158JJAEe90RpCiN17cxxcs3SxTo0cBXW61rkvttmfW6Ec84cPgZfW/7+iH
5WNMOoS8DGDbYwog9C+OjHOqpJ4BJSqOb6olrGDBOKREhjI6f8TkskRTnnW3puRM
h+EA98EH8BLfwz0DHAciP5FEMrOJKWKYm9bRPYFw/jTAQgVVOIjrqeqLfzEJOOcr
106E1aaI8WXKyl1l7e9lURa/CLembGx+iAI3VIR+c7zYUqjHXIP9QbQ1BWlq4PtG
QTs0ckUMFvNOyngsnLScLODNYdAmndxh37L+ZySWWdGblaBNhgCfFmH7wnY+yFL7
YvmVjmvagI49bQQBEDELgP78JrjVAPj+CnY/xmCaHi53x6vvu+SsRw0eWR1/WWBh
cwj95yS8+6h43kUmNpWmMgraUZomZvefKE5LqVvwDwjJwT2SlRfDub+nLpgmStnS
qorVxmCNHz7eGnJ8QUQ0yoWm0dQoQZXMXR2Fy1I9aXJLJT9ZZ8eL4Wq0pMqPul0X
3totPTz58ay0LynW5QCqe9YGKqTSGr0rUVzo3J6hvnEbpPoTyc6DZ7DMcyUW4F2k
/JMzWCOtHknpgE5OzF8PTRJCA0qcGapPR0Vg4PVRyC1/E1jjrP8IQUMlLxi3C6h8
rGOcigBTgy2fUKLQAsVutnh1PsCu+Sw6x3fu2RG5pEMMDUOmE0R9/CO+1u35177d
3OfJvGp8V38+gUihmqFY8eCyNVZygfuc1/Qvlq9Lh6LTl2F6FCQS+UVrpfXvkaQz
QFKoo1w2bgfFPKyf4NmIpGrs0i5SC3IgWyU0d6yZbbLkz/p2KYb3M1g9AUaiHc6i
HHaQbZtGnD9MuzihcEyTJZbEET0ZdPfhdksqN4atN3wmGsJjL938i+PlvGfNFJTi
WGuKiBLzzaY+DkKUeKiLGhl+lehXDncrtyrp7PWDWjNg3kxyhJsSOxegO+jKt8ty
DNlqZWKziipw0uOzcf25eL03P1R9M0eRs+B74UfwZQc8yXZeRCzYCOnFOiKtHA2m
dhZkI6agxKfUl3l39fROiiT1B9vE2HNBqqa4DVK38R3gDguPVOfzhrXvnEFt+016
86VeewqGCx4o8slfsNf/dYXUtPxLrmfKJdiLulQh2xZnh1KcPKbMeB7eHVSM3WNX
ejC3maZNm9SEUxB21bM0i0ilhhMlH5AyxalXOENQSD/TvdkR5+QNyr38w18qhkhb
zFbR/MZrCKPmMqgMnTMcajARZ3vgrmJBva/TES5Xr+/w5vdl14hVgzrd5JP9S0c8
ECGJGt4nFpupTcaomQ1QB4VzGaJXqrGT2gpVwuKiPO24Li0uP6v4zTNuW6kdnP0H
TCmBpEJyGyLrSHXAf5Rn+nFKtPaK8IuOt7qauwZlNy+TeafoOkc9ZtwvO92Fti9l
wXIusGeQcEXHdZQpX8595BHTdYjx3mQLfKP7wF5P4eyaMbrRNG8FvtMsJ0LN/mEf
dhCKowH2GFZkOYLofy2BkQZlHID76vTiYbNtQMNBLC7hXSm3GZviTnStiPdr3JV5
V4FGfZbqUVvMst6mszDcodoWGvIMuWFXwdc4apSg1ADnkXhjdIs+trhLXK8lps7D
33PZL92TeMYf/bEP2sBHBwa5SwROuZljQMtbXfHwTLKPPCkBc7VvioRnaxC00NRj
zU/K3KDtJsUUUSbVLKw4BVHPgeaJu4Di4zuFtKmUWj9wbkD9CAD7EDFugx+A2kU5
lpgp867J3+uTLZs5OCa4HBIfiP/lkLMvQNTdsDBGl/mU0WgHbU1/3LUbFSLJ0srd
nt9XNCnAC40H/9A+tx5gTbEwQqQje64z3mPjVQbfYp2z+7s5Dhz14k+T81p8OpYF
6IxVA+HFWMCmTmQ2dmqsCuei+Ac1+EXMs9lEXZUuzk23j0iC3A2lWPkgB15jaxJ6
VmQScgn9Vgg4wFBiX2XbmlxjpvlaOxaGGSSLyh4FNEtJWl1Vm0u1WfszvsYFmc22
Hv/Uq315wZPeuxVbZ+PhthrtQvsmKu6tGOEEwrPgWaY/PhiXOaQ6VxggnDfDfQjI
P0HFKA64FC8Rx5/GaxzRQCblMqiEs9IowhYnjcRlfEfsaP4/N7niovGQg5FmomXH
OB6jfCksPmN/hVygTiqxy7GO4yVpYlCYipSV6oijaTjWhnDJkvE01HATxx4XUfCW
cL6vo2Jb53FowuwF+LU9+wAuU8qEGqNFvc6TwgBA6/pxg5AbzZvGQJyOHpxGvEq/
WNXL3QUgDdtgdopBo3XOcHD6UTyFN+BCEo8Vn7cc4uZ7sk6EI5kIb6msk2X3a3s2
AcV1n3lObY1joSKIMMUHdp5RkckOoZaqWRZ0tT50jFA8Rv9rlbt3EQ4Vi8EySV1D
yIOoS6brJoMkpxL3RG01Z6DA2Q2VhBFbaC7buW1f7SdPruqkj5pAQOMj5dz07jos
OpLKco69KioQb2J71Q8D/S7B93BxGBfUisMuuQduBuV5/jpYoQhqSma0pnQY9wyP
h9dNeCDntaMXc4+Be8Iky9ldcTbr+GO0yS3TQ6DwCxjnrNoHU/S8FEfrWuIWK9NV
MDq95wxaV3NhsbQp9Xltz55eCAF/rOkiuKwRFNwfkeEgQUFHPBGndEPER9rW828+
DBxNY64UtKjyQGWr4EuSqeJlUjGlJe2xsMh0W1aq5GfTmd7THpbg3US6GtczBCAx
aKWjdP8X2SYeorTwXK/2RWqy+cWr4uDwEL8jThuT2L/anys/bywfWT9eY8t41bez
12kWxP0MUszqxZp+/daORTviLBNvKZKTd9TSogxtItUHKoPHPCeib09dj9Vcai5u
o1cXFeM4huJt9bmhl1rPOTvoPyLydvHT3I1vCtTNSAP8X542mQAnzJ/dO/pAIoNj
JBKeNTH2LycDeQu4aevocsl9L7hCyZcEm1MuHgV1MSnbaqJN5i6iIAKmE7lqPw6M
QmV1ri0WT/DNgo81g2cWz3MeoFWt7vvsq2ThIELGm68yVst91mT40Ou0dKp5gKre
BIcfDl9WdEkQQF02QyMhLd/eAOMsLStNabzN5fJBXrtM1vji+GZsMCnR84+J3lCZ
o82Vkw/dkZ9cvqjaZu/w2hECkP7gbSq0iwaKCwkLZZK3cbSyx+39RFz+0jBiZtNj
Pk2JITh2ekE0p1ecymx2WmPFwgoYpIYZso82zCH4ZpZ4TlBLxJloTNy1J7dYakQj
XBQg8h+dkcD02gSEaVu7Dx7ueI0uRmBkTeXUnBYbbZlpLafASrd6UdDJukOmRlY0
BgrYO1Q2xbycz0vIUF30svaJf5Glkig5Bq8v8tZBn55oPtcFSlezUPet17E0LBWG
unWD9Ig0LC1Ys7TUzveXLeMMXEud3oVHRZh/ZPTZdJM7DqtDz4araE3ZVbTlR6pI
0oMihrXlRhq9DHvIL4SvQVSjKOK1vLY5pyNuRBYAph5KQTBSsosnuT1cwUEhJziZ
8LbF19urDF65jcvObJjLwlmMXaqQJpKcYgw0/R/l198KNuOnv50aHtAHYHN3plyk
oTw3c7mV3QhGKqyhOM/XjzQVvw+NI0sMVadeWbGwiWZlJgnbsFX1Fu61YMWJLt+M
rmrPAtDDPIfaKaJ8yiUYTpjWDb7XhGaiT6tyByzNQy4sScaN9/u0xEmcYbN52qnT
F8qH8HG60CCONcSTQK/H9WtQ8f1Xf/2Hc4DoMBt1AXnx1EKlY5tvfIgAUjjpIF7k
XR+Bw/xdxApwGof1cjB5jZ3u1HjyzFo1SWOQDbfsy1LjZAmymfxw/S2h+A3vYKQj
S5gGf2yV3ch53AvVxb30fL3xX2kYeomtvQL/nAaATaxAllwyV/0tQ2bja7wfu3rB
efIUYIqamfbTNzluok0PJ3McvbWXZT8qdxOMJjB4fMFYy4RA5dWPQtTdcCmxmVDC
RuSXNonubXeTZQBF7BzEC18BTdtKfpjmx7bV+TpMF429LrS51IdhRZNZWg1sKnDk
JWtvG+A4ZFIkFfrbd6k/Xxtc8wM5zyRbpZXoeRsoPEjSqeH96hNqKP9MqEbhUack
uZWe7SolyU1f1IEoEjukIqeuZIohTE7A7rMhDtNB6JJmZ8tYTZDTA6fh2P6HOmce
oukq0OHSW2G4yZeAq91VaN1NnVacixgGLH3IPYQ0SJoQ1W683V3C7Q6JuNIGSrHq
PxhNG1Rr04HvBIUpvK4P5jP2XOsIzQ/f4TqTVGCISb/aF4OjF0k+7wRnqZxsr8en
tk00KdyyApyG+X7yZ5BEzszRGUo1sVNpMw6gWMRPnjEFDr9/xGLaFleyyis3HpSe
psBP0EYs1p3hIDRs81+4pYgvbehDNs+lRlFLlIYaVqgrP6nS/MVcpy5VYwUZbCN3
7zV22LFMNSaiY5VtTdleg8gF+tWVDie6kbOFSzzimko6OQ62ri0z9PQ9WaOfYaf0
9lNmzK3jzj1KahR1okj5spMwQK+jGl4MLc62bCkz3Do12jD6cu6zYqj1RHqZqL/V
x0Ey1DTADYj98t4LH/o95okUe0ohq8FW+yNWOOrWWzrFfWC2auSMVoc6aulUU8KS
EZsDmNT68b8kbTG4+PNyCy6lcz1OKOJJW4VhETka7U2agDnfORBfuQLOwlpsas1w
9TFYcLJIgjPhcCr4xzqhtq3bgccdbJjcjNE9OXAThCaPcfVr+oNdLtk1Mm29gsli
HcK3m7WgSozgsAxsgoP5X+2YQ8zTDqAk6RAR12DSBEP3lz1ie/1HOSwsYSnU/7YQ
IKeVuAYhyEpAED9axZaeKAcCDapeEZFQkT9ynNeto2vAkrUjc/Cx+FlG3R3SA/aA
44E+AOswJQj/It9+E3e2DV9oZKUP6fEfidLTH4w4YGW0+MQqXH7Q8Mq+4TSzzqnB
3NwvhbYazdNx493fQxcvZbQfLgSvNijR7DNTaWr0a/4ntpi/O7SnJC2pNbA9tdp/
6mv7KC1Sec4hMqxJMVmolhD4PxELQL7cw0I/3D8fRMjrn8W4P8LgxlKFs+qu77gv
svlrg1J3V8dTmQUipRMMVH0Xn17meQ8oFRexVvD0BMTro0dEmrpvaxCZbwH9tBm2
NwzqVFBgQ4FVzCilgZMD1l5URBdDsAdQNOD7HGAhnurpkxISu+q0PExNiU0rAxWz
Zd+3uZHKE+v1UOvtKOWwzpUmSPj/7XoepTD1cPcK1b75R/VywXBac5359UKO0GOv
43CX3s2o8ZAUorOmy/LPIPcNjIuMrO1kA+hGoZMS/o3mC+HDGkfklMyyAnCBvF+Y
7+lakZ+BCbVeDnkUvtuywSMqlQLVK3si0pQ7j58yy1vKkfQ/UuvIdhGXgWO8wtn9
go5AZ5bmyvKkOwMoCvc8CrLRdpz7YGWM0Ry9jSWEbnCealw0GwZWyAlIP3ru18C+
KxfLfMi6zV8pj3f2V4k3HnXnXb3P/go2Bg+cSTYEUYYeLMgTPupZa0q4hf+WvqSB
4wvy10rxQxm29TI9gyKRd34jkb+pAKhBVk2++Ap+O9UvlLBVfwti+8RcKLePX6nP
dRqbK7KyreRsKhGaI0/ecqS4xjh2vJwakNFib3T8MteSe2bAO7FwSACbJUzW1U98
XxHNyB017s5PNIUEep15hQxSD7rlSOw8S5SEhqWwf1DNXQXIYLABqYV2lt6Rbm0f
KXZNW7jFKLZjs3rleN/g+0H+kgSYBON/cj49WI4E9wKvzlB48JnQ7VZtUlPMQnmJ
Uv7svW+dt272GKkG+pSJbJOCf9Rc5EMTefR3m42IDkVv7BkQqugaDmbrJgvMTl56
GtVyKBh0MgxdFCyicMmrgTAB4q+Hr2dQYarVFaJhEPn6y4OyhQdjupFK1yh3A1yZ
MpA8brpkk9lNdxRsMWBPAyLZTvploTeh2BgY100e8F9L2Y8MkfQnsYJrXQ33VRh6
Q/j3l/G9R8NnAaAzA5OWS9EqvOUPxXeZzmyhA9rsTGuGIu49fIFGvujAhI1aLFC3
Nbxak65nTbTbIIRMgrOCM5tBRw5DS998JPHcDilImgcvdoROSYITwHMsisaQVBBN
nUMxTmkT+gbY5vD0qAJP2y1QCeyvIVjSMAoUJYRNZPUiDlA+l7WurMni0PhXNv03
WRXF2Bnp0KaxQ3fKZh5dTJ7oiV/biFIb9HuoCP4n7VsU/U/C/LJFNKizvWupnU5p
0ZVW6t1mYjZJxG/WHjGDSI1j4qZCQI0J/7WK/LkUP9EnBJnDhT77Qh41NsYAPTVj
Sm7U3j9Zg8tZTIQasB7Q6G6YcDyzvdyGAk8I4PSngaNvZgqe9OYyO1V+p+DqxvN+
AylPD4ePnULAXI0EaSEBcGAavrKhLJur/G4JCjzrzuuTO1xHVzRg02fg8z5luEHj
fULBOn4Epn+2/NapREweV2RHBo+Nt0Gx9m6Ptw5bkP3bvbAcaJn0M+xvJcu1exy2
4VCF2S6dpQDGmp9kRumS1QS1m/mwvhk/JY5HqR8mJNYmp22AxftE2HS5DnHJYtaV
G2SRUQnY6okEolJkbGhn3QrhZ5/PdKaT6BF/iLIgAV37HM07hwFkZ54LoRdSdlnZ
oIAdQiCafYH2b7QxrZe/CXzhRlOkN1QrfIP6rbQ2Cn1/2PiwB+UTd3ezj5EnkLe+
LJej0tzXMNwZczkFDbiLQxxdD2trcK0WiJsvGwToimAsNgXBhkfvTZHCa1WaOuUn
Dr6b09W3V18jwOEyqVg9WOgH+s4CO3N0xlsCfUNND0c5pW226Fz0F4Ip5bqKdwzd
oxSwaukAhKGKxnKpBchTwrLJEjtlvlkC/LRtuWcw5yxVwxihuDGiqeT/AWLoQhki
2pGIbbBDqjn+K3tn2avOXH8a3sm/17XT9MRIZ+vgLjX3afyiuCN0m1wQgrFpgXT+
4jUl9G2bYEq8ThIOWcGy5krwxPpCsiQl9XTZoFDv6MybO74LpOe1by+ZRmjPJxqV
N8uTgnIlT2Se1FlWHdrxHNouXOIGJgDGPZ4rzKTejhwnRerqqEjpnAvgxOZTi0X5
nYq7UrOG51Gx0bNI9vYr3wqubxLFe2t2i1YgTx8AhdZmS1kHkImmXnvH962Ca4Va
qO9J/CEEVRnZyqw1bfNSw11upb4CHFyxcc1mK5fSTdwkmLNTa6uAmzXIexac+NAj
jvzcLfsOJ1oLlrn1f6rO0Jm6To4fsVbsw0/S/UPNPa5sokeUlzdd4YlGOuKAY2zw
ttL3976oPKKIlPxUHp/4+ysUzM8I2YM0xMpaL7zbJPQmqHCHbcBIu0xvtO3btBuF
CadyudZ4lbxrr8vxZoDhmle0zd5auoACSiASHsn+KPeLbbcUzSSZ2MMxyhYAhA5H
R2ulMNFfeIZovnfIRRFAEiTV6wcqPVhRiZkBJltGw12hb9+O2FXFkGXxgxHGYNSo
9jKcNqBOK1VyNMrF614YSitxLCniNo2cgxPgIJ44ZH/AydR8lETpVppj6Tnr3J9D
K3ea71rCeNtaNXUgmI/K6FPlA4J/IzR2DV3fnoWhKZDOxEf18PDU1A7+1YuMgCoI
eJRsEKkZOdiRmHjHPkBHMQ7WjEkZ7mEVl7rqzKCTG/3tOMmClYdERfrAOuqxJMqH
Vyb/0An8ttHoJJlVyvUNflv83Izu9Sb2vSU+WZ+pOWstpurIZIXRtTw6bvAE3QQs
k+UqTtLLu/vOFcUzYnGNzbsybsyBn5n3UuDI3q7h11zYNLmYAYdEKi5MaSF8r7N/
I/zBryVehi7e2HETKuNGDg+4+iBLbk98ttd0sVWw4iXMbkH1nAxC8Cv9qVUrBeGO
5PpSCJGqbOTuUmrBpQl7aNd6jc5h6wNZk/ipG9xyCI49dPAHoIqD2jhu9SfjXdZh
DCKBV/bw6hbNtc00ZqDOdMND37nNSIoJzrPqgLc3s9/dukGAVo8WmNg6ncdka05j
EZjkXaJASzIOQwxlc57L5CmwdCvIqcuvOeIUkHmypZ9IlXl0CfvPgil9Ic6fbVYw
cuDDXl9rgt0oleFRmSAAFKdCRnZS815QdoRLBWWapmpBDauXrYPpO3R0HxeQ2kM5
GGevJiCegd5iKdLyQEUOOPerJahL//it6CLhKi8T7wx8OBhLchka9+AePi6PP8Ga
PLYqw8/CLZ2FX9rVlScazx91nUVxnalEJ/xKPlMrAJ/w3HgSnVia7zyNzWflqM6K
hwG+iEpU4sYUwFmrgjLZNSEvMcIF9+RJ8wmJmJj5w9udjy/g+kAO0czkMgMrNJo8
NnN2suzhPpTg9T3QSuXmdcRju8KD6xBUjnOJSeptoBPt8e1TGQhPUQVa5pUXFvwF
DhZyQ25ln+7SYfkWbOwwSda8xWwGAQe7LZ6DK9KeFQMhIH9RjY0J7W2oOFzRt28q
eRdaq2+eZSrlzTsUfrJ5IIJUOnL633XkwzFF0lw22mY0cM/BvWe25dDiU8AXpvDM
VKvsmc4nkvJXDgiErqc4DU9RgM6lExvYvgpkTvG0BJWxsmthn8XqEAXe8GkMgc/t
tIqdJnKmMJxpLF/2MU647dzu8Qfkd8fwDMX8KpcTzxIV8sJ9v2ZblY51UErPD/Ja
OvTXIoMxHPc7jGd9GTQupdHE0B2l2Gqe+MamJA/rhAyvbArlj/PIrvEbHHdJI+EP
0uEC1d0pb7Rt2hwPGrSF3Y9m+mZwtSdg++PvJarpymSeEI195SUbrtU51FilUhiv
+yU21NK8g+/VSorzN2KzLbt5h0irw4C33lBxGw+McW5vLFdx+jzkhI1gPjO0kilT
IT3ml4WCR9qDxYBQkD9juBrFhnarATJf1LJxEofViZtRW5dHYFgyCFzSjF7L7lxg
/EJ1xPldIilEmv3NRwGP1Hc9DWvDnlIiwbZN/tvi55Vuxtozov+WDL0At2vaW+qG
T6iImYaHLWGpWzslCG53a6vv5ZZFUpBQ6nfqRcAHAhGPKh86LgHo3P7Lc0WMAhxi
0FhDvRpy1XzSdcZv4UHSmMBFByOMOnMUv6KpYyk5HVo7yWsuJvh+t3OG/IRfKLSL
C+3GGBYTPW5MS8L7wJYmCgdLK4IWtLArWiMb3q9peyibTciN1RkfCEADqSlAi4lX
DZIc5KfgCzRKZuEjQiJpaEpsbz9yJMOGGN9/4SHrxUpZNMvetOf2tHB7HrfBJ6hI
xSr9OsZ1q87VTEmMC1X43ujSZOBW4S3SIzb7zdXxg8Ui3dqpNe6OqHkIv77/cENd
NOGErZh3fIKphJAt1wMmjVmXG5PK03T9HgfGyxWi0qgPPZQ2esN81ldu0aFl//MD
3lTTu+PBNZxsnp4eOT4+z7tqz+SH8udMBFGQb0SAuxFkp3/TTGD1bonmPuD65SUg
DrCXPgVLicFSmDmgyTQ6zV5WL69dst5DyOlAhqRgWqblI8r20/IJf9y0J3p146WR
9VrFEe06AdKI37tdZ6p0Gk7BDrVXAxNP/Er92jMu7XKACLccilJyc/swEzhVQ29Z
tUaqCGea1RtlXV2n1D/0V/86+YFk1eTK1yska8k18cGyb+lSQunFAql1RN0ApwPU
Ywel34E59+C0gKHdfU52ICfmaAF6fFHiu1miMXch4oQBuUuHEMkGBDeCrCAamhLI
M7WWn07tsfoUUJLXdM2kiKaFDH1hqNhjFsCDRBRDm8dXdsOshXR4an7SgfYvN97I
XQfZDXpvfZpeKbPETXuLCSlGiCSX0ITxJIgP3GSWKNn6yG2u4pxlzjCHUQLUy1TA
jb73suu8+U33CW36izYwAqVccG56iTByzTdZIRw4YN4LIGP5VsUrL9yMgWK6maTC
sCgRGXitW7Rp6R9LvSq0w26frHhuwi90XwOFN0sWdVmuSrqANR8zCK1ziGig4beH
cZbDkd0V8SThZP1rjZyb9zYZhJQ3MwGULsUGXS4/leEf56e5rHUmaTs6Oxq+27qy
3UfcPDhonUnhVY7CQ5AR9HyQyFePBuJNxC9uZhykHSPGAJRXeYwVgpBE0bwVDdGV
xAuC42MOGnTr0q0NVu6pBawnh+YZRhfKH29Qh1j613JrU+WuPRBrCNPdr8PfPGkt
dv8b9I47kxCs/VbbpQUA+X7laNDL9ixvjWTlaj08yteeR9ze1bVFTxLc/y60nMO8
NPSSn1q6bih9KrcjQKr+kFIvrE+P5xkrjAHBMtjFP1inIqKcc9uB99b197Bqy/hz
wG2srH80ku5SZOgTYBnqAaMyTBLY4cwYxPEet3Z+ZFfqUDGgzox0WmS7YRLT3y8u
KNsnCz4gGKZqjHn4beIrIDS8WijCCuyuAyetYGzGQlWP5Dv2C0/46O0FqfZqrc0l
DDNVJRWuF9ipSEqMLQRxtCYu0tCFa1QUPklL5+6G3WYBaTtWIzsuRoVBxC+1v2ex
+wGMzUjuB218Rg0cSZLa+HCKSJDelW7ZGeLOHZCU90ZzlniaFEPBRgl0KbmIeHeb
QPGgHKyI051Db00LbdF4Bceb3NUR9kCSF0iqzYmoOhXfCKSVJLPOjJgMFNw6qfFU
CXduqODL8XgfjIyRf2RtiTh1ZcVX60lwqktx1qYx76c72i0PFG5OlqaJdJuS2NI3
yKimsHRRYdsr9xVbQCj0y8W7QdCurPp3ZR/SiGpl+8diVfsVaJYAFtM9EdYGbe+j
Ao6G+B84MQrAox5mvaPddVYAEzlrLKbFEkgPkKVtIC7ubDkbxGQbbz6UQEWlKHye
CuxRPxzPAamy6dW15WYwh5pWrLmjMU3h4pztp8pmKAq+rJEdk1F2maLcwRcip/hI
S2Etwc18Tbsaosnb6gneRQlRlS+mEqGWVSAtrGNymAesb8DaWR//DqnqVmzYZq8o
AL3eG3VWq6/0YC5l30r/FKbboav21yt3DsyfyKFnalT3dn29jlBYC84tUT3qLJN9
0M/jOOkLPWDSbM8RLCQ9IOaCA/MkL7XCd8KETnp80qGRWVGmuPufo2dLLQmeJpRH
Nh6epw96+XwUUNxjnSZuGFgJrcLJjOBDfOKD5MNUOpSNZjcxW+VM85z7FJ48qe3z
kK3cbR1iVeoXZf3lYIJwYDl5PpS6RkxQkxiPJZQ/v615VRqmjB5mGdlpIXee/T1Z
UdJmzg5umomEYSk9hX/0YQFgQFl5EM7RtCT6ThbwohmQ/PddAiMxxOa+puYDAO2i
yL2OT8bOFzmKvBtWG3RShRajez3SVqlBuSA+/agBVgp3UpS6WcFATFuQ117czAyn
+m3XtKcgI8wOgzeWQfN9t+l7DOayw/MapG91+yBT9f7CbCWr7mudMhma7cka7LQa
lkwRBRILyXoeMwJktAOdnQk7msQC+X5E9ZK4cLX9ZT6tqt/yESyUnyfgPGBHiGkJ
TjU4pWgIgOm0gNPDfYLXHVZ9DDB2NPh/MPpUKhoxtnfqyQLdz0PNu10PrXlgr6+e
SbGlmnyUjx/SML90jjDJGEt9+f5TjCsbFt7NuEkiGtzyiikdjx9cLYZfllzdczd+
9M38AHvvrxEAKEqjVXPPmH1/K/BGmOApZ5vb8Y9En3ix47e0d+cnkBckgjpxgN5Z
SGCYX9OBOjI6rNkVsd70rEKGgxA5Vpy4LmHQcFQkMyDYf2B43ZIqT8yrqSgF/HGt
4YmMLjGkbBuLdRImMuHIFrwNFU0eOiDuG4e1yeCDVil4l9PmpsVNCH9FE3TJqQSh
f+cml0xFHGIIKEUAgwleP9LJO3t6x8ESIrAPb6YeBc0HK/ioz846filJkKcN8zBd
wLdi3B11n2hrJUR0AS/f7HQaAFGgoHITPzRiLqPsbBp24hCeomVLErEx1kYADD1X
Ij9HrRFHmX1XExU6NV8Xw/epY9NE5aqd0TJ3XK+1yaYG5Gm7nu2vvHkh+QUZGdqt
wkQNuOuxQ0qPsWOkOuejoLL8FDGsDwvwCkEymXdVk1dG8L/lifQmGbbD7pMbbe8o
88LCPxutAZ/yeW7Kk4Vv++Jr9EaR/M5uaEKQvEPbrhM2yJlfsKVpi3RyCNdw9rKY
G7c9bZ/aMqWPlDYJUHg3YW5N6F5YMXW5N84O95yyFPiqGXWMaFokN9ESVsO9TSHP
zDdXjWHhfflUijaTOskFd7Hr9Txsli3nUUf1TPYPAsmiOCCOGuw9N9WAaFsdLYQh
iJxXZej5YkWc9TSRK2qMPmg4ZO8xnbrapbezSiSNF/EANZrScuhv43MOkympVOZ9
iDMjk47tmOOglNy46mJbGy7qw8hdfw2mfTxHZzxwAbrhq0tVz9J0/ZImzo3xVfGH
xNQvOAcBU/WooeVkEFzzBJu43MmUwYPFpKeRLmuizos7HMguPo1H4NFKWIOaGsve
oOB5AvfVqeO13d9qS2+5acPKnTnA9VZbPPMfWOPtxe/Pps6r2K6w99uopG2gxH5m
MQH1HDWMKhfQfoHI5U7OhXwB5rH13cBd5CUD0fH06a0kH43GvkAS73XifTfPFqxS
1pJPGLkiLzKJ5lPMUjAnYs0UQLD5KFnIquDURFemzADI5qTRO2QeWFNfSvX3b99g
2FyzgjkfjWSbpwoa3DLvJeoKEa8MaPFaBbxAuxwPF9pdAHElcMW0FmbUzBoS7p6O
Kkw5aX2+x1Kl3KxVMLaEKTvML0lyxS+AkmW18EAQkB8+uwnS9taokMs8Uw4wwA3h
HHSuYs7e82C8AamjJSMB3TaTi198GbyNGaY7/IJrgJ+v1LL+moeiawxWkl2zCUf9
9IzBYEJP94DAlKfMw9lZzLlTIxlo6TrbKrUhWmy4H656h/SYJ7Cd4RjzGP6fe4sJ
OI79EE0OmrmfU33zN8oqK9igZEdPd8KVzIIzMgQlh15g6qksIyXMcCs5WtW1sDqI
sTnrUzqKpikQ15/Erz9/6ggAL+SV5eX5sCVAmB9MuDSWSSc0ny0VlMOIQhrnIJSu
bH9lWlqKzqH86eqHmE18RnqjeUmhpKcfL86Xpx0iY/DPA8uDjEzvv0/csXm4sHx4
TVL5edteX26x43OZmUvhgAO6FmDOqNh8DGNww/O4GOPNlrzL4kRdOqxssTSemE0U
tj7zOIsf6n6IS4wL9i+qrBgZDANgCaYnbbnEpx1Na9UP54iXxWTsbotM5p4mtfy0
eyJqB0TK15+NTkhzKVL4eYlEPWz1x0g71TQZM9eYMnYKoB/iWqumH+OkRNNEDxIO
rxj29/1A6CfeX7+olMiR8/yQcDHF/CC8hVU8K9rO2zZw50cNm5oHzORxx/Te0eZM
VL/MhZOXH5rifuXTZjEXjFJQBuBt+VDUV7q+0my7+yjfA/OAPmFcLefgkQMkZ+ta
rpPlhPwKIyj6Qu86fQg8NuTGoSAd/DcZItdM4uxZazAPvdVMJOB2SEzXunApSpw4
Rnp83IT0woNmPdSAoYo+Urr6T5K3R+6VYgMdGHx19nwxWcwE+lV+Be9wCjMN+nIP
PSyKeK4PHrGx0F7kTM2QnICWKphO0MXERCROhZZ7CGxpL7zOf1Yag5vOpDMY7Zbd
bJCzE4L4ulnkv1sYnvY9rtLn0ev+o8/HYOv8VxRNptMtgJZYv23R51uW8/+DLo9W
ySRdY75OOflafaDBe0Laj0Rz0OyliuLEMOejyL2AgrM/O+nwpiwkiOy14R75A31q
TfgX5Y+bIMVjFJza1nU9laUOh3d73sd07icEv2cOAz4s+wWBx8ELez2y5YV++Dxa
lU0RXIX/Wm9mAZTCR8+0+dMzDJbm/lp+LWmaOns6ruP3M8S2aelNqphgaOQCPw3I
grnI9IGNcL40hRaQb4xSoSsrJ7TOkF8xHpo5mNCFZ7pt9BeK8NCiASsO7UPhZ2H3
/kMor1OhmscaYpgMBdim9o8tTzMGKC24BS0byAKzHQsY5dj0A8pdWA8b9FdsTkPK
YzFc/971DGzwr0ZTw+ffEW/Cyiybo/Gnbjs+xILeoLP6feXjdZ803WdmHe7r7JGv
pyq64/KPZWIBAUPJuz10U6Y7/AyO/uSdc8Ix7Kdp9jisvpoFQ4L1dl3nBL4FrSCJ
HVCI2kdpixGQcMkJh7OX2wpzWI4Z04zSlnkecLCq5m1QAlNc+Aptsztt3fGXZukl
qwLP/dxAhtkFR04FLsjNLM+FsQz8Nr+g+BMY0tILA0ZkpUVWMatKng5DQO/13jM2
3af+EvCdtxOFGZ2sQyaM2X1j7mGlhEughf0hALavQ7RB/8SwtR2+FwRRzU5J/Pos
or3xeVcbqCMN8K9COfOU7m/QEYtNYEWbU8bPkgdp9spMrk2YsyyqGf4FR0Vjjebh
VsqxTtFR7ZxteFAOIXnjZnI++7ZUlAGQmyoNrXqWiJVsvbjle/kHtKJUAKuzySiL
s05BCP5wCvxm0zmx265IchcRnobFaJpnmBPtJPkOtGVDjYnjd9UX5Y6sfq76dh/4
WH9jHoxLJnsM5VB7ST5fPNOflsgN/gGDdyx6XEZEqgrCP91ucz2i49euyJYPd8td
VXAfRw0E4wcDC7ycAXg6fxO76ZqVEC2aFJDF9KoPs8+sWlZL5AawiHZm5cMvrx2/
nbVml3H1keTfUibNZEeyklJByDer8ZO/9D4HUziBiJI90qmqmAGo6OHz0si/dI1R
kLjSEVHUjeBWZb5Vq/up2QVR+GEMM+Y9IY7yJqSDBqC9NTwhvgZpj/YoLuekXbYQ
M/S6JpzDYOIyy2qKO0f5FhhIlSlJE25IZqm1z1T564C3ViheSxzHVZXfeF8IuHDv
6dESiV693YTQ1cb/oQKn4kFystBeL8oG1KhKhcB0VwDww+6rP9IdAolzp6lotQXm
Gu7w8i4HYsj5RBqEzAj9KjtskTseribHj7aAchlhbcDFLDQCjINTznGuqPtw436z
pQ1VA0o4yZ2s7DOLl/Hvfrafio8AkpDs8LWQR2/uk1GpLF2HtQglfuyoZolW9qlc
zL5Xug0KmaF4QiDdOJAAdn64WtZlW6KTKJqY0doaw6ZxGybSW4MyxVIlPSrFXkDu
kgXAQ+pem7qpLCHwW/zR7yNPSsKEEhR8Svv+uflY+1CLw8ynAeAnqgwYs03zuZPM
jQ4fk3cscmkvs5y5VeYBssdpXKgP8UrN99fNFzRsYH5jji4psFn5SaV79PQqiWEW
CdY0eviHDmsRa//Z5uzyGuL/aoROGb8xQybI4CyfwT+zXmyXlY0yWAJ5GWH9dZMu
K7XVkvt49wQD7Va67AhMRxbYRO6LUzSXspYnAmACoxE2S4z5LBMmVeB3+TuCkKjo
AxkiS1zu6n/zqEm4eQSD48yhoA8hkiEIAgBj8gn6tu94gVdYMmZxbgAjapCbfJOf
Rje5LzGutpn4fK2RrL6igTRg9+j9YR+m36yKG4W9tmEWdZjy3dDFU6Odn/6Kt78M
gqb2z2faNX4dBGumtZArCikkgtHZdcGneqxZTKwwmnTkGHPsxZeIArixl4mPFswi
/HzS3NuZa+VwnulN6I4TGXDr/8/v42MPWmM7zuyep5ltfhKp382iOayp9ZOxRKGv
Mt+vcJnwPQGXHv9SxiQGVzB9/hhj5qvizBaSfgsWyclqfbkZ1K6kljqMPlZxEdD7
jJ3szBHCkEhO7VRgnBKvLM3bGsptdQEUMlAVYylefUSWK2hbWSPHtMKn8ORbTPpQ
nGWEnijp6a+1UqHGcY8PMA8xLK4O8aZyC7UJc7yI6x8cDXwROBq9bWZFHTVA6LxI
RUXvndjfT9bKsSg5X1jOZ0wONVzNTsstiUh7MDRGXSfH0/zMh1tuhJpnN2Wrxabb
lC4QRpoTYcU/NyJWrHoPh93qCT5eHFAsGO/1nvLlZO7DdoPP15aC4L5sizlWkaKD
mCtkdK0dcRRE5SlXXux3yuJocoVgmuIrHN/L0Fn2rv8MBMHhQyVjVIiRgR8DNci8
STdPMtiP7H6smrzz0VSf5z413mIg04Cx4D4ekMcCN01Dw/4XS9euxmoPDbNgR8A+
+I04l84qzZQ98aYASahYOk8a7v9ysZgtYMqDm2JT+WUNJMB2tm54KKven2iZKd3w
w7aFEEhDVJrhpjFoRpXBGmhqnTCWltdahcks0EcDTDyWRCNWVB2PBi627w3EJLgr
/WIZp0duWumhwo/zSlWkFRzaWG1MLJiAUjl/pd1pJPVP4kASMblcxWkCiOI4n+2o
V1E2hw9+8zC/J7U1vb9xjQRESjgovnTNU1FYtIA1gLc+n89hgJm1aWsCAEwPqhQh
AqEjEzp/HQFalK/YCI4fZYhBQYeS/8cMxFE6tBpMg6IhT0ZWcc+ei+g/bNpdJwq8
C/2Lvj7dma6bP0MO2PSlVL/218khHc2OEjmkZsRC432sOTQgXv0qNQuoZOrXA5S3
dLOXi+6HqcdsqwXt4r+NoLBzno6T7YJymA/ttISDxlJTXSm7Y36JyOr1P2G1nNt/
Zxv2iE6dLPhJyftdmd/bVZD/TCkn5uPWVecr2xmbE7IJOfW76b32O6s3EITE1Yk8
PeBQvPV0qgVjPARFw4QvaVxJ2lh5q/TapvEu4+RIU0V5NjQ9sdD1S60x+x1ejrEF
LgNc5oYLyCVKvUONh0IITLwsHnU4Lrah2itgOti0TSF9C8QzglhoL5BiNwDSIHDM
9506cGASkCc92NbuDxTWYR7qjwZKpEZ4BeKHDGtRbgAie/J4LwNIn6lrD29gmMW/
hrO5rPUK4wjH3hkfJjRufcJ9Afp/+AevcBYVpF3+q9ItVxZcRj6O2btOJXgUYpWn
vZlNb/kzC9edJ9IoSdWUXf5xWkpukzXp4LIGb1fVAhJy8LgcZLXLhafoU9qq7Q/S
gHaVHdH7RuRL2JZlCFcuNKUOGkTdSrmKmHthT41qP/+A8X04U2RFh2nn/VzhqrBJ
NXcAbN97T6DeQDzpFw3+Bg8AZoBE088zeO3AnvgaC8qjfq/Pp7LyT0yWQ+hMdrzE
3ddGv9A6ZmFD7pGt0BFH6Jfd0hGUY9I+wmctZ9CcRSmpJjONExzzhtTuzqov21Tk
7L5c/Tx/X1LecPgDfzV6+S3JqNj0GGrBITPUo8E2a3QhYV3pInM+xxuWOt9S2nSb
2pinLa0/ebrhl1MMOxR/MTfAf2ICUnuJHccbQXdux9xQJIplKy6sy5zS/LWdRubp
DPvcpMIHDJp/66kTDQeAY/GqMM5U5+Fn24q+86DWJPXn2GoMHso39tCdhGzYCZvw
MXdcWcoM6Tb4Z1Mmp3KexkM5sNawzPzDIPzykKTc5kfgoX4LBaRiX7jrNwtvDQo3
zooXg3jGttQPQcynl1LwJ5XA1Fm8sONlejx0YgL8qOHQEF0x64WWBKrSELHLA/GO
sZx9RCNA+eieJHCnTvXiBHfOfWzMHRbZfxslbTrfRBKs6l3OdoUkOeuSI22ccpHG
bRS/ebytEr+1ZwAGTewX5B60nhpYmLwG5XT0Y3FwbxFZcIez4y+oD1VXPvAE4tKs
y+5yQQyraLq5+5q3dg35l2koENL1BrzLxG/MGKjIfsgsye4i/SZ3UNPrrgP6oZQq
z4Reo3/WJLNlYhwICsmQ2qaGBhf37jG0Qb3IBcFkaHukZO0UABxI2vjs7+xdPDzQ
/3MunNpGS+crrKgKglJ9i+aqlNELp6LFowWOfDhk/YgSuQAkV/dHFc64LZwSJ9zH
tgOAJufoy0tddzQTSCb6Bd5Ps4D3JjS7zBElKD3Safi1yzLO9oRjPsm5YT0NissO
6Hcj0NpWWmXKJdrKHGRlfP73/c/mc7DtC0F7tVE5Fv7RDXZyP79WW3E/FXZFrqnD
9FlV4kNA7U9olJgdm1lpifxLb/jqR3W5BnD/U74hbC5ssjVaXDevISjAk66BxLWj
OL9wXtf8ItxRT/LdPRDh9RGJwnv9GaaRNioDboSj1ZK4lkmpNEUyxEnv4OeMlFY5
gGSRsF17xGo47UenDcSjwmVJ4ishmivgdYo7gLyw3tMo3d2pzlpLscrSRcWpevjs
0ui07aLGIL6r0ia83W1wLoomXk8UhOz+dS+n+oxV3vXPEVofsIGfbwcvk/nSJBOk
H9yEaQexqK+ZAllkFbo0MB/CKiNtt1S/vuGjoVI050nPo/uALTw7fGPq5mn3kXkl
Othw099ba9ySnhGzq1hPDppDPXAw0MQhlvenvxLsnFTIgKBvHPwO5DvSiS6BoS8H
IRh0hJjO83CsHc6SDGHtexalsalBSlu0CAL2qsbw/8g69E4VUoah4I4psOLfpLVC
BQWxaQc5ujfcJPFHCjgdw4tb5fOFPgepgX/jQcYZDaRtrn90xXsFR81+bErpeXUA
haBIWnrwzdfjNujVaLiOAgC0nQHhvf9eMX5touzf83Z1j1uNEHSJ9Ik2SPRcouy+
9Co/vfVnV+o1O9w4Nhajt7jaz4XdijoqvDZwsixk9wkbB6VNQLNLXp6zbMCzdzDe
q7Gb3eQHvbs11rOsAaiRNAEDp6ubbkcBQSTuzoDHa/506b3VFahd/nOlZQr2CC84
9I1w18/niMafB7ikVtkhazdSQCLC3VSzmBI/4uL/dkSrPEXLg0H6Hm7z0mQ05aU/
rpjKNgrYYTtR7z3mTBL23WLX0xwhIYkorQcHUqP7SJfmnHh++lgbuiULx+1ZRS2H
DtNSpbgDnpBrpZg/+mMdeAF7tV9xbynlfiEfoys7E8yn6v0eU7SwWhXRoAylbUfA
manmxEopl1nSLXHzFs1GTBjkvs1xttBv/K/BEqoziMMEVhpWjBqf8vgCQ/cLxxZW
0UjEamAiBgUxVgg4xqtfuESVIiPzvj5ndj+vc6LQgPJtndrtwbUViYUao7HSx/d6
aUut4whqw/ikzjVk6ToVyoWavKOS3IpKVpFR7oirUZE5b+d++Bc+gEo+3qQ+AGfH
K3zMvRO0Rvl5JFw+zjxWRRgEjN+ayuDeBAc9ac2pIlDkFLWWmZoUMJOCOoZczIJk
bOQHrbe5oyaML5mwhz8Y3+6mM2ITtViUsF7GKJJj0EoKDXigSVUH6kj6lVLjsXU2
baniczDT9bZzITNoq2RmyrWWASzQVmZAHQ4xDMhdAPUe6ke4SY+yUWuAyb0AhIF6
Lc05Wj1qzGcLenBiHWYRMy/aiSM75tebPAfKakBsrGAFPC4kb5RUD201WlUlWmaH
A0maqmV9rR0HELCdgDbFS7xb/FWZXoPhtDxyY1EfEbvvsDB9LA4Sin3e7EdFqfm2
4gtdc4BspP1DFTouLdGBBrTp8Odj9W2l7E7FbG8tKChK4elaMrz7HiUI0Y1w5EoN
RMx0nOiRey3o9otahCv2M/5V44tvft8aSqq6noKHh2ECMYP/kYDVvNbqRQsgbO/9
YIDFadfaZpIwxcgB61oabNh+D9lyG6P27ZMm0rHDmwW7Ln+ZrSF+38mPtifITAA7
LaziFqsqPLESZ5K219XBgEaskQvxXf0LMEn5Ob5JAOyayk0G/5IxWwIUfqhn8ZrZ
4PT9MdDnRo73OPPA/L1R+2oW/iRkcUn+SJa82hn/5llEWgpYow9QQZx3AML1ZM7b
LR5z27JQWvWqT1YD4/4H4SzFU3XnEp9rRPvnouiek4mw4yKeck11TVMOl27JcgK9
YMEBSwyMma6dkAxZB6PmGCzzwc5SY8D5fJRlk9y1RiYTl5jMKGyLbWU75G6nPlU1
FtstpUsAADlQCRoyc9VQ0t9kviKtsedWl8LSEfxhFwkbP4JTtZjhf40tqifgnnPK
VQOJG5fGyd4bMIPq54IHJQubzNn2RZpvs5yIITyjatlyfl4so2a/pmeOX2siRzqz
ar0jzF0MRvViy2lFiH/REKCYAa7I0uyz/pICTtfPvWt2t1kIgKBBRhc7YzKfEcDZ
TgD4xQT/cF2l1usU1+D/1wd9SViY1ml6XesY7m1x5EfhQmGPoO5IJXfN4zs8okHd
QkruVSIbvEkhUwcSfg0yYjXgCi+Oc6R8nJt0pvQnDDlnZkwTs01+gyaH3hLwDj14
zEHP+cTRuwDoI0ZKHMjggPkiamLcoN/g3kjhdMa1Vn68XnbnG40YN1Y6FGmTjGmk
/t1Hu4rg7WwQDPEBAO07A8kpQVNB0ni9+WFmKQf3eOhjLrqAvUAogfm45kHv16qH
oj/zE6A5KFerNNW4CEEXtfB6CwxNyvVloJl5jiNyXwUHCa7eAH44dwYDdOhMsd69
1ExtMAjA9OTLpeSXRutFSOOXQ4sX9isXb14QmhmZSJ7bDVkb1RLhX659iTmXiMHZ
38b3y7DHAPqsDX49I+oqLJ0fwtDGwtBkpdaCMGMuaIflnTUYrxRCFh3gsx1bsmv0
3GSq/rzGe4x0F51BhuO67beGX4SYavUZv69wYBB6vyJdvdRjuzFlYuZ1Lex/hSKW
/rvVhJSECHLJEcvb/yTUy7LLVDJ8q5MubA2cdTgFowYCr/fjtBxxXO8eh4xC8+It
VhaHTv8IQrPo6hrt1ribfOc60El3X8/ETb8Bd9qTGmV1bKAVUveo2cJnAXIStMGs
omxXrrzcgHYCRJQlckHuMMWWIkmO4shtRIhbKjn5YffkCylDtbNj6b0vxzPliUxk
obdbwmCv2S2IWVlwpOEJKYprngGSgdFq7r2bY90xIcGZPGeqq8nT31nEbqMm6UMl
Dib+niZc440CBDyENHVfZuQG9MRx5Na4mmZuYsEwiAV0D6obC74U1YoO6Yt4CyNb
vP8+CcR0VOW5uYeCNbDX9XKTNQqcrJIcYrYCNhFazAcigvd1F3k92wvs2UQTJMhD
WLlRTn+wv6XuImUnafQb1xQ9CFCWnratDEJhpDkLbUpSEC90VoqfHGxB4/nwIlii
C7LR5J/Lq+ThjERSwzeZ3XKLLPKzQ133j2Rb/8tve1SsnOPHU2KqM5qhnB2u9xEC
8AqfnGARH/7hAE9tZmT2KPBgjgHAlAnf7cWM/a0VI9cdJJrNKobzLAYFJe2Mgije
Ll2Hjx/No1dYKU+IFowIPZXzsRiyzWgYxnMIRt1iC7Sm+P/weHMWSCIn6S7KGy52
CE6eyrI9OgM3yYabm9YZLZH8ykNgZBoVXeGsvx5BDa+g2F2QQ3LfpDjDvbMGmqbG
fRYrmkRGF5ixMQCwTuu3fzj1ExstDHjdUCyfknNqHgxmB5Dcy9819E4q/U7PiWVA
A4A308s6O52KCKnSc+0qKu5BsPZ6njY2uKh/zdveBvYgioF4GEWEbNrhyfte1Xdy
ns3+KqSLGSHJln+hebfhW1nRTPbmjEh3OGAYHs68lYepa0zhUxYzu2D+PTuUfeV2
uMZzKIHib+oQom+VuNX1JF5aSm86TZfjofN1iydbQR/VD/KoCbmaRxT5ZHApa5d9
mopXetXs4ocNXmq9469sCJhYSnC7LPNvgqKXNlLd+zr8rNWyWZc/Y5zBNRD/rwFQ
0Vmf15KfBloVfDgwG8GjRCFJMneL/Em0X0JsUXhvaLFtj6wTu1ZodkLCNEHRCXky
HucEoh/057vyflV8X8J0kxVqx1JPi3hZGohtcnEzlMuFf4mD3I1RGkW4PVrvRnht
u3F88ZUbm1kQMxTSyU769S25yGQBtXnZr6b/rFgWgDIs11ETH8qYzGeWeTc8jFyd
SjzIDHMTyy1e/NgTDYOZA+wwowz8a5Q63H2LK5ojUH9kn9c9tbbYy7tENVpaXj/4
gPwHwpwfTdG8PzCqKJbmoeLtMUIk2/uTq5gI5Fa7yc9CYEtf+0cNZFHisfs+Gyhx
m86bXRhUX20vgGBvoFE3ojPDEdGoaJTdiUyTadePQZBSHeijuiX/2C9X46CY1pPz
ugdkFVXwMpJyglNg6dickp5f0XC80KvtehcuD/wF8HkjkrKvJbRIqk0+mBBm04Wa
EQ2rxZQWCJ8mcQLE7lMqbC27UzUPgLNuc9RSw7xiPfXrpY5Zp1iBnye2www6PDNe
pjj5X+Uycgdf/BCVxDzZZRiqWefEqODEhBmSxcx1c7nyGTlKNHk4VZox7qAaSjh1
mkO6r37Zb9xl1FTH0ilCA86vDOvhtxaZKx+8xswKGybaMLSCoALxVenDAZoeD3pj
fywmUF+RI8mOfIqzZC0dD599O0pJI6DeqI/CMin4sR8cM2A8H7BpimXAdR8hG61m
ikr72YOCvwZyxgk6gXU8NzLSebm08e6wFxCt5Eu68wscf/TNcgvQ8cYxn2CuQOjP
wuLQUW4rJMH5JstpJtnljRwOFYB6J715P7OqWre8U3kvBeHdnD2EEZntlMDbPDJW
rXBpUliDdxf0fuIoE4pDjI0X3uiRcVjHfwA+lBkV2/H0EZmVByJN3YDknhxdfuf4
snD7A0MRhHi8GK38e6ur42mz0AAbXHFPwgQbHLld7xQcfZdITRFjQkfw8r81tF6g
ZqF9E/YkZqyqpDdHDi6V6GHa36ssVPddWvaMcqKQn8i6jTcjDITJsvC9ieGiBMCj
5rEcoM23byLXALOt8QuGPxhvnyBBfw0ig6OQR4xsK00r3qDxd7mZT+l8/DRkuBsU
Xc8YwZ+qwS1BTaPDvAetrwNpHLNfT5o59/EzqAOtn7ci4xg/zNnS7/D75hfhsNvv
WdgMI7ucRG4miFJ1hLFPOLqjDh6BlBCljcS3liN7zWil6G1isbGgUqPyQ6Nc5aYE
K8/DFRGyFbJmAdKZeB1T+EnAsr7zfxgus2GjYLVoS8bw8NEWa/T0WD9ZYs7FscV+
Gkn0OULsr4+1YlP/zP/U9cFzC3WSOfqZ3IDJz2G6lLuaLSCVQfqkzyyJAd0XV6U2
efzEtPDJRUI1uo9C6hCOAts5/ym8iXU02YGhkyp3m5N49NvnC5o9SARJj252hloN
C0y6T9J5tRfoEgSGxFNauV5s7jTrk3mmkn+Lxrn1eBQaL6K/NXDvKvjhklB1wn6f
cxucTICNSLzPedAWGHJR5SaZEo21BoRuq9iOAyo1I+9e0c5e6blsXiGuvSYsjPmc
0jK+EAbprZbe6ow4sWo+YUtdRU6zWQfQ2YFfvSoAm6VnnYmuObmDjNwjo9ABPwRV
//cXdMq/d3KEPEBgRWWtqxmWVPvOLANB87K9pzBeh2HUdk/MAPXkTqCIYjjcP1VX
JsAOZHCw6OO7gKgeAZAX6pjnYny53PN1jNc+iiNjOyBrfk/xluTOv808VZ6ym/Fc
XJog1XbpoKbqoIL8Hiya6ijDFeLf0MX0taaJvR0ODE+B2K1OAd9M4DGnvUTMXMHW
rlhq8IhoyRX2O7F0DLpsqm2SitH2yKrNQ6srn5PmL8zaitIJi4W2fRB4PSK+6E7w
cu3nHAC2anjD2LuY1mOXBncEJhccE5DBe3LC69N3KqnwOonvLG5+moenbOXhU6n9
YKCdlQBahJNir4ed9ybuKQkWXHNORLWIsrijY96fP6oYrFgvubhhQyZvBilBHqK+
SmYE2hHdpkO4k5XCP0egrni9W2lexyQNUtLvGXZ7e+ZYocgAGogxxEVP80CJURCq
mwxT6UOh/xNGkSHQxu3wUCXWglT5yJUMTX3r+e5IHZbZENCnhFZCvM016nuqCkph
sL5V22HeZ29dHBnvbNGjFTJcE1l+EnOXMCMUZCRfqf7w4YwGwKhhBXB8hA6G9eiN
v7Tkol4qFGKR1amJogERiHEtI5feZ5+CFaJAMJ/W/d2upbASp0nbzL0MpFikSK3L
h4P+mUUzpM/y674/g7icYIx+znqtL1zG6CpkaoFH9TjLV0JZSjyy3YSzZYXk+yMY
f4oPNDvbB6lYN6MPnknV8lmYRaJxbkpPlRKK8KXS5+9o/u3KJ35lidAw6BYb8zAh
SKEcyLzDbyD3eKUzovgF0hpffBzTKEQQVL15ToSTo+r7MBK35ONUuz9kEgeqFU8C
DWsn4hTW1rjufFHiKq1Bo0a/f2Sv09OyH4CnsKxF/iCv0t2+XoJOPniL+ipHANIO
ETM9NTi5k92A66PpuiyumhzBxuTx3HfvIitiz8x+MbQv95MYXQtpQMp2knXQ4mbN
XZjkEpdCQQMxmRrfe0Mo2RPHQzC5wphhpYAaT080GKt1Of7kHXkMRu6C75WlbDX1
7UkYs4jd3WeEcOSyCwKMJx1G5ajviiLc81Mt0/YEGaCRbUO1f9sHnx8Z1prsg1Jg
e4D3IIhrIKMVys21Y0v+VTNYFcUSHd9WcZ1YP+pRqJg4uWX0/kGhVm/x30wFzg8f
/8Hl/VVuil5l9yWRFHkme6ZC1SSphqx0mM/PPcPDccItpmCdKqrs3rKWA6Iunh17
fF4pmoDYDVjT6H/f4anShddJpVnZmIxkbjstcX1bqrxVNRr3TAiJT+UH/IDSEgTh
urSq9MrIFefh9jv9RFla6+VH+85XIcZg7PrPpDztnrsFlREpBJEj2NjpUgm73B2T
p8yWCQ/YmTMBLq73Zki9bCYzYSu9Ga0RS1F+++id8ngnaFYN6jv3KyKV1evbjYwz
iikqWtbEem8hLrb8rdJOZCABzo+XXRLQ9amlAv1TG1DFrGU8vlLciZF4duu04PUS
HZIw6Xw9Kg+V2AtWetZQ4p/FkW/TWoj3s3MA8PlUYgXjkAcTQvLtqLNCHVr5VZNh
70AQmtY0ua95UKXbiPRzBR76k10SXaNP2VQymjCGi+PQOyp9WUQZPh9RaZF8Adu9
ezaSlqKbDiA0BJQ9u8XV1xugNbfNtGSw+eQxA+qHAt/qeb+4qv/hH4rlzmsvSxVi
KEAGoYYxgayyh0LtitkE7Q5sevp22d5deNfsKJADIdjCUmwJy1OKOdU6FlWO7wVP
adnxr/fSuS7gw70BjUacVIFxNVnSW5FT1iP/iTJGTcNh4fFXLfhbQGuXM3A2pPwl
Dk2d4L6jeTgk9+AON339zVnMYy3MFN2ZjaN7JH7YIWPEB4TGLdRZX5eNZKT8XW/e
zBGpJEmkQ/0yRdqDgcxtoirq2fXjegIcoLVMRZhgUgq4X6tR7yTTKVbtV7PSvPql
JYaUi1wrp9hJimFXkXbCWG9a7j5aj6wSyiP/RT5aXX2eutPngxA+02yivVfG2uwO
FiADKkKmydD0HtlHqiD9KgcLhxFq1uB6lVGm7gqzMkw04LeQ9zC46B3qbfYTxhRN
2/OzUzJ6Ns9i9GrTwZGk62/RnqZ+deB3KuUcCNdSbl0qZ2nRRozx4MPer7GqUhuH
PE6FQs/KSBqJX22HLIdjxl7Su8c1Hs00/kR5wOGah8U372JjEZ97zh9nCQkrjwI+
HsaWTuw3nIvj+dNQKUZ9Uw+irfxUl0nWuRDGjnl8bgZQNM/9HgI3V9s2gnqb4ft7
7ooewNpqt2Cbudm/FM8UrVTxVKOKD0BaKniwrmEGPnbg+7oBAPrwfBcB3hx773/t
UFNCVOzICNTxeYNCn4Sgd7XEh5ileBg1bIswfZR5KrNsFwnV6iG/KJvw2V8c3NqR
wXrFEpm5fbhQDUzaqFHEfEaFJfZ+uu0jLfAwRU/PsMU2fYS1Qv7tYvAtQ6g2VFsN
Mq0FLHwtSJewr4JQayUatSwf9ubnXKBjdirvveptT8+y5N+vicoEjLNy/ta8NKbJ
1DAsf2cuunA7B7LS8Mn4MnBynscqfHGSk12LftCu7b6D52RZN0qTkTnW6y2WJMa+
RnImw9KUnYzXQaYT7x2sBt/YZjeUbj84Djr46b1S9WuSx37s7i0OiAghpupFksch
FM5IeEohbFB091TVneQ7yRGriPY5F5jslNHuxx4NOAy6jSs/Pxe8WU/f7L6XyBt0
Gv9kHCx1/eKrLjYTEly90ksvGxbmwyGMzZksos4AK84hMCHiXlnzFo0gRpe3Q1yt
+nVtJGz4oH9dYx7WVuci76ZvBHfqBr01H21R/jSBJHiYJ/Ay9xfR13fy+Boj02BV
ZZ781ixCbTgY0t7VXtrSygp7Nb2BuHzqvvSmczcs26EVRsFXtBQiFwu76Njzsa4m
gLRvozm9lg0kvpdOea6hdkPcWMZXAbtyPxlg38sCu30Dl4wxv/eIodD7CUbzkO5U
Gzohz1uHmRIByYp3sazq9FSH6qh9bBzuWqbgilzx1eLS+euuaP1pGnWrpxY15wCW
3bRq601Q7HYhBY7poHm46xl7qbuFFBPigwv0JTPvyEsdSBJNwYUWTOYTemGUZCaR
mWm+byBvNgSfSm9xVvYHmDwzvP6YEQQFYv9SmysPTxJMf36PCNEzBrG0PYcK9swy
9o9yROXUjyDqxquDtsC14jIUuGy8/SmAQtRdJ6UQ9aE0GcCt/rncgfXT5IisYcEO
nCgfZ5RSRveL1lOXewXyKO/eLrcT9nE0Cm/3fK4Jwek5bN71huos9IPDDPNca9Tm
cQSldlb+f69r0O0Pt2gDflcPVDJHcddk5/e2SJzNTTyGqYkkRSZXZ9vbRcJuYXMw
tepPdVl+BrWW8+5WQG/57NIsBu2PlxQ1u0bnHqODqc7hHBnWWLcdxN2uIzNIA1hm
r62FUHAeblK2+u2RynnOe7s4o9Ow+LNUiRqQ72+Rq/GME4poMAJnqEFygOpWfGeC
BGUxxgzueSMpINujx1mDagkTKXDFuxEZ1xFAyDh5yBSsdp8UsNf2XveAqqUzo+du
usQtBgckB/XYe0Cwx4D6F5Hdo+erMsSkjT815X3k6MnQHOy4sU7mPqIM66rX5Pe6
DHoVRb3s4QNRQOLGGj6yb8j1FgnYzYT9ESaT6fOJjQaCnDP/kY0cexUiZe9qyzFT
ekQVLOHoKw97KzJW3RG4uS+h6tg3jcSqaQA62GpRvhuAh8KNEiSn4GL+SMrw8Vy9
oIPmoJWXmnv2vHtigpWAG9faLSTP3dTGzMWBE73ly/EfxevIB99g6EjIiC0ncK5g
2KYBWUM0ecVBRiMWpWo7nyeLMBy21NWJJYGlogXqAh2qTzGe8smr7tYO96ZTsDVO
py1yRDa9FfJTb9TvrfcoI3x8agVKDg4FxvcKm67kFXupLG4roG13QplfZIPPmWD8
CjMOACItX6fgU5abIhqCsqZvZnAo6Zf6PdoZSPfmz47HNpeIMeVfLTKEU+BLxWd/
Wvti34PPAdJ/6hxfZ2Kjf/oOaxGWa8lloxb2NWmVqyzcr/6qAH2vHE8SB6L4C4iP
4ik+3JVLHQG+9Xi8RMfls68ZNrbTvxCiUSNFdGGs8AJNnupBq8DLwexb7uZ3i+wh
nQOv0Q699QtTMXE6uHqtW5rvG9ygUFrHIQKI5+SV4T0AFLKgkqJFth0WeiNpjAO8
JnL1Q32xQ3Tifk8wtgcwUCR48vNfX/8SYSzjZTxiAkKk/VZjVjwzbfV5bWxrAODX
kUOgnVzp7JHUVQiQe68Oq7BKdsTa3ly9z1nPliC1jFrEfxjtJbYA4lBLbMeS4Dv1
rOJQMPVeFWzawIJYiI8wrbUcUeMt9tt0PXXBrzsjqSYNJsCsfNB5Vc+Nek8plnLu
HNlRUpI7f1DZ7t3LxHPk/Okp0PTCW4q6k6z1vcDEt6FRp5VDHH4I0WOL7M4+vh+k
LVwin8RBHR9IlVbIDOJhh/Dbd9qvWik0TdOI6MT1yj8qNmWfvGaxKvVnz0rgL2iJ
XxsfFWwqooxKcCQbmakDIbOqGYnJyndJlUl95vZva/BZPqfjG/q9efQeYzvdeYSY
ZfrwlaSUvaGJdQkSmT75xUQ1mB0veb3+I+0S8Q1qejhk69fA5ng7whw/zlN5hRnG
hXTqr5A7CLbWUXaDMbEU5LyaJhJMxGZgF+UPE6DvXi9g9EGLw77VLsSEMAhuSp1a
W0sStbbN51VxcEO8dN3FxsQXPmEdk1OXzGeqarSi9NBSFbSzFJ1GYrHHmPfM1ztD
TRSS13fLka7joYuWkdCuC72z4tzu22XJ4XjO0ZtuQVCqvv7ltwdUzWEubKQz2zUW
A03NuElyvw0wdhHujgLFDHnt2x3arcoXHvhLbkATLJPtK0PunFmp+UPScTDL/rVa
Tx0JTMP0bq5/lis/EDIvGhJ2SBx6OYHUwwOHQnTZsYES0NeJQEVwNU2ANOYqgU8B
Mm19jKjVZ6VuIGeT9vVjRkNhDlhN8ziqVgZIzGSNdoxSljXsvibhKIra36jneevt
uLLaxfv1drQG+cvJSQbpNEjDEr+88k+7M5VNl8BVl43Ga1ApqMzHJoaIm7tVHEmM
KvOEE4QOt+4UNMkWINOUEZT0eiYoYU4wyZ7BMj0S/0XPImskpLRPaMKE+BIeAKwH
2y/RvF/ddfI0mttNtW8aVsgifw8pUk0BPwJgOfPUI1bhydN++R8gYtqTJavG1IAO
oTjvGGQK75rimBxzNhA3RXaAW+P1eLEupSWt/RCqR5/P1hMVWIeX5ktbfn0PW8VH
Dms8bgOe+/CtMD3tmrk+hOzhQwCdK53HBtR3zMQ3em1gCss8xv5jARdNPpM1GOnn
uq2vITeklYjhDpq7YT0bu9RnYrcE3NAVuhG9ftpu6xYx7tQlvNfEFLH/cXZ1mmmE
OjHXTjkYAqf56QzBzymGgr0DAZH03aL//rA4QOMmkK1ylISpysA4hZBw6t3cVw5j
a4TyANjKkh+Vg7TLn4YsZxTUY154oVdxPqXJptf57JJiPtD/HxLa7LGWgHoZr779
rygsIvy8IzXxtcb+zCgg6jBgziUQfogjFiIFX7sbzdn8Ox6vPN7GYkYbuEy1S+cl
5dw0nXCvdAamGeDfmR39qdrG0bJV/tb6TPcpwugJ+3Av9jdMj6jIaf/EpOrAQRDP
xDpi7CenAdWhvmb0MeFY3M2psF58H3/CL07xjLv77u5HQxgaHDSHc3+CN/1hFIgy
j90Xa6chZwlyhNsz9JW/nkpxkCmBQednASFg6pBZEp3+wp4p6ShUDocAw1wKtwSS
c/5TfDcNQNhbgAg9btfzhgEK3cnpwDXcGSOqV4ufXuT6ydevJXjqZWo5aP1IrMlD
MwOIeZzzaxCktXKp0M26T3XS+WqZ3eUWlwM/wFzxtBF0hDRw7Y19kgb5oIoEygbd
tvUjQdWAiRcOnNYk2FBSB744wFNSzH4E7tXHuZpOaLSUZrGrOUCrG67i5hXozT93
ny7mJVwrV3vIXZbAXQKJzN78ZrKIta6FfOwcUO53kTj+fy1FRURw3gSOSLKoIByS
b3yZLBzBSC0tTIk8W5La4pkGrPc5a5SSlW0xDrayTbaf+piSaRKcgiRdS5fiAUDV
Pf76uqxx3AnytRkMFI7NhaDKGiWh7qsXnCnfb7AAgaLDTFE+GVVO2o1SuyG2sbSg
Scr4Uer6FPgXCAS1sRzk01ICcy/nccn9qAgNWjdQzC1H64RMYC1VNv0RhmXxu3FG
WQMdgb2v3lY8Gk9D+mdgRSZjaaY1d+Fxz2CJInqoEdHwKTLNkQ6f0hWoBsXxoc1b
3HeZxoYC8/cKUus3w83lDCOOFexrDL7bUsAb6uFxmH/BZIZjrkE3Q4PLGxDAv5oC
iFJCOnqj4oxSoMh78uet1w8AJasDMp78uFKgYme5XaxgLmdO7dX/9Ti1DC4rsD2A
qaftBRxk7EGumBbicAmDzZoWw6sYLz1tLRvSPhZsbZ9DKG1U4njm2i6whi/7i+12
6WNW/GJ0KkpW2QNJj8Az025Hk1+APb1WujUc7IOXJo+E6hws2KIX46N69fzZ3tcr
7nGSm46+9f9bgfUgkZ2Hl3v5sKaJLuh9+qGSCdV0sgC8sQe4BaiQXgvaz0cx3okw
Z1DHzPWm/tKffFwlGYvC22q5iTUjJUlvLRQmh5DgNRWRSyDcsIafG/ngqwRCS8b/
9Jeh79z1dNj+dl4ZWIR4rsoDt7WuPbptfAAU+6FKdairSrf1vdiPKf/heow6GWI0
M9dgBPld1jIHGoceWZ8qO9whQj+5LDMZ/VkHIbtTazn7GZTFJ3ce8EL1gtJePoyE
kqATAUDkJL+5pSO3FiplwYUEhzt819y7J27Hy3tHo0X7L6Y4qEHmFJadihSDSE1I
njwBpyA3dsR2sUyGYJU2ZcC12mvGe+LQKIgj1rTAx1wkzK3LzdAV89PbLgk9Giyr
uP6piPtbv/kqa4Thy5aqDcYdvQq44p7Zbyf4uH5lKG3+cLYIVFFYrmDfsQw4VAZv
OPkETZSg4Cew8nLZpKcl4+XThbspmKLXx+dWhjExQx0rm/OOkZmp1S7wITD9d9pV
IvRSnJM6WjqpGeSGGE7OCJHjmYmOZ09EejZKKXrMBPuewGPr8puZK1O94grKpVT1
1Dgp4TDgupP376utYK1Yn/FfoJ8m2b0l+pnHcuw4aaPePjmhi42vaL3DHbvQjyBg
FEc51xvwlGZKrzVTv0jUeXduzs144stRoAAdSXKTOwet0x6Lx6bySkI1Ljf5AXra
VH2VnU1E1wNGxg0GGfsQV32jTBtWKn+LFpmVuAyKPUuZnJrtptH/XmWp9m8La9h2
i0MNYHaiRgvCjF+GdQqJ7/ctl8DBWX4odkR938yqD6vEbVKDJJDMSxRifAWNE42o
MyaJLjQvMNGnujOfYOrBAcsh1Yh7YNqq9+Fr7l+cxU5AycCrFST7NDUapBp7NJp5
x+gbdoyJgwYsQQOxudNLBBp+vDAjlrbzUdUWPZKEJ+5HgbPB+4l0FpAePXbQd79w
IC7Q58Cp9cowlgGO29DnJ4FZIMhEXgGpXh35ZwxvRaoyQ1UrokzPboj9OHYgOCEm
B0rLOG+cvvpdXcOZAERFIRvrVaebQuNQt+d7hoRWYbo2jCmg4nGGvWEEbYpwtPVJ
MtkCyWIZHd2LQYooY/zfAGR3e2Q4sWe7YLq2OKxVb8DAoLQNjiVN39p7bqauKjZ6
b6eBaQGIKdlXqgLQuWNLBOLSlqCX+4Nl2r++Wb5K9I17Il7oASJvS4jbbXURs8+Z
wdGjx30QhNVoVcP1b+ljY9fMRt4hn5AdbGQl/dJ9zVZ4+BB4q6HX/y89KappB6CH
k/u52kbqCTTfrg3tmXVtRbtAWl16ipUkUu6TgIQJfaRTwEw6H3ykq2FhB8FrzG3J
Nr6/g2WBwLIQ8XEpfql+hpoXj6CEMtbMeO7HMzm8ioBdKAWsauPIqj8gJHAMufAw
mFiSG93JtYLAGJ5XNG1RmNP3M5mTzgU6pxsJelRG+0zfRU8pg7VTakRrcA9Ly+5K
f+4kiika9vv97/krZj0Kn7lKknyjRf+kWHENfTXcyS6q4gtUqBFl6S67q1TqQ/xD
vF0J5DYOjvTVqjPEdnqmfaYBnO/bM5oxo41sC22Aki/PyxAkmNAMzDIkOtl0JTni
Ny/gxDCgBEKMC0noFn1aQ5fUbkOao5SpRhMXgrqOEa3XvAoJazxwKJzgyLMrD0Ty
+0FfCJ6Ry2cec8BkfqdmRfeFy6hv0yZd66Acfcl+FD+HdfjzsY4CXM0SXv3qDGM7
6nRKUVyZM5JdFQ4V4/iODt6PZqP22tRV4KMzHISdQ3BIOFFuh2pk1NxnWi6JkY9y
XEtFvHxllJF0KcJCpg/8R5nQFHhXbC/98i2GX/PooQrhxW1LevhSTeJUVA43N4My
p0JbuozYoXx+F1215sjtZmxQV/Z5X/nVFagmB6xBykR9wVR/51eR/UeLRFu/rNi+
kjGxLzam93Kw5Q5OJwCkHf763xsUuXrEpLY9duGm+i8TsIUAHt2TebGEHTTHytDe
vK9QHiz3xhx+YdC+/W3yfRL3awrU/4vWzRNbx0jTsgmvJH9jWtr9XsynIbo5Yb2N
at3yWdmgpvdLZxFUhvJPlYgU6dSnDpCWxNvMEDQifcHWtoxxHNm9RIKgK5AeFrbp
kdjKn25h5uf4Upxpkn8wLJUGVxu98e+9VFEcE8rYGTJtlS7sgFcJq+xNO+LZ1z0A
SrYdUm67GU/q3lJQwVfkPhbgVdkvTcjxnZ+64GcoLkYJOW8MC9oy6AnphLxAP9UA
jMs6CvgTeoRCCHRPZx2aTE434pf/GeJ3UHfZXjog6wmm7ZHopomwKvwREfwB9qym
xSr8v8eSdrHs9R4104scxcMVaBJc1n8NcUB2FYCEXSqiY0Jx5dZ3EI2M+NPGsJrR
FkFP2PHtGFTH3IeaHdxUOI5XmV3QJpI+JSRw9zQwVAVOmN3WlXyOuxOQsoTNuJx8
DBGxYAUrwynBBtFMa38iEkRURp0x3Bjb0DLAKmayw+iA77kKHU2RCeeN7bv2iH21
0UqXzgn/uN3ouYRZGOkBKcZDT9OQBXt53pKvMm+twWkuJ26mVnnSyHYxgthIHHR9
50WxxBChoprgeGLkvd7mfJiDpHUwvYoxMzfd6bHFJm3AKFGgKNRPtRmbiKh7u5wQ
JkZ4Pf5KPR1vImqTrQHCCyeYqdOmPizBBfdJj9rEFudKWNQ5szTqFiA4dX+a9+kM
fqykKLG3HA2XVbeUDRHYHFZysAwvUjISdTKQFjFYgE3MXaz1MNFWEaVIr9SLssTj
XZ/rmOjixwj5/W+ZE8Z56aLQkaGAIUE3mGFoR9A5NBa5xlH2QDcDU5zeoenQSN2C
799m2Be/1WpMEYPOzBTq0J2KvhHQ57aBDYaJfhpekE/eTw093lc0GGQZN5UvGG1I
XDQm/slfMPtTUoFI0lu2EsR9OGTgpCyhACHeNFz5efNkmZ+cEKf5Ih9oEkSLqAU6
3Dzd6/7f3EgkFqpoufA4mipGXXpaZRIqcIW/Z+iZtgnpXeQUnmZ54GdlEssmN3oh
nF5vTnVlhpF4PZTw/pPicIply39zEB/Jras2Gvumj8PbbxuShNYvi7pxVeHhrtm3
R+ThcVDx4Ey1qRpkXvNlh51Q9mOUEIX+7CKV0yGE9Nen7nTiUoquu/+1FrUtiCfo
5vGW33sf7gy01VYTbShugVo+5+Z+o/HVTTW5hnAJ29ZNMMXcvLXLZqW8G+p4Zyi/
oq0/Ycf/C/DSiVEYvLX0FdhWCwjgU9YXlhUTtesfB2LWNPNlL4/ZupLWlYYCYhVJ
MrmEMy4AzKQEFIpZa4xd1CRF40+xbVTqbezJvkdCQNP0/cPvKdg7XSIVVc6sMnXY
zjVsD4quW57vXYf4U+Iw2bHP2RWLvhNL/UazzDGiJV8bNBx1yDMYB3M0PTD/Z8Tg
aKzi2zyfXU2jI22rFLvmQpgYby9+yo6Wqo64Ww69AZ2zuPgbJ9aDb8+XcVwV/Vap
oWEGxsu7ZIeZjtac0c7CFyJOA54BY7YXdw8eHWqmk/zM/B5I90eu/wSWY7sdYutS
yGAXiKdoAmIdYR8CLFascQYTdXhtzQZUqO70dDvjWDllYnq9bhKOAV+M7FIjWsCx
TkFHbxn7+wOfMYBDdWgDeUHm/xzy+0Zwwx9bbJRq479zUpvayydk0IlPh3oLVSC2
F9yCwJaQexZRvwYuZxz/c0narltMleYksraoW7MXQkIVFgYbhD4c1Gq/9PBjGJJm
bm5efeWbb008eigrL3uCPv5V74/vweSbzxIhxzJaQQKmExyQEi6lfCPfgbR/fLGt
lc717YbydKTfOzE9+63fKj0j0iiCQCyeXPTY2ZX3NAW4uRgO66GjmT5Uuq4W+RXi
l1l5LbGLsRqpXdEgycA5sQp+06lUfp0oRHTgq7glHFrTgsAIJhK0T/5tjBqLXCCQ
6PwYXB++71EdUdmDcEW3pdB5n7Joxo7BEy5ZDgU9KKf/kvC3yppO0dWRSwSUsGIG
cnZ0CaS6qErhskl4Xp6Mc1GMczVnD+B0Qg/w0m1Pym/hIQApbCoHKOJCl+Ac5hHM
/zzR0VPyAPLxMU5NX1y6o9PSueeyuBlJKuZCy7V5LnF4arbTRHgZltk9w0nocoTN
Jj1FwM14XlbvZPTPNjbuUsmixcO3hc9DRwFovBmLRgESpm9eauDFkz21rDxCBty6
zF5zBA32W4geYHFnMQ/vHrYbO9Ly4GiFRYss8mZppskdinv+y8H0CmFuagkavqmv
O+ZRRe3iyaaA9Zw+9vmYKq8YF11636zk5Sbn3AXGGoiJyd1pEn5lEYVLYZkRqIRA
eWUBdC//E5ZepPD4iXh7TN77D0DRUnr702Bo5QGl7kQDnb4YVALEBqeqReqRnoKc
T+/AjjssH0RffzK6vdtjrDwM2xOajv5+095Y0HjrZleniQM4TWcSVZWuSJuKOepw
NY6MtMLaiErPnz3zhGC7hGxO3gwES3s+Tmks9KFuNAd7GfqyXP8B8miph2g7nYVv
qAd6nm4vfqoyDJBJ5UYcYKZu+HxaMVejfv8L/SxhIe6uh5fMMtTOiNrFMSzFwHnI
XIcsPTHOQBMpIUPV74Qug4r4JKdxUeCGl0+NzterkkDXAgeP0EVzpj9G5dG76snI
lFTdXLCNUhcuxUaxIMGSsu7nPmN1dqP3td8JFnHaIHJCJe2lCVkL2v2L5J7xWxYB
gbruar58EyYyiYtS8ji9BzhEk7ci6QClwvEN50SWTDF143mrBbEp0jgh1QPd8ag0
yE8i63pE0d1b40Dt/jrDoOnY8uvV7AxKlE0ozJ4RAEto1nnO/KOnWrfoaCPsiwHu
IZTUxz0flRyZOs1c+vsMYyXVamZn7V6XUVqzTLFLTat+xO7t2zkuS7xqmIilTB3L
6MW8iYNa+arFkwzCEfnNw7VOOAhEDNsC0iWPUiejaVXDa7bbjJs3SWGTXVdgKAhD
k0IEmX9EoDtnLGLqgTGtG4EUv8vohaDjlV7DRRn67OxCk64EFgOPOEl2Qu7u0U1w
BjJK0bFWPULDGRA4AhYlM7+mNow6Tx08Sma8O9wN8QwHpNba1/TbYSoDelnLdMeo
R7UoluKMWC1mHkWEEfQToLzRO1rfvO6GzpszgCIJD9G3lBUvAQz+lSNulE75Kms9
kZmy4kdLYnI6A4rU7YlcrKcNJNvBoEWg6QTFqp4ZyB5ZSaNwbA7HDlqORc3XMw7c
95BdaMru1ffax/PJ+7cDFQhULsren7HnBQ5LD+LR2L7V1y2PiPpLoainRjCiFrEN
ztSp9k9YQcKNXJmjgwvZT3ooMh8CcX/G71YP8JkJkTyOqRGG//1fH0uCuA5/UWnT
PDHF+Cod0655vZnFa7mGQ2jSSAMRFQpyaBYvZEKBvXrSrdxGXwzgmo5+ROXhIrEy
HeBTngSgvHyyFcuPl/Uuq9gxuaIwRbPZV594tutRm7mAJbQSX1LbZIptLAEXu8eJ
gwljsQsctgnHEsaRFRVWl3UaCdppsJ5cPAbZFh96FmCfpu2KmRfJQdiwfvX8ZQst
0k8uARf8e/1tpqCV7itH9jLqCC7mEi2qRf6xc7hRUteuLNHjx8Zoco72xampdmBv
MVfX7drqZ0tdIrFmRYGKVDJuVkoPUtQfqNuku7Yk7OQhGoS16etVfSV2XHPoDsXH
xmYHsUsL/3sGzVAy/NW2YcHceBnExF6Ijti8X4t/U8eKabVUM5Y1T6zSbyIiIvV7
9b+18lDTAcJK9nqRgCADjT2q+gmdravY1n5hL/yVd42UELSRygNLWWP/5+lMIsQV
eCV/f1DFzkODXfSJCrl/kn3JYXWW5oWB0RCZ/fTHQgZwvU/Gy/5jd7r67Tf2tTAt
mtTRgcKMu0UjV7dAKVrbnj5eRFvlNA7VDIpsUso1PAAPw2zDa4zFSsWanoGkC4sM
qmQla+4RdBZyhLXxLOlJjz9FaHVgCcuqwYJ1zpbKdJiF8Cqek3fmK1u3XNtP40q6
jneSGFBxF+fU1gL4hdxmAmC7oLuC112acp7N0RhnZ/sXsaQG5RKFVr8+liYZA5VD
x+EkBtSbUZtdfIz/JFz7SgO34dG67S74FRmuiWtOdcuAQixa9q+vxNYNs1Zz9fdG
mBzuz1JnpTADvWnt97pRMb8bE59+fapq+9JYeNVQJXMUnubhWsyXfowEWsab4UH2
HyiiyIA3wt5ZW2eCPewqGNViTm5SFMXlI7qccfjoPJPP3Nfvpdiy6JXJVKtavkLQ
/M+VJwCUb/UPjLnzKJsYhQ7637eWQ4qEEZgTleiAN/ARoF7MmJlin7uEi02qxnf/
rK8RyuAkWxaWsIqzFrNJfzvS4D8EyG6sYs9OgmRfXqVP1kQyWTct0tbpYgJ16qBP
qQx/ULzwbfXhEpDaLnHbw3/XsdHizCT9cQixFkcYIED5cvbGvwzNEcN+O6wLj9UK
w7oX5ClnIpV374+nkx3B+IGppkMLWqt5uNZol83mb7EjdOPExXsRMFTTX+ETDmmh
U5cEfk65pmpTcPQbgH/EBUtnK+Okgm7UbvnTAsb4xvNFTIrp9q3fI5EWlsfi4k/b
Y1/EGOVTuofqB4s/hXYn2fkBijPE8D4W3amhguwW0rXv2MojXsgSNk0AEfm3KEBy
KjqogXusaSmc/ca53XHylNWOeSji09krFp3HMUJqnaX5EY6mXXvWtzfNTzqihnCa
M7WtolbIIquxLHJn6BfIcAifmsKBjgPb9Ra8Kd2fgVkUDnBdwkKXPKfZ099j9jYi
3qz7kfV3a+Ew4QJY0yVjR8kasOL+GfiLaUNWcLjz7l21axY/yqcUgOQNqwISIAYg
GPGTmAZv05W74a/ROl72cbTVpIqOTb97ac97evPFcXc5Snb76UJIt4/OPu0t7/V2
lnOIfEobnxo718qe7JTvom20d6Ztgi9396V81ilWFqrRoM/Pf3w7M0/zoNlVquhi
xlSthgwS/gIh9pVLx0X3nOn7pMnP3EcgJJA40zQd8x99zmUm90n4kNA+tZXR56Pc
VbIGmSsYRmosXSgQd5zLyyKW5Uo4k44TzEimYNkLVjO36t08M4gAfenuKIS/ISx1
dcNBH5MNl6B3ugzCMKug3MoopIv+t/DAA9aw4lT5RErz9SQe1cCNcLSj7547s3f0
dpgY3MLbamlNK/5sOnJ8VZuq9zS1SwKvcLWnVV35WgslxF8ecWD82crFx1xOD8Sn
4cZ8PUFmDG78S+Zw3DpRU82eKEDhREn9Fg0HS/MyDtXtlr1w3+bzUaRNgjD9XRx4
DlYkYvGsBPkkO+4k0PIz9iZsSxUUOEEw0f/BmMcadWrM5vgVBfhY4py/vTsF2HGp
WgnaomOfd8+Q85WPbhQVM8bp2Doecg8TS+cMbz+tkuR84TCbzCiqb6Axx0NNcE95
dfOZYqn05xCmVJW+g9R3j7X6Ak8+ag8NKLB+JWRMbTrO4PWrYYX/3bBAR4pieluB
afR4AXfdcmsdqVkVYp5Byk2+AXiP25UBhp+6XBdBkE6eSgKR8s7q7CSdDVYcFJ3l
oqRkYtQIFIZkmxtmUg7XkJDf8ezKBZTZnPmaa2hGGn2SMYmQKUIYU0k73z92k3LX
JkSTZRN+WTqb0jYDi1meIuZnOK6t9WfFnn0QMV20mVvoT2rwCQU361UfF5VhYVmz
cjZEreJHHcyujVBY23bDe3CzCNboc6X3i2TbymJh4OpodjGrdVaQdyl8uRYTW0+f
3QG4KJQNHtZ5KSp1D22hExPoDWpTa7MmYZNmXQd8H9ck3I4gErenvH2naHO3U9YO
J9mXQAnGGf+SbMGlNJBnNnxTEVQrMu//ehk6r7yfDB52d8k6x5wINkTwUtgrBJmR
gLzfNvy3qlvVxjWkWOKYN6H1B3mDqw2tGs/52QF6pHbrWTK2/DvTkmL/Jbh4Jxmq
/M/xNaMGy3iQ5J1zQPQ4oWAvKDGzoZFR0BHrAnrTHfHd2+HD4nSGUEWZtw3o088+
7VfSuCX4bNi2uZy4o1vJB1BQGCVarKhohWKY/0CnOaV3Q1nTniK4TOCT7SuN8For
TsgDenW7ahtVVKTbGxuXKYkxjglxaO8N5gcReAK48w/1oh1XBuaB903zQHq/MHjP
0+gIkc9hZgpVemF6SC86gz84YsG3/lokUU0kdqR4/GMvI+McN+CgaBFWZZSehZ6r
b2RnShZkxNlJZHz+OtIqFeQvxaW6xGjMkFJ6RvyfW7pzOHDZVxTYuoHF5EwHQlnm
3NyuXqhzBVmVkZQJBC+yiJ1StJ30y4d4QM0WyBW5wrc6YpK4kGJu3n3RGVzGZjr2
uFi+mtgKCMYBuHsK1+Ylp3Co6zl/8nYAlY8tm0BIuoV+Ds1OeQO87cXw9ZDG0chE
m7Cln8a/wse4S6b1VIr834Idr0B2Fhxc0pUOiJePAH04DTijzETrwvKf/nTNIR36
6ejhouea+QNlqqRpXoYQmTWqZaEtucFvLkHsXZSr6xvLsd67xwjAz7JLWXn5UW9v
l+Jmh0e1QNeaY3/KkbcQhKOv+5InATB6TxVRYNRxclNbNUGUCF+KqkKHmHjQ/6Ez
Y2IIAwVklnaHleLxh+WeCMfdoqTszLti4Bn87uGMxnJmV0G55eMIvI5akYuEjLwz
9zyQP54AN0sOhwd8TzH/83alRaLBFR1+TS7RFrZYvRq3YB17LSWMT3CU2yAePxB7
tk06C6kBUzmgSh9C8hBUB4B6qVZX6CJqiLAHjRi+LI6pdhgzF2fgj5rojTlCHF9m
IDgEhTxSZeFuOvihiw+z90jsEbEbklwikE9PGAjjalB38Ss1oMCQD/yh3y+afDu4
vJS7CI1keAKvEW/3QfnYnP8Nb/D97iQsISrHLH6q9iPJd3d8hv3GwyRiadvuI9dM
j4krJFsPko07f466RBP6MoVq170aF/3A62gzLy9HP1Bq6cUfiqR9b82i3m/vY+aM
5tQetZvdBuvXPPKCfHQGeUG6ci2A5qyrNRWbKSb67fOnQlwaCURNzMPzRyQEtevK
dY/tOjNjxWfBDAhiwJmziS91IYho33fg8ZLXz83ZA011x5QCw077h+toK6QFU5Eb
QFi63zy1n23MJPZuiTgU9EG1LrgyqY1b2TkGtRYNojkhiRVwPFPUtxW5Y6jCBufA
CrQ6jr4k1AntqOCYEkXkcex+H1y0uh4DNXktufiHpA5dWcqjIDSm2Q/Kl+FYvEOq
09jFdKdRxz7zFB+vmR4U3fILWhUrrUeqGrH0DoTCUiWCfhOOtX49kywVpfmh6h+j
XI5mShIaQ/jVtvsCySJeJ4ZIZLuAiLMdq09+X1h6GGi7M8utACOVs/g5LtdUbe5+
Y567JiSbl8c/QK1giyphh1hO9Zv+Wd6kQiS79iQt5TJj16BJAfXOD7BQtTU5/bo6
PEZ2vpSChm9zUejGjLYVF8j4KOHPQLVryZAiABvqGX/fxfYKmDG1iVObYuaQgxA3
hUbt4oXFgCOiRROUBGZRyqXnPgM/zWFUFU3/f2aHVtmpzY/4ZMv1fOvoPdqM4Pi4
pbMtpq0IxylTaApjd14cMXZU/wGup2Mhirur5fbkdeOY13rFt+bkM3pQJrbwnpV+
8FNFVsbthX6CPNtOUHxDKKYHuyOTA2y7RKwYsU59uW9+afZhb988uKCgqW0yoyqC
BuWJjoItEYuVTLiji+vquF8f9bglQNdwC6myUD4Vn0VsrFKa935ukPBzvacez6ao
jLPLw/aiyTU3OYK8905t5kPnWtgXDqA/P3N6NhTql6i05S5MOVECZFmZ4qWYkjUi
hMl3vJFPg+8ad7e2w2LBp1v+jZySmJhWklkj2YVrQ8m5nAje9JZXFkJGi/7mHQlo
FMr/rTybmTHOdMc3TgSfYW4biYZ19k66Z9zQlXpy7fMIkFoX05we/A27aeDUlCDD
LS1IT0X169t2BhtrOfvGLaluzOG5fDTk/G8aCv3El21hrbHjpOUGGyi8y1r9iKJ7
Dbpbl+q76ofxYzkYRuM1Aa5ftge+pr89M8XvumRsSZP5QwDsvJUYm+3RwF9twoPI
8iv+mgqtWEyC24nN1CF/+xPkdu/wsyZZfAhl+yZY4E/vtQenLgG6hwgZ17KQ//Sf
TyY0y64EsyiVuSL+EqpoYPV4AN0ufFhX6WWp1eB/DLZEN9Dia9gmyPFjj7XtjkBa
6ATWZiYVkeIw2/xpXWRlyzX53Tbr2GxdK7pVTFVkNH3R0nLObh9JPR2SevUVlM/x
Y8D+EKmP117Pk2c6N9PwjcS5yH09oz1TvBXJlgBJnadL8kG1vozRSyJkuwCIo/xD
GBa3f1LG0scxi73oUaWWL+ISWMtnUjid9R0gdppvCLSRHTxtKhJ8lseBj+W7v3uH
FB4lmPUXP3Z3Jlh4XoeQxXIO3svS+1UxGkYEbjCA3xLi6a4YFLXbIXMQ/Z8AjBtr
JsbiWBZMi1CGYbbJFOcYl6uRkdCX2Fg0b9YYuumdw0ZxtMT2meqiRS+BoRxMotY+
kTK9cVzydxeEDXYc+Y3dlOcXMVzuKG52Wd3W85jUodyYEexHCKXFTYgVUINZL2Da
WduZ50IdM3bMoZAW7NjqPrDTdZJsCK8QyVTybhmhT5+AMosH0KbLYkW/AyKlMy1G
kQ7G4glXJ5suEmmho5zyvK3ARccX6G+UindCnBS06jwmIqPypq6ZXj8r2nANSrCF
pTVhRitJ1c3eAP4ynx4xhtvnDM5HBcfOvuYb8f6UfNUsa+ZpubeSeWuNf3cxwJql
ozdhDpcw7hxcPA9K2MF6Ro8eLpoif1R0q6LeT/1pylRqNEI+mJ2kNT/yE8hh8IIE
Jo0VkpNr1k7fUlHze2/P1+WEfRaQqX0y7lWwRRP3sv7hnM11P9dkGrhcEybZnhm/
NA0uZzky5COCPlRNc7NRT+YGerd5ziPbkL7tGWDGaq7IvBypS8LBv/XZtsEiWilE
+1c9U7YzhUP1dutC9+qyWrREpTpG+Xq7QwEM+1IS/HSFUuvvlSNYRnXti2e50tID
6w1gnCB3sUQQH86MVUxW6I+2XJOYhieCCOBZWQOt9y3PK3YZByQ+N8itKRmMecmL
qPF3JpAZmUDNtWrFrLbXrPibzxkNEGrhnvibZSbLfRd10Ab3/aitdsra9Yl+YbNU
X44MkIT40JwZmohkXJRIZ3d/NQN1HTwkYllOz0OXA3D1NhtSPc8KD6crM/A5FGSP
lJQqyjyT3A2PWW/IhA6kBMLzA8Fu291/CDFWhSpuFMeDc0IPk9+lD9Dz3sdEdlUc
//tdnGcoJimZth/ijoRbQVeYOe+QuV6r16UeCdlixbtkJE/+43pOZPMbiqc+WFSv
1chbLznSicgqo9VXPVmehpsdESH292+08ChrCrw5oGw8Kk0LTrqb1Q5mTKGv5iHA
XKP72NsR+y0JebgVplchKA46pPPzDjjT6jsJOhVK5VPjsEbGDMiR6gYHh7WCeppG
xhOHLkNsp/Vqq41KkO2Be1t5hWpFbvNKAPdeGDhFoeEEidaFwzX67cqUydGcNUm6
PmsGixCbSsDA+Np3tiupdLeJdry20y73mlOWXk9R1YKaBDGlZSmIWYMlTbN7wF/p
F+WkqCSiX5zbzmbQDCo5GdiIkHJKQsBH1R2//15TAei5vxc90vk45lpCjHoH3DPZ
RoL5PyoYqTptNo9a4FM04lpZdP048n5Ktx2Gry1WrXHWbaH2PpCjPZk/9NsyZnfL
4JRKJykkJiP5PWsFmAuYdEOGE+8fS352fD+tuMhNdwFVxSZDRFQGyG5BhEREHoBn
ym1jrR55y+xLRMHuPbf8/oMxbFn2rEggSkCNLmXhn9PUlHkjefp4qS9+BxKVG8Bd
eGx0baNFMF5TbFYD9iTBtmioe28uis3Kpgti1gqavn2yiyl5kWWEvNr5Gqbz636e
aA0scjDNp6uXq0GHoB/jxTFRzFrWWDCHCiY9U36eXQYbV8Tavp/zGLyCLNPEvm6H
T5Jy83qqTZZ0Np+wFgL34LdIy50ztp1qbhExAAZzFA9plaWrvktQfJAmN/JiatyL
KuVO95R7N5JE//l29PG7moU7WaO+5a3I+DSWzBv9g+OBRPajAD5kyFdUCnDr06ch
uKuIydzkPIQSXvn8wY1kkOsuW9+1wzHbbvzsbeN5yv0ZsWkOa9atFEH15spREnAn
Rj8XQvbnKRD1HV+KYkn8U0Lv/qTvPzvtR6hrEYH0DASnCz73GaQGEtCYsrzAYpWU
OaN6JOmySoVft0InlUE2vNuZc+j5LE/bweWkdfEPt78IheH+WA9v2nZgFGtXqBaK
s38l5iOuaB7paNcDoly6KAvnVv4Q0RocaeFq8aGzhlKgxUsR4vSjGWl0bJDS2WvC
rD6D7ZVlACpzb4f5k+dfZdvrW3XdHfM9EHyRHf5fS3vj7r6n/t17SCDUID90TL6X
VNWEoPnoo0padR3cSvJpdYYtbTREEayZkQvhJ6Mvx/JF6/6IB91IhpQDMRfkPT+Z
VtfLfowWlg0kTF1/eL8s4AG3sEGZjpXHvBtuceOm6d2I+72DhHNSq540bu9nqsVV
wzUaY/H6w18C/iNCadeDHiMbZHAPIFcPgJwl1f38kqtdteGHCE2Jl6p7dkbqGN3h
jb7/WoxnLKenWh8WWdk5PJzYf679dGuu+zNYBF/CwAPOt7gdGKU15Q7IwVmuPgTs
yi/muL7F1JLP2mIbzHz6FF0CiePw0D3NZEhRQ9MyjppFh+QWE/3x6+RycpB+SSbl
pWo7wEKpAaW7lXpGHQQTSBpbHg7txqD6awLLEmsyGMYLU5EgX1AjKzx4dkIVGFiy
Pkr8R6eVf8zBIMciSjo1UN1WnVbGbkDHSa6ceg7DVaUb6SnclkkYRy8UFk8JpZZk
UY0LlM581cu5N2mt1Ag3Q8uPfrsXMHL6veGbyduBKxipuIMPE8lkbVwNoaLqZI5i
FfzFB55/88L0TGimO2wLOEq5kkombVN81RNA8j9P/rVy4b/zc6cINS7X0m6p2/Ae
2DpzbE0QpjeacU7noc6XAAp7RzvdtNLu2gZyOu6m9t6xExHMfJ1ZneAz/i55YZpJ
azhPZcdnLHNyGz6Ta0rU3+oiCsGulyIubtXDlwvyNvN08CnFo353+ZtrrIUQHYYb
tbflfMdP05Vbnyme1gXP5jXt1vBplIDKyd55SUJUha4JIHrbvVY1itnJuSQRhNOz
fPzC5MVfZIC9LQfi0zIsax87BvlDd9Pyt1xkWbO6iECxffva7kjwXgSGI+u04y9d
SbBYnPTFsgW95T25OukU/334T7NVx3qB9MxLHhFNUO+qI4qX0HqbWNjQxJ6TO9GK
CBeh3kRF4ppc+uEaHMFWfor01jxJ3zMpR9/JLw5c98uhNqCNmQCkLKpc814r+p7F
HkQINVQttGW0kPpST7J0zTuy/NlZFJV3lKquOy+3Wemj9ZRb5Y6qSlIAOm7v0cri
fzX2QFEaL7mVzJ/xyvv2EC4Ojk7tME/mno5YrKK4yfidp//2UgS3fR520eg+r85z
EgTyze4h4XDaMDkUT501CmpRHZfrwtiVDajpju0xOmMtUbZ2ZJf+AawQLF7UyrAo
NODHCbWC/Ms8FQEJIZS6uRJaj9nQAdPvHgFB5u6QPhpjPFscVhqRD+ZSemunhTNE
3uhyfAEVLLWLac60m8W0sqrhDy6u1VYnXSPjBjHbBgxSSIVFxTRNRznwvxhPxB9W
3d381egijRbz/M+5Z63Uo6uIsfJFO+LkQVI217SYPN+mg5AzWGrlVMKASlEUJ+1H
bcl2VXP7K5xd7yiMm5rYmUeEsSUiKbdlAkFjLagh1hCpPjnNxMKBopI2RY++X8+8
rQNAztQbHVdXoH4z4F3jNqTFHQsK+WQ38e5BE9Eb6qlsjLaCcy1NHiQxKpgXnzSE
LuuxjMaTUpygfp+EfZsZhWHU9yQgIjVafAElqs4Nx6rpIjbsI6oWmplDhuLlIYYa
9JagY1Bvos0WfWgm8l/T2Da97UOs4qnMQh7XcNLIuaOamWKc0ueruZ+BUFo9xNxz
JkorJzhVM8laDWGIUd++U3ODiJprg7VjYjmpJ+uc516vlV5MagLY32KoTnPpYE6v
i164/zqTDrTuq4w6BJ43vfpRFsiysrgQkMnYkS9cykZgn4QGn+dn9kh/oqJ5j2Um
LZgZZU0p+crgxUOMSr3YQkL5ET44OOokW33Qjf9c6aUm2zNTEHB9rgUOBhlkBm6r
RzbxUi+n0UiONgwaimkxp/M9Nux5PcrwMHeypre0f72gHH2WBPmtzQtorfE60oEA
MW4VmisH8KBzg9voP/6Zut/rWi3HxO/SRnLQp/OjLK/Fml4B5qCirCpNsWgLuseR
qVgyBv+yeFiHxH2dN4K1jfZ/oSc/PYtJY2YcahvgVZJ1+amswfYLFIl9aPJ6QTnf
cLuuA1MoxVuwhpsEJBdVP8iI8hjqHRA1HeM/PRzEvE2idX+vmV09vsMMGRr+M3Pp
0YUPYg+0AZ8xW1PdQaD63593MOJx6I2BrHvKOr1qcqWtel1/NiRToZmxOwrQbaMd
LNh/jcjdZjonJF+VXTXv9XZrh+So9fAGGhGfaKW1T4bTt6qlQbzAHugTKvWwRoGK
Mn5f6f3ehneUwgC3mtINSPwDDeyQymiE4ln2JZGRPGdfLYeG/6SCBCv7LrAXO+qT
Do/tJN4OfMDwpjboAys4gq/3iEiufZUraI171bGQq879zlNw2TLH6vCrWDU5Tl6O
o5a9CYCh0S+tw0z0FcMZEtZG9yRJafdq6J5O2l4p0PkKnxXEITXlZF5/7asLyaY3
gJb1/h39s6tMHRiY3zmgR0E5erbwoOwdgxGWhNECigBYaS7p8QC0BmB88q2rGgaY
F91kYXlspsX25g3NstsVInsN8C7HIN7ajT4nmxFPFAJOmKR6SENTRuzw5AFOzK4v
rXgHjMFHc9+sPb4bMjqUMNBsRKhrwM9bQNoueLAZ1x4s3AXVGBh78neO8ZWohuLx
L5GnIjcMU3SDyTbQbxeVDVNKfqX6U53wtV3YphbhUjeETdkxRtTil05zpJ/wvbt3
wEKwMAzon7CfUtELKvqgKB+M1xlK192vw/yvLBs1iDfyVxfZULF2JuQDuEoOiPY3
P3NkthQNbMezBCArDJfHlzmlVs01Lv6Bn5yAX68XD6jW9zNFcP6tQMuw5KaUXNlS
MkrWNP2O392YiQrQxzaEPy5S9cWzf6S1UORUS2xvDpo+rIqVQNDANKlc26zhIW0h
ZJiXZYjMsX43lguSpuqq8Kvd9DQrYJIHpx1jZorr5owAHJQuIS2rji3kiYwfqPuA
x3m1t/rQ0tm/F2YGLRoe9+RgkR73IF8ikliznPbqKeifXBy2SIouu/sSBc0nRccJ
PQReqdJx/Oc5tYes3C5iswtcToZ49y5c2U5P/aZBkRyXuIY0oR4OVTqNp+zTtOou
QoDM9iG+JsvQhC4G9jXHm0bJaxoJpsTQ2aMhkBn/W/Nh3fTQodwUg2HSXV/Eh/UP
9yIn9B/KNEM0jYC5/hwzbP4/A8fEpOnvslDRT89hwj+7Hry7FV4OESNhBK75S1Yj
h3nQJ/Vkf0p+WLxuIuM4e+gk68Adb/eh9vy93pYXu4gGF/sxK6hUgbmBnQvwS5yE
NPIgMamhmBOe8uer/PMZn6CaIDqjU6QvHDflxBavgYzbOSO9gth2b4C/taWd+RPG
9iTp0Koo4uI8RSy0E95vnnHU/8yvS4vhe6QdaZrTYT2wbgOO3jWhnjmahSLE50y0
g25FSBSoJFgRh2szOCmp60OdFuJ4noH4bDEZQIml5ZncD0n9k5cxeYfg+eQCREcR
SdA29G04OPKpngSQlbRzPZlG5pAHv1sBGUlhJQLN3NNQL9O/PxM1VSPH5mlSgEVj
UEXqyrZXbMHowt5IrWa4pQZHJIgD2OkDz0XXsgpI1OxxrZb6kJVMLxPo5bXJGlaF
8X+UNO4SNRHjVgpvBC2tJpZqzS3tyzL/ba6hkcjDCN7CnAHi0aBGuRPAOjoKEY4d
fi3DSoik1qhsEstoBLCtoXd7CvUQ0wStGlqjCkYCJY2dLw59ElBgj/Eu+8S8AXF+
Tc4fvDZ0YuMFA5eG7xjQ2y2WJcl2VR/IQm/yOptKI5Z0DgJh4Nb6VeVHIlguW9DF
0x4dVrER9PJBQ9ZeIhhxcgKBs8IPb69kUBWkIVqIMa/hobvgUNyDKALAcHxgtTXo
k4YEHySkqB0Y8DbdHPxDrR58FEaMrudBhhcBUKqRpfkFngCV3HThy2+lvsLmSc90
XRbie1TGg9H5iL18OEBPTt1UPdOPqNeCCETvYadRyZeZdIw1og9vEVYUPSJVsd1P
a1BLcjuYL36t68sM8becyFRefF+qsdC6tRxm2WNjdEfCV06Z6FwAA5fG5JxLXBE+
ALSGloOV60VhfYrBz2FpXbO7zKY0+kBpckcIoe/YZ/zjZsBsHCqPHPN7z2lGgTHT
ySUdavbheHd1MNq99S0vM1R8sWj4sdqfYuX7jFKIY0oQ+B51CRsHOkn5OZUOuVPM
5clDTx+UyE8YNxd/WD86lCe7tPJ0FmOSG1p5XHlET86vL7DKW4cZ45N9ihx6Rol0
g8p5eRgOpPRUjWdpX1uvb6sd3qFhzbXuTPBjkvmuulOpXqDfQz6bpD0qdPD+ug7E
WGxUHb67IVC+v9yL/MtRs1PpiTRqQuGnfi/u1HUo7OZPafxOf1L0Ade/0kGOy9Nq
7fKfFOKvOKLa9oyzuY39bWMlNIG0doTs4NKp1yr9ZaGihM02g3bj7AR2Q0F2MiR6
7VxWCnN7OxoleQG6uArxNZ0E6/0dqB5ekv4lyukqjVpM825cJhwEPLlX+haVyC1C
nu8hhEBb0ePC6SfNL51+b9kngVVqKYlVoZfGY0ude3VDV6uN19LZ70iMDCgpHIsL
XL18qqqZA0fQa+f7bkEVGqB9K4bZ1aOmqGiwJF0ky//JxQbzPWwx/gRvzLzakepf
Ph2HR7vLPNUV+QtjyB9GcRWphd8etF7kJN8FAkikW/EQzMm1jx5z5byhNM9sSIeE
QJA7JdTkKVoH5AZKFuL7Kjy73dkP5ztVPwxMZoalVtR8Ppdpc4fkovLNkERi0308
aIfyhPOKfFFBrH9rvPvMltV8A+fc47HghXFUMSqgK8zCXGbm9Smgpiymf0mQmSU3
7EA8i63vo7qSUUKSJXtKgGd9wlv+CZ5ImVMiQPLwF+z8a/WHnHL0aidSCkDn6T3E
Sl1gPUG/WBkumqqt0ioLE6odmnY0KciGfe59ymwmJxk3iYAE0FCN015sXi6IYDNV
7DXrHT0mfntgnGfG9pU0lTcYs85RZQ6bI2Nq5b96x5a+5I+8stRf0AWLitNPX9nn
3u7lDPjC8DWZVM4b+j3+K/ZEEGpZb10Uh9rRbTSEe3kok7iBWJ6BHNtBTL61fF7o
XrcSfp+09qDozx85S4pZIuoL3/UMKup7z50InDY0v3bUTsYYSYw5PrUaIEAkKub9
jnlQ3lN/fpwMJ2bQjky9c2WKnT3HqCZVuYBgsOfUVptYFsG/Qr6JMIWxUbiSfoeW
Aesq0fd/g6olAFHKqzHaCY3e4YxwQKGw48WKE21V1aZSOleLp8lDp+hjmRNhyVu/
j7epoFnlj29snhZxHhz9dOVwdyYJAsyz3HbXbTHGvishzsoqvXu8cTBU710wcZWK
Z8WRs/ZQiw5WILcgvtyUKz1FWTY67nosiHF+KMjBpg1W9eAQiaPAHkrXkHQmP3R3
WsUaWa3ixaQu+ORcynmstAwTFHMlrLCFVtYl/lpoOG81+8rkuyqePq/WlbysaWkt
XX1x5yNLNCGtPsLfnlyAEEX6GmpL1OsHXDX8KLi4loeJuoYbmW3bTtlhHQ4/qTnh
gicb47XV3lprTXCeyffsPa2W9ndm5zFl+FwNasVu8eP73DzSRI1k0AaV+D7jkzXh
aVdr0TGFJWjJKuBYoORjGuE9waw/3J5PSU2KTBs1O+oiJDHUwXuthOFP1QYt+27G
B66RO/j4kzgzf84gWrPl3JpG/HYxSV/CBobWQQBx8orqx6VQq9NrH0l12rmFZ2ID
lxWYELq4B6AB8CaQfNYGh5+KpF6upN6DeuhP/8AXE9fsFvdMcZQ2ygTerdJoII+8
ZY6rYcnodh58tido0TSPJsYbgDtxnHJy37iiOSj4LcrNjE+eK7n0bkHPx4LMXpjI
BpgHlUPZwlz1SsMx7lENRte6VHGJSZ0UCiLLuIHBXtl5s/LDeQbA9jKWOi1QdsTP
Bz1EwcmwBdJfK95Pc4RTYerzlScnj36D/cZli0YhN6lW5Mq81SQgoqw9iZNXIdhX
3b0I6GZejFCGJ5N00s6GK9dFlpCBVYm8+csC4689wOjHOCARCbsvE2L+fg4OSrYO
HM+PR1Mr3coJlyeraIuPwhweqo0bx0H2fDUxqMotQkmCWEdmV79mNX/J2/BF9McD
c8s9MwH/HWijJdaHT9n6K67mFKNWrRLLmZ4bn87Z4YhgOqA9NxiLvlYBnsxahYh1
lqswO2o5EmchMPsvkSODlMCYIE4xMcGC8VtNTfjo0RKDKDdCgJ8E8wg4FW0oVckC
6xk7FaivArliVCRNZweLz6Lr7qWGUqkXU9Sqzkzu0gYHGCkIDEnIBWs5D2OUPeWh
QbDOYBIkm+QDUvAd6y/21t6dwaUcGD6ZAK5baEXQqF3z7vFCE2kWE507DP1xbUaj
1yUgW+mU/IroknDWhtZk/7OmKIDeV7fViL4JMsUNxF2FK5nRgoGNSsae8+R+6Zau
wOFR4vdoVB8aXErF9ZNFLIUq9FqtDTsakGTMfla2JTohHlXEv1IrRxKkwRDNAwPp
22Uc0WW4qVd5sTGqPBYmMThtknXgpXLlYAzxlj1xKvrw49r1U/dlM6NGe6gZNnmA
D5RJO8bcLNhmrhsD8kyA+p6T94MQgBo5B0B5UT7XFB7ZX1WCsuCUBE9H8CQHTrd8
jA8w6btnl+f/JihSs14pqtY9J+9cn12SQQS46ZxRO0srC2HXMgCaG2G8vpcms47e
rq6s6MuV4Kk23gaYykUrKFhqZxW5kSS3SwWTkIt+a1XX6+Vq3eXmbrrZuLcwn0oN
nA4NH26Xv9LD1cT3ZjNKDB5azywd2cLwfeeUxLNeUJnva8oB2hJyHvpHDnvyeYcj
rS7490/Sd84hXCkcO0q+qdtmprmBH4r2Fb7atJ92+KYPNXB52+EpG3D2b09JUGCW
Zs4Zynweq3FoxsRY78EGeHYXTO1wrZhkDdMQThS/yPthawnjyQEyOrlWi2UP+gE8
fzX37svsfy9dwdCqIXR5OADBhti1jGFByWbvt+4JA4/CR5iS4eL9lF5NcjUQSB8p
NClcrpo06HPbiTxg0z2sIg2ImMgltKZ8cfozQkh7D3PdfYrnXCPC8hM44jCgoHlY
t4DGJtlivGiwRTmQgGxhiPyCGSIBwPu5DWT5MVC0V4CSb93D31g23NwexAcbQPSF
TAOigX0yrOFXISXLDjQVXhYwVAvvu5nj8e2o1fDsW104P1ltTekW/kEnZcVGQ29Q
bMP/DZftEDux1HdIFqaJL5pOPkNJp90kfzaQnsaEKx3Ahq5f5h5SpgKL+/YsKvVY
tZRypFLeKcxLCdPOZXgi1guLEXEueAHsm/7xTRFvnliel8cOyAWpSlyPgPjwRNsA
cq5EU3iUbW+JhRVOAM1OmUSPrA7b7QftwcjmCBxkJi/Ffh6U7u9qGIipGi2T1MqQ
xzBLM2UmOGGjkg31Phb+7I9ivj+KC/HIDez4wTxsVrvjNchyVIW3ZJtxA39h3dPE
VY9S8+7I2CgZ3R6OawN6wJ/DrG5nwGBP4frCCkwUMGA0mH3xkOr6gbZdO9i4JY0Y
zMQbi8vC+wc5oUETxsqlWsSwJ6mW/95HotJFabUo3N464k8TTg0gOzKDksoX5RRd
weKyeNkuKXITWndR1T5H1JeaQkPXcZ7CvRShc4Hw5Q18YkVndiIGxBWfMxSNBK8Y
D2t3cZfXsO6fEsTpsXh8UgRU9nmrlkT4FAVJb6TjE9E9Z1H5GF52tQ0JJy1fpVfa
5e74lslPJa1oOYNnYD9whHuc9d9hjyClPk1KP6MJQH+buf4wI2822ts1u3qaJgiM
xLbkqL0nw6rasmQ65/Y/djZUn0Icp76L2IBHG7lJtErCTg8l0wNEHw6UDrI279jX
Nmj8sfjhX7suPbaVB15KmdhrGFbPPYHO1gIwgMYydnMjKWNQ1lfo2UlE2/yARTCd
BaxeQ3TK3fUthTpW0f2cy9VJb5SaRBq2VhF4JKkuH1Zz0lhdQfUgaH1K7mTO5yGD
dDedT0KunCV0kF3RXBFAOGcZ/fLibkfu1HG+WWzK6LHblxzaG989ixqP0qfTBpUB
QHLJhnW91ltuepurEf+6aIVUJXg4nBjB2dVz/baJY+omXN7tVxeH5XTcfscRP43b
R3FldCzwlj2uPi4CJtmrC56H5t+0FhGKxeK9J6JnThmzmMWCuDWfy3MW58gMf5WD
0K2pR5cauFKFXftza+Utsu9zOt6JdoYvSN5w8JWHokBLdiRIIONH0ZpKQLghLwKS
IOwxxI2l5qI/vjnWYqXjOCrAdYiSevk4V7tKvV/Eb1T5UFOdJrXbWv+9B7Kwy4UC
yCbdRkTmsLYwvUMVd2FK8cvolBxotMaWKjW42taU30dCAecjdwFFnJjnBExEuY04
oQ4/ebF6QadMdG8U81FGmLvS7padKivGa75O9QjuiaoyYz0nN3BcPv9SYMbQgFMq
eUZjc3qbXCPbidpLKRxkQbiDbCTi0ZOQ9Fw65BnGrbBc3+HtFVUvSsVLsXLlwphi
WVwxD1Ex05Fm+BOnG+/y2FvnS2mqEJyNQtpQOxh4vH4wgXqzJEpHky/h4b2Q/nYq
cXcJEcedKhCEeNsjpMrEupuLeBFNSd3D72+XmAvw0TGnaGyJuw0szEtok7ZXKYT5
Pte5ZGCMjmiqnCaVMkQcLOyESXlKAs/moPUMUGhMk3joXhxVtRmRoC9PtT9Bfazp
Ba9fJab+e2YQ3on+N9beJikp2UwxdmM5CuxvFwnz/DsC1EonQfT+AfYtkNHn0uzB
b3iJrOZ5fz6PShPLR/eQ33tNXrq0x5EbgH2OZoY7uRKlkcH2GNzLM30gnUigmINw
OqRnAy/J3oudgunmptaquovh1ltlPGgWZxifiSUnPa0nVEit/6c/NGKgSaUvUQTQ
8rTrVqpQNdhZrQiPICd3lRA6dFFQiLdkMRw0bAIAKovfgONKsKvn5lDE24M6gz9Y
99yki6qHaZHGe7Out5MaFH6by34bBGRNsK2JDzDQ6eXsnDp/DmrB5RJBNGbcTmC5
fnyQ0wqd7+JAKXtBD0h4iOHQrrtijX2bxt3JSRr8hqxNFmEeH6a3SdC5HQOLNwyY
hx4O5IKSqXNEjGBNYROq8etoSPpDsgTHhGlsjKRfn64eNMd5lHFQqnxeULkTGsjU
L2mrlJwLYMH+1Ged8rC8tPYJEJE/m/Q6QGloWHQkRp0ZzKbWqjHxV7XmhgojjTM/
OPnLDTH9+EyzI3aHLghjB9JQpsO5kqG387M48kJJ1U+dt8xv+Xdl1dVQr4qcXziT
o+0j8/9V0sDVzLjEe3sqnF2oolku0ZdX9XBRKblEPQkNl3IME8nx/tYJLN9Z9PZB
CtU50BQiFW2ON0vI2zheRohNKba+KUU2zPRWyc+zFGjWLu8keoB6FqOcgPgWkn5m
t2hTGE573VcUqa3zIPPi0BRNmIWIawBqN7FbWYej4OmlVzE5c6Wi48ZFKac9pa7l
7YMfKJu3tDuiaelZUZQoEH9PyIu1mw6gHuH6q+OocG7oS4X2e1GvGuoxhs4DKPCK
iWuzOWmC3SMzumjUFh58QTYgEXYYYOhdJ0yjJ/AgzypGXykOX7+FI/gNJfwjcQBV
6tVg5bSoU8S8sKvPIyyMkGRflAC+qqnWf++m7h1+ZPfBLT9dNkdfrIj7U6FW0m9d
SC1aNxcuneLOyJXKvA4ydmw2GkAxjEp/aALb9iunzvOFY5SlSVJ4rMJ389dwDM4T
qrPTuKjSLPNIYUeb2pFZqT+2GXjwY+cD4IOtFZEafEaSSrIFFTEmZiS4QGrxYOGi
KyVNEEzw+0uhulOqfFlf1JxMWX0GBY5bZDU0ZjTgRiZcjhqF1tQoG5urMVdgX9ua
qw1Wms7hUuao/UhuBi/MVlhnbxRSR2O+/pdTJwatI46p3tPUsw/NK7e0T29/OehE
SC8iIlsoSQoJMfPGZLuNZSqLdWcKJtw5KE0t6x6qa380cRvlUjWV0Z8BOyPH8yam
mG/l4PfVwm4WSwPVXhGX97F67opKWDqVXO9/1eBCJ7AHCRueZjVu2NspShZ5fjqo
wGWPLHolJDOcH9nSuhRlVwivp0ny/PWPUvKxrbul/zNmG6Og22pPXMnnmVJCKwwk
TcCtDch5mY1MWy0jygG/tDaaDT8wl1mkO8qWn+0xO0zRqcfg5BeWyTeTeJ250hSi
t/P+odtXJ9BI+FSMrvUyFRynWPapChnvUnY+NyXXwuS8pgdyioVVQV/Zb4ML5D49
wRZJDRgxCajcDTJ+SnELx3C6w6uaguDIMbeWHQZWz/yefF6Vnb6KBL+VGfdurUQ4
8Lx2hDseHt15xi5s39EJOvuMeGztL5uu6BYGzgwOSmvwnNbiM08p3cnL7hWnTlU8
rgAu/PtOKfvUdR+gLwrieaxvgmD892OOIxMvqIkSV/Muz230d1EFCF3YjA9HVaMN
u0bc2+ujmeXoMKCBypgjsrlDSUnkD/dhAS/jBBA5KuCioWOJKIv5C+0xQvGlGz59
eku+8nrKTFyyBts+7pV80R7XI6SB9zs37FvbkW2BQsF09mkzi6M9g3WWjW01LrrA
iGzxkSt8H24sS2+xOud2bh1n4I1CYIuxvSDB7XbWbKtNXko/pqkeImci9sZ3YRoe
Io9Io9L+W+26OD4yJVK7Uzdbx2oKF+v51RPeflEtsxjxunP6BWfyLVCvxBy8dVhr
TMggVWQdkudrjmdLUCyAyk+tJt323inDIsqrO4hGW75IWoXDbB5xp0LkAD8U4wMg
Ib/9keGQBAX7L3v1pN1mFQ3NY7WTlAV9Xum9nZwsR//LBFwRS6E+Dkd15ROHta6Q
zDVJELgsqtp6YAYD93YJbfqG5lKu9ej9uRtyN8MfAr7ezJn2Sdv6Ia49D62y0WVM
i4KKeuDbZQKTc4Aya9xEvNeNfWi6rjlRrdp2IvFc/onMJLgSZyxhzcZ8o1kIEwws
+FpVlwMu/+6u1BB+taDBBj6B6/BsQWOvpVktaVASH7p6TnhinpuXelkrcA7UcUL2
9dhufNmiZ6kntv9KPG4N0uZ2BrT6JfSwd0Lqi/IbUVwajGUFTnc+kTEPw9vN+YX1
FuSWGQXckb6I4hsuecrmbWXhv/cfAx5sqyEwe2NGMMPT82QheEUayB5L0iFiLdT+
xgryXN1hogHNG8fnHmRLuo+Qmrgql9AaSBz3L+AOX5jLdc7kmwhdr8s7UW/lvPco
HcdoLXH2EMdxPCT3pZd7vgTszmup0AdrPAJSi7yWqa7uOGrfCHTGyBWzCYSlpQfK
H9BAkVT4IXNgAOpiaiS3VA1nmz1O/Qse32ZbFuzLihZxNMjxp6JpRYcetRBAUCVm
rK/tP/f652NzFRpQZ+9BG7/akIGEuXt5t85mcBOF0nQ9LBXfwJ4ABji9omoDtZMJ
4BOM+hNH4r5JoyrChfcZGZn3sEP4n+VlJq+JLk28No+HtmbnsSwreu+/MZiHT/Hv
xQRpfPra74y28tVsWXlcdfRBxqnrCJOFpHjQwyeq3Tfd+nLW4V8D7CUwEwn6OLsz
WiDLymPzevDIIrO7nCxCYl2cAWfqM5BzhTV1HZOxu6h1EefsyvPPzeJ5ZQ4szd6c
uBNGT5/GrHXTtycvtWQjR2bHVLXTd4hLGO2h0vpZ+t48LX4cTYKhPE2AdaYaInqD
IqNeRBy0Y4ldmUs8ZJ00vEHQ/zr9affenCkje/sdF2669Ccf8U+SXNpIq40CBfLY
pteZdVVMBdU/PNN0rHBghhweRon9L+Gi0DL/UqKt+8cin85ZaKhXgCVKDnxjFVTi
PKTflc04cIwFvVfKp6fB0iBS2FV569U91Gbf67QBXf9p7Wa9VM1mnRBpwmKbWuCs
zmg8/dGhsj/CYy0+ERo1qo5ljSsdFb59SkfXaDd7nmNXfhKOckzDhW8X78MeDhbu
rjtm7HzmemV/Aj1VO87D2LYZw8eGQbAmgYIhafiUfHU12uI5bhMO3a0vQE0PNhdO
VNzwzIfuKU01lf1yJbuqmbnXIS65UMt4sBcutwV7ZtVHe5qyv+JgRHMvWVXTWZnu
zpNyztldTO5vP9IbUCA5tG1n8DCq20ZMgrvAtfLaRv5Ny2jb9vbXeKB21AHTlh3G
LmXdzdKUtf4VPe04ZQsq9nAhT2KtRz1ZJhUwvurS7Iikpk8UixO5T3pBYiePJP4p
0uedziOBrs5t29sz3b3BfJ9rCslABvVL3K4U9hDmhARgPf+7y8J9xwKJHxUvQ0av
shJrMjCI0/K+QN1S4TGA3qmfja7mKQAkpjZrmDmW1Tjk3f77otAtVjFlwXqNpF3n
VPQMO8hBfj/HhnSFnk5NbYsO4FNROxbI3kpwjbHoLW8K5B3UNpMz81E0tXimWKz6
UTbJiSt+/YO67uKjcZ41kDPr9CySqjweNMnaHJqcOLrEAp8ZYtdWj5l4rGF276qF
EKMTy2gcSkW57YpopSATpgIvoPE/yXRkl22jHbE3OTBE/VC0d28mf3hXDSuzfiHC
HWCfbWNhW2Iet2Q0V2YJXnK6a1dyYQl07oUW9vEI0S/rzAWgVjFPoMVUeHvID1EY
Y6EgtaUv/O/dl+kFDaN1HzLn7/P3TJX56zd2KPEi73rAU/rPi5LwgHc1Pzz/uf1K
oGKzDtsz31opb17+gEyTQvhv8eAS6uxAfgDwYTttAkVKwZX6yd7oXFw7Fcg50dj2
nkMWC8WEAZucy280sEFDaQXtLco5MuUvFjnvwPk60iTK5Kzczydwa3XgWVbZcAE7
JRSK09FfGx0HxzcARdm7QHK0rzCp1m1oq2fRfYmnst+nmnXvb190W0yKd/VbuP+p
6xAx6429dAIBbrGR9gQ1RIGajKwQPBrajSoEIXWkbBPmlgEmxZvMPKC1Zg9FKHuX
igrTdhzgi/w3dVXZeTFBAoITZTE8OEzEi45tLJnODkUJrI2uI6t7ceXGxMRBpbcC
yJmYgbMHBFhRoUcCsze+4md+fewq2/hDRPf8MoJy84nzg2njv6IvAXsuXCNwBxyL
03GlUIcDLe7CR7WwwbzQNzXsVhYDRyGSEX6W6FGf9NJMj69Hwx7AIocrSZMxZV9C
f8KFeVRS7n8sAj79GLuqcfRa3vzr3zCFPu0vQLdhVIe5nejxXcRRsaAn4gEHMEfl
ZHIg4GO3a9tjU5egAkrF1wgZeU06QI4xKyrHZmxF4toVNbFgIBPPUPFqKjlBokLl
5vGvLq0yWq7SldRaU+mPPGqYLRSftmxga60G2ECBnFHft0oQJ9HUOkxHL8F5Jjmc
MdkQebfcp8fCN95TYOsRcOFJCffjFRMrEW8rjYZTjkj71TYNPrX12iPSXmK/o8BV
bwWh+68mXvJyPTjQfgKVc7m9YiRwWdRWUtebYf5xc6XJgSI5F1icwZtx6kEhu6f6
G3JbwwNX541i2UX4fGebXecQ3/IsZCDQNZ3YJ6PdQuWugVoQ/heR8ZG8DVEpw74N
26hXRRAAH5JpKjNKVD4iu1qh8n1/rIHd+M1ywOgKod195e+xvsj2117tNRHiTgrX
HZjAojwK8tSaG4C/SKJjaw0C+cn/dbkSOSjSpemAk/QmVtX4CbIxWP0P4vKvuSEm
hRRUhDDv6Q8Fa/udevNojCXmzZEEj4O4qhwmyUfdTtQhTm/mf+vCoCIhvA03GpHh
1CQluKReCKLbXrFDvtkEBYKRNbsZUm8HquPQ9cdwb9foUhtGOqfsVWgWxsgGHlK/
1d3avBTn/T9OE+nahImkBVDAtc0VRWENj04HRf0Rc1sc3T9+B6C9UxdJEE3KnMU7
nfrapHED5h6uSut+avsiPWTycMCtMUD5OJZxEpoU5fCaeuuLfDxcMoSqr1C0FTUN
bsANGq4M+RkegRgxCQg7ra2LzHTjulb/UgeNQSAwQ4CE7cELz+A4MrRaQMXUgRsy
liUXybugF4UFkEmnl28wxK+2JJciKPY8JtQkom0Ha0QG5A3E4j2eE3iwxUUkAE5s
Eg9/IpLWfxHC6FRu05Ib7PGQpZlr80UgQQMtpiHSPHivZFbpEwB55x2FtUnCBis2
xWc/RJjklEHBgmxT0Z5sf4z3uJ7D2s+NLLos+6IWE1L9yjENYk1r/SMBGyo0ehlI
Ai4itW75InxJaRukWnBVsQQncxk3gJ2xbq+7KCwtq53BWpRU+m7P+XR1XPQFIW3P
AtsUKTyw/rKop4+hJbf0T3LiORmMd9Pxx4G3OswKHpOjMY75CSfUqRJaNF2fXl8u
nX+4vOq2XmKNh48FBKYd71J5iE3Y2v4L/p3zBNHXYMwZBCMOlui6CrLba84HHquA
9haOGooJzFwjuXC7jW+bU9dEBm4kaFFgonaIzNcV+luGYUOKdLsN7W8yLm2LqjNV
S6gQ3sstva5/i4pcIEh3sFMBHBwWhhrQkJgV4VxIyn61jiMAzMwXwC4WPE9GdqpR
Y3kvNmd2N6BiPNdo3OWybHh/bawGjzsmV/LLqJa+2dXhrVXwNm7nwBRTLkDwgVwQ
sSbnT8CnuuSjuQinlkqlDbidfr+NoilLKLmAR1zlQDz5DCBkzVesiNu5htBvdy/+
lrruE9dmXXjbYMffGxgIt15DSVluRwFXW6+FjuJxvMkN/frGZOCw4wAdAwtLvXkd
M6kcy69vn/1jEq1TtUsUTamjau2j5VYzrqVfC2D1Z9fY4GfoLuoebSM1Zi0AenY/
Xf7synSDiPoOQTPk5jLGkxWwEKuX2uSZ9IijJp9IE8X2shD9mHsZtTnacZUTKfJv
5yznQ6XvcHZggZ3Bo16yIfisPcXkHil7J7C3nKgFSB/Ofb1/ZtLAUKrUOB26UTTm
vLkB+GUb839ydyk4a1uYGJqcw3zSxcpnvhFwOOzCnx7KJBlZpF0lnghSZ+4Ehh7L
TMzWBwZUV9CMB/+gqEzHs5kNNEXLpPK5uxS5Q/JEHrgE19lz3e63BRwpfUDgsRQD
V+itv0MZzmMPbf7t3UUbzUKCp3PS19weN7c9pS1DUSBCxltxFK1MRAKyL+5g5hVa
YYg8RtJog1Riiu1ovDANkhCRrL13p1XlxsfocjglhEaeDRCuSDctHVMmC3TNlLa/
a78gyIr5WP1MrGujug5HawVI9xR/KoiMBn8jQfJcoiOzui4mbTPx2s3shW1clqD4
va+alaw6Zb02larKq7TqLCKEb3XI//cQGhQf0gQJkf86pzhbxhVeJWn4E5W5HNN7
u8OrQHxApfYR1HY1DZd6B0obk0nuphsl3QRXUiEX/yr1ZV911w1lV09jBXqjS5CI
FYQpy6/TZq4bRI5mZw2Yvrk5gVQxlurn7NV0PuHevQmvvKhZb8DFiMZkloz0GfAa
IWLUv82QL8OdoOFUUnqV+m96Ze9NC1XfglRhCjSt5b7Z1srgs0F+qzJ4JwGdb/Ug
v2CyQX+CvwqEqKsoYtF1gQnuktBXPuJGtrjT40CAozShAHSGkmY2bInQxCLYpJAH
GeNY0HvG0d1jWAKskSKK7iUhWkCidwfyDCr6yqpmMinNAZa5g3Qu+4c0LwoEzh66
6fraeIEV5jHXcLBlk9EVvApM+4qh0ewsnXwv6RHQnHbhQ3ArMvLHehE5ojasgnfs
GAacHpX4QiTG6dswgQXv6wqz1kQT9pwwEzRbXA1/4InQH4+FkZWSxENLQuwBUxO8
eYjfr5I77aTZlj8ehk79IZ7A8YUSF9FhYywA3oapvers8BJ6rZ8K1Yhy/Ofcql3z
HNsF6sjNLfes6aHKlreKlYTAV0fwxuOI92hD4GTSLq1c3aLCfSeHUTxD0k/y8g93
bpOQDG6n+W4StKpxNzkCqh52GPZUjKdW3cbc0ywemMDt1186cyw2UWemtDDuK574
yURbLN/srjSWJKcuC+AAYe5GikBI/O/jv1wau4SVx/RH6r8/Tk1twL0Zc7jtDL1G
gL5PYHlnD3yxClOLX40Dp7jCr/X9ekL0PsHlJpPvx9zteAEAE8Y2NpLKwoiv/T9F
Uzjfz4Xf84bwRwPi9lsSsNtZ6qpfCWQnjv68VnKkZ8/7UWUP10EbJXKVj0dvC1Xp
d3XTwNlWTIp+lgiLvTW5ETNZpp/iS34zn/XGinEopRCQzSzyjVJ0004ADVkBUOp0
mHyMPhSMZQm3Tu47YV6dnX+5QyB3YFa8FNK7DxS/Njth2CfPRUXla8DA7oOjiTC3
RMsoIPzyE+GMb/WPBqdfMB4q1YLv3iCihyIbNxsjWcrjsb1Scu5MJ3Lfo0Ltb1o9
Gq55g3Ooq5w1c4/tFxgbVgoit6HADo7Untmfp84WAE02Kr0dOurTIj+qDeKp226u
eZe7l+q99x6+zpPwYyGKZKDFVWDYZV7zXwD43cPCgWKBUUV2h/Au1Re5MGXAfXY4
6kVFaJ1Ew8LctB/Bh3lnzpcF8aTdgCWjjxlDR5AQHouV5X/hdlXX4JT0t+nXzh6Q
nr/noflNNRQ/EZWCd50NhRqiZwCa1dfuigSV2pdckQwVCgafKJtEN7fxCObRDYHV
Hqi8p7q2brDZG/02Y335Skzd40KbfxyLUGrSumwG83TZtwzG4lW0CTMhvNpZ/t85
RCW5MgKpg2tV7zVnrX4D1BzNqPNDESW4R4OvU4QmH/mexEaYnwPI1ecnsrwi4M9V
U6QnuS6q3Q/oV11rujRRCMUtLS2/SaaVKGZaJE/SFfCVC5+xzi2nvzCOK1DSJjvK
F2A10bCXUGotBK+D8v8kpeGiygKcUChaOIK9HgDoDqAsvCi1VKDlmvcxaW6vGpr9
NSZXtzoYygJ2klSm8FYDrbarDzZB1ii8U7lfMFr225L6yrBrxWL+zf87s8c97Zvs
RBahQvzCNtNWAt4uj3nXUuR+4zwe76/ohy01m3hSaNxIYK1pbmZ44B3wyRsG521o
qXbkc5LScEj2n3gMTYcQQSrsdT64nULyE2VkX035icQvG0eq/xUtrBFa4KpIZRt+
fyZxKT0M823aU4oqYBaP9LQtxamGNWs3TTQVAZEkoWWFawRnbt5Ffqcd/gCUvZwB
8RkFt7AX4n7L35Pdfag9+XgbPFWOTaz5wpYtyhG7os1xXo6jTgyhzdNhCzpH2OGx
uj+QcB/M5LLdPSB8iYz1+v9VH8k1dPvuEwkkrTOEvY9E81vw40wyRmESiFapujPD
JVRoHNIoOTxGuni2fjBuUv2CZll2MgWXIdTs2TR9sLjekYXajr7uvHpTfxSruqyr
YG1MljDnPxcTPhoxnLTlSsaSEOtF5VlcdcO7+XikIQypGpNGisSDo9QKTZYGfCP3
lLwKa47Q/Z8n9SNmbL4QxAqNIzJJxdqmCmCbJPCEhjd1LhZ1DjksKErwC9/OZPZU
Gl/VSEVe6UemtyOMX2yZQVqofBbkmv2YtPcr891ABFDLeUmG6Gygge4bfQqHIXqw
wNzFO0WphYG8nT+4llsTHnbcXNrD0MGt7bqk7iVk+YcIlpColpFgVYTX9BJT+0pi
sxjFzvsZAs0Gn5uO3BJoLBaUsZIFo9mRQK3g+FNIggJ4L/0t6kHgUmwXDuTfRwUp
eUG/OJuSir/nZml2Dz7sY6CnYHseWf5eIkpUuBzUYBr8jGVZg6nsM9VzRb6NCjRI
H6X/ynIH1j4aF3CwYt2PZJ0bi+IzN6/nVPXX30X1/F2pdwbmHjawLp9jspixu2Dq
KxwMpzTb/LA2xwfKZu4DlJNQvtxI30VDjEImXQbT5rl2+EsFgBgMJiWB38VJy82D
Unx4wPrPBZz8BifRhx4nEmUx/WT16RPhDRcZQT0/0gG910PB5dLPbLhKK9rfsDeh
FnvegYSwHJkXHVyRs+UHdipoKkBgD5NwOvrklduT8e3UQPsAlxT/ssK5C7krT0P+
ul3HzlBgbz6FpERScUQk/UdQcTsbfLlNi9Md4WQZ7TG+VBwGwmUKaf06f7MSALWe
+Ko9cC56xpQ19Q8vh1DKx83lTXGVEZFtmWoq3R0kYFfjdi2Uba53wVl2xUZnWreh
y/J8GeyLHXDCGyeRUfP/cTWoccIfUwfiLhxCn+RNpMsRJC+M5gAuPWiwFEsvvLpH
0bITHhmGi9EaJ+TLRHORuM6clV59Dfjm9/Jzt+PL/UGCar1KPHgJ21480mYp5sEa
GrkRcc2125kPwxff4ilf1pYvt1jPAnyhf7X6FKBLeW0GWcXJGLg1BQu46IkEnKLU
5HoJ3sXvg+SD5VZxoUqqSeuZniVFqbBCofdypSBpTW0nt0Mkk37jBYPPS6CofveJ
sGarQnTxLf0eyxBC1c4Xw8X4SCGwAIa7WfQRQkrZrQ+4kXBksu3sTn5aJ76OmgZd
fitLRFTUEX2goPpjz19EEBG1JO3YQSeNUZHtl2i0eTnhFo905ezmJ5AgDP+3KFV2
Vckx1aGkAW8ogAm2XuhKurtxCZYtYG1jtsGqnNNdZqsq+TSrUDVan9ZIR7I/Vilt
yV/+MHlWG6Ks9Jqh+Xq5uLNSL+tNGvnM7wPnLT7rId9tx/Bu3VBUZs+rRreai4G9
lLKkDmHBtIauC/1sXv3jWtIN4iIePEE1SGQedyr8Ry8WQit2tDbdMOlo+/IqIuV8
wEnL/wlLvHs7mHzdobKAuT1oCrkdwvJt8v4quCNwi5jWnG7ZEHzBLpwEzNHw3Jo6
sQEAlG2gewV7spD4UOb944/LO0t+HwsHmm4AmIbxjmpx2qKbCx68w3xCPAoeRo4u
VGtpYqdf8ka2oZLZqe175KFcmOk19Yfr4HlPG1CpV+QG2zd7Bi4jfQGelLDE4Ffo
vRw1CQMwK9G6KBkplmxqnA4brNrOYkJBhLa8lhpndqL8CwTY+7ov11PBZ6u+/rpo
uEyF1Ci9jSXdas6YHFYiaM8d442lcRbYT8LQHpLnayjvJ3UmEW3exRw1CsYIGKIc
7j0+K9UQ0DiPGJuyoNC2OT8AfAlZ7jvubrUAwLb1c9aQaOQ5Gs+OksKiKUfIXV5O
comeWar5/ouuQL+s1hkdhdFg2tevc+QUQNvzcmbxFhiDPC9GwCgM+jmEBZ2kXe7M
HVhuEboEsSuexSprsxO80sYylWxbauFdNQqU9DPlbFtaw7UzBXrDRB0gHWb5/lx1
P7GkQqjQpJupd1oDx6JVF1LhZm6N6AjKCMJTQV4K+Lvft+zT4uO1MY/Zjm3f1Flc
hO0qRUN+qLqltkpusWQeAPsLyJea2GVu6m1sgF9tRsBdzlV+EqyZt3V6CGE1wOJE
+Ja73t8FnfV2fwtysZObb6tJF67FtcTBE90G1R7je9GjdNtvVNQKxckfAsw+gpoR
T910Kg6vkz0sWe0uOvN9iFRaBU4lY5cpmLXx+QyDwPn3sBLrCxdhlhM8pZAseN05
lEQn1S4KNzzjHiZUM9DeZDZUseLCY+qyXif4ceUluopmerFAWfqkIG9AN95V3hwt
GaKAt3ix7O3PWSwHJzSxuJm5zhDhr5O6biUHnviKVRSA0m1jHw+8Gkk00XgamzWZ
Rsx1mwmwIe6dFNV8ELSPKurcV2eEQvsjHnYWG0XiOaq6isV8te47Eul9bk2aLWhX
Pie5bo7lCfoYnYb8hvkVahDLx7YoMayHjWdGkIuBJ0TptswAY6B1M+rsq1k/PaYo
hRCXayBeFE/+GwrpuxfjuhEIj0NP0IsW+jMwDfY/3CQoJGC0z7naTSyRRFw14jsH
J2oEnwql8PC6aT5rD+lK+jV1cUfJI4JCNpzubK2CMmfRCk+NL2KT0ksBGi+wk6Da
YJEwhGfek5vkfWGE93mxD1uOfHY5Vd6GJ5frWv9kPetlJwfftjsYUvU2xETZZVf3
8gv8UUL9vGZuV/7N4nPjTH8zluycbRhA7b91vTwDf0lC7fxHz36aio+4zWNaEjYJ
82Ms2KsfHm8+VQbZF2GD8cnmgXX4LeTcQPRo5WsAF9NgfDiyEbbzF1h5xbSSteIi
Ibw5FsMVzb9qOELQ5rdoBHL8DP0+Fs1dicJuXjbJkinYXXij4PmSmBS57YralG3/
l9678g06KdjtXcdhKIqp77qzmeOAK0KlhCv8M2qMylyfHvKia1my5TXpMZUHBz9a
NJVTGTuLHwJnCfF1EyOw3SDwEAPStD4EIFkWHpodXkkdURe+iqM6IO0W5I+Cuvmg
sez3BuccxcqRWkvgCaj66SAlDJgB6R44U2KtIz8O6nAgdZa7cS/NKbAw8Gkh0d4N
qhuJ4W5t+4kvPfYU2gVuFFS/zSaAW78DaOi3HvaiC+o1lfxXA++YALkSKGoP7smi
8iR6mMsNwqPhLw5GdTd0ZY4/kDcoWbGPTDDjfeB1dPE4ij07nBb8TQlYJN/nPAO5
3pTTKQqEHTzbJYXtUqJ9qnv35biCG55GGaF8BylJGVT777S/6i7joYKnOKv9b8qu
QMycEd6K/QwZu18/7JjjvJpz2qDJ6NvsD8nQJfV8ahtu7sayoTSDpcEFtM8zMRyu
ZHzgahBEo4oEAF39r2lveGcIZ3xK1RtD4i+fl3zNfz/gdyqyaMTdOdCKgEeVuDs4
cABkgGvEUyv5YsR3PYPodo/W5o7w59vdKvA07QmwzDQxS/FsR4FWzB9H/pmpTDDj
IPzid9FlVx5/A7Bhl6HPAPQnVmgu6sMTUGLeoCduN7aYG9c/e6tdu75M4P/uQkSs
24hqf5sXj7/z2Ve31JH258ho6xhz5EoMQxnyKVEXOpSlG+YaFYnDBMaeQcWnDvL7
XVbVZ1VlkZ+3Lx2sUdUQBJh2FGBuEOLBK6Xztbo0L0tI0NVqHZ8HChQBO1CIGYaI
r5kTlhmCrNt8xnKh6gDN72jB5V5vik7T1D8cowU486K5tpnqK9nxiny+QBlagb3r
oC1yIWwG5lPWTnP6iRIY5/SF1s4SlTeas8whymu1XTosDHM1/7b6tQEd8e9Z/nnz
vJgtlZ1Re3kZxyXvL0iqJBXgGWf88Ig2rwKm8fCoDA4i0zjzbcjfF4S2C5jwMW0b
2RgjmM5yzibi52cwK0y8inx82fO317tcL1jNjBJ7Tizu7G1T5Yk+2hrXfDy8zw7W
MUkbyA0VE583dToUE8m73ZzalzaYv0uw5V55Mi0ZsNw1BHlGBNTUSnwhgrAXRktk
8jO6FyHFMYJHVRfCms2UgSIGol2NAiQ31iqF6o0a8pGk5vjTLlyE8Q3zQf9Ab0Qp
Olvt8+DUGXD5kADqTsQBE7ddf244nqaCjvdPAGTQQ7wdAI0RgVBKgi8qW3l/st8I
WIFWl0uqgGSZLvKLULz197GGO46jg05Tko8lAnbkv9eYWMEBErL13TFff/19lvdL
8J2BCoSZrvbN8sSQOqPYX0mI7TE0bRyChsNtzKFvuBtZ2GbZacsUxaC3kHdfV/dE
lbKuCRu41llukycoIuAjHw2HyadGw7b25Ubf2SsQ1RlNUCVK1reuNI/e2kyTmc51
Mzgw+AQBVsdcpY5ZeJ9WBTSOo7QAQRl9+R02KXACbCOinOXNY/59BFa7r51hN1KK
GNaO7YFEkpPwcxDFX8YDmUgGtHi5DCR/3PeRK7KKOjwdHcPt+A5uyJsOuOZUvWQY
3HuVM/MjG7780kIjffL2d/szchxSdmULyWpAW01jsoQmMxoR1odHCIGrj5DlVqYz
CZeKyvd8eSsloMU9R1QvpU74IPp1kDnHbAO2/BPYCLISPk2/rAVKD4/TRw0RDB4r
zib2/2t8hvNDu/+GWWrWLbByJ6CSjDIfisWh/DJT768DJJ82Rd1tPSR4Jy55doNc
mYEhfevL3U2tIWVIdqu46HMXefPRvt/wu+MagAYEKmiQYhmMNOA8v0IxyaXSAHhz
trq8xr3QzX94D+DUhUWHFjl/Wvp0gyULEkeqtao4cvrN/K+S8kPtJHUA/wV7LrMG
Z7p1U98oqzRO8uu/fvEHCcvVsr5eoGsF0JIqVDAENHsLMD8HtE+WE2ZXLIVPPfof
6+muOMRI2RQSV0ssQZJxEZvDOxMwns0F1YaLrXt6Ray2gGyxcW/VQ5uuOL7NU5gA
97k1sv28Rmx8lfeGfSUhpSeTYg3Yu1OSTWeQ4q9nFJI7il3vuZ1Q2L4+um1Y9dAN
Ijvx9ZZOI+tI3mVaKyoYbnqHkKutgxj/Ol5zYJuX+rurYl0FROrvuGD04q2hcxER
wB/5Q4cUlk02Kzu4EQ766RQ4Hztahi6pm7brqQOrvOb7wu4dxemiASED+JUm2Luu
509YV1H7Kg8MyibUQAWR8zCto6QnTP9aBS4YeXT2ZauUtdlcANyIboTDqeQMcte5
E0R9Sr98jresO9j+4wYEU1mwvW0+XjMhoNhkTfOrorq43qAQIsJvsZipvCtFomYC
V8lyu5AzXe4xvyaMhUUkZ8SiTgVVGdUPGkFu83JEbKoB06AXxCYwxaO99mA2pazB
64cwSRFSlXCZnAD/sOmCAaFeiQwhuqvy5ZD56/1aFlH8L8fqr6ywS0SLEVx6UyxN
lRyvNuWhtlBBduK7LiKDQpia8TE49bcYAEzhKAp1pNrDQks3lylpYGI4VAu6MZeQ
yx7ob9GbbvPggIvCfhUhW37x780RhEuIXtbJp24w9gr7keyJFgzabiiNx7kayPVq
Z/gLMfOlgbK5CfJ5t218Cn07vt/JZHMssZbQxRN9G93T6s0S7sM/Du7X+ronIgw8
AOeSQ4tQVz5X5WrfJb/AtJkfPolbICN94RKvjzliBeMKZS/X242NheiiQRe09sh2
h0QRVf/+XECz+cmYJk9BogkAslfw3Ezf4sad3ssvxQHP9iBzJt59KKtLieNj/Mpu
+CdjJejx1oICWGn1bYM7tyKaqRAlrhc6OInSRxhYxWLDybPC+jAoZVN9vDL8Fqrb
a2P4yF4gQH3tvzphNoBmn0JMo50b/juPGUl32Ld/rYyvfFNk1rBfCrKWMxntpd2G
va9EBbCaeuC00wWKIQTOiRowKxSm3dhCgsCVZifBuXVYbzYVdf1qO/KtFIURkaOe
JV+QM3aSoR/U5UtN5I/oai9J+sBDnN5AArJCg7+abzM7JI6107sOEs+qTcRj4PMB
D5SvU8HA7in/m1d1JRSGw6zNmrsndyWcOEnTbm+kSLVevlVBo1B7vSeBfQ/sbuXu
xg9giY66j0v4rP84oKGQKk9cdj78w0gEBVcSDA6OdqrDLaP32LcRTa8Wo8eUnFxP
SLX5ljvsYSIizvSZu2GuTymVaKH/Pn1Dzdc5NdhaUsgkDRoeiPIAV+pUg5z+oF2H
5nGtoPNc4+KoWNkrbD2/mktBCh+3QGXzdyyjAKu9zfwNwVcDa/dBeUqi3x9Iw0Wl
wsqRKxFhypfQNgUktjhx5g+4Gj6g/h7KK58BCviKZgl3kxMw+hfuFKJ4VqmKT/ij
WqFbUy3iFxtrUt9Scd4dUUsLAINjCwUrGnmuVyrFwhVPxYJsGsjy+FzDdY/FIC/j
UHJqNE89XJqGkO2dCZ+C+vHO6Kax0Hw8eR2eDZPQCNoSUU98UGuZmiRO56Pwmun1
KlGlW4UX8TKmCnG/951oL6Tgh2e9LTjDtIdvTSmgfJNPGls2KElx5sHyINK62Qc2
XCxuwGLlrx0wHHqsmFG1iThqI9wirK1PU1REoUiiVlFbepLtlbIwmue32h9hFwHp
L8g9fohoht4z6wmsyyGM5XBUlY0sZtt2bxcd+vrvVGIOtFnm1hq7B6ZTRPjXaZvx
+jn0E+4EHxU38L7PPoe6zoi/gU114MVr8c/TrhXQfRBzkOnPptc/1VGWpqV9Y/ZX
iE5SbI/efwDo83SpO0k3J/HUnDm1y8YGUHVrty1wUJsWo+12mfu1ePaURXyT0o2t
ta62kAEJO/GkhTYZDotBDLocuzUPjeR09Jlqpi2ESyLaBCZ5gNNG2wQGrnfehpZ7
43vBUt472WCEgqINzAWQGviGui5QAtx0XAt0VkYEv3TlXYXLpsbibc6d4CYaMTAA
2MJJySb2XQs7JFXoYGmS84wOp2r5EdVr6MwYQnHDD5/v0J8N2rfRY0sYui1KZnKR
wLJWXyey+3PzWnDAyOE1VdLOI6avqGwkMTMB8AaiMLZDd98O9uNgmi6BwhioFclv
ad/4EGO9/twTaIxT7G4BxHVPbGB8ippO150bFi2eBb+vp1o5eMazWobAfbUG1okU
t3AdgFrTvOjRpAi5tX/CGEIOXOYmX/AaTF9nyL5EuMNSlbPCqK65QUwqcgNmAYE/
vF/BsiclPjlIOXuyJkWKYmBthXvU2DpCU9vqzKOBx4oZsc3jYj+V9TIkOL+/Kd5+
mxRaFeflBga+nlaUtPlQl/+17a/wPrrKLzYhOh+mdHjflwo72l/cM5AqM9b88l9A
GbUI7WBN8bi/jnqZhUn0V6COBonILQ/wGCwLE7+jWTiz++iqx99WWj/JBTZuu/O+
c3q528snh1BliRJJMd+S/rexG08PoY8auIzN4nD3YYtI8GMlzXC+iEOiCcaLXmvq
Tjlvgf8FHLmF3t8GwwGrcn0np9PzPikZI9iDhMSQnaREpBjhXVVnmwWg7PHBmQxl
SE08hj7qWTIxDlOtKBmNFQXl0cTRD4efA6iF/+BSHjEukbTovUUCukRXnwRUSXYv
ynE9ndvcTBrr4/CczV0M9gwtuJ3qUWuzEKhZq6RN/JSmufODTqV9CzeXJXEgD9O3
W+T8wcu9WgCUx+Q5U0ThPoowsOY+/4Gu7FKG8juo90Jcbc2lpIJuIS6chDlcHagF
vBjUEy/j9EAstp6fxaaOUf2aeSDK/K80u2bKAatpk8XfWyx0D8Kmw4nHwdd/azzg
MWqqNsAIZF1YJDJhWcmZYeiJrD7qxAh+/W/jxqzCDDweyiCCcUOpIp6ETI7TgmHT
JLp+1DqaSEgN6Xo05XBrgKxQH/zRjAsollp2JS6jx7DTWsEgb960J4fq9b7acnbx
QSfl1fU3xIXdRYBEGPpjeV9QGPL+y2oYBmgwaEFWcJgTcU4duIvgVuOt4JjSDep6
eZIecMqY7mPnt3ms6hTk4mAnClvncOG/148M3CWZAH7P5j2vHhSoQMBDkpi0hC19
HAf1FjkhnpooOZzF7i16G6/UFIYAqGE4mdJc7hxIaD+iHmp7tGUrTSCbya3y9CQV
OTikEzygzYlrmIsVKS8ztDVxWExHokIIkTi4Jg5sFjL8Ne68CayG5wwMLnUiJgtW
JVP1O5h1kfhzlWorVD0x5oTD+jNJTmckEVjE3BwfsHEutRp3WG7MZ+d2fARpesK0
xBPMAECp9D0SnI/d4Uk+e6RvCi0LO+fQo99BC/RYopo7F+G45P9bubXRDz5Enhcc
73AmngIMPm7R+CxcVNhOLkJZzgl7pGGjbOw8+zGF7nAvDqKXoOYZDMZBlOA6LRMd
mev0S9S1ASWw3omRHx2P3hoEzobwWb3hbAKl8w7aMsXLynwBgMpZfyJbrqrM4Nfq
hO8JyXLKpwO8ilzVlp7gHPMSMrKeDgXWu19hZjKJfIE1etNO7sKaRBoQ1yvHL/TA
2+IxKEyNSl+oPA9r2bBBUVLVOok+FfBKJepeG+aNmWG+ioAiVpe4zODjVpy8UB3g
xY7hVGPdoyFStWmVzvMHVQWEqijcAy8DQ7bwToqYNj9MfPcDu4rQYHakQwcQvAvo
jm1nje4cSwS9ShWPlz7tYRs64sYOzCJR0bwfEB4dKJfQtO9hC7Ov19wXJBjsj3SS
mTPKj+JfECxw5A8AUmRjghGgD0OXIASto+vNzeUHTg7w7IxvTmNnxcttBi09WJU7
MlrnH5cC0icbkLcHZYlD3nflspgoBVDm7QRgMznHN51tIAARXJFfubue2PqOULpH
mEFWRrELw1idUaHBd3R7ZSfQGIT6fBwGKPiCQc/XUioDgwX74QLSw1wEy1/2goS6
+nOG1+HKP4cBz/Q7WMi6p2TAOVeGEY25y6iW1Q6MBazHg+y3uu2nDcBmDHIRX6Jt
f56T5wQIK1cYpioQaeB3x5ovzI/U6CJSY8+xKALsGcsIKlbuS4vAZgdc+rCyxgMz
5cBW5MH3+ZAzFJ0wTJsba6n/cWOC7qu1x13w47vOOt1gRnIDNTnkSefL/AXwSGHU
yHo2f0VT8GBeiim/mVlLYCnLopdTXf9nxYt7mtBhGN7smApAPoJdKw0HQ9xPb+/9
sVUIfEoqy7kHuahJqkUv1n+5eKxVWeh/KYyGac5rL5D/CmhtbxPevlxF7Z1j+9D1
gNy94QPENKigKsmHiflaB9eKAQGU41DAmS5CUsU3KGoai5l+Eux3eQCueTdelAVT
b4G7O0vtwKHF6faAvMKanPPbF82YkXCqYfeJ/HmyEtiFvO5wTQ+a9vijy/AM71Zm
EvC+GzxbVE+cNuECceoeE5wVbdD7Cc9jscM+P2dzMbBA7zfZQdvPC/igNc3qNggZ
if8mZ69fEIkoy+y7S6lOMsWy2iPtpVbwc2lF/k13C5qjPYIFVn5VjfVXD7BtAw/d
wNt8uiXVP9R/+83AV5Ccvzh3avDd4h+D4byUc0uD2blzcS1AVneDGVk6DY9YuCqm
jkBgzPwcz3IVaUDb93rhDQ6oEaaJ4YWuDO3ztF7Pu3MuDARScGHT8VzTu/fnNO+E
mVLCGE528GzrSriZO99m66VPWze6NAYUlURVJWbjSsIMbu2zZZvdbwA5iLKcAYUu
6b9UyBDP8Y7YSqJQYn3EXFJ1netcTUkwkoZ6N5HTaFuEZEqnEk394MHLabIjtn8o
nwu3eyyIyEg6TF9V/iFf6rQZ+DNLTtAoRWIZSXCrIElPsWDVcL1SUVfg1ounfsi4
5gfgrk6YpsjU95512NcC2pIscNqn2z946YKTYd+wixRDHX04E7XEcI2et49R5W29
u/7bLqWEjjJgStGtj14BgW+x8hphc6JmK1r4uwsqJTkdOwe66T3leD4jmp4DiyEX
YzBi88yJG1+8BA3EYdqHFLX9Mz3Nxi+v9aNZf+EnnWuZQ7l7//1CahobqnIqPa3/
FIXOixiLbo6noZz4AMnuJLpU6thkHtAwyzh473B6hsN0a3Ahe9oDoi5zpyAFTthq
Fyy16k9bJewSZxWddQPdOmzfO/Ov304XNTYoNXZzd2RN9mvidKP9Yb8fpgOPg46m
13Dp4O9eMX1Pbk9g8pR48mNW17mbXG2ATwPLueg1qA+OlXvj3jWOOB7NznAjPEf5
r1r2qvWs7gHWTw9L0+bgT3wNv8TSwz1om847c1XynU+anl76AVbT5d1vb0rptHoW
z6dXcPU61g9kX7I+3sieG5MyvEtQxEGYR9ufNlB9lGPO89Cn9lzH9Ac7YUvCQ3y2
k++SkMggUZ/eySyip/ct7d17/nSmKblVlIhoyZVgySvYqhyLcSl7l0J5KWKCUMtI
6O2diaa6s/ZKv4Mc8T+XmlHAQJ5KZ1KI3AgAiTHGHZcgm2e96K/+7H+f+6xyV0Wt
WPlohEzgyeq8oLPwspV3yk3ccJJb7wA/TE0k2AUxj+Miwdx7SRyQcoaQ2GX0Ek/e
DqNlQRsTtR9kFH1SVozfyJA+PVTwgTLU2+Cw2jzDRNXfQzv8ymtA3ZM4cxzDtFDc
wVs66x9YVlGnpRlc5F5P9OS+TLndj9GFCHTNURGAn/fQHan+4GwhTmY+5EQLnxJz
JqTaB9NaFXgGNL6MG5M1imzQAAVQ6J3qebwfvbCnOYif8ZwCx6lPYFxShvBB03Bw
40F94XM54lmmnGmd29OjN6e5RbzLrDYA06F1no3+hz/LtyM27wI07OmCT/qoCmqL
OwACSrrx94U7swFnu+TWmnsRDzE7/SlMYQ1k+1CJgkRRvsch5QtAKQwvTD6V2y51
OAANx1UXxH3f4cNw3C8piapwCl3FeR7igFwxaV2JorB2UON7emGZpFk5o2Su8zws
TsnBgjgF2JZSUYJNcfkQ9Keu21Ts1kBCmsePaiS2nOutQo7nGc3ifeT0wpVwyD93
xVDnwcmiNzK/nk6BlHKFH1tg2IHUfjd8aEZ2ThR1dL1zNzq4hBIdZVI8podfNo3r
p5d/2j8vGbDP/0QiOMzdlIIlexFhb0tzsm03AbBqMcwcrdJtBdRpZ6cEfLU5XZMn
4/TrKs1DY+ioHe/bqBeHgKCKlFuQG0nehe+LXz4KKF99UEfzv/4Bbjnc7R38TcsD
fPMsOdNqcUfWa0nXPkYLJjnSLOmSOXQ0hDWHjOYukYzbELB8ueGtBfSsyLO42SVK
0kYf5gTxozCtK7uqb6ePzWwFrONkrDLSQ42F3T7Tn2kJElZH2XQP6dJ6+6CQEpZv
JtyPR5Fmg7M1wFGgdWRWmQKwujwAcRO4sqNHnY44yja0vQmf/lCwbyEsQWKQ0ezR
MwN2mE25jyXnVWCddU5QU90A58qLtsvl/Iq69FU7nBXSBobQT7bbguMN/wtmBWdL
EtKv+D9A7zu1LgtdPFRHPlNOio0ooLmCkkqeXTuQjf02r+LWtzcNgaWIzCKofO+p
WS3Hqb6PuUHKsrfk07+5gYh8nVXlr8NY+YNs0dFDjcHUjqe44V6sNbh+0C+IJaN4
L7xFZJ+kzm1iArBeu6rqTbliqTN2IZVjI59lfi564+28Xw2VwSHEkUR11vLT0f4b
HJZ3VPQGhTbz71PhyTKhtAGSFsslPn1//pfKiRoHhwQ35x/+7n9KkGXW7gBnOtuY
Vuy0IqqrKqz0h43HT2gld1/EUZ7WI4kTBWkj0QcRFuZ6A+tEkMJS1vNolDRsTQ6s
o7upOPykxF5gvk2tBdkdyp4wx3r1GzUdhUEhTeh97YGsgJThpMJMq1iYCM2DOY89
s70lCc9Nq6epp3Baq0+nylZ1tvt5BRwbK59IQXQDTc0GDC6/e6usQtTJqqUmkyyG
BrvxmhsAqOm1GkFrj3EVRXHSDKVMPDtqDmTPxK3v6z2J3mhP+GtHsv2vqNqbmUnF
oFYRS81kkQmDTXYAXgDAEcviu1TUZRLu7JJoOLLRnclW1q1y9TWcfBF5hGB3AAI9
WYqy89JGsKFRfWcHqqu6/J3cDIcmMeDMUkWYz3vObBNA1K/a5CT07yF06LdZBJeL
wq7HpxOo5vnFdS6V4T1/FLvm9DD6kpv8FgZ+oWgD81IImxA7Z4gfQFtUfdvIaY52
pWg1CDUI8HEwpRer0kxpTgc59UgellR1lmJ6LbRzXKFP7vU+v4gos8Mdbxoj2CX0
eimjU7k0rffzEL2sluzXFBRav2q/RONcglVOW8d7S4UQrclLXxQNVwNo+KWLO5ny
PMxgRbAhTiwgp8P3MC4fi65wu5MxgcAyAFPKLh2wxz1yZII+jhxD/zuqqKi2bLkw
XCEKetqslPvF/8TzaAYinC2iypn/61roQoSLTSDCPeaGuH/bjEeSswuVsxem25R1
TfjQrPpQ2f6GrMA/PFe6HlPNm7XdFhuhm8ShEmDHAqEJPIYycMUnsxX87mjE2dZc
KTTgSnvhl7u2b/TKYwjdqRkJrl5jdGqc2+Uv360HBs/mk8pRbGxK/981c7wWMw97
0vdNVsuKRLSoQgPk1vTbLhlNRD116sAYdLvT1Crx7qwiYfm9vcwDxYtD8ct/BHX3
Mu/MMsP6rCqtAnPqGMv/u11tjEMSa80xT/SowclvoiHaclys86nnBYlmErhj3Mbu
Bj+WHjS/epLQeuWqsfPoShA10irUvW7bvUqLHO8W7qkBYI0A3cpKdyaI6ZW99NA3
0RKfsX75YZUF3GzeeNJTfHHXcBCTIHkg6YowbsqIQ9OmSlB+gHMuhFzyBr244L9X
fzMW3oNsT00e1gaGqtCb2pa/9riOXEyBwP0A4+cN/JodL3Bh474loNiKQNG0TNi6
cQLV6+DaivsTQGCOT0r1saI6UXQws9V1Bdz8pQldRiZl95IZ3UeLUuMoJi6/WV4H
h+fzDlcoCR7nXcxB9RkNDjv4gcbp9pPPGs3so4ouanaPbCkFTDpJlOUIMcdHQHbY
GBhe6AxksB+UwcDjU9yz8D8siHeL0Py4xodfd8qG2XzbUfN9ZvGxdmSjC/nkNryL
+8xCTG3bJQ7ChqJuEqOimd+6f/NziXwMTNuoMDRHVZ9qCa7YXF6anAwm4HPLbTHH
ou9UhQI0uHYoPe6PE5aLIBwDJmUtDlbKplBhoPCFAWUe9YYKR3+53+X7hZhewkbz
2EsQQ7GUshR8ugDofspYw+t4n4sDrUdfx6qNmHRrBvWR5IvmpTVobquZzsjkEs/C
Y69TqVSjn+2uBoPWDmBkWw5GT37LqvZoqc4dBOd5Pz53zx3BLA5XvKL924evoQJ9
2IacPWnf4AJF/xqrp4SKiGw2xteC5KRq2+1Td7HXRXkOC1rYq3GUm1/RptnXW4J2
mbbK5qUQ0sqZCsiLkeYJxEXiZ1HGX4/QjTdZ5qKHx8EwMwNmLN44u4FIhSSvEWd/
A9WM1hlgNEJg/uWI9HqzMFUQM8H4znepO3tzsYHwbPkOkhDaikf36etr53U2dx3q
i0fUEQ3lVwv/ICPtPgAE3mU9FtJjFqLbW+5+CZFFsyRmXTskUhtiYh0vIwOq4Ls6
LwE7MzQRgWmsEEqxjMoR/PZakPhX9GQJV2yijG2URrSmLF4uBXR/OklpryRS6jUp
UM/r9d+Iy9E5jDO/9mJW8bLxjOb4TRqgMnEJQ7LR5dQvZqDe6VKdooyqUHhz75fM
sLyIkaTIcxnX6bkRYUEqJ9MEQ7M6ye37GX8LGL7iD7IEdYSleV5TZMxvkFhnEl7D
suTEDoLoKN3Dyv2Txv0wJi8jR6JtbtVPRBW7AY35QGZLNypS0bPjSOf2boyucOqs
OGxBezVKywcktIGSULebIlpsOmwmP3q5ZqnxQvuRvn/JB0VgHME5cHlhNEg97p0q
uzQvwOyvK5Kww4C/ui++XewUbIraNmWPpy5DEBYhqZoasaIRf9CNwtkIIEogJXfu
6FDx0C0dDTShyoyaRyuUEj2EGYAhiAV+0NeSIV/p98RG68r+rSN+f7MH1+elSHqx
8CZTUp83xCcs6aPRR/aB6SFaV6oOC8qI11+mYup7fSw4VHf1oSsmQp29+90iaqfO
jferG3PQLjXOhXBq85i69vkDmSxvD5JpAKgWdhhR79VLSECuXL8SGwhQrueekXF9
DRa/y9rPKqUsDEIvKS6rdh64dNZ61eEuzVqiIMhzSAxutOp8wlaZ54004jQKVUoR
E9Q78PQRP0tG+SGzmNGAjerXpmHeICFiiN3JL4KpvaM7uy//xxEBOhwd8Dgo4ZLc
3Jom8rg8NaQt8vG3fdlHIPx2OhzKq9A+xUDo9KNgTZcngd8TpQqbeIg3Oi50NnfQ
11T9pKUU+bXGc17V1ZX+lQZTw8RvmSCNNED3oeoA5/BvS7l1yO8vJR+xoiBUh84t
BG0YtjpsKHWIFMc6WadAxr7Gcuj/W2xf+py5C8AaTy9aVosQLWKCrFi321Np2Zod
BHs29IbzjKACNR2s0JVr5Jhq7YKI6yHALjcr25D8dDJnIa8DQ08vids4gahN3rJJ
6txq6NJwiI5g1+za1UtPcBnZ4kZOSI9yp1Ab5fRQmsn9HGgXW5ZepnHQwuV4pHrF
96Ce0dc3h9LKSNSLiRcmgw/YeY0adPvlzLg5a7Ec/jR3kCxSYEJXbU7BKT6gL+w9
iy6a7si7XHjqX9rCz4EWezOtubyelxABukEI9A7MwXpPjVbxraWSSS5XujGs1bDE
J/55AhS8nOVkV8s9KXtK3z7FUdz3yTa3qL5qFsnno2M0x4h4iJ0FurEb8OI7zxOJ
qz+FEpqquKHe33su4Nu+M94KJYGlOyLFsXgpB1HTzW9PgwezvEC0h4X3dQAMQ/81
OpRJAeQHdlMy/xdn//mrJyYCKc1jeFFhkqHOm+nLYm14dWcbeUvzf7Xoe/sFrg+z
L6Kry4fhWJB5QlotdhfwR+94RGjfgoEVep07npMlOyik561kJtZVJWs3HPv18UNS
TaRxu1WIX1WZv0DhA8YrDpDa+u+HCMNb+770MJfFxfLm8vagljlkNz5c/axKKopf
4Q2/RJ1nh2GJoZ8/1QiT+VV5MYdyfIu+Q7DCo8kD5d+vTI5owk7VnpIwQQXVGymt
N+xl3HYDaFruwVdzcRUpsyr+mxkTFSCzc3JqZusfpM5Vbsk8LyiEjBH+3hopxTeq
PiNFTY6TAi5oCwW+3CtWnw9x26XZcsGmedKia0v9lCpiiyfgkd0Ban6WdczYfSrp
lglAg3VTLoqb+gUVCAZumbzUlzvbPqNbO6KgZgrfwP8/JfVvBYDbxWb2sbncCKvO
0W1SpQ1JcoN9KkQlLHKNRMuahOcLXyooqh9fNs8Xd3+4IM1ZS9A0RutzFU+M2G8X
pVwluWhfhtoa3KOMl1IFTsZJFw0f+cBmDZN0L/6pe2YwwaX0Ikp0/GVaiGlXB/F2
wDZeq1dMLln+hZAzc1U0LS723cZpFl4rBUzHLmcxf7UK5//S1BJUTkKgugwPR1Mn
LEeIIvWSBvn+n+c40Ta4a3DFoumT3ZSTtGicJWD2SS1QldxpFshRv/0nP7ApdjWH
ybFW7NZ9xQGOLBnIa2FcnkrfBWQB5RFB7vLvw7jwYGlXf+28bA5D5SSgEWmsz4Ko
/ehzopNzryYFdr8XV7UrE8ChEgLgxa8WBlzfyqX0ykFs7tSbR82/2RktvVff4ws+
sFJjRiqsmLy3nP4cKdJZAiP9EV/mSbY1mIx7TedYrqJGIkdsFewAYbkl/mnQS/Ti
z/96uq2T3I5z7MrmLw8HM40a4A/v6Gcsv6zIseZ4UONAEqnGHcptKABt0fkHCwW3
w4JH0o2lzbkSOUvPcrD5MRsgVx+aEXcwegzxk4TxAwOQhVjsTBRWr01RHXncZfZu
qn9I609OlmWyGWq7sD21kpXaOQLm2k9Km5I1dzC5wDyxk8paGuelxvmjHY7RPZsL
iBr+zlM+cblCRbuhhfhEGBXk58JHsazB4yIO385QhC8tTtTv/Vb+8zjllUl6eVa8
xjtCb29lhWATCDTZtDQiPZbcR3VLZJzwUgIXe/IQn1m3w/sETa67j2RuzyL7dgxq
jL+qEHTedx871xvNEsMmMqiexxSjnvcx25j3/syQRdbdV0YgehUVzNhBfqQEc4K7
7pTFuAerAYdAeCCupgxdi7Uh0o/7w3CXqFrd8g8VkAzD2KDlYpjGz4fE1owRJaNg
7wH7myXPkciVoHm6MaBJlN+7igasG7vmy/2vKhbokLvHYPe73+XIuFavJiUca4Fo
kUJpgltpdgDCYiEji4a4uyiEjoGzkLBLHqL04bfWi/7KMB0nBkkTOhu45Sv+UkTv
cwQK1lRSbac+zh0+JLXaARbO+Qd/gVynQt5hbp/qRlDLeFGVRu+S7LEe/4lCAS3O
99Jqsvh28wo+q005EC4Hex2baeoEYc6UeHor772L+qDygNW9eugMPDX8g2sM4Hbi
6EepLsT5+5ALchjMHi6nwmjWTXOovtTEx+zCywNpNwx+7sGZru/wI6d0IhlF4B3q
98zaXyA00Fq2dhvXcO5KM+xLgtgQgB94aPYb+GgF+NFocivTGjNvDgmH/P7dXqbR
hHWiZJZwTM1XjAeWgZDAOADOhW7WoukR781S01MkS3hTT7LO1TpMRNkVNsO/PoKu
UE+zgROnm6Qj0emD7qlkrK/3uWNmCk2YUpMClJYHsV7QUyQQpfD1I6TxP1Ooo7Uk
dATvf6hmL2VBoTiDYVQ1a5YQIkciV/MKq6PfF/TsxYCG8ykwgkb8Q0XLygAW6UdS
qKg7I+b/WDbl8lnn3mGmw/JFn3Hk7QYegI/eMOvCW+pTOqux5r4lsXqKrmIrjGLl
G5ADYbKfahMLFpx/64hki6npUEEYTdkq2wwhYq4vE5rrrHVRMEJWtUlzTXyc3OyZ
POI5iV9HgzN9go281aQe0/bSuVr8twlbZP6yf4Ahbgp5FtdoG7wMmfUnXtwRr0LP
6Cy6z7j1t2PAolb9oeqFCZW46jcwDT3yPl1fNHiKL8koJVzO3N93390piVGAAPPJ
aysitV3WYCCgcn29Z4XzIUpacfn9Qu/kXu+wXci/vlScV+zt/pSQpDvVTO9WGqbe
GOPC/Wlw1RXhkKS+dJRI3aJOJiLbzJ12ZiRPA75lifri/VMXU6XYzoTctbLSHXhc
57bnaMdOpIDgWX20yId+YaAesqDCp98MSR5lpC5fQHuBVUH2DZYxTw8eG7vrvDgV
lykRnrKCK4nhwTQJXyIenZymjqghbqKlAv6kTxgbS1d317v1E0xRD8lVacwQ9LY6
IoQDrQw57qgYBFI1J04EomP5hz8a9CC8pavCUAib2Yn/0BQBhyBJTVz12NSeVfkV
HnEpLIu2wGZ9ClaVb4a6USRERtQNGPSQBEMX3dFIOnyvLWPEm7GHgpHoFilpfbvy
WkV96H0DASQB4GxFQsW3Gy3xaew+/bCHzep+3G0PnPEjLDzQt6fZdCjUAe1B1NrC
pncMsw3qeeHKP1AtOXhlMWMUIQ/9QAJ/PuHdHZALutx6Nh5m+mwyJu8lKpgxYzYm
QNDuaBZFlyo/Ox6DRfZC3CiOtRkze3iUUSXTLaFEhmnZZmM+naDhg9hJi3qgB1ne
E/3+eqj1ObYQVdI8MU/mIv8CIF+8ZobGXJOSo6U7va5Y57kjedWjiubmx4yiGhFG
qaGmYQ6oCHs2YVsAzDWqeDgdSFbpI+uhQi15XzOZXCOi8fKH3xPhFg2xzgvgTH4b
SQkWIG/s0b7qTI4Ay6HOGr5ko2vbK3CvMt0/GVXfG9QXoll/pc5z/BTyt5QYJxOW
C7L8JJSQzoxNZ4L1WGhYLSEwaVvycw5Nzcx4N2ZEio8fpVjFoldSiYCdVCXSKG4k
LPIbMgrUvON4NhrPEODprE0EKerigLyRWYZjMc98RIInzqrhwbm0O/1ksLmqmCzE
/MaLMiqcLServKpIAhZ3rKpmX42O4J0uxOgBzHMs1rFUDYwIEFZQOFD8+9Kl8ebZ
46DmvUtfvcf/EwK4GR2BNHk7PgRbIiaVAQfq30RKV3FR7+d24BQLVYxq/0ywYJ3Q
H28yjAn31MzwdQwobIbpOBvb9EX3R8/Zbb6FhKzcpyLOas/agWGtfkmke0jOgQ1O
ELTueIljeUy1mOjjw1x8OU8EI6RYbKm4RS08k9RCeujIojatnLz+dRUp/sxDyEb7
++RANbRbyJeR1lCtnPX8uASV16XnI+DMxKfsYHhGNoLIlWxqgB6zVzfv2WAux7jM
6qg8sXcG50E/w/Fg8kNvxLxbEzt2YtSaB/HUROvcLS76jxTX0IYkBocDn8grvTYo
LmusL3+agO7WMqJGARNRwaQuFdQqndydCDppkfKWHcB4puqsLae+kW+qhfKw2Bli
FKALLBbkIwCWz+VHOYvA9TnGMyrgpM2J/hP+4AH5ybEtjCf3NcVyOH1u9+OiijlM
78pEygeKRG8ZjPiLO9+nXH19GfOSaiy2UbkzvsOiJ/v4ZA1MTFLbzkt4Tf3Uj5lY
1EKi14cvEyxkPX7mnnqN7L1g6qMYN2FRRHBOu64YONoPIVCL8ldaiLLMy/U5Aooo
8fW6HUt5Oqllodmofxz46boGwTwOvkeg5/Zi59vJKQovIP0Zmucr//QjhC7e1KEI
sIooWRCYIg9umiJXPcSVpH+nLhJc65lv/ajcJpOG9scRl5zHY74ikd8mGOy2RmM7
mrlPnCFF1iTw/PvPxnnQVz0FsERSCyoOT8nxXobFUymuxEOS3FfhIFf/dEgsKE+3
8NrtSfzgEr+WalSXYgVptdkztXJJ4udRkQ07Z2RUr3ysqJrjU/sgQrb/rrxo4gTW
RiEqvzix0Y/rOzlxgO/aTwyvZ7zKEiaq+H15STiKX/rqlDYE0mWn5sB+wIy9pZ9m
4PXUvUzb1WfJGFPDP+AupzhJU+crSpsdpByddZavpNESg3//BGw+2JReMiKaiCUh
MSuZZyz3NI0P8QhiAsrowfC1j1X8FTCl9tymkHTGwakwQT3/2vRGNY19C34uviqS
2B8LJ9kva1sh8nLTWsyQ2qM3L7sxDaVATQt+zagq/OzzU5wlr8otPw4LxULLPuqb
mmI1uaoqVjYGMi5ysPBl5ewMGwPfNj5RkxMkulDacsE0lPOaNx6uQMgq9q/2sfbZ
/7h9zH7l1btu42cF/4KDmK6+kawyuVKqABvDGKbwSnJ/anCR20S4wvD42RGA8ZxL
/jZUeuk2qTDj0Oi61S4p/MQuJp8I4OFgvXdyUOnMQUJK1UzgGdAg5pbVLWcG3E8t
+tiD+SEBq5nf9sVbZB01L3a+ni1swTZfbMJ9FEXe6yeMYvr7bkB2GG2Fxt0K6lkz
frZjZNcuKTWQM+FrwdyQdtqUBgqpP5ZyYJcdx480MfCGg5U2jpF5K1Pp12yHeS7+
+kn6XUkI2K78E7k1LsX0j+Yt1MxGn09mHmGk+m41sHKtjmLOrgoIDu/CAoq5TuxV
2r4KwssIiHmwxB1chTvkv4pG4cqX4sAgiASp9Y1NRirf9fHoppdbJTvl8Ok7ihmc
NJQmLSJ8amoRrtfxarYMMVlILBAAwOgUzzRCaFY5KAaW+q7hLfuddeG32bzy75cz
GK4kKBWJT/0kr+fyPiihc3K6mYyJsZAZQxviMTcZLz2qcbe5FVnZLti0Wki02Tc8
djEgSyQTNqomliDJorN1r7Ty05LSaDnY+U6z5TpuXUk+a0YX8BSKwcz7R8nUt1TB
NCuuPBqj0P7gvkIqwExHor07w54+WonoHfgzvGfzrBtD+42M18DAKyaoasc1PuoL
cLe6LoQtEMhsTaTg7rZRUn7CkbMehMSJybUsPRSyXmFlmu1/vy6h8iD0yoXi1Cs3
+QhOM6GosunvBs4T2OZ0ZNPuyTUjBf8qH2uJqWzoxOIvfonPwdsxQ1KXkBlHEXuB
BkxCTtcCYDgFT48EXwKiwVKsuxXYKGe0xAjj3XOlbPTeT5h0JLD29JfScWNZ3S06
BgFTlt1dE0NIrcxpCR5wvdvtftS7/2v8Dhp5CAZ8SgSpFuoqu436LpRAXHNmddFu
d6oIqGaSXKplbRp42z4eUY15EUmSpzRuIPzGq/Il8A/dzoe6UR+esz5uv9FA7L+p
YZt1sy+939nxwy4hUEd5HhtYvg9F7hJpoE/ugjRUMY6neDBU5EpXMZCatZYblbVs
DeDit0WSDZ+KP1nbaZtNvQ0Jq2MxPFxqkjSfYUtsthhiOfMzArfClV3Jzov+4IqQ
/AcT0Gn63Eh+XtNr/FscVWYfn2k93f5iYUxlExXw1SPLk1jGvutHE8VcOfekj8W0
NQVy4FR2BZ6/ZXFxe1DIN/pVVDVZTEkgMTBQA7NL5561ZR2m1gcuTSYyBvjdNbtz
GNoY3HZbh85KqxQq+MGGZXvOzsL6Mh4+IhUXRMgfHQ7aZA82I9M/8udNoDg+FLzG
liBk+jzpLvi3HPdgZlHOPQQL8bNRVIzV1Y3FAB3HpZB5l08tsLUMIh+Co1tWs+3g
Qtzfy/L7lpbI55b9zunisqNWFX3AIbSQCyxAq42q4CVAeQEQPTn+Gs0044RWjuC8
/QhAGB3vnmpHGXVw5zllVcfQMkmQYjbhZyzPOc52AzLt75cHydpo5bSn/CSZIWbW
96ZZU21vwSltnAndv4OV5pzJkdX76VwHaUInXhV6u1vxGcTMvSHo8D8BNyuAC9q/
bQvQk9IqOfIe5ZaWbqbyoZs5qIDCsxKME15/35dEBu+oxT0qM9hlPnTgKYgNwWcI
Upwj+o0VPhRerNpsqWUpzKlu5QTKz1YwuxmXnII1u9gAZ/+Bx0imbsGEzZab40T5
ZXUv6a5KDDRwGxCDBj0l5zb3IY7yHmCss76+kMnVc3viTklrvRyZig46H80/kkMC
RB7hKcgjGGvGAws3ZYzrivgON/pDcJBiMw30rWhMdT5rCtm+vNuQQYpGnE0wnhdE
By++bNBgNv1pNiiG1PadpjnGex0JSDToWztoxEJzwTl3GE4wlEk/t4bmCOOIFMIW
FRK2WVntU4Z2uC8P7gNkwYTLfuYk6qcg5UxGH5u/nI+o3fYIWiAVV6wVIt422GLU
usy3/4mza+k/FISg0IfHVLyE7m+xxf98iy+4gRbcE3i445e01r0pWeS+elRxkXjq
eE7DNxWH8K2VbBiSjmJR8BE1k4s7phJ+hWSOfdshP1v8P6FXRp8ZTxACu8A6kUC9
qehtCEwg5FEdJ0MKMTd6v7XvNHt4ZHA+O+IbsCTcwDS9aNl+5sZbSbWCQGWx3X9H
u0Z2vUdZMQliesi2VYVT/ZyQvmUcDHyRAhG4I5BIISYoNwpjPs53T3n7ZbkEFJHi
phEWxu39Pn2kLuXryp0x2f9hGf2SfBaCP0vXoiD3Ngn6WpuUd5GnI3ou7n19Rk9S
H2aE+JvAg7XqN8tBqyJQVBw329SdwndmVRROLEobmg2Z0A+6H46rqpv+Kl4FvfUn
f5pr+MH/o7efFI+2MBvf9/7/QuCXUyF8G9a2F/1bojMOsrehoFSejqygyQiR6K3a
tqBNSdeycOoucarOFzQVtH+vywjjlG1/grbz7Wm6nIEVTD4oLb9g/2/wk/2DzHJf
jGB8MyImO3q2iQ+nj6D4fTsLJdONbXKFU6AlXUJ1+/EndPI1nAXrAygnZ8JJfgGm
OKFFeEvWgunoUYdGE+IMl6Dp3aeD/NluvBLkkh8+T9t4k7L7vKvccUMT2xKiUQHQ
jYylllcJnt53doYD16C+oHid7BgvBkurdCWTRvtsmli/D+QayEUv+5eifQP8ix/N
wH5DQGybNHI2A70RQTauyFXGCUMhnRNwP6qQlHoDTz6xxQltzJ4pFq/AchxveOjK
cSLpReNZ7YQ8rS0+aBClg2Jgeqs/N7g2/fk+MG2j/NEolKnYh7uPmmWACH3CgUwL
ys43Q4zhG1p6YgYs5AwxGDTb7eexDUNqafSitRdGBIQOzUwwYnL/ruHeJOEj/xQV
Q9o0SkP0wdguqDW6xNfXyQYAjymxbnzC+cufg7vp9wTVAJBpFaDzdIZK3jaiBfaH
XGN5RXFbrw6+JJKoW8YdP+hrUDG4QLQaYOglHvO2Em6OMw+1/rddXBe5EhyZFr1C
ef/chQEFRPqOZVSoRtjV4siTquiTny1cmnD/2UjVOcdAldHKn5v5HVj3EddXW83V
xFI0aYmlMmxDGT42RsMMHSfX0kmZAGxxujfkrfX+JCtXn+AvY3moKKImM8S6J3mL
yH2RxRsqD1wlXKMGmXMWH5bT7n36bACzEzQROgPJa2YAZ52j9664P9lpM1TlcClI
bC+Yu4SKoO5CcN9Hxexl/BHwzM0EMrqxcW1TZinU+PC9cEaGujwExovSd0CVzZm/
dzuhqpVj/PwfrSS329l5JmYN57bkA8rKKsGYSZ03ysoCuIXn+Kx8LryWICNJz8xJ
U74GtJUL635/AITotevtTE9ZIzhG9BHt2EL0gUpBJUtVAGSEzp0jDxhcayxZtFdf
XtFsIN6a8NqCi64sEzma9Rs2aX5bJ6R/OQ439ZskG1T8QizOm/RjxWek2urypXJ7
C0gz4U6rxJ2Tm1AU9dxvwD42yceoOEuGEsBJxS/1Z16IX2RLGKnaJubgSZE/xQLP
EdjTQQOtSTEXg52mTmNMSWSiOOxYENsSYFT83hbiWRdsMhRcnnJdetFvhxtMMOgb
hzkmroTgA5vhvBTSZSQiowXacH7S+2WrJwEz7Ifp6qC6qPQTpkWMLONxH6hhGcNP
slT0PMLeP+nHxn8qAXfCWMdkxTqG3OY9L3WvBStrsoX6ISXwRXNMMNqkm/ozXRTZ
VmrL8vgvAK5Tu2WsYtzCKmG0XQx4McvSENY2vQDGJJN7aTxMQXy4JejIWlr9qDbe
as19RakIy4bAFOyG3ns9mCoBDTzxbj2UjOBSExZndwYj7MNJQARbXykfjt0cXsDI
i/Ea01jJyQ5odERhXLBYIeeotz0oJTOmw3y3VAi21gEC+Au+bjHrSfiCpOVbB0sr
L9GFzaQ+oUpsA20d5fFxXMEO04PtZWMcQaeJuKuevkv0wWDTpdBxOnr5hjXl5VYp
Jsud4RFQEc/f/uFmS+P/qdUe2Ea4LWYzjfjmrZAeTX/2AQB2j5z3kFEZOIxz2rTa
eJ8bpeGNy5K09g0m8zjFCfyCpdsPoxgQC0nuE8VcVHdUjBEBySRWYomFR32Xayiu
wplVe4DKhMwfY3oS3ntV4MvRotCGrSxegEBteP4ZLSZLdR4mITCpPauyDpNt42Tq
e0eLUIbtAVWuU9ng8fj8dM/waesexKmJBs/DuamINND4jolJKVydsFlHyt0DDTGd
f39kEAgYbnLcmHmuGyG0Z+GsVkaqDZu3qn+VWT0EBF361KzBrM6IxlS/BxohzUJ0
ZnSBlAdf8cMCGv0TAZFVu7yGNG8VYsvMiNN0PT9DJPrk1L3GFip7QNTPa/hps0xV
Fp8dWRKiZ58oZKcGxWpPtya+4X51jn37O9DHeTUug3CahjQL5XgkGuii1F9vbxI0
adA0kUqda9ZhVRirUS9EOSopKPxU7TC83TP/dkxl9VUCycuSYid7lCU2gdWYUVAq
hb87llxr/8nkmDylVEfkJ5bM6eiN4qepsLvfYU90jNOoxznde/DX8WGTKQnPxThR
VcV8C0D2dWoCcDMT3Btt/AT18yAnw+3+wAnwyFVP65+nf62BWq6+/RDyDtQ83MIC
9UAAkdBohQdK0mBi+Fk7hwqvnjB/wh0cHW+MbIUv4dA46xjz2bMLqT9F8uW9UjfI
1sKmJm7K4+6Cyqgr78TNaiqpbych9h//k1j7upqmw8H+4/sXzzVsOpVUCUsuNsI9
tnFLMfUfJL+lCwfU5163msYOBeY485oMXiVtvtk07bRqv3cZaY69Co5gsai7qsLl
gQfSFw0UH158W+EvQiShhy8IitmG2Vy8OZW/v4cb+NawCohWJ3dVW7DLowYvmhsN
oi1H97/Bz9rSSm99tXVGFg/jljtEc3BidSSrKAOoxngvZRhEY+5pnR3+jxUdhag1
3vRhfAH1vl7YFNLvX67zT33wd5bZHwQ0k26Zm1wWlKponL1Pn9CJSHCV4/qlFUCA
iSdlJPEwtFEOeNZT9qpaKQx9d445abUyhhNIift1fbLr+beYuepRsvDEy3eLEedk
+Y1bh1yLkALzwVtMw6fjKiDVtAny0ITqWLvdxFZUQ6xSZcKMxFmqZ0I1u3H3B2km
N0UwyL44C22tEzA0dIXUTL4o7zDM8MSv+5aGyjRXVUwh9h/cmmwIlUg07brfZAFP
z98r6rCsXssoa8FVdMN5pcyPR/sukLol+q3p/yUm6SLzmyl1nftogy9slJG907Cp
OsQyLcMetrZ5whmxXrPjfjgyZWQRW2/ZXeEbTW+ieP+fr8JSj3s41DRshSgl0qiK
+xCW5klcVf++1kDmnhYhHinxO2QbgiFiS35moLRXhoaMUIg8hI9hLPgKKKlaHEWv
Mzut2AQ1NZT/Cqlx1hZq/EVlggyfBkp8VwT6RsoM/vXKue7UGtrZa0mh9PfkWZvp
LoCYq5zLdQjnKZ3MzAoyBxA2ZSdhXjHHlZ51PMpjsayWywnJ156vj4l23GdO4w0K
bV/I2WgSToZrOk8R6Gdu7+/LqxaxEk2B2YO988H7Q3guos8tUaw7gezR940CXhh8
X2E/pfn91Ny4fybWBuCBvIjPfCbgP6GhK1zKIoSDt90hSuabGMCTwlCndO2cPWwL
8hPniFaQFciKiZ5nlIgKZdGfmUGaAWJ5EF+K8wjD1+/kakan8T/rtphSx4TE3APx
f4F7Q9YnM0pRWYh4ZJRZMVIbSL+eh9Ll8+hThNbTM/HncysY2b/OswEpMwYD5Pzo
6pVNYO+YoIHc01iecm84z5isqtzU5gy5ceZs4JC/N21tgPvwce9n/1xmgPABbnNu
C+9CSqzfoMNJabEIz6V9U0CN3C9+ULHoX2qejGgPC62mulRKg7v61qUWcO9JMbQb
rHs1gnsDQpKeUuNfYu5weRrBzL1sr/vkdcqmW3fL+YnBTSFgizJk18Y3yClFxzGs
5chUaiPbJyhcmHp3sRrGAxWtxW1A9sdrQytVDnEQQE5zuYRDE8xyD+9VZo/8dsbB
cYwxPqX97FTOkG4SpuDfST5oK2EB8zW4K0OfKdtO9CeTT3tIoHa0Zu0vD771EKP4
lbDAvYEwZn3K6f9mkbekGxwgbwmBVEUXKqPTSEU0nE2WkZ0f7ZFZFknB9N+Np8vv
ypKpbk0bFkz2342vqc64gusLhy9gfqSCNLoQ0zzjkhYi7ecny5vaqToI45GwGcMT
nbu0UlV6XzK71XLA4HesnNBu1pViqinf3HdyyLBtlGJeaPzxYwSjEIIzw6R36GmE
2HzPykB8QT+8DhixuZvXJXVtRcI1pi/1lPkpzuzPCVFki+bcwbyxF5DT8ldAzJ8w
DVztzXpAzstLQFQn7KxNkekyL3NWDdBMfEiPfzfASeJs44LOdvY1+muE9RicksNZ
A3la5SetK0oMenM/5vX4KFefpTnuRLZeSQHiWMR/kB2NCFVDa/vzdRSlBlNQqAbm
r4KgI70zXNQovPTQfGNFl5p+v53SjL+/sv44pSfP+9xaFt66OBPl91y5WIP/yJ2j
kYGxmaHKksHLqJ+M3vWC1+Y1h2XzEfBhwdjkbnfUWWE76wPHtmJQN9UxH+DN6a5K
MM9tYTkIubea9PCCuFUWmMMpxeGAIA1LX/WLLC6A6X+RmZy7OnDksXv1+sB7XBEn
gRZa/7GLmieNSJbqrg8qFMwQYKTxpxI63ia7AdeNVQOHiFzTpFNtRwBO619ZfWRO
Twk3EeMNFnVBaCqGIiH/EWfslt+IbPfFUSlb0aIxJp+KTCK5I6Jo8xwCV5r5W48M
uhq/VSE0PdlHAcRljOMHlrqHLNjtL5JwFAe3xADHOCL1TiPWin2kMVdzOCZdaUWu
9xlfNNZTj6y2qe8i39xY/DORsohMB+QLy+2tN+Ovn67dJ/0JlIxzcvdcpBtQRLmH
flpoehFomPooRynZfGCzxcQCZLXX1tuZtlKf5UVLsux0OVuuWfoN36FzpIDkF26W
IU8bsZNxeYMlGiNKxAFTL6Bnoh/uK7GFW95mw3zk1XmtUrag4cfcBkV6GB2gNFuo
f+ecDXCb1qgOnDvOzksjz03WWE8zSNkxtEHZSZDoesX4oMnN0Y5ndxvDmb/0bo1F
c+YT/AzdgZMr9OhT9TyXSeHf+SxgAwV0vAxDm1iYsecAzSnlXDrFQjaQoybk/SeG
HE7+LBQU2kouorP5/yySdWnb+73hED1PvGFJMzYVTWRvf5YQlupPkCnESlFmc68G
Vcjjfvkb6bpYg6b5lMJvK3SjWntbZSqgGePQQsDJ5f4xePKDEi8rbAYOwN3rE8ga
/1lbyisG8DRAGjYzWOcLUmULdoIPR04+LFf0hZlP/H94O8cOkrL6LbpmWXjJepYd
hPsoeqsQNOHaWu3LSdKhfkRJIJjRS7e/Lmyyt/mqyS+Dg5KYuLk05zT8r/t5KYaT
Z6x0nEp/w9thyxEp6SF3GiAmN9yBpdTMsIkQIzSusYPAPyKJeskEUcMLkl9yVhBX
cFJBc5ob2PEGgowynzmCAl3bqM+x6ac8jLnB7KHzGzS0g31v29HnHSnK6Txs6qFb
eHEyoORVGH6CWFx8BzIRmaIESFleKd3Bz+34UFJC/b5vKjMCx9zZ45ZiS8NUydLP
w+mjWhrY9bVwcC89I0ufF4P2DOZWOumMA8s/3JMt+8//TocIpYfQMZRM+bmkBfDs
Lz+Iv4kzhPXYkRPIg11493N6LBi8ds2OPv3AV2cTq/7/K++/EFqMdDwImdRDWlYI
69oYV0r8VDmAamrKblrPH4S+DOGWJrx4uRFVDa3LHuUOZ1sgGBT/xPjzrHYPx4W2
oHbypiscLQgTnK1EW4DaruPedjnAn7b6PWWIQguL3k4hmEjOCE2JLpWFobjYW5Ok
W67GflubpvNs/niYIugKSpRvu3Dw6Hkm9DWCJH6jDR0kDrF7gx3BFaG4DJBxE1rA
WrnkEBJb+ThtnW84Czq5mZbOJZFwKr7I6Y68i+t1okws3QpXV9mjw2NNBnMlzm2B
DEoctRv+J8bg/Vf7gCxt6z382ziKoXJaX4fb9THrBbr0bEV4hjrHIgijliEhFJsq
UV3obp8yonLwwvEZyZvkPq4xyNqTjrzSHloMSPYlkqeD8LBCw6gLAlE26Ai9DIoK
AsNRFipq2bHBKpYQ/rwlHEb0aFInmcTOnrlCwXHufn18zuK0vD/PELK33QnmF5vy
bc06R3z8LMtRSWc/YeT5x1+Od50Ak0spoCbz6XfD7EdJrqSafM12rqQWY15UKY2a
Bl88FZx8UwnkvV4fGlIvDwMJABHCNaxyqBCayEaFSb89idHvNQ81SzFs17t1Kiaq
Q279R+Rr+bngRWeuvuAkZOnapR7LA6frhrq9IrG6EE69m0hghqYJ0ELC3wCrD6Hp
KGn+v7PATMdaXptrtMlx08ou8Cc6HbR1jqDh5rvcw6xHvOUr0aGZErvjkxVqdBS1
5xa8MYshPGrqufBfO3HaFq7OyIzv8rWnZ+iVpjH7LDk0V07I2UgaaHxGE7UUimpm
j7osav7Znfbf5Lo3Bq7di3nJrmJYdttRizOLcjRnM0T2HKk9J2Hrlnh56YNNoKHV
xdUNKhHogfSAI5RGKtqp3YRDUz+zB6gfAWhxWGy68XThlfsk7wBcxhze+by8Qztm
6fg47W6eeKOvTjwz3rAmvcuQOOWA/0HEZqZcLMh9TDLGEHtl+ZuRxcPhlhvXcRyG
oPBEKvEOt+byvdaSSnfd2NlrRLTeXIFYo+G7OsnJ7JPbACk/z8zVM0Je6XIxc/Q3
Tso/IIuOjt5SBDaqYMqDVzYV276ClerO4qPW+yCUyZLMPIw7dzvTGw49ShHMpnJ2
L/j8mkrC0uHUQ43OtejW4DCN18ZjesrM3TEPo8aQN8OTbAOCt/phKdMGX3d5dy08
kk/T+XB6HlIUzjGpDxFnmnFmeYHpZbZ4nrfAiv5cew58MKYQlsXU93Jz5IEgWmmG
Zxuz2uTGjS/hp6xRgx1T2EOYKaAKmC77tfgnjfiGZWckFO6i9uQ2UTkiS0UzmavR
ovW/64L0Lc32vIdutGSBEm5o3+riGpifvbCpnPg2CzRMzwlRc7CV8rlAc5D7tY8o
cSkK8IkQt1RFNHiZ7uNss3tjbtnJ4+7OVGK6ERig1GzJ/lOyC1KGSk3X47TeXVt4
eHiG+stKYOb1MZbMuJ8VWYRwXDhYH4rIcgxWi3qTAMEl1dBHpXckyaKPx38FUDd0
rqkTlAxhuCuZfNj2hafHbt9gJMu8vV8RfeSpWGczeWVA/lU+5LmuRsr5aSRbQbPY
ezk5ry6PAdGiZGcmh0aF9ojDL8w+H9oVwf+SEEHDr1W3Lb4t1/dTsregkWoAAsS6
Zq4aI1TGLegBmF3PwaR89vi2tnKOdmsDKS1GEWWNP23XfEmklB27WZ5awTGAUJ/m
aHNNw0WiAFLZcTRN4oQLCXFpm7qZmake+pjMFRq92ZTts2VSa1PAO7LxW89t4EO0
szVuJh8NTSUnhT/bHDtpI4J+84macTBRbICBSE/WmCl/pWDgb7kDxfupyBrOJFR0
YdjptpSzNZXvLOep53Q6FM/J2o60SqV6QV98l26B9o4lMmuAWl746qpCTnIK6ur7
7o3VpxeV7ZrLJC8h6XSm0Mv8MU4lUbYgcFw0QG88oZvZBIP77P1whq+z6bWY4EMI
iGRxC51wuDauBPZaoHmBi94Mbz3zVNSX4N3xj8RaTgtJuc4NKC+sm/M/PDbQKWXQ
sldYHJ/yrGUkaDx87GBPXjMe7oKQzZX4aoOq7Cf5Y2Z4o3W+CkOdQdtvhEEHtWu/
uZUrHNPqlQdZTI81UC99Um2Iof1C0n+cUVDNrB9QHwiPG7XqWe8piRpnc8MCrlfI
mgisLqz0EHKunf4X4wV95DAGetPtLMvBsta/VrFnU4wYC2ZoyA1scg4YjqU+TLs0
fmZAKbcLiJStaiKmcWpmL35c2+1amopyrPPcXYOYHvcUxi4wJNOxIsEZM9HeZFRW
xXzXqpoCDTnoxb4LkUNT6x5QGh+yrxj6JkFqCdkGGlqkRtK3IrdxE4yHtx8DRiMm
Dp0GPbFAuRSMmEUWmLseP+PeFBQkRWMbufkcD80Y0ooF6QRM9cs80/1AkWyKqAJL
NNJ6L0CTTMiLaT/UNqJ0/A20UAEhMFoi8rF+xwM5lwD39DYFIzm4xeB4f4NvKWR4
1mogz6Fts7vrdYMsuah1I975fXxUfM070H0DwaRski5o2HirVZsWAFR294XTd57a
g2o2rpBua4x91BA7iHOZGOzFUjRCOqcvlcll9w3GIPfIzUkPwq4b0epGSFBXAkdb
EuSHcVmhveUU+flBQx0Znfn87VA6osNDg5HgwOfnLAChfbQq8XUsaUtEJsjKulR8
KXU24IIAvMzwYA/RJU0lgOukDSU+FXoNzAuNObixENdKCCBBW2os0R/sojXdMNNS
W4ucyuEO5BUOa8rmS3jxKpIFPEpLNCN8tDk2RL50enRgeyGM+SWWe9YQYSo9l8Mu
rZ7no5I/+oQ34CZ7gN8cLhRWpv9z3q6FyTFy5LCnxZI3bh5QgjCrTWGv2qyIUdR0
WbeBFGPY5gnti5N61fQ4EIJ5D5filpSDKAqyGSGAumdGWDU8fkybucbWFXdS/njG
XriIx4F0bXU3NQ870NlXncaS/okWrg7Nsh+dDpiCosCGZ456/wtc6hZ9L9MTo7Ua
fBdYotke/OXgWyxjve4L9moD902RwNbo/J0L2irA1H/BYE283Vp0/N+A7dFpWyXR
KK7RpOXgi8o5eUGhLyihGFz88CHvE7M8V83GZJvfiWr6XcDPhzf+gCixeX89dZPI
TRjddvgUFg2L5e+/Z3ci9kcb+hD+DGax9VuGUfAQF2fg0jmcBZ6qp7BrK8sJO2F8
2TQSKbpfjpLmXEW+61G2nzBC4LEPUUvDa+5zZ7BbpcrZUxMVh4bV2n+ceKKkibhL
I10DgXbqk9xAoSs60Felm4j0J9a1voApi7fNg54l8JTgwgOC8S+JOpL4OqT7p14M
wWJ+oliMxRDlbwKL5yqmjEYLbTCOuCjccVUQozHwljlSZpVlluhzXzl7h+UhVVBj
tKYx+VU8ZiSdMneTsQJBI9KGE2Is0zU7CXtHuHR/Xtiu2V+5f7lnaKoSLazkNX9C
jiQNU6iLok3g67N3qB41mGhuF0AIpk0o0v5WS1+M22Xz9MJtgsEfCNMeUHS6nZcN
1rMJvjmrnEwyV6Y0YCcenmNQMDaza7mpltEstDY+TUQ7puRAmtxu3o/BtG6/5LUk
OOLTp4TOpjHXBfHeVnPDugzl3NYBkMZmtkkVSbpvWl+v1pjk6+n2idjJszPE+4x0
QL2wSxB2zR+2iMSK4GTgp5yPvyRot2jchlW3B/GiDV4pQXRtG7WjTJBm+HFxCYva
fWHS0M8Vo9LeALPyk/xTF/cKcELJ1FG4ukmSnIROjFtbL4Dqm9i7Z4uZzjTHQ7VY
+W+0YAo1wGSFMQdW3UZs+d9mTUF4Sgt53c28kqVeIyNS+7XSE6tejI7TvOnjRpNT
FEYKWtxWgmKP9KlH2OVkTpiHIJR2+L1wA7ScMO9WnCSuD6AdQ2+u/rKgDjjEupdg
khM2tiiMcp1DPF3HrMDHWf16+UvcqZ0iKDnyPQyLCqG7xN6Vohw9nsjPynQlrM04
rZSEcMu8FnjvvpP9PJWUh1Ayk/A22NKzhhYogJ86OFLEUaUN1nye2xsVSIdgKgiJ
nGmShdHY5Q2RzdHOm/5yqLLg0gWKJJtph3hj6Sy/L6TOR1K3kY4t7fSLkBeuLws8
DZrnFh64igOlM60G5zGcrHi2PLyy7KlGO+GRvNhWy0E/gn4ldbB9h2j1BVmUYNqn
Qq46jRjhuX6nBNnAlMUFC9PAud/TkLOpfqtec13HuAwPNePh1i3vR+quW2QjXDYw
dEu1ugVtQrkvIBPL5zf4GcNlUpF+RVjfSe/nOF/STpUAnHcpPn27tGM6e+IFtX81
BY0meyhW9eeDLnl7AfPQSaeelj3QW1AKXXjYuHtiNEQNAe32Wj4okx4dZwXl2jAF
ojdAzXWmduNELd6VbgICyvU2z3WBNhLbM2leYLyxaymtZ+y1f1CfoZrKqNGJdRHK
W+ODGvH4x1xhn2MdgnxfT3q1x7TOtI1xq2ZJWRU9+ulWKnipB/lqtfEf++BEgMe3
w4xRdF4AAGcmifm50v5sTlaM3yH5rQWfX4FM52YIdEC53tpJR156v9MsR/gxb3Je
h52DOPmPRcubezMudbrevdGmTbf2VtOgVsvguyLd5qb3yq+c6fNtzPJl5tiQMsuU
Vz/FIFSp+wkB7yjxtjXrmC8+/WoOVEJhHozkX9CjK9gCqMEGok1SE/WPXscof+W9
drkYEiuCnJLCgukWf7KH0snQPrk6iAzRD1G5wup8e82WG/+7RDwcugJ8vz4E7CTZ
3m8csmXtlH0+DXDxA44dwdgo3+RdXFsjuG2FhL1QgwIc3UyPiY8BAsuHcCWRJ7W3
Ie+3f0Kt5Pp3lVvS231Cwt+FSP4prWrv+qNkOZPb4UhJiVPZXqsJmDds8OPC9pfz
3nkCzo0BG3jiEKo2RW4baJ8LQPlBy38ECV2NMM1C+2JCg6xvuf99aUuUa7JghRl8
5t38mLjenmo4QkkaJdO3PCEEE5x5WpI6ATWtygTDOGtJxdaIHDxXdcpot8hQaZBB
fqYuU8+kJ4WBvsSK5sGK3VSQ93sKaOmaOx8xKqS56Zy5h37qOt9xmrAMTHHLspvb
NtnLar6WNISjb5xeZNzDbzuuHJRInicxm3s7NrW/jTJSZpF3PQcVFD5rnFhExhN6
qhUHYQuUDQ8f3uJkIIXP2VNGcuZ1tjR13mO+Vleyhrz4UCeOrUcmGeRZYGBjxvtY
N92mWmi5/+1IOrO4EGX46I7le3D1ZOoWZMvu7tklkioA3M6e67CDnjcAR6Ii2OMW
zT2IcE0i5r2XmEZvDi6OEZjIIKr1UrZBNUr0u4KWYvvjMehEoGcUV/cCm/Cs011R
+QjQ/gc84RUgPn1MHlYXeoVqBSP30CdmW+VrwkSPNoAnoaHfYQUQKHZIH5CG02vS
jOjR2oOONKAF8pn5IkBf20DqNTAfj4OcMeUWMdqzcYoHqTI+AqOCQoSkVDotLItC
F+jcSOnKL//mY5eYcc3ouSEy/r6hHA5LaC5NMvEenIcKoy+4JRPrvKJYV73jQrkr
LnDKjLkkbdZ5AUTAUZRMups7m/hCJ/WfBde/imFC3wZGMaMzjsfRxPq4FbA3r8fp
r4kIRdQvyFCTFhQ+xwWo7vAaLDMzFoQdooOb0svh4eLBJbKKnSsWPyOfZykQFR8i
ZYRq6m2jh1MnsFkSIDWYi5tc5Q7hDXG2WbHmooP7S1fFUw3IPUliLWhscTx9RGtu
rZwmX2zYVma1vNphqwIPEe2Pt/453I7OvuQZSET1HF6WRzVdrYQxRfYt7ePmXQwq
eRCF6JfUGN6XXFSCG7gUzLjTWJLt7kN9G7BGJxNoeLKwGoaoxOGhXutBLiVm9LcE
DrJsmf412lAUU6qPGFVflsIIqOXA4+hNfTeQhJSNIVIJQwY0bHva8mhZ9BUeQfz5
flbDG+BakKQQJiCU4Nee7JfVrdsAbM94C0JzNUrWVXLlklpBiKwZWOpoxMdo1CM9
QU5LXWhYH5TXnzp7swNuOIbe1BWph4n8OBSXy8qp03xydJC92bpuX69RgphiJh5+
FscNkVlCfIhsbYBxHtUvkG8bVI7iCkZPea4UwMP81f70fr1LXpfsmW6mYMnXRUaN
n2fG2nUEdKIYiMIDk+Shvv3kRCSxXmQxyArHkfIKUAhPX6jbW2+/AJR+/EH33ucL
6JfodqIek9Cd3JbQ2t1t1um5AdK4SCBH3+LfQYJlDor6k4s+4qtfk5JyElvTAp90
3LejD0lP+zPloE/xBkmqsU85Y5HjB12xn0+V92+SqKH+aVodi5i/UpbWM9Zkem1I
+OSk1m+yi/lpcJaWGmsJwEuu+5Ke4VLKzeclbYO9aEHiGl0icwV9YwRti+E4IsJd
pduGu3+DUbptS/adbGbfYLVlFVL6xbIPrru8mV//FFnEWADxb0FWtG+SbdVJBchy
Wvz+W42D7bZThKwXMmilnmNrLVuoF/zKlqp20FApRIkaQojvKprOoVS1sEG/gKy3
bSAxABAUxIB27769rixLEI4objH13rDB47JijYwTkgTNTGlSNVYxCfLOHNbY59MS
C85cLDVLuWfqL/MPZM0442XvmjncLwqsfg3N07IiajY1FKXEqj3/fx8tCHwxfcL9
EB2uk2/l+4mToj6JiKIwm3Zl8bHCpnUjI4gJj6jgsYdVLlY9Cn+wXx6ZMCfH5FH1
EW1/VekEcbuXsK+ONm8KDvA8MmTrOtXUkpfHIuuml8jYawZaYbilIPvZaQO9nCJ9
fCVNll6+WMO3jDu132ahCfQXe1nHvoJuv5GM7DjZIsXU8stWzgv3eZ6MemoqSbIw
HjE41xxaqA052QAY2LeBb/0RZPbf9WAegdhYC06qf3wsnYjSLaaQpv8mj1RjvdlF
O6ksY1QiH9FFODiuYb0x0WQr3QZzIv7x9BRiq5FDYW609e6okfIp1XOTa2ZmwAYn
L4itQHAb8kOagGWfHEA9Ky7i3mJvdqAEGZYUBnWwuHpWzLKwun8tduPJXXQUUBGs
kT/QQK0zWCtSAxN5QwfG/mk6d+VmQ4ZZVtpAk5qtUncPcjMTJJQKs0aEvK1xJ6iH
q2bc1sPScOoMBwlPYfjIAKb1aRKQvKZFrQRCMgX7OulGKntMqft647YiWxF28bd/
LbBc9+XpRmx/pjA7kmFMoYuApt+Yy6HmWVkx905O0Ryt8w5MpNphPOXu/x/kpbkY
19IiQZd0pvMbhPkuO1yRdO0g5iNEfYW2frESCwMr0nERRg6CWUw1CtCHkKFLZWJd
Dh8Za7l901hhFUlFBCVtqlcV3zPs5q4AQmC85vf0N6h9MeTMM/x2FKleG5WfG0NQ
9mZEnhLaj/C8ySJHbP5LxxRM6v9rkzj2Lzffgu8u8qX27bXE3qCyFPTTgFAHyNq3
w0/HdaGaC+kn1mo827wK8yA2FSgqJO7NOEHdC4qDff5xnOFxJm3jBLHEFaXKALzw
HDWgYZgFZA9SLmkC4RHQd+JqS/ox+rFMO2SFSSHCnQV22zL6RnLgjRhv1I594uqT
H4T0XmXnk739HbHPYiHJr1eQHm/WDZm+ZEQVBniq+tfXCq4Tc7IohdOaZgzcCUzn
OV6sCD2Eek2UDq4durcV7TYFm4DaOvQ2AiCE6+WM5/9n7zRcKqwuLc3FvUQ8qWZN
92GzPIxr9sG7YxZAC9xXiEUSidFJh5XKrhqEr4RikSwAcsqog96/CcFkYWfAfAW8
L4tbTOrRfOL74yho0J8gjxuSLRl4s6HuEPyI6Hw8voZPcqJc4iBYc2Y9YWdvg9zK
o69NB73pQVPC8tFTvrzkGgG2UVGfHUH14Lnv2tSc6h/UphYFlv6RrJdbB4Pi/8Hk
j50tT1aJlCsusucSPDrGrPvSY+/6FnpQA8XBzpnO9HG50xt1AT0HIU8N24vrd904
7iF7HGG5akq0TA/xlSA+f9Iu7d34yd6cWIAlAvgyHrOepJIwzwlZhgAEXDAxvJ0M
0FkYmC1F/d+lfLRWASeH8Ij2B9qSOOECPjMHB+GPUMNC4lE8GYAx1addi0JFeGwB
nS0XeBlePBdDal5IgWc0RGOCt+lwl/Rm+CgxKd8/SJ33NHHvY9gWQzwXB8HqOa0G
LW86x7eEKr1mEz1qyKgT6nNm3rcNAY0DQ7c70fRJ56EYoY0h2cqGd7NudOkU/3/a
jgMmeUPxOBGMbIYGw34hL9JGWetPDpDO0qvO/TId9aAMykF8cP6rMdL8SYmtjVCq
0x6HJ6UdBq4asOqcBxbSvJu9DNZPWX37WKcuNHhlc/WzPoztjeA+uEdQF8KDUI2c
0Vd42W51PB5Xvhm+sR/BPU0vQtPa3Bj2bdXQTt0Fvf0u1ZThFIU0TpUxfS6mJZh9
7kdywdoZhD4rgz5oa8bFHystgsuTqG2vB9B4OO7bHVd29IDTIUUQiWSN5lwpdRXG
l+yS0ZA3uWlnPsAId9HyCmJ/XOIP88/CXtCSiVuexe7H7jTRg7HhzKvfL/Dz4i/k
SdGjpp9SQwfulO5iQk7I0hiE37W3jWE0Wsnf6Kvz3IMbaMJkWsEu2Mg6Wxj6BsOA
HwPz/k4riGMSUffxeBQC3C2NbXf/QBiW5LluLoq9W43C2K7WrIlD/Uhl+sfyR0z0
Gje4RLt8iSS8N4tC7UfrUPHk72ldyMxgfBr/6o9wMGfXqsUb2Hnw22QKG+6kZ01P
9iNwgYbcoLYX+Okktg69UgzRTCbY/u0jissmUPMAKJkLc9fxZQHrPjldkvz3oKKe
w6BSQOGdhsL9NTU6QwrwJO2mVhsjdDaD0fDKK2lQNYE//0argV3eKUUjvJGfX9qI
AhURwPiXtoHpQs0xN6na9DyLow6EuaJzT07xkx6IZe0B4x0bimNJJR7aiHNdpkfY
ypDBtERHJFZgDrsYD3Q5I9jEBKV1ZoGHvOhRaHxkgELNktBsWxPbESxPPCgQ6TGW
hvsucYMO14dC3zbzRVzlB9bSRUyTdT3PrN2TOf5HIb/EvqcmC+Y/G5se5rHe+fd2
K1Ku+qxrd1QWyDsZF/9Ml234f0gjakPN8xugsIDNp1arCwCrZfvi/cQ5GZoPqGQn
claiGPuVvP9ZxFMlNtBybVyoYGHf1wLzkCd+3lO2Vq0l25aA90NkOO+7UtvUsDmy
hZCsu7Qx3tIx0BVHHkbC5+GUaGrAKOxMw79ijd24GvtmTIKDmFl2YrGwX/3jJ6kS
D9GfA4zvTCTWtzq3jl80dcHnHQBOhpBOaXsemlgEV8sXzYeobpy+tbcNXtsYT50W
2KCj83Zqm3LtdhvBtvraXd02KMYIb9EJtN/oGfriOQ+UqCZZSS6t11eB4rEGbI/z
yWzi0WYk69dZS47lY5DAwyBTH3d/+83JMZMrceJp165ru8ibVeWdcHEOXyh6aMoO
W/k1Chf1PkdcP8KlEshnhNIWBkESD5DE/23r1zr1bM8j9daHrd4Enl5o2RDgZlZ1
+1+clPPj+x6iPt0lEOEcFcpH/FEKTuZg6oMaPxgMdObXTHBkD2ofd5m+X2bZve8b
BFPEfRRPnFc7X3psjGDS0MIwW4Sry7WiI8HmZXKlnudP/n9qnmkCG7qYKWvGkqmC
Q/6/+4uMooMnLHIyvhDnb8haVBc43MP1q6P8oR02Cj/f1MCAiTJGkIiqKpnwH6it
5ptFwyP60fsYTw5FtL/z0pLOa/fEgLSBYDmaEAFehTGg/bUMijD/frsTCthmcBw+
+PqQXTRisqpeKJi4oqMfNQAKNxDp5Z/H7b5wrmJGJFw4YJxP+vLlFh+1xofucfJD
Q+GEwcWRNN9syLpgG5vdDJ9tEOwTmCIC4iiMdsY49tFvhgTQ8HXd/88Kc2ncbpza
wyxS91olJQaPO49sCKFFhpoA548WmxqBEvolew6e2/Tunexc2XNXmuwJyOwSohlS
96G7lbBL9M4sTiwonQCf3K3xCVWUP0FuqClM6Mo53STvc/reN4UZVFsNuhf/InbE
5bAs38+Vr5qjeRTBpVk7G5NT/cVTNsai7I0k3uomJhrEoQwu8SFUUS31B3PNBZ1E
PWLSAtfYw+ZkxBO+Vp8dwGGLpdUOkaPbSlUIsuthKubPHhCOXH81/NngyRo3BH7o
4nGB1h+ztPc8rJ2vVN53CBhazPCZx/vWS7HVuDAq3dfd5V2FNnuS9hu4IXDS8D+T
5kmNL1DphR0fHPWQsnjnFU8YaJOrDc5ZdEXFcV0rhATCIHAv+4OTYuBPHGYBXhgz
IEGfvGR2PofPRhatzezEwbPPTd3iQwybSA1WOKX/GhVCPa3QSOUojA5ZGJnCPPHe
VKpd0C99BsBcnMsLf3uKb1at/LW6FR2pdMae4StE4opPGM22Yn0/qZT9v59biDsv
nGIGRbAFH2yYIrt3o4gNw9O2gMgwZxta+yLASy6a0a815rCD6SGYtDzuu1SsUKUu
e/43g4OOb48UNtDX7IDAHNnM4865zlcZckW87mcrduNPIe/R98D6DxuZb2FlsLgF
Bp50Hxo7slTXpQK+geUr7VTsXz78vhacaGKnPPyhZ2iAOZAt2I5vfbMB+Z2CK2WF
xYWHcKwOtSNtjyGb8NoSKWnrlPTVT0v5LuwMJEPWJx4MtDEaViyjj8JRA28PTW9H
aonhnn2cKAt0gT4HDK4IgldYGZJhY5bJjC3kY9r5OTdMDirZM3/n3UQnbcsgVpbc
8nRoPnGku2MZPITGmJq/UHnqxBGujo0HKj9iUv1E86z4ir/LCMSHwqY1qXMA1XBN
IcWWCMxUAWAb49lVLmmzx4nczNnSTUG4U3ZUkd+BoutSnwqcGM8jXmWyyQ+XiIQu
I5Sd00gMMRp7GIWiqzs20BdYOvqhSh7wz2JlJMYpOGqxARIP51T7I0sSenWOSvrj
ORRLqou1yLplOUaMIoJohhaDK3xzmUQ865m01+DOk/NvBQ9mZBSSVcU4FpXrRT5e
Nlpgk+TwZxle0Q2PW6ddFKJfxUtcrmRUgWqcUwe0+fJk7Vy38ENo7sbmVEuAkaoo
awEycpfAjoETCsEd0duG/YQftHe0hvKjvpcDeIiPspYNZShkQAt/aJOeD6wobV7n
CUpVNOfeFaT14YUiGTUTdBmof8MC3b22MuKQX1I6pUlnzi2U4ofUy84/66OohxEP
oBY7hHPhFqXCrO1NXCEK7YvLaDT9QzyM7eqTXNeZ5RVqmZoBC3KxvKSj94Hn3wpD
4p78JLl6ioUzMHlf3wa6DM135etA57vboxYv5nNtJZ8+VK50FVqX7lU5Nl2dxCZ9
23+uJPrwLYVGAb9B2YpeNhPwRhhz+W+1yzk0wLGzOBoU4LGXrofRtuPF4qfCQgWH
EnvKVVtB+f0/pg+zFTL9gaexb6ujWd9oBryyeqXZ0u3iuiqovnEU68un1+pAYSF7
wWyrA8/NXMqf5BROz8KO9EIQSx2W8ru6o3F+Gos7Ft8Y61x25OmSlX2HTb/q6yDB
zX3klqBidjnE8Tqg7IK1BcRAY9OVNBdxprooF+apUXb5PRnPMtvb/aCTUyzy3pCG
QbQGVemVixbQfzK3b96KxWTg7oRMuXD57mO9WhFTYbtM4hBHwz81kh7xf7XjSCNo
YQnVEdS3Yx931Z30pMD/6bZmfFj7o/Wq4nOmk7xdbTRbK3rWt8m/eBxgAZpjg3TF
6unHD9UiBifftUL0Tt6v3dWCao3TU+y6ZaWbRv+JCTbGGxlqPpDKCWCxkxzqtTI5
ISC58WWcE85cV/4KYupVxL9h5wGWzro+C6z7WEOAp0DDwWAkyK8kPG2rxppDQQGj
tgZG/w/TurReeNL0YtVECicHoGEB2/swq6gEO/NHD/kI3z5pyzh3fGq265Il4Jxc
Kk+yacW0LIyPJ0rMWykgW/sgViREvjfWoSmUvIpgx5GMuaKI1OtpJouy5yG4HmZY
kiTZYsukaEoCwJmlOhP2NTkIlIYi6yNBGQVIqPwLIfcJGmWfQpsjkBpSD+4oqm+9
t1YYC9q7udcO8hjVd0k2/if+2OyJuSaWIHVBJCYsEXuujmoTdHgKlyvMGwR+cScD
kO8rgKeE8FZvSzM/ZXhN778wxO5Vu8E7zgWBru20G53sDqTkziqqKhTcNRhXYqEi
t873enFiaNFA+UPLzIju1MqbHjHSVC4Ysch/m55wz7koklBKCJVDbn41PXBCVFKH
2Z+JWxqN4y/0w1GkEWQUAMUNRf4m1mR3vJRg8V6DzARPO80yowHvum65BUl0pHm4
TIsJPICl5rOQooIoypQ46JSnMaBRvenySxZj369qz16tZz0aV9NBfz0PXV0NxrLm
KP0W0ENzt9rCKfw+Beulyc6cvaIVmbeu2PmFytyjRcgI2IfN/kvqSVIh/a2+s9TA
w9XBwabZNDpKmQEMCd/PHdmHydywu+BDWe6ECXpF6Uc7kE9vtxaxvc0Va1r/YHGN
WLJo7ZiNz3JodskHi0jEvABheSsDiqmZO42x/YjLov4FrN0aCQVOmp7xbg57Y48V
j6JRhWn00sNWSwIEwB5Tg+paUuvcmU8w1dhCNio12OJpzRSsPrfSNDSZzdN1t705
Ttl9yEM9RT26xTyQj0EYsFnJSP06KmNdHCbJ1glNz1W/+1xkiUVdI28s/J91VsAp
agc1/Dvepz6oat4z/vB/1jWaOWv0pL8cgbAHpP8rd/U4ZoQTPiQSkos0dC4sEY9t
3GuWdIsUYlgKVB5qPH4HHMwJEXlB1w7/B+jP3B248FAAMMWP6S+dg5R7B6m3FgIC
jC/dHBf8z4nn4CPyC9XsxL+YcGzPFZwYxU5BgT5jy+EQIY1uSFeCBNiIzMoXQcs8
bAslvMJ/hIG/fKOvj1z2aBs3G09NwUjy4wPap5PVGiUNs2FHsY8JpVXvUEt8ZIpz
l/ThxUd7quyK2cVkczOuUDZ6MfnIHu3RSBOzzC8ENhsM80Mq7I3mXHNZwoWNN9jk
Zch+HTWRFkk6shmN6+cOCkOtqbw1wF3dnye1rc8jPg+QJpwpA3xgMU/QO1ERzzCg
y+pkX+1NNRrKJT6uAJeDgjxSXdKkpMzy29ghCsQBOhPrYqRA2YDy7zH1+hQ1hyQ9
5YsaVXchF04PwUTTsKYdQRFDSHMHkVS29Kus/yohw3HCI5uqI7YNGH53y5uZt4Ab
i22EUNFnHeEpypU8FnlbUdgem0foTL6NkOo8F/6rt4/R1nqvuVeYVA6JEonjfAfL
Pwg8gp70743FrKSbdap5wSroIz1Ddm5lc+w4SjsBGym+AmyyGy9WNSOtGrX11ADL
cNbLop1E2B3DtSgzF2cU62fgut9a4O9/c7juLQ1L9PXKpA8f3SvUehvWX9A8BKzM
BrLmNiOiNky8MotGI2aCXYC+fAG46KQSG8Mf4jq6ydIUUmFvDsiggRweOpK7k93q
YASCiG9cmL7iCIr9L4oy2TZ5lZmua0Otq21I3XSZRer/kR+pyOHUtbtadLekxitE
fjLN/y9YiGz7ri/D6dgYvFg8TBQlVG821beLDTuEIXtiCEjZRGTLg8Pt4zYKFkmY
00KRdXQ62HxRji3SUYIFHtHIik7SGp8WM2riIa+74a18BzTXtapI74RGLeSlICTe
OP17GAiS19C4CiSAC7ROd7Ta6doUEhM/Mug4LnqwX5g5VDuppJNPsAmyYGjec3qY
hgMyKi3Rn6FSW760f5lJbViRzUqEovUAbtFzunI5Ai2tmx5kAEaRTs+DZ6WzY7sO
SEdN5t0uqPWUDP8Uiy3TQEfTvieGdsXiGiOkzIY6iPn1uddzewNVukZQfG0Grjhc
6NoV8xgGxv/VrkwixlmLehYeeYORh1kE5ML7FxmP6BhFi79Qq+hTqsg4mkB4F3li
52Q2sgad941HesYA1nA4sSEcDayY6grouMSTJ8Hc8OL1BxHqE5YE8vG80En3zmbz
aymfEjuC/c71s+nWLzKkF3BKR8OO+PF4nWBUGbySfVjfejV+Qx07in/+uobJ49mT
C+B4DUPWh1NueyCqzYtFmnCe0z4yQHeJ2H6FYVovysfpCbrjtMZosGJIxuNlOlSs
XvB93FlXpxy1SXbTqtneNjk5xe8kJ3KOIeGLMxbE8M9QU7PM1AMNuWZlCgRNJqes
Zr8BgEMWiQLru8oU/f6kMGvKGZyGoQYg1yuGBPG6TIaItuV0XFX9sBK6Wzt+sowV
V0UzkVSOyi88Brd8og0Qqkfj4KD7EZku+QJNIIIH9NPvRo7PPOjZx4K/vRzt2IB0
AK9q2kbRsiwXTPydygjkXlsFYDbnRtG59z4obdVDVv28b9OaJNw0KaCeVeSkqoVy
6g4yXnsX9VqLfvUut1b0TnUZZfGJ9QHIdEar8DE+zeZJMO6P6+ZKHigu3fUQrWGp
KHtsd1NXjXafhTU6/DVUqSPRb238BHBKu4XpS8jl4rOGLmcdxja1MOA8Uo9xzgrg
9powgKS8+SpFEbnumI/ESdudNwVcTf8nrHT7/eaRT5adhSj0/c2m5+wePRspgYTU
97Z28W0/66E4k1X1NleXxuxiuOYQlwFUHKehMCq6BOeYoqCkBqlPLZ6ILgNGjTyV
PbFKGA856uXzwCrY1wqwYaU1/yG8AweeXVkhWDFkWfDtkLgBlz99fawdIYIHVPy/
46FM6ZlbkyCje0R32KIC3YCCDh0h2nv0sk41p1B/I8izjK0sFWMjFwddTtgU/vbH
AOH3fLHY/HdbM+kLV6BrgQD5AyJZxMFs7z0e/uVIxVksTjr4yVUu5c1knYvYbxXN
AsdJMR+qB44caQRgpvRRtu3I0wFNSf+PTL5DJoZaKfkZbWYVb6xdtw6tRuwPu2sT
yjtwfZ8r2neZRPE2DjfHOaIzBZp23E9aGC3715YT4plW0CL6x8TaWVlDPFLnQ5yd
aBFn98LMc2kuhTKGZacafey+E07g5J8JfrHHJ1e3BsjMMhSiGMC0JenJ8IdlSAlG
Pays7wcuiDjBe3WDpTCH0XV+XmTUfGvNzy1r/PAYG0/4wTULfiGdO2frjSuJNCa8
GV37X2zE3M67HldtU9KZHpq8XfRy0xS5z+v41YiWXRsTvO5ay1/7TkB9c2ZPEJfL
oGTYgrnDGVm/abj0w9GvWO+wLQng4saSpgs3c+3hGbvzt7PBdfEIfIsuZhKPVHLV
M8w6aj4jKuRyGoz37K1YyQbVj5XUmhBV3GMazVORD0KpFoxPBVQaa7i+VvbdHQMO
efUtZV/d0Sh+yqSsjDVMd77B2Ug3O+nR10Rw6T5V4eeOnitA1J3/D2tEep56ZzZ1
apDtxLpnWPxQRkygT8VYBrkSU9ZA+rAZZ6DuV7RfJoQ/Xdj5X4hdXn3Fdawg/5UC
b5nAKpw/2Vh+YzKJsUD1o+Z3gZVEPDtr/mBLTZEt/4EZjolR2LfZ8LoxmWPPOSSh
nekkXoHVw+WpwpdNnMmvSiEbzG4ANOTnnqxl67VsByekWFJ6dEk5qCLc7CsIVOiQ
/A0gZuMrliBbISoul/vWzTewR13RgYIfxnsMJxCzU112oO/Q9EzXUFPQfjO7S23K
/6N/BFgp0Fm7bTdffglQtlRG0hZtOtJeW8ZUchlX3VpKMugKl1ED3cHujaSoBnZ/
uKNvNlNTMjKDw9Dm/3tEpvxNjC7NiPE1WV63XGg/gSPZPIte1mpYRVwf41ba0lL1
NPRA6NsFwQYLAOcFKq1BUywoOdTNVgU+pYUEwmhkckY+rwj33Kb8O7siX6B+CE0U
zh/KH/kgmpvMgNbYagDTfmQqjHeI+652CF/snq2Ziu+C7TnWfBRDkZmKubQxGEhD
ppzPSBFnzVbTOOOGV2vsqmgc7o8ED6WvEzEClBqw33NESe+GMh5Dleilwx1ydn77
zjDjXmn9kGsVSzYfc76BT5Qr1HAtjQZv/JDEQUhWHFmiP09nG/IwMxQ91XKHnXRh
46wxVPAdDPhgIKHNrUbcJxCBQWMHJ/5zJIJuhzlV4Caou9RVEicGxwKuf4S/a65a
MdcBo1c7hGTkyHwgKtrMMmp+/b8Noi16PjND2UJOCrscp+tPbdWXW6WzR7k0Hld7
twr07GmkzxFipzBcJvKb3NwcuhckKnU0Z4UHwqoiFNhalS3KoqbodgMv59/TcLXO
l5q4qmOPlpHjTMuBp/mVIQBNNz/r+Exq2HBEWmyS76EyWZTMyDhDRgSDgA0Om12z
MvLm4U5tt2glTcYt+YNrDnf4Ahvx7omEud42GEYH/9CDK3YJQ3awCug5F+lqZaiE
uT39AxAcs7Py/MV7Pj/VedrNUBWHyRZG7hJAE/TwYlrJrvmgpyUECCdXqq0yYKXy
roULXiz3sOWO2QrjwkxyqOb73MNvLkcGqV0AruXnLN8szpFDL6fYKFfYwry/Wadu
rB+LDiarq/ukspbANiLogeliaOePMLxVdP8cL9zm8o0GxQieBrPy+LjGdKzby/Cz
JsxfR3rttcrakbVV3RBAp859iVpoN4ZEC7lynNtpEY27WiNEe6fGWq5X4unpX57Y
Mo+D1ec5CCBDyZuNW0us5i02OgEWymNUgc4g1oDkonI5h5hgKgdqodt1F8TDivFI
GPHB30g1oH/8kEA7VkMXDGeL86RoxITjErtBsRzEC8OWjQDRBQhig1150spOp/R4
7x8hVDgMxtoDHeNf8+PThM+ad3b4Q5O53Bsb23LmglPWhQ8aY9oBzVEXAJ4OGYp2
Hd8Z+8lzSFwOTzQikv1GeLrnlVwz2eYbvmmpY10IB2NbOvOsjB5Nlkg/YMP1WiFJ
HAHPHsny4o/I+Ih+n5P560tXnHvdt64qz/GOPyLSk7oJBgVXORdnyWCaY/vLJYK9
i1O3QohIvi63kglfKW5f/ZzqzTGOO9TdUdwgoxcHzU/ZAoWjfJg9rtVJb5vbb/KK
7gRFBNS/gIjHb32hVJRSSqyb4v2DQgwTlBtQHPF9DZrsqsQ74SSlON9UHbqReaiX
GfkhGh94cof3wRKD9AYHAg4UrQJRdKY6FDsTNPEy89ulN+Jc51XgQcWGBkKGPy2v
2unwnt05BI0eKNP2UsFdfc/Oz2P15eJWg62aGJ7kVod1JQNV28aeOn4mGnzj6s66
XAM1kp8jMENyL6incoLljZDK6AuX4M8k+ec2UVmQkMhZYhgA1rl/dxzkH/1JzeIk
aucuYZfNydRl5jg+dogl8KuXugel4sdonvJck8dhYf5OJXg3ogU4FopANu1r7ArN
7pFCTPW7rhixOXce578UFOy14CCyu9xSzhgwDZo6zRMJkpERknAkvza5q3X+JItu
EnklYA8IMSR32iqjZF/xFEpt9K4YJCrW+9HnWktD2+U/KaMoOkCmU88297dPuQpW
lbNNZnOx8MA6ZGwZ63JFRROhwv33L7NRBayhzpKReXFCu1zkg+JnbcfFO7zo718z
8I/O+24ASOzoYUjodAo7RoYYZpCvfWKuuZJ/ywN9yeZG8tZ327GQ26m9rTHJbKr3
Q+n3TdEaUdlQ65WKccJe49TgHYvlcFwcuj4tBf6hlMVafQgyJ5ofcpRQag3guUSn
pmAZPLhzerLkic0rwRYAtpQKoErypcoKPgsdge1J7tD0Jl6nGm6TYpyn4Id1YTZt
Lhzps75aKc4EZACcbYWZJwKVk9zm8Ktw0hrKa68oc1zdDmTAZfcyi/+jt5dHrLzn
fDNPnuMflizCuz7b/REjW3QiiQR3QDCtIsZk4E6fUQdtdjnNKHIftdXh+05CDsb1
NDQSso7HOkpJzm3KBPj99hlK/G5lC2j3PF4onPuYEE0Bhg7nfLcrGD5Em35HniIV
oSH9JDOsdah47W/yCa2jwW1PpRVfOZJd2Tu8niPG93aaSHXHprHNH1mnlMcWWEcb
qfqMh5n5lh0LjPm7CoFzwZM9zNccpgpntFT1iFKKqtUNf5rwuJ0AP3XfCvREsl7u
mcKjlvHqFZIE78YSzVq0aXkQzJHPYn+PdJMCABADL83+ajt5pXGFg2Mkc+UNYvg5
pdn7xgOt/LHyM/1Wxgffl8liU5RtLD/JqMAxx9GmqwGNFw890k0kxdAZoO6xqF6E
lvNnuL6g8DQiWeVb8sjPLCiXP1SrTdgnzNz+KIHnE9amZ3u5jBE1VMwlczdXI3Kv
/s4D7vVsvaffMUutGMYnJAY3CVwvXvv69MNMF/dnQAv603SIc+u7hQNck14KD6Mi
OWeSR69pTKPJn4sb9nfS3POI42nG/X1UKhQpbLn/fcf5wngxjJ9n8g5Ttq83jIMh
3TH0aooRD4KD/BL0Zd+CYK7/Mik+n56yARkWckPzPNma0AXN4HCkHBw0w/IxqaMH
5THLhIvSuuDpnZLqWcTwC4g425YDxLQ/wwcQDYC+QJpRXgagYLlsxQx/OV1JW5Cq
MzRxCYMJjYmqT/cnnqbk1F+ke4eIjwkAp6Zza1TXfdy4O4QswSvOATXuIJj/5o3i
e8JvDX3JYcpTwMUUAs+vxG2eShWqqaWwJgxA55ibF1A7JlIzbE8AiTOaLIAJQLGN
tREMiEpWDP4GyRk0UeUQQOT706ICYtiZgL7Ock9228CRtXLs1DDEJzpIupBLw9FC
KuPvRv0CcUSz1T0hNFgOo+adxVTgUQWsw+UScda0C/5zRB+0HMYLTa93Q/5Vr4vF
bhzeqFMvWLBW332FzGjomoOLZaP9b0R8ZGQjoGTWijHSjEwlvmma06wVgNaZJeUQ
XyqDEL9w+WzvkyOFoxhWdUpMnoRBkBcWRwTCXzOWJ4nQMfVwCepz7QW5oFcsUhzm
5v2BnrjDUajMNZV0Drf5+goR10mjQ2R/yOnlIEMfs28TsTMjjK8Ma4quSFCiZXuO
yPWqi+l+JbZaxf+Si3PZoeXk7ONDKIjouNchjFJZR43PR1e9yjzVqZ4n0IVa2RIf
QoRw9K1GlvdvK2cj3qw44FZrAFI3bu10mnYXJZwr5RmNXBj6NGefzObGAMqKzJbu
ao6+TlWuTcEb/WjosOrySSgD39/IQLDMMZl7tmngkzribix5/XHe9J3pEoGCiNRx
DQFRCUFaLVF3896Afmv3G2DqdmqP1a+Qsd9qLeUHXRSA+71lEeXuEMVSieRVlLj/
SCGQccXPF3PxxrzYs+J3EaoJjGm4gDhOnGmxXHP3YXXmGnce+JEQwVkiLbu3kURQ
YLbEi28O2CrwtjIaBtI3Ke71fk4ZeMiEfonSQWmQWftTkzOFGXhJ8YkPH5ynMqgr
n7zctSVuXb12nm1gLwkN58zNx6TEB9HH3b+wHheW+KVmfPMOYU7VxbgG+Zs+wvY6
l5xVXNuMcQj46mE5H1xj7EV2CbINDll+l+DkBQXk+Yu/rhMYOQQccXYHpN8wG0cx
E08//wAeCLwa3lD5EjElgu8BbBxQcaYOzNzt/3biIoTYbhxWUuMedG6HgxYMAFV2
Zh/yjMZco4rYMj5cHgCxNB2WIMAH7CJsW0gebNgwunVFaU2GQwV+laX7z9N9lg1D
lid9ueOZCGYhZ34hEl+DxxN2SxrvqkaX/rInprbvAkpUh34QgDy/O0Tz0bd28LOC
mOPyV9lvkHR4aeWpelSakodjRVX+FNbZQeASNAFLxSiOD5jkJHZbwqoa3t6lSPRu
xkOMle8ZTyFXg4Kt7bBHHJWz5t5RpjEQWFcjBp0bztama1jj9Gq4vkxYXrJPyiTA
4pZhXMKiwUVCMVY/XnSOZtJbmMLC9ErHIed9PkOHXCoC/J1gqBhWjrcnKiy9RCJD
sT03HqAexPtSM2Y/LfBkO0xBiVHHSXZbJ00k1JkOwHEdhpv2saIORkm0+sXzw67r
ro4oHZzm9AeV/KhLXiWLtZvCtZSV7DfG0yTAW8nB9BbH7cb+JEHRBTuvsGAZsKU6
cFyLfEhTF9j1S4kDKHoFkwEp8MoR5rdyw7vW8ArqfZoCG4oZjLAthLCdJ9Ai7MQ1
m0CBwnRzBhvQ1CrmNo2k1yfPf4QYEPjYbBTlxTlKGe9hPrxCxiNiOv0LNIq9ptPa
YVQu+jcI9ZdoaYMPZr3TAannVhX15ZbMNxx/3wQQ/Foio0ybY41s8IQC+kLq2Ew9
zhmcvHfdTaYUlVHXPu45J7C/PcQdcMbEwG4v0o/9+/me5uLC5kwN+/3+tMdZu/uG
+kYtnFiVFoPe8stRp/VBeQqRWJVK22aqeKMH7bklQ1vl4aYzv1n1HMgHDQv/BlUP
YbJOoCiWpccdKnO5scRzq59rpoUonB5yf6BEjogZ5M9vXyjay5qrN1aNJWQxguXX
GQH2cia2x/ETUIWsGqJL0P4iEiqIzbLpnyMT3Rbvpdsl+Yg84qs1MVuj8vbNX8FT
FdUqASW9eyEF8mpvqxhaogAVm4dd3KH+9nfCASrBsORnz1f9HGu3LIuixruBaSr/
6J0lo8RLvdHoav/9YSUu/VVH+xZWHSdINgdoGHxVOI9qyuYZ8M3PJTAzjosUlOJy
ptOkNGsUm1EK+eshPMR8IswMln2rODkhKDPmHwCNn6ApATg7l+WFoznjYYe3y70z
ygmyZ8otNunJcvSb9xvJNMx6RdAXVeYEozdsQcsba5chms07/PdOB/Jhz/6LrWj6
utlE9glTcaEhKnTF3F7GiixH69/GI4WkxPvnnFXl84nAL9XQveSSj5QgBF4ABv6N
e6TS8GNpUq1bJ5se4oMuSsyXAPz04JIhwhuqi2Tl+urQ7VCXwNDaMB+/6+cT8tyE
RLb0AlLfArW4iZJgKv7qmUrqC9Agz3BsmWs+pauf+nIpxCwuw98LYlLiLLKF8WQ5
lG/BlMMs/lme+QjnG5YOb1wHk9Y8eEaU4JDbKYYWBgNs5TjcFgktINnDUpFKmSxM
CW+Y6T6lkwR3h1O4HS+vs145Dp+KNgX/0eg36YZTEBrCJ6Ag7rh5M+a2CzreD61H
AqodHdbR/47edPNRwEpGiI50i517hj1AXf6KrqYOUuQb+3xe/b0Y75u/dHznHVKv
sxf1aJZRQfYfHsZ8W7bl7/QGqJtIEHH4r4g7WWDPFdjbH9IMMCZ4fop7DAyAukaq
3tKU6hCxWstLSCVupzIOfwjCkQHcZwSXR5UHEXiuvBFWow0p9tTz58tq0HuT5B7L
q7v0Z9YLziGKemwyOIi4yN0mNRRq6r3qbqFw/BD3jDXLIgNu5mKgFhMvTKGHpvij
1jWV5ZesloIj31QE3TTNGvqjoq/bKtuZu+rt50/TnaKDfXeT3ArVL7NfAxXPcTAo
r6GB9kMN6d4Zm9Vafaxfg7Om32T5BwK1RKVavEp1pLLB22ThvMfo6XkD/fo9fE5V
sfNz3e8z1ri8XhAAQNuFeQlRM+wvmssmjgVlmHTa/E01oXp2sO+1SuTQC/1j0pvj
Uc5xgxgnbP+GjteXXd4zrCdXzn9Dl0fgp9D74//AaXvziSK+9ltCLJOBr2ar7yt2
YcSmkyHCU22xYU8b4T4StOY7nDuU8QL6Mqj3WWdiMfJn36bZUWAu9qKgtADIiyCx
pHo4LLIqtxgB7MUvWtbfe27PveMZp0PCD8IC9SGW36tta9NM4h9KO78ER92Rdma9
cTvOmYLrPU8HnE3/r8kJXJ3lvwZO2Tkt9eQ8npJDbKZ8uQerHjZzT1Q02658zuTT
B9nO5l//V843zcOqCCuyqfiTLeKtldXhx6WFNdNMJPKw8A8PQBdWfqJ3oyP4QRj8
0jr6jtkoQNBFMD0yUFK0bhyiisCZ/qDtSR/bbJkvwPBPZt8tVMCVTYAETtxvqb94
mfqYMxu6ojy5sAQv39DRSiNSdqcrPl/kpEQuJqL4q+drOE3OWp7fO2HqJX6/P3Jd
Vk/eD4o2HmJ/6YVvEDVkAeCh716oJ/Dz6m05NOhuOLxVsFsfX4/KfuukBjbw8p3Y
zYdlhIsbWrqfpTOhnhPseoBnsK5xoM/1WTwn08g3bUKpNaN6kOAorlOGIAsVkh5V
gLW9QovuhydvVpYVEpwHrC+AX6YVE8/GunxgyaUcfX5wLXa33JKZ1w7qjqLiK3+7
eytypKHYbDMR/DdvyXrTN07vMKTIALzq+8PTEc32MMdxGkVhFbpMN0AMuQKLNeqj
iLTKOTnNoGn/VUm5wGnn8WC7YrfxxKWn8j0wPifg9FsewkcrhZYRp/9ThLQWOMy7
TMLd0vz9QgE2VoxhbMtVjQhMAKmMWwdC4kVP+7W9sfoieDIb8IBNp2tsWccbWJv/
Y7fPZFj1XhJI0zetuYMwDUkrsZOIwHwPX4pJ3lBxDchj5MvRK2SaE72s56Nv55uQ
+Y+eFwWzCVpe4nuPaC29UE6Y7c4lC7iLHYd4wRq31Mmh9mo7Z02ZPCd6UZ8Be2qn
vaQyoXG9K5cmo9IWfmYptsClZ6wdOfF23k+a/suHsagxzSsMBfG4imNVO1SM3OQK
9H6W5qN5Car6Zc2Ud1AUGe7FkCrD9yQ9CgL4xUwghtIe2K/hDcjpNMEMkZeInpea
lduiXn0T/KylyhqJgM2XrkxN6F1Iit5o9k5B32QPS4fZ0iv7PajwhTn1IP+TrfXm
AVg1bQ1P5qrDj9TPDzXGtC1VUTYGxu3BpMa69MdQbAbcYISMKA/1BCeurLVEaGXH
GWxm8+JL+ZKNXi+eAz8YLw7K3nVF4Bsc98rPyZ7eXaB9rtO0hw+fbVRTdCAe91kq
piEBUZg13e6S7IsAetB6LRc9qOUZGoGVZIID6RrwGvwfIndWdhT0j/9a0UoE3Q6Y
hZxmZNVpigDaWYi63A1evmflxt6WTJI7GwT6DXD8aOgvVay4h/Q+EtYDxsrczzEx
w+ukivCoAGqv4ccTjMyh5SUzp4Bmt3vUWm0AxdGT2kbyp12K9Orm8MAIvUDDkgJa
e9zFiYmI2REeRZuQOMy+jsRLEaV7al0+kYsANEwsjaWS15zbFjXNn2r1k1RYkSJp
P0JBjCpwAe7lhJ4kxHXDDVMM+TjEAUdiMFzzunaruzlj9A40I5BeW/t3VLI0p2lU
UPsyyyfiLRz01G1H0poJebUjUbhqLBCBvd7wMoQ2h4pR3qgoL6Pl/RLloDM1VPiU
mJq10dyvWQwYAm++IlkrLPRgveYeix1yflbHxtoJwqzRQK1GqwuaSd9lMxAKuKHm
CPAVVJihBNpQqJY7xyFhzcshKZDSg3psmVI8mS81TkQudwIgz56MdDi+BqP4XNWY
aUtdS/rcVc7F4c6gyHHvsw5SaMw7RVcWc4pCmCKvqROOB3jnrPHOhiKsYdQsADzQ
enl8AjcaRckQpiCl1TI/eknDYD9HzQahpi6t1j88L3HGlC/tWI8WofpJDOUEkKG7
T2xDsgWxWjvkSiUCXu8OJn2kk2Q5/gs+SHP3dHiNIrFgK2/LB/yBUt68tomz+H7z
2EaY3wx+jtrnp6tLcgG/okpIkIaY1M4Q7H0x3pJ4DT2Y2DNEL4rwiZorqVVvEiTW
A/Jw2Un0xMA25wntdCEVRYgcjl4DEpRCDV/Pw/lqaB8p+ZBAk7Jk33d1n9HLkDyN
Fy7t5CUdoBOky/a/rRnWUXiwD21G2SGV4OpVky82qvu0YLgEZrKHdQC+9PK6f3Ez
fUXdKttnz1ZYAdQFi7NZ1XzQbMWziAkl354aoqx5SmLpEKIucShsfvQTGn+m+qEB
J19s7KoMYx9LrRIHRfQEtXqdLoChh6GYuufLhUTF0BvLzDf+ZQF5vmK2cOz0Eh3n
p6LLMKCEk598kBRtzi31A6xvXH0EA5OhKwmqHXZH04jwD2CthCsqPKfsalzV9OWW
V3XV/Gyx8XHbSl+x9KyYjbbLUzkEjIyvQELwUz8rfkM7p2qSzQf0fm9qdZc4NeCq
PwZ+i2s86L/BgUWSWyPKGltlI7Ko/rHf69thTu3jma57dQmanvTR7SatWeH+OpVW
MwYaqTjDde7Uow09Nh73WAwh1UXPH5H9Ce0Qkv2moz9Bi86K0ZOeBc8VsFEy4aqh
DaFyyUysLsRMe8y05TExW/nT5bLvkANOjX2XucnCk2rBT0rOod2SKMFenJu+qKsv
qllCplKPc8MrUYRrZOvX8Mh5EIY+VlsFEFIAN9UrayrAsl00X0n/ae0KrfZBcR9q
TufH5hfrqOHYNgmeLnSxviwwclO6/kQ4zYlJa9p7M6yUxiqh2eLUMNtx3/kcouB0
LEvW7ph9EKhM0M/puuCF5iP5rQyVD6b3G8Jl4FAXxlSYwH5YQvv65/Ovwxz3Uikg
GN5uP/ATU314tNaRC6doLrThi8TJ2eNcaLZCr9fNcZsFHOdKHjGlo/hiVlTXXoTe
YHwqoL84KnNCDoFnbarnr58bkwspI/8kRRpcUJSWDemJ8OkCChGRMtCyzHs5GEYv
NgOf3hAudApanPr2ygcacCEuezvBmlNF1BuvIErPGUQXOYtrH6p8Hdeybjh5aPOW
fD2PiXv1XLT8Rgmc0L8Z/sTvz1d91YrFZpjjoiOVCGMnTvSM6EIPUyajTFwLaatr
K50zmLdbqb8juI2bWDTiVyonN1v+7dhsw1J74wLhtFhspO8HVtuEpLS0xXUAV/Fj
79L4TB9bDhpoP1mEu6JiLLamwI+STZ6wUs2GkkVN7N2WOFi9nHk0llqZ0qamIxui
Zq6gpKQMnfB0LZ7OMcutK+zJKOk8MzwACJHnIDgAZcp3qSNfsLWYD6jbuJMnjwMs
SoAPzSWc098MVl3yTWRaKM2YUQlQv2sJT26BCLsXbh+miDB6iJWiKYjafOA/B+Et
MhyLfMTyFqPivfaS2p6ke0RGsGvGEqyZfp+54YkCgLPKYmU65quhnx6T6Tz3OBRu
2qE3GfGVoya94/F6rYcGo5XtrtE4tvBS433EqGXuoUAXtKRw/OIhZPbZzF476duW
1b8MJ9jNYUuGvqTLP3IqI+p4NaY2JMCNlL5kzIHvY9k9bEVQIH7VrEoP9yfJOOEg
afdAcPWwfmNSqi3ogTBQoDJ9JK3pGCHh4zYKHFrxW8EHjKfKxLeJ0SnqzIt5Nq5H
tK1jULxyYOTjYXF2hM2US9N0on4t6y2fDO70kW9oz7GQFwvH/AwomYFzLirFo3P2
1N4HFsFSl5D55K9L+iP7YWO90gtqAjg/Q7C/CbtM8wke4dTB9y1vSfFIyLJythM1
aZcfjZbPbDNaqMfDXFL2wkxtyTA+wzISNNYZ2YgXHtwV3ScTj9Q7yeIlTwhxnJe6
itXJRhYDVgaBHQZGWmNNRmV/SofSV393YK3aAv2gFgxjb2+q33EAjqmiY9Jk1Uwf
FDR4oH9ojtdhymOfOoNBx2at9jqVO7bKE1ydVhdW51Lyp2Cn2MMaEMlz42YHq59Q
BYf403e8Nd2unRzw0v+t/1lP4ucw299ghgRVhWDijZDKXwASttUv0zVFv0zpJpgf
AY4sW9vztpcZe5VqeWBK4XAT6SuyLmcKmXPuYx/FCLORyOS8H2SrAh5VtZdgppj5
Z/RBA9mGx/BaDfr5jmuPvDDVxdSpgL0Gc8lxtr05wmF6OPHNqs5HD3j+SeM7SbXb
dqZ5qy5Q/Cv1d0rlmWDkoMuwr0bkWTbKBlNBr34kenoW7XgAXGxWBd8jDLeXcxBK
+KFBQ+FwQXMfakPiM038XAxHhz/t6g71e/M5XmtjIgY1e9pwjLm/VFqDI8ErK19A
jZO/BPeg/m/sT4uXmSnVFJZfQd0hoShBa59YYg7NyTMWQzFmZ6bvXCQ8M2WKLzmR
4Mkt+50wpQtqE1V/gsuoa7Eq4kK5yjmupqU3rKejrGkdhuCRhEawsxFCujju0nBB
7hG1Yr0+QeqSYZVTFCG4hRDORQwl5tS5Xt7x2YF5RmsPJE35r8Rmpb+3Nfk8WoTc
MedG0Lud6+zUewBdU3gVw+EozOYQh4lRCGmRCq+/KCANRcULyR3xJzgJIXop2CNn
cbmgb2ra/wk4mI46ufj88oaMN0SlPySd2oXn9z8wqbs+svRL462Hmxfd+EO9v+IJ
U6CWj5VQ6cOxzQs5D8EPAhqSjNrwvbpBfC2QMD+khi6ncLtaCO9pacqyTpSw/Rj5
hzOIERepbSGHvtIGxJlwWYOHe2DJdKmewN6j0WMjY78N1+ZsKJWr49l0354qF2iV
meCvyq8oeleNmE3+op4r9yTIzps9pWeo84m+5kQm1uzUVMf6YI4MuEQWIF8k3mlk
DlNSAFtlnehDRbJjpEcYQkz0W3JGD5uBR1J2cXLcZOYDUEiAGPJh946aEk+RJnaa
Jl+nWrv6huCmmLqukObmat/rE29CoR5aqtg9oy+beEmGS70yFkdR/jbIXOQq8uNL
joSWKH/uSeDYWoCC0/QGMm16jIjO8HBXIMO1b06YmuBnBPLQ3HtV8eW5mZHARW5Y
C7X96UWih5RwIr546BXyqr/K5E8N/6RndTLPaNjw18o8NDFtpnmrBtq7JRD1rLLR
Q8vf6WzkUZ1pZB2jnzciVb/hht29b+NVeC6U14xjuZ3hgQPxi/C2GqrZ0Jj7vDtw
kGud9RVxSTQDRjxZbTpCp+AmO17IAhZvPdUiqVEagB1g7O76A7NBg54cbuWHc+xj
21evhKjcINjbmdjv7yjHTjluREaiLWBOk1BScVP6zVv/sV9cgO6uPGZp+klzm9Qu
aph99G+xLv/cD0+2ZOj33c96k6qwXAd1yyFvm/WmMKQ6niEo5kMutVjO4c7QZwv/
PoyJ3+hPc59RMHuXCq5dqDKkbWE64iARdNHOeKTyApB98kpDU283rlTxkgeavtqd
DUh92hoodBn9ejno9f3HapT0vbWsPqhIdLYgp0b4rRGjd8PuhqcfNcKhBoRxZuoy
7k5Tsk6Ql4YiUXXpC/BHMYFGE/XDO7yjPvKkUJZMtrYMVMzilk58A5yZ+paSHnUS
nBkrfx//XHWdkjJZJLbsMg+vua1TahTyQz+sbTR4cxndDY+bkhhHcHt28wP/lHW7
K7WshVfJXZmPC7TIXLkF2xdpDxMT7T7XzSNNYAIPH2qOSACNLQpPxKT2QRR5sueB
zhCqucwLiHZXFcotZG7eM2o7xLLAht2F/CU8SBUs1wnQBNtaO7+yOAEgXMshAuNU
Qdkt6xn8ARsexqT1z/ipEcMDjBMrzq6qxi2XDHQ+tLd9Px1V62Iv1UfWXzUbe2FN
Aydd7WQ+Esk1lkxmCAiSET+RVl+3ROHuT155A+SZyEELT57x/fb4LXC/KhR9yZMC
tf4So89PFClL+L41/BhL6qw1rnCRvheaZZs/ZcYW8ieEiY1vQMdn9s8nrrDl2AtE
Jo5Dfug/Vg88ZoukyO2FHyWuKSEk6CnrYyo6Ca3DJJxUd+FHyEefBT6dPyL+oMXO
Pu/I4hlLYoe+cIIcsl4VW9zwZSvgj2yTz9E5LxnQnhcYUrnzzz9kg56pd8HINe0Z
osEuwTiejCOGKzj+qmbCyu7fZCEbsq49udPyqoqfmbFFrSI/UrRX+a4TQC+RsVep
Zji0BOg0ajCYN0qu9EaeGTFUOX5gqI9yIw3JnJfPvxxjuu0xNy7ukvm4fc10G/mo
3uFPm7iYsd06YoIrgciQCMYe+uDhQDlc9fZ0U3T19OpuiweXyQZ1Rqb8bOFSYz58
2/I12FOMIV7OLdxdLhr4CBDBs9ulW+GkY6bR2PaR59SSjV1tSA3PCSIGNL2rhNml
CqVF1OT9+2Yi2qGnZvCCeFF0ekx65+nxdeO8e8W7Vc3wqtHar41KvSFWuNTrAU6f
He+lBSKk/NNeTc6nyiWTJ4pqE8Agnge7HOiYWL4NPFHeVedNEImkELRXAsrzrhCP
ZafM0wG8SsIsK4PU5fp5/iHlh8Ab0kAaxrbn41G27Cwp76VW67dZPiDbyDdxJA2c
HQMUBTR6RXJ2xiWf2Pc9XAw2GD+fiMWXBPUqT/FHFYLpjjIlicXLVqiAvOdbOqsC
kgH5eg3iVKtUmHFbmsKY0+ry0Ey1P4hXi3d7h3qoNsvjM1yBBeMvlbwumKjaN5Wg
nDP+jFJeYhGY/C/eLAmMoR6uiqiOjR3ATiZuhkcVkrQeIcvCeS7QexbIp2+x9JND
uSZafeRKYchvLmHYQZHrD2bL81T8YDNs5FJP1gE/udDQ7Mx/SiH/FrT1qomVBAXp
juxyJhMWpaP04oP/zuJ6PDFMYZFza94CX5UWHR/LwjCeMGWyADEiTdoqWh+YzAMk
BNPhH5CweaTXPdWj8N5nsdn7nIAYByyXeS/B57Sj/hWF8aYJa7hMGEb2hox5jlQO
qKt8Z/8AY3uzVPxGUa5eiLUOV+K9i9jzlbfrXSQWaZXELq0bG7q/tN6EL6BHotV+
CTH6afWFEsjA1cgIoQFchNC1J8+JvIM1/LO42Cdg3LLHSA9AoL0FB52GpvdFqzTg
hDL/PkkC7uwFWR4jp1Yfi244jmhw6+SO/PXDTYp7S3bqc5h6hGrFHC8O1IhLH2Nc
uRc41R2DNRJPi6MSxdI2MEUf/0n96Z3+H7n3gU++0+Fd4nSH0We84x4018tez1OZ
OwO+bfWvXV9ddagr2tjbYLSjvSzN3j+U2kC7ZvU48Wll7j1vz2CCm+POROScePZn
yNkAkySK6W2nxPr9aj2jxwsmRoWAUybPv8Im0J6gekJJY2cmS+6uFvXFPDs1FI3t
ugVf8SJCziH6aGI8nqaBunYIQ6KaKsBuxw6o1NXvF4b6pTikpym++/FtyQeeUERW
0QjS1e9aB5oiLByXBhOBAqN9+0QIeBu4yp8kfKPH/xoSTHhSCvL+Bc8M3zRd3Dtc
Hd0Dqt+POP8XRtP7oZzrP7jJMrXkMz9Bwxzmzvq7Brds0Cbna52oVHzB7920gPmQ
HSeyCqDUgB8F7bZ/wmku6T3UhR7XzOkowdsi7aA2CdfNH5reEE5RdG1pKBulC8wk
bm9xjvv73bXFy+cbm7gvB483Kc3/CUcenH51eEdqCpbSaupwsTIKUneFHqyMEnao
Fvnb2+9dGmbEsQBgIBQ0JdE6IhF0B7vK8Q2ZftNzjN6yy+JvZTMQjLIj6mNe8SAj
8SZ0KcAhWr2C495sRvYOSTVtyQS/GlnJSrZCpk+bkMElWKenApOREJmeiQB50bYA
R0U9Xe7nujtx7ZRjOkP9lKEFwcwBOeDNcY6nU9HIi5Ydbg3RuXvUb4ROUZCMvrIV
ksd6vLtXFJI0IIGw6uJGIVArlBU6X4TwKZejtSZOKbGy6sFhP4QK/vykMlKLi4lo
Yzi57OPno2dghue+2Wj5wmZ2wLdM23eIAr+914LJRqU/CPtHPXNdECS0F5qgLAxg
KQy5OXdCsM6VIE/JadXhVn1fVhmTjsyVB7MbOP56dTJvfkUfcyegEvxiJY38FNO+
6WM5TbWsccSkHbWXxEaDNWVpbnneywu1vFBiZUZcl4a+RzpFLKoDXQNzqfYG3OMR
oIoUN+TmdakFKfylJeiqyidToLUQlYMxfNDYq/MSthNpTVNbgsruxl9zfICC2OyY
iM7D23WEH8yy6U2iT0w/Z5sWpqCOI4IkdWBdkgGqJTPdFXFbYmJhQgwnH8vl/tTF
Qxlq2uWxpcWGTEawHfGWLq3LNj4xaor8aH8MzoLjSMF5d1zLo2QSCLXkbouz2Ra0
bOZhk/vr4Hp0ArAhC+Xxj1+pQBjgGC815u33/+b6CCBiyD5g4RoAm4fQ5wctd5fG
UiNrDNtgRr3bwZpsVJlDb6LBjnmr5+IeWBgMCZO0cj35WthaPC3ugxl3qamv8sdH
erBhoJEr3tAq2t1vyCMbmzBZb7RKbru7tXv2VWe+Atv35kIY8E+dtP/PrtQhKB7Z
4oJI/f6Jogo5+IXiseS51eokXEIeolPicwjQIU+gk9x6pNuQFismr5mUt0uqOFSH
aBndDcYjhGqUd41enw4bJ7EmlOwsD2x4GTFuMy/KqW6qd/mCF+YcbIlkNNevgGkQ
ssYVFdbabBHTtBcjmRi+KcIJtOqp9Y70DZyfNJzhz2GKSojIR9i4ifOF06du/OPZ
IBnR9PTJlNBSe8UnVF4zNBWTqlOKgB5yb+RmYKwRGfrC0ySBtjwWhtBGVSlTfgg2
tPWk4IyqvqsfGYdrj1VJdVkcTWhPJ63MJ9503345QiM0VBZyFscsNtBQZXnH0ZVw
37BS3eUC7jyCA5HerTL4rLdxWmFujYAKlOzJc36ElF4ID/oFQsmX0U8c+DTUFbQ3
OY9MnaB8kDt+w610wOPcST2RO2w7DzieNC6ZwMtUwbwgLm5z6c49ujzPzv0bwWC8
WdVVj/Hczg4C8+b0uNOgetNMnMyZRlkhbcYWgjwwLCCWOiQGunlvR6xQ+zP2fV7v
SATchC7NjVJ8EuAJyk8Q4RtXSj6Kr8E+Bpj8XsnXRON6gauBVxioDiXfoBFqh0Ac
29FfXIF9SWVu2mx39iVfYJgVSEkUO+CA2fY7N7egdQR+Qc4W3OVW4cH/CwEMEC6A
YFWAt/ZSf/CjE+jt1LZmEeoKUKqipofw6HHqOOB9obj97NNYlkHAPWIfqmi5m5AO
2ZbP/zPwfCKRZjj7/WBU3dE8GoHP9FyEdXMlG5ahd1YFaqHW6E/Tx0md+5UlNC9v
Kbzx+imZ1m0G+yJm6K8mMHUDyneL/jkosu3F0JDNxBquSAJ29b+zltrUXF0VCo46
cJvOSDHCQNyLjIPn7o58PbwDHkSLLJhVTgRH791Xi4T7b9vlTE7CNHtq391NGb8M
6Clsy/cH7Ip2SUZRmdezyumqYc1dI98ZXFAATbKVycWFtbPEpHIBVwATQitVq5qg
Qur/8WfM9uqf/qAet2/me70yvPHJ+8A0S0N6InUQsx7bDEW64P0D5MD3OIG8nMA6
xhdknxxDQTGhHz1yhaqasjinT9YGyFys5KO74hyk1g1Qh31TgGffM5TVCZ7wG7QM
kpnUrwM1eeK1cIHYw4KIPKrsDHMsQkXSrNcXzxrxHdAsLTfOt/5LwqgnAugVQCiP
V2cQokbGU6GHa8tiEjZSubq7N7T+w0CfwEM8S7SCqvL7/udBNF8T/x5G/c3MnfZ2
6aPRXTYUDI5//PyhhY/57BTM55yyc96HIUMJgqdVweTFOHm4tbzKMdWRUog4FtGA
dvsWSM8n2kKvhicE0FsVetO2PStHSbxNXXNtxMQH/7I8o+AZp/t8kaNb8ck7bXQK
cqc53o0ws79Iji8qgxHqXUWTnRCdlel5LISRZNle3aRPyYiTwqVlSSvYMUlP5q0x
d7JYEoXTg8f+pz5Y1HpH4b7ytbsKxUl4vSAwvtF625wUOAmMOPPibja8M6TxhDHB
P0SY1Jl6a8YLjAq1dYSNvnEqKSKR4rVFM6BuhHksndAzcgLz+L3bUTAupExFYeIu
vx2EoyAUnFV51wEOdl8Aee4DpB1KA8FlozC2AXsNY3HrHhagNiR3jd09vvw2ML61
miZnK/jfkC4RHoeTCTlBGj3TscOs5rVlvEhhDXwIvm/+H/1VUcXAn/8ReJO0iWwR
LNHgb0BA72CDLWgKF5W6ueJzpvBMrjyZ0zLsitsx3vqV112iVTxh60UUZU+RQofd
yK1eKEB43jjb2A05rzx4cTFAAyspkalrl3Mb3yBbhi3XBSQBgtvfSYHI8YFWdarV
MzeuPRInxzl/565Lh5ulRt/58jch/3R95Ii3DHyTLwfBx6M5uP/talBKYyo35JaU
QTRCrPfZ7yvNrpC8EpCoqNetmzX312o/5Ktf9EUqgqEmHb8xUVRjXgr0nwJ2o5e3
wHyUN6bBoohyB5veMlB9Av7Pj3Zc/UqHlMTqZ/VbbVPuy16mkUHv44RymEsdq2sX
DKGFu2YThurd6v/Q1yImpEJLxUUBCImGamT1l2Rg+1NZ50xGNG9dcZhjupTMzE5k
iRWnNn70mMrZIyuY8xXRN3m3tCUfssbchVeamh5ALolrQc2frntNRlz7Rtx4V2//
fKY7gSUgoad6whkex58vr7V0L5ZGf4r8ErquM6+1GKmaNok3FX/5QyJYX3Gpv6J2
FjjQFRhWOPAOw99VqGxwmkLngUUESQ3LpbH6VFdx+k3PVykhpcY7sWBOAIc+h8bL
HHd8VW28Gduwe79I6jGV8VsZq6GE2j8I1fQ8euBM+LA7kkuVfvD6LIeATPfsjjMV
/Kn7mXJiPIg0cfVVGYaf1UFTeOdH4/zyM3PVhQGiefJta3uSitGp0R3pRFAkV6gM
FIDDoKt93Nk//SnrjLCumUcnOatGcbqwnAakVspSh/eAVxLlHqgoPZcgY4S+Smvy
DDKEB16BolCMf7/V8amWjAWMsz4+P3IqbOLc9WFj8WI31avIyohq6N5QjqPdq7vY
ozSOFq/mZRndT5dAJN7zH53zwvCv9lqJ2ZNUfa6wOHhCk0ePlPfpoD5McdbbmrkK
D7Wcrf6qteuQEOruv9Q1VLxFrxGdC7mvyaZ7bCL2CCecbicflEh/XJTEsulDidy4
COar5eQJoLpIIIYOgZut/B2GQmQoUgCrzB4xRa4KNcWvwnn2uxEfBSxlw7/5RlKC
T/FGeyS2kQ2hb4QXobOt0Uqc/f5xINxNS/bVbWfUL/r6ZR3zwLe1+KwogLdQib9h
Dsc+cPYyyfXhlui4xGnLlZo3THZT3XqG5qB09EEPQSwFXZe0eBSYjBYepb2uvbzK
0toS51esm/vMvsegZKMd/eKrdUqo83tbJYZiGTy3crAGjhfCq8eKW1wqOYzODuJj
A1I1+gpHe38dgLJ2sVAefr2xrN4m0JALrEBZ6BJjeZVQmhp4hfaRxI3VoyO55Zu7
56AaJRYcqtpdl/ByV1INGp7zpT+iBSYSotQ0ICnK9ZCLko1H3SvWkjXqmSMYm4rW
29tKtBYZY1GoBTDqU6by/fV0/d6CTMEOXefFAh7Egx2f2C2f4+Yckl2TXaZ7nXYw
YRBG/iwN1Dqxw/73EJCM7y9mmtga4ZCzVii+LvWVAt7SoEccg06IPto45iwkeFFa
D8E/UgofgeDANLqK5VEehJvbfXhI76jpe/zfOLO2AnpwmX4QXMsr4gopBqhKkMoI
kB14GDGQQfVQh6jkxzHwQyv7CPCtaoCdB934a69O0kArT8cAk0sczMSoGXkM3tEv
MwVzcjaLWqNdSr2XgGvzm/QQQO7K+qX5HTCT5WXfoZD1nVUD2WZ1JYshN2VaIPk+
cw7I8ynEaA+1PQiSykdK6zMmoukj/bH+SdvoECcQoweVcVvJqPCVb/mGX4EuoDSt
bfA7N7XmUJbxw5WlPXiBLee3X7JugrLlJSSESAdkspVigVor0AWdpykzLM6LUhXe
IHAuhVEpCXKBRRQwmwQAW9hYi0IG8S+qwebiBiobCWcGXr5aYsTb9zszCuLh7gHy
s11O2BVf+UYE9ja4m5wLPPw8nXKT+4VF5WGLR9acIvNVGN1qpqncwgdxa3D9wjaf
qPIY08vIZXkj6XZDSO4sefZ/uEvWqapEV2HsvVAYghJDrOnhBAGAONPL+UUKDyuv
ECCEBiW1jCzpvTQujZKE5693ax03crTISF/uVekTn+D7FUiVoi6mJRi8w7reCa0r
kLhKk4293qIhch+HXVvw0iZRMmv7NRe5ZPx0I1yYiLS35Kn3gWvYQk4WloWZ+uhI
98ChiaWwNunthI1qKb7aeReJ3bQeENVxXOUruCtYxVLsvEBr5T0MELhoBwN401+n
wYrNx0heps2dQHNnMz13q6rcTpExP0w4QdXZpqWaJjuZ9LQDCcLEbBe4kcQEEqnv
Uj2LLrLWCjMciVh9rZzVy1oTUrFnUBQWs2OfsSlDcR/2xjwyDIskcr+E9DKPC1n0
kOz5i8vUtEitrcSdBMf260x4Y+sI3AWLs1Ksrk0O1H5v7aSAsYNSRv3dhyVD3GD9
1qKf+7lz/0F7P2l4c6ca6YDpmFFtvyG/cayJlFb4rJxsj+gjDNKHdjTxsEnopu7K
/Tf2ccirNmAznc3mK2urUu75fjFU0bZowu4xHCktFLHg8RgX4JWS0PxuZgHPLT7c
AOKFGVMDtN/s4odqm1/CbPY4CMlrcak02muzhJBanof4iui3s1cNyw1WJo+Wm+H5
5szdbSg9J4yg2QgTR+S+VRyZ1wSOl5f8g+XAfaDw17Jhg9Uf1zh+F1WwGKXV3VyJ
wZAtzNtkc7zdAqqz5EnDMbwfov9+jQ/JC560POm7Ds839hMzLIDjpPs2Q19VUh74
5WjK2Q+2F3mIyunTJO5YbKK6ZoURK1qJevnnmrPk2OD5yUiJr4EJvfpEbZYltVO6
7FrNssfbjcFP4I+qeze03+a99YzgiaKfhMfhMa8IBsZwBmZSlhNx8k3QsHR7LWiJ
I4R5G225VyT0E9Fn1el+o3xzquJE88vmg3Rw+xj9g/iNRpUNASQgsPbk5QsA/WLh
xz9odEPmoRUtBheyB2O969FAi0Tqg7DHPYySdA9h00J5qel8urHSTX/hFEGMDRev
GD2WaNB7RUNfCW1iJVM6CBiQzQnQh65kxY3CaAo/7GvYm5Pbuw2sKTovCdz0ToeO
Rv33b287SXIQlXEgODX/T5h/MGTul8bzDjdCiAzhF16h4uJFnOjrpXDW5VhXLAfK
zhmY/lHgRZZzk4mU0Ob/VeudNi+8X5GeyBJ2T325Mksk1bPNhiRDbm9xoI8f3wNm
LhlC7nQDc2/oFwB4b6EtdfxfvfkgBbApIQbH2SbxURc+8qlWxAxJmMKCPo2AT950
43nyCgMsCXnUrUX0SQEmiCKej3Q3EzhbMmJKkwu8s2lUd+y511L+F4ZIdbXGWGCk
TNEcfGgMFsPTPM/krE741O/89LPrSBUZFpVM0kJ6o5tOPjie5skXRkjQaEFUt1Lk
ywo6/7POWy0wazRkm2CTxdCD7cjmCNmBcml+LJbbVfxxC9tWaXx3oq500ltVpZPj
/usaMTck6pWZn5H1anbJgzFoQCF6yzNQQy1T64eMkZmIh2ESRmz7fRXt9m0wf3N0
NLN6ywl7w/KbjD0B8L2/65zqUmcKg2UNNwmL8VPN4mJnglNfFAVu1X8LYFLKnhD1
Psa6MsH5jcXxhHk6lyZHG3dCRNm7uKMMH8+n7QbS54sKKNjesUF7W8VmgwlNoinV
zGPqgolaE5oK7vPFEQpKc8ZFi6viXYI+8hZ9PD1ifSgqSOQzP6HpBKNsENBlcUQI
n8bjcn2vvD+oRQu8q4OdtSd75bh9SDxrlpzot/xNvIlbR3x6uicK3TeaYK7m0Ytp
mpJ/07X6CeRP6/2FgE9l5m5sDfyICCGAWAPg65oPeBrG+XttvQTzWrr+Ly6CZ97/
luXpTGL/hZdoj5TDc5pK5jyw9qfEcq4DWhHG0XJJdKDkb+pV6hk8SMuO0HhCnfCo
cqZdBE+2KQPsJfR+9fHDBg8K2VcdBvXN0ssUu933kmqZKj8FVMQUPRGdLMORCwNv
brwv5JU3B53AsRwx12qEdSR6fLJYzN24Rq+bStsyZX25D4ubQluCxYgbmZKX/MTI
eRoY/4XYaNbBlKfRZgQUxsiUVbcGYNbNzasrKPgFCmxAZJG+oIQqyozK/rMuv8dC
MJ8ozyzMyj8oaAvfS1Wtn28M2Wn5f96NkHa4jfpIaKytbXp+rdzc9anrY0GDM9Ix
7zOa4PUHdHPIZ+ED5nsjXB15O2A9lvnLLcFKKh8dfSl6FLWVPK2fB3AOcN/tiH4z
qZkT0j39rT5TsJ4Rg2t4d5KgJJiwQtoZg8juIwSii8zmHvQqe5CZeZGKJnNEFMzu
yzp0QpUDEDdUf9b98k5Ss3FUjr4nK79dkn8q6Lr45p3e0w8eHQv08NTBpvHSRlHi
MOgfZbjGuTwfQMFOiOfzJhhq1zCWUsJBqh9KKVIyPRv65k2hA8QC+0VzIqD95i+u
nQsYcDtc107JFmNDK9cQFsUpCvyPtP9PasTjaeBigOzKOe0iVO+6XbieSLBDVkgr
xQrWk0xVDYAmL5LHWJ11JVy2HMH3+cZB9aG6gEHqg7D3dTIoXaxvo1qSX2BtfE9+
drjvVm4GMCy6m6tw7qx0zDH8ALqQYD8aJfEc3G0nnldE/usOG8e73hMDuAePMTLD
Gc4XOz6dlc9dinFIDLOPX4M0ZbOoqDpmmYKPq3cvQukly3TRcSHQbOLFcrST7Mm2
NBOVhYDfze0So3L9yZhRfSSrTcc11WaWwqS4QRIjvfSpYyxqIUHonVpeFlj9HY9E
Suz1gWUK0Dt26acS9aGe4UXV0PngJdMw3qYwC+UPcZMHH85dEnk0YLQUrJHtwad4
04nn8KMsx/iO5krdXuloNQI1m6WY057JxvJhYBknZ/0VjvUEqz3DJb0+FYuio+T1
mKJhGuvZQLGqXdnYSOhufh+cu+JSUCtqmvy3EJFwh2fnl88HL6+HfVaQ8ucUSyYn
XlEH+svGkPg66Vgw6L6T0Tj6QKGgBtdnjBXTyuRzhAOMcRw6YTbFZVotjd1UU4Og
/bjI8BKUklByqpbcQ5ypWd8iE09RkL25VHjtsOLs9kZLEvr26055+O4KFhMFqRqR
B2eiEv8NNm7FW3yL7H2j6gaR1VWYd3aTeBxUzrLFeSKr/Jvrh0JPWJn9t7zi26sN
eQX41z4LkwAdfc9I3eAdwqUNhklpvB1O7Kof2fzAxXvq97qWOYOQXoH675dLqGEy
0YI5ID43gYYPeUa47tFMUooXd3Qr0skGnWomiE+vKrQpeu1A36ghUk+Qi9Gyv+yw
UP/GHBbvaLcaW4MQl8CnvQAvn9gY+dQ2JnXU8VY0pYlyv63nUOFh6+H+gILoZANB
6/kLYiOlJWFmJLi+WsSFjbFvc5vsMjuluXXx3ZQRQc+3YfN/CBFZNHhovL75vADq
eW58tnOX+oG5nOxm+f+hSagex2RyeYj3X3J1UpGhL3R+uA44EXQJpf2gSKU+UYE+
FrSIZ09JMFh0T5pXdlOrwRAM/yuFz6/1Uhk9uAq0ZjfammO5vinogvMcPREOXpkB
hGzq9nIXE66cGiDmEm3IqtX/V9useTMF8gbaAoI9v7Q+3cQ/um3eZ5rxMWgOFIq8
hLRtiiyXzCePud+yFVXWiBB58nnxl7sJir+lFTKtYBjOMFEXmrYvkhzNlS0rihEY
7hmDDj3R5nJsO184LuqM2j3fifbURDn9gMxpMcY9Coi3pQOX3dDAr70SxV5YVZ+/
rDapM5XCgiENDpfu9WqLLccq2m1Iyzy8vuCANCCJTqu6X/i36IC1tXzrPl7ovtsh
sz6S+xrHezTnIcbrUr/s8S9hjBOrzA8DOki1vNC+ljPQhWeb3fIh+6xLIf6BSJ0d
OG/SrxFsIPtDX3TtXJuRFjpFyfAAzFIqUDIupiQVi0SPOJFfHTwq9HC2kWFsvSTg
b9TkYHBhpOLiHw1m5LmtjK8zYwNsHboSaWub4yqbmwHTIg65a+rRPaxFxxrI9Lbe
1n4XXjBvTTFBkYikCYR22oNRRGmcbzeP9aUf1kM+UHnBY3F9w/jM/b/8hVONZQSj
egOgql36kBFjb6ax5LEg+696zpUJ7hCNwq5HbTjPA+3D4WhHtNB7l1bVD+vhxNCa
8wFHiZW0DNWuqSyCGx3GX/80OROqDF1T6AMRKomQW3omkxtEYEu+/zYBhbZJ7VqP
xYm6EW2Q1oKrCtE8cCiVhWzfZ5IGZxdXMsposevBXV0hmhIkL8iVhYy9KwcfVVg3
HPPxC5emHdInurXNjytXCMfVZEvuA2h5j/Q/ZYyz+GfSCMEBFjhC1HfNY8EgYvVb
f1vwYkpgk9aipnQ5bdd0Qtv3SbVEYarG4n0qIP9XAifWGJDvggLPdRblKB7bNIS7
zGxOi8a2fBM/NjOiu0yX8y8nMHd/jn4t2i0mOvKr7maibyHG6bTDozIL6frcJw7d
T4Qm14tras/SSPGpCMNz9PRebfEVuNEWJc+VCL/61e8edC5n8Z/0VrzUblQZEUnC
00TV2O/DwhYtsZlnxK5bdKjbekfRj6V4sN4Stq3pFBVWD1JLU/EgNTCdV/nR9kae
Sq3wf4WQNwfc8exQ9DCswSzNZg5T9WphxgYGk/Vum8cTrsS2Rn0epL0a1tcAbLIc
Ml9z2aWrIUG/9fDbtiHMhw0NF5ViD+z4ZIge6lqAvkXp03vdRgDs1lSp+G24uriw
mK0S16zbxXUS9HDm9pDjnpXKF/2YeHHiwUf3JEUQ/nrj5tw94bH3QIOY7kLeCA7v
aT+BY/rbsGe7C0cUpgtdngjZt7i7A/66DC0rCcoaMr0B710bYnjJtPeZYBiATvJA
POTLm5lh7StJWPmZyelMULOkjHt3XOg9ba1eKFEOp8lljQJQ4uD7rbZUIpW5aZuy
Bv7aye+Fd4Qua/m3XhullJUVHxVejrsBa26T/jW1EMiaOIugtnp1fERLtLObvsvm
DxCnIk4uGiBDgp3CD9yfqSerlO4ZTRJ2s/bICYVnhm7KieTWr3aRb3+qMA0kZWJp
/r8Afu/Kt/5shGwl2N/gfLTKRUOksYCS7ni0Yado7yd9xGNBX/zs8yx6cctFY5w5
OhKMAgUJYSq4OqexG+RG7MJkC3V+NXG0dv8zigd5SUHhpaTAQm7nPxnPq3Rt8r0c
LmkjukJ2wGrDbAQfhF1EpXFk9CprITWeeKZXSkbkH1FT3fJqcNSZrF89gFlp/iZl
Ehl7fRH0tJVfhBr66IJODLeXAL+Cj+WHRuuX/05yMb38dhc+iOk2HDQ72I2Sv/YP
TMRWngS6o3qZYXk9SVDd/ICF/POEZhYjXfJP6tm2Q/x+ljQz9QTKaeJDCmOwye6C
BQtUWOFjWFMc0LmytdpEKIV56MkqhtEpO0Zg469MlW8wq+obVqGae9ZnEsbBlt7p
509BhVxXfHeCeO5WyQYLNP7a5dqc4aCkDF/g6ABuauDRFAgaCHCxwZqRae5+QjCq
ZTj4iXFhDmn+TJJkYYElCgbKx7P8LOqJdWpA5mDhAE7QuvjFIZ8QJJZWRr9h+/ev
d6kOyGZBf4HTUZCrhG0y1Q//QAloI2kp8UL+YEdLWI+MSUO3R2GqWxOTVHjoDbvg
JgJFK9JJXEa/omKT9DcQJ/J0EZOzJLBUXdIHLXqSqmMZyFU1ahCAq1RRDIe8xm+3
PtiQmWiKE/loLojvYrx4TZpYEeWYLS76ElEVQE2lqjT8BpvGpSzUfBDzysgHVwVw
+zNFIJ3PH5BnBxle67PZvZHj4qQW4qoLZT5NL+BBzzlhBAx77gRiqCGmDPOiCQuU
YYEcT8ojyova1+e2BRFP9293fPd9Barz7KJ4dZcHLdI0pFyxXTlPIepPJtg5tmwz
iwFKwBYP3xyeJ1M+ldhjF4dTJ4UaJzGlbf/53VbhBOOO1B3MOs5D52C9isAXQ9jA
2DyExP0BKo4yIirf2WmzqpGEzvRoRJ34n1fOt/a22PuQkMtzwMdcsXW1tJNNNGIX
jDE1TrdhgJOupMCOunivlTkUBUYsru9uaHb00XcAdTN35GvKVUwkv1GpyeuToDk0
9YuirZFRBVYoo88fNdSP6Tx0l7tKEm9G8bV8akcHz1tMzr4KZYwBvM1HYXVDHwYe
JRACl/etiLAsIZbv9IXi9gABaRpBkfwGbGw7yYlB8itoxPQ5OzDleq/tpHAgxZ7A
CmxG+A5K3FFPGgWEr3EJFiG2+Vk4qccXBCZ6UXZKYy3xxFALQNmllzBenwGMq7H2
4Gj6IfWcMhb68epa2plpKac8yoUcgYqCcHScOHsBT+tc60m1RR3rMr1aRmDMokC7
vH5m33xD6wULC2StZSr1FK3mAsj2bcfKa+yTT/Dzwb6lgqjgJ8UbeLaaZ7lKUKXk
uIbXhaykRXYLaWqwt4LHmWPamlt9V4Ra/OxVTtS7pN/Bqsl3ohQdaWZKP5aETj3g
MTHuea4UMoU/C4MM+S7bAKMoypQO7Uk69G3fXERrwRMqOFWTdB1F6XvwFGNDYJLO
eyzOwsRShrqXIJSk1JNt/G45HAhfJfFagPQSJZLWry0vjzXMEypagktxScfOe6ka
MBIKKAdcw+hKMcb42hWvgqhwJM43GdGu96yh0qWJrIdHK4mPLb5/UhEwjSraZaii
lVjRUO9OxAt7YosnbrGhTU6JBHgmv0+qQv5Z41c/SrPBYp+TIxKtsc0/sB5rnfbq
eoj/ATiT3+V0drA8a38V1sySsmGJufqwqskIQQJSzqqHPcxhqzNcC+/frHJGYe02
+vHr0FM3eVIh9iRwOtWwaf2bFnlPk5SvmyL7PrDN15Byrt7pzw4V4qoWlaVqtdJN
uGViGmNgy/nmV4W7HoOQNTln+AaSmgIgdKK6jWuItpE9M9pZhU0CfaUWXZlOC/1m
YVFnhitBHU2TDh4oNK+498Eyt5d8ikT1x7NDzDe9FaR/ABauBXOK+lFEAcoLv1Yg
YUoBHiyx0cmqzcp56c3McyTUcJtBv9to696/fmn2/uW7ylGWqxemuthiDwqXECzf
Whmrs+SW2O5F6Kud3yBtMGehnE/aeciU/ehMPvjzhXaPS6hy6fRtfIy8xtgcHOcu
x+4i1v5EzGi+NiFilNuJOvG39GT0qorAMdtHYT8Wyz2/8K3IG4lxXaTO4x06okA1
l6fdrtnflz5G47A3IscxqCDzZ8iF+GXsVODID5aMheMSHdaEOvvjSsJF71RVjdsq
YHippn24DuomOcXBv82CR/50H0UCDx4lwI3U8XR3v+lDgp/qMsNoNtofY10Sw7d4
VoOYZycTF5r3LGfwoYc1u05lxzgwl+QvIVuxaP8nYeclPSoF1u0cbpZtqWmN/mP9
L/G7plu/FOZ8fe6fV/lOzv7FYm4GX1zHjDvUPQ8xY9qCABO7yszbszcV26NNcgUU
BqD+hIaKEIjKFnKACqD9LWX6ytJpgIZYWStA222koPb82UqNRyIkP3JnwNdRsBGb
qUVZJb2Pfb55Z80iZ7knEE1LNmiu4UcXZy4pt91GBywsR81YRTTBvo4pfJs5Uc3x
gFPhXly5G57XHAHKSVoW0VHuqW+UinxNFty9oEHrSQ1w6/eTwFlwFBQb+IkW1EBP
jP5Eb69SbIwSi9RBibWmV4FlxbMVb0uR+0BVVxn06r/5P4Ny2tOJLoaIZTcpaJo0
j/DUoyILfpFhOXJQGp6xgep9XJoAe8hjeiQXNgMrLYR54AoF4MlvEgdoPuDMxSqH
jiU9RN/F1THsgIsdY5icZPrm3C5Zw9+8XSCJg8zG1ssZetFJdbRkvHVvLE9b1OaB
9QccPkBoYv35atpJ4+MNgDGVccTOgNhDjhKI/AnxKaJauLlqj4oeU7d1jH1SO4PK
94QtdebtidzHzsmXF5Roh1CflqSQV45RM2JoOZe9zngn1eA6N6eSkTMufgzpsDLi
39QDFlbKjHI+KKCQCrlv7FqF9HxDF666S4JFyRmxxnZIolCw/kjUPykPeW2QtGQJ
+/5h5PMEeP6kKguWYYlmYMtEo169XZp6ic18TEG9JXb4fQ3aJXOPPb7Im0a6+QTu
fuiOna+zx9Divso6O1qY1Qx1/vLoengY0e2+MK5Ir/WlfQKy81z+PKQgG279xcS1
5ICY9RJBOV1i+eYRrj7bPKBKf8W143OZS+9P5Cky9Pofm3q4rULO5cu09cQY+c9z
Ws1s0fhNg1EAeBAZYjvXuOhkiaioECe8FoaFr8yAenoW3JolRF4WmgIMjjDKlpeR
37rk/OKh6THzJNVHBtlzDQI6zCEjdbDODhxT82CsZrntxiPHcsShYa0NwjB9LjLd
/883PEjLkAl9htQ81YeztM5z2eXRG7X3MdB57oB5p+zibK/BARdmfKjVAj9djuD8
/s6cxojprarrbfnRhYff/qzlX6Lk4c7n4hLT+RHGaB1hQsB1MSR6Fj4iBwBTB/G7
E1HEghaEOQAgrBOvY0jG3iPnBCe0F9vp6bsr0jqj+dcP+mOKREYwfXe5u2PmDAKk
ZrCIcW349YLdWDLaaM2tG9pQm9oJPTjEqh1OqAHhZEQBvuYwHh7afsaWU9BRH8qF
0whK4druFmyMOABXg8AjNgEFEJyEJhg7bn/WOxd4XehOEjBMS8B1JrHwlcMWgGFz
5cUfs0ODR5lX5kG5FRIYBT+CZrYX5iYw3xJodtxbXeY2wGtGXw1NnKXFxG5BM16Q
yCyyALqvyKnEpVP9CYh+TiYgL1F9qHxH7tSm0qc7Xt7UCCj6mEnRSi6Ob85JbfAh
CMxsA7zPpUgFfTXwaNbMbs5ZtIiLoiTK7HKq35XaazeMQ+N7LvQfcUe69N+g/OPF
Eo8+86/DFFlOnB07Q6fsnsQfuthqRN9oBqEPqK06Sh0w8vKluZD1RZNelJPOMm/Y
Ojq7NKX+OvUyOGtXGvnLdB6rP5h2TSsPYV79fnHzNWbmaQt3JZw/jkJY6CQiwAp5
ZI/Nno5SK1gC7UA2im2bhHnFzJtHkubGVsAR72Z8AalmB059Sq6gBPzLZFY+/Kmo
db/xDTpovHpsFumZ01DXl2y8Dy+ME6U5kPbT8YtkMf0t1uIlfrGPoqFeHiV0t0iQ
zWIfqmQSZqDgXN0h6zODfm0N86+THUlBifYksueCZDnAcrZ26Fe8F8Lrb8D7pP+7
3kr63s37BRfB6Q/OcpEYR4ghISqgwdDd26XUK+Q71F8CTfIoWBmSP1zMP7bYlDv+
dVNlDF6RWL2et8CspZqkngcr51nghYTT/ZdcFZgXiWZX5l4qXFBY4AE7Py5uSQgP
e9TW1CdnO51B0rWZWMTX/J+6KuftFW64x1igXVS/H9pbZvv3zAFMy5s4MZBrX/Fc
MtAhQyWAdQ4iEzU0wRaYfL9L5xGPQ+1rAe/Jf6Xf3PQHS2u2v1xa2dgwZQoI6S+3
crlZq+1q+/FRVGcDMp+RJ8vbr1xnTw6bXJAQuWWcpxiKEz3i2xwwQEhPJerA5D5S
x5jiFE0TYOhDIBCbOUyQHpSBrrQ+PfA0Ul9izM7fuJnd+I9cr2lE2mHBjzs0xGXY
zEGsQRhSNscZq65PWQw3RvsravwVmoRCfbXmqufc1KUaYibBR6cgbbMXcgBder/W
Lpwd9S5fU/XtCZP163TR82CPxIrVLK3gaEsg4h1ixtu0cfbIkdF9vTZxPOgYwubE
94n34OzF4/92A2aNyjI1by75GBnRg/tMT8/mXyD20I2f7/JaxryHSeLdiON/L3EY
nMkvLtMOqpHxYaK7RW3Lw5n9VPmcZCpyiVeGXFhZXtL/ml81Pb3vUwE9ycePya+s
sdY8q+9bQX82Fi4DSfBy0Mu1PNetJJVteyTHH13/SZlLATW5pXRH7xGo3ZwJE2VR
/0cBkvUzllnRGcAg/fiWjuCuRXNBLdg/woHAYw08DBki+tmYsFlF3Jgk03XtJNVi
0LjuYOSnzu3BeBHecs6a6tDgIaekr/dBEoS+8L1ng3K40gkpY5mQC19XzqBwcCGl
kFruIHXGflSXxlddKBygxkDrZ7ai84mBn6CtcR8WjBBfgWb71X10YtFNBkxdGEpX
1VYj48eijp7omkfUmCo1F05MZ/7819f6KyoneRZkI6u2fEqUXxTbs0F+6aahUOwB
z2sFWWmnbyMqLsOwEbDz0egu0Lz2qCKO13WyynIlTdbr0ch5Obvi/BcHfbiWE6qy
kwKNhOu1shBbzE6sdyOBiCf3kAWFYq0F4Ie7pCDESveYvj/yJKbauKcASejPmE7F
TtSDOiey5kQxD2qNoHXWQGP9UK2qGQIRDOQwZz6uankBAzABYRFYTkZcELUI9QO6
C0/OXalT1DT4PvEtXs0lop7BTA86J3cSHLdxGbSX6pj7SKJGWcHH7sj0UQnLH4+E
7rItXg3XABJNd5atm91IxzxVIeWxVOl7oRF3xCkuHSWFZG9HYK3GMIFU6iTL7fl9
uTHE/5MIWpv1VHPBnSkiw0zec33c5yxkzaw3QTxiMvj1ltM680wvH6fCF9m6fLDV
X86X4I9KXyhnJhB9XM2FPd5Wgq8TOpsj010z/zet77Z/AsqEP7GCcBp1MOda7tgl
Gd7ymod7/A79CdC/kD5nuLEABYPSulBRDvhGSEKeD3su9xRm0NIrALLtXwNHSLo/
l2SDO5MrTGhhagkYr2TqbAP06kpK1P5o7QMCiJogEJqa9ONl7Qe2fmmfJ2buTeYC
Medp0V1pZOoGjmDpr0+dNOd6Dco1Bs4yJrp0Hyi7umS8iD0duLJbZqmwCgCLNaKB
T8p71GhX9OyqbdLBOoCO7r0oCXe0IoXLucdTSGmbtF2C9crL6W1BaVQYFKSyXW3D
+kobn6+wn7NB0ngnLrBqGcu8wacS2sHN500pbT6EzX6dSWnTlzbQHiLhbI50vx2r
03VV0ba4D4wFxX8Lfs2Ez5ro+LCaWVxP1onTm+PmE/tRDQ8w2FnHnqFYCW0Skuz5
4u3UgB3d+sUe2j5by/3EbOQksbIgul6RLrY5r0V0ieTJ1LWV94BfPUO5HxeaBfRs
axewcyF39n/VUshT3Z9iKFCDpuqrqK/5LuFtYhL3lzUg/T6MrcnzlLWxX6mG0iI9
fyRTZe2NZuSsZqBhtfZpLFB0uS13XP4x4JCKbU3cw6RoanQg+nIoe+bzC6EL4IrK
2bPH18FQarDjafh+W3FO8xhkyH4/G4q4xCsok5x+qfXV8P9kShYYKPbmO707bt3/
3uABuRYXHMJlAFx82XMzDso/SpkqUB0Hyx/EqRjtq1xWJID50CPjAwBGB5gRHrWT
sbnoMGSxxQe9ckFDyJ9ACMxkw5ar6PEa0b4FRESf0A12LRNmUh5hLRzGKSefXmXi
VrGIopGImmV38BOTesHy2yIRb7GvPjGJj8Y/TNcivXzkG4STt9BFhr2YlSl7HsDN
1pXJv3K7rSKapidzt4+Q5/rmbdao/KlcDTuSzdsTjmKLfJU5kIZqE5cvt1xzyT6A
Wq3hyoq6sNY0ioEBDj7BkVby6jygp4kw4DatbymcNm6nbBR2QxJwv/xIxqWLrgll
Xb4BwynRjv26eWNyIbHdWKHw3tNcajGJynIe5zfMRoRQDB+HNEBEgFfBN/f4DmRA
UkX1dfeMn+awC6mXDRh/YgKJGcMr/SNF+onrcJc7lLbOidQPg5LKW/jpaIDa7htO
aQ5Bk0HRaldhNlladdNOp6vHJF6IxYT+GIjhNXJLEQwMY3WgNnP1+En1ZQW+xxIJ
cC+xDJnd2aK6x+ZWIhRHnMb2bMeJhTPbekc29x8YMp0BmHnoyIfnm0sQz9fvc4gF
6q2JuTblROFSFb/ixZWGy0DnXCwidoY0F+OHECtWoU3kteqWarboa7QG2Mvg6Zna
qFMra2geQ8PgEis6JGtVLMnQ8sljZQKB8cHpoXn8z8Ch1Y0U+uk/qKQHWVi4xlZ2
EtBynftILSyC4BVEVzQMivNGtxNE3QhRSFysaDG2dSaGpkVDdvh5EbtE5SrlExW9
LVsr8LM4q8Otgp3HyHRk+69I5eQlB8te3bgXJuHGZyZRFo2+z0Zz6pskPlDPAsAC
JJMtH8TTD3feWeuY4BosYl/qBksG8HPTCWuZfDKRoO2e14PKiyosMJdp9BSf03Q1
yvAB0XBp9+0VDZpbdBj2yDS4xFfcCtd3BAGOY+sCKRx04ejng9Gpg7KN21cIkTOK
MgQzsjAcx7X2oDDzZ9idflWvs61MZ7lDv6pxlLwquDqwmLy0IsGjF2SkPBReK5Pb
cmGAA2fS65FBxeOwxJAKqZGFfCQOjMTvcEANSuOOxjKT5ADGVO4hKnRzBo5WMolv
/upgZ+G8Rm1iagaIvJJ/Xc0OyHDM5h5jKJMok6zoe9QogJmWmxYiMRrD7jyahT/5
50nQmlarKPJEC9nBngRmYBhy2u57SGhKd2dM6H1/SWR6KpOnIIqkKBLredmtqG4I
EvcZE9cRN6eYjQbkgBjotZLRO2owxDA9AXJgoFDDBLzpii4F7jEMkkfzd4WdK3iH
rNF7/+73o2wqqrPIr5/FXVFC74dqaxJIgh0tzLvJNCak9QqeilI27oSvCRJX0Kee
WyEY/SE0zZuEixxkFQwK57cAf7BXzhGmpKPynoD2x1J9W7/Lziomeg8g0OL1Ls3d
Bz6xao9RKtMeFcNorqapWooY+unH+naUs89Qsl5Rc4xGyG+bXX9HypenX3uUAsSX
K9p3+/CHrB/pjsQQlxucS7Qg5p19f3R+u7YPXGm77ryNXAp4Q9QGpfu1Vg7IaCr1
qB/V2CeLqBmPetw4JI87DgeorTleH99DuaDjLVKA4zxn1EovVmOXf2gBxfVA7ryP
2xg/GLrqqiZxXGT2pncscewc9PhRaSvnEKccfBxs0abEiZEk66zQ/dZam1tLnkb3
AXIYvCl7Hd6flnm+DX6h1/9dV7E/1MykvNzHKZFnKRpyH/4Ohp8jAEg9Q5ZYiYJx
WcBqSg38zjC49RfmwNt0VNC8IsAy8gF5S58UHAx35KFPGtIobfM1CMIXBo3gDrAy
AbXwI/dWEK1qoW1PGQtLNtsDLJbO5K81oEiZjWgLcbfVR1F5ghXxv/BuZN0jf9Vq
XJRHTsMf2egv5Y3HT+eRa5e+TWp1SpUi2vJwDMr3dJ1fvUgDVptVwmKM344kD0FZ
edCg7KJEBwlI0JRhTE5n0siIBNMRmQdByecAhw28Wi4bqSFxtxQLCMMOt29wJq/O
L+Mk0l7S2XhuuVA4Vv9dzz+TjOQTex99ga/UmY4QrRrhAFmz5s76gEGrV3fq862M
zgTXYEuLv54TF/V14nv/mzpdI37nhKUcGTCY7g1Y7xztpBrQzIO+tcJn8CIXKbxy
JaQ93h6CCi2+7EI1JYekoAttAUl2A6aCgO2dY1K0kR/H6LeVLjPCB0dOycWnYd54
Re2k7i1cwk0OSGW7Zfbb8BAtv0tWhJP6r5vfcTzJtiRIlgwN/2CHotCJ1lxejKAt
HZhJfPs+dv9UtSxQ/ERvbl+P6nFaRjxYXZdap6gDA5rAC3pP16Wwu/gMSlPjlYrA
qJPFNUXAYGZCi235Gelqri6bx0OI0wMnthXmMKB/ztPu0AqeXsUYuaHUuxLcCCTy
J4aPMI8JGBevC5PuEVLb0/buBVFT3AY4rCUfbO8PbLD9ym1hotib1lWBe81dQlvs
Ba94vKuhUas6yBcn3biCxEPFG7uUZU0KjOFO8MiXPCtRFv8sBeFBRQHn2x5Tra0a
StGqqJ71PJxbrBh1APomNMCnFhA0tWXbOdkl5pbkeAIUysdeiQpehvplcRiB33xT
DZulAAUDYhADR/RvZJvfhz/nXWir2Js0pGBVnF1Idi9+skD4sJ8UFRyWQ2p3hLWf
nwiD0Kwjr+Iri3+zKmEddZ/Pq1bRhpS5jQJrWwIyD4CEksRGmUeBUpS3TN10DyJ8
bPQM8QjpC06cUHBviig37m09lkDKX+gQYwwiJAYNC8ECrZK/rGusVUAh8ITFDhFn
6vQ3bSMaqF7CN1G93v9bsrNqX8TYkvJ66apFBi7nZfS+LwyCLBsSjTP5ewn0/Weg
1j4U0eiUcHRbiKIGySZzMPw01WotcQ228FvrmWYRiH5gcqYIDELXqetcto3RZSUT
Uk0m8ej9Tfw3WobBfDG65AxygTwV9CXMOG1zFDEAwHDzi7UgZlcS0Cs1poimKmLc
lkoKUlP/SxyfDTRMpyAzX5sn+BMfg1bW9lkG+nMPgH8NWhLyCxkE0d79RVVxdPkq
emd3128j3hsa0C5WSyQf2LCRMYppXIEJT2BguZqlLKPtn6RHTpjaOKoxVRZm8DKH
6oKgdKPl2bJNz2EBUluURzFzMAkqKGRhMzukflmYW/dkM8NP2AYKg/PCZT6FmO0Y
rlcP96donl39Tn5sAVf1FulAvsMX4IcPh6JGW7D7mjNjlRLhLFqjXNGEJuPl74rJ
D80SWUIxPB+xGz7XKbhVfc9a/KuuYxWyd1V9eOk/6/1CYyrgZBDHN50+E6FUYctA
LYHwrkIS28kl9WW7LibR7siCr3Xs7lxwDQQ9ueAI7/fKIruAVFeU2tGmqaX6dkYI
6CXXV0BLHNJL+Nf/ElwkUB0fPUfkOY9rsVJnxQNcdO6UYnkEC77egoFKGLdIjmlU
tjm9m1WpGT3IIJfCuD8Y8rcez8tQ2+nw7A74wiaK3rYwBHXqlC2ni5mmi4aatAtg
Vx/IY37Dth7Yb6aGKLpKzR+hZ6cy9EQyiJ7jgvCqSMUGMPcX/e34AxsF4w4bvaaw
isATbocDtM6UNbtN9CvUOOBLSPaSZU7s9rwlbe6F1Ovt8eB12xH6n5tfWjNWQgqu
Th6NqHXt9Wx4CmdDYFOqtW8zlgRQci88N36KjaKVEQWzBPJaSo+1jeZH7cc6ecJN
eh0csq7kwEqJ5oymRo/TMlvjSU2Sz+bWCHBGMY5gpftvZh8HwmK/sI1/00kfOmyj
4wslHhiWeUJm8VcgWxMGR25dQcaV9NHAPnvKdde8biSpf9/SYVbvHS2qzf8qukwY
qxQkRfBefD6Rabi3QsKBd4estmgBXP9PK3X2OKJozIFH8rmsw9/cA6gEnF7yq9+p
5/KHNqyLsUwJSDXthoy7nWfc5UbehnDWncuJWkc3LhjDHYagxOVxEVWrKICAkewq
ymQcII+E62E+TEVzJ+lkGWjUpzVXjsJoQUKRI9qL+9Tu61qnQNI2dCKh27PPJgtL
fNpAJuQYQPzIxlJT4YrOmkU2mt5+bSXGWb+PXS453yvK/tSG2HAhMhmn/7Zc34S1
9tikyS8Nv+G5X9tsjb7o3UllxZq1/uK93jQ9CU427S9GVdyCMhWm2xHNxn7g8JEY
jEHflYhlBPsXX5k1Vmif7ByOOm/yi4WN2RW9KrIdiPM0AIi3F6+y5vGcqei3smQq
kDieYlZcUFsVBKf5P58bIEueFtJdX+m8b/Gay8fhmjIWW1mEQCK5Z7NiUJzGFMaL
ZkvH3JQ++Hl+gpXafjfm6QQrZEwPh6o4qVO0R59MBO0OX8rjili8hq/dKxu0vQ1E
ORvLNYVenP7Ck8E8qQmHdkMYh/r9CTCpd3qUw4InzWLjj/V93jA7I/ldFPjQvvlE
m3/zfWokUu4m12gFYpNTY2IHnsR9ynDhK4QEea3PE1vnG3lhH+vzopQiF3B+5b88
CRCUjnxx5sSTMHug1I5KTEtn7npQYnqKvoO3t3xAWMHPiSBCWT8jfJabDUi+iC1/
PtL4XyRtkLiWPd1GeiBsazIsBCm4CmF58xTAWgFRBBI2ucyoCeHS00rizkLszf3R
3hOOMTJ/vSoS0EKPw7E5RQL0ZUxr03mY6hmGRFgbNPqeKL1V2qey8Cvr4kswjN2T
WDeemghWV774aphGYiMANmQRxog0fTmjqsVlCCwMMPTAJga1ZlMf29ZzLlBgD0LK
DPNBw7p7KxBKBjf6/xek5pLzJRJQjtasf4qznE7QNEBNBGFWjNu1iDsUaf7X7oZ9
cEjcFzlMNBtRd1/QTMEywN5gwRsQOn7u3uKZSkDBYyfg9Pe13qa/f/1hbQEiJP2x
/kvygBIeufj4alMqTJMrxydU0mPp32v4cyosN82laR1AkicqPd1KpHNHVe03YesD
bVcumD+eAfdoztzwGYmj7dTZth2c6fCiW0bA34BdP8YK7Nl8YSdFQXrwRytBkeTe
pEsV/sfpk4qewshupT31e0T2Qmvevhl3YZK+RmQs5llvq/Scfi/itEE2qmdQtA5P
1Pe34lh1e3Yea8KQLvzZUiHplnUy0eX8whwQODdzJOh8jXNQVeNu/pJ69zBTK+Pa
yNQjv8Op09/b328JllhJAmTnQDmR/0xXJ7xzPpm5uoCKUJ5yUl7AHKz5X8IPJt0E
4tvzmUZbxxwm0mVA/IN7HyVYBoJlJBRvzusEhCsQDNp5KLWmLQvDnUx9nug7xBCu
lH7CJPUrufPudIvJ8Tu7ZP7qxGdZbx/pY4wJdTQroH/peVf1Aivd9PyyPQ25IG/O
DJsFl9qHmBUlXu6aenJzZSs7ENBKWojGdmDgywR1B7RM6de3Oz9QX37tUxDnbjlX
L/XSUkpybpahPV0RttKLVsPeIaOPAH6FhmHfd3CLGQVey7CSgPVSJRmcS9qwXaHV
puyW2X87opc1+M5ibjaHjNJWUj5iRINb0/IuFpLhwfH4kF8ETxdut7H+ReCJ2tjj
dZvcca8EKAGCgqZsJVisTpnd9xZzyKaE5psz5Ephgh3waSHoKjBMYa4o6GAHP7YQ
gARR4zmyDW5Rq7BE5NhmsW/yO+0mdIwD8r7owqoBDuqFzTaeMXpOzaGw76r2aIT2
EbR8F3YcNrOafy03dBEuA6ilvHHXogZhRMWdKy/9Z5PSest1y9rIKUSXcVKT0Lqp
Gm6VTvgcOC/DYQnVzDQsDw9MXC37DA1SuCDQxw+6kj2c4V8AAjiZbGAEkryvJGbY
TsJxd74gLpY4x6FQ4cGXAh8lwaQQ2R5h2auqb4wW1L5lrk7C3TsNiVWOjkVQWC71
LDPEUNs4ZfV19YkVb+zOhfYoMdC222HWdrqc9od5mdpUpp7UlLGLEvk/o0JxS4Tp
exdFkiEcADxKpSbSyzcjn7ZN4MdEHyzn5cFneuQPWsOOEh2w53NHIfgxHEqfkSiU
zRfxX42mJ5drQZIb9ZV41ZlkM0bhLDr+TyyLkt3e7mhmtetGA6XMC5v+wPhNyeU5
xJoVh3Qot8YDU+kZpbBi1Zma6ugWI73o6xQji/HZe9jFYOirSpHMkRtCcilw7Eut
9U1SVtX2LGsgD1ZC0z7nzRgSeMxjxrH3u3qHCgxcRJ/NLxhKsnCmCqciUGLmspi6
dbrqU3ecV/pu/YbhLxJNW94OjQHAT70FsNEkFpnEWZVwkRKNE00rqIYb9Ant0skn
YwXdpsbGc9CPAwJW3ycxff7gsvy55iyrjt4lKZkz89ijyfUXJBBT5JSuvfAzoWbY
ZX44JJ7Jiw1m9xvEn/8BP5YhPlq97KdPSb5zCjJm00oYDFomLujSzgwtrCES1CSr
BBU1xbE85YSgFQe+6FQ834ym1ADttB3KkzJPadMLVsIc9scLLiXeRv6gzk8w+gb4
495pI7sByZv9LJmX2cUauOeU7XfjKs/n3rVwH6uPFjiwyZfTuy9naZGRSZDZpN9G
zvaWV8VTJsWzPCJKHGaGFfbJhe5P43lofakfX2mkpaO7EIpdxVz+23aLPXFT6mkt
UdR4PQZsWZauFJYU9VYeCtmOcwe1Ve245EExEcEoor/vnn40f9XzxX8xB8rpzGb0
vfvAC7SiyV97gAMtdLWn8EpPmO60AplVbfd5TUn9GeCM1Kk8ySfDIhUZul9QDVro
a2Bd9GjTva9Cwf4o4vNEehvoPAhSxPko97ooSa9ytrcYEeKo4GjbJZAtXs4Aio/T
Zikdez/UNCw7AXnElS9vojuLAV9kzbbx5oTfxxyAX2UsID2oWcJ5nAeeydjX+yjx
c8MULgg4iFNgaA7r+qq/6ixTA4grETi75sXk9qQX88yjzaNycrG7DQE5IrEVkw/N
QXuZjNeqLyzuNylcsJvUqPC6NjP1xfonoODGrDdPJ5A//PkMPb6Nfst4GKRUTlKF
aW/WQ1w3BNjBkHjTZt0ON8yWoj3DFmuIvviSwX+sTPWUOPOAHUpRcY7wDxP70Vjt
jYPT8fve2xzSnyKd03GxWnGiV5sIWL3Hv8Ejm1RwwPXEqlvML3MHypZmgK4omCn0
w8qcr++6gZO36VR2O5BMLd4Z+7xiRipeGEC2BRbxwLHs50K2YTQvxTeq8NFvpgFg
O5C/fJIVzKHpj3CyM4Xa+z8+NDsZQ3NfTvp9EjcWkpZHbW0qAAr073tnQgJzo0cU
6xVbkLacUWBjmF6s3noidxklmSWbOFa6fKIfaHKGzpsz57nTtALFUH8Bx55CIQZQ
bKQdqqsHkcIR2HsirmNik7NmdTK7rkMzyEy25nq7RzcxfiCTfKXpN/mVzBFt/xGh
rHbFunV5WE8dRAdb2bWP1cwF8VAu4NzCVRGYl+iUkPjYQicDXwwILSyhwctq1P0O
pJtE1j6t9VjFj+meT2MKpKexdHcYkzQOApqOuOca/ylucO9IyzgqQDviwUXGIFDm
epom2GvI213GLXmrG8va/AoWKWv5Fe9uhY2TgdO3wSrQzE092V1KKWgWtQRQoz4q
Z/PlkpNYVtSVO/FGyBJA9BPFQsp/rb/j8AcZxXAs2j1YhVxC8UwkBgyH9R8uqIwA
JZdX7L2jrol6vMAQZzvg9hzhMrcVznYzWyuxAvlCttyzrxfcDxvow/DuBzitPcBD
E5VOtjalpkH2EMniuFF1JHiiKNGgh39Eembd/dBL15ZCTKcy3AOya/Ei/FOBPY2T
x9uydzs9s66gKhm9XF1GdsjrBtb3Jc4acKzE2U/6Ostu47gcfhIEWdWVRJZB4s47
/0A71jIkPkX7ycedpuASg5RMGvZSAphhSIXfk6aq5K7VfQwzcNN2QBhTn8oNv3GM
UPszA7IjLdvl/t1l60SJCVMLrs1jFqWy4KPFJkUD6yYD6kzW4UEIAx+22tV7gyE7
/pvcodbAKm7xWDsecTi4obEkA0JsPN2Po8T5GcbFOYlXC6OQ7Ah7GVO11ttDiExg
y29ruLcNwyxYpqXa/l2lKWISHYBqN8ikJD1D8LY432iB1Neg7TFVuXZo0yLfI4gA
idpIcopmOQLIlVpKK1E/r4z0SqaK4IiihPCIqbkxgaAIDsICLyTnELH5GWZiirQq
9s0tyUpwtWsfPWCn7HozJQAJy2DYMAkw7ZXIjuYwA1I4nx8Jape0QS9fWYcporz4
lzpA15tD2BwlOXAuoX/rGZn+DOrliMQecHxRY7sySnvzA28eRonNaSUw2BX5ngjJ
MumLc6GDaOg6XQyQ/X9fS5iW9QasFsCIxPsBPxpwEXCr4wdH7GAyYGq42Pv0exzY
qwflbbkEKYKVqjHQrnfKDuP2oJDliacx5vO2Iwg07eQW3JEx/ZAQ+4vb0PeS9bYR
upcF4wrRD3TEPuFwpRL19x4zEMVVjCn5JAT3/GHGpx1Tk7zz4XjIs/vrE19UNqse
RPhCWlaEfgLOI6bAVdzjW5WzMvDcYke4VabizpeeLfc5T+j8ZxR0MsEIu4OXmzmE
E7UqCmWXF2ZfOYA03zRESzdriQ57P4WPjtAT7KBEs9E52DEG/ctt4ngCWkYzii1R
eURyj9KuKUURCsuEkDfjD7ogoG1ADeXvpc6jk8yO7gmBlyptDrex6XdFGV7EzarH
vbHU7LVC2IfynJYDd2uRduX3REte3PaUrSJqxt+Nxqo751cn+q3eJi4o9DOGTIxf
Rnq46CXE0U7NNa01SeQufwKSQt3WoAYMvDGEGBtup0p41FvHIckz0TdR0OYr66ps
gSM4KjynP+nAq0pO4WOi6OP6kPK9nxN85A0oYgvpQmsgd4ARxQURvAlOpO6dy98Q
9tlHkm3YHC2gkgHDjxuQwDNxRtfmarF0MPVEmyv59nf1P1z+gKOHKFpNdIrhXlty
eHElmO4OE814cqL+F2krMoV6U5uwPG9fgQ1nX2IzcAXNwBeXkHn1XGtVXtObKrCM
lsEMWDW95OTY059srPY8sVu0uu3Geju1MyTCgR/EvZcAzMXEk2k0/Es97rop9tVA
Ln6ZsUtYd1d9ZBT2XHEFXxW9+2BVIoioXOysQEXlPIBDY55ynLgsi5bnH/CMfW2t
LL3Q7FIluRIvG0DrfukCdrAlTrGgv5mU2Oz42XDPtaR6oRZAgrgUt/nMIa9/WYWy
rrQHKXxudCaD6IJnNqbXwkyNwXKwS4TvYQ1Sev7qqhkgA8T9c2gqnYHrP1wxEd8n
9CdMChc8KMASspyoLxQkdDoa7ybhW+uv/gXMYdrhh86fdESsvvixKetadlPPKg65
3dvw/IRrqw74XGhG/1K1vEHb8vyhGvP7wX8qzZRYHAsW3EXrzzwVb4cRG+JGKMvJ
DHf73LRXChrPqwJezxj8DUQD0wSGqZ2NxdvBuSwEhL0KZvD+LfROYdMPkVc0nQ9W
S63+MpUFjx/iPeTnNtMbj68in8Q0F6u5odSxM2aU9LLtfQNq/l9Z+b1tjdiy/k+B
al2yRiQnzVNJw8foJWcL8jfAtxl/y2vJKi9TbqMO+16pjDtySqebEhW6O/2qe++U
kiq6yUomkmAA+TFzqntTv//yWjRDSeJJGGq7ELQYGTPS3Msops8oC6IY6fsQVUQS
aM/zbYucW282BxiOaXX1CHjGCC0EYdJeqTMFouNlZC6xRAYTIkOAZr8oQzhnW4HL
Uc7HzFeEakCDVUGFhjA+oJZj/s7TulnOjni+vTiys4jKSMW8GDNPQI3/rZ9mey0Q
lJYLaZMPm/RP1jNdPuUCS3Yl6qpjgdnMNArC55uYEnvCC8g00kJrEWU7f9AzG1eo
GfyrYCfszApsyGG5Tgh5vm9GybyTDYeCcDvd9GHi2C/F6D3T80+oWjTtPSYlLu3U
yBRXySYn0qCRDLkI4zwCBhwD83RgTI42aKZyNon4wiAexb4AMEF1A44nj7FArE4m
OlMc2KKHf6zpP+stzO5eMnr/q2Zh/0w96UfqWnl2SzkAyGmrBj7WY/XIfWh/wruO
IlOeK5lM+96CVUw6+7DDyErSQqJA/aKC8HFrKwg7cH0ug15pA3Bgd0hu1jN+tc8L
CywWjQPA3bJwELgnUTpcfibMd/bKHn5xP/qOhV8Nf1qdOhoKT6TblJFgA/1pgXXf
23FNUHrY4NMwUwhihPv5U2akvk50Kcmt+qfTTJJeVUWoYpkh/QpAT6dwL9o3mglM
nCVs/bXaCSoLUlQvlz1pmWjgqCovNZOggD7z1wyT7IQYDax4WWLnhQzPk7HUxkub
4kE7fgXe39XtBmBoXZ+zJbFI87Ur2COx0JhJKFqjKleGStCg9S18bdedlALw3sB8
lxxDpa3LgYHuzjGaMxGD/T9Cav79Qgj/NQFri2S+9rz83MMLwMXMbEX4AdMQJosF
/NDFfhiudVsko3sGfTCukh5VU5LLm0lC7co3gyJEnuJOB5wZrW+uVBHm39f2JbSI
y3oLu1GN3nSyzBhwPX8ZIi2EXEzvAapLWoyd9olMQHcloMFiCX11IU5uUlZRwRpM
8cr8P2NM/9NdsbdhWqt5QF0sspgO+k3b/5nO3NsGqjOeGx31KCK7Y8kOJJQ0vdBL
fWv4/s/6SjdY1AsyL8nFDCVCyFcVtJY1my4zP04/pxOdDeb7DHGp/1AZSB5zCXHl
wBKrOeA8o7IHaZVNjtrpyJcV+QfTeh9HpAZV72EKB6b/KxUfAW5peNxvTrl8aJZ3
ERMlxyrF3CMjc8lSMwcvcH0yftXUH1tUUmDl49CNScJx5EXThzWodyvTW8GB9a28
oRZ331PhJYROrp3HVefz8MqRqtDcqkAAohjuhFDnjNbYDBBWaXG3RZyRCM7E/2Pt
PGqK54heEXrrolnquwaga3tJBGVrzQYt32UwKiSNjtzmjKkYhHtEpHZS/TCDr04U
7CZLQzDuG4tlNAaVOyNqcQv2hv5EzGsc9beWPpAUiKyg+3nFh7n5/E0+QuJbMDt0
CW100Hxl8iD4oaIqbC+OY3lTFG85ZmXtg94w2ST2wB0MH9t4UcMRFJdQYiY/5oNI
kNYfCsHZU0LWPlOl2lfQ2fyAWqAGB4mI9syq0hA+gDQHc2K5HILe83Mf6ma5wdVE
aFqeTp6GRw7be3aIIWdhu5UqxoMEtweAGW55GJwtQ8tfIJdRnoHX7tS/9SiD8txr
la37fSjoFD7iPwLQZs82jaMfBu/S7NbpJjbIAsDavOYtIMnqwzBp2iajFmXzR5nU
Tv+TSyjqYOrMFkuyV6Ex9/HuWQMbQpAYeuZvjtW/ubahD3ux8KB6r69dSPI4RCdj
3SKkqYFmpSsYKS9gzfS4u/KJcUgz+rJL0fBmOWn1xhUJ3/nJaiUcUQOk5wwto8Bv
Qi9faMiM/CpspSe4IdJZ0v6pVfRekkrpL5R8rIHbhhae8Q7foBNaGAeNBWjITV2j
Xro3IPu4aRSjjFCYZNWVL/ARPKbnZQn8Wdu1oKIQ/DMg90BSK8w014rCIdHH5lNF
j+r1FFveSZksBi9L5h0s8Me5+HsRwWsDs8S+Z0RBrMQZPdi1YMajc0a1Ioa/V7De
BCJirTmKVKVz33lokZR3FF6AxZ9SjteBdgOd+99DpCKUFOuNVYsfZ8zwqhAhjMvy
Mtbxd0bZEp/fPJBF4O4WL3Lh49ZG2nX+FAGWoh1A2dLKjlCz2QUF2ZdANT6k+6Cj
A1xu9qZ5tIkCYYU/iV1rFw14o39Qkwj6GQiyM+fkqwWhvIw2McBKMAJRy/Yv9NJi
T7zqCqgsWERgMd/RAZBNFyrrnsAyoDqfUZp07uswtzhFcWTwBPJaYnqI6MlIy61X
nAq/npjwTtvfY201WQDlZip1iNqFbv5i57+psm/eD6DxdzdSSYBl7ME2w1DZz0Mh
5Mv0DowoF0h2/oe6vsUbUghi8IZiK5JXTbN5Lhy0eHtpqDhQ10FwozwvIfXI/1f/
7IuI3xgwIplpV5V4+qH8KTzKoyg9VqS7+cl5HdBFc3jvOnX7kDWKqBwTypXD4HHh
UmEL16IoIL7nO9UFKGJ1Wp0majJbIO5r+Q6d4AKy12QeDJZtk9gDGrNNkxvUySYb
jc/sB8MmoM+2KXwu5dmw3LBVIbMoL+iYtpOERNKxR0aDZoWKp6LPVZiyTW2lTfYJ
WwXUJ6TdJXam+ZNfgLPq6gpwijOBNnXFFvgb17sSgtP5FK3zC/j2fMMpJEf1bof2
zGFD7iVIu3Emfkh53Ac8Ev76R7dIQ8AGZowRZzePlRHN0OusWic7OxD1Jm6Ow2jc
NSEwFmu5+Rnf7QSsnXk/P5fXKqrEXutJXs8YLSBDUQkRkJaMqhBUsEKWxoH+MNrX
9ieqzNXxdWBdc0iHM+X93NttnPFgoz4vNRlx7T563a9xpwB6F8tJ4lrAFF6Ku3pE
wj+vD9JHMc0plvwthhJyVie88X9Edb9R35BA9FVqLVtIDsXrbQyX9TEt7qYYiNnZ
3YSt1Ule1F8XxseYQuIg6HWHub8U0NjMyC2Ehd64Hpc+Yq/sdj5I24KhwGqlhMwr
Z5LdfXF1EKjn2wX0vch/Nq7GF62RIw4BqpINQpTVbZ9JsCtwY9FHIxg6DIKerE0q
S+1wn5oNPxpGRyBWh4YegMaGlI7pG6cuvLQna4Yd0NoHAXIu/8I0Miw6kqPOXPQf
3Mm2LhF+zJkUuTPzTwALq5Q8qevwsj5M7/WaRcssZg1KdaRWiBAlVOWpfLszZs77
wfrCE3wUWeCnBkeX4Le6+6mYIve1CjhUpIInBAcAn/oDIVh7wpkwwfovQhFtg+6u
+r1Ac4KE1U9c8PaLVn539pFO9I60KKqFnVgrGh9/CR6qLhNmkHQYRzlahP88bqdc
H7LNiJjbWK0QCEpI6b57ozj1MDiDZgHONZw/c/WqMCBvHZwr+MdlgazZKZG9Qvpa
V5v6DRV2orTq68zt0DWRmpI9RYZQMJ4fzBDn8LgDxvKoLea/C/RS0KBm3KOZWMOk
WNA5uXpYjcQekn035WY/nbG629is/RtUuSIkFMWuUkT0NmRrgYYkj1rIvfsK035o
fkZ4GcOx/b7B2tTl5TjUozQh0OvI6ih2CHrvlvWrF7tiEJcRK1DrPtFPW8pZqCtQ
KQ4rGXHsxqxrJQB39RJxkm0q8zXBHa9ExFStbLZVDuz+pGheewl0piFv+q8F72iO
tT1St3SaLTAQ6JEzB31cQlmL+adCTioOxXcuCg+nrLSSRVkvyBTf0NZ8ROMxuI5J
OI9Ex1PPLX+Dc6z5IlUneWuago/X0KxqJ7E8J/L4a70/nPzkqvBS1qXrWnJN2SmT
U51inu5zuUCuldjwCP54X/eF4rzzWzWdnJgqWo/BegLyYk9nmPkNV+JOnyw3m15L
82jIbo48uoepXfkESWe/ArUQ+o7Ja4k+wjU6KBGWpjAP77dXOIS4QuJ3ENrn9sMQ
CUkOGMJoJM8V0xCP7BHKkHL6HfWakpQua6TEh/I+IjAJ7FtcxLyZpsp3SFdEK6T0
AV4bZ8eZ/rUuwxlV/RUJppmsBF54hmk1KB6N7NI6+DEZQmF1zA/WicZjHZlIhd/B
n0t/Hiy4YZkN5bq4NpOMVJCChzp64xE9an3kZU+2lxuYdKiVEExMs7taXkOFUyZ+
5052Cc2sSm9aXMyLUJ/st4hAoYR8DDIu63uceR5P5ZHgJy+D+w/JCFlqo6srogq3
KWJwgCICB1ruZmbyJdxtnqGRtvGc5ooyzR2BYOaiLfqqw1m+Rf9wjGsEEtTQLwwu
trRmSpCQwvroqviuVSG5YKXEJxWtLBusrFV8eXnfwt0Qr4rnWTO2RiMy6yQN35xX
rnMnnNFIYlI7c0L7bG6Uj2OP6C9hceLdpHD9Z5JEkfyw1uCnuFdLcyf3YUacU4GW
ChoPdeiQkzaXMVZu21jnB0175IYQxtthiAn+SNJWVlpiWYFgOC3m8d1fgnhG+NYp
w3msTrYOq8XlCkc9eC9iDpeeRrpjFFJY4rfZRd5/rQKtw2E6Ph5FH6aEEROjdJ7Y
IgwGIRl7bsqrlctrU7pn/vSz5lKJmXJCALFDoFNB0anR1lwM/pCaO0h9VtRiz+6F
n0ogt8vwnVQlumn2/gRRV9RMJ3PXmMMeS1mVMARy09j9OZDJOc5rG0wECQP///eY
ad8avuFAmdHUddO/wSLlaI8DTuXlR/wmEtX6LeVdxCbw7wNSEkC616/9k+/rQN+f
ZwaJF4bLvDhy7Zq/D/tzbDSAg8XbD1lH4C6Yp9kv+cUhjYxfapVQQ4yOatvLm7pU
zlwWNapV8tOysGBFRXTcXWic003BC9YsYK/M7YkUzVfEMmI4nC6L2kZQaouua+mi
jjw9Uk4Ag0ekja4ECvNLl7CO+6a4yII40Ynx1hnARlyhLG5wfmdhtOd6YvzXbC6t
62iIqQBmTD09uXRxYqEy4pBy63aiV3DzkI65O8YFFbwRVYOqGoiDgIPKsDWlJY/s
JuNeOSjkrJxgte86/VNygObaj4QrhOCiM5BE9m/54+mqIV945YyEX1xJgHMoXrbD
flJRQcGjPmdQsCFajcJuI2TzOPHE/dRD7Ujl+YgvQFMQDcA6TR0PcyqL7arCSN2J
ec8cKOYD+xcB+Ht5vd3Xjtt4GV23TdSssSUurCSwUxQds1X6RFbNH947CpvlP0eN
V9TstkwlP5XqMwnRKAcY2vz2MGrMokHBbxU2Ffd9QERo36XSRHcxKB5BQdvZVEOX
6QWH7W0VdldpE6Q+DPBqgfRXA1de+7dagXwTc9g/eX0becQUxd6BGJkhchmWIm7k
syYEG0brOlcpJKYDY+eKZ6rAZ9zzwUSwVMogbGXjDp7yoqdmijJ396PNgbG+GVFb
dvVz/7hUPBtYOx3SiFr/QR86h3BlQb3nlHEfnW/lJ1Sy9OMsGsP6/Po7i9C+evn2
RlVCd6IJhN3gRwfEXPivI9VIku9Tx5DpdUvbMCN1g5xm5jVQxZL06fg4bW6a/XMt
gegIVkMEi54QMH7Iz57U94rVu4HcQj4dkLIbdnoXapwiwETdqBV7XaoHRecv0Xbk
zGKK3p78HelZdTYGIHWOT9cr6RECrw59CmjmTOuA1ToBXrCUp1dq5DcRam+Q9bbv
4J3maefHveCKOat/9rdJXweI9t8AinnDHHxk6wWrIq0LUkRuNp+U3JBpn14GL6QS
ZUZc5edTbjINIXN5M59sd5KslkQWjqhkGkLLicq7bN4GZXOSaYrp3Tug8uACYthJ
oP/KVSdxgTYYj8TZ0pGkStt5v4XXOuU9LagqFkFtVTDOApF5MIIqtGA/EcOgc1LJ
ZfJXGe1vakej/nx4ETndTlwOb2h4+2HfgLljuNOIclXUK8SpU6FqXKYkmiAtsGSj
a5/k0sV5icnEt0RkWJWrnm9+5jZw7IQMAz0lP/tE80nFXpcJAlyAL7nZzVuCSizl
38nIf0HZ2MeJJsZlx9M0bV8l8BYspOJ+nbMX+db6cPWpUGfmZ8w60iiCvkGVufAV
p5J0kfk8mPwogvVAO1PAPdcnWqbaDx5mULmax67VPoXYVyQIf9nCq4z0FTyRpQBt
8wn5UyT8ZVuXhrcvLZhG/iUAdYPdSmOYODEgstrl7uCV+pt8UAGNrvQ0IzI5YLDt
/8lyYN9+jx/46yPU4FV5TQbcix2nIYGfAFCvAyLp6gR6x37sVMldksDf8UNRft7U
rgnCM/fZ1e/eaOgw8oqmtYTBkyvun1OpkVQPK1/KSP+oBZ+ontCse4hkpn4Pxa5/
qbbeYXnzXZ1ZN3JXX7EFlawGuNKVDsa/drzToNSibnd36yhAbtfBki0GcCzKHEDd
D/KDQRwR+Ty4V+KHymNBoXjkWTueg4KER6hpif6Wu737tUUk14SPXClV3wtHlsAx
9+3rMv3tSwHt3soAASWHrVuHGjmXsxHnYRAR4bJyJQjUuZtVkYCNBE2lI3VU4UkN
M6K9B0jAzsH9aLPhaMcD7qMTMHQR2aoFWFXsYAzP6FD2jx66DwVGySFtlJwmrIef
Gx01JBsR2/Puk36XdRxJLbQjIFgNtDRLx2iQOEvj7kR4+EfyL2u7Kuc00hiV/RnW
iJuOyf0s/Nn/2QsDZsnxL8BYPl7W++7ORjcDhjOu80pw41jLtjABCRPyVH0PIoxK
cVAAVPxtU5zXqnVI2J9OIuLhhpsDRlrbV/6B4Lew6WW/fo96QA7vjVkyn96W2XEC
JHfTXaLNlk4QXruJMHKe2ORUedonLTtf068mqLbeEdp/sQJeCWP13IZtrpkCptiL
BfZHyTEq70NZsBQD7xXpsHNNHbMlwJdO98d4K1hr5UF/TKHqcxre6FhtQYQ5+2RK
lmmQwDe7svFy+to/v1q8YiAgWSD0EZlBUuEtLMxf3RrSOd9XOzc8fKT1qjlmsPLn
dgW5dzrcEhDmVdwxkG22H4bcC2hcI2Lx2o78RswOXvvVMdMVMM8qV2VDe91a3aaG
TU8qWH8+o69bQJr0Y5RNDbAT1pL/fYId6AF6xViUZRvUfvyaW6KYCqgUDgLgZ4ea
x5ttk6XpQrBzL3mfX1VYcId8CGys/q+05Ayc1X2cJWh6hlY52sueW/471CECm5Eo
HypXjRTm8xjoI2y2gp6O3KTtavYI8eshb0Bk5zuDAwy8Pc3+3Q/MgMXH8XQkzXh4
NHd8JGQ1x0UOKk1YntWNLtRVRHxMf7lOJejpV5su7ze+9nrUkY7AsHk+xQNOkspx
PzGPqoJrn0oejWrT7wCGjyGq+20uDJNP+esOtL31rsEbRk/40z8SsurJPQ3hdjVb
QgAJkB+1lQGuymnYOZl3ZebcPdx2lAUBZaqadVulLJie3RqcT5edDTy02Y5+6nFc
iibk1ggW1K/+Rt39JGto9Wu+Fp4lK5ArXltlsMQ7HNDvqZIVGr3Uv/6UljN6JAZd
pNZXfr3NYLpEaEc/T06ZlJAfpK6UOauwM6eQ8UzsSdNY1jMNpO/XLlaO1DinTeG1
JfubtgVd6C1ra2IJuxkeyhThhGUT+Le2OlqNgMzIENcHIzBoFpaL7inAS8TWUYf1
wEAIle1jjvPZCIlTOwN2lgyW2tngkDJktV0ynXq1hRAcQtfXYKnzSg69UZi8wcJs
L0hc+s68kpmT2VUIO5wj6jx//yigqBwKssTAioBrEepEujCZt3EfMO5x9mdHQ/8x
7lY/gC36Q1k+23PIi9WPCKoFTc4wgVV7DjiBtUB7uxvuEtqDUVJjTHW2qzLqASKU
Snihitu8svxBfp2LblHc2/1H+1ca/JKTdpqWu3L2XWts6W4G/pJTJoDTrjROSmm+
7wEmV3NJ/oS+gD5iwGKPXXpb/yWgkqI3sT5gdQRmdrzLQ8lJc9vrgYqKWd2lyp9y
URypM5o6NlJeI7AJsL/+wIFBMfg9S3c3ZyPtYJPiNod6B6t7hMlYekotTye7rY5P
3oYFyB5MBZ4yBXGgvK6i8tF6dfPJC6qmR+Wkgw9DeSDruYPrkGX2szTxv7HnGXhd
6pyXHakMtG8eqz9ej2XbxGYHMyuNC5esp0yXxYHbJsfyIN+GqO5zrFLzJje2/sLr
z72Tu+UvtKtRRZ6vPR5YZUiEq410jnYu4/1STVzjvkVpd7N5RYB7qQwam6KvvcyA
Kkcy+GLkm2gUSlw06Voa25mcdZGhDZ4IGokkzXpoMt4fGpDY9Hv0kytF3XRcRkd2
SbDsCq+ADcsFMwS1X8+nlBrB7OkliaZkynKwV/wtuKyJ4PA04dEkgt+IjN23/xIc
ScoupxyQWHc9G9yjMqyYOzHBRFhO4TdxeTTQJk2/29/e3F5OBQpud8K7kKWAiRAh
6/LAItnP0XZF0Ady3qk2p0oEwC8MBQKDctuaPGgAW5QISQ/7jiCEYBnoeyvcN3+u
zZDfPd3Krqa4AudqrQ3Ebj604rK4F/8NsZ5dHeoouELzNeL7hLmE0WFpNsZzlf4x
WFDU9N/bnybZFyI560k+S3bUlX1tPunH2Hp15NoHV+In0TKRUFU48wD4zH4RaD8z
+o4DyvAubqQARQVwAUbh7i+YLX71CcINpDjfQpCHCYRH/NzV1Yg9ePMnz6wQrUGF
ltYnL/ezuxBxRbdHvfQGS6DVB3pDsQbFtlSTH971GI2uelnOEn+r8ka9RT3eX/Kl
rHJDWfWdOj25a/eix9QEWyBGI6qIv6pSLTyuH04CoJ5HPtvPKTIfk/ynmbEjm/Px
ct0spwKBYiaGhzoMxEIocxColmYJ/lsxhMfuG5i+ZhtajrA2/9UXGm0bSKIf665+
vRiPKankOKIEry6Ie6B5LgHFrBFUCyqASx9o/kffSLjXrbdmwW9jwzuSvC+kCyT7
YT5ftbx0WEeofiaWjO5zfycnxdtoxr451H3UEEz5OVND+gVBCW+5EZcDBPLUld1A
6selONzqilCVsTNjcr6dQgUTXaAEfxE//eS3yTGEV+NHjAycBmfXoumfvt1f84Sl
ePEGuM+uijQhY0Y2dFczqky77WVDZewMMkHXtIG/UV8Gfse3OhDzxUsz2gqQ0qjF
ElFycA4oa5IrBZ6CfW0Ui2GJmb/mYnjjYYFqs9joUD0zgiKCW2mE3KM8Ecug7kdk
8nZR5Cdme0O/y8Z0kEs9E4K7maK6WVZENSiz9o9ekF4p5tfDmo9COnkx8flf5OqJ
Gpo+XDE3ANqpkajWkLES15Cglcid0PCFb1LjQPGcGwrG3oKHHq3prs7qV52OpEMb
+CEC/a7q3ifTdGuFgVTdm1ugpVfjNJG7BFGLIn71in5Sw65+vMoZ/IP1AflwTd9J
qLtZPZwltWlKxelJKTzHj0PqE66ufQ63aXjKbF5Cyudn/fhtxN7HufSKxLZlcvHo
Z/1tQooBi00rECkI0A9C/UbodIMNPoeMk8yy9cbON9EQGlh9JDhM7MK4jhTeePRb
kLrd2V22wzIoOnt7yWXCj39jsqLVfgmJNvjj+AG0o7odtg5dd+pFpHNr++Kktni2
yHAOTNwEbzmf6f+T00Oa4QQ1ORaMN4jq3lg6hLuhb7CWmBBUS244Pxrquy35BPSN
jjnhIp+Ca6tDoPyAsY3763F7z4zrvKp+21Umc99w8MKy4HCYiMpt40XKeRxcAfxX
Udxt3NnFbq6j5UqIndRVz6AlBks61hySMHb+DMOyyZ6koJgLuFtgy/RT8uoLtYVO
iKW1V+kyImzIxXu1mFbrL8fueV6tsfipcD4NHORcOVymWXMrplOqFeACegTXEJyB
3IC1WC6mgRnYOJ7BbYbjMYOL/ToOx0oD4MGOqmgGJYt5wUDFF/qJRIbERwX8bZlS
vrXYHieyaZ8DfmyhDIanXDR5Qp4kRsS+Cbt7WQ91EPZ6/20EPwOOZ70V9BM2lmca
Vu4VGlLN9XDHc1OTDwNdI7o9V8SBM2Cyrsf+ip4+Hn4jvW6TX8QGZm/mG3cSOnuk
tcW/pi8e7Xq/k7LnEx0Wnwxyhc0BPqWWa++5fLcWDvku3WiF+nrC3kzk/8E13Whw
x+iCDGSLufQTCHrdnstV3tDErWbqCMSl0+E3qaFYoWgIvBxQFk3tDTdsFe2KD3Zg
veIv1vHc24h2iTlyGRCN1096cXvxo7puVaKWq9mrckpYc6eWf8uLKAHtD1zGVFTs
oEYSH/OLL/dZD60VAldRd/S654duMf+nbx/M7wc/sNQwkCnQlLcPE24quYUp8Q7F
hF/y7fwL5C5FlAGyexN7p7htKyFyP//rWSQTQwlVH0JdZ96NgdGhdK0rv9QaEoCT
vKX/tO8X6kyKg4ikhdQWG4a80Vxn68DFhdltmbtrq3/JKzk3ifxKzar2o8bfIx15
1ri3iUeU1EOahRzLGn8cDZCKgYRacdUzB+uSpEIxwOsqkDvw2xsfUAjgcrTYIXhJ
iWmeNy6QsftksurRq53NMI5Jfb+GPQKPxhogroJtmHpcGyVG/HOxRNeEBy1DFPZZ
ioeNRdQqGnImdEr65V6QVowGtS1jSvydDLfesIl8mIDi+tDQNZcHmTXCXMaJwBHZ
XMsCVlrVuPY4KzSFbwIVubjuC2wsvnA/IJYWGSagss6aJ6qKyniuCcyzU3WEzbcY
X6x8C2hjQ95mzclcwM95PvXNeJdk7zK1zVwX4u+tqyP1AtWF0B4Tz6flizhNLCT0
i2W6B5pDQYlqvMSN7arzXTSQXbvw0wUWGwrV0oG4PDIQ4JPjKwj8NtPMlNNe8Emq
l4U0zsm03UQjw8czOjp2EKa58CgiYLDM11/SkJ+LooDQdWHQz4o/+yKPmpyWdclV
QRtPjW7Z0lWvrmOxmWVhCodqXv7kP9A48FsFvxWmr2aKj7PJfcoh3+ebXNXIgWZZ
1Qgm3Zl9Si/Wj9LSccq6p7FaMPF028/A+VMUFpShh4UzQqQ1sB9+IlmNFj9yFKPu
Tz7gbpGaGDJGKdBgNONWgDWQXdYqEJJLnXDD/WdAR8gsbU/xNavD4TLD3eBbzJ8L
/BgMOFSbVByqC2G/Sqc5ctohU9Mg+Ww4KegAjfGIW/bGVQ5chiDPLIHjksMkO68i
hPZ+M+EptD7+vRd+XdPEPqF0a3Api8EhCzFj0rxHjjKXu5eXc2oScPw8RiUqLUKv
KKct7ip7CQx8qjUL79JZ24QF/6ZIWf2A4O/lO1BI2kw2VL1HPBBOJBPIXR1as4X9
jfOF4yZRfZBMseyJ7zBt9wda09N8MR1hyptPInAgaH1zIsBuJBXIt7pMUnwD5RYv
IXjBRIBaXu4yMef1dFaj5k8B4m3LGtJW2oJyxVQTXY8JLBg8Dme4ZIjYOjgiuL2m
M81WEl3ZigNsgbk1Zwr58cqgSPaP+XhWHQY1JpE7c7gc9zN6Q18cbTjoWxtLOKy5
ysDbIpPf63TFO6LomR+WVBCGZ9SQylr5Q33gZcxYR4MlKquT05PcwA/wqbck7b+f
UA97QhybUDBJeZ9E3UUY4FVyOaZ/kROJcFjXCUW8zj1phi5LItYpcyL7ID0Au1Ib
obTorB2nIjlA5fwbZ79H+ayzpCB+7h1nIiVND6jL+P+OXmiNJC3ImMhtixbGayxL
IuLhglcAYpIaKXqaTU7pCHc7VpQgNubiLqZYcLOoAuqVeTKv0P7djVcIAgMt1x76
DA0CqrOs26WRR0aqwYEuAaee/1uiA3K4a43uW8exFR/IQj+I4jeytboZzX9Dz6aI
7xX8z/E6hYmtIG44Vat+t4TxWQ6xLv2VjFDVICb086rFtti00m3skxzOTQi956xD
QzHxcHUNaRlur8wzJrlJE/65dKECbMjOh8GCqzEtENCMy9tQb6F9/zrATvd73J3F
NT1O4UJSh58YOlBGq9iNzJLnnSA4NAgZbZoOifCLkMYQ4UGqfTNvtXdxcDDDv37B
6rUqlzWZ/gDAII3I1nNJbqYMzNOs3ztIEwELbh/llJIRqy74ipm0sLP9M6RUroGk
x8Auvr+dF0MxR9EQ/HJQMQ7VExhZki0WcJVvJ7LHf15htkL7MvYrbGfybSMNFYSM
eALYoRcS6pE1PzXJg+tOZuxmUMLnAkh+k4Y9LQgKm1KoTeUFru/DGn2NRP6+kiXn
vX828NahvefP8L7gMhXsUeA8UbmmjpR7YPADDOe0FHK0og7UMMHLyJnBy2xNzlf5
mj8+iw0SDuoeq76qQYbhrhBlPAnAD2QxXvu/RjIaC+wi+2+AQVHWqqqB7Wxt6lv0
lSUZ8RnlWZWcP/CToF36MlW4eDGPOz9nv3Xa382gQmEspPWUhIMy+SW26dmJR9Kx
tMdYk77iowp+OfQ1N1MANP8Vbq2xoU1/Hx4sQPxg4axfY0HhPa4DneLenZzq06yD
K6HJk1u5MR4U+tjpmCc1LV4NDhKseT6NDJ/f1C6ADx4+hag3mUzq6UbVvSwob6iV
Dk5jjrkt3Wcj3+9Ly1aB8ax3l4NJJHblOm0/2rz0E2AmYpcBk4HLkbuH+llTmYPJ
GJVa/RHBdoWHFvYOpjOfvDv9gUbDLdxnk/71naoawKe1wkBGTd0iAqAvLREYqY6K
l5oGkB4W1ej9OBSURGEn2TEADjWXioym7+UpBl4KDtS3ucLFm0fNEBGXxe/f2xmi
5qngHSUS0bhvqH9UDnkvfRvM/gVK0h20V41sdLY+bt9JEcjvVRdjUSFkiNgo5E1f
xEVS1a4QrLhz0JsBCgq+JilSyiM6Hi0OgToGxcESPw5F32qASzCcv4D73enHCPk0
Eifg17y/UykOq7gQRyLskOcY+hwFp9f15X1uupFAAZfcDTTOgQyFn3PpNvNfJGha
OtbkKYGTpsbRYWieHkX5/j9e7b1p9SgpaxyCQ4w/YL8VSrcs2CyjyDEKeyyvU8gm
0Tg2v/jA6YON2Z4g+QKxNSS9WthImFFnIkpXnpV+QEOZb2ZlLdrdLQ9MG/C6wb9H
9FUiYHIGSecFNjVLTzA6dXLVf5FZ0L2Uk1agFctagw4CNgxhjcEXUiLbW9/G6BGg
k09lLgMdPfxB4ARpdRmsNKs9ntAtj00WfYqJzdpP4AHjCXgOElLEbNvYWeDcZgfK
qoBU/oG6qlT1cVV8d7u4nryEyg5yZ/sRqokHhIJjDv9GLoo1FE4IcOtG09rOEa/P
hRsLMFDGu+5IYHsbzPoFpntsSd7X1xhkhI1WN9U1MJqtzYtYYO93rw5ldDDDX8lY
9OWcko9cFxAa7K1vihm1SoVY85UZbo38wHzLHs+EHCJziamgg3IjLpnYsdvGcal/
mTxn5U9rsk/TZZczVbw2BEe82q+2JTtRbOIxiemcTkZR4keCCQc5CJDJOxHpN31G
zEKLIBnDuZXNDHz/YFzpyHlMuOxXqO3qD03Tu/a8iwjSxyLzuOhBSX0P1WswUVXG
ThLJUdrBNJ+z0OpIOBUY3okAzWmxARlV75rC22DflgGF+QuZWf6vI0gXgA4f7K1o
Uy/4DaTrwglc92OrAFTsv3iXfaBI381mV1gf/JLdzL/iDlHB/3qgUOZG+jIDY2Cu
sWWpjWb+5dozSmr/2rJdZdBZmMjTpzL/RfhyChdsa7i6koP11Rj1jMRqEfDJypzl
K8SBBWKNUrjDWeoRxF6lZBqf3nfrbg/EU+9/Z0rZ+pPBsr4T+qbw+iJq2fr+6vPv
7F/H8d36EM7bR4ll/xgu+TfOuzwMYjMc4gRaebnSg/+5HK6pVYaqz7sthhuuPvhA
te+NUlQkCSfAOKHg70gVD4wyd1HSV2/YvfJDNHu1tmWWL+wWH5FK4KTrOSHJ5vft
SH0SmSOvfZ+O7KSxP1Z7VjQccS9QosXoNWfsWoPoOu2pvLO8S0CBtiNUsPYD6ukk
4sb6bCprzprftmdNTU9jntw5oCj3i5OzWQVB/D3sPVHt9bmMLwleZNjgTdu4HMhp
tUsTw6c2sampOyrK+3b7FCtXFmH3MvouTl3aNXMyosL8axlnBWI823iLwsn8EWkg
J9ACMg3XKq6Bxpp1ubQGpET8RbNyG4X8WChthp/B8V9reK2P654YgToJAgUtzf7M
VSeQXJq8dkweNCrHG/5hhjPFC+0LnfwSqY6X/1NdQSzuE4rL9zM0gapIw/uCUk1U
+Uk8zx1gMNDeCVgaNKNUoaS8PuN/cS+zDo1Gysa6hW+XJOIzMcCfMghxfoqpJavh
cHVmwzdX1wh4Q0/JU+TO8PALnKquzXyV5hWk0D1Kn+k3w3xVJUXd1Zh0GG+Uk5oq
GKpeYw5wXqf11fYItDL7RH2lxh/qmSUjHOv55FV1KkdEMhCK8xNkFomg5il2BHPy
3xQrjuJYdtJM6ODsQqzBC3jsDSZ43O5GUWab6vhkFz1w2Hzyez/W5udBx5n5t/jY
+tWO2RMRGx2fmozcReAS244RVt35Jp/Pvl1PgQHJztRlXTeZsiBVNS80Dtj156Sk
LijzLGSnNoT0B9WvTDJwj01kLX28tC3DIplpPeTnVENGAUMmzrgne1+3f/l9SDEv
MT1ZMFPab8VjGCZqGqJaLmG105hCMKzGt888zHI5NGVIxvieMZweZe2psQP12cgo
piv99y1ooptk0WEazdXm5LZ2DmvjTa3G3yh4z9mir9uqDg7xx6MSPIn99OT2GJtO
W+9Ru6FTWKZMI1sQdPz1OgoJCVqRnCxCfZXLDKbD/Zn85MVaxUVkOKT5EBPA1EHr
n3jxsQt9aoT3Gm4BIkWpE8Z0FjkhIealyjOHmyLD2tBUC+DLV8ovlj+h8l9KQnvX
BKhZ/2VKswZDxhaoq5daXJtrgc/uAqbOEBFe7SSoldOk3cnkIyYs0pnObyN/R54V
IRfZDMzV/HDjMp6zPfJ0oClTKrJhdZhQWn9UgyIGp60Gq5Zv/1RhzVwJcoZXNfI2
QLgUVrMDSD7tJ67HVlsV8o4Xp3BYgnl2FMA+cQttX1lPd3SiCZA9aVzqXWrmmsUd
X48p9nsZkMYl+ujqFKt/duFlkERcdtA24omgbV9mBNiFLc7fD7sA7VN9uLQyUcwj
18Gza5vC7emqDKU7IuO6EnSlrUL4WAphGZb+s2A9vSNFB+MwkcHzAROM5MRs145p
IJVe8M5CICed+fI95zqbu7cblG5d8h4HzYmOpFQUbfvc4ZqV1rK/EX5lMtdGqmXn
83bFWeLjzWuHAar9d93tYEXRVlKTIwyrKjWSGt4bVMXKt4PgoMViFhIb7xgTAYjm
0HMKRjG64ZbypKF8qWcvDrtS0gaWd+9mn5byuaxqIuqWRYFaCoMNFKioMhaBkZte
xUetNeNWZ9IdGkRfQViHEWsxwa9JFTkJvmZvnCwaGy5O5mEE919xjH7D2Tszj7vj
2epAEhxFrKwLAqW/hAQFMS9rRP71wBh2b094c4/aTg8YZS/BXuzXu9qYyTdR7G/A
bFu+RNUlyLiK+omuhr7OwWc66sJlLbPN5hjfBa4Yg4qMgkVdV+NoHhduHji0pwnh
7qsHnRcQaWA3OKxnKzU1JxOrQzanIl3yHQM3eYrajECMawEJ5/JlyCFsyUUfxJsw
RMxkFhL52nIoX4BYhQIW8+lvcZ0sec5NbtGpfjCJRgIzakHMhsk3OfDyzODEeQHv
uey//cjg6wbFH2Wp/skUmsxCk0E0teOz36+me+8hZxsiaMfZ4ZuLrksRsdWKXQnI
sinEZasb9r9FqI2O/RstpCBdVWdXsP/DFiMLdiCTCvl/pyESvkZ2tIOxPTkRuRwR
k+I6yUxiCMIsVcroWtVQJku7vN64hZ77xc0MLTviEEyTdL+6yLlhRUA9h1rXgITw
Wzut7LVdTRDZWFXx2YpRiX5+KiyIv9xLmGpD6KeLgO8CaCcxTk+S4xCpRyc5S+yJ
dUGS1K9e4LV1E6jWD6kg9gBGvoTTs466J/zahL21GbHcaSW2DVAn+zrDyKN2q7eb
t4Cr34G2fk/Z+5t1IIA3ZQUR9M80Ng8KuQNZ4coO0dKKY18pib8U33owAe7i9TS7
aq1T3B30Q7FQaza1nk5tl/1GxLZVFl3JFn17c4KOM/5bChuSO8f94qXiWEceqruX
HNMWds1SQca+5vA+zEP1YYJ0VZbZL4Pr3xtyqt6jlL2RhCFdp0gL3W5U/QPpTsjD
tC3+EVxUtmJsqCn6mG1536d3OkcyauBHYOWS+bhgRW1wWJxLE1CKwXO8g2Ojjrji
TvIKT1M/Emwo0V9w/TVYDemxxFlFVxhbYwny+vKoKnxIp+cMIlsYSDFLLiiJS54N
oZQX13ySgQu+5vbLTsNDK7ud+dLKzbvBVSe9kXba2b5o4/6u/j0H36u4oAToyr5s
KwCbRsev11n2hik3xKLYbsXhdMTAi3Tznt4JIdcP5iJ8gLlvjJ2n/m93le9G4X0/
ux1BBF9jx/BIdqFNDaAXY2xYRrucvqg5u4FQRgTtTWJbjO2xTzJqBf7HbG6F6Gph
I09hkp8RikrI7ipAzMeOhn8qHU0t3dDu4vg6uQ2BsfCr3SyZRjN0hpqsv9MtLcZl
bL0Nx7j1M3ppmlgiPl77EKk3pfF9GrkxfyQvdY0hzdaOYglIjplpjHpU16o8fJX1
ePTG1nElVOQYELoEwCToFTke6Cb7cD+2+LtMbysfkaN8Lywi3go/hT6ysrb1lzGR
R9UTigy94vGenPVHWPrF0dHkQDPSBuJ+GF4rM8g+tGXAcfOvCVJ45y607ZsM29UX
I+favdnB3w4QFKbum0P3N0sNnRruNUMK7xvLg7TJhjDAmoMe6GOnEk+DZOh5a4W/
lj8tldHsPKzYqX/MT0H6e80Ygo9FNsUZlErYCJeOWdz3lHlt+T+hUodn0bn0GshM
FTC/nN60LBS3rrKwc5l9AtlrkLtEq3PcKlGvwOmsg4VYNy33Nv+REfGykvesVqkV
GcqssHrR+58kuO+lDPflJUbk1/n2rx8vvMqTtBE4leJrYiRdIU1ZtuIwnvLfH8OQ
q5BOaQLkXqJHqRqEylEIsskUWHHpwlcuN5ExZWddolxLd1rXMHzj9raTNOi+AWtC
ZUtXlh/8bmL477LNQHOTJoa6ONevoaOQ/ar/05T5i3s+K0Qu4sx9Bty3KPGww+g9
9OgI+z1+DBiA7KDAEvFGcSHFwogAredXOYYbIFmocz4qWHEyhHkl7XHLGbwmV+ZR
PGmvIgfdW15LONvLposC+eNabhvrEXA02sFCyNCqnNPQNksZPkBu4s/ammqixj/N
VIntE6nsCEMGVcMnQF7QyyJtfNNzjD3tH67LnSBP0r1G1kRygZk0MpQL/EFu+ruS
WbhgCJeYXDLH/02UIj31ifXSLaUrbVbQ6ngXVzyph8EbJXmIAFJo1hKT8F5N4oJ8
DYquxZmgseQfXhZEqKCSnYzdua0SiVc64f5N+8khH+COR/CR3OxKd4kACyRQLpg9
e1bChhUx2P14J6GxYNNiHrLK06HSelDHNQgceg2you1kE4zqAOHnmDvE2ZFN29fB
TVyOWkwu7ReaPW4wh54KA0Mdxfowwi4foae8GMTHURc8twqopkHhky2cKIxOmhjj
zplF5uiRJ/iQn2TrTTFwLsAhmOl4jq8DavUQUVu2opqN46zQUfHH56Xbi/s4UeUF
/rlNKMppDJx9ft2TI1f8aGUEy1oSWda0GV1huYW/6gg1j4htRuqoLLLa8BbKbuml
LRTPStTzDez0aNvAZkWiYlL3a/AeVzO7R64HVPp0hOFEotpqasHXEJMWWQLZqSHQ
4ygme+ySL8UdnKjtpq8MAL7WT1dpIB9fooPgHZthx9z4xpM4RCKq751CZwPKkLHd
UpcXnD3UN9l1ndoxR+L8Byh2tZ5mz8+F0FPJbvx5EX+e/5HsHtA6Ij5vuhYhMySu
PtIUGpxtpOJlbTankZslcqO19d5uuGpoHiPeAXL44NBreLv3TnWNJD+9bp3hJ71W
H5u7rPqN21kqHnyq8d4BcVULj50di8/adqd42u6S9ZTdXBkJlqHRQtGMYAoKprD/
n+prk2HMv4d3MBgoppd3ChnrkgBaXcu5B/VnKKVlb/oTUnDe5VyQ9rCoUo3l116l
a8Qq9I6kWX2DYEDR+lNEtuJz2rUjKd7yZs8LhlIWn47byOOU94y0abzGx+sMkvNC
0FhlpSQ3XJTYnQzOZCn/WVZZAdQClhxuVxWi2g8tf/QB27vShUI6zWYVUopr44/P
gg7ZhdWQpU4Pm50tcai0BnN5nLHXY+iYn7OBWixtACVK9UvWQM7GHMmqQMZyh8Jn
m9/m5IZ0H7SSEg1luuDNBX+Nc+THet72YpLB1kwaZNkUBJLu7q5UayZ8IoqDCrg0
2FqMrbyQv94Ee2faW+lqMsd20FYUsa5otOJATPHsa+udxKmu3qiF7M+WD2/ObTen
YFa7MZ84OlfGUFK5KUsLuR3nPcpDhT+kpFcfP1qymzjTU1+rzgsY7SASenARRM4i
7VLa8cPp5negVhn8vGlfapMjVSkn1DH5kaRqmnldXqqm85rwe9wrFMuszR5+zqgw
SOylElCeezox9T7fZELdkILZS3CoSzYqPNFkdh5PMxhb3P/pZvY7/8N+W7n2o/mW
e8FzpRoPYFIcaKJ6K9xKWY5qBazaSSnsDp9aEvbUrfRFpmBydlBDXZKYI7j/MQsr
jo1B+lxztNjmMYLVn8nfX1xyrlc50yy11zr5wzX1OlPjIA8DK3Nb6ETuTM2Xd/af
uPrbnVfwbTsBjWGCc06ZM/JtUllT/Ui/+sNrHfMRo8X+/C8Xg2K2iuK5SJdB3OcW
iM1i+fMQTf0ws7PVE1B9fHViUCGSJ78qKc+diTxDpwERYUhxAdABk5Xsk6cmaOuO
6fPLHfeTuHSFQ6MwkjEmSWlnyOGfPTLx4lU9vRIQQC48AwNAqpNFFZgFrN8sCeJ8
iHp7bgP8KvvxKV/6Diaf6LZuCGeg8AnAhP3ouLsITmTBeCJXbYxLrG+YqfRLdTXS
vjOMBTA+fhftmdfzA7MdeGXmGKSFhWZp12s+oaNyUrDkb1n73zqYTpBdGGQRl5r0
i+3G9cnzxtvnZ04ntrwKfdxD4UL37nH3w5E02kRJ4XPTqc6rhja6CZNS5A1bNlPO
Ppcv6ylUPQLyA3QMW84koLIEdpWsbCC0aQpxZXGCJ8n5YiJhzPYudRf1VrC5LQGk
LdWhe2tVntdq2Zvrk6EqjrKuLC/wz+pE2yVDrbJcNo1ehqSbwBNa5gmaT5LqbmQV
NeHdyJ7cuOPUrL+MtEW0g+yqDe7KMnhmv4Qzg2GtBS1H1mL6jXmWmLRAArSjD8g8
m3WevJ1NuaIro2mJwOPCNlpYPfxio1N09uCdKmMtDGJiT2NX5gu2xkanDData8n/
0hjzfvIiunhyhaGYEenzQqisOUAqy1o5Ygv/BqEZsBi3zLKyA3albYn16pcHSPlN
ypgXywbXMC8OMK04KdcHDZ1E4bOLRm6NAyK3Z8Q/TsF4yWZBD5lgiMx85nSg1pvU
laLwmVwHPTu3N8dwDkNIr8h8pbwliHUmNIr0zapXHJRURSYJYR4Ssep/Ed4Sxhov
jBESFu5eSf06XrTYCz2c0wgXG540ZJK5aKT626zSsHClJYR85FQdL4vhbict9/2v
J6Puk+icdO++LxkmTSQz13FifotGdOq+1pHLhv6xSEHK7+MVfFPf4u1KcBKuC+Vj
+1aSo/0P0NXjg4Q0AaYIl9qattvp6dFXFq0WU2NYxG6EMBxzlMty+TnKgO5NNcVX
NaIVmhFRmGHqsGaV4EHZL/PXqwHX0QUlqY0jivGXVA+4ox/QvznfOQYiCM3L/6st
Zm1YkjEq7uq6/g8TFuBUjKb7I+XLQFmkslS3Pie4wnuSkJ/T6EMpU+MUtdkW6v0q
fz7Hw19QAN35527qgAPgLByv0qGJ94gFJnovDOh1sLUkS3SZNC+eaijOadINTD0k
CfI6JI/sKeA/P7qWuOZGdqwXQnmfUzOKNhEoAjoDeBtF+K+8RNwBrMmNGCaw3+Xi
SuSALC9LSjjMll2Bv0Qsk0eKFrRGIdl2W7oSYy8+el2jQ50Yb1icqCkWoefOyCGo
W9Zl+/zNtYdlRNejb1xZc72Pf6f6hujaGmAnlzCvRyBm2FBhf/1GTzfS9bAf6K/8
EjhBhMzHYQK3kSkcNclEcaPzSxVAJZoPss02Fpj4+hr7dCF+O92ELZDXbsatTTBA
ClFENqgQfnTUq7UcADAiN5S4iEcMWG2hGpmtMpmpeoBwynYAtLoBLVQ5X7w3JHZY
sHY+rIjY12nEmm4lbgjto6+Q0SU/8WzBSMNgwCzrJ5D5cpOkl9u7aIongnwCTUTC
BKmdZKQ/HKIdzqtYUBpz1GJKlXqkEu1i8OFTryKpZHSLu6mV6pTh9IcilMuA60KN
Lvorka7OZhWRccYj5ncERnM1wOvzRGNqy/9Rhbv/tcvAxXab6R0i9o3ltMgGrxFr
V1iD1rBFpwnTapygJyu+YsMokoebaUMGBn7bh8DkCrjMnsk4KSNoK8kGastUfMFM
dGnJCiTmPW61iFJaGD1/YE9cXizXze6luLXY+xWnowIAWOSW1Pa07Zxi22uLL6dU
E34ySHHsLc5/YvLL6Ytw4k01Z/tomctJUd3suAf3uObUzT3/a4NO0uyH7UcloCdW
z9H7n32UHjEYeY3laeM6edj4BMurGXCwxS/PKW7lCLiu69kWIEFyJTVFjqUTltL+
Qk5wGds7Eo92OGnAJMRBmsNV4WUQ6/WtCLBuzeL1Qk5j5QK0MCJXpNjV+1DOaFhR
P3B8fnM9HeKVJvQuSHBGTXtZzw9xlDTMbz+1s3LZdBqB5VnY+TnBkBsOFF46yrGG
DwtmMpeNk/0DHVglsyGYhiENlbVUpIXX0n2mFcs5sBUKOrI7a5iVxRiA06Y2z+wb
3vNGuxZwjUpz/F6g2m/zO2Hti28Ae/EcqUW7FnzBLIkAtWI//+pF01gtXO8Ss7mJ
sj/YHRh0U5l6ZSk19xm63oUOKbuQFAliW1qCmtJN/hLYkMqVKSYt2H3TXULonZjq
cGJpOAW6JQr3ovo7OGa4p6Wu40sql1SNi97SrLwWhaDT+wTGvDFFS64J9Ln6oAVM
qMzil193m4I+0j3Pi3/eNEeVmnOkFKfdT9rNSWnY6m2tdtl/UCZo0HGIuTi1r2uG
2tvVYdxdF6Ew6GexoZh0lTMhHS/yswer3ygVES1NrateQRgu2qwJGGc/RE8GYq2R
sRAKHv888BQmxTzo6fXNoW5NojU13iLcYzQC0DpSWEUmpBkFAKNPpY8f6EXI8Go5
iyr+vv4Kj7eALocwNXIgJAplweFP79IX2Gqk04Pj4yph4PYUDC34pBwaKFmxwdk0
GiUuXQjRTBhKRNOHdSZ0FB3SSjLYdCt1e7M9oNN2KCyyaCEAB94IwlpAwx0PmtB3
a+Bibk72BsULsnkM863SJxOeqJJQJi/3b4WuEDH3V6T8erSd1Yy5jUZWXpNaFRjM
KCvIbwrCVQCkgfoW8/5nlFYSSYbbCTnwWEKKGjBrDrTL4bpnHMWavTd4Bm2RYcwH
wrMMBWZxTwNkAyGjy7/AVxN6V3NNTNL3SWkuDCRPvsQd9Y6vlwzbSUhdTwVUUPbj
2ep+l2mL6/EPk4rNEks6yPLJwcblcA1hrkyZpojzk5p12qKWl0BQvNtWbvw2tp+P
pZa1u3kZW5Q7tC+bRw4k/2SPNpkAxNcLaPrKb63zKHKe9vhMTQmv9jlBqQK5+m4M
ViQ9F7PVE9JuTf/MZ950qEem46UcqUXMMiROXPTqTSTvLwiFnoIxcBBSZjGOrKOV
JQzT8W23MmgVNxZqMwIx8ZzfS+yQhc4tEhqYL25sOn5JzFKXkNeqlG6t0NIN9S7s
CObbm6YHgNIn8TuGPKIajXODJohle+5Nv0G3mVNY1Y0luL/ZoAB/CnCzLJ7/LEL2
3dMdEBsNcXqYV8pFxzX4O2dz/Nvwp80HVPkUT+fmqjdKRezeQHKCT6VNkHKZ0ZhQ
IPo+v4Bl931tvjXnp7apTL92d8Pg78x7zyJfXA6Nd91prR+fSmeJFbDdkd69GaQl
lK2Uju658zWSn32AF5TT7fHs5dDNkSEQtfcxgPXiT2a5KcwAM3Z9Tx466F8rfxRC
IvElbRNh2JJMMzq9bUPGvKrkxLc8RTy/0oQZEotWgfb4k6v1GQHHmuJ6xVYK26bs
kcaxOiL+lm/uT8MlRyj5WZ3wo1/YR31NkU3w1vDdX1uUFeNkGSDWtewehKN5zMDo
lg32lM8usrpZ0xvvVTDX7DmFECsH/0MhsSb62ofn9f6gZcelxXQNV4IGgXPe4RQh
1nUfGgq1vgsGsS4/1LVwfm3x5iwrV5+l9KbUPrGD+wD294ndPHtxMhH6Tfc/pGNx
yAVdIy8ZhesFIE2rwkS6E17H4WNUCIfvvFO/jELd7WCYhhtFHyDva7QuYZUG4OoX
fHw5TfZ6v6mX54ct4COEirU5xqwOcGLvPvWB462ECHdL7H1P5irApKFOky8h1J7P
g6e8FierPe0+Ra9YUidavPC2lK94DIiR3cYG4ZycLDO2HpEy7DEC7psTSGWj0pJq
jwRd5Y8gX/RvPFb9Gq7T/DDGg9vkZxVGlZvE7HmjtbawEt9IKpN++W5V2PIAmKrL
a8yS2cj4L9H1j6+17AR2dEbmFfqjtn0cc3soEjcCJzYKaTi8ehGxq4QOy61VJrG0
Ru/xt4NyZ06l1PLCsu3LEsRFfFFYKG0lvAZZ72GKjZwbkMNFiBbUWZ81TJ3LXM6i
gSfeQg70i1UwJZnZq6qXvjAbKnw/kPXb8OwyhCevnTUZ4HCraNGRiCyqf3U543w7
KIz2MCANZh9YeZJBZdTYByrQdmYZ7ervAabAYkv6Lfx+Zal5hO9wHytg/wOtj32R
f1IFZA1PtUTCYSSucg/vfneE38uJEg06tFEur/EW22JNHOi5r9CyQrXA0F/k17KS
NJZm8YeFM5P+f0J4vTCMhy7Vniy/LTcrZaRPiRKtPKmATe3WYGCn0Me12SSHchVA
YEfs0YEZt+badeAXbV6/j5BdLU+vARwk5ur5DvTisH/i98wt18Pqz7gBD0tZNTsI
ywRB2b5d+IIPVtWgEkUwdKDAx3icv0jICXfBCltPno3g7B0hGi38/BACwJVuZLTK
xE43/QRGhJH0QlK+qTgxs6n0a+38PQNQw1IqDejpcECIwdnhLu06pKSZ/LgpHp2t
EBWn1vWAn9gnoiABLfgXWk0B4D9tprUYMxyHCC5np01kAUU5UEqXEQl9dPUa0mo3
QxucqB1lOT9/Qkim0/qwZwiTIExppGBpwoBgkkx2bPl8MIp3Vkhd1lrfksd574hz
3oO6u38Nxi3I3n1XPKauMEDplVoYy1J9/BBibdCqMjYIbNg1D6N1TLXLLv4QCkE8
FqWMBiHc8ZZBJjyRdXVY6buzP2mDT+BNg5XZE4MGOH/RONXd7nUR9j/jM5ucp+TJ
3IYXjYntXpo21ULz23uQugZ62Jr955sSRMfFieRm4+2apRmwUlJop2o8fLQ9gy1y
8L+JCdcGyTsjRuE78bH5kpQvhQMOpHwvWyzKxP9kEKZidO8NZY3xVCusWouRXymp
sytTprq85WqBs+Td+ZBBOQfqQa6qjPvXJZJ7wMKZmLaWvdm9tO2vRwz1HPedi2Wy
qtb73oG2/r0zPzrP1WJTVXrsh+SKNm87MDSV7uJkTioyt5XdoMmqEtpjbHlVj3cn
i1X0A+tJPga5hzhbnpd9TTqMURYpiI6fXiTzinRpty32Urn8uPVuk2MgrKZmrbDY
+OucyymyInSDPspxElORf1njjgtFWZMBOwaMX3BEy0Yufq1793M8c0a6Gg49O66R
g/rADu2mG2zOpXG5HyMTYTzpLJUMTccAYMmYLAZookDBp09FXCY/r3lrr8cl2kZP
iWyPW/+fpULUEdg7Qb4jlw11VO70mRVJSFitc5Sc4WNjovb0uX8siMEInzTj3uZJ
UV4rLmJmIC69B2E4WLIawnT71vcUu9pOEnuaWZCQSkTJq5OAmRwRvjtzAKqflUdF
QP1b45krFk5nhqwb+Zdx431DhtgsMngy69VikZHbcvFFC4BdQeYaeM/g3ykYT5+9
hjIfykJ3/auZXsGt7Kgvz7V/04i+u66vDTUNxLRts6TzD4KLjKWsjyL4FuaGs9dr
dFeF9ZpzcKnQ8blMENHDcGO5B9mq4+QDobXtrp6GNJ3usRqp8xsGkpKdODpe6Y2F
2DVlIVAKLSRLdf2WK3jZ2uwov7zLt/BFQaunVv04R7LgesPJ3RzkIT/jWDK24Gl0
MkQJBBG18fx2hCZYEYXS6zqMgaiD4K/YIwOtb27appRYxhUAPvwKTlZLpKVCk2xz
laNwupmglOqTFrkAAUL1ch7gmvtAbUjsl+sftVRKMqdbSRjaUsqAHK6WZIxVFdgp
bs5LCNl+treKPghDu1eDZkkyAhqTUYbc4QD1rgZ5uew8gvrgnYcQIdFLHcY153HI
W8x4Cclp9ntjjfq5Q1NmJkIPylXkc8HCINPjsgE8ilysR47H4hwamagMKKPHtlFI
uWcvyYwFEDYPJNbqekkJxUR3xtLZUdI+uQonSwqGiqYpUvIaaRR+fODXkW9EoSSk
6Vcc0YGQfh+EzVLxrOzugE9sXdSExjc1JJ8bhNIfQtRzbeQwp2+/XFXXtUMBcY0b
H2Wh2QUKvQV+MnRVdZV5aBOGWBQTDoyLwG+dl6FGJA7JLl2t9GYTx1SLJgZrg3ir
djh/tRuC+kzgmS78MgxFA75ykhwDoCrEUjTRRc/asUIutqcH4/g7QFslD5hHh7zH
YTkmOl7yCsYAvuhddn1HHJUADT2JhWwov26+UDO7P37B3hJStz3hE3svNLTf7vR8
/ujsiTQ72fLV5fhfbnaXjtlfewegRn/vm4MujcaL5q8eRGD6ffRsVSpeMbwqMAiy
dPwPWh5U1rDuydkoyf+5kXY39XYADOv/jMSfT8aBR2r8xR3bC4KxxyFIc1Mq0QEi
SJNToxebfxHFtuVaVY5IaAfgj9mvnjjnBN4ojEcUsIXWncfZ8Hlg6Ba84AahL4Fd
2YUZuEK/1+X9a1Mafr+tWn/hf7E/7Axi0Q8dECbBJsSw5/IO3rdXKFbSMHm9rxA+
wQysTYoAbFvP39UyT0wQhe1SYzQgODkyADIB4mEX58pEd4utaC1thtWDozcCiQMZ
f/14Cwsdol7GyePuFwDmECC+WC5znurJLdNt5jAdVnhWSnBOlKKnfjJaMb3e5UtY
WZoJTIFrIxda7LoOmweBW2RRcQI9m52x0Ozmkm72ZPaGCppblh7gV1KWmbkFDCmo
f0WubAiS55Y79/GZ3G3adBj79lW1rHZFEUysmj2rk7rE2EJsEHW3r7l5kMrbSu7W
2BOtznN+m8HKv67n8N1q8wZm0IgBTas0y34KeYoZiMtPXR+8r/CZVhITqVkFB2Mn
WIUO1gRMK4hvD6UevRQbvo2oc+bcy3DGNCic9mOK+g4YyYj1AKZVxwXCx4PI/7/K
CjOyiu6wm4dDpkKgeo7ipYRemIIcjMqdbj+ljG2LI2MoJEppPr4/LZQqyVAMD/0V
0wNJGecBha8SEV5YZA4A8C39pa6Wtvyjn6ciHTIfkMffEPYx8n5dWE7Er68wpFWA
vRsZRnoJOIss5b2LNGTsEpadMn2rsXweR03uNkaUW7bTpsvbLpo18bjllouzktwU
t6oj3QD54Z0SWdocSh7OtbZRZJqYmWyGCea8g1dpqEgt+wWzwLbriOJKkPfERVB0
Lr4Ffg4pdvi9FGY+KYrJ08OTkPa8Rjs7Oaeqny6/dlnBn9xf+xOGTqqJkQ4kOVcT
yQy+tinkvUvu70XNcgn4lePbbYX/hdg7FO8erLlwT8JGeUW1xrqKo49oVyc7vizH
KcFIvrsP1lDKsHNJ9qPo+WB6s1VrO09lXGi5YN13lraND7y4Fk1VkdvaiAs7Pul0
Dx/eBVLgyxTrubSQFkmM9dQDBNPKiBWBrI5OReeTTwoAr2d7SLT+tWrmVDF4Mw0v
hfZEX48fXbYU6aGNlnDbBhiYBHNUG5mb+HHS3QsPtx4KGyT3bclcKj6XAO0B20sJ
javvh4zXKbomjAXNA1YPIsj1tKQUvMwhOQJ16bhRY8xKjQi3jDes84QWfB0153+o
i1tguBRuWweY1oUMaUrW3nWmOA2aWSJKrAhVRR4q7C3lN2quYV+u3y1NiD66Mzcw
vnMAUqNldOD9eWB4nAXqNvNLVMx+thOnJU++/B41KWCFK0JGX/RJua6+seB4/SRF
Kbap07ksT/aIwGRCcNvzze2KLfqPj4LfqntaGDbHd6dQVs/kziVzFtYV5k+2FgYj
eEtidQRrj3Q4Trcmpt0DuJgRSo01a/8L83ubD0ApdLbZni1RTjIWMHteEmLWl+z5
3sjWHd1EnF57ggkcUfpVGcVwkqxQk0ONZziL++fwiqKLpXN46BqpN3jgBBq+i37P
AKmLMuIeHWQJO3/kU4hi55mPo7sm57zDYt0i72BvFCYnwdNPu2aQoKzusvCj8SD/
sTnmEuOnr8foU0vswUIGCkE1Aq0ABJ/YoMlgJnV6WOlrUM7mgK+LzGTLnfCHCOgX
YaUIWWpj7JlboX2DgODjPRR+XDgPz4fZapKaxBdc+pdTGcW3JOH+Rw2BMbuuEIrX
Os/H2vLKOMak8VPzMe9SKT/yucNcqUJP4msBxQXmW4cjuYBh0z92BOKdItFtyx4A
vett+8/U74xSMjYRm9syQMIqNlyUNx/l42Jy0UFlVJSpgh4JhAl5HBVJl706nBAy
Ko2O6eSLxSWYM4TeiKZZt6qQgQvwxXmr+avPZg4tfZ6XVXdug8KJaHgOHHtgshTd
YCIBBos4U3wuyedXjoBqmMAe0AKGATFk2hmqJHy8zY0sg5cpTs7FlZ2qMonesaAc
judSuNF1KTEwHBeHYY+Qr/49W5Rf5BBZTVaN8nNaxB1/YTfuZ7c9iag27EQM6rxR
bzPfu9tinx2vew8WyyiNDKoriRD1KjTIgpuh51jlJgBlneqtYXEMd4UqRtg/XmJk
a6/6lAzRRheu6ABHF8GOe33AH84Dhqqy8jJGImyEB/GvSLeg1R04cGcJuqWTAAEY
Fj4OCrh1L3FTRWoyIvUNwLHY4DTQ3uOBV+FcK+qZZIHcV0BqeBRUwvQ/RJT+oVIQ
q23MFqe6pqDZEnPKrYK3mZQz0paAi+3PHFYKm2g7f5wQDAN4wlBJl5rF1VnHax6s
hZ8AiLLeaovxakocvPo9RRyDrBNkWntzIciWQyXm8aq8aHJdGr4ApczRtAuQ9Itm
xnk0mF/FKcRIGv9BWFQEykzQnohUa1GJU3AhArxEZD0Rp4Ub5ACj3YY7cEp/3/EI
VEQdmf4OCh30+6kvxSxjJpxhYMt9MzO4VvTXn0c9neWfBf1/iUZPH0Lww0l7nkda
/wbvBjBDLTMs2yW0eU8n46EKPwA6VJ/CCAEljVJUKQ5W/DbQJC8tFF1s6VDLmyOR
ps2PHItwSMj53tx6YUCKBwOdxFVYm79tGlo7ilNbF1LUWb7452CkB28uFuEoNQZv
XGz2shCZR36YOoMb6ZAPP+asIsx2pUVs04NLC+P1mfpFn0ufgDFjU+nGf+w6VTxI
8NSlgKPRrv1EAkG8h3J+ehbfRJt67rl/hjyTzsGT5/KLfvioPm1Hp7gPMM6+/xl8
nCnGocN8jzH+WazSzm4TSeg5JflnMJsGQzX/VAfxZSjjF4Pl+siuQSd38LJDfn3S
rIMeE8BTfN4DG9boKe+YKqiRE7Bxv6gvKI7wasRn7MvR63kbvVVKUtqszj2MePub
sqF8zy8DUW+zPjWuhzUsGGGSD/3MLxCjL69Zq3Q47+Q3QbsWBe5wewXdIka1Hhxh
mHVIHLTC/hE5l9BdvfCr9WjS6qdcCxWewSoH5UaKFV5z9DscgCsai7vTif6WYqt6
ixsJ2pyt5EUfWfXr7qzypM1kBImTZegz7KWBVO1zsCDfAlS7VKSqUDV80deOJz5T
lFPznFjLAcH/RaSbWpoQf9naHdUMnu5toQ7nqVryCDxD3Lg7viEsuUgK9qc4A3iq
UukQz3re1we8WwYpOKbBkcCfQpT6wuWl8GvpJ3WfHt6DeY4/ziEBysl1ZpXMARki
FsggNdP0bqSCaIohvsQfsQy5rJRMLSj+1ppPcaw3hWQyZrvsp4Y0Qv/Gh/GLAqhM
mSoaYN9ZXKP0Sv9liM8uGLvuMgw6nQvsdBhcwaF66PIbFV5F+6PGD7fO12CoONdK
6Y/7gQ5x6q/sELT6pGQaWQC1qyh6FF7yeo+0dRQqensiSY4ykHBY4JWb+HD6EvZC
LX6Yz54nwxbqGDE6qucpDHMk/R39U7pxmlUUL/JY3NIOqqa92QaDNetIrd1Vetz8
MlZTF3A+6h0VeacFBPxPEnvKpHAJRmNdtSZV+ZdWgVMtUDKk/pqdL0bD9NTCaRbG
FNj7K1e4BFtngNpkQya9wx556FiuhjOdHWVtiEbsQ3UlDUSiFrKsq7lS5JfO1O2E
YCjkTFFfuNbDppl5xkitlogPwPa0394EE5L5Mai3aMx7GQVizkBJkkADN5OBgeTM
CwwnPe5iHwh7tdITs8PyaacJkKHCWF2Mkgu53jGAd2CBr1xlUc/wxqaEQ0s3vP9x
BKqJPqcixWe3Ds5JxIedQ9Z53HacZh5vgi+Yldf/79Slx/0qmdm3xU+96olC0GzZ
XMU4KuF3NLQRiTuhG/DDxMjfoS5DzL/9TRAJoF/UbGRbOzNVfGNhRME44VeeLv+o
IWoFUrhywF+X2Kz3GnQJ9TZhsNMAGxfklo6M9YS6i5uIeJb0bmu2qU3ahUZUK2VG
C68xp58LObXQEa1ukUGfiG2wKkDZWJ/z5WAVn13PuEoXuPmbYj86mPnzigzoYbEm
WAbmJEZ3ncIpUc7HvMetnFaF328VQ2zePoNTSSAHBkwLC4/jNX2Jf8oWnworma5n
pBGNLpIgBNwb9W7ivSiEUQ6zOAEW0VMXZGBdRVXpR1aePyQ177tXoA24oru2Bks5
rtgPGNyZCwi52TPVzYRZhWeT8aUjkBjbFnBDYmt46uei04Afo3jC4cf5ldfUPxNd
SDddXAlud4lCouAW0jG7rIOJh28X3DD3Y31IbzkYbojogRobdkWkaDdbsIR/mc4F
5e+UN+1Gz+AXDssHSR0+0BcOR0DzlHc5QiM/p9JOpLWKjgUzqVzhH+E58Pm9vrPw
t263qQMMMtGT/KVMiLOlX5aCy7knqMtBgCrFMuPNvqyr3H6LHyl8xolBtjY3XTV6
1rM1avSbWg27U71lV6M7YfehRWs2XeV7/MDxa0QjT6/Gp0JLWJNo/to+lzLbM7z2
dEeTvXKKdWkQt7xMtstvTe63ds4ufPex+G32VN9h0tGatLzQmITDtfsQWPTI5p4H
u5Xq5ypgltWolqlSrlwg10bcCHvOJahc2DKP6YyVH3RxpF9OlGkx2Fuio0nnrij3
vympgcjTjTnxeu9QGvwtmgSUJF/+dZuVn3ErX7WKQJ00mjl9ttC4qe+35bHfp5xS
vAn9IsF87P4ToF0b8WNYONL6yUQDbAL/bTh02roH9FQxhgIHS77u+7sVSwdlC4AR
prPESMYVsBL/anCVim5l4eOwo/RSIN5D3rSAp3xPagP9HOS4/RjkeFPKZ7+iAuom
7DxSrkcDKzKazYuFf+SjnJBeU6CdMQ20xcUZhMLSyjcBjfG9tmbYKdgq8wZvk0XL
LekxNPx91Xkvp/fnLJS5H83LNlJJwD6Kuw/0ZPwk8askXgky4j41Hrkg9HWKC733
Wd3JuJejDuijRD22gZImY8fNdStUap1QXUWBGbATst3veJNSQLeu7ufDFpCUOcIf
LVdF69mpHNiLZqF+JM/8P6tr9CKEj+UpHk1FO7owSkM9G/A9Ym8sT+9JQ+y7RHIf
L0vi+JkQGpG8sccN7WC2ieEJKBZaat/wreCh/PNCTK90EogUOpI0FAOJyC43K4SV
QYOR+7HtFa1N+2AdBaOGvi07i8Uk1npnZIiXTYdkp21bIjumvsg+iuw93qJm+0x2
gZG6qOVT8xXhhLOuL8PeajrcXuz/h/ijjH+C2Zu5wJ6BaWx9wK7tXKeql3Rpayc/
5v9T7R7yeiMbR0/nFwpTzNA39v/1ESb9ywVBNJu0d52LMv8UFY/qjqj/OR7UyF7U
c3Z6lyne/DZN4ekzrZ7M7gIfRWu9rb3xfh7lVfZWzSrft5Zxv6tAEgiT3wNRW15x
E6Z4xPXtRXOPUUicIXpVP0B0lF91o+FuSVNY6TLQrj/AKaoR8Ia2F2b19hut1BVz
oXdM5cI48bExnM68zVH36oPIHcvTEycIAV+1Zw5AfU2QzmhYueh0aX8hriLsC49a
u3VStzBPOGcipRItyOevtlx/jrkOPs5gQMA3ys2YrEVIV0kzATB4XWgk+fMs4H0V
yiINB5bZQxJY4pY5FNSu7pEVEGewRDwmxpNbHWVX44VQ5NR98Xbx35QaL0hikK2Z
UeA4DiYzuMUV8HucAD+kFta3htL2KOHZE7XDdCJhXXXogOVqtT2ibBZWE5vVuqzj
DLLDHAX06LMwl//1Icmy1fP6/tggXjySq16dhsBpb2Q6eBy7rsclMTidTcHy7Jqg
a0Ne0MbA1frPJxsemCDYJxMzlH8iKn2S4GZ5W68YloNIYCj/SbIsSlo3ev5TT8aC
Uc0xFsYLrN3wOC5aWwr1mJsI3NiWPL4/McfHdnO2uYCp++oFKoQ7Bi1aV/KiEgvj
6Di1Os7qt8xF8EnWQlBloxCUr0VegW93AaS5bbjFmSVwlsawyK3OgTu2GApN8k9C
HScw5+SKH0xZ2CkAe3GRu7GP39Dk914gt8kDzxF4sedCfWY1an3CL1NWYXRn9Ul+
V3QYn3IGDciQch1l/DX+JHzpB7r3k3uU+stn1CmdEnRf3kc2QOA93J/6Y58H3fx/
YrUXiQHB6zSk+VVcTJ5PJ9nAX29KrlXeZWSKxJYLbDmp1U3YIePrO11aSoR2BO96
hOW2p2sHo9VojWKmotLp3R/RbF7N8dSo8Qlccm8yvazMeQrRWGNi4uqB2Em0yeFQ
rErHgEwrkqPMWFNTQo4TLoXNMIYVz15BM9p/g/Ru/2w5ATePkFrVVcwrNDDXZaLn
eXnLOpXHPQoPmJQBlDjIrN2W3ZdR9eTfcm7RghO15urKS5crPYyXz8f15HHrfXjL
8nKqf3jk11mCgTKgPI3FFloqRcrQ8yLx4pQO9qv93lQ6KxCA7bLjEsL7n1kWNIBR
o8Kes+LqKZFNVemGrZTPoe/W1e9kpAeAtPDu4LFBAuu6KW4XvIdDp1Rz00mPb57P
jaVhABN1AX02tC8USBy18YavlPMZCtrXVUKveeqCncYJ5x6k/EEYPHUjVbRXaTmT
v0NPPrAkCq52mqDNDM8MNWb4Arw1AOGb2swNxFfp7OCvnPxSbeCvIf/5MtvlDeeo
5e1psHqSgQL8tgsK78zH0zxiT9EmQjBBuJa3wsex3yjimLuH6Dx+sw2T1p9XZjNG
gPD3IAgPy80OauI1+nTIkwLnAivrXSA7b+Q6/tswTnV0ZQl/JR6E0KnBleRobpL5
SI321mYDE5MlnE2fgt58pWljQHl9DNsUiam8oe/ZgtM817nD/8BZisfweiNRV//8
Uq74GuhYCS1WkJcVwRM76FHkkNPVnpuz65w07bROKzI4dWSPBwdvCgK/dkdRVktN
rK4qFUyxYWyjJDSvrKBGk5037N1BTaLpS48Zfej2alCLPRVedyyUd+HcZbU46LGf
J/krdxcq3rqBrJMj7tg8zTm2/F7B1ouFntvSCCUZFrNd3TiyIN9yi0NPOGkT+0ZM
r0KoGn55jGExjv5oHALRO3cuVZImX6JrZ8QmEezUkx0oWR0709gA8wDsbkuQMEBj
jttPzNXPeY7QrdtLvzEATS3Xj8Ua83cMamkY1d/c6I4LwZMyfNEJNkRDuIRRFjlj
+5wkQFsLDFenExdbmR6P7SdanY6LwmIm1MF6MCvh3qYh2tHRUJcO5pnXh54pFOGB
AXWYZ+B+FF9K8SoriE8GWMw7xPSAh0YJyJkkQSnP4kOE9lPHCtj5uYJJlevDCWSR
YgvJNCJysZbXiimRxgmA4EJudwQZR7Q60ibo4uJuZftAIfxjwX0IbAUQ0871K0L4
i1g4YIRdVoyEQUvIJto7XG15bTtuDzZpmZTAvVjaxsh+8yLSDmBYTouoCjm//T/A
ioOQOEeXIrLajyDgSwe9QSGwJKOg1wJA6JepP4QFiDFUNtySUOG89EA6VXU8HHxt
rRyR57f3KDm3kZtCKuVqZwbeTz+6yPWp+kIv992iBma5Y12bCd3kx2uvCh/Nuw7d
CO3w7A+BfLuytuSHwPOIIpbEkwOeV3aD3tYTHEIBsMAjnOsJif7g6MiUD6EOeysb
AfhysYRgJI8ovGQpi18FXWbd/iPg6hJ3NIpkMGIWyTOQExTDHDrV2aVGFbI2cuUe
+eyUFoBQ7vzdHfYm1MbKFLahqKmLKpF9p5OcWr2cX04LmeJHi9VCj3zL9i6Jz0j9
Mp0iYOYvTX+yPyd0RRQEn2zCM8x5E8QKYaW/8RsJ2nAWJwhR2ZINfxvtZfesOcct
jUifVT3PVkPbackTye+QsnQqc27dtyE1Bfy0BJDRmuVQb1b4n9f7x9pD+3P+cOYe
dx00kSN+tSuEPAKUBgvmOnC2Uz1cgAKuAyCS12oCyuFBXH5WLs8Ip6t7Dk4XbgKU
fU7Xh5ZGDyFK1HJcKWu4sZECvdv0VQh16WplTzmGbyrbNPFKvJYheEj1p7uyHXZM
cWoen0Ob+gh0PD2vxrZEB1oSSnmxJvbxypjkpNWQWViQf5Brz0MPWElh90KiMjxg
Ne1hJwY+mf6iZ9eETPa0wLbuDBnf+BY/F9tr2weEbkMKPjuwFmHXg/9/JJX0svOK
sa8XNYj2nHDD8slzq92W3xRPVCE8/No7CufM7fnK7mIAq6M+tPa1s86CBGw8OPiR
PfcUr6cmuLFXat4BmM9Xvk+vc1KHbAO3VN6tlLRa6omTT2x1ab/VLeE64L6PMbTa
xCiGNOAaQvZJIU3yCmixVNzHd9TsoRBT8p1bsj12v82vvjENEEz2pcwgit8DAMb8
H7vsv6wf41RbZIYTKFgiCE7oONTHSfA2zjny3zFZksS6CbBTnbbYDRaZZfGdcOLX
YEJu85VPMewWI3UEeCEVO6Ag60tTwaDCnk+Ey96/Ez4lSFBFBpLhSeNvyclELU20
Zdj0GFLRFX3QMLOl3mS50bNYIm2duP2TIwKjypEHMUhgTJfS0FJk4Wv4W4lMPBvt
Byy3ONtp8BDuByR95K+MnHyVQypKwcXPknHGuqXqw5hAQ280ogVdRC/RZWLcsS5C
8NvXKd24tUpFIgs96kJUBKS5iDBh0c4qtFj4LtuMWNI2Xv9qS0SGVIwyyvGoj8zm
rqHL6u/2lmfn0Ri+e3TUSyR1ON6urdlTkJ4hkqmJKrK8raEle3CLjmQkCaAZuBfZ
vZdCe8fqBx/sCe3hTn6QAc2XuIzuIE78VrryBXQWyKHIfQv49DjVr6rcQtbQ7oPf
/XQkAL66/HofjfkxCcPYVAVO73AVcqQPJTgWyNqHkVZq4m8Ou6DVczn5zWfP3LZU
ULQf7llKWMvAkL4lmUSwN3maelcfPfsUuZhu8+Y20pPajQJzIBq0Hy/PoEHSRmjx
OrpFUi1rUSd+WYVbQCvfPAH/hWDMKajhiEw1Uqfse+I86zZcOctQhjNpmfY4baAZ
WNjP3KiVW/GHP+G8peaLLQjE6EtiSbAoCQzEa7p9pK/3tXmUjyNJ2zFIOgeaaVZc
QSfQ5FvjVMcWmuB/SzpAoBY6WzONokRKbm6EOxCm6LVfrQShamekDZo6DvTAMv4N
m4LaoMHWaOkx9ZYgO7Fuu7tz7ntdc/HbLwMuADiJdgc+NZbQOhPuYzFZ6jyHD0xR
ybOC7QbFQWbCTpeX2AB+TdoWYYBHD1fXDTagzY/fOYdL/0yKg/4RcYqI94yxsBUC
5BnkI1S2RR6bgOEdWFJq355HD8KrDKQkWOIzy1HZxSRf13T4Ox2nDVJLJIxFGpmE
j/Iy+Jt1SbRLZ4fti8JCjjRR1D2c9jwBuC/TZ6NKvtukR9ZhoRfVlCjibiohxsJm
lzeFspXKwV9k+/Eg1KxADLNzZBGH31YjhQRM6hcW5E6QQne8B7VaKlx1xgtYb6+p
rsMH+HdJxBmlih0ipKbLouSfsPXP6XoVIHlH1y01AXKDIG6zPF3in9Lg+MqQU+Dq
8PEdg0axITW1S8GPn7goGwmW+oa2LtxtwrrbPJSAOl3clB/iULxZH1zrCbQoJGcN
TZUrie4c475oiCEogYVEUS/gcE85YMzT/XGOj6rzB3jQ+U7nvnYUI896vdUl45dj
0UffC5rO/jY4+i55ZpCknHrQzfJ2UR6QAngXWCQEBSZy3uh2qUXMKHMso7z6FTen
/BVD/v6G3ZoJYE1QYuxRISCwMGJV3+RXeYcuGI8Ef1CBebbNXqYU4yRsIMufc0zA
3hJmJSMy/g6PUa2I8HUpq2sowkqN1/Kt9NS+ucDRGd02H8VXfJud5SKhJ3Cr2JFc
nZB0dHYbP0cO/mhdsPjjVB5tMjgrA2u5hvBPzXaj12IjvCcQCXRePksg3GRSEXHS
Hz4Abr6a8eW8NQVgl6gik8kYewpUFxQWDGnRadUde9qj6j6NTPKvqltnnznevwUH
zffX8U0OSkRdf+DYLH3ps4FS/S6l+Tgj8bVNzuKFVsaWMoLUmljvU8yZ6pp/9wwN
liKPo4mEkd6yEqi4FVZWi9ekrsGzVUslPg4+KKi9W8Z2tdU+Sy7pe+g3Icjq/R1X
ZbAYDcf3KvvMGPTHx5/cuOVA+SEryWvCxMytcojsvW+87DgBdphp8A8UG8j6Ml9m
o4X6tLtZv/qzhsdRqwllwE4x5GdhJT8hp87C7nkJJBBACiNG3KW5Ibv7M2mRXqYz
DI4dMB+vpnCEg7C6hAsrdZDf2kyG7sVRuRHPC0/k8TcO7KdKcYBZco9Rg01Xwr4l
D2ZjdmUddsJwImzJT704mFLolWvqbGUDJhaSMfRCnN/xszg3ToT8vF+K0NT6/ySZ
0dTlPdhrgNO6bnfSvflDRLQecBuQziTA/FKFXK3NWewbMCWCLC7anVQA+XKQfVwL
wVOQuEpcdOukF7cHlz8hh2mAgOznbeeLTdC77/pGTQpn1EgbrX70HndunCNomLF7
W0L0hLOiFju7MpL1yqb4IdED5VuJYU2YmB+XB481dSNmjAytFTD20hp+FtYKNm+I
WrBMpju2jM4QQv1wp8o421yZi7dc6V/schtZBhE+PFJ5iXVr3imb6M4x7gCRyrgd
unPpm5xWfiyG0ngssg9XZMEdqzRMgO9S2+sCQxsRu/ZgdtC09fcOUYr/r/+Ubjdo
hQe+K14G+Ch0I6aEGS+1NXcJ/anR8BaZSE4rb0pbEkjL8KwuuaLeUq9DHFb+Ldvh
APB0oucLe6OQeIH/feqsvXxMDW5Ox0ymgHgYQMrzubDNKcOYHAb/fjPBQr3BEG13
W/OtCD8NujX5/HaREgL5oxe6nJBIosqSYZdqwLn+4bJXnbNrJX0DjPHVJRpXUuk2
t+U8NYI+8JcbLzzhTQmqEZiP97RNjnYlPrsvih4DXYaRyC8wZq3cV1BLuAL0d8++
mMYSy6i7Go5gfRxNcN1qSebBF5Rjx/j4/pmDP7Kc2/0+1np3gbln6RkbmoCA3+gE
ncbtzMRQutWgEQmhn/5QC3iJnQ1Lqs/+p2zjMLBfk/+VDGCbkgwhxrPGxcOL1Gw1
uRVjEhCiq4hjTTuzgLQ5gs46VA0NV3E6XcXmXs2vd392qwUgTjY9HAeM9jP7kLFF
IqKm0pePSrUYb8GAZFC9LKqgnIPwVGxC9C64jJ2nAQA2/30bqycRWYdXSJF3pcnw
yg3mcTJwkGqG/wYWS55TrX94QHSsab/12k7MTHD4YBCo8lSxSyjVesTD+9g3qE1j
kK5y2UsifUWpt/NOdPcgboA+MnrCDc8XADtzagRHRLpEmgS7i5RNBJKolNq4itQu
AK1i6HMvTY7KpNv5mgDOKsScxbgx9lGZKK5roEieBCZWAGB0n84G4h9FMMj6DIJ5
MQL+U94shfG1dQBp742z09LljWD2fp8VlbGAJzFjOHwQDQ2kmA3HP1BYYmDuPP8I
OwPKcQliwrNXIJrg6O9iT33Y6VpmPX0zL/Tpw/prNB7yeVoqW+ql3Mt+/vbh95ph
R8LqqkfhFftNdq/PXhsWgLleRqmIDkqkYWLaoFsFe3Kp2z2eZ6b0KujPFdSoV1Ow
4X+PD2cjS6nQMNpzZiPe6nzvObgQrqZ242XQ5zZSMSEKdSoteqKK5rj382fUUiCk
goiPWbZPWds4EQFW4JdU2UlRFqKFEvPIYWSXMOSKupkdaxsZn5+8mQ/2sDsx+yam
2ZohZljutjnN4NiHU709XkTziT+UEUKZGPpDmIiJJH8Nz733TVdPWKwgpylF5V+M
g03O45yG0a3fqP1tT1lP+2MqjfgyiBNc8NThEspDYPzW+15Cbh+XIgGjBtDcG0Fi
UvxFE5Jjd/k4OpZe9GPA5soqqhNpM6mtAZg80w0shdcsMqJfG1l3QHx7CocUtmGH
cIGVemz+NfTHSuM3OAL9AFtAgO06meulIvhrWbtIdl/VU6Aio3bQva2pk6xELNSA
T74xsKa/xG1drufMA7KyRfX00c3tQAhFaafgN6PWiK42XzgmZDXagI7D4+/w6Uoq
XFb1/LsBVNQufOuClWWW/UEGdi7kEKWi0vvLy0JDRJnk7mdYgcD/BShznZakA5/P
fyFTJL2PKVufVCvn+EpHJbGfSCRepfN8MXicUoOfLmuwbb6dSbZ4fJPqtMU7EYlq
PzbCKxxhcuPgsdlFCusavYY4Q7E2MxNk1limN5354QPEzWCxANS8gZBh9JGNy2Kg
buedDC2+2cNhmlTltnRun5/A+wI7hPxz8rygQP7t6xISvw5IFXAzfi5VMZXbkVLt
W3tHRwSras1curMJq6fh1uqo78ia6iKNlyPdXb0z5NvxHAxk7mj6DvWiU29wxqLn
JZvrXq+LxSmZOnD7lgE0z7Fp1d3Xdfn2OVhaIMGOyzoXQJu+jkHlJ0XzFAGWUIWl
W4IXu8SaTYuj+8sRIdW0h4O9GgpGqUjRIlvRMVMTTOzEWD5ohJsxu+VQy4SHB/pL
1nyNVVq63TMV5kozhDc4FJfg2mdu7EGvfSMg43WM9rQKKlsxmz5WCE3CaRWzE3mp
VR8I1ehgYUNOYyOsmtCDKUsGtnFIKc2Nv3j5jSuxYL+dJ30KUyD7L/a51UEPlpfm
o4rA42rbpdT+cGzXcR1CqcMbpNcKXmtPT1TSbEK1F3n6yTsBCYSPRYDIK7c/O/5K
YfNxSeUvNIy1u61hxyYWNtaAj2AzMaQueYCsS1UN1gUU75CN/UTCkO8AkHU7Mw6Z
MQpq1/rO/1GQEv77rvYNeg6bfDaEUXgnt1nJWxka1EjREHygw8bjR497fTNjpO0o
d4WPGQf8ND/rGBcu6HQqkLylNyY3cLNzbTZ8+XySPztUNTUDRsI/tvIxBqUOIeb3
XErSct3Ef/4cuxUyMuslFEE0wvE1XwaUtHaA+QFXVT8I8JMBJl6v5aEM2k0ru9vD
jF/iHqd8uIwehweBv8z+DmI3xga6uH+AoJx5u5AH92/yJauNZJ+duxtbexdl2xA5
ra7+IiKF3Zvodj6xKW7jtfXbUWH5ZQusNVVL7WDpEixaOOPZYN94CKW3LqcjRIjs
Qa5/6iTerKbPI1vkDp6m9ZhE7hGwDNEkrVMKqIXgKT1nYbKLihiF1vbiOs5ZTsov
9g+HuhU0XgORlQ/YjLPAn+WsweJCMQthti5BVGTSMjgodlJrRJ0bxSoNrD0Ncko/
pvuOk/dl+Ulv0lZ7B7V4gUlHFl8eSS/2aHv3LoDWfkHkK6Qx4ojxJuFQ6Zy2iZBw
sHC66+GWOxaekXy+CA1aFCB2rxfYgFpq84H8i4DmOhF/2MuRVlAJsrmuPw69U5Fd
bCOa36HyviKnDJ4hOr/ex1hbuDAsK1vTRlbafzRBok/dXfqQtkwotXu2ZkMlFEs4
8eKlqeqXC7dkD7qEOQ4K2/McZte5VJkMIGEIK5xvQnR9L2MCQdtqKah2nV7pMZrN
gqLLThAXBPZf6ebB3533MWNB8smlt9hi8Opj3VNLRJVIZsBS+qEq7oz0nZWcIHC0
a47tztlYIu5fbDFkLb2lVbys5n9FmnBQdx0aJLU2Dh4Xcs4YSujPRXsU+rLwUf8n
Ha9vbwWdCSvOXwu/x0ey70YFnLwiLx2ErOwejFo7+txYVb5jxIX8wvKMOnAnljiV
CsL/NwaeDTaznbdaMRjRo5yJJk30fNhhWLeoIDMtR1UaoZ3ZkkRIAJhWY/FcmgrA
fbnD0GWq3TC99w/LP1ncmUoz5ckDDnUwP4lm11QzCWSw33nXbdwdtRhMVS2W99DA
1qctkwo33nwLjQYrPvmuqti6wYnbpek9OgkgLVPxYOT04jkh9vHXpwxkzgMNu0/a
ByeQK2IYBH7izkfdK2dkOaNuPfYS0To6tL+yeSBpQbNSUpta7vwroqSFgHpJUNIn
ObTjfK/7XloFR7KA37qIUHRGLjt2m44qXO+kNL/ej5yyoQ5wzL2alpF5tcyK8ybL
EIeuz/T3anZSmeZ+kRvOgAB6XC7R3o+yAlwQEWqDKhLq1cEAnGnItiH/EO/+VkFM
gb5uJ+wIe5MeQYbl4nhh0YdOpje5F6zNM0t51rJGSkxRjs0ODgZGjI66h3VMCxvb
Mpz7ZImwwOrXBaoRFEBF+debaJ1Zlj98mgC1hoQD3SGimiaIdLtK7p3e6R8vONoc
S2T6wF8QGGo0UsZjsSuIYNdLjS+7fe+sRzXxRNw4jYDvjmYLiUXiVTBu4biWvB8o
Cfta4U/2ZVMug0BUgJkDYQtdaTIle6Ixk20Ae1byS7QjabsA7sS9fEk2Ty1s7Hib
zmSgqt7uqjnVQJ0gkbnMn4hwga7EQSzOBeI3DVkczdnT9SLoKZ3huqGRfWJMvvvl
jbTaPgfiN0UizHh3Ps3+fqg0UTbdCPz56+9g0tuJeV2Z7uChJdsECstvb0Z7Ki/J
rVH8pWacDNbVHlt1hlvIX5wN8FeLxHwcKrirnFPhcQAqQw2UEKvLLSEeBRNJbChY
vrAiIbuX8MsZq1GpnRxFPZba/JjcnYdzM5j3imOpwIbttlijaCtzGey407M1Nuac
NZtAlfIHa2Vhz9Pi0nvHN+EFhxzfgLVDBgLELBle08A3517wxmLtHglVE5QjTOHs
feFezwN31zOxxPOkom7HIDDrwWiburA3wE2wqWI5/V8gtXQN6nWyj0ggf2Y2sa9V
XtLaTJGKYKpHzW7mUeK1d1g6z8u3Lfeb7ssDajat/HVetZiRMeNCIY7NjU84TLZ2
W8s2a96HjphWVuDl3jiniLyoo0g2dhEz0Ndnd0PSQnptu5LqpIH1MbVyk5q7orL6
UHK8kxN2ZpKAlSNRXFgexv01h9atlsVzI4FwyyXQXqlKyArpZB+AFiUw25zqvMp0
mUSC3udhc+COM/D6Mp0xbX0fu7JQyMiFwA9zqkRY7n0svqtOIujgIWo0q8PgGdd3
UubTlDBHQZLETLxx1ueoExOGlc7kIYkpkL/ODSj8sil3ZsI7fCPGktor3Ia0ZJ1r
rMpRiipWCwWrW2DDxlMcLdqmwD+jWI2V4/MqtHG0BJbjyVCnOTfUlWuQZ5NO2rTh
TKKd2/+wP5qt5zI344NOCL6acXkKNzOQlfd58GX0DQwPdZ8jXYozeTm5sPeBlYah
kmKOhezeyzGsIO+5qkP8l+buFzYPhGh0ypY9jxVhPI4d9DWC++pCzRKo5/Mh1wKE
79Hv778OIUyeuGpP9Hb3RFtkbjPIXwibQfhJeMQKPOWm8qGuuCE2S+P8qK9i9pht
IhNX4xjSytUnvZekhTG6SF8nrrdt94+sMAPdhEZYofeUYgxdFlEa7Ju+psemtJhx
u5tpssmBelC0mvsTx5Z40VeZRZnKJvGq86D7zIT1QJlDiTdTOBXqRKjrQ/Ta91Zt
mOihvgM0qJIGS4MAGJrkP45x3Jj09B3YqOe7VUyApnzeOlsMqBgPljnz/npemdFD
1AImWZCQojEaB0nmomq+0ybj7SL8uRXzZmJq2YDzVGudpFoerqmUfECRxRgAkeP/
k3OANUfWEacvcyItEY/f4V/NSzGzXfKtd0GYrwIq5CELmkaGsfjDb3gly427SQDn
8fc9OgbZFhO8EEloYU1bWDfxs9fxtPgdbH7D4kVHYUFE52TN3ASvdevyuNBgIkcP
b9+pLBVAe3Q0D8p8yiBFB3muMRjdMLPcr+svXdwgT/2KFAicEmQ8ll0WQOhcRMee
3OyZEL5Qdikb87AJ7kUn06G4Gma0d6NkT67J3t+mk4KBKW9eiKBuRMuSItrT4rnt
L6JoIAu2TAaKFr1d2w06UDoTDNtfWCRgk1ez/SqoojEenTvgpgFSBISLm1DH4y6Z
B6U6JqYsFtsuPVCkPxFZCoRUymb2T+dG6C7nnHjja+/pBnxXUpduiMgnTt+PcwQH
YoA1pc1iwCpNz4SnyYPVOIeCmxVGMUZT7l5kwg8ekRHROjWrSwB677+0XLvb+E2l
q5iX7rY92cJo0T2dAnVacVX1F8dHy0efHWBmWPGuBTdcEBENQa1LdxhSnariSgc1
7qeh70n6+VljaDy4RofjHUETaWJY2uqzZ1MhCbNWfcY7XF/W0bUz6H+nuEI8Szj5
c/jSkTbNqpQpBd/SlB6TUFBGTNphMl4Ck5aX8SgOEk2iRzwc+ueQRmE92zAb3eWk
IzvPY6fVE7fV4oeQTdlam1B6Kma3iVPmnZ8qMwHVIMblVYYAV4nIzUZArTRtQOcV
ISeliVUb/WKKObb6g81LbaGf0PCtv7nHOwAZJwJHuyKzAvUkLBD82+OSnrOfBT81
2xU4oNp5aqK2Cr0tWbx6DASe5Grld3Pp8MgKlND8JuHTd5WmcpY+35wPTly64YhY
keNzXx/LChj0iEVJWGt4v1O3yyLLqhK35SAErH0CqpJzzLG2I8ZrqIfm5XIHqO1r
5KCNqN1mEQZ+c+lwu1yQH5WCCpgDHPEN5yO9xRsXjYhKq21WsDlKnT8XAab/tEAM
inEyI45tL1hzzFWyKO4qg+ZNfOuIgdx45XEusKZC0xjD2j3kJ/G/EToTN8b0dGxD
T2B/Sb9vkAHxvhhX/MPjjuV5UO9liQJP1PHW8fnXAEDn54AFu5yIT3q35xvSc5i2
bFZQhfkf64Exrn1+GVXmShKJOEiEbgkEBQnXL0HNTm8zfChagzcZxQapcJ+x1Kh2
JedUTia0dv9IGXY5prgncAPlKxeTy3Kx7VxnY8Q7K3LAzg036Nkzx0UZ3Qp0UEm5
GUHlu6pRK4FkXmNZKcmbyg4B1W5VIPp3b2NtlymryVrFRN6sgnIsgV/R8KRV1JmY
GdFnvqsDW+In1eFUjmbH9rf/Zl5QjgvN709WMobDx1pkr9DGVKQ620Fykh7n1iGN
68WnI6Gqjtr4IE5FidaQoKLnMM/V3B5uSP1jaHT37VyPdNoWIG4OWMapU4DdR4Bj
+AyKliMM5uzYnawWmAnm7uUX5gbnQ7TRQYra5/sGVpLHgoxTAkJLrSW1JOFJcL1B
TLCctkPfR8v5L+JhPPtQnPEHC5c2GDHZmSkbMyREQGfE411yn5GmiIpbqgiLZQmI
InqgsslCfi2Zy8IlKYXf+qK93wXZiHPQ8MjWpIG6HUukKjBHeBusfmZgKNRFIu79
nyfs1FDjTta38SziWJQuMAR0Hq8FXDj7TMNhhL8ghhbteW5WXlz15inGVgRVEF9A
j6YlA/CgBfTI9lf1vJksJQF8Cyh2I/V7khxiVMctS1ibFDAL8EtA216ymOa+LviU
crSHvTsa5fjBGRXVQJK5wlvBTa9+K7Ev0Mk/NUeJL6LfoIkXRoK1P/aJR//NQATq
h0q2X8AKbFDffCuyPanHqSYsu1jjrYCpX4OEtUz5EYS2wz9g8MUQUpuaIxXxjbro
W/MoAQp7sbPTK63Q/6JVQoFTxjiGTqMz9yPAfetFmYF/b9vohgaL0VLlfz8cw+Uk
uMWxKsVJDM/ZR/EgEhF8NZZtsD7xyldXogCMnBiKBjp8GGOvjxZjPbErWat9M7D1
YIUNfalU0/DyxS4rhjQv9Q4CEcb4XhRMjnlcFGXxdrFyAjtR7oyMs1b15h0+nNxD
fxbcKyTb98lAkOvxqgBtyjEMzO+pnulrC1OuvLkdVjz+2rdvxm91q/ns4mKz2hO4
JkQbhLE7DMPgtIUlvyEehs8TdzTwYm3jgdNn/J+fboiuq3djK75IiiVMjjbEthG+
0DCqd9Fz1SoJ6s1oWUc5HJARd6Ic1XzcoP/jbmo66sfvaijNQgo+9maQPmsf3TC9
D4mb9OHoxpu82P8ixO0tIFvL9UUSZfnTGuII2ngLnh4YGAmZIOnwn8U5tvLz2HsO
5M2kzyI+/6Ydc9V6vNiVgji99Rjbu3bshohVHPQvsabsp1cui1CAi0eXnro3KLkH
wek44N706Xn9/g74F/HKqj+2QvgijNFWY0q8BsoWzoLIBSokcD7lW6qz3TipTjqO
fJOQlmZ2nr/xH6oLO5qxbjq0btPrM3b6pevPKT8Da2VEVt88iQYqePZ3/9SKtSaf
+2QOQB9s7Q0f1fyrDjOBAFxTNChaoIz5emWCtI998y/TuRNkUh6cxzNn3Ai7b9e2
QX4WTAIFroaVLINBhYKGLdLf3jWuVjyJN0cWbuRtCw+EeG4iqtA9+9Qtu/IGaW6Y
WNOW34LrmnHtXnCADBaWRSEsagRwBa97B6PAFYwLEOM2vPvO6+VqhOWBs8aFm3eQ
VDgklx1wIdyUepn6P0ijJKqH4PmJwV5SZOxLAafEyLX8m0dIJkcmBvirhVOWNivE
LpzaTGBUXKzHrQcTWEvhcHzUZqIq2DQqEyJ/FzIFOWqznM37gYF7OBit+Oqm65Pc
BBQpiZYYeoSh/Zb0x0bf/zEFcpBqjDsXL3nqaRmZ8bPeVPR/mAj8A/u/+FNOWagi
j+XPX1To9kGpmbeiI5hkzJMF5h5sW9GG3c1aoyoa/jq6JNad7cnsfpX/a6RuTvuj
nEYZkJ4tlTpP1m+NoMyO2ix0lpR8CVltu1OCF+ZrvvuDd9qoWMsE7MLF1suuGVnp
2P4Cehn/bC1t0bZTfRgd3bC5r1bxHgrFYmjrfIIwEiF59Q41A/IgKed7A3DI58rj
i9cE/qRLVF3ZJRTshqf81y5qIUrr2pTz+/cuBrqTXBlwe6jOoiZYOQFzM/m6QGmO
+E/jlJ96iuigwR/1yWEbK2GLdCb+xq4Tqi0MRQeZLLjSP+jvLpyl3C4J7WZXWmZt
HI7XfUw8iTNX6LT5qT7c6MwXOdzNNE+VVU/yasq5T/cxvPjA90vanhQSk1EIuG0E
+ZiC95G5X03dHD3OWuxRLaB/cXblm7hsmNo1XhtrP05pd4S2teFGd1tUq0/S5Zu6
toT+tZHrr/cfx8qz0Y9h51cNFggV1TNFljJ96+F5nEbggpPx1IYhKwpLkuOR9rtq
pViCjsvty+Hlz+p11FrozuPdfVtXjjLveFqpl+UKXVYiRUnRMngvMrt60Mm30GL0
2vMSyZwcJk6boOZIZrJ7QGuqhfIasWFSEjX0WP3QOmrhu8nCsjCDgSuBB7B4wM69
Zy3mkodph2vZkrzSiqj8PaKAty5AcvmbDi5uDsdWWmnYWGBeAZqLyecHoYAGz1oF
zdzXIBqYvxHjLyBeDVseDQmVrDc2G9PMfsbNorPVcMTkYZ79lS6BrQOSF1OPYOcn
gdiIg9USsTKWWrK93Sxt5ng46cTmothRQYe/snzEHpKFsbug/5m9o0XigRLod0s2
ieUv6VXY/KIt4d4xDPKy8dtgDUDilb5k5zzHorxYWWCX6zm/WK/PvX2HzyqIEClo
li9ptGnxSG6W8m9aS5FgjScHbiupS7woQI47jRPdEN0qZ8Nph6q6gQ3DtM4sg5Ec
XUjhKbFmns+GELq+xfOvSNReOPGtLom/lug+VKEiXKyQcOtyrtYo5vulwSApptMz
rsJyPElZSL9gRUJ9lyKcMwdTHM0JUEdon1H4SElqDSiBv5NU3H562E+9eFfqe645
PwrqABJUwtJ9GkeCFNFLpXE4LoULg/iTjJaFaCGH6FSTBpl7VerOmhoZySNWysSS
S8swbacGJkupyf7wGCSQB7ESNL28RKCsA6rZPUkNS7/pYGw2ektVSjyOTqJoyTh3
ly2IJ1d1zXlYl0UWfBhAyBxJ5Gv7J1pNvTg3tXOZ7gPyOR3TO9oexTnbzHuaoZrv
RFkwWeuL0PJP+NIIZ5o2wHT9LRxHmzi/mvDx0RKIDUznm4p3hOdBXZ00/6HFQvHp
n9F6bicUyDtPoT++BYs5wP6cnIuPho+BDYDJ5zxmRRKpXggIwEMxwIBjNNumExb6
5dlo+BTX/T1uGmS1b+QWcTausftZnUk47BK3b//te8uzn/68q8Lu2vrAFSlujmL3
ynJ91MYWTC97vUr7CLP7439ccq0tOEKeVNfdQgTSEST3RahjnunRn7xBg0MbLTAI
yL0IpC+llw+Vz6FxHS4h9fuH+yCvUFuMTJfBgOrOYpQpvr06W4DphstRxRbjsgKr
q23JBk6KK77d2J1a7RVkVSHHGyZwytZBsLoNWmD54Dvu68VDCoROV3cMWSY72xP7
abtr/QUIWwyPU7ZYtgR7tkMgFPcDSs5/ExPGrE7hZbc/WhghfnD8vsZRSmj2mFI4
lf0oMetee6aPuPTVFCa9492433HXcuitzXLbyodx4PtANl4lpVxIK/rkSdVMqNGk
dzncEeA3fD+RmRFCEGBV9XqW1Bygq14mhPFm5BMzETxJXTeOJwB4y0pYRcDLdAVw
x4c307IJEEgIanYqJOyc8TfL2HEmmBFlAS8p2fC9zYPeuzynurPNJciv33pgsc5T
JEceLL8usYjG72WF40EmYsfuQxiv01q52Lmmbz6PfvsDnjbmlSwtGYuXqpuElSxp
L2Xb6J7zcTco/Lkidb3gecL2aPISgB2F2yZ+U+Df9giuiGb+aTpJZWKoB97tm/mF
0V5UjaOPsHR4F8S+aPnntcOTU2YlJCjQZdfBYTpJ+rImGn0Sk4n9EQgQ5gkmlYuW
uW5SXf6Iyx8SKBrlKVtmbf569ZJ8jHvemiIMuY+aHu/Vf+sflgdngP7JacHWbNNV
xtFvRQ08NrVgxkA+hdIRjDH6lsiTZklQc3FFSp+WeV2uto9c7lgEHfGhaH0+RXFA
eg7ISHIgyJbM0eI/IgcZyk2zTG4nk5LFlFSkP5HZzafWc3OzmiC1Ilro13BI7zFK
Aw/EL2jYWsj9RUX98ZmqTeQxKdTULg9818e83ILGu65frVHJqwX63bgEjXWDbGC2
lOz9HsCgRlld0XwkUOaXpA9sb8N4gFE1Li5b0hOPJNxn2Bfggi+e4Sh+gsFoU3Mp
/huhPrH+3UcUK15R/2KvKp7UjiyyffQt+eo5vCYgt8hK4CP2+/WLwwMpmaDj0lQn
YvZGImbE7LQ0B4Y2uZJRiQTOvwU0H42NtJWnaPbQCJoKohsC0H3mHrC32TLzliBK
Maxt068exEs83ig3B8t9i0ErjGNqDaLf5zdH4BXuJeXSpfVZ6upZpPDc5oCrWnqX
e23r8RZiZLJ/eld2k4B5IHf5ttwJ8tAtckHff+j4bY1b4uvlVGob6f5SJeS8VMXt
KbtbM8BNaa9I/0FpjSTUB6ggm/V+hpf+uJL+KcjRtJyv1eMYQ8/X3VwqnlLzqsY0
nVY1k+GPElzAXusz7z3Hh1qMNwb192nWnO9Njno4ggLZyQp07cz7EPmgmMHWaL3I
SFX86hlOBJT3zG+YZzOJEG57cTfLR2toGK1OlTcOZhw1Ic6f+6MyryXpIulWbE/x
mnuVQhijSfV6Oo9wvKibmoxxVXuClGiU1WVC8QzBUPb9k3pQdxkudkodSzu3bnEx
sp+rok4HWMD6peymb/n159CbPsk0BSppLTkGUCaI0CVbQbM2kt2Qk1BxfTtjWTCg
Sl8lE+R5YFVb5DusB3sRhESl0qaxNKpupgX15SakAvPHutfhWZh46Xjqm+4vjHDj
MXWrfZPWmJXjzKAHzqqyCDClla/Z7idOB/DMWrDZ9z1e8NdDixRtt5+VqicdHmgY
EulptZS1tj7WYKcR+TRhm69U2OmdZTyIAPPreJ9nYngk5upBcvJK7yHKsKSPgUlg
L8pkgZjBNV3YZfQcnrHuzibr+UR7BxmIedaHGKHjwFuKroAXzg5m7dr8PW0rodAp
uQHu7IGtRZRiB4ZoLBWkssEf0eMopnHtTL52DBRV043qZ7HXl0R6ozByQbgibvf8
XlLwMZvE9h0afSOja4KOUmgfsrqxUeLK3nejAGzbZ4y6s9bAyWvmEgzRTChUXOQ/
OaBuv2rF8OiRKuPXh9VIsQ56NDr9kxtvWLUvDjDWtoKIF10YjJdoAnDK6mde5TrT
OdN9a1MMnOcc96qGmktTa+I9420KLr5trVHI4S4KCM4LXf9ukiGza2x1QmRogjHW
QPLeVdKYkf5jRCFqD57EJfhs04+5dl6h/2zzlXpv9BQ5FkzoJ3E0V4FgFBKWzOv3
FfKZvFyFn6U40lstGUAkNFFcWW4QufSvVhiCiB/US6OlsmzA7d544+XEkq5tZJ14
HZqRci83U+ekmAAwU/zDLM9Sk8tMuMiga6bmw8JVqZbm80TqDJaxiybCoM/+j+xR
fGt9RWOCllMohZPSBwlEEuYZgDCJTojA6/zCyv2IRBjX8ZN8ylN3FLO/7vLqrccU
CkFay3p12uKXKdDzH6osUT3Prdz68Mw4fuuVez/HJFegJpaqqO4znDMfpVE2BwAU
g2mlHzIt0VmTA3DutvJl6qlqlQYbptRqYgjkrj/7ihODga1e7iiCvZiqvFHQV/6D
bvLqRZfPOewUfOlh5cvVvc47GZjig3Kuslma7m7kK0hlBN7nHNEpXsl6unF962Iw
ZjYE9meAeJHvo9UEW/yjy0QtvH8sY6fb8g5MDmzGYCqVGyZrzgdkkS1wfhlXTVE2
3KTnheXIzgoy9qRf/jaN37a8RE52zkhTt8fPTAsDKJa3Rnd6HvGOPuMbEmPXXR6Y
GFQhLweONx5FzKb1YFzab/l/ohKMb2dGmxDVAPkkBOtWVz3rliclaLDXYXpOmWdE
7c4t2b17OugZXr5Mj54/Qvc9SlNqq41vzzSj+DaDW1wSx6X2mKIZwmhUIntX6Noy
4QL9yh6tjDoOE9VTB4wEuYcNUHEVgeJLqDXj2b/gG5fG3Jszag8FzmmiXa/y7KtE
ZZw9aWgUMTcmTbqqf2omMrQ796SmZNGgWP50SPX9x3qOyQwWV3AmR50WVIBvyBt9
F0SMBO4Q+66mye0MevaL6hXGYmli675l10ZZ6k+VsQaJBzbi+HcQkKV7E8BLJlHy
7YHdQ5aL339n8FDWLGEqCoZivsbW/QpiA8yHOR0rRPFMHH8QssPt6JAxSuEVbOJ3
KOF8vfE6I50QDn03drvX98yw0V0XpaLX/Tfg0pLEYCuJBDPwKq2f31PfeG4xO9ek
qk8oWpixbwymt+ik199J3YTGilSxe3uP7HXTHbeYcPfDk0R7S8Gz9/yBFE499ICA
O9tvihB/BSSjlMnQsK7O++esQkdPkwM5nkvQD4C0tLAg96NNgVmVk994L65tIRql
93fhVseNTDBVZGoaMs8DJJ2YtxWeRnXzoJr0hO+zfIQ6wAHLvVtBGPLMUJtZZqvI
1eEBJovut0WuXYDFwubNrPYzlFoXENl+m+EvJasJy1AD49naLdahRIC4IZwKt1O6
BjmFZ0rsgE2mkSdIxPAqpmVyTM0mZDr1+NrDr/aCE92ORAvbEARPuUU+r1p1csHh
eeteI2gFQoDDSG2dGQn6DN813H5FmrECA9AvKDuWFmlhV6MGBW6aosfJXIUxkwqI
R3a9M8wbl2/cPPd9Do03I+mhhefakVUmrRE17et9TpStu0N7vl+2ELXhZidUbx5D
6JskvGNctv/2HxfoCAib7TiYK6sS2Hfz4gKF3KI7p9u48IHI6im3xv5c449GLdLe
Z8N+4n2L4oMb+PK4HvxrglACkXD30cmz6F556d/LPVPYhPmJ+niHzg5mO5fGAe4G
muxsuwgoKc/Uwk2+Xwlc5qO/4Z/h2JMyFAYm28FIL2j3/2354kf/eTezTUH5GdPl
3Us1X8BMGFd5PnRxSwngOrTss/znAdjYgT41PObcCZlLF1brxK5bEIo+RxsXv+6N
AkabgyIlGhuBLnuYs7B75Mg71g/Bu/u0UZY8urNVbaRPkMmp/drsgot20ggOKC4A
KD7Zu/g9kvwK7Y6KlmUU/QMgO6ASADvWg3KuzYd0aLHcgw9amcqRcnH2UTFUsFWn
uBfRjsdcXJYTnSAm4l3fYKvSSiqoORTOHri53ipCe6WQvIi9hcgXDQ+OOMRAiiqs
rt223JVz4ZWiJyjZC/3HtVhBj8peu3ZW2++hoATy+Tr+R6jmPyvIkL+CrYCtmvT+
Ixn0aNiBfH+WbFyK8r8r5URb0Ej1ucGx9KqCOuh+6cTATJVWBmoa+rRMb8sq4LZM
uuRF5y1VX8o33MKA6oXo7NKWDVVvR9FYoSQxFZxpfzP7KJlN9mCGB/23/p+JIANC
Qgks65m0QIMVfWFQEvebkGvMcG5iNGFVmmVEHcINFbRgRwI3RB2AznTViR+ZO7Qv
gBJnNfkPoIT+WO2AmJsypRrVm21d+Nsp9QhE2GZ7S7gSIlfs+yG9hg6mAZz7GxuR
M7DDMvR2HQRI0WaJppvBgOjVKUC4ylcCLDtWTN6uZvNfn5GXcQl4X/MeAoV/j8MM
2BXbUcOo7Z+G8p7A9/6BwL5WOSMeomnutDQT1vrfPMCy9i1mmXWtDi71tUVW14QK
VfDM/1TtKzQdxFFaLmFx+NRgfdqOIbMt8I4FOr1leIvZ3JSmyEZLV5zS53UF7yAA
sRwBmot1OJrBeNg8Zfv7J+4dSR58tm+NYFoIbvfLBbX6330quAUPalQlCeTyWI5J
s2seSIQjJrIdX3iMQ92Qz1CEdr6YFLit6R4zrIKs8ut0fVR8+wJsKX/v1HmnYPyQ
lVJ/RocwL/5iMPhLXvDplU3I0dfaz4E88SKbLZm4+6UEc68sN9JaPc4LAJO9pP5d
9hf9yAF6i7kb6LL3i7SsIWciE4AOQhxoDbnMTPfjyG0eaG0wj+3DPtGg24U60M9q
Q6oIGfhG7b1kfnXHpmaygQr2wR7boMv9NtcilJGBaRSBI4rvz3g78oxM+yKIy1dG
6cQ+6WEQnXCS1nwtGv9hhIV14yf7Q9qS0QFrf50bZoXZn7ydEEro6G+N5yqj8cDn
EvKZMWSfjo5ME8GBzSTMXIlGnIliLXa3Cv82F92oyoIK/rdIPb9qf5v+SXizwqiD
PdTcDdFuwChalwMxNyzlGZAuHdLpt9R9hDRlz1M7DZT4EFn/ArwEFDaXMv4lVQMz
R0i+oXK4W10hWtcrltvEosymqSPq0FVCxt3jAJybjpgKIBarhXLgSQZZGvluAB0n
v6CIeO0WJXAwxXJtxTopyqz8eYWdvgMMLtKtIbFDUsLZVwbg1JiyXDJhR/KxiWYG
PzSQSS4TTU8bUyE5NA1gX92WfyVJqwXsza+eNnFRtJSA/EUQ/71GnmIKy7rt1dlm
27h34BmYdiq5H3FO/uUWIELLgnRL3Sr3y6TjExjdBDcfLGML58j+aVbiFpFcgbjS
UUQ37AK0ttC+d2ZZ2Zdx2vkoRolD81uY13FH9JxacqoI58iVD+LNe4CS/NVTCXuX
OmpTRhVr5oMIm1eZ+rE9UagTxn76VkaCVtJbo+0jfPUoYa3TOD2rr6wdKG5iqMzn
Ppq1fwL5yoFEwg1LnnF7AdMv1CtJvFVyF6wdxr1qemfB0s+TNU++C2lqTetBYSHs
0/8u6qug/8qOjesACfRYGvFuKk9VNDAZR/q69mT/IOM/PqEa0mal7XoEAMYT9k9C
YP7ARWP98D2ZqBLe5ksTy37l2CPk1e3t1jVDxY2P4YqyVfWY6xWcLh8wwUUp+Ci7
MVTzcqpJod+0NjuACsS+Bzw46ePHsiPOjVGcjOnliIuqlgnLgcrqal74ibRuKf8q
WZfzd2vgOYys4pZOtkqtUa5dnhL7VpjZd9MYZTH0GsUS1MahoA/NwVYazfjlt3KD
qiI/p/8qd8hKSW46qimIX9woyxpAH2Vp/6yUbFoppQvT0fWL7w3j9hwY99/Kc7G2
pevGbwWv1jKJkp1YW7Un1AWTfWPO2xr5FfhztrlQbS7t28ik4KL/aIebbVPjD4DL
TN7+xuXakc8FpE86lzg0esTlTJmyQxaP1tFT4ZcctD6YmIpc0FFw1cvGltoXviv3
Fz9YFMdPqrJ+K3/77aF9Y+t2tpuM4hRwri03typ6nMRArIqPKYbZcqXJGEYuQdaU
iabbQq34VinUbxeXD/Rta1oot8wQdmHPbK2PMtxpTjMZ8yZbZv/2y0o9uoTYCYvj
VIV6MTyM6AvKZcQ/nBQjq150EbmQukg22kywV7cXzd1ywo8UD95mSdlAZWOaJdS0
U/htatGNqL8jM0n7MRjS3da8bpQlyPr5IcuzblkY2GNUvw+5HO1bJv0wb4FlBzqi
YNbGnZUNbQOhf9bzc24BeHDnSTZDKAxsXp7B7Yo0bqTOOWRLZi3/77sSNzPqjZIX
YRK4SKesRhRb8T7DfzshqR6B4+A3xYnTdqQ+4E5v4kD7sW9D3oQAc7TyTw+KTU5P
A2PyU79XGj2vQ6urVYlZkMwBiCePWyi+dOxpgBeRwyYXaNw345ZN/94On8eRESN/
vBn80/Myvr7FPNOKyMGKBaip/W2Ms/lHO1YTu1/KQqiCDX7TLAWqvM3SbULbjjhq
RVaO3QRu66V7RzruMJQwiXOEYJBDb+yTmQpNjlZoSYSSWhiEPdxGaMWqbiEGAqWh
sLAw82RxYfldfodrFI5PLrJPvF+C2S4q6mbcmqEJDd8a1rOBeAkvEknvjrGHRUtA
ut+0D+/z8Q0Zg6b6v4iQN/oC5ZwAyCsRT+O47XLTmMLyHaZ8lAzP88LN9ZMtfjVS
UQw2DFqMysxQ/w8kzFCq/eBPv5wykBOAl47cXOkAY4RnHdXoKDwE0OwTlP+LiMCC
CdaXJoxxS1j2YzfKOZ+16cPCFRC74lySxCYlg2TupW8GB0JhYbECv7E+EGP7hzQZ
kq/NRysMdLH9D+vzecNpUqn9kjmTJQLyRYd3hPQMotj768jQeFtfRhMf77b1aPg9
aWLL4WbIaqhK+ARkW7vFsuvbA5jde+wVhu16Si7ct+a3kUhHrJjTaHmTDyiQ/XSf
oZRlctDCcX85JgKT0VOCCyPRcGRiNHhIYvtpiXQefAG02q6as9LResgtTZh1nHvC
zIKbTzUQpopqCdgOj5YSPJsPvs2dOQTeppgneLARpHmNoOG8mJSnFOpr9eV3pcCQ
F2yF08QaoJiBSyn1jm8T3nTQiw/7Gjy3pC2/5ZZP+X/ooCMPgryPqe/3ePx8rwSf
nUoVvDmkMah2FGvHEqBnfc4lTlVy5nJlv9u4jsJ7LLSj8zJpeTgYL3JdT0fxyT0V
c235IjvgyP22+jzZkg1nCJLPB9lZmtioj6lB9CAZjjJxviv7Ze+yTvzs4HEoHApY
BiyXLLfYjJQdogWKdmFweDH7mk9Mo5E7MCvbuicP4gaoRzXl3zP3oZcRi3UJ82Wp
ux3qj6XScbbHBn1sao13Zf4fQHwxJHi7ys08GdZW45efDNf+pZCsS7ggc6hJsfKF
lJCvZvefUrc8UJCGTHdRARo0/WtWjSy2a0/HsnYQSRvx9AOn+4Prq2QjIo5SWkkC
14E35l/0WRttyL/XJf1547UOaQQ8Y9oURKEnrgwZX+AayrE72ddipGTvseCrVRTs
ky5rW/7F/gJM1ZGv3lfshnO4lvM4xpB1+4LlczjuR53udU72otn27Z8Xi2MFFuDp
F8nbhd2NHuP12MNxytJoP4cQE1RCIKtOu60TA7lFymwV7W2ERpSa/LpzbuVuK3jz
9uUTglsxWnMz1Qhm/HdLHCJVKKmMSK4pjyqSYS7cHNIirVHzlX48JB1zCcGy3moY
gOEY/5zcbY12UesVnpYvHhYzpbJgfUn2AUf6417srF3tpBrPk1rF5sj+6UC9DMO2
bGUOdMIpEGM91JI9VDnG+NWmxlIyMA0zOc4F37kZfbsIfbn59UJaSTOrx1CXafoo
qy0S6ZBPhmXasKrGR82uAE1yi1Uq8m9H7q5fywkNfuGi9HtPTfFV5jILMo2tqDVM
E9JkQBG5MYD6OAjKLwtXftNOsIWY7Sh0uI3Bim8d9da2JlsfVB9PFZCSdcXkLjAb
Ee2f/OUB8a37p1RDHQ5FlxHw7auq+xCTAW02n2WqdF2zuynHsrD7sSPRAy5GDDYO
3UzQl7A8/H++Q4SlLYWQf9uL+wzPUt9IoZ3YUmF8k2mBnLPGMaaICTxoyz6FscKu
3DoMcO5RKJqO4GUpKYnkciVf2hOvDVhBJiQVI6i/YURdvYX8ZP+wqUc8Ctdv/4cz
buI1bwHMQUX5XlIGnFd4j1Kc5cPSTFIqC3RnbR2QuVDb8SBb+nzt1FssSIDlfm9+
FeqbPBKAwhOqou1xMym0AaCAGWAgJ5tgkTIO57e5xKTCh9Fs5Yy5lnoXNeQIoaIA
GyQvgyQDUcvvXusrRItUHR8MExSstdkXqM1BsOWnyEq9sFv+Sj7Yxw7usl8QawKq
Ql1uOIx6WuLOZC/U8IjSFiHAZeMKQFYSJqNkKwQTRgVyMAlzOWtc4HRRws5lY2ra
5duVADbQ7b7E3KFFieKBLrCWqE41huwUwSsv6+V6PIF8M23A9DMsVj1n8Q84RHsd
asbcSEXPoTooeat/+LGi9X8nswJbuRbA+Juz76P9WUa1PdpYYU9BIY3EON/FBhkA
G9YnqcPCribG1Ju+qcs1CaFYZd0lkXgOeEPQxdYvjiL1F3AiwKfrjxTMl7bSb6Gn
SjTWZghkk5lyTuaoKbbYtM/Fp5PoHS9zCvKW45Nbvz8vqL2yriarMyC7k1FXG5/u
lfMqpiEZRmRytGSlZQSaLvePxP7xYRXTxE00IxL2n4r3qBCIbJZQKFzRhprPRVIH
h8pEIbDESvgtF9XFr2hxANW5BYl7u/k+gTCQBmePi2/PfEwUJ0eN4jE48ypE2u86
Gblsp6LIFOBFrzPOOdGQk1iORDZ0xOZ2gSpFDWUWm0H7+KcCEBTQqsqsK3m4UK2X
2vhd8Ubg/XRn1TS6Ia00dtG9RUGUZ1DLW+V6hmwc9pBwkUf+K/ZuKQ/kWNoe8j7D
qdSIJS2yc4DMDKgK3tnUEJJ878SvPMKajbzWoXxu1XuGQiXYhSd3fPvmAZWDwqmm
h3SA7ePGTCv6F5u9Sek/m1NIS9NTr4FqRyRyE8rS3kXqYC7f7UqKVyOmA2PZV9be
Z+c+RlhzcQN1cwZZlmgmj10brbD1HWos4fEZQPug3sSgmeMWm1OU92g8VdawNurS
jXuzpBgeF6NQZIfMYiVW5AqswjxEpmF+9JMxO5OI/YccVU+0HCmtoE2EMWkrDXQ8
ZBDpyuCYPiWvj3YpUJQc8vmQYTxNnkX7adkhURRkGRzH2rFS99bBLlkfNmpr0SpN
q2Ra+4jsPBf3Y75q4PQ4rU1TUTzREJNPeYE2ipI/vhWT+6z3k9ORnbhElX/jgOep
ELV1RifpHzFokheWjsUg6x2keotLIfwecv6LjsaA10ckjVVBV75oZZVStty1Dxqr
RCIchwpsJAD2X1hD+rC/AmkaZhoD78v4iSDgyt/gK3RygQzmwDDqsx76aAk/Jtf+
eDdmzV9IABtbI65E/Nk67g0stI+ABoPSwPSos4dgzMHjcZaXXOqfe1EBzu5yhYbP
QwzADH8ogI+TW1uvreLjuumIpNltQ4knVvHR1uz4DAjb/doBxdTA9GT34NkAq2Eb
JHRqKEb839zAF3flK0SSTV6fRF2O0FFeiYZtzuV8QXGLzdohywu1Mdh8GpLAlrae
XfVb2/n1t7z6cV8PTVzhpZnG6Wx6glLvDYeSd0vs1pweq9zCFVf+m0LLLEcZYsGp
BimapDEH1qh//2Eh2ZQimR3Q6zRKW2ZbMd/2gnYkatyOuydUa++HDKlQSbGyfqO/
UZp2vGBQqHGNOG3+/8iCizgkWHQ325nfqZDb7lVsSgm3lKvXJ/SSOEHYaiCDZpIh
tM8x8Uc2lyJcIskdi4cp3B62JbpGJSCv+aA9xmAndz1TAKYrj3hOLz0juqoX5a/3
RjM0SOwL963k4zbQq1zcJyLJYoRBuzrT6HPpFQY/ymDMZvFMFw53D/KHaRe7dqGy
dPQs7PG0QRZ8h9RG+Jlp+YAt+RMo4EGrbcSyAE333Ug2kAcSA5nf1kySAXW6l+QG
Y9aFmaGd/9khf0oP70eK/0/BL76zNjbjIR5UB9Kgf7mrbS5hJEMm9dCjiyHWxCcY
5G/GYFLKlLeJyC2uN2Aztj3wO/gqlusWQEGYTnyCO9WIys63Dq8sUOlYeCcT8rUO
wV5rx7gDWUkQuU+5Ze/s93Us3esLY54vZMt/hJh9ii9T2xZlRVpKjac06ONzM0cw
in7yfOM5R4X5EqFHKiy8BPEb6gAl5r0injBvJaZ+TiY0nuK+0pbGhRTh1tfB9qb5
kUxurfWVA+bum0caH5ulWaS2pi3sLbeMQM/RA7jfzoaY89ZMTf0JILa226IdUOqd
QF7lTwclwfF7mQHpIHwpw3JrNsVxiQBU4e2sXtWT8z2Nn+5uMFaGm7gItSe2wry6
a1x0JSDpzChbjAuRcCOinBL79EcijFwg9x0t7KUYb+DKSnABCKphGmX3SXNwaR5x
qBYAT5zIviwQibzKYeDPc9O3AwbEuRNCRgZVwm+i2a6RWilYgLJ4jRCpYY7xbZGF
KIxmM9rPDwdR7HasJ6YZ7wPPjycl3Qisdb5XcYTfZ3WM1QSooJQmxZs17HQ8nr3u
VKi/R1MmexBvTSvTz7PZDdmQC6BvwupO7EhabPePfp7BTLzgfHwqXprpeJJJSVKq
nv9QDwppTlslfjN49cUOm2Hyj/zvkYjkGi6IUCFN2PUaMZxeerQb5HyIqEQw7FDb
BzXSwwBcaKfAkVpui1wXqHkE7712JvZGavOnbTvKs/WKobE7TMMGVTdaSOrX0MvF
duJRFITezjq5KlSa3lwTNG5VNPkMpLnwHtPdBK6bbp26hMhoYrEeAdnvZ/PZPEVo
6mBARCbc0VBeUXZnrM1H7aPMb6h57/LLm6rRkcywucGXifdo8P2rGE8aY+B9sULo
1mKx+frC24pvdiJV8GX0uTZtyUAdltPfA9xuPDvMwNI4ifnBfANfmK/qspXXofMm
5WrXjJRjEzvyYrle0E7YBtJ0Idm40djIJOk64XKQGSNUYBIXdEVQ/BzjoO7ZVgym
mPUS0vYUdRit5jvbr5sEQmQyD09+Ec2iXYsL7+QeuJmlBWaESZFZ0z1PzDisSD6K
M/CZZhQ/kHFPB7bIr1/hO3CuRU70MVPZEte32KeLoONw3HwGakzgw9p+biv+LHuc
j80BRzWGHaqIEITlzncyEy1XcNJkAf48ScmwDS2VrR6PVgwXbusCLg/BqT2dV3EQ
sxZZFjccB+FfaZZT7noV3xkCPTNXiicgx/fJE3KE1q+IOr+wYwTGiDoUx4LLDMi7
D7N5VyteIKYaolW13TXWnbdq5n8GS+B8x0rgMPST1wV44EmhJNAVluc8WE0FNB86
StQ9e7uX8PmIvNLt4Bq+BPg+Bc9pN88p4l+IMvKloBZnRyh2az0srLYwRfynIQyn
8x4S1aJIB8HfSncmKztQjmOy7hDx1ueAglp9yStsuXQRhNuGQHnTbhVvlg+7SBAp
hiRvZ/D7ttkTwd2uRm0LKx2n/a3cdyLeZ29CdtejMu/7JQnZ1UvngHHiSQP28Zrm
yvT1l1jPMkd+euidKxgCLDS9Ctc6AODc3N0hOXGqU3VM1s3j6bT/lCD4dbA8xkeV
yhXI4agsbTRJkEAkuFMDy8pQxHwKLSSAlmzrWDesu0WctpkHwqJnHntUX7l5MJ/s
QIy/+luNir+TVlHimq13xeEigS97M5lDBqL+NRjC4yPaQmEjYRM/GO5aDCUE6Rt/
cb96jdte7Ezn1BF+NQ9yI563z4aNIj8QyJcwFMoQAWqEfAe1buOUHAElprPaOxw1
HUjKawqMdcwCvcFiOmwugoYAb4OIBqKrTEue1pB3z9uzo+uEEejRDRSIawj+vTHv
Yi0KEzKsy2fL8bCwSJindamNAcvVrMSNikkLxUtRjiRIXpoUE58DxglkG2CdVIxQ
U2zUjcDWOwJdhSB8ps/w7N1sk+2z/eT45HT71z64RxV0B+dv0NwTMvOpGNd1WbWY
4grFUQoYgLljs1g++yu/cUvLu8maa5/G25IqYrTzpyaU7iNe7ZdI1fOYf3Gl1kvV
ps3tBOIX4sCgcKjhJ5X3CyC1GA8KU6sSRBR0AUbJrhAfyOdIkNxPEowqARvM8AtU
NpXlMHnIhXHwkrWbNC/XsLBcdGZunqYaDF8HBpNF1sf1CCOp1lCRffbspTjePSUi
ErLLVXYRPz4pE3ZysEsIdGFbQ69dv1GHyYuhQiwnarXuVFUVhbXQ5feTs2g5JAD9
GaKZnhMqXOfdYn+kP/30LyUbl+2FvKb+Gu0jd5hzRYHpGA5JNfm5DGKcwmcA0Jo1
OgN9RkgouXAFKT/OHGk1x6z/3QMdKzRvrgC6x0MUckxHlR45Lrbkric1VUZhtzbe
Wrjak65SCWty+ew2lTWJ0H6XoOG+dGeJqEJlnhVY+Gy0hw+zEVJT5zut7NNUk/PQ
VBb8/9BUvJay/i85rCiwLs+XWxeRxXeCAg4xuiemqROf9pM4a7ZBSOyq7/szFW0D
BYca8AnBs4JrxI9Pdt1iZZi/bLH92zBb4yKYZSxVk1of2qp6z7Cq0dxtPb97fRh3
ZWklcSbAc3DV6WwYw6IS+ZI4AQ3WTjZi/BXhmsvevHBd9oxClsagiydT6dsKbX6R
DKp8uXnmSyDgC1FdXgPnR8WIihmPz4S1OFqeAF0jUv5AVCmZUqiFU2psNr0Dn7QK
/kV0bFiIrdZDRo9CEPnUWhyXtIOpjNxCPRVmB1NgKVyW1KnMO59K2/da5DpdteAi
eyu5xHQ6Dhxsf69/V69EiMSPUz9xTqVuJnlONQCdreboC7US+sF/UIgQEQovgB6t
zwb+hEB3dhiIoKkXYzv+Z9O04j+or3GvUqpYfXAjBv16GidJk3mo7Vai2OAyeXl3
DkOsINd8b1oZC6m7e8pqgYDa7paNqlHnA4gfRH84nmqmfvQGL9bW6EZyNs2+CQ9e
4ZeMrHgRPTxg5bhELilxn1etj5v94sSTe6siRdw3HeDZPioqIzO4LeXU+35ghXpv
Rhs7J1P4CC6p/q8VusAw5RBq8vX+eF65QCiR1ie3TppwN/mLXsN5DIOwQVWxuOXi
5aY58oSvS6l1IgEdhV9zPB5+yBqWm7sb+HWa5uMHUeJd/WB2/nEzd5sFEikkq2tq
vT7MM+kz84orWfw0kZmVfI29R/Fd5Nk9xUZbh5CdD2N1mf6vvVq4T2/YLJp6cxS8
xy3NKh3+1Y38iwiCw36UyYcYT3KiFcdlviBiEMccA4FuJ3XDnfTzjTFzlLQVCMFm
iObsl28ohcPCOvrLtwuWrWG/oog5Q5rmig4ZHzEeb5qbYjeQYmpKbC2TQZB+JGnX
im7OqoNsFB7kzWQTvf0svYu3OY3CEFKFfFRadOIg2Dd5+ItdKZ39XfOYlV0mGgvN
U8yt9mZkYeXzidNUWkQZj6dwnv2MH7PaOKxJBwN5pyFLdMkNk66QIk+4ITpM3BUY
c2AzBqWnbQ7Mei90/IW5dsVm1XQ2mLQIGOItyQq1+fAiKGkokAHcGPxOR6Zp/3tC
/Yc25bnqNey2w3OZ4YgnjPOU8SDXGaDVucQKyfYbql0tN1JHINZIhnmGSlbKwTBD
n7+lxJPqrOfjfq235Tb8P5PUZi2ysoCbBDsbZxd4rJ7zSoZXfmnRPU8YDUkKcYQD
BNPPLpOd6NjLARXYRGTc6bd/3zgPGpx1/qHQ8leoP3WIr/upgyfBjqnsRPWb6NM5
JXuFlFQxoBlK85zQWi9wEOzRV+IFKdz3d4HFE8cqJuL9RM7cY+P3R1ssdcaJqRtB
bWe4HtmdpyZ88HtH1c2OIrWqUMEeBe+lyyDQMI8FdvjynKU+iUJqGznlI5pr4a/Z
a0RGUlXhoGw4/U45QWQvuhXrfs5fB3FRxmDxvO/UVhce964zki5yMJNHnSoLvI+E
rI6tMgHYSY48iUkF9dx5lbNV8M0UtRAy7zr+LsYmG7dM/cXwv2LVw1HHd5tGs2CZ
bvFo+GZYsGBi2dBhDvyJAeADaG3KAVeZwXIHzEcPw0ZJN40B2t7VnPy8Z/9DzIk7
ARdj9otiR8OWV0JaZnG0E4cwgdToxLZNcyk53pPv6FABYHM4R6ze/U1xubPeOB+o
G1vy20/M5mVFkE9Q+Y0rxgH08zK+gkWKyi1u1rRXrjps8dDVhe8JuaBUf9AN9pcx
3PAyCKHNQ3Bri1a7LuqvnbhzYIfFicWl61WFLK/O999QqSFzeLtBT6jZPFPNjxQl
Q0VDFb5Ka5DUmKRBuWaGZejqMBaYImtUciKhhTaS5tjw5SK/vM0lBFHv4yD2GWMJ
NpFk7bh8k96+RoKWGnSPKoJBKs5aac+Hv3Hu0KBTgknOA3lMNo1XqH8Eag5MNQs1
iPJOcbkUEaLtTEcYkK8L2y+qfvSN1QsiKw5iurvx7FCup0pEycBfbYgP/3OCKu7C
qUAO0AgEGr57XiIb7PgL3MJsA2M0o1dXSLWoI5VYzIQZhMSRsNL+GRAERen6PQpv
LqY+JHhUGIExtiHMF8hbt6UE7MWK9U4CwVL6YIWak2oTrd6uxc/WMKjUof3DjZRF
lSx1OPYhKrSQJXZyswaudlKo3WaauF08Lq6ONjbS99rymvOmAu0aoz/2S7L1QGCH
iQMpDbScc0nw0eQAddVy8wjuZQVQwYejozuBZCs13zir0yQwoAp7LN1bE/hQbKMl
E46Z2UBV+BLGSFoV1qIm3FmGr63h6U78aw1wTl5+F4400jwfeK/J5jqPq1z/rHUf
hTCDhINCGNpfRDEW64WKZlH/abZ2NffPTJaA9Dtuy/mwnh/aa9VtU+FdOKSMa0UP
v85rrKPVeZg2LJmLN9IwqW/XBrE8I8TaQFpHDVFI5sBy68w6TN3KRXvhO2zal/m+
jZw3CwTl3clSgi5wqg4oSPuzlKB0fbTz3n1K0z4ZDw0YrkslSPJKDwXvf2mmz9t9
BVZZuzCcPQF0GbsFJNgzwzGybjkqo4h366nqESueu+NlQk27oV52zgZv7XYQCR7l
Tkq8VN9tZzW9ReTMUuDmGxwm/S7OTdNHdkl+mNXomEJTTPj3OsIPHhOmEVBaAjFK
yihv6QcoTZVvMJ9zmERSXX16XuCxDJHq2bIds4hkC5kobdh303diLU2ayVH2kNKX
WFvPoDVV50LkiP9YaicKUFwE6KziLHLnbuptkqszeNG6yy5xyP1gFjzEe8sfA3XJ
8v0gTcYCl5fYJ3i5J20ehDToYL6HGbo0Fszw7eTcuQ+zu+LFhfTdK1GKFg+tSBLR
bz+FCquT3Er/rqzkMdLzIKyCIy8t+/n+QuCa1uWblXu2y0b7Eq6CBqHRpGPfenax
qMtjSKI0/BtXDNLY7eTjceaGEwZZKAxl4qtAPLBsaaEryW1XgFWEbSSUOkJv807F
tBRI4V9LOVrrvSHQ6WZXNMK8wIZz5yQGOAtpPfKT/RLOtI3TIGeU9pCM1qOJNARF
Qu6Z9eSKU+Vjq3AD/FqYnN2DmLeNxwHhrnkL9iBbn6UCdcLccc5q61w0Q9pJ0bPj
jiebyxogMP7yJ5BpHb36wL0oz5vLITym9PSL82rkavs2c8I52Bl2whkpuXTMEh5Q
y6uD5ZYR51IZemrIKmCOpdpRGB1v6nz9rDVQCw1bCs8YdmDPjNQ2S9q1n5xo/m7H
3MxhQoWkgSiDdWBSerQ5AzlshEw36R/kOMCFEsQe7qnQYsj99qjUZOhFIcb/oFfr
5PrAgnFjv2P2NBe7NV1ZFfZ4BMaO+oHDJ8QJxJrkMQp+Oto6BhhyKOHD5rtosTbI
uMytkYTy7ZTOl0F9OnB4qDJyCevQ0qwK9WvFsNJZU6Gx3vR9q406S8F6ddevT+8e
UHEcBzQx2p9FBRHcSt8mnN3mraY2dhqLunB0rMKVmxXTIbfz6u9WWFnExyP8YnzB
ilxfphk1rV6jzluBzi3+ddXtiJkmlfyj9nSOaUlKSquZH8rHBcOkG2DgUjbKKwzK
rTMy/GaDanwurM/nxgbbuXli13Xm9SNnAkCN7cujj9C7zHrO2hgdhzfsnYUVODFC
aFR9vwTR/IWznXK2hsQa3aoDb/cW2hAyxId2OyI9+ahdNqmNFj2zvULC08Q9d7cP
FXbWRWK8wb/SfoX+0cT9q5w46D/qYseYw0Ee8URG0OnDYJcOXBFlBKIzc38KVxJ3
zvLGxJJBOAsyrljqSe6DbcvxATrlc2i1KIpuW9Dy0dqbNVCLR/uLWvNB+iFspdlT
/QRrHig1tc0JtjfqmbXv7OtCT0d3tOIOa/HDSjdNgRVrXwiErP7k5/oKwJSd297r
mECT/PrSn1Wu+DZZIaN5jR5hf1X8m7KQk+JQ1KMPJfqxUBQoY7zKTSi/AOKBbYie
dsMGULopPYJZQRpb6kRvm1uadyG7BWH3f7tC8VXu1oNLhMQmGu2W/5fK9BtIz14o
9lVbmjlprFML8noF9gwfiqzdCnPuVlxBzmGUWj/FQmdGh21jDcOnC0vMj6jsAZ/h
pzmakknC/2eAwHOeJ0tjcMRqd9pmeKbuLsf0a0TekfuHsigo4nrNhHXR6iZaBDhV
3W9NB1C1nw9Xg4TDpxCyCheF9fDfxvi7vhOHrksEnO5wv/81n7PUgnPEBFfuFEq1
ESA3S4KJ/+LI25FFsBnHToxFIVvG+my9YuPQM7VFXcaM28UfzN3Qi0vbYN7J7yZH
hCr6ihGSSdEikgPSglYrFanVAaLmjsmms/xAlTfbNCFCpsqA6JCCSIjMhiYRPUKV
4f8Tr2WacqfFXk88KETobBvQ+o470NzPTyIyyjTJN7nwzuvvyiUxrzUAUFJiyJUR
nekaXbLygDJy56wb+y5q+98tsbxZ29Z5kgQu3cktcuFJBDcygVFNXGzxdtj8Zn1M
/rgFJIQ3wZOOVlf23HUtM6j3yfkN/pGVdJx7JX0I5+PqZdrCY7nvMARMaJTb5hFM
xcps/a++KtpE0jsaA8kFuShKJqmeP9H/1m5brKXw9xJgzkYo4sHtwMQR4GhjvQQL
I0MicN93U4t55YI7lDgvbMMjkgRB/8US+MXvDaKDi4m4a/mOuFhJQOnKUAVpv8TZ
osknrRZmVk44Jee1ZwCiGOlwRLgbsTC9nZgPV+Hu89asgmsFV1PV85oX7rZ0Tath
I2F3SXj2iinw2XvsnxCMYAReAzvIKhXZXVHhPuSB/Bf1LJo8/lyd2v++ZQuvBoN0
v/nAlkFJQb1vuEsdIQoxXx6/dEXYr2Y3XuT1X1g4aFvpekVQBmHksePubjHtP0Bh
vOcRguOYak8ExsnkPI5o37QIbWu7B5WJbcOWtHDxYPo6q5XdhNXFNFjupsgKgxnU
AY0sFpahV4DJo6hiruAeR6xtJsP7lGF5sft8jdSrfM71H6skMkXvMgB/PpJIECLy
O/Hns5xVYI6gYxsIxtpTR9WLo/lHJoAluEwX2FOEWeNQYu3GtxcyA/UxAD0H/MuD
G4uoaseJiJGPwIeu/RQTERUkoD8YkzwsT6FRXflSVr7vrTHaximGs0d5PKV6/+kY
AJv/eMqWsw+QUOhfdU2yeRclwi+f0PZNagsfnumk3Y/UCgoadI2Xn7R7Otei7v5J
raFZuW99L22e6/4Tgel//WoQv3rb/9bnuRGtkCiqzITPlB0A48B1+BtXMrDpal8y
vupEOyDqqq4ox2VjvefUvVXeaguiy+chDcNRI4tXiBzKNtBz+2Uh30Tx7F3TT24t
nJHfg06CQgod01Xl5NXE5AKJr9RzilpEebtaZqT/pUiQ+QlX/xUxjbwXfrVbp7OG
5GdsYPGY5vMl3mw27Glkc+ambPMzKB2npjPzGptqr9hFsAY7tCWgX88P8mdu7i6c
qu7I1jooWnj0HowQHQg29Nwi/fKvtSA012b8B1Tk5AJnzF/+oaf64rNpbvFiKJht
/EUaQ/jK0MKLC+vrKti1sYMMBQxrupvTpI9aS3QQE1TSmx9JXHtsZLJqut71DzZy
+cbeD0xejIfNd2Jwj78S7hXWuuZ4DUBByre4g50JZc5iaM+RW83Buj/px37ZwNuA
PwvfK3CXBHA7ucKPqJSVxr4GPYk2gdKc9BQPZYMtXh5u1ViNdwBrt15aLgY6BQs1
RSIIPtDS453FWieQIG43W2LJTNqgXNJ10vyUb7ujxQl9LiTXin4Cm9lhQh3os17f
zHWbVWA/+2zLWgEubVXO/VwQjc8NPD8111DDPNlj/Xd4gI95F2ywIwufz0Ya3fmk
ZAfyNtJwTWxiGvzLQ55ZoXqXtr1j31JPPDgNBF38zZzBKJDbZrh7HVEtO3LoLgsz
XXminmu/bDkJd1j+dCyc0HaoDPgHyEQcpv1DdALe4k4D0KQlG08Mx+xI2swIrb2n
mQAy880rLAYFQWAdlz3W2vervlxD2WNgBGBQRuLAPlsYpBclFulsPsFxRT4Ius1P
lvAe+y5H0NLBQd2R1Yw3pnOdw18RXsoqCt1Pq6VtVdRKiQpWLKLUgmYdxHAjdsfD
hdHwiB5pj0loV5EoSfcaP//FQZtjhh5mR7o2HeCOdbY7PZ+0t73ojHnPF4XaiHdI
4c0n5KymOAUtuOgJpoechQ4hdheD10hzn1ZHA19SRMdCVdEYCcBRH135WRADWD05
BP2XgfMKoLCPVprgr4dZ2J2N9okukj3Lx/+KOT+nTAF4EhAojIs8mxt7gmTstkcd
dHhUoSbSDStkDgeuAdBVn3w61wuMWd8D42XYydGtG/nXCAVxKyj8nk7HPpyavDYm
r/BEMfkjGw2IddKRGs7lfxfLjl96z6BOCOrjF1rkVsJsrOFIvZTXY5uE2iqX6l2T
mZjjDyOIB4voPLnirgdCe355gB/GRfRgiamP9aupBsYkvvxFAJX8gYVfvD8WisTv
6nhSjAqH0YGqi9I6Ziiq45ybTi36jlqwTwccsYTEeSGYDwC5KOXg5DEwWe8CHnrn
MaGqtYf7QqUGvPBYE8eoiQbtIGxeDGFKrBj6wg9mYIXfCt5U/U/mSI+ofXq6SAxY
YTDSNfWfsNd0W4cSueMmSqTO+4LVSIv3V4ylkfFIWPBKXJngAuhMtUjb8GzZ7fqY
d2rb/w9zQ7qGXm6H6CEd6w2Ha8oNFWRtSvZd/9EvLuHQjc23LN1OjMAaYcc0pBQ9
xSsQPyanmHrmVjF0g1nw683QgFF0oSdJaytHAxgv1+ZlYDaVHp0gevzUElRBvTXY
cjb8erOcgl0oqElkontruLlNfXZNZ00QhImcG55cWp7fWjU3tuiozVdXI8KJZWrd
mczJTyyIUR+yTCGWK7SaGbi+ccHpTilLLXIhvGZE8ibnmzZV6FfAnRdnSCw1EByY
9Tt5f6I5pdD7Z1Wlh+0hWZsgT/b3jU1VxpBi7nTfS3Wr/r+8Kc0lYo3fBC03L/v3
51wtduyliaoyoyxp9tr+d1dBRIzx11tNJ4TwOzyfPi6IbvzAUXmFUUSaSjtw29ih
gCAHg75GUPA6HFaM329M4e8xq+RH4cdzxhaVu91AnYd6OFTWXM00p6DC81GRY/ZY
fA2/bUNJDruKlbxYHcDxd1LlEs9k668JdVW8pzn+tEe1/PmELlU8cvJU9V2DEJqK
QGDACekHLD6q2VisMj4+v3Qa4ZCBf51wMSyfdBVIBfFswoMshee4tfImHKZSIJn2
PepI/zl/x5KMQpEuBWEXzvkpxGIkl+z7kNNstxp5NjaoNIzCSzHWUXMUVlHmnQFi
FUJ2fRikBJQhUmoKBEHcsWm9cQHw/6ABwSxpRCnc0uQxksRGcZRn/LKyGhzg9t/j
heu7JpPpWQPZ9NGdw4B5vz37stqLTVv8O2n4XZkdqiDuTE3ESy4LegrU9OP1Lcp7
viQ/5Jt3HXTCFHgvARqNbnW5x4+DR2e577rr+K0XmjSHNkN4vYGrvUv+I5MPtvfa
r/zpJvqoLkFSMlSQrn0x4SQcTpv9yF2l6BCuc8ILzXXOMLJ85Wi3htVIOmvOx5PP
7PFX1nwkCjBNHoA0FhSdE9zmQl5a3rJbjfHz1DxBxjr7HQLDYRZyWbwhAHe5Ub+i
hJmSVNxO28OFiV/LYE+Dx+Gr+P9viTG4RUeNXbC7S8V1xregPuOs7fbz53nEPn8P
IBlEsxeapVmU18mRyMHuCTEhOAOWr2tJAOSsEZ4zEFliYdAbimpALmpuMZuoTejM
OHwtg3ChTM5mNlQyd/49UX6+jnZGUTAAEXdAWbWwSpQhBEL+uwalgsr2cLiqrSMY
Zlp7a8JXg8POE6MmCnE0g4FhSaDU57wi2rhZ3ob+69kDSG5/z/bXkt+o5LPC0QdO
9g7m++qFbMrNhdzXf1P/GruJpGqwiPWbb1bsIT71cJZl4715EViur5KR1Wz8ihjM
2SJ1P+hZ6QuF6MxsoQy0hLUi64VTIjjVP2omXz4HsHs5X/cqUM01MhtVLiDVugJg
NfiaF+j7ABeaMCg5RcI0q26VbkWzMdnzo8g0YHkldq9DFduDfO5H76NpWM+pmd9A
/Y+UsOqllH8tKqx3x4PHnW78gAUMJq+uQqHb32aNV+0neJv8P26UfME2lCkIwCfZ
in9RBnTvqFtcHQz1S664CFFa+AgEf+Hd7IMWW/otaa/AwmENRM8WD9b56ZV1ezfO
n1VhSVrFOMMQdDaa/JE2AsAFU1O8kPupwA1Yzz4uKlzQJNqqcabiYEx/wPa7rxZy
bg3Fk6qi7aGfJeIc9LO6NNdFH09Cr0DLaavKhy9gY/kI5QAt++m1InHKEaN0Svzg
wYeHRuT2CubaggdYuKKSjzVD2HR9wiLURaog+nEpFITK63avOuoStiu2agNR2SNu
8QixgRCC8WNY5ysq/mNMXZxUC4J3GXxgAMzr3YfDTL0ystK7jDH/ul5XXqnFHMaX
8QmsRA+B33ArgIvQQpwjJelt1afepJRpNADOWh1+m6laGUD5h+Cqef6fXrlX65vS
HOCjB8jhHJt2JkUpC9PXO/DU+ikc7Jy8X6TgFHtGkEKga711ZFI2OhFmtCRxHwNE
xolZdJXL1GvjjGJWdVmflPvLQZwtvwU6QTYV8gXdeNNWXo+cfNDuxJEokr92rWCr
KB30KVKJsL9X+jzn9GrdhZsZEpPXqgdPYGcxR+3+Aqe1NoJa++NlnbYFCLHB6g2m
zNqHoz4cUD+BWIzelvrLFVF6W9Ru1od7UQJ4PT9tZb3itu7dx1zLyA0VW5FlCm8g
YAoDmuUz/HVliJuUVbJ+tiXCvJ73zwbQcwC1eGtJrSkErA2gIkhdyuvgdzviQYzo
TI8SIwt28Afp5wj36H0hv1Dj3GO81dzuuNI29InmkwDnPyrgk8b6nPVVtJsErfqy
mBNrlAdFQVnuLOreGmr3i4gvyDz5xooh7GFD31ObsrO8LzU8bF+7p2THidkxJ8YC
2si+O9sRG61Qk8oamCFyHnTnzXuHC6NWixYE9DB4dlDCcV22hs5lGutj0fq3Rg+9
3bdPqQxX5MWJiHEccxHlvmOgaC24zO+HirzlaIJOZ0QJfcqQlkuvrjv5CudrQxgR
XWwFEcEFCaZQozYWiaxYl2hXpYODze6WKfIAgR30gI4CfyGCSKg6sedykMbpELeT
U30PfMk4WKgY2qYV+4zpkqi8WXxu4Dwvel0nstkI7Bed1MB9tpWcGpOohKbPqkxF
sOJaoR8DlnafN62qbu13lnDF5ptk1MFt5UGHaF9jlL3BtAUKhpk59YshR70oAcH+
TcjtYniFi3Ss/HVR3mczYIT3aZK4mrmbY+KL1J35834QrjLo7beGEArGnGA+IiVZ
rP3IsJ/ID8kC0IzAqn0suRF/pfOmvAZysG655G10LmjLkT7Wy57TjqNlKM8ZzaEg
1KKakPYLbvxr+JfVSptpWnspIovqaqPxr4Lk0ctmz1Ph6gVpS2jwllV7VMJaRK0y
O78V37qjmfkCU7nNXazK980QO/PnhF2NZU6pflOarolKNyh0Ky4O84YilBam1Xi5
IrM1gVuixyfbseIlxpRD1j2WkRxokcA0JAvs12frBNPzHZW2kqcfUG6C2T6adYIi
aAziHLM6RqXdv4q98UCdgRLH+VZOIGD78gZ5MQAvK8Aw7nW+NxXs8tRH5P2bD3ST
VYseq6oDp6w+oyjfs6DdYkV4IZdZ+pGa7cRLW+uK/IT/9aCs72/73x9mQKLTBsTt
nTN/m068J2ZVZ4mng+UuW3q/3CShem7BpsdLiMAMpXMo49fCHkOqNjEzcM60YuBU
GJtHv0yBoHKZCC6T1Yph6lwV3bK9Aus9V2rImcbZXAULh7I/ohnnDrWTAmq7Qpou
e0kTlHiI9z6mwsBC4/Eeu0OMnjQ3Q4WFDNytktnWR3Qjff4kjFAu+nmcUXjWmg0o
MOOaE+lt1QrfOzyo6ZxvP8Jd2Vh8hAlZsgEmc4ztFE66qCw0TBbbhcqOjl4i9y2i
3FdS+kZxu/t8R20AjXewxxUvg6sj3DzJf+SG4vwjFLS8RpJsJrpqdPEUKcLFwEPg
QNSzCAc+wuqWwwO0TVevp4lbAqz/61gJeoQOuLnMbRR/dx4fLHzA2KC8xHOnsDab
ku6FwJsdNHM0/jEVMGq/dI9R42d+/fPg3spH8mGgpNxq8DIc+N930JQisfhsr2vS
QTsK8wzSSOsErwpJsMFQMPAu5oHebeToJgqOjV39OKZ5qPJLW05hLzIMPEVaq58X
CtJxDwPhYZXfvoOXbA5VnbO2M2Z/fbD+3LNJXELUmWhnATNGssJ3+jZEcFzvkzSy
Y/Kj2c5k5JwX2lwQDvyZ1rD1w3uJ2eTQZZgl0BH5NrqYfkSRRgrlpL8CdJVN4MFd
Qr4Tgjp697CP3E65nahtFEd497tHdtY3Kr+nAs8WIZqrVGwdcH3qY9mj4nwNSVC9
UpGxO7NX39rcnZx2r/VtMpD70ei62ZY9dfQRs6vNOZqUt0P9RfAFvE0Hpp2yCyxF
Rnp5ogDHhvPHohdoMuKbb1JxxfWU/G64IJF4G0Sqel6EcpUGl+8vn0CcNfFqclU9
rwn+g6h0xQlsOOrhyXHB2h8Xn/CfxqsquYFcQLARWdWo+KhWTpNmpOxsAYtp6WS4
0z4D1j0bUfr6IABGCq+cKf0SHmXhVqdV7iuqLLYtbV25D5IOJoQI6c1t8Cy7ND/8
OXrhx1QMEuPN8nv8mLZf7qa1GnCAaC3loti2UXIR49XHpDXlQim12c4SalmVxz2n
eio5zoq6Py/uhUu4UI6jcmNSShKuhaiObeUXdz0HOXwPyKPu7bhYugw7p4y2KisK
ddUdHdYxTGsLRgmK2YNNQ5bQKH3yYmbREfYGb7rARAy8IhY/fROnPaMIArZteY+4
NO/Litkmh6P5YlDKJE/cCeVPaMnjEiKNr3hgLbUPj3GJMk0I9P+Pou9ctJg9+cg3
xEO3nj5bcrz0bSSVuj+xLqqGfygkgDb2KCXs5cLPQV+AMBSAQDN+s5/CHwY8Yzcy
ZQdrr/I3nSZ7mktwLw2L/opLn4E2+64Pv+noKCQYhQ/dPFR8YnlxQKAbxf0xGvEV
14aZjGpl4S8SLZ3BsOS61ZN67TNii4h3SlHCTQRBx1mDmlwQ8JO7m7xoC04YgwtQ
tYCJFb3htJY42dY/1ESUHdQXM/CV0g7l6a/JP7b+6CTbTlsD/Ix7MdYDZ0hpNYFe
XUBzhRvt9XIn5HtfTR7aUZy2XKCib01yRbphQadwUY4wvF8hSIarmr9R4PI72ns+
adMLfNZk+PlF22nQ4mw4+BKyTP+LVBaCthYAq0i4kYiqiVozq8VuzpEzXU4WITlc
PSeAUGaaAMz2dMTB3YFjVUBkZijfhxvKEWGSyii/35APXFN/01ZQ0S+kJ1mgd70m
a0PLKZLpYgqjWkANegE6ZigYOqKunnRDSy0l3grVp718YPjY44iXln9MwH2J3iVK
xT5c9FymNlNNU92f9AB3N3cpT+0KBGisPatUWTReop2xB+tpXFFY2mw2fsm/Hsfq
Px1j9heTmv9dUL98QIynDBZc+SuXuufUoyVqh4FJfmqTx/LC+IMxyWi8fW0M7nUO
Vt16CV9dv5+IwgfM7t9oV/R6NYsJsX+56uN8+2rT+HQKesiy2g+R//uheOygfWuf
LwYd3N8XT4fb+rrPgSCOHsW1Slg/jUPBShyL+haeIuDytfnG1TA6ZtR+HPCWSnGf
CqfiEDK1ESZ77N8nwdHKiSjIIzjPa52uO8K/sFVhCFcwdfSxoEZdalZYvT0+G5dv
UfFou3P2Ccp3UORqpzpAQtiPDx1DdcnvU/o0XJIyy2kG82KvpVFXOhCJIr6MpGEn
6Bhruig+xlgC7QyMqEPdgI+At71gRexV7yT3iukK/Fr6xmCtzafjgUkl5Faf8nDP
Kmj9WS6k96n7zdbQGIHtu/sU6vQCCWY2W5EDQWlaf60WVLl24i+Gmo5FLJpGZW0l
1KwBek8agk+u32N/dJjKB/08vMqCgTm2SrSRvdlHsBTg0hHDPRpNozAxedpjaKQM
KUKoubtdDuKTHDmYvRYuhpsfo9uI2XMqidbHIWDIb8KB2VA1NTztB+JP+OwByWLN
cl2xnNeTk/AxdacGJ7InxdDuaOGpWk4xigHfCa1xRxVYNx7R1N30LBxJczcuYhxp
4PjnlmbQpy4Czo3qY/SvcvwePlK33ksyuVfqxSPg51DrT4iaZTO6ddhi6i9OPIrh
z3rpJnyBMDlEpAfUgfdXH4UP+yMhe/t2ck2qXIdQcES2eb3pLimRVpd6uSZgt0YR
SlqdNa+mad9EDzZWQCkq1IliypemlRe07F9bhoVo83q+h9Z9TPuOAjTmlmJWBdcC
Z2aULy+4AqgzUSxHjTeP0ypH9dTJzfViNrFvdyOypNYFRDe0fucB/36aS+iIdUBx
HYOszNgnvhJ+JYYqy/tiyMkr5/a4uhfj251tnWjPv1jw9Z9dDbr9KY9qD1jcfj2f
Nxnp30RW4xbie5ZDPI+Ld0QKuQcHjz7iUMi4BgDlvYolgtnrxxAovN4cJhW5mUee
DkLWLzZRXGyFUyTNYch88O5bfQOG6rab+ixbb3BhilR0d5bAvAAxUI0evNR2WUmC
fDLktwUpFo1IcshdNFLVOHa1Uuf7lzVhOoE/JbzHxxpy4S0YGTRJt7PAIJf0IzGy
LVg9eQHrW3HQtEhJn6FX1GjMNW9JFtECHiVUmBvamy+2nl/eaztXhvHYJ6u6pRXr
2FjSk/mWCgro4JJH1jQQ8tPTUFwhbvxeKz2ffqhVlIHD4GiDB3naLhBDWBFkzeAh
89buRSlZZt+z5XbVu4g5a+IyOWcv7+VwYPQyXKG3ZAPX39b1CtE95Qj4fjoapOhL
eJIx60qUVOgG2TVwglaXnUPNKrlhA+oWWiUiRuWEazzLPxzJc6JPD1M6szC11T0A
7DOn5gw8EIMHk89yrQss+YyH2Qft4Td7iDOAHZZ/E+YDPKp7DudKZJn1o1nOTkDp
RnIG0C16+4nVcHYlq4yXF0nVdKNNGXYMCnyShXR4TRNW2ZcejTYOAGFqpw9a/JOL
uRt58Q6nYqX7O7R/1e5Qy9R8a4G6sj+FpUTl3+NzskAFwdeJ2Q+QrYT4bE0hxt0W
CXEvqlEaasJH1cLQ+nGDLSq18DKdoyPE7xlOg2h+FKmOxDl+cLt2dMozyO5Ugdgn
RfNlHJXVcG91xnoAuJ6KsJN59SPrMgir5TUJCK1VG091WJjDBUnRJBwe9t2pswC2
MWxGGHkj7jrYTyNxqnK5sTVBWyvM/3EveRhwpONfZPS3wR6rC19iPrsrOaIG/QYY
s/uW/jgOKrCFervwCTnaYbFu4GkO+XZMQws5RKEHF2z9V21zOPGIS0Wl49nIUFvJ
B2xRnU5l2/VUyJGV/XxqMwQc/NICW+HBIJH8PYlAPx90zB94BCIVMD9elGmjjVdF
p++ARCvuBXA5NiLzu8Smn5HEboP95eyb+i48k3vb+jQ7jnHD+ZW1dbndvkszO2n5
QybKdTALqZRb1tYSpiEijcXa/n1u9pzlM4QWa9PhOuWdOq2KOtvWAUl8iVy2oIJk
K00IkxmTWEio+7yKt+SRjz65ge+cq54V74GUaG0VhCXEiMFb9iZDlG4vrzcnPMua
kaOk8BUu7I6aZKUW+6+YSx+32ZCBlcgwq3fH2iQ1ZJddPqH0KAdXzyHvgR/3so++
5nzqLo0TLRjWj+a9/KmHz3vjG9NEpLOp4u8CZOEizp1p2hd2dxYvFqPk68Bq7AML
pN9xYFcHljsWaO1ibo1nOyPAKLeairmVzMfSBdLl0rNEe9p1+tczroJUmHYeybHJ
bACBtVEj7XtiExBhB4jFdPEVgbCQ2XLNhfhC53nI9CBDGneZaxLY6JrtUTYwjKKY
sClnw/Y6sndksRylZD5M2hNkEPbfyBKxpgwp+mxHFlAgG6Fm7YzxLmW3RrhlolET
Hy1DVP8iSenP8mBEvFjmGNVSNVk0H/nNXBe0sQSxb+nPJbERDU/ZfQuB53ajh0fg
YnRLSCi/V4zJFINstfA8S7FXC0SsGXFhzGiSvryE0f3u5c1f2TuZY8ryEgJ3GS4P
pRbSDi5WhQy5eWG4W13lMlwo2i6D9ngGNwEw7t24TdBbN+jZcW2s1d+kHy+UnmP1
Q6mWVqjGduvZ34xnH1pHkHMs4dkhvU3deGvXAyOb3CtxKIuBN6Eg7oARWOT61Ehw
t6+slNi4U4QMbzAjusHC9juuznrZBIT1uVQ6pMclCXdVGVnvfrlpUrnY0NUzcMTv
Pjo1cos7rw7kW3svn6xw4CH/mThQJvQiZaoXFstgcrg5YONsWgB7IuAF3DRmkK8e
+tm4nhe6pqzfPIbJZFOjxVOAv7y34wLXr9sI7rYEfJYCts1EHxqCSPNzfNsQx9x8
LZYGTXkwSe1gEluZH+lCOt+ox2SluNscMOdj9LyKEhZ/ZM4Aq4gVY0SIYfJ94Jov
vmLjKuH/Kd3tsv3d+4xIpJSVnhn1T49yHDwyI5totgZfXPdYwNTJnJgKAa9WrcT5
clz6I2NxRHXqpD9PJnROoiilDAV1Hy2oXYMQBY5NyTnqk+m+zn3d7JQ/ZqAfMty6
zsdevH9V6P9XLw3XCusImEZ73yfTdDQueAriy9d4weNXtUJdJWyoc1sYECkNc7Gv
oHxNbBRktwFuASgMl/9zoudfSTA4+bDuBWaWZjsdv4Qrc+vtqn0t6M7+2Nf/s76R
g7slM8Zipk5Nyih6Ihp+Li0TZlH+D71qM+MAGUZmb7VPtJx6umQw3TMbxzlfigaK
jiuoeEV9RjiDBBr4o/8j2e6FMi46UsI8ICS/IUl2iYcAuMs59ApR+mT2lEoZGajr
8kEXLOfn0hNOAmB5E+KJulaXa+VnAkrQtMSpaF/huECg3XzJjpjzsA/lb3P0hpwT
WQmbv0k44KiCy+GECzofAEZ0ec/8M3L2jcbWvx70b7zD6rs59jG/Ez22pbzDSWPN
J5mFIkkopX1Kz2ISM/l9Tym9K4eXcg1hiG+dB2iaVI8ImyvnhbIGsbzI7RdApNIX
N3xy2A11NYbTmng2fDZllLlLUma8f3VPUow2yOKvXpwCZov8Q4aiG/Q8MhzMpE2J
FBWMmgRB9k+P91YZqiEDXw3luvlDYIHRGr1b3Li9S9OjGnFCmGdoEadxwmBPZ+Jd
QlzAIA1QhKAGfiz/x25sb8u35yP++VGlc5nTrUPGfUs3oDRkGeg9ABL+JVBqSlYb
OVMkWKynuK3OU344l7c/Q3uoFPruOP+Sn/+qBNdrf6zLPxdpQ+uN/AwZKnsdcK2t
q9L8ouEwWbw2kF329FWpwgxTn1BixgnRyjCVcAXywdwVzTNJ3APSq2Nf3T1Rd3Dv
+0RH1tN5f6pPSu89MoXfMbDI3IEtKI1E4m7OepjmUfpuYCa19iyFBWqo8ZF/CHxu
5zx/e7FlHzE83EPeVGHq240TQjEb35Op+dHUNwGEGoR8WdSDi4ZD/sv0RDlqARYA
GwgKF2n08WTDxreTmfWqTuT4tvQ4uePhLf7of0zS1DkBZ3VahM6072/Tk3At/V9y
NATBbYXo3kwCNfI8HofLaqXK1j/XC4fokDDDQhDDDqZRxMHTb/LnGfEQq3nt7y8A
IRWHF5KIg+kwxEQkqwWCr4WKNzq6si+48Rt2jRAHGWKj3d92Xu2Tarzpxfoq2Q5e
0YiVHvX+oZudgyMBq9kA9XH3SnobZX255lUTXRKtKDqUHF56y5MuVE8gK/1a21CJ
ko6UYeSYWeZX+5NG/U8Ldi1odxigYHtEJzxGi0PYNBYGB/fbO4bXJ6c2YQh9uulY
dj9Yk1BlM79ISH4DkPpkiJweFMYPwYCaGJQMwIF/4BqH5dvHdWJn2EkkXw0SPUf8
w20wN5ub8jRm61J1JRR6hM8IWMFh0M/XacQFs6hxPcqM4iMg2EiUyEUvi7iLMZSo
6TaKf4GW7TJiJaoVK+RZddXNizH7HHWGXE4uuSmRYftX+goZpNbx0adT5Z/Jhl01
N9sCfzQXz/XW+fXSZTKMpMUz3Iw8Q3UkseTSkeVi7sNinMg+BOL2ly2Mah//d/AY
86jGPDo8GwEY31j1XOZozNMxo0FrJeqpKYamyLoPwo23QwUBc/zMEUn3oANlIHld
InmE1jRGlEBHVBBI5LWA3bjxYqBgBvpiq7LfDENHD2gl7iF6TJIXPDTmW7bvVxYX
XvUSmWZFnKgIwPe8juhNs+N6ugIJDGhiPf31vh35/6NYpGOcB19rvZq5zH65W111
3iBMdCBtr/IC+0u0MVgTDICMuxoRhGR7k3EeZwXwaXiEaFPrA3HJITnasda/A8Ra
VE6XmeAD//u6DlQgpneyNRAUIHngVXBKGMmUZUDdmL7a9AZ1m54jSE2bpjMMRgcz
qQysaIwz0DcO7+dnOSHpqnlIl84gSvsD1R14VOY+naONByrrEIF3QNdyABLgz0Hr
rj5B9if/XyvgbfzGl6a9td8fJ8ivnlr6G3RLXBzjMpAN3Xo2szXHSreVKm7GlnR/
vj+HaBNDEXDvk/7ZdX/UB3NbT9wafPnMo2mULjA11YwdOUs1ZfEvPujNiN2va4Dz
R6Y5hYwrLGzYNU8PAV+x4kPAajS3eCg5/qa2I/Url5mp9RgYNvIdmRU0HbnpI8nw
aEHYX4hUs2/IEqgpr4fU+dvOc2qdyOCgpp/9MWwo35tHvnwBhP1Uk9NZ5I+Q6aZp
P4AgIlh9ZDUmz9ZW7Qx89a8TWxLHMygX/yIHrenxYE8UZNG9BeliNWuFtFAzF+yk
uMAN0oViEPXcugMLPP8EPMKvtB1ViNVlXAYdyeJ9MBHWwNEYqs1PDbXCU//9lteX
+eYopaPQvLIXWH5jHzWpAMjmcskjf31eFQVeYh2USk6r6UHTibYPOzYvLZ34yvTL
wNkaszJOTwWJeR7f0CRvuyDpn5R/bIl8mtY4ms4yGeAdgQwmPAhPTsE3/odH/s8m
tyGLw66ApMSksaNASDVnbrj/An/HLGoCqc3zwEw6A19uATm8rWj2CyppvS/Gbfmc
HSNVO0Nm5UE8SeWZQ+scuVwagcotaRZpi+Jxfo7zMUtdlZ3H0rzDB6pZpiJHjnIJ
CAvWwhBws9VUyqCMqKjKKNCC4Bc/5UJrqIoTbW6fTEUbSj0Epviq58ZozRYvXOt3
qA9HrhzLdxfB41QDqOsLQQ2fNdwPLTNWg0wsSP2qNLfFEUoixeHdQ7jCN2beDDNz
mHdOjyxjmkSWpdOuuYIPayJQExVCRvEGnGUZP1B55aNCm90g1He7UfUWZFY01PP6
c1VvbbtVns5iYJyPoYSELqKjyy5KcClCKTrrWtmcrV3+858pyypa5iyMN1sS7atH
uGvxz8grdpeDNlb8K6jZKPPE//N8xZqvsSa1a7mNwuBgm6eicUYgEU75a/COo2L8
V/yzmvOErrosafhvqAHMheR2oyagYnX6SeDDw4LfMoeO+h78zDtcvnXp6ZYyS7p8
eIRHP7hBbKSkhBxcWJxMZnv+EyaGbYKCQPp/5D9cP/vl1ztSZvDXEP0iGu3u+ZGl
ZlcbXAvqCSXWrmtH/6nybKa1HoBQX5nZohgt2qT7a22qrmPA5ltGUMePgYjiAbFq
ecrE2viVIIV0sYJDixSgykZ3QhOPP+fY7JS0CDG3aIVRHjBzbDGog7So08L+kfmj
voFrJbdwRHa1b0naaE7MKMGxLrBydVj3verJFIpXKCRr+dTMsSvZR/50sya2GHp2
xHTc0+dSQ+pY5Xe/XwIrUSmjVsAj2xXiEluqbFKHjzDPfGVwn4UQfkQrvOzG7Zf5
In8d0Mj3MQJv12BqoWvA0h2dDgo6mScqAd45klkfyeDg64vNTSd2T3xTONTZOoA4
R/cKgdxeQKe6T17hS6r8oD9AUIuKzuaMLi6E9gUx4w8pDi4ebZWC9OrSJ4/X2HVF
ZO65mFdF0Koo6xxlxu16JGWfYoU12lSSgX8zFBZohisgR6pkJq1pR83WEUmtwSo0
eVVGb38wI5vUZ0vqRc8iRR+bCAyVtFk+ry6oKI0Cyr4FF75vSNnzrHIXW51hz/8M
G5J8rSZ7AmTnu/6aD3IemtOoALpRmtibj1vLYRfqBB5RgNESS6ZL3f1Tlc+4CtxY
xDs5R2SS3GoYthPA3vw8b7t/RjPt+mtLPrAovga7ZFC02Z/Yso1/XRpSbQMYv743
t2c51tyfLPAi39N2nKnH24uksRx5aNlPBhiokoQonrlFVo4icp6vA2IH48gtnOx9
NfoQMiORRZQ80sd6bT9zT4iLOaPY1x1oraR89DUHeFieK1MlxTdV1TCsDxHem6Y1
XW3fteRSZ3gpwOgOdl5n6KWST9ZnuYt0N7UDQhOpO1j9+MU0h0xslDxyehm8hJ91
NhbRbBymFT/dpdmjk1AEc0xYa4kZ7k7vyLmaRgy+dazRFhWJiNVd9LcyoJ08Ainf
nzzdd/z2jt2VS8ky14S2LVQdpEO75iZpn+NDcn9UgPy2YrwrV98w+odWvQNqI33x
SbOxLynIuBDebSF3Xt+/uj8NWdqjnJkgEtrTUfKxG70ICN2KJk9L+KIMVBcBREFr
QbwTVsKMsfHl/4REq8WzDmc9WWn4IS6GxCaWDBRcJxrF5OxAG+RqwBSmSChS2FGZ
hazE3JCNHkc3JBGTD6e/GXgLWbefz27rhKGuBlSZ4jIlms3N23/KRduil7V6qGUn
qzXMflcXZ4brO2+ydVOPAr2YUF97w2QHoU5VsOsm4fODzQwMMjZVvPWIIGXOP0H8
2JlBQbPqZ0LfgUkg5tmVtwPG9Sy48IyovgsIvWc5Pu/Itr+fld6IxcgsFLTDbpP6
HuFfr0QUDX9xQ3iQQgIllqIahaYCi/HdiiQGD+KRaMcdG/Q8yI2y9xaQBBT+vjID
cLKcnKx0BDbBVpVMxFANNAfQhLVDPZmFQsOjbhdRjuUjz5La97RS4vkY8MLrkL/B
JGy3ZSbRGKa08m3pscKvaYEhvIYR51d/xL5eknX2NDf0RrLoeUcricYk2zWxmU29
FN6Yh9R26QSCYnAdoBhLbNjkpLtAbjuYs2/Cj7Fv9Ub/cQzlUjiwqmor+YBSYIud
u6gTU1OHfohDc2h0/2uWWDy+wSSgfnKNO83uPrc5za+BuygSyjCeOEta+r4+t/Oo
eTdqxpwSkuU70JYITZZrUXAjJOrKQsxdoNnklxd6voCUR9X5GCQVC8Tytf6zYfTM
OyUwJproH1jb4IOYRl1a110du0KPzLp5kCiGXBUPBytzNssrworPprN3qHxn6rU8
tqzIHclF5YMJ+x1hQPWacAw7B2B5AEblBBkYQg0O4LAOian+0wDmuIipohc6d23D
5/sXYXlyyVZbjWjWc68xLFK9n2tqUasWl+Rs9Cfeuwbm0i7FiQIgdO0skk8kRZvL
r9klWFWcXc63m7/un6r1cL7CYWoX1LxkaUnAu4ms3478NJpQJeCpctSHDHbdDpmS
iaXpOS4Q7yjLMwgLAX84JiJoG+4QHne5yaCucn9RmrS0D9lUXGwRrBb51xffvC7D
BHlSjNVllm/RmwTfSmmWsobH5kG76CS+APbAyjRuKYZWfyrA9HEJN6DoIcHZy23l
ONWXZSYvQdU58KAgT0hJrHrAaLSKeeliVbkGrgAR/5960Ax/hKMQhqmMg+xkOBdi
RTnHq8djY2y7lxlolzIDjEreZqZGGZWoqdZfdZgjfFiqdYhdV+9AtG6XH3BKd3ar
DZolsmv2KQk4AM8F7PrYXGJAnfzOmW2MQ0iNbbFumqq+eup3ngEEVqIBVd+/qQq0
h3LxZTBkwuaeNdN7R4msxDdViZnmBiliKaHFEqeKWw8b8RHa1JJl8chTpr2Ob6Fz
0To63or4zOeXtaCmB33TzH22TRROEYjzBhEKcw+ghJiJgg/6P47TlA8BdatWynyC
95+lfUNEcWzjAGWyXsdNvGmuqU4XT7DunPT9AqGosgc1Py4V6tlkMksvF780jpv4
NjtQdEZJbTAr6J0HEZFIKc5CT4R9i+GOEYgXA8GlqGS7nOMXbOw8xHmyqk0uf5sd
ul3O8tJ3J9o1r4IYAhyqK9+Fry2vsHzCnbXmVi2EXQHH6ogZlRRtPv995rs639E+
Xq+p7/JfF8daiyD2NH4GjOyO4rAxy/JDWxbqB6A7Xmi4nTk6LJaOoXJUjT1EgPp3
SSgAQG1YhKCxGlNbP3FJTH/Pbs7vaQy32Rw2RFK6BG6PsSVQx6KvkazH0UGcRIKR
z4QTkzToMCAEIVMtj4vAPjOEL+stmWscJ58u3CBjv1o62f8esASBKwPOk8HS52yo
X9UGhGoZLw/Y/FVyuFH7zIH8EqFEXUN65IUE1oFuP74cRw/wOToxjM+v0421/TO6
JfuSIIlXALA5ezfGaucx0uonClu1wQpNhWUblSple2xeEcUATS+LlpWApPBE4Ar3
NlcSgCB3xjYWAeWyi6q/LIcNDDLCavdwjVJGcMBtLyHd53q8ejJNsYNow4Ot/KZV
emo+VUkq4CLdvcMgFJ7R27uZCX0wnStDuNaXBy3sl5usOTnxeGwf57zn/NjYACUN
BxqrUMsbCtHUvzmkNcICcKFAgZb3TqTF8x54J9nQWsXw0I96O3IMSo4IL8pjdjCN
j134tQZX4nmjh/CzBRi6pi7rbRhJOJgVchQxnK5b7s2AF8vuUWYqfNeFFXa+4AyQ
9AYtgWLsIR5mMxtG3+hQ3b0By2SnlBGT6gRz544rAIebqJFCDFYowijK2ndM68tG
lekpnijqKNfJ7G8sylgONI/81pugmPLR2s1mvAybQCjeP5BuaDvArmRqsGWjqspx
4ItAdzGeVfh8y2xHxD7Wkzb4xfgXMHkXPFVRKV8OHIfyq6dPR4zNO2ns7db6q8Fo
SEmnsu1oCu1ITjfzpCskkGDYXX5YxOwz/ohAXjBmzU0u8Ra+u7CoOpGg2aDTa6UK
OcO3I8WnzcUxGpoUivSV5QHRnMAzCSMIwtDn2fCYq6m1x5JzyBaiZ1AgRCZkEvsL
pQBx3DHuaVuyWE52nt2QuIzVR1JTV6fUnuU8Ol9LugIAUmvALKN/bFmE+tU88tpd
rDtUFwcDFvYCT6PnmTeGpqQhZYE947Q2RmtkK4Ir1sMRwXoRr8qchBCxFOrHKwnh
usPBiqm7dOsAIR+TnKhisFmzROHrPjQUs/vlwumIy1WgIQaf82sgPqKb9qYc6vM4
Cwdo+cSmRonYOipnf6iogwhdCM3nFKeVF8GqFBPyCZiHrDv7IAoh5MG0vbbHzEop
Xc5svWBi9SYBdkWCUkxeETFk8Gyy5afE/FvNbDCYsBI5aMDQ+HA5bNaxPbo7lPSs
rBTEC1tvrpH/jXxe42cCisJgoZa2PP5z2k8MLUZz6kdvDSttC40btyE5eLqr2BK+
s5M25k5AyGf2CMc1h8xvAtP6/+s96tfN/5LuQeoPwuaZVbGy6rGUaK7u5p8xET3T
ArQ1Fnt89awuqOfuaiR/A8sb0zE3bLomnF2NLIH8DSdswjdv1VHL1yUo92w++512
wDBumYhpaZV8oEd1JkIICdd1Xb+ez+cYXHTzIMXdsKQYk+4bqO6CIqv7EfiusT3I
o5yRy/K/Pc9pC91QR3Ej9yOUm9edFokbw7vzSAmiS/t22sRNkNUq7Y/pRKCzzf/G
yLTn/mQvYMCimv+vaOQwbCegYVEfLjo5gEf2TPfkZODwldYwvogkib/j/2o2qWMF
IwMn3L00VOEBIBejPk+BeEGB9/vpHuV1X/DFiuOrLPm8Sm6uu/rrypt8HhU0HOLY
PRpPeqoolfmApAuAjnmB83CZzp8dUMACyeoe41yfa8eyUcW1+uYx1j1KXieDEeFw
hcl3um7kyS+gZpemqOfUMdZ+PhiHd0pQT/+kpoThAiWumHanYQWu7ePHf6f5u9Hi
iLX+tEPC4Bxd3biIrNcXRRWtxKyJhLr2Mlk5EENzS8MA+uf7RDzDQgvS3F9uaaOe
AqdsXuWusMX7fb1oaHsPLQ15wgDFnC1Liupr1/T7zXOLhB50ha2W7p+nB2StoSDr
pAnziVugu1aPr8d75+xC0q81dN/NWj0va+iYVvfLgzV6WBr3NHQp4iCojvJyj/v5
9l9yD7iYjUifV8bkKGzChgCUwACcLD4y2f/Fqh7dvjlixDdjQQdB5Bz4MvgHlCiH
3MQJwoOslTywrkufDEaBBtetEE2tCFWAExupwRzHv7jbkzjoQBl3B9V++5qhdksF
HFIzyu++/CTx60CeU8CFC+uqJ8U1TjKnSry1S34srZVo2WxTxcTAI1uprFiL2ija
GTu9L939N4BER3D0qxWOph4BTwbnBwr9RWh7W1Dz94S4wdvfMffdJH5eyC9wX9GB
jmGLflhQlkYSN96TKwmVvRfvG9Frc2r0+hqXKbFmJmKB83CmfO9lV2fvZ2hVemHM
2crKnF9+eZ9pxpQIKo+NRtEhk3PLVQx9nkVe3COPw1mJqtfu7uQQxc5pEm1Dayji
d3iah2AzWiKAT3k5HbpTUjMJl1+8ggMyiPfnFu7+o1xPm8RO9fJGXnDhfB9wuQvb
CIxCDHGzqDimUiwYg1LoT1tk/nNnsQ5Pin+6XVuN0I6/9UNLs95fvsjQBTqGPE5t
GD1L9pFvhV2JoxXaGiEVvm689kpqs1CAyZpLnThDKHtRUNJ1SuuscdvUF+xwaOAH
zfEMUjdqT1jlP2Ms7HsdTC6RL80dGlanEOnzm2KlnSPgGu7l43+aq1RGvq2ncWzy
tTADMb0fcIQWT1zqlnkPCpar1uq2OibQ3kNdfGJoHdE27NsjM22vKr6j578pJgMe
658qDQY+TNNlH8huFs7KLPnjfZYLv7gpOljsNWYchpXdUObi7Fj/3o54tXb/kh25
xJ40UM19+6sZEw+IZTcF1DM5qXDLE2S4R0ysHxICIvdZy003f0LyRxpCtcP78wMa
15AQ+MsezAw47NBUdbF9exbcPrRNgijmUgAIZDWURC73WgDcBmRuNxt1mnCVDYcI
nEqiR1CKxvYlUWOrloO1cZTOir3OXgbYU2Pw9tFVOzvl4V2xZH7NupHUkad4efsc
rnxO5heY/irRlCaf/dehgcnjyUDl+dP+3oslQN4TZzJVk2ZSfXlZrsCY8/KiW6V6
a5Juaxr58ZAQwmfWgiNs0d7rFh7mqhGRPr2zbS9gYQdlmL7TXoz05jDThyszz5TN
afA2I0GXAC0z12hz07wSNS4Kd8x8tNHs+2jG9fAUX/QGNelufiI3IpjdnwWSUzil
S/KJj6xEprQlqZ6hPE566ZyoF0WGd/I/7aDk9+WE+cZ+rFxr46Y5BeUPnBOk3gH5
iOGCJF+Y1+6kcxBBIYdJ7JDFn97Qr6mVvLBXrZrbaMsiQ+V6CLNPg2YxE4kDP3hx
mszfTMvaPkbQ89T2kJbList5DwZqxcr1m3Hmb5TI0Q8jtHt5aWR0Pxv+Jvfrcw3o
vDwgqDj3CB2UFKUax7EA16oFH+Tb3SI0AsKyvdqBTnxuB+Gc4NZ46epfIzj4nrMh
Y//HKsCcs52sdtVk66zjmjs9H3UuPGVrvmsHUItEvCGe+4kIwRV7H+AqYlrV5+sm
QmcISQBc/4MnHdi0ubn78GDSfr1DPxpAf6nTIRe4Vw1M0GPNgTpZdOxzYviCeMBk
6veWAaIBd2QFyoqx0sO5jZkHGdJPzbEW/RipCEh3O/IVwB0z7PJ42+wFigRupKli
CZmQCVbw5VzIsNdMvxWKhtFffe5JjE1bbKciURs8qYvSdk+1PCbxteH/zq/q+MaB
zJofBlobnqVZY07Ls7VwF0SmVr1Pp/m5TvRik9UJIylmTzxYryA7vZpb0FnFhJaw
eZ5W6I4ieXwxLTD+RDujwnvasCPTikpySko07GfPgBdM3h4c1hgz/baiHGYHOei3
ftxUXkG/MZkYjZIesAHFLqnrZgvDiyC0zbsr9JDWObG9fvRwYKc5SvNr8T1V07rh
wABjI9Q4YMXKLHVkkYgJxjfoy3Tfz3HoZ+Y3piq66F54W9sUUk+8GIPjeLDjBoJj
KkAGuakfxiM9C/Dp3CB7oJSCwT3GtctNRE9Nr2hWy6xfWkvwiHHv/Sl/XGIwxM73
USrM0zl/pATwdElBLEoUwqVhhqJlUUFNS2eQxqHfAMsSYxw+DscJq6kdW/J6mLBD
ofdbBBWCQMBvb24q3H7A8M6nKR5INiH8jgZCYqzyzhEQ0LqAOmnvjnfy6lisfguL
+PtbsEGLjcSlAKCV+ISkuE39CNWsar2+F/CHghTiyQAaiZSJIVCW5L6E0Nsvz6v9
Ax1l1A5o8qNB1Hq1ggD0Ck7zS9TCCrWKuIYFWOzqDqYp5aV7w9SlV66MhCp6jwXS
NmMf8kF5QMQ7RX/evYE9FMXA+ZuYhPK4xJQ3oFSyjhKjWY1Ot3RQxVtJenWLNc5j
GdrmEEAX7s43ST/YEr3emCAq/cfAAl5MFJWXg4DhC9cYhFBH1B559uYghl6SRrVS
+FXyadG1QvyIn5TIpqkEAJCAyI+R9LrE4U9uatSXT0vlbd+6YFak7R9hIG+estOb
xWxbZGsDSSs9pmbFn78cxNmyniORek77x6gsIBMpuiO67byDJAJjsNcmcfLAiDys
wapWaTDH6bzADSRVgMGycpMG/iQ9mOrnrGlc6O5jM4XeRQERNuwxs9FyD+PTn+pq
qf9qn0ZHQsV6XVYrRuY0k7KXl9dUm+g7GGkHvQ6ZP4QCO42mpM4e/MKHhs8cIynV
YDCLEwHBX5PDkAORO7k1qfmWlN3CBA4aUTZnKGqM8O2qfCSyK9mfnJnnK0QRmxvL
eZc7wBQ5Z9Ac67ejKArG0jOe8ouaI5J7HfR8K9XkMKTO2upb8ILEAd/ANBZt5jGy
ODbgpJ8vJieuR3CDGkq2jpka+AOotemICYpt9578FdaU+s//6ovsJsQd3uElwvJ3
dKyPh/ZA6Oz40ZA99MJSwO5K24ZIRm2gmm+ral9tRiuQuwdWrCOYDDjY3TTVeAo2
QCUcdTv8/yyABYB6N1kjvJv75XJaEo68XioMhrMTzNnpogC0zQQj1S2dBScV09mH
lMIm+M3pBcvtWOWn6XbXRt7CWX6OO6MzKKRad+A3I5MHcxd12K5StZ8bgn7RrCu8
scMyuV9mgddWQVCXu0m/sYLq+Tb3Qk+JRbi88Q7mQPPUwDK5mPQN+tCEjscWAN/J
ewmdSB/380GuzapJsZIX+m+nj9NG0E4nVI0LUEFPJj7jF4FyIRczoJTkoS2uSokx
HqHkg1SHDerfrntuqPCmaz+1rhe6sqXu0WgBv0UO0/zDUmGPnliCrYhC9uEDPR6Y
dATSCnNmCMXwRwOHuUXedXoBVLAtoZbYS0RtLw0e67qFquCcz9+4TDgQpr/qEC75
0QOJ9TAeZZPIJqXjegKfbaODF64UX3QFAiuwe07frvskjAIb9RtkePhfcuFJq5zQ
wFq3P9n3Whq8kYoj+B0Zl3IBa2KLtzJ3v6LZmOj/kuDBk1ftpMxYUP617n19b2er
q0fMAfL/9v3KkX2RE6f27OlDXQZkpMUQ6LaDGyKmtEGk9s4i4KvESFyC3gYPnkNJ
3e/x4WX0c2Qphm4AhgG4REvNnPsiJceKuFuNfI1mSDB65iwZIYfk075Io+KQRDaS
OKJIX7alziN+MpeDI0zmkNiqq+pFibDlvZOMO/ts0+TWZJ18ljtOhKLdDWgWsSF4
dSB3VlorL9PzplIhWwXWM+pbQgK8h/8POFdutRybWGwmH10maQc2aL7HxD/Cn7l7
Xbyta7nLDN7f+sZQr27BETu6G8+CrBZYDIhzKB9YyVz59RbfIuw9cnFYBUXHokvP
6XFrIRVkQ6S8Suz+gukV3c5jO9I8ElhHDCvWIXoHo/uNIo/ydDsLmO6toTgxXArb
WL/0IkvAiAODIGhmErOCtHvqi6SwLF+c9/naEj2/ZZF6eqbW6hx5iC444bX9XfJk
dJKh1N1W+33lq1EGA/74GRaYKxzi+CPUD6fcbM2DdA6YuuDHMHAqtwWwVT52zDNl
O7QSt6X7MbEX2tFegKwjj+iZeQW79z5E43xL8b36f2JZYFwPWeMM+oFC2g7Qwd/q
jrFT7rmkpH3XQSKtt9nuVfLeeoO/FNc8qIVd2DLFtE5iju6V+CnFEXccsQgB2zSy
cYACDItPECav0ODSD8CvU5JGNKBprpRiFvZD55OOVcx4IJjPUc1dK8q8m8+OORJd
7KIstf1aN4jQr9fM98IYNlr/MDiVT4/Ci9hs5xOFxv2U3KNihEWdN6XGtlk2I+oN
hDM/09ljQJ495Pn9WMgKLB3s1Ualn+qMowByYsNI6SnJPIxnAopTpqdp5VnM+7rZ
GgHH5HF59tqvQVPcwtPMJYo+DkHhtDvkia4k9yj0kziQubxKWHRTWr8abMTUyM92
nqtVISLyeoG1ovoB17t8I6hqCvWMNBsw0dbjSdLKpp6e/CYvB4EjaibV0LtlwlYt
4YFe0bN6Sw7O7T4JEINtDHqICGID5uMEXwOqoE9LwwOADfgKC3esrvNX/caCucMs
By4tYtIyklmdVQYk3XpqbfpfWPvL5BZ7xp1SF/NbgwxzVe85MjtI6PZRp8PBwJtE
MrNH808mwjJyRQrrd9eJhlVblk9VkN+XrQtJIYv67JeRBt8l+9elimjXGLbX2myh
wLjTsRKFQ8yha75W+R+Df1FVwSwd3q0MdX5IGQR+mA/DaGJdwgKE+tKMHsqr0l0r
xZQcmHZab047pzET5dHlLhOxLwLjHIrK6Pjd85p9WnAP6axtjMTLO4SxKwQLWsG9
+/ydzMZ2TYwuAgW99QaQlWZvsHHYArYLuYm24nN+2MhdN4KHvagHz/2lzRaqo/VK
rKyqD7oopIITm9akg57fa9vjx1siruLE1VEPkjdR0kelK30IFbvkr3NI/gAOsw7G
r90G9fNPGWK8iNcLhs/xIcMheJhoScGD0v4kYp8+C54ST8Ept/DHw0iLtiH2N2fR
kqCj11pp4+zae+dMvMrqbhj6lGfZhyN6BAwn1SWEQ/abjKrBEkBLLrEN16WoTUoq
moI790hNZ8//BaCXrOEgrkwWxV9l18OBST0J4pFbP6qoN25XC3mUyfCMt8715tYy
VRIBfJdIZg5jyKsFDWfMvDJoMcm/rD3SstLwIIdQyKm+lFczLlhVJhYV6WqazNzx
kszKNcH3/RXA6N6ZW8EW12M6sSOpfMfgtStuvsgMbjknhBqMdeqx0cjXEEwxyUgK
CKC8Jp/iEO0H+chFXPALqr8SbO8JVPlyKVj/qoECa51+Z35T8iW1G/jb2c5CBL/5
NAmEcxjrtquVOiQby9ul8jI6fSqnXmWOZjfbHy2ASMgK+hGC79CZROsm9rVg5aw0
5Yfk5hxLRsXj+ZE0hzsme1PmMizQRIu8t1W5K6BWe1FchgMv8MtiTJxcDXHWVs8l
SOlMcBjFjbyBk/hJfbZqsDjLP//IbES6EUyTgJ8UJkxk36NP1tF5pboJwqbSCvQc
iUhPIXJHIepmDOyxP1BMaIlv+PAWjYlrh7PGciH6y+lDN4RHiYmy4iVMM0i5aHQT
cL80xbDPJQKvb66pBH5m+VcjbwBjX+XNjg272ogp2tHUl3xj8p/vH3a3jrf9Ca7a
nPoMQz00nVbDkf4pSl4IA9SdH65EGO6eqfsi5TcC5tYtXX/scYg4TYKs3te6p4ZT
+Bvce30SWvnaOZOo/EvwphZ5Zl9ObgGTig2U0I8aeUzJ0v5Iw9E23T4E48yeC+dh
iyfg709OpGge/MLuHpTUVpDqwbsTQE0AppfHjTw5M7kgvjV1HzbBZZFYgmBN4Ck+
Hu5R83FZ2cZfEujQii5bJgFSx0+nJ34odQ5l2ZfolILCaNsYbFQqXzgMBTAJA3Qb
XmgFbXV2sQKEwWykRcba/MIHmONufXhkcThfkNJ3P6ApmaxnPvdlmrNQdVud90tf
fMdFB3K4An6T3dK8I4Hf0jYL7MgvoiVVzZUkVW97xDYxME6xlBOjJ7bt5MN1oq2v
n6NmIhdwMxaVVwBI5T8AcJlS+3AA6Bio/JcHQzBkSY1xwvv3f8pJN7ttRqz1S/nL
7dzOzjEY6HA+Y9Un4kA6zGgUAORJzWHg997bZLmQb28j4sAOYtFEfFIs79mj7Wnq
TKdo6ourQun7MJeTlbJ5bAu7w9Rz78RJyRcqe1rX+yvHepOEPkn71G+2mpY+H8ty
/Nq9r59bL/t3pY0SNy9OVTPU/pIrXMRBFo7R6lqKoxvq1Aonw90tSMv3+ZmwtaKQ
bQF+Wy7+UX6p7y9gPkjeuNMg8eypsczzW1wv9CgxMcwtZJibM2cJyjWFr9XGT0eW
GtRdNzCJ8wgqE2DQBD0xEX23Xws/Ljx4txTonfL2btd1y+Vl3rjHG/+wJyD+xpf5
2t83F0LSuDi7/2bNlUza1F4XYBpumQ6/ElaH2HrVvkleBrQ5/NR2PO/Ca6nU9JVw
4fN8rtVmzH/vfUzHVoD6GkuaRAlnzjneKANmJy4l+aq7BidEaEg4RPWwALy17RHG
2jHnKisWeIRrZ7unZzfJI+1yHgoNY37Nm72xA1UhL0fswUkA+clg6nkLbdu5lE5B
IxvZgrl/bCtaSZiZyc5fGqK1j2b4KWFQASnBNepWvwgEOP0VqhM6H7uKXA5cn3vq
Ah7BMr4nJ07HvZnUc3SKUPbsL/aahbJLhRclQajvGUvhj+h/0E8HaXez86JVglJ7
2/Hi5/Oq463ZKBNj/gYn82fq1XGWtzbd4keEg8Kqo48HqM5NZTkb9oOyCEonIzFI
UCmnUxoRCkUxPgqVafZb4r0nuJarcjSRDKaJlbZTBFsmz74DeX7sSGgzjcEJPf2I
RHeGGRLuhAnBRfUjI9hNSFZHRk8vIc3rGlPT9ZaVXxi9brUNqn+tbvxHoRbMxfqT
fWBWKMQGDoV0JJ99YrxL8GbAqcvtmqA9kYhH6o+OaNIwmgGyo0aszbRwTMc1ppD+
1iEO02jvrBS7f/Nb6YMcX7Wk+CkYBx8PIEJkTcdLwRAW5JwUMfmNwnjwXgd9w5AY
EOKc6buIL4f4d+TKl1cuRAC25uU81pUePKK0vt5GyxjMKqnkbjZaE2IqujN2+Cu0
Az55iIAmH603hYx3GQp3LTcqGdRhS+g8nA8kVqMFiPO8GKYimzAbSGZRgoXt27Ru
og+34l/pUCOgQNAsuja0ZuJwgTjjgY59jY7giMdB8e8NueBcdpQ4BNQchNYfFpOL
KE5BAQfPtq+FJnm4JlbhdjIt1sOBziTvpqNt4wDWB3aXMOSukBk0NT0c8SvFbyWs
h50XP1D8e2J5ppQt4nJwjOthafekvEuQqUh+TLqACBO4kRb/4IpbYrG/wGwQ6ItH
AoxLPjeG5sMLrLTx0FHe/rQ14+9hpUgOLNNxGw+sSSjvCb4pE2NdV3XQzWv+Yp6Q
dW2bR2j5//IkhZ8Sj4n5mUZ+p8tL35mA8EKNO99oA+Gtqp3OZHicogCoiR/1BVhU
bcw1SKb2Es6Knd5ri5LwbU0R2jg30eb77mM0yKflD/mRHMp/rqqtzPWJsSVoaFkb
vK8BHQOsgUDFALGpk3kIj+oBptjQNM7mzSTVsHKz5u1hBgeTbWCz+0S4/3AkJPac
5b55Awq5Yr+MTtkIFIi6pBVsj53KU4/dpWkqG34qPVRfmAp/4uUr1cNZLu17w1n6
JqKXoka3SN1UtvnUTqphAFKDm8GHDaA7LsdeuWE1oOisKO6pr72pS/RDaD/NgH/3
nVTtJaMRmEnNXlnXjX8uZjtcq/bhLDNG2PeF9i4Iz5/t/cSOrl+Eb6SEfvfh4jx5
pe577zZOr11l4q/MJ593rLrusQPOhzdvuVfTiZD70AlvcAa0bjwxObBb6/cRAVeV
aLZ4zFdm5FOSh9lff+HU1LcSXxU54Wjx8/t8N2oFQZOabA4j+5u9ozvRGvTYD6lq
ug0VErMkdtdYle0ocIN/x9r3H6hHJ0Eq4mFRWebB5vRfrwc9r9Obag6gTOP38zUj
8nrUMgsvzIhIkG7YilTAQ5VBH2iu9howC7i5hz5QIqvSQhbgjcqPGd8yKxd2A9z/
sQSHRc9oofb6VC3XnY85j687sdXzAEYNvvETq/BD9glMlqDKa4ux0/l93vhYTZOp
hzw1b7PlzsnBgF52yhoGibjeDwPqGScbpmdIZj9ap3kEGu5EhcJXEbUJeMAG9ppl
xiSa3BqRNITvqVXm3wkus6KetvwCFvkKBf2uB94K0A/KfUt9QzZc5FjKs6DQXJR4
DqeUvVvmSVOExksXMTN2Rue5t7ikmeoO0tUt7thPpif42Li5wYm+e9wLz0HqJc+Z
XilZ3PUhGq6b9IQOlw50m4sSML6MgycKcQF/pEDHvskSRo84/TPbilLAW+gveC6p
cwGPddH3dlpH6dO0ud3tkl63mpTTateiFW+g+2kKbLary6mltvdeBkqmEiywj0z1
398roSob83I4d6wL/BpLucCOopB1sdgb6WbzZDJHtzlGzHct4YAhjbMLVD3ns6RY
9PM3H1FKmM04VvJh5zvkq1wTq0G6vz6paEadwI+rPXGY2tWZpvgA/uXSu1mq5f76
vAZA3IHsNmLTGFB/UZlX67wFAAaS9vEV1+ATq0U1ygQNoa58pwFvCIqKkmYnlH29
brwxgeB/RDlwW+Jsdr2rGjnIBRtDq/XvjbTSxi/IKlR0xsUou3lutJKmrhJoQXl0
o/v1k/FNrsEyRXYxeJAZV/EI0+q9JXgp2m4PJu7PR/lSbnCC0e7d0bs8vG6XRo/p
BsTx48bwyQ7a+74ICFQKqn0tmSmU/kQJwYZMin3Yk78fmkEJB0+AIdFIMz6Cco/S
ABp6H4y788na0MtGwNH6IFIe7EAR8lZr8e8zPJvJq6o4icpGu26/o/gKJXiuMd2S
L6YZxOYqvgYZqduLKRGJpp40ng5sh3eadCpyjjGIMEKC2w+5AmPg3O+VMHJV8oBt
Cbh7eXi1EZpCSuM4sgSiDPHVTX0PknPDD/8grnxeGtXoUSMrAvr5WzmE+xZzbYMe
0ANQ1TTogUKDTBXkCPHUZyPzg/UNPwec9+HQ+kB5hUuyWAtSq/f6nQa9SmCnj+2b
//vW2axqA5Nh4tgz9KHJWLe51G4Nx08Hb8iDuyIVInMO8c3ve4ppDNmC9d3BlQjR
iwvAFjoRbxh+PZ/lN199cIvMD7xv6ZRa79Mieewor62KINAP5KvTCPtLsb8yyK5q
jB4JJ/rFzpZiqLS08VV/PNv7qyLvosBvbtSp+5cLJ7nulVevyiN7jC6li3kXLc9d
+4fXr9FvUqdHqPxex9QXt9oamzqz9VKr3o2x9HrmzyXkRPjBzUTIQSA4NzMlc3Lk
jUIic8SiAvng4JrBX1uutxq1idvHcrYYxmcGfPlzUEcwYTIWdLOFVrC7hk2YCGPo
XY74F1+vfsC3zn/z8Ve70D9ByFevH0c1PkevpDPFv/UYpFLVOXRgYx6R353u3+vG
hPjmWM0G6lQZamRcl6Awbj/9BNF2kJJ3rofk0+Rsk3LjlvBih0aVKbIY9fO00312
XMRCpzE00rULGlKfsuVjMdTI5pBVrTZWTMMRLZS1gED07sQyGBH51Vz1zVYe6ZzQ
aFuGNtq3uKeeH4/t1Do0WtG/BSieTJ4xzbxDqIZ/S+Ae1FMxzDRhh0jhE8fKJZ1f
st+yYWrHJP5SfgfbhcoYXSbE1o3+GaZMPYKhcVUZRF5c64U2hEYg85T4RqF0I7G5
AnS5X9qfQsSKUxW49j9NBQczs5qN5wXe1m4QkJqgxe6/f+z3CZZ+KvZ+Hk8gtbZh
CDnz7aX5R6aJAsxi3Z39czT3XMJ47kh933cApqdmWMccv7iuuWMPeYgKBqPFSFP5
AWIMkB9eMSGu2N0QOkLZO+YyopQ5CbTtAWX+Nifu3vzJjaiEDn1sBdGcpgCZQDhQ
7r5oHPzSDnJEFgFeSNorQS4CLqcuj/5Q8VAbRz7TRPPHposLCIUn2ultbVGZJGpJ
vkVMVqEkYxwAVyhaX1R/y157sULgCYSsn7Vs57vopfyI+YJqMY3B9K9GUmj1Cod4
+ZoV1i8GbA1B70LvZpZ6jEM3ya5pmGGMKIa1twe0CnmOh4gr8VABY37dh6m9Trc9
hM9H7JRz0doG9O5nPqCzTRU/AM6i/YyI0uQ4w4JLdd0dGGWac1ZJ99WT4duhcTMI
/WADhC6A3hbf1PqH/if96ccsGxYjA7XEneO97wwh4t0hxSgppkOFNCDEZjTrDYgU
VuhfYXuw88/MwsuMT6S9aTGrjAr7R9rx8+0ykY51LgNdsqszgsQFsIMD9t838y55
v84DK2ejodljbz9fLjWkqGaMpt3iNYDl4odveEmkHERvIGlAcNnyY9NIYgGh+rUM
lpgbK+noL6Jo9OhNe62F5A5ktAPuxcWoikumXcQ07NUR1GC/W9y1cb7yHgxy6J/r
y9BZ7lH1NvUamxic6WpCHtWcLktPNnSGPuROOuMR2uYPb4ZQXkwN6k6VhhorYbiw
FdqxDkRtL6XYS3Rs1ik30ziOX/dyMnvzcUk7tli1neK2DV88VW8hDEi83xiSFNnI
rcjZ87FjhSNpL8vtfOyPE6ltkJ9n/qr4ZCrbjtiPXbOAZZpGN6EQyDD6b3F6b47Q
8a7U+FV74VfJknBFcQWLawy7ReRN4zOM5/e4xnYyc84x/4TxnNgNBkEySR4FOpLk
JHxcRCmhcpy0TQw0fUh2IYV0mxlqKOS4We23hRGn4hGvZ8VOpUjY8XcIybKPbzsO
nKNo1YO1fWgrNDu63vsEXs2YQhKVblEDzuLTVrn0LmXIy7RvrVl/IF9eXE0Pe2NW
yOOi0VkPPuiiBuZP1cHyXr5r169CgpbLAankyHMlNC48tnuEhoqhZ0/FlSIWomH1
y26LIgrxCMPDSeAXZhENKzKY8ZWBR/MNKj2xGfpmAJaaIC38STD+Bup0ZeTdfZbe
8AFFaQZDmOYEJlez+GnHyF0xyjO7QCJTws18WX1/NLAEilkChNLXsSDYj5cv+YWY
D7DIiPyybwQw3PhTp5km4bSqBWicF0Oei8BNYdgT3TxSQptiFZy/3G2eC0UE+h56
Oh55n9hrLa1F1GRikNZR3FuIdszv58FD4+BMaxNZy6gLA5bx9wwjfT2lKRUH8TvH
eBv21ad3vhspyA1CkE7foE5AZig9/0fxISGNZUE2XdhvGO7eXTXeIGVeZLoBrMzP
4qaK3gHWsGx758d82kOx75zq+w1jfTx48pJgtXDRaHPIK/CjahxOJohrHaqapHUH
MSUBHjgBAAPZxD3rF3FnsztTH35LT2ICO5iJWKJYrHskaLlnZ++FKgwEDVL++vAL
zkjOeEWu7Q7NC5vCLR4C4FE50cmpzAhBrhVXphs1U3jwu2YN3kLl73jiXtSThrnn
ugV2lJdjznwOPozfxNiRU/EQVGmCr4CESAQ7mEmaw8aTU5wyTeF6BFwhSP7igLTn
K7NjWWTXZWwB20qOou8mxYwnZAydLt7LzKvby/dj0LvM7jtrC9gJ4LNdg13iRZ7g
XlnSOZRqYfCA0bAkf0Yj3j0tvWlIRinzp/CjSZOQd9/G8GHNeiDof2VTss1bYfiz
wTcwqj5eM5CavSyJyuZnrK26qjn0pvwqudeifLDlehM4hxfPwWOB93bfBqzht5AT
UKMv1plL255kD8W1wDtuA39STquIi0vu2tjFkRQfYcPT96sgVeNNv1T0H2sjm3pG
uv6WFrOyH/mDId/UiHrlx8stNZ23pz8KGQ1cfAbsaKd2ryhBBJmmgU0TMOSqHd6P
uon05C5HyFMvb4RaPmzI1e/8s04YMVmWoBO7W1kKVtl9ry1KqqcP8gsFHfDagfk5
85UzYDKsE6tDwQEmOPAakdNBGJGD4gAR0chGGwfbckj/7sD+WcKo8tr40YP7LJV0
f1XO3ycQSZ61IceSbVDK9Et/Zt+KWnHalbkprtk2IXXLKBYL9335nePsx8W9vgI4
Db1ryr++bVi08UqgOLrUZEAUikWx7TTYF0Opikqc/NQpFpRaeYrHmnNRJZW07e5N
p3VIqTiU/C2hMENGml3VF+J0uE9nEwgEgDmBmCOOV4y8v70q3Xx2PBxBqMm0NRhO
KYAQpdWpSCsTE7cijAs2eZylR3y5m1uzCjfCvShVj5VxwlIPCdESvajgPV6JHqDu
7RjWpzT6X1K2XcJjouRDtjEQm7glMVXH4oEvwsayj/uVSAoEwirrW6Wf7g3Dcz+1
ssBs5jCb5MHz060tW40NXRG8MuzP2g2c9w2ILh7h2/k+hM6p7bW9WWw8AMEFv/pt
S5dg/guNMozXVf/crbeQo5hh3gCArkfl2iG2QJK7kr6UQ9GhBB7YZjyOqXrL6Pxd
NAl30J8yU/o2Z2vuYJhMl4whSRWBUPmUxzg7+mOF1Gp5QcuweKef2Yux9wialVBd
kB3z4pLW/WytgQ7XX6UgCGtMrIjO+Z18uyjSSriThcrajGoY7v3smJk3RBq6HPUA
0h9tM0Si8YAbx6L5dnGgGMz9xk++bG/+S5PJy2JlmmNKaU+GXvkxnTX1Phk7oCrU
4WHGEfHgLMuUfsXpOSGPWLVgk+Pboe5CkEuPhY/7HdPuianmUoVOW+LgHr3+TSn0
6jpttq9KA3zdgfSSju7rnWLfu+BhLV1vWcLvUZxmGWBzzinea9iviik9royuICZ3
+oG4HB7m3EV9JfunX9jx0p2aqzrQq55uJa9/qz6g9GZrKAFSzM2iafhl69t3O5Ig
RDQ+CmcHxgTYbfii4rXnU0EAMj1vG2jFo0VA5tQJP8XrFQ95GB4kTH36BcomyV07
vKUMQoCOwT0ijMigzZPAIvGKZcSnbFI7bv56Aha2QEHdQwOIWS7yIkXfGYme5dVN
ImbGcEzm6tkUHObwB3NUzlWYMmLPnXuBUW+ZYcLHz3vg0tDddN5wpN21t9uVMKXs
ICnfWK7cNer0hCHcT75SqJrRYnhhS3GtaWQzB9ttlxTm7bcekws61RYm7ACazEto
LY/yBx957tNeDLZTB7eEUvRojLJJipvt1gJstn2K6yAGDE9K2pbSrZx9H1owi/4t
bqdkekWHaj3kVxIbbug4orLvqywa6hRns4gjFge6ewxROSknRqMwTQtOJLk7Zx0C
wSnx5jLjXzZqzvNjQPoXOpRphCPUywpR0B0AFwVhYiETt1VBzRHiSGq1bzUZa7s8
3ouwbW47cb0owjdk0TEqTuK91bTr7iXNKXqfLJwtCy+28HMAZiOs5XyLzjkgGe9M
P7fGimdQkoDnOdKa1hsx0bAJ7z4VdMJEYhZfLH75LDvzMFjjesW0mlj+GdRcyagJ
zszzDaZ10U/or62o8P9eoi7CdmEuJOd9s3QhK6HqJNsMwdeSjLJIxzn+Al4nrjcV
/qRPBgChIWvjGRv8luqA8zKw47AQleBveLDlYPup57cVup3vR7IW5sY5jsPkdrvc
14C0ha3h6zK08954kdnJbm+O7x+V6fVKkkTGpmnaYfEHEZyW9f13d2c+zujcZPsP
YdQiBkn69dXJdfevM4UuVyqYHTo8sQl6Wde88ED1JccvHV9Y3NTRSIcbwymOKNNf
VbgqWdShiT5UraSHe6iVwAwe9/TIExEvd20BEDajdnKT/F1xriEyC0zOP8DS9AoJ
HXav67Sv9D3XleuRpdWrYvoTUpiFUCLNUZbvFPvITwru6qZBb9E7ndHKcuRy8n4u
kQisxHfkowtPx2QgaC6dz3fBZdg3Iui2ImoWScBYKjTaXhFWk9q+j+Xyw95rh1TX
8u4bgucoJE1Z9MsCSAI/KoIifxORaOdAit6aiFOZn3Tjm8WkC/x3+NqoVwWqIyZU
xzKTyF5fdEMT8mV1L9Vp5DL3Eqjp5T+ycVLyjJgf0yZJAjAC4kd9uewXaA4oGprX
72iu8R4w9pqCG7qmSBQHLygN7mmsfMTK3byhBc6e3ErmHsA2RpqXg2oHKxNYqIIp
yQsD42FT+O4dTs+hIjKrwNc0RsnktAut1a1wcBsZnMQbOQ1txVnTMgmdym5a3yXM
50ahC0y1T5x7uzr1ghDuIb3EEQxM5wwu7LQT8tRM8DZptewyw+mt4kv8BS2VpHlA
Qs8bDd3uQuuZRoXJ5LHtcKkDpOr/VkEyEtENg26EiGULx516StcrBE/7z/biUR9G
bxgBm5BTL1H8PNieIvkNFiqThhD5YahVBWe85gLLlrDNVZgKRrxLbJWiRXaIHzCL
mgFVMe6CXP1VDnZmn50xsuyFR/rzThrnapNUKP1OZeW70hGlo3IqKl6uPMb1iAKU
wuMeVPYA2KNE6ZLi81hw5H+DdTzaB5JL/HFMp2/ZpDJ8G2jQVIZ2kRNt/JTFx9pz
A2Nc3JRyPjog0gIsmnNQTX8U6EpwDtXbyOkbXdapky3kVSHuo6LX7jsq6bu9mI51
r3qaVZLL1NUzv5p6rygkj4i7PY3f5XFkX2UYFiYG4kiIK9deV1pDFypT8TbXOwia
enJuWXPDQu/ejSyZjZ69YKr+IcP8eMtRPzNPuDiLTDTRvmxMVA1VrFfw+89NYaAY
LpQxI2eQqRpZo+buhajE2csNgWNA0WX0tO4fQpp6dqpNK+LcFUmuK3iuUTQ2nxT1
psrlvRNTDeZnCHnN1mtuRtI+onVo+OC/pU2pmgmWlQekZL7tjA7jxLvfuJCg7ryA
6c1cuHn19XNmkpN08W2HsD1KQYHE1CHYDfN0fF1BH3/Tbzb5p9coeCSm2quOrpcZ
p6ITwSeWwFHjzwx3N5AsFw/ZM9c4Pycrj3i31UUmVeANWstQwaFiEtMOYidd0BHQ
WKF6/tppA+w85sLCBQf9kEpYIuwY4mLtIiO2XX4YMI2IdzeRDJNuEBWJ00EdVFv3
dkw3aHzn//xEgudvjzPAN6A9J5X8EYXLrskXlhviIQ95Ny0ZW7AODnFEN4GNt5+h
J5FznkyAqnp5Oz1xH1uiOwnxt68gGOyUnER5WdoMBqP2tjm1IClefFstViDJr1cA
0oI0K429lBNdMM+CGEhePMp150wWE//7FlQXSX7vCqLWnSn+JT68dyYO1V1tKiaD
DKCGTXS6tLnxw+CtzpsFHjLRR91z58WTudtnKYVzg8gqGooZZMjnVET1zK3GgfUq
PZ+Ke+TvUyvbSwvAjkLvKHv3XGTF/MuWis4sqZlcCyjnyrWwoAV32GZyUIuweU7V
GR3ncWeSBOlG0T/+76nhsq8HsV7be/IiGTX06mIW71cYUvLifgeHlSbVE79zaqXw
fWpjKd+jwkcZ8jIO8DC3waq8YBe5dpj76OpMsuC4vhJTRMf9I59n8YpKR7Upi2GH
eU2FmiecDc0L+njlcFl2Cc0K/jae6+HDyTbsy39oVrShx7u7cfwyW+lr5lVx42IL
TytkwsZNCrL9YLdAGogMJNyY0SMRd3gpP0KPulomzneh00NjRI8CanwB7Jm2vcmF
O876yT7no6PMnXNLyLuGj7FDW6mkhtX7vUF8xai42ZVs0HX/GRzTX6al2Lev3SuD
eZCn616DV5H+kc4JEhtSrR1PaojL370F4t9OESmw0Vmdwtoc3+alzt5c8aQEcheu
V9ckXpsJ2ErZ91LL/mar3z+Wz09/sq0iDdkePZCma0NV+he0YCfszp9nF7HMXAbH
sHOBoWqaptARLJm6h+S5NCJi9Kg8Lwy/je+3Ap3Wxlm6Y+IdI3HllRCd4GwUFDv7
vtnY9BgaR/92G7GRl/F0KtTGRsflfjNnJ34MmhekGEUWDGbqf4QklOz6EpN2wwQG
0+84ShUtA/DGhmc3X4rJM0TANyeivYvAzHfMFi5qrWK2upmC3+Q152TiMZpw3as4
2M4oQxK6ll6Px2+UAfxPK4kc7Z+4fjAB1c8myM8LYL2zlCIL8EDoJnEqv1TUM3MH
aXLjsFcgBRCUDCxOBurMQ2wTQTrioEPNsPMpnCiK+K69c9SAxHoNGe6rDvTGzlnF
bwvZHM3JqOGd3GI7PZLE8jFnzXWqgKST73QeMobsNAE6R/o02EtTFtMV4m8KJsGH
+y4mQMx1Qa/s4x3Ly/Ty7qHRfuvzMuG4GpvcYjkEYhd1HKUoecG0Wr+kYFSlu2bg
wBrl0fpl6YVcksSi1C9utFfjUokSWlPYCmuBPB/bYfSIP0AYfwkvmrLPEtD3iQVi
v9GlJ5kvK4Ef5dF95yO7CSr9SX8vSxYU7LdzaCXt1y7sXWtdUfgj9OVXwcIHbAkC
HyfNO06Z6lKC6dJCe/A6H8+JunJtzWuRdTuEbJPXV9+XqpUb8xQ70wocL5983ktp
kG6hmJOTCFbIOOkocZKKaG7idqqdNUcXDBbjPG9ahppDrpQZMkvkuElnyEx3UDwK
EBm4yjMXGqJPmzFY3Xk32TIeqR2FZT+HNTiEdfCgGfpM+kUMFizji/gnkhx8T9c6
Or6ORXn0XAsPy+k4SbdseuSssUIZqreggP+QsfI1c1oN2U8t/2n5ebFO7TSkFD3i
/+0F3Fv1/oOmNq1MHqrDrbOHDI44B+3la57a5ytHfl46ReyY+ASYazv5gSiMJILh
8W/ex7mqVC8s0LPizrrGePdHcHLhTNZnJMQvnigH5o45puhnpqyfT2dyw1rmtrB5
LjsQG1vCTb2YvYgAmSYXfhz7OrTU4yS7wmXcrqtZxBv/EdWMFqDhhSA+3hwGJY27
BKRqWUGeQCZxcWS5h6i3ahr7W3EYCIlA8xQrEaJe3VeHwdZpky9oy1Kbdr7FoQSv
+Yvv6hgginiu8OQ635+IGMdoh/uoomn/Ows0eONucns7AzmdW6fPEdpc9SFUGjI9
bpMIt+m8yk7qx5WQuRMxr1039tvaxfhtTfVN9EIfehXjgYf/qgyWuDd92ju2yvKn
SxfWI+J1PHaOd88xshsltTYkzmApUiATGCnSh+DH6vVBN5MCruCJ1X+/BygrLu+C
Hu09FNnBSiCTYaO6ePRwN4eLMXTi06YS0IPtIefjfYLAUsH7BTA6SvYn/PmwwXtG
MExvDqg7r/P4SZFnuJNY/lyMQgHQROl5Wm/0dqGFGZXaoCi8NH0UjavvZwd0/Zl/
r7++v5XySqbku8t+13CJDIxvs4xr9tVrHlOsD9WewtgcoLZ5kdKyqVTCQ2qg0v3Y
gFGgG6eyZtsYA8uMXOaKy+Wgv3nx54ZWaBwESuB2cz/BJpRHjwB3jhjTEI7AvBvd
Kiszaux40OpSHJpPf5QeSCmGk4nv3lnTta+wa+0x/PqlPrHtop7pYlIgTeJHjO2U
b6K2GgQA4xyesB9CAfGgI0D6bNgWM8GM2dZ14lQqUuhhS4nrNFES893btDrg9lRL
8n7rwTkLiEFHRPWX7v/d4xfFkA+WdP4pWJL6vt4hPPfj0t23LVhRzueRS9E4dymN
CgvbFMUPRKfNzW2HmUjbDZRE9RKHDOvNAYFPClrELFG6GiLhWf4AEzfnfCg23rBZ
d76eDyazx8T4UFSxwpYXcJRJpjPZ9ioF/xmAV66TL8/qDVmcVhhhy59DnD7retj7
XXUu1jvDSHv+eGmgOE+osL8E0oSOI3mvR36aqCFZRViWe7UILG4Qd/xMiwtjDdKS
cX/3XRT+8aFkj75Xf0QI45z9lcZ3FqDM+lXQvU4s94FXFPvtU4llMKLkALmJo7m4
6zzvZPYXc/M9kC7Ag+gWK5N1rE0BcqTWK0RSu/Nkfz2xF1S4oiLfey998hqVJii9
KmoEtXz77Cvnp+7Z/ukOUFNUj9oW7IU1XbwrcYSWLTMFx26OAs5GhD6BrpU6uXPZ
rlSmnS6k2mpa59iZDmC+cTy9OV4/TDGn9aNu696MUYC1HjSYqN3mbF3bhfLYzc/p
IiwN0gvx1QcITKJBw5nVniT709fobrW+J9jcyhZt4G7+2HrRXvAevHHXb88fjv+X
QDptHYiJTB1ALYUBc/6ZNox5nAYeihDhcDQaSNvaWJcYQxeR/RCDt91MUCyiu9tX
lG6EzWPTPLELnACRSAeCTJBZPC6e3kCeY91UIgHxAdKRLqlPcK0dJNys6ArO/3O1
MzjtYtZNohXezxm71/kQfhHEwT8qk1kqOhToJBhu+9DqoBBKWMyLsCMP35nT7TDQ
jJMt1fpWpNvC2/OMB72WjbszFa7uVvm2Rbjnhbgk3TsPktXrmEeZUkc+KituaeSz
0zO4jN+t/kEum2FI6slMMjH0XOH5eBavyIQl1IQyd6WaGJVl4OskWwsH3BOnDgIN
eQOpWe7svnRxMD5ID6kY0YZY4EM0+17oWMquTT1yynPNJ40NWQ8fv1OnSAVD/NPD
0KBcQeDk7fvII5rShtodCDESR+T3GgWFqA0GYfGKr515zZVBVXgqebfrUXlUKGKD
qB5Aw89ogi/NFst3WS/XzErtXnc9EmIGLtqcrilrmn625Frp6ypsLwkjcwxqvkUC
x57AS8YaQEvCAq/y9lj2d0TYwFoFym6cdlEybTkhwHbWx8/OMA3LORjKZJdUmnod
ZwY25+afsZxg3pagwcbDOHjjBeY2nBQgzFsJx0+lDZ9PCMW5R1aRK06D1DI2wdZA
IceuL4ePS9/pMn+yaPMkF3dKX9TVkR1wFQAvXn00k+bvYfdV0pNv9akjyNkWqeJ7
sIi22e6kY0/X8AGjexDcVnXDYBXWlt7obE6iLxTabPLYgZtQL8OYNkzVcWsYzdvV
Sab3X5dFY1L8jd6AfU9eiTBVUydqyVnGLVgtB/bEMY87Im/gW2m7Evx1j5cFsvb6
9ZOI7M/5g6uYPEh8mI770w8apKje70U/80XmV7wBzORfj3U5fH/B/1oSLQwoYBku
fqQhxWRWpnFo27TJBKB0E86Sirc4qxa85NxulcPT6OyVy2kUH9xYwI2Bor2TMdFO
fPY5/1QXD3hpjyP1iyI4r+7wTDnsDd1acj80GCXduoCyTn+AqB6UrzA4GHxrYHaX
6NNtQxikaRfZi6hxEOpey4B26s2d1azoeSLNtyleIGt4vMg/uVkdwU0e491ZJ1dT
krJtJPFoEqbepBcJaONEv+7WVwVrPIRfdZNimSJ1n4V2GWbHLOpRhmCpEAJy/34t
uHOogKNT1BEUbT5nqnecI7L692jMry8vX+iTUCvLjL3NadTaougvcZamexVsNpKG
jce0KwsmGUZ5Qp0r9RXeMklsaDwDyDzN1K/7fqsIgYj6lVR0TtgCHSc0VwUKWlir
2TwRau9AWgQrb8467IRNdZ4UgUp4yByuG3VmeH8w+Pti3PAhCJc1P+P99k7aXEYo
21y8gwmEZh9A2pjKuFYa94UZ2SLLKY/+w3aBvZyDsObmAqjAhAoT7iqQCCHC+UzR
Ha3jPzva+fWHY4wjR7eU7YafPFBg03PDkL1xwiNf69WQxBZkYtkVd8z90rRYm+ME
Cs3PDx1SfJPw5GKQ7Tbx3YWBUqiblC0QHt5KJPcrt4V2O3dyA0REHY/ZKt82egZ1
Cs6jKFaQ6SmHuAuNVweP1BNNJuT7piD1VynrJDvARMbUV4uiisaS9zSEghOJJ1jr
d6a2kmi4hp0ILYYOVqrGPMAk/beBPvZe4ONI1mf4ZGSUxriRLn8uYJVb1/z3c8s0
DxWGCj7HUjleLSAM14W8gApdt6dQzwmOm3tC8SHq3Y9n/wCg+eQ1Q10wy4J7zUvs
wYEYJIU6fYMGNWGGc2n+Ap1LMQYZU/CT9Gt67y7NCBVGy6TGNANk5/uoieK2W0//
tYN0tcZNuyJG0fWuxGvba2fYypxPKidDckHEgW1Bk1tqRMUfL+CCWVATxwfPIVqK
/ZtzJqKMEgcJpf+pguic32+YlIrdoUy4CUjoUgBBsYOYcAHL0/lBq20knuIVzK/l
1O/x4AOV4ttsyzMs3t71m6t8wEDx8xJHamkfGB7fTG4S1aXkmEX9jqgqA+TXKLAE
9zQ5oRsWnGkP11WyQ4WkVeLjAahH2O2CrfSi0dgbwoJMCRfFTVnYqWa3DLeTEzss
t4DyRb+MCZsR3z3Alq9ucabnqBdlaYo558fv8v7sBTgALhytdM/u6IPFJcbHxOi9
AlYEjvwL6nu6LVSIH+Uft2f52xOO1FQAbhaZqN+5x0Bi986e4DA0VI2vQBBZhQ+O
hfKUHoXjTw8anWPEIGbspopJgwHeWghnyGMcN4DhHkgzBjriv9rNv9ILwDupyBn7
z3bkcUx95+x7Tnck6FnnaABIx85Cb8tzP8scjVxXosj+zekYvBsd58zS+6tg+lma
7WHRsiLi7//0vdbnlNNZ6ZC9FgFrfwBUOk7BAeKyVJ7uBZiT4X0119vCooJOjvx+
8OUxXKsf42N8WowgzzMja9F+uffNVZefJJq5anhMTHaWm3fw0hTWhvWb4W4ogNvR
/0u8keZo9WkJAIowIfGpegD7oSXBqyLWL16a8D5jQw1Eb24XH2pQxICGstOCFbdf
LU8kLpeb/n3/pWJaE3pMt6fZ4mQ00zvaughhvX7wB5hWhU/LYkwKWDiMix3XZGnl
NfW3rC+p47VpxKWfPog2BI8DSzgngt5dIIJiK7q/ukt41O2fgdZ9KOcNZPo+Rr4l
KGewSZF34q7T+wImMwr3UJgBD4XZKYKJvOSWa8fcCwg9BPTISAlgiBjwgGRxK79l
isEvfupo3327K9xW/rCFBBMpwjHsPB8ftmDEJPqBfEUxgGcDCPU7UqXf7dVotBjZ
4MX0Sw9oYQjF+a4UzHBkq6ZlOovxWIOkka3hLx6VNgPTzUIxqqueTOhl2t6k2P9g
bu0+ZvARDx4JZ+CUc10k3n9HSkU8+aLfsB30dpAwFhDXTSPoN5XJbs5vJdLYLxbY
QVq+6Wnp9Hfuv/oa2B3IYDxKeRag9OOZo/yt1hZpOu6bYUrZsBRABbmFpEdUpE1X
aE6/x8HHC87K+h/Mg7jlfq3KyrNgUv37P6Ty4XqKSq3GUbFZi4pllN5hZPvupc1G
tvGZ3JO+C/VyfF5lLZ738PhFemyaMuveuuapyPMAkxm8W+MuQikgELUgszjfLOhi
Kj+0LB6IW48K4d4e6g2DfnG85Trbe/buLfrnt64aaM81QVlYa5ekMZ4NfA93yw4J
QnR2BfAKqiYByc3bXKmVBwqSn54+tFhNNmKAvKVshZBmMxaM6QmyWeLUPtc6u+GT
vudto7Q7gwztuLnVal/uMo1AAunEgvttN6jh7adMvnJBdeZHAhJp5cLQZOBgXhdx
whDmYVKJR9brvUBehms6z33gWJdhAxgYs7AFoKUNcbLojIYopRP/mSbIiEcefj6E
zpNIsf3gaTsMlA8VVSCeEDphqw+tzAJPHkSzMAZx1nYv3Nusplm1eOpKgt75autg
KPdf12NcFaRt/WFC5EfP79Q/tA+tNNBNAX7+liKugllVGv86eJLvpz+gvg/LEy5y
JWHVd1Qox4RRKpVeqMd43ZMHpc6Gkg77wivM+ojdMbeNlpPNNTeIJYXz/y9Rz51X
3gS6i29brgucoIxXXtWydc55NsnfnL5AfKRgr95A80hgHeR+yCDEA0NcuAx1qck/
s1aO45SFpk/7mHyZwCJD3XLlBD6kqh+OVp+ZoIykZq1mGgwxMuOxskEay/YAlR/v
wlLxE11wHNTQKMkir80OZU2SiVx2pEn+axj4JPDWSF48Pg04RxiMR8MPDOPHgL4z
gdP09QItaILLga3oE6Wln9xOwwCN7zPQek7QgLhIXwIThhi8R0QuObyH3UZfMEkj
J7ho5s21oRkS6zjeMtBl3nbD8uA+9iijx9OCUEyVoWKNEzXAa1jerZDpwdahRpkU
e3LemCg/zw9DKJe/0AFKaIoomm0SngWfVxv8bsWaxv16gzR0Cpa3gWBbud7hObsy
ypsz0//MEe7VOfY1nURBnQWbPxUgeSODQxT96SfJcCdjmeCryD7gTSaTCGrL6ZB8
TaMi4ZH8IJ6szCLfjYOlgRls+cav7MujhD6QFeBo17Wqz+s+NZe9YYrEABe1n8Dn
+hnIDpExa8eL1SRsYFj351iJj2n7Dt9Tgts0AkUfbhbr49yUcqumvM2F2eravg12
HcoUHef7QSq37SKurliqi9nvV2ucEjUOQaUH2ZLgVI3gzzBgYlw9cFLILnGXbPC+
5iJ4kVA9gz02sPI+DP8nZ9nThwotO+5Ut84MdFUXy5kfAAUmL7pWUS+6RiqqucZo
cCr7HYVyEiRBIPwt0Z0pqrH+z+yKBb+cEUQihc/Mj4SPos+PBIxFjyZsibprEbyv
MEXe1BlsRhqLb/eGj/ib5W4GB3geduQk83cr2O4HKYaw9icSBxmmvpMmW+k/39lo
9mqqcjgIHy7JdU0tQcp3jJfV1Rzjs9XzERJizXkC3wauV842jooYbLu90jZBpNoi
H2xsqHy3bDJC0XbX2+V95um619VJlK9Dq3AfpOOWtuHkeXGKhOk65byEIcWEwrdU
06S50REhUcL4N6sVKnYOOMtg4qY+q788gJvmKEuXKrf6SL7IXzUxSN4yL61kMO6g
RyOByWAUcHlOHQtepeEvwFrnO8FO7TLQqCYYNo3TVOgbg9RWF2IJOaTIyWIoKWgx
ljoz42LdXE764OfrTbB6zKb5KA69b2Z1H9H5gejGxFt4h+oVLakG6yekRC45mzIb
n7fdgz5NZ1hn5049TgdBge53objHaJYBIA5I1aELsMwPjl5jA01tjPBHGuTtJnkW
KuGwQt1zWvrJ5Fn/sZpXCkTrhIcXdbxR89SaAk9COWRRya/Mfg2U7IqSZurigk5S
MlKsNyMkgGU5T4xG5pF6Nc6FYtwJU/30v+BNxCGRHrJIJVlB74Lw2Nzapb7z3YBe
aJ4Pna6NKkkt0ZseICp5xTsAP01FOIbbR7w9N0D+38NFrxSN3pFlPKKXiGIFT8SC
z/yGSccyJ/Vjb9BRnUYgkkHSL2saN40x3XcpN0/es3HgUJxrFEssxSQKylVK/Lkg
pBQs/xLpZhGhzMYIAY1hdMee2UnNvGubPbK5rj8xH611N36g63mH6VbKnUhbeNOj
KxnyB4t2FAVUxtWPzaRbi4J8v13A41cJDmAZ/TiP3FP4jsFjh80OxI2xga3WdJ+b
p0qL6QS2rgRDmoxT9u8das6IHhQXavXqGTyMZQq9vr+muj3qwsqi0PTJ8xJwIN20
THgcODS7W//3IBA0ZdWJHIOuqFCffBBJbZY6WchKw0quBbl96Lf7IRF5m66nUO5H
V7MQNvaGN2lqyerFFftLFCBizCIurCggzP7hSiQDWYnXB9YoKDrMrOYzTRgB6hO1
sOGxFpdeiU5Za0wYHOMTkQEeQ5hU46jhEZuhE7Y3+yh/ii9LIhEO4g+Hq1nKVaLm
zpT/CtBIdEzeACGLOa1be7+eTQsPdhGH9bbEWVuzrMibcwmHF+5JWdA5pUzcgluj
yedMSfK4oY/Nocqxb8ZRpFGDyW0+LXGgLTElwA89bD8X082xER1mx6IWphu31A0b
7pdZIBqcsYe6L2eR/baJhl6uyU4vdXSAyLyjUQnXi8KVrFlxFFNPH73BBcpdP4Qx
9Ra5fTXPUycUauviZ03BIkQrxaJaAXb7StOllGckD9tjRTk0fIEDlTyhtNihtoJ8
exXG+aoi6OzcnaejoiE/yzZs2iTw6gM1SP3o7gfv1HXgl5PzBZB4fhJ62FjBLbU8
6B6vXGx410S3kB+OeAhYoZkw9uByJu1wFcCOsXeJBrM1Ycc15XWQlow4MclEQ0Z0
/A6RQgwd0AnOmHrKKli/qyJSGQHKsjaND+p7bMWdxJgA1yBOBvlud8eeHlywqhmt
GDV/7BXT5wFuQYh5MrjV2OOJgcTOkAropa1WEQeqnu9O7GuvSkKBnlButL5Xlrb1
sKSy7Dm3PlqozIMBKiCos6qZa0eXU57Wq7Nnou+43zL+dCtr+HRJf2OtyFbCCsIV
/bhIuVQZV/QPAdpOHX8P0ge3ma17FrQGOvYgj/kNbXQ5n9RjoeSD6Q+GfY++ZjUX
/nISWDoHjgfktVi6D3jSQ9sEz8ZFnDE2teZ9cDY+BaLGuAuP7cIio5Wp7xfFGZWo
tRrwNflmQfpsq2Btoiog8SSQtEVSpTLUw1UZx1p2/y6XJuGhkQEsZdGMZud3Klmk
e5uY0zCdsNc/8/wfKbPEnD1NaRzy0f9UC9lo79cUdeRvaabQ4+ULGT9BsB8XtKzx
xYXw7QtVdTwsbfxd4jFVcjBkwFqfKHE3U7Lm14DUImpxE0MkJdiaOIiz3gxXaNBn
S3jWDv/j/fkx9JXwEsTXPBtror9Zi8yCbuE/yI9m9X03H25/VIca7xxAhx6K93qu
jOwlV5pbyXPwpT6H0Ltcv77Lc8Orp8I9yangSVKyASzf3GP6uBU2SQF3nIN55iGx
ZywsXuB2+sp0GsPzhiKg59UsFatGNgxvQmD8UfJioC94Tx4nilnu3nToA3ZCs/dH
7arP7ELitrY1sw1oLf95O7H8IM2PG0c7jakepB0Spev885DHNwoiZX5IW337Fd90
8VGc7r6BZ0DmcSBIIrm3GR8zDrv/OAjvXzbUnflgPql4BRpzoFcERiDq2NdiqwgV
CXGIkaSrhES6O49QbL+5SoeQ/krM3FeXVGbiA3SvpauHmcZIvMlgev2rN52pWsqI
r4HEz7E0/YZrevT5PQFB+MOAUcMtMuArSQcd9A8aewYbD2EDNfyBGnm76aJZeX9V
Sf04fWlebCU99wl/8Uh/ysFnmWtEH7XimX+f13tcDCzwc2oKwbnsARabUhwh7ytg
Aq6Zx5xGAE/ZNf4+Bt7/jMdhBzF7oeW0+aHf3KGVFRqnUDpizW8PMeJ5hjzNS4/e
hbRxkighOVRmPt/2vHmbTmMQhGoxmKKDloA3ywFXwStsFip+1wWL6wVvliOQf/yx
g/24p2ObRoiUMQb8aubl0k3K8w04RuWETeFkveuDU0GJp+V45stGywew/Jg8MUHk
YllAxK8Qt9DAjejL/OKt2R8LMCrrFPi/8QFYv+Kp6PLSoEVWY+75zjtetKqtv5aH
MGydYWdS0Bp+c+3zBfyXIs+aI7jto7Sifmq3v1nE2CxOp9qYZk513TSUke1FBgUF
s2m5RshBQMmDXy8rpbezOkBMVAKlQ0XCsO7vK2lr2MUIYngGTm3+HwLG+KGiAkhl
0dxdKvoV24h9Da++kVhtgzDJEO2oHHS0aYFSZHRh9FXLnjXPX7b0jHtObtwRaUO0
QxBHQXWRvJkV8Hp2SXPwF0cNKEUGV+eVM6kGs0BSH3RRruNZyD4q5W8yXytbil6a
EbOTU6iMBxJZHV/nfF1m+rdxsGxW00qmjjpTmO0/IzewGKIQdXtGgJ2qBBYQqgX3
whwz0RqmIPQmkbWwDUBn7v0wndbzPVqN1g97R8UzdmAC3UWZ4aFgcj7VkUMeUGcf
alCYmGPMt+x1EADorknpFh1iLzjjdPr7t8RFD8t+U/mOBbNVHag/B/OOo0wBbQqI
2S8GLHE9bXkpMw4U3P2MF3P03UNa5bh5xT/ybV3LseplHqftwmGIockVxAjCjGwm
XKSd5hD5u/siRzfu5PrYUASHtDxEnspTVcEnhxmnSEWdds5vje9EP0oq6s0jHft1
LvFEIpS8N9800JdL2WqVSL9aHMIYWwwHh75RuSZNfVqrofr7V+R+qge8X/fTnLki
0LLFgBsQn0nW33+07ahCRydHOc/WCC2R3mYEKfaz3OpEqD4f1fpxSKyGq4oikggF
X//zV9xU69oSEGV68L5a6ppcfG2m6yIvWnUT3E6uHQoiXNtdjrTzIote9sAgvuLr
1AUSZRTFNhqIWhVQAqss9NpVaspnkZLheSYSwuicwR0cIB2awTgMgC+Dr8VyA70S
/ap2jiWrlMxeqhfbxuLodI4BiqWyoq3xuj2PJ8VcJxhKg+ElH9GlA4DRPsPeydRu
aOPp05TvvUqBsqgMK5ahZKWvKtPUKJLLEe+t+SJGXU9I4i2T0swNQ/nOZ+2L6M2f
MN15Gt0IJajJ63qPRfB+1TcU5zlobx34x1CrkXPk6fshMm+u+15Bdp8Kt4Snq8tF
KND4w6E8/lXZK0o4qGD/IHT+vx0vt6DgE3H8pKGcTQyEad5WLNja5I60CRwbEkAu
2Pm79yTFLaRSbcmfEECbmbf85mTLk1KfAWVwP7DD6vcpafoYTx5obg3SxPJfJDQQ
fY6Ehg6+YFDNiHQWKjt4XAz+WlkfJlvBM3tJVlgZzxKYUeZLg7XQpRHZXXwcOWX4
oZ1AjQ/2a+Txe+tX/bXjVtxd4iMrMI+Hy2GYZny8arpfRsqfAqBxg5UfhiZ5cMdV
aPTiQvZGgcm6GtvJ2Q2KnDF6zNuQxip3evOQty9frSRXsTIdR+pUXAmltroqt3HO
bwMzhkVMKKMJFvLsdH5mUGBT8dIx9332jX5VsHqWnEBjeF0jH9+okTwd08Wns8br
cgp/RQ0y43BaCWDslFrAN3SDT4CTb4qvpkGumWgpcu2P2CNIvuqfnooSAAHb0DY1
es0t6P6L6XIpy5jwbtKbQZKV/6ZVza7XwqbkVt8bW6gquttV2yPWfXx53gElvLoZ
3jnnGHiO7uphXaw6NFotP784/EP7uelUyXezv22uTpQ66GFFxQoTcVjuX5J/XdAa
5AOhH2VK62MdzlHAnwK58A+GhcZsz04p5oX6tUSWCE/g5Ojcqo9EHXBGU6E8MBr4
EefMNMHigrDvqUmmGZJSHYYDfl0fyzTHC/ysVvFsSavE8R4DLq8HE1DdbOCN7kBw
vWhiaeLNOR7SUlavvB5G2ZrINj/RUDh+2ucAHAY7qUUNwbtU83uAMH8P0z59IPO3
F6YaEWegFKNgv316uWPx+fWsuBU2Y+2xUAthcMC3JXzUQbkxUdwtqgckcQyUbXCq
X/4M3LxOgQis0VxUTRIDQEQOOknzd0vSWB4XfjjLQaU79K5x1fAGzB23exVSzoxY
1r8ZP7IJFRPuB3Lj05ZV1qYHntRAm8rNjdARa5jx7oav7J5qK+vZiL2IJVVQ0hAp
tpDEGVnnLuBCeocUVGj2+AdeGvEADeeZK7kgBxVVfjjmkB8tC08FItolvwZD4aNS
iA46JteSAeyLL8FV9CijpGkBnBKPs1BobGXfcGjnBVK/0aJJj0KF2u1UJqAmhL0w
Pcbwq1o/PN/v+DsS3I5eSb+pOvS8T1enzUAiT6FWpeE/zh/MWhquCMF4cyCreWWM
tapUQ/YFSzsaA2FEsn0d+/Rb3poucqd1GmWrWUq4+BP1Sneb4re25fS+DtvkWQUB
3FjLNwa54fG3QPYMGQDBZJZjCcaOEnFJ8qtLS5osfFppyabx57DadtkOsnG8rFUY
CTXxPLUV35Quc+lMbkLxsSi2i1oddIDoHWefDT8oTdPBBlLSfAqQ27AOBivym4Xi
2SQqZFsKF6A8TOywpifHLKlSXQ/lub6vTLxpJQI049jrlbeu6k/uR+31yQ8N9fz9
eBCEkh8mS5cK89Gyx2FuGob/JOQvkUL0GMxPCZR99F59nqxS7yjGZ5LM8FlwwDho
9DDu+yNMCsATSQY6tq6+0xkLh7HPrbgTEnWRXdMYZUqvVmSlSkYDeh/32QZwHb35
FYDK4w9jyYXoLKSVMkigM6XeBklS3YdEBE02vm2tbgylUy+3poXeWeEIUUWCLF/H
iGDDy9ZJiS0nLdDsu786xz4Rx9Xi45EdljqaefMgEJmE6wMPUr9x7dBRtEUuE4en
573H9l7WSqW8Pcd0Xzca0kAdEv3rjIjTIBDtUjoEx7H6GlzjkSuwOeMt+iVLfIIq
KBYEx9pv272mEWiWSeETtoaCsvk36t/b2lgMgrHbw32zv1fczWOM/xeTzlRjJxF0
WzGAcUwxmn4ofzqMtRJyp42V70sfoVmZ9ZUdCeBewYsPkENpogrpTgl9rm2s4T+6
36VzhP0Y24SVyX6wwoY5gmW4CNRiqKxgFGW6GJBQirr7bVWSI+SLWOZ33dqMHgTo
pFS9tieQEIX7tcOOqlm3Kfdf8M5wrKCq10wAW/RyZ+jabfSXMvNFR1F1hMp+bzdT
koGkD6AGkSKVf3i10zsxavpbhl4vaXQuA5dGtRkWKZpUp/2Njmd9kWG6TliiU2d/
b3d3lydQFVvNfUPzYOZDxBZ4jDYnKq/ohqFjKXzJDkHEIvpVvicfuL74cz0q7ep8
xfc06KXmmOP1woF73TyT27MssrGWs1/P20zLRSHFET2r53pckIbdHFrSE/KogMzX
iFKD3JlKPp6CVCPNJoF8Le8Ll5Q4badmx7RNvR/+0rndVzidw6A4ucrnDVB+genn
9c0ggC8Q9ufXPMnjEUvfBhTxrgyarCnd4cOP66VNp13WLVpkVFt0Wx3R2VyGvcud
6uoBmHMJK9jDxjbVFgkmZ4skKwJFTPGOIZn4+MnRoKL3iKAC7pgA+ZtnxkI+I/fg
ww4hyC1yZH/nUjW4vdef7hvYMTmgXd03zq1nKYqciV/lT72Tz19xb63XRXpDrB+j
Y9MUug0POwWjfvJZ0JFMnQWNsSW1aHfabmd1FMrIOIrFJAHe4o/M2FU6PGAL5wEG
V/S9RLweAQUxHRBTFiF9y8Hti6sUjr+Bz9NUKNEpnrR97lMyGxFw1lHL0Q2qCx63
KBllviLD+1nurczbuyVw3zTFmh11vfiEH4B9svmhhcKgqa1Rj1o0zp2Y3k7fS+dl
bhi6gkGApGd6jK5nY7w4DLAWS5rEHeIslmtuiH30MeDV45fjHIkRcVB2L00atdO7
IS2yzMjhPfTId3cQCgSQ/G4bI+HAUKZ8ohjmBmhUZwLOqbfNdy4LHF+FlnHTyZEu
jkhRWH5vUA6t3obLot5y0l/Ml/lupyZBNvCRdNc49Cs3VrHdnz/fJj85iXCqgU0a
ebr1jTPzrsVbjQTNBr0kCNHNu+Tne/ojVcvD1VrljDMCN3Ean+ewDYMIB9gevuBO
78PGxVDcEl6nJzxN4FkYTlzJnOkqPqYZz5FvKfjqFlB38N2P2jMcIPAfd4knHlKi
1WErZojKMPRxXIlHQLo9sYBsBM0JwiqOx3qErySkxI0ZWlU4skSJtp0mDUkjy5pL
qVPfAfgwaED4oOgVAvKfrmhiQh04ZQGBk5Z1TGScE/hTiJwRzMjaF/HjZPPBt0XJ
l1ckn8NMbzxrF6NX7uKVSuXsV6tUzqV46YR+m8iKjBY4bXF7phzDbjuli0i4Tmw/
/6UAtutP1N8Py31Ky8wAbD7gxMWVdEHQAJi50/UU0FPr3icLugEPdsJwKj4IxWHY
Vp3orwJVOWcZgO+EaNR6xi0EEa7Nw7OEI1Jlm5MpURL9bZUyt+2qkLjBje9hA66E
ILgs1hrjP77/PmBHVBL6myf7ck4+1FL7ifmh0lMEU4hkg/619WkV9nMm6p0RAGr9
iNECBpJxBnlgJNoLv2PD5KLEghhBNBO0rLP3b5VT44GZ5dtORRa883UDYttWhPD9
HLMUvg6CfOcE5muChLLtp6edVvZUTT8oIkI2K+ylyn4lO16Nq5QLuoCdwtHhiHV1
6KI5tcTcKT0hO/TpzT+nuQHhPWQuAkpG1vH79B2qK0oiqEwmNj9FeGkjFQACfnxI
nV9/iavxfxp3QLXKOtn6DPkjytGkjXzO8h29BOtbGFKpSvDlSi164S3sT93A9v4c
HV2EL/tOeyoNlEfHBKWyrJdsxxqyaxsf6qIyuVDUetXkRdyhwp+e+Hpg7eGAOa+K
F3W9nW0JjRsGpcsCapjtgfRFYiaIoV+e005AD+BlJJ03U4cMmT+VhmRlde/Ko6gq
F1vLqq30bajQaA1fAyw88j92PKWrLsozDmLIwMf/y4tKDS0euPk+Kgm70BzTxHKI
yIWqGymgC0JAWhJe1uvoeeYE4EeKuuq0NQC2oow1CVZQ5jRZc7jOzddjtQxW85Sm
PUjgHKa2ooGN8fYfUJyguHkKV/SARJpcGuD8SN4sDfCXybKR0UmO/RKjA91ewMOs
pdZSS7kpdXsRG8hUBCM7fbuKJqq55ublzhsSzvb4ftf0J+uTumsNx+vgBNTgI4c5
mdYyRehBh6S7mPzF09D4VLpepXbX5CoWKRSqRydLLHOMTvO/1Bmpx2mRqXTLSFkV
0s2x61ieLHM4ItRHHnJp6qlXw1GvMPOURph/Rh1I8CK3nLJ2bVaz31qrHFVSm0SJ
klyOJZWPLLJZqbhqZNg7T4sh+2dFAgUuo65kwBihKXkgMzZ1ihuWVz0yBppNbPiu
UiDaSnAYIqRdwIHeU1QMNYz7HaRIkZw2k2za3lpe/6WeOFwr4ocJOzg/XbBo6TTn
4elt4lmKnnBVjVTNQf+JXeBA3i0U1NBHiWkij8etOSTh8rFuL2qoE727pu/X+K1Z
Y1zQy0AOheLDTfaoO18TXxsIaBxXwUejOPA0YBLHVH+NW4J+1cuEYopzcQA1i0vF
fRAghz/vT6kQYauj2vretKtlRe2HpiC1JSX0XyKO2wD9GviSzJjd6joxVORyS4J0
23DbWhz92VbDvxC8QABrh2u6cUHPhBSggSfUf9N0ACObpwFRPSa9/oF39GKHe+8W
d40K1s/5tFhKNaYy+4ML+J/vRnux6C9WVVyyx9oOU13uaIi/UGAkuMScymKN/lWT
laaC/stzK/3RF1LiGE7qUBbcaPbLwqc060QKOy6wyJdlFyM6/AIKhfH+bf5EiXpq
4BRrEENpIuQADg4j1iKcEz1Uc7mxBTFdZfILgVi8twAnpbUtTEr13j4N6ihVrJNq
kKSo+Bx7pg/ovHLgKmJ4BUfVXIpQKp9q8YYAg/zz0M5s4Nuebtkp/p+1mIbqnzkK
CZO9E10hP7wHc9kEgYXmb84YreNxiY/lGud3dzhipfRY1RKh9yEvL/AtzD7kgYvk
X9Y/qWWY937Nr/tm+zkubZZEqhUrsQwjegv1WxKMs5jMSvh8FD8tgxIwDhcnXOVI
P/VtS4xVCk8GKJSUdpf+iyzWhLBSUiUbl5iLD52uuwanxmtnPf3dIyKkqA/OI5DJ
LJMPSFkGB4TPnCTFuabMAJbfxIk+MkHKYCmX7b+HXcF7gvTCYxZc/xEHRXOYZQVU
vYWzzNGaI9LUJ6O5iyKRxnULbzyGYdgvpIxANM88zOYjp54R8j6wEXZixbqqm9XE
b8mCtC6DDE/GmQ5iAhSLSvSbHukGZ6g2tREhjcZEqKRS60rwVsEdHqbSttXw1iFh
j14Kj6BMKzgr9xJxa+zLPwnLmAKstenhDP3H2vN+fe/LENgYa0DOPHV5XQ26ZAh2
XQzKYjJFH+atgXkcoRij0MExyvxJy5J+/rjfYWvL659qMER5SteZlfYNMJPIErKL
pp7pZUVX1Vt6zGXxOJUWCf4bBLfrkgeDk/RAUyxoos8oerCyjTRULpdHwDFn3QyK
GpwjmeUkyRNXbyzcMlGY/IaEkm5vzz+fcILSQO0ey5M4irPeBe6tFWghiKItlGij
SLvWzo4W50fNRWBupBISPmpJ0T4vpv/VYUE6Od/keiDLbqkYy0w2soEFSl0Z7eWF
rmR55fdaWEZ78zePEPyFS6MnvO2273WkgaOgLqiSj5kJlvnrmnlxaOuBr4PEQE7F
9bXCJGVxvMPOfqcw/Qv6xUH8YKmQhb0du8zLsf5JSlXWJlNTZKvmBGj3Q8Rv1GL3
J7CH9r4Amu9Hn6Nchdk+sNtjiEIAj6s2+WBml1JXrsF5X+iiKZ7XXhuD32lgTP/X
PgkGmw0FeLNfA+u8gHEufLR/mgFKIsj5VGeTJ85+9lAgnj0NhGxv13EgA8iYROyZ
FyRh0hZnVRTJX3h2NBBFT7CF7SzdEhtAdVi8uvxxaVpESwXaB/EM1ocWUccwkfPg
V33yr2GfsAP9WOeiOTBGGGGcSZHeFKHdHBTDR+5bl0Mv7zNtvAinpNBdY8pzx2hm
yYWls3J4Lx2JGlLpl8FpvF9CFaXO9va2itlupmX2BFbAeP3eibq8V8hX9HMGC0zt
bBpMMVybTwlAEUmOycUEnK+7DH7KAhiCohFU+85reOM+IWXAsgbhb5VtAjevh7hQ
v6HSwN7NDPWSJPHtAOLZC4SYSTdk9w3tdNk5g6wcivTbNHcF3mCvy6f3v7Gemg/V
pFRGW8i+TpgA5VNkfuFIsYCT5CbMxIY8mijcBIIueWRC5QXYT9r3MNdzcEbtauyO
BcfgN6VKa0qLEoFY38nz4SlKA6FHxhJ4zt/a2BNQPihOd1MF19rDcnqFmwjoRLCS
rcuIW/fFLrjoe7Di0ZBtmMAG/B1JF1Dzn/433mo+FVMaLx2wwELcQlsYuH6wHG0l
Lyzs0e7QOr4ICpaL4w2tJkw8qXuz52bgfED1NwJKqX+TEg8ipmJHnBU85VNFtZ7a
AJ8APNB0UgN66JzKwy3rWyU3IylWsCOEZ74HyeFyErcuZJjRllvSPY+KoQSLjQBw
t7x+lngOEq+fe7a9fWYFUfOSz9Uqr+0xdXPENRKE/S2lorb9+TqtQvSouiFgeOn0
KeVrpuZ8ytIFnI7LossO1Y18pfv6gzLgAjlh0603+7g7XWnVicDeVLLd1JcBiTsM
CsrVVZdwxzkY3Ko6WPSVna0ZLmpwVPc5riXVITPDu+/C9HfFr4mQmTmucHCUKja2
muWmfyv7HMJcllDsEn1bgGxD5YNlx39K7PJOlPfMUSvlE47oFAatxp7uCZ+lsDqD
nROcxE9qHRLhybj+OddrZqW4Q/Db0WyjL6AdmQov6Fs5m3SWtuX2O4tdpGF71U5G
lgin5UKdg+M+VqWzhPYT8DmEJs/4hCq6xKMUEFwQ5UoAeaC6URYVsrf9QMQrH/DF
nSb08B0f7vlL2jtsDs7Wt1EjAHRpK7Uk9yXUNmTkE8FWEkyESAIfyVsEIBlP1Ef9
oXG6DF6YToG3HEAJ86lriyCiQvFfX9xk2fhUgeGrak+OsFeAETtQFkoHCcfIFPMN
JD8rnFnIWSoyVBD+PzDnNJ5lNoUgNKiYPDfsCXWkYYdX0WplcdgIRdJT4+nTf4v9
mHNHCDsfbQyqqFSSN5xeuAYj5JUdkrGK8WdzkUKvaaXug7z73O8AS/k/71ePUW1J
xwnCrz1XPQvasYcXLlL9IItHslDzJlX0PfKAYR0eF4cMYUYcqGPWBIvpuTA/aAAb
J2pgiwWBCTho561ck3PMPLB/q/B1VJnaEbzr7YshfoWX/vcpqNc3oOuhAB7703ei
a81DjjZZhILO0Sz6+OiKUJdnjH1Ltm7jJQ7vjSenh/qMX6XBJE5DX+kgIl8PdRUr
m4Z0kgZJwG1Ijn2zE7mA7lnB7l6xHXZFqGx4L/wX6xDykbLh8YkaEd7wmdtmSFZt
88Q/zhPNOE7nBj2dY5M6908NXiEFwPCKEbvrw97bZoo87C9Ji8dsf9mw4C7HP3vA
SZhMIU2vZNXks9199uePtv86Sd7OQ8TNQgzvNpd3MtrFXcyB+BJdLlB8iuxwCjFy
urC4APjdWUKPKiBW7zDoNYwxSlG6XGdJuE0toaf6TP0hUxL0f1aLjV8XKVLGcEOa
L1WsccegBs13sMUNtvQa+4U76r0BtITA2rc3UG53ixDTPmQygwQA4fN56ECD/2Y7
33Qg+Rskv0ib+ICCtDimDNoQTnyJbKFBi/W6uSbaxQU49SKLp61GaH7T45zbAX0E
qTAsJinXU08yJO/fUGl+7vMKZZeJS/FUKn1LTHW74KAsfo8CZQev31YoHo2+1Lio
DikDgmbFFuRNINAfOuGBkc3s+wW7Y62+xVuNALdLa4AcD8Zorf/gLi1w/2mZqUIN
TVMFdRODvFLKHQfv8dtJhB4hYqWGZRtnlOtfjaEwaenG1hf42SXRwBNX0wxpOblG
TKhCxkCijZcBea+Ev6dJ2Q7TQlQQ4Np07fgxDyHxt4cTnZReTgdIvJbKQBYEZcBJ
jpJ1HM227+4lghllT0imdmvhAL/dFeZZjJlghtClHGyXHO8yod8Gm5+693KNYH6S
Tq15QasWwMLvAUjUtq6aTnfKnwPo/qAfyeHB1MZz1g6dAdGa1iXfpmXg7D86eAuK
LsC7QNFs7xwtJpsp/J5AycHz15YFqLmT8Kbkf6ibFRffsG40vYsjLGU0Zbd/hXs5
YHS9lhd49YV7Qr6bqFju8O+SzNhjOB7cV+7JcqKYA0eLsWEXVOVfBMSqXBZvXjBm
fPjHmmkUqmxUGec9+/9XURu4CibDYUmmI5X5U8Lz5YJGGII8Y8hH+/O205aIDkCY
iFgnJbb6flUx7YAFiPBG6dqlTnhe1R38GMxGF2lVHOlF7+N6fsptN078xWLWkJJf
AZmp9P0A5NsruOtP3HY2GK+z4qDp/OoyNPjdmJvuRTGh1LbHRplj0wxa831xUlRC
3JJmmCRLgDsKrY+MpTrqcWFe0eTqXIvObbGQvpIkrjpzuP/RCpxKgb2GOhjdPYKH
ocUTOCubx1j3i0qB9/0YzkpFjt9/CoZl0tCDR5UYuA3u+7ifbhM3gzJDt2Vh3GoE
XNkM+yQIJR1nKVQa+MOpQAf/cyabVRvZMqiL7vPfvUXIiOBXKpT9MDoEu5Z7lF1i
qPt/jyokbOnGSQcg/rkmq7hopy4PhqdEkf9Jq0Wh7aBrYSccQhCEwCh8qiYfbYec
fe4JM8VWgmI9CsKtXs+iMLT9FNWly0Y3+5gdq+d3H1YAjDCWpWgZZewJVe8uGST/
of9dl503Dm9Jb3PUW30p1MvpntDqyCAt9aNni9ZKmn8dfnJYr9slzP3Drje37mGF
obO7KUQgasycJ60uTkC0R+2jhPM4wMWdnwsWuLSntnO0xnMdbzLacgvxzKTCEZg8
L2zreeOAdv0bMAmtvFjdH8dZwDK5gSCN88N13P2dZVbx90QLt7GgHjh7cgxnVSm8
58fjI79zMm2ng2tGBjHKqLYcVYP0fDZis/82p61IuR/OuRCFaR0wpUlVnNwChDPS
v4xViQTo8UlfvB1bluUbhaqeLhFeaxVfc44Aurhvsb9LSz/XJ0Oto/OjlpGywmiU
PYRtaUpUEX1dVaI6C7OBw1T4lee+mOIumoPFhr7zZQ35dM7WHCBf1BFIWfviM0HA
SynjMMvuFOIsC+N/aDxyQGPWNZZb0xZG16Qh/MonWP+W3T1Bff9oeHhDvLwR3ipv
ZStZsvWO9VAw3S5aYshmXA0T+ZEoiJow4qM2QmJYzvSqWLz5/w1V5h3jniC0vgEa
Dq2LfY8SJlLXU+67jEx5zENOOGe1L2JdATVPYH4vUlkWGtdhrzHsAiVcbwJUFiHR
IBdgi2xneYJ8ram/21Ihu/gUOhD7Kcgw7SKoIpSzn48XnTL8yR3Rhc/zMq8CKEjR
mh+S1YdhexrqB5glEkRqD7nHxelk9enigmlxDcEbK6GW0ilhvp78xLlVu+JewPdD
O4a0o1ggdInf35b32dO5GEc6QopgblH5HwY1fdZGb3K9QvnxSZ/ufR/oxmpdWH0/
4AYiSkL3Z0pG5G3NA8vnpTkgSZycahy7OHDKYSUQGkScsfjIFjAckdYaCigphrSj
OgxnbLcZ5IkKxFkuJ8O4sIR52tGnq22T6nwk+zRFyUczeA9TR8tXNtVCI8HUjc/P
IJI49mYuFFrIehvgHzlcjZ46bEXqZT26VS503GqkhL3jb85JIaDdJ8GLbcUYB4bF
nquG2rGVQlzZ5Gy7T3/pEebBxXBduQf5mxI8f2NZDfK3hH4ylGThXjsxVsHwJCC3
YqYX1UbsipUfSvK+B0uFP5EG23B+2SpzoATYT1ROrzkzd+P5gL6oQQJawHzNFRoq
KFRBdl69wqEc/nFBQ9TdldEbvPYCwM9K8EMWW4EQAZKCqoxjeKaui3U9UqxnZ8vS
cck1MCP0D+/AE/ww9vKBkd4T5VmQuKzmA1LtTJJznuFtIjr7+luIN5NN1K78Mpo9
9qoft7h++dbcHt4LOVP5l0vR8mjPRcFvDjT/1IAy8yJVAgFbABn00LjT7mEn8L3U
DFVfAPv/L4BVvn17vOwXhTY/GaA6k4gcg8MYQZPNc5NCCc75ApE5ASBWvzt4FKu0
y5ZbGXomlEX+GmLALCUmpC+4cOHFJ6t0220Joc+uYdUOtC34tCfN/eveBUL4ver6
GaPgVQPjKPUXENvaL+KhbLRULNuhrORQiIEsPm2hMmZ6dLqzw7kJzL0NWP9jCat2
mPfysat4iaS3bEfLsCmYsSEXkUEV2A0fR7+HcZpiSyvY7835T4N44rjb87wGzY0R
5l3CdVx9zlaroLPqQD8czLnfLJEh9rhYHMFqUD5LXwDtRGenEtSEanlVQbA36n+W
9n23BnCtYzrhsE5OGRH7nUeSr5egdgDX7p8WBy/Xuv6y/lFeBqS7PH1QcjAnChxS
mAzQtPlPOi+Ugksb7zG9TKrB4Ez25DDm5pJkteAHuFxxBZ7ouoQ6C+3XF3I5ixSi
wSzIKWgTICaVZ6BjsXQ8GhdUj2lMB+jLyiA4/FyVSkYj9MawbBL+XU2cSAle0ycg
KLY75dxOE18A3+3R7ugq8HK1HeuD7yPKq3DzwDdBuVCG3oloNwvqzUxp7aXJNMvv
DY2TjiUTPJtSOzASYE4W81QksooPhAUwmHwa3ZI6I8eKmMQKkioQtFoEHgy1vTx4
T+5BTnieMJxEwG+mgbbzv8nExAxla4269EaomqXwh9qHOwKtdTHC/RF1rSZECdWF
mkghXWNRRIakM41JSRqj9CDuDXXhw5g4y7rejRfG1/bTnLzxqr/2HUjm8/4/EYXm
nLM0uk+ub9Bc7KVg2+HSCL/JBN1VawQPgQtGet0nYSXs4qt+nCSUW2W60p5/P3+s
rNkBNvJ0i9/40U5pe7gTfe9v0t63nDXTglfGf1KRPkJlKvPBME7Dd2+0ePM6/asK
a28O7vRml/ugJZLFvFcuqaDhPsmM1ACl7Hpp74zVjBLLkZuxsV4PeCMk6H0hPt78
UvjE7sAJIaemEWAHYZ5huSdJzC68oIEYOJyKjPiO9iN75tPnNrntu0efikEWcd/w
7r4JxUedKRyzbDBEKznPtEek4qylxJUu80Xe7KpDzIUzjlQILFC1XumLLPJ3j8KB
jv4BIwB6S9O6sSmcEKVqoEMtHAqzMjaz3Mh8vvtFo7nhmIThkXdtJLAf1VImFIXL
IJGUmtAFsAQZiii/w5ANSAtql7lYNYJ3PiLmDKyq5+V7lisrR/dBoIr4jtOnfIXQ
V4kpvGbvWveldI0WOYl82CnK1beOQAonWfmNAvH+ruWH+daBBrfUvKtLv+8to6rM
3YxbwXRRcLozvWUz4is6eL5YOyuaSwwcnoQxuzLUg6v12Z/Cw/EzJC/wk3O0WsnZ
fcw8+KvinAvlZ5Kelh0uL74qw/wkgbx5ydxZNfqADRw3pMH1qTBveNFgGJZN3Tgv
mXiBFupZbeR9fCelLdmhGVyntvH4PxH6H3rYOEmbrsLy21oK0giO9+WYww2V/gA8
B9UiI4dNYpE3tCpcVmo1NSkhijvM82NUhUx2SSTYLtQ67Y/5uBDcDksDhllJ/Z59
5+V66DMzymFB+fO6GPvY5hDeFXD1PWU/r4ypDF0ilGdWe1hrtnOxnvak4/frEU+J
IcdEUVurjsh5Ybv8n9enCDJW5gC0+aRBHW39CVf121HsoowdpqQSb7x48M0ucJtZ
jkf2WEZYRbFImDVg/pdJ8K5NEEMdi6oB+KkFalsdjk9/Fo0IUinyYYFIvVWrGX34
YNsUlKxn2+1zrP9kyKxYk7MpqX8I4ee8uNyEZqYS8D7PtyDeXgzFBKJNjt5DXhnu
i8Wmpf1i8UoSHmCa5xqDjUIhtbLhNH/jd4W/H9IfyCB9hKAiM5LsjdiWJRaIj0dg
OEw5qvXknSEJSwIzq4Ea7Mt6gbTZmpuwf3MLvaQN7Dds0CJeD4fMnA8/v6svrmYH
87EBvEjytl+hONLtBdNZmLrcM1RmGxg8G21z1cR1Y3OmUx+krOCWky9JOWs3iMgS
EEbKymQeJKbqFwv7llOpY/7CusfB44NxkCoAHHY9MycnmsJAnq26c/HhObIbPgE7
OqnH3LYKxKrsRGBjFRUGsSlY82BVJQRMXKnd1Ljsu/OmMeRboDEJV+AQRj+gOyag
f3gzJ2Ep6zlQ9TDFM1mGA9Ac8XQCxnr3xBZ6q8Qp5KaAGuhnDfkHKm6CelsD+zsy
awrzz7hfKVX0J4Z4wUuEeNQcPXzRJ4nXUIrNpXiCHGkRa8JRjiy0zqMaYDb+dil5
FZoX2T1Z8sypyyEPJHMWO4q4f0N6r23xrPqfPDWZNihz6+ZEa5Zn9k+yquEc/AK3
SOe6DpKfPMLcO3RGpK6KF8eWj30jGYepVr9lFOLzJTz/gx20crfYiWQkTPbGj7h4
3URp3Z524bROoHwkp3+s/QPVNHnOFt7NNVUTRHjW3cliW68F2qRxPlEEyqLyE1Mf
63XmZkeJyipyIyDFFq96Eu3ypjc/jrfSJq/pKyZFdBWXA0MOJoknaeSuZc2y8Pd5
58MYJIloPeOHcnDrI5cM7+dIl2BavlAceCe+0USpdaan3l7xXOAlgMaDV7xo4NJf
BpoD4ehRfAVNE7TZ2zHBpsWJuX25yePNcG1Vaxv0OjHCYueJP8g5mXimLuAsNEhY
twvTfHPfV6w3Jm9gH8kKznC3TfcCySxG/qzR8moUnvRBEgB6q+vyu2OZNsnPs4yB
lSc54r7wwNBlWqlCijC8g6mtmSTTNqFh8FUX4/lspAsxmdcHUj9njZn15mYp40Ev
i6LMmo8RMaofS5Q9Uo4xkyQkRL5faR8W3Oo7xEvcEoDhOhxBKxsUy9s+528COwL0
JOGWQ7bmz3Gaa1wotgnI0Ehn1IR5PzOa40U7at12a2cnBY9OjDgz21kU0hra74yk
BLWwB9iqF1qro9NkntXmjmzIlwN5+R1YIbHjtqBoBR6FaS3elxu0RD+lr6dpNZ1i
UXCKnfJt8AyxoJPcnreHATDFt9Patvv0s5SquvqCNwprP687VhVqhhMF4hnr/aCl
aRrmJ0mclWZKpZDTbPyoKSTbehTpbu4vE+8l46KBbJGFK6DOPvilwTLK4fUmbLjc
aYtZ0mwA1mehNatQVI/kj9JKFPVrvhSLnXT3wqMGNkPMwTaLrk32aqroaP6dMsHu
sF84Q2aTIkFwTuQ5Cgw+rwNwy91Jmz6wfvlGr0tJSrsSFHAXIssO8HMhfQlxKKCB
jOamzkTd/fdHZU3IjZy3d31qTUpW5BurPL46MtIWvW2zn57fhUdOUFVRlj2uYoOp
OBwL7I4nydGiQc3HuXw4+Uvtqkaph6qINmZkkaXrzbrdSVhFOr8Ap1+glnQfr3+B
lQ8vupMTJ6P9BQgfhkQY6mPrg/IbW5UQmCDgJ2rxI1XEY/3A9thUAXxVEkypNflZ
blrN617/Va3vXUV/Omb7RMGp5oXnKBUOJMcB5Av3VR1uYO3GWKszjmxaqI+d55h5
uoVspJOeoHf6r1g8UM3zT7AAiyAaLF/Yqm/Uhn7XUyegXMxA6ZhPhnA9qpHWmbL9
PNFRJz/NviPX9NkaGnSj/a6Sop4EG+O1s0w/VTuMqtMkJ+Xfq6uw9s3WTl1FJMuD
fmZuYb8E3pc3+Ttgv2af/0j80hQ4TByn3aor8naBYmQetkA3hdjE3L+nzjyE7XV/
r0Lu4j0ulJ3a9ADaj8svspUuEvyTgRciE8lxZwjvT2jVsQXA5c6yAFa0x2vd1qbp
2q+AiL+iDLRD6a6U1H09WYdmBdwdcITqwLKcynfS7fe/MA3Q11uaoyl9rbN7w5uw
fUVuDVG4SKqj3XagPs68IYjuSqaxOYKIttg1xtmImL+AXLH/V9SWC8/tAGrJOw9s
9fJUVAZ33+d9KAgY7mbw2FABGARt8LQYKnQqLKaJzYat67gC9ac8OgTzQD3ts1mJ
OTBWnHw/cF3KbseV6iakVpzKd9t0s3iqftBYHoZ8OgdHcITU2oVz4c5PFAfEnra9
ZLfJe0nk4xQBNGpmIzclRnCJqEIrn7l94KlIeY6RwEcsOpcEuLPTEc/mNIxxkGF5
OUJId903RV1rzoy1PsYy8rVqugB550ozVCzjVxqdLafKMDdF3K5o/BrSl072plyb
hfYll7X22wrYDWjj09B68rMENMbOVOvg8vb74bU9gwmiK4h8KT+hn2IKxQXKBRUV
pkid70AmjIkI03rE910aJ1g/OqZDFsuvieiWQHUmeH95PDvVWjbyuXrfVuPOfvs5
wsVilML1lIqVzySe3OVxyk0OVyQ9WL+ZEVnLBVooGDSkUvIS8NXpxDdazn2txIYk
CfTwAziKNnikEf75JmpCUUIXMJ/bSwjCpuDP3R+/QriFZlorhRO/RfqSLteDStX4
+Jii2uurCIod/rMbls8Pre+gJ6fTJBs7MUD56S4BSH4+JZP7l35fLSrcvhqMtYP0
dwx5XGog/lbyj9b9ZmFgU3VhJW4j+GyxxAWrHQouJ+Swm5K13l0vVjYpuDJC2Eli
x7pnBcR4+myt81L/xiJEnU3qVISUG/nbXYDJu1nMCUlD8efOeWre/4yxaZKUMs+8
xaR8ZX2T5US+wpe2YDlY4Sj1pf5cAR8+q8jNVpnxBuHc3lGPWoXzKIg1xKxgBHWZ
z4v4zy5OFXvceEdmWAvAyth/C7xdOScIn1dsLKd1GdMlX2iJb8zS6LF7yYCvONKv
Cr/mJW7m2bilx25tDFBBr4IMhWQUSJ5bHojMvRTKxNBhQLJ9hRz0DQmz/rb8jL55
OyiEeB9s6JbBMZQvNNTAXzg04z1SCMpYzc8s8nykdNv4O0shC1Grn+BkF7sueG2o
utiENU/OjALvcpDcspZWPf5wOEidwnKVHGynazL4vgXOoT6CMM0c/9jGNdiIfcG8
ZOdXizS9RS2FKtR9gBI3olK4C1z5uWK1oXdIt+aH+xumSxX8QxT7YywxJAm37FlO
WsJaomtxBqRBAmCAV2vw+592YsjsMWxS7/K49fASTbkT0Gc5pykc+QXaKviMIc79
htbzxcXBU3JyaWsJhNm07cYgFl1PbbW8WXN1zO+OsRCxb3vfwPvZMTzVLtBjVuJo
AYsXCDnGZvsQvf7o8OcWH9O0+y7dngrRP7NBv5rRKkTPcoQZxIJlAtuknqJHk7WZ
8ICtsDMyr9H0jjXA67i9vBEn1HcHajH00EF6/0AOxApcLj8brqXzXDOC3jUcvQP6
ZlHbJtkSq5fbpUK33wIbD+rVeReMFj99xkE4280hvUhEBCL/ovUHJtORJmb+kc/c
f3+1Z0tsyaz6fZzwYqB5Ao+pxWhCYDey9KB9Aancfla3iYUvbjAxjcw9rrHPdPY4
QEI3NbNQGv8MOWXiGArV32V9cKs/rDOEbBOZGfzWmwPOpV1a1nn0oFvLanitpzfA
iqoCUMxpj7aI//YIeVKZ9fVpz66BZPuDc1iiTotHHs+NcSynbLmmF9C0pNfVr9Ql
nNoUG/cPA34rDyHH8eFD7Zp2Oohq9Z9Dc//U12O6YMuHjHkZ+4PSIqQrb8I+EP0w
1eEHgf0NYSBuIsNq+0iREeooTvQisCy/w5Z6TzauqSaIxJct3smct5d5BuH9/Afm
uA8ti5kI4ASoPvNHr2Shtuf/aurSr4dW2WhOE7clXiUv5lCXXKKZRSnHF14dhkzS
IlBt06zBAS9P2CSFFgOF/S37UnItj/MWhyYCEDgdeqtB5CtVashncgpTtQNKoKKw
utYZoCYrbUSKjN/w9MJEKqgaFU4VhymvCm6+rNkK0Vh3PJ2qf2wDSgDvgOgYU2rd
W8ctXH0sdn99oBXskspk7Tf+82jZ7L5y0ql4HcnEk4J91Rejg1Nxpwm/kyFv4nG7
9lBzm+NDRdyZvWFfDRoNpRoihq/JCy+JzfZYVUrfsRC/tZuLYoR1O60tmiX6an6U
7SRxZM0N6ch47n5Ea/i8PCIIai7pSqfvqFBIP/i+BDOg15C2UUPviKKgIFeJ14f5
eyQWOhPqFcxzAeI82LO+UHna6OPZYhUHkpuL9DQE5xEVq1ivz+b5qJ/4XOWykBfM
Rjwj9gw+z22Y2LGxVfaM5ulYNy4rB2HPZflK1YGJLjhDLwAnW9a8wZaM/2ECyb6J
VktvvE1UwPLFGZGu0Nt5oZtpRTXjHtW0rcrr2oAQdksCqOFAD1cB+k72rqQpB58K
7DrEm5xl9vXPSOFvwmskjv9bbetwm3o6XB2Ze6kG+A7nZUWZV28LBhO+w0p2nvDM
aoWZ7UfUgkU//4tgoCNEDoZrPykjo1mXhzHcVJ05w3ae1tZhRFpa5XuhfAE0aALF
0fjEAOjfWqwrsID7sQTAPET6pRm13vBFkfSUU7rZuLKC6RJP54Uib4CY0cW/P77A
Rl62N1aXILrLdBuBM9UOrEHKtOmiDPkaFOK6S+6xsJEkgHz8/u58DkPaiCtj36w5
dXgECpw7xMmzJg4poXujCbqqRgM42nERBLN67pkNtqvbwzKHzysLXLeAdDeprpWQ
2S2QAu+C/EiMKrO260ulZGoCT+TMSX7gGsNCMgUVmkY0ifmluLSzDeZcmofhNnLj
HLfchbKp1XEvF84qwlwjI1T0425pdhh61eJB1BjiBT0/TtO26TbJnFe7fGgF6R55
d99MdjKLfuOGPiIzvPWjHiTXDYiBP3+frYej4QpD0n106/4QdtweoZ1M69jJu8WH
qelYDmpiwPa379BCX1JlArBCXn57EA5zVUJuT0yVNJ9vIOMJMXWuzJNeltdBH+2N
iX1myyhhO1OEe7Rl6/rqScMs7kdzj/eOgxpvtLWlxq7frcNb0oiQZ5uFmy6JBYMF
cVyofj70qDaAsjXUfJCNm0UbZdU+8FopouF7GTPZb4T0HEeQlfVSjV3g33qYBiSd
sRtHp1/fV8mGa5uk0ui1N1O6hmPAU28T5YMHF28OdZw4OnB1MGH5P9CONoJkcOi8
RGiz/5wT5NR+PwYrY7hD0CtYHUC9yLSFonyUoe3sqTnQ9E17cDwShdLLOoLOhHgf
euIbCPu41s+6+jdN8M1xEr5Dz8htSYfZQZ5y18jXOjmxisukmWLpw0kXvfSXMnCE
qi8RJ3L5YRJX8GQJmkT2FZ4NCsah3Y5AMPjjtHIdY8cmUNGUARm53d/CRXGP/dSX
8pCLZ2/EoR8Y9eMZtD8aPghMUUlQFDTil4qjOeolcpfaloWSjfc0PFGSjaLGidlE
Aqx9Wnoo4hd4qdvhq8Nv7amX0PTBozs3Li/ap9JGLdgwSw82pS1uE5X/a0slUP/P
ntXhgdPLjT8+BTR2omLLccdpHlI0i/GiQt3zU1FrVYJgttmvjd4gUPjO/jXYM+mR
OgPkpVZ+XfGgRoSKr1nRdc8pJWR7YD2ovWcy9Ts3F6MhXdiCI5n4ziHeOs1KO2Da
0bUbQe6XXazOfW+5BWjWgBEk0SXZxyxaJ2eOLHCsCcAUA263DilyuEAx++hVb27s
ApOtxpEBR0LQ40BsDWNf8wjvz3spkF3+N155rosEFa+BkTixLduzpO3H5cdmINe6
kpL5f7eFWTmfVkTzDcTDdSYoapyg2Q+65lBccpljiCoMgY2kpyedmv+Ib8kMNQRK
EGhS39iJJN7lT7G5GFVJsYMwEgHbbD442YX4riLDwV6wgMDVaO7RNBhuwyhDFta8
XcssMPiEkr427ZIFiRmmNYCu5tRiPKt0XhKJCYbuVg6pSEg1Pnr0lrOZUcV0o6Sh
yC7m41BZIQulQZZlEROTvIx6nmCb2BYmw+TqDhwPzYUH/r22XZauF02Op8ONsnrf
ySG4RzInU+yV4qxFfXRnBOBQ+uCc3qX07rtTzGRl/XqWmTA6U8sXwee/ulNElwBl
S7uHnJ4mwWY60hXoHDJHCpYXAENJkaqk99ks5cg+BguU+mVKCRgEMz2lNx8iOILD
/KJpc8aODv2c32E0RvtxzbclrUOkOvPKuUr3GTQVRXUTTNI6/ER+GLupeQ5Y/3mn
xo3X5eY5RtJlgqh9UFTqnwKsgI8Oz0mX5aayMxjsMHuiH36lWCvf/bcJifd+20zI
DUlsE9PMPZzd5kmcNu+OuuIp/3c3ActB0RQovefMhXM6wGdY5cNsQxfaF8DKZlg4
1E7V/WwrInmayC9aEyHQrKemF30TZorxYnrTv4bD6Wrvziv56yTqWooqpLIbZd1m
K0Qyvhj5RF35vKKMpkJ2COUvn2UUbXR2z+gy1Ob99oxqXVcHlD0zCf32Wv/RPvZe
XyrkUIgqKhnLJPKuQ7YMlnY4b4BN+NJmNCreb6pNpRZg0uIwrW/Uf8fYUVpx8/6R
ifE0AG8jAriRwp+PcOwqA1jR2VyUd2xq6p5dzS58aB6o4vuMPBddAGhCMK3FVdqP
8LgwInWPFJH9AMY20btmljMqJmHgChix/Xjzjhce8LcheQWrWaNID3ROJKaPxPjS
Xx/kYCGa5G6fo2/bEletdD8vwAROuNPgDdYrBikJfXkm1to7CFSi+4TAC5J9qkPF
jjFS7OqHSLPJgJZ9Kzi50cNwwGUFMfnDp8QjNzJY133PiOBob+uEQ4rhBI8SA8ck
NoIKWK4rbx9MEpp9xGVoiObFwpk7Umnv4Ek0CWMlTT21kD6B0fuhawoFemv738NS
2+gPTfY+rkD8GDM0gk3Z/a+0Y0P5PN2Ijqr0hn8lyFgQ9mva0dU8Y9EZRvih1MAH
OQyfc4TLUMyPcZb957WU+6Z36u/CgqiwSzceV2TYXm0MG6G+K03s0ffJqnYjXY0U
MyUznZiGkEiWhw/QCCM3SMx7BnkqWHA4nt/o14S8GCzIpsqCxmsSKOn6BQXxtpiV
IjJJ2O3AyDjYNr98JaNnqw6P2/ShYt6ba9+nKH2j62UlGG/iRg8V5rkOcyxrmune
fjv0ArF23+6i5aSKpq4xWcxSbGfavKHC/4fKxnqIzuG44vsfcD2tisJezPdloOGL
agiKf7dLi2Z8TgcALPL8B90CQ0IjoGC7WxPtB91tPhsuJ2POZIgNkVXa4L9BN8Ep
WHjTh8OENR8+fN8y8Z2tdi1v55qcP/NSwlK6yNdYMDYtHSZAyHlMbEjBr+ZibjbZ
3MaV62t9c3nDQCM1m3Pt0jUQouIB924ucd0T69oH3RbHOAoCvF5L1CxgWB5pxCU3
MChyHjGe0QX6M0oXdnpTiFBbOiTPR4S//p5ufE9eRT7U0UIJs7x32/fX0ourYimD
6peoMMqHoCrRhb0x+QhV+1Nio+uG4jMDt0D7Rj+1eaDQCnmbWgI8zBXu8vnxUcUl
MnwMuBIVWeCnO/P5yA9nXv3HhFfJhkjf+VuQldk2PL67mm+TyNx8SCDUvO1GDqGD
XklpWVIC127lOdOIKsz4YBFsWJsHUId0EwVDc0EPc6VglScjllZmX3m7kRtwmoBN
MO/p2kunnW2O+DnSxNuYnN3OUAmnTOQdmM6vs9mDQlX+4eX7PKw4PmERAVHWeU6l
tXgGTkH2GxjE1FbJfZVe2s62zi6R24ia9aZRuRQ5zjWzwythVoOOZB/HtRqPZjTl
MNYrS2mxSOK4pNok2pwkFNXbQ0sn87k3ixRro5RpXIYxUvzPwXNi6il8XI2EIJeI
pjcRjtOjXXnNZr7uRUNSZOZyEquLzLo7PEDaKjrYKns2Yyl0HdH/aG0sXm/Irayj
XeEf8Du1b/Tjw1cjlxIdOgK/jTZCNVJ0HZHOLgCBqs08DpHg+oS1w6Dp9prVlI2m
Yb3GFmMcA/DvVf16iP0k2x0yi7BigMguuQmSuGda4rPCXmWp6h+siZauJomhL048
Ehesf196tsotGGUDDW+G02BTfcLZJubIfoTsEt3EsowB60mFtyTlkxyiK7RXqa6r
h2VYNRpBW88+RUvKv4DYkIkvj9FsFfh009DkwdxjL1NsP92jbXEIHBquJpxH6eN0
vYHVjhlLr5ftM0C/Mcd+D6H4dapTwwXAEx9W24n8NpZNBthQTriHdtb+HEPwGZKD
3OqonKJed3Unmu0AoY6mx4JS0uGZL2P1mQJw61UPlCFNDD3TVqoacuyEfxaODNxD
r1uFoGhNf/kkx1qhankXSAyiquWSWUT7excHn5OU7PW7H1SAWwPP8E4/iJ1DnDUL
H7MmOO2B+UL+9evSlx/YTuZoxrIVv+lcBSaKdiZpDw4wT5LOs/AxZuVrBLJONFyd
DNJrtSaSBWmfriRWpZ7pf1wMb6Jsk6AjZpYjDV09sLNnMlU2Vackpe6Uzo6uBZLM
hhZmBnGg7+dyZdGRVGSvqAkExtEYrJesPp8nZotJ87k8Ycu62gnfq94aeg6tP0bE
xHlzWCdQBYSZ9pynT7caj7XHXcMRUEvjOpWF06wE+ZdMVjw9SPJPbKdoslOiu/Yx
UDwXiEkXBXD8SHYE3s8VAwinbr9VXGJ8u9okuTTxY0sXfbP2cpWDCchRG9OR/BHO
jaXkH3qCR7LWrdonGkDUSdoaA4jUUprculfR9rylLBbmrTl4tauKvoqxAF2+aKcr
0p2+0xeCLSk1EvCLzKezecaMUovr4bqU8g5V+rdvDtNOd4Fs0rJTG3KyMTqKSCm0
US0H/WO47VdA5XBNgMY9+gaFC/BOVbprDtTsDcRQsDDz6c/PrBscMCh4xb7gkA/L
6YHpDnBuItU4tlNN543WcccbsyAGanX7f/E8oqAwYEgoWTXGw2R9+buSXtcERiqy
RoBJ+8S2qu0NLfdP6hlh6ExedAIcZIofdqM17iPhKChtiXIdbIifMPODnBGJDo0W
YRMVusOVY379eQsRD7U3YgoY8Z86ydasDhaRWq8N6v2CXsY50zN4WkZVjYvpqRXM
TV6kox5qmbVUzNg2b7oIEqg28KPEuY68kn/PE7acJ+X6MPc+msStoc2/ZhJpiTau
XfAL22DMFhweZCQl0UYPrnpi780N+sV3rYwNrdjbbv1TI5EUHAgWRpcU/hxaaazy
p5ffY32V91UDIM3lixfpw65vDS0Ydun/6desD1xsltY/N9FLfRo1SzDZNGrexnUa
etfbzCCib5ajxam9JWpg60uIHnhX5Rdw85yP61Ln4i1GfbCs0hO1owDIGIQgpakS
MOvqzCHnGnAw2X4DlY+x9HnwaXaE/hgGCuDUT4YmiaORQRcWlmIJKtjFEUajqoM7
MBZQV2+wa+E0shGiNok1CDCb6Gtnnao1yngCXZKs7r6ljeWuB5pCGZMn3Rx0s+2B
vw0bMHMTJNkUkvL1RNXtNk6+PejPRiQppRqstp0M5/N0TZb/CAO6MVb35EZL1xVz
MQ7hx8I8nuZVIqS5CmNYITLzgHwICZ+XeCY/+LGz6sTdX2vAFHNqma3HdpI8wUA1
R3RUKHNYXum2ZaCYvnSG76BqSr2FFwVaBS0EGgQ0jx7CPOPDVqY/YE2jmcgTz97Y
SIVIZy2dAVBxjYnQd5iSb9DCQTLlmMUUvLlLgl/bexElFO+pjcSGw5OsdGfNAmGI
MbA6r56G3QeUocr5CifPHVH+VdA4N4eznr7f1vIoXz+NSu5Z04aBwR2wXpVIHqdE
4XoIn0GxDE+uM+JW3+Bk9WaqH10IuNSW2Fb8YIcKE6Qpa3wi21jnsgDFq8HPZNU7
whAY/wfCH5/P6WCHw0AB0T70OwHDSUTZJaLxoZpPd/hVSIUR9/fRW3JYmIY8BaLE
F9w8xUNLDOBaW9Ylia9kPOc7v7eN+JzKC1AsyUodu81KBEGleBKUnCPl2OUepZnZ
0G3aSBoCC6TjZOuFh45o6/1ffRTUvu7G9jWYQYpzX75hNg+IbeeJHmWLrb1t7UBX
8JaO8cZoMVYEzB+QLFX3I7G2jlzIw3mU6G3dKEQkaydrCOkHigCCZmYWxt5uE375
4kqUfib40LYdumTOmgXGeUKOqgxztjmM5ydAbStlH2EmdbOAyo9W28eONpIREx+F
7FrqzGKt7XedSpiZwVrVIPUxq/vYTyTyvB6ynRCVgRVvCoa1vEV5cD5A0U8b8bt0
tTdJ7f3OEqjy5fpxTYNkoqjUH3ERTFSVWRtOb9QtouYn/mUaG12eORyRvdLyEvGI
D13LQp1jbW7OwjUbDnU6MqJOQGm4Kwfb8KlTD6R/utthbvs7jkDsPxS51VXnl+6Q
OxjzyhDTNWgBQXTm+AShG3sqSvGj0bIRxesQurRnlwDgTc4Yyj51lKqciI3B+ilo
t/X1xX+HNWqqL5McOeO+Y6sx+0ehZJPUSVmAiXOrtO4Qemo7PfdMI+w7CsZqyXSM
PNWKxiTD57u6UCCvFMsQzfaY3TDJMKkpVx/1ynyUiWhw+V2Z2Kwllwo8JNtGUqNc
ab0Fi5TgJiODoOub5sJA1fBAFIYU6Agi8s8OW4kuapeuKf6E9hWlc5V4d+CWGmai
cosKjv7CUCh1maeDJa+yyGb93GOMBG8f/oWvsA67yuK9CWIBeCQ9vYyWeOLHAdJJ
eOyEke2YpcJlbRZ88wWEeUCXOYhMvDl7SS52VNyjvL1re6bnOECthZdjOLwgoGu/
NOxZ9OCyLjZ0vqn/1t67AfCx/FDERuee2lJe+6xUWeZfv/Ek6DLwUHP+TANVif/p
t6/PRPeewKz/AiCL3pP0o4DT8j7ZmB7oHuGjFPLKOWltR74m4e0xGNUVWv5lsj6+
0Ehb0HjgFHPze5qkd6PUU8LoYwc3kEI1NhYVU8YMoTeNp6bW52aiSBiSxrUbmtej
dz4lNJBDKIUYAF8zY/ql4qvBi8WySWtpRoBzZjgWmMiGN1WWy5hRjo6UymLsDkVb
CatinB8zdDlhVhNj4eAE7DUkWNrCGtM9xwelCvD+C4bCz4i8wkIiOly4OF6ciRRj
cY+d+cqmEpn5o2RfKTmyKK0AR8BKKUrUv+Z/sDNZhkvzscvIU8OG99yRpvitmZ1u
kO1LLO9DmAHMcaUssDcOxxkwyJQGyYyoTPNtB/SF5hHOuxwCQS3iV0BCMUlD4zJk
8l8MANwer0/pzZkSZ0Gnxkf2vJRmSSVlnZsjKMVsEVDLqQOITb4UVrEMVTdjzbmW
kv23Pf/XabtKyTYp8DY9z15f0KypLaUVWUlv2d7yAImV21YFMFsWzy89ACH9AEVr
ZXiWsNHjbxUo5+A6JnhlDPA8JuTvE54SloarzmjD01zfOPPjsvSyKwaQUyrHr9kZ
pz4z3FZBhYdZI86dH83Bkb3o7FpYPqFeiFIUPnz471FcNJyxDXh2+SQOBUvjvrs4
1OpPdyxen1yxW7HRp7Uaoo8VkCDnSp0hAlkZZ1F4ZaDDiEwYMsDn+1toj/o1DUWz
FEdJHX6fFs0abNrxzmj/RKPqp/m72bglEN14KmiRtCHLzE7OxkHcs8l8LLN1eknq
zs4atk0vuRqxPYTsDMVo00jgZUYmw+4DKSKNQHzpfBj/OWTBlG5BBAZkg672bdGI
fHIoC11oU4z7wyf+CfcRvXxCkyqrdu+uK+Lx/sTRyl5Yh9lSyaWLbGymb3a/ciD8
CBBPlGSgiFRWf+Fd9PsbLqrN/zgCJlslFqikWjo3AYs03YEmfwoWu1DolqMRd4VI
kdoHhZvTwgsvihStcq/M4LYxH8JedxSPql3z0POCBpa2xAEjo+FtzlBuhlBZgT5n
9rxdBPvCgqzXu7qGNvcEfMAEgdfnHmD3YN5+02cgb821fktFRrIGafL5Wu+qw5ys
ZwiAawAulopSI7w/9pdEH7Qi1s6QgIQNG6LWNV1HrqEGbOSX9rU7WjllqGFR8ldn
kT+J3Ot8MaaXZ9FG8L5qwLY7D8QItfbu9OdfQOuQDg1zintpv8Gl4EanJ2WqRedA
r04IaLoux4KdUbgr6C/cRpMvpJPukJE/N7XD6+JvGR0dxwbXqN+jm4fesmEhHirx
q6jOQsRS+pebkB0IAyNq+u3/JCBa8kv8UNVX+/h4hXaOnl/F4oLGFyCHp6XhyDU8
pC2VerKBkp3M32FoNFS7xUcVbfy6sKUfH6Zn9yHo0mtiWi9dzoca2Silsl+m9w2e
Uqm0tUvAaFEBnEXtIlrVQFg0lClpDpm7ZOsI+kS3My9kXRgyrYyph9bcNtQRsH3J
wnUIghuaEpPPZM+4oUH8kVroPp2/XJY2uVYWGlhfqYG7XzD/LKvlJGULWrPcmFvL
gS9SsdrLvOlcLYGNZep7dlzwaSos9x8/XlA+SnAXiVO2mutSd2FbpjyYpePegF+S
da46+qngro2VUqBxB5BcaXpEutlsIx5p8VmsezlC94UMMyBTHSCIdEio2VjzT/VT
43EbsGJuSGOksJ892Inq5RpUQ15tyTaWNvxXoU8yQ0n450Xwe90CNq4M62qVXGyH
ntAxptd/MPH+BaQ4bAW30v5wu0zAOexrhXmrNpXA4Y/hwQLHbYNoHr65Al+W6a5s
TTejSsImgqccizW71lrqwZ4P2CUsbNXrF/VWI9BJWbGAutAG2g6dWP6ABe/QRESM
rP8Xfi9XHNZuzR3UDG049d2vvl8UcyvQHpweMzOraRxHq7gmilrL2ARJHyF9miIz
vA2Im/Uejn9avxNtanr6pRwqNZZOnOLQbjEekNkEm9mPp3DjUC0d2dj/CtxFYecb
CbHPwhTvUea566sBTJCm4n8yTJJLb3JJUU5bx/T0tIutr/b4pJWeNXxArb5FsGVG
LCunnCDkx4lUF1HUSizK69Xm8TuDTZUs6ZclCQ/9cEWBXWahpRkDlJioqI3tn4rE
kmHHBXTnKfLXFYv2VT4L32My+ByPCF/TSl2o/xH82Vo/a6PKclwO9FgYtzo6LCHw
DHmczs9uNM8pg/8DkrGGgvSRZOco1XKeV8ps9WliL69ajIuqob8Ajwl6fmYVszvf
KEClxpoqKeQxJ1Bb/CyU19u9gMqZB+U+7xCG6toDFpgq1pZck/1d2UKvvXHe4hzN
XBpW9ZrrX/cEjVZ++8h4v6GV6HoCNeOir/RMAIqhfqrsE1PDUT9FP/iebyoTdQdg
1lqbI/EZbhoghxEvINXvA8j8DJTg0k3sfVOftuxvaiVA/TFpHRjyeyUH9np9CymO
YwRk1Vg45BtUq17MsMMllI0MyjK9scVKTgG9Lp3D+3AZCbXmX8O21n7wLOWEfRzv
lY5OD8X0us3ScGdHjHbmQ6nhPslWf9jJdeJyrma4UN39fU2COKDQItDMEylOtT4l
GMuzR7MxqsxKlSRi+qPTz0YskfNHl7lfwbrKLaS4LSY//dJl9tj0JtK6v3bgwtYA
B6668qHxHlzPIJnoQM+9L+Gki5zZST0hYQj71IZgAamzpGJ96ItUdW4NcHGa47vF
0tqRl7ITD1rXwi7yswTWWx9/sbMWQ+qsHgELv2DPpmd+gIFNVb3E+5XK9PBVo4u0
59e6E9mKsB6fw6AcWla7upgYo/A74AexJ4CZ9XjF9qGWgbFyCK6ocHsx9UYEFP8/
ofHCmzPgxQz2ZdQuHzTy2DbHZbj1/FR3LF6RAUfphkvGVYxJUUoRFeAqrPimp7+A
cKKFZ7EiEY47fUUGoK4CjMXGm6UXIFx6b3i3fJuDVk3vwVWV0f+lcJeZHNMb+TK8
JWyobL+/vt9WLjp69dmN3C8CgKlgppIOwftKgCCixFsbkgVh7pXpiAiKJphZ2HHB
tw1R+qd3puWfaKmjzhlcUl20bBJNadAQQVVVwD8qd3DfipSEEcwDDPA+VcFBiTA6
OjEEgqNX3iG01ZPKyotKZkTQIVwZdobUIoHgR89i1uI/im4/QpMwWrexFYAjZdsM
eTCoRi+9Hr/u+daspWjS+BYqZj6yJlkPElqzSQ+7mWyMw+SDVt/brDi4VaCHF6o8
g26pXfSD0c/CzAQCsU0tl8xDYQtNTwCQep1YUtXzMpyXTF29n/A+THF5VJTMXNAn
gYTdWLKfTuScUmqzBroo3nHZd9AirWAEMqKXRt5XLtTCfBWHoclPBNB9AInPQlvG
Q7FV9ustU7TiWMNp0A31L3f5vdAmEyulPKnEiUl3BB/erYExh1afWV7Kwmrf5uIH
UCOnpPKbTRtdLfkpd32VqH8xJP3Tmeo/oSoCbk/PT2QuhOYwq7AJojDJz78v48Op
Xgc2Ecos+4PM/8n5m5P+AWAuM4dhym/4pq56ehQBWgT4XzhXfDEmXNi4uIAdrdD7
TnvHG2SJxhjFptsJh08/CwI6bDog7f75eY1ILBJcBKB/3prMtOvu/FC71hckq+OE
u+EsDHC+25W+v3zpOaWkPoGwbHhv7iav4p1bUx43cQylIa7w/mu4FyrvesBbbbFL
Yq861fU/gWu1T5pUQ6QO05HZ03ZQFVVSDfJFv77gc7XNoDvEt4zet3zxNPxgzCD/
fDreiz+IRvnuIabnmTSpXpRMaFY9fHjs2aUF9fbXGtTOaohUO+fth8zFfYG809SQ
W2FfeteM1HlwruckoeuD9GDJsrwdoprPQhdsIn4K3gKTQNYEGUhRGnimd/N0vu2v
cYaK9uoogXEGH22WIfPn/Rd67ezylj0YsMb2O0prrTz2v7nXedfP3dftA7/HzBvX
qkK9Yw+iMH+izp+KQEw9SWiaws2HrxGRIHMPj7hjv7DK29a+KcbswXjVnIEMwxVd
bHhc3OjzV1GhJg+JQBtp36NzAe4UEHRLXMg7ZBO9euZQZ3WrLL40EByD0V9atkIl
M0zkqk8GRQADz67vSaTBgBENyW5MeivkzsSwCSD1434H60JVHUruUbS/hnw44X0m
8X9FrN4y4FfKMx7hKLy0ikExJ4csNOCMJCbc69UFH2ddJ4Gd2lQFmvv7zKcR8kiq
oGBRdQkadG4C1Q3Ax777q1WCkmIbM99vKGfJ+Kjkzt4Z12QkfSNa3z/ARa/Fb9XF
SQe95Pyxf2BILnY2NfBfavXdWqoi/BMrSeW/QgyztKxmrODZpmxvBt9WrgGPFNTQ
OLTkmPBJ0UewbQSrLX3wypFe10irFf+QCRJwPdpfXspAHjptxvqlQ7a9SAzXBpuk
K9AWqNMl2IPKZHe6taJqYoSRVc6HOsDilDP5MjQdFN1+RVQX2feRcH60dqFE4FUu
NUJrln6rdAoyH/+Z0s1MDVAvkhP3i9uFKML8yJPtX473ZFUMSYKACuvU9kK+aLIP
SJpEUBnuqhvEuROzfkNIZC6aYASrVFargwTFIdw0Ug8b7vvUaMhRqHN6EuSpvB94
J8BQaCiboKzk6fjB9hULv1ertMlAAq2qQ8JruG2j5SI5IikvFJw2dqaFcDwN7orr
MV8MXPVUyf9cbswJTWqzDMvOQ8Ze04E8O2cF5xzPQQS/KOjvznyEMpldVV+T4FCM
S7FYHTV4ADAe5fvpT6dgcr3PuovQszOzns0ufEOc1Y0PJcpxZ9FEgVwurx25J/dx
Ftu+PBj2u/fSYJQCqJJee7MRtN1AMT1OZZmU8xmqZIT5AOXYGxXdkButuUM1H+Xe
5PFJeIiW2lxAlpvvXzZ0QZRpMrKRNAVQG4MndkSAWebIVksOMRCZJ8SU8guKfrqw
i2gbwJxoScmyJ5/FUPsPH1xY50cb/HFq7GkBOCs1ZeqxhBhxmYT76/j8dZWbKajC
ccaWIyDiJZbcxeMzGBrTEulqoWtLjVYTagmQqVZEgg/d5Nk8bLMFcrvIo+LQPINh
TUjNsyfE0fktd0F2RGsX+c2dhgzlBv4z6ZrzV/AReUvC970km8gVnrF3lpmS5h8+
UIhDNkUtStsUBfdgXla5y+g7cZHoIe2dBDRVmxFY/iYuvEtLfDRh27/D8TaLIfFV
UKANQuA36/A+HHB3Pi1G7JvNLD6YKfphPEAFkLTxFkBZBE9LlAkr41K6JZGwHESp
PjBmH/70qZmCHnWj74dOefLQiH7ywszce0ksb3MfiLUfuomaBf5LIYt3ycT/M87c
+xFI6KdU9K/M+agsoOzKq5KjlhFtAXiKmN9ZauRbpbVWnDnu7JT4n7Q5g+48FEGG
m22b7hKSbAMAfKGXo4Ksh2Y1U1ZYyQJ6kFloip3/Ggm5EZkgQrB663cfD3JRSvoP
AvCv1X1AjgfN1iqSRJalSUjJyVQL9qMnxc6Ll20dFuGklOXTdMe1qkah/23tuXIY
yLNiiF2S/TM4oqy7J7/3ZNHdvQ+QXbDQ9RTZKKednderLJo0VpUFVzfdeQa/mJQa
IPQ0sPA9zXf8C2n51waNtY+3dlnw0befgBJEiPTX+AbuJYVhZoufVVjmUAL83+Za
pTtjifUx+X8HfUXG2K4ZQZIJdxv9oJYFYnRph+LxuB7VVWkAnBqA/JLEHznYzbPc
1wlLeDWN8o7kaQJvbxrWnG988z/j5hUdriGPKWrB6sxXiCifgV/lzHO6eJy/TAPv
8vgNso1QQ8xG2Sqfrq68VIyjI2pvsqhIALRseXAD16h5b1cA1UE7XfgbNApL82o+
cTiiUTDEgUdZRmX7MvSgfqHSYP7WvJFZ71SNNYAF8+2SusLahrExXJT7VC6vFhmX
WzS2SitBmBN3OI14E5bAY98+GkIvrIwErIQXB+wagBs/z+6PqdXDs1h5EoIbv4Yl
AJu0xvgZbiNhQxW6zZGTTT0ZYd2/VnJqji1/WGs/wtiRxcpVioHHuFlBhDw/gAZY
ytUshXKl2BWcy6d9aE4ggDAstRhQ89UlQRmYKwr6azaA+T0MEY58M7t4RtxGrACG
aZXkooSYejHBEYTEbV6qLlv8cnX5qZ+VvrjJdO4JrQLDtW1mN1fSg0th+uqwVcIm
fwTfk2eZbYvtgjwSHbk8DyosayvArw+aTYCXn/xRODByhq38t/hgY8PuRDrEZaaT
ztaqxHq3Nnq2esAUBItipqiJLE8ttajkZvr9y5TPJKydckpGSG3krH6gWHD0BLuB
nQh3Pi6adTxEQYI/eEKX2V0aYbxpvPN7V4VIGeY6x90R1p5pUIY6W0UcscGSGePe
zriDMGANgcn/ixTb7ZprGlhm7rXUHkLDZpgt9XcjCcghXB2VuezhZPW/cqr516K7
g61biqPCY3+p3/WWeZwuDhXeF3Kcw7ruQB2qgbRNv5rtj1q0zvRPNyD97RoQkNe+
UvtqVEV+8FM9n+8/Ur50CoZQzE2HEC3fS9PeLN94VieNHPUI/JbWqSGMv0VxQvFf
/E6xTg3CI4l8NNe4dkWYawRYhhA1YCBP1An6U1HzNDcIMZfWPMxjjMabrloAbJxb
8xoVX1kX0IYWHLIJNDQTtgjU/kY/A99lZI8g/8Ggj/Nnzc92x8/Dk2KGt7CO3UlX
m4jCSt6CHuv/aT9AAwI+f7HZvYE77b+J9omMWzGSewmxRWHc8GN+r8VA3vQsk9N1
43Vd/4/wooX2JZ2Oe2orw4toYlk/Fgr4wFe/YD2hYiCotCZnAGSHKMReTCzbg2jO
TQsX2j6Ob+gtovgoIivzUXpP0fN6nufWpNsJ1Boqmg6ZhUh1Dziqq8lPjLyrknsw
MTYFGxtho406y/pRZVXhYihvj7yeGr+STcfe0St06iwCa6foSaHxGOsMfLqIwEmg
d3j8EJbRMdOYhZwGARCRT/ZzwWJvmOcEg++K6AXGbjXkB2xeCW+jHh0KqnwDVqxU
Sh++mrB2z0R8Wb9qTI+LUXUPr8kCYDKetqqA7vmf7Tvkam5jRLLQXcOKxUDiN+pp
s5H2xhgxFfVKMvF1z8FugRinfNEZndaznQlArdtxHeA+Ot0LFboYVEJVvJSiWV72
J7J6BcmrMEwrGts3lot3/QgcmdNjArWKg864RlwH154nkx+pNHLI6X5q/gmvssxM
czFngZz+CMscm3iyMraHdnBFiERQm5AZ9HtTk6/JLDaUp+t3/ltj1rQmQaWo5kfF
pJpMT4oY4RdcceK+45IlMkzjqn9GfUt/qGrPhmSChzKBdKUsBO0SuHYU2646SrKu
zVKB1r6Wthe/Ozo01EwfxOqA66di3rhfZM3ftDj3HJns0YPYCPQsQbj0TIxl3Oui
2bE9LPSPRdVqGjaQuFoeY/FH0oD5xd0xAznFeNzmsSbV9OXy2hF51v8bT9i13m6E
V3ZWZbfZENDxlFnpwI6lnvsCaHQ0l0kLcQPA6082YfxaQ3/0k/9zfJ/H1IFpugRh
U/0D763GIobC4Zsa2x+dUy/3YheUm5ZxDxDHyX+5P7lLX07TDgZ5ofJg6pTnTUzv
aw92xFf1XRUJ9VGcrbaJ4/ULKbhepGA0DwKASfG61Sb96UP/b8OSu0RWbZ9zrgVE
XEHlbhPVNgegWR44uZZT+3eZeo9vZ+vU7uCBduTEy5UHPdJC+M0kSfXaLTxLKxUi
CIPV6FvDqQk7L2v+Sg51fjHsGbZPcJZL3QoRtIETCRPPiZDWyY7fERcGy9HgzdvR
NBo8UsqsRIZWcPc4JGErApcdtk57TLpH3ot35v/eTiXythyFj15HTwXg8MEzxprd
JVxsK0PBXxdPi1QIQbb1nzSJjGdf1GIvrgWlzsr9g7Jsy37ltkjYr3YPKF28TYZm
PSGPHRODy1LjgSEW6lEg+y8vZsujMnlYzrzhW9bY9dswliFmhqScP2ROcrX19rUg
1hrXHjkF13QSBH+vQSGdzRS7+AHFwGwEPBKBt0swAhVE5KqW2spZFGl2MM1QH5/l
HdMZvIWtnKO0o2hiXp1024CnTwZoGDZd8n32JG80lpTO5GqmLsnTCF/euCQR9vTs
YjINu+YDouKD9/W8Cngp2XPKYScWpjlMc7T1aGgg/PpmJa2PFZX5vPVuxsos456a
rE6yys1HtopgL4TQ1GhHChyN5nTGmicGRZCz8g7u5yiZE3SAM3wLWrvPh89yrSlS
m4qoRc5//j0yoJVMsbcalEha6JtaAhUIeEisTFOWBsuhegMWgfPx1zjR7VOiOB+N
RYQz2d+OQjMEDIQ9OpwMM7hiwMK8poDapH63xM5PWqUQnJMUMPxvfytI43PdHpsz
dcgBGpy/GinZq3kwVtcv47iQdTAk/SiuuC5FAl9z7U60EfOQuTbQHLLop+ID0Ik8
4mU6l2qkgjkvuuHbIvEgws+gI1TFvjuM3bwtNd4zx9q/GBbYwCdEWlGARUzue9ZU
Ejvud6WCBPlPdihBCEKlJ3KX419HkdHJ/tkyFkJj5PvaKL/kkYY+s/ZK+mkUCUOU
Wg5AJunswWUe6fMjLrBgW+QKyDYB/t0md162qJeN/jPkVMgkpkjYLb3Shb+WlEHR
uudQbmtXL5+BEBUXVBBoEenenXlzV/eAN+zwetPbi+XF5kjxOU7pLWDgC6B3GFf9
d/I9ouEFTohqVAC8ZWwKjAtasJOadM/Z5BfE3wemBw+8QQKP1z+6QkMw0I6UtHZB
YqKNxyTYs7VCO5wVuA+rOOlmpeMAXRQ/3br9L+w4gxkoKrKhrEyfsXS77rqja4iE
aoYTRn7UQQKvFPCCIbDYPfE+s8we5Fuq+AUWBcx8tvx2We7QEh8bY2MxUNZE/f8l
b1fG0XUZUcXSD+zFNcdsIpWGmIGuwGHJzxm9PwO/ls2qGdT5CflriyFv7FBTP47e
MNNkOaosHvIo13jGtv4VTlmo68f5Uq0tYuK8/9vBwHtvmK3wDgu8CqJqBjJ2RM/k
ErDvfVKu8spOg4oIC3JOjiOVK/T6Yz1XormOyJKTr9pwGmB8da0TOaAp9OkG8EIO
SvOFjLuJK9fbQPZbBzDT+sU+0kSyn9QoHc1rhWiwqYPiV+Jl/+yQ/8gRKelP8NZ+
fYAzzZFjF0TMuhACN9hy+y4HfGGJtbuI6PPh1D2kojqLM3I4bcucmP2+zIabyi4u
mxCiRCv3RaWfX2rlp+59dirUdRfJmwCbJL9pkOcFjn6u5Otm0mB73yntHZLr7MKK
IW8N7ntXlZO246fmD9dpI2ruIdvWtRalyouWN9PKkTTgUEjTA10v6+aEc5JkWbIn
7wpiQXyFpR/XjW2wuug6F4Rb22vx8catJ1stujhPQ+S/1pszYNOtrYq6gf5zkNtr
K8vuLe+jILrIIn94rOetAZSrI5l6vhVDZM+qJi1Angg54jWJ2QkWDC4NFnFJYtst
hcKI5YDis4cIQhNsxc9NkWBSnN66PAleA9FELjn1ODNaFg/RRJdB3TXb8w0zXn2w
SXKlY9xft+7Az02gLFTWBoOMhcC/nOTDJsfEpFmB6tx7YOg5JtPEfullGw9He6tg
1xRBAHGqr0UeTc/lHSdCb98Y/+bnvQfAK/zWTB+nAi1T3peLL1LnJQwTGN7Vtz+t
wzjFg7tm+kY/VBFWAhvcfXfpi1yZulmLLVqXmpdia7rsTNPhHHjJMAgfARKudU3F
lPHag6Y6yXZ3kErh+2jSYUZpE5ttfspSxiNG2doz32WSG5Y8pAPXnR5SQaWGrZlc
igKkLa7JvlMGPQwa3rFJ2hgu/J93h0GbZGd9QvVYbrUqCRHU8RQyLw2Q3u+ZuXmX
z1nVXK6hF4GjqWfujoVFgiOzO3YBUGyiSpJBrROFzu1msLZy0JapDEQDSD+Y/Ld4
IHIQ4l14CtCvtOrqm/Ol+df9jsB1KeN+wI87R5L8UG1Sm/kp/zfyBnJ+WZ4pG+sI
TxEwIeJNzEbU2OfA2lv4z961XpqUkU3hy1+VDZ62y2rG31vNQcjfVYSJoJyZjLJO
KYYtjerhtbDNjLzKC0UpxtqFX0nwhnBC+HzaHy69xNS5Uad8jjkCBez2GvNviwHE
SNztgP8UHSFS7ELu3MGWyGIDZADVjq35KRwyQSbi+mS/EbJ0Iajf0xYbnUjGJuJj
/qa6vhfei6gQ0yXsMgUm8OPEdsczR5clZiP5pPn8rfmyFdepDoWCbc6yqFTYuR2k
1HowmTBe528ZGrP9hS0iii1Y/KqCMiz2qy5QdAQr5CHtI3EokhitaOXEQ077gTUr
zlbUhg6QjbRbA+OSWbELQDgl54/EWuc/jk6EVWZEuVdAkfcj7HheQK7b6wP5H9Yu
83TXgVtW1hR+blNuLMLTOoseG3BqrIdR97gC+C2CPXr/EP+lGLCTJ127tL67rPbU
r3w5dw9+y6ZzAkoS0OkpzBBaScTCQIEOpTw6J8DJMnRQmis8gX2BPcOWKe/1XK0Z
5bIOXg5aNWfV94jZg87gdNew66K9ItJm/Wolei5AzHsgp/IU3Nn8goUHDtOTmtRp
x6CfT/4CFjqRUCLUJoa2IXwxuaHXdape2bDMPUOpELF48+VgPkHsityLP4VCcvp3
MEfd6AJjumveA3jKdJ+xOtSawLZuDv1cVBc3Chi1aOGjPI2q4SrVhmlcy/7e4co8
fp0nVkrirWE2ELrQJ5lrlx6N77wvYwfDngxhD8TAF2UgCH8EFhPD12GUjfLxk4+X
133GNY9n8EMmXMh594qiE1B3lTi4mCdW+eUq2RUCQlCWVoHBQPP2929HI9ncmQzp
MM4TCXqZ/0pxl0iPn15TkH7YyAvkfzW7tqW+Us9GQueOL0eEq/FlLeSNjp2OuVSP
AMJjVKCRZBM/G68/OKSqb3FBxk8vuCGIXr/xDxHw8cvAJoIegBSjppsb8iWgSxEE
s0FEPLpW5S1noPXPVxSd/2iWN35yTM7vNaJ6qu0kopCpHVyf283F8sUSFfPGSC8i
MpRd/ggNt+KxasvLF7UJ+Jc1PfkN7sSQUozt8Q088rEdL9MObSkdvbh3UGr8hnZf
93L+AFTcR4EqbYy30Znswtyt3q+HWGic2ePz9RVZYJuKhnVtIaQa+vbThgHLAvGL
LmSjv5RU8GnWocI6pVpuzjrxXS4zVFZmASDu/Foyk07/fi5GY78UgSgmYWjDZAVg
5LyG/aQt94p9zwuVgWLTCY3mX53XEqC8jfdpn+QuJNS/FSgUE6g4kSLtqDoZ2XL7
d413SrQ8Pf8DbFn7ionwNZIOYGucqFCaVMQOinsoTItFQHA5RIUzn7VPeBSnPPIN
500m38c9madf5e6AKXxdq1x5cHIIFOm7gTcXox2Zn1YFG9AULoVrIf4goVbxcFzo
7aiwSoank867ilfGz5O13K4bKW5DO+zwZZMFWWgS/IQ9hZtpuU9uIgUr7Bqz69Lk
LaqC9JT+zI7kKkcke7NIgj+mKl4GEkx4y6v7NNWe9OLZOei2gm/XXGdjuiUDsXOc
+RuiFSe7jTBbHQovURCmX/J/pE5CB8LsHCHopp0PF5GqtMpBmLPl47hPWUV2NCme
j1/m1QkiFqj8iFHk7rci8t8+sQylL8fgIWomSkTsDJUoCp8MixE1UZ8h3GyIe0Nw
09GYbnxmA1qEFXNGt4S6zwfn3yj63uriPUP5PsqAHg3Mj+aT1r2NXGPiEzbkfbFE
mqBB8J3/X2H5pt4WOlOxtZ/fDd00uD4elte9z1j93FbG8ZueuMWGfc1yDlDiLlO3
NGGNkr5IGzTj6mLb/22B/jCGEACl4S+ZylhOhZEdbU13VuMBtLPNyrhr5S11iQlB
wkwV7vMqGMKR4oOz4IZ4ENH0qV7IzdfpqC02cGljGyUxohNCQu6RveLwbOEhAY0q
IzALIwbC6lLQz4e1hyITgDw+9fdtjJnriz8qnfjx2mMWfDZq9geWqwxCmqIa/j2o
JRTqIbTyBf6zkNWJeZZGntEtibaR+ge5rlx3MYN3e0ySx2WK/5+jGqJzKrx0dYLS
3FoaGOsP9wbuLM5heRgAUbQfFp0gAeV6H7OPJqiXD/oon2m6d+PtgK+8yEJj5uZP
TKJzn5DuXWdLSel9yZA8cFErxOuNA2vWwmBJFWSJWO98iyKcDl4wqu7eHU+3L+0/
nqihDshtAjolfNZKTJU4k2WfH4flnLAELOP2mon7R3TAYNYOCRZBrlqNzb/eLPvb
lCM7YN2gnfThEdK8GKQPza3MIg7ArHGD/UWIl1t/B9GQ+D3iewgcqV1bylxu+NtJ
r69eZMmRzB+IEfkdyAv3JB5SfzBuUl+ut3pAu2LCS9PEBqT4+mg8ahRFAXDvwHOV
mUSnpb+95JNonoo2QszQXmPVtTEHGBVWEpEs1mfbvRVLFsKdckhCrB9wbNnOCjy2
bVbBJCo1S0laKpqgoFqqsnAjfUzIRa+n1esB0UVTfn0kK057BV8PMXJAlVTsBj5r
A51j+oxu+hWBAODs+uUGu1gVAiStTTjd+3Ym8NV77rWp+Wv69w6jdQVTAUHzloj6
onEKsZADFQQdmN/uy3zUNvlSM198KT4/U9w1M/yS8wlZqDpFut4FmPOMYkNH7qsO
8Ez1mX6V9vHqIUieldfjlYO3xx7uYNW5UmHq2IEyy0WNvX/P0Uz775vVoyQDxsGm
yPFUN/hJBCHd1JrbMqtR6dQENuYPyceucZrlxV7nuD1neI601RvS0Dls3q8UFdb5
d9AbTkH/df2xfSiR+sF1PsnDqjg/UnGhZ+je5rHnmT1PvpH9eRij/fcfsFFNzYPw
CDlvv50MlbBS6mPdGFTAQKPNIPClBztqLCYE09MmvHsqWm97rfKCRJVVG7wt6Y+L
griOxXaDIDc/bglGGiCrB6cpTWYbgtF0NeSWmZ29J43npRLclrEzE2El/AD0JrOv
/bEvH9evQ5FI8gBVD0Wb21scMLRJvxWfq7xe/xXI/GH4gb5dwksjH1NZ72o83Hv1
gNBUf45/PtubpsYKP5e3P472WImX8uer1r/4AubJ+GT1xutPx9HZ+oF833bkOOUA
5hpXS4OAdNAAXfgEfIpkvSbBrUlc2UdMrikSksLUHAW3oEqLomQ0CIbVV0i+oDpS
TukHTYB3gwFfXI2K6kE/8Z1GqbJtvIFi7A6aIKG/l5HxqIpfRfpkAASHaDYC9jt7
ExCwEt+iigKk8Lz11KZl5rKdm1IShdoJOV/huMEks6h25I8RJzJGqZR69oEhgmxE
8QKkAvmH375qKVrWLH7QCsgQGkl2RI/uj4X+cLaNWxcyKpcE5mSlvOJ2BvfkOy6j
lOwVe4/FIIvU9yHn4z0bnvqb9EMqXsSiu7yMX1OjDcfCJBpixkOdLYy6Cm/8w4kx
5IocRvJFKjG0luXexXcsbv1SPgCYpN0bcEB3SNqsl5DNwrFMeQS4gQgXR/ckMui/
U6wl6DjckMroPhfPSZAS+9dnNwTYjeU3vZPhg09xNhc7UTqdrihqdfIzK/OZiXlL
qnnQ2MH8GQjSR3Of+8JDqDTcdWHtuUUae3nGurV/BI9GBrao330YfVc0qD21ewh3
tjP9ara59/Ao+inqiLg4iEuoJFXdjXSlBHdtLWRqFtUbZU/RThbN9L0Z7IQchowI
ZUIMj/FW9Zs7pMdYCqEKivwhQEu6KshqDurOOpgBNbX4oxWEPA1YvKIyWZpXSNXv
SBTr57Oxw7mpPq/8htu0zp1io2S9OYxOYBpqqGmyrAOiX1W/qmXHqeuAVJY5JHF2
52lFKO6wMKyc8iffRbSp694MaBebxCZ0lx+OcILlH9WFqXl8L03ZKkA/rd2J4ouW
rgtOn8Hs5QeZkr2+3lyxeTBXHu4uJ5VmytSGHdFqq6xacLCUSZus9nYwBluT13vB
E0o888fKakn8+FlgZcqiaCrHyopivznrTegKfTmnL7+9c7lsOlaLxAgSZd+l975h
WZZ3NYXwa7wbFDrldaYhCDxNIeGjzwtRfPR653vj2N54D9H7W2LSOGWkI4T6IPec
ArY4R9IjLDsO1/TNtrsA1FVntW2FYD1cyy87Xd/q2cNryo71A7pKeqWhh7QhC60Y
A0kBFqLPT96ax48h6KrN5xTj3WNHrpG3DZpkO2N12Vl1l+uTImMiwf/g6LZaTY40
n+/owiuheuah7L06+irPh1ci8VAqy2OJdmFMXwK2JCvo0jupMx8AeXs9W25hTvwB
q7DaJjQOs3EoxjtULuupq/Fv0JWeMPLwoX+JJM5Y1m1Lwi2JCJC939IVeTfAglwB
VoriDB3RgmxoBzCpSNk+CQnbamqkYJMKlP/GXwkZZPIt4SESbfM5sqRvGITqFZ8k
zZm9i3MfNf7RdaLL3Nf1iRzf4OeUm23tYVOnCQkEBNubTe6GH3kYjT/NmC6iftVg
+O/WZShTSKhh0hhPMbHyx1yGxbFRyw0cUQJCdQ6FpDaOr4ZmfYjKkSThho8rYnpz
UEjhdg2BexbKjhMngBt/BIpdBeGHFK+tzq7IqFENJNhLkSNjjc6aSsFnhL3PDfo9
8iugobhyTSWK5dXkDmQnzNY1g2K9V4u9YAabiL6v4pCYHkaoL8eNGhcdoR+LZNAl
ePB6r/m+yts9TG5TZEbQ/WJVPg/Dr4AlZsHbVxXZV4JnZkHqL5J/p6fVWhyD6+bD
oGuqF0fMcKAAdeKmyk3A4x5Ea9cVhhqC4v1bZRwWFEGLGpr19zzy3RSbNDUda3dy
hUzhMChUPgSCOeNZu6jy2CJJg+ZYkhX0M9rbgqgk0COJl/FuF/Ubdkd+3T3DbsvV
jqxQDUscGciSEWngKsTMbkC3Zhqh8vYkTTc0cS1GqvtHy5ROwNtpLm6uIxAXipum
KiVQIE4obNhCj2lRFmEUZBomiOIWZgAPQKYpq8abEO4jWkxOf+gfe4z97fT3mdy0
OpIuu2+/txNllYZUHhJKvSjGS+/UVIWVtEn/OAKBqMJaHTKYaiHP7TQ1I8vPbeqH
8ULk1pSjyS3HL6CfYGkCrLdMn66t7hZw9N8ZXYh4fLlc1RIxuXHWffT6P6kY00M3
Dnmd8VdR3FHdn/kkhb/GLL6GOLeEZ/n5ZNoiLcrse9b45U7sHqy3lxmFOOmIkrYB
d+XHWIIy8F3Q6vx/u0ZnqkmWc+IuOgv2EmEZFas8umh5H6WPcnGMUjA5J2BjmyI/
L5JUagAXC61bUnC1meG5VSz1cq9Fh+7ZqbKpUPsmG3u7hjxkD58xvgvZrTUWUdCz
deT4rDola5r2yf1w7f/54Ajlb+l94KLYvy8pYP5Iv6hONm1ns4Ez/NcYFIbjqUQc
CqEysunkGZ7oX0YFwx+4jY0jwXk1RgcsTWeErqWg6FaCFQWXp6rxhHiyHo/Tr6Cl
Zf/jknWiZkwrLyZrQoojzkKbZm/QLFKqgtvbUUfADYMARWJKuExefHFodEp20VUx
qf/LwM899vmXBdr/QJqtFj7HC6u9paTxA2IbLPCv+Q5qALD2D/KFaWn4a3gFCv/f
I+MEgWJQnGhbCiGd2iTtYSwPkRdN3CZy8it4ZxBVyFj7H8q23KM2z2uJmSFwLmUf
qJ16byjFmm7TEUPUiq4pZ91wi8EFA+rm91KiVRI1oRQnSQzy5IP4jR8aqHj6f1Bs
lzXEngaco5OFGcPLusyixg0fFjt+OYx49KkuE2P+ds/kgOeFX6BQ43Gu1L75QiI6
DOWFRXgg+uqJwYRVU0K/eXPon44gW4EBn5mxwO5Q5Bxqk6KOxaYNkqJ3kkDISPUC
2fVndTN4dS/CCENrQ2FEU6WhCn2esizxZBZSfN3171ylHqurDY5qnrBPrvZ3/Xee
gSrOMU2t45bvGfhFqJBAlyyxIBFpynEcIDq7OpMPQ13oFLLXtbMe212qIy8x+fzA
iWfJdxMCkiBu4F75b0B1bDZwJvYK3Z3bjBneGEIzN3TSfiHMYD3LFG7OGb4tim8G
w0rS3inqxdbHn6pJAY9qwzSi6Opc+7CHEjqzP+pKinWy1EXvfSLOfIr3U6ABSWS1
Z/mESPTdFRRAEI+PhY/L112EVb+oPscNuju93xgk2TsSPRhLs+YioUYrsoQauf5k
+BckV0VA7Knh9z0NpV3EromLqvCptl2Uetu2PtbTTBAc2Dph9PhJjth5iWD6NDWS
WGyHoRRv00sR8J+IP1ftrQilFsSB7DuseVyfBHtZ++FBWR2AES15tD9vMeC57rzo
690zX+1Ny+z6feK5AWJpVHs3AieulKgI0Mn1LIoEpeJDYreJzPhANvUlHE9sLuDQ
O3pQJo1hxcE9sQZVO5tDIIyBkhW8DHIduFy/icbmPwUtt4mUjpvmbeItGUBw0jJ5
whabpmhsixK3iJvtYZBE+81E/zxt0CF4vsZKkas61oRSaye+tW7G4LrbeD3yuX5a
guFVpEjyhI30YFx1iI6CIH3XqHUQGev772/IYcJ38FX9f5FgKudXY4vYu7iP97s6
NeGPveXswxNGjT8GWG/tnbmr2MB9ZclEuaSXLuw+eeH8EVMiOHseJ5Waj8vVACIL
tr3nrV4YLnKtXeigU8TnXn4OmBegOOKRc7H1qUee8sxpVe3bUZxYZDUogvmZe/aO
r9M7EnEv4EbjkGtMY8KVyZ7lJnRum6mEmPV2XwCqoU8/Z6ZVuhuElw+ewQvnrRO6
FZ8KJ1xs5B1h78OR9kpdM0tUBkfucx75hzKC52zAGC/QgT8+oPdPvOaIF1xThtIs
dp8BF8JUtGWMJqREEQIfzYIgkG8i0gK1E/s2z2ThjVKmTVN8G6UMv5Wl0Iwwo8vy
5V7Rv88zC+e/WR7Va98af8bf3ps/d+MEKIqpGBOReT27xA/jWE+PKYKxGGwHjY4a
b6pmJK/T+kYZwqfv1+FQY5Q/slQrhBP2LLDOu6loj2GW9MCxoeDpNYA12kE2tWAq
Wt1q7M9Dd2GgsFRGhfX6czMAeGSz170JjpTgBz1+ywiJkRzzTZxjjWhxNrySXNhq
V/bamwWliHb+AjAOLkX5+IQIzYWGaa1GRvvqxc916KnbS2vY2nL41c1wrw0snYa6
NHnne/XfRn5ShBLw7jfoJ942F0wReaNWMa8iYyHUAuAJdu+/l9YGeZhEKvY7UBRm
WS+BTPItxzWfBhtH6IsgLCOqsTVK/P0sgVBrZkgG3E5h5P2zBFSugulsB/f/hjbK
nZO9WMuk0b35UPPc2eR/p/NBx42Zy31LDrrokHmp8iKN4PKu3ZFvR25AjVJoNXhc
b6iIVItTRkD1glgH0snF9KrllEv91VKmoJpOY0PmeFmuuU+CPZVs9TN3rEtoiNBd
rxXTMwFD/oIa7Cu0WpYTZwHmDsM8upML67WXfDoRMJQvMV2R70+kYFSJSlaTYojt
aonbaGWWt2ZYNNzANrwdBi/otsIjM0qItOrzwl+8bl95X0R3XBCnDhLmt/vXVrQ7
xq80TKGDhgx0RvXcsVXu4PcxX5ab5yTiK8uE0GL2gm0Z3fNUFhNTe2psCRL4zJJk
IyH5iFjuSbh+lBA32QIMJTUd4ZGhzbuDdZIGGMcgigIb/uYCar5jpEFSZbKQZngk
1dzuPyZuguqfkSd9G6dCkfmo2d1Mm3Hti4yHn/9wlPXqBKqdU9mETgT7J8+gODyh
aQbqLtUcYz0wOuW/nXmoeBWZA8lTZra4zjCh/q7CsTSO8irOhKeyvOmywVIQvF1M
X7xz1tTgq1MXCmz2kZy3kya4bg/TeKZbSIKJPVyO1euFgMTbzYPue68ufC2sdzGg
BWeefcbtbud1tHiC8P7fyHS5GdLauJDLPeseunZtYMwkLh2adQOnVlBRhHmoCXZj
oEV3ony8PxiTCkr3FF441VSikKW2SNYnhVyQETdb/TyRxIhmIkmO0VyHCv9IZ271
FTBsrOpOssf//HsVzmwVCl9GJu7LlII6H2KE75ARuK3rq7VJrOuc13uJoZ/mfG/D
ZMaiXdCA2cSUG2TmCW3fSeXyl1PvqmiMuDHjYe/pRaj4OVy11cKIwJjDDqZBfvEN
t4wF48WOSD7eqU8/jKvQTdMCOgMak/spirkURIRGSiRgSMxQMSEZqoXLy+cdzZmp
rvjcUR42X+h0s0q/N+rFclgA2X9HkF5C9QDg0HCzf09bRGclJJNn4yb936Mys068
JegqWw35/4tG4vukdtwIif7qykeiR6TMJxqTxKUr13zFO7a+I6GdVOhGYUuAFMgt
AtSFWVxi7s8JRSQQwCaSaJ82UGS6JA6BavzcQCqpkBGgmDSkAv523EM35M2Dp7Un
z2gePmPQ5uEfAVTJCvyiD3dKAPfi434wUDXYIM9E2hcwF3SZMZaXDSCu+wYwxn0A
/pTAzyeFYy4BQYUEyCuA4p608ovolOIAsAQsJCyyMoNfpaJDw3oEQaQZXalPvLC3
X532fvpE5PLjn6JW9+nDtgbUIVjkKQs7gYYnGzAhNMU96mtwr4ZJW11JeLBuLBgY
TPfZp+AXYcfncVJZzsGSt5aJmaadLv3/zxAG61DvSA2ubVS9X9U5Qk20qvi82XMy
9sOPgsggzc9hzzB8AWDCfeTjccI27DKvMRp/Q+k4PSieVERt+bGPq4t4dqteAjO4
z/5hOL2L83lgDpiDHPWjSGBLTEGSPYYyPYuZRuBbng80l+4nxSDLHqkWew2GjXt9
vnneSr/ll22tX7AZElh/GWJLNKKBW9jgW34Lum+PqOKJusEMCbsPsDKWVpnT3CaR
vkJkxCetX8sdyDcdGTvrS+AVOfYcEiEMYrnHSzHHJh5PP2lH4Ryga98Uoq0vYZoc
Z3L3aPFBIJ4Ir7NV+rrm4RoYsgm7YhethC+dkYUYRFQWFDQ0I/Rcb1QEG1OqdpRV
opOSynJY4Y4zpY9FfgmpKL6+10W+wvVVnJn3BHQuZZREjapHmNzuMHPotOdMivpT
yRY46tGNAB9EEHAOCFf8RXAR82Qm2hFdqtrQCTPKYls9FW2E6Vq+nY1w2xuI2bZ5
w0v30o8eRzz9t6Lo4UB9MDa30yD/qNWi8/FwYifM0kV4WIjG5SzxYoazdJLjGJj8
o94zV5qo4oKHZ2rG2Hyxv2IHBmDZ0WaIvU4XpH5l3KMifAT93Ep7HAM98Jh6t8+g
6YpQO5nGJhhmY599N6tGzb0kaSpI34KSbfE09+9idzW9ujkgPR9GVSjdO/s68+Br
6wJnhVW/PYL7ddhYS0sl10y/lzQjpqaBHqS1Vz0MWupVfF+efrh7u0nomdsCGM0q
exPNlDIdMhQpcgFYs/uWSfHbePNNzZ5jihPVpYvA+WmQTxyzcoGpc+XcFooBTWLh
RNxejpkeA3Ga6BjYU1DCzkWZjHNlYjJIAEunGVHRS2jbxYYBcxntaCefXOGutfRj
Gg+cSKNxRthq31i97EBqLYx1cgaMt7rVtelNKRRGh+nE3VPW+0tUQ20qmEXvE37K
+jDwJekeb9Kz1R4jN2XpM0i/6qoHHDvICMjISwYG7lATKr6J+EhNc21k79OkR5Qk
A28u0Nq6NAtV1S4/Lh3o5dW9ZsMZyeDrt7jN/Y6Lkc5TzPsxpXfC3zw0AIpM6jLa
EAEuJjysVW6vVkgafNrIO7w2RxZ8+zm+RlFxA5xIsLrQDmzzvCDsVxw5NZNr+wWx
lAIaL08MwVx7xrxN5mihY5RNU12TBvHCRgTXW33kRSDTxAleVmXlITaJYpv2IsSW
YsBhdjY05b9gXeD4n1heGJz/NyywdjTiceMSwnxcPoUqnCEv3ZCPS3uViISxizBu
9HVAzMuyxoCQ/I+SuZetnva9JSakS4OJ7jY33Ry1FF1B0zUoLZckFnPoGbBypA8p
LXDhn7pKHGFxKGU86e3A0ablg0szhiwZGu719j/Cb8r5CsVgSjx4RO/hseMO9JRJ
MOh16Imc1mDU4ZO2KNw1Kp1TUSfzbMK/Jrlp+MhxgFaVTacj1LbwNfb5OQ9iYFnH
Ehtbh3BkM5Yb7lKZOqIZRy03i+DiNImH72VsS64MFHnfRXjlMeSLSR1d4fjxqcPR
lCfZCz7xLixKQ77oPE7/7FCg2+B+ykLjqC1YHY4ufi1kc7FsAea1lPgGoMDvF5in
tN8/MN4+iFhtgEU16roOP2yPynDCYPNrWXdBJujLhNqwyh9aQEO85m36dTKTbQ9v
tcjFEEm97u94IbqXw2VBBfZC4S5OQ3/8p6VzgFnrQ4VqBk8YYR7F06UN2d2FiTfl
iOfu32zAS441Tabx7Rt2eA563ZYl/kFGwlP/evLFS+1yMwacKXF9ICvMYw0SC5j5
Rgj4Htp9qgrmpMrztu2/7MWRLJBBC9dlnSVEpUPbPJue5OpkZcCRCfHYhrV+FTGD
U3ENrCtpDko4so0I39bBHOjcUbfnNCcZR6tAxb2YzxnKTvhxoy/BoFTXMqfYPDcX
2q/M8LKCgYFA7eWaM9TB/PFY3eYMRQY/uHH6iXSw7YsCQXg6QBeYAAFSmQbokdtM
HM0Uhb6q8nWQPsZ/iYJqYMYFftn29XPRnF1Ab9GJWcMSw4+6PliOEIcO1V9f8n2y
XhiDHGXC1NoLTPNFwXxuk2OewS2xbzbYI7wUCKkTvM5rv+vOQX4sZdi+Y/85zo3L
a7d0kWbwXH1a2PwmxJV52VfXt+M1uEL8ShrUa2yQQdvBVB4DUTIIoR7Qhc3O6gJr
uXPgSkdZNSuQW9rkC2k+HkExh9RJFdM++IKc8AB0FjCdGNaaenb1RjucD7NKCuDB
nCozn73PONfqfVXGoMG11GqQuKABSo+UXPV9PF4nWWKyqWea4LarydcZS7nwgrpE
GXDx3p+2nOL83Ms/QFexqFJ+iW/2lb14XNMvhGMvHKIZfqCi2NQD445jNN+c2GG9
3Jp41W5iOcaam1aFo+6I30tSmfbCeJ2Gg7VlBkfSNZAKyeGrHLAYKrpP5o25IlL9
Hl7KgId5/71LMRr1N23a2tsJU1h14rUAjUUVrI/+AutWB5FbPTCZCxgDcl1gS2kc
MvWfJRRXoBQT3HqWn/Xj9A3epsqE2cFyHySPtfb8QMkHulMxrW77DtUZnZxNOySn
P8VzGKUcmRCWGgIWouskvWlHBa41gigf7sr1dU8nCv+0LCXxH6kcJRLuKgkGcFow
xShCdBpmOjQwEwf0RPh5VZYdEuwX68jQICUNje8GU7GigQgHfOwxR+J77/Lcuqhc
m5yHAtCTdJ8gqr/wyjXqCeJHJYIrA4Dueuq7UYsFwg9XPYz71Shb0W/iFoMI2NWl
auOcBMyHSXcf60UYrapwbIxi8XuBAv/bZ2qWv7U1BblH4414NreU4Khqa/7tkdlv
DotKSdOkXNlqDSE8ezazfrvy8h8TNyQ12AW/b2GlnoVkgF4sCoCcJK2KB7O2X/Sr
Yjnci0uGzJJnhtCCmZoDp5rP/qf2LkOaqj4x4RJwNF88DromyhDr3vPKGxlJdk7H
j1sWpuKRX5JmL08vjlj7D5QDErMoYip6+sGG8TE3+aYIU6oG5XYCTk4Fg9S2RSqx
hKQr5e5F+bIvOUd0GoV/Z+iQTq6cpLcQAlsU6hzeN8S1I/dYUmRwPkD85h/+y684
y04owvBOZs4GDm7rcePBGpCLVisn4hjv2Os7MqWIIlWoo+av41aXo3/7a4840gHD
R3GdkdOOo7QF7la98VjU6jHMNNHDDj23Fvhs3E6WuqMY0/338TAKBCg5w3sdtK5K
fQsHsgnpKRKgQTxFPcJ4jzfLX3bmbGoZVfNeDusoQgztS6GbpuSeSUB5bPYE5ETE
1peO53nxB76SfBRl9tx7UTebVdDW4Ecmy3vzagzHns6CNxDMUX2W8NWY93hEFcYx
VYnLLMTzC/XMbvVJGhWlEogiMi5aM9lwZehWP04ER+SmjBjMGviLkTyiompGj5jk
lEUTVIJxk1Lm1m4CL2K6t0TglwW3r/rNIFoTcjZrp1YLmK/E0YBDDaHvFUydhxlY
q+d0kroofuU52Lxup84VY8nNzcKRNG1womE6MP6iYDCjoUHB/jvAKdN3/aNb3hUL
4wvRNI9gEVLiBZfmsoTko/6n4MHWYCki9eezIFVToMT8nCJeAO2yK/GSX2qa55Ul
dEztNCiN4QBrhvSJNrOax9rXiey7J6O0VPeyoM0As3k+YVjecbh4yRMsVKZiiAGT
+Jnq4C3NcrvmiAmWf3DkJ9KITh5b65PjG8mvI5ZtM00uwqIpJEoB+7Tex7z1efMU
62wvqwGjwhx7LWYLXknnbxewuXCU043cQHiBQcbj9u/PvKCP0orRPGos5SQDelzf
X5DWVI77Mf/0tGDtEH2VRzaIZxGHtjKqKR5WL2teIojuQ2rjLH9Xa6PbgYIUqJwI
DTkoyZZaDudV/F/2AvftV49kOwKbEZnOOI3K8x1Alh131uEW5rgv+Pn1NWHqkx33
VWnLPhu3VQn7RR6ZL8A+RNmNMJIuv4iFgW8CrgP+L5gFNXZMGmBUxW9KX16+UPUb
aN3hwGkJ5oOcM8vQ6SiRAOWBbIZ12O+uUqQpcp813fy33sqQrP9Ask3CoCVX68Z4
Nyu3W87n2D2F2oc40cwecJFpHS21opKVAhMwSehGQvY/W7P3rlCfjsgrCcgKOevD
TI+0QxV9P03lxfgOFAS5s9fD0yly5bZob6KLspv4o8iGUeupXBDqCoiItGcAeCE9
rKv8x6WGPh6svNACN/w586pq5TZIPo6tScco7phT6MI4/6i7phtFunrulBGGGMr1
8xNgTcWwLtZqkeoUQTfOA3PYtJ+risRIaybcvdkB8fjMlXQl8iU4fxqo2zwSFF4M
xe4GylwTdT6Qaj3Ai7tfoFMfKK4KBTP0wXjD7BjsDmdToWTUAboFQnVs+nBHTScy
9j9JvsUBwQtVw70RO+1kBR6DN3qrkM5Kf72Km0N3g+abFz4/yUUP2KyNXVO4P8BK
g62KwD9VxzUoDiYmMd59xqgzMrt36GAc/z/AxbpR8sn6JwBVHzCo4GM5VN6UP/3s
HI8z3BdTZvufCtn1qQVTA+UpCkDlIRb3dmAiJJAmrK6slQ+7f7//3s0aOKnkPEhL
eIjI9/1HaiEWLrHHIsaCjGvRBGABVRVaETpnewi9OTCUfQz87C4GIB4RQPO4U67p
TWsisBmdnIza5OqSdzl7SdPyQgwN0kbVjfhsVlj/QhbFJ/HkfhpQpYTNxo2sjrJ9
mTCSSYGU+sXysVrxciaLXMh5grL985pL8DwEVHk80t2xg7590MSOWBRB42Q/sk9T
zIrKpU5R/JSRJzhDc/GMKgwX5eKvGMa4pDmBT04MiDwddIL0yBRhIKy9Q7foyl0A
byJede71r58To/7sUNz8sN7o45otyXBS7VHNDN+HaPXR+bkmMV+ci9Ha5f2C3L0f
T71WF5izDZIIcD31pa/Bz9ghQLhZc+fEeEATUd2AKZcyM+1vVCOX7zQh4DDumOM0
7FVzDiT2hD1yRq0hbA897y5REP6BfHKFr3tFzK/pZXZwlg/95ndxaITMgV52I9zT
r7DKqUFJ2182fs5k/bhUqVrmC/BVl00+qORzHalmJ8ViuMO7dEDNKhZkgh42D5nI
3SdS0uJVWQXXqGs1fmStHw0BS32miyOuWSwe4SaDUKRUPHzAkI4MYqvjV9Lbt1Wy
0g6yDg+UThkWk+IS66fl3h8Gtmt1j3WKg2DwhxB6IHRBBO/fZD7P6kKf0/dUb2yI
O11deeUS+I/7CE1/+J2yqzfqXRKvCZImo1noTFZHmmZj8zlIbi2NRhtCm+PVK1Ke
GJ3gmbrbMEDgwSRLCtZlwF8BamwIIfVIv0eRY6zC9Zq732/DZR3VZHX2s+P15LiX
w4Wq6yuRzEUjGxTFAbAksZYjzgAq6XvhK5DSsrY73y0nEI/Npi6/diUX08chCBQD
oa4ooJ1JpA+RcDv42ACPS/bTbjCZdgaJyWccOuuQdxLc0SbGaTEvLB8Fkw6oZIu4
X/v58sBrA07C2pdxXhug/QUnJrkXAGpQQ2Et+gu4I97wnIa/iQJyMCt5LhSDTKGS
6aKwC7jl0Okk9ADtaPaubQMSYKUT7k4LUznyc9sdigXUagc1ZYH6WsdHlvpida3b
UG7eR28wJ1B/JEbrW6VCDi7OGMjQqGMb0rnncoq3RD3TFBcKQOEZ9u8tPawQq/OJ
eqX3ALX/P5jt9jGhVuxCy27/wtDzdK90MOtm/3VOl1QEgift2eXTwn+GVL7aDkgE
e8yLyhLCw3vqJ5EdZcigUkIv2cR208+N7QbI9GX8X2cF0LxVpmpjZtnorUPNzMir
vAVvaVc0zIvcU9X0CU/IVgfRBc25NLBXvfLOePrhh/WydyOOAfPNT40G0gY7mE6p
Gh4qtLlkrOD7loSY0Ptee/39g10c4PeNwS5F4EiFiY6Emn4fqwU+J+a9x8IehXNR
uvttIZDuZ/ZL+HZgex8DyhHbaW8w0cJWmEjj5/QJIZt8SDEDWVaAUcgg6DqeOGFw
zg27uuYPcTSk7/bo2SYJPXAlVRsUeVtaOOdB+G66Nsf4qdS7LeTVcS0B9VK9xlZD
+NqdBFXjYCSiLFtxDcvON6aVoqhCYn1Zw7e+yx4V1eZ1AC1E9OWyp8kPIvjFa1zM
IcUbwfQRudmEu06+NfRYEh+TAbjnRo4hxqp2WIg4aMf2LRoTQPgWcS/tqTVfcK8J
EXK/hR1grGUf2OXorBEVdk8USmSZN+HiyBAxA5mtgURWwlQoUYMl82kObgWbyHad
PKngiBf/0J8KJuKPuDCyjq4msXkI+Qu1u8nF7kciXMKoRYrV7e4KnSLYcDmaArao
JAy4ixTpOeYye70eAD/x+InD3N98Zzd9P0AypKJxaCcWEU9qzzFWFwG7OW+VUgyj
BkzHvjZ7LH8H7nxCMEXkwWHUyUDd/ZFObsvuUoqsa/qNfK9aGcAhbLO5YKyLaxs5
CsRHR4sr1H20jTM/LHrGkh5VWyFEePa5u/e2KdruokWmzIBfkhm5s5OdELk63xLa
oCcxSpO7vBTQ2lld/HY9e0VHd9bg9HXJrZZ5gtUJIjZoPn29xbZ4PV3flWD4SoVV
VvcHYFg6OWyqA0eVGYR7ssG6TtRP1sp63H09rpushByAdKG8WdzwxIDXjF3gO9ok
1ditpIekrHJCDJsMviqF4PBP7SzG/4855no6lojsvCxS16Pj01kIbfgw0xUyya/j
IuiiaIHHlXG+M0hscmIGfBx5mLLOqR0Us72t80KhT4RJIxAi3cI14QJL/SfxDvwg
4SEnCP6JviCxZecp6dKnibe63JixdwXyyh+r28clvykInOmkxjtA7sVLDpH0k07u
ex+Ae8Wn1RaLPbnvQw0PwooSkPXx8AnUJH5wcg39wILQgocT/yxjgsE9mjwoowv4
KOxcWapyLvxvQhYQRwpFlZpoez47V2VbjTPU52LubR+RpK2hppSB1z++VT3hP889
vOFLglSXmsdd+zQVvEZvksc5XS0Ly4zparG1WWlGwuD6bqtnOxAOxH/iHn9YsneP
tXNYByCrQR+q/g68bo+GfDk6sAb7vOrW9NTbjRH/pVw6bV1t5WRg62Z7KdR6XvSa
NEKize6Hnksya/QoVF9z8yc3uEr1kDWGXQtuyyaqh9H0RKV6mioZ3jVDUxWgNxz/
dSYXasyRn7AayJfUp6I+BJajkF8ZUO0fT4kfbKZ56TBJyOLte+nUhSjHhSlzrAKc
ve0XG271pz5hSP0XQid8Asb4qOZ8OgP0IinqsvU8L4Ft6wGQ/AMM3+ikXl6qdhwJ
FwqQWj3MVuPnKcjBn57DRnyPUMvmbpH9H/xMCPtzGpApzbsUbGwVMi25ZaugEeu2
DLozburqorKpK+T0qdbyGVIW8g4cR57lmU7SrAgxSRmmN2ICPq8KOpuHRnIB5U2d
jEi3A4jybTE1QN1UjVcdhOujUdFWse5ZHqaWPhvyK+QU8XLiCCJd8WY37ZSwyRIt
b+Cvy3LiPvw1aYxg7f29gtlK+1WAPr+huyp9JZjlt5EuGDjgEhDoTAWcUch1g5if
WrTfMcTNgckWI4fcdXYepzbP6AWcbZIfNh1hms2tZEoL2vN8NaO4FOk1HuSwgfeL
noHwtch4T4HYHRkWKy4rose3eDAAbd/l4LIbVRSWQRDC0h2Hq3wjtLNovT9eXsSX
pdmoJ6UUOQAqUyI/Img2EGBtLzmiRSB45b/RXR4m9tvma1amSHNkPevPzqpMJAQk
VPbNw0scx8ALjQl4NxV8YIrS6qy73R7j73gkNxrMICe0rLoYSD+rEcLC/ab75Aw6
dlgqx1SwsVuq3qt+0fcfB7H3YzauJiLkXhYgElyxcUv2TcArCL+LqxQqt8Az0j1d
l4Iyx5j+b9qJ+Ec+tZbpIAdkIUD0GP2C5XU8KrIPJ7ZJGNRV6kiJtshv/IJq0MyI
bMl/fGQ5thVAlzi45HFnBrE9WrlEYnKsbNaXJD1TClzftRn7T2PXX0CsOpmzmREo
yiRhYgdpsgO9P2LHIcdAIZFi2/v+PVbwz3KIqo7ArJAXQ8xG2VfLbErlyd1kkSCI
OAP0lOpNgBZHdNcYW2fT/4k/sn43DbfDa9QTdbOsZ7ZEBCCact/l+gGURoUCxO0V
jxGDlDVRpVFJn8Ov8ra3MsWexpGH+dkHrh+KOLLxhNuomGi7y9Oiy+lMnywDuIdn
MxkWkaclTbxAqSQUhftYhiiqw1szpGlXGWrG8snpWCyC8VrPVpiLD0568YX4nNAG
TSTf4CxVYQAmaDEYhYQzj08Me0itqcKKZnkP7r+iTuY6dAlHWi4fWUCEG/fiuIIW
1Dcv0HvVQIswOnM+ZW55Ls4dZpQscD8n8dsO6JNJLmMJxQI5MjSWcl4hdIE8kFEf
Q4gQYfjG81qYGqdZ/jL6n09rXyPKR8tCk4zlstMPtcUwnZktcecBKboscgTUC9CG
/RllEXbS0JywjLYggmIZECtMN3L7c5DxBwk/G4fT7vWETdyAQsWlrlmq9c0tFvJR
zC7Ky9gJox4vuBbF+JrmvqQy7L0f3QqmBbUNFQLUpe2nh1S3SRRn3Cqq0xQe2JK6
MruUh+dOsZj2kD069FVfT+bdw2/UsuQHyS9qrx+8nQfaWZNiw0GayT4zG/jxJIeU
N9xkTX7MA0MgETZSpjj3syS7WQK8m/Ya9lzSCHrvbCjmCmL9ciKUeSjPbrJsXZ4E
L1oSw8mBc2cHp7m276AAOiEDDaQQJRjnpsKwzbz4tYQ/dO5RjKfrPCvocttY6Zs/
+Uz2CmlD5t8fkL/LgEjhRwfQrBVcxf9FJn5nJs6BN97mB5xOiMn/n4NzdmXjjLP+
FuoFQrYBnAGejk39jRCYzJQKBlU8je+MR1YLPPhW6mZvVorCXMXTfVRjh4wPeU79
+014s5AqedNyDL4zu3R0bPnrBnV0ylHhhoiEmnBgbfBwE++KkZNSWPQB9Os3satW
ooumkn0cgtmBLhN172E7QgnEjWP86kh2ceH28lztCSWvxipj/ZrNqqyK3CY52MAB
FwkzbvWRKTya2uJXlLA+CPyXGYo4YJECDBWaEmCTaUMl3/WzmxkVLsl6TPH+9e0+
p8elh2fKkjk+fp8+5vQxZ5KlLhddc5AcuMhiLXtealVZDeRIblvScVY7MTboP7Fj
iQDNSCfRn8drfc5iYATQ/u63H9JKZEnzxgO0atFd214JBjq/oHtDc7ip1bob9UR5
xhEHGSvP59eMb2Q1/n0bGqC+fAyQn9GzOIZFVrffVvgaNw0D89oV91KCMHf+hXIx
AcoK2eJkLdekv44hVZTbfxEWbzBC6kr4yqEiC/wVAi8RlXJdfvktO2rxX7zx6lDZ
CyqEV3dDSK86eXyB9cKfzS5FbXhL+0f+gZcA6GmsN/sYsfqBmQxC+r5BGXotL5Zj
zkssS52LP6SxVznRHGT0FesSECYxln4PwOojcAvxPhTANo8l+EWYvZXX7003QepE
/YxWk04DHLj4akQ5+R5GN8ulUGafbM2kB5Tth8mOju3ghpg+nC2a4DVtTYt03XmG
6PbW+Esb8UcnIfI6+LTMcLYqWx6o9eAMN9sv5CR2g29u53DtJEDnLnwpVTY7Azbo
TfrVyDEa2mK9BATFe5x70r3jBQZ51wsu2tNXMKMNKHNHPBhoG5xFAumzBeg0WJKy
suCCXoD6ZKs+c/fATpq77oTvQ3y2sFfP2Hgi3i9u8bDrVzrolM103Tq/a5cDcHD3
Xt2mYn+tmEVw7UdfDn0TANpai97hsDnlL1lYrh1qWzyh8c8ez99sjCqJtREWCg70
Rl9S1ia0ZYEreaZRQ+r8kwv7Dd5fu5ZVarexwjP/2Yv/66UdEwHuf0X4vBm1e5uo
c7Z6scQpZPOgbIGMuvgLgnKumbCYbzjTiN4zCkYg/3j1tU0ray+zcC6pwzizhqQe
QWBILh49DDQBOyYqzQD02BYQoGxQ/0ZHpWMFDrqhAUAcc/IxYxWvtrDQQpTrSmJG
1t/ACw28DAHH2J81Wm+gnvb03+/zorPiVXXQpPA/v7bY9U57cq9EOHi7vMRMUiBy
GElJ94rhuywCxm6t6ZsTMLtYeEAYASJPINifaT4NsLXmaTXGPVU0ecooZ20ktN0c
HxrSpRXuSrdg+N4i0gwFvqb1NPTJlKW059Y3iB1g0BlIjJvG6q5b9+V30B/i8BKr
GxQglDVzo+GOp9g9xsg7OHZROChuDmpdcp0jsEYUMLtu5t0jVBCX5ve6U+lVxz7r
FarInXL7ybHAdyqFZGPmpl2IL+nxGfDevY0BSwd2OalE7G95I/1KWlkSJ+fOzZ6D
tu4/nMihwP7IPUDD31PLh0nqvHluJj2R/j5M2E2jzBoWddbuTTTohXgbU4Fy1Z2F
bO4VuBM3irpwCt+AaukJVsXWqXBDUNmmG2QaCvD2NMlBHu2zBg02ai0IqZV48NbZ
emTajARhyhyGh2sQLcjJ3Y5rLFDzDX9COMfwD8HTv43BXHbDn/mM0G0CO2rReoox
6tunbYVGFVCVOWBs/yWoDZJ4Xa23oKZfvsB+PgmPkDBoAyrLptFq9nS3CgTTUBwZ
yK6vr3LYWjP8/ABprGKIGJBdzSJ5fHFsF/zKgGqWspjWkyM8U5Q5SvAmgJ+NvtS8
lpfpPZVC1xUauHx9eIKe8dKcaAqeLpaWdl1MsQDCMgaHOktOUvyFzN7cCEQX78qW
mtA3kzRhnPHudSTxbOtw5ZibRpBHLsvgXsYKumFBe0p/QIoUwSUg6tlerzfDxNS+
/6T+T/YsH7NnUWM+dR6r4ExT3/qoQkmq9N+V9dU/UStO9uXgFGR8Ru7vAHCMN4ug
Nd2LHXTwk1R8WqALL6z+1JMxRHAhTKIxZtAAsb0Rhjrc5yepI2Tgoo5WDFSiUBMg
xvdf9CGLVLZ/Y0efRmkkFBRriN9ANFEj543FoXb4BCaInJb6BZ0+cQG8PZir2HZQ
C/2+Jfg2ucACH6oivrnAbbBiJjstrApNIeTa/hAU18CKEnZuvZq0HgZIjkjNP7um
WcMC5D5qFtyveFmSPYuUqY0GrbF8NpPL89ne3yq9IUxoMTuvqXqFGs5FcmK/Jf7M
GKZG+fac/8ynIXyROXymEHJOS8Rp0fjXMa8HChg4FSdVzfO/OcwgSc1sOwPuKjq5
naTCNkPtekJBRglyQc/l2ypSC0wb2Zrhwho8vvw2XvpL/JJULqppZAHBWUdQT6pU
HnS0vxl7jViSGFhbcqsq9mEHzP20miaNsaGUZlxlIjCMUvnGd8OKu5Ul+UnbueQS
OmC8CPEUWqCz7GWBn+m81hUEqQY2MjwpNcJf9Ce5ntArm8vS0i5OCh7KvESBapFE
sZHCj+aR4FrUScY7G6FhPLNxKkV5FUpvvzKdFxY7MSiMFnqaXRpI+/yNhZPXUHpd
OMHLh8yGV4ugDRCETXx9RkOqvNz38oPBN4boAOg9412XXWHshU7tYmkWeFTv0UC/
H+ed6mO30bgYtrcyy482ufUZDq1qCFrUC2gaMDMJWv/4RtrA0kBHvzEmtHz6TrQ2
Hh/EOCyJ3ib+MzOdwFFnOxbo3Mjh9sqfnRClgY/Vp2ZkIlXUnAD+14cMX7MHAp+N
iMnS96nqX8lcTdQ+objoUPyjkh2dRWxT+WMOvcGjqUZvebkuGseRfb3MNkGzvykg
4R+DrPdtWrqRYka6OQ/43tNrKoqCwyBa5VB1O730nxxMJalXYr1C57CjBi/x6csd
Z+PS4r0IdWT+6dyrilH03RLbM9eIIeGcvVgV9kae8iExdXBUBGaCOTQUBa0/1rOF
zHCcL/Xp09o/9jugmaSccohclbuOqXttpTzWa7g+HHUDNqXQeovrqSoPJMkJSrXC
ZIY3SZ/XwIh3ZhZCbVuyvZaVpeLc0NSKBo+0Z6jGPuszb98MkmFu6npHnGMnlzrX
CduAzyM3hmJcN3WWF7eRxGcbCeFy8l2qPN6bO8dHDl39QGgM54h+m+1MaoH6H6TK
3FZYi/qsmOLBcyRDJ7d2g+G476n1CNGirPU/AJP46MNtlUWnBlTDMWtgxqErNUFh
s49pF7FuBD8BKZSIB1dS5vZM+OuV/3y6T2KBAfQjax04/kNi7I9oI32MqdqyUHqm
S6uZx+Nai85qna6EE893sO6Zcar1bDlqO/JwOj1tOaLGxZN9PbL+tyWlllp2MlqO
46m7L5hJe7K7JyHkiNsbcR2N/YpuMVeoQI07ooVuMvfLsfcYdt45WIt9XBgqwpoC
gDBPKU1/1IuIKV0j9iZFWL2lbhFNQcjn+y/gnBhZcDG+Gjs2DYlfMrOty1ABvzTI
sUswURGa/MUEtWdVIjYuSVaEsAg2sCAHWOoV1bjx5pkferN0BShhAT59fP7zK/Wz
BykPDwYp/trE3FaTp6crZyENuECF8Ry4ZPGFaMG9+VKNSWy3eNXZsDh8XN7Nz71c
xUH5E2OQ3JMsBKwPjp1+AESUOceeFpJT8QNfYu7635b5BBHvl6ZtGwzi0nrokDTE
D6dpi7DJc+wnXrLmqC89p1JmjQ0obnREiYtdGreWg/oPvoXVscCq/X9IEaymRo6A
aounLaU2wOcADWd/roCPNfH1AurfHBy05vfU34qRTDFBrKW7lngLqTEwHn/Z0gFL
3zQkXbkHbCsbUfQKwtunQVkdDvde/d5QcnZt9JlE6716as3vN8M9VDB5umV7mjkd
lkZzD2Pr5jyiiaOG/UZDMEkKOzX2GD86F16yG5BaIR3HZtKq93b/P7f1/NoJVIXl
sac27A6LJ5Q7O5htOvhHpa+tp1tfNewQp0upAy4jopRlJI1h/IzFbP5GKhbdIsEN
m6x6JfaDgQeN5EV2fMtU+sY/XHOOyKEisc6L5HAWvv37mYp0A/XGdo8LRd4LWVpW
8bQIN2CUPBETQemudIDl106UuUHAI8g0SXHtED2UGJbMfCRZOj0znYEWgLYBtsOH
IwIZz7UP0OqTIkOTWE+wPP+54FeZeGgzul2o/d63vAIG4JpIsY5BOwgfipt7p4ML
GA0yy7wVzugnyvrtfGSbeE9JY63SN+dQtlIZxRZIT2/w7k6qLmyWV/6VuPPDROyv
IWiU3zfxjURwXhwrU0/opEUr8BKL369q0o9YvBptqTkNkmGxU2cvpVkYJnNJrDpj
Yu8wlFx77j4qFSBsxTPhuHPIljwCQC+MHVMXADnUub2CWFb4XGe38F6dyUGPPhgZ
nQS+MV16oXtUkVo7x6/vN7+8FlNWPHvlQQLDAznj2CB56dOMi0y/Gj5+C97FSxZ8
EDsSifKJiZ2XdPx7NK/kDoUuZHglBrWGuv7nUWznKhPWgU7TorgnVB37DkQ7ABXp
fKxy+vnqnyWZ+YN66rlXZiOOR17FplWHoU9t0/dMXESqOfxaFC1vIG6MorHk+7ie
dIGk9cNosQiKrYHzev7srVd5ZO0sqaCpdpzUqRxAX1MzSw4ejnldiRzLn+S0nOx7
ftYUZ4wa3gt7r2BHyyPTAn9XQU4W/qCWzsSEefR03z5qCLF1+FgobCMuX2rJZ16Y
g6aLw2mw4LgAlcqvVCTw/ohY54LXt+kGz70xluHaMYqFRFzN70vfKW5Eax6xb4dY
GMOilxHRxxYgXBPZ2ltp1wBN69XXwGwQOaR7DhzvCpgP1zKNTEPdR6oNCSznwyrK
d2CxjjtUNcWLif6EWOvD7ga6OcA85X0PTQUOG/ZgQWUQq2Y+TMV9NF6qyYNVWYee
7lbsbjvPBaB6HJ2BamCUXzT2dilwUDsldtVR1TSDBfAGnWF0pR5QuaI5MlFvz8cC
cB2U70q2k4b6KAixjlMroozDObe86GkVjdazL/xGCoiHZDqnPykKy1wFcncu3J59
XbxBsiq1QSBXgI9P3Ho0aBzv2Yg+w8gu3UJtG3epKwz0kXa5SzxMl84M/r92xAsY
B5JFogb07l21JfCGfhVGsHHX0Oe/i2gEKrUlvPdm2r/RD0IN8mjuvLWZivjMVUac
Ko9t4hM1cbEvl1IIE6X9np5Gd8OAb06eEh6TxNFhVYfyGG5wNZNPpX3mXLHtRKCn
735tmcBQDZCy93bN0Tlldw2PPdGCx2ScC9qeAylrkIibtRAaD23QED8xsgy6KmTH
F5l+eHYM/4zeBLSj7IiuL+LJ91PO4tefJpCLuy2SRynwyJSWBQO3YxZd7fqqTyzC
mV7kVOGQ+QNRCMZZEm53HsVJB5IdcgmgJS20ILAKpkg5ZNe5+HvtPBQi5jF5Ktqm
21ZClAgWhmJ9Kgw1bYZAIWd6TyGkqxrRbkN+0tWzIMrR5YeThSC0Duqx22h2EVdI
gTeJ3gkZHc6LrDluRrh82zUrsgESNb5h4AQR2dmSgOPlYSIirLaXCw1zaHGbxMK7
C5/6WzhhKHda1YWAUtIE+t1j1jbZ8EQtZgSm5eS0X03ctKPttZDqQLxVo5aksGkS
c2wW28FCGrjnXgCpF4twjZ28YBPlQ7ScHkaWfeFOsriyoaG5ejnI8cikiv7Ig3wq
7SMMvk60flX9GmA9MoboNQ4LNW/erzxFNT83IMtOCQnhd6rauSx6Lw4Ls6CwM1nH
0oF6X2GuFEq/1Qj2/E+Cfdsf/7574VL+HTNtR/79GVtcu8ied4caMIi/CxCPYvpQ
k5y7UJ82fQcRUB3tV/Jq/dCyAhsYWop3Bb39iuEZ6f9myJNECItOYuzUJBZ8MH4t
31SVc/7euHqYnGr564aLQk40vqZ+12jy8Bb8enwC45FwlCyvHYe+VKXs2UPGhSGN
aISY3t6C0SJSGQeDtxz28nvYPtZPo2nNCm9cquqLlIBxhDCdfPsnlkcwb/VsgwIq
7KByD6lNsbnVA3UasOVycTp9euj2YTVMdnyyt7Jm+r0GnKbN3p6moS+n9dGKSPe8
o7wDEkWHKJIlq2t0w2Qe0+V22D0hWLOYHQZkyOwEIIacEBXoxWiHKqveQMoVr6cc
a9KIuyrLEmIgBqYV9ZY2yJIrOc82DyHCJWCZPJg1z9X5kYYkAPiEz5H1COyuJfN3
0Md/EjpH/FqcWwZFZNg2J6/D421j/LhyB5jeNv6g8L2VcRKZi9OPzyPv0rDoLf1k
Mr3lGbF5SngVcqV5L26aXCl3MR9kqTMnTOFifmuNcl36pXeSmQ8tww3/Gx+ammPf
0bmcdAhkKcLdvjqnR+XwxPDpla2qjnkFTZ3g7LkFaLIHXD/z01LWW/hHY6AHeSBf
JjHRoHWzyK5DLSVaSeT/Jwyi45qGnELyXQa8awzkWeBZG3pGXS0uGdPoL2jBHtSY
YiLwsm/FtO2N35oKX71aUoKSfIfBAtU7M4LzNAaBCIYHQYMMBJDlz7oTxzSJPRjG
pn/m2/G1Xy7CLpD2bJtWeQY90EA9dJVFLk75sjwOi+VaQwCGPMJcT3nTz8vtf8xd
1HzmCHH3eBoSpIn9a0SyYDf9dqhx8lJ6RvLprwEpP6ykP4nCMPuRNU3OG+wdgyHH
kiJ0KqnltGrvjM26ABjabZhF3NN0WWfgueP/L3MGapIKkWFVRnyS+jBDtvt7he6I
WXambcgl6GY7qaf+nQBQHZvANPtGu848okMOdN4EkZoCK4jl0WJ6bEIH8G/5UsTZ
gTyJF2IbcHw+BgxOGTymPOZguKWNPgPtABF8SFDfRAJnEvaVm4VW6ZzwmKzfrdRw
khPrUvdy8X/b9KCTmiN0UpKbco3zh5BoenX7+SmtFDkgT6rl332SISmo1AJGjfZb
/C6jDbbSHYGmypLBJ+CleVStTUHFtnJZ0Lh3Nr0aKKW0AWqsqOdWsBG1AfjqMkkm
C0/axptzNaH1y9zK6DV5CWcK8Ap7x0Y4YxEMvM2igT7i27gwnB1hUbR8IaAlRhN+
oV1boIHiTHt7vHX1ZuLWLGg8w00OPhZpxWPhH+XYmNgfQJ+vVnq4c29akxZcYz34
c7/AAq2yaQqPjkTZAIP3L7O6XeFEjGw8+bN+cDyGeOEzFvixqR+Oo9QuaUjWGQU8
BeFNMkHIGZxcZCMhVSnYVaURZw4ENHvIcTaciKPMIEd27IJnG3q4AtSzCTP35Nfs
2Yys7Q6+rKztrHNgllO8QL4OcHuNz3mMYhHxRrJGEsi9M778zyY4X+rBCR+PuRgk
gnFD1NZp3s876lpC2hhEHsHsPMbaFEzIIkFktZ3s8RlKJ/hEbRWl6KTLSY7mWnRC
NQMjQih01HRbLPQf4QluOAGuSem21nsmzNpPDBxH42PuV/iuc5tXiRIYgufTdTjv
5V/dzyWMwW354PgdbMwFqivNoXy+L/EaiNs26Wi4LUbe+IgEQpKUTJYRQK0Ftzuj
mMEmE1zSCg0Uu7LMfPGh8Dz3PtvDI0t9wtX2bKgbluxLLXBTHBelfCZdJ6BTKw9R
sDeXWIFdprnno0VvwzQ/8BW7QQ11yJ/CE9dzNX1MhghVGwT3kt+vgtlOg85QPYmA
4q3j1jjCcEH7yYwxp/pCG/xUEs/NqU3GUnTSyvoDgIvIouYP7aa/4234igQ/hxn5
n/ozaWtz3KtRFbUDjH3khkZChPbdWOiuIkm5lIuicopDS26Qg1bsrrdkmheQB8os
Ialt+lucNUfzZ6BwMEd2WPbxCVSIiDC3lTAutW8POt7XM8vOD20IPGMEUJEP/SAW
NaqR1cKZbQiowGmtfGpbZKvVMg7RyXoyZzdfUE5BJ9PGRKEa4A1W4fk6XIxxAOlr
6q4MSOYR/SF1XS6o5RldCkARdtxNxYXBVe5CuJz9aKwgMxza5o5mvWn4Eb11xL/7
1Hjl5vMxwkupLER97cxeGBw4eJy9cCXCdrEiLh9LOfLbU+yr/qKHkM8mQdhUCKFH
WbTsTub06gJmXh7WxAMUCvd7ZdEvEi1T0FIf8GU4MIfLhrf7I86VtHmdjq/k/YRA
QM0zyERLR61HwNEfxec79dbh5/UNNFlBCHSo8Nlp9lUwKydHUIiOMlvLOfds36XK
yyUd9VtOTJEbO8H9feLXycT3kUhYoRVBYvU9CvAZAEozu/pJHDU2tT0cydeSoTFg
+5MYtNl8PjTITC7Zp/BpOeQOm3l5pcbll9674lA6n1m9Xx02oZf3ZNP9wRbyJ5fk
Alp/sn8EoN5umja7auOG9rFQAb8bNoTN/vTCI2CmJerMawrNiozDrolnSgm8lDBT
33sCJtpe2nEUU4W74bi6Kkf26UG/zqOb+zud5HyGUhYUXi012GfdV/jEIjUDfwwr
XBMB5+MmWbm9QHZlpmw4VAduWPfK0UzCN9kUNvpZcl4qnrh2SB1HqWBVFPC8R0QA
gVbuxCbfyZzeiUBFNpcC5uTvrU3MK3W6SgzbXFDo0rPch2ZHV8UKsCeKrMCMn9Up
lpjdEHhXQTvO26134oEpZTrntHSnecl0rQgVXxelPGfWohAUVHQKyXY9C1boxdhD
IYrKGFG7Gtg2vJN0oXC0T1comKD4xNVWjzlSHMScpUYXLeKLmbR9myDkRAlUE2X8
qd1FxKW6DIteWg0raBsSknGSJ7vyOx0mKh1OmO/xc08fw3cTLq8ALdhqRTAOnK/t
o5bdBzUHabb1XLLzVUNtM7wakVi5Txlxwz1yrGeAcW6AY78QDoFJB+HzgxAQp3Et
lKpCEnh2hZERBp4GPgy4sgmnVB2cY2BH2R9JCX3ozUVxGBk9X7sPusyA1L/beaLW
Oa0VgM/hCOxMNj93ZhUB0/YsaqE8Atd9yuoH/iH71V+TNlzIToqcKjW261ne5r5Z
t+H31FpO3+lznRaespMx/5lPPf6a3Fj26ftZA9kCnQmH6aGvAF8H/u6mm80vSG/X
Yvq5Y8k1C/fSgZPeiMk5sms4lhV5wlEOddvkd8kzhgEoRMucBP4zDILreoFNJheH
Iyn29Viuy5KpAAIaT2GEVg/63I4bYPTAEeLvPsJa2IDbrfIeYbpHYkl0Fj4A1db1
T9osaM41bJkoMNlk8pnzuZO+oPDx9l0OPMp7AQRY+h5BCiX5Jo+6ACnZ+uk6tXKn
zsQjF7ekKOaZmUNHO5wgUoCUJRwd6ctoxzF9OYuR+EJGAfQCHZCK6cnwCvrtr3P4
MtZlUTiKoVDjz8hhX1VRXd0n9agXjtTP9zoYReBlNOmGn4KSJLrLurWNcESJIGDp
+aHbsBaCOK/RtQwj+WEncvt+U0GhKORg+oMg5tPRtfFc6qG9jcUFnL8Kfalv/jvA
jKjbY1XepuAggQtM2w8Y2Ifn6dMTvBfeabdwoCs2h2hwvCfmodecbHWAiIEW+6FN
nr6/nPSXiRc7YbHEJwa9ly9LXuGfbBOvDZ/O4jfz0xzvzyILKifZ6JOgbo/vEtmW
sa0++N5xlhlcjv2LBrLfpd0UK9OoOpNW1cZWaKnoo2eMCLuoA241yvvJ19i2lDQJ
dQz9Lx7uASr+6kzNYNSHyM4R9JRw/b0h03uykzntdYmOeLozryZQsqHUM9buA2ko
TA803f2oEH2+ujw2/QrAabDFL0/a5PMLyknRZqeIgtYtwpV6Jvbf91Tl4tVlH0Qk
R70S9Z5tUoo3wi/lLrAMWAUHAs2Otl1mzaitoXC/qjc/SnI95r3GwPGo1raQk21+
4gF3tH3yh/DWols1Xck096K8p1vQDkHGBcJ8ztJGkPug9LiKABuiJButxlKoLjig
TxVx9EgpxXaebmj1mbWtUhHIdDLnc5ypZNLVGO/2T+YnMHOhu7hY5/oOq0+E5tud
Yi5sI1AvUHwm80gdjVreblEE1cB2YXOGrujmOxTRUXvB+4rXblsVuBtBQxnzPjDC
fcAR3l5l1V7IntuokEuLV6e2Hk6afx2SbByi6vpPRKo9LcSMAgofF690H+mYW2cF
fDGYHfD92lMhjW3CjXklnC38/fVHoegst/LlgqpkDcyaGGHGs6lKkthsq+JM5wRU
6oPhwOmwetv2+DULDiKuFeE9UsFr+AOh2JaWFNbQiXKrbcBf/6MHId2STV6gFS0m
dQRM8HC+uamzKxTZ94n5gWDAvpiHKfID0WVkF/qO97Cd8ZvWrpFqmPxO++LEtWgg
Q0AYMTcE9F4gOc7W8GVxbRkM9nrPj8rfEs4j5amy3YNFPqKF4rJExnyKa76iHTon
s5ljOKmva8imn9MGPJYi4zhfTSYthd71egut83z3mOtQyLY67J/Yc8HbKFDB2vTN
tSKtHkzufr6eqrCCbOQtdBn5z3V3BMTZYylmR/nrKWo//hOMqP/uexOPdM9mBoNf
svXVK+6ZrexQ0LOiLJI8hZewarAsXkIVuOjCVWnvWQbD9esNYN0BGJAO/NwBRfQa
HVxKxeEeDEKen5QyPI8v7zTADmIaKma797o5ANqXCueib0+/Tadve+NQ1VCcmBki
foY0iXTSxz9OGNZN/4KZjdlDU8kFiW/f1rWg3+7hgvbrSgs7ovXOsvhCwe9C+mq8
Meja+aQkdrc28kumKW7X2m3tN+M6sMG9+HRytoCGAWyJLpJ15MW3rwjwvvZanwyU
YW3Z4l37Kd8xD4TpeQ7KATwuFbQjpmoUIsFx4brVNmSD8t3Rrt8DVTS31XRWBok4
brFpoO+pGMo81Vep0a0Ddl190pY6p8nKN8HXpmJvvsZDMzhz1qrnNDK25PdgvgDj
3h2PBhR0YE8kRir06n24Io1Vx0pkmk8LP/E4Q9IPZv87nWI2bl3/0ZxB8hLLyhQz
FMjCyD11GxQkEf5lXLQMaZ31t0f0/74kmVnGmtdsZshEkc2d939A/Xeo8jbDB/Z+
f4Q+lm3k9qkFMtM8306esaJcyJvZb0hSSJ686A5C4xGBdlxrFyHL23I1xr2umORZ
vp834BwxDqEiGkqFCHTchExiry8UAaCF8yblQS9TE8bRjMFaGc5vaQWC+w9epgtL
NN47dPyVY/p8A4rlOXzbdHsn/knE8vLDpC4Nio+D7fUzKlX1BOkWUju6px0+s0+Z
nMrjBAmhI7pmVHxC1KjNs2aSdnJAzIkYt9GLueNsi44K8stdGolqsNVN4C4+F2vJ
IPaNredAxeajXS4S4OVnaFPLy9sB/V8HFfnk/IhMLjwdxsQSbnSFGM5iKCZex5lt
6saOkKcnMUI/cL2akaM4pd7Ks5bX7Oh3c5rJtzwgaIkZUYuStXhSQkOiMYK+cIQ2
Y3N0c3pTHVSGB4WpLbut6Z4gAzURzeXUQFIazvBcHw6ibkmmDJQ6NSZnAWWTHrW3
ufXHwn+emMvbZFz6UrOzRM+jNhc6B1D0NLBJ+7y5I+J6IMYPV0pzbOfM/aqVXv06
rEsXwVFt6YaiiGQs12r8johkWJs6uS8DB2VuanCbswb4Rc7B6TLGdYdajHRbT8RK
RvLBQhM5C4og6km2egrBJFPPehRRuhGl3zm9U9/wWAuZvHbcD+VNW/UlY6u4LlcT
pEs1YGbB0bZMOTYh3Z83A0yIO/ixR9/A9abnhL3+ZeBvjY2y+RaiX1/lzShpCSlw
yaEJTnQ7gGdhuhqqjOBs2sgkVkcXKWB7Ll4RGD/BuYyDX+eXh9SQw3Jy2xWfMTer
KH/BB4QuFyp5G7w6r8mDk73C9U3m/cBOf/DX3mIuJ+FuT23v1YIFWL5IeclvmEr0
1QRhMx/54AUr8dChmDUh+8/VJ5LELzm96S/ob8eq7HRkByEZaW6iuo4/zuGMxlsR
QNOLlvwm1aQYIrToRZm1rmU8gh0irfU/YtfuE/jpV+P195fc3FA0V29HZnzcxIRS
H9PHut677Jo79l/2IUc5sw4mkWCmfg3lVL3UhQequ2JIF5egvztaoZbHmPZQ03/B
1cO8dduLYjDZ6cCNvLLBwFU3PDsBP9aoKVITA5sxnaSD8TRFihVZi4AefmQWGjvF
2ptTZLHbogfGtr16DT0an7n05frZJM9WOdAwKfZH++v2JcBByWbWvoXV0b6IMt5N
/nvSc95FYNfDcZkdSn5hCBRzNADgERn4GQ0oYC1pDGWnbwHTstbFIqwQGVtZ0Y+7
kAcJpQQx6P07jnP/hGAL5EY3IRYdrALGwzjE+NVmRk44Jm7usywG1FbRyPDAEGuu
wQVGWhBZM5PocTPMpfNDqTrUshWTXTKCKld+m+m6s7PRW/5yA1A7/etVIK8PFI+x
dtkDJtEDvCbM1rbDod7q/z1oMrNJPnOlRCJXDJhlb0Vq3cKPFoz5juosiBEvXvWE
7kzqJ1UW0MlBvbSJl46rdOsgjXKMh9CywCcYfenmaGhxoPxYZQFkDH+seKLV2hQx
ZyIF6AJWQVhwsWEQAmgoPTjcXgTG+AC7hzIV+66+sMBbEflVhqBoAOTO24dgZgT5
kIaaQUI93PeyiTEaHotRCuuWwqFX75e3Og+lz63UuzwNSN8e2Bi8hJz6m/WlRlvJ
88isjb6toAfy9Da9QmglYPALFVG6/TcyQG6u0+XpH9EoKHx3ZtHXfS9L4aL8bB9c
+Y6yIrMMc3wVVaI9Wcw2HQ89y5VSYx9Loumx9wRbWmzoE+lN5CTJaMxqZKB3fpUL
e/Vd7OlTXwnv26CIsoNI7aV1fbsS8P86UgxkZS/LZQ1RffSr43ypxqBSUptaSJ6r
dmL2eItj37w3miry9saIlxXPbqVUlnXThBlsYErh+m06uA5VHpOYhjqma6pSnCqU
2wxkNW0Cf+LDzahOSXhyJh3kDpFWQafqDtUrWhldNh3LbK15JfjHfhVZjinkDXrR
L+eHhUJhciULuaHbr170XMzByhdyf7eg0HHogzCwHm0CPIhGSe071QhVjKWQE1oG
ziU95eZ3ZajDEKUFCBqFa2jtxSjRG1nqCeIMNasNTSq+zm3uDUrxVq3EiM9TzJNW
DX3A87pYg0IBUK1DXSF67/wtfdqulA8kBA4PYcDZ4QiWh243x92ufi2tqbASb9Sd
oViv+0ZXP24HtLXrTYFzNiTsabrslptWnEyUZAkSuYuFsnF3tjqJ+uV/4xAABtkq
bdXMYh0n/Q8j+SoqTJkJlYtF0kYhqKz3wsf47kOwiYBGqqXX0wFa6MLRll9Z2xGF
gsZSJxuUq6W9T6JC3wSqZhd/L7rU+AaWFxBau4fL33HCprzDd2l4cYNJ3ZEmj7tU
vVcznpynnB0rmzaWIkxH9ryiIdT7PNF9aMad5hi3Je5ayyXgbVMBUTkH9G95b+b/
FtsV3pFSPv4z2yhzXtJEyq1c93o3NEWFojIjFMedsnIrgYjqphbusZs0EBDUeRaw
IvvSFHzlQCIl1Jc3FY7kx7GEfo93PzGCI+f4S3sTo8mvefxNVzbZqZDMYcpFV6ZJ
vA3ioqw4jIZjpRK5S3PrSalAWs7+5bm3cbI+GTy+K4cS2JdhO6NBTXkPodYGD1IX
1ulmG5ZlYR1fgABbDa3jNtFkJAzEma/stWpcuHG6XZ1e68jvfUmS0dx8pdIiaKPp
LD14fatvzl48YJ6xJgqDI8wsKJOWRbE/gvgM4kcjbbitReQwFVr84+v8MIKLuJeV
7Yo03E35b666hBKjoPz6axIkJZyvFCPNSBeAzN/8drF8SZqG4GquXegRw2sjxwwi
bjLClmJ6CAF4MkjoYtDhaRD1cZprW2P6sRtN3SPeJeDzMpjFHrwcQufJMqO/XjA3
NL1u5FbJP6nfyeddlKFhlug0u/cMEBMpaYwCeI8sUC1eAabCaZkVLCJE01xXR7f+
y9rJx5+0O1okeiDwzcvCCJi1Cj8bnNWRcTyps26OCtND1CWcxEW/TF836UF2j+lG
w5RoOoZ7p5MhHIhvs4ygtYMvDMa923Q63gI0hFVXH+h6n9MQWw5kxzIdzVk7j1Pl
y0zJL3Vms0f1RZuLa6HPxn/JOIY8aDi6DhZlUZ0m1vqEMYyY4kigEL6FVl7fwdvl
dS3/dLgFWql6yyDPI3bsaddJ/G3hPL4KHmsgSVEKyLR48Kl91lpaM8M3yFrEDBOA
6CIJnzxM5C9iT7+iISUnb8lD3xH3/x1EuXhkByUIgyFfsWeNaAda5oTCbXdXswuI
+bF5mOa3tRiiSlwfSJcIu6P4Wl9FrbvrLMHUeCdN+RnXsxIt6PfyeYf+59zKK6oS
lmBIgbZLkCx9WQu2qJ146scVZ4sFqAKnAEgVqZAAykS6JW+sUlHZ9Nd1s+nthxze
GqGMBJ61+2pzAhUjI0WeqhKT/rP7hrQLV3Ah7rDpTXbqqw16rOxsjzNT+F4dXA32
sdb60Oe0rOgSNvaUb30iN3+yC92+Byol9breVGe47VMQGVd0rgaD00Upj8lVlDkE
/5rLM3Zf5APXD8/n+ZX7dJ2ivJMtaumQ/WjmnWrTB6YjSXMLWw0bxaDW95uoZVFb
22Yoln9GjIJM3xF9G5PtFkJbEfmlGioka/fc9bMba6capY4+A/vYbLD4A/cW8lc+
2m/0kurPuCV2CYPIFH6CB2q6N+LtkB/Yved3BDvohRBDRTJDGP/ssxwj11yC3fl+
2OnYH9tUWZkbSjHyhNLDWPHPXBY4baL1ZJpwIDxjBHe+vcHlAzKr7UY5n8EBC8OP
z6MqP5bLcci0xU++IA9RJgrpxL3VQ8+JX5bCuk9nvT7R370ccceOJJpgXkPtvI4F
uO73nBXr+iMcAKp4rQoNjPXUbYUn4NeEBOOVin1G/Xn158jbcTgNFMZ9pxmTvCDK
NH8QQbKtCSbbyEWqftb3jhVTeFLiZwgLJP//05WmO2OLzJgBXmfyjNqCOyhh2v/G
yZr8+rtxZ9drXbwb7HutJ02DeSNRSLVNEaGGHIc1T+dktIN5T8nqe6y5N76xh9DW
nzXFCNRgmlvo/wHp/2DBM9zx8nK4SsF8QqVm/dVpnULCrixhqsno57dCZb7f/Vw+
wYH0vfA8c0zPAyKBtW39AXjGKlgKuDRL+/4m4ZTbc/qqv1xtaio0/d3CbU+zPsGP
UQzLEUQ5U3Mu8whCrQXv25XsrHAZgRwFNCR6RCbgGtGZcF3PWNUand9ZmlpeJR65
A96BMU9ZDZfpWDyUIYLCf+vdUyhu1v/3amSnylGWPMAKemWByXALq/J6Hi11kvDT
NRL2Tjozh7M+mcdqsp4O7mDiQH+ZZDD+jEYSb+V0pg9MFIn6nlkMR46yajHEA1Jp
pWYc2vWIznby/iy6Tu/4qCehXm4N6nyZz0XPMIRglgbkNncUP36FuthI7eLZX/5I
XI7yZ3eVC9M7b7lkYHnks3n0gb5lqpmOy/fyfilYby0EdeA/leCdT2HSn7WoKgZE
kamExMIzzCPYCFRd897JZyhCOC9BT6Zh9fDCedYxSyDzgDMIgcy0znK/bO2wcrj4
8LWZHbZ67dCWKHJUav2TmM0Q29DnzIGG1ZYvLbmYlKv3a1WSC5fNJk0xLs0ceGkE
wl+nvVFvP784jBowe/aT6aPoA2gKwaJvlkr215Nq2PeQVxhZiTZBc28h3JALF/Um
vS3kHy2g/7T7yR149SPwI4K9c7ThFI5c0ZgyeCNKi0B4FGfjkZPFm0gwIdEspkB2
uY66Jz6s6Y0T7JSVrhTxW6KZ2BFPai65dOHFqIKsVFe1JoZ69cJ6RT+Zr+vnvgUf
0gwq2sIZAHVegH7X7DL351VtQQKSatgWdjGPTLzQzI/uHwNyYzsL3tjHyfEKx6Cr
coNvk52jkzwXMIEJif+1r/0UyAYC7cazdGOEmbE4tR+MqEiF0tMhHACWCkJ1bTSR
Jp8SI2rfefWZdkArIn1t/zAPu4WIF+tseJnu4kpYJH7GXci5t5DIgZB+hcbcn2lA
9xGtSOdYJqr7mvX+4PTNs9Mrpzwq/twDOwu9Oj5ypU9vaqqevwWuEBOU0Ro0Ow1f
/WVHQEjwsvDbx9OxWbmasNgjVhxa3kuGu9cOkgpzaDeZo2ilaejPvm5r/o+44qMO
8KHVvAcx9FoL98J3qPlzDMe1N2NUr5bWQ9ihgEDU15TlGWxW1h1UsCN0wJJJGxUi
4iiBjy4ScHy98NNH6VrfXOou4kXnYltbwsY+VVATYIMsnjm1V3o4HprFU/uGUuM2
TguI1WTduIji9GIFQAspGdO0OU2JbsQoX3wwr62KIsFIHgu874Tpa1xLoqTY2l2d
bY4icT+PLPraCI7diYROfo2EEPmYsbTmx5yi3lDlRbxxviFrRIcZnYZ9eTLB7EX8
nVvJNiE+phm8uuEsCdZYbm/JD4AjDx/Q5dvCyKoeQGMofex+ohkD1KLk4ip9OBbw
4kO3WNNk3wHiVoqfLuslBEny5HjfifygH3EdHVxnm2bKJKcGBv6LyPRe8sl/tMvi
ouborodfzAaabCbLPxhvQp66fjw7CilPwbr6zjM/AS6MyylR5pumCxKjrGzPdGhq
+aYv+bidkn1SaJNvhj20YOOUDxMZGG38D2b5JbXLYRsQcirUdYerthTaUX1Y3d8y
THHU0zmHQCJuCjF3nHx13iSxpbTRcy8TEtsUn7HyYpgj6QQhUjUwR1doXmNXWhwM
9tQhYf7Y0xHPH30RkK25xDVBXGIJjdaabqsiuVo6Mohgzw2b3okAswlQ/dTlXe4F
R1zVI5oJYwyB+1Mye7xh1T5bp3s+/AqVHWQErfPN7bmTskrj1GV7ZA7NyfN9SMbU
COc2fbxKIHbW8wSBURzpmoLRXixU+vUYomaquwoEQ6al0NsPuvS8hrErWdBLgXNc
/6CP/JNZ+Ee0vQewKyNkYSfpBYNBXOsuEFCPk2ckyG2wdFHjpHKMvJFRI0h+Rw/j
lrHkuWNXajkmXZKhSaxan5QyWzlegURqYJEoOCFGSqRKX+4AX3QR4npbjo1Dk9Ty
0SaSm4V2XQULIzkUA5bxgN4DIJbL6CKuHe7KQqZLMTWsjFJrr159R+x5zVgOyvKs
1CEYRU1b67VG/no7e0WvrhKfLN4noPU40HyVWULQHJVEYz3h79VbAP3GT1Mj6YVX
dzvejq3GEQPb5ZmSWcCqTKlXZueDyAwrZec0pkzUIfPOoaOxiJueO+j093gXxpHT
vZ1zrTC6Ui9GRfVB5jfHki6ufPjQIuhQP08iMmIIJs68A4ORjxEQ3fzyxGZqiSqs
WzuqSHOreyC3RWj9ktACuKVlyVefgei8lRlMPI0+ItCaUMNwL5yKIYh/LGyla+9n
ObF8P22cit707i6DZsmJEm4w1jLjlep2VW38HyEg/YlY5kea7r+t/3U3XzgFsXCX
cDGtUeuVXepiqMOlTAV0eVqlb7VDrF3qPXYMlV69jOdWfxkkIYRn7lrlCE5ACIlv
jFbWXM5E9O6ZHQUzf0HZYf2uP/T6IyVSywYrHGoSSdzzZb8k4S+mGlsRb8ZY2FiC
wSlh6gUkJMXKbdARPy/xtg2fliSbB+UjIH+3kGtWXByjcr++sYoEgWFsHAquIc/a
i0bjO9WM4EVmHzCjedqH98yiCtp55R+36oPufFQB2qru25Tb3+0pu4C43vtPB0ZF
XnFnvAQCqXn4rP0iR5IQuEZkASb4m6LT4qIZ4dEdNVNnXohdSZhuDAo7GnT9ZBy1
NEMihr31N0KkgsCLshl3FwNNTkyi3YfFtAMdvWc9wRJudGOkovLoZs2rMRfT5JG2
2IKa0cx8WOPr5vAb5sX6sQiHtRwQ8pQYSnNgBEWnoG2jeDP7q758kajiBZRTXukT
s51Wonp4Jo5qSFRPkd0p3pximkSlgA7/OB61l817O6hwVRg674IIMeCnXkwVuSzx
BilH55gKdtbk6WlKMDC9G6O0I0zubn0JmaIz+XlVZ8xE2ZoVabUVvgv2wy2VfP9R
Vf7hi8JHV5e9BcYvg3UlNnMBvyxakDBCB+zHiDGgzWek/+Jz7CGcyx8b5HT3mft7
0p32JK1YUwdkTRBdqudhJ1SX7OcmTV5rc5EJPDTB21EEboYlhiplbC70eyFEbJcK
Wa998AesWEb8D9vdPOTwQDYUGoVsUkrOLWhYo8FJimQ3e+sijAQeS9vsE7H9OuWs
BbunzSWkg+Xa1BqPodki01HkEUGRyVeI6QURdGRtLD0TDHrs+0+Pf5sh6E2AQnJp
L7NbnCbrIdh20QyeTrd4HlWYjCmClMrDT48RcNDKj/FGXT5Rg7KSijSzQ1ckh2L8
vMBrhS2QtTXlM9BaSBU9X4aBQ1pOPySHujoN1pkRu1mbqf8XOlR0j1K323iblRg+
Bsv8xra51aqjWcuJHRBnzOFmVwuzq/ed81la6+0fDvxDJu2TfYIK2hlBjtQ/awGy
XTpcco/9xzE4HjLEmKDlmV4B29zklXNgVy0m5YwbNVZ7bBrsMV+dCfj8rn2E8yK0
u2GUvvK5x4+9tZrhcAWOTPGZKjpP2blcA7yIbqKFnXvKUGxD8N5w5Zbsq8gottCD
ebJ4o5L0mn6wJGA5CqZg1FtrY3Hh0fqNWbxet8f8Wdf98iu2K48iza7lQQ4WIt2K
MybR6e8/P+9TzSLgeJTTVX7cl9fOGySAELFfyYygg4gMfqB1vrJBtToETNee89+q
WD9vTkLUVZIsjjdnSYtCaTlXCgeXTNwpwZe5N2YvEQlV7azYoczMCwKRiPFfJlB3
ee841Aq1/l34JSPiGdx9sNWHDzf1SZxYNEmlWt2rPB7jQteRvTcMaAE44vsIaEyI
XAXH9naGRQxti/69kYeME7Zcmr9bWT5azATeoHXLx/wxz7lFVE99PBxCczvaCURA
iRzkcoMGxGLqgWNRAJuJb7c6pV0HrJi36nFyfIJmGs9Q4l1lCweIw0d22iM/fMRP
/gqS5Q5/yDesYZWkg69LlHiLI2uUjPkw2YiKJ8Vlc0PE3RoMUMW0kEGNLKdsH1nh
37oVmbwROaMTtnwRm6EGYsnCM34/salPmPFIrfmKXBzVEmEboyMo5aIX9J2WYOEN
kXD6vowtjhG9DqkIk05eWSJaaifH2DbmVZ3lCmGkvcsj3Ar7WHLYpKTM3n7kRv/0
6t+pvRAQuo/qCkRodTFZP2SW2OCIgXYlxBPLRh8GTZZeoyix7zJyb2FWjZXVSJC5
/vIXcdN86qQrwXBXbSqEQVYt871WKrJlrYjUymXpV7/ca2fXL0N2qnUSnHyKPV8n
LiZ7nZFFMJ0khJcB66HTL1Vm88NCWI73WHXf2b1N82pU12ZY//BxloYtA6kZwCwU
d+NQdkZ3e/OzpVz1mTyEylsSr//VCL5KxqAhOia+Dpt3Ouji2nOhwbP5ugCx9rp/
3JxN2e0ITpttSAU1KZkEJ31XP1jqAZSUlOfl1bKLxqtcYRiFBza4RZKNMM9omikl
yJP/bCn7s8fpghvqm+eXbreo5tU7HIVSAUhLCSOmT8vYEdCKVjlazZJsqkFNqbom
acVgCKcxmeXZj+UTYRR1Y8bgTMmodxIj4SHNVn1coiHi2/mSfFgPtlNXc+A/6l0a
zpaPYUGKGscncpcszlNLCyNEmtwnA+qyU/igaMgEwkiWk6EMwtxqvMSulO9Ahf7q
LGQgwJOOLPKBXyx9EHB1OYaNjjFeOErRDyW074jMTa/3Z6l3DskPdO+W1xksUqjL
NaTYIWnBoR3+kKsggkNujPeTKWgmAu4/L1x0y7bO7Q0XLY+rVBbhCH9frh9guwxv
us1MmMkbvbT28kgwxnEFVWgRQvOtl1YB9IrfsQcWbWCcvkXeUTst4Fhg0JE1CVN6
tp19+iPxhJW18L94UjDeqMQmB3tPSg5jwStjYQHAwAsd6+KUVi84Wb5cdviTK6R5
KyGX8r7vba9HtUL+PrLTHrB7BuHeSj66PQRkiVqh8E/19/Txv3NMMwCdrPccuQWX
maBw2F873J9rWO5f34gXrKa9ufS0tYw1BuPs+lJ5nP1goASoXAXZOPcwE9BZIKPZ
t5S8+e9mNmYpQIGEWXFY1pPrQwTkIWlqIjwnQMQatQwhufRgul2wpUdZqHOWO2C2
TgF0DH7owxIMFtPQ30+hEz0pQW/m8iYoVuaVcUrD/xULmAF012D7FIFq7h9nutYe
S8QG6/ZWGgi96L44/hYsbJG6h66FUmSoGxXY4V1a0/1VEmnXbwHmarELT9hT3FvW
PBgNLwQjGBMF3Zpyrv9W5DB05NmF/fSGtguj3yASsb0CFNFY0XDmRwgNgh+xeBZA
wIYxSM1m5AhyraCngMY8/hrbDDDhg6QqxfQtSHkKXSTd6HWaQb8pWXq6E6sHNrF9
J35lgAh+Elj99MKv4VAQGTmqjG6I4ElonpOVMXKKtfCRGH2KLUj9AZcbCfuHB0+e
XP5d9H5sJVSKRH2+n+Ghch4myOuKW3WX9ABCD+/DU6GJHynr/keSAOe6mqsQxqqN
NPR3dNVBSYIgcrRzEpwddoFOgJ1NSDXhya8aiM0xcyNIIPGAzCNOAHru/PKhbfdw
7MQNoq2T1YOhYO9CaAd5LUnMA6d37cFLFi7VPf3A99cfrrh3J03uKyX1aOZ9jmMh
bCl/44RKD1DwUvWzc8CNFDnV+0JKkRe5SoCx0RgvBZfERG9JLnrKZpGuSmf5fYoE
GWaohBfb2Mmgp2qNYmHyplCGzbAPWskUbZ8oVMoJ/OO97n3C62nwre+Ybx3wZkc8
/zpqh305HDhQtvXA2ji+7sCp6vK/dn2s4l0aX51aZPxIPWS3gENJ98tC7Vzwquq5
1rsipuP9uWMt9kJTaHOrlvSXDhYcfQwQi6+D9FdkBAKulc5Z0P0oNZFQQ2cz6hHs
9VHrv3JtsWs4j9I9Sod3zexXh5i/yx6b1n3s7f1Z3UA8tUGNFPnQcX2jZEhxU1zX
Ejhs2uASwpmfb0KaCgc5agvaO77o8KyzVaFn7LWb4wEoIu/dvb3toFeJZjmRNDKo
S3WH/IkyYfzgeFprs810XwAHGv1uQ3/lBmQuREEk9LSVq55dN1l4Uvj2YLPNUAPp
+jxQIgYhZmrhX9e8PZQF+jjoY9UDBwsi5JOxvyvvY+eNqK9wzqR9WECh3ZFBKjUN
QAyRp2aKZnxiRh4o9pEfjTn6hVG+m5guypMzf2enFbsnsg1ypprT1biuWUH0aTJW
Sl386L6Rg/h4BCFkGtL4QocAVvp0nllwJtBEoDPUqu1MiSqaFSm+n7XM+jGIztSI
o75TRyy3GYocl3b9p4YCgtvvsfRloCoqLGUDvjlC4rkYuGdd2LBOnBpYmSoIPtPe
hQYqpPJvSSnF+z4PXxVjy5iCLGl7X+Mxt70ufwJj77l20LL4tyivs0bUVwT2zBls
04+MD58J+fZt7e6UkJMB+bkCOiI1HlNU+vh9Zc9N520Ihla6xb9LP87M1GkIOuZo
vYlijXU643Q6LlqFGA2gs26NT994+XmXuHxFqvTcQpjX6dx6rIngol0/OUSpn15a
1JN6LoxSM1xDsJWhdV7cufCq+GKcskwXb7OpWl2UWkBPetigLqX4f679l7Jqv9rc
abM2DLFUMfOJA7LVmkXQFOOCBJvItAFARN6rllTrAR2QJF+DWmw6A0jjN+Q7zwVp
KjcXWSrYccWZXdamkNUcJq87q/+qDfyQcpFGcDBRIb5mNvIYVq8GFYKtTi9G3zOV
BiBChtgBAcDjpUZPj6RmgQ5LlRwXmX1CekJbSaSPonwRYWwZqpFOC0Ql5T7nwvXd
VvpGl+jdHKwGU+4VdNH0fdz+vyUM9spJlhTSXzzSMMKz2bcV/57JCd3btk8SznN1
877icQaSsgVlOv3W/aDKwV4C9i+hli2T8ZqLxcAsVw2v3GRcN5Udu3U/uZsi/8D3
dEXzKLImQYtrxaKw9m2gODDd3QCpF8eCL0IHHdnzudhdRbNl+EK7tVQDWHPrByDp
lYzKWSw9PvE6Tzr6cA+fchP0wBMrDkxG5qllSj//ja+eh5r7DCM8DGz5RK5Dd2T6
H3Z+CxWv23titdvPx7yD3VVMjmr0vJUZmEQAAovUzV+wtOyU5fjl8sq0+OcEUr1T
f3rIuYyb546EwzW06e19fBmfuJmEHz6+S+RQWV1kk+gqB8tgEI0FZN41sy/iu2RZ
VsKYE4RsOwJgbm6Y5hwyDxYEhuT4pGnJFB1h1hG6N5z5XEszcYPYvHu/OiJuNty9
K/dykpttmd+ZWpM7UrhKsMoodfao3d8CV+GO4PJ9X8T6gaAMIjHosOzcxnnewHD7
NvRHrHYeIzaLKchYsiyvS8kx72rJALHP9wFinkw5RVYJntNIxLGybbI4CYHDXxcH
WmBRD+w4jqj3+KuDXZnTtVlklqo/sEU2lnVwNy0cwPzPDb0yb/KyGR49rXHCGb/m
2UsG0UNuCYfQ5Ly/zXVwYnnad2T7jH9GUj7YbCGYp+pqgylZUBcDupCHmf4fJLD7
gJuNyW5JEPwsJXHXbDaQHOGkarQs7NnfOFcekGdx7KMI7qYKWGpKVIUozfy905xz
li9eTeWIihAS1sSZ89Hky9zDeXeYjLE1bAixIGo94IrhgGAxUmJ5Q3OX4Jrr+N4H
CKY/Yu6ZQEDvK7S0uyeHL0s2YnfwbScabzauG8mXunQopH7qRShfcnnTZlbiMpBE
ksYF+8Ic2x7aQgF5hHPNpS+BF4l8WtQ+GhglpZ0+LVZ8UiVDCAxi0Hfrs3r+LCVa
xTG2tFUc4MqKz6jpl0RFyZ1nDgNjUpavlUfvtqaOMM0wq/VrUGnWd+/Bdp4P6FSo
QiENZ4MBpwwmXEl457etTKhjtPkVMLqnlhptQpQr9Ugj+Zu+YxjvOvZ4MWO1KVJ6
RFR7qOyU60ou3p82ai7glinnO8zpt449Ebu4ENgQw3Ihz0RFaBMTyim9NOKhYvRg
mMuZpPyZCr/iHkIanL1fE06+DOGXl8ZOYDJ3Cd+TyztsVThRMKBSMMSN8ysMLHQO
zMcl4Q+tSiSc1ABMnCYOCnpblBbpI7/8Y0o7YCz1punmWLXACmc1Ckmphi9RP6fx
BEr+gHBJ3MYtYc2uY9SujWTXBxG43d5y8zguLW3gqSCYkbQK2aKIFIsTPcLF3p0t
WXaDTn2/YhCJs+CFhJagGFFhBQ6RUtS95lVfe/VeTvaaq9HFL6OY1jGm6qiRtcJD
nOS2a0Eh5wmgMdYdGJPfHQY/PlNQlOiL2T0eFx71YW/316FVgX+6SmeANS2uPqlS
uDDUm30zW51nX7R2uRdwVcYIz66oAuzxq1i62UALCEOtQV6L7Mb4IFZrKQ5ANn3S
Fvz/qKCYQQpPq0iEUdBzSJgOgPnZPRAA39+fWqAujv4Ijw1P4TFxGV3kpAsKQPmG
5aUPyJkubYsq55gUIuZCnUewertdtJemSfIGJvDLexXeAEnm2wCgjqbTBV9jiPan
P0ASCYAJzppnkwUCacKE6rcXQ799nxQzTLgdxbe8bTyt2gWRCeE/EakPN7kPbH+G
Cv7Zxw/tKLBuVjWuKWGNAUmAPxRhiHH1dMvPC4y7VxN1ivm4b96vi+wXj9LIcDyu
410Rbd8SYKZqvf29gcSRw3sIyhWQ00dGPqQo4s1aVOpDBzvHGJTtuzVZHIG6ca2x
+RC1N/ZpGSop9fzg5xtGfSJlsV1CV6pTO28y7+LGH1CFfP659IGh4gxbUrzeOovq
DTSMo42zGMFQTV+Z33PJq7QCNSaj4ddy43S9Qh+PODv3O/zgJjhtTWiwSF7SYMYT
hUq/eYxN75AEf3Q5awzEEwg4U35hItJvQwJhp7/2NSm1jgKyPr6/48uydEw1q0Y0
GdNV3l38eQ8505URv31xFA99SMjDEunDkQTJnYj48MihGAGtpvKi+/cK4vsH6Hw/
5SsQFIrDat0SCZ1XPw7SuWTDKNEUwp1fA4ij/XbH6W8sG4WOarGXdRZEkQJd5Etx
BZ3BVIMV31ekpYRcsnEwzSWGl0ozk4+RrJDviraVitCWpoP9XtCU/oAT7NKdTBHx
o/lA70sJspcR0DVpITzqNzwQbUlh/i9X0Lbh/wfLUaDRfwXQ4Qbo3E0XPQ0EItes
w7jcGFjshezTvVMGpg/j9e46B43xfTGyyIlcIsl0eSssfJyTr2+6PwknNsJaxwEQ
JZ8tY196qo3n+ZZSkGqQcU1vJIjZ3lbDc3UawfokfHrvmCD3sauZXGmTEqF5N8uM
ifByGsnUwUDwNk5EG/86mfHRlSQHnRbSL4KOULUuax9DxbtHAJ30v9TjzZRD+Uyn
WLjRSavTQt6Li9nMyaPLg7B5OCYp3tXStg/t6CsjKERHk5sSdO9JuRBEcVn2N70Y
euO5zla9sxdzJDjDBB4ZwjCX3QlLUhocIZSXSAf5as2mF7kFlU0mMOMA2sN2y7mK
/u01WKyc4eNpm1wQWjeCX6/u+aLq6IuHazd7FajqhUiQeZZoKXLOA4DoalLIvfoj
tDdn8QWzs3iVU2VxM8fRdjy1+0VuCZMQ+KGpiH5iSdIqhjb1vZ1T07+HK2DwmZpt
GBMoeHCW3rmXHZwwzoz9LHGjfnKpjkwzpVY+t9potE/1P9PNxiU2mKbwVi0S/5Ij
urxOk7/wM/CClm06dEDF2SfK2k9404nLtx4/0qk51LV3298JKRwFklbDGiAbjjiw
4dxXFK5OtR9OdCjRGu2r4ahNTwyfbzlzKbYJAEPI/CVZRDegd5c7VYoUaXZu9ddP
Wtw5KnWySoGW2e+u6DVRuYRqaEKH8CUw74TVVSoWUEiXU9MscjC/9KDmpREGGQyA
jFqJN3A3Fqb5smsIBQTtwgnxxNTOlSaviHH8U1Ft0KtHpMAwYkTcGJfOlJ8txsrv
cwqdrXfww3IewtYZNv+0q8DkTJQsY6TGIAKYD1p2ehWqhJddetCugxAamFDrgzLu
04gjkbG+7kUB5+J4iZ8WmHacr+KLdfemJ1GnCZ/QbXd52pRH0oI1hgWRQapsJir+
CAa3RkSUzTPO0NizFKOtiRySdGaF75q08TWjV02CsmG7WDsPkWCaF+uzhf7G+jfE
UOBcIFG9WCtAiyS96g/i9Cxr4HNmmZCOdHwrJNFuaR68DD4D32C/Wk3qSUsGirqk
k3BShJJnmeMv3lIZOcZX6niEQROlypSSoOMSJWQVgP8NTjwqHQ5yz5CyrSVkh8y+
CwDXLQ1yNCCxT2kB0OP/970FZb7vqvyUqqL2ch06NAk/EdLaPu0fEUszlZWqtON7
W/gr2ZY3WyKEWBFpSxa8ozdTrRXX1pmiCjHZI6BAxCQtXYPjPPTW+2oJ11VAX4Vg
7mQ8GBo40cj98SBG113vXelJALUpJ+fNbyJinnu+RLmQBOc9nu1BhOWdZO485z/2
k/se5k08vWrdi3WRgfNrzNb1F4DuMtfuczguwswsGJQOL9cb+xOK+Z63wl+5OPTt
wyS/WhoP1YiFbjPbeBXg5uhE7wOAL++RNwysZOFlTufrUAuhNv1ZKKiq48fCF1mT
uBTAU92+ExPHBCvjTJoaAI2hEMK4zKIuel/Al88zpcOg73WCMuPs6a9EeamBT6qk
MjlJmEQTxWMJP0GJH9N1FKJhphrej/seTycxzfnLREsTnRAu4WO+DiDIHOgitn7V
tWrYnpl81LPNV46ws1XkcMTh70u3hfLDvCgLATIjtwlPN9vN2nP+feMrMgYsdIzm
hRp9Rl7WBT3UCalfrthOVgsuLoocMuOY1nSnG7nfOM/i4yqWVLgzp2duMkRm/95v
DxwuqPWaEu2R6G2k6Q6hxH0o3WIbyBhhomXfqY569JHWuOmkH0U/SV0aUYhKFSYd
nXBeEF+GC3hMVb3hfky1dsBnDCSFurKOvRdLXQGviV33oNWefY9I8i5GN8HDI0lZ
hF82XZYiNDK4s9ePYwlwsOxYO4xkCvvOKr9UefoKemcciCi8Nfgk0VJbrh6ZQkA8
kzfEl4QOYcbtwQPsUi2i7jpQ0+Q4awb8vFRtsRBB6s+6XFwPr6ZJ0wuiArljlxdS
Yt/xRSYfSyfjJE/Xumyqg7n6KTcmLn8bKpMPsgPZWVCZlkRJ8/lE+vdcBAk+10rR
/DgE8wLJv2jUVij4IV1EuxdbRf1vA/WuwjQLwqXE8g478j9ILqGBStYcFRuU9d1V
ityYMsTgDSAwzUJ2zKXgU4cC5uQNJfbsTlk7QZvUx+D2x6slQKmjqzFtfb+OHX61
fzOHwysxK1WCEW1IwDatjqz98UCXzdrgRNf17zFDyQkjsTcrp2c8F79qpopM9fVS
YyUP4QB9CwitTI6fhjTETleTdTMGGnJykvGt7gEaVGvQJ7n7CxgDN0B6G9wo4yZw
KzJkv69++fqG0oN7F7+csJzWQ1CJXV3X+325eT2rQFhk6IKrcr3QE0pRFkGoXQD5
EUPztMXiBvw4H3IopT4YKeceoy+YSX/qHXYb27puAVpYB70h9Cws6bt+kDzyPYR2
shureZnNFGqWtVqnb2ED2cm+jCpMpiYMIyIUDtlF0AnRbwki805AFDE4PczgZPJs
WuuZmV45X4NB4jLvCGnAfBalxtfod/kZciSXOShf67V+sq1WCVLAMT1DsmF5m70A
Fh8I1pzUi/eHYhaMDVi5CQSKF/BP79e9dv9Z5Cz25ZmOYSzwJjbIDb8CRtrF1ptO
LzX6Wq+d4Sp8hw/v90WA4KvOEU3sEaI+DtG/1FPOg2t3U0vGdrPKPwJW+e7ro8mB
PlHKo6OOIhVlq6m2weHkgroNNWrgyAc3detcqvDGy0rfxTzX7+hEckcNHQeibGT7
ZzP79HMWwerDDQHqNUYPxEKyM+tjXTxsVccT5wTpEWC28AF9/KtE5bljnvwtBr/t
gTviDEnt2a7zBZsjAjZ/RAqF6bwlIbd5QOvJsQU957noltNy5yUq54tNgJd3D3LB
xBy6bvGd00G0yRj5hL2l7OlApbzReyxfZkPZlc+nN38qj0akWFPy+X2IT9pIvWLP
0WVVsWSqzVCHYAyGFDvVrYF69Ga8LsqLwxedmazu2ErAxVi6FkUMD01lDWU4bXAQ
cTPBvGowW9g+Ihu79BRljz8L7RyVVj9yYPNXI3LNLSLCe3u0c7XdfXcyzRDTglVg
1Q/e6+IIRUGw9SUtcE1i/vIkYwXALO1yvAXVBbiPyNrZjHzUElT6q19n3DOperLk
huKG25gtIjxyaaSyKRnIigaY63aq1HVVoUIcDU69sTp7lai9JPd/v6PUaUgAQOwK
x/e5kZzE0qvLwE2Wdw1OqYVKY3XrMz+ASMYiwtA8sp3gaArLmLBy5KrhPh5tEmQu
U/asfzJoMjcrOqjvjH9pw9ZmjfNpk9cJkXPx+SG3YpgmKhp7dORn4/uVti4IbAAG
jqlPJ4wUya/HrGKbL9dr2uujPxk033mK0heOw9YMWit1lGeUF7rd9PQ8ASVekJWF
d3ksOkZ11lG2J2LOI2oJeHh7OznKymSZgPIrhlNYwHonhIp81mlCbK9HR4LgU6b9
xDNVfVvnmIKNDwbBF5vePphEIbE1u1m6y5QVt9ZmMEMEoEKI6RTgcPz25M9D6NUH
lcYjhZixOu9jrN6CFpCA4OfdH5tyr2EZ8IefI36lsfODgjJz4dDs/MBwMh/5y9FR
iPgG0RdWBDSzoWEZ1ORMEvS1BT9eghTObI3zRgZwRzdFpNOzVLoJYGwJbGK4m/9V
5ZPfsYnav24mMdVm4WdCZH4Q+Y11Z9jSwLdk5V5Mr0uKeIHpuY1DyWIlw9wybC8B
pcAj/hM6jxdOC3ev66n2zTdxOGfKl4athE8bVV7FeIzQ7Fdq3Qlel4rS9/LbpaTn
IQw2dewKBmygp4cO/QORNyGUhs7IkD67RMrCLy4PvSQRF+39Xi4gTLBrpa49RWTN
9zLgrzbsRHe8TGGQ5a4xZj3a61IbQr/nQfVuaTQpSpU1/RU1Fj54XDxDzCP+xccv
vKK6gPW+Dhl6quE+7m633MLONXWnN87d+gR5JOwk5fibizD6hy2Vi3n5n0qug1dZ
d8woNvL2rBfM1O456X7XulW8m6wYKIPWMUL58YAD8SeEXUcz8DFgVi2WDSnIeaHR
rMekAe0Vi7R1YUTGX7LlAOK6Ugi+h2xV26l0NwPBnwpqoEw5WNg9BENZjUoU7MEk
D8ZZJq4NmkgsH7oOZ1WDJtAUw6qUg9G9lLQufCT66CJJNx0aYQ7Xmz7udBgfkAK3
RkKg1VMBCCKnlA2E5csOdXhU1Li1GyZdKzjsyRavvCMrI56dIp46zzNgdNOwyu6M
Ae6AhzxDbHGFYBHCqJC8mLMPl9lptKWoKuqILYPtiNMV+dunbtbZ/apJ8lHAFSht
MmvMHXQd2h2SKbWbyIYjPa1Iqphddok+7/k3Rtz3hfcHyIiNtWFM+EUvmLDamKCP
NVON+ZnBRv/Aiih3kleOrxVaA0HYQLjx/owU4nE76MAdIMlKGz5ZUtH0f5o7iwai
IelAWt3eyoR/9HO64hkNA6m6w222Q8HBCCDZuO2uOKuCiqDjKhpx5GD17U9aCGuz
U6N+3Lx3iiypfldvZfDDG1RoDRiqTgfabc3FztCTFgvvCEADVB0I8sWE2IxULuMP
XEeU5OAzysqrorIHvF8whm9xTGiF4Yf25tC+kTS67U9rQWQety6N9k4j+rQoIK+W
Av8lrblpNSynXs8adJmRlYML6rNr5YGlNbpWRF1rKzR1JbCkweD+tH2c/UlpSlPV
GAnjGv8QTkzHBpLugLTII4lw26gFFAlqk25oqmkITuxfTpTZkwFAXFDFsSjfEekV
nyrG3YCWjzKaIa34p04kgmbaxC1io1FThdet3nHqk8RohPw144KEIPriapS5KrTT
69g2RI12kqyB2D66o8dYF8MzGQBDGrEcCpNnSw+Qu3nL2NecxwfI8g/MpkQfuzLy
KQji3yInrPIv+1DD0QWTXTv4vfY43o1GrAZbN+CchAVl++lYEW40oOtLwLfQ/bkv
0ircxOYMylIRrdHrGpbZ7Z2BtoMaODqvFRAd4/yW/H+Av5B/w/C5+0nh0qhsuQn6
Mm5rSbZLY+Ta73p4Ceh/eMNOA+R2HCkpRT1dOM1NYQMcqycHWaqoZZSiq53QNvPW
ilsShtVcyDzvtOIbyuGKWM8pBJRk47dC6RnVDFI/liL/RClDExQRlclQepbGdADk
T7T58LG4eMFIH86x2uSoVeHZNv74mnibnHt3oWLJuxr9gHCeL8WNRQJ9bEWg5kOk
0M65YWKHPTYe49MQZdCAVK+CMD4QWfR2SBd4YMJQ2B7YA6UYOyVUg/5Kdn8vBwXi
zij3WeZk6F/AZpmaRz6IeYcSWY1DXGqk3iphEPkGJ9RTYGF0HswpdEk8G+p8C6+T
kuAB//GfQwZYbBS3LxpDAWYdFv92jO+k9fyO8qmMPhtWIEVdcM+lM3UoY2APv7Ju
wcYUHyujHv7lqp305gfUQMHNwHUQ0GE2o+es7/2i1mHf+hPOQzdt+iBvY9LTMPfE
yo39qaTyWYks0YRYM83VDOFeuZd1mBScTBJWDBeLfyzQ0yFsnFXx0Gm7glvGUmcn
KsWm55XWB6rZAxNC+8UZjJFQWEJu10QDrgsRd7CbwlhGKTtuztYC0sDJan5NZZ3u
jKsaXofLT9yQwQ+oj87fOzJneZB9h21AYN+TMlFVUyftHlEL59emUwOLdqvE9EqA
Jh4ipdqi7j/rIcHY+ruvixH5ifEIxqUGjk/jZAIZ36U1Ji7QJcPoKgKwlY2VxD9w
UqpDZPHlLY//mpZAkI9VLF4EXYr+HOVhygRuCwc7mtI/JK8ygvMMLz0WdDhA2xh5
uTuGn5j/8859sk5GTqiDIXwGKFwWMgUSw2rhBhEAzZemh9qHrr8R2C5Qyv5abFUi
U7Vj5VsLkadEGUXL/1XD1XStZkZzW7zqCDhHlOMr7xNymz3dv/brEJdYhmGGKXfX
/shqd4H99gRveed2U2QxPsqYQpV57NOT7U0NICtBES5k0qVT//BthSm2oNj2gYBj
M0AocxrfiNYYVd3RDY9q0xrLddv3lUqeZrR7nwpoHUwDY+qKCmWowkooSiAb+6Yb
CsPP3adu44DKtk+1Zh1HKVPljOKpWZ6wh9aRZqCxw3jeB/6yT4Cvg9R1Wz+CFHKT
5R4Qb6S3Bz8KL128STC2KcRDSwMVdt5u9VbeDl8uAcQ+shPp3VPhFgMyIRJHvWyl
M88h7kIg3Yf6azWNQiB1YsKpHj1eB/RWC0VgX4uInqJVksdCMXb44hzgAXQqCsCc
vhvRDDhqEmtMYYm4DXNOcnpWmLz5IPLhU6WdgKLdzXonuVhNquii7OAh63favsmK
IuBk05og72Dbz1SD9GBwimG6Ia+3brMuHEWIxz4iTq5UqHgLBMjthqMBFAtIN6pC
+F8DMwrv5P2GdsvoRjstI/S9SbNLmD52PxdBuxYmTwBfRd0tU8Eh03WfAQWc8dTa
sWPIrusibGpMBl48MAaMGH6dWYvjn+/jKGhcIBwabePFG4r5nxYLXoLxWROgRcbA
nf47PPZl4c2l8GpHucIDdw6wC5w0KBZc1mQU6Sdj5N15ZIVBM4p4D9/5YxGH0WGZ
f44CNcS6Npn91ZlvDln6OeeX3zmWLPO+sa8KDZ4NH4abgNjyENcj2Cx7W7tTtl6/
sH+MFT1dlrIM/GAO3CpJ2mcQnHtz6zXz5VNWZ+wKXMliMzn2Axl1T55FMC0lEgLJ
MdM6050OtlO1a5YSDMvI+bumUbmURbk4E7Fx/ifGQnKJoLH9hpXRNR8YN6thdeSJ
ORVgS0vX4EmbU53MpbEoPxxLTkdW1J2d9QnsferdKSNr+rGGu50bVztoTOnBkHAB
4FV+LMiuQ29wy6tS3sDjOW68wdu/pdThzBaLnHho8K69sSXnOEGjm5ZC7l0AzVDW
hW3R1JPZRNb28PxTFCcxsqT+x9lwV5OrXsifJarQoLP4NUtnU01/EPvCUjDIlmH6
N3laWYYS+8MNNT4nvX1UQPa8UsGPU9e7ZgsucCTaTkCNVS6m9dmjRHnIxbhOaSh4
weYHS5Ag+xPmycBLlXHoLRxITboeMX9k97KxVKHlEf3AStPmh4i+20YCrCOn5Ywz
Fxf4QnzyW7QrfuG2MZNAX1z2hHnW0AT0Zmx9A+xE4thV9w/4KlE/g7gEWK7JFMrm
kMP2k04ae8AOkGQHrNGkjxaSnmMEmmq8/2aWUw2FWV41CpC9hR/8T6i/lWLxrReq
YMZb0N2JREG5FhWcDn40oP1zefyZtOwLscDJTDSYz7S4BBKweDrGVdCE9bVbMoyl
ZVUd2nDQzBOF540AiJlYtWuvKr91r5/QB2naufYk7O05/m+a03MCI5XWo8CCIBkF
/PbZmp0MEEcTW+6tWloSTzv61lkPUV46QXv2NXdjr2QeaHOuqJDOhTUPsdb501cX
yvkvsGba5+cPI/lTG8d8teL5gIVk/dJT1LKRRyp3kWbypy2+ePyYsRN5xnrCiF7a
XL3nO9ARO78epIHgnoZmuiJPSg+WkQ9byd+HuKMhCGMXDPTzTWVKTUB77PNe6cgA
hVdlEuW6rmDQ4634XQ9dJvSQOZdeuzOW1EzrxuaKZGIB8xWOL4H1WpEFGdJppRLD
5+c0NYuh8lPGwjHLG6HEBOEoEqSYXGTyxtvFLBWWEW5hn1u3ECeAazrXj5V7Iswt
tnApEnoLUQmowD8I/AsVVg78iFs4P8CWf06fh1hERnPPbZEmhOkc1VMSiLX8VcLa
eU91NNrAlWOLILXsRldoohaDeDFudf718ms9gyqiXK+UnbfM6W5JDghzA0OrD9i5
ruk765dBdkvv7a9y58Yc0MwpiOLKQmitZgdNp1KhT9iSJ+sstUCsEfHs4PBB/SIF
/kpJ0b0PIpBKNbgnY1iECMs3XnXYrhLu2UxJjezWaMDkb9RJgeIOzr+/u0LALSpo
EgTCDDBLcTh6c8PTtR6XGpfl8LtmBpTVFyfMVQH3ED4HwtDv7gH4ceXDYua0MGwW
p+RzEIf7Zc4GiZUJ4jRknzkJZZIiBr8jeDkgCiINyOsLXdRQ4fDUtHGhnTOHxfnx
lAfjOzR7Cu9ootVl1biZVUvsU8tT9BiEp+7/1lr/YQKr5PTDhfQNm9by27emFhhu
C8waj1u8B2/AfKUesvaketnS7J0xX+4Uuf+UvuL6Tqs0uJCBcN5Z/6FRs9e60Avl
iRYu8MiDWDqrXt+QYimKWZhlV+4CvGPST+e+LYssFU6mGbEae74UvjEHsW8FiGQq
kREl0p44nR1BYNVuXPx1eJuLfw5cYX+THhLSw3HHB5RNpTXImD8Keq8F3m+MB4PI
Qk/2YWNlzREHtTNrj64+QS3U9Sgoky95LX1TPrVAuJf80Ft97v/Im+mB1vGHJxjc
FK0S5hQG396jobkTnqZi2DjaYYJqeyIkN08AiXnu+TgquZx5Wi1Pbp5oK9mz5Xgo
eW+tcTJD4vIcbp9JlwMKZBwF47XwjynxdbHgotgDre5un+EF9saI652oC+eHO8Dh
jIzAb8tfCZRSf5egpBHEvm/yV8X4b8F2C7h0mr52g1QFzf6gtazQBbAxAtzeojk7
aI5CHpBw2Nv7GVRGCg6uTHpOiUwrH/yJuVsP0NkD26SZILM2OWO/CunJ2gQ+rDEO
Eoe4/EU8orpicmbpb3Zlm+l2CcgZf8y1YQKRylEwDQ4ZNcSpLU2fjUfB3Ud+AQkP
nK/atz4Al7K333fO0GdMhzutPzomJVnGqI7VVHk9nPM25xEHNf2wlgUP2yyLewCu
oK//pONxKsFfEwn353i1jcL3Mf7a8+0b6YVhsEWNRCNSTmG1lVP8BhIFDNFhmzIn
gT2Hzw0/QR/qb/9mFJkONZu3G2ook6NT9qKsMzMCDTqfZ4H3kPx3LQetfEL/Ey8S
4Bz/6L+I6hfscUyAz2tZOe94TOkf37BTacjFZ0loGTfcKhJP8kK+JFCC2nchSUKs
lTYKxIwIzsO0l/aBQuJJzA7GXPyDqwZuM6BzTkJAIVInUNRZUX7QLEEB9OD6EqyJ
E9Brnal3VdDmQAftX/l/DWz8VlXys+EyNb8j5nOVA8GUev1aLkTnb8y7EojGo1F4
vwegne2TY7624bWKYQw0prVqjraU6rMyC0mg6/fOf8Bhhk7NtVMqruQsV5h9SkFr
sbAJmdFmpwYGY5saLXWw4dx/2O8wx9PjJsdLFJ7rWNUxMENJOa475dXD+frYfdqV
r/H8Zymny2SD4BXhTMMOCKkXOgmMe/vsTgjeRcAd+VBGF9NNCZr2BJSACx+44PyV
vS6+Vb1y2zTvDXIVNVYBS8e+w58ofF09odROvFdn1o6Ohe2fIvspbs/469oAut+H
Bt2LRd79QKZv6pwasx7PdkOF4xDHY8QbQJwyIn6uY1vdTXc+ADf8MhRTdVhYyWIo
KVaI26X8MHwI8zVInGS5oyiKKxbukuJ+mR8KMLzbxOzCAd/L+TANpDWgVlIkR2se
Ps98ZvBifzelT2F/K+/TewF/0k1oiZJKft15/30AaAu0V+MG3jq8JhSNGwcebBfr
bb37SxtIhCC0XLcCaPjK3yMN0O1QTnudhfB75gbhPD3oCHvpXjE08OIodOfZDBwX
G6qEs0azITTSdw6HS9iLWc+SzNxP7MSzcE0o4wees7EX6ILMeKLTp1kuQSDT90Qg
rvimT9H5TyCieRuMEBzLwpGBOmzXST5YApoEMotYgYyAS4QSWEXriDWhLwYDAlLA
Lsa6bZ80/ZLiL/Bas8mKb+iMopUuzW0y9KpCreP3srTjtDrlO5tjelq30OZ5JzSU
CJR6NlsZpA1UAOQX3L0gkrTNBqYvEzeo8VaiqIts0qm8MTidZtb/djbqR4WWN2//
EQS70ctGONKXitMGdHM0XuYepiBqxXfZrFcAO7ixeF0ZjcaqRSVkyCAoFc3lVdPX
Fc/YCgrjr1HLHUAWKvczgAHHdQ0pcPMyiD9xyWyLGdHCUGnWWvE0X79QREkdMX75
O7WgMLzdNx9bNNM+mgawHBbqSxasylGZYEpV7rS4f3P81VBk1SD9SYeRyErKs9jt
7BSam5NBb+piRujOw6xbMYFU10EdNcEB1tscVl+TNqk3xLl4rXgbTpLsQt/f2SNf
DjSBaFItQP3Tmmz02gLrCOtqnquEqQXF9oJVQjt5smIL15dSdcixyrA3oPpnJy/+
glztntgpe32nW4TWt8+EvvJaOp6r17kyq+BqOduugX7seEBbPivbFVkMF09BFDAI
UMxLNBm+X1LFDpoI+oe6XP4Er/iIKp3bFFDPQqnEYK7i7KdsFe2dtJ3bpYq+XrS1
ee+L5CjKuXNeEkcQnsUOEVUv3eBH1Bfq8BFo0J2L82RX/Hnm3z9WnxkMK49Ug6e6
+ApCw9sYDuCPpfL7eMWHQanFEV6UVMEmAhwicnFGuz8wu8JT3A98j1NM/KEDKw/0
2+38FtbWr+UpiREK6Ct7iQ2uwCMrT1wrgy3WjjbBXF8mlke/YRIv3DaGUTfdo1A6
XkgZEyTxocYWEsApH22Tgab0TU7pbadc0sZ4C/uAl1nuwCjWZJwinMfzntV1qWFZ
2fxwH+rV+Muqy7PRWtpvEkITrZwL/11Uo3qXFVrKz9s9Hj/nwZyGpDf0yNqINJzI
xJu2QIkVCM5W2w/4VrgqO2kJ/qSIhXd+8qGvHq859xGZs+Xxifk/REMBfGlC5XLT
KqFIinXuPVt5AilnNNUTPR5/YnXqkF3I5XkJ3eFtHntA+M+XUPL0HdapHkLPvUPb
WK9xvLNyYzc0q70OUsWyK6LXL/y2deerai19FsQgg/r3rDB8vJOsTmrI/KmLszJ3
goPYOTredisKkpLMILm29musrWV0aVEhWyFbmal3sr5kL6yvu31/aeIvEql9oWen
WU+Q9wzm6vMI9cCttwSTXBU20EDxf+Gwmgtxcn5+Yvo5FWQb9aU2xN7B/pvH2DvF
KL8EWO2JWA6dNAkC7B6n5khWA7JJKSE7140PDkQYQCfyZh/D57b2C/Qcw2RXr7nY
j7h5JXhw7IlKTiTPMSVjgIldbeI6ZxIVLFZii9pUyg6lTgS9kSiomLYM897KHjpA
N/ZcBQ+cYWAX9AnCe7HY+b27cL4stz/hOLqsHwEEuRQ1P8uxaclDpir6eL9mx/Jm
HDfNVe401cOXB5+qv6998PyYa5Z0aB4Om6Ahs1nVr2wsxdgdjghaE03TOQEDBpf7
kZp6bgDVefAg03dcyFeL+WMukeZ9cYLnmQu6iun8pmSrg2h8Eg0F+5PDGopZMWSW
2v0bF5FkZdsoP5vDy4W1ZY4A/UwTVKbWLYmAr3JQesTcwnoInopabwx2bsUJT88s
WHFnpDl7UKsIBCQSppJQat1nf1yeFIpSf8GMGv0e0tMEdmrGWwAaWqQfZJEaXk5P
UJwgh1BasOXLxFHKdXhuFrNx1s0DDWn8jvENw/3RvKAvUi1PvDItKyxBI51HQn1/
ggpZpCbvdLhvboOACqBT6jHq5frEeAhYXW68txqtwnOyzmDbaC4SNrxgda08zV5e
F8rxtj0pCRACB7weMSiFCQH3bEnMLeMPAT2tBzfamKbxxnklCJKNsOf7nXmO6xB9
52a0EgoOr66ShcAC5cCGSrHapQdT8sR/pStnSeLfHaqKXxxAdDQXnsUBjMXA0+sv
19+pWMMEtixoD4+W20s8J2gvyDaBKoqhkJyULdmj1cvHAQw3iR+lh+qoCRFeK15u
/eRnnA8RFJoxQKaAkkPd7RwriUZcAaUBV0CKKZI/fcG9Hhd+ZTRBHhrPfRDDU5EH
ZvOt2SgMIPFOFOxuKu9MVS5N+yqIjueCoMrwTIX3jrpsDtzPdw2AfP4cF9t6v8HQ
E8aO4qaeP1Kb/4Uy4Ss7UL48oyLOcfqm4P785tJZhipA/pkpv6ossedWPGEni4M1
/RuAJqHwYTrG50azkRNpZHa5gDLnN1OXss8beJnkYSiw460KbTKQgJUUzdXcybNB
LBxEYrqRzfz4oo0ytaKxOGc81zXAduG5tnX4DnBp625PULOErLos1xZNzurRgq7J
kT8O3rG/5NyBPcewpqtfT1R1MnKnpLlizLDi97z2jJcNG+GM82sEPmG8ut8VWqzR
fqTG7dJMrrj0RhnhwAmtXaF5+6KpDmuqorGQ4M97LC9mheWbVNz7TgB7FbW9eX1V
Jz7XyhU/N7Ags4skydRdGWVKKMqTP7VT6wycXfM8bKqT2x+SiCm3isNeMCjkgL7j
tMrZ96n5jjJfuTTsI26XQXr57sY4fng21FKLzmZPLwrgmvvHYknxUVBr8NELSvbP
DAOgppLX0bSC+HxhUSYN8NgmlSVCzLDdj8hs5hjikH6p6jKklvIaNVOZ7nhub1t0
b5IAvNDgn/49gogSbQyM4EHfGvTRxy0S8WUWraofMKMZRvFE0tP7N9PuWBCblRcK
LlLgbiVxe5n8CXZGkjpXIgtCWgq07d2AxDIzvzKapfrRKDa42utwR4PYZ6pjtxC4
++ED2AJrCwQNpdzB72M+HU8/MlpuiBd5Mu6N0dGIEz8DuNHDe5jO3wS1286cKT2w
4BLMyDkTPtlgPQy1lf1R4srrpaUAjJ3Tzd5FY9TwiCXV3lixl+td4mq4Fr66bv49
otvzFG+KsHp575cwiM+czeQAyLDcTOJW7l202dWIBgNvxn9xdT1GfoRHaKmYBicw
0ipBW7siPBsuFXqBeaLPaB4E5c5sunjVlo7oLq5MzJtxcwRYYKaV6BjiKc4Dp7yY
syTWf6y/3DarC3Im49Ozwvrc4Dhh5mezWmYO3evaUOpmwaQ90cc+owGU9LcLTe7I
ikmMQc7X5qBt2VKO3bB8wLsZ/9xlkeqjzzrLv5D4Py8Wp0eYjkY1WnkhYA6CpTEI
nzTUOVaX2rYrzFpjalKvvIzNG7lbYivuUaTcojdjPcjCWsFGAicILQKRupDqiOvJ
nNMZzw8BM1vFmF6OjSr1yBlDqTq/VVvDqYjPqlNzAqwFCiLC2RVJKj5CBajzz8ev
ayWLEmm3dBc7CnO2e1vBiqbG8qzqQSWKuhkm4MoJ8penbxBc0yx5p12DicQaByCd
9ECHff6h0Dvu5Vv5NYGy1QtBrVQ2dtBgWCuT9jElOaRoaZiNBoeJIAuAZIZf6okC
XMX7lgxcGXXhVftoR8xFdLRf8UZfsiL2QKux3dhqiDj89LvvtgvhYQF2Z3ZJ3rtM
GW8L3PNYfR+/MYKasy0Slu4m4h2vG0QDpmDVb8aUrwhQaSn4hcibr6wWJSRrajt2
+rGd6YuUR1xUkyGCUrgD+fOqflYQYuJm+3SLA1HT4IyNVHtDc5DHXtSecyoulFv9
Af0MuH6TkM6FfA+4k0VJUGHvDhjN/njBVrMpn5BT29EsU2pujVveMGITSfX0WkNC
0PB5cYG++4OrCcoQ34J3NtFqngW/1Ljsw7dyxpybaRL677M0jeVT1oD0B9M15Eh1
ZhJXW+wYc/g/30ufXfzXeg5ec/THUYJsivKPDIFv0iBXS5tRTT7e2ufl1W9sDviE
ldm7uDmvTghLlmxrWXIs9T0xUpNpyhv7Mpy3/r5RO/M2tOYw1Ts7WZ5NVou0kb9x
P+fHOGPYYDy669JHkcEBIbVhxT7GgBHcaAvIyv6GIXvRv3b2qN3/d0zoHkdv6vha
56Q5c54i7FkomgvG+A9vPtLv5e/LOn0x3HIU+u3yxAhpNEtJlX+Qnis90ibwA2Hs
pYbBDybOFCUJbcdrfsvhFrAS4vHa++tl1nJ13LOwzDDWD7Fp7Rrvh5okKNnPIgJ4
tCarSH7YxQFSPlRGIRr3cCfwV50guIxyGXtQZNBZvUQ7TOg1TcMu5SbutoMW1SXM
UYyOUzwHuXY1yjqohJJkXG+FkRXKVAmwS4nPVS4WO479VQJK+T4tUj1U1A/yqXk+
agiuLrQY5WNfDNfEb+AB8ziDlV5aqUfMlYIF32zpyyK7fZfJYt6xUwIeMBZq9Jwn
uZKfAjdR9JzvRpC3N+YFTLA0wRYGtGCiKKBorg/kdq0NTsiWiemay52t5PV5SpDx
6Ka7VBvEgKsfXHEc/0uddaPaGuw5Mo8W0LH0LdX0iEBUB0Tu+bRaSXKfROXcNgj5
EZWu1kfiaSbnzIJkK+xcxLfDYmCywkUKWmZq979mEEaP47fSsQ+Ge9Otk2FKurlD
cF8uDeoWaVA0A7gkgrj5B9v+tbOp2JR4PQ5irfdZmHoyRFdsQ+LSYY9l99ilDoNc
hNex9LJXEQQpexVdcywD/y8treWGWLQCRKfklerVU725WPhYGHYISkmbUKb4vIwH
rWmQScepGmwFFT1OOvvOwd398HjqixtMYcTkBuyQzctNVxJ1RSQ6lBV+A8VfOgm1
/pdEucxsHB9of0DD61RReokV4Elr8E3Qi9t6lkiCn0mkzlYcDAVVIIV4Bd3aZRsn
t7PE4v8Kgoy8fpIw5/KFvJxhZh2QJWp1Ov00sMCi/z4I/1EWXIq1WgG7w6sRkzLU
9FQshFpIQyZfn2Q1GRvzOzIlUrH9/hprOiXY0ZxdxNpH7011ozycpFhePM9HvUdu
sxi8qEUr7n3vqH1SaCGKWts1DAuIyv6ZWjLrxrcy1K94ZySjsgEf9tjjtdt8X7XN
udSgfoJdFg/ZWbu8LPGEvbdSt1CneBGbdBASvljWEMGStefl3WgNlb1RpO/bAYk8
hiHoQzR7ZGEZRTWe8Au0Jo9rjMZNAT7LlIqm85K/ITjvdkGZF488Okvf6JGhNu7m
Ctpfx3DEmY1FSBNR38CwBIGgPrQDjQoJImzQ8oGmKLIexPtPRaFmxnAtifWPncsV
Ty7W1pJ77dvWaSZXrhYWqUQ0dTNmfCORo2d+6HR4b0ln4Nj9VfVgalO0KFVy7uY/
nA/GgF1lPsDztW2aIpyFEXBds3wP1/p3LAWdqLFCVOjWpgmRpKhhJwgzOhD5sN5p
WIG4fK1EqT20MYZuH2uz439ZWgrEpf5aNrOX+fPOylYdZSRyWENQNSWK/TJnHE1l
lYHho4PIsZQvrvpXEeTw2NpxrG3rmKUBQs0vVMxpew3mDI4GVn5mY/vrZ48yu+l3
Mzufx8fk12GR0//J6DWr9UXchXcXxsJPLu/8Ppdjvh26dpPCs9qq+dhqXGDsCtnB
6Wqz9HJ3QDso+FfrkZ7g3eeyljJDtgMFb5t3AREHXxBhlYaD0eq/E5s55QtyapWw
IvfYBcmL64hAlS0UBnOGMs+ElNi6g1XX90iW2zdvWgidmsVwMIkYg/GR5p/kHhhj
PVaQmhlUdRabcss1bxyVE3ObN8Y5MxTt//g1XeebK7oxKbVlnwYtoV2tZcSpMc6V
wbSg2FkujaKYNYXqnFWZvMYpY83HvujF0YvwyPsTjlnTywQysKkYjuuVyiI6vPbs
qwnYTfsyw0xxHdwI6HkTui9HwmtK0mtJqZWL308dUmZUHoUc+Do+MF0o7+f257om
4dXr/vFQRyAzY8JHznyPxCvsyNci6OudU++I3Yy2HDOJXSoYkkUCtXbegl9yH9FV
tcYfUKgEvGXmQuKZu9vDQvUc8lpi8qbEeEzWEKxD3yTpwa1rnlFUGq4c5VXbjVCu
+UBP1wODt2gc6rCjVXiqKXwOfZ1URMslYYXq1HrXAlgxuJ1KA+D1yjM1fYFJBHYC
nlS0xyEWtdnwNDIsLsy330TAIPMIWBlpjuEn+w0/abY7NFLgR3YNq7kTn8CjZCDE
MF13FieuenWmc9FyOBtkKvCtQ64VTqcxe4uT5m2zS+q8XD69RCMcCGhe8KxRTC3y
LSa36xZPlO+vGyTI9Si3yiqCkeZntbRJO6FmldzQEof6TNzYovoqwILt8F9wgyiY
A1ui41QKWKv2g2EY3VowDAU3oOIcaKTxkQ6fzP22eMXT1az/+T9rU3sqizfvpCzs
O1f9OaSdkvrpFGrsAvb3C0NmOF3/47osGperlci+ksNvmaFggka/uByzZC9RkHyo
fXDEWm+Oqbu1s4zwJzkybQ2RGLOWKVUxC/8ylojRKcO3+Mwss0Qy1WqBhlwhGT14
lmM0hsZrjma0smtDfFNRy37Gwa+x+b1zGyQHLWrLkC7/Myy5bkm+fiVffAhCQ7hv
ac/1hV6dV87/z2+/FIUAkGmXX/Jnqz4xWuTxXiLmdrmxoAh/q5uCV9GXooYMqi0k
cprgW8cNzXY2idFUZMPSiQzPc8R+j6JW3uJ38LGMjxwxMTp4IOZgXsY4T1n4iFgY
3FB/jD04TA/75O61tMpkzG+8r6N7gAWUZQo3cwo6vDFUHO4aXqO7H7+IBMo5rns7
obZQpwB9fYLchn2+Wuof7O4RjFFy85cKsxX0PHHJxmKghaCiEJjXdsMak03BJB3E
P0EG2S9UapR+xsVpaYq128DZeUA6HyV9SBj/VQHJSpCZ6i5g4LZtPYHfUyRK/Dq0
Lcfw0mgw7YEANoLkP3q5ysitGoAIzQoehBgijHODPgrTF+FNL0BV6pi6C1qco+tE
TCTij44jzhZ/edN4qCWcPkUdN0AG/ZTFQJe3LXaAKTWV1EUbyAyYTvyeTgAsadJM
fczQhmXFFz/4+wocLiiH+UjAOboUsGcVPmXx8XC+GWNGvKFUXXWgDB0WSAS1u1d3
cRLXG5PBrCOC48g3+/YoO7m7QX9teKCqO4QtVZVkrKRX/uZLHOGnod8ybemrcfrr
BFJZ8atvTU4pZ5mBTAQCrETsSKNKRlc9I4Sv50XgKEQdz5iasNRtriiqpCuXGNC8
2VFlW5NZ9CyilC2QXZKJ+jvExLixbXNqEcGK3rlQyIlFAmHWn/LhaGpS8JTP+VW6
b4iRtH4gBVNwe+qD4nuBlIz8X0gHjPalh85xmjaRepKmdwPqrWJckAyZK8nga4Cb
uOfsJ0P2mQxN4kWZtsMh3PSXAfmHJl2Lwl6V27DNkkaATD9xMQHewnlgllcuV5vP
TTknzHmPd69pzCc2vV2dy4sxQ+hq8FaplWQxeabR/xCk8KGuzYklgumxzeouNz6p
5J7E+4e38VeJtdua2v2dtDGYTqEgEHRdwrxcK7xlYszfJGg4rT3W/LcrXhKxs2S8
X8EQtnBD00hjRsSy/8HzDSvroJ5RWNcjm62yYexg4cPV+FTznWzgZcIlbLgOjeXK
UMcbc3829y6CqdVxLmmHbIuWHlwKxYiSTjiOGlKvTfi44h4+3kmbdLiuZmswblGG
bgkWlA7AZejTDxK6KYGWvMGHYyLfJSphCBDoKkN+UdJecmbIoVkoojNyXqaWvhFx
6e7F6SnI9/ZGO/7gbnUxyL05qFD522dYKzC9+7gPQzCC0TASUTcVfgEfRAbARViu
mlTeJsZVFz8wqxlBCm0vWqlA1VCrM3v/fRULpi57x48KChgxPMZtOg8dzE7SPk1n
HCBkdo3PVxIuzR9O44siWWcZMsyLTRuHvtufhl5JxxWXGTQ4RdDAmn+3r90WkVxl
xEzWie5jQex2FML8CTzIGCSysk6nupo6T7g4UqyhYv9CIKxmxD+agC0WaCOmEHV1
wywpJ5JUajN7E8FNw7kQegHD/PxH1AQyoy+PMefjw6VaUcNf1QM0xAGK8aAFSJGS
/5j7nMAeZuBjt+XPLEjoHb8V1u0Pu8naCKA0qoaYRNvNhIIb2rb8vS8kojD/V+I7
HP5iV39+8t34aHrQh3n0ViJLuh14bRR3oGPmETA7wfeAIxrGudAcu5BsLWZfJlDW
E7a7EgJBRVcWz1vpe//bF5W9VxnkK5D1RjBYDJjB+UtODd3ztI3BfPCjkKW+j4tQ
uqaJMcEa58UAJhzzYatV4nHuNDambo8Hm0mpDw/0qcl98xbHI2DQrIHajSTnxmJJ
mN35Ue+KWjaREfpNpnWTaTOl6fz2pDW9nOi0zijNFb3Xm7AbhOlpG77f1OWP3SYW
cBdxLML4laYi9uF3/JYvQjW7oZiSaXuuwbCh4OnrDq6h3bwm8MVLcPQJCnle49R5
4TYIQlnmn9BOgrDxWm5wQTOUofgz6uVBJ0Xog1P+6++dNjYqLQzkmr4tGNa2iJ5b
JH3LRFrPF65QBRA84rIgO4fN1PRTqsXEZpk/OB3lS7MEaKXK8lD92402X7RanZvj
Agbb4pweWrwacd2fx/bTLWISW9olwJ2Q+wCQgjTk0Af+3F4piFt7FM2oYzE0Wxnl
cbq4fHsI/w3uPilT+RxfLWY4RdBmmU2v+/W211PoYzJ4QSM4PJKwlgDhO/Twy2xv
QR1ZazzXg4neqHbVVNuQ4OSTROjDJEjMotB8iXykQXHCMNLmw4IpAa94Jf2+QyOp
yZyaBc5mO0SbYUEhgodwYFONJQKi+4WZRUv7YCkIJhbYJhGJegtutRAjsHYqPsOn
vM91W301Ki20sA9jT3kyD4eeq606kczUBuw2U+K9lpumuLIZylir+PSCsZTdWB7E
6vxX+8Euz7dsBcuzfmv8ULedsoOfPqImLSZFDH7J+29XsrelT5BbW1qnutAtuZZk
aCMXxpdrpwq9IJGykfeGpEiAdiJPgYZXtPEujTOjw5SB1lYFbxr+TM0OuOUYhTEr
iqHiGph3uFyAP8KN20GoZicBaSMkyrfkpEQZ7p9Vgd5pRSmcJlHoEa+KNMYXkK0/
gKUm7ml43DMD8BQCL9aGAB2mSiMryODCSGZyGXbXQN51RjewwKUvbEvMoqI9ilCS
Niov1hibcMUPUcM4gnpI9DFCGRHbUzIgNbVR1kfstTYK8/xDBSYdjyGV3xmtlf+k
iNk5i8WQjNM3918E2BkCTebAMluyPlWcwpQFN40TWDX70EqpqHTGutD1ME30GWBR
Z85mMc1orG5tK0hcyUiDcJvOBCoYLqfKPe4yx5dJKn+xODe4c68uKUrHfhMWvigW
TGfU5YpRpsDc/MeiQ971mppfEsQ3beNKeoqEhFmIWc/KZk4bc90g7LziF4j/LAs9
wXqznPhK7hfxxJnP0U2hU9u3MNXfFMpb8qcMfzRS4CJLfTFi03SxYcYhe1c0ecZ6
Mg95Z9Mps36xeho1FuQm7AxjVYK1eaPcsKamhRAkiQTd0OUT71didkpKtrnl0QyY
qBP6fND6f87DxVKAHpodmPZzac7LwD+m1C9UN2vHTE4StJKM8UF1fQ8IaiGlCShZ
YtGoX6l79gxbEXK1lqTI7gSqPmk8RFOy9UuEJx2iGQid8ORkPDcsdw3sfKE2KWLU
hhVCZ+QsA2IltNb03q+h74GIDAyM3mjexX4faxvuoaVA8NLAx8i4Yxr+L/u63AG7
E8Lrbr/EFlsu08X2LrwJFkZtunDDF+3VBraGi7PHhu4yE1e3LkG/9cTd81MuxSGK
2um8RILvYKVmDYlj09O6mYf8rrAs8toS1R/dPGSp3tFfzHlfmoOAklyX1HCvHUX+
8vDinmDIjBVHXQ98ohZJgimS57mynFMjzws3H9XVsqYL7HneRvfCGcUMy3pXZ2Yc
/K0Ex+YP7bBcPhr0Ss7Yk2eKftqdAPZp0E99H9arKnNmEZjS1WEHeOEDB2gtAenX
q2BJA99KfZfoZxHqTcs6nzfjwtqoMftGCHxqE9vt9xvkwYFZVp/UZevYP3y3/7Kh
jJy+0e4Q7jKc3BL16zJkWlDFG8xnqXm5AX1ro6KQiJXxz9T7KKUC7ay3ZQLjVUlP
UmunI/S9RA82pPZYusMQV+50hSZThnjv0/x/iUMOKW7+Tg4GJP8LQU3sj9P+tj1H
wWcs/W9JMjiF7ozVgcmdlyybDwCSVOue+eg8Ub8NMkQ6bxGR7XTuLCS3SiH6EtL5
gOg08O/YyYTok8EtV+vmVSZVkJD/3BaH84yYjUo0gy43vNKBrpEd1i6Ad2Ml0jib
cFk20VGwuDZqS+T4hlJjvSoqI9TiX+g7fZeta7BROBx08NV0UoahQe4pzaSgYhyJ
93MX308aXZ1vJlhEA8arZkeV47G0oo3arzYSW7bSOrc+8aLcHBp1Er76//AvARtc
ItxtPN3sF2+7JtQYvB9tXuzmnrUS2Lka0EloRW//IFRiv7lRJy67TgUqAM0ECbQV
EPFWeCyWrAkLJn4BZncGlo5pLDqJok4keBb/e4okXQpDE05laAnmvz+7Q7Z5eaOE
FR3DmKIhGc2JUVSG81SuZN+15WWX2CQoC8N7PuHsA9+qVxrtw4kUd3YpIKO1jL1W
/ndjCOAiX7Tjn62meJQpODlOWVZOls7b0/s8LL5qcYjUjxSbLKacI7dW3GgDg18e
CnexPRtuTAVAbtASKBo43TEJAAz8kaWl3l8Bd0/EHymc+3+OLcZmPmR/L5pnEEt9
K/iDPHaHJftZPQzCIxXKwRpwnkXr17epwjAwqy2VDH6k033iE8qwyaNLtHa6h768
LEpVP+BV6WrXhgBxUdijCFrIi8tiVDZTjoFOPiJYQmM+HI1ewnXMnTlkBwCQUzEd
4ntv1iIWld+kV5NKDIyA0TBmONiv41LuELUVraP3vIbyqnY+kDUHrG3aJekUh+0q
vjT+D/HxUCtqWHf+/IIH8XgDw+lobg/mI9X7w7n1p7Gj57EoXDy5kloi52PmJwaE
2AeTjMJLJ2BklpdB/bSJgIhDEaYz37/rG7NILgiwmf11onefMDZ2majKi5+kGOvw
6YL//qb5Zbqhgg+HSSgOQdXfelu+qISgezTyFjhIN22iWTmeQz4NsY4dA93pyQX4
ON4z303v82xmkbwF1Vu7xR8sYgKnlnL8qeiFa8zTF8QMSw79eKastdr2WtHog27v
MFKDaQIl42tW8nWlESdzYRO1vHhHP+fHlFH3c0y9tTaYx+ThnLxWEbTE2+f8Ctc1
B/o/Es2xlOBJNt0s9YJoqZMmw5cQUIMy6Or8LwZL2rzGuMTLca9EBBANW1uQHzZ9
DO4J/Yz39HY7w798rMbxfPu55WNxlb49qabnFlU6z2gV34o4mNYjk/NwqGvtTXOp
IOs4za3tyV2bFKVdqmzq30NMJI31wPMSmtxVw1ydljAI3PU8N2+YQwxaXSXIXFFu
fvzWZ1SIcWTFTcJ19OAxD3KNPD85yk7OU1UedlKzF9cAjd05j6lQuFjMaydo1Oaw
0MwrotBYD8oFL0ZgavmKUYaB637gn2y8WfvUZvhneqlFvDeNTqtHyLzk3QBThgGx
o1aW6hou9zMzw9CCA2aRpCr3btUaNxIpFrmSxym4ah/cQymWpVEpKWIZgwXd1ftu
md2CtKdWlFc12bN6JYBDpxJNtcCvgfsOnSx+f7jSKUWfwQEayn/8RLgO2ntTr9mA
VMREhri5qArpPQwRq8eMiakw4e+zqneUioATUK2NRKYuqbM41PM2iT6KAZQq2OyP
G9m0HnjWTQ0aBRquXm6kQKitx16kXiNLkUCa1WNCVWpF4i/AYxJGo3G/YOInhqE6
6WnoKh2Hp1YtQKDvZxnVMwjERfQ3ztTOTeEhqQBssvpIxKsgquSyqZHIAPlpMu1k
iUPXNGmFiwImxkhlhepaXqwkCrYSClDt/hEo+RFH0o066WwtQWOyqoTf4L6m+rl1
fHrXhm3Shtbl+TxldP1lT3T0ljeqy8bk9tGOQtY3LumIP5lZkCGnEWzlRj8/y8cL
KViJYVRAb23LeSz82HjmEks4ibwwGnHx2siBjE65HLvwChg5+gtW7YUYP2sC2B9G
MOm13v5ATMxtQG/wquZ0m+enaDOkecaUyGeA9tlTuETYJf+PF2omxedA2ZrsFArb
5/0LUMtMmWW4b1z1BhFfI/N4bWRNMck0eGsd6nOrvaF9XaN1LcpOPfppZTPv7lMV
1/3RWJ2IYUh/Mh5a2b0GcSR4wzPWWfqyys0t/0rLnFXnGoxkeaivADz/1uzbizuk
oLWY29CkYX4JJcLesNRFMOB1D4iNisCqjVa89rFBCxgWyEoso/t483Wyik26fb6C
IETP9sBPn0KTyygKT6MKZ1j/z/3iuiDAXC2HDZDG/G00bV9RxmBDH5ZvMOsj4vyk
O6KCUv6nvcQBJ/WrjNPsNam/Q8UFUIbaSzw3KG8h1zqaNEI+94O6Hg+1iwMHu2Ve
LUSF6BbZ60CbrZMVGcA6dG6nze2CmposP86IRGlrgkkHvMf/lQ64J8n7jZb5TXHk
YGholILYX+xukw52d1TWoapF7oIZDildAaJ4+1AUYV2ZuqQv0fncifb0O8eq38FR
NOH1021G6lQ4+Clrd/RZjB1QyRY6E2nOYIoRWAMZotNB7hOhgNMrEuV7LIY20ZOv
RRGd3b0Za4s0+elnJcj+U3o6wGEXaYSnM/3i5BWqhKBLaw4FnRCR2hAncGs/qE+G
xSXrH0dW7ROq0+T01lK3OttfZhI/jCNSxUC9Ipn7fyw1C565aoXLxQGMTN97DJVN
4nPOWmPaktJTZbSF/ww/2Sn4i4iDgEzE0Wc6RtT8/kcQpP6GM1H23Xdv5E1M/KHY
PTklFsoeFPjGHwAwRQIRUiJ1pwf+ZA2gno3Oda7KyN2FAtVNr4LtaraN0IUQolid
simysuVhF1OfiZ8NhMPVnmv3z5+ERoKeqIsH3t5pLnUkA4plmSh5/UCc2HAyGErU
6Rmd90T84W+X7VWaIEq9TMWVZdiuGiqnPx8qeepgfVsA6VugaWLVedBWDbAG8xXb
vWo/IuIQo5x+0nLUfOSoOj9A0wBQ0l9Tk8FaHQ1swm/Q++JHiBnrNTEUF6IkUkWA
EUocRRz0CsY6QCux1JWDwgTcuC7lCnIqfKrDp2Y9QRUFZVjv0sKAliIkzOS5Yq0j
QKu9Gt3eq3NC76b1YmU8nHhYJh1sCHAVgNaBM/O/TyjydtttZ1cxrkWsYqsmCE6m
lbfyyR51Cly+GzVKrNvAkR6VAgXNlTKIYNjUl9kQm3XbdGQTe+XN2M+abwAu1KOJ
ibgY62kLWo/wQzSzstiHoR10f8YbjANRM7huOtQ+E6nUta+/QahxeC7HWWEq99Ky
dq+Kkzg9dkI58goHWuMdE+0FrBRmuvLxgy8hyhk8CGAXm5x37+YD+vKvhrL2kRHG
R3HcwHtAN0HEdtTw2Qwk1WEHNLQgiz+4fgRTt1uVhxWkkchV27Ucjd4fYf7q1Wuj
B8cbTro0eFtG1pu/cm00O5x0Uh3kuTSFZ5KcPNc0tXgwXevswBOQO0w+UC8KJbQe
714QQRiyb6jSCfXxdh7KArSNOlBjr0CGDu2hKSSmBmctksdLVQbUsDLVnsReXEB3
IAjHhcLLXwsD231e9lqqFVqLUY0vbR/Xvu0sBClotGmw/S17VXSoIdtcrQwi4zjO
uB43pwvqSOYxKylOlsd4iIsdoH2pGlLlSj2DpvsDd+pkx4Gd3gbpGbTop/KrRjX1
Km1Usi/f7avY6DsaTqYXZKKC9JeLp6HPrwbXTHI7iaH+IY2PjFaEPxYkEjq8NQH9
R70jXSZqiZ/MwhFyxRCBs8IShkUkvmgDBRnMbxZcffEUiXS20pRffq7rtKEbuVrL
cdxNgLNoWaKYY1uWvghNCtNaz3zctgP0SnLJANvIi8CZBWmDpv1rPBO+COvBYEMg
DUy7INyI3D2fmSTT/akHrwPu9ni8YPnn6BIF+Saqi7H0YUtb6Czx4mI6bFyqCKiz
tBPCmSYofSFv8ZTYX+P7U25nghBh25wsVqkz5vSNwEKcNLv3N7NhrAHRikskY8ez
KOgr0tUAE3oC1jGrj793uTyIed8dJZfeO/enc7Rhz3wRw4XCYRZr1no/ILZhyQaW
Jt6UzDLWweO/3qZt3JonuidEMF6sXAuJUC60Qntww/hZb+JqiHV77scFHYfCB12/
zPmi3YRSXruiYywduAUQk3f4xN36hN/RnWAFGZmg0tuoaiWD5V62tw8BE1HFO1I1
KailJXmiC5aXKt5XIW58YxqkWOX5p1Ry9on+Glw0chXnZFRj/OZnVRPKkLMJMXxM
dvxSb0rwXZ4zL5JX0Ex7ZIeY5wn5IZ1iuUEBs4U1gr1Gtt7qlSFf6h9jEXHDhIT7
nkJGfqDB9F1zIqN7qA+nVl3EqT/x2EkTu3MVzhUrHY8O92mRvI9W0kNFCQSsnn0T
iQNaC0kA/qac21mo9pQ8xsQ6bj1NOOZca+eQciltFX+gG2WwWgxaWLC/FW7UMbqA
ORJvibLYhFT2gl7Kn/8RL1W4ED3VH25MRaW3bUt37azNza6KLzKiqO0SGHqg6Coe
dc/9a4I3TfkqHXEfHkr871zTYfXm/JNFg7xBEFZoX5uzIiOFMm5bKc7SIyBwAjAH
AWtqEfFLayKfalVDFkKqTXyVXA4QrbOiSmTczeebjGrbTzNpu308rgIaOJtisn2q
cIUAfFz/ZBoMVOYhsEHzJoWOuFjdi2zkH2doGFJZyj5SAXxLxMRi+u+RfJ80Hj0D
3KuGBJKdJ1NPhKWQKOJhzGdPDvcWN87pAy78Cl7erQIzxWUKWtKSRxLbFzfOwW7o
qcWWoD39Er3UlfMQgABRY2OBneNd8U7Jq0UUQ/vV0/Pq9to4TmLh7iFMUollF0xH
zBRDTb6TIdqzBVBVsSdLOCnEgFxiE7O8syLHh95/xl1fXoerrpNhtwQrryahL0iY
ukeImdK01MqOUQUYL0sS/KWiGU8GoNkEamo0rM5GTndECN/xv4cDMF4WE1mQH4Gu
8VhBaXodJTy5UqIAI5MfQOCeio69LhQIzS03SOjbGN0ar51lp2YQtu1B80Xncr4b
o8jP7sb4eNd7l1IbSGO1o8pLDUranTq8IkKFRKNM9+SQfBSk5npJYO3qIZ/VuETv
OfXtEo5DB9gFuv4v/2OBKmrIMYeaB6fJTrUpahaL/nVZpb73tpvCL/7Fxw6hx+gj
UwLzQXg6nO6nBrUk3KpcXCpg3vV7cG3uOADIWwk2025F0HwkBAuPqIIqzD0LKvKk
L8zaX8ehjqW4HRVA8G76TSMWF4NM/kj3EqvmFlUufWTREJ/pmUGaFtK9cxbSMS7r
/iQiXnqfNHveRWM2IOoSS7+ePJc8mbEA7R9JKv3NJS46X/J1BVFe/zxw2gR01Qcr
fPsZ+aHy/w6tS3DC0Y/k6vwu5Kur6LipIyc1ndXkfWyq7ly4fDmQJE52Q4E+RwTM
YBpjnLHVaGdGwkzCpJitvzhD4McmjMYqDFdT00uYoX3mAL20v/mYNT3dOfic7+YL
57dXRlOtc0CrG5WBvMusj4TNgY2ua+PMl9jixHLcxU/XuxZN1/7TdTBfuBpDsfLe
5085BWXCJgts3IBc6aKLxkol8wYIpnNtUeAwbTFtEeJB/inxIDBu/etkYQ61wRS5
kncmFKlOKSBgrAulusYVMjl06s84Y/TTiY70jMZsEJr8QLJmOCsxrsByzOUmG9p1
cMdGarx3SvfX7NU4LMZf86p9VE5eIv9Jg9xFCvX+NdlMJw/lcEUsI4xL+69FlFm/
fuy5qA+E3XTmmjj0UaMOqjYabbfFfxJefCaOKfuHoIQ6a9kEwUMAqZ2U6STgejZ2
+LIJFH/ZuUzbR+3K5an0IJbHArxEhMiXvad6nLiZ4ap5v1G/BJva2Gn1H1UtGCgp
Dhh7mmqf86qcdfUgz4+RMjEx8KGPurtnCYeLW4LFgDXq6sxCeC/gWqJPQFPM1Pr+
f1/jyVyJ2Iv/lEkjxBJeyYHlT4oDOAxzEChgiovshIKka3rnQV5Lcrf3r7IDrTYa
WMS4x0BK0CZdCRotTMg/YaKJuPmgmX6PlhMOYnri2SQIHCTbheKfs9OBE9f277Gd
xvU88xYvRUnx1pDZxE5PaueyHh/FpX98R0naXvNkMnRHh2o1n1XVmuAbxjwCnMvE
v2hmWVWoL/MhFGwKRTw1FCVZdiS1twLG1R8G+/T3r+M3mLGTVwaQDJ6mErTI7w9F
0zz2K8avWlLVj/FNbizW67isIhJCx5rBrue/eQ2aK7wRy0X0uNUex7kAvN6jS+t5
7DBibu/Er9pKYRClJcOgb+o9qW33Y3f45p45P3LcUyXld2cRbRJSYs39HCp0UTRX
oxZdMoXISE9jNIdnfK2JEkzkVOYZ1Hr9o2APe8M0C+HXWOxelDLvYp8QjJ45hege
tOag+nLsA4TyHtAEtKpdWHQLTOK58Q6NKJJDkEYLUEY/yVublbP3K93MPMfNQF39
gqxTTTu/IpzlvuOSc5+7AM2odkgnbjYRHzfmBClkCfkK0JnxkW5N6FF5LOm+2gGo
Xm3CBvaUsN6qNPxvu4moTmSUvRMtFjHg54t9r+nxQNIi9Ec5rUKGwSbPxSTZ7CJY
FO3vX9OhZyQ3QarCsBXJlDKrmv6yKgZBW8xgWvB93t7qFZ0YvPqCUxerJY6zjU35
maZwTLB2ECEbg/UBnlzIqpT5hOndhzeajWmgLBti3mjlbppVk77QuYQgs8Ov15JB
XD6ftbMVLDnKbCSsDsTuh2Q5sNtebBa4xPGdQ9wbxGeKm0qeqHMzzBvWnjewYmKo
+qcmPlGE3Y501rR26hHq+IgWIA1V/1qSXOqW4EfuAP/TNrpMO0CME76DkSN6sSOX
Fp8JnxnglQIvloeIjYtat6zLDQ3tcKj068TkFAZ9alozN0hrRGGLZq+j+JLosNaX
vzD8O8o+tLGvELj1g88FwG2AJcCMgUwJ3sMeE0l0rTWU8WTIgujf4vOUflwRVrKp
14MJn4a+gHPVQZ2R9tBe3XthfOVIfhCIpAZ6FOecpnRpxDRRE/s/9Nu/hTHuXA5X
jyy6uzKcmXE7Zm3+po/RBMMXDVp1nXhC7To2CIvnpzq/CQXz3oiPnptOnTv0ty7N
4f+zXMGWO934xvowldvkrB11wXeJcx31/aAWE0nEYxYNOv3q933gXfJdxy4n+FeT
Mu9MZUEUaEm9j16dbuXRRDY8t0pLoIxkkaN7NvfkKGqYtvvMytA8qz5RtcxZcnJX
4U1udLSdA1hopi8j0S/pyfLB2SgOYpwinyQ6Q/AVBYY4nXIAt0cqyYrpBFoDP9sP
humRzmUN76BK+FqXWy9nlih7oDFZtLvY12ZL1xQUTaWAuy6kRcOIovEf/RrY4tYt
/g5JYkdtNMHASQYg1fIy99Uii66XLpeh7zowfyfQGFBPxpeWvNquQrs5tNvye0ko
WHMHE3TKA+0ztfg2HVS8xWCyEVMFAYiCNwuErHz9JGJmIzE/3qSDBHNngkYss5I5
yPf3zHtpZs/VCPZV2lafsYLfIp2RzDwUXnSZEdbiq9vC1OwEOLodLNq9l3hzwZg8
IJtpL8QdMDuZG7CXmpt3EoPAo2WSCIZUs+cxyeZQ+U/IhPZpdvvMbvelIJZFOhuI
EIS6T4CNE5EEvT/4AA/T1SASAEcTNZzNKlDU0B2k2A3h+WRWokI4Q/9u1EebDLYB
aF9/QXTJlWXtU1C3E2QtsEmN2EagbzUbulbEJemZx8thAbSKZhTl2HqV825L6Md3
fP4yuMdMY48fUBdcBxtWDAwsYGthkwatZtq1uXEs15ytLvtojGiX3gx5q8tOV1pt
/ENG+zUdfjSuiyPAnPjEBuvB/b4751Cx/1YNUH30o3fZDUr0MzRQsEMQvfKryNEW
+Vx2zdmkhrptsajuKH5YhKoeVJNX1rUl2fp7OycteqbeBV0HRbC9d7Jm9Gw8w0XG
ZKYbDu+R4MksvKAMRfl/h0kwNOEGZWon9e2Z1BbNmUj1nmsbKGS3hqPa8+Sx7FZK
udR2nFvpQg7Ab4yqmVHUH5zxBUcMIqCbuBDgGEqoSJK7mX+Yme/QlwscEfwKcrIt
ykE08xYYmhljF+itn+uMhCkOiPsHdEQalnKuI5VsqcAJmvXpAEqRMhOxOiZU1FX6
pr3L5j0bxK3XdBVnGVPFIHVFGH4tUGzV0D9Hdg24KCxHvK5gOL6HN2U+eEODa5OC
2te7ngo8YYO1lc01ERcxTI4cmjNjZYE+ocBmB9pdoeuoIIMZpDGgRu3bMFg/hteX
g6nZnOdNcAU58GZkIv9ntBA3JuT6uzikVbDf0wO4qxNW1ZRqbQw2TBxRFCB55jSU
EQq2Ota+7oONkU37O1stZ8/LkbEOAWdnADqCQv6YaLMQjI3rQ4d8PQ2ng/SUn+F4
F2x3CpCDREktjVmhlqVwwR4DTeigUS4avMzqecSceqb9umisJiHlc+4VHiQs1S/w
C0EFyXYvzd+0H9jyb8HoRLlVYQdJDHXW3WdmpjkHjXB9D0sKOoFQwK0jog2lCZXy
Oo0g7HHcLIepbHkke05L+ChXuS7s6HkS56PolQ3K3F3oG02r1MB0ZcSg5fNiPdsJ
xbxqT/t7e0PJgmvn2qiswz5laecQzrHWpa/sqgeMFZYow6UeorH6GeXbo1zWMfMt
b5TA7LPVhnfxx0ZnPTHtryir/SGvKHKd29fG1j+kv6n/q2ked+13N6JlBjKsvrGT
k/kkJUuWACSSlRiLj/up3WHd7xHj2SwZLVTiSoI+0Y+nEm3LdReMxoI5pGCErxmI
Q6RS6d46NRMrVSkVkMcp0z17BitXv7WKDCxjiEb2rQL0F3Qos1RHWekryqRXDkdE
oZXwdbVsMWmPfm0T0i/1cXyRlQHXHJTFHTVPN1hPU/aOgafvFH4dBbPT3HThOX7v
wb3T6X1fS+fLomd6oETBh4DhhaeGbKVTEAIi80gsO62ZQu1bJJSS1ezIjGPp74CL
PLKLmjBPqG4U2h7+3dCPly7MNbBMaoZ3l8OEXZ4j1c51VbtfXOlhvvuP1Y9bWNbr
0V3VVzXqRUdmkJybCf7F5PKCzZ0q50EteLjaSJe57IOHjZbCK98vymF+29WQ3ENA
b8Sm6Nax5iIONcGfJgEYhxnbTascxByi3sKxfL2FJtewkIkCSd3I7Vjvnz58QOix
yE3epN1mnEHXTfjottbU6YiL8f7QVKCq/EqJhdDFw3R0YnTQrvnhGyWfm0vT/ta6
IBX3qVpj9S25AVXGwLqS757Vqy1hbqkRQPicgXEbjVUwmHyZ8w9I4WPis42Kp7yM
Kezx9AbmlEHz/KmBL6tP5RuPLwb2LNc4p1CImeZrauEUAYkey8fhzG9HskqZZmwv
yGbekpe6a36003UjcjYTlMzHBYZcVlnj+1d8K3mTcuSYF7d/YXet4E8SrEqwbcF9
ekWIfwYvWbbkILJ0dAAble6gE6o2g5p2OAgfX48YAnyE1twZj1DMn7n4DKTEM2Ms
kzULyEeziLUTETy4ajA/EYWaNuK2h1OQhAY21GcEae3sqBRwF4zr/llXL7xvcxq8
XfO0caVa1MARuBuYpRCqzrUPWo6UZ4HB50pDYW5u1egfNDC4nMgV83putIP4NO3E
HDhgg7d2CHDLsW9eJy45Yrtm4YGJT2LfB3BaxuG6T+jCJ/RhlgORvmreGYHCr6E+
dVv4d2kvTxJrq7HQYPG+cDCopfvvPQfOkLV17h8Ef5rZtNbOHs5hIkOIbyJuW4GL
BlBJk8B3KfgIXvP6xfSFKGr53dJC6foV1xfFZOv9dd6PVHJqrMunzZyA562M5WMg
Oe6lUF8V5GjpmGMc+HUmJZ3N0BdXeLYZbx4Lp5BOQSZ8+kWkOMnhvqR0a4ZRhSQD
dh+HiMqhGTw2ukXQKIB3IJKzmGHyE3VMpdpqmGxLpW6YfVvgMODlDu6nXWFGM0Tl
uOLQfz2z6PK/lOqgcSzr7C1+H1H1ctCNwveAK3jEKNwskkxqPb5IJmHwrqnl/+0B
uSqNKh8OdnTQbywsU/4dv0cAECoEmjVywyEqU8SXA9+mkn5EtVe0YN5WESQ0zdwv
sbn9MHhonl3FABHCVXVkn16qeRAa2ETIxB2ezgvLrrbe3KK49hGmd+KcZQ75IBi8
9NFnH2OZGjm3gPIvBJJ1t3jreD2fQ9cAlBsWf5keJVxgWQjkgJMMcKjrZGdh8Zww
phLDEXxB465h0504IjJPF+IRsqduMiZbY4oEN+YKdrcjDhQj5MFdfcrLQW7jQ5uL
UeNojsqArsaPxSC/Tv+howOYwCrUmzbqRRtAir0K5q63u+3jKA0tO2Dde4SmTt9V
JfInFuAG7HpTjESaSaxM5fVVA1RKqBSI3Nrq4S+uBImPaM/tJYI8RIcXSmqvxyaE
cLi3D1PEyA21e/MwKJx/Y1enCovcPzfdmAeHPblhxWkONULyNCSnhG3+FdqQFef8
CTQ7H2FrjHlZSBi1MCalgLsq42xXOMj9ZA8ib7rTTGM64j0gUT0I8zRHxEFIXyft
MJBKJ1Qmr7QrkghyeTpG5zb7NCznszAVuAHyKhqOVozKB9gRteLyHSxGrDHh5qlz
eL1nKo5mJj7CJC7WN49b3E+BM8lbrWzzAW7kie+Erj4+rXkAHlcec88YKQSr6CQc
z2ZFxcPSepiCWPENuIM6nel/fEZegoe9JhiNUrYWirJ2pdwJOrzmk7DdUyn9bkq2
ZRarD1Jxx+C9xpKZE/m4wvXdsbcUCC++PQBFPMFzjr9rGHvMx7zDpo6qrBAXdfML
ujGOogcNYQmN+/heHA+hfqOiyMoNNotpX98Knj6kx/AZU9S/oE//R+3L0t3SRBup
ySafcw5iJbTBIqFeCJB2gmJukwVaUpWKMWrFqK7SmYxqYalQgQSjakc0SvzEu+j3
XacZMFQOTzd+lneyMA5E0mvl1SrrWrX1Yd1LsYAl9Izu5b/0Plz0KyUG+ws2RP90
NfKrjhcBUOqG26472vts4CerL3Lzmyop/STJPP9JlpVEzHvfXfHAuPfWIas8Gr5M
Fgfu8xXde9hC/TtkXG/ztyCk/TN7TIaYFqyihVBVUQb3fGxJ/H6dGpA6FUbFV+vW
yKiEkTSEDIptgHT9t3wXl/zJNnLqMGqpMM+Poq1rFi4cyp/HrT+jsHwxVuqWbjhk
xIuDZJNcLbAQwqAcv9f6YjYpZJAI/Rs5C4uyKhIrdZOBFneWs8iSIrF59eTF3qu3
Zf9XY6yhY4wM7rk+GW2XuWqa9AScyj/SyRsmPZw/SSjW35tE8j1I/KCIpaydu3+h
xLbdpwNSqW1AWSihqwhSdUMGXnIcuqXH2oKWKEbMXyS5oXu7cBbi9uzzPQ2YuO5Z
wtgxZz8V1g3o/bkd0126ZiivGTMwcZ7nyzh+4a4+3x3OEYM3ze5CDJ/42lXOLGdS
vlRbU8ieW+MJkoK4i0mn0J3Dy0rIM2e5UrtEvENMKHolnyXD8WCYqFVePhAPKrM8
5W3JuAPZiJ8dWu7EVmu28N/YBhNK1TL67Il+NNmq6JoyIz4E6h8AXIf9DLIYcceq
Fx9Vt6vknfceNyZ+Xl1d9i8CQr9hILBgZrzhaU7IDZPaQoCC+3hFw9oz64g1+0yM
nQymwgaeOibI0Y6Lsm1GVP+86VAY+U4KiBe1xhd0OE2tnm9646fTbEqusxZOIujh
lzuOvZS/rcmV8CVIb1LGYgvFZ97A6EoqgfmP/aZHl5S+sMmY5rMAsmZ7IDqZx8M5
GKbblVEjJ2D71cmkhhjeEiBlR5FM/LJpbznhY6ENXh1YLqrQdqO44ChGvtFE3bsv
MH38UTN4wKhZQ/Pvs73xArtjPRNY/XurdibB867pdCUgZc46ZfNDRK+NnWXFZwzJ
S5IIZFeCgmthLLxqipkVMpN6ZeUxZ+ma21Oj35Q1Rp/fTJtGnyQUqIJY1vyeco27
U4yF0vzuJuvloNQz+31MN2ISx/GVjaUGTkXSoZooCFZfpo5dFli40/Smxh8luRFO
pBkigG6AVGG8NytCRb2CvEu6vmobZSoRIHqkD/gIFq3Y/m6kn3Z5cFuq98+V5kac
ab3H1XuYYmI3NTdhIUL8pHa1ocqA/M9GdstNgT5qSR8kKiKZaz2P/hNU72TEHAk7
ZjJpd0YHl4PS8L1dBcHrwlfIMSGSt2dVO/kzNZ7F5iL6dDBWaSZR2O+/aQlET6Er
9kmQxcH0N7PN/sMhXldxtJdy3YXg5UZXQC+vnAV1nsaHOY/02mL2pd2QyMjcemGz
fNQZQAfAcni6Glm9DS8zZ81XkMG1Dg4Oiu3nUoJpucM0I9+36IUvl894lmNz50o5
FajaOWWheDPc24kmQvoC0USnZTmm2QV6iU1v79iXGHQoMZ/ki+9r16Q5ZRRTJYb3
2VyZ6N7IRhcDkdtzkMIQt8zc8mpoAfqnMVo6ssO5/5RL1DDlwvi/NJ17sPiYe8Dw
mMHIKcjuA3ppuk6leHJFEe9qF993LjE1jv4Jlr4vwqHpGVlsxg+NsooC4dZon80W
zCsHigwZ1XiTNTTVFrdEn8mKSLnudxYE7O9y18QBlxIW2kKbS+bFjcQ57Hkiu0j9
mDLkmG0214NaSkxenuB7Fx5uUYHPfp/5fMFxETnJdbnJYDO3nLrNW5+4xv71KL/n
OXxC4AquDoRKpn5ud0VzG/bcdXwoGCWc9YiCI89qJ07OAVonhHF7lqXgqIe1nsCp
+YEMnVA6KrvW8eOT+cc6hsQkoLNFixwALoHf5jKBlMWUvLLmX8ElCs5s343yFh4l
ilLmQUga8AnzTpgYq7HGFcCy1B5amFNyuRENu2ejaUKmM22aMr9xxEDJz6XeHcdi
MimOCEbN4jKDvIc9MlArvajTiNBP6yt48lJSX5X5IN0iUPqXFC4dZcBUpDm+01aw
Q/pBj13JG7coupfLFCmYs/iAZgMSmiL2igOcUigarF1E2C+KL9Myb4m5TVxJBJtc
B1O/rH61OmcykQThqnLJqVvuPtEKEveeS4GkhbwNmLtUhaa8LhOioXZbEwyM2hPX
Vqaar7xUZB/7M8VtsnUkieG/T7GzoncI4BbK1xlvQo+zZazrAK5i5+x13HatOEVd
YNOVUxA2wuE4kMhM0q8iJ85PfHFgBboLj1TtUtyKEry0FhoRAL3ZAIIbh1b+JcY4
mALZYMtYMMYCw4eLmudlYA+jMPbymkUf04mvNO+k5oNMt63TPA7nZ5Ha1d0S2FrG
EpYVi5uwB19/m780MHBiEufJqBEJsmkPCxApX0NB6SnwyP6Sl+4gXbZxTSnuaWKw
O0gsZuFisLz5of3Cyd/nXWXBw4uVlGc8iGz4h6VMqRsgPgnLDBB2VRL3lOABI/R2
pIRaZ86PlXMgJcPxq1GP1oEaVoFXlD32/STIGGhrmt4asnUxzInxy8q4b7WEER0r
PGd4sLXKyMmLI96ekpUBSgTD/JYCwYjnVQ5XPKpi3vAXOqCZCwzx9qm+MdeZBS/Z
s7Znp7jZBOJU3M436wnjz6qvhNayTwFSP+cvxALwe+z8c4gR1GHJxF3QU3j4VNXl
5SpT1AOVPMnFEj4TD/dfMyFwRNoaUTiZzeEBSj+T/1dIr2Bo5qbRKfla/gXzE5a2
0gyeFV60eQQ7LwAtot0+XQvsZ1ElpT6P45W4r35xRrZJ23kZ34JHDQnRvTc8shVY
zHAZvXFXIQAusdLHINMt7cRyk4ImMOrq466bhocgkxaq/hAcU43s+ulZpKKKST/Q
nwBRvB4TN8hAUOYVMM9UXM9CCIogNj1i9Jc+iMlBgUhInSYJeyZu8SpeXe+f1d06
IlP4d/xMtCq73CMFf3SGyhnoWVQqt+DN3467KAl586rq5/M+dllKHa+INJYiOwX+
thVF3mHopJKN6pyVLa2EP7Xw6JthrmfCMZ1dqPWSycThzzU2roa2NwiCP0u5fy72
99VJiBLspenTqeQBNW2x+CZsa60nssz8WYEPTMzXtt11EZRDoYI/I+b5PcrI8xCJ
4Oa9ta5YruZBRmOLZQsmeSvb+sPfLendQsHHh9F/379H6SZJfQecU/9EBtw3NPny
PYIxQSopCe9iioxWPYSgPL4rpkhM0Yjqiqk+ZnzeuMpoP1rlm8H0LMl/EV55IBRh
pDDLcxsfcpqop/kx58koxSBfUonXzl5Wf+j3HpZDg6jU8bUthwQO+t+hUmeOXrZd
w6PAHveZg3vDCmyFKuXvEpz41H3YtLgrzGjiV/C9u+psjrXnFSndcLE45MfQY1tA
0TceuasyYJMYrrgGggRaOU7GGvwSon42M3NtXgrxdLCBNCdZJrUwujIPJb4te9DH
1f1xQPHpCE9YuXGLfRxjPCHpzQQR7t4zmL6JHT1kE05oRdL9CKw3KzWal6z1a1SH
nAtSt98olkvP28qx/q9vMTJe7gY3sw8gazrtuh1G1Ch8RxLv0XG+w7jjWGVb4m/9
mgM7DXCPYmpdRzxXwc3zBajWemxlIJp8QyIEKBztuRdyeES4nXla3GXtMAaBtisX
CwIqbFtTWL+qZ/pGZhiM5SZ2M8Y7j8sRHTQ/3KcoGY0Geqkwxki/B+blMKR9NQT5
7hTj8rhheP/objOLhiQ4LqjpqfQzTsUI+04mWOB/Lb89ORXtbdFrG1VyXIsZqUTt
fBEPl5s+XQO49eRqgwfXcUCVJD/O5eZtQQdS0T8qKM6mdOnFeGAQ3ChIkmwjcnkm
OyHN10L0bRw3Xl18yn4y0ZTS6P4yTxs2jul7k/4vzc4yWdt//RL8eGU3blgOvEDI
eOUnI9oCe80aaXqubIeYFZKl+atm+QqWZHVwZDqejtHD8boFcJwrm0mG0BhdDMzc
JOWZu1YUf/FWzBzDn0gFMVxEDn5hRxaaBYWC3ddAXkC4sVr77MOK6j00IVQqn4jQ
TsFqEDklUeZy3+E/aChJ6rUByySKOSbj1QNsmCIvEke54LdqbKQXijd905j0tyCn
IRoDqzriF7nn8B/qJNetHgIRz1JmP2m0Zxiyq0f6sWkCR2c4FWzid87xpmBIlg+J
MzT61K+fS+w5awFaUb7frKgZrHd+QY0LmXTBL6tMQhFj3Iy+HGKlMRlf4X/6aEw3
gcjQAje3WXjlUE6MQQW51gJJ5E0zzaQKTbTSaKXrG+SdYW/8Ert4SPnyHX96rEoa
/hdtecc6X7EFpme5dmGQ/+edLBk4Zj6kAKZMzmSyr3mntmk3nB30WbAxiP5s3J0V
OlbkCDYuhqGUMd7uYq/ONXFweupuH5G546sExyPkXd0VJ6OeCLa/+gqvEhGBT9YD
yyAffErcs8DY7NBTKtZtz0YM2B0QKvSrw0e+SjjQLWPXOcQ0LUVeAM4aOXiWkyMx
RkEHzBFg2QYxvpbN+2n+6xqRdXjzd9ODz4Tf7BVbg9NamMfsAXHn2vpXyyoIbSM5
roKhEmwdAaIOa1AjJLBEMbyNesXY1xM8F4JoJWq3SilxKjCcqsy8TIcugaDVsBSc
/xIX4rvhAOmu9Ej4UOVoR2st5DoJMVJk9n3W1zAD8/c2787j+zMvYId4WD92pXUn
W1UkklBjcUvjAX7qs8M8rpPTjIn9h/i38QbRZKW2bp7p3akV6gxTPk6mXGCdeY9r
SWbt5E4MkFQWsREEsRVV/diVQvd8bjzOzbo1BXLqIT3mRRuUs/qg5ltu7ieoLZgo
Az/3OcDmjHkNdvTL6PY5peH+Ji92FD1lgnthEj2Cb0FcmQDIqUtFcQfhUykFJdY9
wAmYBIsTQdlL3FYGu24DHv7GrlHkImDzIfGobmqYr6NmUilhiX1yLJTmouNGQeFm
3ec4J+qv1CQxcS3jcrrDi98L9Uo5GDojeK8iuZu5j8nk3C7xDFkDAmigUeAf00gE
a1LpsTmCsZFRa90P1gFBB1GCY0lgFINdGVyGoxIXbjnVTJ5eB+1zMsH55cVpjDaf
+nWG5Ku+pJLJSwTh1gxvPefGSTdR23DaTdNHT1NqfeYeihHXlHgyBUF1zolr7c8n
JGTqZ5m7829HgtwsUKaU7uDS2qBjoPZEdxDEcbzGcUAzJZfw08DpJoLDpSDKlwsq
HPhK08geqyWmIMP5UQJ36NggpKVoIcVVe5BkjHmlySu22+BEUfRYr76HQHqkKcwL
xiAx055CinMgFheSCSSvFvDCrIhGwukTxhzOFfHvIFipB79BYTuOW9yD0kO3AV3o
kS1fTLIyBM2RETOQiMSNxPpiqQjpPN1yvh116EcZipqLKLtUXtxyk7///Iym9Vpu
fnVMAT5ZayaOBljflWJ/z9OfkpAbIewMuHUZhGOj4jutELobsqnTMKQ4MVFBRaeT
nDxejIXfI2/p9ZeiAgXraGUD4ig3JEYaWhLd+rUV2jJXdcPgQDaBgBRw6ITI/3g9
M6FtWGe3MCIo6Peub+Y+XNHuGxmr4DGclpG54R+cLtyzvqNg0lCGC1k2jRDFsfmz
BLn8W7KnT3Xp0EjPphJJW2Zw+eEn5K9VboTsa2OAoYMGlqv5MOe9YL2YOMc+edGP
onatWkypAF84YU484lyt7w4K6HE+JawfW6cqt3+N+bMz4ZnA/UAgv1OJO6NJftiG
HX5I+XdGPtGe6q8Aqiiwq0KQmuuym3no3DkJAyoaHZP5mgpN1eoBmH5i9Jo4byYO
KgtoeM2fysj0nAAzjxTSroe88sNzrcUdB6BF7l7FzDdQ7VcjYj7wp3OPaWYGi2Qg
Li8Oej3xosmeaUXhujAEopxMtdxDUKs81yLTt/ee2iERghyhs3l4LqDtRFZB8kCv
1fskdkcegUTjnvZ1314BOsPnjfcceJDBcbLTcr3AjZt4kcY6bznJvRHbBmPxLFyX
MbxsbStgJmDyIjmboRuDwpA03HVntb1aT7TOyS2HpJfJG+gvDPYj2MJozbWpMrhI
uQi0a9xNsgc9jZLBjEyL5T1M6eF+p4/1KQoUcvSM2GTrNF1D64CffYCPG98GyrU3
b6KmlvL2NGU9JAagWbJyg4fBdCrJ8V//b2jEFlYDVHQb4a6RQErcGcHgcpAQ+y2V
XjTEaZG+LNdcn+iN0kEjGpfH6/Omz3/web8Dpiy5+3kaVJTeQmvoWQH5QkWKR+zY
kB62N2hAxA35DgpjlD7CYx8pJoAAYersceLgTBK0usbUnNG0ivwfq5jZ7LJ4Uvu0
ss4B7DD4haRHar88vbvxcCIDM4PMeqGCmqZ5lGW/f8czMf59lFBa1gIcgC/GdVcH
hGbPCEMMDrFar7UICnJ753xjNuJE75WuP9XgEplfUjkR2Ko9hOuylsY4sDtsD9U9
fmoxBr5xOsfUEkCtcAkhLeRAnBJ/6OahP1tQ7rw6ZP4/t4m17HSR/I6MZF9H3X/p
Alxf7jwB8S2A1O6DK5hy8cek/NwGDe8v7ATVmAa6akgYHI9ODBnSYDP6D039669k
iUaQrshE3V1AwoCuGpQ+Wx1pwHEFOg6WCM3Ve0GzHFW5J7/YB1fYEmtoH0AKa/ja
YYlh8Z93jfPZ/Oar97VzQualtNx21LWKZbMVkJhlEavik7dlarX7winhePOAR8W3
yfKzsSiR6iNf7geTlH1RfPN78XEAez//5PHifiw7NLyhVL1LvWeif4R6VPt8Of2h
fIXLYkDdNV3lyOE7orl1NZyQd7ZE8GfRiEZcGI+hYSPNUbUwS86har9sOQjarWQ7
KvCk/J+u6rZQ2ocfqKEfVIau9TnXobFbwu4I6NAB1MOrUQCEoPLdZBQpcjq6zxOo
alluhlK8gYAVB+tT3rdxQNwoNg5eMYpL5+Skbo2Yikr6hcv1hrWU6wpBL/XB7uSi
qOryVxQjp3DQ2VdkJ6kxzICvIqF98q5LrKX3n2C4kXiIDQ5amG53kp5l9fEFm9iE
ZdTuNnAM9bEDtNvqCD+AyVfnhMd/tLcp2J556QsNJHrdNmCeXkWPiy4K+O1gVkVT
mhhOHr2xkMdCVlMV+hBJn8zxogQOpetc3S8M9GgoKfTbcKEPMljZGmUqzHVWHbAs
nZX6KqvI/OyBRuy060VOmWqU9POM2YoTsJbv9VLZWJ1fi+EHYo8vMaaV0eb7WT5u
n2xTLsj17+rJk+YyF5paby0Iciu7lxxuqq6fWzUntX3ZAbfulvUYXVNCN4S1V8iG
uX8MjZVspV+3Z7SGIdmjW7KF2BJDmHSE2uTqmhL6cMz+7Xp874YPgLC1Xtt0vNWc
PrdZ10CqCYlyM45FfD6r2Ceyhb1hYRvKP3u/RTRhd16RhbOXmwnH4nIQ1jfjFyUJ
hVdREnuJEoy/g1kI4umqJ+a9xQiDhD4ktlQ/f6krS0xWDpos6ykVBJ9s2GvuUMeo
VefOORvX058yyG3jsvRnab1LSViqLefwtDQVI39zage2ExRR/hbIlJnGlVGIkWD6
2lIu79cpIcmhFUysF6FflYPiCsAu3j4M0092sewPYX84wgbWWnn0th8/a1R0z1ec
/tpzz/I0RmP8ribrYUgr8gokogwQ0UAHZThm0B9u7xbkZVKufurAaxRiVEwavNqQ
aF1KBLO2f/x1xkJ2OlMfK8Cig+2CIreCV48a104EDdkd+qNtcHJTOMX7BZJebqWq
Dxcs2NdwUJqc5maCNucBcuZPaUb13tQW1U2GWQJ0T4zq4z8ePNI+9ERGNs7gSib4
4W3vhkrsjFmferH5H8Ci2LSRZZ/zzuntioYGdofOasS1CSDeybjK6gUMLgwFDF/b
T0zlRXiMCkgImvXIzFXtR5cSlylKUma9sc5lts7+TgqBWPJfhus5ZBaqrDe9IpLZ
aFXCo76ym0ZofCB+S13U79sxbNOWVphJ/vLHp/BfijIpQD8hbNYJiosJGT0owQhV
cnjqqcXFi1N8S+/V2aYRiIrP12cHdq5pvOBqOM6qytQFH/wJQCh+VdpuOQr1IJNd
vr5riwSTLKhKEBKCUYu5HDc/A+C81h9H1+hxSLdz2dU9P6op1+xhs78eiSdBeBcR
jKwxz2Zf46jM3//0vsCTWAr/nx0V2Nc4xqDHpDzGLsSVmubrWl02Nn9EqtcjqwxO
xnXHcaU5+AF/mRl5FGIc45pJBmE5KgGEZJ3HSXoCbI4y7WAFJdDCcNP+uMtinPvT
N4xft6ORi/KZf4/n0eyaz2A6mZc4pBBb2BFm66O1e+yV9rlXa28V6o+hzbsV0dfH
5ssKdjVDKoyxU/OuMdlw0O90y5RUzV8lQciywtzmtH+u8virOhioMnRSpEvN6oLj
ULbQto8t09xRhma6V+oJzG1gHusQ3gOGaD1zhkHidDhC7GiFkak427de3JyO3urS
bFjAOd7gRxKQ7ldE5D1EXCc9BtFww3u+Ypk/A0XwU87yyIVHzsAEM8Irgf/n2fUp
B2x1pBWhlUqlGQzjJ9ZIFSSr8O9hpVZZ1/Jv+ELq3H3EcGgN4BzrFgkbP+4W3Tt0
Po84MCU2oL6qzjrbnCW5b1MbwZylvqpRWZjre3VXTItH7GBfeh5tE+6oZbO2PaWq
sUElzFw6u4MH6K2MQTRVx6z0wyXjAhjxLkJ7MHLZWv/ERsJao99cWEau7c2vQfIh
oDq2g2qFvFC6LUUUr6cLwiW1XeCRUW/hIlwi2vc3vafqmOkj/S81MJqDc+LLH6Lx
LDaTeQaS0lcp4nm4miHfrF6QTgAsPZQmOYYm/EgTI9uf5JxgOb8jPsScUUQ/OciM
BWsYlQNC7zVd4oVS7n/uHPmz0XZ2/gegSmJanP5DtGFyFUCjz8dPC3J1K0lh9IgY
weecBjRZORnW8gY6y++18S+QiWRH2NuBBSLVu2soeF8aPLydXnebuaMkeh7O8lLj
75D6ykmG7YkNHQaPA3DbPZIbEbBO1lTVAFqBORjcPuDdStbdGDGRg+E6qXNntzKp
ia2mIeQsZU1MNLE5b3T4gtBBkaiu4neeaGYpK79Mmq/gdPgh7HNF3tCMfQuYlR9U
+Y1Zp4NN+zQwdr8OnG21xxmEp77J+YRnrc9CDkfDkm80eYh5ihgS3GbTn5Gap8WH
NDEdGnUNzhqEtT8Tn7vfZTBwQtHHOdHHeCxZpkGcpv+uV2nqc6xba3M3cuBr0I+n
HeZ0QkPBzpJx2WVi1Am58wNVhnZaxGTjFxUMBg5K6+EMC/H/Zs8Y7tmxNInD8su9
HhUbjpZ53Gz1y//207eKfiakCYaFjuRH8CLWYgaM1i/62U4O+KWkA4bEQZ9BrCCA
vKK2xC/0Y6E0/6MIZMi5mhlg+Eb1TTkM+3cJ23FahASsLKQh7aN2w4oHmA68XakS
uWaT8wO3ZOrbIZOjvj26uivE/8z6+eTxvw09lb5rzNltUHdbWypRmugeN0J9oB3B
OAnqNuuC5qceqhTMe8GwRHaYe+mO9Y0Cs+kt6WyrUhebdYE+/l+tT9iWuSC+AemU
NrNf1soPZ1NfWllFDJ5/f2Xq0D23faKtmkt/SxOIX473yZvp86SLX4ZL0V/MSWyR
tg+ay+oPBkuGUHLkIqcDg7ZreaC89bssEpQMLAPX2z8aApodfbR7GMhkfp0OamQu
DFEcCORHF9+Q6mFjz4gIl5X51JrEaz+VBnmNHzGqMYed74tbLF8Rv2gG1lxoA4Zz
8sDhQEOjdCkYEUfCXqxGb17n2ngbVEby6Ha1Q7tbGr1l4TIzzXxTmzMdt2jlKtz8
BMp4hOBmxLqNdE1m8FomZ96ZmO5lmTpPMb2/BsZ/VDloSGe02SB2B50B+2PmVcPM
btmKfab5yK8xRUb+7gqQohBzzvZMqs7TkuU4/un/bZt6dwALMD2+WtsXguGWqfQX
XNg6nMq1JYxjqhlIQUtyWlxAapFjzfwqTpyntio4yOAET5sk/RJLnYrMPqkl/L6g
kiq1mij3q1oWF/5Aw0+uHUDziHUQku09eBjr76ak9EJg+U7Sq8/bQJN1xpCsTQeO
X0V8wUs7Yy00KchrmNjvGyhpBQ3rLZ/snrOGalmS78veGNMdWIaqVYzYsHkELUor
ChUE9/UjSTaOrTeImIfxjVH5ON8YxxuuUvyf6OttZ/HvDLsLbMmXVSVv6c2Cx5do
okypiSZZcdvJWySO5vuDYSZtQBQqDHRwe7n+R3Bmd0QY8alwOol7KAwUwQV+ZMeq
rDxRPUsfgJ3i0SN7kZ3pLnk30M4cWdbgkH1boCQgBeufox+42nsk4QXuOz/gWIp1
t7Rs/fgFt5fSBcTOHkLX8m13CcdUBTsqzjHO0NC1msaQct+ht+NW6j/sq6niIbRG
hwrYBaeBpzlT2jSa31TzhtgOMadopQyqnaURgeD0JBm8XH3k8CKhMX3Duv+Dizwl
UL/d0Zm4Xc7PaVtb2SkV3zxirU5awBcL6UxU3HVApSW5z6cTOvHv3R179/JK9fVE
Tgqt2KWQSCcY0WgASXxwzCDunig2jGwe/E0ewMHQV3elxF507TFz49lGh2D98uRD
QUCwj4L890MZfcjDjFCD2+96ptmWsmUMLw0Kkb/uQMLfRSF+/VhfY7bYqEeReV6S
Nen4VfczByejiZpIJKBjGp/KmCKa9WLFQfYdTU8tRhor2nkodz2LEoOYKhv1ZRyf
lzNraVWisGK09UEb4PP9s8wNX8Tn3e52UywQUbmSOEtCtPXz83rH//7R57bKvTRU
AjhOP3C71Rqosq7mwAyLSCTOIZS3BJWBRymLhOOtnub+FIVWLBwKZGPtIPu8WxpE
U+bHNn9L7xixYkWSMyym8f3MSHNtIeeuLquDuRHvmOsayaLEsi/PKo8ARKW0Kbyw
cmy91S2O0lPkexpVBIs+ebGtSHtC+Jmv/IDAiEOQ/ZioQ9A8JqXA/C0XvUixStFR
CqVTUHmouCu+5qthMK97qntoQEcP+6qUmHLyRmvP9mlnFugonMEvgiFetk4TGgak
QXYZc186vTQYgkvFnu/nlJzkvV7QyCqVYDrPyr//dEqeXyiEV2rupGL2kEZhipu2
LLT5IYyIUojvMYhWIsDFDEGcoC2By1vWNFc0sMVqDqERJ9JHpz/v7IbudEqe9hlz
suiaD306SoiVftS8PP4RNoOg/NbfZANazn8Asdpf2ZwRKsGRzG5ldVEcFMRZEoxW
6be+ujWJPPhbAHwuQ2kPbzI2wz2PJUtDh3+G0eXVDesqKYCNo3d4P5DtTofci/YJ
UsFNu7mcoXgPW6HGmtgcM2cn7kgzvJeqIaujW65pYbMUNDfDwf829jMPf/+57EW6
oFl9YjoaOcKAPu9edZHYZ6884S78IWePTN9KgNZZ93ZQpMXNtj5Cj6POLZ3Z+AEp
FCRKMViZfaAXF23rpmGUty7/9yI79/We2i6MJ6XDUnHVOl0sYC3BHQ3DPVEyBRPw
/9AGmNhYQ5XwKZNJRwrPlWWmek1WjpZQgqGe/yu9OmqTlwlhyXHrU/wetYeUGSYg
+ngFxbtTxajL7YZwL6eTUbrTBZDOCs8xO2zXTmKvPcdMcqSLwJ+f6fXFmpH8ae/3
YuGXV3DZgx3BUt2MtHMbeycLNAdO+37dEvpCwbGtk1NzwLdL3zpOiTC3+A1ZOkqD
YSTnNcB8TY5j7GDJLFbqMtx3xpugvVS6cvW3FnYJin4wnrI3pTVbWaV7bbMHU9DN
YJv6Vk+ovy3omgaDaWcyBTWCNiwvnERv1ZAVP0NHs35Z6XjzsT+/Jo5ikgIa71s2
b/MG2Gf671s/GmdO9vPiJ/jQiScrUKW8e9wrkAufYxuk8oZlYdhAv/yX3Vfh57Ai
LXXpUvPFAtR6b9nFQGs/rjyPLD/SlsZHyt0vNB4r95kJU6HBARdO/Ks0krl1V8Mz
AK36lB0BUxx7j1gKZxtXLoPli+JwyaCmac7KXa9/pEi1w5THfuIsFg4CkrYe0z/H
gapN0RvaAcGcOgYE9d24xXAjquSyxcJCUhq9KaUy0x9zVO5uCtuX66L7XNi51tup
E9ImqufUWs5ntTb1Bps3MRieab/5eG4b0t9O7xwbUuxsJFSn9dyDobi6X30iyhbv
fNB2fFYsns7N52dMLikV2zRIplP91McYW210H1GGxFnVybVZcSjlGPq13NezOHjf
BVSKXtrsvcDf+yQEUiELHwdbXuzzFEOiB9QZZzDFz1Rfry4tOF49IF0sgLlQNkcA
PVQBlwrIZG2hR0jRcKWysYyytEUfFWwyBYA0h3tgx3QUq3Ts3pQI/DyOj1D1eMdc
p/kR9+vks62oHyZ1G/9AyOQAe2DrnB+hC61aWajdAtwCQtB9xP+//Bmb6dMrmspa
r7sWcsI+/G1wEQXt7QyE+W2BgwdVV+ekYHctY+WKxR44aaNELIHvJiwG5+okff4O
u1vNgeM0vvNb7ASry98bfjYkFr/wx+7Jkof9tX5sUGfcFaj7HRNCQLYtEmbkj5+F
Ppx1tJxxNnVtDEGdLfe1oxjNTKTPiQxxwHM5uUCXqLUdmbNnNfNMNEy275Q72p71
uxkjO2HVLhjO+oG3Zb0JVWaxWNSQWVfNKNvBh514ajhYZUfXrjfR3mlXkOLEFaUo
/wMP4pMz/xOgP5MHbYtAp66XsD3aKC/E2cnzCwZxZCW39Pm+RlswI11Na9ihl3z/
prkxqlHpD627vwRWzE2L50m4PDyewsPZorJuSmcN6PVyQDJaBd76UsF1W3D94Cqm
5OVNCgk9Lg7boUNj0q8/aHRzEUUwf8Yo/YPgrIUmHkUNno2lH4wgY2Md/ciENaLw
2nH7IiacxDYIGKH28f1UaharrEQLXcKedrytdjMDUQCTnVtbluA2kO3s7mHqPoq9
WkGMK0oAlffclBehYa4kruX9bLTfU+/biWEpv7U7sn1JrjziKTlFIC13KARxk1Pm
JcHBUrJaA8iP9bCOW4AdB/vZsbckdsXLHPRNZve05ZEHsbtbUcV72MgzjgjKyvv3
oU0RgyVTI1kQoO0NMBTuwwRiraBEvoF7mPsNCKeq1ZOfzkZPIv80Dkre1VYRrC8a
I2tLujKJCe79avkUVgaVsAR7VEYkoOeetnR8JX2m+zJjC9az+Tbm/wFmDLSDrWP1
aDFJCh7CU4c1XnKl+Hpoj+qjL/brGPyjQegeMVvPCoiKKUyRwizjY67s0RIw3C+9
WGZ7KzAuJ9xYSjmYYH+E95b+1K3m6WkjsNI5mEeUrfsUqsjw/cclYSeAit0AniLK
761mP7maJYOEa/Ws8FqZKGZQkVL+5nFru0SsxSmjBuCSYx+jyQSw11+wDJpgjNjN
NxMQA+BD4dgPj0e0KrnY1yMSjhhz+iPTvhVGANe2CEUjJgZ07p4ZC5+4hxGkQ5YP
1ADlhDGRG+D2QxSk+dY6v65+okQ0Rg4MT3aqQgT9clX+/+3z8mUVQzQaQZ4a1u3h
OkWb/O4UcO303F3fjtbCC5DXkuP+1VumrhexHfet/lTSOkHzB9/9DOWoGd21ovyt
PBP0DSv3vddrimoWu20iOr4rT/sb60Fh8MbNMgg72d3xSKhDC3HLaiDAdYlrRG6X
QrR+rJreGtVAhVvp19mk/F/53u5ovKVc9bqP3NVg2Ja3HbGBS4ptnX7gKoa1NR8S
I7S0Xz156k83blP32i6+sUNyKKkcVxPNUNTgrJmj5aqEXf5GSa9OT1ZUyiGJDlBH
SNtXwlzl0rmEYF2qz1yjEBjQaf7P4sgDueXOA3NDsxV/TBSPWdu0Z7jfN2V7zUpW
BiO03HxieDBh/QkoDOuDwD8Ndsax0Yw6Q2hpmEIN9XrpZQAHtAVCxYwFXt3n/4IN
MpYgkLMwAVmc5lUUCYKhC87jnN6ATqlHAfORDTGlc79SJT4jDslntOfrEWJQUq4o
Y1Gy46hdajh9rKO7ZXxWhLHmCp0nsndOOBnpQr8gAH0IF46zecl40/0JsRpDiE+F
bBTBCcedsD4M9UPnRX5akCSNVw6+qiDsykqD2mzLTCQWwd1itHQGVP6fguIoD3lq
+CQggErNiPx8+f6lQQaeHm1gJxxmZisFZP/0Zz6w76UavJ2wd3AQ9qS1i3IJlZh6
9a8m8RaRHPlSpE78/u4h5+ugkRvdTuCaTspxqqTLsFl8QdT7jshpPwXgjKF12Vq1
4Ny5yyJNS9owE80P7QX0qLX2KNO7h/V4wEvROJLu8jBN9WGCJ47e+5bQg6gbAuSh
wCKn6sWDhMkG1CH8k/h4D+bdpps1cgWAGQneUamgphlXRZqWkqouwrmmG2sAh1Jk
5Po6MhNFnI3CzZE8rXPLeE89UFE7lYXZZ6MNMrqNrVdmmxZ2FwqMfH9gvJbw64g0
HLiWbkltRqkU3o6m+xGRUdLJ95m/1xjoQp0XWMzzMcCbcW9Fl5phQ0J+gtYGa26e
SB87z1TsCWx+6R5wan9yz9WfQ2SV2cHUk33FoSJGIMKqBPsMBMYQb7a/lR6veNo2
mRzj2p+Bulsm/c/CmgXNhXfoGdGrS5BN3F/4gZlSIDFJmFuSqpWOL04PXD2iqnmP
1c509iZCKQdQ9srFs2F0MZ9TpXm0adfV3FfAyZAr1Okdv6vlbfuyemBaq7KL80UV
QdKV+W1cpR7IoTWDGw7poRju8TFBUM74YxlxxcojikXWFoaY3C44zu2/WQTlA9Tw
H2p6ROW+4uJSdU9bVUmWiEPtfBPpUVnYjgZKoF4UXXgzV1z3+JgZvq/u3KQxq20c
OYG6dZ8q1Lc6aXgLwJvjgnlKQxj1d0XigMOAxsyiB+oGwyrtwKFP97i/By4caC8B
rUBQrYLV9E8VmcYrsAK7fnK/uUelTvgCciTzLZwdtrR4eQq8BsNg1RmZmoq1EUjm
O1GfY60WVw015xKATJmYZAjX0oNAwHIWEXRj5EL4MGaPsRNcAXtTlb9njhniY9vE
HGnDobub6qY4v37RcnouMAhNXLrvmyhVQWgriCySUhFck23A0R4M7yda2j6QOlzX
hyonqB1gsAc7DD40j3cbWlLnuE4LzmQ/KSx9y0vKTbAB3Y31ODvvgZK6VDeGNfJ4
MqleSddJT+O1uDpt0YIfm3KQ+I50roxw84nY0rrf1iJRgr57rgj2K3TPD5DYQlpa
pmeWkcm+AXFWAtO6Kt56s47KU+uoNf9OyJE8Gp+il66wBLe4y+kanGmj84ixcWTI
YOD/MXUIZTqq8S8MsKs4bBKXXbgrmm5R9uQm6YBY6DTPaQzLyR+KTsPUeDMWEfwK
o2LO8XiU/3W9pMofCEaI61ccXMfPaTA7brTz5cTIQt62iMEgxeqI+ZKZASe4Eue+
DH8HguUrXypL0a4fdDuA8Ybv7DnVGnaq1CNQqdeY17piovGEYhfYAM7JF8v2DmEH
6RflfUN7taw72RsjZ1wZPTTAcBvoy51lPhh/eWLK7QulO7Zs1e03nmZwcra+MTgY
N8ytFOXtJv/P3Jke+0im+i6f0/jli0yVjjGDonMH1rOM38O0AVvQovO+VbtxmAO1
ePaOiUwPCCIzFR7F3rkM/W9+vqt+vNIapW/eTQPoCwmEX6kDcro7oEYnigeHMVun
jlr1eV7/AvAhHuLrHmuWfPjlxHPRn0BSMTbJjg/Dgf0zufEdhRvHe+9e1NHczW42
Y9m9CiIegMsqSE85qcCDBVtYWVjLThF0Ll1+RxxD3RD7ecYszJs3EW5jNLFk4hSb
I5QLycrJbq+uPjKJNCjfxRtjk0o+kvL5RjTi2aksa3zheuVFnuJC2AtTY1HsKzEJ
cnT1RPPmh5aEuL6HaB0t0Ebj2jKfEWG1m5luNZmuHRjxn2w403iZS7TvgOLhdAzk
KHDc/c6n7hVu9xdRU7IeqL71vtT6T2cxd24ox/wgysB0f2F0xWlWbkMWqjvPWTzF
MLS0PFeYlkK6sQy+pF82VtX+RHqGVeKkvueyh/oikUoPzHby10p5HvW2JS7AtqOf
rf76+9kb+NaevNKYEnk0S2LMje2g6EDmsER4r/pH383lWhMt8yLC6WnhM4pTzpnq
ojeTZ22hDiwmWNkEdWoVxX2eUtOEmtvRAeQYmIKJPSMVvKqN3Ote4LTLJdcOwZ/c
knzj5Oy2TgqgthX/JV7olBnzvPUIf9xqWgEzCXfLn1Ru8dqbgw+MbIBeWmgUi3gU
rbfKQTkOV87++F7EOZ2RVnINjY14xCN6qqQ7zu25BNVCOAwKaKT++zi/MkOFQ9Ww
ZamrrtXx+yrApyDmaEw5SXXbDjJiev/uR+w6nC0kVnT2/ntxdVnynk1H4REkmz4D
RQWG9gSFFdUzqGU0mB7lTTSBjX19DG5EiDxww8DSDezrjiQD9dI+4rAhcx20Iu0D
MRFD991JEqEZXmkU63MiWf89VtjNw+sTLXrDPkZN5ym7+MvKnErInSlrfEGGAq8S
XTwWlX5/irWo+WG/ua/8vT7FH714V2G1M94wmBIbiGeELZRqoakHsC0titkT1vUX
6pJrUlqPDI7OseBUMdvLRDua3EZWGonCs0IGoJyiH+ILnUb29J/boBHF0mUoAjny
dd9oNzZTc7oHuAAEmQJ1KcFTNtVoDgs7+dOCRv1oontpTx73RbcgA7CeU14WPVRW
K73i95PolnyyeHczc3DNApucLvUDbzGyC4r5Tf7mthAYouDF4o0QQ1gcCC98SSjc
QS6MaQM8bqX8Dtm/ngvGBLmn3AeEkK8eJwqh+lu0wWmjf7LIiKINcOps1ofhXbV6
t2ez6Z+XyXeXIUMqSDHoSg1PL0OuGRPiwND5hXS44jvGcfYlMPyvlGaeJMbY1qUa
YXIVPsP0n9o/d0zIH+WxCxqXC8rNjjmYsZ9ZzTF4tzcpUcPWDEgBxL//dvyUhmQ1
qBBdNWnYH4WQBf1zY6iqUQOoGydvz0lZ5sBLzVpFN+tfjydu2WYtRViidx2X7UV7
c/LOEuJD6sfsUmQvKXVrqt1YrrD6P3zVErqr9ENl0xnuayczLxIXJ90kozOnHvln
wxaVrHKt98ZMwUxBN5LZbbvuK/OwpXdKYIq35v8VQb8YC9z7hoJIFL3Om+wLj0x6
7T3zPNhVFP9V8g2I7sk0lDftPSYmV1uXQwp/egzPWOAGBqlyfpIA/aUvfR0s3hFs
RsphdilBb1RvqZi06x+xEQ0SAh5tFmsySB4jhRf7zMdW3sRuimNepGHQxmjBFm8p
pRTKe6velyHxBXVwx1dOAqYMFHlT+bhMl9ET8zi2GrZBNpMxbZPh2KCWMuROyeES
FPPv3anuhB1mMlMTTdYadM5EwPmoTR+Q8lb12yYazKULzDP/ME9YJk/a0z9hCRao
wXkWdFmvpDytadEAPraouSLqddsGaN4xMu10iIq65gE5gXR7PORzPN5pUJyh2IZv
o3FO1u1bnZrNgPMKCTXFR9sX115YjLqLQTDMVhDGea+fVt+nF4XIT7sZ9l/Yb4sb
gsHo5rQ12SyHcG+ptBd7zU55RhON5ASZWL6l+fj+edfmHbR6fuEXZWVtv7ApQxf1
/8UkxrUl22OUwgG5hArGprPI6qFN9MhEQjTUSgoKpHXXs01lPu8GgRARasrJGP5s
wrGF6g8YGj7gHvk3pmji6sTL1IG5czzXVPO44poePV1FoOXArB8Rz4XZvuFIFDHF
80Ox7AMGpqMDM0J607hbuWE5vQ5mV6+PMffcDpiwkxKnca927RmBLJnTA4jF/Lk/
V3YFVGstI9ViHq17FQAfsL05QV7cReNKz/xr4ANVskRng0lQgDDtUp+xPaV8qnFt
JlL1q1Br2xny1zFUdcdPMImaAYBEQB5vMEp0THVgqN6vlI6BLloy8WPStFicWi+B
m62nj3DTLgJyXAT8Llf7xYja8TWDkuXghVPaFxYDe+tq2aCD87nGCQTJH2yUaTRX
r9nZHkEAW/C3Ws9XzOaK8pnApWfj0a4scoqRLLumwfvNasvq5ctd9/lpHH98o0Pe
LjtI1MLNWF2G3f0Yavu1cNxIWZhdS8H0G5efXin8o5P98DFEVVdu//Tk5ScLh9Lg
WiyMlwoEGuZ2Uti6k8/5bPIQR3H7oFDbgKhLdAyY9Z+J5ZV7OMLD+xklqYDUU4+J
BWxtz36PheDSGWZDrQslby4I6upwrcejvyzhyW2jiKm/9CaZEePeGE5Pqx20hEPY
oAM22jzh9sOUmRNoy9sQxumwAPV7dkQRnTtQYixes261u4CZt/7a6P5T2EtD/wFW
4ng3QZRjP3ZmcJEQ5e3uRnA6NT1YgayVWk7iRtZikLGPw+vgQ/yYMRCgDNP90wez
lDj/Bi+l04+jnu7y21GzVZZzPLgGLdLg8cuD//FYYFeGYTztqs8GZRYinsAHobOi
AI177nC7Q3dnwJ1oVLktwXvGp2C2rv6f/zUPfUGL/cLbDh21140CcmhTwPOIeDSl
rlTyPYbS8qfHVysNn8MPlMJ9GgaMuNO6LZHC220nSkk2iEKAki9aJkV6H+Zwb3O4
UL6cGYVkka7QGIsM8SJ6Kpzn2vwzD2eZ/TcPYJS6ShlKPlpzB+lnaEhfIt79aBoL
Rbb2hEt6eJM3v7GTnvh7zXqCAwcI0grLqFJdJXzjmZwpH11xYR9pf6yRSTwdJaKV
PksJULLpZxjTyHd7Q3NgLDNFvCwTateNCH3tWf2wqx/SB5xgW8gSxSvu9oMiDoBT
gM8i51wxsSOxV6tElLM6AYsJy2xWR0RHA61oCnHiQGGH2AzMG7Vd/lQRlIR++61+
Jg5oGfx6U40M8xUqEdeUjrKend/MusMY4GM7XJMYK/2D4mdpiNhCki5r8uXHK8ib
XZH6tf+86yeghpGNuFoLr4rJWJCrbpYTcyRQqRRNUL8HGBWfv4kQEp/ayXwZ27Ag
R3Wg2cvjFBytAPvW1mV5Op5A+snREDttdX3e54udj5+efTSV9dgREywnMZa39iFx
NEcQY/3M753ccfLVLlsFsGIr9hgYg5oxIejr41WwZUnG9/ivY6vuP6uUz1DpumDV
hOqG7iA/c44XP085Og1Gh+CkhTcKCglaJh2SCngueRHtM4jIEBGZiz+ma1e1VmIj
xdQyy8iw9uG2qL4pvdFELFogljN52CsrNxsoXE3OdQ0+jt9QXLL51uS3Usy1f1t8
B0p/i1jiuDRV6sqBrSX0PnBmWkpbs/YTFvyCNJRVhvZRvN224Ei6MnGrkDMVEO1f
tgcQyLZyWsyX9+ksSdclJCGVGffdNXLuRUiC0v+DafbtHzsMUEvqik+VcNoof2IF
eTLRC+Ra4GQeJbS3BtksuGd1yCZxgdUtpmdjBU+d1s9kPLt4NZmpUrY+jYeOuSzq
c0lPPeUBLjyEWkpSOvg6zxh1Ozx3+ifxvYpIxsTmxDx0TQqBY6+MlqWy+omQu3Kd
wHC0cnkuc5y/aKKqiMEKMtqy0G90shMX/2ICxPwBBYuQMcgCvfr6klPgpmYFOtD9
mp9Q3z9SujBK9g545Y3/1mhlPTffbrNFLnt8ZRn27PcOrgOi4/QBVGOizZbrR/mJ
YCrQ2jVFLhjxOKBdBFl+3tvIlxAnj1NuuaEQi/h37tfxnshS/UsbFigkt6zgSCW+
B/RkWCQwKPR2AifevZI1zazlv9dDStIMlrE2Lf6IDhUGWkaYCFANoSqz2X1GVn8k
xXcqxg/HbxvBVGJ0LHGCVCeZvxYXeOZz9fC2lGR0UmRmfoAtISmw1PyCCvdNSHpq
F1aSgjrdpVb1PwIcMIzByKwonZ7MA5ko3l1FJGBhPyAsmzJRLzMYqNrrDNaZQ9Hj
k/3iVpm4FPOppi0mQDDplP8Z5JkGnmEvXfKojLI6s0Y/W7ZSdLKF4w9uPbvbG57P
MI82QVZfTrqABT5QdswcDRg5nUmsFDzlEufU0jMcJA/n3NOoI1a1jZcu4ahGbQ/n
tzb/sStw/zI/6EY1lTQWmU62MKTy8J6scrhi7KPnEYUziadVDLiwh0aKRThNnzVq
7bJe+BjjRGHszJIA8Tic1eYi/odVAjHJvK85Cs39gjjkfQS1kdyyzXRUpgCgFECW
Ss7WiATzRTVXuc4wO9PBx9DKkhmnn3GdWCNYQN7E/XPNbWvJbSYigvVE5S4+W0o7
4VwhXjRpWdU0U9J/HFZwOPEjRaczK2kzLlq8vOq+cPAg+jpVlz2YskdPCJOMXuzN
Gzb4xkgae1GVGWEJMwV8GgcE5Zaeh7zvK6bnbQN+Nwxxw1Ra92/j16B1bo1UyWFx
b8fokFwFwsEECe2PnSToG+C7d/3JF4u5SGewhmnnKm+j6+FbvUFTl2Qu6SEPlVr3
fi4h9J4H2Lgc9tsMP34mhPUQUcHfRIhU6dcW3IVT5CH9avRTUNwZ7uvAj+hBNThk
gFVccBfq/r95axN9QU96yri7Bz1gKstwLTJ+S6o5xo6z/lS/la32FkyaTkQDNAaj
LNySntL2NwyUhwuTcvu4r3GahTDuSmMNl3r5MDoLkkBkD+pvgah86wuUfrj036l5
QyjkFLlXHv2lCwXKJKbBQ49VtTfse2SWpX2DXMyItELenzsPhsOzoAZ+UaDzNfGJ
qBf16+9pOI2oQzA3Ty5VKpnJCwpjTLjFlwnQrzI7NpQcuacO0ql41nbRmEDOLHiM
nBwAbjHEHdZt00y87QXDwyG+su+LF2i1SmmtEn/EztgS52FB8FQQBCZKmEqvVwhl
nZb9x5MbDt0/c33ZFLEolWUKwkcO1r12khuKUEYajiRZhrblzPvqMl3DkGd5qHA/
SsEILtVYUB7QpTjq2sXDDVj+guYvciUK1GTze9xj6kUtj3t8T+JaTjL/kMqo5ZIT
OegjMEWLl7b2XHQxH1r7thsePA8doO8HEoF+lHtA6qGV6GgEK/NSEFb8t61K5p4Z
HmKIwgdRzjaytrVWEVxEzpiDB1PqE1jiFN3sQdth4MeJfk/v6xv1RBnVYntwXfCu
e0RQbk9UckrvXtO7ijcPmHsLFuyClXCkenuGSKaPuoo6fC0DFxBied7Imx1auyE6
WZLI/6FFkpLv/53/N+n5dO2zh2uEod7tueJ/g+JteB3tBdhdVz4vSDIjnSVjUndw
zQFcRzWpvGqoE92VPf5w6OCnsBAvtJEREnUDvo7GR0WG6fil9CyXuRG7Ru0aTzz0
YlplpTxXCv1itDHcVKXSjukJek7f2Ator6UF1loU3PcqF4KEeJjOt3J8liugh6kN
mXPdEEl3SYjkZypqFrDOiPBEuGhJjvh7X3+vao61+UEnccS9/zlLtSd9/pMAN66W
LL1ywQFar8v9ObWCgSVHDnKlyNSI0vY6/vUPpnYQA2l5DOIi1kLk9jO3KWd6SnB6
bkOvUPyuPJD6Zxt4hS4VR+lCsztV47PbMVFquC2QJSY58qXOn3DjeA7a1CVcDJWk
DIgOtiRQJONXDUQvHDKYEqHJQ6reZtGrcYiPkeFObhhbjxO/rJLQX715tWeb29QK
wgmyXjvTlmto/07+ORFwnj1r9613MhNObsaE7Y7b4DKubawwNxcVlCmg6YoF7o5W
3ypHGXr0hZf0qGQyn9MT8jdBGgu2EeiTkzmj0zCh+XTPy7Gik7/afyrb1QMZij+1
DCIn6eE5E/nfeUWiEvDDtYayrcSPRmdvdBG7Txc7WCEITRDk744FcaVaHVJP9ZFZ
OMCbNIU2ucUUl2VDQ92RI61GJRmYbtwRgupE5aZrbWJuoA4l1AR6q3mHIYYcJ5IB
OzbWKr58/RWmF+i7LpJU/+YbwgGZuJiITTldMGxPS3EGbIB4np+HRxNyS3QA/vHb
mF1z3UYdH+pYy1KY4HoeU9OPFrzxQm4DXlz5WjmHKVJerYCd2xlbAFA17jq6IcmZ
Pk28ofPBqmlGomPQ3OIzDH1ihWXEVrEd3YXfmfa+v9UwdoDtgRLhXDyW0fc6NBKm
ZaKqD4nhLuooZp5bOxHq66rGpt04Gxk7Hi6XUVV11gbEoZZNhk7r5QyWC0dGZAH8
HjFYTB82PgqGTUtoPc21P4HaYZLqZMzoLNA7m532/U3WxhYXYGmFb3hL2fs5moTr
q7/iW+wo3ZyalL6tqxIdBogUd8mleZL1A8XLXVllDYoTFFQ/7ISi5L6VBqqrS6fa
zojmpqCpDUqcC0Irv1vDMVtiFxD4S8zGYD0WdzLF9GbT4/QM/lAkXM9bodlkcYP/
cUqTquoqGcTTiBeC3WZqIDqcpgonD+VnSVCKdvEjb7ehfKxtgyxrLAYRHeexyibc
CC6LJjoSyjeN0VzJTDTe1hQlV9IaEVeb0B1X2vwtLcy8Ucdmp7cfD74yEJV8wS47
HQRNpmnLh0nqxTgmZ6U7BlYtnKZEXYBd1zdwBsmNN176OGNw9uOEjtfKUbpG1O/8
Y0aBLuxzhA3OAziSvAemu7CPa4qZcOYf2rvUJl1k05mMk5Bol0V4STL+GDFENvRS
sTRTfqvr1NafFIsApBEo/CR2t2WV4MTOFqldRtiNiFMdf/dfomW0xISolDGI690W
EiRU5icJXX0Yif5hCgD663fffBLB1mt5wQoJizW71FRPf+ZcsyhwLtdZzUBNMvwb
xfb+5vWMNOKoo2SW/eotYpiW7MgIUqQFhZZy/APaz3aKSQlaU9wWWJ7SmU+U+2ko
ciimrCPyCH+e3EjTg/2p5YXuiI1b9kGi56ZnU/5ku5gKi/Y3Od9Pkv4tgGVpr6pz
ij7kI1B2P2A5xR7oygyoOrl3+rGB1R0YNmW/kmWn61r9GSE29XosMX91yXf7XtCa
Bp6T01KnzdNqeUHyN+OY4LqPxOgAeGuOMOtocZN8EjpUN9iviyAWshFYJvLXmOV5
pZuHZ9btz/KxvUZNtr8xoUS1asjlytl9kYiEbOQ7aHTcscqrfglDxS8iUZofLuIA
lq/fWX9sqTkh5XqEA828Pbwxb3AgNoxIuNz2+pT2jTvMCAwXEuLb7vVXZQwHsH6l
4JIM5I1OEThpzMfk3HnM8xJHP/oiRDBNz4iRs95WMCRjU/v/0kXJiajsl/hDTVJ6
IgnU5uudA/Ft6n3rSWa15ql9ywx2q8DLeOP3A9BI3SKGEJ8QoI7ul4g/wLQqevOk
VoNf9gyuKRD7yrkWwcwuGLY5VkYxx/BAWJIAA24vnHTKsE7Fb8WI4HflaE2Dv5Hg
s66X06ooHif/YGYKNWXwbldeKAbFbAOKUNvzSeviq+MClNTMSqGf3kMi7whYSSiz
JScYcKysQN+o+n78/+nAYql/lWV0oM1B07rJrLSudfu3dQBvYcCv1qSWkKLbDRle
610ySUnaohqZ3MZGTDgVWLhVrQid6/XFv40diaMJD9VsTzwtAcLo6RDsEwbWYQRG
JOrPokUq5iaFcTGCJ2q4UxtoWm7TqyV80fdbvq/a4Qjga3bOXCwirbCN6+xtr9wD
oOxdx46UMb5WWwkAn9iT2wWQR7kbgtYzfw3B5QjCxOGPODq6S5/Z0N6fVWFyvwLr
u4BB7nQXVIm3kuHIERU2gpR0txdn77V9cJluaWyghscXULPptsxJ9cAYK3+ZjPSy
YfvdLrIDAAS1ecZQSaHv+Cv4oxky6aY2572KFLauS+U/LmfDvuH6j/YB29vzw4Nt
mSlKcBekJdBXfgOXHEi1QnI+fKCnY/izqvAnWqSwwLwGS/LaG2omZHokRwhabGTV
snET0IVYb3V9xT82dj5XYXAdXOs++BIAl3bwumP3TeIsb5diI6lcPppd143NzgS5
mJpea8eJRep5rlgWNwn/1w6EVtnb5atG8MSOiBPAe7vskUW6+bb9y3Be4hM8fCIr
Q0i2b1X6dLuSa80qrgVooYkAR7MTFihFRuTCzDoTHosUssuuNOg9b2nBZFujajwV
MWOIF6Ixkktf1e6OynSodtXBc30Fpj+MAgxmO3zoYCHL1+1hAkiuBOLHBrmDRwK7
h9mv3txOeY6WL60Eh3D/a+xPAZzp6GlYSz+MrXOhkcA/44jr724RqmEobBtWAxuR
6bVFtWMfmJRQZ8L3hyPG10D27CffYj4Noqx/D7DEDxtqbBfNzjeEIPw7oZUGfYbj
10I4CLsNBQr9BjpG2N8W6uPrPy+7z093qkBdYUGt04/TD1ggzk0BBb5kcljTquzX
MBPVfmn/BiLI11AY3Q4QPveLP62R2O3L/Qj01GlkEtGHZPocAU/mBTxXcI88HQA0
iFlQokYOzKGNqcj+7WsZZi0kKlYJ/v3m3l0VUof6HEqFiDg1ybbbbi/YbqWAms4U
ZGG3aZo+j74RZjRGvPvF/qxQTE2WMTr3BhFbY1/hKO3E/CtZi3rrHkFjPx2i2kjh
YEzDwntnAzqY5YfqpNmrTv2jaO3LFkiUd3tpOXUVHlDQZzxAdA4Ysf1e7sOplvK+
AVCSXUWz5XL8tITIXgKn82/lpF5kh7ytwOlb6cMB+LpdSLHtMIKOkJh7dATN+034
eocba7DCzvFop/r8F5R0kibHOGpaTwISFbr4TTvf9i3BgydOCQQu32BUVfwAn/Fq
s6q/iP0I1T1qCJj7/fEgKfQfa9wjjVlBq+vSHu2mbYofaCyZ29FsfkcqgTyhtMM0
RBkluR5CakzJrvI0xuhjzhj6SwEoHww4ZM2Y4hDZIePzTYKzFrhXE99ywfAFAj3V
/O1n6GiUEw+8WltDVzgoA0aT36GyT2mu0nh10rqRCzXbzE6d0G5rtXzUcQF25W+n
jaR57lf+k4L179WRkyQsu+8h9PY///6XI1LpwjwiuK6FteYaBD2qbrFdqq8RqT7H
S4umtOQJalQ1iTnlqatHLm+/Wxc8+P8FweXqc4d36uQjv8Tz/mhPIZ6k7t4B0rDJ
iganS3Uzi2Pg3xdeUA+B4qfwLnYv1fV6ezKLzNyPSX42qZkF0VKaM1jYSSuYGiez
GgAu1lhtoT+HJ8c5DY1V/BHhGosbGIahYruHRDU/Zn+/WUbJ8TYv7cscNaNo9z7+
zkFU/9nAbqL5Sh82zsd/+1gGcNODYN3n0lTSEARalBj1ySkLSIDDCawXpNS/SkpM
w8J6x9wzIbmLDvTrs/sfuycHVo94eFEA0Y7cIhAfvWJsA44w/maL+06ThH/LFYRo
1wQeBjibqUtSAJqSctW5aKP4dHcX7vFjZWdS5QYpY7iBQPPWR19UcRZhf0HQ7mjO
gSGyg3FIhhxdqds+i33CmSAdmK+a9GYmrDcmykyzXqjwC6LFsdyvT5I+YS2VtiO0
YZDa2ew/FuPbN1nN5CGbBdFP4gx0G3RHrugLmeusWRcoy+3sepRQlB41Biw6RRIu
yg0eU+ym7F77b/NqLgGaBZ2vo5/2HUKnnIrk5NIw4A+7QKz8QiO6fZI83S3VN+k+
h1pciCBxMavDhoPWXqSeIsL1Unhk4gXND+WGXPNlYa7oAqNGRaC/tLwFvNT2qrfi
93j4yo0iqhYwDZBgf92Urcdd6NydkJVTLqxJ0U9+Ap1AcCo/3TLZEdbTDJZk7COv
QtcD/zMsrpAkxSp/CyCnmgZftU8iDzmWlJLruTKcxGnUIk7hj6M9bEYOHnJNftI6
XXiA+knRk56dqqCInDWgAcPptX6huJVoWwLWBMD+cjG3vT1zl+I83AijXs49MNpP
BUDOcXk8X8NHYpk+O1ur6RpZbo9attALsLBCUtUswsIDCLv0C866dQYs0+w7Toz+
J5ACORgMvd+su0Z151oSmhdyufbTyTicw/T+Z8GkqyatziR7OYTUrxWy8mVy2jfI
IALfmEWYQqKZHq2L2vPCMtS0/UuCo0wNiuwyYN+76mXrb6njecfHKhQQ7sPl6Rio
pcFZRXnhkeqOBiUZ/NgjxcwJaYoQIuLT4AS+abMlCSMu0nFGhXmmdxsKobQU/O8S
jRmJd2yKov1uXciG+z4FEEYJgChHENgVcsjO59csKXWGlA6v1voYOiD5WgY5qJ9g
cF387eLEZAQbkvL6S4caTjqlnshR1AhD/0jYIZb6trpq5khA98TFe7WAR7RYuMci
/mYutqw6eXTNBDCgyZR9mBWv/PGLoUuCBJVeu/fADEtLK+JM01DSx03VnX1tKkby
2legjutVAs8gUbq/Noluwwc6wHE3A3Aha1qISuzyyKIio5QkQMl4U48UxCRoA0aj
DAPM4kYStnmvVjXe8bq2SAv1mrK3SizqScOSO/wW1GsFOIUIA2M/A9cg54wqEoGQ
TD0RaRykg6b+aU6Hg9L7z/Y8RK8/uMsboG4616KsdOEG18DADL15XJegVKpRkrQ7
nnA/IVPy0z7il7wFQp04fe0sFgxiKHfByHjPptF/WLxidcnc+hIoS0NX1Fm5fsLx
0Du7i/W/7msO03iwLqcDi1u03CDOjKaJlq2aChVta9bCanyxrK86DbQ0WWfR3zSC
qk9aywWpK+9z4zWLmYuQ+EZvhgRZItRIG33Ju6heFX5QEMAqdt8keQLrVCCc2wol
WbmXD2wMPU1Qh2nYlMo5/izZRs8w5RF5ZMYDcWzzQ6krHwtZrfVpT1WcN/cw94pr
2CXdnJ/i792FuMl4xTflrYm0GuJujtZ5j4aTnxgkkRlz25uKcHWUhf84ftB//Dx3
jqc9Hh/Y38cxAkQornjYXQyd4yFd6SBr8/2grgHISCqi9kp1HQHcyy19/CJRnXPE
Sy1QJDg+zl/dTfgfegwDrOhyKfHLApqmqjIlOggyqtmh6E0+pOZFIq3R6AKLzf6y
lcQrsKigBGntFMbjfRbvdlT9RojkASeE5eR53UpkZdPHxcLpw/6nj0dNTBBbo7gY
5P3Y3SAP4KjJVP67by9t5QlS2okl2+QtflvTdFBftKwdKduP/VI6emnXnLXja4cr
yhYaBhgiSXj2lB3Nbo1lNR1JsA7dQ5bbXbAXZdJoa1IiLJuBzfJyEUNe5NI+iX+S
uzNQMLfEeyIyzdN710Byzc8leFFduwrasuDQYRMFFx/9JTi0PHYEewP48X3UeA6F
TWZfu71RWvEN++GTnWwmFgwvPdP3HzXi1J9rWZIfD9JTsOvsRncwZO5ATgYHKsay
1pxkac/Xdn0CVHVlPj1Q75AeRoj10wvrD/hlKi1J290oipLO7szXLVUdLTsLlJ5E
/zSJBbEW+XdBKBfPoBr3LrSPENycBZ+e866sADwvG7nTIpQga0tsGnox5hTKna4d
wvTTggnbNYB9BO7mo0k/Rqsaksz4THeMgSoBZlA2/4ztWzmO0h9KEAqvHQch2gI3
MGN/nAKBD0jar8+nIYlrhXKInDdFd+uWLSwCW25bsBDjHyduLYqe1ieWDQVJsBKV
BObZILHyHpLz75KpMGJzzhdAmW6fGdC5z7qjdOG1S5jFf7FMiEWGrfbQlo7PeOA1
8klfy1PRA+tMfLeY5z371SOwwh0E613z0DgGgs+zUxdgXEIAA+5VaxmBsPVEoEM4
KiTB7705cnif0Lrptn+fTxAcXGhqM05+xAafyWdomKFpw4ZxJRurAVCiySlwosCI
qnzwqu0C62K/ItPq83qEfwhQ7mkvkNRGZqsCj32CyOC/dpwUoho1uXg9UCXa36jf
zgCUybKww+6+uRg05BYe4aMMxEtDcySbai6Umlpe+qEx1438pqac9qdgyPSAEI97
ULmUZrsqxfGmsUcGE+7tKk8iqcOMV3CJZEQ2H23g+yz0g+YpgShk8lpfBCY4pTIJ
gPOvW9fRBT/IxAh5tWXzCnJxJGDecFRypZzqyV2FVRZaPYbVIntNgJaJxXRJuSP+
vU5AM9WfGW74R1ZmADCL9E7aWvpYCleDJSYt+8yT1if+rrR5D9OpyQM2Qk7wMNYE
nd0LOtS3xhy+cjn3BxRKZEKczfxuOKv3LGtl7I3M4FQ+K8W6rQLggIG6GA2RaHL8
LnIY+MABUsRjUqrhMoZOWRp0cdJuKnDPgQ2e3TQ8Zac/bDQ1MRHrznDwP5TRyVBx
cjliViON7z9he1TD3YhRcYyO98rmlJNoWQmkdrfbn/x1l4SlR6spLYKYlFUTAh42
9l9SS/Pex0o1Gxb+SstaUfuIEl2esMeqe/N0x1wUnRsGT41E2PCwWxDfYA2ivoRn
9ycHV7gWmP5z0ZBBmzYSMs1ujLIcRBsa2yD4btSWmb+ezXazp8r4BpaHIEEIWYbw
npjex6im80tCFsjPu9cd3W6Rl1/vo6F0JUyvX1BVkb32TbzPhO6S9ev77nxnCCXe
fDE8cDXxf4AOMt3Cd2mc1tqiFaJX38cHkRPS79ESeogr6FFvNnXp6ZABeIeIE5QO
j1ZSjdjFUBN5sxm8lI8oulZE0uxeejNKQy+hcpCI9yfhhNWE954dMopWOSOpA8FE
a4O4QE28la7Rlf9qBfHsMzaZSWOEgZtM8XecEYmq3Zf88dFzyulf6a9qtHStfuLV
fadv2HbRHmL6siEWB+rhD3VZ8qrAb8DnGjCYjsl51UcqZM5ASlRLYNV59HK2XfCK
o8/FwZseLRSzHxcwwEHU3LiaJA+lN0DJee/oWyIcHgQEYugfOqfOyO8RWRP/7g67
oZKwAOrQE5ZZGscw0duNog6IHvrbZ2ciMGoM364RS3HKd7o8vePj5ZieDN6Yu7UU
RNnjViqJs/5UzkemM6QuCRkbULtkYLbi574qn5JnUz9BZNUQqyfAXk3aOzUJ6CHU
ujdwDlCGfyhT0p9GPJhoEVqVBabkQRKSFNGLN4kJALjinLGolAZhmi7nZKeGMpu2
FasFmXERcO9/K6e3hSLglTRmaij3/7YBB/h/6aPQKZ4j8DxStgXgln4e7TNj8V1E
gW+SDIpJjBYuVW88PICUEhqNecVveBl+9s82Je9/y00fzPqDGnNla4C3+i8iJv5/
lIUALlZ3qg9kS9Xc/MkpKY5rmBie8ouMHa7geeUHYkWSUyw5IFHmrCQaL+Bp6kmX
/R4TOmwJXfhDUYBa2v3tWpP69sQ5W5cFhjy3Uh0wmHfjqcsxlNgncPPG+NpXTLE0
i6b1ixLx090fzMK9OrGOr4KOJQhEBgUUgJmqA+vNtALZ1n1AkeUfftRgtK0E3dr3
kjkv8n2IxzU9LttPINaZWdI6NzBvSGO3aC3dfhds3+9Je1RqLBcFMo2p6dkcLiHC
31QkU65tjw4BmovqRE0A/ejrWjuZV5FNbqL6og+6LpjwXh6uyaD2TiGkc6Sy2gEU
OGKCCT6EmGdrNVsdt5WjybjwyIhQ5Y+t6dcx5OROiq74szDWz70u5Qsd9rjpwFMg
WjFcwy9zrSvMQlHODGNTOq7ifYfTV/OZHuKuvqE8v/5XquoH1S3K1gAD7Yh9nrev
ssMxQmLjz4k7C+2WEjLmO6tTeyCk+xxo7Hh9ssULIanZMd5krIfY82DGhCQ2wbjv
Pcf0KKSvpTR7jJhY+Zey796IkC0T6VCxnd1PI+QUOXocQDxElWGwgH+uZeYQTBCB
5AwJUMyIYuKRt9P+kE8xfKM0UzYfhgU7JJwtDjei0KyXm7GA+G3hvCPkQEssEnWH
n4tERupVN7UI7Ez2bF0+Lv0LC21mFkoQFzC4Y5FoILgY9my0IIF4qEI0wfqTxki0
aVUZvu9db+3x0x1bAKhkouRNK7nu7T2A8jFsK4WG6GrRLDkPuKSnzb5D4efiYokr
e+NAVZoP/CDF536YClR1WuSIWzEsg0GSuAaWvOYF+KwwBqevfaD4MqsSd5GHgbt+
q17wQbKl4GJDHoQy8L7jDiAb4cKF6Ta+HVrvOTmRk76fmqJYtenRTiDGxZ2ejq6d
A4XqG8xXxIdk4zFOmK1uQ3MVKp1kBl4d0kIq0bktUjIs5fCdjp9z/mdDr6NcdqV4
fY8cZpU5Ru8w34dm9i1etYsHrOGYMCQvxfrcd/zAS4fGavH/xHZT5CzLE2yVHF57
ubose7Z6KD2ACtrPzr0FdEbAD3lSDckiEV6Gfu01YiWVflh3nud7c0Pf/0oSE9Q9
ktUDu+9BVPeh0AdJM88L0wFKPtl/kUOUpvQEumhTGh1AgOu9t3wvWbgrDDinVVmq
jW3eqwxf7Ilt95683iWoM+6//BTP6wOmqOHjS3UYVja57p9ODQj2LLNKt5b8jg5z
ogjbdU+uBRYlpJHrNA2Bd4KPgt6omcMYKIBiQuwcfyYUiuD2oW+wfrGRyIqbHmWH
DQXZmQ37fIN3R5hqGsGTpkq1puo4xhEklzv+lZyuNgUnbN7KOQCikC4L7zQZCB37
Z0VpFy6lYMf2jat7X93x7rOnK6KCOBFpcCB9NPQDHOp4/zTf1GVjEup5pYza+tSQ
ERBks3wSdbbOwhQr4GxrimBMjq0Tjru6Hez1zRgKlQTmcswOj99brBWBF1iiXD1p
Ozr/CyENPD4Jk7eOWfEpZNd7gRJQ9jscsbSQdtFgnTZuhufWugLim833HiBT9Lfc
IY+wqZlu+dgkibxp1CARqCSYhHW9sJkZ4/9WoTlD5xYXsOEtjzLESSKdtAmBA+S4
9/+mZFmKQ/dfenEyT0bghFQb0mDfUyYP+VUuNFpeJiA6HqpMFbtdi+Ez1W51AbTy
u0fr/QM2zRySRYUvq/7FyxmqPOdwLEWNGMY18nw2c4oKIUUCC1eK3C5d98k2n+lp
E/77HsCr7mEQRm4s4GPTQrEXhjf7EyGcjpJF3Km5o8HZHF3beNAA7iK8jQL/BW9a
CHbWAUBSAuY8DY47jXkmBbNhrKFXAI1hdGIVT6wu6daikifwVecLf4indBhn5Ybs
sUr7aMK5kiDUchyHBXJcg56HaBUuEhscmGCsOA51kS7ls6GmxA16lQ6YnL1Im3u8
DqTZuEObID3gvY4ippZwkmx0waJccEDRbRZjht+eI51pXnwSloltUXOnti6bMST1
H0UzaUWqMSO1PrZZn1qnlSy0rqBaexSzTf5+nXpD1CkME3LVJ327Oyvr9oMmm4RN
yOvl8otfEefyYylt+99fRgTXYIkJyw8Fz4RcNrI8rgfgYkfMeuUvbL0e8pRFveGb
REg8AbI62j+yyX75id3zAUgCXFC1tAnHDKXtPV4Dkg13j1IGMWxOEVzol+5BkWQ2
B/TpQXqAHvmKS8r78OxglhK9zWDNDjs/w/c/46V4gISJo/3vXCv0rh+WirPwbkS3
POLIda4zp0hf+VU3uVMj/Fvrs1+jRUBKbq79/OQIew7gI7YqhSXeOgbN5W45A2GN
UgHjJ3lYbIBpunmrwgykelrnyvMz6NSh0rzcb8PJN0zYYkx/lo/1JMoQzsUDz/Yr
15BZY6FEzDSbOOMO5KV2vXOy1udtNjHO48+ob91eIM3YVub5VGiIxHQO8u6OfLiT
ONvPuvCvcNeQfsn9d0JD+sk/8Q/PedRvOVOTwjIv41tbfWbyYiwKOL+n7QXoooMw
LTztDJzMgDvGKcUfdI/C/j5E+E5YMX1eh33csGDsGxwGawu7q5R/K34XTQiKdUz4
eg9faiQ20w+f9thFcn6J3kSZAFSIFOLmgRkVu4CBhPfujIjR+EAHgApLLzoX0uYw
suwNwIfepDy77CuLRSIurEixDrDJ4ZYCiklJtn5IVb8r42GowF34ETHmgT5MNhof
I1mHzj7vcP+hxeWo8slfKIxSo7tUgFeos8UxK9l9UGrZpq0/xvTdIsmTWi6zP32K
yeXbAyyr9EiQay65dsWtlBBgcLV2soq7WaC+vRHskop/paht0Z/DhL7UlQo0eH1y
evpVvB5Jt6Udo3qTHw984YUj98DxSKwP13FGBIwUu9+B2QdVGo9U9SnCQfVtd8cM
paMNnJLhRW/p31IQFvsM3HciI+QTj/3raHsCqxKp3TBaU7NXXY+LNRCdjme50aol
/u52cpfcWmxUPqejl2jMT2BGcjwQvJq/K0/0vS92/7qm465FaarW3lqjABS2PaV+
Y2GE5ja1gRmsD2i/Kzhqsfs60PXJYmrIyCJL6BnF8jBflOLzDklWoCYEcIVFsRGG
U+LUNdTyat6iRBIVsRibrTl3cmv2pCJxLd3guMt28ZYCsnP+Wzmh/G1UWRk/UPPO
q41z8pQtdDpA+ZoZE5yhqiZ+YPdUbBWf1gCGzFeYiqD1eIwE3V95zuEJovAB5Wuf
N2YhiRe4QGPQZeROuicaZTsHOstCSYITGF+CkQEqyZZ8m2v93jNG/AQYz3U24Hc2
HH13KdqaB1jclRTQEaw6WRHp0nSOceQ60rGHXHOMWIRciWjba9aIfBxbn6byeYZp
oVWzsrxrSKyygtv9zdOuxRkKqzIjIa+Cqr+n5aeV20AlJjtUFGDb7d1S7bNfh9ZT
pb0wvCJ9y09P9idERLDR5nMmfjdINGXXI3VA4FSCWxfF37Gjr0Ii/VmUwf3H+Cb4
MI3b8fjE9/XLJYEB2G31XgJD0tXNoZue0cR2mXYyQYzGTbLDr0vRCGZv3wEXySrZ
TWyRuyCqhoyzR71okZ6M1F0wiBItD5xfYi42J5vyrvmmIhxfIz+pCZSx81QF9cnZ
7/4Yjcz+41Kh2jgudONi4wT4K5/7+2NTvBnGJJvgYJfu/+wgmFfHeCinl4NLyVeh
ERqO4GhYa+wFCzqMiUsblDhTIM+sGpcW9NEdSn62FhGtTO9ZlybhKlXP8Zn9hV2H
eCJ8MB3VIQUbEfjar4l8NstDqb0H4ADgH0c2OGmPR0cpIYmQiSc3ssu9bULM0uXV
o1qF5yNDyPJKHxpSRI5OurdR4TmNdgPUBI6fKZ78Ug57sZGSAvNWY3Hrgs4kbvDv
YhR6UqfyPVBjqB182TKv/smIaK1uwwX1vq3Q+9jiEu4HPmrnfaSmCWhOQLKNF1TI
XphSaE7Dsp8gCUEIZymt8fmgr99bARnf3WoVpgQMMm/K9+TSAn8Ey/8xW6E9GCxr
jCxGH7YANXnk+r3YwMu/D2JJL6OGsHWkVgjW4ZgaPR5ayqRLdKUW4j4Scoxi0KF8
j+6YNfGQpET7BRwjTWBbsFnYk5t41RSRuOJDg1u4UUznUFCdocN6brWWkYi0AcMM
vrkMBVy2JVBz2YD3q37SCYoqfE5E9DmGaDtUmaVaA3XecFRI68kDcea1wZIOddYc
6uuKBQTlU+Np+etwilv7SHlZxDHU3fyOTlmc75Otrr11TuuGr0EtVFZC+CclaHuX
oTfzZajLK/znF2S67CwRHIbPxgG7MwAhbJwS5dKlnLzuhmeOVBjEOftuetU2XUvI
UggP6PYhfj3NzStpiFj82EKBKa8EIMsmrcDuQjFexQhN9GbX2Sa/pVgh/rHr5zLD
BH5ux5pW8s/ASEJT5ShTibjXCY1LDjHmGLe2b/rqLRgjT4+C9yBt08SVhO7W/j6y
dyDA3b94qWOa3QvdcCBSGzcEu4Ad3g2+bq6G+4RbfJM0ITOmsGOvMQn3YaWq7zFM
9+tutTKjl9EOCOOxpE4SGKZQG4GuXXu2VuB1re69cR+5v2WiqeBKhYGIORDhTSfm
LJ8uEMQVSwMbXc5PybJCf0H4cWo4q3q8jFMe57ovz18pmLzPiLgArOdAj2Y9b4xK
JCn/RyN1Wl3BWNQejM8O8NdElddgf76AG4YmnB5bs4SfvRiHF5D0BQJo7+WjvPmy
G1gvaaFs/E63IDZmyu3mCY7NfSPic3QVruQv2Iph0b9vdMSwJUdT+fgrpAWw1d3J
xtl8ibz77I6I+EUPl0o2T9I9+Yna9+KnfPCXDkqf2lUbUrhp2qps371BIUoFIglL
fyEbjmpp2OQG69KTtc/RSxnIVwJw9psYxrKO3ZWCiOEWcoGMNIa5NZqpZbX+Yug+
GPO5YCafxnQrzFfUOVEaTWW8+XSppJgY4IdhcgrYp+s762PJD8YtZT9YAukZAUKC
aKzG8yu/2akCSa7de2wwVu+DJjzAXH+uDKJ65WEkXYNfbilcnb4s30mOAkxShRqN
cpP1KjNymLIOw6azsBNeB7O7wG8lPGIGruphsWc+I39DhcCM3+xt3wXrak5VOH8S
OZsf2L7Mkk03MnueK9VMF6aU81QPJgIauSt9kC+53lNosNSnRhHVp4nSjEw7aZQL
hJ4CmXJm9DGRaI3kMIyiSSGWe0ql3qkLsDeBevEIgCtnubgNUWJMX58HShNoQajB
jJApLvhmmj2eDvBsGFIqg/5Wv9CFGSxsQtKNCA7jcu7JyQGwhymm56ptiPp4WerE
LxMer4yR5c0KpEcdjRZZr/YGbTPo+COI9qbBD1JdKzwRRQNK8s/nHVOxfM4sjuJB
Xevgp0bhTSg+SGG6q8G+aWEST6Ewphkq+7951yytWJCfD0wUFeR9be+Ag2QwjTvJ
eAxJGuNbny/tkxCQsi4PWaDXQlDiYxGPPdW4+cs9tHQECNEzOqqu0/6wpXIjgbWU
iYkvSKMt76JFF393yL/Rh8mohklC/rY0h6ow4NDKenauzt73j9yz8yYLTT92cq/G
c9NCBuz1KTrjN695wUW1UvRmxJYV6ZYzEWLD+n0nD/+EvS0C3+dtV+yC4MYlE7rS
9m6JHYIoD6ywNvyZMLJ0QyamlXWwWhjm1fec/ClTJVWeq0eG3caAFFfGnFImK5vn
JzxatlAbDrAENd+EtbDLS16CYcmQ6XEwS6712rrGGwWRsBsl3Wb5LkJEjbtY3n+3
uqeal5wfJD+sSTylhNn8u0nUQxp/SVHHaUYP1p4iNPG50QQrzd7NlXH0Wlobiqf6
Wr+W9fD8lTRSHW7AFVEKDeHIxQ3ohBVLBQ94Out4CW/omZVX34xykPKxk2POp38W
0oZ01LxDy5FpQhUmMXt59ZSNZpVYR/JijgANLEKKWwmvNIMdfcMNxhUL/HLMkmOE
7zbtgcSsn4z7tF/GdmFiZo3uo5OsGNDI/MMCC7QV7jU49R+jgL/dZWuVr5fbqqwu
7sQYewhajh1eTcjC+mmntWXzcGR/paYhXFkmtbA+ucXdNdnCfQ79TCgT90XrPVJ1
fPZZ0VWSrp1dDVUSjiGJ8BA2b9WQMulCVo6jxLPaffHDrX9Vz2c3Q7Nd7kcB1Yj+
x943tUhZ4yzYM1PlbhhYF3DBCP/9pRp5Nd2/Ss42EIFDcWzeP0gmto0GLdC2ZqX9
A4dzpCUSuwsPe7mOl2BDUhxrw9ax1GMbmloDPQyG14BDj7m/Telw7Zjo7srs+DWQ
rEbVg7tnfqI8t20L3iKYi3GAvElTZo6iClci2Ryt3o8qjT5zm/AbIR/mLn9cGnzW
saOc2ILh+17wGNM2Vj/qk8w5PVNxQxYQRehbzj0BuAdpkDgvb4fwdhGIu5wlXzRH
2Kejc0ENGbt0vW9wgTxkoZYJ1pOWROn9Bpoc/SgSF3TfFk3XwBkgAfQZ6e732oN5
jkFM9Igyfq3L/nc+99+wObaKggyOPqHIm+/C9p8BFPCtO9HR/2qzuDgWI8Z5JIba
Zzzacg3w4Wp5rK7hzjH0LZtgVk9Td9vKW3VFUSRW3YYEHaTqOgdm+nuWISPga9ov
o7PZjnrLW1Bec1Kw+6CHgUzuaDhsxbMShxD9jLdymBGsh5ZpEPc1x7d+zzY85Emj
U08IzrLzZXNT5fqFpDFoP/Qj/PdcotU8sJ9zx3Utjzayxaddeb5LJ+xfLb2YCY5a
/U3RqA+J46uHDBKtQKMj1miK+IIQSbSoHkyJnNebwSZUMztr4fH2GE5LHZggRfFw
A5kpA0giW1UV+HG7gZrOfkpE0KADWU/d9oE6HdipOfso+ZuGIP2oD1BOHBypOWFB
DlMCHO5iulOMad35daHOVNjER1hnWBOjK8NPWGy3nGTCY4aPg+zheza4C0e+ZgeC
pNKFFAlTjMTNj/zg8rm6EhqvcKSDcPMIsj1thdiNiS/D17aAJ2+q+OZjY2dPTXdz
72xCVCvotf6vfKIatwzSTHTA+1QtBYRb658mm+hgrron7eebUT7vYHjgEx9JRIRX
DjkpJzAcJlEGc9/nSnaFEfwTX0qw5sy2y7diO3p7ShtZfwW4iydZwHQuEQQHwNRu
TDlyOCo2+Med3/zOMk33NGde7uOxBwDQrxEnT+KXNEywX4NNMkjAaMcb3z+SMbsy
joaXoKVadl67mW3r8mbxrMyU7Gm8QoeFK7P4rHbC5aLixul4kr+t6aMDWUC1RO/V
u7HlTI/sSUhyshMBTzsPf18ZsfOnhXXMHkHXJSJ5vqnbDE5FIj64J+QdMf4bw249
jG59CFuvKJ2zFppx0SR21m0lA3TRfP2Unwc+FJKSpRTSsZXYJMFu4Z6aXffEJw27
HsJlkzt4qfSh0I2AIuv4IMdBrzl+ndbYrTunGO9F77Vf9MIUeRyHHxrFOnnMKxfK
BYq+69iePYPc6nMsQlUX5byDOqviXL+X7LaWzcRwdDjJyjePqBE7tc92rV/yTEiX
FzDHlvcUZBMNuQrFMy/POn00AdNmtgWMMHXZ4IXiEoM8r7MRi5ONHe3u9kZ/YJWE
Dlrs55CSJ3WZAeh/UaXi0d2Kmb+WUKiOhMwUPoGTsnjGRwR0y26RlaodgiyOo2uj
LbhUXfAUtF+Yyd+u26/IEmPj/6Xdw8ybMKH9hOP0RX4iW7DJ34UfphJ6bJ6C29UZ
UPpsOKDAW/ysRr2uauecfyr+7Mz/tom9Ew9Kl9HMZRs1XBieD+QqPy6E7GRPKGw2
k2R76gsiA8Ik3TJfX6p+vovXTpHbsfOanJvVLnmHMYbNsE0Pt3dNzXfnEn3HjXww
hzBPBvQ2oDN/yYej2o81gdVJrp8Gmj89knuvYkkB8h/zz0R3Ao1Mkhc99eqXAltI
bdWC9PWzSNFZV79exUxxziZSDktSIQrwofY+fhQTReuFNVaR9qaHL4xYB1s4bc2R
vBu1ifGjoiJ2/K01jEyM76MLklT207BxwWM85kN60V1cAciw0Nodnz+bj/nR9FCc
RAHAqqrKROcFLHak4yd0p7p+7J9L1Rbo5iMMC2+SKsULn2BWKKMvdM8UnPbYHQ/K
8m5UcFDGd9Zp4/WXlW9v6Vcor9ULqagmpflTydUQxydbHYUUvyOIKfp7KsKZpCky
rRbkjSdpX00FVThptLUjUPE9uRhX5oJYjuE774nuZZKg/uszCkriv24XPrZ7GpMl
9wHl7XHBt2VJSDGgfDOOPKD6R1aaxGYIjPPUtSDT/RJCz8872srQ05S8qDMnVzGD
mpPexBWFzBGF+L4OBSabvE0ZOZxP0mqvmJoyqAcDTtteYSzoj7bnyJ0UJiqZ08Ub
4Urnq7TZtqpN2xHz/Ts/Yu4LvA39tocTyN2kkw6VNcfyEcU90mST2PIUtumDwtas
F4/J3coNrV+wRC2t0/5tfQjiVueEo7Hm/llf7R5us2Nq64EhLiGWmrmROFiFpWla
A0XutgARuxtnxBSipV/nRBPE6ACqDmcnh3ct/XWZQ5pHsYEkobYYthgzQYc8qtvR
nzUVDeds08bT6v37HTCl3NFr0MBDsIk5wLsZSMJF096Vk8ZA/HQkuhb+9vZgHUGU
vSiveDOfSazIhg/7P4URBOsESMiZXJ28yr0PDy18ZvLTR559VlzpkiomGvKm9w9e
c8B/oVf9Dk42rqFANJHnJL7kPBkfxqaD8GuVYj8m8WfgQXiVWxW+lhbPo8cnTzUU
kWOEW3AG4fdbeO0zsaS04BcqLVdsDBKGkCgoy00vNKKTqOmczyTYyVyBSvCqo1lC
fQE2d/7NQ/5s14j5rSB/0nlSNGMX9AAMdQRYwuMKVfYj4UAH82zJcy9PAosYRyJD
JCwHeh/LGjpWFwSx4SsKiJWPXi80EbxqKbWDCob7dxrv13cxa1CMoBP90ZZIokUA
EKz84TGa1TuCKRGihVRNeduJTUwWtOlObJY+tvQ0uGnOQTPiWHTUawV6uohAt9S7
dFjK5rGr1PjmM35UCUgiC008+vUnkP0gKqmOdQofFrPsGhUHoxK825AvMxAWRzlj
KSGSjLjZT0IRw7GQyZtF1nOUsUNyktFkjeb8UnMTIkQnJUyk1Nx3FLj980xb0Lp6
MRJ+l9Jl88yFA7tMwSeJ1z7Po8ACNKsYhBQYaizcEdM96oF880//X5d7b91H3vYp
14ZaTNQyACA4dnLjBtkv5gMw8EpGcyuqWYYZ/E2u8wSHxNlzXBhFgeNTJ2DuvWct
n8fV6fo9pZeiQzIgen2gi8YxJ7NSIhQ8lA3T0EKomsadwVLz6vFAXU/Q4JbEIquI
3LdfEVbAcGejik8tuiDnw1ai+HLWFicjK16081GEX2ma8Lihre2OCtgH8qZzC15M
zDWAOJFoMS3YCKA4BBh9fhEaeCExMYehlc+nhmRdk/JcueQeao5f/7pfpuNkBhGG
HF+5HBKw+dNLtQLivbeIP8sG3lL9xpFcD+tUthmqBkEAqrA/GvgoeJvsOep5BaBS
H3R16zPBN6PdHs3szxUoTA2tZH7OQUHl7IqOQLN7Mp+Qv8K7meXe32FRl/2cAtna
iqnMCmzGw+xC+WyMCRuKQQ2kIn44+hSxQivTxL/9VFXogeql0tso/K24BGKktXHe
t2WRxP5IwvhHflSDGruaAEr0GSnCcU9WtrX2++oHFaBr2Q9V+u4YswfBwItCK7dg
7uPw7qyE6cJ32suIGmYLmfE1Osk6pnFtUUB9M7TCfef8cEvJ/xYPd/Za0McEe+59
690EU4+iu/vtHFbmvFbCrATNZcPZBd3QXXEW1ZHBQE1M5cotYHgzHUFX+sngF4d1
t4IBkHF2jpxJKAS6tAyRWAauH52M3u1av3AXbDQ/YwxzJkqTK4wtLmabiMgoMa8k
fqwVb97pan2oJhjHd9bTJWSfh597YJUydEgdhQtN+mCPhfjfgw3uHGUoY6qffm7R
q2v4L/FhRZLuKwGu03h48qb1+QPswjAetVgOctoCG5wvZ5EudKm240VmMZDN2QS0
ljicfPEQXMDqM41gNmQXsOnJ0YRU+9rIGmO6xrR2S+hKyVNxonXo7aJ+/YIBwdxo
9I+yMLfKw0A4Q5UryYuPOMI8O0x8q93pGF8pue/GKbbKkk05lLjx2P0ZMjuko+bz
sXNJzwhzwaWwSEFUcrARrNVLUSb+nd7p31Ndq32aoYZ0AWkVquSYwiN1MorjIqDR
LXlkmlWy+kHQhbg9IlfCkQ5tnY+2LJceZqmJYHxex1SI+0g7Vj5PwcWsdrJ5n/9d
fn5hzAwWawS5VOo2TI93IHHMPRQc9+E6zPtFZFyAGtiYT9qjNMd5kTm/bGNAjyvP
xN9ydO77EDypn20IQSY28R0LE/DYbzd6LJzLHpAnpL5QSn4ynTUOUhUZpZBuvbLg
SA/ce4yLye1s3nPLhHE1xoxmIpYln0Zb/SPQv7/3dsdg9GIrKdyT8jXK+q3OQhq0
Y1gUF1DiRJylvNuoizM3cfGIpsI94ow6QgMtW7u9UT41x9UM87HjMvl9NbSx4u4Y
7orpPTl6NlN1eFCLxsZCYaNdbVJk9+vtNGY7S1mS3nlSgDfQLyUoX9M2UNmR0plH
2tNbkiazUdkDJMp9pYGPiweSDJuil23EU5Lz8na7PfXQqyyy4Jn+cUZQFjc9gUWN
/gm/AoZNssNUwspIQ+ChkY8WiIoOUefY1vUn1eEyyeHxQLhGYjtnPJ/eSASk6UpB
sRkVRxYHf1trtAnyzTU2zKIOFx/gDdV/skJIBnLzuV7CpLvNWY4rF7SZLh2pFLBA
22Isnn2UNzfEQVxMMnoOCtko+bi9Qd+J1vQU44yzEjz7KlieGTO+9T5oPkyLGANJ
tb346NHYbSc1mYM9nhNPXAsgK+KaZ5ybYabF/aZ7hgMfP8T+FRvlXZ5X0RaTUnwL
nIZ8ruhgTPCYlK93fsuuPKV6cPXVP3ubRbaB4aKMjA/k2yFsIc2cY0xx8XqbR8x0
rydauZVfbkL1Rh57bdlIvmly3cyZq5d0fvs6SF8hPbHuffYxIkaJHPXiaZNK/92y
RnfvAp137/FquzsUycF67OnDDr6/L95EjCkbTgYG6959BFtN0sak0fj5/jGeDB2c
04DfDTNiAo/qm2enp8HUkBjPWZCJSBPZIlSB2fQxhTTx+jk7XewMcvtZ2rKyShoJ
cosgIUrNPYY3hAPYg2pLWvjAQ+ZpOuOR4p/8oVmkW3fH1/LpotMDw8p8JlY8Ynx1
QAz3N3e8hVfgynR0/Zixm6q1btuKTqd8ARsqRqwGudjZhpbkW8bU0rT05Y7QEWWU
Ov6IHXnlVksMSdiJ92ryGxFPLUpvkAj6NvtwmqczZKszGOvEUHdcKiZHlN1BW32u
KQlASIo3mPaj6LkUAVFa5kIPjpehVMC09e/a2hD7LI0A6ES3xxMULJ4RRnIIGpD8
0RIUVlUPMQBvddJLAJbfNavszRn8CB71guTNQE7ijs0H2iDNgO5WCzreTEV+uf9O
+BPfGgOHjnRW33sOrw3dQu/mtK34poRoobo2l3exVdwVsnccR1H88WHbyy7xqqfK
4MTtADu+Oyu73/42YBfYtgVEfBOhFWPo8vzqbvisLOsZizF2jTXV/c8kMpNsXN90
IuUAn0pnjsYjRXoKFa0kfJIQqSCPcMY7TEZ4OZGJrMjc4HOy6ZFDcMOUjG+E9K1l
r+x4DB+1Bhqi/umHaY70CX8RGvhXsfgQzLGdAt0tzjvtmEqv6HSy18YoFIByYM99
GPT3W2ZGR3m8tAkhsHQSS8IyvkxRaMEV+xoj2zeYFIbzAO4B6io6oPUdRscboG0C
IJGTpv8jIRIZ2m+ZJAZrBPPYmjs7IiRRbuS2fZEc1BhcRjBqbIJ6ofQnHWhmqqZS
2G/L9c2UHdCiDs0l7ruVn7S87Pph630EItfK8j3DdLKmo1WDrNv5XFd6oPV62bxZ
qPPlrQPBox2VEtygvkEotBOI8OFpJqSJRCyc2mAeQbx7siRlluwMFRLik9gz34rr
pMUvduL2prNMc6h7j1G6qj9k5+YnJAHSkQP6TC3rr8KRIELEaRtREcKPA9+S5zrt
C3eI7qFaDWAk3vH1FpOnZ+RJ7YVHngqHmOwaw0U9FOIIRSOc15xpFbqIUkUPBQ1k
XaAcKUf2VTkb0LUdowbcP7ca3ZAHhC9pEUrCQi0rOqOXrlhsLIu7bMx1XYM8qTPB
u1R72Vw03tpC6UUTvvCqRRUO/MNXgXh3n/BFPlx/bKC/jtHIhYD6Y1y3L2ny5sij
4wgQ3Jx4cZJo5iAiZfPJkhrJ2QPUW06lUET2+ztmAJxtQF+nWY2bSJP1fPN+GA14
vt0hUvZ8Pt1A/KULF2PbljJytxlW5HCNodxwJmeMKdtBNtz1UX98pV86hCCGO5JY
512uS6mhpaKT0c+74ZKe+qp6L186h2e/8rFP3X66E0tMbSV0c2pc3T9FFzDP/xtn
gQ+9p0T8HU8PztXadMYz4EpGp7IpPT85VF0VlB5sCTcpmUXDh7481unLLeF/fqOm
08SG5IEMU4+OFOWSfbVVEhwZWIyGLaRQaDn1FWed6AXk0fI1q0hTAijSKrmigZXz
RFzWCv6roiqa6pdvbg59U9KcKyeYD2UPQS9VBW7dpzWiOviZjiSGuxzfb2eBtogs
o0I5DkR7NJxJgAadHMJFwEhJafvRKD1KMP/dN9Vl/enZ7gjcf4EZ/Sr9CKN4UxIX
Nze84rjFWdyGnvyCSHK8anEkogVOUftKVk14HTpA9Q/YqKPkQKQzLWEQPCsmepYf
f3DySjWV9aiTot/EXY6K3iWeADgLFlh5jd04obzEVvE2B9I240OF2xlnCPd2lq5f
RkD9f5q6bw/39dLIheFb2hOg2p1rWeqRmbKJhPRIefOu+mCMoPrjJU+n6usDTC7K
t3F52R4vUew8y5H1T8aqQwhJnCxZJ2qpbA7mJ4/gPOeWMsbtALvToVqKNI+7TE7h
KSk8AUzY+GXfgNxU4mGnyp+5Wm9hY6VHFSvrjpB/VNuLiuAKLbMYtpnO4G5De1up
YKVoXTAC7/YjgYiO7GMKd/Yu9I1sWFnS1ILaegly2+u6X+jJKdJDjAGzibqXraYH
Qmp0Sx0jrMuZjdslzNb2uEuSpoPc4SvSLk6TyvljKnfc0hcbYNOSeuTBcsf1ei40
BU6Z9UIiccPIQsCiO5emMvugRDnKfgwjyvhfxAyQUx0LIQxBt7Vm1C6Qgyv1hoSq
S55I1J+si5jXBB35NZAUyifl7TO/BK8HKTS8Ygft1lmhf8JaE9YuKa3DetJNuuIB
FdI3MHcNbjdl+o8ZC3JlMS9hwWenMStB09qqTol58T3Gq6pQJDDmnWn0SdVE9NFk
wN2vOYIjW9gvuTO/6oCE45F8WEUvhqny8I+fQE/GgpQvAfPAQWa79zbfuFUEL8rE
i3NAcQrgTzCubgV1Fd96hlpS7JrE0hIAwnWjlN/mr37epAWs8LBC/WMzWEgCMQ+s
VoZs/DlFL0EQWRJA+z0npMYpS58ib/N4T5Ydc/G+zAp1Yunet/fB8UtjxsfOk1Su
EYz29g7lbqCZgfJBw6RC18MVyQtfO5eLNEq1fG46tKpKGpoFul0dyXQtoCwqy6hq
ifQvP9Jdkq+Agc38pkZGeUC+dFiY5f0JzVhII8UA17Ks2K2IaOJppELiJw3IYCO7
BFu5tIW1kUtm9799diIa5tIFaqnYD9OOrEaKGU1dUzNSmkVZxvcmpku/OxEYxP3M
TPa6h+4gBDFppxgkVDNqZQKcGYotRDK7IsmTlYpCjBp2kdxcPROlMNVM9kkwlnNA
BxNa/Nw/bPC5bTsCcagYBcIZoXWVkJWdJ7qe6aF/vKMv2jNqqXCqw4Ps/qJoimHj
fa02mv2MxNT7gNMzUK7QKQn2juw56A37KhyQbqjBLit1zqz2LnT//C3/qF0FrKWl
ikAY0kKiFMz4ACSaA/mbyBU3zW+myw/Q2KqjQ5LCFk+On4qcEeawvSiJzjKWSM6n
qmncf0cxgiyv8q11WVXonoVAUTXrCsFYOgqK3BDhHvtlH+AG/DHC54ltsneDMn7D
ytaYdWKsRYstKtz+kueA1krpWOBzwJ3uDgky+h4zZLyt/0Y2mAsMooUSd9j4Q3mn
9x64+83/bGIsu64c5AH/67756Yzke6yqQVRokmyrKsmPd0za10KOWQ5eUTXS+kJa
WDVX8sbWYBQitogqTQIURVOLnjiaVM1sdLvSGLF6ZR93TGfxdJT+56WR6GAx8Muk
SsK0ym52VbW4EEtz+5C+j1ZEUXKoDaakCuDDanBjTSTcIt7ckVYJbAKOqr73XeyS
pElx+sUzXTF0Qj2/nB0FN1Kj5fb1N5Kp3WAR52Q9jLicCW+7tMOabRocyeimLfyT
rLvl+TYJIZGiqv329xoCUSPuEy+arVLAtUMA61wU83wyGNVkKFh50CefNh33Q05j
7swPlCAXHG+lEN2iGWyvhN5oX8pY5rDsb5FH5KGz/eRcTXAs1hIaBxp6n+LOM4Ie
CUqTztHnvD0ExbsFFdpEre9hcVXWOUtOxRBAPgcPBc8fVqiJkumwLGcmIHHQB8+p
kzyNUgJw1gLsf7ZKthsAXZTV/R6zQFlpiCSTBhUEDvEDBqTkl+rQ3k7OvvEEwDCj
55vzeb3onNvnH425JITNX60Jh19ZQdGtT6v7CMs9tw4Kzw+Vzgii1JbrZzSXMREf
KjBD2+YN0pXBWTwjByxvHv+6pvosO9eFFBoadTUPxtIoCxt0DEEuFnpVXEIwpxCb
92YIpA2fNKLLcFz1GkjVbMZQFujLtRCF2CIlSAqGoUYkPqDowqhgykKcaDb0RX/2
i56EJijOsPMID+KQqkDtXrscARIW1cMxkIPAwL8ZB81AmLGjI6r8cEqPCiNX5W+M
pwLmfsrQmZ7LeN01GOjtu3LOgvBROYgsIQNS3wobL3ZerP4HeVAknniEQjPVOlDA
S8BVs7uyE4GEk90pX4InpLzs08h/ddEU+zmP5w+O7/GmBpTo+n1hG4pxMGzFCyYZ
d5LA2rPV2vcbfH1by4h2aK9wkRifMr8vk0Xihwl1zPf/VdAFFJD8NutKtvVJvAmn
BDQmXxEn6Y4haS5RozXBs7ct5je5djAj+cPU3uyACOr4dqLzJP3VO5a1oWaCSaHf
x7CRBtS+4gcgC6Lo3W63mRLlPUJGYGbOw8THLLOoAlbqqQ1fmtgSkj38Dh29EXlp
/TOEQrKLz88giufq0Um6HOPg++5QaQXakWfYnLxIeimymytRfW0rPdR59K9qp+ow
+KdYfDuL8dxJjndHkH2OInZa1QT/SvCY4pYkI/NkZVp1Eu+WKdRwRU5OxRecTO6+
u4gu/r35bAC7tMGdEpVjnre+fMAnmYb6FSyxldf1cOkuCcZzGBVvUWQ6NU5qKsGx
SZ5vwIvklNIU0DoTtg9PKYxYM8LfBpW/9pN0HPUDKerI37RJ/aX5JeD12TFtlNCk
sW/+So9Kzr26Keg/yRTAbISwiN8rWYtTlnLJwYbMVxeMnRfcOFdww91f83a9ijUS
DKXJAMJ7IINZfB13GPyaqNBO3BK/ZYktOOzIS7fxvioCfaxtczldIP/Nt7BojS1I
pnMfyPOP94bxLwsXqqLeHh7gWHO679CQXWAkPT0YSbKaDRPE0mdLDlubeY9SnQ7m
ELR2qOIgn1XqewnHgD2Bel8nXJd+9JnoBJvXSYGA2Nhoa9bW+FMUdFpcSZWRKwiA
6/Vh12P831b66jKzdbnkDDiAEISMa0TM2qFohE4tEwy8GhPdLZrvju0nHi2w9Jhv
2cldikVuTC44rOA98ST8A0rNk8ZS0tRj4lVUZPXzPfDHy5kVE1rSESTnucguVgd0
KL40axLYRwl1SOWB+Ou+aKXLcmWX5F/R7UTov9+wmIkGqBH9hwTgl7ba+pOjL9YD
PrYJhmc/ly9qxd7qBgaSmahvKJkoRqWhtK8LuIlxpBQeZAA3t6xlYRsUYHlAkZCw
SQuXZnOtZCvXnnSIhyxcw929BBvaF6GxEZ0O317/VgeId+LLXa2heYAmI6oXQJlw
ii3Ifcx4cWjXl7N7DLbks+ISRKRKSVTtUU59PRbiYciEzn+o13SmoNIP+aRbJTmx
h2QH9k6sLQ7yRb5VjuaTXfQNjcWzzEjz9G8JN+F3zrp5SIOumR/p1slJh4/batJG
ZagqJ95s+HDmiG+mGAg1IgkFIDQq2L0psEoLfWqFBwXeVPKNL3DV2LcQCqxd493n
TU31u/nhVpUZ10Uv25/iu8hrNfrnaTYQMU2dVRTeBizBRnCDDAIqpNIIjgQ6agxu
zcEGixumK9cm8KE0Ee/TRcvhbwrSTDCl1HPrsVC3h6poNpebjGc9O3crIsjBsPx5
Vzp+H5GsrqnELKG3oijLYvsU8OcN/FEOKRDnVx8/hUY/B8xLuCZzwzvsV7Osyy+Z
MJH8qsmgcgDQQPJ65KykpXB5qtU7MbdFnHIduUtkFMJ1cZNsACf0qpE5P6xxO6GH
qVhT/wxDrm9nUAqKjTjsEcYwVas0RagLEv66xCfDkOdLPM36olMHN7XLdjJ8KL8t
I1+r9evn/5t+0Xa77TmcIPXyrIJYtihYzR2v9B5mDbK9gypOpikRKNp9pGG5i4mP
E++B6Yc/2zIDxJOkkQK+Dyj7tv6gcHtFLpbnJOBCDBf186ez/mKhXTtjtzn2Z7uy
SbYkPc8hSH5q7QydxOZDALODOLcssi2g08aHEsRO3j7bCiNOxfPJ5Q9+7qu0Mh5Y
XuFicJ8zcHjWB5rgBqS/uptlSypn8wiqW8ONUaLF9trOo/rlxxvyj4ArvqxCeadC
R1pC6zivDYd8kzGmAyooS5o3CgZdXUljuOdQSHNiffhlvs8hGqI6KwKG9WhyR0/B
uIoVAYVywra3AsjZsJckaNgc06FgbTjedC5HxvwBWkF2hZbve2OcOGGqcIg6fRe2
gFl/z+4whxip2vapnK6ebrzkMQANK63vrRucrFuizjWZHXpTtGY834EBvrTaPhDc
2Uww545Ub0iqZ6fSXMNFh2ZkmsWbQprMPB+POYpH0buoFQKDg1jFcrEAMloN+FSE
IdGlbj6fz6nND4o5/Z7MkChTehF9ixwl/WkvvfYP/3B4+7NAqrnmuKRgIp9G0D0X
Sklj6YjBN01WDiB8MUz0LaK58SBDqx6+oazXNFO8QxsleOx7lqfbGI/ZKYnMyzAV
wzXy9q1n1YRP0PClPVkObJGF9Y7hhay5ahkTJZYr6yYIMECFtpaRmgGA8JdamEco
QPIx6X6qw13ooFWRRrNXfcXn9FJC5Ppdf8sQAlFC/5tTEDKOGoKyeP4FitpNokrn
DLwRPVfVv284aws3oNNNayZREZkvwEC9eI5dCFywdRf9h1lM9hfTJ95D75UbU7+T
UnuaqLJMK7rcFHIO24/4vCGwTPFJKjmI7DvUHoEP13arCHz8/oTbhv0drFUvdE+p
BOwLIaDNwpmV+XGv9U8vOeHa7S8dHWsZnuHVUhMD84dpE1aMZAwQ2Ez5yEYzG3Y2
BfcggxoLkNeZWGo7JFmD0gb5gm2++xiGIZ9xRZNx39gXSM/nqsP9Y3/Mr7BozR9f
bSBipU0eEjMSdTg/woyBPaOIreZG9p0W8ezUiFeDsTVblDTWEegr8OHS//8WnrJm
Lu+/YslB81zJrTLmU744JyJtmAqva17BLZ0fvobknnbONFwfSA80lammEbM4k++9
Sgzgj7WxPkIoNEQ6EUDl+RJVr01/K4ZqjpCrV53eg9vm2sSlW7L+nk/qa7koxYIu
XH8knNH4GWFrNkf/V1qD1AS8wk9c43BL5Cndm7/DwmGtxd8QX2ma9ie6IyfnGuik
zRDQYSyPbtDTtr27xW031G0FB4faSGnNGft8k58W6eNh9wBH2CsjI6IeODcL/E6f
7pUQHUlIfmxqjUr4u/A84dfBWE971iZlbyzGG3E/hxJv2qnRuaTJISvuychxTs0U
k1o1pvuMqGgbGvncmjKnF+IjkZyp52BZy5f6OKR6B7on5XOGNzu6PR0oa2r93BaP
C7QE5cEw39Pos2r4lGmAnQsbdKHrMtt4U3fXY3WZUMBuoYp3AHzs+Dx0SfQDqZIS
7zrp/WTLtNm1qmWsbLaxB/dBgVTPmu2P5Obqa8QBpQBMgOpc/T6UofN6ywo1MKGb
DtlLeX3yF6BRC7bY7GSeo1iG/l1CMLRJfKcDH+xQEfGV+IPz0ixSotY6baUha8kV
3dYfA2m9xSh1Tq9DFYvQIrAhCW6P5EmFM7oEGeV6d7mCbJL3EvSHGPyb0AutIPav
cx1pXJb372sCWSC4QdnJwdbOsXi+LvbsJYEE0i9semB7uxYa+zPxNAHF5ulC0BRQ
28mEtDJPHyHn/uSyp+afJuq7mgkGgY1PeoL8y3JfvnEuleIJd2LQ1pukt8hMN4Q2
r3TxnRR9Vaqmh2PgxNb2L+1TAFYJEz9NuIK2igcGE+LrX9udmQPH/zxzo1l0JPcL
OYvP/FoWPPhEyAZtZqO5xSvgyBqkgU2WlsYXZvewQIIg9Q+/H+Jc5OFqgrHMXdCj
qqYKj8ZjCnQikzRzq7RJaL7EvUwxZ4a5bFFTw8+FWLZ/UWIIemLMH4wVEzVv1sg0
QIkru6RHmMDVhasUWq2SfIAvmWwr0Gcz5yUOqMU3MmH0CO3Bxi6qAPq2CT04zV/p
PmsLJF9MKO9RML7QCp0Tuj6Ab0RmHTJ1OkSP1XXO3xTIyGDFoq3BK9QVtz+Y19Nb
1YcDB/1dNgZFwDspQP+rQzjyLO7ewM2HgqzSYP/HWfXA+dzD3CrtbrkKFg1iwIWK
g3kfW/UA5hlB0+f3lJNZW0eEGIpvc8oLPym2BjhZIGQkDO7aOClqfjizO4NSqaKE
pHmryqC/VxGTlaDUM367fi2EIlxzdAedCcbhz/Cvt1JZ8cC3YuILIdOYq1mVdB88
tX7rCxk09qnfb5hWPPYs48dIhHVw4A1W7yUH2uWBEqGY2cp/j6RPRt5/jM0vmpWU
Zn17qWr5Q2o0aOSsIRsFzRGVWDUr9ExGt1M0VIVU2ftM2elz6lXD2hUuMZNtiDjU
HB3LY+O1DZFd9q5aULhA/qRBIHsb5DLkisJJJqByMWW1E3fgw33dWRb0QeX0iLrJ
ShgSbpj3UOHYxFKKM9cSd/LnfHzkGPYgWiK+K2cW4PK4brJlTCZMPtSL/1izg8gr
UvF8L1AdeQJITKjScUFJwM/kOAFopwxvunmnl3UXjOqDmTLH+YCU6ETCxi+2JmpV
8A/df36f+KkKXy8vFTvY45dNJiK+D0GujA5d8BIDCqnzYMrjP78SMChvUi0qZVjA
HZqnVohc5nlcRfJUXrz3E/7UI3wjR4bQ8n18gUr0Y2nCvIbJ/4sBjkzFtuHboFOn
plP6VXwV2Tn6oHO8gKMUd44YPMGDkMSCsOvovwavqX/YIRPUvZubdhf0gtGTyZMI
Mbx0uNhalTCkAZl0q9UtiOzGFn4lPCtDRMeHi6YjIEYjvj3XynqgYfWT1UjQCIOj
x/xYO1xOSsuTVgIFergPKIjbFSgdKNlwbxxCeqjlKBH++HGQFM3w8nOwsAltE/SP
OSIcHToad/mmlpUOkD/+5v/cxzRtVEP9VMi2V9EHYmEF03DqlwMbZm3oQkqU1M62
o+UNg59yJXxOUjC0GGVDi4KxYuWXE5RFWRiRXgRz+2Fo2If/uzXPHCFabSOndxBS
m9KfmDEv4TKSj75ZupVtrbBK2Z7pL43nQHXkGnBcZG5BpD6Yv8FY8tGNOmyrAcOm
deNnrZlajk6homHoPc5UIOwIGV7wU74nwbUjD/hp602rVBdtHNCF99WeGItsdslt
IX/EwCvpuCVkRJTqJ9F17qsWbqGeUOTlFBeTOOZP2FYA5pBOdUwVWPogzpaZ762o
thTr5yDv0x0oCrvSjdF10qjfeYeqfAMjvLlaBjlOVwmIVGouv3ina3pDz0riVU/Y
5hDi0ecPIYVybJFKJ2SMcbH7Hmj27yqBiFylZXYjTSP0yEgx3I0xrZmiJO+lFMU8
YWR/Fg+4RC9ItIpHMYcJgWFaz6AB8hdF6OOL9R+zZxxMCx5VuR5wDFUtWxr1KDHl
vl0ENGEdxCT/cHxDbqGqWBRSRtoN5TmPeFwW/UOLUU1ztfOlhqKp/QAHew+UzlsE
C4/fHkUcsze6EKBaKQR+C+sUjZ+4c/hNr25o5Zxbg0A0+Q++1hWSFpx6KhgdgPs8
21HhsI4zDEKJrRLDLM53vxE+wjOQLA0kCbXcWmB/vp+pt0zG7h8Bd5/+IO8X51ys
uSs4P0SQCZQTEbQf2mmgFgi+IOrwSeyDjBgbcE3kAsOct4MbBk1xiNKVQ7QuETQx
V4hyxMiHAo5kfS1l5L43b5pw2pSiWgCY01l5geHalU82mJo7bVW9CP5ZlRdq3W5u
vJqGPuWv3jCX9vz22TqTYhu8C9Mru6ypG0cpx4e+DiiYmCWFYkyZtoRTSK5F1K4q
8mG8EFSgULJLVmfQ7X9e0ByEZjX3ts11yrjV+KgaH3eNphlg8ozOcEUQwrHTyjr4
4yhteEF/MBhcvzjeHid6LYkHFs8fB37vfkbjy5lUaoA3tqrw2kYcFzSUqovpniCQ
CEZ15lCsuJFoBOTwHDCovT5kR2KAdY5cuKiGEEECFfkcu4+5azCHHHhYACX2OieF
yF5mugiPQWvBkNwJDwDSTE9tTWh+5UPWezE+P+0w/i4lutNz58ZJBYK7qsrCoYkz
Ao35ooAwHk0MBMLz+Aea4Gd9kA2xX26nF/lK24T7vNDbVFjqKY+tbV79iTHHcw4l
jheTwYYVzenRjm9p3W0sQS6SaIdPTyZqX6DzD7Ay5Jiwh8RlqjLFc5F3IwNub/8F
bfTAzbktyB9PBtjlJ2dLxkNjI0hn/I0vCqh9y2BsRcEzyA59xLt7hRoRg8a249CJ
DnUJFXLpEf+XI61eoQWzmWXkcLGrd6ZIeYatuc1qMPY+Ra4Ve594FjUo31xqHXYQ
V3mUt2LZFVPCg7tHwHNjh5O83i/H/7Itor+NArnQLJRAnaaEy70SmNJDvJZhOrIM
L1c7e2+Wrq6pZlcoT6w89pUFrJwjwG5qdCWCW2F27BF7HP3U17D1d2oMy0BrufRS
jeWraOv2dztzFf01ixDg9R91YkfwnLcIM5RGZ8FIfjttPMoX7uK19Jeys4jnNoo2
PrrM8FemqSfCFuCyCsRJ12rYBepAVENUwl68d5fWjWMTUF8rY6BkUi4vf/6MM6jh
E1ND/dmjc6MsDDquphf0MMDAevdqbrYzcxUn4558G6NyYWSIvyxFLwaJ93oRc81x
1i9+V8GYRDmu+WLcexMfV3xFnf5WJYUPyberKtYCIcB072IHSiChce1grIz1El/h
Lx3GaPqrOvFGFcmyir/QWuIaRPCreEvxRNMo77QLcsguc9aVjs4MBK1qngw3BWXd
yn1TFULGZ5/zgA02sgwOp53wHAVWH0Fp+OxH4efQTQa0puv4VOMHLQLQHC0/CejL
YKBC7i4l6SRNFp1mOIGuq/OyE8icnJf2CjKIoQQad5U6dhJQRow98YfOCyQrEUvq
uwfeiKEflG4C3DdqSWC3PJPGfej7mkN13XSoaohPxX8WvsMm05TRYPi80FO2KCcT
spIKFyNuVjNAwFNI9P1PZxms0zoOqMCsUCtWFnnMaCcOx7pDpohRJe3AZec5qrdG
zywkdRDVO/Rsl4aC5Y7k1LMJMH56AVWeKuGb933eyZIZKqp1h+HPexkrdIKs4oav
Hy5AQ+VXGHZFT77i5OendM7c/ZpXmOYMeKhIUFDejbMk3R4StadW0k8DzEMMju+a
MfC/yCchMnr8jPlwMFBZnOgLEIO9U8XpfBSqiLMd2LLuZwRHs9K/KbmmQ1MnUAhb
06Yo6nTVqOuiwtGxmk8NTeA72ovjYFlUj7bQ9oZ/cO+CO8psl9AUoEOvqDGTZ9TD
oGlO0ZO4srmjh5RpBvsRoRGNMNc6mqAirZS4W2158aPQdTIeIcnobJaI9fJUynAm
Z/V11bB9U2Gg1Is7lSaHQMKwg/Y/9TW6QEhIIGGRQuqS+xBf4ibClSOAKTQD1n5u
3oFqyuXst3UujE4kgy4TfJuFInTRliaACUbsAyipOPKhPnXvW47fTvbqKgZht4ds
i3PJtAKv66ucvnaTp6vU6PTN59FqSELCOFl4yPrfaoSlWb6HxLIs2t6NrZopKni7
UIr32rMakYIAAU9ulJLHwBcu7uP1xjuFL9VTxj2q+RD/BsSgtNkkxQ1MWqj4rAek
KfbARoIx70RZzbsfhF1qU7R1mT9dB8RETZrprkjmtOm5v9uZJ7mZL5MS78sDjrHD
3GNU33F2VfINc8k6EZnu8u5qr1IKt8IAbXOVAE9RSuYwJpC6E6P/qL9m1/zA5rkm
3jTTVw831zIciaKoYkEvAxQ2ofrFjZ7CV+deWYGZXlit3is7mw8Q3bqcHbcgGRzH
X+CfUDtTY4arQUg5eFf8X9vWsuLL8XKQAZ5w4F0SnCZ92aaboMHtttEPDTBu65YG
xBN5zHzn2SliiBdlGk/HqNXpBlBrsYouU3D7jRCQO2kjxlUlar6eI6NnSO1V2RJW
IXaieslSq2WoO03TPhW1/z2PyzAOxbxLblD+GNGOvh8KvfRXP+RhZX9TZgGE7q3E
Bc2s/xco8seNoE9yE/MX83pdSrVNKH7KO21xPMQkjneAtzfQ0vpXNhSoGFTlGLS3
DJ+EiNfnOwkmrSUZx1vtAXTBjVQo8BACucrRazmLQw+PNvtm1ZSin6OzzKDSBzyt
SWw6wdfu8vs3hf3GbePsaW5Wfg4HLmvdSH1pQjfQ0NL+lBHJRqtxke+frCTaiUZy
K82fBMyueAaoIDRpqQsq6UPvbR0wG2GfGUD4Ot3OvEKsMD9ldIu/yvkcK+EW7673
OK3V4/KwyfRZiEWCbpffV9nHCpohpa4t6H59R+01Pd5RGTHRDYlz4klMPF3Feq1W
ImEAeTRLHGizyyDlKKpN5QY3PiyD6aUCFwOAn6EkfnFCcC5dnwC0YNC0M2l/nkyq
JAZZiqg8j6qREVjf1B9/4GqXhS2zEIFl/p7CL4qbdITVY3sunCxetzFEu2P/BB6d
oSa1+qEqDs1/QL9N+ctKvumVe+3LiLGkzvxT8qAuMwCNcR7Xl8BjnI8d+5wvy0re
/8k20BcC4tnjWVIHH5jLa3h/hKChD2LTRD7K5NAthIJLDter+lP89UGgZwWM0ZbO
wr5Kg1xdxHEt95GSpdtmm3wFoejotdUf2HpO6JP6o2DxlAv8Cw5eEv3ktbqD7Pml
vNqdSugknHnnIUFIAYJj0ff3xOCxU79s5evL8DK+0glJdd2p95nevtw1+b3FxsZR
yhaFu+Usrt8jBrYR5xGRXxQi0wv2z6zGNNxeY8BDtXNr8pPWroEjid/8kbFnIs5F
HO8phjP5k1xI0xqejegjFFRG+QkpFEjBKdbSuILxPPkLi7OjFYAw9aAEiqjb5bdu
5L0EBHnkTZDvIGVvESOkwdR0XT7gbHJW7Moq5vBxnpEPNrcOXit+8UWGmI/1A1I0
xobDQziq+KgFnaNHkyQRIqY064iXy5x0WYJ7E7bn3KCQ9dw3ftgo8r1cpjkdd/kD
I6c0Nbj39IqoH/qPJON/2nrod/qwSa0hddt7pAyxBo62Sh7AfKIOwENIr3VjglLO
aZFbfWFQdb/JRP5/UsFV9xLNU3wEIo7IOOClv2rUJ+F+6b0xB4ItIufCYC5xEioM
Vxn2HWQb8L2JWsJ/ht0DFZs2VycfIKINf9kYWuCwxNO7eiYS3/pKhowqkA/APz0Q
aMvbOZJtUEi+AqS6w19Qm826uwng+o2XlYdXYG/gLHZppq3mu5uejcfatVMKXBGB
2hyvncTT6rfr1WhPLd5jx+nABmLaHt/lDgvLXE3XRqeDNm//qhB+UNkNZyILOQ48
wQfuT+g/WsiOwKvlKXXE1XOXqSPGGwXlGnuRhnu19rWVh9o1RN6eSYrpvmdKMSpa
ih/BBFcFFpW/94pAlMqEILRq2eL5xdx0I4iRUCZwypA7BK7E/Lp4+M+UAhridIvB
dPG7QDRadJ41RIm8mONTdIkPKoaq8eKUiiAk/U/uFYtcCo0iojj9C0rfIJ8JXm0x
KWjZW5529dO8VPh28n3jmQoRmBc1qZLsgeVOXBdWZXfcYUZYt+nQJXzjNlhIMWGZ
ixTUwQczJMq0NvfKSZwYsOxl/lcAoJM4YAV44QDs82JBv7huUw9X548fQKuACxzY
Md4PAa/Hh8pwjrJ4LdYZjq2hN/FGavUW4viCOZHe/1LvjDDUrLB5NSbYrm4RF8TH
S+3cx1CQV26uyq4oYkUNG4XMjPer53uaUpSSLkdEWFcSzcVl/K2GKxm0e20LcWgO
oG+y750KVoqdIOrhNzMewUQ3/YRE2s4A5ymvpnxStlKutIIbWsyOBPy9vtTDGKIJ
KgFLXl36HVZEAb/18lnzg5awUgkmcuVtrJPt2RYSNrj72qwYEvN3FgL79HNhsEvN
TRniNbekTCJBI5+LSlac5iiYUPOVGDu+uux8U2N6dCtIMeTBZ5xA7jBq17ci8DCl
bI6WiIbQeRhZrjgUdedOa8mjBnNq3BqAkSy1XXlRjtRy34KkgQsgI+WT4gBoI06n
wPpTySwzuc864ywCsoKgIDtdRB2olhp/hXW5xm8RvBoKRVlFWWl4G6s4d4Do55a9
dW0fAg/riNo0rpb17+OJ/puNoJ+2yUbsjviaq/1PhRMr/WiFJROeI9gTX4CvacWq
I1PQM8YSGImsJfoeUB01t2Na/gKWqfTmZt+Z+1LBumYvkmSQbypOTd3SfVSUFB6n
lePlZal35BrmUZIXnoSLYBoG9jP9z4L5AR+iPfiD89mvA7LAvVOSzuulnk7Ima0U
T4ATXIESPRkpsfCvL9pvXHN5dCMBKF7X0DnKS3I7ZUC1wGt95rpp6eDw7U1xA+sJ
3g+m/ZgqMP73DBudAq9LPOzqdlQS3CNeRTBiMA49rpyMMwJU+qUapZaRF+a9aewk
h6HQ3JO6T/aNXAaHrD8s/xYum9cTHh3eRBLWecIySVqKZZ79SEGKVxFNT6FdEOvD
xFeAUK3rp7oc2hgTF2JMDA8UONr8e7drekcIR1m6+wMr0VS8jF6z5rDCMeMNMdNw
aYbtzwE9q0BZ2G3ceDYwMCZhnPSl7H4oYIGXPGSM1xlfnnpCe2L6aLB7BwAjukiz
n3ekqyhiEznItuPSi3PSw52gCUoQVxrj2TpaOxHD8UvE3bzMRR2WDswVqaNceG5O
3D+1IBbC6y4jAw6M9uTQGQ7ZEAnIdnxyg+OqGq3IS56Uk8HHH9yLuBaEtg9kDqaL
NzvQnv6pq9ik6PmUSTbHfNO6WPXef+WqRiHvP5NnKeb/F4r4ozhMKnOt9XoQ5mNZ
LpgQt6rXqHfM1w8Fw/bmR/HOYnCnqaTxg7pXdjZk5psLINniQIwQhnaZYA9WGuXP
0U8Z1DxGxlEjmap/FQjFMp5JE9rjYMNL0+R+Lhp0ppsUIo3MuiX6NDPK27PkJPCh
kyEFp8NvhO4fpHrVf9xxuFZWvSapL1a65po5TTHrg2fHJbAWA5e1PxM61Vz4eVKU
5yHbfkztgZ1YYYcVfnEDPc393+yADQzHTTwdyKlI+Mg5ruUjs5NHcJnk7We719x2
DJSkjOPegHTlTqDPjYYbOtV9Dh7QR1awJuxEQhqWa/DH1OK1EeT0kKmBd1HIYoY9
fb2mZmyxUH/iDa9luy0vEkt1uwWjFUxG+0rwhQY3HW0hWC4+E1ZRzuiEta0aXhd2
LQw/YTK7grf9Z0UQaKwzNlzete+aU1Cc+4gOZPy6m+Jt3bbQcnsNVTWybR016Mb/
fDyjBaITOJgz8Bifncm1X3lqV1LDqs9iMLPf4h1M+gWvLm2OjCDdb1U/Kb0cWjbA
imSg1E1YKyxvWDMdU1aWkY8t7DXQK0Tv1kYXv0pNfaGJTcYvdzgEXX6keH/I/D77
TkxYN3C73eNjLSM3xNeFAgWm7OpPgA30Oh76T1pOgKBe+be6QuBFBYJ2796FlBgX
xm/K2hSREB1eFXmJXA8aKKAgej0MUlAINO7uNT5EqTWSogzsQbEsbzYIwSGBKfXh
b5t2/fssT/7MN9Yo09kkAa/+RErFs6RF4Y7FqEwU/1+7YtKN/GeMBJohECM4tiYq
wyLyqxoFjJiauPX1da06m7y9SrxMLfXFvNJH1wcyt4m5/qecNb9LFQSpNi8jWO0E
3zp4fy9xlotEc9RhMb/yP35xeDRfn/Hzvuzb7kKeVgZ7DGvXrGXBNc+mib5Mr8iK
sF85mJAraq3B2uaNW1wbAT+8WdrPNJnSW74Nd6qEpm5eheb4hpFSCcPtBBYuJN8M
O2cyUtHH31sSVe0jG91u7BEIizjju9Grtt2vxapfk6p18Wniaow+F+DzumwHjIkr
jg9c81zSfvWARZ5+CK8HJEzoJW/6ioWauY67NjlPJHGBgEtq8cVqelVb1cQi2Ke9
bPtbsQE/R1BVjQfy1u7WJemKcWKMQHddg/jOnfaFCv9DTKBcuXn2qtGBqxRWMXb1
4MKTKHERVV5QV1XBoZi33nMCaSLhruaql/HNmJOvUeL9oDsXbpHgjNN+W/j1jM8e
3W9qsr8Vr/97k6YtDgyTisgBupZKja+6MfmFWy3Ce8zbBZXZ3Hdurl9/02NaFZ3D
X4r3dFQ1lCNn+HnwDZtlCShGjhLKc/qo7f1m1hwln42+EVgEVZYCbN1JFq/tGiSS
BtXupKLanXccHY8iOw3XF5ho0QTqD8hgXt/E2UZQtHxpGg3kWM3kdr0NDEzL8IGd
hH5uh0UIyrZ87uDLeO4az5j1xALjSs6vFjSdnmhy3kLeNRUpABHllZ81SDj3Nwim
vsXPglXa0KOKa6sPzfP/1dTgDMQh4tc8WD5KL9NdNAtS/6JlVpochvIPY6IwFRSi
T+fOnB47E7CO3Y/1RJE94Aj17f2zZVIYHvycrfCZzFDdC3q7vT38FC5SaZho3tPX
D917LhrlpXc7ucBs2tGg05vaW1VaaZTl63S6GxjayA3oZDBiwiU5gqnFAZVXzrip
UMotOMSmhCILJDMpbuD9lIkj5+qW3iWNB+5iQ2I/m9FPxpoxt6xpksHw7/bHceNd
G1pttcKcRXG3TgFeYoSGWMwaOweBrJRXdnVT6lihYXaVAEiVn1OLzdx4fppjWN0l
eNOXMMnpmrgdUdqxsPHLTQyyo8H9NW9oSAJqt5LQ2QfOf1ii03KJ/ocECjBdM1p5
W+FkgW5o6dkM8L/dafc7IwFQMt57cPMgc/ygR6yvZgXQOJtubzq/Igp6UgUGzPdk
tJPuGRL9/KHSViCjsJPsu7QoR3EFMdI90mZ+IOmLdJBt6cbhN+MqDjio+bUTX7iV
uu5s6Am4MT1kV5KukPUoSE/hIMzZgI/TqmaFR+/qjg/y5ohZ8aOdVc1XvxuvvJvT
3LeNpn+iP5bj8l6jBQMXInj10TwOhTWmR4VQwuk+e+vSkgq54/r2zFG06B/6IaiD
FyE8S38AJm4vDgjtPexDbCaMHslOB+21xaXmpPUyb/+Nh0KR3qgflHuf9/M5njcW
taajOJGlp5Ji1XdlnEbm+jZTxt6aV6j+GUrU2UwM+C0oH61eX0N/PIkkN6HGkYWB
vjE1m8vXXE4mGdceWCXigmbJMvQZdBcuyAHyz1I+Colg24pIEhQ430qD2pZqrSwP
K/qyKC7cfHLrnTrUPzeMB1DXxOnRdUEHq0NFPMt2/dTf3Y7jDdIdtgP+OFmDpl3/
ZG//ZjL/f6ItldXIdZzw76yohnyMjQBky/1nJ9sa3H6fM2w/KI5ZWoO4NRzWLrgV
vI/zPMRuTUBaLeQCmmb4LMvbyRwCnJFmm8myXMTm6L536Y/Qqx4/LLifO++bKunW
lCDAMOapDAbRaFJuSRIFxuI7xzMnz7SbD5Tcd++vLI0YAfUztHlTBqTR9pZv8sq/
ejKfAQfjzGqPI/ZvG6EIyYQwVVzv5iSdGglu3Z0JRYkWJz7FXIySs8zvubbqqfTC
VCE3PP4Ehn50lLm/6SuABdFIkh4qrBgADTQ9q7x7mfYtETIYBfBVkFz/vvRt5aw4
IEimjT6mWKui3ZWNFv+C/KE2OvrRECqU2PvtQkb9q27zGui+oDMPP7PsruGl+L5W
LWugQMEKHve14JcXK48tgiQZpRAnltz79YigBJaG2cxNUG5PUiqLAYA2418wEtro
3HEEK5X9rvOz6u5NltBTEyLhL+XL+e8CZpTLJPkrzY4qwXT4wjGqQfV48x+L9bCD
yV6aaNELBFMGoCan732Tfl0gOL1A/PG0qJF08hWvhs4KIzuA6o/vTbOp1wDz+Ip4
gLqKsyIh/1L9Ag2Qjxb973dpccOENKVr9V6G2UuCMbAcOQ+vr5GN0HcTj40AySrw
l0Zt+nXtWtK68bVWSNTgJLgAj8usS9edJRRm8HevR1uFXEymnatXr9+TttJaLcdl
GQImM17w1rdwj708Xj7SBfV2UmUAo7Q6bv6ubDj2E2lPGyfhXmiJhxLPlBbmxLXO
hqA9S35jzVkzvyjvAxv9aB3VNS4r+/E2quOno1oBQHzK4hmcQ3zbGAE1etyCy0JP
J/Tj2BlaiaRsiVYhl6EGu+ACHwa2Ma5VMtQ1FPlTIK1zXRubKRURD4Ur0E9yA4C7
EZCwkobmu+7aSxdtWQfFWizbIszZFHtCaDfk5nZZPSybdBwK0HYv0xbfzBWryphV
GjiIT37RuDuC0a6Rd2urlxD/i5ukKFU1hHbkbj0LcLTDE56Flyh+e0NECyvX0ygk
rHxZUkp3mcw90Fd/8Z+Tvx3xr63zZvVEpIFctOSdrxiWZFhJyHLfO4NCI4L/flwg
HgGftWZgIHS8THhxTVVIo3/uxn1XpafIT2v/YHhfrrCsoq/NSzX4d9WRTXW4Eq1G
83/NOtS9Sn1FMlR0X2jZ5cPIo+012M3uOjmlYkLhGAKlp1aBCDG0kpb/gGybY4Bi
itbAqK8KmYBSs0OIQdlOcK56p+4zrwylPmALAaO2wU4/ZtKUX5j825g5SUAJzL6e
bCOGRdEcEk1b90rCu/5n4Wk35vN5cajcwkywBKn6wxfo43rDLZiQUVGufKvVSWot
icEb6HfjGOxlVs7jZ3iQjjZPk49F4+LVmGXyPjY0q6Bpshy05SJmJ2jm9BVnGdkp
HGuNWfZZ6sdIMKbjbPXsMDpwqo5EmkNDabBgzDLWTOl00t5DHlx/Gkr+ZcRJ8g9h
h8dQ0l+5wa1oJYD5CdArFq8TEF5JE70qn4r73wpiL5PPmsGnNsN4QLF0pn9e0u9x
anHFMA2+ard0P5sxCKWzjxyY0tvF4olhVbuECy2aWtRVsmT59qg2rvatkVOpkDZi
VNgIQSk7FlKu9Ebocj7D0hUiHdMw1u2sOGWduq7/ulv3+74oMz6mSE9y8FpM44mo
0+yfwtNyzN/dB8a28zipBqVKfbFcVaw76wbafhMUzTMvfJTlS3i9TTi1vVwLlaKy
5VJXRELPU0CsqXobAfZ4vKTUoFWKdcxRNKtYtKYJbHYpwCj08zi5MAZZwtDhU1H4
MPfuj838CZId0W8/hBS8Y3EiLajCnou79RKskEXjgVySa3VIXupRQT1ktKmmXzHv
AbbBmz2O7QcbbnzbhnDOCeLNvyifSmywbNqhnpsFnjEQuw/yJ5vc2mL3FRNjesnn
T/+7LGScZ1BLejFzCd95PaWM4cpn9vlWnbMaT30zxPRBbA+epamM58b8+09g8NhE
prZjVu9YHhk9XOGCLzSvwJ0yyKCxvirenSQqr0m9mBo/XWlsh4TL0pHW1zkOeRo6
v4BSQurgt0AnB5f7s6ji7Mlqx4i9fY+kjXfTGzCRA6XHRVERvANMWROZ7DerwNl2
IPvqaGRHGz6ambg/EQxQkAkrv+nqvipJM1BMr2mGDGaf5JwBnMw+JoakwLAReNLx
jGshFnED4FrrjHnJzpJKPddrumOrv2aPAjEeA4DRQ9BEdG6JH0LdoMSjA9z1jmKp
XsBSioda8oFVHBff5ie0WRIS7uZ+cXBr5EBfAMX2vhNrKHM/L/n6qVdjkZKOuyI/
/okCe45dCNpeGAF0ZE8sonpu7hZqfygCfeoAbwD0VFCfTx1VYFe9cDseQcuNC46Q
YNHAX/88ubvp+nmn7Y/WdElM6LBmSYZFrZ3Ah8Sm4yDCeWAxI/Xi1U7UMoKLJxuG
8awq5wdikVaAz26cPp+/rwGm8+by6Uw/f7CBIbyxaIEzxmjqKRL4UBfV5WhN5hon
u+EwfM6/xiX7wpKuT8w82U3Sx8CKNcWnadVQnR8Q9bkJmt4evyNXB7JoH962XzGN
RBjfAJX5A/pVgcFaI2tSu6Y73n947fz0tNwu/H3Sru67OHugINmEVfR7c8d9uvFU
ooM1eWkeOhFBZQDldkB7R9Gko7rg+kUb3N1FQpnxx5U8WUtfSiH8L0+91XecX/g+
gnIOLTMedH8Yr24wVoccUezfz0hBFJD/sIe7Y18G0OspEexvBvzZd4SLGSXJ8YjA
F96c5bDq4SU+FDeIJmseF53X8X4fJIwySuUUOv4aeu8HxB3ynPwNDD1OkPrl3Vnl
yTuFANFU2rrQ/d4Heyk3VriiMKPUohz3OA7kMKTUTsiGMOPDJ0A5n84FM6DZrPHB
8+YYMrVj8kMvEl5xUVd6LsDmAuWGo6PnMiJIq7ISeCo40l7NMfz7SlgZYHnM1eVb
4Okro7QY6+nXGV7MZ3vR5EDTAUDwD1J8D75DCxHRAAX/lfYYDuyJKf9GZ8BZ2vFK
iWHvZjkggTDB2rYQJv1jIivtMyrgp9whccu1Pm5lBe2ZvmkqQLiREF3Sfy0FTXlX
6PBCt0bL9vV3PK9T4896f9K3fsIb9OrkJ95peTlU2yIrOcAS5Uu++sC9SVFhNhwK
BJOJbSmmTYVQBaQ4hkoIIX+t2YVZbXxE83j4fUeINRWY5KNskPLp3L5eD5M6PIUS
1pr7pWxTufoLjbhjid6Q4FhjZjgcO23jnyCEtRnViMxVgqGvMmP+cMR94UMUrFgF
TlFPXFyA4NjGGq++p8QQtj4QHOSuOFxZJMUDmEl81TsvH7HfrQjeGvQUAdU7phlk
7j4tEr+DO//GuhRKl1n+G5HlJPT0qVauLrxvnijEAXBtGtSDG+IJxlQtwPMdnNdl
8aY6bixilETxsqII9Mmp2x/z+nFNyqNak7p8laeHfpNNZJBt6VRSA6fB1nsb3inD
7GenMnAvg8gXo0X2QcRcpZP0Uqa8RTlslwRc7/xtu2G9EaOUSLtOfGzZP+XvEW9R
+Fv+eqEH/QSJhSpXIpFDrtMTmM0pT7OdtDHmI7/lMjSANoAxNBDFsgqEelUUoTHh
9kqrKK7tvGQsglSC+/MnSIX0+auVE/dEXQUsXMkTjTrbWV4jo4wejnLdpIx36wUZ
+yRMZcq/lqbZh1PIpuFnX5h2lKNVJ6KthqxTzlp4ft0mC/GUzpzQNDPWWLfSVw0O
MkxMjgz9FAzqpuNlofi9UGLjHQApEUkDA7axPUQbLOKCxU92/eyI/HdAU3wQxYm3
38GEEGJ6RjxHwe8d94pP7EEafW4AA95HOPn0upkbTVZot83VaEmES2DKRoSfgHMy
K0jqx4FjN0QSNCyTBvLGdossRBcjjpCM3aiZJAZhX1SMImaC253rCW58ScwyHOtD
Uhxc+p2a0nL4DzgjqNCSkbA+xlIP7IUOVkO0NFf2C5dz3IogYqeCGYxLTNpdMWhB
Fba+up/Ioi5bF5FTpp5vr6c8F21mEIfPwZeYQhQ+Tpx/9csrvUyMIJIOTG8B/VYH
kFr8tOliWBCl2EfcSFTjooMRrT8XSviN658GKqUJvZ/Vwsv7B/SUnDnYPjglBzLt
hXGjguZMkFV8Tr6wiyV+6KZZRnirUQhHAh4RpA00MUu1PwryI/gdFWWM+kZH7jy7
6T4Ya+0vHhEYs0XC5O7RNYgRJGD0tSm7LM9Zoz2JfL7qePc0JdGk7CHiITBEfESD
VUaybbckiIlhE4VreXtMEsUvwdlVl7fF8PLSHLQSmE5nAi9mFMS8H7Lq20rh+oYq
JUsv86lNV97feL5Wf395ZJbPdFJZ5M4ZY+LpYlX7Ozy97hx/IePHotqAmrJlzO1a
SU+AUSZgg8u9FV5190BE2RAdj3X8hykND+QisQsRXubO9PYEWctNC9sQGICbFdvZ
wnXQgprwM87mRkjonH7N4uJMmFxLEZHQNdUE6wewC/QK2uMjHstEJYnHkdGGoyN8
LRYSWkBUb3T8JICZnJQRuC01e0HHF/M7S7iimru2VAax69RZ9hyxKymtk2KT7ugK
wrS+Iya7di9EpAveWxIOPzSbf8gcNyJkwreIJRads9mm0pM24za/sEL9xZ0S6lCQ
v2RjZIMGxAFdOg3LHTiIuQvdYXesEhfsO+9LfRXEYQHDw6AYrWDdAMLqmCKJULXQ
MatSL7PwJZ7JOJVsmoV5A7UorCo05FhSq1xQgXlULWnnK4wA1C1EEI3P490xKqKf
IJjLR5/1Tyyjkbwux2G3/OvA0TTVeglM6Gtcb8XW064g1WZ1burMusCZJQrN0SPZ
h487C6HBds1mSgO18UAkJU3RcZygni0tlVrH9TKnrOG8Iwg1Avujz0UoighrxYRW
1PTzrTjaz6Pv9ErOIJrDcs+A/iO4zWcCA2Ewzcr+K1d6eNev+9IJJJtLY+ZHdgtb
TbDx9/RazECcyMFcNX0t1iCjViruADNfQbALrjqT7ghc5WrHAq1a6HOfTO4VC5mc
27WQBQFmtYr80t3oStB1MKkOeYtqLs42ok3O8mn2S/4+5xeuHXsUP45Cj4J9QE/B
5JiqBlZYhHmMy72yp7A6SdCOOOQ74aiipJNnw6kd+UlOLlJAfDKmBbPCTmEdVuP/
WHTvxwnNru1d0Qdgw9N+72TKgN3HP3t0CrddS53SgxcukpCedJCi5+tNeEZ0ZEgW
Cwe8BZW/IQu9mh4GfQvvwXOF1ukPlVkT+RcCPcJ+zLefV5d391ZFrT4MZ9z6v92L
sHznLaUFz9MPnVwTEOCiXb/no6RN3YiKLhxo9d97diD+TifgdrF3kL8cv9xuluUm
keH/7z5HAQBvddhSDWOtfsicZnAya/dj6ANlceHdjqRQPYEa91XBtOkY5SrfYO5N
ZpByLWIq+19dN9OzmjMAzP+xlbTUDLERxRPzx1mAZhE6O9f60MtNsLqjHFTEb/vZ
kFYuVdRFjX1F9xcOhUQYVG8TGydLmv3S7Gdr2yP4eIaJfUeLd+kF8Dlqy5ZMkBGx
rnnkwzEUVn7h0M/mR2CpEL+iL42Y6MOkmpiO9Ld7ozoqhuKN1v63NeUXw6DvjvN+
C1J38jydxHdF1XalI67ynsAZmhcKwv5TnZdoybhAoo0mH3v7PbJDT/acZKUAX1ST
eMsNQ5COhavKVabyFwHNcCcshWXAzKct5yQ85+z1s7eKfoGyXKwuvsaYur5HWJhT
kBJhJ8hlndMWCZtb90JRFswYfad4SEkAvgQ+e7IQ7xch2Qhs98gnbLHdTkK93Lut
H7ZsobRQV3gyNe/MiNGZI3QGvvIILm/KeI8+QmSseAQPXhE9ajx2/xASwm1vTe9F
jjU1c6fXucZMl8Vz2gMazMPPkb+QTjEZ6lGyWh/iNMfVqBezZFxd5XL/nqCQrLbM
Z5seCOEI+aLBYpGZ4vAofjNJkW9Wt9+Ch3sjQJDhVAA2MuGJqbpuesVjHlubXk50
4YSWTN7obcWrxxXeMoDVEI2F5XpBGfuddVnUgSvcWMWpCDIBqeXfnyj4H8go4PFi
Qatw7ASNkBFdS7/Xa3Uh9baVR4+cNUBIg4o+PJBD1vwOLLrbKFlUSgOnqPyDLkzC
3+/+Y+YJ7aJxIBf8vib89NieVSaLJxmtxxMf8GUOItpdtyW5Z3aUDLY0YMKGDeAy
QkppE/OLdLhPLyhPizfnJ8Gl9EV4abn9vqPmUEtxjl0BU424R31DtFErOdu1lS3k
ohWk14PJgOWZxokxDs0saZTm99qoOsVdtSgDbZtQyOnE7M2HqVg9SvIHN5O4L6W9
Ng3Bh9BmV+4trkUUGSvASjqLucogL+MbFRb844vMk8i5X4bRT6o15fVT1fF5T2cF
yajoN1/HodaUk6G/fZ+nmO5+uQu44oVxXxnMHJFuE6guMUZZCEQC3XsrG/x89UgM
VhjdQPXrHPfLXLFURxJA1wgjdExE9PSVkBxgX0YdfNDE8SGJ5NDmkN2ObDdjTnPM
4FbvblYjirdgr+eKI2KuFdrNOPAJ4CGKpmtCTvX4MNio8xHECjRMvINO2VctrOcx
HWfHAiDRN8hACgn8Sz3NSqTs6nxzAkR4Y/xJ1NeVnVH7en+z+0aJOwOwNuwQn0cA
00JNlzbJ1fvXAGuask5XuaIWWuDyhuw26U41msILP2fc/rqfILn92WwQvTrbKOJd
cTd1vA02RBT7CxmUJH8IH4hrWHogKI+t5wk1PG19mVuH0m8DlTvg8X/BeV3KxJgP
s/EV26V7Hw6CcnePFJ4Mi3Wvp5KZDNF3DX+pNiH4lo7K/K36T57XkYxWqXhPN+zq
/0sX37d6H95khyrdhS4B2esWY2U9xO0TOHijhQiRNEeGzRb12n/n7Kk8xrOj+9+I
ksazrrkOSmlB889T4m4bRJB3+VfUD6QaT1xZL9veWV6bUmEF/98Ge86vsTXDQN2H
nHizBQamU0sTnYrZaOC0HB4CND5x1aoTqQtxipb3mCRVy+D9bY9NEVJY1AlpnJbV
1MKfHLDRbmw9TxwIiKq51dgPUplxOoHF0gBMqIhbMcsPurLD5FitUql8li1rZzS2
eOhv6t++zqtondlujrGk0Ye8OitLSBAo1cEcCzVWojsr3esVBttfBiv4hQeuMAlV
6NKTSadFBkKVIRJnvTzESy03mM2jZh650CLN8VQd2bmiqmYk6COu7vxWmIeMY0Vt
0HsbqBSBGCTjH+ZpEEjDeMsTmvQgIT0iJSFSwR5kQb7tIVlqsKI4HqPm6X9bekuA
ipp+4MeGgyoh0De/imiJCRnPkZxJojxvM+77dpcKdYJCFX01OCC+RMrDtj3z0FMU
lXSkYnWa2uto7wPHR9WfGwL+CGU2qlUox24eG0dj024j0tdoSoI3ScXEVW9ug1Lb
CJyPfBpEATebynyA/DBNxR4Py6QaQxj+DQQEVZ9BG8MLjRPRCejfdF1EZNIDAbCL
0ifpCl/1DTNxu7rVjIvRBX45v0DPkkv5+6VZbSSGauDAu81AS92TUhU7iA1PFGxg
OA9bLpWhiT72J8qF9aro3jV2WxAAPrWkx9lR9SLoBeJKTzxP3zwNaRXkYuKzkbG3
KGL7s+nI9TK87BwXFLeZIAcyoM7yTX49nbUfiVRUtxe9rn112D0gyFhipnCg8UR0
6OTTvPUI82YYyzGYbF+qqI4hPJWtM8IW5PMwB976V0GwtD9cP1O7WQ83t7lZzIaJ
+X5vViDcizXczdjlYQ8dXQ4aiwj9UhndWHuyPudDcz7U3OKOkJoWnJaDqWj6vNUR
hhZCteuVMkabHO6YGuq4U7Vy7cHcJ/xu2QU5k3KJCatXwba0EkXl7NADzVY7unHu
MMsKkXNl153o72hqq6fJFB3q5/b64DNiUhrMKb48HEihoDqTGp+5PGAYsP9iQHoV
nhGLr2aE5Hvm/iLmzETz2zYf/HelYOIx6rViAoh4VPvRXaQWgwONsIG3HLFYeIG/
dtvQW+pVHWIRPAFE448OBffNBjGSR0Sbj9PUR3nu+stp733zaC4sKv2C17/2wuN/
Z4Gl0JGtJMB/4KM1biqP/Repe0/sYk/ykfrjPSKlaS2CVv1jhkxKDEqtYuuMBPsN
F1nCjjB1KfDOrXGseH/v7qNK8BkQ4lG2unpentCNj+FtFA96urtRhXS+d9lu2DE4
7c0t2GnA5NyNa329Yw1MxK4B3vpWGTJZzIlbgFu/9bZg07AyZyLzckmCwoRZfkPX
tcrUFhLIoGRXxISILGFJIijvG203a/nPu1S9D3al3qsIGbNzWzDyKm9cQwlolGT5
nYJ6l8d8tr+4oTAR0uKUCjiVcvvDhBvvwyRgpRMDG8xanlYj7AqSRHR9HgpIWRzW
+h5HZ/kG/RexQ4OrkZlN5Kp/Vypf5CvNtcasp5we9uyVqbHBctfq4CicfzhBcpvI
Cq8wBw5nlHTcH5MvkLFv7gBoQiO7AZlB5u1H27lkSLsqwq9ln0z0A9DnNj2ZHiT9
HpwzOrQ63shE/4oFNrF2iiZmXAJE0XrX0A3DrZ4fKzNV9m/eLWJsEu1b4Cx1qFU7
8xwAq1Fifmp/57Iz8GiWR1wwolNWPQm7CxQfLUd56A4v6oheI0ynzD+tO68uN4CB
2zcffzIC1/YxdvvuWIo8J9VluuPBMp5IqbzlOnTJaJpD4QwwbZF07/0fL4pwC7kW
CC1ptyJzsoSrLqgFq4RpA72LXnsj0VwC5Ds7UIt902xMHtLKPGybWcDMqjnnSfXR
vDw5807/ioKWGw5S9/30ll6alamz6O2uD1EQGo5sv+Y3B4zpHL1trLVqpzfNZPre
sRxBiurRjPmBAds1669HojTfNc7P221VSyhQptuX7ivNIfciWt+pSQPC3w/IB0v7
lGhDUPYE4ccPFQqDQcfYchlTCgInkkRp3G2mGm6c/MpWRNtRD0ReI5lZuBJri2wX
6MG4q/CzOrbb0tU9bdsyeE32S3xVFSTZxIjAsvLL32Ay+ceGbIMFKKDsF+yeCVnj
vVi575XvvMv8RAO2icN96C7Okndqm3seKyHzk5nIok/cfye8UD+evbX8p1DmjO6q
nENcClluf/NRSqPHXx2OoFhVKC7xbkgDzHibgzaFpAFYM9U4jQ9YSEGQg0ReTFar
5SLxtR6Tm6dcisPv+ikD0Se50EUBLnp/VtNZentO5cVtnGSkTU0VTBgccr0cDfsD
wAZ0Rq8PI7dfE9lA9HoWQ2jPuS5gLPdMqgt99zMuWWwm1Vsb+GYi3U5nU8WxJSdA
dcF4+hKMkOPoTa98adFrCdUDUogpr33hvTKl9otN9+Fz8SWVR+GwtWiqHxvEW4vF
0TTfTlwwlHI6aUi2rJdfyBTemAhgtnhruazKo0bBCkSG6tvJYGdxCVc9LiqipeRm
2OwGK+90dx1yg4d7jPO8k5aq63MsR3+DJAbyWQl9Uz+yPckrWTLqgrsifFBPSRp4
SraiojdEQ5ICUUKzZD0njyMRWFdd9RM19YMCskLKbKa9mNMojNvVIV9vbhS8C3o3
C19ynHoNfhh/0yZhqG4CaDQaUsBk1NwuJ/OsquJD2dsl+iW5krPybN5bAePnnt1D
MKFmcwD/8uc6JlP1a3FJF5HcbPHttTLe6KWnLeKK3eQPQWsMfFzIt8zN7gfO/I9f
As1KAuMQMOjRU6RcvcZIFMsjYNuaE9WRTe/PbUwnnc5fvtROSQC4LdZWpox1eHep
Ns/jN8lKrzVxGftLvS0L1UcvvCdvSs4DQaD+ZwmDROrrsrDQbS6ubq2xhqK9SCLE
50t6M0nLHnmGlo3GZkU5gb4NvYJrNAKlvbafqi5cJf5NeSAJXNuk84cHs0JXRrme
Rs2UMkHlelRqNKjPTYxnrvSARBqCh1nlD1sL99mwWNSRLGTAk3R8/Pz6pGWRSlbQ
71vh/WHvv1NAP789QNfbltvt0dFF2aHL2zvoxtKqn/+tT3z1SZ/Hg6YOGI+H3+pY
3/qv8eN8DbCwUm5RfLumq7nG07HSbre+kNfPBsWbFR5XkUkVBu2qSZXKcNp2KTOd
KfYsN2eOu0JfL5EJt/Req1lnH9k8KPLCsuYlkaGiJvomNuCEyJtYYDPFt4Ha8SVj
fIERFpAg9xjd3M8X+6Esz8NNGNGYeInhs5OfA2fuY+lhOoyI2iC5slQrueF5IUbM
PQDdhYajboer3vyyUJSdq+2yccPUJeXiCvs28DirdIsABkDSkmWUJ7pgvXLul7Xy
Yv/LClXMOogBjvliVAnTlQFFwaHtpX2F7Hn4zT7HE5DdWaIfH1pITqdpjkCDOs95
fPpdVsEbydipU0lnYkwZ1NM+QW05YQUrGQbUURaNnLT2KIhb8tjTgXrzTaHWDa6J
op5Yf3uxhH3PWOnBrxpzYZmI87sH4tyEehrKW6QYDh+s1biLNuGyuahwp1WHxMk0
3q8ij3cGHj70kJmLIDsYUdVX6OcWAAxUD4k9obDm3y6ZdNNe28QekCqAQAM1pc52
Wm5Yj78K/f96mRiayXuZqGvRIX7aSWlI5kCHwSC2pk/Vg4ePm1rpdF4o5vWghZ8i
q3CyAeGl8TzRAsPsLqlkUnycVdNGegYIf0HN71oXd6Hmamu2DafGqVOmpoiuvMBF
oSApkf8ua+t9fimBN5tn+zsOSVLcs+/k/QSgcDD4BGuo2NVRM63O6iWbXnKNI0TN
jxAS0PV4ToyiMO1a8+t7b7CpCd6fHZbocVjI5Lk5Qy/527oGjrz4BwRGDG2JU6Tt
5mn+qDZuHJIaz6e/o/DuDk2n6c/svhvPRr/b+4Dqb3iiMseFM1uz+/FYRysAK56o
8TBjwLsLn0krkbq6SycOqB17KFW3Uf9CTXWB6v6zOzWFd/OhGUkw2ybK/4mCJ2ra
s9Pr6mttTl+PPTAYn+vX/oYCkjXZf0P0fLb5dpTQDVk62T1tf6f5Ww0pgC8GLMcp
FLmjAH+ewSDY7e3h32azd682hMJblLmOTA+KzsmLqfKnEpI3jzx5nuzEpCVOHlBr
dPetv3xyMHQb35B+hB0rWfmNVSiyLpJD8bRZW6vBxDMXL/dwM6IQsX7F0+ID4pz7
QmtIUNySvkSjb61GvMWo+Qpio5eYrmnZixVeD90fxlwBA8/e9qTjdOAHRkqasI3D
A5E3TV7rfhOEzyqKbO7cvr/qx6SZI5WNGZ8oX1jvDdUohXuxxgb/GgML1kYG9aWh
4uFA8kyxArh7hRo5ILZvAXPFP5S8WVfW7OYggOspA2RdC7HyapIFmyXJaObrV7l4
uaH3If7t9sXamHUDXHElU822d/6NbMDXlmGFOaUwZei/VHHh+Isz9MQCjLgjxQJF
drDtAtBlQHZELLrhOsLr4lFMlBWWpRVAdxYy8cpLKwK4W55mccLoqFn3IxS6cJ36
OHAoIiNXt5TQOpVs514vT71T0iuAG1aLGBvOueRinp6J3Fg3f3hfvfjRB2R4jiX1
b9R7jrv9N16tx/Njf/KAOYyDGukluYA+FUX9mYJ6BHHNsHRJY47t5CqDuuP2fGZy
V9jBulS4Q7rGcIHS8p7XMBx4t0bVdGgZwzVEY/AA+SPWsAtVqo+vVaXge9dJIFQZ
CMUyUNw4PDVq2A7T5coxpXz8qH9Ofg3F7GVRQaIgpN2IksZvcZhZIcmNpctQhGqP
6tFNIqG3543i99By17qcus1Pd7hDyL+yKUS00tiB7fMrgv2BW8NTLVY4B2zTl8Zk
tIFRiktW1vj1pmyTxsJ+f1qn9UriKsInLrE68/Th0KE2DnX+TZ7EG3hNuKtp7WPW
yUHwZUV+EcHEVr/Upnic5B0o4nB5CFXuoa/OMa93KKxe9lDGCh9IKfSdg1UVtunI
jDoNHv6jOOa1lRfEflb++KfGdRCcnn8WhsLT8j3x37I6J4cv1tQAfUHJCXbNjodx
RGGkhdAYzXHl/CDXhe+j9LFteh0aT2X9bvXkfYzH1yf8UkWQPdugk0/sIks7c18G
oHkgqTIjeernmcZDtshboTqPVBNssg8dyiCL5pV3AVC2MMnwwnnnbM+WlyW3nxw/
0occSo3/O/x2b1rAR3CA0sQPN21ovM6r+Ob70Iu4DCOc7uTOzC3KvNDs4znAP9E1
ME1W52CEtYYv/yCU8NTY+c87R8fr/TlkaFzHGJ4D73XKOJGy8HaAeb6ELPjVAlVn
9WrHDoUxSdON13ZG9qIX2p8ng1Zxqe7lCSaaHsZyx321ThA3AYmjOtvH4kQDOkr0
jYjUmzLiH36BssT8hGUURZh1Q09FjJ1jonxWWZeJZAwwYwZ0gf5gALBLRuIYpINV
YZjwCVJ2bow0o+PpaJtVVPxSug4F5n6xy9GkZ5+qpj5kD0XG6uHc+/wiT0jMRSmm
7zvrR5H/Bw4jITjweriNtVbWjh/2f+jiuRk+cBOrSlT5ZL0PWoQdijZMdi/DLbkH
8YvUkF3GNEiJ0ht8hs7fxLd8JoxwV4ObWyZzLBlqQU/Gdidb9MIM5TDxwwmz7AjN
SHWL4L3agpMYX+wreAkjQdTxOjX7rAzU7RNpgqNf3D+6SHGerLTzF1i2WPF8X1Zi
xcKVysXY5m/62IqHQIrOaMHmDCgZYM53WRK+Of5zI921TLljj0Ml22WTH6DhrPPb
rsn+25v8z2lfzSvgXPLQT2/QzMyml6Hepqpg5YqGv7EzfpnGAR8EXhHR8HJzdfDJ
OV1xcC4/QoFhNT1zqWuEXYKeD+Id2EbubA/993nC61Y88VuaN+j6raGlmfGytJGC
mVm4BxlZPudRF6FcLPqhlYl4yVdkvrm19NzEvp++N4GL5S2buEIFIpk+CFK63Fi+
rPCdwOQRJ7qJbcvU7+yonRmlr/C6B96mnspu9Fb3HLKNLjnGG4pKpLfEUvXyOWzq
mZquBmzz+3EHb9Q7+a89hJ1SxoyoZkXjMQAzj/aPi2rWqwP9ujd+Ez8r/Uqmm7AW
5OjFNF+FG9mGuaZ42YUnS46ikwR+ACmnJDOJLiMGNxlsd7dt10Uy734fTjcDU9hf
UD9+TEjxnl4QCiPxGYPj0jaaIcyb8VCl/tIL0hf2RuJYtsmK+0gtuWKulEc4RPIL
PGws5Q5e62v+M/FJFEMA/GXp0wiCT5uL1hBoDeDTyO9TfHo+csJ7PBSu4WI1f7dc
SMlr/yb9g4wcTfZh45OPckU7ocxnfFy8lKWRarmtMdAeY1TubCtqm21Dc/jPWzI/
Wb6QUA1oJXKZf7TN9Mo6HaWU8bnvQeGSq/3hF88dBnwUIuZbpxqRdfDxO45vzWRg
0VpeFLEz3miMdGYpDAf397Cqt2aeSi/Z64HEPsaZyQJpvHDM1ZqHNrWbxpgu0YGk
a5M00cB2s3yymoyt0AhSANOu+sYKTv/JkXcAYRHP3QW30HwIqttZ+af/qnJ5nJT+
5+JtlJjsBqLWi9Oxh4sI01s4Cv89XiIHSptQqAigFYXDABx2m+nj+RTbVmeSxM1Q
xZC97ssnufR5Zr7pPLmPkJgZTdXmVT2oGKmI/kWsaebdFV0Xh8cM3/IYAaEjFN0m
PUCQELmLHfoqDooh9KRyeaygVtBUxqtuBqHexPL2V7NcN7IoZqydweVItDWJ4Mxf
dyrqQ0YFp2YbiDSgQfX+nCAFogksMSv9QNmFeClPFUCGhrjGNcijG94I6wmSRkiI
HsCiSaUalOpzIegQyV5Syc+Ts3er+Lc8LcvPN3MgR+ixjovNhiOkTjOLQktc+9Os
bhxjhlKDEgsYU501gPPqHYHvhjWaJfFJt3+2qCOQ9L/6SJ2FikUwWM34YjS8MSqv
hqt/ox2FplpBFmRuWcqw9vi4pNOMSNyHm8kuBHjm7neI7ARlxG3PaKNsh5DY5UF1
Z9wxwvVORZgq5lGXn1t2HkV0mWDF6q337aJR/ad4nubJ+adXT6O0IO7f3+XWoWdt
S9EBylVxiR1wIKxQhBB7ABpaD48d64f4LuhDBC6USDxcGSJXXeAc/pPRO0IUNmrq
gunYoMl5PAiLJP+Mlwn47tdI6w/ezGzQfki8DXWxe7/c5+V3mSOejNtfSv8WeFo9
LkYIUVYlUS5ih3DH4rTyujrm3/y59MBiZtsrCpyhII3GnDjJQEMgN1j6buavIKyO
frihS0F6u2RZrrja9CywA9s2VUNiykqwjYuYQRnGyla4sKHc1EDNBgHIvAK4NMZn
E6bNLi4Re2+U67zvtGm2sCVB/7U0eTOChtsquXelsn+iehErpViEVNtAr2LWCEZd
2x/wa5C2RvJtmZ7Ef4qXMi9LlYVamCIVMLP2U8uMfNhaAxpDBl0qNdf3QTqY1+0m
7wOy/WC7iMigmFOBOvyRg2l9EeS8SFYGOIdJt2XtuHgMeSJeeJpNji6IsKv4y7hA
vYoQdPzRXw8LC00c2cPzblR+m55Q3LQMABu4pc1+6NoLIxT7kj3ooxda7kyg9ori
xg9a6+k3voeBNJlU8P6h5rg7nC4kCHg2iX/kYId4oIpniNdcv4mHSLaRcyaNfi1w
KC+zD1HWDhmg1LDbgfcV7LXzCqcOmGSKPC9KfRYaTYGw4awETpzmnxzXZ26nXlTC
Poo2dVaDCKpKJRwX94ucdgLQAPIaCa1+5VJPP8iALIQjZlTNMFwzRzSwKv2Nt/lK
rJtY+JDjsLi3XFfZULhheioGd0lVyKpxBwZ3L+lqwkwJN2f3/yjSTqYMh9A2qVVq
c7sx5uI7PEjrrCA8Dqp+j8TxLLg23sUX4U5EF9JkNI2gdCwcARvyCwTh9y8sHAx1
ZgjkxYWeHa7zT9zUnzU8EFQIi6CnQeWmxO1w+Rhpd2w//XhknGzkh7YncfSWEzzI
F1QL10M/DwuYtnioTOsgoooIxQ73Os6Q7BmJWBro9F4NPm2QkMhBzGlTdF7Mry03
dRd96NhOrbTUiLHpwStqWChGLOox4W6WxFjJgL8Wf5jOQj8Dz6hyujoRxNfhBPT7
1q48d1ynQMlIOHrwpgKDTS2PbHfm1QAaKsM3A92r6951R8iQMZVDt6KDnCVe1zui
NqbJg0qGuiNZxepMKEfAVvqB3hn7li464RKvFmieGVRUu3M946+o1mgcHjU1RLYQ
dBP1od5Dw4B9ZNeMwHbTAWc+5s0ByR9pVmV5rTEoQmIV+zb2BcQubKYqRrP0ylzj
I8WcdCrUtHUDvL9flWD72TwS0wUvm4DEsFv4ORvWRzHYTJ1CSJllQ1lavDeehsb1
KgHOPVBtCpXHn0VSbgULpYaOIibXPLHh2X/ygy1UFxM3jlhEL4jp4f7gzkSGnWHn
5vTCZIBz0QYOR/i33GLtxOuES6Qz2AgFHjq2As1fXyER+i0pAFvA6RXm5Xbaa7/3
iyvp2r/2WTGbCIh+Hw8L54s2wKAEj1t02Ro9x5XKM1vYVIiXj2gfERwf6vPyCc/O
GL75fcSjBS7Yatg2JBLKJTc2FJ39fbWQ2ceGigxHRI0tRsp4DzYuDaI4BJzeKFWe
UicY4IjKGrGS69x6wlfM/q5bAtEdKYku+tAtDQivgBe93k4bOdvLP5Ynzk+gADWE
+PwabNy6TyqchVkYV8u4nguOy7ivFkHGCsEKP6rdF5RlNvo9wzcTTDyv/CKIJkbQ
NxyR0bwcJeIj8HwroW0M/nv0Zq0Qv73YHUretqzmeAVX6X1RYI8NdCFnGOxl6SWG
AylJdWTIyVakL/D02OkXibqtlwD3dow84Bx8Jo7NgsqiDB21QI7Jx1tdsr8EmAe9
HDKmgC09TkeqF79HJszR7qJafajqZUei55J9eBg89q6fCx1tTgcprFRupegRcd0y
Sjd1lip802lXY0Syr+D6c9v9aBtpcwY39NKKx3dujgHi7tlzZxjwbWnr7FWcNqix
noUoF/yae5A7KsS5ieWjRjpb2gI6pZTUfz82TWF14ShVWa/BuFWaYlUpbq8avxxo
PwlSPvUeM1FJa1NrBXsbLyTWsK6QrDUu9LsRaZOWgIJjuUqCtdOKD+gPAW3W/LSz
4VUNTxgpVamjpzmcKKBxr0xvpZ/8sD73gMk8TBaWxIYxaaaKHAkH285y4dQzxXel
QyQ4Pwvo3YMJfjimy+id5pC3AIBpAayG5KO2XY4Jxpd6y8c/ouisolCBKZnAg+3e
D0Xs4olK731CTwOT6RB9pnRapcxlHokUMItrAy1+u5v+O7BKSUDHZuX/cJg8CHG3
T/Ti3fJnjEoZsOztrUOFX1dyZ5KlWCSX7yeJQ5CDuRdamwQ3gRdpo0YQHDnsJ5D+
Pp1OM5QmdDIrqI82OeG2Ynz9TsYp0pxwzKtfKxdxi/KJD1uIiLLnh6ygnwIJsuNu
weEteeEmre3Mf1LuhGdOyPlsHNW/ys84xSkr6kT6jX1CEHjdOl9KphCwkEvDBh9J
+bB+6bOsUGGFDEm6fyDOyKT4u0+6f0fbwFpmHe+07KloVmSCjnbsxDol+18bUAd6
SksDgWbCUJaXBC3J1TLCQ5jH9KqmF/fs0rGgC6pWs5Hq5sPrXYL+OF+qA2B5kX29
MAXTr7twZTsDDc3PAXVZHlMty8aHptc60SStY4gaAzVHKXDA0JyCI7olTHeKDsuj
iXJuxXs9qjQ8hN4hLv+5POUmvGCFgv2TEi84OcuaNVLdmtWm6rTqatgPKr8zYOq/
LTYX56mpGatNjI4kSeAWQ16Vk4xFxS54q0p7kPl2Yj5gXPidzYcIHnoPmavByia/
ZRQZD2jp6Wm8yKY2EhmHhAkUIcpi13fsEnDyUZzRYEfJXkJ5OSnsA9GSaZqwTzlH
WH5+yye9+QX9l1vxVuXrM4jYIM1AglULoOk393ueb5PEb5Iktuwtoy8yp3Pg7fRg
ubH0uawruFj/YmvIF0ourPGjjFcJD1JnYgoSrqBFv3HfKE8ZY7VQGwLvD9sIPG0Y
zzfLlGRtbBRprHMJXJHCRtQPmvQ8+p7l/ybgvi+0gIcno+iCoBoB0+M5Z8R6w6OF
gtNrBs7bFEe0SDv5f1jGjNfMzxMZElHUgUzNTKvofhp+hU7pJ08xigGUC8MjrotN
TCZLxdyAYG/exG6ZgXrKMB1gOkZ3StKjoLKs31EciC5/YyDbWWCzA06gaK0aUEX7
93mvDVv23mYbmsnCkqPToQwZfhuVztfQCSxsec15Y+lN/RLOuqZDkb103+4lZLIv
+U/c5W7SNPZN6m3PruXgATShGGOkT21URTtqKD+v93DzJ60stYH7kgLuN1dpTOMP
ee3VYNoHp3zquVxHNcmG8xEdqcbbgHH2gryhNhWswD1FTMaYAyU8wcpBnaC4rFIz
eM42os4cgYNsCftMjdZRkrUSCG49AZmEYzrVrbbxRzkjl9NZDqv1crTtgOI4ujgI
mwJCJCqQDHiSce+sc63lx5N91042m15oP3QLQm1pojN7iTcT8f5453/LyNn8jzQj
McY3tDSvdI+e3a5wvWWbMkdXvDMAc8qIrWOg2017OYCcfBrRvnST4zG06LTHTM1e
+RhmgIzwXpBKxgCPwM6zO4kQvuUAtojFv5FebPoc6ebdy4Bb5zBRpgMwxNa1DG+J
ooVJD2pVyqWCcLyIA95LAm/IQc7t/lLSI2DpRbZcFmz8ZPsRKDZzQdnA+iV8AgjB
71aqnIRWcWmVzyBnClzl4wsoZfCAPI5DndEBAh57zT94+qmS9KxMXD608e2elHvq
7Jp+CTmfs5hSMoC+u6EG8JVwiUCzaslXPkZhfpbeaX5OQKdATly8nOJKXKD+EnCY
iUBbFOCJq9bHOPLsdTmAHzY4wuw9tcHse/9iDne6X83F0YqlJ9+PmohcvJuEaORv
bnd8g1H7nFDATUWFgwy6lRZQcIXiaP/eY6kxkJzVEq42HXUfuoOTVlqPqCFQspFE
+bGLdTNtLx2KI8vazRqB3xULcVdR9hX6845bpRoPBunC/Ih8S/eKAyOcmefgvmj6
xUDyt2XhlT6zCPRtaLsL5qtmdNB6dFRJZcd4Gj7hcpd6k8dAJlzbiPFgzJms1leS
sdd61mpEvuFc+KLhCCjhgaZRhTQuhsL4QKlehuFZXXTA4gMeuKq9+/EPZRWzN7Lf
0d0YUn4eBnqQ/i1HTcRutxmlC+xyFdnRAQm7h7Te1b2Z9mMHqp55C/VH40bZsplI
/lwwYfs5I86D291Tnms6+mO/HjCU9nvBn2w5BWAAekuYj7OUxD5vuA4K8R/NN6dQ
M3vUQjBRSmODMVLwBBxYKaSCYqEPhFclbmh14Ms+wF5Z1xZqoVNgy6n5JNu7Ztdi
ySQf5qFGbjyqjsIDfkHdQhJZ/t8Hw1VXHcIOjigqv1w1XsW8VkQS6QnUhZO8vjma
o5JO0i6tyoC7OO0JqHleXNfpRp+/2IZA9nH2e220IPxuci+roCiMNOsufGOY+0xb
ehJk7S9H0BVMF3RVZXi+mtd3D0bAj+jbGrtQ1RSRA1gP4RbEL8cIMds+9iK6BfrU
/VWxL+oonDn4WRYSVAwI9c/A3ZnIgyMu17b8gIKK3yNJVhOhXn1SHok0BFSZWjQF
PKlDt4FsYsdDJftquXwB6gwLasBftS43OlOTsR5FijFOr5PIvbCPjvQC3sXBe2E5
thQGTfZlLkabKzvA5o2hlo6c1tOZ4Nj76kp29P1lMJWO07hN8rxnLxUZ2bduTEVR
AlM5ABbOAEJW2lyHtLC04WMHPFL3lYT7cKC7OEXJ5LaCi41PGUTW1wFbvh0qrf5S
q/Utf6b5Zj7xLkyHK/5scZRbrRDKUWHjdc4yfFaVtp2pYy2+jHHzHpTWJmaUlv/I
hi9w7St2ohsbCQOTXkH/TpkL3lmqHE4AHdBAoXi1S1p+CF/0M2ofmQApdh7S+GS3
4oVFsGlSRfvNpE5DVUPylEB5jrLoSPTDUwqOA4xKa4mv0GQnsagFCelI1BjqK5VJ
X/qpZVPhRCqjSAmVCdHYZpdAFj9uosANflvJLaw7Y62RTmIOU4vYCrGR09jTnhFZ
b2evr8Rd6trQsHRBaPtVlYELt55/XBEIjRueifkj873hgWz0D+Q1wCUYlhOKKoRf
3sYv6sG+GG17lNjH1ovtB75rDGf+H1rScp4pbthTZcEZrzCeJGoxgUS7VBG6P+lG
hepONP7QWo6XOyAUkM5i0a6WM9fdaMKOHWq/JWEZIIEoF1om6bEp4Z7h4H2FwF8E
qqp7RtS/OS0UZJTw4o9KJGv958/2x4bjvcoZc81fxJCB9jJlb0bJ79urJqekz+tS
JZWXQ1RDbkswO8YrzooFbSkZZ86uWan8s6Fxb3ST48Xe7KOwpi+leUUw/bj6TjmU
C2Um8smmlXRbE0VmnmZorrDjkXmFsVZKWu9CQ/p854N/kFlETrQ5iMHgVqbTsS7D
hLK5rvhF1uRi5yvDekxr+kL5PLHH8llTgZkrfoZcE4zVtPuR2MOSsjwZ6Gyt9y1Q
zW1fOYncF9d4i9x0cKeQH/8X9p2sdXbtSEjtRPuxLDMMPW5D5CbFFZKJ0c0qWwwa
YAoDhpjLKDQcKYLncEYJbuFrUlvP29UcBKpOaINlDmGJnBZQgUkBZ169abfKWFqQ
NZCBBJiYwgWveaUPUhbi2TRPL9s/hRL1nMJ72SnG/kBcRDlaxjL4LGsXDqLWyj3q
MsAekJCURSztEMtZAd+oQihCULjpPh56FBonu27hkE2Bbc5skyrLLjNA3j/mwYsM
TbDH3ZXdG1sUkt+cyKLGuY9Brq+Vm5ft0110kLXFIU/GCsfcOyljyzf1QQVy22g7
1QwHm9j1+oHO8KeYFjQTQCsGELxZwH12Mt3+2X7CtWosaqIWiZPQUt85dqsLcvYl
QKnxLEniW3f/PIeTLJ7s+gCVjinYXadxIJfHmgGv3/vx1zahdX+/ZJTHuKNZSinP
ohiOOh2VGTgwHGPQygEBAiKpnNzwEcL8F3RGpH1I3JZuN6ZxcdFbeYJo2dcfGs+i
D15+XHlQRcnC/OB/P6nBZEkraWbTBdfCWne1k5hQ7tJ2/a4RJpqIhhtbTduBaljo
XnLfTQd7g6TjO1u8BLDl6CK7gEt9q/yX+wfsEfT5MOioz9g0+6kdNoyTtmuYEU6l
Y9DKxmCzcL47OKW8G/U5t1K9eUe3MWlReWDTQIEbCuxassvHYCBFalGytgjUdFkX
cT21M251CS4tNzoyQ6pmi90c0oyIRU5xmyrzet5RGTHILP5LCeA2Lj73QV5XyfJP
bNOc0Y99ZyjWOajYukEWE9Du1s+GLzdozGCeQrGkX+ybJs2Tge2ZRd9j4FQgxaDU
MQ8cPKT+EIRjALnwzsRsKLeztyq9rzIjX5bDbKnpt/yEdyJS0qE9775OBzaoh+da
lvADC6eHej8B7vqmjDsL2hhklZJndi5cySbSRnaYKGm0gUGifIh+ucRDEOGqKbLR
1BMo2Q01CZ19JE7jh4fbCtzvlg1LpPyBtMP4GxKcwPRObuyTC5Zg70ynBgq1z0yh
pVtTEJv4vkdHTjz8+nxww3bNxQ6RswX0F3mmImEfcSIyinfpbCo2gZeN1X3wxeQ7
+Yw1F2aM8UGEFbUNL2NnP0yBryHavhs2FSAJ43VBDx5hengLlovAJ0Zp38PMBSHU
GKVt/gE9xgX60nFmqa64UmcMNnpiEYK1YFMPY9yUyYmanXEsa9C6tYCfN58gxDED
ySjaz1pfgeGwH7kGF915dnrLdYlLTHRlU1lU651xIfrHnZGot6SaGeFYyfuLHLBP
f47YcSKu0i3KvRKHqFTeQcyknE8RwSExFRnx5E8eSsxsEUGS2Z9bZUVSIPjGWS2q
LeCm8rwTAMyLgvvYurqC5w8VNrxmZq5Hd2elQIGpJB/4aeUFLA4+8Szh3FAp+xDj
W2BlrOONxZzhx9MzZdvwM2OkSyDMRH15ZmH5bUwXzvsATyNkSMbT25NHauNphqPf
xMS5Blkt9bLbVCa6YRhUPT9eKHvy3I0m0OHj78OiQZI27qh81SfplyYhaKKD63cm
yptqrzBSjysPONyWt1mX6J9tgzm/xuVsV/AVEEiPs1G66/xIlKtQ7lMgLof1hTGH
UgEP6SlnjL7R9MyczDasQGjnx0X3entPLNKRXQlajQAzyiMP0mhvyZ8Bnzntzkj1
JL65PW2kRrlkXkrlA1dCRL4h/4v9khZu65ECFRoMaEOimcNHogX9Ak8V2y/+ZChr
WdUh/lDfpAqj3a5OMYBCBEJSVNsggVksJeijtW7Ih/ZOuIL1rbFRil8Z6rg/Pz/2
GYK9l9iGR0qiT9HOAJVwloAU0eCzhVp7UpxsvqDyTO2e3DLeVw7CUmOOjdGPymuE
h70VMLHPNGqwLBfKScQCm+gFWQXQdVe4g0FEnGgwg+c68x0Aw+BTrLS8hihIlob5
wpl/8NegS5Annw1aif5yV274j+lftlfSZLaKbFbcooiU3DfXHTqsQMIcSnOUUFpU
zHwzK8vGmr+IOsdlhqHcSes0SIAFdVkI096LeLjybwFLifS3zaa7OBZwCHbisdgi
bUh4hOb+r5qDtmBH36EXWdwEfBQwKRw4aSTxVjD7Kt3CVZYqZnHkRNp5iqb2bcZD
Db/yhdrUpRGBGrijUppMfg0bOZ0wIcePjm8uEfRISLvy1jkye7NvMB0lTC7dOhjp
Js2cN8G1T8nxQRjrddqCWIJ7h1P2NqX4ZoUAZHdXntl4mEetbJrR3CC7kA+Shw76
Mx4RSSoGcSoGTE+lPN44CUOyeTHEBa/BKizTgGPodRIoUbxgd83UGjMYEVpxQCyN
PhUdW169EoOpqP/gc5D3xdGtRdZ2+e4xON/QfJfBYB4QwZppRQm+/QUCnbYaHUHm
Co98VfLlkijSNu7xFbCQFkp5ct/Jf1RzuXHAA4BrAnoifma/fJmnNEXgsadqq9QG
mCNLYNeADixcZpTz6pjnmNb01pPz5qgZW+d2BU/Kgj6m3XLKQ9XrH27vgO8N4KyN
0MZPequVDESPBzTt9jlzoVwRk9WzZx7S7CEM7VqSTBN6psQoBP2Gq4ktSbx0/27X
s3Sn0iOWfqpcZjYgl0XNlHnAHHWN2OmgomUEN4/d0rwEy2SnG03j+F+RMa7A8gmN
kf91sVEVwdz5+6SoFqp7RzCSzpEuBuLMuqxG1GNB9NGx8Qs4SXlZxMDs9yoEh7r4
1Tzbix78Z0L5J5Ju19Sv8O6nmW5EI/6LfMg7CAyyBAvQWjh+aFkwmAxIf2sPFV9w
sb6BDUu0abQUh/I9jlT2AfopRDbUZCMvzmRo/DKhVmkffjYGqu3ARt5B72H4iEMb
3wmEfKWltLeOCuKuAfMcB8gwXYJSYfWRHgTdevs4T7rPK9bjupsOAoEGu/j+sZxt
ddHbw3gl9XPqXQ/JH9hx43jQrfTMcAo+XeheLENv0dhlSyGCzQXeDFiXA/sv242r
2D5j1Y4aB0SYbIYhDa+TnE8zSbsW7hK5GLsCyYp2NNyOjAApqOl0Fg480R8afx89
mJ3QcOdwUG7AwbbBK32lpqKUFfZ9I0yLtryQQitpQz0WOPZtrSoKjKfh/wNsEukb
LOEltGJ/1UK8MHYHwSWTYOpJi7TjedOQ4unoj8ZlN+uhkeb2gxGxV7ms4h1yhDts
K+VaKOR7PSD/TUugMQ8Z1mH7qEqCruq+abwMIAVmfm1XWN6ayDXR2b47gK5Q1jfL
O9KFPPmvjA/aGFPAu1rsRuq+kjPxFSy3fHTcUmixgyMniHZEtVJpxDlCHjTDCHO4
X/vgZQ/Fqjix8Jzky6H6kJaW/5Sw0FBI6tKkB/RaoC37GiA10rWuka4qBya3YLPU
LuMBSm0LDuxCqHbpsm5c4Nk2njTC4eKdOpIJ/2OgHK/vjkmJXue+dpz62KqF1CwD
p3Y2giaXkvgesGwVAB8QUuBKeKu917cTDe9nznsriYeZDDL2lGgue+/Qt0PESu20
miI63urwb4ruEIcp6zSQOriZpYM6AyGRPuBH4ns0Q+pmdP4//3WDhVhpvM6rduDU
9k8ySUh47og8pPJe1OkVrMunep6MvuMDHfLdotnQf1KjBceBcs7d/50hSXtkCbEc
SXEZibcOF5cz8g1UW5PBsLAqUBUGKzoNHA9M1H0tUNkoJw5oRqRUpdYE12QXV62c
UG6yzooFNKLIup87Pp/X9oTVq4Z82sZZv6HtZxB+Bp616hpt/2cnFJYY+4BWDX+Z
r0g9AOsc06ihySRKTwMrXRKIuG3V0Vv6URhqo5fjTb0I7tWj/Ouut9g0oEY9JO2K
33J1tWmYbITP6p1P9qE7BTUfyTa1JQP7kOenBt+uT6w6Cfs7jOCnhEeIN0RlkaUW
zQlMGzSq1G5W0KA6ZxDlqi8TnqreHUd6o/tcSyHVsw4DsRIaS2etyZEwaBEj1TTT
SUlm/TAQnABwtODlaj4rLs0wtc1PWj28m78az5VfnxVKXOnaszkSTEa7kDKW5/eJ
in3H/B+CXv3kYqwUBoMjBH0FfKtsaGb8V4BhqlT+Akcby9zAgmvy/uqU92IFfneg
cFboOrEhwdSFjMogB/Hg+GPUN+pk6AtPhzbF/SY/S2XaWCdMjDEpYt2KK9XVKLPv
bw+aEEBt26hS+1e6v6gjWaLQm0tCLnM7iUV9rMnMEyprfUcat2spBs33kqbrZVpr
S+hBpirznN60OKqidGa9gam/UVn++zfhZUZ0J5Yh6V3KTGl0bVp5A5O02FgHHtch
k7UxZTRn6gMdUUHBxX0LJi72kPPSLsXqabjOgk16gs6F/LT+b/5NC/3diiGZtf2k
Lo+TUeOslXzc0fKCHf3Haq32kwUQEO6OObYCUQMFs63ZEVFc/du1E20euSHZFqEB
ruVa5qYMWQVTjFy7XU1qKjG/Y8Hh29Ghu1prrQ0a3212Vp1j2Wtx2icm8Xqj4CBp
i6Lpmcqb40h4SJl/TLxQLvR1LNaDL6Ek2knTId6iVl1tQg6ZRgyfQYnssa2uhMsE
ZOdVi+Ii44xpZ8FlEt/HTiToeLiicUnY7dpX2W7V24IP0XxVTtK9VYzmo6Fx28S7
EkA3XMdg4O4ZIRQCyRr/EWXmU4xNPTiQNx6kSm+a+FQDSzs9YtrOwDNfJgdUlNMa
M6f17QrEYAK+hPfj/jvDkOtBn9d7sUd+Rfzmk9FL2Bq7AkwrUzA82ICY8tFoZrdR
LnSTNxdwIeFeijKs2EhqkSG3VGje/enzOLeJHAGqyOIIuPp7WLJC6m89+eCgWJLn
20vEbsbYXBwXV55dNkFIWCVa3haSkeATuqVL9CR3TzRlUpRTa2jX6ootE3U15Mhn
t06yNuR/i1qxEZJMlAngnf2I02MiLmEut/yI0N9R1rWsWnhrKkoFn54fAahCYUyc
S07L4MbHYMdMINgj/sAFrlhQBBbhQDPJ1sDMyIu/pgAyxpgIBx5zaBRkR/QYm2Ot
vAwYe+vI3uRarfuzUzzj56yZkbN//cV5oJn9SM607uBtMlovNZ9pnhemEbOxf0GN
e2BKZabrOd+75YhqAQeNc92467TnZXMVsIFrLN363HT9D2ONUJw+HqtYSWFIN35g
+N3266cRLj90rsSLOxZpjpHATDAoQl4bolbKgEk5iNy4sU+mY09eQlH9ObittLIL
Tew+f7Gb5Zk+A4PXWOBd1P9Myo6dDCJEProj87lw9VZVv7iuWQRjEToBp9mMaToA
XXKtIVlr9RLSGLcWKOeINpSqqZWDOF11cN0+WltUhx75MMm8AnNdM8nblVtSPt9m
0OIEYmpQq0S7GUjtADAmVLLz8LqSxrXRuu8aQr3OhIppK84SM+gzWKtBMelp5MId
8OXlvOrT4L9tjlBWi4/tlOVdz2bhKfWVeyGMDQxWh6l8JBAqoEs/zU+KFAHIsAOG
WLmhmX4ZHeyzi5Mx3TBHTUTk86Brzp90LP5MKmLLBK1KXAls232B+qOpzWiVcRQW
mkOjlrous22VfLNP+Pz6jQc1G0uS/uis7W6KH+DAT6eoF7Eh3yp6xYm0ejwbqY3/
1R8cQGZO0m6LCl+lSuLfKQicy0fLfghJ2YVtA2/P4jmQzSQQxPrzfSHERf+tEMFV
oTXOvgrBVuqSqD7uc04xb71dRpg7DNCQzh3eQyJG9Z9l/tsXCwLP2iTIUOpLXCRF
PEfKWDPvMTqTS0ALTU+porFz0hq4aWodkXsfM+jYrzUWTSA3zmA8FeTlDu+asnLD
ljd0b3mTreMkCAk5RnHqVieYggyHi5pQcUt0iYqRVAV+KfSIzk+A5YIO5ZE33DHh
91wZ1Pu3BvatTYGG4qtC8TXWaAIR6bhOZ8PSNbPZ9SJTSTa8GmWuo7dcFaZ4GKCU
zXWMGv/kzTVTE9FZ/VPi8ucFtEpKec8lXD9EZwTRWLXPEM5Q+JZH5DJaS3+RK+bK
SzLb4AduE6DzO3WQpaf91zlRqE2wWo8ai5ndaKtiSp24zKybwjJA1MnqMiBWo2uv
bT2zvHClxyjrJ4UgiPrPGA4D+jjqhMlekiEMLA3mT4WGmTSA6x0hbNkfLGx9SxOI
+dmhN1+IpK2Jc0hhfqWgi2sKUZrbhjR0DXIQtQvXsXYESOgApyPZCZQTIAaYKp7d
Ty89PvJKxxhbYgV97JgsF9OI5LbKYgv852sve8jbOP1DrUMpZ1PwXaZkHOwVm1BI
dDSg6qKpYr4oLr/BjSAioCRj0AECLvuyMqpMLlwXkmWY98g0jayt/UQwpGvgkY8Y
KJ+AqXk+GIpsK80zGn7Ud2fy+191wCGKtiqvA0aYv6X2WnFYG4NjsWsM+Np9fcLm
8mCNCbkvK8WPJBQc7Uik2uLIAvQuNoWDzJ5KWxXA437S9wBYxhGJcTkzJ4XTZ1Xq
3/MZmeb1PgG9xsVSTaL2oLjXciqX9Dn9icYkKiXl8s//h1TYW06jWTRN2YaoGSpx
jlLwRTahAHna73LrvPDMs4+wAZrxM7hhT2qFFHop4cFyDPuYu1dcLBw4eVlStSlM
Wjte2uoF9ETVFsWeJ/IjAgYYtjZlsHbi2Qu8bLYtvVbmVxHUsqgplnQ/6+uhLuK/
6dd4ni2b+rqUeU6CEKLiBTaiVxP49kNlUBlRQwryn70GFyKujMFw62h4NcciRYWM
RVV2MLe2/8o/zILk11WYJFtpEYp5xKib6AqiW8Jdzw0xUCD5vU2MP7CrBXbJvk9y
Mqny2jB1zm/gSmmEifXW1u4ceP6JL0SA6JrPxZ8AL/KPLZIg7Xq9ELjRp8iEdb7H
XmOsIaOjQJDUvgd94F7RkGURWU3hNNu6LL1mHZ3d+5mrMLk5ZqrTFYNdomEzUv2I
FGh5IhBBUNooVWHgz69NKISyFMzey6GBQSfnl02wnObtIJiMeMZU89yXwDsPrOcB
cMyJp5lMINCcjy1WD8ZTVsq20h6S7VJx0nkpMOxG6AVi4PyCBuvQqkWtw4lzrDXo
zAtrrj6euM8nYQTo4F7cKpkSBjGq3wgpQaWZGLqfLLCPbTbn5gh/lCdNWhyubGKi
y+rqcRq1e1sEMp8iqZ/uq0hnOA0kYwEZrFK6hWo5W6XGbPnsraj9IEhkLPnz2EVy
NFgorHt1oBAY3ahFBlHe8mByOlP2KncH9yfbgrN3dDL2py+dkRoChuKdE8XgskVi
7pnBXtTmd1B0phGAlyYKAxwFW5vlq9oMudZSk6yGQWkkni/6XAIllgbBonyxsIPO
j6MPlIhQVq2kc2eRD++O1hKnRe4r2uPP09sjW/CUJSLXQ+vfxmnbCbvy6NE1yhOT
GL4+vsZd2sr3zvij/QOnLOpwH9BWg39J/qS6UMz81OWb79e6xPo6we1lzpEYzPa0
wbYi5bZumzsEillfLNeH4QB8c3Bimc3YBzFU6AVrcwhhmRcicGiuocVeift6VclZ
V+ak2uIrNWuhkpyngRgUFKQcqnqTtIpUts5F8zRJaMtOBEWWUNlVPiSxlKVOxwkA
tTnqNOqcxBegITR0gCBhcmm0cF9Qr1UjXV+OaVzuCzKuUHUJ+W+VDjxD1dwQoubs
K84FSoEIUC5bXWiksAQJNC4PI4DnHkKxeMAUD7TmnBEuRz9qgwFEHTscqCumAeJ1
7bvSHp7yEtveZ0OSwnjvzrR133ZlDAl0s221ZSxaImtnDU0Jv3nxeG29VEaylF/C
BrrOGP1D1HtN6NQbJ0Fv+YTzFznwDPLLt73y1gx0cprK1PLI5z5FWC2hxJED4uaP
XnVE3WscJeRm31GgKex/Lo3DF9suK9cVtO6SvfyTvp6XKQktDj1vIArnuvIsp4lC
d8hgYxcpr+K/BH6dJ2C/b4b/XsN2ZDqm1/MwJy55NiJG1flFxUtZBvlvPT5b+Ac1
zQ5Pde4pjIvfENWs/QGJy1adKCuIVKcDOnunnm4bV9bbby0EQxpWkVSBtwBsWEgI
0K/Mt9YREvuZccsOYsNArcNdC1aeq8Eo5zFpBC3K9NWSQsloUhNUHGRCHgebmd2U
pTNp0PjyPUmBr4MBF+3MOjVeVAZtzxvtcUQ5xmjwBgaIiczqlWDIjTUocx/N5r8q
H7WP2uMGG8sGCy/EGu2RkqLohQnD0DeQ/4Ed1oipHYPna7Ctqup6lA28sk/hT3Bu
J1DcUAxCvpzCs/HfkpzWVa66hoBK29NdvMZcct4syAU+JaxVfQatNFz9scYNazgG
R3FxX+YjzN+Vukw5VxCyXZehtgr9D8ZGZvCI2Mz3Ym1/9QFMhM1IEv+DLLLngOcC
VURgP5fSIJClmYIRHvC0Ill7KuWNPiGUaTL8QPky6D2NEEeGgz3YoB1Uk/HQhfan
D4sNAV9BBGkaD844NEx+8VqgV+aWR4B4b8gR15Gn5T7gndMWrcU2PGkj2vlNGI1E
b5okPy7yHaCcIIzQzQk9Wfi2Wdgd1ubl52BT8IgxIUe4xkC8HryJtvfjH2tDdVDm
Hp/PoOq7NMDXP/svmFtmB08q31Yorn/rePSSs8URrbM9pt6Up4TFpAfRNyONpv3U
iMSsbq0hbvNwNj3Uxo7o8rGcpXpdLGzZimEf2k1u3f+EdRQBzkcbzc6bK/LzNM0c
yspWfX0t5tg485DzwgEOi98hY1L6M+na0tUUOFR3KzQ9ri0IvlJP6+ZrFEHuychZ
kh7XGWh5Ag7LFxh6aTkyWZVFrAH8pVNu4hsTOThtQiEQ1MHUzukQVNECB6jYNxG7
7u/7oDrmhY6HuqA4pMYGeNEgtfeyqFebHtqqcDvQKl2+VrbCJ4tDfztSl/Tp4SRT
6yenaGvSQvOIS7ayaMzXxtIzJWbupuJAaYSuex7BPmEEt+VW6ozT+zb18TavzyrO
B+s0g3hpYzMt4dcBVzzT+lCS43dtr639QkKhx58mT7BgtY5iTF6IVdxeETqB5BFP
EnHSpxoHRywWfoGKza19UGqUYGm8clxo1d3igVxoXisQl65J4DLiSykZtjd3VKvn
YdzAk5DwosF+15dr8o9rvbevQUOcGAmoIR4Xcy00VCx1m0DsK7QtWOVe6vPYDJHd
EnGltIVsF+Vv/MscdhMwx5FY702vuSKE92S//keUeobzwip244ParaW0ijbqW+mH
ZZykW3GqX7AWePcfX65hs7ilaRi8+NT7du9S4rS45AaHQdT2XptFLese2nC6hFs1
SGmYH2YTwlP9Vl65eMsJna2toczY4gokGV4ox9WbeX2cTStvrBrjuIydMwZ6mkh3
IzSVPUUznpDxZZywgjWlWp9FsoOWLmuZ6GTFfSxsu9VMUAJuue5eCHgF1KMfTBSJ
6rNnzO/9/Z7KwtgOlTCxhx37GgWeKQRqGVoWVIB6USH1j++yyS/ZZRYczmxvfx1n
3ZULpI7Vz0XG7YdO7TISsOCWT2kh0ULE035jWv4374PUxij7PO4Ju+t9nkDdC0V0
NoHv8VrXh78gQ4KgU+HS0MsFaaQGWosfRsoEZCcE8BK3Bzij/Pzt7K2sbS0QxNdH
UWR5eR1mAIbP6K3jAAOwoO2pHj+SgJ3bjTwInfGuwNLN/1gCYUCBQSq7a/yEoiZc
fXgDfB56sS9tTrwGfQkLGvyWHynsir5xQGv4+adp5xDGA16ioJ6X2F26HNfCsAEx
1RlqcdyrpbAgT5sut6THqIjR5+PeUXSKMl4K1u1BXB29WJuWgdPcUOhxwzFGUY45
H1CZImzRJwNr2N3OjLYOsxb3S0B8iP65b5PrjuXW6KBt1KuBRw39N/D3Gisjo5HM
p5ND4gygGrR8meSlKhHoxjKteBYmULYWUhvZxS02r+KzuHS+1f7dcFg7sRG5g9O8
CWKZa4tro2PHfBGsVK394KLiKKw8KJFsSpzDngcRIYpJCPHq+j3eUrAevK1D8/+B
V7saQtlBdwPerhCgzBGLJQmgyI2ntQV6F7U57FLzZSyORGCM6bUFb8MvJptCV88E
pOuBnAFtQeh7s2tAFJFQv4KRthgVOHfJg3y3f+qZdRxf0S261vg4qrodJcecw1jU
NjGG4iJ2HwRAG0wqiRqGhF6C5WXK8ktizFAE4i68bRHRyi7opjtP0KHmxNENilT/
KkZGCm4vbhXFuq00vjHXLRPzGX5LXJbA935FFP363KJyhoCJMeeP9j5KhYHXsrNj
ZnsUHPpCovEzky05l+IsR7NP6e/D220c/ftOryRx5Xz1laj3zwyCL5GdDUeJSmyB
cLZYWO8xAcdRH82MrZz2DXafiAN7AC4GJDPUNT9GbmyTQLgJqJKd7dAFxxCB08Xx
hbXopbOOypvIqlMzCKEzyrcfVylpbvHsTBc42Pv9pF7jIE/mS6vfUa376G4FwrFE
bYxim4MAy0Z5nQe5wTlkkrMbOSrbmPGIA3E8sgTrgR29dQNT5IZ+Hql4Q6e9GhlI
o4EHJoI4naqNzFd3S94QFrHpavAtG1layKAIQKFKfsVXXXzKJ00SSkS25NwVLB52
PLqPTsxuxnhDscJwQPfonfgH0f5fuSSL0cTB/cUzTZDupZmSvZng/26uTTNodWvm
/VgAjdy1DB90kOBofJcgTxUcz1WDUlkpvsCf4BXt2VV24mPxJ4nSZiiXCgYXqWih
Z/fxM3m6n48QW5GcqjtHmOSgtMaL4qy7l0FQDzZMautX7YifRyhw+tUMcWMakvS6
wNizSGXOLxKIBWnVoND30gCASikU0L7+N0yGIBsEpu+y+TcVRXQwe1/gse4jOMxb
tnAAjetqzmv2yr+nLVKoK9pCY8cLsgoL6sOv8FldnDDATn+9tsS4cls0cHBAKKRK
+Cuq4BKLTw9IWKXdHxdFENmOn9j6JfWrmpvSw15L26oZgWhZ4Hn6xc/5thfcH9nz
gtkzmFEqdYuA7vqKR+/YSlAddYTAbYhCweQP6bebrs5i5b723bGaTcjAL3qWdJm7
5AYD0IxemMlFHAx9BR2qQBljS/TOldM0eQZI0H1WSK0BJO/NzLRE2H84R/URph4B
eGykM5oySutFLxD0ccLzng2qW8eIN4ryVimeRkacPfTXo8bh6U/9iEnxl+1B2GE+
p0oj6tMKsDJPpE+nwlh3589kjK/f2emlqAx1w2xUdLcqMOztngbELN15KIuN/ARK
r7n70ktnb1YNMccTLkQy63LgnDgemRKw2BoHZTeHYgQZTtzBdZuHC8CMi7jmnzja
y/NTDRvaXSmkUlKwj7Rj4vbeEDt2GSQQ4Gq24wWQDhZdZBvKuxRseDlZmGauHh6M
e1hvdXZ5mkhYtevyrV1HJ4KWyRjM3EXW5rkmOBEN8WCvXqHqhEI6o5XtkVFztIRW
qMXz4AivFsENTQ3Ur9g7aAUhGdYOR71Xh5sa33ZuwzlWKlpqzuSmCLIN41/rrRiL
vQk42gKAD+ez4fu2/3LOvg0SbuYKguCl9evxZKYHRywRETwrJ576X6MeuHY49asK
/X/e9iETB6A3Z4A09tNTTTjhPWfkzLNB26ugUpkVeGz4K0wn9k4PrEeluBxWxoz8
6w3QN/RxuWiqMVCgy3+Zp8z/wWYUxFs/slU2IDon0U1QSlMnHlVzfam1UAFtkWyb
2XC7cT+ifRtwmIPDxylA2nkgta/NnEz3wgIRbgDWuGwYAfU79IASLS2NpiTgLa1v
/Iqj8L7FNt2C+IGVI05rM+2hXcsYWU5qYUVFM7g+QVCAQ26OOy6CEz0qcnSOk2Z7
kHJguqs1qqNjR5zl+K0wP34Wjw89oYdsxFRe6nmHvNBp9LF1DWAaXwWYQ6pZMIMB
Ou1JRsywDRX11mao4gx0ZvWSRNUJ02zyAIhE0dTn9rukht189i32Jmi4J5dLqfym
ZraFWr3XchA440ZXD2Vfisx60stYPXpAmNVtOnsBJQfN3EkeNc+WRri3aq73W553
4LW/MVeKuSLrYoS/O4uL+4wRUIyqkPwqjPkx22CE/Yw6MJvpYkaRVT/4zZ9rf1jc
ePcYqAWAQGXjkzY9AICojNOPqyznu8VsrO4ugemAcv7e43YDsfqbdUZhC02ZAckE
8boIRRgVfH9vfYhudUJjzFEu05sY3aswnPYKHMpdjDDJsV3viw06WXG+QBQvOO4A
VQ3Hn6ArBRhezUzfcFLH6XHQXZogsu+HVep6Bke69j8ZAgbyew071j4VyIaDNjma
1ddA0I2hHazoXBtVxbYuQjfX8OH20GwIx3SG3+1TAaLlnlLU8UtCZdqEGxnBmqm/
AmpCMzyE3yuvAaz/Gpy/qp4cL4jME821vEH2qkevFaTCpv4KYSaHtkWjKbvlSn7+
tWbkf5V2P7Cu8mjamyk6ysnmhU8kUmAm688GFOtMPlhyksmAlEXLE66Pw9lm2F38
xjHfixHVEsV+PdzOSQto7ZNO4oGn9Ig2/TPUhOvH2u25sSTWzty5KJHdl6FENm8B
CjN3B5vDHTxMfTj/eJ2Rflzx5AExP72+TzkibNACCCJidM5/KjLnhO8SIXXxsvau
E+h5IJ9EalWhTs84PIwF0QDJr+4DeKyGC37kPtDOpt0dgXBMYTafQHPq2XsJwTdv
CVolSkToSFiG3ur3A2PoXRqaXLiae8F/m9cfw+5FxR3miKk3KBvoziZSM1BkB3Ks
Isusdpy+5SAUOIn/YufkixGLU3rhRzVJZZ8khksK1icuvkNPJH6uCdzObXEnxnGc
o4RLXLuaZMirY3AkMWGqn30xTEsiP5pVykwuN4hniMSVS8o1oj4ydfeMPid2Nr7l
hLrTP/3qhb8gWIDj5HurHNnj6Axoq5gLHg7dF28y1c9K7IleC/xYvZdgtN6P3654
eCQrFLuDMEIb+XC6jijG9txGOHtl+VeZVcKD4aEwWKnZBVgXZ3QJ1gVuCrHLhqvJ
pYZdhiczxHtQ9JUsCUgikhSo5OvJQd2RHIjyGfumEjqfwuqEMlhd73h3QO+RXSCE
FN/ojLA/J/2DJuO/PR0DXNamYbcfRKipUS1gBSANCRo1ylx5FfS68KIx55qE9GDG
Nzj55Zkeqq9j2tWJ4SzxF2dHF1V+Qp1UY9VTS9MPBYpaSxcZvr3+mMdHRWFqDamG
mZdSLjNbXo+PLOkzJfQIhBge9lA0GAllZ9TEMEzGlaj/66UKg0YMzfuupARHNq2m
/QgavhhmSRR4shvlIFfwjgknO2cffPoyOkDCQ5Odex9CDRuQElDUf93BwtmRGf1R
K+JC+YHrT2q3YQ1VqMTFGylGDPEe+UtjuJLB9B2CWhIwqDRqGi1Oc3s9iqCADUKz
hhJxVswO5UUeTCwxBKieJu5yn5Aj6sNT4cylSQ45vlD6KUqrg8SxtD1KsSiKqD7U
NBOHk5g4vjKPVtUWpLoiioKABv/ucOuGpcSBl2MkeHDLwtVkfv0qn+F0CU/7NAJf
E8+jYrmmwB0isbsJuwR0UUT4dTcG6iIgEtQes/koP9xUVlobpkJqwGvmkzB00CfJ
jI4VhRE9TDpv9k1muHmkMIRCVNwaXNzHlyf8ao/+UTRcrOkn3NbNj6ZaPCR8Qu9j
ybbF+bLj7Bxay9rss2fUC/aDY56OKJIHEeTC9MeJCHzNVd/8v/9LLLBiZYrpqpfs
lZmopBU4eaPqdPq9rYR+gEMXOQcmygwUBtpX2A8/NxvmklS3b4lxnJ1holVAdYjZ
6Jp+Gy69cCs44Xi4Fv8+KyWtpW2RElcatIAT5lbwAQxf+jTvc+GCQTHJd9IqnSuN
DW7EPtry5HhSNAOGZ2BvExdpJUDU1H4s6GmQmovocNkWj9AyP6CiRThZM5SEeZFG
cE0R/W+5N1SlUtXcHoDM501OokeanqnymQUKN0fqe49sw5D7puSWgCxu1DvVGREk
NaX3WKK1R1BYtDofN2HE5FfynFLL7UO548H0cae/uzokXm6Dlrzz2/w2CKwfYLN5
WupwJ6dj9BIAGa5DT0htqAE/WRKIPc6cs78mHcWU5bc8UxI89cauWfsFKqYOWlpS
0YUX+PrjIUEUCiGj7RJL/mnNB62VmYg51uALQSVwV5DpsKAq5W6P0RyHB7b5LHdW
rL9BKxT0HQoJ80PTL/WslqXadCZEdwyFuFt4ve5Ylpt92ib2/QG/ijvTGBztIAwo
GjSe116YXD2ccyW7QSSnyEZ5CHWJuZ5xuWNVQm+roCta4wVohzIoz5jg+y2KcGGV
EzpV17zalvDDLUNtdMcX5TZx4iiXLeHWJA/G4kNHcQQNR/GtVxwWxRCAKZ19Qcx0
Mb+fC+z7171w+QWE34vGt8vv7M4lV4I+aBrp28uRaxfhacbQ136bptEJ+ozokf5w
giSlq+/DoAYRyLblrpQBeivJeSO6eeVPznR6RTDHLIEWuvh+dKYEiiDleRWA0xvP
7L972WisKqT81vRQdd2rPhzrmsESmaQVKqJgTGJKNAEqr1RVQkmXXUwaJ29qYK7E
0s/EOa8t+bOuiAgPcN2a8ltRNcKjAVzUb05N++L0oHYyRwOQa0ZN3KucsoUssQQp
73xnOgKz1KzxIO1EOs6ObLAGWOrrUkG0kMW7peuzQDmrzeDWdc+xuUyHegQ7Ssnu
rTKzMsCuIdfGNBfczKY6XqicOgAmkh5euv0tVzXQuBwkqEFYt7N1gasjFV0Pc1kv
kFofkrtvaclYlELXIv6vRCquXO0iuVzPdPnjgJTluIEPpUEjPjAx73V9sM/7H8UO
w3jFgnNe7UYJhTx1GRn7AstONulPkJh09f7lstvlNv3Yx9nSRNTZY0R/BiKLx5A6
LvfnK5+y+glKzsD7vS9npwCwD/33Zp7T1sgPXhwnH9lkQW2jOua3IjOw7d54u9N3
w/xu3DGNyKGG5alFbipvCp9g5oSQjtLV2k1ZRYnzrYg9UnePHz/fN1FMZA7Ry85W
VGn47QYPKk22zVrVkB416idRcBW9wsyBq1OIaz3KjoaRwni68Yne7LTqH9ZXTrXj
mJ92Y6psbJFWyZjuIq0vCrtpPzuMcdUhYFX+ttMuY9uPD8n/38LelmmsNu1EcG+e
Jzk2c+//fUTDjFP2cTOqC/5jSirVRP5ljHZt1QqoSV32TUSlI3+tjwB4Y1/UGiU7
Axr73wRRkGl8YFLwi13jOekvCXhGIRCwx3xxuv8U0z2tBnVTQSZK85HSXuZizfOa
Kqas5JXwdQczNlqBiMoFTs7fCKARrxRm6cl6ur3oYQvTgk4+bDoqdI0hHXtmzxuK
lHh2qVlp0fctzwejwUNeY2kiSLw6PBMjYP24OtEAD5U5WGc4f2yY84n70yvJGuM3
LjM77llOF8aZg6Ov+vRjYbP+4mYKmJrKs+m1vgS4WodY79tZMRvqMK7JPpZFzFXo
mHx7y6+VoKYjizIzy1eRN4Ywnb1Xwr4pACUa0GHmP6P0UuxghScmHXk7DdZZCiqQ
XUxjcnaJL2gTY+V652Yi54BxOVMa9VDNzGgHbRqEjbsf9MVozW/qdgOvlW9sHKOs
GDM6/gLiDkjBmNjvI/h71ULOoz3KgaA0TQoUo/UmLMTDtHcDV9E+S2S8JtzBnC3/
1YD4LS8LjGdw+l8f5Q3QvgsVEYEK6iB4xdfPC+3LC9AQ9TSktLARE5/75ljw+13p
s4xpsxPzuGlKEtxcZD2vv3QS5fpS9a/BKE+yFRq1E8fHs1klMDnQkL9VMP/7LAc2
Gug/z/KAft1ym/aJBRPLxz6a6xJmZ+MChrYkQchzDYjIdPIsoZBSKolCYuQGxxHl
bSYo3zbo4Sv9smTNWgv8ziq47vryKqtakfU6atIDGtcTwcJWSjpSMllK1vkiXfTe
bdTYGjqDxxvxkG1SizzF9JizOP5LAeFecX1Ocycn6jz2YCvKtuHkbgecnWhI5XdW
PPbbxWLMp6kCFQML/dKBJLgwwBjIQ0MIHCnH8e+wNEn64N3xVkxlMVkuW9GLc++z
dWl+lmoOObY8hoLjAPfGSfVWiiSl7UJIZmb/r1BFTMhp18npDT2DxQeK/mJ4HWBf
Vz3AFFOqfdgO6jYUap7hfoxN2cFpnTQm1ECWBIcKxgm90F+zcUMdThgWJBzQ7F4z
8BMWbEcWPgs7pZ/8jqpwmgHQpbHZ5bA+lkOzoRk8gFeV/WIzaBgSip8KXY6xO32T
VB3ydVsluuOcNE1KTmj037SIZkaDiivioDSZcKPm1z400bVaw6TV+ud3SSXfHnVu
e4GJwiBytNt6S1EMG9YqwxcWC4+Chd6IwaIOjXW6II0LC08jlIuwm+0IMAVRgNhA
cpv+JMJbLLIc/TEL+0MPMJmBZpeeJN9xaY0FZkv5cpPUo6ohJ/MiVaN0JS1GsMBS
zKAKq5G0AWJizcn5XdP2v+Ad1jbIVIi4WT+NCJuPDjXflQ/FLLV7OeMQV93SiB5R
HXCd++bCSXaUK5ZIHGml9uLG6bXe1xjqUx8jE7QR99aCUrnRUQ+gjKtjniDKI/M7
nE/snOYa7M0ZMJ0wNS2Ld1dz2Wl54OMLrvmUOZgkSDCS3KHgpp04kzm0cFmTKvmj
z/qNX3CA7quyYz0R2ExbfDjN5Ou4HRVB6r0wf0MBh1jYUCvJgRd6/REexysd2L+I
jArpy+XMELj7VX1LoHmXZUjcx46i5+Jp4wnFi1xFcmOhrr2quATyURONziG5xSM/
EjKirP82rbYOWfQChfehldCawybbpP+oRMvYbU8V5zUE/vdrwvons0gDcrzpJVGi
GklraNXvi2iFOy1QAb0YxcX+xRTPUm3AqhLq02V/ThTNCNYA77Yvt2Ko8e85mtE2
F7G+ab+Yd6J32bUERlcQqOhali/xINc8MJJnN5po5LGJPw+Kkk1QgiZ73UF9X/gS
M2/col3kwvaTLOTxi4fkL69kLiVGLTVx/259d8cCA9Df6ziG0xhSnrxijYaCclyz
zZyAqf87EY6N+IopSvo+7f2PTwflu/IsADgkeq58riLWFdshNimNKZ+y9zIKWQ38
KwWi037D+CSNPDgsv1DF9QrOZeS3/0P6jvXYolFyQZscrAJZNJgO7N7JJakseW8V
EhGwlabZdcwPdlikc6d0kwwFeEMaC3XpSWE5ZrbsWX8u7CvVMMc+aTswSlGGtBI6
TDrqyI8n/5Q0gTG2xSNg8K7w2r5wfBHVVYh8TYpqdbDA9axynFz2D2pZegDRPRi/
ElHq5IuqDFsNpaRw5h34aFPCYgHWhudDepVLQCPsSkMoQqJCx7go6SLlkb6b7FyH
BvsVdAtUP258TAfss4Ed0MFBCcLzJgb+L+1brwd5mkpGkzbA/WbqBm2a8EQ+bUG7
BETzRXBDl0AwiAvcAzBbVFBXDvecoL5LC7Sjtp0ylqYX57K4kTZQ8hMx9LVuh5Lh
jmyZSsHu0E7zNhT7bc4XhJmrv4dWEqNZdznmZ5w81fFWdk+ivqSEIpsQD+DkltrU
Dh9wYn8Puok7oIdCxqF6DuwJruf0uIoTkaU+kjqTwsR3NfTVQIIQ6xkCCrHEy3xF
X++KA7C7rICTdn1bmPDeSZLRivYyN+w9Uu8PMyE0lotmVxOccTMMAgkbRH9uV6gc
QZmbhuN1rRaZ/rY3UdqD22LhBCkROeQy4T6g40rVKT4y3vKzxrtLJ2xcsbvyGm6a
BQxEEc2sCPj0Q1HoyWd5ZJOShhpJJiYIgOt8yav/BkmOZovG3dmql9JQDDKqyKfl
xwX5Y3syH8653+LGjYxBdi1DCF4x3ojioBwmkzczP0w0ih5Tlsm9rTgDH+O4BUJI
X8jmmaj3IYUE3UsfnkJRWeCBshkQkD3bpcFZl82kWAg7m+RVrgnf1/unOhDRT0hf
hTi3j2hIDljCi9blMxeM+fj0KzkdnuoMDgCY7l449kmDeb4aESXVwH4ziOzSs621
c7cAOAGkUgU+IXNlya8ugM+mwGzo3wV6g0bbBM1eIemvk1WuJ9nlRSQ39emV/mdU
GlotkxJYc7rkmA4ne1diMGFP0+gAarL4MZuVe927HUOMpTH4CEAg+jbYmvv8aqd3
grN5ujB1kmH/L/bafn77d1BZ4C7de8ynC4wDQuHnqts160tuOycoSO/JTX4Xf4rm
ZSe9tDaKMWrVvysuJmKKBr04JtOGBvsEO+CDj5Y9aVwRzawN3ReDKayUcCKavDht
uvF1yMqM86oKBlvf9tlPbxBCbuhZIMnlf2pNIi38Ksh5qHZIeA/9FMkMzoHA1Pvy
liFfQZj8EbPKRCG6DoqZvSHDpLKkXwxDeb+mDJ8H5Sz+iht3l5W47fYcdTn+Wyn2
8o/E0eZvjdwKPdGoXgmpnk5e5VR9PKHvDSC+jyiiqDgBCzQwnBQcyhLwK/CmmzGp
qJYXLH5i8PTCcfJPbe30TXaTuHX7DnN81CoAAPcMTw0nhVpOJS63+ZOZ+yQmgsY6
hTBTj5Kcx75PRYzkrjAXM6IS99H4UoHkS05kT29Tz+4lbhekh5R+Q24yq6B3TzDO
d87brDLZUwGVcsAcZdJsThQh2lDxK4yVb7kdjM2DBVo6aEWXEnNpxPtMuiZ9gqfy
42KB36AF8bve/RQxbF237y//ygBPx+8q1VsxIBe0jr8pGuf9FbUr++nZA2e7Ksi2
8fLRnj2+dHMOurgL9u8eLDzmZx7vvg7B2TAjuOjuAiX0T242j/yBdU5ZCevytIWN
H5WkWDYA5yKXI3eZG/O/kwrdCBluE+kmdOEPKIAKYcexEddb3QQZqWc24BT4uILe
LOEM9rKEwqXCeaQLCHEDYK03O0AX6hvgbjgzj6V25XCZ8ueqY8WLm8LE7/nOjBrI
TYEEZxMGFZIExLQFtBUTZpkrAgZqOwy4x8TnFSz7tDubw12OVa0GacuDVOuM5fwv
MYa3dHzFWLLMi8POOMs7T1mLm4+d3Ow3d0EHk13k/hfFDhBlbWU+zkujLjTxzOi1
WZLS2zw4Yfwuo2JTrjzmY8Ti/femOowzSyX17ZfQiESfGSMe7YNK1XCKwvZMdG4Y
Ie2jotp0GKXa2/EU2XkC2+NTeW2u+vHWaoQzy9F5zykOUWJWV1TgKznuZfv+mcWX
7DvDaoRNrdCKyaonK5dl3N5VlIV5x4EtaSmqqADsFgLFtW2rwnHZM72qlCfGtO7J
IhytUjA1SIW53u3grPQZUqXv524Si740LV/QVvFdso+EzYpRgvUATt0H9C8QiK7t
Y55nenVBOK+Qfp/veG7uAg4Y4ekxmcsL7q47odbArBwPoVkmfip9Q0uv5LGVQvI/
jvo4DAx2+WYmQ1ApC3QYpTnydUf+oU+MlyBfv4TlaGsH2tTVCPmmvY7YqZIUgxmY
+5BL+pFXR6xFKCYU1OJ8ZtkPEqdFZz1fHj9rzak2mprdTE3tq0rMhOv6JZ4r0D6W
XaAuNpmFVpi6e8J1MxuPXysibxtVjqwSA4TDwNvXbH5L6mYM8C/mQfvdMHg6ZaTr
KBq80R727Fcxfbu17Oh4RJhVbge2UwKzG3JGdSy9Hrl10tM/yXgk3+LApkYX8P9G
H9rVGY7OPE2Zm8MmsxSybhpyytdyxaQrVzvnVH/8o5N0eXQkeqZqK5nR2XfjUqDF
+WIeAQ0cbgbmYUcVcrKWdTMSORwFzTRjsr77AwBDrQmTHLYdK8aTbf+5snG9QRMX
7HqGlVmSakbpccbsHGiCRkWgfLRnVDldwzENvpS5MfZAjuX524KtuB6shXZSf8B5
pMnIvewIIZwIYFIj3XKMyOSoXaJTvfNS1k/PHlnCPCFkPTEaw5eTIjNyG/K0SEyt
kNEZQPMNSDYH+2Rqcux96ETwz5WlWlCg8QKcgDt9plWAIFc9FKABn/zDqicUJ1yQ
cdJf+zgnSbfnA7VRs1gmAmIoIpitTAp3IpYTw/f4JPiRcNWJ6d8VaPL/zevLwDPc
MtbLNHisC/AnubJTWmJSIPY57sG7TWYxlTXwaqRTDH8ptiae6CIG2bvC78/iNEqb
1skBxS7736nC/1LtY7r//3wS0uPTvVtHGGwGZr3mB0QL6c+iKTVZgN7gMOv/rZMc
mTG6j/wKGCe6MBN/HYLDEhcm+DtYc8UivSQwFi6vplwG2TvpbT2/W+T4DQU6p7PS
Ybi2P65vHCshUbStJyMafJBNUhAj5o9gJ8YROUcKUjO2HOw4W6sf9ynXcHKot3Cc
aoPROy9NNa4gIDCy1lfmgtsjEuYuOIuLIk+REoqFX+dp7J0YIiiBoTE5gBbESZSB
ORo7gHPKnsvhAGsroFo5Dgu7iKF1eWV8B4FC68u01uqJ+aFr56ySgjm+Az+WIOxa
R/vSLUThHqq43dgjN58YaqOZ2XT/e3da0akel84AFQnqF3nJTFj6cRXwczxW4iMf
SX3jVvcNA4HvVn18WmgH6Q1G6RPJNgB8tUbS00/9/XBBxbCjqT8IE57nurJUGBd3
NDAFU19CmstFbqFgfdJnnDN1Z6itGbp2H3KKz8AmOX51A92iBCTPgUQ5gnRpEydk
qJAOd4wfZPQ6uL1FV54egB7ObwiWmAQpqHScdKUzprDFTgJq9dYnfZDoUrK4K5CR
7W6iWQj6dj2/bJWRqgAZbOoVwkNudO7BYBM6upxktSxNf5QQ1Bc4j1VlimykjKgD
8higay6GmySUnKz85W04nsaIf0TeFqGA8cGVvc+Jwe5M+DrR82Kkh1pogvTu4/5s
k/vmIwr6xhPm8hifMvTghKoQCXthZWbs0TjMT2CfDHb2J/Qp51LT2Kwgldjfgqtj
c7QaLy5dF21TseUBhs/oSCEcYMbQ7jFAri9jZPdX/LP1hn3juS3iDBN8+wV+dInr
t5vKeYVJ9YbPM04xIiJyYwO8Ec/eKs2x4gcFdhlaNG/8tHc6mRJPDtRPu03TKdyJ
YOIyG+GrxwLNwSL7e1s7dAmnR4/oD3ecPLF/liXyvqzfkEIbXpMFcVL4SuxJty+S
msEOmVRg6RuXKDzQy3ROeQlTvtZCOJTyWmU+aumRq7LwKlM1Bfl3ux6ew3PfbEzq
C0aRue0esXMI09KrYsQ1SMz9MQjFYqxjGXpoF3M5aINaImh1sF3glJc04dE7+ZIM
2iLVbtRODnalMatDdSkwAPf0/G2sOowljU4dHlo4KF1hV9zhWW1Yzuzml3oljU/G
/ulbq/ASXXJgWFKiiMP6gazinctK1gQkjhYCAL50uQUF+rvJjmeNJKrrn1WLvpOK
mnAixizM4YFK5er5YeG6tJb+cnVl5azIAGmlANQxvbtg4Z3dUiOLG7pVisC+eUOB
FS13uWg76hpyK5jXYQSwX7aJmKO3t7MZPLyzrkH+LerbiOCPyrXCx2IVUqRRhIjx
E+/XabNLH5yhLfsKsw6vO6Q0rmjcvoYtKGlp7anZtF2XbynDWxSSykPwHYrZbxc8
L270f4S/WoQzTLYF1qPMvHY8NcQQMGAe7vThwyoud8qRhYTH8GrUa4hh6w0mKajf
/dAJr455b5xe9xj77TYTyZLStQH3Cb7xllBcWISi+fkJsx4Wcrzb+holToYEOg5z
I95dkWnDPDQZxb0V/oL7wMBzoMiPdkuvNfP6zhJsIlvQXGvuk9aRYNGMqfyawlbu
+NgYf+FJhGsuXWKQ5crLEZeMzGKE9oXt/0bdrQ/7IsmGsYnuAsTEzUQteK1KvJNf
MhmP2LBBI+eijG80gw1MWWdDfEczcDrkdnKgt2B0cOPwLP7DQqmpDi9zjBfzoSrc
LQ0+9zUEXC9vWtDDOKaX4ScquQFP5pZ2/jZOYb22fgvVU4e2MJsLoaARk5NrijF3
JGDjkj0NSHJKZUzFPVhOmU/lP+DAoBI4gvwNeA6x084MmXh/0/lpVoTRnPblo3/W
xS9D84F5wTJjra+fSrreTM+efkPeAxxRurPZIXTPBfAkUuPKoIUjXn+Xyuf7MtEK
Zkw3IaDznVvkg/qxKEfe3+e7RHbnXbLnvrLXMfN/J8sT7qkNAlVu6jWe6NpX+vUP
EfK9nZk0xcvhl3EzZe+k5cJNgKSwAZYVjfc7tpL4daUNJqOtYNtdyMJlFmHzKRsG
rpq2ZX8eXvocX0yRwpLXphCXxTbf8tfiiLreKr1Yoi8u9UniacccMJ00HrOrxhkx
vfO/oFkT4k1Y2mGzVjbE21mISQ/RLgsFzYnV5KmvsxMmmzr0mdSJil/g8MT1XZxm
cFdiv3+3pcSsQgcq7KFdOePymZY0zYaKl3zDdXTf9be72RbV6QQn3hV6KjwIoNGW
HqgQZb1eQwKZnTZZNqtUuchTm7wfBv4lqp3qsDVx2gEqJpGwKjt2HRAfHVuNRwuI
xEQnDtpY78upD77bVVpGdqdkntjc8BeXz7cB5IuD1zEBFcsXrh1qL/fcUBe9orEE
cZkjg98dOcSWvduq2vObi7WJFW4hfb6gG+YlDf67VN/gyZu4GMXAQZUOGxQMcPqd
rmi+SubG7jVkYzH3DobPaj2Vtdi2bPNXYVmzCC4MMIGQKCmWMLmTxW9PUSZ9yCqT
xb2k3uK+xc70Al48sDJddN3A9BpImL/q891AKfRnM2YYc9jZ9R2UTdlLs1SfSekH
eelFF8pBk8Dhzb8Egsukufm/qGMLSMPSkiZ118AsGr6HWbKlqDDEpCOTkUEhPV7J
jsFYXt3ogS/DqFBG4S7tATUhlRYhQms2PTucIXH6GRCR9h/0a64A5LZgfLfHcfnJ
jBXGygj7OmWUa4pilYb9T2E0piU3kjs+i/x9FcSVOnAIa7ZlB+KelhLS3nBBJ3sv
3oYH9zL8sSSItQBXSpsmrDMa3CfbDYpFQViH8MQkSkn2ZA6zb7o0knQkynNlUjPt
HWRXxL7mCvZMtf7YR98CJsx2CgWe0JmIngrrDLB7CfGD/MgWb08zoqWREjX2F6ES
FQWfuPV4JwcTlomI0XrmCrtQ4lXqYjR8vt9NvWcb5nIkYiV4Wyr9RqoDwyJNMHos
Bs1Y64Tz+EzU7AtoN7R57UR6XXa0eAtFM52K/3fvM13zKIF+PcykRhb74DItGpXR
TVMU5/GIClsR0K7firqR+6DNhRjRSuoKVc1ZQinwxHuda0q8JvcUgnyUWBzl/shv
gnTpec6zE1/pmW9kVcGN/xUhNu41H1dMIflfS+dnkJWHHzf9emFWVSQPdsZFUpmD
Ec71Zibgu1TP+eRaKc2tBdSqTFjIq+rR6qNHMaKEVKmjjc8tq7WzSAjarnaU+CJK
WTd37kLyRmZRbRGvEipsVKFS4qSnP/O8AE+2FyIC5VsHJd7gNr9PJsrLi7/h625r
85K0qjasL5LQ2U1nO9OI4vFyhrVzTr5lMBoXXDj3AHLFxLnerREiXerNA2L9bghN
juJZc4GhjLtXkNJqN3leHq7TilPo/75UXC8GWsGOXuFj7RWPKvm6Sj0z0SY3XdUT
Gv4qUih9eLS1zarvSKXMJLGjTGSHFKWQbcF0Yj0MG7cIreI8OBAK+a6yCLoTDNBY
zDbil9p5durCeYelu9mUfzbT+XMlPviklLo0DOtdHkNtknQgNe0y45UCsSa4cgn7
Jpk3S3Zy1J4PDC/tybmGU8zAYw8WU0/ncS2fCWo3gzst8MP+tQRPTRtVHWK6iKbe
PWpInzKl15BGUXf35qaQc9A/FoeCjQBla7CrFiXL65yj7MocYFLGWwljhfLLcKTA
fIsgvEBJHd144I6FSufpkcxAl9zj0fM/NTfYgiR+6VxO4z5f0BSKNb2XdwP5ViEC
uppZQTv2p63D4n+2bfGNyshGXq5BI6e4o+k+bK8eYFLwLF1pjMokxsK1tfaqxeEo
TYmfYKCmV1fG0rNmh1u2e3ZJFQ89HciihJc0KQpxrDbdGRhkUpIHDGnZr6EECSHy
1lwML0ChQG4k/eNNvZIxCCm5YZ8aBqFLnTnXD+mwK6b92vceytqaE+Ybh3w9AsYz
vyyq4qwl9g8QOW22e1PZsXvjC+VC1sUgkmAaQ9FdLeQ2Im21RLL9VliNO8XXx8Iw
/FNYSJnlIUcdKPhiX6moiHfEzpHgsoQ40EsEkfJ2xqAdFkAO1rShnYHFyA++9Htr
bIPMHs9+3yrHaUO2Sp6AsbC1vD74uMNQ3sRnLlKjXEIrS65v/DJbcu1zIC+WCzqB
JuacrXmLPxR1yISkKqDgt20XtYlGJmMgkT2fElHDxoMrnlpMp2jIRDbhXJ75wvPH
96JLADF0wPm99mLAlUHf7/T0/geUUVbeL6XmXjeR6Cx+Cu1b2Yfo0CWmdRAFgCdu
V74kHktzUJetROEAP+9iIHi7jo8mEp8LQi5p45aQ6pTcq/2kZ26O+iuObRuCpHll
UIr2ku0bGs4sTggCd3cZ0ELS4hYCoEvAiKA+vxb3b2KCOm+/9c7Xr4GOUbXGUnFE
wf+1DF8l6kZa6v29cFVmMy7J8Rz0KdSC+G4LAKIx8akjjJgSmcVnhZk5fFECqtIf
kh1cg9I/pQC1TCRXdtcfsKAMbB6PJWe/sVxWXupKRyq79H0D2Hxyq4WAqD+5mSwV
5d6yM1q858bcfMaubuD03eoN8j7SobcHtrwvIVa5PthU/KzT4uxlN3+VKfKkkqSJ
G+pYLU5ipT/dAeC3OoYVfpHfWLq3aYA2kA1rAC6uToJAu2Fn2c16mdWFzkYBuhD3
LcXyy9+qg8SNLq7dW/po7zGE/WanhgaZ9DpQ1VVfLNV1I1tAKxKUwiCx1ppkWm0U
kdhr4S+jv84VERBY46EXGhpHTN6qOi0ejZmmgaNnB0yIm7m+oQ/f90qYm1X/1RyI
1/s2M4qUpXPT8evbrphwEEwY75GH+5Xh7EtFQtgrhe2SrLaKusQplTrTAps8Mks1
xwfXQWEOwwO3D+oCzWDQcwwh0cmxCvubWUrYRuQ5fE0SwXeCHmomhfFAK65sFv4T
/j1oRpHoLGCMEmkpaoXkNk2HKDLqvga6BwJ6iPEvh9UqBld9zPY/OQWVLIryjygP
sOe2dXu5vZ2Z6sPbYizp6z1s2BIi5G/0ltpLXqZMBjpZ08Xj4pUxME7MUIZ2VP7s
N0ziIdVAX8V3qi3srN1A+TI7zZxLG0tezVqTkUqRSLsUwUf0oQwxpVUinne7k6YZ
zPwchYx9Ire4/tNK4zgTiFLZxZZgUw7dXKComvfnb+FbnylNBGvkSvZT9vT2Ukw3
dug9WC3omCnZ+Ox4sSc4BoEoZl/2/yQ/ffTYOO/0hnKjYGwoRuNTBvwP01IFrI2Z
8ryKdFQpD3TY3yPzPuHDDo8JR02tlIbCew5soZl1abPAgfASAGBfdFg2Hs/m+fWb
TaBVeki1zbZ/9R01+Im8JGZdKxoLiaRp73JyRrE3lmaTq05mUWRgkmG6GcYCtxQn
DfAOmrKY1DLAl8xWVuCd5kwh6ncigUqlCbOvtGSvqSzJzlG+B9cIatyTeWpY9FOJ
SKekbTHqHrN/HC3lmug9+xPkhcScyLXKQVIex1+Q3KqHrFnOGDFxMACNaXr+VhYM
4+HpHS3B61GL0/6UPbiN/b9X9H8/yM68E8yDeY6bFfnOQe/4nNeK+uTxrULGV3xM
63aasCZcbd2s4qrp2W0scDiDpNxZW21Lpe5DKrlhlvVzTZxbTHUBKWTEqU0VodLM
hlkVHqvivytPbK98ln19owzBqTnbmwHjWqnjJBKpJuv8rchdhZdmYxmC31ByFfCy
NCVF4UAxgI0zlfnfwnYnwad3rNFqGSMwr56OqNw5n4covA44aqWREKFMvyTKlxam
vBjTtg5ezWq/K1UWgO2d+4yTAahaeX6CQD7kzVKJ9XbS4wyfZtknEoRXV5RStVhX
1yVN4+I+RteHX6CJXRqhP8MGn4rSg6fBEc/CBaX/zzCP+bbON6QZCDo0WkNIr5hE
enGCrhi166S6GHSRKh4w3flWirfgTeNZiYIktTr+F97V5fKl5xmmWhWrCy+zGnOe
xdplAdlmRFbX95HW+VvhloI4VRC+vQtljkEabyMYC6mg0yEza/TdHZYQFhY5Zjq9
F5/NiFVzY48YzO8HnP9mSZqxbRHgEU+mxK0SrogpOKMfkFkNoy610p7J7MZ9kjRE
q/8HQPPZMBAyir408q4PP9x0mZwicFgG6nbglrTXFQodezg3mcsslZiyoNXQsydO
KmK9ytkAfzf2/GP94tS8NWKY6Cur6np1NOGcx67Vv0n6Sa3ouPf0mni6XiVITPDQ
1jPiiO9vyADrTDusjVTIpQRYo0F9yGSMMhVkTxpB5muCITAbPgLXf0dQSvaWMnkn
6P12SIwegZ9ElMQGPuoBGlxj4Y6XsBJiTP1erQnGWg0Tj5OvX1k1y6eC6sZ2i0Gw
ZNDzooCtL8h10XcyrlIfyof6TACW4w+D5VmfPHQWFviukJpryJfhCk8/pefnbqG+
CzRmMn/wBFE0dEqhK0lQIKFoWcSWCS1iD6429B6C14D8qO6z7WYNNYFqouRDD0vE
5GgyeUPlNNWJtO0G3ePu7xj8HEOVKJLSQRrseiL5pXVrzmQugD3xi3q4FhF8ZUVT
0KYZoUawr1oaF8ytZrPPB7a+9VfwxQX3UX92jKKUjsHW+8OyhdPme0RH3dPDolye
AVasVx9RcfQSdTWlJTMW6NAkjiAQS27mjQWck2ezr92g+XYMDqGumT3bz+q5/nWi
GXkEzxraF6oAq3xf1QBrzNj2DdduND5c+D9zxf57w9sJxFsiY9zGPfbIA8mN/9st
laBDi6N8e3w+p76JVJBeb+QriIBHURL4qUuyWcCJliVpanVCkegr96oV1416xM9H
VczvKL3049RYbdv7Kq5n4kNjRiAraGJZi3Y3LkjG4bh/AmWV8Wy2mQLsa7r/mzqW
y6dmvU+Dj6aQrjSIgHxlyzzVK4s4MNm60BEboK84kTK/Gd31wNApr5QjdUaBSuTS
XQWNsQxlr17MqUNjIsP3MLQtcEcUNstmtIlgpJ5shGIC4g/zmsmfjX9A4NUTJ+5P
I79Pfslf/D64VPf3r/4faOjl0CsweDu0MBh8HHmmFgK2VsgMGZ4ybHXs/B5MjtJt
zBP2gJOVdpHdJQqy6ZVLj6cJkOuQXeGpZI9T0aZ7IypnFQX/nm+2XATMIevKQlCz
AohJOqqE21NeWWmcZbhkiRLTn6unHTm40suVZd/Diznj8HQHQw+RcBriCFd8KeSc
r3dz/RSuBFNyTk+rJfrXHqk1rWlxm1nrja84QPLZi/Aw2HtrCkuhJIc7uUvmNrUz
HI0sVZTa2woC8JGVXtyMsomPvM5e96SWB37qQXSgDJNZCU9qUfGq50E+ADchPmtU
9J+X+DzAA4e/JgYz6D4POsaTTnup67TwqnnuJbZFlvz5tK4Bsn1MWjhDnCiEVifx
WkbbAdkaV5Eo1b8r/yAxWqaVRvcQLUsmIzvjpLFaTxU++jmVcHwpqCYGt2zRvftn
SncW4hDB30n+49V96GYjBkm597byX2Eji5JN9Ro+YRVWpXqceNojZAtFvzRHfjmj
hecAYcqXNYeV4Mau9EvLWrQiuybD9EDSayVOJCd3yC3f8UQtngsQA7NMS09IdKbU
gOFROFxnzMuYY/mL4gHY548Z5bbY+TohtX2AhshSy9zn1sQbjrzjan++dfgWyQ/R
YQh/S/5RE46VDGZXKqPqX4GN4iMn6wpE7QDI0+7IAQJfG856ZoroZrYkktDnQDXp
J2PCD99MZljXYuge+bAZIL7tIY0vTBMTAuNQUVMFBfgvxvGeEWNqVPoWTcaBbTld
JYKZ8nn8t3xXpx5brRi/nHiwnNIdctwrdGGcg8+D1TTDaQINp/FAygMAvVC5wIxG
gOTXznkNfwOCSgppYDZAQKBcszhK020dMfj/5QaTEp0dnWcx0ncUB0F+4Jn0t0xR
SH6qSOSm9aKShDKrvLSnnWAyKhABx81mzvL1pHqy+36iii/kiH9WXseL7S7zOJvv
6ClJTg0Ihi6+dug7732gdEB2AqBlKNgZ5/LN/qM4KK+4pW8xN5y4t6QfTtWDLCfF
JKg4pVuoTPCFWs+YYEhzVvZj6mLd6pQvoBEf5QyDAb+g9BYrJYFivIw/tyzw2a8Y
bFFoW8KufoBMXY+m+ScExOoG3MuiwijUywghrMllqOSRiGFP/ak0+EMDjOF1J+J5
64prOKkIDsAjwPpzzD8smhiqiXTJXeex5DwPcFdb98tvg3VFw3Lyxjoyb7WpLOTP
e+jkh26DOsGnOYkWIJZ8+XPJhcnPKZhe+BBikkWALexDei+ASDSjHK3n4VEm00IN
OPEjUWG4DC7KNx2MEAy7FDnCXcaPUB3/crIVlx7TwQHq1QmowRNhs0z1CiRVoOXZ
1ujLrOxAuKk8TgVK41pxGtnwJsJOIutwk2dvzz4sgTHqPPNciNZaET8/yOUntExm
j6gEH3ugAZMiQqvrY9oqs6p/NQffl2RELfqJSaNIaLm6eHhD8iXGuFCt9shC/dej
8jP/rl8Nbbg2VKyRmVhcWjDIWHTMNYUEPSVYP6rVD9aRmDZ+dzmXqBn/Hag1IcW/
IhF9d3Z71yucUzFB7lGbPUyG7lRG7s/oEdj5s1i/+QTtU/5k+jIICSNBlStK7o5H
1xdLCnb8tVzR44fpmyqZtVzcmCMBgeFuuT2Xx32tToDDm7DI9ohoRkFNo/zHAqH0
64Fu1M3JsDWoMjT3MCVR3QrJSpp3FEDO+aFWs7D1aDFBjMG0bxafIK+CavbhA5/g
txqCiq0FG4dKvAmKavMsWt3PgUoFWF0VGEfrGNV9+6OfOTxeg89h31M7X849qAg/
ab1zXxXu+KWUzYBtY1hydPNCN9FLw+hycmN7nONcC6UZK9ycmj5Gfx2QQj6GvE+u
Nti73E6r8caBF2/06YpP2UjsKYDBeHHt2xdwYDT90WbJxsRyXYPANJ1vlMFztsGk
Sw0UtwaUxSwgpIRVN86LT2zDI/K0Vu1Ed/GeeRIGg0GolThX5EVcClT4ua3mUyco
JYjoFTN8h/e3iKPFLhk6KOntvTqGZei29yG94thodKmEPkdu1N7VpbKynwzt71sM
c5dnDBT8nvlHDw8rs+b9tbrL+0y/2k4p/0NEfRjb9JuJ405MtFwsJBBLAfkKuLu7
5tQpTHrCnvcb7Aayyo+eOgAWrKljujju55X2HAukxishDNM4uWmSGjN/n7XgnSwY
HdKzQmGyCLpyZsvIxBaygpOtSnUejkef+lRQ1DRxlYgDzpbqShP2pG6bjc6kdUVF
FfGFEGNuYxCdEQ4ubzhbqIcfAzmX2cwnBOTs3xIAK/o2VovboyPWRql9E8dsJLwQ
IvXRPephELksVGsviRE9IEC7o/6CXbUxQ3thJw4neX7Nh6thf0Ndb6F4Pc9U/AGN
aeJoMW1d/MNRlKAJIGFpND9m69n58DnHm6Kxg4qzU4y7PbZRLnBA+Ji9fkAhoWa7
VqB1LSZfQXQdCs6Kr7EU58Y51cAgMyP3UQyUORCZ4NpvN+CCYtguNetBLBCJoFhr
K/sudh6HmoN66veleaEMTW73mKAsUHLoKIe8qtSeRzSEBIEKXTXAgu/bG6rhAFPl
4e11PiJO4JUdrMnkby1xKEHRUI57N4Rel3XupSRctZkb7IS1Cvde8Ra0dVtIacks
7kwZ0KQbFthaM1KYLPXpVmLFG9wnDsZeJG/N9uc/GKUu6CvuoN5Sc7u7rvZs99mo
8Gbb1WRidBOrJbp416ju4KR7xAM8AdkETXFtB9CGFV2Mu4cY9v33ePXwhZCHoHAB
ruqoL/NV4f76KozjCUeso4r8KNY35XejtgUKUADz748g9FUbKt2xynJPuper87Mz
3QcZ4dSogvji3kbjmgXt032O4vzfLMNsAxwSBQnbYDJSWFXC+63O3A1keoRP/lYh
pD1Tv5YuR1oHK+6MwosMSmF9ON2Gfi3TcINUEhSIlJr96um0a93ieEXR48qMGBm6
fJEF22TmoqXGrF6WtESLwPkSv8V6pMGWnEZuZvHTd3nWWp3DDy9y12GIWYtiUL4K
o1EXpRDb6KQ0eyoLOJvxm7IWPkIIZvOX3bycF9DrnbUZntO82X+5zew+dE+Za8lR
c6gnR1cs1p3oBnU58ZKDBbqJi5TVmRWA047HTdg1fESnJrJwNABqlDgja98v9mos
eUNwCxImCNgPelYx3+jTPQ+ugitZYHuGi6H3cf5/y2I+ZE6B+pUmvGpyIu/BVYxN
esPuCxUvQlHD7hfcO/6SCYQL61feFMzcwMa+jM306L8hG735vJfkd6Sn226Tqh4j
IEINf6bKYCT2i3L64TAkGm9WwVr+TzgfNUay9Rrxn8/TUDrc+OlPMKGdgx4SM63q
RUUqvdHbRlyOblN4S4KuuRQjPss2IE0mLpkiaREiL3cRF6oS0K+KHI0o960scKYc
yJRPfheoj8z5+iryAtZnAQexFZ2oF8p4ohiGBbn4tC8vnW5nTIgyd8/UENHCCeyD
d5zi+vp1mPjbSviqfUwk3oNgQ5iRtnFdPdqx14DVazv9FHh6UUmysqhMuTJxkj7y
hXZkEdho0VMvS25ycXCtwG8boRKFSMOj43hzDowIyYBrZpwiPOGCOXq4RSMU4OOc
c9SxrnqoKek1mBIXMVbJFtcNLmGudkajQfXxdcRpFRfT83eCtT0uwbJb6QkenwrM
Y+3x078JzBhI3bypZYqpncTzQSmhDwjXdront00yAkb3/0XWRy/XbTBxDgxkl9op
U9n7sAauWbyktliV0opCQ4D//dPiSoetIwxpAEQCAV+GcUqEy9lDT0dUdJ+FJxHn
vPscm9CbGIeoRd0ND3n1lpmr2idtO+sSZQEVCSkQPdPRy0m3R1U9YeGz0c01FArW
29BTtUZ2Z4Nq+SISYxpttcJOzs15eNAnhPRU92xlwdj91qXY4+Uk2MTRNnGIpdjQ
RK5ynRGPsQrb/FfM4FXXhQ1We+X5u6jTWT7OXy3pFQHNWPs03BK3vmPIxuTmaPZc
u2lfdjt2LL3BD8Xa4JZdw5Bc3U3SMp7U3AGc9EGDFWHoZVYON6g+meWoeo5Ovjrs
oc9oZHeK7CYUKJa3fjPJZpg8ILZR3c7obYqiA1ic/lTbZUu4qpfq9kFQ1CopCbnd
60UnTd7N+d+KZ3b5nKlYWgezJ7DICYwreLib7qmLWTIQHxvBBRMIZBmbLgcqueRZ
r7o7u41qY2SUz17Yx5glSB+3LBxg+r8NtWrXYUDYSjcf2GEDdbEyxl2QKjZ8WCs8
kXGXiTWy2DAbpQCi3p5P0vnH/2pFLoXlE1cO0F+YV9Kn8MLS0OdWGNznpxipURir
TwVoTTrCBeUJdFssOY2wZOk/Zyuiz25dwmPx5H5o2okFsAoGqa4KpzG/XttEMFUJ
Xu2fDiJHtiSdu5NtZMwvCcheeumYXfl8OXQvTL4kRgQ8CdYS5VBT3NPUgo4P9JY0
fZR4xc6l9sisiu74IadXsYqu9QkQucC9qYnLRZm1sZgnR5lG0SNyhWyOpNNcW9Cx
3Qct7ppbXv1kaTj6KKqEM8FcXiJy11GxQKgfR5lAxG710SzRrx93GfyBNJC/kw+A
tLbetactCwuBz1h/xBT7xN52L7JK3keO1F7lw5sRYX5KfZUhMLER0erK9Os1boLf
FG1Ll2ngH3CqHxmAanS1WssvJuGgsYO3iYgOfOeXYh7fNZaPoGyMTe8VkssiyR1p
BtAlFfHfnFCCOLoNnb+OYhM3CsJDMaFNxcGHSEzI+d14MbSV+3WyWQFIcH/LTL6H
RetTwPP/mGMh0ftI7cqZp4XVEwyiZhhAgqWPCSPecmnbJYIN3CAiwMFc4TIsH+Xo
5DNQfF+haGovuL6CO4OzFEYxSKWa3H6dxg7l/XkJH9l/UkIeNwx7OQMDctFGYYFY
X1MLYYsZlF6djUM/I920rFQUtMOWn2N9p864KqSA9ihIhwrO4o1bZ8XKPVfhec23
lIChfgBjdPbbMN17TTNNNrSyzfCAODpRca12gV0Y9WTTV6ENxG5pJUMDrIlyE/Ic
OkJqVRmDdTo74o3ClIBGl6Ote4OKsZ6GljtwQkdsXA01t0EfxCPln6MLCdxHfU7z
LxW93+0j72ch+8DNmlQb1wYJBZ5UD6yaL4ae2WGs88HdZmwGM05y8g4xBWWO3RSR
HU0nOosHQ6B1TIe6niH6tqfSQrViLdwgD176Stt7vwURABAyZ7O+GO0dxARdAraN
ODlAqMHTcenXUYTxfa4HH0yaD7YpRG/XvzCoDg2RqB4JNP+CrA6uMIY9IBwxxGag
tKre4CTf64y6qMGeLlwyuTI/YYZ9h9T8Qvp4RRepsvHNKJ/T821oSCA69FLMiUg+
2bR9pofPunfG86t0mECTmTKOLVAXxB5KhSTVEr12SdIzzNgg9v8qapES3p4T+tSI
kc1TumjX2we7l28lUpdHAJJZkbYCzuHzeQFW6Po0Erra7EwADhQzRuZ+ZTUVsI/M
J+jihyXjC90Qn+d9dgbjTd/6GQ8Eq2UIyZ8RT+9Gdpj+unQCtcqhpmldtWS8eVVc
qIfARK5RLFKQi01rji0MPkfM2x7cxNDylCUb+myYBSMJFqU7rLOA6diOP/vYzz7U
vVsbRZHNp3b3TJNAuJiuo+3T60izR1qQOv3inks0riQKVXBja7HXYBFHfXQhdmpH
KeewyCNujM5Cmz7OJDJmNnGmnXIKOV5MvCD+Et/CBEy2XiaDOd4SXKv5EbLfGEuG
MFdTVNIaAxUaW7tuZjyp5X78Ja0ayUVFkqts3m6H5sB+hFoinaB5618CUAnoe4Ln
aI7jIYfOwgIcrwMZVZPGcc+Lp5TmEn/CwXU5vhcJ65eFBZYwsCxbREvVsX40HMYd
1Uid5Ccp8YJdNIqBGafFLtr1tLVY+fK+h8VpZklI3YgBVXZIXOaamQsbllrzuspE
cWr0r9/lThJHlldnsBHYoc0e1S/W36Pmtzf33pKhRE9ldeLuW0scEfRJNEViBtaB
If4JJuYWj3Gy/2BMM+kJyj7cN6xHL2DpkLM/Sh2kO0nnhVwr3TvM6n2OIMmNIzq0
cWf7s5zw3g8muSPGrvwH++t4FJUv5HUVwa7Puxr4tAYhi5FwyEutQxaAnkLoi9FP
sr66yRwXFinxsP3tN3gj8ZfOOF6iXMChzqBN127G/6FcWrQ3cFeBEmjFvSBTnAYG
ydQ8ugvZQWYQkQ3QUrV1YdJh15D/NvahUuLmU1csfJP4kiviNUz9hypqLXCstz2e
vmcgcAahVY1oonUpAFCvrBURc82kfsVBcu+lq8zq91NUdCV75fy/cPARyqr8Rxqr
UalJP0IJqgHyxWawToqIBtjGHO0I4f0A+674QTBT2OXctgX0eHG5SGFRX/W6PMxl
wg+enW1Fc7TT122eh2QwuhfU/av1784xQLSPk+05UZ+9hKKSzGjipTLVcXw734th
YpDAUuQ0cFd7PK5FQcDGZ/osGBZJqMlHKvRZ0dt6LH+0xozztfqF2DO011WrICGQ
GR269I29Z+c34GGkfrivGSdHbRVEOg6nNx0H0ckc8uQTPrtTfg0Sb663MpYIg/0o
LrQVvF4590szcy8eomIsLWmwg/lDQqWITLhirICkz4oJLSkFPyMya6iv0inbS1Gp
FVsy5RJNYpUeJMPreAgLbUIkZ3Fbmg9Wzp5aA0t+fO2j+ASxDWcEstyNY9B8NbGB
6SXEKx/mWM9lgeN7zQ71d9F2liTv4s1vlEHZF4CcUshpS8h0B2kaUB+3lP7LqRif
vu+ySTvxPwynYl6FKs6xqzIb+C6f/EI2Z6alrCya8In/LbxGgmOybh7NeXo5Lg5i
encPetUzX+CK7uIVOsQK8J6f5bXWn7qyLQimYpa5lkwielMpQB2nxtu2bUJeT7/N
kGpoCf/nbgB2LZtsGZ0EJB6/+Zazh7HriwPHO7EclOyjHGDVVCit2/RQmA9ZiKMT
DOWsO27NBDeiDmzpbkO6sktcQ2P2az7/k0yy1hSwGgXr5/GVszhXrfG6CHxD4ws4
QxMD70B/K0RgIiLUk2UTxuMhbv5VlrNdXq9oYnjtc+mn0tM4c19TxLFexpqveUYE
VE1C6cjrN32iyiXC1h0RRWLwJVX61EgBh5hZvx3CIlZOa3zqEkoDUCL3apMuntT0
vaUUZIeNKqvNfNhtaDZjKopGovqViMJ86fZlqK1iCltsx0mgKGNgs1edDi+o0wGf
wBw0kPtuPF5EOQtrxHCVM7b3IMyb0vfxHu7Fc/1/zI8d/ZvmDVMkanfrELZINExe
j44AvfXa4hj+y7FEvTEMBAeZSkMpK6/L2Luw5YHRSS6RA7Xb2e02a1Jf9wxPGyz3
bjrrrV/u+anXyGEu78ccYvPKuAj2x9PQYMAViIind2v1OoV0bTUp81hlgBsB4t/Y
6ootwTvCRjmP4wx+m9csR3HvmXyPhvYAnFGtP3Zt5Mdgq0NarMJkAu5qb/zZgVyz
1ei18CLrNG2FvkYWV93qVtOSc9hTCvfM3u2Yn6xXpizDPIFM+zeRE8tv6kdL4o0b
+vrLDsV3+w7yKY9r30TEUvcWmntvjrmMoeFvZUu9btZQJ8VrFO6F1Km4/KMaZPtC
ilsG2xVaffD6NJSHOegl/MFpxYvxHlOijyusWNNsegpThShiT+Kuxqil6ntgUqOB
EabNE7w48snRWGCgmeOl+47JqH4qpDkKOEhR5+GarAPR8JR6OQhrayD/Twr+1Z+9
zPp/Fws6QLdXNBDFs/QpAf3BtlrsaABYLW1w0ENQPnrVp2/P3ECZywpTDHsJMU9+
QCaMHVps1uYn1SX3BpoiCNCJtHgiQ0NdFn28RCBi29mMoFjOJ6JCzcbLQ5/DlUro
D0Db4/oylcpqRTbC3DWrN59Ow/Lcm9AuwY7JEDl8Z4PX0zeRLwMopTOyPTjO0f5u
zpGRzlvAwOyvfQzie8doCDqEsxGNmkthlOt0TvPcs06XK+cDMoFh4p/QozRNm0+I
+1PzcBha+VVqoFYk0IFkwyxFhV5cXtxiARvAyC/MeyDwn6bhGt3AUFsewDemy4kK
gw/QMfthSMtI++Ckd6rE2w5R3tGRCGjYK8XkXJFoMPjbT67FWFZCaKYg/DrmO0rt
tP+1ZyOLx6H+RdKKOBOooqAHugcQ+3Bo2D3eghK1AobUzuBV7UTkbPLPM7lJUQ6s
VVdOQ8sIEg8oPrm1VkQubJdvDYQqNzWtmygSgLKIvIajIa7UcTTHyyR5vcTr5WRY
0sOdJu/XNXzw0IB/TsTKZ607tAW5K2hDDmW3UR+WvuTU8Qhm5j0Ixo49ANJi3pmH
SxQ5y9NdSDEKj04WpNPoZcCHAK5f3rLaeZg/8Zx3ZZl9XWCCbl5X6mc1UL/u/zz5
RBAF/ztADcTT90MrELNGXBf/SIyVuFHVqmsoN/Ldx1PnDLg79SozvQS4w2QdB4bL
hTES+K3q0JTVX0b2rZmJWUtN5HDYDEaCbhbnblmBOW11WG+t4LlCqxGBDsAXQT55
BOdjSrNKO7xjjA9M6UWcjZ9t1f9eFlomh8oOTg/yRVM3Zsrs5Sf3RoR6Y6gr36Jd
cAgRvt3pvll+bkjocVTN4qzt5ZcPeruWsv4PrNXz5ar/C+vGnYXsZ/yeb2UH9+fR
hcBV4CyPAzgPJWFGTNfzGuCbiTbBcbURn5JGujKL5YABvsvMz/6crn/Jdb71Ji5s
+xrgm8Uo2kXp7GYzC8k0QsbcuvZzFWsV3aQFbZRoZN2F3F7qB029Q6GCyfVnVfUK
lOmu4kioaOVTMniVBq3sop8XAQj0E/dVqW5X8qqrwF/u1/gvZWU66MuTiB0H4rNf
cRA5QRf9x2Wm0Ai7WA0ZQ+Cw9ehOE0cpevwdp2nwSdw8fAJiWD8bHVxEHJv32YlC
gLUmTGbbqgnaUtnzRnow1wcqOc7+Uzy+lHqP82xTo6k1Prd+CcSPSI1YdRQWvB6o
qkLcdPAgQoQBtjs8yznAW6sAc8VMYUslWmlxcGSLYWi/c5iurPRHdrHqHdsDuq/t
nXRNLuVWfqpcBsCJVVWHg08PvPHt8afD2JaKTXwv4D7CkLBJ4Vj7wm8392kWgR68
YTud3I2xMFp4bnTApm1QfoKW1NJtt8Wmir7ixE4ycERU2zH6gzpGkx0LCvHAiy5R
Q24TtOvdAkMbPnDmnW7EsxIhOv6AoEGvhIWobUxLiFmDkE9qy8OpKpigNUdeiEU1
+w94NyByy1FoeGXMeTGrqe3Qin0UV8zVoL/sA+aEOzKX2fjoTp7nwMWDK7Sm5+sg
TM5+huhSBM8Qf+sRaW/+gvofr4AguVZ5laV7zt6cAHiQatl4xUqZQHT8bUjrldqZ
9UeIvsHPwBjCewi+q+70aycpza1UiJ9VKmwFuuvPUXMvJ/2EdetYpdk5Td6Z2oRG
XU1VCt90acaY4huZ5zS+l01S2PlfwI3iaO2M7yrH1s1AW9MiDShMio0BU/f0WeqW
hWXMAwoNlLfIHhbPAgLcM1Orm/4RGTp96d1TCcMlaBq9QpNpcxjL7/6wp40+slhM
Wpk3z/1b0/aagK7yrPhjIZMmxFFC8n9J6CUeLfhA24ZWeFb+ULtWcaFWTd7Cix6k
zJh3PHUy3kwafGQl041pFgXHDjm7vRD2L+uYvacl7U9zaA1vM0ZLUmBrSZabt3VS
J2VEGVvLQkCIX+NCc4nKYQzJS6oUps30k0PZJB42ZXZ+0jyitQmovM6PZcIUiwK3
eeTBOTqIc+G2NEZbgxpxkRpSX4yw2GwSEZZ5m8y/DkX+huXsAkS0UOoJ9gWldY6o
pGQlSfJfsO1UrTrnJXR2sWi8sw3PCGXKvn5Tw7qXuJeBbB1fYXv9D8UXI/806IJ0
6f0PdPuswHkhtknmqrM33keKVmjCFORAScdg3d7bj9V4yoIT6ipQUAqs9t2JeMvR
sUo3fnEc3GsBI93Hhq9YYIEvMaF+8trXEm5aWIed+jp9lcs4hzNs2lF4NvqGU76Y
5wqKkM/rGK2s6s8FaoYDESlu2qK/sz67rE/LRz+Xw1XMq+EMqWP9VwCF7jHCVeA2
m11vdjx33Jjj9Tp1jZt4ded6vMMH0Y3NYnvHe/F8vkM2H1rL7Ej3Q+Z81AFCQgqO
oJh8fZZHcLV2Yih1nYoLoY4HVK47/grvtbRlnDIAUD7sCFKDjt0hwfZPYOB0K1uF
uN+5jR9shutJ9OJELAKtn/Mmq8+gS0YmNrprkz35bVpVqjbIAOZQx4Dc5H1gfkB4
JsBVd0R61lSNlfSXDDH8vgIhu/Z6EpVg86MDZNA+O66ywJ2ebb4xymsQdy55PO1y
VCyM/5J4ojzanG3wgIVlCB1IVU5zolIwLzqFhe/Fpepk7zgwFaAMv3KMqScDk/cR
SR7DE5e58NVGMAy2sPfntEtI1D0LIhdShpXAsklFaW++GcFXEo6Ryco7DNB0buwA
KKR6mq0ihokiKdbU89BmLMUpHH31l7aUJsw2ANz3AoZzIF9EpEpQGYQdDCAH6X0i
epA8yiBgIVvGfEkaP4vQTToAYK16tAKgY22ycagJZ15xslfdF8pi+QbJbpnjwnla
1JNkwPqpY21gZcbz2y5WAfIou3sZDJJYDS7iEsc9f5TTBiv/UB5GTCdr8SBXCvKE
XHh2ddWFVbsY00Oit0G9AdJ0l/SROnJzMmxOdakMZ1uHgJbg4SemvD1e48LwWK5n
1viKI4HuRZDB0ELMLnNduGTudl8i59tDVRiP4pX5FyL+mzSxe9KhvpkrRZfKSNGh
sXqVoHtPgdH282OuqHqwtnWW8ZViHSW6tnPXlG/KJFbzV/IL9riNHp/yWM62o22A
L8OWFAzIPKEO47jS8dRboO/6IaspnpicY/k4p0Lm5qKUtUiVKxnSqt5uqA0UmioC
6x1FwKv/KgzdVpr0fSM0Xt2JFEFGiqT0UXvlz2oF0q4MpvzMzqi82KAhfFW+S1xb
fC9s6Lbf1P8Ve/cXEkiGyzMTgvo88LDcuGX0ngdeocA160qUHCsV3D5fScpYNvfj
nO1XKcKm9h06QcOZEPIzUrY5dOv4ewii/hSqJoldfm8yse3bbTIvp9UwuAmvPknV
b4KPh7/Fll60s9wROBcCLR+KBEPL6YNQAak4+3MPPTDBonRRPQ/Q8dj8uLVLA2MO
rKUTUhEvx2hxDXv9SfuDXkBmGvulmDtjQcyuKChHNrq9AJXd26158z8r/4n46Yw5
3VSauqVgjvx8ZbAbpeyiIv/vPY4NMci9/tjKpgaRC6VrTyE5HrDDfs5ySBxvM5f/
KSa/mUvHOmKQfqbN8QckLBbsH9Nvie/MOO7WZt+z5nS2N4RbWYCxoXd7g64aMpHl
KXlvHmCrcXzuyIgFx3Pz810H+2/NBaDgBRa0AhcaV4R9SdSUoU4nPG86ZZjwKHTK
eD7eP73dSGF4jl/F1rFd1COo7/Z2hTpdPY2WJEwagmKgVBHv8Sz5Oy01glhcaLDm
YrrTu8Z/POxQpHUzmKIdooRLwk7Zd6e2EXQNAG51uDm02fpaPYHwGXcn97KR8PDN
sNoOhVnMosJV0nqoTbBgchCmtyDbu9cia2hrjwotC6umB1ZbApvDxT6W2JvbpTDJ
Z7fh4Z32Yg55ABnrpfZLKx6g7Di4HXfBIy9HbBFeFDXp0PBq4VsoMmLu1wlCDsDt
HLWoV9rnC9jzCTgiKAJTKzVo8DRXFzLYXufb2c67pvNV3H8XUMOyZoTwiSZ/ANug
tk5xDcYvyfJT4XlYedqN1Elnx+8vsBvjj1aXiNysaGb246Jh5HMw6jWbtsB37zlW
Ex98LtFnTd4vAtAGHrP4MTBRDOyD8rx4jWzxOoaxIwUUnypiHrXF40wNTE+9T/pO
vAqII7nOCuc+Z9dzFDrVF6IiXuTw9x5hUapUuN8i0UrI0m4+VdDm1m834YUstSda
qMzsUj4H39kkO2nSMmpGRerbrl7Is01S1EG5awETxXBWKJgPdhmcRA44CjPrrhYX
e/jlMlDTLT13BGRS085cRDxIyzKrmcHGQ6ghzMKAl97LwQfbXVsjvl/SEspdj9hA
6d797xSgqI/N3RcM8OYba/Exve1uKA9zQYrxb1ygGZtttx0z5MCYwGC+E2QHWbcr
HPC4m99ExvCo9NSAkPS6F5YQVBdIbxtxkmLWkgcWHQsZFy3jLfJRsYeV2rUsSig3
RikCjxiR1r9Kp09y7uPhT3JF6K2I+zVHETjQn/a+HOETeaaZgIIvQp8u6ic45YFd
74H3nvdofU58TLWOCo7AZOkPU0V+X3EW1P/p8J/EtjKV+2bCjsCZK6hi45uxDc+J
tC9NRsM0J1blR3R6ukLiKqorBLfqO3CnE6Qrh0TTHg0PhLi5g+5yTWoJt/BeR7WS
Gg5il4PgRwsTgqxVMv9xHJMFJz55svkOmk7cZrijp/Yud4Fn+wLqnlOc+Aj4YHr1
m4ANxmKZKyZoT4m/EW9j2KXzhrqnLvFjl0LRrcX+PpdV4I4NnpO95JThd87IWrnf
qRvOqbjt/T4NaQq3CBWj57L3mPVfpdUFoJal33qPsP/HAOaKDLsS/qYoyfasWcjn
yNebsl37LgdmwxNdRNEyx4zj5bloUa/37cN3dKatiw0SBmsvl9VLZhVrGF0FHDE4
qrgdEZgCnEiqlGqXHUoZ0/x15DsUD2tujhhOaMAcg5sBw7lL4Ospaga8T5mKnW+m
R62BzLTUcN/9/NtpUnMDZT+dBHm8NNTAL968AWMMeRfAHcVTZDeMGP1WVIvoDi7L
jo5URtCS5YTaeKKEshyl0/4eJtFAhJf6QADpFkSQY/yxW1e3BdZEowBwLkaEUHDG
T0C7enkkfdCkAusM5Da9FE1hkgfr42rpshWkFi3xaSe9dcUteHWAzr1U53y/Al5H
ica8cTJwX62Kz5/hwAUsW6pZZHaIaWKL/zhFx5klUIQvDp9yENPeoKGet7hkF4id
qopGOW8094iZU5XPeRe3EWJImZF3vKWoZ1hvK6UXn4cZQPRCCerpGaKkdVafGC06
0CYmHxHWe1CGixYVnJ/f9mbZ1KgjDa67zoD39vyfUt8BqNr3hIEHkQ0GBqHQtx0M
AyieD6qdM/NKSY9rh8Yn95UgVusfCKNkJ4brauavCoZujSapzncrQxxBJAgchwE+
myVguVzZpSrcvWlI8Pfxg064WfH9+/hLKtDkqn5CWqlWCqS+DtodQAl45Lq/FMOR
AqvtLIsKvRk4eSK++Yz59ojGESpleIwZScqbK1C/FLE4hwDhczwWV3s/ONQEC0oJ
06Mc8KiME3P6hi7ElymNLj0Nhi2+5IlZU9MV1on9aIyXBe8hnqfrqyhuqECqwP+q
MoYrBYKMfvPwfs8onnSQMP/CSl62PZ9OHg8U3IMBSExaAZzj7KG1hCFdrgT+fVjs
Jj0QUpQuhiqZpYOKEQlT+kBtXQoOanmCc57oUobLninXDA1KzK7GU3dNt2fx++eT
8Otpd8Dp4pCUOmDb9nxaVdzbiQS8vwE8/kFD8OuAg/s8jtz3eFIepwcfD2kdrUiM
5z/ipoWOyKDQiaka/3ckx3ov+pLFPk3iZg9kN7NQv6EC6uBRFKHZF+e2YTrgYuVl
swT4xXp2DBgnYde3v+Tr76cxYYnCZORHZDbxFOiGIbM2xtePNY/8ZQftTS1BE75m
1qfW4B71RVUO5/s/1UeFINk5Zi7kw94s8ciqCng1EQx/qNePdQnOXpIZDOHlaC+M
bpKLoACr8GMgOXy6eqARZDfq6PTi3RiSUYpo6he6N3PDdpGedAEiUqyR6ZZCYoJC
9r+TZ1gCoX4j55vnJ0Hs2DIG2TDipId5spuItQ2fry+r6wJ78ZHhqHlz5/QS8AtU
7Rx3Ih9ZldPlJUEOxc1dWcuvfgEOypwHX/0DGjgg/9RLz+s7AlTsUVtTs3Up8Otn
zZj6udn2H9osUGGuRksqu7mRsaZiDjfYx2s/8VDOuciu8pFfCwVxIjhF9CETv2f1
QJCDOLBSqxnt6+LHvpDHPlMcBi/88cEx88cchm+gHQZLD4chAHWIU9oUjHsau0zx
WxqJkfo3c/OkphZxxrQ8jNXPRAEW5tL8aYu7Iy8SJz1LOfvFJcHVO6mgcp3ghZrX
2sMJdWJUISHt2ijHjnS4KucDI9y15aa0d25vB6MWF11JxHWMpj/3B34rggHV0Zjk
u4COOl9kwZdgjnmrDYdJHGMxxSUO7UgD32m61h8OCO3RAzlmlIYAgP66B3waXjHm
hEO93hEJcMMKX1trWku75/8eVf5Pcov62WnVBSEJ4Wfm+yYI+leayu1lx3Ag7NVA
XZkEl/j6hWhEKSEXj/up7TQK0tOSiW3rE7q44sKfaHIJTbV1JPWUrK/p63co0fJ/
/yB4Scd9ogXjhRBa5+1uoC8NLwgnlJcZIy60HIXbB1ksCpLL9npfyTgvYPLI2ltj
2Cr48g/dsqSzoAnvUSEspXQ+oH9FLzaO3tdU4xsbOnQlHd6o3IfiTQUQ5rtda0M4
yUMPyNNZUOZNOOdAsROMGyTKPoMf/EKMQ2RSnFOeW5yrxAFiRKwDp3vi6zrh6kXV
ZrmigNyrzo+2TnnCtWHDYLRpYP13U9lJ2JiYnWAKKcERVX5DOx6v1jsp1iPV4NIm
4qM89pKLKsO6WlOHUjvUxuzY/FIeLj0H2Rz09QN4jiH5ftBUzfnrDYi1E6mXsCbC
pqWMxNYWZT1wnNyCJlm3mMUkdC7lsfImKafPlmsMHm2HVachs1qv2Bdeqo4j4b+b
C174+4imeahzaPRDphHnPGWr1kUeZfuhlYVrxD5eDCU37zb7FiGuKkAdpn1pqOWt
tT44R0T1ej0WrIEoDS8MGLgvHNtUDGCMqO8uMYbsxKbyZ0lyLDltyxL7qNWAYzY8
HtMyrQNzGikMptzu51zxmKxBsrrw0hhI01qgF9NuRJtDuQskKUlv27Kd7Sjzm3Xp
QSUIIIaExkhOYfab3d37H0U4Ro6wUNGryZDgi1GuPUnSKrLbtVywsZ07mvtA7/XM
EybnLTotUZA+d2+q8dnUjJfdhQPHS0X31r1Fv2Rh9gwvSbEcFYb3TnMqb8YbX8fC
8lVIVFmFMMTw+/gUCzhFcQuvfGe4HpOCMyiD1oyio/VVwrq/P+X8x8qXSt57WsdL
LE1rSijRzitilHgc0XROBW1SrKPqkZk20zI6bnb9k/BRAOLGBGactuawJSI4+A3c
M3P2bSWrGeW/6M9BW1sbYL5HkjBY5QfVm868pJCF6HwPDqx9U02s99oNH8ofyu/M
zY2LH1oEor7Ad/4S9cEVBgozaL/smzVtBK6hsRA9KMp6Z2f1LVtNrKR60+fwFdt+
aqIoo9YCTNfwkDYpD4pQWy+QA6i//Ha9dNdR8iVTljpADD8vZ/Slp7KO1zwBOXtW
u3wjl6d5WY3vqqkzTt4LibI0/T6zJ6J5+RQH+koxGVWUmI15/+1pubbiFBtLrfto
63buHSuUXjOlW05ixG/D1K/njL/BDsqrXYXbOWWpxEbVu+Owzk9CX6QMAdmdD9p4
PSZpPl8MunoJkMPPKRGOMUrO+OCcLhWxAmj4OMUdM32pz9fpDL1RmQWoZHrsAAPx
Cl0xcp+JbXikt0uQ6B106nECl6NHnI9Kx+eNV7LNG9Vcx60P3FcnC0o+/MveDb1Q
G6QSJMnScMyfjLpBku6dYvWZ0Q85q/QNoJeNixJcDl1YbuRedvlGC9axHlJy6WWo
v2z7C7mYQfVfXrSmZ0ZLW7DyFIQcdBy/a4tG6/79X40axdq0udV/DfNtTNOGBQe7
EfsuMKlQfL+RStA1v7OSWCbcLcEk8PMFu/rRvHX1OnWHgF5dGAh/3ZPe1Dg0+85c
PawBguEH4QTmFQe6ZIl5lui9l6HdkiIMawciiLOCyVPCTmEOSEIlv2vyXkj1vgUD
ZrPY/32Pcd8fmg7BWj9mwr40SjXQO6im4p0uXsd3rMLQfkbx8CRjCGCadKCatMy/
OxXzP1frf8PjDLgRprsH9A4qHa7daahYkgokfsFebNxG1KFkk9nGD153botqhYcF
dK5i01Z9UBQWeys5JDBz9XuCE/+09cWzdJ2SqSDZ8T95uVUvGCdVAp4ps5PFUPpk
FwK6OKdZz3zI0WSV2DLIjIk0It3k/7a6DkE74N6N6e6f/g3Bg8xjTTRJ/SRGDBZa
fIOipSsu6qpmf20iOeQkder8y0MGD94m4dNUzSHgTyV7/Wt2eobH11XZCKdMLbA2
Nq2brS7K5NoShsdxQe9RTYtX2yGePL5VZ3gibAAtg1jaE85NQVUKOPHkmFR2Ke3O
5AK9wAyaOuTZidXRAjFPfhmPs0apdfTWYQ1awoBspbVoXdvb36rQNZ1++I2J95B8
TomEKs/RsxXgqTUeA/4snZynli725L8rArr6xdFpEsQF82NCCLmySIiCmKssYwOO
3cfNnDfiT7ohYZ3auXty3gtaxdheQJftpAZJEo4vQ90WgxsJyLaeFtQABgPWwMFM
DXp5iIVRr0/VRt9xD9SDTlr82hY0RERvrTUzLy4byszzSE+PuzFUGYCXlnfvGd15
bvSPqKFXMog7AuJcMdiOqPvSbsSLviw7vzSDsThb4GfWfezx99/2QT17azPZm/KC
TxROGuVdxUG2BCotG3zpncpqbxjAMfycGeoBV2aG4VDMljwXgOxJuaY/2bwAaY0g
VQUw+/rmvvULYIWuAfWdX/K/4VTAjsCmc3JDaru4iVX0OWMvz0aQWOVtNhaQSKMd
MUKbID8GvoGtUhPGZ1R3biZt0kLlVw0zS3C7KbZMrbcFOK6OFeto6tgVsIdqVqih
IkgqC2e+fFH+XH2eyyvJUP8AeWKtoXmIF9lx2XN795WwZXlbf1saM/OYv3lYlf3e
TfkA6l3yqps4JlWgJZ2IcEylpyGjuneSJtWarpo0uOSQtz0F8C8FX25lMpvWSrYR
B9DooFUlmcSTfl45j5RNCM9f3jkc/g0AHBt5X3GHm2XEJXFLJOpli3H0omUJVWbm
lWkHBl/0mQ8C8gelPtiDt8K9pKfR0IpLxw6qE4o8d0NJKsoE2ZwJ1Xw1KIuYKzUf
WMtzwyaYFgXFITFX/2bUdNxrzCvz3mGKd/cg/fT8wG8pMd7fizVFpUlz/uSSpWKV
1PqOT0XBAE8/LFe1xUZxOtd+3nDcbl7prEDql18UOcj//Rox/QNEw/fDganJI8jA
N37Cd6ipFmoHJoxhl8G/W2t3bFN44pyjr77ojCbhzsdvSC8+vdn2nA/Ti9nzetC6
WHqBJIYo7IRWZxFnRsg5r/PUHkJI/+iEWohJVIk3MfOb4Jrb366RHaG3BaXiotM5
zyKRkgZrZgTqHD7GkKhG/LdLrF/Lczj+5iDh/2gtd3dKtOyUT8JlJPu6VYdJXAvq
EHwcUvkb9+HO5neuAT9PUiHGrcWs9KJ4ekCV38FRHL3kmpI4x+qHnGliiJyR3czD
ZKp5+qSkamiB1/pnYU8NKT6urWBSrHK5JrPkUbfW1Vx7CBDrneWWE2+mmf+CXlkL
ly7aJPxdS9dpzoRs/Wba+m/nwb9F1ih++Ey8fCJCyUHxF+M3zM/fvi81jold0J+t
KOG2MPY/r/z3jdeBKKEk9O5JjGvFahKaO+YxB0dpVlcy5p0d7YrHVKLIdK7aSCaF
/mDWwOJKbE0I4kf/bcpxOkpIccTw1+skG3QdCAVB6alLcvYG1kwsPQihjz55N/hP
E8WLebO6SqNi42UPax8ShaRclD9XO48CPEvs9i6SkPgagCndLGUdSkF5EBn9B8h8
cjB27v/4ppfintcO4ouaW7A3Pqnxhf51Tgv2BNN6PHSzi9xNNmHgd/1Kr5yD+Wte
wxQhyjv44Vg0xaOM6K7OjCLBg985r5/pO8GNV3A0hDyw5pjwZFtbw4ymJKelBoGV
MSinI0gUsTRgaBss6RU8vZbRvpoNWNgbJY3NrsFrMdAHa7YUxdQ6zl6mosOcnACl
2cSLZcK7aoQximln3yy7j494LkXb+BSqfi5kIn+/QHtCp3c0ppV6dIRfHARz/sNf
NvIbojaqlUemaYG+GM9w6qgMYM2Y+ymEOpfoJ4oLrw/LCaveVwlFSj+AuD2GpHi4
PAk5mMoCcslBqg8rI7bdchj+/Hr+0tXX2FDbpRElOP8cxfM5EKCEAW77TiShY3PF
2bKh4D9Pysv407BZ9i8PgGA548hMMwh6dRIZn6gNZXR7YuSulZe2WT3/Kx4Ke7PO
2csrcaXs7M/0EFRQy30+LOmrKd80hb0mAmDHhn++5rW+6Riepj1rqj0NhpjvwdZE
cgeSC6wi2OVqhMFUq8Z94nP47Umi2HX9h7mTtX/VXFXTxl+sfedS87m3j+eUkl9+
RtUk6qG5gIybuSceDzAe6PwKRPMxu3qenga0U0j+mWJ7GopzLgln93haK6vnvkbN
mh0N9P6lIIvZj/2ABCknAmrn3kcH5mBCU6q1upmi8D2LPv6xMX4hnS8IGSZVsSLU
I/Py1uK7QiSqaihDgIFYS8V2YmZQHGBEtKyg5vixz/rFZqxilV6D39Sdqos7ojJq
xKgJ6ciIT+pGQxOrU63acbPBi82QOouYzhsbfRhrIOym6EGE6XrCC2h999YCvbKr
1R+8/cCjVbn+fgZFDtdP2IrsOYToGdSHEALFyXiHo+8hVUDHCVgrUUmJFNLrW9jQ
FKMOUx5DXqueioijCc+7JLV3VZmvcDK1wdcDzK/X8AyLOrhzexMimlAtNiin7VI6
OUYXjum7JW5GcAImLJTL3yjHsiEEy69O75ZxOvk4O2QydPfvbBSUL+s+ARdB2vvT
RLp5SCgG1x1mQixf31E2WwHB24YhiMOByhvc10MZNtoOmWyJNQZdTly9dpWloF1H
1Bgl6uCWVYW8+HKqXTfU5N0aTYmPxdHXx0OcfjpHaRBpg042TULx8ykkXf0hlGRI
zguLdp4NWoINBnW1KgRvx909hqxLDcqOlTqSyFQAMwi1D9P4VXQAeu3MiL6bAYCW
iEnJsKPhXxzG2hfbCIXCB85DXHuHl1AYfh+o3sWBq2pRWmZgVudcO/kmivZNnTpo
XgNnxI/E4RBcmYf40WZP/jnzuxTQDl9SGxVlgsK/x9DdyY98lqLxUyAtxAU+Ohrm
jrXBzOZDD/mYHcvdf6MPk8d5JnBXkE7bjApHwN7z8NQfPOwGP0Rv5KvibnKiR/M7
ZpRiEDygqd4W36t7lcz3YP4Y1PLcFvCbR+8UNtB2mDPszLmzdSTO9xzBzEKWK2O/
oYmSjJh8f4r80U/rLLsjgdw/fzIujfpyf9hWfVtavcY11nga7szctdeEfE+xyMNc
ca+ocYBgub4K0bFPxYd7DeiME4cIEQN0WOfNIWMwBkHum4QZW/l2xIoz9TXI55rf
hxUXyPNINGPiZKVsJEgsg5p3ZyACYPNIq05WQlulAWjSkW3ClYIqeG/613eiZPDp
dOZFnKZ9zOtzoR5lczsZ+umv2KCNu9Nn8ZNhPhTI4B3VJKcVHo4yfrPDttIO53x+
m/NIyiXarbhINrh7Lej6e5f0wIiJVxHrE7VVuzJlbEEzciReUqGuzW1O3pR0TGRe
PP+J94OMQFHyL5hG8AedP2+m3C77CGIkE2+nx6ezTojRQDzgxvVgb21BY+f4k8Cs
AHwV96T65z2pJWnKdkktHZU3lUB4vqghrqZNHO+UzN7v16he9SRNmAopkqJ1LC8R
DbsfTyOgH89XeXJ3g1ttXveJwXp37kUThvRKa90HF690d/63yI49dZtbnlu+0+Wu
PaCuHvdS1tJPq0QRUax5lOWGh25/3FzXgrb+l1q4fkf9hwS0XUmBkahG585dLQI5
bRnI/OaNV6Fm6vOBHgfqzlh0aiR/C0m+xX+7A6F0P8MB5viUySJlG2hjDyA4YX67
OpJPh0LlEuU54hiRsv6ozfvIbvPogUqYnWoN3Fgy1urTN2Cw0iemv7LJLr9dtc1K
l7jZ23QNBhdpTExSCkJbN6VvosbgZCKID7IkY2wkEsJpgMUH9I27mB/bi2lj8bcJ
d9N0g94ssFXK8RNEUd6y50nVLR1Atp7CfQd04A4COc48z8+/vb44giEYE1KkPq92
JLLYeh9M8O8ItAT1nM/9Bwq1TR/P1K5o0owhIIcTki3/FpajptQSlAOpysLqaJoJ
zSLcH9AooRlqpX8r40tyM3ftmGKrJuayU7V3hiHqIBYqM7+tp6qvH/Ot1qb0lGrx
sQVgbp40J4KzBmmseigooYoT/RhQNc8qz1WPzuVtI/MZivtepW+dh1af8RkqEytT
TmDMu6v73bVbo7O7H2M8VVYr/tjBDPRmZ4Z0jnXCM9NuxDfBqqoujMqOYcmj7nF7
am9j202Dqdz1g5RmAq8yM0VatFT5PeDBnsKTCmm5VJ/L4FHKHU4tuqchnxc+hooq
UKJX+YaaIUQcCX1wlpOqqdmLXxpf6sQRZe8MH75HN2loWsuJ+hzmOUU4L123rsUI
FDuQ9RC0IcWBXQ9UcfHjYW7omqNynk9c66/lYeFd4zYDJw7kXvVZKksubpiFxQq6
w7RVo0WqV+Hv+kwZYbjfdWaMXadwGrqFxhvutp4Wv6W2e/kJWdCmNLsEjc75vcLU
5WIeyOjxMtVMhFPAfnlIa0u4sxHYY1YPjZjkAPNv7PsPT/6KQVUEyWeILFpKyaht
gEjYHaU/xtpHjjJ/tSfrPtMzgG6NmggYzAr/JZKPdNE+P7urUEHodLNvCWz0kQwK
UQReCxdEQFjIwhvpZ8kT5RSok08L+eObovqq5c1MVqOFWU/ssqu+Ki0aZ7XmYmyU
otqWuGzD+NdqYcLfdGfg9ukgcPa9rrBY5j3Ek5iZtIqX4z2ynWbdFKsXjTIUvRPW
JBNY7DafPiSReIXUe2nRHQmevzwGhex4jGGW1uEAPP4PKnDU57y6zlE1ZDsGg3gV
xMhLajhyB6c99OcuVQqu5CthP55c1aOEqHN/6rFsHnoBQEBukUOzAUiRNatCHXh4
BtS5lFE9Ta7ifh1YFKbZsht9os/0MspcBtjhoX/atmKbgCtSgWkNh0GZxmYjjijX
BnKR+4FOz+FBFTDfaq+shP44taFI/vyW+tfbKtzGvsmsbRpPuetVJJ32/QOvMhes
yK9FcMENkfacDucPqu2dE7ttpDotSdIiXq9g/D1NZ7Rd2qyv2nBZWaoOqhP3MCQZ
Y9iXW1nYd28PS3tlLKr//RAAO/vBNQuNPu0YJcPNRGANC/PvEpS5vDNjaGQgxCfV
I91OKxlNa3sMmiNd5EEmJaza6e+zZ6rKJYN1K6pHJrebQTOhuKhcI1kNRJfNrcQ9
D3dd0s74I4+ggxTGEw+EpocS74vzG/8j687k7TF0rVwC99+X3SxhcU037hAxzTkp
Sbuddmdx9wzBai3one09N6b8bWHPy4NA0HUaenGpuT/qFk2lnVot7ETe4/fMtCqA
Od1Yawa8cBqjTKb4uaiYrWXuvQS59+vSyq1f2uDWtMJ9q/rj/nZgEIJPWVk/Fi2b
7/qW7+NjsDeg/xsBnKBHtHy3GxFqk2iaW+gSgnd5i4UE1WArvBuyNsbVRhWq7dwk
i5ol7Z8aIt96dVDX4KoM3wya/xj+Uj+iQKqv+G0qUW9LeFoeNqDLJ9wBvQNKnYv0
e/hJLqp52+xt2Fwal44cV9WF1enhbXk/9EisLH5jonEV9+YW3vmKs8QCRGk6a6TX
alNdht9DMR7enU5/BkqwJWrVSTpoApBWtfhGaN7dFSaeHyVbvYMaacxDg7NUDZjL
Wx8ZPGxniPnZQzSw7ZhtpSslJJXOSbsZN+L8cD1TfgSWwi9ZGH4ylbvT4um5feaP
6cFKYri56Z01o1Xj2jHg9n4Ergy+oe8YacQmHz0mmTH2OTy/sqe2TSfaSf1UrUik
fP6AjJoTVWdH/5pOZfdvrzcexG9mcnfGNAYx3RCSbvVAFekdR42E7CQxETzGygmf
hifh0uYnEqasF9js6EZ1DW999DRckxAEtWS9tZZlg8BGVN6aqens2xKHRLPEv2p3
nH/t7cmfDBI1xHPPJq7dx0UTPCYYFb0G+z8B7MuSL0m57hQOf1HengVwEChMTeu1
zgHt3w3O1vQUGF2upOOh33YwhBTW8OWkDJbjIJIm/xfP1uqJX0O1pX9CDkdFnu1Y
M2B8tX/jcKn0Q2kHh9KoikPe28kA6yMc/ufv+wURKj1ab6d31Q6KKkqP1G4vOX+f
nyT/rCvuibG7zER0apz5A3KlBTTkR81k/0JndagUm6pnFUTdOwm4tnesloA7z+M/
Wwe7zaIMI8nBt21hrBM6WHkqixXEq8v8V2O9E7ZrRv/eJywPihxTkH6Shfm6zzFN
WO5uJrnqv0wELEXvhOxbDWQphZsVpnxTcNo89/2RBobRXUtKS07H1AJFxkyhYKin
w6eA4RnauFFgYG0xK6tI50WJaM59dDu3/DeCUulNaGJ4bqHxzjjtO+QIi9d/pxgr
OMhPX4TqcYQEtXBKQDBVKAQdgxfOzhnPEb5why231ISSYelosU1BPO9jUDXbg/Jn
ofGvLWwmAM1O+QBrbYlOmHbgri59VMocbM+KXJqTwCiLgY9VZ+97E31PULj8fguA
BEY6ai3ZLKhNfDQoQ2J4W3h5tegRG5wUQt1S2XYCClgwOYlfmKbHyCBrTo0c5RKJ
r7LDpW8hd6bg8o2QPVHvdZT5yWyJQQGEdToSa2d6GXxilFL1d5PzIvtFyuFqOUS8
15ITMNS9wEoaLcoUqx1qQm0CvKrPmqUgLouzlik0VG1cI0lNp/NNRYlyblSZOYqo
jsBiuXaRKAW5sia890JXQUuOk4vBhjYkARqv1DYUAofVwAAOrn5MdT0p/I5/K2FP
wCcGpdu5iY+QUazg+MAMrkch7CqNhhv4DjIrN22SUri7W0CET3q1WQS86BWb5FYS
HeXyykxn7FPgUBDcfEM7sgYDZrX/Z1ndlaOyoMQ14J4J1yvIppjVaMwq51Er8qQ7
cpQlfutTb5174G2fkutLZFkrlCnWmxuw0stZf5KhyQf3x822K0z90se4RVhdcTuc
DytpG9QnkHgsKpfhYczAm6l2y1qcSJ87J8oMA2EzS4LqudlKpnuouSArC6GYoXGk
pomvVF26Aar2Q5EdzAMd5izgon5yrNquO6zvzkUWyOooNepCluUmlclcUO3WIY4f
fIWJZInVImylVj6ABDIlHhzvy1PMius3oxSNolh4xmKp0GQNDc74O7s216gjgw7p
yN5twTIckn502Q/k4WwsQV6n6YrH/3g1njLqcUu00rl6xn1byoRUNKPXQ+gPsit+
IqnweVTOffgVJhECc+vO3FyQbry8hyNFRgOB0+JJy+bSTWXdAb3YnpDRRi7sRfh9
xnTG9FuewhpVdRk0VFi5aHJu+eMdZoFKy9CSpexLp3WlsCa1PceyR0Mc3dIVDHxz
VFmKzWJ+jKtpocHSq7AN8fFCZ5r1J1flFvNUTcUs7utKuN/xxislEt5YPbHyfm7T
OmLRA/I/kAiruneme0r/Z57Aw6YxtZms6XYM3p6c+mFWF/YYNmD1NeisNnTxO4xI
a0EbP1YRjxd/h/pdHZpCS2LlRkKNTmWMDrmEHmA5yMtPf4CTj1TzfiAiP3Xe4fUa
8XJtX6fKcwrbpi+LK0tLTOqKNO8SkpAl5kdyIfF/i5TQBUnpjnKw1R0zw9QoxnwT
OpzlpluYcFmmHSRdtr6HvK0/5Vo5YFQ6RGUr43roCtVXipQoE1GsvwrAb2RG7Day
7eanmKPzxXUdwh2lR02maV075SQPvi7keZESSz/vGt6Fedw3J5d1hHHl4BvtSGgm
eJH5+AgEDUHY1PSfJBaqFsiPyfTdqDjB2zzrHZdge2Ln6f3t4rzqq5nwB/bgOkp8
swhve5ydZhcqksPYzOj/JWe0eq00QJmCUVTnbu9ueOyvIrdYIB0WgQMKZ9uglrpy
E4uz8DK0k/tYK/qNGXCnDxClGPe2IwKETKMqJbSsuscLFVGELkwrKWAojLvyycLS
6UGNqZ+kH6LCZpir4ESfEKqzwkMe+EDXwD3DvikkNAvcwzhu7W9Ps/3pW00VO2Kw
8PGyfg4NKhuYHYwSlCV1w1kks8fAO6Qqc1evPTsaNUJFsuw8hkjYa7iiJjwIq4h9
mcNVQ0b20ZHQxVw5FMVoVYtiarcjB+y917WK6y2yghmp36g8AGPodh/OuUl31Awd
8YqS2MCxlxQRG3LbTtYEOPtAGWlM2Wd1wuyMlLPAd1r/MJXw2a7zmxZZK1IRE70t
r7pEGHjIBYs9qu6yH4JgelKTKaC38/ZNuaHuUy3kJvzLLHFncx0GXjW5H1+ejkK9
HhSCVYyOMH4wxtBAF3DpScYJNBKiGz1pu3jjG8MwHoFAAD426ifveqCBvGhMHGDF
pX0I0JBp/o95BLe0UIJYsCxUSYQgitYEFuzQoqcKVUvR+keq53UqlKcUQG3/2L+V
1JnQQaMowy5s/929s9OhRUzCG6HKEtWaKWwGyKCR1jGiQbML2L3K3X+GybPeyf7y
tWR9qAukq3U3F0OXcNCIJ5x+WuKqnFlf6MynfMEX2BVlFmBjuza+N8pwxzhpHVgM
v7CJ3UAc5a1qRqbvYPLgzWZp4tGiR6tUAxPQ4ow+nAG3gBx3g2I641t/SdVwt9g7
/xt58QyE03irrlXMoPFY/jlLKJL9QIS96z1/SdKDldtouHrPUyjAcq+nAeT4Txa7
RWS4tUhqul+tSw04mjurX0OVFdEH8kYTq1ga7xZ6qWafS/llTamGUji7l9MrwciA
55QLkV0vLU0KxMlOYW8x4B3W7VJbaCfFqBTTRyI7YVTloZ0aSSQW49ejuvOs3uzq
tSO/aHXW7F2PBfHSLj3YJYcXzkl3caddl1CBWzh/Ny9MdAEpuvOSNiOsJ11S7kF6
R/0xdLphENdhfduF+Am/oI2opfQE/XW8VW2LLkaR/2NSB3XEG9JsigNpeuiBAxmZ
SfbEBQBjdrfHPG7fbWaE7PuyYbEfYNygvxUh+4VebbJKzf5c87teJOubmj4P6mmT
P0APFxKhuipcyIw5VoV3qUuo5sYPt4kEhBMSZBcOXXujFvfNLbkElMvGanXdrXTc
RD3GDnDsbr3P7FVCYZB8Mzlx7QIF6SGRGnaV1n53tbqVF4bEVV5uHINs9CW+onkA
V9Zpke1W+s/xpWWA4RXEC+ctAR9rh8dizPauk+/MmQiKxePz47m1a1JDHGp232ud
/JjPrxLUjysCFpiyiWBCrHjzOL3uOHTvDLturZF7HgJj5rnfkdJbz4yCTq+hbuYE
9e78oVvd0ZehOz0OAN22wgyKYGwMIW3YncA6HIWeuK2NbI+iLwYzWRKBqc9PDsU+
QxJr1wc9bcLWYhOlaSbEAh+GAU6obsIEZ3282Zlk0ol3qD8dsje3WZVCIe7G7J0l
TOTksBs6jqwPdQHIpOoNaDz1GE3hrVMWCAQ82+JGXtnPjIux0l3/hJboDC+NC2FI
ZXrPT8IcUBEUi9wSbZPUJ1V9ebhbeSk+ooaIGAr4VLhY25me2MDLNfJR0rP6iudW
7EDTuViFvJIDcDVNDw87fCVJUpdNrEIwc5B9t/+aoxp7YlmYoKhJerClXoRdDgOQ
6KRU7KtkDCPRYcsB2Xhn4X+n6EJK3Ws7fqD4/VPxVn6+uxaeyEKo84kKFEUxYPtD
0FRh5I52yKJ4Xe1oUIg2nFOC9n1sYNBbZLOOqXPh5E4KuHM57xSOJp2SCv8ml3Hz
HjTKTvv0wLGYg/BYwL2ZduKJpNSznmK/7hiCDqKYWJaAb9Ys83LxeLT54icp5UNb
4sGrmI/Up6we7J26tJhex4ieHT6v/8ETGSdfaxOQ/tJILU73oodnaDqQdVsMIcrL
sP1M1LqxtIMAnBHS04VRWARykg4fyzlU+1xSZ81XYYzRruuUP/mvbfcYB7Oi9YUB
z9Rr6XZSWrct/1EJ9S7j/UfO9eMqWaJ/gEhqpbW0MLN4RdQiR9ApL/nCefio1M/E
HqboA1UUoEgrDHvLuuh7tmE9YTMfQOZ9O0XG5wPnKRzqOhCA/mrzSn+wjQWs/WCq
R1uhfrUtJ/IBUbcoaWiT37URD+7tfDDUGevTmnL7bYkLEQlfm2tBRiIb6GnGQciw
A6OC8aBvj+cM9fl7XG2u2IkgcEPGGBauF6blFuGKP1kPaToI5xg1PaV/QBXngHJc
bcpzw3K5unQfWFN+Idg7OkwzuU/cXODz0tnAi5Wk5fnSFL+ImIs74nz+ryMKd+AD
1REtXJnlztZu8zJj17HUPZEFUeqj6FiNztMYUBqKj0NaekLJytiGt8GbPZO52Eop
ynThOJf9iNEs+V62L4HB5Nlp8x3NY15gU0mdw1h75MPMkyHXZkjwVeNwVVFRg30o
9Fb0yn2CJ4MeQTFV8DYdRwpw/QXEAyC8pm4mTyuF5IppDFwsHCLLhd3EA4ew1g+a
8M9ebsfBIH1MbQn/EcH4pAileY1e3RdOqSGyxYnlRuYm+pD4P7GlSY76cgUd09m5
HiepNkLGC/M2vE7IFdovvOUYvwYBllr24cMaklWvWIFy/3AMMZLvmVo8SHZ2ZKvt
7lB07s+nJGHH5BcugW0LIZ/5e4dXpnNTTqvdjx1xyFOgDYURZxg4HjDR8gU4blSV
oNU4S0ey0LoSeYercPMuiC4ZSWBqOAMmhKQVUdbS91fnp/uQsntMB9PqN8jmldmY
Ya6K//9nn/SqfN1LxKMvu4JSrgLyZ9nqvzAM1eI5fOqr/JALN8YLcIj1FE8OExzJ
ov++zM4HY80ugHn1BQ6OFggjan/Mlye56KemYnZy26hD/G2QJ8cG9DSD9Fzklwha
pjFhlZ85BUOGuSHXTkIz1pn1ZsGdP0oAAa3OJWhl4xB3kg0htMJsHOsE0J/HAdbk
/IVgHIpvjmFg/YQT/xt1omQCNnSnBP6gUxURlECqC0QRk2VTNF3k/4u/IVlS9mt/
MhOig62NAKECJPwLiVJAN8WMpBT/mLfg6I7eXLNzSOoGNCBfh96kgZn0BFvSw3ES
BpualtzKt3qCdRAYMidtuU6oSrxoc0bdyqL+0COGs5W4Pia6z184WlFQ0ODRkm5A
nD6apnfdMU7UbPxC0S1qg7O946jdP2ezGKcoEsrwluUUcNVZ8oWUwTlAC3n2eIqs
oZJMR9cVIKGtRbGUFRJQEKyO0CHe5Nkd86uvljuAFxYL/4HvlJc3Kc7c6OZeQIsQ
YRiCpPIvo+fJ9s7Dg8Gd9uzFPHqqV1ogUQuhZHBhAyOmw4KgrWIhpXX/QxQwvqUO
6nd8XPN7PM73ZcLyxPj3v03P9JKRmzXq2vmy5CKcFbbT1+layIMcmlKNPYgwkHNg
zU3zOP2dI07D3VX4ULD0t93HomN/KZv6Lj9+7r1jz3PtbblcEowORmQCooSB2QRK
pcIWaUVKTjegHmBaOC15dt5zYHTSEAaP3tnMEJMs5psERaYYJfLjdXfZGTtBxuDE
CPJ49+1mHv2BoOEqcecBUlTCtGLpg5oHLxgTbNQVTAa7WXatihxaTvSK6b53TZA8
nGhDtQoh7xdK2frfw44J+ttAI7m6O3qGKdcdwsTTnyJ6H1z53sxVfOvEXytV80ac
dLjMJhTD34KMsKtErNo5ItLCzXXFnyIwfStv/WMc3712tzYcuSTyJkpIepiuouy/
0MxrGKQ5KeXNLXFYRn0zwDskLHnuIAanMP0UZk6WztQGQbFKmgM2lNrVLbelobUl
MO6wc+c6VA94OecVKZeXVp0AAxxDnALrYWeivUbZeGclE8LNceAe8e5CJxUUQF+d
moGN3fH+lSIBR+DeKSo9wVw3HMnNlF5QOI8iy+0v5a4Fg4kD9AH8MPeGTXbux3ru
+dalbb7REjHgQsE/rNnPrksyA9va5KQoxKTpotQlUh1QPgnymuXtoRTtl8x+wYBl
A0QFDWklofg2haKFhGoKPVP5fxtyYmn+gEjy58L5eXQZe3J1nTCaMmMzFeNYq48K
3y2JM9pTNSDTbZoSxtu7TWhVRqKCTSxny2gLCtMXHjQSNDxC4rPyRpu/VHVzqDNg
hV4pfWMlh/Rn8KwZYZyA9ntFxih2yqvzPNLut7izaUzOtvK45DytHCT97FE4+SvI
HRr6iwhygqVvPv7G7DvdpCrAuEgN6gQrduxmkCNEDhobK1zpZYNCJDEnT+ELPls7
U0YE2PAFwNXhNa4L4maS6rDn1l2ybLGXqbAKvs5ebhp4huT6Uy4k4hRMNNUVDYrI
3UDzNyEnc0qE0c57vqNJ1dvRkOMf7Pa5n0Vg+WUExEhyAW41HqLjuztVQfBYZVgf
FYM8kxSPFXC5OBfdXYzL+fjVGkc4gjvZpHnDUuuVnw4Pv9NYuQYoVR0cmUOK3SlA
lSeITJneBgkqNFSJlPswjmXvStBYXsLYOF346rpj7YeutFSgrZFKpxjrf7zXXn7m
t2ruhwy0aqZyICL2Zw8tYmY/g+yQo6x4biKH6DfaYPXB86gQ5Akj1CvgM9tjbJ9A
Yo6LgNfUVfKOTwjEvmSJC6uKcJ5CxXxHtIXfQxxM9VheGuB4iDbNCBxJbIvj2IsU
5eOrlOZGoBc50chk5FWGYdi060Lsk6sCQ+qoX/7YWLdv7AvA9YOcCR0Y2s77Lzgj
xkmYpcxiIX0rYu3TBdNGr/wMGQW/IoeWvREwJFDPgrF0rzfPsBYAbNQkYuzKJKa/
slCCSDW4PzJpdkYWN1hEkpauKk77mdesSEuRUKnwkiIa2VFvMPfbhO4ZE9R0z3/8
Ifs9UOTwwtpa/G+nIy5UUhgKIuPtT0mifCeSYmj7P2mFTRH4CVoWB99+CYN8l4XF
SKB5jxOmn7bQK704MY05nt5OGPQ0533kdBGhm5qulZKUOZFJyM781V/ftyWFoIJe
vENf/+ht4AjUgdQVrdT14KB4BoHCDLgGGnn3px5NANLYlIrexQ/AotmrThUKXK44
tWLiHDdvUoX/S3Gg6ofKwG9jp81sgqEceB4MUQk4IsGWXkdfmMoDGEjNsRTkmhom
KDPGZZOMK1pvoSOK+qrRC/9lJMP0XFS9ieRqTj2EGBbwYxbil8hk0+7SgFV42m7K
s5SimKtrk2OdgR9r93S+xKRsze8PGdn7YPHGnFTMCtd8c3WUuji+aMpWo8tYYYra
jPPrzlgo04rfNXJxsy84e1m23DWifEydIK6wZmzKlskXXqy+E7F0TTot4OV7N7JG
GqemsvMguBwF6vN7WlNtKRM3AALFA4HbIBcH6qV1LfvxR1rMDcyXlw3qnCGn30J7
w4oF1beP8UVbDCBL2F1Mcha4gXiTl7B5atpad2Z/KXfAhKM/SkLhp0lczrd5YPB2
S+cp7kGNqE1zAoMme1dQQn/Lb3bqE0llvAiOM4tHznN/bandP906lcsTBdKinMUS
OAlQR6hkhQS1ucxN5tJsE9gWE0rSJTz4FGDylatnkuzBZEYoaStNDGnN4+TjCMKY
EHRdgGgKm3Cz6RalWPARJcH+6eTjn4kSc1eC3m47iT7UVD9ag9AaFTpfz2E3Ni+5
zjsa0lrY/yKGI+OOVl5sVzdTSp8z4W8AgtkSyQ0MiUHHXLPP0MNObH2fvLYPokdc
9VGXoJ04UwgGc+eClTb31RWd3xqGIO2/+wlZdYjRhB6Z/t9BLrPo3EByxLC7IoGn
CiRLvyRXWUl+gowkFTCZQfGdW0BRSlb92xu/01DLH7OQk2/H17Pnz+8JJ5wEqqwz
fTeboh6wyhNjyhDlehhzgx12AeoVyWuRQdSDP/WL5Jr889eLgCdKkZwiMfoJh4IT
uotDVphJ53WCZRBNNqn656+vJ63orxKzjeD7palFQ8UPQ9wupPFDTogqSzeDqr7S
fYNoUOWVzf/t57GRXyapTr1dqMktRereLeLvuF3mLeFC9Tj8D1fPk749Hbsjejw4
/luQRuk2ZAq7U0i+kUojRjl+uZO7SN7Yjo3RiVoJ2Hrc6facVxJpC3CdHbccb+pv
2gULjNMCBlj0jmIfljLbDyZisTycfbK3jwfDkz2mcafLIMGKvRKkbeNloFWQK/7s
+rfiZKqc8s/Ez8C2jLtAoFgkiifoEgWP7L7Ossvixbt5PBx/ohHQIijtvfq9OFrN
qMFsHvcsGesbAFAQ7MAycIXr7B6Ct+OsPvMnA7rL8ryDI/CWQ0Yk8ilqwx6+IWcA
QmJoSlV7zeNLRXewmbYDOeXS/4p7TWI2G4CXKk0oI4sil/nEa+tKNx/Spbr/yYOt
H7VRV/HSJkDTlO9QdjuylnIvClcrBwp59g2Q0c70sfll8l1QxKRzNukQ7T98OHQg
s/7m1gMlgIu5pruOezOePQ0NGNEX+uNPT7Bkbz6hV2zFGjToq2L83Ivv4n0WPDh3
o4RQLDrHnwape58ffEc8ODDYe+Rm7f6ePykEcNAvIhqs/53x3leqYD/ceW4Aa3TQ
Drpk8B//8xWjD2nOJtRgRM7zlBCvlOGHWtw+2+IXS0M/S824b+SUiw4hgqz/ZrNB
9JA6X9ggWxXDVyEKb07ZbPpkzYlXzJCFJQn1Bam0BgoVdjt69n0eH55sdT68eMe2
AGe7YtfbKET/0kA2BuQ6jveSmr3dP6h6woyIWWvn3DMw0YxFhWSmzGg59RwV8KjB
Jpk2NWIPU8Drthz8xqvDwZSOhrbj7rs3jtpjTR8v8rQ1FoR8UNyuQEBaTatL//zt
ytX8YgP78V3I0iQ/j4f/IsiYq2+6ndHB1X447q8NQWaR0lKcoH7RKkrAJwJ5EmEy
NPW1xkq7T0vqfM2U5Rxnf3Vxei+gEnghlTEgJ7FMW3Rxf2ksyi89bCqciLNXlStG
NUL/iXCYkrAsX+LCfU7QGEXnN5qoF7/xLyjiJH2UdVz2EHbB9ERSRNLcfbWEwKeO
yJhetNFXVPtSh4j6vx2mRy404WGRRgX7h3qfR0x+UpGhDreCnBAHclqVe+L56OnU
b8In6bT+9xyRW6k4tW6oKiTrQST86wSHtimQNqNXvrblv3i4j09fv6ZYjARZrPy+
pfy11zoWhQGGejBMS2metZ0I7ym1yv54qzUTWphuBUqL/8YN29d0iRD6zqkw+ky/
+GTK4m6Ys1z9+ebQW/qeYGdORjYaYJiGTyko25E0f21zBi1Bn538jc2394oFY1xT
TjICxnzNaI2zBFSVuaDZ76MbDxDzz4Lhkq/ehUc6NFW+uj/K1MyBZbwMgsJdl2Lj
kyaiLHVYDMWq1WvzTusxXuQgtz6Un30A+aH942lpYr/94i1Wo7CKjE9zemjM6HdX
sgugcO9eOBDXZUqTsgLUMLiTH2PewH9RY+m0G9p595S+BCyzvu+VBOXJy+FW0YkW
ELPgznxlA91PYJzA2jMXvZKuQkt4OaePr4Hr8SJPnhhbH3jHKRUJvKviRdksSt5M
2HgC7Lc3c3FwgaVJTjGarZvjbBF3B3BmdGAcCkv7iYrDLGiwBJiTGHvnh5GOtCjL
0s+BEqbzre2ioeA3ZIan7+IGRQIMe6MzJUiWKWzquTRInp1/hkpzu8wxmgjy87re
0XT0AzxZpRQOAZ7WhPwNFYRqoDL9ID6Zpd83tah6OJNf+aSpeLe6kmJe12DTOxw6
MCH5uT1OF7sEQs0hGHTY9sugbWwkJZ5tj3mXdfEtAS7VbTDoKT/y6xVULcy/0te8
mQkpggQpEHPyZf9HQQPGYN8wz2OGsMsUT6GDyh0ci3YxeFk0wT+WK6e4U4fPuXGx
gv3JDYAoNLQXPKG6KTBeN/D+UB33IcIaSgxJ4ZSazzCqgFMEmgc+dTrtVweR/ZD9
3Y2H1iif7Ik7qwjxl7Jhi0CbbuDl7M0QLM+yXmY0XU3JduzNg27stwG+cLsi7EoG
M2l9Y7ILzuMOpiujGD3XgIxULpzJymYXLe+tsL9i5KpGXvXTPe67OvCvIO8V6fu8
toVLo/92HeVoJ7yioRxiC8cpUqY7VkDTCQLEHvTMv641hOCFXR3zm0Fg34RDyFrv
nv0bxf2vnzv+As2XgL8OyeCWsB8rsetnKXXnRpStKtxVKLuDA4HZVkxQz9dQ5pwr
iQztax4WmPUxgaf3biQkL33b4hyzqiMzwN+koIJ0ReWnpQCJta2sI7Bt+UHzs/lg
h0550B5vE7r0e3i3e18mjs7fOP1ky1fES+Ukv1qRP0MVjG10nN6LaTm7cimhoONJ
oo3Rhn/a8pwmqzegSqpriCkg5s1MwhM58GedFk3EOd6oRk7kVc/5N1529k/RngmL
Wial0wzf/X+dLYNrAxJvl6w24Cq/IZh01H1XW9+T73T1mS3Qs4dTA7p+Zk07M0b/
kInpTtuI/MHvG/Fe656j8GhMk8JjqLeIRKollMtL1DHx2Z1OLGLOCGYQ5X/A9fBI
5KKyMMGW9TXmVORiz+WbwMwyo+/qS7Yx2ogHvmV4/TtulEJs5c3R9ZHfyvn7dlZ2
rj5ea6hlbU/tN26/LaF1fGAg8OTtoO7ThZT4bd/x9RrNgiaR/w1Yap1pePpFIkAo
uwNBS6PcTxwewe1cRRBmK1EedTfMRTH9mNxNk1vjgqKjXe+G4wcheIg4QS4Ia+6T
c/9QNaIZt6Wrpti3AL9DE5ozt3mKSs8wjgdEcqs5AmUQ0mtqTelNNa4ELt85rwwh
buH3Wms2xShGPZ/OBd3tQKl9XM+f2h+bXrU4ZIbM+Atke08kvQp08btwpaf5vuqQ
F/Lk1i+uVHnImZif4sOXOTrjuNQ3NfV07lYfuVFRffUIUpNvvnkP+DjgPQYhUihs
/gW45L38OUOlDQLpX9tQzc4Be7SB91wu1MQkwePzll9IYFxtLH816aBWcM82DGWW
Fzfpjap0aXje2Vwwx5OcGuzcz/ms+Gm78oWkHlVhQJXT/VypHLHdBm5+/DG2V7Y1
/RDwTEIDP7JPFQF9g1Tf3yQ7ME8dQOhFHhvQJGuI4uaUyNzl5aQBi5PkLVORoe5E
wpA9AgOhAjyjp+ehSMYfKVNwTLEurtheKiRRdskYWtfRlidG+3j63r19pBU8We+S
o5Qur2whNxMfWv2EI+6LzTtNfxvmYo/fLX76JaxkhbkiJKNd1eyw/u1DmXRmpwx6
4Hr41gKYZQDiaZ6qFl5IWSyFVbtkzKzWKM4CVFs/tv5lojSbMNjXs2bRavTQ1E3i
2tde8bb9qMR1fwMVq7FraWG27wpzQMclw/nxXar6i9PzFJB8Y9GolfYXpUVQMfX/
resekT88gWju1CMBIneMN7RWS7174wQ0M22gTrluuNJn5QLKQCRtmXWDtSdAg3J1
qY/DmF/ZQlTKpqx3/wQd3xk/RHCVXal+oBuuZzpyhfgIdnHFLYAIw/3NRF+glsfO
5eIOle/2kjFgVxq9zoyYo2Ap7mcfx0ZoXy/BbdA8ynka0ao3KrQnGcJvDvvq30+u
c7XdmrDx2G2YjsH3OpDMRUgmsn1YyevXJalbIjvt9n6sedhyMmnLoSVvhrGCWd2G
xUMFs/HAK5QGr+0U+ioBFuZK0Y/zOSyemLKGehDI1Q4BBOkeRY9lu738CgFDUknA
/3SD7/rbb+AiKaNb8lHS1jTvsx5TSB1ATC+ovrRxqpDROdPsQmjXezwdzpRGYEpz
foqWLf8iDKNauScXdYu8of/Beavt7lbGvs0shlaPO901HtLMR64PxiVZ6ZQE1Dlj
1j8ZBlJtZhHbtAgkr7IAzM9VSfJfFMfuMh/vLZiYb3jhCHZANpdd6cbG5pjfiYo0
QzvpCy6cXBq+wzQV6qpoQeuAKvqhfe+dJhHUjV4hfbt5HIcI1Hfax9XzgoaTzR0G
lYWPiizHEVgipEeC2e9lU28f8y88TiMnFbm3WVYrUqknn4LLv+vGeS2Br33XyxL6
n2n7iTNJGLbe+MhUAEDXyXjq4Nlr+ZY9X+JD5aKho9AEzzedAdrs1V6fIw1/jwi/
+exgS74VBdOuYeFpecm0pNtOYebOJE7x6gSH7CStmrFFbzMyM0RiRCLLY5AfvUXT
24MARS3nwzjaNw/ZgeJgPROoCZKqlKDxG3MZclkiN5B84MLY6fXRfKDPI/tJuYOu
BrQOMFss7qxr5JQHjZTS7oV8DJqSZJ4FV9wEE+s8FysRtfQQ5F7BvxIJKZfr8SaV
X4DNq04Ank5u/xalL8vm5TmdWf4KOsUMiIONPkiOn3uT/wd+koQDQZp50Nyw7NZO
FtpU3ZmZGcVWv2Amt4JkIqZHC1+2W9lspw3gfvtxDhTKonq0shKkp478ZLLr0+6O
OpRn5KqLzrmK4U4qYNANesIry3j3LtyxnuKZCm0btsIOzpgt+xCwC6YctLxnkvYb
jINZDTJ9fu+/2y3E/F8E3ttE52A8haNrMXOG361lwoUOxIIO0HRx7lJZ6lNmuwbm
HDB6cMF8w7B08owWVV+1sH+5NmK6d1EQFnoIgy1p8IxqAAIw9lI9sZH+VcPyEdJn
6pKJTW5uVKJvVeZz4j0C1irSqbTXkUipv/nUFIxhN5oXHnigssWPw5GkiB7zak/b
76v0Nf50RmxrvINxn7wTALL3iMfcoWivN2QfaH8id8G7+TDzE8RxHZ7RGS33PNh/
O9VKQxBJkiUb/0LdQocb97sY3wS37vEZRl9gLimqTC3mM6oJxwzWe9liEcoFOIzh
e9f7n9CvYbzZ0+yZVTx6zj/rcvUa+fjNZEZBPMk30sNBGsgjD2U+Je4cdzWW3pgM
PjaADpB/av52O/XxDygxslbN8ksX+QLGA9jUGnUrel7Du8BXjWH07gFmfPNterkG
croIp0qxNa1coUW8ZwvaVhPXFXsuKScC5GgunqV608W2HTlWvFiFR9yAX21U2KaB
elAAFwm8YfTInOvOVGzQ2WaaqjdRSWeH4HmS7TGrODVxReotd1olg4/NJgGOhYim
BoBddrh1CAhpXtTKZmWms1WJ7bMSJVw81bxVmpfH5XRCWSuuw20/T9JAs6YUblvn
JbwAsOmA/7qF7pU3bGD14zy4rf8TGbeCeUdG95e8VsHLxZyYqGF+twUpHTx72otH
CIlkNL+O8ReMq9mHpH5/+1x5zdfjR21ikSYld3cglr1MXmt5+k5X1H9PHLgEZcm0
H962qlkm/cO4AxFDDi8Yn9Ls6BoNy3BkNIBaI/xT1eUXgYyYjisjXsWudKqwE8nU
9PKhAA8ER+vTAmcPZIqtoFWaoYBHKQAzgib9Ld05Gff/e0jEeg4vHkdY3GrA3+sv
kJA4YxjttX7Mt76SwR9lv6G4nLCoU+Ani2F/VO7amAC+YsP2L6rpFNSC5IpUuFi7
tsTOd75L9YBHe4qy91O8pG1akkAz8gAqj7JnhgXmwh3DfS7MERt94tku9twpdl27
5G4RsSRUCsaDl2aOlVKEDvKuRxx3phtaPb7dpucOeohUyxlor4LNJW1vdZj1qgi/
C5Aqdbf2G89hjufGTwIR/tcSL0cbk3arM1hmPLeMnBOUTu7UQgWIpq0Mt3yl6R80
MhGw/56mqZzt+Rs+yR4Z0LfvsuC5trlVNn9YqQbzs5pIGe9m1tqkx1jMv+RLLZqB
8c2Ppgp1st96e4V0zFNW46qAgRGD//LW0HhsrmpXf67rnE4kSSOCrwBw04LS1Ili
2SE43o4yiG6Mnmr4jj12upnYNOilDw6yBPs+claAK+iuXDmlE8sa1rGeRc0ronuh
vElvzfOQxTG6Gtjefu7T+s7+Lh3mGz1UWa6VqQQ1D6bXBVJnY2iFzs411EXPmAVx
MNLqtt4qNZeRco6uJi6LEHsqDaB5H60jyAkG8cEF30XdVn/igk3TOJjjBW2j8Y4R
10pCZCW0ayB+6jkHDDp+Y3YpHjVluzW8T0Ygvwa9V2ZBlVCvEd/Fg9gq2aHe9kVC
Bsq/K8M5A2pv42UXGsHXqSyFqVJTCDeRrPW6eJqB2m/08j2Qg5aQ9FwYRmCVSSb8
nBFKQ82xY9UL0ClIyA7e1E/iTrpuBg9i2IPPe8dggHpvGEfIkb+pO6x3dZyIUWL+
NX6wi91BJhDy8hinFt8HIop9nxqhR1nBYkPHxn+Wz9rBH//i1gKre5K5WFM7Lzol
2LImbgve8RyiDHtFxA2LvbKv5qcajhUN6btaA/Lu59NCBPAmzGp+F3I+fzvjOltA
3BF56hgy9jHhCG6i66Flz40FUk+FquFR4JG9BdTlcBht/FNMek20XP0stucU6Ze0
aOBHKwQuR2Lk9VZO/fT3CqYo3I2X5qOGQdnPBITrJHekIC0tEdHfCItq+q+vKtkZ
VYhmRNp3iVFEoF/wsIzvpx7lfC/lNqyOqN/RNeBblQ/ckb38gbhCZuQuvAChvefx
kbuGP9GGqfvlEgPeIuLkaD5Fzz7LzmXrCsInMdBghyeIKqVDqG0usXzL4Q1CLABD
1gmHvdmjBRbL6yxfh3ttVW4wGR75a4kzKehJILMY6UgHHJgLvXjJYmokomS8BWwS
h6M9G52JhI7x5IJ/TBK8UrBqI/tx6Xr42v7LBu/6Vtn7v1H0qMyV9lD9PjQzO83Z
G85+MM9BYW5W9Q/oUUM8PGvVr3sAWJbJq185Ry29C4BVovRhX0RP8xFxDG7bYzV+
9Zb66MHucG5JzxdeOzalbdtvx/Hf5/ylO+tmL/90f+uRKpSUEoMKwuDZ6QPfHUnN
suhpvDLEVhSdV/cDx/wngdAd7GU/fTqgEyDDrAFjEL7pdjDUoVmtFW2+QhF3b9eG
snbhAhugpikk71K4r2z8vmNaaBYNUsRp764C3uFxs3Fj7iGot6i37jInJm8sZH02
B3fblLd/89d3IBuIgMiS5qItlVWPmuGR+gglwkvssYqNkgQNfRZJsQHpPbI0J6w2
amBKOQ6NnTjwL5SI9W/Tz5NJQCo4G0PC9ZTX/WOrmuZYbtQCW2/kFU1K30fN6bPl
AhArqDpD9xeApNvNCjtI3RLUlbVOr2kPdaf7/LW7vaR/Ns9pFsb7K2/M9gNywLl/
p93wj6bWYBihEsqRdDg7QPg5Q4mFsTZpDuGPL4dlX0VPQU2+DeYEi50tj8BKQJnw
8OxRlkqxibXBZs2GrfhFvkMhzCV89ZdmL/AO4BjjO5WO7NurhFCRlgKALdp3n8H5
Qlpe/70b8J22wo1KNZR1W6rIaMlP0OYpBYWdY78oelp0845Dt6Q4i9BfxKd6c6wd
dGXECcXxQLfOHWvmzrF0Ou2l5060C1nF/jLHF98WRbeIG/wNp9T9rhYRvud2bL7s
w718uZ8MHwidSDrzrM8YXHQGDlGz9jnk5zqvfiMmexplpQSi3T0ryRiZlnsAD0H6
CJtdJJJhcGG3vVTn0zUPSCOYgUDBqMZY7CH63phZbsVODg2Q3kpdgHWgR0snFEM0
fAiI/tluA9Lr4Qs1rXIo+KFINDbw4YvCgk1tG20lO6LyaqZ1AwHA50qq0OvdcivE
n/RkHFWKrerDeH9Q9vKe7skU2wPhEiXxG/WTJJ4AOa1eaeLFzOFlP7oyAntuHXz5
UgkbfGUqUUxUT3e3YH14mGeUZAzdXGORngQ86iUSYg9VUuO8WVmXAyszZBnz3819
pz1FbghfwSnQdSy8FtT3Ad+U3nk4TJngvDY4z5S/9rfxldVln0uyabh+OYGhG9+L
r6gZoYUKul1dwhQAeBD4hzAqgPtm9cqo5nD5glQDFQ5D5pBHIfr8YN3hHbHpMYcm
M0QZU1SjA9x6R8XN2uUwXii6/eAaaerTUcB8SNxB/oiOL7uOeVaD21FDC1Otn65D
oVyuXXrOOWyxilV66N1UqiCljw9OqnEG7wVQ5EifHttzM9Tmwv2ag/koXgoBxcAP
/JDsy7R5k+8zeiXuh3w8OtVXGLSXfWRQp1LiUmQiJq8KIOg4MMjtv6BNYTDZccpW
n4wsGcrOqoMHOpxQl2WDi67IQPRra1/wR0rDoXDu28olAQNCufMkWoO+PEFBv8M+
4DISdTLJ528a3IwrC9ohL9BjoK5H1lzt52jk2sMzv6z4L8vOZrKUpOrRl4ZB7Jsi
ovzCRfdYLfWPSpJdsz/SKF5hPQnEqXl474Ek9kfZuzuNMcZSvlzqVcNBgjR9MjoL
DakB0rHajKIoRAQ7tQGg3/MASqtfIzlUpUH4ZM9S7qgHgLMND54q2kSzK/OhLrSu
Gzu30wwceWw7GuXKv+ywfkd9Q737OgFABE0du6O8PoNMJlPMLLIewdIeyxD9zbQH
HTYu3Yg5xc0v764LIwnrW0h02WR1fOhAdyoRg+n8p5taJkZ4Aa7uSL9gsme19e2J
MQ4QYrG0q5MQTfV1OxgqAPOS6F0hsOlTdzOmhXJSFx2crHoiiZkX2tzBTE8tk1XS
pF8zlsr8R+ssT1dgyUKLeYKv0eFCTDfbVtLy5MQVMJPNNaSJxHFKWefhb+rNCHfq
47nzfhFCSFDhFq1VJHX/3dEFRT5CFj9Q7LIgBzPbwfyYmzGfBdYI6PzdVTttPYTx
CGQ5Laf3H2IzfUDeYJOqJ0yf377PgzUXFqPKefCtIKSRcmOB+5vJj0iqPRd3zC/U
95MpUVOvVGb3B8igjmTD7LUnOAb7zuXzRZUp/kRDTR49uD9FKQwQiX1dWbFGkCub
hlpMH19vACxiYPh6J/mxzUvA/DlSeVgVPfg0oy/GmHN21Zb0QZmOk8bvHLGleliz
7YGokNWu/Skj42M8ViaIIbqsUFscvI86M8D9oi5Ijh1bMGZ4HLfh72m/RgBwn05C
+aAr2Mrn1GOCjVOqcA5sD87Z8n3YXpmOzWXa0CVYEVNw6K5fWevXUzvECtfAXtZy
zcnb7sCUv1+8iT3/UW5Ppn3zIdfZw7DyxaT/FlVY2ew89EX/gPG2kWDT/42cz+LW
q+UgPoSyt8aM13OwY3js4mkdmAVkDXVlLD6W5mnu6hwDo6kqTdd++sBWG6UGxQMH
mEqm/HpFmjT84cet2+JfP8u9elQLk/mvE+uzMA3pWO8NUS7G9CCoDF+qPiTGdUKb
6sD6w2j0n0oZptLQlhaQefehvF04Kxwj7ESGzDjPXm0+GYkyslBwXfeiPNCY0G3O
8zsEMVycpRKOXXgZm3UHNABQpOxBgdrEw1bLAAgdZXV3zDkrPld37ln1Ctr3C+BI
W/0/Op4PwVmy7MDSnq7La+hpJc/E4eslNkvmTtGJ5JVXJg8p/I/J2y81Ukwuj9pb
fB3sQaL3jAD0NPjv98IOJqzhI68gJY1XU3oAdFosZajQV/SwNkdwQPxgsm7tPU8w
NaRAwlWDdruse4MPWrWO+kLL26xxwlc5ZvJJqbgAHcsmwDlp9+81NZP5JJUEkyK9
J0RyGyXJPdJ4DaTcL6ytfqex/WUWumPW0rHikpyBuKs28hdsXnl/1GB7ewTIKrUr
Sfituwt9NGIIqoEME7uwbm9ODS5uESvUaiUaIhcy7dkzjngftmDSIIU7Fzvkdt41
YxRoPMZhWLfmgSBb30hD9QIO+ZFw8FsKI1m8m0n4jIq0JDP6Tx7DV5U4QVzqK76p
l6cD3BrQG/uMm4G15RKTR6pzethW78TM/07v5XL6V4uvcgDVyE6GecRDcWjLz5XN
1HrwUm3QiQL+RZQcDIrDj5eSGhetorZRrnL8bSVQbbiQ+IR5GqJinT6CPVnoEhpT
0oY4ckr/P6coivtxzp05oA2cuCDrc01sOoTVPjfzkV2zUMbTpes7R53EzF0N/LG7
lu6IJJMtLPLwvqQW02BwVPTT6N90fwo9AgXkq86q6MNBCBY/xrdc1W1adJhQNupF
mnIOUDUwYsvdfh2wkd1DPo3rKihpILB3Srsnb1l+jj29aYtuercBRYCERpLNffnv
TT/n5xG49y6qTV8jXlYFcVolM7/z41yqMc9DpP9Al55B6oqSRWAFx2H7q5vGADR+
5imvqItB6LAbsE0vIAd4fPbmrsEf3VIyFXsCSOM5WbywJl1BIN+Wd+5rqdvYKel2
GD6o76ATQSwrGHRdS0dOq8+5xULXcJLJSccnbJjsntZTygpnjIe1GhfT2hyCY1/w
wLMUYV7j8oyMs4nz3NzNise9JDsEIKMtLLZhoVqXVA6TtklumbIh9Kh8hvk+o6OS
r4/HwMC6svOVVbQzDxMoRoW5Hjkt7pJcE5Th6jGc9sqfR+gje/6rLWP0svWvxGuu
aMu7OjbNKnjP2hqpl/lTnzRCVUrGF5RhkmrATo964s0Q3PjRgmmVwkrUuk678dL8
g+FemKeW8uUhaXWJXIm+SbOHcvUIpXOK/Ua67A5oElPctz2OYNaqGNYwk58XefaZ
T33sVC8bMc7JH4pfJM1TbC1NodCv5qZBsPA1ABRRhfV2/ZBy82BPggDBpPq6ow2J
CrKmpihEwyxFp7FknEhA8/AFLH8RpqnAxPFHPer+siXmx2ExQ5hDaeF57ZCpBWzD
oeouRloubqu6qNN6WTnIaU9aXETMMqPcJ25gI5vUhmzPuwoUoWc+HiAhUPO8Ho9p
NHfqnALBr8/vBhAAOX0s+n79IaiZVLlS9jG1d39A4Fj5jtrZiDdcLr+yGTLLpKR4
+TAJR9zvOMYB2T+kcC3K2cn98l5moIiEtvJx0P10/DldL5R17gc1e3e0mfm5GmYG
WlgM6jIa8XdU1pqKVaJnsl0RcGmG7dOscB/y2gRUaB/t1Gczp2ZMj36f2YbIttr0
EO/b+Sw7XnRLKXSSdvLxcIfUnbYyARpWNINtoz2juGHsmb5SXrPa2PpGLbJUlNsc
kaO/r/iWeou3p9X3L2cvBP+HqJpcJ+4lk7JxgZao/S+EwDmBXNA8/sM/GneOJTTE
Lr2MmckSVgU2dUqJZwajd5C5LljnF5LxYc3VpdgAk/fbJjJDW2U0uV4ZUF7FzKZW
yPwfVQ+Bv8x6SsTv6HTiWJj2PViqVQmUMgzRoH2V84NcOAazrb9TMsGSJvEpVy0Q
crVSQadFPTBh/MIO36kIaR8W9xik//2DhmmisM/y4SbDThm5LS1Mit2ESQfybQoJ
uzt+jJiqiwsn2tmkGsMq3DsOBaMPtPYgo9drscfTujO92OcdivuAUsKfQKqJ0eXq
V4pkrwNKaGoBSStXt+/8GfBxLzdtDH0LidcLlBMTz5lRJBYt0013OFbkKMGiDHoU
FZ6lJBD7IChG0s9TGAnqDGZ0tVjp3G4JNjlAcqZ1DFEH3Cavr+BfXPlhCa0gvLXc
HWL4n+GmVWM5rqO8UUh9xx94C+XfO264Hsm27d3jXfVhL7zhVnHUr3NfpX+B/aqi
3Es2gdWAa2phoU17OAKC8dViF5BgpP8qvMeVvtZv/xGqWl2vwcrBqT9ZNtP2RoAP
+RlRNxsPDBMrA8wH84VAxthk7Bg8+0bOan5jPQx2/bjjI0orvJv/CvbnK0oI9Fch
rvLwiVrPijpbN6c9UMMsUTvbmYAJKT4iqvG2g6UBk4tX6D8W1MAmwAmjjWduGWLS
nIitK3zJvFdUB85qYKC9kqaINEDfDuHVvp+OXKnW7JaWjS/iOzBU/IiINB8t21R2
6ijMhpVrueul95gt3i+JyVqnLsY42WfcISdEJC4vv5PtAPef0Jn9Xq9rw5pfu7Q3
h2ztLoelTz8F+JMC11BL0KHWC7AD1MFxrVnC2HzxdAGzVdhKM3XharlVA1javDJ8
F9HL2a7dTEopyeOLGaVJDNucn1RS2ETS+auPWbRMf4yn1N02nPoBM6fXz6QoezPO
k2WlIoq9k1mC351Vshngfy/Loa1+fluj+cwNhiVMVAxrX+DWDIVVlYBJwXOdZ23L
7BUs+JfPAQJmAVMHblQmH+Opra67z1RT2GW2nsPgt7QSwTOp5+Ytpmvmww2Q2xVf
F2l5W8jRDqknOVxrE+Hm2CUxtYDoOva319LnN7EH46jLU27SXmzL1tvYoUnsTEl3
V04T3p/Nj7EXgBrY0reBMP8FIbvW//OR88dheKjQONMmCWf/aK1YK08jsOpGSm2i
Zhk4rpxm45gkGEEHYiceQ2p2xaaDNWhfYr9jCmh+UAKLsewa+GB2SsZnEzI14UzE
nVsl0hDTjktw5wFNPufoNL89fKxK84iz/mXGVbyN8F5uavO3MddqRGTQtZnhwnwd
7S5UIew4YI9axc9vsomodHnTDw/pQldAQEyFwNyV9tuJlSXK3hq0p4egDgw76rFt
k6XU4pbwsdFNzPypGW4aG0rA5AA2xyiuA4fpx2xhoPPj1RPL0uu0PKjDcqIWop3z
APHg3Si5PZAwx1Wy3xvNWvuLSG+uPjt154qrO9J++EEswWSESIVTUKvYn4EvqUhs
2ZSJoljVSdsXsY6GXJ1yGCeb+jJLDxWWVM41zTHG+sqoy9eao2uDLK3Ut3G5RBBA
IXgtneD+6qdp74NUJYP/L2qFgIV7ouMcW98dSpEYWhB88YrFEajnXLvXibbIy4/0
jv+/PguED9MuAFdOPtC9mn4PIQwsdVO+CcWmyT0qACKvfz4lJxAlIGIrg3xuGe8D
w7OWgp20JGh6GQ3klzd0IYjwlPhfMXDNztCtg/+g8x4hN473w3J3aOyCsd2YvHBn
8CoZuQg4ORUcN3vkZKO/+5m2/hELJRJLqRYXwipYoBZD3fLws9PdziIPEBLSQsAO
iIScKKrvFJUQF1NGAJh8m7VB57muLR0xOlKntvI/P53AaJBHw0tbri19/k/7EaM4
cabutHPlQo59ZY0YNz+CiqD8Cr54Nrjs1q2j5oARUk9E37PR+NJ070B1PcUVvDA+
LLmcYK5ILnoCGu8JUEDvEziSUzc7qIJhDPMjHmmR9LTP+ukxGU20g7kOlLbN+OhA
fI/6b1OOsNSDYMYliXm766ikkCt09F0s7iLES2S4aXEp/nRw2gwkJTzo5PZAn0Cv
tetTGwMwJjP3cOGrYuZP5zDaAlaW901xkvXi0d7AkkYQ47SltX63jOaryzsu++d0
AFHkDGml6sbKzyPO/xVrTX6r859/APMV2Om1JOYDiytTMxCrKx80YwVfldoTByvC
rdtJ4ZQyRiGnWgaaire3Y0L9o7kpf2NtSk/B6Iiz5FOq9LPCeCT/m3p4obUNHWP3
PdEbPmVEyWanm/wNXRsem0sy5JX0Cluya3zT7SjikBz0v0HUuQFef5BEOhZtw1c8
x/Na3g6J16SdywwDgXPN1K3DHcKRNrOa5I+MhP6BvBMtAF/4GaN4rte1i7Vgq662
CHG28MSX9JCsi1B/Tb1a0tBoVZDrO5PhZ6sm2vs6Qvt+kqws5x9Viu+DOUru0gAu
QCZx3ld9SAfKZbbQI5v5P0LzLhcsk/5tQ/y2N3U8qqCx/cggiuyir4X1PmZuWc7v
4xa85+zd6yP5TLuEi+6HntOAtoJf8SwlTB6Jwee65gZjlySgqWh6XZNZ4fWeZwwJ
EnwnpsPkOsryRd0/aYkaW21mNc72y9oLIH9lbxjT0d8OuR0pUPlfD2MFbStkwVvy
U4PLz3CnPE/Gkw5f4RRyhp+r6VIxZ7i7HPYyfhJc8inYbjkCgQB5+myyk83sVT78
X50/BsK2qLIJV0XuZByGSQfgJ1O4PQoUpsyDCCTFJYgh5t7ury/ePNoQk+JCFrGc
Qn6WAdklWFq5mq6Rp9siiY1LdIaw8sxdwCDdWXhQCKadp+7O9zrAxRoppsUsbCrL
x8P9WYn1Kv1NcjwiwC5wSzD5jWey5myirIi6TPMEc/pNlk4jjQLP0vsGVVgtKB9H
tvOp4Nb4x566Bg3Ixl2b3x0kgd+mUn8VpEdvKrtGEOU4n5izWAdfryzNYuruScMC
ObW4pQwxm4GxcdfyoewJnuKhwQWc/WC+LTVR3KX0+MMuYKHR8o1RsSVYkJhrDtGY
jvuXV/QWPQiXjurqMoBFaNAFLMHSbqL5vOZ7YJlQNu9H9cr6z+D1W9luNt8eSdg5
b2JhIJF2Lg/GDZhScZzElQedZA+Qm6W3F1V9kJBB9hjW8bvcd03vYPiP8+HMTRK4
aDjfTYOdE8aCdcb2/bB5hTxfaQ71jFNKHokuT+7tmElzsBmlCW+K27L9uCEVZXgi
J31kA0xuT/pRgjR1oATNb9NADc0QhXNAKpFdiX7dfI/HNKtXxCCWkHSxU+wFMC71
0iq58kTDPssgqu5orcToByY13iL9FSiCF1fK34GKOWnT9Kwos8xq/nZn/khsuxmn
8niYvgOjGK0W7yS51RVYaab2lacFXzzskuRCBw5fu9Q+oDXbaAQtiQxBdYw+ppDP
86n62emugTKtp/Cm09w9EatiIcWeX5l9KQ7KKTpDnQeZ2bmSTc9zmpe5g2Jh4SUe
I/OqJtNxs3pal5Nt8T//MVHcRuPQ4kfeYXcBPo4TMtvHkJt01j+6LL0JFaS0ddD1
2fS1Jq2ftIbYDpOKAzGGgdobtiRCGSxABaHFzEG6PowDeVA6//VR4cr9at0W9xIx
x9vwhH+CvlvParxc1ndxu5tpdlA12uIDZJk6xjAHhqqAKzUNTMuWnLP2jUDT94/1
BGj+55KNdMvRpd6fJGL/QQU4rFIsZrza6x95MjNHJKBAf391V7a4BXt/S4WIXj00
CmHVbTh/nkEHYABeANIx7azqjpl+5FxXZl6D5GVhCjH11QIYVkcrDIBfGwdVPscg
nVjEwo9S4QgEWlUM6boA3hqJN8GDkSKiiVLoPz+HRRrWofNYnJNBi91siKH9CNs+
nqHiqpERugfawuJ1K4cicbcPkzfhyfKTUrvmKjNmCFZLk2NyZNpuPBSLiUYlk3na
ATtNmcYZmHk/sz1q8i7DuawQFeV0g2xH6R2Yk8bZDe4xSsgdZQA4b4BRJKaWbPhw
eVfC2Ou6aUFr7DMb6AGeo+VEF9aF2VCCSRkHCjJnb1IF4VjNUmWNM1tVkMTOqjoS
InFh1OHvTevvMIUzZ3Zop/NJy9myJtduTGUYNnEX7VoJm5VQ5MVAq60ooGVDopQe
v2xY2urCJJcc2f3nI4tyQ9GDLTlc6nBaSUhPzVNdSkTYuzSIcE8Y/yBnBRHfovVK
334iU6qctTM5yFsTbYcXNasHHGJvEXCGEb0bHSWxOzRuvApmPtRBXjytYwIzmWWb
kj8T/ZyuD2Cjk6sifT5vlh9qOXE4bh8uSlnY2f+yUQqNPf/FERLVZWhkra1PJ5ZN
MQ8r4cZI5mCIA+bI82OqkWBXdeuGFHr/vHjhFWyKirywVlnfGyVOKf74Do6IBewe
3O1UTP/BRv0Wtc8hdORoME0paru33XpnaB0QwLQbiTl5n0wTtuiFXHRWt7OflWl8
i8MLqFR1dX7gI8aGgAPpAKEGfuElSL+eqR9HsI+J0O+rnvy5T0eKOi+ZargEdaj0
rrOpXra7VE9XB/ce+Ztf74k4TNul9+Ap9Qk0IOPdODNPXCvCkVl9vD8qIjgNzQHz
bBxz0AR1VzIvA6NHdUSz8tT9Vl39EnxnjjmqEZfcWAB9zeyaYO8uUZ9F93rG+lTK
h/iEc6nUdyh1FHJFGEP66Z/XGA3cq6mgllyPQde51al2EGe5f5WIFEfuZcb/yVua
xxj/lF7R2rpHwjERioS8JdnzAxzewEfg5PEGj2XmYCVy/5Y+tsFOMaSxYOWsGUn3
oGewj1k0zV9A8JlPz1mxYtRdkdczvLoZEi7sAAeaxsVdzM4/lr9EzXxkQeOVPM9Y
qPoMRhTnduzF0RyaqC+fuogdlHXt+MyjH4z2EBj8w0NFiTNcBmHDCjXewkOq6imQ
J23kKQYBPhuW9nvH8zPBEPy36p0O+ISX/vY9rwyiS4M6p4st62hV1jh+FkyB8dyo
GwnSqRt1WMwoKZ0AGdQQSCCyKKi6fPK0ZYfnChhkDH8y4SoSaVSqbUIeUJZHwBlE
6MHmim/DV/fMk2WrS6vdeUgp3Xq5MRGrBpU2v0RZAeMe/yWn7XAhE13JJP1Qp12q
Ec+flf8gdIDI3AiIWSbfzAT/SeLW7Nh7DLkxpmC8uzdFK7565Zhozc3vh4bMmdLo
n44oHHaxOy1/OYCmRjLtGlKu81k/RkU7ieW4nEORzHrwRLyPiPNZ7ZCGpkz7yE5L
XmfcSrOYu6KPd7WRr93XUAFjUTy/SI7lQirLzuBYRO3DK+w3r8aaCiz5AHdM34QD
70MtYVrUJXpfISWtCH1/2qdengE2jiNnhY8eCYiG26/qDH61w/s0payEt+Wlud7D
O1Ug3YQ73l6K8PBu4qlTbG+wfB90PjfFYUaf5g3UPmOpBSlFYY9wU+oRod3mtVdp
ABRh8dWWs3i+MmhBWbpynAfmNcSDZ9i+z9FFkQdKag1ZCrKooPyci6sxN4nkFQZ1
SZZaJbMcyfgGIMG8CXjUWPjaumtMIBjwIALUDC0KBbJexhFQ6aQfvzUD6LI/+rR3
Chv+wqgNbY80novJZxtsUi7/tiL6ygX7BuRXoi4cKLwXXedsP+YABr0XEvARVYC5
tiP66Mz7uA8EImAQblhJbcoZq7hKPlOyVJWl94FfdEMwV6UbEpVQzeAv/JNly53N
8wOzDwLbcomv4oG8znsDBg4fSzJDutJ8HELvcxKzxRT3Op5+wuRqLnkPfF8zw/Lm
4th2fet7+3RhnLftVAZaZMJH3BBPpKJ/M0069aPrxJpG7F40KKL5VFpGB4b/m4CX
lXBJ321GGrWn6h91LFrQWLDSkAx0shdsOoQy38RieB4Lxcst/K1bXBpS5Ky6COf/
3jAtArDfBrfFDROpADXskhI0uCZKQ4a7ys/hCRxDYqjU8T/c5+21/+ISfhavYx0D
pNDl5X/nM/rltwdjweIrjSWaAf8cE9VFGbJR2QazUwFtYqz97otBhe2/X2mrLY30
/TMPfkI57lhTB/mFtAprO+hhmZJeN0BNFsMp7zWCzFWQJ9giZHLtZbKcXsPlbMV/
piRsL+gbqdM5bxtmSCIz8r1i6jQup619CoQSX7BNATLvlxVzvNru0OFq/g/xQ6kj
LxwIlB8GkSHY1Y+VRNpv/aOhV59EAs11b0g2gD3V9QhEozLKq6xIq45F809OPS0O
LpOuhAgwiqHcc/jWMGhGcQ/uCT6Y3zcy5DmaH+GWL4uxuRUY8sGumYhI0/aycITD
7f5FFw5aKlwDg4wRhUTGH5LeXt1l/ZNFP8gBd6LBT4ZVQ4OIdqlTy3UB9UvriAJC
rR0lzGSDjUHcZ5rtgYuCG45+yrWWC5mr/cPsaQ1fzqZS8UREpHLL6aiGG/n5/MVy
T9bLLtDk92UF0vqBxshf2B+MletgYylEEnuWnyGxcDbq52qiWnHhVCQi0BXHKHQn
evLkwlrLSk4XlZGFRLbq9iMiDc37jeR2oPC7hI+Ejvkq5IR2B/h4DAibAAXunppC
ajtOrIyTlFxDZcn1XG41tINVfX6ptTmkw5LMxykD4BT1Sf9Tzty8StS371nahjtq
eYZRxvFcrsrOUsypZMpnXsDbMUU6OuqTmos2MN/aVPA6Kf78mBKF2/KZIXQC9/5S
urR4rt97LGy2P+XxyFSRMch7oOi6Z3cCYskN8VoT+EXddeVzognr3rQzEjHXYZC+
fmJT1MYYGptIrTQwLMZodRVyRwG8MbYdZkh5cx7Abp8E3wmwTtvy2vTL4qVQqNeO
XQH6Y/4E1y7RDzbLWVgnnmUhE2Prc8cAPQOtvvFADsCMMBOhvxitHO6SBbSV0vzE
vY92BNQyA4jShZwN0XxTHiFhZ0OomR6sPPFRDTUheT3cCgKj/+lwPflNS2cJUZDU
S1jAK7vFtPt6vacSIudY9Czv8VNaQpOp1GyYYVzDxw3UeSqPS50T4VnQkytwr+rm
BG5Uy5XKzNeATp6uRc9nLX+JRbQVVhVCm3WRP9KkOS4ipH94WDMXrvYu0PcnR+7L
biXHsgvW6GkYPiUlZQc2HOeJYmUHEF5wjDWMmbReX6uN7U7EK8mlkDL8p/aUrDNw
ZgqSJHJHVQ9IqmbF7uIH0uw92TKvRXTHxnuWQ0SKJHOBdZOpbY/bh3oAurnryo/6
yRC3/0Uc02nwoQ8tNHL6dmEF74b0FMebQQ5coXVjNBfd2ZVmH6I+2ADJJ1uSxyYK
wYEUo07FUGK7eUoSp9MEaZB+VMJKKCjkOPOWM6i9ibBWIiNF11OigwPDzq7Jh2x+
fBhJMBPT8Tf5FzKICIcCT6viwW7dbuV4SwMCvHxHZPDw3FxHok52IzqHeB92f+1i
xIEexDye1hGy98CVkoMrCNlUnDHBBsS0NzAde+bBmU5p+cQh6tTAyqZfXbDC6nc8
gd08m/PwyFTYxESVavLbLEZ4K/UYeAKFPzVcWY8Mo0dK5Jfd5o/Msw/S5hQcXTup
WNyDJrlLLNQia+k1vye6pC3qllvMfHETXQOZrk4GV5obpXLxqwL063VzC+oKGhdq
xPbxuPaDjqLcu4+MoXEAIU2EkgPEIBTmH+9HEQES7W+3r+r3/HzyH2Ybof0uZ79p
UeLAM9INt3zZM62bCy+bgpZdjsh49PAp8x4/4AHYKjs6+MGuzQfCLSmVr2W4upbm
OcJRVI64RpZl+dQSO5iA/LnoO3SHLoRwNORylCwrxrpA03FiiNKmNOH2k/tfD3eh
wP6NqKuzzQHAI5WRY3UMzrOpRpV4MsNMC4wMp8JcRBNlzXGtFbdGB2KVNd8gehdO
pH6qhHNam/DcMyOjIlryN7JrZJErDUhwcqaWrIqORyWeVa2sb6TiprJrxlU1bpIx
aSSQTxjGXwi6fvpUlvSVW/NfJbbPLB3RfgyCS9oAFvElCOTu7UG50991zVULbwjz
YzuZ0L/bZS0c6qt2/jMEHvoZnE1m2HV3S9651vksXdx1GPkr8xQdkQuMRpz5ZeUQ
8hpNvz41vxL7o+IhyTKr5Uxwih3Vujen4oPoNR8vtlx15mMPkz1/GQ4vQtjnIJMV
RGi/TrCflauUqHJJZaHxE1uUBbm2UqLcuj+GMx6sfaDGJGffaLOpr8BmhgVs5e1R
TqDySIpV0NwIbzOyLRp1W6ieyrpeGjJsQgXrODDlkIn+LSKlUMz6EQf9DAJppO4Z
yulOO6fkclJAKi2rdM+Z7o4Sgm8BNCyaeL7KYKeH6lcxLXQonShoZKPgnjDoe8ok
lbM8mjqWI9OwivinF+jmFKnblDAZ0KJiafzaIQxrI11qog37vAqcPl5IBZ+GTwhI
+f+iMsNl0iY69lXjfbhDsJ9JjhEH2/63ofkqs2Oyu6WIN9pzV5gOzyiGqe0mrZrT
Hv4iVE7hiU84CJS1xqa6fbqyIUScWwzNA2TXZ4cxIW+RSk8tGVrMehZVDjYgc2hq
g4iVdZAa9xnBxhV2BbBVpNTmnkBvs37dwbva+L5xhGaJd1o0TPlqoS8wYIy9JVhd
S82GSWlEbq3A4XI8oJlQADdx1VPMjcKgrr6UG2K4dS/zozeLezS49W9c6+k8hiQ3
n5c6RPjXLFilmsl5SmpySgyfYgkb4ZXmFmK6ghXXgfMMChV1zRHo3KRHBr01/2oj
+CQdeymB/PB8JZY9ybN/f09PtnClHKO+3ldDTCDE/uYAFAZW5cZVgAU6vJYkdmoV
APM13ZmAUo387HfbxB3nqUNXtY68k2zOSBE1psrbGymDr9fqhZy3ME9aFbr6exD3
YVFzFje3/G5WtV5MurE8wJ0fJMaTnPW745I3ynEBhEPBh+z1QZhchTaHgRaP5y2R
RupE/+TOSUf1R5YolscEknYtysGu+cJ7ea7lhc8rW04h16pvA7snKtiKHI5S8kIV
5QR2fXKfQ7W+yRTN6PCDBKZRLEamHq5RL6A7Nac+JniLj6v9snnt3WNNwX5eoJv6
E7pQzy+1sgWFq4lhZqlyEtnJy46fBIkHulPK8cukX9T/0Blq/O1ZF+fit7ULJ5X6
9bqcjxtOfn3hajmNVAh6SSE56aMwZKSgG/BSKt71ZwzkOE4xFnm21K4vwK4fSxuI
Q+gASoxDBMW/hrRK88aGEqepEKol0kAis4tuMow/y7qinRsRIaQJpotwrPj7p1lX
f6HvXKBcq/lcWw3MeDa3gVtV/KqcxIDitym8AurdkQZnNiYx6cDkuJaEUXsiDBTb
qfi1A1ehZFLktXvdFfeufTbzkKqtmNhcLALR0gTlspWjxdVGqMIDDC+6eRWSmUkZ
5DPzvNyq3I0qLbnm2vXCvVcl0nV7vEOxan9nWEEUZe3exV3fLnfwGqW31MHwXliG
4ADy9eUWeB/vNuQKyi9kxshK0TK/F1y8VFfr7H/BJrD5nQNfpYsa6a14hfKtPaZP
DLk0KkMNUK2hgTK4wk/ERseao9JEMiPbEkLm0MN5yshD7/bHHej64bpj7ktYRvXB
DQEL/pV1MhzT9ZLAc1jMHufKq4TB8Pz2HDP7mp0IOjq4oWnPK/feJMuXQ84wfJ4G
xGuphDkyunGcn0vd25m2f/YI64N+YfrtFk4WVcV+nRYOGB+1WM6iTgKZTvoKrYK/
HdekzpvC5DCWDoI2oTibWDa/rPwpgqi1NuZ2CzkCcRBxW1dpNBKT9A4EiGRBuudz
RkxFm7yRJpysYWpAew5um9iQzZ9ki45lBcyqJwnX3q2KRSpv3YmCnKLBacEr6NSb
usnXZafoCaKdNbHFzgMa5cGpWfuAIdCWx98T4r3dBG9DxEBvLVOl4iP7hjqeY10H
oqplclKf2elHsF/fs4+8EfwvKtT+sEzfdbJa46vGGUj3V99rVwoCLcDwIXp0drox
d2v/hB9pJeFcLbZIz1MJLY10n1VBsDLHs/qzqiGvBEDU0TrjcXZdcIdOiayO9CrO
xWykNuN98vhB0dHsWhAHShbE0VXzYUE8dyi7SbSBSx3oqT1UD5egAN/aooiZaGW+
uRbsiMRQL+aLeGX9Dqm1+f9x5mxP0nFf0zlSXbs0v9ZUfB162qNMZDh5RQN2Fcpk
9mewTskvZwvAuahmYt/cGGZD5Tftxo/VugyvB16NaKSVcUbf3I8hylahMQ+PnUYd
9Nc52jl0imqDxa5Yu2xKCHKZziDFs3Yg+xEMlJ2t0PM577d+yYrPN/3bQnkFdSBr
L84plz/EXB5ifbR1slSIYA1Us3QW4fxtPdRKh7neeXG5GBKaW68vCHuu6oZ2JHKs
RQlC5eqJfvmiQxzmDMo2y50tK7XzhJXHGS/PLe/4O9yhepbb0pbt1oVF0LaKBoHv
PUatmv2Duth66iYHzW7g+G/anYaQFXqBJpMl7vaBK7493b/7hPiLQPZ6G+A6Fyle
Brzhpa/LYiaXI7vG0G8bYaP5bdHHK5xGoaaQkt1l+KoX+UBAr7EXWUbe0VHTg4L3
Moy8yc5YRDilLu6LeDa/Rb10ZrbegVVXX87mkXzEd40Fs5EZ6kEY2KkhF6K9e8SZ
6zF44lIGZ4+liMB89A2uOwZEtf0CWEbFIRAMh/NlHdc7gen3n6pSelmC9VwTm6xH
5ahr6NpRYx2JZ4JJh15Mfna0vn8dlgNCQg3s98nSAW5kaBzY1OlMOk2mXrwnn827
qOYbjGRV6ui9ynODwbP5FMasnzfrsXbH9zsG5onrMlh1x5OsE57fAfj7hMsSEAEI
6ifN3q4PP8dhn49MynFxatQhD8POnB93X8JqY5+kVdRe46/CCABvxRRTKojezm2c
FNa3AYoe3Lj+r/PJoU13LDPcYm37eeYYBPPBBx4NT+Oe8tV8g0DtuQHI/dujB2W2
LyaO4AVzF68a3/Ra+hLgLwYQtn39HqnRu7ApXuaw2kwabVU7eIQo8ByEbHAc+ahw
KNdNW5NlIHkfmEL3gWzTdg1q1XBD7yl3lR8XCQ+J76EParAhZDne26kEhBmzDv4p
nTqc5wtywlpNpVBRA4fBsl1J1WQ1JsKgiU8DcFf9CglSCmKLU4M/+mBXiH0dYiUS
yj0ngXgHcbdNA6a37l6k9hDbCpfHnee+Go/WwzdRj9WXTIh1ilQtB8RxE22UWQti
T6LvkA2lJtPOUmOHktHmOyb84+rRrFhou29Nz7CZUVBSsO4asfU94XcTVGBGbcnb
I53dlH7AKheVwnoOowQ8mivqg/UtfsN4qFkoSh3hhSzKA5PfP5iTxoYt69OPNs/q
p1yrCXDAT4Umhpi7gy/Y2BZmqN/8hFIgVwnVDvfZWpnGKcZbNy3Qg+WoxCGUdbP/
RZGsb5QiOUecSiC/3CLlXB3LVe1rfuHwiybE0RjA2w5V/OwiOqfHSW0N5LtoNsby
wBDJLx0lDb4aYzNJc0oS0PU/wDHmMbwRwjpAbx4vU2KDqAXyP2M1O4uIdD/Y8+Wv
ZmVaE03/Fegni073leeqx4WjnQkcMYnIJm0reDhHitFqmGcxU1jDYRnX4CFmKceu
gVI2Z/yuu7id0RettQtPowSzwK1Ph3py8wQoi2mJO85XQOnWEOvocBsz2leEjidr
w3Lf0keaME8uViNQ29EBpdLrLd+w9MK8oe4PQm+OC9HjIgbrEpC9yGjfasJLGuMS
p9V1vw4LLGlrYK4Xkcxs6LA4xgNWPt3s8vJ7yRTPqMkwCrX/v28oLGxgFzx70q63
P+2TW9+YMwDlFx0BCOAG/6aUnAYJXPZwXDsPulaYYBB8+H2FtorpiJU4i9gHwnSw
uz4Q2PjrtWM77ybpKt1EA5O/R/k7yG5Y/v7PcQLL8BmTwoXGcdnOC7Ak4nqa7pJt
Ert12TZmBP+2GgUVd1UaAS2wMn8VSSQl21Kkfip6X8s/vU+6TGMI1vv/ZuwYwLQ9
S8AOOwgVzvVTLTWwHoW7USEUKDbK5zuerwcbpFikQfKXSEeVnhaJ5X+9oiHRNOex
N5CX2NsyCTzBi+/gW/wtiy/LOepckEXdannUTt+oGASwS1INS3agbwyFGT5+JhO9
ReB5B7K32IEZ81Tr5XoyxlNEADGHgj4Yj29VgNnLr1e3HGB2u/DYdgXb30p3gdjw
cZRGtdvted7wfoD0G+Iz7F6JmAWJ8JDrnsSRKRTUWlfvOY94vZBdnwnSUWHYUQAC
TcbXbD4bxl7haVaFwwALPE6bUK6mri09a1fYQI4gN0c5JZPmYpoMnut8rZcnf3H4
xHQylrPcs/PQ1faB62oUDQmUD7g5aIYB6vpMRUDxnr1ZlVxeOrF1JSMNFYmM2rur
B+mGOk3fiXDRM80gAONiOFqZnwjLN5le3viM+y3TS+f9EEnHxli1fL6HJmCQj5lP
jrKnDJRK9IA6cjjr76ZTiUm/R2MiYFwDoAqlQa/nGqwLuC07ktzp8+dGQvXqDwkk
qaxoRftTr/xty2OCc6xH7hEx/F5FCjYVYA5V6jOy4bCpH4oNz5xFo2Wb5o74HaC8
BPmBb4Gac1k8qKr/huM3LM3uPjvCIyAB+ItH+Qns0cTpLj60E7P6cvNQTzG6DjQb
dClGKEuZXEWBWQYYZhp+dVef7wvAVF1I8miK9sbR03vqh/qenTSO48Me0C/u35dc
WUNL0KZ9puWcjac+WiWEq+1t/1i5NaVW9hnY+gQKYZ/nX34+ctXDJgHP+RIvqd8J
4Nbp4YOh/NIplpmij83RJv0/teG/V6kI0iBNvWLNmaEoe/uTeNpKIlTmKdkQeaIL
7pZldfi588MMu32BFd/1jlgOkCMRWAg5nXqugX6ln6zryaTPYHI3K4e/wjIbiGE1
KI7D14uiNQ6+HNMjsXcLnj/2fZ78fE3g57NPxOItF8k0K4WEmSLkkVkxviExdY0v
We2f8p7IjKiEhlacEkH3niAXp5Vcd7uIyRMRaQlgAwBnnzPOR6Qrb2fL/mWotxGn
1lHjc/Gfc+ReAC+EFzfNuaVVDJH4UUjhY9NjR4gAlcx8N9xByyea0IZUq5o31ZZW
+JCE3KGAj+IsNxYMu/jgapW0O6MOrOJitqbYTvcrdPqc6uVB8BlW79wi3AY4+XJf
DdWLYujSKao/3DKEKNEeT50Sv5WgYR3BCxppEPXEw0G+0KHo6Nuz3y9hcQQyB03d
PMcpOtw+Ftv7d9tUgnEq7gaP4JA65b/umi4K6LGEYv2NN2FOJKu2L6Y51tvqM07R
LFezOyQ+OwNSCoq/FjLEz6fDLh3hMBF8gc+wQoxXLumxyz6He1fY/YibeMm3dObF
75uXtRkZe0zUvtdp3fhn+b8OBMRuq2xatWXueBYz29X9jCrQI35drCfRw3u/N0r8
GdugHL8R3IHe+oueGrF2XNJ86LyalNCqarLueF4qF3yppYqzG56GGgqb9B0+Qa20
God3Ozkesbj4uTPwdhq3sDi8BYKa9egR+hT3pOykFHNQBUmNYOhwbr+ObPG1rcnE
QfCbwk3tPCfIS9OOvRenxpyh+aMlw82KmnGoFrd/SXsyMMiEdFub9QxokloP9ZKl
JXCPNuNlA+o4xxCRyjIiJMPCHVPfbn+qrgowspap1YLZJYQ86LoiVPfffZAqJk9V
5rb0VHEK5P+4TNkI4iWgy0sz2GDTVjUMgrsl6oOE2Rx5ku9jOC4RGm9kV81bE3W/
mtWnQfi9uSo4nFAa9nyh+4HJ0ntbqJT9d3A/VvMxHWkUi9URyoPF8OGK6QU/afmx
gk+oUJqqJbDQRJw8NMKVPmm+24MiZrd904VcXddjDFKwjM48KzDjviuKfxyMsx0a
kzbOLcNndAtGep3E+VZI9pMtzZboXTCzCAVjGxP7R3aXPgRVS7oKqKZX4MMJRKsZ
EyFlG3XsVdBq8l3TkTlsvXNIifOP1k2BvSEl7QEMqbZ0rcmQvrtOTu91vykW5FRP
YK9AwldpHkMnYby/5ZE0Eq5lJZuCFDtKk7jnMMOQ0/bPrjBzk12joSUb7UbYSUOr
5nLlmwbU1hj1GzJTk6bUwOrvgcgONB3BbtR5xWJb2eU3HIAX1l2HjwMj0LBck70u
zP9DN3Tgt8Gu3VRalhnyya9mNJgGZLIvqVdiV6IAmEjWjZJ20f6D/RqRejQxxGAa
lLfXvbK3x6ntH+QwuGpv4fv1ROrxNy6e+42UPyxHGOSUfPk2gEXIPnjy9YwZkjSc
fWtj5SjggPYDfMRfML4yu0+eWuKEJgJ/vfuN9j9qXREp1ivO7k3tOgqsfPHUbYQO
SzGwRYBZnWZrIrwH09n8EH/OTlbo6AlwmTADneVJiyL0v732pWNkf6Og7LFfWa2o
xDMpNXvAg3Ec+gfHsBYmfxtU9x1E67OGza7P+sciOseRbO+EPqLIxEzlDpQkSPZT
RwGvJdHrLT601L7Jlvd3bJcqh1qm9UIvwHwG9xgIc27ydUZ3V25ZSALiGNJYKwNF
nVd76TiBmwd8Kk7qXN3AxV508bOA/+oRtUjx1qAzFd3A7vEalfVw1Q1rhsVdXYsa
y0k1azBQjQ5XHZ5Zdb29EfdZnbm4tP+wKWOCNMacqQihQqgzXlgOxUq9ABzJzOZn
sIZ0j9lTkYohX2FkXu2dX7NjytvX2gzfaXx+qptmbbricecOfnq2DdeadiLgbKLT
EYTLjtiuWllcw5STdyehwGnyo0SBwLngkkO5Pz6aD/CTvWHSzHffz5/72csmWWYN
bHwgJKAUbelQk6sOQJXDOABNOSsWOB/g7+cOGCcn9BjvZkl5ePl2321Pqh/OYHql
1HKHE7qF+v278ZoIQB0l/ZAY4f6omPO4pkNSx/OylGN5r7QGeXO+jbhEIbTjTPuV
BmhzXn2lNhfRLjr7xEEFZ5S+YoRkIo4M3AKbijPxvOe4GLVgTSWaikEs1VgcZ0Bv
qZQeB65qEY68IBiatAb9E4DSata3tbeu2vAq1HX6BcyX1Lqds+mT4AJJFLBYCBeH
WcWERcs/VouZ9kmmA+sHw4H9nyJVhqlkqUWkMh9wYndCgUJ37o1Pt0aahPjZCvDP
JTagG4K93dLMTjh7RoEorvwD8weWyrFcNWIlzvHFKy8G6MF+Ks9moU/G36B7kx9u
h+sid6t+hN3CAGE9KbffvmCXcmSv5fWay8phuzQ8WaNh6hA8qnkVc6CzqvabINDc
jXcUHhjbU35aU8/jHoP5BEm9QMTGtCrmFt+u9F4/cTkKu7XMlGUJTjn8TCMiqRZ3
4rQissWkRGrndAdGAd0hoP68NgOx8XgnMgnw8wtAuW68XJ4anz/Pp/WRMOhIzR0M
RiOuAMO5qk1Y4LDZdYvTbyUlB0I9FJVn1U4o4Q5GVS4WPKmmSCKmpZR7bX/hfTur
irkyyBF8QF+XGJAgGFIzqnrrnYvoLI8BElELZk7/xEM7dJd2QTekdH49b/ubvWEc
FqfQOb/WGCaUVYgteBoyTSUW0jOcKdFjYKs0HimZhn5vONrWU1QtiyxJXJbf8Vgj
uDuzgYkNkccDEtZhxsz80XmxjwKcXtK0ndAESrNzjZvY7S7fUcld+TnjuxePOFX0
a2CJr7DowvnI2QUCq0HVtRcHOvONHK558iVzXX7R4yQOPfPxp7b5CM1eM5aFJQ/n
8nYp+w/MWNq9MXFoAgeq71L9Tjv7e5dquJHODFdc2D2C9Irk7FUVFTpAkOLcGKgw
ak2dQhRwSZGnqz44o2tcXrsoFvthpsuLFvWeCGBvFBy28Y0z/v/CrBHKlLlaRoPG
CscT3TCnUhrQ1RA/fWXlY8aquGlPKdBPSluHEykf+wF1dvrNYErb7O4rjn34oLib
YyrcCDjMnlxH07KHGfMBOBSzmvu2AxzG1F493o9Kv8BJCfezxLKMSnwNIhOEneE/
33PNoLkVCpQg7YKw/wCuqUn71Dajjlgv5mpC2SqFE0qO7p7QCidihodymSt1riIc
IiXDv02dDh7Xrgu4+Lp7k6v+1xtHl+aMUveW5OsSMoPnlLuY+OBnVns4uUbrce+R
/iN6k69eP6phoIFSwDEgis+ImS9TJvZ5kx3Tuk0pSyxmdcubcvBeNdp2IVeMHUiD
Cg8eQgz3QY08zyrxYLbuBPg5Aurx7QrQ2G+MmLKWp4x3qtoeroewnvAhMAqKwJlz
xkzvc9ro0CG5CZkS+ghXlWuvQRUNoA2T6VD3MhqjjCbQhtWdv273Sd3YmyAGyihc
VrfI8v8+0I6rso1DWrCFR8I/nsWK7OZwul7z5De9WtF0U0McyihyRaGJfdUM465X
6pNymcitl0qNke7Ebp65xD67d725qT70WzkGzwznWsZJRjMPUPrO3M0VN5iAxQXe
wW9fdwWm8PGIU7r/uJ7fMKSxOvMKO+U2TgXrzF6/ZC2Xe6ByuMt1gQaoMMec47Qx
aQPSw4lrkiHHfarzVS0GS1SMpx00+6OApWOAQlYJsckPM0lwJtQvq6g6H3Qj6Fvd
dB5XwydBGb6lLcNxpYJHABCkgkmEv1WZO2ZuNNSEMKyCUZKJfyZiJ7k6M0aIjxk0
T8Anle1n1TNCQJh21IgBIOFpmEFwdvCcmRWorr7ffJ71q1BRwx+yj/y+3bHdquCX
KcTIe4+JU2HDb26RqpOby6xqP/+O5Y0qxpEtVDOPKbk2mKzSVa06An0Mh1pRs5z6
KYcT/04XxxUY2q8fwplRWWPTLvzajkDx7WErrlV7frrEyKQuZ9+ZpLrbt+sK7hDu
ilc5OXA491W7TxG7UiT7/ne8tSzznyLo679IVkEb5SJ9RGo8JjVMCssDPf/e7Aib
e/4q1/9nRkLdcnbzPkEZ2WDqeaipVJvXe7kki6JfjyjcwGI4utVTUpqWH8AxGHGp
UXcyxEysp7FS3l4Frmyd77itvgvcmZC0dlHbCeJU5InHoGs2pWfyCAHkbDybK6Tk
EgPLTC9ARW8I9YhSJ0ZbaUsiMuAklQtv/a32AN3M0GcBS2MwBKwihv7NUE3MuPwz
ScKgg0+6ENaXgy+7Wd/k6GkegPpeolmRPn1r/HOfHoTWgBVQnyHrjIGjnu5hqLNN
2OsO8jrvCitrTE2RzHoZBRZQ+xI7+M/1TVWvz0btslQp1c6J66deo9+047xXmC92
WwjSeY64M0M03KTx0SXt3B5orUctO+e86cx4T9wQIdf5qVlTx6M6YniZhv8bimLD
SbHUBy1UldBGMgUngIYjyT5ntrMb9V5yBqYM8tY1FGFaqLmsl8J7NSAg+YjyXIr+
erotDlvr7XPeRHwIA8RmOXvaOczAisrXeCO6OLhRyKvxCsdmjeXbmJ+bcqDv/LuT
cOS/fUTgdywayQq+Jk9ZvPra2luHQ6BZXwTQJdjiYC38jJfL9EVm9GMUC7zXR67d
jzB36290Tt6doe9oWksXlsI8Fbigy+9otdaiiVHrCheLQaDHDeRaV+9WwVXMMZJL
HBBqmbyUnFVmAtDl3fL+gS7hstVbrLMGcydudFZs70irOkDs3IldjyDRdw5FsFRl
wnXrmQsO2OkcFLOGWnxfseOE9eaMJE4+/4AtWq12n67+j9zdNd/w7qGmACN7+Yek
wBzdguw7zaLbWKbKORcknpR8vG6JGvszJ2xJx8zIytP4r+JeCN5KVz58dJ0zD5Is
bYVcTK1uAjJ1393cHqkJCwZVmSlCwR2zhYkp5o5Ev7lzD1XtxKCqf12arbmDcfn0
4RVb/dd//GARoJxch9jdH9J+7AAjDj/n0D3nSNvz1B+xLaN+YrSunbFo/Jb0l4Mv
kkbz3V+sLNyd330DayD5P8OMzR9d500yeafNf/wVtmIgWFM+AhINmbFlxJrZe9zy
Epz9hteUgMLchDmqQwhF5iT9dJUMX9KsBS0CVgsWghL6s0ZE6TyhWDGNFcaMpiI3
eQIdf0ANa26ic930DJ1TTjXZDsEcQ9aBo4y1OFE9/RvcPa9BVqhT23T0tLppMxpv
oiDU5buRgnGGOpEDT+LreGj2kPMHTcnWKSkw/WMng7pBuK7US/qTzlpZSzzIm0yN
KLjseLtN+hk0wTPsUbzl+I4bTLS0Ku92BRJ//qTFDTNZQHIJy1P1XCO96OgWjZVW
PAD+xSKkNk8g5+hyAtKn6Nmdp13IaCht89Y9g5SI6Qb7keQMvQEWuqwYVs+O391G
aZPrqxcJo4HDHkNftyo5AzS2nrgp0GS7yUb/umQC/EkQ2sn4DyT64GOGIBOYfI38
+ZVSZcmvh6zvpoxOJ/5PkUVGoD2PrGtRrjPzZTQ1ANKBwbMI5BebMAVVmdsxKzOG
k4ueAH6LH0KD7E9ARgKX/Q8H6cJsMSPhXnfWexChLPrDdhXiWnGJf2AC+VF+uOe3
bhqL9bWXUQ5w4aXAB1fdkPm2v7zZS4Uisy1SUF4sAaND3K5B3arg8BO0d2CwQQ4T
Jq9IJE6YFHN9tM4ZD4lO8Ll/0ZiNwjQLE0mFz52mFeWICiH3FudfzFckPhgF12nE
rvrJv11/uFPbLyvuNppGoLLP4+GXGP//aZuvnCkMNXXvn3pBbOjG5ODG5MNTsjgT
TB99lusH47CQZSgmZtekxhvJOixBNrclL0IKucnv9lF8FTUbGH6TwW4o+JSS54GY
VwIyU0Z2M/HR+SqLNCo2IpTOR+gOoQQKJgd9BaEQVNLn6ktvvTOP4mGV4YHVtZH3
DAST42E5vx54OZryAg/C8WrI4wWksnvj12V5h87mx/n6jH/ZLanvHWbnG9fFqfoO
o3i+Am5Vo45BLoC2gsD2syXXgzUpKW9/kSWX2CGsqGrsqNsK3OtU4xGtfL+vw3Tv
AmqdpvCdURbAR0ByqZeuuvziRhMawiTHBECpyyvAFGS85SJcFcySFXTTaeZxgB5c
b/wrKseFT/YA3mtgs7n08OMnnqQmL3ZB9Iw5LruOkaaSjgoq+gXG+zAGDkuwLAc5
AeuqC+CydU5ViBAsi3nXISkAH7pqII24Blib+HLep4NHj321IoNy+kK8LFoTumbd
ZiD9fqKwoqwYsHJfoSJubp6J4/2ztlXyXYOzwou/WOVzpvI5Kbckx/P+GjHPyRax
ABqDnhQVPWczHBVXJ9fEs1A6nPWUoz0xQ5PnnQTU84Wk/vUv03EpH83dp48dlAf4
VWmYhzOAWzX8sZI8JI7fmO57nS//HHOp5zHhMPavrUtya/rWdPyGjHxSbJkut9/N
nGdvj7LlZZb4LoABWKAOwvoNAX45wgrqtog990b9V6TF2XE/PiUZZRK0mIkq/mda
2P8W7phU/i0vLf50XpYz0/YeVidO/SPubED+2a95gJJZ63H2OHnJVu+QA677g/ku
k7tSMAFVoeh3rudKlkmAK7QOq6QWnD0vOTutqQ1JQ+/nYDriajmP2dowjDFV6xR3
hbXKrtRvVOvaP0IAMWpp4jl7AKJrhSz+xTBY1b86BhA11yLBJj9epod2JXzN6HRo
/NbqXHOHD6sMnP847ZvYVJOuThlZR2ZR/f+ngaBsUpG1hvoYfTLs6kVNxpygV9v/
Ihj9BNoHjfuXz1JvmUyAV7XbK/QZm2shIF1kyNpPV3b00DN5LkSq6VTx1ctZtplW
UFGTfJLkUIMCRFTRedc/ZmFCDSpvlSpTrFtdkvMAz5/VLbTXI/E3UnDTSr7/e5tj
IuzZ9zUcdYiYU3ZDmGsrW02cNjtgDk/glx9nv3S7RdyXKTlFAeApqQjFIIi+2Lmd
XZ7QqmzTT5IGWRuZU4/2EyJo8NUXuOjMIPXhZ8HvJbs0Q6Jwq4wJc2KXEFhomWPb
+YfSG4sRFyCoZeF20SOKEd61ojMU4AVpt8qDzu//kvDwYyD67uqNWMT+owb9lHWV
QKVxkHj1k1ILjjkjrpV95vrk7dXIOEjLKDKx7HmykvMrjb0gF4giHgoKUG5qJp70
QFhASrNM73csl/70KBlNoQSVHRloQLXLpPGHImCPJJOs7c+Qh7h3keCHP1ANOkEr
G+3mYo/s+CS2UJ0on9A7HZYQ4nPz2Juh/afnsVX9mucGwAwKz6BD3ceEDAweZxd/
Ysm2dt1nDumK9HR9kPC5lzRFF7f5bWGsFX8qjOPjgqY4+yMweuBq15n3xQb26SiI
gCEmlJ0UXEAQY1YXFk73sxmGkZq39w75s5ykvHcQZIVjSK97yKWrlAtv3kSAaF8T
ocHcaeN5ODhF3wvvdopx/N+jteF3X6+D10AnNbl5uSDiPUDIvx5CJt2BRNVJh6/l
9duZCvUpHKJHbcBmbx/vsOJgBSy8CIeTkDnvvY7Jqn3qnGyG05GH32GSfgdLBI1o
ICQ/+RGVU1/7bLtuS4WqeCEF3p/nLSg6YabQsIzkUhAB/Mk12qhdv/FAiydxAtdS
z4gkLuDPNMpsH7j2sHafkXTgQi7ktrNgKQv4R8ow/sTh+F4nXbS0uRMZzip5XQy4
Du/4CW3GN2rXL8zwZ9/3ModTdFtAGrQ/34+6pWfzzAFN1blxkd8xFxNC5X3zSzbl
ilb/xO2NxHW/yeyOWQXNmaPd7sGjH1YixKhPqt9JMdS0L5SstAQS5C7+2JkqDuYa
3qG6bS212dC2KY/sHkMpKpes4KCvf+jnq+/Zf6E1wCKoEkX/tiY93u/SLUGNpCXQ
8N8pu3Fi0hdcEhOYmiVas2BEdWLMBQkii7afdXAmig332MnFuDf3MbhglOcBfOQt
5GgSmIt8O6vKKSQWq9si2TEiy3vjZxp2qD0TWrLguIbugbqy79VL6hWsF5B5gAIt
uM6a054vI/vbbHs7CnT+7P1qa1o5V1ucH+WP0VyNV8SWauGhBjEzBmOviXx5UZ2T
L03Q2qq9Jein6dL10xvd0xWCRHcqWdrV2umvA1FVJeNUvnyoYKF5WRbuKKWgdscy
v4h3AZP5E6YeqmwP2vk/0GVVM8yqBJNxCxY2hqHMnPj24eH4bopzR4wLPjyAJgcj
tGu2RJo7Z74XvAhgm6A6erm4T3Wamagoc/2lxtAJcnMM0rH/hdD0+I8LxzXgYB6T
czrUDsFVQ6hvhZ1vTuI/p6Ndscpok9Ij0Wh6z0t/dkGURjvI0kx1ZniqJo640Pge
G+Voag1JpoBXJXqfnZ5DpGINCu+IYoY7jmVVFRGMffhu30VmsJjKEWsC4nXYyJFl
QXBhFgiJRfjJrfsFdtoYIdGmX5oSy12ALWR94kYqm/q1h3tQhozMF/bRNur96F8P
6NnXAfnSUBiNiqHcFAsq4Xsh6xCB/KqJcnLSwRKE+hdQ6nLVGOCcoihLRPDyHf4k
Qwe1eYOpSokmYSgKBx+U4zQmlv/sH80OdFmmKewyZXGp0FQ/DfcTk5EErC+ufAlk
ioo+vXVibusC1tD8AkMzcxlNj7UGWJZIxrHDk0IIVck8rE3WcBvY3EHx2sK0KB6D
5dECA/gYqog7cVp6KGeelIbYcOK1/LPTfRugNWWwZf2+YgWi697mMv3Iw3th1wwH
RE1cMnfV94oa8arFUM+rAis98bgFosWYW5RE6sT6uzyBKCMw8T+mkLYqkit5rdTT
uoVb5NrE+026yckowQ+Qw5GB0HwjoP0C9Jn6rpQ1j3FMCYzSVaH3dxEbYBe2E8R1
FYhtx7O7oLXieLIeJiMmoZwjrf01VBcCXG8FKHfD/t5kwaJtuOj3/+sTjsILvqwe
+Zf94QhYD2dynPUUvVv3/APkH++Q5xXsRv4Bxoxn6Sap8EpPi0sO7MTW4Uv9dmeP
yv5RnAjgns6oGB468cfnDUxqBpoF5x7mrlN3KosN2eubfRk6NK4WRxYhb29Gc3iI
amAlq9pTLmkz+ZMkqwh6twiPWL30ufBRt+7VqQPvOejpKO4SK/llikRTP0bJxhNU
LZo4xv+X4YVzWTHE++dueRIy+441nBEBbBInHSvZ/ScO4w/0X8b4Ev7Dz7JIL3oS
RsDsaS70qoP6JoSaFQy6rbdy4Jl9W/zXpx0tOA3IgeHFttAsL/qHxgRgY+V7T/v1
ld9PTn8YFaC6bqEfwBOvrva+TAJ6OexiSoLhA57zcXnrM/Vtu/B1t94TZ8NvvLMb
j3d0bvMfjCNgdf0M/SJ+WM5Ku18huhXyAPWR1ZyYNX0ZKgV9cTpwp55Lw/bAlbvh
xehtWJpsPj+3r6/x40uQhnVK2AQYULojFYAG59WgxtNrZDqTNDgzkF8AHhHlcUlY
v9VZ38M25GS+sd4Aou5BgSoST9eBDUSd0fEjnUfn+jedZkB4pJeJifj7tkdgIRKN
3peS1tv+fvKBlncYNhTdT/kA3sk9/SkbfzIaprxUBOcssSEf5TSLQ2O/lre7zt/4
N1dRAzhVPIQrjuIrR147XBf9S7jesN0L5H1AmYISUeD5sBnVNCEcRgjmtu50Vy9u
km/b0OrfVML8sjZCyDQ0STLjXYeD+M5VGrYfbMVhpUELGevNZmsO6k0DnKDzApkx
0bfRXekeaPjj68cO3g9mrPtY9xB7aRQXN+ZlmfMjAa51JPGtHhR4UVMjBZ7S3ovr
N9bgAMXbTdjd43RJF0U08bzzYWnG3020xpMu62EfUlwCINqNSz3CbTIN/VzkTyho
/ok3yjQ74SUtJIL0Za2ZpjdlDABaYpxzCINm7qVTCnk393Mp1cBxyIXX7x8ANDYk
bx58vf3XHr5rDbSoNV4Ag/vf9ZORLRUJumvGuXtitCzq1BbeQKbHgKsobVtoMt2b
LTk8V/K1s1F8scBXxgVrMwJJr2Te5Hqpz1+24TTe5HXXEkLSzioC2wRzIcuoTq8S
XHk1iMVjKeJx9gaftMWWezTDavfvn6x3Pf+EZF+YrVMwMzVzxlU06JbI81/7Lwbg
VPRkDihsOWijTWuserpfbGx8TR25lMC8pHgKiNdRyt2zYgg0BZmrBROrAxsmopnp
pXFKDjYpBCS20VuNnHnEkQGLozxzKW/UVYbRxHop1ghSojJCkz0HFfBW87ZcZ6nG
sNshWZKGcwLEVocgZvAQzij9bBrt1s+17t4NmCX9jRWTYsPSBs2J3y7nqwqkAvvL
z9hxYnP+PQc2DIXeY4LU7RUyFdB4AcTgLzLDRN+Haxkv2dsAwTtQfegfPik6RUYR
wfe1cHjy0EvnrHDWv1nVsedkSyE042MuddzDqKri1I4LTT+ddVu5E0LEfuCdeSAB
duuCEOr+asDJvUqbgBMMBpBSl0TXjUVHI1hQmkUVxmZjgmQGdCsziGzV9eaCFVEo
94zRfR038iAh6xwxffcg+aLwzKFEodrDPJCFZpE5awaAWQdHqp8xCWDEcqti44dk
Bv3vdKIlPlI5sW7n1opPXMSw+tTDEGFXfWwBfU1Uv8eRJs44tTfj8tLMVd9+6y5o
DlMAFl5d9W3qhScnXb/qvBsmQhHCpirJ7lDZsDz7hphlDBqvVDlTENQYTT7/FcX7
r+ssVqLZEEQ+CqdAEoQ636iXdOUnzARNCqct7bMKHwz5M/ZwbajVhq757SE7R3RJ
8WXTflt9sg35vWuYk8a6kt/VJqrGZcJ/gTgFf5PzcVYRytFgaFKsKFZB1oQSv0/m
4LsiqHQZtDjrwgbEpS7BSEl5IOvWWigxAWSz0qC5PjII6d1byqEnirkm6ZI0S1iQ
kCHS9QEoZiv91Nw5MUaEPzBloaqPa02BWyPc4qFxDmLH4CsrGLjoUnHUbd4SKmZH
ZHgxYHcWG0JZE9rkuTLhbeBFwIb1gwAIxR1jvXqstVom+Prh5Gxld1qzrhfZJpUc
M6+U5KziZUZDDwqgihhVxF/U/tMsxsVJ6g38UJSpAGYxUiDE+uDgqTycxzixYYAs
8KuDMMER5NiBgErItACMMmcnX6ZLhTm5TMBtbHXMMfLgRpghCOpQvbIdSCHwuERE
nX//PqHhIVbOnS/fcWBqFYp1KlYgqyfP2utO7dg3EF2uR3uF9BzkNzSIkLpFaWC1
ZN+S3dIMjOjoelU9nD9YcLv56MD4pG2HVN6vocjHvfPh6sJ2OhKK+MBq/JxjSGmo
tYmTQnegyIV3c5tztyRTxPHj0m0GrTYGJQJjAotu6gJucc1S+LItI86IB0T+m2Gd
uSPnenRKfOB9O0xddWr/cG9AYmBMIRlCpnfTWI2F/esIrtga7n8v3ixVghsLXyi0
IAexBvPiCC0pBNB9UD0yIcjjtF47iMWB+B1V5mwGAiqarHiHdsjIDQvlHVueQe5s
u+UVLKvCMG147zRSopKyjPlQR7pRtv4vYMnOorcRswhuBC6zaDm3xOj1bi1qoLK6
df1+fRrWi6rV9AmjQEtPWfK2QRfiwiKHVMcz8DXLpx6GtwDQHeisJwZ3gzItyIzF
jhacs3tHemaxcfvJ5KFctvzxqMADjzizAUfr2VN6V6FFBxaT8CpdZ2DwqgEQUY2Y
HRIbUnY8+5iQIe++pxJB/wKe9wbeLyUSfaOpPQ4OpkfVitrixgK5ruhPZfKsVO6x
5daBxfsNypE2/zpZYRvl/BH8U2aYGBIyvuidHfDds4bYzfu3GRs4Lbis32ikTdoz
THSJSbObB4FMHg9Uz8yYEKd/pgLKZhGLrTIh0WxFLCIFkLUA4rw6i8hn3HQvzIhT
rYv9qu1o+v8NVeGVUbCK6zfLhnw9i4GnTEgiIXxnF4gpiDWgXS/z8bEsrTcVVLJx
77jJzC0KLS7RbXjUKUKwmf/6RuMZEBGRkpMwk8/R/67KdJg7c4jp0JSBrDWgTQFy
6PNGsQyuFZWC6V1YMa6lT19OgOYu00/4lPXtgUF2nVRPDEvJfeHHyPBZmZkUXUBl
XT2MjpdsLCT5ByS9c3YDYPFWVEw4WAw5WXeFCQIt4F55gnKOY5WPkRlDZiVxmNhU
7OHacSm86fA/PfY+RsVxETNGO/jtTXhpHQyFgWglSwmLCSq+olreA3dHeKVmjn3C
2CTtWRipw96dHENfdaV3Px/1AmxQdOoON+IL7J7cM0JxVfokMaZqTx+q1beIWvC0
HBrrFdLMqpKmpRb0N3v27It03wpQd0bujxsD+pDTpxiSN3bq+dl4HVlyLx93+IJq
QUoXe6R7LqDOR1IVwVLHldOfnkhLCoNCciygdIJ4Fb33dIQt9+bWEZieLhcRXYUt
9tVCxB1OrIPHkjes9sswPkUPdHS4CCsy/BL7dZvVsTZZh9xn0AJ8Pl7QeOiBBgw2
OW2znS03hkmV4wQLWbbSWVrJ2aq2FTT3haJiGPpvVwrrr3JrnGR2pwN883PvAnWB
JfnJfU+fHMDGW8lgOB3/xUVZDq3rCB7SNkmhkl0QShQHeSGHntasUxxg8oXF3tbR
u+WIUnKIgIzuMwDA741Oo0Llto0bdHF2jCoRkZ0WbSjrKF18lPNoGjS0Fp+nbuN1
nI2DR+MUEai/1dL9xTA9+uF6SM4ZJd8D1TFgwg61r3VfDnZRRH42pD6EY6KTEcDr
1sOIlJ54EGKO49uACPT5bweXJyJjwJgle+t9CpYRogzT6AoD31owXzb11BK0CcK7
eCFzQPUT73gIekf8Mrl3gPSqyY0Glw6fTLPthcpmvqPjW6O8BRtaMrrFxXh0I9Cf
QC1d9K2Ydb551hyiJLp8NnGZtLktd86Zkdc2fFn4/JwL1Tzq7RggUH5sgILIOnKl
yDHHIeIGjCloBLRGp5tosJ52XKBQalr0IYxXRg9u6hSnzMTbCmsyK31lQdcoD6PD
6kb/0ZFz8lsqIcna5173V0uVtNLjN/UnMKhvNb4o4BEXMD6c1bsxgMFkQi4YiKh0
bDNqMjRnpNCkyk3Epogq5aBSFhdCRHggO2OQAH3jwvVQzUybaS5RFJok3f4mV2CZ
mWLdAkl6rJ43UXlfMZV0bauT0AaCfMcaa/5cXxPOK+lD+1PfuoBiVQZ9QX9IAKqr
83keMdPIMPZoh9WjeyTpz8BYep0du/LshdjQrGBGZMrEdoxYLETW/4ScqtqfJt+n
bFtyJzVh/4N9NJmcZWBaNlCK4px0iy/cxnfWdanEInITMuI+0svJv4BJ6nz/mgy1
rTFFQmN01faJbj1joAz8UQS6p3k6DHxXj/kvOJ0LPAuPPE6SgJDQbpvhFVZL5tru
9Zo8KmB/y7l0ESefSfhjwEurYYjES+WlERy81SinFLOfiX8ejrWjVFhRMHMdSz0p
TUDkB3f2hEfHyqPFG5ElCyi084uGQw37YIGfidQSQutHZjMLeDSlftjgrJRPwFtT
p0BaW99dPdCVnCpi56vvehFDAfxEm1c/Uxx0VZjT4wQOPyovEE/mdgDWHt3M/WDc
qnTrjT+cAupk7ZnV4VaLQl47WUY74MRp4DHPwiqbvhyVAlGXO9t8BIxm31KbtLuQ
hMSKmpQG3WGcFYlEO3oCVtHS9M4kiOOxihmjS/Aj5uX23abmXwrqu7ZLnnslfHV2
tjJKlZV1XTvPkSlda6QiqQ5IzP9FWpNm+MPm6PX4FQfB7Pl302Dj/syE2zdrUXHe
iot9BnQBhqgFXJDTTHYKFDdtt3fSb2ajBHU133eSc+mu3UWNv6d5hwXEWdBvT+NF
99+/+38BD3KtDLsHiDge1u+nB9QYwhQITTBtx/NNhlgaD5yFXpegavwDAnh+H0Dc
Mi+9WUAr0aWEuFB9c+3EN+rALUod4LlXmxzzbr0fn71UmsdlhJ/jhDNJoU7DRQ4b
nI7u4wnuLbk/GcWI6jBkObuBpG0A2/YsWP45i0Jz+DRp0Qi8BGxD1eNsTyO+8y3F
jf+CsBqBExizzRiwKtTIVgmpBiGThPPuq3ZDwbGUIFHKocBhJy1meI9dMn+VTmdk
4ygdxbokumRgHP5NN63WOh8foJGIplJgkpJFa1djJ8WL4wIrl7H+8dibJUJPdh/z
xBhefqxxsEs4LJopFan2eerDlFjYjHeTszp29OEYZEJVljDDOEvwo6wLIPL5d9oX
wLzby5bjWVPv8M10D+SHT5NIVpUILmhQSc3RuzE7Vk2jP8CJAqv+ZBHzvDeYpBwv
V0Txx1QenV7mCMueaFPmBA4ROs+SlpN/j9DgmnIDFgD6wU4PQVkR/3fWcO6SI4LN
tFFXWOCDeMC8TFGjGI1HucZtLmEPTZ29Qm5VkUgXmwzaw3Lp1/ThQpUefwlR0Vrz
uvs9qa9Plmx6KgvxsVgxVGoltoU0AHrm4a4TABJhZLd9TyKxOSZZgAxFnher0xUX
sUDfEBahfzQcyGuyMO2pfNkFkpZ7VhwC00RInoamI+NyDvOEjXzrVFWKRmazwr/L
VBlGUBuzZ/oeyfk5dY9rvugNs6UD8uPHUDF0b/WuW4Ta0ooW9zxxVzAtku3YdajW
DTKzYmUVDPol/WQIn7xjl2kvYKEDHe5+dWqcDbPYPEJWyRXXBa1OLW9V/XanMZ9F
02Q2WJKWQgXZYoq8l8h4b4zgUhBHCROyneEWuG+HKO3wez0RFViVTHUbSLxws0Di
m/Fn2Hk+8jWXpjkRdMskwGAUTd9xlFrpkeg4xwpTnJe14zJww6B3kIt4iU2BDO9E
nm06NJHoikh1NLGCtZKW+lsUgA3YPpbfv0pY5rbByvu1XqlYUTyExysPEfsZ48j3
nPqTxp20tg7zI7bjfQ5HZJ3p3EpVB4X3pcqGnbYt70fCkZ7/b7uM++3BxkShFOvd
A+i3gx9Ok44RM/0TulDChsK1jJ1y01OctW0uTHzR46lCaPrRzNeS9c2avXwxUHkV
RDNTg7iJ1Y7XMbyaOYW02DKGMcUDzREtdxDN0kjxkIpnq4+A+KEaE4L/OdLqMGqU
maQsXyni4EoTFEMJctwa08zUtAQIZqGiU+aD8RK3b1aQ+aYyo8lwZQQ5sCQLM7uu
hLr9MKTX88b7WpWEDU+iDOo7CeMbxWLWz7wu1ck7h4nxj3s01lgR6kJqjmsQ2mlK
6DSwlv8Of3UejonhoYPy+Dy3hrcbXC5gVVU/QyfZgsxDwsiZ/O5mA17aWQpmRF69
KGm74jDMwaguEwd52hwoew7HosGIbl8ny+0AvtG5dvm5bwV8zdedqDrYsv79MLz2
DEbg+Igzpu0xBTShZmRWg9rt8MU4uE+lhsrVpNsBdBsS9FU3KkeVLbKVDxMU1NyU
WJIN6R6WmzXOdZtH3dTW8O8Nr7+9tAFZtnfy6TQnOpJCSLjxhWlZ0TzDuUkouBc4
XfNzqhXCjGYuAcDHxngnbvS3MisbnGxmIn67+NqZaqWNxZ+SfynpQruaCP6eMFfl
YKbvPD9OhJw7RbixDGzh5QhOt8mvca252SkHK5RZ6nXBEP9ggbyYRGmFhYzvwO+O
A6c1BZMgIfPTGPqR1vnl0wGJxF4RM4CGTGP2CKmqauHUVhh9RxiHDYAbA4P/doq4
LgKiDhjHDE8KR58Fux348r/j63aYnt0Xm9Dxga5sMjNt8xq7yawKkKB0p5GUEeBg
Sl1PX5f00VRgyosqPHTt5IuTu65YoqqoQfID87ub0SZoKcuO4GHzFvYRwF85QxVi
2IfKDU1VXqdsQaHqu0TvbwHtbPT/irfAAriDwPlt27Uz4xx+gKB1NCwrBuQnb+w8
uh18qQM5E3gh215SLl+GG36Z1kF1dAY3HU2mz4BCy0oNwt8aIINEvrvdP1tV1ptu
ZjbFVzNvgEui0OwbpFbhGfG94ORIIWVhDNsaFCsSuJkSXYuucaTr1rapTt4fBl/L
Q3wGsdosYebkzKQJhRAJxeoP6oX3G9+Up3QGOSZpI6BMpVRAy3qg2YveEOlFh5wA
qfReZLYjrZ+QaNPyKcVtitc+UiivesXIvwTzJ1K7ydq5bw8LMOuPB/bHTpk3s6+K
gr2R35pobugYDr1uTF79kAZV6p2tPOq4MXmennusf4OHuoHukUegZB5TLuh2R80f
k8QMclBgYKQcJF+VXFmaH51upTVlghIsmLczzdGFYLew39TUyXAu1itLc/ZVpxNf
nzxRHg51kAMAXH6sSBWiSE1LCFHvMGIhOrUPyF6nXUaehZFiVvmZ/v3Ruzqb8F/O
FXISAu3gpUabwAtjbg+JKNjl315XcCSSLs+4GmVj2PXSI5sy7yh19lL7fp5jJoco
FFEangZIKj2SZC92KCwpNcE5G+WXwOAVim0HC+1PXp+5P1juR3xMkcRXMNVeBa+s
6xGzJ1WyY2w8pf7+2QF1dwOb1DKewTaXhPQDQCPLFYy8wAq4ey94njaB2wQs6Ga7
4UvffljEqfNJ0Vo07IxMXTg9UQIubWH/1gE05PEKRlzCiEp35pyGooqLRc8fyMGG
Qcp4t0Rkzgt+3o5kSpPovQrCURxcLjfmHBAiA0z/x/8CIOw/2XX3LBSFhD3RZzqO
9zd62z863D2Wd/V/uTUtN39urLThjGcMW2+6V2uz0b2c+9Z77jPpjPLDns7Db5E1
UbpOOw/6sWjXNdm1RXX83hsYeaNnHyz1mVuavexG4KpJrhmUXYHNRGM+MJvXaOaj
1TAFG9gabKiMsewfgJkXMCyYDEeyNFjVFysAZ/uT3TKUvU5e5y/Sbj8tgYvZ3asA
DpgdYet++b4RzvlEruwoZ34JP+gafJlDZzO3yoRttqLNji4uscbnHGshev72utn1
puu7URjSkrRy1momssg15GO/YaYowbSsWw+P8NX3JLnmDl3otVBbIm3FOWY8tWCA
V71CcboMOCiYbv7m4Gvoh7pZBqoK6gdTwMTvha9ubjqP83hxYjo0eeDArozAj2qg
L/mA9XDYNYrb08uxF5Iss6EVUWhM5HGQM9OYbLumhX4tNf32FocIBDt9wSfmPg4I
MACgrJXncSGmsCPq7FSDe0ZzAf46I1pE91c3fpiL2Rdos/tzqLR+OBG/c6ffCCzi
kxAxFbUVavqIJAdahZ2KY/cOHfbEHm3yYONjkHb1OSRyfHurXB/nkgnsS9jnD7hF
RrYOV/J1lhqunwzI0YBJhEiGqS9arEHANU14GEkeiv61rirmRzchtxMznpMUQJR/
VcKcI3+FmGmZ0r/FvhF2idmN0cYnDJBhCJDJGOozFFDYlr7hX4ZJA7L6SEddr5E6
6R3zm3kQgJMzE2JFjVJo73qAOPTQbr4rmWHI0JLoTV5J3a2TLb3E3cuiM330+SnE
TWWc4fQTPAbCN5yBwTH1HMDLNIfBWpRGgQQCUVhMJQqaVXi98snE24PiZixWUHQy
MWEE31ntyoC4krftUvhX8H0s7NTthz9zyRNgS3hNYL2EXLt2Qe31dSc2vs/Vi8WB
A9+R+wLNeacNKu7H4+SHnISvwZRrsHJgR0Q76r2ituL+22tTOTb6jLMSO93e8rJH
HEqd9wnFeMbNAairciAldb0vJ8GqLwgKJOKtJeANc75kuGpbL/SJiohpWdfO5Z6R
I8kRfjYHckG68O+4Tk/P/rRefju93s0B7PCp+iyDuztgGYfPMZFuO6rBBjl+RcQM
c5l+ekxRUKgdQ5ymeIth1bLBUvB8lW17nuvxI3nvh+WVbVtWM5F9nt0wZ1U5U0kd
CTsAZ0/Vc37WQpBYCH/h4lpE3ekQ23cmkDrDnhmvIvAtPSp7c2zpFrH2gmINMrpQ
Va9bpd9BNzzwzNxqBNky3me/23L1IYLIT/zfvwMI70j481ZHgJSEKUbRZSvJ0uZB
1DCK4pgBdsaLznIyHh4pJN+LvJL9CPapMkPH5jbNb1/dfBisWM1lZSHGtXnoIHd/
KwV9blcG4qHgT+mgbDRJP/PL1tJ+AAbxOZyd6cCsaZjDtw7AakxHQB0D6BbUDhMn
gAbKyOU7yzxAAfH1MPa1JKGCWyXPtAg9490uiSHBUoFYeoaD6tdQOqgy708pIXEY
e/MV3dgDM+4yij2oyIUPUlO0bIYZk7jykOH7JRToXrSyLUqe/nI8wW0SSO5Scizl
khMnTcTeY8vlRQslLyUgxcFgSmJ5iYT0uyTcGLbqXoC1R27f7GeLBrSw5Tef6NY4
5n32thMWWHUWb5E/zu+PVrnGOEOQvw94+jgSYtX8/PVQqG1eFi3pwadmIXedB7ru
Kd3e0JznMPqHp0HyOuf+MUonerKT/rK9dpvTcwbIP/7nxHs21dm18d5IDqveQFdX
vsEk2nhs6nj7rZv5VBU2XSEIhPDMW/94tLLcrmjMtqrnegBUmfisBuyyTmKRm6r1
jlxLg3nqsyoSZaAmLp8//A2SiCeRGfWu2RdosZEVp9w2zpeuXolQk7lWMMd215Gl
TuDj4D1UHNZlcCT700i776RK0a7Nevu0qrbnQownYFrtD/RtBt4+MduMlhZzku6w
P1e25vn3JfTeuy3OQxhylHfo+9/jrP2VsXBQce3d0g4nMDFKfNj404uC6LqpVxLN
qPMn2bDxpsV8R4Pw51IHRdd3arYRUTFc/XCje7jQhtqf3nSdGTvMxJksNWxpdQvl
HDl7xVkIKIX3UWpTDQ+OBwnNgf9xnl/P+izAd2x+nVDkoWknYfI8sPs/OPS1OAiU
Vq8nPuwXIGZGpAPiOhBRq+Xt4jHupwSsMT+Cvb00cCIdjyEApQzDD7Gv5QD1OOWM
jpu8Y6U2iZaIvdwDqa0XIZjCJq7CPfP0Hwp61CcyyzaBGDZDd5n+NfbETeOVjDVc
yPmry8XWWaRebEA2fs+GSBXjMpgpA0IX9O0epjOwJNa+jJ+HKYHZeIGYBBQUQHed
Z0Q2mIK9Eqoj339iOfIkWL1tzL3Lp/6ipqZd9oAOXU8eBdyuMS1Zu8v98qD6//qj
ySPJyn2aEKfolfCXbK6PTFI26Mn22RoCRYVLeFvCjTHDtlb2oe3EbnXwj1nFZBhm
3+SaytQQcLkXWXtBHCxrc3IwS4HnHERi8AG4U9TDduNYbiGC2nz/yIRTnkSV7Lz8
RcBazfDprWLI62wyxIedKhFq/WjqgvecvIlgyzUM0lzy1c6Q7QDXtW6W6YJuW1Bm
niBusxMcRQ9+ILzWZbjkJ1ydc7+hEF1Y5TVnGEyNR+neciA+NBpFAN1T8sp32pcd
jIIEBPosnqNNpT6zUVL2YiZSYYX+aInU/bEn99bhDVzX0WVFnr//mgAzceARM1Vc
PUMRwVKScQltg36OsMx9Tu5FRVDlewkzVVd7nL19jRLgJ3th91/p00Vp/+6cUUfg
GwxtCfjF5KjJ4XOVHHbkOXSiNKqlvjaZO4Hmn95bGgjhd0OvhgUCOrGLjX50Pfht
qp/eCrySx0g0/aOpHXd0asTzpbMFD0GTondyc0mFXzdU6KSUapyjKo9IlKs6O/8p
4/KGbWduu5qy5r/7NPnpBiasBjHjSrJVm20m79DvTmRQeXPw0blWzV05iuDGJmNz
4QUBPwPGFD7CLPGJ6UFHOndRyJ33UxHVfokrsJXlSb6GasQrtshOPP53EGXlbUoN
Zy8n+hHZo2fJakqQxw/4MMuDxNaJuP61T08HjzjWBy5ffyyYT7G/NXETys8rIRDm
CHoFIEQBWD9GklqF8ppcqHyU3DTh63xgC6FM84QooURl9Orm0HGL4sOa9d9sS2od
3Hke004oANhtbnDHp5E9oju0mgJDvn7hxZBGvqE1oCVE8lM7610Ybt8BXmgwq0+4
0/7GMK1vYZ+B6Qv+eDrjCrlmPqJ5CMWadcW3C/kDzzj7buhhDgVbFFMb2nbZsefd
SPbO/BJ77gEZcmyuOsT6D8QsOuiiuqnmjtdRKFHCt/pCMPlehSzk4mhGFyCcY6dd
CY3NU1kXFND2nVdChflk6scrcrHlYDE77Tk9nOkxC1AsMQAXZd8SoB7gqHkEdMN9
LQ0ESzvmAAePntPS1IXTCcsS+1ax1+B4oeSWyWD6K5sbKMg/U9dHx5rOdVyF5Dr1
rYUfOpqpX17d5QvNNaO5AblF87sa44QilQbf6bJyeBGPdV4ycDdRIpelOhND14j3
iXVEZssQZd9hTkmg+LaIIM/ZYB3/roPPiu/kRHQ8TREqHdMHAzXiEoXGt6XPUu+i
9jvAA6FbtEuSfbbGEPoo0UnzbgHCSSLUx98QHHl11fyDBrjUofzjUnYcpD5rPZFt
2cLj98vBXH46fpiZezmZLnxqk7YfU7lXapVBAUEUEpGVBc5UAztR1fT/VvNWEnHI
57k57w9dgMM9ct/nXQJkyzrJb9HpfMnP+QKAc/FPomk40KwqPw+4bWSAOHRRAuxn
53yI3liYqw5QQNgXpCX4doyhgE8A5qdJsNpDud166qJA9F710gMukr42+c1IzZnG
ECaWnawRo5xOoonMp3cgO27WqbWouDlUCAgkH6SkTwgo0czINWSbHvrB1MrCQakv
+DAPNS1avMXeQYcyBWzU9qCu/fJd76TlxmO+krJEwL1C3TXWXStIPFGisB9Bb6hv
KVJKwdzV7WTOEX+bIEgIWGM1SPPi8ixNWSN2loxnIBOAR7ZmlRVRXMLrERVlOMRa
sQCsgftWlIpO6FMcCxiDoMuY+50JQ2iUqfc3XoNYjSWO+Ua3KzGNLzjyctrM5wC3
8U/nUOM5uM5/Grr+ZiUAgmPuDYEg1p7qXKC5szs020fKf62RpXx9L3Pz+gISD4ya
/k2rTwkGGHZ8fZfhLBxaxA1B30Qh6ebTf19wlKsMSs/uy4I7AIm1KEz3bqdZnAK+
4dIXZ5bu6bwQrMQl6sP4eDZINV5ZCruO2aZ3e8x7EA50FuRq38Q42hjE0XCD+S8t
B9YmylawyoEFgE3X36NNXKmb6Ov3MoYLG6Z27/pWQ54lIp0ni+uKJ1KtOaht6XWq
0PIIR59FQG4RpoqITDTyO/RbRDzh6uG2a2x782vtj4mRtS9OYgPsBdqRtT5sAzLX
RR0v47qv/ld55gqgZ3xwH2rlryxl/S1ELDc2wZN377uhu4I+X7c19gcmldmW83Pp
JmnUcskoVwMeGCd193XNVLQ7PhiTWr9XE7KVMXqul9RDT1tibMafvB7t9AVHgd8u
EnpWSj1Qonb0vV678gAvjemBfrSaAqMKVbgDXWL+LA2LSzKwq2vWRzduzLaZIV5J
IKkFfpti/GqLKag0sc/lg6fK8rKUozLQ7fCJtSW2MpGNULighwwUILVnyJOKNfly
jcqC574AHPvE/XyUSJgNi5eNtOMedPC9I42dKF6fAHABr7xyJ7MpWOD1B8nVJhp2
DDXvSCK+CavvpE1VDItvosyJKajb7tAiJD2SOt9dD/KmxCyhmEfF1csu/DwDboWQ
tOQwpIhI1p9R2/iGLJUGzQ2/jEQIjyQqY8ku/bq09TgUK5QELbVg/CrKtAyP0FLg
ZHo+KIH7V+kRkiHq4/9z+jDDFM+Gr6NUT5bVsUOQZHCCNTiT9zPVgDwqP2OJMMXM
hXa/jpoUuN6pjSrJpHNhShdQIFZYHMNyjfeaYTq1wmkdaAwA4T7BnqltFQeN9A6F
iURQtSq1mHJ4FJaziJo6aYGHNMCiVNLsqHipPMSgyabY+ORRVO6qLr00rGCDdc0c
o/Ky6bKjTrHeKtuuIGNbyx3mpsV+/ghKzNzLa7xX3LtHQhZH/fNvqG/lu47iy3Wp
zv2624J82nnOY6/FjTzbZKw4ezlncbMD9UYByfVxCtt2UqBkt+UDS+XpfFR0U18T
r4vDln+x6dmzCtGQx1cG/O1vw5RuH1C4xMsqmoBc0F1Au+q28WtYIsZQaK9rNOwE
rV6toQY+uTt0YT+qcnUdt2zFuPZ11iHi+Cqlv9g6825imXoYsejfDza429d4xB5d
IX02ZRqGyJsRMwCmm46AjVGsoxnQovn4oWHDiLGgWz+aSD2PVmnoyYndfjw8CNeI
Uf4k4kPgj9ZPm7+4sYRPsXAygSpcgSo9jnuhQGW/0JqCzVJGskUCjgqY872qrNC4
/DyQTHcUc3u/e1ydAwHWltsMmRUfJFOj1/cAy81F7MFrIuKdXiLoD4BcxB49yzSV
Qs6tsttAx6jROpzt2efm7qPsRpCJvnm40YQzNVDDno/eORi6Fd53jmmWXBoR4kXg
pmAANoLKzZBxhw4Di8RAY+EwwDQu/SKraOuc3MsqcWQFUPtk2CXlZaJuOVWV/vor
lXh+PyHl/a9uXfL03flXSJp8M+HCsE+tettU14yi4K71t/uGQa1jqv89aQrZwykx
tLREAPAsbwuLWh+UAd58nUwMCeYKujFw6HEJvfD0BANsdteg5HkAadYMoYDTW2zq
It0BaRAa9ExeXHcU5LYxTvMDjcVRmr+4uMrQKK0wEe7GEGEaNFwzR6AlZHXiS5Bh
45t7pBUe1lmwJcGhfxNoOKFLuaTWdMP3CcsRt8To6UHd94W8kemsdo1pdPU1YBUQ
xC0lWk95BjjNflNVILBkW8YBbOKc/yvj+Yh2WFKlKj5xMK2Q4IR/IFydqc2WVdpD
glelJNhDZc6fBAMN+Tm4+mhMEENqxJf7Kmb7kTdbrwG+zxnNJEt4aiWvrprWye3g
VwZiZzsJ0Itr9Pw/lF2JVsLCi6ZLy6Rz4KCU4owsFjlHab1nw9yWqA1wKbB5iDao
vE84pQo0cKF8IpYR/YsIeYi7emHXPkpSLOF7iix5Ib4cJJVe2skuM5zcnIAxI92o
XLqevjoH6AF6cNLpghZ2eOT0Qof1MxkQ/0BaCeoGgJX4dE6vO5Xox0z8BxlIGCYg
vS5hc6ASUf0DVaSP0KR+RFA2hjK7hApbgP6IrZFQA7sOqRSDsVb/tdE0e3hlPvYV
36MbYegbYTehpte4E7qIG/l/+HW1BPnEJQMIl2tHOXF8fISKtM5wyuKtA/qvB/E/
ttPJJIx+zgcVLnHaKLggMNHatCSV6n3r0AVZqckauFhv466LrDWlodz6xJ3/swsd
cd0b9GRvV9x0hZh+P9rKGXEuNT/LtKMznoSvBb7hIC2fQ/hPgros9hr7gKJnXvEX
Tc3MB363N8AJypF6IRiUV+5j+X8+uRAlEVEaKMj93xg50EXF0+OEVLkHOl9ityIk
f6vgy2EsUF40E/W3pzIIsjwx+jyzL1g5fDz0TpElXJ4wTln+cHz00O0kptSCvfio
mne6L3jBrdxKRe9J1Vz11IAF6ldLaGwN4vwis795dptL4BjGRKP3LurExeiUL5q3
u+psikUT12gcZ3G+e6ayg/V4vpMuirmzSpH8MBYbcULIhTKf3jNzQ3fuVMTPUNcJ
TSp0ELll6hoBFXXqd2c5hn6pP/MXRUfJvaPham1HxXuzACxTl0ZbT8NMxBdJMY7y
mWSGXVAUsGgzQb71TQpP980D8YzwnYcb1W1dTjqbjjhEkjHCeu7D2ShQvwiQf47K
O+bmtDqs37cE5Y1FwNM5BAzvdE7R20Q9APXxzeebBKZuWX708hUjbzR/1L/MDZHH
PsjxMqBtoJtoVoHfL4+Qa07OenHDBWXsWpd+JQXHmJwlPd14Nv57IbRKNMrdF2MU
p5xXRIJFBkLCWb/pnTPaG1nK80XS9Qs/i4S5OSPd5C9Oga6/jS2YK/9hMcexonAd
MQHd2IaBxJ+ugjW4a/j257zTEd+CQV7L8gOVSk7urF0Mfedty6wEUQNWD2iunAsb
80krxbIESoQezcl4CcYi1nc9HflmA11896WotPoW9uGINOd6vnETCeJ1l8CGpyMF
LKC/JOlnxCvhAiRQvPoRGNuDJXCFhS+quJ2DzQo/xkCK1RQjc5jc1yJHWmDnlXH9
Dc4J1p3k2gaXSU3ekPZ50rwROHrCWJa1U1aVzLOIC5fyvCvEQAM89129atvRGgUL
fITdSDK6TTAWOD2S0SpGLlCMSm6Rh9AOWoC2swlZASIMHEW2creo8X1yBJ8Wsa2d
Wg3gN8PzbRAlR+7XbIDecl9XPssqh3b4wByMIytYdbnxeJevRjK66DtGCM8tGbcu
5qMlcVwJAS6Te0nObKeAg+J+AWTq9CeTAvGLUjvPIO1nsk8gsVLzMB+B9OTl2QH3
e7x+wCmEkw0VBOj2030vWBHnGnGNv8nBKB2+PhukFNVhy/h5MDdvMS73EFXzX4Sy
tGHKek4Z8YLLWzG7P57DXEP03qQdQXi41XVbKRpS4ro/VJMmN5tg3a4pvXQvYM1I
g5P5f587GGihKjF91PU1SJQxaTsP3jnWkirIS3aErW+eU4POG8FZk7cY9ETN6oZM
69yx4MrePkhsAfCxJbO7DaT8ZxEr2csCAVxJ6DrZ50swOYXvJ5uv2fQmHt0T8XFO
YpDJEkaFCK+3hfxV3aHBuw8pPuF0Krq8kSCxwvSeX5P0F+HxSM++MDEhrRr40hdQ
l/9IMcT11y3h+u/B55Oehs5tMAX8JI8bAy1NfdTyIxJFZKGWONvUwgrWKrmIAZoF
766LoABRsNnNf43BGzYX/An+1vtp+SLhabXCtrXbmoSL62nHfwJOYIndIfNlGJNg
0cGL+1MsdMqzVQ0JOoaeNsgzdaFCstPSUDUkMRG6BzwDf8it7o85vNihL44Mskm9
fYupDQvJiFTdyKplfjsoU/3S+xgv9Ol0UpxakdogeQIzLEkqjkaceI8sJ1yATHyS
1wDR89aNQifr7rptbp/tVV5tIF2bT2L2/iwLOh3MWnfymt7kyRMSpNYQsNoRGs8F
uY65fMyknRa2zLzguJ6UG4F6sGMeNz996OH/8w1I/9uLiDUxrDi83CjIOe8+1KYF
0LwAQH3F2sv4gVQ/31M6PcxYlFIeTPQ0FNYieJEGAk69F7EZn2Oa3zfbWz1MMcrp
KmXY6puiCQ3AArRFQ5XPyFASU6vtJ9kJKfS24MOmvZ5yl0jMtXOx6ZEBj/HMiGUL
VIcz3ftQR2Xe+WyXtUIXqpxFHnaxVLQ58MPGpODOUV04zu17Dzom2Kp/Z0YFjnZ6
56GxxR/wKHNViv93M8O1OwAcG5S7wiy4Yr8JBdTOfv/kH+dGOujVvXROD06V3uFd
HIR54UrBb7zqoDfeMjSY3K95K/PEIOeM9IUDZmbqHuVfITl9u+KvHjPKVG/bKsV8
LJBc2eZlOsjalfwDrdf7fMypFSY3mtOKuTvLKwiu+44imLGdd9PfhUzT6h5XIFXY
e0+alQ5IoGWnU/zLB1m8KCM5Fx/R7xhR/CQx2Y65IFAk7goxNZsqqSAZE/m+8Sn+
jSofOntE40CUzfL01nc5AKqH44Cowt16mNwtcZUl2an3s/ZEvjOeizfh7F2WThdU
J6aVrtCsBM8WiThAbc9YYTFhGsDvjXT2EF5Yx/rTYqmgIbIt4QoNpS5aWLQ5QJH0
EW8XZ8s3h19CO0ABPFr4bRmzvV43l6WmiwWr47crBRpVtZul6/apa6e4Vv3p0LY/
bHV+QmPni+sT4U8xmp7Iqn0qV8+1aDOx7hnIdeQa5aflw2LyNFJLSlBDBkJ5QJc/
yNNs+JHqiOFvgm9qDEQDCRF1b8wpnnWplbkbc7D85DSipOpz9tIKBWp/bGEXZBHV
x0/LbrLBh8kXNVZQUmxjWlfZoyWDzvdjELRYsqeoK13SNYjIwfAA0YACNfHhhY4A
8F1ozcuAAZ0IIvGrUcTe1oCW4670l9neiQX4HTig1BmiGhkUaWc0CmOjva9ji+gL
WJgUUwP3n3pe/31oSOKGodhOloYv16a0JDyVEUTvsNQy5zmuYwXC+d4dAO6tphqQ
VgXb6Y56Bs3KldItVCRJ0ItYfXTWECxuIuYYzVFhesCuNxoG7yMfRjZbojPOBP6X
RvWdrmJl000Zvx+aiDqdMYbxc7OUiqvEPAR2Xx9C5nIuFFe9FUJ03j3lluaskXY2
jmrs7Tf38qn3+Tys4Su2zmJzkHmMXgKTdwUIyM9VZf8B8rL7bZuI6BUNPQG0oM02
8BXMgzT1d+JSAZlmQIomYrcgCH+tLgnzPj27PqG/C0zaTxLCX4Q+4V+ACXqw8pQV
CK8eAHqdvGMHhpclO36yrOlX4U1dv9TkLoW16JH7Uocgvj0ALgX7I1tDwnmh52hZ
hmWhVKfhO7FmvnpBNa4He6ug4jiV/Wg4lCF3sONe+iOGehSJYfK92ppKr+8shtYk
maNBJaiiDgUzAxIZlTriJETBuUOpHp1K34aVjXi8vw2lQEXw/E93tNCSmWIOhdlw
qvZvw9Pgd6WDktVM5TDPaomcg7W05QVz+n1qqTcttlROnUeloysqyR+EMrAKW6E4
yBT2h6j4YqJz+8odrhJ9Y0ZlIZKYSfqpXP6rtinEr4AtDco5eYp66UN7oYYueVNU
/AvqIUJexEKND+DQlDL+KWqVHjg3tHDJVe70VEG29v9CrO9vhm2VNtfdv+WYhfwa
KGYVyox3vF25Q1s1430woikFg+z8Ly38lCjS56YP5PPHJwPxeD+w8vphcvL+yxM1
UWXCvs0+ULORQRwPanQBcAeK7gnmVgJBYCwtw+0rjJBjak+yfvfjHQa/yT++LF5N
8Lx13MYdrt8IWL+luXmx36opQjV/1ByKLwdMzoew2t2ClhqBRQU1Gd8OIRAY6p87
djslgfVbht+u2zqt9UDtP6d16kv4PHiJAyqS66mW5H5t685Psi2BmyLA4oYbxPhf
nScPoaVCidvu590h3u7WD9AWZCjRN/9u8G8eie+bQQiVt/6Ze9EaiEZrTQxZQH6M
W/iPqoCZm1dXg6yo0ZWRdtWM+eBDNvLwbonI+RWWIAjfi0IpQpPFw9EVXdbU28iZ
Xbp95CCxp6RzlDHuErgxIKy/hKYXuDlXbWQOfXwTdviY76q3ukbVPRzJVm7Ru1i6
9+JEwxTg8/DWuoijxTea8iR5/1PWMQnBea8cBDKQqq/LnIEk1Uz1gQUn8NAOxTE4
Leh/JzHXZd0nVtvqf+Pe9prUPM0y0uR0INdP7NjUrKBF2K+D/a2vo50pY4M3AUhL
hI3DhAyTOcnqToUE1Yo7oQp4tfEA+HzccPaeO0KBRFZWHEZel3PNh3RSQMNZR9WS
Yv9KZUPlUild4AXX5cqTC6+WY8ELLsXa1FTNtL7VMxSzyRyv1MI83XinoyoaXWip
h7IAxbI5TxGf2gb0eC3iXHO+Fw0+pQeWbBxjbIP1UPT7ymMLziiLB1GwjZSZWbuI
0xUUTUCrYZFdNAG22UZdBU7gTFnfpvKUwqRe29JaXhx7vrygS8kR1JvjrfxORANY
s+cQMtcj3337joBLv3arcnlBD88Q2KMJ9vn+mReRnQ9BCZI2NxsDtmIE7XVwCquj
8If50QQZx8EqcfUce4QpbzKPwfYkSBQiZO93CxciH2IQiRY/jrKNZhYX0WT4WQpY
0kNODw5DDIfe9GovGd7qK3eFygyF8Hw4sITFy+S8KLey5BblriSR5AfsBPoDvudO
LkbBP/4n6M+4AJPnmwfGWnJUr7HNamKThNEp0QL3sx0CrS5qfto2iEFtJILR9m3H
7lFjCMKsRZeuqINbGA1eUZAZLJIJ0+eYrFW6li4FePrupSpYKZfJfcLoD9JHGYb7
kcFqUSqieQXX3LF4s0BQ5OLQCuEvJ5OCiNBrqlQGoxuBuCm/dTKwgviCFnd6Kz6A
dsB1i7UpDGtLPSTPq/RrlyRkBWPwh3ccyPo+CYr1gzbgIUqMKB/3W2CP9InqL6cU
tWiUki+inss/TD4vLd/e6b0pG+JnXrsS3QZ11KvYNia/O/1AjRAuJvCqeCLy0I8C
0uEJUWaHiR5lnCPAihpx00Rlb28jLJXTZkpXAKADozZYDbBnYyKdPJsapylL8AuX
QxHMfQeTx32Jrrrv5mVkch5a1tA5dsV3yTsZ8HBgj3snNKB7XbX/kyzhkHYPcieI
LTCS6S6eugc+Q+kCXXqPLpZ60qqqfqzcD1dRhGmiw8w4FCxkgQBUR/MV7SB3d0Wb
WwcfInYLlGG6OB+saAHJZbffvLUD5IJwcEBc+I/2eT8b8049Dlu/e9rgF0voR8P0
zeq2aP3v0/Z0PUn9oBBPw7Z5hbPReDp5TI/IcbgL8rfa9uKWi5gGT4/RP7HO+YoJ
EcMCFMhK1TSEZSZu2RAJ8uVivia/ts4heTujo6dMk5D69iPP5p1SnMZJT/Jeyy6X
v6AFe46fGQ9DgUt+1X8n7rgLtQuAlsosVG3aCT50dCNvJbPMzwyKGNHPf4LK7uk1
BZlHecQTCmxhO8ZiyNZui7rRia41BO1x30i6v/tIbqj8kY7rrbIo3Xo8b7egCGHv
RYZQF+r8E4bCXZn/BQo4bMmw2B1vfDlFDj0QX4HWhFmT0SbmGMp2JMJmfLhn7k+T
bJHdLks8W9ToJvR0FXBERfg6tsElVOb8KJYxWe+gaImaSm72+v+mqs3YnvJEopr9
eUmRCGZ1LRJnTqq271uiKyymGWQJRbY1B5UQ1d2patcM9jmOJ1T80nmWarSLXh99
4R63UQyX3exY8s/QOUN7OHcfWoHGB2l8Tw7NXEPxCDw/7IBOyRW4V+DKvNTfutr/
vrYuFAWFos0K053oaHKTTQQYE74enWcbxXwCJ/4j41/mcRxIQT8m5jUTCp0VLL+Y
WSqODZ3Ixj1pDO32V6p7dZdVsAB1uYMr7GnplscTjR5g60lNHKg5bSxGTMhDpLEn
e/vYrErBQ2CvCLVHbayimW9J2Z7gTmsNC91TkE662IcFmQlr2OpaiJKOuPaIWAyG
dPNGo2aUw66QnYymSNL0iJ2xpQGK8bJ2bjd+FFAXRqI5ZBfQo2S/dCk/RhrTK7sh
92Cj6BqOXOwx3PlVyV1ZXfpInK4k90rE3OoCA4kS6/HiKEcSyorfmde3M7CV9u/4
B/bAc8Q4X9KdOOUtUdG5xLoP/UTZ7xJOqw6GbbVlfXGVvZHCtkrSfOlkWKj4xIDz
VjpvaJ7dqILc0INV26KY7G3VtfJ0hLWGDYkPQBYtLfmaei55Syu5VEYVBT3VGOaC
IrZUATdFgs9+GF9Autd2zSIxMl9yEDDwejLBRoevpTHWMGL7U1P4cO9nyRhvB68R
vj33XiwBggM0XUSrtwGK9HjXQNkmcNjVvk70ghR3qxLxB51X8ApohUbBCfNAuJ1x
dnaRWWJwrOtCH/dutL3mGdOusqmWhJ1tn/4uWm77SvEF8DtP1rUM5ByYcOB6viUW
YFkP/3AuxIXoTnz9KxzXLtSospXDLKjEmHZFUpVGXC1qQwuAv0iKCc56XcLSLKWK
XrgkZXoPy3sRkJFpzqJd6aZnSx0BSsHx/YAdqUvJhmNjSpMLmnbVzl8beDKGujde
EUdXT6UxHtlTKxte1UkQXhw8nadxmlsZcvwlXfiOWdsk2mxwsuiCIkQOXoqDaLKa
flClV0tAG/Dn7kyv8XTcPs5KOOZcIGLhQRXuNvAFaqk7O15s3DbDJ5UFi/JUxfUF
dyiOtL7WgJv8V/kupVhhDDOK7p/7WV5lrkI3/nSJKbFlLX4/wmkSYK4E7CKRrzeK
ye3YEtBiF+Kmb7o+wtWpTnvKdr8xaKpY8L2FoAK82teVstx5oBDan/vBKSKXtldj
ZMGHSPncRfP4LKDx64Gsf97DM9H1gxgCuZSBaI/KeKwahWST0yevd2aZ36R9J9/G
FwzNuSe+Dx1vXLgiHW1stDg48kmrkhmGv0u0Ofsdvfuum+WyP9EMEtnX9qer3Khz
EolOm3OMHz7wHs1dWntceNz9TDOwWA40QjqOtPnEqy8eJf1BYO6IzdsEY3+OFBAn
I6282Le096V5SfHLL8EAartk63A8x/2mVGfUKkHjUR7aTcxH9t/cQiz8dnCz4Ho0
e56lZ01HQPqn6IDrEDJFaXq5SL2XetIElivPzBiZq+0DePE50fvv9/ntgOG/I5Ms
XjikAL8ZaN71CfiML3g4xtyuIf4vlE7K0AIQA89r4zwAGInRMIFxLw3xITqMOwVk
Ry1q2zuYxL104I8c0XC3tna5hyyRPxqWsRXyXKV5cDU8N8e2178bxykrjAOaUH00
L6jlMT9aCkxacxM9G7oakaY+m42MFFSpJRZ54js5ChOeIDyUkzrilhlQZFuKEI8g
gAF8pv7NqC9BTP8itzkP73ZYnXGI7VHWvZ0Baj2j8xQB1DvCBqOfhSnSFpJufaR0
qeiXzOiItZYsEWDxJ8cZy0rnHjHNiQ09Fx+G3dbRAc25Fxhct7XtcW+iUeRTHzvS
BROtHsO0mdj6WV6w7Zm+IkJYe5wUEetNJACYsYn1ES+HO0IYivCURrLHYniB3f0z
DI3M2XJB91JjlOz/xXMJvFMOZvS15OeKqTdM89yUEVvuVgT+0I8BqGIzXqyhx1Zw
ymeO/qI2eJpkHNDvr4k2rcG6QI1cTzBMhDDLWMZN50XHd2ptcWv4P7NOQEOFf/De
uzKVytXQuqIs0U61i4RQ9EuJxdun9aOkl4kH7FyQJynVWNh4G7P1cfD/jGzqv/nl
02jLIjSsqsm/id8KaoBK66nUuS4CrjG5RJy/FXbe8FD5i7FuTySerMH8YS87yWLo
KfwjlceaTyaS2xDGdFmOi8vp+FEEosU5Qe1fWHyw55i53FvIpcVHrd3wHUojhAAB
5L945hHBBS/7bNN5gZ6f1L0V/9zaR4B7RvwhOoNdYNOKQhyAruq9UpxOJBT0/qEw
ldLjQ9MlyhCJHZ8B6sQqBGoR02WrRRUTJCXTPUuhf/CTjVJsP6V4saGUbaN7PLHd
jsqOIkqoUvLcKdCmyzMltjfCOj4mlq0tW180jcirQzrnajSPN7djkZRiF9uG7uSP
qKBZ/T9U94Z1N8pP8Fan5Cl28kW+YJTSSyEz2GsQifu6Ef3z7xAoZEQ9SotMWlWo
BuN+VDO11M8Vn/nhYRtMtIe3P1z1yIMoLg0waz/vC4CgeVS/3RnRjg/s+hxbN+e6
ZqBXB9/yrNdZR//rEm2AQILbFR7EhAgzqRPUriBHRoA+dt37rSaCawFGvIr/CmN5
mQgCH62hmJkE1ENd+2c+UGClvUIv4BuXMn3A8HhovoF4o8UTNAVz7d4TGQjxmu3/
52uNBlI09xlBv/vZD7GSU9tyyq8VqZesrAtQzt23uYbLZONxjpmhSY1od/4GQE8C
NAvDy+64ZbZCneAN+/35S4fDZqQHSETTmGuh5anM8nUyCJEcztDMKlUgEOiXNx5I
2/g8ythx7iwRV2KqW9+MJK0Gg1TS7T5m5mxl/SDSC6aW7kxcWdu1mgXTp6YGjPGF
lL/H2EC5ey5MkNblqxNVOH2q6NPevIPqOIQGpOBolXL0FPtqJM0wqdDb0vkYADGQ
VK1GSj2OiHvjfrpLrB1Kc/yBiEcPKclwsJwFm+cgE6Xx/h63QoUYsxo508MhAlcH
ogUHr4q+6U7Lw4nugbm51oiGthQRGbAi7mIVI9BBjCV9TBv0gIieF+9il4QOyL9k
DxesV2NdFiTKJyVe6WrMxG6hgoeOMyW6oofTdppTjMXP8MKXs7yyinoMdUZst0TM
Y5TT23nl8tprBtzmTTakGVIObjHhuGp3u7L4eW0ydtVxiSt42s1qNa0e5GM4z75z
vwpUOfRW6GCFxcHBd9Axqec0qDAT68tTSMsuQF5T82Bkjp1oMFLj6BPDvSuhWb3U
PzwYXs8PrF/0kH5jQ5wVpzCfuyreKfpwOSBI5aFCcNBgTeGUmhsIwMjlEzbQuUng
axqSWBbc6opKGF0vDdg8CF6laxVA0och5wDabtuoaX3+oae9lD2IrZ9pFLQnoJBm
2DiTO9LFnevmK+n16XUnoakHhGIwt6deUtfzNsCIeILkleBNWSRD95Uu0R3OgKHn
oG8WCnhP8Li+5K9cZwX2ZtqUqIoeUw9LGU5dyF19xQrnLC93luUnkr2irK9Qe9do
zLZ6vz7b96rRhlT+IUEg6zVHjeUT3OhUTEkTpAw54t7qcxZqK2FISw36LHvtMsNZ
fxFKI68Z8fZ5oSQlIoe1VeEqGsQox5iIsdd/Tj2l7FjeTyp/itu7BuSbJoeSWy0N
+5XvZO/I2au0xsCsKY/BZ4mDtIldILShk3XQkS6ZLCbBLzgC36rRPcXo0ttPCB38
cQ/Kku3zpUbPJW7q588UvumQLyn+y33LyHyMVGhz2q6zx92fWisc2NvOAeo5i5O8
1JlYHdYFe1/xotJcyRSADgHm1NWY8aHMCzX4zgedtqOGOhr3B0FhRlpHbfGJfDgn
o1dsUEsHfXpSta5Y03Ovvuv3D9jkb57Bidnk/UJE+eqHzrJQK7d0zx293fRZ+nAd
TioSL92PnxENO7vZ+IbZcv5JzcBV/JamHCTGb23jASzHZ3QB3v5bgX+QJTj2Cdzm
4ocbsIP7fE+vLtRXZrImBYm6qIyKT58tJFN89Afi8DV4w+kJLCQz5K0KLjBc0kNx
R+BvlUMdK1fT6EOuCiL5e3KJ+M6AbcnsA7DXJTXberTjb3Ft/VkdVIOpYTZA0i5A
24ZU+O1w7eraTTtVI+m4iw3lMYpOEevO6QwqhHs5nF+lH4K/1aDcBVFy8kExyXa8
OCpC9+igl3WIvH4t8EWUZaQDpWVxPt8hlFW7SPs0dJ0pfpKmymHsfDTivCdCIGXN
cGjOv4Wv1aQMgPmgATUYiIuDWCNv9xV7HwYVkSJ43AcPNAQSwcMjvcWx0AHDuOjY
YMhC8BPtzeX2CEkbaEgcUUrvCZL7S4xE7W1ox0GV73Kdv3HDmDNu6jG8QIunDxPL
cP8K+CVm27T+La9bPmh3Y+7fIzq2EX8sttMYi3aiB5GchX/bOoB/Qi1FEYagGTFy
shMEATVtYtWPlH2qhQk7u7+S7QqSQlUzM7cEL56TJ2gYPrl0RpITm9CpLDYPwvxd
KnePnuDX8NM5Cy8QdfnZMru0hPCnIOKTTNaR3yD1LGwJjUuKrGqMDcAOmbMQKV2g
DFh3XlAaFahT9HEhc8s3LzjejDbEz3jMB9YlMvyz9l0e2hyCQLv2SzO0gXN7krG5
kGbtAixaVt6IG5D3QmwbnORG+cPwelNJK+jC+Hmw4Hwagx6dBONSLZxrit/Ww0/B
+RFiGrtLU7AuWxjk4KUInWGxPDyd58hK0MJYHmr5CriHZ7mLbOVUuMJ1HpwbDiU9
L0He2Y+RUPEjoFdcdDlTNDYLpuL2L2Rl5ira5FzAcTbvbI2cygjo9TXVsL4jrejM
f3nTLoYgr/vo4m3jAwQ+87R6RrtRVrgU4rn8ry4siq/f4zN4aeaDDlyD5rFVqARG
pEOMBqX+nEi7Bs/mqmoOpqOepDrN7XCvQs7QOXTrzIpAFlsKQ+uj4tBCPXqgGRm4
eP+Cypp6KYuTBWRmXisRJa2x+RmfhRzC/RdXu5jE8V3tVP7PFo13KnUm+dnWiDUm
wBBSDvqpUJH7uJDyd2BiQhRczju1dUBwnftvKcjC4jP1t23CJFQwMUVzE3NNoDAZ
5tEc6Ij9JO0g1SQcLXvizCWRVB16s7XEuTi8t3XSpzIRiP6MHXOVfFWJ6sj+4Pr8
/4J6fRA6UC4jMXVpX9pBgQWOq8heFX91Jtn6O391O8Bhj99wpR8W9cf1ta3Aw7eN
5vKbokzszCoj4BldItiuWwvEIkXuI6xHh5+v4E6bsjdD0btjngAzRzS6BTJaWROr
b5OU19K23oTmCbza7cgRiS2r6eZ06GshdqxL5kzIF7dq6PypyyXcUsbUarFkLOfr
EopcwAcLk5WJ8laigJtaFIBSBACG9g5vV2wndVX7Ye2Rv+foYsgwIG64t82qAj43
TwBalks+x3CXIxDRaPUOIBnuOXVc6leeU6fUZE4hRkYXepoGIowZVMouy24Aowlw
sI7qUxI1jx9A5oku6LoOkDfBt485swwMxPCOhg9wceYkuMxGLEDsT5ZyDqp7H7WF
iSsVOJYjezwWNqDdnf2EPZhWXZQv5l1NZtbq9HUOAPMsOXBx4GB2B7vDK/9CCPyg
Nrrj834Y0xN9PCUgdvOm549H9YZhokIH807sXtAqTIUqWru38AhgaHuc2OPCHcDR
+0lp4v4AKzZCoyMvUzidI1bCenA+WgQWm9RatvBlTAxL7Vk6CuKRjzefK+p9uOdd
jXTzW39aIGusez2+pK0oigb5dfkC8RirU0dlDZmGTGB4WEW9CBCTD411X2tivfCv
XL4oRKhOVf6vyYdVAljy4RQNyJ5+j4v/rAAmVtn6wMjPa65zyqnOwWMCtHwI7GRb
619TVtQ2rNs4IrqHWomg0q+GMr6Y9fOsm0zlBA9KWHMtGoZ7WFVYYhZVzygMSPpm
EvB1jwG6uPnNdmjoPjzF2o9SjC2yx3AfsAUu2LmiarkdookiZinhEc7yPlMPTpLx
U+dy/gIo9WDjuHMPCrVRepBQWl1Hg0lA79OQDZaM3c0WO/wC89FyXjZ0ZQM9jwgT
pShpoqoOiVrEnCOPjI7d9ZQiXSJsShl2PdSELY9WuuRtE3WaFrS5IIV+PZg7RU6J
cj460lhEoQYwsO9cO6kgOK7dVSSfY5omKwv10wykQgnFq0x94vx0/mLFSi41JGVG
14fA3ffp2weG7pyZKd10sx+fWf9Zro2pdlXaVdAYap3dAwWqSmfP1UXNaH0rOJ6G
GHVce0AcJK/qhBNY+HiCHdMvuPuQrzgr9aa68r8kSWGHuUK7Vakpr5qQT+71nP00
Y3KzMk1qsKFw8GNNxo0/j/2HD+dHEwgNgS9A9k/Pzb6yxH2ZQksOhHAV33svpIq/
t/Q0RqUDDwimR3aZnUJxBTBmdZLkSMRgv72oK9EmNZ8ST+Ri/WgV6pide5UxBd9X
5rNlNkhTbMDLESfBFlX/D9eptX2Zx4gL7vIZW/sxN4IAHvgUvWXlpmRKOG+Isqw+
DPbs1F3JkRnSeSZ83lMp4URvC3cSNQ3Y1MLaMhkZkTUh/bRih5VTL06m5bgARrSv
juB0kvVBZUicEGKddVl/yEgAmIOSnfMNm05jPbcIEzg6bGIviG3GSkusF/2pcbkZ
vivynvBmU04WX7RkccBSXq3N/i8mR/mDhPCtTsIKvzSqddxW4GMs2zGb++hSjbTn
bT1zefhK9+9knzGuq3bVgSFtT0lI4kWuGV5ZeE/9/wL2JdlAJysnpdHmELSH20E+
JH+uLl2gFcnH9/9vkRPWuP+qGOqFh9g9yFlD2BFt7YsqOcRClECRYyEtk2s6Awxl
/31+6w+urPY/qDcz9/tHomjAQ7mhc6XTIh0JMIe/cOn2rHDoirHAIZqCbqV6rDv4
HuZTikW6egzWn5ixw1SkBCaoaN6uCrAI/eKeiSOMQUaJfz6nUY27WmiLxV729o/v
uKnN7lwYjEiLMkZxcOhIUPqLhw0PccySv7vwyA6SPm8rpp9nF+WkMLW0jMMYY7gz
cYFp5cQaK7yEw4JrwSEynup/HUrcuIzFeD1Z9JwfoPb/nuq/FqEUcVQirklo2yMf
iFYY7xro+CIfWNa9Ol8dhOp0LNst2RPQsYcWSUtpnECBvz6ECVxzSVHEQCAgp4RU
2KBjoc/TpamiBeFvtOFMxvM1gSBgyty/MaSAtlBrz4ZnXXKrEBRJ8g+cLlQSlFJj
3Q/S/w804kFFEcdkFYToRmBs9iD0mZMBNPN67Klg3etwTx61ySz1bZaaqwItTH1Y
unbQs5sIG0sfICHmq94uVGwP52D+bGnSuCjzc0Ug2VD3jtjoE62ViRSmdW3mD95q
8dAhO5I+QrCzXygl/Hy6rNEruhRSxIsxR26C2Pc2sfH7W8A1LuNL4BdkkJArAbwm
fzWlsoX7Z3EmzsUCP88TkA1hoORdYR3ZgmJbZ/4KVd3khLHIG4h3NMKzLExp02XZ
E3eZbUIWRZvaGgHsFSt+UroZAWiGMPTz4UVeOqMO+0nGABbZKXeDcbmANCqDUGeN
HWThEaBz2YXcVqcjkZhi1zBXQMU42q24PMFQXPsBdro254b6S3JoZqQ8FfrfAKSq
tE8NjEDOIcCHnMCBCRZ0QzNfRkAci8AXl05c1P98KWDFDKEvdcliAnZJxhD/PJ82
u9P/eYUIwWmnhQXzZ8skhJDymmsUqIyXUQRMAuS7+LxzUBE/iZeCwC8jsiEU5VRI
W0kQXb7ics9nPgn+Eym8gwJlRrCktVj7fO2/HQC1RiwPicRdsKupKWj78H+LYlo9
nQ6aCNQ1jihGqENiXgVxlZEpG1y5/yuBWK718FzHmtYqoskt+oArbRmxLzObaqQZ
4a/x2WXcKzBSXlunzVje6UX24WReYzVuSnfm0ZUEDXuXHrg0bqKIXcrRb61ibHb1
Ock2NfTv+cTTTMISMmw9K3LbLKwPUviIglr1d13/3Bk+3vwGd4ec5LOfHroKqh+G
+gV9hM0A5fHF3q2UrN8FI0YTFoWR+7Pwq7381lqV+wBVUMoJzPfp7hqDOvSI9FH4
F2o4CfbQgz+bmPFhi5CYZSj7PSAsg+WY0C01ilgLSEtUB9QOsu0R9CS4w8vyQNq8
3t4PYw8IB8Gnxkxl/2RoTgr96foaIeaEwVLobktFfkgWdTKEr7bLntm+xZ6SrnD6
rU5RD1JVaoFdIu7BXgF08RP8grCQd4blRiIDETZq0ouwSnndFXf3Ei0u18BrS7Ny
DGkUP0I0kyxujBppCUBSkje3yvTL/Z+FFvHtyuD3YlJ5wh1SmMkR6/uv4nGCNE9f
aNr4YUxGvFVj6KjOO5TR5zvc/ZOg3QiuJrOIyLCZyIYYECM0d3Dw1vkl7iZ+kPUi
MG9SI/6O2Bahhgx9oeawCJov71s6hvf72Y3G2GF7p8TDDcArMjD9qnUjOUmtmuwu
wqfRvBUWLzpL0BrsUSCl1vGrmapyoJEVeku6lixdRBNFTv1Z5CAElPHhPT4fxAmT
/Pl4i9xD8kL6PNyo1HAaPJIYbVldH4eI1MZOVaCjt4HOKkKSa1SLq02GEs7gDXYB
Xz08hz0Hc/zT2n7BK6peoq4IVXPmSqMV98y5Ig8Wdf9hxn5SqSO4WDNvvU6RccKD
ZY/1yfMhtP4AZxyA8kfY6aNxywqaWx7utBbaC2KlzSMNWvsQL2C59sN7fxNoAZjB
7OxmwyA5VoKqWI3OIX9AxtZCo1L5+lmiPFWO+QEbM66JwLJ6q5mSOPHWsEVt0bhf
k21tsDe5ST+0QuDFDGEVexTW/1fa02/PmDC7uG8MDU6YHlgxqSpQLyEg+UAgp+1w
tbZFHgkEGveavmaAQcuYaObPYuFRCpzg0bXaYO5Tt7Dq88tAfODf1GhC/6puh95g
rD4OJhUhxLAQEIB7LINx3PNgDjSI/N7+sRa3l/xBn0TAvhfyKc/TA1z6VVgs3p2s
39kZemqkNxbWx8MfZR48BytRjETTzVHyau2+V1OAMRMudr/DajLfx5Vw2NUzPPxk
xNBt4OhyG9n3UD3yqX2PVWHrC2bGmCVtlwDRN5ZssVkdJtcOGBuGDWHHwrH7MIJY
SgK1bbKtMC6TjVWhbV9gd7PHWpgwUpGU/LROdb/RsC+ccKcl+3DgwLgaYHStdHkh
t5glvXo8jV+D4VJgDk5dFgrmqycf+WwT5bfz3Z65+jxfr5rSb9qLCJnIrkhIsfdF
jze7atYmagm7Bipge7g2PxBVs/sB8xcxinaEnDlHz/3/+ugTPVUZckjTtOXNBJbT
SRNZZBDjcQcI4rbSS2XhT3tVfG4LY5w8tpwUZ0XdrF+Yjk3NHbIqHJiJeHbdl15M
JK6+1D1IMQ8+Qw7Wn256U6nw1pXpyKjylRYUYaHRokyoZ/9hxch1+DVAQ47a43Iq
VJrfMPl18g3EegfRvKMcBDEUUUURxYwx7TzgDANaM70RkCqmExiajYrf/M3qGFxQ
m0XOo7WjE3MJddqFH64rIZ0pwESycuUcowP3T+v6QfFyhH/kB20KZuWLLUhBjtRx
4oL3YeH+v18lSvCLucsYyLuA+w6WFWP1rZbc9ll+KMMTX8uSeSDjaeQcDY4Pnz6p
LOQY8PtqheTMKQiKekKW1WZs85IeBufDayNgExOQUNZ+uvmgpCtR34wdLTw1B/D7
F4qs47Kre+9onr21D6QFA4HW7ym4PF7hmZlZlmoSTn3hvTl08XrIRHc93WDI3uFn
1POe2anzoCMKxTnUbHharTM3bw5Y1ygfuHMkL9Sdq5NckoYfWAOWdnEcKJTYB6R3
H3Z1dmb3p6Ploajt1vYPPvK++YZgP229pYQu9IJSfcm2NX/PhJtpSNXBjhaLXWKd
YeMBA+DJIE9ILi9BjXzewjnyB32pzmI+aslrw5D4ScCpNoRYLBdPXiYrc+H/g1cS
CjHGPMUr52H1QKv2XIckJSgkhU3nnmQHErwXVsrmSYEq1+kCr3PXJexI5CcU6zXO
qn5UxT4xa1VrQ/nEWaY5enu8h2qtEsjl8tFmswUMPqwz+NnzWT5coc9w6EVSY/0D
Nz2NO3T9L9Tz+C/UzM67UvrjglGtERxGW8SaN/ZMOHWne7EvaOwU58/ZYXhjfEVV
sdy2e3lVJJkoNuGOgqxmhVcenylXYhx3VcpL6WIOkXzOs5tz0aIzY0vNsqEeEXUu
cjY++k10e4zyWBQzXsLuOSesxXORzgDAF229SdojPAjujR213PnDH9kqogOvkP3i
lbSgR8M8DAlejvNW6ao1EJCbRY50pXTV4c4yEkvMK0nKCJYl3SVmTx9NHIPHi49L
eif9X6GaiWQ/M4i33slVAxs7oDeyPg74OI5Gyuq3s9o5tmzh9mCyxYvaUfSyBEnG
bJI7EOAJ8P4CgGNRl3i/NnCsYvCWDhQRZCZktFZ6XtwKBDWuH8Ku5nCXdBjgDn40
lLYvPm9P1TUHpIj4UpVRZaWF9KZwtFqzxr3WpRGH49b7FGH4mcOkxJp31iv/Cgw5
cy4yLXRm2H65ywTf33DwmFTLjFQ+oTwJZJogFbgXceVYyiOOEXFJP0IC5oRx6PCp
YlHI3mQotDDT2QXd5KuvdFp2AEV/lnWGSqlGZtfmZihbNwxwSKGCnDEXRdM9uNnC
YrWdHdvBAVnUACWYtWvxBoQ1mW8BzdyDoHITBelfFr7c4/u9tdV89hq/B/uTqtzR
TUygQosFfTvdnVuq+K3JUsPeAjhFJ6dwxgrEZU+CbLmff560jUKWMgazgXetVgya
wwn3TTFq/GsxWgOrfN/R2xgMwqz3lYHZeT/Y3NOwHWYLSiFxmaONRQPcYwAB4TC8
QnZ/cjwVo8a3bDppzoymu45l30i/75ThfkyH8QUvsHCO79rdbtGiXfGGmWxloOiK
14M3ZiS8UzhaAzgM7ZlN0hfUBVizbolfN5daAy9vv/7mLJ3PmoOx51vr7n6p1hke
AASqYyhSE3LPF8jmMze+MIWlPkQVJd0L6Ay6qUKsy5WKGB3Dpueq+mmYsEQnPF50
IyLkavBiCA/Y5s3TwLNYVTCWIINaq6rXMYBtsWrXIi7t1mqu+8PGz4bWbkmSY8qK
lmW6UpR+j1fBkjeMwtBXY5QxfGXnI/syI/T3tN1bJtkZe/TiRyZgzKdoJj5jVOH6
fWVR+ZDAjQQmHYFYvFM0x/ApG6+T4s8DMSK0/55Ihe1brOJwk1r0MGGm3uejiVkI
EjnU7TfDWn/OmGCtJ52deZ398XXfW06AWblWzJovcOzETwrchV00PL75hZ0pBQzV
GRzMx18qjrDR98haw/vLIkBuZojBUeSbqDV3+3fAjvPRyoSpHJl/GDbAjBaHaqgL
kH7Ekkm+UL5+mQx5g4oUqAftvm5BQI440uI0apih2465uT8Zb9UuDwbPT+L0nj9o
f0ByL09u5Z4nrQLBb0ujg0uBbYlZxe8va8RUjyRPUapYmQrGT+oVQDbKGiZn6cg1
B/EdfM1QllZyVuW+/9txorTRU+ZglZyN+xrV2K3w+0YmqqzF4k1sgjo4gJAcfYdE
s10Xpc8QrP7zqUZEqbHmiFOG2rnxdGjHMdTs6HgczgAODzjZQPw0+Qrwt6oUMQHH
J25aVEgNJLje9ql+4jNXv0xXrM0JoBzMV91O5+ktyJbMiLfk53OglnaxuF5MUNVm
vhxm3BZlqURaywSP3OmyxGBdeRbsPse7l41Ixv2mThhdqWqPDxeVf7fhNKmMkRjL
xXdLnVXfkCsGbLR9thRt14CXkK8zZqjREd+gf1OROPkCxM/WbhW9sp16Cmi/ecZN
OjcG5kFx5/XJyyvifHDNIzTfSrp4tulD4joCG/iX8Ie+x+2dqjj9P/qBMhV/UjKU
4XBXXgNg5xVsJiFR2/KIQ5nSEvSYkBPn2h3VpGM3A5FrKy1NYsCwhshW1Ceu5u8e
wofya4VbL3ZBBauo4x68m9kApeuBidljxNyVDxHpz8/1FgojHyN+Oq4FyBD5VAyw
gH148PM+S7jm0NrG8tOXzeYYu+jobkdOpcAAGFs4QOleSPvd981Uc8NwcqGmqIPe
erLbwm8jvo7/dheXMemNcbMj6/J7KtSTKxiEFAOdT09ds4h0fVnvvsix9SprFygV
GUsabqhsjE2UY+TT1GVt+sr8QQz4FnE+gnYA6E7XKA8z+nO/WLDPmpptZp+ge0oH
b5RumFXd6m0XCXZscmJDhweWr+uAcj8XwZ4kg+10z8DoBq+0hYHeNvusjRRxTsGT
ga1GTiONfKGXkulaujZ+5krvVdxrHSUV70X8WYDk+ngDQz9by4+ibkNDgH3fBahm
KubKiolELW3GfZVqIDjpSvxSdZO8cdaX8aqdfv5cQvXQopeP/qrBunefc7oyGnU9
RhGn+bqAHwH6F0rg8YI5hWXxlJ8aAd/iXYWzFOXn5hKE4VUc00dfAtzCfihcMdgw
U1+4HhKBmJOQQRJuEKK/dAQSLobFNx7u2vXBKUEg1bwU69aFKvKD/xp11AqGzM7e
vZNR7tuH7z+jJZN7JJlED5VwqjX1FlkrfWgEU8seBPM9ln2twDI2q2QWK3Clu0MY
6SB4v5wFmi6N2wKUkrF1rzaKvgbk/y+omtznjI53WFEVbssYVXYPdCT/k1jLihBv
JM3Lx3d7Er2Y+ZUSKiVMkBnA0qgB66DfFSRfjxeSxgKtHAekAZfSQDN18P5mKsKC
3iKi9PyDWrHPM+0h+b7AmO+mZx92MTQzcSM5gFlCGFhpRKficnC+WgtnFEzgh7nu
diwtn1KLEiDq/faB3ZkCc3bcY/Ng/fBJ+YaJ5BNPNB4u5wSlHnsa+qKILNwbz1Fl
QWfVFBoVtHF6S4TshvpxigNKtCmF7u/r5p5IN3FZB3774g0O2cP/osiYJ73s/3Hj
hB2nGwmUxmbEXdbHhBm0khPgiu+x3112VZVTw9NsKOLiFhRjk6kS4YTMog6q2UI+
54tYbDnvcmfytwNrB/KZOYZ0+LSmVgFbqcrgQ/QhACH6Qk2MViapE4tiJii4Zu3L
jYItfxyBnK74I+kQlfI3JvFMuY0gvUGTaX+YBQS/Ur31qLSddXhqUKcrPGClZVT4
ATlFqCazNHkXfP3L8bE9feclIOC7nRZMMK+9Sp8ewoKu4OxNGZPmxzajKtdjw4ja
kh/kIFmCdFlg6Zo0ye6aWg06AGF/YT4lGB/YTeftmOwjqRYZkCahO8jfrklUodZB
SeRypVmO2buoOOie1a/oUbTtX1P6kbcFnxm3Slv0gRRXkf/yY0eHMyKbqroLR1vc
n2UgVlb572NnPrcaVi+C9HgOHXRHuH+p/7qlVo9RLaOxxaadUot5Lbi+/Kdaq2SF
fakZ6XRzUzqreaWntaZrPHLc/TgmdYjhvj5UaVumaga6ufxRk8U2woqYJXDF3V8g
Z+SLgz4MUFpS5OTEQIio98Nvdb9SirKcSUcASmD7b0yM6I+4MNwbAfxFRqRNQX7Y
rwaVhsLuIbR5U61Udrly/OvC2v+mYKslg/uYNdJIkhEQZNN9fHWeSO5IKnBfQJ2B
HdoHIBeKhzZVyqX05w5jHG2ttM8lyruddtiMDStDX0YPxNb96PeD5FXRICQNQZT0
TCis67Ocrzm2viSGHWUFs179kRCHMMwrA/x+1Hsu/aPmESNq8CtFtvh1likg3Aky
Vi2brO/6H/WaBCWX/APcopFr/fAeEpiPnWtRIPMpJ9Pn+lIznrYd2xHG2zbVaAHO
Vh8Fq6zzoXZTEyfSakjhFA2G2WRbovv9ac6BeMxn09Iw5L+9pzDJropHwKDLdfvB
OejCaNSKUAqMHF0YqS3rMqEIzWDI32q1kFImo3aEau9CfZX5gh2TRV/pG/HPr9I8
yKOzVwqljVbC2GMfqWCE1a3W3Dq8MJQYRqZtZmP5V38pZUaV/mUe9FmJ3QeQK1Sn
BVCxy4qUsWSfOPVZPeoB1+hxliVgMZHuh9kwtaqCUEfqZ+wBa/b+XMimwrdquAFO
1PL5SxryDC5zfJ5705nAFWs4ppOVd/NDN6L+3/yN70en32mYUdNGv9VBdQxJgTqS
4YI/JXtKnj/QzJNASt9SfwXlsbu1daneSu2NUeiOqP6ruh/jSdfaAXKnHU5Wq3mp
6Of79LxHVpou455z/Kz9Nv4yvB7G5HtQwB9pIc7zh4jr3j728WVX/QjW+IZv7f9n
s+PpVhVA8/CUkSRjyEwkS0VAhqOpsO0yjGzWza4yHOT/7VqJ/3kLg7eyru5evpiA
94OhAPVpjM/tlwzisnhe0h1wJxgCLFTIHpHrBBIB2Yq55jBYBhaS9urR42fhB3QH
X2bnHk3fCVPLJcgat7L16Dsotbf/vFOAYragCIogpxopRegmowPh4v8cp7s8LSut
MEXa6/vq5B1g5cnf/CSonxN3n7SAhOMJz3o4ssWdOKgW7gNwwiMZlO7FWn6yUfyu
7OOPNybzqkUZsGH2EsILZHg7nu/K+/NGwgsqUP4A190ssp3n56a7sDEFvXd+0Xww
WNk3ejlovccAAV0mxmOuyY3tVNuavFkMtWp/MLJhn3YphFZ0TGCmx8H9b8s0jmFx
VL00OzTIC8cSDrnD6r1WJ08Cl0fQB8O/Vx8XB44fhyT4uWA1IISb93j2Kd1CrSG9
gVXUnkHGBXkwIERFj8UA/w7OY4BaHnUkIKILyGcv2xyNEz10td7seTRYM3tYzH5o
38SSqfFAJxh+9kgSFVUuPssOKao1DU2Z5oHHDMIXbI5JdhG2jVcObBFjP7NbYpbb
p/LA8qXEfh50GU5GcPccLs2Iq5WSp6TnWnOPf/Twv9bX30m/zYCIWexh52V9vwE5
SWbBD0gv+Z0/6Bn2ro9t+6HPUKGNCApko5+42c9C8aii2a27DEXNgYcTB2ay9Dg1
rEDPSNP5W1qv+GJ3PRuScgExNQhljzTIvN8Vzum7s0p08yVFBhct5n02nvlXc6yq
nMSGKZQL+2T6uix40FtJPZoalqcVxkWYV3RPIghxphcQsQR3RExWdrT3vOTjUbVt
/YB0v5cnhxu29MmopGvqHvHu9r56yByS1scrQEMYFwgvUrksUKRdUveP7Flo50Z0
5+Q5KQNxOBd4hSQ2vyvI1frRql/bTj1YgGLNUUr45r6HNfZaxpcS8Qwu75UWeRqY
IQDb8koAO3bACtFalGTcAiNidJmb7+BDDiUeGRfW/d77rsedNKq5W9ngKRtizocc
xORq/mTtATpiPwwkiNpULiiINBsKHA49fGZCXe6KRsSZuJTfAmxpxEluX2RtkIBX
ZqWSVIPiJJ9czLQBmSLDSABarscBUjE2CxBNtf61gK8o6zx323pRj1K7LYVuuMF8
Eollf6QQSYomK90/+nEVYCU+0J683DMrRsYYjorNpOFzI9blPp3LOY0zW/ZWYlRI
vkHZdSSVjIwX/TpEiaQUilqFJUXDV/Et9fzSqS4uVTwOAaVGLkhUnJdiM9vJk62S
s5rPfAJjLRap9mAerym+LlmeVotTF42a/+aNZ8y6YNYAbq0cw4e93X1KrSi8AHwj
jWeSFH1Hhwdj2gBEDRWKonTaeXm0/LxnoagJFZp2UDZewR7S7/WUasikpqGO8Q8w
m2sEuha62G2fsQJNYQ+xYs6xzARkrWoWMWFeO+VIlSW5dvJbushHwDJKx/PJ4i55
/lCR7taWKrgH6P4+wHVWdgvWDEIPu3erDLfXByyDaJP3dXt+tnbCM/yWMNt35yLO
uEBvZWlf7XTrTMJqP5BLGtHvhnkn1g8SuPU6ZkDlL6jVNjBT8TEPgN/Kc8jV2hLF
mZT4bBXjhPDLaCIWVNJKSY2JVZMTn9NAxBOdyCi/ZqkY5DG3zgGFwMtIIpxucS0D
nhOmmIqGK+GzTHWojf7VYJcszQoNqSR7y3XVQen23RWdYxZzhxPmyXAoJrNZUOXY
NiL/6PQibDErAgzALqvCFz8n9CJy0d/fBZ/1Mq4le/JC0i1+ipBiFHt9K6mzPR8m
gcEUThdgpkyZP7SOoNLaGxWVN5gcbERRogZCL12ogNiH7h3a1EDD8cjQ0Pra2ky4
r7mJh4hbOMdQqSf0/dQlYjEQYJmB1YtjCH8lYOLkaa/RDQLdwqFK28LDiHfu9V3k
O1LqhV7I5k9ntvijd43SCEZ9Tcl/xW6eH4Gw8hE2K2Gj4j+T0TIiPeXVXlap9X10
3B2oWPwlNgzAWzUHvTG58ahW1sezFtwSr1ofDQqSudSIm1vGrRvmgnmagXOUNjZC
NOa+0TxaZMflp/yLFHENulrQak3TueriOziSzNIwNmZL2LaV2J2Z1BBZ8u9WQz7S
AWsZBH6L+9NNhV6ul7HZyawed+klRHHM/Zoz6zpffwzzuQfaAntmHlHROTbmprog
NErMoX/LzSwYzdkgvoKBGZSxWtBRlyxpq5nNvJaceK0loc2KfqAIk9P61yATARh1
4XAGWy871flIQBmzOZH4BlHBAEGATZRx52YleuxA0XsQJGUBc8zva4JSvMm4ErJt
CUJBuTICrxtiyuWxUzPbjwZ1AKcTF2jn2LoM6iX844AVGuL97nZs0w3zUZJjWf7j
6o7FcVemxDfDMaYpcB5V/XsdqJaZpvzaVHaNHx1SBB8+GYAgESn/JmkbACMu3XaM
xULk24wxy/nyc3g30zgiGTfq9QjEx8nv2hHzmqeb9/iUYCyXODgIJ4IrsJuGA9nH
bxFt55vrmGVc3krl4UtUbSe/X81TyCzUPxGGquDHSsWyKd/hwYZ6maZ+8ukUU8e6
HSJm1o0xem+b17aDghPX0yhymCcgDVZg0sDvy22xfAoQXrd8Bd37UJ65PZLd2Z3N
uAW1RoB3WRdZWrLjCt1LhwRDHbHuf+kyOurl3X1XETGQNCjmZaRc85AHnvcTtfMe
EYRVbTu/FNtBX78gMsfpd7+r1UGGHezcvgixDOoWheNKuQ1bo7ydxpIDR+xG/a6x
3nBcAMipDX+AOR47qeCPcjYBJ3u4uHUxa0iw5QqnKyQvoS6u4DTSQzNKBtaPKib5
5PZJ5hOoItDSgnIMTjQXsOtifqNpNKrTPwFY904Bqbt+WoJPJm/oyaKf44JXCCg4
W7lxy7gkdOHAOxID87KdJ2fJFqwuFPbxulSBFpSew2W/uBpBOqokd9Nul8fpnnPI
zLKZ8EwTOV4tWAAgbHgl1ZHqHQtxfd4Xs5/f4pccYqZH3qyh+mDwOp0ZG1i60SXR
rSsaPmNpjVnTME4UPQn+9Pcmd2/1c65xie/rNHuDkmTTReqz2zmDJGcB9PZZwXzd
/g5NxbHT9Z9r6OjFRm5ZiCe+Zb0l8NLdZT9ERopv95EOAYFIdMhQCPuQFlSMk1S1
AaMKSutho/YWguUPqHLOHX9Xt0EF+inUO2rSwiQRBhBvPSvfRYYtNOClfC5QV/su
ZokKLWHzVtnKMLs8/utJOWLSRJVN4Jg+cgJ8WZvqY4owUsnP9DHCsprgyunLhAQV
ZP8YP/VvlczXs/suFaYCyowyLcIm+8ivb6AvPnocdhKaL/rcek2/PbBGpOgvCtQO
5QKGIQYI3IiapJlxvROaGcCMPyto5YDaOrVRTVMxVoINb/Ko8iHnQ3TqRjLfHYSJ
A1WeCaHTeu05zbwVZeInPuncDcxkd+z9o8i0TlLN7yfj0g/lfFPpGBptvodosU/Z
YkzgBYVuNs1I9UPsgtHHn+V7e9/xKRCag09a6kpmKz14YpHS93COSPDIOnOoVcot
RYVI4vnxeeGI/3EYzhw6AgnjQhYEPDP/PSZPtwZ5+Skvpi/UXJlshEi0pfjS/prH
+RxHTgeJLhXRm8Ym/afipMCQps3IGBSRfWBU6U28KQiVN2jRywAQCfPELoVF1kjD
tMyE9VF9bqujo8Ln0tgq01yuIV8vYi+24xiWqBWyAa930X5G7w1KeUyQPUNMNz23
STFXG/fL67Dcs0+i3hSmP38N1vL91fT0mCxjEv7X2rocC1D9HTkZm2PX6IJ6bq4u
AX5o4H7Y5xxXbungYkIr3U+0sp5GhdKh2ZQSkJph9Wbn2A+jgGMS0ygpM0ke3cVo
2pklHM/r8RW6y+WXBnfflweAj9vUoHu0t9zcbVLnsv+v9dhyIVjrn0fqLCk8KIF1
DAyKaCICdAR4xiNDqTkaiIK0Rena2ZSLRd8QnkN8yGLFY52itI8ES7b3Fl0o1gcD
nXWR3bDD0kpgNzgWPFN1Kj+Dy0UahxJ5yL9Yk97e2CH+HUOfnev6/KCQrXQ5Luqu
I1XIy3Uyo1Q4dj3zFiAYrZB2syNHQCXjBMzjsloBmgPNmP4xWJ/fNMCHxRDsWFJa
Bq3CWTiJgq/UcuXLFdExPHi6df9tu5WtCajPcX1Bceht6AUL32kaa+i4dPmWY3io
cwTL0CQCo5T21CvE1qzT8Kf1su2EJMhfd3uBPnYOQ21hSCbvDJO5lgpzOiFXTKTb
iXdk1KvLLINTfCIWG4NDm2JOU68HGcmPrYnvHfw6btAjK2oocaltjBq+t3NCIEmA
PKikXXOZJMxqqha9aukDWHFFGt6SspNA8AiOVBEkZAIxzFxhiBwnYqAkOsYNtlQl
7daoQo9ft+BhXIM/Z9LqoYDgdDeDYyubDC80935TO3NMMliYjEMmo3B5J+zIE+Xd
axzA+K05acYUVWa9fwAOssZVjkAnQW34Uq+06gfcE4GjYWdGAJwSDIXIKgnd8USj
EDGlds087F0P/Z9NO7AXpmfeUzaNllRzBhyaqCYcX+7MUPbmFjDmRcwSPZJGqAwO
aarRnzd5+0jDmAuhfRlUebUTBBsyM7nNkqGG6bbEoBfmP2LZ6kQVNyLp3JQLNh6f
g0nlxd8iw55/L5wrU8l2PXu4TGcJTLky6+gPFs3vjw92vXaaBvA0A7Qrn4Hv8x+b
B9+E+yARbZFw492XgJF1NSYsTgdoofJIWE6RiGzBbYWMxQookbg31sziaO01hGde
MeIzvALPTQx77AKo3RjVSgN7qDItqM8fRuUEGRl0w7PKfIaSvphl7HJS87YGSc2c
JgVDF6qWmE8y/5aJOHYciP/IW+6BmRgVk3TuSwDDhYYkyKsLZfZ+H385stj7l4fE
TjsHndhRfOI3LFTd5d30ppxoVLqOk/QlA1J0iwt04cexjhBAtc79tjCk06fngZYT
pYtimikJwv1YXy3hfeZxC0+D2zt48QzjAdMlhtRK2nbsXe5bqJw+K+68uIdT5k6v
B9te2ilFnhzw2fLG15eSP9Qyt5hozR+A6QixczlAeRDr3i9+W2rRUL+04hwi3IMN
OrJS275bmB1cBNEECZoMNW0oTLsU3gJE1ssq6EWAIjDLSGPnJodoLUshlh3+3ws+
Y5k2y+3BHXFrSDcmV63nAIl3IyfWOb9CJEdyFIxcySYtabgn4W2DHwLamudZGzlX
dr/Vo4G7Ho8PMPZeSJThb10CkwfBEYPYcKdy3v83MCCMgg1rT1UzbF7U6jf8hEgI
jamyqBK6WftZD+38HmwqkJtKhNn3V6kAWruTFjcWI+0iC6INUEE9v/bliedPKkHj
+2rXvE4t2TDpwkGFPj2T9AEFR40X+268M9T7FtPB3MZnMSpovYDJgOTdZ4NzrDAg
eOSCQFbO2jkKVnCllMVI5YuyGArbNPgI7E/mHkKnNvxKGF95Ym7D+f5m+9nURr6c
wCBpfOihBzFjYNWKtM4em4smGa1oUk5wCxRrxhnvKLKzkzvuA4TxuWyoGTx8WaZU
2uHF1JXVGoKKSiiqAZ5A2/voeKJW1Bzv6La1mAmFvNtF9HdvqNFTUGIF9Q7M7oHu
a7NMT/nkRmsNMxz5gZzqY6mTVYHtoOSW8MF2zOq9ewSqhAGsCWJ48ezJVsSBej8M
TdpiBvYEl5oX2/Vf/PWUfu7U5GTCBKKwqAtsJJb6urlqfSEG/0NLG/BGeYuGmeDO
t1KncAIRJvVHxig9xnggHOooG3blV3i9HY/xlM51CpipgKcUmMQIm15B0LxX4L5W
2QleJ2FlAXhexIoUSyrcbZSqkdSS9Pd62Zasbmx5sGoI3Z63N9moHzt6GGfMXPmj
Le7BgxyzP3uKGxwQzOt6LN4p4TPgkRG+fRrSoF0Pc/Pw48at3KWSHUqfeVr8NcAw
qFHsNsbgoYya6B96q373/lyuF0WX+wxwP+zJdLPTaj/+kVU7KAmfglueYZi9VGmu
MATEh4M1ZAX8amo996QU8dqDue1HAroNoxHH//fSFjLSMMynkXvvCxQE/Yx6FUZS
n/oSKsSszo9wFSs+2R84nwNpU9Qa/XyX0/hUmm934hfutCI5pZXLR9F0GyJ+PIqy
uZHv/LNWoVuR/fESaE5b6puT6E91ObApxTVLN6Jhs6kjWx3hujfCbIkB2vzjxBZd
1CqzBpqm/AthRUqbXMYX5VVR6A+B/Ptgmwq6tSlQkb2T5L0r/05g2ten03YmBuTt
HuyuG6Nwn4aYa20/I9cgPVAtLeQymZ7w4L5GZtXorrL4cCnQdLwrkS8fFygb4j+X
JIRrn7BfqfJfmq1aXQgZmAiV/iy6vUty1nAJpQ530vwy0AN/v1sQn7w24zoRTcOc
4QSEP8x08Juu2OFwjLFbCqek29pG/p4UdDmpAreWceIfNI4OP5fE6bXegLuWfd29
b9UEBHGv9mt/LN+4ZEMTUSKqyYxeELy0gu7W7d/aLx4Urfs5Zxsg3slITYFe4oOX
GGEQkbLlSzdUGcplXMrwb7QYkts23OAyw8b8cpzlqt07eyr/pKheJhYt+X2fHEQY
HQD22+mq7rESqVTBj99tk4TFvhU81YNQOygxxDA7/VJihNhWQd90IJVGJrP6s9ls
hucxahoM35CmCZs+uWd9UO0+wRz7xJUm0Qsp9E/nzxAO+1qu26fievB4Bln2kt76
xbqA+ZCbAxUnbTZbs6XcGUc4+n21/Gdedtji6UCjP9jzulnpnBFM3dM3i6fMEZ0y
py/i+Jq+ViZM87poVSvoXru5ciIZye6Zd4L7Fh7ODf8duDcv45yZoSuy+StTkqML
iwgCPld/HHD7QFDDQSX/a1tVWyr7n4rCFoyz8T+2iRnEU2KERo6/nOSGJMVr1IhH
ILpvb9NLKuIq3PzWaCLHcrqZif4+IAVx0s2AfxCivzLc21mb13oKDDHZZU+Lb9qk
5TeXGjY1uHkHXF8Y90cdcei24lsUh3V3ew3E4Zqnr/i+KOLASkuQrWo0dVISajWl
cnWZIfqfZNGRpHiTgQV27vqI6XtnDEqJGzbjutx57KkPSAa3LsCPdD+OvEO4qEYR
tGnxgTJZIw4o9GxFPV5zuHwWirmoLWCg/JRQdeSBZvUYuOZIDD15PsCBaVCm0OmL
bdblm7SJeMz+65zq/rXY2/w3usoW9NMHGkY6t9PzbwyWlgN0hK2LvSM9uJDOz4sF
LrIz3qPW0cP8+o35UzFsLQAg3Tm1hrxCLXec+5xtGsMX3XBY20K8yL80HFRjF1hm
9hZJkb+pLrqzGsArdYj64GVExtXKRaJHUmi9bjd40g55K0c5QAyQSMj4wvCjQ4Eo
c/YjrxjnMbMQCKsXoinWgLQETA8NVn7nMQRANUohKkdBGv2Evuawkg3P4RFtEY3C
oImtsIuHnEKwZnVhB/Q8vbJ6S/LS8YaSwafLV5MCcMG8YBTaOIGfbB8fGwVDJJHJ
EWeg4bNvvIeDteJgV5m/WMXPJtf/xaMNFQITnLTKUPYPGbBqPEHE5qgk1ywDG0K+
XDh5dbSAdCb/6SZz5k16MK6KTwIK6Y/fTgxzUMdM+S/6jKElq+laVSWr37iQ2TmC
tvPqEVS4fidhUEHa5nUOc5L8/lJ8BIAg+Sd8TBB4qFFtDE7NniVKeBSeOwBugQq+
j68TC+5ZrF3V96wL+QewWmXxobCReVM0+FEUkGDrYlXIuZl5saSov1ffklHAv8FR
HTXmxUABeFUj9KdxeMVBbZSADoZMDJ9H1RhPM9EbtXToYnRcYqvpRtAMX+u4HyO9
StIU8gvSyGaSkP+K8XKkKyywhdGnHAEghTIjI5sHwy+IWNPLZ2aBuj4iPdrcNx0h
Xse9o+xGXTiV7yP+u5O9Zxjb/C573lV04c39Ig5BXSxt5kN3CQ3hXQt6vsNeje/j
110MhKURrZgtYTtHoQM8ZQi7FuT5OZHuPjbg1QAA0b/Bnrq4aUNGneVX8FX8v+BA
QM+N0KWJ11TkDcMjA4l8EqOl+Kql3WTDD+aX96/hnPWpGA1uEpARy0JK4e2fLpf0
bX3tQyBtbE1vOV5IlrE5RZVgxWRcAFZ/JpTEgGlz/p+f/IBLnkPRFHA9AG0UiHKv
opCQ2Na6fGWSMDnExjBnnPFlBkG700XswYRPbc/Fv4IqNOWe++siCgq3r5Xht48/
glT8Bt7mc7HT9I7bouUPMozdDqe1AZJq6ltmT17PpRvwoPe90ufNn+iWZTcaBsMO
g37bDnZMMcgiz47BfA5BqVaPq8WGXVLIiE9oq55VNHOFOQEjLsZ6O83JnXBhNb1N
CBz1WXg7SKylPspwVrbGq8IPFTTG8w3ho4NE2ErXAYjfsnzsfrzbdzkoyigUypXn
bVEQ/aOxQ3/AJuyr273K3g8BNs6owrlPKui29Q8b0+tBT76gk7v2ibloXREmrf7E
fjfFHHS4NEFi/yjG/3lRe4EmR8u43RJh6Oje2dk/5aI4Viza6D57UYsceZzGCXnY
2qoUDqIeVqyUR017/dGY1c41+CtUk2ubBZpdFjxcLufW1SYVfIftDjFltiuh8jz3
hf4TdkUYIS7M1nITxYXVI8GCjLPhZrj13WpzAkIxHPB4+VDdNRVH56mTXkkYRLMC
zHa9GnBmHUsbKvs8h7F9KQ3MGzBfOm/nuh1a1tsNVs3MTHZfjUjWITXM6Uc9I4cS
FEOqVZrPoaGh2VhxShodPwXcsU8Uudb0l+0eS9hfIeRN1rxKvwxG0nNZW5XPFQt1
0zA7spU49MgKyoaeaUvigjAtsamPDlYitOK9EYexsS9nSJMviIRsI1+mzJ7rlU0L
/BRAav7h1KVJmfeKlS2MUx0VhKPtbo8E4vx4oqpw9R94sn3GDbx4WOHCQBExnl8T
uHUE6CDG1f4mjJaQXz8fYIk5y3sT2OAvr98Jd+ucYzpTWwKM6mjpBk7O3e/Yi+Uu
nGP0a8JE5ZfeOuM27LH91+zB4LugfWTCqJCt6JV8ZsA8zVIJlVEzKje7iblE7XzO
qgOXNcXEaf8pGlww9VzgwPW6+fZQAsSXfnOy6bw6i+eGAcCWUBZjiKlm8ffiZOck
ZWgg1vO69C1W4Ed3UyUQ4YwKXMD5k2EaQ+6hc5bU4P4B1eo6Ct1cKHxKBmDewhv/
5XSjHJLjSexRSLQJK4OC6/nB30RJAogGhGYZJlq7xXZBOaQtgGW5alnPeks3AbjR
EMq8JfdBqOhjXUuL3SsY2Ys2TECfoEwbuLh4C6FrA390rnqOSAh0L8WsFQuZaAcp
1OdSAv97WDQkhhe7aIUTjosNvCZ9vF6J96ZcKJZbpqaR7Tnz5ksL0+b3IllZqOxA
jrMe5Uvsukzi3AzBmZbT5wM6ZWj9T//p/k3Y/L6dFni1Tg9L4RDq1iH8qavwughf
0KUDHrZByEU3eG08OT7nisB9SibjAGe91k0bEtmMzspV2Vo1Qh4iCSViFhrFH32B
6qcl3iludHBpCFAjMEoNK126/4PSvhM+CGpuWXHn6wlHcOM8ue8nh/MQm6SZjpBd
a2POUMd8qDC9t/A/EUYyFOz6/BNpm7YviaWXGWxznv5zL1KwB1+xI1NGts1LNsQD
aUrNoqNnXTcVxZ0A6T08/5JyTWSi8AgWDTROxAf/l2fdcNPAM3+LhyK7UH0ccDm7
1P7l5NQtcWMr8RrOaOfE9kJ9D5SZ64ZDbqhMlpE+E6FBfnqxPNpyyfA0HLZQFbKA
PlgdJQL0rWr8gb6mOePLHlzHx7iie01GrzkKPJrZD52xFb11qc6zEWOVjoryVZCw
ImTOjkleiimYK6VMnfHMA2lguziYIVTmzK7xiDyuRr0Q+LMmiInyVKwxsZ9zi61R
ELt7v+VbpReWX/s45s+MhZv48RP9JMF3bzK5rCNepxRjyEFyAkCEtcvR4h8CMPsY
06j/PTPuCL+WuXWn+EAp6gMCL8SuyhKXIF0MdldLHMmaal1SBxuwQXS0xGQOH2ZQ
mInwD6iq+OsDngabtULy0ccb0LvKJtvock8Csecx4QAPWvyRxgCCgVBfhAJ/w2kG
T8FeNbqNF0vZXXhvGZodCq3KWBlbvoK1gNO2F8vkrwBJHbjGmzXR8E5j+oI5w+7h
pwv7t5gJkM8w1JeNbx813pzweEGUq+ByehvAL4NrorkWEeQwNlv+qsGK3qZjHANY
3efg64jAZSIP3+dEl8oQXUCqgoiBiYwDzZtKtc9MzyV9OKwyXF6t4ulv82CN802Z
4fns7tBPofKjePqeOAOIjSPddPq2jV7KN99FXHdoTUqnZ7hMPmTlVRNA8g8bQJ55
sVchcPqCVsdFNm8cHXUGlRsaBOXSOVQaq+qdTBZGZuK7st5Ot0Q6tlhC0MtV7drE
mzXuN28nQWaW7845QBuXTcPGHhGxORFkzCUlroQG/yLcHTrMDcRp/TpaOd479uNO
bEZZL1w7h+rnbk407QepOXAGQgkj96q8buzSfOd3fncvqrr7flaf+mp0mLOdtRrB
/jmdz07EHuSBZ+fyh3kC/okHr5YRlFdvLDNtMGTm4y+bCrGDqR6Koe5aQExHh9l4
EBc9BNAkTjSrhtpk+fOtVC8PXBVHSL79wbqpnVzIo2iHcQesbFW+G7tJp/zsFFLW
v0olbIZZCu9MqR3TNJ7+uLYbi0ROH2bKCP+dmz9E4rIH6AYOLuG1wFCQUiIdsr5O
2+f7WXXwVxI+BG/hmFTixS73OWiv2xHUnOxIy/sTqSLyMhVS0mlNJTYXBRjfoR5L
Orze/spBvwa0ZPUxRnScRM+K/y3aE65cysZhTLnNjBm4Gubpaa5ShzGNpEAkErwM
ypSsXMHToU3HQlzgwu/7k1F59qMiTipfzRFjUT5JhgQJbrZ1wmIEK5izDPtgvlW2
D28f8ZopJY27vAkmX8ferSBc3Ch10LqNWVFhDY3j60e9V92Phs5hhEVeYMjTCWCf
+Sd7XjqDqmWGXLF0DJi9QB8Ln4Ybo19sGBUoOiySKVCCriLvN6svb1UmRX8SorOl
m3rToB6OpcxxqKaiZ270QuhK9gUDVcfmbAI94uoBX4PZOleXJpX+yOKzJY6Qh+19
SKyes65RGuf5jfZen75IYHJHn8PL0X6AORkAUbWMXz6hHSwPiNdOYK0V+pDF2hgT
zO36sG3fhjSwuG1UYymbpjdNFG5UlyjLTfSIEiUekejOJTFmYmYvGPEh7Ovo1sMV
BTzmxnNvlBxOTjzGIm3DJjzTybQUTSg+qi5D/N5ms2oGPh9D2AO5NedwJg7ZFliC
LFDO/zVPQgVI1NWYXV4irxhtfx4kMJysRgtFsxZq34xJjc7bTUzI3TccUF4PuxEk
66gWHoSJzwIiOuVBKCJ45AzXPmbJhkoP81rxYbgeWkDKu/aHgsgar4wmhsHJQ1ui
q/otyfrBguH65NRc8yUFHai6ZNLTKrvy5wfs5fj5WkOghY/wKRJkZtdAaGZH9nHa
JOQVo7sRbLADgCd2hDK4gSH1NO4lMWW2ZVMj+afK8uBi41x3W857bJxQ733NGpRY
Gi1AbhVFS23saTlLulLS6PCoecd7NBdrRD5EPdPkeqXP5Laka2BaWdOxildP7b20
jmjnR04u1yMRe3acAiEBPDKcIF/BtqUsuV6I199Rj+Tn6VI30PKwf2k4WrxM0CbK
TfpalsHc6Lag9CWXU2frawYjAWEKxSt/fgpqI+RuSotWpFxvQ8xcGh2ZnXQ/OaOI
oOiOR5ln1OdONnogbaDyNqd1iSpS1nQff7SD4X2Wd0Tat0YV5E+xd6NvGy370jUK
wYKKlJzWxz9e98Dh2b+QI0fAmOfiTzibPRVVuSbcAHApQqb8+yHWCNEZqTuNMyLX
322398lUBV8eO3dQ7ZX4aic/TDvf3dXje5debvsYcEBZsn/KNI9pYZSiB22bjmZM
81wHXjEAxqFeHRmACU8Ncb0e8+5kNsUgEdzD0KBxY91ysDCqqhaPGbYqWocIPrAv
Tqwhv+Xppkmv/91XJf8hgWoiqNFKuFvjLOSMef5sWzp+RIIJ3Zefj51p913ZIId1
PC0nNgiMOOw0Nu79ZJfCviNNnwnfB01o2CFmWPkZd8flIxVGJ03EHURmZZ6ZE8Dz
XAEqbPR6rf+lnjoYicgFBUySahxaKO9TzaSPWfN421edLhaj2gje4tulLQh1lnc/
OVN+ZjqzbU6mMJW5HFwfHh5XK09Xe/f1apcIN1tzw8yWFdsgI5owbnWoDS4jox61
DV5ACL+GK178r84+eJgDaZgZ9BeatXEg05ewXYZ8tUfT8CfYBkyVEysP4q1XBN1a
EbA2kq8ViUvuvibO9RFP5p6r4grcdoznYSLA6iB8V3ih9hU7w7h+k8vEoY8KSk23
ivXtdvs2Cb9aH2tx4xqnJDHuD7D9TziiGRoCHyPX8+yz/+QQPEKQQ/uF15gK+ttT
uL20XXmaujHgNFJjNRvfXDfKooexwwqVGhzPIhxlBNeRJ7FzT9IVmy3VxvcGbkGv
bJgp/DaY4Kox+cj/rCYZJhPO8othhav1LEwce4S25HTQ3Z9oGiMUwFO7R0o32iCg
8BrCBR2TIvrLlmP0lZEJ6cGBl5968kt0CjE7RuqCAWnZew7FtOuklG3xuvJX3oZB
XcB7c6tYg3XAwaorMUDmBsTK9Du8ysXIndzqZAR3qtl4Rtdc58GPV7Oxin9HBr9H
wrvRl4GKDnwI4igRvgzHxZVZtOAWu+iR5h1KMJ02rrTMLW0T81CaS7+ULZn1QrSp
9e/VLJ4khn3cyZCDC28iCyh1oG9nWgCD32phloE/7rBJ0uTvllNauSFoLkOi3/TJ
VJaGyHS5lS4aaiPTmZHfD4ex/6uWnFNK8+ctPvPcJjJ7RrTRBbd3XzwQWqQ76ulk
zYVZkUcrwH5UD2h55jfvDHaFGdYX1LHLhM5AN6PKDeX7ftYKvHglWD/Pv6Hnn46I
Si8QTrxn3vjWx9fyxStsUYmAzV+cNZxkBNE49OpHqYUyRuT0FhflbvtQOQTWHoNJ
z8euTDBpem8NWX5V8mCRb9lOPgz+jHmZS5Qji1Jg9DFt3Qb9quMzLFc9mNKCNxnc
3ExdiE0cjxOxBbeAKBCFSzx133LKy+42AJ0HUCQn9n3bz/YP7EwbnZ4MLzTHOOFX
YXEbZw1YWnHRVGDo1aYbTTIx4kTD+4eN8/NyzRrhhaSrCrS+hRGRBV0fPKRpHpbb
7zgx4IpSILL4hH34FPsy2WspCbOhAE9Xxld/1gFFxY7TGjWnweB6IoqjS0Xxqd+H
l3Ilqeyos3VwSpVqavG3Dwf4HxhkajsJDy/JE4FKRWnMYHpIkBP+UhH5JqEpnnsw
3PiVtQjOR2NxpM7O/86Lx1f/q6fnqvhaltbn8FP2Sgv8WMoKMHLZAYdG3oEygzDN
g9Sf/+dO0hnyAu+HpE7Gj6OEe1OeLpf/EdbUFewQBTeN5ZUplVlERmFmGPWc9taP
knoQEZdlGWLMkBzh7kSoaMbRfI68v++WKgZ9url1oa5Jpu8OmWnR7zK2jEKijvpi
rjP7QZL++OaTiIBsoHahztAxPUKRdpVF2aAPi4Fty71YRnDbzM1OoLX3e1z9SVHO
ADMYbs9z9s8DNQAeA34X69LCnirH0M6oEXND2dnM9+8sMHcRyzkMIP2rUWzDVYxq
2PpGYb6nY609CTJI859bPAudhYLqj52x0U3lr4U770DjlZpIM8tplAkfo4M85qRU
mtuIapTEV1S9Ca7ijGjkWMEbmyir1innnPiICmo0OXUTgWSpbek8FXxTqNiU0VcH
FLgnk406tPV8k3ighto7XtUWzJECyWw2hjUTgr4/6dfUQu5nk+VmBR1/cgQZQkH8
BYpXGYOT6IaHRCnJjRs71BiLwqMSNJNWfefbyBpcCNJIsSi6rE1aSvEHVhd+EGeK
eEyiOtciEB3Ic2WyORDE880eMRIep0b88sdCsApGIJ7Q09e9otiXpKmzOEIKVgwi
SEnWFeAS2Jr5Km3zDxNk0lxrsY/FTjmLbUYUeslBgy7hW4o4GUMc4Y/SF5NCtd3k
qhs5fTk+c055H8OmuhqqsTFo040HU9YPfIRKP4r2ajKyv7upMR+9gj47qQ6W6cnQ
LUN3t8XCF9r6sLc7xv+iilZbgBK2bScJJlY2+SmLSg0BDW1k0e9cap7E5yrpTMSO
jU06j+9TesRhbRtPBeRIkPvyZPnivZEKY5SmPIIdNVxj6ZPqMWYdLsbRN5pYJcjw
ydujhWubCjhU4RayKt/Ym03m+lkQoEBaY2wpMvKl6shDMP9M0beNLniZRGSQbyJc
/HQgOP8ogF9NPl83xjFRkmBQmTmMlW5lBeXoz5y0QJYBrYBnIo5jKsesABUxcNsY
lAvbgI5jc61iTg0v5bq5FKbl1+slJVDxEV12Cz1jxFT0T+USx/FUl8iKkrg04lI4
vL7PrUUaYduYpdFDFn2kWha/mnfb5ENtCUjeK8Hm2KYdcDWdtvB96b9xGkij9M/g
4zrcMerQSVawSynnuhf5t53IpZri0kEEHzyf68ngtRzjUBKQSvWKjpPgL+MqZQ15
hFDzeH6fIWFi6FE8XnYso0jD9KodkSsL/LhIihHtCoS+QqE2p0wKuZSbptN/I3zT
XPuG+fwSTnsRm0bEU/vS5Po8x7SZghJ0aPVtSN3UIZbEoV7c7mbFJBnRSnWGwZqp
E5TQ74HMQ32oinC5qgUaZg54F5kPkEvfzXf331ijsWZ1Cj5aK2c180s0n9gOWzzL
1ozfsPt5MhNEB3JkqqGQxE80aZTZ1O/nOt6O4ws1BBuUEIMNvlzk6bXTV8agnC3n
FpCjCNe6RZN4AaDNXfpcDX1vA6EYzAw6huCwOyPM1Wom1+nga+B1Qg90INJfmWqR
GeJyqrz4aBz6/wAvpcJwqySMQjl+g2/loRlvNTiku4yuKEbXsD8rY557dz86Pfdp
58Flr4VwMOCKXJm4AGiFeP0jio+sKJmziSxb8C8aLQWueo7uoIbT9ZRaJeofiwBC
YO7tF1XNVKhj8tsdtHy22qwm0oza/MM/lZqrHrotvodSThYAZsFLVQ10FgiqDU+K
UZqd6DSBZAlaMorUb2UbgYp7vLKWD/X/URbAq6tp2RYznSFVJXLxV4qOyMz7qPsV
1XvqZ7w4OADqy+p8ruYcgrdyPJdGzbIDTuCNwhsf45MyJAAx8aV+KOh3LMeHEAdJ
oOhNSwpQIRfTM/yZ4JctRVoHv20gr5nAyEMunKqzFf9/HHpp17GWpKy3LAGdtJ7h
uLpf3AO7gPoPuLTMYHrtW66y9mKrapy2lZYWflQOiaSJSS4SKqrEmsFce6/ASFqm
+FPqF/z/w/aqDkEfuEBx0mRuaOJQJgP5UqOfgNsQ5KA5+aG4ljNg4xzdi/fsV7XQ
okTpOiAxzmpbNs/G7rkAgAMdVQaQfxxLPuYVi6Xm/o1l7TPeHRGTfTDKCJW1D7rF
MYACB5nwynMXtnSCOWrIdlBxRXI2lMSGMnx1BpSobYk++q4LCDJuZag3cZM8ke9A
cIhnEViHjkUA7LCpGIROeqfrYGDKAXB6dUgHlr8zo2VD/zmbrNsEhHz7VhRsoVtS
NLMM37V2ua8ZiHkVDko4NnxpqXbhhgw7tRRZFuVCNigM6pwDhjkvvae8nVBaiBF2
Z/Z+KAJvfdUvPFCIgFawUtkxkSGx9w4k2ej3+eKmKHwgMwb36pjh7FsL2JBQzCN1
gVcv8RfxeFYpdWe5tvGzBrhsi6PSFGiuKRSChE+uYUPOVenkievCLUj8JERA3PBX
LD3FHa4Yu0gLh6bDEUiED/hjPddav48/P2Q//TKTjixXLHoqkrQlomIjb0LJ+g9e
5Nf1n3HyLeLTL4NywL6h+jyyvSgTJxmpKEdoswVDsSokLvwtA9V5RM72kbHrFsq3
W9RUZAobCP638+uXn5G953bn9prIQ07wsUhhlzD1qE+q3eLgDe+aDoH5/VbRshEs
5ej7H+Amtvk38QHTxBXfeoo5EHAmylDXLyBntU9N6yl9SzZ6CyZm/AYa//9RgvO6
vJ/WLuYDxSuRMt2Qj+tI+btwcVTfIum1ylXzhcjkNrKceEeZxHGqtSmSG87fcIT0
ZOCc9rGT8np4Q5+EI/9eDSz71u1JeVl5XDhP6rNvYrGClMeG35J/+ZeJa0abOLId
0YmIBDZhsnLVBL62cT5JnJAN6x9E+TZ89n0RZLBZcUOWqSKaviy6hIrFhcEx0PDJ
B30NqqyBaJFEZBDpLF7yVobWlyYY7NpqiMvlOhbpr/oXhHSNyh+KrI4szgC1frev
/UW1zEUVqgvfi9lCu2hijm1rCZQ1mnfHulaqTd2si7GS8LOTAnoGEfQy3CjmL2IR
4Is/93EAZ9lY5xEMWABXbtXjL/L+jo47tK7h+nNcAN+3cpTyBFqCCBQ0GJmaFSEN
yS7fhJY9TDNlhWUJyVfUk5J3SgOYGiyBo48utudQeoC7a1ILvxnXCYX0RGCoPgFH
kk6tqI9+6KxA9CclOy2oWQ8Qv9CUJyM2FAldpiSUcYUJ92lHJ5pNGCn4XAjxDoax
BLL+Zftt01Un/daLF1ssc1BrMQdx2ZNPC3wNI+3FUsi01UYBKkUVyu+9qAZsw/nb
zvb96MrCmLA9pIcvFbHpdyLSCzNKA5cyBr7hlU++I+D1Q0YPsUMdOSER/yohlC1K
oUgsvXb3IK6Ujj1N8MHpQ/AfcCa0AbngO8bVFV/2yzSynfP9FBxde8Q0TmmbqdVu
CblLfRrSEGxdm2+CRGTHXS2j1M/A6r164B6a7d+jluXnoqO3gQqs/oBR4spRBqcB
OwYfj0BB5vhe8+bq8EJXUKFBqMqng3T+e7shIHPMo4f06mLElBCYGSQ7tnoREl1l
xaLlSAQIGLo+oy3l5BV9orlPc6ntvyRlZAbAR2SepSa+wUUZS6xB/NXR+hZKm1lM
OWu89l/JdPdvatpAZKmlI1xxiYVUxnKgH2+3yLkpszoARZcQNLw2McjvyCXM7H6k
7oO6m2+upVMxsb3fOicNu+Awb7iTrakKkjCSx3bfwGwIDcBDv362NXEdUhly24eZ
Yytm82E74z0sf+ny1cUTlsH+jMIGp0FukDwQ6Dehm2tti6EfGyYbgwE2r/CgHg8A
GWhrDLajk+QkPlfRLYDzKH50x9leX2vcMx/HldgLB8lpmiv78ycLlSM6HgOfIHs2
FxaIhJiCHcc6w1ArG+4C0/lRWORbTqz4EPQUajdfWvJoJWW5BkYhsgzwN+RbrswV
HZ7ywTX1dYMViglD9cGI2e46Twno6MS2prelebkPKnxIxHkXj/7ktAr6w0BFdFcU
DEncqt0kuksK09tJirK2Fw3rNE7Xigy6rOalaOmNIUiKZkHZW4AhLbXzTmeSAZEp
fYypj/LiOGxfBKz41IPcLndMlyyWCNbg1uMW5/95A52PkEbWrGY74KKmXJU51sIY
8slgSh2QpkBolkLf6mP6l9T/Z5jyeehFAGVTUBBAv0JzjBbHZAA7lrP1bpB7rkM5
uSAS4UkymWUnxj3epzlr8Z1KtoeNKnJIw62ZsizR97e5W/qGHQjmGKEc84Nnq8mU
813eZBPUfcDfmzfJH5/RYfaKN+f5Te88YTx5L4rb2Ayz71ZAQK06EKz+Bk/tvsEJ
20wDyA5aJxNMWsarLqYTcS5zTmk/k/UnNclZ2n4USLPlIP73ld+m1MyIKWWEEQNZ
RJ8HkzQhMPpSkl0GVq6GMKSTo+ZhBRvuLJQrNXDwOXkVtBbJ71EhVId1fPI+wFmk
1al1JeDkOK7yKeCZVfpL+WzeTiADAaEH0gsNuQnRBVS6UD2M/VftEyCPDOwD9ZVx
qflvp3l18KAB2TV55DgVNK0kRijgAUR6FZFvCqFZNB8t3E0ixGO/Y2OsJaeeZBuW
1A7q2RZo0TtPFHauX1S5tIA0I1I88OxrswzWGiTwEc8b6ewy8ly2HJ9EyuOrwP5k
N9OmmiXCFGplvWjIfx7EnhDpzs4wLD9OFuPd4OJHqqyfFGD0NnIy6apYO2RSJyMe
lPLubd0QPYHFS6yKyRYosk4z93lpNeTYYE1BvKUKh8yvx0HaXgCxGbTkq4BnvZOV
QFDlVIXUrdOyhXE7llGLGrR2Dd0vRRkk1GBz9Vk5F/rcEuHv7iB4HHQzVkL5DO/U
1mHb8MMNSt6ePTwfN+UJKmHto9hoVl3dKfqXdVnkaLBWPD0BUW8AVhLmJINV21Hj
RvsyMQb89GGpOA46Hlco2Qd1IelmK8Fg+jlgjQRhiGN2gusZoZOWgWHGpZhGsIfL
Tb0fP33WDXKTY+pLTBzUk1uk0Abq5u0x7H1veCPqH70JU/ETRiUxiV9PGi6yt3p8
mDmyvgiO90pdfQ1FBWFXPfgdsKhf0VYlZATVeixXiqXn1gTdNl4+XgSmWQ/Zj0/i
wbbpPmciW+DJ6okuFu1tJR1d7ucg3ZcZbu/LS+CttSunsIhnXuSpYnhDe3eOHLTJ
IrZvUL2MF7WuWb8HRz/drwabOYUEhvYsN1ZuC2enoB/EAQVuwkBqnhj+/sV53KmB
MRVD5FYd6t1cwCRJ7nEqBq9thmPtN+3o2w8xB5ks4OaWIgaGYw+5/62QGKGJslIq
FOk5o5NesAIr6Fcc2Kny8aouLhGlWy9yDmvL5kSUZYmyAphWFNXiuJTvYeUUsEi0
2s9Y0HHRXaKRykO6kIWGsGRekZ+qh7SMzWlpKPLs4Oc/xPOYRc5WZSiLy82WLZWx
lxhLxS5ItkaN8BFGB94BxYV2CUBHrULrrpZxZM/y3mrJzXRdEcy9BWbZcYfwTprJ
kAl4qY05rwsOo5tvoEY9nFOQQ3ImCDpAv2vVdRe3CN28yB6wydrwPjb9MG2J2R8I
fRkEiW4PGbLiJT14pUWrHTKzKN12MU8/mzb1ueruoeiSayR+nR/1RFG6iQzwWoEy
ABPIjROHonKHW9NsMSXIogkvBpdq+psTQkecyh+PMVSbQVYwmhfT/4CWuI6gQlGD
WtTWuoHXuZ8t8K3o3zzfamDKhOGYDUrNzOLkzwJhSUJPt/FgFR106xwZRqJ91BUL
/+4InCWk6aCbRvyWM80+G+i5w+jEfRcADNfr1iBFJJvOtlJ02MjBWpaJUQhoTyVi
sw89TaRynxogut0sXmwt77ApdMqd6kLHMTMRwiv88ApFtWCIoGQX1rpdmTHMxpGi
jJqaMW+1mmM6lJAGPCGe5AYh8nkNnmdWPERaE/nEi8ijdTGn2FOmTfjKK9Ryxjbm
YuPgrFZ15bzdWvny91Gr2PsnNoASTZenM90/sjW2ahr53BKxHqPHZaRUFBdY6wDk
Psmz4fOllZ2MWpFO50/IPK63LSmGnua90SVMdchrJ8fudDDGZ/434ZE10WYfjYOW
8ql5qspy7OVbxJLa1WNig4CxLPWbhpoh/o1wGx2aMtDSuXHMXvXI8TaoOr4sOa09
UkS+6P+orWHZoE1bQAaSUoXfx/o0jtpjpCwM+fy/gHT291zKLhU4gpgEHQx1GI59
WGNoOEO+wPfsjByRN+QrqEJxcv+rRuTs6J+ti/4G6ZCgp0WdJDSGnk7ISFG3W0Zz
NgIQ2xrk0C61+bvvTpGaTL5HQP29E6bEoAwbqtQdMnp4JhX0WVlCc3OQawMGEEqA
/YFGFlPl7dsoCycbZB/NNWVTBV/GADqO/q4c9uxuIgeW5VFa+LArRQ7HnJ7bF5n/
SvJGT6LyygLxZGSWmscnJAdPR/mbQN3ke15JzSf+zQbNcEtY5c6r9utpPzu489Gl
CHf5MBBnrpK4kJSxdhTUeMHmxMG397s/94o+ZVUSXK60nNkHdGiPSpPMCiOxEhO3
XCZCne6dZVrphy6jkfYYPWWX7phV2Q1dTDuxXUlk30Lxs1TJCc9nThNHliZaz8nl
Xm31RfzGqXfuermXdMKf7uEvtsGYP5peftj2o1CxRnRT+T03Grufm0m26CuxqymR
jMvlR8IOhucto7Tsb076xsIo3r76JspAkv1Rpj5tLFDFytaOs+9tHGr3kkZoexGj
dtjSniejnzsLpXNrDE1PFAw9N1/mxN6+LXJuyAbXP7KFUgvfG/tqc0rHbXRUELkV
ex5r4mk7JDdMS8ZbjAPhJqd+BYR6n1oF6e5EVTKrWBsdwqFOO16gXDK85LmGQz7c
zAjmCn7l0oieiSubYRZL9WbX5U8gQ5SnvSYLUdOXNPoIkkAeUAtBUfzNeJZg2OZ4
T4rmaj01+GsSW0KpuHimrKiJPgXit+BGCpr3Z9BszpGxeRFIRmuAhDAtOJd3Y+H4
HCQq7Mw1YtCH1FbKWdOQC7PsuHDyzJXt17qhpGz0Dl+M4p+J4mslMgTzwjXukwBm
7zIOgN39/StzIQXgPUIkQSIbwRorUrjnZdMwszbP27ooSS3YkVBqxSoP8sfaxmkh
giTvFPiQWh7uyEyTRPPKoeTdSBv0RZe+bMlUESe+hHcs/R5oJHvEHod/GO7bDVbs
htMXI66feNvt05Y0fiYgUW3SQmlsiwC+CqT6tHmrKReG76uNR6AYX4LqzdkBFBT3
8qDMKF9Ufhmv1MM40yUAFoJTWDIbpcotGyHBXTD/zmcrE4BAGgLfUY0ni4wWLuy+
WTEV+2dxjKpiOcE7twUTWz+clUMtnM4m8U1+tX2Z1D/4bU9ik19hsiymUyEX7cYp
62ZpCGwzDv9o5D3W23m0nm/fAS1SD+ZQuO9o8vm5wzo2dLOoKYZ1QxWDkLOmAnHD
Fa9Gc7cFvqzNR9hgNRe7fjIF1z5QTR+NJ1mJOILstTBeZv/Mz6VAeg3XZ2uIBr8A
Hq3r/0AxgPg+On7dJehswLJGo884zHR6jL6qyXKUKyAd2yDqETm8xNpmkznYkE/W
G6OAUxCuashxFRMLE6bFesrbwbp/7zHyjv7rrqdSJgAEB+jjvIMTIAeVXWd5HbTH
sjuv2Uop7IuOybLRcWIh+0QCgMXZdjcXL9Sq2d7dROblMqgCD4G/UheB4k1f5Jee
pFqEu0Nrzytbm2MtAwPhRk3zptClpVOXtWPnJAdEI3Lcc1VTtLJF3P54ZaBuUsFg
Wm0KA8F/mXjWYW9NunW8axI7NFvHX8PMD+aLNI4QP1gGSdx1ej13lsYJExLrhTd/
EHyGRDMf1GubPKBwdup7kesZOwIJfsLnk+zx0pLmGEPEOjdqAYuU1NYgcVTKGGOe
VuZ9wSxQHFjnVWpnXGmb5ykTVxOy9jlZ0jBMvheWTyKJJbxAEzusuU5aeJ0eOxJ6
+GTu+MCCnKPbtecE+JDpueeyIyYAxyP+aDKZVFyTTuOUxCSyBhZ0NjZ7hS1CfOhj
hrS230jeklwxpPUmZRn2kU+75zXbinQ+yJSZkneNyLmpuErki31CGJpNVDUCg25y
m0bZoBKelosoykNWc52m15D1vrWnwQLqSWMIrbh91DpchT9TsLVFgYXyvky6nAm8
udxiSA40CUVW5PCLx1Q5MGSSLty5y0PH7vOf6kfKPXzskZqz3LZSxw94K5qflODU
o8fAzdsG544ph6GwrstxIVEQfdM2CjpL4LKhW+0/4bCgSU/vilVH0dmu5OZ5BjrK
ZMxRJGcseAF3U3HJzE74ZudTN9gYkp7xjH0/y5MdK1D1bYnfvotkzSKpuaVOfqCZ
JMME0z2hvCvXR9B2Gza/Ldbw/IkBRCWojKNEGaEaCPYaEEp0Srs1ZIkPeLiIuxoR
FoqKGJXEy8dy0nOIA5z6jWIPdQr+Mj+IpGcXB/ww4AUB0GRZAEhSuQLPgDhAfQpN
r7JlgVKiZ73tpyhHyBkoeDM5NVgbztXBY1o1356Acnc12Bc4+GnMFb7HnqBW+1Yh
FSjAakP4gR75YDdeBtQS1DVU/1I9f1/ZOqP9BSMdYmCj/bSim0vWSSbDju65YkD4
1oCa5EQWB9/TGhNSuZmfTymXt/7Q2WfbUTOVjubIQzmR5Cuny7d6Ia0z30Fr+jqZ
9orOOV2hPYtrS0NvXoktA/bAnG6ilfaPAKFbCbf6XfLAS0fi6f1Vu1vxksmGRIsy
fna1LeHGF+FYLWtGqHCXGrIWRzrJfCR3zYVbVUFyfS3pZvZ2DnHj1x92Rm9pUDim
KtCN4hilzulS4Rft2MaqhjVDVmRoxHmxgmD/cLYbfCDiWnXl0NgUJnKYkCaM/I3k
p4xyH/rJp72Ohx/unUwnrMaFSZoWcZAU2FGrhaSK3uhQwIqm2kFr3KP7dIQ1+aAZ
VWOKEp2+KYjfIo+jFBNnusmqwCKWi9ZxuWZZD5L+cS3hiN2O6SNI4hWk5uLxlQRT
AtChZ8xRnp92CbzraNVDtLdfk6GdDwb6hnqOCPYuVzqePZfRF0ADuMeC67wF1xN3
/ZdTzIt7cYhVf0gmHwxi15RxA6u5E3gOxydYQVCWIhAkSi/GehSzc0qmdf6+zJpF
1QbNeWqfmKWNsksgB1dCrA8b/PXq9kXXu+wDg7o3Lce8OUnfvwI+cgq9Gq7OT5qO
3xWRDbt3JRrlqA8cN1IuMU51YkDln7AHabe+Fd4BILXPpjCISM74JbeAXUVz1d7k
xdOBPmZaVTmMsWcjVwdLcKaCLOnNhCRlEPdXMlUoAGeD0vTvWRLzAowbU+2/6qv8
WYKcnbmxixyaFBup4u2C7NZ6skAOt607gDev7Jt9RXW1VnHuMtgwsN3J9himA8Uy
pnL9pFAfCF45iYqC2RltOW1o8G38bST2GZen/fZjWUxrmVul4SLA4HxquJ2CyIHg
swTzlcM565zlPYOXfg5iwE8WTrOr6to88wY56oRdaJq4+oVb2IQ269aTbf5LIZcU
EafVLrtj5S3vFGXKMcrimGhVvzW0h/nwq/POQZm0F51qAp14ZXXT0nIv5B6S83R0
BlVeaHIPCQMwfvB6T5srp0IY/BUYOgvotAgV++zJOORsXhoiScyO6MrICCpV46No
svZuM/tyA/oWOqvWzGp9kT280F45mHSjbxnMuCruSpD9YY00XziZSh6cmk0of8W4
AeonLxy9dCTf3AQl7KwqfduBvac3ZuxAU+CxasKlsSi8eNR1vh5YYOYhGycdIg+Z
yrVsSyLIDrZ7ELqSBoPXroHylFoCjzCDRyAYtbX+FFVy2pImLWCYartq50f8tf01
upeAgfVfDJebNDuKwOfmufKaggdUz9Y0RgbQhVKYBO9Dn6QiyZ/8V2U3XF4LBj5A
SnqebF+TWWJC7mai1C31PCzyaSbPeo/STXkhbzdbRcD+UTQKaAgXx/v48TCFkIRZ
HYyKvLKbV44VTfrIIErVPLIA6zGKfsvLDD+tQXfdm++pbqVjkfKnh6uwjmT1qmBY
ORirLSFzH4HPG6vAt8iS4AOMLNEyjlnG4ZjnhfGbKMS8200VUnKgW7VH4leQka7X
mSR2ISEzdzE00IWSLDLyyTvHgO9cgOs7irwdHpY72jkF5e81JxdOolvIWS6VGpPd
asxTxfPo9g5WIOJJeRMlTl6DUfeZwZ6fCwgDreJqf7jls0QWmE4Hzfi42TCcQB+g
XZh23zEB0TJx0a9WxqhgH4z2hAcnumksh/GZu9XeOcdL3texMaKGg5+2w6W1bMcF
LU1NAgya6DD6frXMbLJeM7itEigLEIzAE+FOlNnIrTukOv4QffCJ72Xi037ti+J6
PkCZbuBVXM29LTTRx0a5CWcGHZ2KfAGVEkrS81yrTzCVAnC7CfDaCgwnghgMSTYp
t4+ar9WN+CkgoTUeMRo5qOO7/qhJz6ZsUcv35I8Vyk/f2qg2dG6RjXO5DHWmLe1W
qHt7/a1tmXMd/U3g+E45QVjA7ExC1pKKyVgiFMVaBKSi+Se9ZzuyeMjdWVY5wqh7
VrAzMVUSoJn72Re38QquN7GIwxEI8sN8t8KeN2js0iMKkykzsIWjkgf3vN5y2/1G
5rTV0OdJ0OAVVawB7JqpHLFIgDdecC0rlkseiuTuuc7XVYi+0SNmmJXfKa53UerO
+8D075tgPnz4/mPYwrvPHYPsGwKDv22kIOignquMYHrOIX4JzqoS2TSMlDDnVoCo
z0qsmH8K4YpAcxoBgET5M858g6222hls230tWqZAkRuilEiUCo/urVXPt7dRfF8C
N0NpXU7RMUAZkdeFpZzUq5jBrUuvdgFyqCE/PefDB9rA89BVbsUSjEJ0tOBJ8/dP
eXEJmZ26HOcRaAdxb22gUuG0xmzwVyztS6ZThkKAGm7U5FBtK5XQucPULVlEbhH/
SSshnwAEbrmfUUjgcpxWZTo0v4OarKA86ftm40QwVj6rBrb0mGdXhn3bGjOm3s2f
SbiWFk/WhdTG2qO9UN0kJe2JJSOSf9w5lj+bXI09zEUQoDAdNcLWRdVXfrSxTSKe
vjrqszBDp1YjgCT3xUz5obIFZFYyzWhTT+3WO7Tm32ub28cUGRi726DRv+WYOyOl
CfwfdskkCg602cMBTCGlBLS7qREsPLnlwDLVkqTm2kOPfevIwRbOvY6NHjilbGDs
amQ0OVJe74fbag3mFFZpQUSv1mzF0PaCkXO142gmrLZ3zN6TiBi6s7AFpJTv1D/S
umR4kltmeMV+3zeN+daW3nKdiZMkBb6VaKCEkU+NogtlWdpX2zH7dpZ7OUG9zFCk
c2LiFXyelD9hr22hPk4jUc52c7o1/wku5Fi44vKYXjft42fgNm2Q+UddRHjRQOIC
U00LLp/qW5zZjAsJ31x//NxslwiqIFlldv5z3WRiZ+54g/CzK4GWlQdN9VUoO4MO
hinQVjiZ2lBtaf33RyqUhgI9ag8o7+dH86JGpsPoTkfSHgrUnVaeXPFX9aDOMckl
4PrliVawIC3YL8STtp+vo9IcbL5ff2ijg8hYUkdV2dtNDOw3eMQIUQa3286KUkMp
YJ6h+q9hGKaCQZqvBw8aYvNfwSfT7LaQyplc4ER6f1EHp4zgQqLPwkjo0nHIsijP
SIB4nNMnE7kM/d7iiv7xSknZKaOL8WRYOvKyu82yy3gMHZkkzF2PJDV66saEccKW
VvWOvKi6B7iXXG6vW9dKLJkxiXqGDYMA75UrprbtQ7nKOAVmJjTf3sFHSDry2xOE
JpMeyRlowxygnejdl42Uat54D8uM1fKfKSxGSbR/Q8J7ViRdtAVx8xWHPOATMrEK
Li5VO3JK2dMAkyWqQCKUSTsHdpJ6ZudZTgRupIJfxMY8gVGLZtysMVijjc15gv54
nnaedspmNFaOlKa9H0ldSIDg20+zvVD0f66gqbiZ7DiXteN8JfQHsVgnDA9hMbp0
V4n0JaCLOlpf6Br6kTvas4n3SSQ2JyIiKMWnhDrcrDhaDL5aPHqXlDOGXDHEbJHx
vrkdHcefhBJklNGh+Ra5dnllKpzBEtAEih7xno/MjnArjvKBappduBpeC42eJw4D
aFwZPt/ZN1Axz4NYWUdIZQz+hC+drTPWsm6ZWzAIvmOBm4or1PcaTqbdFEnOI6Au
IjUpB+NadIFs3JrG9tg65ePjixBslDllQMEeA0a9YJIryuDAHRGeQ2yJ6LLo5AmH
yyiqmKXixKZ19h41BNfCQy4nmHDssZhBM9g20uIwcV4UbSDPt1tJalpYHtAuo1Yy
lK/I4vSlZ84iwj31Rh82WAmAH7JzRzkeclMh0ZOutlSwAg8MzRrZwcToSfYgN+Gf
TBFDMNh7Ejllo6HRdEtbZD70hmj0Nh/vPmS8fnWdWVfsQFX+ucn7RD5hvtOw1J4B
T3XqTDgcjrgTr3mYrWuLs2W+yIhvFmuZsvCqyG6gwokgMIA+2ydTBGAEtOeIA5RW
JQrP70bwDZMOvNafTHiFW219mNcudvchSk+8gRD4QcmZyeLQnVJzQcEE6dNwiBmH
DTLanIGL7s9GWplW3iPxLh1+cCb7oXzIDC/ko61RiE2PnQivVEE3dMwu/Xr6aNN3
526CseN5nqb4pkcUbhM778i1HxMHF7nfN4A3UWyEUzJdgNS+iV2nUMkAW5bRArpK
Tc6XKMpBmOwpUWAaLJXPqEPU4Yq4KJEkdu0uZBiG4tIHJWbJ2CTpxF143qLwdZPS
EtTbp9E/GpsiG5kCcf/Z9etH4RgNqunMFDfEbm51XswmZECN4JWEeDXrKyakUSmq
d+uH6ZDijg2nsXSOsOvVRBgTkdmLdpuCBsrhbTiZoKZ4I0sGknNvcbH291LX1efI
bXc6tSpJ3d6WkVIC/k1884WeNWyp3VE5doSpixaCMAhuvEUSPTw/yHI4JzeBdoJ4
pA/n3IOdBi9mHVI0Kfc1kl5HyMHOqNgV/q1k4G+jAwqJXPNwqJ26X2pjr6T5qaa5
coLe6LqASZspkZKI0i72YwI4X6qw4Jk13LT3wNXoD6BqXuVtCb0NTWXtFCxtdHVN
yLJrNllPP6UeQEB6a4CKlWo+NyQ7ySlCB2IQ29Gb74YMYJu/zCesHdDdP60mQe0P
C4EReACKzFl/ReX4V5I6T+wg6UvCAzyWEcvTDH1Y7btWJjVAtf9nw8IAB8fl9zVL
BZePA3JzAYYbWey1umnML/h4qrSJcnBrncFv8peppwYNtW9liYLpXoUS/0r0byjQ
VwfrV/nJFwyUIVb56RFq5QKCTup8+2/kgGE70HVQMaY/Ieel7vkPkWDSASMIjJm+
h1JA9SqARoMviPxbdMLqW5g4MJNIY4M5HT1UHdKC8PoTRMRHxJfkVTNCgNrQl5bf
zDvvd4ieCg/cWSaX6g4asgPfeq1m5hRX3rPUQlAOPZgZWYRoHPH8k3AcIydTl0Gt
ISC7Y8POvYnsVl8cqSSuxDmvukSu1BnoZ+hlURjcvnrNhVe2UtttfPjl98u/3LrM
PbBag9qOt610OobLncYo9Oqwwvm/YxBBS7bXkpbRzGVKa3HyG+mqg0J+IXIe80W2
sicAL1ZdBsnbMUmh4o5/fOSXSkH99XfCiD+u7TgJoJ3uUTuiKwrMtWJfhrnqcfwn
E4Jyd59zvArPAyDZyAVF/wP70h1FSFHHkb7CjNkFyOnAUkIFZof/U22c7qW7NIY8
gGgdtyeQuE390MA0z0w8hy0n+FTM1CNY4YunK41VPDioILcmUqAaPWghsoIq5ZSc
MCtl9bEvfI7B9v5TmRdtQs1WVd7axqdZfM2whN80ljPHi3IM6ltTrtUCtUnsbY+/
3RnjB64tNMxcj/5DNEqqzSmqWey6D8esUL3ix7Lj2eOk/kVbZ/rd64W7uovZ964f
o5OW855ezKf4/ZoX4iWfp2S/aeb2CMefZpux8uq8hmJC943B0/RbSRV7OlmHo4hu
+A2wfUR/L5RfEoC0yfI5w3qvT+0wQA/jKdRkpM1hiWEL+pWrCdGLr9c0zgq9CszL
Dax/6TQXFtyZwzbksXRdYJtWg4RNaYJvYo/QL7Xhqsam9hAQc4X2d8a57FBcUYPZ
UUoKzFGieKYvHsKmUsE6BzW2UzAn+9btU9SS4GqtKGI3dzJ5d+1eIPSBPH2+D14Q
VjP3EKjovBjsB6V5KXIOV/M/Lgf+t5bC1SSSojTjcUPtsWJ3WhxbBQzdsYQjfjuN
2u+3WpxG2dzvr3iwPE1BZn9DGKIPs0XJhqffxmueqNy0IBtAJhzOeXG7USMXNOFy
AMqN79PpOML61bBXTzcA019U2Uly5dTmg6JN2OCxaUNPw5bpAHc+aZBG71VUujP4
dOu7BKRt3rP2LWHmp0pdw6Mv1xgdOyv9uLkasSrfqtG1gtIhsfWKOhW6DMgF/QiD
EO3cawidkSSJwtGeW2DBymEHFpXAmAW+eBH9OoLhwgFSv06FrqjHt7X5UPbWr5x7
JUnu92iCfZ1Npd7R/c1vpWM+VDqStfnSO2OtrnADr6NPfRF1oy4KEAi7jYpitglz
pyuZYcAvjGx2k29/33Uui051vvQxRlGD2KPL3ctOGZfhzCRgJliVz+o4C8bjC0Ke
xMC+6n9GkwI+dxauHo7+sN32IRsk0BECKUJxb7wiNyBbPWDJZWJxc0bOMEtxB8B6
lJGZsx+yhca9LUvhsQgboKaagM+E0v9ry0q7uf6VQVWkgzUdYtLTjLUG6Fs1KNVs
w3eGoNbpp1f/0lN/o4nVQO4pZB+PUcHQnDHDOXJCGDRaRMiQ+YAFs0DvLj/O/2/T
HHcbxRuXONAIBjoPmL/4p9dgbc6udOCk43d+w+AAmZsOLlkCI8GHGeP6vcJp/nXU
VRrMtQ/+Kp16WigIXedfTRjeb5UkYztwfLMR+ddVsWnj4QNsdJfr00O6pvxuomtZ
E1yaD5NOl0e4cKKvUy+uTHSV0Z52dR45yprQLDA521S87e7CskxgkLMKvac2yTap
BE4CKAK5yNONJAE3LaI9J5iq4PPmusMbJ56aVKJ3ajRbFdSAHejFJ2FJL3DNRU3H
2zTd5blsZsIdzTLUeoFIR2DvI+xhx4vhYpYNbgjCIhUp7v35aMzLqe3OSDBGWhMP
sMGgJaXBJE2KeGR1FmbVGH95vEmb11m168pw8gF9s8iFllidtPOctEXzttet3mAX
gPcKhq+Oj7Fr9N/vMGaLRf6AdLqS2KFOemufz70aEkOWxJpaPIqrmUAaCSbT82vv
el6HIVw4Vc3q3Q9NMzy0AH4FEAemRXqE8BnNFF1X+wRxKrrE138C3RCiV1T+LSCL
67Ds33iz3f93+UVPU7AuMOC6zJxCq3DMVCB9wPV2Bnst+YxqW410BZQSIjPG6q/N
no4bFaPCodPfrT3eFpktiKFI3mAnW95Rghea/NOO62Kf0d210uBi6b3C9ix4tC3J
aeFiH8W/4EPQ7N7UMJF2Q+gGZpVZDFppqyZdD+1l9zlXXOx74gZ7Xj05n9wUYMtD
nxD2vUlySVICwhxat1avFdIV/FZlPB+1UNWTQkT+/0NnbQctSCqY1wnWLvt0biYf
ifBDvuLtXTxGn185Gj0MKClCa84h+mCMC52pG/9zTouTniB2l1urng+jRuKiAgbV
avM3DE1+mjyPwfLDPTe/rwIXfvQ+0Nv60byvr6fUZV619uttykgJ2I/oxkE1QUEW
6zBZZ5BrbsKrXb2YJ9uCI+l1B8t8Ysm0m2GoGCvJZFCNqa/mR8srJAr/6iv+5v9H
eQoZla+7feyLrWbG5wjOG0hKSh+9Azv2/c5W0Bro/oXiAIcFVY50eKBRiPuJuUtu
TipbspXlO2OWAZ9VIcAh04L32o2ozR2nDTCgwxfMdjJxNbtKeYAxCpNkMSyJTZAv
Mlgo2bcfs6OCLQODr6TB1gnpGAL0rPJuwcqliiOHkfp+slDd0JE86WLT7BYYggto
y6PYYRIYoqkovBc3WVvXr/KiC73f4nbESGfU4ST2MuyTAFzjrC19c+ErvBWZRo1T
eEEuE6ljDHMRy2u9AErzf/08wGPKrO/Fveyhj70/bE2Ak8xz7GJRU6BoPUCH35Lx
qBe49J3t9DvHXlBwoML/y0VC+RMBjOZQ2mdrK/h5k3jUQitcH9hDVuEcbNxRsbHz
En6Mf6MGQoNUkTRkUlzwTc7lnYSjLRCeyLJoIG2TP+5PxSHbJQQgQnmSiiWEraE0
+Fn1h/Zj4hk1j//15Kn9KQFa0kGhQA9QarXBvoSHdzxnX0zA0SeNgm7WVp8skCxB
Vp6o/OR+9xlUTEKZ37bKPTgWlhAhcZMz7wJaJGddKTuHqS7v/binvtLgQyUtY7SR
Uod7Q5/bsKUbRL6R83l8IPUk6EmojbqSnKSnn1eaX4VGRYPAkTVk986Jf+6+AQME
4dyyLwWYjGHGIwKXBvxCdXVrquQZxBabTC93WL6QgotJp+daNNR7JQugkkCHoruq
cakEbJdqtxh9RF0DgfteYmzvESJjyyGX98YjIohwcmAybaSEfVyrq/BbX2xt6P6Z
0nqLoyttDehl6ImONlwNA9VBjdUiuO936HBcZgjyAXNblHaJ+ufcwExpRRa+G7VD
bRKPvquduyAH/WoqJ5V7l0Io16iq/w99HRvef+Ds8AjbSEHUSkXX9cWQTkXZMY9x
L/jx6gc0yGDS7BLDYvbm9ngDvYAzn++b61q1IzMZqySZP3Y3FV2TDuYqjfoaIVch
7eJSz6mcF3AdhPkfjOt9t03Yyu3bR7qwtWmxYXPYVhL5RFPmLNyIqaR+K2WlgcHD
Z+Cz3WCbUV74c+FWkoEIJAvJbD27QoBCqjTxLAppY7CW6nJU97U8Zh4XeDnR/PVA
sg6G6nWugxOu/dP1n3A5ek0LAfdYOWBqEomw6WVljgnSq63G3NJiqEp8FUI81LbN
RyUGROW3ztejnuWJAK2mISXujXS2VB28w70FVGBbZDoxwhgqlEPUoFXc8p6NBnD+
3rW7sZDLIv1YiMdgO4uePzEcI6VgBfRJVSFtcssyfY81UcUS3q4AdSXlbyurm4xg
iA/Yo0HeBvUakXqw79eYmj4LZFYK925/n/05sMjtneAv2hmHw08OdQVQDxwmB/DV
3MLDJ3vbF2qxBEh9n5l312AFdPW9uJsco8CVTTBNvFhFpwrkLSIQRpqF3JJnQ2ts
oJ/PMjVRMY6A8h547N3b+RxMXIkkD3dRw8+IMAkC8HKqwJE29sRele6KKtUn3rZs
RNGZAYhLcdjlZjALNV5MDVHi5ZHmxGSt9QpQduLoMFUvcSEcq2UypYKbu/otlPPX
rcrl9bOUS8rOQ2OUUdXaoNvnf8sh2je/uG2tf1JFOcOU/vth5gdwLSRyePCYKmBE
o1Dg3PhvO1WbPNj46NPlqr0IUfjIMW5CaOkrqRJ/BLVpqq6q6zG2Ch5UD3xfnX8x
8k1FkrKJvGmRvfpiaQ7PCpMQaNrdoriPTrKUw9J0+yBzEcL2M8VIFr1DMU1sZVxL
aRwuYLhYOoqJ3yipZFOLLzKC3BZTKa1xAGJL4hVXOxEQpF8N1qU/LCOtv0zK+G4e
jXS33p698gH1Y6YlOI3G+FCOnETo4Vs2Z0AFa/EGfOsx6DvENb1W5TYrdycwRcCU
jAf+LAKOFPA2JwUIYcnZbeHYpVPsZ+RByiZDuTtOCj44Ik0ckSjqD45bPw8xipAq
cZyj/inaBOgwarBI9hXdDRCIKHU9ABfO9csq+IXv6bstnEJfrolHN+EBuBLvH02n
nxy9MNRJ89JdOca8VBgRWFyhGYBHQUZNt8/bi40u5e5u1WQuaSFZd272YZQJ4prf
VijIa4gpdazrMJbtWnZEZPAxW2J14E8Yfuji/LMSCx8Vd47OwCUcmwdFNfxP6cx+
piUE+CdmWvWB9iTCSU6ijH+tZnhrLMof4fdkki5b/ehvjXR2+yXGtt7see/ueEZp
DSsUA9TEhQnVfT8Ddk484edwSdR6HG78at1yTPUM5B4G2jhfRZjMzZjCPh3/p6wJ
ceWOF/KjaCVfuRrPdKOc1g55dV4kKXxnsUl0/6wqQ3F7PNZOJhcgl5PKCWCopzu1
j0uiWWDoubLRybDJ/eTuvW/x04aWhjiKs0H2Q6LPlzFZIgGu9sjKJPOHKfRKhrnK
ICgI5ay9MbHuMD1HI7ybyAxOimC1F/fdejTiqMxf0YFkuIb5sSCZWhyh0Jj08uvR
70Z52WUwzM/4ROq55OP9IMeSf/TITXofJIVGMaUpNgocgiWhuyv4FoVAEMAEpIJg
LcwDwMyMiZu1hJu/p9KCbRkTVuW1nSoQygcJDosmVJc8TScOwRi1P8VhkeIaSdS+
tOVF4P9d9a1kNdaRokin7JpNfxuiwm1xL91HUBFuUZvDqEYmvaa9pF6M3P94pep5
/IL6l08Z0601VK9kD4tr8NnLJHdYykYHCHJt8YSC10iMY/UzmbnLCNI9OQuJ3Y4J
H3EL7JU9F+uPdIEOsmjIFXF7LBFE/kja4Rv7u4UaQWplIV7swXCxlG8nBHDBT537
wkOpRox+6coSZqms2wYaGF6BArOeuiXOyRFRcu6ap3BmS6JYc2YXeqxImegIJ7G9
G1HluFzt2PuZHby07Ijngrncu8ArisMWakSwUZrv3yOrXcNr6s8ok24HwdO7hmYP
Q4/imP/e7jnwH98fSoJdFoZAgX8AJXtykW3e018F6wnN6LdT4u51SQohpreYtx4s
4hAOIzvDQBQlXRrb1ZSFEpLet0e00/lWJIOU9IZFND8t4y07RM8+YKMYVSdfk+3q
2kaP2dhADfT7i5M7ed2dcLnRjOEaQbO3wp9TJtn3thKqmopGaL6ytH6qHmJq+TTz
HdY3Ma/14KNd4T4Ycb8plbBwK7nErC4Mp4H46PGEQohbQm+y5WbOoTOfMfyFC3tv
/Z4RfIaCYNEN9wKh5Tw/FZIDoBZqPJijzcS2vGyx7ppHi3TXQ8XkN4Z7ZZ79I2I4
bhHqb7wXop+Np7FUdHo8O2TCM0sPECdtNaJqGNlE9UNx+uGIeO18kKJNTI+sfG+2
29rufXRUcHlZfH+xw3TxhviNEhJhzw2lFoP6ssNPEZYr/QATNtcF2yvki5OWK68/
IrQm/XHH9ltven33nai4k9g16Lqjvs7p5cNA6EWKur2S+GwF0GBMu3K7u2tFYr6k
gXqE+MWw0TXxQQ4rniOYBe8FzTRrCzpH6n5qz/WxOUefYOJhbQuGJSF9xHa/3hBR
0R08r8wfBL9kRKCuYDsWqumKZjT4R0dBa9W8faP/uX9rMQJ9rfgTR9JT9qOynC37
86jMQ4u2mlAeTpkiIL+Wm+86IK2Jowjfktn+tkBBfp4pG/yhap5/trEPgxlnMquU
NJDZRJDAQ091EPH/uaTKJZ49hFNxICyfWVWRWXVa64XdGeEf2a0LjkYVoq8G1v2p
U+TqpHCeBMpMdfOPlGpVdakXULO53DqNvzZ1BpSTUsJ1QzASbHfofa+ls92IDvrw
+Wo0fizy4ZRt7P5JPfDYvXY+RgF8NhmB63+qjmoCin33z6gUI43cLwJUxzxBJpLt
d6q3AbsdWLLFNbFEcjOCsmoN04I2yenF0JXcZPPDT2A66symLleKktdNszTd6yiW
dXHe1lpLGzLQYLKIoCYtg7AgT13MI1B5e2qcIV8XRudSlU/cpCcClOf4zaWDoXiW
g01dcaGRZnrQkLTJ/dK4iAAKCU+tYDOJ0mmcdUQpLiwZFLE7ETAAep3g97G7rW42
Tfwpag3FeyajGs/7WM7aHM8EcJUc5UyPhrN23Q6V1S/kTgVduipNjSubAuNDU4IK
w1jVCl/BmBfwd4XX4XRNsHLFahPsLvXgBDMo1HJa+Wll7F6k6J8JZdPpyNjOokAS
vFPsdLfkQ4TdFSkS9/wxWIam7aF6ejihynvu/Xbtf9tQqOsChKGNckRulWVW7vG+
DlwNqCSCtcJp2SphhcZHXSO8WNepoOa0PUAnUcQ3bJQ7GKilymoKIHeradTwjvOH
HYDWdThc4ue2rBlyWp+MGzNxexlIbvgAnAu7LjttTnviirxIxLPCARet3oXmX5Q3
i3/b3gv4VOQ4eX6LCpxo6L3gdtgQXnN4w0QUeg0mKIvTZFtCYz1tcTV79TwRrbnF
ljmjukqzMoP4WyU+rknADH+pcUt5IdWE2BN+hfpfUm0SbfViRNN4J1UGKG4jiLrF
z+Qrw5fkjiyEmuAeVl07y0Wd9j3yNfirA5Ak9cIXa98vq/flcQHmwB6ICG2tmZVe
/7Vw0SNTolVaLxAZQdpTrGc8xkt/7ZJlk0a8pcMC/x1xI+d0N2+xtssCh4/Aehyn
sKGbIF7/Z9zPybEiaGCZmx+ypIsJXbSJReQ+g9kAJJhW88PXDV8e4q9uBPx4VOKf
6yRO+8E1s4xfu5JPpcD6STAU+Mbes318HwjbBz4ivPba1WkH3pjs65zvMfl4pgT+
CePag50XIw1bxYDLl0YiESzEaaZbeFGyiMK/DcsR06U/dLSdh3XMZH5zs9FuUVEU
ZiWKv0NYQgNVoJ8vf6MVAw2MYwr4+h6WMkrhY58RHm2uNJFKz4Ggj6Zjbp35A1FE
PC03hOMwcEuf7pwsztFRxKmuX27//f1o2NgxIaBsUt/awPipXWGf2vtOa50o97m7
7TGEup6nLaNEQnyVj5f7E4c1roDikVlXRmRPfzd3pzciG7OADZreUihiN/M4rwrZ
YGh+oQw83vGo34q//m4lTZMzeDqJNeEADuL7rD7KlnqnPvV4zNXW9wcTVyAEQ9M9
Du2QlYewyla0ompKEWpRPn+fNe/qH1WzvdQ2876YgFAQfh/wAW40QT9AIpJ0Bk1g
35xhfNZe3OD1ZOW2RLVTbudt0u+m7IbeyupFxF96Ki7rW7GsO4G8n0iE92R/hFLL
/f9ZeBMAloOylh9JcP0LTrsQuGGRXd+LPWqui8657Zdb7EDp2mvi8czLy23el4ch
vMxEGMgKhuBjfTvKVzTT9W55PB97r+ERez5Q5aHLLV7xELp02t4ShjMGWI4tPHcm
THHiOfdVxnyUwTVy4djHuuyubSRzsLS8zvA71zxmEF9U2PwdwpUI7SgLmzXpKZBG
3N7w9fpjcpALFU9thnlzzMn0sUxCl/cl+007xjfI/xYMQ2PYaW62sUtYkaMDRScg
r2tS2e/9aqs1KC8ATqWJ/UMJiBEYFD3sf3mJSPLw//f8O5lKd60zaCZA7uL5V6DM
Ldk13zE0Xi3e6FIi2BI2jKEXdIPk426McYAKakBI+fTjuOdd48wnT+5D6qTdXtp2
LnJRveoRb6tQhAKn7JKH9iNl27uqRqSRby9b2MD4y2pJKfUqG8ckgglVWyOVrgYI
pPOXeSyHX9mn4YKJOgzvf/CXCi6U/X5bZjLBexODzZbg+GvNk33n/SN2NqR+bB3j
ZBJIB5X6EUY7umNzTMzmEoSEW09NfFf2nQ8ol1bomi9mEkJDnkfyqhyumGU1ZMxc
Duuwii/Hee4V1yBbyNROvJQfO2z5p2ZSp4OysuBERvmL8CseXjtZJIJKP0OJUHMz
u88FODaE5ahPH7h3Xc1MM+iDlPrhnfJu5dGE/iKJ3Wy4NPfmYnecOJoF7UBC6XiR
NKY0yziGPAHWNvk1IDnrjUMzErNkP3eWJ3TARC5Oub5vJbrOrdue6lIvsW/OAI7s
8K/1ug8uKelX+8Xjk6CJzo9/yx4bLicGZtQN3gH0beNW4UyqhOtzrFRVRA/BBC5C
fRREwvgTWyA3uSdpAXIVq8wZOQ3TOhMmao6BeQD4jm5MaUwrMFhPC8Utxepfd3eH
sew6PPlt8oKY3o+prg7LKfL2RV9g1DYfsxu5b0Z4wN3C2M+A81Ro/YJaF+duW1qW
aRpXW+8wIM9ow3LrnPJir1oSh89h1eu/dxejTryQQu8KEVRD/uvM+XRmHRpv5Abm
+qbBTxCJDoFgFjkgOa4J4LeRX6nznw76KoKW8VQci+PnZVKe0CR0ll/Erz7ORVc5
bWGdc+TFQfUnveOwAe0+id20gK1592dkS2HNS2bS7dMeNDhSw1llmWvl1AXuNP0n
P55qja+yffGzZmqMaQTaa8SETe8OLDn0R6QPv4otDb9QJMbbGiGGdNxpP7/GojCf
tHsT8nJU1pS6OtZsdK1nTqgQRynBgR9Bmgub7i1O+LrmNTKNwXHGJEMGhkfBBYqD
Id2MSHdG1QJUqRAelhkE4ep/h9Kyo78kvH69M9k48Tf+kY/xMn6ZZ7EXDX3qBawm
HtnVgfefrGo5bE729y+L8k/DA8H0jBD+n66DKvsPxkpAo6sBG0gfvcKEgeUToYH5
NQTV2bH9YIjiBKFwNKzq8kPk74jPQBwybQKbSQ2cUYyesw3x/VIF7rDZJknTaAEB
IISgR2FO+Lhb9yzOrGBABI5hLYf2hHiQHocGriwiRcHy7yZwj/UPrrfJHLhHghos
5f7lfiW63CqY04VePlZNHAQxzO4wVlggryJbAhFMpz7HLE3YIMi4mzRhdmpABiOP
NAqu6+ydN4ZvKVugogJDhRcdtcOCUsBmwx8U6zyEzI82G2Y1ASFgzg41nmjZ7+RT
zuGiXQsbLzDqefYaBvOLxdTGw5riofsMA2Ju/RZ2leRbeWT+o+/DfuSUjLgfzmyt
2VcZL3v0Q+jk4DJ8XAJqYXjFUMpPpID4Qc2+jlfhpzj/KohvkOv6/5eISLf5qyKF
AZ2YT3sIJl5WnWiNgOlD7tw3jNuz5hqdkipPPTvcLEGZTAfPa2B7lDWXE1FXmtA4
nitncYM2e0mbQoGQXraRYqgKBfQjkRb+0QMStoqKeahjmRQLMGm1cCPI8NjRjiPo
1fCErQSqhBinBtF4a0GiPo3UhEDJh2KPdT7Rs5h0e6NzCTqPrwa+mpsPVpSbqvla
xyCKwS5geUsDLRnxsWeezWz+/Wi+PUXSDfyQIRPVJV/Q93gb1qLZoFzu9ZK6nvr8
TfdXiWnqVuuQbDhd4IZVKakruIn+otVNIdQLvBUiIufBDFDUh17XFdu+HCtBZPSy
j3a3x8wcDZQpMjG0BNhn+JHOw4meJf23WRkt17vX19ZB34MQfOI415aPvuSVNXEW
hN6bsPHEOrizRcm9Zj94zOiDDW41q5uMxW0qojT1aHsDMv4d0UprCRAScoXNkAj9
HsCeb5v9lBb/oxuT6qQw+qnw3tkxH5CQfn1bQP3acCadYTKv4ev9qqIkK0pVcDJy
L/rzT/mgWAd5iYxUmHJqfv1OMzZGu8EObyY32WB79DPbolzWp6IZ9xomQPV1btHz
ukMmeEOE9pJ9tqzbzmbOCTlNeisB9U9g8V2b3Zt/IlPChQ1Qzuak3+m4z39h4z//
zkiJReNSLzTxzrkr+nWEMRw0SDE/xbSOg8aMXISXUXFrrKYRI15ojyEr0K0f4Dq1
PMByuwQK20gKGz0uCbaCTRRnxhuvKXTzf3sUG9OCM4m2EjcfaXXynSZQkrD3iDKB
HUHlSUkvhg97tBcUBdiTDd04UyNHV8OlSPKwGb9Mfj0c23skI0K9W5OAbKcdh7JY
X4j0qBvpIqsaSeOuark/n53Axwg2bwpcU+7A82ZKSPzGfnWoMNXj+3kdXK05LqgH
7eK6aPFDgioc7thi5ZHMUDH/R2rh7CrD/ZiZPMroXcowSy0GAkuohnbUqiBajtDc
FGcpfJKHsZ+3YdFFAkTKjW87yNQhWi8xcImsrXAYcs81Fakhup+ADRuNy8/Q5AXd
8aKWcqkCZI73Td08nF7LePzFZeSfCN0yh65JxNxYpOg00vyLLwKxKId99Voh/dm5
9ihP7RBt82SpoFAPbeMhr8k88jaXapCx3ifvd+a2AzXuTVOE7LWKi9jzvYGlcN/q
yaXXmf5dbjznWeBpXtiO9yJ2ym98AkT00Jj3nM52QKXgdwCwCcsnFr1wZifRlSVB
rzBad6MeTBvl37YgFqY28abe10Rpy83W2xwGSs66JM5ielBw8CijdVWq619dPzZn
iv7jJv5rWmqERkeksJe59d7f9GY8sBW24xSkMJ8q7/q3ZWmPhwLBj8iOf33zl8sN
w60VJ8LF6iEy3FC8YwiPzYiZE0Gb/4p2chfjuTyX2x3rrXmXXZiJuZNAHGdOMaGX
x5IH0gWEWBfneASH9uGWJSn+t+20cYySMWdhyWbE98yLdOAveSLPWEAdbvRDp1c+
dgejfC2bYDJG0myfVskE+n+fCecwjFbS0mCoE0tTdlStdTITZ4G4kJ87ZlvHr28b
WjfQOAeVLAoge6V2wnotwkRM1ckELp6DLSFYyB9MljCWtlhnB1bfV7GlZc99xMjB
M19tecLmy3x0LcZMxdi2qzomMTaGI4PFijqmPdI+08uX5mMBsN+iHSQj7BNIl4Np
UmyMrmGF0lxVWYr/2689hg2Uj2elYF0/Nv5Wj07tbgkjQR59hsb+IvT8+y/Qk4kd
s59LiT+7ZxLweAk0r25VsMk9Y0fJVU5R1ZXyumcoW6zqgx/3kyFUw+V4qBaQlkzi
f/iozNPioQn5I9KsQESty4VMpF15h+y9mPHHGHLtap0qCxHKBJOvipVztP6pEzmi
EJ2nEEPbQRBlOalO6+jp6pHjtgYkbnEiuPBUn1JyvPxoIVqujaccdtT6qqYtFmiK
VU1GP5xy5mikvg486gqy6DjPRCnbWGzMk0c7Xr8cnFOZuKZuR8evUgD7OxSIepb6
TMSIM5dQZ6xIST7xcvKARVqQi1qIZNmqXys4nAI00wUBexb4C18+vIzI7Hb2ONst
Pxg0E4cInk6QIA9sv1BFLCEPtKcp4E4MtWWBA2+FKTpzYdmjwuAmr8Ayw1fJhhs/
+E4miL8/cpqJFXAAOhbATqa6PHtfzhOQL6HT0Cpig4FajH/TbqmLDgI11ImBMhEi
LIy+DIw6q/iXXlVHM1m6ZBw5qhO5Czmk+scYswOC3BjG8rCkgeC34cwmJhIXiQXA
QRn69K7eThZVCGBBG1TaH62w60rSqH1jIO4mTFEXNh4ceUSp5wgAkGiUVRtnLwNp
1eNTJUmCwc9eAuUdx3kM5Lk1aHTESgDzdLtbbgmAn2ilGhavSFEMCy+VKf5y8nQM
LyROEcodgbB9hX62Y4KyD3Xu7via+VE6rSLfBmaDysr8d7SU5Q5s9d8q/tZqS2fw
EHCYcu1vDh1pxEH6uFGjmhIEDvQ2cOKnOr2+xYLwaJCBxgIhfzoFOx3PxPN6j9pr
hDux3vj6H7M2acSAyJEfewyIG5R+PEAhYjbLnoOtAF/x35FyGG6hddp0cBQa7Ana
h1a+EJtRQ+AcgpOUIPA0iSvGa7m6FYHg8xoS4ebvtjb4VCWghFpX7eb6ZFqieooe
QsknTnZpopzApWdwZFnMYUqP5eLEmusX5Vlvx5WMKmrvil8djWuhCcSjr9qKkTBq
913qDjF3UUOZ/HWdlURWCzjw6/iITBaMPkfs2LqQgSeKJWIqY03gmm+gKYqSrGGT
CcJibb1bf4WtNnr7nihK2OL793NBpOrj0+20QXKErXsDBYurO7P7cVJqXK+BYlAM
1esC69WXPz9GwovqMEMeW+rWPk4f98JkcvJUjixusjI0XI4zxHuUZeUFaNndd+aR
qSW+o5AvmjO/nuLmD5ZpCkHAbKZxj8GcXvzGVvKf00rJ35gOc3RE07OGxIZk8esT
/TVsHG8AXLdRWiC/YWNDGd13dYKKGKs/W0IMLii5tqUNFoBdq/gpSnnd2PBgGM7e
xFdb7mhHewmyu/1tBm4HAHd+gO682fZ5YUh39K2sk3zGamwXZvvV7HitSRAs96ug
S1G6kWwbNtqTVKWDUR6Ww8IYuKQ+0c0ifdlNqfJ6qzOAA4+C3ZweecfMXD/G2Zyd
8gyEBUabg7GgbjBa+CaHt+SEh7GDjpdqFANpoZQWRDowGRhILJ2ej/GeS6d2/bn5
+o2z8ejapZpLzPzHIcMdqDE+TlEev1tQIrKf5pFecSVNYy5vxhdwBFEJ6g7yMk+C
syqRvCnmxuM080UC+MrTF/iKHsXFQ43a7+Q+Kno4TIIgwJFnNuZ8IzBtdHusGm+w
bJj+9WdMWyhFO5JLNFe6eZTozXamloUK9tSwrL7rKkAQJ76PrwU+xlS2us6S3BGW
iU8ybxcXxoahqhS9Q30xUc1y/fWkd1fS46Mrw4wdjr3j6H2KkfTodDaSk9L/CuY3
488N4PariZcsb8Gjouuhi3M4UEJwKgMT2DTc7SeHm/ShVVFOZ+ZW4mX6cL0UJH2Q
QqwHrH8wU8pfI1R8I+4di4G8C04aGkRjpv3cI/Q7NtPG22Ij1SSldfY93uFEw4UM
zi9TQ0iLZnqKNrU9X5wERlH9yRFz+Kd+xypU5MbpbNepW4vHu5Q9/4knZGfFxV5B
U0As/xId/KNy+dxsinQ34UlnCBj4L1OBfruoaGk5/0UTpS9bsj7XG37+eQkOJ2iA
j3J31liT4vy/RmWiLC7BItocqN8dRzbLYWrmlirhbqTdGBi20BGutKVi9KofsoHm
FJmN3KCKOuMSiEbx/YfnG07oDjxBxRNMJiMBs7fIhJbNGjPH9urzRB22gG05zfBH
n+p1O+rmrSh3aCHhLX6nboBVVMiMxvZ7+cJCO7dHOE+jVORpMj6VJnHFmacVAF7J
eIt5rkTIEjAQom1qO/AaV0GZLkjWmHqCB0+wRoMSxiJky48Rp2SaM9jlAcF43hK6
P4P8D4aAbbp5dhoN7miwG+jNJhdaWDmusxIKR6SOKJiKCkpgl1KFiCmvQQkOCtfV
aZBrNRPSk6815BAqa7s7UTFjsspWbkmBokAmHm+b/a2V97Ntu3dTGdIoA1r8MHAE
jpEjywDT9dRcpzXkfZq/rzzXrpJkJ1M+DzpbhyxkWFYDmpcTA21kE9ExAvVLrY4l
T4VJeDfsMudHxuWPiH1FPn5JlanQLKy2LIaSz4o+HEd+iatQ8HjzHOb+6huTRTad
V7SKYHDGuzXsSSyZfir0t5AbCINSyAck41c6JtjrrJGEkGK5zpeLOkZSkTvgc+JS
53EJ9rWbt3NVDtq0+BJRJJkP2xykr6MXpwQBSVfp77AJoAweYD2KPc5nbidy9hsN
dOknu0J4DJ+kLez/En2MIfOr45BP/+fZe7xWM4ctT485oxcZiY6PeFUN1aTfkXkq
62CbKe/ilYQoXME/WmSwQk+YszX90sN94pEEtKS9Fclz/1tyhnAdVf57nhStIOyI
CRFG6pdvhbvoqNWKIkB/glA67ogV7/bvUl4k/DCc59XRi3mT4DEUvRxDnDamLo/s
uTfJdnzgph8aNtILA9qh9nSTus8xjojSe5rgcTjbZfgjEJhK3UOijRvZUynAJhdd
w2D7mIFImpIy3S0lo6VoCU0CWKvIrrxKwShISeJWApYGrysqmw14s788S74qYt2I
mPWMIxfNPL00pi50MOFV0cxVGZ8oHaL7FH3zIs4pmy9KHiDTWabY/efXpHTl1S2h
eOpIiw0/If06Rwp1Rvy6F7HzbCE2VofgbUpQz514UiLqscusg8PEFMn6gGrangod
cb6Ns8GWyDYdYtr0azAVJMDq8Xb7spqx5xM4cg855V43rjnDNnP1MV9U+EqXwTb1
+9OOkGTnnvcPtbhlQeremna/xL+Te0Z8zTEwPIR7TwpRQa6ASjkj59HMF70lEuPM
7ElynSE0VJorcKgXO2SXqXOl7No+r98Nkrz9Z+M8VFL6u8v/MPW9khOGSTrkqTrP
y6AqIa7D8YEY6Xbq2BF995JgfOwABVD8HJUHar9z/bH3CnY/7XczLx/ZW9p+Fy8j
7DK+Mpx6p4RUz5hOF4Csj0I33323xsJL3KAt1vTo1NrtFNfnKEikvvv/etSFD8Ij
iHzzMlmzR4CM1RjckwkxiXRaZp63Nk5uLmwfe2j/Vvb11BPDy1voqInQ/3hNKZRC
jeWI2VnYp+qYZWjDr3E6cQjsNSZJhdJB0gT1ZbBpHUUcs7RexHunmRJ7r1F9GIlA
Wm1chYA5jAl+oQnnSYFzyndYZLiYqL665anjThtejUn6MLBvVoKbLiQNrm/+jqCS
jY/lGvj1qTImCdLwf5fYqxtDRo+8WZGQWI1L6pwzeMASmt/mU6JSYjJm7GjUWUMp
x2sWuVlMtaAGaSbjhMUHRqbmZbgXf7o+OXETel+J7GcabkdGe3YDrCrX2qpvC/7v
lGqqp44eKEKfCMvdpJT3m6x/SdEAyLTHq9OCFT/P3LIeGQo4SiFWH1DTMysv3y4u
BgQ9so3KMWk2Yp36BgBE7muD5uvzS39P77R6ZYHnFLwvKmpJAZKfnEYlsDNTVTyi
jUq/W84RSf7pKO6mo3ikj35usZTNHBkZZdYVX6T7xkH5AlFJSGdgdYk3FbeZ/+8V
J39dBOnROJObLO25kH+uwf7Ju+XPG7b7LVLd9TW1mTrM5+ljBBAMPirK7aQH8lGf
us4OPxDGbkMYCGhnzbqqUcYl5lNBbcEdsZtrWmHTf1077c1DKQYiY7xxgp0ADEzp
CKaIyzhI8LmUQeDKno5GUPxtbrdjDMoFdsoaQ5YlS02CvNs49GVBmfgsXADZwlKm
iQb4B8XLPHJktJ/86fgZhu8dgsqOIssj2Bcdmi9BTg5B6ogNXB1LPTbv/25oXg6B
53feNsrYTPmbPqIIDCt8W113RJGi76u21VcQzwhrAxZp+hV3cH1cC00PNiYtT1rg
7EbrQ/kUmBUXDVbAFs9IbCrogj/tgdjJhR8S5/jiuJJmcuaGlhdzmAVPcgHdbKC5
L2Z5NOTHa6nvfWn3czltiEwsZoZxE2jYzja6I1xdCmX0fFb24nEZoaVpFRiJakM0
smtPNzFUngP/tYrFhtmJxKJxClQK3/pl4xEupWIb/o0KB6Wv7yI4+HBqXjWPA+2X
sl5YiaC8UfMjMNG8I8R1UbPNH+PSnCHFaDwWP4HLGbI2kL6/vYZ46pAmmP5g4kr2
TWmEB8h9WRR3VWozc4WXNG/CoEBIM+UTjwF/VZa3wywVrl4OURXErCDi0WnseNrm
L3j7fg29t1haYY6vu6p210LUlgwrJ+NvLBU/YjPknDvPHCLAurdOFk2YDBpqlK7Q
wAYVPtBmY2+ChlDp59qd4F/3086rCgh+IHS90dDOo54SWnP/2Wdq6fqmj1uO8/rH
GD53RqfnLSc8V8LJDkqPRgnB7jvkTQwC70buYQYmkMPQpqsLhsT6SgtEvRF5KKqn
0578bhDGxb64dBp1vJQ8zS/+MPhRGrT+RVqhq7RtnuH4hbcNsp/xSuqF0M+aIxNh
PAccRbbuelQBb4gRnfnYwNQgHPFqD/jHljXz/eMIvq26vkpa1v3cHhDqlyq5hTix
49imcvXdDgcUAlKjTAlHsXnzc1ayHXf+pKTsqVYj7Dign3QOJTjtXXgxjMlldbG9
KxqLx9HLHEGv3hAOuL8i6QQl6fJm+j8P31cQoT6DdKVff0EkVS49Cw6C2WiYiaG2
WlBmD8ZzR1zwOhBw7LcbmpWxhhFJHOB/TKWMD/8H7PshApzl5ZY7oqHvB5wbeTHQ
Ot2/207ldc6gx+EfYdIaNDDwnniGN4C6UWuZl5AOnjsQl/rg8ozm9bY8Blc2KBv/
Rh7a1qWnTZZ0VqNpgMyZuxiCJkbeRnSTuuOwNuYPZprmrsjYR++DKg/C3q+hvEUO
lArzCNSFJjkxcsOVN6i5SmpPx9DeozAtoUXOfpQrf00GRUT2Fe98J8QxqPBV1uhZ
mm7g8YyhbFy4ZSz/FgFE+yDmftGj0vGiC2t8C49EeGI+p9Rp6uVDJBcs4nOdevA2
SvaFhE2WYgSx6EaRq0zZ0hCsJ5AY6foBSWnuIcgAsYQW6yXWt7XJiTV4GSood79C
ooDjrFGwSOq2+TBnBBTVM3DlKgw6+ey5JPMgDSGUzjOzg05qcxzVsJnzdnBua5vO
YzOa+TvolkoEQARMNEgxtdaSavYQqlJFy3lSrsWiKABYUKnl9KuUrViPFK/L/MgB
T2S8/c6IO0GTdIBU0LOZ4WEKDiw8KNL/nOlfLP15zeiQB/ixBxQcnVW+dnr8j8f7
wdOHZtFRxql1Z5lDU9Q3RSkcWrZtSjoAHilkmQRfFDEIYnPQAbTY5SD76r654Pac
I5MWBoK7uQWI9d9qkVSwPsdExlGD47AJoub1MD4gLuDtmNyCta+b2zJyjIMOiCqg
TIMHbS7FE5Pyl0y3Kq1JPrJwFZ3gRz/G+vFhH0SnVg1X8oxrqemcr913rStVth+6
jzTjiO6LpIvOSH55p6vmk0kd+YuBBkEckRUi6ey4AgnaJaLa8OtQARdz6I6WWXbn
65f01rIb/EuBb/52AXZeuTnaAq3UKUeQX2Mk6aCe5h1KCc7FG29ZtWmBY+dGHx1W
ehgZ1MMjA99qGvLA8eLyfef/hrb/NukOsMQ2/iC1s/19ToVBanDdLOi1iSsZeNnf
nB6jz36N3Pk54poeT+KFVj9UA2iP0qKqQBRffPWVCiVtFO96F3JJJbeYm7XNUby3
fAOouKks+SNKS0ebsVBHKkvyOy6vPVXRY91ZEGzjkaQiIKx6kNxi6+82IFGFzV80
7EEgXK10BclkFr7zohJ/Is9TKUKc5C2gtyzQbNwOz3fMTRZ1YlUM1DGxVzmXV4LI
ukhn6eCwA8daqEGLIPLxjmwJmPEWKCJ08ObTnSA2vcPNTt7N/hj2eqvEucKnpmVu
vVUuN8GykYkBA2SLi0yzKY90/wUiJVPaTeAHHt463vqdT/KOkMTlcil1VVkhThNC
U2CSrgs+CFwF50KaHYk35y23DxpF44RB8vf/ZxoT/yIo8IN9LStt6JJJCXh2q2lc
uM4s+2lHXzyGY4L9+fdYV8uwWviEHSOxOpeBeIzsFtOgm5ILB4HUThJSUsTVhHpf
MLlrbQn+DsWKeHKHhG+KV6FTWTER77USFsN07z5wK2frV+CUwcwyq3KUbdMXO5oA
SHJ3IhCbufos0y3oXuokUAeGt2SYuLuHAc2tn2w76eYxUSMAkaOOOmx8rL3EwXCY
0wjhIR5CuNwQQbX0qyE22x/h3PM+vlaPFa/ja/a6YSXKMzdoKNsUsxt7cQXNWfqC
AD6mknT4Bi337LFot/shYQ0zchkOHFFHqQlnuDunJv0zrdqXp2DASz2AQp7h/aDs
32KvWQR1JzhyoczFvnkF8RsP5gJTpq/zsY774HK7c5UIB+OuXXsQfNKsf0kuUjc5
mnmA4u17tWsGC2OuJH/J4bSo+x7BkSuFG6CuDbJx2PZHh/DAKgCCTr7Xq2MEXEJm
Vg56WboQB+FwlYloRUIt2HPtceUshpDMqdMGq4E4P4A+20TmFNsaqYK+RxiD7TCR
QgmhQ5CJFDb51ElzgC/2ePt9RuH/Q6RhYNnamaT6Xh4E6VzfTNW5cabEArfS7aVd
JFP/4Pu5Sa6efL0vVrHBKMTWPYCcuozYyrRAe3KI1r+qNDfTvUKmbKpB03CCwNF6
WcMqJZYVLu3quvYxN5qc2jCYZ8JK7h3lBE3v49R+/x1Fg427Qy3st/ShfCXFaDGU
V24xt8Hj3K3o9Ny1C4nnid5uvgak6wrXVrKBF9KfZiLdN/BdGvJ+UotAMu+Q1ujc
uBppDZA/uS29/UsMTRAK/kijSDyQt2frZF8Ct5IdbNQJqHz2ZXMN6xrflY2b/mjo
TwoN8ByYx1fYH3UiaxQ+DsA01vDsCLaWQJuRkLRQA4oqKrn29DKWHqOAPT4W5ueP
LJzHa0Alwi3ftZ75N+IP75ZWtJrNR/XvuxPyHC4sS6Z8OCrp6jjFhk5owiF8qCOi
Vxrb5Z7O4Sk3XrvzPMSs77984UatEzzy+MDUXRV9Cjtm8c6Qv7AVQKcUdOmZjkJz
+kkUwLKHcZDTgL9lni8DLVoml8dJRsd80WUj9FxYRM3nvA5dCHWEf5aTRkAufO0K
PN7i0QwSz9/IsVK3oQBkNqIPA2cZtn6rXiNDRVdzgTy/sqSWzmrGojNOGWsNBC44
DHAKSfEZFrPIzsNOHFj3nh7Y7qVDo94tb/WsTbdWERUXr76lUA2rf3Ck1gTyqd6U
2WM0fZ/vTiRQTEB6o7T7WWxipfgLc16ObeYX7Eo851ATjhV+X/ndT7cPn/2+c86a
SoEIJvFrO8XOmZQCWnFZp6fUeDN7qCFg0e7qYw+Da8+u67Smgyh4HaPx2Pw7cnmY
J5mN1IyhFeSaV8GkTC7WuEx7NOtSrg/xRvzDHfkIfNg8l4r+VFygg3vbO8ZIZxBg
a69khwNw7hDlihFIZzCWpXrPniTt3JC8XdlnXqE9Xd1g24T4tD8A+AiuQ05KKd8P
/rCcEwavTlDoRxO5mbr/8V5I+hxKfHzFT84rYFyqBxfAdXcpWUDdTGuwHNoKDliI
xkl4IYX5+vZ6tBTTJyeEpzjZC9qgXEJx2yqh8Kjzp8psf8m5bXcIDDQwkJzyMDYh
n5/L52DcXR/wIkc3AZtvUTWvW5l8Bld6LDSTBJPIY1TskkLM4GMmGhsTu8JddMtJ
9vwRJBt1F4nw03HMcbeKXKFVY/EYZ/Yf0n5W6spqg2jUzE9217Yz5swFP3kqWB5h
O5lmnR0uvkNBoiy3vdqTupZZMIrIVXpR5gbQPvK9DV8ErXhoyJmil/prvHuXFxod
RdubZ782T81f6fe/GhBDS8Hopa5y04BKRmxOI4NSKoqjxHZYzWNT1siCup6SRp6F
kZJPZqY1UKBHHv8St0jORX1XHTOiiLXPKtLI69BHHUemm9FUU1PG7WG7gDYlKgBC
FH78LwkiFpNoeOYR55HX2W7nAOKE1bB3+GAXADMOGkAApDX0AA4ynZq40zGbV68u
dP7XuOrxUos9wKsXPFKPggY+0qqoCj2oK1OUTIKCwROtueeHy+i0MAD5fvl+NIsc
cEIzkqshdKJ1MtVj63A4PPOHW5u0F9RxYZdaSZ8+RFbF0jXKe+H6Pc8Wq1KkvjWd
DGEcAlOReQqE2vQBe/EesHdIRXwmX9wTTRzNz1bFcCuY7+g2R8pGar5MaTOpS17j
h1A84NIZcNWPf+yHGph9sjWDu/RX3fGuzDfvOAbCNphOjQ2DVvclUbWGcUEm2Mc0
3ThEFpa76tivgwxJZ9S0LUTM+4F7VpCoCq0gvaFS2KERa4lmKri/svG7HoQwJr9e
ueCL6Jb/Bd8QhoOJOVoNSJSNqWZLLINV0LEErjBL9jWxdfy+5hYTom2JTi4kXCwy
U7ugj91PHTBuB1Maku955Lor9tehD4gXTfgGpXrA3dQcuLNlXkgNLV0xgvNdCRUM
zlflPfGqtkZgKs9z4cLReK/iMovpiy8ygT71m2CM3m5PrDaYF5lIHSTwc3U/MIia
PlAkV9NERc9auUiPGyO8wpCPEy5Tb2BHhjxPRWynilsSSPRPal9EY8IgLoYyOEAq
mUChTabsAZiA8ooQitY+IYloOGYuRW0FNh5L2ryDVh1hYwFJfEx2GDUa/vsvA5e6
sluDFI5+nU71h9QU3CMsS+hSA/jOfSDbl2grLt5jCGMuVmaxrke7aq58nMSY8RD8
Q16WYJbKpx8cdVbFWqqYzWLenGSKTWpb5l+6XxgTFMXPbQ8DN/ubQAXTonMDpZ0S
vZMgiYAqamyOlwq7ynJVvlMEHyrJ98kyOd1hy4jJe7G/xHa3UVJib/wyUkJooBkI
cWPuSuGxrZJSKZruYmy2AZi9jB5lVLlr0+XTigRYkvB2+XvHn9VI9MF7UMip/HQR
GBnzWrFHJUKjuMG0ng8jfaoL1L8LJjU8B+9YC8Qxli0DUX48O/n9sS+Ov4DVIKoW
3CgPHhXbqAhaNW+3sYSFKa+H+0WOFJ4Ftr7bXSGO7nXzKew3Vju7kBQ4Px0EZkdi
0RlnwLXmNA8FoHBYiLSsa6sa7cs5tlVApkH/AcfH2SOEwB6c55kQJuwBNJiMmnC8
r3o70rdqhio+GAq4ECdc70aKJpYI3vmjVypr1vKfv7q8LEPD5PXvtxRNhQH9sLgb
U82KBcbTS9D/blnvQYHJEwi2mwVCIPqn05vnLGv8BLJocbJdegiMflP/jJ7iUR5l
eDWcaMwUqx685S6CNwBbBmaP+dn///WPuQzyaTuuMoy0f68aC2JWRQRAhWt2WJEH
styohdy6UJ8OS3AMR1ejvPhaUlIz4xIB8TZj5qswRynLz4jFUoIha0uzUmJSeeDE
FItqXfOaw3nZXtVPjP0kZMRTFJ8lbt9/epPbPQkAcEW8SPN6VR8uWxR058Q+tAhl
J19jXXBIRNT4z1tfjDxLjP84gSvwwapacnaiRgXFHQYpWvE6bRSGtJX9xFrCkJVy
I2q1c04EZrritK3SMNdBwqtLgIeZNPVugkYr8lmzbbexdoZlfuomSafjxTTJmWle
fJXI6b7IA8NHWxLABKh+XxGnazmcfnPWOrEDz/3WCRBoeZ/ipwGnU9BL6+GLd0+v
6haqV75N0emUorODVeURFBvSmCUjBvZVD8FN6PPppKgLAUTl7dxTNk8G9pmDeenw
p0tbP5UQ2+RJ10LzJhI0y45vd1JznwSBBfboICNLgf9Zp096DP50CuwVMdcjnhL1
LMvJ7kmFYHs0hlPxclBO1XsmF7M7JJB3HhycYdNRWjgYZc9MNhsGQu57iljBUtHL
z4Kv/HztNXcrgSWwxA2tVzkkVm48W7U6p6gl4JhjjqiLVao7AS82lBf8GB03zJ4M
k5OaaMx1XDTZOO/APmHdAk4FVTwiF9D4y5Flahz7nnwdekUKCp4hQjdetPEdvUmg
P7tqGEkOJrcCVMDTRgv+E2qNmP6Xj3sqtKxv35JBat8Y0hgOCJC65CotaYuth173
84X3+erJNoJNWhre4kJiBWnB+EVBKOCTMczHR3LYLNnafAfhO65X3CJRZZJCVDj0
EblUliGdUZJ4RVP0TwlzJY59Yr6WReKaVAFcNMYXQPSuvOgTNvafLfowPKDwwUma
NrPXVx9EGi8HbhzbN4F3DnohVM+v2mG0lQTT3eZuzIu8De1IRA68YC04HFEjG/AG
UWRrGbCXh8ln2ig8QYMkmGKmjNkWOmHVb8X8kopOtMZk8PpB3OT45sLE1e8A12lw
UoQ6M4VsqZs1ZQ3spgWInguG9S5pHjG7am5Hi6yBi9RqXavoEKyoCdpBl/DBu09I
dPbHdEOIkO+V9ksokcBuxkfVeLwR1bnrU9DQE5dnDcSEBxUDZYcWsHI0ya+K8RVD
z9QIOT43Jv2fU3r/fFplFpHsUbyK06V0/p1MJ8ajkf9hL+/FWq2WsCzpMj5J/8Yi
Ln2n9EKzK8PMVNmYSet+UqxaLZ2UBWKSar+fr3MrrlVN9dNdfJZUzaNqaZuJuRkl
VBcM/T7lFmVUlPooZYCnq74s1Sf6ZjbztYm2WKeuSYgDeYBUbZCRXBNdDEm4/V3G
lGt8/SRbDQdvr1ouCOpcACzXvHL6NdyzKxiX/nr4tg4jO1w8hgVV0RqUcXfmkiiv
OuBvMNPDnrxShruR2SSB76jMtjcC+MYz9PGxEodphgTQNYYZlSCtLBqIXg0ZDqpC
1i9D2lTeUvacxUUFf/p8qu35Bbb2nhhhRJ4wnYtLHNVEGAVnyN0mD9DEGq0MYyEl
HdGiiv+vZ9w0bRsY4OqnXrGBNbTMeyBLVBvn9M4TPUkBPIa2T2+H0zfAVFM1frsV
L9A/+TV+a/Vnpf8WrBxNbLixrX1Ute6RmS73udXpcBrYqYvHhSmo7XXe7Q+IP/Ek
g2AqIJ2IKwm13vCL3ZZ+/YUrQYXiq21SSbse8ahucZSGY+2lADJKtfT7pVseEkYC
yAq6bwdt2fzlpsRWVhCF8O3E3xiao3/KMPGaYYZGAKszQdE87v9nLrqQyPpqcUXS
bPaht5Uup32TFAC5LTkq6bpIkvAtg7R1HHgzvANqrsnTz6RwH9xHRf+WORdYR1sp
9VmmVX5KmZKKBwZa9ipUlmOATAxwJ7s4l+gwfZ8iyF+VG/Bpmr1hc+DEBeyHg7h1
ScCAYiETeHP6cauyjOFD+KRX+Ef/xVDrm28TIzh+t7eVRMByzHnf54e4ZhL5tExi
WtFh0dads4NG67M+hbfv/JwmfEHYGsLa6N5Rn1jK7l/zQlUgzrgTIG0WaeOwhZsI
hX1q7ojZWzvWjiL4UYFou+hSMHQ/4y8uCSnAwTA8BLEioP2bMZmZcEp2JqZFg6Ul
V3veFZCSW9sONwmyX19hv2iprF6dpnVbYAFp1USAbXxURW64vfVYl3ABK3XD5BIg
qUwQdebKs4eNDv4Pb4p6UD25Kqm8T+E/fh0aUwbeQ76JDyL7QX6ubePYf/CGssSF
E9AMb1bSPrHGizq/1l00Mu0dZbGpPLV5z1q6yeIan0BLt5TSweT6t1uiy8gzOULa
WW+5GdPpq+WAhwV15Jw193YYB9N3/fUlagakHOGzh9RNIB2VX9AYNMJVmp5E+/a7
gVKpK5Y5e0jGxAYgzdLCBEPNsnnEqZK54rDutPyPcCE2qseuIn8/YjP69Nor5LIt
/wKGm/hFTp4J3t4Sisv8iyZBj915lvi3VqjLD7np2bv1dokytjebh7q5VTRe6tQ6
Swhudfm9lZ7G22DS5+29cR2/BkoYv/0kujQRVj8jBJFG23f/UCzP9LadkAD0/LMx
iN3+AFlvcKYivEvZ5uuj0/WqceI2ciz5N5kMIBCNcNBlt9SB/thv0zzBqApuaw9b
MI09jwXnhqWQC1FBVoDuDFRk9WPnrEzgY76p/Ss/2wfSrNcrw373TxAQjP+cHG1a
aPABIyaO6Ojuc+LEsbYiD3Q84ceDEJic45ImVrwGY6kS3mtkTNUJ5WTSOCTOqkI9
+ghyMBeDoX79wiAyL76SCB6zpxqTn6dzE7D5m48LUbIGfOEMnxbcT7TYh+xVuYMq
Vu4UWBaHaigzNnX3aAUmHept9EFElo1BxePjneOUG95f8hEDTLkBxHjBsjqhHR9y
WL1exHYyqEKWnWrZ4Ljcl6xZn81T6cGlTjnee/llK318EiVAITW6on+QKq7WJME9
HEpeAkjfE903gxiHBBSX5QnGfI2aSSgrT0UKNUCKoXfd4urLr9eHAWC1m7PQUCYQ
0pxxv7u0jqSP1tNHx4qSN9N4dOcjyr1ER5NEy+GPkMtDJJ4OXbyEM8V278AGraYf
VG/WooxsYdqgbGPYeCXmBYq7510tVQetW7PUCZuDPFtLub80RZNWO7MhCGM5u2wJ
hgkmtnk8YvpjHzcvUTAPKn58BPJuuQsgsMT6cJQFizboYYbzPjat5wpgh+XCtYin
JjeHmbjbTo7iXYR+/zELByGCNRGvYzebFtYSG9njXQ9UCgoArV9N/IMmEfFyLv17
GYdJuXii4Qac5B/J9KritG5+sg6dGXcuZW39TQErNoGsamZ8SPAtgGfXSUPJVm5P
uETaYQTvIEsqjvMPI/cKUqSTj5Sw8Dwg+lzu6YP5fS7CgZmN0theXHeylty/VZVN
N9o5vqQSvftaprxjOa5oS5xKPUonFQK9rQJ4hCF1zvKRncffh92dWjHZQDiUWBF0
wakg7WIwzfVPT8jZLdiQLA4nwBgq5hIN0SP5n86mP5GAOdd9EY6HWZYqflnJE1ow
QkWcZeTpiCLGGCceczkObCml9KvSHDWDOl/PLomRCEy7MDXEHEcWblivqGqQx5pc
1yaGN/szxZGhO40IgskaXJiIUx0fnLs6+ZiQW5MW/+S8oQfkPD49qrT+KD038ghB
nIWQAMM4i43vS87JjciEenfsX3Oh9+iHZEr/CetyUtPvqYJ4C5qOhNbm5dlkzhYk
yo2s18wyfIoYaswSeJBU4tqiXNqJqprzM9ypIkJmGpqfAhTr+X3JL0hBla56ysom
kSzeGAi+KG5SaRZDsH2zm4djg3wsi5j7Yeppqpvl5fBm/tdMjI22kIZ3WqLIweCM
MzjT+dIMpTlwsAD9ZDlcWsJSZXKH+5HT2AjGYA1yfrg7QXKyu5C9koXtxmhR0mvy
/Nhejy8NcywET9zn9KCI5duuu0eydjuDtiZbbDClsISmvXQekhpX+ISb13OxIJDN
q8fFXwWkK2rkJPSA+C344HvLwmamZ3F3u80ZAJuQ/eZm80ob3va9vw1Z9ouWw5Cm
H32kG6OqBVWlbXAnMOC2ElLEXE17s7mEZUEbmxHxjWwifFEyBKT532qIa6ZcEg25
OQ8ks8E5q1P1SeOeRIlNAurNP3UEdVaJXmMdQ2W4mK8ia1cesRTOQq/8tKZkyF8u
yywig1eu9MMGRSEDeCRSaqE+XNidAej9LQkJ2w3IFh3PY6j5SS5sQZzUhMrBFMKt
z8+apBE6jHqCG62B0f30MMonOWurAcAVfWT9ZZlU4AaboqrcS/PGSanMxeAaGU2G
j7gm5abVR1d+dVjq2dWFbwZTwzoCqjNa5MH9K3s+nkMB4e1K3D9aPRpkcwyc/S29
vaFyb2U30/h3ig3yJpu2IidCjjCiDtovoOaN9VhZFVHFkOtfbRf9kMJgtkQbIDK1
BEHSmJCV+RiiQ3nxhz/oZxW2GtBo8o2Nz45slmiAOhi2A95dxJFdhewBoHg5J76z
USZ1rRIoXFvNXASvov0Omq/gK2Eg1ZvEgKxeY9NOjrRfOBuGhpXU/9PkYiX6Nvr3
HmVVbsalFTr8jr7Tghy6uBJxd/3bKfPE/S4TUWWKvFGeDOMym+ToeycMU/CF3VXL
t0ojn7COL9SdmF79Kv5kjJr59/lW3fXxF87DmE2OiEUqRWtQZhv7GGRZS3Has2hp
dujf36yhxmEKlwLyfAryauwPn9n5b1z9OgRtgqSmrovcD5Ru23j6NahyKTY1S/xj
QE5cXOaH+9pmg9NhN05MPUyiqTKnW9M7vu7/PXMKG5IzD8/7XQBQIm7NbKHNdZQT
DFzS6t9befu8md1BMl77Amz/b+QYTQ59D4rxCUBfwdM7LR5GwoWflNnNEkF+7H6z
TSufC7g1Gh+TWdXgrUOZl+fP+aBp057mrd2gdAFOeq5Xx6rSanMtd9PldHtOUy2V
vPabbI/CoEqzxcOkYd004QSer/rGbVN0pD2l5EN79C7RlKXUtj/kd0+OTIfujF3s
3l+7plqoaIzT06+hea6NQRchNCQz7umrr3wusLt1Zjrovmnx+dFnpnU75MpKcCY+
EKrElWuqPE/WcgQxqQlsxevfBrDGAs0nMS5oHbHjP0RIFsmsnYDPopHspw5l1+US
iW199pBDg1lagNfdFGyyr3K+2JJi8KUeYkD8GIThCCZgl56bbnm2bTWIbO6q0SHJ
AJu+EqYQkQ1jr/9blO9RDzxmhgrw2U94Pib4LLIPaBGhcOe5fzMuhaiIXBSnkKWq
jmFEYVDA2u7Tm5STNqlpdNLcxMAlNnNUyHabQcgVVTv0AcsUjxeKbjud7NQG3hV2
DorZSOVI0YSUujEcQbAG+lZ5D5p66Ie8+zreVrbKPiX1QXGw1aNE73u8p1c3rAYk
2wiwJ6ViVGV/mkJ8lRO+bTVc0ZWdR106IPCcgFEc1H7uLq1cnb1RXNcQKFssv9IM
9vh/65EhOXj44KHgQL3OsLRKUMZYMK3I8xDM00CwHNNZrGKaTgcbLD68T074vReN
SMi6BzjYcGDHBpa8knpx0YY5xue0o/+OAESakg3eR+r9v0Ig0R7fNsnbYBO59k+H
qCACtiXesd7bQ8MTXodaB0oQcUKoDtSrxQzkHN1YnO5HP1mW69BbEdZAQmhqpUNc
pV8pXTovXflkMufBPRQcRI1yCVM9gb+Rp+rtRYplWo13XPPSYgd907wkeUY+0I7n
1ZII3em2GslxVbtZnxJGJd5XBBHDP02h2MwcrW22ODcfLDEweSED0h4/fKijXeWq
9ngXKdZoLg6it/tkr6+JdCLDtek1oHfc6SKeMxH7RiJm8iwQ+z5U+K9GFxeJGuN2
8kQHietxIwEMHNP2rMKqfB3RrxINcgqfnlSTwXgMKup5xLHc8TfViuQC9Yj4/aWZ
FMJ+58hFk7cJ6Fl9kAnnAfPugrjXOjMoPqd3cMOWvGA6cdTkjxs5ndTiuvCxksbu
fKj6QgRUrfjpYdk1fUN+KjTwy6qIabYw0ehvzPYnEHSHZfNRJEBV9t7VZ+RDF8lu
6MJgpG/dHehqfMWDzxb4LZyi5mRQQwQ1XzJkOwRU/yJymjNr9EH+Ob8BInhwcTiC
bV41kshdcZx4kjl7lSIcQbZ9t0YKrDlkdvkv2Tm/aI03zLEppx8ah5xW18zhH7s0
vmz3q3jyReW9dKhN38eAwoljdxTuG6GDBAPAfAevT4UYAiaMkFY1rr6BQiI9X9e6
xwxwB8G3yUEW3B4C0Ps5rN1U08pLi1Brk4m3luHmKiIbYMsqv5wqe7cFc+6SfjCu
L8SEZ0eoZc4fJZ6JBknte1zhTuJB2rG4HWzkaiD2P1S2WbYGxJFcoZe1/Mhcwlqh
oTOM2EM9sSZHbj5KgGTgABZbIgBItMRSB8M9KrbfFF4AcB2+zV8/+tYnKsRAHOuj
NFxTzVFWBCh6o8GaVJKyuqEbyjm91q/sSNnYpllUVlRC0OoFxo/RQylzvG15fVtJ
W/daDjuE059ocgcxzSo72l7uzvfKrfP0+ZdD7UwvdchRVwGoVbvR+wlh8Y0baD65
Sv7ephtbgWPSkFMgrpAljynHrFM9HYHEzqD9Q3eWNse7AU+BGeot84HzfYolMZGl
USw1ysufrXBKacEQniuGcAhaqc9SegqPzMlOE1W4wdE97Beb80sLlpJ7myRbAx+W
CQAC5m+bn+gcoUCqq67AU7JT8srN2EK1zovRhO/Od+naiSB9tHL7RrYx7O/dYczp
AaCNxUvmOe6FnjATWArhk5mwY84MabIV//ZFG+PIq/a+PSI98XKCOXcmPdwVWf4c
+6A26BJA22gwRgfZM6iub5aNCL8skwHT9e5iZGaSbT9Ir+fIbq82lnBuwbn+kehc
lCkXgM14/oXN3TGrTw+tdt+VHZWHRG8Fk1Jljx5sDPqMfi42BGTwqJjqjkpQl7e8
yiMtV1oVtKwNz1wyd/Lw4UWjXTnvStMhvdXN1moyK13NHFUtZ43B385SNtamXgap
si2DrJlicUtoPltjdTOud55aoGkhBui9ODJBvpr1iIxpL4ks/teb+imdFetg7Jm+
DhnL1P2uvWlN3ybgzW05XrUbEFllSoTavwN+SLnc9oH24IdWmFmrKyM4jhebimtN
Fj9RnDOoPM5dXmvEo+z4nWL26G6GES9L5JP8jduI+5LY75CZEFDi8LVY58BnbKO6
KyTZ7mubBZhuYTXa/ud9Y35msWB71hPztWbQtW6wU8CU+C9ESW6ggiTN9pPeamyB
J/SoKj4eTN2X9fyQ8qzsr1x7REURc+f6D0kLcol8cHmIe+/iV7843dxCVS1pDZFE
a3mG529+h6Sd2+/hxhnuf7k8RFA41OUhxf+hAHwTIXjhbDf5nvqfZ2JESnnlJUUd
sKJKQ0ZGJbQSlSVfOrAC+5aXVSBOtjGxUMdV4LjFiFgmY8Um1kVY2CCER6cMYPju
w/qXj1PHfK0hWOvWmYcLC2pqk1hPRF1djn10jZS5XXGZD5bTQmkrcPUZmvJHoXU1
6rvv1iCGzD/jfXpdtCYLqternK3KSrA+jeH8iimh984MDApGDffYMsYZwykNCAeX
0mC172Q0fgeZLd+B8pDDTuR28xMP3q4Os+F/Fete7wEJD8L/x8VYKpooX2J5yKEb
miKAqpujB62Cnv4vM8/PzW8eaVJI9Tp+VHzkzU4XiBFwq9jFNCGktiWMEVPSTFkq
grcAC4m6WzS98RRQg3ZKSh8X/nUQ2lk01dO2NJX0162xG+w0i8yP8kp+FjWGi8C3
yC24t68IWPHJZOdSXoHFMwOv9EQEbxP67gaCbkh8jBSy+Rk8BsBAWzoG+e4anKS8
bGFOkHF3hKWADiojN3YVNctpLh86OjmCtXF5W07YCrscmzDczXK50dKM4oEUxC6G
f6O8t6DHU7IrAvHke+1p8JECsUGmGWVeWe8jzH9ubBvkj6V4t8WWOwmxuNTwHTmp
9Og79sctk9OInmJCGPXu9c0GYjOp5WxXwaZkgxAkM0tXG++oGRCV3vrscatA+q2u
tbB8EyVRA+XgUs0i63C/nvryWmIcWFTpAZQboSNPogB560AbfUVFoZIxp9sRt+s/
SHKJVtZcfSRtiHQndExPe8oyHBeE9ZWqoh/oYT276r81h5y6pgqogVoAGJWn+Iit
Exr7wuU+1L02rUsy+SuMzDSSonWKux/BsJSTI2alla8v6Vaeg6LG2XQR9SrJqVQZ
soj6L9pK/x+N70XrAX6IMLG31C1cEZoCYXkS9HmcSq8ok1aXpEY8Ysl2sGXFb9Th
Ua7oAEBiOjzj0nBVCILoxZuVof6Sw17woG4HHFJI8rT1l445lSyDverfLwonaZaf
YJH0Vx9jmFqnMEo/nXlKt1qE+DFNLj4+8m+vvg2CUvR4jJ60TCONzTp0GUc05nbT
en0Bh+Dtx22tfgj1gJ01wWHOGrp4RsxkJA6rBiGifZI40xkIxcIF1c+HAKUIL+RW
7kZaXoMjEjC7gedXfukK0Xm/YKS+jD4C2yVy0VORCKmTeA7r7X62rq7telOsmXoS
K5ZdLkjHDxxZqDAwTf6Hv0rKzDP7iGmBXwSOWhDOXOItSZw3lASc/+HQ2Thoyhxa
48ZxazdTozsQh1t3PoQtGeXUKuzMAZaQs+CetS5mAe8CvwziKSNs9RtmLR4jbJKa
DpBgMS0VWmyQRuZhcyFOyWZDSGGj0H6oNZUM3SFC0sd1mEtPm74DbjVM27KmvG2m
EASx8pNAI1TI+LkriMf3oABV/2vjjrck8MN9C57jUUJCoyNChMPNjjVmNZZpkn+7
/V0aY9s+MdSHgrUUdVaYvDPDLDYmCkQXO0WFY1Om1WG79Xxt2w1/TuhRvbAWfDSN
GWewbQs24VAkoY+zqqG9Nk40PJaYl34HKOkDp38L/0MXsy4fqUIlBVw8lyk/MMdl
OXc1aJErkx6BzGhAKinDeGEBvekUU6XmvCb17lja/WVx6mF/MoiEvwUyxsVnxsl5
HvlrY174ApmDaKKPYablCEVkqJPO5PJXWmAV0r+6rDVm7uxFbsP49MPE4qhofv74
SYzhOznGOJ8OePmczf+XSYxSGSdke+gl55PgwmZPWp+JyGM2XqYPpe6GExmLN1Wn
jHlyzIi7TFrMQayUgTQetd4310RdciZulVH5U54FLdSrT81VnhoTrL103qufj6A2
FACR0DqrDlj2TDa7spdsOl2XBhKFyn+BQKJ/DMABl39j2nXoGIJrb7eZnRL80LYf
d58ODTCmUl2q3n9Aq7OPqT5mbyAMFWnaTU90U03Mqs1omO1Ld1PU4Boo+A0oKKnw
eBoyMclMbJCl8JXrtbjhhK3R3FsO4/ryfUHNF2rzG56UZvSBVRjlFV5wkzABmb1n
uneXTqVcsDNoZg05/KJVGxWj1EiorzaTOIsJGA8pCtSHJq9glkRP+CUqUMIGqDyj
a/cjglEDESwyzcm42h3pSNrHDGVgdIqt5ZxeT88Be0WljM3QRx6xyC5n1XW9cges
BJCMtLAv3iKi3bZBzFVYQmQ8AcnpSInFZtOinC3P2b7PBCoOS+ICWNaD6hE87t3r
Nn4V5NtmG6hmLkF6YAEVe3TmBLsSqRWJy07KwmKHJ46zaMweeKQWblJ3MHaMwGxN
iVHQ28KXdz5aXk/QkV7fj/ICia6VjulRFZTLJpXuWiK18le0z5Zy9PGAIUe21oF9
RlqYdeacSRvMIcRSM9SP6i2AgsZKZsFuT82TjdJ9AlxlZF+4OQv2bpEL+KeVoesq
aZx88faf7VEaUdqqtrn772+fo3JCJCcw21ky2hjQf1SAMO4IZu/o/BzO7kOAgto6
rJ9JYZ3l2UlahgT6v3d+iIzGePBQH25PTOoiWwB6xQX6VPXW+M5WwzZHob94g9h6
z19AxnNQzibcywQZ8is4bYI8AahTymzsrTr3weevprIB9LMSvWsMMqLdEsRnF89G
sxjYKcHpTImTioEhwxZ/GvjK6cZ7e4P2wu/8EvEmjuqPNG0d8xmEo8IXOr/VxlnW
qBPANBb7YEnuAUkRE93WJu2x9q/Mg4HNRoqf6BvsEoz6MLeQACMKFdHqfpHMKdfR
2LOpQdGCt1yGu0NPbVQgO6H/WsRCTntvvCUaYjD9/iFsL1e8X4yCW0JSfrEkDMjF
yeoQND71l5kcq9/z2iFfqFlk3L6Cv1sEmqq2Me82K31eACzf5E5T2lugvd50TBxb
Ma0W1nviq4PNW0EWCj7mQ58QP9Y7IUqbxH0cQ7bdlC5TMaA67lNqVmrLzh/Jhhat
hcxpo0x0mANcdQ8A0NWq5UoA3CrIJEe8tHjSw0OdRdNwe/4tfAEI5BKQTVnTrh+j
gF3XKN6JEqoUqCcyfQKkqsCtmDwxWj8FTBSnCUCjv70CvMwLbMgkImY9jiaA1Hwd
KqhvQM03+0ytRbj7HTXJBIn8RHpOPIf7I0lRiYTYgOhxZKzozzRIKvxDyYccCih8
hhLBTeSFi1PmvR0xv0N+8HxXeUogDOVRV4gWDnH8Khblv2QJE9RQMtPB2Soks3Cg
zK/cg4ctdpryYeASRr9gMciAcpaFQj0FEXUpd+FmieeYORnmsyNdP3z0/Q5kgCf0
+0D4Va1fEt/LA9fiKbV7DhQQYxwYXBZXJ24Dja01uRv9SQmMrK2nYyFQX+ALO9ka
z/FsHGxqY5pUbyGB2fW9NZjzB/DHoMPKDnW5eAN8Ori+m0gi2niVNdI9Gi0Efhqb
2J52ieFD/mHLtXQb5PkZd1MD9mVyCXd6LZ6rS4o0VcweoBXa8IYcUIHNh7Dz9KRu
G324cDuAaQyrae+hSHD5CQ9MHn9mt0i+BFAdq8uqRqChCzIgtr6IOBcrY9PIGXC5
/JBIpuK6Fqdfh7XevWS2yB0b7D37ZWVlHadg/IPMMZt8jRuN/PJJ0wFdXi1OthF6
GpFNNJ8Osm6XQ/+WYTgBJjsljOXH3bpYpv34hlM3ycfhMgHi3BTil/S7IHro1aEt
XY09qVUQTyHeDaes505TDskSKL45gWmjoub3iuBLyeAqCEyGxh85OlLa8Mn6mG3C
49KIMhXBlCx5EKQ/8rH8FVlHIdgUAm5995DEwebuoBU3Ymhcx7DdaFWKDZGZMOvT
GBJLs+x2wVnQed725jidTDUtoaFsBYrnww4w73PBS/U4abKA8tmwVhLEsKF3yQLt
xTqv8HbHUOLuq6/Al/0Rf52c5+lmDZwVkcwmQCX8bpfecKWXWMXBVw1RYTQ4QjAE
YyazgxEz6GHt4tCt/oigncyEjZCOX4yhbM89/t9FaCGJOi0xQ6UUzexGlc8NMHqp
/X4k2zVP03yA7QgAa/EDxtPAzgZz45jqieOrdzTSWk1SF0tRZ2uw/ssEg3mn460A
HdVOodxd30Z7XfC0vDO+02z7lXIQMdk/VSULKOYVzVs1o3Gqxn6t9HyyaUvICDDQ
iI/SM2NYYJmTH0/CqA4cHnnqahJv3K9kfltvj60Us7mMGUBT9OFQZElBI4GexN8f
Y3Up/rwhcAbVFBTHikEn0lh2VR5dhZ2BjYRCvzU5Ju7LqeweygAiN4P8mt7KwiUh
cnIJIphTj1z3AL+bV35z9uGPhxbTMqm0W/pZIb1JqIieFfdznRxkX3Fh2iUcbcJo
tEoQH8we06QjSZgxlu+a53sAI4c7LkAmFMx8AfnnF1yhFRsFe5Z3xl0dQ+zKVj2n
FqeJLKuP6sDm/yzh3SmPTrZMMepADIP2A6F/RDgu9QqIatLJ5wGnyZ149YiLrfAb
78b5Gd9oO0ShjDbmg4Pt67vJ872WM5soVbm/FCKvHLOn3xWjXWQ5XZQPMwptTPQE
3qXeWGP3/Ul8ijx+7o+RawsrJl1xQjeIIx1QRUrEwpfWRl+XFbMERw6rKVw5dzjV
wHr2ROxks9JTiOBTtJS+3m+byanF7E9A/YPgezR6VWBfmwbN3ERkHROmnGyaEkoW
f+vZPks4FlX5yXrMqXoinOezSL/XF8v//qncQDdreKxDqjJhSM+xIcYsruY5K0If
WGgcDRuRhiKaNvYnYpXYpnOsmj/D9OYRI7g4m714gNDctd5Sun8kPNTd5o0VO/vu
bCVwb1r4csP9hYXqV9eGv4ktD8gvXfLIUtqnogxJ1dwgMf3cpgde2wRK9BgBbSO9
P7tW5XfSqcDuAkFsFrP81Xwh+7VDwRpOyVOyzGZPiSuWnZAzqGgGyzdguKHjjcj0
MypGN+pUhk/IVjaw9xKEBO9Wi8RTMgQf6Q0oXgVm1Ynwr6BVGO2bbjgbNfbg2DdF
3llF+L5m4EskBoGhIYwdSYavOBEFDQkw+MeeTgwi3W7YNDmD9eAi81D2W5/Tq8zE
jEJEYsMNJP53la+aCS7pMRRphUcIp8lMpZORfG2HDCTWD1GO8dLKLc7SbXNOyH9W
qvfMxT5aYcssgTO3I07SmK/hZEeX+AAebSI4ZRZtfHKzXpejCokfpk2eSQUe0mmi
qWGo4v/AbpAFK8vuGFg6Y1Tl3HoeUjj3OX2rpBaSSqrxJneeU3N5pFpTd/XVpt6u
10vgOF7J5aWjwNkQ/JfMqvc58ucS/jUUWawxNLuO3R/8I99J3fxb384PlqwGzTId
KTr0eOFduLENgGVPfEb4HCahtFkaccVLbgrh969NPkmh0aK1QYm9gBx6gO2mEPdz
PZjdA90iebWb1whwMt//TI+MgyrZoiVeRqjisKN2ruB00RiKFWVPoQjOt9u4157I
u3bXQcM1HYwmgAIAChVJND7WVeFTmNxf9MKzMFaa6qmzIl5oDcixhmpONNGuoy47
z2OrJdXCNOCiDR13t+TdxGKo9Ag2Ba/+EaTOoLNV53+7PghBTCSrCmaiae8e4ltf
tqj/xCT7bXgzV1kZHJ+WGF6V7AKL0h0bbQboHO9gAx+ssGIDco+zk7sxUFlHem+n
Tp9FYlfF+0rRwnBPwLTrGVWKtcAFcuQUB9/cSXSuakIY9geGHoMn1gXKr6DrF6tm
jG5f0YfHgYruoWBo5jLdZzighogAGH32uxf2bNj2+leEo5QU6/EewEZfEjudhieX
a6aSxWr++3n3ZYgrd7W4i0raGCRVoM++uV1yMd0tODgz4oyL2NUqnOQLC1aD6VXv
Cd1XErzlCN/h5m370PwqtjYEWdqCN/dnpuZDgSwsg3PKAi8tqU7UVSbcX0bBj5ZR
Z5J8xDUfoCfm9gH8umgqRIUDmTLkcQJ88MpflMCMKBCawM3eY2Y/v/npVD6DYnOa
DvU13WBoNGFVGjb/Va4zQTufZgLvtVqGfDDs2ChNvb2maN5n8++Pw4LG32sTEfbv
l/lNVYVbW8VM9f3pS9cRhtX2aJmBvJPEP3JU4EVXT9i4/vTz+xuKuf3uUbl85aG5
cRM0P4+wCJ2YnLLtEWuGKnuxBdNvAGvpEyrJmOV90Cblj/uKPHnr9q1qwYHbdFXQ
8M7jenm1gxWrJr2hSOz6YR+LYex6BkIbebzEXJTeR+UWDzHflK5J4gi8PKmgg8fF
oPS+PX6BXXXawzO2L9yFyVyn7/OsxITfWoHbjadZ6cCmzzXvzI1JdIkX5xPs9OjR
l8TNqI4sZ7fWY1pU5x1KbAhffEIghlnbsoumr0665UEEuBBLjYkvscmM/p9G08IB
YowMF4rnOA5kWWoW6zbePScC93fMzZ2DFLRXw11TuanvDFsSH+oeTKOLGsknihw9
YcIqkmLT3P/p4+MocHUuFUS5eTzUUule/N5NL3/LijlYkZh7v8MTV88qGw/kZv1e
dL4/3zWDMkwpWGFu4qjQ1DMnOrNevnSS+raGQ76RVnJrGQSIveRHbsYXb19/X2Ke
hGXCZgG2zhgkmgY1SbFOV1F7p+jzHHFdtIHLgkBtxzOuf6pQ9drqOPY6gldVJVR5
jKTN8cCO7KCpnWjzuLon0DE+36q2QM+0GWmlNxb9lIbVH9Y0JYjsj8azaDxwXC8c
vcAYCMlvpE3TWWTN/iz1uQ/3JRaMIqc86JV7VAC3ACTt8yYNu1nBksG4CzPt8o5B
d/tscoq7xQTwjisvdIlOID81OSjYHkKsyLVaIYn0pQqmK05jfALLZcyTgSJuCIFE
AdTgIMpNEnqmDv3ClOGfoSGxS7XVsb1CeERc0EJUIrDm5kl2eaT2RgKXhm2odG7g
sYFyHcJloEmZFAHxLM0rQ49jlKDlI7MZ/4OcSpTA+BvjzwyCzl8yVC+u7YEajiCR
nGvNIT8dWjazL+D+PbRX063H8SrsPnPbAMe+Y956hQ3ECZx/biwBNAaJd2WCdAPj
gPN0lu5u/oJrCN/csG98yf/9YgU87JTscDag+Oys735MeWkX7TdAhtWDQ9rqvr4c
VZVC21PECPPoT3PlNoQaXds2q7GMSEV3ZVKwh99E+0/Vo+yvdEmxGX5GgpYWygvn
ImTVw5v6p625RFWH6fnvf7Gyys57wGE7r+tRVRmtntIUO2M4secPmXmEbiMWXpfk
AAFR9WoBdrv39NSuqvnVqZOerUQ77CpoUJDQ26fPiOXBarf9F841/m+IP03ckCL4
4OiFlhT65bH5oGhXKVfcn2kkxCYvEVSH8VEvvQfnpwIBYlVNspP1XOGQVHDv9Czm
bed3oI0C9rS8ImpdzE25NM53Tu489Z94s6ntVV6GW+1Ye8XJ93k8YOSomR4zIWfC
A0Mjmh5EpnVJKn8jfRcGxgGAb63GwBQn4xwwVFg4dC9+urM7+Jvd2pbndf68+RUQ
j5WDH416XgFyiphXYUTEM4WeIRh4zf1M8TVM62+ZnZgl8WpZvgkErAkQocpCpSZw
Wgx2pbZr8KoFVDQcXaSb3EFHtF7RBuhimAkJXQHi1UEfnMyr2RxhFYO1rg4+Gui8
8GBT4ETf14x/1XMe++yKVkb0APwr66q2fGX2ZfzXU1/tP3e5B9VIdcp3xqAyXqow
BtLmAc7aGtfv6KPbeBtAnw4iyuh8jwP7gdb9+w6qpWJ0BTyfXctQ4SMTFAMrb1w4
2K7QPBnYEne3qt1lGdAn6UX9yInd6KCkHH4vXbdB5NZ7XyOEfCr6zJMGvzbL3fh2
BQ4UOchQr3xJjWl5Q+y1Oq5rTTeQ4guvldCqzBzJyRAPs1vS/Vpz16Wg8gSI7Jc7
RxbM9wYIjmzD3CwoNys6aUDj/itohzZHJW01OZBt1NELRVrRvELF9/Uj8yas8EJQ
JGABjhc/9Nnc5zyu9yRV+Jp3XZ4J2zNgmDAxvQ4dtqPH5HX6JbHuz03HoH+ujY8u
x2FU5rfqpGvLE26dB3g5/BHjX85ozAXMi8KHpoB8baaltd4153YPTUN3HlKmraPK
zmG6pDajBpfzSnecrZZvLSloqAOpkt5mzWfY+RmbAvduur9sNLHHGWppq9QA1W35
1UmE/egs9Wv0p5ZYB0Okpbcu0unLtugCLz1Mefcoajn4+5q9jccH7yyV9X6CkKJF
YWdcMY1jpuu1DB3fRpK34zOkBrFoJAnZCQ2qNPCXXmcL2PfVHIYbtiAyU4GHhaBX
PTGT5KxVp1Z9R5Mqiav2TuMJ04peoFtSNGIOECopjOs2lqrOPV+KUv/7j3prq8na
lJtN0KMkppOsMtQzTDHyFLiU+1WsZHIGIQDw8Wi3uh2GFzgxbyOAqx8mOP+ytyDU
ziVXVQh+GRUMrNH9nyq2Jupyj2OFHc3HQ5KuUReIfyjsWBogqzB5zbnTq/rTe94S
ywEzmCLogXHj41iaXcM1XUyU8TB4r6lGsT4UTFRQT7TYIHRS/h+dPGMbOE905wv6
1SeHM+AqXivCFzPXlX4XXDxg/r1tn61jUs03Ap6tsPs/xAs5nX97pOPnInYfN7LH
L9ogdBwkoe/SF58hafjHOP6VbXF09xYisnhyZypCpMC/twLJbmHjzrcmLXkMaY8j
y0OF6egO36UN8trGG8b3OMKf+g/TMnSxhf7x6bxnCSCDw68tMBc+aWyoOGVSFoMv
e3i7Xkpx9iTMwPOtk9Z1fQ7EQYrhFphKveXoO3kyUOV79ihZ7lDOBJ3fag3Ef22Q
iFHbucbdlBuKEm/HbcIQwRytEJ1O1j5xMMClVLJM/e6xc2nHNscjPmkXLFplXr6Q
TaMz7RTNn4knG8Gv7gTQeM/nhTiPMVquleVl26n0MVB0L64pyevJYd96i+OVEHdD
zVL841Oj4Ig3XCCZn64nJBa9+nUS8ARpzMIiEb3GvL2cTBWz0IPA6RMw0CEb+ZsU
NJhs9XnaRVLp+dMQyqR78aq00Yx7E8Eqi18Ma8xGKBrzy2Xti4rNcnQ5Mvo/wSRL
mGeCgynjAkADzTeZZMMNSvrtxdguqWIa1zEltCo/4ldyrYNOBEjq2QJzYcr83Uwl
GnlKKcz8czs1NzVaDgfA0eL8GegR28Huh5VL8/Y1be3Jz3O4oDAMsR/qKk14/Iox
al50P5S5S5c5OQW/1rjytKHq94hcbkr00eDvhu7mHmW2b1h1GH8wNAogxRSJNdbg
DDh0ihIm+LtuSWgDaDtJL2/UA0Sj6Z+b0jNIIj/gmuAXQKUm2P9jBVTXHoc99PFv
RHEFD0H18mvCq33g+QNfxlXcEkcl6RhzH+gQPGJguU/W0hSb4j8gebNbp152YEKB
xm2WZLuAftpekKYDNoYNa2UHL0aPTQk76yW5SwAkwuLGUzVwm+FUnlx2uJg9NJQ0
evy7MFijf0vfxAKbrJUIpjjjZDLcudUpA/4KWYJ5Ny7B35bc17ONelwORezI8vHM
Nu8HMwrJQMTRu4ho3sWh3p7p0+iGT0gb/dpuPGyX3m4ovw3TspjGOfwYR3ISqEHK
KAEs8IwTrpXy3os5urYZrKr9HqNY2EdJ7vIeJiaikjitakJvthh444fv9ewBfqqx
TvZbGcObIQabCn3NO1dtFN35lwluAtcpJ0GrgSCY2ycXOe8yckjDfDZtmFfetTDe
qqcm/9w8xBHevXSw2/snyWU/zLT86zM5oCA8PINz0JqweTuTG+0fzp3IclOL7t9t
p08WXPqJn8EMA0VA5jKdkar5UuRWBznPK1pzNQP0xyNfYgk01Vd3eYm2lo2N5g8Y
pQTGUh++Q7xHXnVZFvjAPLJ6IYLpyamrQFJuagpoHI7PsncR+xJXBcQMfZmOMU4E
fLwXMqXqwc6EkJXS16NWFupWMOS9YhTKEMz7RE4NtNWYkgYai5pcw0dvUcAba4uJ
s0/YskfyyknnTlE9TM1uRO9r6FGFWjvAhZNfRyxx3h1Yqw2y81pfTX3wmVt/0Aqn
NhycVpdysumg85PBOfF9yRE0yjWTcSR/FcoLZYt5CgDkN4ZmvvoXHT+VV8Nu9o7t
vSpCmuEp7KMaML2Rx8IxodjYwn02vX9eVSKiRsJ4idc3ml3fJzmb4jhY18luoh+3
3rE2UgG94tFkOf1l2jp52jf7ctD4WgF8Wod3OhJlLMM3EjdtMD6E3T+iFW5j5cWj
oQuXVhZ9K6Cu6ELWx82G3w2qsGSx3VgYF7JuDtb7UIEhdRG5RHumqMHxPFD1LyP7
G7s3qTK0nCEZ7oc18q5EHkNwhPe3/W8PSRZ8MFuCSH5L+YpmWWf5UNviL0lkihM2
GqXrHTk8Iq4Ta7jyVBwdwtxborfMjyGjR1Tghc6r1F423/1RIlNMzcTZ4uIUh2jj
MlYDroXJ8lw2F/8Yr4MukN5M8eMtIhpaS6zuY3L6TbpJtcwOQqcnp9/u11Uy0W5r
t0c5eTqnYRxJ9mZal1EdEM4f1FTywH/UWqvuT+QYHgVgwXcVylCkI+VgupKDjcX0
XpAVXjW/F0QUui9h2vNIYw/UPSGcdvLKosxUhiD0Cz18ypkhdRTqC2VznxmUJ2aR
LilHfByJ7BDtz6yFzYGrB0HcLEAe0hj6es6nmA5rKvXDYiQb8SGYHbk2J3xoJL5M
sqha0VTR8zPT3YaY6jDV9b4DPrIe7UROQKDH+sRnHOpNNeRL61e7Xg+jGcd9u4+0
XzJvY9qtgcGcDoRnrDnrcyOneUXJE55Vsa2+kYWCAxZHmcuA46lWd6N1UqkMDyxW
Cbp9KT53pGA3rMMnJtWcE1uCEF6ztWWv+h+kGcjocEns7bqW/7REbnnLZ7haDAVW
5HdAuyTTNGonaZDye1jJBGOF7TNn6NG2b4dX+IihkZEkc7pUIrOVbElpyNkxhg2o
/3sqCl+437de9Va8fUZRtwRXIuel39jTz8+XRx3NcugHUPOl9nVEt9wBZ869dTlQ
NZ9GBTU0vl54WPAAA0+BlOIbQaRI/3jA34KTBFUzi711IxIbHcY+oiF4+vl3XnIZ
qnHTpAbO6mibr7RM2ssmasP+wpk7dmUdGE/W7NmASLZseFoxKAxUZKqUP0oZOrX6
fZd9Jkvb7vfRxsiiUo3XrShYEAy9vfHLEHWqUkjr/6buFZxDspK2k6ay0hM30dPc
QMqd0Sc6Xk4a1eWfYSIj6ZHvRdSSYX4X4gpOpkP64wRXqAMSfl6iwWZGHBTKlZGA
HsJvLh3bQK57qwiB5UCVYKgfA2pRlECMhEnAzc1InXzBvsZ/wvX4ZyaBY0ssRt8H
J6szy5G59Mlr0ehqmHSTnlbRtqgC3AlcRpoJAceb0dJ6yCxVfxJDJnuuDOKkjQBH
2qXH51E0ygCqKSWHkPqRo4O1OMO9DIbPzUM0l1b5F0t+2z++rRzA38NBaSIKKsZP
WXABsMLPHUiUHqB7ilejiBu02Zsyb5goO6RR6LDh/lNfxkLrsZ80fxzSirp2OSUA
MOBFYv8/xqLsxIsUlP5OwBkExnPkcacwB5632HWZc7fw9oBeMeHsfucvrKShbLu8
rxwhPusxR21QguZLbdiZzI9FAGPHEGnEJaCCg72RBRkOiByWYPeY4SQ/sPk8lVFI
H8HSKPyuiV9anyQ4N8NxkPO3Xpg6s0MI0nLitaFoT9dPEDVVL2rJ6MRLIkoo9sV6
HzJfOk1LCOCAN8VdKYf3Nte3E82xHk3tjso6u39uUE8koRIbGkl0MS7SeWwbUamw
H0buZmJ/q3FrN57huf85YE1YtThzpfT9eO02m1SxBNEi7aiuaPEOmUNXQ3kOtaVG
mb489IrU0GAeoJ+CpVlRRORCfDheV53hPkVn0taHUqjmLFp8zfTGRROtpHCmOHIr
8slSmHhf7YnDZEpedKpE+AI0kkmt+XxUUiLGh9l7Oeyc0ursdu+uQD0vSCjlOgaU
g4LuWVJVJSMy9JgWUPaaVzFLvcZWhe6m3WELTzIooGcgz/9xW1c9W7TYbzrREJ0Q
3FarEn3ac8SvdXeajaPZvg2MTgXSG9tvXfgPeyIK7mjA8ybrgolYw6LSJ993p4GK
buqwc7K7jkr2yx2zlzRL8BPfttVXtkNxchtzHm9gGAeHKtg3rw05g7SL3aFm5Vqw
IY2qHTBlqOY1H6Ufxc/wny8S+7pXk9HnkA58xs4nkV2APibek0Vxzcus7msCCE5c
bR9tyXuDNTLLnT7/NEmPhftHRXXjSQmAFXWuDf5FJPaTz2W1zLIzCHVua1dGOVkj
Qaj97m0xJpUZV7HUooe47Z0QpKdsAGKo/N6c3XD+37PZmqD6OtMrfLOAKL4/i6iC
oh/IDDsbLTWUKw6hYfliBg4VGvTqy40SYaIRARWRpyW1Q3FHEYSpOpg3+KT8oryg
mPW1AtDqed3B+rUVE2sz7v/n/jn4rJhP4G/8NfO3oXYVrFp5GGKyxSNLPQvubyv7
WnG2ikeiKONYFw/8wKhcITpQQz5oOaPlbJkRR06Jz6U20mOPe5Z2Gr37IckeSXDR
tDwfbfIYdU/Y6LtMASFplwGBlGdTWC/cS3HW8BiqgKNSt400YlhAa+yed5oX5yT6
y+6LWhZmqjiKoAxcEzALF1GxFiZc1g2RyZrTGDuN3TOsYVOHIGuT4qM2LZc8oW+w
kwl1pbJpcYjh1+IwOclYIlLGntRmVDU/tJpJlRJ3j/5yUVzGgql0oLeNHB0U3Wpu
ZJcFUQHAriLW4j5sXAmE1jhj5O4d3/DXOd1/b2eXYsXH/eNFfuIjVkDNE7kW3mX6
d4tCR9wAW4q16A3TgkTayvcKEdwhAcUFN2KQSTaQugugFnapbLNsxjcWl0QQTbOD
ycwL5iOl7GGxNHJhUr3w67dWf2zPSlgbjINa7apbpLja7umkJaKsdzUlC3yrJqYQ
ZAweKtguDgkKBDPeNeVEkOTk0KhoqpFUZYqU6ajHsykOKMh9Gct493PM8JxCwRL1
huHz4kHVT0NB9KM3v077ztddFQXLv9I93NfZ/FLUhSbD36pX0B284ikygs0/YmfL
ZicTETY6qGVTK39T0YG2ZWT9klXGb/pMx9Q0sygVrqPU9EUTAK19sqV09AWcfExu
yStNY8rmrquAhGST+RRw7zURB68nshtdLbWgEA2adBYiCx6kRJPlxaPaPUaYs8zr
KUdJiwjOmhgaZaOGK12gTMUiRvAc5mjeRkNxhUWo5BTZbRo0ZMyYa0FtQCYnnNEo
rCYTgW7scf2DdajRFQHv1DXY6YxDwwNsfVQ7lxI6gnQYkywo09GNBqmjN9fK+tHd
S4AoxOGIq1GIASyG7wck81InkvZcFNliZcwS53fhA29frWUyu/XOtMumvctKIAv8
KlnP/xRF4ryE2Ugnm14nQ/9vFYYHeWPaoCtCA3GgLgsaCQTkFEuncORaIOESeP89
Bj2XtNd7DKk7zQoDpJgFVsrF9321XVXRZINc132hko0cwnOVJM75ehxiggSR534g
2lee1IWWaLRRHoiCal4kqkpKp/lwIaggvopkBkcyZ2BaXxhnan4xWR8q04mdjy6n
+hVnCQi9TQukDlpBY1hYV8rxFpl9Q7XX6bTRNbImADZuOCx1r3Jfv9EM9V5zxRxf
V6w7FjhTMX414dFGc/0AgKqId+TNwBvMv2Qiy7mcvoCF3QQksEbHzSYiXnRi1dc1
SOk4klMrGZ7lrnfEJ8qNZqXKp4uBEuZkteTzYATSAO7sgCjHhpViLh4EUeeDhp7K
nwRt0Iu1a3DxEHop/o6I78qZ0QozMxHtJWG+DTGvKv4R9423jPu+ue2ARrUKMglE
n4dxLUXPLUicxKGi08JRrL+AcMbmcGFgTKxN8/V5IfN8KeoW2Z3mj2gYR5zN10YR
Zs6QfTFxUy6V5nYRhR5qBk4PReVNGRlMFamhNXEacAUdF5Tor1omDTUVXhw3AaJh
4+aoJcTk7sXsmpylkU1dP0+ZqG0cq7Go75o/+RpmeQQpLKFi9TD3SRszQXl7QZ0v
y12U+k6mBWRMYvta8IlkBYsd+jot8pfdKywaZ+iHku6guTRqNv7oPcEcVPfLBlX/
sE3yq2sgtT1NjG+uBgm6gD7rsWV3lOZl2Rs6mLsdeWzmmn85J7NN1RHWvxSya3TG
wOGKx3ZCj5c1bV8DiVXIef6bAiY9cBSSIGjrX4gUpb8WLbmX8pnLEyaPcyXkYeTk
uK0m7Zr9yr4GiwbPVUEEXDXTvYvMIpyGVrGu6m1wJAhdCLl0pP2O2CCAL/HIcNr5
EeXYwLp586XgCD5OcJT6bHXqQV1//gYQbqCMtO1AM1R1JcmYhFqKu3fGvqhmtbyO
QNaUuj+3dwl1lRaSbKPnzPFzoR8k98wzTAzBXvlLppzcVNHB63u9yLCYvAe3RqdW
eb2b3Evb4z02us89D02DP9CJ6QmbPmpVfhR2KdX6N72J99Tc+qjmVEKsoBJeIJ9/
qkVNrb4Oc91GnP3r3o9kYaqan8rQMidN0c+/C1+fco6RzciKehhIKurUmCTVwe00
eybgr+bWuTGTAgQS7g5NgohTLkAinSrvVDYTAWL0lXwBJXGDc9IF7WapyGUaz9ly
tHzbjL+mqPmijl5gacpFkEWTlJ4Ze7at27FJPU0S8bX1aeIZtBmf/iVoiGmmeRcL
/Ym5LG3JxfqZMqv9/GzbuFX7eOd9AdepiyC6SSrMypJ0oG6jleNaYVqfrRkVkh9T
vHcG5JERVdT5tGMAKuhPYQyB65NMkAwVMsMNmvwOj4fiN99CulvswhEE694K7v4C
3paRPrdibaplMvlZM/qPa3I0Skj4JplPvkYq5kSE9qjzyUqNcrqyOeVc9KU6g7Gu
HfMqT0s2dRkYV8/gLSyi+buQd8BnDq6SPUlpq6yefKDdvGII+TmjuyEgvhlnoJDo
OppVXLcERnXfzGPxklXtYa8aa+oP5oagpej7fli9IAnZgOIx4CYgr8d+ZZRyyK9R
4AuLZ0Z2gU+kezjbZsCjo4LfbxmhhS9G7jvuPaOtj8JEE9jSgJh2F3/6rY/rgUQB
DThMpvGpkS+lHEZtJs2q6osFwE903bSAoLJVWeZh66vHaAZpqFFlNd8rZiJXh6NF
CW4Rcs/7MxPa21qTLSCSaG4NpiTl5QGK1RPI0aHdRHf0+fVtZWkWcZ7hijZyYrjv
X/VsGjxdoDR3rtb84vCTTvHMl0UXkK2rEqQqL3VGwd7Q6JsgXi6yIyl4FLwvQB7T
4FYGmCgK2cgLzRoufqx+jDU7FvOggjFv1yihpS/mYfrP4UTAAcDxiLefyuj/8MHD
RGKxRTm3elUYhnxx3cK1zOCQ0Ioq9RdG591YXdhMPLQQzWdtPS19VV4ndG6dlfx6
mW0AcjIuhUvy+nAocs3DezM3IbJwn+CZhTTv/WFopw8SjyQW5FXawgX3soZaQrZ6
o2vfergqA/HTaJkPTPTEw95TJSd3wBD/+SGOVEcRmxS0Gvn9kiu1FOFo2v7el/MD
HAiGpWuEw++qy6mKLC2TqlZ85wvDlI748hwxnBcqV8ZCYZGuSkspIsCxJIP+/kcr
JmjCAKpsNGdOqKn2BCa06+JxYiqT64dze8ZtYzhQIS8Dmndh/ljcPbx003hX1HYA
pd13YYyBqMNNsFa4p5TqFHYg/tPKWCYhLxSk8GOCR8QLUnAQ4c0Vc+QyvZy9w27A
lzi8EOOcdqvL5uRiwbDguvqDL0KA07WzdC4qwYfaM3Zzc3lOmdnF2VZhQihcex/C
WLd05kbK0oWVPko+kog6Ml2LeS4CQXIoek0R1gG6p4I9TMek9t2V8a8LCjoIgKGK
pe/EiHRQUul5cvM4pOrE/awvW2Qo3fDiu4i1+zAxAjDpwWKnVpvI1K9Aw3SUVezU
DWyH5RsRSzM1zIz/oQWso0n9Z4gyEuYnTv0OaXmZbQPAEZJaS2yDStdmvSvsrgOr
EYIP3b5crojDXXjMYUpnGzXv9fG5Ki214t6cLdizar0KCXVdI3vh4PeGQEHC5eNB
1PX62ViuTrWUDqQYEZh+U9WUDBo5SmrxytlPx+EWvo88jdmfpej0G2PWfJtPS01s
ksq0fvxShuQ/pFUygPL4hdKZkCOFCPnxQsJUW9v4I+nj/1sppGnHdWraSNxzh1xS
k7fUS0mKp01HG+4r2Sl+CNTuiPG6wZWYw/0frINldNmxYQMrz7hdDnpT+AVjjEJP
lv1ldnaS5GAhr5q4lHxvzoKJVCXKskVFofd4xjSgGqkXNK4AItrMVe8XwBgjt7UP
8S8KeUZlIFqkJw69NM5ckHxIJ0BEqems3/CDQKYAC3MHt120uNzhwi9Ksz8qU26X
++41AzKcfWGZhrsX+FRgSwaM2L0Snhq5MSDYz3bLUGLvpuym6yjbWbAulW55WQyt
ahIIil/Uor1WcI5xDYqRYBQAvWS83s3GtYrBmaXQtw0ZbVGgKbf4OKNKsLHdOcTr
vbtyYK90C/oSdRmnG5HGW4X2m4iEbbOZec7QfnKGJaEdunG0vD0tLZU7fP6CnddP
YqJKOWrDmnhlwwFMK/jkoA8pXe7jlQ2EAwB+HrEMmNas8j3CkdxZWnOZSnA0DzjQ
gccw2hXS9FyJulHaJATHyX6O+sWy3pdPguAyPk1R4hNTlz4d8YfM6lFBTtCfFZPQ
lb0zXhosQ4bhND3z/Qw/MRqhbgYdbc4gWbbLugCCckNI/PzJ86SoBZno9qNwg6JI
jpQJ9N41Q+G9iYSUYQ7VrDhdDsua0sqgYUNsr+n6GC9teEWBEfJvZttj5Fzu0x/w
XztTRzut04dXiam3ONJryGFrVp+uEMVRxdaMSTdSNUwuoKBWGQHObtMhBpm+tuaN
Sj42cuvaZTPfmLhjqKLa+BaN+sKTmSDUR5XriX/8CT5QNVOWxT4ENl26TWGY2Yvs
/gIoInO9VjeZFoDAKQDl4qC6u6rSzVsNL+B9dVZHtz/eh5ig3hYcVXTSBsMJdnjz
1dAaw+/H0E8iynVMbWtfTp5atuo6KVlyRyLiKjuqoiI4gEXuvV2Lrccxf4GyRmrE
QX0u/+iFH3hZK12pvpJU+xwmFPqg4i/KQoTsGIXiGlGxgzl9rT0FDvAKRQLBzSyk
NO+rVyjh1UgMAG2P6J51H0fGSDy8tucX/0AtreRXANo5q8aiQ0LN1tUOX3h4OC0P
oXiP9L+olnb1wO6ILA0UTwVL2zo2IEdXK4DaV2db06GAQBWemX+sfMET+iY42hEX
hYUSXzMFI1357kWUTPsiXQ+fGWmOYZamPtbfDGcOfVd1h1RDPIpKgiqW4TF5YZMg
vOv3pyXaYJ4Um+U8sLT1ufnWBokcLC8M22Fi3PvX1Od2tZtePI4lpJBJxySOYlO7
seY2zhFDQ+aNl3GPhjsXYsIclTGalPxo5TMs78SvHiOV4EwdhqYeblL7HtYG5kQs
4etMQ72eg9iM/qrcGAPTmtyJb1QOmNNgMpCECEkZVarlSyDsZbdjEJTSeAzRKs8W
NyObskvfvrbKx/u74P6srFLf8o4KZPCLteeRY9x9+UuTmJhUV/wd2/2wP+LCl2l/
QMdY7Oc11Aua+bLzt3qMa5dqrzkb4zW5z3YovfYaYq9xLr+PzVHOlaCA8J5ltFmC
FKC6T7FwHHjWt4jM/MqwP2ck8HFCZO8Nz0alWBkjQekwUUSqRxBhVe9dV/NYrmbH
Qqo8oaXGa13WnsH1sx8KKsE0FgJx08E8EPOpkC7UOwiLUF8S6CHwnCqia/B9LCdI
8M/CV6AdO1p1tYWN4heyiGKX7JV6/mjJVBB8KZCXKEd41GsjIpttIJKrJhCf2s6v
HK+WZuHV3QJtFmmbQ/b4xGYiHltkweTeak1vqI2ww1vrr9o1vSk45ifLDEdvTo/i
o5D4vrSefJKBl+Or5bzadcOnNBwL584XV0iEDzSmcURRjkl5qq95FsXD002UnxHR
w6BDUiK85DBSBl30vge7gKEsFnMIOLYuC5Fnb2FY5lqWJkHBlkosZtJnRL9/bwJA
aczg6k0o83pYrzH60iacfWIjeg8mDj4S1cHWcqXmGhjGD4zXJGmDitZZr4baDA6D
r291tC+fv5z2JiN754c8uuVRLkDfSYxqQK6fPDmVAQul6Gu3VoEmvWDDlyX2TJ0x
Yp1DOV75qoUuTE3e/c6MgJr9ewn3JlooVjFSmyEmkZR/k9eZCGaiYvCpE08RjKQ8
i6IER4pOmE5QhUOCIpzl0m8HJQO/yAr9bXFBzhPiPPcvnOqpRAq2+h6EuHY80LjS
9zr41bYxVt/grdvQab8bWWRRK7Hq/ctfgedEg3lLCs1Kdl+xhGE6+POoLsRU6Ss8
+zjeHC5nplS7Dl7zzR1W0z2+BidOUwnezEZmbvOQqOz3UyOGnRctEro1x82czMUf
mGZjeNxKmSRUGbVSkwRnF8SqeAHOjiekFwSASHXIn3n0qz4QHMriRDelwVddWTZN
XZsiadZNdFGLetYwP7IDll5bfJlW938IDKQV3K/Cqi1SSpgGEliD2InRu9aO0oJz
Xy9w7iKW57EDGUAG3Wl3n7NNnyfijNcksE8iPcTRL8rUMEo2O8NdaWQA73ZaN17K
uGzxPTZIyJEzoEYQw4UxdKgRl9+0gjvoCnH4KGd/i2yDqFqrQERSTW0UURQK8Rf9
4oeHlu1FoEL8c6NbBetJzbKmLEfMwJEWmoUHjfZ9a/6F06ziR0w+2p4XhHUGBpPt
iULBcl273B+h9SSAxwXv0NBm9kLCboN246TCz3W0V1CY11PKrH1vCLLA/0hbcLOS
rmfeTaePhfXj5xH7mB/pcW5EEXRS/5NFsLdf8ejGi0yVdH8EQ+nyQF/6X1o9vttF
ILLjOx7rLKhYl/poZ5MS5/Hhah96qkb1NE4UwNHLrQSqCTDt4Ox126T8oVcLxnDs
8oXhIGRO0kF/OrdSXLABqrVtN+5xWp7BRE2cgjEsBzoYKfW9r6XbqlrrPOTOFp5Y
bSRso7p4RtkdhFYZgUjEPzbzV9c1QPICkfF7SgOjoS52RF6Pg+MYp1u0yukCVWiy
FED+two90Vh/uj8ep5zTuq+/45oP8QadPqkYjU8lfjsrKDSfA+fOZi2MDWYF2OQ3
8pyBQ4k56N4pz5ua/p0QM2bTeSEL7YQxhfPtCAVHsdUnrWhDrR/eU1x0HvHInx/T
q9ILnbkeLM7D2BpJ9HHv9/vJkfxFuQh9LCrcYpFQmm7BwkOhfKzuca2YS8qcswNB
4nIcI4c4XqStEcM48XdiZDWZrWAPO7FkYqekPva94/iJjjQCDkRO1L9HOsecs/Gl
mAkEN04cUiq9EVR5FG2IGwcQY8Y8DRZXBi87G0+AoQiTP1zBmYVLZ80mJ0+ZiTpR
Qem3cPD74VDhm3Dxr1nXL6GD7/xAthxX7XkEw49INM962lsi/axiA2KubyXOPDaR
cAbNei5NqOhQCUZ8KDRFgZ07ItnZJyoif/TJi5HNmqSH3epotpfEqYzmrf+RN3pF
Az5hyuVN0mlRzzrhkUuDVt23pdELmSdcf4RF9XP1AiYyxdoc9BeSnNVR5UN3YJ12
HEyLuaTomQNhsV0AMCJ9gGS3/77449f8SILPWuowPhF1pvAfUXh5MNbv0tDxlOV3
RVb2fGEOwWTbObPjIjahvAeuVz1Wp/Rac8bF2sdkW1LUeSoGjP3iRPxNvYvvyrJH
1WoiUYJLUvpwhWzUjxvU018chf1Vm9ELI10E2C79/xJMafhyFI8EN4C7ymW5gwlw
if0IdvtYIKVBLlAuIBDmY9Vp36JC0Ri/05c8i2rCTlp8F8Lz+rCa8BL1FROQHX5o
vrxc41reVgSpZBtqkgGNy8tUoVRpBhuKy+L38nrpeKEhXWr9pGPC5sIvcjswWypx
KMVQ1oZ6upvuUqdMy4+JQ0Bpi9rDi0WlUBU+MQzaG4R/vMr+bpgURhQDr75OMQqn
uM96lEntGTWFfYQ4KGD9bPmhD/X65NGEnL76VBQMiC6/1mwHn9B2OkUpMhtpRuIe
C6RBUSZ3IQcmM4bXHhIOj7Ax8xq0BDLWPo8tYJNRAxdobploDaYlup0+vl2lAX63
B9DNze9PCc4qKEE3c7RJKm3SkJVCqve4U/OlOXMKFRAsJP1oOWVK3KknFEopMRlB
H7R7aFNBuYBpxdGzIRmrSxnEjAgfS7RA3v66uCj1kAemBt9J4qPcCPoKu+gPN0iZ
idQKc1ebaBqVw/Yfn5/PVTHSWrG2RjKkLYNAnUTLQ4SMJOoy7ab03+LGHGt1F0Dj
MYdq0gP4XJL9swnXAlidwz6XjmkxrlIKcMxCoyq9NnoIrKWsNY+vzGwyEaQWYmh0
LpDgMV5nD7pjZXd8oCFxCtnGsO3fkQrUV4DEnONKXV0bRIVTQ2mVVPjN6X0TvESP
DRMd/a7WDyzMFkjWUeV7lTtJQKdgNIwajqZFxU7R0QF5SKybyVo7c0NyFL+Kg05K
4YtGu9PH/yc1U+EcVDQgOWjeRGSky+OEdLluqf7f/d1nRZGhwnQKcbWM52q6sDaM
ab4xoVIsBkmQymah7GoTFd/Ha2x3udnhWpES47ixtlrh972nSupCj0/sp2r3ZZJO
P1mvhQZ1DxkBHhNx9l1YUh/gA7pDThKQuwEAwADhkcwFTOAPyOpdfmQHk4d10nhM
qJn9oAEAaaAkJnFkSKv7sAKw70fxPf3M+wW5cphPeu3jIECcvtq1S9bccBX6T+EV
LK7F9g3pEXJdNV8qEJbBM3oV5Sch8GBIWBfGk8fkJyx5wW2yiUyXTHCXjyvGndu6
ONMRunK2AFhV4rJbdf3inca7UvYISV4gUiTeytOppxSNXLTCXXrIA1LqLRw5AP0M
9ceRPc3skRA3JbFfJ24uvvRgka9CsfGr453/GsgwHfeTDz6Ac9p6CLSruSQhuUYh
C87RDpq/21b71ygULboB313XvTG999UhCGZISMp/SP8qVhM6dzWcwdXvclK1venr
SGG+wpugzyWumVw4ZMKKSdmL++9zIl1bMhY34bWEutmhtG1ODkBW8OE0n/63YIs2
AFkEVNsW1mE7vj7U3papYbcFiTuUUDYvzSHdZQf6U/9Z2MzQr+wB3GvV2zTMd/Pt
Od3teumMpw/By5uynoYUtJGjNSoMjy/SBsxNV6ELtPysu6BzcBppMJ81ESgNcPyj
A3py50jF85ggOJ7hfk6PcduscMibw0BE63c6xIuR9PqZwtYCy8+GgQMRVnAakE49
rPbFby0I3L720iKaLu1QmmuO9vVSxrMDnulYG7X8rY7vkwfWo76qzBCAk8manQd+
4CKBhEzpKpOG6VCoqrPk+aumATd9EUzR9I71/TO4mMrz/UeemmtRs/6T16rItYw9
j+CxEvzsmUabpS5Zsua07XU+YO7fkfHr0vEpvPF5/N2hX0RJHUa/4EwVn+UL2dNd
wVFRLGNsv20GfSoOFIW3hkvjvbFCt2psj6RZFITTZFJtOMeHG4Q3BVnZbDqJkzgd
N00JWCGj4ou+H1+K7aAE8MjWDguYfcSpzkvIO/sAEp9DzTskwWX+gzTDKQcOgxlt
PzaBsta5+9c4Ify4keWD1giWT/oJEgZAvbFG4okLt6AE8Ugzuzlt1bYlosD8C4LU
i7MHkugyfr5uwsEbtYFliHpdVfNohNoV0OzNyaRrhvPd8Xh6jNbvOKUWlNNGDmvn
t6C+yB8VVmfnJlpXU9lO/wSLkFVTFZ+V8gQwlD+0i7w+PrRH1ulakz90u6AbxszI
hIUXTlderg8x1DNNtZr+1O69tJgTR827jTB0NrCyXkYNo766x+GGnMK/E+Jo96C1
NB52/blQHpPVCvSdJjmhBp05C4fqcO8p+vB76GrpzMEDTkZE3tS+OGUX9OOzwly+
yYw094Ka52iaKzToUi7ZLkT2W9xxJnqRvMzQyYyaNkj0+poxUpBngzI8FQ/Vu8tY
jF5t4CnKR0Vo5vmwjGxEtKDbhGyU1/irpuJovtGXJFynSXwmk8TRT1F9TiK25rfx
9aFeXOyMXGk55DnEk+oK+dkCI/rzKvSEbTfIeQCDWib4gofLMYnFOOFGxE4/MFXp
r7l5JtGy/Tyl49gkmy6vHbtNMTIk77usaszTDydntnDvVa6GJBx9SdY+AZR+e7Zw
9Q/Yk461RFDELzGKXABSOy52DlZJ5mMp+Pev5HYIfoVJeJJYWtoIbIw5fR3QmPxL
jBf7ur0XQIXY3FeyYqbH1Yvx0eFGxfqL0TDuX79oHPSSuu6z+NLLbFbMWfcUzcYu
57GveumX257AR+heJi7Q+pUPrlgH+yKylhbcYHXk6FRPVIQuUmnpJgzYCAZjtlAD
iC10NACduDn8PV9ZW9qUsHrzqzPyyQ/yQVSjU4t5ylc3xm+9HxVh2MjFmNm+uf1R
yUrK+NP/akVcNTWur7ANpiX5TbCFxA1tGPLylSRA+EYYpew6zSS3crMuzlwaiUIg
C9sh42AGP1f0BXH2b5vg1oOkZaEARpFgXV56yKgqJplmv4N7hCmgOxo4wiWz5vFb
IvZaEhSt2Gd/JDnu4SJb9pl1+2tjXXz7UqolkXGK+vHBoqrt69MNpSyu3X6aPhuf
7ukQKjX7ff34HGTQo+fmzion03l+UOhWW0Vzor2GowtLYcPgofFCHxFY2LEhKqsU
6H14vxBWn3VS5bpWsm6yAmqCPGbN+uIOj06zYfxAi2MyD6a2ejEmLHSEgVWIy6UQ
qxnR5mb9JpLeWTVv/36ni+ghflUjHHk0VtOiVDBQMVz+HrTiKE+pjDZfJ7KnFWZq
JUgCFucbdcaodcpn6gskNBYi7xprovrB2gGqXBKPfQb711qI625uuzNKhiNd8TT4
2eMMqK8BzHkPXKAurCbofhgGC+/E4ODRhIrOIFdlpjoYYinO3LvQ6G1Y2p8trP5k
AeeMOU9CxpML/FBkJQfOzhH5ytqVXt0/xeXGL3I+Hqyk5R7Rsy6nkpWGwFZ6hb4F
EzOMVLkuZOh5E1JvSn4TQAsiq1L9iHpQ4OZ4Oiu4jYS7KlR1YevuKG/sS7315kdo
quxC+oIaz7QWQSrPzGm8QMqWJ0k65eC4dZD849OWuztgdYUWEgLut2IK+qZ7EMmk
E0zELHtOFqkQBGnm15LJ/W4LNUFgfiXoNTkVWPVJTsZp8wJ31EGRCM1KPxEt60xK
peVYP1NEV8v4Pw6jTYk/Ob8ur+QkJFQVVgW14mScG960zMS/ZaeynEvGWrP7wcqo
wuKiUDd8Zou8ASB9MeBVOgr0gAzlDTxbiGwWIx2N3aWSFmFVdBV/qb+L6dsjL+3v
gnGosAJKbCeA/OByIW9AZvTUVCRIsEGqIPzoIivwdFguXnyqla2qqS7s74u6igOp
Gk/41rBQPO9Dt6ytcEiBJdX/MyUt9HLr4rhRwpZFc5+GLebcN5Geg8PM7BBEvUPO
CcxFf1HhuiI1eowXXSofs1m8BxA6II+3yVV3XcteMFK2syWtPhW3nzK1wna308Df
wTIJwNRRKmVf7bPE8Hoh6IwgnCq+LkO0IbU+GeR2GCpewT7Sg/SFfGryVdLORxR2
dFvwpH5iEYfYT7beSsfKGQm7JB0g/eD36rHA6QRcyexrHjQcsqMtVyhcNmAunFo9
UckcPSDIBVX5XPd6dE5oJIHw2EmcQuVhVXhI/orv5XlMOTHfpK67ZA9puP9C9iYE
/V2cyRjoNanIBOyAknyWWaEB9wazzls5ah5RDurGiLH9ZtebMOiaFNZrCnBW23yh
TxLuqJRTPwl2VqwXjRRqAZOVuN0MfnLkySQtkp9Gc3XV7jsNky8a4GB1x50zaGie
n65XeT2J9jTMOXfX5etJMrmfpU/7TEWVloMy32i2RDdKcLQ/Abt/EOJy/2jwG582
7ahz1kKHdruqnUhrx7p+Pfgmwe/N0bkmlsADsRmmQX8dXeSeIC6KsHX6GATiLBFG
LUEZLuXZmm+ubwPuYnByKr5Z9ZhxRwAB3nBXcihYM+kkOWOi1nVJ2EXa7w+3W4eM
bDZcseduVanvBi41f2gc8utU+DyFk6ndzusMwiuJGtEm7GtgHfDc/w41iwT+KtvY
2iM5e0zAj55KDTcdfgIg9OwXwGJ4NshGNwaca7KN7OsEeMSdhYi8zJKiZllovFXy
NFqU1kq1I/UBam7JLWxd6bNqWyMFUBtmi87f8arIT99YrQLIeXTWPeu4IhRVxQZE
VM1j9CFvPACCG7MOIbIvboOGJq+U6NnyCkv6e1nu+AM6H41bItAweZINhkxnjFov
VVuHLKtMwdTSqURDLXk+BrUUSQUBwznD9xZpvb3Te1pXUJcvn30QbNo5LIJRihS5
1BVll7kyHcSoplBLaySSrZ+MZ5Wj1CVf2/qNIhnh2DW9gDz1U6HyDUDxNGaZsAjB
2m6chQw918mLeW5p7gOB+l69n0fRcCXXYRidrZS/zdn7DGA/jxTCHIS89jgDZfJ9
dbf6Uoy9t+lm9NAt+CQ2QOiTCsgBAm0lcCfxTEzf1wfFxUMAOFmCOTgkpD7MW2FJ
46u+phwQvJFicPP1fOJd5rkSXPR4XnTPcjNP2H1xqxMhhondWosXOpvCICaf7w8o
IB5hBFSaCBBXyM+550VYV1G7BLvtsqOXRwME7A2wtli5NaBM8nc5L71N7TW3XrRU
sWwjHdIsvi0EMY+En1AfWLpoG7726NFLe8RpgtSVPOUWWP/NQs92E22pe3trHAKA
KEQD/zt3vDOSojItGO27ZYiA6ULiW7Zs+hDB97HCmoYy2DfSOyvQ/+b1CzGzLTpI
htjQAzWSthy5/56zXZ57lwNsP1IYxAOmDH5bDdb7szP+14GIBuccykyxOihn6uH6
PxY4ZnMYH7Y4rYMDZtuAfDvzF9EgygMcB9H1W28nKeols14s93B9HaJGPeBLMDF9
E7911Li5PIciqyZEUekFG+H61IurGyJq6KA2iKDikcmSm0mhiu51kll81GxLQ9v/
kNS87xpRPMde/TRgtb71//Bb2CrOcxr1N5tJczAQoQdryB5ErNcNTA5sqRLp8/tP
0X0hDi/sW4/cYkZPaJC1CxiQkhgACEvQgeO2IJCPYv1T/aT1ainswj0L1uJsv/Uv
yB4xmY4bbU2fPV4YbKKw+66X5Q/0UrfMudi41L5i4cnK0nnldHtwd+08VF0FgrYF
5gLWvILMJRAawfjTLrGUZz8eXxukha55SP0OvKU4ph6nQx0+y6KC286//7iZR6lt
PSs3jbnQYsI0DIuUn+tv9HaP0iBPvvBlAdduKEaQrudqnpT1ecaeGykyyNkV9YFB
5UFsAQqHMnx5iKinvg+rQ9S52rulP26AXwUvCkcHJAawqHTPcwOxGACYn2GNFdkE
DZHidm3MXVnV4ULXbAaPyyJPVYN7xpMPxVtNTuSM+C04P8EVyYzEBJ7XEtH118jy
jq5BP8UMPEnhd429vatoqqv1+rZTx0obQs2wVqXnm9yxpPPCg4mLXLWGRb+IFBFZ
oIK6KzkSM8KdINLJUhpWitSQsxClqu6MbA/hZzsgzbFGDJT6RlvpYJV/XVSKc9A7
3O43+WvZdq/+MdLyQtOQc/HOW/cE2ZxtHFa8ZIQshrsLdRdflt1B/yzrNL/2ezvX
OjJX63ryZJ4sZyS9K1xYv5LQfbR3R9MlxrAJyM28/dgSRcL1f3iyUpQK2ay6nEQL
+tWko3M2w3p02e5GSXA4qqKop2A6VqN8Whvws8QobCepieE52VotDOWxGzGQNdOF
F5S2/fp1mKkStb1GjgfCp7ZIWKhvIovLllzEXDIvz7QZdDst6WxKlzXc60vWnYh/
R6CIzzL74uqQK90ygCmce+sBDJdTIs4+pProipnydWYIhxTt1lhN/RyYdOziJ+/z
Dhi1Of/RoLhEuxEAo+t9KxWTgabdvHHQAa1uTA1sF2n64fWwzBZzy3jJQ+DXxbp5
IHHuT3Y7rUTDauPx3UxNb4If49LCThgfft2kKbmCfB+zVIWSi7XFvId7Om8h81if
HcHRD4WMlx3nlOo9u6sZSTKkYM1uMpy9/9TMmpYZRWCF4Iyh1eDpgxB9en5kaNSG
mIFEFhLvkQ/RkubeLqD5IjTR8akk/kO7vLsucvqWR/JBUcK9Vqw0/P6rFDu/oFnW
0URItl4WLNPMqtOWKYExnjnAYJyKJOorIu/eD80uhG7NUDSdgALuMEDJ6rX37zAo
OR9AHi8OU+e0pKoIsAJVy1aLFJG2VNtyWhQ5FU/2dCFTOUA+/xLbbS6voonMtGIT
PoB+HmPh1/RKW1rJcPXgXQz+PnPaL9BtgFI5Tlabi+1zXKeaym/q8+ir+eZnhjWx
K45GmFgCFSMmop3A13g3ec30ETu4pocXjgfHF1oKAX0yqixF9Xd8TpiWgQxKOsCT
RvkV2+4ZIXuXebMF4J20k/WBZcyha6ULxUalBrsZLKhCL+MelQeObXnon93v+d4y
JsWMwTlsRZ4RobdDkiXfurvqy+edBns1Qj/GJK+d3r3MgLoUZN+q1GHuL7G5SnYl
OBf6hrdyAv/L5TJfCLJOUGhkDXA57/dA+e4LV5eAIwpW0OSzkOUxPkDaY+uKn2Hz
SSpvbk8JOmTu72WFBVVE9EDOFHrj5dAe8KhIQHoOMKw30OllysVD5NDYq3CWHKBY
wR+W7CqYVNvOa6nkecOoSFCeZQSaSZAEucHKQvacxs/75FLMtmVZEc2Te9FKMK7/
Y/WSiUYwXAg+miBOBcI2FJApTMFyIpjd5MYkFoGKMV46anjuf5hq7XZHaU2Ionpt
HrptQLk/eYruM+CX26AHJLLpHxkp6Puy3Xig3NPpu0Tul4gvk87+0ocE2lJKZt4B
W1M/0kBd5Vorcg33yQJEZJpnrNhr0GEZDGQYvDY9H06gTpi8z2O2PSzf+ySgjbh4
n9TOJ+axakAeHIqV5z5/P2yOvaudXGzZl6KZIT/aJ4dZJaUm8UlDgQJ0L5Ythfi/
MoM1aW+WpMF7JBZQNRA6eS5Kt558cmrSDPj92BsT11hEyH8JlqeGPQigO5KAj2CP
xxPMYYQRbFowqJ+iG2r4Mk9HmESvAdropLNCyc2BC9UAogDPzH9/OYVhS3fKwIvU
Nd2SwwpoWe0b2qIO+I7Kzq7v+nvh0m/85yfps/HSACMmSv2WaNZuzMn+pkMXgACP
O49sUTBPiD2OsZjKxfG4dCqaY1v+oW+M+XqO03MJ6Oa3HgFJrYrfJBH917Joco2C
tN8umO3flMjEBlvPTYdmxL/F/UBeS+aIn+g8OZ7D8uaZ8vrF/muf96T112N57Ve2
rDhGcGa5Xn+OybL+i/nttLPLzwTBr49InMo3tihaad16xnG4R49p00lvykLtxHRR
F2A1hV632oen4Sh16He2HtnQOcNOOwWip5BJ1TPBUZzgS1iv8Oqeyh+FjpYP4UU6
GB+SIMDrT34z5vN+oqV86a3nebGJuwszYJuCAJng3EmtJ2lFAtomyIyIRsRpgaNd
efrE/63vJ6AmKcXHPGzHvwDGNJE/ynDfVEu/YAFrv2x/Jqzk7hx1Ysz4P/Qw+HTY
7TkQOS5C5aEOtW/zR6hNza0lhIFRvV9zTJB+4CsEXCef1PY/y4cppmvjDUt9Zz7S
3ySSAc/y9eKoKAUGniIJsSkEpABnNrOhc5G2rEC6xAWCYq0N9ovyLIZswaQ9c0Uh
4Q96LGP+HSW3cZMhJxn5fvIr3JI3arta6IqiP8u7Qp41pYZAWHj7UoBfkAoHy8fh
poDL7nZFOrNHvhYHRQtXBV/wwdMNCPAbYnXKMlCKPXOkpzZ9n01WKiB6Ti+ryDMD
9J4QbckxDlh0SYa4NOOsbhgr0ojxMQHwf7w29WOzQ4KL2t4OR/LcNYm3qdvwkTm+
gdu7Eqihax6Q0N/GJOBlC8rvRsz5ZJB4EtD6dpDAb0Ck1yRCWG3NQ9u+RCCsfmpo
lg//oXwoNeRxfqrI5ECIgU22aulA/cPotoy9ndr4SKip3U/jDawNKoloiFiWhy9t
VNY8SX2IM2K/DNdGoqS5SZmMq20f845qBxqDpL17jPiCFEF6CA55xvukN7JNp/2m
4PO48JprVwlwv1riogsUY/qO00TLebj9HdqJtb9BDtCNTvTRAC1GHkoAxi/3z22J
QfZgeWsI+n2vezyun6x/cEWmEVBD7tI058oaFdrMHrOqojknxONCL7fEpDwDd8C2
6WzzqWecCDmxxMRLvnrvD14aqxhbD8TC9a5TVztqFeNf4MKMZHdiKDbedjGn7JMc
3pQIfQRly+8Dxre9lh8a7u6V/zkUvEid4fQmi6zfRKHdyBqVEXK8cRdfrIsn3GSx
O5IBhVBfUR/xtL7N3YgPlQXVkJ+/7muCYRHWPj7Bu+9/oM8vlm0vW15gzbzrMiHw
SmilTMcDVq/OlhcDuoH2O7eqmweyXtMsD6lnj759Zv052NnoscaLPKPYA40Ei2IM
Aq+HUIZnVHvRLAxvJ2NsXh0QQUUvoDTdo8oeNHB6s86sddffIaT3W3qK0RqmKKnJ
lB/dsX8/pVUmLS6n+FctmTj1kl00wL3QlXimhNreGUoWJ519A2fmVd0rbcwtpTvr
yyHvixRIhuoA/nto4VEHFMwg6aQhSOr8YX6FQGyQer7x2Kt6mkC7nEASr/kmcBKG
tjQpAulSyf5eLFLJUK7Q9Z4I53iLKfRhuId1bbxayJH7e0VMhIB11qHOsaqXeTqh
A2vWi8TKn4YM9WiEL5mlmYwmQZNzXyldrZ3mgb5Rt+30adcbHa1dtY0wpvX+2OlL
ohPGazIRJrDmaW5yxME3HGJnd57FWkE3FgHuUk+ESdvO8dUpg4ZL7fNVyv+pYHoY
UTxzO7ZDF8XQgpQkRSl1TOZJYshDQDEEbFwE+mJ3saFIxkcWvD1o82xzrOJo9Zfc
MezA4GPBdlFEJBOf/eKeLj2b9Ss0zCXJKx8VPtGJYQH0BtH1n77OF71aBLsgGPYW
w6K5kJs6x23dtYayA0VZzAZ8grOYTsfBGR5GAKHmp5yqk+7XMVyk4nZPt4x3ap4z
UgKX/Bd7RWAWEm4Y0FJ+ufl889NipQK1kMpDsG8Xnji6zdXFODtXpGbuT1MtRSTq
b7pRWP4ubVOcK2Z6Z3HaCEnXbcyXNopwYVM/DpPVEUTM49HQupTb7j6CqUR0xShm
dBoqeW9BT66UfppujSWnkvzbVjMisbWZHWe2efcPeZGEpMjmFG1xNrtubHmnuJYA
jA/wsqo9KY7u2GBBBhUaw01suWZOLbmQp4+gUHgAcfeCbL897HcIAN6gPBc8ssr8
IQosc9I5N5An5CDPQg0ObFObBS5Pm50R2nbbZsMfFAVfye9mI7k92qHYa4mepcu0
5X1K68k4yG0yEsoOteEFJajfoiHc8+kwvPTgxgneoQTZLIcYzr7TtJ4+ndYs62qv
NtJmIC2WsoiqFRshVMaOUodJ2qyfTWx0xNEIhSvarbUqJgw5FEJ75glDE3leibpo
FlSocJCTJ/j1LdDJRy8NnNqZIyrRKl+UAyd8rbcj2rf3RpnannqNGD/h5T3AmLLe
1PQV/2YzBbyiO8jvuLENRaKVfYpYWu0HpKF9wevb4S93SzVHY4oUTvEDUdSeWm5r
c0UgKVU9VySYBR9BsxyNlOZZNQ33M4kGSRslkIFcMKhQVrDxTqe3p9P/ciK2Yb7C
2iMsZ+LbuUfJgxKrl55EuGsp37gn66eDKWzA5mcYmtX9Gt5ABy4X57iGc50SJMoc
qL4caufWDSX6gI3u7VtUlhzAdXRQeB0BPmLBC1vkYgLc1Z7TVeTkdWYFqKTUbNxa
jPetskaO1bCT9mIrNt3cdThWptVdMWW5YNr7hgdizNxmuq6sud+Pp8Cg+hlRVzR7
L4iyn3S/zjJwDQOoPpDWSpa8Q8Y9pQOSseV7miwJxDoWji39X2p8YVEhBxlcVvlf
e9Z1nLOORuGAEjouSHfKzTQGdpmJ7vBwPP3MuIwU0QJU+w4Rzo6a0V1Q3pzJ+SxO
zgAePY7m/0U5HEyIOLrisQ74LJXPeGhqklj16lCSE8DKd0oq9Z9JE1ktaofWkbpx
ApfgC1qfgHSVzq10N3FBZzh1IeiCho5yBxDA1+GiYCoR9qzPsaMuWNagsDX5kKKb
HA+HkDkosykq1tP60QoUaKfiQhkjPvIIu4rjfeKLMX56R4NwupUEOwXAINXGTRy7
60cHhC5MEMA3s2oxjdPd/QpTajV3/eLNF9G7i1B80bDn+BBd/6vleilMCMsJeGDx
F4w5UPMZxXziluwfJ+5hR5pxtOhuDj/sT290xY72bV2GGz1R+b8CIbtZZkJQ0kxx
zCFerEeODC5LZkAyGKVzuTGTPEERNvC9Df2Pv+b4Ua8af3+M2qokZAMMDPcUdl8w
Srx/+feNr5/GkQRt28g7PLc4B7tp8/mrynV+W0aUypTFUKzojmXsof7v4Ykc8Ulv
/3P7RN57Wh3ImV6mgQXASHAG4qN3tbubVJPrC8dNHbUcCv/WwmNtxkFvFQzsUmAN
iVlQi+NsLWMRcnf1koyYg6j6r0zUTHPqfRUJs5YYi0aynXMolpMIaNh6dsI3mJzG
JzI8ndyLNvM37CYtFUMd7dkLGuUWvqhq0skDnu51ZSv4WKdl/CzRMvZBGRBuHXnf
+GSRYIaUaVTGNtRECDx80JMPs0tYynu/1amcjJDOPPxB4GeO9lOyjSmekDsmFaxM
H0guX4qMtpg49Rz/B05aq6Vib+zpOkpQ8R/KDHB86faBRaAtsiT0x+3ZmCxBnS5z
ocJl/Tnp9uvbhktk8L//6ZwffV8tHmSGk/FtgGP7Z8Q6wB+K9YXy6RjtnabywQCx
r/hg0GBTkFKK9aVzhs9hLL617mskJykevLSBFGlip5RHDp5CimqnUXOVDI+S/ydO
ZyNV2YhEW8LyGD+twMBpfP2GmFJ1w8bXXPTPJ1fhUIeaqW6/d0EwaERv47HZYxbg
dt9M0rKKdd8/KMvyyQMHoWMbNBuO18Nfp/0n1fw7Mcfor8GUOrIWz2u6j+f73SGv
/8rL/0E2U9JPWJxIXejrIIKCCpVgwyW2I1cKY00PTzGwVU1Gue73vE+jLe8gSrZ3
DdGq88d8DCSViQNiq9Gg1bjhsxlaM4SsZ7joqm5a7RBSuC+cK7sgPj2lRsmgSLA6
224FbhCtVU888rfspNAarD/bsULvpbYr16c8V0egJoQdzhkJSF7tgbDeXYLUGTC8
KRtqx1gXplXHU+X2skirghX+6Wva23Fcg8inMi9IE+9w9Kz42mK2rqBXcKvDC4Re
jINkDkGF+gqIvh1lr3QzFi1SuPMMGMV8cQaUZ4eeJ/uWN0GjhAw8rm77WR/HQxHn
viBKZ50RImKwzn4X55q/D9SWGlMKO1CAciJRwVSOYkTChhwHAYIF0wAWke/etU6b
1yEA21mPPKKtVOCmvHnwzwgRzhJ7n66LLAkEN1C5ir5CJJ2mch0EMi8xP1F6AM6e
7opW4mlUkYV9Cl6ArGJyA/psvYgcgNS2Xi9pAUXqxtoxxUTHwwoxgfjNH79+beeP
3XZcYFrX2IGB6Ucuj3pkoZSwF96qF8RUm0af0yEbs+oXhAQxt9bcz95piiNLPp/I
6DRU70Uebru+dhDvKiIwl4Yj6cfAXbx4lgYRLvwZVC/0HKRYtVqzsQYldz3BlcFl
6VMyD1DOcvaC2OrSlSXUFJdor/plO0fkIfI88zKwOX3PFM9KFuRBwpMfQ+UoARoP
7vUsJOK9rpyQh+G7pILudW2vdX/ccOe4VxO8qIdVnggIkFdrTfLrz/53UmLCp4XJ
sJmd2y7ZphLM1F8SL4spxeuqAxT+LPX15Nhdbrwkax/DIP+TlG7Gr5RhXrBpatGG
2SAihjkpADuDIC/36elN5dbpGfqucijVZH+FGoqZTip2PYOkFofLNuh7WNAQU5rg
+h/A3O/RbGKc/5BbcGc1CsUe0ovwLSyD0sahYSk9se3rPyzPCN+L0UrBHn/C2npD
lfuwwpwXl5BMfblvbSc7IEXH4WZldClOfCHFCoXS0pj2MDa81FpEM5GcUHQ2VgH4
q0jIv2CgxYMvg49TA66tU3RVAJb+/cK+4ooOd+/XMlYFaunVSYNnKaNsvNICH2Ws
J/AaxBGBpbhIaHPrB4Qdsu93/XFVNRz2HTzUVielAD1yhwyIBCex2xw3oQZG6dhi
vNzStC6nydMiuNejjCdr5MLPYlFjWB2DYvvUOUu3iTIxjRbHmVzatNZkX+xN7+YW
t6uEXyUjJyZIkMM4Hzm7g0K9PhA4RE0yHQDVBe0yzr+VVJ/z72PbXF0eK2edPY3t
YW1MHpombpKc8lmJTSVStWmx72ILf/aoNhqcdOIyYqr0guauCvuOjzGQkPqGxfwk
6xst0ntjzP/1nGB2kID32bu9t6CdyyVVs2tBJTqDag6UQScfr/pdP/d234lYVR8D
wJttv4EW8W6HazECv5wWUhQx4RoRYKosKCGA744wspEGbYDSdCyhnrvNUufm3K9z
rWhwz2QGT1v7d4yngUKIh1qMN8+ITaw6wETe+3M2/ttvv39QIORn/EwjQmtQ9+FO
cnOcbNcv9BBFP0io/5/TeQaXtwYeNbwEDtgOzyNGtjKl8AHxTvWI86mfQWlh8+Eu
qKGTz6FtrWMQO04JeekNlE0Qz556fv3nKwXqFSdj+7wwOK3/OmjAtT5xsIQhFXO9
kygVlkilz/wrRAK7LhVMUfggDPdBaMg7zU7hBBoJRUtzfSdKeAedpfNlWzXOm63c
teh/8RiYu2ibsZaAogyygTb4R9zr3iDDa/kwQfA88m8BsBO9JndHQPzPtsMQdqFd
xFuAcG4b55WlXsNu4BpSK/pdATYi96E+hbpQjRmB0Dgc9gP1X0DlSb/bm3j1rAJp
mzD4mQOL/J8BOzS/BVzJJZXd7TsSbpz/7HoJLKPZYaMoem8NwmhDycX7MbIZmpmL
x3SIx2FgB7RFqvTHXWmUhbVSDmDUe4YcD2ZTdjWOrCUhzoE+8AFAvp+cCF6y/zg9
ew9VWyih69jcDKUdFCNHKNZJTdBO4SPDRvvyPq7xL01oTl0KUXevYPZ25+FL30D+
TCc/1WffzP9cuoUPPvCJLbWfl+s1NICGaPjWiie2j5kZt/S4TPoVQzyrsVssSCH3
zhqI5EUHrktgiz3Vm1Cf3MNNVJv5vgHOlbf3VEXxYRqOmJj8rzj1zEzgybPOCeZ6
FSSLhIJXFvnhwu25PMB0NBnserLPEWXzN84sQCq4YdNH2Ddn+dparjTE6co459r7
8qytGy5kiSADbk7WS35zOw8HiENf3X/kacoBNX7f07DtZsid8ukU0lxRHsZLmD5F
W9Ns/YsCX7l619+p4fYS/KUiVLjElyRXQnG1Ns23b1YGGALVLD7nwf8BkaFpjZhR
XM0PHIAnnXEbguaHbD2dLmg8cPx6CL5AuOfhcCPGTcUqI8auC6iXKOpzrUltHFun
YFJsHh1EmE04Jx0nB+4JnwMd29w2hKMBfkA9mpwXTwsrhDb277p/YN3HJ7IfXaQO
qgUHvXUdw+Nt8pZ3/mCRyAlG0O15lrCUZkdi++dNkRqB4eM6I43qEnoSyeZ+cZgA
YY0JOmcmLH30KiwqJyJT14anR3g63RM4YZUw+hHoWyreVqWW/LRaepaD3hbgLJ/C
7740hrtZ+YVsX/o731UULP4SjQoVn5R+iW0jQdIwH5dDLpkEPk/cDPdyzNzH0Rss
2koYIDCGgzUXcdrJCCeViKdHpDbN5proaojALHYna04+qMSeDlB26Ti77ZZtOSiR
TBu/5Gu3pqBvDoeQA4dx09S6oyE5VJC1/GtBsHGQmf1L/MhwukR+3X3N8e1WbNCv
iCHXo1L9dhLfSMvFsJMt/0XmR7Q7uQKlkaiE8xS/kD8hy2FPQEHG8Zh9HoxIDJPh
OCoowxjR5jopSCSrouLRRyDspxzBg9Y36muVXX0vS7POaucDzy/M1bX5dWhK/qF2
akxYvTqlCMJ9HTLYkb9UtONMsZFyfnHqQCfJk5FuFKR3/97m0oKyuLRrbvfR1o6j
v73bGYOfQKm3+IiMYAMcwT4aTOl09nTzJt2HkYY2H5TCpL5xDYnlCJvNMVnqbYFC
YW0vk0pPvWpvTqSIcDnrl936OLQ1sqs8Ktj6YZXlHnZGwWUUyokJFE0GRixu81Be
ManB8abRcHfMmPdgw9ASwwaGzoeJiSSb1yDS8fXMVwxJ33XkVHsO0T5LDgjUiVmN
lDJcHrSYMm0BKfJNz6xekXLulFt3nhh6/ma1p98NQsxgaqMo3+vnrs4V5GjK5hqW
F3R4TtB3pSeduZVVRKb6hWquPI6GHW5H+8/cKSBDhKBEus/A0rUnAPPXx+zdPi7h
wwE674MP7M4fZqX7TkbJuQnf7R/zX31MXzvOGYqaU41bjrd8ikz3KrJ1x/wTWpZF
+z5v7FPbo7xqukF2uTjmOZOAcAxtMHvXq9VWkfpIJCubjp0J0NzsUS98fmgITLe4
gXVRxMn9tgn0WSpIEuR1ck3RfFzPtkwlHy7BUKG9s0aJTIMGMCD7IfBxeveYc/PX
N8EzrZO7l3qmH3fvq9BjEFCbEWY6xVcLJeXN9hFclU9emTYE/2rnPqsZtn/IEbMb
T9DyZ+TKjKFOD4z6iU7w5e8sj9lGhX/Ki/kJ1Ev3X6CTTWTR9t6WJ4Kf/1VNpV0X
KvLg/wyp1eUb+MYngfO9Hy7DmxUeuggP39EqKIo2JE1S2+JVp1n7YrkmErl/VJaQ
HutOUn3LRg9T265B+xyguPNlRFdGfWYlebFbYovAPZZF6o1FXH1O+V6+MlSZ6zJ4
UaWoDdGftq8PF5aVqTl5xh+Xlvzr70jV0pMP8SIZn+D3OqE5th3MlJWj0C0sCmMZ
Uj0ULigPXpd2+20SM+UAR6tbPKlYDpmEOxU0+ES3alac/T3YG6WT5h3v7msDmkrl
oVPFU+q74Y3gqcFANd5KnA2L0a6he3Q0rBwW44yYfHzPHFVwMiIPc0g6IU3fJ3pb
YXKsntQUw9uvSd/atWN/PEmsCl7ZrdbCDeJJdSjNGQtXbZi9rL4Kt90s9ZcwwXja
GeTnbz6B2hwKb6+4RGHUiUbSQ2UxPTrjXFpjsWG6bQhTLNPvlIPS1DtW57rtjCpi
uYQdpI002evOKXZvKnGV9HV9D3dcheDEtQcvfWDgR/QQ92+3kEh4jMXn2IrsC3U1
TihhWb7n2V1Hj+KnUYbOVdLL8r7mHXy+hWsQBcREyRyfhespFGIeb+Sudr3dYJoj
3Ucm0FFDBvf91ewYtgyyJYU18Yxn0nZywSAKWfP+d8gmvIshnCz6m36LGzEpWQ+a
f8LnuoaS2oGiiKYoEm6zlJjQuGPANStVHo/MYJgwv7SnOgueU0w8d3ljAqzcpmE6
tzrJ7594bGtt/i0I2EHjPSCThvC87N60myTfUvs1rglhYCTdp/keEVCTPWVJgK5t
1jSUVBUbpL7blfMCNH0JoXTQ438sNBYOl9mEHeMmGq9juU3TKIPzrtDz4ug3WLru
OmtZGswi0cXgmI96ysJ6yKOvNkVF6SGLiLQHbpV1aQnFl2fF/ScC//Dk8lEq88uH
8t19odwvpb0gxQHsw8Q/5JJXgA31QdxC+pWA/zSe7CsczKvJR0cSwwjTAUYBsAUd
NstiYPwBvCMrPzLyLld1dcq0LHJXDC7n3gmw8INz/LViMSu4qFy3lxipAqfaxzA4
Ju8hxD5tNuZRjIIFyQv+gYGOvVaglKRsuRbSWKNQQt0The4KpQf5Owt8KoCQm62h
pfCP/hMnBjiApk2o5aaeIswJIphbmgrcaT1IYdmMyW5MT6xcMVsYDGezFPYF83MY
LMJwSaMvUF+T5yj108DKZjm4EhBK31RYtF+/ld59/kk70sPa/9cpR9SaNG6YVpgK
nfWpuY+QWJCwKs3bXvGAhjYzbaph4b+Lp2KEHQSKDoNMA82j48027lGpbUn/VWng
SulgUyYmYo/b8IGVhtofas5A77BGJ33fbfVoPc38+YcCnDLr2MbiwNYl201vsC4e
s+9kxQZ9I5Y/p1B9MzlIoUrrr3QaTezxOPKGcn9vncPbjCvDKnaZjmsjHJTct3dv
oQGMb2hopLKfaByaFxwjOaSf+pYFwIg+B3zu+Y5arDc/bVve0+ye9GOlHUg+UZsf
5rmUNCTdxFeJwr608YRs7AlBkQ0oIuokirj0SaoTYB8k6/Zaj9fgsm+a57NYUBjj
zc1WfRuSr3+94qvRXN2tVQ4aH/WH+EqeOOCwA4yfi24TBdVHaPeQf/4WLN6zhqZg
ls/FpWdLOHLptmyA3j6sF9E3GG6qM/NyRd45/jpdAvCru20bZR0wgF3EIWorLSPi
eb1A327y5B/XjbtATlQd1WIBjJqLgDj1E5GQIZbyof9RqqwlIPPopZ3dTzXt+aqh
RhG3hOKHgNdmJz7ZDuDmhlHZzbWQM1fCwmNaE6dEOUhOqN2tkL5O2XMkXwOz8kw1
VYCtyQz3Ft95LQ/WFmjJ6mYNqD5khG75jnJwtrkKqltkcCgfsv1XSXKPQIBNxDek
C5SnCnZ3jUWRQJxKXQuT0WcRI4G98SP5/7OKoMNTASE1TzGA1DYzSg/PyMXYYo0O
rkNqa7xeOj3NnNgtStObCpkQqTIiEJfdkQQ//wdXCdnuAHnWl7vH8JFZFfDHsd4t
ggv+nMc02Dn6FW/XqaCwVl0vu94qgnV9LbH0xvOb+jINrvufemqIiAWxWrbcq7x6
y1jTMimYNxy2Q7sWxva5HKh2DWxMNp+2NvJPoxLragm4013rE5Z6zLOHfN+WKC52
3kPHxwNqkovprgQTnkBYZjoKvHw9/aB0i6OzdCr8LFUwWhSjIOrLPb7fcoLt16Oo
uM3dSrP4roV20vkjAGGf2aQ7ggyG1DrW1x1lCmj7BbzETLBjuSuscip41wi06T/f
bMk8pLj5yxSii3Tp+MyoJWDx+wdEaCX9gaGSe816HiYjwhMv+ThKTQbWbE+mtiGg
xBH77hsq4qPgju1220cO36GucOw+CXQYBEnOb0Ifj3MLQiGLEU2gfwdT7cPlPdXy
rdU0DpslwP7pzmqq6mALFIxBXDVpu71KJU0/dJcBviS11VC5jKGWaafzpNLPEQkX
KHht5aILvsZ2xWBxqFj1sQ95S782BRZn8c7peULoMNTbLJjr+tCQgTQ9lwWnKvFe
jtj6Sa8cOA7FfDQ4IDHQKNtPx+0Cu0k0sAGCQlW8EDFDEQuJpIu9fZc6RT9XnoVc
GZCIRo65rz6LXHMRGRxGpp+S//Hupiq+EXp0ykvMfBSXWY9UPqPf6vlAPQF65dHE
HsWyaxqxM7FB7rwvzJJnhQ0VkGW189TAsdvV5KtZGR7G8tTpSHPL4hP4mYmoRpnI
CG6RzLZtKVCJ1K0qv0XjwocHmf1HjIkHDs0dj5yHNziQ26A/RxgYIZEbRp4zgS4s
o2eMFH6NFZnVTfNQmi322VyMx3b1uMjVw5YeswWBzlLjWUuzei9tZ4E5oaOZ54oG
toYT+BeJY2Pxo+1cj+c0VxRHy2ftEMDkJu6NTzFgRZP92dVjh2gRvi/n1PmnT4lS
TX1239ZLrPK2T2nBRnNTuJTXfCxo4XQLdFRh8udP8BpsMMJci+w7HssUr22C9W9p
VYoM/mUc97+oK/N7Uqe1qXqQAnGUothIGiCkIGg9Pe55lznOWfu5xxTETQGMYjHa
Wh9M6vVv6poTPyyYzRtSniSSuyKO1AVqULf2iVgdehsJG896Dvu7QTnlwQc0rmzs
Bj4TkOX8S3ZyjEccDiN33XvSYPyKaQeRTw8WEzs6kIuAToSHROuHx1rfzyOtWIJ2
ZuyTLMHJg3Jf2V5WILDKn9tbokGHO2ztJOke3N6IUrenqDTKNXdiXFmktWPpKlHe
nBs9WWD5+TMZkB34SdNqOYqmfW8xuoTnBKRQMeHPScpI95IloCz1GnBglzRFyFi5
UunuF9z/1hNTICHwTvX2c8TiCprC0mUcSimhVIjikujiJTXdfn0NBxrs5OawZHgl
VBC6g6E0uwlEmCK7qRtIODBb2h8cjir5B9IQi2d4hrAdxh0rH0+2llGrahPWuCZL
8wJ63PXA0JzB5p5sa207uWQp4wARaAVrjrlJ6QHs/ND0Dn4GjaZLrCr1n1yNMRmU
dd+C+Scf8QXj+89/TazWB+sGnG0H+hNwr5GOZ47q1zGdvokk8FXkW2mS95vMGXcl
yidBfozuC2yWY7vOyGfq2PNfUiaP7meIO+FZMZerlTTvy72Om+04/CMSIibgcUfB
KstAEIzD6pqfLviVQkUNp4I/W9yZA16bqGvVpW9ECJTpqARLCbSxphX0GEyr6YnE
y7945EmjPfixLvaOMsiLzOCxBbgEGzHlOj5S8GxtvuPYLyo6lTzsfvTBM/+y4dId
fYcPBfjcvns+S5QZKjzVJRZOaDy6jKQv6/aoPvXXGQBG3JZl2S0nyjC0nCk7xHH7
GuPUYB++NqpxPkIl++1J18VNdGdu5pJjOEHUMy2Sl7PnNFCGsWeSyy4zLQIUim5R
axm1QUhcwsHkai83/Evd3fhZWa1+smV5ytOu97f7Udxif+7Wm6pzebpxWgqabW2w
UBcLLJ2k0GvIKDCgU9EUxICW8xX0RdE7gEcRnPmsv4FULvbUbqHiAm3Ne2hB/3If
xVciZeSPXkQQflArng5MVrZayExDXRRxHJvns+EDotZmf0joSZ3Ks/3Y8+u9GsCM
R9JFKj6amhC+YETkrKZzYYBmN3TFMDjk8eSO/98+E7J+LPcl+ZZbjuQ0o9Zhin4L
SF4bEK3rjDsPXigKvrf6EFYNK7F+jxa9Ft04kTUzc75L4iGDxQOH0a5CKXmohJTX
2xxsA+SNuJ+Bc3do1ANKm7L+OvDmpXQ38Sk2nhO7i0GhfBE2NE+wG8g+ix7xGpsI
pNJ608r49/tUoIhs2SFBthl8N3fjDvtCS63S6qQyeYde2TFm+1Q3EZ5DUkTPq2H2
n5GKvgy0kP1dHo5QzEAbsfb5E6cYS82RyD2KCujGsBfzAKOK81z3QdAKGeYzDaC5
5LJeJAkuJV4e5l17+oxocuNcvwA39Lh1WxU9vUxro3VUgYC+pJkqxQWkZ8QPlrF/
/M+oH31WksROpM+2LzwCL24HmEN99alztlHwx1lgTwKEDv+56NklRXlgfid3N4DA
toiiqxv8CZE3JvP8sLxvtmfcm5GQrpR6RZX+lKQbLbpVSeDiwLQtBskrUddnDBEs
hnVv0TyIzKB5JCgiz3oyTRgzpTTqi1JmH3FUXgnLU8COlBWLGeE7JO+qpBZi43gw
V7V8c5N5/3NniLUxDk62FY89Fp2NNorb6ly50Xu7Ar+mONhdCCD7sa4EF0k/rV54
P6a2+0ajqD8p4B+CDao7bvqaquFclJrHmncQd8w97MNwL/6KMK8Clze/1CHxD4MJ
iQfHIX6EqkK5K95mrNo+uxQNUGPibU1ZfTysVqr2WzXskVtYj68goCj4TlchC0rP
avqxCbqACIOP+M2R6uNm/Lj7vQRC001BRdxkcvwZP0nEv/1XreK3ua09/6viATfM
D3bK/duIuhS7iIUDRp/4te3CHYiCguuP6aEn3PO718f7ZlRs6HYC+k/VG/E+njEz
lg0H9DSQennJ8D5nPtJsEEKwLtlnDAuUX3sHuo6Dtf0/wbRkVzFq8xwO9lxz2oL3
A3pmwBJAQe5tIQnolya8hY2PrXPwwP1ZZiq9B5TOz78oQrxCMSGhFLNpZA9UOpok
ESCQ8/zxmtTFe3c//O5hx0GVns/ubyJls8Dzcf1w4cRXDXdjRstHe5c/JxihdVmL
agP3M7sCmuLsJ2oJYlkmo635q9/c/vvR/riwMmYm7seeGE6dc5iAvFlw2Bz7TaBd
VGYjlkOIlmenO4JKf+STxiuXn+Rlnbb6stSyjQtrT8cNN1OtxR2WHkG4BnQVZFD2
hkog2A89Z0mxB6k4/HECoVrdJXVF3vJmMfysbPwyggBnvvlwcEJS2kDhjUwVxvPg
R5VCTyYhrGijv+QcugOOi2BfsCqEJavKOD1UJqaUAI/3BGpqVTn1RAFCVQnQbQBk
XDITPPF9TSf7ePHNzyFKHGF46ddAR+JFQm25AgPXz3JNlAmAMKDU64NyIQDWdc55
uXggahztygfqd+m5FMlX0qTQU2AgacT20owJMfuShLcZGvc9Y31gouv1H7XsK5Bp
1QfckVcYIfAjdY6FlOzAPZ/heGl/5neHdzQUTFvb164PEIeArcjRmFyv2HqoZoNQ
/SOSwKv0PXhp+aE38+NFEcfgu5QSfalzTesGMBa1XwZPcxTi181Y9DZAEaQhPRcq
arApOJqmvOslS8ZvTD2OWN9EEn91xVKxtnYiE1Zl9HTZyLPjqPyZRFAlfjb7RAAO
mI7XxcFGRJNooxJpdN7EHFssH6RuUlVmHao1ZpsKSp159ulYIN40Ui/ko7dG5ZRH
zKOFl3CqvjOo9dFcrtO83r0/FmLeX3CcJVTpN+J1/gTQqDlAHuOWkCQ4ARU862j8
/a5wAU8eyn/xqdImenIWjJhoUbAd2Xn0aDfSAzuBu7Oa9h8OXd/hfhm9Pi4eatwL
OCXSQQqZ198Q1Jxtq3w5U/QwHI+VD6gDx4tayvG5hi/gXFh7Yvjh1w5aXOfgGCdf
X0isOgI3oOe7a4CRUbDsOh/pAduMo8tmSJApZhP9wyrW0+BLn89f9K2RDqyCQKDR
a89JjeU+ZNGjyT6ee3sEt2ZeOFhtbsW6DMrO2zEQ08iR/WH+/7QUDVYS/fTD6rXH
LexhBmgiqpVTLdrDTARSHDem8cy7eKKcnHVAs7J1GA4pjWvExfjcw84hUblw+tRA
FY72H1jgGDB/8vJ1nvE3aHAcs4LQwO95xlsV2FEh4m2ZyO/81HcTin/ypxIOc4wo
kxqIf1S9oTDclFGqXgFxlJYK29rDIz8bGmctXcApHmmrtN62oosBG4TsU0e54Qch
MrrZ377+/xrL6HYu5yEjq5TUJtzpM2GXtaiw75F/nycCd8XC83//vzJAHvlUVM7s
37RBlnOaP4ZvJN+XcyRMXwvf01vYi8kNLZFkaglPatwW/xZUYIVFLoEpIjWLjY5m
3AgPmHNilLuO1oHwGok0TsW7H+zku0N+eW5CXH/v8xbIDAZoJSaHprePRYZo/rHH
K27QLRse0e4LYd+Ih34holTW+T2ybrGzLQakyf9D379JfAqMqxpP/cS/elbomx5M
oQ8BO2yA7R9mBeszftqMKhZF8UJ97GxFjTHjiwio9ALGUYuXGnGz1p+NpGFxJ9y/
H7NSa5+syY7zDceMOlv8bOhD99KQOWaZxkwBpqNBvEal8IoBB86JsyyfALi4bb79
FAvcPKGTPqp8htH7JQ8nnmttF6br+QpYpACEnVg1BoKE/z6LuKYUjKsMP0SZaI4T
SRyraj+uuE5MoVoeaL3t78aWdSNL3yI86hcURakTOtedGZxX7E5gHwYpdVnPjtzF
FAiHtp0lQegQpqWgxcpXE6iEJ2vQDaKYMo7h2mehQO4ablvITPOyxPa/66P/saju
pNots9FBxyI3WXAWfUXVAWbyNARP39LwGRxkgA05T+U+sVoloYJe9rOMksckPrV7
tM4KpnebmkKu1Ojx4oeaqGjGcq+C8A+NefuwBTactrepr4xnSHus9VfiLz5O9rOC
+D6yEd+TrNgugosSXSrvU7p8CSEWVlvJ1y75Pp3zL8VDwIw0ZCXtdmYETC0NxVUE
pQk+HVv8HjgVLrfhyGgc3r0pyONB+GOFmCiSYWXzDHkjTHVd3AoL1RNE7I97Tnee
qGtqVy7BAu95ikljNpIPJFbvrv1+M7DgKBz71Hsek9aSFlXXEf39UDn9W8RHLbdV
ae6prpDAbtNI9gs5pzbVs1IocvMJwiBPswpfbOk37dQ+GhH23j1pBtlEuv/QqtUL
CCDHQoNYIxjOHh4WAhFn06/3fgOcapqGoOLiRhi2QBMq3TjeHFX19iI18XttHWhu
bX/O8GKtlz+0zZGXeWamD332kIcq0lDu0kDlv3171/LbA6e5lsBV2gjS6MfZIJmt
gDqtHBIQctxZBf/Vqeq7xmbW80CBwlnoewJ6osA0ewKyuV6f++EQfGnXB0QQo85X
L8CzFze1YhSmRBLRtaGkkvHdpW/bzV+quoL33P4ic/lRvQDy7SHZpqhUK4jHOKgw
nXUz2mrQ7g5Ibn3BhdaCPATIJYvLPppnIrg41r9Nzk7KvruGYL6zXB6w78LwXtSQ
/4rttw9YAQPeeSjUUCfc5SHqMN7sBhVvZ1ARwHmXDGCI05YSrt7cqlWo90j8nmOA
+1Up5G1/f8p8p5+tCwFaOjxL7cxmVbReLs7t0CioaZtmrZJsRPEMID38gQhftOPo
EPV3sw6AyzOScp8078/dapokLlBCFSqnza2/reCq2+rG2yK1/pTJtK5fJss0JBmp
duO9de5xsxbRNpa2zQqGfeIriBLgURmf1EoMhYVAJpvOsKMZvaxyeKQSso//wcAL
tja84R+rZUmrcKyJ80aGpzsnj7Wqqo2a8HFt89edredCAZZ+zNN5/S0ASm8APaf+
mqYzMTLZI8bZNNy0JLnlu2Zg8sJnlRp+DWFtrxauWKGzYB09x9nn5FYzF0a5AqC3
vfRbmW6FO0c38wrrD9LPzU570ewvhSMUVWnc9lYpvDtVTifvAAY0COhRVIFRs20k
OnZZamoaSOrIZ0DQ/CI/cQNJQo/4/xdiTPSvNrxcEwwaK4jvvAcliXEpgZVps9ca
ZeTme5soRoIaJSVAzb+S7XCZCseTc3NjuRw2kOzl5LfgsIodEbjOBhNIEJfLhP9K
IW0icsXf0C96Nj2osJrZN/RtvKc/uqEhh5WLP+viCl9W0d6hOKkB00cqVSfRh5ea
2nYL4ZI+MObQ+5pB8zWRjjGGFTaA7wcvmBFFQF5ERpKIoiVS/ttItRJ29mY7nY21
HQDFEuU/HdHznKTlgz7G7e/th9ot6V2vyP30kxwxlUNhKzzxDbYx+p1KLxTvkO7i
MjKpc/JKfliAWKjXKnNCRIf98GTYZU6uBQIJIlR1t+5deCdzr1jk4e+jr7Nwasx3
MBR1z3tkfdHEVlZPFm4nUfwNPtp2R9+pzWS9QBrO0HYtyiMTxacSj0iWQBzX/XXu
loCsKjYpcVuaxOSvq+sO36W6S2WEjQC6ukPg8vDEYaMG7XYxuLvY6I5w9uauZJhX
9Nb6SOos92SoiCCSVejEm0dxlvcL0baHYN0RvsqMI2eAlmFm7uBaNkkbltee704A
qFniYmPxyBJMymkrHfnlCqui5TpW0NRcJQccGPyx8NISEnpnyBBaAbFq46KKHQMI
Y2TJCTx+lPHQFdXtJNVoKUlGma7UbQjqyRYoUKHNUaVVCddO8/KdzydnBhZk+DbX
rs7weiGxDrZXif/JgGcYAv9eW93C6+hshBqWxZZAuHto7dkgy6m6Gl5HvCyKhCZY
NDRscRY5Q0O8vbEHlxW8FuZWSPCHHTPXPAHlZD71B2F+6aXvabjI5HuLAUcVJ6hZ
kTlH4qqNx3EBtMzqfXtO32XT5tgX/SvquxNn6SULwaUg8NZCMJhV3sSEIV3E6VGB
fuSufPEGi6ry57MeBgoan0dVcTtZu/dpRYoYGq59P32hMENePQESZZfJIxdBioCY
ghnH/sJbWfpzPnwWILhz8UhPB0hvqTIZqb3ALkk2vh95UiZC+9YUnn+OYEHt2CaR
o+jTmI1LnZSni5LHnlDRfZGYxiLhmnr0++c0jgJavhTSzFCcnjsyM1xDZg0CURFt
1Gvww/AHqvuT1lwgxH7jpU7B/ihlhs19MIhTFO314ma3EoDrEAceIrHDx31RV9ad
wJzXQUdvuPtihZSwmRpMayFI8UshhP+N1OO9Phx9xJZ7Iv+PryzLAJgxc0tQsfn6
uRToLRoTSKlyroqOCCeVnE5j4HaD5CcyYpZaMWX/vh34+rXtS4BUZvWcHlIoKpon
pJ5K/k4MwFBQijVKupJPkk946eEv6wrD1K6pGjWRBnf89QbD1wRgh/xNSPAqau/1
4x84W52EfzFFi4+6hQvcnG7LjDZV363axLmrjBCkWhG89p9dju3SSVToGZ15w+GW
hA/WUyZN+K2ZCLx2vQn6A1IiMqyHEU9kw/Z7RgYW9URINjOW+KdgPXmWQDoaV+pb
73S4KoydClAFfVqv6WeF08OveTvb/DI02DNf6hJgPrYK3wrRxOR7/KLYxd6V7qXP
4s54nZeZV940mE5TbQh5pq4TvemWc3ZcfDDLeJ905a0hIL0cyJTX88SXDArZcBtw
I+BRYzsyT5yoygTZvOioCRTXNh0kE8pzSBdeR7v5IO5zUlTUIIkAObDBpXtM26PA
XRU3cYZtKmLKPj/+OD4+S73t46SLZ7UD96nqQk2idBoR30wX8aAn3T0OgkW/Zq/d
9G+5nL4nh2+B3GCFNEek8gDnu8u7OYTyCmAeYmB7su5XJxgnoWQQtLCmEjuKciZO
RC7jVFGFfvlIn7XMcE+PWIJUhVX+wMr2tzlkxQIAxQD807mZfp8CA2t1/J+Gv59W
NxaHR85rXRwMX2LEvlpxHPMSq6O2LYw18o4rvxhcvDmtsYdnB5YMvNr1lUwAq5tS
eAqO7TvmNgzbc3nIkboi/nk5jffQjZqHmuQZGJRf7d3fPbQV6AZ0/nbak7GuZM3f
fII2sraRnECtbFueFk2ktaTMzwjEolyzilz7LkUNvkwXClOX0XbKTImgKncztoqi
uzVTaD4wNzBS93JvwiQJk/SGhHiq/FlO2dkUYvwfmtOUj5VHpsDH2lFJB2yQlM23
ynawyX1C/wNAFzjHr2oW/cP5KFTN0zyrPaTTXMc6l0FR2NeRvLYNaZy6m4VZ1zlz
B2C98kv9samCNOflNrneIY6h3hoc0j1Ut2Wl0V3fq1GF6oK6/zK9PTzKg/H9XBD+
06d5j8dkb38J40Oj/GptOcF4JWQF2iSukinzfAQDgc8VaIlWVbDwwqzcgx9caprA
QughTbYadvlQQTpqUKPq8T4mmGWPJnag8cE6i84iLCpIrlXjBdYCG/FzRGSC97HF
u5+EozX5QyAFI4+Pwy8stvd8Hs0pqvVJCyL4anYQPJAePfpQPRR69xgVRLkrCq8s
M+qdePnE2TOjUsbhjt19hbtdBDk82vur4Hc34gYJ6q+rPnfCKm1rngwsfUcj+Xhr
DmF08sGsxaVrhC1YYJcS7ajRxHkQtafj8MVnnTLjjybSzuUd5Pc5ZYTjeyMUCJmw
zCF+mVi59F/mcd+4O27taG94qttPuivenH2qBMsc06N7VvbMMna8ubm2BOR2xFWz
ftUQ3s+dmNsx565KgloI0G0mLUk9uNcpNRVmNMpzrFwBen33NsZVKNVWZ3lK+Bez
n+N4DvVHmcyDvaF1CF2JRbTIj5B6XDzlHjNiN6ihpW1g1YymDxVfmNXcgY6RvKsy
n61GSJIctOs+RNvxVvYMd4LtXcvyLgz3NQXx6aSJyZ9i/L6DDyVZOoxdkUtI/4F2
jqcsj8v3hnWTwbNi3uEYu0bUw3jrDKoIpCqsgIR4/0T3fmgSoj7sLrUHq7IjYruf
5p65BphWw/2SyfjGm16UUm8Gie7eLGGK9PR1LLu3vnZa5gJWh0g1myFEZhBqKbjh
WJuNT9X4qwAUvQ7vKUkR2zy6ebkJUlFJhvSswaNFDHxIPN2Tcv6W/EZ+HidjLUyT
7cTbE8buENKkatvpT9bYpycUxbuMHmy+DvVW4Po/65SyxUlasNjV/NvsY3fhObUW
55SZ8+lVkT8k3YcNxJJexb3Q9bJQ9+0KvEPfTKk82TZT3VPFYG4lCz8541SSzPX5
LtJszPIjU/iHjiPW81BGm6JyZZK+0+KZftyFN8pg3f8xlBxdYQgcLCKYY7oC9RXF
b+XrmvvyBy2qZdLnzSQORrRpbtb4NSqoHzAPQ8izELQbDe55X8FX4YD8QOcZxY5p
SDHFbeAcaUcBG7w2/jdBGmVnjvv2q2uQEaayOKYmC23sN1pizvpydvC9dCP2xebr
jP+X7PNcF8ockw3nWw239Y1kWuQo+OwW37scPAqz9O4mpfkmDq8EeAt2ongfrUX8
S4bbdohJOgZSGSjMKfW2cSKrMs74yrbGGHp5z5rWRCui2v3KRu5ES+C+MluK1G8M
wfmL5KI+bMiNHDN4/jiLqfW7Ldj6I/CtqAIHTOZQSVTMm7w6+/W2srpf4aMzeCBT
ZNNGc/10sZHVGEFcQIxCmn6UN4+vhcwWCYgG5QwF9ZJVpIrBWWy+r/+I8m5FTU6D
kQ72ceRSwiHfRKdtPjAktUyfQRWbhpuKIjU0LhurtAsjTH6Sr+43w7moht41pldF
dl7JIeupDoQxkdZTBHEo9acrz8Xti9y4+A53zqw1y+8g5lbmO1INUaSl9ZZMnBxX
ifh7poS5otQWp3svQi0cHIxdwrGLrMEvVm2uFKq72l75B8QAbfiaBT7bCZFfRoRF
RpDkdXf5WaAMaZ+5thvMTGl7JZgqeQVlZDipwsb7ta4+sGvgwCRprtu6COzSvjWa
I6VDJXypFJFWRCv3omMrYe0xuzm+1KVLvNimSu02PVIxUDJh/ZNkSnA5Z4t+7FPS
KuzxIEwZrqZ4AdHM6lM3P6GWkp4CxBFql71WMPFxMhlHkPlGle80hqUUpDZM3/82
9jlksWi2PN2Rt0Xxyr9Z4cmNtvGM2MB0hHJ1cQh88syPo5RzfOnQLx8Ui7d0mj28
Eq9gZ4ytkmPsfRajG6agndz+AeJvWzYMv3gvwkiveS+bJipnxuKrwwrU0l2480Vp
5wJ6EF+ss9tXAngDvYY7DcL/WE/ngB3AhE1jXseWccVABDpT629Bk4Pjh9OHZQJf
Ui0VCcRBwktlW7UHa4Uvq0/9Fc5qZNRmJzO8U90NP2gTYlJooIZNuXF+k6m2/iTr
4osKiuf6yZqduwJ27H1Ir1Bnh3sc2s5NwZ6hEBYdGim+IBZl2RjRo8saeFbSGRY+
45qTjF96ahIo34oG/vcNq41XFHSLx3QPUV1P8tYq+YUDlymMwMKBYzjQ5ZlyjaYV
ofJSzz3A1KLsh8ONXuYD5HAW7YrXXfEhx6mxYaW5QqSrcW11xUdsV2vYm61WyTVG
x5iVycnt2Rsmwbdey9XqE0ZEzIzqgbWpkFeFPP5JZqKYkX9W3JWKCxg7nSqu6fVW
a9eWlHho9lrraNsoGqc3a33c3tQzXLpHaG7ZMr5EFEPkcfX5X/84TSE0qxT29vO1
xqLBj3FzrNcCymt00ydrEt1mRZweyqbsHqoCGFt0gTlYkQZ1B5FgNLR3S2fPnlTa
Wj8GwHBPxjjZywELnIaExxfrqnHrFsZID8OWrXX4l8EGGt+eY8c0tpMnWavJ73Qr
3XK+bFMSeWoKXwh9uEc0HVosJf2OIeHmWoIm4Cupj/vAcvFg3kMaGFjG13HPTRLb
GiP7Z2OAOtIjlruO97/wIRBL3iNY9o63j6Lgr6qPn3ec3yjYVfpX2h2x/ypmqbwZ
cveX+3vT0omz4eBcWOmw2XJb2JxWffb/qjdcvAdKnbxQbQpYYneCrzKiws/SY81O
doXlYoTHwZKpoIMcBg3N5weDESpCxH/nT1h3lnLdxGu6DqdACuPyh4SwLGbDP2Gq
M2etU3YGdLMbfYqzVWcdF+Q0Gh+9+hYghwCf4K78jhTJQVIzEg07yUCDx6poAkD9
85X4mz2QBGwqeagYgxOv8qX7fPhP3ntadysQ2ly3qEzLcunizRZfqr/G+ThF9WGH
0CUMOWcpKYPvFquYnABnTeOg91mKm8DJb6DxPNqq7bPWLPs8XDj2mIZqFSZsKNKv
+M+qg+MBl6gf/uqIq5hKcMa4resxE79REp+vM3ereixAWwLZTjrQNVmrbM6oQviW
iZuvWtHaFS8nR/TTo6YlNZuR1sh0SGYeImrGsR7K45eF8ZkM6jD5yoTjguB4U/0l
V9hFNeWkNhQM5kP8m6P4x4vMY5MKiQsG0UX3D9Km0RG0kJjht5iHU7vSZfjVBV6a
g+s5XAtFAY9SivRxGPhm1uRaEt84/1vbIpQvchLznO2kBhp2QB14Xs9gJK8U0hpL
B7ndeo/QJrLVmgfyaGUpEvtuxQ8sfwZaxLFW5isgYcSkzbtJ8qMIkW4P+ft3ZTN3
vQCA7sK4+4JEdhC1yvEHLRg5U2zYJKq/zOEGHObrvt/kz3TAbJu7PKHdwIQRc5ly
PeV0/3CErK+6aqESvbOYY+PX1HK+Pax4LI1LdY3Y2nlkR1cUnvBDTs3DyjYc1k0w
h8Rj9nv3FALPE/CcL6gCCLQfN7xAQf7zfNDP6VJMfBhVMrRXMk+51Vy0FLGRIPTN
jR/O9nfV8GNimvR+DVELsgCMyWy6fj3BQY2h3DVfzlM+hS8Zb3444YLNd7yp2LYZ
CeBui/oqKFosl+Gw096xEVdjsZMa12GvoaN5ETmZRaNBtF59pWRxZ4j91qIxvPsl
1VqswiAS4T4qjHXhsK/l4+dEPM1dF8ywj3WCBtFflS1U4WeIEu8GrlxSK7dHQXQP
dXFQbQovr5fLf8RPk91DWG+7rVsvWZ8TTTPjoQUC/t0WXZ4iMFwW6ixr2ogvLNx/
ACXP7ViTosrZhCsSWFaEdzJpn1gMir6eY10yAPc8CZFtUzcTZMrmmDwDler0l/uY
DlrZERTaB13REBpsdfT+DGhD2Bsfhh+4uJP6ZLHOKWzJKfZJypUU2Mal6fea1uSe
uOQ3f+JhFaHuQsiF6uFJUDMrNu2tKSk+0pTJUV7buAQYXhe7kka7u4aBvcu6DyMF
FN0A+iMyqwc4LJCAhT3q5csYArCia36TZeWlMUNDrj2QAeAV8NQk6klMRfKr5sQW
xQJF7lqoWyuTh6fOygSse215MIQn1KTaa8ZgKoZwTasJ/MSW+gA861CYiT6o9arz
L1rolOSv5sPrvDpGmVHGXusW+J0PATbXp/N1Ahd9JLzqgiA2fAGzErn6kxbLQloJ
R0c/E00u4BXMyxD1rW5X1Y929peLZlsPkOGMpFKrsEDSNZnodn6e7xWAZ6IYAI31
VXJNXNKSZ7O+mBIHiSVcejv99aCfVzMo0iP0wU/8ExF8KGLhOcprXZV4tWuxCACL
ty4H3rIklrV1o87vd2h9lLa8D9FbQ6Iqk5QvCJfluEF3hNiKusQY/6ZzHIC8ZZdG
CkIp8G8R2PyG5TNS99rZXJdlxlnspLDCm9LC0OiZWu1A6tuMQa4GNDOD6+j2Pcax
y++9avmM1T9sOzbXMdKAm5Fu5CQ48GvrL0D58IrzDkGCWCFOLSpHqLS9ekEhFa4e
xG2mwfyIqfcRrldY/ZT+ycCgBenS3kaW62TPpB1Z8NE++BCBr6fs72h5+47Exl3L
mfTOe5m+s9zpm/MYuf0nJYwfNSMOc/ytXsHTgbaFCgiU1HLfcV8bq6miz3sssBZ7
kD5jRqH6tYgQ/T8/NF8IvXpsRrAuZ3H5NTH5Sf3F6lEst8SY/lheHw6C8zDKud8E
HIRA670Ci3LRYH1SMtVgm8nSZQ+GXxQPeasDZqwGtLeLykhkUO+EJXd+qI/h0HvG
akUx6VtMT4wFNMdU59fo3BUeQoMGqU8l/I6Hi8Lpoig5FULFG3mqeh87sn0Efx4t
tzrui2SidxcxTmBBXWyYJ2WAALDVqHW7JXGsvvpDTo9nuZL7GkIofQ65IBN6kJ4H
UGP1H24WqtZ3P6qn1TT0m4aJElE6uuVGDFJHPDaYPK6PK5kPAinU4G2omzCKJmxV
X2to+dhi5b17LdVRdrLwPhwRnkeLYnh4aavmbkR5kTLOa/j3/7R8FTiYA6r99QK1
BK9PCtiDSyDe8nvga58yJnLEZ97Uopq/3jCZwHqq2E6lGGZp4rRsSVChnPnNfuwt
vLFHNFYCytfO6aqT98zfugs4Ay6xGeXhI1xisr8a5imJonEcHURHrclIUK6Udkzd
Kz4YIPRYkvUOyE7iQkgL9wP3ELX/ZFsQob6Vbe42Nko3tq+/hXrkzPPwDJn65zTg
nrdsEtOOhJUDynGJCt3Cnblu3l5hEshhV7/jx7m3SD/56ml6wH157hLi1dK4XCmd
ZJ5K0OMnZONJdQaCa1UjSoOQsnqNZXuTiocBNb8SZzfMb8IHp+iLjViZt4fBn9XJ
Kp9/GTMfN2fJwf1rGE0qEJJrPDgWu9OpSZ6gpyMMug2oTsdg9aGYB0CMCSmfvzMv
Z5osID2xMecEIKdTSwchNcIVLWNo1lAIxOeteXC3ce/ymngP6xmHfZ7FrLa38kQa
pky7Mk7fQsjFambcQOs+DWtnyKmqiPqb//iT3K33tsMsUYNQs7pDzLAevojwAaRp
CSucPWTG7hN8CTbBkmzgNV5p9H7IDhD57t6Cm0aKYnE3NXm5YPqD3cJ6yTd9Z6dC
ZxCB1j5ev4zpaXflNWZWGrWSpn+Db3JIAWXzWl41K9d7SYtfRFE6lmm3MYMlZhes
TjXSotQqA1/+ZvwzDpkO+tsosA4PjUV341Bgq5GviYgeoEZBAcnd1divP47g311W
UvDPW1IYKWCUCB8H3FtTj3tFJ+DM25sFcvc7dodPVC35LWUSKFft4vtnslxjBLBq
R7cZx+PjKA1FuNZmdVy0cqxtxXcOVRKSc+qHjaqTA2kOl/eAnX4blaA/yYb0AhE0
x2iNAIEzvu5JvqPhA/nwuunH6XtMYE0pqUx8b74bMH9y60zurlKIbKTe3H/LaG+d
gTaKmBWh6uzi20sVXcbduaR2x3llyNa3C78MJSPysRcfvAVVGcYbqcB25u/llbUn
1srGJ06R98H6A6uxlnrlna66ATKzv9gRYnOl96zJqVBvUn/wUBP22rY1gpoBKNYc
0wPlvHdPtn3ZW+Ek0y0ZwNl0uPTtVRhQEOduHrzL/PLXwd5p9nOXk08UZYpYZlxY
1Z4+b9YEzuscFb21VUj5XNTjqLuasjHALnZRJR2fvLiugP/3ts9GeWjSS/nwqOmH
D0yC3N7UnueFgCajHY07Mnfm52cLA1Kq0WsxAR+vlmMKeoXyHaRsiz3wZNvQp5TK
/bKgHeR7PogoZT3ZjP18mE30hGGmIojl1+J9Ocz5/I1/1Xtl8gCNBUlOYqkET+oO
vY8kjI84Hij2HZ17L8LeZwK01AfE9VVf6bfSE+Eld2YsyMkh8dcXWI68KIHVKk+9
7+IGtChH9eyD8q47Cl4aHbSyGWVqCG5g2Csvrxg7rN3dXJysVfuiPJVoLcrksobt
PBjvwwOaSInM8dtRfRr0bxiWQwPE8BvUIfVifgq4ngLRgcnIvMz1dhGuPwY/L3zN
WBvZECWwlhJ1lIGgO9FxWrnQRfWHxkPYqvGmtRTt2rOQDYGJx70astb/lETl7RVv
SC7WY8q7MxVccPaLaIPs+zeiRXgCwnT7rH6SWfrNQs79Jb4y0f5jmiEc+YvVgJMg
FNR+IbTu0V4ZLA8Od7P34bltDmYl/kpLMwCDvUm5z468b+RFmGhEqbBQSH3HbQ/0
SkqZ2HELkkRhKPvDH6k/5KpY6zvuXadHfgfrmJWqqqU1SSfCEJTxWS7IWwNhMQUr
bB0WHb1KXmMGeAhVfnHyV+VeJV/8nklP0pQ1cw0wvZc1J157/52bhHRyBuIg72OG
pS4R7A1xTLkWnCxva0md26pGPVlTDkWlQvahyuHP3dB/C+2+oIWGQfaJMFFtWx3M
3tsf2upsnT+Go8cgG20LJk02w2ojRAMRH0zNIOkyIdi5Hxfilq+Or0kwdrMSOpA2
86lud6ZS8s43ERJq8HgRPqqsY953RPuXX15rs+d6vpDRHaaD/WkqtlVezRIMNWgk
IUabEXSxD1ajGWJewyAYhd66J0pVPR0PqxkG8wguw7a5A/nqcoAPHBifrsipY57r
PYZDfx/hc4mWuEYxIgCkllJkO2mJFPFVc69xYHQ+KNFPXJcUIUUChmXcg9ub54h2
eQq6Nb2r4fzSBEYNjVLKabCvSdp8MvHx82HC7neYLeHjaDHOZHIi4NEEKCR954H9
JJkLrrvqsCWK8wdXyveQB8PYfZ88tLgwHOdF3HAG33bi1Jn/Q5HTmb621pc2gj8P
DDBR5DEgcsdXcyz8tdLZLZo4/canQzeNEgaq4qaxCdFYhRyGprbulbuSYZsO0M5N
GVcpMQtcAHspUh1gGAduiUfWgng53RU3vp66PSerx7u+RIRP3+TkVqCu5nPE512a
KHUcwThynAO1hUs+9dzVpmn6wt1UHZ7CUKY0a76WRsoqf83HeYUlbhJqE1NWI0y6
3O3Hvv2nfaRiRlm2QiztPKk2qLUgBOfAxfTkZrIg5/kA7M1tOKoxciZXxA6wHywt
WiaCWvUz9qS1ZQGRnsmkDUEWBtoMEwQFM7q40Jt1gLbLhABlUFKDaCBsoc8zdTaz
lxHvq8ZSTOUqxcZUiJJQr03YPeswLx/4HRLUHUqlKEYA29Jr1uWppiH//esBcpns
vk5c244jFp95nr9jOG8WSEOUQPy4i+BSo+mzrsXvjQ3iDhpiKu1xjAMsLxBkmtMl
uvASZrY4TMOT3wQ8TL7R1rpFpVRv/w3Vomg3PcsVvVIML84d/cQOE89JZhj31Kfu
igtRJYBtZ0QjdFYMDOj976h1UmwP8gSlYIvX96lMlTRsxjmqihUJlvXynel/m90J
pv3C0Hx8ntw5Vb8xt6jF+oQzOBvgKXzTRhFbd86x6EWeKaLHySIFuEVyWZfOEF7H
1iLuIVIeEcHYbOOoePS0Nl+GIftIjeQ+NsQoAfOS8fvMgUOkJBQ9moonC0vuXO4w
BJAIgMTAWUXRgLVCrBZfZPfZP3rvEB4wwBrgrUF7f6efjB+XI0lGTYbKTcq9H0AP
npN5QAFiQDgQU5erMCIHSmCmtC2aA9kHo7/XeJdKtErT0DCDm7nIPA+tjbogu8W+
zZrMHy0Vg6CeEj6TyhpVqvrBemsSiRNHpir/zqqwYdPQclLHY6LYVO3hpvAxqkWg
duI7M9SgNntaZsqOo4PoFUitx5XS1vKhoDvjdldO1oLpQpYJSZaV2YSa0TLOKmUd
f/7CUDR98iQKKBLnmR8MCRstcROprI0EykEXU9gdt2C81BN9CoZH8MGdGFblV/22
8GOZQ9J1GfwnfbTtRlkFWjqk0xsAGkrVJnS7JG+BzLg1nXeyL3R2zbJlRB8f52qT
FiAKyXtI5ks+F6/+DnHTqlwpKwNIIDVfEJYShoWxgm+9slG6UYb5AOr0YKVxSdjj
w/HRFvdvgiuzofjif2SsjiYqDjz/4pc6wzGmCAWHxGYPL7rRwjb27p8zThd+Ot08
0utVkl3ST2F0a2eDd2Tunl3vUcwlEaAMHZCUS5TRQ32ZL94aV/B4F84hHe+2Vr0g
lv4rGIcl9U5zUdETom0DdjmLjyt5jiz/0weGV6YCSIxgPMSj7POF+hfDabBTa6b4
LvP8HQZPtd18IEeTMrsB4W1kUVwUDQVaC7KwR7yH3FsGmE6RRbikADbYcP7vBtiP
IMfip4ry0msXX9qfQtejRvcQuEGXUdveAKiLi7c/NwKmZN8ECjUtOAxTb7l2Eu1o
pW9L57jWU1J9d2uBWnfsBf57i8upTnoCfUYQdR58Eo/nTab+ecNq9l1JjNjZ5QMP
eVB9trFc+keyNo2D5y/htKKfchHXGFin36zrNMBWeZ4IyVn6CZmBV1y2t/VGJPWE
8GMJH/TnmcEvb381gjZ6PeqIxs3loT3k8p4T9rwjb87+3W4KE7JBw2Oz3RFwj5n6
C/QmdFf+oGZnd075Y6V5c47qvkpNHKWFBWsg2MZgchFPJuvtPPscNu/DB35/34CT
yJzO/K9dUAsHpHwu73QOtGIx1Xc0BWXF37ihs4rbq4OZzoQWY5vDgQidQgp/qvez
NZNpX34IKvlppVPy30puMNIk8X2HCmWFsz07g+99KsXQntn2g38eOFYHhW/xvIWo
z0bKwdlKL63ZV+eena+mNGirTnzPWV1c3S9n8vYtPQyaT6BWMffTFOL9fjXPrsSy
sj4Qzhsu/Hf+6iMMsypxCutIaJWcpqKytqI+SZE7+bTQu9BvBV5YOGzOdO5q3TUx
Y1J2HVsX4AxnhtgBZE3+WNF2tNv/yVe9OMHc2JTB9NiPzVFjGKiVhxsPhAebQxma
RRHji/b3CsHGyfnLA2Amnu71rkmDmpQ5CExSmBoFz1zsbjUukHcBqaUbJRrzf3GJ
UoZvwFJKdwlScGdLMPJwBhxZXVG2D/LHFWoD0p3eHCI4/giK1Wpezw8naYIpiCa6
81fOaq31PWxxahnJewHjlUFvyO9j6XtkNAkKb6HHPVqxmmKhlR26TNF1/bUNt4Xl
aGPR/lbgyBnWpt+3jmilFX3v0opfPYZz1jrHVNv2sO3z17jGaCPzrK7Sjxnl8JL+
zuCS7uFyzPBYSYsQMweDVlOhlVKKC7C5XBxKmtReqg7YgXOG5A5ixsRaNtnZfFWf
DS/m3G6bttXyAOmD/4P/wCEusCQ4fsA+6jgTpOvEf9RbjTIO98suQyThHfcShRkL
0Z4j0IoL3t+82ImnUrGS62QmKHq8TKfjbss46xHkui/N28qM1J4ifRaV5l78dezv
8Z4gYaVhXxcbza1Wqepr46swyjAp27FD26JG4hRgv2OPfJNztW9EN1LtOnnql8TO
Oa/5ykgin3V1BhBlbj4P7XPd67tZ1OMeT/rAAbMiBNYILFNyrG1263CEzLaluUnp
iiYC1HBMz+iYlyI2tbm5/Ee3RJNd5CzVe3ZvmxjRYsm+7cRoLbmJzUWl2oqxgoL8
MuWFUswXYzBeVRiHt8Ge7yDp+Xiqn7gcpePR7gKoH4ycA+wyWwOYIO9CLcACFdFK
vQLYzj+tuLTbRsaC/sP6TZjgmC5d5YOrucPpq3L3S6iBPuX3UAf45fZ62tK50uCe
lPRwXgg2GZgeoAJgAQzR0VhIiy6Hc090boidnxe6i0MwmgP/tX24kJ5NxTwSfvrp
qFeyOVFnDMXZeIBNKfgfx9aPF7md02b1Q2HRZp/BadKd7PJucOHYbBvp98KPBz2g
K7siAxQDJVzCnaR7pzvesD95wks4AeJuRczcongoGmAk+zd/nex87Zt+6xFxZUFS
xw9N/ShE9XjiM4V0kG7rnR1NZfwKg00jYkcDQqq5/xb+sKuZ3EpDzteZWV0Tb0h/
QIZYgD7t2R3F81VAOCCGm9Uhu7N8Iwzis6nT/TEn2ZvToCNsfqwot0oS+0jtFhSb
gla2GWW8qMHNvJNu9nTgJoz+NPMZf/n7+Ns+4sW3v/Wb3Y5IyYcetdUCvLEXc/1f
2tlO+7xA9/LMr4qIRPme8oVEw5MIq76KN2cJl38vrBPK2O4D0aCawGb5FYOGHaxD
t0F79rr3J2eOoj8j5SGcdMSad8QMupXiKE19wDFRRFnskFg0LSf1eKUColJ5v3FF
nNCsBRkLpur0+JQyX651xc5NtlkRKqcta15Isah/Sq3YedXxlk1z72IiL/BUii42
bnE4B+vfjO4tvqxpuFXGCmue3AE6HpWf9R9y32V0/I4Ne992oW1tYCeoBFFCRHSX
Qhj9lbn3UrZ6ztKQXMMl/mR1IvsQf5hCvxhV7rwagMySIl869a3XJVcermLJ+reC
FOxoJCeM4DaWPO2UnLVT0rj8ynARQW/xgmrTwpfTZ+w3hHNt7Y5gHBR4+2m0ZQQ1
3qornkNRPtbho3TEIT4yAewGYeT+d7eJBjDowz/6rN+Rryt/HYDQv1seKzOeVVLG
9HVCYEB9QJ2GH7AmbA+iZIbU40d4c2mMFd7kAEliAoOIlADlF48X0u9SbCOJ5U05
njTh4JxVLPnWNF23d56PQOJ9fxxrBeGQJppTtENrtEKWsQx+6ua7kOjXFos86uwv
01ra47yxL9qA/ZMS/O24tvKyearHwUDZL1snv2bsSA1uXRvsZrWtbuRWv69lPe23
igTnpB6fo4CqYSttHmtTuxNGw2YD+msiENwRgT/UZvi3CTSzxxN2SUmFamJ3vT1/
liMwqD09ANNyJjHxKUbtGdS6iitz1QcOrSVOWkn3t5wfxhi45u+f9QUoPbBNYJoZ
eMV3oJrxqS7BNMjxADX1NpA5lXmkHrcuIKNty+xykXrLEHJn6+Yg0gs+JPdq6trf
ZNk12c/HPy9LUqU1Y2y4MOaspHKn5OI7TOT643PYmbHeav68hul/csPQJOXR0C8o
d5IY+SNLfWHckW8k5Nix1zdcGyROgsxzufyZPnW2i4v5FtoiumPrNWrL2wGlgs/1
35EIPQ6J9c9EuPDr93MA7MlpMw0mvCa+foe8SnA7183/Rr8O9Yv0llrUByBd1/Yd
Uy2p7LiI/3PmFXOz7D3VS45Z9ILJdufSRF0ukmnD1jInNDueQzRJhlSkb9m/i9o8
98xyofjuNbZ0HyxpM6WV8c22Ds1upUwkxMgVu4mg8j4FQhFJURttFF1KpM+j8Q7+
23HoD4/f2nS+GTDm5nNtRVjI5gfLtg+gcd4NmowGTkrqyqHF3S/MWiSjFFChczWI
c1gi6Tu1eHWv08NzIdqJypVzcGx9wbIobYMU9o+L+9rXoiPMZ+KcBYbLtVbFoYkx
hBtTYMw/gdEoPMuQeW3UaXKzenYOVH5ebRgxZQ2MrCs7H6Vgklp9nA1V9eZCSKwE
c/gt9rXNkg3RabklM/1AL0W4LOQ0Gyyye+4TcmASjIKm7H3NVS9MXoWWqIT9I3Ox
shcAj/nl2oV5v4yYIiJL/dGHf/W4mt76KzMtbFpSEUy+NttgITciihpIpy85Xi+L
zdOq5Eu3QHkx26DIFNOJ9pV0U4Spqiy8vJ00/kiJj1Ix3z5y1KCp6AkY1G/DZx+7
fMGZWs5//GwF+8V+FBEZAKufvgzYpPhrXm50KnlY+njPy2KCOA4FMYpbfa2dRe8q
DyF8oY/MAH1uJxQYyOndaHKI/zNOoWG/KfYcK+HmcCZSbwY23tFVjNqkNkXCRgPe
+IKn2krLtng2VdkYimfPjHxt/Rip0glNKa+9ZFtJPbpWwHGYJ493NH1yrhH/R/Z0
JfsmDSR+H3ZUtfbWTT4VvobxQ7pBDUbjHc0glPmzLVKWfTb4SvSPxL6RaGmCW6mo
QgCu8i5aHG5CQ5uNtvHaciI799vsWZAVEyDBBHCsBlCFMavgTgC+2vRpLSJcvp6B
zoCXUygASCYmz25mY9idwLxPfDA9F8X2WION7BJkTb+6C9RTxRwAYlN5mFGF2dL+
J6Jnf9r3GazfYEJZ6kFUJpe85LuzA+OZ2tMDfgQ/aHBoJ/WUDlXokcFRQSdguu0b
l5+/G2z5KS/UQLNiM9bH8S3QC17GCLoNbQEiEgsl0Sn3WZ3joH7+Jeqaji3gTPOe
mtCdVEtcwbYyQjl1gtXxN7cm1pFG/VdGw8kbxkbyGDZmxGd59GAa+s232rOGmU2W
9L8R9xZ/IOzGaHNQGrj06/6xiRni4jTRxVI2XgtTw7YEeHTnU9qdkB3qbFvgCj1k
KywtJuXBdMPf36LynRYuWjB4P+/HgHk2/bEzMkqymyM3YCqo3Ycr7eXdtBNoPlLv
PHQPm1yzNShcaAk02l/2FlyhJH4ofPhBQAsJnFc85qwhf6nZ8aP5s1UNgCJN6RAD
t3a96uIbPn4esycbMdsFxm/DKl3deuX3AAbYjxBqzC96cUa9VtcLV2yrDln2Ymib
p3BKDlByHiU0A133DXQYx8yI2UzHMV4raa72ImpKbWnB2osIKhYlrC/js40sktS8
PMxv/KQaKV7LtnIW027sj3B14mXOi/vBsdwnMbf5tqJLdesvDhEIrwEsJo9qrox7
2ORGtryuiBAzNkvaDDG+a+He8RmqtYdA8/IJfxy4CZXy+iMU9Q8sGiKsPMYp/r/Y
pO0tchtMikbWbwh/7RRGRs8oTV3RkS1GdOePPbKHInvB66IWIecyGKTEcYX0vCL2
jgx0S2HZSUkjSOjaa0nWZuhMRWrre8LaapEt++8mMqxotX/KdjT1aKriMuyW6/L0
gBpV5Xk4IBPiM+NWWIuQIzfsioVlF3/zt8hMAYZZ0uPZVOegCSrZ52VQtHFRujyr
7QKnEvf7djg1RQ9S58uClV5Gi8rIYJ6j2NrOFmKU39BkcNziiTQU1FpjWRWMsX1g
ZowQXW9IPqSB3ROVn2GhvJ0bRfb9InO1Zg4V3ZYMDNFNJsWB5u+Hc3ZcJVyfpFzR
32oIS1XvjElo6tAkXMoK6xxMk8bwiGb8Wcxte+ylOHAMyvajHlrE5Fl+cxPbRGvX
110W1jrvXiV4Gx+JZVDVn2jgYafqmhmmWGRXhY2wmYYbguM+jd2yjQEmkMJ/SSMD
rDZECYKWx1DnK51F2YAs4yOWm9QseVEhHGBFFhDabHWlGbc0qmBv5vgw/c0AcLlF
U/iwfz6Z8IrBBIS3MG/8GTKlyFJCNC4B2lTBwhdRYOS47WzbYkxY96K0ZaeJJn9k
NbgnIv+5HfwwRZ2gkfUAOK4p2pdZSmDvIssIuxdOEtjfdAaZUcvSU/Lmv+15WVZG
cfVdlmh7Cv2WkP4evX8d1OX9wTDDzUDrTqEcMo/dU4+tnCfcW931N4cw7wqXLKBO
gYNPbNJvBbKKDDRxk/kwCoCkq0l57VlCFfYlwV7x8aZq1/Qj+S/z3pfASb0YIU12
AZuvj3yYXVz5Hp8UhTpS+iLfYFpT/HTfih1ISi/mvmPIju7aqOxlurDSDawxppum
p9MXYM3h8Es6JOjtfG+a0vMJk7FZQ4LGUfUtBMbJiKO70o4VF5SQAYSRCzB3TI39
o4tW1iU8c2bk6Nn6I9p3T4FSJmbQ7VH799u8xdSfj0X3x83lcpfWtj4bGzdjh9ss
yruyRZwnFG4myhBiLynCQBi4/n8+cs7BfvNpqhEoYfW0UMELEse0B+jnMAmJKAZY
0mDXV0DVnx/qRkBptqdU1o/+sxqxUB+waQaImUGmtnP+98Ylr4xKC4Lz4W7Tme6b
7q8UpSDXVnP2a84a5t4W0RUVWB9ArxaVCICu4ckKdGCBWisSguXaun6KX9oejG3+
hTeKu42sMZt6vmf1BURCu4srA4wmk8UM6HRZaCjACJMFyzxPyTV/Hozck4LtcNqJ
TWeoLZ+1AzNDgVyCfKwcaZmkGVoXJ27sCU3woPmmpxtm5N7qZ7lPFQJmys8fcAu8
wR8gDRRUiMdezB3enQh8Qrs768sgeTz4eOC+4AmI2PHcDAtDn1bJfnjkxEcPE42w
iYLJmGRu2G/8vSkIMjluLXezT+DlRyBrQSaPLdfZAhuO9UZs3uOIjVmnpW6U9e7c
hQHC+FaLbsxUHl2yUIxTss07C0pehfsY+XcPcgQKm2qULSmxRm1sL5w8bMsqP90V
xqmjk9iMhKVpNZS9FGGiATfYxHIdMLHWYBpAbm07Ka7rEVs0nJ1DS1/UGO6w9zXq
BHSebPpNyqE6XurVi/tgNfa2dwW5CINJleX07TFtrqTdPOQCL5YW2HZhTYdqELJI
dLNqovjQFWT7XTmHIwj6b1PrBAVIjFz7JyHSiW5QPEvx6GB2zFlEqzEemyD/gvkp
in1JoH44010wM2r7Prm5kU36KrZjs6r28ER2o+wxxgz0AIHb1/Ob8vxg+npEE6ol
LtuLueWzdTYiPubLS+kHjVf1y3QRXt+QssC0Qy13SqZt8nKLkA1ugfDqUVARpnYs
7X9BdfNKlzJ2pDgOCzKYa27oBs5kOgr0iCbhr/yGV0ATdI6wo/2Sdr8WBiyuhQ+X
yNA3Ri+iqxFH6vf63g51uiF7xoESPh1chDH0yoOq1M9u22RUXoDGLsnaJVSuGr1o
D/F01VV8OvS42vvOuale99cv5HlXwscpmn1LzJvnosEp7BNyNEadCsT2Pd9MTt0j
kW3jue4poNHeFb97+nOnTDSgH9WmNX8ZXwfpxDGa9RRBoad9D8E2tQdLtf44V/OO
SHHxUrKIyLUSHz+pESr8DdBu6J3Xtc7clP1P7ZJKLfgwj2OuAjDYOv+cmCG/I7v2
IJQ5n0ly95/1tskLwIg4wct/kXIxUK7i+6Iky+NsHZ0Z9GjC+wuzQyYHyLT/Rw4X
+b8NNxp3fMK81gRrnAKTFynh4n8yYI/gI5+QoaOAExnNHLXaBgYKsILiI457jjki
sVa4pLpLfiRJJQieVHokfaDEKpvT9Ypd8xLtvVEQYH2tYWbDKvQ9IJBZh8809JIU
i0vyI5u1jA+JqiGhsVsCqN5t0bo+IFLJW0EYV0h0PpTkshq/PA7dH+FTvTPEeL3F
gOqKAKTj0QRUbCsRMM1nwFKF/GiQZjtcvmQDa6LeBivrbLRDdgq52w1/47FUxfcF
Hgj3ed2R3mCSoqr1N5ZmYUuvdh8Dzk0Ro+jiEarcNtufX+LS37/8ALSATcqsyfdW
yO2Ox+LOtAE/q8WXjaQEQKeKFCBXx6CUJuoyDC/P6OEqvI2G97o6ZULYtH4NzPZW
5FkMyNNUzNlcBV/oOYfP6B5b9IKEPBaNc8EUU4J68+85SfZ8deqF+yYCwo6NlYYV
xKOWaVhn+ypjS2XaGhc7/sk0SeLLCoRxQIdQAHGBdy/I46KvJ4S9UdKQLMo3zTZ1
T8rRCNevMn0aaDbXUpAe+KsUEdJCcmCdm7CmJV5rY6lD7Uyb6gFRbQsa2HvTbpeS
6kW/b7Z8gHJGTLhTfFHolMb6+zJgHLUuZE5Y3fSUTwiUfnfl1WV3KMXSjKUp95cL
AUSGf5DxMyJjhy5QSir9UFDDkY7j+fp+02oMUVaRb980EOnQ5RXZ7U2bojpMkcwY
GTHc5naQklYcHj9g6+77BzG1nqSVbCK+7VoTU0z/Uae19I1HZS6RK6WHDmd8z7e5
0ytBwv2MP5VzCmvuB0RQLbj/pr44BdYBsxst5DDBs2ARkdXrAi4rvMIPDEoIbzni
F/+0F8YuYfPJQ5UlaCja0UoRIDrjuUt0GRvPdEo0vQoHxK6ZLo8NjmW6xTCAgw3I
5oIJVNgiwB1HdV5WUF33I2XxIoiM1piGTPD8YfatkHpOXvMKGGVPyoOz0hLi/x+z
qmxglnrE9q5SRo/ggB/QpoLlUMaT8CXMMjnvwWuL73XDg8emFKvz2FO2GBbGfmGk
aHLZEKrWYtTRzIz/cGFLbuR3Evwpby3072Ysuu38EPYmU3iqO0Ogzj54ONDqOV7h
oJf93IHlJ8/l/HeIpihFzlxP1aj/Xrm7A9D9THFC5X3YM1/fJAbZ+iRCkUPrYzls
43Srl/4pgvLJ1Mj8ovantE/jZ1C5m/J991GrmmyDgB+tWnVxFGo0SdbWHtk1Z1z1
UjA62lYVP/7N7PziCpm8oUStM1vK0/ydOdxLkc6awZ/p7Qqhy/Oir8iEwEdbGRKB
wNzEBD0nSwJGxeBcMwRQ883Cz7VFb3iwbLK3dz1ETTmXh0RkGYaLIykInROd/HoJ
5r5XXMnPhuhA01SdTmOnbqNgdWsMAp3XUWqf1iV4msgLt8B73yLye6sT02gD/5HX
7m14iyfDz9eR69oB4PO+67XZQD4jcp3T+ZMZiZAFJBVA/brzTKZpBMZKGVxpC+GN
W2wiRcfM2OS8Q4V5FmBuuT+gMLnFI7GYhzPHqCmTP33FLIYjd509Ks30bWvrBMZI
CB1lhQzG3pOCqN69yS1DfOgYB4sGIi5XtxGJlSvEwQdpI5mVC6QNOP6Zutw+OeBF
gleZY0C2fJPr6KXXjjQRe0ImBgMSjYbWiK6OFIoq6Tx4KeIhQgaGjWgUK/zCGhxn
EeZejE8wLYWviSfEOnQBtzv4n7JVzlZYSlfv6PB5KJgaMKDSnHLILMA5Xr3w7jet
teIUpDwBlA2jfTn8w1zfVSWWJilGi98PiH5gH4pIwmN0oBr+eL67dYUcw4nER9JK
qCqlpZ5OtzQBIgi2OMuDoRfg3klH2lSNM2yofnBpB2PeE6iz/szzES1kdKMVoSW3
1SoF9Yi/IleIHbY3n0Mn+N+Ba3Sx9KOGRKA7t8O3ALCU7qseh+nzkPUmP9Lsy/Fp
35ii/8iVvDL+/FfflOEGCDEm9xsL8OimF9U/udUfQUop0ThYqX+HQ8D8y2pAaLLc
llZgxH6usJRkDJDPBx3Gk932BRhugEcWkiUyqg/q/N27hhWFE5g5xSvKXDFbCU4B
kI4vn0x5St4v7qb9lIAarZl6jCnykWONKVow4Bv3c0cLY32qLJ8RxuLDYpuyrsJd
JhLDNz37pkQXiMnesemuLqKh8jWeQJNzoLC+0rPsvAy9C5oh9td31dPsmpAQkKz4
gHkV8V+2CcNK47y2VjH3XucH7Ks47UpX3Q4MbSNhHeytLyYVKB18aB1o5sTEF/gW
IpXO0Qqa2P9Fp9h0SJx3arzDSz40KbGmcE2kjh8c/0WKQ3e19LF/n3f3voeAjEGC
fs3IuPPbkuUAPV/vzpHnEKDZ77FlO9rT2I+NOUAb4ll758Xa6VDQXKAbiUOIr5Os
jUT05wAzwF0p42kyOP9HrzI5j8WkGV5JrfyQe/8IjfhceFlnmhQObaAkiFk4zjnn
9zQFacOacOAICqS+6UtWdAuH0sBY0iars+A6lutDSKydfCYyGMpN96lW7FVdR4iu
5fnf/skDNES0tLI4jOe65YdmZWKAdujxlDA2RIqqQTJNPyKIvk7otrS7fU8gP1c8
KYdm04lWL90OUVk5QOKrVvLA7xwNzCvZLYWyka0hozw/luCrIEPeG3o6uN3+7+Oo
aU8R7MZTNmG7VzaZSA+WDdBtpFD9nWqqVMq78cmpNFzWD1Q+xzBhA0k7LLsyPnmK
w4eoVsrfML6oyXNN7XQA7tHby0oHH2a5fRl7XP7k50jjiUahb7IyobF6YEC2xAjn
EvPgQAFsMXpcvRT7uq7s4fkEg8YJZPKCoS51+zdHtKiuqJAT0xoHQG/4QCT+oWNa
buSP/uvY4IJQ16fN7TCBUKQZu5RgklADCG1YVa3wZbmpmABDjUunmNLf9dSf+u3l
0Oj3GjVG+m6gbOEFWiT6jnmOLVjNpfsMEC14OZ2n+crQSlpBDBtRw78jbMH4X57/
oUnIDo9fQSJlBOtktK705AFAm8ZD22aXcJlNsdqeTZiW+ProX5QMuZwAEfpgMEEU
DaMIQkWcFzM0uSy27DdMGe1SNILmmaAkzZV4WGvshdYLFutOtVqyFBRVTf/+7l5p
07Ik3XW4tc4O7K7NpNVLqGG3x/yBxaqEtUmrTUmaSFumJfZPlwr9ikf3OvK0FvJN
Ke2wHzpxggBAdCBLKbEF7lOEb9grHJCx2+0iamDnVBgXJKeuK4LPk+Af0mAZX74E
gTm8cWt0ZpjEV1Xt54hgQZKvR3PDApA/g5kPwyAGEyRSgQOrZmxY3C3+T03vPQEB
5m8fXl6ACOZoHdX3iklcddswSSKxnQH/eGtz77GJdnpqWwjybzBHopsIbskWrgYb
iPwJhbLb4frjQGK40EsgoZVHxL2WX+JHMiuXJQOtM/fqRoh3Zcws37ocdlNdgMv0
L3mZZx+Zax1KoqXho1H8mEChI7E8bKgtuvV3Rl3BYfP3vYcEmzsGakBVW5D+VgKS
uEKi8KeOa3IxrYtq6KNOh19R/SAWOtdi6Baseouisq0sdSQPWaFQ/4QdxTfkdcke
uTYTq/UXnHCQIw4NlncxME0HjkeVYeYPh4U+G1SrdKeDw2ZjFOi6KoWc+LipCoCe
o6SlJ+FzYeHDj2K8gUxyseuATrutIqQfpL5JU+cBzhIFfrCKORmNo71JM/QCub3U
0FIAeByx7zFFEgEqIMHnSo3NKOj9kdH089Qhd4FjwUWG2RyJAItKUSQgsvuYXFOd
cotVxsPS4kzFkGYdPVxItEZ+zxZ7iEf1CBv/109S7RDtxH+D869AcVcWrgs+Gs7m
72UNMdLSWjP3utsaYxbOPSvQA1G2Irg5dz7YJk/7Y9nl7bXOLG//uzHlUWrnBfXx
4Hi64DSm1+ywNwEenUBMBYpdIeGmp4ZTcacKpHXeke9/OcEFQlDmcsjayTIbdMDh
904pZZGHwQZq9yRwci+lmqwZexk8ox4iCLw8hzfrVglaU3GOdSTInTMwvofbT/a4
6f90VITO/QdUHRFC3Lbu24N6SIhhurKtaNZv9wLupMDqrFSYlbItBkN234ldQfhb
63evmiMEDj3sHEagJSq5nTPfjvPEXaj5ImvE7ZT/LycGex8lJQeX5SHtTL6fkEDt
/5hu9e//MaWX0kIidS6zLxSzFig94Tvk5ar7QQ42pQbH8DsfiXllzn2DmC5n56O0
SCMfoY8tM2yoGOouAGaP3OZKwX8epmVaggeSME1N2CZgFnj0Fxyf16x51jsUSIkk
nhA6Tehuy7GHPqRHW4uxS8tCLSygCrq2vxp4Qj/4sA9P/3B3tpetWUzYbMZv6opp
U37K05f3LHBMtjLmgU/kSk5zWM2Zcao99kjhM72fieAE/KLkm4RV6OnTP8KE/WN6
AJ50GidJ4J5z9xyPGt64Mdo5oEIWF7QNqFFGPD91Pf7aDCWjixIkjq9/nOUy1Hi1
/PLHRQcygQZ5WZ4I8X1iruqjSVSrRzhPm0yDEIBM58JQQ4ByVk+RvVf5vOI+AOaM
WMCBIRTXBrAKdvZbMDmx7VMkO24Y9ypTx4ykppEfhQPNiO43HUiE54VKOvInTym+
9ROILit0xruZPLicyfy7Jl6hvS6/YWDcehQlIxl3pnolyD8Ts35xuUR0zubadjfw
dSkqPbc8XtoUCbVdoQnq0wYtMot9M864PCn0oAhPtDalJBKIykaf23u55ZwiDuQ8
9ptv0UVkGAwbf5Arus5Qlcs27rvN0DT+5dt2v6vqye0FU46QiMV3jrXZUgx2SvXz
YI7NHzbyOW9NsQ2pC0VVvhFWCziN6CLAnBLOX67hsEXeRB1lv4wP12Nj+us/4T6h
nXS398SLMp7u3AESa6JrJHMhHQ8UlyFyABFNSmjeahlZq13BMrU9PtUrwO5eKsD0
l31Msf71nFNhonXMMZDaXVFrWPIJy+/d8w17QkLYOhNgQVTZQSxPcU2emw8qpRcy
fiVzHgUC3Gx08A++s22sNGBszGSkT8/JBayTSQHuXXgOCir0nU+nzr+hV7MbARTy
Hcg89tPOJuC1kVKO3YW5a7FONZXFes1uQ8Ey+3z9l2KaRG4XksG+yAMtC3IoK92B
sy1b3Olu12oBwLByKfmU5UiM06kLwKa8OylYwNsAQZAWxWRguKfiZLM6a4Jn2ecH
JuFkGtO+6GsHu+/LeQBXkfjrzFnk9Wp9rejMHfXCFo2Gc5TrHnROA6NEtkfergqm
WwHo0jCa5PIypZLHc/9SRXugPfGHPjG9L6lp0yYbqjPOIm8wkdpxeN6SvMjqtJp2
iLLL5tzgXuI84lpAtHW5XEOs4BOHDOuRUj5TCUNxpeGDvIXYNtV7wHOtWqZX/5Mb
csPZ9ccCvWYOtolvLXSHp/VcxznSViYRnifHun+uh/ZMPSkBJI0pAc30wT4J8fn0
5q6I4R9b7x9WHLkEgW7+wDyOlaz6eZL6NKl0rFznF5WT9A1UWWsXsSIUTp1EqpUa
z/IuDFCaYiWisojFcmsvBL931iuGHp0UTENKjtQvCKFjibI+7VnZ9OGck0AQpb8c
mu11HpqJ5Oo81ns9U/sDX+CHfvzwkfQjzstJ30IrxKoxg8tnsIvN020i6TJ/I4ik
5UXdalA+ALQG+F1ykMIOXdQvZj4AwsrmfLtKFRNNnvb5fKa86YeRkXIR/VJz4Kea
mJ2s3wCRL7y5nHhcaTyaMvXZwBBQr+M/2HQ7tICLk4yW8MTy/LO6EHFL5ZK3+PL7
RllhYT2zn8sWX5wzxQxRYRNCGkXoQLxko2LwEVQcG9nLo4stCLNJ7t8NpzXStS52
ngxnqhxB3G/yN4vMDVNRYHjdDwkE9n3XqnW+gkRa93DyFosd4Vt23Hxke98yIgzE
8K44zB7PfqHRU1r8INHILXpbKHTBi3IfFTj5EIiaiCIibdz+VMjcSRBuaAAU+Ny/
Wh7H5mRzRoT5fboyxviU2W80sYg3TfwA5ykXDMTu5P+ADhc6bhRwYwZTxUX5JJp3
LQ1ciL0Kh12BjOMPpuWWB26xN9K1wnSWm/FYzV4JasNzB8l6uFE89TcFkaMooXOf
tUDA8Jtmhco/CSxzrmtNrjNP0uzLoD2UpmzRXtbdlilpHy6oRmCOnE/HUzYdKxFq
C75FTtQiVqAFPvdOw0eweNjQGXTQxAxMi9vuAsPSWJqu3XwU34t7/BwNRZD7WZxX
w125qdIu1NBPN0xhMHk1zTJnjamTRBYZA3YCNvNpfcTAUPInsFrxu8ULOI5BObyD
hMr55cMVChtW+rLVqoq+nXwZAz2lR/ydkDIp9ZsvAnUliAZaiEP5kr3VVQLDyKRR
UTkVlpZGOw5Ddew5Pn/I1hecx7Z47KyveocZ1e592LsZPLVFqf3RdLvPBtDWFcon
GKr/V1LuajpLKmGnzYvovyqUHfHfNu5rvxz9NYj4Q4Zn6/evNjBEgoBUcXa2b2+w
o+kNBDqk/5svjbcJztOLbp1LPVT2orAOt8QYl6XGo1b5+UHc/y6HoR2kAUdNRE1j
ta4HhHhEb0asyUOtV6pSO7BYjagLWV1c3cDsdNPd019N9kHVBFGYu7AazSfo66F/
Rqt31S7BfFtMykB2NNegRPxqqwQTiegL/lYiZVgPGiBqiU1OwThhm/5gf/Sl1eb3
jLvkAGccOEg70zVoypFfN54mmrR5KPILy+9mVvvfaiWa/Vlq8TWJpQR3eBW9kTQX
EribHKzNJIw3yJ0NZOT/hyy9aD2Hnf8U35rcQxSblbVx4ZBcVbL5ZLx1A83Itvlq
i+hysPrP+vcDmwRPzcL6zdXHvvAZXSp0XYRVeRRWkkS5L20q2dzzDL/gwJ44hLNG
1q+yt3kPR74KKrSia7euYL1nqYntTSHvA3GEmRRgL98DJmCpen3mUrqfKDYzcMZb
EPlEgL3mdzwiPIyw+h8W3jLpVXYAHjNgVHh/UQObL+/kfy6qKLS7vut5OLPG4wpx
P3zeubh42volQCh8L10VbJc4Qqx0yygX6H/T0fLOxaCebPhO/zgQeV3Ed6Eiboxz
pjLvEe50eBCn37Nn0uGjD7lt4+kkqsGqNojwDklCp5s8JytOdBZfaSqY0T4x8t1Q
Gljk0Rz8S4ctZy3UvqQY0Eof1Sdx89uwbvDGri7gt8Cu3C7aZfclSnJn7T2Ex+0C
J2csoKIKyniZ2IHDOq1IOoV+7bOGFGDfSfiI20y+ChQJ6T/PG18WS1TTr+6Ocr73
1dkfgE1MkGZgrJT1GB73YqyoEqfLmjtEUcPxbD8XLehNHiGNMYZWiCGxuwFtgpd/
Xsz6PuV4MZe2AvqimQlgIqg/Fo5dzr7wRXfygFibFNwAZEmETIDdbkSETPGcoo1O
PEPAjVc3a01CVcQQybTWU6n8FvkeqIT/V0aeBfs1SygVD3XyFajPnBuHiTcVcj7X
fUX4/s9PxANanXn3tpeF9kQPA1UQEu16SttpWk3dgIWIdXgKKwZY0SVxU4JLQ/6D
rgsWqc3Pr03p//E8QbIyhrmYvybQZTOb9ssdESaZPQ64hlK+Rro04WkraE9t8hz7
tlrmRobuwqtqCy7l6B+6JZ9jaYRupcKM8Uv68eQEhdVEsg56mF7SYsEp04D0cnlm
h8Lg+AIg7gn9Y+lUopoZ55rSXU09+guiW6aLgivD4gE3HCZZCPEn883LoVOV8yGQ
wQNxw5Im5YyaC5k+/dp80dzHoSz1p5NCeYORmSJvSSFgDwVLSl8O/pdt0Vwj5C6A
NF7FeFEEQSs+vAYTjHb/7Qf3W7swGFdhdn0uN8YHT09f2tS+XigDKVO9k8frnWaJ
5pPXDqcxSrN2f4DVp6yqrCTqYPcPlooYretJgDcFAjsFKUOp8M+a9EHulTyErnrq
w6BwdwOXphWrmWBZiohVkMoJ8ej5cOWYYBj65IMGVWE9GkwNpyUkJ3HOesIP/Iud
sa+W+LLJbjXQacpu5MnGdkd2JSMJQUbPJdqMFIZgdH9aF5lbnrtigKWDp+rg1/nk
Kzjg5+5Di2OMnqAQO6/3CkkGJQC2BBQ9+Ada9SbEKJ0ZBbXxMIiwubGQNHgf2pKC
d46awJEQq3ZBYCGHsnM1Lk0LFt/7xVj5/Cl01OhftBi21OjJCNv4Uz8EertZ1JE2
yuYZfB4F80khgtiEkoAPD44iQnEq25hpCHRc1WvKc2Woby9J7lYUq2clhr9DwHec
IS6QkNN6BvJ9zCEFQP6I1i3zLyb90h10Pr7v6s0MuYlRSbUbBgS8mH7g2x9IYrjE
MucXGgUiCkxfhbHq9gbW4r/B96QysND1+s57BRM7WNinR8UqryLsXEt4lnZ32lK1
tKwBcSK8rGGvweq07UXr79xiSxEN7n2m96Qnqz6908MTjpeWXM1dbzw/LEwQSkY7
Kg/CHJ1cl9S7e2rWSOgmEHEjfSvH/OGkyKaZyiFdmrPN/8rg61+ByU/3ijZI01Ek
M95MFWvwG5NnD7+BsLK+3iDGbXT3jk2W47bCy27ui7Q4X7Ec3eOw9ytHXVM0Lvn3
+vsgvs4X1HnuqC5iX155ziAJNDh9XEsV/wJj7EyT7Jy412s9bROdOBKltPczCWUU
IR+Ig6P/k7UeqPCmVUqKXayyVezNie+AexgBzvpOURLmDUxk2+FSNc0ckevLW23M
qXl+AoG39q8wdSF3jXmtWQ9MDBFbSAwXefWiYoFVNIfxnBiTQjd8YUxA5VZRKJGt
fI0mq0MvaSEqh4V9Mq+SRGu1DiwZC0NyAnqGA560NwUi7gg/P5z9j3Rj9D8JDazK
fdaPrlecqsxW1B4wzmRBOLJczcoRb0RVIYHI65Oary49vTaoQ4jHW3h7PEU8unHS
lNRYKlggpVtjHGgP84qs8CdpStA9Pmn3QV524AqTFA8u/uOZGe3SxjdaEqV6Xngf
z43oAYVjmNSv1dyi4lXP/J9fcnDu93kjAVhXfgJsAgOEKdu1bBGEC/yL10I6Wc7A
nfpd8iVjnCopo/rc+W9SqLly4HhJ97bu852pr1sykSP2SzWG5exZwJ40obIJTjnK
gL4smDYotT3mFwJNWK1mXCsemSlUdts4n79HKSvANnf8svVYW5PrrAXrU3ti868W
wH2lkVOdgYDbCoZblAJfpOHI2zzGt9LMrc5QolDqH6wihPMBaBEUSeZEqeJUBgmD
jp7dHVTN9yQg0MsnTCXWrEc8FhWlrpDspN9m9SYvksIJhu5SoRa02zRleemvCq4D
j77Aeed+sKnM7OAHVuim5kADmx2N4ra4wsKi+lHGliqRpQd1ZDpMvSu+pamhqlVw
dAFaCLiu/Tt9ZXPoIkxlNx3WoojsCEB7UDUroCsBZpqvHCtlMW7l8+9Sdo2PFBss
xDzgJr2Ij4Yx4sXEvF4NccFl6W0KjEChNYh+pxROm3xIWjaLVbLu2dMFe4j7xraN
HFPFjJOjgTY9WpLTWXzY5VxAJ4cq5EhgyG7xdzHBbiIN886FpAemEcSs+FqfMHjm
prSsE2PZYZ0T8nR30Mg614ob3i4vwM/pSPIQr8WIySzSJdHX/bvTA2KN+HYMh4ve
oPmLZTWENn1b2Xpslqru5JC7BHFFuGsTIJJF68NEuZHf78TcHh9XypPlxC34BqAw
4s08ItOxGokSxM3D/ulzp4BLQzDllVsJBaHRc7JcBuLmYs7jd9SnNxeQefc3w2zv
ZQiw7tORFUPW3u0i1NAvvGrVYfBtfQDvlxZT5MCiFoRyc5Zj9LvgwN2qGO0akS1I
iZrpUTkzTOd0YDiAFMhNmDswOqvwl6wI0un55m5ynlXcZj3Al1YPu2BpEWysP9Xp
OMg0bPc2NGJghs1KjL7OZPE1qyAKd+fVlad4sa1Id3oyVbopJSzyJbFyfrmSO2sI
dZ6EHR+9lYsGYkjBhDsEOowjhyI8EytM0l795OaVYg4OhqxkANYdo3Z4JIfSJypY
q3+5VBNWQrrvYQC/bRPp2c2v8XAu4Na+7IcmnF+n2fP2BMl/wT8Nc9napXsReu+d
2xUU8tarXoAknsqw9CzvY/AWSSAKUC4oSFF9bfQtUR2HeVH8SLnIkUep2OEa81AV
9wB4DE2eQqHKG9Zo5A9vjWAT3IOxjaAFyA7+skzECPt2tTa1vPTv1KtODGQ7nCjQ
K8D89ATSNiH+0xCQanKRGfRP/ltWz4k+r0oDFcFYCWkIzdWav8kmNaYCPFtSD2dC
OOf5Ppqjp/PgChMSLtNtNPKnQjKlB4Xr+Oexswjeg3G5kwcPiL5pzLINK/QdQKyD
f5YpbHkLtIXCikmNlQbvBFMp8jwjTdO/zJw/mxVGR45FCZGpLjTnv8IW5S2QVTN2
4S4Wd98urPQKwn4KEU8uUzHlCMthkK93r7pL95IE3jd8JPVZpN1TvU/iMbM8rD9z
zff8UNGhTfpgJQnbX8edaApSWsuVVqMh6Rf606XYwgUjiLm+nqzVs4Ido5Nk+dUB
HKQbrTDeQDg26+FtCQK4BGKQ3TWdd7lJGiiQdhAgty7ou77xqQ4MTkPZ0hN/TWIZ
su8g6TdcIHmwgVEjYrsidNhvQ6rcmVbrdUmZDFcCVJioqifQwDur+QZSA/pej73Y
oWFUmJ9r4IUgA8Q1gRMQ9WHnzWiewYT5gpn50zwdqvrAJkF8Jp+nlt961jDx1p17
VaWX7j9ZgYfcLAISpkhz2LclF6QRq0xaxkFBguknb4Sq6zW1CWslRT4smCxyONS8
gIoA0/iyU+2pMk041f91Sk9ETnDHjNhjm0jzdWDqYo9iz4e9rP0/82c30CeBunBM
rhLYm4whxRasOMsVwww64xUjyc4ulCshZO5PZvzh906UKlY/DXRFMJ7mJlavnuU6
7ON0bMvc4uNcquklx8kbNRPwL62xsmIQ7eY/gEUQhBZJVFEqUpa2pG5MMtldO/il
KcQf/XWa94IOo1YgDojSjGArb0rmCiV9izh9eCyJXs5kzTMqMVk87J3fbMydXaLp
yJohUb4SUAY7/G+/eVDIOu1uWS25MaSoA0mNjrgjdePwSXbssr6zd2UHzWUoWPTu
/gv2Db4dB8KxYxK2v+mvjR3s7t+sZvpJAtsvF47Ra2+41RKZW17fakFK/mnju4eu
DS85oVkL/vp+dxNZSd8iABc8y43ZxMFo5wy4ustQ/15QDkfbLxN1eYqQSpR0++bU
7TJqqY10FRdLGW7ZeriFsO2UmmaGxPw9LLJJop+kp3DmQqdcnVkN+IrZCgNgvwd6
RKz2A17GTtl4LZPQ9Lh6GkqvwHlHPn6waiB8Ui3XnEMBO8z6avSuRkwYtwvwXltO
7q3J1zTIpPzGY1eGhvioZ1l2IJBPihBmRxLCNNRr+sbZaIr+3SFt9b9pRf6RX3Zu
O0aR9NhFmq2tgvcwzUYYjN7M+MQ5g+Uhf6fKWwOKRfS28CpqHzCCM3K+1vd2NySd
reXtl5ab/VG/HmtMYX192+u8Jj+InkbVI4BT71QwZD2lqxR6C5ex4TwXNFpIKZjZ
5OsosD+afEcpoBQpuO1m+1daUwSI27sxLNdS6YdBIq5tvURHE1UN1DxbsOm0eB8n
iHV2y36GUxoZsvSOUUOTAzIY/R1qpclpyKt3d/XhWEcQ47rPag+C8K6wOZMFtdFS
QmpYomVg6QCzZCQutgNJmLXq7H2UeBBBSG5ffypePE41ci9DBzkfKZicf+fz+eXK
MVrhLXQpuVY15rweCCTTyvnKd8hyCGiA6mkyqcemk9Eoym8/9ICI6R+InErFszet
EokdZbIbU0tDjHLLR47dHy8EAq6XnZudrkZ/dW+k93wSGtzbDxMaiBJtj6gmMG5v
sDhfBdNC0RRSPqxr4F4/gf8hj8ny/Aci+T5aultM4wnAEkrfaLYE3HbWRqnFx6t5
FjzK+Pmuweh9k3myX67fF3xYCBpFEy55yM1DH2nek85XEk3+OPVvpVYquaVs4XXz
7gHZVVzRAONT1tJkDrjVYd6OX6UggyKEMDz4PyppckkbTRth9JI0Ri/RNZZGlJW7
Y9FywP0HYsjhH4xY8qOGk7uqc/P+LDxwp6JilI+ftu3kFUgS9aPYq8a/dZSacctx
VXV1wzXRKou4yAIUa+LooXBJLQNmzp7plb1hBfyr5CraPXNpjtmbs79hY8bg4ldk
YC4Bw409gWsiGuYBE8b4ZetQrghiWIjFdOc8nO9usHvkoqgL721YbedhfqUN6xer
LqiimkPLjMGnggQep7NMIjGpGvkVQQ4IG21oGXHnGT317MxNbQjwL/T6H7RlnkN/
kV4oQQzpIDDM0KqS5F5xs1MJoif24qCwwS5RP7rx7qoSMvrNQBW4G3o0xH9dABxN
Q8d8q4jOZ/nfwQynyDjql68JngWQjTwn7yFneVUTJ1/T7ZUjtNqh+LK/9g9Qq8X4
ze/sggIHNwbcnZ4tLSeApbiB5Yj4yi3HUJl1lLAauMOR8gaNr22Ya7j4ySe7xavl
uG7QhWCtvtdoh8BG5osXnOf9APSO+AAwXVsWIMvAs8T6YSsxddYvFOWV6sarZ1Kg
QMFkoWHwpg/scuC/iC8nH3ErEqW5Fa0gl2rALBwpclOfGugY7zHjUoVgOVDawL8v
HUgc2JwOozs6x7j3nR6vuVRp6QW+rla82Baai8qQvhZEbmGOxWZLP2H5PQ7QRg6p
KH2iZIHJ8xK3do8ef8BXbMtAeW7DDs655+o8vm5NBmNpLqx4MiprSJMFw86YMVfC
v1mCOJE5j8RnvU5PF6wH6WlUtzqAGLbfxPx6lygGcjwBTh1swPygVISCINF6xXAt
2IdiedTMVKQfxXXVuz5Kc7DRkISntMn8Dgtvu2or5DIyVpK42SiYg+r+5PBpvEsF
VQtPrFWGVVjcL/bhWgrnMsnlihjqM832o5bNgyPX+kaf4/BMywbC8pwtTDPiAx6I
wM3HubhqtLX2dsMHfQLYNuXhMr0mKmqVbsnPQuuXssSIbVAGZSQErf40tnzDd2LN
R3TdowiHzmDvwSvRyyr6I2OkSLRCFC5/iHnwauofUI8M3CEYNCIOvZFcRjfr0wvd
Qx7Dp73WFRBJPKbKiGJihIzZaDqMyLyNE4uER0RyER4fHZn8xfjUuqMTk1uekcUb
qy7LgHNVtCWzmm8YTliVYK+QLxlHofa5yHtgq9/KSwR650oiioyCJAKAmOMxUX4L
Yx/R4pVbCu8CGNVoWP8hGFPM/Yj5Bl1BoEr/KGWkJrsFUEbEIlzsdBtytgoofLrS
T2DLLQA5YVpMnTMs/SkNR6qjdNhm1yFcBlydTgWFfsrpOsmWLw1UgIWIBH9L2WVh
GRYnYL/v+YrOP6TXShSGhJDRqU5fo/rYeioelLHGSEN5lKt/0REsLuw5G0MnfK9y
xLip/bDmaK+586oFrDLgzzyMXKxSHkRjtQ39+qSBGMDdNi305A3aekTWhRQ3/jSM
D37l3EtGzq+SjMCtDDSpjttm+LW+I7bfUI5FrUZJsxoo2/n9P3lQexRhDJcjdlBr
Y15mos5i18TbVLwAfAi2fv+fNsphF+1ocfWlX5KaoL+FEFqgruUuE4KlFFP9YsOO
Bxr0SND70q4bFmohS2QSfEv+RiIYDLym4B5jYoHEgbz3ZwFiHMUYpBBKvuUegpuS
7bGXOdIFQxBmIszDCNUgyVKKBa22ZUN1t5B3upgQFC06k9WN7S7I0GrBPbGXm/vM
6IhPcEN/nkRt1lzzhggpP/HfEidSU12nMMEpTZxmYVzxZzkgZxiq7cwTwyaADBIn
bL/qG8cRwkPU34BsAfeYxS+ZRRFu93tOu9DhRtxzE8yQfHRM0fIAjfF0MPm3mo7E
fpEMifiYTRYZ3tPNu+q0rrDpezb4nW5PrIrl6KInrLKw8qTyOW1ZvtpZvGCjhLZA
4ttBZpUulhmAzo2FxXGsHH3Wt8BNSSiDmPJgEnwjxCESnEeBaJn+Nt0+aYUjLZ3i
E56ruMjrBc5fzGXE9y1/unwPlAuhAPLdQQWNmY5ccjHz6/ZJpQkWXzzepSKm6Upa
xC5xiy7x1j7HT5pslpziz/T/TUEAiQCAZSivdonaRGKcXyW3quIbvmgkfewOkP0a
oytnrqWemHeEsHpG/N15awNsaxyMK9sK6uopuYW9Z142fk97IqXu4tGIRjrJhOpM
v1xp1Xri2x56Gsmx6lu4mrdux4ER7a0J4LN0LQ1mfcaBm1Qzwxp607HC7C5CuDyE
vYjpQ95mdfX6NW3P1d4Jgz/FldYcLhgiFZQ1cGv7cNiBPXLMXM/sYqiiLbD+HM4P
2uLOidQ5MVz1wzObiuHDrNJ28HzdLpvJg9NTmzDWoxYxarab4hBaS7v0iUCmvtyu
o3mQWUbGj8s02ZtA2ETIcAFHk/xct0znOLcJxFZTn1GnwLraeBklx4ln94yJTpnn
htV/jgEhANQqAPaDZoiXyPxQ/0iKMNRqKwqugvmdjCF13Xk4B/FUEgEalJlGwttR
ECeiaoPFvsrsI2Ko4yslMPFoBvKjsiyJJ/oCkPUQYR9UwaAvnXlIYNxexR7LUWqP
gRIR3ZG3DNtnasPCbq56rWS001n8uI5OlVrj0QYbCMnlj9CO2+NQWEPAytLy+jMW
ZByFjcOgij+mIih1JpVc6P8wMa9/GliqdceHoqW8mbLCwL5qiFszYXoQ2BjYJxt0
JMMWIX2Cc7NKdOlVL84CAE6ch9l+G7JF0cMBHOoBeOja4SRqvYGN7NeQkTsSYYCj
FGEN4nMbrpFCY+Cdt7Cnj5moIRPru0YLXy1d5uSu3pq8PtFy9aCENkxti8c9Zj1K
PqUeLmZ8oLjXmFxhW7GJN32cbh59a6vkwqAucbaVG2CWerNI3mSwKGGZ8ByZy2va
An/yL2BgVcEhJ8W5zqwHs8YIzfzaTD4wZXatMeGe1f6m9PuZMBTDKBbwgkgXlMph
doZ75BeeGTvnR/SPhEdhQtEcdEpOZSsP2SddAk9Cus9sIHnkG72rryWoCb9020JJ
ouxZNXWN1E/PB7YujxskPdC5215YX+NREYax0UkBVXFuG4F0nK+kSWDSXgoTz8L7
ie+QoCEv7ahJTikHrEeleHi7D5XFuKaQrT8u0NlstWMK9LDfckR4ycPKDRdbFg4n
MbSwpuLpT74h9YKC2IABV4nJj3W2ljYElyyNr3o5pOQa2ZRkdl/QAQxrIntkdHrJ
k8WPGFP2cJOG8uvPmtk+z0PkS7b71+yfUYzTFownxkpuPEsLeC9MSthlB4Ktmf4H
grt/PvBc6zJ8jU9ibQJGoPgpmM8UBrT8aUWXXgODZ/9ufon731e3xA0RcvRHJaN8
HSd5NCRVw4HULOCXkBSnuDMhQUyxcdHFVQKjl37Ly1Sa8pdHB8qAAG7kXlgjtoy9
060uegCVSxEO7woeXiEwF80xRuwpQgp9/F/YmA/utf0nGaKSsRGQACnSXWQs1LAL
sp5Wl2JFIveYianYWmsoM2SArelhfHOKQSn1FMd9kjUGCDAFbtryk+Bcx7tmbVB6
olPvJ7fJh57h11REdDuBbme0Fq8kXk0oxtjyyq8HucgHFarCL++1etKn209XuJld
s7qVsD+Z1tJOyUT/PWb97tdUxTvNVCQsn/Lg3Ixo5+0xeF6jLbuZwmE4cwh80pJf
zBI3+FsuVz5O/VQMsp0++ClbvJZ0CfWG7YDwFUfhUvMBLN246HaG7hMlvxM+BtGL
o1GggS56FBuUN0BasO9We5Ex17DtDriGQ7+4R57uUg0SOco4VrDScFJEwN+TY7WJ
MYL4XNREj5B8YsPcfbOW4SYLHgqfJnB2yot9vBcQMkkel19vFwXklUJMDQO7z/g8
OUg39nuIDGMlrPm1WZHS5yAH0necHq7g2I8Wm2PbnJvXpyMKrQygsANastERG1U0
S/vaBKirFrlJfU/vZ/7nhBKsq/SE9QKzL+Q/PbQgP2hYNfP/UCXfWIY5S66XNxCY
HKLEbsjQkc5F5RoP3nLOsAoFeOoGwMmb6+Y+xdFZNuljqAlds0oW/z1LraQJMx1J
5aq3NQWvkbsyg9Hy1l9eEZJ0AEB2CVqpMxYzDZSztV5s0YMFEel7T4Zen+oXbA7+
zRMZhbOTB9HLzUewKlf70Ky03RGDAX+IeP3VmoPQYjKUoGnGotHj9/aYxwu/a16C
rgWBA98GNsHrxQx3uAifp7ryS2asr4QfDOgDtI/r8xT3t6UMehnFVBWLe2VrTRuf
IPxNHfnovBQcoaledUb4kK9+IxQRf4arUaNI0BC9WTIE/WXJO0AlET774WY8YWST
1hoKCo2eq0Z395k4wdbynDYncz5GqVnG33pGfQFoaQ2qnJKQwQLDnanCksBb90Vo
ibi+ECvA8F2//FTSGGiOeZotQjsej+jrp42YHFa8DJAhMpVp8kB6cjKBWCbV3vhL
Ea5B4BOyU6Y+pwzTec2i7wkoHX7YR0X21yA6mT93QhvuTdYLNZXXeZov7y9heSBj
/g7JhJ0QYVNzR5YGMnPmJjjzqpwrtXRzvUrzWT6n6GFlXrjf7jsb+9DwgD8tH9cY
EOV8R4Cyw/uGGwV7Y5oysdTMUz0H5lFeo6Ftn+1tKohIwvLqL0jqX2A35JHUu55K
laGbK4NB94ulBg2BEzn9+NjU4Z4uctRBs9u7EXGFhZ3OFpY6rWQ5FCII/53j2Czr
98mjEyuiIuGpT5U1AojtDk9KKb1JnVLoGFAGRPW966mQm7kpMggY51EoyfGWk7Mt
zAS1jeXFAB1S1uj6Y/tEXsvv9+jRj1ZxqkKbVxSfM2vFQ392y7CuVPViF8nltRol
bABxSXKXlyLo9bWjNm426T0OZg5SfckraJcbyaXb5Vnpqvocd9nkptJxE5LRIHkz
`pragma protect end_protected
