// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:17 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JIWEyE6kOw0hiBfGnHuDeYwBIS8qlDuhlIsVBqgEglNW5mrt6vWxtDW+EJtXILSz
/RbiyiJ7VfEPMpCw+1bWRHJ5SClaVJ+wfSDihZK+1LGFqUoDAVVP0F9/smWS/83k
7rC+EuRNMwnMqVgp0GaR7W5WyBQPuM3Jb/mGPtzieEA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 58768)
sLjamwWMUxXtwcjygoIP/4oHoUcMdYSLvaQ57vVHPQoffHJXkwpD2d6aVFZ7Gb9S
rfgAgG8QXpOHtyMyO+oEg9OLZ79KWdI7Fe8925YiyxYakftJDxVhyKP+XeNz6g/G
34ZAKZ2wdqvJ3O+vJJ1h+TXan+so0pbQ2bG1TgaotnHL5cN5Ptljr0/m6ehhgXqf
Gg9yVpKIVaMeamExWdT1DfoTXsZtsjNl95hQynMroqnRfKILWlpCdiaO2hTjOqxO
Z++7QBhxXAKy4gu3bGz8djZc+lHl7ZWhqla81DJHmqWYv5J//DXDoDw1mxfyYETm
dPgky6LT7fmFfxwGyEg8PJtSJNWuWNf9SkAso39soYqL41fFCwrstODp4nhIAvHS
g2uo77ufTMxSYrg5ZsLo6Hg8PXgSJXK4y489ArHjBPnKD7ZZ8mv4HSRTRIuJQYVb
aLhBJpW8fgZDKucgmndJ2fTjkb+5oFGsNRimRqwbfce8fYzXfsE2OL8KT+BVtd/1
yvaV9IvjQCpB7GhwBDxc878irr0KO1TfYZ7L1l95S/lTyZbTxwJbxe42+rQYKALe
scvq0gK9miUn4dWA9+yV16oE+QrUnDTFtaNltigyNrVrCv/ZJ09t6Nscst6w5zC+
tLXML3Z+zhsDXIDFsWjVLPQ55aguqmS2iAXJLzfX3TSKCCO16sj3SpxS4ICvTEpL
cyu8FKQTL33/K5lPB0ttcBM/c7SLyeOvsPTj1NobsRiwOptFmViXbI4YZTEd1b0J
uIVQaSAqbMJMdEnd3rPLp9BV5wcO0WMTbJtgwr8+BTxDHFhIVOduvTtZhpYYKBY3
kO8q8/uiQbgWvUb3GL2GD2TeqnFSCQgwFvvMQh0bDrah8u/15Ta9iR7ylLdZ5rt2
JGrngaX9gG1opXV0l/WMiWr9a5LoUwpZgeplR/9hCs/g9mTisRK5s3Z/a7DXYTgS
/zYJ2+LG2KtLnGsUN+2M0JUuIT3YEUoUSdu4mkE5zMlKI8LRhOvR8ORii0W805+I
x4k3FmGabUyOs5KtfKATEwwf6LXJlykjw2aG/NeVsxqHt1dD59YrxKcNEj9QSI8z
PCD9nzUTpnyCo2Cmm3mVRxjmj/o32/28v7pmMfel/6wTmEOD8umvcWZUT2bR5jiU
xZVddyg/grw2Nj0ibLJoitGV7HXrQNxIJyV0L4Dgf/xSr0z2dRHt5g9sPG+I1j/g
GKXhr8qDdZ7UKsuE4ZUPR7U768rI+kPpwk32FlwvxvqgWs4l8S/jF5nPjnZIkRxC
KHcYqWo2gG8voB5bfJLzzbdbNA05ETfWzWMXckRm6n83CWqfoTuYyfTzMgjR0W5u
CMLnZApaetkaUxYHixfzU6Thys2G4+CqYcP+1FL1K9nUVkIYBOTSN0ja0YIcMC1O
CTC5mwyK7V26vfrkrIGIL/kuwcc95eTF9Fj9UklzbZPbE8w2l1E000/zpBYlYLeq
Zqbk5I6p6IM6ecd9KPv1D4h5pCzGmxvox2INT+OMeSBKJHFCfZGXpj5L9ubm9+9s
Zy9QK9XFHmt5JfUGqjxWplxHlRZqpPCwgDedVFZEnJFAu8Ti9WRIdjuo5UixKw6E
5EtCG1ZY0gduPWFESQgbSheOLTlNEU8pXS78t5qh3vY70MmzeCEMogcWLO/828ka
5tW4VxjcMd0Deni45h+e3eRIlgyfQ1CJRXDIf0WYOAKdA18LFpfzyJDX3vD/KFDr
CwKKeCYDLytbTDO0r8Zk77DV2bIL16SOo7P1eZanPOiDT4NswiUyl7yLxLIGQSGN
Dh6DlUR8xU5yIsAL9Akk59hNRA8LR6CETgTpmCkzRXQ7HBPtjpyL+lT/K7jAsqLj
LfP6U7FVQl6mORRUayqDd2kQIcdWSdDpilOHA8kVU5vJpBLU0x2x0UdQaAIcmd7m
P2D9NNgj+c8Cf3zQ50UMN3I8jX066HfzLZLzy3ThyqjE9dvFRkeyWGGNJpoEON69
P+SgLBpdLLa/h8u45Aer869LwiOLRXhff06VDCafabEOV1S7Ohhdqa9IwKSfiXMg
0E7xq2kCBAG2q2EbyISu3e4arpNOd9xO2/AYza3w1NdCUvSExOW8nm4UJ3Mkj/q3
WV/NImezKQd0x39AW7WDzM79ZD+aC5DgHMW9zPKQRzIbpQEgN3ab9fD0MwO6nvn/
vMaHX9dYtI22OdxldMlvLee5Z90lvNruflCxHrNa0e8MsiLrQFHR38rcwFp6N98D
onLzyOBWzbcWeqkAzYxPDI4Ls/HHKczqyJx5MYjppv1y8rC2pkwGh/H+mI8i2t+5
gl1kw/hXWB380XmOBE3UEHsgkxE1Evxw4FIklBg6Idt4T2pgCl4F1+jGwc1uxkxE
iTn/NGMq5QBEc1RjJS0X3znJq7AoJUY9Lf+/jExAq3afc/Baz/HPZ4ZLjKYrg2EH
jJc0ZGKmXMNvlOnU/Wpty05ZRlGNKQDbs61+Bf5/jU1CThaxQRsQzKvbIvsvF3id
kk4iq2EhDqS+jaMVDyJhHNFiv65L3WYt1Qy9FSfvxqM2SmeR/ZQbdKGPfXtrlXGR
PcU6ubIFhwhZDxdAedtFPrD/wvaj1flItHAaPaAcQJE2swiGfm0P0d14TRIfDdGd
2ZL8yjfpDf7jkmtQuf1IlIf5nOO28hQURmHvsbzEpjfyrVTFDDXFpq0LBiKH6gQ7
bcFLTdNKh5BjFZiWlReIm0DpriHMfpt9aeZ0H62JxXVHkGG7OqKbd2E/bcqlC5PN
NKSVwpVuXMExajQIJUtkpwOfEQPIyf+ZANY9jSsv1ASRGQx7qAIOoZLM4W57dnWg
xbKufkAJQHRc9jOXiSqHqsVUyrUOYHe0DeUmTDJzcC9rL7v9N+lU3hJfVco5tPWR
wOCGCC58QTVEmnimDAQa8/j91GfNQh60Tm9M4eutCx+EciG7e1pW4I9B+Afrt++k
WJzD4KehqYSwJcmNhmYJ/rTIce8c2FWGm0G12NjgF8ja1q45evatLIXkGWVN9mOc
gztyjhbMYIsTJW2uDNU1KANobicCMUgPqTxX9PHa2lrDXHHAaAjDZYEVv5iJXXb7
EBhTP4pQogaV8U0TDnEvJZrqa/LTzKYVetLBfuooc30bv2buIBJZ9l/HJPt8ib8h
F1YrXev49IsoFx2yBOmdajCVcxfwaFS0j5jB20JM1hxJOm6UD0e5valBcK5okATw
41e0r15rIZDpr1OKEJx4oU9+qHWbCrDeEMZBYZfmoG5ZrMYgU/XAYaGhXA2Xo483
8/fp9LJGArj0bZZV8hQeaofWmaNTBANoEr0zTGYnGNhr1mzYdV9b5gE/2nFGLhTY
42qAnuqYcGLrjeFyxJvXh8RL9s8C3nW59GOgWN7wVTWx9+AMDLqRblLcvJeMJBa7
9WhQ9N4ZszoYi1Xk0OPH5JoxgSZbG+9lPbrYlHxPL4VXz2AbLLMwZn28KOAIJviB
hBC23I1c99DyLcKXE64R2TeE5ypPVHxV9Qsl43ed7tyfbqjhzmF0NTrQPwQdpw9s
8IQWNGv7ugnreZzWZEJn+JekYmwhG3tGVU+Ip0nNDwmDoN97nXfMYGTiXWuA64vJ
L15fkbVOGPrm1ltCfPa+q0dnvisxvVACtSh1PY8YwIhGOQZg8EOvztVNo3orO+is
FNBd0Uq8XqNnxJmCTZDihLpAiBfT+pAD6GzUaMyH9nefZ4hB6zeWe49U2pPTnaXY
qVFIdhEmPfzUjXjWPyGzR4nzcSIoYncVvc7GvcbDLm1wYsXsCrAAoffvj5wWc+Mm
tpYZn+uPlcF50/i2WgwOnoD9GbH/BKto8H2AOC5AtomK6+6Ai8bYZsLBTBoAQE2r
U0xfbr9F8haI1ywC232+jXs+eOgNS1WWs3kWXzK/JeJQXENjSGoCxRiPH6+/k6+Z
+sp8rQw2FAExhLKkd9Tpgg0kZC+Va4j7fGo3U0SV1oyFvqFXv2idYcdqNDfTbsgQ
k/haM6RNmzf+XKb1mvBG/pn3Xsx0D5QVV74NAJlT6X061WQRS+wipH3L1ajK9MJU
rcynyyknAaNxVd4IIO08uJkTV8IXnUd1DuATYb8pp0G3ttd+ch7pCzJ2PfVV1d4R
Jnfdjv5bDL1FYUvRgZdXYVRHqb+2Al4FUbawP8fhQi9W2YsUj2rLmPKyMbPdd47B
UV0cOBysg5SYZ/iNv3jZ0GaFYDdeioz5QDhcNCrnza7MSJt/GdCUkvLvkAmozDKt
U2ugHTBCFGyGGz0MWbJ156gY8ROYz8Uusij8bHK3YRZoSJZ+2jaoGOsOrciE/5De
xKg1Rmd8gjnxj915xcxVm2UlDTgU/UW6omZL2aFCaz5IwNxX1lYbUPCAwJnQKAxd
Zb7ulGHcZQpGZenKgzz7eFQxZDrm/k/sSOsTY1HdxqphmhF07/gWz0dxU/ZIIdnW
ApphcIa8TmAZg4UNTvvPy86w1i6E9sQ2ERNdzwvzYB1yT9PmggLga1gmxr0H77Cn
msatyop2IaKPd5YcP0xlTo6jyZ/w1gEhBLcvFgeM2MSeCfZBVbayiwLigRCp0lbK
T3jLcoZttSzuvhsmhR3SXqcQ41fQvYPplIIJmVA/OEFAazcOZDOoQ4E5UCQdIOe7
dg9REPaS0H4NIgUdSe93ZCX/9ZfL/N7IieOhyuIsWjm7qFkdZFM9ateu886RyRov
RbJNv87yWZ03ZOz1Kzp9R2A6vRjgZctWcUUiaSWHeDuI4jb/kJ3b/Dje6mvQNylK
R0QDnjBE+zT/hUi2n0nk8ndQKWMXIr1Ltp/b7hg7YtpphVyFPvxFZEnbcDgOfotq
iyxENrKvdrTK2eQi2tTQd7Ix6MLFEyJXDEEyuLn9K4BUwnQH5cSgUyqqWkFH7sfO
s46oDRNNtWKYg0ZAxsjecUOx5DwAjCBKE24pGqNtt/Ez+wxozstQZdAEANDgCYBk
EeqVwSS5TpiluvO7tzSwe4axxzS34sRVuqGPAAtotktJdh9pIPIASXBsQZik7VBK
zZ4UdrZ7HpiSOLHBuk58x5Vxa96WwlnGBstjB4QxrAaZc9P9xjidE++LD7lfQ6an
XQuPHquq1BsvUlScoRV2tkgNYJVvQfbgH2K5Hr6CZvQTjstNaY+IqNGakUgU+f0h
iryLiMIDyUK1JITY2lonsewg6Q8CXHHL6DOuXf4uW3OX8l6wscisG+gmSte4yOUR
bhPF32RjGLIewfmz4qoxeo/eZOBKyO+GUcuo5mdNwO+dEtPoihHMU36//zZ/SGBT
63qN1dFYhOdLE1ew1/ftNwf26WveYn2ySCoD8ZebbsYoOif/dOB6HYD2JPY4bQEf
Gh4YRBlCnUBFK3j9bdGen8rIVWy4sgrr5JqmKN4hYfTRBl0QwRSbeJsBlX5fVq0l
60f7HDGcrr1UX2zE4os4w0KHpbhOl5/G39qjl2C/r0UquoZi3ji3rMDGZX+rERN0
+YOdsKkVJeeCwm6Um2VVhlYI3Ghwlkr2Ebvl0DG6AjDvc8aYkKmnCIrWfcsZAY/y
ytXTD6u5OyGEJbhSWDbjXItwT8XhozUfwAa/sOrX9wmNPobpSpDffi7q28Fly/tr
V/7igSXi38vz2Q7St8GM0qrU6DyFxQusPnN/9cLyLaFagGZLrh8WLxT32QOctUl+
JlfVMTdozt2XoLVRsYWcuhUy28D9ck/ZyVuGy4tne6cam1dYG6D//aofQTzw3xvQ
tKvutvoBklzlagudPbTbkga3LSKq9/+ADbIs90OIpx0OYqmMRD14AbX8ehlQD3zG
rdlrPffNA4LjFHywJTOkmfi+gtMPLy8DEN2mTdLtAgAJDZ+cpqYxcggL6A3PEqP6
QJ8xZc5r5+p2Xo1rcMkW9kb9X+PcAPO2tUz2ehtxEvR0GBeEcn+ac5ZVRmVMHEan
0mfitG7i/vpFLDAGpt+JFayPu6HrwLpyvtJP3/2u8xdNMnQwIZt6u84/uu7stSjw
5UBHqli+Vwr7PXIU0xnYfAYVEB5GjtzsAIRV/5eDWuZ1CSaSa3qzf/U6oFlD17+4
dEKllqZUsF6EHT3Yzlv3VxsIK3LIuUiz41wiTEravxWexQylS3uIshdWw4BjDLyt
JD8IoEpFWCbWRgNCKr/iDG9XcHClogWL5Yd6iEFup61vYg6bP/vORm7RJUF77Fvy
QseHDCRps6WMqIydaZJepUkyEwB7pUW1S+16XPcbvY4t7IDtaR7TVIOWc8qH6Izq
YL7dOVdUKszF7z+S7QtyEtYwE+ts/1qUMrGtMkKANbK/ieCHCx3ViIq4sVup6Erw
XSS4Ur7r/KyDgOHKvJk6f2lovTnusa7CGfL0O5ahId3lME9q3uewydrfv0/hCVPf
B7wtRbPEx8HErtLYt6+l0BcxXdf3/Y/+krMdbcs5hvAv54joP54cHvzD/ojfx87e
AdY1neeiQNyti8uQp3nORHY8htsObG4cpM60OAyX0IwQXcq8/KXzi9JsMKShNmKF
Z5Qm2XX5DNddDMgrKR2LH0Dkx+yvnwpm2pCEhtk3G5WRaJzXhHK3X/oMmbtthE2C
yOmXV01imyJRNlPf3NlVvQlcSqT95f46MI80klQlUIIKelU2dbJlhv9NnrDsRmZy
KJjW5rzttaDDpBIqcCtB9zvP/tpTgljEuj6wDxdzstKXUuGFWom59ra1Zk6ClWN7
b1R8f/0rabLPCSmebVcQem2le9b0hfGnhvC4ERvAFD9Wyps8C7SFgY8dXl394PB5
FZ2WXn7mCjeE6A7AnbieWx/CBp+0kn2CzI5lkFNGh2BzhwVZWBsHfnwLvTtd2aY/
//rW3f7/z5vFzUg8FAGO533/yxYb3tP/VVhR29HpoqNiPeiuTlNuxdvFxVJi/78h
gFv6Nr8KbRd9uZiBFsIaK3kUt3Gui2Ic3QLAjuhQ5EJ0WrB06W2ylLlxNn72IeH/
ToCHkxDKqwnpZjH9JWQFbCyWsF6MBh2h2HDaEwVKWfRcItMg4xC4nrFFgqNFw//Q
nosqlqUz9pyGs1idiXbJECRd5tVA6g6ma3D0nrzeuFF69Ud/4y6aTsLnWFoUM0Br
lVIR29P1HUqkm1gVoN9g3ya+Uy3LhlUz04ljnhjbX8gxEGkcW1abkM0U4xFX1k6Q
gqWuDNgCD9dJoLroj4YdtWTPZRYas2hBp3DdzDFO/rkou9umEpJMlwY3Tcr4lMRP
7NmLQqIVZSMIpfk8UwDG/IfCByi2o5r9Acq3w8KIO4HSndvfGOevS57Aehdkcka7
pRhYAOd3GQ19hiqT0/aenzHB8FJRbNTQnAwdhfL4Fd4RKGBfgeD1DigcU8/T7bYd
u4bkcueC6nSBP49OzJtxo/nScYD1MLMgvsGRUCMtTMUxISGxA0cP5VzaYaIXLfKC
kYupK0pxWfr0Zl6+BASThDaUBHJhxzl9pxDs/a9OoBYTZC1oGUPKA7jxZV7UcZoE
8DQ/VPrs35sIgBww4px34xCosvAlQwnWUXcZAhEftVvxCeye8ZT+57HHEI1EFKWJ
9Vvh9nTO2MvLGYfW4iDdEXP3z8UPuDNOqZ8ggzajdnhBDK+k7PnGMJEdTNhkMws5
TcbAOpsvzejd3VVNJfs/O7RChZ/GnBAA3e6zxZaR9Pdx+Mqd2TLzp/7/PaD7Pi/z
JRCxcwOSemC7nIZ5tJNq7VZvum2F+v8gUyvmGSTNO9W5kwCBq3kQnRti9MpyULeG
+wSXXXf8PZP8Hqjh2feT94Csgq7qAa7KFDSBxWpJlZiU9WGGatzRhBn4F4QBPZHD
+9DIUvnT97PKubjm2GuBjEADra03jtGpmfXCV/rO5ccu0+YFyw9XjoxUEGGe3zN5
lpVSiH3nK1re7xzcSTmbakX+7SEsk55T4YJiER02cOzio/eg0gUgX7eDs78F9RNv
pBHtHyGSE0NlNAc7R7ddch+JAZaCrvXLYK12jYoDnDqyzIN6vtHCEDQ2+tIKeLs6
mzbHMrn2EUkIwwqSchH5N2+l0OnSBgKbflz2qbjgH+bUlR3c9YCBh6pDoQpT3y3x
GA/exv4Zria9ZxcucWInMnfVR6ZHQopOfYmlWqnkGnwvVP6YQKjNWQwHqseaxDtV
OnHGOeUgVteg/27Y3Hjzfxzm98wN0YBOYAAptvkD7rU+rFxES93v3F1yAu9a1QF1
GUpkezd6x4KDJXiSGWBrJZjbtogBYpYvcD0wdCH9QQHhbYsfVATwlYP/D1lzEaRu
Gb9WWl6zWc1Dmrv/0LTmr2URpK6RfwIvj5tGu9wZMHG//JKcQ3ABsoeQPzqxN6v/
xG+XoYc/Av3I4bMw3Ai7Wa4yhih6wY/y7+ktxYDgHmGytvbPojuiUqYPsbL7N6ZG
QyFtAq6+1QzbGxoW/4iUWQzEOpM6HRwkCEfDrwz8HAq2C4aLa6JtWK/RsRz1T5NK
HBZJCieCwj6Uffmf0MmhA5OhyJ/bHRfCUZoeXZBjoFhEVABJSbE90RIVhpUQoHW2
Wz+AVkP5jNuD5Td2ptbQNCcLPLlqAn9qnpkMCO+t+HNfdCbucDEROLNYmEvxMD9o
9C33vHvtkeF7Uk05GkymhbojjJHCnW+35I7fuqsf6I0v+1y6OcOLBvEVa+yZ6SFg
+5okaTjFQFz2Otq1NIFy5MOkkQ/gDm9lvrLz6btqA1gC44WqaK1um9xefCgb3sRI
x/w1Tkiy75iSJ1UYoJIo61JuxP/lq5U6NAuJ0SFdaro+rPwEI36bFm2LyQAlyNCk
4Dqt0eHm7ENpXHL/hsLAwF63WPiHj8X+CKkwLcntSfuBJ/ou1I5w5ca3EJmD9jNS
A0lq2osFoXKRAFqXEcTs/wQiWmSPK4olZVZ4pZ+wDttHSjNnZ5HNXoy4tAHEeDW4
HmTuNkDwz23x0Re2qDCh6RQwKaNzGXn4FAutZbPUOBwPIOVIcCmLn6txhMeYs4yR
hWD9gae7E8cXHJshO4uCmI7osRqCuOmf4K6kJ6uzuxv3aMCnGL7skddSoTA5y6vS
wa0wQs2isstgQ3vpyWnVg38p1m/kUWZHC7MMdu7f0JdkI68ROHtRzUmAr6Qg5mzy
5H1SU1RGFI5UsGNCJL60YpSNftP2EaldoeY4/0N9JdW34Vz4rZpWU63nG+3AWzyF
WV8/8zyVw3Uig8+d7Aogz49Ao6F3gAMZFj4D5+fuUfV1inVI9dqJqjnOr/68ic4x
RHyGpf6aynDUtZXP80uViBgFjrRbcYvOD88cmsurvQoZNj+yKtI/SuHmwg/mEvJp
jghP22+TKENAMLAcrVxgPR9fuCHTFsz5EBR+R5jyieEE6v2NRpM4IY1pb2J4WpxH
IT3ab3A0OSOKlu22lYeHtMmFAKQd5jPg7HfAFuVPdIvzbaBDCtB29x8HCplRZPQy
SrIbSOrMZ9uzjIFm2C9NXGon1R9Ie8wKhgGa7UwckftRbxenc902OFdDA1dgwuIR
CE98BPhzclkQd99pERdK8ShADnKbSZq1ToM/G8jJAxdx/kqHCbo+2AXxRCrHoIvK
sFyKYanONfXqPW5JwdUicOiNpobdZFZGvKHAKr/77S2TjrHZiKWHMpLBsRWKepCO
wG0R5gmUUFf7SbV4ximP5B2kMm6feHgWpZ3qDR94clPRvXwIHOWBDTt+W7wbcUrZ
Qbl8AcG5b3G7cpa7mC9H1gb+DBQyCrPJ/7tiWnindcQzC0ti4gIeFUvD5S8IN0Oy
TadaS+5NZU3KtUb2bgrQo8ewNDOtfigJNiXk3U9cz64TLtrSTFQid6Zkc2Uf78QR
nh5TqZEzSoDFDbeJ8HDh64E44VkeFZB5sb6ShLpWmTJl7Dycq5yCx+ogOv+ZVSZq
UVZXO480CcyiqKgMMpRTFSUqNDr9/M+5UOcFwYAKazByqR9iovBfQvdER9Vy5aSN
GHDwA8lmcinG+3bTRwRbz1wEoL0o49VogbePoR//VgpVQT8LpqzAA7t6l/LodFIl
5H2sURracc3G2F67e1xDO7F9mpSk0r2HDmA6lVzceVjxgeIE9klZNDgUeTnQgMyS
KJiRAhzJBO7rnQqJKLVBHLMID91WFOBRVxJkiLWKzDz/1/XsgfKjSQAqi0SaSjop
H6D9G7aijGAMheI0aSJOCBanUgQ8Jcoq8Zb0m2tfk2ObnlOnTnMSehCx3R7UIcS5
xKXPjqJlS55huIvaalQv8QD0PlVu9NUdpg1HQ2K26LHgfPTnNFgpdvS/h8JwwV+5
z2kn8zfZty03Fqvmk/cdw3gsB4iYrpjG4YruQqzyR5iE0lWzuvYyfvv+j7U3i64M
9BULhdYXT6MKfMf09gOixxn9SmEs6Vz7eB5+TL7w31BNVVkKNYiC5ywEBzy4NOyj
KoXLHx3v8qlFmIhnXyyw3EJiIYe5a5crrUPRRexRD1Yq6/ovQV3I2vKnlyTBfMMQ
hb0AzcvTgd4s+AF65rntOBT+TJkindNiop+PlOHFWhDwfped5Z0wZazXmZl3dx64
0htjaWb3UamM5rJBha1XdfTuU8l/kv/oLsJYOX1trUgqD3hEZV47CVsAF8uPHmG9
CgO45ar3B5xGXISY31XueINFWE03aZ//2epqOMC3cOZWSz3fWGnocnOfNROrcjqm
4tooy6sA5O7e2VEFAepkzQOQKr0iJdVoKCn5KqUwTOCrWmw2/115vyxgTS8mu33l
xpyzJrB6Lb2iHp89D/lwCUDLwsyrI2+nx2KT+oLt5lxEDMdHGEhIwNzX8nYc/ZIq
7xC8oxtlEV0vYLBPHBu7Z7T4p5PLBN+IQra+v2K/6ve2UYuWrLtkOOabh93R6zfw
AzQYJjQbHWTI3N7iX/JdP4vf7pJcRrqhc9leal4oXRxfW2MIBAIVPm65vUzHIkqO
AQD8zfyOVDQoJM5zoaVuPYNnq6AAQ+lvhMxMvckx0cLaX5d/3cYcxkEQvNPTW2RY
i/w4VQamcKZteTcJXH5BUzaQ2EccrwYtiw87E9tx9yMSpZ5kGkzPPGob4Y5+rAk5
b7opHrfG1nIOYhsRJB4ynYeKCxD2eYbKIh3DHbzpyntMLg8nilgsR+f0KoFK3u93
+/cAn35xo9YeD6ImnGYmLOXgQJEZx2PzQBxTjoCxV8biWJFC3VOEMMyAboekkl4F
RPlJNG+o6S+stjzyEsSXku+M7Gehd062dJkBFmKBKHhjsYKO8mcvnXIcf4mnZdOc
WljkSdsi/Xyzsn3uX9qADZhhY6hWo8dN3QhWWIJT1tbTVlfOK2Zk/WJ4nzeHfs+y
eHgr8mks8CHgTW1No69NAum63QcrKXt1a3pxoT/o4w0vlerB9b4+IggehsKArD0S
OH9T+jnSMHIbC0CJe4pyDbJ/TPFeJD3zBGTJYI+yiwj3s0hYdgfkSTjV6zeuQCda
LWkr+pIxANqGLVhD1rwMvlaiP9gwbUKJ8509AEU0eUeNlQQ2ndTDtACWQsrQujBh
7hTAwh8ke9Nal7r9okB7QZXdHVPDcL/pwVdcXBRrkwTAFirQaFaDL+UKC5hAorPT
okuOfF1tNwfpRAjNrVGCzinL7wW2tMm8MdTnUXFlQ8TWrmtpsd1Ug5mphAwQIjBc
T3YDkHfRjA9Cv1kuCgaX/XfYHNuJpzMPlYbiZWPmxC+6XS2RvgmiuAP8jLWRzruA
ntdjk02HlF07F0TAQWJq53SFBPGASlZH+hBOFGzGcieiZBNPihfv9cme6uDa9o5z
SJwyydqJps4Wwn/coi5/V2Hom9uBKT3RwkYCVkckUucUY17m+P1qnBNvkzW8lduE
BJJo9ZoOVDV12SQpLj4pn/VfgmKc/zA4UsdlJ0bOEap5mWbCmZ0RGuJzpfhiYgW0
ifN6q/aVUQbEmJumZQdnTCGfSW6SreHfCJVzJKtXHzO4pNM44Jl5gkvMKNDStPZD
1IvSX8goiWhrsVQ19wN2ULE60pYdeR9yqlQVin0crZu453T1yGhvM3CFPSr2g6XQ
PDnsjlPuCW7pLl6wjWumCZw5KER4fb/Z7sWTj/HCt3qEAQoCYp+Dvg0QzDX60Hxs
QMPhZeJAnUKwcqIWHFFDWBt2NRZJOWzFr5IO3tTvK1Ob+dg0BIsJNbxMqrnvfPCk
v76LiM8JtncZEkkH1VPx70HlsoBlTbHP18MM6uDVlc4EUbS1ZjwtSL3+MF956Zaq
syMHJQoNwyw+bLTOfYwmNNwkP33/91CpRcdsYYlZb5Y1EJwvt+0ic1g8DAqQQ16Y
q4o+UnjLEjDUdAlK1xYAFzP0g9cwi94n3+0LNRIXEwOHt+71E9vyyEXd6wGf61Cr
N9xndtbjQqJUzYvKvm/dObF2bhc8KCBmaJ7QMEun55WJSqGESXM9kijgn+e4TIN/
7eAwQaWPE589dwbFcFuopcp8SGaobjdPms24rLcTct7BjG3RTmBGVnkZodKUugxc
Pl8OhMr9Z5yvYYQ9vyC53Xq0FvTpF0lK4XOR18VxmMllH78jqffS0fkf7FhD/PLC
hqnnZR+64B452uPDc0OHc3Y7j31DB7tVJZPELklXKupybVFL8da9TCY66SBdZ2WS
UukfPX/9+8M+no2oym0xaqF5+ElFiFQ5Sos+WyDvF9GC9Q4U1uQUgWVqNU5PBDb+
c5q4UJVfQTdyvDQnKYk9cdZsH5zhSAJcUpEnjCNornkn0j4ClaMOw+7SH+gJdHtO
I6IIHfHFoPVQbf2CZoh6g8wYQxHZ4DobQ6H4VYUZ0pALZTQqhqsPjsUtbfzJ7N+1
qD+yUfW/6YWZQqMdONBQ6Vo5oBIDefq8Tlfcq3kJw/JkIDoius3MSh8tl6z7WsqL
3SqBf28yEVKfaWwFTCU0FWubT7ws3G7HRpf1rE3jdpw5ORr8/uEbRw64EkuyuhAQ
B17XLpq8+FBYTss5JDcGOX24bZNvyGscTpx+2TAqQuidHx+G6JSra1SHwf2M525n
EMM9islmlu4DTdb3YIuRSVRmFxJNFZo5Z42XgLcpb4EEFJge/mAv+62Wp34X+xxy
PnfuoCXMW34Cw4gBM2FkdW44/1yuNqwDkS/oA0Kw5LmPYz1gCV+ntmHrfFCzRP7H
QMJzIwSvJOOXxPTOtxHNhqkIvB1tGjb4Hz6izizGDUy2ffaZLV731VqAp39ovbz8
Wv4K5iOwLTYtWreVloHzRSAIr5Sl9NxFb070a0cTioLK1J6dnsR68xxbJZGqHYqi
R9ARi/GTXaTfPAqgJj3PjEePEkJgRmZStQMwLOUI+lUZw0Yy2DxSLC7vQ8kTlb5+
WngXVpnpTz4b/E9CmidjvQ43KZQgjbT+fmJyHBU+k9PwTvrhSbYqyrnLxBTBYDjH
5gwxV/dLqb1hMYHQ9XlknkRKQflEfy1EY5urCKVNb5nlHnir14aTRzcQKkGZcpsO
aRtio76IqRr1q9Ebn14yeLJrKOm292AxPDjzuYkH5dyjmksQxr8jh1blgGcSQ0uN
EuRSPwametS2VbRcUq5CKziBVwJ8ug1BfsYd2WvCkxQPCMDl/j6XPwl7upUTNLLi
7nwGkIi8Cyv9EAoStGUuxH4ArPlvEkpHRKr7XLzMVsmf7cZAXKvw8MSsf8BDBgAx
vzvjVqUFK7aa69RCmQXkjCU8QXNlBhWDb73s2vcROTYm68xJITKhl+mwXgMC2HmU
aUj6pmdyvT+veaNGjB5HNChbV7jMYPi/EfGkbs5qUaddoDdyVsmpSVipybHKK9hJ
e5zbAozmn3NFfj8/raH73Ti6SNbTP3Cb9CTE2fPhRfDhj7Cwb/HTy0OpuqVvdGi/
30uVPKu1ciaNeUhhai7JCO13YEGvpbMzH0k+4eUAonFBqxKNyL40jSlhGPwwTrwi
evOuk38Dm+v3nMAt8dz471x3R2F0DZHdwy/RWUwbiMLL0E3h6HZAnEyrHCi4G2Az
2X9Ea/tvnLFDkOISTlZ417TqlIIgNtl7zOsa8jk7tMz7bozgT0ERjZFZ/tiu2mwu
TH6hK8CS4UcjtXw9E1nHaFGqCzCkzseHnVI1EmnmdE/EEZ+D5N7xdGmoScAtvzwh
5hPzc4DeGAgPQ4MEDKjEe0JkG1cQlLLwgJT1EfsI/LJwEVcxk1gI+3U9cLxB4HDO
MojGKmAsZFZZvsqXZ5Jh1q8+Z6KdDo+0jw+0IsxZDo1ZEJ3BBCfY4ZnzBMhFj+Fg
bEVnfQDVRv4tUbSabdjBrbC29bZSeVqXEDFLw+a91DFZVnsnl4R/4P9O4Wi18riu
gUbpsvbmys+d+eVn9QsCpVnengeZ0DYZ5x0vVWCu5a5boFvsEXCyvLjg1L8d7f12
P/14by/KPXYWUGyHGQPkWzbg/Cy54dftLtpaapspE4CiaFBhvfWhNuYcLFyP9z8O
Y86IiuV+QMnj6Sg678Vr8V7r+lSFG+TYEXre2D4UOoJil/GJxhSD5iOQNK0THGpG
PpegW8U09de1ZY4/GuQvL8nsQGLmrKsu2AxSucb7UxfFKMv1xQ1snqSy5nEr8Auw
wT1w61O5iGsltfXXz2BxFZ29Y0rNrNeAz8x54W5bf2otp5zkAB7TQuRhBHLPhyvr
fKHBBOkehQH+QWdAXBcy/UsEaUMArQ+FiXcX4T7uVcmN6R875cdIoNjHmq4c5NiY
IHqXvgebpojTX41jel9me3TrV8sOa1FJGAvYozbD+ad88dhsfYiNNILyrngObDcq
gBw6Cta0YbqaviDePk05LuYyhy+UWvitEI8Iep/ubCZnVBku7YuEQOaR7l3SZ41Y
c5X0sk/fstJeQZD+q/RdHiHGFMwT51D9Hk/0nBXgxaefaeb5LEBzsVhcp7F1dwRe
XyibyS82c870AY9+ztD1DeGfQgAkbL4eStRKp5pQXIqe12jS32jHVyU+zkzgEsez
FwS5ZMXHsFDgghbIKmJxsisbfSvZUWWQq+3qW+RfEWDYD/Q84kvwUs+o7yKr6NH5
4cilc8FdFU7d/g3zmaulC6Q+nSANMZieiUJ4iacvSEqwPFKSQ4Y2MKUsHr48mKLP
PlfGIWTdzLJpbFyHn/XtqOn7WH/5NoDY7sF+71b3U53wZ6qDfh0pBGsYcqrSSr9v
3hepuOgHJxkNcNszDdy1o8bpHwVLZWji7nVseNEJ3xzfOvLf14Oym6Vbmv6AJgEI
r8AUYudQV95Ri8sity/WSkNW2x8BFL5slAzyf+hKtnWdShFCiLTHQVoEcFsAyoP6
phkwxZq8tL2/QifNJ35IK+vx4HPXm4Hoq/3LXgaYxyVsWhgrFPZ8ObcPGykT2eCH
6i2LmwkDrHKBOgHauOR+WsWZHepRCHP0Xr699hgQ78baZzKo69KHc4zWj7xAcrZ7
KF+GhU9bb8HnRvYUxp1T6iaUlPs2i3g/sKQ3eX/fMBVKSdPo+wbaaFS7PDpVPC9H
OOwlwIr+p7BYSW1I5i0YKSMPeEOolzAPrRt1EfjluJsUJDQ3vesK4BMYcZ0w/hq7
RZ0IwmKbyjVr1hHaXo6asyhV0VsEZHokZ/vFkTe1WHdKHDTzBI8o9otVUwsnO0xL
ohC7JQNy445NEP9zFlXXgm0rFtpK2hBIUTxwiFZvckuJ+pDylT/yjBRQzwHwkc1s
2/2/C3FBAtoh5wSwt1w1vQSVaZ1RKscbQzQvImXQCJiSWz4g3bqP+COK2i7KYv+Z
GAe1W22UwrH/jjzpT46oVBm2+fwro/7ni6qH36U6jXx2MRk36mH7p6FAjz1x9TMS
XP83aFsId4k6aCsvEhwWI2iCnkmRg+aX7KBLVfXBRDLWdHs3uPd1Ymp7LFxusZuk
VG32wreRejlGpDRsiKYfnP7kyelFZiVdGcaW8ZDG6WTRBmUncWNNaadH0AolCasK
qD59UC50H6Xw8HQLhhHZpLgM5nZ1m7r2ZOSI8cAc9ayJ2FOSGpOr6t4DRGysZYd2
IbWKPeC8mbiOSqIf2RZrdQpNHMDGiynJ6Ezxt26DGNA9n1CGt8jKS1Ek/gGgTjts
inHredIm0eZnwIA0JUvZUg0oazB+bZmCNOl9FHYEBA83+UzGUy9XDcycLps64Re3
gK/zY0R/KsYD++9BePKfwcBm4zhcFoj8JWHC0/hAl3nOvReW+7OJARggOKJSM9ZE
gAGT/NuaZYFytnnjvjGCq8cpkMaQcltqC+6imd8PSI5osU9Gx5M/XkSZnlzsO7Kg
Te4PAgbOqKSy3yytLDIkKET5fsxp176E6nv6YuBN9cjuXt2RdCzGQ6vVLEBeHmzG
qO9Eu9McG+n3e7lg1+nuOGX24GsNYZulTtCvWI+i9LboQYNzrXQDzdQtMXvWQw+D
MG1XwEUfh4eSt37uFQOIlQ35HRp+e06/BIeIRgcFb5iYnJNja4i8mTthEH3/jk/+
S429rF0dpuULOjh2vDzXV6xyepQw/Zh59vpMkFsMUCQBhtkfxJUcvTGOf9Tgd7ij
e/RnBgkRwT7uBFPsfGHDqgBYGYAPrw45jeaSJPGF2C90v3B/EUZFmVNkvx5lNPHI
sfzKZ50W5EDa12PfswpeZDHCYJeu5Le/yqaFWr2iXnJC4V31C3plVu+gsiF5b7CZ
SyCRZtZsAQ2LTu4k4AlnsZjq8tpHMz4cLuEJLfY5Qb6Arasu64z6ahpKBaLKCbWz
Ps16YcI7C9axzfzK44RauMegRRT7dIL41yBtJAbNhzF0fXFvGEazeQHN3kRf8/Ey
LcMhMuWQg+9RCWZCnZcClwva1H593KrxzaYLsVxlecmibZVT+ytYngvA9GPwhCIB
dh3jvmUOLR84Fr24YVrpt9QlczMYgowRgvFFpLRf5Ty17ijsNw9mSWcATxR+r5OL
ttLt3mPBHUfqVs2M8xu0cNvA2Cg7bPF90nbQowyoF5qXLnqUMaJJJrRH5pNy5auk
Xr4wAry+ysmRJzoUR0WznnvAcC1voV+1cT+FTlivmwKxQFh9HpflEyeqESnxP9od
teJ1mDgPW/gXGnbyQ/9XC726xxj0B2BQxVQyR9pHAEqKGKvMU0Sh/ihAGiMzLOlo
07IVz7nYZY1IGb7WhFY1voL0me5DB47tK/IA+D61AfIvFEprkv3J1ao5L1spX2iT
WxYHqvHIxD6pgrTe7lsnEBYo+u6Fh/Q4Mlsw4RMRZtqSaZ4eZtDjc+E2JoNIGOqr
vfUENxQQDZ9QMWESfPdgdaue5/M4M2S1u/JQvceIJpbGzUJc77zB5+5wliOvzheu
6tEwvj3um19Fo3Lnkh4vCWjr6/vtQQNdV6nDXYVlup7vWgtueBlDG41BrUizNV07
CqM9MYinPqy7TLNx8JNIPP+5wLattV0Lns2L5VbhNVunfsPJfPM1ZfvpIJfGquHC
zuQP5mcMlHleBt/tmTaG1YVDyKyUHmH1/dProgfoCulUut3PLqu4Nk/zfXfr6lFX
J/yCm8tjpkJ2RJgISkVuIN+JRR4Hk/646+c1/RAC3gEiWdPT3HcGxsKDKwBoIOPM
ENJkqJdeghNzHJVuRpNdUHmlOhDEch7pI4/HaEE+zGu1CpOxjGIV+rxu7EhbED+0
cBDnzaJfmWAsSrh0Z1eWpghEFXaXyxaCjVQMQHOb71+eebLN5hBiTzMNYsIeXh3p
JmGGbgKKbK71c89kTzHBsb4SyGYvqdaJlHqltK9Go0hHkScwm5gB5IAkTgt1SILv
ptUdCHrtZqtc22lwl+0vecah69XnFx+PPN8n37wS3kTkSPdNUng431rxqasw4goq
tF42LjNfQ6xZIsCnJDRfCulCQauregk1ZBW5N2V6kL8OcZJ4X4JmTgy31EKV7dax
6MvHoRPsaWMNzXTLslZJCNS/e1ZLp5KRUg3kZwNbZaALYh3tlcSkD+jXEGAwvrmP
USHKbPxahZOqx+2CLlEolKjSsS72rI9O5qZPpkJ99TNj/nL+6s8sCviMMvoPDzax
anYEP27su235LMuoAM+IuUqXwZSmfhhC/k+oiW47V1deRxmtjJdlOmpHXgtXiYLe
rnjJDvW41T0+CsCWi4jJih7iNeJgBU0B7PmrwrOyRzNvxTI5JrH1RBMjqN+xzvuK
1TjqkQ54b/7oIIBisN72E6yV1f9+yzhgCjitdUxRzsyEaZJmR5tlWEmRznJZ4kc9
djZljtp3t29CFP2HQrRWcIW8J5Kf4Sgf4sWmDvsNV0JzhsrZLgDcu9S850QnpumN
Z6F/kOGSkdEUCivjYXDBBWvYDZSgnUg2ElvGEm8ipc38/0tMS/QjdfEd6gZR6Q7R
g/y4X1fvSFj04EQ2i2NGNNLZlzCzItTb6Mj0gh7y2R7KVtDwTs36xS+D9GnZeQ1C
eJ+Ksh6JMJ+0fgn0k5ooiyiGZjLw+qLymnf2M6TyGXFrCY6rb8TvOS4gpyw8fk/i
lHq/mIUd28zNR+ejB4opByCGK7NL/12iKG66MkE/HrgyM+SyjH+5mvKcGuA7sQ/Q
08iPhhonllSIezDr79D2vs8/SvsBTt04xuahT1rJVnR2IMjxQR3axbJLy69UQcoo
9ZGxLlG274M46C15Dm6gUEipFUJjHxFQeNRlNbCru08pl8yNoT7h1ZQDCKMV1buS
HynnQs1vWpU0zh/E8D4QmBMW7yafFATODtmVPYC5wuBnlXCSkZzdcayQ/VZoynN4
XNwerK2BhjYheqkIvioRmlmpLpgxzdpUtlpcT4EZ2TCoQp/bVmonGCBArIKwNmRL
7Ciat8XVRsVcdgYzySzDdptkApHop+ez4fUycfkcmksv0ldaNCx2zC+GkMluJDaw
4nQAROp9c92VmSg3q/wgi1UJmsGRvWPm7QvDY4vj/VgAHZ8h2n6JKfUfMUMBMHOL
htB/bnCYK1fzHDzrwG8d4yuS0NGyBl7caS/k+H5hokJuzThQdWvyxnNGx3awD2yT
TZ6WcqQW4guicqB0A2aaQ8n3zQyGJs8QR0G3YtxUEc/p/Sd09Ejdc5och3NUOHoV
IMuoTCMxVbVvaEoAT9lDlx+vEqmxJSbqTXjC2BLFizxeQ83oryvK6sqN1sXJXnnm
8nkMZkMkRNzKE90bsfvqqVEUZYNV8Q41gdZkflWUFRDTWsRxsHQn1CKaT3KHdP1E
mKd8usA5QXkcXNR+WG//9evfU0oAiwW2PuX2UzuSXKPJ/SmaeP6Rm9w34fgt3VEy
pZf7QG7mesG31BK5Fl3ezcCSGkv5eBSsei/eiRTThVwzeCBXHYKB8LCwSgv9kaz2
mVrPbCu1aR4p+lmX2mXQM3J0Qt3QvrVnJrzI5CtOb532A6/DucBlIkeARQ2DhWsw
0czRvCT10yiba2M4zswNgYuj+ZEZCwF8j4e5RmBWYRbIOGKkw+HwAmGdo+oaymHH
58Gl0hp0wnCZCJSV5u8XFnCtf6fjG6qvlMq0ryNypBJDxSsnn9Bj2QysJlVVWxmJ
GVwZRv3XNSaCDH1DhPm16/7LzAwlEcmDDit96Lb5wqIEH569SEmPMz4rXNcAdsWw
ztYcnpIDR560H1JrMkuQSovpIapHvYS9Nd4Bh3fCTwOQdrO4gJmICB6vjKKr27dC
X+t6pxi52yisL+ClQABu7VKfskWAL+6mHX3VbrQLxVufLDiRHNDZq3WtjjnE39kg
fa+YGipF1a6EmzYkBz6SXPbckwi+asgiqkzR0KhohVTEFc9ZbJmYJJZ3ZDvhFgdo
KeaFNtu0DVAWHKuX1qtqgmUj6kpbxgyMePp5rthxA9hyYMtphQAeNuSmbuDQD1Nu
CGEeDACknO8NzQeJngHXuADDfRDupn8k9uShoxUqNNxY883x9SXZ73ctte5/kmIG
bp6B6FLCapuPB/p8nn5deMD8oznTL/KmfDTXcmldcwH8MdaimVQa0/Z8r3iamPC8
rcziRwJdaNknmBCziJAlNfyIYuEtEyt0JBZqTmD3e0KQ3bQLsvvqeUjrlQLApmgE
6Y/dHdygnOtqIGekHL3xepPbtrsgZMTl+Zw42mlgXTcx6tkXuI7nEFHQpjta5Ldl
SoF0TQNONvNA6GNttKry2ywHRF3rR22M4moXLNI112k/zDNTOUvZxuUwsl5/lWxj
6CCDmRMX5zgHu27fT7i5MT/Z/VzT5NrQe3/5XB2zm5zR/Z8wFWo+OtfFJdjAOSC1
K3tDY7aoHjT7QhrSTcmPAyOo6jDzUoYURQZqHPQud17a/82NUj9j+vZ8gZyewV+d
ksSkCyjjxm9/0B5FUOydA2p+gVHvxIYBJtTSyuM6JEWMTbdjNQM/uJiUepxAH80Z
9vfkWheLOPSnLTwjtWRi+fSoiFsrD5/d6mq+lhO99H/7l3bJLd9/5YL5svKGEI9x
VDMOwQMXyKHMK8RvN3tPfJPhHqtUbFPi08+cgpElky8xDlm89mfvXB+qmsoXDnus
WWjYfzZ8twyhER1CdWBO+g/7l9QGTkrB7DSQ0MWVA4Ama9fZw0mUNshtOkP3nI+x
JF99Ln2LP/saGLsIPAOAEffFCfH5EF1/tOKNaiELlibexT+iq7sI2+KOKkjukior
nmXUfosLeFQnosgn9VwWa0efxbOwdnumUMDBbry8HWnt77/DHxb9lIm6bCaCuIUI
5n6kZ0OSPzfBwicmr1u76BMqxXyg11aR6cx6BzGfdxpTfQs9kPv3p2dKv+3dETZo
6ifwznis6hJjmSL9dU8C2xYDSvmCWMwgsCL+mbFynK2srJZnhZYJ0Ox2LG0szDlg
VtrK/F/qlcFQkCl9Qt2Occ5EXP7QPWfGrgTaMBPCQwumlPryeJVCuQl5ex7NmIYR
YsjvvGUkfWVOuNWPls7KEtizFfpSq9ozsPf+1PtbuccgTEQOO3mvcIMOK2vmddnw
kAX9R1bpHimZdKlwQcq+GfwezbHQHs+/c3WgaJrrezRUEDpZDvqWBJT1WLUh73AM
nCUel14+C96vst3WsSLJcnyn9uDIQwKWwkJh/93FduKPbnRnxBk1lx1NCQ4TWQEW
0UsopFgKWDWfmYLUM0/oyE3oXQKfaCPR55mxpZZRaFoxjuzO/r1XZrS9dQRDaSwp
5or0gY8g5O4of7+lSzf5kjfBF+Ay0oJgIlgUnD0UaG6mp7yjM2q/LJRo+Q4OOtqc
tSt74sJDb5IZUi6dLHjGY4xphikS6+/iQx8lP9ex5xhEPmNGO4PbL3RcpQ9kwkqY
QxuOQNKy0s1PZ6NmEj5ufTxeyGnOkou5SgqKCrC3bzPzuP8JnvoxtCYizDIHD2Eq
wKfLsgMWC6oY7iHokVWhCYdPqJt6JlHCSsa1+XLg32KBmOHyFfedR50o+W5GcwWX
sXUWGPJSPo8mFXwOJSSa1CZ36lNsecXXeJxETXQiGfltDQERU3Y0ZlfX6MEpmn/4
Dgu/3u5I18UO6Hy9JAeob8iJEvoKK485Lv7B3P/4sfXgtwdyzTGxDmnDqQKo8g7o
dRmEdriZgwsQgFAZrg0pc3BoPudobAGKEqgikp9BAWZNBX1/MU/kkmtXaxNZUx5Z
IjabEULxWXKpjhylarz3ywi0PWFn06hKl1QBL4R9sSjRWb6b05Cc8KryXr72nGUd
bnYWUlOBOawiuiaRIvqyDXz/omJnHE21f/yauWdUYpbKURzpM9Z16F7YA647KPLG
i9hhBMNxf7TbNsGBeKOesFYTgpl2L4RJW4Zyuo704btrfhM9SCpC2RzTgIqsIXOJ
EfcNpj/weH2Fsze5f6wll8v5k+zVIqqoZ/2fdKUBvLZqRgAnJOFBuwAVeV3c1yHG
b70uyUmM5sN5lVYvUUX4wE8jITUcFszmZW8zuhZSnS3gVlc8/o3l7ecGwbKG1m8O
9Pwq/z2in1ENjnKcl/NHYl6CEuf5Ty7/ecq8BoWSH2d1nT1qUd1IBHDLdkYabFT3
plXcOdbE7bSMjCYX4cqqgYaTGUExhubjY3CvFEGtqYvcuHUl00FRau5ygMEWqjW2
CQc2hloKZf+zEGAqsaVkAefP0t3AzRiP/vA2pNWndtSITsXUxjzLF/sCHzdw6DpG
cONM3TTX/a9YzGjGXu++aTlHdUt9to9P+uNeLmNDf6nK7LM3rF3qW0JKuIqmRUNu
y9Q0CuDWYpxueH/QJHuTYCb5FLMRBhaKMkz1wcQZdNoVoLreGQZCiW2mwC5c69rr
mxBYejUsBhryEWMC1xdDV+vGsyB/c6s3BKcTnGAcgxObrNy73bqk8KW5GLTgQTUu
GGBAVornu6dNS6Aan59WKfqfXvCXSRv3JJjjT0f73R2NpgIQh1TBvfEfMeu6E7dl
fS7LEIbApRBaTDja6sal0jNCH6FvsgQH39q2aFK9/CTHv4yQkEJCzDO0H5ucxl5H
YqaIfO4ZNQQJoLQS7glHm90kbyDFw+WnwYXdbtLJ87hPjGCZKFH3VJeoDL+Zw9NX
UZrG6giGKBtdR4vLMNQvZi9Z+gREppH0K5oeRltgw2WXlFc52rNU/Q1JmF7C/8hZ
jWD9nNtjWAlNJPz+W57s4FrHNd1VDla+EPdN0L9CayBbCR7oFL7A99VZfV3+UwkS
4CxWLtAMu6JGUQCELa4DrTT+mZYEUsTb0T3nqNl2dCbUgU34UHgruy7efbUstnqd
4yY29O5g18sf+zfAz1plXOOZTGIuulJYPgK1W/0oMx4v10/XEQyWe5kFOVcKU05r
qUuY3cIdmFlqLqgb0w2AaumHFa3CjI7y+zMKYPkbrEMe1uUyi3TxH6EKhGkDCo7f
dBJo86L5Ql3phuLisTZ9WTGThFcx/c07KOX3BP/zvc3SElsaxPKr0aNEV8yy596E
4fVtZir14ZnqKexaG+oTqgETlaspTlMRAzAnz432MtLwRd68gfhChP+SoUVR+/Rx
swy++1GFPGLI/9Jzb3fcR6lWqFegpb+WYSds0uiGqoWjNOTTD3gqzvxXyKzppq2S
Gfi7hS0L4JaoAK8DU+hYu+EnPqnTdWdGmHSp7Oqlwy6U1j5kt5YS0KinWsIIWjF0
ewLjgpwN2m6Rt5j8CaTmBYtawzRlMaSJSBjqZghxIpaXAxG1lemqlKkbEyLrZlT+
9bQH1a3X8Xtl2tG5/frd8fnh3bMpukhRpsqedWKQvSmlbiew6GzlE5uD0e5ZP0Gw
TVUlPpdz9w7qxeYFa7MIniv9JZqtPTxM9AzoQCx9V4SQQZd+LNxW4LjNxvklPY0N
iFwJta0UD+wfSSncGyf0+DZ2o8VUaGoOfZKEMdTadzn135ilh3Xu2Cng61f/WXjO
hlXuFmUtxqJ7dj5pSgvjuj5paF0XLVsugzEoGRW4qKjMOA7lutcrxfMsdoX1qPqP
9wyU+HXWyQGXNfBLO26/3kVgs9GdpqnQF4xWYCnO8rq3QT+DJ34uoBEsK1DGffC5
MBBxjoSDwU1Yju8IJwRxdSepd37L3bslezFbzmv5jgjDXzfua+3KRuS/aW62JnBO
1LZrdQ2wfJ/4RfJV3orgdFxjHNHrCCJUBDw3Dmb7psb3Sk1qM4JlTkrct9TTSRPU
m9fv9H7aU8LCNyqPm3vf0JeN9Mzj1sgtb1xpJTLW2KuOmWMZXdkFzCsJBZEBWueU
xyv2GxY75/qhdqA503MUT+kUstaPZlknrY5ve4adju+OZ0QkFEUjAwku258HVe+j
h+ndjQb1K3BpofV7aF3FRZC0B832RN/HUQvMZp2yWVYXr251TK3Fa49Z+rw0tzoB
Io8uYqo6f3AngCS7nlG/VzEyPGls2WgwTN/oHw8NoaZpoaIwMFFkxLhFhSoO1HCk
r2PMPx3lwwkaEpg4CnqVbsDTW7AZotqq3fcHzVB5vbInuguwklMsx90kCWdGBnID
swRjsJTf7BLDz4YgqSHAnHvdKDEkKrrFjAKwE/8GvBhDYUQ/xeKNDmBBT7TyLPNj
8XTowQYFiKiwi68n/6ajhPlIt6cvQ9d07rxCGHrIfyWmOhVAe3FGKKqx+UK626xa
MQD7N7XNh6LAzdSe3L1PQB3w2mnntMOAiCW46KYrxhlaEgLXaiwloLG+pfezPa9u
+AZZnGqsNG0F1YtALrBTAhidfRCOGw3PnZ/Tli/DxQtm3KR+Hol6UhfldQmquSv+
bqalf+U3lLFnJxhT5NoKoDRerjFKWsQ9waSecHWRgKWzYfXT0fZtRhGHQAt+Z+8t
pZGHdYMr+Wr0ZgFNc2j8VdFKwB8U5C3MAsuMB7YdeIgAntepByJcx/Q/vpB1BtBo
cyCcbG0Zyta72SygQLCo+OtG8ZTAj0Sb1oqya2HVzjLSgB9IgXpB1PLGmObN8RNp
OhLRDVjyZIed++jPzWIjMtE6kxzibCyW16CAN/0TmKKbbRjKLo1hEecSP2cFEGqh
b9lryt+dadYERbpvxQi4tGZXDfisPyjsm/PP1Qa1IfinLPHHCSbgJhKyjMT2E1UV
2Iv3Xb2dMrAqC8PsFojOenA6+t7uIJ+fGoRUyYMRpjkKzygueZloL9/zQCo553hy
MDV+Z97y7mQtddlWz/P3JL+VhE7QXUzVNL+x3dJe6x12RrCByuRry8JT6MPMv2uv
lNs4BXeBBj2v2xXzjU7a6F4tXgmsDnkJ5Q/qaK+Qil61Br/jSN5KlwUpvkhcclN0
ZaD5soImxHPIc/MFxo1KmtIPTAyDkMiyGibHb/QSxzkqAb0rzm99LUm4g4eADDq2
ncCI73F54HoKgAzsS1aShWbUPw7p0+aSJhr1LJ1DiYfb2+9CBMeIMkCnFoqScVe9
H+13qdpDR6N6KvOHC5PE+ZNaReYSkPW3afQ/VDJ2nVFgq4yD388xG45eGBjM0yPw
3HtM/AysVLDGkJdKaYXsDfM1ySOILX7o+dNt08HnOc5dY+0GzTyks0yqM9ZC2WAu
jzWO39u2F5vA9gSkT2xycGfcUURdLjUtEBK3Qa2ZPr6TvinsfYnp//vr1nBATgow
ZneCzFZI+aFsdzHretkq3moJXffLujxfc4N5qizSqtZHQAxPpZVsYC7YusbNgSO+
CbNRprlk1zt+uGsV+evHtWPZH4oG9Ysp+WdG1ebaki/V7Nv/5oKsb9yEPyfxcmU8
pFKBD1i0I8PtnIB4ahC819l5n3U7w4eDXyJnKDFBorWVma0hd7/SbO7XSkJyEInx
VGMB8PKSm348H0fSvO+GjceGosyqhiIavm55oWAZnXTYglF2pD8cBa3kE3owlDOM
nHxkSD7uVNCBWElpmXQ9C32unqUx9NKwpCxq57A3DjRJXzFUN+gb7C+SY5KIpx0y
N+pLzo+Kjz1k5ej+HUPRAUzDeO20G2bqMU4PHhzMuyh5j0TSP3uAXFIDXZaym25j
SF4lucLvObuqHnuqWHHSSyZM4nnplAvcAbH8K/xxhT3ew+O5iRGLMR3Vfa2/6stG
N2YP2A8ooqvFT1PWHjN9bm7Dhcw0CDz3D+Ft6jDL7tCOtqKEAySzhJKJc+YYaEM5
Of1IQLgHZkCQza0WJJ5u28Gdtwa8/DkwktxEAN4rthkbEmvmO2z/fYUMMJJBo/gF
OpxYC9TcLc+Shl/pGPSxXZKRkku4pmMHUTPe6oCGiQg4eD4PW1ZBANqc9ZyyoZfO
pghzth53J1dfnEGbt6h4gXzKARq9bZWwUkn10dVIqxTeTuh46PtcicnHyGPomWBb
j9UmVX9sv6xoSkzZzNhEFvheUDUzr+l+ifb42ViTAbz1R+n+ySuEiGUm5iD8zmFl
Ud+JdpaThT7gHgBKnO3iv7YIQsE+rhepHZ1MznsM1ImZ/nqA5jnIdOQ0Tg3FXvKA
greb7sq3czbsr6u2i/jAYP3kgbfgBEQoqlozhbFrflojf9BrE4ArgNzYOKagUzLk
VSrLuH+KoVBX4Y/PvmL3exCE8/diZSa0Hry+rdk9wBvPcQGQJN/Buf54w/d+mPA5
uN+Opn88UZK7z7Te2GEnvo3OuKNhpnpmwb3TKzYZkJLEW2YsJEybfDuiSFzORbBs
+l4Ve8vrlsuQ5lV5Xua5UoXuMLNam4VpY6uN2WsnIfRWSeWOjjrIVRhl6PTKkdzh
uleLMW0VlQjBCW8um6SGDYCU3Kn//xn3FSMqYeIkaXhDSYvCRcyMsgYojfDZrH9L
QtvQ1in4NLhARbA0VZ4MUSfnZ2yArGqUtCrkfg6DPx0O7I7w6/bdt5b/IB/Z1JjN
8kF+fWF55JQQ6MK2N0qAoymdivI9Hb7qiiBxDVQHTN6BF+IWm2CfzcJgvqEBo/1t
GK/po+isIfPytWUHdMA44F5MHVTAFjLvT7B/lOmUSPMZoNTHiaF60PnPNcJPcL9Z
ZqtkcbHnf8DHV2ZqTTk2Y9M0Hd7tbmBlvb8r2f2CopRGZM5ZxMtGwEu7TKhNgOAv
4HmO+QCv3j+nGqq1bnJsT0p8JikYehN7BlMAkCX0zyg4dD4R81h+DOrZdkZpR3LF
AgHgLEQ8UEcVff7hzER2XyTCbh7HrK4LxQJNy6eqrYgLW4wv+HNFbsmRdffkky+t
pgiy1+ymZo3AbwbvGY1mKc6Qf4z2hAWww5mg/ws0BW8Q4wA9CC/WFNEcE4A0rVhN
GoG8vrfHrQnWNphBr/cJ4Exvaz99ypOuErNfIlPq8WGFV1emunAUjTnXeD04cm/X
Xd9WQK/rJukBo8L8vyvjVy6mPqiHSSoBgfPUXmJOt0/VirH7K/F08R44ts1oFMIt
YeX/H5Wkl7wcNvRHLi8+ALQbomJCyx4VMiM9vwCjWeqAROUEow9PZ4/v6TstbV41
6fVQuh6//ll5XT4fmFQ6jgBRVTBkk0bJWW4Fi/+upSqMlQVCTMXYU/miGshAkx0e
8TBnWHLo1sX2tu39s537Wn6pMSTWrqFFRdeX5AyKWCFsijmHbmZe2WmpZNc0LjJK
Y4RJ7HOc6rY+8XY/jpyVHMBWgfya1Pw5HS6kxcMh63b1zODCMbYQ65Td4DnEous7
/L76/z2afnXUE+DtNZpcdmrso2dxAWfWxUrQ4vIXxzHW7F07Gss/fTXh3Hb0d9ir
J4Qfjn4NVsxjOHHbD4xlX+HP7n7sR41Vrm4CU7I2SKvDE97dIyIkARjN/zfnHNFv
MZZLNbQdysNDcIQxVf/sE6U9sVlfqcCDp7UcLJs2F7o+ve6t0T8QH3End5ftHeaw
hAJfpEm7aMAofe8HPAGoHOIXhCF3bsxuo2vfC63XpbQxJBZLGUnMryvCOyBJcywp
M8cWGtc4z6y82wxdYDXcVgoW9PdGQ5CGe/VEHyGN4HptBFabfTk8+zkq92oDUROT
EGGlE1qKJHU3m+Jm5fSB7i1zmy8X+RgOWCBvnPIckVBwgJvySiHKH/puuceUeEgK
Sc1+qAri1yC7Z489wnbsxFWECcgCwhZ62V5iTzNfxK+h6HkJ88Voapa5Ct1jDESH
do/BPv1puZ/sl73udu9GWEfN9F6eoxCizYVcWkiWR15pvLpgqyFl8QEwGYIvI+r4
qnjnI/DfPeTwT1KKu9A9mvxpFNYsgXeWGO6i/YVERr5CALZZ0kotbYo8fYrx/tuT
uOQgOY//Qcy04A9MTn5dMDGhHo7kXRwZhL6sQpPI74s870rsgtLwtiA4FG8wLMrt
N8s34mNjql4n1EKOezFtRTt/lyraizRuWJYh47j7sBF4/LKjHsmf3+14TCRZGVtx
JLPKdkm8goENOpd7gtzysi+WHT7DbxlN/zYHerk7wVGga+hrWKMd/aaMJwdO+JrF
UlAtTv9KXl9wdstdJ8JAJyCJ+eSpO5jRF09UdHwSDtPKXzAVIcY2tvE5w46isl12
/Zy1iSB2KpIqmxNXQqlE/JhucSiQyVz3kJeiRPm8/EMaN2QlxcwPUaqP4e7BoDr0
wKOmlWn0r7ekuZ5ZVoDmE6ChuoF0j5oe3K9DlozqoCFkgkXK3UIns/EWrz02ERmf
sbeYGft5QFlOOf0nBFVyWRiP+zemSlDAfu6salqRK4uMxGCtfJ9qifG1ObHSxpxh
v5Ap/tBaK9+8SfxzN+oNs71glcle1zM3bfjIGmRtnwYvIr5IcyYK6O1DGej5Hu6/
Iq6+4lgRcw9Jr1QsHDbkdeSVz/NXMoipzhA8fMVNM1oJQxzLkhScHrMjEjrdy8co
geVDjLgzDLHfu4GzjNtAzWn1vE9wvFkVgV4F6NI/ii7++vkx++W5jh/B4iJlwADr
FPTabBq3I5wCPl21TizVY3vXzhJsfsljXCaWUwEsUe/W1SzZ/mX3Nksmnr1tguUV
ps74XZkFhT5xhzk9GKlI0Iu+1sSsnGIZM+aCkkE8s7j0n6mzKa6KUuXbcZYGOV7n
cC2Vm0yU/7rpIkLpTM0w3SsEbv3u3WOBSR+jTybgOv8wWy/BsfzSx9HQGV/Dn9cy
Z5rsGBwsJjWTwCkyGDYzRPxxyy7VO5/L5xxXX9XQ/I270eoVULDZvAxypCGi0hYC
P8LiddA7MiNXscWIK+u8Kx0AbkF8IfisO6XLEB30tlmpJcDVv2k1riobhMDt8gye
/BIZDxyeVyDLQ0M+mz1xuvjr3NWXZhsCWdI4vJk353ka6KMSQ8KAYY1HhbPPsFMZ
rqMkqN/4shHhZbWCsCzLkMJhEq5dplGUR4phaE8qYO9N37DmKW1HFwWcVLVDWoFa
BJicZFgQSmu0FQfMmFKi7akqHpGS2FUGvvXlcufcQs1z7zTRvmCMp2Ez4NLc+Ivq
YnFae6Ct/V4SQX+yLIvNYyaggfEKtLMYFHgbgdYoQ825nsMTacD5reN163C0C76n
s8Pvt84/NFu/iyH4qdoxprLVPGu839kC84J0M+O2uZC+yaw+dnKibrK+Ih0hncD6
dwfji5maIV7waug22x4Z/Y8s7e+7o+5XOsNounOPA2yvsfSZsVAFCNnP8Sy4ri4B
AjwrZkVftiNWp6VhA8FQufwnI61t+/dRVWs9BVc5DRbRf/Z0U1Hg3gQCtCOAtgAO
5j4e8nr/1JWwszisbBAwp+uVx1n19ghqv/DJ5XKseaU+C5jy3Lk3Y8mCigle0rks
0waCBiodvhGn76jhE6HazkvIU5GEjQ44OqkFFKTcCUx6vP7CeiCsiu5fX8iEK6mU
reVTIKZP+Ox3Tb+eiadC4cW/kJmn5CbmG047i3NTLAFaT7gkU5VpyVLtxh6uauyU
Uk5pD6TMaQfUg14fZvs5GHaLnri3Xe9KzPKGdpQ1BFZLpNuP7Yc8HMGHfuhS+hLf
jPCKUV+lnRBAnqzHSoGVobaDGZQF4dKnsC48IWUa45a+X+73ZXRkvF18K6yUq1lh
o3xX+VJwW3hfuKlxdDgzde173Nlr86nAg5Hh1H5i+oUyT6ubPu7o8tQ521kSsw4g
OtU8RfEAetk+dudNIuvZGD4WbCJ6gLvUlaDdqZFbBCnGcPk6bSe1zyuvkYvD+8cB
bDosSl+UDZF2GbWlVW+sAl6xUstLn9Bisfo8u8fvuzaaF1DuQOEb9L/ZJr64KqpC
rimNUwaWvEJM5Ssy5CZDCDuLxRj49JY4NgISqrd2DvM3nhrNNE2TmXKvvjBx5bNZ
yaS5BKck5EbM9OI3RPDtyE6pG9ZK8nQ7s38RzsRO3f2QydtE7A8OD3O6VtV41IQZ
OpSxj+lzTN0BSlqdFbERx1z0J3DvvsSnQlwQ4cQgR8dOMoHONJghBDg4ixMPHSAo
Aqh75RnqLhq0/y/ArriEEUHzFPFnZ99o8u/ZJRYEb2ITc5HtZ1Ah99JKsBC6JCLW
aH1Lunwx192ZkH4p3pW/IQd/k3AcjIkx8wjpZtau03z9ZCDlFXQlY65n1iPIch1X
hw+fc2zC02BGP1do+CmCK2dHM51Lx/5HHmGSSZcYsTD+bW5xINQSe6O7DHKLy0vv
8U+de/vVqttwZxB/jqwBx+UD+dDPAxCF7yTRgYAh3Qa2Td4N2kfEZeXmuE7eeJaN
MhMnbkn8MEL5blyQ4gtvX+nRpAZqSbdBZe6V1JTzr4j2DhFmqCgjm9ibJBYlfuOo
Sv0R+M3f/w0hr1/IqlyURY6z44t3nxU5Sqi32ssdn1KaAegqNBfuEUFl99v68IHn
BlDCP/WjJrIcHHnrBuUL5/jKJqLzYoc9U+mnasT2tqu5s1TiO43FJMPewQeqQ8go
6EgyiuKhzUV+T9UpHy5cAEA+c1zQ7PGVjDjA6f8dm7gQXKs84NR1pcd7cnK+o23b
1+UTh2WpPKEoPO419bmE80cmP7i0K272nB9HEt2E40XBaZ6qm7GgqJ7pO+ro/k9l
/gx8swARJrV74Bqmp6bDKQ/397dFxSokWcbrnjJ6fBlZN26Wuwjfwm1XgawcMb03
k0s0TeZtKIvYqEJ67jUkFhJxVnvqohghf592J9ckRkDavhM7/RQO/NlLQlJl/3dd
Nxejj7CTiunUJwS2c6Sm9qt01KK4vsabSNnyi4SrgSn8QR5vyGQ4cycAoxscAKRW
6nVrMe2j7llkv2YkjNxId7DKj+SqqG/eSWqkFGNEi6dDSV6OBSFlYlksSPy8Vyjk
EhdhGtNy7zUPp+M6vCtTT72LoyN1/qxfaDYrtPNUDWnUwkrvU9NeOHf1kd+dPO9+
5OrATd9yotwWOVIG8fmFgOpt98HQaknyNjHAJvUJCQbzGYgN/yHh/R1eOu0tkJpc
7Pv4oxBMppAsPDjRcrR1Jgku6HgcN+zJsvR3VUcl416pMd3MpsTKDtBrvnxxnK7t
hrOz/hbNl3X3bsa3brYUaxtHtdFNSXrNkFyFEmvtXcNbrUOOnmdW/x43OzRodXQp
ComV02DPulvk9pVqDDKjZaloCqbMHjYFxfjZHbNZH4iDjJpOB9GswvbWuHlVcot2
ieFAcek3cFXtj5aD3QRjQJ87OUpo+P3h1mvY9su/FKWatZejeIftQql9Wk0qhzZe
60rlABI8xS0ZCNx8omCS22OnjnY5b4Y3L+Q5uG6Dj0SWUDgkz+R9ES63f+C7WJah
XDNcEsyBIYvvY1wyuggARDu99Vwinr8t8KGyLoV/+JbtBlgmlXPpaFQVB4mXqNTl
JQhnKaAmWB+I5yvhWt0Q5ZKlZ8POyMs4qFCYl8i1n57qNrA6etYo2FzoFQIRVhhp
j06wDOF8ej9CE2/AYmfZIUaAylxwXI3fUUSl1apm39GdcmG/a/8k7cVQwOhKvR0N
ew3INZPLFXDxSpGdIQZpnjlNlKoaIjEOAlihJD9FZ/igwFuwlH5kxQ3bfyKASD1M
jZJnzGDL6S9dhE2Mr4V/ZKDkP+jSVTENoLA9oAdFe8fiTuFGJ1ntSwPIJxuuGVZE
DViSfIpwQOOA/1F7E16j58GOayx9vRJ29vi2rdtIQcojnOwrvutO7p3wpudYuHB0
+/IIPeOTJfYyag5NdN7hP/gJpqdC/7S7gbCDFqXbcagxSa7NeonM8eE071GBj3WG
rrTEvldH8c8iEdymtSDzB/HuE7Mb6r3K3LVu6YOh8edD4A7QVtBlt4EYpfkmed68
xJKIvTfY0SDgj60qtYQGxgsiey/tgLjN6CJEopS7A9BHqcFvEtzzDnq3IkrwAo1N
y954e9a9OtOU12UiJ18VHCP+dRt4Hlvwt8WODa3+GMB+j/LBfEsBlMuCwYlEOQcw
0oiROzZyaMkr+TiiPb0G/m8k0sG34iXVhHTfDGV4ZdiDrDk8t2rqagXTI8iJ9qvI
RYt20TFYUalLk0ZExUS+XQkCj3A7+45VMNcVLsBkdF7eH6KBZrU2x/HDyW07UE0Z
ARbyZp5dK8xQpc83djGboXAUVHqI7EyTPPJW8WTnliKCXeUkxBZULhuWsLOPaRSO
e1ScDkLBENQQaR1+dZkVP7GeSvNfTAyiBYbjnG3ZkqB2jGB+Shm0hlhXX1/q329e
XVqK1UFX8B5R2hOVlevgxRw8NCi7U4DUrRDkPZkn4gDd1yEehE7Pj33uktLUq1mP
Mj5g1YRcW8w8/V8bZcxbSFoiP9X2O6BM6+HhmanTgMhHufgwfgO76zjbWgZrLyFE
BEnPSooFauZJ+omDG5g/8ZhhZTuSsfdU5g8ZzZNuYqozEKjOosNsm9VZwbYxV9g7
plwtBlfaq+vkTVuSZPBbHLWrTgZ38opJR4ury5eOzqyq+ZgHycWFY8ZGb4EE+DVt
ApA/yb3o2n6Sj5AT03d6tEl6TeN9kZ+qF44TcQ9GUiVPmHZziQNk4agLassRybiB
ZfHzDVoccT4MBt9dnIHJarvpp/goq9hxzgKkAfW69sr+sV3ZMiZNMCitpIa8F8nr
E4fzLVpZl1pBB6qLd8sjP7UY2VZozofCpfzzB8OqoRZuTrboAlJfszpZO7XpIorj
PBbjijsgeKLrOCx4oUgHd08dKmSc6L6Yy4SEL9CjN/qBbacZas81X1j7SF0FKy4m
fsSYbtfZ+GlD6OPQRnq5LDz7Vswt01209RpqxmTCwIE4O7SBX1IYYm3jqgAdp/2J
n/jhGHvFP8/b7neM8Nz+UzgFlMO8O7jmPYgN3JVA7c61IBDsASDNK9ViAt5mk8/V
FDqmBN1gV3S4ATiJDHrv4yPdanuSPEhiMOY+JTWcuXXTFKccBI2R5LI0kxBgXtvr
5IKUYr8uowEJ7nEEFjzI5kxGUKLYq4hT9l1Cpl+Iq30dMeIWi47lEDlm5VkaRH+y
cEj3bKDk9OpJc4woHmkFn8JEgLy3OTO6M+kos0mbH8+w2MGD5QkgCGQ26sTex/pf
ws+bKBILI+Qd/d0Kkxtu9jjHB0z++VeFa3RNIM/8Li12RPN4ztiIr2gojwdHv3zC
LKLl/GzL3dB3FUV2Y440HFqHa3SULaYcuEfIdMj8waexQ8v0wU3Pge5BYfcEcGyR
tPPX69LDSuWSjPXxMgzEX8r/huhqzkMSoRcKQRRSTw86tOCd39tvO1dC9yO/kGkZ
1npBVCM9cmjgxaFY14KlcwbP5l0judbowLMZA5HvGS88iBcPkpK5qCRkuZnM54qv
krDEbzi0QmC5Vjxl15lXuQDjYTwawUstZL/hXi5NIxP6fu+Yt3PgyHKMEeuQmlFL
aIl1jYmVyIA7Q/fihEvGeLGBjH1Z2s30crFdm8II7gMqDrvDHrIZtB47UfeTV8kQ
A0pjWpQPsPcl5lu5YtEW+xv9IkgtY426ByERPcyJ76LB74ZhdGpcUZD0OZ6L0RuC
0EndVdBz9hSya8y+ScxwfSjDRjz4xO/XoZ0/MI57x3D9E+MPfOKIFYyQsIDsK82c
MFJnmSEETWdhWDA4UCjjQtorVkLX6RgppE/k621MPYC7cgCCSxlH/G/Lk7G4TZxz
diSp+VJvGziFacLJQT1mUhxIVh0rvCtLBNDKGG9twE3WO+SEzzCHlnBfS9PJm+LZ
L11bEkSjFzh4VrPNIj2/m5TEMOfShUPwqGynRrZOp1Ns2uVoybPW+JoFFyxjOGwG
NNzEmwyJ5CehPTn94o5jk410h3zuBQ30KlHM2pJ8vdeWN7d2efXHFT4Fm3kBNkSc
mmurvNpH+5jlI3iS10Uy5Ms9M2KqM+Lz6u+cI/4tbDiRQupc5+ANbfDKqmq8Wh6Y
HlwwX37SXSXLx/Tp8Uv5yXceuVzjx51I4P7y6Mk5SOhcGIglwQiY2l9u/oNEgA69
d2FNNGgLNeauAGtc4rBQwHs8UTS5U5wisblZHZeocFo2Gw+YTsTe6wv4kx5ZL+bJ
0f6TnTs8r8LGAmFd8x1aQkDWnW1Efg2GPrcDnR3HuOJo/eAJM+72voaTADv/oGwY
GEQJi80ZiCQVZFBYgLPYW17P1yx1qO4e0/T4URoX+dfmc5hudVsqZ4c7fniLnULA
UbJ6QSTe87zsIB88+SmHj8v9qj8xmnWb7ShbDUp7eapWnfnBDKDOA9wH5fg7JAQz
PPmgQ0tfxso2F9c8EqKemKbz2Ilh7LyKc9dHPswcddFFxQiH9Mj5ip5ezKRTMuhh
hg5lz5FSBwdobMVIqEFYTfPs8JTQJ/Phis7oBNqk+gAUUzRUCRNxnb3HllQQa5z0
rzXaXN30R6lnLb6Cb9CCZ9URsJCEZOEpEspiO0YjU5iui7t2DCh26+LbPw+DNcy4
zighiDPWk6AVaHL5q2FTpKM9P5pYFV47KOQvcL971Nbk0zI75PVee2N5q2TITsta
2P1qM1t6usyEQHXw49Cid5aK81Kotu5B2jEpFe3IfT5uA9114Q+4jSW0l8EXWPRj
wQrvrLGbp9gAAu4DMumj0GZhXtEtN7O/W6fqMB8/sUlyrvS+lmFHRWcbwgFjO8pK
ey2yFO46vu5YHvpu6qzZFKBeQfuk4yjkCCdAOlQ9DpiOwU2wIQzPRBLIsZlPGU/y
YilP9/466BX2Fql7Vdqjr+MooWY0T8Y1eN5mwVNoM3eF0BOEJ3KXLt2ruDvU/wA8
FVLG1OIq11BDKiTY3Vz2+6QkdQwwYSF//PDq0FMB6wYMp7yem+lwlqtrHZPeLrmo
QlD6QPEOA5EY3rOko3YIDQYQ5/8ozlSWCpXS5fqMIK0cm9u8DrlFUjuJ7R2Go3pX
drwoTOaIoDZcGpz/B0KfUm+CEW4S6I5TNGZa2NT2M1RVsXHw5FEH17AeSHPfz0rL
9I8SW7l5L37A/K9rCSq8nw2Agf6kpKgcFb+h9sL2oM2afMjMpqOenL0Kf2Byesg4
WTV/aFDopYXWcI08CrnFZ+pUX2sPmUKa4+56lj7YeYHrrRD//OPZYMaP9iGaboiq
U0iSoETLpuGdbDL1hQve2y63+1v4Wy1MQ4s/FqfNnWTWLLhuY20Kp6kCIAqjPsmN
1Nn96M6+TxXRBIKgxjIPieLFN56i+ARw/hPqx4I2nxrvBy9GskiiFx6Yw7eyTqqg
/NWZz/jAHNMeDfkI6gL6o6S0pf4KcCiM8jodnknO6o8fBwz+F5eM7mKCZNAQBryq
Kh1efWVEW0I5k2w3H2dayc+R47JFZJ88HNjmljb/+Swpf5Ky+sJasvmRll1Xc7x/
yNYxt/0kAC/P7OogN/R73QwthW5z8c1osHCIn6Z9Q2z6iCDJmEnkDCySsxyJgfVb
4E9OzhDjE3dd3BXliRHzGmMlUoG4f/eWD6mJLrIG/ZNw4fUqQANfzZj9aNFH7DyK
myf0O6s3UTFp0ER1guzO/dqM4MWgY16MwQF8p5RpVQtUK/cKLbhI9Tix9fpPpjLi
MT9gzOkEmaPMgdK8tyrxGq1Bi/urO12b4neP09TANnI+39Vc6XcesZTRDOuftNyz
mMXKhaP12dGUpnje+tVHBVG7sh8QPVIWjIbqhkOSoY+PaRytDTdh5bYpu+DQkFeB
X7fETipUhOx8ERbIcdE4K2lvOiqDUjDixcTfkk8JROzb5zVRXmheZWah5bq07O7v
KxFhLf6OLjcnQ+0RQ1cYm0B4PdIPPi3Sk4DA1ctKnajSnrv0+VCEkDzatcWsZ01z
/aCybwgKQvFrveJouKufQDC4yxh3bpGyI3VS1DLFZIidSY1MXekaqRzfrcfH/REP
u3WpIQ6mNNnxKOcGgiij0zLAqVBvFn8ylKutfnmxtDJ9uhov/7rbrXtb1zJYY3NW
3nbxhL9gRQ4Vm3ox7uC5NTzbHptjanuQq2gxET9yyUEcBeOEuzUNuxJ5jESemJIu
kyD9bbwsohTM/K4Ff4EC8IXlHbuLvIMIh6X/iGUxdMBjiCxpYMQcemR3he33DGvk
mnGmy5tJUJkqevMUo0kGejPI1OQU9lKbkFYFBycjeyOuTMDwtmZCp7FVwwaZVaM8
JVAuHYrCPWzjnwRXLz+ZtA5iF1Xoj02FzAEWgAkfY8xFhTgk2eVEulo+EuQlqHzF
6H5ulEb9fVmsoI/BkNnzwGHG27F+5gOsf1aqCHwZGJktXo+QGAlGJ12qiGAg3OKh
0NWNCsNMehkz9ZEl+HqSJjR+wh63o8LAHMnFKvqgmqA65AMHit7NYbzuDwo8+w4T
dn9GbsBdtIPgNjHrRKq8fxsbuFnJyY5N9m1RmFvVNSzd2c++4R1HotF2UlnVz0J2
jMyNgcXmk/Jp/O9KnHsRC2Y/b5shVzKjVcghhR46g7ENtJhYsU11pmNud01gfLrI
6SCWc4VD7aXAsWA04dBnGi+EVM8+K6zFFkwTaQppayoy4NakzXfefopkPmlZ8XIV
pow+hCbLwZpmngwnrMfEyyrw1HQQ/UeEvN/JMpF6AW40/nh/YeQaIaJFryOqLord
8Ky5Q2cdtXGDDvFvoPD9jSY6G26pkrbjxElk73X3SytNd8IKi1BW7aNlYqLinEm5
tjQPv84pqXSokhyrvpSV6ZNvevRvlpRwNAoMaLYxLovAyYHtDJ1odN2XvyxwLkYd
ZNjQP4LtsitsdTdmw/G0zOMM86SKFxAaNJvmfXhN8K0Z/zwGUwQXdZtthA+797JL
3DhvTVITmtGJMWX1gQqt3OKjLO+T+YvvJ5xTl96wj6WuUHTwpQ+UMCOv2cKMoLx3
+xjFQBa2nLKqzsjWmVNuPzvO9W6awoQ4trMXMrosh+/to4IB3gWFB0wMytx0YqMx
WO2kL33N8mniX9VCqeBB5gWcS8vbnNlVNTQFVHxwrlvsXw35WTwDq/rLJv70duah
NYL/aWUgebbD8vTR8otkAByw9v1QrqmFyARIp4PoAlnYCHjtzJobASQZLguS5k0r
yO/iZspyVdJqJtxoTeEoWMPd5LEoY3S5HhHjpoUnayVZ8rRkPXpB5+FEdh2kgPQR
Il/tm9LGYfEFRR5o1WZPkdczqTttubVipnZjeFt60O0r5aIem/bv2aFuf/mdRqTs
oh9fHi9W2QJ07frgYVWAcefITAYMUMe4EHP2vLxJT0sFbqf8xTc3YGdfjEh+qurr
WcoC7GADvIz3PbCcLQkjiuf1VxgJgRSzFp/rd7vbKu1MHJw7jaCQsIgThaDMrgaP
3+1w0Uo6vAJR6etcdHQNRayGpkykDweMV78qjAoMMpA21/yVAqttne/hccJWo989
kW3TiJx17qGtW8IPENTZt5k0+i5XhyCn5CzAsX2+CHm4JXJFtoP+a1fLrIXoSVa2
Yn4QyD2B+61ktPoyXHOeVkcJYvgL0MzrwIOQcvLkNwcDCQKEAg/+u5UzUQPf/J1Q
yk09KQ2vyz+t+Mm3HScc4gtLTzvQxHD/wnSpbEKREEsMrk+xjefmG5M2Zz5Y5OBH
m1e3GhvRQkTVyexDjz8XGv5Q0N72IrTy5IMc+euMsRbl0zvexAZjg6om2M1okAas
Ux7H0J/5W1nxwuzg5jMqj55AxRjm/tzVFWaCcnP8iVgRWLaZEv2NIiFjpa8KjvpR
wXqrokYIfwa4MZ4aJEOEJgpch1IKPDyLCXDkIMzOLWPxHN8FiC17KTtfC7AvzD3+
F4EfbZlbP1a5ZD26ugFPs4dnXkWkwAd6WVrg7W9gi8+ERav0u8Lsb7nHzOAdcqhG
SMr0NIBP5sEs4OuSlT5y18EXsEBkJFFOod5vixou5aYdGjj4ZiEvnSnmG7MvSdKK
I36bE2hGp4/e8Q+2CoaJR+f/KN6fLPi7SIlUKGH62jhOnT0PM4maS2f9bxLmP1NL
OwASewJ2w0q+m66+COqk52+RBjPcpvB05IYTst8UU87NHx8OZKloU0GqXTmFSEgx
vZR3Jusa+l0/9rpM9D/jJuJjWUXr5VQ46x/f3fow29gAxOQe1ltvWKfeYQthPKdy
iORCeLZcfSx2Mt6ZBtkClahZY64lep8fYrijYJuWO2f2qOlTyHLI1t3VP2imlDRU
ra9Dq/8+BoFTnFJv1VhdeNqzHOSMVPiWW0Ypus53lAUX17ttOE+bkOdmxiSiuP7y
uOj2PNOnSjghClnQOunheZj+8U2/XyLbXgfpNNLfJiJKWzZ+J3vaTDBmyGUJ6nny
lAdjU3dhCduSYtO4wdsao4M2dR+ySY7U+QvNXtFz2KRy9x0t4Cx3BOLoGaNoAV3b
rgdL1/C06sevSA2DS9vAV8GJfP/4E3AsVl9X/X0fFVzzoiyYR6pD4YCSIqnKERdg
qiwG91Y+mBGAJTvjcYmO7+u0VHMI4hLyVP4jtOu+n7fVB73DrAUZBvO7UrcrL/FG
DMdnnpVjg4KjQehHO44nXZtyVDTgMzKByijx+QwFkvC79VD5jaJijXIISKg6G8Oa
2N4DNQ8wfnhHRPJ9r+Y73zWrGdugn3Dof8vXhyQZSEqG/D6j3KzgezLtvAeog/3Q
R9gFZHvg7hZsoeC+vyLYBNGsLjf6A++3nXdGAmifiB8w/eTqkSBmlLxCWvM4+WEK
WiDj3F9a5vgG7JolL759YWQoBPcoYKQ0QakSZNsTo3caFBHyOJP3RAgYzvIVq/nJ
eyjrBLCYoSuUrTfFrfJ3i8p+1ee29B1K9AakGxSsbsDS+D4Izl9TUU2FMKiCOZiX
HrOJ67MMydqKWs9Wmu9kDUp2MjhIyTKvljbUVvZ3jWqXH1JRIDzp9wHgZ/wKZwOD
LOt4NhMBng58c9QI/g8oXasY2HWzmf2AkAkFMm/tpjRcpIoWGrmuMetlW5TM2vJw
CefOGvJhACLKwjF+jYML51zviOHXwQ/8RzIB49QTDwLA7qOUs/JkWGK6CLcTh37d
Zc9mbYWWSBRamEcx0oqTPejFoUbMlBo9gqJIlJb1G3lQ0GMInnFODneGttVaMfap
SMxrnFyHlLzGe+K+QAhlnFLzHEcRi04oh1ITq0ZlLajUtMrg6XrfH6EyKpDf2nqP
pgtwHuhGT61PX1gBwkofBqBLa5u0ElnWdgB9DDBcftoWRGn68/xqxOH4V8AaNB+O
zKNxql1LqN9r/Wm63GMpmCGBAELZjhLcWDKU79sodZHgpacyd6/25crkmXtnvjuA
jLU2ZHsM30uaX0xoMfqk80IwkQxZuCdwu57QjqA2KL2Wga0QYwBjC1WGKoAxrmd2
iyVqRaF/1budWuwQ4H0q3jUAodc6fNFSgvnKUBhqdsC5HadLByqmxxZaUd/zwdp3
NeiUKKGBxF+/4tpCWDyx/cEgWsB8B0+g23jMKA51aNF+Gjr3Maov/p+zLm57dRMA
n55W+Y+2wedaBkJpm2V8A7zEi1vaWy6ngGqhMYr6u9MSe2YZ+sCflmCb94e+uU3G
Ptoj7PWgNYxxGg6sPTiLS/XtomSyxXfRcLK7aiWbmDtdVb0Gi91UVYaQpqR9C1H7
xnL41B+RUHuBqhNX5Z933OQYGS71rg/X/3wfP2gCWTA+x7bTYWaLEKlnLXDcXBf+
bfBrRO6GQq8DPOAjMXLRGatHjMGEkWTMisdfka5JgQKlBTOo4msrGzHjbo3BQrHS
K8eP8D6M9O0zjRctfDYu7Cfww6vurztQShw0u2sGbE3LV6TyDVpg/4T1GEY3KvLJ
ZaoyGgm+o5VwybDS1bq65YoCoKO61bWkVW2aKXWLAEQKd/tyctumGUvenMzf+qpO
QWaGg6CbRqt1VBdpAheDuttag4uyeXWf0gMUdQPBbkIMBIxMXvHv5twUF6XbqFHe
7Mp4J7yskmlWExC7alsqQwUJojKE73T+i3FplFkK4tt4L0X0/OyJV66xHyly+1eG
HiK1dSbzxcHukJ3yAzFSeWyBD260juUeWHpyKvCsFcH2/9nd6rHAANdjf14cN9jy
mnMyqDUn9K5sghZfAvDR+G25sMp4estW2QlsPuwjdkvdJPG0JKucsLm7d62UGJaf
M3dtTMy4hADiKmmoZ4uRoobT6mzIeU1ccO5ACzJVYD7U/170otWVeKZuJf77NqMj
VcxhtUWCjeX0Nc7LX/hwMszutAy/TRTecTEn7wniut5acPCI1vZIUjDH5lYz9eSH
DzYH5sWNnIc3nksopU/TOsUvPKNjxGbzxSnRoDXe1766Hu+v+E38jVRSfYlRxIMA
VUW18r+98cjUXewt1wW3cNajENln5n3HkxB5wr/JY135cK7nJYqto2IAPNusdR/K
3mTCeP3W9ys5XOiQWvNRd9RKhR/INtxMqIkWqav8ZJeSTXBdLKOJXs/VXx6SwQQi
3svNKKdX204+66oAQEss7yAXY6JAKrCsPMNm5BlaTp5h/BNFosxS3iLVT9guWROs
hStSr7n8C1S3fs7RzQCk+LtfLdgGVYQmGd0pdxyk2WN7yU7l08ajcoWLqYQcVOYS
xBvMX7YThHqqSyPa8JBY65bWprsZJvjyTzuyERA0kz4Jozu1BBGszBT1awWn+RNB
ex0vr9KQJ7foPFdZUjtasLbqX/PMpBSIjBUZFoz3Y4A1KmCDSxgQGxA9//gW7+FK
2H5Ad6J18gymGHWZUq93RUwBGXxu5fZs9LIz5+5xK2U+NpNSU0i+6RZNMwqDHGp1
mjWZLzVS9Sm6rtgcectQBT32uZSyaiD4aWghY8oskDkOYTn6AGTuIDDlG7TZiTGn
Cj+a1yhc2AiBCmyuAzlW94iUBAubEbtrFE54rY1zIoP3aiKqrxdZm2g3DRKOIW8b
5z4b2J5efiOgSpW4iKb/JBNACZmnmyn2+iR1DZtreoOXcieNfEKVBjhWOoXs4F27
W8IdlQH2ct3fk+6J9BONU3H5ByWNQanz/VNNqXQLpwpExxsXC0qcvqChRzhnYpue
kscF2rjEM2N+FE859u5Bk3y6+gP9y0nZsgGh4IXbagxH5ZA2J0FPIM0s1OKkVscU
O06qiJGxuGdPt3gGoOZPtpYhJQ5cI+ligoop4E5W2kxXz72katRGUohExSVgMDua
NMrBgvgcE1ffmsPq2brhNjLztNoCQCgp1CUuiv6l/9KeCj6QdavBTzhM2wTzXLUR
1kqBty1RiiqcFDxaXpg2m0E62hTLbpljM/fKUlcivplaYJ28w/fyFCxh8LuCF7Lt
k1sZHZ6oEOc5RcKisf/PQud6WaIoWrRdB4cEEzp2xgEvHwgqcSfadudRv2SDCYXL
aUPpwlVBwrM8HNtGVNwKspIo66FP9Vxoty+sG/P+O83AP5NyM/0j91POj+QD5l02
AkkwcYlZd+s2i2iLbUV5Q7fSdRxou5zeG1n+b4dniL2IIwfeHRBwgwPz7x8/DmlD
5onXt3n5cV+v+mRRMQpXmv8VClSNzS5BvqFjp2G639fBCr3PJHYkecJUCkGuvb99
ZmX4ShfUMh1TMBNNX64q4a8ZE/Dova0zTxxNnhyPFWZ9hA4Qp+/cI9qNr6l7eu0Y
36PBLTLCLa1/hKbW0OfZpfVhMn3QACqQlU45YA7g4IGY2O6PuGhPUXq1iGxSf6Nc
DvQJvw79tPuhH8eJrrD9bBepBVzIgDPkDZgUc87xKdB/GBScfP/cFI77z9bu0mCn
2/K87L6jXbNcD8fVybrd8pn1jxl9XxJHoVcEB1TmQuRQxDMgQIFzlexYhZdWfJPP
qvJ08SaLGpX3OXsR8fQenLH+vprk58EXGMUP+FgWUkCfQZmTReJs/Ba2Ov+tPJ9d
lP6RiHKXEPcUvbuC+JUSzj/xmyx9T6C9W5oAFgeqQiPti7pdqWxY/KTW6BjTIjTi
Xv+2/CBqamimuy4lYwRY6AThIZSD1pKd0LYn/lVcsc+ESlolPvbt7NzSDTAom0Jx
xfS5JhEB/9LbDtq6Xp3ZvRGgdMsmY40GcOzAoau9voz7ugH3O6mRzmayAnikAZDu
yFey6li+svMuYG///QwOlseCWK5fXoa6z+M2aq3AKFfgcwVcZq6+Vvw8PkWRDMKp
82VXTj6vwPT/T8R4gvDb3Qah8gjw+XK/lpskB0VVYR+hec2fOZ2q/RGyKr2kiVVO
oBGqtbjHR0fWICu47UMdtYxEvw6F7w5fqtMAxsVLiIwzP/klVOSNcPW7BTWdMk+h
z+L2M51X7pgJNUrb8KHSl7D4ThDbXzIh+F+JxvqHRfwJo+cSPF+zAP3KcAcyYK2r
qf67/S8kauxloLK+XIWPO5Sc7uyr9cCtX7xt7vG7LHZKXX2NFWveL0BUSuQFWIB1
IJ7poQGOiZGzI3ycBjW99yLrx2rRxCbsgDrPJOYgqjPEZXFzhPOcNAY5+za2PTTx
wWQy0kAlNLVHoEH5DpsPnmsEQU8WX3cX2aJAzE3Yf8Uuts0wSufRC0QchQmfPilQ
3HenJqxBiBqO/i8wwxKLO2b3Pd8fVokMP8a469dAO75iqLQCaTYcZcggUQ8aZ5Dm
B4qT+Y2PhzIzO2B4W61MzmqxBjBuSIFpDX+FL7dcSMU0XyydpL+SenwnXFpaS480
7IlcCekVjgPNnUMAZDYAro/Tow3o5+aMviEX9rVZ4/a3Vz0+nOqI8AqiDN38E522
ESNXBGUp/5yXbALMdB8w05xKJTSOHt+FZ7AWYGibOO8Ss1lEVvMI+V1hTfUE/lqy
9cXxXTMshQ5e29E/O9Emypr5ez6pvoIXHcf3YaYxv9plREA0lid5RfiEQD2x2mI6
x4v9F2A/6FOBfCWPtS1zLwGODKU0nokINBVFvZyezhQEF9JclyPJE+iI9JT8KBSf
yWoEEZ4GZQR2CYPQjoX1FgZ2dmNgR4jyRDIItoY/OSbDDf1X7Hf52HNqXOeR8t/c
NJY7iFPIvlyzUaoy9MMMzVg3WQjNdt3l75zb25fAmm180krZdH5xMLHq1fMYHOPY
Q9LbtD/hS1EtAzSnO/reudCYAspoTl6BVcFrdEBRadFd5AwYvo0x/DV4vNPrpyV4
jscjJfYKZCxicD0RbK/D7XtkFCAdRDHCPMAsdE81dfUkZ7HgF/EbW/7/LAV9e3hQ
KWNtguVE+dakw+9rqEAe+i0xhWX1ZZRQAqLeR/HlSWJ8VN/7/tROECMAXAGrY0cR
No1lKvii6T1ZuEKs+jMhf8ma3XmIgu63sAwClVVMdRNTfJSzuPCK3SsltZsmA93W
vjnJkEtCS3gqvx3oXATKbN+gmzdj2TmnA3GfOpjZH8OVU14dw4vjEsz4JKnls8Dr
WBWKTlf1ENCPuuP/TpayWtouPpflsaiF+htawKW5wjGCMBx8UbmKiQVW9dkE7ubN
UcX7/qfkznwrwUwUets92VYQkFjnVguWC7xqetjqrRbk2mo40fjv5NcMA6aq33QY
lmY/PBj4QueDKYhrUBWUokKS5D9xeWrY8IlXYlEhiLWNuXnJ+uB56dGwXk3Cz9MT
zV3wyhXxEj3TmSuMc4QjBVPFEfLrFEm01Uk5vd6Oal9yf4Zni6HGlZkLquDT9TZc
P4Bu9t+XSD24Cd/4zk13fXtG9/xC/PMsmsoquajsjzFANUkJVEUUdVNr4Swlqutg
r/yQ7rgJlyE5AqrCQtIYAHiix9pGJbaiUP+hp7oftujWJeWO/Yw7g7Y9FObhChfC
jgyjo6yx33VwsE3afBn40vXIuSSLsyWeG1k6z869csPiypHWeFfLqXJLHYL0pjxF
kD1STExRn1LzwvhsYARt9nO0NsKc8xxH1F1ta/uFNM0DZRVt3tiUSpmpmQKocZIb
MW3mcycZ26DRYFRkH1BaDur64MzihOwa19+bAOsfGzOSS2P4z0YXiO1dhpi3OAs+
pRLtfj7BTUwp5EKcJPDIY2tsoj3wS8j2SzAtKJ6vEWoEDU7nPKnN9dL9lSlMe4uH
nclwiBFWe6p90GoMuu6JHgdGGdZiUfR6ntzyOu71dYPlbqqnYHZP9qs3StW02D9T
/hd6bIaZ1SDEi54DC/xaOYVxk1dfxv2E5PX1LXqZSvvHW8MpIM1NQHt9QjKagW5I
XYuGqQS4cTAxV5/2vWF1Vm1makFBx4hm5N12dH1u2DwKCfXaRq7psp+QqC/sEkv7
UbXXkLjIepCWMZurra9mPKzxjvhiao23HbXjEm2q2oMOt7ARa66TWuKgjnjSEdOy
doLxPCxbX8tcjPLoysSM1vHoJ/c87TOtRxLaSwlBhjFhYDHsZQFIlm2uCA5VTgCp
1SjMIL7BHwSauwzctVy35S2Zn8e9PozW9lHp8z5ghgwbmnRtBr3A6fFThjvt6Hsd
cJHIBBMvbAwF5wtB7c531vSXTCLjvBTKkfM3wCqanN41IoXcx4iISSlLCV/jNeMH
R/+JFuiiOo0XfK9MPBcRYblpTQ509bFtTS8bbIaJK6UC3Ni/76UixM/l952Guv1T
EFKElFyKJ90NQn5PPxQOm/W4ytftGu41hEdcGmDMfWKb0hSmsLWunB7dFLC+Z+wo
nDq5gq49ACVm95VO3A4IUB1mC3wDw/dJJ2dUtUjHFi5cMq6PA5AH5YLTSX0PGpHg
kn9KUKAhKdCFKLRxhbtTpAYE03rWssJFNYmepxcq2hxGQHMVyJ5emsixsfiWLUZi
91A3vpXnEGxfXZtks9/eiYbWFgS/kzCSLylNHjvYyGW5PerB8LQEoVpOofVJdasi
e2iJBLBpHEEQqtvdgQleN4uSILM23FV/luAvBfbZJoZY3RyUsc80ugSKP1eL2SUI
2G2xRNaRv82w+cS5CjsHLuQffmGzpEb1pmEMc9Xd7FKLBDV8WWFPoyDPELRCowLy
qEy2h93cJ4of7Jz2KgkPMNlgKs2//7608QRTyJ6ILNdsj4bbeS31VQsUsVtsGM7M
2n3pNMwiJ6+PVx870S5FcNVp6xfqzsichcv6BnVmOd+qRsn2IlgiX2Kw7vtSwbLs
qGhrzqPGkcTnzFKQMyRDnlzsc1of8EGQQYz48S8i4R2asGYcSsZEYbl87xWjf9No
Rmcpew7k7qcY12NGsDHBB/rtMZLEvyqPDianbR3po6T/lYeZxziuSYRaQX4YYFzH
1VeBmyQsqosYwIquNeaTeGZ7rBTevdItQiKWWPf/2FzWJmKuJd1X6R533L8ekdu/
zlKmCF65PJBM+aLtlDXEXKDu4hcsBEQacGdEvrM3rbNIzwfXopQudWjW62TR6QJK
I+LxCMNjw/lGt817UxI+wiWbCxlCxdDhSzuXajlazX/hAOWAM9zhbPoiMmLSR4cV
CemB2RBDgZ94Kz7rTKoQVSd0q1FkM5K9KQRkYu5HMJWyzu/6+vRM1FgzTdYxHB9e
zT/1s4c47+Krarjv1mz9X4AzP/ThHVfuWEd+7PTTqb0RinaRnbOBHijh49b0bYav
4QmeewlF/DdjE/0yqpq5+yUbteFpCD6Pg9GZtTNLsiDQBccJQjqWnlGxW2RPMWAE
IJQipX0O7jwTSjWfVd1DEtwXS05Yt9pgAvdFw/zIP6Za/amHBipegR9G6VtRGgaD
V68hz9TXtyNtwnHOzvb8ugsKjh/QQTbhLQnzavul30p8/CUMuM0wK8Lo1uonxiv4
273IoB7LsXCyxf1zmzvuG2ctLpQx7xc2edEdrb4goWmTqmieZ7/JwbjCCRKKt4Gj
1gEZw7+t9filV9qBstwtCQSB4NLTVXO2WkoLecsYS7Hm/PsJScE9Sa1QLkzt+ybK
PbNvgZsFlsP7bhNTn9Z5SeeIxBpAfkpTNOI0FqASFBmfXBZ1jJazvy1IbaY+LGa8
QspkDaXtn3kvAle3BK5Zj5+2/T40niIRPRGq/HqeM8JW+jZosdchiu8mVME1ozoC
q8FL2XuUTipuzYM8LH6vmyreYblrJvi5aFmFzWGb9j7ste2rD5o5q6lSoy/Nnxg0
ozweub0FQ1nfwHxiu+FNg0o6nW/jY9xDIKWBxIhoP5VsqYsbTfXrI1/Gi66MtBX/
2oM8ymCYwp+0g9AxkZyULU858qFAQL4o7qODnSxjuTIqDCSSm/VvY5Es1hoSj+TV
rNDfYvwqyjZKjdRJPJnHBKr00tVe04r2bSxn9ohBf34VZj1WGCoBX6+EyvAJ2qcF
faNyIBr51AKmwp+LM1RrAo5+8LFruezNUfpoOM6Gf2MzA9NdaUbmL/JxeZVMkSIe
dmvTXIxlJbONnJ+vYm0ZSCPZlRQZzbNmaJV6pSlgb5HVPYEEkBzpfFnEmSNjjOhh
td3sEHdAZtz8AMXrkwohEihiUEK9N3aCxKtGf9fp3Jkdj8guxBqShCan7PqI+15h
NYXqZ7QAW214OwK/3I7zW8XMRZuAzQoJi67OTLplNpEWLCEPLoKVRGWovX0vsVQp
EuJdcYRhRn5BTeXf4a9q2576BH8mhseQJbVyngstJpXO+gHdYdkqd6CxPfPdfqKa
F8PQUP+Gg2PX9T/0cMRHJ8kkQFywImimxusrEL0Qz6EqNahuoQ8GG9waRt3kFF4x
utD2TCiUBdYUuhPq/0a0upqKnFPwukD/elBg0e78jSgw0fHe2/VXIu3AOSAtFMsk
0wyMPS5tkPgXbcXQc5yr4H04WozStl9FYZ5/8l928ibkU7fl6jeEANwGwAiV79HC
gaBy8cFhvRWFzjr38+wbK7OCXEeec7UHj7STq2/ZxX3piNazEPRXbzwpfUbnCOmz
G8MEy2EoGdVrDoC963NGkmPxsZEAGXFV7ezmbaEG+JtctyDWlX+maOhaRsXKmrX/
TUfyxjmjFYsXSjjSI9BHoUMIDCyp470d+FIk0dyBzU6NCRt0QEUWX93gPbSBvmeK
2xiZmWYbpMBdWRq9trpxMObYzR7heDE0KCnk0lwtRyTW67kDBQ1Y5oHhEwW10qYx
EfoZcYyteVFQRyOzHgff0QKgqdUZeyetwrnpkHJbACRjEjZstBb/gqNGuuwUBYC3
GGV8RYBdKjySoto41IZc5ArckHNmdSeeeURCT80RHO3l7LHhOVyCRZAe/oqBJS40
lFOhepKz1FQZ3bshPUt3zphWVICfS1d/OT7sUTLTu3G8Z1TajSnMgHH7ROwLmguX
XDWyrf6X/34rvUKulshgfA1aqtSsYKBJ/IwTTHYQlCSUnUD7FVGv2wfjcrCtEwnZ
wbJC0HVKvBaiY65aZrWqwdzCryJYJ7qKE5jwOE4K6AAj6PYcn8kdxBjSnlTY49J9
g9Ko/dF389/NB/0ItxkL/c6npYSLzBLxXMOZ9yRlorqc1hsmWmHUzG8bd9VY+MbR
bbdkq56s+THI1i+IVji9k/qk876bvg7ExrK5yXeVa1YmaIrUJB5DYACZiVImafq+
BE0sZeYQRIV5Cn5bk+13+aMNE0psRlJTJsIWmuQd/Y0XeLgUAmMJIWe1vzIlVoXV
3AJz3s956gfgcV1LgHavR+UTcoKwa+pl07PhnSa6X2/psL1fULkuRJf3RfM7CuLb
gO4MJQl8eAi0m9kNqiN7Occ7bf+mWLwQ0sFEVNq3s0Xou1N23/nFmBzssMhZbSxV
wKU9+xRxhebBXsRGLvmpJOkgfHFtOXBSzywimdlGWUhmqRsTe+wDFZpu0LyYZK5r
ZLwfw8Ba1dbh0tPLAZFqZSruWIjU3GC6brfUHMVGVXQQCOAOMcdGggfoOFbelTjI
KIlGTI+wURXsgzHQEL2L0xM8D+FFrq6RorR1DaOZ8QpODP1q1cTV/dbGS2W3wWan
ULyamTsyByAZ5dMXt6qv7hSa+7O4OeVvP7Bb65IUWxdOxvK1bpu9jvEK1Sw5ypFn
+x9wxcOFQGwmC63I3pjB75tLKJ6bMdyHbF3FiP05uswR6yquWUoijVu8G7j6CMDQ
NbSMd184AaQ7VrMFNKwJ86hrXF2DI3w2T6xUNm3Pk5l6y76TXsSSV7yekMy3REuh
FB1THjm1IqMs3QR8vDCUrHOmS4wnVV8zbSVQSGPpbmVMW4WB5ZVT+907ACKWVyFH
xbkqwJNCk1MKUD1KZc/SxTcs+n5NYybIrqzWA7lYJTK3fxw3aNN9OJSOs8f+LdPj
pX07rDixbKp0B128C3P8ZJZnP8jvjn9tZO+e7SHfdjgWTmbTzzhF+y5rcf3fD96c
X+bMLppN1J7PxEk7f2TW9JJYSdzmJsfaBLXVr+T/IcD94ld28dXVon+6xY+9cnL6
s5n87hzPvsIEs6d3NyQAOizhQRG+cqfMrNBLMwLIER6ZVyXAMh6uirfroYtf3Gcr
/x7Hudyw0UXTGyL1TggDzm5FpZQiEQEn43q2QLp/Z2KhaXqIjiIxOgZ8Gm7bzkJr
9kVBDFuyPpkTy0GOqy1jzZKmup8LW6E3X4ZknRx25ba/EKk2MH8EgWjTZLVZXKK8
++J9E5rhx4ikcfowDNF/YwMaeAQG9POFwbN74eQQ+FacQuB+Prb9hWFPQgxG+Pdk
tS8A4iVGUapeXFhz9Tss3q6KBidDzuI5dMdmKkJJeELg1oWV2wEJ2IBdzmXZN13W
MHN3KrvuNI2tQkOPl50+3MHsFJ2QuumiDawcs90uwQzhxeYAgnD8B7gSDnPRjMku
boqmW1k9850o/vELoZtnnuWvEFPwlXqXKMif6/L3eIBird63e7G4aYoC9+WJ2gLa
WgQbpWdKS+e38VQbeCpQgmOu9WtdPLnreignozqzb8LO9aRIv9wfpVhidhGzm1J3
xlhPAuL6Dvxe2v/oPZz6Zx3zOTn8N5Xe8asBkYW3d60ora4nFCp5fg0bgaUqxvP2
R38HB7xbpZZ05ZRfxTFI0qHBFI7iruCRpJe479uYDw4iO83vVF6imMMuCL0NS8oX
mNvDBbEgeSQiH/A04RMyhSUO8ncVgzl7cBxOAwmC32X/j1KLjCckJy5PvTZzGTAZ
eOfm7w3F4uTNAxWwYydo8P6Fsm5h4MQxt4IW1ZUbBdzqz3Y5cxj24Q+e8c4MPHt2
0vvTYCYsWSjt+SSHO9yPAQkKPoFLE8XIxQ8UNfqLiB50WJ1Gx8Ckm8lUsHP3ook2
ChG8wJ5mrNMqBa+BEvf7jYGyrOZkwTeotYxaiUvfUYiVCRHjuly3QC/Jj7OFoOY1
hmFU3GQxqluwbbX5TnsI9edWeZjT1wrXEzgKOLymoqTgW8Rogz5dmGhupunJeD1W
0WuJldKdgoo3RX3TaBVozUk7CTZflPB+QtNLfGSNXkdEaZq3UdmlXSEaMBzKIb/7
6LvLvnywmIRdQOCDErdaJCY5Bepxxc2eaD1epyBfoANmzFTNdWKQ79P3u8SOn/rH
gPQ1ORBYkSlCqIlYUsx9R3Fqzm7R3y65gBj1v5An1RvDQyk1Uw//g/CXRn3mX0cW
0ExNPLO17WTlfiRbNOC71XxAs8hS8DGeWPg4LHZTz8d5Vhr4fOxQ+0Aporyo3/nI
aYOtjweXdIMSuH0TdLHNNh3gzWxNBlGOfH7pQutEm3YrPNo22U2q7Gofi+GiP2pt
lttZguYi6ozf16Rk7ds4ldg/FiZo1x2nGWDLLozGWix89eyGJEjZUsi4slsakkSw
eWcIjsuyfMxDjmQtdKL9szB6fGw2OXHp8jjKnDEg63LS7q/MAw3SFf1XG5VqIE65
Ol0BV+VFW2+cGAYkbp4W6Bh65yiqWqQAwXk1DEeh0rLAfNHa57sOu+7W1U7u0/Vb
iF7i9EE0IRrTZmQTHKE3ppImlgFcHPO++plQpnIr8v91/57W0iFQyzI9tzzUZj4k
4YNzpIsQMR8YgbWrnVFHtSlC6WMuoQBpyHkbMqEA0peLk7DGJAleu7be0ozdGoAL
viPQkUpv0Q8jIcT2iQz2/cMGz6E9vM6vuEn1F0lhGwAVRc164bTLEoO3NtoQD5i5
cBafZwHsz4naVVwxanxqAeydkBQAdzQfHUtwD6ysjGtD097tyRCA2foLu7myry3K
0WvaR4LCPikXcL6coPutzlOJavLvHjtYlY9yVN9yXjjGwdq1zJ5VmU9v/QUnelzx
8CXBdyKW0vEx7CqEZbPJoOKWwsJq8mdVAj9nsDYflGoXHqg3JCKF3OHFCA8pCDnp
+LElI4ji8OiUVR8WfVRId1okqOcydZdFuLkLeJFEiCVYkF2NNDJ0n8+qeht5/1lq
aTnMoZ8a0c1YQQg/xiURoQNPQ+jzEwyMKDByPaHFn7GMK4UvYP5CLEzXdB3J7k7/
3J+rdQkvdHOUpM6qiZnEA6W7LMf2c6MWmmn6T8FIUFZyXYs80vsKpR12v+QPdu2d
GI4kEg33xoBYvPv6uLU4Dv8/vsmDtRm72+apfp+MvC6pKzZs5iRGZt0zrWxRc2k1
ATA1AichlT4YYUsXU6th8do40s0QN/mg0URKw0RE0XlEuOIUh7smcrHPsHDXPM/8
Hd4PZQwdS95tfilWgQl9NsIg3Mcbgj6/KsEQHMW2cl233DjzpTxvlimHNOd3Vgsh
QBDgK55Kii6+7d0kzwlpMJzLxbKgeIiIfxkUif8oOSo6eXANmh/CPj+BBorR+VPZ
5oV2XuzpSIQT1ry554pVLiXxvLHajpV29S6AZWpBxzT0OUl9tok5XfDIWL90KiD2
k5NHflI0/SX9+zzQT9xx9SlkCnicwsramIXsvySkCS52Ex+eY90UF/XRHJv2Ppeu
a+mag3Lvz2I2IHEvyailzbEFdyOaKBoBRBqvl2WuUx2esAmhoYeroYvoaOYiyOwC
cwh7+CQAi0K+9CiS8cczuGJ50+rLa3JLF4ux11/mN5G76Wid0VEGCd1wEzfbUOzn
Pu8He/KdKWMEhYVAfZo88bFvZzxCFV3n+dqdWFSx/pyzbP8myl8L+zBTd2F55K8s
ag8yDJEybuZDbwEuu33bI05dIFg7w/U4GRRo3wRAuWGpYsXRLFrhGd6A/t3pMd7f
pvW6BWsHdbgyJThZJ9a/Jzks+8lA/Eij+ZValKWKfkFFia9si4rTx4D55fp3sd2H
GxDakru9awHX/u/yO1rjPPXPnN0x0atjy2y8xKKw91/mLcxxOo+MM3o+QEh2oM0q
gwv7/yP0W6wrAHm1WvANPAUOLrPHCzfaIcyqwJPcId/oJzHO8hRwtthpW5zawYu/
cHplAWXdZQvh4LM2UUQpDMwZcANmmodlOFo51gMAeXCzpcVEp3a+kuWmHfMGj6hI
QgOA0enN/P3V/minN6kgTo9b0RS0wS1bYamK2Rr1ZyYqcda6SO+8b31Y8Jwoz5oL
Ts5/b4OoIjHvOb3mVzMrYFWl9BSaUYCr0TdRD2nBkTHvTb6gYGaNSY5WHJ2VLsbJ
fUjoBdcJiXtf/pSVAB9GhWjsa7sG1OUyu/I6V59i0vUcB7FuRsFhclyrDvm66p6R
7Asu/rhEzvaHyX0Korxxz+dcGVVTtCEnEVudeVtgQsFGlZATwyQ7NUgIKYxxZo5a
1kVZ0ZCgiLOKMssaD2YYNcWhS0QMGEkr2vopODRMhApb0DqgtfQNIyALqibgNLcC
KwvtQCBmdINkPDa7S1Q9n1f9ulCSAIrBXW4OcMuidJVwDdQ2I8I0B1A1qvutB9oO
yX85s1FLDAIcMU+tPLa78RrInGq4xzEuzuNy7xZbF35Hon4r+yAuADGUq3xnuu/v
5eh53FpmcYJbxAlFF4HR4DVV8I/3rDNAQioii0iNazDdajxtQFKewFhxFu8Xu0DU
ZkxMu1J0L0VRbmTlT1QRR4tHYiwtAJhjpaOKXbJvIgyyuxA5OQx3ksTKiDWTQSkk
34nAN339miTFyp0JorlbJ6Z0ipYzVEsa7tJZ7Mnnf9LdXNH2KVsniN+tnz+mAgsc
r3QYd93Ur67Fo8czs21/KgGL+rmWAnTYhb5iV44Xrp/K1OF14CtSjKJ3oIxnETym
0C3M9O1WMovfkd280HrLayonISvYtj2rEoirV65cIkcE593VoLj0cifxx9TTUmft
myo9ZcQYnAawEQoLCBITqgtNFYqSEfpHhVFdACWELgWQ/Juho5JXbQ+e7VmJfg85
TcStwxHw8N3XsuuATshmMU6VwvRCwdw/1RLyGLn7GP+OkbzRZW53IkuNIKxdUgEv
vXgIll3Po2D0PBcaUyajsjQRSPBFuNIsnC/JTQ+PNI+2XW8mX6dknnsArf9BAq65
LWyyr0b/f6pEXSaCWEBsV9mUrs3ezT50IVehg5dHr9pTMt2btan61pFdCreNVSLd
awysOgDiHQMMK2cfbEDSvkc1ScarC1qu+MixIorIHyrz1r+xhZJT6WX/AG+Lbx7v
35RkmtjrjNz7fIQ107gb6kXefy/OuXTtqLToJq+W2ZLjHRTNGYTL2wRRsSYwYJig
SR7SpT24pR5KXmbuhzWqVUB4U8+25OwCZ3tAdFwPiheK7ydEsctdRx5BcMaxpX5n
+U6Ico1kc+DNbhcFiNOXXDPXMgIeccQ4WqO/YWQi5R4jbKrSTpgmtuXDm5gNJh2K
2pCr6JHkl+QNkiaRVhGeo6wTBhJHdXsA8G6VYnd/6srWKf5DQc0DJ9w90oEyD6lJ
Z38HOUibhz5sIg94i6i7EEpc2PXuZk+syh3Ke+ZRqJmhQstaAVuZSxFBC+q2FMNt
QBnO5YUi+cn8TokmKh5juO221yy9TYJr1FLHJ7sdRtzaEy+c5Dv0pVGxiplbn+l5
zaJj7f7K/XJuwrdjk5/O+qxUET2aVHqiqlWX/DnwLebwpKghOR52xzE9XPMUmyum
r9Uf/2Dg+favSvLhZ6Qj4mKb8XkJaDs3mqiM07hKXsD00+IlV0edu7x/BT3k45Ud
nIpez+5QnVjGGRFxkW5YlqwvJ4KNzEQcCWz92aTXS8/p9M4qz/RbYzcktKgGxVTE
l7ydan72zDhEPDAxYuFSf8Ck6WD04iOOvQUbf+GdrEiAUYUAd6ahwTsW6wposz7H
wqloImDlV96X48iukAnnwafkrk0seEb87ioRpqcyic7MvLj0UPKdenMfiLeQyJfu
M/aRvukNcRLyijW+keor628mMi3C1KkY3W9505zetsYsLOmtQxwmqKPGtKZc+++r
DiWOcMsmjXLV66Np4/cP1fFRHG1hNsNs2E1o75u+RQlZuCQavfB+DWGr9CgaARS8
n5Z0DyxsYbvO09bCjrYHjb1SWfpvBckX5hk1C6j3+1a2eRIbmyxfay2AevtF4pO/
UQq49uN/GpaVwBGyjIcH5t96+NhxFj7TVJo1xbOroaPG1UkBCk3NV9OUCK+SwMXV
V87Ei8RJOWybXb5kR/o433YttGeFVaoTDMXFqqrs9x5AmZvov+penCcPMYGguE+S
PKtJ1nrorSh59QvU0DwiqEEIgIkqR/cUqK5G4jyvRtBZxu4VWPFigE9rF4odt8ms
ZkK7jGPJBEg7ed+dPlQm3x3Mk3a0fTKzt9UjV0p878PA57ytbPlNFpG1483jmTpL
bdA7FS3y0UBkNrum0pIY0eh45BnX/P7htBa67LkOYQqAPV4LBGn7fHjldZhRYQGc
P98iPCHJKZBcdg5eFUdyfAMAEUzWEeiEi6yVzwSg8qZCUh0mt7UtLKqVZwvJU7l/
jINGuRATiUoojUCsz4uIpojaE5SvjqzNSuDkMXTB8Nib0dYUK3Gxthvyel5MRsRt
C2l3AGjTWcIE5HI4oYXznSKbSikk4aGgYnyOutQJXkw5vE1DPfAopV0cJGlFDSa+
XTchR0XHOK38fO84yNdUR0M9ZYdK0obmXgCY9b+BsVwP0gtSBFpJEe7bGRp9t8Aw
2m0Tru05GyJDA3LZHLi83ge0WT6rAXsRQt4AZki8XUqHadvD7SIjQFjSeHjv7Ec5
7jIG7xnam1gJSGWE0inuzHUVYwRz7WAI/VOoSHRmcf/orgL6wSKVy3koIdu4NcHb
d8fjByLskgjjZxO1X+5jl2UJktD3ubIfY7Bls6/0ZFkv/DPY3UUEeMOHRZ1U6SUm
kawspAwB095jEb0kQrhb2bjC2EhAxrYwFIcW+wJOLZoSdgMd/q2O+k6iV6XBhfpV
p6EiRjpdjnck6efaLbmatx+Ig21FfgLqR/iDexF6txtPv9/p8hzES1kJ21keTH7D
V7pOTbQiHQtSVoX4Cwkx8tNHtFjCwP2ngLVfGyMoYO0QIFgxLZruQGs0Pxo9djBW
8fHCkXT6nfUsVFoHvDDIRF8n8lKA0B37GkQt4tYT2d5Yje8+ivHh0Uh0cs1cdx4w
dQAOWUbJuzxbOhXlRbWlz3dZZRnYtA20UdF+lHDvPLUZ7ECxYw7/5+XjKjbsooWm
wmQgniLyNBTvobRfF0cxQlv4G4bpperynkOSaby7I+1Q2BmwxIciyD7Rnk70kORP
N+s1yk+Nc9rB6yycvxDnQ8uL6PVB364Yr1p+hcVRzNhnsO2siaLRRP2HONvkUcLL
xm4JxepZO85rnnG6wIE1occrJ4sueGPt4oVd3JOuWES8LTleen/PnPoTxT7mn74r
4GU/2fxZE6PC8up+OiVnm/qC2fQIEb+SKCnznoKntkxGramr5iAod1XSygWvwwie
HT3dqG7QaaRZM6RsNa3DjT5dsnk+iYtysgCAMaCeirpVn54iOc8U8lFad+cW3JwI
gy3DsAMKj4zsGXbmvoUEyO+aFWlTAi6Cn+Vn6k1XWxt0WCLy0y7FdtDXO426KFBh
3D+5HEML3TYe84HLs1lbAcivX4uRVZWtZlhAND1TAX4p+pcdb+XqyjbHHWmldIZD
IzCFy21U2L55yXXevwsdwTQJETvIP9H0WqyOl4s10Fjv9WyKfcOOvkcEGwl0LP/J
IukrTCUyofaUDwLUw7ygX45cwd4dP7xgPouwHR4szi+MOKOwo7NgmD7HPjVGrWFe
t+u/OVb0XS/hPDc71MLJkBEHLJgTE99PnjAw8SiJfw0OlpN2feb+8DaZ/NltWEhI
XJZojUV237Q0fpUyypExOHJQroc6Wp1Ms1Yrs+H8ol0ZbsOjbc/UuGAJzV/8gwNI
9BGfHXfjivt1dXW8vSYCmk6F/9cX6umn2APsdlHrFFVInmdGWeFDGcS/JEhC0dLZ
7pyR+dE7JazcQuvukfrCHbs73tcrPJMrHXpPiBI1HXMHcsFacGsbJ/wKTRkCJL+J
V9e342U1Pn+GI8RscWRnKFizLS8xqLVNeGPuAS37QlbUwMoGMSkxuQlVfVBZ9Gi8
SQE4Gw2iVZPzRNflEROpXWhCoS3kkE+muAIbBiAQC2CrdTrM9GeYlJknHbnObBcX
dIvbVrLPvNjgVZQYv0kLKhuY3w7ewOFuywQvAKwR59WNZjDsDFOTPTiGM8ZpnxSG
jHYOsQChlp5Q/dYFLd16pfc4SHcvb64+/2AbaOZZ5JK6r7rwqpypFnZynKNp9yCw
leh3ZalilNd+yc6O17Q3clFWoUfCpJQQ+he7TQS0FKnManmseE3QSy/J7VkEDMB/
+j2fciXPOmH/xa6rkNhEyQrYGMmkE+KqDedBJeiXWti3QGeZrMEgqXbpGDYCLL0L
ULZg9D3x7Pgl/ABtAzRFFWZGfjZLPiGstudI5Mh0QHSfYBAQTNJFtAWb4kMO9m+c
LBEbn3H4ury8l8wy/mbRxyztZDmItsnBWASaar9UZjtVL8osbEyRRKRuFmV4QvM4
XkQnIuX7AwSImVDPL0sHEIySLxbXuQk5L7Y/WNy7FlZEbdr8zJMpcTguzhKRv8YB
gqN1OgDcM6euhdo4xUB91Ru+n7+nl1qVzr0idF49/xDUSmh1yGgFw6E3/BVbCMVw
haonQxufFUg1gDGIKrji0XhSSDxZ08w7jnFI56MLC2XnA6O6YGNBguOtwjtTEbCT
unr8ZvnRKCUxbsB84mOIbOj1JLIT6Q10oc96DutNvo7dNC8Qo294oc3JtdeScavH
yUd2DaXEmjkoSsnpTM+j4aIGEtRLmYdpaLFvI0Rz4jh7pGy4/EdYsoMQZ1sXLVC2
Gz3dgmOOd+t0jdfq3ZAPkuEDsldcUCzmLUIap9xcqP9+AJvcaGORAynRfF0DcNte
WIC4QkD8VBNH/M5JI+QTodYm2h61Z0IT6msqC1g8g5pQB5LjpzpwKDihNQ6Xb5/P
DrBegnWEesJVHtON5YeGf15nv1/QFzB51PsGTvvhL5pWdmvNSEA6GpH2/RY5+Bu8
WBDttsj18wcUzQDfjnzcBU2qeDkOoTglO4UjiCnjVTaCYT6vuXvNZ4i0x/Ud8Z1K
oOpUX4UirStP8F7di8vANFjQcxE33U1friLlPWK0uyC76XYf6TgK8lVrSAc6nm/l
9MyFmVTVmAfYa71FNVn8s3N+b/HGYYAXu8Tmd690ZD6UzA5ISItjk9wxCSc7Tb+K
GF+wZbj6ve8XiT8KkaZ0dEBWKr1tRagownRAu30PQ4tOO89YddUM5Vm3oVFOKFgK
vEEUlTYG25G87C/+EAdjiVdzXIr6lohFzdU5AV91V82q/yk06meiNt4FBPi/AeNi
AZydaaZF7q3iI8n4qYqEluncJDKs5t02HEuJi0lBxtUVHT54X5Qu/GU2MeQt4jzc
bj6ahSVxrYevcl2UXAgxnPVCmmmhhyC1OGz/TlXePUJvdzmkojwI4vjEXpuyndbR
AKbMYZx32RQXp4DfWwr3L8dO2R7MLWh0/+0gKvLdVkFprHqJB7CIiUW11QLqaWNe
XRh+Fi0kZHo/rtU/28T7r8vFAHXoNZ6fD/EA3GT3KTClNipwCA9iO922hmlOCo5a
8tlV/OnM0X3rfcGUZ5klIDymqedRWjIpLl7ODiI1kL4FIpztXCKOYlH/5OSzTY7c
B9XZqgX4oHZrPmzzShSkTEXo/fe+TUe9sNaD3HEMF1WyfzWH/+6SX+Qoduw1xr+3
bDH7ZR61jQ+vGsFxDWiAlM3ahrrd7BkRdgfosYEq41ZgF5O7ET6Ws9P5GfeUAzPc
DOi7ZFN6JFN4u2p3YPcJ6HjWmmPYkC6MYwlXjoaDkJgPZYtVvaacWlGJ5ffPySdf
s6EE15wLosJ6Pmu9+XpIESDmvgv0fdyq1IElZ4lkUwgnkOTnilCbQ6tNEz6O0UMN
zssx7gRbTUW56tS7B8pDc7aNosKLFI89caj+ZhSkGXfJZq6AafYNcQZGrXBQgULY
l7bRAMHuBmKeDIhipaWXCNoZ5pLEdLl/uyIHRGawh1pNfqpOYLvAFUMmitLUUrNl
oJdvlxnK/mO75b8KjfBjRN4kayIJZzqvCVuXFtGEsiWOkfcu8vl18Ny34Wge2jls
CRZyJYzENrvKrBLtUgjHR8kv/wWOGae8kpPM5f8a3qWylfxOJakIKXRM5Dhhb5kf
cXetrz+z0X4dzwYaZAV5ItzdQXN4EqnBN7EmiZGprioExOSO7c61h7KXeGAIdMYd
h2AKBjFigQIqbkHVFZIB8nVdf3ZwyXEIS09DZzKJN7TiGVOQKS5Visl787xsETsU
wh2QLFsSf7yeykLV6wO++EJzaZNUjaYi5qTxpwNc+TqweQiJhwTuE+410YKrXQ44
o+6a3E7FPfopky4TV2ur9crVji+QjlO3b2kQdzocvv4EtQl1pviPcNswmjzxv0SI
VDqNqKGJAyCNwqw59HcmLLQZj++LCsX/Q7yob40/F+/3RyBqrU0HWOxjLtF0S0sc
onj14llzjKCBxt7bbI55Y/nPWfK+ABzx1PT7GFAFI4tyExCnBkvzA0ACqeTIpcfD
ndQX/CQ99tSAji2TUutphPLavg6wsxG/BML6YQS3FRFWY4/cFVBxdZhRoQKpGSnF
h1gS+1ODnwCsakPo0tgHMETgO8/LbPAb+VX88q+Kc2EiEoMdJeToNBu9Z26s2Ghp
gn2OP2fbAQecEi6k83B06wevgxXnvPmJxV0me1sKh9LRC56hIwy5kxRD9bgAjvh8
aZEJTjSpy2HU7gJ5/mlcyw0ywbOWbDN66boxp1kda2wYWyx1NYicQQWinM8Vec3y
4yhR9nICbvpqKJuTjwkQMr/ariW/tRoW81+yHhqFGVTVrdx4MpbTNVN9Z+IPdsRp
6vcMzURWF/hoEVLVWdlqnXP/Gc9dLpTVtzk3R8kt2ZMwXDsoEYHXSDw6JGWmYlZo
9IwWpS7xPoLWyRpgoRlDRYFdDLEL4Cuxq1ilRDyDChAkHMwBKPEcFG4QayPlbQUd
D4Fs4I8vymgt67ZmvDksUkLNCWisBbuAlzd4Otoqt42vkTtmOdh+ob+8J9D15fTb
T+Z88Lc4QOif3KM1WToCJfx/DtVQ519E7Me8bt/GaMDmQF34sYg3yN9z+VRn/9Jc
Q1BHQ+PpFenBDAp7G+CyowpwLsdjZxOuQUr1wcCUiuYQiQnUkZZ2s6jNvQr/8CAh
qbscSjQ3tBCy0mxZSYWKI/ECMsKW/fgcbF427d7HZXR14l+CweoWDN/O1oMmTueT
yxn0oqWzV8leqyhXXy4vnWuGliqUpVLOGKUSUBys/cViDyE5OYKYtRghAZni9m3+
yxOGmN5jpZGCfpvIkzmX5xux1HCqO+CV1CgtPgHjjT3lPuxBuEw6NsnQL8Gdm0FR
FOiPf3QNOSPUOkuVPCRk8YUlI+m1f1W+YuRvlIdDUIhsATKQ3SPeZkmIJMlGBIkE
qANBuD4eeYVPMP5yoqN9hhlMK6XMEWaSzY5flOap9cWDL7gNMNMKOvUCwgjp/Tbv
y49hiQLUHIanKvl3VH/li/XlfSqRyR0gWkuds0wxyuJ2KeCyWabC3c/iZxG36XzP
DS5Fd75iwUFTcXOpPkk2/ijOBP6ElZOzMqqxVX6sKK1Jolem74lG4+zsiHFeTG1G
sXrQ3ce9OKxE6IkM26QuEcpq3VYbvLkV6LoTwrTpSJZxMB5s3Nb1q24BHJqAVg5K
xipe/ICu04PftCMhl9i+u0ppOdKPYu8ku+IU15XVsXw1iLnWFtCtFS4Hgti37c4Z
IlE4kyuI3wiCs9AXoWR4o0NL/xDFw6gDXHje/rgDvx5dYJPFN8zRtcRH88aEci9i
dF2t5nIo1cXY96Kf/kmr9yUesBlAhr635RaJKIfZqlUoB+g33tVDzNbG5tV09c7T
GO7bezpYq1g+ilHA5i+NUTkIzajzwoXFuKtLiVDD7xDUGkShRN8a7W6GHRVyrJ36
3WKqR0H7BNb/2BsbgPHEbJEWaf32HklDxN10HYPiW+UixqNgU7cz3LZFoMS1r8Ar
IvpCRTpdK2vvMnEvZXwxPar+su4q94vH97LwOvj4RbK0L7efaumRIxZMPDtTlN00
Odndb6I7ezbFcN7EBlFZTPY9X2fd1dxbnW7jHkeWEwKyo0bQXh2+GF4/pcH9oUZD
Akw/LvGCku0kUkHVsXE5MoOJuj3wruggkeXFhxCn5+4dop2BEHLjHxPcRGL6zSgw
AHxMUPnkiDSFXZgOA1wWa8z58lqoiU83jVJ/mNSqay6kMGwB7P2KAi+NUJdHU3ak
phKbRe/+lEpiY5rj9fnNn6xch5haBGOllMp9hNx9FKrkaQQPsXEcg5sJoay7TXMq
MgkX2vi0qSMGuwR56jhFqB8x2Nb5ATe+/8kaVMCXSTyt1hCy5QIcxyGb3NRQpM32
nonW59GAslmKyEpBOdaAROeeBfABNgUmFp5c7EcsGbe4ahkTUQ8T3NZ7O0Od3hP2
NiPNdorv2v04PdVQCWKEWwTYhSO7+lynNetOQ72H8AZXpI6k2SmB6CbmFrymvGBm
YyAp0f3Re4MGigsyASmQW1UC2JDq5M3u2mgkWptxbKX1dmU1sdjgw5v5q8vtBllr
0pAijKnjZEv+5iYiDKJjrFIay/BYfE4NVYXrQs5nrrMHqAcOBMtbZHoc4GE0JXH8
PVTw6nEBOwxude0fjwBy/Oz/DhDQqVdnMxoIyb+J1muGrkcRutXLX1LWtp4jKHZ8
+eeakuHOK47lFvKNp6O2QyHUaBkNdOAcql0Gxn0y6SgOlIxHO/jUDBJj2ygxoL/v
JtbfwgJvecZbdq4xSTBHCLg5kbq9Iofwaio7jXqRW3aNBRV8WXL7t2lI9yuk1tul
iENb8KVlfs8pDvyigZQytf5HIdzUHtuDVWo5f0nDjZ5O2o08bZI5ZSJ5HPpRB07c
z9s9rma8NFl1GF040ut5tAGRM3cqG8c5UcSCaOXOLnt24FQskqsPX0BtY9wKIPGI
hZziaLwL/GsTR6iT61lMAtDug1XXaoNInUfanO+3GO/1NSKONAPeMmXfSh4FxlCx
ru2cQekF55eZzfLfZULtulr4EDSJTZ78wQpofeBCn2u64PUp6CGpVO4t9d/c1Zy8
HmFpMbwa/1TMZpCc7ghRiWfxRT2hGTJrzxHyJ06A1YVokXjxUIqEa9GTkOV/2Mq7
CPTpzsSpdP7rzRD1u3eUlmzepqckCWkXmJrcDilIyDuJTgsc1hdDOXg2g1mGAsac
Ek+AGRgQTDYW51EA+pobxvDzXwr8ZbHbPqxjl1di1djwGYr4zfT8KqHp7PgUXAWm
krpittAO7y88oM59l4+YUlRRbEgDd7+URf5Ct+35OFBz7B66UpliBsO07wlLYju7
egOeSd8xGwjwzI54jH7joEr/z/6BvVTVRFrWWBf1trRoSFJWi6sDlx8zih/H/zCX
J+F2i/YZBqnoA1P6nj3QFihzZjU/CwgY5a8i+k+sIuCKcHnY1a8nx9y7oaTJEoFu
c9jNWgOWNdyaVgQ8k50yIiM1fDPtyK+qcU6hFPK+0/Si9/IJQF79rZtPTLDa+EuL
/4aHcN2jdGYh2NkGoKuqpQxOAFDF6Fr4oiF2vbG1LJkAO0TZkMtGhhVvOk5kS2hP
7vWaj6Nd7FFXhTzDK73oIl2T38+hAHFAesSCV9xO6q2kpIwRcXu8JZS9KrFbzRe5
W6JD6pSPcLKJNb4ytiBWu7sk1JaDPVvt+3zJsbNGBMgAznam4+HTYE18wpJMHrOO
0PfuE6Uxhipn6g2UwXa++/k6RmTWJHRgCdgarzUsqoxph/yYL5DuZ9bFRGk+FPPi
PSzQmiPaDhYzAp5NkLrRW/Ne6NJu0sxSJ8nIVZvaklKc3+yNO5PeAmG9BucDJzX3
ETk4Jq/HKNCNvQd2bUl7d61/8WPrdTWoeONudWhUzGi3yHgHiUgsrmqt19NWaZjl
co5m9FD1AP9CvdL0dI6p7j+nLepDXFPcU38z0UrHdnzQQROGSKQ+L1al5CD4dVWf
4jEi9dZ86yVBKV8nQnTackSNkB/eT2gTAPXsLzN5Jypm7vnGFFOz7ZTzFYe5R04g
VmDgnM4vneKzmJ1ueCPU1DM+7ptWI6kE6CaqTCz1D35830901kaTcUzq/PFBogtg
yao4Y+53wK262EsBs+Dw60x3hG6rT9dmvwyXjHkmUCxI2LyI2fsoS1cxZ5lsZVN1
tDqR3agK0jN3jjpjydwjM7SklIm4KwL3ndz0mQ9LCMHwo0FJLRKTApe8gWMCspBN
GWouA1ulifiT7c2PtsHXEZnWbWXxb9cDW7POrojZjofwTPa08ffjFeg0h2kSDlWE
tcfnHH8mUIAXXCyG+FasW2M4QlmWCOEWaD6GdbGbGUVWbvPRuwZhavQ8sC+0Fc7X
Gd6to9oSRL4IOKAc76KPRAbMGr9zMpurf2RnwOZDg/y0AK9CViVpRYLNydBJthZX
ssihQ/7l7w184M2s1sS7uTkWPGIUsmE1cUkVC0XkYBPcMYiCS/gzcfvyIPjCXFg8
hT1MVvj8U34pPaoATlwlUOBAS0MYiQoEMSKdC+gejTtEWS1leMuhlR001CjaD2Du
K2rQXIg+vPReQNm1BMomPKpFBM3GlQh+vcZmjGp5QdLVnFedLFkRY3hToTto83LZ
j0w0kCETsJnja1sXsxBqSnKVRyvNMsKVxBOj92JILWPFp/2+360tJ10HNmFNUfqs
s9vigY5CShx9yISVreKDZTbd6GFEYLuRDxo5nC/3lqCXARd97jFNd8iA29vF0Q+K
xHZYd8aW63KTDrV5WMpiyU67+IZyPt49fCgY8J4SXenftGlzvuceE04J5x0ag0tc
SsBHSebv2znGfVqxEN472MsugDf9IApTab8ztZfFWRhZTpL+qbpLbPcqD3FKChGB
SahKjvdaYdqm9swnQwbCGSQigyWCeyqsL9yNGU7c7TtNLE966KVbQIg+rU7XDEip
oBmahR+fnEYAJc1See49s7T6yEYq/m3BFz16iocMPPubUzLn/Njw0iDoGpPcb2d+
MNaAbh/lRb+mw3WX0gxs8VIf06TE/CT1iMHYEdNdL9dDukAUA/MlGxnJdOrkT3Jf
EA/S0MfqSYz4q3Lq73hG2wrlf5vTvqVB41+lyA7Loe8msgPkU2ObjzzYXWXVGxk7
FDULeGi0zbLZeN9uOCqtdI/3mIJFEFKuqJIGAtqAAy3+wyHs1NhGmW4RWjfUhDhp
PUWvXFUaO2uF/EwKvRzXo9bL0c7eNejrjx7M3YQBbwa7Yhy6eWg55BwwuvYLYRNw
KehgYVtoVOu+ENQdhfRchmNAizCYqTMgzfmpMYGW3UqAji8oSR7UX8nEfFsL5zO5
hgsWFuf6m31+OX90okOuACjJXpy9V5UlyhbNxBGXZzp8CJPQ0X1/vyatG4oVmOLr
KdC/el9693qK2I2ZZ84JN8dy9iE6TKdl/5SloKl/TjVylrEy1zjwxoBVcbjLQNAa
iXYSx5Fvo0os5C3BvChnBD9fUvuquo8ImdKBn7ppbspE0apnszw40ejCmtRUl7tU
s22Jcs0Ss3QXxJlB1G4SQvlrRtsRm4ukOLkdRnqHp1v2bXmmmhKU2s5FzOLMdT6e
TTy/05cgb3SFNVdAW6/+W3SKiKOAm2sES6zMqUUyvPzfbvieHQvyOaL8wmLG/FMM
z6qUxK2GI2oBlFr0Ug8Va4Uq808sifwM7B5CZMdVGKp+uWa92vL/0naoSPd4Mpy/
SqmLzDzro0wq2Hi2eeq9PlW25RZVfs9Jn/3hKXzVks56pmmJhe6ub5EdJDtHDtSW
+tYnYRReYfmV58vr1fDi3VxZczoEGgKKGrzNiRvV/74j68InvKEUtNypUUzHY+bL
8q+dz30lrbuBfCp/zXwuyGPILbDH9Av5sAjEHsvLwux5dsldYYmNGkKHADdR1Iun
9xQsG59DYu+oUPkHLVjvEiT7E4GTYp8jFNCLFyl2zG2UqsR5wtqMJEIVMJwA1IW+
LpGawhDcmoHYZtzcweSvoSFoBCI6Y1zytqep1N01Cnj6JJINVz2idMDSUbny3XgO
gYziFAhSJDTLAN4u3CDkc3nOYlse62YFjIG3tVDN0mTnBe64WJ8Uu8XmBecr8DgP
XgDtBxEkbvJTN9w6wQ2M99pKExby38P1Jr1IOsjpiUe1sPEgYEVxKDh12prbLsHR
irOYD90VZzl4oH5JkB5XY+bx4WiesLsXW6uI+wedWi+3f6Gxdqt7qMI4aEz/whhl
QweXPvqQ69HQhhv1okCtj+28gt2A3k2pYxJKxxdIgagrq3s8EcXEHX+RLM/NAbK9
iwzN6GWODKaXgfWqysg5fLjAwZUIixQek1bMxQxCFsMsxQmUx5dZm7Z+Y3guGqAh
aJ2MTjDVIrcCsvpFkeLwLvwVcPxPYwAiDZ/+O9Z8F2xvYTLt7smdJweRDGQeBCSu
597I0W67NDcESaBnkyObSIxcM45tDlppYkvDbWEzBlzYe6ebBbz2ufH2IrcEO35V
Ajr73j9aSpqu4VjS+hF6T/SNyvfASkPwgZzLpSRkbKJaF5RscrUMTo4jtWBMCju2
doPlp6u7+R8n6XunU2/0UnqQDi23nOu1/OVxD3DRzXvX5zcn2Tqj8zsIoV0ihAeX
CjAw4rF9AwjI9/UJgOAZBsqmnzkjIGMTLm7yWwmz7CjB7Bsil5f0bwHpg97RsVfp
R8v8hR7meK4F8p9Hvi0mYxsj1LMI0VjMuf2GvlKU1uB05j5kbapOGfblcSerJJKx
5UXXtZU1Co/oe/anfOOrIOupLmlqPNIFCnKEkGVA7GDRpnk5ihviUdJPwijdFfKX
83z2dGXQNIeUQja4IWRTUDuc/1xP4+vcWNcA62je+UPcXpaN7mEcKe2ZtPkFXiDv
Qlkfa1oX2CZHNljybKiWZPsMCmCvXTlMCmHto5g9SQxDsR1zpRe/lyeb02C2Aimn
y7VZTMJholNO+9deqrJJHbMRSLh2gC3PAruH0rKmwLivAlUtv6adoZboWoWx/K1C
PI4wmCpoJQA//iO2fQxK1Vjpa+oSUAoPPvvPap2x+2YOorO3A26ywXRovnYtUXSQ
zLUmBINKR5k5wgQtW/0wXEhvFwWVxq6WHV3iHzkZP9NnND8asSKVTPPvU0PeRzKc
5WhGNeTt+AcDGKu0EjhIlZYS+cYWe6CmVqLyrvMqN3CZFCoRjFrcNGGyAnGy8QwB
OH4NdejH2279kjAVhPZYZ0Wq4ZsdFPe98dlH7XAVFS1kbtxS8HQIkP36kLuYr10K
lYcGjIw4F7KoAktC9oQ2HmvNa7IBlYO372KY7uOF493LviEiATK/KCJkisYmIz8t
IXIm+FpikuvJ3VB4pQ1X2JBlmrRO85VvOZNaQacyJr4z7MNBP6Q2LiUVqIbUbJyy
ZoVwQuoFr/cQdarpVmfPBDTDGnhQbiyTD3i9Kx1dFtpY20CX0GNOt4y3QD9MqfTP
JdfDQ9ToMXBfurElAQpoh2kfYxVaH/snNMskCkiWLbPahNuVr/qgpRyg75C+y31L
sEHQAhugBkVQhGNVFqQsfGkPI3cNESBj1zPeW2jP98Pbq5P7SPtOSQ7BsVZubKeS
ULqu21UJegy8iacv0Z2puxJiwJA/d9UjHl7vPZdSfVZCerKKvy4D7cEymjQrMdus
btypKRJJ+pVNHwCqGwM4GZMykbID+1jPMYBsDKXUhKKjIQ5SVX4JK5a9sgKuPq1X
NnatShXfdJmg0LD7Y3DiDJxWN1Npjy9YpMkam+8Rxfgxd+XXIuRFgbYhVLylIsIZ
2DcHMa0wYdJZ0JRXgEK126w/J0L+N6JLtHib5W6VbUv+T9jbZjV7lddW3B75O1uq
GJrn0gH80o15EmP+KOwGh8cpMutoc0SXTNU8gk3yXcd08TGJSiVDFmpCA+fG82TK
SJ7eNBPxPHycZy3FXPJMv+AZcMFrIPp9BjGWjEMmhtXLlf5inIVxaIo/U38XdsR2
UJtKd3kgq5758kRLlIPy3x5Uss0/WhDnOZNdQFc7OZkUBTNfzc0N8P0ICapocPwH
VIpO2UT9RORbw3oHLYUhcTYx1+AWjzS4J3O7TEK4WZlmC7bJXUdQG8VxEuUYN0Ph
xFnrQEeh51Jz3FBqzP0uiUjwdz/bk4FYKsIqg9TZkHeirtv/Z5rBw6PdOcPpBeOA
8EHyDgZbC0E8UTTd2wNHmB88vPQCQYwS4xSOTuU9OeYx7QXq2hGSXOGWnXi18vwh
z9Y1Nr6m3QFnKRLES1XsExnYknfCWWdp1EnmJjkKAnuL2RXjXJpFFwi8xdsSNysl
rDGYV9IIDAeP+SrQt64NUWSTQGP2kBvsbQG4oXYlGPNJt3QJ2IvOAxA0jAQ9lPCl
b7VgJnDLVk+4rG44MrOJGgUZtFFtMOrDcCoKkKOJdqkWVG0cZwXyA5ij+HWYglIe
cfszZnPBfiQ6XXS1eQLjo1BMmG0zuqZfMFCGxWCYPdzbepy2oN/FavxH4kYiocMR
clWRF89HPOTs4tWozo2Dg8yq1Q060sZeOGbB2xxDBc1+eg+tRmLJ3WI3oCrDUIfY
5El2Bd/kfE1ZK3LSEoLrySz5Hnc9hcFFyLI602skCi0WAg16InY5P+0/9bTLfmd3
wwXJeHL7x/8IpnMCdBXsP4qvSzaGOKPJWNpvowqfO2v1aaEUmbPIVE/6nSVDIKwI
ytkKl3P63P/jfbh3YgMP55keVu7lrXQPwzzvy9pez2S5sm4+Y4Y/TdKC5fvgXVy5
0iFJ2y0GUVYDi08CK/sI2h1raAMTq4sRohvTpvUaajTWEu7o4IbzLtId51P8QVOJ
mm9bpisDEXzzLlPXKE318RX6FMd+tnPutChUyS6FK3KxnmnyLSESwtRLrGK7clIH
EHLEzk90TcufDSPfE3ZhWVcfutzJqbD1DOVyDpmGL5vsckitutPU1ItD7LBlLYAo
sgx1qyIwYLhvI/m8ENlZQoofpKmlr+ETWcitWk1lJIlcEDR4vkDq24+QQBEjVVFd
q/g3uRCWwNHlVC6XuyDyP7GWXGPgwB2msnpXtTDngIxBxK64AsEezPHaKmNMDRzw
QCjIisGic+sJA20i0lgBCcGnDCaM2G2jD7l0GDi+vB5SDra02/aXJv6VlMFaTtXs
XwGiZF/c8S4/27w0AGvglRkSIFh/QTTD7tkOR9dhfMbKtnSjkfQowCsxR1dQxEdh
RaShQ9AFKDK+T+HUuxCQA/Ge8/rGm5lO6bKc8DXL7rQPdB8SNogJSLwxsO0/N+V3
1k/jxSVMxwhdqz9KwijbvZ284k++9eBSCFhIFroZSNKLfqbBqoUSm5f8sn68JfpC
qiEayt5uhSKcn4/G/qfCQ8NU18Vx5a0hK08HaJajFpa+6WlTjGNYPJqlF1PxGSRj
vKa0htZMtP7mB8oSz8VOugUh4CmlzA3Lr0Unc8EzdHKO2/B8YzBf6Lktfo4cUJqO
jw+TOOj6kabsX+BloF+Z9PY1WwRd6ZBYoDDoQj9LlDN8en6flzEjIGIaOXHd7jHn
cJPZ6+kLSqALGQzYX5azaef4VwMtp/w6ep4aPMz5/HQp5LOrca0q/il6+gF/Kr7g
uEHbzntEi9Ix0zHVK/6yycoECA1hQOCMwgaQwQA0XY9kSwhCgnkriK7VckvfPbZg
37MCAe8qw5m6pJJUJZq6U+wob30MIGGo8ubr54b0Xc0yDrdg14m4S/fOaj7AAVx0
6E3td8iYraI64DUYBbA0EGSfh1pdfY8d/sy2Et40rk7eg4Jl0p49NerC2Q4cnxA8
IjYu2fn53WChgoO6pnnyTgIG7vA83TofqbURi1b+n0XiL9hD/RpXUAgAzlA4Bo8l
xR8bqeRf+qhVMdRQLL65+XMxjEUnF0wa2StGdb0gX7NNNunWZjgxak6mOpNsrH4F
KVChNOdty/tQHV/qkVsfvrwlSBEZ2QNN6cHuPY8Z1WM3MbfCYC2AyJKppDKtfNwP
m69ihWhwJTktmvHMfXgD/IQfbcFfvqpd1GHWVVxAGzcOPJxlcQg+iqHXIfm6hG3C
jX/YBt8KGxV5uGLDX7lgjpJjhAbAeBTtBv8RuiRL1lqc+bDsPTsk67yQLb5VCko+
vrMaM3JJNkJQEVT4J1AYn0fdX5FqflBofx1gHGDTnLDOwkk1CLVFo2GzrJ7XizII
HcHJXH5IZmXoIrEElEsPhx0DijNEyx7JJ5W+jo1BEA4wfz1nci9PdPThjsvj2Ti3
q1xpPXWaOJeiNs4ZSTo+QAUf1g3s0sfVNK06rycElpbYwtIwntswfRIQDWytc0p0
yOl/6/uexheiTHMFZqwj4L5KFEGQN2iKqm8LRSsnCB6wEGhdGo02ov/FsyzYf3r3
EG3VqhPC0y94uY5Ghx8ZP0ffSLYyEYPv02iVFpLA+M9/Ulk2ew5vr9tyEGOtTf2E
UUHJEI5qhWg9g00WWzKoMTAFZwtpJRgs3DkVwg8R4yobi58PUNUYwOcli5ViH420
yH1S4UEAEMX7Q+1g3SoeiIs4qLQF/fCVI0OnJz5oZ1GolALKJRp5kLYW4iGTG3An
7NstDTRDEh50IhbRm9TufI1y89UhNuCQspe6MpMseqTKFjlEsVUiEgdQrTFz+TkL
DJWL9XGcmIfO9M38T4LO9cE/uS2+BcDO4wZ2PKJ7gvxR+mwhbmD+PW5gHzJXt70a
TD+behABPmI6NnWyx+SL2Mx7EYOVo28mRMDl5snVQ3TKAPg4u6D0OfIz8fuOsBK/
qIrMlas1G+zupSCBZqRh06KmUMmuBNnzVfgjHpsO0iCpmTECG69z6hB4A0BS+Ivg
VnBA7LP+vNzxAU1tt4TzGI1G+17SVdbILByH791Nxr7O2xGshySJHa2vRyspBx4t
xz4VaDy3gS3nRPFKK3dW48DqrvSnNpH2GN5BRRISiK8zDMB4w8CnRHh/MHZ5lC1r
9BcF3YTBKenWt/sO/UcEG9OPYueWdz0bNueYRVUQUnPgXCsDveybuws+56sZhQmZ
6j4zWxFSTTMfJViE2G7TIlrrBdh6BbMYIoMxJ04tzdqgQoBssOHB5u5iWh26XRaM
dRwnfumnTkwQxkX1pzFMkTcQbunOoNxv0fqHMHBNc4pkQ94rsveGspzNPNWxnAZH
blsPE/jcE4HtAX1t+3xSD2AFMz+c56vTgJXrzreoQwosnuvC9FeDCNtkE3V2+Z/X
5NEZaBDJraI9Xzb3U14u+3qyXnLWyLcxvb647gLopp6NJ74tSb6G4oOAr4Szd8A8
5frMaFHKn9Uv5UryrdoDlqoogIWq/YuBLHpBEFeozkrj7rVeQc81ojkYblFwLaz5
4UHZo1O0sgajRodVcrbPPSckGyxC5fmUzX8PJdBqfWr8MrLxZPQ7PF7hiGYcYgzy
vHzeclT+NDWEvokyrZovJ00dqJfiDhGqgiiP9m4Dyz5++1qMVb0J9mEf79/Q6Rqb
Zfcu3KquaX/I4wHR1ZN9WH/5C/6uRslOYASAxg6MYGCJz4fLyK8EyJC0i3lopSXG
ZCGespUVR3Ho3JCjOUrvwXX3pO3iEiWczYwyBpJ4SQDgNplfS8IVy1jmhrFNpgjJ
/A5vpND9iJmHN0Jk7zeUNt1j4NjPCCgWWpCIjrjMM15GubzHede4qyZAadO8tqih
XUlTZjLQoV7bPnOjvaac4z/k6ml7nFld9mITMmKLrSUvN2QT13awojBe1nvcckVU
8uiz5fWcFJK4QXcYqURnrN29sLhELj8085c1JQdTw6PaNuV5+ZnR6/egZgh+4PRl
4waGNUe6DSQf5ivIZWHQ6BW4vKCYkhM6CVNPb255/yQrxfUmIDyCRB+QT1OMMYH4
wkgfcBRmZBR+v1URSz52pGm3DpawDqx8WUEwVSTmrgQezIEeZksPrVk1QNV/n1zm
uM8PI45yN74zbBDwe6vw3zw491qjZA7iRIlG2G7JpqSVTK8JiJ+1ovmkubz3mdOO
fw/MNHUaH1tpGFPH6DfUPdhDamnmrHAOL3S3/z18L1RZN8bh29tnNDmCqEcaXj8L
KPKEje+fgY/awP347r/K2FGy7czs/l/xuviw6kOjIFNJFhoVHBIn7T2Y8LKVSpkY
IaVHP0YtvE4FfBvGVu+V6T886LSE/bomd8nZklzMZrNfaZwsUO36m3uCCZRcaJt2
dipoPm9BRyFREAafAVooYXbURRDsUPy+DDX8oi2gww9It21usTfGNmYr5kjNJ3/M
l+YEJPWzI/rXOUbSmd9SV8OGRJSdFeL5yu+eAPTndjyWf/li+NHTfQw7H6v2xvoL
W3l9A5tuqb/X/E6y6u6uQCfEsfga6pVM0+u4XRr6Jb6v2n/P7jKNG56RbrISVFx+
sY2BoIlsvqzdLF/36Av9iavtdsqhoiBRdkVEHKN72CqzMrXVHmwhdQAKLWnIwkmW
x3S6wrc9ezekWO/bSeZftNNkErCajrLK92rcfPz5uuhW66XvItepbSaOkEhnqrQF
maVzoGF6YcP4Cfkw1GExJsqpOsGCjWAjnyyASuUtpBcqooYM+wxT8eRp548yere+
hEMmhZ4YzqwVeeET20qBT2pvUqSnzH+CkW+RV/+s0+xwu2YMrw4gZkKlSlp8WCdL
ABmGGh+2BN3dVvCHzth0G+7mltijV16DwtHvbKIJvlJWuRrPUej/u4/i70Ty9KPa
EqQLc5a+P11xBF4Rc9syFGjtGScUE7DLlwcVIPLzKDX695XBVOF7k+3kkkKO2jsa
TOpAeNm4EySOcHlvC5cIrctu5Vf6z5GGLGc1UtBWfm1nWX5ACMVO/C4Ex8cp1r8Z
+/I0QoklekEXqUbSy+0PfoAUC09g13Az7q9OIeIa9fNcF5xkTXJzCt4jkw5pPnT9
inxwQpk8ZEgmvLyU2FOwGW0CwBL6w8qvReEisIKqds0uq84RxlmXaGCo3x9TyX/4
X3lyWAb6Maa0EdqjUPC9PGWE6een0mX8G4ntBNOvHgY6suCVb7/d1DTqbnNliCUm
aParFyLxWnq3ZZNendVyulfFXCjsLuH4nvZQQt5kD5MTfGBIa2iyQA5r3H3XPhBQ
IaGeKQnTZPMz3wTx2eYjh1vi3Ezz5lAJoMg8UBd48vcOyoRWeQIwDKD/zdRMK/5z
q9JnemMvEG+cXvel1cggBBvpBPwq3LnpuZ9BZTHWF2VIjpVla6gLpu1ZaX0IK/bg
ipcwhDHKhRWfO8GEMgAMqvDK0asxQ8nj2ACjhYj6Lc4bBkMiW8d64n91Sl1IoxCH
wzCk6v6cI4cLboyr/eNcg7JkJjgwfX/5x3+Wnglkh4dCH99cvpZMyLYG/74BilCa
PzCuSh0m7Kvrf7nbIjOoKt9zckisJsiQep3EXvrse2LaD91d3II/v20SKcSnJCwg
75z9EYLsPVBQ65KZB+RJ4i9t+N9jYO+qhf26kUtUFXMLsvsLUFDZsBSh8V7OdYgN
0P7gU2S9C3dND3dtK/q02S59TpWUSwxnbBwa3yGykwITumlAqr4mdyCBK3omdAIU
qsfWGQTP0frJ9KuISEdtB1uEGvjri1GdkUXjmh2j/vrJEpNMlHTpZyL1sD7ywk4G
cl9WXHu8GqOJdpMLAAzKysOtufIb4uD4qwvEXNCh/UqmV6vbr2g3qCBZxaJHuwlE
amgf3b1E7oIHK22/FI1OQ3nIpNrfInXfbnS9ajxxd5xTDZsaumOLGtZIvQTSr9DH
9WbwW+zCrVpcAUKH1S53T+0bJfgAjspAd+1F2dZQY/L1iG7Wz8j7Pk6drDi7A7Hu
+W/wq3tlDWSIl2mmDKMHYh1OBgC6HsCyyLWscl1TFWqLvIAsOeo2o1gouGfl3PmZ
WKGIidd5IpF04ALkiT879wFbBlMXudy9LmkOzc2TAgFY3fQFH+VpAToLUqnnzXEd
W1TgoLFnj8KpLVx1lz2H3ibhqvM/beOEBHN6idfbfeOAL0XdnL46figQObasLkO8
WOt30Lcuvb5Vs7x+rZtvLRhNoHHvDiShl2pfhkbZlRL9hog65r1HX7tJSWCUj1se
bM+sTVoVXnziKbiQcCClPPobGD5SyE1OMrJLArwJHTKXidQNPQ+3nVx/BBp9ZM/K
Ym7Ja5SjkhqCWbqYa8L11500fT4KGzd8pLgt2k/WsN0TvyfkXuofr8Z4zzM1UXo4
o6Ly1hBB4fyMeCJ2zGv3DpVK9d4wNws6Mx7q1QDL5mnRpJunjP1fQ8rGDHZubyy5
dUHvHZm+wttL48I934Vbv3B2cA1evTmIafwzJsHaPmw9aaph7fXsT90o0x1X02ne
OKgSSNebhlVOYUZ+tlAU7a3V7zDNkNlp+GS7FOYNtUbIGP+yf1lXpOJ4SI/VvB8D
j/Zza5kk3pqQm8/5oZPjow1lARKhqnrcIt8Mgy214vfplkvyoSlp9eNjDei+03/I
VX2uNy1FnSPNTrpHadnv9M3pjiOIVhjA6DroYT8YSryohvOLXMtVTJUpb+b32suT
BpO7K8/oKl2uSPGX0xmOzH0VF890kdjmzfDF+e8XdkUG/YGJzqZOKafGlwHCgtOb
tfG7QvYqc6WgJ3Iwls2MACk3LO1RwQF5yZKZ3cC/ZC1O6/TIZuwx7kSMnQ3rHj27
3qxAJprdTpT1x4qufg7eFMu/6zv3A2Ta8WPq7PP7S+ryn1ysbDVYqkn9ThJVjTOi
/JH4/RaEQ4L2K9I9ugSVsHIBWsI8gjXMKDFTUFhcs7PwI+O3LSIWUnG8jUZbgjx2
vXm1/odPugQYkMrBr/m4efTDKBMD4LGy486+d7C6wIaA930Hrw+yImXGcMf/lQ2/
o3yUDjM4nvxw/JdW0wWRbOUS3EGsF7hV9vZ/1oPlhiY9dtP+36nXf3Wyq0wvOkO5
VhJ++JY40teMuEU08PqFr784J9lTosjohGQ7Ae3oGyrj+CGxdKkeGr9pCfCX4kIt
XrKPBvs9xSg4X0dKNDViD845kqODESmDfQVIbHIIVaF30BQy4iLkEAWC73lJgCL3
vf2QYs6fK+mKbxshUlDeNRRsxjzmJi/BUs2ER0FtkDc1CquK7VPlD70zhHYEOQI2
uXDUFC+nGAtMCQk06tGQn00JmqKmTrhS9v9yMCCeundt7ZTCcHREx+OZIg9iUgPf
3ShV6P2bxCI1LoHMkEksPuX7ZkgWoqdLBGE0IlNwsHGWq7D3crt0HWllTW7q25Of
CWC3yVJzxojgB+iWxRHJwzt0I6Q5ePL8Hj4Uie75xah9VEOu2Rs8leRzD+5/zE0L
fmMWA/XVMqdnL8efiChEBg+DbNClYoRcJd1LnwN0ONrqNwYyAeBmbUmAalC3wecE
KVU0uUESIbH3nyVyzhV0D6mirmJQeidg2VBQuMUgzl3+ewZoV+/xJsor/+a1PQ+G
QFEQL42yZm0DiIvzKRM8TjB0x8U0eKM016h4F2PpzsHInfU0rhgAccqunPjVVWrY
r/suNuoksCcj0om61v5C9MWxRFWThQpkJKzjkO7vhyICpXrKrjoRu8hYhX0qD713
OCx4rlixuzo271khz9dyYAv9ww42+OdkCgo7c8YIhB8ynZ1NcVJ5aWHWMHY87rqD
sLPtfkfqMUHQXOVZFurxY4hPX/uZJ489sBQSFkqgz8d+Rrq7/W94ARoNKCW9dRqm
XmhDOx4vLo+WX9LiGucBzoVg8N3ZT7kqMYJJn1ifGRRTi9eGpaoS/pE7wkbv3taI
SVGFFdE2rJNfd+6GAnRYYQmkQt3Mayxm1/iFmHZcG5Ap97ZuCyUhoCqw4J9B+GBI
eOL71XckiZYww00+1PBDC10OJ9MqvlO4/2cy0FdmJfNQz3b/4WNAVbBJ3grAbv9t
qtD5E28AazGAsDUUdvPlTo7qEOLKIMwmTzGYyjbUiSrrjCnbG69M7cjruACWMePk
waht/wnyVdZ97Pd5w0BaJwLO6R9GAthwnMmJh1f8tbpg81snfkgKS/hLE0Wcn+RB
jrGEE0oFJmxglodLV54FnxvfDyVX/aiimJtRHnL0ijF5NM3Y2wClhJVvsgfwig8L
7TFUPQiPzfzuFEbeiaWf3cFJqngvtvdPa9S0QnJkq+4GqsyJtq8SwJfhYao5QI4W
jUzq/NRAxSyxyPZP7ofrzy0wmsvbl3/Wg5t6g1x3kKWE1VtOeA/5uRiAnydu6UbZ
LUZYGA0bZSHqxPnuREv1UmSwkvr7ybbl7kJNU9uzIbhQvhtdzXEt2sEzl+xmm/jf
Iogx1gbvjkSp5FpH0J5Ov2/htbGsCCrfNQWq0U2M8YgDzrmgU33N7q1ylKsSfgKq
tEinmhJHfcd8QDgyam8GjfuWVOg3Jl+65Ff/+FoS/Fy2ncN8uqOZ2Ou1xmAatmOT
BmOl2G7gJxZBfNyzeFElHaeP5tdWK2SGAT4hc3aTF6HaFuQACnmqrudwgM+0lEUx
zD3vvGiRUJzEAnIDbLsUNXjKKdqCc+Fp5M0ofliM3tF/k9HGPfWEvbyZldrcyly2
blR3dtJObYdeLla9GlFAcwe8Y8CKqhNr9uBBHHpj/UUldhPoyM9Mx0SJJSPMpZmz
uiIuoV96mRnKLsmabKLvwXa4+sJhb/pzUSohazOF5Vh98tBRTWteB9eHBt8RE6ha
8cwEYzIGqIF6/3ZlcKW/E/KDE6n+Taj5Bcbgb1mitIvIAxJ6OL6aFU6LSQgixW8p
bZYi6rE27OWxdelQgffgZFzFgWZ8v5CQCAh5mSkVHkPI4ZPVHDe9R9w/0h1HA2UK
bkUCoFpClkLA0OsolUBqrRwJM8oDr+eJ4G2N/ZV+8meDji5Gxvo0HzSWKl8MXNuR
/F7YX3v4ZA7T9ly/VXyEPLO7AEPfwClzkOQSJe0hYkhge/wnBROKFg++oh+y6Wsr
y51BWLcGCX0mkMzcS3LFXES78Uits4kpittp+bv1ElthSNNmGUjEwlQFkt9b1RQN
i4Ov4p6rWzRAqGLIYyimU69nDaowEuqMVf+tMTLYWaCdjyBJUfCj67r52l+iSeIH
pJpxN5CVbJ3MDBAoqyL6Q2EWEMiRewclgTB7o1L6ae0VZ4u/piB3GvrAIuAKjErv
bjCj8sR/ePkCJDXS3bJZF5Yyn5IaEp7AeHOxQ+QZJ4cQHtpoV7Pp0cE1Cs+n9DMt
nTxF95p6rsRydTwjP0RFDshI2dhWJU1eo6O2u1rXyXn+lLYaT1LzwE9fJmRAKquH
i53MgSBdg5d6gOE+SYmoe5lAVlrnxUWjzkNyicK9ha4DFZ0m+SsEBpSjncofrl29
NMzbIlUT24AxJwcOmm13rgzSt2V4floyw9l5L+YdrxUWfuvxGxhcATDzFNvUTOS4
X3jqVLYqfZKXbBjJyybm0jTrSPjdpf8EpqTQ5H/3NydcRwheBYC4qDQvT2GX3tpY
4KNanG9tET4+mN8fnGYxmDJjU9uDFzwUx1nH4qYbcN16+ROEXaEaPOIV/vUHriCo
eek9+Ir8idzUXkuOkDt/SktV9UlBlII228mevNBeuhzxXXBGCJ97XdV/RkxkIm1C
cqQku2cSNqdjWWoPYOCJ3LvPx8ZSVzr0vXcK2HzsGUCb7BGHJ3ufNwoW3i2evwlR
4ujLm/tymV2aCFvIoPg9VwmdzKaIPH36N6KMJrDn11HasznMOJJ4T4MA+NVozDfk
lpA0BaBPFZ3X+Fm1vQzFqVYFsv0anQiRkmq5FTisZ7DlYvsQHpO8AprERqBaKO5b
ao28k0be6UwOfYzlr5Ttrhsahm2Q0lG6oEOnV27d2h2eAweamfEPtIFM0+oSrWJ4
J786cegi8qwQr/UXw/nZj/Di7LSmU4iawQbselidIbDr7sXMLtpbrfSS1Eb46a/X
ToGRIsbOzE73vgaoCbTWSPu/W+zxLzHdlE+uqZoZja+M/bb39oGurClIXfb5mteU
UeLhRCYmrutpCEM8TOd4nDguCc7SliHxYSiT4oYYb/e7oOy9gt5WsBC7o23oVqIn
p2oyWTJ5Knl2/ArnaBfP179PwHgW8sMz00aJa8lmXSO3o5qbCQn902t2pMWUP7gI
Ag1/h3sMrxIy1DQWXEx842xEJ5lxs5FuWTNMDJCmhxAAPBwwBwwu9AlBN5ao0noj
XaGEIT3KL77C0xFJ7KpT9fOatSHOvbNQz1idP5QidEtLE6XTLAkZYiuH6rkFOmwA
lY+wN1WJF4jk3uDtgvf1xjHc8lL75f183fECFqDsa8DIpBwwH8FLF4vzfYtbOSpQ
b6TVB+pdOkhnGU9+qUlFPLv+HMjceHJ/1eUOfgW42J2ggk6Ls7s3RwkZecr9WmtC
uaO06eXb8dVWOsMR3vnBxCwLc3FuX6OFF3ELy16USpIG0g4H+zQ+GmAma1l9s0ap
QqHXAWa/z2enhw1Jfvy3V+QmTF5by1VlC/iOvYuTPT7qPPQeSnQPvN2Wm+Pnyf/H
exg//Y3ZjnkcwuI48gYBEm1BHewEJ7isupzAIArP8uYw9xqchABXJjqOaeILYy7h
Hfh9kJWooOGLzBAJxHXng8xJwnaxfdt2mu1NT6ITNomBbRluMAMHeDkZgKuW61yb
yMooyQ/ILcrrbtyMhzvfp9oCM4vTb0YzPCAZYiPho/Xe8c0tET6gZpvRb6JUjBMz
feT7d3YASqXFEm8mInNLKss9sNaWlixKqqtKpLe6OkzA9TfQ0Iy3wzL5qkLhaXbR
7uNbj7KCwUeZi+8qdyKI4A6IC4jAmQKl96fG8Llj2S+OHzhBawCE9wwhtGhDoEui
BDADt5wKMMQ4AnYIdI2Rq06ZKT71I0c0gXXOV6gL/qEi52pETv9/pgK6T3RTsYk9
4c3ktzoWpUa27UYyYe5P5v2xhopivkBmujuKtAel8/NKcsHpLyR9ZWn7yBRXsyOA
Y6rrzbfmQZzamCf/0n7ZO+h7binLVDYRSzxsL9R8C2TgOuH6vwklpTOIcb7zuEjD
8Czf8AyJQFLHhatp5quxGhRQWuOjleYyafHRX5vbl+K/M1IBYNF38rLrbdYK/H/k
zYtTMZjwchypOWiyhKcxh80R2qziocgtURUikxPdlXMHNWBnD+kwlVM8mMv8VxIW
cNWQfnBxSdivk54jU59ovI2OMR7Ba4FHn0+URceCdvYpV5uRn0w+aOzG21nH7JRK
wTqQ6/Xb5QkvzrE2zIa0SzgOpn81z0h1dRHtZg9CIfaxO+BpSGdQaLwlkoBTXuhb
zBUZvhKmIgbVRTsaxmVY6rqtvVPNaeaB9OTN08BphtOxnR7xRovPG3VEb6Y9N0S5
3gqbSfTb3o5pMBw6ZHHOtmWoYwf+gUloqwW2J7PdOudaTRe6cVcT1+EAudmEpD+8
fFGHb3Kv4DqLVpyrNq+lt6I9f7p6bu+fT4BM1o91l7ABZgTqsF9bV9K6vRUIhM2R
gehdDMxiPh5wj6YWAUKUgyY7urZWyR/rrdfBo0n/rKOI+QQDVAukhwG5UXyVejsd
ovubjO2n6rA2IwDALIZBtx8xWMzraXS8LFcsL6YXn7uLdJ9pAnJcAtkXA2ZZYFFO
o8aS7jfNG5bAFUvvdtGuJjHDqLTyP4kWFmPtq1vDZvZEWYpAlwXhEOn2MqT1B6F9
kR8h4htwAXvQ6e6jHo+dn36/ez4FsUcTuettC/jA67F6csWjaDi23Xxb+7Cq5OCh
VssBikKjvq7FwD9PAW1ms9MoyJEpwpXcXi6POg0rOe76TfZa8Q66NNj0ploAVXG8
GVZaJQv6NALdxJU37fr/LiMi7bASbX8qB2UI2McqbnLlE0jTDj3f2+3/2Lv6uPKo
RL0G9a+T1YmKf8T8lZYNMABPHx+OjHKr8a21T0IAjrBvww5kWJDVApH3abyETIZY
opPlb4t88jCjC7k7Pz/Rw6ZoKB9ywSYNImJgHPUM711ifv4w3VXaDiWRs2EO6CII
TeaS5Ffbg9ynomGgsIrW68+Y0MAtFE59eQVRfKCII4pVHWsE3hKEHeqiX7mOUflI
3NKjOHPxBGhsHJxNRvdslvTZuyGmNzlphLQnznPL+2UmrbzmUPISL6pPf5zTdKTi
UtfFv0NQ7Ta7yZCdIYYKaLlSg+4JtfHQk0Alfr+EFPQLe+cj+bRXW513TohTRjTN
vOjtwdBV6EZerCRHf9RzUfgeW84zKkF3VBQ//9dbcVpAjJiTBy4ME4L2rpnpPXlH
4knJwl0MJSvQ+eH+ciIAxULtYVEv485IrmBskg5RB9X97Q85PcPiMCiIqn5Ei5Qi
mRGBcIw1naOJ8NoKMz0LCLgrPUYOEjjJrRfNQGw7WFcyoAeoKYpt2Mmh4ilDJ9Oe
lBJzyWMjb2RqDL+PgSjzSiPklvGUz3B/oPlFlm3xitT05pVzm7FWJywGKIvwo+vF
7QTqquQLw1wg/4w9TQkzsE1R+PFLUkLQvlLsrEzn1y5a17ZdeB6E/Qn9rHOmZd+V
JDFfwXwvBPaWhOBiMKlBDVKAoJYdsarWONhyYZe/zFg/tKFOs8Au3G6IzYWQLRM+
kVbK5SKZDL2KpkUL8O0TB0QqG/kuobuhXm+PQcfWDaWigEjcYWR6Z5v55UobYN3E
137KIC93iLYvRMhixY5tRHsHYHjb/FhQ0Mbauakyj3YqGGNjCtiLVsw2VOo/ZXH7
SPGJRco4gF+B78M9zOpXDsTvAavSCIrW/QbwqUPXXmJ6snkIhYoXqC4Tl1SP5l34
19eX312bJyQw441DpApREc4qkVCrKtU8lauf4qYYvET1mWflsFUldAB0lv7WVJ+x
hh44xGC5OvtCQqo45YzVnRH7BEldEmhhBZ6ic5bpK6EYlWpiLyOf39JvoOjAPW8h
OmKpOvmFmRo+2+Q4p7E5PtWT1OM7UZfeRWLEEHOd7KqzRFIPwD3Uk/PtNT5VCvf6
XEthBCXd+EVGQ1ZMT+DjRduHFMqmgzJ9Md3gJgOzBTOOM/p6rBR6MSgTkRix0kTu
f/p7/pgqdMIr9oiITVoKAT1/ksG4xGp2eUgHAWwa+cnmG5f0/8bXdSjB+gaFoBKm
TpYYwMskQSE0F1C/D6/Rfp1Y1X4Q4JdhsZvz+1Z73vBVii6MGMWrNqSitu0j30nF
pgSgB/UYTG461/zR/FOh6sWzCBGGQnCUFB3BzqAIPOKRk5UR7EX570iK4iNJq1Gq
f/vK8Nh/nFZ/cSpuNB2jIygsDLRfp6fI+OQX21WCicMUMECHKZxhuVMYeS2o0m/L
M7OMBRd9jhP5DeQAu2jto2bm5NLVDPN/ypab58EfwheE+IHCs1UikkiQBW6v743y
17IVVW7Sb7/AjF4aP1iGhnW8j04I/DVL6TfH0qm3J9cDhnMyLEJnVeFuxFYYJtu2
5OhOOdOHA0D0TDwytdI4cH/8aT2a+Ec5k1Ky4wWKmmkSCOIgghAxBclyQNJsqH/h
xHzIxraXmOPdSvUlQ9Cq0p8TGLHXGWm+LpKZQYwTEtcmQd4KItk0ixEhCzE6+uwY
nr5bxrZQwiOAYuVKC2Z9wxeeU8L3SoRS8jBhvLu+xzIRBFaeG12WNYjaXdxwqVgX
Tk8mB9qFVm2WQwNHxFvHrrtRYVkYlhrxJlA2aetM0N14/jGIFPO2zd8GhYoNrOcu
wJKnWwYCVemj9rx8B9tNVHSJ2JvSQfvy5R7hqWEEoVQS/oRVYNHDtqVSSo8cjjr6
GUtLbJy2DwbZadNz6vS8B7ObNKxMf2z6GH91K5k7RWdFvcGzHELMXmPCw7be60EB
uhBCVd1sfX09VLYd5gF2Qg+h/yX0C+bPjM1Pvt1FpnP3DsbzxjvcuT4m0pGVbago
it87z4lhiWy3bEJdqbKBTRROyUesK24NVo6i4a6ZBUoHi6I4oL50l9hBkNCs4asq
vvyIS1F6rDSQBDPtNeJ5l5RtE21aHsJxmVUqVjyvvBejFpeRevGsNrrcj8bUmUp5
muUCsM9h6Sk7TzuKzt1LZeh42TwlI2jXOWnXmhIdJvvjaB3hrZ2d75GuQdbNLHsh
YQxFariPoeY7tKFb12fy1oV0+AtFYsT7i0PZEmP23cB9NPG4dghG/JQ2bAtxVirc
HS3b/usKSMT0yLEcKDivlQ/E2gRUlE5xMhlPr5Fg454Ht8bDLPXCx7/36iOfFjr4
MTG9aSQHxN3pec+ros1XCyq/d3hTr3f2U+VOA2gXO4AVfO700qFpFnvYvV+k8Feh
WZASzo73fO174nvjwPGx3V3QkmpWeH1fet08K599WVBlb4z+6LE941XK3jV/qOGU
Gbfdm/T5x/nei4CHOhuOdg==
`pragma protect end_protected
